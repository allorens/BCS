BZh91AY&SY�˂Vۃ߀`p���"� ����bK��         ��U!�J��H�TIT"�%*P�$DJ���PJ���(����"
�A%$��U
B�%JUETy�U)"�T"
B�QPT�UA%@���R�J��AUUU
��$�I)QU
����J�_` (��RU%0����X�I
�D� LH����BQQ"���*B*RP�(�!"E�%(AUI�G)UT
����  ֲ@�O��Z�A�5MJ i��mU"�TP��4���%(e���I�J�[V����TT�IJ$��	A^:Q@ 3��@ �à5At+  øt  8��(��s� t�]�� �Wp@�  �r��P ��AJ�)�UJ�$P ��*  ηx :=#�  ��Ӡ��P� npC�,W  �s�( i\�R �K�x  =8� ��J��"T�B�
�zI  �< :��t�4mJr�@Y�B�sG8 �Nph ��  4\�p :l1��T�4��@)uRE �J��IR��I$  �^  ���  �Wp��f���@sK���]�)C�Pl��T�Q��G��4 wp�ANe

BUH(U*��<�� ��� U���P �` (q� aER�,�F��� Q50 k@�4k� �� C�TBR�PB/)�  s�� t�� 1���� �d� � 4`P�h�'� �  ;ET���� �UzI@ w^h  (���&�F�,�� :� mQ� -SCkӇml l�EIQ(�����t�JP ��� 8Հ ��lX
 A��:ц� 5i0�P��4a,
 �i�  �EE������y�E  8� ��@����� 4ņ�Z��� mE� �`�2�  ��    � �P�� �%J�A���h S�0��MH 4    )#Mɤě�4hh�шE?���&��0M2h%<��J���@    �MBoT�RhѠ   ��u�İ�1�*������YIVJ��l��]u�=�ۇOη����@y�:�tQW� A?�D@U�PW�'�t	N]��)��*�~IDDD~�@m`<=���ٞ��&�`2ay�a�q�q�e�8Ì'd1��q���q�q��Cpa�Le�La�a�a�$Ì�Ɍ8Ɍ�Ì���'q�q�1�1��L`ƙ1�1�1�a�cfCq�1�q�q����d�d�d�Le�Ln0c1�1�1�1��2�q�1�q���La�`1��a�Lc&La�Ld�a�Ld�ld�1�q�1�q��8��Le�L`1�1�d�a�d�La�d�Ld�x�2q�1�1�1�q����Ld�a�Ld�`�L`�&`�Ld�d�d�Le��q�1�1�1�1��8��d1�q�q�e�Ld�a�Ld�La�i�1�1�&�Ld�Lq�L�Ɍ�Ì8�c0�gxÌ0�.0�0�8Ì8ˌ�Ì8ˌ8��0���0#�
���.0�dG� ����0���� 2����!� �)�
�"8�.0 c �ʎ2#�(� �q�0����8ʎ0����(��0)�E�*��2��� ��.2����aT� 8�.2)�"� 8Ȧ2���L�0��
�(8�2��
c 8�0)� � ��2�2���"��2� ����2�����0���c2���c
�ʎ2)��� ��0����*���2��
c�ʦ2���c*���¦0#��c�¡�(�
8��20!0�c��0���
8Ȏ2#�(q��Dx�.2�(�
8�0#��� 8��22��0#� �8ʎ0+� ���T�"8���ʎ2#� �8�2�GQ�82�� � ���0����&2c
&0"c2�c2�c�DLd�
�2(c(�Ȯ2+�A�2�c �®2����G8�.2����"�����ʎ0L"�(�����!�� 2�0�����)�
c���&0�0�.0�&2�xq�1�1�q�q�1��\d�q�e�Cd�q��a�\d�\a�c&e�\e�d�\d�q�����a�\a�\x�d��2�	�38Ì8ˌ��c0�1��8ˌ0�&0�10�c2���2�0ˌ�ˌ�ˌ�Ìcxˌ��c2c0�L�2�0�0�2�ǃ�<`1�d1�Ld1�a�e�\`1�q��c`1�q�q��ǐ�9=����~s�?��gz��))�_:�=1�6�n#��ƛj�#Y���U,�5@-�ֱ�� �QP`���� it2�{sK/r��� ����i��w��M�)��a4Ԫf�@Q� =��Ch^�jD��T������-XL0�d�6�G(@�j��-6�=WE�
�`�t��s���(^چZ����i+zѴSm<��,�6��w�ٛ������'�v�gT0�r�#�9��`�����mG���Y+�n�c٪m���.Kuml,m��)U�,���۶���-Ա��7��\a��\��RAE����N�cp;ܭVݴPL�b���V�F%���Z'18�j�5�)P8�ɥQ�fR��jZ��s%ѡ�%�v�$1h�
�	In �Du�a+VGy���LkeL
%HC�	Ԙ���+m�����uܠR�E����cLL���Ѳ*���f\�с�Ƌ��_f�d\n:1dBT�r� YHVM�y6�M���1�r�n�U�����"�w�YvM�m�6(��j�#ee�"�{-;�v�ǂ�j�ߞ/��+��"�錻+6�ඒ�dኳrS-H_D��D�JД���Հ��Pҗ�v�0P�bi��������Z�f�i�@��rU1��o	MG@���3F�4��I+y(̶�L����s.�E\ѫ��1SS�  ���YA%�Gj�ش��V���:�ڹ���-�XĚ� m�Ӡ�p,F�J�,Me3�3wWDB�ʅ���N�� SBX�Z��ޛ[wb]05�$�)ol��7+�F�ʔ�x%��b2
5���p<v��1�Q������l��{-��W&;��Qu�+�Én-�$raܡ����&���^X4qH$���V�r
݇������rmm �Wa:̵)h �9ueV��
��)L���䢴n��A5�,�IbP��T�ز���1��V}���NXw�n�Y��%�Z2��!��Õk*����(Rù��e�Z�t�paQB����yHn*�jѼ[�&=�غ물\�(R��B12�V,#b+j�\3�V]�q[F]�D�Deaf�n�͛n��3v�wj�^�q��k��i�u�-����k�:�kp���t��B�����N7�ۃ)[j�QS,��h�� /�N�т�!�����
Ū�Ș�i�ӱ��޳]�tۙ�Λ�`�f)���̗
��ƚT��JS��5��[�m6�ir�̪	�s)�-c[j,.��)u�oM<w��W�N��j�T��̠���t^,I�um�����Z-���ݲ�AE)���.��,�a�R5e8ʘR����q&4�=]��ݦ��
%�;D8��de�J�T3�+E`t��*��O&3(�B�e^KQ�YYX�!;J"�5�����[�����˙�Z #J#񐢥>4GVřK,�hj�^��,
�����{������Q�\4U�L�����1i!�u����n�w6��)���3+ r���M�]Ygi{t�n�g-��n���QֲS�bP����*���0�$�2Ԙ]�+T�oM���{�d@k����Ê����VQ�9X�A^wWd�b� 鵇n�K��qU��H�R
v�����R��űi����T �%-�X�� �r�Vɽ ��ӭJ��dĳ��Y�1GW.�S�[@�#�h��#�^է7X�1�!�B���Q"�t�Ў�f�a�x@T�N?�ZB�:ө���h�8�F	bV�nf-oI�s&7�ۡ��#N��^��#�[8P00��1wF���{m'E�����t���5gIL�J��s,9C�.�f˔�i* �4��.
��%(f�j�\��}��.[bOX�%ڙl-M�����^�`3���oDn�#�����0��fkij,ܘ��1��F�/pV�8o�'�	�0��	Ѝ�uNKT���=�mF�;F�-˩V-2�;�v#Xȩ����%7�\�+-D�D�$`�q��c�zU��{���Q�����2}���V*r��̷�CD.�ĶQ�*�a�N��r�̭������o
��`�*���[X�[LGa+F��3t6�c�X�G,J;���AG�k���	�M�ݭ�Z��6"�gĈ�1.�6ɻ�L��(�%,[͗a���X����W����@-���{l	N�l�DS�0`�S��B���V����Յܵu�ّ�Rܲ��`ނn<7�]��PibVl�Z�Z]�j�p�>��)�eD�Ju�_�|-n���T� �ʦ�Å�)��H�ƍ�]��D*U �ܕ�!�������ԅ�[HJV�Y4�9�fK�hӤյH��Mb.��x6VP��{��h=�O�����Le��aWV�SjK�_�EJf�ͳ-C�
����eh�q(8�|\���L�x��� �(^��[�c;le,�@;��Tخ�R�x�]E������Z�}�X�+��Y�xEZ� �iݦ+s.���M<aSaȝh�in���2�jc���d�Ɓ�'�5��݊�X�bS4H&n<ܵ��`� "���xR�l�$yD2j)�E�e��J��Q�����Uޭ�
�jh�k[���V^U�ܕ)!�wqej(�R�E��j_a3p2��c�m�Uñ�T��&ݔ�m�#,O�:��P�a2^5�i��-Z74ީdM�*ʥ�lN�Pfö�����"�39Bd.�\9wX��	u64N�%��jQ'wR���&<�2�P���]n�0��[���w�u�iB���PY13vYlP�WJ�B����vG�[9�1*�*$���������c����&�Ö�F�dş,
��hRu�'@�Cqd���)W�� Wz��� R��PB�L������1��%Ṭ��f�1��h8rB�����B��X��k@W�r���J,�J�6oᴦ\��5P��DQ�%=�P0$>,���!/n�M�w����	͔�n��x�aZ��	m�U��&r��s��v�)(��Q���2�fdZ� 'aೄS��S&�U1�{��;�r�U�yw�t,���f(sf�T���
Q�p�d5Sa:e1K�W�5��)7X�*|�*��B��Kn�m��fۙI�y
��'V)S���]���j��j`GEmbL��7�"���f�n��[u��1��"M�R��փ�LR<�O�K5�.�XJ�{Z�];z�cdR�,٨J߲�[Sޤ�+%j�z��CE� :���ѫVbeP��Q��Mв'k^+,эܻx2aZ�b�H��Ѐ�1n��x�ٴE�4�mP���uibw)�a��ܢ�4V�&�[%]���d�,I,��q-�r��F�h�k��Wkvf�8���c�shZ-hZ�f=���՚ L6Z0�I`
����֛%(�6Ht&ؠ(j&�`��݂a�6��gSA�	��6�J[���DJr k
���3�*n K/��X7��L�s_74�*�;��ѳ(������f;1�m�Ƶ�6è�E�b5
QdY[�i�9����R��
a���ј�j0��.Q��ܢ�f����eAM+mBv��m��Ӈ9���Mٚm�5����D`w�2� P�8a�R��س-��J��u��JoZf�7�ۨt=�U6�l�{���]-�[��R���i��En�EweV�in�=E��pp�����^��؂e�qauz���[��J�0��������:y5�����Nm�*���h���Z6l�r��^+��R	���^�n��ɷ[�mlh��4ӣ�6*:����$�0�A�F���o�
Uz�(JϵP�SV��:�
�dB���.=��M��l�T���n[�t]���/�MQ�w�ٗ�d�{D]����jX�A��Upæ�ʹ�U�ե��θ���QsF֪����5���aTv��`S�AmY��Z���niVsB,��Z�m�OA*���U��0XH�ö*٧@��B�]\N]�,���R�kd  TU���p$	E��;kVU�8���Z�h��V�*��K1�i$��[J��;J�@NRL:KD%�������K.٤v�a��moom���L&�v�S����)t�ƶ�&�0���6;�/V�U�Q�RG�{�#��N�ö5P˂���v�0,�sd����gE\���:M�,P(��HU��#�%��%�4��L)&�T1\�V���4텏(���b$�0���F�T�x�{v4���b�<ܭ���/t�@T����j�S��T,�jh�Kv�����}��4̕��'�=4��Mŀ޵{�anV^��L$ /K��t�I�+y�*����-��!�sk\z�$��3�QZ�J楸���mlf⡁�i���p0������J���PX��Hy1+3h�܂�I�صG.�6�d�ʆQpk4o!��w��&�wyN��>h���v�U�@y���/��kn+���J�ц�;���dj:vZWB��ޝ K3,d.EiS3�H�ȯY��ܛ�R�볋,�a�D����!�����SR�;Qn��f�L��L3kj(쪲#�x�bܔ��TM6�n�^Z�'�(&��jFh�y6t $ �;D��1�N�J�\����m� D(%�m8,cIݫv�i��.��6�S-�x��-[x�Ą�lb��}vu��f�A�����CU�=bEN�w�����!��z�
*Ɍ�m�Ad
L)�eV^6]iw��5�f�&�������"��h��,�r��œ��Z��Y@Y�Їη+ig"�MK����
Ң7{�YF`-րƫd�7
��^+�7s"�%�٥mc7�Ұ�tf�?KPfY���Oi�9iZĩ (4էt��xo5��!��z��%{B+�͠�~˧M�č�����  5gv�Me��0����S�T\@1�#�A���]<�{���`��^�s�	�ґ�0�u/]J�[�jm\ً3-��X
GM�*�43�S���7i�P��Oٛ�(أ��ⱡ���`�$۬����p���4�aX�mB� ���f^�]�����'�n�ok,m �4��Ґ&j�:.��`[wn-X㺟3r��N�|\�EW ��V��M�[�Tƞ �,��-�dجi]&�Y�(孉�-��Zܙ�SÔ�jo:�G#OqY�M  ��(P��	��Ӏb��3��tqvX��BfT�[V1�K=X�)�j,���ҭ꧉�Q�0k�]�5�K�4m�f|&�8,�T]�Wȝ�B�%�^���&�DL{r���N@s�[e�M��²�S���0o�r���n�!�f��`Mʼ��Kv�x�%���m��ݰ5�ՅaO`"��y41iISrdF�=˔
T�p��@JD�30�"�U�P�ຉԘiuz�Y[{kx`�۬i�5�i�7H5���j{�8ݭ��fOk�h�fب�]^�ͭ7Ӻ�ȥ�F���;�Rԝު�)��ܧv��&7��O��v#
N���)V�f��4�7e��P��b�x�Kb�����-�W[�P�B!�Y��ܤ�kC
��Չ�"�8��4ԶN2�-$Q2�d@��/j?�Kjő�mM�j?��ʳ��4j�z�)GL�n�
���˫�!&e���t����ěܰE�D�+b𤐢��0Sh1�*�b[�Oo0��^�5�E��hȑܧ��69%Yd��ݬt�l�B��n���%�%%�`���Ee��v�����R[�S�0`7& 3(��+�oHTl
R��6���3."[͗#��#vV,f��zj�7�2���n�VٹSX����R��-5*�a���v��Mh���dQއ������9jR�"���������l���Z�;Q��Z�v����t#��	z�!�{��j��V�R���& �JV��Hk!�km�y���MmjՋBB�ԡ���ɫ{�\F^��n�j����X��6ōd'��+�n���˷�@���%�4)m��J\��MQ�Eʺ���Ix����{7���jݚI��ْ����QR�ʾ1J��x���e�)�q��`~�u�豬���V�(��^k+w|5д\>�r+idu�8��]��C�@�aV_v�]v�'a�\d^�k�vJ�(H���n�u�����0�Q�m\Q;�p�m*aY��2�`DR�Б�B�5��aocOŧ�8�K]Lf�tt;��RH��,ڋ���r��R�+3L���Щ�q>����5��RK�;����b����l�k����f��8t�{,k߲���m6E���y�:\3"���!��
�l1��؋�w��#\+�0i��p���PWo����![���V� _�0�A\1한pq�Tc�ښ�R��z��w��v}�d�|ڤ���c�(.wf�Ōy��b��<��V�t(an��X#��B�fy}�;��2�'��3�,���t�=f��F�{9嬅lCp�)��]h��Z�7�Qx�*�a�U^ks�a<+��!�	*+YV�t�� �����u���!�m�2����J��)�уhZ��qYd�Mi\N��6Qܡ݃�+�PeJN�>�E��Ǟм�Lm��2B}D�Wݮ��7������X��ϕ�m��*����� �T{V�8�rm����ΰ�ѷ��lsr�� p��}�o�����OsC��WWD�ÖI/���6���vHK�lRZ�X{�^lc纣r���i_V����	њoQ����U�Tt쐉�w��|^]0C�k8?�]�4C�yuu�y�З��IV�v�_"e�&E1��ʋ��yd�d����|�f]9օ����:��*���Na���q&�a7�f	c?��~���+|���0}�z�D��{��+�������������𝖳p�O���;��7X{��Mv[��*�%��CF>�a[���G1����՚w�{b+m��t.�ޣ�����;-Iqv�T�ک�Vv���V).�t-�/���ׅ�}��{9��� y��gJ#�4.f>Дݓ_,��2�;?\��w�t�b�3˷zla�����=B�$�w��?]X��_t}Yk��r���+���i��5��[KW7���{&���!��hѠ�`338ovw+���JVnu��\�m^ZɂE�AW6hNK����*�2����7�Y�'�E|����v��t��rtp����^��a��V�2��e�ZLj�n�
N-���wÝ��r��it�8J��G�ٵ�JvL�!,��V2�;���1�5�5)��4kE�QW�,��Tތy�96���7guv9cY�>3�B9���VVX�/�b�qK�)�xooJ#h�7f��O-�t�wp0]v)@��
������lM�ǆ9tR��\k��-������h��Hu�8�c�g;/3#�J��D�>s���]���c�)�ufgfn�j�.u�R�N����[�5�ݽ�^Ί]�o*�:�8�i#���G'|:�]z�[������Bm�]���i��)�ݡtJ�u����F7Q;�ʦ��^��{�_\7�u�r=�k2�y+E�ӟ
ԝ��xd�*�o|>CU�eLJ�����r��Pv�|P�k*�����CY�u��X�m�厬�g]���V���\9�Di?<=ڳ���[�;�tRH��ãvV�t_ q�Z��v�O]D�Z���K%��{:XĞB�V�M���u�3�-���jgg�mY�(C<U��h���e��#����ݗQ�P�֤J���c�9����o+֏Lz�{Ѻ윐��R�k+mH��UK^;St���qUv.��2�	�PҌ�]Qs��,�"�B��1��f�pvWkT�9��n�8R�K����*ZOe<�>�� ��0�c�ս�f������QR�Ϥ(�1�=O��{U��:LB�:�f[t+
�;�D�I�j��W	�Ռ^��i��c��q���k8�t�g-\Z����=n��V57�L��@���p��X�&Wfc1.�i�v*;��6�Aͽ�݈]�r0�� :��nu8-fe�dN��7�1:E�UӐåeѼ�>�Rw+�~��=]���C���W��Q��AY	uwζ=0��ˢ{�vj�͛��oj����e�����7:8_;ʙۼ�O�V;!�Q2v
�v��I��ҍ-�	wD�2���KpUĩ����9��\��Y������L�r,�0m1�yZa�v�]:H��-�k&� �@^	Gf�����Յ[I��;v�̃�YDɘi�)���>=2���%͌�j����Q���O4)����\Heu�s㓺����۰�舀Z*r�w\ͧ�h�Ů�;�h�2g\��k�߅�O+6T�ի�f#bj<�R�t��V����`��\*�>��liC�=yϡ��R��y`;�J��90U�G��%��w6��vh]wG�����WD��]Ea#r�)�!�F�<H�Lѥ��^�L���]���-�|�#��+(�u�m�^�ڷj}�u���_1��2�>�Q:����1�[ėwX�ö�]�H�un�hHFq����ؚ]i��t�÷\�c���:!��Y�\����;q�7,m�SGR�]�E�u�V��Z�>�tbD=�ڴ�듷W5=�}��8"9ط$�6�'p�;�~͓i5VwpM<6wh9;�9gms�����1sTyv5/��A�ag^�Zy��#���v��ɴ���s7z�&4�;�
�6��8��\�r���:��{�Q���Y�P�J��7��Z[!f^T�ϘM��γ�ۓ���s�S4^�Q���\Rݤ4�h��}9i�-v�����{E��[�x+�\)Sܧ�i�r��`^~�]��3��uv���*b[}l�Y9\�����ιWD�Xޙ[��[2�r"�oG��b%��m�kː8�ɻ)k�zqM�qQ�V2z��8���m�R[��Mn
�w~�uq����ׯ��*^�Ft	ڰ�&V�)��:{V�x�u�1cOVue��}�L�	�Ǯ��%��\��ےk*Dj�E9�l`r��y�t�4�f탰�t��Z0R��Y2��;U_ZO7��_ڕt>�L�� �K;x�4jtYm]�Z��M��Ճ2�.ךX��f�+J��Wr�\�h�q5�t5���������uŵ�6�M-iu�b�;�k�O��4�yE���C��:]n��Va�Y��v��D*���ԭe:�]���W9��� �YL��(Y�&t̏���e+�	)4��P���]D�[�w\�c�t=/��{�]��-�M*�������(� r�h�w����nմx������D{J�n��XwV�L6Nz�.�$�6���M���w�3H��0sZ~pm�R���];�w|b�>��VnK�����[�\a�(�F|��������7�<*�,����(c��m�k�J)��z]�7H^�H����Ɓ�r�Kg"��V���u��P��-�:�M ��V;-�MR���<i��rs��X�9�{��S�(�.�ʽ�ji�t�wjj���Z���e,�R�� m�R�����D|+�us#��&��R��eN�+{p���$�{�B�E��l^H�l�t��%�fX��$�()��.��T𮺛�&{s7�;Ր�%t��m�G��n�c�M(l�fvˣ���`W�%�{76��-L��̈��o��l����R����\D���#��b�[B�:���V��ڀ[�uɤɎ�{�;���>�C���Nk�;âeGt���lI�Qt�\es����6��C�ǸJC/�V������ĺ�N�v����V��;K�β�͍ܮX��yGu	<C��zK;l>���-�j�B	J8��2v���Al9W����o���>��g���ھ��j2�k�DT��(q,� �JƲ�۩FZ�C��M�ˆ���
�馥K����gn3K1�X�����;S��*އ�1�r��bt�2%��e݋�ϩ���F�|�\�Savۢ��Eu�rMY�2I��Y��c7���](��\kln�� �%.�s)�2lm�,�RV��S��,f=��_Y̠r��μԴYOt�Nl��� 4V�!�msX!�;U�&^��6>�S��/
���w]�!��֋5�yd�R�W�5_L�4
ۃu����紩��R�w�b�Y;+�Q���$��z� �l۽�	�p)�'tXL�NٛtsS��r2b��Ū��Ԯ�)�8y8��'�0,�B�g�U5kx�.�-T2�6��Q���'�M0��]Թf*���v.�����Ȏuu����Hiu�;u:{�ЭS2�=F�]�i�5ۼ��pV.�����G͎F��қ��/��	�Z�֒�u|��k(r���cU�5[��0F��Qd] ;h���z͵+�5*��N���T�Mzf)8�J���K �eǩJ�ْ�o��:��#�ŎmrI�.Ձ؞��L,���&c��U�;���Ԗ��BH,7�ΝW�]W]�h�;n�^�\���м��e��.j�N!�	i��Jr�i��� e�l�s���qޢYi*�81R��ޣXS�p��5�Km]b�-wF��rwL�tA6��dr�^��#H�vP =����Y�&���d�W�i���'�l*�>�v��o���Kv&���5�������,>R�g7z�[7�U�0�ջ����úgou�Vߥ�۩����)�u�b�n����*,G@�g���SB��2��F�K����+���8]���y��+�MO_͸,��� 㠑� ���ƶ�n�d
�тN��w9�|R����zRӫt����cϡ�س%X�D�6���g�N��ɱ2j�}#@���7ɖ;l	J�zc�kMeNLMy�;���r���U��*�����bO2�ΎuclY�.�!5*�:��eޛ`uv�4�h�5 �xvS]M#Z'i������.o��T����\�4C�ա#5q�'N�2���;��^5F|\�݇���7�F$���Es���|���Ƅ����x�zt�O���u*��ڴ�¨,�H/BU�z�j��Q諼V[�t	��b̝���mY�]�k�r��3�S���Gvs�eZ��fŇGC?"��oU�v�է��:8���L��!�h�m-�a�Ի����uu8�y�4�K��թ�[ܣ�W)�
�!�m��ѫ���E�w!6)B�S{��
��vK��mAv���u5\'Z��W<�ia�
uʯ�u�R�P��e`�F�w(-���֤'g��x�y-veקbj�-xy]�J��E\ƨ�}]�[��\d�#e]�U�9��) �����i��؍@��5��͉d���-��T�;��G�rtS2`��=�5�u�}�cS�9:�+.�v�#�T���S�O�[imi���M�Gp��5-9h'xk���K�z]\<�im��we�v�|8k�\.;��H�uF�S�C�`_�޺fRR�{�P�Hz�\kz�nf��ܮ\:�wus�I��h%c���U*����s�!:��snDc���v������=F#�ő�.�N΁����G(j9��)'�YʺU�ᮛ\�;oy]|*���:��Z��e�DbSsw�9��έ��i����e.��<j�kd��޸[��Ĩn��s:�M�דk�� Y25�t��H.X�	:.�_t�-=�1�%J:B�8j"�k/�uq�ą��ܕ��`���^(u<�n�=�\Z��hR]� G^��x��K��� ��F����peu&��V�s��Eh�&(�Y��hm,�O�Pt�X]�=�j���+i�lݴ_���:��t�e
�3fs=X�W`�aQ
�ħV+�_]����;��vE���{Yk%���t������M�C��T��؉|\B6���^���n�pKΫ�U��ꔹsǲ�3-uv*Gu�f�Uv�b�ҘR�1��IG/�۷�[4�`�(�ٗ��p�V�ʐ���M<���|�Ksww�wu9��dlp�Q�F��x-�W��V����h\rAY+*�*S�F���N��]Cm^k[�Gn��M�*��U�uDw�*ꇻ��ٵ�(��
�������#��q;@+��[����^R�P��X�D�餓�7�.��t�K�����Ra����{qi@V%٭�r��G�i��B�'�Ɯ�$�ļP`�4�����y�Z������*���P���[��m���ʾ��ո����Dp��
e�����ו��]�����f��Ԥ�7��	8o��Uخ�w���'�-�r�7�_\���{��oWc֨�����gJ̢������n:H��� ��/L�ꎶ���Q׵�b]zU��Ͱ9�$K���jp)����Y�n%�Y�^S��,���ja]�JU��ق�U�=��[R�-���'Z����t:�N)�Ӥ���pZ@ý0Ԃ1g������]��y���)���9�t7{�u��7�����X��������S(LJ���/�.w�,���y�{�2�JN�ms5�S�!�")��K��g��-��\��]�{`�$'ښ����m�1��s#wI�n�7��g�W�s�ˡ�V�\��j����N�)�nl1T�����iY^�f����Z�N�X�a:}�yQj�=l鼼�O�f���]�\1,�I�aIy��h�e�jHVj�Ǫ5�.رٛW3���|�:��c�pV%R��D�+fyN[G`�Uh��(�K�Ǳ���N��9��c]���Ojv��\��y�ږL4q��ɇ�3ݻJ� �O��*�)]��c�[[O��ɹ��bUj��uo�2�����e�I9���G7S��K�nWl|W6{���۲uwN���:$�t�)�G�A�<�T����]�Һ���5�
�S{]r�/�H܂�TK�;�^� =�o��9���M�vu�s�N�ʊ�Otp�s�&��Rq����r�7p���#�F؝�Ԩϻ���;���s��݅�wwrO����׽h����oh�o�vK���d�fT�n�ʊ�Q"G2��vؚ��ctS�H��?"�|Y�ԆZ!��ʂ8%H��.��ުSҪ���ؤ�4ȠA���c���Z��uU�)
) �4m ��"�rK���9Y`|���9��ƞ�[`P�9�f����Z�,�]j=֝��U����V}��.En��L���D�-_� Ah��	w�� J����J'�ܬ���5����ME�'(o4ā3�Y�-� B�I�q�%�� ����VHR�᱙C	P�v
H	�a�B�h�q?�@�k�S��.�4�n]ʲ/�f|�YXh�DE�tA4@q$>�����Z��h�.�z�����
w��\�r����!�h	�r�_��8͘��@��b��׷)�JѦE�GJ
���9@�҉'��!��$ʐWM>0�g�,ۼ;��)� ��$�/��RX��I&����xk6����Q�B@�ڈ�LQ����).S�њ���5�w^y��vm��Yt�-��ϡu��Z�(��|��s�{����}e���5QQ�_����B*
!�������z( (��U�~������?����VA�����F ���0��'�ý���u"���^<���d����k�c���Vm��Jy����k��X	?�zS�� r�Ic���W�l�J��R=n���o\�^��*G�|{�qt�C��=۷�X�R�U���}��պtV�ӏ�Zk���r�=[��8Y���k��D듶�!�C]��1:�u��K��\)Uީ�"�P#P6��ݓ;��X��hUs�|(�nQ�eu��Ѐ��@��m;��!��26���E��b��Kl���⹍Ic�]pm������(���hLmu�
NƯ 6K��J[�6Č�,��m�+�o��Y���龜p
W%9�9-l���Gm�� �̣;�g-E�'v��n'��G^q�h�}�4aǱm��c~u�k6A��l���Z[���8�z�GK���y��z��}�ҹr�^�CG�s/T�b:��i��R�����=��fsj)�B�meֹ:���@$���K�K���ٳ��ט���+q�	N���*4�V��g'��b�����Ô�3�� �J��i]��:�ͥ'��.ur��y����d�+�ޭ�	_U�� Ͳ�k�r�:��W;��U�L%!|$DT z��-��#G=z��ݝ+��n�|��׬в��fP���W�z���׷��㎽==8�κ뮺��]x뮺뮾:�:뮺�뮺�ۮ�뎺뮺�뮺㮺뮾:�:뮺뮾�:�=8뮺�㮺��]u�]~:�:뮺뮾��u�]u�㣮�뮺뮺:뮺�ۮ��Ӯ�뮺뮺�뮺뮾:�:�u�]}|}_____]u��Y�]��O-���[��,b�Zo[��oC��h�Aٛ�-nv�Z�e��"�\�J@;�iU}1��b�y�*�IGC5�R�����ї[:�|�� w���S��c71�v�+Qꁡ/� *i���O'�^�rN��kk��x8f���έ�Qb����H`�vYf���`m��nT7�U�dYRX�q���&�����=�f���I��/�r��]ՆJ�<@	^_ak�f�krh��W���M�T��W�]U]e���d#�Sf��}���V�+\ݮ�V���ә�"e��N�A5.\�8qVG��-&��V*nQ�o6��\�֧�I:�:�s���f�4�^��d�-���E*�t�N�|qs�.�:�m��M��⡇pV�{Y��F*)�ss��ƪN�}K�-�Eى㈼8���|��}�F�(�,����Z�_mF�_:�Sz��'��wz�'z��WZ�xb��"em�E��)wrͭ��2H�k\�+���_>ţ�Q@U��zp�HK�/4�.`���B5V�	z��#��p�i�Z���!��n*���2���v�7}iFP�0��,S���&:¢�d��VF��Yh*���jVAT9V��;Y�Yk�fTJ8��m�uߜ�}�����뮳�OOOON���뮺�룮�뮺뮺:뮺뮿u㮺뮺�뮸뮺뮾:�:뮺�뮺�ۮ���x믎�뎺뮺�뮺�뮺�Ӯ��n�뮽:뮺�뮺㮺뮾:�:뮺믮���G]q�]u�_u�]u�]}u�u�]zu�_^�__^>������G]u�~��{�4Ʒ�dU݉`���[�k�}A��0�3��ںڔ3@�����A%ݙ6	ƞ(�h�u|[����vR���":�
�Ca��yP2�ǚ��yhӻ���v!/AAu愨S��]4
u�3V��5��K��k~�E�'8�fKȽ� t��6e�ңW]�&lycfK�u�Gv��>bAt.j���ж�ol;�jhd�G�̬M>w�Y��t�w\ej}o-	0|���;��[Eu���ӷ�{Pot����;q�j`���2�_Rv{�6�g[n�b�ײuxe��[��bם�k\0ٱ��.��u���{��lS$��N79Pӕ� ���6ŞoXڕ��b*"u0m<�s�5D8��kFCDRw���_�{fي)�krQ�X8_/���y�B�b�M���l]1XU|'n��q�ZGP�x0}�e'�����:���シg՛�G���e�s``.�ܩ�F��ݬ�-�t�6�fR��m�(�T��yڗdt���2'�/p�n��E���QXd��g=��T:�i}�hqU��+'&Ȯ����f�y6��zh�<��-���\�3���]o%�}��qnJ�j��j��-j�s�]������W	�53�-8��ʵ\��b�*�ˏ��.�M\~,A�G��Rc�AZ[�=������Y���ǧ]u�^�u�^�u�\u�]u��]g]u�]u��G]u�]u�]tu�]u�]u��u�]zu�]}u�㮺�8㮺뮎�뮺뮾�κ뮺뮾�κ뮺��]x뮺뮾:�:뮸뮺믎��:뮽�뮽:�u�]u�㣮�뮺���������׷�]u��]u�>u�3�7��̂�`��ں:�瘬V��=��g��Z�s ˎ�A�1`,��{%���t3��b�}�L�.Y��d�ŝe�̮�-�z�i�\�R�Gp��YY�)����
r�ջɻv^M9�VJ7ܲi\w�&�	Q M��oGA�K*ő�\pϻr
ﶚ��w�ͩB�U��
n[��n.�Xe`�G%ay�O��CQ�5��B�S�Ża���A�9WM:&vJ_>=���(4�ڝ��l�s^=XZ��u��KwT�&�r]nff�Tyv8L4o�M��u���úo�c��l�G�xؕ{���$o�v;��u����Μ��R�3�Jg2Q7&ko��L���C� wr��뭤z������P��Xs9혱(��E�����&�t\'�2i�i�o\��3%5h��im��*�BlE��j�ݕ�-�#���d���b���\/z�9ʯ�^��9�>��
:k������M��1@v���:��Б��^rL�.��]�he�� � �t�hO��1��UN�:�i뺾�w�To����t�l#��r���n��ǋ���JQM4�3�,����n�oR;��|���`�j �V��QG�qg/@�cu��*	|���.��KC?'ư��%���H�����Ct����JUaX��A�6���kh�X+���'�+]��2���:q��:gV��fP��:�s��]Ɠ��&��ٺ9H_Tٙ�'M�=ʄq>,o������K�!>�ҾR���=��\��O�Ws�mG�nt�Ի&Y/� �T���j%f�{v�����8.8�Ne ]t���4s�+F�g��o�&���<�����ޔ�ڭ*��r��p��t�f}B�
�ٓ~���;j�p�`�D�i�2�ٲ��Ĳ���L��=�P��i�T��w3qv�5_XQ�ѐ]fVm!	�D�����ĺ�ԕjq���.�n�Eϫ/C�	�;;i��d}�˩��u��fuw���S�oz�8,.V�{W������:5T�����c�}��"�+s�me�Z�U_P�����\��rwrH;?+��t@aK`�{�Up��}������8T^c�5�} �wY�i�ٯ���V�M!���	�M�9��WT�� "�{)����1��<*�
'eO�eD���zv�R���맺;��"�����ٹ��%��M� ���l�2L���6�Iy�̭�e�H����	�Թ��Y��G��K��_6�;��B������ϓPo,���=B5�*����M.��y:��W�t+b�B$eF͌2�,��z�����K*=C�Sr����u���vs��N���;{�wƖ��\ݙ�K�/��V�[�Z�V;L��؛�y��L�W&������t�����{2挰���iQ��=�k0󒪨��B����,�T�\�׳��KmnSCc�a�j�
�Jp�O���L���M]���n�댻=7��!��������ō���I/z�ٮ�z��[�;wt���]\�<�˵V���1��8�%��Y�j@&� ���v6+E#�.R�\�l�ʔJ�7j�nUg#`����r\�w�l�Ol]Gm2&ǲ�u�R5�����1M��ݘ���f��:4�};H��*��V��hi�$*��Dy���N�\ݍ���ڹF�/P"�}�B��9�9[6��|�������м��]���c9���>W�F��كٜtx�e�"�����r�ȁO(ܩz6�P\�#�8��7��<ލ���ӹYz�1�/e1�� o^i��K;ko����ulu�4��Z��tr�e�i�`*����͕�����'T%�P护J���#��Պ�.��m�������[ד�h+C�˗u�D&�8��d)9�t��]v$Da'�-@��v�n�07Gq��a�N��s�*� D'2�4�k!�a��Z��oI�Ǔ�ǹl�f;�s����P��R���>Z�Ts���o/�
���ItÊ����}����O�����n<ޮ�5`rZN�{��J{��=���pM+:;m��+3x�R��:�a�J��v�4NM5�oqJ�Y���Us��c��\�*k�_u�1Y}�@�%-�:�u��ܽ|:l�m^��z�5�c���3�|�浫)eJ�I��7]UvJ�\)���V�R����<����	�a�m�������[�, (\�̺UӎY�ۥ9LI���q��4+��6�fj��X�.4�1�c����ƀI�k��]Ƈr��y�h���׭��8FwY�3L_L�5L��v�Qr׷Y��f^#"��$�zË����x��z�`��T�:��wB����V��"��{s"�[��"�Bre��k�ݡ��j�P�W�M�t�2�l�]c~����/�]a%�Ԓ�p2-G\zt�����_W�q��s`ܪ_?�Z!i�#m��8�<�o���/u��V�GPh����h_W`wϕ�V���ʺ�8���r��͖�;�26���T����l�U���[�v��u���������+c�+��3<�n�����r��ú��#!�Q��^�h9���M�W��0ej����"�&/s4��k'e8pi%8U�E�wU��m�&(%�,*x�*ni��ׯ�����.wF���[�fe+z���7�٧ofۘ��r��j/*_-Tg�Nv�Uh�x[ɗ>�.�rl;}�^�@I\8���vew0h���b$+t�/4�7�A۷�*�_g%�0>X�y���wJ�m��<�(Y��:5�H��y��υݏ,���#�O��}c���U_V7��P&&l)p�n��y���d�\�xs�x��+�9�ٯ1X����i�f�h�2�i����#	Uкk(�H4z��I��#��L���'�X�H�B�[�0êc���[�ח.���&���f�X��.�ܧo^7��ɷ��˛AωV�پ�؍�=��fH�r��U.�c���N���%���|Lʋ���Ӄ8w��Z&X�>ЂΎ�&nSM�c������u���T�9
����k.�2�DQ���ʳmT�?:��8�m��v���x��\�(`�!�7��I��fkL�rJ�f,-ǻSO3�뺻���xϳ�͂�A6\W�hK~�XVw�f��b]A�ս%ؚ$j�"�u9���7{/����Yo^־���'N���
y��.^�Z]��"����%���q�ЮyEU˿�Vt��}���MT��U[�[m�j����%[�+��}�u,,��[��C���Xʝ�L���ߪ&t��k�5bF�`�<ʠh���לD���`�ٓ��1��{�o�D"�&��{U��W[�8��p���2�:��ޮɥ$�#�[��/�Y5�3ಒ���J=��_]�t�C�=������o�Y�u
8k3,���=�
6�p)Mզ�+�{:J��:��nd!�R����w�b��b\�[��S����i�v�5��J�"��Ě����J�wnpN2�����c�%8Ũ�9��@LVgU���n�vv��*F�F���@T"�[x�P��1�wJ,�m1�i�q)�մ�j���jl��\GL�;�)�� ��p�F�+5�}�c��&�|�W)]r�=]�C����3��q��m���ΥBڀֽkM-���e�j�M�f �L���:s2[�w��L���v8��)erq|G-��2��u'V?��g�̼Q��b�y�wtj�뽛�Pw�j��:�F��ɗ��	Y6Ҹ�s��N8e]n�dF)�ֳ)��:�ڜ��+ի; 39��V���F+���!��U�?QODC��o%p5(�&�e�to"�C��蒗JőP+ota�#mU�2�������{S�sr��W�3y�utNX�!R#����w�ԟ�_j*i�݁��j�.�X����&�)�}f�rә!����.}�D�̮p5O�oPgv�����[�RF!Hñ�>Vժ�trd?p�!7N�yF����ϸ0��z��ցn���^����w&շ��u���� T�z�)��Q���@��D����_,��9y�%W�� �,!r��D���ךּ�qZ5nB2�����e9u����)��i]�ٰvO�5Z�f�F�HB�u>�Be�t�X�><�������]an]Eף[�{�'�Ɋ�\Cꓫ&w.7.��J�&q��o�h�Q�v.4��E��\�Ly��H��;ᭊ���,��i+�iEie�pq��\Tw��"�8R�gd���w%	z��b7�C�k^�936�O]�*��p֮޶!Ȧ<��@�+n*q�[�]{�p9!�7Cb���|n*$u٭�_r��:�E�>u��$�kZ�E��E���{ 釻�-}�;2*7�c��m��OnE������5@��S/Na�P�qkheA��ӊ:/6H�dq�Vv���L�Վ��:��+�fm_��6��/��+wsu���[S�[��=�]D��|�J݅A�m�XB�N�"j�.w;+�'X����bӧwDK�ZWtc�M�`#;�� ^MK��5V�Ǚ�T����o����Q�G�������'a��ˑ� 2�ʐө�3z����̽��}S+%up]��t�]�ƹ��,����\"<'�N��z��۱�t�6��_ڌiBIK�����5mq��\����]�{�=�f���
ʓ�ѐ���LT��Z�1:ÔR��V6Ŕ�kC�v�R�(4��N�`m1GKJv����(�� ;oV���i�w�l��t.��YwX���#(���@n�*f}���?Yݝ�|%���C#�s�cι�Sh�s�Q�Y8��V�b�����v�h�[�&��8�ī�Q�:��q���q��-�OE`Y����9�lȭ��s�3�TƱ)]N�n�!�ό�4�"p�_kU�on2n�xB)��E�:��������R�B�n@���bu�Dݼ�g�cp�3�9�m#Kf�ݪN<0a!= ����dP�YpO3S���疧<DU���n5Nt��zZ"�y�hLK_eF�uc�G6����V�:7���Օ�:�%���S+�m*Z��[��hr�wyК�����9���@�|0B7�M$F̼8aE��"�t�u��n��Wt�t�_-;��q�������}Zh��{fъ�Hz��O;���T��3��|��ՇZ}�^�.���e�ͭ��䀨Q�'Qi�
�xPz��Ghs9M�w�ZY7�Q�Lev�\v��mVY�yw��.��A}"��&��-���ǻ�'S���O�w.�W�ݷ|.<�|�IU�R�t�m{��ڜ���.d��Y�7x�B��P�`��I�J͇�e�M0��	��X�4qR j���? mnx�=�6~������\2��[�;X����,Id�(?�vT|�ATN�f�ܜzq��������_]x��\�x�c�&�#���~C]F�d&[��E\Wf*�w��vq���-ά�.����ˇ.�8���oooOO����g�b7��*��ʸ�(8�B㚊)~М5����a�!�[�����==���~>>>=�?G������=��.$��.J*��˄�b�¢��/� ���_;#TVHk]5�F]���ԡr����(U�ݹ���%ur�(d�˧�M��p��:v髮��"(��jI��E���ya/G��MD92�HJ�f�D��NL艨\P2�]����c��6�$�cD���b�`I-S���K��k��Q�p�s��K�t��u��׶��&N�"��%�u�1t�aS���T�.4������7X\�k	l�5�]�v(	�5�qpM܍�؇��.��ӻul�Ӂ��r�������o��E�jnU@�;A�n��0,I�oor�x>yh!F��x��\j.s�Փ��і;���������,�`Fa<E��77J5�G(iҳqɝrR�qX���|m`�-�<NMJ����w�Y��}�\�I�|ep2�o.Az/�y��@|��_��Ə-���~^m�!�A7�c��NK��}eT��8���RV��P�O$�
�d�J���v%yլ�7$�&���ղ�.=���M�󶖼���i���/������&���z9v˞�7���{�ٟP���U��k��]H�������󞥵%�ߺ!y��2�Z����z��u�	����οt�Gm�{a�"��yK����L�lU��+�®��J�bϹ��b	l�|�}�^L�����^�������G��2���ʯx�>;����m�w���u@W��RJ��v��u{=�vV����o���+�>���އ��[�D�W�_~�k�U%u�o�0v��2t�T������ <\�^���^��a�ϣ5Y�|j�\�*����^��^�f�RR���=��Z���P���ƪ�}���yÞ�&ͥ�W�='��c���vO��J^WB�����v�6w���w���϶gK��S�Ɨ�.[t���3��V-]33`U�~���?��ۓ(�?CӶ�;��'�v}�e�W�ײvߧOpMU]m�eg��?�����?mW{����v@����&��38B`�,K`�5�x�����e���'�P�*�p��x9�.���b��5R:�%�!�����j�{�|�Mr�7>�;�J��6�p���5%�s�wy�+hu�}P�{Xٗe%[�ɫ�b��J��Ww�}D}�����$z;e�`;��=��N�{/۵X>��Ϳv�S]�}���ic�:�3I��O<�?ּ��li���l��UNm>H�V�q��n��p�B���6��0m�� 4����ݺ��[{�:��^f��ۖ|>u��_a�ՑU�*���R�*7,�Ogr�}���+}�Wv}I����;���R�zz�L�>�͹V�{H��/w�1��� ��٫�Z���|�R��6?z�����"�x�{���ǯp�ck�^BL��z����3�ӛs��w}����k���Q����Ϭ�w��{\hM=?5��%W19��T=�ѷ�SӨߊ���)y�][޽sŌr�x��L������8�C���*�V���GϦg{����􏯴�7��轞s���Oy<�_�J���ýo,��4�us�sV��s_l�@��OdfQm��#:��v���Ӗ:z/�;�
��2��G�^4��q<;�+eq�55�}mS0������~�]��tñS_	*qy���g�.�
q�n�eK=��UyumP�u�x՛�����>b�~��0�:��Vx�]]���o�a���(IN���i�];���Xx��۽IT��q�X.����:c�)�}�ǽ�2�p7�+��Na}�^7n���5���������Ӯ�m�#;\Ѻ��_T�ꇾg���j���S}��{���+�`}�Y����J�>+��~|q��}T�Y �=Yˈ���>�6�UMI�k�nyy@�����uX�v�͵�E���kWo�����U]Z�+�Î�ʡ&�ov Ǻ��m�~���6.�+��.�I0gG\�s��x.?��W��ީ�g˙�]�wv��1�c2�{�s�}���/�ثy��U�_�^��-���wglF���9�3v.����:�Fr���R�ϝqtq���k�b�5^Y�޿w!"��}�c��dпf��k����j��Ȅ��x����=��'��K��uw�r�K=\�[+�+�����j�U��o(�U��Lcq[�/���~���֫�E��#��?g�������Q��8c�<S)�e�d6o"�8�4�&q��"�����������^�*oU<7��9��մU-ŞĺX�ՋlC�<���WR�O��8�lN�f����xz.Kr�Vfr�B�@��}�U�]|�,��v,�{C�S���CJXΝlnJ9�~�{�6�b�D/�b���_?x]O����no9�z�Y��{{��!���S����?w���^պ�@Ϝ7�5m�7����*|r�������ޮ7pK�X�a�ɬ�-p�>ځ�ݓ]����^؈�" ��zh���󼭦��2�ñj�y�v��]�1&�o����9�>~Z^|u��rr������ۼ�Y�{�ͅO�޷G��iw���z�<����_!�P�l�f�����<�ػ��T�i��׽�	�,�Q�+����m�}�*�{����o^���yqڣ��|���o.��U3�ǻx������T���������Wd�k�v��t>�3����^����_?�=SO|�G�yk��s���"���s�{>s(:�&���&��Ha��ַ������`}����1?�٤;L�q���fl;�4��������}~W�b��� E;(�Kk��v�x�T������y%uiMG�8�!3ItA P�� q(���Ml��9w77N���b�|n�I�'wlu:�Іj9�q!���m�:��-���:Ώ���\�����ޗֺ�u]��|}��OR(���a"��D�4M
��(v޽�\�I�o�b���zɮop������;N�U�����^Y�z��}�m���C������҅A~�ʬ�����s4r�ߏ�>|�����m�uv�n��gu�·�f�'�����I�)w����巘17���~����\��d��о�t�ޛ�Q�|�P�2�1|��
�[���"��s�\3w���"��y�Tߧ^-��B��o���/o�{��W��YdC�5�T�,��l��[����}O%��I�/uy t1�lU��,����c��&*����Wz�������v���P�+��=��Փ��Y��	�~3�;��{Gjx�z��o�K�Rg����뽑��Ư|Gw�Ĉ6�#W���鳜=藾��f�����k����u��-��MS~�wfz`O�U�=ǻ|>s�.}�9�f����j�Q���T�����$u�n�N���/���!�%��G.�'K`��t���nh!� H�w	�M���&���k�&l]	M�/YX�_*����"��z4,÷Ա).
돀�����d�2Yt�빚`�4�m�X6��ƞ��h�;�t��`Py��}����;<=�5���]��3��C�� �F!�;���d5�sgv���,ްo��ރD>ǧ�>;��û�{#�C:��lbD8�g]wk��0mש���k��W���k���^������m{�����ѻ;S��}�c���)k�F���ܖd��<�)�K��y��:�R�|h{�wM�}���~�r��Ǘλ��uD�c{>,s�Y|����rr&�?t�՞�BR{�{�~=���Ӆ	><�1U~�nG��W�j6�3�O]�M(nt�x�eL4z���ɷ��Nj�������ũ�)��<��r��t����Y�θ;&Ǥ�]B����{W#�׽^4r���L�����Ba���{w���
Y��;�-j��o{��z��|�Ћ�7��R�G+B�C�2�x7�%�w��tr�4&@���4�95U{�:����Y��~���F�a�<�F�-��p���e�d�/J���5�N-��Xin��I��e'���U��N|��Yz0w�uPVL�L:ؖt��N�wE�+��݈1�43�"��,Kl[�e�cS�����k�	
�*t�Tw��߾��Y0��\ޣ�/Th� L��A*~��3�<�����s���ł���/�U�}�gQ�zg����j��ɧ�>��UݖNZ*�i�ޞ~p{7g.G:�OՇ��w	ȝ��P/c{*�;du���ԁ�4����uL�u��b8ݓ�죵�;�}�z�����ڃ;�}�N��+Ƚ��i���9�յː�!Z�{<��l��6i
���꼝W7B���G���O7�t�/9]�IK���y�z��]d�|3ʙ�V�<���D��|������ڸ�ٱL��R�Z���'�Ľ����Tm�>X$�����ʧ<3=�M
���xwO{��p�/Ͻ���>#�(�h�t=��y�Y�7��s��!@_;�OYI4W��8������3����xi U�u��#L�Y���sY+���o��|����_Wv۝�Ի�ϰP6o���t�ٛ'ܘ}���Z�ע���EL��>{�
8�	I�lR[ú���m�-[���4ܐ<�2��z�{]ICMsm�����c��s�`E,=a�֨^M��q��χYIu�,�U"�t�=b���#�s\�[�� ��lr����ܣ��l�Uﭔ*/4�/<����u��=�6��o�s)g�W'~���r���A| �^�S�<��w{>�Kn��v�cN��i��oKEF�H'nl����jgp�ϩ�%�۳u��%�X�q��K!���}�[�yB߁�m�,�^��yW���u��#��_Vr��	ѫ{Λ����}[yC.�'Z�p�(�~S���o������ �M����4;|FܝyO��wp��ރ�G�y��@�W�u��s�J�[�tS̝��P����w�kʕ��^z�S�<97��,��~�އ���>h������ߘg�g�����o}��=��?{ƪ?�8���k�d���t;�vG\���͸sCi��=�1U{�o���U��͏Q����K�����}��=>Z
�ϧޔ߽t(�D����yt���U"U;��f�p�|<��$�s�q�M�z�wg^����gj��ZCc;\%Д2su���Nds����y�:���6��&N��K"�)�c,�`Y�k��]�e;�s�↕ҭ�An�"��J��s����\;38�HJk5q���@�����f ��R�N��$H�P���|�ك�#Dl��H���3�����9{�'5�<�/�=6�ӊ�n]�6�x�$��y�H��O�{t��ߏC�����j.�*���<o�W�S�U;��m�1�g����d�~��<�d�ү.�kϳ�;��J﷏f3t"��w�==Mux:!}�ҳ;���������w})��-����Tޞ糨�h�}�`�C�T�/�l�ؽ�k�w�qn�W�z'�������v(w���1U~ᕍp�5F�¼�yjw�8�oϱ&&r9�z�'w��Ệ9�7~���;���\-�lY9%�<О�Kޖ>*s5��u�^���gε�+����'�M��W[���zx!6�*����͉#���
^�~�Z������^�E���7k�8���׽}���[[lEg���|2ʠ+�oy�w�������s�շ�6��h]l���9x��.�m��ѹfl���2H+�b�=Q�A�ܫ��.��Jwd<�eRDh^����8v-�eWh�YM�[�x#��e���{VnR�\���۸Į}yQ0~�`Cm�R���vZJ��̋���l�V��א��1j���ރ�S�^�)���ϸnH1ݬ)��̞�}-�t��ǝ���&Kh*�m��zr�w��������rɲ��|u#�'\ �K�owz������O�Ux�c�߸`~���t�ۂLO9=�"�_��3�k�y���j��kb_Fϰ��M�x�.�-�zY�Ϸ������9��m��㹥���~�{]�_l���j��G��_�}�7������UC��ʧ�9��v}��������߷ϡ�t�A���U�j� �y�C��[ ��v��׃=xF�w���mt��		�L��[�$\��ڙ�x�]��~#��]����>@��V<��H����W���77�.u�p��病������o/z.��^���}�>������C�����
��>�~=��t�J�'��~{��u�F�|�4��X��r#��	�d	ےn�|��m@&�͖�x���cNWJ�4�>Y2��`3o�J`����S^�g6go Og3��.]�@|��xzk�N�lڼC�]�Mǉ�@�uq�X��Z��Y�i4��s�HgB�u��/*��.0�jr�Wa�)v�CR�Ftj|{*8���Z���6����ur���y[M�!��4m��*۱"铴��C�~S�2�m�z �V�g
@䓟 �F��M���:�M��2��P/)���P��v}l��t$Ӹ{�M�5����u񺍹D�U:v�e0�c4��S ��\YԲ\g[��,h��^Ӷ�����)�L�t6�����F-,�æS��P��P����p0��J���J�0�}����V�U=��z���ñp��MN,d�Y�t�j=9�2�Zѫx�Q����K\������Xc��:�G������V���:հ�C�����֒G=#2Y��:�����Ј�a���o�>��ڴn3���ݽ���(�v�YN;��Mgdѧ&-xժ8cz�t(KZ�;�}+�(sɻ�V�-��}�R�7��
�4�n��X�-�R���0��zW q��oܫԝ� �r�=���s�%
�D�,���'S���)۰�kOz��Wj�j�'�i�.^Ӯr����[=��*�2�̮Ā8�3F�k��W^��Щ��JA���A>ձF��DD雌�i[�D��n��$�Q!���Jњ�DݔU����ok���}�9�v�������9&~�^�cM�{�7-z��@k�OOI+=C�m��7���	������4NϏ-Ȩ�f�C�D
�_EX����(�4��e��!���W<�.l�S�^�T.|�u`<�bCk$�wt�iwX����WV+Dd���Yu)���4��f���7d���X�b��1ֳ�k%�)�����e s��nB��kO��wctlN����Mhv�jT���͵sv�*d�u��u�8��o$k�HB�^R|��O.�\�y�ٙ�c<�b�V��0:*���u�+{�hڌ�ev�-�ۡ)��)0�t֋U�)Qi��rb ��>+{o�=���5z$��n�е2�;<�'':o�b�;k�|�JjW��A�7�u�E��8Eǳ��`Q�9]�����q��������d��P�������Vl�c�\�~�� Ze�Ez,�<tB�7�m������wo:Ι�<��D
_g\�V��x�AZ�=U��6M`�F0�K��[	��v��U�=N���sNs��kB�B�:h�D*r��rƜb�J�b�W�6l�F� �؂�Z��2�-�xce��J��v�k�ܮc�N�I��jX���6������'0�y냻�����Δh��cܜ�L�c�J4�Hu0�v�tC ���8r��N׫�PM������{��*�����<�./�n�8� ��U�7t���Q�����s����>gO�����Ƿ���~�x��8{&g#�%5$n��2XsSt�5i�!5!U�qffd�"�����n==�=?_�����o�����Ͽʨ������\��R������A��	q4RbeDaV}�-BR"U����x�������||||{~��������!\�s��IU���Nv��I���Û�8b*�)�v���8}�!�py���DJ�aF	h�k�X���."��-{mF��y���T���K��S�u �8K�V*⸚��
��	ȕ���d��
'��eص$q������6�Ua�������&�_���Ρf$�E|jZ��[$�\pWN"���U�Ez�6,F��z�DU�����=�l��%9���.4|ܖ�	�/%�TQq�G��%>��d�ےNX ��l**���� A������o���xߙ�׸����O,)���ǔfgV�j��oٕ�g�w�W)����;.RJ�X��3�'��:��}|�?� s�y�?_�L�8��m�8hk� w�<07Dq��ȏ����v`a�MA��(�Lj�M�fn��D������ͥ����<dC��bo軟9�p35�q��1>O<���.|�Qu��<� W3�>�9�a|@��,���n�3`��7|�"��[z����S��ކ1~ߠ�,�=�%�b���S1��n�q1VVr������0��־�F1>� Ϟ�~g���ޱsgâTz뜦���d�;�%MZ�����`H$��|GE�$� �����p�:����߄�r����}�uqc��|��y��Ƽk�_w]W�Ǭ��f�^�fO�Srn�o��8���Ug�(��.`5ᖼ�j5 �@���oQ�W���R5m��'��Yx{�E��}q�;>v~�F���?k^'�~��(�@O(�c��m�� �F����/6`��m��Ά� 4Ϣ� |�L?���I��Ϝ��+���m�dVʹ��#���bQ1%6ә]����[z��Dw?����L�:�X�җ>���ooE���v��	3ZcV�mIj�-(��u�U����v��G��1��l����	g��d,��Bwa�Z���:�G��U�9V�*��l�����X����A����Oli����%x4�1��<�d�R��"���|�wK�+A !������3{+�N�ɺI�[h��3��s�#��$t��wxi閭 ��_p�&���2�67�*U��u��S)���=��w�ϻ�D���������}|r���L8��j�|>O���i�hM�B`A���1�v8wmJb�d_,��0���Æ�ƞ��8�{���n"�5���g��5��7�ė]b�Ϻ\�<<=/�	����(- ���_���|�Ǆ��������x��� p�v���A �Y�w�E6�9����TW�F��_�  ��y�y��Xf��O��4�Df����a���=���ӄ�!ی�p�����c����'"�����Y{�����ŧ������0�|�$ap�}�#+Y��m���7�: �`r��y�%CM�H�{�e��v���u����΋�c��NY��y��������G��,fFd>cѹ�}����G[%5_�'���܂��S1�~�Q�	�y/�:�͟�|j��<xGф3�u6Q�h�𮖪�����-�E~��6�NBH-\�ZtI���8L|��,]����:��ɢ��7�W?~5Q�l(�Ɵt�i�q����h����<*q�|�Iq[q��o������gb�B�){v�ڢ��Ƕ]���z��9Bsg�ҭɆ��p�a��K�4z���N�?���N�������ʠA��z"��f=#��JD�
����$�%��d����7J��S7k�܍�@s�����vo���{\��>.4�vu�ITc�
y� ���H�ʒ�dD> 
�)�Ě5I�*-H'����[��������hስ�}uW]⋍h4�g[�nr��I.�2�.�-���@+��*�@"�iR�ңI!II����<|G�x����zu<�"�Y��X  ㇾ�`��� L���w�@�y;Z�9����Rh>F��VP	M� �n�2��8������8�yǧ�׆3����@�E��=�/��&M��+��FE�t�����Z�C�{uc[�uҬ�\��֍\y��<�L��@tvTcL�l���?�=�<l\��	����\e������L�=���E=�k�����������*�F�(��|9�|�� 3Y��k ��j :gwlG2K7ל��DR��8e��Gö��m�t�+lk�vyB������ڧlΤ�@"@O�p��(��)�:g��OW�Y	�^��qt�Wt	>���a"����]}��Ϡ������p��d�^�b#�CA�Q����)x
�޴&�&!�e�]���*��;gf�����X]��Xe��h��*ߙ���R��b! =d�if�$��Z��"\	* {�5�'���FE?{���PqSf�wl�;eD�y�Ӹd�z`>0rOzC�=M����;oG�@8�p� 슉(�P����.f�/�"���Jڤ ��/'���#f8ߏ�b�9�`Nsg��8�-�]"&6 �g%g��`Sx�;�q��7m?U��wH�{w���p�C��}�=j��E�l=���מ{ �w��H|Ȗ�ʆ�*䶵��&��#L���/�C��V�\����]"]�D�����F�ڔ�B1�ñuݍD����K���XZ���l��7���e���_���)����"�/<�w�~�}!U/x�1?���VtFx�5�xa.��3�0]��zSAle!����G��(�ah���v���Q<�'{9��{�w)��`�Y 9�eM�Y�+�{�;P�'���G��J���f�tA�|ܧ��^�md 훏���}��mdv�]?�F�@��}@Z�+�.��%��{� ���s.�L��p0@OOɤC3{�De_o��/��g�+�X���h�_*�z��5���K��5���4`3Q��G(��a�?�(�w�/΢H2�jŵJ�3�ש�1[��(p��Y���ދ>�	�P��{�$M�m�@�۵�B^�E���!��0{��]�8�0@l>%����2@\Աz(�B�ȟrp.��[ �_��
f�l�>V�wf�Fo;5�!:�b�������i]��z< (�%@�鵌�H6���E�aG�K�-E{z�'�])k١���� ���ȧ���kvCL�Jv��m���5����,l���S�0�>S�y�� �1ըk*t�>�[��$Dsi�9ցL��Q��Z�|w��f�(� ,�x�&�l��������B��X�F���Q�1U��n�.�->]c�j]�ʌN���8p7)�j��b^�����e&��w�ٟ9EY���O�7�׮4q`� ˕�sh���	�um��>7]��qZp6���rJ�Urh6;W��7yu�h罟���g��r�9#T�@�#hofvu��<��~	�w����-��9`8�wtsu�~����9�lqk\s'�4���/��t�mM�sG�l����ǅϱ�7��ဿ��:p7�nHy�D.tߟ.$61���*�u�S��T��/$�z�7��ހ,�o02�(U`ҕ`Ӽ���߼d��3���� ��>��R�3l݄<,���<���םW��_0��?��}+�[̈́xO���0�N82�|'&q��g��������na�d.^ʟ_@�����&x�{��*��ޖ������՜kv��v�a-�f#��^un����39'�H���p����>��\XI����f�
�O�,Zҽ���^M�`3~�h �k9�N��GU<x�iɊ�s#7��5:�v�޿*壧6���r3�	�b ��M��Q�F�m j��Y�
���~2�_GU�k���qm���Y��r�m��{)ܟq�)B'rp ���54�yΘf�:�U��ʜ����Ue�S�H9	�l:5���v-�w�C -_����l��
�r�g+�9^	G���j)��h��;���S��_�Х��Z4�G�~�-�nbY�����u6�L��uo!wy�Z�Ϟ�HP���}�K�/^�X�3�0j���d��]J�;���gvcÒ�J��=@�V��q�ob3�.�r�f��V�o<���ۺ�:nJ��VU�������[���ÿ����@O8R� ��|��y�{�?3������@��p8������e<�#�A��i���(�歀c�*L�����Z�V�h4�<�;��"6��Aq)�M��F�ϔ�dpޯ,�Y;+-φ�y5Y�EI�����]�a'C%�=1l�Db/��1Mp8K�FKx���H�-k�nyL���5L��vh��m�z�l7��.F�TmA󰁺��[ �C�:֐�C� q�S9Fw]����	ګxЅT7{YP�-�Ž�o"�`9]��x�:�"�y�#ç�>�O�;��!��q�8��Y�(Wٙ���T��Qj~L�Ⱦx�X�)�Л�l�^Ǐ:��@��=�1&�'��	�'�d�u�J�2��`Dxl�fm�мN�a��%��<^Fr�2\�\��0�i���߼�?��ٯ�ע��8 �=v-�]y&!]v�۪p�jJ�}ɦ�SC�G�cty8��g�`>H��{{y�7f�^p�K+�V²Aҙ���Y�2@m�em��K��ƚS.B��u,�awLؗGdH��Ü���܅ьO"[kפ@w��g�1>�&���
rj��"�y�-y���ƶSC:�kQR��ο�=�{��Ў��ՈM��o�G���w{R�����3n�8�.��R��ĩ|)��>˗d,T;E�(4�Z.Vk���#{�x\���֖�uE��f��A�9.�b�)0��:���;nu,��ە��_R9���&E��I��N_Ͼ�O���"� �Q{��V,	E�R �b	{�o�Y��ʎ<K����� ;�t���SMX����>��#�<��qd���3��(��{���q3�y�/^�%&��v[�?�]ؽ���oʼ�;/�K�U;Tz�gae{��G�!��iPڙ}��nBطf�QN�õ�K��,������V�❀���b��َ,���eR�����(�v��EO*�7Alٿ4�ݖ��x���K4,X�pkBi��2m��?�Z����7}��ќ�G���f����3�����P�����v�b]%��E[�[ �?�^�L(&�xQg��}����諸�O�2�����n�1��T�*�[5����O��r�$G��^��nȭ����s�S��PH��}an�q1K�����΀\�V6�J=�+��P���}"a��].��9�V���;��N�s�M�mٚ�r�ͬ��@m���҈���s75��X�NϹB���4[?���b�q&F��.��I��8�8�ɬ�5�.�<���jl��]<Wg�ȍ"<�2;\�'���Q=�՘|z�kSs��D��`{��lhv�&��Pa�>����r�z���z`��{-�V#eT�fܽ�%���e�\=��ntofd��s �S�q�Ux^��x�7uC
4���wz׫FwR͠�S�m�t`U�$v��-�m�s+���O�ﾯ�|*��<���*RR��ݙ�-S�C��cMЇ~oz�}b��ER}�:���Ϻ��(�%��me
��u�kz�ܲ��boc���Ȃ\2|���˕O7:}!r���a���O��T8�鷸�\��4/b�ǵ��k�v�����pq��`�Q����zkBr uO]����ڄ�X�.~�5��-�":`G��C���3m��+�c9��SY	�ɗ���Y�X�A��0�c�78�'�DI��"�%yF{����/��^t�q�>��ew'�Z�<)�����z1�E��?���վ&ì�kq�bQDމ.�Fö5�Ш�A����L��ٺ�塅%I�q�����Kݰ���X�z m.0.��n���kwI��9M�Sn�kղbC���o^rd���F���"����ac/�Q���B��a�|��O_��Q��o���������F50Q�g�3�oE@����ƾ�I�x@��{ƙu���W������W���U�W.��;�U$8b�o���*Ͽ���1d?��NM8��g�S��Rʲ����ά�8.��uN@���Gp�lX"Uo�w�g��<zʭԺVюwm�K�]Q����z���m�����厮#����)P��f�DZ���&�3a��/Z6����$��zB�AO�H�� �$@I�ϟ~y�����׵S�w�L��/��q)�|��;BUM�<��M[���r?���@=b��۾�Uro����^ H��^���dB]1�7�I�
����l�4���1L��6�-��L&,'�MK����~(��!�0�u�\����r<�m�EWf�\�.�(1Ak��/���a�	�3z�$>�}Z�=Y:�3i��x�k���08�jN:���v�a��>!�ʓ�Fy���%�s��������J�4�=�w���t�t�EJ�P�:)cۧ
�8����g��g��M��!�Y�et��T����z��be�ԙ�|6����\���Q���c��F��Y6t�S�gh�9[%rY��˚y���0���Xs���O��y��	�FI6� �]�.�=����^_��9��o|ƣg�^)'\Y�#]�F����k��;�.Eo��X3�C{iu]��< S�=�����%��8�0�N޶&��=�2�FP�q�$o'�B|��j��dB�%���� ��%G�\�)��F^7�����2�����5đ!�|�G�	 @������F�&�<2�D��R����d?N�=�X2`�[��a��B�#���X��]׻ys=��7��D�j��/$�B��C}����w�����~�8��4�w>3�Xn�j��ht�#/e]z��^�ظ��TǷ����oz�o�\���,�oT�i��8���Q�Q|[���3�A]߷?��'�"����ջ�U����	�4Hݎ$i\�@�[R�F��w�if�jvby8�P$ւ6˽�5t�wj�΋{C-��;�6:�������]�dn��&NӤ��UZ�vs�sǙ���2�O�b�1�<��3t0��MV��YSF�b)�<"-2�c�9����B9U�2�U�S/9�Cz��o�h�y LWy�ߣ����bS�5�[�Y�$ؓ�����Wpz�b�g��n������i�Lx���=��l�}%�D��E�	N�f���9�2-�K*���3E��k��P�둕잺df�jj"C�X��<�g��Q��>f5������R���!�뛨�[�9f������q���F�\��@i�Gxrz�;VL�6�vq������* �m�⎄�7[����&,���,�^�b �AP���[��室����h�.�r>��VIۂ��C����Ǭ��5:A�At��u����e;)w=#��IS�׷�lV�`v����cr�d�jV���:�%V6�r�,���wW�S0�e ���
q%����ȝ�Z �^w�쬟�*D��j���iŲ��r�7���SB�v��`TU��S�z�J��t"��;IO�v���Ӕ�/�2��%��7(��B܃����V�G,ER�7���[�@N�3�w��'��b�Ȑ�Ӎ���7�v�4�GO6�x���;������;X#:��.�,mZ�Q��ܺ�wh �R9�S�;�����.�K]0]��P��Let��Q�`4�Ÿ�N���893/Ծ짒�#��U�3�[��G�������#W���@�؅5�d鈼����"}ܫ�����V1���̺i��U��s��|oZӫ�FD�w�d�Ԙ�)�l�5�iʇ���(���q!O�(u�Bf!����Ѯ>���ou�wcPK$�b�ʜ�o`]Rn���&�.�������J�*����N%ßSa�X❷��N�2T�`���#����#1�%e����2��RFR����S�_R���U_w��_a���Z�4͗�u6�T�G%ݴU�u���sUaAU��, :5���mvM�]�i3ۋs3\5P���_
��aa��F�2f0b�!��X%�
#�t���ՠlm+GDe��%�wg6�<�V��D��J�U���ʾ�˪�:a���$N��cLR��v�,7b�>�t��n��̄�ə_�`_����P������-�%)��z��[��<���j�Erc��n�9sJe\=zxᮡ��'oEd
�������#���~�I��7���@���1$k��qmp�oV��B�Im4�sg]p;6^�A���u}/2E}6e���	a��R����P�H�꺼�3�Vi�-�Dh9L�ε��}85��h�(]��i F3z��L��:yf�R�l&�w[1��[fj���� �ᠧ��(�M�]�֓4�Ӥ�	���7i��s^�L]t7�裵�A	2��_[�@���b�;�j�t�FAkiY�<��ѨWhz�o�#BT�y[�B۾�wO(4�.� �p�0/t�0𶞱k�`���͔�뾩���oF3C}]Դ��-��h[8�u�B�^u�쵻��;����U���V��t=�q��-ʹb��xrvR%��Rf�ρ���C��}ӠX"�s\�ovYYv�Jj���u�$��Y�ͦ[�ڶ�XŪ�ܧ��X�M;�\��A轢�\��E�(��rhwӖ��Lgx|�fӡFcgW3F
���""B
ly�yaҋg]	��N!:Rs].��*V��uZ$�.V�0�&�Jod��fuɒ�;,�h�;�71�nr̩9�sF^=J_����ٻx�Cl|�4���P�QQTFR��j�e��e@�@��I�� �01C�1&6�,�H-	�Q�E#M�ЀV�r�$�Wb� RI��tUCERa�.�$���H�@���}gQG��H���U5���
(*�x��IP�����B1B��>c�vv{�ν��~����߼*
"�Z�D��(�(⧴���<�Ad�Z	RaO\�v��\b���x��������||||t~�Y���}>����/9��%��8�=p�U�/_|� ��DPG:�0������q����{{~>>>>?G�c��g�?�Q�U��J����Usk&dqDPEsqDEFeJ�TT\T\Ms]ɕ�i!a(���TUښ��d�F�3\�E�5�6�!q+��4UU_|�h?l��8���q��+�;H���}sEQWTN��=l��J*�8s�2
��F�T�㋜�¢�����AyX���㓒."PN��QCS�x��+���24�YD�~�p�1�v��q�u�\�Y�V��	��lv��UA\WATqL�u���:� ������#L}D|��JRXh���aŻ�kɇ:s��f��,)���۫m�E��\n82�Io��rc�'p�͍`�|��¯w��vje (����wn���ꋓ�Ü�s�b`d���S��Ҵ%) x����%���R��0�r�?��o�9���FߜEQ�\��]4�ב����ڛ�	�ˈ���z�T��-��q�d�� ��/����}:���5&��������vȳ+���詿kj�����A�j����&:K�q �^�rY1֯;XL1�[\�.�S	Έ��M���m3�v2�[m�ĺ�%�bW��0�0�:��@g��1w��gU�rh�R�(޲�-���ox��3�WT��:��tf���d)ty�����Ņ�c�<'����m�wq��Q�S�X/ ;���4�����n���c�\����v}�ΐE�tO��YE~�����0�]U�.�6��/C�0�>�qp+a���a��j�@�p�ּ�5QN�:��`���53����L�н��>w���I��}�Դ���YΎj�kb��]Fr����/G�\�4Nn�Ѽ`�� ��vJ]�l��ne���#�4
q���ɑ�����ۛ	n��W�ڼ�ܳ[��}]�V�o.��y
�#�GG��?��LR�����=&�t���?�4����S���iՐ���a�4*roQE:�X��Tj̈�)�W?�{���%WJ�Y꾋nn�*���B�"��y����e޸DfD^�:�!�\�s���
Eb�gN1��̛��s�4�@.zv��{k�{7�b��珺ӳ,PrQ��	܏�Ȍ2��!  �����7sS-V͖�������Ae
ƟR��>�qp�Ml��$�
�PvI�C�p0����@��N��D J��F�:�fp�Sɡ4���l*��ʞ��y¥�
r��J/��'�J��Ng��{WۦNs ���{:��w�[�����:�*$��&��ּ��l��9��&�xB�%;=�E���@�W>�	ԧH���j�!cA��cGjsm��:x��:9△'ad�k)ٓntsD��
]+_���kz�߻�y���>Z��u�o���!�B25�Άq��H$��j��F&�C�i�mr�b��S^�E�����z�y�[�-�zvvj�	}�e��c�y�4�sa��4�{��tC���$��T�ut9Vf����Jҙ=cxM�K�K[dt��y����5�9��Y�t��l�A�Q������*�v�?��*�,�$�g�#uŒ��J)�˶�g-l�������cj==*�c�] �FE�	�o����D�6*�y����\�Q=�]6{г��:�Nx`U�*n��=R��잣wO2��6+)ִz�<�9�Ҙ�!JK0f�ͮ�4I�כ��W�m1݆B��SP.�<�O��z�J9i��vӣ��L��K����C��?��G.&�Q/M�S8]�%4�ɕ���3�w��L��xf|����~��!O���QH@R+�Sky�ƙ77����4�~a0�'�v��;��\U�q�jL���0�Q��[��"��M��,�5t;͘b�9Ƶ3��Q�Sjg#Ll���J ����զ�5*2�r�7�5�0"���Z��v`! UG}@"=���yyl��a9-e���з�_^�TN)+�'<�%���f�>��WB�Z�whĭh����ڵ�x'�~�yF���q�}a������p��8�fs'��d��{�ؕ�g4-��'EŸ��������Y�e����kr:ϣ��L[Q�W��^(�j�Ȋ	L#�z�Y�i f�z�|$c{5��(2��O"�[���"�r)�.+v�G�Fy����К��O�;�.�����I&h�ҽ��0�[
�.���<(D������p�s�*4�b���GS^��-�P֛�ܭ���z�<g��s�j<u73?�\��8��'�q��u1_�lv����_�I�]eV܈�5��QC��d�9>�X��N+3�xX`2��o���1���3�+A9��;I��4d��B1�xWN���y��]]�>��8��ֹ����i�V)�*R'���ǪtP[ɣ
ł��,��k�=���%�ˊ�Λ�pɓ�����d�9we�V���dV���Mf��m�=����9Ϫy ����ʯ!�
/$�B�V�A�'�Vo(j�e��ˉ9��n0��C������d{�����Q���+�{�.g��k_Ukt?j�"^�Y����h��~38��X/�Q��|��l#�ul�Fvh�qVr���9��%���̢ħ.-�����D�=�H����s��݈��=�8�~��1�J�*�,5��żjS��k3�����_��F�!r�wk��6j�O=��+��TRf�z[-O;n�����j�n5�߀kֆl0��լ� �����(�oa���S����0{�:��W��O���;�11A'@���0�9�Ra��)�|i�'`���q��w�%�-�Z�>�2�_c�n�鶄�R>��<�z:�7�3͔��ȁ��w���cI`O����f��M:�Ӎ���v6^��ez�-����oE��t�x(�������ۼ�9���gtם�z�]^�yh�<��P�gL&}�0�=�Qa����g?�B��)6�q7U�Wf�!����Zض^�r���|˨�{Sɳ!�C��TS�->�	��)Xܙ�:f��f�Py�vDVE�V�'�$>כ;)�|rۤk����U�O�5}��"��)T��d����?yv<�}��z$��V���D��{�wd:T���oxA�t�Z�R�i��u�)�$nf�s�c�����ҫ�����G�l����9����uu�U?��eQ��"� i�|��[o�%S����T�dꇶ�o=�=�G�79M��@7[��2�K����U;�]ւ�rٝ��uk�h��C�|4�U�#���^5�b#H�4�"���ϭ���������Klr�j��(ot����u����l>�]�.I�f6E�@نu��8�D�OkD-�(UJst�@�f�E�#�I�׭i��^K�+��ʋ9�Ƕf.��d����e����	��u�/	���"~α=�1>�Z6���H���O{��=�n�ޥge���c��(��.�8�Z�w�\ӂ�GL��.���&�>t�	0��'�tIZ��m��[M��6�s�,.?��ώ�H�|Hg?:j��=*�ˮԆ7�p!,g�q���q�9�f��m�-�b���Hv�q��[��)�y�c���#�)ɤ�2ٗݻ�q�C�?��ڼ��C��!ωC;&�������3�3O��<l	\q���TO<�gNs�t�B��mntkY�Mn�eD�;L���`�0�-��F'�b�>�/dǣBMJ����#/���X8��@D���F��/n��3��F�Q� �����L���ѕ��'��[t��Zͱ[��*�;Hyw;uə��;t3ƴ+{��B�f�
���}��2�����¨�� a3����`���Gs�������o<�g�s˫����wE��?���/�
P$�EB�H"D�4�R �/������v��>>�9�a&@���}a�1{���ө�9���X[�>y�7��	�^�bv!�G-����2������q�J�H�-�C��D]�����0"��;^�#Ayn�ۗ�5�D�����چ/�QgN����f~MN�hh�,	*��sێ�L[a8l\̍c
[�h�Y���R�(m%�*���ʷc�|�Gϓ>�.{�XMļ���ꆾ͙�{�5�ŵZ	(�������+E*���f��0�~k����|�k�YΆ:���}��{;5�P�PZ�����������l^J=�uЁ�=6��*<�Fgt�S����[���ͭ{C1�� ��@C`+Z�{�W8mЈ�gLq�c����4��l%��{�,�%�Ң1��"�o(s����̙�d`�vX#��]5
]���gu)�(r����4��rC�Y~-֒�t�[̓[3�aD�<�T�w����6З�G��V�ާ�a�y�d[;��c+z����'qt��̋���_C����gX�ӯ^:,�IMu�ba�4�
k}>Ln~�^|��˷��6\/g�?O\���Ȭ.�0��ؔ��X����D��m4 �2�*�Vb��iWp]��L�{��4��זJ�T{�!:��4ڞ���2lAz�2�fB����:�"������u�E��y'j�XXz�ٰ����HeP�Q<���Ph � �U)@/�~y���f�	��{y�p��0�4��A���0�o@h&�ؓ�D0.oo��بB肯.�����,��O�fv7_��]��Q�?7]�I�T�|�.�~k�R�)�d��B�^{3��>)ƏCm!Xk*lYc�7��k^�&<���הa���Ӹe�7�y�:�RN�#y�.90�"�&�lm��13V�ͧ f�Q�`p���-�l�,�U5(�.���Fn���[Ř;�{a�bO���ı�4�Dy�rq"%��[�p�k��KP.���,�C��n�l윸Z�Ӕ�,�	��P��&��[R�"�<3�n4�3�v�2E���Y��<e&��k��]ys�=Cz�N5-�[ȑj�ݠmy���y��xmQFC��Ǔ��]��Y��DTJ���-��¹�$�C1��<�i����6}���V��=L@+Z f�hf�Gz�4�g�-.'4u:����8���#Y��݈Ee�2W2ƃiLQ��
�p�V^SH�kr�d �Զ+��1�5��\��=�6�
p���k�s"))�snR�;^Yw��G[ʚQ?���1��x����~�U"�+5����h�%�mY\Vi�a2�=��R���A4La�H#�W��{uк��_� ���T�h�f�\�ټ��,hnd�p蜲�c�6�K]uY"֧6�1���E�{x�	�"�L�GW����:�֗�!�a9�G�!H�a9"	J�
P�����6;�Nf��FDr�"}�ʷ�놬�9�(G>�O;�l1���;�7*�M�j@j�:ۍz9���_���a}c�b��Cʝ>�]��\��X�zK��Ѣ�7
ms��%���O���{S8�h���#y�3�X���[Hfd@އphU<1���ꥏ��(Q\����s�Տn�+0��|H0�O�Ă�O����Ӝq��\�pY-ECAE��H۝�X���|Do}4{��3��hbvUj�z�la�����]����k�h6���_��X�<�VGx�r���~o�����HA{����Ao�|�����G����%y��m"@vK�L��f�`��Y�]��2T�"�
dܩ�j��tԋ'��9ڹ�� �;�.D��/�. ��<`�m6!���-���w'�8�ۑ�a����UV��-�5�A##oEc	�t��3a�����g1�Jy���oV�{��SÛ]�h��i��ƻ�����C��iwCf+y��dѯ�ckY�;P���K���S'�l�L��ˬ��$�{F��RfU�]��
���P�U���r���o�r�Ti���=x�y�&[ߎ��2�X
�ؤ�F�s��ʛ�Z��{��z՛;�y-�8�B��[sJ�!����8��0VԐ�=�}.巷ܦ��v�۽�lwn��� <L�e ���BA8�41%� PЅ P�^_m�ݤn�[���>^����K�y�
h�P�Ɲ�r������O�� SK5�O��.6�6
ފ��e���I���y�]8�ԽOc1�2��IF�\A��W"m<�9���ɮh�{�p��OA4m-M��)�2���-�p4f�*�������QB��[�'ד�/+uV�u 
	\9�V���d���:l��b�N���u���V�
Y��K*jr�F{6�<!�3�k��2���	ͨ�,�L�*W����Q��C�G�79M����	�ܒӹH+j�����z���3��b�f�.�M��ـ組�����kL7��uٽ���ܭ��Q���Y��������e��v����4��%��&ȣ>ep7�����Miݧ;v0f�K5(�C��'��xG5&ju�ZkjF�]WX��V^�Ƕf8��{��OR���4�I!���,|S�ȸb۹�CBd�����{"��#-��n�N��Κ=��;��qX��:go �slO��4��!�n7'QyV3� >t�/Ʌ��H��X�1���Q�梥�mGEO��U)��]/a��Y�x�|�SK �L��<z6%*nVu�����a�e��f��EG:o��v�m"���i1��+���zTX��R�8�3��8�yu%��:4��ry�AFr�o���G�6�ͼ;��m�=���~�W��0 C=p)�R���@
>yח��޿?7������^�'��.�y�8\3ng3 c�jzDV�6���R0�#\snq�WTMU��p9��L����	��<���2p��޵��'�rٜ��kM����:�0k���!�[#+Y�3N�W��8�J5�w���]�;<��>8`5�9��v���gq�{NBx}5�B�L��|L0sq4��_���H07�]���'� ��;.�*�����y� G���i��dS��rp]?��N��Nխ�ve �oUsB�����o��	C���{(�,���ߡ�����MJ5n;D�tRxGxk}y�/N�V^�X�*}�����*	�z�E����@�oPmx3!?&�]�9�,��z��2���w0�f��n���ۗֹMs
kW.F[Q[>�",�=��s��{�Q5�ӏ��D����}��������G&�	G�u,��i�w"F����S[0�i���E�}���V�����SMn�����+�^�i賓ג����{`*롕�y.�bo�|'���>И�w����-��t�Z�g5�^%�)J�X��ovUTw��-�*�8S �gPe4��o�n��;���ׯ���8S*�F&Zv�S|O�8��2��iœ.��]��O`'���h��b�n�|���0�+v��C�(􈧐�qE�`�<��ee��K�����o�-a�v��m�h��u�w�������V���؁��S�rFo��䫬_o7Ԭ.i��۱�/K��e�Y��;���k�&А^,�� ��7f���㊌iӄ�K,�T����j��y�[o^��x!�TˣB�Dn�,�k�\7'���_���n��F�u$���� ِ�H�-�=[�,���ϯx��ŕ#�<��ph�S�Wɒ�.�`���K� � �n�v31�g9V3Uci���a�*�6�E��@���v�i��!�UJ[�;���Y Ē���4\8�д�e!��0CY}�����a��vv4WA��J:�2ʰJ���*:-���R+BN�-Lu�-��Ha�B�����	����wz��6�'���Ch������鉚L:�[<�=�g)Wji�\.�t�ۥ�L��u8k|�o;G��-))��ۮ�:��	�I�	X�5/��s�6�P���`�eJ"�52�N3 ������o��%�)
Qq�*����S8��ݺ�����丠���f(K�g,C�p�\��
�]��nR|�.�Z7�8$��r�v��ul�ݘ�Ϯ���:5�y�Jf��L6�@�J�
�.���`��	�լW�L�=EMpp��,�_%@�妳v��˕�M�Ai`���B�N-�!�n̶�z�;�7��{��Sr�~3��ͫ����G%�.2v���Q���GfJ8] ��fͱ\�y�|�����/&$�J	ff-��D���a�\C3�$�f�z���h�+��	氼|���D��l�B���/�J7�Sl�~�j����*YF���uWoD��v��cޫl�*3F���dS�Պtkpn1sN�x�_k[Wa���vx����<�2�+��>��o�v\�><3q�Up6N�p�Y8K�\�A �;8q7VT����ӣ3�lɎ�Y�U��R��cE���V�g:�S���pc��I��9x��X�¶��ɫ�ml��<v�w�CM_12�<i�ӳ����V\H�˫�ˤ����\�b�B�#��HY�,h�\T�j��bB�p<��޹k�f�@8���XA%�U�w!�/F�W�����3����
���h�)5� s^�6�,[����Ò@�3���Z�z�#�;��^_>w�|Q�d$qPD_�2�.
^�8�����3c�����m�p�*���nܓ����=\r+�x����ooo����G����=�8�񭪪/�f�c"����
�������[��݊�)����TD7�㏏o����������?_�����h�y1�u��!���[#����;�;;wUEm���q�TG��r�G���8���~����G����m��î���p�!�94)P�'��J�Yyd�~�5	1��E�,pEUI<uiW�>ﻌ(���2|�6�we�QE$����j���F�/A`���d�9 ����z���R��ys��������5G�>�U��������XUVHy��/�@P����+���b⢪�̊(#�d�}�a��눒�)9�ɬeB�3�HrNs��>�"
�����ҽ���7N��\�QpUUQ�i ��j>� *�.%yC��K%����DG�$UW�Y���嬧�2Tv���j�Ԫ0󫘹���ے� 6Omͮ���ǲ��*?e��0ΰ��w�����e����1falƅ�F9�o��Zr�r8���=��2 ��0+)���R%����}�<�]{��>�ѯ��7��iȽw@h��DO����F�� ө:��Nݹr�Y�,��9(tE�����Y�& 29�0��Z��&�Z�4�S
�Q�O�lO���,�)���o5��Ȼ�Xmn0JJ2c�3�N��د;kwt��_��싎�3�7�U���[8'7)�n�9��Jye��at�"�Q����1;��ߌ�E�OI�ڷ������n�m�Z�%om��Ƚfg�X[� ⑞�K���4^�1���H� ��8c:9�8���t)Ö���|<�U�3��	��{L(?,㋼jw/����I������4;�`Ns16Յ�s�L���ݭ���F��jb}y����z6�S�Ck�^m���J�Nt��.�u�f3��λ3q��������Ե��|�,O�|+�^O���)�-7��-vg��z��lb��i� X��kb'���tIt���1,nO�"]��"^�ޭ��z"�9�X�z4em-j�S�T�� 4J�f�ѿz��Z#<
`����/�K��xP�	t�<U�	F��� ʾ��,���HP��ݬ)_��8�"��~�{����>y��ҳ���[�ѭ�Vc,�n`X4iٻ8Gn(-���
�GƚZpj�ZU(��^n�]�	�!�չe�'x���tk�R7��v综������*���P���e$ p`@}��~����ӿ����i��ژm;��;�l��p�~0���lX��H8��=_��i�TF��vB��ap1�$�����^
>�OE��E�	]P��]�=LJ�&��2�gl��[�tn�m!��Y���:�ꝁ��n@R5���Ot�5���\�<���M�)��OR6^�y���,�Rg�$_C�/D{��b�@�B�v��ȉJa�������D�<�za�b�3�uֈ�'�n#�8�=Z)��(b :�&�k8��-l����YbN��=�o�%kQ�_�y�������ꡩ��̓��L�㎩��:���1�m�S9���O�M�ձ3�,�އz�A�.���>���ȁ���Ι��g�2,a����H�_�!ګ䃼���E��c�|���Ml�s��	�a�:Mǫ�8p����	�-��,�b���$��/k��0������K������S�ę}>�q��s�3ތ;��{[|���VOZ������ۦ�&)� m��D3�����Қ݅�k}L��;��EvPN���]I�=�&���kwwu�73S��U���|�c���.�x30~�V�=����oۥr|��!�D� x�<������E���s�Ysl�io�)�mXt;DA9�����-��z��q��-����y���{�%�,��w��i�w�A�M���[h�Hi@��%(���\�� !���)��A)��)^�v\��z�������dW��t�x_��*ФG1��1|��5�j�
�q�8�g�5r5��s�fs���
Ş���>�Bb0�w�\��v7���5�ϡ\my�K���.�:��*NOs���p�ְ��u�i�CW�<;]P,$��/�[�SG�^Y���d�g1	ѿLLY�9�(L�WUl{ �״�Mk1��N{�Q�G��6���'���ڧ������O6���0g*�!nXە�C�R����<��[yNy�F�D�O�<[-�r,X��^�
���mx�`Bt�xm����5<5�q��&9B��d�x(�7�@����K���\��d͉�:���vr����j<z�Z]%�;�������8�x�m(�m��-2��Ʌ����v��W���y�����D�=ߙKyϣ���F�y?xݷ��m���-���L�bL<�↖�͒���2������#{UGCH�L Z�{�<�6_����xn�䰥��1��y[��f�8��Ek�����׉@§j�f�9��.��A��xar���Q�r�ƫ\��?Za=�������9���m��;�|�v�%@����s���Ʒ0G5�3J}�CU���\�y6d�"�b�Y.�Z�^)WA��N�>'L��n��=9��N�o_3����|�7N�;�����d��"Q��'* ����V����iPf�02~�s�'���lߥkvx��-}v�x9uВ���]�C�5��n��%g�� 0{���X�A�l��چD2)s�V�<y²�n�6�rx;*����)����kX���Z���˚D���8�I��a�m�����{|�
���-�d绝��J4F,1PTx��{��>9R���aqMK�^ڈ=��Bڌ�;{u6���kѳf'�m3�A�I7 �f0XP ;*m�O�f��v�֎�{�b#��
�!KH��
��|�F��M0�sȇƗ��
���ʈJ+�
�g�
�+18V�>�$�f�T�B��= Vǟ׈���\�;�P0��>�y.�u��a���X�Ӻ�����Qq�3��7uy�>�K٬+����w�l%R�i�"8˲[�ҧwM�1#��s�;F0א =�M0�@0�R�,Tt��ǝ�2w\;g�ʤ6���]�sR�fAtS��f�����	f��v�'@����{4˿�N���2�b �m�en8{��2��u��M���K�H`����S������c�:i�7�Pl֋�_m�._9�fj��X�qx]��(�:޾Z��ˤ�vP�-��5���J�6�Lɛ �����w���|��\�7#�=��S�aG�p`H�P�H�J���'�2�jm�����M��;�V_�(���wv��T>��ٻ�7���%{�ɳj��MY���|oUS��$��e��^O�ܑ��i�߭d�*݊���Q���y�
�m�=����up�ɯb�2c_�n�z95��L'ɕvP�i�W"F�k3�xQ4�6�'جg��b�������ݡ���ߑ�p4�ȺQ������l^J=����2���vIn��U�igp��:
vL��h�{������k�D=�Ɯ�M��s���;���N�dMe��ѐ�t�nj.S�ʹ��'�~90�֑�M���0�/��():��F���]��ٴf�R�̮����k?�c��>���C%�O��C�0����a���<�d�U�P�f��`��Ͳ�km�����f��J8�F'p;�`p[Ho3?�>sH�|M+3�6�]��)�km���u}�\�g6侎��3�w���O1vz�8���3�7�w(8Y�2���Ԑ�ᰬ�%�EX�/�Q���i�/����˾��P�v�1nm�
����L5�Z�+iڃ��ۈ�/:&���IC��� w4V�9���5��y�����N�tBӷ�
�����y���,�l�r����٨����gp˝�]�����:l]]��i�'0���ƞ�,.��Y�F�J~o�|����3�IJ�
ҩמu��=�{����_::�3��;뇚ȍ���&�	%�0�q��u��L�<va��60u�[�'L
,���-m��z��@x��&f�a8�"�ǭ���w�|f{��ƫ���$��
�{v���5�d !�,��.�� vv��R����*L�Z��\����׻^p��6r�"�m��Y��W�6��к����c}lDz	j,�����SH��4:����SS��b�9�n��������6���q�� �zfs�X�-E��y�m��v�-:�뻚8<�K!�3�l�g�y���ꃭ5�	��(�씪�ª�˻@�'��+6]�d%��r�d��c��Xq�z�D��v�����e�S%s,h7�*� �[�0�]Eܳ=��f��k<�X��0�B.*�2֟d��/Kc�=��Zu�9���V�i��p�K.&��7g_��s����l��aFP$��u�e�:35c���X�k
�V+=�B�H�;��=��^d��E�si�5(X�hBp�=��v�\{��G���<�{�{���)��ݷ���v�:i�,����Sg�^�H3�{oSem6����uw��1idp���D�u�m]Wr�v�R��L��\)�*T�����U���e-��n���#Z�^��&�wJΥo1aC7�����z�(�9Z̡��� Ѣ�+e��3�W(���������^��� @��ws���4wIiŧ߼�l���:��Ү}����P�����g|q��a�[H�@�(-�Ĭhg̪��3��&�ίW@� N�i���:y	>�X�b�0/g��,�;���mQ��j�u�[\o5CD�{�iѹq��\y�Xތ1�f(�p�T�i��?fdu�3�"�fP��č��2��m7�6�����h5��ݏI���p3�/;ע�9n]�sscR�tAvG|	��bm�q�v��$@O|�l�R��Vb��g<�Ö��e�t7'�Ѻ*�T���k�@�:�M#��1��wcjYɷ�1p�F��ry�&�y��{SKv�G</+����� ���_qq������K�Y&���ůY˪�t�8��n��fBy�%d�՚��R�@@on��[�o�؊)K8m�.�u���1�>��m�؅ ��gxn��ћ:� ��_$��X0���8��('çO�缇3�~�c;��roj\���|��z�����_k��n�N�\2���"�Q���*\>'T�۠x�s�F�̜�ݯ�f%~B����n��R^�ʰ΅�e��-�Y��ϐ7��uƘG@2C�"ju��W2��F�J���3B��6��j���f��:<����wc���0���s';=�����֬�N0���+A�ӼVr�O�� $WdDs��_���0ȣ�B�~��Ͽ}�}��Џ�QO�x29�\��f�ӊ�%0F�d�g[O�]�ئL=9|G��9�Z;%���Z�NN�zo͉Wb��H�9�ѐ�@�M��k"�D��a�<���N�v�k[���f����a�Z���4E{���������-�D
{,���9M\'w��)����FE!��y�Z��)l���rOA��6e�#L*둕R�n����7b��(B$y��pj}�U�e @�x��C�� ,n�;K^ݰ�rۡ%��5�	�>�A>$�}Ӝ6���4Q�5D�gX�B_��� E�T(dkf�zv�k˺;<˲<ע܍��j������[��@���X�O�)����D:|֘hL��Ki�΁6
}�0��&�v�^�vy%��k���nz���n�ތ��-�3�3��M&a��{0���мr��|��Ai����쪮�a+�t��g1�Ϊ�ax��E�1|����mme�qa�B��H�ߠ=�Yze-���"�=�C��ZGc�/�\�UyJk���_ޕ[*�Q�}���}[O�V�;Tl��tL%ss>f"���k���ǅ������:u�A�Z�d\U˄5�Zxv�k�_+�;��d/,�3c�-�ݸ<WYF󭊽���B�ь�[kn�s*Τ�[��gYMi�����X���9ǧf�+�}�����!�!�D�������~w�<��������e�=>�}�9������Tq�������h�}W�ʒ���[�<->�����W���?�?
i����17M��1?�=�췚��j�S�P�\����֚<��?�'���چ0�o����vK�P��Ӣ�\�W�@����N{��fv|�[�1�g��{T[�@�{�T�D������C:�ߢ�gap�h��.��񮧗}�t��o�4[d�[3�eW���)������ؿ��\��������]����H�u@ط��#����~M���T��Q݋d㡨s>3V�{Z��Smy-�H<�xL�)0�]��b�K�>!�K���E�|jh�TXTlf�n�{��p"�Ι�7aJ9~K��+�S��qJ�Gm=C_���H|����-�ɫ���_^YQfrx����@��\��֛q�����y+{�?���P���r�����k���ag��Q2�D�&j/�ƘmkM�/���Έ���*X�5�K�ƙ�jΘŔxj���mH.����Ƌg�0�,��8�Cf��=k#�+�y���)���@Nn���t��3���Rg�S�:��2 ʾ�jsho=v2���B�\��\GR�
*vs\)_*��Z���řd��]�̸隅J��p�Q�G��J�n�i6�U���\�]n��K�}$o�C��_�/���~H<C�(�R��q$���i�Q�R�E+�"<�)��c� �X:SJ�N|'ͯ~7u�8Q�ae��ML��Uj�M��6��u��Q�B�Q�I9^�p�:t�'�hWˀ���p<�<;�K/H�a�L�����}}�w>=?xu�i�7�a���_�������wb^��uowOq��b�K�Ce��ڈA�i�5x�k4�S��9�[c�o8w:�y����Uu�;�@��^gsm]�i��� S���Qgk�9��kX�qdʗ������-cuvh�XP�.�"�1&1���ed�Q|�D[�k&�L�wͧ����f�M��Ń�Fj�i#��y ׷�K��f�3��ɨ�!�$�@�.sq�kxGCUv�0p�*Z����V�ҍf2%P�|6̬��+���(���Sֈ�J)���ɇ���ěYG#|�ewH���S� �3�)��G��t^��'�A���SM����~~��|a66,z��E��w]�%�1�5�S������[�z�(������e��ȣ���
lU.��r��L�ȭ̻2���,eH�F��)\������1cw]mխŴ1�F.���u���β:]xLi!����d��_N�뼮`.,W$���O+F�x�������aJYwһK�[�ʍie_F��#��������!f��ͨ�X'���tt��������/+n��]=9��Ug5[Xb��@f����?lS������V��c��T4	��/�jeʶu�5����6��� ���*�;?���)}wj�]���}yׯK��}��{��ߕ�죺�rh+^��R��ЫJ�lo;WM+b�bw�Fu��"���4�{>�}u��r�<@k�5Q0�A�ʰs�|��1�˸�}�P��˕,�b�ە50
u�(]l�3��c�M1y��t���n�T�ɗ���A#�ƬV�����`��t-�Ǌ����×W.�i�X�J[׫.�r����6�Ƒ50gpQ�}X��r�b��v:�l4�$^����%����u���9��w6>��ݝ��4�(��v���®PgG��5���SJ�!Ʒ�Yׄ���lRw�[�e�je*s����1^Z��u78m�RmS��g
��Vʇ���FƧwY��ٖ�31�mq��"Ɠ�3{l_Q��ä�p�)���Wh!����Vs������X�@��}��"�$��4	&��V�>l�w�L|G�i�%0Z�UjҬ���ݶ4����]*�d�ڻ06���"K��Z8�cMg�>�B�؆r� ��1�H���읇o{Fqj%D\u�e�C��##���~wkɪ���[�z�����dݮ9z�]�	��o<[�
�4A֥�]oC���P���C?h��1�Ux�2.��:�1]b]���кSr�9zʹM�J�2�Z҂�v�"`���%f�s��v��n��5L�ځ��i����ӷO�a vP}���z����1%��}�l|L��_%��[���k�Nѱ5���$D�S��s��^�m*�>�\էY7����)|���_d�{\�i8^���y`/Ew쭝,'�5�]���c����w
af��`��xhWK5T{���[���`U��[iH>�I���<9��=U��ӱ�G{��$7�b/4g�p���YC�K�r��\�w��u�6�"lm{�n��4v7�n`��[8�P���/���{&����Y�}WDM��r[P��t��|�*���
���!z!㦗w�k]�Uu؀b����X	@�=u��[[�!u�@�u�������M��5S��̈́-��(�ڛ�p���.���q@s1��tJ���L@�J�:�^5�%���R�G'\К��Iΰ����03|1����lCv`��|���8NsF�/�)4���������EA�ӡE�,�N��·�j\�*O/�J���x�]�o%n�b�*��埝���F�5Hm��eI�,�Y�a�j* 4g��᷻����}��,�d�0�$8{X
.\��
��'�+�x��i�2%���yrb�rz��8��=����__�oooo������3��B/�Hu4g#i�z��PO�$\D<�51��,���Ǒ�#/c$���?Y�o�����������~�Y�6��� ��9"�#���z�ɇf|�1ET$�rO�NxW��S��Nu�SGWW+���8���~=����G���ޣy���i���z𢈞{hxʢ2
��(}�=qNv!]�i5�Ƣ����F����#�c�`��Nz/�e�<E��(SP�$)rMr֣�&�+�,O#�9�ym���b�B�I}�؄QT$���>�*+������Պ���p�>�"�s�js}�7�h��
)�c'�k���_)oP#�9��2�S�|p�9�̛k�\�Uz�jEY̕.��BT:!:�E�T����gğ\%�VK�u�FC�1��93PԐ�<y�>y��㣒"��^���(�d'�>��x��n�>m��3=��S9,p�����N�	9"�;a�)�?S���:����m�9��Wr����}�h��#z��+$�B�L�UpW�,^�	sa�:y��6�5��г�"7�M�b�
A*)��.��S���O��a�!��U �
�T��y]V������h�GJ�U��kRa��Wٞ� �<Gs�6��+Y,y9��\�h�ǄW<�{����`�^R�p�jݕ8����;H�󸲵�[p/饒&�������9uik��pvg׷�{�}ՖҨݡ��Gg�.��]�8v_��j�����"���F�վ�r/seC��D����Cs��8ny��򅍦�	��'d�?��6�s�ՑK�J�4J���!�(�x�H�F�=M,��kCx�4����=������9��
��h)>MH��ꖡ�HN�g�L47V?���4��O�'ӫ�8p��r�1�^�}˚�/q�{9����ʘ�p�� >:ƘhL��!����&q>�m�a�s�3z0�&i=�E�[�U�-��[�W�`l��@b���3�I������>jn��5���݁�����-+Td�;ٹ׎Iv�J�ϱ�����6��Cǝ�#��s��4�m`�Z���q���u��i[�[6uLRt���4�lG��~��w�\1;=������Aû6[�r'j�M�A#�w곘.�B����EM�
�e��f)�4k�	����ɯ�eBlb���;����.���w=�zxU@W�1I��r��x���Kt�E;X{�T���qv�u6.)�����.vj�;��u�ZѺ��N�O{�����2��0������I&5�蜿�O�n���,���%�H�L:iֆl0��լ�i&�(P�vkS��r�uE�>�sH�v/9�#q:�x��0�!M4�L*kҟ5��,҃C����ñ���[�0߱� o<�v���$�[^��W�y�FhM(�j�u�m~�r/#y�k�F�g�S�u�f�OE�w|� ����f6k�j�z�&��@�i.`Ǟ���}|�Q��}�VYe6=ݤ+�2T�X��B�^��H+���u@�Ͱ�e8E���6F��kb^(�c�J��l��V6:�T�s�l��r|����cb�b����6�ɣ!����Sh-Yȹ��M��wi�en�hM'���}�#�cP��ϻ�����^�aq����`��0q|���m�DE��Ge��qo4<]X,�7 �ɻP	�ލ25�r�����*g��'�̈��0�<�-�˺1�'j��!OI��!��g(�뱱Z��se�5o.�[�7�t3N�3r3eܵ���!ΖfN�Fb/גC:�duHY"y�0s����gҊ	t_��3���f5�~�y�ٶ�ڭ=��0�<�~=�y��y�qnL���	F��X�T+v.�ʹH앳�w;C�=�?gwu`1��m_m�ۼ�/���3z1��t��Vr)l�n�i�S���(�絔�Ϗ�r囇\��<�4��S�`!���	>�s����v�?}����7��sl�����D ��Y˦\�-��2ȒGH��S�e���cwl��;o6��Ö�r��O��i�f��m�<�d��o�qr1sфۂ)�s��9��HB��t�3�u�f�
+�`>Nخ`����^[��y��p[9��j/�ow�� p�Td��>�߷��/ƕ�	�h�a��'���Z|���EJk� 7��Ô�����SM�^�4��Ey�=B�}�������-����c/N���.��<�%���w;�`�<'������� ���dW���U�8ZH7>�4r;XV�m���T1�Mh�E�F�n�DK P�vGӭ���Z|�P#�oɜ�5 h�S��WE�7���9�~#�DRYv�4�=-�(m��3R�}��4�і��G�?2+ޔ�W<�F�t�����Aڳ�w���h���W�ʹ�}��꽭{�T�gC�@�v9 ��I1�/����5�K�V,�Q�N��a��*�k�Seˑ��U���e93ʌ{>�⩩l�c3F=���̤��n�2���v���Wq�n�+DJ'ܴ�v��md�k�@s6���w�8lr�-N�a�Jޕ.���i�1>�/2�U���X���¤BPX�r��5u�U9���j�/%'s7�G�����2 �F�=�z�])-+��[���0�[7�;�H�؄�,%���C���޵��%Tl4>-PN��RU��V�a_g�0���dY�n�LC�0A��-8^f�n��>�P��j�y+m(��2��+�K�g2g�t{��-�h�!Zi�?u�����G�8�f4@���ƀ����ܛ1L�|"�͘�G;Q�O�:��93ڧ����Q��P��P������s���!��p��M�&�����	I�a��ŃYޖ��t�).�)X��$B�N���ad����:�i�v<�T�2���&�bm����L�4��&w�ck�ˁJ�O�Ѵ���OA�ä���g��XǪ0�T3J�wŵL7��D>�9s��}����n�6-��`zJ�^o�ў"��~ٯ�x��D�=_f�!����P<p>��Mm< Rl��^�S
���t9��3�y�s�&V�4�W�P��q�`�2tᙳ��Ɛˢ|d)!{�]�C`0���r)E�����5�E�1n���g�F[;;j]&�b�49v^�r��.����y�È���lm���ػ��#a��d{�(���Z��l@�uݾ��/*팥׀s�%jJ%�mhP�c�}��W�u�HӠ(�%�?q*b������vrҬ��Em,3_r�/gL�Z�cQǱ#{�u�c����ާ޺΀V�2��|#��`�l��mب���C����2Ύ�N��a!��J8}��2�S�J����a�B0,BQDމ.�Fö43 ��ƟH����D��+��R�L�J���;��4Fm����ul�0-���yׁ�0-k˰j\��r'�Ǡc�����ֲ�jO����e��K9���C3��a����R�3��^\��c_��U�ZY��:�8̔Uj٧��y��=�w��/3M�1�\T{K�P�KH��<��炮��o<�2��\<"t�	�V���)�C@�����Q5�©��{Ŋ�ҸS���=��2cY��&KP�X�*z�զ��l�֗�L���M.X�tX�m?C+3&����&fs6u�Yz$�I\#���~����*m&r�L酙��@E���:9L��1rA�Y��z�mH2�����y���)��O�Rum��;�#8�����n'uJ�%��ر��H/|U�{Y�̠M�^�@|����6���<�������6�8|s�{���� M��px���o
B�fG6�1��C�2����	���s��t8Pl��@o+z��$�8�_������Ƽ����5�����P�m�[���=�R%Ni�{�E������'�j�Z�-���X�n�ʽ1Q�ϸ9Rvܝ�gj���G0W-q�[X%�ڼ2�mⵋx�؇'�r �R�av3T�g|��-κ�?@�a� ��N�������A=E��1��R��u�0�̌�g���c�T����cOشo��DqO{?�B�;Tm�;:��i�H��"=���.�q�+��S)�Cq���`'Z�@cgSHYf��P�p�ƪ�9�UBqz�u��~�U�mxT`�� Jb^f���#�&�Y�e9�`cYJWh�su�%��*�Y�H���g���4�_l�����䮂�"��EqTB_�����<F-A�m)���E���5������o8���� ù�t�7]�Ŵ�m867oa�9UJ�tp�Wm%���{�\yN��7�H����b,��-�1P^:?	1a�����,pT�c�͓�����LS	���b�U?����f�`A��h>]��[�'T"q�w<�n��|�@O��#�]ml!A	K�xCk���\e���U���AN��f��(�o����6xܥ��1�..`����t���r����r&E��g @�õ�z�@f}a2�"������[Qz{�z]^\��Z,q)��C�&��E[U{�Ysn�h���cF'˦Ԉޯj���{��y=&�*4�>�s�L�/)��5�P�:m}֗m��s��v@ �:|�u�x���FQ�vV˳��x��ͥ�p�=af�.����CL}s�t����))�T&�DN<@�ɳwO�NY�qd��a���(	$_�<��y������~a��u��6'�g:��u��X�$�9���@���`]����E:�-�!K��Ny��	�pN_(� {Ʈz���R�� U�#:\I�W)c�}���P��fd�'�/�<`~���(3iae��(к��9ۦc�#6asu���-z�/u�����6�&`�F�fښmd�^/^jv��da+�h`u��p��ԜA�l�ͺ��2�;~���K�����ڋ�������7Qx5i4��T�,�_���7�3�TgH��&�f��[��]��A(��ٯ�w���MY�u���+��G��x�d��u�B�zS�v1�S],�:��^q}�N�����1����È����oȍt�E�7ͬXn������M�
g6��'��Y��D�Q��ǅf�;��)� o���ޮ7df������Бc�.�1w����S�I��Q�΋:sf��!+�6�n����b�%#b�A}���m�g_�}��a�G��X_��b�o�N*���m��k߸�h�5u,�s	�Ի�#�/��r{ו��VN�`�2��8��mQ9���d�{u�eAZ�����Q�Q�t'�<���_.������5[�/�[�5��r�_'�l�!�hAV���ξ q��q�^�^dA�A����И߀x�x�HC
rB��{�>o߾~{�^_�W��睠��x��8�\���7��XӞ�j��@��r�2�+��#����N�'@����W��)�Nó��[��˽u8�h����Z�(�k�Z7cCi�,���'��-�4����\����
�V~���5C`&ͪS{:r�s�����-;j&՘Z��)��n0de�=�|Л7mk8;b��B�K��ؾ$E+��Y�����O�6Y�k�L�����#��BM��yw,�9W�Y�
\YV�~])�����dy�A���eۊ����k�3j:�6w<���p��I�i��կ^Cԝ^{w߶b���&��+ιe�Z���{�5{];u���v���7�-#QR��&���XO�cܣ��$�^�a�h����g�W���_�X�X��%x�Ɯ�x�)��\ژ=�
p�����x�8ڠ�<t�l��F����Dm�d�S�j͝���2�)��.�Ur�U�Ͻ/�-�d��Ϙ��ˣ�����;��oJ]�ܽ�0����`\��ކ�G\\��M+��_����\6�Fu��(�X$�.�h�w�f����A&)���v�v��K�3��(��z��{K�f����ź�:�g[��ة���R꼨Vl��&A/w�ӓ�3K��[��c��!��DWw}�gUG]��_�2C�
z�h0��1��UK�<�/���q�^�H�t�a������q�z/�P���=����N�;�c���}ǰ?�۪^�7��R ���,�j���p�of�J1PB�0�"'u���F�v��k�fhxMQ���۶<��J9R6�O��6f��!�{^����5 Pj;��68�yWv�Z)j;�b�}B����l�o0�]�a=�v�g,���޶�y���L��a"5{�F5�/ϕx?+��Χ���n͕��r{�k�Mg��XM�͍X���Hr�8;T];^C�Ȧ����M�Jx�@wy�Ǯ�1����ARڵ��wb�� %�CW���3�Ȭg��6� ���f�,��Oo���a�b^J~!G�]��bE�zB;\�DN;��h-T;�wc c�>&�Z�st*f��pǛ4�"+�Q��T\z˄�=�K����;W<t9M�e��Zz�|���1Ou6�e�h0g3��ynK�@�%sG�������Cjk�[�_ҲH��G��޵���t2�֩֬U�r��V�@4��7�ɪ��YhM�v�0*C�E`��AqK D��Q�Y�&����A���HcT|ia��͢5��ic��wԙH�L�J1,j��:r��jr�nWUS�=�Qx�J�<>6�l���ɴ�֎b�H�9;�b�RSNb�fWPF�e�u��a	,U֧<�����z9�Ϟa��w;�y����!�x��A#��nn�Z�s|��[����G{��6�z8kɨm�d�42v�����P	�wm�������TP����V����To5y��6I�[](X�j�=�#C{�`5,��Y
#(v[GY��<�)��=�o[.����SS&}+9�f6$������k���)E�U9ګ�At9��8�-�"�w9b�5K#i���'����Y	�=D�Zj5'TN
���U�Ő��0f�tUmk�����,�S/��)�45��������0�E�^+c
�*�.�b�U��斨������C���s��"\��a��4��	L���4�iܧnWn�8�5���$�$�L�^5�?��;��F��Wo6�>��0�$a_/
h�� �5�b����&We\BBA��7�d����5ߥ�ol�?D�O?z("}��3�Qbn
w.^��VDT�_&��c�b���7�_�>�&��]ϫ3�F�7x�~(�a>��Ck�6ʆ�l|��(��_w0ܞC��UA�>��Q��t.=�)�o
����-됺X�0�4a�Ö�1�j�j^��0o����U��vs��T�꿭���VWU�m��S.�ۈ햋��dIv\���u��ED�S�[�5�a�LU��@ܻ=n_q�����-�b^�A��݊��Y]:c�_$�oo,Δ��z1ݻ���J6���܅m3�Zԓ�;�7c:����!�*�����簶U{X�yE�g�e5*c��=���h5����wS8��X��r��B����F�3֑$�OL2Zh�ڲކ�{�"n�j7��S)ҹx�5͚�q�Ek���MU٥ĕ��'l��'w�p\wV��}M�w�+��y��H��b�&n.��3_"�a}�q��+
)gWn7Xx��n����θoj -V��k���ڽ��.��m��N��2�:��0KB�`v�[�w�C����r�<�5'c%|#��Ȫ���D��Qq���֢f��[Y��ת�����7��#8�]�d��ͪ���;̢�ڛӤ��wj�k��ӫn���als�1CX����Wl�s73���d��WOeu���}j(���w/��{g��X�!�e�2;&�5|ui��r��lfj�7D�g0ZT��xz��2N�+z�q�]�o�>��s�Y:��DDo����]��1��5�7�q�[5�a���-fvJ=a#�3	R�g.�@� R�7t�s�AC���f�}crZ��<C�Pw�`��y%�yw����3�n�C;@4Z�˔)�tH 1ô
�YZ��k�p�7WN����.���,�͠���{rF���w��T=�l��镔跢P��$�YR�Jtd�{*q�&�+k+9DrUX���iX
�\,ĺ�[.�-؅���D�{��&Ieo+���Qh��.|ᠲ�^ڀ�y�U�T7cb1.�)0Y�����bֹ\�r��96�hT!LX��:�esB�Z�-�YA�L�1ѧ�&�{}�ywh���Tܕ�Q��!����NM�Mlz+QY�!̢�b����C$�7���E��.�Q���ԫ���\D\��i�)����;��Z��2�H�m�A��(�v���!���qh�NS�P��G��^Tw�� F��Pۿ�{{U��z��ծE]zv����f�|$�f=�d�{ڜ�b��Mjxúa�X؊#n�����o�',�s���ࡼ�9�N��I�Ψv⤩D˟�}1��cI`�yS������uGZ�շGQ�A���N���Q�����x�5
���I`a��YYw�[�U֡�(�.�!�-�ql�Afl��2ޝsh2�d�&�B .�Ԉ�%F��a#��)�[��d��)^�Œv�J�&ژŽke�{�Q��*����{��)�����.g�t����Z͓rƬ9�>���\��WsȜ|L�FabԜ7Zt�ۯw��g95Fs�ÖL?���������������?_�����8@�ʙ�M/�~�:��%"���D��L�ϩ�;~E��z�{���&vx����{{{{{~>?G_�ϼ��y�'Q�����!��&�(���h���((����a�Aig�G�=?_��ooooo����~�;�����7�HY�G,��c�q�9���$7�߷��Y��Σn�V�톸�jj���*��dՄ�5.m����Nɞ$8�.zǱ����"�R*-'�z���rd���2T7��W9�MML�64�����+��K�T�<���cn�$�Ŵ��]xn�"�*��ϧ^#��2����:���Ϗm��b��#�_��AW)d��55*6�S7u�E�ՑԮ%dݻ������8#����L�7�TlFI\'%@�ŕ
[	fq]�@]�ܺ. �]u�rpO�-������ӻD�7S�Dzq�iF�&v���Z��{`/,EF͸k�z;!�c]>~�C�����u��sN�|����uE���SN|mTZ�~1��4�~�:������mK/##LTGR�rrW�Ƌ!X��{t������ ?�wk��,6w+Q�5"g4R��S*im���#�=݌l]M~u��J�$��TA�	\����r�`+^<�F����,*Bp��qW���^�1N��.�S��,��s�d���-D&���(�$��ƽ�/4�Vρo?�o<;���M���`KjEp��uP������Z*�2XV��%9a#I::�d���di�ܮ')�ʹv[��q�[�,���0e1��l��F߉��3��1�!Ʈz���BR4�U�#'d�����we�-��^���C�N������y4N�1�M�;��z�(�g=�[F�c�)u�;0�Iw]y�����|���vA^s���ȸ}�'`N�l��2����/Fލ]�̇��4���҄R���V^MXM���S�~[�� �Q��=�4^u��5酩�qm��ht%j�"�n=�{5���_�;��xϖ�1�P�[""�b������r�튬k�sO[����]t�B���Vћa/��m�����kG�=���wRuaԾ�V#�hj��cy��ɹ�]�yKO�[Ns����ns������+zTZغ��"Յ�if��svN6{�{�Mz��Ϟ��n����Ϝ>t\?_��ha_�f�f��HEK��i�<�e7&�{gՂ{9���4w��+�Pо$�2j9�´���n�t�y�m2�/~#�)`6�\��Gs�i	?��S��5%�u
:Q�Z�U.����Y���0)�y�3���8b�5[8(����إ����5���w8�NW��BM|����.�v��?�~����Y;��T��/���B�!���k�@�f]��f��1�m�3��ZU����������J�Ɍڐc��.�[�督}�o�X
6�CA4�̆�*n5��QlX���r����]�g!�u��p�����S��t;[t�������].:Tj,��.��Ob�|�nb��{�O��E��[p*Es��9T��[6D���˱��߯w_ld5Y�{�K��z`��s��l��a�O�� d��t{Z�|�h,�#�����A5;90��nJk��W<L�S��|�/E�k
Mĸ�x��l��t��%�W���٭����ޜ�ت����FCQ�i2o��/��[���p8�	�ݍm��3�}E�����^4N�㝗ǝ���א�v��S�Hn�P/��\���`l����cr�����=�lf��i��U�:�t��)��"$����iv�W0nfs��u�;��"莣W����.��2�˺�\�p�8��v�V���tk��Z�� ��B%R*P�F�*3_���#��x����{��fN}��� .S�둚@�j؍:cZõ�ȭi����l�w8kԷ�b���9A]��t=,!r���ǡѽ[vyB�ΘG8:�Y�3uf�!�X��q�5����!6�����ʼ��
�xd;T�~��Jt������?��_X0X�w��N�3xY/�mm�Uu1]M3�8+��`���Gzc%<���j EX�y����6�
I��a�k�$"�h��. OSY�2�<0 ZH%�[��"y��Mo��-r�}�M�뱜�7��'T4��M�B�A�9{j�^�$��@1���)�a��I���C��m��>��kx� U�;�7JmPr��LT/RzW����@g��&
�����9�*��k>P��v٭9�R��/{m��_�^Mp+����WDq�y���Zۥ�i�* >�d7x���i\cͨ�0c!�*WE\f�aD�A:��A��7q�շ�y�G'��J(���]5�;c����1-/R�.]O-957e.�u�K���/�������u��2;��z���/u�++22n�g����niq~����E:N�:oi�N��7��vsV��x����b>l)+��WQU��p&"�Q :U�Sϛ��/���A^,�[����O�Y��	�y:��Vu����b�C�Z��]�.�Z���6W:��<�3×�/wξs��~�Og�}Ж֤
�	����l�s}c�i��"	t���ƈ"�$R5	ś�jWB����F[?w-J;�GeCwY����#��}�,FH������Ap'�����I�Ny��=U������Mb�����|ޥ�W�&�dm�;cIN�-L��.�I�2��f�~"&�q�Dw<�f�3d�7}����:��FO}){y|l��ƪqT�-���?[���^]d���F��'�nf~dF�Ͱ���W��w�z7����H��cK����]�e�[L:$��w@hͅ���6�<�i�	B���W��/�����4���|�n�T�@�!zRw��"'��m��zTYkJ��;�51�x�Ҳ��f4�����%�q4��d���9�k2���͌�ȇl�vb��S�"$I�R�� u�|����OWsaAR�%U*�۰�$b���c��r&�9/���h8Z���dj�ٓ0���:�#bb����iC��XI1�F`q�g =�.ٰ/����d�}�ף:�\+Ja��<���o��$5}�m��Q)Tf�6���U��zc��J�3���K68����w}��T���1]��0{����]u�cgJ"�;��2��ɠ�r���Tgv뭃�PK�����F��V�ll��3On�[�~=�y��$�M;��IDˡ��O��X��;��6|����m��m�?%��8ʲ�1�㝓�U��3?T������� �&��3�ζ/I�*����?�~m�$�5��!�UR��3-�0�^�����bq�M�u�~���8������4;����3�ZiL�=)����d��b�`/
��Վ�x��1�����;����C�^j���sO1w���K��޻����*��f��+Z��/$ez|�|�{�+���ٓ$�+Wkbzq�i6���ӏ�\9o�u��~:��V�{����l�[t�o�����5T=�_��Y�L���({�F�ƹ��j�{��W"m<�9�
���F�����&jZv����y���ٝͷd(�
�d`�M#5�Z�i�6,q�(�i�9E��vvZƯI�݇e��NZ���D+:{��@�m�s�V�f\6>���'G�dxM�W4F�.��L\e��T��8����g���ʗ�\V�%�iFf���j���$xvN��v�1���\?2�3Ж���ͮ^�x�6ly%㲚� ��1ު��V�]��*�[dL���T��a������(��0�r׷p8"ɭ�[��y��oCa�tI�E�]c�J䍩��Ҟ�a�k��s��D^Kk%�����`<��{��ʙx��o�R ������Dc-k����v3��f�,���̖(�LZ��Fͫ��u��lt:�ꑀ��g����%[���gZ�����I���C���_���P�»�w,��B���uQ��]R�s��������y������0~m�ht���,��1�řhЮ��APW��7ƪ��]ET�\�*�y�����>�^��%θ!��yx��Ɩ�Dp\�EC�{1�ӝ�&�ݒ,Ϻ���N�n=l���U����P�����!|	��q�������י;�C�k�_n��n��b�ʫ�G�̨������t�0Ôbs�3��3�_�oZ��P)ȱ����+̳��*�VN<Or��o��Z�f]Z��:�%���Ǘg��^,_8�1D@G@L�C������T
;�>�.�4��Ju��N�Ƒ�^�Jc���0��T5�u<hրհ =�&s�O5m
ڟ!��]LCR��;lxV�WO������8ܭ��C���[���vSo�ڌ
z1a9��v�
�r��2���:>H��$�]�U�o	�q҅ܓ��;0�[@_������Sjgv��8�m(~7�1�ѧJ��Ns�T|���2a��ܵ[|��+C�+Kh ���!�:v�;�y�Ok�so�N|#�^X�B���~� �XRɥ�_/�f ���7yL�z�6Ì�ho��z!��/t���dmj�kb�oC`�0��F˳㝪a��KԮ������^�ȷ[z:�3�t�-�5�23��$R���)�Sd,���m��-E��/��fp�ٷnrY�*$�Y�	E�$� ��TLa�kHw��BM���wU�%�!�j]oUVg"17��r��E�[Q�`��S����,��q�׫�, (o���z\�n�T?	͋՝�ew[$�J��J�u�ʱ=7���*Z{1)�ZӞ^v�>��/ї��]�r"�&���7J|_5��}�6� �0�͖��ɕ�dۭ���>f����V[d"�p���lՁ��V�SG5w8�m���\���M�:F�o&�f�aD�����&�{���5�ʇz`�ۭ�%���_t�w�D�V�|�g�at�!a��>��+�k�3�����.�xq��V� ��ck���i�\���}y~���eU�b����3����h7�����~i������0�D\C1,�kw�Qd�i�}�#*��=�L�z��}}��W)m��t֋\��II�bݰb���Y�rML��|72��t{�=	�
"��m�������g�L���_S#/����k�T��>�9�9���rz�U���b{��{W#X�j����{۝��O��$Gv�߇��{g�;���TC��m��-��»�C��6c�Rp��͂��#����9e�p��aj���Dt�ҡ��X.'��q��J��3C�l,Z�pw�p��Q\��QCr*[y��6`�}�QL��`�N�=p�Q�k�7�s�{ �tIu^z��}bX�cb��y�5��T�~�-I�.�(��oB�*ˀ歸�tŸ��w!lS�h\}R�=���ƝnNbݳ��S��yy�G�l2c�N��l���`9�h=I�=u��ގ�GyT���1�mk!W׻��eЖi�w\;��fO��ts��Ti��]�p_���4@V�������f�1�&g�ZW�k����j������7�	���"��S�ic�3zT�4R�%ݥh�ú)�a��v���\��'$r��$����Ċ�\:��,t��w�f����:+�Vcݦ���$yH6��z��mg�h�Dr�GsBSGd+�9=�N�g�@����;���		���Y�V���KRB���xd�]/�ѿ/�i��=�g��m6�ϤI�w�Nʘsgz�
f<�~={�û�k1���m�!��.o$��C(	7&5���E�Ma���)6�]�Y���j�N�ص�x�Zh]z�I���}�k��X,"����ɢ�U"�-�z>T�b���1ˡ�hhh-[V'2�X��m5n�����t���)����$Dsf5�sE��򧏷�����<������m>��[����O��D��)5�?�d��	�3����И���"L�Ydk|ɹ���k�~�۽չS���[����b�ˀű�@��T���2���(8O�ۀ�9]L�^��?KZΪɥ�R},��|�}���㞹���:6��|3�'7z8}����%�峴���B�v�V�`�ǆ[ ���BY��a�����2�}��G��������r͆��~ �Q|˹�FN��j�Kg!_���ʽq�q�8ͼ٣��>~���hȡ�DC����.����0mL���v���N�p���B.G$�-����a��gT��f9�\]�$�����mmf��]!�^��h��@&�l1� � D��ne��d_�[�[:�q�/T�^�z]��S�g�EKȦ�ŷ���+4�ʗ�N�8��Fg�C�1���"_���6��{����)����k|F�J8�;�+[#���M��#a߃�-T�h��[�����U���IZ��K����B��e�/*�:ۋ�W5�\v9e��bg<1M�jn����ui�Ot�Ժu�W*�5�zş_�}����}����ee-~�{��j�VЧ]l]p�^r�����}�Sr�ǎ��Aj������,�l�iV���7)Y�������t�Z�%6٤�)��
O��m�����F���*�ڨo���涼�<�3Y�=P7y�]�Ի��[M"��*݄.y<k1��n���EkP��I�9��V� \(��b������RY���MQ4�C�E]0,�>^K��K��$Sp2���-�xR��.�yX��M����ۓ�<a�F]�5��S�?�(3���M�Sd��.��Ō�[�2 j�sK�����m�vEi�˷m�I,#/WMY4��.Gs	���� �u�"ö�,Q�݆o5jq�-�C�m)Ra��Lh���0�Ϩ�Y0�ס��rG*��fcdI�Wfִ�#�"�F�y)F�\ʯ05�u3���/QA���er�QK_O%�nh�e�܌{f�`�'�!���՗�0�ܖ�S���kGd�[)n/���S�d�F�������i�f��������b�i�+�\�����wn��W��M��Z�-�4΁1�0�r	�vг����0���~j��/q��L���<�
�Ӗ�f1�[���M�o��-H�iz���n����3 �qߞb�e;�7�����3/{��6˭�g'�퉆����c92��=��3ם]x���k�i�ӑwک��8`9գ0�K�F�s�_n�b�F�XP��_e[�O��#���[�/3��� ���nһ���H�dԸ��Wٖ�:*ٍC`��F�I�I&��*�(�E����1� �0`�d8�rN�ro�9����r[gC׼c3�u4���w7���qƺAN�����QƗM�(򃻝���qh:�����Vi��ib��.�c��k��M93�T�`fhzF���s1R�H���J_spuu��м���l���v��W+7�2�0*7�}h�w$��N�D
�6Ч��y5𩯡�rp��Sr�ʕ��I�g#ڀ��ϰ�<�7�>��32`܇P���-o�S��m>u��JUc^��,�Z���,r�z��@.�r@i�=[n����]�r;og@E0�\E;�{Pk�9���.��PiT�U��w[�G����i���Z��WG��t��ەf0���1�,dY×ʀ�8�Q%�_VFo
����:G��];P�ss%6��t@����.N-�L�=�_>���kM�� � �6YJ��R�r��7X�WH��X�v�^��*��G7e8����>fì���oM���lt��>XY �*a�H'�h�u���u��TqVb�
�R�t�
��I�i�9����E���W*�֮�ڷ��V�+�N�XI@���Hu��[]j���A���p��j�~6xP�)nogqw�8����:��4n�;�ܤXߖH���WTXNy�2æ���.��9Q��k��F��H�F';#7�,&�+z����#gb^���Ʀ�[�է��*>�ycn�mm��Tڻ��c��K�+5� +x1p�y|�WN�u_ �Se	�u����*ҙ[��C�B�@� ���P픈�}]�5;�G2�ݷZ�>:�Y����0R�j\:1<�u5�+��JD}��m�@N�΅��zf
��BYɲ����w땹0�+5�)���}X[c�{i�8ڸ�k2�ߺ�8
TWvwpC�M�;�}��+ގa�Yxy#��j���:���r+������o�bJ��|��<�rŵy��Fsz��X�B��s3	n��@�o����z9���Te�j�P����>�V�wO�u4�0v����(Eb��
���ٻ�d�N��:7�gf�F����"��f������KY���P[�	6��2L�8��<�0`h�����wX}ɻ�|Ü��C���;4�]t�ة��!�͆����]�G����Q�u��gMJ��}�x�r�­�;�mJ��Β�ch>g��I㎸�< ���&�+Z�Q���M�ag�?w;�壐q�S��7���N<�k~��i7���x�r�͸A�D�Q�ˤ S�B��AVe)h�^�N�~o�����	����R���qsPwtG-mE�\߼^]Ows0Vs�,s�+ノ=��^�����t~�Y�}����p9�dN�
��CtO��CG��Au��'-��rMq����ns����������?_�����9�����pG9�▧6'2ABL�u͵5�@�m�����Y����������~?G������p9%o2��Eo��ɦ��oY���P�.s �[cAxƧ���3I)�N�dʍ
x���<E	F�ew�wk��6�O�k����ot�G'!�k�iz¹��Qm�ٕfI&����1A�������z�MTR��7UM{S\�rqC}��N|�4�EE1�'������u<�|y���e��wǵ£F���5�`\���͍�Hqq��Iv�'\>;�+�a�D�*���^n戼͌��j-�D�d��L�Y��3}�ul�ݟ���/��Uv̞H7w6��Q�*wK�O9ι!���ۭ���p�c���ߝ,�&�Yx�=�2&�;r�Li���6(f�$+QT�窯�Qݜ�wcv�gT?N[��`�H`����S�<^?��7�9��N��M�g�����|$��88���[V�@o��)ɣ�)7�x��:p�;׷ �xRŚ�ݷö/Uk.N8�lz��s�M:�ͪC8ÌFtQ��D<=MB�ziQA���xݙތ����"
��	�}'{��0�Q7�]����v/�k�wN�ve7h��{���f嬘�vvXZ
,�j��Ɲ�2�w@xku�L��)�Fõ�3�h�Io ^�q�<��!{�p�!�ZM�2�@��CH��Gh)�+k�dQ���%�y�3<�������SE��� ��zk��8������-��k�٫.F;�l�91����NmtK	��!�c[%����*,�v�`�B%M�6����z�-7���.��wV�~�$�h��pL�Wg�d*��˭�(^��^��[��kkL�������cֻ�v�v��%��y�g{M#��c+	G�u�ʎ��y¥��0Ȭi��c�\�d�fl�0�wT�8;��RR��el���o��5���](X�C�vX���<o�	-0��6b�����Ҭ��;�C�+�ĝו��/�!�UvQd�:���Xo<N�T+�����v:�U3U�[QF�Rܫ�GZ4֪� 
TH��G{ۘ��uַg]��ݏ�wQ��������:m@��,�9����)�p�y+Zm��U⥸��l�r�������x�<}�w�WJMs��8�ɬ��I@���a wR�"�.�)X�:D��p���Y��)r��C�r��q(��ɍ$�G0�wI����[�&qF�	y :i�O���~#.:��E��0M_Vfm3�h�����ǀ�Ӓ	d9��ؚ4Q��*�\�d���ؕB��uEŇ�l��c7j��)c���f�7���^]p2�*y�5U�ta��2��5�b�M�jɚz�I*�٦ۣ����lq����s&��<�&�y��j�����n�t��4���,Gut{�a5�j�\�0)
�o3���Z�j�@�.c�D�ǨRz�]����ؑ�t����9��5m-��Aێ����1[xը�������bNwLԄp�%����?s��a�y�e�o
��*=-N�vL�޹��7���aֻ�{��3����g�mޫo�qY��3��}Cy�&=���k_ɔ����)�Tn�6f�9ӥ��2*-�3x����)	Ff�}v�,1�x5��ή�!m���������3=���ߔؓެ�Y��0F���S�E6<X�u�#a���Vr�Wfk���o�N��)��F���s��ª���y��
\���N�i��ibJ�s.��P�s2�f���g\��X�jc{���i��*�[�U���O�)��|�JK���JyU�z����q��V�q��U����j�	���s3�3���~X�+�ԫf���jތ�h��bwD��X��3�D�<.�u��.%�-��'aZ����Ig5�ۛ�o�^�n��n��	�L��zn@.��77�A[6�sf�� ��-m=�1337�>�>Ʊ�51~�U�8i�Il�=]ٰ�͟C䦒&U��ʌw���OTv�;a�%]�䒺�uE�Ѭ�
��[���A��v��4'�ᬿ��j���E�L�$����}V���<�J��{W-Ԏ
eC�'i�+��ٓÿcb�yo��l��b��G���V_��:xM)�1����/��c^0q���o����jr�z{mۣ`h�J_��䉐���D)qo�6���jk��B�U�窠F��,k;E�r�x�c.�i`�1I;��5��y��p�Â�y�:P9�;�p�]9���ir��*��Y�0%`��:-��9��rZڼn�K&�ȶɱ3�$l�3�.� ���w�O	c��cL���l�RB�X�;|)�ѷ[4A޸�<:7�B���9���Z�4s�5ﻞZ#چ{�E����(x���5_-����G��e��%sn3=�o��m�39sP��xup3���AS���O_����#�N?Hx���ѼX�1�������/r���{6�����T�e�d���vk���qu�s�I��IsR��KE��\kOBܠ�Q|��U�v�T�&���˭�u�V�k�21���˯���*�z�O���^�)�
i���4nt����]�)�E�}�
a�5��t]�LzT��ս>�[�YA%��*���=���-�z����_tӠ٘��H��YZ&p5%vwyO�Ǔ]�U���Oϧ��iK�wN<]��|����ڰ��:Yý�=N�N釭�2y�5a�|��z�׬�:��l�[5Ga�6E�c� ����ٲ�E�]M�b&]�4��<볊���\Z!WU�u�J���瞺���ڬ��5��-��w{�vuY��Xj� A��t�? �4>������s; ��b�;6th,z��F�,���[Ⱦ�������ۋ�w,�rk���`�*O{o�`ܶ�hեY����h� L�d����QlX��v�R�⍀�+�5��w~ڕI'���O���`U��y��3.lƘc����ظ�8�̽`o)L': Z͹��Qՙ[۝f.z�l�j�w���=.��8��wW�-�[�����Zw:������Orj�������8��alVϚ��#ʶ�u+��[�>�۪'K��?gX��}��)��k@�HXL��g{��	<�וТ��\E�4�+��Q/�c;v���wJ�W�q�k��깞�F�n��M����3a�B�~��,�[�5��HI0l�]N��N}����1�X�FaݠL�ͧg�~��*���3R������T��s]Y�TF��_[k�V�$�!j6`5ư�"1�,�m��Q:�z(vR�� ��FZ�\����;Z'FS�;���f\̀�{�m�<�������i���H�Y�zVŔ���;�E����H�,�|���3(�m;�VqUL�K�J�T���u滲�v��Y�Nv�[��!݅j{�<��a�vq�+�Z�4:�g� �o^�Z�GX.5���f���D�۹o$�
]����w��h�P���觽�.�M���55r�=VwA�U�;���O�>���K[�,nĕS��כl�N^�wrK�,�2������4zE^�)^{�����clIUV�5��BLw�����+�fw+S��_���	���k��7�7ek�3�u]m���f����^��f�oP=
�fdj�W�ʖpnr�8z�M3u��M�Zn�&�9���0��"ߝQ�8���6.[�˟udb��Gy�/.wj%��2��mC�'��nR�V-�]�r����lDz��35��R,I#]�<�{�1����9�;�4V��r��Q�Lt��~����S��{�*�o��S�����hT_��au��S�`�گ��Md,�nx1s�ݘ��o�v������8�{�e�z<�ys<i(
+D���OGI�Jѻ3�fU���7W��+H;N���8���#�?W{5Pt��%�屋�A�ڀ<q��8^]�:&���D�cA�.T��&�|3B`X͚F�Y#�Q��!Ww��Q��c���Z�� c���P��q���?`��N�;+�vG�#dt�gC�Et->錞`�G>u��W4\�Wp��
����f���4t����\+���k�Qs��U��έc�c�<�%���Mu��	���䈡G���1x*�	��J��L�n�(�[��� �����xL��H:���lx1yy��Ӑ��%>=�C^ L�}�ʾ�v�ӿ��Wx�q�������f�0�ڦ$V���/4�}�ʦ��*��,�=��.#�>��3bˇS
�ۑ�]����3��~أ۱�9:�W�J}ʚ⬨�@��kVe<˂�55�a�C�o�+�z&붬[>wP�}# �2f��ȑV���X
���ÈL9S����zg�+�
�����vl�v�K=^�b-W,C�������>�z�97z]txڃyA�c�s�Y��Fϗ=�ѓ��V��5�[�1�]{�Ӏ��#e^�������m�wY�!�����yN׵x�-��ƇV���̄:�=;�Gt3�G�u�[�f���!��Ol�"vV�x���v?uWe��ո�Ǵj��y�2�s�u���\��[d�m!�]�u�Xu�:k\�ț�]�Bm�>k�WA��P��^��1�$Vn�;�R˝O��r�! �y4�� ���[�ؔ<B����U�;l�8��j�Hƶ��җ�����}X�m��rtf�&�Y�F�Y��[�P�M���ӈ>�h�F;^\�S��z`c9��m]��U��ߴ/�[��-���|Zl\��p��+�l�1c��볏>�Ǎw�����VN�)�$5�tk�>l��3�g@[���
���~j��w�	��|����/)��V���_1�+g����7����_v�٤!���&&��j�vû���*�*c��E��|�Q0�Z�<ԣ�o�1�P}ʛU��[CNcy+���@=G�S-R�^�����$Kԩ�kh[y�.���L7oMC{@�U�F�	T@�,ψ⦲n[_z3.𧖉�LF�x��ϱu��w�ĭ
P��Fa	U�y�LS�lS'w{'wj�8�$�Z�\t��z�)��A˛[�X��TR;*�k�{��闗��VF����Xc(����D��]$M�����Ί��������NWZ$j��9��3!l�H��z��ކ�r���y���K]؆���M��J"��\�ؒn���K��`?D���~�NhN��u��H�M^����t��mG)��n�1騫�;51�b1�roab������@�މ�	P0�Zݝq��`�;KG^�Ȼ���Et�v��F�K��D��t���lxS�5��X��M�W��m������Lm�nIv���6�|.� �� ;-�ҭ��n�U,l;�^]M�w7],�.�]C�+1q��%��vNj���[Y��P���~>w�ٍi��kf�]1wY��f-��Օ�:Uֺ���^�2;�X�ݐ�ř�<�V6)�v�)ݾ����B���C�E(��zZ�X�m����
qnX`�h�ButZ�9�<��,ǃ��oF�V�l\�TY�f�+^~iM�h����	5yPй���5��`Sn_n�蔇u�N4��-��p*�"��lS�[�9�.�U�"���96�s�4��e���͕.����=Cc]*T�u�S&�x��;쩰zC�"���w���ȭY�S[0�/Z��d'�$���t�7�k��h�bO6q/n��7�C�*��ӎ\	γ��E���7iY/6���U	�9Y���(j�,&K].�8�dw��g;*�q@g���m)�V�E/�:����.,Ai]X��j��H^�yEX[l_֥� ���v�v��m�H��̵ͣ4��a��Ĕ�ބ��I�q{���a�E�7YLF�We᷎,���ls^Bf�*������ ���ےŚ��私$�;P�ޗm���U��z����y����iۺ�
U�L�*�ૡ�)��w>m׆n��=�)�d�xg�0�U�nZ-[pdY��A�L٫��٠=W�vQ^��گ:ew,��]x�46]ǌ��j�����O[v�wpk~�q��vV�q�Ԡf�oW�o�e-���Y�Zٰ�K�dM�}�f{�nz���ſ].z���X�ܷyW>��f�wS4tpW�5]חV��Ӣ跙HpUǶ}���x�F-�Vˀh��h�8գ1��N�kF=ؙw�=�zG9!l멙P4�Q��y��:��e]\��ղ[u6�'�.�4n�V�-�6��k�r��l���n��ؚ�k'(ui��x/�r�P5���s�v�uc�N���),��.v6�G5���5*b��HE��a.v�	�r�J�҃
U�j��9�-tjcSn�4�����r��=�}j]��=�b������*�opa�iΧۆ����k%.T2ڥ�s�K��}�x8*�'p�5�[N'1ϖ�匰�qP_
�:�uL��4���{�5�/D���ꕔ���4wu���E��=DAegm���p��1�8W�yf���j-ЋI�^pWq�I����]O3<4���{��d����p-)b	�(��&c��ý_l��C�/��T��$%��9[X ��Ʈ�]4�s켕k�P�v�}I��-���0�f��7�4iy��
/�p�I�sj]��c�ٵ\{{��[Tl���ܡ�����2�@���^�)z�N'�`�OZ�.�� ����}k^nNߙ��m-���|
oX��,��ÌV0������(&>��ܡy��wjKZgsSw�*�8�f�g|����:��c����oh���r��eO"���o��,+�j�ַ˰���E�iV1,ȟ�UԖ�YP�*ڜoo�!�,�Ո��L<�ib��op��pȇXj�*y7�d�obƏ���W�!�t��5+����U��ƫNe]��	�Ҫ
B�(-��&ڦ����R���R���p�����Qy�τ�5��3�.9u�y���R�u9[G� �h��&��*�Y��W�����a���h�6����X�b��ȏ��y~���M��2HspCy��7E���z�*%-�]])�¤J�-���l�uz�e갻�鑰 �P�}��$�)��
�S��\T�"�7������巼Y���Z]t��	o2�f�m�F�Z/�"T�S������d�$��fVB9�yr��;�1n�R9�Fo�Pop�v��Y�fN�K.f�_v��,v^F�����iTw{�^�wqYQ<�R�UәI�&h}x)↦o]H�<�M�)�ƀQf�<qh�3�hH2��n�Χ�dݡ�^7�C{�h��h����0'GF�C5�0
G��X�����>�8!�j�!�^ͻ��Ha�8�E��q�Ŭf�+�ju�PN�Qq�쥠�2�wҐ��ͅuw����sGA��yMF �!W��(j�
�(�Raob!�t�I��m�<͋CkK6s>\�7���Պ�9��a+k-o��J[��&�O/����{�4��E����!얩�m�O1���u��1�Õ��ۣ���HXdma�TJrS�f�٪�������3��{��d�ҝ�l�Ϋ��9>}�2MΏ�}Ϝ�Ű��z5���W��m��ԣ����#�p����x8j(:��H���9g9˜���zz{~:������~?G�?����3���jJ�[	��ڮ#����� L��!��}��S�9^Q7}u�������������t~�Y��ӏ�,�.s�{ud����p\�Z��`Ԝ�Dm-w2M�\re/��,�s���ϯoOOON�����>���ڞs�\�s��)-F�nPGw<�s���Ӑ��:�BI��T8�9�k��i`�Ib)�.wvn|s��\.�j�Z)��Ҝk,�<�׶F,����zb�1s����Q�Rn�u!s7t73	��W>�wkbC�8���I8�^�>�&�!��,�E[��8(~I�63� x�k8)������CgQ&B��ֺ���*Q	6X�&鹸���~Ms�l�,Ȟi���F�k$��������҈�eMC�"���ऴ4B(�"���(�>��@��o^m�ޣ��t��$��]��̱�t���+��
'Eռ���n8��{��9/��
h��h�z���}��Ȟ��m�忇a��x��05��Y��B� �j���Ģ��~����5�Ǽ�)����n3T�Og{�d��6�8��ՃZ!T�1�/��L� l�qw�ޘ�^�y�s�>��"6|VS����R��^���^Bt@)V�z�2�k��к{���[�����C3a믻CL8�M�P3��H��c�{�:��>�6%9�l�h�J�\(����1L�Ü㖠�N'uɞ�glM�Vw=�Hu��c�\d�>,�����ǅܲ��j=�Y�j�o�0%R��Lr�Y���јڽ����%��Z�о"��~��0׏j���Ϫ)�<�Nd�j���UTJ�3`�OOw;Y�&��v\]����uR5R�	U�ڦg�f\��7�}zV�xV����M�:fn�i�_�l$�:�닁�iHޅy��k\_6t^o�aHc����Z���W8��� 7���f����{*�FP���N�J�D��Uj�>�m��P��Ǉ�����`" �O���R���v�,;)vZl����N�=7���8Ǯvr���g�d���D�6�q������vջص(zo}e��ٽ�l���*Ud�Ԓ�i(�U�ay�w[^��s�����@�ʤUy�9Ю'��I����׸v#�]6��k�������`4�v�uV�j|��x\�c�_��B�b/V�6�M32�����:����۷��|�8v�z� ��js�\�C���]���i〓��)s����Nʋգy��3":ۗ/Pp��|�p��a�]�"Ry<�.�����`�w���YߓB����t���t�te�7[��Q�֮�U;�S�j�m�`6�/��ZA�0��ܹ���1��&|�#y��R�V.v�|o{z6��z��*E+���Z(�7�\�����S����E��L2��m�:��­ݱ������a��.ʽ�n<�fJC<��ްsmOXZ.����M�\Ĵ:;n%�)	ܕ.�ts�*c_��=�*X�Qݬ�����w[=����bX��>���c)�2�4���R �P�|��>�}6�f-�=J��ـ��lC6*ï�}f��X�V�,|a�V�M��<Q��U�p�*�&�ܹ��� 
�T(�(�(IQ��������۳T�g�"��o�r�z�zFO�n�*b����N����֫j������
Ɏ�5�71*W���@���	�o!�����Tͮk����ܿ+BfUu�;�k�����p&��U!�>��r9S�E�I{���o�Y��k�2��!�k�pj��o��^ڀy�u\��t��Y;j�O<o��(�竲����܌����ɶ�|�,��`R3��7#��m�1�5�+���n�,��~�v�K���uVP�S��^�h�i��U�,��P��q1S���d_��J��.8����wP=
��S�m��3���e��W���oDa#�l�RƼ�r%vp�޸����'lKl�d��~�#\�>� �����᜾�g��+�Ǟ�f��;Բa��O�������������Y�~jՙp����p�~�8��=�0�t�.o�mb��e�uf#���v�����v��et��w�Жk�nH8��NM�[�R�9V���C\̔�	�N�Wwa��7F�V��.�g>;.�Rْ�sO2����=s��G�n��s�ڗ^��;\�gWGaĕ�=���X�uel��a#sͶ=5e;���� l-�X{�;�_���>)x�,��ޟ\'���N�u��[�Փ�вH��~~׽���V�l$�a��������[� b�D�ܴ+5�v�*���{S�� ~��O��6G�.ZϐF^˄�Dg�E�穳�5���boNevWݡ��z��Z�?O��)�]h$�^��c��?~�k�\q/x�;�X�4j�\��O�hś�Ve٪����x�jۇ��*����Zs�1!pj��-�/y���)�ix�k;{�ɲE�(,f�?}\�k����1�0��ҥy�����l�s1�Z;S�ٰ��?/Ĺ���zFi��r6jB���eVE�`�����w�i��U ��K/���@��*��48ɣ�K�U�v'M1g ����kh�a1���F�_�r���T�<f�<z�_�V���eyCR��P%�9	�Si�t�7���{ٹ�f3՚�v7��ٍd�bC�C�ŝ��g<�SCo�/&U��Sf���7���Qc�+��L�'\-�X컰�8z{���|�ݷ����?C�a��w�X�APԋ����������}KS7y�^Y*�6C�����\Ͷp�
Z}�q��ջ0���T�?�I+j9y�ax�e6{z�B�Y�����X���3J鵓�neö������$����%s�w: ݕ��wrB6V���t�o��*� �ǔ��1���v�f]�W����聋z�Dc�ћ�[�X���k�w"ټ�N�+��P�g4^[_�HC:������8��������ޣ�-|���F���z�<Klw�y��}�$A�70*˜�^��ݐP�h��֚ez���v�*�6j�ި�n�[Km�O��=�T4�;ruOEN�G5�Ì�B�z�ʹӱ��X���4��6m��a����8%��2��M�\k��4��41��mo>���W�s�yB�ѧ�����b���8�82�<�4��/��S7�o���������%��*J�~ZN�)�u��QȤ�!P����������:��)�['X�cH���ܫ���g��������s|2�"�.�x��a;��R��ɇQ�!���X��R�:��t����_�G� �T�����+���k��Lw����$o�\�).����L�s��ō��*����*��~�㺣�m3�R��z��5M5�񉮦��������\�$䊮��D��
�ސ��W+&��L�,�Q����U8/1{�i��Ureu�׾V/_�Y*��%!\\��i�ζ�lb}�c�{[c6���:�&.ɽ+�f԰�f��9	;K�w�g+jw2u��!뷌���S4��9Ю��X�ǎvl�ls*3r�EV�z�>�.W�N���jW=I�_F����oh�1�9���*m��z�e���{:��Q;�l����*��l�ӼI��Օc�5�����^i�n���ؒ������e�0ϭ����Yl��j5��F�{��1o��꘎po{�L�2i�{k�`o6o� ڸ��v��t�t�lg{ ġ%/UjoJJma���j�ϖ5���h�TS���Yuڵf�P7�������Ȣ��N�@���/��Mq��T�V���ѧ(,˝At�
�i��Δ�q�B}��ی�b��� ��	@f���e�P���)[-đ6e��}�  a&M�V'�0ް���^�����\S�����V��ܣ��m���t��QΥv�����;��"�b�=�`��Us�&{긠 �=�ՅK��k+u_�����#^��t*?�q�αT�j���U@Ӳ�wmP����/;��2��Y��E��,g�5�܋F���9���r��zK%G�����BwJ�J���,�V��̎�6[z!K�r�V��-x���&y�e�����2;��Ku��}�?��^܉J|�=����y�lD����3ҽ2�V7�W@
�E�K}s0��͞,Zv�e�8�];3w"��qz�^ejP�F��5Z�Mtu�ޱ덨֤��>��H���m\b�^��_���y3�L�h�|{C�Κ����Ϋb��{_�3Z�y��Σw���j�ws{7�f��c�j{��6��?�B �\�^DŸWGi�x���"�H��}f�����x���w��`Һ�磹p�t���]��-�t��x�V��Cԫ�}��mb^���v��f����S�}��� ��۽��fv2�/Xa>�*�5�]�{z�fn����S�[Z��p -���r�b�����IA�����op�Ux�2j'������3�үI�Rf��`��f`�s��zF���q�:�1�-�3������v�b��uH��;��{fy�zs`S��;�vR��w��فZ��n���7jb����W�◱���C��n]q�7����oGVe.��י�P��<���8�uQ~�v����AK�\?m�d'�Q�nTWUl�KO����z�˖6C�.s���[�����OAM�6Ku����̞��N�k���0%��#����|�c���lh�p��o�;�� O%��gH����<n����g��}L�{~�B��¦�9�2Ǡ��{j�;p��*o�M�t��h��1��{p3�t�B�J��C)Xs�hX�뢮�W1�{�g�y���iXx���Ǥ[�+��!q��]\㽺��8iu�Xy�������5�6��A;tn'��Y��4��Ѯ&�f*t ���4տ�J�U|���CgQo�m
3�7�\l�wg�*�'��-��{L9o��
�[�Wf4]�U:o�[��S.21�u\Ǘ�`_��^���G�%���xtt�who�m3��Ǜ�s�`��ב�Q`Q�1�E���ʷs��1S���|��^^�s�������\��gُ+�}�[]�/����ڨ�v�w-��[4#�g�~�(�^s��\�Ԓ�V�9έӴD�e�.�+��ul��+z�y7�u�P%M@��&�D���0F%�Jw����,���̽�f�0*���T�앺��S�x�Q�6�&2Q�����{�3{Z7����Cv�	��_�l�p�T�s%�T��wC�]�k�tԾ�A��c ��pl��ѵ���ӵ���`�6q��km����={��*(��Ca=+����rb"$'=M\�uw�=X�ۛ�����<�z�]{����{Eㆰ�4�Y��<�7(���a�k�����t ����ټ��K�`ug�:��o�ֽ=��P&�0N#Y!��z�,����J�:x9�DAu���Ve��Mz��\P�fW�cEa�[&=[�'�������}���*(��˓�h)���=�S0f�;�v�p�XȺצ�N�LT�Z���u��^���������LV�;�K�nle/���x�#���e��,��HP6�p�����$���ݢ�+{M[�� �|���v���z�7A� ��7�2��ؾ�_sV\�K�v�}(��ߠ�/�_�v0t��{T=Y����u��FFo��:��i�T/ױv[wXgmi��70���nt�����P*��ݰ�����g�h���~5ST�Nmn�qaSCg2V�����j���o���Kl�|Z�^��'��݀���זjd�pS���voD�p�#%���C9-�����ͽ)fq�g��������-܁���wts3��<��y�~n��tOdw�XW9	+U^�5~���f��ٮ���}�/ٳ�ǲ�+xZy�j�J��m����R]+�[�dj�6��F5�@fhwS9��9e��4��f��̱��BqXֻ c>�W��CuCWB1P訮}��'!��q�۲ժ\M?'B�\�*�4%������Z]@pͩB�V*���.tt"ʻC�-�Y�z������gt���<��o���v6M��H�+�%�m=�����l���8�����{������vPy:�����/��+�'l k�`f�^,z0�wF�ޔ��B��;��I���v��u.��2&ޭ�+�G[�JOo��}z�N&����{s2J�&�;y3��
�)ma��XQnY�����fZ[��kStKmdLt���kk>N�jZ+#�c+T�@��b�q�N����9՞�d�:a��j��K�Y���
�!f�[Ԯ��8�v�M�9h�*�&�R^�%�r���n4x������ҭV�K�(�]�����w�.�V^�Z.��bRt�uN�j�u��R`꼾��Y6+XD����7VjD�;���ܲP�^��-l;3+��ܶy�ݡpG�A��i�0�-t�X^C��_H���姻>�!���a̗ӥԲWf]t��#��k��f�AD%���K�x�|��bh,������q͵��F��&�Wvtm�<a+8P�xR�Y����_��'a�aS���v�D+����Z���5��-����-���
�f��0�ܷ�ٛMwP^�,l�ڢ�{�>��fDb���@T�%��mh�n�� �kA=�&�8��������]���K4&9�h@���i�nDF��[X�(yr��!B��m�6���)�l}^��'�����R��t��j��^�"�B�@,����㩩�f�K_^B(fTk<����]ں��@�W�Q�
�n�l;+�FOe�'2��	a�w�x#쑺X������"���n��-�������P�V�pf�@�Z����sj��Bsy�M��M i��)����b��嗜���q�| {�u�&�(9�2��V5iW׳�kI���^f��ޠi�g�w!2E��y$zl* YY�ks��E<}��r�ak�tn�����k�ĩ�����&��9�/��1i�r�5��}xq&/j�9F�u����Th쵽��ؕ�q)X]�T+��j��myxdmG���Z�2|-��T':<�^�G��e:�^ �3�N}�U� R���JɝQ�,�����6�ʃ�0��'�::��ΐ���*,+.���� �J��u�����BA�H�cӆU��7d��^iU���#ї�:��b�,3b�Ѽ��+/�z��F�@ﲃ�Sf�  �ߘ}�oi2�z�a���Õ	����H�FVۺ�{�FK�],��P$k�3�y
5�;��cHlI�#�e�ދ���)�d�����yJR����k�1��
|��زE�Ħ��g�QYo9fn"��7��r�n)��׷�b��];���Ե<wg;D�����ua�[QB*�!J����ڬ�lO7W)�������xg/�N���D�U"H�b�1G��\�5�6�$ZF6��;�ݦ�o�[����.�Cǵ�N�������H������6�
C8[���ꦲ����.:���ی���}{zzzz��s�g�9�>�K����'u+3	3��.���D��'�	�G(#��Yώ�8�oo��������������>~��r�EѕP���]�CPUږ���ec�8�W��g�����������}g�c��&&4LP�29�m�#^Zf�~���زBD��.#�A�F��f�.o��\���"ȷ�/�,.�����%�O"s��I�1�]e���� ��RW%۩�;����wo8�^hs�X��v��Blo4�˕\���&�2�s�lH���*�8����NK`�:k9��	��O[�#{wu�'�|��,,�ŪeS�Q��Q��cf��痒�wt�a�|�qP�O�:��x��	�t�"WX|�4^MU�sG5(��b�L~n���gl�m93��8&I#�S"ϑb�2s��۳�Z�$���om�Y�y���w��w'�~.�U�(Fȕ�tmYq%y@U����ܝ��I9��6(�--�5oU�&�Aѭ�%�G�}� �� �ѡ�r�G{i;��j�M��v���^ �<\G�0����F٘�m����7��[���,�Vݱ�s�e���=� ]�)5�N;w���7��Z�)/mw&��PW݃^�r�����3�s�̏;f�Ε��u��_�u�����m ����_N�D6^@�Iԥ���v��/ns����ŭXx��̘؝��T�������v}iNU�l�G����t�H���Lھ���r��m��7��*�<�]�]k�F�L	ܶ|��ꇢE���9{�q�$��Oz؋o�k\�Wm/Z��7�oy�br"y ����oV�l�����H"I&^��|i�E�V����CG4%
�C�]2��u�6'�mU�]x;��	N{��+�����oY�.bƪ�+�i6"��#�f�η�˼<�{8�\�תƤ:�V����,�h�Z�0CAܩ��۶�]�-I����<T�ʰ��c��V!h��,�Q���F�K�m�k}�3�n*��υ�� t6�{��;N{�\uy�>�]���V
J��iߢ�Z<�{�ұ����f���(팲��G,�W;!����ޮ���Ժ��{.��챕LT��ulo$����&���aO�^�8<X� xx~-�<�e2w~\�p{fR��F���T�Ŵ��ss*���'K?k�`%c��y}��Ӿ�3Z=�� ��UR��eZ�El4��Lrk�6��g�d�ew����U̷*ht�0�@�q~������y����ë���!��{���ڜޮ�ֽY*�@�V��̘5{�p���4B}�Y8���d�08����� �]"[�Jn�%��j��i��6��h���1BI�WX.�zMŵJ��Ӽ\N���k�x�]~��]!�>f��0�π9jj�UX�n��]���o��tt.V�sj#ӹ��ߒ��r�n�YM���^�z��MS9h^�,)��JB��tc�tG�_\��%s���Ŝ���1ug\]���}�g�5��"W6��G�Ψ�eי�.���Uq���˳[`?k���Հ���y�i(�|"�귅*^���+��.r�6{������u��W!)fu�V�)[��ӫti�����!�Q^�LdrֹT.���P�YHB��й�y[Aw`�2�3�{&u^U�o5#j��.`܁���˾�[6*��(Je�/xh�j�p ��9���R�g��eG�+�27��u�+�ς��T�m�ǽ���G�NƦ�3�J��͙j}�s�}��W<�qy��5��}�tlk)u!9ğo!�V���Ny����Q�נ��Zј{���x��@�ͺ����A(S��9~�ӄN�WNI�l��7��\ݚ�%b&���Uc��§����j���z<xlmMF=v�=�X&�˭F�7��a��6�n� �]�C�K)K.���֢.1��R��$������ꑹjf�[4��.il �r�ɩ�p4�|�'"��gd�]	PW[�$��i�M�*��[dXڷ��Q$9|k�m�c���-��V��1���PKki�T[�юW<�]n�&���;{�R��geh�:��샏�}�0�-K7���ȖP��G�Y�����;:��cs��h����
�!]����6;{}�ұ��j����fn��F�l�ƣ�VA[O/$D�n ˈ���TƄM�@z`�~���Ϭ�����V�q,H}�Y���`�[it�k��[�g0��7F��
֤�]���
ͰZʾ��*oE~������=��tV�Y��7�G���o;�����������E�ƌ=/UU�����$��'��YS��*����-��o��ܠ��xř�5���`bcԅ��Pq���b�I�&1|;���X`sK���s�r��v����m͜yG��\��Z����k� \���M�5���m�������̉2����}��ҿTs�ʠ�Z��Of�vO����z��^�:�_$�~���g���1��U��t\G��B���e]��;��F���%]����q݃v.w��|��ki�c����j*_Hdf@~Y��9BX��T?wFz߻/t[�V���H��)�`������t��bk�m�a��2�{*;'�k����{U��p��4���/�c�]H�9P��k�Mo(�|��%�&_r�}�nb��[8�f��U�d�T\��z�֋�K��i���㘿!O6��L\���%���-���mN��.+�1�B����m��o�HH��B�noe_r�����VW�f�ԛe��}���:u+o�B���8��V`�4oX(�$�C�5m���k�tNc��76-�N�� �xj�s�oj�a�h��ݛ;9qIq,5L��H��4���%��:��441T���{���8w����_�pw�/�ws�r;+�uS�޵��@�L���蚳wU};���ӕ4�>�q*�����[��j��Ɂ�g6��\��Qq	��U�D�a�\ȑ^����0���j_9�"3+`s��D�}�����������ڵ�K$��<��W5���c7a��(8���4�͛WZ�5��o�vFώ�ZKsBJ��5�֝���4k9]����������l����z�9�z��ڬ�q��[<5�9�_O5���2 �gP��|��G4A
�"�:��U�RZpzѼWώ�饄�)ia��7�u�cG��w@l�j���_E(ûOn�x��]�>���}}k����ۃ�Hj������or��z=P���<oUN�V6��3��.w~�i������}~�=��t8W�]~�x�{���m5M���Q�g���f�.�B���O�m!8��]m���M-��/v��зz�_7�O$pNV����ݎ��Y�H�]S['���u�-�<b�C͙�����it���;�KQx�w%�n�%�r���7���:z9�7G���'�̧`>�W�aI�
��hڝ�,xuc��bh��+�7���B���ڀ�b��f"�
�&0���Y�5sPw��{��\�E�f���*7J�	S����j�Y�2V���z��;��x��~���(�����w��R��c�)�`z�_�tΕ�M��6��3wA����ވ,D��·�S\7��S��	!���Tr��1*��=Y,ψ���2u�W�J��/]Y�S%�˘�����k6�I7����Q�y�-NJT̎T�4VA���]���Y���RE9�εwf�pʈԽ`z��O��Ok($�e\��Y1���&<i��^e��B�T�U�lWx�8+:�M����E����[d'��o�C/G�~�p��[㺙��qS���G��(�O:��������7����:F~�5�b�_�j#t)"Z���|!�̧�s�ᑝ��Nu�C�*�h)�1:�׹+7g[)ݨp���Zz^�0X�R���{_3�3�u���']���B�����8np�ױ��Y�=#�P��Z0�g8���\]a���wh�k��Ln�����>�z��;
vi��0n�+[�z�JQ�si�ĳ;��>���/OVU����W�}�"}��8'�� :̀�H�7�K+'���n�jh�?��w۩{�x~G��z^5���yt�]"�
�Q��W{ygfZ�8v��͵r=׭���t��� �Zq�|b3�1�qޱ�v����1�Cy�߇�^����s}ս�x����hm��.����[5�c������D�O��4�NTh�Q���^N��r��M�,���=\��3[U�Y��'m�c�\4?R����ŷ�M��x���h?C�l��fb-stD��ݗ齏&{��k
Yw�٩��1�������j����58�y/NP޶/�[��!2��ǚ�����6#�uT�NeTV�j�Wg%�N�{{�D�,�Qܯ�~�?Y*��T��gÕs��<�F4�<��������홡���>�&�Hop�o��(<�Vl���)V�,+s;�C��=��ʢI�N�h`}��/���ԓ!�|f��ζs2BR7'i�9j������4r�Y�ښ�T'Df;���q�N�^ ~ �U�������������-�uq䦀����^�n�Q0�N�=4�j����:�5���o�U����_r]����SZ�\�!L	��jb(3�N�}�t0�lI'
���c\����i��/�[�q�9г+;��u��K��E�c*�Z��{n�~��9�]�o�m�V+�ޥ~͝�mS7���|��h�y~���/b1�]�&�ّ��&a���}�O޼�y���A�bgeSn�O}��I�t!�݀�n;I�W���7-�������۽e��J��y�Y��UeGve$�Y���ڬ���j��u�={9���ى���a�\5b�_r��v�޽���q���#��D�?\�8/pC!ڛ��/�[`�w��i�O`�D	J@{jk��ѝ�z�37��ns��Gg�P���F��q��q�yRs���"M@zU~�kYo�@��ͻ�j��v��޺)�Ќ9M���n6.�����������Uң����n�Jl�Ž6×�6+�[4��"�3 t��A��8�7>��Y:�,0FWm0��f���|���;Nd���Bcƣw�2cr	�sKw�s�W��p�wK�K�*MÝġF�*A�j3�0gvf,���0$y׉�C-��O����H ���4}c]m�ݾwKH��SB���\0P\��l6�j�|9�s/��E�e�؉��ku�+x�WY����O���B#��O�ީY� o!�;�8%�t2��}��{���\�dDL��7z�Y�Կls=[�('�GԽ��e3���;�Rk�mWo^뼴�K���=��q��~i�N���P�Ϊ}�t�mm*��ê̶*�.J���ޛvf�n��4{�%�}X��5ҹ�B��Q��UMc�GL�w��ܞޚR;i�=VTA>���[�[��&�F���踀ҷng �ms^�c��Im-�Q��j���C�2�~NЮ'��'��: �	O�+s`͇&孼�7^p�*������y�����^�u}� i�m.��L�8kk�}�[��B�pw}|��+�����9>���PV�ZB����k�_7�^nwr�b��=�d{ڊ݊��ht��0I�H���@Q�A�3��q�����
5�%�ׂD%�m	 �ز�m�ԕo~�-�v;^܍��N@bװֈ�\<�%��ي���כOuAx{��7�7V��k��Й�۹�����8�*6}��@K3���Qz�h�7����Q�Q��`�Glи���x9ώ�g�fԬD`��e>�{��4�j<7KUBUg;��4��a�8�`���K=1��p�C��`H1�Q�CLF��d$4uSꔕ��d|P`6��Q�a�ty¾�EI2�g���z�����8�S}m�����8�\t��\�[�?g򮋻���Qfv������E\R�������,��ϬF*��,��v{/:F�<�-�2rjj�38�]����cs�����@Qj��HM�p�1q�,����A�9��u�Y��T3{��((�X�U3�GV=h�W�2Gs�[ec�Tb;5r�.��`6쳥�l���<����_<�$�*��"�MZL��E�u���؅[�<';�eP�����NT�-�Z�R� ���ẙ�t��tD��"KȔL���ܱX��u�@���>ͭ{���sz�[·��\��k/RYst��9t�Oo+��23p���_u��N�;C�Z�Rk=Su��S�m�i������I�(p�Hr�����钁�r��x�����!�J��X��/R:�wt�˨���eWk �JnR4q0k�/(�s�v�8k��wՕ��;�	�ҭ@�'o3��t���+���Ow{xY7��n��]R�w�;���V˳�͋ڽ~V3՞~�p+��	G�/�ԵOM7ln��.S�Hi>ݮ��R6��[�p��r�8(U��䰇X��u�կy��рV�]-����\"��6ˎ�*�W��쭼|����JyM֮pbvs�����+6ڄ�+O��Ύ�oLc_4�(����vpv�s/���MSΞ#"}?��*�����;Va�ǵ�u���D�Z�79��XbTY�1N�i�&^.��R6�ʎεF�NjS5����(f����d?7c�uմ:�V*�u(�m�!��tM���J����S=��f��2w�=y�|�V�;��M�`sju�]a����� �^��>���uw�����dP�s*��$��)��&��:�*	;��_n��-����BV����C8eҮ��0j�p��<��4"t��Ty�Nsi�P#צ�z�){���5Mb�gD��4�K���F����ʈ���@htVwr���
<ı�V��yr�Q
���m�S��ZvRQ�s2���t�A�n�љ��%kYA�kۧ�-�y8ݹ;�\�8��� ��r�0�"�p����� �Bv��s�!SO˲�v8cM{�8Zv���$����.˘o���mخn������5j��z����+q�Z8RBT�RSU�&x�ͫ���sEImf��#���h������J�Q���6��- jW6����}*b�����ؚif<r��n�FQ�d�G�|Z<F4�W�%9ރ���|��;��݄4�gW#��i�R����$G��t���ӱ��K��j����&r���� *�c `��²�5�I��L������8�-�����E��ǩmNqꎄ2C���t;���8�s���\�.�A&�i�k7Ю���d#�wIc�Uѿ44�U�n�r��V��v�|���M=�X*HI4��X>o��M�dZ�婼.�F4�CkB�Kq��i��O4����0�Z� K:X��c� uvZB���[f9܇����vE��P|ެ@�C�V<ʺ�%r���65��.E�-�����VXt��ٴ�0��WX�v�q��zx^R�Tum##97zpT�^��uS�@,e톅=��V�ͩ�\�m�}$9�u¥t�������5�HcI�e�.����>ŒC߬�^��q5�e��GȒ���wwV�������d���Oߎ���==>�Y���Ϲ�?Y�uuj��H���ֹ�n��;�MͲ��Q�3[g��.G]s+�p�|Ϯ�8�����{{zzzg�qϹ�gӿM�Y�a���*wk��n�����$��b-y������G[�����������~���==?]f}~��7s�,�jM�u]��L�s����*��3�J+Fgw��q<����/�5)�D����t��d�3��ES��Q� ��IPy�tR�ؗS!�	ԇ�m1(0ˈ������jyBS���9"�2ͱ:�ڟ۹��yI�.� �X��
���VIS�(;d�5��*)3�?6_<�9�Ge�n��8P͕�G�U�Re<�ՙPje* �F�duˮ*��.�v�Y����w4ք�4�ԕ��r��/wRM������rSL�bK8H)���*����ࢩ7����*�⃍D�9�n�$�6ș�[Fa�V.���-XU�L��Ɣc746D���|8'&곪�[�����M��4���p�
,�n�}�/'Y閚�ܾܬ���;"1)�T�4Q�<��#�nˬ]7�^�ee@�ݮ�i��v�]������tB��3�+��d����vd
���SA�^M��,�mO�DRA�u�ha;^.ܯ��ڻ|z����7�ca:�Ѽ�
:���F��s^��Ӱ�5@Q�[��5��
�é%Z������Jj�9yj�Ec�O�8'��蠆�7e� \��{�?j�y�Y�t���!@���s���H�u��\�^�e��Psך�.�w�����}~�g�e�[h�h3<:���1B�Z� �̩��^�=x����!�5r���Cl�97�����w�����F��U��?e������o�9�4�'����GC��ӣ'��'nW*��W�{g�o_t����� h����ǘdhY殸��|i�a� �<�D��+�^ud�}�_�8�9�]l��L�!�,��u���/�~��/Jv���1���o0�
��=	����<����k���v�d#��Say��S;��ug:�t3{:m�+M��f�s�-)ٻ���.��N��
:j�F��'���	�����n��5)�?s����gu\�Z��^e�^����P:M(N�&�f�v��q[ư�V���^�3s�SS�ښ��r�&���9�3SDȵ���/C�v��ۦ�O�=�[L\R�Ƹ���)5��|�N��7bT]��h�K��u��uLl�RmK5�M��|\f~��է��~�x�E=EG�6ͥۢ�u�_)����S��d����z�z��Wx�^�RSAӑƳEJ��N={g��]rX�ߤ��¯|�͋%�k�V����6{
�8Բ�d
�Ӽ^-vK1�TgB�� �So�O>�v��z�7LCV�K�S܃�C�m�m��	�7�cDJ痪�Vҫ|�%���R��=�w�sG��z	��̘�["߇7\ɷ�"��32��T��5���r�X�3�-�X	{`�B��c"N��jz�q5��f7%x�gq�U{�?V=�;Z
�o_��L0�t�ct(Ԙ_�n*���z���H��y�����ű�#�I����#Ro7��\����z�JV�ܸ��9���I�/�ْ��7���:rY�==\�dY2�*i���Z��21��H���'M�b����G� 34�gRd'I�Y��ث�>N)dFv�OYQݘ��.����M������aN?	���]�E�u�Aߺ�"#�5���Y}���Q���7���p�͡�\�:��y[O�~�2 a�p��"Ww{w}Ԕu��-��eݙ�m��p�SF�S��|!5���y�mn�·�B��`9̫y��P��SXܳҬ��=c6z����c}����r������Ш�b{�X����)��qѩU�?��}NoN�/�QކV5�O���"�Yr�zg��늘���������������Pژ!x;���c��d��'��K�J۝�Դ����L®U<׳yd�ꋕ��JY�:k)��������=���6��Qn���&�v
馸���\RtM��<s��oU�ʨ�筌l�MNFcu>�����n���3.T�6*�J!Jνk��J�[�+��C���4cgw�>=^��D�ʂՎ޸iC�uZ�:���������A��|�JQ2�|�9��N�^�4ki�n����F7K��ǹ�Gbz{:ct���ݔթB�X��ET)�@�Bcnm���arl\�F������.&ͮT�q�������^*�#|�A�7�^h�e�9�ܟ�j���GR�r	�z�{�Rm�S�M�ݚxީ/��Э�ݕ�y����["��Q��yb9��1�l����Tل�����m�>�5wf����J�ݽ��S�>�yl��5���j
��k���U��Ӟ�����L��qP��.�Y�cU�!�3-�m��xW���Ԅ�U�Yq��`�Ռ�;�۝R�Z5�<�o3bN���b/��1�p�ѽ�I��r�����˔֭vqy����l�u���=�{n�+ۆΛt�*e���r�w*j���S�m�{�:Co{(`b��c�k�+맀�Sݹ�&2�o6����g����zY'=��t������3}�`�ze�&J��7ꚿ��_)���m�_|���Mb����>���-C��� ܆j˱�xѿ���!'�Z����"�������)�+�v*�+0�(���ZN΍otxW�2�H�Y�K[�=I���d�l�Oe��w��uC<��]�\�w�X�)vA�Z�Ʃ�Τc��Z����9/�߱m����eڥ�I�٭Y���MiI.�Q`o�f��+]��*��y�ټ����`��M1�t]㎘���M+{�vͽ�ō�2�֨EL	�B�����R��\�8,\���z�I����N�e)3�O���Rʔ�C��Z�F�k]6�Ik�:�rY:ޠM��K5	Etx��μB��y�я�㓃�ݵ]yfXLX���<C��OvWw��{�NHJ�gܩ����~2�CfGl�9e"lp͚[���.�gf�d�	-ٮ>���+'U^mW�������B��ng�'rt
��3ɴ,���Z����Z9�^��m^	S���92{5l���OM���x"@��m�����8��u��;�d�E�ɞ�n�!�jcw��̎x����l:ފ|q��Y�d����9m�j�x�·�g�}/[�}ݴ5Ӆf.2��Y�͏7.��KE�ƒ�7Բ�
��֚Y~Kq'`�����#GL�N��ig}���'�V�v��\8Eq�_RV�`��_(�1�fR��������9�����v�]�.�ʘ��s����Bh�8���y���	jyR��i�$!���9Upz%�����o��Y���~��9�G�!�7�Ǿ�5�7҅p/����+��Kk��_N��H�ξ�k���s���vj�ΏW������J�b����m�  X
��n]�OJ��~gzk�nt�nv7GX��gZmHu�D=E���C3��%�e3���8��Y��/�Wf��vw_�I�W��¡KM�h�k�e.�����pWNj�Μ��js/)GI?������x����u75�_��KtGT�F@ӵ$ <N��G�{�DEgd�ڻ��}	�k0���N����b�R�5�t��CWL&������������	�6��]�O�哽Qs��S>�L��l`fkz�=a�5n���;p�Y�����q��N�������>WW	M/UZ���*�f�o UŤ�e��/���5e��.+���1Һ�wR����:3���,5BY�RÌ�g�s�8\Uz5�Z�\y�>�����l��s�;����Nr����X��=��[Q���eTGan22��u�RV�Gܜ�Hb�oUf�:I�gq-m�R?Ǫ��N�JI�'��kSp��&uw
6�Vcpȹ�V�i��i*-!��C;A�x��K��E�W�?w]�	���7�v�q��G�;o�#�ϫ|����d"+�f��gFY����#���_Z.��5-����Oq�G[A7��ڝv�[t�=Z@r��ЮB�����ֳ�FG�����,ۢ�� 4oY;���GYg�ns��n�x�=�r���ɷVC�;׀�*�܊w4GF[3EZ�������\�K�V��*=ۗ�,Ip�3��NCS;�aN�v���l��>��F��vW����v{�����ζn#FTMf��g��Vd�:wĽ|�WҀelz�_���W���'�ԩ�Ȫnl��zj�(?0�p�(�[��W����@u
���WW׌_B�r5�{/4K݂�
5y4�xv劥�����Ʋ��%'wY�\��1����n)�NU냡�aW{��ү���B�F9G����_��	���: ،�
��6�BqNN��NE4�g�MJ-��ޛ,=x���^�!ښ
��K|�ŉ�1��ƽ�{��IA�s2�c�<��c� <~ $A3�U��j{�`��t��A�>vR/����n���-�@���>�VīN�C�u��IC�v���������u��$� <>+�7�\��#笪�Q�2bm.����4��t���o�A�8�ë��Ws7Ax}�P�b��u������nls���T\����v6��i����-{��ݰmCK��<��UEP��Q�ʛsXp�K���,z��K��f$�u1�3P��3<��e�;5���
�=���Lpw\+k{���4��h��oW�4�r�x�*E��,�z: ����ϋ(ੈ[��Y��P�4o*�{���ޘ�g���yOF���_;kw�En�]٘"8rU�k4�n���%��*d�;X�m��Y!�=�O*�Ӻ�S�c���2����͉���30�r���5�%SDd+혖h�3�Ɉ���C�/6X���w��Fl�|�ί'��N�^���.���iʸ�̬�m�ja��FQ	��6���*�A�^[VƞDa�y�����1���Q���������n��@eН��97�}΄}���o�gtwx�4�xm{�I=OP��.}���Wz�ɜ��Uʊ�}�ݠ�qA�=t��ꀹW|��V8"fj;L����q;��r2}�,�	�
� �R�w��T��4���y�}�7Q��ym�4�䡜��wF϶+����fvkDt�R˺�ݕ�s��\�;�)��ֵ�9�:C�#1\���R�j���玷���zv�y�wK���7������lM+�z�!��i�e��b��-��o�Kr�o#��O@�Y�Tb�e70ݗ����gC��l�[R����͙�<T��Tg³�=�
�ҭZ�|���N����+�4�ݖ��k�eKV��&q�[���ζnL��' ��gq}�ˢ0_{��/)�oS3{�Muy���<���UH���d	���a�Y7���g_������r��J��3V"�S���^!���4hȹ�����וc�>��g+�=���Z��53uə������K��gTm�=���'�,��ވ��]�㮒KV�\[�ʹ��_��M�&�:"*,ܰ�p��F�0�T���� �M�:�K��;�b+7�/I���v���U;����1���6��rӭ�03�_k��
5b���K�7��Hl�������98�pB���o�)��L]���ڰ��-�����=��+��u���<�d��:'��N�۷�k����Sl��=V�}�S�$�����t�<���S+�>�8���S��V�,^j.�#3jt٠M�}���3��5aۋ8��S��vX�z���ĥ<��/'���j�'��5��wFw��Ѯ�]y��n�"Õ{��na�v�"q��������ݳ�/uV�\:n�7R���"�*}}��2���R����!þ�}U�{g���|�}��u������﯋��P�L�D�L��Q��-���/m�Io��:`nt�a<�#6�>����1Y-je�+6����{k���my�N$M{Z��l�ݛinhUL0[��H�gw��m^>��c��s1��Z�]�ey�l�s)�O^"��p�i|\;�Tf��'�����H֚��z�,�ʽv����Q U�X� �����"�P���G�<A1{,μ���HB he�$R�!	D�%�I	�)T�	��I	�beRdeUa���!�&0+��"�P��*J��
�"B��� �!BE �%BA �%B @�!u��"�B(!"�B(!
�B�!(�B�!�B�8�qD�@!	�@!�@!D�@!	D�@30�@B �! BT � PB �%B �%B �* B��	B�!��2�@$4�B�B�fB	H�!"��B� �	!"40�� �HBQ!D�$R�HB!�!��P���Hh��CHB aD�P�%B��Q!	P�$B�H��|��A����"�� �����D@S�^��)��4�wl��=�N�0��Q#$�]5��fF���*�>9�U^��*� tAy � y'��Ԇ`��ۜ4�ɮ��%xn�����[X���$DKc$QP		��	dBR(@��	X@��RT$�I!eA!I�!P��	!�H �I$�e`B  BD ��H�$YP�$BD%�HX�$��J! R%�	a%B`HD�f �
&
A�ZU
��TZ��J���F�JE!P�D)�	�R��%B%P� ��P�"D!�HaH@�A%� @���	�I$BH@��B`BD $�0p�?����O�UTh�@hR�@o��~�����~��\B�.��wʤDV�� �n��b]�4���:0gҕ�t� 
��oN�-x����*�@x���z� E��x
 ������OC��_08�����~�X� 
���<vts" 
�b$@ݣ �
�0/O-��C!DVͩ��@uXa4*��qH1$&rs�T�;��.�-$��h���ą�]i$��Ԁ�<跿��W�U_��8��*������L���$2O��
�2���p3�f� ���9�>�����TQ	
�
��!R�� ��E"T�PPB�!D@QP���	H��R�B��I)T�$JP�"��(�!TI B��l�IT �`
�!BP�(��U���R�*��"��*�j��:�	u�V�TB��%EZ��u$��(�)	*UP��$TT;2�ʊ��P���"������A$IPT
��R�j�R�D*UJ��5�LJ+ٮ��  ]][xtnu���7w`�a��KwZSkmbf�u��FΡwj]�e�':QWgvX)l.��]ԩۘ����kEʳ�:n뻻�hWv�UN̴�撒%%EUkI�  6�
(P�B�� �QB�
([�{áB�
��
�����׶vt�s-ݭrWWwsZ�NZ�[vQ��t���:�Էp)u�8�T�V꫹e�֝�v���YR$� �"$]�   ��� v�	��wY�΄��;�v��:Y��v�[u�].Mwmm�fV����+wk�뫶ڻ��n�]��a�m�r]]��ݚ�We۫��r�k����v�*�IP�U"���
x   ���]�W;Z�J�ݦ�V�wjڦms�q��Mmn�Mu"���]n��ڔgpSWHV��\:��+\��,�8�ʍb��-2��RI"�W])<  	���-��w+�0��U�s�ڋ]kV�6J��[��u��m4���;mSm�]ZUh�s��hCS�X.�T�h�vjݷSWjD�5$�R��%���  �Uz�n�����wZ����,��lзl�ù��s�S9A����v�V�s�����֭������&�Zu���Y��n�����$�UT�*6�TN�K�  ;��UPM鳹�� �� �Հ4MU�  [�� S4�4�� $�K    ��J�tEB�B"��  �� UjP��� #=� ��h �S (e� c)� �t� �@ 6��T��R�*QWY�  G� �J�  6�`  f�4 ��p���9�  Ɩ  �`  �� �$]��( 2���*.�a"
�  ��  k5` (� �;u� ,� � ��p PR �  �Y�M(�   �~@e)J� )�IIR&  4"����h �)� ��C@  jmU5 	��CA&�!2��h 43Rֺ�(\f�ؖ�gu%g&a% �NP�2�����=4��N�b��sp#� $�f{�!	'@I$$?�����B�PBD�$�BC�+]��x�s@R�sV+�������vh��kw�T�m
+Z�	�JJm�#RQOT%�8�'T�,��,YԤ��r��=@
sG�2^KA$Ԏa�w7or��4�F���[*���"�b���.��r�!D٥mf�pYQ��V�ۂGf^_ή5�� ���/�*c�<,1/-&av�j,U�t𜩘ԬZmj֡�b��u���'��Z?ll�{�%i�|��K'[Ϡ�tm�$ݣ�*RL*,ũg��/6 �dei�*�][Y`
L(�tNu1�µԫ:M��;Ӯd[���������RN�V �¯ �D��N5>��� ��6�Y{�`����f�732�k�bm�B�3Fc�A�H����4]&U��I\GR��K!�ZV[d�ۧz��� 7V�qZn�$y�c�dˀ���w=��\�S��.��Gne0��z�7/i�����f2C8�ۻmBI��P��2��u�3t�4�׆�q���Da�#�Yw�� e��+J���;�&�-^V�$(G�	��T�Bm�(��a��B��^�H3i��wha�v�k�:���*M(*�H�edbe%��J��GVWz�&�,a�XLd��r�Y�%��@��5�����p�fiE|cɓV�ڀ\t��(ei�eP�VSd��E�K�փ�M[�50��{y�0\$ŠPx�����wu�Ȯ��b&�cx�;P�[�e[�͡2	�.*�-�h��+�s+��ڗ|)wn�L-4oZ(@7�r�iǖ��T�ovj���@�p��ܧ�ښ�+�a^�N�S���Y���Ah��Tp��HIZ�kpڼ��+#H�ݬ�P�m tl��e�.=��4@K"����&^��XSZ��R�i*mnc�0ABJȤ���v]^f��m�m^oX�0]HU��2@���v^�[�j��V���P�����)j��n�O�a5 �o*�L���$3���*���o(MkJ��U�����4� m)hr��<�T��Z1�BV��z�9N�CA�-cp;*鈆�O4��Lyf��0�Ԭ&�;M*��������ܔ�CE]
�/\߬�w��g(�)T{Wa��'Y# j���ٸ��5�+H%�%��+���?	R��F+*K�%�u4�ݷ��o ��woYV&�ZI�2�R���4!�AŹ��V0�9qk��3k]?����Mb˲i߬i�
� M�^KykR[�3Pdr�M"�րE�3�oP.���L@�d=.���Kn(�WOw7"��X�L�*�AZU��Vj=�2����D1���p�2���+FQ4DfT�P�[��G@���řrS!q��2왁n���M�]F=��I���A��fel&��Vw�E� �JQCB�$��ʘPH[� wmY�q�z*P����%]ѱK���",�y����eYȮ��j�ģ�VbWv����i��m�v��
�%�z�㡹X��X]cc]˦�0�� v������r�j���QL���� �jVe��@3z/VJa�����j���k�����m��bjP�[*��e5��x.�Š��^e9wgh�`h� �(�.�]���Xqm�CW�� �5l�dģ�ݼ�X;uaa�է�w�`�r�:LdR��<���0c_ۻ��g^��B%�,V ʦ�YH��ii:���7�l�h�]ţQ�Xl��k.	��LW{����QiW+u,�J}w�-Q��ÊQ���[!�Gb+&��t��cv���k� օ�@hYO]��`�F�QL�A�tkeۀ���Zz/u�[����+OE㣥սlTl'�oi�J�Im۸7!���PLi2����L.M�)O]�e�I]
i�Ԗ\25gtݜc2�b&��HˤdT^@�*P����e�5[ʐ�6r�Q��Vu��`^[���u�K-k
'��� M'�x�P�ۙ0�3��Pc�nbBZ��щ�ˢe$�h�X���y�L�n�yon0�M�T�x�-J�����bB�m�{�]�5���V⿳*#
Ð��F�yx��&椳f�Jsnlz�f���:�,wz͒��ok&Xїx&T1�-M$I�I4�Kku���А��feݵGsY�LX�.���̤�h[�m����1f�AF6�f���8��v��m+��ZuԤ,:�m�ۼ��n���۷���0m�M,d���y�V^˛)*"��t>� ziD"9���;�V(5C6H��;�AU�9Se��+١LёELxU�k>�ri�$^TE�nQk.�R�w%0�DȋUϬ�n��b�DL-FI���51n���2��y�6K�%�R�L40F���H���i"�У�vh��kn�MXމ�A��3!���m�Ɔf\��'e�(
�������q��[��$TW&�ktK�y����gP�x��b���N�&�fJY����ð�zop@mJ�\�b�i��,T��
�!��ո���h��PN��n�k��h-�^�I���U�5�����
mm��c�:EGP+,�b�A��u��V����rڅf�iVn�6�Tj a�B)�"X7s��N��jƦI�![U�eZ��d"RV��%�G.�)�2�&�u��qn�������m�(���5qޡ����{RS�N(6��	��. JKt�lV
Vڄ�T�kTu=����nm鵑Xc*�zY�"�[
���n'K]G���G�J�6�ާ��V�m,���Х�5�M���{R��iV�`�����36�ӘԊY��َ����fkw-�w$���� ���ڴ���o�y��8�y5 �{D�:�,�u̸)cM���7�40n�@ؖ�ӄ���cz�����76t��j+�sq͡q�V��
�T�iC֬{�e��Ӵ,ى��XZ������)���8*VY�DXm AT���Q2�1E���S�t�0V8JЊf��),��]���-)³ө`@$.���7U���r�j���k۽i�l�i�W�u��#�G,Q��
�e��3^$�溘�0#i�-����4��ou}*),��j�1	�z3	#qY� ��H�\m,Qc�n����]֕�j���zF�bn��v����h<U(�+�*��1De�"5+۷`��I��l��%��޴���6[�7f�9�m��iÑirX�k�e���Zx��
Z�dn	5df�MZN�)�5r+��g/k37����6��͕�F�h���\O*Ƀm�1�Ë�9�S �H@V�6��C5E�@�gd���V�Ď�*�"�N ����t�P[A%6�<��^V��l��%B)�ѕ��LԴ�����B�D�����5�\�Z�0v��n�@�M���kܺx�u�Zڲvm๩�T�v���¯F�s �˿�F
�j�'un���VU٫�kDc.�d�F��0�6B���JkI�\-l�*�4���0]��x(Sp���k��.�֌�b���f���@Յ��B���-ٽ�)n�ZK����9�Ѫ��J?*�GXp��]���� ��X�����t�1X�J�
h��GN�^D>����iJ��N�w.m")���@�C�:�XU��W"�4X%�sU���Yi�0���ЇҴlUye��!��FD����(e+�P]"e#�Ǹp;
���$flb\aDe=�Z>�\�T��[t���[���)�4��~���)�I&3,4&�>;Y(��n�;�A��qx�>FfGvʠuS�uu��\���{{ڒ��j4�큘��)����tFǉĮ��C!��	f�ِe���ǻ0�o���Z�W����bPєofnn:X^3*%1�M�|�S
�IW-T�����+����zڌ�� D��n)Y��L�GD�A8���8��BL >�wx�KZt���Ɉ�U.Kf�O�eSǸ\"\{F�n(i&��S'!�C���.���T����5���8��u�2�G
�>feG�w+͒�c+j��]�
Pر:��t����n⭹8�8���W����FT���ä臚U`��-m�e�1�S!�XM���%�b ʓA�1��{X�Rܨ��,h�e �7l�*���B$���YR�������L\{wZ/tPq427���ĵ\���{�@Х��9a�w�Z`�ʺx��"B�k����)@��O\���N���M�~b��4�f �k����Z��۸ɩۅ���-U�nXY7C��S�e�Y�D�Q�m������ñ��w�h��']F��n�V��ƠF1�.k{�/i{��m
���U6r�QpHBZ�ld���w&їP�s6���(S�fU�	���s-����;ba�Y���.ѐc�0�N���|���j!��_�h,&�<����oH�v�#�pE/!Te#�R�NM#v� �4��.F��"���ur%���[1V��`�|�h !X��{B��n��֨�2��v�Jͺ�tdq[:�B6�%J�@K, �}���݃iݨ@y>ʋ�YJ�f�z.��u�L�ܛv�$(�&^�	*��������ǚƧ{B%��)�1I�l,E�U��;�N�m�u�O%��$!�(��/F�,���(�)M��*��/ [nn�GY2*ɧ�̦�̊��9�+5%���ޚ7L,U)��Y������l��+�w��r���v�)�J��,�+�i��*�^�P��U�V�) �E+�X�1h
�`��[�L�ǎ�u��ʛ�m'Y�f<���)KmA7`���m��E��!�G�`Fl�4�cY���]��yt��l�L��C"$,xY�QC.&��m}{���㣫�*n��)���xn]��Ut��K0k%`�Wl(�B�g�-+�,�n�$0���c@�hV,m8-�g֨^|��C�����x5�dj/6��MCNvm��õ+����B!E��R[K\ �+f���cb����m;6U8�����ȥ9��&ލ�.���V6�f�Ȳ��W�؄��6�,�&�KT���=���̜>‬�5ΩIQ�ʷB��1j�gTV@Ò��Fn)"���R���h��b
N���8Y�����9MZS��=��n+��J���c�M)�4��4��&�D	�V��<�ZYK�Y�%`ʁcmŢLt��vh��`���-S22)��c.��b�iI�.�(��NXŮ���Rġ򬅃Z �F��:ǷtVm�B�pDU�N��(�.� ]�e���xE������}���x��:�,M��7aʴ W��s�NlmY0��蚹�a�rBsl3Sk"�{:F�3k%^@����[6ho#6�.�h���١d�ƥ\��MU�hKUҒ-_��w[[�
���AeHl݂�T?CKF��^����n��Q�THU��4���0XZb �{@AS/4* �y���gM\�,i��L�<��bSj��uŐ/m��6��4u�#F
{��i���h'�� &ަ����Bh3����5t�"��x��0��E-W�J�\�4�X�i�]\N�e��\���fCJ�i�Z�7�	A����әJ���t��齭
AFj߉���1j�n��d�pD3�sTP]s��.75��K�r^'�6h��d�[ 4SC⤷r�I��j�z�̽��ۭJ�LJ�6k*m�#qI�ptMc�٩��/+n�@F^�Ha +^\���͈�B�/�o&Q���Z�q��8��zQ���WNë�aXtaZ)-A�Ӗ;�%��V1�"ޑL*×L�z�O,&��<�ѯ�D��K����=�Le����u�tP�xF	eņI}���l�M�3�����x�B�Gp�9�X
��Z���{�2�nn�]��7���l�m]����k�������7AA�o1�Se޻*���]!4���W$�0�nX����s@�aV}���h�9���-c�zD�.�l��B.��^�ښ�TU�eIWJ�T��v�5���VK��9�I*�{4jí;� ���`�,ݰ#�x�l-t��f^A5�2��r��!����R�n&�ч���N�Vt�u���tL����R�m����B�t���6L�+]���`��G��H:�Fi���u&X���{ se�,�M"��$���Z�iY����)���-d1j�Bՠ�姹A^"u�ou��E�(;�BC�y6���m��-ѓ���ݠh�Oֈ��m����F�J��Z&lQnh/]D��2��!����soE\rcsB
��B�͙Ku��Q�KYr�h���K2�KkpF\�������-71^Z�
�����&�)�v7��SӚ�n�2��5��Cˑ�	�5[�b�H�³6�U���`�/K��-)1�n�� ����΂����j5�-���;n��ہO�ɏd3]��H��\�kim�i��D@LP���;N�SI�Q䍊��Lϑ�e��I[�*ZW�ժ�U�a���81��d�Xn�7x��d�7�&�e^��^
v�n�VM�.]I-�5�E������p��%��ƆmZ7��7v�Һo
��)4eXU���2^�
�n�z�lZ�M!g,J6��e��@Ь���LD�6��^��le�KN�8iccwkKj�"��y2��R�O��DҐw$���Yĝ�(i����T-8ea��^Ҷ��lm�%ł\Y����2��@��H�ћ�acvytr	��,ӠȈ�Oe�\d�p[Հ��Y����2�c�66�W �)H4�ZL�u��n��Q����<�&�ӹp�%��/_Tz�wV�:Ώ�q�����;���"
RE���f�[�sPt;���K�iv^�Q�9ޓ\>����.y��XGh<���͹�m�3w�ٹ3��E'�!c�����v�sՏ�vK�wky:Y�kW+�c�O=|ޙW�YX�c�a>ײ{[N����k���W|��I�Ҳ�.�f\`�"��T�ug8�<b�`J�S8��QVRܴ��ebޙ9Ǜ�)GV���ܥ���l�b�܄��#�\���^�m�B���,E���6=��ܸc�%���gY4��W����{���Z��}���z�Y]wT+"s��9_��4��--��j�szHfn82A�Lm����>[�]����Iv;j�N�m�t��3[ܮv��=##�H�jI�M�7b���؏\�z���[��ƫ;�)�Ky;lV���l�k���ҾZV��Q��oC޾+��Үs�}��e�|����k����8*-�zr��c��[;��
)���A�Zմ&��4����j����FKY�p=I,��
�������&�:u�6C65E���Pփ���u�iP}�X�3;G&��O��Ld�Kn��bƅ()e���d�㸛��f�C٥�Xӓu|޽�ءJ���ڬ�g�H�}*D��Xqޮ��Ls���+7��.n�0�`��Q�֛##�$��`:�/n�����Mz�(T}�p�v��� G��j1�уjk�P�.V�e��� �-�.&�w��jD�(EJc��f��D�v���4f�b3O�a7�r�=�~w��{w�k不�J��;5c�p���ݭqyv�}L��'`�`�x���_<�e\�"�d=����|n\���л��+��Z0�e
JGX���x-�ƻa�*��F��$�Ȟ��;�W����pL�ʾ��\���m�UW���ky>������%R�\tuiena�����S\����-K7T�����g_�+;}c͋���`_=&��γ,��f��E�Wa{��\�5��W�ʙ��>�'�H��e@]�]�8P������v��U�L��!ZMA3�`=��|�py�i�����O1Jq�d޾谸�vM#!�����Wn���v��B��l*_(�_e��d���	ǟs7RY]�(E�K�e8�fɇ3x�I[n�'�x�]�T��ws[�~]֭�l� Ç���7|n��;�_L+�p�Er˷e��f�f�"�$�d&��kwt�F�1;���$׵���u��J1���o!��9����y�]KQ��p���V����c):\]�"ڏE`��2J�إEc��T��,bsM,���ԅX��f�3���]+Q�ԕ�wzK5���,r�M��*���c��Ʈ���R{֩|�o��/x;�'WCv�9�5ekʔ����YW��0ɍ��.ASb:�]�a=��#�,���;A.K3�q[:E����ef�����CƧ:�yD#Jsݠ��ld���{C�n���ó��՘�����z����Y��%N���bCa��N���%�ڗ9�w�%"-��1"]s݊"y	��N�.�w ����jP}ܛY{�k��j��7���J���钦���?@��ܫHͬ��}lҰ�u��Q��V{6���U坫ls���i;Uuy@��DX��W1�+��^��m9O3:�����^ryN����|���cp,�%ex.��Qu<.�>�wyi*=c���e7�q}zz��fs�M�@��z��Ї�K�ce��h��AܷRC��*�vS��Ɉ���E��ӎ9��^Ǥ�
gS�����!�ge�ZN��:�R_D(�k�:���!QK&�{<�nڼ�4��Ó��X��jb*��H�_r�����Q��lj�\髫�&'�Q�����u�'��ʒ>��w��L`�]�3n\�l��,v��3�S`yJ����w��p"�An�W5��R�U�:�Z�\,.qK��Mjރ6�^�6��N��Rd�ȩ	�Yw�%b��=٭��ս���9��a�v�3)7���	!�:u2���V���hB��\�iԽV�Y�>t�+�PZ딆����3$$
X��l����yî�:yٸ��8�<p�LWr
!��j�}/��B�H����rAL�749��������vyThv ���r�`��Y�↫2�=��f2�oo3*� ��ʭ�֏q��7�ǣ	��2_�@�ݳ\�1A��شٙ�_q_uۤ.vp\���Ե+��)�G���o:5�)pJ8��+�-�Mh�s�X�oU�;tSV�=S�1�r�H�M��	w-��r1h��a�$��*�hכ� D����F�u
��N�4VM�2�sl+9O4�	�T�;��QO]IC{�h:Q����E�DX��N�o��f,A��\@R�����\w�ʀ>�'�L�'m���\�S���j�n��:c���h_8t���Uʂ�qh^���S�ju��բX���|�7:����7�T
Qwm�qQV��u٦�D�w�b�9=WM�!����T��T�� 	�����VS�gN��a�������kǴ��iX��ۦ;(u�|�����EbǬ��%6���׳��׷u��R.'j���bv
ؚ���K{k����d�\4��.��ʒ�*LZk�\�|yӾ��h挫��n>���̾��(v�����ص1�ZK��1WI����*�W:"o�tv&�|(T��h�α��QH��m�[��W��$��.�T�Sk�W��,E�C�ܳ^Xy��:�f=����LgD��Gco�f���Vub� T��t�q�əx.�E�}���g��A���)��6��
�8����NWo��r]zm�z��x�u���{�@gC�N8��z4>쮨�(跻L#z*���V���N���"�x�=<�k��	��STnh��p���F�x�\ر	hũr5TJ�ѠA�5�o�%�����.���z��Y�WrmJ�.��X����4�Uz�ҟ5�*�5Q�];I��Y
��ٽ�і�oQ��դQQF�5��:�!����PJYq�#���P���L����1���[.���Z�DG��Ȳnt�O�Jю@Eu۽���;՚����'b/o쥜	����U�l6\SM��	.5t�j��fn��b��z�_3�j�]:qB�u�������E.JD��'Nܫ��W�y��+cC���PO�V3o��O���u]��V��*�┒*�V����{y`�����ԯ
rح�������qn�J1,	X
���-�Zt������lV8m�]���(8�s�ގ��7!9�S)Г�C�n|r�@���dlE԰��ab4�����]S�ڲ�h޶���Ӄk���tC�V���p����u;j��Z$�{i=�+k�����
�i<�r�����b�ى�A"^�yJ�x�V����\��v�����Sfp�a��y<�©c�1��E!�����ށx��bCe��{��!2\��s(�U�P<�jd+�T�:A��W�����x�i��-ֹ�کN��[h`"�1�w݈h�����ҧ�;�7C�X�j�c��	�Jvu�O,��cqܲT��Xŗ.���1q�-�$����bѱ`Ʋ����'K�����[�//_��E����ORwpÒ+�� ��j�%�9b(C�W��v���K
まT��3�3�^Pa����nӖ�3��Wp#B��5y[�*��@�|����6�+���o�]C;LSlʻVSB�p���!�q�d��.�Vqń� ���썷�S7����ث���i{��3]\ʽ��H|�V��)�j>����ݽ����\~�мw��M��^nu�\�D��}���껜��{�[Q0[��t�ٳpeE�#�������,�^k	n��O;�@�l�`󀫗f����wh�����Ta��p<I�W��+0L�k�]aXy����p�:�+s���>>���6�0�f|��*r��ڃvR`�r���bB�9b�I�v��5��"��B/p�/z\����&�f�������2v�y�*�ES+:] ���kB}X�Mޭ#�k�Vӆg��+�A)x&�z����j#�q�Qc	l���Xf]�:y�#G��V	��Ư;�@�^���.wǃb�ɚAۢ�a����#k�egler��E'��8����W�'s=����q ��-��,�+�R�n�-w�I�Ko�� �r��nS���j��[7�[f�̑;�z�h����2������˫ݑ��շ.�XA��ةł�3`�S5M�ǈb���-�wsu����\�L�0R�<K��ҍ�x�Q��}ʰ����]aTzz�%��B��:�1��7x�wA�&���=z����(}�R�:SQgJ붜�,3�͍��%���vB+_O��hV�ЌJ��20�sQr�#�f���GZ�*�|���v�+��kv�H�``�f�ȡ�mɭ]xsjj��+:U��*�=L'����`��!� ���Y�]ist�L�"R�wf�RӖ;k�;<�iIL�Hۇ3�Q�Y|o�D+��ͷ��a�AzX{9��	�V��Z�;�#�%�[#P�Y��s�z�*7}[S��(��l�Ȼ��]4cnf��ZF�E���p'�Ն0��{�n�
`��4��;��F�TF%���Ƒ��"�̰�i��[e_Z]�D�l����t��A=���{JMįw���5T�>7X0���,�����g3x�����c*�%�1�kQ[����q!0(�a��nVLBm��qh|�������C�QhcT���f����L�T�Л�A�c��2$�%"�1/{8S8fS�qU�ܷG�m ;�	W�%,�Ғ⶯��Nr�D��c�&�k��� z^��(n��םۭ��Uӂ�v�X�s^����x��d�3a�/n�zcbPj6BYC(&�ە��ڭ]��M�Hz�6FGו��6*��t�@sA�zͺ��nsA^4�r�}n,2��f�<5�t�F�C2�����5q�wAJ������]	��|��DЮ:Y�r`3�YoM�v��fG�F�j���i�d�+�6m>�ь�l6�'x)=�z�٣P��];S���]u��9�Ry��C1��"��r�ue��3#JMu��`�߲��b�� �e�Y�J���Y�]!�}/��t�;D��Z��{����f��ӆ���0c3)��=��ƆK3�KH#��6��/yA��sK��Aj�J��v�a���-���B��:��}3�K2�$�@�$�e�����Z��Ív���AO�/����<
�V�[8�+���zuܻ.V�,�\�g�;�@�{�d�X����:�} o1ϕoP��;����C������z��Vf��cf)e��_xu)��#��*�`��w� Gu��k�ݴhq�w�}k0R�-p�a�?�um����g�֧�Z��{��&žG�&w-4�^'��ېP<�OD����o�h��;^b��9/��.���I������B����*�qt�5w�3FWM��lW�9�R툟'��z��� Q�ة�np����K��+9죒�+�je�Z�w��DCl ��S]+w�_�kƮ��}�"�F�g&
}u�Q�Z����<-6�2��7)M��t99���e�r��/��ki�y<�BV�ЫZm���{�d��cb�Hg*K�Sr'n�1d�`�н�ftR�)br��;947c�u:j���a��JzƄ>�;��2�
�E(XԮ�f. ����T�6+_Sہ�k�MI0�h�g��f�2�*�*�z��I��T���);
Վ�gmw��ȡ��To���ׅ��]Y�-�
�r�;�ğ8���Ic���&H���hҷ�>�Q}�n�"����Z��˘>P��
��,��:H=��I���󜒮�d��U��x�(�s��p�`L�i�����2Q��K�l
�ȹ���̷���PW
J�K�B�V����02L컗į���*�)�������� wc�tv]�-��-'��V�XB�v��4H�xP��Rݩ�^�q��\g!,��B(�r�hT�80� ��]�����S���ղ��V�1Oi7��=.��=G�r�ŋ1��Ǚ\��Թ]C�o-\��K���bd��kon���t]��jj��2��y�q�`���<h}�I��:�kzRܙ-@��Ď�5�|�0�O�Ǳq��u���]C���dS��i� yr��+�Uw0�T'</r�.�Wj���9]�3�(���'\/(_C�i�3���w+�]'v�J;�Ti�a�6��=�kfv5Ē��P��(շ{h��j��Vo���ݻv�x�v
�8i�:���*Wvv�Jw�
x�Z�|��0kqT�{`�1��H���s��F�4w$�p���ժ�D*�a�^ìuc�y&��9��� pGZ�f݇���ݦ^1�A�<Z�L��\�����f�)��qK�mE4����)¶/dH��
	��"&U�0�}���Bt�r�D���&�9ƍ�v���t���*�T|`�Bq��X"��5���jJm*z�m%���p빇A�.��8*�'@�g���52`o'c��yT/]���*��twQ�}0�K':V�g.���=�:!��ڔx�l�z9����]�&W6�>���)-��Sh�WB�9�����&�.fkb�X�Pq�X9�FY�t�Y��<L,�C��p,�)�8s�ioV��U���4�Α���Rێ�_
*��[+��˺m<m��4u��
s�+���4~=�eʽ�
��s.���L�v�k�*�+�Oa�U:��g�u[t���l�}�Е�\��KFۜ�T��s��qL��p+��s�}��Mf30+2��l^[oi㈙���@�I!!���$��|��s����׻�@tƘI��^-��I��i��q�5�ұ�GWjˎ��Ji�Z�;4��4Ҧ]gV�����֝W��p���_�A��4��K��
��N�Y���Z$��q>N�.Ż�+��/\-�\�^f��g|��w�(��@��}Yf�t6�XH����;x�*�2���նR�)M��X�Yݘu"G�m����	�n8als$��`m�74v�W) B�����8�U�:�y�9m�ňzm��-C�3�+-SN���G65��8uc}�.�yJ��W�ʨ7��V��Ó��	;�qm�ք���g4�b������nE���9��7[�J�NG3>΢�Z/e
�����ٖ����=,w`{l"5�p��7zX�:v��h���K!]z�j�m>{��
˽J��M���Jۨ��Gc�;��(��R�)�����Ŗ.��EX����rǒ���r3&_����R�؆�m {$�7�B����>��[|XMy+*�x�cF��*:ir��1�z-m����l�u��o8�1h�
ogwJVƔ��MKdK�h��kn�̕�;.����x����D�)_#�� �������N�U�9�&�a�y��}�'����Bؖ��رSc��cx�	��}�1-���΅�faM��hp������Y�Z�����J�(�Q���Ʋ� �/����X�/d�"���f�2���Bq�o"��	
�E�Ne,�����Z|S.͵`�R��"������_�c���w�CJp�wuaH<P���{0�J�.?��mS�فE̬��F�FE=�+���L� ��X=(lzV��]���"E,�m���NSF����v%G�%�R�v�S�{fk�uw���˴dm�]e�܌�JҮv,28J��u� �Y�<�Ur�暊�Z��j���.�2@�$2WT�_ÚJof���}Y�za�&a{�!���Z����[����D�E�{�tqn�[�hI;��ըK��fQ���d��>˼A��z���]樋ʵ�M�������f��:8'sްe[���[���V��@N�u�ž�Zp6�z\�!��k2�4)��V��]�Ɩ�(�2+�kw\�ևcK���E71fL�D%
�U�F+������ו�`����A���QǕ��Y��_sR�-!K����(���˷m���bNÙXY�mS���M� ՂY[I��)�^��uVr:�$�%��K���]����\�T��r$�qi2tt��������Ƕ�2 ��q���-�t��nY������3.��9�}�Y�Μ��V���H�or�y��
�Eĵ^����䮶���Z uӒ�!Q��f�jQ+�	]Y����^t<I�}�"�m�Su��Ϡ�T�r�K�f���JLube�4*�;"�o)N�b�s>W��Bq�ҁq�߭iה6�nH3��G-�a��Wr����݁�L�w37E��U\��';�](�u��94�zQ�:cy�DNV�K�*ÙcDH^uYIY|m�7x���.�(jig$o�]����m���.�3
�]u,k/�Hf(���n���`� �����1|弻������ی<�y�1��T��%�W���or�V([�}de�]ۡ5և^Yn�a/���6�V�ZUy��r���x�]�ȵs!���WQ��/[ܥ��']ıD��ome)�5���K;��'2Ye�K�\����sͦx�٘V^[�=�Y(|Ҿ2�栘�{�a�y,��T�sԶf�Mw�r�3H���'Kvr��ewlv]7�]u_n���ys{�Ej��g:�Ai�i����Wi�H@����mu'v�c��uw�`���γ�>ll����]3&�W�v��
�����]���)�j�_q"����U�n
y�O��1�QP�����T��e��h=�D7J�sj��m�-���i�H��mҽ�s2�.�5��n���F��U���0L��_>�D�4J��8V�v"�_+�l�)�����؏f���l�#�Q�C��m7��\C�V_ʙ5 XWQ��q��N��&,�^�}��*̂(C�
����kh��d���LV!z^�΂�m8:�Nn�w,��-����*�Y����o�,̍�E5�MãN�]�)T��m�n�nd�:�NZ��#��W�.�.XEړ��>�;EH��Y{w������,j�+zy�O:��� ���0͉���lU1�Nd��.`��cㆬ�#�M�I��"��ZݬE�B�rX�7����-�o�Y>�b���`b�i�\�Ҋ�[�ԋ��f@�Ǚ���%䁿�j����,��7�[Oh�βl�Ό\r�×�����4n�jLYڹ`U.-{e��u�ɛ�'3���tJ�����׼�
��+���5�m�t�372AdT�3����.�l-�:���<��D���X��a=�+�e�kK�29�^G��]�HH�VrKm���lMu���p�P���K��6,���Oj�\��1-{a&�ѻv;��/��խa�'uDVem�'�Q�/8����f�N��^���q��{u.���ӧ��0pԷ,��M���Y�u�c�����w']��y�La;֩�,��JA��(�����2�A��S��V�(Ә�5�yL#:�2)��Pp�:�M+
��(<�;Ku�3^
k�!:�qkog;nj��ݘ�2�.ԥ�vY���ԩ�^mŏr\�G��K4#�*ѱI�'�Ĺ,La�O.*��r�]��/�<�i�K^�h^/PY��5�����|O­���8�F�	�ʎ̎��-5��L�e1�5�^� �ǐś�(m���:��˹�<�b��E8�ǆ��Tj��>rs�k���gT�ʦg��kR����+D���=��W��«r8��PK����Z2�03)��ld����{ɳ���>Q��s�ݲd����T���
r�g^94²���ci.���&Ky[ի���c�i�)hoN�|��v9��J�!����V0)kZU�S�����1��r�d��
Y�>���k�Y�C����Q�2��s&��t��m�AG3�	@�x�l�}�͖Q��B�=Zkc��:uXE�U�cy�UI���Iۼh�_B��G�t�-N���[��a�=�h����ە؎v�B�|�4�V9�ҵS����z�1aZ���h-U�U.���^�5:S�s�r)���٣٫�]N��hꤓ��P���Wv�E���&�R�r
���X����MqAۮL-����Z��Sw+�R0�
[�p�V
9��T��ǩ5�2J:�����]]�K��f���s-��)�{���X�߄��y�fi,�[0)��!�]1�"���2"]��Va���*f����J�݊N�K�y��Wylc�YzT
5M���t:�i�Ջ���0��y�����GG�ֹ�e��O��뱹
1����
�wm� dn<	�h��o{�z��2�u�����6�<] ͛*�t�X[`ys���wݴhѵfXp75L��Սg����To$\1sK�ǁ�V�:���{5ZT�D2Rӌ������ba�J��m�m��߹S�x�K������p�/�t����Oy9�w�'O��hs�Y�� ���guŪ�n�"�)d�8�w]�vv\F�1�Jl���>q���o���������Ga�����X��l��Ot��Q���Yz���փ<m`��ᅉ�s�;�؏e�ť���K���sl��}�0��ʝ��he��@LՌe�W]Fą8��c�^P�v��`۠oc.�im�6ЇP��t�i]��3uX��K.��N�kX������n_n�L[��:���)��,����j(�c�Ce��f�Z�FT%���>)�E�ϳ���R<�lҮ�����k'���.!Q��;�^�	�ʻ����:�N��ɀ���>�ֈ9g�e�W�k�1�3׊�V_N�w��squ�N�]e�2�EMe' �c@��>��>K���i�cC�wS]��^`��p��D��t*�n��_	nv�]aRJ�D�#R�vQ2DĪ���x��y/d����+vZz��#M϶$V���\�mn��Q�֤���%�����
/�q�4�OC�;���MM�<���v�@�x������C6�o,vٌ���;�����lդ�̾�۶)vwB/�޴���,�� �_Xh<�y[h+�墮,s��ƣ��wG���b�z����Dٱ.ѦD���z�QU�ق.���K��@�9���Cz+�����Cs8j�;� u���A�`�fT��9l[��qn��Ky�k�wv�W ��wىM��Oi�ݼ�=�P]�e>������FK*|~��x{�1]��,�^K�Mncp�ٸ�{mj�a��,�\�2uN�c/`̘�CK��E�<v��yR=ӄsS�6"T�M;�
}K�̏l]� ���aQ5٦+�:%}���!��e�r�x��Y]��C���]��FLǃ!�������SF�W�mwBm��*w��V�T�t�����1�q|h���[�s����)�0%�N�cy+>S���;���O �(#z���6Ŭ*�iZ�¥�[�;��l2�7>YX�v�y��7�`91x�����X�����t(��b�9x�}��q�@�*L���5��ų3�uf*Q����+5͂h���=X�1�M� �E
N�(�[�ӡ8�Z��  �;�m�����6�[��6-Di���D���,V�. ��ۅL&V8�ټW'���tN-Qc��
�՝� ��	���b}�sʾܙ�u�ܚ���잼�r�"�L�xr�%���M��;�t�>	���-\褃W�҇x}{Ɂ@+zp�'�<��LZ��p6��Ij��NjS}r��s�g^�b�*�ER�L���niag!��;��n>J��5�V	�v7�71���Bg|B�N*}�]����J���.̽C��MW�;aYrѻp] T�̂8;��o��p�cz�]�w�j��EZjn����+UsYZP�Qv�K��F�n�T�g&��ÌO��7Ё�5���p���j��y�^J��;�N�8�qΜGz&3c�{���sӉ��>Ě*�Ea���nnt*�+��a�q�1+�Z�w"�����N����ʹ�w��hd�ބ4裊�ݬϵ
��Y��8���z:����X`د��K�j2J��h2�>8�Z�eq�՝r�J5�2�wH��b��Zba:��.��K-�=���R��V�\���֚kT�AZ��W�b�o^���%O��}i��Rn����
�A�X@�������OGP�y�v1�q���Kjqk�E�1$�;���Q7�����$l���`��M^�""�n�a�b��b�H%�]��Ӕ��ka�Jǳ2e0P�o�Q�|ք/t@����d8f��z4jX�a)#�b���p������^��M2)!Z�N�FCS�}o�!���$���'vu;�lz�aa�}SZڳ�\ �Y��Ec�M8 "�>yZ"S�#�����k�mM����(b�R�l��Ρ[!/�_c][�Э�Ԡ�ˡ`�Ǉw,���I�`׭*W�r�32j���
��=��+)v��elO�*j���m��o�Ϊe�nv�Y���ٙ�o"r�M�,;�5��{����m˝�5��--��Ky�R`u�\5)��2���b��1�Nh%��!�jK���e�S6c�;Fbf�u���-�s�,�y��c8�j�'F۷%f�
C��ա�+�_}k��t$ޖB�����#\d�˂W�Ժ��haj�:�7;yj���3y�SB���V��Y�\+���A�}e;TQCI��g���h�z��V�:��n�n�2q���,�X�+_F�[{�s�^I���;oON5:���p�y@X�4-6����.��h�V��P\�E��T��eiu�w���'mg���2�qTO)�qb#�m� ��	�2EÝ�7��e�'NedT%�t��o>J�i<u�.��l*cSuq�ǅּy�Z�.)�n_�)(��io�F��=[s�����,
]3eҹ��@�m*&�J�X.�n	��c/��E1t;;n�F[��B+V��/����Jj���f�KM=�������ӧ}x^�yR'��{�F��TW`N�5���é@O��=�L6�Gb�x+C�ӄ,4���ڣ1h�n���f��@���D��˭�����ُ�ֶf��|��F�L��
1��p-S�����L��m�}w��%ޞ��<�n[7r�:a��U5��8���ܚ�d`Pdu�S���Ә���l�F��,�2J���5}g4�����s�We����]mm�|-J���Dh�j����m�M`�����M_��l��������wmʭX�� �����]����s;M����c��������+Z��,�<���wz�놛N�B�<-}|�3~[2���^�P$<��{�Ԝ���5V��+Mʚ�m,]���˾[,pI�Ɖu��qį��
����Vw��y��0"�m��;\-C������%p|�v��K����tn�m8��n��V��7:���S],�MBso.;���y����+��ϥ��F�=WM)�;v�0���*˓1����KfH:�M�8P�k��E��(J�yQ�,W�W{�ci�ck�*zq�lT'i�R�e�Y��7�4����b�"��mw)��@K�\���٬�Y��9�op2k�*���Ѹ�iTcz�J�YX�a��Ev7�K����b��$��e�`����z���}�� �{@n�vv�WR�ʛ�T>W�!6�13F�Br�艼e� ����y�����>S-�����C�m���1T�� �o�l��bwA|Ӫ�G1�g@T�2EZ�6˻�K��/#����0t��\��K	��s]>Nq;���Vjyo==��X��T�n!k�
�n�-5�swY(�����Rj�6�^��b*�F�H�m��[���zkq*3lY��k�N�R�{i�n�M��+��ukFv�7Vȧ�jwZ�n���׼\J;уB�zr�����L*����f���us��4�$�ر���mÙ��P�(�x>�a��y��g�6��![�k�t���I��9�:�^U�m��@.p�]�ZYVz�9�/��:��ԚV�Ѽͣ�hrmb�K,R�Y��Co�K��.���W�u9��,*C�E�����(E�C�/�eb�@2ɥ�4R�w���Yוe-p�F�ջ?m3Ik���t;��7�.�щ��`v�z��F��8��0,���e����R�u7Ɍi�XF�UY�ec#T��fu�����H�B�^��i.��HtҘ���v_ դn�d67F��	��K����W���z��E�3��;�Fy�>�p�C���)s�����]�ܗ�2�]k����e�U�����ts0G��$:��6��'q��&�RU�Y:/F�`H�F�s\⩊;�0�Rv�A6�#7��oe�"�!f.
aJ�W�^�>�Df�d�A�����,U��L�ȩ��Z ȭB��S-V�PTVJ-�Eu�\ʚ�X��IGZ+R��Le5,Ac)UJ�V�b(�-�0M�&e1���
�TX�B�EU�ň���X�EU-.�aEƷ026آ����"#6ب��*��QUPU��TE�S-DME��f%KJ�ۭ�`ʕjX��C(Vڪ����+QU�Qc��9V��af����q�A"�Qc�X��-�mh���J1�X�k��
��cQ�V�
DUPSAm
� �Z��r�j��**�Z�(�*�Q�*QU2�\�`��-(0PDUDAA������3+eUkE`�YR]�`�����US*R���ģ�5kJ�Ac6��UQy'����}�|���$0�3�Twاoa�{�j����x�<�������c�w�q�-ud9�RY�����}�c�{�%�hU_���')D��]i���,��.���/\P�r�2� .u�rRφ��]i��
� ��HJ�f�|�����]9'0�=Exi� ;� :�5��ƐJM{|q<[��9�}�{�� ����;���V	A�Kt8��JfH�;Wy|��K+{�(��޽��#�Y�8)����6h4`��KF8E�]gao�7US�5=8Ѝ�B��g'���YcU�z��{�b�ϱN��"w
06.c�"���e�A��}�:�����x\��1��e'�"F�=��Huƪ�-zoE��ˍwP*��e<������ᷥ´,�����y �x��@8:׃������	��T��<�y�#�$����1�my-���bb�ֶ�����G�lT8qx���:�z�ƶG�_�yR���}u >�z�tz �q�L������{|��c^np� G
y����trb�F��l�y���]#"�ZE���g{&"Y/f Y27�V��O����b���7\q=~v˼�AFb�CMj�!�ow$�V�����rz�N��[�!���F����x��XsN��i[�[�����sٲNt5�/(���z�>��E�Ⳉ5�0\�͛|#�Cq��3�KuWh���2�F�_b#���q��tj8\�C@f����/Cw
��Pf�O�:�8�rt��F��iɝ��-fm�ש� '����.1�ͫ��=�: d�	��c�3_=���T�HpJg�~��|4z�um��ȡ/�ٿ69\���8�6sݒ��Yց���k����jd�a��Փ<d���A)��۵���<�T(�VI�o��U}�.�� G��DB%I�P����Q�7���8J���<�I����Ԫ"	��U���n��X��^��z: ?����S�^]&:��>�K弧s<��CV� �ʂ�u���\'?>2�+��:0����3q�ђ�u�=�Y�)�A;RHO��{ؘ��>��_`����tԔ7�9���	1OU}�&h��c���:ʝ�㖓A!��u��.�ڋ��q�N���L �a�&�������"��(Q���vv��W�}޽�<R�8�9C��}��W"�՞��1�U� ���C}~H�wWC�M*��+j�mN@Y�Ko	p*#��oQ����������)s��r-c$�wC��n���zh�<�|k*ڙ��j�wo�w5]�o����t~s'+��]���ț=t�Y.����A:������ӳ1u�xJᅲ�˹������WϊX�̇�BW(�-�3Bv �pHe�{�Z��Z��&�e��u�j��{ư��ry��:��I���#^�nP8^�����d�=`Ϸ���7K��Gu��N��yMU9�>w���2�q��|�|wNQ�h�k���S�y��7����h��qT����K+s};�,a+M���鐪7f�?g�ļ7~���'vB���S��݂C�=U{�[4�|�.9�P�7.�����
����̡�eYAt�.1Ľ0�xyU�.prC�qd�tm���g����ҕt�1���� �1�8�<�lZ����lP�e�ffWXE鹰_e��B�j�3�YW��j�1r~���r�q{�A�Kv��:�(���);�Ͱ�,��d����EgW�VW�tbw��:YB(����Lė=�!��L9��%ofG\�k�\a��gQ�r�ܖ#Dpeȳʤ���t@�pa�0p.����ƟGՖ�
qZ�ۊ��1B�y_��.�b
;�'��Tw5�b�ΐ��*g�Op)��ҙIbZ;pa/i���S|�-c�-�G�pw��)1��-�o.䄯D�]˫i�ɘ��ᘶ�m�$�x@��F�|0�os�\]�̋+����c�|�U�f;��π��ਯ�a.��IA�r���� ��t�1O�$[,fw�P���Frw���]	ٸ�s�sD�ٔރ����f�>��=�uᑩ��>�������d�y��S�ug�yb�BPQ�D0ڐ�e��!O!ky������v�@�	�J�͇�7&�R{�%Ӻ��ܑ����ֳ���17���8�Lw��8wUdJ��(����1�3�a�0�צë����({�r�ɾ�j�f�7ϝ,�
&���녍�j g��7s'��f�CRI��,��!B�y�lmf砄�pe�����vF����ڨ�R��[���r�^�n
?p�ho�컩.�[�j����:�{jX��Q��&cEFt���jC�����*zc΍n��O3�+p���?��9�<}MX�=�,�a�L��F�p��p\�@xL8��<�nc�\S�)J�*�ɝ�ָ���U���'���j��&*5�zk��Π�$r52�3���҃�ǫ��'/fM�)]-�{�1����源
�Db�n���̊�)TD�|�a��2eĨܺ��(3V������ɧ@��>i�aMMqY�v^jX�X2;��mj���h�G,ъ�2�B��t��>T}g$�4�t	k��)�[m.gV�!���S�#�P���n�3���Hk�Yz&�²Q]SOc��Ձ����8�~|��]V@�r3��^jGR����at�����#J%�d�+8(-Ps�
��qf�.T��������N�iF�|t`|�$a���_�~�1NP��r����H��󫣤]:�P���0�6�E����6\�	z�ieyÌ㱯����"#9�H	�R���A��mu�܇�\ځ��\<�d�r��^��=��\.��lCw�+�͹-�%噲��9ߎ�k.�W�}0�Hau<'����̔p�Y��R}V�PD�i��Z�odvࡀ~��]�0%%^���\�G?��"��.���|��ȑ�6Wp��#<T���J���Rf�]V�6 N��UFX�A�Ks��V�N�^��	�����hT�3<,�o4��c�E�(�n�C�g*l�� u�%�vXڝgw��!�ě�W�l	�yu�S:�j�>���N� �K9(^�F.�S� ��Ol��N����t5�.��J0N� C��e?��m���f����աA>���;Q�_/K}��W�f��
Q�$��@�o^q^�TA���Q�t �ƙ�v���a���,��6T&q��LU�%Ӑ�w��[��Y�&��^�������w.t�GW|u�[�)��ݽ���\ݹ(�e�I�;O����i��2�u����:k�´{���mrs���Un�� ��jC[����CY�9d�ޫ�b�Ŗ�k��r�Cx���q����ó~���[K��E�Q�5�!����G,�Q7���/B;�z�ˎ�;q�ۦ��.e<�@��7�R��圃W2ϳC���|%�k���[�p�͹pҫ5�����z�81hņ�2��x��]@B��uF�o@K���6�};�
���ȡy2��>z0��qp�½�=��u{j!��j)Yvo��=&�S�m�U\kt
�U"�lDH�:ˬ�x�f6����=�.��hf���z�h+��v��x�m��q�Y��P\UH`�,GK*W�Q�����9d�X��Tz�&>��=C�g�]��X*�bt�j(��7�[8�}�;�AۡY��P�1���ٺ��1�Zu�����SRD�ˢ�!��:>�8����wNl���ʔ����hcC@�x<u��C�Jq�7K����\����@��i��
~$E�S	�/(�V r^`���8n,.�"�N�J�f��2ܛ�on��l7I�����zfD��w%��Q�pK���0�`�j�vS���k0i!���`R�Z�Ss{��n�������u�eN��7���w�^�k�n�q�����K����;����TI�b��&��S9�֓��
O�t�;8^�B��*vbӟ������ �y�X7��W�ln |�6����4߹Սu�E���}g��n��
�<�+��:�*�҇FA+1��	哖��,K1㞪K�MHk��{q�g~��3�L1��K 1Ĭ�rLnA��W����ò]{��o�Rxh��b����̿/���ux╏@�nP2�aN�Y�α�h6� �@�b��ϻȋ܆y"6����*�J�V��Yq���r��9��_n�ohE��h
��q�ߡ�������Ɔ�H�;�c���N�/Z֐�&}����;��8r�]2��ߔ��=�	�m������q�+����U�Q��J��'R�m��qٺ�\)�+��8Jⴐ��=�Ϝ�i�:P��]>�1リb�S)�s����`��p���T�&�Q��SY(s�V8(�0c/sr��B۞��N�W�����uZ���<$�5�����n/�T�X������F?-�0vԺo�TmZ���@�
B�⤢{���ߔ��[�^>>�J�1�k�o�[k�v��.�*�D�[!���\�R�v�W-&��A��C���ͥ�LMÛe��¹�Ϡ��
�j�g��obn�VVVW)����Q�
�[��ulЪ���@�^��(PϔY���)q�!��/Ve�w܀;f�*���P��EdA %4\�TA?f	��rxy���/I��1yT���qs��]{�tپ1�K��P�Z�uȘ{fb0#Y��b|Oa�oF����o�޵��Gd�5�P�����ƈ�m�ұ��*�����B�,+�@ˬ���/�M������!�+7����]!��J�6{��溈J�����ZO��S�A�:O��t��[Q"���+K �ul��>��I����*���QۉE�yڇN�_�v����˥{-`���
��|,:�oki��^�#�ܱ�=�qzq>��ມ�n�R8�%�̓6�ܘ]�m1Q�0A��L�z����B��5�u!�oYZ�q�U,�#s6G*l���a��+;&�"�+f����o��S����z.Eژ���뇈�2�x'�߷�u �`R��𻖶�m��Gh�!�ξ�7�k�ܮ��xA��e�ڨ������F�Wl�"�{�gV��/�8vP�-��5�\Z�G������l��)u����\X�)�H�c���++�����ud?%|GR5��u�S/o^�6���\�vE���F�ݢ2L{����{����j��(�y�4;Jb����:�Vg�U���٧V���H�6�=�ٴ \^�puCos�L8yqW�CT�J;�YW�GOךe "Da1�c$�q3��bl�C/S�¯OmKu�iNƽFߌ~����Q�����/F�ݴ�H�Y_QW�Z �9U���y}$"��z$��O{�H2�ƨ�����TRon�<r�*���Z�UnUs �xڛm9��bR��p�.7��_HX�f��^~��� +���:�$��Ж��WQ8��$��f@FLj1a�ߊrv��h*�-��6X����B�ɉH����[���)��J�fGuo0�NC�%�z���	-V*v�ѣ�:7��K�:cMj XOP�Xm��k*H��m��a�p'�r9�^�hAq��׺jQ��N���:�*Xo�o�-�!J�c�[&��V���CA�6�@�.���O���Xk��U\)V��W#O��&Q;��k�,ngip�xF�c I�P�����+b������c����Ae�:�(���?�V<������\�w�V�I̓�c�|K��7,I�jF�S�[�4e���2@uab�cb��&M0W��x�k�:Ƀ�L�%Dޭ���/L��Ҳ�rY�rv�7�5̊N��*��{���d�B�3g*�[8�k��4UG�6�
�ɾ�t���cR�C9�Lp���Zr��[Z����'>���W������ÍH�,B 7�T��Ϯi��qH��"1c�=^���^��-7j���8���PU����0��Ið�V��6���״�uӌ�Ep��j����y���D2�wJ�����H��E�Ψ
��S96;&�i�S�3�[�|6랎�y���n68����"8]B��A�th�����W�b��7�l�203�88Om�el�J�Y}�HqY�]����O���0V���C�1��P�Oۊ�pa[��]�D8�c*��������k����F���+��lK��;7�..���H�FiV�s��:s0�ծA�鎣c�5l\a�ۯ�MCr���'�-�������/]��9k���reP�7��
�?����:hu���i�e	f,p�1}�
:��Q��.*��j֥]�ۙ7Ʈ�J�*.y�/왆s����<��u����;7*�
WEڛ� &�'nv���V�}F������ վ<�p�~V+���Z%���#���^Ts�%y)t���m�X�)-�n�C�HrzԵ�p�_J0w �g�uub[M�A��� ���N�Gjl���5s�,�]Cb�aA����Gq�ӽ�wu�\���ۧS5��ޡR���� ,�'t�Gh�u2�"s;�n0��8.��;ᙵ�����B.�'Qh�N�Py�@�9XL6{(V��l{o�^����[W��7a��\�1�;\��j�<��������*F�8 �x;�CD�O%��>��������@�0�퍌��%�0�۽�nSȐ�jR���ɺ6'����W�ev�H+��s2�_`��U�^U�8He�]F�h��ڷ�欛c��Q��k��{'b�.u4�y��u�ZMc�n��Sg�wqE"0ڮ�}������ T���Thhn�v4kbY-�^�����_I�~�.� 706��M;ڱQ6��Gi@�]��V�g�|Ε��U��=ػ����m�Ա�0s�]:P�dv���u���P=Z��?X��.d�Y�L����:-v�V�Nek,�%F 嵛s�vini������uݚ�\x��SO'�]:p�b@N^����Zhj��ޓ�&)�pmb�vV[U�el�c"t�ά��q���BL���B�� ��u��J���tjRoZ�厎m�R���}1}�R�7�1hS)֌���p��R��y�'�O��5zѢU��	��Lu8Yݎ�D��M����J�h6E����f:dW;LtW��+�Sf,3��b��h�M�ԉ!�,ju�7�c���Dq��sR��ǜ�;U���|�- ]gT*�C��D�tӺ�K��J�r�`N�����8a��n����m��S6TzC�\�&�����Ԟ_bl�y`nE���V� O����r��jb��<B��`�캒0#A�Q�N˩�M�;;��mZ-�
<kcllu�@�{�y�\���b�9���}�Sg,��+���x��IyANh��Ƚ���Q�Q\��֖/���F,����u �ve��}/����st�$/j++���H�����]&�P\yN�u���ZUu�̬j�@03��Z܊������S��e9�3��B|oy�1��LKu����3}]�v��x���N����n��VH����U��N����."����R��r��ns��y�nԥ�V��p�[���X���b�;[���}gp?CWVz	=�T�͔k��y�U��i�I��+^����.�
sr�y��c������u,L.�e=�#��q�骳q�L��YA��:��h���-���mA[�*��a�q�}}¢v�^:�׻f�	��Z�$:�}ϭ��Ok�O���+MN;�qx7h9���MC�q��;/���qUka5�B���ca3���v��m��. ʶ)qg�4���h@���v�LIIf��v^0(�S��q0��ݥ�I���ޝ�&)r��Ѯ�iԷ[�٩�z���Jk^
/��]$��X�v$�=�h)E�;�w���1"
,Q:�\ƬjUQE�F�X�jS�Y�,b�M�c�b�۶Ͳ��*B���V���8�D�+��2���A[E���a�� ơ[AV,*�kn�UEJ��,E�h�e��Cm�ETq��+U3)�r�B����e�\k��U�Q��	["�Jʈ���QQb�UU�DX��
1id�icR��bkQ�����ʨeiETPD��[j�ĴmUQm�����QkX�̸֨"�jRثX5���TE���b�E��U�KaF*�%���e���(�U���"Ȩ�(�(��DV�B��Lh��MB�*�*"T*���(��M�)I�Q1(�EdX�)*[J�V(��b*��dF �A`2!YU"�EZ���iB�X��EF�VŖ�&U��AkmZ�l���UU*J�R��Ĵ��(ȵ�R�@�5�M��y�i����R�����f^�+��oKrTjÝG�ws���*M��8�7������#�=��3EO�qn����[��R;a�g��dY�SN�$D�?��92�=�-C�v����X��6���OP*�b���O������W��TDI�xG��>�DF�\﯋b�8mT}���_��u�:C�&*O���I���^�ߘf�V}��>q�Ag�ݰĬ�P?������P�:���/�>N0���$�C��G�8Џ� #�����ab�߽�H���~>���MMCă�Ꚃ��1�ܼMI�1�'�}�$~d���8��9}݆>큈Vr}�N!P�1��m�%H<��)�
��"'O�x}#�vN��:�x�>��X��hxçt��7����'n3�>��H*Ó�x���+����Ɉt�}���k%eg�����H,�yf+1%IY��r�RW��?S�oL�b!�" ���<%Nt��ǋ���KΟDq��Y>�)�O�+Ӭ'hk��c�,�RW�/�6�=a���9���bAz������c:�rM{@Z����@�X{��|�C�D)��������h���� Dt§��ӈq �!�u;����T���J��ɉ�(t��j��=B�2w��i�]`b�����1�� ���rMJ�U&�}�������~�ao��1~��Ȋ��ѣ�|D���6T*q���1���Y�x�CR
���r�'HbA}{CY�vLC�(z���*c�rm�Aa���n� T�!S���8Î�~��C�l��J1�zk��W�T�P��@x�&?�>=�3�� ����+g���fP��0��`qa�Ğ'F��=IۏGv!�Y�(t���*NuCX|�!�tyx����>"-��ٕ�k�~cD}B>�">����+?$�+���I���:���biS������+�l1+'�+&�ۆ��+�'�ǭ� j��i��ÞS�������d�1���0��fI`��mU.�{��	�C�z��{`W��u���?!�J�����3�|�'���}�H*��>���Ax����+;IY?}�v�CW��;ߴ���K�ѶLO��#�~���S�n̟X|N�^��Y��W`��O*Q��7���³�����m����i�>\�d�Z������"�U�7ـEG��٢�R�LVQf��zY=��C9Q��Q1rس�a�ǣ�P�X���t���Y�!�ͻ�6����=H[�xkCW��[Ӫ~>���C�:L���R�zɉY*��옐_�u��i�v���|���|��$�1���+<C�bϾ�IĂ�ߖb�!�����
��_Rb0']~�q_���}����<}';I^���Ö�����ĝ~�9:�����(�3��z��I���?!�'���ܐ����3�x�:I��Yj�f����J����>��� �����jO��r���L���5:9g:J�Y����Ԙ�S�3�%a�WPԞ�_���?a״<I������Y�%g;�$����8np�|��ͣ�Ǻ2�lӈ�X�!���Y��At��޲M���Y��
c&2�����D�?��j�^ -L6���@�P��3�>C=�v�H,<a\tǄF��� ����c1Ѥ3U���?ng����t��g�+������J��0��q ��K�ߺ�$�
γ�{'7�!�z��`VV�����g��+%W�`bAu�?'��0�0�E��<"G�����SP����s���v������Af��1><��jAC�>��8������c�
��RgGh
jNЩ�����N�8��a��'��w�k
¾�`c�X��<C�ǄdY��P��#�T{7.=~>ʍś���~σ���3
��ݓ�1���@�=a�ruO��8�Y��xԟ!X�qĩ?!S�������=z'w���p��l�=x�S�W���#�>��e�&]J��gN�w���*O�WS��7��>��E�ֳ�J�e���'N3������7��|�?��$�~�>�u�5 ���N�7�&3���R~~��N1�""+_q�-�Ǯ���K�+.w����R�yd\gl�O�1 ��>9f�I�bA�g�xÊ�IY��=MC��<E�$8�g���!Rz�y�|�ί�gg۞��+#����z�A�/��-���6��}�J��w�5H)�Ϻ�~LN�~a\ga�a8��~La�;6��H,��;��*AM���;MCp��XT�j<�=J��/<��M~��} |��vF��d�q����N��R*ێ��<����/�M��Hr2�I޽���lp�p6%�݅C���\��?
�5N���;
ً�������&P�Ѣ¤���Bm̭=�x��X��:"t���O>�\Y0��@�>���aXW��N�sE$�v�ɍ偌�����6�?3��C|��d�<˯L
��<q:�q �ף�$�
��嘁�� ��DGo|{�cd���Z���w�߈/�;C���;{a��Xw�5���bS��d��Y�K��MCRt�~O=���C��'G�Sd��tßs$��ۏ[�I�휌1cG�D1ᗵ3��g{�o�G��'<��>�q�2_�Lf'<�b���a��t�_�w?{��C��@�}�>u�����ށ�P��d55!�~�e�!��I/��b8G�`��z�ќR5G{�]o���C����'��WY�%�큏i�&ZoΡ��&3�J�����:T����k�����W����0��Y?'8����eCT���w}6��掀�X��򎮝������z�3��$�IPY��Ѷ
�Rt��58�ɉ�T=a���Y�ݞ��+
��^P����=O�gO�
��_{�3�'L�g�߰���/�Oݘ�e�2��1ơ�m�Q���}c��D6~�8�S�Ă�^�Ğ�Xpϲ��%I���5 �@�3�0��Y�cgo�1���c'̪�P��P�=B���|���xɌ���rwNm�J�ǭ�+3+�#�ǋ:g߽��AO9����!^��ɉ��C�g���k'=��u72,��d��]H*�D͡��8�_�u2�5���S5����׆OI�j��W�$iqªX��� |w�x§�:C}�!�Vx��u�>J��+���i�����������Rw��hq�����ў��%ea����
�2T���T��:���:�:�S{��Z�`��C�����z����<��<N�=N�OY�z��r{��U'̨x�!�}�1������I��Rw�`jc��9��k+%W�
�ϲ!��}�ϫ��՜����	�{g1��s���F������׶eI�v0�~�P1'�/�92�Y^�Y�����OS�ă��ݕ'�~B�v��'�����$�N��Zq�0�R��,�A�tא[�����!�>�8�Tމ��te9R!�$����o���
=����ݻj:��x��zy�J�akǂ��ڳ��%ut�u�lK���0!jf�a�̽����[l≔�eXu7D�Wn�Ko{s7�GK��XZ�+���z��������_!����d�Y�p��P�<NM}O�3��cٖOSQd����M`����|���.<����t�3��v��h���E�dxp.�� �5��h
�E�E^�j����#rzIɍ�^<w��t��A�߾�Oe� �F�{�a�剘��tt���GE��Hpӑ;��&W����?��x΃e�.�hk����p͟�u<��Y$<nvF	܆���mSJYH�1a�0��N��j@|TK���WNOV\���PC_BU���j=t��vW	��cL�F�*�F���,j(�ng"xs�L���싵����Z���ٜ]�[����G \�b�g�)�p(gN�5H	��ycTj"��;7�X�+�2�q�x���E������B�[V���҇@�8k��a�Q����y{�Yˤ�g�^�s�Ww��l�l�U�ᔼ������[�O=�|8~x� ��!�Uf&X��Ç�9z�㴝h����P�zk�N�.paِ�wX��_�!q��UAT��-(Z���ܛW�
�cZ�Q�^q9&9�-A)Q��w�iv��jB�����p�e?{-��u�\��Xiט�Z7�V:����Zv��gFۖ�J{��CY���6��R|���e?�ĳ��hvZ5�k���6�Na�|1H9>ޏ�N�p2ˀF���ʶK�[��J���4[�gL�݈p��l@vSx n�&weݾ���.3�Ԉ�r�9�h�=e�|w���V�kϨ:�*"�b�l=n��k��I�Y��tAq3@QZFE���L�z���e3��縰���Cͅ�W=]�M���0f��W�m��t�SU��|y�>��X᧵�9�y�7:A{�f"�N��+I��C���'�,��TJT���b���:��[纀|��byy���ip��8crF�(ئ雅��B1�#�fm�����K�ksZ���ih�������j�9��C������.Tb+��dāΣ����; Q��UM���Y�ǈ�9�0�'�כj��/���3h�9/h���"��T 8��D�B��*�7��ۄ���`8�}��Y~���d�n�L��>l�J�����엑�
{����vo#G	�ͪ�t��V<���]P�a�^��((
C�mHf1�Ce`�.�f�6D�*%��󥔱�M7��젫�Gfnt�*ΊH���T,���6����b\)�8x\�����x���2vc5@�`	�z.q�yoc�ř@� nT��6+yn��Գy��;�x�&빾�
7����iTUu{AR�3��+/e`u��P��!����r���,y�Ϸ|6Bu�m�U�{����٥d��_F��f�b~ī-`�s�@F���s��C��zG�����(_�;"K)�:qzr��}s�\�\>7+$\V&ӣ\'z��t���](\7Ur����	�)�'L2H�6&�šu�i21w�`�]�;}���d�b1���2��vq�q�;�����El�~MQӣ"%���ڝ�tȧ�m1�k��O�m�3���1̢�-��>�k�X���$t�u�(~5O�r
\mo�p�.��N�9��V�d`���2��p��T8D�(��޺���w!j[9E���wg�*���׏��g\1���0�q�\��B9��2��C�m,(q,X��t�j��p����k���k���C�h����
RY��-�C���]�W�&wՖi1�Me��K+�7����2�1��:CEzWZ/����O�Q=ȩ>���3&ak��k;�����w�t�X�����Pپ��c���>�#Q��q8R�ɤ7��;�4w�8N���$��{�c�<���6eW]'^��{+\�m
�DGuܽU�+ŕ �����>����3F7��R�� WU�O�b����m1Nƺ�\L��lQsvP�l�;l��I?�@�!L"9�K�;�q9лe� ٬�
��6b���������}}�ȼ	;q�#�joLX���K�}������$�c>ٜҝI�]��\үX�!����WV_�m��&�_����u�lu�S]"�t���X��j�м�8v�wZ�pͭ�S�y� �X��E<�1~�=�ᴆ�b����*�<��.���.�Ku�Cp^�|�� �C��]~/A����Q�d�xOʟ����
���CS�q��Ƌk
a�ID�!�B�T�*�c9�6@��tQ���;s�6��څq�NMҠ'��̂{���ʩ���-ne��d�QP8SuXB9Sf�e�2��I�:.��b�glԖs�@�;��ת=��KᙿSB��y��d�n���S�'�8o��I��3D��i`��볳[�S�D
���vtWmEaٕ|�yO�����b�����q��\U���㞆�75�%�^K�Mz��1r�e*�D��_�0�ҫɹ8 ���!ʱ���\��oqS��x��Z����s+�ۚ:���]� .YaB�&k4�֌*ʒ�@���^"a����1`�+s��5�v�t$���\o����U��L�oE�ܾ�m8���4���D!�C�K��)^�W����,�]Z�`��z�X�#u���]#���6):tn��� �\�ڬ��2���dִe��>��}�;��*��Ϸ�G��Foc�ê�iz6�X|���v'�<����.��:Z�cgOWg\N���U��㬧����Uѐ��-Y~n����+���]9l�PGw{i�L�bi��w2� ;2wOXLwy!�O@�n���b8�wc��:�PB�U=�&2҃o�o=j���{2E��F��e���9��M�|6{
}q#��^�V�9�6ɱF�Ǫ<HH�K�*]� *�#b[�l�	*�s�_	��S6Кy�Fvݫ{T��U����>*L.�Ѹ0x-��T`���\@(;��(A�&$�Rֹ���ܺ�!
�HO3"E@�鈦�5=�2�|gԺ�N|L1�ܷ�Ʀ�����B��"j���e}r��(������@?��r�����d2[7�m٭淶�U̗�9�q(f�L*�O+kTG"M�"c�@��;�=4��أ-$�#������������ה��\�&M.:��B�r#���Q�*����׍�O���߭Cwq��E��j�;�&z%�t��>�V�����w2օ������%6	j���%��t;:��5��c��i�-�sJ;̛� ��[^�5���llw�����7��(!RK�,�]���Ҍ^�����+��m��l�WM��d�Βzu��Q������\c̭i�]N�g����#Y�gwmQ�o!��;Q�Yٔ���՝�FC�]Mt���y��^���Z%�����
���xQx�t> S|xV-E7�Ouw+kp�V�] b˯�8O`k��ȳ�g�}EeM>�A���ה�j�Y��*�c�Nn�<t ��g�]p�����c!�ϲw�D���	��u��g↫��JwM��zq	+>��:2"�f�L�����~�;�7(h}rx��v�1qN���5���U�m��L������
��Yxn5:�W�1q��N��El��u{�8��7
��}oE�L�Y�C�xm�����s»����{b��Ļ�@�|������F�Ǿ��a�`v�pk�N��yN��q��zhoS���CF)��4�% gi��E�ya��?.5�%�v�T�EKt�B���^A�
�F���N��msX�.�纻�6%�4�Cϒ�~2��Ƙ�޴ަ�8�y�ne˾r���ޚ�!�i)�dͽ=�2���뼱:�+m*�ڭ�6ȕ��"�1P��B����޺�i��%ihykaͨ�T��W��6o>���N�����^l��P2���x�QwʔC�b'���2#0�����n{/vjmQW��^蘮�Y3��sՠ�Cv�RF|ˢ䋅!�+����s9��3���T{��7bi�7�OY��5��{_��%8���`l�޸D�T@�욓�W�������'` 6��;�b!�����odl���]}#	�Y�.v�����LkÙ/��R[����@/�ׄ��ڭ)7^�V��C��Å�X|-�k��Cʠf� �d�;;�]��o0��ՇvA��nKG�UzѴCDu�� �zC����2�q!�e�����:�DY�Q=9�������t�$t�,u�eU��ꖬ*���g��Ɋ���%�l�R��@	](_*�`_Ѯ�:n!��"��0T4$����. ku�&�ji՞���,g�����@	���]먌��8o�{b�["�]��ь��B�D8滟q��H������Jj�^��r�#LV�����%2�Ўð�u��k[S�#6�Ń2�cqO*���K��!�*���;m�[��Lpu�2�/i�ԆP��v:�8��[yU�J�DG�m;VL�q�[n萛�}+~��ܾ��N�1f�����m�5å��1�'j��YY�T{�8u�z6E�Sc����w@�6�"�\)(#�;&�&���J��VR6H�y@��ӡ�ٿX���	>�f���h&���3�^�����.FŒۼ,KtZҨM�N����IH]wRk[kud���=%vmb˻s�����y�C[���G�9�Uo�m��ō��ZQG7w���dǼ[��hBo��b����_5x8��(\�J*uv^��'xu1�v�!���o"j�T��g�I����=��w��+�Xdk>���+"�ק��X�|Dѵ�(��3�R@́�p����P�7����Xr�+U�]]γL�]O̜�RѴ�wG[���}z�0B����Nd��o�|�_k)&���3�X�����jűln9r�Iv*'ru�Q|�ou��kh]��4:S���M��L�{�=y��V�� E����@s���S�C��)�c�һ(�����v����
���P��Ru'��q=+fR�Ŋ�z,;�2�g	<��e��C�9���!/���-����1��E>�jҳ�iDή��c:���U�xL����9k����F<�:k:���.��u
jPr�F;��7\�f�n�\��	(Mķ*�(�-\VBDu�����O(ݗ����ے�������������]f�vc�*���2*U�l�x-3G��BL;H]Gy����mcx*�d�R��n�m��\�+8b���:���A<�F#���^J��v�r�a�B�V�	6�h�K�D�����f0�4
�P6��]����@��Ո���k�G���xԆ19VU����X���	�NL�F�)�>��	�+��L^�
LU�*ۮzug6�`�2T��N�R,��fQ��r�7�D�e��Q��Sl�S@V��[Cbj�u�ҁ��$uT�c.�g۴r[e���5/$��޳K�eܛ���ƶ��j*�q�v;NGk�3o�B�!�ˊ��({�%Ֆ�CW8�L�lܵeq8�ջ�/�w]���5sF�zH�����D��]�"9�9�����>}g�P6���8�^F����:K���݊�p�׹8`D���&E�y�z-õ�������6+;*ӦE�]���El��]wQ���b�B�"�*�A��<ʌ�R5F�s ��ݷ���GE*�F�퉫\Y7��#����z����m��[̘-;�`�Va���Lp���*̎��7�/,�IQNA���[���κ�7LoL��F�O/�]N=4U=r�n�vފ�2©�Q�γnUҧ��k�8�B��-V<!P�.W2�Vh��W{�M��I��G|�A��q�5;��}���h#��:V4�W-����|�v3S(�+E��>.Z��v���T�fsn��SyT�{�_n�\�w�����m���q+"��o���^ޝ���TDb��D'�X�)�U�"��`����i��eE�Z"�c����m"�ŃkmjQ�R�(�J�e�5"�Qe���*��[B�6щ��E�E�`���U���EGP�1&1`�*Q�Tb��++
*����1�"���ch�UYR*�)YPQ`V�
�1Tm��T�r�*�0`���J�l"�.Yf5kF�bE��*�J�QTQ�̅PdEE&R�R(8����IR�����h)R�DTEb��Df%dU�`�Y�-m���H�ň�ʲ��DJ�er��TAA-��
*�Qb���PPPV�

-���mTTE[e!��aKb�qȰP�D�Ԭ+U�ł�[r���* (�UUD`���J�eUbȢ��E��meX�Z"���`�b,DPAR*�D2���kj���R#�,+
�VV)+�F�B�:�i����g]~{���]5�������j�����T��B/{g+w@^���d����;�E��r75K�\�I���}_W��W�Hۨ��*��d��s�:|��!�z&\��
����*�*��%�}x��T���x��S˛����M�,:�90p�a�Y� �m.U]��΂�@J�\�S'���X��»r��i��S���
�J��-��CB�wP�\�P %;�s�#}*[�4gf�W;����;֠I�\|�t�ن�����t�M���d�`s��w1#�7��U��ms�*cz�?�dL:�C�vK�}��J��8B�iW�ț ���;��^d��`���ˊ�"iL1�ʞ�B�\��K���g���d�}�ܻ���R�sܕ[�gjO���m/i�T��׉���t����;� ���C��"���<ܫ��K� �ZQ����5�w�LR�o�Ȫ��KUן[�~O��Y�^Wy�8߱�S4���iof�k9nሱ�wcd�I�(�vl����¤^�*��p���ꚺ.�ЊU%�g&;�of[	UK7 #��S>�r�Ϳ�a�σ�c���:�=Wn��ˑ�=��X�ں����Ɔg�I�癨���]D�,�Jݬ��>�b��D�}�M9�#�3��g�Y��4 ��j֭V�d5.Ś�Ԫ�
�D$+b[![݆��'y�9�����aڸ�fC��������� ��]�ԫ��{��[�T�g�^;���.��.��@��±U}_r{s��g*�o�e3n�>j$��TL ��X%�z���fU��4������};=Λ#^ڵH����ƽ[�+�5X6k|@�8�W�W�'g���Z�1\mH{q�h g�Vn�Xh�yX��Y�U-0��p����r���ї���hL���m���V��k�'E%�>���C�/OmKy�V��?d/gY��{1.XB�u	��ΠܳŁQ1ٓ�-$��kQ�%�ΎG8�?TF�xo��3���|�p�������G�����X�7�d��M��C?�z�����y$/�[P���� h�7M�ܱ�T�=�(�u�F]�����7G+G(�$?�� �"�EԺ`Y�ю0=�o1�Uw�O�tɮv�7���R�=#�*/x���T��Q�[I'|v��	*�p�S�8{N��4Ѫ���Z�Y�-#���渀�����D�(���
�DDdu%��>�6Q�)��qf��q�gJ�Ӄ/زPRm��q)���D-�h�n����2^�ZWg4��̖�[
��Ľ�"�d�\�����.��g�	_��ǵ�$��1u_.�k;U ���5c/�7+8�*/^#��Jnps�qT��hj��r�E�>�����.�;��*c�MDJT�\G9���u�5�!K�+��9�b:�x-��TiE�F�R��m�ǭgWR.��cDJHS�U���)�7�C I�P�г�]q��u���$��a��Vp~�_2��,�#�-F�l;�R
�����X�W |@J' ��4q�ط������ �VPc�����aO�\0��d�+Z��!q�9�dt:���س� ��K}2�n�pU[���&	e\2Q����xS���S��-�����@u��GUҵ���ٔ'ON�M
p���h	�_�+�ʄ*,�(X�8k�J�����b�����3z��J��z��:Cܿ�Rxk��d=��>�D+�}�B�����t�<�Ž�,��\�<�����7|"���.1鯩,��r%֍=9P��*���')���b�q�����!����D1��B���+�GM�ݢۼ����k7�Wf!x0�����\�W��W��CD��)��9+�J��.���{�9�a��1�Z�r;��1y���s������ް�Cʯ˳�&�Z�U�]�o5�����@�U��\[Τt�8( ���+v������6S��7�����|4�ƴ�A춎��R��}qު�K��Q�T�r����M�ɱb�&��x <:'+��G��͢�+1��b�|(ϒ`O�;�Y|P���U|�͋�.�3PUUj����s\;������)�?B7�ͦ�
�� '�}��}��*~��.{]	/k�YُM[󄄭;�X'���1���0���zˈ���})R&��1��V���������!q)�GX`zdTغ�q������`g�x���{|���coڶ��-��^q5�A�#��n�n��n芀��"���	U�vƽK}��9�C/|��>X�B�j���\1�f٩6�@�吅jw�%�	����{��GyD O�RV��v��;���z���]9�s?=::K+yJW���.�����y'[U�"n��[����t8_�`��k���jɿ.�4x=�߯���^ɱ�55a��.~�P��"S`RӒy�BU{iM�\��C��]�[�厮�е�_Z�mF�ϰXp�l �̲8��چ���}Q��6�O90���W�aT.WMJ��5�vn�"��p6�Y;j�wx�1l��gB���>��a�u
��0�|p'F�Y�jn�����?���`���� sw���3��˂��'P��nR�sJQ_��ĖL���e�8��L۸�{�y���<�ՙݳ�Ќ�ѡi���\ �H�\���z郦�[�B�NthVN��s$v��=��:%jg�N>�~���g��b�xk
Vr�([6Μn�������#6�����v�	�3H�|���pwU&��':F�sFG�X˗n���j��x)�]g�6��<Xg��Wj��ʖ|<,W�yZ���5�j����_V���$f���]�B�ȩmsT��bv���u�P+dZ�N�<8�!�e��
��Ү%�|��g��	{��cj��F�<�2��b�a��][/Ģ�b*\���D %�����:j��t����z�;����\H^����av�Q��h�7r5���7��R��@Jh�@#��sisY.��ݺ�����9��l�R����4�+�5�6lvɁ��o�d+�N�0���t�8��hM
Us M�`�dL/�X�9�g��zh4r;M�2���.}��7�:9��%���W�k��?vVWB���f��.
��!1˯�ȉt��'����R��9�������ˠ�uB��ڞ�{����Lk�(���5S���̼�a�PD1���#�I᫆�����A݌�;K&%������J��e�\���H�kX1��NB+�TjAՙ���/���,&��%�u4E
�"��ٖ�u&�a���� �����f0�� m:�~�������;j�֩�I�:B��]�Hb��v�;����8�R�I���g*�Ͻ�{Ȋ`m�ޟR}<f�t����s+Xf���"v�ٮ>�c���)]��.�
n�1G"�j@{�Ug  4�S,v�A��y
����+��>�=�Һ	e{�[���JgY��`�P�Xw�M���L1���H/[6ʟ�{w�̰6���H׆:��9Y+�z8��ݮC�=��17��
g3����K�}�\>�S����I���4[�V�.}k¹�aپ"��O]�ǉ�����:�1�ӷ��zI�'���ڮ���s�&�h�����n'�g\Mp�'g��*a���UcC�t�3<���&x�yE��+�U���[���p�����R�~��/
�.�&CDl���o��M��{r)=��O�nڑ�ӑ�a���hqy_\���gH�5&:��>�Nk��p臞a{XU/r3,r9�*��J�r���tƋ�Wף+����6��Yu�k�8{5Why��l����[^��Ң1m�IL㮬�g0q��u}[��;zr;�o��'�{VXʥ(�j�^�;o�Ա���f�!����f�1��������0em+���M�
��;*�j.������*^:}���t�.G1-qs0$�_� ��V��+��1�1@{�U1E�bBgV�.�V�]0��Ǡ2������]"���w0��Q��dS����ypQh���C��#]��EVӮ��O_B�X�^+�Zm�X�wG�n�B<!�ezɥ�sh���(�m=ňk��5��t��Ю:}֋��fQ�>�ꮢ� � �6�S�(���>1w��<�rZo{O>F$�y�����!�t7z���A�6�CD58H_	�Ձ�YڍT)����Vܪ�`�cj�@���[9r��py +��d��a�v�2p']���t{��w���\�5�w�y��r@�����mP�^P��8򎘾�t���=�3�4u�'��O�-�Kz���\��3^\u����"8��Q��|��ŉ{&����ǣ}U��%� ���7�9,p����b;\�3YH	����L�on;���4z!��x��'�b���醀=g���&�/J��,A�2�u�ቇw1H��ߗ�����lӟ��a��e;�&]�nӎL��6����sI����j��7��:G�>��m5�7|�I{a:2�[�:��j�n��!$rn�7[J������ZU 0F5����l�:�1v����;!�yo�� �n�+3 ��꯫��V���a�0�	1:@+�Z/��"�<5��kEw�#�ӵ�����\���@Ü����_fm�������@W1�����T����	`���F��7���Vsr�~��S;~���C��d1���&����P���2����Q�/7�'3C��k�}�e%����X�X쪰/UBܙ���|���4�;	�eq�cf���m���yK\O+������G����[�F$�g4����efK���o�gx+�d��(ip�.w�y�l���5�iC�'>CT�;�y�=�ۦ�	��Ӿ<���;p�YYP���뗭Kbc�t��i��l>M���k�ϛ1ň��U0��,�e����貒����6�6`D����s����Ju�r�� `���3;���0�2(]��\��w:貹S��m�n"��<O3�y^�k����Û�c���tE��Bu���޽�[%N�L�Yj�Wunτ��Vv4s �t�+BM_����\���w(i�.b��ӻ�v�ya����/VUB�̅6��{or��X(���s"n�O-��9�D���b�mgZ4c����XB�S�^6��u�$w*�efD�e,	�3��5��B�4�
��Fmb�˸��8����Ж;�z͸�eΗy{Dn�  .7�7LE[�$!�~��/N��Q�w+yS��
��}u�����-Kv|��gb��`.���m�ђ�7]s�uc���r������T�͂�£��ꧭ�U"{�����MPf,���F�A zïn{�_aߖ�q!\iey��9��y��u9-jJl�2�T0�j�q6��'/�8���N��6mVÜ3��<r*��02�,G�?�?z,�{HN� H�r��*�`^�@鸆s�� !O�T���mOsp^����,{]�.�n4�c:�Ε`_1�8��&;:���u�O�kss�պ���4�+����p��+vkY#���~�/�ح������'=�	�p�F: x���p==�myc��(2.d�r���\�J��K�z�!�C&_G����%����3�:
�������m#O�2Q�6!!���N��}�0�;˯w�ff����c���_S�_Y���/�����E9cT�pTz"HF5��~� <@O�@�Y���hG�]��ъ�zj���m�u���aS�נ\eix������s�A�Ӛ��81KW�XUJ
͠�2������9��KR7��)��-�X��p���Og8u�������.nNr����f����$�^��K_ ��{2��wC��7%��ʯlVvPhat6��zw;���or����QVK%��$E�Q|��w5]f�
0�����r��$6X[�����پ�01��Tg��N͸(ƻ�V��+{9��$k�23d�T�I�� 8�5���;�3��tw���[�ws�bž	�3�䵇��6\+��F(sĹ� �A�mz�I�GE��Y��B�WB\f�6�I�e�6�Z�|��7�nG(��^} 5�@�v��|��qۥK�g�ԧ��W��3�B��v�Ԅ�,̷����D�mJh�M^3�!���N����;�U>a��V�>�F�x
����T�'/a���Kӂ�mp�[�)�,E
�� �)Bx������x�ixnJ�ܠ�u���_���X�z=�)�`�)]+��-�J�Y�D��9��]Fɢ�5�JNݴWK�{��th�eWi�0��M��;[7���LA�p�tֲstx��y�n��e�`E�7[���2��$Պ�!���^΢��ʫ�3�G �P�]@�9��p�J���O35��%�fƂ��+q).9`5,v����]�V�i�V6��{|���f�3Pf��)��:��ܿ��/�{�kV��32�� 跢N���R���5�:T:4鬰��墒�e.)�v�}���l�0JaNu�nZ(�ȱu���q�WQ�6�pM�㔷�W�Z� �˓�r�w��*��i�U�"�[C5"5ݩ��q�D$F�RT���W"kd���>�>@)m���CNr��`r�X�z��5�l��"�vV�9�S���z �qnlsi�7��#��}���\����D��'�r���Ojz��e�&�W p
��r�wkQ�;��,%��c��t��xev�̠D�įW8Ү������fӧ��(^
��l��2�k n\F��uȽ1���
�	�p��qD��sR�����۱k�n�6��e�@�{Yb�m^Hdj�	WAuv�+�/a6~�}��h�H:��t:GK�ݎH 8q���un
�w9� �P�66y�f�n^���ٷ0���܋p�-|f�W��w.�I���H���]��de��yY4_>T�qB��̻w�գ
���S��M�P/4e�ŵX��k����yK�˩�B�}D>�8l��r�Z؂K���n�j�l�Uu�h.��L}�]����7�U�*�YX�see@����H���re�U��"�N�׷����f��f-�������(:&)�y��TX��\T+��N!�;���
GA\��2gYJ�T�¯��/Uɫwj���t�\[{eWh�i����E�M
oOw- d�C�lQ5.b��_w�Y����\�E��f���Q5�}*LYĞH��s��2�-��2Q��ܫ��ȡĦ�F��jZ�ym�
:����*_j�(V��9�l-�����A�6M��B[��;���l�c2�q`�4	s��5u�x9Te=�#���F� ���Kt�Z�m��V3+N��t�e�P!q!Y�9�z��VUt�Q�ky���d8e��i���q�7}8��{�w�B��k+���8��-�-����R�p뢖@����ه���܌�u�]�Ͱj�N�F��Z:���ڝ4akj�vY��?4mQ�xЎ֖�6U�IæF������=�Fi�\wγ�Q�pv(xVљk�h��=������F���fVl��*���v����P�ٵ�#�$���-ZT�	2u�c�n�'F�l0T�r�	֒�p/;L��8	}���6�`\"�b�)WM�v�e�5j���M�5��z&o.Z`��(�{tK�����t��!��ꖩt*�n����p=�QҬ�KX��)N'�H���!`���t�����V�9\�k���,��29@��+%Aj�����-T��U�XR�µX�����֊E����"��.1���H�2�EbȊ$D"*�����c��`��I�X1�`*�Q��U�dF
��J�X��̔T*E��U*�[LLATEI�XʐP�
E�ŕ�k
²��QbŶ�"�pDh�@�XEm�#XQ(*��QA�J�dc���$��EY�+ �B�CU����T��P��
+"���FTF6�YEUD�"Q���!Y+-IUm���
�Q�Db�V���B�P��҂��QjQR��6�"�Ulb��+*,mU�����ʪ
�رA`�V��"��"�D�*��hTV1�bA-�V	V±E�(�YYQ��T� ֊[-VE����
�s*�,X
#&"�+?^n�r��_C��F��*(z��bq1��ڧ�m!��� �(\��tJ�݉v��,q7�h���:G��ч�U^�������%79�ަ��݊�0]�u�@f���gʸE�N�	W�[z�.�\��i�c�u~�)���*M�]�}w-�NP�k/�g=�F/�c�9�u ��S\�]oܜ�Y�7Nu�՘��.3�u2ˏ�;zq�ږ�حO-�_|��ˊ�V����1<ީ�����[K^j�8�CW�1�j�P�r9U}Qy�Jf;*XaMmp��hV�OW�!�,��:z�����M?�W �r��1]Q)BL�[P�8�ZcD1�y�b;��p��&1X���{a�s<vg�ã�`v]6�t���]ы�)��M&:���8z�F6��f�iĸw{��WS��+��hOBo��]ꓸ�~}%����$���-��]L�=/@�9�w^���v�^�<����vsr�j-8�Ҫ������F�:D��͠GZ�R��U���3x��6:���^�Goј�U���=~��k�������Xit���1,"[^\j�n�>JgO�T��5��ݎv�dAi��Ƴ�[;;/�^�/	�њ&�`�d���.��X� ���Kq@#(v���s���Es���]j<%ꕠB�7���*�j3W���ϝ��
�}�;i��״��] Ucݮ�S�5�]s0,��y�պ@꤬����}�UU�I� |��:{Ƴ*/GWa�Ǐo�wz¿�f���>)�	U�<&e�[��Vg9�yo(l����nW�vһu��d[�2-�ڇ���2���$�I���}�U[Lע�i�ν���_^=�z(4�Y�h�|V��o)rg;2T��wy��~ˋB�϶����3H7F����}���pm���!�њ�����^}f���QZ;��7�H@����8�����R��:���#�c����o��������l���\�ZVƯU]VqV(�Z^Wڛ�=܇{���1չ����5��ZuK~m_�hy+�(��ݤ�/��*5��i���o�	�b��8%weUod����3��.Km�&������D?j�健3}���O�ǜ�f�wϻ+�kX�.��H�|&�ؚ��^�Yy�Ŵ3����E�$�HI����Du�����*d�ٞ׼�b�K��H��b�/`��0���L�(���X���V
�I��V9�5�m!��5�S�0ɚ��!�9�J\���߶�םQmuB:>�A�b���SnIq[i��F��DU�3�} < L�O�Gs�{7z�JK"7�8�N�����Gv���BN{8,��h@ާ�v)�?��{�����ꢟu�&;U㌘�H�7,��	U΋vr�a��s:�f'����*dn��}�q��n������N�|n���:ŏTTo}��c�)�������%�X�H:���^=�����W�*¦�Ev��}Z;*�V�D��p�������f��6o�9���	A�V��uS��C��GF�cG�m�{z$s�;��@Ӻ
��]���˚��۾�R���\�7u����ۇ�M��9�j��xuוە�u�U��;�q,62���s�BWn�IqX�����p����u�:��u��/��Td���]�{K^��(��a�*��yW��=G�˷�4�~� �N�(�֊vr��r����;�"�)�q{TS���b��1FM��v�d7��|����:'���e�e(Y�lX�Z16b�2q�,��a{%O/!xg%�:
�zb��>I6tOj�,��WǞ'��ZY�t����}Wq̒n����ظpO����$�vރ�N�yK��}�}_{�LL��^ձ�dO��m�����qv����:c�~m�Y7k�ov�u���v���9�!�4���Ǉj`J�/.4�X[N��H��z�=��QL��ng7kF0k{����}�b����`>���	tM�4�8�����1��qV�M�̭+�3i�ȩ:Lꙅʵm��ԴoW]M9�4F�^��%�j�#�T�.7nW>XWw��V��kC�Ƴ�����[�������E���h�k�7(�l'�m���Ƽ{v����E��[uTGT���iI��+���=Aj�}�wO��	s�W��įL�[��s�±�ǿ����Z/�ѽ~��+�=~0��<J׆�$~��=�o���4_A�ge+���_��9�QZx����W�w4���7LU1'�>թ,��Cr������>��X�E��|��k�����k��l�{>�}�+�4*fwΜkGo���ǻ��fy��9h-��9�g!6�`��ņ*�5uA�uA�w���4a�h,������d������Y	���� ��C��X�ep�D���5���}��3:hۉ��k���;PcT�q�ov)R��7];yNn=�n�q�n�dB��?�8ؘiz7����T��ј������153_,�6�i��Sơ����-��ͻ%H�5��7a8⟻�����/�7��E'�R�aw�����/���s�M`ܛ���):/j�By�/e�oF�6�D^NTb�9�:[�S�U�U�B(�t�ѭ�s�{����p�,z�߂�|��OQ�}S��ɸ�nH���?C����%�t����X��5�t8��W78��n�\�U��=��z���Yˡ�:5����s1�~Bw��8������5ix�ū��t�Ȕ�a�k�.�}ֻn]vf�Y���ZؕN��1�:{k��Bo��4�՞u_;�T�Ҟ.a��\��c%0��7Y��E�]�2�0OCaّ�sD�kh\��1�/m�ٙ�h¢tއ�=ޫ[�m��A��K���a��Rb}[��z�Ȯ��������G�ݤwW��4�Y��X�ƞTv�"2!��e:3�23�=p���u�n*h#��eX�8�����X�H�A,`���pfR�V�� ��v}ڴ�u6Zt]�t��+*�ʵ�=b��[f�-�j�HU���d)�[�!��8�{۫/w��f�o�p����9o�2�B�W-�2��&�x�����}�ˣ��4���rw��8���#�l��5��c�E�Ց,K)y6={��|��\��7��<^w!�5wXt�CEȱ�sۮ��k��z����"��q���p̿CS�������k�^-��'�Mp��i>��yg+�R�#yi��lC>]�l+���*���6�����!����Ow���T�YO�	��s�?�.��'1��oXWs����[����*<�5����e:�l���+e�y�y��W��S3�x��kgjRM�S�a\�6䨯����T�sÔ��r;(�z�f���KVR���Q�]�>�QY���t��orj���e��=�x��Pi1Q��l��9w��e��_���9lN�}�}۵�l���1f���� ��#��,'|�=9lh�lpR���~��^�հs6����n�]ǲk�����oe��:�@��/h�D���o? Jnu��u*�g�p�-��*��O*W��]�x�c���8R���7CO{���K�4N��tD�/%�57��'`�W_��着�	������^���������^]S���y��_|{�]�Ϛjp��cȇ4�F�y\�Q�|3/:�9�-�j�³��H��O����#�u�h��0���,��S��Z�����%�i���sD��U�ϫu����8��y�Ԫ)c�-�.׻}�ʬ�nWvG$#�ʜ[�Gv<�,H��y�x��T���S���u�{��2~N��a.�	CP���z�|]몦����;�+�\�tV�	�t$�瑧r��3]2��45������R��(@�#3N��Ϯ����U��+#P���������^�R�U�@ᛂ'\%_Օ<�ypfXՕϝA{^�
�#%�ޞ^輊��1��U��*����td���o�4��곩��N3�:���Nv�+eCЮ�4$k��=��;�ۥ�kƬ䲍�m]_���z�p5�&�U|�{���qV_��Ij��{�.�s�0 �G3:�/�zV�ܰ���:��hCi��t�SV�С�ZY2MO�3�(tw�2�v�N`NV`����-�UUU�/���W�>�̟��
�D9����
�w��&�X^�|wO,n�����>���?��ՠ�F6�S��\TcC[6��T��u{qәPN,��s֣+Egx�I�H�݆�0F��^J��41�\�p�&4n�;R��4u^1=T�ߖ�eŴgض�R�����zݽ#5�=��s�t-��)&����g(�3<�ujmב��l[�0��,�YY^���ʯ�]��)�mo�E׹W�uچ㒌s�B�u�m�Fk�e��Ж�6������ړ�z�l����%1��bU|������R��ջ�.q��w���V}��ZН�׺�����[�5K�;����©�X�;��(Z3'\S�%uF��_l�����S4����o3��2���Y?|�?m�Wie.i���LEn*�ҷõpMTԛ�.�nQ7LC}룤 ������72􎖪�d��\�,�-�r��2����6�kf�CN�-sZ6�n[�V_��zW����1VzRt�j��ڜ�Q�f����U
��.�X���.w7�t�C� ��3����VH����1��kv�Ö�A{��>xx{��/5A}	Pϥ�|��.�7�h�?�HC�J�1;��W7�5��Mf�8s]��:&��Y�r��e�#�]��yֽn�e`�T�e�2�u[ֵ�lB�[��mwEln����C\D�m C��tr[��EQV�%W۬Z��{�do �6�������ȕL𹖷�X'�yΦd�ò��f�("S���]�qc�Փ�AjbvP�#Oa����'�(���ҹs�]�u��;=�S��!TR����r����'�@����r^�W��g��E¡��8^�`�k�=쿜�����:��ʌ^b1A�ⲲgY���2o�ru(]�ܩN���7(����.��r�F5��NgEX�/V�`K�L7[}��;=y�{��hI{��qs���ν��u^6�&}Q���k]P����}^��}�_3C�\�N�u�k�����T�kL�g�b�ۧ�CO���F��ڎ�J�K4�n����k|���o�Ҝ��F�+�}Ր��Vq�@���Mv����% �R�CEK�"��庭=:�#Ep�����HC4�Tm�`-n9f��8q�"��fv�������:�2��^gUg�9V՜ڋQʾҲ�7��۟kTGk��]�`�qs\p�Y,U�=V�:�Ȼx��КՍ�׈���9u�)妟vD;z��d���ڽ���>�Aի�=�מ	p�;ɠg4Wk{r�=����J�XS3���R�!����2���pxc�b�y�yz��K��ӓ~��ƶn�'�.6W��܆��Ր�F�u'd�j����Y�e����m����75���/�5�(�q�N��N���}�Q�5�g�6Z��孚���뿠%��v�[�;���C]QmK�M����⇺�n��ssVp1�Z.V�Xo2�+��.j�
L���>�ZSx#p1EK�eΗu��n�����%�E���F,{p�H\���A<�
�u�>ݤ�h[��{�	��*{qN�����3n�����˾��(^B�7����7�;�lm��4)*6�v�Ùc"L,M��Z��VB����,�,��P��wҹ���;��%����c������muN-��Lf�Ga1x������BV���W5t�	b�n��lN�aMAs#l[����=�+���I4	;��)S���K�Ǣn�4��7Yئ�W7��[�ݑ5Õ�"��@�����d��Z�cj+L��]"z�r׼���nLIL��q-��X\�db���Mюv�o�$:�[ãu��� Ksӽ�J��G+��>;(@N\�[ytT4uD3D��t�G�J���B=���jt�gU��Q_-bڥf�;.o+h�7E��2�iK���V�ƌԴaɬ�襊��i�\��䳂\�ÀO�o�&����Yu��!5M䳵�;����$�P��5�t���лU|��i͵���^d�mm��ܭ(�ײ��f���qe^�s�}��,��\"y���m1��V�u��gDʼL��A��uWCq�^�s:���]��H�V��+Oqj�\3�#Ue��<��LZ�T�O:�.��v���^gW��}�g�z^�^ؔ�|����T�m+����u�um�z�e���)i4+�Ǡn<a��}�'�0&��l�=�t���,�V�y[NS]GD�ٻ03�3(YD�\��f��>�)G�ۿ���N���v��*E"R\wz�[,�_���f���X:\�˽膀m`�a[����\	U�a5�J�[feb7q<oP��h��w���"��l���N�<��N֌�ŷ�t�K�Z��7Iu��;1�ާKo��S'ܨ�s%vw �z������s
@8hd�B��aG1E�[��EWldl�ɲfWn��7e�`;/�3l�)*�9C�kN��_�!ؠ=��5�>���K3��r�(-��!�Z`��e�^WC1�}�;p�Vi��������f�(����h���(kn>a��ʘ��G=p󙧱�q��	�����i�@_V����D���\(�:��Ui�������u�w-���T(�@�m�WQ[�۹ܛ'{G�g"�'m�]p��;�w�+�Xha2F�C{\� +w^�t�%��̩�\����n���˕��uIƜ��+w+�{֮�;b��iI����y!����8`�z��u�+*�t�VeϦ����!G7p۬N�O�'���I$Y��t�MPa�U��	N�^R�D��c���,���*�֯�������UoQ��s��o"�%E���4������������V������m�6��ޡ�ƻ�Ņ�:�Vt���c��7��{0����b�,&t��㷘P��W���hU�1�Y���K��1��H0����@����OG�e���vo�gN����ց�wf,�C�T�S��U7c�T�¼=Mϖt�m���ptRZ�������:�)�G��8�광F�3˶����L�H�G�؃�K]�ޮ��]�ڈ,Fx��m�Dm�Ub�����E�lR�`��bR�+�E��#h�X��TV)D��H�#o�+
��ŕ�aT*TA�YTUE"��X�j���FE�QERc(�P$XdX��AB��i,m����J)XKl�Z��YJ,PY"��E�#l���6��f0*��JőID��VE�D�VJ� ��F%�+R*� A�Qk"m�����őbũc`�R�Ȋ�# ��Z�*ĭk*6²"��YXUH()X)R�aDPaX(��2�V�)P��*�*�dU���J�VT�H,�Jʌam�b+�6�dPD1-��d�",�d�<��\�Lk���u���{Y�3T�Q	�Ycb�[��u˯��ۭ(cq�ћzl9Ǘ���o*Šn���6#?G�C׻�%gQџ�H�oT�q�^}�w׳ѐ������+�H��֮n�Ի7��N
��A�:����-�򧝛���uGeA�b�ggZEl�CO5���o|^-�9���
�z����?u���7��-�+ma�`F�E-o[�l:�w��T��ڡ|/��<.���s��kg�e�	Lc�J��|3�`~M_���\5�s㋴���:S�M�x���T�S��ŝSIm֧Zl\�vor�����wp��ơ4+9�F�#���.z�qzշ�(�`国�����}M�;��z�Ġ�#�Pbw�b�.�ΒWʡ��;{X�&��R���F����ݶޣ<�pX�)at-���OVa�7�L��D�����R2v/I�]���H=��YOc���0�,-�l�c�;��#����Td^��������B�Ȭ�^��}�_�T����CU ���%�J�uS�z�]#=��r���wS�᮪�`�Y��h
1%�A(�9����=�]�Ed",Ihp������%*4����d��{ki��Qp{Z�n����+6t�ȓ�	ջ��M�we�a|p��d%�ո$*��Z�T`��D}|�bͩ�*�wY�q��G<����	�����/JZ�79�OD�H˱��&�C)��W�
�^�Nv�z;në���s�`�7Iܽ��8�p�3Cpw(���:��ieE�+�r1=�{Z"�EU�As\����#q��m�/�����i��l��Y���˔�q�qnbB���'+:^�LoPu�6�=��D.i�q?
��u+v��K�9�v[�+ܬy}o�ջ��\ZlmD2�f�N��զ�V��>4�ԧ��E�����3��Jū�1~�]�\��� Vd��{�!��Wk��[&A�O]����\HQ�}���}X�ς�6*mQ	h��u˹�]^A��>w�m���c�U^�To��uų���>^j;Y�mfc�H���z���:��wٺ��|�Aݎ�w?E�!�t&�������̡��.�1�����ٞ����~;* Mi��l��vk��˄]`���6�5)�y��Yit��Y/�=��}
D+[8�k�j�An'��>���m��ӏ)f`����uÔ�V�D��]+l���&�1R*�l���ﾏ�=��p�p�l��'oJ�n��or)��R�n}�u+�\��e���G���{ٙ6��y�=���iװ��/��n����kE��;�c��j�ip�@��;����o�r#��s;�5�׹t�V�4h�ʪ0�gQT��]�aA��д����y>v���V[����,����Vj���:v@Վ#�d����e`��G,�����HC�K��C]c=)rh��O7z���#\n����e��$5.u#�z��ؗ��ON�])�7��B*�'ܻ�}/�����¨�aYs�nw�:�i$wӽs��~%�N��x�I�����:����*�ǖ¿�A���T�L@�{y��O��wn��O����~NgmF�\�p���s��Pp����U��.�J���$f��ڢ�i^�X�ޝ봸�u@����J�xqT'. ��.,��Ջ��u���Z��
`!��ut"���n�:��J*�N%�
��z,.��b�v�.�X���+���[k6�)V��vѼ��s�N���T�#M�blRy�#k%e#����>[O���w�C`v��v*��Y��=��^NV/1���9 ^����z�	�ݕky��u�|���/��/K�X�E�>|P;)U��f��f�v:��|[��]�)΄3]�Ŏ{�jپE_;��z�%��D�(���.E�ެk�7��]K��1�6��.~x����ѯ�%|����u7��8�u������M�gM�����F��T�c���y��F�|��䓔:p�:��Z70GuOZÏ�螯N5	�Y���V_;�R�'z�����֞F%���<侥��ˈ�~���7ʲh�\�Q�pWkz._W��_Pځ%���K��}ʖ�^��}נ9��]���)5 �+����W5j{1��4�-$�VU�NS����_rѰ���4���wc�y����u��>���TS�N�%|2Eu3O���dsC�^��U�+(����~�^��%B�R�_j�C!�"�D�:������:��N���da;������J�)�@#�M޼�xd�z��.�5�R��w�^��޽{y}� K��}�+���(ltH{��؆��N������e�#�b`#9�S����@N~��GW7���MB�h�A��K�[ך��iy}&�я�,�+s!;��+�a�'��L�T>G�.ع=���O��Ӛ�ޓU3���N�º:�͋w؄59�%�V�M����Uh�<�[P�Dp%l6螜���]��b�b}U���=D�b~r[���F5� ������}+L!Wh�������^i�4o=�OE8I����KAF�D�ҝB�.+P��է�����\J�覴.Do�}ʴ���|]���YWo��0F�b�og��+��h'�F�`.��c��қ�et�O�WF�R�t��{���{8\��5�d�ݩʎ��;v�9j��
��e�aU�Ocvͨ��|��#}Vƺz���D�w[ʽz|r��������u�5�[߫�V��_,��Wc�&��kV1lY|�Y�]����J`�L�{���́���[��oɴgcQg���h�L�kHr�v����)�����XR�8�G;o�=�Jo{5�kz�Hlr��F��.M�'�@����bT���P�eѲ����S��s�s�
+�5#�"�=V@�r3�G��<�sR���9��z;r�;�\������%ׁi�2���k���rV*Z��|xK[��;��5Z������t6���(�+5�uP�x�nqPUͦ�I�/2�b�X8�$Vv�B��[�4���������8�J)`�\3r%������A�Y�$Ԕ�Z�}����������λaJ}^�^�O�u��W��0yٯs�vt����[����ve�:��U�������_iF��X�R�W�C�+z��B���l��|-G���kc������D���[I�.㩻�sv�p.��m����7S
FnR��]�KaZ�۬c-�9:vʇ�\6&9�g����4��v�& �l6[���[��"��׳�o5CCvs��k̾qF���{UZ�EdF��b��;��}r�v/;kV�8��v�Iq�����,{��rC�y3w=��n��nF+V��V��c�����}FV�2� S�/fQ��KKw�{o$�����
����Y�Ⱥ�����5�t������|��F��U�@�h�&۶)�}���R�u�	�'fpR�m�#�E�am�����L�����I�m}U_p��L���=���)�q�[�W���'���5Wr�u������z�t�Sm8;K��k��ɨ��� 3*���WJoit�b����	�U=�Zܼ{�ѯl��_w���36�y��V��z��9J�t����
m��u�]��x���\�Z�f�PO��s�-���Pޏr�s��#'�h�z���Nt����3�@#����>�@v>ܞ��9[i����g0ڵ�*�|�K�ށ.�(���Τu�E�,i�}��o�߫�C���d
nghĥז�x;���S��L8Y�pKbEv�������A�vfde�n�VE尙l�Yg�Y�*�j<��n���&��)>v����t���]l]W:��oB�1����W<әP�&9_rB9*�<9�`\�v$���ˋ-5\����5���\��Kj��؅h��@�YS�;4��;z�Y�n��L����՞3_�<� ^b%尻��j�]�@(�vs�e_:�o���b��Ehu��ws ��uÒ�M_C�ר���Ч���2�Nj�ûM��Fu��j�wѺL�M��ftnl�#!��O_�
�\��έǅ��m���߆�P����c�|9z�T<� u��Ւ��3s�l��l8<6�^\ݷ����f�ux>��Ŏ����p�q��T�
6���빽���X�4����>�X�VO�}a&������u'E��tj۹���[��5�U'����}6�]�xb�aw���od�y/����K��yZ���9�aX���%����;��xo1x��Ù��.�Qy7��ЕDÇu��:��Ɉy�4���nQq�Pq]}oR�w���Z��;���~�����z��/KU�}����R���/��������ֹ�?�����]�yo�ud<��w����z	�ʭvk�4<NҨ7��i�u�z�9O)[N�7ˆ�����#�ލ}[��Y��Yy��W�z���s�㶞	tkcT�>��H�#�������5�b�Z�sh8�82�35E7�'�07'5t�q��Ĭ5�Y6�'Vj2�ʴ0�޶��
Ĺ���`V��އ;7�?d,W0;#:m_w��$y�O�s�76��9#��9�fӱj�3�zL}��P�m���q&��Dʛ��}\��I����8��O�zS�ՏW`�@� &���m�-�N��Uk��ngb �<�k�;n��(l����-�U���5�w'�̝6�+w���S�Ogt�wս͡�71_���������ѡٵam�ܙ��d���'�^�"ɹ8�]3�*�SJ��'�EG9R���㞅�p�)�w֏C��m@k�n�zvf4]��>�[kp�Gsy��s������H2S����1���AYv�'�s�:�����㠻���޽)_,S��t����v��E��t�:��bǰ������h��S�v&����5^|�j-�3B}�q�U=��;�v��ɹ;�؜ҧ�������-�*�AWu���S���Q�ӗ�5�8ov+����Fo��\���ܹ�S�bb1A����P�T�sÕ�����=�o6z\�h?3�5������1�J�J>�U�KKH����ޫ���b9W^��"���b�;U=�pm�V��Z��S�	z��\O%�#�|L}z��S;�KW9h�n�ab�n���J^\��CM��#�e�n�ʡ�QnN��*�ѯ�_WصOt��S]\N}ܩ<t���a�cj�����b��v��`��o:�|2���I�����o��}@���N)��w�Խ�Գ溲^x0u
��v,砑���w��i�vq�xz�5KR��o���C,����n�e1+�f�~�OW6��I������j��mF��>��#o���c�����
P�X��hN�4�e����R�����K��bu�"$�S��û]i��̡(vf�{ZƝҞ^8{��څ���h[_7�ۭܓ�ʔh������N�a�AW��+7�t�b�x�.���鳈U����y��n3!�N6�R������3X7t�=<��N��mw��.	��:�շwS��f\c�P��s^Ϊr������2��U_DJ�g��5�#8}D͗�,�wo:����������\�E9ds�����ۿW��!��ry�v\i��pۨ�G|U������谀.o��4�#9�/2���eܾi� k�o���]:�F��K�1��rkb�Y� ͍zR���/,��R�ڬ�4�۫s� \���2� ·լJ�l#�5;!��䅑�-m�47[@9��}7�[CA۵5.<�m�z�eՇW�_Z�xU��t�����Ns#u"�̽�������ե��0Ø{F�lm��ͱ�U
D9�}�l�	���o0��̩u�W(	1�� �-�SdH�#r �0��Xaʌ8��4&����>��/n�V�ұE�j7�as�Eu��T��+�y܍CKhv��E�b��6���(�s�m+3-�(�[6�ҝX[;�;��n�>�w��I��T�hh-V�1���*X2C��:�sxu�qv)y�X��S�l��#��ի���R�썮���܇��=�T7�Lw��o�I�9�1�I�3Q�٥Z�YW٭O�APU��Wa��ҭݗo7v��o�W -�21�F!�d�ǫ�Zs6���@8ښ�d��#��O�������ٵ�e y�8����R#��P3��L�+L�jĔ���g8��,mf�tN:��.�J��]lFvrV�R�	��ґ��<4t�r�OJ.��R���>usz,r��u�f62;$�5��7j��Lt�%��u,��'dWt;s"C�U�フ��{�p\E�"t���gn�\G�E�r�F�c[��W��sk���T�[��m�ٝ�4�.y	�N*0P�<�pBK:qQA�c��6��9�
�SUy3b��I���t�7���3XE���vnRy.O�g7W�k/��T�Q/,�ޭL�6gX릩�/>�lw`
c�u�"x��ۡZ+2�����T��3u�����c�4
�ҕ�a�!�n�ND](.űR��?(�gDMU0�I��:�y�җ}\���Uh�C� ���Uwf豱L|p"֖�8+�<)f��_q[t���!5M)U�኿��W).�	��a8��}�>y��ϱ���q3G!�����`˺��ݳs����ZH���+_t����{��\h�s'B
@���b���V2��J��2�.�}!�Oz��"�a�s9>uer�vS��˷E���b�H�3����epN�&���� �=���ֱg4]��n�#�A�n�ηP�ڬ�3��ť�J8����58d�y���5wմ:.�Ȼ��MeJӝF�,ڏ"|ޮ�i����� E�G`ņ�U�#E�{��f!i��>�OF�X��#t�&�u�
�	�p�,�:�N�u��u9w�>�es|gq͖m�%�.��{{Ke�8[y��;� � �Ж+4.�ˢ��U���]��-�|e�M :VSp��6aS���}����C�Ƶ�a7��]m�;@Z�k_pB��Q�g�e�Wo	/���O�̻��#��9#��w�kV]:�<�m�U�bR�9ܗrK�u�]2*�f0�����QUH��P֙J��K1��@֥[d�
"�B�VUX�`�"T
�e�@�B���q�X�	�EQAH��V�fPXVT�(b�Ȍ
�YP*AU���X�c+Yn��,C�"�Ė��v�m �&�m�T��k*�U��Eְ�B�*ZP*�(� �����F,�D4TP*c!P�����[	XF�Z ��Vc֊�eeT��Ԃ����J��"��ZR-E��"�+��3Z�]��S)*E�UF3�P�6�*AJ��P*��9q1-�@�1�YeQJ���TZ�"�V� �Xk��m�eXQ����d�%aJYYEE,D��Jʊ�Y/��Y��-��y��0��i����2������a�2�Y�rC�y�t�F�i4��dT �g�W(�^bxV�ӕm�����w���xΜ`_f��y�q)��57b%[1'�v	W�}w����j������l=�Y��7q�w�.N_C*�p���j��K�y��%?l.#=vL���B��Qjo�i�x��􅚤:�=P�A8�"�YwG�n՗a��}*x�+�1��B�]^W�CA�-�u]`=�¼/�`�����1׫&���\����z�츨irx���81�����ap��C�q��M59��n2�=̥�W|�1g����u<��U��s�˧e>� o7Q�|k�e܋B��lWOlg�s��j������+l��g����3-x���c���-�m��VFm>��Q���qu�.�j�|߼bt��߹+�#�\��A�r�⯣���n�9�HLߧJc��R�c���|���<=ǸH����%�V\�:x2͉���xM���#��Es��Z�)�>{���ʪ��F��71�j���#`��`p��(@�l�[�E�m�AK��upYW�.g�J�͕jU9ӫ)�aJ������u�[�:s#��;�5�솞[��d�)q./c[YW	��$��t�bל�sέ�OI��GWj���ME�:��5n���|���S�}y7><;k�JC�#=-��������C&^�ۢB�+^�EpsÎ��)9{�=�Gq���a�MO�ob��h[�n�W#�Y�Z���Wws�õ^8ɇt��x�^I�
޷H�;�F6�T����;�Aּ�9zUD-}	ޅ���5|x�fU�r\Uj�ӊ�ٹ�gG�m}|�Ў����5�����|�D�=!j����>�"<�_L�yu��v1nM}���W��>��F��7_���*����m6�&v�㮯թ��|���SO��5�7�,��vo.�\]x��n�B�-��5�(O��.d��]eexb�c)w��+ƩL��m���QK^;�W�nT2�|��w���=�����){h�G�{�{|_/w�rް`��kA����ئl>�}����to�9�z�B�v�G� ����F��y8>B�vI�w\���@����+ۊ���U�e� *[A�M*��z�cn�p�e݀�B�
�ܭ�>���U��PNB6�����>��y ����A�2v_t��(wu�c��<Y�؆|���{(5u�#�B�0���v��Dm%��k_֫ݓ���cT�Q����j����MDf��m��z�k䀿p�ǞS�g��ᅿ}���<�WR��≎��e=�j�y��8vG[VZ�AN�O�G�J0?6���9+�8��B��]{6^!�ʺ�vFv���-�8M��2��Sq���k�o8{��C�g:�:���j��.^\T��5�Zۻ�y�wg��)��z�ΰu�[��'��م����5����uz���7;j���=�m�2܎/�T�t-�:�����=C���^g<���0�;T�>��b;��3��/_��ܽ����d6�m(W�tQ!t�Mf�Q]}B��r���b���PO��M�"6�b�#4	:���wSlݝ��ƺ�G<�鐵ٖ݅�տ��Z;5����dR{��:�h��x�G)r+͎z�G\��"^]�Ȼ�'��Y�En�xR/N~����|/WY�]��v�4��{�J�g�sdV��з"p�*~��H]Q�x-���n�S����JΖZ�h-2m.͂h�5+Jo�7�fԂsv6��˸�B�K�D��1qG��Rٝm�`l��UN�i>�,zه��\�{h|��i�����?k�*�������8��ڎ��������9��m���Pe�:��4��1	�%�p�����wj�\T���;�7�:�!�&�mCS�Ѳ'��u�C�ۀ�ws�+rO[���䅫��u�r�ǐd[wWu�'��y����� ��=��/V]��+eJ�=K�=G/��L��JŵK���_K������«qØƻ��^U����q�=���AO��}�V�\t�M�]Iָ��P�f��\eVZ�T��4R[.rt.��{�r������.���T��mtF㥹��L�8��<O1�b��d��c]u���UG��qof1@+C��<j�)��^�C:_N�T�ޭi��q�	�'��CȞ��ZD5*i�'0�ٚ���̛ヽ��H���^�u����و>�+Z��ݐ�v*�r5U	3�<��U����K��1˱3���Me��<�y���v���� y�`\��:���mmd�/r�0Z}��6���t�v"�
�u�q����p�,l���wԬ�i��q�e��vy7Ow���ʑe����o"�������+GK�k6�}���.���p*��VUy��@��5��W����[/u;n����fXS��t�b�㝩<�槆��"���$%â�<�][�`��O�y�oa�bֆkEWH��FK�r�evn�k���ȇڐ�վ���6��"�J��G{�f�+p�C��n��T�2��{��ڹ���Vf>}�Ԃ��6�\쾧3i�/#��*��Q�]��YX���o1�,{��<���k7�l+ސ�9o�uC�����,4mڢ��i�t��.�ҽCZ(��Z�8��k�ޠ��R&���8����ݏS�S����|��=W�z:ջ�U���Ǻ���*����ˮ��K�Q��%�]���9�u����uD[�\t�v��Wy�}NJ=��^QW�7��BsWM���)ދֆ��s%;7���j�� S{^]6G��|�N��r"7e�;#�ok��wRh��C-�#ᕒ��V%�˓����M�0�������]��#��j�Vqr�gZ�}�+9�ʤw.R|�V-�.v�2�*8��B�P��yI�����&s���]���<��WϪ���&�ZZ�B�ٱ�nz9S��ާ�ӱ�{^�1"����6S�p�.���˱t޿���}X�iy_n(��n^b����ꅘ�oK䙪�U�Pn�T%nޚ��'.b-ӫ8���f�������[�Sݙ�����"-X����u�`/���Bh	�u������:�\c���6[���ewoCQ9�j���O�4{;�za�Kbk��.^ש������C佶9ؚ��T|Ks��;�z��z6�M wD���I�IB.���s���� i��w�_=�x�ף�r��y՚�t+:�:9�����}$��^�z��%t���hs�=�/����O���ׅ{�Sw5��f��)�v��26W	pD�;@Gm��>���Ƚ�^yѵ�aח(�����S�3`RX]��#���@�s�pe��z�f/CR3z:��w�{���2V�Kxo]mАu�Zj3��7�VQ8i�,����=O2��ѻ�+�K;8H��P����0G.���!K�^wݷۉ�����g]1�.]2ii�����N2[p���KF��-�'[t�V6�ޮ�0�g+�s�T��yvF>���z���Q�Gf��G�5n�h�����g\S�095(o-*�>��T�{7�ɹ��X���v���Ȧ���y�������`�xq|��*��5�A]��2-������Hȵ���}��U�ֺ?��w����%��=���o-ǕS\'�8U�ĵ���[p.r�A�z�>m��{/vὩ�|-�y�ȵ�K��c���5���eG�H>^��ճ:�9��5����_c×*��^L��\�1�Ӻ)��ڢ�yvU[�d�Z�O��r�M��5)R�*z�oY�
��,���,u�j�.�m:�Rᮽ�����s]��9�8���u�3��ys4����pU�TMA�j��*���:�"��|�^�r���xW-�ɮϩ��7{��x�a\ã�9I`����§���.<2�O9*�+��=ۆޣ-�QX�U��:��V,��V�D|D��i$�:vCD�R�4k�U��gRó��N
��c1I����x�e{յ���jF��P��{9Ll�]���^����ǫ�p�*��8f]型YÄ��5��"�L��(DV���h�u6L��|��V�U�"/1�(�����A���}��C�y<^}M{��GZ�;&.��x�Is���5�Ӗ�#�ە��xH�f�p�h��a_I��}�=��od
�t_n�[p��	�$��������(����!����	ّ9!n�>�۪���JΩ�uF���m�*���ov�ViPe�#��P9O�b^Z�!�چ���u��j��sr��M�\S⋱��	���:�4����(;�`C�۽��zz�ܺp2ު0Sj
��5�'�=����=@MWF�����V�zߧ4ҷ�X�y�HY���5Z6�>Fȟ��
��jp/*է��
q3�β��י׋1�=�wSw+����Krv�.o��f���f�8\T�6��*]���վ�X��LVog��z鰰�R��|��F��w<�V+l�,��
:>��������w9���7�?gf%X-݃FA������Q���$ޙ>����'H��dY�^�:�B�{2Er+����9j���;Yd��,�����J����z�;Q��V@ua�NL�`�؎����n��x����zM��_ ��p�1�1�FE*��׌�7]��4<��Y�(���Kyӯ���}���ǥG�cm�����{�ݭ�g�f����j��&4=^j�'��|0�$��v����dY��>}�`WvS�o,u����J0�@Ή��f�6v�n6�U�4��k��{�3]�/������5�md��C�V��Y$����_0�M%�"�y��Eu�^�#�.i�v�_�%������5x���P���v!&��)=�V�maf��c�sw��&�����v�|��J��-}�����	밻-�ZeGwi��W.H+b���qY�-���9�t c[�K5����xZ^�V�|ֿU�����ۯy�J�����.��P:��Y��:�����7�E�.������o�w�*���2��W����dd�et,�Z�X�BZ�\�8t���"c*�[�bD	m�c��4K3"�Uʻ��cJ��0�'�8s�;�����U6�2�6���.a˛��{x1�2�m�ѷH�`�7dD�6���ޭk�D ؀)�(�}Y/sW�1q֋���r����}�h�B�~���m���쬣�M���ו�.��x��*�����OM,��Δ��1�9a�7��aBGTvל���
���Z�')]��s��q��T�]r��h��8���K���qZ�G˷�m.�7*�k9&^�P�Sg�vVW����w��n����C��q��
wFڠ���[��u�]]��{in?\�XO�B3�UC��kޓ}�^A�{��k��*{teat0Z�\��o�%+|4��=7��Իi�-�����yw���E����{{CC/>��1��Md���6.�s�W7Ԭb��`��j���e��]ˌ���{�"��]F����K����K�ֲ�М�~�:���4�a}i�v����w��WS�#8ջ�{��,<�'��&�[���7������8�E-YK����c[E�v;
Wa*BӃr�u/�c��"�$�:z^��-��������)x�gv���)w`*�E�F�e�TL�X�����9׉^�SM����4K:����GӰ)�ޥ]5����F�՝.1Z���V�/!�xw[�P^&����3�E^���k�J+a�TH�iW*p<�ҵy�L�nͱ�������V]>Z���/V]:����p=VJ����-"�c�y�Vݪ�:��MD��*��tL�fi�mS�")kxw��R:�Y�miqn�v�B��ܷY�\���j䱈(n�Y�Su+U^���j]���p��nr�#]@�.�q����+5���z��+�b��bU�����dD�`� �FH��swЀ�e`�݂��b�A��M d�X4op��&��s,��n�� �Q���rV��7�����׵�M���Z�F*o���ԧFv��L4����ul;�p�}�9��+k�6C}:�t#}c��V=#.]L�3pr���`����r�����^\�	��·,6���ɷ(�v�رmF
��X�{3��K�������!{L���<˸�c�_»l��<�캈��n���n�e��BN����ʙ�gDL&4�����%m3[x�i�/ ��h5|�	x
.���MZCYڞ���������Y�u@�+�e&�f���\���sf���˗XU�ɀlc$�G�+�T�"Mh7�N�3�w��x�Ưvq]H5ݭ �H������ީ����9B�U��$i�Mㇻ��i����1�Gkn㓁c�ɋ���;�gp�(��r=෴	��m��+�[ڡdk��2_m%Sm���-��,Y�Kc���N�R�v������ًh�AΠ��wJ �h�1rΩ��n8^u3��I/����%A�_ٚU�2w29#���Kn�ICpU���
�� e«��4R=��zS���5��e������-{}Y�2�e#��_�cCo�㥵ُuĤ����;� �����d��o;[�N�[!kn�ݰ�.�o{�T�����LXԳ*[WX�\��]��r6N�C˭�����̡k�B���7��ǯ����Ԃ��͚����Uf�_\9M+#r�\k���U�L�&�:Ի���)�\Cw���z�l4������45���5��Va�F:�N���>�®�]��ɉ��:Nc!Б<w����t�v#߂V~�;���K,��3��D����B�^TF?�R/*a���`�E����(x9���#Sר�,�xw>%�
��:u�*j�y��s=l^'�|�3$u��֋�z-2���=L5Ƹ�۹�'\s�5ut��N�uPv�"��6NNj�S.�J�bĢ9���8Wq]�L�0�U�{���u�b��b��y�k��*�����b#*�8�V��k�z����ow\#���'�4����[����A]x�H����#�֨_2#9p��y�N�=��5�8E[��r嗓��È�@f�,'�Ⱦy�֬���e>�8�y�<��ߗ�_�v����J�Y1�5"�PPc"ȸ�m`(b�JX�a���A�b�J�a+���E�TP��V6�VQQjZPZ�bJ�C���jcaZ�嘒c1@"��q�jE*VE��1b ,��G)`e�X(���d�b"H�C�f0W-�,�+"�T��X,�h�dR[e[BĭDu3*;qr��e���jX�1˩��0�h��1
�(�Ȳb��\��U������%�Ȱ�q�36ʬRT�eAf5�h6�0��H��
�e
�K��`-\��2�X���(��a�7l���
�XV`�Z�e�2�+aUR��a�aPSVkU5D�f0�X���k�@�)hT��v��̕AA)5����8�b�X��EʵZ�m�������\�<��{{�:ɽ���Ku�Y����UM蕓�&��Sa]�����]z�b�}Ɔ'3��DSش�:���W�1�~��ymXȻ�Wv��x3��8�r��s��@��G%��/7��Rkyϸ�l˝�Y���t���[�-}���1t[�����1+�)b�|��sg\�vv�v����n����`�9�R;���g�"����)\����^u��D���}�s���>�왇s��=���-[8�4^�.�P�Bi�"���@wA\9�<3�֬ ����E<�5��t[�^�'�v�]A�9�.UOn k��ڼe�l�n���&���m,T$�����\KﱨM�8T'�%�>y�w۾��=K���ڸ*Y��9w�D���Nf�6�v[p�q�ƴ7�eNü�|��@V���}�R��[H��	S��_^M��b|����¼;7*���g����C��s6���yq؀,+�%�m�,k�v�Mu8yy����P,�R�0�77n,sҋ#)�EtU�ةk-��4�!��\e���C>7�)�\J\޳Ga�����F:�"�*9R,4�B�2�H��2�Ye� ���}�
�����W���t�>[am�X����DX#�<ߒ�Fjzc7`���< }T?}��y����_�����M䯙�y+��ft!{j��v�ɵ�پ���z�����^��s�/}V��^�;�zZq�M��t�sREu�@�&V�X��η�ե��������+�a�`/��4N=ޚ���fw�6k{���;��i��������=;������Ǻʖa��❛v\��x�>:��w�ʺ��"�� R<��m0�/գ�׼팎�J�پ�����q�A#���/n@�0�c�P�����w��d�ۊ��Vt���>چ�+���?JE�ep/�����ս��&�<��/�+�,�;�#�l�ٿ�M
���a�%���a���p�{�jd.���f���sU�����g�ȯ�U:#�G���)�"i�i��0�̺���G�ܹ�[ږr�p�܅G6���ȹ%<��������@l���y�#��o<���wx�y��־�I��'���V.s驎��)�s�=a�Q�u�<��k���b��&=��f��,A�+YfX�vU:O�ul����dmvYt�|S�!*t��U*��!F(q���)I�5���aСDpc7kE��ԡ�V�'�p����+D+��y�ي��f5�ڮ�|�[;NA�1�E<������Y���U�(t��:��SD��������M�2ϯޝ�r�ʾ�Z4N��y�ř�=�}�=��=P��+tǯ6���<�|�������S'��<�m�ؼ���N�9��	�Xi��xI����;P��{���Zo�/ǧ��5e�p`��c����{�^��k͑؞9���t<������V�3�4�N����'���K}.)/C�{�r�i¯f��jُ\��������z�#�j��7�o�����r}�������:Zxw xO\�Q���݇�|��cкC��2�W����~>���>�[��^��sN�-��������V��`��z���o�w���%��c��Ƌ�B��>g��y�O��X�7��ƻx�����kT�sD�I�^��ǋ���*y�+�r��X^�Vqʟ���l��c�xr��X��	Ǻ��w#Y~��O��D/+>��P�j:�7@TZ���#j5��j����d�Խw��% yi�Bt������Ie��!��>��dYݠo%��ن���qs+t�W�"av��|�Zޣ���Z��90�'����J��$�%Qvef��q��ۉ�,��^�m:�H���k�X��[Z���ފ���]Z^͙�5C����Z�^v��<�@�K� �_�;kf�2�D��aT�pV����Z
j��Dgv�^�$�LYq^��#�~�ex���uC�e�^�2f���T�����-��NX��+��W�ug2�)\x���u�ݘ~�%���#�9ģ��H���DkʧD��6`�����*�����^F�W-���XoN|T�;��e|��dD���c>��?L���\Ͻ��Ϩ��Vmz�~�Ἥs�i�X{�u�\LO��m�}>�6�ۍUd�o�^7��j<lsV�޶,�j��3�;��G͋�43}O��W������\�k��t��/O����Ls�>3�inyu�nǻc�m�ܜk'7�j23�7 zQ�L�-�3c�o�ݨw�^�q|L��?m�^ꉞʇ�^�]�WT餚����iC��py���!%��	��ߧq���7������V*�^S��}P������3����fTV����|Oi�Pζz̒�zP��J�,�������w����k�������}�^�Jcޯ#q�Tm��nx���⢰ָ�ne6�T-�����n�<>��U�@g�����v��*��o�����m�����M6��_��s|������Q��@�j�U��ς�5�&�Ff
�)��T��kJ{�o4v�hx:���E�L�Y,䳻�����H��/n7V�I��շ�\�V2'Ϝ�����m�GT{������j��/�GkV��mȑ����y�4g}ռ��?d�M��};����a��]1q3��L�'�uHc����sܝ��ka��|�zV��Q�Kj|�nZdy	A\=��n%N�&��������p���yP��{�Ћ�F}5�1����u�����w�����uj��+*Y�z@���`>��`M7p*����x����:���C�<�Y��۸���i�G��q���s�~�qJ��� �������*�Y������l�ݻ�����϶|��i��1��
���}#M}�p�{k�X͘���zƾ�Qy*�׊O���c�N{���|^>��|���;�y��cb��s�!��"�'n_��׀`�;^ǽ��}�F'|D=�T����W��A-܈Ǫ���l��r�
�/&iu^I����+=f���C��"��Jnʊ�=� =7�c")�m��{� L<5�¼7c�p(~F�����p��֟D9�<��� ��*�뚐�z��c�3h�Q��:�Q����n��䭮Y������G{Φ�{΀�9.���v#μK̋����s����������?�?3���Ͻm�}]�u�*]-UfC��;rM�+�OAq-��u�8�*�K��y�Y-kwt�� ��(3�#����(�%f��І6dD�AٽN�+hP��C!����7@�8����@j���T/��EE:�N�\�!�3��3>��A*��ls�>���ފ<n#�W|=�;[�?�Yzs�O��\+����NiKs�����V�âp�,Q���J���5[�ޖvT{��U�mΘ��� ���p�����RYHnNHgn'j;2W/��@�l�=k����p)���^��8��M�4j���i���ZD�������ڇ�����}$xf�� ����$�w�}<�y��̓>o���/R
���C�w��v�=��ѥNQc+�;�ɝ���}3�E[�}�|�LX�DkV�皣�~�Gq���w��PÛ�V���s}&�l�x糕w�>���ѳ<�9�h;�.��>~��������q��ܲ�������E=��ѹ$���-�������>dY�2��U�>���\z��G���~����,�z=ca�^7F�H��w>2���o��#��~ N=��}�¨����������w����k��W��mK4�^k`4/�x�Y�[��צG����T�*"W�a�Z>̍�j���/ԑ?}?S�j�^Tȝ����f`����E��^˂�ZG0�1�L��\��J,�Η���n��
�����K����x��a\*E��>�@���MsA˥Q��},m��N���_p�#��k�V�2v��#)�LV>ἠ���.i=g9�Yg�X{k���g�=膬~�\�����<�#�o�@Of�M
���a�Z;�a��5���{{/'7�޾��	Q{~���ݹ7�<
�z� �=�E|��r<X_>P�1N{N�#�dr��w��|Nᯒ���>�f�s>g�r%� ����s�#g���"þ��y�/!�ѥ~;!a)�t׈�B�FEoN�� ����d<�^Y1�ޡ=,1�u yT�J�}���x��<�m=J�ݰ=x{�u�[����z5΃;,{c�Y,_:�����=7�47�����g��>�Γ���b���=�K¤�w�z��N�y>Ӿ:�J�~;����m�7m�g�|��2��E:��:áv�l�$xܥn�̿k��U�V����� �Q>�ٖ}(h��ι��}6��z1��GzX:W�v�\?i���DW��i�X�֍R�k�R��sT��笻m-��Ib�w>ڞq�VE��Y�{#��K�q��Z�y$v��_�Lg�Gh��|i�@�yY˷�o}���_Lz7���#�q���o�m?���7�c���m�/N���=�0=D
w������K�d�\�܎�
���G�>@��\t!�����K����?{x����U��F�:N�mw��\[f�e4!�Z{"�o��I������x��;��8m�dh�a��-��Kn�*�"TT��je\�.�Q-�k~��0�Q����y؟�M���D�}�>E�L�Q����o��3��ϼk�u�Yף����y���y�ɇ��TϤ�.n*�	��@���p��u<,\t�^��i�]2��Q^��{ѕ�f�a{<2���z+�n�쉨��V�x�ͨh��j{��1r�t����⛿>>~f�Kc�hp��z�-Ue�\ ���`{ӑd]Kv���h�j��@�c��.��A�����=O��r�������w@?O���0y���db�vI��4j��Kp)�j���{�
Ndl�o�a�K���G�s�G>��Edi��p�\�+�8�3ٕ�J����?]�̮��*�p�Et�:0�Zw>�X�Kև��W��)�g'Ӱ�{�pj��*
��^���UE��L�ܮ����wǳ麏m�x��j�����X��VK�|Y���K�����,2>���~�	���?0XU���8v�-lW�����?i�ᢹX�0�^%��>��w�.u8�Eߥ� .��P��9@Ty�(�|��l~`����~b}Pz�|��j5����J��Wvnݧ���[Ϻ�3��e�=[x�X��%��q���)�s�I@���o;5�/B��'��ϕi��3�'vgQǯ�Q�b��.�{uӥ�З�y�0dV*�x�ok��r�m���ی�r��\�%͙�.�������T���4?W����ߍ�#=,5��Tǲ�V.<��r��D-'K������#��OX���Ը��씬���O7ft =��G�3� .���۷C���GǧE�z����%!Ϋރ�O�T7�U���׏abp�#=*8�6�����zx���>�1=��M��x�V�Ks�.{���Y��c0Ζ7&w�YDuH��v� ,S�>W�����uڨ����h��Fg���U7��������ۢ�9�O�t��U�X�����p��uHc��~�i��+~���Oeߴϒ;�ׇ_��1�ْ�'�)�Ĺ���D�X޸w�S7�,/s�N��?r��
6ע}Nޜ�^/�=����Z� �e����r�{=F����iҋU{|x��_��>ʩ�2>��T>R)���o�����3ⶥ��d͟:��霱玺�s�Qz��3ҫ@��2��s��I�������F]:��t|<�FZ�p�ufO)��p�U�zl�7=U#��~+Ar�s6|_Wq.����\����(�F�n�2����n�W����g����j&��אn�����1.i6��r@��e��mr�Lҩ�JQJ$����jg�@�4�Ǐ�D��f��yv�S��%�G���y��vs\�ݘ����ԟCѾ��¡�	�E7ivhȲR��ƛ��,o/�u��W��f��Ķno�LLS����Z;�%�#�|
}WGL��]{Ϻ�w���@����y\.��p.%Pn{>�騿	���մt?ށ0��F�E��{5����D`x=�V�z]�ϋ� /z����s�;o���W��:��"����i5ۼ��z��i�>��q�v*<�9Gc��`R9�UZ=�;@T>�Iuqs^�D��m��~����y�5-��^c}��bj6X�3Q����,̇�s�>���<n=���	e���l̛�_�/߰��Z�|��ū������K���.�'Ei�=��K/����z:^��{j��wPZ�nu>��*�Mo�1�x���Nx��;Q���/�͚�k�7��SmU���߀6���Oe{�~�+���D'��"�������FYUFV�;�WY�@��R<7.��U���m]Z�oN_��F/;�U{Ԃ�<48]�6�F�v��RT�2�]øɝ��l��p�㕽>�Z��;�ٞk���#�/�v߮;��k���(���N���S4��d�ݪ;�~��i��;M���/�p���`ݷ�X�08��B��cgc���lO��gO]2��Z�pB�k:�[9�ov����[���z�M���N�c0S��R��Z�9���n�TE賜6����X�x�ʝ�I|킾�9]��[cK�����A��;}*v�*Ȩ�z&#�5]�tH�zT�2,��%G���R�#��� ۬��j���!�B�$2���+d��)��g_co뜻4��w4��
��7�y˫f�=0��2�5L��io6.��HAq��l�7�;s�N�a<�n��a
�8.�+U�W�J�R���[o�jh\떝��c�+Gf�8ɍ��W<ǟ3�G$�b�E�̜�B���gq�s��J��y��0˃�v�j���*.4�T�6��fܼ��X��r�<R�Wni��>�Hm���Ϣ�*`�� (4,u��]�n��I-�D����oj�e��6�V�N6w5����p�bq��]/�aǛ��2�{�\����I��GW]���
�Jⲥ��(ުK�r�7݄P)5��b�cep�_gn�׊vt���l�it��]}AG�U!�� ��#���O�T��ՅM�֗I�(�m��d��G6:��,���N
7)�	k�ЎM�\2���'_X͈C�3�u�Ƭ1���{oR�0�T��^�u�Lߵ>�V�n^.0W���hn�F[.$��H��+k5A7Zg��1|B�6oT�׭vk���N�"J�L])dM{�;5�ß�U4L}[/�u�u�suw��������ffɊ�q��(tJЧ.�Ӂ�y]E��*�Oh�%���ʕ�s��WМ�X���?[
�=�*�'�@�c�MlrN�p	�P��`6q�'L��K��U�6��z»;Z�*�6�r�{��y�3o����j��b$,Vݒ�:��O?���{��&�""y܊�-7����wN��ac��UMTmvKi�������Ǘ�!Cr��V3�ʶ�;˸����+�:l�En�A}h�_[�n�'�Z pz�蓕�f=�C���mD9��2<ڍ�cm�9@
`�6�	Օ�#��B��8;~c;=Į�9vQ�lZ�Y�����V<�i��m�b3�V�3R2Fm�ʐ�B�ni�y]r\wb�)�:8�c2�U�헽6Yj�hV���K���9�QeEweJ9���7sS�]楊�W5w�jv�,Z6��%G�M"�+&�*rŘ>b9P�!=.n���̮�7q-�o��Wu|2L	�vM8B���(K��2蒓(��=�	3*�R��ʉ'V�.���m��n�67mS�O�6zS�;��_�N�]�N٠��́��*�ֻ惬��WV�7
Y�������ʃ�wMk��!�P�jlt���8�`�\�X��5���%�np���_<4id���[7�t+s/�Ķ�T2�$i�J���kYYl���0N5<E̪_.L���"
��`��DCn�a�I�Am�J��b�ݳ�0֍�r�Q-�7)�pCK��b���FVKE����傦7-�
�`U����XWY�B���J�5����ܮ�&��U.fA���Y�����`m���Z�&Pv�Z��ʅ�Z�UUP��խ#j���w1�1��1f5�h�jji��b����ذ�*�V�jc�m��ĬD(���sl��V�u�R"�5��\��s%�w1%2�v͌q36�-��Z�aTZ�2�,�
�TQb�«#.(;fa[�1��c�ج\EEZ��*�bVm�b;d�؉v�2�Tf�m�;����j
nY*4Q"�Ъ4k�m�J%�e�TX�H؟�޷��.�w�;3W0U�[b�}�V��ҍ+�xj�	���T3�ﴭ��Nb.Ζ��QU�8�@vwkD�RK��y݋1ҿџ�锦.2g��s�㋯i~/Ǹ����^��j�*��dZ=��uj�J��+4o���W?T�"�|�2��Ux>���\z��{��7��ϖB�<��]Ůɕ�r�w;�F�8�dy�z�E��d
�R�]f�
�z�x?9c=Q����t)z4ߒ��u~�׹N:�k��D��UHB�%z�����"5׹�{��g�����Z��D��w��X}��5��5��y��8W��w"߫�p�#L�9��@OfQ��_W��-��aW�C��엻���r�c�l����G�"{����_��[ ;�e�)�9"������x��)�r���H7#�=���6�F��ߠGt���LTz��]��zg���@]�`U��I*�h����Q��A��Uʺ/[�y
�.�\�25��l-G+ӯM�\G��ǜ�I����R��l��^�v]歌�)��I�>����S�ͽ����5�A��i�Wܪ�b��t=p�����f���Y����`�+�j.���w�G.A�g]O�잨�_ѕ�a�m{����ge�3����}�?w����$�Zq>.f"�d�O�V�hֹ��u��~�v����s�P]f��� ���`�
N�(�r	�A5�T�S��z���Owv��yϮ&�Pw�/wjP�$E�-2���4�7�n�v�M�@t����s��S�Q�H��޻.=yH_��@�����{^A~�^��X?1��f�J;��V^��ynv�� {j��?Nx��W��G�v�_����~{G�dz���t�N-��9�d��'���N��n~�%��K�;��<v���p��<W{���I㣾��ւ�/}���t�=O�vی�>��s^*�gzcY	��#����
���F��W��(�l0��P&��~�睖��a2�,ǀ���||%��2���Ϻd*�L���>��^�_z�VF�w�@�]�t�:]��{��a[�f�\�.r*�	���@���n2e�����b㪟�D��=��N\LTM�ֳ#�ܥ�\w�	ׇ(0�P�{�=sp\�dME�����*ԯ[0ѓ��С\H��n�s:��s�ﰺh�O�vF���_C����,�5,�X��2.��@�q�ֆך��?�7ǖW����A���H�/�x�;�:*=��џ9�'�0[:����;qX+3��dr[O���E`,=9�>��r����o�EG�#��]������dR��ŢJ���]��q��y�;#["����ݟm��9�Ľ�b����G�z<j�s���	U�+�nk�u��Α�C���-�G�ΊW��;꾁���4\�<ډ�[cML�4gj�<���i�aU�g�����
yNP�<>0P[uH���<΁��e}�z���O���_��L�K�hJ��	 {5��%hWZ�ǳ6̐*=3�u�MVѸ�s�ݐ%���U���~���e\����|L��O���w�)��.tq�w 7~/�I~ӝJ:�O��a�K��U��9�uxh0�����fy���
ԝб�J>~�=n�?�O��vJ7��fǴ�f�C��k�Q�?H��7>�v���*�=8L�*1;�c~j�|E���<n#ު��g*l�y	(��������0Ë���Ú��uvr�v�}m�-��qP}3qŁ1/������^�{ݷq�G{ީ'��{w�zA�V��M�wyE�]3��O��\d֕q>����On'�*W����I��qF�X_�:�����!N^f����^��aՕLf����;�z�w�MP��S +S�}As_f��a�iy�Ϙj{-��'���}�%�q�zJʨ��WLa:�FL�'��!�����q�q\�|�A��u~�>�^��m��:��Z1�M �!�
sq.p79Q`O�޸w�S)8�όg��C_q3+�������
�{Ջ�Ӱf'sC��j��fgq�Z�,�K:sb��&�ܲ��:�@���&����u'����E>��'-�FmS}��9T_$5�#�Aa�w�y/��p��E���yn''R��Y��Ud���e�m�c�����*���w�+�v}�4���TY�yQ����(��z��u�^���8�犎��}�K����*;�P��.�9�O�q���7���~VԲ�L���H���kҁ*jp�Y�+�l��U�Y�h�l����;O�ُ/]��;���n�ϪauW�#��������GG�b_������*�&W�Å��̍�}<D��3��\����a��$�x�����ȨyU�:�ِEG���,�b|Ȁ�ɔLw����	kgp=Q
{��*��󚘮ܸ��[7��>�g+�Y���r�C����A��@xv"�&)���v��נUg�Ņ��R�Q�Gz'O��)�t׍�}@{�����[��*%W���͆6�͢�d��mNmyrq^�>��.��qZyP�{z���΀�9�y��<�}*i��x.>���W��ʑ��r����9Wy���^J��S���ɨ�Ǫ/����n�}1q�'Y����{>(��V�8}�OoQ[=�+��<��ڕ��D�1���ד���k����*�ǂ��\Gz������6�;�]N��,rB����lf����#&�U��f�7�r�
�Փ��N<�K�����,t�7���K\�,/�_v`�So',�[N�6/n��nrr\�ɘ���YF�
BД�dX��|'r�	���+�':�ǵ����Ͷ����'��D����<��+�X�٭7�@��뼢����G���h��~���ķ���NP�F���F�Mh���]���8�*�ᨌ��w�z��ƹ[�*F���S%fo���f="�{�+�g�|z��q疇�;�i{�Y����L�-Db������q���ίb}gy���#����q���9J��]~�\m�]�gܤ���H)��]��9O�n����ϸn�h	mF�2g�b�'Լy�qu�9�����~�q��b��knYX=R�+1餧oݷ�q�o�MOu�ʫb��-.2e\o+��:���zV����\�fWJ�������\~��S�4�_�_�t}�s$VL�@�W����
��V��:b�19�9���>bR��-9�@�G�~��·�p�4�nl���d�RÑ�}�P�����5s�fuw�)��hz'��g`�)�=@10��쑐嚏\a�� {أ��>��ϯݏ��Q�"���!5W����+�7pc�|��ľ�x�+�Y�_ �ȯ�U:"�·��Nw�ۃ=�Y��Q�H�bw£���p�a��Σ\��@��dkӯYC���<4c5Ⱥ~z���;��֕�J�tf�F������p�ti��v����R�5��	;mle�ѹ�m���,I��b�Sl��HKJ�V����#;�熤]��a�7|/��1q��Gt��4��G�!�]��G��Y���}����_��H���
+�Y���L��V��Sy��N�u��i�[���^T&�^�����C�r\�?y�ؚS���@���5�}���EԤ{"&�=��V�w>&��:�ۖǑ�X�t=qq�*o��߻.%��Z��	�M�l]`#�,��G�|�dOT{�+t�͟i���3Q��
P6��^{U��V{��}U,���2z��!z̡�BO�U�=� j�����L^g���?m�&�u���S�H/;�'=�7��e{�n�������(��ge���}�N'����ﷳ q�7ў�:�gG��Oq���v,u�=[�\$|�TWG���m��k�(��=��qw-E{Aٝ�kK����1q�Bs|g�n9�����|{�����n�3wb���
*֦}��ZV��~6�c�z�n ����U��2��/#�B�3�|����1�-V_C�:,y`���1z��֏��\n}�>0�#�L�K�e�EU�5<�~�����O]	�o��M
״cdNnO�b��J[�v�	1}�Q)��`v�"�-��� r92�{�ܭ��Ʋ]>�p�l��+"�de�R��D!	`oM��d��]`�j�iT9���{Na9g�Նl]�k�z).�RϝM�3��w%�v�Z��o g���gA���Jq\]�d{�=r`=艨��7@U�^.�����<,��܃]����N>J����F����`h��z�~��2���J�2�"�%.��#�s�Q�����/vc����q/֑ȇ�(�9��'E{-��QkL�٣I��o�F�p�)�*;詑'gx��|���~5i+�Z�IQ⸔oޑ��{,������>�3�_��教=��TOxق��U,��}+N��%�C�'ԯ���)�e������m�{�c�q�ٯ /�>̃_G�iQ�D�Ϧ��ex��j��ƹ�������,of�Te/.����������]	��@>��+�<m��U^G�麇���a����5^�P�����%�x>P���>~t�T7���Ĕr�U�����چ���V��-u�.���l���S�>�Gș��l�7�~:���1���:'�j���!%��	����w^��m��ߚ:�?��LV�,z����y\�����������ݸ���ң�=��t�����݇��^���I6���I`�1����5�!�s�*�ɘ��3
�(���Xk�p7t�i�jp�t"�]�{�4��`!�}�,�GgT�5];M�-8D�����Z��{�ceE6|�e�P�+��>F*��+�^5u�H�Lt/+v�e�8;'@:<~ /�o=l�=�EeixX�;�o��zX����_���{޿27�>�Mm�k۫�<��Tgq�{��3�=���)L�k�����;�z�wR=���d`�ѐ��3�nVl�㾵\:�����m�0��T�tq��X���ɝf�&||��Y��ߞ����S"���V���N��Q���׳c~��A=�4�I����p޸}��s/�f�W��3�G�t��G<�w]{No�x���V���e��z��q��Ѹ���Gna�����v�ў>�=�\
���CE}��qΒ7�O�G�}����D�˖]�L��Bn�9���PYw��}���eT���x
��c��#e�Wա��lÏ ����Hmߡ֥���Q"馏�рqҷ�#����򳃪4pu���T���><��Y�׋:�Z�	��=`z<j��ޛ�u�/�v\/~�φ��r�B��#qn"���� ���@�<�`;K�sfi>Ѹ�)S����V�G�)��޾�F{2�y^��r�5=�2�W�14����ToD�~~�,*آ2�F�����&�&�E�XX�|�'/���:�3*�h4���6�m89˾\:�8�A4�df���Э)F@����$Q�I�a뙲��8�}C�%5j�E���!�r���VkNwZ�/���Ӕɽ���1�i�b�3�)� {�� 9��`W��7@#෠͆;��Q�����������-�5~#=�]'GiTz8�5��C��sf��@y�l{�g(
�<�%��lw�R�����fs�h�p�&�����'Q�,i���W,ˇ���}1�q'�}�U1����r(<[�|�������Y���}�'�����>����\�j6�	_�<3�}�:���}�	֭o2�l+ܡ�*}U���W����n���"�^��[�/6kM�7�,�| qHV]n�RYz�3W�+���	��Z.<�Wq��:�*�᯲��秨�Q�2v�����]�w��J�+�<�uHCoڬ
�X�|z���^wHh��i�.�{"}Z4�����=��k�n�Z�P%�z0ϙ�����e������#�/�v�~��6���ǲu��
p�K�10 ȴ}~'�K�{1	��U`L_��ד+�3��ȎN�M�;������}��U��b�lf�5qMi���tVU�������x�Kt쪰&"��>E���Cת���
׫�67/�}}@�ð=v�~˕c/���5k�7�i(+12�.��z���2Ӂ�r�]6
��cA��]�on�ZQ����M�M���}}�t��Cݦ�ү�g�<f�q�O����=�3�|�G�T=[�,����PY_A�f�]M�Y��5u]wn�����N�٬�q�2�o��;#�@{�U"�e�E�^sY,*�����n�{�.�d��&�={����;���~�ck��f���*۪��D�RÑ�}��8�|'b�.�v��FM�7����Β9�H���_�܁q�7�L�9����&~�n�o߱�Q���^�[Z���q�)܁0�]��5���{H�=Z w�DK��D_�5�ޫ�8�:�­�v��P�{����D�N{N�l�%�K£����s�8Ϥ�K�_��`����U��yyD�Y7��#�*��5,f�:#�+L��\�g�e���X�w�m�_?z�)f[��w�Q��#�Ev�ڥ&|�v�=��zO��Ծ+&���ѓ��k\�3Q�ǫ��VK��
b�[�*��nyN[��c��OK��r�^@J�~��=�=Q�L;ͯq����ϮB��fS��]x��_&�R���=��X���O�Ұ��{�b���J�2x�D�3�������YLu�%گWm+I��$#=\|��龤 YN��^���`�v�и��5�������b!���;�Զ� X|��N�1�͕�j�M�%����%�N��m�{:����N�����2��M���)Z_$�~����B��tz�nE��GvΰN+w������*_����L���uշ�D��U`˴�V�u��b�W��gP��kB+c$
I����.�,�̈���g�S3U�ť���]�>Ǐ��j��c��z7��Z��}E+��.�<�
Ϳ��%m�<ќ��V,Ӥ�ϵM��\ޠ��%�]۽e�ai
�P�J��
�l��
Xja�{���[��>��%+�+ַ^�ڱ�\V�u�_/�vP%��"v������K�|�h?K4 x�8�voc ��X��9�r�9$��b�zK�*oTשŵ(*�A�����vv���^I˔&{��Q�d�$�-���n��d��m��WD���go��0k�&��K������T������xo�	h�m[�71�7�lt|���8uő^���8���G� xs>	T�H�b^�mBP(0�Ge�ڝK���Y$6��?�I#�۷��tB���-6��])'��&����4�ww��9�Ӧ�~1�uu3jg�"���q��6�ݗ8)̓�Ͳ���)�ݺ��is&:2\��ޤ�]&_"�C��n��c�[NH���w��ep�=��$��f����:b4�ݷ-^�ɂ�T)�l�9�=XY�(���_DVd��>��]�R�.NQզoL� ��Edٗ���<u���[�VVM
Wb+��i���i��37)W	raJ-l�mJ&�}G���x�rļ�j�Σ����)�m�s���t:���2�k�K��$5��I�ɫ+9�6l �^�n�r�p���f]�6��U���p��MF[yS�Pr��Yfm�|4s#v
��N�;WZ˾�6C������AV�2�'qn����q��R���&7�f��[��eA���h�k�}���7��#�gw:�0cn�\���v�^�Q���=����\�e�9-˔�����Ν(�ys땝��@7����E�:�;G�iC�G6��nrԜ��9��D�Ӛ�aP8t�s]�B��^���XXw^n���M>�w�l+U��x�|��d��ж�ܫ���U�Km9>�ti�h�dY-�f_�e<ȹ0�.Z���
�=֦\ё[z�|��`�qru�սV6e�u��s}g-��1�.o�ZK^,�f�Ս���;�VgMU�:D>ͪ�(\�Kkc�T��Z��}(�dU�\�syiY���	�Ynn�b`�447�we:ۂ��0:����7������[bV���U*�A���ØśUx�:�I��b�6�[ͪ��E����1��L�k4wIO�(��̀I��9r����d�.v���I�v.�QCh��-�A�����\�DU1)JQ]�\&&��Z�m����2��f:��"e�,m��j*��
�lZ6�TpQ,��Ȫ.ی
��PR����1��f-�Ҕ��C�G
��Ea��ves����meq�r��堡�\JșF�PF�
�b&&�p�ZDJʅKeQK6��\�УS�V壗32�Z(VW����j,��-��J���s�Ȭ�kB���-D�u�3�
����Y�*cZ�ibؒ��W,�-iX����D���J�R��P�R�����]ff�b�U��+iQŬJU)B�ۓ*��G5.V֍jbIv�)�FV���31.9��[(�6�QB�m�#�#A���0̾v=����|��p@0�Vw�9��L��p�M���V��vowm��3�F�<p��������|��\�{����C�\u�KW7��7Ǉ�f�s�)v��^�B��MTm�.�d�������G�\��y핻�-�D�փ�c0Η�d��b��No��m�?g������;��
��8�5���m����_y}.�=�񷳤�r^ւ�������c	�{&|��B�3�|�"�*��{�^oz���.9�޳�����vyQ�~rN2��*�	����ҙ�X^P`�N�j��5���R�����d�z3}�=�O��WH1�aw�H�J���>���M���W�$�S�.GWTo��V�6}i���Bt��|'�v��������U�Y{�!��>��>�����L"�^�[w�Z�{-ߨo�6�-�6��Q}��RE��:�88Ҫ��QhvX]Ef*���b��f�D@�9���^@,-9�/Ư���u5���&��n#ޑ�� A�1�t�̕9۱�eo���@�w�[7����"f������V�����h{>�R�Lz�ϓ�&��ye���k]3�:���5�ɯQ��Q-ɺ���W����h�k��>︋u�����P�H-HA�L۩���E�N���\�-���A�n��B�L�P��4�*���-͚2N떦E���V���+F�.�q�u�Ɋ�j��p�a�&z�0�{`��Z��.�J(>�H��0۹RV����a}C&A��է�j�@ާ�J(�;ui�j�-e8��������#��;txu@y�h���=�M�=�Zد��f6�����?t��ҽ��uh�Q�b��j�|n������1%�Ux.�����)22�7�\��Fyu.<=Q���/�>j�|E���<o�w��{E�Y����q=ppߊ���u�������>�sᗎ�;�'kf����!����d39��G��{�n)����#���'{!�y�y��sI%��:��N�y5�\d�V�dg���6�<�_,�g���"R�9�g�L˾p��p�6}�7����^��oEw�}#��/rkK3�7�wR=��zw�F; e\����>����=����b�B���>�m�1=�M����=��]1dγX�ax���f�.���Z�{B�}�!�n��#�����~���e��r���H�=�s�5D�i�5ݸ�?�������M���e#y3�&y��Q�.��c�'�=���
S��eK/#ޠ)����L]�W�&�z=ϔ�|lȠ'��{�'/L���;�P��.�9��>=�7�����~jp�`�ߡ��v��f��&�D�ع(ꇳMՑ.e��0c��\��[x�F��Dlw����б^v�}�5�yNo�]ʃɢ����3	hU����Nu����8��<�S����0Έ���:�30�_o`�����/��=��١#�L����Y]u�+SY6n��wo&s��P��y�ڦЕ.���G���
�:�<��l��}ï��{��"������cO�on=���c�A��۪��ex�8\�͟W�����1����ۿg�֕�^�x{��H���H�#=�T<�7<b|͘(=��D�����9��-C�sj����y{g�#"���j�K��R����˂��a7���n&@|j/�bc���7�ށ���~^���۞�>�u�0��rb��׊��ݐ]h_����P��p��T��س�?g�y���B�U�kK��7^��b����/ސ'J�2ǽ�f�C-׍c�/+��v�{������M3~����;�=,i���Ǫ9fd>s'��t�^��b��\�wvȝ��#�y{���6m����9������u��^N��z��3[L	���뭟�o�A���|�]%��׭�����W��1^�"��I�v�v��O���6kM��@�^Om���[sO1�U�oĸǬS\@����G�p��e�P��i�碻�}>��VET<9;0�4�Q<���]�+�*j�$�t�g-B >&`{F���[
�J�7l�%s�$���s�E�u+�p����+z@��U�wS�8t�讎�ݎ�rAa0�H����7�5�2��NgI`�\e�|���wj_5���y>��/��]2��?Lݴ7����g���~���b�i��%���RT�̽�z�}���lW�r5׬w�N���;�q��L�L�����9��o��׵���Ԣ��^�z�#�ֶs�)���v4]SpS}+ҭ.��L�zr9�|S�q؏�׏�U���2FV�O����}�QG��H�%H�����DT\�.2e^��|G���Y�Tr*����9�Mz��eK1��]΀}�U"�e���]d��P:�c+���J�l�_��ﳛ�1�E4V���j��g�����nn ���U!
�^��{w���Q�P�om,m��8��Mw��ޫ���q/ԑ�~�@��X+����~�x�<�#�l�ٵ�C%�뽢�u���<^�Ä�wrǼiwT;�__�|nx���썺�O*�;lL��7�9��q�9!�p/к���=�s��;� ��7�£���=3�>��J�G]Oiq���yFc.t���>���EO����xnzH�\�2*5���/~�b�>�����Q��w�b�<���ČX��a�V�n������B��%ҕ�Jճ�����u�0iv��
�m���魹�yy*�u9�����[�6�47��۰�z���k)KX�NImѰ�jiD-d��J���苚2�j<�e�wPec�lu��t��}K�,ZG���ǖ��Վ(����[�w#�1IG /�]_y�zJ�R|���Cܝ��'äֹ�f�i�K!z��1�n�w���-��軋�|���3� ���	Xo�T�=1����0����U�]��9�w�C%��$�] }�ϣ) '�ձ��T����2z�����^�HyxߦO_N�<3)B����|O�c�������a���\א�[�3��`�Օ����Z/�h��ԯ���ds�#��d���d�\�i`o�㏠mFs�)c����z�#y⸣.K�_�`5~��Я/3����=�%�h*e�،���2g}1q�Bsqd{n9�<����R5�s6�.*ب0�\��'���͟>�p�jJ%�k����
-�|%ZY�-/�}z�����S�;D��?>Yu��cѫ�����^�q�\nC�����D�%�EK��������ҙjLnR3�f���G�������.:��F}�>Gn3޿��b��ת=�=3�.x�&��Y��뮒}�Gܫُ�W������mG��l��]$r	���P*��ᐧh��#L��e_IE���^~��+v�-�w0�'��4��Q���ta�C6�+�.�(,��Նv�v"T�����C�ݴ0�9�v�$��|��Ȑ���J���N�e�7vP�;�Yѓ�Wj��rO���D���l�c���u\�ZA�I��}X999�G6��=F����W�R�#�_F�4j"����l�>�G����f{.����:��	���=QO4]q�O,3����S 3�>�XZs>�~5}�����#�9ģ����:s�{c"�O|��7��+�eS�p|ȁ����?S��џJӰ���hz3�wA�~�ܾ�~��1�>�^�؟O �<��e\���\�C���14�mg�wl�9'��Q	%���I,�p�|�����^�C�9.t\G��	5~���#�7P�'p�u��i����8�%�«�����]\v�.	𦪧����wc�v#ӔC�(��W��_MG=�����OZ���b����P�6��/���j�Cy��5U>#},=�Uh�3F|2�y�,8Z�׹�R�糣��U��<.��j2v�oK��0v�l{a��/|�r��v�mz��,�ЖWo����M��We9,_d֕��p�k������ڈ��nz`��T�S�}4w�~5�H�7<�z�7�yb���T���]�"'�0�Ȫc*2kK3�:��oR����J�Xߗe1*���c6s�`�&���/o��+���F�����nXWC�^M�"�rˏGj�,��y�ǯ�k�ñ��
��sn���32�'��j[k��mqz�{���!}�1V�f!ѝxa�[����U��F�wE���k�1�$�9��(z���1OO��ë�y���۔b�{��'�0��Q�5��^���]Ī��rk�w���,�~�>�3����7_��^�|w�_�í�Z1�M �D�*%��K�s��c���;���z4B]q���7�>ǝ�5�״���^)o��Gv���e��Q����U���������V��	�}���NEk޸�ϓ���A�=�h9H�=���s\��Z�v�S�圪�Ǯ�+�/�J���<�*����W,yia(��?Sf)^���g�=��BR�9�Br4ײ�����4�l�0P{UHU2�V����;=�L�o����ަ�)��P¥"���Qsq�U�{.�K���ȿ��U"bb�W���k�v(�ʩ��o���q�f��tz�Oq�/���9^g�|��dP�7�TSG�d���G <"�O���䴕�:�z<�)Q���=�c�w9x_�B���K�'mR *��,
����!)#���<���Į�m?��g��sO���=��o�/MG+�T�����r]Vp�߫���R~���GLͥ.�fP6ߧ�X�;^�ޕ���*)Y�o��r���/6�,�Y7���B�E=ל]p]x{� Zs,.r#�jh]��mMkf��N�j強w��o=X�6�dȏn5��Y����]����s? ���'ô��/���ֳ�O��ic��27U>�y���7o}�W���6=H�!��~Tl׿Ie���?�{'�����>������f����ϓ3R';��귵�-�Y����k��g���V*߶�L_�@Oi�T�v�jd���p����y*go���b�w�;H
�V��W���;adue�h~ݭ�Oi��H}Ul�Q����9)�^��v���BU�;�{�����X�}�Z�H+��C�{����g�g��B�,�Zʅ���z}����o�3���>�����co����~����1�^���^�N���\nw��U�p~��Y�lx�\�_z��d�s�>^�fC_qu�8�/�"ߴ���8����+�o�mS�}
�\nG�����uLܷ@>Ȫ�&*yW>E�%tj�ܶ�Y��5x��/5��h��^�;����\��,�p\���ʩS-�*-J�u|�_��1�]�bZ;� �_�z�x\{�v�}މ\{"7��W�=g���P��2�'�=�����GW^�_�*a�*�O���;_�ݬ�J�yK��&ﷇ�Ah�ee��(���x!�.�AI�۰�U���̫9�&�%U�І�WJT�^d����ǝW�a��.v�2Dq��ke�L�8� �����ƝP���F�97ROR��#�mV��I�+��L?�'��26�ʮ���R*��/"7������џ}��wdyK���<��#{6{g���[>�4*u<8O�e�&�v��ܾ�x�+�Y���{,�c���"�䋬���=�=u=�=P��fMQ��@/�t���j^�*��l�J�����ׯ�{�U]�/ѯ,
���I
@�=st�_��#�r�ȭs�=� ���\3}��Y�}�kv�dn�C��=���%C�r};��w^������R����a���j/<���~8��Vl�n=�W[b���p�E�\�-�Yy� �ל�~�g.A@g~�O�����en�v�T��D�۟r�S�
��Wg��F� JV��!�����O_��U	����!'�\z����9�;&���osR9��>��P�#6�MƗ����
�����FGz���ʑO�և�y�]�3��^���`��a�RU,�V�?��](����8=B^sg)��Y�mj �x*Q���w�zev�+ܶ��;O}>��VES_d֗q�;鋍r�{7����wi{ʆ��[�� #r��j��pŚ1s�U쮧���e/Ns��WmO��:+p�[�Fg=��Js���t�r.�_9tp��/^�`Ÿ����&���MK>��>�;��S�z�c;�:] �3]��eDQ�Ip��}��Oi�
Tg�b�*��I����m��u�ӄc��d����ӟ~Z�=8KeD��g�V��crgY���./�_��"&�7�Vj�� ���&X�9�;���U��s�۟Y��*��s����2��(S�W�P>�\�z�ុ>����GS����^���D��g�^:�A������z+�n��_�_���H�jF�EE��V�˿�f~��T���ks�p��E�g �ׇv���_��=�(�]v,�LGc��1>�{��6���n|rx�EdJv����d��ﺡ�K��r������9#E��o�\�sY^�=��O�L��Dg6*dL>������U�T;�mg����@�I�\��v��T��?j'��.sJ��tD�����}�  �b�L���>��rc2&�<՟Wv����Q�zz�ǽ9O�'� /z�y5� \����y�^&)��;<9�^��$�b����Y�Ԇ�F_���ᷮ���>=��z�t���<��� ����⪽�dM�=~>}�7ƣ�nU��4�ٌ��rk�+K����Er�L_�ꏍ��<����9�^bJ9��#ˊ5�����2����|�s��"QC�b7�'
a+9}���,嫶�x�	k��n��NG��dԸNo&#��bu���WY@d���$�9&�������t��*�4m�*�U�����I�:�a�wq]!J`5�_tG�F�Q������sh�w�z�F�J�k�t��������a�-��{Em�)��REO�6�|�v�6+1�3�L�Gm�m�#��+��ڲ�����j��q�Ǻ����>����ɏSX3AJ;�2J�t-�����2��o��j�7!��Ɩ[wY��1T����t��"&�Ԩ�#; J����x��qUt�+�&�c[�� ���g;��w��S��p�ZO`e���A�ٻ�K�H �����Gm%�ܥ��W>�3�	w�];ٹ��q�-�֭��].�-��r����i�F�j[d�Etx�N���������v��Yv�sJ�^���L`��528!��W��,�1�7�E�n>��]�j�ޤ�E�Mc�j������p"�ڵ��i��i�|Ga��mnO�--��u�f�8��W�Ky�Eu-
�����G��'��H�V%��]A�u�ʃS�ŷW�6p�٧�"�Qǃ�u�v�|շ�`ޤ��n�B>ū�L�Rmf�<$�ԥ�PZrv�}k��_f�mN���c�H<��[��m�;�й�P�3���~G�ۃm�lӑ��d]�<��6ƽ	í:b�T��$���:����*�u���� Wj����T���ؗU�#Xj��|����vK�Ui�n�1�"���;�Rt�gWY�c�,%R��t���,��9rN���,N��6��.�Z����M����`�8.|�EN��+j�-ֽ����;\��:�o��RͩK�-\��Һ�+y���OźB
�g�O;Vik�d[�uEǘ�à����ݚo�+i�%t�Q�����O��J ���|���+�iZ{��v���7��nq@R�#C'��s]����r��9��z�q8y�^^C�gi�-���+S��ή����&��?#�bS�dGa��)䘅�;�u��`/JZh�9�Zq�,%h��L�;4DF��Wt�U�W@Y�|�n5�z��\���ܓk4)e�28-��J���J��#��Aǔj	/����o��xM�	�<�Ԙ����V����GEoo���e�Ft�.��-�o�J�H?dn��U��y7fּ�ղ]u䂹a�'9����Da��@��Rls�2D%�?�+ �'M$}�}y˨�Aˑ!{h���N:.9ۻ���$L�[q��u�ե[�.�e>v��
>,��1�4z��x,�pv�bZ��kѱX�$�qX���}���s���u��J-d7ٹrn*3�l�v!j�d �>��䒹�be�ݢ���s�����ΐ�� Œ�f�vR���I��x��ǁC�R�I*�ov`�>��q-���=�=�fpIi-^c����l��JF��I��;�,CO��p��\�-h�K�1�R5�,�1U�"�)r�85Z�_2����pĸ�1�3��%�(�,��*5�]��F�APTUe(*�er£��Kb���,A2ت����)�����m
�Z�LL7m�\@��Y]V�Q��Z1f�(.R�,uܱf%2��+�m��e�Z�����ܮ��Ԣ�m�m1*���R���(�h�m���E�
�qm�wnT[mYlܢ���SY��+-����Z0mYb�,[J�b�F�h��"*�P����̸b����Թ�f�pJ��ƍ�U� �,���eTUX�[r�7-¢"�6�e-�r�f�
��DԦ���Zʔ��)M�������R��1���TL�V)-�ʑ�Q����L�11��EAFel�N��xn�|�u���#�7I�,�b wkB�s�D-ڐ�]�.♖��K��c��BJ ��&�%����{�T��BG�ݝ�B���co�)e?���5��=��O�xo��O���3����L]��>�bI�.���EmV�ǣ7�ɜI��{���+������^���s[���c<��Y���pUU��G��v��߲,3�D��+��JX�.U�����鿵��M�`h�k"5�t�u�ޭ��D?;z��{�Ѿj�n{�Q�x'��O�aK*��3�����Yj6.�7^�k�~ūV!�綤v�i ���~��e!��{nQ�{��9��%LǬ�a"L��k#7v��9o��bo�=�>F�g�<��w?W���μ�l[���������{�iNS+x]��8ic[���D�p����q�,/�yP�8���������_��իc�l0�L��������|�\R����Ϩ
��t�}9����ϓ���A�|��&��I�}'�q��c�t��=^QYw�亽h��R������f�� �DUH��]0*.X�>��Q}Z�t����/�b��Ӫ���Y��_��6s;�0�{-�<��3혖͘(=��
�ex�8\��%N����f�鳟XԶm���R�����������s���՚���.���|GB`�Gj.���7��k���ג}Y5<�e������s�� �Ӳ�N��$Σ�S2�~�FןC�-<�\���"ַŉ��1��y5 �uΧX����R�6^P���R�����f��=�L��G�Qsy���=�<f�_�O���ۊ�L�c|�ޜ���rD����v��3�Xt���_������W�Y���ِE<�M��T�SF:|gѓ]c�dd���E`1+g(�H���0��/
𿟕_��:��΀{����U�V}�C`Ou�8/ܺ�� zt=����f���Vɭ/O��G��	��5�7�:�׻eD�u��K)Mt{6���\���Ys^�}7>q�Z�mxN�4��icܮ�j6Fr�}�3[u�|�R��}eL.蓧��ᓖn#ߤ������T�~y;��tN�\�|�k����7۷���BV��R�c�zs��}^=7�{��U��s�/� '�ߪJ���+A��&.���L�M����'\}�R��6������*�����{�5�����,�8����l���`]t����f.c=�b��q�@�}R<7���s��U�����/���Hw#�ʸ�:�Ez'g�G�jcs����h��ȣᘪ���3����	���co�~�i������R:c�=�0=;S�:��5�����ѨS��|'+�;-C��W�����{SZ+s v�V�r������K�s{���yފ�Z�m���"��F��Y���s���gor�.W>�������Y�t���y����ܼ9�ڔʑĹ��)��^�ӻԩ��U���Փ,��P���L�}�y2����>^���4qu�2�oh/\e�y׻��u۳�i��ϑ��*����嗑��-�fh��DY�,vL��E���S2��4�R��1��-��o���sޟq�u~���,�f��f�>t쪑u�L�@���m,�k�{�#�j;�g+�^��w��=�L�Oi�����_��Ǘ�bZ6K��F�-���W�^B��{���;g��y�P�]w._�#��H�o�~�r=��g{���?=�К
rǃ���H	l�2�vT�݃ǡ$�}-_��!�^��N�C��'e��fh>��<�@�S2a"~A*_%DO����wND��1�~W~>9^qw��1������V�r�{�R}=�����s�!DJ�=�7Lm�z����Fƽ�ρc.;�9^���]��)=�?_�&3��P���������r}%����M�=��oC����:K�_��f׉����6��q>�f��yz�K�z���t'��<����o�@J��>G{��t5�/*�QǓ��0ޔ%������I/8-$m��a���<]���Ք�"�ѣF�%�e�Q�x��cǙ|����~T��u��e>�}��4�p����c;pj�ίa���,r�m_)+x�����"�v�ԜzT�����v�;&D�j��N�u
�͝��&�%ѭ�˩�����7���ki�%+��cUS�/{��Y�P�O��_{����t̯���qε�У*��=��Ï���}��q��-����#";���q�ݺ���i�׽n��O����ihv�wΨ��q;,e���
�'����7��}69�
�g��t�Uh�W��d�l�,y�'�Ȼ'���_��=m�[����ZY�T�<�yM*�8�]M3�6�� �xȫ��koB�����=��wO�j�\w��{:Kg%�h*f���,,��o^m�̨�9���/_x�xV�x�d:�OW�|<ϸ㈿W�nb��ϟ����!Tʓ����6�<�Mv�^��3y0��ґ����O��a}��z7�}�TG�^p��2 �.��������e���u�r5���TE%@T[�ˬ�j5�v���6�x%ӣC���*]���8��n2n�o���fOzh��8��M�,t�"�[���-nmCF���~��~��3�:��;���d�u	�u���n�ǕS��4���3�H���,-9�/�������Uٽ�;�3y�7\4��ܥC]� ���dk�x�4vҷ�B=h�F]7�;A�J�0��1���w�Jk���{�qA2�&c�2�b�J5u�[(�c������Z6_Z��_g(�+F\!V��E.���v;V��tCf�uB��	-��2��knh�g�9��Qϟ�Edm�
��N���l�A��"f"������ZvkT+s]a�͇����Lw��29��0��s>�N���0�}$*%��7P����1��vCr����[o��U-�;��{ʬ���W���{d��{�7py獠fg��ǵBD*ܬ�s=V��/F߾U�a^*�:�WGW���X-�n�||��s"�|�(��uLɗ>�sY��?'��'�/�C�	��ғ����+�~-�׆�US�.#}L3z��>���5��=J�o�^���p�$���Zn'e��NQ�\o�,{�x071g�=�X�)�s��Vwf���'O�Օ~����Oi�l�1��MiW�O�i��#}$ڗ�N�%�w{
Zc�;���W����{ԑ���qW��x'��O�aՑT�Td֖+s s����o�w,'�����}��>�t����-�� �گ�}�������Dr��<B[+����*:� R�I����ᛪ����p���72�yR��9���#�����~�st�~�H.�<�Nf\
�&��i7Ķ/�/Wu엙�H"c�sa�}$�ӈ������vg-���WB�W� *w�����͔=�t�t��������ތ�k7o/!��k3�)��ou�Ժ���]έ��鴫�i�ވ��d\	ռ�1�hZ.�R�}}��'R�j���ެ��T�65Ϣj,	�w��f�ɖ�r{q=.����x�Ϸ۞Q^�E�{��3���+ݘ�ѫ�P�}���� ��@j]~���S-l�h��a�.�3)FǴM����ied���W��O���VԲ�L��rު�u�W,yiaF�um�%�ٿl�gg��h�}�{��؂�_3��0ϯ�쇰6\��&%�fn�B%x�9��s�4{�-oV���=�B��pw.����i9���{2��S���̯��Nt���>���u�+��Ԯ�vLzm-8K{;�����q/���9^�N �wL{�s7�^W�G��������_�<k+Ò�Ԑ���Ӵp{�u@�xyxO�?*���݅ր��l���;��0���xw�ݩ ����3c�sd�^���K��7�/���L:k�6f������.�%�Χ��y�`^���)��\�L�r&��^Nz�g�/a(���~�ݰ��ShB��qx�yoEH��s钦=�qG���Z=��M�~%��~������u��Z=�D���V[T?���'��3E���#��g%���:whZ�~ߔ�|��ԛ��5��'��%E�n�F.��.�����9��t641k�)\L��3O3E^4��P:���f�+y�u`���-�pV��ӳ/vh�i5�f�F�Bs�]|�V��fjc'���,%��o0��c?U-�%��l1�w��7�˛�vՊ����"����هc4__���"����|:=L��٭7�W���Ul�|���2<��{��(w��5���WqwU�V���&�J�vy�dRvg�BOջM��k�}����5���������/R��=��=���Owtb˼�/���h��K�T�Qc*1]øɝ���}3}2���{
��/�v���3y��-[}�2q{j��|ֻ��jQY��]ˬ�U`_z��L�1�Ҽu��@�)�ӹ��|����}�|�G~�z���ۆ��+=�3q� �f�Ϫygȱ���{��p��%W�����Wu��h�q��9�������q�¨�z❛>T�*{��2�:w2�gv�b�r�1�dv���6��txr����
Ӫ7����#� ���=791q�e��b]QL��T�s�R�����'��3�j�ZE���l��y�E}~�r5��=��)s]���}83��;��Ā��qJhT��9KGw��uC�}~�ϣӕ����g1��soxD����(/�y���S��uʛ&�wa�~�M^�^�<Q������g�"���u�.���[�oT�Rޗ���Mk+N�o[�Y��/��������Y�nB�!�oa�{�B��d�Ŗu�"�c��"�k��;/jt�V���v��e�Bɯ �vY�����. ���j��{N@~9�A/F%�q��8I�Q���!�'خ�w��疔M�>�)T{�`T[���r��d�1���=_E��"�����$.�k�)��{ڒ�v�>�Q��S���~t<�"\�Xw@�����S�{"n���V�~�;$�}�ą�/�
���kiIU��nϲ=�F���zht�VA����z���]�^Fv��,�n��S�az3iq�s��� d%~��g�-�2z��!z̡9��Y�>u�y$��<<t�����f:����l��/ǧ���,v����x�wؤN3��p��LӇS=���]��>�I���N�.�*}��gC==�@ڌ�`e��T�ذ���~�r��jnw����U��������������9�eSQ�Z]���b�\��`�^�Us8����~�)�@�yS�\v"Σ^���{V�E�ʒ�s����>��/��~�y�3R7������g�)�ϳ�A�>����߫�nb����Qn%�2�q���*E7�<:�0c�?C�7ГB������S&J"+��e�T��tB�<��1���oFCت���no!�s���;P�he���0;����S���h��,d�}���ˆ����s�Cn�
T���%�>8��s�����}�y��}}>F�e���xX��X3}�<�^J��K��U�<|��O}c��qE�s2�������g]�Q5~�z���J�u�Pѫ��;E�E�>����K~^�,W,�v��+sm�E�'���2<���P��2.�[��}����K��{��@2ƺ����9���W{~�'�Z� 4l�l��S"b�q��ә��x��<����^Uוܧ�����E{��i���9ģ��H����Y*�/�'̈<�Du9�
Ŝ�B��a�}ۏi)[U��ߠZ���lʯL_����O�@W�fA����Q�^`�:jGn��'8��c����۷��b����{���j�ǳ����VK���s��{�"%΁���� ��<�bz9=��<<��_�]�(?Շj5��u�j4�O���Er�L\sWs��@�(.�?����[ц�G�}#U�����g�z�!���M�x�'��0z���~-�׆��T����ͬﶫE�o���P���:���h�y	(�Ǫ�ZN�/~��vrzw�/Ǥ�GћƊ�d�g^��.�z���;������o=c�n^�����X��f�$	�u�4�m#���
+��X܋(`�G��<�M��v�=�\���5tfr�y�6 xÀ+'�����1cǕl��c����[v�]@�S������G�9��ڞ�F�5Mh�����=�Q/ʧ��$���؝�2�*�+�2|+M��;��[�WY��Ԗ��;�i�6�� T,���ޞ���۞1~z+��g}T�t����L���3��c�_{��S>�{�}�G�c��b�a�W��W���V��E6TKI��4r�/NN�{��b��{�UF��T�Y9�d�sr�$�^��ϼw>�W�_ʲ��y��'D?}Q�áe^^����W���N�"j,	���ø�([,/��G^Ӿ+Ǻ�5���{m_�2�s��z�5��W2��=���LӑF�����g���!�q]�z2�l:&�p���� �w3D�}x�MK�~��f��:�ET���L,yR��:�߯�N��Kܴw8C�/�oW~���AN��#���O���f%� py2B�����6fո�tb�������s6XU}\ħkō���gӟl�Y�"}t��g�O����}�!5d^��w�N8��LMn�ӐKGwØ��,\J�F��0y��;�q#�@B��!	'��BG��!I!	'� �!$��BO��B�BO��B����� !I?�!	'�BK �!$�B�PBO�����B�i$ ����� �!$�pBO �$��b��L���u�f=� � ���{ϻ ����|� �)� �P ��  @� ��H��U	"��JUz �(�l��T(j�*���EJ T��UT�)�R�I$�os�f�0�x������E	�0�mRZ�Qh� � #�"Q�NxP�@]��UB�T�� (v;�J�WFgs��
�M �7RUPU	
�(����!%Uk";AN��ʷ&@�'A�q����Ю��t4�v]��C��� ,��"���E�E��\�Pe-ak�2�Н���w1�5T6u�Uw,%�n4J��H�h�l
�Xhm����Սuٌ֧q�H�q�����q&���s�Z�P��v�Ye�ۃMD(H
ىVڭj��Q�5Jkl ��E�B�I!��HQQB��HJ��JI \ �(T�R�UveDU
����TPU��[j��� ���v4AfQQ@�H�(%%��   &i�*ba2L�hd"�)IR�    L #`20110�L�L��!)U&�       $	�@I���454����Bl�i�*��H0 ��4�M4�13�>�x}�z�`��꽱��1��b�������Q��IG�*"��� ҭ��UQF���F�n�+���?�C�?�A��<��1BH0�""�*�(�(�,��$V�QG0=���WXǬ���=�^�o�ӏWH��5Ju�j��/"�dhpʏ�H{�¼4Ǹ��i���3�>W?A����)�i��NW.Z�	��)ظ��t��U9`ִ�̕<�X�HL*��%�a�ٍ�θ��/K���-�2d�l͑V��7Qޭ���ta��e���a	��^fvv�Y�&hG���w�����u�M�8�#�6���c9�N�����T�P�C�u������3���^H01�39��'Ŕ�Z�l޵Ւ柕+�#�R賷 ���^X]4���v��\��1������c��ӗ��k/W]���4�ar�٪�#x6{*}���Z
��&�T��]�BN<����qMa�B���e�E'@:�5݋J-�v菶>\��n����m�:�i���;�n���f�yH���5t��;	I����l=���;Of����D���[(<!/3l���n9��t\��ji}�ݲ%�����s��tSm<��NK4�����A$Ԣ��ܘLt���:��p��&�����Q��6��Sx�-W[f5��a�i˸2̆��	�sY���߆_�>�X�4��Z݋v�"��UMҬ�Z]��2��[���m�ȸ�[�C�φݚ�%I���-��^]���\)Bs���,���.Q&�KIML;���N$�T.������.�E�˷p��M�͝��-�@�%��ob�9-5�S��š��#�ˇ�Yj�]�\��#�* H�.�/`�t�C�e��+~J�ݻb\b7r��)��N�a+�k�9^&�団����k�4�˧������2�� ���R�V�.��B�-�����(�[7]��ñi�dP-4c҅�0�î�^��ں\f���p��:a��9��Ln�+������C`ns�V��IgW��5`������>���\{���ɦN`I��nn�✆�&g`�|��we�Vܝ͌��wHJ�ef|f,�"�朝���z�=#�<���&GA�z��޺�\�X\�~!B���t+5!���ޫU�7H���$�v���*$v���4i�nF�*���tl*���gWx��=���u�9�0�ʎ嚞p����Ni�岈Gwc�7D�)C�!����B��ϕ_Ma��3̏N�����4Ԇ��B�(��4`Η]"�n�E��i�n�#�p��"G��⏷=���ܴ�`1��S𢽯/,WV�&ݱ�%{�4NѸ�|u���z�0�� ^��R���]��AaŚc�[��I���f��\��F%X����zWÕQ������bW4ܬ�����Q÷6�G\A�V����8wp�3z"����(mZf����w�w�{n��y���Dr��@�C��p��$m�6髊,�����R����f��F��K0�}ƼQ��.15k4�wr)��ii-.m8�i9��ֻ��1TM��
,;�P+'�}�	8F�Ԇ��ԞNz
�&E�6һ��>�N���=�t%V��vN��̓�x��TE�eyH܇c�Oc��m�h�]�s٠��D7����&&���RLb,Z�Ttu@���P{�Y�_m�X�7��Q*�iov�8ꛅv�K�5�oF����W�C�永�ǒ�΍��ŵ�זH7Qrz�io^�����	V��]4�wf�Բ���t�ݙ��s-�i]��^WuK1�6.5�D�����E��`�:�"n��lY�9ۀ�ėxhӴ�t.�g9Qt�;IΛ;홁���8_D���ʹ»�:�2������p��G��F!��M9��g,��v,�ٽ0f��xi�/A�F���ٷ�y&d��%a�A�;�6�,���W	���0�@��ǊHe�̡-���y��v�{�ռ"b��gicU�w;&��OX2:�-R�c
��1�2�cx����QǃQ�+�
����Hw5�j�%b瑩���[�ok���}�%q@��oi�{��Z�u�X�ே]������ҷ�bSi��sݻ�2�"]L����H�sN��32������	��)���.�M��q�qn���m饧;&��A���^Yz��9�����R��j<5c�KA�_�=��i��%�nM"qM�������&��`X^{3=5��A����y����㵋ս�nSc���)������w1�kf#�S�X�tZ���y�&�W��9������q�8H��f���3��<�5� y�S؞�n���pAfGcz�`'A4�G2�W]�2�?v�����:&�nA��`kAg�ۏ�+zs��`ﱙ�f���\�c5=&\B;h��vw�GR�f�!w�N�n�:�ҧAڒ<d�zY�s�.u���m2��
1͸yMӜ.6N̚��]�N5�w.4x���OD�;y݋@���VA|Z��M1��w���9װ��r�<
����L�(�m��RIq��GGi��O��E�P�u��ΒO�eô��F�f��\�O!�{�p!o�i�1g���v�=5�n�e�]݃z��
g8��x�Rq��6���y�vn>^���h\xp�oB\C2�����K�T�ca)�0�=�%��]�����ϓ�PJ[�C}���EӜ)�7�&m�"��, ��3.�� �,�ѽ�ssK�4l��FP�:����[3��Ę��	�n����������xa�3�@�<QW��,W������ݛQ&D���#�{&)�{�7�k�صř��8���q�t�5S�J�쇸tI�kst���W�um<-��M�����M0�(�;Lc3�5�2��^HsWlC/;�^䬝���hթ\'ۜ7�D��l)�{37m�����(�d*��t�)-ܹ��ǣY8�5`7fi��p�{��QݯH�9g+�=�Ix�y1q'b�DsC�>�����NepQ�e+�Lg�1��+��1�\�7U�6HP�Gc�'X��>�˕�`Ε� ��-9�W�̶�Ƶ�e�9�[����W��#V q{7"��8�/TxF��wx`������KrJm�I(�%m�)��$���m�X��b��Q�J6ےSm�IGI(�nIM��%$�m�%6ۤ�t�����n�Q�J6ےSm�IGI(�nIM��*�ֱtnKSt��o���_=&蠾ĥ9�-���'Fw]�x��w7��՘���M@�VXPԂ�n�	&_X�L�V,Te��&����ۭ�CʁT*n
���[�S�Ҙ��b�L.��3�Zk����N�6j�v�h�������?D�	=�6�ʛw�Wqy|�&��qY�,)�#mK���)�|pmO��ܳ���6�$vp0bR�!����k>�o��{_(���+Js�Μ��U$W���^���Α��a�E�`�%��O-��T��h�K�����d;Ӗ=�X��hY<C�=����h�X�r��4/�X)��=}�+��F`NuǿXf�4w(������K $�w����8�1r���Y�D,�9�����C��nz���^R/�߸,�jk���6�62��ɌL�4�`p�|���4T�w�[�eط��;�.g@�ۊ�Iv
�u���F���a���x�>#��<L}��^��;�: !��_����^�X��P��QQY��}�{�dV���n��O���%�l#�8���5�h�� �:iX�T]
X����f\m��h�����in@��M�rhQ����&� ��:�Ĳ�裏���������i�]�!�z����IQ3���ԱĶ���%w�*q�s�)��Ю�(�
�b�=�0�3�=�ڢ��V-�=�7<�!���]��n6떚�6��o~�`?���N����A�mh��u��T[��h��U3�2Vs�����f�ڞ�����Ԕ�\��{�WV]c :ݥ!yd�F���Jr�{$�t��v�6�|�!�ؽM��6Ly(�7};��@s=�̪
��*�s7w)H.ӑ��h>�Ѩ�O_���䞰c���{�5�M��!����q���:�#C`H�sf��`&�4P1����*`C��,\{h�nK�L�1=�s\�]f^�¼��aH<?]��U{��9��=9��д��{�����O·��������b�����'�֯�KF��A��$�n���}F}�����!�3�:�s0�tB��I��Kw-2�ζ1PޱGY,�)u��^	ˢ�`��%�����J�����;\F��'E���շ�9�W�DFi�W-�yj��7��lo]��:�>�F[t�	�.�[�I�1+Ub��]���g�.B��!D֜�=6�z���/~r��P�m�6Qsn����{zX�6���^��sӲ�H�Z��y��|���,/��u}o�ɜX�ܝgB�s�uF���iݹmB�a��٦��Cȱcϥ ��k�-ńV��b�`(���xu�˓$-�w�LLy����k&�B�.�]��FG1���z��6q�)�4�STow����V�wsFl�ݞ�V���-�	�����q�n��/q^sl:pJ�31	V.��D7v�cg3W����t�X��#2��A%Y����w	ٳ�ί�s�Y�p��~���9ڻH�3��r��a�O]^`�\�b:[֯{�wf�2=�Q��N�#%��M�\�e�Oyof_2S��N��
$�z�#7�3�lzEm@�[�z���Mh�p��w��íf�Z�N7Zsx��8�:D�},B""��2N��I��R��n�L�M������g+��gC���&,�pe>�#�=pu�J��p���Y �շ�ŗ6i��k���<�	��b�q�,v�u+����[1�u���zL��gn���G�Ǆ�0�~����~�My9���X�(��ܛ�i�k����k���߼(��t�����_	�ObS�)�5�N��e� 0�XsyV|����ځV�(��~u�B��{�`�:�k��G��a���stG@=�%0/I�<m<����l�h��V�2Ѧ�v_�,X8w6�� �`'E4�u-�z;U���@��k��Y���=<`��]�s�޾��4e]��N*W�7�s>��U�������5�M�|g,5�y�	E<$Z�&r����o�Ø�ïK�(Ǉ���e\>7`�y�љ�༆��ɂ�f�2���^ ��]0���9׶���2�.Ǯ쁜�|�w���aU��f�ȷ�u��w����A �1*�G.�z����H�A#F<�B�ct-hE�Z�-�0��a@�dC �ݠi$τ����uJ�<��.������Ӿ�Ň�p2��A7u.���$�Ɗ������'��Ф�g� �)�%���T�B�=�$m�SE�iv- f��ā�����2݌]D��[1B7d��Q�4f-lک!�r�����\���B�1�;�i�N����+s6��@/U!���)�D�}�}uu���Վ-��N�L�n,�/<�$�#FQ����2�[��ڢw#޽gnވ,G�&���/M>�}P,(��"�4,h	�u�vg`�X�Ʊ���)��R�bGo�7Q;�cd3{a�˂	Wv"�]�9D熾{��H5�y/%��q����+���S�pK"aj�OF3'����d��pr�'�=�m=�SQ��� "OD�+`���7>��aem��f�nfj.բ4�]��S��uF��FR�
3��u㾅��\�[���_g)�e�<s��F�2g���k�������å�Z}�E��SG�)���{�2s?xw͑�!�OoOQo�:���ښ9[*R����/�!��ga��&^}}C�O}���p����ګ�p�Վ���}���aZF���m�EG�u�S&oU���˚1]���mMs��GQ6�E#�U���3.��)�6�wf�4�϶��Ys��!eW�t��z��n���zA.C$}���IY�QǩA���,��.�:�'Op�����[%Z���t���c6�e8n�&��&F�J���572��G��ڶ#���2�)��DV3�c�O*�#�v w)���IH�nIM�M#"�k]�aTrB�j��I(���$���?{�#�?1���Wb}�(�(ߔ���AT{�P����v9> o
��?A�#���o���'�#T�`/������gt���j��܋���n�~h��q2}�Y]u���͙����yHYgu��^�v��o�>�[��7}2Ȥ-��������Sݩ��F"'zs��\.�#8�4/��3%�ȅ�6/"�!]
ٱ�Ǫ�����p�LU�z���Ÿ�?;w�l:lOg^T�r�'x]��d;�[�h[[�k����+����3e增͑�G��������9B���ʹ�9���\����~�'�b��Lb��+�S�n�4��hSaՏzv7�����t�����k��T�#l��Pǭ��񺱩�+7!����L��b�����{�l�Y
\ؽ�ȵc��o�F鬆]��ir��>��z�'Y�,`�$W׼Or}�ٗ�=�r�#pp���ܼCȇt��:E��0 qr�zp`�zA���\�t� ��0MV7���jV�̺3]5�s̩���Ma���a�*��.n[����u�\jM��o������w&ԧ�F�-O^��S���HP����vR��_c�x����k��I�`�.¼���x=�gK���lmaw3�Ƥ��`aC�b0��_��vV-�bn�����\o�Y> �CǾZ��yYi�O��-qW%���1���3:Qxu�yfR�(޷n�Vq��0�A4{rok�t�M��:H��h�_,;�J�ǅF�S�Nl�g�E`�0�� �c9���F>w�1>5�ڱd,c�ѸN[�{��u[�|�RN����y�S��%���+�'⎙�� ��l��ٮ��*��]v�X��ܡ�6�U�C<��Z��5"5l6"�h�w���fِ3��e长b�>�p����c����d�b�U1:�5���m����T�
w�KQ����f�RSv�v�J�r[3�{<�6Z!�;Y�Ғ�̬�|�_b�
T�+�f�=\�wf��e{�L���H��ᡛڗ���8�����B&&6z<��oU���2�R% �ӛBMR�ĕġ��{n�\.��wj�nt(Y>O�E��_],Wo���T{���ﱣ���p]�+/.��wf�Y�/�J�&�s����^��#�3*t��n�Ý@4�(�b�B��{�qcy1x&��� �,��Rڼ��l𖑽���k����*|����d��ysU��<x����p�$U��,����]�ie:]�m����żl~�ʇ��	�g=i\���y)2��LE{�\��̸1p��%��
+���Y�\Go����50�͊�~!�_��\žf3�����q�Sv���vgrۇٙ寖�9q��t36vI�x��s�sJ�5�#�b����4�Ţ�����yy�.�iơ^B��+�>�z`9�[:ϸiV�8�y�x��cA��cY�7�~L����[�JChP�>��,�����w�w�'೤[��U|cM��n#�n�g���<��N�.�='�g̙�s�����|���c�=qL�S��JL!�y���-��vQ�;�W45w+ڗ�%�!���̻��}r@ �E�%Oy�j㏐��
�eW�2N��6�f.�Gs3���&��:���&��%�?H�v3������f<ӌ�>��eos�I�'o�v��
��j����EFO��pp״��:�B���W@l_@hK���/�=V��q��,���q�7���7}��Vw
�!Z�!�Z߷|d%�0��S9��gU�������Z�x4}Ξʒ�N��Ps�-��AҶ#�JFsvY�H]�6��$�=��8s0>nx�;��|��{wJ㡜��Q�g*�S��}j�HE�Ƙ����4�h]�T�k]����	$�;�c���8:�-��Oq軭�T��x�|����K�<��wI��Q��͸"�9�}��4Zz���l�ќ��;G��6
�9�bǦn`�?mf5���~R��W�V	��v+!�e��_h�'���ؤd�g-q�Q̍�7V�t.Y��\k��o�T����s{�ȵf�,gf�=�w��m��7�"佅,���sd�L������I&�*�^Q�������{�r
+����&� ����﬩:����ɵ�G	��J�Axa�Xn�QF�<��K�6�t��zv��0=�X��ދP��߯0�r���{��|���WbU(��{��y�'D���Fi�J����<|GYw!�zo	Uշ܁�6�Z{6��.	{Z���I3���ނ_x���.�~t�b�o�����U�����/}}}��3z������y������<Od{%,��o+ko�W�j�w���Z*ڈs���g�y��g�v��s�{6���M��R�S�l����ъ��^>��x��qi�t��k�,���3��G�ul�����}�zè��᳾c��X���h�8�/-�
�.�9cRW'�rsE}��
�2��0ї�E����=;o�Rݙ�Q˻��݁]@#k��R�$���h<�Ռk�'^Q�Ov���`i2HC�1���L�=�h^�|���#dn-d[�g����b��w����]\9�\ݚΘ�÷g�i-WE}8X���g�W�x��{�#n9��o�7��������'bWM�n�!�w�I��^ڧ{uw�˯ǔi�>�4�ވ���okLHexZ��r;��e��U��x��]�	f!�ޮ���$�D���ׄ��Cwn
Ϝ������wx���f\�r/�cq���������>��zHxx��J>~>ڤQ.���ǃ�{���X�o��3ʝ^���>�͕�c�Yb��܊KS5�Q�oC�s\hW�P�V�~rl�=���m-�#_����E�o�ᇯ�.�$kk�s�G�t�i�z�e�nֹ_w����NUP����$����6�1S�+�m��IѸ�nU��c^����OpUfq�%�ӧD����Z��}��x��_鴺�ry��c�bÑ���f�Y<5z�!��ac���+�N�r{����M����qj��x""�H$�z�x�C�uJKС(\b"!��Yퟳ������d�v;]��z�]���B:�-�;�w|z�܄��9>W��Kr�DB'`/�h�O���,89#ʅ7Gv#d�	��'�Ϝ���b;l*�βP�c3u��xiq�Y�mN���:rj�·��<��K�Eo0|���ܠ̟T��bs3Տ�O��W'���5�l���n]|wc\T�֖��;x���Bg,f�㯃p���wE((�3oN=)_R�k;&vl��4�q�eR��[��m��=�b�>z� ��WB�;��ɂ]u%�}L�[y�8�hئ������ķS-U�+&���n�#�ִ�1?s�5�n��fTu_)w��r��M.'Hz�r�yQ�.	.99c�e�{���x� UDt�9Sb]����� �.e)tiT��% $�T��_!@��I
9�JKQ"K"E(pA ԋ�Щ� \�S���C��D������bld2$b��ݸhhB�q!cK�dm4����*Z�&.6�>lقd)S�cI�&a J�u�Q .)qB@���j�8)�M�Dt�DY�$�pkRB	i�! �&�!��q�er\��6� �H$ĸUH�Iy\�	?}O�$�F
����2�JE"�|@@pt��Ɯ��E5�Dj�T�/�>���y)"|�
�TM�mJ��t�8��}��$�����z���0�$4?�?���)�������F���1�3
n����ng��8.�
t��V����x_�e�
څT��'{ou��5�@ѹR��e3��ܠ�sS(�~1�o�UÇ��ưQ��=�	��۝x�
�et�t��sx�o�*�y�V���%W�i�=�.�(Cy1���������<���3
U������5(_8�i�g�!���~D֛g��P�w5S��ŵ��@SbNw�R�d���������M�����aC:�J���ϼpRSb�pd��-��A���4�(o�u��l�I�%<���u��1�\w��>kچ��x{)���4;7�����BhZ�<oХ�q�ao4��|lT"�����+ϭ�|�zyE���A����y��<S�o��K��8��u7� ��ɞӧ��cq�MGe�^�]�V����6^p<���W֓[ �]�V� ���q.�ua��gWw��se��wn�/��q�P����w��<�K���cZ��4u�Ǆ:$Oy�1b��PѼ ��ǉ�_��
V�U��Z��{B��ܕ�{�yVP�\ZǛ"h23�X�յ����D�Q�&����4��Ȫ���|Q��{}~&�d!�p��|BU���$��yֹ��V��P�Q�bL\R���2E`�ݻuyb�,LF'3�Yu���:gw�q�b��&7��6�Z͝A�Zo���
�zXi2�4Y�ݒ�i�'D����6�2T�M�ì����~��Xqx��"���c�U��H��f,�cϒ����/ݞ�YA��i��뺶��XZl롇}�X�'R�k�W9:2�8�Gp���֘!��L��г�te�����h���b<��.�)��UlZ(ΐ�ckb�.m�FNˊ�wn�A�a̕�;�OD��Ǭ�N+��w�{�X~l�2>ڼ�z�?��mw��<�<��-	Ndv�N���,Pu�@��|S�V�)�S�>�tk���֌���5��8H.����żＱ=���ف2 �2Vٿvh�3��Xއ^AĽ汤�</<;Wg�e<-m:Sv�PK�P,��<��*n�-Ҿ<_�l�GDeq�v�N���>~՘�b� ��z���;�|Z���GƝ����t za�ZtUf�cjWG�i���3�d0���4�P4\m%��N�h�GH[���T���^xL�f�s~�{b�������ھw4����ܬ�
45��4�g�Ζ]�qi��H��nT*on"Q_8\�h��̦{��T�~�j����o�D�o����tty<��T�6�*�:s7
�����w܌v�1~�$ѰA��tc=C,�۬/n��!f�����Vhqg�ş><�\���M�ݥ�5�}VV���]qYE�qȗ`�$�������H�3��]Zþ�u�Qh��բ1�ۘ�m>��������J+��e�����ڵ|�7�슞^�p�y�u<���6��֤�^K�=Y#�Y�J��%sv2˰�{Á�kP�It�_�5�=�\;�fiN��v�*l:�L{���J;r���}B�K����-�[��WrO=t~C:6������S�r�lY�q�]�t1��CSS4�F{��������X��:*Mĺ=�z9�i�@i4�@�Ts�{�>��}�M�[8�J�����j�u�0��4�J�>Y�M�מ�1o_`c�R��Ols��|��1;1�̭X:`��H���؄���[�i(��w�Y��L���,�QЍ�i�2���=�T�b�E�0�!�O�ϙ����P���xdvzr],����4�\<�>�X�Z�=]��G�sx��#Ӎ�,������;cl�9��Ҷ޾"l�'~cg7��np)k�G1<��7J�S6����{԰�_�����+�j�qnC@U�ʫ[zx�+���2�-�ò���t��u��>C��5���7ՖJ}B�瀫�őq��+�g�M�:��ӕ��*�hX�u���g�R1��b�Zr-���3s�Z�29HkNijD��Ȑ�M��$�ק��y�'��W�ʻ'���QJ��ϐ}�û<�+hgV,�L�aG��Wܸ�s��μ1j�j�/�M���d�To���z��٩�T��f�8��Ѹ��2�؛4�L�x=3m�{��^�Ӣ�-'o�GNi&�c�`����&� ;��:7��r�)D�l���W���v�i-QJf1����kTM�>��/(�	�G���b�V.�o�9)Һ���و,�Kd��y�k���ӺNt瑥�$y#k����z��Q�Һ��`�&���Q� ��bTb�
��ٶf�͹�A�j��hI�<[��8����9��lu�^}Rg��n��Z>��+f�Ƭy�r��F,n����\>�es/t��lpb��ix���-s
*`�q4;x����
Rv2m����qUO�x瞹�ڙ�Z��e�����$�������c��RwBkN�Q�x��Pu�1p�����7���fe���p��B��t��2�oɲ�ٷ3r\���-	�o��e���e�����c]&n�w�j�u�S�j�9�u�w�IP컛�M������\��ڪ�z�a�׎�G�G*<�-�P�2ɩ[q��I� e�ԸF8����+:C���z�u>��e�_kol$�޴���b�����V�����.2��%+���1�]B�qь�e��}��؜��{cf`S8�����=���	�a�}-Wp1�[4,� u��k~���0+Ɂ��jL�����y�w���/>�}n�4:a.�R<�������Ȇ;/a�l�k�Eg`��(Y��^F)�7G���}�&>�_|�&��[t5DA�l���[�aT)��iI�������-$pf�4��Ӻ�clT V8%n�R�y�ڤ �shd̷7ǋd>b��ͷpl����/o5ff���nk"<qHI�n�ǲ�Y(�њŎ��Ԭk\�(݂"P�.�k߬i�J`���IA<��	Q׹��qz�v滸�ăoY͒�br����9�!����R,b���6�VA^�E�)ϕ!4��SN�1��S�����d����b��6��J�!��9]ʬ�w+Ea%� ��Z��)bIb	b���e�1��w�[��Kb ��#ĩK� Ld&�\�"	qR��R�rX���$��J�L���!
P �a-&)��p���N�rؠA-�Bѐm��)$аh@�MpI�E�	1 ��J\�&
8�G
iȒ	 @�!�*�SD&�. ������H�KR�q���mH8တ�#��
�E�$0"K�M&��fR;	Ό���۞�KV%��W"S7z,X�ض���*�����x(IL�j�uZ%7SI�W����fx2z�2�����=��~
�M��F�B�S��}�z���H�<���9�������{���9j6T/�@q�U��3w����l�ߐZ���ߟ�
o��N�s��WG�c��w���h柿z�)n��<�Y_�1�A}��sU&�N���p&�`�7ګ�G��vAFF��x~ 7��)lWG\�����Q�s����_ڡ���H�Pz+�w]�v���t�=�_D�TU ��2��V��;���5�Cg�u�|���|�U�_��kx5Pf��t?�s����G�M������"��D���=��G�c�=�)��Y�"�����1n'�����_�ϕYoP���0��U������|^~U�ʋ��4MZ���/~~ʏ�G�O�Nu�Z�?_q}�}žn��863���V�������֏�o�x̎ߗ��s�.�!7�׍�ɶL��a��s��DX�_gS��>�7���N}����l]�B�R*��9U��YWLy�nW��$W��zXK�w���Õn!����X��0�1')�Uw�}U�q)C��6�~�}�k#��F��|s󇌍��}^�u:VR�}�*K�x���W���j�<kƅyl�N����4e./Wd	4���qYLc71�Q��G%�k�x���^�0Bl��D[���1�V��E�vkp,)���q�Yjn�-Rgk�u��v�t��
�Bco��Y��;^x3�ZU^���~�|�HL�����g�����^T�����	���G�����Q8��7X�����$d�7��L5��E/#���)����ݠ��������ֹ����bJ���EDB� E�K�_ʾ���7��f뾅"�Z@qp9�:��H�l���#�N d�QP��s4�0�� �]�J���/0y�^��x��;����n)��)��p:���FwK|��+7��z�
:���bکS����Z�0�м�����I��Qy�hC��[�v�c�]t���;��=@5E�W���Bؤ�Z�w�Aa����P�I^W&Oo��K�x��pH�;��+�A�Y��Qy�fu&hCQ-�	x��5�k\����5���� �`������n�M�N�%����<A5%�B�)"~ܔf*�����G�K@��P�ԉ�$8�n!�qMsJn.�^�Z[�u���Hj
���o�;�5��jb)���	�7"�h%��'�"�CUA�P�7�n,�c� �-���ڨ�M�y���+�8θB�/��T���q�m ��A�����Y���:� ����o&L�u�g~���+���:�a(� �Ɵi]���G}9��WH�./��#�2�r��,����5&����u��wUĤ������;"nQ ��L�m��W�3�Ia�P��B��/
�J���ٱ�������h� -�1/jT�hz�j. =E3�#x�G����{�Ժ(K\%�j�K�QZ�#��D+�C1P-o�!�,�eG�I{�̧]���Q ��(\#�
���#�Sp:��W�)SQ:%b�"\I��Q�z>�ϫ�Ͼߏ��)qD-z��]�9��Nⅎ�8�L�m ��s���Ak��Y��М����D����P@^����)��\�T���x�%�)�Q���=9�i�߹��ut�b������id ����j!��QpΫ]E��)���:2Yћ���b^!{�"�HK��4Q`��E�S���\�V^bq�SdB�B�N�����f��B][sb^�-���k�8��� ��n.E�j4����$�T��ܟ���{����
TN`��r�JZn�N"��Pn(X�����9��W��xM������h���&b�/7-q�6*�η����76��b�j�D>ʒ��;�zRiM�'`Yˋ�5�ak[��܉���ų��]�;f���Ł:����\�/*)�C��|XCpT(KHMy�� �$�����%gv{y����l���Au��z�[4���P���!�B�Rs��P�7�������Y�[������"n� �P�u��I�����	!�R$�����tC�k�K@8�]P � �(q�#�^���g�F��da�:�Y�o���\�C�PH1M@������x������QL@lC- /�!�o�z�]o[D�:�$
ƬE�SqN�!���9�. �A�@��*d��=o�ѣb�<c��S�����7:��TΨ9���n&���M�dB�R����T�[[�%
�Q
�|$�8��$,u@��/�T��:����Ք��V��ҧX�z�yꭝ�P�����@�0�w�{���C�	�jຉ�8��x�m��K�z���\�k���qA���܀�j"s1��\őAu�4�b}��ހ��?]�ƾ�߶�ԩ�#@Y��T��חr�,�ķ&��iTƭ�nvb��Tk6Q��D�9U}U���2n-�5l��rt��h/c�XCq1�n��%v�1 �W��5K sC�k�j!��@�]��W�G��^=iF
z�G�����ڥ����;��W��mn[Grs�3�5�*�g����ݦt�3^ͥ���^�5O��>4X��>	'���cj����&"FNaZ�Z���Û�IZ�S��s��o�+ޢ�m��hy3���|a;!��1�Z��h��5�S���f��P��t{����?��~�X���{��^�{}*Џ<�M>T�/��˒��IV$ץ�]h��{wE �8$~=�G�s�z+Fn��3�w��"���[���������e0����� ��	���a�����mE_`��~�y�����>۲n>����#���q�\������b���y�1L��pt\f@�
�tb!C�V��Tσ�gxl\+��5�o/$���BR��y
�w������� C�0�:����,��c���R��齊�"¦ɣHgow�W��$z$�Y}��)�|oص6{"q*���	���<9�;�C���[�NI�s��E�+��ؗ �`�Ȩ� ��k:�u�wk�����3#�z�Eۻ㗇��+Q^��-O#w{���A�[��S��U9zV���}�#IjoAp���[�W����Z#w]L1X�f3��g�0�Ae��=n��eEs�Ǔ��V�pJ��0Xڿ=����`�ж�󥚻r�(���m���E�A�琒(x��ɂv�}�=�x��¹�&�D�M�@�d�����g����4jܖ?%�&~�;ԩA7V���"�9l%���q�|[<o�;(��$ddD$@$T�D$EdE	 �B@�|���=��^��B�SY�՝6�/P	#d��(�h��</?���?"��|n0uDq�9ܗ1��+��}r(���������W���泱/&�GXk����r�xS�g��2��X��:`kexi���Sʈ5�&��|���m���c�lT>�\M�E�4ҹ1Q+*�;ػ�'wB=^��p�FN������oy۹�#���G�sb�u<���i���ӛ{J1�+��J7��wg³÷7�Y7����۰�}�v�7�9fĮfv֐�i�6��͵1�d�)>̴� ���B�P7V�Ro[��ݎ��6�Ea��(%o"��)ګ�N�����89w����OޔҬ���M��ޤ�J�y���p�#6�H�pFo�=:ʛ㻿+����\f8_���%��S�=}/���]��mU�X$�m�\��O
ؒ��x���4{������7���׎���*z��c�PB<і�t�p[ܹ�K�CWܖtw$KϨ;b�~=#���b�$�\zu���8֫f%<���X��|�eWƈ&�&�ov"L^f@�\���P���mt0�ڤ��4D��BĲ�/c�$8�kL�bi�1��C*f�$)ʒ#SOXGu�N42=Z��{;��R!��_YO�trq�3�qd��4Q�ta{c�kS��b����D�Țc7�5XxNQ�(�BM͎�w1������r�;��ԚC3'��x��³vm�n;hT�7�e8����q&<��F��7\;5R�A5*dT���Qە��l�Rcë>еT���J�q-�u�r'ָ�A.6�o�n�k
:JY�<�߰�����Q�b�K�!�	H�$
Z}l#�3ƾ��� @�sֺB� Dh��&C!� ������$@
ZhH!h@$bj8�RDN"aQ	��i�2$�����L�H@��"BmEH�XH$##�,�(��U1����I���@4�,h  4�.��BJ�$j@���F�� ��6X�Jt�i!��%�'o�BK.g
)]�H�8�i����4�HVC�@`���r�5����%�W��GxZ8=��4��'f-��y�a͒a@��
��	)b�G�=����E���,�_���WI�ӿ��'�9���;�:�k���6�F*�����:K5��Sڻ{�h;�"OQ�y�"�j���f�r���-^/�;We�۞ޫTa1�'�օ4�y���k�^*.W�ݾ�ц�����S9���a��#>��Y�#Ե�s�i�M4t�G����r�P5���#6b����{S�w>}�=;֟e^�\����P͇hmF�q�ɸ{�Uci���35I �1oT9�bof�Tь�	�������
$��obԇ��V H9Y&y��>>�1xy;���جѤ�y��09*u�e'g.'���'O'�a�V����ZojR~���d]�<�ءW�h�{:���կV��F�m�����љ�8���^��L�ސ���^﹞��dמVӽ�,֚L�[ݸ�f,���^���
D�N0-���_��_�t�~���}��c'�;��*�Ѭ;���i�9[Xd�GML)0���)�oP�����cg���{����[���<_f Z9{Qq��F��������vY���Q��-u*h�8��o�+R�WP�}��Y1{�G��aW�*:�W�gT���]���xs�F�&��8�"�g�q�I��7;�+�q�2�ߊ����6�q/��NT��HJ��L��vL�(��)�F��un�Pˑ}�I�M��[꾂K�p��Y%�;�Q�!�;�k���@�n�bov��$9����xd��Y܂��`�*>lxI��{���	k;��5�3*۸,a�-��و���!Np����������ִ��W�x�)~�x6l�W��l�x�5�����ȋ9�,�@�_��2�Ō�z�g����:9�н���$j��VsM�q��·�H��I���=�/8D��kX���E�mKq�u���9���%���aV/O^�t�ޜ�<�].y���08}yiD)fbP�������p�{h>]�k<R��V�l�v@����4^�7�Z5�����'x�zm�ھ<��a��\s�mtmd�Y4���s1#�/R=z=�z"�ů�����Gm*f*ج��/����n���0j��U�zӌ�aהu3�R�k~x/xfW`���XJ��[�;3��}.i���8؍�2l���(�>ܧv��Э|�F�yV���\�Ϯ��'�����DRg0��z�����:ǽgm���t���W
4+X}���Ȥ��]A�oaɏ��C3y����ٽ*�^|7����Q���# ��kh��ʶw0}�VAs6�6��x�ƌ�7!u��j�r�_}UU@'����a�{U�F*D�aςл�8�K��ɳ5���zzm��y2�OB�LE9�*��x�	us�35�Q��8'�Z4���֝��2�������O��&v��Q8߰G�ۨ3ۛ������<W��^M�=\���k�O٨����7G���k���4���UPT��MC���Su����Jr :�hOlb�h�=�-��j
wt9��9�?jz�������Qacr����dX�q�GL����G-G�Քw����U����D����_�$y����b��l���`T@��o����i!�<)lp����p�=�]s��s3+^�T�xFP
���Fճ� ����P=cr!�%i%�~(�r+(��K{�&,�1� ����7�%Lmŕn�W��7a�Ͼ��A魣�;#ދL8X�L�����#��J>|4-܎NY���7eG�����2�"�����ݪ�:�[	/U+QLr���A.�u�
=�UTn��a����T�{��y���}`�2��^��4w����sn����Z�P:�s�WQ�ވ��@h��|����L== ޺��ǟJ������lT��s}����{�S=/6k=�B)��o'���	&�3K��&{I�%�U�F�w��J�TY��~�ȧ���~M�����6׎z���ktMl�#Hi��y��][��Ȳa����
�܂ù�۽����w��1ޑ(��9�tE�J�L�)�Y��2,p�¶�I�ݚ@�ɨ��""=����� ��(]��v�h	���9�;�{ղ�}�t�,�B>^��½���e�C˛�O�[�Ŝz�]��<�.��e��D�X0ҿ�וr�I�]�=�ug u����50J�<=^l�3��ɩ�B���z�f������[�Axv�wln���������I�J��x�gV9�g�:�yЬ�V=p�����'t��Y�O��)�%�3�s��%�}�e�1e�)�²��˽�sLf[���8Է��{����>�]ފ^�#��ޡ����*g-�F�q�X�J��w��*2�ڶ��燓g*X��e��uT��@��8wI������O����H�����E�j�+�v�oq v�4�J�F;o|��'S�FkVZᮚ�ڣ��k|&���M�ͥ)����p��x+�7F�[dhq�8��t篻K�~'q��n�%�_=�5;��B�[���W�:l�s�oxb�|6m1e�y�;�5m�%��z��d\�p��i�y�؆R����}�c�:xƽ�C��*��ݤ�jh�7
i���>G{0m�~�2�s��d���b����,sF���1+�DY����]�Pi�ৠ�뒄X.��3��-��)U�)ϔ�ƇfԸUݫ����n�j�>�	���S���-[����VOR�7�_'�Hx�X�1f=z�!�j�Y��D����${�;{J��O��5�^r=��P���@O�ʬx��q?��h�[Vh�ݚ(�*[��}̽N`H��6|OϮ�Z�$�I2pl�E����6�5֭Pz*Dk��!�.�h���^�e*`Ǔf՗U%iR�X0�����u����8�0jZS͔bl��#�qk����pݿsN���ʿƺ4�G|�$�#y��r5v&hCP��9pE�r⺞H�J��6�ͧH�#A�tA���fBe�UlULَ)d)=6cfQAi���[���b:��f޻"�ŝ�[@�*�XV;�$RDJ�D"�E���E�-X��۫���_E<|�a �)�&&�s'XH��V����)
[��T)" �\²,\@���g�R�[�4�fM7F��L �4�!�M
8�T�Q+�Gx�%�6�~CH �&��k%0@���T��ٛX&&C��T�
Hąc����Ȋ-� ��8LIH��.��Y�ci��p�ۉ�CQ.P�KM���mP�!�dCG\�:��/ye��bI�:�%�D0�ˮ�篏����DX��k�������f���8�^��iGvf4�Ҷg��c�s�)���^5�>��~�z>����\�z�EEg�s���a�u];�/k��.�����K�Rώ|W�f��9M{fȒ�O��+���u[�Vv�t�O�
{5�>;P����i�)�L?:��y�j�F���Ç=;��jy���fL�#���Y�j�Ӥ��ˉ�n�=��T��zUd�ՊJ�`�Wb��џn	���ҥ����FI��ܝ.^D$��hu�RhU�Yك��k��JT��U�%(#����O�Z��wOz���h��W������RS��M���"&�7���}_}O��o8��xx��l�4�l�-]�r֊躾�~���e� G�������{5�5�{˓D�����޽�v�J4f��m���M{ko�4��vX-9ܙ��i8֞3]y�.}��x����b�q9�oMG��u�
�r�}���[�(��jN) /��8L)�y��n�q�j��Ʒ\�^xC	
:��7�_���`��1�Ƿ�:*^�I˲�ɕ�=��d���neaB���k����I�xI�H?>��g}�p���z]���k�ԋ���}�W��';m* _�Z�Ҷr��%���g��/�}U�|Tp�{���Q��Ϲ�y{JR���|/�}�{-����6V9�e<Ed��4<��B��	��n�>a\\
3s]�o%xRP��\`��>��'�������;<i�=3�.,vJ��E�q��fzv�]�Ϻ�Y/��p��ך�(�=���xy��a�%IC�Ҋ�O���#�n����ۺ��f�uv�
L,���0$��煏� ������}�S�N��h�����P.
��"�ǅg�Y�f�&��I�u��ź�\t�����癝����G\Pu�����'�����%���Qs����FG���;\I�|xv5D���k��|���2�B���<�K�l�P�C��٢يv�0aX �&1h����諭��$�X��6�e_�]+�R�J�ӡ�`�St���+:�d��3`4��Fk��Gwh#EZ��)OךM��u�����S�N�7viWZÇz�Y����������%	Ӌ�î(AK��u�op��ՍX�	R�%��n��t��B�ru����wDd�|����m=|(X1.[�
�h�,<S���C6���q{�~8a��cٜrs}Լ��V9{����Ӗ�:�z���k�{�,���_�5c�0�d�V<�邦g�/\���,��~�ł?K��_��|i��r�Wqg���s��5�?k��$͓�.�w D_i��EOR˕-no
2�.�MN]����'?�!$��\�z��q|Ɍ�$&�d�?��e�����KV{<���EHGN����j$Xw90u�o��5����;.WS�[��1r�d��Un(��k���	ƺp�Z�n߫N#�i�KOݞ����vn�7�{G`LJM��/�*z�����^j�6y�����O��xU��?Q��Mu��td�/}��:��}��s.������:�q|ˤ.�ӎ���/e��,AG<��U����{g�c��w�>;O�RF�˲H|�|��n�t^�Dz�mi�N�[�&W����}fB���]L�|0��}C�_ej�y��^��}�����g�5DZh��!6����ۓ�cݎ�j�X������s��w�ֶ����rŔ���
*n�ԙ�����RZ$ZG���*GG�K��ZE�/2��tc0���:ғ1�W�-�&�ݓԧ,�us�q�mY�|:pVtG�N�Y��]�
/��Ϛ�(�R��=mUTro�E��s�8���{��[.�7�1h�����U��c�Nm��x%�#*�L�&�&�X]f��Y٬�{ʸ���rIh�����������7VߥG�,�פ�mh�{�+E�X֜r���y]���ʱ{�ؙ�&����z�t����9���l�ߑ8��y�h�J��2z���õ���U]S�c.P���V艝��hY�u�{ވ�ιϜ�}Fe1���PU8�W�1�ku�����l���W���4[�S��z�N�^\EOkVU�Ц�]@��Jzb�E�1�O��c~��)�v��K1�]��>9mj#�k��i1�h�_�{��̚]�e�8�4Y�i�M����{U=��CM���\��yr��ӛ{3n�ش��aO1OV=�̾�Ӱ����l1�kS�����D��D��a����n���v-�3j��w�.�Fa"xsz�n���d�y]1h�G*=QF.==��*�u����-ƺ���rڜxte��֯��e;.U��O-�{۹�s̓\�v4��lC�,|�a%ܡ�q�� ����
�\i�C�"��?DDz(`Ө����ճx�xX��	��zl�d�n�S&}���*4�����<k"���W�����_wT�$J��N]G[��tf;"���="k{}|�_CϦq�]j�vY}{QÈ�f���k}��E�$��c��R���zO��w�ғ�]��>7�s��f�eT㓓��|�-Z�=T��f~����)��+P����R�;���LP�Q�hM(prp�O��CHX�[M��7^ ��M��}�{e:3�Q ULL�*ٍ.Ⅸg��ؑ�x�Q�l�b�ܪ(�D��Os����ce���:�F�!�Ox�Ōm�E�zm��F\͗�-��fą��3�E�I)GR��@II��U|��ΞU͐�}s�"�0U֨��WE���&rR$ˋ0��s��bb�єh*��ӳ�1ƹ�������;=
fxJ ��4�r�l�4���Ŗ�����˕ꍜ&ǤO��݊�q�پ�3�9�o����%���S炜��>8}jO?Y��9�F.�fL��ʰ<F���7���F�;�1=����yE�K[��^n0�e���,�[��e��y�_o���I"���Vd��u��N�M���Rz�_w3��K:�ļr��(�9m{�rٌ=32Ӻ��ǐ��EI�P�7�I����}�
��K&��;1R�nMUb��O6����=�N_#�:��6f�@Q�3z�u�f����7vwBY�{�������s�7J�D�E��d������w�9^�f��ecJ���5�����"K�Ѻ����y��u���Փ�Ӵ��53ܤ�:vO,���o��c��)0��8֛n�ƞ8��Хnʭ�aW˫���y��P���"��L	�7Tۈ�:�G>8':�a�ϲL��숸�i��yOu [#.a�㘅Hx���4�/�~>>4^zT�����{�V��k�<3�"���q4�s������-v.�*�^�{���醙�(�4.��K�9���K]M�5��9��-S�ƛm)�/�w��mvM������h��}��id�ɱ�)�I�u3�j&�C��eA!���ފ�5��.��9,�9�A��A.�����b�� ��6��q+��G��OokC�zgrm�M]�|���;u�ϢJ�xr����)t�Ź%ʼ����vI�z���m\�"&��w:���eiD�H��Z�n�1j8���ܩ��ø�I�i
���>�8zf�&V�1y�a"�P8����<+2�Mr��7����-���uK_�QO]fn�M���������������ˊ�d���֟��p���瞑��,t��N�c��%iWw'lc�o�Ʋ���gr�'dC�B,��k��hb:��{�ZN�I$�KQ֦ѷ�1�����z=�C�A��G�s���3�'������,־�$��=����cx����R�G}k�ǚ+�k��p���xPه�'2�S�rm�Δ/Ot2eq��aJVV_�jG_K����5g?F[��<�,���7uѦ��[Wbj�Mk�Ǉ�H@�����6o��L��N��T��%�s��+2�5��vG��t���ͤ��o`7������CN�-:*�i���T�e�|\T��w��;��ej[�>�j�̅[ �Sۊ�
���I$�H[qL�$��N	$�ڑ��	��D�o����� (���!&؀n>��Z̕(�%�I�e�D#��RB�X��ƧZd�v$���P!/�0iɖ(�i�I	��SU�5��`�Ę� �;RE H �nD� m�M�Ҡ9�R(%�q����4
�)���m�B1-��AB?PdS�h#��&�h�&�¶�(l@�`�Y]�cp<���s�)}�\�	Ƕ�Z٠a�����J&���s���� /�oϪ��&M�v\>�{�X�q�e_Z4��b�t�<k���_rV/ox\����<�S2��!�M?	�+�{�߶�{����:��}�Tpz�_��h���2Y�����C~�.�_�eN|�keb���~�z���խƃ�k1��aѧE�k��v�g�yxb�H�~�X�*��9SgD�n��n��Ɩt�D,zN���j/9+�Q��F��Jx��d�ˎ��b��a�y?-$�__!ʪ�+�����簕��GW�:22^���U���>�"������݂g��@iGw���5�N�t��h��0gM7$v����}T�yz��G����+�Q4�fs��P�B��M�ztu�>����^zO��4���w����[��~�M��Pb�|F/g�{m1�zu�T����g}���0�ypύ,�!rÞL���3�{�o*��k��+:Y&+i����fx��}w��<�'�>�bӅ�3���7ޝ�.���b�0޾�[�^�Lm;�"�z#j�ʧ��_�n3����ʕo^닽�'u{�����#��xe����i�zJ�XN�zIɯp��gwҼ1'��c�IT�s��l�����'�\ZwB�[r%?c=�x�YI"���#7�x����:�V܏��c+�\w�kލ)e��q�����G;~�~,_-j���e�|��
:x[��qWU�e�����}����ة��z�]�-o���Bn���Y��/Ί�rY(ds���ƻ�o�������OL=�o�-,�FI̏P���{(s۱C%�6�];����8�/�>�������S8-5�����Ḱ̩j���YMc�]���W��:Ro����K�"]���^�3�uuۗ�xY�0[ջXQbx�H��~��H�O�4f<k<�Yl8h��8�K���}���Wx�0�zf�#��o֮)�N�<H�N��,ה���.�3����h﫼�5j*�~��3uѴA�N���`�R��OfcPE������K;�z=`h��Oח1�k�~o�Oٚ��<��̯o�C?Nf��q"�ŧOG�Pt[��ң_H�E\^X���/��v@4!y�q�'�,]:Xt���]{�^�c%��΢��a�i�\:H�e�}�l�{�}�/k�)V��3��)B�I,~�&.Vg�O6����Y���l��ܧ����7辆�3���Z�!���K���Փg��w�����
�V�72���=BX/G.�T9;Y!��J���̒(�����}>�r�L��91�Q0'��r�ow5�@k{��h�rh�Ecy�&c�R���=W{�x�5��ZN�{���/]�Z3r���$��%�Yc�PRjt̥h��"��v�aQZ�v伣��	_���Wo���}w:U�ҹ�={��B��*z^Ο���,���s�]���˲��O�X����
�������x�Z�O_�E=ǻ=������N�Z/�^�o�20��=^�>��u�#<i�Ҕ�y���W��B��R*�٠�EӍ�W�8v25��R�Л�>���[>uQ
C6f�.�FJsN�f�NΚM��y�8E?#�~"P��5;���E�Nt~N��쮬}�D�'��+o;�����,�WrCu8W�1�5�=��y|��/.�)�}{����:wWd:mT#)�ocQYNhn���Ʌ�o����J�Z�ͳ�����������ӝ�v1"�FoMy������H��	D�.�޿$�4b��YB�=c���Y.ǧܮ/m�ݭԷ����t��B��ܼpb���y���~{6;�~�?k^2Z�i���(b�|� |q��)w��F��M4�\FS�gZ�g*��s}}Ƭ����b�Zk�[�xRpSM[�S��+u�+%x�U.̗��=���e���|�K�S���(�Zץv}����N���w�3N����Xp��^i���=.n�N�~�r�ui'0�ikJ� ��o��D�3=���TϚ�N���o��-kK(@���{�z}�͛��x��u��u�[B8�7Ϻ�T,��j�A,��(���h"6t[�'��Ip���rr�_}�(��g�_����ն�ީ���9YK��u��բR��e'�V`sӂ����ڛ�m0�N(�FR���Ƹ��KӢ���w3޾�u@�LvA�~y��������}�E�Nɶ�[Tv����ָx�tx�5����{Z�Q�q��<�%ʶ�i��|�����_��D����5�$�,�%�%�^�(�s�jp]�J��l����kFm���,�3��wo\5mvk�}+��11�fӱt|3A[Ĥ�K��cs�YXtN%ٸ�滯K<{�(N��/���/!p�h�xC���fŸ��1�v-P���o0��s3��#�����9i�?�UZ �VL��̮x/�vp��-�Dpr�U��<�9���kN�P� �sVf��>�JN]��v)KwJ��z��C:__I/�d��,�	4f}�\��f��**D�8W�*aJ�iOZ���TP���fϽ��xF��c�:k:<[Vi��e��o.�O����c�V��ӧ���7OOM:S��Ѝ��3���us'OX���0g��k�D�[^���T�Xa��a-ܩ!�)]i���x�iWw��s��B�J���k�q����U����e�u��k��#�JN�뮵��W�a��=�C�����I��M����7zlt$���Ե�>�'mp�iޫw�
ؐh��Aa������w[��*�'�1񥛫&/==$��}qw�Ƚ�s��`�ɖ���峍a�N�VC�/W��~ק�x���C���)��(���̹��s&;׻Vxg(��iI��ǽ06�O�J�Qo]m7Q̢�7]`> �Sމw5]�c��F�o���b�XU;'ޕ��$\�+s��v��t�{)����ظ�yx������>��tl�iɗ~�DxXw��'��;:XƼ��Κ�=����\D����界(ć��֪f�<55�����Zø�J4�,�[>��.`C6f��a��]��^މ���� ��Y�8	��6��k{hk�%��y��Y5��nw�)ֱɋx)ݬ�)p�#޼���0��1�USW땴������U�C��}����?�C�c�O�޵�g\Q�ו{ު��r@uu��&7V'Ƴ�0��������wr�H�3q�=�jOy�:wfg�IUP�kt�Ѣ��.�N��EuF��C�q��jcz�U�x.�J/Kꈳ���#�zi���@��_/����y1�q懈�b�L�F�x�&�^��N��ﴉ������*���I�3�-��%F2h;����FFL�jdx�Z9��4��5�����bk��X�����x�����"r������>��A[�Ba���o����M�RDImR�3�\���TY9\��E_ʵ^��I�K��6A/�O�&���ܺ��^s{�L>!���W���n�|���ð���[�	��~&� �z0�o0�\	���/����(ڃ��b�,�IY��2)�t�ޱa����Zż��[~�W}0_�u���v���-n�o�������,q�3k�*{��i��ҟ(��g�{�D4�B��[{�<s���1�z�0��^��%�����d�ջ\�a�gT,����V��2C��Ae]J�9�;N�p�x��;������V��r9|�[�n��Ǎ�6�`���z0�~�	�4ښ�̓a�l2A�K�N*��X>wʍ�>�z&ޞ�(<�4�N�^��$�&Y�s�u�ZJ�B�Y���<n����^���[1��nZj��#�4~��]t�TAV����=���޹Ӧp���x�C<�"�|�c:d�5�;t��*W�ݼU��,yw�+X�̝W!m�歓�[����W��Z��Sh`��8#���B){��^���+G����[Ѷy��������{'�ܓ�9��r剻|���ۥDe\�%��T�zO]��^v8��vxp&)�ˮmq�_e ������SFL��QvM�ۻϣn���|�}
������-Һm�(�rҨ_a��n�JC�l{#ԣ["2lJM�������ڛ��S!KL� 4��a�$JB݊�� 2�LK��2���ff"�=qB��@�+�@�C,je�@��*F��h� ����ؤ bL�53)��3*h��QUC��=t�l�M��5]���E�4D����vS�lCe�B�JI>�Hę$A�r�@!QC)Re
��L�)1����I	4ۀj���e,�K|]��`����Y����˷{��r�Ph��r�66��Rq}�f����z+����4�b"���p�;��Eb�>����?O7/���Zt��eI`��	�%�r&�LZ�I��M#
���f��=��,?x��H�B#ߩ[��P�vt��xW{�[�8�Z�Fsy^~|�y����$Zvbe?>�+;=)K[+�W���Z�4�&�}�<H��r�%��>ʣ�7�^���u��gf���������x��i�������/��S��N�$��Gm��u�j	�{ݴ�Ɵ�6��A~B�F�8x�tx޼����j����o_��a>ʥ�n���DF�毠�k��8�c��x�|�����wOL�vm�񋁊����(����\.�y˥�*�W#O9�I2����}Hp�4X�>>ۯ����B���-v/M8�p���lʿ>�j��b�zp���2�z젞�7�����t�c������0T5�+$~�{����(��'�M#F��xӘG����ܵ��cmd	�բ��~vD��	D{�.�&yM׻�}2�������ȱa�u�͙�כ緝;8@iZ���Ek��%J��e�Z!V��~��=���m��xW/F���ӭ�W���Wɩ�$�Ys�o�N��TQ��:�؞���%Ql��N���K��\�-<~=���zz^o�a��f���Lţ�M�h{ѼXp�b����<4k�^���LW35�α��ˀ%������D�;u!�!�+�] ���MI�gea��j���4��D^ ���응um�@1�8��H�ŋ�]��͋,5�u��e��p�s�=g7�y�]7ݐ��M/vAN��9��"�I���e��{�h�r)��W��l|���z��kAK�+���:��{G��J��Q�I=n/�N�������skͧ���"��-/	�Ҩ\��gq��c�U_����f5K=:D���S�M=ᾞ̭���ќ<����M���]����,j&�=��P~_x������@�]���m(��x����n��hea���ְ�!�Cf.zW�`_��]E/1gJ{;���l}��4.u3-�e[N�N�9�'�����5��4Ϸ�v(�P��B�Rb|n��AW�,�u��,�W��v]�����t_Q������F�]�t``oN�R�L)�3a�:p�B#��{l�߯i^�*_��>{��̩�J���v;�[������X�M��O#����<׭���\a|�*�ֈ.ݕg �ra�HN'�6�g�מ�+[�
�jaK�����|��&tXt�UV�����/�4�-��WmQ�ܩ�X/.�����E�-]S�(��#��ϋ�������{�o��>k�u��T(��k_��@]Tcާpf�*Vtbj�5��f�a^���X�G#�% ��v���?�k�W��L��J�N�ے�2���Y�{��s �7��6��pWnK�I����S��sJZ*:�%p���ً��X*7q�*��Y�{n~���2+�#!Ӟ���n�<����?�~�޻��CN�x]:���Qױ������0R���b�a�u��_RXX~��S���sUw����o��u��l�,�����;<�,��D ��#��ح}���o�dT,�dNN���Z��:.ڕ]�s_Fi��<�-[u3�;��_E��Z�j&|$Ҹ�3"���R�;���#x���;A�-�*Vv���6y��)�xD[0�~7��Z06c�����9���I��UV�I���}����8s�4Ru�8�s�s���O�ҷ��u
k@?,8D���������z0z�@�d��!`X|D��B<)���vy�漅޵d����9���	� ��ۂU#j�_�"��܇=�CZѿ�⟶z�ď��8+*�
��}��V4�ӊ�z�u7��ʗ��H�s��qyمc]�3���y��ֺ���q��4E}F\�1��jFYۈJ�Tk��޽��8p��q���������Mi��9P�:�a�ك.Lƣ�R��ұL��6����V�<	�ͼ���t��'v
ŋ".��c�ٝY۝�*�t:��0Ӧ�B�q��K�U��R�p��1������>��G(2�n������'��(�9�	.\|����R��2�������G΋��Ή��jyT�S��6�aH�rt_��s�5���Z*m4i��i_�{�K޼�.b�ײ`H��t������Y�OR|^Mt�ы��n'du��x�������m�󾨺k8�)�0�n�J��.^�����g7$=7+ơV������a�Z�wOs/-?<4bss�e%�x��`��e=��� i���C0@���<:I�q�}1-��U���=y���j<X���bӥ�ɹXM��`ݯ
��F�sYȤ�u+r{3q��d�c�`h�5�ǧ�p��J��&c�\[O�M�*4º�����PH��jeG����t�7���m��ى�S!��Y��Ɉph�3k�+&3p�9Gۿ1�ݛG�E� ׍z��km�3�ӂ��j���{��)�q��3��x���r�k�x�D>-�&�EF�I�Ooޭ$��-�k���L�L���V���r�[4*/�)�	��|�ɘ{s��[4y��G��0�.�������p�X~|��~����#�kIƴ�d��W�V�."�}�4�w�¼��Κ�����7r��2��>���W���oAY6�u�;ѝ�
��/v1�I�;'dƵ��x^�/�I�5��HA�gs|�.y�u$+��ă��_����}u�,=�L^0x�tW�_���ԿQ͍����2��dz�P{�u̚��Xa�w��Ji<0b�j�#��\�+ή�{_}y�
�����>�N
�#��>&v������j4UƧ���q�=-WZj�ۑ��ÿ*���ǭ�c��,[Z�-�ϰUϴP�us��<=���+����o>�t�>�{��{>m�!��9 ��N;/������Nޛ�ʔj!��2'�bk�c].�*l�&s�L���qyc�=ƙF���S�� ���0��k����p+�����WG�!d��z]���M�|ogI�]��=7]-�m��I܇� �8@}:4kySs�ݙ�jk��}Q���v):\��7��$u���Og	��.0�f���B}��_p�N�n��@�r�����]�t�R�iO���x1���i.�ӝ~[��I�X��ō?J��e����ҁ�\WWJ	���^_��׳n�u�5��ɗ�_w�i�\�:x5�2Z^,��N8��WJܵ/��ײ/Z�~���f���5CE��{��O��0����c^�r�_L$�Z[��tK)�p� E0�먺��3)��\��>�Fm�Nez�	��.�&|����p)�5Ҝ�����Wz�S	�|��,��7����vY�L)Q����J��(��q4�#)Wz3&_W���X�x�N*�~Β������;mչ��Л'�c~�<o���9�{����8�X%�a���;K#]�s2�:��]��f1�oY�������3%k����4f܍a^���:��A�h��.<���z�ƺ�ʺ�1�����&6�@��w�$�]8��c��Y�c����
�ׁAx�;h�r�MrAk8:���nf�҄x�ґ�h,��҉�S��jh{5��� ۔Vs��b{Z7�p���c�[/�04X���vu�-��o�KK6�Ni"�³n�S��LeF�1l%4�mHl�E�T�"�s.Bf~�^�6��r7J���Ur�D���׆7��7�CPI�{f�
ËS4�ݸg*�6Q�S�nl��U�ju�jC�CUv�����I[QkDb� d����Ȃ#�5M���k�#D�Lr�S7^4$8�܋)�� mܦ,VI��wn��l�J��.=4ţ(�aAn����+љ`�]n�
4ಅ��yN|����Aɬ�pû�d��ܶW��	fR'�*�K�D�һ���yw�2g/.����um��e�3L!D�@hR�$��2hD��1pjF&�����NP��!��L�S�5"� �TIM�� 6��>i��.�j� kr6�
CnD�\̢A:cE��( 
"I�')�6
��JC��GN)M&���b�C`�2Rb	��Orh
�MJH��+�8�Ĝ�) $6!4�ېD��Q#r9ɉ"`Ci�2?����ж�ix�0BK��{��و>�7�:ھO���{t�D�r*ʔ�g2p�<[��֊��:�1i�'.~Qyy�:����eA�� �e)�UW8
Μ0�k����3���೹+I��>vr��"cLZIf�=�H�n�j��N��C�A�a����vD�Äm��g��[��J�<0�rX��mX�Xx繅r��V��kI/�8.���^�$�����۟O����2破Zuq�D�N�z�c��o�L�w�3T�,g��X"�yفy�:�=BzC�ؓ���'�~\H��7Ԣǵ1Ӹ�*�t���9�$��ƍƌR��鼄�h]�x�ze\�����=�=+��1��|��-�RC,\�i��w�-�N��W��>�W�R3��^�{�{8����˫�"s��ƺu5��X�{*E��)��LT�: O�fL�ZUou�YO��]�b�*I8 K����y���8ξ��5�I��d7Pؾ�T���"y~.`mN�z��E����}����^�i��#��^~���	�wz3�H�K^b��WS~:�]���(BGq0��з��Ψ�z�a�gk�{�����n'��JQ�e7HvA�<�fz9�W�n'�k�>T��Œ���g`��U�w�<ڝ���5���Iw6�>���Tr��{}�'։����&.ك	���RAY��k&B���ϼ����k>#)2�M�L-�*�G/��Wdf����3�хg��w��yQ���j���>}�oo�C��L�=�rb;jni�^10�t!��moD�U�oy.}�I��U�6"�O#�5Da6�n�q�en�����]K�y�������X{�v�\7�(.��(GPp��L2�3���e{�eG�M:��y��Ef���FouoQ*���E7�f��t7j�E��jcH���t� ��ɽ�6��BQw�.?G��F�>�ux[�G����U����Q�½�lI��mo
/��O*�6�гapH�ǛW��-�/�͒�"®4É�]�t'Ct�\p��y�̙�o��˾x����j�Q��7�(�k��t�)�P�K�K����3�	3f\)�c��;ۦ��<�T!80�,W@[D��Q���JeSB�N(^���n�Z99���90������.�)J�72���/�B�!�Q)�ר���!N`��9�54~�T� �,��וt,�{F0�^|fʯm�c��y79XA�G1��e�́�2\G�� �����d�ЭZ׼Ge�=��}������M�ww:��Ef��t/"�U�M���ӎw��9��id�H�0,)�C�/:tQ��.��L.��lZ �)�t%'
`��՞�,w-�y��y�B�T�/�2ܽ��Ʌ����+���ჺ%�\43�\ˈ[�e�Ώ.齨&1�a���̾�Ď�|t��
dwݘ����%�Ap�"��'���Un�/�3q�v�SHk��v�I���hݩ����R�2�P`���*%����T#m+Ȼ8��S�{�*E@0����<�M4�t)7E5}�F�q�^�R�����g�n�Ok��÷x�Xw~���K��rt�U���VkU�$J�ׯA�}�5��d�Y�м���v�I-�*�Q���ctg-5W
�I�n;������w�1���,��꣼Ҏ��`f?�X"b�l�}D�z���p*�X4���}��,?Dz�	�d���믟W�U%��2�.?��Hp�ӝxw;mp��ꛌ�l�+��n��|1���R�e��{���To)T�1m��i.+ۿ�ˈ��`~/I�	W�|���*=U{�gj�lV���Ӑ-f���f3��D̈������b�]**s܊���W��'�`>A��x
��
)�3�n֢\�����Y�_�&��YeߜR�3f�,�׬�i{d	������լEQ�w���M�D�F���.��3!��@�[����~{f�vy�N�W�r�����|t�E���(�G��?IQ�A�E`�q�o��d��o�YX#K&�
��s�&�M��\Yx$SS�-foM��ٚ�"�M�v��d佃qZ!�w�]����bxSF�2�X�GL�d��FR�Q���ge�SNbјp�j���g	�q�n�z���"I&,j)�+ۮ�dz��6U�<�f��i�%�ux7\�O%�ܬ��6seM�l�2�� �4�ӹ�kL��a���ް4kj>ώ�|���KX��v�7=�wXӤB{Y�UF�d�d�D,r�ed �=��TuC;ʂ���X�W�� ��̼�W'Ί�{d_�d����uu�ݸX�滜x�sӵwYww^K�kU���Z�RMQ�{cǓ��:��g�O��dN��9;Ei�g�a+а�%;��yE��A����;��`�����ܟ�����l���2M/�M�eq>�H�����S�8N�9Q�� Ԗ��I���%��ﾤ	�~�߃��¶�lX9F�M����9���)����L��~��c�k�y;$��s��=9�(`�o����-�_n��g��-3�ȼ�SY���aA7�3�$��+�Ĥʍ_�\�笑�nj$�4���h�Al��La]vLѺ'+Q�^��T�\�����{M���r�^z?��ͮ�ڏ`�'�VY�,��ٕy���AC��	�1d�PFg,[%����幸����F$9�˂+���;�yK%�zq����0:�
�Jӱ'����޹:<ko��)�Y�ќ��ʃ���c�
0�&�[��D��U��S�����a���f��EPz1�A2��	�z�l���,�}%@���淵���x���5���|���ba��S�e�So��͢u�0��:f�I���N�nf����މ��g�p��V��)b�9+��@�#��®�X�+���ۆ��Ǒ���\E��Gp���J��DDE���%Ϭ��b����@9��tL
Wl�;�uK0Q���-�ax�X�Y�d����ٌ�KWwD�Kʁ��^�ߞcd��֧���Z̒JMM��E��A�+�6rIl�~3dPg1��r�̉��q>�[�_�C%�sYܷ��f9p��6�F�����4����q�4�ʚ��L9��9�!i�\�nE�}IdkϢ�p�"X�i5Ϧd�&���A���,�kZ�%�"�sP*bIakN֘�,�Co-�/f\9�K�S4,9)�C4A��?�Ɋ
*ѣKG�V���\I,�)�wB�͡v��|�<�K��z��b9yO���1�l8��0nlcd�m���s-��O#,s�CDD9�bQ O�_pB8��A��R8�ITH����!����"	&\v�P�-Q"  EH��e2jSК$ԉ�bʕ�Q�L��FK��]@J4QMV�Fr��_ ��h�"7�R� 7�q67!6�hm��@�g��)2
�#�@�pL�ɜ(F Z�H��,�@��D#��������o{M�ZJ�L�6^�ȍTp#X���UU9��wf��>���T�'�c��,�ǩnא�}������g���`����J�S��R����/(� C�`+;��h�vu�j6�gY�ћ�-N�v^��kY5#��DɛWOR}R�l��٦�轘R�����V"�֖�Z�F�x�#���\���jm�/6�+�ʃِ#����fF�!�Q�ƿp������c�w)�����Q��A|=���+�'���k��J)Ǣ�JO7�n<_a�Zл����|�}_V�;x�KGٖ���N9һ�G�]��$�m��K=o�� y����;c��Tpپ����X�YOxS3X�K�@(��bu��py���M;�S��
%3���D�41u���+l�Y�W1A�p7�s�=PA�l�-����"EL�[Lb�Oy���rX��'#�-��+,��m���KӾ�]b���=�s�v��|�S�gO���O��ͷ��u��>�y� ��AÊV�91T�1V�kL��E�q┌~���p�����q��܅MF�d��G8Ѽ\t͗�������]��^���4�w=/Y�85�d���+��+�`�Rt>����4�u��=���>�mu�����O��Y�;��9
��߆:(��
�*1\��α{�W9|�H|�����y!�97#�,.�mH����wF���bo<�q;!���L�qgEٶ�ڼ�ۓ~��a��p�X:x�&��ΚJ!�J�3�ԓ/��4{bO�l��?DD^�n1��g}�1+ %�y'���:t�/����{�\al�Z<�Zz�ݯ=����V����!?x"z=INn����;��<��]��1�H�;a��ğ���e���X�g`�#Q�Ʃ���^M�%�����C�{6��t���U��Fv�ľ�AȪڻ��֚᳋�7^Sb�p�:� 2�S[��-5qEY��&�fqJb��û\�9W��1�Kx�*���0�η�h�}r����v��EN�Q]����2%h�htS&�l4���UT��_�QM~��.<5J�=]��,̮a�(��Wf�3���
:�J���)ׯ��D���5���/Pe%	��j�1X����֞TI�Gx��l�GD��Q��w�eN��-/c��ϫ�.k�K�)оP�^�MC�`|�kWl�|�z�*��2�S��4������Ln�Τ#�VF}ݔB*�8��6�07��z��ɺ�@��w�h��<,�*������ZR������l	�R�j�x���o!�f_.�F��y��'/�_Uwg���~҅#�t]�r�1|�b>�<�Z���WP�E��� �}~�T��]�.����70���s]F��u���jY����n����Vn̵Ǚ,Ь飫���oc�l\����1���h0�B�`��kǑ�y�:���ӂ75����I��ZG�(*��ތ�j�Q��n�0�h�M���_0�R��F���N�H�`L%��\I�"��;�B�*���3�֙��4gu�����@���U���N����Y��Xb��>�\yЌ���&�*,+][���ۥ�&�$M_�V�{P��d�,t�'˕���<���K�Gb}���]�\|��^�����rO��;��y�p9e�4"��3�Oe:�]�Y�yB�k���]��!uB�d̓;��:B���h�*�Kz���
��k��<��\*W��F��E��6��q��D���LN���]�����,�+�'l���}�p6��z���(��P�E˛W8�I�����/t�o/@��Ԉ���\����s^L�����42�m�_tg��T���5iXh�z:��r�<�Sȱ�Kmo^km����=�<4�m��Ϋ�z��
��s�w�Abc��fo��!��V��Н\k�b�籲��fx��/���2�4!__1�K�{��N��������ǳ��p��u�W^'��	�FM��ř끩1�)>���%���v��r\�z�����������[�l����ǲ�ʷ�7]E�6r9t�}����O���#�ϼ�`�Y7 7�G�h�?Q�$�W�K�53<�P�E�s犅m�cY�sQd�3��7�܎���(f��;�α��3��<c���{�] I��./����m��g�ˢ���bǳ|M@c���3�����>E��g�Y�R�m�5��lLL�yy��擎���\��5ے'��8�du�2�vR�
�<�ܘ�B�ʠA�����t�z"���ǜo�q�����D5�IJ����JN����@�OԻ{�위�z+��dJ�ԞxtvV؋�\�� x��o(�T�i`�B-��^���� �m��6����G�9Lx���=�1s����&��Ϡ�4R}vXE�;֒}՛��cq���/K���ix֚<���;d�%��X˽��Mkz��O9�ϩfg����}zM���{ʪ�w`�������$�u��}���c�Z�WW�w�l��T&4�� ���R��lI=�B�.�q{��35^R�"�Fv�?ei�Vr�|��7_n�8�t�k-���7RƠ;�ҷ��3�
�Z�M�:�p���\��Q��L�X���C1����RE��0Q�dl��`p�iJ8{�_M�ksS�p<��fs����[�#��u5JI�ٗ���o�M�ܽx��3�$w<\i���Y]���u/��;(#k�v.�$�-�c�\�"�>Z���@�����j�;frz'���u��w�Q�,�灰v�}Z���Br[�j��^!�1�]E
܋��u�y߱��,�e�p����I$��\k>�i75c!���\�q����kF/�Ǌ�cL��ǛwarH�h��0�5p��e:��4ߞ.$^솱hW5hWL���A�0j��bYKV�4K֭+�v�Dqf�1(�d��ی�.R7Q�ʻ�9�${b׹��GOEZ����y6o��,��w�ãc�2\�dÔo�o���udT7̥��̘�e��uY�^��GU�ޕ��p�'C;RI�(.\�<�g/2�r�32���m�p �H���T',d4Dd�b6Ƅ��n�!�BT4S�201�`�&C&H�L55U�&��$�M1��ܶ
8ӑ�#ޕ(�� �@3�@P�M�B��H�T�N��L`���BQ���@�n]o�N��6� �ʙ� �(�4� �MC cB��Z�e� V&�M��@��L5N���r��m411���	��14�i�	q�RR� �K�1$@��%u<*!
[@M�-��d���3�YQ蘳w1����h��~�Tސ#zި/�9�bofܽ�d�8�����ϙ�������8��퍙�-���q�T�����e�����x��M[C0�g��OE ����v�m�����P��b'"��,Trpi�L%�Tb���ٺ�[zZ#(uz�a�*0�A�y���{j�E9����k0�Y����{�	g�Ӿ��+ˬ���|��;��s����ǐO���t�͠�g(�K��g�&�zp�]ھ���� �6 ؖ�gPjc�0��:f``��bW.Qf�f>/9جڀ�`{Ը����	I9�����VrűKְ�ŋ���^�/e��C��9b�H�T�����{����l�.᳆�)h�lw�u��j�9�v���I��з�(�:qqfa���0%L�s��*�C/�ܰ�wb���U�tpie�&y(֥NE$��</QQ����Gg9/{�'����a��=4ّ0�K//V�_�c�l\ �`B��lQxy�㝼j�jf�-�� ���Q?����<��o�j��Fd\\��⨫�ϣ�����s�Pu+OC��ވob�O{����m���ŋ�R�F��F�e�	��K�P��W�>Y]Ƥ\/wBskE�	<��C�Vy���:^j2�}�(��`ůY���L��e�L:���|�Y�ΔWgx�rw�+!�,�8�����Y�@�u�F�yW�n��ܤ�i�k8l�b�EW:�A��S(�cb�O�=V�]EhM�p�z7����<n`���(F4��_��I��)ö�\)|�G�t���}��C���)n���݄`<t�+&G!j8I���S]d^�W�}%���Z�5v�n�5_���mM�~�!�	�Nnx����ղ����7&�����AC�L��X�����o�(��F�N�-dv-=�q�Z+(WU��2��C;��ffOk�=�@P��d�����d/��\{Ԏj�͞�a���^Y�6��K��}B�S��5n���� ������oa�f3�G+T21�fq�
��,�t%��\k��v�Y�����0ٓ�ﾡÉ�~���������$ұ��7^�1��nk����޻�����F��<�6�a��u|�8C�Z �L�w�*��!����u�Xe��wz�>yV_!T ��ّ��ᮟ�M(y��Ugb��nn'o�3	�IA�g+[�_�K���{�2���-a�<���<�CPa�y&7��0ꇗ`���U��Ob������k:�T�Xae-�������J��Q�'y͘�m٪Q�#��>�R�g\7��M��E�o��;M�kL�#�����G=��˄� �e��7��������ᢼF�3��6{W����s�/*�|7�{�@x��~�Z]��Fei%���^���.��z->�^o���S������&��RYFW`�[aFvx��§<����*o��׉�n���������������0���m���ֳD��''��pg4g����;)�m��%p�\���O�9G:uB,�l3�V�M�pFm�h�\e��ʶ���&��^g�["���?î�ɵ'�ª,�.����d��z=���-U����W��Ev�� ֩b��r��
`�(��f0(fX�m�����#�v{m�T�5�H��vbܑ�'���da1���Ӯ�[�b��
W��3��&�{S]`��}f`�G�N����ۡ���U���N`
�TM���FG�C������.k�#H,�2��{0mr[!�&����}��Π��ut�9 Ų,u�Qp�8�rs��,�L���~�2�;nG0��,_����_���)Ӯ�2#�Q���7Ʊ��S�xM'���P� &l!���J.����
F.3{۱�u���æ�C�w�hW4��5�K�.����	���6�tK��Y"a�ʝݕ��X�1�崼��u��:�߈~���Щh�j�\\c1��hqiv^ŗ��i�۹�����*̜V1�ͽҮX誨��8ܔ��x���Z�Vr�4	-�٘V^t9�3-�Yd.ԏ}ჷ_~�����!���Bye?�h���$J9��}�n�w�3�.K�k	��,��v�ѐ�Ru}OWp�<�#�c�O�ÁOj5,�{�-'fo�]څ8����,�wta��T�pzg�����i�j5Ţzfޛն�>��%��z�ͼ����AiF�C��@),�8k�ʅ
�LF��F~��"��^��}7eӨ�J�Z�a�F\�k.�A*V��+#��MVj�y0@�7��V'<|ؓ��P�I����3����9�T�����lm�d/�d�K���MZp��j���.��ˡV�"8���S
f�!��]j,.ؠ�qv�l���DXݮ���T���=\[���=Y4��yY�/Ii�U�{lwY<�ܙ鴤����9٧��d	�ޢ̢2�5�b�1��g ��<��\�W��q�J�-c�b2���� &nT���ջ̧�I����7��MW	���{�:�K�D�����^�8=�b�d4˘;1@����#�g��s"]G�!B��T.����c���n�*�M�[Q����^��r{�{;u�9��ϤU����զN�׮zgx�J����T�d�{7�.���-���^�#�^zp{��ެ�]\j鈔���5��E�*�x���x/[w�*���ץ�.}�Czm]77WP6<A�C�l�ʘsq�Î�g��;���v�*�P)V�:����[:�Vd:�n��uË5/&�=|\�[8�T��u�.���QGK������Q�$�I$�r���2�i IL9�L&��y��Mz7m�:Nt�y�,ͮX�DsOTo�V�m}�������;v����]�zd#�����9�;�vY*�����G�.�_I�4�Ĝ������s2uO�G�s�P�*���Ytl�!ѡ-�.�����.�i���G'<lX���R�I]�gt���3'1��MrWex�B�]�d�Fs�B)����r�䣉ӝ]\:��$�p�R���)&�n��\��l�+����X��دv�M}Qb�W���ZP���s|�I5qt֘�GM90I p��*ki��o�u_�2Z�R&� �Zp�>RR�!�6)n�E8`C"�PƛjZhvE�pP��J4 ��cT� �4�H�T�"A
Z���B�7 G1ɳJ�� ��	T���̥Md�JnЙ"L@ �4"[A��jI�L���H�$��U"\C  ����$#�L\   p��b@
���q����! �"�.K�Z\ $�s)@�g%28�!p\ 4t�u��;!).�-T�H(�� I��M�1��$1 ����#"�je��)@!Y	�!*f�*7p�1Vb����5Vs����:*�Z��ﾭ���ݗğ�,���KN�'���.fN����,y�{��f�+i�m�2�6�b��~[�X�^��	H���oLuCW3
�o�[5ePi��l.�@F� ��� ��ܼl�J�d��ܓ��'�������M���t��R⪶8	�5��{���{���ռ)�D���[\��+EgL��=\Tv��^���9F1���Ol'j=��nY��������S�yJG�3%�x��l�\N.r�k�pq�ck�w���^ύG��G��O��Ak9���|����F��L%��f}ٔW�����K׏���~G��/\7w��d��o�M��Qf��}	-���W��-�k����U�챇��i`& >��'rC^+���V����iXe�
{nF�yBZ�/x�����ފ��Ǐ1�GT����sg]�e�'B�7�cem�b����3�Oj�0�uݖ�{ptU�u�� �n1�,#2br�
�F73�"ʓ������?�����{��am.�S<�{�<�c������Y�ӳ6s�g&���b�B�ȸ�[ŏrS����Ԯ
�9�N�4��� ��Y�k���[���">^/>Dm:��:��D/�ٹ�=����GynƏu�����w�ߎ��س�H������ľ�5R���.��ɳ:�f%Y�상�nf�nn[գ(���f�F��I�}�9q�������)r�d����ۀ����X;ǃP�]wU�wR��=x0�c������3��ݔ�����/i#����Z��􎑮���7�a��G�'{2�"���k�d���آ!�G�n��^ۊ�Dg3�mcڅR3cnTa�p6���mtje��2����S��9���4�:+�];����*=��3n�_��ip���d���3�-�-$�a÷�ս7�y����d�2	����`
.���%��3�/}��;'{���~��Y���!�BwX��31����qT;���홥�'��s�/�r�]ē��J���?�9��7�p��b�vck�������Qf����&A�����TdH5����&���p���6�e�0GG��[�.E�=�x�
�+�<L.��.�S����-�2���zw�c�qֆ�J��v)l+���jř�;�f1U*a��;��F��0�������*}�l���u=Ù���f1:�c�ͥ`VU����īo��uu�C�q<�|MdK"�XIu�j�ō�[�3s�������n8�J@?}�p��3��s>�rj�':��8�ϰ���K}|]U��Ü>���kr�
�V����X���1��ݚ)��y�䜪�:����;Zy�����==�#2k��Z�_���ޫ{�������(u��yalɗ��}��=M�Z��!LZ��VA��nYZ���W����L��5L.5=}�ڃ7�⶝>��P�:��=���S/�:�jy��u�Dd�!G��Y1�Ζ%D0'�5P[��p���9
J=��$���\Y'�E�Ծ�a�}�s����k$n���M�h�W�Kd�A5�ѷuZ�>�V��(ŝ��6m����.9�{Vv4n�[���N#�}4��C�D�3Ή���n�<Kyª��`ؽ5kUN�\Yo�s�,�h���%���Y݌]�2��kR�E�	��:�ۨ��)`�4�N����gu� :�Ǣ��F2�Qxz�DP:8EU�USIa�wlʨ��K�M�o���Ch��ۆp0�(���jT���?U.$���{|O#�M���p���۬��_�,h�􁼪����4�r|h��2ޟh1e��)ئO�vM<�ep�S����+�!&@מ�7�M���<5>2�I�L��:u�ϗ��V#�⸝D��a��̗�`��5w.o�0R	P���O�J�Ǘ^U�G�*�-�_��^���vߍ�vjӔ�{g.y;�_=ƴWp]����S�K���F��L��IX���30��1l�����6�e+��H���ܱ����f֭�X0��P��{|���1'�j��2��εX:��4-WIn�;CĖn[�[�Ҫv|�TL�����`�X�}�)�6��7���zʷX�TD0�]����x���K�t�,�w��z7�,�����k���A�#ݵ�h�!�æLGKz�Ί\o^n���gwn2߱;�YT

��]p6��j(�S�93�\��t0İ����M�VGt�(�vzIL�0��WBgkԏ&z�$�H��U��7�B{�L2s�Ge���]�U(�Uᴒ���CZb�V�#*��H��t�|�~��V�����x����h3���8��uF�rѲ�t��Z��p����}z���x�"sص�Fnq��za{�I�G�ҵ��7�:��v֊�9�<˚D>�es�r�.l>��i�`�{��<���Λ�*��-�oY���}@W�I:*T$		$�ZU""(�Q��A~_X��G���d���P���֫�-����s_��*uv� (@TP*(��PUB���6�!E�QmQ��)�3���C�7�u�0������m~���Bnx~u����'Hy����*�W�,y�ס��k�Z�j����)_~���$�#�T}���i����������_��3���=�(�?��2*�����)l{N��\������?��~~�(��[�������0>����{�""��u~e���$����K �6 e�4��jxA��b~��h�_��Z���B<<�|���#��.zX}�f��A�?�����3x�1o�W���	uQ� ~�'��v2�H�+��F�o�����~YC��|��""�s�3�Q��7g�~��?jҏ"~�Jv���ܮ:<.!������~�)�������?Ύ���""(������!���>�?�g�w�vr^����՞T�(t���k���3��W�I�<D�?�}���|���y����~����"(���ǟ�����l���ć��s�А����QQ���G�?[� Cp��@=(*�V�>�\>c�� P!�`O�;�(����i$#�l؞��!�4���.
C�����C ����ͪT)!��*a�K!���؀U&�c���~�ꈊ;l?O��>P�O0DE���q�������?e�:9�;���@~��������;^���� X�'���k��D��T��	o���h��P""����8�<g�'�J��}>?�8I�"(���?H���C�7��������;> ���Ǒ2a4A�$�J��{��c�Z{+Ӻ�����Ϡ ����g��,i�#�c��^�"(�}`y��ߴy���u{.e8!��Q��w�<��x{Q�^k˃tJ�(}=��(�?����`��<���3�׫�ނ���C���ޑr����r8�24�Lj�U�}�� w��?�=:�^.��rE8P��c��