BZh91AY&SY�9��٨߀@q���"� ����bC��      >�&���h�dђ���d�M�Vլ��F�"�kZ%�m5�U34�J+MUSXU�S@͚hkF֭�B��iJ�j��*^��y55�L�m�k
���6�ى��SMƵ�*Ķʖ�J٤!B�hƉU3fʓkD�j,�%-�	U��%RT�Cd��b�taSm�kS��UK��m�F9�Smi�c��j�T���K[m"ئF���
���"Т�KZ��6e���X�S4�ڍ���W*Q�KV�l �   NC�Phe�m���83:
��aʨR�36�U6��uku�U�S4�wj�b�ʻ���V�;]u��2�ۦ���B��v�l��AR�  �|�������H�{i�μ�t�����׃�))Zj�*�ly���-�.zW=z�n<}�})�I��y��SM{n��N=)������-�il�������fo  v'��o�:[+ool���(:�q�<�Ʋg�Z�ޟT�}8Wz�����>�w)���QU�/��=��g٤�����)[ۻǯ�>}�J���|�އ�E��n�UW�����*��Z�+b�� T��J���}���QM}�K����kR$�y����Y�m�;�l��OZU�����t6�{֗u�p��^=���ס��s��ٜ����6Ĵ���2H��ڂ��Q[VU�  �K�BP�m��M��SM�s۽+�RM�����iI����{iG���+U��4���KM]x�����j����/V�h*��V��je��k�E��Ulh���E� ��t�*+{�n��=#m�'p�w�EkݜL�gWf�D��T�zҥSЏzv���w$��
�*�[��{�=5Jn����کK{�罌���v�sն+�fJl*�jma�  j��i�����x��-�!��]��W����3���U���z���A��8 z{�pttwJ㮃^��^�����U�C�ǥk+m5�Т����   =�o�R����=(ѥ�������y\��^��;��(7�W� 
�ޭ� z�W���'��y@ �OsJ����ى�%�M��k*DSm7�  ���Ѿ���QǼ�A�z���� �Nq{��Z��X� �n^�`�Gz�hG�� O{���z/^j��R��6�i3,b6�O�  	��vƍ;  ��� sOp���Jc@z�sR��z(��Gi���= qѶhj�=��       P50T�J@�@h @�{!�R��     O&!I*T h4 �  j��@��j�4     S�=UT�� �h  %"J#IOe0M2OPhh��GꙢ?������+_��Z�o�v�:Ȭ�YQ�Ӣv��fXz�L�c�����{������~��VAS� {���fTUE�;���3���?�����**������UQ_�T�)P�g���_��^�`�,3	��fS2��̎e39���f09�̮`̳!��f0���a3!�d3!�L�fC0��&d3���f2�̆`3	�L�f0�f0��&a3��fC2���L�d3	�&��2�̆i��&d3	�L�f09��L���&a3)��fS2���fBe3)�L�fS0�����L�fS29��	�ـ�s��f0��̆d3�0!�L�fC2�2�̆`3�d3	��f0�0�0�0L�0�0�2�̹�̆`f�*�`�"��2�fL�)�s.dRdS0 �Lȃ�s
aQ̠9�0�L��s*�e̊��2��Pȣ�s*9�I�0 �P�#�@s"�a� 3	�Ts�e̠��G2�� ����0�� ��U3
aD̊9�0�DL�3(&a̢9�W0��P\���@�fQ�0�\��Ts*�`�0�fT\Ȁf2�Uȋ�As�U&�Ts.`�"9�2 �eE� ��W0��E\ʋ�A���	�0��+�As(.eQ�"9�2ʫ�DȀfLȃ�3
�aL�a�̦a3!�L˘L�f2�̓9�̆d3��f0��`&̆d3!��f0�̦`s#�L�f2��&e3.bd3)�L�fC2��&a3	6`s#�L��09��`&3)�L�0�S2��&d31�L�fS2��&`3!��ff2�2�̆e̦`s$�(?�}w��Ǩ?��^����y�]��<��ؙO�����4PJnܒі%R[q�xsu-Ձ�X6X�lQZl�tl��j�:Fw�\H�����Wo�7�1�Ų
�n�º�&���ۆz+�fG��r��m�{$�͂Lu����;��� c@&��2,��^"tm�%����Ztb�J��l��L��j�`��2�T̚��R�܍��'fC��kí���m^�,�f˙l�T"�#����#K��n��J�e6��fm깩CxƗ�ui�/U˼����LT�.��V�ī7q9��<�B�2Z�U�E�nP���5-ɍn���X�z2�8ő�+Y*ˬ��r�����:�zi�ڴ���/bӃҷsd�Z�Y��r)�����`���n��[{���V�Wi�L�j|�ӱ�ͳ}�Q<�q�wJ^��J&�b�o^��5g+\v�V�!,�[V½�XoPUc2�:u!��nEO
T�fn��t�֊�2��`,���ML�"PS��X�3�hf0�8���l�kf�z�k�'�VӫBionSte�����̙�5S���.�0��;{t����6�ۨ76��q�8��o#�C�col^��]����6feB\#K��j�&�!(ssi�H�J�;ƥ��K9&k/7z��0��t���-GY�TV���"ʷ2ń�DC�o^P*�[C-���������j���1�j��&�@ф^b(n�ѳ5�VF�t0�)噠�vb^�J�QL��<�RU7~s�бH��Y��'����X
��v%�[�eZ\EZ�[x
n��)�5u�:$�bW��`��E�B[P^^�S�����M�����a�fK�B^�ә�	��AORK,�Zܧ���T�,�5ٙA���uiܺdG�q�DLĶ�w�S�03*#^6h����)��$˽���Z�M81a�Fsmˣwa�(�rT4^��Z2�w0���P�T��[c]�SA�/e\M<��/`q4��Ih��]�DnOX�"�� ��(���XLWGr�:&�2�,�2��+h%r��1aÌm^cRZ�S�/:�r�Z:q�Y��,���K�2��9P)YZ��Yt����z�;��j4����R;�Kɬh�%SVm4[YJ��mR�if*�R��f�I�Fo\+$2�-p�F�3�K*,7���6�f^�w"���t�Yt����\v��b��c-�61M�C��ݽ����e�)��1��;,;".Y����M
�/v���f�#^ᕬz�����`XrF�n2�9܎�(TCX5����G[��ıw-�3f�����Q������hP��vj��rn����
ga'���
Re
L��}�m��O	q
�!*�࢕^�hb�y��i����}��Yh�0��5��!v����"�d=������1��N蛭�:����]��$��<��6���4�n�I=����U)�f�8��s]��J�A�^N�͙0�(�^�k͑j �Y�ա�Y��ͽ3uY�srF���&A�mob�h�E�-�X��n�[�fZ��(T/6�v@���Ŋ�"�f��f�-%1��z��WGT*`ai:���BS�2�+F�MK��=�1`�o+�Z��j�jm��SBL	L��GD]��f�iY�܇m�
'�bl�׮M����	S&♊nb�Ÿ�DB;rV%2͆�"Bk��+��Ѳ��� ��gjl�A�C�Y�j�KӍ��aQ�{�(�Y��y�f�B�!�:���r��gi�x�h��%�U�:�kwDˉT8�ؙ�l�U��c1cݽ"�ݦM��'��-n�,Vͥ[bh|F��X�}���	*������^K�0bܰ�3��,6
���QK�����GV�}C��Ehe�|�M����5X��4o&n7�%4���o^�&7<�&�
�������{�[�ê#1$+#�63&ӃoF�kF��6��`�{J(�Et�ZI���VW ƭ`j��jug{l椵.k��L��,�YEIQ]��1 Ĭ�X�-���W�"IG�Pze�a�,,�ZvH�%�����h]c3(�ڦ�Z��`�ʶ�{�;��+���b�����u�C+&cyImhZ ��g�=�ܲ�n��Ch�-eՋ�.���Yw�C��4[�� ����d���QÏ
X��Sz�nբ\�SFY{d:b�ˠ��k6BͰ���bT�5��˦Ƽ�L��K6U��k�eHU
�%���U-�Xt%1s*&�K��h�ttPzʱt�lO*�-h&�m�y�k��D�iWl�Q��a����ݙZ����C:��1r�땸m��Xk[e-���	5l��Ò��ڗ�[%Q���&&���v�䩷.����+C݂A�E��t���)R�=�"���Ւ�����5��ű;��[�QVc�Q	ZB+��vn�oo_F��w�o=�.����[��\ �r�`ҩ��\N��:��X\��c�,y�Ă
Je9�t������M��B���ѹ6^d��f����KUĕ*��9���*wy��R*٥��t�5�.��6cEY܇(���ʠ��mQ����΍Fc̷[n�LJ�j����m���S�-�Q�EP�᧔�Î��]�lYyX��y6���hG]˿,�˫��̵[�`�1�\L�]iv���!b��i�b΂��h�q��%Qo]-
��{lվh �}�gX+ @4�"��ף����7��@��	A��V�����O�̮C�*8Z���ݧM����ݾ��\�D7�O$m[��8��1w��"`ջ�4��S[$�u�223Q����4éf`7IK`MUu"5,�۬����[$��z�Wϳ9���t��5Q��uɲIX2���*�u�6�:F)��\\�}ʱ�U]ԛ�LM��P�Qy���zbճn�?F�R��R3)��j6��&�h����ڎ�-e����Xfl
����,��%��82j*D+^TkN�C5m� �z�1����F`�r�`�1X���[e��M�1�&��zd��Sp�T
�V�Od55�z�NַԷ���E>��6��o[��,�lE�ܚ6ء]L��ݧ��7�3{l��Z5Y)�[�����J�Q�yX��q�,d;cv�I�.�@ɒ�Ƶ�����H����ֻ�pǩ%�B:������2�D��Q��s��c��T��n<�b�k.�/s��Ypeլ�b>���.�`n�(u�#So���*b��L�-D�2ֺ��b2�1����hQ�D�#��xsN�ҷ��1��]�J�1����&���F9��{���T�"��nU��;�37?G3�l��0T۫�;ю�fVLC�T,�W�m��RJm��8�49�/)E���&SI��n��`ǚB�NY8ӓ7/-�U�9�Gh��;f�����&'�j����n�=t��X�b�o,�;�BMF�7���p1�6��oE^e��-<4e5�z�fٛx1<�5�^ͨ�`���&�e��M=��D�	vf�u��q��<Y��0ފ��~(-�Ho`�ĺ�u�۬կv���:ׯO ӼH<*�.O)�K�h�t�a���WZ�^�6&�v��$�5� �n�Xr0JYl����d�^�l��8e�#�d˧	���;���6�ɷin�̢�mlbk����0�71n��8�-2�a;�+8���%e�`o ���y���q�����o@xд[��V��W���L��YAa�SɛX^�k�e�2�K����3rQ�Ԋ���/j�L�܈b����p�ч	^[{j�ⅷH� �̡6��B��YNZ�!S{�m���ؤ��i��jġ�fBk"�6��y����wZ*^��9O$e�L<(�V:��ŎM~R�y��A���6\�sM]��jS�dIi3�Y��y��˹F���*�b�Fj�"f�
��mm=�l)ԛ5A0��5f�y�#R��D@L�;4�,��h6Aţ`���&B��<)�t��˂U6�6�Or�Vf^�X4N��^�9����	v���M5�IP����D׼5��f�׺�����[��(!�����S����)I��$	C�-ܴ૊�T�mA��9yx��ThM�H�X�+,�E�ժ�gf�k ^�L600��e�գeH�dQ@��nfS���Zt�JflyT���7D*�wn�r�Z]�ҫQ���B�]T�u�ȒS&f�MF�e�Y�Y6�Q���t��1�m+-l�'6f�sB��ѷ�v5�)�X�b�����ݭ��P����m'�C�}{�j7p��Pu�2OE�b���|�l�y��wO o�k-�ٮu��ʵe1��`��ܑ���b�`+U��%����OSf��
���w��qpJ�k/�8�X
l���K�(�B�J�%e*bð�ZS�e�b�یV���h9�ZPږ�n�Z�v�V�U�r��kx[٣q�Ӕ�yf�[T	dAym���ն#�^1u���v�:�V��V�cj'�
v�8m������b�+D��`أJ�o5V�ȞZ�*[-���E�NA�l�d��=t�hܫ��	���X��ޙ07�-bش��ڼ�Z�^��K[o_�1��M��A�e�U�R �',źIZN�R"��˛(���7&;�t�ێ�;�a"HP���Y�k�3kQ�m-oH�Z�O��:�h�h�pc̩���3[�vi��'2��cM<��c��F\V5�tF2Yd݃�$ku�k@��O�T�rm\&�Sq��j���n�ܸ6��#�;F�]j��*��Oc��c�H��kcOr�n`v	��w�Pg"�P�^�L�Srݽ���D��QcYf�2b&c�vR�LЌb��H&R',hj�y�Og����=Q�d&R/p��sK�6���=���35�t�qYє��Z���H��2쑸��l�ٲ�y̊�ǊZ�����Y�z�/r�)pi�yc4�VE�jV�%鼤����S$n+v�J7~ǘ��H2W�+���Z�\�5ٱ3&��J!=ۍ��j����^T�"�H�i]��̑#y��fG��n딷[�<g]�Vu�X�6m�H7sV����C�,� {R��L�!��u����m�n�6*X��˼��\4P�n��0��E�K���=�|i�+Ay��������ⴜ���hXSX�)!b�Gk3m��e;��K̹6�Y#ҵ�&��p�dӽ��1�OQ@��E�EգMR�!�03,O�SK�eӠV����-Ŵeh#zý7�u��V�Ee	�)/�^����2�i�bD�䔝��*���l��sU�=��
�&B�z�gMh��4���j�-a�3TZ��ژSNDfi�Sb8�r�/S�g0<���Z�J떳���l���F��A�6 D�;#nֻv��,`��WKc��;��M�A��7B�*��q檇hhVk,S��`�`#\�E��6��F��� Y�\�����Y��ud��U7�yI0C�-JJfx�~���0��(�4h���Ց[u��E\q�#�7˅�x��Xw���U��dp�C�2��:��cY.���h��K���8,T9�X0nR�������F��\Wqu������;���al���֕E��]���{�b��,D����n\�52T�h�E"�t-�hce��u�k�LV�dxk-���(�c5zh@sJG�kX{�cyk��ճ��<�8��
%�hj�{x68�	Q���]D`8�e�X˙��v�)��P�C��>`	z�a�)֚WKj��8��&��!gF�h�"	�Njծ���3kO6'+���(�i�N�!���q��u�f�~9X72�ͧ�l�M1ʀ�'L;kHSB�ҁ�jx�t�`����aۓLrFf����b�Z�s���Qj^zH�2��2�bN����*dvqXY����k6�k��8�faVb���iQf�q�{��SժZa��d�A3ZV^�������5�R�A�Wfn��-]�!�U���)oKش��4����wZ�+/3[ݐH�ɰ���G7dTz7K�ݲ�,��(������J�,	�{��zIx�pf�*���b��N��^�:�Q��sTOD0Cּd��mm�ֶ�%���`^н����7姸�<X��\��&^!�V�v������oS`P�x1c i�܃��*�7�e��	f�0��l��F��[X.k�0�Y�Y��`Zoq��ԁd������FM�	ۤ�r)���VH���-�.l� ���Ee���.�IL<��p�F��u�c(�ˇ%J�eiuжnhO	���:@��z2P0m��$Q���sԆ�9Rg+q,�Wf�A�ǚ�,�kh�jKEKL�76�`ǬL��H//�G�h�XЃ�e��qu��1Iٮ	������&>ރ%C�G^��x�V��Z�#�/�&b�&�M{��^���]h��F��E�����_���Y���`��p &W`2y�fa(u���R&�Vn)@�M�����4��wl꠨��p|.@���A;$ȳ�L��"^F��yX�f� վwM���B��ƀن�}���#�ۤ�t�WW�s�a�.�Gh.-��ꈮ%"0�d�ļ6)��k�iD�/I�ːes�m�2��ڸ�#8e\��8@�P�8���8LH�(�P�#��Lpl;6�t䄳�a$VBFuG�jt�c�o[&17�3�Nla�{(kX�{7+"s�l~�޷�p!��һ��P�#)-�ǆ� y�g��I������|	�(C�.��_�ʼax#���MgåN���RYZ��z���"���=.���<�r�M(��1����C�b�V��xM��!d�8M��Y�B����+�Qj�"����q�}Z��N�:0�oH#���uǠv*fn�ҴR�[��-V$uZ��H�>�����7���/�����y�߿G�¦����8TL��өrA�����Z"S���+��Zvq*�8n�.Br����%��b���wZ�
i�;*�-�^�*���k�,ݷt���v"��I���8#ǜ�ECc��	��!Ъdķ�=�BШ��Aҷ�Ufˬ�A���MC-�;ý��4��� �7�<�����d�-K�b��Ӓ�0Kl^p���N�#R���3��n�|k�j{ȍ����[�@YO����ז��;m� /�u_uF�Uӣ������"�Q�1nR[��{b�P�`�\6m�s����aԯW0�k9�I��B�S�Li�9bk
��l����%̂ɏ��|��[�3qu�d�#x�V�̏��m%����m�<k��rw
kZu��\r�t*�P�qś���"�M��7]�;��qҕ�pm��t�$�iD��Xw�x�v�<���{';d��MX�AE�/F�͝��G�6*�Uh�ѫ���,W+3��[��m�y
�F'�	�հԖ�&�QU�h۳�8*���������p��o��r4.U��|���q�=�;�=/�Ө���O�f��R���]���Uӹ<�U���wvs��)�5�
4�{��[����� �/%oHieq7��l�U�eoGvo�:G��	*�,�q�Z#/
����!�݉���kں�fa�r��;.t�9&��<
N֪Π���Õ'K���r��T5�z���$�,=//�o��M'Ѧ�J���enYS���F+�TV1]G��Đ�J.���!E�nZy�w�a����]����v���-�ge[�i�s;f��( 7IK��"�#�4b�vl��H<����w:��۴[��z�Tʁ�
��3s�6u`=���8ս��6��+rb2�_mL���,}-ta�̺��b󂮻��[�/P5%���R�s�;��\�ǣvNU���F�yr�7n�h}s��3-jt�L:�"�Mt����e�[��w�Nne�냎�d�T�,���V�v��c�g	+%=�-���8ө�p�8X;R��F�8/rgV�b���6�̬:Jo���V�ns�MZnbT������A����|Vx
���M
�M��k����j;u����Z�ݸ��,�.u�������Zr�]�f]��6��u4�P�wu���i^��o<����)�˵�X=Ϭ6�"�_m�����+K��vNE��m�  �շ�`�9��Tϸs-C�=n�%�9q����^�t5]�yŹ�V7y���ۥk&��gf<9 �[�]�M�CTH�*�j;
�]���os)�@o7m�XOLys@�"T��Y.���-g��Y�;����֔�GU��`�ϯ�ʎ%�������q�x?'���d%w�&��YW��\t<�&ZW��i�c�y�6�]��r+o4)��Z�u��WR<b��u��c��ȩz77���q�Na,�!����K
`��-�,�g�00t�p��7/{y�²�!!�r�G�M]�7[�w9Nr'��hn�[�7�i�m���{���Q#��WV�D��_��rV���lK�9���YH���� �|�^���/wZV-�M#�j��}���dY$$�q*�y=+'+Y����w�VC��.��E�� z1:VZ��h�uj�q�K �|�.�9��9[�0&�(��U�YZ6T�7�W��6:�M���2N�)p0K��ţ��؄�L���]{���V>�d��tM�d{�,�PƝ�̓^'�')efMKy��so��7v쾱2��`����}��l��*��M�)8��V<��}"�|[��^����o�Q�U���:��ɕ�mMw�i�"d��^A���������/7T�)2���_V��[
��8���c�� �Oeh8u�`���o]v���:�ΏL�Q�u��n\�q<���4��C�A\V��a�Ep�cX��gK8���o^}��ڊ�rH�� �b���P��t;��5#�[���ڴhJ�m3����U����Q;ZF���������\\{C�;���+�Ơ/7�������Q�494��ݣ�-�sZw*�R��m�]9)���G&�`4j�B��U�,:,փ���;�Ovef�dƵ�I�j�9��B�<��]��@䩑N��s-X�Ȅ���X���	��Ո��'[(��;^`�\Yx-4����h6̼�{d��Cm��x#|��;���1l�u��× ���r�e�:�pn�ݐƴMԠ���]v{�{��R_Q�M����%����˂�M���kXk���b����E���/�C
��p4)�6����x�>�rN�����"G�31r���Y}�Z`U٫)GG�iQKI㔜��`�����Xm��J��%r\�����{���u���=��G�'�L��p�Q5���v]Gk$���`������T�"��!��H3lR2����Jp9���ՇH,]Ӛ²����h����ؗ{@-�TYu�"�{]V-�ضÕ76Whe������bݚ�o���߳'3�6ǅ���v���q�}�'EF��a@[�qVqb+����ӫ�&Լ�{Y�S� �5x �c��)��=��IƦ�i������mҮ.�os������m5�#����.ؾ�3����bV���'g<���U��K�\*�M*��^�4���5zPf;��l��WA�0^������QQ�j�v���380�z�d�'� s����-swu�������j�ge�(�)��w� ֤镙o%�͢4b��y�ڛ��g��w��w2	�]�P��nv	�n�:�ٺ%	�����Pt���ҵ^��drI�W],:�;ʖ6���̕ ]r,6,ioTxW_M���]ٛ�*�3G3���l/`)����f�=�w���ՠ�`7���Í:�;qEqo%����bv6`ҥ;����͎)'�'���*9��/K�F"��%*oDz/+{�D n�Gټ�$��i�Ҩ'opG��.��wvzqÇ�
��N,��Ve v+�����F-�*w4��|�a�DpԪ�6q�.��|�\#�u�d���� Ԇ�o��:�{���+��ۼc���SN x,�vL�x��@Sk+AzK�W�->���FlY���ez�EU΂g^��wWvK�0��%}`���.CIYD���T�+f6����r��9�n��O�@�s1kwk-P�F��,�˦x�y�pwP=�+�ƥ,�>6�hwSi�r���&�2f��(�y;�@��e;�2(��[�����\�Wr&�,e��D�Q3g�Њ��K6M�Y���Z���s��Z[{k��)Ւ(�qR�ȧ+5b�kV��7j��5����`�-Nz̭�ո�1T�#!�qǶ�>��t�F��ԛv�]\�q�'u<sȚ���
�����tH_gs�)��2_����o/P�oNE[l��f���oM�1q���'.�ڵ/nJ��1u���n��n{WG��&��U��^�e�^�7�� �����@��]��zS���	SrweA������4c�me)q�����+*V�2��qe�T{��b�k�!���R�eͷ��X�4�9�ӳ!��4�'�w��Z�\��[g�3Hk��'k�L"������=�[����Ŋ��	��s�����t�c�_6���#O[Zm룔Ȝ�ލO��v�����0�gce�(f��b�P�L��Q<6ܓ)���c��l��N�-t�}�y�5˶�s�N�v�������<���E�Įx�-m�s'�����s���
�|G��Y�H�6��w�M�)����Cy3��;�o{.�UǊN��J���;���u��Zl軻P����^���;N��Z�≼QY�wgztμCa���4�M	����GR�똀�s�Z`����3\��������Hq19�����c.�N���pۣU�~�)h$j�U�.�WWՅ�H����ͫ0���_o8��<�G��P�mv�o(�V��sa�8�5%7|�GW8zJ�X�]ڮ|U�,=Z�WMwX����٘Վa��ej��r��i�弅ъ�=��y�]����Dxإ�n�WZ:!�k�Ar^��;���
Q�U�؄<�ڸ�3-�!MK����z���?4��b�{�[�d����7\֚eA�c$��mWU�y�њ��fNSE�J�kq�@�-����#'o��IL���� }Eֈ�嬧�et�I��+���/�"D�Es�HORo��t�*�}Z+-к��O�����8�`�w38'��6�y]�<Dm�;��i�bR�5�_T��*ⴽ�������hn��(�ۧ�����L&�I�*3D��hK;#uu�_j�{����m�-��lf�V�ۼ�L�/Pu�h�I�J�ZX���I@���Ի��N3y�K,U֊��i�K�4;{ v���������.gR���[X�e[x�+F>����T���[���֥2 Y�bE#�ï�I;苃]mt��3
�XaZb����2��!;�3��o�̨�=�Q���$��e^<(��-�ۨ�Vo�>�ʌbI���@�s�[��-oz�$J�l��%"{4ЪCd���f��L�����qV����ΐ���;Yy�ng&�_]	�;��t/��������.�8�&���ubg����-N��<�ܒ��r�drV�g	�TkSp��"����&p�2�7�ʒ3]��udQ��d����h�o��][�I���w��E����|��¬؜���Ҧ�8���r�ZQA��m�5������[S%�{k��<�vl��!��-����̔�7�՜j�o΃;��T�G��ԕ����K���hy+�Nv�����3a�n8r���b���6Џt�wq����gZ�����5iUݛ8u�(0Y�!W���k�,�W�(��mԑro�4�gD�ٙ�v�P�k�m�w�t��kr���Է�C���zOc&;����p
vk0��5�F�/�����՝[�Ҵb����ؕ�P�͍��L���g.��O�Dk��iVs�u*���GW�{r��B����?/,񮛆|(i��V��*�6�=�J`�S.��A����)0��x�g�et�ʧ0�vj<��Hj����Xx�+�+X����Jē��:I^w6�q�5!�KL�'Iڻ�W�(Ft��e����4��u�)Xk4��f��`�D���]×v,|a�u=jjP �K�=\���kz+���Ց�R�=��-���Y�ۜw:��t{�ք:�)ѩ\�(���&un[��O�ʩ��Y�霕���r!>\�T�lqi+K ݇0�ޝh�T(�ԕl������\N�h��ݗi�d\:]t�6�6m�:v��[�B�(+di��.��G�o`�LOT�Y!���VMb�.ٔ�i���ͤ(읷�ޗ��-sVV�
ҭ�z';�BM��,�7R��&.<�:vp� �o!�n��B��w�W�tθ��,^CH�:����5a�#*��jk#|�ƶ���6� ��G9{����G؍P�6��]��tD��E�(�kjh� �N���Ƞ���Hs��چ��рT��2ͪ;l�Ǉ�� ��0fJ��VX������w"��]�:�̝���9]*�mKi[���`3�L�v��6����^��@m9B���w������x��A�m�䷻�M���ʋ��<s�ue`�}>.�b���$�S���Z�����D��~�2��X�Z��RS,�;�j�#f8�$G]t�G���B�S���5�7f��Tᶀ�h�<�]����C]�=���Pe�9]G����u�wQN��ls�r:eL��j�u�]ʔ]G��N�u�^�N�u�����wz����7����n�K6���g����o��ߎ��J%�r�"j%Ƿ�����B��P�W�s@˩�k��=}Y�
��7i�����^�[+����.�n^@�1S�⬼����0k퐛�!�f�����7�GYѵ��{�l�E�e̷\/]ڍ2F��l0��5Rr�8r���]r{�E��[�X�/7�xd�hSb���ͺQ����\Ia�7�]�|4�b*�5�+���˽�i�}���KT,���l"�V���F@þx�_<Ɖ��!r�K0�K{ y�ƙ�Mֻ+6�@�Y:Q�yCrj�e��BB�,I�W]{�)�c�Z2&F�uDT�9,�W�p��!).���j�G�MCJ���{��f�sV�bXyb[3��O��2&mmC8L�u�k�˂E%Ƴ'n,�������ˊ�eK���lU���Ky�U_Qc��1��Gt^K��ۺ�$*4�ܺ$2����=�G�k�D�O;���=k"�f�0�8��4{�����9LeiW"�S/�X8�	*�ʹ��/3�9"����S�&tSe����G����I$rI$�I$����E��$[��#��y��ab��g��#�����T��\=����ߪ�Tҫ� �6�k�T	��_�#@5U�z���]�a'�Ȳ��$$D@u��%��C#�+��1� ^sDƈ������\_'��N���/W�-'��O9����c篼�r{�М����]����gx�}���=]@}���o�� g #�+`b(~���^WeX�p
��VT��**��P����'�G��@����KL���J���"Q�������=pدJ�S/�ǰU���G/]�:�����:�Gv� E��S�/��� w�|������w�⢂��?��������_��~���z���W+��0o9��38R��p'��`]��Ѧ*m*�sq��n�GHV髗R�;�
va
SY|'˵���e��)kV���ʽ�.��f��oC���CD���9�R�&c}B��7D��;M}jTk�;��C��a�.b}O�#xy��-PΆ��3���̫���pY�z��\2X��˙b� ;��ܲ؄�OY�x�읟Sg)���n껂��fB���˸̌���Mc6�����@���!e�[p#k_\��°F�L��0�P�ˆ H�0neUޚ̭XS�Y.��&�J�����3N%)ʗ�n����@hw�����]�`5����&Q��C��|s�]����weXL��%@"7r�|��;�y�ުD웠W_���HW`d3/�tuW�a�T*�����ӡ6���X����!@(���C��'e�E��l�r'�����Z[Qm�j�Ep��a'_6P��FU�ܚ�iGV�c&�Kq��a���Xf>�E-ܵ��sa�.�tkAVs�G��^�]nU�ui�3w;���/�8��C@S:v��+�Ģ8�Ѣ��[�np՚��lW4�r�崹 ssB����Ch0�JK�Ջ���j��V��:��f^*�	1XY��7�2�&@Ό�Jih�8��s�tj<�}���ٗ�����}��w������������||s��������������������������������������>>>>>>>>?������}������|||}�>9��������������������������������������������������������������������������||g���w����{}�~նܝi()��%
u���(���#�czu+�{��Zz��uSW�e�h��&�������f\��v�k��p�3�+e5]�y�vݗ]oѻ8�q�X��T�*�4{�щK̼v��,ފF�]b��ݛ֫Ks3*�\���:���ft�फ�v�lj.��}S�p�p_u�hEu	�)gm�]%���n�_W;Z���}}ݖ+Y����r�Sp�/o�
��*$P+&��A�wn�5���n�Ꜵ^���Բ��t�%�K��H���WG��qșKF��j^�t�8jiX�g|�vԡʻh��)�������oW��!��:u��΂�T���S/��!,P����:۴%�Y�K�D�5
�O\���>[ٛ; kVEY~ySt�}��D��fJ�e�;��6AŖy5�fY
�1.�vNaٖ&�����.d���nu)kܞ(Ry�ܡ�Hʴc��n��{Ev:�[�ɽ
��\��W�o��l�g�N�d��˷��z@��LS�	ͤ��Bm�j=z��6���6%ײ���t/�/��K�v��_>NfNv�n�jv�Ҡ��s��cvsx�œQ�����O�Y�y|�t��;��`�!�)�	j���vk8����/?w�������y��ώ|||||||}�>3����������������||||||O���O���o�����x�}�>>>>�����������>>>>>>>>>�������������������������������������>>>>>>>>>?�����������������ǽ=��w��B�C'q�D���$�t��6m��k�Ů������z�k�KJA84]m܀��j��}�Mu��N<����l��5�oM��wD�C@���2&��E<Ȫ��`����iw<K{�]��p�ѺE�G�����r���V���+��J
븲���6K�Nrb�7gp"`{��U�j�S��=e\̗Gx�;�K6�E�Muoh���iV)��w;j�p@��z�t���K��3n����6��0x�)�բ[$q�KM�%��2�^�WwIB#ws�"m��!k�%#^�,��3�ݽt�`yy�M��cE��������V񆌝��9����E���f�Y�l%�^�^JO*�
����	�o���q#+m^G�D�^���Z5o�WΎ낟,�6��iJ'0 K˻%8è]2���J�W�;�@տK
�c�{���.��0.�w�B|l��[����}/o9��78�7��U���\̕"��J�*ë�����1]jp�
���.3#Ϋ�/0�jH_o`����}�k6�s3��B{�G�=8k�hn�4%ǜ��.G���h"�ҕ��I:�W�Wd��T���D7X��L�L�h�:u`�t+^Vc�ED62�]��ؼ�:
e�ѭ�VK7�Z���ou��)̺�ȊIq�d5�)p�v��T�M��ȇ��2�R��h�%�B��D���4�3]vj)�\��0�u$������]j��}�Q��K$w��++�烋=��%��R�^VR�V���N+�m�k[���ͫ�֐�-�+0���͸m.�)tzd���=��H���;�Q�y!<36�e
Y�l6S�g*>|��S��o��ZYW����ɣqi4��nN�
��;��Z�f��=�³"\+�ˮ��Y��y���h��6Zf�cm^�
�n"Q�Ɂ�������|�9�ZT��<���m��nAϥir�r�⭌�m`[��h���ؽUCr%˷-��s^�����՜zR*��ঋ�koZHW�I�gp�Q�/��TC��Z�יN�QH�7��Q�4D.���	U��u��f/C���ѢZn͎�O����&���W��9�u=����s&��ʫ��v*��Qy7oB��tq�\:��Ǽb�Ū��:4��Vъ��T�b|�.R�Y�+���(�"�#�I�Oj���9��Yג����2����&���݃F��ӓH�������Mju�K�6�.O�]�:�]�;�v)8����B�{7l^E+R��8�kR=���F�^�����5�pj�(��r�c�#Lg�ټ��z��-e"�f�XX�f�ۺ��%�ou���@n>����û�;�'	t9+��7���8�����U�;�1؀-�C��eǔ����z�QV�P��S)9�
ѥs�4��)YL흻׸����s@t�wR�x�VrYu���f�L1�9�5֝
�'Z�L�u��(M����s��.�!Z�N�T�s	��B�\�Lu�)��c��3��KU�&�Pw(cXd����0��n�k{(GQ���f�4��v�-T��RZs�U颥�Bw��]}:�w�c�mas�N�����u
�w�(nj2��d�qK�EC��+����wTT�b#2+�s�����ZT�t�$��4��kx%1,��x���%�Ȓ��v�KZ��;�7l�FC�V�وfB%��u좝�M��E�}6�VS'����~��j�W8�;:m�\ݙf���j����pLi<��p(�g�λ�AasΠ2.މ<��畲�N��֜N旙�7�%Z���F9+.�5Ī�{t�	�[R���K)��,�����^�֯HT���3qx�2��\mv��.;��m���\@T�鮹H��u:h���u�Njwr�U���>HX)ɢi��Ϡ�Z��l�Մf�T����X����`d%���3�|�t�L��(�Z�$�k&�ܗ�*��J[�c�x�-Wjjy�/�(L}a����˶�iJ{A�Ni:���,P5��Z��2'V��
ru�`6�C��{z�[���yl�i�(��4��&[�����7nM�;����㤥p���gca؀�:�D�S$���.��4��*=�*�ѳ�v0���8N7�a�$���9,i�%�Fq�ܖumv�(�_g4�'M�|��.�l�F�]�q`�7��M"���*�<����Kx�)M��F�*ޙ{����j�,Lr>�x���/M֓/Y�ʔR�zT�VNA�ը��w^$t��*���h:�Vu�-�8���`��U�Qiz�'< 
��lOv�`���7�1}xVsI�V=��m�Ə!�oF<��JR��r�S1V�������Ǵ���~��oU���#���oOi�2�8�ܡ��w�M#�I��}Ӗ�dl���z0PjE���XIk&:"�8M^�/]� ��n���˒1���fU����wrL�F�] �Y='nX�m]�W6(l�kY��_ɦE�Q#+m^tx�-<=ZQL�څ���W͒�hu1l�0�������N���`�H��Xv��e��-U��ƃ����[=�X�(81Ѽc[ޘ:�X��|hf�{�3�����z�!t��D�qbv��,�ƭ�쨫�{a�gV���R��lݝ#��~�rvX:L,N窠�QK:e㍺�x��R���"��["�tD�#䲶�WM*��A�]��\8�@Ha�佣���X��Βۻ��N�:m�ך����x&�]c�ײ��@:ʧL�Oq�����]�ǎSmv��w��f_*���*��[������ަ�m�3E��VgwRp;�%wBm�A��{|�.��:(��@��ӷ�' T�j�053.�C���NSWS����+�c������9��Z�6hȘ˩e��E�r v��r���v�1�Ç-�6ͬ�zq�$��e$�74i�9x���ɍ�&��qf)�,Q����W�9�N��5�u��i��.HY��[��eKr�'�qiLoZ�K��s�X�uX�Y��4$��4*�`���%etf����%2}Þ*�R���b�&��H��snZ��Q���(��X���\n�р 2�YY)�v�{\89Z<�E�n��)�5ȩ�nov)����3E��o&V�WrU-�F��0vի���p\�,c���{�n�g��q�ը�P=��
�M���%���v���He�����֏���(>7��kL���h�\e_�hM��kM�r���T��)�ss7 �e�u��%k�bx�>E�X��;�ɍSk��Y�����c��,-rY��R�.b��\"�����֢���JX�F�ge@�+ �놧k�#m�������5b��2�H:-�ק.�V4]4�B֝�W�*�`I ��1P��2���͐�׹�j�t�̜u��:SfԾ��6y$��n�չ*.��7����vwm�T8���9)�J�By�`�[�ՂU_'ƹc�HZK��������;H�mv��X}{/��19M]ڣ�6Zw7�^�����7Ocڔ��k��=���#��\��Q��oRt��h�ϧfm]>��.-�EL��)M�u���߮m�'����jh�:�e��tL��1U��6��}����fg;�z�
�q�������bq� 0�'LU7p�t�W��2\�{5^[�x�+�Ó�=�h�ׯu�˗��R��`F��LJ#f��V��ŜgV�I�X,����{{��L��\n�ە]fa�	ڔ7Bc��!ʱ]��D�ٙ�����/nIW��qm�E:�����$����R���9�WW�iz1�fؤĠ�p�r��^����S+k��刓3o,ʄ��P7Y�P�Nᮮ�J�3���������.�)�|�������c���N��TIԻG �s��:����Y�^�� �wuy�&��x0�f_�"��}��õt��䯄zKr,;����V�ט"�2�7��Q��o8�|���u�w+�.P�;N㾊)RgpU��m��.�_Rɬ�x���bƾ��<��|�hc;z�2�\:ȷ������P������c=Yg?�E��u��"�ʽ����8>�����:��$���Sh�-i�3c5u�cŦ���Zj�Nop�;��
AT$g�F��G
b��/�Ny�!�u&��}�Z�Ux���b�;Ƕ�d�-�3P`��]���כ��J`�P�i*�r���=U�cZu�0�me圼:�U䶫���˯,�{)��u(Z��
� �\�=��:��n�n�uk�m�v]���cF4�Y�,m8'b����Ói�����>]����yd8��&3]�1�A�,�iY�u!	�h�_�z�r�t�w��.��J�K��	{�"�P[��d� ��x"�v]�,1���ܚY�	�ڧ	�����QҥħV=-5=�!��kZ#�b}%H�w�-߯mmFX�	��[���j���풞K�.�IWMx�Ss ���.	���^�w�R/P���^2��V�T=&��z�[�h`�����I9��*o�7��B�K��3A��8�29C���Ut����MUq��W;ral��܉�ʜ�Yha�6{L� keR^��*U��vJi�-=���h&�Ug�p���Bt��w=`ާ����4��<Q����w�:s���)��@�.HJ�ǧ"��`����K9U���Z0^V���3m��` ��w3uB�����mv�[2d��Ǔ��+�x�'Ϩ���}%G�������Y�B���̭�wkRp�y�{���
kkbgZ����b��|�QY�˽/�����TR����s��k���K�qͩ�]�$��RVΘ�
�5f#�)����d�O\�Z�lQ7T6�Ul�԰��]��B$��JLn�ea��#ћ,mqe�zB�������8��u k�Nv59V��.Q<eܽ�%`[z��}�[v�����L��9�v1|�n�y�X"�ZIԈ:��B��2������"�Om�s�=t�}����4�T.�BE� F��k)�
��nL��,����qW�|빲ֳ۹ݳ:k�i$��5�+9���9���,�?�CL�'f�M�t3nf���&,�o����M�dc��ӕ�wJ+��\��sć��z))u��u|���J�����ν}̮�D�{wݭ�h��u��X��m�|�bf�$� �B�K*k�V���]�;�y/��*�&�#x/6�H+Z��A�'_P�eId�p������%j��.���M�v�ouBQ�:�d[M�۝R�@��T͍�t)N����5,��d�r�i����r�;Bv��efO3ܺ�{�!ҙQ�$���T��B�?\i�CW����Aux�Q����-|���]c�Q��6]��Z9t&b��o���Z�����^_٣���o��g��r�������&��ۏ��{�1�X���d��~e9#2H"��F��2�u-Ƨ�ء!~"2
���2ES4��)D��dT1���s~Tv�J�d+n(,$o�a4c���%Mb�ݻ-�d	�8Ag��;���>Y��|^UgB$��۽�F#y�d�,��?�pf�OlK$8q�V�����n��-н��u+�64p��0yvK�~\�6�KL�I)�y������:%g,�b��K{ɧs�6K��x;�-��k�6��j�"0b[u:7��a�D�2�-��>{�SI��;R�0�]�儯\�g� K\��r����h��;g�o��a}&j}�Tt������I#X�Lԍe<p��˫�����+#�)%�nB��[�W8�����n''!n�ő�9�Y�7c���b.�����G�A�=iqSEQ�!N�zb�B���cʶux#��5kWS�C��L��¶�pf!��U�S������Zr��H��ێ-xY�����H(�F~��wE׵�#��g��Dl�os��b�k=c�:"T���kt��'�Gr��hE���f��ݸ��IB�[�6�i�B��:X�x��k�<��[ژ�����Сy谹F�<�8P�
r�(t0�#��vK �X+F�t�غ'%&���-@��@pf�ص�i�έ<(��{Zp��JUȂ�02�哦��a?!ҁ��;��n�+�^�!	�����n���j�(�wv�l^e��'lOgsw2Q����k��uӶ��AN8Ç�,5��h�!���F�&8c(�$��r"P��UB�*"P.4Q,�AP$��c�Q�R�DAKE(���-GD��)��	�.8�D)�b��FM@�����(dQ��-�M0�� ��L�YF���e�&6��N�kʣ��
�Cq�$"bA��6Xl�Ie6�rm��AI�����$	�AW[TEQUE5�hd����"�������:Ω:~=�>�������}��o��||�(�*"����("��j+�肻�IQS|ƚZ"'Ƿ������}��o�����Ϗ�MPZ��$���*��<���6�����*�()��������I:�L�UQIPMTA�`(bH`��*���"()��b���5QId��˛Q�뉤��*�
�`�&��������ʹ��A|�&Z���&�����Qu�Wv?-�=�ԗ�w��B�6�f6�<��u��ӁlUP\ξn�%���5ͪ��q��U��)��9�_|��u�`��>s7Q�;��m\�W�:�q5Om*_{TKnV)ֱ�Dy�\�6��cZ-!��kh�h�c!����c�1s�@Q�9�v3Z�F�Dm�ՍPU�j�5��փU��$Ef6ִ�F��6�c��-�m;V`�E�ܶ�.5D_78m�����Z`�9A4u��f7�;����Ap3a��/��B&�5�?)⮸Sw-����kX��C�'�L���8M��lY}쐴Zڌu���譺!�5�嗘*�Ν��^6L?�`���&���)B*9�̐�i0Ʌ��������!8\t? =P����ͣ�G�vF�q��FJ�@tu7�&���v��H�=�8&,�S^�aǺmzo�
��x����Dȼf��wƲcg\��x��d��싹�f��et�1�BH�%ꗞ����~��"=[#���؞5ǌ�3ڽ�7��k}�1e+��op��Y�����+تT���\>����^3'N� \e1S�󺢔��Btʾ��q�]~��*���z��0�l��6@Q��O��L}��y@�ɕt���x[Z=��r����<=(ov�{�s�G�K>�y��}�s����<&+"g�+�j�π����L^��N�O�"�;\��|�;�o=���]�������.��TӞ��o��t�ω����N��ӖOuM	'� =H��%�.��Ls��ќӆ�״kO
�q�<eM�}&Um��o��#ܥ�i��9�B�%>7�êP��;��������Zj�k~�B�偝��ĪY�eMl�B���n��Gh��spYfL�ѨQ�æ��R;�;��sE;��M�E�D�4��]��+����Ft�s�:V�@ǛY�EN��Ǣܸ����͑bŉGND�W�bJ�m����?e[�N��U�a?�5��VvP}�#Gs0Ƕ���O۪Hy�o�Bk"��SڸiK�x�`��g�EY%����{&3ov�]��(?|���c�(9r���ڤ�:^���R>��W?>;�@�w���wɏɳ\�Q�}{����.�oo������i=�u6�1�zK��T�:瞘��B&6kn<t����:M�4<籤^Y�#1�ݴ��;,�f�r��9����h��/��5�7x=>�Y�3�c�/8'��qzҁ������{N�w��P��糲�Am�.i��m�=fh��t��wt��=Px�˰$m01�QA�������V��Z
�Nܻ�2���ݦ�74<r4�M6��t�F��c�F{�5����]׼���2���
�T8�{��s��1�>�*��\�ת�lMp5-t<w���9Ӻ+ɽ��aY�y-��l��H���IL�
����-&�-Ž�*_'�c-���$����G�A�O'��W��қ�7y%I�Q+�W䭺��v�6�=��q+��4Mڶ����钜���m�e�=t��Q�8�odM�	�9��o\u!�p��ϰ��[�����7�0:�Jُ�ݞ������Q[��yg�<{\����{�;�9S�����@����j����"����p�#���%{,Ye�2�w�������������%
�ꧢfv-�E}r�������j��I�<��K��b3|����1S=s�(�ئ9�h�ﶯ��ةؕ�j��E�m�ˢdW[�����-zJ�W=�_AW�{ʀ���܃����Wa� �ӻ��Ef=�ʧ��Dsü�W+
���9����uVb��Έ����1v�V9����7�Ά���9�n��ɾLQ��㞕=���.P���&�o4o����:W��՞d�dO�B̮׺���{�;տ5�ڧ���z�!����٠F�cH���t�a��U�A1络�vM�������r��Eoۖ�m�=	�M5+��I�ibw�q���^,Q�uw�ryW���z����ݢ�4N/�(��X��b;��
R1j�(�Y�t��:cm�O}avh8#����^�)�;��U0��\b�4��"����i{}���(P�<�:�	:I��~�GS7�{�p(�Ś&}�u^�i�3�����=�+��#��1���L�����'gN�tK����5f]�T���Ɖ�K�mj}�kF
Ӻ���t�Mˠ���%�Ʒ��8�KK�*zhz�~�gբ�Y��3h�l{�{^zO���J�H�kkQ��R��bkp��D�.����`V���h��1CM$f�z�4{�y>�R�+��-5�U�f�D�"̩6��A<|���ߺ�N��Cg:��7^�,��c`�ɞ��!�~�=>)���>[u~b���_����I~rw��q��"�k8���zh'vM��S�J٫�������}�;}�%���Jx����/��js�|�O	�-T[I�[�6�[E��fl���m�玂`���4�˟�%��k�z@��;�aú��N�VJwLa���F�q��o��ǜ�@�b���م���c�g6�.,N��T���%�/fV;7#�/J85���f�ۆ��2��
�g='M�����E��F�^�]ӘRR�
A�0<�]�.;��cWw{�]*���m�\c�����k�'����I�â���ѕ�G��?k ����{�f-w�VB��\�_/x��U�����w�=�lN��5�Ӱ�1�ͼw�+�]�m5[����yXR������\uF��{�	�n�&�)��^������d�Mv��Ȥr/og:�]*E&��C��T�z��/��W&F�9��qc�P';����=q��G&6��&��x�:;{�;'��O�~8gW����5���d�!w
�Ǆ�����ˏ�D�ο��������-�ҭ��n�hIk����o6Lz�A�g���������m#ݰ{g���̞(�ƽ�O��|s�)�݁��)��E�u��z��6	9���l�C�������s�p���� ���zf �o����X��6���qb���z�{ ؤ�
�s�dϻ����bt{p����?�֍ѸŚ��*�ʊ��0�v����z��zg�������ϵx�]Ǣ����������<%rl�̾�T;`��o�c�tPQN�P�j��IH���:�F��X�d��Ք�ܔ$wf��+�!g����W���5��.��H����^}���>�7�tϼ�y�xب����n����앒tK����p�!���&��=y�87�<�������3S.��m�����O����<{d0�2W���矉�z�=ԝ/��5,���uM��G��L��X�[�#Y��-��M`��4�_���&�oxܭ�WGf)#�zlC=�r4�ԙW;�G�	��=��^L�&t,^��=Y��#�ʤ�ﾸc��Hb���ڸ~�b:F����y����o^����4�W�,�,���y�`��;cC�\ ����X���?�!)K��ު�(ʺ�����$m��$�N�f��-�Nzz3x�0Ɛ�*/z����*D�G}ł7e��Fv����������-�pT���r>��3ۚ$7�Z6�44���d�n�3�lpz90����X��Y�l\�c��[�i�[���"����9�|46�N�\;� ���nJ�`v��T���7���>h��:Pݫ�a��:;�)�O�q+��Mt��38H���3u��j�ql�rђ���p�{ʸ5��zH��]_=db�9�BPĻ]:�3'�v��bV,��ƙ��>�}p���w85���n���V;4�l��C�;{���f烷�Ex�۹�b~ͱF��ev|}�b�!AL;�ܽ&��vvAx�l7A����ēT�z.\��:�����٥��W,�CH�5���o'�բo���g��R�ʏ�_Z����kX��?W�,�e{� ��#³���h�:󦎛�~��XQ�����$,k�ޑ�)���j�"/���<|���+�'�/j_��Swq��1qI!=���L��X��f�B��Q!x�*�{��=�h��Z�}�s��z)"��R�i����b�o�n����jS�R��K��yC��v�⌚� {�;�s���\?.��B��m3V���J�8�Ǣ*��	��Np��shE� D�T�Z�~��	��%���dڰ�|<9j�o��v��w�pSy����p1�7QL���=�dӴ*�h��?���8��[�ԟ%���i�{�ѡp̓n?\G]I:�kѧuX�=w��.�S�z�e��9���p�:f��}��aIQUn���0��bI�}�fm����oS�J���9m��Zװ�2VU9p���[3)�崔��=�W9�lU*�l�a���㽓j�oV�o`�1.,�j;(M[K��&��A�w��8��{��1��1�Ŏo�5^�sS����$nڳ]�1�F�f�9��}E�h�N������e�P�M�;���=O��M�p���������?���l
�dQ3Ο�@��N�Oc�#,w<"���Z��Oq�>c���}�t0Hj�n��h���N���π�Pb���{����[ۚ��z�I�@�4�-����HƢw���0�[�r$��!��CCVk@�I��Ɔ��L5��_e���ƣ���
{<"��5�Eǟ��u�nV��\1��1��5�79/e���Ta�S�R���&E���W\=^dz�>.d$�vE�7�~Εl�6nO��:���0�R��C�%�o]3P��jܢ�\���%T��~�M��{��&��,�r'X��B[}T�=�unH��˝hL�����d�";7(�Nx��uwm����k�wvΉʪhy�zIX��x�^��ߕx�Ű��ٻ���|��I�W��Jo�~�i��f����W���vm�x����꺡�ksu���/��"���=>��b���^09}�7뻡O뭤�?w?Kf���voOP���e���u�mz�?Q��{��<U���X���zC���1�׸/;���4���jq���=�3�j�󜱫�&7ݔ9�b�M�_/{�o��6��`�9Z���{z_@7��ޫ�#r��nK��W�*x]��`�O�I�#��s}�3}
B�l2��q�Y����奈����|��G�~�gV�|���Ԫ<+�W~�R#*h�{h�T�:��;�7׷U�+F�M�'�E\��vZ�c�P��PѸ�ޙ��_mo�A��U����='�&�;	�lڱQ/�դ[�5�&&s�\��J�Τ5(����t��~(&H�&��S�y&�&A|�xv��Q�gZhlt2�l{����H�u�u�u-���ÎJ��w��eMf����@�1�(X���`��,{f�W���;�J�Dћ�H�=;S�f7f�초�Y���j��%h��3��B�AaJ�C�"��|����� _w7��e�.G�0n`����}�xqv���e���>��}��NOw�AsۿFfd<��L����V!]_#8��S�½Yח㻸�z��;��y�b�7�f��I2�ml�S���8c�5�]�}i��Q��U�����+�:�Q�p��65��y��;�8���,̤�	���a��@A����~��&���}��eo��jzL��x�V��N5�VVX��c}�#�x:���{����;u�M���p�y���Ϛ������fjBd�*�З^�^7^u���w�M4�r���K�UNeкz�v�ä�f�wuuH2w���Ѭ�q^4w��EwS}nz^���,��`^��ޚ�o���{��OPn�>�����/�@8�ۘ*6۞ �GW-�@� ��v�q��ʐ��cm�W���y�U����,������Y��@�g������譡mt��h_-��Fca�`�)t�]��H�,W	�&�R���"m,�n���b��$(�#u�Wz %ٓ�kAN��5��x��WVs��v���5��2��6�� ���7�b��J\�-_s��j�4/O  �M��sjg�R����p�SC���,Sٛ��wd%�wkc�����{֟�fCB����}�7c.��:P����uA��DWS4��D�׷!b�����&rZyH�h�I�Tl�c��i���H��C���R- a�x�[z�G���6���a[��ed篇d�j�=r�un�*��\˨�J��m�/i
�b<V^6�c��'BB�UYSV��WMK���4�S	'o �������b��ˑJd��8��F�^���Uyn�����s�c+����[RF���ōۡ ��9)�+��a0��s(֎��D�à�8�Y�<Y�Ӊ�s�͔��ݱ�[�	�׈�:��%q���Q�m��3�Y�ھ�Ca|��^��j�c��p"�����-	�cU�]�J�35�q��=]�b��c~/�����]1�4[���EY������a޾c]rAޤ�65�X�Fy���6Z;'��"�9�K�k��B@F�tԋ��ӵpr��杗����|���_��Ct��\��x����5d`���a/�7�<������
"Gl@ያ8=Y��x|{v������X��Pԣ�ڼwx���D�#;[����ý�7"��b�VKz�����m���S�G��'�u�^�K�����D�
:�E-11�[É��vd}:�����2�hAt�۔W��z��lL���y��y;.wvb���`��1Vz_E��0�%�p<��t)]����|ȨL����V��W;�}��T;L��=�,�J�)Lw�&��C�/�(���������X��1\�"�mf͖l�}Tgǧ��Qz���^�+p?�n��X�_\͌6��j��'���2V�=+�4���ms3fr���4��r�GE^��mi-,.9��h����Z%��˘'l����u3E�P��=%����;K�ݛ.Og�C�Bt�J,�[�f�������Pud�+�>�q�on�YU5#�v�I��z�-��o���[��0���b�+V���#L4(;���8w�;���َ��{3/䲲Ha3-f-+��y�(T��G�3�o��V�}̛�]K@HH�G�KK��]��2��m��v@�ZT�)[�ĜEV!�X���u����.�U�Xܹw�+����W��dva�ͩ��;�J[���,d�o�L�@�[�h��#d2�t{��T�CF9@���\�ٴ�r�t�Fp.�ԚMrr�M;�݉�5.�Y���p��(W��m�cjъM��j�u��+bض��j�f�.ZŎ��ÝlEh�A?_Oo�������}��o��������>�9�ڢj:����A�+�\9W��έT�VϜ0s`���j"
��Ehq6�O��������~?������~���>չ�S�W�A\�k�b�sĹ�y�EA���4�D\������[��SV��ACb���X(H�n����M�D�1�t��EP��PQMU=EQ����LT�U4��EՊ(��oPu̯R�����yi���S���Z;�u�1�MT�uY�:=Z"���)(*�)j�*��i�f�����A���SɠӮ��r�����l��E��4W'J2E%)G��Z�*�(��Fb�.`�NE-4,k�K{�:�߯;���m��}YQ����]���-��AB7gaݜ�8�V��LJ���+����{w�+��1u����z�{Ø�.�:�`!�)�����%�:���ӛ8D��O���<�"��Z�v"�z�$�L��r��tunR��A��`jϾU9�+��Oǎl�$	���A���8�AU�5O�b���"#�4�v���.�a�x��KE<��֖�&��[s���^�6�S6����������9Z�껗Q[҇��HtL�|i��Ο
w�`qmâ�"��Ԫ��W����w)��DcC��Y5l�*��a�|C�_�S,ޚ�Fq�(�E����V�ʭbPp2FH�����:�f��h�������CǌG��q��?  �]���_��KmY�VS@M+J�@ƣȜwp�֠ �#��ʿOxz���A/����'�9�M'9�dS-JSStt{���`����%s�D�D��҇�s�eK6G�͞���f�8��4��yNV�	)m��<�^�5�_L��)�\,������������^�5���D@�$����X����bl-�����6k�W�����x�+��L�������X`�Y؎qp��^7�	nќ�Z��/�>��G��Є���[}��0c���SlD��!ڤ�̨,��M�[y��4�N
�����j��0�4=�)�����M5k[����4;��تI�b�̦I���h;|�0��� �՗x�@]kэ������ )�i��]+CǜS\���`}ʿ|�!�yċ�C�H�ǹ[vOƦD뀨OH��[+pt�uFa�Wé����F1���~=ަ�Q�U#+�Dc� ��	����Ѵ���~��~��SS�/�.�]�!$��=B݄�0�cɽ�c�O�l�sH/�_���`�Ԉ:llo��k
P-�1�}���Y=���Gg�-��5_��U��8���K�����1���+&��މ�̨f�Gp/�{Z����X0�bac�q��d�6?ga�48�j�.Ÿ�7����a�,.��orcg2ǇݡW����"O��a;k���m;��R����
����#��
Q�MuY���W��3�MI��zx���2�w.� ���g����?
I���H>j��g�ƪR�y��z��׿@�!uD�ß�>[�!���(��sRG�N�3���ه�Ő�v~v���6h|��f*"�B��E��=-��7�n֡����Za�sY�BT?�@�4��z1��cd����#��'_i����ŻU4ﻄ�􃚾
5=��ƾɇ˒`��o�����P�0�S�w����	�A�Yp���唑.�!�W]����l�{e��kg{}JWv�����}�[��4��;�>�c�o8�c$a���u;�#��8���+�eBx�PqI�-]�M칷Oh�ˇm��LPM�j�A�ݕ�:�"i�Wn4��m#���?�xQ{��nM��iW�w���^�� _��qxו|�St��!UM@p�_J`9��$�ħ6-'
�,UW�Q�h7l���ƨ�]O1�G�ޘ/Uŗ�����}�CC^�[	����i��*L��ż�\���˴��
h�'N���k�=��<{���p�|�J�0��{�e�#�D?�^����7�%�_v�O�:��=&��x�O�|�C����2�.�8���+�gj��;� ��? ��=Sܫ�@K\�Sch�a��mRM��Ȱ��󍑄��	^���[��O�x���PD��$;�!|z�%�g}�+~��o����ӥץ����*�<fo]���­t���ӭ"Z�Zk����'!��b���O��g3w�����zH+���y��1��R)hs&r�Z�PK�mr���������̕�gƚ"J���zh���þK�o2����+�%�6';�`{;#�kh�J��]5�c�880�)"x�u�]q��[/,�l/i�3���ų�0���|�L3&�eCvY�{r�����Cx��-f��]i�`7~��B��ŕ��"O��$yH�-a
P_�~�����]�kܳO�{���zVzܗ��L�E`�Wszj�s`�l.�ջu��3NV�A�O�}f�f��H`�W��a��%���۾�N�^�]�����)F�BoA�� ��d��gDn5�zT��������+j��_���>>>�e��h�Yb�������C�F�B��A���i ��e@tM�1��^d!]���3P���`�1��.Κ�=1����Qi�v �1���.��M��My��]7C�:�tS ��;��f���a�{1���]��z�����>�g ��>MF0�쪖�\`-~;2��^m:� �zp��c��P��N�*{7�p���Щ������F	��#���0�~کnjJm�d&T-*��4y���b��j�_�gd/]>�o�uP�V��+(� pqfZ���e���W�'#ɹ��	L�*~�5�e�7(�C�\��;�0��!^q�cНa�Z�Z��,�@4�YB`x5"�@��+w�Hy���é�k���c��fy���D�.���)�JS�|�u�=���PH���C�Uҵ���E�x캹��:r�����j�{�醣�H����Cw�Dw����%��	Y��=n��H�ʼ����5��ne!7T�M�|���*��]i�?7��t\y�)T�E�WJE��̯<��>�As�8Ty��[ZDp�c	�OI`[	���Ÿ�^�����r�a	���߻�;/�5�nd}#Y�5�lT!�����B�vd�"�yo)�;2=�E��S}[�����7�%�lI�[c�Ơ|%�φ�쥔��Y$��i����Q{sE;��I�k���5}�}B�Y���q��rF��D�J�B]�����y��������]jr�N����}�N5�-#���OPAǂv�l��V0�б�8��4�χp�l��<z}�t�|+��N��� ��
�c�_�@\w���y�]�1�´Ͳ�B�Y�su�\O���9̽��}8�LsI�b�-A��{�38���ß7��b��.L�vy窓�(��U�\���%�^@f����lc�^��xvQ1^:��{�@�GD��ńM��Rd�k+��!�<?���5[�Cz����7�4�B!�Ë@"x�v-��M�؊��Ű�_[D�1�k"�5�cs:�"KO�mi��I㞱���O���2�;�%�RYA
�����\G-�������p�Τ<z"r�)i������aq������R�ʟ��z��!rTͲvP`b�QO�Vck�q�zal��ݠ�3g�Kz�h[��hq�'���@�c�j+�K��m٦�D3�l�!����Q"1�y�ZщOʌ�
= ^=���z^|�����`p���x,ZGx��N[�e������<G��

��8#����.~(�2�~���՞4S\)Z@H��C8eJ����3�Iȧ�]���������9W��r�ѺhGt�')�9c+3]A��`��Y�y
�C�Nn����;�ftd�A��Yt��z��Y�t�|�W�:�,��!ymtQ����ےc41�nj����;Ϭ�;1��!�3�9U������ ������:�ZJZ��[�W�ïDxp��@s�DJt���r�Z��I�����=z�m�d�l�y��.�ū�w~#�?�G@���1�0��Y���&H�I8�'+9�R��Xs_]���ܛs���z�C�>W1Nc��=0#��\Ǚ�l?ܽ��=��%� M��\�5��ӳ��v����tF��fC��k{���@�a'���C�=?�҈����U	�(��O�7Q=t�/�^hQ�G��^�5�^��|q!�Y'��J!����{�� -���L��R4f�bM�����۳$Z<�X�J�k��S��FM���\x����i�dฏ�@k�}�%ѻ��V��_�k;������bQiȾ�v�@ 0�c��G����A���>��хE����=��|G�5ƈe�$B��O�-l�۔�Φ���1�Y���sW��a�bْkr��"vh3ܮ����`��W�Z4:gkAAi���c���V�ן;'�z$�q�nd����J'��K]��x��ϩ��56����Bh��"&_�+��6������L�$��fU�mz�r�~�O�c�h�����Y�c��+�U/����g�2
y���a
�uA3���
�a�[k|;�B�q6-N*���T�8\�1�X7S&�ss[�6�J.�+w�e�.��[Gqp������f�*ݝ�(|=�����x?���=�z+mY�X�5���5V[;����]��rm�j�&]�[�Zz���`D�������?y\����/����p`��f�����|!��z8-�����T3g�����)U�'$�u�ᛰ�*��M'Y[���s�"nc�M��[.t�w���Բ���V�ю�Ƭ��s^�ѡP`b×�֯HFv�`ԇ���CC�8������K5��$�x�?E4޹��d_���vu����i��b)-1Xݕfya��U��l�P�o_�)���p�vJnj�'b�$dQ��rn<�FѾ[[���z���6�{"��oH/�ς���.����b�ö�2���˞ȡ/"*�I�#ݮ5�u?P�z9%�s_<�Ѹ�±�!�1���B1���!�شQU*Wۛ�|�s��&���kͣ6Ⱥ,�����Ӯr՟�ȃ���~���/��[F�~�}Eؕ�ĉ�(y���9ܡ9t(��E�Pes�W�\��T%�a!>�@���������b#�&�;4C�#�6�!5�=K�u^�T,ߌI�~⨰�]<\ا[!!����Z	my����0�h�{�#�A+�I��eQ�X�s��ڄ䭇)C��:�®���)��v^9[ȋ��\4����p@��^���:��bx���D� R�3�E�43�kK��i)���sD3j�m�ܰzͣ�N����(�X�ji������C9� ���ϻ�>�?:��Cŧ�͌�e5�}zhZ��N8�����^�Ĩ�[�R�a�����a��$E9XK'����_1��`,k�&��(�,9�R�K.�ǘ��ޛ��1s�_Rl�6�]�׷j[��ށ�x�+���p��2((���&	m:ݖm��{gSŮ�mlpȞ#��)�sƺ��Gب{�#�
�������ү���C�ފ��X\�����5�y��5HCƞ�ʙ�Ȳ�C�A!�(6���f{D��'I�`�%��K�����ZgF��NӲ���·�6�#��&���_�$<1�d^��"g͠\e&zBs�~�#��Ѯ�j�S+!A�c|��ɯ-��5�U'}��>{;2�eKQ���z��\���U��_��{��ީ��5�L�����0L�q�Hn�u�Ϊ�-F4Jm�d&O:��Άbz��g�Z�{X�� U�;�B�w^�������-�8��S!>��_�j�/V3E����,��gP�q�_ڢuu��>!���Yk��Wֱ(��*`x5��a黯�TŬ�5���A����/l>�/�R��	aꍑ�r �r�ʰ�CCXQ,kd�.Q
��Se���G�3���!���]�2�)��0�������n���V1XT�!G^��I��#!0�$�P����&��H���������W��?�����⒧��=�y�4z$H�3�b	s�x�E�y�)�$i0��pח2����9�j�w��|����}��_��:E�r�=7�D��i_)�dh~�~O�����G��W� ⫙^�:�Sֱ�~�x�e���Є&T&n�|hQ�a��*���z��"��8¡2�gI���ܵ-��9��c�]���������9mi�!���GAj�,�^ԗ`���V���ͮ%�5�b�:�ȴ��9�;��ޤ&��,r�bP��#���k�1-��h��ɛa���VZj�G���b$��:��T�sJ��m��l��(p��� ���� h��~?/�mWtR�ʻ�~�<{#��=I�O����㤠���Qa����38����;��&�Χ6n�{5���,�Ħ.g2C6O�e�c��8��&+�C�z�N�/�<3�/۶r�O?&�IM?�����������M�X��Ar�5�6wA!�@"}�ӱm���E�V�Z����=�g���ŭo��L�3� ��{d������ޡ͛�Y�� %�5���xU�w�6�ݳu�j��n�Ճm��H�
���X�
�2�4b��N��I����y�d�f���Q���ny�}GKZ��$,u�.�
:���P�G)�A�gFd�ѽ,�wn�ɪ�`mX�7$��)���'��v�zc������YMѷي�~�W������������ X�y�Ĥ=���?�͗�^m�����>vi!Bi���7�>aE�Q�Lۼm�ئ&��+=�=7L}�\�E��{�Bf�5CZ�^�^����:/1q����	U��UD���֋�5�{a��c>���LŘ�馜�,�4{��U��Qk�Á��%��.F��U0O�:��eu=,�A��z0�5�A8���?x�4�����|9YMM+J?@ݨ�C{�^�Wt�n��C�OT�C�|$1W��U��k�Z���G�ۦl�����[rA���;��U��������C�Q�	ŵARʹ*�O5��q.�P̓'��6�����)�#=��^f|N���v�g<K��63��#ϡ�o�>�"U	��{<��1�J�ia77��;+�;ݹj����c���W��R�>���i��z�����G3���sО5�fṏ	0lX[mK�q�nAB/�=yw.,Hw�H���o�%�0�������vs�e)Jv�"�&���k65�1�%�dյ�BO�q6�bJ�������磾zڼ��"�/"�Tb
I�f(�@�/.���U�n�=���� �:���Ur��[�+������w��Kht[j�Y%�wJ��Ӽx�%f��&J���Gu�q��I'q���i��A*�Cb3o�&u;O�݈Gf�*�*��M�ۻw��W��,r����|:g`�}��8! '��\wS��^���7�����y���W7�;���R���`:�9bo]1֗|�;�f���K����*+�sv�^
�D�u� e2\�o��h^	�i�^f�(���������;��
2V��r�%�UW�r5q�bwي�X���#��2�H nk�D6��ᄩN��w���HɍNkNS��3���P�L�C��F����S����ْ�6Vѵ��7B���iV�� � >K�h,e;"�!'�N�fJ'��7"�ҘwD��U�I-瓛���������+��ܥ�J�w�����\v�e��hF;C�ۚ ��Y���d��uӡ�p+��%��99}'T���t\���Hw�	�Uw�xs�Kt�@��\��/��
�y�uq��v�$�����T�����ަ�C��x{���)#w�z;�����n��v1���tcى֥����bC�gv���5�%k#�K���rr��2uz�ty��]{��γ����6����ur |�[x��l)�� ���f���.��sd��)�A �7j���Z��-y���]@6����Y�.ɎR��S�4	��U��ò�Ӏ�?~����ޖb�oIh�w3J�ݰ���3A�<�K�7���]68��n���I��=h�}���"Ғ�����N�mjm�أ�����u���c���re��6�md���)���VM0Ⱦ�.Sv�hwe�
��&n���Lr���z�w�+]��&�x˩�tk��P��H�C5n�ؿY�����{�=�ȴ
�$y�1XyI�^e���\�əD�-��M0��@ǺM����o�_i(���l��s6NP2^Q�dܩj*�)��:]���}a�f�6nM��:4.+t㋦�Μ�h��S>��⸶[:�����.���5 ,ZT5��t1�MgFCZ����Ճ���N��e��R�KADu�Nu,�h)���*v�v��z� ��	�šO�ɽN����W�;���=|0�h�O|,?)A&Em�ggQLބ*�Y�o���R�ŶN�f."�I΁�SNb���2[�E���M�rF�/e�ʒE�BL�>bwlm��lS�{6.�rfY<9����&���ʼ��KٽdՌo�6K07V��9%����x��oL\��}�Ȥh�� 8�Fu�ͱ#���7�%�;��0Z(���P0�����;K�@)��tmgY�܉*S�j�@�C�Ԛmrޠ6��B�t�c�D�$��u�(AT%5D}�|�>��)���������~?������~��x<��i)l�|���:��Z��@g���������~?��������{�A���%Ri��J��@R/ �c�K@��-)I����b�)��KM��ݮ�Jħp�i(e)��4���uI!��4xO$9��ԯ&�9�N��C��<���+�M�;�S��f��U%�E�5�4h@�;N���w:�9{/���z��&y��C�Ɨw�ՈJ��w������0�R���-f�
J����	�� $# �ԋ�P$����������3�2Jʁu�� �c�湗i,;x7{ �֞��v�E�"��sN� 
��a������ږ/�h��?�?�F�2�����Z��E~$)U��I�
P����/_�{���Ǉ���ɘwڊ��7���u����	�SI^�H��������*�/��:�K�� �X��]>�3<�����+h��o*���*��zr���=����,1���Ӆ;�?D~Y ����I86s-�qOŤv�&+������i�L>2&���Q_�T���1�3"$�/\���n�:��ȝ���خ���������
k�[�h�cv1!#�E�\��z������"a'V&.)��ϙ�j�ٗ��Or�3�9}��q؅���)�.ֲl�wވ�Xo�����)'��I�x��["�S�bPֺ�«"T��h�ׅ㈚֞�J<�(����O���Vk���b��Oܩ'c�eq�E�����	��e�J����[TED܎v2��֦�J	��:��%�y.�g��|jʋ�8;�������&�m����`��4^�n��D0^�~�i��B��T�SM��:[O�v}��tk��8�_3�ӹ�d< 8 |y|�؏{$�%�4:!�Յ薟U�Y�J�/�j�zznϫ�Գ��5�Ϝ��].���L?���}�B5�~�d�5�ѣ����Oqr-��o4�nv5����ds&t�.���L��L�u���}�)�fX�;k��ٙ:Y�e�⏈<5xyу��D�^�s���%7*�D��JŎ�������3u�ӛ[ʦTF=؛똑V��T��;L��I��w�P?���U����W����{������(�gso�n㛏�n�E�"hgӾ[�	܁#�j�����	�G>��*��;u�Uģ����E�G;M��<���t�xҸ����A�K]_^������z#{�o9jyx�,��^i�O�xi0�0��֮Qy�%�;1q�O.�;!��ض���{��j^�Hh��y�^u�	�B�x6ⷊ���G2�J����O���ef�}���y���+���x�	�L$sm�B����[�c�PK�0���6���^UEv�6;�o(`�n��A�	t��G�0��5�%��Q8֬�-�����ַoTdw8�qҸf���KsQ�\
3��h�y�R���p�D����-���mU�r�{��Jv����V��Ë�~.����̼��-�{�[9yחt���0�=�j&�oT6�������#�u�M�nW�L��_<�t�C�Pi��I�ʇD����N�
ְ�ތť�NBP�\>d�&���{v5�ِ�xj�AzJ�!C��g��t�< ���q��^���5�r��g���S����깃�r�Ps�=�b��h�"�	o!�=�gf���&��ZI�3�-����W��J�+�Mj"z�4�F�'3d�N\E���w]��*� M0�39��MV��1�8���j��̸�D�ݵSo�e�AD��
9�UAw�}���}����D��?}��z ����q1w V=�5��UKc.P���*2���z{/��te^�Ej�˱âgO�b������t���cA�A�x~��ڨx�	��M��qz�µZ�ն���"u�,]�瘠�E"������!��Vϸ5���e(�8s:a��1Aܺ�=�9k'"	�u����	�T.�&��Wڷ5V�(��ab�v=��]�>���W�Ԋ1cʴ!ս?1��}I�`/Ȑ!���Ѥ�0�����_�[��Oyd��7һ�o� ��P����%�O��}�ȷ�}tڜ�Lk�n��r�бk�z��{Vr�[A�١��f�}��逛�_o'qUeWCа���X*��q�-��D}�]`ϧ<��Ƽy~A���0��0r��p�n�ėQ�X�'(]���Br�{O]��z+��C�U.���A�2<���#H���A=@t<6(���-Qi�x��dDi��o]��/YS��9/T�R�es۞��:AO���:�9]���e>�3v�������l�w9���J��+4��]�;GL��d�:d���*�;~��̄ɞ4��}M��7! ��{j��w�1��,R�����\�K�t]6Q2���:;O����;rU��u���o�=���G�ۿ�z����������=�瞹�}럞v|��/�i�d��1!�u>Z3�ǯǪ�V/�<�f�x�U��������}����\��%�>Ϸv�6�\�~��=%�@��:"ص�!����.���g�=�x��ZD`^hH�s~P]�C͐�y6ÃzY����qh�1�ӳ8�ҽ7{M��u���s��_?�"�]�+�sCPC ��{d���^=���i��4�5��,9@�E����ʎf��W^l�#�5 ��7�C����
`X|a��?�Dde9��G>�:׸�;Pu�Ȍ��|��
�q\�˫�EW��o�՜_��o�g�;8��R�W�)~}NV�7|�q5�z����ٻ
������Jm�f|���(�'�*3�(�ǫUj<��$0�g�������߯|%�K����*1����q%�~g�K�ҿ�����՞4S]�n�emY�L_���$��(�Nd��2�O=tD�I��bS�]"��IRkn0.�GnC{�gv%veO���.�x�O㇄���\�}	A�<Ѓ��_|�/:�{�Z���̜�jL;2�'S2��WGr;�2�vJوS����AR3Y&H p]Hޔ�W:[���U�[������(�P�u�fQ��P��y{��!��&��R�����H�ǉgB�(X}���:�[�j�	Y��w'2�Uֳ��;]�_�+?�\�*
�=����ދ�]�w�]l-��#6]�f�-�_LC2y*-M��cG�xŐ�
>!x&v|>��4_
�i�e*]i^�Dgnj,a��~Xy���ét�	�?y큰���v@���]�fr�ڙ�P�UVy��Gl�b�uV����$kz�(�I{	����ď�������R�u�뺴tA]yU��6����BT�n���k�wINs������}5R2�-ݛga�P{ݺ1�dY���h�<�;!�Y�~���K��L޸V1`s%��6Ʋǿr��m��2$�s�de���'���ϲ���Nh`#����ЙQ��V�`��-�d�پT#�n�pm9�a^�@�b1�Nn&K�|ig_���؟�h��MXHG(*4Gc�	��!e������Vz��x�l4�g#+��_Vgs���E�ߌ��dW�z�_C�j��W�m�\T&��1g)y�8&�e�a�;���BhwO��y�ި4-aƨr�Pk�"���	�#E�I�0]��,�����W��x��O/fִ����rX<[��<��ҫ6p��SSʒ[�����|�e}��+g�fad��z�dy�>{n"�_:�'h%��~�}�0项��w�޳xyn{��F�Y��-ح�OX�زmM��=�i���E{jm�+L�[��A�u���K6����_�2�z��H.��TA��u+u#ky{����;�ίo꨿_�g9><��ý������Tk1Q���dR� �O�u�NV@�4�V�ю��5�d�RO2g5�b�=Vn�̺ˆn��O�kDV8ژ��>Fu�PɅ�@�iA�]��T)7f7J(9��[�ysy�n$6��0��Y�U��TH�~k�.楴hf� p�33�g���e��d7W�J&:���"�̒␍�a=�m
�N7�������O�������jU�G;��k�[���Xn�E7�H��^K-A�[F�����nvc��NN�z�6��,�,h&����S�(�^↖������Iq\�8{bd��f�תk�6Z(�L��v��]z^S�zyP��S	�fW<5W(��RX��CxHO�����C�Փ՞�葴�&	��>Hq�J�N��e�q[�Qak����X6�����g?Q�=[?<�%�jZ}���ϒK��"��lL�c�Gc�يdemzm��������u�絎���U���@B�W1��/P��M��W�k�\�.��!��n��vR�|5��kIU�0����>��_�W�`a~rq��� ���5�1�۹���>������v�(}��tR�2�K�I҆�F�(�x�lU��nd����vl�PV�Wf��;�w����@�����s��եи��:б�'�ӈ����0�x��s>2%߁�h���m�,�O)�
ڴV�#����/f�2[�Xo<����*��G�rW�Q'����DҬ��л�{����"������0�Ⱦy����� ��S�PԴF��6��Þ8�JR�?G�7�oR����bO��B<��'b��u鑙ǚ�M��^ҹP$ך���ۦ"z6��,w����T=C�S<`���愈�����a�_d�6p>ϝ
���xz�\��z�P!ub�g�v]8=��Mۂ�R��ޭȋʖ��GF&H�9�lc%�0��c�40�����pa��]��cH�5�J�'�G(]�_�KU}��A�VQc�͆��e	�ط��G=5Y;C+wr�~��qRY�A��E&Y��)�ʒ�5EP���S�"(j�P��bR�����p�*��=�T{�+sG)�	ξ����(����Lh$i0���s<`6�F<W#����ҋQ�ck��2���"!0I�K��| B��.��Qt��]/s�1�b4�����a���Ţ�ul��v6����[�(V�7@��<�۹�2���Q�yw�N��QQ<Û��������{��� �1�̡��׼�i>{�L�wF��L�WE&�=}Z��4�M���-��a�C~[�P!J��V;iQ$�%�C+�������g-�2���9@�������p=����� ��b�#��}�SO-�����Ù8c�h|{ ��
�z|���Q�LU�Ƹ�U��&"3v�;8�u�ʛPڝ�-@��x`>ϘG� `�:W��䟗�:x���
�l���Gu-�������v��u��R��s��8��bP�f�߹~�����p��
,f�r��q7j��ک���M�C���R�^��sO�Գm�`��5p� ������啕K6�ma	����ļ�[�ln9Rcl����[c��<{Ӂ��۴7<�LB�zq7W���20W�z!�LO�Z�V���@f�c�/a�c��8��^O�o�D[h�o\R���lfn����9Ѱ��3�O�.�J>���g��"\ߔ��>��;Ӭ!���- ��'���+VY���n�`O���zf���bY�2e���*���U���q����|�z�x��z�Ú̮��	η�%�(3e��r���j�1�������<�囟d�W�'��A#=��S���f��CŮ+X�]A�gNsױ��:��`B�XO��c�AQ�V�cM�� ���)d��9Ǻ���D]��Ge��ː�j6�:�x����{����
�1V�z�%=���7�#���F�$����9f�(D�����62��iEu_c�·5u����8ȱo���q��?��U{��93��
z�����^z=���=~OmC�=/l1zk�U��dlm�zA�%6ߑ�5Z3I�*3�(�^=oV�^���v���*w�i���/<�t�p�)h�#dL�|y�Od�(F:�K���s�-�?D��~�n�F��}�C�{FC�QYx/.�x�����i1�����'+�i����<���'��%9��)���}��c�?L�~�^c�z� �'X��h�8�`cH���hJ���7���
�gЇt�[N�.	�I�*�ë���B!������wE6;��-@�az��y�=���3x�M�,!�n��y��U.����Dg��{%��w4X�v|��<o �������i���@�`o�sL/ ��Ya���G\����-i/Q-�V���(�PY#X��Q������U��_���_Wn)޻���f�o�)�A������2%�S�(�t�[^�$��b-�6�j�Ъ�|�q�ͩY��lj���h�S�40�DXW�D;)�K��M�j��o�1���ܺ}[f��\m���Üm�u*����lS�1�Ȅ~՞P�I,���u$��s4�&-4.�{�6�Y���vĈ�W��9������>]��_V33�PG_�ݼ�
q����%-�
���dmړ�n�
�kU�]q��ĭ.����>U�i���#���3H��r�
�5VѝW"��O��܌R�/9�7�j5l{a��=���W����x�� �8����+b<���_2_�̊�\1x��+	��)��,`���ؽb`c%[�_�oq۷e��6N��Y]�\���ޔ!Y��baط�pN����O6D�za^�q�"&u�)�r�z9v���X��R�\�%>�^Z�=�y�~�l�N��6kɎSj=CdR@@���_�6������Z��<!��|�	��R��ZҶ(��+d�1���8]�e4��.*	���n���$�.H����=0���NKͶyt�����PyO����J�����w8j�V<�e���]W �<��"|�P#!��f�a��/�E4ۥ�tܘ5���M����jv��5{�'�T[^�-�N�����B?�F����)�_��p�����7�盺�sS�tN�YJ��2���ٶ;"�t�z$ƘM�$B�,*�E��5����Ý,�#���7�>�iJ�&@�LR�t�/^H��X~��NRd^�|>Ϗ���b���D{��,���,���T�7�%��ls�/����^���Iq\�Q_~���V�Y+�z5���%<4�C�M�n�=R�T�ev]w	�kq�5J��V4����ws�چS�^T��9�39M�v�2�T΃��b���{i��z�I�-#Eڛ�6�"��=Nst�-�s���p�йؔ.���˼�Wu��+��_SC�6{\!̺�� �P��
�Uf+s^��:�P�D��p{�Q����r��C	�Ъs|{&m��s�cj�f��2�Z�K͚��t���+yu[QNV[Wm>����cR�IX�+]abn):��K��kY������h䨩��/����ȅ|,]�_����Q�Q��^��%*��X��p��+h�v�a<�����{�AJ	�I[�f�������SV'HW���H��.����82�ř�:��w�S����Y;�'��q#�˔==�e\��S�o�T��&�[��-�F��3��5�@�_Tg����1�Me�(؀mt���pv�����d�8k6q�@Sn��i���E��b	�:��ڈa= ����rzY�K�����pM�ڹ,�䅡+��a��w��!������)N=.��fL��g�l�*U�t1��f5<��Is_i�ˇv-��S��N[���k�X� 2��tkD��OS��=JVv�GT�ݨ�|;��������H�&Ju%��ر}�jj���{X�Q���f9�â�K^P�,S*�#G����]ԧ��f��,����n�d9I,�k8�a���97���F����P���g��6Z�l�;0t
�w��؉�Ѓ�M�'�c����r{�����h���	;�1���W�_;�IJEjܝs�,ZM3�N�s�L�ÀW[Y-���q����<�"����m������lv���>vkYԸ�αN�^��_om�cv�=e#��MѩϏh-������iU�7\o�=ʶ	����7b��V�MD�ݫ+�f]������lm��c�N뙵w���L�B�h�oXgۛ3�ﴽN��ڸ�Qm�}e;۳k�q[9���=3:mɻ��h'�k��%$�Z.��w�V��ә�<=�{��.���Z|W��5c��1�آ��V�����n�����L�؅����%gI;B:j�6��"��p�g�����S�>��Z#5��#o�ަ��Kq*h���}t��u�fr�-753����Y{��,�81�8�쬧��Qڒ���N�w��WvpZ	�A�g
ӷ9��7xMC��X�&͘�k���2e7���usx*��S X��򒁕7$]Ec�<��a�P-�W��d��[�ӕ�"U��L��Kƥ<�OZa;HuƵ��	
��н��+�y!̊��Lh��{q_c���V�fkk�t��V�sz�sTi��ʻ���u�֞�sr��/sX�嚴��ޯT��kI�euQWݥ*����� �s�����|~>?������~�_���:�5�4�0�(h�c�V�g�trP���O�������~?����>��%��m��B�h��+��N�Il
�44D��hM�h�E i䆮g�s8�]e1'^d��t:�����T��:�us�8�IWV4� ��Ɓ�M5s(h��-��WV�B�tدQ��)�Ҵ��T���/�d}��� �"Rj��&�7�i�@4�)"�y�9/P�9�Jj��1!�����4t:܆���Tʹ�y:�t�CX����mݴXS���NZ��s�:��g-[%���O=Np��%}���T5��lEmì�#Nn,ަ���?o�/����8�?��xx{j�^1+�~���ב�$��_�Oo&@Y��B��/7⤱Gf`��tn:�f�������X������{ʄ���Oz��0m�o��,*�O1�Ffy�3�Ѓf��Wv�!�]&k�+AGځ0����5���&5�09�oMV��w{	t䵚�(���OFwj6�T��*9�����r��A��?��j�A��/}3�Z65vҋfqU{ٳ=�q�c�dr�kɆi�f�O@��{�A�.���x�	��*v]�*Z!��e�wfÝ��&�uCvY�GnQo/�q�c�DȌ��/_�1�R��]�}ݖhF�\:�����d�&*�@�F���
��e�7i�^=���Hz	@A�r2�'����nu�ƅ��%Q�U�~�����S:�:9�"��̆��E�{��~̏x<5z�7贲B�Ǹ=Qp�:�;�Y݇3<��-y�0q�P3���gD����"�k����5וRp��!�;��M(OػM����t��^�P���{��V��	��T9��l�O��Rm`+D�g`���a~��z�.��NZ�9�2�E�
�J�=�HD4H�%����ٳN��-k�p�)^_����d���j��V������VU:G��;S{�6+��V��,��=X�Y��Р�wn������l��<�ɑl��^b�F���|��QA��������"z�db����>?��L�(���ߟ���ﯾ�:=�-���%6�FB�:�J�'�G(]���2�6)YE��������?���7Ņ5��W/}\�Q.� ��g����c�%��!�C�k"�gtv�j�j^��)��aމ���	w�y��������g�������u�/Ⱥ���#)y��\o5�0�[7�*]���R-gz�[���$f��A`��K��#��D�����EL,"}t��x�=��Sh�����ͭ�^OvexokG�d����=4x���!7T�M�/�
6҇@_�t(q�1I؊��	w_>�X^�&5+���Zq.�>ߘG�y��֘��~�DIu�m���ћR����[W,�:���8]��z�N�r�@�>T�D��怃�(�8s�x`n6!���}:�}��L\�S!7�c=_�J	{�TX����E�~�������"�����!5�.��=��^(�����e��reO��N=�\�,3�5�a�	Q	�7H��A��0��H~ՍW��\GV�3 '%����2�Jr��Z	EjLZ����n4E��љ�8!�]H��2fdx5 X���T{�c=3H��W�].̐�T���5Gn��[�����g��I\�69�ƱW��`WǏRY{���^�Ӳ�<�x�U
�Q���uJY�����fD{���:�Go���'6�� ?����?� <��/9�ֶYW[3c������@u�����Y��M�G�ౡ"'�~Pk}�At��פI��������u���j�&�x�;�e~�輁��[�������~j��&e���5���柑ss���op�m&iB����9ϒ
E��VՎS�3�J��G4���4�22��_lܵu��j7')������TͶvPcK'Iym�+��ZP�)'�:蓿����>��OAf���OW�V0*�m=zA%���,m�%�=Gj�Tf�rͿ^��\��ۭrwu��DK��Py�A���C������%����=6h�uN��T{3�J˵eyM+J>�G@�(N͙c�*ǩ0X7��/#�LxOEלħ+x�K�O1o��r��x�������L���]{���U�<�D&�m�1��E�����!�MRҜ��j/2�ypYۜx���rk����t!"���0Ơ��K�������B#���)��n�NS�D)F�*��*9�Z/g�KYtu�3��g�sT���ڡ��#�D���B�@G�M�=?���,=Wi�[���2�J���j8v��P
����_]pQ�����t"t��C��P�ܩ�3x�n�q���R*��̛�l�7|�i�V��̳AmǷ�� �����'d��]CC���z���e��P�������x?�������eԊ�xV1����^�zh��:�w����F�J�5�ćA�/�F窷�ʟ����{}�P�Z��;s�^���="���=V�czRr،G�EL0UP2�#sr��C�����gܑ9���/���������GVH��v�>#��4�\�>� r<(��^�M�嬌���F�]����E��A_�.������/�����Y�K�6+S�DN)�*.��cv�Foj,��;k�(�j�c�����G< Te�����00���ܠӪ�WQX�64+�r��\�2!x���w��ʾ複�*���mG�l�J9����b؋��QIS����:��kof�������1����l�Q����'��Ώ�����a��I�6
I��윣������K�D+�<��5s�W�gc�j�A��%�CRFu�6-�6�D�>�W�f�m�:q�f�C��0�%c�e�0Ci�$_�7!�򢰾^kpa��%�Ս��A�)���	���k�ذ�T\-��J�p.!� ��F_N����诺a��:�s��C�����엖)|lŷ7hvd}1Q�ȹҰ�O7�[���r �:Q&Eܹo�~���o����A<�va��C7�F�����18���xg^J˼��ْ�v�y8��}Ә��)�8�be�cYf-]�w�B�M��R�kMKt����P�y��k$n�{ ������}��������E3�b%�tȞ�J��ܜjQp�1�="z<�Ⱥ�I�}{,�/_2u]Z�Lb�]MlWv����9����%:�Q�jªK}2fm��E�*���	1� �s�j�O���u��y�,Pb��1 Y�v�oR�� j�4J��^��4�p�;�0��{�}Ў{�����ɚ����X��y�%�x_v��)�S.s��X�Gf���yIh�%�&�ʅ�TM���x@�M�A��x�R��k�>u�x��U2��Z�E�ʒǚ�-P4X������9[��>CL$3R���<�q7�3�muSƅ��8���+%���i�ȼ�ם�WR`�����+S�zA�OO����c���i��X�����Gv���lv��,�q�&*{U���Vn\qdF�4�@��xxlsH���U��TIŰ�:;��9B�2k��&
�ƞ��%ۼ�Nq���XHԫ��^�H��p�W��L��q��gд.`� �W�,�9��,�#QaC;�My_��0}���^�E�t)��M%��>#^n��]\EU�#��UE;AmJ��eje�����5�`y�^ܜ)z��1��!FU���٭�nk��>We5��M�xX�Y���e�g]uHt�Փ�G���	UZ$����&��=�oMrܼݷ�L���s$���3����~�����?�������If�;�#`N����?T��/g״H�y�hwH$=%�F]�_����&Br�n�1��;C�֢��	oH>�UB/�O��߸*���u�S����}O�Ev.�fU�w�e�:���oJ7r|�\e�j�L\:�vzm�� ��a�s�Ȫ|��j왆�ٚM/����W�~�=��g>�܂��X�į9�ׅ��	����k���g�~��������o`*r�x��]��ٸ6U�����@?!)�ѐ�Z2%?*9B��ס�Y�j��v���i����Ne��ͳ�]��D!���"E�{�Ob�j~BS+�S�*K�!B�ѓ��5���jD]Z3�7�`�x��0�����*`pjo�	�5�ޙI��,����7�H�a{��h<fv�1�g��O�����fR�p�M��j����8�����A| �_O%��+ɑa���:���c//'��d��n�x��̗mF9jw��iAC64��	�&��ТvP��Gm�+u�k�!�n��FI��F1g}��	�t~n�P*s��?��Dp�n�	���l��pca��>��[�8�2��v�g�1ѱ2��d*��k�,�6K	**���
��2ճj�´� ܗ_}QQS/��;�ufr�PӨ�A;�U�J�(knU����;�9ҍr�C=�n��`p'��p���1��l�������f�ު���3x`�F�!P�j��È����̟
���K#��Z��^Y�Azp�4(�����u�ܧ�q�|S�r8�-�0���J<���Z¸�Z��+�����I;C��]!������h0��M�Ta�E�
�a08G��G��óm���M��G*LVx�|���q��KگE�~�U�_���B@k�7��s5�(��TW��S��Ig��,<J����~����s�j!��Nf��D�&�&+L�Wr�B�ހ��a؄}#�R`��y	�s~V%^&�z���� ������s���º���HLo�'��F-�A��]X�L|��F�3�+-���tdVG7�eW�;�}��[!�����$���YA[�0��{6q9h��ֆ|�-,�t�6�ۅ�&���9#�dwNC��ؘ,|��z�� y�S6��A�,�`Z�Kˬ=�zw�=[¡�)+p�7˿TWhx�p'�N.>�AUcoj+�;��ڌ ɍ�4�}aY�"�Я"k5�'>����c^�F&�%#�d�,.b!�l7ъ���N9(-����~<�%��#�a����Tv`ˠ���,g�/"�����ʑ�5�v��7mq5��t�}�N�J
�:���(�vrx���N�ǵ�Vv��w+�����ٺ�P����Ļ�6�9uss!�ŝ���������y�Qʍ���b?����>������E�U����R����}j�{d�Ҵ�rn'Ȝ�0�r/��	��U�;��*:��w��w~�q�O+c�E��3f�vO"�:��}�Y�JY��828e�*T�5��1l�}7��կ]�L8F�y�!8�NV��YAm�z0�y�<�-���M��S��c��^���8�Õ��Ƣ�0�v�rt�Qi�g��%�qyK��H=�Z-���q}���f��:�����au�V�8���«Z��>�YX��Py���!�P���JL��ټs}�(���^�G˾���	�Q���f�z|���ɷ�Q�~F�;ine=�MX[�f�LKش��� �.�D�~Y;�$�7���0Xp/��=Y˗�m���/?9������.;(�{�Y�lP>�~g!�vֲ�.��w��-�%�)ɛ�~2�Q����!%�`��[��m/a�@�s�;h(M�*1��M�v�U�T��a>oAؕ���V��w�y�D|gy�C�yg)i������ճ�g�B�+���4���T㴎�xg��ݪd�Y����!F�gc����ί����w�S�GH�rO�^���N�W_T�@�ɒ���+M�p�m�Yڅ=Y�3q��=#��`��\X��&؟ƍ,F��їi��#1��������<��8$w��o������g#�<s\a�W�L�#M͖?B;k��)G�<��^b��J-�jw|��om��9s��ۭ2�a
�`��|�:R�j�S�����;�X��l���x��'� ��|Ǧ"nA7��^]'�vN�Q�Q�B8Ȟ��4����7P���ե\��v��-����]���`�<�������נ�]\������4��]�usz�S�tȢ���J�O�1�C�� �Ⱥ	;q�c
ɇ3�=o�+3�Z���1�Q�L��$��1)Մ�VRN.�f�H�hTN7�A�m�/rSV�]��/�O`p����}[,��C�{z�&X�LU�H���Q�焼��e� �9�v{����G�9j=���DcH�A:�0�_@�T/�T=뒞gת��P���4!�.2�9�U�����{{�w[��d�_KD��_~AY�{T�L�R�˨Oz�z��ȫ�>P{�w/�s���1ɵ�i9��߷ݩ��;v�<⇹z*H=�!������@M��^u�Oo�d����ϧ"Ǿ����@_.���*���҆�Lq�X1J�8�0.��uS}V���cL_r��ѭ��}3�1$s���|�3R��PZ9�r��t7�)�tMQu<��T�"C���
܊wf����Q�Ƶ�n��<�4?�S�������/x���gVor��%�ʖ�������L�OH���������Z噾WV,�������CX>�z�yǼ�ؗC��>�a.��\#���69���Ԉ�)�f�_*:�n>���=�XsDn%c�e�Z���	�nm�ar��x�U���a�7��^��Q��![��a��U��f��>�v^�v�z̻O���5[�t'"�Q�޷]��x��Ҕ�Ap&_Fr�T�B*-�ݖa��|�^�Hz	@A�޽��!�JgWn�dm�~3U�����cX�~Cd��r�Ⳛ��c�x8}W��X�n���gz��=W��"Vu@��5曌�M^鋇T:/���'3&�蚍j:�Ib���볎�n��E���!s��B�ݫ�^%'�>�[sձE@bÂ�5���V=�e�ճ��&'���4�`mT�41,�d&@W��£�.�Nk�G���R��u���K4?��]�����xLB}}^A�v)��~BS+.JtT	�"�]���u���0�&T�VM�o�e��T��uL�7t�h�3���KR��Y����::\�阏j�N��̽B��j��f�3vݮ��$xU:�g��t%���:�A�TLR�}k.zmrq����i��ȹ5�B �Z9�"�EB��p����;3��ز�$�3��."����n=3��5�u6�����2]���CeB�D]�S����X/lщb<����S�Ւ�M��]ihP�7uf]�Pf=�%I[z��)yJr=x�w�n�IYq��u+�1U*�6wZ�(n^ֹM-��;j����X���uCh�M[��'8��v�)\�FV(9��@�f�5�67��vt8��������VЛ�o�r�%MKz��y
��']��襧-�«���ڈ�p΍���G�|��G��t��јd�ז�u'3z^���n�H-6�3y�O:%{ǥ��w��}����J����M�2��m�����0jX������`�3-����67/R��Ρ���rSe��aH-{�߶�Y�7[�t����-q���'"8v>�.�M�4G��)��(@��s��L����&��������5;7:�ҝm�!jQMf�����w�>o!�[t�)���;"�*cU	FP�M�4���p���ػ����y:.򶉖���91��m�iQkP�]g�j�q����� �j�
�W|o{RF�I�e��f��7.�^���<nV4$�J	ڸΫJ���*5[���э�G�l6U�yoU���73������yW(F`��B�Hy��e�Zɮ��Ф�����A�|quEw9�����\�j�%3�V�Zz塛fz��0��9�f���oeIWR��ϴ�W������'Q���0Io�&ud��Є�ޖ�nl�BrS(�|Bq��S����j�P�����������u��
S�"�������^�˫H��кwtR����$4u�^�M�i�1���P��U�Uq`�CX �U�<�O�ȫ��:@I������z���ˣq·V��D_����黧���}�q��L(��`Aq���N�]n�U�c��ں'�j���dfC�Pr�Fj{;6h�F{����*�e�ef��-$�`۱�_R ����l_Y�ot�z��N��.��.sV�*��/rwZ!zF���%�vu�-h�Q՚If*�l��Z��'	����T�\HHv���0��ʓn��ϢkA�0c�O��s�h��-g))ќ+)v�M�I�δ=e��v8X��V�ze9���9h��E~�h�MW1�b�.t<�e�K��X�35+A[��lD����r��� �8�h�)5'�����r�J�ś]/w�g%a\F�䱃vR�jp������\ay2A�7o&oP]:�n#� �1L�P�Vσ�Д��=O#�'D��SAA�IIA��4:S9��}?o����?������~�_p���9�K�)�)�@Ё9�������~?_������~�_�vX��lhh�)J}$ �Ц��(
y��Hh���S]@��m`���T�m�i6�	�JM�9CEr9	�ES�I���s)KT4:(��R�N��K��"JhJHQ���ѡ�-)I��R혱�i^�4r�ti�'!���9	��Q�(�:4��ܽ]Bh5�@E���
��)����l�y)Ȣ����r[�=]\��W8s����y�V.�ꔣ����@khit�&�`�ڕ�R�0r*�5�x��c�E"d�d�
�.��-7��mN�_U5�NC�.�� �M���aC�%�s��wdj05GLou��:ٴ�=��b��s�a�b$�B9����FKRBQ�Y�~-4��&a,�\E��3߼<<}WN &��?��S�Q����J$!f5s*`x57��a�f��N�<2N�n��9�6�Lt��K�~���x�ؽB�ϳ*|�֘�厦h���"�%�e>�$J�Y�� _Ey2,S]"/�M\�/��nۻ[�Iמ�#�=KƒT���8n8C=|�<�ʑ*L����++� ������h�Cв}8��pX����Ļ������&֡#[���1�/0B��۹���my~���NN0-^�8�Adw/U�t;�|��}���9V�vo^�O;X���Ʈ�$��;\m��&����O��:N�Y.�]Ү���E����#��#�z������c�
ئ��D����ϬG:g���z�?N/yq9�Ī��mgԮ��G�OnJd��X(�P �À�P��j�(%����z��lc�^�e�4�Ɇ^�0�ϋ��/�_Wj�����Xh�8� ���g���\ߕ�*�7oP]�_y�19cFR�%�!���@��D�4�yh��kt�V8W�x�_~1�?|�i���2j�j���WV8n�Z8�gNE���v�6�i�fw&,VtQΦ�hK��%��X�YX���ER^�u_��X��O����2�<��Z�W!�s^j����Â��G���LC�@/����т�1ͼ��Y0t��;^���������cj	�õ���Ӛ�%CZss����yA��>H)��m��6��ڡO�$��,���Ҧ������c�5b�2��O�1�O���!rTͶ�id�o�AP͜j�*��*1W�����^S������4�z$MǩW�V0J�ڊ�q�7�A�U�4�ģ8��������I�}�݊��^��siګQʾ����L��"X\��Hy]��E��z�̄�D�N�#+A���]lS�S.c���y�M|�Y����!�t�դ��*$�6C�/��'��y�u*��U���w~��:_�Ә��t	c�*Mmb;'� �.��>B�Y�nIژ�[���ܟ-ވ������e�2K�����"��,9���>G�c�	� ����d2맺o��<P6ں�K3�h���n�v���/^���h����u�)�a'�?I���7�M4-�{�?�-0Q�"�D<7kקzi�8�0�e���}*��W�bC���#Uu%"#��O�]��˝��v���y�o��@�u�zE7W�z������4�Q���o��(En5�V���+�7t �J�0��{*�г�BҬ���m�+/�[�p3����*ԇ=����(c��Uk��I?#���j�EL��w=���&3�bn������s���͵��ER��MU�m]��ݽ��^��8Җq��+�w���B��K>Ki��`�������J:�E���̖�`˧����7�dN�|�r�6�j3��
����_P�n�6�qQ��ȅ�<��E�� i/<�үC�)�����yփ���Nf�qg�=�\k��^>4QX�"qfh����c�����+��w_T�,Un�my�hG����1��|tE��P�J=["Rѝ�1Y�i��n�/;#�y��/	l��&	us�NlfϠ^_P���#�����0s��wʹA��(�Ƚ�SSM��y�:�Ψځ)=XXE��/���ϫ�6��l$t��Xޒ&f�L�1�J�;������:&q�{ [9~)U�@�!�"b�*&�{�*l�^i�x��B��d����F�s�)��w��
��}�EMz�'Б�P9�2��v�Ӭ��9\��Uwۏ::��3�#n���������ָU�S�*�	d�'���p�m�cD�-�
��C	-md�2��-����4]��1
�M���2NZ�^�����6���#�Q�çة�͔���=�����ͭB �7ak�l�z�(r�T�3E(`}��G���W�qږH^PV�<K�pԋ�y�6vv�V&�0Qe+��&ueY��� ��I�:a��:��
o�JV���e^	X��X��d���0�*+�~M��s"+/�,e���m���y�����v��QM�? �a�2�[,�4�^��N�L���X�(�LL�D��幛�20��(_p������Dc;��L9�_@�W��0����P�8Ⱥ��9������u��z.�+�|���\�$�����`�݈m��K�~��B��«�e7���uv��o7�;�Vu�Ǖ�)�#�ȟ&�}�b ��!|z ����~�j��F'�)��w+%��I���mG5q�g�x��R�S.t������+AF���Lx.5W�Wc���ܷ�T~�V�2�ڄ1[���c�Z��dd��Q�+0��=�:k���@�!�>'�2��2[5	�v��e�uS�'��j�jT��{&�����Ksqe�Pg����Zξ�����Ә�%�LX�S�~���uCvY�{[(�>�ė�����c���V�
�]���z�*�YX����B4,��R��Y~ѻD���3�h����u3�����mf� �[g,*;��r�>�`�Aσ�!d�������^����������M�X���f�c�Xpm���u���=���b͂�dx�c��'<��{��EU0���K�{��%+��f,��4�,��Ϫ n�����p�3��k���Ƭ(+yS�i�g;n�`kht����2��������~�ܫ)�**w~��=��||j��)��gU[��{۴�4<4�.���-��+���������ơ��0��ρ�
��軚.i�������ݗ��mg�������ƭ*{̋���,�u*<��zq���1��gA�ki
��f�F�j�S�^��BG<���+ �mj~BSm�	�Z4)=����`{�5���U���ӖtF[xN%¬�̙��b�9�:��Cv(�����V^%:�T�	�B*��^�gC�
E�5cG<��c�O���
��߅0}�zˇ�q��0����oUs��K=v�f3L����ǎW��j��,(<{��Ň��j�ڴ��=�L����|$K�}^Ifr����!-���
�x�ˈc����S������R��	Q���'�&�	��ji��*j�_kg36�Oe~~�i
��u�����x>�B�M	J�}�0�O�XBmk�j��[W�h�=����+�bm�-��|��Uz<����rx��|7 !�*\�[�=��>41�Ͱ�����KA��G�?ꘖ�%���gq�X���O)��]K6�. �M��TiC5������61�ֳ����i����s�%��j%���;�,G�^�(k�u��Fa]L�͎f�h��P��A�
�c��Wb�bq��g��΅�H`��u�L: �.
IQ�8dT�TŴ���7^���{�೷�BM7�]�}�WV3@����?Z"�!���u�%Rca�u>Z2=8�V=,�iG2�.���܄w�S�fԢ�;w8f���x����_ܻ'�͓̐��E�:��L�Qʈ��ٜ��Y��=yQi�LW��ύu���8����B9��+���a3�_�~�[�j޸���r��kXCOt�\<�+��m.�ױhdK< ���2W��֮KK�]���Zُ%��5��73MvIa��s�$�M�C�ڃ�
��w���O3?FJ���.je�H�-Q>�mn:���/X��	J���!^rVΰ,���͜/�ym�+�'�o�~����>��sF�Ã�h��D\{+�]��^}����~FPd�-���@�Y���ߵ`�늞Q�w_���Cx7� ���i*븚$:�F�*��A8ݦ`bM�Bj��*k���[��=��"7���R��$�4]�*a0Sz$˚W�[��e���]��r��c��L'׭�E�R�����j��\:��@/�m^���ok��{e:2��-��C5�zz��n�g5�j��'�­;�[����L+XS>�߹�����s��������Y���JL;�l�}y�fy�ڪ��G9)c���t蒆eӨ��|q���a��v`��X��܍y�@����t��3Pu�/�����rc��R�1�,�`d�a��3��,X�n=!�"��Xs{/����h�4�2f=S���4���'�	��81��ҟ}�K����/C�Z~X���{��oJ#��ދqq�n�������d�>�i�E��ְ!�s���Z��ޚn�S�Vat�%Z��a�����}sl��c^�;�R�6���lH!w$J~1~�:�5"���=V�{ғ���J�����F%��1��]���.�3tW���y"u?,����}Bٽ��ez{n�s6��_��<���`?t�]�U�ym��~���+B��<���[�SK�0Z�X�zrGF����nk�bԥ��O���
Z+��K�6��1xו���OC���V{Ո?���_.��t��o��Mw/|#~�v��n*C��v�q�b��9�HDYz�x;>��^	U�M+���n�`����t�"a'W�l�7�>���8t�v��� �#.����h�:"U��8_pF��q���f�deW�c13�|&��22q�|��mz�i�l�g�tZ9;<Ɣ�E�۾k��������%!JG��p�j��AY)t���ǲ"���a�����;ּ���JH$T�g���2�#(�z2;w`�o^����-�3OEZE>��� ���M�#���l����m�������Uv�>s��_f˰wr0�ɛ8}C YMO*I�c&��~k1Q�˃�ȥ���"�C�Q��ca��喘�_���:�V��֬ܪ�����͈�!�3����=�&���)��b׹�`~��1v��/U�E4��N��"�ۋ=/P���3���]��B��W�+-u���)�]�ײ8H���~k�V��1I;_�¯�s-�v#&�﫶p�n�r����wU���h�ƅG��A譖`85�@�7�Re�`&(t	/�Bq�Q9V�3��y�눛���1�<8F�溦�+� ���#}1淜Q~Ok�xNoMӉ��nφ�31H���I�
�)�T�zo�B�y�dV�:jl���wv�l��^7'���x��ת��!ؖ+A��L숀��oC�uHM�h�sK6���"�e���.�6+�[����:�%�:g�T��2=d�ôB�@��� *�uݽ���=�a�nB�P�`9��(q�Z�T���O��/�Ai�V�rs�i'����z������	�D�y��حd% ������TE��r�����}��D�{E��P��p�ue�"�ڵ��6��v�'q3x�ګlwJǜ��r�I�o����LH_;M\_\�Zu`�|_�"œ4����W����>>5T(�]��ǧ�n���Ib% ,� *���|$L�^�ٕ��0-��*�˦��qL�����_m�?6ɤ_c�Z�n�K�x
�R�pp|�QFZ����y�%/~�]�<��y�ؖ��V�J�7��	F�v߃|"ϘQ^Y���a�г��-ӳ��v���mrgg0���|�D�9w��H|�w��f`v`��3�1�W��I�w�'�}���OE��:Y���ZM:������嬄�rB���1'A�d�g���C����
b����_|��f���f;��0r#U�5M��[`\�.{�`�2������bȨSؤ��p{&0�H�܌��c0"Y�l�W����k���;���h�L�ѡI�Q���x�y��uTM��TZsם���{ghl[Iq-s����֧��xBnO	�I`�\���2���c�5����sa�Yi�VW��J҉Y�'��Bc�'�_Oa�N��N��\���O�v��]1[�������ˢ�
w0������k���kצ/|"�2� ~���z1��c�>�\7y][(�5�M@��7�yQ��w$��YR�f�V\��_j{HK���9�1�x�q�tL.�]��wB����ƈ�Ro����{A2�AvZ�M���`}c>�M�-]�,c".3O��'B)k3v�v��v��w�V]_�{�������� �d˙OK9�Es��Vxyc؍��r���٥��(f�&����L�wW%݄����)�Y�K�q�T�zb��XA�9X]F���c�o�#��u�7]���r�6!�.nN�k�&vyu�Ҙ����������3IP�z���Ӈm��'�V'W�ѲBc�$t� ����;B�]�Dg��V��(%�S��u��J'o�Cڋᵣ}��2�����ALz0��'S(����Λ-s����9�k��)�2�>���~�;>�-f�ú�<`(��N�Aw�?)��<�J-f�q[�����~w���I��(�J��Wߏ��g���ܧ���a�Ʀ��.!����ϥ�~�1�*���������b�&��#>�!������,z�����5�k�cY�| \�s:�t�;�'ڰxs�Ӭ��yԽ[�^mE����W���1�������,r�Pg�	���5Fמ�����+���� +���1�r�Vw���5��rQljGh;����x�mN^~�I^@	��,��oa���hH��{Y44��u���ϝ@�mZ(/�u���T�SǃL�B�eK�w[d��L|0�\睎pu�N-�(�^,�>�[u�[cK&Urc.��άLwu�W�1�C���闏�3+����N���<w���yq����.б0A�l��U8�c���V�ܣ8l�R���e�ru3X9�������.�ξ]�Ocx$9}$��N���x�V68V����b�Lq�(Lo�����k&̨�5FkK���kvl�H��QCfVKx^{���3��@H��J�`*4�j�zp7���pqVB�ݎ��,Q̽E/�AW3;��ޱR%��V�1�,6�,���դE�}�\��G��������k�\-m=Ӏ売����l٧����+0���k�ÙA�w2G���z�s�vv�dEK�/"K,c��i��!L�)�u��l��6�
{l�9V�`x7�o~υ�f�J��aVǖnY#u�u�5���ɹ�m8p�2R&�d秹�«Q
u=��1ݝk"�iUh���QC]��&X�($&:��˷8�9�KlF���7r1!�p�J��役l&+w�p�y�u�$�NpT�����7���浠��d���KV�k�Y�l����%W ����G�e�
�գ>�A����޲�!�z�'���Ѯ.�)�5��A�6M>ޫ
�3����_r[��yt�b��OS����W}3�-�e�Ϋ����?K�o�W���n3I�/j�X�����2#�e�����ag� ��`t2�j���|��&҄Z��^A�-�]��U��ڽh��]Z��,\�Ď^�*��WaL���	I�W�uC*g[�s�LG7y�ۯv�/4�R����D���ɩ5婼�Lw�!$�U���Z�ˌ�yn�u�h�u�֗�*�d������Fb�1A��2Ӛ'��7�L%���E�W���(_;��)�i�WΜN�
���W8��"�� �c?�*^7K`�w�g&s6�3��a���L�W)Y�0�P7����</b��s�����ۃy`]�PV� ��A��X�oL�L�S�0I�+�|���к�����.#t'P�H\�lݼ�M7��*;�v�Ae�I՛�l�
�JCN��5Y��p�T�ʑ)��اv���p�u�'v�Q@o���+Lk8*+xrM���РU�)�����M��rP��x�M7��}8�Y�ʵ���ձ����|5cLj�k���>D�L�o6�Sfe��q*��E��/Uu{����=c���SM�Y�)0e��f���9���FL�X�FQ�Udv�kiV;Z��Y7N;�I��>V�1�uJëx۾*��5.in�ʜ��෍������|��/��9X�v�T�(8��j	���$B��2���W�ݻ�3{�F��(�7H���.B��9��A��4Q@PV��	�+r�x�>]�܇rh91�{�H����O�������~?�������͑���M#E	�+UT�9/!䆃?^>=�>>?������~?�����(i(�:y ht�F�A�x�r�HP�O�5W0�5��ԁHkI�#AF��%�4�4�Z&��H�CHh����/y!����ԏ���)��JQFΊ���T:��@�"��>��R%SZ�҆��(�GOd�&�)h
��v��M h!HP�0rT��I�h(ZV�A��(Ѥ*��1:�u�q#J�͐�(j��P��h��#������ՎwOT�#5��w:h��L�L]����ɵ��'U�<�O�!����x��ۡ���������;s9I��̗�-���ȷ|-�Ò�\zd)�`�Kϰj"Sm�(2l�e�x�hI�D�82O=�{�T��n�"��b�)?�Z%~�|��a�.8���FJ�c�;�F��y�+�cn��ν$c�׆�����(R�J7}��Y���ԁk��l�D�LSA�=���5x��+sz�w� vQvM��I��J|���Lh�&��G\�싇T:3�#�eJwUI��N��������d�T��I#rz�+�㗡�;���T���z0���lf8ņ񋵘��{�����!�So`G�s�h��'�-�x���#_%#|*�R�Q�o=�gtz�b��+?
����T�9��=�;�-\3�
�2��Oy�<>����x+��O��{�9��bB5BF>ز�c�1�����E��P��X�	�Q�6r�.��ׯGc���^<�S��߽ C���7��^a/S#+b�٣��<EF�����G��T�9��z^c�u[{�_u�
��a���̱�x��Uu�s���v����@���!71%��~���^�;�X��B����� ��c�]d�:�	�δ��BB���3�IZ��ꄺY\N��5��*����5�<�8���jpY��}�M�}׍7wv���n���r�1�-�#st���8���L�D`dSט��vo�%�~^o7�fm�?Y*��6k�.�̊�ƽ�MgJN��4Ë8�%�X��^>49AL?{�46J�WW�0�:)����
�,	�Y*�ݠ��ۆ�1%ڽ�]�I5��q@�/���n�'i�f�wB�����I@����J��Dwֱ���?E��	�r<����;�e��f3^���}Ğ֌�5��/�V9+`%bO��V����\�Y��[�7^$
�gj(�,�n�W����_��o&��(��r����XM����Zs��1�t"uש�B��j ����Z��ֶOK KK�Y��c��0�lS͈�!�w�u[Ԙq�u�w�g:��Cċ��N�i�!'�$�x��ʖ*�J��w'���魞��,GG�mtS��H������ydt��1��od!7�[���&I��JrQ��S)8��l&wj����j۸Vw�4b
u�C�G��L9�a��e�H��*�,c1V�"���'Ҫ��t��ӕ�m�͖[�
J�A�_�@���:��)��Wޤd_T��C_)[�$əT��>���@jq�d׫ْ�>����~f��_�9��z�Z��ś�`&����:uӇ<�{�c�c�}�g�]�s[o�:�u�'R�6GP�ٛ����ͥ��N[�d���C�O���k#���C��9�QG]���eW���P����<�'>������rw棪���'�=����L|`����l�TSE��H�ߓK%3�/�
�}�%g#m�3=��S�Nj,:�xj�Ί��q�F��q�ؖ,Ad/����yS�|���c��B���Ne���U�8�xWդO��0~�H- �<�� ���u靼@�9е�2]L�oz��d��ҵ��T��%G0��'Z��ߎ����<�R�W<df3�k��+�v�(�G�2��+�|hiT��r\E�MKs=up�B���n�-���X;�_0�(��
#-t;2O�fC6H�TXW���|А�E�!eD�?Y͛����=ղ��~��Eߜ����΄U��V~��Xf*�Vc$7�d�7���E�y\���	�H!�fA����iẀ��y?K
������ޅ��8�>V��n��N��-�+�x�ti��l)=�ܹ��(1|�3��L�L\-0U��r��&�/�L=���z-Msؚ�*��KcP\�.{aU�@�JN�z��&�)�L���}_K�3c��u�&�KҶ����4YPY坣�A��1��un���;UH�4A#%u��P���S����Y3�A+m���1ΰ��%����SKkT�枅[݆!��ͧ�K+D�׫(�9+g4J35u�,�e���֔#��x}���T@`�U�sLVav�@��\��q	�-�d�f���Ø�M��s*ҡI�G(Cu��@[��ܗn<cT�2�Z`Z�P����趐\K\�D���Gb�f�!��Z})h�	�����_F�}�2�:
���T9Y|��LG��}�@I��7�>�]�Ժz�n��k=FTձ֎�a�h��b[���5�&��?�ˈ��j@�s�C!�\�냎���D�)	9���.ٵ�=P]׊�N�XF�\�,Vt�&;�0m{	W|�h��7k��>>��Z��N�X�lha�o�i;�����r�O�Sy�{�>�B�M	1�n��ѫo^���s���^`�\�������Ϊt	�՜r��F�@�R�Ĺ���a��^�n�s������#{ȸt%@x��H`c�����]t�Y��n=�t�ј�5sj��Zʿb�r�����}�D,�` ��A�'��]�G�?*�;�"���2�WC�Eځ����$��=O�;�?�Z��
Ǆ����,��۷ ;?�t��^a���K�|2���5�7)ݺ�a�ۦg�ӳ[;f����J��Y�e���/w��}^��Th�l�;g�9		�����}89A�Ђ#���d�i �D&�v��{	�]t�wI��k��5�������i��� z�tʮڢO
������?�Ʉ>�L{�� �m?[���恷C�+��g�_݂⒐��htZR�1B���=��;�R�n���u�Al�V��`{�W��c�w�H�-�Mn��PT}��b�U�ꁭ\NޝR�9��h��v,S�[�^mz//��kzKJ�!���	��-��
�w*G'vf3��g�g9�Ғ�i�,zqmz���<�_э��S5���`Z*�P��f���S���a0=��*"����RP,!f,:/".=2�m�9/^�j"nধ����-�j�f�}�<�{6'^���0��ǫUj<��(0�\�$ZCܾ%�@~�^���Ȉ�h�K%�ǳ�ʙ��s�=��_����~�T�n,5��jiZQ�@��]��/N���*�d��.��Ap���G���d��ħ6�LJR���u�o�#�7z�91O����}�V��X�o3��
�i�d�S0U��0�I�I>9��X�J��E�5��.T-�t��OUc��kyyהS�C���^���7�$��.�V�$��Qi�g���oy��S=����ow�t���9�G�4e�lSϝ3�]�������׀*(u�L1��k���3v��E�osx�6k��,ֵ�(A��cGRϏN������ �mK�"jγT;kS����Fr���[M��WJz�e�F'�5ݦ���XD�d  5�lP�=���TG��Y;ؒ�U��n���٦����`�]�?N:�!������ �����U_�ܢ�Տn9i����bj_����w�4T'��8C<�#lYDG�d�B|�n52']P��Mʇ=̾lwF��d��j��q�����G'�J}T��طvh���#�3���˲5��}`n��ث�z[�S�^�4-Xu)�6�5a��ܼ�ɽ��O��[*��;�G(�Ҍ��fu7�m�#ô>6\/j	k0nY�S�~e�L+�Zeb���c�-A���m>��zx��"i`�M�b8@Qt9��&���c�ٌY���o9��ވ�r�*�y���$��'[{l}7:ǧ�֬������ �-�?|��~?mVmR���Γ�_q�I�_U���J^Վ/=�S���bcw%8k���C6�'�E���Ƚ���U{2q�Z�M[�d�UW}Q4N�������b�%���A�ɲ��e5#�%ǠE�ڑ
�Q�ډt��1%TqW����د�I�}@�5�Za'��|ncA.�g��q71Q~����(�.�>�����%6��܂�.�A1�0�Т��bM{Wo���=�ѥ��vᇕfI�7N.���w�Vm�h'���D4v�C k�g;�Zy�K�k&�F�,�[n>��k�p���W8����Xkm���7��<oU�Q�X���~�R�'��g��>�����N8�F��]ٝ�ӏ���v=ŷ&?>ze���2���(RXKiܜjꋇ�f�Z�rb�f�{���ҹ;:!7��߄ߧ��xeH�7�[���&I��Js`�AR�I��(��Y���]Z���.�ҩ���ƃ[0��V|}�B�k��+a �0^��Jd��i�2/��MF]�ɍ;�A���AUji]�"s C�D&�T������˶_Ucjc R��dþ��hӡ�)�u��H[�#h��f�cc�l�����	rܱ�O��wC�V��$wfGm!G�K	V�s�U��^ʏP}�%�H@셈�6�L�4g܅B�U<roUvM�!���yh/�N�5�N!w�y׈�o���\�՝29R
>�f�;b������e2�%�v��X0�t���dR�9��(q�Z�⠗��Q�%m	ֹ&0�-��'uv��y���F;�~D|O���5?B$�k+�m^�J��tֽ��O���kX�9Qy�Luy�rZ�;��[[ �MA����)!�De����&�9���A��U�?ud�*����P�[��'#�w�yh�ae�|V]^�Ĳ����� ��s��J�er�z�b��i!�Y�*=�P5dՎ+yd �V�����4�'��eY��sc���bq3���6��_[�z_]w���xU�w�ܳ¸3���'ahZ5�o���y�3
��<P�5����a�q虐t*>��Y^S�I���cB<�j|���+7�7�bb��w�E�Ef����tas���W�ǁ���?�R£�D�p��'�������7�-�U�ә�	ȴ�ٯ�V䇖 vA�%��g͠a;����C�C<�q�qP����vn��>��C೐Wq-D���'yq����Pe�@�JN�z6q�H��"7+�2����i�Y��.�����p�m���#�|�1�٘a���M��L�t�.�0M�n!�Z��݇W����x�Ui�J�/��f��a�o�����W�c�9�?!)���f�OC�^j�i��/úS�r����v��G����ZQ!0<���_K���8@����a��sI��{yyQ��~�Q,������n��/��w0�j<���d=T�`ɪ�S^�Q�Ҩ1A`�f̗y��Rt��5(���c~��Q��-A�6�|��\)���ʿm���o��%�0��kY�I�M�=\���_��Ƃ�0�sRq,ȉ��,T�ܚe9�w�=*���O'�B����B�Ez*��+9'���9��t�ŰnoM3�I��:#�-�ںU$X�d�����='7&�)rX�go]�t����e�y�8��3Kc���e8�f-�/0�hw�/�r�)�7(~�^5C¼E���&�̧����{#��4ƈ֑	�θ�aͻ�h]�Ta�Z�c��푣"ܿzӮ���+��PW� �b5��0��Z�~���S�)�t�[�]��4�6}Hħ����>�˵��X[ �+��0�|y@���'-AY�l�0�L��'<Wq�"�7���Ֆ>��1W�y񟽷	��P(�X�=Ð軷5�ȁ�n�A˶��~A��{���l�e6g����~,�I����������q���S���ٺ��h=�� �z|��+�͠�@ά"����- �2��4[�]���5I�D�о�pޚzS��8<��	��J�z9���f�ޒÒ�e8�N�ў�p��WP�*j�����:�w:�x��jY��xᨵ��0 =ŧ����Ɛy*f����T�(�g�=����^����ݐ�t�*�� t�J�,��輈��
f�yQ^�mFdd&R��A&���,b���Ū�z%=y#:�3Uj<��6Á�w=�(r�N��	������B��z�����Q��un���`2S�M�ڵogZX�	W�� �����=w~Z"�~oM�uu�N��Ol$�%0֩Kes�f_������1>�XȂg[h�.�j*�u�ދ�jΪ~��Q���3���a���+6�v��z�|�'�%�r�K(]"[�ņ�+)��)B�
N���o[��w~�B��h��G�t�_O�:�	�� D�VT�cE*Mm~�D�X�z�D�^�d��[Y��YT^wk;�^Z:��FY��S[�`hnOC���'�/C>v9H�A6�x�1.Vs���L�2�3�S���S#�dY��3���p^Ȓ�|��زO^�����ټ�S.��fckQ��F��!���}zz!�|vC�|��ׇ!L���ޔ{9H���B*����sQ;�l�w#���<y��Ϲ|q!��h����B|�=��������H�ǵ��E���VJ�k��JqB�O'�Q�1�k��x�+�ix-�2���}'�����A6��B]2�^��9�è�e�ˣ˾KB�㒏��U���b�W�������swl���c�G�2�/T�|;΄��]Ví�e�LW5 _��gX��'-m�5>��.��n��C�O���<B����0%Ct����=�B���k��D|}��s�$��άFi�˯e��*\�_�xum�.Ɯ>ݵ�X��eH��/s@��7�
�Jh����]K!Z�|m_s,l2�j��, #�ga[�L]R�k�
�P���΀��7��	J�c�g�Gr�.�rl�����i�n�b�F!�)�'�.�Q�{f�[�d����?-	m�-�\�����n1Z<cg�
�\�<M��z:�0n�L}�
��ܸ�����.f��0�;�i=7������!�����]�թ%�R�E��N�E��-<�e�[��$v=n;e�v�cZ�oT��<ܦ� ��^�U�P����Cl'��|Ւ�m��}��o2xa�w��,�u^�����E\��بS�\Jn�����;A�Z��Q�$��:cYf�I\Ռ��nci̥4.����e�7k�R�wHp$UĻ�
 e]�2�5��LD?�閲E��j6�r� {ۊ�ہe�0CbFb�)�Su-jqᔐA��6˾ڛ0]�.VK��l�OY��n]�́$-[�e�P��fh�g��[�����ܹ3��Ft�����aj�d|����B�]L��ܔo�Q�>��'��y��鼬o� ���|�*F�f>�]�*����q{r��vV�qG��x�_J�ظ���ڶ�/���{j�w����C/_�'�9L�4a,��`�i�*��
�U���qڨ���pZ����fÈ峈"�;R�>�M���i�m��eܙ���q�ñ׳�i V2��2!�&���!��{5�%�n�p15`ruD>�SQ�]1�k$ܚ�"N��$9NKsf]FUL���O�{2�Cv��ɡW�۠�@�r
�Ti�]+u��ڗ'B����P�Ĝ��[�ov봱�/E] Mc\z�.+e�I��u,,�����J 뷩PQv�ؐ�u��t�+��e�J��]}6���i7�d��oZ;�N�]��rr�N'���ꎓW<��i��'��=��M4�+�;1���s4I���.�n��V��Yd�8w2#��:u����m��ܧ�un'�*O�������+WV��g^o�ۦ�$�T�i�[5��f�����9U{-�S�e�6M��Wb�[����*��w��V�
i�����L��Xx������5�n�n���85�q��t�bTf<�3���ˬ����^�,�3z�N��?��Uu+#��X���v{�Y��}�D&�q�hr�:��G(�6{Vu5{x\}}��e/e^��4;y�qԭK�$V��[k�Ʊ{/Ch��W �.�Ǡ��yB�\`L}G&�I��#e��Qk�T�C�ju�Gw�'b��.�\W�+��6��a�|����O;wK&M
�k*_u�3��	c��-�[O����//n�I�� �F��9녟�޻�}�ui�>�z\��=$m�f�u/���`\p)%U���\=� ��%�)�d�B���h�JL�����~>?����?��������}l50U|��X9?a�B�N�O"""��г�����||~?������~?_�Ґ������4�O�h�hJiJ"^�������hJC�tRҜ�͠����(���SI�CmU��9ADTDW���A�i�ƹh��F���t4��h��*J
F���{�AAR{��y��Jk���F���.�0IQ1������Gw*[�V����.�D41UQ�4��KrBU>ܪ���'�5�|LժK�]N"�a� ��E5\�PG��!�Bj��������T�T$KLCHh+C)TEG.A�׸�CAQG�e��"A��@�ێ"�V�}L]�dw%�ͨ6�.������^ƴ�����j	8��]e滳����M�"��t�b.��k��hI�0I$��ad��@I-�ə$P�ˌF�$"�m8�	���~ �~�Đj��i�4���}ϧ5��V��$?����C���I��k���_8�Tm�^l���&�any���fh�]���u�z]����Ęu���حߕbP�	X>bO��mY��%\���S�&z��d��{��΍A�c�Œ���$d4�ɶM�aL��^��X0 XM��e���i�W��8�ܯFgT_��
'$yQX˝'�㰂zYX�@uiU�؄��V�NlTk��.}��m�%����b4e��f�ɏr�: �Z�h��uks}bԩ��ۓ�Q	��:䳼I���Y��̮��"5�0d�˨T�7�8H�����2N��9�h �J1o֙9֬������Ӳ��l�'c���������?J�O/zD���2o@I��z"�҇7;�kN&��C�4)�+�����~́#ZB�t��#�E�	d�Ai.ܒUg���3�\�9��Fcm�1L��g�������T ��=S��N_t�lQ�;!��$UOj�&�D���s	C�xj�r��*\jO�ø�vC�Ϝ
n����n�p��R��l��L�ǀ8;T��R9�`v(��)K�A��T�)����G:��x�
�zԱ�k�
���V���#N���- l�%o�7��IY���T�4����В�ٻ�u���_'�d@��>�LL��xkH�~J8E��;�0��E^�`����8�v޵��Ĵ<�[�De�^����ha��.��,(]<�n�k	j��W�����7Tv��k�`����(0~`��eb`c���{�uŃ]+^�PK�X����\{̡���wC��a�/n�F���␀|��`�4�~O0���P��/u �]5���8��ݷzWг����v!��R��	`dl*�W�zA<<�Й�2�_���8�S�\�}���3炙W�I���ȮSӰ�0���L�:"����^G<��\W�>�!�=�܍k�'Lݨͪ�#�7��@q�a�m�;��0i�e�A���x�������-��*��L
�"
��π�8Pa�1x����֟^7����;#ܛ�h�_i��P�k��v��sB��-u-�F�d�|�Fd�(��/j[�)��Ȭ�(8��4�m?#gl6v����¦*�E3��@��X0Za�s���l�0�;��&�W!2,�����BT�Y�+\�n�V��[�+��LՆZg+(�vg�c�t��s;P��Q����x���0`��Geؑ\o�����0^�1�ʄJ����c�׷���{ƓWؾNS�
��ğ���Y�닝���s}iʹ���m�z]3��+�Fb� �׬�<H�i�lܑn�I��;W).�S:k4�6OW1�*^e~C���{���`���Z�/\@a��~z'_��I`�~t.ܐ��T�±M+J�,��{���"���;��~����@x�so��aU�	L��ĲOk����0���p�����7��A�l�;ޞ/jf���1�/���
G+�iN�W�"��J.��[�\���6��6���L�=4_Z�������D&!�q��B��4��Օ]v������}fr�n~�ܡDץ����c����@���}�|_��=W�������:�Ñj5�x��T�w12������A|=˘�[ho�V��A`ZGizD|�Ķ�zv�2���`��z'M��Wo�l������.�R�8���`�φŐ�v�a�a��Q���9k꫽��D6[����iun;is�Ρ�Ƨ��?LU�>3�k�G����h�����b}�K�&��2Μ���vN��b�1zr��Ҩ}~Cx��W����4^���[��}=>ھ���=D}�B�q>�3z�/��l��Ռ!���H~,���i/��Ѥ�FGZ�}�@��؛�n��Fv��!��Ʒ+#/cp�Lӕo&�����l-G�q�_��]��bH�8��N��*9��'�Z�������9A��
O��}�8`��qZ����`��=@�c���ؼw6�q9�*�귳��/������o�1+��@�}��x�=[j�/�^A�}��� C@"_�?ߋ�\/�U��~�9��oO?�u������L{�$�Y�kă��^1*⒠X�2|�5��j~�T/`/��sr�F�O���y��su�^\���j���3g��κ%�5��+ʲ������y��`��wb9}�v�k��wC�;;��7�Sm���ɨ[�j�~�#ܮ�Z�Q�B�+��b%��b�ȵ\К�SD��	��<!���:kS]4<�����%��5��񢚓IRy�[��ds��w�kb�D�-!���� +�m^Ǧ����ƊT���Crˈ2э�	훭�g��CP��@hY�ro�@J�} ]�0S�=$oR���b��IeF����B��k\ƥG�u���A�A�g�����yȄ����/|��}���iȁ�n/o廣�P�%<�svi��82���(�s�����χ/�,�[7�7���-A�>�Z��ֱ҅�P/�_�U��y�r��/�}� Ư��,d��W	����leDW�IP�bK��K�L=4
g��gU�$kp�u� 9k8)'��1yw�;�d��}]�1�b�O��|эWo�Y�O`� =¬�<�X�8��pR�]�I���uD噄b|���p�NW0��JO+��2�jYK`Bq���]ʡ�������Ԍ����(np��]K6j DC���v�@Ԋc[*������t�~��cZ��x�+�i}�byI#y��1�[������h_�9�+���~�=]����[���e*�VF����Sg%���wSE0h�scH�,K��ϒ7�gJN��ŠvQ1@sVӖ��<��Џ^a�y�Ր��h$ڠ�bG�):]���n�:��dqx�e��S�#�*� �_M�}��ǩ;���_��KA��Ϣa���k�#5
�S�2cZ퇓�73����؄���އ���<��I|k�P�-?V�J<ğd5n��U�!
��aj^�#MuW�;�;����q�iqzY��!�RY$5$d4�ɶTG���J�x�bks�/��Ko/�U�����D܎Y/x%��ԚK��U�K�a4�mkni7[s�'�������*眅�!6d��>y"���4���5�.ixT���9�W"���ղ�RV�3̆J��lP�I�J�gu\\�$�vM�#r>�G����K�g�U���v�(���MJ�x];؆6q��k�3�oHG�Cǎ���E��W�B�s2WKa9��;�A�l�6�t�u�
6�,-
�Gg������es�"]��]��o0n윛�7�Gֶs���+7)�{�$ZHV�
ky�@�웺�7���i}gso�Kj%Xn��x�m��5S��p#!�����z�m��U��C��b��&�H�IZ��뢷�t6zXc��T V�뱖�K�{y��^(p�ob8ĜJ����4�wI�t��z�*E�Yb)>��\]�I��	���8�z���w"V�`èE�=2�=n��'��i�*���Bac��]^�lSziS�r7�ڶ���L��"/{��O�;��Y�{;�Y��4��8cz� �o���o���&�_N�Wk��FwoWk�Ʒ�ݫP�$�|��K>_8)����b�/�U���N�.0tqn�& v
��nd�Y�	�X2��m�'"��|���*����n�	�$��X��^n:����D�\��[^��i�l<=��d��S��m7/��eK���q������Z�X!z�����#����gt�P=qBkt>4�v�����̆�엔9�e�_r{��NT9du��B�f'���뵜S�<S2���jإ� ̙�k$as¼��=�����'u�4!�y���ڸ�+���ub3O&��Z��B����=ovs�,]��`�� ����Ѹ�魋�Ȯ��)�/�chk�̕rvh��Q3���r�jni�vKǁ�XJ<����Ͼ�������%c�� W��g�Ӯ�x>h�F��RiI�;W54�E[8��n\�8�8[�]-OU��Ul�YrD�lD�~rdt��k�$�^�ieT��f�o�ޥ9|R<w^.�ʸ���6������$�O�����{�܊����S��3=�����P����[�$�6<���������'[[�[�ݩ�D����ղ/zM4QZ󦎢��Jޚ�C�pl�9���G0S�(^���(`r��b�3��g,�]��.2X�}�˚ʝ앂��횂7ύ��0{�7��o0[��ceX���JS�#=���QҚ��4��H�����V�a{;��w�`�*�9���Nȳ��1�-t�Jn� z����WP����~G!�q뙳[7޳y�ε�(Q"�1�A��!�Xd̠����Vb���w|�_�Y�sj�]O�U��9.<:�g)e���F����������K7[Q��=gv>H���f@`��(	�����0"�0b2d-��5uԯn6]v���k���5�ҦW��{`�����*b�3�{�]�滳;Y<g�#�nFRl�{˩�K��H^GG�S����z�m֕�ϵ�-?�-���_�%a��J�����S^����4�N�<�)���NL�t��������g;�]�*W&�z�u�$f��b�F\]��3��oz�W^l�>�ƁW[�.�d���D ���������s����r�Nͺ[��}�;S�9+���;	8:�R�Y\��6Y�@�X~�w7)hX�T6b�F���n����r ��EI�z�̑sNd
��h�s����r�����1�jP��[-��
��Vat.�9w#U�X!�yQ;�q��%�������G��:���=���IQjn��+B�n��ɦ�l!�\ё��^Z�'���~[�o��?���cʙ&�Ѹ�w����1㫧���s�����ds�U�����y����Ž��郞����k�ΤU���cs�:��K'9��!N�ɊXw���x{�½�=�Ծ���=qvNN�U�V�}��_�� �d	��j�v��BK[��Wm=���g.�N�����ǰ�l�ٶA�!l�6=��2+So�L3�Uk��w��v7\W�6�¬�����d��n��]N���:��^Ӵ$'ۃ9�gA����;Ϩ�.��h��+��m��Kr���3.n���u;���OB��1�U��Էo�d�U;=L0�m�N-��>�j=�7�����Q�X�㤾��O�P�vP˝���+�e�憸��F�u�Ѐ�=�rG��^!t��\_���z`�e1]ި�g��E'w������V�( S�\��7��_/��}�q���|C}�R���T��A<�t7���&|�FC:#E�����2�Z��T�~�X+�w6"�PĊD����/cWE��h�]
-�nh)�6�6�;��
6���	V$6�o	TÆ�hM$@�q��X!�ⴅ]_�<���.���#����)�9��
ۺ�o�_Qư�2��,�) �	s��O3;��$�/^�&S��[oc̠N�aU���x��gEx������ؼ7�Ʈ*�Nz���=�f���)Y���#U��a.6Ks�X�cV�T���`�!�TM����\V�� �o(:�kI뉃j��==�6q�+�=���+ޯ���f�%�e�p�X�kȣ&̘z���gMV���ϻQ�r�7U+��4�&��Ԡ܈HV�Y��>��{�p�M���ϻg�n��`��=ґ�n�̑tB܅V�� B�s�`����bj�k�Nd/6ؤU�8�Q6gd6z������1L�"��:U]��^����08�T�h�%P�q�td-��g��L�׶9�on4Er��^|f+�H�Su|�VW;�iB4�t��=yR�P#9uʱ�r�etl���a�u�j!)�ȳ�T7�*��b�n���s!��/;9��a�K�D{�P�4�/z�������7�z9�ٵP1U%_pm֛�V�v��T�Yl��̋��`�\�)p׹O�k ��Ys��H�f��.��Å^�(KYH���Ǵ��S�������
����G0n��h�Y:�J�8�U�f����m�Y�ϴ�Ċ2>[LM��%�q�j.�݇�����gRAn�J�T�f��4����j�;&�>�8��n�p�E%�/��m~W���-k/�8���T�l�;v��$��K�'��Omú�MUv&���]�P�{)�M
�f]�_E`sj�u%JK��޻ǒ��H{]e������V 	��1�WE�Ҫ@Uv�0.j9;�<W1���3���r���5������T�'x5�q�y�m��a��N��v�����K*H�LӒ'
�>����[��qlߏ^ߑ�
�c�^̸i�c�(>�؞d���yǀ�nr��U�&sj���۠��:ȕm*�;e;���Ȥ����:�澗RQ�[�NK�x.��N��(�*.���[�P���;���ۑC��J\ �c'VQGp�8�̖��+$���tZ�&o3qtR�Y�U�@Q	0S=r�-�����:H�9J��tiqu�u���3�B$=C]f�S&�Cȗ=Ha��N\�7AU�a�ĻYl��	���6�ź��,w;Z�=�x���g:=�۫�P�0f�nc�$���%���P�����X�8ýbկh�u�ڣьV�"�B�KI������<�����ځX�n��z�8�a��^�gσo
�>x�IO�����J�׸f_k'Eṕ��j��}�s���:L��3�&+�A��)�W��J���J�Jݾ�]q��q� �/>ِ�,-VL�d���������A����'�r��>�V`qt�Oa�Z��N�ح�I�$���yb�j,��-M��4V�i�ވn�In�].�<˵�]����`�L��g(�3��mV��Ь�-��Ю@KP���*����0�ٲ��A8�!����*��a�N��]�a\4����/��]"l�u�;��=Mf�E�D�Ze:挫ں��8�T���Zn�K�ۇo�����zԩ��PV�
O���v��۔MZ|��^�Ӛ�
���f�٨]��峦^��C^7��њ����W�Cr��s	���C�9Z�tC��v��t(�y�l��ݾ�Ö�66YJ���Ơ��� ��|���ѕ�q�p�yR��6&�ԅ��U�qY�<�N�x�5slD�W�h���7B���E=��J��.Ol�XnP[��.�a�6�oj�oFeءtSiʃFu�G�F��tㆃPּĩ���֮d������-��*�k�����bϜ�n������Ef&X�%N���O�Ӄp���tr��d�f��]�ۻ�oWP)+���F�!+���}���<��*+�ĥ>�K�(�B"����9:Zj�jj)
&"X���)��5A��^�g?^ޞ�o������|~?������%2��j*����
�>d�B\�uKEQqPU4���z}>�������~?���}�hm�7�0�+����H��"^A�&��� )j���h��9:�����f9�r��UR�����"hb�P�=Λl'D�^��M�d9]mRQEIT��QE�����T�AUAR�F�
*'F���F�]AP�KT�5I�i��I�!����h.�����oX�Ts�9�����'SȮI��h��n���"���u��؊�"����f"�4�LT��h�r0i�q��(�)���6�OQ���SUU4z�(*%�
$���4TE2E��QDDEQDMgp�;�xᑄZ뢬h��ͻ��3; `��%Xk�<����f���Pf�݄��׼7�2���Lek��q���g� �~����zy�Q6��=�<d=�n�o�����y�(�@@��i�-�S��*����s=�����q{�Y/����0�Y�`<e��@ڞ:��vn�0Vơ��U�\yo3�-�>&;��s��g@��_�m9����w��*������7O	�$q,pN�?F����	��4Ջ`�b���uכ����"k���+CO3�<�J�É�~���*W�t)���LucՅ���At�f`rXk�]6�%�{�a�4@��i��75Ы���*����}���Q��j���a��={������+�@)7 �]D���t���H��kr6N���uW��j;�m�!r�>n#|�#	W�<Ʌ2J�*�YhM�v7�v���/:���FГ�+3͢nJ��) ]g�%w�����59�dD�u�<R��h�l�[�X�'R�Y�����zjev�.Ʃ̮ͫ�N��2j�9�����:�iI�������Q�*V�뤍ut��ҳ��R���Ǔ�g7���mIc�u��kT�/a]�Vw+9��${�D姕c�]Lg��  ���7y�����#�Q5$(�@�-͞J�4���&B��k�d9m�i�f��i6��̚�59�P�[{��;�4
/��z��C==�3���&wWV.�جc3���:��w�S���R#;�9\�n�z���ǌ�A�����>��>'t���_n��F�(=��g��Z��U�^ol��Χ�]�u��{����y)�}�#��dGS���V5�M�����b�r��(׌����QzOA���ƾ��h8�P*�-�_��w�}�0��`���/I�9���`o6Ԏ���h��d/��+ݾ�~ݠ��H.��f�Ҽl����D�,b�4SZ2Dv��]�ۧ��O�T}�2R#�1]Acj�Uɧ��W| �r��.�N^d������n�hn}R���Il��#b��M���B�5O�"zq��A#u흙��VK���^�ݥ�m��N�=-N̦r<����J+�^^��rB�}ǭ野�[+�Cs^�/B��bK��+D=�{N��Qd�0�/��F����ceۨ�`]�۷��8(��n�<���x7�����s�2f^�n�`#s��E��G�vV�][ܯ�	`DٻZ�^���;䎴��R�(��P7^���m��Ce�^�}���bU/>�5s:�[^EI��]r|{2E�9���)cq9
�6K��4�4��u���O�I��e���q�k�T!t�9wu5�UU�T޺�#:���O���r*|���_.�t��=��D��3��ڪ����+�-��n�N������*��Ng�߲��݋n��mr�2-i8�մ	7Ǭ�1�m.���6=[�hÙ
$.��q��{��>�>١��>vך��D��q���L=��7�@��M��h�P��ji�s���㯴R1^+�q���L0~�ΐ��~ɈYy.���=�4��A;	z�y��>�H��ℷmNN��r;U�X�:��4�x�9@����b6��~��_VP�N;��8FO?RL�1�WnU��M�]��cRg�v�U5��=+J?&�}�}o��C�_��㍣��>�:b�RS����Tl͕7w]�]x��g�k�eK]C{O並:L��N�,�$5(���gE�HM�z[WwpE�#{���܅Б������}uW��}�q!��gv����}̅t�E��l��%��*:�����������3Ś�*z��ݾ���2�����	����Ѻ���`z����t>_f��2۱���t���$�o��;H@ϦF. U�O����˿�k�L#��ɫ$�Gq�1�
@��|��	H���,��Ns���S��Yl^'f��ݱ���1 ��P�����p���A����Ԝv�)ʹ�s��u����cѫ"�gge?�c�>��S�}�옵�f��A6��]�T���m{a�[�����a@�Y�i��9 `��~�����9�YH��V�����y	���<<~ٱ?��?7]���i�M3�@Pm�[�=Z���]=�4[�����5я��QS���R7-��7��=I	~�	��9������u>u�.�K���"�1��;��ܠ�ng�u1#JmcC����cnf���U+J:1I��+��K�����GYƯ���F>��H�9��2u$�.�*塖��w��S1�i�6i'G���1��Oa�R���y>2�h��K��B~����5�}�v�ș�*���ڻ�"�y�����#�//�}�E�.��j�z�6�IZ�q�\�[ϲv{��7Dmf��9�)����E���K=���z������"�w�KZ;6�YM��̼��lc���t��D%~��p���U��2��I��3R6p��zw��5��$-��W�55ߑŞ�Tiɱ:�h;.�9q�h�MU���>;�J�+�@�MѾm��7������̜�w�d�UnVŭ�2�3��C�F�t�.����/�8��=��|�5��AR�I}��ҹ���k��8��C0e�=�d���%�v
��ny�^�9*��{m�{��`̀��Њ��n���Q��'��D�%�SN��
g$���[͘q��fk��E&�������'�9����"$u����g99�����[oz̜�Mܬ�����X�!+��ɯD�Mf�%r��9��c��
#Y�F��wGm��v�����J����8I��df�����a`��+SNZ0��l+��݆M�`������b�3��wkڙR�ߍ�W�7voLRU
aŘ�:��n�ʕ�v�r�S�ܻO��d��i�2޸����X믫|<=u������v����.YT�(�u~��^���b��˞�f�ob\a�FwD�.Kq�`6�%$E�*��;5u4�@�g@��p�z�#��o"�k�cY�����܂�Ѝǒ�IU˹��e4��n��3��؁]Qp{���9׹�W 
� oBK�F��H�����L�S�n��z\�v=�Ky��~Kk����
��lrK�߭-��D��k�)�����f�Y���y{!�dy�����d�ղ/zM��Ek튗���l37�4�}7�Z�Չ 8ٕ���b㟤0� 0[��dhFw��v�d���QJٳ��f��w^��͸�N�G����h���2<4N�N��l��}��ϲ��K��w�TT�1r;XZ��w�X䶙���b���.�2�����=J���n��*(�'h@���:c��'��}�0��+�`':�~[��״7�9�S�a�͆�%��Gt���L�Pc����]����{8��+���f��i����cvS�W!�H�U�rK	*�2h�ؕ�;Et/�����Ec��T	�x�ҍm�u�w�z���{�yZ>ﺷ:�m�P�Sn*��<��+E���� c�~��s/Q�zdoWf�zѶ�R���i������W�`�����_�=����IgT^�B����$F�SSVc�����c5�7����0J��s����!]�%AK�W�qM��]V��;�pwvA�%ho"��S�Ng%��D �R1�%]�����̪ ��f�p��f���6�JV�y#�>͵ ]2��p(1-�7��,V�ڬ�=ƕ+J1��Y�!0�I��̛�r������â{��m������+��L!v�
5�jW�J%]�]3{�ǎk����;wd�q�g�̣V��nj���U"R�~/�k$G9֛wbnI�c�w�W�x�w8T���-҇�ө�� Ќ�T ���� ^���'=�\{so�|���i'�P=�|ُ��C3�B��߀Ծ���_��9�R�rG%��]�ͯ��1[�p���S�#ȭ,���ҷpI��B䍮�X�)u�h��+���܅���3Hf�w�4�k�V���YoY�F�p�d�NՑ�:(U#|�%�ߨ7��Ӛ{x�^�cz��X�JtZKa�{вT���[�;˥���T��K�(����&-Ⅵ�DoOU�Z��)�>�}��@m�?+�/z=*�������o݈9�cO�Ft���[�M-�R���|��N�ҜVsK�<�DVka�h7Ű8)O�n=X�7q��e��t�َM���aM���z;���PR���|���������v��S�":��Tgv�C�vO����g�A�x��%����
<ϵw�,�9	��a�iN=����ʌ�����l�02
cт���4sjO�*�k6��GmϪ�^_D��	�(i���oա�7@�ňRs���L��~?��Non���^� ϒ�
ឫ��Ӧo��ɫ��w 9�)g�����S�"mudצ�%�p&��c|`�������-�}gU1[z��ؐC+�-����N��oW�ZD��*�|o0��{b~~yS�B���#����Pdt7u�XW�N�j:�"b��Y�.Q��ʽ���X���&k\��D�@ŏ�.�L�˻���Sm�o����x{���)\�W�4;Oۅ��Q+$e���$o-�]�B��ap���kg���x��͑v�[uJs:%�Z�=
Ȅ�V�8�NN򥱹v��T�݂�f�����(�rv����?`�ݑCZ��8��y���Ód�� �yyȯY1��I[rEXn�Q;���R���26T*s���s�c&��anÄ��W"4�U_g�Ͻ}%Wl�65ѕ�� ��MQ^-fa�ٓ�U�o�0�HD�Gt�ouq��Jk���H�K�����qY�9���f5ik��u�٭h�vC�ޠ"
�L�=uCyr��Gх
�=��u�ETҥ^ǺX>�f�+��u�"�O�9��Lde�ϳY����	kz1���W��'�Ǻ��W+�.��A��7ͣ��ޏ8��m�����Bu�Wd3����J��'��g�NL�t��f��1Ámh �.��������C��t�(��kkc�]n�T�Y���ܽr��}��Qٔ�B�r�0Jhw����Ҹ4e%�[&����E�(�I��iwi.�
32�&���+\����D��l"��1a��ī��$�Z�����{a�:6�TI*�7b���[�I���F�r����ꁓA�UN�.�*��KʻƁ��]��{jJ��g��J;�0�Zq:�Up�۩&^�"zn�xq���&Z^���Cp����6����ޣ�N�{�gT
�����sZ\�cCk���M6��f��o��8��P�� wg����>dVQg����p�_zN��GG%ve.Ɛ/-M�9�6Y��=c�~�Vؑ�m�Y>��V��G7b{������F��VW{(�ʚ{�
�|��SPu���"~�����e����p����R��ǒ�!%M�W�]��Y�7	yw�w��=��H9c��.S���� oJHEdi��s=��v�BW�[��=�U�T�"�=#q�#�5W��gO$���Ҹ=������̝��#36Gm�@6�S��f�+��*�k�᪻�8U4N�>lܫ�{���C����3�x���ů���{�vvi�C��h.�5u��3��bT�g�����`ibV(���(����z��J+[=���cF�Y� r�܀���t��C����=��7�yո�~s+f��	��u������ⱉ���Л,WX1U��Ս\�2�+7[��]��.�;���5���� ȯcz�x�S69�ц��zN�S�頳�3K
���T���+v�f��v,'�=�T�,�[qY�����HZ��Ĳ����Z
���]���]�-,���Ưq@��p�o:4�� �eJ�j#�M���$�)�7C�������o��� ���xDՙ�x�(;��Zk����}��y%�j��6ѝW��)�3ظL�>"�p�2:m�#C�ai]���X
��c:�okS��fR�h�f�NX�L�`i�75��*�9N��K1`�2�1ή��R �,m1�j[X�;�8��Y`p��y�e�\��PЮu��t���t6s#`U�Cz��y�e�ngB�U��/&=2��q$UZ� (������bC(u���$)B������}Ɩ��~;�X5��=WIi1�3b,�޼��]�ͼVd(��z�}(�'mP/dj��iV�Z�#ʦP�5O\)Y���K^�\��4���9j^�o{�E4�WH>8�:���������=;�m\O�x��Ǧx���'8dn���Ƙ�;��t�^��,ԼuQ�{C��+��9s����v㴦K��0U��8���f�u�̭�[�r%��-d,��r��v�}���� $�\]�jk��Fg"�A��6��e%���ЛCT|�5�!R�� &p��ǚ� Հ�O(�ua�4���q�Y�G�Zj�kJɓ^K�.���K����d�r(���dB8MY|������>�P*u6��	M���>'N�����òv��DAx[���s�Y�S�lM�,�<C��0�;tf�/hCB�K�&L���>ʾt+8�W�Fe_��`�p�|�x�;�Y�|��C�{�np�o����LF��D��:t�1�C�ݧ.��,�2���MJ���W�5yD��u{2@��fI�ڻY�/�2Q���y1�:e<�|B:,�t��ЇlF��n���[�Cфꤦ'�����q���"n��'%:����Ff��
4�ѵ݀.�9�OT@M�9�F���c���(m�wFbuѷ��m^]�n��Fm5�Q�w]L�/pWtT�Y]��^&�Lb�))IԳa&�z4( �V.ٹ��ާ�.M̱Z�d�d�
�n#*�B��2C[pl�2aFM4m�S�L�Kp�%���t'*Y;��%��
��9ٙ/f�Mğ^p�:Nb�MJ��HI O�Z�>F�(�=N�}ΟS��.��(�����u�9�������}��o��}����������`�*&�Z�(��:�Ij�&$��Ø�o͊/��?�O��=On{}=��������o����~�1_ri)���4U5G�-5U%	@_-T�/�)���*���b
&����`�u��E�TE�	�#�MSD�s4�D�%D�zƧ�5���"(�&*O{SGq���10{٫�G7\�TK�i�pj�"���4�� ��"媮X.lOv+�E�[�4Q]�"��`����*
:؂�*$�{�`�("��#��Ʀ���QIE4�����lj��s5DU,�Q��BR3���F
k����9���E�UEsb+�m�4w&��������(�&��E�R�U1�ӣ�z���5I�h�"��mlU�?xbD�i�0��b��E�'��.�����,�m�|�q]b�OT��O9螺w�<ճ+;��/5��4ήi��%DV]GPⱺ�t�(IQD�M�)e�	N��[p��HaF��2�B"j��߈��"��)�J�r/2VF�
�{�k�7w1nE�u�K����7��Z$ϗ��`-���
�`����V��Z�3��kQ�8�;i$�VQH�y� ������7Y���8j���E\�yY�����@�8�$m����ʳQ
�L\���7��蜥7�	j�0�x�'a��q�u��?(��t{�g(���=�d2|}kWKRJ!6��[���b���A����|	�hJl�q��z�s�ͷO�E�ׯ��f3�W֗���\*��gwG�a�Y���3׷�&uD��v�i?���J٩H]�W�R��ΪתWX�(0��WG˛t"�'�f&���	^�X8�t�t^j��̣Pse�
�Z����c�<���l�\VQZ�2��;�a*<$���%rBA�M"�c^RWL�l��Ym�9�+{g� �o(^�y|���까�B��(*Y���9����n�7�Y�WM7���o1Æ�S���k,a�[�2��;\�@y;X�Ĝ����w��|��-�`w&�dt9�[��7�;j�gW�7tGE?��̔켏F.���;�G�N��M,���ko�ޞ��8��/GB6��=��G*W8;��z��ۦ���5�pDmPuw�.�7g]/2~P�F�	O/4�؈��ù�cu�˹�nf���!?�������DE�@�r��3�vkkf6�Ź�b�sNb�CJp��?Tyq��q�LB��	���<{	��-�uUƺ�Wgs)����ƽ�=$���w͘����[�=8��d����ηg$��-ٮT�_�������������['0G[�Z�h�}�C�*DBS�����-z��P+�v>j<p�e1���S۷},�A���8���4:LQ~�ʯo%4�LP���W�FN'���n͛x#)�z�!� 8H�6��Tw����3b��ķ L(��Ջ_Ct�;�3dS��o�]!�� m�7��ξ��Zպouȸ���^��UPE�$��lϺ��g����@gVW�e����5���j�ō�c�Ľd^K ?[�u�Bs
�~�iS�KM�Hoyf!��
at��ӏ幆*��]����=��5��b�%����p�;.Ko���F�y�5a�9N�l�����K�=βWLR�33
���avݻ�{������p{ØO���w2�,�#Tt�y�ρ<�t+T������4�������ϩ:�)�|>�����]
��D�F�k��t[��d&9���O*��o1�MP�F���<ﺢj�f@X���I�P�V�\E2�O2Ų^$KnE�����}J���XU`�z>�ˊ��ɋ��-�� �;�;tw��j����]�v.���7P�.��Gz�TJs�x��	��ߠ,�hd��n-"Y߯Jn�=LzM���oH6d���s'�4�M@ z�HkՆ�����r��m��p;�ϛ��la"��$�]-�uݘ"�nѢN-K�o��������M��ߟ[�f+T�(�H��~�@�~�<+G㞐�e�C���Osw�?R�\j�&G����*��h�t�^]+��+K��=��(=V&�<z;v&�S����'�B�]b��W������J&�d�4��kn}�{<p���غ�/��Ҳ�9Bs��/C�^�i&��V�"�--�h7�a���`�ls�6�F�Qb��r�q�����=f��R�-��]��w�)��e��7�4��f�J��8t�C#�}��匚Z)U���ZG�����8���+[g>������׍��]��}[�肧Zx͞��B#0ʃ ���`����;y$�T���/c�,�m�����\0+��̢F�~���9'���ݮ'+�DV��i�{�)��Pޚ~�F�goM�b�^`�L�^����a��p�j43�4˦���� �<�*t�v��"�Ψ�ӗم�
b0򘕗@@*���p�%ضQM�K�`����c"۵Vv���ڷ�*����#:^����ۣcז��'Ę>��i����׼�Pw��ƹ<.y|�i�/>B�RV*Y��9��x��n%.~�k�f��v�p�1��݃���=�?5Vs*U�AB�t0ٻ�\Lu���\����7�����aܥs�j
Uߥ��7��2.izF�E��p�Ҝ{/P)��7S���RP]�PɎ��<��FU&�����s"��X�z"X�6?K�S����aq�8��>���9�R����A��J"o������E;���q�ϖ��E�,�Ȯ䫧0�n��y�:y#���9Ϋ�z\��D|����`�3F�7gQ�M�z�R�C�'/
y�su�N������|�	+Ը{�v��
�%	H$
$�߽��S{j�p��b��Z\����:Y�Vۙ�|�S>��N��˾��l>�h
��0�W+k��$��#^[=w��;��;8N���I��l��s�㫼���¸8�9����dd�J�8�Y|%�Wۗs��>���=��6�`Ԃ�Ybu?��>�A���ӳs�	�����r��E���ڊ$������a}��#�^�+�W+q�T���|��*�y�+΍�gֳ�`���oV���O��c���82A�+��_aw�:�t�@�j*S����R}���q	4w�p��Mo�#<�B.@q���e�t��݊�iQ8����d^y��/y�G����wP���{�L�@���lȊ�'�-�z�Pc�W���~c�.@fc��ۚ-Ns�_I
@�g�A�Y��Gt{5�#/+z-�?ܭ_�ȏf�����f���`Q���[�Վ1ռգXE�qs:v�yV�sFx����
5։�'��N��\��߭C��sa��TNw�Y�����:]ƭ�ڨ��S�e6�V��9V��_dGp%��Gv�μ �^o0�t�~�wx�sD��r�ӧ�'E��S�6C:����KK���vf����5wK�v��(��7�RX���n�c]/L�c����1w���-uas��X�����P�R�׹��b�&ѯ$u�6��2�8������7��v����L�B��w2fɸ|�B��)A�z���V)�\"]_n��Yz7&ȹ��A��
��O�κW�J5v�1�w��	�i�[���fL�˹�ng�l�/���V�^���YuO��:xn�Gww�lf�%Q))��Q�u�����_*�O���ӹƟ7;)�ms��UIXn\hy�������CC��zk��5���Nv�+�Ѳ+Km����('�Y���*GsuᶏB7��s�-.#����U� ��7���Mr��)�ܻM'h�/SY���=w�F*UYF�e5�����Yn��yY+��!V�ؐME�B�v�ʿuY�8N�Q3���d&�F��Kh.��Żˡ�-�8RѯvJE�x���mkO�N��%�A��Su��)T�S�v.:��g�����r����u�3;���+��#^a�@s��BgT��W0�쭾J@��b�]�����u���w��ڐ5*E� ��o0H�u�m3�����'i�Yz�v'e>woQ�ʔn�2v�n�}\C�#Pj��N�a�U�&`foy#2S�n?_�~uO_�Uo�����h�s::"�K�y����L�_u�ӛ���y�ڝK�%����<�D��S��m�m�2��l���B�:Þ &݇���8/,Ď�D�"4�X喫-;�D��z�;f�/A��s�B�lkݥQ5uC3#���;;�2TD1�3+�`L	�2�X�yCw���z����ӧ}k�t�<X/�	o�.�0��ۻ�/NdTE#�U��3��xF9��v��t���g�vם�e�	e��Q�ꚇ��uM=���ح�-�RR�ɨ<���t��5 zk�̺9^�L*�\�L]�V���Y�-�E���xf�4����gMr�xy2��Oi�Oh� *���2��Rޔ+zmu8�6��PE���u���s�J]�ˊ0�;ⷺ�I��K:�,���h�ݬ7Q�yY.u,
�De�Q9ڡ�(iU��
��'w�_��Ot���l�Ԓ��QR�j��Nϲ�P�٨�tK��,��'�O��4�1�@�@���Q�7$U�IH��o^*D!����5�����N�?�|��2�#cզUz��
�*��T�}tv����	�h����u]gFZ����nN�a����9>~�@�3��M��.-�ܰ�z���Ƴ�l��|��ۍ�p�d>��������A�Ӭ��;Q�dk���8^��k��4��W�:X>�!�}��vM�c+v�֡z�ޫ�>�v���nT+oH�Օ�w�X�кF��n�`�3��ŔŴgAd��8?�^�.#�|���t�gi��U�Uzc�6���u_��0�^�L�ݶ�5��Ȍg���>����qZ��1��ݒ	�E������͆3�7X��Ok�pɃ(�f<��:7F����������Ӽ�f2Q�N5[�L�S�����x��p���yY+��}����cg)<y�m@�N��.T؎u�o�}sޕ����</.���IFood6�㳏��_'��:;��֢}�PwLS�`ocaT�S�vB��\yf7����@r���H7��G�xxy��{c||܆i��s~l �H啀�~���^(�R��D0o�u���N��,���6��=�M���Bsd�"F�Mu����XC�����体���U��۷��ޣl{y.�v��\��:���̄�E婹�26Y
-X^d�P���N��{��k����Ud�z@mAe���Lmrں�sNə�N䞇u��Hm��h��m��c��"{Kr
A�F���P�����������h�̩�����?�+��O�(�Eo�I�L������ǝ�ݯp�nG&���]:�ph��pS��r&�$iC��W9���ܟݯ�P�>Y�#��C���A�c���ʼ�A�o]�<I��-gc�s�����S��l����{<���Ϻyk1E�e����������њ��+��\��F���k����l�X���'��5C�z&����y�˼�U\|�=4=gH�
��Y������C��XҼcM��eL�u��j�Wa�f��G�+W���Q�����Y�7MZ��]�Ic{ک��iueX� |�Yg�fB�Mm���NDMN���Ⱥ���7���GK�J!�?���:�='_g�w%���Tūi��c9��qU7� ����>Z5� �1��ׯ�X��[�]*�g���7���d�ɓ	[�%�;����c�6�l9���a�ͤ���z.�d�I���7�y�b�W/o6�/�;E��z�@�g	ف:)*v\�ZF�.�9z�~|��q\R\���s�˞�e?;��^�+��X05�..�{xd����W��ޕ��)I��<�g�4;rV�.c�yq;�F4�7��f")bU�7���X7Q1ګ��J���\��u���:�֑�jp^�m�m��#�[Y�p,"�qAM�^���D-DI�y㦌RPܯ����P���έ#wg�4�T��
�u�x.Ղ�F��AOM��hs,��\3S=�wQ�3�z0�܍V�= U��.���½<}���|-b�kWYT��uNb;�1X-�)Q�R5J�u�<�9��@��:��bT�S��ѕ���V����J�Ƃ7kp�9�['J�Ywf���1�qP�I2��d���.�ڝ���N;7��Y��vޠ���Ŝ��2NGl���w�\OA��N�Z�æ�f��3x
�^3[�
�vw2�e@'��8�F��^�#+���f����Ӝ�һ"��*{	��L�g���_s��lZ0�4�Ө�4�Z�\�#;ge[��*
��vtf�r�n����v(����(���9�������	"�L�F���H��4�Y�<�i;0��L�2�|��s���C���U�y�;ח�:i��}�m.�[T�*ɫU��L
�����k8����"�T)�p흕s{D��>��-��L`�L��\���k��̹�7[�5��B6Gzl���ok�κ��-X�2��>u�zi�X���TyԴ�oC)8��He�"�j�j�������镔,�㮶�q��q7�]|Z�P��ޟ��(�3;g1�k���^����m^���:��/��-i�^>�CA��y�Ց�
�U����]\�}%��{�@�ޝE�Y�7@�f��Z'N�wŤKX%B�.�Q�uQ��	O�؅�#�F�0f>C���<7�����ڈXw�1�g���5;2�!*Ǣ�2a��&�p��Yٴ��&�-����#8���s�����M��ӾG��˫
�S%:2c��^?������t���s�g毘֭WE�{7Y�[.�*v�nsXK�
�z��ڴs��}�� �:҅'ԷJ��'.�%��bY���;�&j�lN�*{&�/��b�Ov;�����t�քK�	�c:��#�|�3+9Ώ$ɋk ٌ�e�<��;���|ַJ�eY���4�\���a�X�Ho3B�R��_YYK��A�N=7�A��iC��5��Ĝ:�Jsۡ�im��}��-/������}E��N����.W��ʬ��򬅅9�Zw6L�ެ�O{�o%u.e��9����iK��SsS���Gz	�ra�ڌ���V7��Go��@*������8��u�;NJ�ЙV0w1ff��\R>�L�C��e�gC`t%�z�rN���e�1:搗��� Mh|s���p:���L���2C�B\�1�v���enaU�*�wpwf^�f�Q��;:N.�D��7��{s�p�o�	�{w�g��!��;�Y]"ut����mWlS۾�0ȑ}���G��B�a���UN���p���I<�n��K�]�RSQ�Z�-;�F���+A���w�ë�
"Q%貊���K�7�g+u���kFl,�o,�ԓ��x�֋W;�sx�.ȵ7>�*T��Ǻ�@=\��z���h����j.���&������h�&j�֢�3L\�5���:s�����}��o����o����MN=����4A����?#5Q��r �����������>�O�����}��O���?_�~Zf$��TAM_��4�"�N�噪"�����O�f"�5����*"��������(��88-��:�PMQQ0�%5w&��X�u�& �"����?'UEz�**������
�����9�ͨ��"(��Q�j��Zu����DS3-SLETUT7�U]�z�Ԛ�j����C��c��MAE�6�UUAE]�E4DLRDDE��-��	�咨��1E�$lh&��0�����	��1M�*�)�mSQ]C����
(��ADӳ���M\ٛ���LM�����<؊����l�)Oy4�UATUUDDA4SUu��-U30TO���u�qT}��U�w;h���kMlf��]�9w���=v�"6��u��r�vL{��gk�=D>�6�2�����:y�����������%¤Ug��SP:�7������H�ʋ��X���k\r�$q6(�+���vu+�r�.5���l������2��ƺ��}�\4&�m�
o�Mv7vS��.V�{��]eE���v&T_�o��=����Q~c]�����f��7����(���-����-9z�O�gˡ�c��(g{����﫡I&;*��)=��������w#H9���F����8�7�̀���^����5����5~����)|6-�#��p�uP3�P�����7�3�t�j%��h����L�gv:c�p��E_��k��J�ŷ��4�I�3�Ǉw�G	kx燖Td\&v��Ѿ+�ɷ�����n-`Ϸ����h��Fz��L��c�5X��qV��`*�1*$<�5��y};���<���r�������" �ْ�݃���;L��׶Tڱ�� �-H�H��]d��gí��޺_n��� ��Z�M��	T�9�_z-�
��r��8��j�mJ�8뻖�������;x���d��������a���I�1�/��]���o0��xq��=<�-�@!�tBa�Ѩ���̀��H����ڙm�r��>��͙7z�zu[��g�	ڪ:����O�S<���k4wY��q����9,�4�i=qQ.g:
�Lng1�;�T<�Sy�F��;�<�(Ϲ�Y^E6dЃʀ���:i�����$����8���.6DFܘ�Y����mI"ΗT�<j��jw-ӻ,<�p�ݽ�z��.ȋ��@�#ս�l��GRE_����$M(���g:j۵��@�aq%�ס�q�4p�WL���*��e�5�U�](�d�7�\�dOl���R�u�|vzXc��VX�t���z��U6L]cE���d���b+�9<l��w��gp�����@M .n�����K���6[㪭FL.�8Zt���\Gi�������q���rΐe��0����t�es,�I�k��Z�z)�vuy��i��%�e��s�ˍ#��t΢��R��F�Zy^�J��P���X9��W0��L���t�k���c��*\�g��U/�ɳ���^�^ʁ;Y�;tqF�5��<�y�M�.� P�#;5��)v.��Mlve5�&�fb'�������~黿D��s.��LPQ���/Q7:uN7���+�@��m�``b��/�s�^Z�"��3y�03sh��rD��o.����6m�����M�q�[[},sp5�,����P���*.�����&x�Zk�S��5�ﳽ�}bF�U��t3��h�xTj*������DB���͓u����m�j��}T;����C���!�3(eC�R#j��4F��%�Nղ�\7�����"v�4�"��ɦ�Ԏ�x�L�PI��n*1���Y�zrk�c�*�F�)m��|ڐ�cO�-"���j9�O���ڪp�#�=��O�n#Y1���$�֍���G$�[��"�[E���ND����/+g�q�rv=�� �ˡ��$"�+��zt~��+�n��B/�g=�ݔ�&��+��ǔ��\�[�w�%Q@��C���5��l���:��#�+_w=WC#���/�Ҭ���Sȱݚ�o]M��ߔ�w��ݚ��ma{�=B���7��q�ښ�wl��K/'e=w�;	��=�]t7�%s��1�1���^j{
�b�E���}�/�y��T0�-�f6�g23�J���k�R5���[Eu	!E^9,�&�6m��mQ�j5�G;�62��|�g�;g��C��T�;p[�O�7|e��*b�N�5u٣�ʜ�5d�QZ�4��e!q~��z���l0���D�M�&3Jk����t���3�UqE�y^tH�&�I�����lz(�gN(�m'�9G�S��N��Y��h�\Q����*X��L�h{������ا���Q�^`��8�q�H�����~[�/k�\)�D��{�c_$�E'�fǻhG�Cl���>"Ѷb��-��5;R�^ǭ��3ٽ2�9�����/��j+�������_�q�~#�$6e�F/��Ws(�葼���N7v
3�O o|��(W�����'{��8�:7Yi�諝�ʺ葚OW��'������C����_V���+�-2�t*�ovO+��$wt)6U��|�N��8*�ʻ��{r[�b��{��*e^���X���1Z�L*,��u��-��!15�/m�c$�����4M�����.g	�ԡZ�)o�^���uك F�䇷bL�b�����ݵ��;~v�3'/c�gTM�U�.H`hi=�O�fQE�8w�fUJ��{�n:e���qA\a��E��1����(&���?\�x$SD��dl�K����}��X���&z��Ś|�&wm�6��5��^7p��ۜ-f�j))�F��V�j�� �Njab�;�6g��w8F�x�5��8nw_��7A��*��7M��u#K��^#a�BSQR�����C��al��6�$��θƾz����(6c��3�L��L#m���H��2	X�6+`֦���9����ml �T����U�gz�4�t_[^n��tRT� 0��w}0�L�-[��|�k���~�cmw���^�����Fc���n8f�!���"=��S�W��侻�κ�$`�� ��g�?'"���w&���3�3�C�y���bۗJܶ���7r�Gƕ_��1���E�*4*�u�ƹ��)Q?0�т�=LP�,�f�\����[]��ǻz�5-����`Y2��1vH����(�ݲ���\cQ,��k��nH��?���>���o���X��aΈ��0��Ay�L���_��<=�����b�V�Ϻ��c�(r�t䌽����������{skp���7��5��'�C
�ao�c����\�+#���mܭ/��0,|0��J�0ݏeƕ&��RE�h����x��wӷ^Y����c���.^y���=�f5"�ꮝ��rt���E�7n�)^PQo���3��.�Fd5uC1�:���`��u���u���n��>�����뉂j�礯��/�6j������s��(wٲ��ñ���{	��jM%�'�"�K9�agA\b=!�2��T>�,��7�N�U��y�YH� ٓB*�v~̮�SF!ȹ��r�S��wpǋuƱ�F��m)+�*�F���-mm7Y��S��O��ﵮ͝�|>8�ޛ�pd���H5h"w��-�m�Z�]��o�/��+��C�F[Yռ�1��};B����|�>�+���M�ޓf����Cהx⹻@�[c��=*��H�Lu�g"�wy �l�r䮳�r���Sv�e�.��x7��eq$�ŉMt���C�����z���K�'`&h-�g�����o�xxz��9u��#�U�ϫs�i�>F��E!vڱa�]��ײ�N�.a��K���i�W��]=��j���q�4ܧ�&�3�����>���a����-b\�<�_5֘��f�t�l ����G�}F��Wq�u��_v�F�Cïz�*,xh]�ʱ���vyE�H��#��ǕZ�1R�e^�Kl��׸�e
ɖnS��oh1�3�����s�PrnF�YD�qr�t���$U����Z��3׿pe�p��A@@}���+E�lMdͨ���f�װ�gM��nZ�Cl7@�fA3�F2����\X����ڤ�#:�k?m]W.����y>����U��dh��xRn*ѭѭ��g���sU���Ӵ�y�j��"+�h��\��|����B��DZN��c��F�gs\�FT�����@f�#��l���Q��S�OC��77�{p�8�.�ܫ��i��k2z�M�1�{�_�,ї��S@,2{4˖޿V�}&�(#w�2��%n紧�VmG����yB��z._N�J	���4J�i�\���ڐU�����re^�o*:�ثox��W0��{�������&�^���D���;�i�	
��	v4��S�r����a�6+=5y����-����z�Ks<����P<��hʥ&�AV���d�E_v�s�u�����_��VSp=�r��g�c�nAO�B$]\�U�]��k���+Q���쪱��<&��u�Dd�Q\�ㆱ�c�X+�O��ٻ�ۥ�;���\��D_Hk�R�pi�[���W�]�*@�ŝ��f�h�'��V�ޤW47d��i�|���2�3��3TAO�e�f�i/s�b��Vfɓe6�Z󦎫 ./Ҍ���g���S�ƃZ-q�R`��4�}�����J�����S�v*Yԋ��6��hos����CP������Ҩ�S��h��
&�߇d�[1��;ݑY���@�,i>�Ϸ� �9����"GO_�mǅn�*�?O���q������kV0�)81i9;;L���/,k����2�V])n�o [͍�*9i�;��:�窛�&���Cr�;íΣ�m�M�l�� �S6U�킶{o9�@L�C�<�#H��#]���
�+|��;R���|>��o�t��"������ ���Yͣ�|B0�fDu����ٌ����ȂYi��˹_��N����F�h���
�Pc�>���=����m���wgns�5�3��7�}���$qHH��N���Fv)�FCs<�����}y:�����E\��W�rX����~���y��Β��I51��JTP�lT��b@������!�c�ct��3eC�̴>ƫ�0���e���s t��W0��R��n_(.!ho&/?C&��R�.�_�T����\��q�z=�]y��š��s�c���Y5"�0X��[�/�e��k�p�'��T#2r�U:ʷ�]9�B�a���Nd���C
D�Z;P�H�sĩ�$,.�t���>=]XN˛������!�����h�d��.8ѫ�$g��� *�h�uT��7c*�-{Ujۮ��)Lϻ�_"����}�I��ð2R��C��j��e�ݪw"nV6[uhz��N���tJ������0.�SeY��E��� o��*|7�1� �3@}�qd�1:��A����:�!������w����0�nn8l
�5���dʧ�r��c*��C��]���b�6�?�Sɺ[�Ñ� 7���zu}���V��׎�ȭ,VEW���9���}!�(�(�p͂@u�@��"4��-�3�I�^�x����<޾="��)Le{m�{�cn�
4�ja�p]��[�[�}E�Q��:��2c#�匑��o��'�0 MeK6��6Rm�*�r����!�*�,��rE�]LvUqn�&8�����U������(�˫��wN��:�����dzS��>WT���� ��ki����Av���^l��αj���A
0_Xx*C�#Y����H�����i�+�n'�L��T�b��跿р�!Mov����fw�����r�CD���}g�\0�q5&}�ܽ� �U;�O��w��{������DDA��c�Ċ ���E�?�� ��T �{=n�\��'x�C*�(ʰ�2�2�2�2��@��2!��C�2��C
�"0��C*�"°ʄ2�2�C0C �2�0� C �0�*�*��0� C�0��@Ȅ0 C"2!�C ���A��ĎFFE��A�E�A�A�A���A��a�a�a�a�a�a�a�a�a�`da`Xdd`aXd�\�=� 0�=d@0 2�0�2�2 2�2 Y�������(��p C C
 C  C
�L2 02 0 0�2�PPi� !�@&�bed	�U �ds�ɦU �P@�ea`Df&Q&&f�A�&Q!�]�$� �L��L �0�10�LL�M2�12�12��py4��"�0!�C�0�4���Bi�a �!�n�C�C���G�A���~��*�@"�
 ̟���~����~��$��������'�H�����$h�?�������?�_�������UE�������C�E^�eETV ?�����P|?C'��?�?�_��o쇱ETW���A���� 7�z�������΄������b�� 
�� �)�RQ *  R ��@� A A( C BB ,  B �
 J�"
$ @�(@	", B�	(�! B!
�(�C
�BH�J��JB B� D4�p�A������ZPE(
��Q����_����������?����?������?���y����a��������:�������>'G�UETW�Bڟ����Or��+��Q_�C�!��?UQ@W~��#�_�'�����������/��C�~�}�������ù�_ga��ڢ�+?���?oਪ��@{J�������O�:��?p��'���{����������TUEp����!�R~_�����#�
~����@�t ����v�������=�?�2��@~������ϫ����K��0~���E_�s���������O��PVI��x�����` ����������}QR����JR�����U�E+MIQJ�T������
�UPU$�JITTPve	#m@�TIUփ�-�-�cZ-�EJ�kEUU�@L�R�Ym��1+f��YQݻi�j�U�v��$�kR��S ��Y*���iCDJ�Ye��fճ6Ƕv+a��wiH�EDk6�����b�+X�v�P�mm�14�Zmf�ɵj�J����6kjkVQ:��k���JH�������̵[*�%�5�h��,�[U�x 	�9b��u.���Ŵ���ƪ�˻en�[uƹ��vպ�B�����ٕ��]���:U�cN��l�g;��n�̮���h7u�ut馷4�v�m�3kk����66�CZ�5���'�� L>�
CC���
�x
(P���Cs���(Pz С�o}���:n���uu۰�iT�rv�]ے��]ݦwN�]ٺ��u����6��u;wm��Lw6�㝶[��}�����N�.�wkZ��� a�om+��Ժ��L�.�ÝvMYWp�Q�ws��k�����km��ҧk�,�6��ū�L�۷l���+'w]�m:U[���v���[b��g5ݕ�u��[e��ڭ��l�F�6� w_uʺc��WK�[��v��uGiݦڸ�ٮeMX��ۮ.�4p��wl�jS:�]�����9�խj]j���k�1���pv�`�r�6��O�����6���b�k� ꝷ�+��[:�\i���M���kw�s��նn�E���1]*�;Z�ݝV1�+�Wv�j�w[-��tB�mժ�l�bڲ�D��e�k�  �����ۍ]'j������wlv��}wY�ڻWk�^Ǎwu����^����M˙���Gu����5��Cf���˻�u'-w{��a��֡X�-�k��@�  ��F��h�(t\mv��k���ΧmVq�uER���  wwXB���  k5ڸ :��n���-�n�l���3MS1lkm_  �� �[qp P�=�Ѡ�;�  �  w[p j�p N�M� (.]nWM �� (3�2V[���b�l��l6�U��  �|  z� � �v[� �ڝ� ��[�  ��  qw   �㊧@��\  �w �wz�v�Y���4JUQ;i�� ���( ����;� 
r��� sW �;qp t.u� u9�  �շ  �4�� +�O�L�R� �)�IIR�h 4dS��PU@4  ���R�   S�he)J�  )	0���  bz=���y{<��Fg��z��+s|Ȯ~khb������P�7��Q� ���O�!���"����)������"��@�AU�;�3z׿���^��*�1��Ĭ
Pkp
�Gnܨ�]1���kof�Gdi+d��ʤ��wy�j�P�fÔ��!)ҭ�
`�)���і^]��+M��-�m�t��bu�=���U�ʗ.�i��ܐ�ژ� �n�Kp�6»�+i�߶�Q�#��8�˼�3em�1�q!:͢��4e��m�����p(�1;ҥ�B��rM��P���kPY%a�xMj�e��k�y����SM�Cj�(����Ԋ�K���TQoa ���P閴���@����ӏG0Qn�N�z��ڻ�����y�525��;yZ�d7�3q�0�Q��R��O�x��P�E)2]֋ Շ��,+V���*1��:�iz.f����V�[E���إ����m�-ػ�MsM���
�E���F�;z�3NpX׀�lmfk��+I����f+� �4a �����9�6@3*V�ӡ��h�D�J�yPӂ�v8�����W5Mi�+2���F�Z�Pb�`n�sg�\�6�n
9n+)��0X!BwkB�Q��c+*]
+�i��-t�S�,��[woB�V���L��,m��dH|:���E��Rhض���)�Dyb�	��0BN��"��D�%�7P���[�e(��sA�R�1U�I`l�ǢI�}x`���q3��h��4�� ��&*�Ӗv��th��r�Y�U�c2�1T�$�b2� Ey6�pU��۽���=��hڡnm*�Y���2�e�鱍RaN,n�7]���Wv�	V^��i��eA���#�­m��ǯiP���;71h����/-�ȳ�-�Z/0�#L��h�nV�uh�n齧vn2��̍�YWW��Ӏ�X�ņk��6�(�1U��텆d��(�oh{gkQB�[E��Z|�t4�.�A�.��0Q��VGA�b��LO�GSn�S�Vl�kE�*ݠe;S-mf���5)+
����TҞZ��m�B[ %J�a᥂�8J���I7b�7Y��b�j�B$"�*�aȁLV8��ڧ�Ɇ%k�y��o�mG��v2�ݖ��,j2�XF�1z�Ō/��(S��
���5���uj�'�j�5{�+��,�!�v��P��%M:/T�(�0�hd3u][ٵ�G��Z!:M%��w�)��6妡7-��UK�q"&�����ú؝�
�4�N\��b��O���+s]n�&i8)el[���YKQ%�r\Ki�rb��p]��q<wfLɗcv�թ���rd�3cnb�M�AU��)V�yv�Pe��f���Vi�$�V�:����KL5�-�Gp!��d��u���󥶄���Q7QkihEJ���6i�e�J���u�$���8�u�&ԁ�c�"M��l?�<�w�fY�ʽt�F�.G%�a�1e��6#�Ҙ�t�nc����`��J��{�1=�.���.7�=mi�iU���ނ�x��3M&��ç1���Yc^7��s��`J��&��WZ��օ+
�3B@�A%���3T�ĴP*�c�@L�x	�o"�
N��	��oᖥ�6���"��J<�����a�d
���Lv�����kJ��<
�* \�6K�E�dq摲[����1�v�М�,���9.���N�L˂�Ϥ�!ZY�mM�Y A �;�&����sc	h������!0w&���+�H��T�;�J%Wr���cR��4֒u�Ҩɱ��Q^0*a)��XVs�v�P���ˊ�oc�
C7�p�
��˴Cm$0� �����RXJj�8����!i�p�tG�W-M�ҡ*9�IHƉ��+6���A�r�E˥+t��g�¾Or�*��=�P*=��������kD[t��.����X%)meb҅�f�U��R#ᚲ��e��XYX�6uǺ�-�3LK!o�CiK�ݪI�}�n�t6�;4SC*cǩ��S�V@���X����FL��]YU�%[f]Ean��i�Md�[NU��LY&��@v7T{�v�+>u�SV��Ij�6�]�����p�n]��HX�R�����xo.[�%d_6[�V��ܽ��S�f)u�lC<N]ʫDh��qf��6���JV%�^B-MH�[wi%����l�lL�"���;SN^������&4�I������R���^"���`�JĶ����� �j�(���!���:$P�[�agn�X0�tU��˖��w��_[6q�SYb�RZ�������(<�7`��7)���ڔle6i� S�37$��m�BR�U��Ѕ�����KS�7�����*��n��S�#T@�"`v*��]:�ߕ8e�#4��*H悱07`rd�uo@�@�ի7i���i��h٤2�)[:�%�a=:�a�մ�PЖi�w��Zz�6��6�ۥd1����N�L�#.�@ �#���C9N��n^<�p�*+Տ�&v�&-56'q��z�4r�q�� �u�xT�|8!�f��5c�B�^�ҙK7IXU1U<������P"E��[J�]^[���&����wVB���W��ʚi�)�/1�H�i5�V8&5r��=P޽E��]����n�����Ӓ�y�M#�eU��HRF��V,L	�I��qnR�޺T��c��Az1 f�Owi��12�s&[La�Sf.�#V��z��XؖbF�e2\u*Ƃ�VP�b��-��cV�J�f�2D��H\q\,��v�дD���D;)1��W�	����[��Ȗ�Q˻�6�aZRhN
u����r� ��`2eJ�i�$���v�Ol,ӑ-�Rݒ��:&��n��p��3kb�z+J�����z��2v��h�o\��M"�AB��2�'P��F�k��[�x��q?��V4)��`mö���vB�}t�nb/2�MO-�D���Z*�[xPS��zU���-H���H|k1d�x�M��R�N-!hsS�fS/&0XCq���r7�r�O`�۬�b�P���f���f7_�<[n��gr�U�0��6��Yt2�-��[�.�;�l��3��ֈ2�����c ���1b�ÌU��V�3����-�Unb[ i2�́�Pݰ,�B��*�N T$�X3mIFAvTŘE+ʹ�ɦ��Us���%R�ơn̎-���C^�4Ƹ\4���5x��6�(:Ѵ0CH՗�m�H���7yO("m�ݪ�8����%�(��/l��p;��r�%��n�A����u��[V��Cn���/��u#q�5�C�,�z%<��������Y�5����v�淲���e�M<�����ux����Q�1̌��4EѼ����6�vO(Ʈ�@��%�X��s2dT#O^�ӣ[��+����-��r��5\حP�E#��im-�i�)�ь7�]�>mV�E��в�7�#g�F�f�!���
�ችd�B����g��)f=�]GҀ� 1��o�c�[��CM��R�ۊ�5��KR:[D#���ر��)F�Һ���o,h�p,vR��ݗ�n���z�^d�Nзv���C��?	zs.�ݔ��-��(n%V��1j/f��B�7&e����¡q��4ӽφ��<:����F��%r\�h��H�j�^-���NԂ�!����b�j�]wn�^YU����576��r2�=6s���t��P�Kif��!�#��ᛦ���c	X��&�ےd���)mh�+i�2����Ȥ�x]�1����̩or�"�I�
ب��B���1�rh��I��@�k
`����Z�0Q�NmL{�n5�S�G^LA7D�n7JR��kb����Z���rsi	N逬I��L�/n٣�Hl�8u����Q�x�U�
[�����nMޥN�{ABh[om)1�L�$M�ՄQkc�4Z��m�E!M�M��EF���r9��KnLŵ�m�a�"���w E�{�PP!���eঝ��/f�Ǡ�j�+aPu�UbOq�Fc�b���$FH�Y(Ԭ�cK+^'yf����Z�;j�k!X����t��2�֤d���h�VnWk+���"����0����!Ǯx�si���L;��/��R�P�f��Y�[�n���ATw ���sX���ۼNŬ�CrT��n��h�����hHG��Z	PϢ�A�md,��F�� XGh�2�M�xh;�-�p
����aƌ�.6)ձ�G�V�IX�up�0҉�nJ���p���E���wP��7[3E�.��Sw��QO�kB�YXo��(Fe�ak�Iԡs�����Ln��7t��H7���ۢj�y*0��Z��n�m��Df��u�m�F�ʸY/]=x�`=�$��5vPGe��x.����:��ʆ�t����������3 �]*�]�ҳ �6�<�e)�ɘ��橀8u:SvnB��7J���ț���ج�0�m�h�^��KOu�4�J�9<Y&,x-L�qP.��)鹁 [[�^�Q=6�'����r�&#J��-R�\9A�Ujo.dr��0���ݘm����5,с�]
ڇ� �4۶)�M=XيSIz0Y��Z�Ocоkr���n�'I��X�@�R���LYB�J��S EF����O5��ҹ��h=�V[�M�y6�ò�ln=���l����.�eĊ&�r�H�k��nI�8 �h���z���'z5�D��.�+r����Xec�e 4i��6u�.�GUZ�y[Ii�Ja�ʁ�2���V'�ޓ Z3.� ���ĳ> !x^Pvӣmݣ�,���Z�3*�r�[I�)�<{���25��l�`�e;T�]Ϛ/1M L� 4�3S�
��lJW��f�sX��lFK�ff��Y�Z�r��ia�u�|b����kU��6��*Á��Ɩ�k Ũ�.Ѐ=i�h��2�e�n�e&���6�ш5����U����m�I��_3Z�Ƅ9O`��le�BI2�f�hiha UQK9�ǲ��1�_��3^@H)�92�؍�%�u�� }j�(��7��66�M4d2�V�r�yܔ;�4�Y����ƈn�����u@<t�cݦ�:
[gqKLi��f�`�p��˘��5���WCXsY���][Z����5�ܖ�F��WF��R��9�%X�N�����SN�6��Z��MlsM�&M �dR�JU�kV��5l4ri�h5�/v�Yk�(�$Щ����n��Y�-\�B�ux�ڽ��a��;Ŧ�m�&
ĭ�b���n�r1"t�RdВ�,D���9y���w�Bh�oK�%nU�g	1+;�Ϯ�̕��5���L�Vl���ڢ�k[�5u��\�8)��"@�YI#J��K�i�-�7*˲4���AE�5o.��q�T諭��Bqa�6j�l�uS�7M�[XF�q$�Py4ݎ��@,\4��4cНҸ�h�ֱ�T4��0,���P�5��&�-5pYl��	�6�����hM[u#,��`:�� ��u1]��j�w��=t�̚�8Ln�okm,��ʀ�i��؁��n�bm�`QF���aUZ�]�cC���"+��L�7G�ݡ��gf"]쨴�H�I�Ȝ�B�1�x�
j�d6�ڦ�������(�aʒ��X�٠)��,?@���{w�)F����V��K��D]f���%sk(dQ���k����\
�mZ�bC�-=vCj���cR*�B�;�Y�Yh�h�`&NV�%6����n\��,�&[���ak��L���k�d��0���V�Nތ�ۍǫѨ�yi��q�n�s%��6f���\x�)�L��mmJD=2�(+!X����^&�&��K1j��2m��W{Ae�,����LJx�$pQ�r�����`ۗN,���[6�*j�/Z���Ȉw����2�� ȸ\���W��2�z�-ʱx�^CG�J�4�v+:�5�Y��Zu�@l�He�̔
�J���kF6ٯDH�)\�Nּ��C��7�����vS-��[Ȁ-T�xuø&���Ґ�n�]�,֤�le�1>��%��w2�'���0���8�6;*^+�Rf�cu�j���v(nW-X��w�3JAJLh�5ï�Q$��$/m�b������F	{P�3YG�Y��˙���,Zɫ��M�4%z�l4�۩DR�^��5�t�߄��`�P�R��WL�����k(P]�%��	� ��5c�@2Hm�	ޥVo ���X��6:j��E�P��3��yb� m��ʚf�Q��M:�;0U�z����Xs(FT[۫�@Vۙ��H�e���LV�ֻ*�i`kq<�T������KH�3W�n��n*�����;d	�"l�1�ЃUr"�^]���dh�0S�c)!�6�lU��
٪�#w	N�������ZS��؛KoR�͖R�KU�f4��nV���'���ӊ��C3�5u��I\����O�W�8	6�!����C,T�.9)�j�����ݕz0G.V��1�TF֝8*�v �qKԑ�ڻ�,�V�O)*gL�L�F���oA� �1PA�M�㴞�b��j�2�^2�L-C)��{hV|�[���bX�M�F|N���"ʓ\Nn-ىK�ɱ�����jŒآ���WX�-+s�Qeмl���������n�J'Y9"$f����^���/e�/"{��O�qKA荸`@mh�)R�EZ�$9�x����RmYn�wpKO)��9n����w��`Ո�
w�̍�h�g"�*����[ӭ�9Jy=�{/��&Pu�,���Is�G���חw�%Zu�c�K��{�}�B��]#�x�N��3�N㬬B0�! �6�q\�3Jȩ���Ӣó������h��q�Mk�	N�*�ĳt���]i�5�9�yd���.��k��:!�G[��p��O�v�K�i��ZU��ᰟa�N�hv����C7�Q����SZ�p�W��ꏺ�ݍ�=����U��h��e�W�������,C������WR�)7�9�����b�e	���J�4�|��N$�M�|�u,G��X4s�dfFv3Q��J���]��������Y�@�敭��[��c*
��;�]2�M2Xz�K�\�)�z�՜�:ѝ��s�&�ct���f�EHoqllu>�Cn�Yv*]�o�n�ޅ�k�ǳ���<��PWi��e] �+�n޾�:�n��K��eo�!��,���陔��\Ua�KE�i|���}R�"�{X6f�寷�#��P&
��2���d�6��W��n6�sıf� �9	=+FcjR�V�ԙ��p�N��CZ�ܺ�%$����I\�����*ȼ�|�u]�M�YN��܅�꾺�m�$1T���mm+��6&ސ�o�����
@89�v�z�tJ���(P�j��Y���� ����ޛSe�X^Pݾ�4K@�s\��s�:�9,��<	F��nھ�A�]�j�V�pa�N2��3���TrIvlfg|Y�Qj��#j�.U�!��wwf�fN��2�Sd@��h*��T�ܪ�p�c�	��}3�]<��w�l"1C&�]�Ю�h��ܥ���W��;�ޫW0:���O�js��D̰�a�Ή`��طEJ&���|�,䴬я\����_>��mk�q��K��]����]�E-�>��'��M��x�b�1��]��7X��Ju`줦�|`�)�׳wT���!|���5 ��,���QEn������7�,��:g�/7�2�:y���rw��']��瘕l��N�ɹT��֞�e�j�Z��A)j`!�:C�I��I�t�q�K�k�����^��A��nW.}���1W�Y(Z"�2��qQՋ�l�WD��XqN�7��U���/�x�8Ak�Y����Һ��	^�w�Lz-	��u!5qT��r��)r��"OC�B�8�7�`J�sXx����e�>�U�#�Er{�՜+�q���ΰ-�������t%�����w�&�:I��-Kpm�A�c�7���ؒ�Ǹ��8D(c���7��퍣cl]�\�a^��u`Ն)�Z[�\��R��1�wl��rt���I��vmt�+d�7��P�ͫ��üzj�!�*AS���jq�F��i��]���hG�|�� ��$w{]�+�+_��>�y�r�wl��Gc'\� #�w����1�]VU;��=S%Sp�%��h��D_)f�j����0�.��0]�E+k�Y��K ȧVU���u¬7��`[	�Fc�m+�����I�O��ۗt�u=J��Ǹ-
RY���q1�m��ѻm��z�2�He
}2Q;c��I[Ieb=�>:�����,+mǤ�-��uP
T��{���c�^�c&5OoP8n?�<E�����Y�V�4������a�i۠�ki;X���M3��kV�\�D
������������͏]�Vz\sU���鉌ok%�m[�����J�A����<J�񵻥⫃�_n�Ҧ����$qW��]���1�[��h����>�%'[�qfLc�4�Ch#o탥�֣�䣘��U9u����\[ύ�xHMڗ�d@�B��n�s��b��I��S{WA�1�lunu
��p\����2�1��c.cb�S$ǣ�OXū.!4�Z:�Sh�����WѴ���R�]�ﳷ�]D&v�?v��L
?����+t7[���X/�K��v�w��X��V�]�9eh�E�����/��\�f�QiY�v�Rً��/�O8r23�Gi�dZ����3J��t0-�Hb���ya\��v�ؾ�iK��|�>�6��ü:�[�����:�tU�p�BѰ��4e�<�y�rQ�}{#q�Ŝ�M$�DIM�ڱ
��3@��Ψ�f��c][IR����ͽ����
7Gp��A�팩z��>�"h`�ۃGr���"b2 �II��k�	P2Mk�uYy�1]rŃ�P����I�{M$�WQ���b���;�$���I�t	)�P�.��3�8����0�=����X�:��07L�J�9����5�n�T�$�V�ɣ��ql;����2I��6�ZT�)�ל� �w��;��-f�ܛحe��qweL��������S-�٫-	ȚK0v�l��!Y�r�z����h�Q��h�7���F��5��S(P��s�F�]�*�
�S�ZsW�CvMվM8�p'v�]�k&v<J:�(mWi�P��\/�FU��\^�:n��df���֑�R�xGr͸�7�Ni�X5��rb�.}�r���ŷ�̧ٙ�&��+k���6��\�7-�@��`�׷f�2���XX]D�,s�f��Tl�f�cHU����ފ�EX��C��W�GWs�;{Z�a*�N��/7F�u�V���5�jl޹���)�[��Zf�s���ZM��?�фUҥ�;2��تB��E=��=�AW�����\��vj�K�R^l��X�ĚF�tm9.�[��2����%������2�U�h���X����4�q��i)S��%�˶�X�)M��#�7h���`�Վ(t:w�x�ٗO��7�*��;��(��˵�����id��^�?j��[)wRPm�w9���*��sE{u
��N�
 �*��3+m0��]���"����3S�pn�͐6�%s��|\]�NPHw7����nʉC��H��+:`Y7A�HN�8Bu&��xST��k]Z p�W.�\������0��mY
�=r̊���1Uf�ʮans�v�<���J��U��{��m�Q��Xi���ue!:Z�9c��c���U�NEۉv�m�#7v�����M�:xBu��kr�F*��.�]Au���3�|��й@�?�\�8x']VU��/��5��aZ�v�u4]���&���|�bs�xqD:����)����R�TLU;tp"��q�3r�R\���HI��wKC��nC]�޴6��f�O"�s��(B�8���`�QF�tꛒ��xˎq�.�T���kE4�m-�լV{G�>WA�Ü�t�!��O���u(�]�h2Щ���sy���wB �"���s����������=wwop�6�p��t0=799�U3�+�(����&lZ1D�Y(�9u��#6B��(æ3C�٦;���:epօC��e��ִýX�iseI�^k��¼�sK������5�AՒk����Mڝo�����Hy���wF�\˭�d���V��1��x!�8��pҺ{���c:jIV��B��7���.�&�B��r���f>ous�k�]9�v��4~��UA��C+�[�>��A���74Ԇ2�A�G���u�ӹ�����,�Ϡ2�ۛ��[q��f[̏ {VQR�mWof��.vh]��Rm�TY1��f�D�XR<��z�[gz*
��t�`�6]�����z��/4�Yo{�^(\4Z
��3��7i��v뵨難C��Z��l]p�A��(������f���wb�$[�^)�x�	3�
�u��c3��KT�nAfu:}Sz�v�Ю�/jZY��R�����$x#u�zYL��W�kH�����x�l-��&[D��HǠ*9\'��oLMwu��KI>v��TN�o8l��y&���v�7�����3aP帺}�;PT6��;Y%]l*�5֫�ň�e���{�����cj]p�����D�5�)�F����L���:\J
��h�W�fgq�(�0,<oV
�w|����2�2���y\��w�My �Y#�ɼK
�l
X�}}ϡ����]Ѵ��C���v��!2�rڕa��!��@��Q�%�X�Ѣ�y{7˕�	��%<��ۙl>�u%w+(!չ���U��g�.;�O�/��]��ܮ�VY���LsI]`�e���_TPvr�@�ta�itI���f���������}0�le�r��B:�Eg:���gܘ
�o��峋|̼�����*���2�-n�{�y�OT���wK�[̲�����W&5�t#rZ'J�������IR��o����ҫzV���O\j�\,�L���/��vB�mʅЛ�����C+�6���{h�g��Pv3ef'�v�Ȟ���.<���fܩY\z�oG�^;���n����rIm��t��Y��ˠ �����ΰ�h�M��U�)[�
ݙ����,����o�G�vj��[H!i���xP�t�] <���|��{���ĵ^��%\n|-G�0Z$�.�Gm�C�h�yܾy�T�vo0DBQ��[�x�κ&;�)������ʋ�W�J��l�\bk�B�i�--�l�4J�z���YJ����t�˅�3!�4Q���z�S\�nt���՝X�',�ilT:wQ�;�ܗ˫*c�.jB=F_`P0�n��j0|9'����e���l��Ն���M��r�Ό&��f(��rf��k��;�d����ޓ_n��l��'۵ylV��_VU��K8����t�����6HK<�	�9�P�+Oz5]P��M��Q��]�G�q<p.�������ܡ]׎)��Ժ[\�:�X�Yc6"�
��y�k�2��6	�}���� v��1M��Ck3N����ph�2�9�+C �	�ۋ��
CpC/����O�ne�=%��0�O���9�����d�N\�R�^���\���+զ�팜��6�m�Dڶ�ҪVQ�0tc5�؛��ڶ����E���R���A���n�/7E�
���MOT������F��(�e^���)�X ��&4l%m�xN��ux{�����k�C�`d���"�F���5曒��RR�g����v���¯/@���un����9�	ݕ|�6c��H�Ί^Wf��Ru�pm�6��hY x�Ѩ;��FwI�Y���h�J�@]���2c�[���/�U-�Rt�j��	̮P���E.@�i�A�,�K���<�XFXbXE)U�t�oKM��v��-rލL��Z_k&�Z��쭾q��^���,�3wn�\0�t:��
.nZ�ee8��Mou�R-[x}����.������ܮ���LNg+�	�k\=�h�7+W�~(sGq<�ȫ$��9]h+�z�ݘ���HpY���2���΃f.�����5�RQ�/��妐���xZ����y�/���0�� ;/+��N�i>����S`�i�96Z��JT{��K��d�|���A�|�#+1@���Ew�e�*}0����΢b�0i���J��/��i s/$R�l��`�.`〩����̴ǓӜ�1�y7_MǪݿ�w^*1�||w���צ�6������M���Lw!Ԑ�����X�Nj���ֽX����T@v�b�R.
�Ve�X����㏫A����F�v�,��/Ff��z��U�ܲl8i�{���]�XbqI�S��ś��MD����S�Z�e���<�:hT.����w�u'o��Uk�)N��`�x5Ju���AXud�Co��E�}�Ns���kg^G|r�hڅ��P����%٨Ŋ�Yb��X��8`\^
��Phz.Hwsc�ј�.���(��m�#�+���N�L���.��
����R��P�W�AP�ɓH��igfbR��;*u�ڏfw���5;)��Gܱ:v�Zr&�.��w:����ss^� Je�J�����x�"�g;�h���7N09*.��N؈ۿ�GE3�Z�p�JVoI�Վ�R�t�!2��h[��;G�p]��}�kf�<��P�2gT&����Id��d��=ʫ�4���Ni�����E,�4:�#���3e�p"v9h�ЛV�[T˺���U�#o+�_�j�^f�	�oz���c���MR��]�wr޸r�E�퉃�pW'�,��� ����9��^�*��GԤ�a���"-I�a�X��]CF,1�(��앦�����c�^���m���WC����ޒ���mN�g��7*�K��ˮ���#d��f��2RD��t ��=E%�IS���5!�!o���βgݪAy��.R�b��@vV�P��<�AfHE�=��0��V�N���3y3i>�������a�O<�B�N�꜆SqV���d1�؄���BL�!_u�7L��9�޼[X��6{�V�f�;)�疙�q��x����s(1�:�,5��;�����	��rl�g�f��I�m��8�������\��<�GK�r�Vh7��'czƻKW9��T�{,q���Z����v1�&tyy�oyr����B������u�&E�}7Y9$����W|�ZY9�S�|��酜� ��o�۹�jPr&���}F��ä���g��H�Q<���}���:�<eK*�󩑄1 ��'��BI�X����6���#�j�|;4���-�uK�.�����uZh=�3WgKw�����0�3z�ŃT����Y5jf�ڡ7�J-����I��׼,ɩ\���]�g?��&;pɲtr��M�U]�>�;�G��>��O�@T�P *=�>�]�y���VYx�?�?�*�v��r�� �����B��夤�x�7�����D(��Z�$�W�d��F� ����Y��h���Q:���l��s�tb���ゖ�h�U�g��7��Zqó}hnS5i��!j֘��+��M�Mͭ�Y�b5��ȍ���A�����_&)���M������z�9g�D����Z�A}{��A���U��}��I1k��mr�)���N���P�m	����!3���j�����`y[�+:>͎��1�#/��j�D|-lwx7�TpE}�
U�s]J�������KA�{crMk62�e]c�Ż*��<�a�R���K�߹!ԫ���׃8<�"*7]��ԝ���⸒�1�$���o�$����>9|��	�wamS�f�K�h��H��P��f8�sA[�]��36�k�.'EV&�";��T�<q9]t�M[s*���wZռ���ܛ�r�m�'Iz! L]VWg�Xʠ�e�^�V6�u�脰o1���\���M�ٹ�%�&�X�*�AB��%Ʋ���59�����y��&#�Tŋ� ؄$����y�5��w�5�����2������]Ν2�V�a,���}�A��I�k*`J�Pζ@�ѝE�38	�ܸ4��,	�6�6uG�_�]^Vs�-�R����ݚ"6/����,MҲ�Gz@3OK*��_�ѹʷd	r�a�{|�=.S���r�W�����Tz^�Z��s�DҐ�n��K��|�V�j參2#ӱ�6��
��9	�%�\���v挛px���tC�bl�E�I
��c4E��$�M��x���on3_ʘ���{ҷq����c�vWԻ��V�k(o*VB��x�B%3���s���]������V-�\�p�ʸ�gӪ�6�8m�υ�A�BU���U�:��kaӲE��[2��вk�6o��O���$��a�����u�b��"oq��2�
��M�jep�ڊ��F��xg=a�$�kn�
�8'8F��J\������>T#��groN,%C}`Ԅ轨P�kM�ˋX��6%���_!pnkY�W2e&{1�ܪ��\�Rjo[����2�h��t�+M��j�/�y�d��F�v%���7
�krF����t�nn�"��j	�<��Qi����ر���vxy�%����]�ҠP�̹M����ǡ^)�Xh�5J�t`u�ظ�vv9iP�����x�h�Xs^ҝ��9�9;hR;���ai��m
�]�����-2�]]�6�U����.Ѯ7Y�%�!����"��1�Jk)�z��y�<v���C�s�H�F��ĭm5�r����#�v��ߔ�(̫�R��)[tt�N�b$v6A���z�Ïr�Ğʰ3i�D�K�T -����9p��n8S��y��8���������rj������(���Ȣ�L����=%`g�&
(��c��d *f-6�n�q��ok�ѧ)*R�)+�43v��S��Jܓ��:�㓜�2^�Z"�C�݊�lǴ��`N�c���}�Qd�넩��P�j���j^��}}����ID�ǐߞ�R��5XF�6Z��fh��.�*Z�ܺ�vo��X�v�b΁^����]�{S�IT!���.��wALSO
����EA�GfY�+
ulg_2�F�A�5�b;�zQ��F�ʔ=PVڬ���=����T�6���0ST�)ymd�©�Br��J̦��^42�/:
K*�T4��$�ج��v%<��k)��7f#��j�^Ƅ��t�1�i�NM��.Cqen�r6z�����'��2n�I��/Lȥ��]:�x��p`Y;p$�^�vy�Q�}{q<5������O0Ŀ���oVV1x�-i�x,.Ɲ��֤؋r�i�W%1��}b�zҙ��l�{*�@���夰m��u�0��/�*ק��5-Yj>�ÒϖŨ���-��^q,���YWH�Y�.�V'<kz��gY�%-
���R��K��u���f^(@]u��h�LK�dL���v�ln�Գz��p˥���D�n<�����t�ӈ��
Dh��0L���ܲ+DpF~�����ہ#��JG:�1d�]wj��]n�d2��CD���]��*o��ݳ�����5�Nsq��
v��J^��ٝQ�Q��Zl�6�,!^�,�D.PZpu9k���R��b'2��@��[��z�ʱ�9(�Rr��������-���*ro�&�1�t�}�s���?�H$F��Cb&��9�o��G�9}.�1��5\y��<�vr�Ce�؝0�i�������f-W���U�4z�v�R��u7+�����v;9s�+WM�� �b6Q�6��/����oGR����'#�GhP��5uMEQ�I��?�7�]������T.L�gb5��:Ҹ-<��Px¼�p��Jt�ۑ����+fw�8��)e!��UV�|�ŭmbe���ow�A,w�X�ŷ��bk�X� v��d�:��eB��X���[��5�ʱ*�Ue_f��$� U,S�0V=�-p�X(p�x G��mqS��}��p̢�$z���-��>V�t�dl�WI1�f��j�:ޤZ�ڡk#^�N�����Z����w-u�h�r�L�Y��OS2��V:G.��["n�U�f���n�'j�=3�7��R��e�7��m���ue��LMѲ�E$��!�# �G�&-74���<�sCh��Y�0�Y�隑ǧs����o��I�kF�J�eme�&����{4�ӇZ�j����)�9��3�>�P@&UҠ�5�&D�tq��)ĸ���|��<PK��&��R����t��i�,��fL{}/����t٫}HP�\����f�5�m���f�,�6�-Y�]��t�1i&Y3��|��E������U����s���ֵ�v�wr�<'�%%+b�V���)������LV�>8.��m,��G����M3�"�0�I��s�<���{�to5mr�-��E�n������g>���Y�7y��B��k��s�G,p�"�)=2�v-����+�o9�*�ee��*%c]kY�̋j�j�dL���J��h�qJ'��2�O��0Z[��]�1�A��kk�Y�k��!u�H��CC`c7"�#	��h�z��"�wc�gKx��/y���G�]M�Ht��톷�-�$��@W}lȘx�l.ХuԚِ7�H+g��c{��&��h9���cF��d��`-h*ϥ���>�%����I>��L���N(�놸���\�o!�UE�>3)<�,�v��)\�R��+��݊=V ��{��+b�į��7onLa�ho3i���rFw� *�L1�v��i��`n�jG���< gj��knk,g��؏#{إ�	��E+@վ�m0�:#���\�`�ݥ�˔����(`앉 ��ro�Zo%�(Y�tK�2Ȃ��M��;��@�	ؠDݷ�ت4Goc&���y0���	�/��r}�Q�=�5\�+�x[&ebY�1�@��ū{��z�S2�R��m���ʵ�Qw|�4��ҙ9��O4�ݣ|�֥��	e��Y��\R1*�e]���Ą����>����+�I<���ycZU)+�8T��Y����6�})յZ)J��0�X���gT������;l��w��q��;/[ޱA�S�r:B&'�y��@T�pDpV�S��dy4���BM껾���9�n�M�V�2U�i+��)�)�n��UMyC�"�F.@�x��]T�z1��´���K뎻Ao����!a�ǲX�&xˠO]i���T�2�r[�)�j����D��捭��Z�a=��|/��E�җX�7R��r۽E�`t��}wW
"��X���LA.+�Y��'u�v/�g���(�ȴh�nmhX\Y:*�8�p�˭��3�b\Ŵ���.��.c[�n}:)FiUg'	Z�N�\��SI�a�-�������e�����&�R�M�:�z@�k��&,r�Z���T�Sl{r�!� ��F�C��U9��-Q�7�ĩ��f���Jˎs�q������*����7T/�R]]#2�lU:��oG`vi֘�>n�C�:�7f��ڰT��^�N�n�����/:ܧ��sR��5@M2�j��i��M��iм�Ꚙ�Γ�Ѡ�������92�ܽ��uݦ��s����;��Y�j)�u�}D42H�v���ƍ��Af�g���o^Յk&gsX��'a(8�V�zo�j�#ݥM�K���iZ&@���'��J�.[T"�����#�;G&��n2lN6c��Zo�v���SJ��c0,u�h�buy���3z�[�i ry�j�w�ʻ�,������щU���Sn�T9��}B�\9Ҏ]��3O>ï�a�{�K��p�N#&tݩm�B��{�lF.y*��]T�ze�Y�[�:�m��O�X�49@�9�J[���h��k���Nf=�Tm_[U�M�q�a�r��k�C�eg>(郹�X�)aL�ʌ>AHtd&S����B���%�}������`�t�''EE(��hޭH%.NG����gS6îTr��GE�TR�HY)f1���|n��8��
�R�{>���ݛ�BglJ��.f\`Ns�,��.�r��X1��l���-��i��i�_%�z�#uu�+�6���WV3����u�z�]�
��!A7CT��b�8��sN�5���O�v�&=�	�-=Ѩ7�KP�74�T�`�bRN�`N�|b���y|:)Z��f��[3�3���..y�E��.�:b�u�F�{�7m<��
<�!4I��mX�;�����я��U�M_N���\���L;�P�IF�ա�e��2��Mf
��l���+�ўJ��ˊ���ֺ���jr��X9K�TJ��L��р��@�!A����u�nC*R���<�0-��ɧ�`?:�^өj.�U�� nZywF���puo�Ke���uc��^?��̑L�)x^x�n���ʩ�,��k5಺�����2-�&�>%7r哥�!�am�A;���.�x��ai��y:�0>��xä��;�4{rfvܹ�t��X���5gsk���|��/Gl7wup��նU��Vـ�)����0Ke[p�'�ө��_S�.�����v$뾟<�J^s�*G_/�Y��5�x��ē�tNgE��e��]��㮁�7���/�<-��Lu��z`t{k�д{J��m\�e�f�f���i����H*�ط+��+,ݮ�O*WZ���ގǣ�9mi�Wn�e��v�p7Y{R��f�eFt��/�Ru]�Z��u��wk/x6B߳')�'s!�8�h�X��v��Jﷲ�5��[E�*b��r`AR���A�=�܎C�&��0��	�u���Y9�/��`+Ul� ���l�����6@��0�}y�����2��eU'z�e�v|���]ĺ�0���S�jQB�㶬]����QYS�+��7����+�<��z�Rɒ����)vK�9���sls�yBغfs�ـ>n��Єk�h� �
_;6�fq�D\z�*y:�Unvt��G��"��H`J�6*������َ8a��ʚ�r��`����޺Yʸ�n�d�Tra���$jn����Ӽw\�Bq�SwF�r�����CC\[Mܡ��A��7t�.R������M�X�v����k�Y����`џ.�Z�tgS�3�Y\�jm�֥�=��r��4f8֞w�{�B����f��:Рmo���<&�(�$��Oz�{VkQ�KDtw�. tAݸ���ޜ1�2�fwp��ف�Nrj�1Lq�b�b�2ꫣn��D���n�Tj �j������6��sp`�����ۺ$�g���[J�7u׫ �X�).��F�N������ ���:��Ef_\ֳ�wVv��-��S��鮺f�)૛K�*}kY�i���&��k��j<.�P�-	��D���w��v�Vv����N1�iɭ_���Z����8�,r��|�;��kN?N*��<�4�fs�}w\���l.t5�	Ɛ٫�$�Ht&Mk���Q����]K,Gg'�x#���b�B���b�ٽ��d\��ȹ���GV�������ݰ�ٮ�>|������Z8h�9-Im7��e��$q�ɍʕ��
;��3T�1����s]�6�!c�(��>F�yd����Q v��<�</usk�.����[��;1����;o��(q-8(1Z�4��� �ʮUkUok���E��f�#|hrƪ\�x�R�W&�f�m���vr�Y����q-֊���`��R��J�],�X���Z��
�2�Z�J�_4�*��V�e��{ŗ���\�Nv����&�.M�Ȅ�����l��fK��Stk��4�a���#��K>fk���֛��UP�y7IC/(�,J�ip畭_H�P��ӕ5��n�YP��!®L䷲l�y�©n����X���Y��s��f�JV�
�Ž��@��d�:w0�g�K�K�:�)�KZ)�V+�A��#ӷ�;�vﻡ��cP��OcR)γE��WZt2�=\��I�ҟnf`YT:��:[$QsݟO�z�r�tl� +�����w���y�yx�����fƷTD_�ðշLe���g㨮S��͟��
Wq$hd{�m��~C��C�̍�z�9�%)ûһXu��k�S w��>�5d��fW��������>�z�?v�՗��.́o0���$�z���zc����}��+ke�t�d&�Z�ƍZ
6J��V�M���3�ē#V5��nCr�i�H�ԁz޾��*�Ƹ�^\�t�V%Z�-J�]W��P��;��B7�Q9��,*�ZR�������X�-~�Jq,{}�COr�� ZV�wTwڳ�x�Nht�|١ح�2�mD�ވ�g\샐��|^oZ"ƨ�W`��A��wj��q�)y�i�)r����U$<ߗo
��;)� @<���T��@j��}1��´�����B�hݞ{D.س^�p��)�v@�GiXڐT2��,]��~'e<��&�lT�%;��+�oJ��oi����K�[��-�%w�v��n�[@��U�c/�|ԋUn>�%�4]��6�p)H��|E�F:����Z{�!�9e!eB�gHf)��j��h��y�y�7 AəY6�+��b���7��n��i�ۼLİ3���ӝY���%-�{�	:�Z��쁨첰m��f��;CLj��<��Pw]r�#ג��(�2ma�Uu�=������"�U'D�#���_��j!_3�%/n�`�3;꠺�p�v:v���i�X�s9��w�[I��N������Rd)kW�5Xu-����a�f�Z|;�k���f�A@���#���3��R��y1_ U�����,�((�)�(��
�
 (()�s����u9!AC��QKQ+@d9PVXUE��%!@��9�E	AMRPQT�Hd%-�UD�HPĭ!CVX�PRd&M- U!�cM	IJ�҆�2�J�����8CST4�44R4PU
��d�IEBR4RR�f4T3!@�R%D�-:��h�
�5(dLM SM#H�)M$�%+��44�U@U@W�:�2�ڽ�^��yS.������T�Vc��C�<m����Q@��v�7���y\��C�Rj��7�}������v�U�	����a�F�n�DJ�_f�tsp`��N p��]�df<d�}�{�6��4�qB�z��W��v�����t���J�7P;�9'���Ӽ�+��EC�=��{n�����~�2l�i��b�+@g�6���������N�gյ�)�y�"����ɯq/��{HϤ�]OD~�s�o!G
�	������A�5��f)[�~�j����{��\����ҪW%4��a�S��ONc�]�MyV�G.ѨzOk%Q,�8��T_�%�頋�֟���&W��ن��h�L������֔�t�sbc!�<hg��u���:k-P	{MPb/���Ss���1���%[���k.|������^����]r<I��Yp�q|��2��
5��c��B��f��Nc2桖��[3���(�]�S���/�z�<���C���w��V7sbv��������Fm��2%/VamIe���~C-�B�m��`<]u4"x5h4�ܷ��8f���n�"8��ձ4TTg8}���'�p�A���+���b/���>xm_mM��S+������H�6-��f�ve�36؜j#�V�_N�{���-�����������q��`��S^��is�����h�Fu6��.���D<\�]8Ac���x���gŖ0Xj�ijN�����T!
(�}��6�	5���暠ۇ�ޥ��Ea �p6P��u��t�����@
��^��^�K�~�t�q2�ݢ��P��}V�z�7C���e	#P�BMZ�D����d��<Q+	�?��?yǯ:�-B�>!�ߡ�z�X9y�ycy���!�X������/`�kT�u>~'h��x	�T��w��
������ig�\��ps��Rg�za��T��lb�U����~:�g}�07�<�ɪ�%V��ѵ��U;���}��7q�BuZ��
q��]B�������.�n���ixf̭4�v���BH�c�{w���U��[����s�j^.�s��[�m�G�>yf�D��B��p���-�i{���H>�qS��%�m y�1��`��]=sjhn��%7��	�v�����ӓ��}n4$���O��Y��Ҋ�{��R#�
ol"}�ν�Z�����ʗ!�g���[9c卟�5�sX�;��n΁ ��]v���i�����772n52QT�m���lI������n�\�I���!|��rޡ��r�n����v�`���[D�I�`���ȹ#���i��ww�ղ:��G�ғ&��I��L/�V�_P���Y���H��>K�����~o�ت��b^���ج
r�*Ԋ�*R��S'���?z��AM��5֠��x ��~5y�t���T���{aH閺�j{,��N?c�LS�m�ez)���! �4yr�V�	~!p�<%5\��>�+G�-x'H��\�LWޞJ���0����{3��� �ϗ�D�kh]��n����
d�*a�#����B�����[���j6rQ��|r˃���x�)��b�v1�IF�Ý�c¬ȸ� ��7EE�'y�Y��ƥ�a�@�bQW]J��}'J��������z��O�H�z@i|*�{��0�뺤Ev���mI��2���먽g��/v�eN�|_�����lO�_$OZ��R����M�b��>!��"�eٝݎ6��W��׽�p�ƈa�L�
|SH�_+�8h���
kh�Ѭu�O��ў�=�8%0��!�a�%Ḍ�R��Rb��f��s��T��D��p
��v�g-2Y���29�(�p]����f��Ff<�i�*����*[u���q�t삀�M�x5�]�x���{��nđ�Ӹ7��5��t\� nKE__0h��o�Bǧ2���K��y���Y��7_Xo�z��]$G)�Yё��Gu��?w��!~�me����J��!jwr.`9�nX�1qR\W���=�{�'��suu���-
�e�~k���ظW�5�X�.	�߅O'A�����0lz\;�y��ҫq�0F.^�����4)��6���Fb��o�B4���3�6a���V���!��K�G"_�S��WQ:�ף_����lӡ�Q��tv�E��O��z�އ6+rJ���7�Mn�m�.��4�d��w����|�L�N��|����a/���os&�h�w�g;[�u�k�s-�UM�w��:R�[���{:��6���R_�l�p`����O�f[�t�u2�Te:�|2h5��5`t�\z�߽�צ�ctw̦��{Įח��S^�������٘3����鰑�	�I�Bu{�j�+}�joԭ+��"�]�dw���,]O~��
�L��U�DH܅�{�/�>Fq����hh�s�EI黪�w�vڝCY�'��ͩm���%WФ�5P�C�q�y��qz�{�4$��\1���Qowg�DR�C8%�f:
n�ur�S%+��nV�N��k��*2A�Ct0�P�y���\�TZ�K)�л��M�֦���E�N�:���)꫺�����]A,ްz�[:��VgP�e�0Vn#.�`���7O��9��[�|7Hf���ʋn����9 E/��í <���϶���OMγ׫ɳ�W+���Q�����¼��G�AY��r�$�bW$x�h��\V�qN�l����H�#�SxL�2��+Oؖ�"ڲ�L���Њ����V3���x���^es5y��8��+LN��m�gh�_jT�~X���UG �&��C��I�@7P/�O
4�隁��OG�m��PNy_{�p8�v�/:(��ʇ=�ے�8����3�x�t݅�R���s�ˌ���p�� j+!5�ή�"N����c;�W��j>��]�M����DW�����Rsþ��ON��p��^S+ӆ��4��{=�iC3�2Ǵ�O�3�3̾��G
p�W_�)��Lx���9�S3�SZ�΂��nn>/�+×�J�_rSN\�7"��_
,��14������E_x���_P}EU�+��t�va~`xAc���+�Eδ���L�S��v���/ƽj�@����U��#h_XAj-�N�z����q9~���=�R��mfИ"Lᛥ���*�v+;Y|�|'�j�:�6//��r���BܮK�7�Q76�m�EuǤ��0r"��19����V��7�*y�J���+T���氹ĵ�{�+eW����*���鬵@%��"�[$T,��컻7&���b��w)�'���oF��;�>���p�w�_Dk�X��W�%r�<)�6-s2T�=�I#�z���Wxח/��sG_�&��pq��W�W]4����T�܃ӭneI��}��Bj3U�-�����ojߜ����0/���|O�Yv%q�Y'���:Zp
[?Z��Ͼ���P���G>jN�>g�T:�B��(��Ʋ����i���k"��
	 jټ���y9�ᮚ��?d�����'��.�R�<<��qF���B��� "�d
��oɣ���k�?��UԾ�� ��]"`���*��1�RZ�^��ŗ(���.����������I���c<�7�z��C��p���m�ő�M�q2_��
bX�C�LB�(��%�S�@.��g-�fx�,7�y���$�û���Np�=��{ݴji~%z]WA.�|�$۱�ܠ�xA�bj�qx,~��+,vl}u"�n���xD����x�v#cej�W�~��s�y��	8�N"p�<��N�� 4uK/,MP�뒖(X�8_5R�UI������y,�h��ّ�K��	�/
���5�WWf�Yj��,���A�{��gi�x�5.��橫�^��Xj1_��;�c��~rj-˫׼Y1����[�_2gTo#��_z�uy|DӴ�y�č�+�u���`�y���ʙ)���O&��X�ے��t�v�<����5C>괅z���<,����yׄ�l[���'��{�H�<��'���2m��q�&�'0�l��ΔUa�����#��|gB-C�mդ�^���(`=�xd��f��/�n�z'A�-�q�!�|K��.�o�x�P�@�"o�X����`�e��]f�	��&�Je�C���M]�{�pw���&"M*�ty��rY�P=����ˁn*�yeE��aü�$ ��ce�=,T3O�g��/{>�V��.��.�G�u�T��kj�>��zn�`{���M�Y#��ʘ/��O��(ZsMT<ҫ��Y~�ݪ.I�3-y��^h���'�.zH�*ah0����R��Y����p�^�rO.}�(^A5qۤyT����bw��WÝ�b
�/��~3%E�;�S���Z3�h+���T�,H�u�$m���&�󸽳c����d����2����:.a��7J�%�@��&���I-��[�v-�f�H@��H�LG���B�ҝS���Q7/�\B�q���f��ф��Q���&����K�9Z�quۋgk�k��V��uFf�vpO��t���`fB�.�5U�@zK�8(�>�hF_=}�l &-���_9��z�i���{���x����>�2J�%l� Be�7/��O]̵���q���\ٌ�'�2���:LeF��FӘ�[��K�O u��!�Tp�)V�H7+����+��o�5lyyV�f����懼t]���{
8�`w�����a�kܯ�,{�4���k��ɞ��/�a
�B�\�eʵ\1��p�ozD%q�I��_��ԣ�����|�s���
���tUL��ʒ�c�Y�HMu����G��ULA��CZR�i�~��f\r�5b�C+dhS����;�Q�uҖ�CVF���g�fFm�V��ʽ^pÛ�<I	[�ę���S��WQ;o��%z���٦=
?��V��ڷ�Z�d���t͚z*ڄv��:\9���{p���S���*�^}=3��k9AaI�΄Y:�z(��K׾>�^["'�ٜ�^1�W���:auK5gr�9�ԺL�]��S�a�(��m��u�����鶲�`j�xr�����A$��`PY�O�8.l����^&��3|���ƍ�|����*���{�+))��WJ�
6b����5���:�4@�pI\�H�`�ګ�T%�%ˠ���c>;����}�D�8�o�;��V0X~q�*�Z+!Ǵbc�c=>�`t�_��g}�CҪ���svg���nZ��<:j�U
���x�6�3�nQb�Wb��F8�C� �~۰�׉�z�x�����G]�(Y&/���2"܅�H_��� Ww�$+���3��R��9��K��X^l��u_'�4J� ٨���*�����D/.��lY�����9j���q7���ʘcp�!92��nȹ���\�HK��#���M��^�t�ݿAQJ7�촎|���-;[Z7Щ�f �)�sP��>�wv�T$���cnz�֦4��.�o}�Ɔ��DĜ{4.)�1�2¸+O�Im���j�>[%Xu�Q�1X�l�n��K�+Q�A*���i�8<���۔����a���jT�g7m���vB�n�W�0�^m*&+�a����K'+�F�i��A�w�V�j����w;-7>}^��ٰ��\�5��^��&2Q�?Z�N����6����uL�A���Ab�g=���ͦQZ���=b�x����,����N��t�D���M�bf�o�\���WYli:��G=�{ �8�Bb`�N��S)N�\)���h�]�&㨁;y�*�&Ӈ>ży��F�R�ډ-�ɜZ��M^��Xs�]n��)�\ȣ�$3��]��9&�RA���f3�=E�˄��^��b4a�cn��L{��#}��ރ������#k�:�,��s�5�ϰc�FI��p��3�6�Q�F��R�]��yC�z�W�@��Z:5l����������^���U9)�7��������{��ϯ�d�gզ��eV�����8��_0�������s�?|=�2�����$������]�&o��П���3r�MJZg���Abt�FZ�����x6�j�+��;u�� �:c�x��^��~����ˮw>u�"�N�����Ye}]PQ����XS��Ml-{�g#Xj�a����LÕ,yM�����;ܪ�^hC}��7�Fy�p���{�������t�NW$^���^>�x~����y)����4n����]��׻�0=B.�;�_J��x����}X��j�i���l�m�B�>�̥���ٹ����Q��T��ـa�"��{>��B<���؇M_��.�,�E}_?/V����R�V���M��uyfӾ�6�:I�(�C�]�X.�aՔ;�/
,`�-7Jŷ�2�:�3ս�0� thEf����n�u��t�=�ir��0j��n��b�bw�ר�`���A&[T%ջ��F*�D�S��:�d���(��MoXֻ98+ffe��C:� �=�xk��u��&�<��Ƕn�`Ve����떤KU
��U�u3�t�,ޘ����o�����2��)�#ݥ�Q�C���1t�;qZ��J�����{�b��|�_*��]�,�SdQ��䢠wFT-��I9�n*���/i2!Z2���$����I�.�� ��i���g|6�(_c�Y�-*���o<'ͬ��ΡY����w��vy���8v��	��m18��2e��[�L=82���*Yz�#R���K�Vv�
hj=��xtN�F���z�a1�l3`�,��	 ��(lꝍL��ړ����X�]�Z��d�l���v2�r4�ب�T��Tw��p\1CӵLY���CB�eC|~2�ù�VWS���愦�9o��c\ơ��+�余ŞDƠ�&���Q2�T-���#������Op��8���rJRr�Z-nT]9]��$=˸��ed�/��EL����S�8iS~Z�p�d��۫O1�����O��nST�^��sϭ�x�AS��L�.CdW��C*��}֍���\=w
�:��z��0u������1�{4���3W����j�
]v�n�
e�5��GS�z��^�<6]�Gbq���E*�d���OTA솅�r��	`T�VǺ�1�u����(���cj��.��M�kt��SF��(�T(U#��r��Pѩ��:s�,��<���T/���̄����ڈi9�۝�>|	�v��1���3�5��:�N�sA�<���9��g�jܨ��X��hs��)��s��4+��Z��؏.�t��nJUy���9|,�YM7MUͣ�j�*�K�d���ow�ss@�ucOyboݔA�0)r�}۷$��A�����X`�pp�*N�z�n�N>N�Ы�
#Lwpݔ�u�N�g�U(z�b�����="�ݗT벡����މ��n����P�4-����`��f�"�'�يU���ʊ2.E�\mheCD>=�&vt���qݰ���5�5S0��a�kZ�+Ow^.�`�O>�7K�^E�0֝�Qcs�J��kcS�������c��%\�Vr���+f��Z�o9����HG",�6�j��Len�,�#t��,�c1,7Y;�K�C�e���7t��i��Hv_e�R��cSpX�U�q?wbn���f�{��!;۝K��Ju�7eNا_�:B���m�����/(�r��\\WQ:C�
���W,߮�oo;Q*�������2���M jr��_n[�.�q��W�1�	��� AmuÖ]��p�"X���\����"B���N��R!�((�����������$2B����iJV��
i((2�������"�2��"
C$,�����Ȭ�\�2),��
i��(�(�*�#Z
r�ih �S$Jh���C$�MB�H`�R�S��(dfFLB���Ԇ�H�
r\���))r��Zr�\���hR�\���%
U�h2ʓ L�((\��\�!�(C!��U�������v�1���=���q	gq�a��e�{�	��ۦ���S��ۍ��tHU�Sj��F���kb�r�l�S��Ǻ[�������S�;�asI����9�&��#�5�05����y0�ܺ�BV���b��A�:9����ϰtf����{/G�u�r\��"����<>c��V+�.�W�{w��9γ�{u.�U��M�2�]F���pNOr�c���BS���%��M��5R>���#�u�'����9C��=sS�y&��9>J|#� �G�.Ѷ��*>ٚcoB���~�?y�y��&A�K�?{͍y�R���r|�5�����~�'%��+�!���}���pL�A�1�u���Ir�R�>�ѩ��MT�!F���1���1�S~�a��w����ǳ�<�A��_?}�7?A��z|��A�%Ru���9�������F�K������$�����hy �;���u�.�P�|�	{��ʘ�G�1U^h}Y�\f��h��?aY�:����9�:����\�w��~b��T���6?OwP�s�'�Z�����r�$��~�ԝ^��J�����A�nO����Zruw?}���^���G���i��`��.�y���[���~��;��9Q��x�pn���tf��.@}ta���O�r<��n�]F����7�e��w�lΰL��΃�y���?BS��߶��-M��U|P��ɔ�t=�����7���\�	��a�?I��?�Pt{���5&��;�Z�U?I��_���/p�������kA�d��5��:y��}�'%�u����e�5_}�p��G�"�^�)��T�/];;��sZ��ɨ�<��%?y���%�|�#]���&�B�?c��9�ΰz<����Pw}:ѸJ}�����}�p�O��A�A��[�o��Ф8W�M"*��������~/��*������fq����B>�DG+UX~~�C��cB_��{��>���y�a}��<�%�:��A��w:�x�P�:��g���!��֧��������}�w�jC�|><�?]e��.�..U��Π� D`���5����kݎ���j^��s�غ���>���*���p��� �%��_{���r^~�#q�]ڞ��`��K��G�b� ��1w�sn�~7��Y��۝��/��{��m펱C6+y���ǵ�����G\���3Z�������\�m�VdȘT���+.B8�#xǘhEu�_eX�,5���':7�4�-݊�!M��Z(�-
6��]�����7dZ��{��ki��u�:�_�}��㖞y�[���C�A1�~���Q��E���z���ښx{ޗp�>q�{���.k��꜏d�{�����Cs�}&���ϴ}P��N�ӗ�<�R}�y��֣�u[�~ϵ����uu�Z��w�����rw!�h~s��dd�]������9�܎F��ݯ�{�d{��={�B!��	�!��1��\��8weC�Oޝ��[���|�P�Pr��p��A����pFI�l3Z<��P�������jN�ε����K��}��|� 7�������?��t��"���H���YM����辯oǹ���{����>׺3�'P��sϴO��%?_����W�jfEq��K�Zr8k=���r�5C��غ����O!)�\��r>B#�>�f-��{q3�]��g}�9��w���e�>=ޞ����ڞ��ߴr`��u����9]GoI��pL�ϰkX����y9.f���s�(3�=��ܹ��c�5Q���=�r�X�s��g��G��"�Ѩ���{���{��w�{����w�C_G��>�F�sXv�����{�'#���Nu�d:�{��r�׸&\|Ò�5���a�)�r����c�}��9�����j��E��x}|�C�{��9�?=�Hn|���w�6�BS���6�?O ԇG�kp�C�?o@o���j�?g�N@w&G=�q��u��p9�K�Y/i^a�lL��қ�\?}�Tn��y�9����.@k�4K���\�=�<��u>~�K�}��C�~}���L���>ߛ�9;�BW�a�G$��5��hwEq��{���X�w����{a���sRh}��H���"Dt3�u��18���%=���^���.�g����:���}/V�����(}�.���l���2�ߴ��l��G��W�~���^F��m�w��B��#�D�����1�ё@���'�`rw.k���ѩ5��3�n�#�:ގ��BQ�x}��~�Ru�ZM�����䟎���ѓܹ���ޥ�?A��ߺ���k{��^���f��*n�6�.yC�;F��`6��!��8�|x�K�rĸ&.�t�s��҈�5��ۚ�
w�q��]`�ݢF���u.�uFR��qY�R�imh�)}�\�ȩh`R�&
�n̮*G������ﾯ���իX���}��G� Gߡ�Q ���5�u��S�r>�wv�~�nJy.A��:���nL�9�P��A�N�����Q����9	O�\���~�`Թ�uR~�!������x{�s0�㶷:>��DH���!��ђ~7��2>��P�:~�G ���}�~�ݏPr�y}��:���}�F�u9<����?A���:�kHjG�".$���A1��k�n��1�*9ל�����Ϸ�<�cRk�����Ԛ��Q��zu-y� �%�/����O����]F���={����=�A�BUGG�i9��5E�9.�>����G�>���!���B�)X�7�E����z�pe�>3��B����w�y��eѮh�^f/���3�O��`�zw�m�*��~kp����sX~���{&���sz|����v#ϧ���D��5�}�q|kB��O�xy�ﻝC���Oɘ��������7�d�'�[ǹu�e�0ܻ�2B��O�r2_m{��3���}���䔔�y�zL���}&T�����}����9��l���Ͽ`��/ag`G�y��5��=B�(ѨJ><� �<���jN��5Rdv�XЗ�?A���n�^@{=<�rn<��Rtg5�5��{��=�gP�B^��}��:��ɷ��6w��Gfk޾����y��k�d���OϿh9A���{���
��W��������N�ɩ�5/q��&�Rj�y��%R�EG�j��a���{�%�y���BS��u�/���R+�M�}�f_�f�G�DH�� #��ݯ<�������y��꧹:����d{/v����伇pe��}��:�
��5r]F��9�nr\�^�#q���e���a�*���~ߏ�sF�}�Ьw�Gզ"G�>��_�>�?G�j?<�폱�%;�����A���p�O��䟠׏�lM�C]���k��'���Zu���GA��˚̐��bPj2^�y��w�<�<���~a��/��{�����T}�{~�%%93P�Ƥ�L���h
c��?{�Ǟ`�>A���m���5	e�Pw:�g�5�����'�g�n�Q��Z:���� ��\������M�b�X���Jku�B�&\��P���^I�f�Z�.��/�� ���J��u"����Y:��Z� ���U����ڛti�a�;'�˃*[5�S�l��USwxk�Æ��ͣٴ��l=[S�M�rŇu�_�}_}TY������=����w'��Ժ��y� ��+�N���u@oxk��_#s�rܾƉ~����ևp�{�ӯ|۪���x�����3�#�����u&��H�2��G�G��H`�P���87{��~w���*����A��B[Ǉ��϶�����p���'Y�����+����s�����]{���s�;�r���^����:�!� �Dt��� � �Y���sr�^y��o\�˯�A��u���N��s1{���P��.f����*��15�����[�2}��k�h���Jy�ty'#�;�R~�&�~�/�n�e�x�h}U׏kF�j���k}����:���|��2}��.����?�톧%ϳ >�5�dd��}����\�� ��))�<�C�j5'py�����;�Ga���d��ϯt�����+��v�3f�dc���?�K���}1���P��>��ѱ�,F\'�b�4�L��1�6&-�XwqR�u�[3��֏^]='NiL�m����"O� ��0_V�P����h>�jd��~��v�‧t�z�b�Z�~ai�7����^�y����M9u�e6��yQ���/����j˽>MvxA^��B���
�����A�'����񁣘����=Y��A{�~lO���bQ���d<����i�`w^�ǅ>�gaY:�����y�_�P���[���bs��oʲ���R2�p������G��a�U�n��l�W[��Į4e�Y;���s�n�H'�l	n*i�n�P�^=��2Ћ���(�[*
���c��v�w�˩u�g	�Z�Z;�Vp�ݚ�ΦJ�d��N�S���L^LJ��TyL
�[디���Aގ�S�UW�}�0nƸ�xG�e�o�����~a{Ρ3Z�^��mMh�I�|� �m6;�W<G��΀ȡ��ퟐ���B�*�BJޟDk��Ӄ�=����3l�} �(��K�>�빪ʛ^�ױ`Xd������S/�n���,h�c��5'�3��T��TZ���7������恺�]8�@��{�
w(/��h����2@�f�X�v��5	�4K����
�?!�����8�����#��p_/<Nz}Y�W���l�2bُM&� �OJL����0�c�2��8�S�@�0��b6�+71}A��Q�T95�n��f�E���@�lڙ��	�:����/��ˬ�oW���r��l�7��֚�*�Y4m�@k���5T$�:��e7���g���?AK��Y̑�
��^?zw)��}��p���v�y����[� �yf�w�[�^u��)�%�mB*��,6ڜ����.$o^�j��X$^z:z�v��ʙ�����J�hVW�b��3.�a���P5N��j�xW>S{06	U7}9�"iD�x��[_,�=q��0͕�5�}:-ؔ�l�� ������#v.�a�h,b�e��",�`1W��[]Xb=�|�`
�����jw����|  ��5~Pxh�w�*͖����ϻ,$+�nW�d�nU����u�/F� �[�=%�5;7�l�0�/]=s�����c��ոГW����_j�â�x��w���ѓx�^�װ�po2ȸ�u����Gx'�t0?ju���|K�˸��{Ru�x�~H���^����9Q�o&\q�,�j���~��V^��i���h��1k��^�����[���X�{���SK�V� �u��E��o�0^6ܦW����!zq3Nغӕ^ʫɽE�-`���
���bbik�2G������}�����|.��q��0	�S�m,�~z��L�{B�G�,1(�'A@\�H�ӟm�D�����xX�aP��kx��첻�����	���,h>4������@�3d�(R�&��e{�_h�yEA��FLg�f�\�}Y��Y����� �*�sA	���SQ� �O�!�8�^�5���-�G�����8�,Ќ��_�'�G�\��Ϡ�W����.�A�S$��Oj�c���O�!^���8"Uw���/*ŽػYd����P�b`鴚��Yǹ���:~�ؙ�񚈦&JkP(�S�=֫�ms$n0�Pw���s��%Ԗ��a��uϮ�w� j�t�N���5�_^�x�D,;��o6��E۷ݢa�������2KMz���
��W���l+J����I��}��{*.Ͳ\)��� �g�kF��n�W�����v�\c�lӽ���5Ԇ��ӳFۘ�u:zsp��L��$�J�ba��ْj!�N������ˍ�/�V�+x7���{2�}/ngnt�E��w�y��i{9h��Y��.�x�t-V��,��^WfV��6��4,"6of��/S+Eg��Z|�z*U���^4����;dhS�<M��f�eB��4M��-Jmh�w�>u�g>I�Vo�t	k޿`��ݞ��3���]\&X5�}G�L¹D*,[S��:���M���q[U��KD���gׯn�M&Y8(y��5m��٢�薧x_0�__9�kR���a�ޤ�]�D�����g��Nc��oop�r]&oF��wKk��]�G����A�>���+���%Ad4�;�
�`t�{<���{�+;��.�g9��HM4��Ϫ����`Wm�v}Br�2�����gto%�GC^�h��
�q��w��;�ǖ��8p�C��L�R����ɍ�S�L2�n�h��� <�d�s<����Z���3+iJ3�Hb�,a��Xm����ms]@�f��l�	&�Q���ޭ\A�Jޮ��olV��g� |:��R�bO*p!������ګ���H�%Q���2"������b+��ڞ���5lB�����G]?k��c�!x�Cͩq���=�z��5�o�}C��:g�X:9(.	��B������;�/߆鿊�cp�92��#��ѫ�L�!�{)�/��Ӟ���H���?��C dFP�ӧ/��"�4�j����>��:,l+Ѷ�����KP�Xh72Y�u$F�.N���1ye�ei����V�za�Gh��7w�W/�o��?�V�:OJ�rPJ�҂�4��py�=���|=�̏a��fs^f�{��4j���q�%C,5��%:���F�i��A}q�����+��!-υ?6��1�y�C�	��7̀�D7,/�42˳�Y;Q ���M�������Ҷ]��&�8�y]Yq墑�S3�0�'w�е���Qb��m���J�Ƽ+E:�.�`/�e[�ګ<*_�_^'Z��O�玵Ԍ;0�I�c+��W���~�ؐZ�+��Y~�U�&=���.zu��^]z��K`�)am�$>�A�^�d���e�R�v�P^�a@>���BJ���=uم��v1�_]c%�{ �\w� ~)V�ٔ�N�od�x̡�EC��fB��u]&�%gtk��}�3gb;�پn�(�<|M[5���c�5l�P'K'����5pJ�.����{�VT~��jz������(���q�.���{O�va|��M項�b�zo�9��zQ�U����~l���.=��x��ύ���p`���j�H]�,U^k2��bMf�5���BC)�+�Y)�܇�bs��%o���a'�wŕ��qM���%�uQ��0��;
��Xc >�Ub�x}�����3�1��W�B�0�\ps��ƥ����C}�`d���&
:7M	���oN�x\a���k��X��LJ/P�Z[oֽ�A�{��Hs��IO�uI�N~�X�aƬv��jNAp�eU����S�����uHB���F��@P!a"�%���r���uo��|���l�'�mP�Z:8v�q��~ɲvy��^��Њ��4*0x��ߓG>Du{]X��L���L�~�m����[p	��r�ǃ&�u�[�q5��N��5��A�^eoM�0Tu���	�W��8��H�j��G�u�c�x�M�.}���A�-�tI�n�5b�`�Y�1i��/Y����C�x�Q�=�J�+��z9йr2�U�LN��yKƩ*�>�{sn��}�gby4���%$,�}���`�O�j����3��������=�"���w��J9Hv%P��Aj� �a*����ހBfj�����^���\��ⶰU�R���6^��Oo��P�:ɣm�Z���S(�+Io�O��+~��3
��f_�v��R�hV������R��8����jwhǢ��M[� ��Z�EVy!z楓P�棞�>�-��|mg�s`Uc�ƽf���	�W���& �������nZ��7���}�Q�z+�;>~�*͘��� ��}�	
�[��4�a]�@5�1���E��o�.�Cp�~^~����6tw�|�b��w�{���A�_;Xȏ�ȉ�G���jÝ��%< w�l��i�6Hb<�'{�]���P,���%���,����.��:k�Nfc|>Q.8X�>�@VK,��)���������l�N��
ֲ�='��IZ>�L?���L��+��`yY��d�E�L�3޾�����l�U�����M�	ۖP�3��q����WIk�+$~|�r��������y�Wվj*{�qb�P!�eǥ���H)�,�i�rtf�e�2�����@]�$K;[�d���R:υ�ѵ�`�nڂ�]��l�*�F�Q�.� l��U���q��17jS7rN���I.��E3�K��br8��id^[��D��Y�[�cbA���'���-9I��u��+_\�/ w��͘�{iI)��d�ۺ2\��k����r�#�1u���Yn��D�0�6��'L�R��eK_BĨ�C1�Gs�#��.�9�����|�ijv�@se�\H�Vq�ك�1\�]�h��8m+�X'��;j���1ۓg>�,Vb��ʖ![��dݭ,$M2�b�P�}J"2G׫�~��V�Y�5�U��wQ���U�)
 c��kNL�BU�ܥ�ˑ<OvƱ��������
����Ep;u�s�H�7γ��`̛׸)���:�|�ĩ{��Z��z�Z+@wlK���+Q�Q����^������ -��;2�X�l��6`<�L��`䌫YW�EQ�0H��U��t��K(�P��s�Y�)1s�b���Tz�a�1�,v�i��_�U,�9iDVF F�Vܖ�W�_Z2Jx�oSK�U������m侉#�nm;T�9}��[q�`k�d++�[N�˫�B3���ylV
�r�݃.��j�@2�>�Qr+��3���H��mw&x8{]�,pCth²���A�-����:/�^�2FtVӓ)��x�Vnd����� �n��>�:����R�,�	�]{�c���{{n`!Mt����/�Pg��徱9�|J��Jo���ܘ��z5�Ld�T���Ė���8Ï2��.�R�wVowG[EƷQ�tʏF%b�������bE����2�'�l��V���7�������5^Eq��
{n��P��S�3YqMDڔ�j^'.Wib�y�!�ŋ��v��EWa#\���j�ح�K����޶]��|���[�èY_+И�W�m��m�!J��.K�>��
��ܻY��}Q������e
p�3$��a���fd$=x��i��td���ꎰ�Ȋ�ݠ��L�DE�iwN��?�]Y����:ã��z�%Y�_R�ֳ�燧ι���VhM�wwS]���5���b���˵����J2LbE����o�+��#ʎ�t����M^1��ߩ��7�:��A^l���:���wn�5w?��U��!�����=�{}�Gu�U�LqT�ua�� 6*=��
��K6�*;Tg h��wco��:牕�7�\,��K/Um!i ��E�®TվJ��ڱϝ���YR�Ǿ��6�+Ȣ��*���V1w�]����4ncC.ٝ`��H�V��bws4K�r�M����nʖ��c*�wr� ���T[��>ѣ˥Qv�7�B�׷��P�����e�ީȆ���c������Ng?��}�b���)�(�'%)S&��(��2(B��
J�Z%\�B�"�T��
���iJC%2
��JA��J�%�Q�BY�ҙ5��J�R�J�BP�BRS��!�R@	���b�R4d�Y+@�.J�f4������A�	�J�4#�BD�QHPfcH�FJ�PPdY��C�J�I���9���Ug[D�蜺���l<z�A)��]N����<'5/F�c�TҖ�V��}Op��C��^R���s�����NC������+��07�-��P��.8I�x�!�*�3dt�^� ��&c"��En�V[;t(?�z�0��>�ƃ�I۸~��@�3d�(�2.'/�l~Z1K��A��%����7��'�R�w��Ϩx�}�vɶ`p�P�J� c�"2�?9k=�*�	�F򤇺���н�4#+c5�BN�>.pCg����� ��V ��d�����1�m�7K�̽�;��	��RAY�����S$o8�����A�s6�~�� �p�r��s�;^^9���	��tR�zv�Bǆ٫��xs���U��~�w���1*�֫3��~/�w`7������L���m�¼��q�����J�%o�>�����/\�U:��-�M�����C�
��s�	o�Vy���q�U�(,���vg���zz�ج�CΦN�6s�\�U�f���2�Zr�b���Nb�}�u"�N�9Sƻ�H��/~���
�|:Q�֖jc�<=�2�2���@!�4�15u���F���Q������͆r�(S�6�cc)��Y.�rQo�Չ��^s�ړrNk�n0����h���2<��(�TԄY�ל�T�˪��Pa�o2��F!�\/6���s��M+;��ſ���Sh�]:��OP@\fvS<&�{b�'+s����_�� ���]w7+Ǝ�?�[��j\p�l�}37�nFS,��zq�j�ۆ�Y,n�f��r�Ҫ�l�xɠ�6���6n|����_q<��/����8���c��2����گWN�^Ƴ'=�j��O�{9��v�(J�r�Q�2��X��)PEzM���-FCn��P���um��y"j�=r��C����u����P���<l�R���}IP�i��{�M���-�b�;u=U�:�{L!�9{a;��SS�h�(�����zaA¨z�aĬ�'F����<�7�}��w��?"����\<�����^��z�'�� 3S���֍6��m�7�Q��&"D/X����M\M�2��*a��#*-�#���i~�D����]�2�@Y�|��w���3��t#,li����#A;�C�X�'e����f�Þx��<�J�$��	0�Y��u��,�;Up�V:>��=��}}{�\ϰ*%+od4_u,�mZ��ZL����g�!��ސ���-��I�������z{B�jۃ����]�B��a����8VfT>�����gL���{]lؾ����\BL�p�k�Bbua�s��]b_�ˣa-��5�S�Be�C ����T��/��B�Qő�ǵ���Υ�Gpyi�3�PK�&��E��h������>�#�5s�xϕ�#��i�?Wɪd�,~��)�D�D����TTJ�`�����%��Xk�wJ�[�鍈MUɱ�@b��`a~
he�]���w�Z~�`�C�Y閯_�;�~�j&�|�]�Wf��tèX�n�ns��oy��D��f�y{0�C���ْ8���?O}x�kW<X�s�Z���=�d��g�B��^����֌�o4anH�/�F,84��A�����>'5�]��=R��5�ka5j]?m�z�Q~�7�hf8�x�L��p��*�!^����va|�����V۵���gst��{�-�G��~�zSe:���߫E�nT�,����TN
�|�'+�q��Y�}2c����@{͚��/�2EB�Mλ�#TK������ne�G��<*'��H=[�/׍s����+�*x��f��g�Sw�O�^�طMp�J�zRZ��.�
���sc�˨��U^�A�����9X,�l������_�x�A���vJѪ�!&��Feݔ�u�t�h�J���ⷽ^�������!JŘ�.�2�tB�inq�mǋs/.�+?&o����p�Rx*�pB��a�<����1����c��k���1���q!):��0�s޽m��Lve�Y�+�b��eY����è�_���}U��}O[������8���+� 0#N��ZS���&]9�Yc�}9�� ���h�4{2��^���`�e���j��W�Q�@ͯ����������u����v�z$|p�|�����}�S}n�G��'7��Y�K��P�;oచT��Y�3X=~�s]7B��!�Z��v��a���p
�ՠ˔L(f<5	��-۸������Da#ފ��q-*�E������e���?z�j�Ó�����i�0XC�L*��S��f���4��R揳pg�x�p�?S��^V��s��p9�d�@қoģ��UO�+�V�.r�V�ۙ��r �,�v�v�J������T��- �N=!9�fB4y�޳V.�����^9�!�n�\�W��E���[(*�½f���W���ؘ�´	M�N��=M~��u盭���t4��<�=�EY��@� l�3�ʰ��4�{,Y-�"DBǽ�{|m��@^����|ƺz�23��+��]!4���k��>��R���;w,]�3����MD��ȟ�����FX���~ʗе9	}��!�nr�k�+5�bA���?�r��6��ϲkj�3-�����Թe��gE_L���-�s�Ʊ����x�7y-�!]��i�X��(�Hr����ﾪ��㮝����~����,��G M�F���Mz�η��N�?ju�ﬄ��u����{��A//\J-�kW,��	�U3q�1	%�Z��)���4~������ƺ��=�xkl�����5#a�$ר�t�ѥ�U��F���hV�(���C4����~�m�$��������>���G�x�8�P>���D�$~|��ʘ7�~����p4���W�� ���*8��!�Sl���!?#���(�������6�[�bj�y�s^k�{�+ֳj���Ώ�~��{�|rౠ��v��zO����b
�d\H��f�ճ�n�����׆�)�x���n�E�wONboF�/ʀ����<����^�U�ӴTsj��`x�m��}�,��(-5�BN�!�l���x���.�P�O���U����˼N���[�$U)��Y�v���8�G/�g�{*]zϳ����Y���&or�B�s���,y<$:��e*�J�?�*�B�6��Wa��C�}��X�2��5#����=��wu��E���{+ 3AW�(-T!Y1��e�V4���V&3�F$�g�}�+������n��r�չq�wz��u�N�˰+��n������8���X�j����{�qj�y��+��eQ��h�JA�!wV�~��������y��W�#G���`����6JfЭ��Q�c���/�V�+��w�#�N�<��g�[�ӻ�l��|ܰ	��1��O�t�IA!��$4�yy�g�j\���i*["=z���YbҪb<��e5Lyb��L=��V8�x� ��_M��_oD��0�R�`^
(�YC+u�f�2���MS��5u���F��XC|�2‱��#��715�0�'p�/k�n��V�L::�~hx�o��_��O�Y���^�)��������ֲ��R��#f�%�n�_k��3��E^w��ULP;�epy:x��z�%�wX�~ܗI���}�Y�W�XxF��<|����v��*c�>�Ѽ�*^g��	��
�Wyw���N�ɤȝ�p�"�u�~�7�b̐^�]�o�5�������}�����&�ǝ ��N�xmUօ�raBI�~	�Y������ً���yC�?#m�����3���q{N����d{�f�2W�'ޠ��|�� �)���T}�����=^��oq�WWY4�T."�3ft6w`l��T�c�ā��W�|v�X��9���g�ne���t{;D�fY�P��U��刑��)S���=s~�,Nvv��^�¤�s�ѧ.�=�;���Y1F
[��X��}S�_W���}޻��<�=��6�9T8��Hy�eFuOLO���ʼ7���{Ћd����	�z��駓 ��a�@p��0Έ����Ob�{�i;�B_��5�,ļ�mnwa�b��{΍ϫd�,q'�W4Ema"|��S��i^�G�a���®�^�I�]���6�W�Oa�K����A.!i��{*�?��]^�ьĵ �gG�^��mj�K3���C$����N 9`c����u?iD�
�����Q�B�w@A�N��z��\Q���B���ǡ5W&Ǚ���cʯ�m��>�<1�s׳�G��8�G�><k����9�m�C��Hv�V������{˱�oM��[ٶ9,�Y�&+X�ʡk�:Q��>x�%��s����c�D��.��T[��Q�{��
�����.�ƃX|M[5��Z�ѫg�Ai�77 ���=O}����P1�K��83���<%�3����߃�Ќ�U��EV� ؕ`
�����Z��]�RVn����sm���%�t"jU����ǩ��Z��u�Ԋqo0�E��E̡YZ��@օ�ە%J�X䲆r�7��W8 �/�;��'�%�����=M9��7�,eJ�#�f����4Q\Vx���c��V�m��eD_� |�(��D��h s{x��Z~�z!�69x�̓�-�\{����>ۻw\��nʓ:������yš�_����i�Eǋd�Y)�܇�b˭g�V_�jrބ B��Jb�i[�n���e�<'+�1�k��}��{ᮞF�[�}�x�����*����?"�rٿG��먒�u^�4%��+�����Jޟk����?!�o�9�@��[ʓ��ƄM#�(Z���%#V��w/�ձ��<�O��E����V�b_W"��yAH�Lz���垿�HJ"a�W4�z��'H��z�g]v�
�Ng8)z�x��V�V����K������N~�`#��G�|H/���3�l����hp�h�-{P�}	5h{�.�1lǃ&�7X�Q91�䏡��l�P�2�N�*�d��Fm�>E��ϽHG)����Mւ��4�,!���vEa�=&u�
"�IS��Ǌ��z��6�ϲ�崬�G��q�s�>ϧ����Qs�۹�g�Q��{f�_;}!��}��5ڱpu�\�e��b@L�����]J��]���^����.�Wd������9��-���8�u�E�u�$�u�4u��}��l��r�4��_<��ML��؎&�^����{�?㦼hk�N���U}UT��:}������T$��W��F�
t< �;g�}�����k�r��xS�T䉬�tMRS>j��o-�ro�C>��*ΊpE\�R���r������R[���=���n��ø-4�7[��}������=�U�1-��@43�HW`�!0c���S��YzrG��.�{�@�yׄ�l�~�*�rct�g����hIZ�v+��H���"el���~�vS��f='}B M��"�]Cd�"�N��D\O-�~�1��c{�to<+>�ٽ
1��̝��w4����%<�=u߅LXd֩L��w���$E\�a�ؼp3��V=W���*b$�'��%��KګȪ�S��b�p	b��FF�}���>Iޕ�$�B�����f\%���� 㢸@�W��$~|��ʘ*�=~�F/~��K��!�wSC�AJ�sMT<ҫ��b� �w�e0�/G��{é�,]yB��	���|�wV,H��u����p�����S���[g�WÝ�b
;��xmtG���\x��Y1�Q�T��4�,:'�e��)��O�z�u�D��ģ.aDs��Y���f�/+{0,�^-N�s4��}K*�l�;���1&�y����Nv�Nȟ�oR�M���c���Wn�=�%[���"�����.�mE��|7Cy�>��B�^�Я�)�x��t�3��Li2�������<�Q�7��>x�7�UU�{��݋��q����f���t��Ce��7���0�*w"��/�����"_�d�*6����& !3�Xl_�0�f��1�m9)��&�TIB�ֵ�*��~�s��5&����P����C����J�ժ\���\B�L��ܿ	��Kمry��[z���¬�>���<@�1Q|����Z���
>����0�
���\�4���
�zU%�'UW�kwr`9�nXֹ��wRzY9P=1�0��J�xc�)ȳ�����H�x箤�f�/Ƭ�%T�,r���&Әa��4*�)f���x�=�u����ІU���4=�j��*����g��z��xM5LCG���N����ݪng��_����>Q��Q�%�@��A;f�.|�g���w��?<ۖ����U����72��G3���)�����c?U��L3R�tO�)/3b|_1�Vqp�U
��e��~̧�y)T#��[�%u�����,z�,��뜳!Zlk�)��7rњ���ٻ�Y8[͌��W��[�7iEI�Ӎ<�ilə���&6�>�����/��	ku��Ąy�N@F�N����C5U�Y��(�b�9#�|!P���킎9ԁ<E#S�G�ܲ�oY��=��%i����s���W�-�دRq�80��b�SG�ƃ��pL�\�Z�r��T4�u��Ä�]Ĵg97��C��Gr��V�(Z�]ט�;b<�� ]��lF�\��͡�$��y�����G���`n��_$��h������y\���%�e�/pXG��[k:�,ж/{�a&�� �<L�|,-��9$U��y�{��+��t�]�j:�rP���nY|1��R캳����s��D��͕&d�t���v��Vz�V-�I�,E��n%�U���y�{�u�R������gxAI��H�K�s��n����e���R�+*'l|*�J����
�]6����9�Ǐ�����T{�ۇ:@�tP,s7��4�#V����]���H%�޴�];�^rn<n�<�L�Tzú$����QUm0�#zF/��-�'I��\�z-B��-�w�9����l��J�L�ޝGc�*�L�7�b������O�w�ly�u	�[�x�2+�7�3x��'7(h��f�I`�R.� �E�g]k��پ\-+�Z�ɒRt�	�5�m��@L�����s�ud���:�!�F��9���޵ٖ�u���qW�aٻ�k��u�7T���Pe�S�2s���1��s��u�R3��O�y]cF0���3�!�t��s��xcߘ�Z�o�[ɻk�Q�X�5ݼ�+q�uv��f`�yE�Y��+Y"o�y=Z-��'pF6�6n�z�R�$^���b�4zu�ѭ�f�
��PԄnm�o�r�|���lx��������?�u�=	I)�^E�x�x�{r��,QB���Fn2��[�)��}�H�s*6��ֳ�P.�c�ފ�5�}nvW!���6e^Z���%J�6c��pQ�ڸ�ֶ�ң��ɚK}��LK���ј��NU��=�y�N[�UId[������{/x�h�t�j_%D�!�2w�Y��j��|�����N��; ���r#i*}1�zXˠ�kz.&��t�]� ���|Nn�5���[[ 2�}�=/�-;�`Z=����lYE^�9��%�(�6��Q�W(9�C8.�݇"i\�7�=?_
DlNt�WGw}������]����$c�����l���&�u��u�v�VK�	ծ�r��J���-%���ʋ��H��1	=�8Ok}�!�QB��[g	��@x��u`pӛB���p;º9L�h�_W<0Xj���F)�u����u�GJ5���WdZj�&��C�"��Hd�99#��%%FA�4�d�-T�2�
J)Ւ�:�ʗVJ�R�-J�45ERP�&Hd�@SJ4�BdR�BD��H�4�T�	HR�dd����d�@KJPRPS�9��RRT��S#B�MST5@č��9.�5#@SM��R����*�0��)������15����KN@�)��T�C��dD�.I�D�IE�䀚��������KV�K�t��,l���t��Ϝ N��=ݔk���ۤ%�P���z=��]P�����ͨ��"��iphȏ�}_U|Iwԡ���M��+i��tE�!;�c�� C�FP��XxF��:��q힦��2/q�1��g<��U~ܱZ�7P�:b.���:�ۺ�B�U
����`�R�4W�f�Ǳ�n�#���P(�>EWP���݈^�������a_� ��n�xn!-N���0�$��;�}�Gf_�\�g���yѕ��7�q,��V�R��!����~`���~���Th�n*��M~G��N���!p�H�Ә�ӱI�����3��rd��Û���U�{�g��qZe2h����wU,T��B��t��ӧ�E���'5��-�cK0��I\�i���#({���K�W	h�W4Ek�#}�����W���fCȲ5��~��t�����Ї�-�,����?��*SJ�r�}>���4]�7�����EX����ݺ`������Y[;G��R�K����}`Ju?iD�!x�R��؀N@Ӫ��`��C�4=���+k�N��>�]�Ӏ�<�6X/b�q��<��:�Ý���.���j�wi��L$�������p�	靶�e�DF��3xFpp��J��.}���(ve����ٹf��C�/lW(�ԥcO#R������b�j崴f�5k���p�|�2��w����cj�N�.Gm�}U�Tr�8Q���꿛�,7��h�e�����1�<hBĝޟB�@:>=t���v����e�:����gE��>��Q���6_q��]l}���g�����c�B���<$���D��3[�Z���|'��ռT#(�\a#PJ�ӵ5^��g��>R�[��[�O���l��3��m����%2��7"�_
zsu®ұ]z��5��r��ű�ߛ�عm�G�x`��\N����C�l�C��0��߫E�n5�}��}��iw�DLKX+���۞�qat3�W� �M�^��Kd��78����u��򬿪!mԌ��:W���f=�G#{-i%8� ߗ��"2��
0��L�4S����ީ��0�e#�]ک�7�����e�8Cq,[Z+	��O+�U]y�,�~���e|)���"����z��Y�M�:�Cqc�H��\hd�/`P@�dʫ��(Q���Ws������'�`�b|��	��ҁ[��|(Pp��r��gּ>���t�Dx�� f������zb�r��T���v*�	����/�׷��ԭ����t
�t��,E�����X,��WVl���q�!��ΑZ��4-T6��Ӓ]GewW!�O; ��V��'���9.�J��Q�lEa^t��I�R�nr�k�O7%d�՛�L������%�|{����|��u�s޷k��q�ߓ�[^��No��������]P���$EcG�E��nΪ�$U�
�|��ې�&G��V��t���b�%7>%��M���MetXO��?_M������Qr&�#�y`o>� :B�`�Y���>��	��R��k�{�.���{����9/�#x�����v����+'���5PE|�:ɣBT���G2mV>�n7Gj��¼�n	c	,�]�;r����ͭ���<�pv�vzfe����:bZ��f�ds?K*(��YP�i�5��V9���g<&�%4v���#��/� ��#���lܳS��}O���<�=��Vlķ4��3�Ϭ$+�@�Z��Q��-�=�5Eid��>��� U�a̓��둿zZ�Ύ�/�Պ�0~'���ئ�x.=1�s�@��'�o�r���~(�oV����|X�-�����~�ȣW�I>x��?8�Y�2bE�d�>�	�D�ǖ�Ϻ�¦ O��_9)����2�"��)�>\�pˀ&i-#�U.�S8���L>�v��9�G�y�*�Wc�g�Z�AT�!�r�f[�fs�m�ҝKC4�IR��S}�@ͮ�U]{6Э��C[F���é�V�[j-�x��]�zES7�ݻ�;_�>�!�ν��_v�������h��1hX:4���l���b�X�|	��>�Z����8)�f���-��n�˂���: �8H9tW ��-z1���7�A�{w�����5��k�{�6bA7����:C�=b����������R�*���-|nU
l��mA���D3"��G��y箮�Y
��##�Z����9�W�'}�Ϲ�Or���*�������^�@���~�|�w���uSW8��F�=���������`%F���{�����S� �DN�����D-5v���$C>�_��9(C�W�dz�_��om��uV"kfI�Q�'�l� ��.��8�n�7<s�$r<���O��9ޤ[���P]��Q���va`yU����C��e*�J�?�r�P�=!k��莸7��,u�p���ҿH�^��	�f����c������}��a-W_܀��!�m{��ā�sTs}��Bܑ�I����ѿr�{7�{�nx'�/)z��M�z�y�����XD��8yzx��\n���V@/���R�XM��20c�C�7ۑ�寲nZ;��.z҃W/OX��p��8�>s+Z�ВufO���9	yp�غ�3�"��˱re�^�^�VL�[Ռ���c�O-l|�k�(�DÑ��i*>��Gޖoؗ�������VSǾ�ו�n�)yk9��s��Umٺ�J�yU�^�ɾ�a���1w�i������k�*^i�^����WM7��ܟ7��jT���x�1vt�����
2/^���6T�����=�yX��R���y��R;�պ��Q���
�<��i��^�(1?qw�̱�?z��v}q�`�{�ק��6��tz!g��J7$]�{d�QƧS9;HY��b��i�����)����U�b�=�_F��혎R����O�L�R9�Uiw�%J�c~�y�ʆ�˅>�p*�f�Kol�>>�����]⁧慖��躉K)O���k/�U��>vT\�>S���ዟK�i�]�E��}�ρ ���C���.y�=~o*o�:c\�=*)5n�x�����Piz�5,?��5'R���kcn�*�8=���ԇUڥt58�� ÷m���a�H� ������/k���Kd���5�g�i�i�85�h�3�G>���Eg#e2��u������r��fS���z�m�ۡb=�j��N���6�ڗ"��q0w��2�#X��o����W�}�so�6�qzr�%{	��T�������{5+�ؘ`�<���g�V��*p��խCz�m�ϫ�.\6��?mv��[��jJt���r��g��Z��Oh�jL;����o��[��R�/�Q�����n_�=ܷ6�͜�~�g��7�ֽ�� ��b��9n��Z�EV+;XҪ!�#![����;�G9ݶ�	<�	�������6�g�������y��s*~��gҒ��g;O���E���u�߼���sej��pg�^�Oܽ4M�4���u�.��{��w�����~����;	w�BOva�{�S��=R�f�v��5�Xu+u��c�c��2
�L�[����-N�=��z�z�r��y>�{^�_/S|��_jA���Y��RM8Q��e8J��W-�$ߧ�����Ϲ^�Da�\�y�ۦ��$��������q�b+����B/�P63z°�v�Ҷ����E�t���������ZquұA�F�Q<B�G#�w�t՛��U������JDp{��F:ZE�**.�Mܭ��v���o�
������6.�}��#���O�D'���&��?��R^�‪<�+�c~�y���������3�Z�%ҁwΦoxVT��]f+��@�e�m��>���q�Z̞>G�? ��1[C�^qoV[�n�+�Т��CKo�N�㏔[b����r�{=��E<�Ϟ�eE�=Q�+�ٳ	`�f�r�^����YI����ܿ����?l7�*�P��"��-�����~ȕI	Ԥ�v�5;��Z��hʄ�W�ئ17�E�;>�k���^�t=m:�E��w�J�Nf�ĎRZ�z��ႂ��3�Rʝ�^�sͯ{X��B���m��m��r�������V���zCM��ԏR6lK[�����y:�}g�ߏ�"K9�"|��$�!�� ���u%;Nu��Ûn��z�zu���t.���wZ�T��2ы�X�p�Ԇ���+�w��.�k�x\�I�rz�)��rk������d�ܲiK46�/(v�%�{�i�=t��{��)2#�c����ը�EIM�"|��m�d΋&� ��oX0օ�X7�h�X��nG{���x�����,^=Nrҕx/�j��n�����S���݄�����C����.��Ra�K�~�r������-��vg���Ow���m- ���t��>��xa��ӝk�;�*F�/A���`��h�:�c�/�m5�1�ˆ�e���v�gOb�����Sʋ�h���N�Əz��w��tƭw����Of�`Ev3�1�k���]`�]���r���烖�~��NEf�uuAǐo��i�k��քzb���_W�V[q�L{t=���6}���㩮�̣^O�ކ�o�M<�Smؠ���Pw_�2Iڜ�׮�h˒����|&#���'��=:y�㪞�n��ނ>����'���s�g��H���(�gR������;E�ۀ��z��ٍn��Z)���p��~�6����=�^��T�fc����ol�LJ�e!�5�i�l
	V�Bm�\[?Oi���r	Fg��z�N��u�0�Q�s��^l=v�hg����Y���Q��E����x�Ѧ�'A�I"Kuʯ6'�	�:|�I
ꇦ|� l���f�Vu:FZ�.��\#\ښ�����t��≏��]=O���r�P�t0��T�.����{��|�}|��릾m9Yg�{\���=^�SE�r��yQ~`3�k�����y���O.�^�*9�ׇ�_'�k�i��m�;�
�q��xZ��z#���y�]���f�s�Z93���+v��jtiyÚm��g�c7u[���`��M?M^����l�~�_��M�/-c�5��.�>^U	�Yzs�{�6��E{�Z�;���=��X��jy��~��YSU�Wo�ۙ�^Ӎ6Jq���6�ޱw�.� w���|2~�~C�>3�ʊ��D��gK�e>�g�K|��-���=�J�H[S֖�8��Uy��F�?@��g��Z�=�@������'`�����k���o��`Q�e�E���X��Y���^9���8-_�-��c~��W�婽��g�-�<|�=gN*B�r��E5w$nq枃�Z�XjP9Rj�{��yl��/!�ؠ��=B�(w9.�E�F��.��0PU$���X���:K�����ؙ.�V�j��'.-�h��6CK��e򶖸	�9�-y�_.6و��6�G"l���(`�w\Ѻ���n7_�V0=�������+�7������yj}�h��*����:S/t8ZlHy�wVԖR����Y���ܙ06%��Pu�$�Qԩk��Т��g��:�Jzj���!$�O���[�xܕz���o�{ը%�]�>r����ߞ��F}���y�����(��Л��~����a��'�
M�Ty/ZԶ#�� �u�.*�)�W�5Li�<�3�{u��y��l��5~���I�%J3����)hJpcN�����H���D�zj3��N�f�Ra�qo~
�T����oгr|��Ԇ@�@˘9�	��7�+���i�4���n1�llW��w�>q�^zQ5N>nȝ�"���dB����{zfKNI��oL��t��|���+G���׽�w����e�1g��o;g���_Bw8��xͶ4��.I�0J�cs&ab��=����jR�nh�����&16qkx��/0м�2ғ@9Sp8��̧����jM��6���X5�ܻ%�����hL�)f�O{#���zz3��_#�.��~� ���&n�������:rH��\2���rV�>�ٶ��1�G����ow�W�Wgb$,���HQ�R��������VU��g ��JUoaɪ5��:�˷���HU �(l͔�&�-�_w$8�tt��T��ID�Z�q�~"��� 5e�j�uR�ut6�u[|���1`��������x�>U��뭓F�bt@�N���ݾ���H-�԰��%˞S�b�z��9���ׁ��� ]\���~ʵbŘ�q�\�x�Uu�IZ���c"� ��7��fKL-qV�C�+Œl�+��7;RЧv��ZڤÔ��d;�ҡT8��eSysr�_T�ӛϺh�e�DU�E��.&��Z�om&���}�|�ZYBi�2y����U[ur��gF����k����$D�:�t���ϫ��d�\]>�|^@���"�J�6�؆�Wl�{S�N,TZ��.���o`�9��H	&���h�l9�TaV<���޹6���4�Ƃ�D��b�0�8�+�Mku�3$�P�m�� �.^��䙊D��	��}���*Hv����Xq�t�*ya����g
��y-T�JR���+��f9��֘��Nޭ�s��Ò�i�2��$4����(;��:��
Y�i�� ���f]nt e̮`�)�u�wl�V����c�&��n��|�¨���d����u���6��0=��>�8�[-ʽ%�V/�|��U�8.X���b<�p<2ˆ�u�K�VaS�ۻW�Ӊ�Q��XƮI�f���ՇP�lMY��4a�gf�Ͳgκof�C �N�5�X����[��6�e̲�����+3�J�_1&�sFs6L�Ii�c�u,��q�fu^���rw/�d;�e�qv�s&u*���Nwgu+�ah�(��Yz8S��]��hN��ڞ�<r�������o�J������% ]��;B5�D+T��҃a���si-s{W'ͭf=���81L��܎�-���R��FŹ��V)μr��F2�"�bJ�7s��{��QO�m*n�&d�t�`Jh����7�/L�R��l+!���?��nw:���z\�a�x h������/�	�9)��ٽ�:�ykw$68c��l��ZoBy6��P�>��3T�3���FG�4]`�5��O��iE��Y��·����2�V�Y�y�p�N�A�k����$8 �om�-|�r���6��:�=�����Af���蝤⹃��K-V�d^���J�tM�(yQ<:[��$V�M��
;Dd-:�:��/����m���/����c�;�����z�ߚ��ܙ ��4Pe��D������J�MI�CEO�#�"��������
*�!
2P�
 �&�� �:����B�!�-�4���K2�9)�1$TP%	�05aB�д%I�9RR�K�P�S�T!MQ�2V��ʆ�i�(hJuJ4R�R4̀�� ����*�ZF��*�Y�KKBP�)BR��!1�� QB��%�dRRTIAKDCDNJ�E,ELE-P�9TM4�ER�P��De��s��J�����r�s�EaM�a*�T�y�<�V)Ve�ĆJn�{�m���w�rR+q�e���q����WmN��8!��dpl�4_�6$V�&祥{�Υ3�ݩ*n��b=�&��^�����u8�5;[4�E��:��1O���Ob˓�k؎ߩr�Ag�V�_�����G�hO>�����OAi�v����]�[�l%��=�ת��P+�;9_e(J�U�ب�I��6���n��bݻA�_��;���f�O �{ʁRKʟl���V1�p�

:�͇�MQ�V'�eny���+ ɂ�z�N��#��c6?W��+KW�^�;E��o�!�����4��͘*�0[�
�V.�}��K&z�j��X�mT�y���W���Q�gs��}�>s����i|2��;T��w	~�s'����~����{�ޟz��td7t�,ǩS�_x��O��9���X�������ɥa�w�	�@���A��%Q�g<!�	���afW���=e�Py��T+W��A=�Z����{*-��)V�X�w�^G���rn����a�ٜޅy���Ff'(YD�n
;��u+~��n�v��j���[J&uʥ�d�q�O��Uw�.X������|����=�ayC��NJ��k_yi�Z�~�އ��;^�Z��YR�̋��{E��_�Cʏ�
�`���s�z�7=��Y~��}:���9]���~���7�W��DN��k<�����nY���I:�::��ԳjR�֛�^p��m����m第���}����rЦ��-�oq>���u���ˏb���d%/o�öE�5-�H:����;�^��+܎3���i�N��P�����W���������O2�S�8�������A7�ӳ �,�r�57P'X���bo^�֛��S��][�ne�7��^^�ܚ�S���6���fXy��צ>�Zg�wY��f�/����z%�s��v�	�zy!�`�X��}g�}�	~'�~u�x����(�-�e_�vA�������ߨ����UuyW��A�%��g�4�w.��jX�v�뾈�w<��֚�\�S1f�p�e9�����ˠn�&�����F������ {0>I��m��]72��3�����KC�oR���^�
8C�|�:�]HmD^n1Z$��A"��_Նc�ֲ݇�wΫ'/��U��~�x��uN_OOv	y®���vJl����� e�sP�V�Ŏ�躉K���}^���{E����M�SX��&��Oנg۾<��J��{w��}��^z�����w�]�0@�{p7�;:�ϢN�v��C���&>f46>BOI�ut�U���/���n���v{�o�'���U�v�����{ˬ]��j�i�Iy�b�N5��BoC�m�a�&��P���vX3�iy���s��L��Ԕ����j.�=�Q�0ۋz��tF�ˡ؉ԛ\���6oxE�!{s�R����9�/ �$����MV������'�ކ��+˽;o��Fz��y��>s�Y�Oz���o��Ǎ_��\��P���U4�Щ�?N��zW��ڝg�XE�D�aV��X�l.��f�P��yT��7��ׁ�HlM��/Z�xW2��}Tv$�0!aΫ"��}s�#P�N{:+��\BRe
/�nv)��d�Mf/��f�	���ɪ���z�PP���B��п�V%m�IB����i�Tn��3��/��jAߠ�|�V����7��F[��tB=Ũ��Ny�#��{ֽ����o~�OQ!k�Kj����{k+6z��=�Θn��;b�r�S=I�,G�:&~��/BU����7Мb�SS4+p�؏�`^�F�����y�?!�*7�M�:ח�)����F@S���n^�~~x�� �4��%i�G��c��5j<�Si��J���2�Z�P�B!뚼�C'��pC�#u��R����f��c�7�us:��B��i�٨L���I�=|��]ڷ���2)͏7U���P����
}糔���l_��jg\+
w�ك�K@y[�N�쓃c�����"��s}v{���>5�^�ly̹�!Ll-�%E���jm�?�k�*�6�o�;?o�z����7��fx>��:8ܯ��W"���� ��k2�"��ׇw5�rx���8�n=衡�t�-�S��W|C���:B^�ݒ��#IVˣC
�&�w�Z"��'�R��!ǋFM5��ж1�2�6��*�*�̨짘:s�:��2��o��9�8@g�΂�������E�=¡�fp�Kf��^zj35��&5c5�0�q�p��W{eJ̄�0��cW�KVآک�gj �e���v�Tj��}��%(�@=��ߵşs���}�^�]0վ	��/۫T�`��j�<v�Le��^�z���#�J�q�ʄ�U������]�D�ꍥ��\���.�`��}����W�&��A�6=�;4�Ken��0HV��e��S7�9���­�?V����ճ�9��'�׮�üc����Gv'��pX䎉�=&�,~���7�V��:�������}����UѬ�"�3���c��	�^0L�Q*r���j�^-�ԛ�DSok�̘O��E��wG�/����o6�rꮰ\�FU{�^�M�V�jkkP�J�=�`�p]������g�k_L�:��¼�^�y{��a���z�ӗI��jL�`�8x��A��`j�V�����&�Gg!|�� ��H�@�U�C��,��l��[Y��׼�m�N�k�;1��7�}}�D�-��{*l�ڬ9�|�S�3���p}�۱�d��(iUȎ�����Aۘ���3��~��¼OV3M蠦f���u�.+�-<Ӛ��-Vۅu�VNAI�U���ۋNR�w��x��̸;�NC�v����D,u�V���/v��y�opU�2��SsY/	'Zù��2Ľ�v`h	�X�~Ҷ�hʄ�W�x�ż�ۑ���߮E�G�v��}M����+"~�ns[�s����:{��o;�T�cx���C��B;�a�'�*�5!G�\�|^�й�u���'unn{�*V����y�/R�Œ\7�MBn1¯F:#P�DYP�˹u���캣���sW�r�����V��N���
i�)�U}��cو���i�sT�~����v��dk^�i���������W�������$[��Օx�oX��t��g�s��i�Eh���W��Wd�o���.\�Y���+���sm	����5������v83��Чt�J'�	�A�B��a��L(c�M�J�-Rqs�:�Aj���&�u�D�{�YS�4L냆��3�%u����r������(��x��C���/��n72��U��o
��)ꮩ�Jɬ�{����%�Cp�D=ʋQ������=�w�s Z�������W��e�<�����m��Oj,��_��Y��P��U�W����j�+����7�{���>��v���a�����J�w�z���Uv�m��9+ҏ���v-1�o�^��������;��`~ƕ��]g��u[a�WӃ�E��[Q'~�J�ɿ<ZxT&�_�mT	2h-�T^��G�i��_I�ݯ|7��ކ���R�PR~���<��y���zVa�̓�W��K��f����I����]����aS��R=���ьN��>�N'ª�l�f\����������[|Ѿ�^܁3���ќ��7�W�{���Q	�S�r�ZB́���V��{C�N�ݗ+uk{9���7�װ��ئ�~��*v�ʀu��.� �{�O˱5J9�I܇,��5�]��N��mNlֶ����ڠ<�Y/r.w�Y��>���(D�1���u�Ů���ZT�-U�GIZ	vP#�WN��=qu	��Z57d�x�e�s�����%׽#KP���L�,�|"��w���N��s��»��_'�u�6q�p��tF��t�M�݂���׫�[��G��[��EV>Y�&�K5:4���n=������o|�gD��Wx��d�y���qZ�kֻ�y��>\j���N����+������������OrA�8��S�+<Э؅�5:��z��%=J��	�:�r�<>�Ďbq��5�{G^c�n��z���{ʢn}Bw����.=v��1�b��i	��a��a��s{�O���o�����E^U�r�7YIl�1>�j�ԺuEz׫"���c�Yә���8������B����QXq�W��~x\��X��+-_�b�f�����^\B���W�4���ow��^�į.����3�>h_AQ}�(;��7��po������b��5Qt+7`�Q39�ϳlPS��2J��,��x�_\����6E?
�:��u�wٙD'���Tߵ벐�����I�;�]0����љ~�~����/��妖{�;����l�jG�L��f��bI��p�zn�6����S	�����: ����������oh��S��ྶ��ŝ׎�^ :PR��l����tJ��+8�R�]h>�wh�ګW"���:�A�p�<��z��ͷSD����St��=.�����9h�#�����آ�^���i���o�� U��#�
�������,3�&����P�+)h�q��m�J���y�����^�KG;� p��ؘ��$&��MN����f��I�p��b�y�u�B��g���3���y�8/X�P\�5��Y��jZ����z�ˏ4�(�nkh�;�ء�f��\FW���_o�_�,��h[������ ��а�b\�L`z��ʸ�t��a�{����{�F�)��<��N��M��}��s��**r��1�V���[p�Ú��=���~ ��̫=6�.��A�I�^�I����j14��S��nj�i�R���ý<���-�T�en��[��SФ���WfL�F���+Q�M^�#�������[/�Y�d&� ?�柽V$���ݿo�">Z0z�^R��9��3j������^�aլ:`��n�A���������ۓ[��m]9��lX�\��g��Q�&�4v<��'\���=�Z��I7q���������ew^�j��6��|�2�t)pws��_�ܺ��//U\�<�c������{WN�6�/o�n�3P�g�q�G�Ks�{O ����������>x�5&��({%�~�v����7�'/�|��61� ����(�V|о���\�ƥV�N+�����R��L�y~����k���ꮰg�s ��ͬ�q�8�k��5K_��>�.3S��z��T&�_Цۉа
*�/i7�F�m+��00�嫢�Rɨ)?k���;z=_'M�*��dO��)g������gPq�N4'y��7��|����-��Ȭ��0��2,���c���
~���b�X(,wzV��P�J�?c~��=�,g���v��6��S�/\�m�/�@����5�ug��s�z����.�&w�B4֫72��A\3l;�*P�G= ��m��c��{�L4ܲ60.�ݐE�!ù�d �R�r\���
UsP��;zWp+97}�V���!#�L㵑��E�/�Wj:Y1��$v';��*�nb���Î�JC��*����eX�m��a��3'�Mw�I%�sR`:�y>��J8iP;���U��h���3]�{�&�*-�p� ��ie���W_Y׽��u�V�N��U�s���]�lHVXb2)v�upd`pZ#x��M�\0,�U�e(pj�f�@���Lev��1�^m�Sm�k1��Ȏu-Jʎ^��v�X*�p>I3T�ǩV�˒,�Q9I�x�U��]ǰ<#0��{8v��8��_Q�k�կ7�,�P���;iW���C'��.����򼴓��*��=�]J�+];��ubp+��v��`�̧�O{vj��5]����z^��tS�.�TT���v�^�cj�[�T�V"�y$=F�)1`m�[M���y���^f�z�6 �.�դ�� Wؚ��0WIY˦kHQ��*�[��tv#Wh��ns��hu��v2�ζ���V_K�Y2}�wn�rQ���Qң�C��7��%���aw+{t3�$�w�>�*��)�l:��v����:��.��@7.T��L���5�MY\ ܺ��G��1Y{��ѩe�Ht<����yX��E���ngP��4�F� 6h��s={�S$�0�sؕ�,� ��i�|��w|1�{K+��g(�͍�t��m����[�A\1��}Z�;1���<5�t�2��dhw�W;j7*�{T}qe��y-{�Ef6]I�J���eVҗl����u�1�QA�$
��P)}��FU+���z���v_JOE��睦.y�����W�B�7�ފ��C��[Ko��nb�8C}nQ�2��j僵Ι`��֕%��v^C�\��J�s�ң��8>ief9��>{���F5�3;��-B� ��_>�0um��@�e�C܇�j���»-Աؔlz҆�T�X�Y�
��E��R&ɗ�s��8�X���D_V�U���J�
�q�bͻ?gW[�r%�W&o�9���h�6�Z��	B�(�����C���16��P�MVqx6E¥�U
7�����2�Aj�%��J��:
�	}pҌ����x�]֠�ܡ7�W�͓zp��A�x,*���c숁]ܖ�?Y�u	�w|�JtKڜ[��c���d�ӻ.bzhr�sJ�r�S�]��\9]�C�J2n.á޵�e9�N�Y�P^}Od�e���,,ԩ[YM�u;��Eu�\�QM�3V���٥�ոjs{گQ�&�Uuub����Q�x�ΥȽq��J�] ����I�&�&�Y7�#{.�	{w�t=�.�����l[�bŶ��M�B�Z���<ӊwm8Y:],k7�Zc,�����=X]�]�c+�՛�^fΜ'8FY][��^WV�K�l�����z���s�]��o�3HD�G0\���b����ĥ�J(j���H��������"��,��"
��)���2R�)(����F("��������*��3!�*�
30
� ���������h��J)�("J)���j��h�f)ij��Z���*����I(J
�����ZJJ���s��h���	��j�(i)���(�h�JR��
)��)��"��j���*
����J�i����*	����()*j���ZJ�����ZH�Z
)����i ��Z�j*	�!�"��������*�"*����+�o�o3?w���y�پ�����"א��X{�1X�ns�t:L��VV��k"Iڷɬ�1�П�M�uJ��cq���S�I�M�P�_B{F�5�&�m�;�+��tDơ�+'!^϶�|\�iF?>4{�:�N5�~Ŕ��jruyÚ���~�vm?\�#��z����8�h�B��՜��;�G?r�Y��K�͞(�Nj������6���4���Z�;���S�P%xz����k�S/���j\���ǁU.�3"�ݜ1wW(N����[.}�.�8{b��U�S�0^??wz�JZv2���{<4�����w��!��8~�Qf�{�v�E@�^V�.�m�DZep�}Q~���Y�c[)��$عm��e��^��cv���]��osM5���%�\Zħ��c'b������ۉ��#�ߺ!����yvMiߖh��/$G��G��eS�qIR�߮<�<���7�l\߼6�ˢ��*M���-&��\���6躔���'�p��L��3"��bÓd������)���h�m�����W
�����g����X�^o'0��p֬�m!�g}�˽�eq����U�]���b�6>�{$�x�xn�b7V"���Z�ΣL[���]��7�,�8C}L���"RVp�[ו��}�-MF����ez����I�U#A��2�����z��������v:g�ۏeB�>s*|�S�l���	��A�O'!��������JYm��N.>��ؗ�?x&��sH�;!m@�`�+oS��L4�{���c��K�:�-j��w�6¿��L)FcJ9@����cL}9;�Jx��]����m��x�z�ѭI�ŸU
� d�L��=^͝:w_{�m��h�����O�=�i�5��n1��Pin����N�:���/*u��1�س�m-����o>�=8�V�$o"ٛP�+t׫���^�ݞ ���>�O<>[U7���xe��+�m�[�pC7��z��s�4y}����5T���߲�.�É�z�,�78w!W��ڻ�؟[�:��:����̷���7�$۷JJ���gڽܼ+�dS��\G�t�P�=�y�H�ۨ��ݬ.��������� �5g��-U���+�iY/CM�&���[�u���I��i��Qu��SN��U+&�Q���+���v��@N�e�s�&��Q��m�w.=�I�DK��!�׎��T]-�1�YΜ�v��w��|/ܶ{��n<]��\�eэ[��HJ�d�x�+��z������R}z�����g�R�w���t8���y���__AQl�������N���F��MC�&h��-n3z��AO� �+稄���R���)z���[{B�o�]�7��_�<��z���w����l���r7z��<m���ۇ��Y��j�7����������[��Vw��*�߳f<��P���.cއ��G��]�2���{�����z�m�S�r�I#֌dy�_������}����ɸ��ץ*Y�*!&���6-���}K���Ffr6��v�_�����7�J�Mfk�Z�j�u7��~Ѵ.1���u�>JI������Y���<����-�m|NA�o��P�~���?�s�xI�����3e��rƑ�Jq��fw�[c�^][�5�r��+��Ѭ�m�Z)�bZ���uW<�2�̬I�6�Ɛ�B^Ŝ������
������+��A}viM�S�m�!���/�u%+p��դ��+�U�n�&�q��}�ȝCb�{���Ӿ��޽����{�W"qs��k�mդ����Ûn���U��Dc��iw�gc���b�o:@o�v�W�;g�絭>5ݞ�w���zh��x�up����\�[F��]���ުS��-�G��Y�j����fr�k��_)��u�Du�7~ܧ�~�I��'��=��El.cc�+V�׭�6�}�z-Md�5u��v�{�w7����J ��
�qϬ9��v�2�5q���lB��[S�ɪ��=��Y&���t����k=3ϵB�x���k�o��s�9�61z���v�~�2��g\��~z�4��Zx�-�W�]�+�xM��~]�%����{P\���T�P�yF8k�p��O.߽Hu��	V��b毰ng�%��}}C^�<G�)־2{q�}�f��y֩��r�[՛%#�B���wŎ��b>B�ˢ[3F�x�����G;o9
-�����o6w�i���{��rU7X���ѝT.������o�;eU�(R�s��՗Kp�p^�8�5R�y8����8�fcĖ�[بw\�(Ot;��<>L���[���~n�_T�P~k����k�_��<wϴ{Ϩw�t_B���N�����KL԰��^�d�B�{1���\�����
6g���S�wc�i8G�<����J�=����l4�ɐ�4�^;�Vi�Y�I��a�^�R���9@OT�9�2�>�Fq��',8ׯ�bv�ᥕ��Od���n1�W�C=v ��~5�sZ����mz.��G7.}�>�Ӑ�dϜ�+���xW'�Hw���c ZG�����w�m�U�6�o���׻�~��_v��%������!hy�ǈ������k����1�n�Bw��.߫�VR���zvg���W�~��|�����^�硸���qCݼ���ZZ8�������z�:��`u*GG�խל
q�'�	��Z������O)�H[S֖�5n�bOO6��|�Nb�(���3[��w�/�� �]�4Lk���0J�˩6�LؠN�!�1]�U��Ѽ�i��3ecg#l��U�{�:��-sX�;�er����P�Q�/c��v�6�r�K�JкBٙ\�����W�hn<�롊��h��NL\���v�ǃCO�H4�-��[�N�Ƿ�+�cv���7���XrY�Md�3L�V��+�~��E�*7�/[i��ח�^նU��a:��	�u{�N��̱Gܬƹ)s R)����^�xT�ƵL�8�F���h~�xG-go��]o��{�9�Y���|������z�sY�u%>���}��ǎ�Q���OR�b}��0��$}���;��Į3��^�c��Oc]�U�+W�'j�}��P��*q�h��o���Ϊ/W�����Mf-E��?b^���_Oz�%�P�f����~�Cz�5ƻ��kXR�����J^Z}���p�������+���;V�|V�f����S�p6䥳Q/}5��E��\F�ÿ�q�pƿ���1�T�@��*�Ԫ�jW
|"�����m���7��|'�(M���l���n�ۓǓ�S��X��]�����q���n�3��M��D���+6��1�^/J�[��>�K亲���w��&75K�{v�:�d���3_�2u�=�2�+^l�}9���$x�@#ǜw�I�qRB?��ҚY�Wi0lΫ��v�=l0h׉�̀��g ���ᏴY�����uY�o?D�=kO*�~��L\{�x���#ާ�^�,�.���x���2Ϧ�Z]�a�ټ����]{\H��ל����p�b����8Ƽ��S�eC�n��z���{˛����Kϭ'��SO���U�V�T~��zz�kaD:�ۆ�2���޻>�.�7 }_{+�$� 4}Y�}yz����{'m!r�e­�Z~�t�J�����/0�����l��b�y���($�]~���P�[�C��fn�(�gP��z1ϼ0�?}��A�<�Uu9�\V|��TB�v��'JR^�}������)�a���Bbf�ɷ����տ

~XIPC؅�=���[ݙU5�H���ۓ�Ii���8k/�8yQoV3M�
	}�g�tz��i����'v�AH���=�����^�W���{*-��2�@�����V�8�i�٠�������î*yh�%U��-,w����Ijxr2�s����
[ w�a�����Y���E7��5�p����^�R)Ƹt��Ms��Lk����P�۶��Ŏ;x�.����w�u\��0�'���mk(�"��{��L��;՛X��~�T���i{Q��o�-(w�ڞ`���D�f0/:݁QP��o�q��m�0K��rF�S�+�[���J�e�l[�[��L�B�&��d��rz���2�xJ�r��޼��}��9\�����fuA]i�v�5���kei���d�M�r��g�Ⱦ=���Zu���5\�q(L�pz��_��y/W�����b[q�O��1�e�u��ȓ��������;�����Sϻ+Z�]Z�Õ��O�Q���c�M �{�`�]콝}��4}O|�O��o�wg��R��4M��n� ���p��	����^���ܬ�s֗��3�\�����~�e�k��YK��y���5���Ïy�"e��p�<�����*積���H�?z�����c��Gs��0��,��y�������yQw�y����N�	~=��]M@�y�e2�F��wQ"!�<��\u�Y��^��]ҹY��˱RM×*v��-y����0=|�/;��������m���q�j��.��l�OR-�����Q��������@��U�(
ءu�duw	㚍�[�i]͆�[�m�{쿵⨏m���& 끊����/|sv��b�-S����Kޜ�j�5�M=���Y^�[�]U�r�c˳�.�} .(y��������5�yx�_��)4�ʶ�&Í�d��7y��h3_k1��ۢ�R�_���X��eG��{'.f���5y-k���mc�n��_f�$�nzs�?L��~�^�(���9
��ۡ��x^#j���iz�5/��cԁ��
��uޭó���y=��\�c�o��3�
�7�_At�"���k띻=��g��S��q>��Ϻ)4놵�BoC�f�wz&�;H�|��.��[w�pnͥ���xc�SW���Q�yY���NDkLKn<���$_ڃ�	%΀V��dk�HG���{�?-�&�ز�mZ��:+��nk����:�Z�%~6M[;M��v�Mߛ�H���h�����1o��]�;ᦖ�U�;����Y�s�@�'}���-�tOY���DbZ�Uو��ܴ�7�)���<�Dޡ�5�,=��t�勠״^�yBwll|Z�A+R�ql���i�~�o*�{V�o��ic���\�p����pˢ��L�<֜��9��Y��/�vaŲ���pn�絅�.nw�L{����� JE���y_��AƷ�z��=��7�]� ������[�yN,c��J~�o�{�i��w�lz_��������k�}\���;�c�k���"��t�U^*L���Lf�ؿ���v���TG��*)��N3ާ�l�8�	
~�\�m,���y6��^�Q_r>�zO(9Il�V�_q�'����I��4$��Rwre�ϩ*W���z��xX.ad8���I�w��ל�R�buS�g�s�|�+��2{u�"x*�?s)��rg����yQoG��n���6`�!&!-��R�qb���䭻P���qp�]��4�{*-��2�ȅ;�l����o��~0%�������\����ep�[�=sD�!Z��W�u�e�.��;)�O��ܦ�B[���	t=�]�h/�ǚ�#�7��@Χ˷!��3*0�����xF�"��l:�M.-�ua=a�[˳�B�ʇoF��U��tKt�a�	ԇk��1j倮�:�jDi۲� .�M�cޫ��Y�6�Tazp%C���&T�VT�k4Z��f����+&^�1-`�^��|,q��]�^�q];��穼�Pb���T��s&�6lX���ka>���v�>,@�N<]�ȝG7fĦ��_6c2��3��m��jO�j��G�*k2�/���|�6�p.7'k.Yc��t�ZY�g!�I;�>XZ��C�8���kK��,��nvR�y8����	 B�ۗ�C���c����Oxۢ���/i�����f叨ѕs0�I�.�˭�J��Ѽ0�j�v�&X�&j�[����A�t]�Z�]t��*�Յj��jQU�yf�4��ΰl�k�跌uн����]�hVQ�����7	tB�5<%���Ӛ���̝6lt��{U�ܣD��Bͫ9}�u�٩����؋]kM�׻1[�Uk"�\Bs���p��}X���Nj�l#@z�5W���n�f�ڇq�agM�T�N�57X���ї�ڱ�oV����u�:��S]kT_��K���x�Y{d���S8�u�T��|:���-i+N�F�`}5h�cNH��#����T�[�p>p%vܫ�\�/�)2j4��gz6�<���m;�c�ҶU����Q��L�fJT-jG��.-e�s\~K��Au�JK]9�*�tw�,sy�:�\cӭ�i�.ƥ�օ��م�܆h�d��0�M[�6��-�4��Irv���lb�#y��H���n��N��A�b5+|m��s.����(m"��Uf�[d�5g7m��L��d��w:;}N-�����[��t�@��&�GGv��8�Yb�u��<��c���84����A�@r�d�"N����T|�f���\յ{�Ħ�=2�\@�Mz�(d�,̫����2v�%Y,d�tz���Eso� �_v��l/Q|n�:��K{@L���	ҳ��.��t(�dy�����������G��N�U��6�&��q{���� e��6�{���N-����]��K�[�)Y��Jbh%�ژ�����ɺ����q֫��{:vP�2(�u�I`�jKw�:�kj��3���Mr�ƴ�B;��m�{�Yy�m!�pDsyzޫ�+B1N�G�nX�w�����{�o�·�A�'-֞慊�.lsd�� f
SD�I���{V�iӢA����9{��V�����Ӯ�)K�˦��c�r:�]��kl^q[�Y>^j��Wv-n�d>K��0�:��U]m��9�9��~�}s��y�g��b�)*��*%h
�
Z������"��"���)&��h��!��jb���������*������""�j
b()�

ih"P��*
i)� ��)�"�����rh��"�i
�
������"��(j�����I�i��i�(�j�����������������(���h��������
i*��(� ����*���)�
��
"bh(�)��j*���
�J��!��qj!���`�$�*�������
X� j���"�����b������������"fbf
�db����� �+�d��!��ˬ�O�5�:�2_�ϷGg��Ż�Zb����0�ēu;���Ť�97q���+i:u�N;Z5'����_'�ƀ׻����(wa�ǩ�9�B��|�+�F�����-��Q�m|r�k��~�)yi�%�Cz�m�a�&�[b��LGo�A��u�6���Y}-�m��E�{F�&�n<�uZ#ʲ����O��O�T���0�����g�s��_E�f뷩�0�I�b`4|��V�n��nz�J~?p���i�f=�ћY�s�s�	cN�yB�u��$׽��.�O�yU��7X�ȷ��,�m�d�	��=�"�o��+^���mWו��*_�58ƽh�D>�W�Ѻ�=���e��+�y�^�+��+ڳ��c^ɏj����>�}=|���]���~sV��R(���mOek�6V?�#�yz��<�i����;rV\s�'��F���Bm�˚��D�=����/Su�+���($����-��f��h���6(��ɕ�n|#��61��c����Ha;əT&���_N�ʭ��*�q�½t6��=��=U��*q�f������.���,vy�\���m�θ�홪<���HQ/#��`�[�"���7d��<q*(R�)f��֍3�*v���W�F}�o�x���V'nM��|�J�1*�7z�ΐ�X�:�U8��߯�=-?lB�j�а�+��JNT�����L�����ѵ'�ϥ��ǜ<���m����4/��d��#j��;��Cg���%�5^��cZ�_���uIE('-�Yy�������,�<�W�Vޅ���Yi(س�'�*����k#��q�5�]�����`?y5��~�),��I�l�Ɗ�f	yN��SN�j�M�o"�3(�У"�A��W;mw?!���܃^�f<j�+7a�רU�k
�eǝ�^��\7�P�hȨ�Zt�ֹI{�[\EB����gڷv�By�i�5ɉ��q��tF!�ZʈکY�f�����{0���T����YQ��js���n's��1�xo��[�J��yL����bi�����`��]P!8U���o��sn�d�L�z���_e�7�m�rZ"��3$;#�
Xr�YՕ�$�����U���S����Ɛ��Ү�k��E�p�F�hqG���V���zvz�N�f!�-�l���G�L�qݒ���;���su������՞�%����ޛ�CݩR�v��;:���[4���P��=����ծ������f�AF�벙U~�]�l�Wb������u�.�Ǣ�(����/��t/k^�2o[*w*��{u5���}���q�p�{#ίu
<�е�*F|ے�7k�S�o=�ۉ{�x��r|���^�EZ���^YQk��2���_���i�i��^նS�wo5�p�iQx�o�6�S��$,�L�N����8k�p��O,�oJ��5�د$�������|����o�~��[m�u����my����)ƷZY�}#��Fʼ�����eK�v`"��T��)ƀ��k�_����'�
��Rx�e98	��������:��b����v+�~2u	�\�}����z� L�nc�>�!�j�M띙�J��@^<�����ڋ�����A�'0;z\)�,�eH2�)O�iV��{Xq�^6����O���ٵr@�2��^D�^�&���hw3}WIS��-v6bTR��k]6�xJ���.��n/+��+W�\�m��������P԰�4+��<�|�M~��o\w��l�-�]�����3�8�j{ν�x�Jt���k��wڦ*�T�Y[�g�ܢ�\�Y��尿�*3Yu	�֘����+��DM�Z��{��ibZ��&�__�Ȋ�oy�|�M<jw�o/W��ې� �2��E;ay&s*�����3��m(<��o?D瞵�ǻ=&������-^yLfy�aGh�N�[赤V}����ջ��B�mn �z�פ���rt�a�ġJ���2�/[֚��^i�q ����8�_�nGh��ӈ��s�����r&�벥6���k6��|B��o��J�()|���L��Vw�%NA�{�.6�S�6.[x�o�	�Z��tυ�\�2�t�'�������;��($��hVIH=�7ޞ�<���g���g"�ն���T��ugiHk�%�p���.z�f�e���kXW]�ؗV�A�i��VD��˳�@s
pC�.-b�ۡ�:�����u�jי�Hu�*���1�$��\�o���n}RW#�֕M�j�\+2��*+Y�"���k���JP��wo>�\4��^��E0W{۾�����if��]4ޭˇ7��PR��*W�VdmY��������W�c}�v��k/�eD[��帐��`�Pt$f��V�}��_E���d��e g��S<�D��@g�[�{K������_�YWZ|7��7�$;^��vd3k�wQi ��{�������"����+&����^�w��º���~�n���NW�kW�oC�f�P��r��$����[��}�,��X��_\{h>�C�>_O4W�OW�L��'�ZbקF^=>כS�;�����'`���TTK��2U���Iv_��V��J�l�����5�u{y�����F�@u\Gu�{��Ш��H:x��aaӓ஺��\�<�ZR=_yL��������-6����}�������@uʞ���뙼��Q�����2���w�ڱ����tŴkw��ި(�~H^Y>��F�x��]��s7����K�r��&ڣ�0��%��1'���;��[s�(M���b>�-�2��m�X*��W9��=�R�"*{�wur�>��̭��q�˳�2%���ѱ��yG-!HF�,�x��`�P9�+}�\�g{e�m���K��1�O���ϣ��N�~��q�3�p�����a|��ػ����y�� ��(;�������k���r�p��]�#���ﻪ�﷯Q��/�g�Mӝ}JU�^%�G	���<��8pӠ9{0)c��I�\�p�GoJz;s}V�n��I�G�ep�ŕ:n,�)Y�~ ���WU#q���fG�u�X�E:��^Yfܥ9=���}��\9����u�B�T����9%q�*��E�n�\�5^�wbN��6��3С�Α�糮)�[��^���]9�I�X�C��C�ۂ��T���v��ǜ��>�~��7]�bo[��}�O�8�r�j?�k�{���8 j�������<��	��u��Q �<.#]��=҄��h�Վ����'߻�\uݳ��;��/7KW��w�=� n�f �$\A+����RW;`w���պN��V>��w9ҲN�V�=�u�����F�9A�b�um���؄�i��-�v���~Q%���*+㱞�tD�g�י/��Xs;)��尃eN���h&ÂB6����1.���k%�ac?f�~���x�1�,R�w�m����2��k�k.�|�e�u|Kˋ�������Ka��6��:#d���:l,C�V�yM��I��虄���wJ[ġ���U���8WTK�s=2���H�K��7E�ʽۅ�\�|��ܿ�w���]s�ez�F������H��k����c�`���	|Q���`��Dj�О��cwT^��]8n�Br��k�G\&�����&�wH���_�=�_)�T�K�Fs�;����eu
�V��دf��q��p��0��WQ�t�;o�,�i����(��V���y�~����\�}O����_B�ZN�6��˿��^�}��oK�UbT>�1�2z'�nd߷8�U!ء����҉�`��}=�b:�s�-� ��W����'�أ'B㒸�csF��?(f�.ϫ<�;q����]e�k�V��׆�k����r�^rf��w�w�����K�NG]F5>�|��e�b���sġ�/��S�(�Od����^��ў�z��P3'��]q7��=�}q�T��j����4�Q']R\?7%v�J���ox�U�w�詜ً�J�鿱�Xq�<
���|_u���^FᕆY��Yے�焗_�Z��oU��%���PM��V�M@�%���C��ۍWa�t9��B������zw�����Tl	��>7�;�Z|��Q����0>�}�n/u�4^Z3�>�oF�W�AS1v�5Bs���-p��{�.ţ��i��՜i��b<:��ڂ��_T�5`���gk���蒥���FR��������c3�3����8�Ek�� WyB��7VS�c"����%Q�~"E|z[S�z�h�[���y\ʭ�F�4�{k�����c8Y��H6���='�|ȁ���8��|J�
a���B�~Ϫ5mL���z���)�m��Z9�Ԇ�~�7����2\� �q"��nz{�}�`*&�6g�חf�RC=[/r�Ѷ|�Lf�I=9������X}=W�o�s$�P�Z#I���A��T�1��ӽ���>g{L�7Ѩ��u���O&��P`�!Qs�μL��]�����3=�xTK��	ex�F*zo�]R:�+�1p���7�={�Q�X�lkΞZ'6,�-��K�̓�2���%��DKYx=��׾ͦ6᫿=	�܇�#�wg��΁):����������-<��g�[V��U�b��o�l9�?s�q�r�e_�'�GNu���v�>~g����o�u@p��1�vй����c�e�^����^�p��~�+��z��d{5�gWCl|��%.߼��˯�j�N
��\�Bk/A���ؾ�C�W�0�y�^����x�Vy'��ʔﲲA-_V�jt�h��Ǳwa��ҋ�[� ڼ_tY�I+g�wN�o�]�ޫ�����Ը�U��#o3M���^޺=�>��=�UWa>N�.s���'{}z5�}'����.e��A���Fx���b�C6�g�14ȓ~%�w�W�sO��]8���q�Ы�j#ǽ3��t�9�Y�퐆c7��c�PN�r��]A)��2�W��i����Oq��\f���1���W��Q"����~�[	f����pg������#q��2�L��:`����ﻩ�U���g�OnV
�>�Q��=�WA���K�<vΒv�3�T���F��S����7���:�m����=���bc���wQm���|�ԃ�%���$�3�UAl�W%/�Lٹ�rSO�����/�;5��_��q�ݴC��RG�;��w��u9 j�����u��ݍ�r���fׯݱ�:��>����\M�u�|\��ӟ>��o��F\uճV�Af��w����� ���O��X����#<��5H/|뭳=�m��=9�����\u��nyc��r��~��A5��� ��_i>SC�Nw�y�񪑛����Tx���ڟvy�A�dU���q1��R"��L�ܠ&��	c��n�8��(=��z�X:=ֺ����TV���_3S�H$b���|i�Vr�L��҄���w�V�I/��iJ�cD:Y��*k8��v�%S��l���J�뇷��o�R�kr�\�mN�o0���9��b��P�����~������j�[Lu�kw#���w#���t'L�g��5~���J������TC��K'k�d=7��TW�����9W�zfk��&;�7����[V�r�WF㳨��O0ddoz���'h��7�k`4��J�#�N��2�I��ȩu#�����ܿ\?|�]��{�Q�ˮ�}��h��}{<
5���F�7(����N�}4�0�{tR�2�n�I���|n=��8�=��V�y�+��q���7�3>7>%�}u4?���k���DΎ�87*}G�U���`(�r�p���w��ez;���[B��'�i��ڌ�m��S+q���t2���p���f�ho��/Da��H���5�����л��%�KX}�u��?J�L�_Y�R�0�j ��;��n6� �l���ҷVG�����=���b�wu\Gc��;�w��?}�hp�C�Z\�݈��N����U�(�"巔5z.�ɝ�/��(�y� ��v��k����^z3�)�G[��u�A��]D9�Iڙ`/��X�p�_�@��w�9�[�xh�Y�
�CeS��{P|����Ŏ�`�\�+gȫh,�s�	�.�`�v�
>�o�xy]o��~^� 2�F�>��{x\ݡkPx���R�7�2X���1J��U>(��b�k�Y���B�k�e��w�cS���iƔ��,�0��{(t�]y���WvũX�\���z�cmf��!�V�3���Е��	ͭ��m�o�CX�@��hPwt^��
M�W�#c���	��![ei'>êud�rvd�'jf\:v�sI��eJ����J�����Y���O��>{�U��7)�m`���j��"�X9�&2tXR�s�⦠�s�ß�;p`����֥rBT�Z�/�IY{k��X�^7LWP��u0�\0���V&i�
�_2��k�	w�M� ���f`��W]p^�'l�,t�B }՝��ڢ��>U��"V^��5pLޜdh�Lf���ё�ۀ}�Ui-�0L�І9r��W���Avi���:�A�K�s�a�R�B뎅h(���ﬦI�757:gu�����S�n[H}�ʺ�A-�Y�2E ��:mT�[�W\��n��c�a��:�h�LU�$_&�ہܲ���t=9���_-m_rYEU�L����w���APP�;{��*ΖE����ī{;�g�r�u��nX�[��}z��u]������0�vW�F/t-����ps�jK!kف��zR[�]m.��eBy-��ZI��]B�����줣�ݲF�w�9�]�Jx[E_UņRCo��7��׉�\��-���=}�'u�'���&Zʆ���[��ɺ�����cn��6
��z�b�o�3���4��ίO)V.�Ʊk�F�3R��-	k"�=�j�;�Pٖ�Z�\�B5v�p����P�]X�֪S�K�R�ӗ9�ưIx/rm	\ơ�*)a�k��{9ە�4��I[�w��V��M2h�F��{�\`��9��gPzjig���H!΅e�z���lXB��9}���fL�,�!�v�y�Ϣ!�h���)	l6�O�YSq_u[�{�W.@?�����4�9g�^
�@ }G.�-U�����w�^_2o��Q#�J�n\%�VK��S��J���ZDd2wFd��W=ޫ��R9ܞ6�>]�:�S��S�'q[���vsFi���4���X�@����ɍ@��
eu���;6�1׀���}'ֱ[[tn7�lV�t㎀&��AV�r�=�����'3�Ž>���� �Ήs��+���]Io5t��M��.�fЮx�d��u�WX��ԥ.�#��Z�ǈVx	��D^#t����m̀�������z���ˢ� ��=����rU�R�Z��!i\�<�i����������룦��4Vd�J𥛬�v�v�Et���EƄ�N0�E���,�:�n�{a�|�2{�q�yO/T���a͉��ݳ�o�;z�k���g�u�T4��PSAHPPPSU	T�LKDS%QQ%%R4QLEB�QMDTEE@PL��$AU5$�EIMD�U-QL�Q~�f�h��b��"��h(����H�*�b�*f**��a���J�")��)�*e���i���*������jjfb����)*j�b�""b�(��*�����b�(�����(�*j*����&��"��jb�	("����&J�"���f(�b�"*�����*���*�
�)��j�����X��h���*�("	(� � �&��jh�� ����h�"������d�"���&���
����N3��y�Y��̫
Ō�7]HO-2�8���G���0D�1pǨVG	��u���4�q�2�ʸz�(�spΡ;x?������-}�w?�X��n�O"x�.#:C;�UM{�x��ϳ�eҗ����U{{��8��$)�j�:/��t����	��C�~Oz�<����>�ǌ�Ȗ�����X���{�zJ4���:{$i+���,+�ֆ��tÈ=�ll�_v������>X��Q�{��pt�ԭ�M�%��D��1?J��7^��@U���0-dt�Ҽ�N�7�n_n����J�%����_t�]Q.�L�Cf��1/k��Qzr�=alW�{���.��3����*6㚾��ҁ�Ƹ���
�T��R��	|F���}Z�c�Q]kL��.�R^�Q�+}���z!�p�WF㻨S��W�����ݕ���-[��,���V��im�s�o>u/�[|+ћON����	��1��o�= ���,�y�<������������'c��X��
�i;�,s�r�Ç�����>��/�˝;���]ǜ�ݣԣMt�|��X��n ��$�]���x����vM`��+��zn���g�/duP�1W�	l�yx,aQ�z�e��Iy���X�m=�����z`ƭQ��U�v�N����Lh�EL͡[1��8�����e@�q�#_i5b��̉��c�iK�A�wCPPD�}�i����v�WonR⚙Ե��y̶q�S{���.�e{������.2�R=p���pf�A�P���V�Ծ%X��΁7
�z�&z'F{T:���̢9WR�Q�O���e�x�$��sġ�2�h��+Z�7��;���yE?g�yrE����g�;����r�����q^��q����1��b/d��w���|5F���g��H΁2�����V��q��?}�����<^Ǹ�R�y�^E�U���[<e��&t�� ��,	�b�U!q�u(�SBs�}|4{z:��gPgm����7 D���I<�T�j�=^���x����X
D�=-����Q=tߴH��{�w�k���:~D�y�`V�j��a^�@��ϯ�:,�9���0�L�IqW�CGۖJ�k�Q��ח�����J}��GNW#����o��FuU1X�K�D ��� �:	�4�LnRy�>Q��M�f��v�Q��[g��4������^�s�|f�s$���zFP���c����"x���V���Ӄ=g��ƍF�&�����Otϸ���`i�/��{�O�LʵB�^O��n�V��M �GB��"ξ�U8(��^�It��C��5t+[x�M&���hJ�W�&�ia�si,wI/]����왝E�7���-�k�:���.8�y��z�qx��6������:B2��T�I�ͧPP_����(��.���n:�!�\d��d��P̎ˀ�¾�:������KË�Gt>Wrb�>�F�z��WF|�z�����9�Ҥ�Tw���d�N���n��W��^e��5��cZ��Ƨ�r6�����ɽ�b>�X��T�p��G@9��(toeH:x��=0���W�uf�\�<�U�ѝ�t&��������&�yMo`���7�C�~���w��6�s���̨s��t�Q�o�S���J��U���|zO3q�W��꫰�'\9�wQ;��ѿ?O���g�×�L�H��n|�^��V��3?K_��݀����p_dˁ�ʣ�D�\Y.�3�;�����7���;}w
3݉W�ݍ����eW�e���G ���|KV|�t��>���;�v�3S�&��
>���s��j��a��T�,���P3����F��\i����Lk�3�ی,�nz���8swb{|s���[�W��k*Y���ό��
�=2����S��߬C�4׻�Ÿ��\�AR��������{�y�:[��:� �.K4ΒP0�\U��e5k��ˡGƪ�=��qW[/`��!/�K�a�R���sYW�G;Q���d~�ge塦�XX=�q
�8;����H+kD�救:� ��\G�k���c�:-H��ٵ�\������+6u�AWv��a!&1���	��1�o<�<�]#5��Sic�6��'�}쨞�]}�ˤs���De�]��K� RC�g2j;�A����<���ۇ�a��|�&���H����V��x��u��ul�$qt\��éź��+��g� z1΃�y�=�e��J��[f<{6�8zs	}����o�h�y�9Y�ǹ��,�#���"d�SBY�>؄g��ƮF�ͫ���Tx���#��N�oi��8����|:� R����e���L��;�/k��k�Y�����GY�
f��W��е�Y�5��t���q/ç���w�]�4��� �zG\Ǣ^�a��+n�b=?y��¯�sIn�e}�l{���y�Wu00�fhf��A�SĪ��鳓��`r��m��o0N']Vz:�H�zor�p��]��@u��Z�.��#ޙ��l�(�w���z2���X�@r�\Ez�˅t��9��q�qމs]�<�Eo���%_~��v{�w��~��U+ʱ#/#s]uњ=���P��d�w�O��4���}i�Y�^��K���]c(����,{mD�	�K��q������S2*2,��+�D��}�� A
��j�mW]ބ�[R�e 	uw �+l���Vfূd�)ѻ�ב�a�݂|y�'%t���5�.��İ�Տ��	h�5*�A�F^�OB`wO�\�$e�xgh`�V5�H�M��Ut��F����T�E��;�Ȱ��5��4�^�4����!��?��[d]46��o��S�e�Jý�H\bʝ7g�J���;P���om���LU{zD��=�U�����������ޮ�v��Zz�m��'MDI\hʨ}��6����%>V6��z+�`7����oWa�#����z����Z��.��$�p4q�r/+�:>�{�t
UqS/g������MՉ�����I���:C;~�p���^��љ:���.��Z�k��; �t(�({����Wu!7]h`�{����'��k�=~޼��gV��~��WG]�0�=%���5Q��-�pJ�>�R¸�ֆ�GW;c>�$�nL
��g���c&c���պMǟ\7�u���2Y�D@j����+�h�Qz{<CwG�y����kc=���^WKo����U��=ԉ�q�&�uh��P�zeX2#I���F�=�k�Mv��wݶ�Uu����	i�������p� g � �T��SngE��|Z�K2zH���6w��-�c��k���ݴ��5 ᡲJ�=����eB+;fH�.^�NG�i$���B��Qp�y:�y2Zؗ*�Y��M8��q�ɶ�Tr�|Ӊ݊�[ם�w)�\��{Jf��h�-s;�{%�ɭw�!砑��V�ʺ���Z*⧑�7���7��ˎ�>wrnJ�h�wPވ�e��zd�-n���غ}N'wn���Ћ���Co�|:�V��|+ћOMƻ���}v�=螢�����3T�v��כ�2�k��#��G��d��za�X���֓�ͦ:�r�Ç��^��bԪ�p��w���;��Z������1�붬��7�0�a��W���A�X-� ���Kr���z�rS���U�zWoK�47J�{)��H�<O��a���P�U�zpv�篇�u}����)�nʝ�m��uh˕�B���'#��Z�>t��B�/�S�&��u���M�4o�NS\���K�Iތ��i��ʁ��6g�<<N�r���E��q^��\f�o��S�:6�X�������K��I�ho|&XW�L�1q��sx��=<
����>��n�W^��{��*�ʝ:uT�a�+�w�A�3�O��,]J�/n�Ͼ����F>�=�Le^�� �nq��NG(��h�}��-�ǫ�c����X�J���H[S��Q=tߴH��7��޺W���}��X;]�|�H�|�<���,�'�b�D�*��vMhgޗ.��]����U�:�˸�;�Ք�#��gP[���i!P]l��B���wO�W���bP����{�ݩX�{`cG6m�k��Zn�[#����u���eoH���}}qށ�<k�DU�p'��i6J�X���ͪs3��s�O��F��gk����/!����Ԇ�q��#:���Ir� 55����kR}u
�3�om����g|��E扌m��Gi�/�u���_���,zC{ZWMw�^�{W�m�[=�RD�Kt�]Oi��ⱣQ����p�yǉ�'�XO��7�e������m�ل��r�f���u�xTK��B�+�a��OM����ܘ��\���8�Vwռx�Y��7�c\�K�TdS��$�Ȳv<a�	��k/S��K6�֪�0�v�@����N�Z]WH�*Sq�<���C7����U@���9��Va�W/O+S�kڊ��5r�qi�^��A����.��q�2��c�e�Mw2-d�r��|Fdø��*̥qX.�a�ѫ��5>�p���\o�j�zUv���㵐��K�����	�d������Ј,��
ngǠ����g�W�+� �,��^���/.�F���\��(.^���?!a�;Z-ޣ�[
�3�`_�y=A��|�wEW���"���k���v�d�;�Ѳ,�°0���{*c��JZt�ԑ�8KWG��K����r�c�<r-�}&����ZW>0乸)��씳.�.ڗ�;��~i,��9>K��r\�\��_d�^|�O����;�g<�d�O
�z[�s�W�-t>�F/T鸲�H/�Ζ.�y��A��49�g_:�^�
�����7���]w�OP��uw��;}ב������:��ƾ2������m�p���w����J�R`����p��=��B���gA�|�h�ۇ��i�R(�r�J�0�I�P�9:f�ye���o�3=��w��C��N���ۉ-�x�#��}�D=>�${���]9 j�BW�0�(4mo�tM�U�@^��zyd�h����H����"H÷��#/����B�X��Mf����ۜA�ѐF�$����Cބe�q�R�뭳=�m��Ӏg�]d�`�Y�ݓ����������$��H��(c ��B.Y�+O�_kB�y����F'a^���Ӄ�v=7Şs>�{���\���'`�]�	�/g��k�J!m1�=�Q;U9peǥ�iygR���Ѽ��[�\OzO�����r)d�!�=��^�aG����pЌ�k6~o]��.��o�����7Kn�o���f"�mm2�#����xk��n��]��&���>�?^7�]5���� =�#������B.[��!���;�-n>�Er�Wx��˜�,��Z9�w 9M�1a�����aQ�NYRܭقX���b�f�Hj��7IT,=	<��utm�PW�|��sC/{� �)�T�;�D�V}t��3}�:��8��ɉ��tg�/���]��@u�ˮ����ţ�w��'��H�J\i���l��?*:���q^�2�WOIӚ_�WY������/#��J�=���I�$�Z�ə���H}�A�u�,O�����[�~;�CiW�s�-�{����]�Lͤ�$�\N�]z4�(��7�GuX��ѽz�e\��'2��?P�E�����N���� �9'��9نLw��vç�꫞�#�j�p9���u����H^,��qx���g�v����H�i��io#R��������l����_��Pн��C���:冻��ᾇ^�.!�T����N����gsFZ9S�����8R��9P�����vgH���g\>S�\7νh?|��v�����M�lO_�b��I�h�$�/]K7MՉ�밨�'�ӜC8������I��=4&}����U�� ����k�y�C��O�������C�޶��oò�_����`��;i�a�7ۻ�i�<�8�	r��$�X�(��{$ujv�پ؛��ek/I�j��p��Z*�/j\�mE/��zл�e�����(5˄=��vZ�m#��MF��\Uأ4I�2��.v�P�96�j�J�oG^�e��q��N��� ���ƃ�w|aŒ�( j�2L���+���K
�Z9C�AQ�]=}U���K�c�V�07δgwV�7�냦믮&���" 5P'I��][F����yx:��9���n�>+�s�ѷ�G�B|��D�c�ߟuh�_\K'�V@26vH�\�)�Bj�'sw�[���r�v�񶘨�m_Q��p� g � �T���ۙў�r�^�P�o1�<g��
�j�U�R��7e�]��|���<��Ѿ�7�̏T�i��G_��m�/f�5�s'�svh�P�|:�V�[��^ͧ�]]C؄���ފ�7��񝨟�5���U�F{��זo�_���i�U@��W+��Âպ�wٴ�\n]�p��<�ώ���g#����=�<�^��%��c�6FW~���x֭��S�6�`��hk��E�|ڙ��� t>�|=�׀��Δ�XH�{)��H�<O��f��0����[��nI��joyǗ&x��	q��MY��wIκ�j}��H/.�B��9'n�C*"=ｿ��dᆻ��8k��\�mk�-輍K��l�n��[!ю����w�#ZF�.��⷇:0��X����W%C4�*e�}��<�΍A\���pj�1E�Зu���ɢ+6�k�pm�����d���e�o
��'b���ƳT�o1󡊍;6��z[�t�㶉���B�3(��.�͇Qi������h���Ll:&UGH������)c'l��l]O5M��%`��ڵ�+yR��FU��y��rck^^�\s\n�`i�|@��[�7m�Zk3{6�Q����of� ��ki^9]���yQf%RbP[�G[�3w�u�����)��ձ�"�Dp�w-ZP�+�b:�F�mN�ɚ�Z Ăڀ/-��?*�{���_<H��җ�h7N�*�ҝ�V>�4�aCi'�V�ԣ�(Ʋ.h����'hܕ�]�^����͋��Q5hYJ�� m[[���$(�Q���o��p��.��b:�9V	�K��U�Rl��k�۪�Kh��ǣ��u�y�\Q�ҵ����Z�s�BY{�K�H��Vœ(��9U�G-=�)�|s�A��ʒ^-v�+C���MQe�l�T�u�'5Žs�f����Fϑ��T)���Y�fej�]s��Uo &v����9���t�����]� ��MЎ+(�n���Hvp�f�I�R�.�f�j!:TW��!+�]r�)�Ɗ�Q���ڹ�vQ�R���P�ӥ���z�u����U	y.��s�X%�fPx�����֊����i�T��8tH}f���x#��gbiN˵��)ܳ��@{rP��_rmS՜0^�J��2�5��-��'����;��E�FT��r���$�'1�����E��:�ih�*������J��R��H[p�P��Xv���qt�/A�`<��u�So�+/�r���he��*r�7:�r[k�K��V�m�d�;Ṫ)}>�&XJ*X�T{��) ����g��c�H�W��6��RS8Í�k@�T���;(�K6�۱7#���[��(��N9�f2@���M��0�5lF�q�2Nb�.�g5.kZD6�m�%#?��;���x���]Ų�;��3�N�3u��2Z���99��9.����\�u��r�Xt��U� �R�Ϗ0c�f�i������I�ѳ;�^:C�!�Q�5����Cbjq�/z��-c��Վte�wϩ�����l�eK�klm��u��+-c�$ҫ"�B���;3�4��
r����黥��Yt���Xtu��6�[���	ˮU�\S��cq�յN�JF�	��&E���r��-]����$W+�.��4'6���p�y^���%�譌��iKn����*�K-drP�9(e�̾������VSY�4����`����45c��Jl Ѯ੉�u��_b,�T���E�H���7�lS
[���( >����"�"b( *�(**���j��(j�f����&�b�"	�����&����
��"��������"����*""j���(��)���Xa5LR�QT�Q�55D�QAUSSFa�SQ0D�A�E5DUMUA�$DD�QPAUMIAU1%UTQ5�M%ESIL�$IQPUU0�EQ4�R�ATU5IQTTPQDDTT�2����E!E4DQDUUAQPA5TU�TLUQ$QRSRD�Y@QDI0�
�B��LG��=|i�6ɀl&�j<����pd�/B�J��@M�'�	��gv�ǼKԱK���)?�����Y�w�e��m�����ν)�n6�6t����&�|{r�㸿G���7л|�^W�1�7���;��9���{$�S<@���*g���Z�7��?}�����<^D>������k����".du��:iEq���{J�Y�� �,�b�U!�S��~�n�M���T�5p�a�z�J�D��b�z��wQgn;��o��q����YcI(��"������Q=G�ʤ�]k�"�w�J����$�^�+�Yʎ��ԁ�>���@��5�"��0�L�I����teg.~���ïM��T4o���\ur����w!�!�߻�����ثs%�B �\o���(D�gT�ȞJg����`-=hLv��
�o���Ni�9�NV>��.'����N6��a7�tUa�3����ڪ�I��RV�D�J�B��>�2��4j55]E|�y��3�'�꡺�X���	d���5���r�d��¢\�]+\b���WT�����++�~��Iɜ[���KӋ��\l�=ܨ��ѧ��>�Y;P=0�Y�}-e��[��^�6��Y� �}�o6bU�i�;�?z?	��g��I)nf�W���n�#�hN��MV�w.f7ZO 1�'-�����Oy��/��
�h���Z�sA\��mCw�]���en�}�RP�ړt;�nJpJ��STe��>0�u������6��J�V���N)Ԕ��Ϯ�_ݝC�o�� ��.��� ���za��
z}��~���������+��|��h�m��y����}C��eX����ީ��NT@>�Z:G�k�~�p�S:�"�n�5=���ж_�m���Uv���<�bqGn{E���O�Ó��~
��f�kAJf���L�86�U��	\J7�p*<��w�\����\�+���$�Sy���&�F{��{<z0ߥ`��9)/a-��_����/�aw��'O�iy���w�5x�74���\f�;�b�eN��Ĥ �c~��Gi�e�49����9�o��f�s����v1��=�O��]!��ב����f�����0����T�Dr��K�Uk{�s�烳��w�!�o~��y�8��#�����|�ԃ���|ΒUG�a���/��\\b�[�\�j�s�H;�:!��'��{q7���s�}�C�q�TFwUp� �/F�^��"'b��u�N�zV%� �OD�`c��2�eXh��+����H����>}#����j�m�-��mV��˸� Ġ�V��Ge��Z�FJ[���j���6����\�lbG�ݱf4#���WB�E�qbiG7��+�/Y[r��]����9�dֱ*չ�g�����,�-D��O-n)V�Lڝ��u���Qتn��+���ZM����i4a��i��@�փ�B�!h�cT�s�ف��H�OgD�Β���u�}VOD>냖���2Y�RCQ�G��SB����#<��\���y���3����=��*o�ج�q������2�1>F\��3������Qk&�_z�ZY����&`m�͛m�K3��}�nC�]ȿ�u���O����TC�N�2��ި�ߪ�?���TN��Z�'uF���DQ�r��p��$��z;�]��P]��a��޺�r�)N{M���q��&���2�����=O�]:�7�+O#��/r�p���>{�Q�ˮ����9��W�6����U�r�OeL�9@��aF�^�j��:}��߶��{�s]���
ɬb�k��t�M���y��l������Nu>��J���!m0+=����g�c%x�c�쇹�ݠ��W���n�7�Q���T�E��pf��,]zk� r�z�ULuЬynĺ�ΐ9�\J���s讧��+��ﻶ��YS���)Y�~ ��At����AկS^�c�����$�$J��p���A��9�sg."��y��ݗ�,�[��lh���r�Ж�Z�v�J���RK�hR���j˽Dj�g,���i'a�۶[�FYT�A1����y;1��7�_�Om����U��i��9[rE�j�A�ϯ�ޣ�Ӈ�~3n�z4�ч�ȿ�����p������u�6E��<n�/�t|�"�����fS<p��v�.�����7w�z��:G�θ|��n�o�׭�p�ȹ��g�}��2ֲNs�	.��`H�P�*e����f⛫��a_r�������nLl9����^����+�ѫ��q~�����,	�)@����z�����HM�WZ3W�+-�n��N^m=�'�Q��=��8v���.:�هK9��2O���E�J�>�X^�xg���{��mz�߳}�xwV�`w���պM���鿫��&�,� 5�'I��][F�||�U��nL�1>ט��)��k��j�x��=�ԉ�q�M��㯮&��L��Ce�����g��V�K#�{)Q���r�v���1Q��j���wu {�k����9�
����kuxGJM��l�����n�8e��p
����;�����ɷ���7�wP�tF�ݬ�J��2}�Z��Rz��Ozd��c����Xہ���R���{\+�/�w������1F^�;:2hLn	���z��;F\4�p^2���H�F���ؓl�h#G�ϰ.8����[)ᩗ/axG}�v7�~s�f]������}�dt��Bk�ieFH3rJ�+j�����v�S��^�9@�<���w�:"H cnfi�q�q'+����$����$s�li��C�zyla�P����� ����7{�ޞ%P��W+��|3�n���f�׫���Y�|/=�g�搞CwR^�c���X��^1��>7���qat�+��UE� ��uU��N���9w��րy��zW^�]\�^G:���oe!�s"���̳0�n��'Hm[�A�^O��RCfw�:)�i�5<�^\ ��jȵ]K�OT�=�� ��-�9'e���UZ2Y�ʮ�y{-��N�+Ơ�TmҪF�6�s:O@~<JE2�;��W+��K)��L�kb�@�毰tb�I�q{$�%���gC�yLdm����X~�4�p7�G�ñ�^r��xw����b�Չ��[�[���m��Y�$ό�$E��T����S�E�V$�Uƹ�vK̟G�xyUӱc��:�g�;h���>w����c��Y�gI*��& ���mNMWA���`�s�j����y8�uf{D����Wes+#�;q�@�}}qށ�<k�DUa����� V�NUp�ع����H�$�\)���{��'�yDt��}:0��2��ثs%�ɂ7���纳%��uŀ�-��k9�R�*lw��4']Z�mjV�Hܦ����:������;fAq,��I�Ϊ0��}��]̻�2a�v�Ԭ��T�wv�mq��;���h�a��J�v�c|�S��L"ԓ��}ř��tϊ�g��ɫ廽� e��G<�@=���#PѸz�F����}zsOq��;�� ��\떟gO!KT�K�^�zg��X�U'���"e�!WR���i���Q��j���Ȟ#����ˍ��uIy=�W��d�D+�; �]��U�Q.w���Xj�S�j�ٱ�۶�^���R�j17�F:�Y�p�z�9��=FI_"���{	�����z2�v�����*��w(��	If�
��~{��w!�H�������b�{*A���U|=0���aWP~&bE��(��LN�����?�K5_ں�5��ӏ�q��V:�}������%���^�n���V���X�VBS�+�ѿ�K�p���߶���C���|�p\�LN�z�{�!�<}q�L�&�����*��5�僇.&W����Xl�ģ~�p*<��w��><Nu�2�^�7֗w�=��nV�^���7o�8-t�9q2Ǫ΅u=G�t9N�J0��W��)�ڮ�T[��m�6R�ge��f��Y��YS���)\c��bI�s�A�j�z�n�m
�?z��_��E	�4�]xe�Z��y.��;e˾l�$GL�z��NVZ��MV5��i�+A`�����V��1��0���b"Uwf����7LHx�w��-5��E�����'d� k0U���On���� ��)'#���mL���
]9���]���u��ב�k*Y�����0�����z1�A���^��vJ�g��V��z�?i���g;d�����i�:� �g�J絢����Ǳ��z�>H�\�ڨ���uQ<\S{q%����9������=ʈ����yC̙�^"m�����ĝ�٨�������l��eXh�)��I���=�aؠ'raL�"��dw�mV��L��i�25
Ҫ"d0���yh��� ���1�=�{NVF+������c�_���0���\���4.�f�IF���M	gx��Lx�x�@��+}���nE�϶�c�{��>�q/�:� W���M#.N�	�]bw�+藵�i�0c�5�[s|N_�{���RS�^������G�]ȿ�u���<w�����N�!�k�ɪ���a͒���B�]�GN��>�<�U���7	v_w:�/:@�]��i�42�{� ��}B;\WR�J����m-]�\���u՘r�i�+T�7�~�~���|���}�\+S���Ȗ	W��.Z.��bWp�z�k %R�4婘��hΛ�K�d�yr��v����˱�5N#O���ɏ�%ۣ6M�j37{���WU�]L��Wd(-T_�H��7݊��hV����˙݌�C*�t�Gi(L���Q�H��C$�{������ޙ�,t�x(Á�z�e�����l�7�qޗ5�`+��_�B��W�4UW����ܝ�J��y�㏙��99L��߭���w���']7�u�`���K���*k��{5)����U��#�����7"���ONc�x�P�����֬�{{�J��]iܪ|�.���jbp�u�A\���O���3�v���M&F��/���χ�wo�V��c��&w���*�7
��D���F�"�{/�w;�ßU!��Zz�nR�7x��w�;Vv�Wi&�I�4g��FZ7[.f�����oWa�gH������#���Ϫ�M'�gӹ�p��5oFp6N�B��'��Sje����f麱7���}�O�������zsl��J�BǸQ��N�o�<��p@�@�<ܡ�^�|g�P�мq��;�;)j�w�{9�,<�KOG)8v��w\��f���( j� t�H��O��3ڏ���v#�W�^��WO��h�Cݶ4y�;cǳm�ϻ�t����M�W_\K�����I������N�`�����F�1��hi`|0�ϭm_�+pH#2��6�T�B���k_W9˩Ux(U��Ǖ�JlM��v�cv���J��J�n��`]�$�[�� ����8���'���:��]zc�o��4�s]�A2���y�7nJJ�G��_n�y*��E)��?���G��7oW��q�==H�����>��.:��j�L��n룧&ѽW�s�˅��F�:%�To�<=5���lTm����wu {�k�ހ� ���P��'�^r��MW`<��΀Kg �𨗵���>���^�]��g�C�\MdJ~W�<&��+�f�lmp	GL�v��ɨS����clt�uԬ8.2��
�m=7��p�E����er>Ͳ}�eu��^>v�v��}Ǡ���:;�l�%W��FN�=��u�녽�ڪLl�9B�'.s'��k��+����.�^�F>��/#�X�v��f�=�0���8�G�����3ѫ���`9��| �j�/�W^��˥�:����RW2/Ч��y��h׍�tv5v'D��G���*�W���;ĭ���MQ��':�5���H/|�-��v2]�3+��.�.��}�8�.@��P��
��V��.T08
ÖN��|��6S����+��o�iE���+���������N�K���-�/ܪ}��/)��=<�=�}��؊~�j��} �-휖 ]��Y�[�TI6�=�o$��' �V+�e��T�q鉩x.p��m�*˗s8A�M��]U�Le��RpSt��C���5��攢0���%w1�tB����np���]�T@�E���nb�]�J�sL����4�j�5g�����;u�m��Y��d���/�y$�C>ۺ�s4��2b���d��l��Gv�=�Lgl�q>w�.��;�=%���$�X
D���yWu�k+��дֽ=�u��'�.%����\��Tp�P>:���='�|ȁ�vd?F{�A���F{b��^�\� ,.��h��QJ{���t��ϟRM���Ϊ�)Gq줺�ݮ�I�o�:י�j{H) 
�>��z{�L4W�P����,���{+�>�u�}l��F�={{�離��$�3�R)�����+�/N��e�h�jj����#\6V^����P=>C�>%��3�'����)�2E|�\�D��T[H���V|�\�_��ӭ#�A�w�3��*��^�}"�9��1}Ϭ��=9|G�OQ�Pd�Y����TKYxT`�V�W��氎���ƻ���j���'�r.u������E
���Rd�;_L-��O*-�I}��󊮤b��n��{V����~�n����e�c���~��	�mʪ^R���~+��'ה�fΚ�Qx���K�d�O{��2��F�c{ݐ�G���k�ԝ�[D��U抍�\q`5����9�Ld�Q��[�[��j�D'���m���a�".l�Ӽ��
�5vM2�-�f��΃w�P���	=�V9�Vc[r����s�dԶ�QP�.h�.���&�a��e'�[�ݥ�Dxﯾ��,�s�J��i�v�]��ХeM��ECL;���_Q]�aS��RP�������+�zU��r6R�>��򬛦��4W/�Cl���䖋1,��F�VU��uhޠb��p7un���q��V�	�o��A��N��J�{L	��:]�]�k
I��7]�Ul���`2��O��B2�S9�ͽ_R�FܮMPľ痬wkkj,���ZWN(��_�p��7+�SyWsL��G)�&������G��ں�����j�`�A�x/m���H.�����ź�i�b,�(�5���#����ʒ����讒�Bu���������3�+��SL�B�X�����d�
����J��w0�E�Lh�u���[t.���Ý��8bz��{�V$Nj�C���f�i!E%j��
���k��:0�B9;�$��b�8�%�+it
�x%��2�o��g;�cW�3t�p�$�T�.���Xä���y���lGo
��1N��98��-].�4䙽�DZୡr�	������\�Om�j�\�p�9us+s1k8Q�E��=�Ww�����{H��<��b)���ʮ�o;�W\��D
�Pz6����{�྆�e.�+��f�n��˻�S�m��#��,��(^���=E�|��l��I��R�ĞwL�u�)�' DU�����"��mP(P4��>ȉ�K��� ��h�ݸ�#�{��ͪ8њ��s��4�C;֬�DUS�r��dS#7J�;��ջ�m�r�;�C�sNE�:�\�7Ӏh�4���Z�o3�AԾ�X�q�!��k�JfV�T.�aΩ���)����F�D`O:֍���a�����ђ��+���N��<o�Z�wo��@�Xfe��ٻ'��gv�u�r����cQ�q���$��u�N'ث0g-��%��̙{a�x�(�bu�����	��u�*t\.+8���y% ���&ܾ=[C%}�f�w�x��}p�f@��uej��Eh,��sWUv+!�m$,��J�ˊ�L�[P1V>$k[�m<���Çv5i�J�J�����XЎ��Ӵz� ���P�;705�bɥ�{.�D�P��kz:�}:Y��z�U���A��ؐ붵�+b�koS��9�D��e�P�V]9�K7����j=�;Tr�vcX�*�)V��ױS�h��'����I+��I�oZ�û�2�u�x-]a1�N�����3�t�_$�+{��><o&L��{�,�w�g��o)u����}�[�T@P|PQ4AU�DMDEDPSUE5TSCEP�ES��AMU��%TQ4PS@ДPPD�RQQCUQ3ST�AMTW��3DMD�1EULM%�CT�ILLA41PSBU.XAEEIT�AILEEE-,M1D�E+E5QR�0QE-45ACBRU-M%1E%AH�DH��!@SM% D1CT�REUMUEJ�5)KADJO�9P�E%S@���f��鮺�5�=���w��0-�V��7rf�:�Y�$�jM�L���g;�Y���wg��Z"���KF�i���'w�@�5��2��+ԑ��K�p�1K�q�|=�	�:��#��J^��:�Q��rͪRk�vz}'�X>>dq�n�U�I\J;2�W�\�;�.i��z�o*=�h�O��΅
/����p���+�7���x���	h��_����^%�;/��1`��{-d��w=�R����6w���o�^���MŞ%+2ǫ�gK�T�#�=q�^s��}�ŋ>�45F:�B����z;��^�����1p�R��u�^�u(I�o@��/ߖ2jө��
�y�I;���!]M�j4�^gD�9�$<}H<<�ԃ�%��eN?q��r׽���1p&
�qF{�WU�b�ۉ����+��8�h���=ʈ�ȫ=T$��cnkqU�C Q9�C���<�n�T��ޫ}O���Ou�C7�a�lόn�1�^ir>X�O�p�}��FZ��5qdT�dL�����C�FZ7�R�w�������G��p^����+:�#��N��9}w|h\C�,ҩ!��mB�4%��뮜��fj���4wSz�r�y|���6�����\l����i�<����a����5��Hp�4e�Ԇ�3F�IЛ�T�ʒ��\�z���⤉�ѳ|�tei��2;�)�˭
�$�C�fș�2�٧�ƙF��:�F���j���l_wm��|���Q������ꌁN�D�#.N��fA�1�`�iT��q�;=c���3�G����[��=TG��F�,�ç���q�*]���,���>ڎ�J;#�GSN�(�	��=QSʳ�Ϫ�P�K��{���y�R�Oz 9��(ޘܴ�t�ힱKˮ�z�;_ഌ6Euf˗����/M�n_���^��Jk9�{X��m�ެ��ոٓ�����_�}{<
4}<�����/�t��>��|o�j���ȟnb��}U��H��a��W}��%_����q��ύ���'������l������铔�9+ZV���r~ۆ:z�z�u^G|�X��F��b�/�8o�E��pf�O"����g���Wٲ/w�<�2'��� *u�EĮ}��_⺐�=�(/�eN�JWy2��w{�/{�5�b��> ��ՕZn6��oD���a�/���s�\9��C���Chi�bjUȭ��^��a/a��$�Q'��2�ўF��� �x��?��>Α��θ|�Emu=��3~�1K�X��n�����@;���)k}Ɩ����ҋ�T|.m�φ+�]�;�t�{92�+��)����w�	'�s��d�R���OA�hr��XCv��qWlm��4����p[3/uV��NNVm�b���줻�%���סx%ӝ���`G)�詖�/n�Q�J�M�w�]k�1��ln��~�'|5��Mi�}#�߹\=�t׸���f�p@�Pe��n��|�t���e�=�MʓE���/f�1<�-]�m���;~�9q�v�?@��k�@�������������r�ٴ��{T+j��å�y�hh�us�=���cs��I����M�]}q6̖Ph��sJ`U����OI1ҽYF�=�
���^#|��OR'��pq7��@�����-nz�*�o{U[Ng��zB$zVӣqE�ʿ�n���ۆ���>5���cn����z�����;�x򜖉TR��VR��~6�b���v�w�;�4�?bw��yae'#ҍ���=��{=�Ja�5������Xp\e����zOw3#��k:��\Oh�kgz/��]����o�= ��^Y�=�|oO��醬e`w=��MI��5,�$�֔�'�����7.�87=�
1���ݳBv���p���	�ύ��s�/��3)|��{������u+���CV�I�Rm�����K�_n-6B������)o�сP�ڱ{Ȣ1K�8;&�J�>"��hǈsŹ�K��|���r�Cm�[/��ǈ�ܮr�䨛y�n�Wa��x"�Ml�e^1g�uֹ���܎�,k_;�����w0�yN	�!~
&��.���+`�U�:��к�t�sCt��//�#�O�c�&�%�l�vb~�N.�1�5�n�]z��j_�K lG�VE®��'#��Z�>t�WٹSl�N�}�>��溯w�f�Iۋ�%��~4gj��9�.3�g�;�=\M�r���K;�6�������;e� ��i�s=�bá�$�%��	h����U>����ژ���Q`>��=��),f]�u���x�Ǹ����v��#2��7{$�,	��b�R�>��Wc�>>��g��.�\��Չ��F�u1���,���q����c�=%��t���'����ʃT���Q��$qr�Ϣ��z�h�r�^.��W)>9}:����O��7���x+3*��}7���3`�&�	L�x*����W{���}\��C�CI�wQ}8�Z8���[{P���2\� ��$�h7 �=�#P�z��'ԑ���=��N�̓��f�k��ՙW.�m׀�U|f��,TB�-M��&_RqR���i���Q�����y���cmG�^�k��}�?�����k�>���o�d�!mrF�j3t�Z�*�6Wc�"��į$'�1#�<��\�򋅙��mW^��z�����Xw���Z{$�N�h6zZI��-�[Yҷyq��������A�ג��gz��fNGsFV'��B����G��}��9��"�˝�L.�
�;Ɔ}]+t��:�s�6�p���n��{Z����;��wF-s�4{�@�_Q���d�9��lOx��P}H�;�Xt��q'5F�=bY��e!�	]�p�}w!�H���9˽+{� �d�:��YpxמWfF��[Eq9�%i���u�U��F����~�n���1�3vU����4<�O8���\o���T�H�s��D������D����إ��ھ�%�v�xg)�^�#V�uWe�_j�B6z%���н>���`�˂�g�=8�^��pjW��e����\~
~��E^���1#�#�x�������4�w8���p��^#qo�8.IÄ�pN��=G��C����X|��w=�{b֩=Y��tqw��e��t��E5q����Q�*t�Y�R�,z��,gv�^�g;�ج����8��ˬ��xl������up�}���G]!��ב������:I��zQ�z;�{pp�3�o�ۺ�]M�x;�ã:'��v�m���}/ԃh�if����=*��|�N
������h�e�ja*��<��s[�ϛ�o���^�㷂Fr��ڗVo��[���V@"<��Į�h�Qo`Uי�&��k`I�xh�:�3��9�Wtc�t����g!�<=y�a�@2VGy#�Ůř%7�I�fVhg2�;Fa@�ʡ��e���w�����n[���H�;��!���o*g}A����t�ȧ>=!tw]�~��r �5��70 $w~ޫS�q'��.��x�{=�剟�Ϊ9���aۈ�u���][4��PF�S t����z��s^�B�Q9�b��~��c�ն��|{6�#��K�>莻�4.!̖jIX�"~��M^�Bj4v�R���{
Q�U�����kj�0�=��tϸ�1�\Ĥe���L�����R��to��K�1��J���5�k�[N��o�܄��=X|ǀ��p:r��[��c��n��o�~�>�(�>8f������ձ�zm.��ﻝ]y�U�u�z���s�� x�\{{��D������4����|������7�/O#�j���ܿU�?7�h�o�d�t+�/%^�^�Yw>�����![�羰�\���t�<5�Ńҝ��%t~�t�f�~"+����F<�-P��ΉsK{�Eo�r��W�~��||������˙���8�I�$(����3=���)D��#vEe
�У["(ҧTz�]�����+�	�|yp5�z���w
]�U�k��AM��r���;�[5ܹ��Ղ�G`�BM��ˇ������-�ǫ�6y%� �Un�oYu>j	J�>�7P��<�ydvKu}zy��	�~��뽦�r�֫=��U�������S�p��+q�E��q�~F����T�O6m]��y](��5�N��0�K�E����s�|_���ﻶ��ŕ:^�q�{���+�N�������mC����>��28?�#�����W~��C���%����ō��ˊ�뚾���R6��t��_�2���n�\�7U��>��^!*:�UQ��Ȕ��q��t�F9�л�l�Ntv�e�#�C�[�϶��J�I���WY�2�݋�=Օ�g�ΓǴ��_mB�5�=��f�p@�FX�`sr�+^}݀�w���p]����DV�!.z���Oz�9�)8v��pr��ه�J��Ur��n�;8-	7*H�{�}����`�v��m1�ӘOG���뾸�fK,���P;~�}7�훭��j�7�|Lt�VѺ=��)��m���o���z�=�3���}ՠc�Ɂs� nzi�zG��)Z�d��F����/k���*�ݸ\nb�nW�o��5����5V�����L"�d��1�bJ��SjTs1��G�Q�1Ԭ~�^�z�~���q|q�z���xgdu9Y+#	�����q�o;��o{lP;Ӵ�Pof͆���gTy�}C^�-:�Fv�
��t������mH ���d�U��]�c[Ӧ����?<��Li���2��>/k_�/�Q�R��j��Ȯț�/239�w�V{6���g��=� g �i�8�SG�����늕�����R�w�s����}3�R�'R������u�1�{�]F����Gu���g�G�za����:��fpoNg"}��9��'seq�w����X��������X��T��aD�%�=lG�NMoI[����>�n^�Ҭ1W ל�����:��t���XH�7����*$7
Fϻam�r�zFs�Ne���Q�C���Xo�R����L������I�ǳ&�{�z���{ߔ�?J�݁T�����/��)�;w<Jq2�k�;P�����s8O@OW��.tt��#�+kd�f���q�_��\n�v���>���/d�����rO)��t%��Z3�	�@Ҽ����y�Aw�ǫ�������+���;}]y����Aڈ2��y1�$?p��t;Ʋ���Y�tu�ml�-uX�}\0-��c=�mv�;�����(��3��~�N<~�]�IP+�J��ۭW�Sh�5�ҲZ�<��7��F��p}v-6�yz/L����[�mRHq�^"����/�H	=�l��w�Y��Q<�u	�v+m�Ȝmf�6�E�3Q�5k�V�[|�k8�}I�Wy������vSk8!A��Pr�y=-S��	ok���D���ޟ/]D��z$l�׃�����r��o�H7��뎟q��O#��&v��j��q�� ft��%�i6J��7y\U��/!�W#����r�[�X��{c=�r��RdguݱH�� r�$�h6���5��Tj}M�c̣R���t��M�)8�UG�h���/+��׀��8�Ib�T����2����*^��L�=�����v���9��j��g��9�6�y��tϸ����P�!Qs�	�ѳaD��4'��n�B�D֌�^��H���vٮ�t�ާR;�UQ��Ϭ��=9@u���2M"���{.Fc�|*�=�DǙ�^��\��Q�����]+{%��J���B}w"�y�:��;��;p��B��R��l1�Q�;���.��K���w]Y���i�j�=�u��������ʱճ�ض)����J��;���G�J'*�|l�T;��\���"���ھ��U�J���!�����;.s[*��_�=㵝�#.yb��T��g��2��w�^��k���/Pߪ���l{�!�ї� �@�ޫD����+�Nط��Y/�ŀѵ!�F�o�Χ���'m��)�w0�$jz�t��l���4S��v��+jl�b�Im˩g�s��1�T�6a�x�97}�R�\�D����T>��y�3���T��s�?�3����S�Q��u�7��3�q>>%��3�I�8���>��~���3�׃�����A����@��M��SW��׬��bʝ7x��b���Vi�hy��}k�zp��3�U)Z49�g_.��ﻩ�^�9z�#�YR̵�Fً��Ӯ����}6w�I_�63J ��+*e�q�t�?E���{��:'��v�_S�i؋�եΝ����:F뚾ѝ��t���1�$�wFXۍ�q<n�ۉ�n��]#��{�|��"������"��S#���x%Ӑ��,	��@����oU�����<�;7��:�J<s�s��*}��ϗH÷��#/���d��D(#J��@�ntD��������=m�(�i�^�6�~{�%�]m����������]��ʒC�6���w:�>�1P���W�����s�M	�x}��񫑷ھ{�ܬ��tϸ���˘�#,mDD��4,g��q����7�
��-��#�֣�z�YZuDV�L�\*���D"��������� "+�����PE��"+� ����PE�@��@DW��_����� "+Р��5 DW��"��@�� ���PE� DW�"+��(+$�k>Ɣ�0�k�B ���������JH��k�@�	P��h�(�L�*IH�BIET@	�I(TUQ���J(���JP���H(��%R�UJͤP�	�����b��i�c,m���lhŵ�5J��B+��:�h�6U�k�l  �  6�n�U��0���@R�.(�6b��̛5eZ�6��-����6R�%
-��.JaZ.�ۗl��p�k��r�,��]��ۻ�[[�E"C�8n�G�n�wZn�V��d�F\�]Y�]�ݱ�]mwwsM�w6��n���@	�m�6]�컺v��mfh�n�v����ݻ6�:�\�k���NQ͢T��.묈�IK��gl��f�+2�2��C6͐���3h��T. ]̡����V�aj�՘�56ZMfR�W \p�kd�)�m-��I���*l�bj�b��8�jj-d�6յ�R��ZejcQ�d,5�      SL�I$��   ���I*���`�4 4�ɓF�� �0F`"��	JT�L@�� �2a�12dф�14�&���) �i<�4�b=FM46C5'���5�]~������y���ֲ⾹BI������ ��y�D�@0 ��$���?�?�i.!$�I^O��?������`�$��C$$	$P�ЇjBHI!�.B �	I!����z���r?������������;�¥�˗�a���hz��?�~����f��E�`�~��~�}�]�&e���]��o�n����Uj�gG�i��ٴ�ݸt�9���WJ�Jn��1޵�+h�K��Z$r�M�-���a&�6&�#������x)ҕ��<�6Q��V�� i֋��|�E�kU����a+���b�uڱc�X�#E��4i��-�Y�ݶ��ʗb���Z��u9Gn�r
�+�ѷ��݌a`�e:�r�4��~j���uv˝kCs��P��B��r!/����In���m♄���e�����H���=śMm�5��Mk�n�wİ�¹�Z]g���m<�^:����D+��{t��ڔoa�1L�@��\��Ӕq��x��b��a��Yf��~�µ`.[b�t��lE�:i2�b\����M!́�U�J�h�`�mm5�,,�k
j�����#0�mR�(�4�B��Q:/'׵7,��F��H٬�������Oq�q&ovݰ�LZJ��x2�ev>�KZ��yMwkZl�Y��U�oX��cn�ͺz��JwA*�;�������\J��L�tb�`�������u	qXɵ�ee<Vpn�^�lh��a�ׄ�����E���Q�M�(3�L�P�٘n3��Z�&F��b�.β�yYh^*�-���f�s]t-��9�:�/9�;�1�b�U\ӵt��6+4r��+ͫ�S�����&��n��n1cv���5b�wM���G4�6mZ[)�>lӠV32�fX�#�m�k@E��":�k�Z���	9 u���vvPUT��^.}�욺(�:7��T�J[���ee�"�.	e-��4���m˂�0�Z#v�\��DS5�^�t���P��UK~��L��-m���Ke���̀�KkD,r�2&s�!--a+!25�5�1�\����P�b�Ve��1�˫6�6�cv�9PI��C���")�ĘL�1�2ݦ@���*lm��Vc֜9ffk��@G�b�i�e茜+	�V�jn��,�Z�cY׻������m��J^ed1�U�;��Q���1�X�꿎�"�+�wx��٦�:3	�\3,�Cb��%l��6V�ݬ�Fב��&RKU;��Ԟ[�N���ސ3"�[�flܬ (�:r�%lT�9���L�ˈ��m-�\��|A����44�r��5�h����G�	�i5�B�m/�f�f��_IdӁ#Y�wl֛5p��K|�
�fړ0Ҥ������;Ô*JcA�E�n�:&�`���^k��kvQw���G����h�,m%�C%h�r�V��XԮ�&�q��M�]d�1bF�2��Thk9M;)n��-��TK�uƊ�8���:������tUq|C�M�%<�B�ũ���l����+)��XF��z���կ��M�|0��*c��q$B�*�N�V�Q�X�Hx��n��ǒ�odC��;�1�XR��*�ú���H�]�a�i,�6�Qd؁�f�FX�"�{bd+ɋJ��!3#5y��;�y��Ŗ�sF̗���ݡGt�����g(����&IL�c��m�2�:��s%�p�!M�
w�
�?��wF��Vec'UAt�{J7�6ۊ�YvF�
���"�Չy��ǅ���Mi���Y��P+����i�&�����cY�V��WoA�`W�5��Й��D�{3�K��WB�]=�싍u"U�(1�D�r)z�Q8��)Y�h��A��6�l�m�����bՓE+T�����n��xNwn��?��^��t��E����p��d,nn{R��&[��IUxƧ�XEKl݋�vMK��j�cRoi*�Ҁ��k�f��I���	Fc�*J6����D��B�j��=�$a�a��q lb�RA�\fe��鹼�hmJ*�:<�%L��uZ�⹚�v0����-��	����n���c{Z�O>��,�RȻ9��F����A2e�J�ְ�.�w�3|�T��W[��6�t�M)5@J�u]�Q�w�;�n�8� [!�ow�l��7HmYy�L�^��~���ak[ϸ��ct�@���E�e2��6Z�7����j���lY�c6��E����7.�$�W�z��"Cj�^Q8�U	+]fꕣ4ei�GjU M�wH�ذ�!���ܱ������R��xl��cͨ��T��pT�v����J�!N�V:Y��b	E�j_^�M�kA5����bL��%�S��.�+:�Y�Ҟ#$���{p�,E�1d����kE�P���i�P8I:���#,�m��o�>���z��2���4���X����k(i�(�/ �\��������B�S
U�R��y��F4[�V�Y���Ŋ�#ͳh��B��Vವ;i�xv�Ǖ,^�ɑe�]�P��P*�cm�I-�g�	;�7���cc���9>Bj���(��h�{j^���Y-��̲�ޛ���
�g���kL2�����7B)tJ��-�ys�i�Q� 8��p�%�n�5��n֍x*i&[�lAI���eVGi�Te���[;e<�dS�̺��@ٗw��ڭ��CM�ي�"$�M#}��<��?�B���B��[�*�-5�S:�%X�b�Y�Y6,����]�gX�τ?����gޟ�c��|�F���?>�ϥ��� &���{/'�������yqX����$�I+ �r�C6V�`����If!*TU���B��s����1��b43��1��\h���B
RV�d̺:�#�Û��b�>���ky?��Bim���^��R�y�{u�a��4�-�S_M��ǌ$����K�m�&t��Odc��.r�ϯ!��g��pq7���*:����e������>�h���Wl���%��:����q�a՞��f�z�
Q�k�1��3˥-�9ƺN|o�ȴ��l�ݑ�;hL�ye���Hu�+H5����k{��2^���X=�Qz�
��3�bV���ի'��ve	8^Q�ŔW�Ld���n*�1(�����E���-g�� S�h�b��8���[Ƙ����-ږ�	���Į�+���Wf�J�\�+�x��ըU^Alp�g��R��b"_a�,��X�,?Cݾ"��s�<�˲�ԉV�W(^6-���S�Fm����Z#�\�n���%� �z>Mu�Ž���c�䤛�t�e�KC)Ny[�$y����I����kۧdX�0�h�*�wG��j�*S�b��;v���^�*�+��7ms�4�)�	:���<�>�gu��	��;4Z3c-T:�[��C�4�3hڣ@�-�]ذQ ƻ��]o�iJ�II�i��=eU�Z���ݢ��5�}�w���;^M='��=�:��=&f��u�Ѥ��KY�X��ذ���ޕl�XP�����@�nwG܅Gf&�o>�V����k�a�c$�Q�S`c��&IW��=�{Zet�ѵr�0T�6HkC��Y��7X��bk�x桺2��f��e��pJ�h9�娯93�S����;�C�>�E���!����eof���/r�7��4i�-�����{w��I۽|��c0)�}]�Xߖ�%��� D�:�M
�Q�똫D�Y�{���zp�q*2^Q?[#:u�)��j>
Ϊ�{x2��V�\�EH�l6y�����0��\�vǐ
5�XAJ���a�J�<��'y�R�K���+��g.J�xP�n�WH#Z "IyFd�ۖ3�Z*���&�CD���=���Ny� \�I�1k��n��}B��;Q��LչSn�+(��Wq�ũjڻνE���Xz��*,����;3��ⴌ�"
��#�f1e��x���q�Db2�.�\u��&��5�D�u�B���[J�U5M|�%�K��GYwc�`
l�U��+/d��f+\ F��u��i-�'u�R|�˝*m3���YOp�]N�o���.���4[�r����0���s���h�.��ﲂ!��i���ܺ:�fɄ�v��rW]t��6Gv����K6m�ح�G.eA�fr��q�2��A-�5����e���a��F�����9�q�f��(򭢶�;<.���x�t��^��׷�xk�d�罺.��x�àu9�PH�T*U��`觔RGou0;R�P��0T҆P���:��IR�8d=DV�Ĭ�a�*uML�I驘���蔷l�Pg��_�R�u�fk�(�yx�""E�%�'s%��˗�d`X��.�P�ڡ���1\q��xT�6u_D5��J2�����*�����'t1��wN�b��t�!��Ӵ������'V�\�:��n��'[e�nڢ����K��n�M.;�V}f����$���ù!*��ǔ��u��7���9�k����d]���v�r֠"@����5�m]�z���v������[��:�w�rJ���1��w����,��K(�R��ȹ�
/^�Ox�LzQ�@�6���sp�8��bv��ZM���/��ƘT�W�6�{3&�j���fN+�����]�{M�ujN��跄!�X��4ҥ�wLp��2Թ(���Y�5ΖwD}yi�y�n��2�s��"����t�*�J ^�4��wp�Xuv�A�ZC��JV����Q�H����"�M�.�"���O%�y!�������,�B��	�1YJ�j���͝�^�RX���������QH�n�n�K�i���p�-�\�<��B��)����퓮����-*��@�+K���j��uv�����mط��t�H�20�O�k���i5��;]VG5[|%�n���#Z�^��PD==zw�N�͜�h�KK/l��ҷ�#X�c:r��e��ۼ�cO2$�D�qn��<��9�5(�����e,~�{��{XR�2+;��1�!�.kU�㲴m����u۵z����[9��ޛ =z�]kn�%���f�[Җ�C�K�86�!��.�nSVI췽�15�{�X�/e�)�������HW6ާ�4��lٱ3�<4t���]����oVQ����gL�l�0kU
�,�r����.�b�k�f��D�1�������!Y�l�s ��������5����V�q0�<��P�n�d���C'q���NSb�'aq�7X�Zc��g)ïS�G��I$�D�I$�Er��J+죉��1��͘\�[w/�`��$K��\�4��s7�{Vc�t�o;j^�.�f\��<�f�I$�H;����DT��'��w�I���wG$�.II$�%���/�q�B�+d�v�Ғ9��I*��Vo�9$�I$�I$�I$�I$�I$�I$rI$��$�I$�H�I$�I$�I$�%k��/����������oտ����BI��o�	$ 'ծ�$'�C�ߢ���C $��G���]���П��h�b�Pk�Wna��]Ru�NN�Δ1]�#	(b�=�rb���ç�W��s��ͣ�X�UHun��E�>Bp�I���ػ�wX�{Д2�v�3FL޾{���1��L����>ĶX��m�������}�fڇͷG:(�D1:��U�Qк6��f��T�ʻ�5b�j��ӓq)�Yp�S5�ʱFfq���Φ+�����h���Fb�RJόa��c%�{{ǁ̲��\^͑"�&�W8�U+���QR]�JP��lnbj�nVur)Jys��.�}�V�f�!����d���[bm�s,�A��������
�*\�F�aUڜ�IֽŹ�S*��֗R��/���e/hۧS�mms��D��u!}�U��a�a����Up /:3*.��s8�]X���l�n+�S�p�Α����.�}�R�>�(+禵�Z�v��bh���8��R:܄=�`/P�������2��ˊ�w��K59ي��=vc,�s�ΊC]Y��۽�	��+ Y@7[���Oua;ϛ{G�p�-U�����ڸ����|���>��l��_�\�o^��Ѩ��q�52��1�"��5����7u��%��jJ�\A�R��bm "븝o3/�=vEo�(�έ����2귱�J��D�y��ǩ���=X&�Ix4����GUn�����EDgwA�q0f�ݡk�I�j(�t��:��K�ؖ���3VМ.L�F��ǥ LČOM���f�o*ݦ���|����N���7�5
������`Y��â3����yLv f�o���6݅Ïyb�
S�&\���ͨ������t��������#X: ��ɇL��6n�u��M���c=Hռ�/oF�(T'�����U�� e	]�'�q�#+�w	���4���tҞ���gVAM<0c���v�&���٫���t�@%�ս���v:ڼ�����Ĭ�� �M�x�
$�2����k� Cn=�B6�C)99����ۻ�2��uݦҵ�n�'���Ku�<�<��2���/�"ݗΘ�[w��'�l�[��iջ��sG
�N��&���v��26�9d��y�ê7F��m[w�;�z��Vn�)�6�L��Վ��"�O�>z���t����ϯ�Vp�e�(Ԇ�'�U��HLrhD�1Q6tof�0��Ô�ĮO��K(局P��e�f�s]=��oB�t ܫ�f�����EV�k��$��c�]�i��e��X�F��Gyݔ��4f9}�K�F���Ą�r٥%*� Tc�2�F�֊I��J��n�c�
�i���6�a;����%L���Uw]�Gz�s�#p�c�p��o�$���`��N*1Q��"��%�)��׹�YP;�/WU�op���S���u̢����BLh�Wu̷ri��:D�G\�gt������B��Ӵr�K���ՅVN�r"�PQ�>��[,\T����4O���*�˥ɐx.�Wv��HpL��(���6����]Mf�)��
mS7hΊ�
=T�ѷ&�hR!RJb��Gj�yWKM�1�=O�:��V��Ou�+Q;�2��gp'7
*�v2�QL��w^JSy����-f�ʟ7�w�����װ;�d#Ÿ��{ڛ;3��\�B�򶡻�W�s&�0�]D��\E���Q�A�5���*�|�����ZPQu�v��Zw�@�%n�Ӈ�4s�cz���xhM��ج��+6��B����+���Uu]����(N�������If5����57]���	�����yw]�˭��ak*ĉ�X�!�S��U�K8%t�����R�q�;��{�N��;�[�ݑ�� ��b��2X�f��"l�A�fB����t˂�N�h��B��ٔ¸�h�[ʶ�����$�n��B��6�Z�U�
Gh�gPL�Wo�*٭��&�N��KRD��f��ƭ+0��\�0���׼01c:q����I�Qg|l�G�m��͓N<{|T�j+�	�\���T���_9B��P�+�S)�.�Mu�]X��	a��=��mk���L�
力LԺb��dj���X�r�L&i��o�^�[/35��k�Ӱ�ư���U �c'�c�E>�WV�u ���e�+��J͗�6Iޏ!z��WvU�֬{�����q)�SpK��r5X�P ��"O��'<�t��¦X,��٧t/#�Z���k-�%fH����3BQ�����f�e���±���L��4m�J�M���E�ruϋ2���nI�;8wYͷ��-���K�N��m�+�ʺ��*=���V딶6kA�!��%91)�dbVV�u#J>F���}\�7Z�K6�:��6�kr���sI�%uR��+��|6�c����r�ܣ��٫���i��}|�������4�Yڪ^�EX�T{�j�'�j���GG	���)��;�����ZP�%ݍ
B�xSG�VEyU�1�$�3YP���W�S+t[�00z��T���Ǜ�mɶ.��nӚx�7�Xt�k���
�-q9�����c3X{s�m��������Eza�+t�Y�u���+��9)w&�XP��[��%�y�Q���a,�V�aO��+a�����
��L�����jvb{P��Ϛ{7��[�X{��ֻ�X�Z�w����k�O��$�����2B�`��p=�Œ�Bʏ�:����U����j��Y�N���K����#�X�S��>��t&FS ��W�^���:B�Ӿ=����1�ɧ�iE�j\7��V�KܣoOZ�J*M��늕�_]������ת��K	�����,h#��r�7rҕ-!�w��]��l�34^�����u��r^vE�����#��+���*�in���:��̘b�ĭ�Y�Ѵ�si�sH]4.�[�IC���֦]���^���xt���c.����-M�,��gG$��$��Z���`y�A�e1b̡�,UAU`�IQ'ZcJ�o�����s���*��.��LQLX,SM*D`���M2���.�
*�m�a(�M#��1T������M��UR��RE��-��Kj���U(S�/�d�P��U�i,WIi-����H(�2�0���U�n�e��9�Q?ܮ����{G�[�i��E�)0ۛ܎u�'f����kI���u��4�����E�|u��t8�WN�3�sܧ�k��G@���C]�!����,�d����Gnu�7U���q���%�Af�{�/&�N�M^����Yn�p����z���4���"�绊�W�.
�E>;������z���
�v��7zZ^Z&(@o4������l;uH��w} ��������:�QB�{=�����_%����H�o�l���nj]5�]��+@��8��G����ga�.~��׹בH>��}K���[�O��PRo��1����]�;�l���oV��wo��j�yV�tb�Z��R#���6�g�I�[
n';����X���tD�[��1���M�.�3��nh�U�S̓gs���E�o�p�tWe��ǟ���~�^��i����f,ehl2Ԇ��{�����{��r���W83L��B�}5v�-Q��Nq����z�L�]��׫7n��9\5�p w�V� k��q~�g]'7�k{�~��5K�~�H�o<9���b�˜Zmvm��e�zm�>�q:=�d�'����]�A��0ȝ�׹�w����x��J�n#��Mѝ-_r�=�|iE��C�o3�k}��h���n+ �$'����]��N�޶�2q� �!�i�b�U�W�w�i�qwG�)�#N����X53��$Ԟ㾛�9����+kZ��9չ6�/.~����o{�]�����k�M?5B6�<�=��������n�L�h=�mU�6��W���Yâ�i@�W[-����&�'5�)ҺH�z\�Q{gP��mdαșی��%�վO�;yk"�_b#��s֭���Y��pd�R�30p�Mj��f�4����=P9�y
}���U\sە�!�m�;;�+9�V᩼����Z]�P��5���|��8m@��as�~�# ��h ]n	<pj��s�j4i�K��+��Jjp�Sd�⫈;z-S��j����Wp�E� ��{}���4��g<��(R��2���
��[�N��F�ܲ�ukox�tv|�r.&�����bݠ�`^�d���'u�E_h3�ݏ-����
��^�T��4�=d`(̾"�{*
z�ckl�Z��U`r�Ζ��N��v�N>αاso\���ui��4�;����޴�fG��>-���{k�u���}�7�div|�?l���k|�9oz�˶ޚ��KcAt���t���s�8{-��AX�	۾S���yhwH�����n^�JɱRR	/!�1�ٶ���оw���k�����N˄{�6{m۱/=y��"���r9�Z9���D:�FU��U���yv�NV�G֫Dg\Ȗ�����*=�2�ҷ�y��z��_���ۂO�tszx�A��&x,��C�6�yVqh�xns�����w#�=���We
�9��T�E{��V[ԭ�{4�[��'&�6(������$_+Y����&�C�A喡Oq�����+����-�U����n�Pr�q=����[o) F�8ʰ�	:�C+F�ױ�ɗ/C�����3����#w���� Sj�Ϯ'�۪�׿|�U�<�>X]�{�K�ȉ���{�Peڷ�_>׻��Ohy6��+{�s��̎&�1�1�WB���3��H��a�R�%J��Ѿ�ʯk:�z�N����@��]��o�:5{<�F��n�R�ٶl)�u�G��3]C)���v3h��}x)rhރnTu��\{`�pÏ��� �ζ�p�J���^uwGe�r;�1��;ǔ�m~� �gb�;�:��f��xp�O���)S∺'�\�mX��s&8�}��W@���58�{d�\�?��9�(���MS��#�7|59��Z��^B�%�<��3.��Wg�g�w7y�7�����q��l�0<�����\�~���0V�w�9�=F籘�%y=z�����C0��Nۅ�K��l�AΖ{5^�][-�V�	=�.+���OV�m�l�	s���ԗ�M7��-d�$��#ff�5s�;�wj��
�Fib�D�r����8��*FT7ԛ���ع�jB23�GE4�ȅKoU�']2��Y����|e�og�<AX�mK5��2�K�)(
��D��Ǭ�ӎ-��42�%���
R�'�<Z{s�#�֎�����U*N�H���tP���a���Ɩ���6`�,*]���,��k����U."�.�U6�̜�V2T�}e�r3��h��f�`�c U����p曣���R�Sk!]��NoF��2�XVF>^S����s�Z�:���w0G�mˑbg�M���h����ڹwi���uf��!$Ѫr�|�Z���c�æ��kU�
H�9���u^�\�p��3M̗{Xjز2��fue�N�fc]�k&�*K��*J54����b�h�洨��'L|�g�� 4
ݺ��ڌ�}��ٽ��U�P�1˱���{���C�3����&�Œ��\D{W�f�Р�!��Ttn�ֻ��n���ǜ4�z�}YR�����m`b����m�A�Z=�
)�s�F��kh�3+N掩��B��z�� f�X�\���&"�M.�+A�ņ��k�	��]�r�8X�� �Nݵ�B��}Yz6��4��b��k8wU�J�F��*��IJ�q�6����5;\������R�ѶJ�#Λ�����'Gg�D	��eANb��;���Ģ��f.��f0���u ҤNM��F��C��������`�YI
i���MTЕMuK-�SI�M�f��e%�U�R����ʐQe���e+S���R����"!IC5t+m�i��J>Q��UK
��5E�l*��ESIih)�*Х�Si)�P���`�e1AfZ�(�Q���)�.�]��dn�"�A`�L����B�hZICuJUQP�]2�Jc�@�"�*ꮤ��0Ҧ�S��,�a�]$����k�ߓ�Y��x%k�(���vh�^Fr�<]��}� ��a����?��99Nڥ����~e�\O�:W��B����[��	g�����y{p����ġ����ˏ�ޅ�(�ׁ�lk��ٸOvl-��"o �v��
��<Y�ӷM�����9Ӯ[���L��f�:���΃�Ų��N�m-�O��IF�Ѣ�F��3�眒�0.���7�6�vc�S�g%N
�Q(Pٺ	(�T6�|�5��6�D���U�\�r�JC�r�佘���W�[�o�k���ww�DX�֞�+�vU��5����������龳�D�m�o�0��"P��^��Wy�*�^�-��\�������s�uu��8(!G=�NC��KR��OY���U��]�;o��Z���W�о(�Bi�[�W��t�rF3U]������зu"pWP�Z)_��4nيI�7Mˏ����O3��^����k��9�=ۙ&)ݶTF���o��ֺ�����Rߘ���`j�#��e�ٔ�Gd
��Q�V�D��ݐ^���C�i��VbM�*,�a����+hNy�d���U��F���9ܬ:��8����]�a�7�|��z�k~]��=�5�]^��%r�gt�|���篔�gX��W���[� 5A�X���1�<���º����������^��� gq'��\��Ԏ��_}q���~Y[���s��5�}��M������nw4��g��6�Ѻ�UǷ���<�^�é���	K=�& �{lS�d�́�T��L0!��&P<�d�$�9ShC�!�5G�!�omw�>rRO��C�$���a'�4�:�2É!� y�߾{�}x�&��yPP�I��L5��2e�lL�)��@�k��|�}����kIB�RC)�C���|a/�AI�q��I�@>d�<��	a� [�hL$���`N��X`(x����8��c���>vHm��$�SL�@����	%����!��By��hY;X����)^�{ʭ�;��[�bI;\�v��&�Y@��e���v��D;�hS��b���襽td��{���B�3�|��-���Ha	WP��J�(}�HC�Bٳ4}C^���o9�n�4�(�<�J@)$�����2B���e�hO2Be'X|�={�^ߞ�{�B�L!��&�N��? ��d&S�!�L����9�o�ֱ�[	��Ha��g��T����) X���|HL��q�{���`,!6�|�4�l��d��W$/THi�� Pc9��z�|��ж�����C�� i��'P�h��d�P-$Ϩl�a�������[���	2�a����
I2���HRd!�M2d��XI����~�����M':j���d��l�A'�!�[�$��m���{�Ϛܐ��6�0��q!8��P�,�8�M��,WRC��y�U���k���~4���:�q�
I:�q�pd�!N�i$�d�Ha�������'����}H!'�,��<�S
��#���+��R�<���rɂ�N�nۇ�s����{�f��B k��k�C,����х��:�/�-y��C��(���N0�{����;�vE��,�@���P8�i!�����C�I,� u��sؾ�����I e L��7P-�d:�>0�)���!��9��__g��@8�L�y�y��`B�P|a2�Z�d0�Za�Hk��V59����B�|I1� �'�C�!L%$��bC%���f�C̆�w{������@�T��,�BI3ʁ�M� �$�d&ɆH|��t~{λ�RC�d2��h��43GXB�V�:�`�B���g���>w�����:��$���- u���f��a>$��2�i������ߝ'���$��fA��āĚa�&�:�2�ad��W�������{$8�����,���]�!�:�:�q	l��4�g�$7�[���^��o+���KfP�#�b"�V�fyx��K��?7��%��UoZ��I��}_W�N{�Ϲ��L d�b�M�C�O���AL�H�*aA��5��M\�] ���*Gy��Y�� N�j�
Y7�c�kc��Y"%���	@�%P�١:��
s�S�D�����L�_h�u�{މY�k�.Z.ݖ����M�ND�קm:d��k���y�g
�2��X 5�2���뢨�ч'oo�2��6v��\-�&+�k�œ���٨�%>��Ȼ�qS�ݟ���0�u�1���2v%T��x�'���sskw�{�¤?j�y[�в�̽��l��y[ﲡz�w.j���\���xann��V��k���c rv��<��ǹ-ù�{[�'���P=է��C�T�ټQk���x��Y.Cl��1�u�s���PJ����m��x��H[�h�7�Y$(�o�p�B� O�1z��=��lH͊�Uv�Y����~��S���v&t[��ܰc�f���z��^��u|�[��c�i��ھ���}��+��R.9��AN�\��ffB��Γ�i{�ppK����2}3iSk�$̎M>E�(��6��2q�ҭ��b�!޺�+;5�U{�wi^E�kf�/�GG�ޅˋ�ͭ�y�+l������ٞ�d�//ڠ#��:�=	`y���v���ԍ��f�K]�����r�"��i7��&�z��N�XN�������x��"����eq��s�m�v��E�v��x�
�X�|�|��ͱnx�O�Y��E_E��,�n}���3y����f�a�kl����~�k�2Yӵ>��lKP�Vy���R\�X�f���sS����6t�����tgu�9�2��Ȧ��Z�;�%y��b�n~��f9���(����&�K�͜��V�w��·9��om�]�Nw�W��_�0�.�J����vN��m�ԛ�����v�ֱ�쬰�f3��vi��l�-C'v�S#�¨c+F�.���fh=���V�ɋ��:%��ӿ�P��Sor�F�&�901d��y[8Y�9�M� .�ʔo�Gc�wL�{�k��Q�he�a���-ҼD�6D��i�ҕ��i���G0�8�3�0�_c\q�}˗�+̙|�R �C�6�0{f������t��Ev��R�_�_��߈�ޫf�_�-;�6mu9����"9����lY+��v�eϜ���v��9<��U�.T�Y�sv;���@��#O+E��b�GP�����k{�̻R5���Ӕ����M�uNWW���B�@�T�Y�{�N��kIr�nV4Dz�h����ɱ���A^gMN�a<LX-oQ�!�r��9V<eY���%E�u S�$�g��k�d�u�,�4���˚��q�q�&N����K&�f��L9�{n;x�께�ư�m�l6�e�`9H��'G$��$�������ߕ�?B��O��*Ke��
��!�i�Z��H�L�Ʉ��a�2�T{�(,H}��L%�Xm��H�Yi����M��1D��f��!�BkUH{�}�u��m��僇�kh�㳔fK��-vY�����yOfw߭yY�fFM�v����2�?�����:$W����\�NAmu�(��,��ܐ���z��:p��9��h�9V~}�c��&n�Y�R��@�m>+��sptӂwn$c�]-zuĽ��i�&�sp�73�����B��c'��\:�o6��F�}�0E����d �+� ��$��c�+����n�ۤv]o���o��r��^=k���7KVws4mm�M"�����������e��b6+.�z�vϳ;�;
����b�����&�R�3���c A���}\�%�F���]������^�8�f9��ZƥL�h[��4�r��v_b��VCڴ�{�˓r�ngvw%�"q�ؚ7h�[t��sd�o�5V�{��dW�R��~��g�4U�3���s�f�!%��Z�oo~�a� ��m5u��=��W�2�-��ryU��  x��v*�R��R2��DR�{��w��ˀӦ�}�hI��{��/�Q.En�Qm�X�t���G���U�][�8��u��5�[��Z�g{��M=�ވ�;O�O���.�_n����y1�(ӎכ�^Ws}1����Dp�Ζ7XJ^dJ�"�Jp&�u��.~��y�ٷ�Z�}Z��!u�f�ׯ_'�!q�XJ��NYrs���\Kok�x�y��'�-�����_�+w���i�J	����SD����t��^[gwi/Vm���%P	�Zm��y��r����˥�Ye�R�5^�]Vu�F�pN���=��IW=G�צ���~��p�=iżz�Y�A>��(�+^.����^C���I)3kƽ�^�����uxq���	e�!T�gP��]4�8�r�U��iM�(4>wӶDb�ӊ��Y>�Rz�;�>���J�1o�..@�����u]={�Uõi���^Q�x���7{R�'��r
���yV-�8D+��̕��"��m�%g_�4�v����ۏ�gp1�5��G��c��k��q����C�HG����-���ya?w��[Z�{u���9�"G����]Diw4h�@�X�b�E]_
"/%�|�=��iV�V�r~���p�mЏ�}�ȓ$�y.�B��-Ļ3�{����Դ���mP����I_]S�����,
o��"��@�y�G{7zVȆM"g�o�u�pwN���f�!�;Y^�P�{ɬ�E��A<�Vk��O�'��&w���+A(8�o���	ھXF�N�+���C�0��F�����b�ܩH]~�qC.�EoE����ҟ:�t��۞�:�|�|�a^��p�[�&�R�I�ޞJ������?VޜSVB���l��*8���`GӫH�'5��L�Y��^asz-�=�"�Y:p>�}���C��?k�؋��9C����;���d�֧m��&o�⪯�X�؃{]eD�a6���oN��pp�V�����ɴ�T�r޾�=:���yd�S&�i��x
�k|���M�ݓl�1�ʻ2�����t��,���ɇ��O�"w���Z��I|��Ͻ��4o�O�k��qO����45��)�ݟ+Un�px.�"�eG�{&���;�e{��F�ʺ�@��]�{�6�8���]�>ޏ�a�ݓ��d{��o�������ΗڮGа'y�����ϼ]���]h�,�¼�߉��ٓ�W:�L$k�R>�w�mߍtC֫��g�w�#��:ca���I)����G{��k���V�+uK��NW*�A%�{������s�:��i���Xn9^,6&^NF�p�,e3�O��0��V��u�vf�TK�kۑj�!'gy���Q7ܣ�;뿜	{��o6��W˪MY�[�s���yڷ��8��R�\��B��gqoY��MZW垸��m��X�MwÏ7%���Jƽ(�����J{�z�F�.��,g�U��K����1K�3ji�oQ�1����o����E�Ch��༖��������[��%~.�kس������j����5q�̷�{'	�ݡ���)����Z�������V�(��`=��1D����wKp���Y���ƌ�[��y/�	NŔ�5�r��]S�j�IH"*�,.�)�U-b�S"v+&��';v��sLp����E�����c���9�Jj�_眙�+s�����v�v���Wp��lH��H�����#�Ƀ%JqO*�6���v5:T3MV^���x�ۣ+��ؙ�ON"�8MN4F���jԻM'�g.T�-Ύu���HUrX� T�f��ݨ�⛾�5��+�b�[=e�3b��(�dәۉ͜*tb���e6@-c&ehfn�Ϸ���kC�#�"�F��@�-ɒ���­��G�Y�Q�2v*����1����J��Tf"^��V֧�8��͜���;��\��EĶ�5d�Ǆ���*t��;3+��jeK��/���q�[��H��ٔt���N�e�3 �]� ��m��O\t�]wN5��\�����F�y�-|L�ڛ���/o�2�C��)Fy�K�Ԣq�{�*iN�9����7VS�6������4�J�S�x�g w���'aX�u����P�J�7�s�S��e�h�yj���Pwy�{3��b�p��W$[�j�9A$�M(6ʻ�K!{�s�F�8�Z8�"�r��9֛ȋ6žۦ�[��
��I�Z<�̡̲D�Wη -�^�86��d�H�KW$�qI%~�}�<"=�Dz2Pi��a��C̤���RUQ��S6�)6�d�EQH�Qb���Vd���%�)TTUF��4��D�m���(@@2���-�1�cf6ǟ5��j��L������DqZVV~�� �Z�_��H��V�1[�yU���G��(�7��ү�.1N|!u�0L_N��4�8�Wgω��9�u]ga�`�
u��q���^��[��>�F+�L�rvڻ���br>��R�R0�¼k{zlS��e�v�Mp�ODy<ź����2{f����8΋UTGL����\�ɕt�czf�Y��to$����Ś�d�X%ur�g+�=����V�i��J��� ��5\�yȹ(�l�pq�#j�ժT��tf��[����eC>�^E~��.�;��5ݎ�M�R�F�#9,��]�l�n�U-:������<�ˁS�/sq��3D���w^U�\�5;漵`NG���V���Y.H��y�+Y�)Ԋ�J�I�1�&!����ff�՚��i3\�#i�uc1Ì��f��6�6���|���?��#Q�~��6��r�{����}@��
r��^��R���.�b����y����t�`�VN��䱽�q�(���L,��]�^����B2�ڙ�ĺ���3u�s�0,'!l��ݫrf�:��/�E�
Wt*�Oy�gw�25�3/C�i�Θ��tm[D^j��P{w؛�>���]܍��E\�Aؖ,�ǷN�覨Z�n�.�2���ǻX�f�${o�����Z�I���k��3O~�J�?#}�	']c.����,�J{<G����`�S_�*�m�)���7k.I�����M9^��]�v�k�>�j��}�ѧ��X"�'�ry���:��o�cB�'="����p��<Sy�Xz���
V���v�S���o�ߨ�(��	���u������CI3[*���̌y�0���F��{�g���ʭ���az�Vr�>0����&��w�}\����W柋4k�͊W�oG̋��Wh>>�\����^^)�>��Eǳ��aX�\�����N�c�I�M!y���9�ֻ�ui-��кG��q�T�mVҌ��c]�iǢ=�#:f>�hb�┃���ݕ�d�=L��
xl5��������x���w�Ώf�������;EԸ��rA1��n�3f. 0\�����3�VP�7]y.�f�p�%3x�7T�7�m3�o&&R����t�pW��K�nڶ6-b�WU�4�+]�,�H�Ƕ.7yw����Mҽ���!̩�5�޶���Iw?+�V��˲܎In~W�Ѫ(��^�٬^�{.��k3)��7��C��n�L��ǹr��A���V #D�]X��'�
Xn���OLG���:��.=f|OP1{"�NYe�$ʏl�g�"�ǰ�;0�F]gc�H�>5��
x�G�"{�C�,�S�d"����P����Ӊ��5⵿kKz���r���DMP�P����S��S;�!�@���������=j��z�[^�殓����=ʙM%�=F=�Z��h�U�x�@���=W��ŗ��⺀�J^��꼃�:J�d#'8a���y�ŦTo�+�~�������`J��p�PsP9:�����q�<���7c���2���2���;�¹	r�)�e��˩f��,߬١�n�g;���1�^1���ty�-�e�F�< c�K��=���}q�T�n�ѣo�
e�p�k�	��;Rn�깋��Yi�ܫ0�Ӷc���_\aj�NEǝHs.��ؘ�1�7H:�O:�º�l׃��b��^o����/%xk�2��Y�L�
l����N��J=x�^œ�ps���y1���f�mS+��v]ZC�q_]78�r6�t]�d��(K	���#x�*���,U6��kM��-�Ӗ����3ک���-�����U볷�{~��a�p`�@B�k���/'ۏR;e��Mv�����&�S[��/��곽�\����b�
X*��G�ۗ[sEK�y����8g/K�6��q�^+�������ޓ5���vh�;Ƽ0R�ik��w:^3��Ѽ�ZC���f��v�Q���v���g1[�L�Ze�E�1ڏ*������ӹlU�68Vq� U�G��ځm�US��9���r�v\Jj��6*.ȃ} ^�-�Ը��@.��R=������/��������F!���i��4��ۿ+���h�C�h��
�����Ƿ�׵�Ι�gyE'uWU*�/�ݹþ7��ϱי���)�Q��;�Zp��J�}<�{�@]K��P��c�r��O��Sx�h�7���f���OuF��K�ۃZ�+��:M#�{����mRV*�vJ��������k�.��l�q��j�����p�(��z�a�s�F�)�Ԋ�_�;L(^���[5G��7�)�x�=�ns��{�GOz׺"��*��!�{�Y�R�-�J���V�-��gr��;h���gs��M=����5������� �Ǖ�>�n�^g�gv��M�^��.��]p��"<�^��>U+�cb�a���;{t���D"�{}-������о���cT��4	3p	s���v��!@u��5�p���vM�m?K�`]z�������7B����w7E }5�OLƀ�i�^p��e� �.ҧ�購\�cѲt�z 02=y1 �@�kX��;�f�n�����8���nّ6ʛ�9ۙY�hS�QC�^,x�>�]��/z�y
��R�W�Q����u�:�B���V���Yr�xl�+s��[�����k9-�}b��q��d�L��u��<���;1Arʩb�ݝ�@'WM�JP���|P�9c�9�e:S	���L�T���n��㧊s�]��P�qLޫ�X:����iZ�G;P����fL��[�i�.\G�v����3&h���ˬ������8n��vl�[ˈ��P�d�q��eZsn��K&P���H�9W6.F�$s8.��hl��X��qҺ���aUjU:�݊p���hD5
(�^�K��뼁F˫�:iΕ{?d�.���4�Q{`Np*�3A��͵W�su�c�%���P��=h������t2�+6��$t+f�'�m�7J)
�3����튂�:<�Bk�
��uյ�c�l��5m�jHKU�S�L4X�k��6�Tk%p�fnn�N#Y���;�M��3�,��Z���iX�Q�V����n�$�7�R�>���c�_v��:�j��%jV��FHgr�k��s�SdŹp2��N1&M�9 8��+[5��Nk�Ν)+�)rt�HڒH7��5_S,"�CR
B[$�L2�XpњKa	l��E�,))�	Hi0���9J�	L
d��D)\��,��^jKHb��C	�WJ@bL��L�k��</��k�p��[�_L��ivd|�s���_2���p� ��+�u~;���["�A1e7�oB����8Mz�u0 =t����^{ZayJx���RS��^M�y�h�������CR�˥@����y^$�6��8K�����4��C�
�}��O{μ+	�
l�4٫�\ l�B%&ǜ��5n�=��u��1�֮������J5��z�������`�4���,�y{w�<rg��u�wA��k��]袝+|��&�Պ3�c]�l�	^�>GPK5b�W�f���e��_�������aQ�5.�}3>��nޓ�=��{(�>���Q�ݘ�*P��7�1���9;6�ꪡ��u�z~�5��n]UB���z���kN�u�7��hyhe�.�X�F�S([(
����Ф4�!�Մ+ p�4Cz�ט�I����<>"��Wf�<8R69,����=��[��<�Llz" 8q�L6ө�3���&���G��@�EFǔ9��:�}y!��
|�:&ٮ�����k�������GN��t�ktZw^�+;�o��z�T�!K��˩�J��Z�]g�^v�\����4�hz�n�r��y�[�t�{�{�$��}cZ��Ww z��Ej�ob��F����9���}��,�0�Z픊��r�w~	��n>�R2Ż�hU�׋���PV��}lw'���۴���ՔSf��v��{淽5�l=�ԁ�c�s�"=�v���3��ӡ֚���f�5��_G���yN��i��_Y�r�KV�k4�S?fo�g�>K���!��"�4�@�ظ��
��a�Ù���tU�5Q>#���ee՜�i'��\l1M�+�p�b� +<*���fg��U�ŧ��G�u��lݛ˩mx���}�ay�Y�y�q��V�3�a��j��j�{
b�f����-r�eeZ�3������TǗ9˻���Sn}��$�H����]\�V���JҶ��q��_G��A�VH�t>t]$7r,�~�?4׼`��":c�� (1��S��7,81���뿁���"���?
�fi
���� �z�M�Ar��CY���w����}Ʌ�\HQB��Al�hФ>��ѶlVQ��N74a��1W�C�0A�8�1��ww�ldy&:�{\�ǵ���ة�K�{�#<�">�;�e�k���AG�
��z�i��xAH�C�+,�>f���۞n���O�Zk��]K��xr�����Y�X����m��J}e��l��E�d���9���%��G4#Ձ�L���5<�ϵo���7]O����7��qۧ稧�_��f���W������_ׂ��8��
���J�
��V�������>9�:�>s��[ǭ���ǌ�W�]�l��(�ר�*n�_4ͼ�K{]�ﶼ�Cl�g9��Ux[4a�H�] =Ef�]@���G8u
���·��oƛI�w����+�i�)��k)IN[�u7u�9LW��V�_`ʜ�^4�(Q�*<�T `ŷ��(d�@�u;n�#MD*�^��^4J�-�mj�Q&��vV�6j�CHA%K�����bU�����w�԰�5�Rz�%5+�b��è���^�����fS�du��o^�E+y)������?����[ǉ��u�h*ۉ�����r�>;ku�	����g���.���u�0|��S��x�?l#��t]��!Y��L���P�u��Q�9}��Q���+��g��>q7Yb�w?�u�Xz���������r���Z1U6P��s<uz���`b�����^��.��
��3��� ��(Ѻ˗.|w��蔶W��_�tk���m�lz�ۦ*��y�o�ﯾ��X��Q�u6͉߫�ҙLj�˞�e��g/��.����&�V�S�O)�����N-��{�n���z��.d�,�o�w�)��:�+ӧ%LX~W](1���4c��Y+8����U��P��G]��M���1Xj��xx(0��Q����NA�uP�����W_�M��͉��
/�v�J�Mbζz�Y[U�������w��E�@Qq��D88t8�{<������ңL�"`��r'%@.�S[��:bS��d' � ��.r*&=��\�1�����4�[)s���M�F�#Z5�9��G�X���۹f��� W��tĿ���tcƍJ0!6���"�wW
��BMzxTT��o{ۘ.#B�a�D�OwX���IKht�-��J�}�2�F�k�5U�6^ܸ��|s�Ϲf}Y�
|���n*��st��8v��c~���OyV�h�+�]�#�)�

P�e�[�ZvN��<�k�R&=�A�VeD�4'�[O� -4�~A�����GMyO#����jm�~�h����7�7eS��l4ƽ7ǀ� 8��"�J��"3�F:��u�_z�{�U�0��/�_��+T���Q'�����r��~��~��PMK4t�h�o�}�5����*3]�ԉ�b`DuYc��*�<y0;��wG��f��yZN	M���V��Ҕ�Y�f�S��� ��/h`ڔH�Ul��I�$�%JU���-醬��V�s/�#��E���nH����чA�0���z��V�$}��(��Ђn�o�4Bbة{r���GЈ�8%�M�x�x��hj�6'�r�{�b��K��3:��[4��@W�5��z�E���ٌ��>�)�.�o��4�N&^��ݙ9���o�v���O6�+�iI�p�;>͜��SL����0x��C!���6�;,0�gc3���P�>�2Q�f��]_�ʡc���H?c����j��J]�N&�K�㣼��Gj���-��8���A��T��L��Zl�2�B�A���^ކ�;��y1���,�j�S��=�*�������\�*�tib��%՟���{�������Y�~U�En��L%9o��Y���[������p)�У )�P��p�|i�^,f�,=W��`K?p���Vo�O8����@�T��W��+3�Hp1oo�{t��Dx?Y5�4}�x��kY�p���^�����V��L!uj�3M*}�����^^��;�-y�"���]+���e��}ﱹ���e|4��]ǅ�"��m�}�׺�)ˤ }����Y�AY���VjVx�j!
��®�(`��x��p�|7��C��-��������T,���G_D����K0 լ�/U��W��Һ�iޡ��fB��bi�.��غ�.�is�[�V�E�a*q,��^󧛸���uDh�_5t���5l��������Xw_V,9�����)����B\�zq��j�,����ر�*{�
4r�*j�]�B�� �V{�i�S:�woy!b�C/�>�]�+�]�$��ԫ��U����E1�ĦYr�.ɝX"��3X/(e��'us�g6�痊o�T6Q[����f��M���[�����\l&��%��ĝ�>z����W��׳$8�	@H���>c���G���9o�qa���9���d*Tm�5��(�l��|.w=*mt�	?�:E=�oA��X`�ܽɷ݇&vBpF_�pB�z���X3�9�͖�îv�|(��#�e���Z�;��3U�2�C��w�.wVdLLZ�!]���(d-u�y�n	�WM�M�"�����pS�*��y,��ks��k�]lJ�S���	%8�[!��ܳ��ٿL��o�vS%���ƞ|���R]�$��$�}���q�)�����i���]i��E���"ŋ��P�)UEm��O�*�t
Jb��*�ETqE2f��Qp�Ha���n��������EUH��!�Uj�[B����aiB#2�j��M �EX����f�fX�iH1����p�*���}���˛}7*�Tу)�k?pT�[S�����!E)�tD�0yO<��8���0%"c"-�ղ�2(p�.�y�g��^����`�P����Y��+�,/U��>i��eQ���{�6��)����i���;so�l1Zg��x0�@�Hm�����v0��j�Ӻ����Wk�1I�3=8f�5��<\�dLh��+���p_T��%A*-��"��os+*�����b��ߢ,1]S�����P6e��]6����G���V\笱3���P�=��
c�������Z�eG���s �Al����0s��ٽ�r�\ym�k��[��s6��Z������[�>7N��뮿1�)p�w��Aٱ{2~H�JPu�@+T� '*q�2j�*�&S%��>p"����`��8<�:��g>ְy﨡˗��MWl���:�l�o�<�\k�ׂ)N��j�8O����Y,A�F�Nݱt���Ш]��O���;�P��Ƣ2�Lx�=�1 �5�2a�X*2�	�;@�����r�&�
���v�'��g�ko���b����7�~��U�ozr�n��z���w�/�}�<���V�Ɯj+8�BU����d�sX��<�8Ԁ�h�ײއ]�	U*�PF9�ԢV�n����|N�����c�qQ��x��Д��FyX�0ʩ���wׇLn�7�Y�ۄ	�5���5�w�����.�2�?B႘�>"��E/FV��älU�4Sd�[uF�c8�PQ��jKm
��Dz;i�GE���^�T���a�:����}�4b�x���F��B��=ISٽ�+oE1Y��0�P��#Q��V��{z�Qg�C^8e��K��N&�\p�q'��:�\k.
�P�kI�qѣ¸G�9�~��k��]��'[e�5��ֻA��Q�笿x}xл���y�n�'�Q��}gnF0i;Q�Of�Vb����t�kC����XQ_ꪫ��N��.5����Qc�ϓO�tq�ǟ1��y����d��H��N|C��sPv�q�[�E;f���#=F�V��:�ye���������U�*OO�:/�v*���Wlf������08�ẽ ؜�"2%��}��=0;n�2�][Jy�A�>��LR�%b��s�ڨ*a��CA_/��&���.�G�@ЗyW�o��P*dTS�!�q�A�	�Y&ν��9TP駮j�F�˷�cU���ߛ��{׻���9�;ef��\=m:�����>�l���Z%�y�7yQu{>���|��b�4�]uf���= �{�@s`��.�R=;�؝W-�#�����=�km!ߜ��?����֑L�L��gYi���4�3Rӽ�A+7��N�4�8�����-&��+�׺�ަ~�R���C��w-�3�B�^U�3�n���r����E��O��*�������iQ��1�	�slk|�ud��1R��}n�T�)C�\����{�evm�������h�V vP�������z�mM;r��T{�8��5�v�R�9�kF1��U�
�GEǜD*4%K��8W^'r�G*n��]{��<���U�:GT-����ٻR�[oBo/5�h��F�'�w�=R���]Z�.�/tB'&\8n��xo�i|X��ogwZn7�Kx����X��u��d{	��٨�W![�kx��>>����b�-���j�4t}5ֈ�v�c��2�����ӈ�N���_9��xg��6ӱ��f���V��#D�o��p�m��k�[��ZtW#Z5�ѡZ��[��A�+Y�n]xt4j�9i��zͺ�i�k�=����7��e4�_^\E91p`�P�{�<��ȸ����@R�S���`R�c�S-\�;4ٌ�̡b�$�*�>����/r�i�j]Y, �SNذ�!Ⴂ��
t����%��z���_9`�\���W��F��o6L�[�x���3�n��gr�n��=�	<��f\3�o�W\�f�&�g4��O��u松}g,-�z�f�ptv�]
=�]�x_s;g����tm�mz��i6<_g����������t5��u�5w�W��m`F<�U��_]�ں���%�w��M�hV�r��`���+ktq���8�r�Jr¼U���wݶ4V�ÂCQB�5��CRw�95�'�'f���}i��\M�*�p���n���~�%6�z��ۇO�����~�o��:o���օ;�Rc����lS�PUė����a���`�.j�f�P�.�V_�]@�/,��ۑG�I�`AU��ˏ�������g>���W×�<�n��0UlgS;��Ӌ��ѹ�!�F�^ ��Ș�uQ�ټ���@ȧ 9��*��"=�7���9��.6�uNC�Rcr}Q��vԵ�*"��vG-�w},�[=u��jΥa��foM���{9��xg�X�h�}�p���n��z}|Lrky���2���.Yb{U8��/��)�u�z��.�7N�|����÷N^#��-Fx�xS�VIB�M1l�H@�)���=��]���,]~~2���n�G]a�e���A.Rwu�v���rF5/,�����+�:�V�:ޏk�궭:ؒ�r�~U���]|�v�_���>s��~5PV�{L��M��Q����t	4n����ƕ�¸z{�4����w�WB�U����7W@VE e@��/��2m(1鉀*:<��Mm8m5��{= fu(����mΆ�5�/Gٕ� ����Z�W��XfZ�(T͋�����z����I�/%�N�a��݆��H::Z.	�[�����wY��:�hN��M�~:5A�!����r���+ȼ�g�P��m#F�//�vÿ�Ԕ(_��������y{ȹ�i�i�|�^<�z�_r] �0�n�}}\hN�@��(3{�����a���Y�m�.p�5 �m�;�C��|��G�|<TMt?0�w+�S渲��;�r��i�N�{�+�p��N��}�A-��[�����b��
�W]Ґ�bp|6β����!@�S��cbb�WH0	޷�z��s!�ӋR'�سɇw�`�*k�y�߯�֌6�Ҽ�J������D���"�<}(���Of;%��@l�r��&D�ǆ9�-�xֳ��Ez��|���'S/�G��e���P�:�%̑@|��~���E>�r��i�b���ڼ3��I-�j��a���U;��L�,O�Yh9�M��^NOGt`�4L��^�Ǚ��\C!R�qà�<�C�E�h[o�a�Y`�+���q��ǜ:�,R�����{E���e���bqJ��:��"0gJ�F�[�=9G$dbCb���t����U/0�ʚ�ۤ����L��R�s^�I�l|���bKN�e��B&��I�|����6�]z`�c�ϯ{�u��¾�A�[�ְp��G!�wt:|���7��Gx���6��{6����R��S�/N�K;0(s�)�f��.|�?�Uo�����+]09��!)�u7��u� s-\���o
qQaua�%2o�K��� �-13o�B�;ݼ�v�jp�t���w5���@q¦V�\8gZ|>�<��0�8��^���)+
F&Y��a�[XD�ά��ൻg-[���ۨ�v^�A1������ȗW.�I[�f�|�A�Q�;y��o+q-�'�t�����j;�ђ�˄1�ۙW��{3�s`c����Q�$��$rg�E�RP��T"(��H�J�Li�# �S)��@��Ĉ�4�������Gm��EF�U*�,uTU�(`�U
7EE�Mؔ%U.(�P��M+��Ab�*�U%]R�J��ZTb�Uj����p�VSJ�����tSu)*���*�MT�4T⭖R+B��X�c�B%4�J�)ATAQD�3����(�Ki��_}��j7�t�SwP���h�Ε�	����%x��@�ٟ���]�Dt�2���]+�SL��m!Yg���K���Ej�T,0��w���׫�+�t���&<b��@� ����-و��{#&\Q0�wI��6S��sQ#}�]ً�
��o�b�]J���Q�/��ޛ`U�ў4jE���ߜ�'B�uo�r.&C�Oq��;P�9���+�0�Ҽ�E������v���k7߻�������.��v,�ب��Qx�X��fh�B=�3tN{��J�<��������:��8J�EVw,��}y�z�t/����F������<䇟z)��D������3#��fV�z�#���r��[;�qv��q/�xS��S�J�u�������+���\|nP]0x�{[��m6�??|�g'�/��5u��w�U���ex��4{��p�l��4���>|�g���5��i�����m�
�����^�ސjT��)�%��vw����>wgcj��X�v���Ӊ���x�u�v+���H���
E�O|���;!n��a��e%����r�R��γ�G��9V��Z�8�0͎�%�އ�4�7�OtlA�z��ݻ��}x�׳a�1D����ݛ��~h��� \T<.Mm��\���N�"6���8L1�����{����u�~7��#�?q^�5�s[ژqK��s^��%%���ץkݱM�T�t7e�tx��2�ɽ���Nn�޷��c����~�?t�-�+0�d~�u�K�ɽd���w�[��u8w��:�L�!J�G ���v��+yυ�O*dnط��X�/���g����*�<��[�Fu�]�{H���Icƶ��������)��Ʒ=X>k��eJ^��t� 3ʽJ���Y���ݫ�:��}�;�e?+AA��]mZ����+؇kp��U�t����7��jf�筘$u�X�8���!ַ���rvu�UR�tI������JS��l�V�[oWأ��}/���}��[� Gi�6����{��
���5աeON<���ԝ�=}j�Q��n�;���A⦜��;Ѱ��mji��b�,��g`E�����cg�.w�A�&���沪ۙ\3Y�B!��`��\�-�kV�f�@���\���m|��M����zv����G�@^��Ҋ�z���{����sx|�w��U�)�\X*1[Ȗ����}OG� ���(�j��D��C��޾���~�M�/��U�$�EOW�>B��,ܝ+Y���[� �+�S�g���e�Yrj�I�o�gOs�	4�^t��=�<��qPl�C&�^��~=ޛ�M��j����:�yn25����}M���F��w<�
;��{���DI�j�iMΔ��B9Y�WV�\�;~�.�o�����(MNQ���Vw��F���ʲh�܉~��,�ş�����ef�7��ԟ�cZy^N��y*�P���I6�.g(�+ke;�n��[X���P�+�;`^����iV���^�\������o@�4���6��lqT�ވ5�b%�=��:{�Y��^l_7�OM]'�]�ƛq�ّ2��M�pã�c)�l��3'�-�6�`���r�f�gMT:�-Ťzl�ḯ�v�!,�[6�a��N��8�������t���]��뿀�k4��[��!�'��}�R}ٵ�ٚũ�ԗ�e
0V7�}���)	}�+XѸi��7��w��V����[��n�n1r4�珅��3`��v:^6'OC����뤊��q_�>����&b����#L�m����7���x�v߻�3�|� 4:iP����|dK�X����y��g*x�V}���C>�5���H�ٔ'a�u]â�JS��|F������W`��7�
�{��X�2�e�ѡvu-��\�Y�2�-�1i:\Q���=r�1�_�=t����s:�9�9�}cR؏D�ϬΚ���-���X�I�T��-vw�n8���v����GM����[�;��G+G��A�ٗ��,O��,>��/!᭡H2v隓g�b`ܤ���C��?v�8�.ǻo��%��ג3�#Y�!���r�<]��{�Z�;�ݚ;���T�I�0g�>��{N� �T�B��G;q^6�sY=3�}8$��b��%���Z��<����"�ז���dV^�f��#e��{��G#�4���(�Ȏ��h�y�i�����x�l�p�,���tг�}�+3D; 7}�6��] 5�Sl�����6��V(z�6�rtf<�5Yg��e���	g�������yR�#u>���uA��:�Ε���0�ݺ�*ߍmn^8�o ��j.�a��]�7���⩖N���̩6E-�	YI�Zw+7j�����Fv�k�6��9���n8����u�U�������Z�Rǰ����P�u�2�0�M���Α�=Z�NiYe�Y+C�w�2�[�Fj�������G��R@���L�9�ɦ�w��DŞ�� ��E!�ͷ�%��c��f�/��m��_m�jQ���zl�� �0�wo-���D�1�Cpj���{�e���{!J�T��e�J�\M��h��z�WY�r�5,x��bh��En��m��V�W���Ɨ-�u�uC�V�}�rj��m����7\����%_lu!Γ�vq�qN�ռ(9�8@�]�#cyj�o�=��m���ˬǎa/;YV���t�԰���bN���e�T�S�7��8�;Wy�l�.�JV.�ܫ� �Y�-�B%;�t�[	f�d��{[c�&�wt��2SY�pU>S��M��8��c)�b%%fu"�lscqtrI"�I=)
� 4@� �EG�,�"�E{T+�AF*�p�ň�*ƨ�R
�VD{A@�Q�9�B.��DQ���+Jj�wv�J���ꑈ��eQ�)F1Z�����Z�R�Dc�U"������T�iCcEUE��c1T�-�SJ�顊",AU�T*E��TP�աuR���)��fG݇�K7ͽ%Fk�s�=9\��W��;�}������j��n��b�=yI�`s��/� _{WS��8+ �6+����+}�9^���gK}���jsٽ��2�M���ʯ��76t��(�t��]���\y=�ž�r��]t��K��[۝ۅ���W@�-n�n579��x4��n��آ0k��������ʦ��X�:>�Ư���k<^�M�a�˦zc����q��g���-�R�8Xu9���>tS
��KxD��w�&�����;�UX�dV�oL1*�jJ�7��Ǘ�fe;��5}��f�\j-�[9����\DmMrU¨�x��^��p��֦�R+} ���y<�z?hԾ\+�f3�pqvBw�̠"��qe�]#޻�gL���xm܍�%��x�'�����qoEa�NoA�V�d�ᵞ��3	c\�5�h��?<��K��ݭ�'f�;q�S!���~
��3�"��I
���7�8ߜ�z������-����X�j��/�o���;��j���b���L�������4ɴ&�����٥���V[��ܙ�ߺ�7f6�S�⺝NWz�ilY5��&p������C�����YSڼJ�-zC�pJk��r{�6>]��8����h��N�k�p�P�Wd��:X���x���92j�`ټ�U!���׌�}���}�]5�Ws�֡�(��OwF^_���԰Z��N<W[�:�W�! ��/�����ڔ�:��F��	��Bճ�W�$�c���"|v�N���B�4gt_�e�w��;8KR���Z����s0ٷ���1��{�8)@˗!�h�P#9�4����p3���W������C�،�Qתv]+L����x��sE�K9��/��ei��'�=N�8%�����B�����/�Y��{�ٜ����Q]�����W�H:�ջ;Ks.�5��uˋ��zH���W�t��"O:�;k��-b�y��-�v�|T���{�7�?�o/^���4��UV�W��reF��	��c��-,�Q�vBN�w�t�إ֫5�tK��3q��ǥwt,�r."�/Y�݅6ZU}�L��m�x5˔Z�U�]��n�}ئ�f�.�uL�b��[N�y���O�#|UMi�O{��w�C����K���NC�;su�[�jkãE�ʞv��Q����Go9�۶K�y�S�;���;�n���'����!�h�i�{;�w����vU�b���v�潕j.w\�t��͒gR+$1w�.Y�%�z;�ѧ���
˾͕�cU�e`N�S��ϒ̃|~^I_��˞X��*���<�S�����R��x$�
2�$;�:���]��E��=��7z&��3���G��D`��ך��G���S��m��\��W�^n�,u�R�,J=~�QYro:.Ug5Gq��8:^�����r b�s�¥�(���N�S+D_`I���s=n
2o�;+;/�Jl�/��B��������<5�7ѫԚ��̧#���Z3���.�g�	3������8q7i�̬�Fe�, ��&G���dmܹW��+<�U�ɝ����TVm�	�>���/>Ȭ7/;|
�feE����vQ��sqQ,�.��꭮e_^��ĵm��㧦���Xv+��yb��hk%j����#���>Q{�1V������ߒ�@i�V���v�������Hܪ+R����~�{_G窬��銏��"3Kqu�TxE]G��R����E��1ﵩ�Dx�(>ul:�q�]����$Ie�7f|�ɋ���%�\��Ǯh�n�&���F��v����+P��&�ًg���q����ک�l׻:�x4��j�$��_΅f��-K�R.Ʋ�V��*�ʷxggws��t������T���W:�;,ԡnY���u&M=���~B�f���X�i�e&{�T�nm\E��z��	o��z�f��!E��r����z�;J�&��7��/2��l_,����\����3 OC�aȥ��t�jua��6�z���_�#�u���F�Ȝ�K���7?\>���&��p<w���͉cx�4<�x6��ۣp�z��P���-�]�g�Do���վ�bG����{7/�92�G�o{�R[Y�|u��dj���5l�=T+v5nj��i�]����M���& ��}ɌR�O3b'��M[76������o�i�6X�+�춲ػ]|���x�Z��bۚp�9����mʗ@7Q!qR��Z�+;���
[�t�X�� �]*�i�j���b��{Euڗ�]��1����B�R����2 ���oi*�G0˨4�b�+8Wc�����oх��8�v��-�Yε�^e���9,O���,�[I޵Ζa�SY#�]g�����бeӷR�Vv7�6�Q���yǫ�r�r��ө#fu�B��\�;'c�<���r<�8�w��ӣn��	M�&͊�}��c�y�5�vm�N��DJu%���Q��x�^�(˔�t�yŎ�:ՖNnl1��(�=�c �.���#6<��,=���fN���_:ɯ7!to������ad0�<�c	�3.�J}���t�w������p䢾���\/V7w�J`�Q��r�gM�-�8�R��.Y�ĵF�<k�&+�nWk���	u�SM���7֕XY%�������,��o�E�xsPj�R��%MΚkV_;�0sC^q�om#��j��C{}��+��չ̓��O���Jb�|��Ȍ�q���;o������$�I$hT(P���ł���T�)��M��Qz��
�0X#
D
'Z#��H�TA�JU�"�ZEQ#"1U`�1�+W4P�Q
����R�*�Aa��#DV���F"��fZDYԦ"����YtVZP3E(��Ep�1`�,�`
*��=�5�o�?Zo_�tY/����]�����|�o�+}�������Վ�#��7ϻ]�b]v�h;*/��8�c&)^��]c�]�r!�FҠII�G�K��^5��� ��'� *ߋ���O?KwS-,�ء�������sU�o4%˷�6��n��O>�^�喴�<6S�8�&H��|6b�CY��B�x>��y`8�	�A3�K$[�]�5��E��:�)J}n�OQ:-��l�����z�T�������طoϘ�p��Rx�ʡ�_�/� mA����[�y�;���f��]@�e�E�Q,Y��G7-�[Of�N�>Sn�}�t���}���¸�H�;�/j�)w$gX'��x˖�}��.��lvd4�<^R����V�cwf7;U��n�Z.QH�f�6*-����,s�����͟E���?��N"�t���0� ;�V<3+�D����|[�,G�^���@�5��>�;�Ӊ��4y#y_���M�i��L�\����Z���󸙙{:��#�dt1F������y^�썭ZY�^�s���DF��]���Rq����Iݽ��܄�7�������]�eK�[�|�k�(�]��!�D4^˅X��q�Um=�!Ȑ�&�3ʷ���Q��N�ܷ9ҫ�RL��&]�{��
 ����b;KJ[��C\h|���� �ᡔO�U��7]q�tF+�i�<��m�YO�Ol��d��������۳#�Uj<�E�gٯ0V�ы�\�P�1&���s�ٹX뮕O/nyrsP���5��Y���t稾���rU�9����K[2��5�O�5���ަ����X�0�o0���OӺ��&�a�t���2+އ��ey#��A�,��ZV�l}���l�k��*���N]��R�k|&�����}�F��M�S��q�j¯+x#�)wu�ڝn<��]�q��{kt2��Yy�����㢇)e��z{I�iV�d���6!U��Ȏ�WB�ڸ�qP2y��l*�F ֒/ܺ�蝀��\P+Z�'��]Z�|�G��@�p��,����z;x���zߘ���n�S5� u�۝�L���S8j�W+��Z��v̞[F����'��dײ�9�F�Q��X�-�a\�4���Y�E��oi�ǳ7B��e^�]3uws�Ԟ.N?R���3o�����z��gI�3��Чy[��+�Ǧ;{����鰎�%)����PxB���g�6�#k�+��g��
��N�ڑAΙ�����O�
����d���wl��{�B�ANQ
�&�O,HWd��<��`ʨu��Փw���wu,䷗��˭�&���{�3)H�ҧ*���|D"���p�̓�z�!+��w{�PëN,�X4/ �z�\ա�7��������͎�I�,x�O�l�U��\��\#����y<^"F����v�����^��\ʍ7�z�Q���n�M�Ž�Ӽ���F�׻���[�a.3mY�*��M[e����_J�o|��;�Q��zd�yp�V��B;��ݩ�����8�o`k�me��˗Uׇ�f�U
���n��/Rn���<���ÿl/md���&��^Mr��^[7�N�]�N�w�b�R:3ۗ�*H�:�{�^^S+��s�:���b����}�	T�V��d\o9ڽ�T�<��^Eu�U4.t��Ph�+{������Z��pd�m�ڥpw�u#Z'����n�b�v�%/4��|��a��A^��Ƿ�R�c���Xc.�aޔ�����B���{�jv�\7]ʬ�:#Bs����U=O
T��bX]�N����o��l��]�Aa,U�-R9���-2�u[�R�$=2�eĻ�Lȗ�K�5��K���_�n�/�[=5��o�f7"�4�gwt��a[�	0EK��|�X�Q<(�����x�0\�y���e��q�f��ǥ�m^��V���wjycR�d��v8�s���No�o��
[�յ�+��f��R'h'w���Q���`���O��Ϡ#�9G���s��q�r_��nV	�=�{Ԇ��K���g9��ʼB�ݽa�^Ku�=+�Ŕ�H���׏p�y;5�vvtz���Q�J�V%ז�jrZ�&�W�rx:���%(���I�;٧��3��H`x�P����K��vsw*#��k�m"g�}����2�mr2��G=;UȺoh�ذ��:���ȶ�ՁG��4E�p�m��x�v�c��㰙�9Ps�wXN�6w,(���û��Z?T�PY�jy�GV)"?���su������Nɦի�ηg��u�Wz��)��kX��D�Kib�o*��[�Rv����������d}ƙ7�����l�q���O8�uo��sq�C�i^.��ƻe�)(����`�f�lր��8�]�x�I�X�# ��٨�
�.텒%�6��(�Wj�ej�����*�gQۭk9a "�NCja޾�6Z��D�][�Mm+���.p���V�.��Z�e��9�u3R����㵭��|�uge9-.ʊsu��F�NV�3���s���7~CS[���RW�G[ע�yApknf;��8�澻�ew[�|oy�n0d��{��W<6K�,J�ѝ����m3(�/H�Rv�V����R+L�4�0�ޫ���n�V�?.G(��JK����,���<�Q�ܑuJj<Ra딖M��e�&�L�
\ԹYFX�z'u��ݽ*�Y�Hn�Ǫ hZ�1��t��ݫmp��t��!�9�N�@[��Ǚw]J�إ�,��ޢ�9�n8��:9$�I$��_�T,�Y�~��v�dUU	���$YTP�u)UKJUrҌW,)TA�"��*���E��h�#�H��J+ULT\�%����F���X�,ë��@Y���D�RR,��SUK��0���d���E�ET�U�&,,QA[�L���:o�~v�w��-���h){�VN�5�ֹY����W�U�I�zEec�:�BȦ�u������vs���>�dY�*��qWR�On�22te+]�Y܋M�NR*�V��I���7=�7�uQ#GY\�O\sf[�����3ع�b5���ȋ�"�Iz���KD�y1n/T�Wr:1�4�G=�m�C}8^i�&
2y�a���׳�T�t�H��_l�B]b+5U��)�|],5(밟���s9�-�ye&&N͇VG��+F��G��������\�@�|x~Vb������\N�v��Y�@�9ݶ�����!�F����[��)i�I�~s]�E8eY{�Vgx=��#��d��Z������"�j%�s�%%�,o˾���,��cf��
E�Db�O!�u͵~~�>/��qey��S���Y�wu�o7ҭ�:ƪQ{o@��y�f�ًr`�N]G�����{�ofk���j�]_lW[��jԵ��c���^g���D�u�-�z�gV��]m�lWd���W���T(�{$��a�χS��yɻ��s8s�r�=cl���El;��s+jtf������nf�v軣*�/A3����:�o[��b��Y�62�U��(e�E�}:�ʄ�7�0��x�L���lЃȸJ��a��d��1v6�;Q���?y�Ú�z���m�$�)u�y�/�c�ݪfEY=��,F1Z7�]��aG<�<Vd�z�*� T��P�D�ڜc��A�=��'�������̶��oQ��oCkrn��B��d*�z������$Ѿ������כ�T��4����$Z+F���O&ɮ�y��3���>�㏜^s'82*OuU*<�(���ɭʖf�j`e�J�\�_;W�Up���#oQ��ݽ'�2���4�v&�GZ��X�m�ܭ���-�.v>��[O�ZB�9��9{����ym��si���H��nK�i+��Cc����ܻ�jO0��Sƚ=��d�V���7�cw�>^OR��pi�����Y'Cls�񃷽f�i����뫫!��u&�OR���\)�M�6}��5&��s�P�8_��wS�!F3�9�Qu�!eSo	��|�/��ӣ�oro�h��g��ղf��w�~�[y~W��j�FEu&�c�f`rZ�y+S�g)�����9yP�r��V�Z��5��/��f1��_��^���+{q���1h��e�>��;K�w��oݧ������f�Q����w7S�R�dCݱ�@�##0{"�9�%��w���V�v�ۏ���=eNLs�q�T>7��"B���Q��S�+�ݒi���yg�T�?+�]ǆx�W�E`�\+�U�:�ua��ƒ�(�SE�)���Y+)�]oel<9���ܷ��n/b87���U2�y����ά%Y���yk]�NуZd�������U�Y�6�95���[�8d�>9.�7��� sޏ�+5v�ܦ}ڻ�������g��)ѓ�p�E	�gw۩{K��'l�C��or�Kol`�99R�2ZX^LΩ��Y��G˳��!���Sz�HM����_I}te=>��-ɴθ2^�˭z���S�e��͓S�vc���M]�������޳N$oO�H�4���~]��l{A��{��f���͛�W���!�vս�	"�n�|��&�#X�i��z�s�� z_$G�.if�^2n�1|�Ҹ�&-�'���R��Ooon(�:q��-L�b�n{���K:��2������9~r���>o��/j3��O�O1�؂�q�Q0�y�����T�_4���яi�ͷ��}ѫȍ���)��u���v	{�]Ϟ���n�7~���2�ܩ�F���A]/�j�>�2gqQp��E�_3��8��U��zn�fn2;g2F�9�Dn�(겸ͩ��X#�t��nN��Vқ̓��ùm,۾��W�n�p���N�"����F�AO!�&��u�����>�3wȬ�XQ�b�0���mh�oE�z�t!Х>[d�9�m	��VC��I�9!��\�N��{�N����]J&�?z*L��=�zl���j��nG�=�
��
ݥk$��SyR�ƚ�H�7Uz��&(���"���&�v-�b��WYKOf�z?oM3���U���{�-����+󞠋��d�;���շ�������,����	Ev�cgqW��F�(�l�V��O�}�����*~SJ�AU���$����"�����t��$����F��
�W/u�1���C�0,:1�<'R�P� �RI	"�w��/;.d�L�
�n�aP>�&���?�2���J~��3¤�T?����$��/��	��~�g��]|�!�������5&L�߁�xD/�����._��MN�Zܛ�a@6X|�2��~$�$��؇��������'k��D�`��@�C���d!	$?��%��>��\~�>������~��%�����B�������~!��4~��B@�C���ʿ����H���2�2I������ܰ�k���d���Q��B��B���"�>��C�?6D6�?��a�ZԻ��$��J! I �>�%OD��Յ?�y0B@�C������N��R4J�Pd>�`U��C�sf}��}_	�s����T����Y(����	����}}g�?�!�U��~ʝ&C��a�O�C?	�O���������G��5�:>�Ȍ�II�d���}���>�G�C��?/����h�Q����_mO@�
�?��+���������>�2����?�>���������a����?2�X�ȃϿ�?QC��L��!��� �=�C��
U!��BHI �XQ	I���	�rr�j-��?�(>�$���PH}F@?�U��$��h���	<����3����HI!Pd�Rd�$>��I�1��{�0��I(��Oh"B�ԩ�`$��D;6r`�_���ƂHHzXQ�������!��$�p�?a'�$�}����?TI���	����O��'�����}d�HXH~��t�CG�OԈX���	���=�0�0�$%��}����C��yD$	$?��n~��~����QD����!�?�B@�B��9~�y,�@��?��>���>'�C�>�%�Q���������ҌD,%����>�?�� ~������C�����O���.'O�g����D$	$/��H}�5~P���������#	�v'���	��X~(C�Q��U�p�@(?�2H~ϐ���@�C�!'�?����u	��s�3��G���$	$?)?��M�C���&�9���9��ہ�wy5!�Ab �?('��H~��	�훟���"�(H�v 