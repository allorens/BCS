BZh91AY&SY��j׈_�@q���"� ����bH8�    oz     P QC�    � AJ    P         �
  �!A���*� )T��E�(

 �)@U
P(P�"�P��A B�� J
O�
�

  	((  ��*�� 
)* ��� �(�Q@U P(B�  �d
(��HD   �g�@�i� ��r ��t�T k��h 1P4*�R� �@�9�$ )ET��R��  =  `l��E cS �����P(+Y*U)�X��h�`P��F�@����T����� ��T��� AT(�x   X�xP 
�G��t(�o��4�Fi_{�ү`��{��AA^j��� )A᫽�P y�� Р�7.(�P�+�P 4JP
(��( S� n�a҂C�#.��B�Tj����2�k
�J1��h�j&Mj j}��iAB1` F�V �(TʵR�U����@
�
 ��>   ���
�P9��@+1L�T��T�ѡ��5H�P���d��K���f*�U(YV "}� tH � ҇�  ���@�� )T	��"�P06(hP�L$S��-@�R��V��d�� D�i�50(յ냠  �P��  8� MB��T���40� R�X �2�hUR�)�(�XՑ*@FMI
�3E�P�}p� PR�(��   -N�RA�X�IUaX��� ���T��Ƭ
�����
���DE��
��j����ۅ PF�J�("���  ��*Uc+
E�-E��9*UQa���UP)eZ��T�J�*�EL-T �������)@
�� �o�  _U)�j�QUd�U
�i`BԘQA ֪�Vzn�UEU��TF��B���	(��    
� 50T�PF  A�	� S�Ĕ�R M4h  b)�DM0Q�O4��6���$f��%I@      EOޣ@�I  L 	�J�gꤔ      �y�τE{N�/,i�ٶp_$���_J�q��c�L�1�/�A�Δ)���� �r� � (*o@x�
� �y��S���_Ǒ����� Z�"""#k� {�@�!,@�a.B"�+���׭�*��
=�
�a��p���	�%�A��|�?2�̩�*|ʟ2��)�)�2�0���
y�>eO�S���~d��!�
|�?0�)�0�̣�
|ʟ2���e��>a�G�A�e�G�Q��~a�_�S�Q��~e�W��0/������"�ʿ0/̂|�̃����	�~`_����~a��A��?l�2��� ��?0̃� �2��!���T���_����?�D��~e���>e�'̃�S���~e����>eO���̉�"s*|0�̉�"|ȟ2'�	� ���O�2'�#� �ʟ2'̃�
2̉�`��~e`_����~d_�@������+�
��?2��*�ȿ2�`~`�U��~`� >e_����ȿ0/0���*�ȿ0/���~`���~e_��d_�	�>d�U��~`�E��~`?�D�����2)�
0�e�A��`Ty�Q�� <�2�2*?2�?0
�2��0��0 ̠�� ��E��Q�DG��D�G�EG�E�TG�PG��U�Q�UfA�T�U� W�PG�@�P ����E������Y�>`@�U_����~e��Q��~c�U�P���G���~a_�W�U���� |ʹ�~d�U��~e�G���~e?l/�#�/�������/��_[�x���p���Q�m�H8�tޅ�-ۭ��J�-�z�0I��HB�8D�зj��8��Ͷ�ۖ Av�1���E�!O6e3����X5�;Yxw�t�l���G6�=xq]+,�iK�D@��){���&e�����I�t�M�8�1]9[z�8�H6J;�^SJ��cv�d'	�2�l%��V�a%YZ��&�b��=x���h�o_v�b��r����<ѕ�u*S�~ToB9��35��]�.�d�l!i�U�2�N�x,^��U����.龍�RN�g^��2^6� �Q�{{3Q���,�;�Lɭl��v��w5XWKm��n����S����6�����6ѳ��\��@R�^�;Rk0�p� *V���Ȗ�U���0rB�^n(�.��ي��iá*�,����OmS�6��y�$bR��-���K���z�jv�α�Ш�<�U��u-�e
 U�[��@�mPg(m�ɠi�mm�Z��퇮1�6��V�,Mmf���y��M;�~׺�[�P���v&֥XF�u�A�ceajӮ�ϰV�r��ۣmQ�N��U�W���zwdY���P��f��[+�Ք�u�����^��#VY�w�R41T��C���H(�� ���u�,1-֠�ݕ2"U�Mg&�#�TTͭn6���sS��i^x�׎^���=��y�*�D�ܲ]o7N,�q�f���U�fbܣ��kn�ب�l��N7t�Xt��e�V�Ksu#Ya��#��M���$�E�����2�Q،R��!��e"�[�e���Wj;�U�T�)�� �9Q[��VX۰fn�*ΗI�csp�/(�{3\>����lj:��.Tc ŻP�l@�2R0��^�bc�F�
�Y*��q�x�o��;���¤"4�z1�'��]���Ҷ�ôj�\�Z!��*���b�ɂ�ʉ�y,�RU��U��;s6�
J�b�]��/n�g�{��Kneh�,��wWd��I�BY�N9
�HܓEaj���y�1X�wZ��BH#�j+L���iwZU@9Qњ�Zђ�ر�&��i�%�Il�o7���x�fn���v�z�֢�d%Q�6���JU�A��89=�n�b�e�0��H���i{WR�մ��� #�p�s�G7r	@]Y������2�9Eߴn�IS�����Щ@(Ǥk���{i�l8l�h��t��LJt.��M�6�j��k�2�R:��o*a5�`��Q��e�J̔ޜ���:��9�DVCz^��Sa�Z�r%Q'w���
<#D�nm�`~a�W*J������Ƌ�^ҋ�Jh�PB˕s4��4�9"�D��zt��̤�-�{�)nU�]�[����,b���J��׆�e�I�8ͭ�V�l�u����f�Enn��GD���t����yM�
�$ܢ�Z'�u��BY��G�e�6Ě��ЀB!&��O+ r!=k&�GJۄ��S+J�S�4�z�z���c�t��QT(��Wo`�bl-���lP=��Y�pһ�K���q4���]!��.��0��V�͏mm����V�tJ�o4�x�&���X	����ٺ�"�Z���KlfŚVf�w����iM��U�r��e��J2a�oG��V���ͭ����zH
��]5-Pd�{��RN�w�M�2]4�Rm\`��xn�\����4�$EJ`:��"�LN�w��ˊڬ�n�� ����r;j��v��EknS����Ӹ�77vZE��l������on��n@��"����D�)YZ\�V]�L�S[�<���(��ΓyY���Q��7S(�,Z��7�6ok�k4`�E{�ޗ��̿I��n,$�&L�V=���\��&+�E��^�ڶ3�u.�XB����8,.Y�;�e@3*��^�60e�f:B�ҫvv��6ԣ�77&ͣa�V�m�ٻ-Y�կ3FMv.�X�a?6v��{��`�v��4�Ĕq
T7Bl��b8JXp͢�q���D��^��T�[eL�x�� �UaڭL�jԫ�sH,�x��N�1V43���Cz���Ή�2"��F�۱���N��M�x�l�jQ�fe���&��Sq��e
y�Y8�OT�a!��7" �z�!�񆡧��6��L�IZ��1��/�Hז.�휘��ʒip�l��#V���̠�9z'���t�ڼ�hmJ�
��afٶ��zB�^�x[�C���&T�)e��Q� Z�0�O��2�\m�si2/e��ux]n<zp8�)Gn�K��Re��A��%{��Ib��64���NZ�f�2n���0š+e�Z&:��v��ҦH3r�Ж66��,��V
�)l���	fj/��sS̷z�ڧ7wI�	�WR�-�J֥�)�f@v���2\�hi�ۭ$����z=©d�gw-���7N��"�.�&�X���ݷ���x���R;��*�lIiˀ�d�OH�Z�N�����(a�Zf�TrS@�KN�W��ɣ;�jX'\hwJǍ]��:zk�m�gFX�e�7]���#@�6�hS�2�Q�Ƒ9wW[[E��K]��2�J8D���%Cu�^m���8��p0�7Ct:8��(��ƫHn�Ê��y{{Uz�Lݡ=��	�w0/�T��nT{m������;@
���ChE�u)�v���j��D�eг��{3]��呗w����2�n��3r�0
E�]4����W��+/E��T�z���H�Eh��*�ՓS$�Ĵjf����y�p;��6��fA~N��n�:0��?m`y�Z�����ޜ�t�&�nmw24-iE\����JW��8E���+FݫL�lש+͂Z�å�ZOCz21���8�mjnsc���P�M�Oĉ����t$6,� �V=ӯ\�v���++kݕem�eJ���^�.�Pz(ZšHnѨ�H��F��4�c �4mb8�V�3n��V��u���/QN�<t!U��� SsE:�un�2�֦�V
�܂��h���V�hX�4�W%-�̩�vs,@�ExQ���X��v�=cm�hM��1X�R�7	�L�eဋ�F��Jiէ[o-d�Q��U���ei���%�ƅ&��*Z��0��{j��)M�tI�I�U����w2+�X2��Qni�,��./Dn�*��e���f=�L����q�u�v�=.K;n�	e�X�37FࡡP[4c�B���4m���69��^(&��0Mv�D�;��☦1�F��$㸖�N������VT۳J���#�!V��/.q����w�9��͙�X[x�	u�DM��U�	�E$��q�Q^�Z�hF��h�̧u�Z9wb�儷U�ڰ�ׅ��	�ж����V���h�Ҁ཭�=x��ֆ�dUZ��f7NR��`�U�'^�+h���d�/r1tkS��t3.�ƪ�@)�Ѵ��Mm�V��ea��᭡y<D�͢e
����B��+�1��+g�8��!��ͅ�FC#Z�bZ�2�A����'M%�Z��`u� �`�&�[�F�t�j���fcNM�u��AՊ�M���W�sn��4�I�\Q�΢�@��:�:t�[�����`����s$s\���,T+�Wj��Y���YR�^��jkFh͚���N�/iU�m��4X�Sۨ���q�,k4qd������r-�z���=b�6]Mi3;[yf�7p+�b�U�$�\j�W�4��Ce`��D�B�J�`��ۼ5�0�"�:]���Z,J{�R�oU݊�l�ʺOl�ѣ�\�ܵ�wCi�n� ��Ս%���dm�k�Z��+�z��hK��&���)ݳ[J�ZH�R��	MU�2�, ��/=����V4���¤4QD�e���5f'N�Nf[+̕��qڸ�<��W��+!���@m����n��V-��q��p[�:lT�-t)m�M��l+��XSf�H�aسr�єu� ��yB���E���c��V��+oY!AK+^��B��r�,��Zuf��n˰�i���[B�^.〺�mr�V� �r�nި���P��[)�vr���=�oĒ��q�HV��a��B�ˤ����Ѥj�%�0�Z�PȮ��&��{r]b��;���D��``L�C`�\�]trQ��!W4�9a��.��V,7�ICM���s�H�k5��Ѱ)��]���gr��^�T���m�F4�ѵ�È�o\�Tl�7Rx��,��)�
��f��M��g1,�Bmj�g�\��4h�N�Ɩ���ɷ�e ]���{%��`�]ZsT8�Sh^�M�,��Nj�o�p,J�s�7�!늮�����3fY/^�w4���W`Y�ܻ	�EACQ��^�ur��mTs2�.<Z�]��ʌ�'�ֽ���Ѯ�ɔ��s�#l=R{5ހv��9�P��ӎ�2�5[�na��`
�C��{o56�U֔��{Wst�Efx[�۽�m5�j����nhgr��]裮�8K�]X�Z+^��˕�(�K�X���NMiJ��&u�U��4�����ذ6�ܕ����Sa��v쪲6=vme�bKV:�Q�Y�̖weQ3n�-�^�l���!��c�2�����#���o2���n��f:Cw�5�N�6�v�ەudeMa]ͬN=��h��`���	� ���f�tX&��U2�^Y͡�؆�jPc�tY�%��6�iԑ�S�!ʖ�`�Y/5���)5*"Ajf"�B�gL�C�)�)G�s�w�2�I���S��wGwV��;0��P�����1r��`:�ɛn�f8�c��f"�zc��6%n#������0��G�T�9�,f�52���]^(*'5x�sjm��*�銎�3yF�ӇH�M��	%hH*��'j[�9LÈ��h����v�J�M��� #-��3+4���]�m�çW6d˻�dn+#f^�m$����L��!�3Y�Z��c&����Yj�d��,��њ�q��m*Ź�.g�"�հF�m��zn�&6�%���ڨj�ǡ/�r֣�t��1'6���Yڃ25[{�|(f��ZT{�M��wD���K�8.ۋ�ܴ�hӳq�Whe茌�YD�bGn^����9Y4�p�tE�y�f�
�tS�	�kk�ŵ��,کd�Zp*�v��Sw�䧛��hS̭V(	��E��ʻ*ed��J��$��_��A!`�t�Yn�ssC4-����e�U�^�֛m͒���P����-Ĩ�SL��䫱wm6�H�nn4���,�� �H�v0nV�-����\ʉ��jE5[���C!#Ѡ,��A �\���N�(^�+4H]�a��5��%V�V4��´<4iyJ�W�i�zH֬��7n��Sֆ6�M��	Y�%j$ʋ�UN�DP����Jٔb���w�)i�;���u	b�8.��(��$�L�������ma]���Yw�o0䣛fDu��J�Rݸ�Z�V��"$i`6����M'4R�GI�aV�������y��X���9 �D0��֔4Y-H�}7cU�-Zi����/ �������da��"=؜cv�E�����R�EOR���3u�pn����HAT$dTZY�/}�
J`�j�M=ݼf6]MVotd�����	{QL$eÛ��!v��,�ܚ軷,ӛ6��Y,謽�Ӹk}IЦ�g�ODt,���Mܘp�E
��Y���o"h3`��,�J�ǰڲ�����(�be�;�y�`t��;GU�LbƆ�9�@q���
�^���Tt�)dL
�>�{���������X���yn���rlE32�j�[�4,Iȇ�9�l�,���5�����z�ņ��"ZArC���a�lqUݬ��C�l*y�Șщa���Ú5djdP��q��;���Hj��SX�
�t�^%[DSHMyy6�*'���i�C�	��B)���5���2��^���5��^��*��I���sEYT=�L�34ߜgh0Dj�|5<�2
۳z�Rɲ�	��x���[vdy�q6]=���B��ꌖ�l�Q�M*�0��n���YV�����&�.����6e�yP�	�l����#�Eu�EM۽dV�˫G"���=�7�A0.P�r���"t�!YP`���x�0��{��͎̩����O0��੓�嵸��(���;70�^���2��9��X�kL~�R�V�"y�)���"�j�����J��ܫ�]���6╒�.8"5�����"��v�d��4X�06ݦ��`�dJ�!���Bkds{��;�Y�?(8���'LT�
SV1��[0�%�V]��j�檔F�:)e�v���zsE��ْ�o�z��
5�b"�``���A��B��v,5mn��1zRz&�h�
,e��)k0����暺:�,�Yl]�����I+����Em���i���FLJ��/he��m�ݶ3������m�u�L�v�96����T�l`k ,�'��c&�ӆ�V5��f�*��1�nژ��َ��e�*P�3w�<K��v��f�p]1��$T��'��	���n����V+&��:fZ�Y�y���c7���se2�]B�Ѹyp)�h���� �3a�b�&ƊbJ�0AI^!H�u�!h`�t���TLI.�%�xXN�d̗e�A�
�樊��rE��\�3�FHa ��V��Qp=��T.�iP(�D7�>-����V���:Gg�F�Ij�"�K�`��xj��%e��(�P (@�j3
�(}*KE�rl�	�8 Atf�c�m�@"��/��|lEBg}$D��8kcl�u+�}hi��dQt^��C,H��5��j-e��g�e��n��
��D"��~��}z�7�3{^t�y��y�2���4�o����m��m��m�.��v�]a5I�4�f�4ؒ�i�V�Y9lkm�kL�9�ȉ��e<ǤfE<��6���r�����{�G��I��;V�ԦF��7Ғ^���w�ޭ^��N�"]Cc��X�X���NK<�IR�Vhf�����Hif%[h��r7g(�5P��;g/ma�����,1w��bp@w4�$���"����ќ�ڽ�޸T��rY~{��6�A�&(�,�qT�I��d��hmfwwv����b]D��{8n�+��t� ��\Fվ��[�n��5M�9�qen�u,(w']�W+�J ��3d�a��]份C:�Q�͒S�Lo,#+��7y|:gN �<�`2����(�{&o��vk.�5e��m>�Cd�G��Y��-j{]�(dT��֓������{Ru"�i�3;��5�;H�"�
�9]_2���Ux6���خ�oz��<k�]��M�.��8���۫i!"�n)ՠ��ւ��8n��]�Vż]�Ww"P���Uu;FS}Ń�Ey�f�f�&��Z�a�o�dM4��RvEC�QT��-z��S:/���݉��!��Ƭ=���g3�j^A����̓ȍ�&�]��Q��t�{�}]$�ۘ{-�A#�V���gjs�Ъ&�0.�:u� �tޮ�:����V-E#�M�no5��oٷltܺ=��n%k5w��	Jfh�3i��7v!٤ށ�C2nV`#�QSr�IA։⏱�Z�������f���.\J��)���b�4rn#�[;l�cV��Zؤz�"�D�FE��{����K��Uj��w]�����C�*1֥M�NήwS"�iΘ��9S�q�.�PTt���4�ǂ�t�+B�q�Z�����b��+�sEwo	�S�qV_nuP/�Dwu[\W}Bر��[~��`�M�G�SY�R���xW4���o��7}ۧ����X˰.���vi�z�٣9,L�C�;eh�Q!Q֬��F�Ĥ����;�&Ze�nĹW���m��v����;���Yr��zgb�����sK�@���B�s/,�=����BVf,���⬓F�s�)�˘,h�1���{��g.��;w��JH��|�\�R٫bC��*x�R�t�*r[��Y!ٕ�r[,�R��MYٳ.`�ݶ��۹���h�K��(�ن'[�W��U2f$��"�����:>.���|�VC�e�+�KG@�ռr�+���uk]�F�bM���'l}�/��K{�V/�p��Z����Y���g^Ӵ�'`�إ��o��k��eѮ�D���wr�[�ӎb���[0�,)�J��A��
�K9.Cq��m�\X(〕F�5�Χ}�-��{&e�9��ylR�(U��qs���-�zb�h'|$�Aa[�TK�#�!����#>�H0U��ٜ�PT4Tw]�)�
���)�������ve!�<��B���#��o0�(cA�5�wc2<�{��K��3���u�E�x�	W���6ݜ��Ʉ��8�ot��Z���Ð��H^�R�w�����Vn�fO/��9ʺoa�,�趺��.;��o'Q�h�A�2�X�J>�r�h�T�6A��!s���UN�*)Ҝ�ƊUu�C���ac�{B��RM�89K��h�ʴW;��g/v��{�	�&�oe�.�t��ֱ䃚�L��$��"�Ys��V��<�nn)TpE���}�.���vNu
�u�օ�����3n͊���K9-�Щ���_/wA�/ga���ӽ�C0�.��Ơ=���]r��h�fV�g��w�k7�q��&��廒�����mq��u(�⚝j�V��6O���h�#B���ɔE�f#�3+n������mw �w_1ݝfY��/Z�}��;ۙ�ʺs5��mpw��U#X��h�M��\�˓��ҳ-�*L�� ��1{��'q������DsK3mmn�!�҂�;{❘0kߚܮ3y�ZkZ+M���(�ϋ�Y6´yf
;y	x��Hݪھ�4�w<�J
��g�nT�l�ɕ{��8ǭ��ƹ���ܬ��f��zG��A������y/0J�&�PN�=������gy�SO U�ܭ5C��Ze���[��A�<U���{+ZgF�YmeI�f�U~]j�è��
f���W�=��{W�y)ڠN!k"�mFh+�-�I��0�`���y@�e��8����@�����;o$Ӡa��YG��S��ػ�&Y�=6�Sj�s��T��W\�e��f���/���!��+�[7�Z.��u�S|!��0�CDP�P��8D���J³ %�p�9�3R���q�׹b�/ַG�4� n�,{r���y�o�v=��Ļ
u� ���<�+�ˑ:����i���I�=3.������{�oHovfl�r]��ƨYL[����uX|z���m(˼�t8��6QT;;ZVÅV2#ݢ�u�� >�N×[�/�u���` c��Q�t����N
�9��Hm��dm��C���Y��V���y���כ��l�wH�#�Ʌڄsf˱՚�91�f{V�
��^t ���>ۼ�9�wV"{��ћ�5p3�n��n�xV�,�t��J�W$R ���w�Ї�cz�������-t�Eh��6-���37����	�T��O�T���]�lިO`�`�n����a�4أ,:�5.�k�v��(f*��7��ۧ1�]j�W��2�b�/v�����U�ޤd
w��cV��=[/���	������Ƴ��/e�ű�^Q.��赳���� \�)]�s��i�j��֞�{]�I�Xi���N.k�WEĚ�ټ�*��)ue�UD�F�C�Y�y���,R�M��&��K0���5-XƷ}��n�FYX����;L�g���љ;d+mʋ��"P5#P�G޻|"�"�i���]�V����wW�WK@K�PmQ+�����1��
!F�e�s����QS� ��������޶�M�w��t��8Ԝ2�^�l���K̃j>[5��F��Gk	I�X+r�9Ս&u��` ��ƹ�'�Yʇ��\��c���q}t##{ ���' űb�`.��v��������75�����a�\4
\��
��
����E�{�0nH��jڝ��'��5����gZ�@��$�˺���],��#ȃC�q�@t�Պ���#�FD��U��fuk��u%�����/ra�e������Q�8<Z�(r�jOq�6Z3��̬�5v�^��1����h]�A�V��*��"Ĭ�˱f����bmg�tM�-�{��8�[J՚R/��j��a-�kL|������� �g��x���P�g:�B�R
��n�t���U���٬����#rQ���&�}\�Z����ߊ(ˆ�`m�v�ĳ��<ܡ���;�����h�Y}����-,]E�N�����WŪD��l%�"�f財쬧;e¢U��j^F[��[�Ǳ57�G'|x)����g��K��+p���e�kY[Ƕ�=���c��Kz�]� +V2���澖���"�t]k�X#m�<7�4\�i��`���VF���G�1}��z�`M�KGSՕ&CP�X�$
.n�wl�[�w-�/OWj�<�y��:�&��R�K.].7�{˛|T�w�-|gi��7���_	ݩ��r��*G욥�V��[�g�%�s��(�vd4�TT�uz�[yP�ʻ}��t�J�J2�hbђ���T�.�EЇby����W,��Iʵ,2�y�+Oݧ���u�A�J���iN'��.K&�Nn�b��:U9���L���Y؈�9��M����M��w����l�T�b�ŋ��^�A] ��wW�;"�╄ɻn�ȳ�k��1���*5�p=ҕ�/_evn
���Ɂ��3�P��T�[pWͳt��Ӳ��K�X�N7�n-N�+�HPZ� 'kw�C�����v��i�;�F����=η�6�d�8u�YZ$�Ի�N�f�_L/=�3x�%�]�X��v��X4���!ˋ;���G�=���T�Ǟjt���vQ�3pa�M�r�兔�p��{�-S���o���n
�^z�[������Y��+��9pZv,�	�xF�6pE�f�m��Q��e�'t�qn]DER���y":p�W}5����q�u9�c�y��y��ˤ"o�OFVL�d��8޸+�r�W��\_N �6�Z�'�m�^ʇ��h-&V]�д��][���.��+P��,�oJvR����r�s�{y�n�괠�Y"(ă��Q��j��gD?���.�:���间^�S��cC*a/`��ew�u�&��zx	�wS�'v�[�����q��n��$�W�E*.�ڹ���Nz��kU5���U�m�Om���ne��-&���ۘi�cs��銏v�NF�yM�4Lmw3�����+��_V�&fy�Tm�� 8\�깛� R-��'gb��$�0}H�*��Rb orv]z��Cm��렺�.Ɗ!v�^�׊�Tl�n��ݽ��6�7���w�;���Bӈ��6��{�5��γ{gso����¬��e������-��J!����,x���Ҏ8<y`�^��yd���ށX��"���z��<�)�QT�P�f.-��zH�0d��'��̬^�}7^i�ۗ�
 �J8@$��9c�ŭ��7�&Lǚz�Z�eu��Ps��0	���2��vg^ǻ�ٱ0��E�Ǥ����Ky��M�;p��xP�ً���7����u��v���,�v��F�32�fd�����ddb���h�0�<^��\7T��6-f�EL�b�:�C�]8��-�]���A��l�'�|�����n�u��*�Kv��N���������Y7]������Emƒc�0�x��{\s��ݭ������Z0�+�����q��7�#�j���$�V�xr)H��hB����ʠ�@�R��SMN�B�\�=�)*���c���H�d:�A����ía�np�z$���<��t��t.���D-3f�;օ���1�7�K��陶.��u�u���#�۔����u�������&��ɘ�����黸%��l�v����#t/�vWue͡xT�GE��	=إ]����>���م���6��m֮����7���~��۷T÷u�KeYB�e`�'�|��o���k���E��!����0fa�a�8K��N�i�g7pqv�^�WKr�i*e��؜LEe�e��4��V�C�'x�U���A��������3W60�ʱq�r��hܻ�J���G@�����|���;�j����V�۷؞�]�I�/.�d�Y���5�Nb&� �2����}�Z��r�U�HgV�DewR���ef�0]��\5�B��Y�Wna�w����]f�c�V�C�GMS^��0�+AV�էF��WI��[�W)6@�nm�	�����Q�rSMn�Q9pM!��1t�*JQ�9J���n[�d�AG*����usUYOO^J��,�����1��u�����[����gPu��l\�X��aʼ1Cq�s��h]��a�9#e˩Y[��&/I�3��:c4�kd�&`0��mV|w�k\�CN��!K���i\-�s��1!3D���VQ��r���5(SA�!�����;b����Gy�V���{Ee��F�eӴ��0�S��uosJ��̫�x�L��؝�2�p����d�3:�룙�S��^w _�r�)̾�7rw�"�]�v�M{�\c.#0���N��v�[lwP�f��yi�/B�p�*5���ufx�͇�B���s�3&)ytyvr��Zi��د,�ʱ[�v�@�K{wb幎Ӯ��Ԯ�ס+���|)��}A.^CD&�,�S)n&��l����)rjt��׸�vg'�2�t�������ʄ������i�e�Uf�*�r����X����;�#F�fD(�.��n��p��5������X5��^�շ6�m�c.	:�^;un�Qƛ���0�\��t��2��ȝw^Ԯ�/k �1e��lǝ�rDE���"Ħ�}:�9Rf��n���9b����	UGt�q����|����b�	*1^��qvýש��!^R7�-���0X���Bw�ah��>��H��pL6E�Q�\�<���\�gU�:��Z
�&oie��.6�a�_U�k�\�2�Nڃ�����m#�V ��ٻ��n1��J˭Wp�Lǖ�� 2L�H�d#ǝ��l$M�e_s�@��z.Ѯ��VmCYմ-�i�M&�>6��:h۬᳴A�p�{B�nJ�l��r�E��{Y2��T��R:g��2�T�NHq�oQ}*�&>� j��<�Fʈ�tYcZ�<�{V�w�كZ1Z�0V��#X��e�����AN#ufo'�򎀹:{�<�JՅ��r<�e!n`��3ۤR��C���N��c&(��s�jb��JU,����պ6�4&�d�.)o	ُz�x�m���Z�я�􀁴�QھD�E��7�f���(���+�u��u�L�Z��Zg�Ő�R[�1�I6��ӹc�d�WM;��;DӂX�b&�jԪ���e�;�y����nsN��m���)���Z��Z�(ocC&mwZ��P�ª�ԦF2�캷7�K4����m��m���D " 1�z�������z�����?p����O���������G�����K�IA��� t�G���>��*z�?'O����# E��~\l����f��4��M�TD_�����&���T�[����s�H�)�7�1�^��ff
�5C��H��sV;�=7�q�,*�@�7V�e�6����)�hڕgft�kCnTvT���eʘ�5^u����ˮuǈ��Nm�����su�;�-�9�U՟�I):���tȌ�@H��*ch�W���Y���'WX+�H���YA擯f�G����=�������Uۻ9���)^��f���j��
�ܧF1�j.0k��7q
�ֆv0�P�q:^�&^@���@��nXi�;3(�)��/"�ͮ����YOf[f�H.�\�	rq�Y�L�J�;N*��m-5�a�V�b��b��\7�b� �6+:ͼd��[�Lj���W_X3��@Y������o�ޝ|���N�T���6�\�n���^����t�痷���MZh�yW�U�<�\ԧ
�[�N�%�=��j���JTn�km-<�z�I�Ù�F�Y�P@2���,�����( VT��XN���E��4�k�d�{��j��Vs�u{e��
�L���=*�-�����5X�*�H�	�Rh�s/���j��A�b'�Xz�WM0[�F�k,<>�Qa8���G�;��d�T����h�a���{Rg�+��G���Yv�]E3�SW�x.�����׼o�M`�@j�3���tV��R��T�=�r�ܟ�Q��dG�k��u�ܵ]E��zî;o`X�b�î�5�u;Ԛ�۪�I��*�����{(D�GI���[f����)���Ϯ��gF�5���GQtk��e����u?-����!���D�&N�,w��d62���a�]\�܂�cU���&�ojo{b|4�s5��e^�I�.�=�j�9��=�76�m][UR��7�������/P���G	@x����b歛��ɋ�[u����U8e�HY�}�E#�f̦���n���!>�/��u�Sɹ��5�k�Ź�o3#[d<K9嵶��tz/���
�il�1.��x�������b�2�^QGw\��N�bJ��O�膭��ټ��&M��m�3����{J[uAs�Y���rvp]��]�0�Z�G4�a<gÅ��	i7�]qލ�ÑST���x
Wǥ��h�=F��;��{	=A��ƎQ����x���wH{�3�{]1`�x���y*1d˗�J{M记$ڻ�J�̺#Z�m(L��{��l{��J�@m!بK��U�=K+˯_E�I�iu��=��kz�
ܼl���;|�j���������g Mܹ��^%�Ր���35�eDp�E��n���Gd'�\
���nM,��ܦIl�9�gaH����hU ��v_���v��]��8p�f�5J`'E+ki��c��JJV���hou�o(f�ݲ��_���7�I���)i��81�t�(3��Rl+�
o����e�-�.��ʸ�ol�Ԋ[���y����q^�ӫ��*��x�*@Hye��5G���Z�p����ҭ/en-�T9L޽���xi�F��HH{����ԡj�u�L�yu�e&o���\�V�a���*2�g�gZ�7ڕ
�4�jQŤ�� �{������!�WAR�S:��_\ ���WWVߡ��wyn�5�w��C�%֬�J���Pݧjr&V=08#F:wx�-AIP^�[�LE��+y�W�Vl������Y��5{�-�p�s��tqB�ڙz&{�v�O����Ԁ��=x�����H�)h�\5���Fw�����j�F�	�;�ܫI �[ګ�|�J��]��8�W\���E�"۬Q-$ل�Lǹ�dk���Kݰh��c�����u��U�U����k�.\:���R���Tꚡ�N���˺t�[:��J���,A�+r{q}K/*Չ���o�*�<tWq��~f�(IY���ZFv�u��IwK)s��@۵ �lfu3E��F�����;�CMR�Xo��%�{�%e*)E����j|f��HM�(ޥL�*%8E��JѬ�)4VΫ���A=|��F���\z����rb�Z'�+'s�����i$�7�Kt��ȵR�Q���8�[��T`��ۧ��]\W�E��ܜbRs��di��چp���Y�d@��jÔ�U+Wy(����Н�W]�z5wݝyk���@�7�x�P[�&���]w7r�b��gT��SU����������� p�D�M7X��e�}���Th�F������h�������ݦ�<%�Ω�.�AB��P̢�E��lO������3u��}�׻��r��M�����˕�������"�ǙJ,�N�ʚ��ń4�]�`���H7���fL�a��g��`P����sCŨN��!��^S8���<i��.f\KHb��$�o�&�&�/��\+Y���j&�<p�4�
�B�����T�AK��cv�B��TI�������Oc܄����������+�c��5s��s�2��9Q%�f��n��7f
��,Xݭ�㇮��;zVكe�#��@����^=˾�{�q�<c�c�Ҕ�.f4����#�k`{&�!+�6�A�E-�he��V���cE^P3.�1#��]ܕC�}͛3l���4A�q\��o o��������ހ]�VVɶ �;2��f&�غ��9"V��X�̻=te$V0�+�d�u����͵����+�޾��!M���[W�Vd r㙉H�h\8�؜5"�JE"�n=:��D��&�����t�̋wjV�;���e�qr�%*b�1Dʤ�:S���[L�5��w:�q�E㭒p8�]��mVn��t�C�H��ln�FjЃ���hZcEB��{R�y+�F��]8Ӿn��_��KyW%wyY������t1�Ԭ���t��Ѭ��c�c�;���2�X��F�*�ӱ���xȈ�ݛPJOj霨���u-�s\���YmB�r���e��]o;��5�e�@�h�גz�u��Gj^�z�c��:vs�w�P�vE5t%�����&�9)�a�y��}һ]�/�V�2���*�&��9-�![�\;&ج��v՞$3EY�9B��j˓es�뵒�g �t���Z}SG>��u10Ǵ���Kvm��28���K5�Vfe�x툍���٧v ^���͡(a�ۼ,*��[Vj��� �P�3�������Z�ם2�\t�k��v��L�2�i�ʺ�wi�ټ
��Ž��i�t~��ԇ9u�C4��w��`�ZN�&�$-��)׈�7���S*�T
H
u6
А��Q Y�|N�Y���0Q��[�ΠB�ck��U��w�F�av�v������Y���X�vF��f�$�B&�_���f�Nl����^v���Bndq�ц�r�źO&���sa��6Im=�Ra�V� 0�U�+I�WJЂ,�d)z�4;q��R:�a�;:������޶yShӬ�A)cS���b4*�p-8�k7qzMc��j��ƾ۩t�E7�B��;Duʨs��Ye�籌曇��F��.p����y�[��L˖-�5R���M�4�i΍�M���]���pL���n���u=Ld}Æ5ڵ=��K�jq�46�A��;jws�|�����Lh_�囶Z�&6�M�[�(^����kSF\��Q\(�{�i����U�nxm��^S7xnk�����X�w��]&rʺ��u��Fڢ����V������du�!��l��){�g��i�˾���]tt��6,�J�6�K��������\�tyq�m�vc�c������nʉB����z2�(RxVЫ�a�+r��u�oZok&��twn!�g�67��'��q��Ƀ�ϸ�,��U�,Î��&](�!�aS�6`�%�y�����x,N.�R��/�̓٠��Y]ίj	N�^Wn6B��Wo.���w<B�*wܷ(�)�,2�v��d�\^e�Q�h��]۷u`�]y��C�|�L�xn:ce�Q�<�����(�ݸ�9���ޝn�`�4�KŢ�z�kZ��M�=��F�nԓ�j�۲d��55f3ʜǔWr��@ �yg]�Nm���d�ʵu�����di���%�@f������Z�5ό3�*V٥M�����V���ݣ8ֻ:�.�,u5�6fge�9���5gc5��7ۗvMJ��`WT�y�V@��++f�}��;r�U�@A^`� ���&�s̸�:�n�7�������tv�s9s�#�f��Q�mn��q�&�6�����l�ejZ4m��z	d�}�M�Ǖp[��V�W��=��[LVTsa�vx�}H��ڕ���;Y����JH]e�o���+���h+0���(p�n�f���7i�c�N���]!�+3e��d�:^聅܈��Mf���uNUٶt�F�e� Ǩ�]�7$ᚧN���F16���Y���On�j�7]ޙv��+1��.qv���C�qR�LC�V����%|�T�;n���e��z�a��v���hUʱ��]�,:]�,�Wij��bKB���uub(D�H����wx�]h[�S�,�PQU�81tkU�;og��դ���g��W&�@o���V�aK���J_��hZ�zƍ��c�E��T�q����e$�d���MW9+��c�E'm�3܎v���+��-�m+�4+�a�a1u�ẝܞ/5�(�M��^ݍTXv�B�WI֘�[:�U��e����1f�������cK��pɌ�^nݽ\m���~2��L�׆v�#������,� ����#Yڭ��y��^+���ݚ�e��=̶&f�i��H��d7��n�M��-��l.�2��2�s�9��InCV�")�'n6�ƊEd*��(8.��\H�ƥ�q��P���_�i�[�g�f�L���.�(��4`��ЭYG ��"�`�����>e�U_�4���ܷ)�'xн�R��(S��ݍ���VEBL�K[����	��Kߞ��*eܺΗ��6�u��JK�܊��H�<r[�����3��7ܒ��n	GKr��Zxe��BWs���l��}j��h�0˃��ɉ�gu1iνy6�5�� �+��k{9�&b���V^��s2WK������NK�R�d�{wr�*�ԵX�z�',S��U�e��2��OX[��أP��7�U,sj]�V����U9�.�k����R��N��5l��:P�:�x�)����(3�%�4U�xQT�#�7s�kp�U��AiE�H&�1]��º\P�q��E!ݷd��9�A �Yel��L�d'���W���j�r�g]��X�ogwbV��3#@�=ӡ7��=�f�n�n�9�0J�W[t��ں��w���L���!ݰ����j�l�D�@@�d��V��i�|N�o�w B�����2=��<
�06+�j2�#5���pg-V�{$�r��R�8wvhhxxb�ڨ��w!L㆗J
Ů��}��)���V�*:3z�m� >��,U�ʢ�R��r�*P�	�y�eٹ�'gD��Ln�kO�rih���O�x h�4Ӽ��+����b�qWzt�u����fe��8r��s/7��X|fK7W�X�Y-�}��j &F��b��� �'+$M(۷a2�#u�T���v�#g;�Z+�<{�6�<�܄h�K���l���n�5Xic]\�(���*����!��&B��f�=��/;�̤҉\�f�<�4P �sc#��^�{��!��r���[�K�)n�WX�/�䔠�L�yxQ*�vp^�,��v�K��ȕ���B�NP�ϰ�-.���{���3yw�J�E̢��V��)!��-�t�z9�y<� ����k��Ly'ZY�0ݎ��S�jc�s���,����|k6�f��)^��;�j�F���Y��VNA)dݽ��{�,����+y ���ձ_1�(�,UI�P�0�J{L��\]�j�A���*��B�n��go-˿�Y�N��� �G�O,u&��u�:�N{��U���]���|C�z�.�e=K6�k=[d{��fYt�*�u+�m�6�]�3]����e��L�1�+W����X��Ut�����LB�P-gٔ��!�r�$`�r.���Ad qfVG4w�N7��}�L!��9���1%4/T�Rn5�IdMZ��x.��y�ʼ�N7ˀO��>�6<J���3+�K���)H���y��(�`�Z�b�YP՘�*�:}rlg+p��{cnII_r�]:ˌ�9�Z�N"���ܬ��'LIl�-��P�q�)D�)f�PWm��7'm:�WI�hVzY��8�7�ʹ�V� �r��]��.u8����=������M��vK�~��:"�LVպ�Q����.|�PejV��|��Dd���Qbc΀��ks�NZ�{�ݷ)i5��lI��U٤j�{����j�+c��f���Zd.��saǌU��J��zvI6>�k��/F�-%��x=��S'D똍�Y�|���9L��DfᔊT�����F�۬ѕ���on�7���o�6ڲ;�>�{��+<Z�㠎W��X���Bb���	�Q8��Q�a�U�t�ݫD����=��-�����`��0N��kC̃A�*C�����tNOR'k�vڦ*�"��y�tn�W������Κ��^�E�C(����3,�+�2e���+8���������;(�}v��d��u����x�K�:)�t*8h�a�0c��WR�qA�%�Q�Vb�Z�PoX�(�[S)��r�x�u����]V�>>�^n�M<׀"��NӐ�ݬ���J��+Ue�vUC�I=f9Y�VP��w��f������D^Q�)�ٿ[�^qd���;{q�G����Ӵ٘:���bTǯ��w2f�%���ǋ�����P� �� =^�~�w�z)�<�W����z��#,��,�nݻv���6�P�"A "S�AF����!���mY�6��f��y�G�Qt���ۣI�E� 25A���@0i;)dT�-��z���D�Y%�L�h*M�`���|�+��z��y�3r5a�0���$�n'��QV�Z�.rح�aC�6mi�ʻ4��H�2�Z��"1['f[F����]M�2�ђ�ܰ�ݳô#������3o��c�����'Mh�U�WneG���ev�C��-]�U5]8`�!p���X
���b(f�J%�J�Е�q�ٛgtPq���{�]+���]��*ؓo�-������fm�چ��4&��\�:K�E�ы�A���S0´�N7�c.���7�GxkS���[[�4�vB
� ���Q�P7��M�t��2��'� �z�d}xm9v��h0�b���n�;t��P#7orX�wf~ln_h����{7�8��v\'�l����{���砛��E��5�lO����T�n�g8-���K��E���+]����a���Ε`����Mʵ�ġiݨ��\���$�9�vI�zc8h��VN���Λ[jp�V�.���s��`��
�0�`ъk5�;�2�.��"���Up`�;4��ur�|��<U��o�)$�骕�O#�q���yc	5Kr�V/5�q���2+Ki�Iɺ�6C��1%���E�Λ�!�ؠ�]n�!�4qu˭ޯ:������:K�ۼ[��Wl��;����b�/�-�>X���ǫ���_����N��H�@�� ��!*%��I�h��@h���&#�:A�^m�Z-L�!P��m[)*�d�TQ�$��:MN��H5E�E�
i
 0�*�4U�����㫮#��v��ǵq�d�,4(Z��4�4�R�i�!BN� ��,�  �@�SHi�T�`)4�B�0Uo�������Ѭ�LI��UT����6�뎚/Y��b���QDm�X����a�T��STD��Q�i�l�W��=V&���<LAMA{i(���S�60Z5/�UHU�4SE%���f��6������i�Y$(8�*���i���E�%�t��6�Q��QMQ�;f�+�=4:*��l�Nƴ��*4hӊ������j;c@Pj�,F٢��+�K���F���5�E�D�$���1l��j���Ӥ�5MomPO[A�;j'I�(=�@A�F�w�5M5��-uF���th�Κ�Bn��닣^��ɪ���km��mb{e�ӈ։5�6ͲW��{!� O(�H&]E�S���"����1//%0(�Z�j,E=R�
Tj���'�A����2�pDS�om:��mj�J�B:-��L4uT$�E�N�!I��"�i4�~�P��L�0��T��������]t Bh�p���+}�noS�t�91��r�p~��Q}:���tr����yI��Lvp�^s��\�3�ڹ����9цt�}��6���}�WWKX�;�Y
�w09���b��q�Z�<���՛��g�cG�3����-�5kJ{�}�����cj��.赊[�sU�l��\4�ܥ��'��\�勽�jT�kz��)9-*m�Я���a�w�6 mp�pr�\��a�븻����7�&�+�����U��sw�.��>F
@���r�!)�3W:��;�	��|�u�_̳��:�亳�.�C���)�h8(6w�V�X��p�����ݗ�R����\���}��f��o5]ѳ��r���aCY���W.}����s�U�����3C��;"%Y�z3L1,���u���V�V0�|��	�^Eh�B��7�'�6�޴��EƸ��w�L*�&�d|y��9n��b���ozv^j�5���*��c��n�
Z�����R��MsJ�ԫhN�LEH��"�!��M�E�\1hV�b>AĂ9��׀��`�h-桇�)�|;����3��m����T��ptD�d?�d�c�oOu�n)ɸ۔�A>P�r!����,6M��g�_U�ͨ���������s{0>;���Z3�����:đ�������1cV��ʣQ�'Ff�}g/�6]`�$_5�e����oEO��6��2$�AN�y�FO��E�W:�K����P�g)��(�$�}��g;�:��s.0��,�d��;�ʹ;�F�8���ʖ�ň�DB��1�h�œ{[�^��4�O8����0Jݵ�ב�P{]Lm�r�b�Y���r�m<�C;�zu�����o���&��2	���z.g���
�<��m9�sa�W ���\1à��������U�}ū��n��B��z���ܩx.��X�f�t426�LZ��EԆ���!"լ�V웙5�8�yQW���:�8ػ��	k��T�'[!��|�[
�}9��P�^�Q7��
��,�i��oON�۝c��4���x3Ņ��Z9]��V�v�ژ���gz_v1�vo���Nu��Ȼz��⛠�i�A���`e���n����h���_u.uՂ1��w�RUz�{��R�@f�\@jn�%2޻Ս�V��c�O]䫦2��0��F�鷷����Ȯ ]@��%�� %����.�� ;���J.[r�{�8��s�=��[�R�X@�� ���`z�Qw�Y�y��cP��aKrҭ9
	�	�ⵁ�+��K�!D�΄�k�[�X��1�"��'=�Гh���s���ӆm�V�<*bA
.d)ݎV��p�ڛ�A�pcs�����<�$|ι��l4�hdcSr�u�3^��H��8���L�ۛ�ʰ�A)�Ĥ�O�����=wJvn����Ӵ���!̈»+d�?d�
��G�#3��Z�Mm�}�g�fn.�%��Z%��޻��5�zw�o�ˮ$���n�Ucy[X��Gf�jJʝB����n"4e拭Q'L��@��R�K{�_aF���ט��*o���8}�P�eU䏣��ؙ[�f4�n飋����t�&�2�:�C4t�Y�%�E=��v���v��)p��v\m�K���^�v��ѥ�B'0�	����&������[��y��}J]m-����B�o�7͇4�����.��w݀o=�L�=w=4�V��Y�hȻ�v[v��ηD:؋���H�$�>��I�Y�ry\	7S��v�D�'��ao�a��Xtr��h%}ݢ>�W��wHn`�4d���YW�����d��6��+¥�ֵ�|��^7���M�0���3/6���wwR����g�5j�(U���_K	X��a[����+�8-T���q]<蕉ȯ��V���ݮ1@t��v6�5�O'j�v�Q��6�h��+����)���m�O��%��K����?CT��C�%d��ۜ��YҘ3]��+^wOjA�|�w7o�PkV!j��1��K3�&Ӭ��c~̀��c��Z�{�B�)�����紾)�n��W�*�v�ɶ�` !�/�fr����߇4�$��p+�̝A9�y�w����)�U3����zz+~�= � YXz�����������r�Ż\mL�JZ;���e�=ݽ�v�/��c+�wND-׹�=c�S�vo���/n%m�z�IO8�b6/!�sQ()$�ͱ��v��ֻ��7�T1!��t�_gkK2��|bk3�{IkYda��B�Q<W�k���7��HN�10�S5�V�Z�K\�%�]����̊M�23�VK� hu\1���e�nu��`�o��w�&&�1��ƈ���YF@ا3��c�P$�n����«S|�i]���@Q����[Yg��ï�Ο��>f,����f�.vsd3���۫�R��|��B����Q�p��o���}���`h����3��73�6��zd�r(u1�~�����\;�G_�{Gs�\�X?L�Yy�B�:���Kݰ��^lM��pۦ9l1�k��wt���5q]EL.�ݳ�E<��7y���H���U9�f<�NȎm:�}���FUvC7}|����s�|>��Xn�� \�Æԡʾ����Ygq��,�����E��g3�}�^2NH�t��D��y7��8q_��C�fj�����9�&SΥ&P��r��X/(:J�aU;�v��+m�4���oB|�E�0jRU�I�(�n�EԔ�,¾+��,��`����u�욥��b��(K�142��CF-��#��C�T�{��w7˥.��0h@ߐɑ��sz\�}|��L1��N�����c!�q�u<亰¬v�wuƍ���,�;��s.kRw�!Y����n�`�����]�ݱ؄yq�L"֩��/]�B������c"~��	�m�ugg��sΕe	�]%R�]7Ӭ�sĴ�sL��|�C����s����7_G,�A�P�%ҫf4��f��xRM��9�,&���dc��C��\�vF��$��7���\�*t��8��Y�S�#è�M6,�	�߃#/�5��*'���\�*�
� ����.�֫��0��ǡ#_��������s�?aΰ�%ڂ������<�[>��(uW�CQw!�2ⳉ����=l����.�tYz�^��[�꾺f�����2X�+��(���o�G��Q;j�3rͭR�KS��*q��T��Y�浸���]$��K4����ˠ���k���R���oK�8�Z�mQ�e��y���Op����s�[���[�:�ҝ2�}�L9u(x#�f��e��7rk�=J�aj�a�j�w\7B�K&�	���-�Si�2�w�n��y=y�<;hh��lQ���'yq{���{�b2l}yڧP�O�� ��u�+�>��[�C���ؽ��6�we�X��9�r������������I������X%jsڢCS3�}�R)��&5���{	�{"�WOo��V�J�v�wς��z���w2p�w�&��ޱjO7�e h��zi�*��r�n�t��yk!�fr�^��j��^F���@��¯�xٵk<��uٮ��N�A$�H��x�-��l*����xK��!���v��^df��ڹ�d+:Ho{�OujI��vnߏ�)��a:7A�3U��S��f�6�q���v:O	�Xt*�}(�9Ծ���ٛ6U=�*�4x��|z���ݧ�)��X����"�+�8�"q`�j]��	j��3��oJ�NXD#��+�je^�p�kw�qmh\��?s��J%�oM �i���
t\����3J�\*
d;�+2��f�ƭǡC��x����r���m�W�UX(e�×u ����k˳�˖��q��N�q�g?�U���x�Tι���/�ä�Pdc�Cj�3��r���s��x��J���:�"�gW�O��8�Cw�	6-�w�@�k6 �L��5Ȗ�8Zο�d��~�k�C׃U�3>�ܗ�I�Cgf��O8[��63�o��Ɯ����sGu	ݹ�o `����{�f7����뿑�lg�tï�5ϞAf��K���e৺ko�+wH�J�K헰���{;-���l�sƫǳ$tӚ�髻kD��ξo
�z�	ে_¹��������M7A$��=�C��.Ÿ!�v��ms�.rs�Ƞ����T���@ꔫ��>|u��xwD&5����=x�|nz^��ɣ������V)����ߕ�����5�1ݽQ�*�Oǩ��o�Ij�b*�OÇa-��j����ᛑ*��>.���{��vU$p�'�(�z���b���Z��l�K�k%*�5�c�$�(�w�s{V��1��W8��p�׆��;y��f��F0M�tIx�]<�nw��m�,��)N�Mjn��T;�f�sv��ou��;g�gWf� dT�ț�M]��-��*�ouT���板�R38k}V����]聀�?i��y8�Ƣ�&:!5q:J(v�ER�oq�*��|�g#���ՠ�Ƞ#s��2���jaJ�l��S�4fr�uk�`b����������W,�o0�M`6�B��M5�u�Muv�=��*�?p�Τsf�%��烥Y��6�Ю��x�V�Mr�ut�큅v`�J�G���#1f����$:�n�Yl�#��y�������1�1��duQ?puC�5����y���d����1،�V�x��P�	���|�� �εY.�4:��	��}(;;�	7�{���j���&�0��p��PÝaVOZ�����5v�}zs2J��f6-��������υm)k��M[�ҹOom=\�(�C9�%\FI��'ur�a�v�dJ�CF��I�GИ���u����
��$_],���h�U\C�/(^���w���:�Wbzfv�l:u����Q݃�M��vWX� ~Lq囊�.�
�e�]�b�`�D�k��V�z�Z����S��T=ZVʋ//-'�A�5!Ι�w#6�"��R/�I�8�(��Q��89����էw;/&���gSu�(-b�[��_�9�����RJU;U���*�o3���'t��sb�Yp;��\2�(�+宻�/�d=�t����Y����,b�A$���5S��8\'g�L%�ζd̓3W��Oj|jqžu�I�zO�L���>���&L�&�c�+�O.�ț�\�=w�3Ә�:�����.�c�0w��TQ��,���ɂ+��6�	���w��w�,�|���\;�է���UX���ڊ��Q�7�.�t��j~�ҝ�}Զ�]�-���^_8���قb	�<��E�ְ;#�/�QL'BA��r!]�|��R*GN�X�i�S��a��?h�0��9К:�U�C���tg�G���M�gM0�z[���g7"jf�Gbpi9��n廣�]�ά��������6l�ՖCJ�'!KZu�:6ղo~�4nd���V�Vܸ՛�Yz1���C�U�N�S(��N��Y�2�����A�{�6��q�-��fZ�3�#��n�d���V�<T3)%�Y���J쐩����,����rD���0<=Ϟ��0�Y��R�"v*#n�a�0	{4K�J���.cќ�{���r�D�����7V��:�<l+7�D>Q�:��t,�d_ٵ�|�ׄ�b�u
t]�r-A�*L��8��u��8���sw�,��M�1� uC05�_g_ ��׃Wl�é$Ck	>�GoF�J�0[4�Ѣ�-z�f
�U3Nu5�C!s��k�i�m��n=E�3�R�G0Y�]D��\3-Wm˗��`"�u�`��-7��Z'M�o$�g��j�wmlI�7�ʻ�]-��0�wh��m�ј� B���kwC���EL�0���&u)P�,�:��b=��Z@��'9SK:�mf�G�=��P������Z��[f�yrw`UҲ+5�&n�e�lg-��آ�JT,K�S{Lx���Ύ���}��۵�7��u�h�;seu�uC��Y�X�T2�츇�rs>�����Rqhv�Ge�� �Y��a���P�H8�E����fu�̺�{g�wZ��b�ZdË�!3i*��]���.� ���w/LF� �u����:+����H�2�ʑ��7cXfC5mM� �)��t��uf��M�5
�v�X��M�'����PU�!���|i��]�G�Sq[T�=�s@��R�Y�`�S�={��Zw�Ѽ��n��ڇ���,f�}�cX9#wG��֤ŋ0f��XԽ����.�o
�H�Ձ��Ilۛ�#Tm�R���n�0i�eY�3��3����[�6M���̼��S�+1�HV�2E��S9�6�Ԟ�7x�oi&�jP�|ݽ��ս��mRM�*\k#"�c��Y��>��Ē�\3MD��ii̹H�E���v Xa��މL���cz1A�+�ɹ�e]b���}�b:�-�Ԇ���2̘nRz�����آ�1��%j{o��u��}wdo_l�A����vk�%U'�l�d�π:;v��_:��;��N��xK��2�{�k�\�)oE�G�`�'<;P/L1�-�=���tY��etD�KV����'C��L� �BhmN�s�)�{wz{���*�3#�����,F�^gm�e,:���l
��قC|кY[�<����c[V:>6L��f5Vn'l'i�mf��Bm#,/��u�ş,O!�,�£��H�ы*�"�WD��H;}��xɤ���}����m�ò��Z��;l����d��5tX0uM��v3���M�] �o"��V����)�Ճ�vuD�V�Op�>ܾ�Ħ*x��g�>N��	R��hP��ܷ�f�FN_�����/�쿶�T��5EA�4'I�֪��cEFʹE,[j	���Dt���j�TZ8�j��h:Jm���C��T�#F��(�P�mc��Qm����&���-��,��b.�V��T�l�X��Jq�*�e�111"PTE4h}ا��-<F������&ڇQ&�4������؞�L��ѧ�4�TE��h�T툨�Dckf�lU7[�TLZ1N�Pi�[��]�E���ݺN�����"�=ih-Dkm���qgCA��(���m�Ő�����%n�m~��cv��틤�G��"�����Z�h9�q�v��]�ͷ]8�;��U���q�x�7�{Y$ף�]h��ǣ�"��7��w����=��pqX��Kz��o]o<L�� "���Uˎn��������tfi/$5E;	$���![V	ԄeJ��=7Q�X�y�^�y�
�1��4�����]���]��=�,�N�A���l�HrC�7��b�)�ߔ�Q�/\L}G��r�@�z��������c�^����Ӂ�i���Qa#��/��5���B��K�����p)!�ZxCCPi�f�VFϕs�kC:��֖�������sb�}<��ɛj��S6��/�U���LA��)<�&�"�;r�v� ��e�5t�w�`qm���Wz��8N�z{��ޅLy�Yp��׽Y�/>��`-��h��Fq��|��[yྲྀ;��@��D����~݀C|f�x-yU>M�4�n�� ��c�0bY'��>�e�L�5؈�|j�t��{w�R�.�-�8!���3HY�1m��NÐ����!�J��S��צ��]"�W�*Mmq�<�"��8�b:�=��`�����cgx|F�͍��>�n�0��]���0�Gu�;�� �"�-�Ú��.r�Kb]�]]v��}���DC��� ��;��E�S �&�z&-?,��\۴75��q���x����r�Vf�H�������y��i�9���k��M7X�U�e�x>?��F���w~v�}
���#ʥL"��
���
Z���n�e�}�$�3�l��Ѽ���٫�M�EKKb��¹B��c�"k����{�G4tNXv���j���.E�ݼ�qYƒ��hv�>
_8��3�kƉlf�J�&�ۅK!�����>mo3���M��j��p��ô���ga�:@`��"���<�dȦ#���rv���u�~ź�=���].7�8�"���������X���4S���H~B�jn
���oշ���s��eI����/J<�@|��{�Y?9�:Q��0�P"P�/V
q��f�#5��&?p����C�&���>��������i��
�-"6�&+���8?�]�	K���/]iV=�<�{b|� �b��(���WABG��s��4 ���&Y�H���R5/x��)�,JZ�6�� ~��6�;}B����;#ba|��T�m���绣L�A+��}s��R��^���ҿ��b>�.�o�e�m�����F0k{d^f�z{wb���$�l�������a�q�Q�d���)�Fq��͜e^�Ξx�xxd���a�����䇍�F���,�����/�E[R1������Ӎ��)N3�P[��Օ��3:
����;���E��ɸʃ�>���?��&'�i�[�|uϡ�>��p%:��$�T�SR����u>&���k`��)	�?A9���M���������(�%:�L�-ܶ�̀P
���۷��f����/E0Lb��CƁ��V`q�铍d�JÓ.��Q�)
q��
���>9���tc�;��k�'2t�J���.�����O	�T�m/#�ޛb5��T�q7tb�c�4/#��Х��`�f��p��%���$�����4-\�Iŷ��TRɛ�s��+;*w�ic]Ы��!G���t���9�m˷����T�c	�d4J�wNA�H�F����O	�pc�e<?�`܍�AƟC�O�&��Yv��7��~�ʝ��+��0s7y�O�;yb�'X�4�/#h�\���ώ�����П��鰪hMq]1�WtmMr�0���,(�.ycu�/%%�r�vû4�|yp��!����.��$�X��n|�t'�b�v��WH"�$�%S06�y���V�����Y�l���
����)��>��Z�"��������	
%���smv������J簔��G0��:�=S4�:�7�Gw;z�P�x�#��PZD�涥�m�,9��R�StNJ��LZ��|��g�!�N\����M��fGǀ9@��:"}}b�i���*���Px����T�$� f�;�[��P�̨.	���0��g���G]�&Y�^�3.�tE���-���˼@Ȫ���L<��6nq��G�׸3B/4Y�Pr�9�in�&����눺��P�<����W:<��U�_��m�Y����N���&�cg3k�U���������i�;<�wh勲]�IWM'��U�s���v!�{[8���mq��5}����F�iK/�T�X�)SjX��Z���`���Řn��x@�CׁPnF�l��n%�{c���dxV���Rp�v)�ލ��is�j��UE����i��<5� �U�G������t���:(��.�����SGg}��i�${�{�w�]n���1�F᩵0��Z���:����������O�����Y�r�b��})��C��.��S�����nj��M�	���}����:Qns����j^$�d��Hj�;�C��S�; ����I�1�����#�O5y�	L[�x��ц�,�^�<^�g�&�BJ�ߣg1����	�[�Hqm8	ʘ'�ƀC{{5�K��Kfָ6��	�]����'XbY'C�YpIRaA�/�{����EQ��@N�úk2qAv��T��zH3�u��-"MvR���E�fpn�d��7p0i�W��k�p�Z*��Xi抗�EeF-3C.�0In��lg�P�`�&�0��z_�E�气�[˥C���8S �Je�3�ZMd��K�+Qز�_�NK����v	Te�?s�*�w;y�|G	�t����U��t�����_YpY�g�Q�-�8�x.ӫ3��;J!��.{/uKkK�+S�����N�p���������H����q����>0巗�F).š5p�n2���i,�@ǲs[&$!�o���|u�J��x���7��֐��kq�P}�䯺���y����ɟ���L?0�a������4ڣ��2P��"zW8I(%S{eo��O���c�n��E����@�:_xS麘S�u���{���Hķ�ڝ�����^>�)�z&g��w%�׌Xgcc�D1�&Яt�ړ��3V�Z�ڧt΍M���vJ.Yx���7��x�zb���!��D��A�xl1��f�e�^�LH��nG���΅���I�$���;���oN��(l�j�*\}���-c|=r���gJ,5��h���0֘{nOC� �{9���7p�4W���4
�r�����p�n��~^o^3���'>ٽ��3q5��\_�R`&22�ߪ���[�6�5%L�c�:o�&2)���GK�w_*am��!�f�みD��u*���«����*��Q%V�F�b��E^�e����l;�,��ݜ�5��5������馜 �����%�Ȉ�nm���չ|��I���9�����≉d��Fi��J�[z���|njgO����A����yX�S�N�U�w� w��L2�bT��N�yQ'��*w4�ŗ;f��{���7.�us� 4L�M+����1���oj���u�؄XKh�&\3"R.DDV����c�N������xH��U�jZJ�S�Vbڈ��53��lX�|bn��m��!٭L&
N4���i۞��9�K��H�PIRkg�m�p�,_���˲̘�5�v����W��\3[L,��=p�{�L8���aĜ�+���)P��,'���y2�ǒ[�uZn����OQ��a�G�M�1��}�<�^�uL0rt������#$o�굜zv/{��t,��U�f�_��K��_�=J.���11�:��CiN��SZLLc"�^?(��Y�zAcs�-��ą�W3�<p%��S��`� z>��f0sQ�vN��x���&����NZ�k�G�+�@UR͔:-ݛg�a�?��  �\]8vv(��SQ��m���M�-�eu��i�j�Ja�Ʋ�����5�E��|:�!ۧ��Wty]��B"��N�&c/��E�-	��D 尽mC'��!���Nf�P���1Q�z/��0��ۻrVn.��Ձ� �<`�`�N������{��y�]��ɘn��p�mLi�«���Z׶dxB���]5�F���AzU�ɯߏ뮌�����D�dE�����4�l��{�ڛ���F�5�hѝ�b�P��t^��x�\��ؘp�aR�w22�g'��Q+��d;�<��A�Օw��<��[����m�U;��^'��n�)�`&��x8
�v�]*U3A����xȺXQv��	��������x�~SE�d fbb��6�D���?xζ�(õ65'�y��^��x�d!���|�����"��r�l�;�}�x�(8�,����A���z͜eY���8��`d���͞�5�2�x�*�-.��3�,�H�s�VժO���'�qQF�����Ƭ��p��oPo���Pd�n�M)Bx[FG)�3�XƯ#cy��e�`����(ʤuŰ&F�l�nU+3�M6p�Y/(ts<�-��,�Ba'�;�w!ۄ��M���~s�ZF�����QG�ֈk՗���������g"���o@�Da��(.�S�.�pi�醟wR�ɽ���/���3���,덎@���^�hg�w�xa;�#�!��>�!������Y7�kV�;��l���vV�r�C���E�ȺƲ�x�Ms�'�����=��?P�5W�w�fH;��w����g�? :��+;\«�%s�Q˔�QIAbF��o	�xwf����66����L(c"o���!-�=QIћ�GA�:��E�Z��Q�V��݇֡�n�f�7������7���I�f�bF�PE��j)v�I"˚��͑�F�pM��v��ĳ´��$T��F����J;n[�^E�8�QP�����S�5���J9����{dõ[�9Wu*�q�\H�Z���R���:���8�e��{'�G#�x�������t8�_����^�4-'��;�~��a(%픿1�{��*��'67y�t�`@S+{�#���h�A�y�@z@9��f[C��j�Ԫ���pX���{I��{���%�,�����s�ޟ}Ӣ'�"]��t#m��T�$���r�{�ĳaW��if��o�9�v\e���&e�	 �cC��-���.�^�^D<����ؒ
흻�
������Ҙ��CU3�d<P�C�Pi�e�A�ʼ:&�׆�f`0%��ha*f�������B7e'�U�m`n�0�Pxj�#��@!r5�q�>�w[S���E���<qJ�7\H��(��a'w I|Q�]~��kj�����dm]
EI��{�XK�g9wk�>��+��a��b���g�| לl�G;j�N21�M���Se�d&M��d�_vr�����@�+��߁����cռ4Ӂl� Ŵ�8� ����vW�n��l[�܅h�9��{ww�"܃��Ғ�5BJ�.�Zs����z�4c[$2`���>��1�mp�&s�k��^�i�k̶сe�RصO"��8�/��i-� =[aS�W�u�I?V�U�)�o�N��%5G�����`ErYͳ�^�pK�;��,��7�ѡYV�T�!�]UM��Hن4��5J��Ɔ4��33�VY�0�9El�4i�z���j����d|"~:�^��s��b�Z���2����M����RJ��y_�F��iН|��╏�w�埕ζ�m�"�z]24�]�[���Ȣ酄jQu��)�yi��?_��omA�6��we�z��EN����.����Y�1����ТvT8�jv]�O̓�$.���w;v�T٪jT��z��P���=�P:mi�p�n�mMVjq�j�oD)GE�uz���uO��D᜜������܎��6|-P�񪆊�TiW0)��Y���M����dy���>�I��
"��s1yӭO{I�^����� �K6���:CP=\��WԻ�����:ƀ�5E,���v�]�:x#��ڹ�H
��)���G��͠�K1���0����=��g~��K�+=������ې<��:݀ͽpy���zHz$@:K�>8�L�1�\}0ޭ����L�|}I��hE���\O�T�x׽~]���ci�C��H�@;I}�ƣ{=S�G������<RU�ԯu\M)oӑ�xL&�l��T^=��w3E_I`ht^R	�n�{�~x�l�64�ESh�^�f�r�ں}#��YS��2cfq��a�_Cm<;gm�V���SU&�TۻP�ż������`�V�0�+[KK'"���+0�e���F:nV��җ֡�2]e�P�����E&X�}�-��ȕD���RW���W�u����F�(����_�߿���[������sͼ4�^Y�������0##)��z9��)�j�&vmoU��F���Q�V����r!�:)�{]q9Tfk���~�r�J�5aU���t�y�`�a��OЂ�ZjX(���*�K���: ���eMBњO`*��E�ս[�z��q�0D����n�O������n��Y�՞�Ez1W5y� !8�LK$���ebR��b#�����=���k�b�&fZ^6�k�\�
ׂ�3&=� ��y��%:N��:+�S*	*Ml�q���Y��6JXt�>s��/hx��e�jc�,�`�°��H�I>1I�ԟ�-f�ki<���ڹ6���Z���z��<�!�[w�P���M��pnO5:���M��C�r�蜽/u'+3a_V�*/���I�'�܌�	���XE�3�
5�����mt�s{QE�0h���97=�ڭ��O��2��c��3�qxwj��T������K�����P�^�CĔ�Wla/��ƇJ�k��M�ŭi�f]~����	r�
P�C�_{<}�.���uve�,��,���ݻv�e�φA��vWѳ�Y�a�r3�z��vM�i�5:�;z
y9�AzdEU���}C/77.���3tqbŐ՛X�Ў���d[X\{��C��K��l�/~��ml��W��SD����r�ڙ�^��p�7n��aF�@��E�E�w)섅Ò��Q���3��1�0+Jy�{q�V��D˩f��Ϧ�h>�5/p%Τ�٩�e��p��`� ����rS��L1�9 ��2�3�a�ncL ���s�1Xe�����d8�q��ڲk�sT��xG@Xۼ���lfnL.`P���F��)�I-u�j۩�bj��d��r�5e�5���]>պ��e��m���;��\�\i.���ӎ��{ǒ���6���-����LO�K�C��� �o���wY�fIC�k�3�|�r�!�������K�9����FEwjfE�-wq�YM�귢��F��X�rR�A���z���ʎ��a1��d�fy��>bV�J�4�]^-p�8:�flyb�%q��1����r�mf鼖/GX���ƅf���}�w7�淄
�3��{ˏV64�z��
�fг6R!�&����b0`�hkş`N����1gN؎��LA�x]��ٛ�X��\��q��N朼�V�l��4��v��[\줝�^}X𼁱��&��Ί�[ZzM��b��A���*�MKdV/�h��2F]swo.��
������[u/c���H"�c��A[����I)]��}�"�b�Ogfe74BU�cg/FX�c��^��\�n��oI�
`g2�7,C}���%ofqc�<õ�>�,α���T���U�{k����f`ڋ��/����{[Ӵz�.���@3��z�R���ؘ֪�Ȳ�NC�O\<���v���C�k1d��!瘝�]���{�	N�y��1Q����������Ĺ�=���{��(�l���Z��"����E�e�8Ѭ8��KY��)%�'F��M����o�ǈ�34�qv�6J7�5�j�ǖU��N�-@����=�e���Y���0�at2��X��MlI��-�b"���F�i��6�u�7�B�3�k7i��⠱�$R��{n�;����gÃr��4-���8�W[vxF��N��%嫣�ᔗX=�A���۾�L�|y��Wٗۜ��Cq�trQ���mQ�2E��X�25zkm_Yg��Z���e������C���֧���ۻ�h�4���I=�}H�Bn��՛쒸FUZ�bj�:����RӔZ�컵u�_{�Ŏ�� ��hVQ�5es���TZMQ.a LA�(�yS/[զ�fROo�TO��Fc�}�og��"ǡ�˪mfҼ)���0m^��*&�Ⲫwu�/T�4�����ռ� �Q8�� M���qN���i�ٓ��� y��i�u�t�wt�mu���u�vh3ؿF=��q;�pv=p]7{�oױ����Na���Iĺpc���oj�[�9���;���{���-��4��j�n7ln�rv�����y�={�w�G�������]��^�v��GHq���9��#���.7�1s��5�wh���G]wc��7`��=�u�uۂ8�&&���l���wۭz�Z�d�����2E�i::1\b�cA�*��{'��x���]wj.b(��\�4b7�ѳ�lc]F�sk�8����bC��ɣ�����{�h��q:si�0t'v1�DE#��]��q�<cTSv�X�vz�e6�Qv.wCWj�m�b�Aq��b��wi;�EZtt��n;�x�S4P�[��N"��{j��<O�^�^��۷v�Ύ��Ʊ:M;h��7l؍[ktPkZt�`�F���tu7F�-����I��wwfb������T���2Ѥ�m,$
�-��j���G���1F6�Wm�D0)�O�8͐m�/mEH2[$�k�e�9yVK���ru�'�2�&�#IQ%�ZL�N�$�E!�]��㫎����7z������-BP44R��������Ǆ�����\��hf\��0 @��T�v��zK���mv���a�Ʋײz}]`�W1n�������ۄ�ή��;��R�5�j`�Ã�<`�ŀ�t�^����v��v�pm9�a\Z��1\�aɆ�p�3����e{��o~�	��>�<3ǂ����"ac�R5����� Њ&h�7����Ц��]i��3��6�ڣ�Ď�^���l�wA���~g�I��m�9���evC.a,�
��y�ۻ}�Y�oK��{��eM�D�v�o�i�m��	w��
Y��	{�d\����l��\j̆�k�[���Խ���c^΄���2j	\����>l[-�Ο�]�����x���3x�P��x-.���p)�L܅я4٪O�xa�j��k��|j�aSr�J����#m��絻�9x3/`P�q����S���!s�� ����F�7��R�S�'*p�tO��,��Փ�cX]�eT�o��S���"-�
�]	���!ۇ\&��� &Iؼ'M��aP�Q�9թEN.�o8#Nӑ��f��-��c{�#���;�*�6^���֫2��ע���5��\ˍ?�Q�<8m�����*v�j��ic��"P���3{emE3v���h��#6���c}�:$h��xn#��ط-D�V�bF�*-;r�mB��#R����zT80����f�!�V�"�uiȘ�o8�q8�*F��� �b �)�H�"Zb}����}������_����{%���d�@���4|�pgӾ7��Zq� �cL9	��0��r��zZY~����S����O[�f�c�K�����;�?<�{h8Z�Z�RN��W�{�=��o �4S�/)�ɑ)�q�	>9+�Z�r�'���Ւ�xwh����@>��}G��s}�8�X#�O�ύ��`X�mEs�5�,ى:���*vZ��R�u���a���n��;�N�ݽu�z@���`��P2g�R9��i�jZ�1��~o�����	!o��J�#!d�>-7�y��==89�;��@a���F�k�����Ԁ̷�Kn�Ԩ��]dI��yR��
����F߹ݣ&������P�<�	w���	���~��,�:oB�م4�h�gF�c��|���N�Dėj�2�נL˱��ǫ���4;��|.�I�ͪ��rx��i��N@�7���o�Ȳ("h$��4��˴��n�16�ծ�ja�ƙ]uk"�ދ���(�,R�,�Ό��;�Mw��} \����5��t��#���FV�9�	���9�fԲrbI�l謞�9�M�ȉ�Ӽ륩��UdS�����p�[v�y��QjH�!q��u���'R�̫�6�˗��ɰ�ܷ[\I"��-R� �H1Vj���o�oj�*[%�e�K1���{X�8���A!AH�$J�B��)2��1*СI������������>��s�1L�8G0�a�q1o�sE�1��NT��JBװ0�2�WB���}5
>�ߑ�����'dm�T�
)� BcH�0Za�#���%0��w�!5���C�����Uo�sQܑ<�'�%]�,���Bf���S���,�{(u���s����ŮIUy��\���&T�K�&S�$�]��c־���=���ɒ��=�g_�aOzEؙ����n��0�XZ�S�脜��%�u�,1ijRR��p�]D�}�:��II:�FO��eV�0}���׆!�{��Kx����]0�#R���)������,F\4�C�م';�6��.��-��75�BuLx��a�D�q<�].q�?7�眷��0y�l@�F.��_Wa�|en%������#���֑#[�m7���1Lh:v�7{��r����Ret㵇���,S����T�]{�4�����W���= 8u�յ4��W0Z�7�Ml�i�^�6�\n���7{U0[�+��PK�<��50ur�G�::��QU��ƪR#=��|q�/^;&����D�N~��Ʊ��eUF+�(��������of��v��b�]��b�Gt5�w�;I�8�}G8��RN=g���6�8fK=��wQw�]��4j�-[�'a�2.h�c�Z;yu5�'��>`�N�]�r�\k���}+8�5�i��
�
�B,�H,J�A	H������X�y�������{M��T��	����W�����P;��hņv:w��H1��w�W8�I����Fjc�y�X��P���7d3l�I/�^=$K�(r��Y�!9詎���auҧ�;*�*�<׬����\LJ�/bv3],�c;����Hz$@#��`!W��0���J.�zvۤ����)��d�Q��C"Y�~hjdv�I�-{c�M��DVk�@���-�}p'rln�Q�tOכ|�VW�wω��]�p���CBz�sK�6FFS��}<�7&m�}I�H��p��-@���V�jD�k֦�&��V���3��cռ*���[G�:/1q���*�]Bm�������X���yMz	����I�Q�a@�^Vb��/�p����s���sV>���u>��[�$:����E�9�	�bY7�ZFi��R��q��\�Μ
N��k��IɅ~K}9�����5�͙0X��=�y��%:O�bS���ʒT�`'GndO�eQY�S���K'�tޡ��3[L%,�@Lpe��gd�q�&Rv/)�ߧ��-�yΊ��rVRJ]�_lsr��
ͽ+
��y`�c 9y5�M\��C�0�Ǝw�5S��ӯ%Ir�gL�]}d�܎����L���0-�%,�b2���K3��uu	Ðu2ws��ޗ�Suu/���O���(s�'**��UW��xiDJ"@bQhQi�X���VEa��_4ֻ֛^���L�k[\v�Hhy��y��m��U�MA���y�C�B�Ȅ����'��]�Ows�y�W��C<�g3���\�]q�N�2�K���:���	���E�>O��r9ĳ���:�ɑ��j(���W:�;�:Ԏ�/4H�R��wN}1!�U��F&��������'ol�?Nuî�[y6<JT)?_�H�Td�5߇t�喘4�|�}�Y���n�۳ ��XJ��!
�կj⛁�#�>�o0�s�T7>ׇi�j�Ja����x��WX5�JI���BV��ZeV�����]�i���	�1�p�X�!2gnlO�Y�r�]��� v�pl'3L(� ������OJ;*����Y~.09�2(9��S�&(:�,U׌��������s�pІ���Of��.�3��o#�șf�$.����9��l�wI�?�7r�"bӫS��彇�u�2�Qk�Z��+�/.�4���K����ޏ��ִ�����8����%{�u��z9F]�MvSU�f�+�+�b��b����fdԕ����g�׃��U`�/�a?{<}k�#A�Y7ꂭ�QϺ�3_����v5�X�]����RNR�۲��SC"��B
�J�Jm�(��d��ܭ�:�+��N�S�g��T��=����3�N����,�3+>7��%�[8�4�:oZd�ҢNk�������nś0Mɮq5�M�x�kjfnoQwB�@�
D*��1 �"$��J�B"��7��ι���b��8H�cvn��{a=k60|�\�at�qW��vr�Ol����6^���� `3�]z�I�1<�#L�&��%sߟ�Z�S�]"K��#��E�U��]fe��ZÚ���uEê��x�	�A�k��v܇np�Y��"�K�x%�VE�#�|��r���&B��U$��b�`�hUӍ��#G���i�82��v��#7l����-����	����mu&X�b�@���x�pgӾ[�	�#�!�B~oE�fb��]of�.�Aƺ��5��}�R�Փ6Ⱥ��敥�m�\���π8��;i�W�VTE�U?�Ɋp���t!�5cЗ��R�E�ga0�9+�Z�9r�ե%�-�a��ݘky����Ҋ��u���' �$
���Ӄ�+��KϤ�>%V��]<�l+�o�
���KJ����.o���z�:�����K����.��T�n�2)r�Z���+�	6�+U���Һk;����l����؜e�ρ�'��a ��2� ��*;�鱁�evυp����%�G2����L�dج��z}�'���~%�3�[o��Kj��we���zGY��ϋ�=ܞ��[�t�k7(^���"�˸26�MN�	`^���᝵.�n�Mٺ�q%XY��m9�4%M�TEb�bQ�ðr4ͼf�Nm�M�L�*F�M� � 	��1( � Ȋ4 �� ���դ�U{������D��	^�j��U,Z���轆s>2%�8��
x����?q��ɢ����8Y�I�ΝL��l�1@�Qo
&$�Q2�u�f]�{DS�Ϲ�����쫈kb�*��n)�n�3��XSs�� ��{2-����T�܌;`3�l���[ٚJR�����V��s��3!���+���mzn����_�׸MF}��U�C��3z�K�]��n����:����x��ڝ��7�"��OzE���y�ƞ�9R�[PԤ-|.�&��ud7W�!r�\��ҁčp����n�y�<�&Ƒ�a4�G;N+��`9�5	��QYQͺ���Π�� L�ʭ���vN�ϱ��=�� b�Bq$>P�	�����چ*oZ��<�C!IH���
v6��Ғ�3��S�]��}Ǆ��|w�!Ű)��-�۪�;%1�b[yd�0O'a���I�y�K$���W�T�7=s���N�Qh��n�wV�����p�s�ÓԹ�Ƒ
�ep$vW����E�7E2����=��7cͪ��_�����P��}ϱT�dp�����S��xp*Ԉ$��\�p��az����QdV����Xk&�{ѥS��hFc�s��1n�w[v�[�ƥf僠u�L�|��ɫ&�p�J�7���D[�kdѴۗ����DX�iT�P�F�R���ZhTh`�[���\��U��f�7�����@C!�D��n��B��M�a&��"�� ����Ê�U{h�3�[ܡ�S�騸�����{�0t��!x��=1)���g:�8��YuJh�ud���s�N���@���ON��'Ua]�Y#��Ӈ�p����Aí~�6��S�M��'�х��X���?Z���*���W=���إ���m��`�>�"Xt'���=V"݄<�k;�}Nמ��mxe�f\�� [+�I����Tm�鷢fy��K1�b�;0��I��U���;�C�r�ݣ���چNn�f��K���zHz�"��zA�[ f�46�d[ݳ�<�V��T*cB��b]�����ĩ��;�� Mx2��`�F^D@!�������v�.�ݾ�NʟE��"*�"Y�!	���9�h{d��T^=��u`$n�ho:2��f�]�
���lv�W"�P�8���w��\]���| u_����rV���܁��uD��y�:�M,��o�m�-`;��6 0��E0M����i����P���߷�疞b���q\㴼��K�6�0�H4KK�;Cwׂ�/#�P����j�ܾ�˭T���,���ond�RE��E���U�>Kj��.+9݅E���X�:<�K��.s7G�Y}A0����p�z�洩T�͍6XwY�!w���0�b�ҿ�!"V�FD�U�`��	�
!��> G�y�g��+��}�$�lX�9�O2}�>��`��;��"g���4h�'Rb�i�z��x/V��t����u�9VVf��}���%�w���w�q_5�@'�,�ߒ3L�R��`U3& ���˟o.��l�I�������Aq���͕+Ҙ<�4�; ��)�|s�_��ɼ�%��oEuNN	���R���ry��.P�� �5��JY��&82��v�z`�I? �m�n�k�'e�N`L��5$�B߇,�3�av��bG�9�hLpm܎i.˚Dd�f7��U);}���R��̅ �%���bXa�ӢyC\U���IF�*z������o[ݫ���VM7n�֮e�Y#YK�J���\�R� Lo�c�PeZ��tZ�$���Օϱ;Á�wf��J�Ru~5"��2k�Rr�Lz!\�<j��+b�b�JHp�{o�ͭK� ?@��(X>��
�;K��:�����y�(�a�ƲװOW���W4n����B�ʻ�u}<l���P�m���� �����azچO��C����a9�`��?�Y�Y��]9J�I��������`Q��(OpU�Dzd-���V����V�5 �/����0����A�!�5���;ۨ��&�	�(ZXD�s�ۛ���t!(��\/f-�R7JL\.�K7�T+���Rfu�˞�9/(h�y&�-���byB0}���  *�!���"� �R�H%,J�H�{�o�^%�c����8�,�gN��Na�4G3��D��;3���A����P��袻[�<I&߅x>�s��:/�pt=�`o�[]��8\sLL$�6���m�[��;=}1�4㕦}�i���%ڼSzm�j��[cR|�o~�{B��A�5k6vE;�Ȗ�<8,`���=�\���b�����������^H�3׳gW���x}�l���TovN�y��]��: ?C�=0ٜ��1��A	���a�-@�U�Q�gRc�d��`v�M�m\�9�l����\g@��	�d��S���!s�~�c����f꛺re5DD�$�Gv��uzUs
j=����i�$AoG�f���N��p�;%75Q>���܂
���lyӘ�����veRN.�8�@�h]{$��C%D��`��;?.>��r~vA���a��ң��`&*ۻ�-:�dp�6S��!#|��F%���gY7c��X���M��xG�W�S.�0�;*Jz�f�X�C��6�:��5�N��Ϡ���=^�o�������{��w�������^�uƹ�˲�P':�fX�k������mpJ�gYgi[���\Ǔ1�Kz�L�;��+w�C��U�o1��#�
|�q�n�WuԻ���� �w���LI��.a�q��H�sn����xaѐē1�D��;Ҥb��%�k	�]��a�������:�
�ŵ��9�Voa��\u�z+�����"�^���gi����	D�Ƶ�He�ݝU5��
��d9Y��m4�FJ��,]q�3mʂU����:;���a�4B5�-ɉ��N�:���'����P��0�m��í��m2�	�J���f�12��c4Fk���{���\�u|�u���D�V��ɢ�GD���3Kcdڴ�
UmC�u����K�{�!�����Q]Y�;�Ϧ���{��a����2cuS�b��'-b;s��C�UR��]�.]�ҬW��K���r���^cg5�|F�;��(/xnf^m�G*mu3���A:����w	�tnb�X`!Y�Ci�;� sU�HУҜӅ�s����Z����s�s��geo([���[�P`���b]R��5<G\6r�s�9f���mbݶFaŶ�/�k�\�qq^��P��kNS�Aߣlr5+�;t���'�:}w�eY�W͖o붼��{�^U�̶ʒ�-ϸ��OB���8�E��3�i�Ǯ�,^*%�K����#Z˺qJq�aZ��Y�ma��s���k<�F���ö4�x�|A�/3�8�����y�u0(Ф�ż��l^}����v�@RR�3sEՄ2u�j�kC�u�,5M]-�3�Mږ�~��$��YG���F	��1ͥhJAm����M���Wm���۵�6�
ʛR="�i����q�)*���j�S��h_��e���_��H��l����`�[-C�cQʆd��*�&�nAodXq�I��j�:�����3/f��oj`�1wR,��(�vK�\���y�)���(' �;-��.5՝V�*��!;�a�zD��WY�g]K�{.��//�"��s�˩EҳyLn�������"�'�kH�F-��̃�]4KG$�=�ǖ�e����/��Ī��u���4^c&���Zf�Q6ŉ=y$�ˤ��X�R&� �t���&V��w�Әʔ�\)n���u*��.�K� \�����k�f�J��>�����ڼ�iA��_u�[�ޚ�K�%�	�ֈ��RZͳ���^��(��^�*��mNג���G{�h�j[Y]�nH���3�8�֫�W@����o9����V���7O��[�m�睪���抹�Y�.Gx>��fofҵk.���+2���vU��e��p�b+��M�y�:�*�vh��5���:(,�@���xue�]�'���Vd�lF����[P�����ɶ�j�P�6��'L��u���r�[����&wu,U�j��"�P� {�Q�!����ST�[i����-X�m�Ί��)me��θ��늈�S�\�����L�TRX���F����mT�ZlFKcDo�w��TSI4C����E�b�".��h�m���h�EEEZ�kb�D+b�c$]v*����)�����+c��N�m8�L�N,U�8�c߬z)Aj͍Qm�&�6)ֳ�:(��:�c[m�EV���ED���+f�Z�j�b-�����j������M���j����٬^�մlj��cE[9��O�!���Z�N���k��?Y��VflmTk10V� ����譵��֘���TStm�kE3��DC1A�P@P)  ���_�}_t�̸�隃�O�����+ǣ��R��[���r��ٵ[��&B�g(�k�c��<�Wa��2�����|� 7��DhQb@Z $h"��@�5�����c&ԍ�����伧�]�b��n��]A/H%%�-�aUd>R��V���ve�{y��^d�q ��uEs���l��.�TXU��e8�:�xFB��ц�sܛҋ[����ؽ�B��4�?��>`����
�͵�hZ���\����<F��ѧ��Z�����}�����e89��v�@�+�8�9ͩfZj!���4Kvξ�8�f_8L�� �hO�Z�]�3I�nc�,�j�����-�E4���,�ȍ���ڶ_�ږd�߻����,(���^&Y��x��i:"����^F���-G�K�|�?b;�N�l�H?𬏘�ӵ7��󽲾���y([�Xݎ��
��O#.�tE���p��8g[����M�5���P3�e��Dd�)'�u�m{��9�Hxj���*� ��Z��TF?<.7�r:���Lϝ�W�����5h��U���
WG��N�۟��c߬���/zǔ���E��CEK�ilw^����
�bo�u��E0˘�s[��hA�?���*5����d��G�	���H�SU]F� x�MFN����xB�5��q�.��49�b�t�LY���5�%���c	������L����DMI�C��b�q�6aU����۲�Ɇ��+�^���h򼗨^�4�0�͜ݗW��˓�KW"�t��F��Y5��4�)hw�o��XH��Dh)��(AbQ=�3wK(J.�ss~��/��L��hȤ�%��]��ׯcռ4�E���cBq%�L*0�	ki;���:�~5�N)��%1�1)�Pw�T�[�]�}ɯN}�fT�O�UЌ�.����a@�
eψ:���~�p��^��|��K$���RJ�
~��[��[so�QER��{�;��O����y9h�a�'�	��r�.�0�o%��J.�7E2��D�Ⱦ1/<��A=x��A��d��2!<8zh\��k9��7vt�38��sS��-FN<�^m%xު}�&�L�.��A8�x�e�{���Bmj8G5�ėZjq�hJ�
;F�L��q�:�(�I�px�ϝ{O����pF�2�:��C�Z����Q�|�˕�)���cT|��Q����	�\���O)���K6�������]��k�
�]R3��٭��S��⛠�̪Lo����ϧ^���w%��0�v/�q�#lԭ�+�gxjˆ@x!�yO��j�n��;���Q}�Ǥ�!���x������	�S��$���'�:�+7c���gr�	T�g���ݨdV��J�7�f�AyV�VIF�ʶ�w.�ݜ�+��b��F��U1�v�(,�y�������xٸu)|�S�Bb��z�n1H�a���3? �����hQ��R�,�u��zj"���p�4��wk��L?����D���;��A�+0&�]�]����m��/V2^�F�˩�y�[�]�_�%�<��҆Ai��I��Qx�p��!����E����jf��e04
�r��of���o:��a���	�FFS��֩�h�|�YG?/.1�3m@�T͸aG֦�&H܇��M��X�dS�`qm=Mt]\���+��s\]FǥT�cnv+���%6X&Pd�-����0<�o�ޭ�yn��Z�Z�iĻ"8r��Cq�h�an��{���EF*��A8%�~Hש�\�I�k0�-a%�.�%�Vf)�νY�l������{:J�.͔}O�)��cH"{$���Jt���uy�e��o��^��5�V�#�&�����@�5��ۂc�)���I���)P銫��Y���O:s�,n�Il��	�.��}��a!��Bm��ے��0)��a|Gz1�_)j ��/����zO�����<�F%���-��� �G��%��n�U��kS4��c=��W	+4չY���H�72�F+k�ul�FS�IV�U��.i]��m����������{�����B��Vnӎ�^�ї|�l�\�u[��+Z9�OQw��X�᭠�N� ��Fl�K$՝j����팕8��k9�����  0�����<�f�钛y`�xe�@�xղ�Zk����^Y#YK�Q��1!�wו0�D��Ķ���^,9�ij�B�!�0~�vK�ƀ�\���Ɓ�X�}ғ���ɷ�\���6(�{n�X�Й�6#�-w$��>񙈿:�C�A�y�;k���ϴi�j�JaťG����Cϙ B�3O����a%8ꇮ��d�B�C(p.��Á|p|/B/�gt���.P�/@��>eT�mv��D��sQ~�����xg�"9��(-10���H�JN0��<!UB�բ�18�|�C��D�ba����$e�sͼ��8����Q�[��xK��7|�=��^Yf=��w��2ʹu��v�9�t��m�ִ����k�Xɘ~��7꼣}tbc/R�����R`��	��c.y���i��ⅨA�W�W(2F-��-���ʞ�펺�)�������NL�dW��I3L(	��M�E[W�A	��a�еY���{w��{+�q'������0}�Vܴ�#�m������ůZ�ώ��?B�������-¢Xp��Γy>"��j�ֲ-���,��Sa��q�;�S7ѝH:{�N1Qr�6�m�c��~�h�o�KCc�6���\_DeȺ�t0ɗ��b�dU��]�s�pǐu�A۳\X��&�܅ݥ���t�µ�2,na�h��N��Ά�ޯ gq={d��︽���R�)����8%tV��V��K�^_���k���rkM.%]Q��>���S��~�q�%Sd��ħV��j��:q��E�*���zA�i�:A��[,u�wX�V�����m8nC�݊!��Jb9�n(��}iA�\ŗ�|��K��x�ֹ�r�b���8�0��1����p鿙�q���!�RSՓ6Ⱥ�09��K��=5ϙ)�K#,�l��]�����Æ	��9m=à��Sފ�6o(Q�v�
�rW<��)=XJK�4�sA3,�wEi���}���
$�pߍ��ÚU���TW:�YB̓u��%Qa�^���ܳ��p�ݶ[��󅙗�<�vT`s�&�����DsL������ƇT�m�OQ��Uvъ�o;�J�g^n��q�\��%����a'�N�{�#�0~�g#a�Г���ᥜ~w���vs=��h���J���5�c�;N�5-�@�/^/a�ό�w����ha���N��p�u�x�Ojg�����3i;�XQ1%ؔ��T4k�S.ҸE��Ο�^�n��Ȼ~7#�Ԫ��)֨���xѩXs)\��x� EN���tM����[�m`��FB��wT�ߒ
FD�3Ҷ�J9S���-�xQ���@����鰺C�n,�%_V�'O�[T{g.�*9��E�͗�Yr�s�هG-L?�Cs�ymr#�}��|n2��m.��jP2+�!@y͊�����W���FdYx�Hr�ˑ�mзnzL�bS]����%�m��o`38:�B7�u@J�r�ei��	Q�&���`�\:[#T���%�wվ�ѝ��<<�Z�<'5h�9@Ue/�*�?�7i�[;г�����TG��0|�i-y�����k֮���ң���M�T9�n�n*ǅz�P����+�u&��^ϙ������R�X�x?!)�ɐ�P�hR{�P�ј��O����>Ǆ"k&���^b��m�g!��	����6�!)�/	�Q�(IP����5��E?IRX��;�l��i�{#�;�-���@L��hOa�wD$��E�n�d���_//
꜉���U�}G%�i��ïs�G�(f�t�s��ݍ"U{��<��]0�#R���x��c����t��oj֤0�C*
9j����� ���p��S7H�4(���"��qw��o<�6�ɜ���e����wJ]*��ƙ*�Uc�����A�:;=�Ϗ���쟾Ϝ���s?%A�Dgo2�B2��D�ݹ��A�2v6b�̡x�V4��6n��r��n[QV���䧓j��đ���{+I�Pl7ӷa�fu	u�R��y6-�L+z�0B�)����U�yZ`� ̩�GU;mm�9Je���C8���| ��vV�w<��ݜ6fE�T*�<yK�{�]�ʌ����B���s�q�Z\K�(xR��@u��ћ������t���!�{*i�B��˼�V0'�k�I}�n~\}q��`��΅	Ge���`�uU]����,�^F�ȇd�d�6�׷�+2�1��:�o�gӯ@��j;��nt��G=��_^,��7��;F�f"=p!!���>��d�^ݐͳ�(�X��ӝ+�Z�u�}~SU����m-��b�^��mClC�OD��X@��\H�Se�ӱ��`rh1����5hU���	Q�ݔN�z�~�'��~��:X���EC��,�� ���2Lo�'�Q����PpO������~�B�wq�h��,t�r��of��E<5��<X�iiABm��/ �r�ޘ݅���T�S׎L�U׵�չ26��&��P|U������\���
��p�4T���y����D=󽿠ܪ�oӱ^��%67'�bS�Tgz�{ē����k*��2��9�/��B��[�D>,�A���?B	��=���d�^�M7�M�U�f#�z��F�y$�ܽH#�k��[v��$C�GPw-��d=�d삛o��4)C��N`b!�s����	Y�i��J�f�����V����0o<���َ�eL+��vn�kx��f����X��B�ٺ�&��LT�nS�n�x�W���c�}� 3�6o��ݯ_������ ^��ȧ�x�$(���Ba0R;A���{~�N��+�,�Z���QK.���9q{Z�S"���y[���fǨu�= �5�z�m���=�.�*Ԛ&fU�?\�h������o�����E(t	K'�kw=�#ϲ�lA��:m���]W�ll��kWv�pڽ�u��j�n��M��1i� �+����0����`pV_)�i�ԭڍ�8Z�P����%��Ji��Ms]��^k�$k)z	Gs�e����1.�h�\�1ǆ�[6��=y�Mʙ�"*K�y�;'�C��s��E1����fwRN���d���\��+]0/��n_w��az��{#ٺ}�����?���K�>�i�j�JaşYc��Rr�e�PU���v��j���y�8�/C�z�;v���΃� ���^����i�.���0���^"����C��>����t��m�c����v�;ǴG3�e�%�]k�n#:�N���mգ��ϨCq�!��-�B(���D�1i���Hﺞ3+�����L���!��>W���B�Q������QU9��im(����	[�tho���3]�*U-��Y�bHЙǕP�S�Wr-M;HI�옎���e��H4Ȟ����}}�V��i&��ٔP�[n`�Ť�1�)Ԓ�^����\���3�Vţ+�X׶���u\#��~����[W�Ǯ)!��5�=�_�N6ۜ�����(wI.�E2ˡ؋}kO��c�kI{:��ki��#��{�/af� =ŷ'�Us��ݬia ��Z�W(5$g�Z��Ĵ�v*Xr���,b���t�N�9�`r��>c���L[�g�C�!w��K�OѩnZ��g�UV���@��#Ռ�u�6K�:��̂qub$��6K�;V�Q��5�3l��PWQ��`��4���+�蘤��
W+=i����Ʈ��uo��"y9�k�Iۺ��z-qx�0��)a�=���؅JS&��$�^�HеbU$�ߢ�u�4-�ot��[o�C���썚e�ܛyd�Rn^��6�D5t�LPc1C�Jt��s�_9�o ���HZ\
�t���xx���6,C�Ϊ`�=�%�v��ʒ��6Ⱥ��� ��x-�2{�+��pS	�|�r�M�,�^w�|yp��0Z�Cw<4'�F�i0�8�M�-G.Rz!�{R��u���h�o������E|�Iyp���-�\@M��uEs�5�,�1'\o�_O����7Փ��f�ax������6Ԓ0½�Kkm:��-����3T6mn�YQ+���5̭��t_k��x����LT�P��g6��b���7i�L�jmݜه��5�=Ў�{���x./.��¹,�y�Լ=f��-��B ��ﾮM3��h������M�����Kݾ�sۇ�p���>��C��W���!��6"����/��=X�ڇ�q�-��<�Ԡ���*�r9�0L��+蘡�S�W0�V��:�['��g�_��<��,�h-�Ú��@��}�Ӵ5-�G�az�{=u��潷Z^V�}��鵗ө&��r��[w6���-��w�7�,�'r�^��,�^��v��/���8��|F�cN{4��Q\J�}�s4T.ǅM�y/�6*1���v�e�;��T^\�f{.$�O@��D���tǾ�+c�'f���gРJe�Fd��*����Q�&���B�qQ�g||���s�Gp�D܍�ךn6�5��u�,�������J�ϋg��P�Z�3��-�<�ȓ!k��2�Z��*:��oN0�su�Mm��0[/�S1�lr�i䣙���t���q�/�����F�'�G(]��׬z���Ol��X&����t�3+w��_C�e�%:�逈�vW�i�b�j~BSc�X	I`��$�i�W6�)�1�V�[�l˳��-�e���w����zzz{�}�^[����O�<qԚ�I���Y��$��zm4�1ux5B[(a���ΪS�PB��۶kguZ�:wfg6�dˈ�&�vC�m�@ӭ
Ӻ݂ӣ��oE����ۮ ^F�+�;��>�=�y��sk���m��Z�[�zYpl8+L�7R�e�1�p�i����ɹ]N�=��\B9eY�$���92j��I\�`F��1kU��1�&�v���r���&����yvr���inb}Sba3,��Sp�Nu`d9Bq��9�u�U�#��$=��ḣ2\���po��nԝv�S�ٺ�b�r�����V{5;��	+t�u�=��cբ��gj�KmfA|�Y��:���'=5�C��w:Ʀ��g���{������d��.�-U���umB���,�t&�M�Ne[�\�dxf�^d�p�x�����uwRWr��o/��ލ�{8���:�gr��-�9�����o�sΦV���s��+������4nAc��[����n'\�z-u^�DemB�KD����v��ё0�����-�ڪ�$tn2*�uV$��e�u8��	XeT-P�N��d�>��A/t�2^�_k�r�mZYJ��Ot�C� ����ϫ���ͻ5d�}�L��nAٲЩT�J�b���ۼ��{�f��̩(�v`6�Z�=��/E˙��e�Xx�{�P�����.c_��x
��X���_��oJ��8*�:�H����#7nķ,��r�Q��d�S�M�eR=���y��	���bj�"��.�]g9�>oV�u!�(��A��Е�����ٵKfe�MJ�,l�)-q!M�i�6��,�n%zę�{gQ�~��Q�'�n婢a�0��.��2�U��7*�X-b�AY���|�@���q��JL6u�u ���cv�_Y�c�ئ��u����F�N��@��ʒ�L�j՘%��lc�%����r[���7n9c_H�o,:�E[��b��mc/��/�^�	g^��)<f�R3k6��W`,9{'ݒ�$�&��d�|S���,^��.!�֫8��9EW� ��
r�晲�]j��h��h���wiYX���R[�R�����s�u�����D�xE��w,��J�w+t�}(����oK m]�
* �C��,��ma;�j���+�}�+V�w��`��&t�(���Oz��hD(��s�����v�ݵL���4�a�DEݝJMe���0R�j��`�|Dx_�9{]c;D��vo79YmB�Q7���C*!���̀ {o�4�Im슲��~�bjL���[��zbv��V�;ӧ����,��1�j!m)6�ӷtu��sx��%�}Y��ؘ�jgw`S�;ޮM�������u>	�7C0��3����l���bl�j�X�m!��{WyW�IV�^ܻ���ws���n��X:5h�m�ʽZ3��)}�]����&���(
 xPMDà��b�(���GF(֒+[[�=������c1��&h֪���b)�uLA5�`�V�S��T�QUAF��PQlfJ��)�5���� (-�4S�3$Mkt�*n��鱢��֣F5�I����j�Q��E���ͪm8�I�
�&j"���Sg"bMb���U[fdڭ�mP�]������cZ�10E�"�j"��ٶ
�ڣ*�'m�
�������qj����F��lF�l�SF#4�EWZ*b��V�",�0D�UE��i�ţKU˷v솴P��'��E�Ul�j�6uUT6�Q�:]F,QQDSm�����QDSu��mj�Z�E5E����DPS��f(�j�����cTS4�kU&	o�������G��-�I����_�!SExy�+���ݟ0t�g[���H�Jr��bSA�XP���5��s��DF��m������ޔ�ĺ�v�I;{��Vn�K�*T��V��f|�۱���ۺ;ֺq�m�WwZ��6�{ǎ�%M�u��>)'�S�. �9�?��;Ǥ8��H>C���h>f�}��I�/������t�Qv�Y9�	���R�9���s	����$t3d�O���s^��q�J�;(���.�\�E�q,C�Q]9�[H��cƎ���9jw��P͍"8Bn����v[��<+l�{�C�u�[��É]�J^�E��I�J�栜K�{����M����ǜr����ډ2<�_�Yjj�hY*L�YΪ���s�Y�|^�M 	�J�30�nx�]Za��!�W�M2W=I���U�j ��Γ���ep�q����[\otL�s�I�MoUH�^�Kr0�E�C�yAjنn׮͛c`ʤ���S�z��=:��ssqt+{,�3��u�E)�w��臓�%�{�3 �<�]�5�xmC'�ݐͲ;%�/��S�����C{6�1ٝ��O�-{TP���y7�2��vS�� �h|.Y|Q��`�bU,��O|n��V����Z���\�y��M;H/����0�y�BK!�Yڇ���_���0�p�u�0���M0ڳ�,Q�Hq��x���em%igW�I��Ym>:4�ǅ�2%�V,�j�� _xvP��]� >�9�ʙ۶�]��j>��+ۄkJv��囦έr�b�r�G�sSʻ������M��J�A;��74M�����	MWWG�o�O��Ɔ�� e�4_I`h���w��D������E���)��(�B"+�j�W�m���-||�39�����3mZ��m�a�Z�`�R9A�ٳ����u
��ik��Sq����*�nm����*��W;=�D&�����f��Tg_RI�S�u��[�s�{g-ս[�z��t��0D��p�{�A�����'	�d��7pf�~B]��'y�޴[���b#�����=�Ǥ!D�f���`�v4�'�O<g;F9���\���rǚI?Q�sk��P�)%I���9�>Eê�� �5���}ڎ�m��ͅStN\f����(`V)0�}��$��*|!�E*[E�5^��}������ۢ6�X���
a�`䖤����������2�K�ҧè#4������y���)�U�;w�Av��gb9ňxc�Ck�����5�e��5�����3�irb�z��y�bk�X��W�3_�`R����C�~4U
���H�4d�5�/ߏ�ˡs���6��	v�'����]����\uY�vC�+2ô�j#aK�2�%�Ѩ;��=�걻<Mm۞�Ѯ��$)͚��X��NQ5���l,�K�{i��іլ��8��Q��ji��X��d뒺�][�2��]։��{��b�b"�JX]
�   ��M.�}�Yq>U�1S3�	q?Ex���ͮ�綡���i�j�Jaï2{�Ȕקn�A���\��{�O����sO���Gϥ"9�P�kh�?Q�>���͇������ث�q�p����!�<�s4"��sP/��j���a���\��w�kG�u�Q)�y\�t<���A�4"�3Eؘf-��q'EoN|��k�X���r�"���N�X1��"`�=1m�뻧���4��$�W��d��˴�}kN���E��E���V�7p�܍U���N�9�R� =ű/~���u��Ɵb���.��	A�l�i�W;Wx�r�vٶu���U�6%͹ɚ�G�'ޒ*I���gヸ�QX�9G��ZSQ9�V��=��"���0�I�g�o�C*.��ft��\fLO;H�:ɫ�k�Q�T�`ت/��-��!�s�}���(���(�*�
j�q��k.!��g��^�2�x�pq��'n6�gv�����˱W�73s�I�=�v
�J��ʤ�[�[�hUӍ��y��#a[��Qv�����5a�j~/.; �B��ʺ�~��-�e��%�8b��+���an ɩ���qp�ooꋷM���$�4Bw���L�ma��S��4ș����X�q��LQa�څPA9R�L��m�����MMQ��C-�[���-<��5�(�QcE���{AĈr϶�ۃntCg�uL��`&(t	O�&`���l3���<���:s�wqi�|���`G#a�/�0��ʻCO�*Jz�f�@���7zr�<gq�od�mթ��=����`��r��^S��B����U��疩�!��.S5�����w_GJ8����Ӱ�'�vh܇Ǘ����t�����TW:�YB�E̸�1-�<���ks�[�Cw�0�]<�o��XH/w��k�D�#�8�Tt]|:�+%�7�
��)���!��9�^1+�Nd��J	{e/�4�:��a߹�
#��[i������߯M65{U��\^Ǩ>��f[���sQԨO�Z���I�nc�,� ��sMM5�cM�CT��wV֡�[��=��͌�f)��K7Iܢ����L3v9&e۫��sk���B�n�ޮ��.���C�	�g�F�
����lǸ��`W��ޚ��w	���N�F�U��ٞ���42���=�-���6�ʶ3����E�#2R{�T^�Ղz�~�/��?X�Tf��yBs�E^[z��B*��ϨI��9sK�غ@�V�2�ҥ�W�lcr����I7Xl��t�u�U�f�<2��a�V��E�jN��H[n��zX�̭���tƛ���s�Nۍ��p�MXi�p�TidP����K�#�K(;�L&�t��!^dM]�[Fy��Hxo�!��r3�ۍ�M��ޘZ�g��"úP�$��Dyp��V��s�������R��yHZ�]F�ХiQ���.b��ؖxBkL�Ds��+-<���0���8b,��'i98ˣf�_���~&BehȔ��Wlf9ǫxe��Wt�i�Ǎ
ز�КG8��s���TZ�s�Sc�%�c�IP���� ��;5Ҽ7S�x��p���Cd�Pp��#��mWW�m���W�۳$��1,X���j���}[�S赊~Q~�ts�A�uӭ��A�lwL>K��>�i��0��n��Ml���i��Q�X"jSm�cG:����;�׏8zhAC64��	�y��;�J�"	�*��|g�^�~�QNt$�4a�Q�].q�?2O��t�~j	Ļ�l�a�6�9g}�LDK����/�<[[�XR�s_R��	�;B������uV��z sIzp���I9����W�-�H�h����!'�ښm��Z�ά%8�A;+^������?}q�����~�y�+]���X*	Ǹ�V:z��sH)6��.���nRW��s���p�[�x��/:�kE�WSZW�/-[��]�-��m�����Ot&!��O�����@����56w ��.%y��y���YϺ�­�Lݼ.�!e��]իsUOUa��.�P���}�Թ.�ex����@�A�{�mt�2a�q�s��Y�I��������i]�]m�dO���_sz�g<�_d�w=vX`38�`>�E�Ѿ�w�*�=-����lߺ^C�=J��U>��}��r=�9lHk˫}�V�C�3��,#�C�q1*l����t��>J�oW+a�X;��|S:�h�v��Hz$@"G��v-���6"��� �xBKJ�;D{ޑj������~�O�,ώ�䞑�۸i�*�KE](r���+��Ct�f�Kk~��V��s{��R��kb-�>=��S�/Crfڵ%LۆdE��	�7!�f�'��e����Z,k�o{������
�N�qm���ǧ�I�`���{��MzL�ɭ��y����f�WK�lsᦫ��L�|mwA8��%�Ȉ��[ ��<��)����5g1��1��8���=�R��~��|njgO���A���K�eL&���Y��1���bv�oU�Οby�|����E2�$�5���6�Eêq �5��Rͯ��z남3m�AQP�Ӌ��,�)H��65
[}�^�)�F�ħ+��|�f�x	H�<J���N�����u+2�&]n���"�*eܫ�BDlR8��[�Wpn6���5�4q5��.�9���^;��K鳻n��Y%�wF?|>�����L-���1�� ��8�)?9�NP��m��c�u�GPh��C�&rN�B�,4�-�`�27%5�uL4���.K�~A@�t4�^Fi���l�a����;�k_��?0���4��8�xc�[]4�}����"�|�|5�� �w;�i��ٵrw]_R6�%
�wh��v�6�w=�v/ƇU
�VH�4�ƾ�J\n^���vl��7�[�e�d.�����02W+$u�P��U
Q�DUiE��k���b�P6�l<�����W����-x,���WX4�������;�X��p���<P�Ŧ[�l�T�W�Ю�3��N�~��M�Y�N�N
n��ؐϻ�gKz0t��J�a_�����b�:��6���R����퉩�{J�k#}��A�4"��.�	�b�\��:"��E<��L�����շ {(��xmO�*(�Qb����^6ۜ�Fe�f��K�6�5r2�ԭ���v�=�f�Vw����o6������N���K֊���r[����Ƒ�,�[}~J�;�T�ңy]��/~��	ޖ��%*v��8����h	N�/�QޭRk�qP4q�w��ü-^���5��v��Y,�y��d�:�oE��cs-P�	ŵl�t�ؾY�BKڵ�m�����N�������N��И�4>� �yם��}��g���޻�D~|����Y�ddO� �ᮭ��Ȗh.��f����N���螦{��F���V9�0�z�YQF���u�5��so��h(a�̘�v�U��]�,��yZ�C��D�3�b�+z�A�����4)X�H�ŵ��ε��ڵ�։�	��vҪ2���~�n�n��L$�q��`�����	�{�Jui�U$��:q�c�B�tMC�#�������!��FF3�!ñwn]�4�t�H�I�1����mi�#���Z���+V�<�O^q��Y5��}�!4���T�#�{ K*�5>�)��3l��ʫ<���x�6+xk%��y
��oWEyߙ��ك�Q����/)���4(���`t�!S�,j�S�Ff�-/,����%%�;0�Bxwf��|y��l�t�>�	��uEs���Y��i�0['w����:�ĝqw��Qak��I]k�O�������9��	P�g9��~ۊ����r�=Q~9c�Դеj%k���+�'%�U����(���B���߷��}f �㻣2T�R����0n�t����TSq�9��oC���/2����/=u�s�j5��N��#į($¯�^��B����y*�6�����w���Y)��5��b���Ew5Z�>wS����%�ܛ��n����ʩ���\�}R7��$=�~}���[j{�̺Kq.i����:���i]@��DH���>�%Ou��M_�sQԨ	�k^�v��j[��/���D������8�g��w�� <yL!�6߲a�'G�Y�|w(��]�1��0���3s �K��KZΘ�![C`[?>�;���^a�>0��s���<�MoM8̣zW	�Ar9�:��_���#CI&]�l�tM�1�����j��.'ѻ)<��=3[,\��c�vH�>���yc  �A��a���B��M�ۦ�t�îyg�XG�:N�&r�g{��*=f|3)�{l��� ����Z�%�ҵ*:����g�b��YU6�_���w�4�Ҕ=Qp�I�T�.ӊq���KsS��,!2�F�'���s�����j/ۙ΢�'1�m��-z��s�;p/l�A{�0��;�W������RX&a��v"c��׫�G<;2��A���nqJ3^��3�[G��*`������>�I���k�;]��Y�':�#�1��g����6�k���N}���a�$D&	��^��tC8�%G��ӄX�W^�wiخ���H��v�Utv�S5s3�r�5�Ɓ��&����z�ڳF!j�7��&�1��n�h�31�Wvh���wo6m��[�Ѷ�$�ʗ6��A�۬�[x}J�X�I�Z���͙ϖ�n���eR�zXi�����LwFN�|a���L-�]ye��MCu4噃kۇ��3cLp�ܪ��y��I���ݸ���a�oö=J\E��^�r-?5��ל��P����]�����	��r��M-��^������ħZN0-@��J�.B��uV��z���zp�v�gu(G]^�ޖ�!�")�K�@p�\�ڜ������V�V0�OJ�%��إ�X�0ξ��s�\�OV�j���l��t��qy�;k��vm��Λefw��E����vﱦ`^����T�[��r}�Wj3��G�uh����,u	��t�M�=:Tz^%b��T�E	lϘ�;����K'U�e�tǤ����D[��Ǟ�, h|.$D���ar\^���w�g��߮_N~ݬ`�#�	D�ON�_E���lEC�{"Y�- K��U��[G�Kzڬ���ֲ�>2OJ�����m�R�}%�*�!�9�=dRt9���Uj]0�J�9�K�ʶ�D���\X#�Ŋ1���T�y��fڽ�*f�eU�Slm��X�������2�˫-�e�Z�ϧ����������f�����j�c�LYJ�)�iuo^�����*��ł+���<8

wxG{۽�^�M����q%en梜�C����3PH(3�U�V�us�e�ub�����.3:���s����檕hWm٫�u	��>r�R9u��u�����/��;K���O8[�c���s��O�ι���LڵF��\��q�6�����uc���YB��i� �s��F�V�,�<^��o"2�Y�0����Xr�Z�W������Fw55`<�|�8I�RZ��ݡ�o\��j��s0���-;S��^�w� ����쐛�V�:�"ߛ�N��+�#s9�0&���T�c"e��^��$re�Ν��
���Ukj.�+V$��z�aν�6���e�c7��F�T��q�OI[�L���9������s���uxM���1y�E�ם�n�}���|�]������N:�զ���+3[������Y� �jU�ob{�3��jt��"�֔�6�e���]t%����Q��n&�^0��̦��`��v���̧D�ۉ��F���HJ:IS	��E�,��J�1�n���:�
���2�XУ�0���̝4m�����5`mj��l �GY�*K�L�;�.��j�'���[��X�N4L��S�,�iE&Շ|��K6���[һk�M���u��XO���<֦��;�dȞh�廖�Hƚ�q.��E\�9E�n���Yu0(��Ik����Q�����+~�0���J�Ze��Jv�7FS�1���}b�'jđ��-�����"��AGr�����:pJ�[���=|sl^t�������q)�Ԣj��w\�W�Q&�3�^�FJ�f�D��mG�)1���Ů(V��P�;���&��2���"��kR�%]��sS�]:�Q�B�>�JAón���竪Õ�
=z/wL���q[�\���|������ܭ����\0ŹX�яy$�!��bmUNFWh�wQ1�6�]^W"U�SI���e�g�·Oj�y�Ի1�3��ʌ�!�8��v�����i�%� �[iĊ�=k�v�V���΍eX�`u�n��i`�Ypg�-"Z{,^ގ<���@զ%���6ōj�i�[7��
�ɯ�d�"CoVJ��^�i�Qլ��u�8�\�\AY��[��Y۞�k7y��ܒ
��^���moj���i��.��p�KwL���F���Y�@vn�������,StY7�[[�]! �
�7/��+o~r�j��%�k\�)��,ܝ��[#�Z6��z�6:���W���6��̱�=���n	�W1�<6�o*���gp�W�Xݧ�r��c4�(kړ 
���rW)wY2휐����l<������f��dZ]���&˖�����s��2D�9�'yd����|H�O��ݫkY?T���󳸌�(ق�]�ɭ"*�j�N�ěcZ����)�߭��ӝ:��1����:*�j��kAC)�Ě1h�h�LCkQ@Uh�hr�jJ#d�14�����l6�*#Qhj��F��-6�ED;&�h�)*�
���l୵i1TUSU�T��SPAD�cmD�V�"�����
)$��h���C0WF(��b�Π�
&ѭiucQF�U��T�=�PTA]jJH�֢,cQE1�b�t�BS�AUF6���EQ]��U�g[~���F�*%(�m��E��EU��EQTMD:=u=���v�b�h���]V��m��[8���Ѯ���TA��(���i���mU�����ғ�cF���*-����`�V-��+[&�f-�Ψ��b-�A:�DIBh��Q��:�%RTQ�EZ�F���mh61M4llI��E��o�O�����M�l;u�2C�N�jL�����k�9��m�Y7y����8e�$!V͗�u�$Ž����BV�j��L�]f�l칚'˧"��c&h��a�y��OW�V0J�b��D&�&Pd�c;���j||Oq�l��)��; @�z/�oV����/K��HyV�ႏ��g7�a��]�5�% ��N���q>D�2Oa�e>�IZ��ޖ�Ưi���|��?��@�T��_��"�av����|���I�9�N��ħV�E2�T�����^�p�= �5��01��+&�M��o;f�,Ԅ���`��q�&R~s��м��'�k	�.��}*.����iW��E�m�����!�#���T&m����TCT��b~�����u���wF:����c�楆�M�-`����[,kL9���k�]^�`:�ګ����Ad�e.�h�I�[��yʻ/{�S�׌��ݨlc;��0~�vd�zdO:�-�5�f�aۈ����dϝjT��ˤ��]�~�ϠU,ٯN�ۃa�8!���^a�]ǕQ�>�W<㸠�O��Lwb�k��
%0I�Yc����j��u��uv���}��<1l���;�sL��AuLKFX��з��!���X�(eL���lc71�u}��9A�٪yu�*�����B1)�P�A�"�^T@�B����=rɶ�J�,�/l�]ھk�_p��[x�*hQ�p^ࢱ&s'a��R�ҳ74�3�o
��Σ�N�{:H5]�/"�'_�NF���(�;s.���ߎRN�3L8���LW1n��tL�j'���<b&"��ܾ���%�Ӣ=�0�OD���ye��[�o����j&Y�qr�3�DY{v���!���r����5���.���2��0S��T�m���>�fY�h��5�a��*q�b����h�i/Ψ��)���N���ּ����N���#C�["�U����wV��P�p��F�����ER,l�lr!���42L�=f�2��-�<�zw�\fI�T�9>���vK�U2;=���u녽ј3�k zO���NE�ʊ5��u�5��o9�\gA@ɱ\d��:Rp��#\15gI]��BS"=1��c�+!s�~�c�1I��4)B��Ymŷ�ڟfу�F�t���x�eng���J
ˡK2��.���v�=�����2OnbS�HеbU$��GN0g�j�	P.���t�l�V�h:ށ!F4��D9�n]�4�t�Ou*L�0a�E'��=0���\��˞�_WfB��vl���"1�C�
:�#�F�ȦW�K*/�r�ӗ�����	�d^�]�*�t��ǭU8��1#]*�j��ma����m�i�ck����/��r\v��br�=x��^|YGv�[u�N� H�mC���!Ì�c)�O$���I�����!Ysv�
�G:%|�ܼ9ً�	�/1�����'�r�8gM���#Wki_-�++lUU�1��r�C�ZN��}���zw�~y�p����z�����4(��ީ��F�c����'��PYr��PX���0���������+'��zM,=>^�\,�斃֨�f��55�F7��x�ϧ��a ���W��2�B����To&YZ�vLOp�q����[kʤ&��P�j%k���\�9/L���m�֠���Ň�S��=���S��F�O5@t\�گS���Ú�u*7Mk��C��j[��i��H�<=-�ٛ��|\�:z��uoa��;�A@x!0���~�2��'W�,�#�r�
ė�v�f�r�Vmq�J����A�=U1�o}1�����.���:�B{a�f��v�zr>
hRٱ5��v$��9�����O#.�tE��WE[�`3?�>B,��̔�n+�ѐe�Z�s�}d3�Fd"��.U@#OO���M^鋇U�L��XR���r��I�VU�8-.�4��TcV؜�kj�d-{�A�WB�Rq����	1P�=��ds֜	���'~?�#�c�H�'�v���g�R�3��� ����!�#I5�.����\<�]��/"��n|H��l�+P��bg,,�؆���{3v��B��ŝJ�r�z�`+�oP�V�% �&r�>97���N��[qnۧ�ἐ�vM��;2���l���S��o�L�S����D�3�~v�b�d�NԷ5,\Jl�	��U�B�ؔr��V�5�-��5?�oN�&�s������4��!Ol�t[O��/�&BGf��CTb�j~BSc�EY�iܽJy�yV���O3�or�V?y}�*�k�2���z��Qr�`UEև�pB|�c@"{zL��λ��D�^>�[����bY'Y��I)L;����7m~2��^u���+���;��Q��!˲��0�7��\�QX����N�Z5(���ʖ���0i�3װ�� ��#scP!�*��m���	�N��(qG���O�~JС��jO�J���v:ϑ�n��Za�/r�Ʀ�!�����sf���h]�Uz#��_���z sX�W>�B& ���՗�\>�
��4	��H`��������`OQkd�M��g�K�}�]�ܘ���v.�K��&ɲ��Ҏ�8�uK1��l|��A�8:ǈ�/0�ra�d�s��X2�1���OQ�(��������t	��w%����͆v2`3p.GE�y���/nY?MF.���` _�\2�ϯ�Y���c��pfpØ�y���XQ�{Qѻ�"U�p�LK!��
O���8S�]jgC=��0�led�5�`�9j���i�2\fMi�2��-<!֜�Nl^�j�2�c5F�������ۓi�j�7�-��xUn��h��g��<�Zx���D�LW���-���D�ǾXhl.%�F�d�9�	&�;1W:k}:�NA��������H�D��ӱm�)��h���s����x��x�Dy�G�`�E��y���w���Qa#�X5�@��t�Y�0��eM�3o��M��g:�����<��s�<h�id��Nfc�Ϟ����5%L�c�ʭM�Mw	�Z��[9{�^�l��CR7<&�oO��٧�اx[G�9/1q��X�+�^�w)��cF���buh�XH��D52�қ�M�v��f�Q*,#ɼ��؇jF��C�&��e5���~�Qw�y�}�	�bY'HĲ"R������9�<����H02TI� ;d1�{2������v�6Ӱ�0��$��7=?D�Iؼ'Et�d������^|��T:=^�?t���u�����v�pω����6!0C��dq��i'b�t�Kd���c��%4!f������|�>r�AaA��smLpm����t�T�4���i1��c)�x	��=fuvT�%��͛�VPT����r��c�[ԃ�.�����V@�Ѻ�����o�/�FEq�+�9��\\����2��K��P���Z��}�phof�#l񫰩L��zo=/�U9v���u�9�7u�iwd�A�N0�B�y7z�(?�}ӡq�,k�1�m�υ����l,�GA���Bg�T��yZ�8�������Adc�9�`��V�wgG [%@1�q���ױL�#�l����D;'�C��s�0%��[��g�!���]U\�۾���kʍ/̱6�=�5R͕�wf���r�@?���,e�*���4�aa]�������i~Z�V�S����w�����X�z'�x*a�U%	q.Iʯx,��sM�9B�}Rc�������㴓��İ�- ��E�c��^���tds͸�v�7%kbBbb���S�Y�e��+��v&�w�c�������e�/X��r�Us���x�9�oi���i���_�Y�����iH=���zbC�S�Q�P9D�'
K�|J��!r�����9�xU�N���_��["�꫟W^�c(���`\�V\��wn�����x���3���8ʲ���zw�`��$�!��tĿ2I�JtL�sv��uf���@�mG����a�(�L�k��|jʋ�6��P,�=n�U$�ic�3��a]h�T��^9 u�W�r����Õ��`e�uF�v�<b�"��;�n�4���:L5ǌ@���{����7�;�.����8X��U}��Ƣ4]����^.��-�qSG�v>V[���{�ҕӯU���.sq=�{c��sv��S;��9���A�Bf�(��DD�d/�W����� ��LRu�ȔeRa����'��]��u�-L��{H��h�oF��k������v�#�KsS�&Iؼ']���j��5�WJ%Z̝��71���0@R�h]ހ��D:AĈrNܻpis�}�J�,`&+���Ⱦ�ͣG��ŬM�,�ϰzz��2vj 8���>�!?T�#���2��ިhu������ �M���=0s7G0u��6�:��4����=��������8Z��!�77�u�8#އ�դs�/˥e�$�4XU��-@�I�(,J;P�S� *�G�|*�?��H**���{S���cD�ʊO�eW�u��%����]<�UN���o�^��1�z6��͹ܳ�������'M�:�r���"�J�`�{�s�PK�)~`��Z��F����fg��E.�f�B�0>�3���i�R̶�h�q�����z]��1F���o�f�.iu��b��^����9�3�2%�8��T�Kl��F���r��|+�||MJ�]�=fc�[9b�l8g&}ֳ����Շ#(�*a؋n��v�P��M�-o_n�ᡳ<N��:�ӴC����޲N9۶N7"�CۛWݞ"����ث
&{bGnt����{.�-̔�T�$���7F^��Bԩ�6�A��֍�A:�[x�o.� ��Ϣ{O���u����빋�+c��؞��M��@���^a�>0���di��0�g�A�ۉ�!�^(�F�,�4�	�k��p{l�6&���}��fK�O��@ڎ�U���v�<�K��77�x��@���n���,Ƃ�T7��4���M]1p�)�od���[++V������w5�2��b��u^�A�Z��*:����nM�Ϟ�,X���'e�t9@�3ǈ�����b����$�2V'j[�����LȋF�'���2��e��;3�fgm���z�oMl�h(��'_*`$;'�6v)��%1p���x�a*/��/!���./y�l*���S��5����[@N�|��B~�pA���׫"�6]��ʮ���l�'X�%�u�7E2��&���40̩O~�~y3L�s�Wq�he/�aft��Ύ��N��&�)C�<�L7��.���ҿo��/��J&��B�;�zK*os�f�����42�[hL�Gb�F�҇@⮗�E��%�yt�~j	Ļϯ���AΜ�L��'���_\\�wb��L�͗Z�ꥵ�� [%��5�G�e�5���{/n�P��l1A^	hc�i�V�}ƺ�
�����h��0f�F��=z]Ke�t�.�64���l{o�ޤ�Tq�Ҭ;/^�.�QJ�X�.Nc��^�Ǵq[���	γg���{��w�#��4��eCj=4�g�N�-@�w�Uz����:�R/�[s����oD�gm��{��WR�SӇ�c`8!���?�8s��1-�:KS#m���{6�YH�)4lc�\��\g5�~N^O�Ӈ�Q��`K���"(Pj����}�uH�?��hù�Ӧ�e���w���ғ~�~k�+C���N�c��LXgc&3����y�<��y�gka�ͣ`�u�1���;��,�f3��E����׉���lZ��;�;�PB!����Ҟ˄�9��H��/D�u/z�h1��X�۹���J���}u�ڳ�D{c�9��������r�t4Bii��ZD=�'���g;�kn�h�}%��t�r��˱W���uk+i��Nr+&�����N.$ a4���s3�|�7A�jJ�������귱l�ڌ�ν$��|�Sm��G�s�3������X��&._��H�;�a}Ūw�)���GGvn�PG��%65Z3I�ʌ�
���[ռ�|w��W�M0Ɉ�߳����On������*�,�ܗб�8|�?rL�A����ۥ5��Af�JJ�7B�[;�R��P�s8\�=|�E4֋�%��$y��8e�"���`��I�{��yi���Ǐ9,n��W���3�Y�/$ȇ�-=��78TiUYO^�Kn1FG���4�6�4����W{:!�	����I�1,��*Mw��ơ�l��Sۼ �����;���b��3�C�Z�L���C;$��}�N��s�Z�ʒT���3������g��iPz�Zq���8�f��)K5C��d�#�L8�wQ��6�zC�J�-��p��󵛮*��E��^מ7>����G�:�O��i�q�%��ޘi�M��zO�5f�Yuw3b-���.���D���!ý�&C��c��F���ƚ(~�+g8:����y��q�!��������2)z�Q��c=s�2BՀ��Zk��������"��'$e>���.<���V�=����!��(ɬk�2���`��
��j��+b�b��8K�_p���*���^g�����x��K�u��i�i<&��k-rz=;��sI~���:�;t����r��UEN�ݽgHE��æ��6���v��v�pm9�a\Z��sQ~�K�,�s������;��E� ����&��8���k%�!���D�ba�X���n����w.ά�e�Ye�-۵���x��#�q������z�[�����ۮ��>�yY݌v�R�pK�ҮŜ���ι�qy�SNɛ�Dm�Ҟ�+�\R�T�v=�w��mb$_��]�&��zF[����ܷ��f�Uݷ1��U��A^nX��t?��j��:��f�OT5��#`S�3v{��hG��N��(N[0JLJަ�˝®������P��ӏ��U�#h�v��O=�3�m����(
ȣ��C�vN��˷/x�zX�Ukz���;�*�"
��Q�{&��6ĳ�R��n��~�,���.=�n����\��u��ۖy����})�\�{yE
w-��ÓB:�=!�N��4uDL�yՒ�FE���R���sZ�@s����[�Å�e���љ/5�JcT�\#wV�!�@+5��\+�Ͼ(n=�b�f�(T��h�T�*����
Ωʺ��w��w�Rn�ZW��X��#W)u\�����A罚+	�>%E�RJ�| K/��&RN����G7��o��qMNλ��	��)Y<�H�,�v1	F�x4�u��c�Yl��W&F�v���z�H��f�b�N�87�Y`��˩5�0�v�B�u�tb�Ȋ�X[Fg.r���!���Kw��]���t�=�eBJ!w%���T�@4;5�^iu���̮�V�{�%��Z:�b��X��׊L�+�Hu�5����S��j��p���T�9x�m;ۗ���;];vu��{�����R�l�f���0�W�+�?*�x��-_F�I�͢Ћ��K�wg���l��{Gs+\�u�O뺽�U	�jd�jܗ�&��p΀��p����;r���
�d��X�17�?ҍ�k^�ً�1Xn�gwt�n0�.�	���7���W�ˮ��r��qu|S��Z'�om���3yӒ6y�k�@g:��)�=הw-�\X��2����w�#RZf)��Y�L��ٔ4b�j��ͭ�JS;%!�sP�S�����m�����*���v�!�LJ۩y��zX��Qfgi<���%�ּw4��CY�#"�R`�;!�R�y�gv�vF���L=Bҁ_-U%E���W��gmv�����L*�z�T��ڛ�H��A�ҕ�|���i�gM�z��Z|�R#�;6$q�1K�ܚ�!�*��"������˖��쩭^:Y�(�"�*�gBe�^�}|PT��V4�6C��>�)��.�lڼ�4<�	����2�9;�oK��͓�+̌�k�֖���h�'M�쮚͡�i��CL�kT�@��y�'@��PTb�ֶ���S�"m(�ԙ��*d�iM%4�,;��<D]��v]����u�ݓu�MƎh�ج�a5��s��u�~��y��*���be`X�#0ׯ:�˳�^����"֜��v�R��k�����v`WZEcg�Dj�N���.M�z�����/��Ȁ�V�W����j��Y�(��ZJ�&��EY�V�&����
�m��it颣AX-j(��U�جc66�Qz�Sƚ�""��Ѧ"��EU.Ս&*KY�hm�lbj���(�b�`���:
�N��b�h1,Z�E%�RLD�LAESQSU��DP��"��[F�EIDTQM$Qb�b5�mӉ�ݎ�SLU�l�ئ��WC��뎚J"Z&:����٤���"4j ��j�b* �������0N�IN�q6�Sj�X4�klӱ�X�3KLQU3V�24�T�ME����������#XMh��A���m�*��
(�%�j��
���%-Ԗ�T��!lV��A0U51���jh֊�����+A�э�Ѷ��[Ql(*��*
ukh�5gQDZv�ѩ������""����TE�O��Ƕ��7N��0�L�:!2��h �N���_�V�ۺ�;鵝{r����oepK�����/��W1t��vX~]{�ǗW�I~Ultλ�%pLЋw8���a*�Q��
�W�{w���f�}��x��m�O��l��������ޗ���۰��PM�}�P����=�Ă�w��M��-���&u��NxwO�2�3@+���{��A���u� ��hj�0�o�i�����}	�!���|���f���>3�rK���0�T�����	�a��Ÿ���3��3gV@�t��&hh���L�&�P�s���׼����S�,����br*�S��3��a��YQF���u�5��sB�3v���\��n�{u�:�DN�5�.�5N�g�\���2ǿ�^#B�ʤuŵj�b!I�Q7��-oSg`a��g�"z�,�^	;Hܗn;%75�L�ߜħV��i�	�m��;"f�v�r�V��q��ld[B��o@�ca�&�[p����!�wR���h�E5hO�%�θ��]�1�E�q&��A�/A�-ᄍ���0�'���C���ʃz;o��r�i"�jL��W�K.ڛ>Qy�3l���Ҵ���zk���3�Ϝ=� �k�9�괾0�gE��%ۼZ+�p�?!��(�m&@�yc�	=%ܑچ	�ݚ��!��8|m�o��5 �)u�g��ؾ�
�-n&�d�}S�����������ݝ݊s�%n^#��D��]��6��Z��3�� )����̟���x6�;��Z�U�E^�Y�b%��3�(����M�ቒt5���&�6͉ʲX�)�������X��7��60���h��cҨ�����k���~K���k��M�u�]>��:2'�B�Y1�*6��;�Rw�x ��,�i����ͺ;MW���Y~��~J	{kTs$O���Uo�Eu�Ŧ�Ύ����� �t�gG��k�\��Cj���Ú�u*�����2��&=s�v�>�KO=0w�<�w�����g2dK���	���~ӗ�O�7q���"n��tw^��Iw"�y㝗f:�L˴��-��l��I&���"���;�[�E���ʾ}�-� ���Ȳ�]�	E@A�v�tE�����5���	����!33�k��H���\>d�/V��v1�fK ��/���
�r3��\m�j鋇Itt�J��5Xk_g�g�`��ht\L]�cߪ����K[iP?a�7ίP�i�r�--�T�Ê~e����{�������1P꽱L�-�c�i�8�v�S���;R�����d�L�4]�B׼��;�O��Si�)�[c<9�S�͚�ɶv�b�0���!�>!�݊y����P�^����Z�f�:e�af�FMn^NV��P���U�I,��Su�m�6"�")�8�*Մ{[TdY�FD��i)�u�5Q�)=��	gYG"`�͌�B�~;�kT�uq�_Y����l�&��{��c�pߒrw�h㻷����c��&�ZRX&t���������Cj�N�|�0N��Eő�$@����Q������
�W�#2��c�:�˂J�
�|��a=k�G�fΗ떸Hjٽr�SlX�mԺN4Y�JGcz(�ahԢ�tSZj���y�6�Nއ��IN������Y�
vmg���	���vl�%�vۮ���i��(,k�t�~h��fg�i��ynmV�ư#aЫ��!�y@`鵧��5����tf-�c�$Q%Q��Q��g��n1�ؾIv�]�[�4[��4�	p}S_�b[V�Qke~R�Y�V��-̴u�'���F�{�r{��Q�&�Y��?��St F�	��n��LB2_�K�=��{n�!v��j�()U�l'������;;��K�gb\3o�D"��D���3j��0��+�S1#�f��mC*�+��{$����\��� LP��lZ��!��ûZ���g�_���sz4�p{.Z|��f�,�&����t���=.��)���?�&_P�Fi��BfnD�!vT�
�(4��]��$r�e�1��wW�i�Z*�.�Y��꘲��&��K�o�{���v���1�V�S�������˔�Y��ScNh[S�iL3)B0��-7���E����I��ַ&8WgS���z�}�V���%_�Nj'�1���2H��I�/�wW�2�3Gt��w��(�|������®�o&֊xk��!4���y���sb�}<�/fm�jJ��Z卶(���I�W!�+�p�N�	��:kz|gb};�Ëhq%����)����Y�����vq���_j�;�Se�eMV�SׁFq��|�o�[�?�P.lD��ҙ���j������= ЌU���'	�K2Oa#4��)B�(�|j�t�)�ݣ��"6�;L\��]\��	ٕ	��H���öv.�K�1)ե"�U��66A����A1Z5s�U�"t�>wK�8g����Ǡs�[T#,����˰[���Q�$��b���)u]�ZB�;�d�@��v-a��f3�����l!�^r!6��m��^��O� ���:��ŬL�^i�»`�V�*/���->:^F�=4�{�?K�'ְ!���8;�lǐ2��7�Ƭ�ߖ��~���^Xސ�Cג��X�;�c�;��e�~�M����Ue[nuf��"0>��*��zJ�}ڷy��'fbv|���lJ�e-]��7�Kh�I����R�mi�}��H��c���@�[՚A��Guf�;yk��v����S��u��,j��m��#u�kE��P��6)Q��2��n!���Z���d��4:�1���^��`f���Ư(]�L��������_�5"�+�Uc]���Ⅾ�M���k��wf�vCk
�Ú�a��hʝ�1:G���ν �m�BՅ�ux�k-rz=<η6�l�v؋�5v��TU,�kv8j`�pp�b�C�%�j���4:�vR��Xo���LQ�s�o�\�E�������<�_�{��3���0![�L��A���K�;F�2�ۑk9c���L��Ts��E���dw�CG�\sO�L$�6k�m�΁}/�w���ޛզZrc1ۻ}���(�P*B "fK�Zz�x4�Pv��`L����w�zS�-�e�^�n�~��^�mz��CsU�A#!�׳l��[:y�x�`P-#��be�\Cv�j�D��ݳXDG�g�q
��j�>�A9�����bP�{"��*z��r��B�g��|���gl	��<�a�]��&��\���X�0�P�hR�TXS)Ӎf�7
֚�ν�6�3�t-������0���nH�=�����2/~s�o���V�ޥ���-;��BLK����*Oo�:��5��JO�6�u��ʎ��ޏ�s�H;�;�9���ܹ\ ۹�o7z����EAΩ���7��*��X�bC/����f��R�8X��[�ssd�uz�:X�Ux�H[�ܡ�kGբid܈���}m7����NF�l�Ǧ�Μo@����;���.��v:{�o_��N흤%';���<��)��C�_=;ݼ0�qa#D:O��G=A�Y;T�u��:�G%ڹ��Jꆓ�)=�Ⱥ��	�-/#kǦq�D�ҍ?P��[g����݆��\Ƕ���T2s!so02��/�ݞ'�R�v�aTrW<�ʄ�'��T0����ɟ:�n9G�I��o>L<ѱ��	�=mE'&nA�vN���,(Z�us*��������QS���6�`��5���Z�З�����t�t��@�4-XQ+W��\��^ٳ�gZn�-�d���xQMH���/ѝ;2�Ё?u�	�x��g��&�W�(�-@�T	Y=�ތn#ٻX�ʝci�vϻ������q����}�!�������C�����{һc<�)w����HMB���w�F��/ ba���̉:"�׺����.�����Ƅ^�Rg��O�N@���k͟�`X�[�/�Ȕ9@!��L�I��5���2�O��O^W��~9�7�(��=�6f��Pe�8{q��M�ڰ�̽����}W��iS1A����w;��D����f��L�[N�~h���̏�H�]�w(rnu�t�7�!������-�mk����+�O��<��rN�/�1G�]my�|��ƥF,�C�P��\����5�q�������Ϳ.�oxI���=��h�aA�q1w4^�Uz��K[V�!k߰��T�U:׳F��<W���Po�ȟ�`mM����g��ڽ`�i��ӊq��'jXH�!5�n��v-�]��}��^G ia��&����馴����lH�j�eb'ץMޜ|1���7{q�j!.��^�&�'�t��}��e~�g�fs�й��㑕"�W-ֳ[�W7��úRV�TɐI=�`A�!��O�����USz0ɧ�������=lJ�u�����iww[}�C��E%�b�i�t#<�����v2����l�w��O�6�;��K��&����)⢻V��?�ȥ��ͰR�09 ?�r�f��VI .�Cf�����i<�2ݽ���o|�v@���Czo@p����@GJ�G���3Sf��51��`�ɠ��g4]�����Wgk��1�@wc{��︚˖���5����40��5n�F^�P���[Т���@�`\A�F���M��t�zF���=wMNA�GZf�6&�[qX�,�<1��i�����c���^e���g7{g��n��"jaX�s��w�v G�F%
�u��J0����HI�csrA���Sｼ~>��04WX�I�����V¿F��=^b\&)�u�mBg������t����߯+�;:Q�f�
g�7����M����ugb��(w<��8��j����ͬ��{mq��Zx�{+'o�Q#��WG��]�{8]�;�H��e?(�R�ϝ_iZ�G�+%7>5hu\<3=�>�v�UlH��'ڰ��Z���)�qZqA�J�8ӗ��Yl�������]�nQjل��q���tG?q��yz	AM(3ǮS���s"�&yR�7Z�d�4��8Z�$va@=��Q��Zz	l�F0�܁��Sc"��+ה:چg��S������=!�����$������V�T'`��}f�z��e`Ծ�<#L�n���1y���̜R��+g*�BV�S�wa�&LY��̮��̓XCi�s�ݥ ��r)O��a��:en���p�������'�/7.Ƅ�x�x����S/(�tVT�ͪ���R(�v�li��0n�&������o��Z{ �]����ͬ���<. �e6����)!��]M��CTFs�Qm�_E,M�Z��S��n�x]�Ab؎����|��󱻭[b&�{L�����P�I+�.M�~����Q���W�S���"D��U�g!�vs��V9�ɻ{ʐ{�z��ϸ2Ƃ�-�̀.�8f�T�y�O�h����m�x72v�2�PUxw%4�ۦhҀj�N�3�Sdjdr [l��uZw7xPāp��}��#p�.St����Ho(u��]ِX�����o]vu�u�oW�=>�ZM��.��d�=�%_��џrn�v)�n'7q�����"��}�@�g��ge]^��p�x��]�A8a�[Q=��M���zǽ�E�c�^z�$_C�R6*Ѻ��f2��I:�+�$;��8H�
"<{�=�msӝ�<ޏ?�˽^GQST�0��|�m��{R�����/���������:1Q5��mݝ��Q"w��2PIbB�
a��ɶ�ؒmC������g���7���[�v0.�L��ҷs����b-� zxh���"�,���y�G��cr�Ǧܗ�d�Z(~��4�d�F���ٌ�}��<�ï�!!.��j�S����������[��ϣ�"��Uzf�oڊ���QGOV��Ǧ�a��9ݽ��ׯǓ8!\X�w�m�b��+�J3�=<�Z��vJ�zx���{x���M�tG�s�HF�k}���������g
��ᦒy���'��>��G'��LzE�S�Ϣ�B����PrF�W���u�w#I�䒰�*R%�!��Z���:g:E�q�C��F�::{j�?���7^�O�R�Ҹ�jKK���o��^U����q�5�����pcƽ89Ov�jz�ؕPD����wI��T0�`ѐ�`ڧį$�K�]��Ǽ����Vq �eP�\�Z�QAV�;v^�
^U�s}]PfXRa ��>aǤd߻U�k}����q�,����w\9p�-e�Y���^�W������|�y�g�ckk�a�%J�B�.ط֟C/�>g��wj�����ֹ����X�5��;K����J��[JX�r����`[���IǙ�t�Bi0��7B3�Ꮶj����lw���5s��&���`��3qu<�+#A����}%C[�%c���8�\M��f�k-wt�l�@fmw����XQk���#6��<��[�ɬ��!�D��8�mK�G�ٮW*���V��]&c	W�;��J��Y�ʄs��X�A��\����vA��MH'�b�UXw�,;ws�;�1!��u|�����汴pe��#�]a��u����n�r$����CU�͛4�9c2�vSE�!&�4�Y��y�iҶ�uIQ�����b	��kgQ��Zw����o^n�~6G+�v��ݷ*�	��<Ҋ�ĝp��,���f�{�ok�u�1Lu���lӞ�������Q,�%A�7�m�3�q"�+�VBL��P��8+�}���'�]�]Z�n؁�=�"�K���(,s&Q8w^��95��c\��1�j<�����h����ӺZX�6vON��l	�˱l�!�`!�Ve����ua�V�R;9.��)n��R�l���ԯl^t���t��w���A��8u�Ns�[��S("w$I��%ovT.6�ZSm�נ�,;�ć�#���';�kxa٬Ȯ�NW"�)��S�wvt�<��R�6#��w����;b��u�� Y�1�<IQ���}�g-.�����(R�H�I��H�+۬��ҀU�,-��Wq��_}v��ٖ������&��:�W&*�N0�Td�&:8ා�Y�ܯ$�=�mA���n��2�Qx�tU�[w�[�D�FOv)�Z3�[���漹d��,C�x�6�͂��Uk��aћb����5��U#�hߡ�:�t!�2.vm�8kH�vޞVh��q���ɖ8&��	�X{�Wo����  ���t�Ot�3�u��Zoq��W�|��M���6�a��\��L,.%u��� )���ٲ"�Km�p�5Nv��2^ӣ3��)�R��Ս�e�C4Fr۶]p��ۏ�Ѿ�"�)Igg]#vc���Rk/��^��ͬ�*�-ۺ����
����h��#srY:C�5y��O4p2ZB��eE"*,�D�����+k,�����'���=�݃M��1C�d��(0�uc�9/{h�WH������Rq�Y���p�\�wk#3^�[-�**v���[3��dX�YY[���wnL2uK�Nɑ��Mý��E�{@�����7�h�P��q�WD�T2�JBa}-�c:�6�0u���͛���A�v(/&���b����+2�q��VY�s�%ev�.u�`����[�������Q�ٹ������t���W�9.s�n)�:���S�W򪒔�vk���� ��,
�#�qBk�m�f��lB��u����s��]D��<@�Vz��<��U%����(�����a��j
6hƌUD�8���L5�����gL�R54QTCx�8(�6�MAEhT��SQ~c�sU�E���F�4������)��"��"Jj�(����(���h���H�tm��_���4AkPC�U���h5m��%@V��U��D�U�c7A��kY���Uh�U-�C[b"�t�#�%�0STEE�UQ�����E�LKAm�z�A]klSCT[b
)bZ(;u�MSATR�4PF,�STĵ����Rk-4UD�h�ZI�b"���q-5TDUUI�18&��
6�[f�Z�)��"�;b+Na�CI�cd4[:�?���* ����`�IT��d�btj�td?�0=i�9���?f�16��>h�'z�_]ۡk�S���u���#dv2�y��u������"��[�X�.��ٽ�{��y��9)��}���+��5��x'��mm�o�T�����ݢ�myɜ����#�`@�c0�Y���<y�5P9Fe�Fs�����{��s.��"�t{l�L�>$%�݂�tۙ�g���t�N5=6L�Ry�2�ŕ@��6�������tW܆R���s�{�i��~5Xz��ɖ�!�T���jF�������p���$��PU>i��[��}Y����C
�=ܚ�����ԥg{
���h�7ڝ5F�V�ri�w�[4����8fq�]1g�ޓ9F'�)��j�x��H�
�6��Fc�� e����յ��ɹrC��ut�3k�ͧ�H����J� ��#@�P��S���2���ֲ�.�!]����m�o[�"	�:؈|��I�w�ɟI�8d6S������<��m�}};�����3/���K&f�;)�%��9��rdN�C�[t7��A�r�m�I��=vD�����L�[æ
����{�W`|ɤn�ͮU����f�g�m��к�;�Or�mf���X���E�aС�2��ٺOd��P��l�����j4�ޕ�Zx�Z���aǞ����V��,�!� ��V���4q9��Cy�ؖ�`��O�3�Z�7 oה2���}�>��C�aP5]�Q�6��̨8"�ײ{��o�R�"�.�>꿻���WI�����y�޽�Ե����@�`��ٗ�z�����6��L˺f
�r2���q�W-�ӳpϋj�u���K�!r�(��χ(o)�%� ��
�pm���ΰ���N�Q��3G�83|$�c�>���y���l2ܣ�/��d@�(Ԭa7��W��v/l1�:����A(��%��t\�	�wF��2rk{��KZ��#=`�K�S>�]�䕃7���.臗�̅t�L��]��*�^:��7���yM�h7���'j�h	���?��[�N��\�TH�U��M�q>'�+['Yj�mEMJ�Y���d��Du��R�N��ui�^i-�W��v�qv�:��rb�����W�4�`�I��m�7��o'��s{����d�QB���yYK�I��E����T��F�Nc5���2k0�s�nrѴXމ
E�*rT��Ē&���i$���.�dށ��(����ne�v&U�R����t�E�N����@�֨���s@��{�ۨ��YOp��N���x<!���Rd=�BQ0��FUB3 ��|'�a�ͭ�8wwM6r���� �~��nظjG|��%R�*p�.tc\F�F��vda�n���@"�ΐ��)���ۜ��{�H�DΆo�ϩ����·s�.��e�m+��6=��V�>��4��`-�z�*v{o��A��Yl���sw�BX��i�3Y���lP����JO�ͼE�לqV����m����0q��C7_;zm�K�v�|����L�r�4:U��rSKt�x�5#/i���)�ӾKnY�7�e�ĈP,#S���4�+�j�'��vk����m��F2�/N���ѫtk6��j�P��*�c���\�qIʺѦ�XөV�X�Gc ���V�5]�a9���n�c�s��,�j���*.ЫWg	��1������(������QK�{�>W{ׄ#�5�N�t��)����:�2����y[���>�|狷�z�6}��:�����|��;�8�P�W�01L��w�ަKO#sL����e�h����꺮y%c�r�x[P��V6�kx���7��L?wtC:�G���5�׽�,k2fdf��K��땑|p��!���H(��=���yY�z�h�]�����᭣*��5V���]��3WU�ˋE� ���'�e�oiO�[�v�M���J|���ƹ�H�������/U*"�ldT�K*��4T�����~^!�<�Z���T���v7�#ö�W�;��V����*�=p�&s�Ϲ�ix�-��m<g�W/fs&��м�������
�-��k�!����յH6�O�y0���$�>Z�n[�́I!FZ����Q��?*1}��
��rN���V�JD�mh�sc��o��%u��U~6�a%�0&�?��ԼeS�|��b�P��*��c�c/�e5I!���tss3!��͟g���Ùy�w��4 ��[��K��7�4>ۑ�S�ʶ�[�dx��ͳ�5nN�>#z�g; \Ή�ӗۥ!�j��T&�X[��tr$����V��
��w��/���[R�\��Y�99Y��^���by�!��\����Ξ�����.�� rҠ-wH:]9��&�E�{G�*�;�kz���%���,:��ْ�Q7�<;�HMk�A�s-��=Hu�+��M������ᅺ�c6�(
��2�2�չƕyB�c��q�Q9�zZhÁ?<��g�m�3�mr�1�Bx$l�o����*��}-SQ�0��Ǩ���~���2{�{������l�s#�ԣ�o���G��h���H9�ܨ$��xv
�m�;q�S�&OT�Ի2�R|S�!���=�һ@�̶���<�Ĵ���j�Ӆ�%�F��{G��K�7�k>�b���������i�* 闛c��K�g���r:�;m4�yu��(.����^����#+O���]S!5Q����D���ol�op�2�W�Ϩ��c��0��oy]	|cmX�Z��u�׉g%'3�n�m1�l;�8����&# ֺ�#sq�'`��k�:�6��ž�XWF���_	,��jCy�\-Z7]�"�����h���Sb�3�dou��,��3���n~1bOS��53�EU�t.��#�vh7@�J��)Ѭn�TӚ���Y7��!���qL���M�[h�\�.����^V4�%:�w���HgX�P�2�(����2Ms�T��S	@�b6��t���������wo�K�)�&�o��i5�\���h�+��]l���{vy+�*�u��x!�L�fH���<׈����2m�S��,��w:M��[�Z�m����ݝ4z���OZTR���uhj�}ƥ�X7}��^�x^+��d�j�V��<{���������_v�] ���n�t�á��'Z��d^H���*��a�TU/Q�*��~���2�����e'��1�I�$�z}��-]�p`�\=�<mgt�''�o)��I�:Cl��ޏ*���oӄ�=�)�.���[g2�՗�m恙��J� ���%�}�ۥ��魨.3�q`Aj���C����*�*�;��;r��lÎ��85��039�(I��\՝�3SjQ�:+k5�N�9�w�f^��4������YTj,z��i������u����O�Q �{����h�+�s�t�Z�n�<gd�f��kfܺ:�zz�i���c4
�����Y��	 ���o�{j'�Tj���M7/.�<���De��W���j8E+��%^鼣}�Huu4��9����{wo�C��Q�hO"��ʟ*6�nY�c�	�U#)�Ce8��]��s{u�p���>[��4�By$�T8�3mH�e-@ڔ�L�e�.w�~����"���C��m��#Q(�҃ǩh=���zq1�fK�(��pc�7�}��4 j�/kW��D�\�W�1�ѧՔp�NNu��R�Ump9�NEH�T�q�v.�R4ܽ)u�c0��!�]ڊ�G	i��մ������������y\���5=�4����RrZ����2O.&΀ُn��-���g��#��V�Mn*	�@Oa4��9���Ʉ��,Up��V(�J'kLX7�q�ɭ�d�5Q�3S�������͉��B�	��)�9��V̶��{��	�,n�р�E��+h�
����Ճ#c6���*M*�X�v�̶BS������\\!�֤d����OWc�_�Mx��@1�9���S����fE��kT�M��oXt�B�2eW���������ca9mr�u�n:�/c���Ƃ�hOs����~�ή9��)��b�i@5C�R�xd��2/i�o5o]v^��5G��%.
��vP�4��5u���=�G��V����t��vvld���e�����#u*��;�wx�����eYs����^6�~N�ú:|v̎�����M���Мu[^�% 9�0�<��Fn��m�������tr�o���E�8�~/���g�
��s�mZ���[G>'��'X�
�l_Ϙ��C㝁V˴=B��|evk����i:Ɉ81~����w���;���#�*�K�ܭ=�z3%���w	�{�˜�R�8c�]U=^6z�dT�Iez��4P����Q��ӵ�1t��&!j9�aS�/��e��n�Ɂ�*ͦ�Ej��;�l[jn��x�
�(t5���)��,f9v��wۯX*���W�M9n�U�#q���%J�\^C��gw^m��S�B�e荰̞��fH�x�=3�L2�J-PSw8�fJx[4�"[s1V&��{�ʹKѬuǬA�~jѡ�|�B��Ϸ0��o����.ש�4���m�~�̗W9y�("����יs� �3����:�A3wݧ͋��0� �R�M���u٘$[����^,^�O�otnv�@W7�~݂M�$��J�����j�3��X�7�іhj��}���i�p ��;���n)'�\�zR��<ch����J�+��H׳�&�d'C��#��P�������*�F'�������RƘ�m��'*Ly���-Ҩa��^`����vO�Mv���r=�X;�';��"c'����l�e�s��������`�ڨgR���4f
t7�^';_������ �o=�hs���:_ ��F}�����b�eGct���Q��Oӕ�2G��dv4��c������ӗ:�\�'��ٖ~���d�P�w1XU?n�}�`��`� s��v�$��ODH����N8q;]��!��`#��w�`X��zu\�;.sy��x��L��0b��5'�&^��V��<��Ky��e;Q����)����ۘOt!��AFXW�?�s��)�����^&H�A�&7ݢ�M9Z۩M���{v�O6����u[~ɼF��;2���|H�� ���U�U�{�ն&v�-�ޮ�����"�8#��ԕ�f���s0��q�[����D͔�q�����j�]d�ʢ~���N�����7N�.6{�R�(-�[Ժ���2PK���SsNge�
z�wLyIg&�2���̓�ά|��9o��i��FѕP��;w"���[62}���
ʞܢ!����9+��s"Zt��C��r
|z�y'IN���#�&<U�D��qG�w�x=���_�A=lF�Ғ�0�yl�����4A\���_�9��͠n_(��#��E�P[.���<��E^�u��ۊ�ő����u*�Ѿֻ�3�B�k��Dp���w:I���tz}>^�/w������y�,��,�nݻv캄f43��/�iEoF,d��Y56�Ae���šń��&v� �_�!�Y���mn5�.�39:R�{]�.d��fK�v����Ȋ읖A�t����v�.�
����ɛ��p�fi�q
u|��F{���9�oCY�cV��	
��̚F�{�j3�:<J���>ვ�S̫��S������f�썗���2�G�:�G	N����:KA춏�g��-�Q�t��1WQ ^I�{U99t��*Ň��)'��Mh���8����r�L�m����ER�Ar;�rGM��<�K��B�=.2	��z���ݒgGr��Xǵ�P컥"-��F�Ħc�f�n�Z{Tv1Z:��↑+N&���Twt`�����M�(k�3t�1#��Ǟ�aZ��h��v�t�9YOcoM������:��:����i�9Y2n�]�=�Ρ�7l��jHJֲ5u��i��՘T�p�ǉݚGF)دE��w]8vt��9�1�{�oNʽ�7�kN>�\V�o�<﵅��K ��1��S�i��e1{y�u0�!D17H����!�zt�t6]B���8�Jf��0�B���M��mƀ�<�oG8�P�MU�]u�+#S���;u�\=T3F�Z5�5c���(��B:�A����=�rv�Ol��j�}Y[��ܒė��v��V��,��0U�K���ַ���l�@�wm^����g]��]�R�;L���̢�j�tu�Bt�P��n�0�r�`�m�FҬ�9��Y�Vi5�Q�e�E�7���P<b�l�.ö��L��J�k�EI��N�c(��1l�#�A��E�{kzǶ쵉��Y��s�Ӄw�ݫ�œƣh�n���U��;�6��`�cU�[�*v��,�*��sm'p)˖̻��u���x\�f�k	t�o����W��ɼC[3!�bh�޴�.GN#N\+���,|z�]Ll��t�n�f6r���1��Z7(1�7��L�ŖN^�9���A�r�`U����� Wd�ܝ�s;#(�{O���w�!�;��N˰Ctr��O8Հo�9�K}3�4�E�_*i��:�_k��d�B�EIE�'��.��/��V��.K��}ϴf�J3�f��m36 a�u�k�u�էx.�7�d��G�%˺{�f���zQ.�R�-m���i�I���nvU~BI,,aES�	!qU!�&I���d1W�`a:5�.Nc#\����,�*iA�K���f/:�MK)o4m���'V�;oH��9�'2���Wm!"5��Z����  �̙�x��eT�8����]�ax;)Q\f��������V��v]X��Gq�0��|�oi��R1�lvN�����/�����!�*��Xk;�Xy��.�O��������-�78[�sQ�ɖb`բ��:p�Λ�n�U|� ��v�3++2��u�}��%��$����c�ْ�4(�	�r�9t�P����Z�ӻ�Ɔ�/���A�٪R��M����j��bB �A�e�jJ��"�*���(��t�h1��it��()(�Z�(��F��PkZ�CEST:�˪
(�)JF���N6�PSER��Ʀ��Ƶ�*���R�Y��ER4ձ�
4�uL�4Pv0�ACE&�hֱ�Ek1�K�U���t�Rm	��_F�t�ݕ�zB�4����ꈢ�Ӷ�ض

I�"!4b ��ED�\D@�d1R��1QATU���*���i��5�b���=���h���MP�6ޏ�`�c�X�EQ5v�$�Iۡ�A��sUEӠ�0Uv7��U�����d�Y6��TT�^���kv�x��g�]�T��:z�*�6�h�'A2QE�Rz1�T��g�?���z}gǺ���P���
dfO�����U�z�v��vD�L������V����C����	�v���R�4�R�+�ȯ6Z��8��^wnD�`�٦�
I��M��>�L4B.�4��Ǎ$AH�n��7��]�y��ha�������jʲ����Q���+����K���喌�V(WuB���>�ٔbB�1$�]��n4�7�0މ�,71P�;���H�F��ӄ��w�w�B
�*0l�ܗP	SR�\]{)>�����9n��i�����gw=>���cdnH�4����a���0|h>��YB�s2��Ffvk������D]�3� ��o]6�B���<.�U�[�dF�S���$���k=�j��E��³Cg�ѽ�\�R͒d���v�z�l�����U������.��*2P�k�vu�8"O?W�����hO"Ւ�lS�,��� !�I~�ˤާ>�1>�)7՞~���s�E	�r�KR8ٴ��L�e�0w������R���^�wn�ڞ[T`D,%)�{iv�����h���ђ:f���Z(϶u��nW���f���]MD��+�]��X<�S��f�j���VZ(K�p*9�5@��ύ��خ+���/v�NR�J5l��s$N�P$�=R�H�Xs����m��=y�I]f�I�=]'i�_H���Q���νR����(.^�;�>m@�&RH�Z�ݜ�1� Li6{��n��T�[?�'�r*D"�q�v.�6�D�TE��uTw.�5��`ᷬ�uR����]:�0�t�y�(M����*zM�hnm�R�8ܝ��|����ei��x�ۀ�9z\?t��iwA��M]ی0�Ge�ʹ��'�h�j�9�@�#��Y�c��n���ۼ��C�Ǡ���b	�Q�;��[i)仧V1f\%ނ�{��8�t�?7�"+!�l@B�U3��M �ʮ���]lvz)k�#�w��+��TZ��z�J�`��`����t�O�"�7Ҽ�B���߳�m�K�xϗ��	`6�B����w,��+W�g��۟��Ÿhvd�\��E&�P���G+&:A�=!��6�i�u]~�^����xXO?8��P�9�p�iV��Wh���>\�:�����������5��c���L˽8��vt���+�I,�&�)ѐ�bn�Ä�m��y������B�\7L�=�ʇ<���\��������\�ݧK���z�K�`�7v��h'F6?V`��>�]N��x��(YjWG	��`��D��c�G�U�(��n]���4��\&'y�Ӻ�fZ#�� � �<r�\��/���;k�k���p�C�F��U	���f\|����AT��.	���Fi���{K;��ׅv{gʣ���=T�L���R5%��������;p����ns�dܒ:�5�\�p�� �p�jϒ���$�!��i�NOX�cܒ/�o����p=��6�&�"G��
�P�3$�sS���k��9痈^����H�9���S�$�eG�nc��"E�0�6k�%��wF�_[rm�p� ���7`�9$��$L���|�ʱLt�rx3�{!,�94F���L��c��Y���u�XzWmp���gq���r�h�z���I;�Zo���C	r�r:��3݉O qtH7K<���]�j#���'|B��G	�	<!J&�W&�n���W����qˮڻ�}�D����O��N�Z�7S��dZ�nK�%'�6�e(�k&m9G%�Į������z�ġ��)��d�t�`w�`�gzv
v�2%hk�	6��)���]
�h�[�����g�@F�����'�+���|}���w�SZ�'&��B|t�3����{��Q^T}�^�ކ���̀�_��]#'�J9J�ϰ@5e���ԟ��a�價����r�����/� �x������/��r�����q�A�H�D����=Ѳ;�.�^������I9i�Nt8��]��!t����x׉�	��g��^6��h�&�sL�j��vX1вΨ�U�͇D�PI�a��b���ΏC'w��cs;i�਷�ٴ΂���{W8��ñ5�.4>�6�PQZ��V ���\/Zή�ݛ��^ڞ�x��?�wB	5�_�}�M��<�r�)A]u��=}K[)/�!�P�jR�k�X.i��e�
qA��i��[f��Cͮ�&_q?d�Q��!_rH�є��ʭ��\�i�����e�Hȁ>�y������;ؼ�R�k$�*=�b�Ε�*�|>Mgv��f�M^�pc���|�|�	;�w�y���(CҤW�h����7oWs,jk/o!��C/mY�CZ�x�Ϧ���%����1��A��$ލ9��-�y���-<�mo@{��7��M)��DX����[3""`^xg��Hh^<�"�B4O%B�N�w�P]y�b�v�i=��3�14=���������>g�]�0�-�tt�7���nd�7�ِ������ϵ�
bV�G[(�Yxvy*vX���V���u'���u��Wn��C��&��z@߶����R�������U�W
5Y����kC�㖮��괉���B3��`0����bv�a��Ǌ��R�|���F�PD��1$�ɵ�0}�p��^gmMskR���Å$��J�I�{��׻��H��
�æE��O��Sυ��.~���.�pb�s�#��J/;W�������gu<n�f�֒U��a�_jb{S?�L�#�̌��}�[dvO��/�.��eFv�L������������h#�=�xVk�8�n� �!91�o��mk�Y���Y��x#���4\<B�׳���� ���.Al3����U9y�]_b�\!��>v>4��Q�����x�%P�_�m�cp���u#������v6^�=0J!j��nj�N���/Q��8��b�j�]Y"wYՉ�I&~^���}���423��Y.�3�t+���#�ƫn#�ޫ����l�ڋ�s������V���h��b��K8��̜�E�z���V�4U";Y�0�a�(���c$K���	2���6nx�G�e�N=��go�-Ͷ����yG�.�=��+F��'Q	Ap��R3����ٵ>�ռ��i��w;/%����D.�5,�@���N鬊u
�[������}\�Ú��w��=y�"�?�������[�v.\���rٳ�Ou7��	�Ѽ�Kt^:�$���Ǻ���\:A�(b`S5��w��wOC�2( �J���X�4d�'�Q8g͘�6��!l5$3z�g9/�1�tnu��������k�*���n� �Vs��7�S��dE�^�f����N���tU�~�������֒�K�}�����T�'UsE·�.杤L�[91n���m�6�^��Kwq�7���\�+?BbL�E��<�_W
�4*�Y{ϐY�.Ua���S�U���:a^V��0�i+���ј��� 6Z���m^���ح9ʊjMl�6�T����^-��`xW��{A�<��\d�߫�Ѡ`�W����cXA�n�#fR[}������8�l)���7��3����j�cW�a���V}�^�M4�^̎�
��U���ט>��.k�s�!kl�j��p'h�H.Pq��>��_��������a�c�ӣ��$�e�z���bŻh�v�����rt줕��t�d�p��Ē���#���EqQ*�i-��N����r���C�ĉ(�=������]!yY��Z+؍+R����ហ�5uY�h��|A*P�z%�6١�'KE�]����b���{�=?`^�9S�͞�ȭI/f�U����y���j��^��$�)�����%�0�����+��1{��+O��l|��);Z�U7[�!�<i�}�履�d��ٵ���=\7�ߊ��9>����-�Z���8{�Ҳ��(}�0��>��>Q2!,lƙT�8S8�s�fB�y9��8�uF�C����Uw���ǚ��-����uژ'py�(=1u�|tmc#/[N���v����u(�)kE"VT�����w�K��6�H�9&fu�G�n��������;�u����F��U��R<��:����\G�K�nF_�0���%���B� �[p��v
6�J��*|�2kv�C"Zz++�NVv��|�G�p���#clʡ�^<:�=+�Ԕ����݄�b�����D�ڣ���pG$?���fz�ؕP����2�kMg��ry����ӷ��]>��P$"�� 0�{�!q��~��8{�ap�|b*�r�;w��������~�ؕ��A�	;G�@S��]l��{�;i�)�k�хrj�'�����6���oЃ�����Q;�E��V�`��0�YF�u#I���ݴ�P�8o���Ť43�l�xG��V֑�����xW�2G)�k�$H���vL�Z�*�׸<姏}��6���q��:��ȫG��:3-�n�����s�0;�ȳ���1�	5���桘o�k�o{���xfJ�Lf���q{����s5��kv�gxP��7��m��,��I%��콊��'��i	wibs'p��n�S���r���J��d'�teQ�cMUј�v���ix^P�b)kW�u�����Z0L�N@
��D׵�ԁ|�11���X
�q�E�/}��ZE�K�i-x����O4�k�X:)��}C�<�Q绒G��]���H�,�ޓé� ��Yv��𠦕)	u��G�W����e�����g�����p�p��R����|{�+�Q�5�@[w54���ز�m����Ȃ:��ӊ.��j�'݋��y�'QP��P�U�YY��S�{WF���Tp��@(8�#�o��t����$�5sʵ�7�n�����9�ɺ���k��q�EtG�X;G�˭�w����V�Q�g:S���|䇉����T����},[a�8A{���j���u�ۉ��^��֟*��a<Jh�T�m��{�wI��$���a],]�����!�t�d�6��7v�fүa��.�-D��mv�a����vi���c�VMM��=us�lJfR���������ʅ�sqwu���Y��� ��l�|�:S��!0cy-��.�_)������'fk]�^ڜA����^)��U��. W��?M�\�qlv{v�#5�lL�+06a�cOck.3����9����X�c7����FF����^��=�o$MM}�wCc�������EuUfi'���Mxv����p���}(�����Õ�~��]D:5.�x��H��شP6#�z%��{!oo�Ǎ�Й�9�ۋ��͍���������aҶ��b1K:с�Y��J:{ckQ�ܐr�u����?C�~�]�w��ګ%�5�3���;Lg���q[o?+>���׻�F�@�B@�Ze,�xl����Fq���"aGk��|ˬ��r�T�܋Ԑ��z�M�I,i;Oэg���V��_5��C�q!mu;�":ɠ"�$j!c��I�6�Lk��CBܠ""7�|Qt�%�{o��J��<5 P��z��MkF�U!9��u7ئ������mi�N�`n�U����fBr-�X;�|����W�������e�Ye�v�۷e��ff���n��V��1��T���P����tk-5&76-�tsm��ݟ�@�#���+wN���v��Y�����]�Ku�M�؁Uf���ô��S\gR���階ޥ��v�ݒd�6�^_:F�f'b�8�5	q�%�����,h�2���K[�t � �0�;V����r�{35u�hs���U��35���!��H$��q`��[�`�)ګ�����۫h������ޡ����0<ʽ��p���\/7�=��Ƕ,9��(�ū<��&a��5�R���0���w�ݭ����\w��:�'����ٽ��I\z����L�2�ë��S/���"Bvb����.�(T���]c�R+o0�1Y̽1R[v��Ol� `�9����uw��skA;�n�R�.��	�T�j�Y�.�/%�dܬV�G[��R
���������;�K�Hէ�,�w0n��j�f�.֩��B�]�X�J���XiI��"��g����^L���F�b�)+x�Dj�Ѽ��g���6�lȟ^̔.�:뱈�P��d�ztil��J��*f���q!���ae<b^ۀ��͝ Q��ډ��Q-���YX�T
�CqF��Vf@�^V_2����*-�Ӭ 1�%�Ͳ*�y�M�Umی�o�	�H*���W���Gt�1J�Q�7���D��W �2�kU#�m5���v`捈y:f�;�1���V˖�ͺ#x`u)�{fp�WX��d�ٖ�����j���W�lpqV/m�ԓ�c?k��oy��l��T�V��gZ�YB���mt�
�;�.�@���kCh͋o����qG�Rم	Y�pT�S�h��Ò-ۮV�E�9�xC)n���2A�ܡT���^n��R���5����Z*�g�>���j���N�`��a�{c�-��w��;z�^�� 7z&$4�`��Ս=��_�;��]�7:h8̢m��N��h���b��[��Ɍ[��u��qː�;�(��ۄaױ{T��pd�t2+sG�^]��R�Z��%�rV�v���Oc�∥�6�N��3.M���Krt˵�j����&���N���S0StT&� ���1�V�[ ��d�PÓ�Z<��T3C�V7f��5�ĜN��t���Ҳ���WWHv�N/z�8u��w�KK{U$�v�N��4�:�TS3 �\�i�p1�]r���T�S_l��W�uYS^�e@n�P<m�Ǌ9r���G�u
���J-r�X���d����W���{�)v��y[,�i�Ei�`�j�c;q+
�skt�һ�
��F]�d�0�	80{�,�x��mjg^������r"q�#ɴK�(������Ob�i��T��ڒ���w�eGn�nc;g[����;8��Wf�vl�#`$�)t�
�4*eۣ.��F�m6$^V�F����
$Z#���6ڻtTGGq�X���jb*Jlk��(�bh(�J����j�Y����k�QDDEu�^�=���h�M�PR[�����t��1]�A\Vڊi�$���(�
��4u�h�&�O]%���OZ)լPjb����(-�TTZ��w��{��td�G�E%�q����.�=*����5E%I�ؠ�SG��$��*����q:&bj( ()(�
�����PQQ���i���:�Eh�TMO��KAELu�
*���	5�����t�s���Lm�
���5���m:����U�Τ�����
"�.���5U$�ow`ѧ55�@tiӊ�/c�q)�w�t�m��/�IP~[݋���壢�U�4U!TSlh��ѣ�z����U!�m�h�DQk�d�#��A��Plgcll^�QEU1Q1�y�߿?��g������3r�Nf���=�eݥ:����r�/�sl�ׅPrݼ�|�oQ['1+e�Dk��(3�B�e�dGu]�o͚M7A$�+�J��פ�����Eǝ b�s4?6���6��5̌�'��I_���gĿ.'�x�mi�}��4
���YH�Ǝ�	��pA�������&� �B��F׻�,�uC�[�q0�}Tן#�	�/��	�bφ�OWb���[:�SA.��(f��$O�Uj��r������0$�VY�h��ٝ]Isr}ܗ=0��Pŧ^��q6��S�[q�W�0YA� `�	Ԏ�Xvͣ����)�hL�l:Mf����׏���C��`��5#,m����o���؊�xQ1�LZ���q�{�t��>�V;����̩�(0���%�sC@���OcgW��ٟ<��\����r̞�;��P�3���p^+�f�)�Y�5�9{gw�SG�����e�.���wO{2�y�$IDG�s痎�����M�S���3l>^7j����i��-�TMgF���;�_v�N��+���'��a�Q=�m�i"�A�U��k;�Vv�_3HZgb�M\��.��:;�г��^�S�s���c"�Ӥ��d��x�j-�!i-C����]��?ڟ������Q��h�L��"�։W���/ܦ�F�ߞkC���pM
;孫ta� U=T����ϏF=�fdjyp���Q�n��+I�����q�wb�\�do�A���#��j��ٝ��'7�Ds�PQ�7 ��xz�I��P=�>駁4�=C1iQ�s���pη����7;�%���I�I�UxC�%P��L����0�50ZeVek�i{�"��A��� m��	�)�MԒ��,��(�g����	p4�|!���fx!�.�#cl��/��J�����"���ؚgm�4��n������*κ���c�`�
�~�B��3�ءS�I�����5}��\6 ��ZԷd�ˮO;���K�K[�q`�w���n[ٳ)��b^���8s��l4�B�S�W&�bg�Z�Q^U�opt�q���͆޿�/�;�&�	�_Z��i�B˭ӳK"�,7��S*�5<�}�]�2�s�]"k{ 53��"M��c*/����L�붩5q��5�`���Bv�S��T�@U7�OA��)���։�R
��c`�`������G��W�����^t�
�b��/����vt���� �lΰcu���/��
ρ�[^�RS�����A};���������sM�G�eC��޸
�e�T�h'��c$��p6!� ���V7mj��^��$ST����	f�ZI2	-�\d�^�/)jO��ֳ�F>�vD����5��7�ݭ�D�2zb�՘��m�h��ڝ��D9��;�qb���p��YjJ�j�5���^W{�Ϝ�vIB{�M��s�^����6�w@A+��Eޤ���#��S��dL���#%�0��R�Iu��W���ԪzY�g��N4^q�;ۯ��V@����Ȏ��ty%��F��j$ ��W��r��N�^���P�nd�",j�;A z�	仸��t�q�{v��F���ŭC�R�>���;o"`+����u���@����i�����򼬚��)ht;�f�k%/�(�݄w��.�^6\ٍ���M �u��΃-��ީ1��3H_���W\�{j(P��o1 ���f�����9q?��o�'�v#�vɊ�`�[W�%˧���h',������\��Y���Db)�sS�4���}����q�>�����Emzx(l��)��uFV�A���s�:U�H�n� ,�?u�1m� �B�T���+��֮�����؟A���'R]�˓�f;[a�u��Մ�쮼{������=pxW���W��;D��I;�l�k��z�קS0�7:E4���׺e�X��TL�f��5�~��R[�.���S̻�b٤R)���4����/�=)}���렽v�#`"�����������Vm-G^j�<�O<w�Ӱ֊v!PN'���vJ޿��G��������n�ָ�jI��>���t����x"B��<�=�0��R{�MN7����&�v~����Y_��H�A�<݁z�=9��h��V���8��q�Z����񕒂��6k��;�M����-��b��Ʃ������Q�7�D��q*F�z-+�0��$�e��),��c׈ӆ�7$��Rf^�����Ɯ��l-&ܛ۹Z<C�F-��:��?7�9�)�7�~��>��
طǎN}�����j��rv�4�E�W�-	��p�d�D�h��U���b2�Ts�j�4&~��z�5$$W dIRGS
��f�l�oI-7rz�������g����D�\f��%Z�l�3Q5ڳ��݇Ƕ���sN�Ty�Q4#���b�����|��̭�����k���v��Pԁ2�FFN�j�\[?�NEL"�5��a�&��M�e�,�'�뛄�q�q$s��%R���~��uz^M��ng�m�G��p���������#���ƛd�'�Q8d6c���v\=�|��Y4�������m��[i�m�����Ǚj�|���6{�m��7Պi�0��ǜ���4-�����ئGZ؞���{{�	 l�-}����W��D^�����	c|
����
�y�_!���{QG}30�N��}/�RL�����P��U���p*�'���C�����I�#��n��;l^e��F�G�]}<q���=�v3�Q5jŲ����.I��i$7�GU������P"��)���(8
�ִ+-1��ѳ�'0��:����J�Z�4\)����Qܺ�����4�ɧ�wn\�����h��2.��}�q��:����M���I��{hf�m��jf�v.݌�͍%���f�[|�e?yۣc�c����G��ʯqc��c��Π�:aJ�xt[Վ�kl�-y9����Kǃo�}��@�>=$w$��M��F]�U�s^Ċ�TV��Q �W��f�Z��v����a����r��ԜL:��r�Iy=~�Z���hoXQ
0�h��]P̸�x��w������5m����6"���R:Z��	G��z�͞�f��b�.��!F�_6��l�8�=�r��E*�G@=T�氀�+�b�%Y�*b�q�O��'wR1p�`� Q�5�Tz�=�Oi�6r�3�i�H���movu��t�R!|#�kd6���1��"�9&���*����L/,�א\��3�I�}�
t{~ab�g�ģm�%a�V{=;7�'v���n�hk��o�u�/\t���v[�uvf����k"��6��:̠��'=���tϮ=�����y�*9�.�ǝv	/-��Jk��׈��e��h�{N����..�K)o���x/�6Rj�e��DZ��g>��:1")�.A�<сb8\Nr���=xs2hdѹ�0��យߩ�����O��q2�������x�x	��z(��}������]vCr3���w�ш���}��fzVm��I�׎��T`��)]��B�J�]�t��(`����]�0Z���B梥�.��W�v�ER�z��Oܷ@y�پo��I��[�	�#�Q�"g����l[MMf�J���
�e%YʕyB�=�pw7��c�ahy����/]e�հGx�	�XE�4;%�5���'R$'�5� ��r�)K��
5yZ\������`E�+�d��f�6�ˍ$dT��5e�B��������א��/��/��<*5�x��|l����7�8�M�KK���>b�}���EC(kˁ���p���c�ID��c��V&v�4�v9y[�I�	8���p���{KE<l3����J�r�4ԑ�$UX97F�%�Խ1WE>ܥ��6�U�<�hq9Yԑ���}<�ǚf߬S��5�R�g4��U�g�l+fHXٴ�Eb�R�z�q@��J�d0M��Z�\yt���ǈ�}�9�̭�P��l��"�'p}r��ݩ;��s]�37�7Ty-4�HK��^Z�sNx��yn�&rx����2����,I��#�'^�IU�*�#rT봑�y�&o{j����uVև\,��Dj���?_:�tcε�9C���k���oZ�z���e����(��	G\p���"�s�Z#�U���E':�p[Ƽv��IM�����k8"�Ί>�[2�ə��5�yݐ���Q׎�%XF�V�*B���}>b�)�A�E�kd�l��4Ƌ��w�<	9�4��x�V��y�uZD���!����G5mx������Xy}�/U��`u{��Q(ąx`��,-ll�3<=�B�/��V-z��"�=�к�w�G'a]�g��s���K�&g��^j����h5d�u��a2Fϲ��� �8#�o�2q#��H��J��W��,ia/�"��)~x����JÛ'ؓ�݇���	\K}�l~0ha��b��,��ī���2�Ღuѵ�@
�;�*��.��/���u:��1���y��ϕ��5-�5�VF%�t�!�ʛ��y۾��u$�d��ԛyt!�E4�ַ�9�<��v�Lt��!�y��B0�f@�ۃVV^k9+H�(����^��w|�2ܢ�<?#�M��=��z��zn����R)�M�7��	3��nGp`WO4{�Q�lS��!�]ë�}-�1U(�L�DW'�V'����o)�w8M��IV�r-Y*4���u��70����g62�âj�pL��vEΤ�rI��������G,��7��tƶ��m�e��ła��aY5#Q+-63=���y�ڰ��4ؾ�]&�y}�M���
*��>�<$J԰Tt�=���}����n�6h*�2�$eP�W���2{-�ճ�.��-�:��44_v�9l�Yb ]-�n�h�I$��?\u�B�����ڍ�x�jn���s�KS.����R���$��'	��w�Ǜ�ou����!��f�Fre�;,��c�'��Q�rr�֯��Y���t���'a6]XD��l����1
Ϟ0]������8,���}�tU��Pv����x@��n��5%I���	�bYz31�ŏTX��[-5�\���!p��ׅ+�-�#m<{l�4	����]ԙp�q����<$�����@���8'�P�+v��}_\|�ʠT���d0,����]��<����4�Av��C7˩��Wk��������|�o{�ōr�q]c9.��?X�Ьf@?W��t��<}��a�`\SJ�J>���7=��+�;����5`�X!W��_{a5͖UaE��ˌx<8f�(w�l���A��Ŏq1�v̎��%6��sB2��U�J$�@���d���z��o���C��B	���h�l���GG
ݬl�����Mp2�Q/��T��>�	:'xM���^�VnoãMz��d�dw54���u��4t��w}�W���V|�k��t}�q�\g�6����Mif��ƺ֗�������iDh� *�ޢ�"�_{�! ��
�|`�g8��������&F`Y�fA�`Y�f� �FV`Y�fE�aY�fE�FeX`Y�f�aY�fA�Fe`XdY�fE�`Y�fE�FdY�f&�`Y�f�e�f�VdY�f�d�f�V`Y��fQ�d�fE�`Y�fE��Fe�fE�`Y�f� �be�f�dY�fQ� � �F`�VdY�f�e�f�dY�~w����� �F`Y�f�`Y�	�f &�`Y�fE�V`Y�fQ�VeY�g�W0,³(�0,��"�2��3�#2�ȳ�0,ȳ̣2$ȳ"�2³(�0,ʳ� L2�ȳ"�0,ȳ*�0���(�2,��̫2ȳ̣0�ȳ"�0,�ȳ(�0��3
̋2
�"/�DL�)2� s L�3��U̪�� *�0 ª̪���=�UVa 	� &Ve 	�U� dUf �UY�0 ª� 2 � *�2��*�2��*����  L 0��*�0 �0,ȳ΃�2,ʳ �)�dY�f�g��f�`Y�fE�V`Y�f�9dY�f�dY�fQ�a�_�i� (i>�@F!U�DH� =�
j�9m�_Ӏr'��T��֗���t;����2yEΔ����m�yͣ�P U����Ǌ(�+㔁PW��>`�}�A�������=��m��H#�ܫ@�`�ܘ��Q3`)׸:����*�� �(�*(�D"���
,�!@ !$�� �	 �B��+
 H��
�+( K
�2
�� (�  U�:�A��������UDE�AB���='`�}��xv@m��,��1߹ U�w�:u�oq��P��] ��As��K�p� �!ڇrtٯ�(�
�
 
�(r r~a��`�UQPV�à�B@Y �q�����j�P(�Su���K��V�ʐ�TP U��i�v�yq�� ^A�)�V�g�9�w�;�Nai�8���	����r P U�0u �ǈ� ���1��BQm�(r(OM�r�H6��r�츠 �t�"`0��@����Wf�:��QPW�ـ�nodQPV���fw]�:����d�Me�����f�A@��̟\�����RE�2T$�k�:ԴiJ"��$�P�"��U6h��R�(��J� ���di��ERScRH�P�Wv:б���AX5�eZl1X�m�[f�ҦmU-afePf�Y��Y�i��1J�h¶jkT��fk,ke��m)f��l�i����PvGh�kb��m��S2��iZ����m�����5�ffH5�Բح�KJ�V�kPb[[ �֋1[f�kXʖ�X����������YQ�[-�  �m�w�;���H�=��P����zw���ӻ��zu;v�M��y����^�e�;�{�=^z]���E����N��Os�9�ν{X<��g���=u���ѻj�Z5yv@�[���SX[([,�   ;�>��oc"B���B��ׇ��(P�B��=
(P�>�E��}
(W��Ϲ�X��T�JC�N�=�6�۔����^�۷�Z�����z��e���ON�����ճlz��i#[k-�jcE����   �����6�綷6�u�^�zr�락n�����'[�;��WJz�ݱ�ڭ5OA]�yurt==v���z;��C�V�^�������v��Ԛ�^���d-������n�m&�L��#d͍�ԙ_    ����}��U�^��/w�����t^�zz��GU�[۽뻗�7�y�ۻg�C�L�^�w^��{�u
(�8P��: �ػ����vv���bգP�k[h�ml��c�   �A����ѡlfL	>��֗ UmU�"��Z֠V�7t�[PY�Ԯ����	uK�8W@ѺsR�ұ�VZ��H�4��  kިu�Z.v ]�θ�Q@3 �wneUV�.�p�Ts�GJR���uC��\q@��dm��
\\U�Sm�J�l�&��B�   x O/[�5A��+�7J��2���F*@р{z^k�  ;�c�C� ��p  ;�Z
V�0J�+[l��mY|  g��s���>� ��� t��{� �S4��=N  z�� ��G@�[� (nv�ek-�کZ�m�R��V�_  ����B��w���@���z֏9��z�t� 4� ��{W ��-ph= ^��� ���[� ���GN+���l�hٳm�m�  y�� � @�ǥ :h��  �L �:��� �z  k�p�z�� ��� t ��Oh�)P  "��F)IJ� �����E �)�F�JT   5<@)Uz ��R$̪�  M�������������?�e��+#0�Szf1m#*N�0Fܻ��D[N��+����<=��������m�o�6���6�6��6�6��m�m�cm���O�߬���Nѿ�%S4����)��)�)T%�����
D��2n�B`����*��e=s�7y��u����6nVp%��NVh�p�)���ܥ.oҚ��ĖHp=�/X�N�-;���z5�Q�e�͋gw巿hJ��zʦ2K�2ȕ�5�cn�wL���yF�ݙIh'A�J0f��X����u��u�s:��I���``�N�V$��12�!�-�%R)���w��4�2��Sm����	��^�A<!Q%9���e�Yݑ��QY�#�FU�Į�(K1K�
���1�M]nبI�=�rűs.@�����E��e��\*�cX�%F���3V�N���%���S�1V����.�?:�>s"����"�R�卭f�;@��E��UHl�m+���tu���͈���j�P�5S���\�����[ml�����/���[Wηxk�ì%pǬm*�ߥۙ��v4V�tT�զ!su /:��Kd�y�K�[�������6�#��-��H�pص[-��2��Ѧ�dq0-f�bsP�.�I.ݤ_�潤���o�̲�nmaO��e"SY%*��`���M��d���y��ʱG��V*:�ʀũ5d7Z/3m]��]�52O��]�d��6���c��E�X�]h[Vf[�S7���6��;C�(M��7/7r��zssR(��'�hv�ۛt��&�&n孩��i��b�Xv�1J29����Prӧrf��ũ�� W3$��52�xɺ��b�Ġ���p8��Q�-��Qc�oX�@$�OKnęz!NȨ:���(n��90���N�\9��;V�M�#rėk��P(��r�뎂��R)�3s%�B�>Z̫��Y��Sub�$	�[uj��7fM�[��`��[����;�.�d����ՠHdd�y��c��[Ff�I+F,��ցi����q�ΝPY��φ�[�E��u���ڑ�v1-�܅5u6�Y�k��V��Z�`�"��e�Z%�øj蕄j�tdqKե�y��Jv�:Om�w!�g��3Q��� �FDp�Ʒ pdS*��8i%����2Y��K@xK��]vH6f���fDFY�3w����T�o2ԡ@m,b�o6�p���⁠�c̔۵/&\�&�����Fa4��	�6fP����4��Q��iT%�F��n{r�%�Jql���`3��%ج�؀l|X�į�}�N��Km<#�>�D�u'z�R�7r�tCo��شҶ�`��d�v��T���
̡���R���%��ZH�6U�ܡ�{Z�s,�Vܗ(��Z�L��t�q���Y#xf\n]`�����/�4ܴh�>ҵj�`��C�S�N�I����GF-�ڏ[HX۔�/FǸ]L�UȄ�m����X44�q�Oom�'�.�v��@�İ����ͫ/���-�M5n������f�N�)0.n���^3��%�������ʱV���wn�/����$�V��0)-�M+1|������b��I.Th�y�s�F�;��԰�e�B9aL�tM�Դ�<�V�L�2G/MeҤ��(ӱz��\�G�ը�{j�;�ih�&�� �\.�ڦ�c,H��t���z3q����BQw�1&P�+VKwm�lV��!**T���R��eY:U�)�o~h���h�\� 4"@ш�nV\���Y���m�"�B�T�E��H�KW E��܄[�қ��FJ ���f�=��y���36��Ub�"�m�**��0��i�i��XB���j�nfPH��`��N�h�dU�6Hl�(:�	����Yϕ�)I`��r�-���ee�����I�.�eԽ�<�t���:���VI�U���8�*�X9�mY�u���p�\/H�i0��U�E�KeM9r�'�i��.��7��\���r<խ����X��%UpD2�N�3n&�ȫ�E
�ñ�ZI\MV��]�]�z��y���F�utr�ɦ�w6��"Eu*J(As����tU��AI�-�I��utә�}��v�n\���4,r���e�;�{V�F�ie(���Cn*�u�h"���3��hH[/r�nܬ�ڝƚ����'�/��E<�Q+rNRFk	�+���c��[Ȁ�D�]�n�H.=���:n;7`�lfҷ��vⱅA
�Rق��U�ޜyY5c���0ӄ㧕�%��ݹ����F�Yȳ#Wz5�&4���F��0c3^�r����ǗWo[�n������Ɂ�����X�Ռ魸�c(娐[X�`�����B�J�)�"�� �����s1(�,�z2�R�%���ܭ�D-��v�naĢ͑[��f�LP��ʱ�K"@�9�w)�����Q�s�gb��33S��ڙD�5t��d�7NƇ�F��̐��,�ܠ�YDӺs��3E��a[M�A�N����r:�&#`�Q��PUTVU�x��7m���*�j��jˈ�pPx��R`�%��[s]�ƪr:߀r(�Sİ��+u@�7Ri�Ǳ],�pYN��۫t-
�+`"��!�����n�Q�0�CF�.�\b��*U����T�֝O�-A����@��N4h]JYi�<�݈]5��%`��׎�![O(JIi��uzv��,]�Wd�RJ*W7n�c�̃6嫅���^㷈!-��w\����.�;�-*�Ȭ�m�r�����&���e�&�gt���NP�[�գeY8lHN`�D:��V�ś:a�ꊮ �⠮`���N��)�MQI`�[���#�i��M��f�5��)n6�M	;����SR��:���)���n0Z�{S��Ք)��c��$6�9k4+v㕯�@b��)81��K����E9�՗F����E��ci�/5���j�[�;�4��e:��t���J�B���ma���K� Ln��͆�m�i�n�e
Ƿ�JA�,�J��S;I#�@]��
��1Y���L�t.	��4�}58�����E��1�s2S�۟;�IN:��l�[Wu�J�������,��4t:��lKh�`���8@a�w�#��M�Imc���i렐���a�Q^�ZP4޺����ȬU�}Jm�j�Ջu�$uM!�cl���}7���A�^�"�--�9���b�w6��P6���X���$���c`aHTZ��r¿���;b�4�ڽ��E���Y�Et0]MUtJT
h4.��6�(��X���(�4�ڟ�=Sz�^�l�ȴK�+*�Xэ0ݩf�9j�� ��CZNi��N��em�Z ��MB����Jv�k���U�n�����E�iY��r�v���S)1�F]��C��0�����a�3	ZŽخ]�w�:�Uhlw,�0mi����ҫ�`���M���D���8���
�F�s��6٤]i#
��uV�7WK~f��!�R3XۣDڬ@	�����cNIp����ƶ��R�V��L�+p��^�b�:�b�ZU^�H�A؋mMֱ%.��72�4�Z��R��;��Ӱ�P�I�N�p̦͜��D�Yz��ov���T�BӸ� �\;C@�Ҳ��H�H���/@1h�x��7�̹��{7�����`�����rM�,m���ʳ�~��T�Y�&t$Ab��%�˴�*�2�yj�k͸쨴Е�&��q�s���G��V�j����p�!l��Q����[��L���+V����	��%C�#ݻ�g��wk ��z��n�3j�ؐK��A6�ræ�e�����LW��߶�!��&LhV��=9��I{[X�����K���Z���8uC�|D���8,�I�=❷���Q|�O�:#.�i����I�j��.���*�Au��+�[��t��u��1��l6Vo�J�l��#U���� �����פ$?��AbR�Z0�ml�'t�����������KӁ춝�&ڴ��-�0n^m;�ܫ��ko/�4CgRѠ�ic�h��[4Э M���Ӟ���ѝd-���slӱIP�R�94Pā���f��aS���d/J��#Z�����H^fm�v�G�6���{�Կ�����\N�n3W�Y[z�9A恓r�ra�Q�1��Ģ����A�`�����V����3iH��[���@�U�^����T�Im�՛^#��%�cA�nRŻ��r���J���7"��ՐC���Acz�<�A�!�V�/Z��&A�0���fe�묨/F�n*XYRl�Z*�]���k�d��Ĩ����t*�L�r��v�7�n�Uo.K#ئ�+l�3���TQ��ۧ�k�U�a�·@*:��V�(<���Ce��*�KstM9�K	G���[+"�ui�VS��L=n�eBeI8+D�²U�gw3CRر`<��I�m'pR(�i����;u�w��X��'��V����9���IJ�6���
�ie�u齘�l�*�5a��Q�zma[�U�Y �ڸ�P4V�UqL�du*�V�],4r4�U�Ƥ�4�b;ج��M��`�N�rbhE���i�1QZ�!�MX��IXn��+Z�6�q;�b['"eVJx����,�Х`����-�ZPױc�I���f���#30`�ɪ�bM�;�i�z�X�Fm�&�	Ǩ�ڨhW��XWp�Ӛ1-�K�A��e@J�O76�Y2N]+L;�i�4X{A�.�jz_ͭt�I@�$�c���Y�=U5"�"��쁬n��f�^��T�!�qmk��5�9�5kP�;yW�gq]�ҥ�F�ʅ�g����ݽˇf���u�{3E0��w�� ��:�0�����4�0�r�cMk-����[F��t�ՑE���(¥n�Y5maR���ݚ��)�F�nR]�/�S8�6Grcd��Ph���-K��Lb�TA�9�V��r7H�����wff�z�@0h��^�+Ǌ�uM*�����b��4+L�>xe*�
=͑��VX�����N�1j�X��aQff[���6ɗ��&�Τ�	�o+.;͂��?AK3]t�f���j͉��q�˸�6�n�f��,r�U�nv�#�Ňt:.;Xp��jX��ŧ��"�����v�����۷kl�n��:7X0&ؖE2�Y-�,Q�Y�ҮփR[��dU�OY�`XU#ܼ8����e�K#�awxȕij��Y�kK*�K�-��[݉��I��0�������Èd�1�5cb���l3+$$7!jb�R�d�,DX����xt]]p�L�h���e�a��bReےN�e1z�u�`�DХ�xa-	��øS-��Ji���g&�q�'+ l����wS#�u9�f�lH3�f�hea�lE��"��T���4����A.����Kvn��j��,�!B\2�[q3a�����Xy�N�	)7y�I�������0w2i.�Y���)�O>4�vu<&�M5r+֔�u*2�����*���Jl[�r��ͼR\&�ClR���V˷���$�#t�6�ST���jcmmG�6��PZNn��6��ڽ�v��u��ؚr�1�{&�rQ�ͽ��[���a��-�0-����P�r"��):�W����z/����@�Z��{j�v�Y�>�����S�h�2�n`��M����c�q�67$i�-ieJJhb줍��Jb[b4i�MV�3w^��7t�R�zu|\+,
:�f��ܓ�,�WP�(�xP�9��ʣM,Ɩ���X������h:d]�֕;�L����яi�pK�@��n��HY`k�ǰ<�L�����IV��4f�-���)j���v�f��Nfi6Z���#,Y�Z������s9�1U����ڹ����6�HV�fJ���i`��kD��.��{�,���u��z�X�֡p}wai���Y��l�4n9z��a$H�b�@@��c�df�T�'�y��WI�܄�#��Yh�16ہ�d(��^���d"��2�Z�e0POC;Xۉ]������/sC(a�]U��ékF��1��"P0$i6qR]�Ė����C�T)�U����+E��e,d��e��Y�3^Уd�*YY��n��7k"��ܼ�km��%=��z��M0AK["�Ē��؁S��&�Y0��͗��bp�\������3%Gx����4�ü6�4
��IZMe��Z�	�I��7oee�{�]��F�b��kt�p�oq>��[��e�b���{�E�m4�2����f��i^��oh���yS�6�B��S{&��9�5 7#����3��R`�<Jl{{t2�Q1�4�{�lj���;��C���d<y;E�&���hҚz�K��
�V"%Zxt��V�?���@ $p%m�l���t��5+j�cSo*FXVQ�At2�v�"�f�Cf)��E��m�':֛^�p�kՉ��f��Zא���E5��9�_��̐)OF��E��[H��Z���U��@%n#��,Եe�ٴ�e�i�&
ɥKƖB����M^#��4
2�$�6�[vA��٢�'�q仍^I���PU�ֵ�,8���%�n�ĳNɠ� ՔZsMU{t�l�����.�CL��0�U��ކ�p��m��q�%��Dc8�/�T �谮�G��o[�"ΥxՂ���7��[��cUb̟!��n��"ƙ��ʳeR�̊�f��I���l4+.f-�%��:ъ�(��ln횱��nЧ�z#Q�)Vƭ�Ď��{6�
hä1�����ef�P��D%��	(&�V&�%�f^%� n�6u��1:u�B*��ۥ�G),5kuѹz�VT//d@S۹PV ��ϐ+]�l]�F����e,C1�h_�´�L)�I6R��	��ǽ9�8]��;�>���wC�=��8�__k�f.t�k�����92�f���Z�a:&�0��
Z!
LX�F�U�]�N������n��
+WulaYV_;��U��&CԜX&��}����������1��*��"���G�^��g؝�P|2OO3ˇ8ӧ�>�|��Qn�ju�fgh�Ɏض�\):
�v��Q�PuL�IZU��tz.q�}�l�"�!Af�m�Hi��t=�%�T���OG�)�=�=d0Ƽ뛫l�d�Eٶ��+h��ٳ���o:�-����I3ZP饧*�Xtл�j�u$���!:��N��U�̝/�@NT��1�����<ݺ��8t�2�\��E�>����r���l����,)�� ������ʺ��]�oj��ut���G:Iv׈�Z�������Q L��������g�Q&@�.��u��Ww=M[�ُYeCgc�v&�i��������op�R�3i��R����T};��	n6{�6��9$�R�B��o1��#mfn�:�R8��������V(&`SH�N#]-�q#'ח�m&������A���Y�g���G6'k�Y٫_V��*Lנj�5T�K�\�]���������J�m�Y`xrQUm/9|oش�A�&��[p2���!�$����m��]ݦV����k�����6ܲ�p"�`Һ�+��I�j��%��GX�&啄�ț��.���4���Y���D$�_WT\�v��������;�<���9X�M^djfڐe��:�D�K\�	���o��5�� fT�2����=�v�7�,�x�k��%k�"򈈲��ٖ�,��s��O5<dݽ�^�a*�u��k)�S$�����y�n�>�~5:;�gӈq�Bd���E�yi����ݬ��UK2��bq�0��Be�B{��t8*�ՃH�:�4��s�ȅ4@mɕ ��c{1,7p��l��l���weJ�(Р����#4+�4⳴����
v�qF�"���r_-���"^�[�iZ���3�WB�q�+��B���t��zZ.&
�z�*=}ٖ9E��5�iF���n�rj�ЁGc� �0N6�'��K��Z)��Y���ջ,���	�֠G T�5&��k�]fZ٤�Ø���;"���ɲ���ƞ���'���=���
<�f�s�Jov �A�^�G�f�$��l��A׼���G�����@�)]���%8�G���Y�;�m�XyZ'"��x5�Xq�X���T8��T��F�of�����Z5���4ڴxwc�suv,`p��Э2t����B��/��.�Փ�E����[ڴ��ųo� �WSgt��\(�a40d)=��>�+��F�u��c�Ni��OP�[c&4��́K�C8�뒯`<1�Gb�wwF�
hִ���H\ �IYR�W��בκ�Al��Ñ�J�ޮ7p�&9�q��gL���3�����0�)���1��f,T2�dC:��gziK7���R��S%kaܭsu�;5������2й{���汣��dl)A�FW�͡'S+tT�7xg`//��jƪ������]�ް���k5������u�ig��5�_ ��G��i5:R=V���:Ѷ�m;�өJT6rē����`��*�B����dH��He;�P�Rͦg!�U��B��zrV�܃hP�K�nne;���Fؠ�ش�r�Rp����z��,�����f�ؾU�I��\&6�BD6��1��˫��%i�M/;1װ��V���7qn;4�N�B�B0P�+
X��z7��ɪ���#L𜻤���ZH�͞4*��}���JW��*�s6�d�[zԧ��J<ݺ����bn%�o�⺴]�	Jε
s:zcKoj���c�}��E�Կ��b���D�[�u.�6�_��Xj���
Z�e��sz��DL�s�+��JjˀmdQ�6�r�
��i%��Y�ԭo)\r�RQ��ʝS��u�eW*s]�8sLtѼ�y��ҭ�����)�1��;�hr��9�J�2֮�O������'*�K���^��/����Q�����pu¶�Wl�<`]��jn�2�p�/
�1�Y��� �]C���Cm�	��ޗ�mp����.����gX�Ғ��յ�!����T2����qm�ӫQòނ�5�j��@�5����л�=�v��|�:;���u�5-w�:��p�ɨ��jJ�;)?��zC"Э��-z��a��C����֐n�%�ⲷ(v�ݔ��Ӭ'Ѷ0K��)�g:���]�)vE,�Il�bT/�pܖ�da���I,{׭L�X��{U�cz�m�)�%��GY/j��Ⲵ�F]�X�1hN�@$�ΛCc�KF%Ǝ�Ε�
A�ñ6���q�u�WJw]n[k������s�#-,�˞�}P�n*j�5��`��L��!T�pG���Ғ���×�͕���]K�|ZNe�l�{5���/j�V=ئʽ��ȃ`��C�wVe&~̖�]cw�'���R���zViZ�.ں ";�X�m)��k�0՜C�R��yGǇX�B;����C�:��ˮ!W@��F�&�^Vl�w��d�*sL�}����9b��M�I��>��i�O
��,d�:(���N�8lU詽���(ł��nT�}�4�@�oq']	r��P�(|�i��Ì�tmu�<f�$F+�]�����c#X2�u)R��V3xu���Ύ#���K�]�#��ђ�6���t�^;X�n_	T�����	�/klVW���qb8�%ڹ�r욶��ne��H��[�ͧO����tQ
'���ב]�s���p��Z�-�zlJEi��x˚s�fcx�4I�k,�o`WC2V�n��̧�5N�Q`����Mܜw���F�ۀը4Х(s��+���f��PL	���3 7o#0�o앐oR�[8�:���@їZ0�s'M���`S�K v�5���u�f�f*��xݼ�ފ|��|ĉ��k6wm�={� �87�H�h�-��uܸX�˟�v����:�P3^.�;&�:G�[����5a����;�&v�{c+����U>�kDt+�V��tX��݆��H�J�yةh���jw������ǻAѫ��	���-6!{��'�ֻ��[Œ**��WV#+^�}y���*j��ȶ�(�G5�$�Au�r�yY@�x��R/@� 팃�9n���N��/���G2��;Mr�\V!�H��G�����'B9P c���E������G�����R\��<�:�L���x� �A*�<�����Q��MM�i w/������+��r�w��+
�v�1OTfP�x�<�E�)�5���c"�4�H�e�s��S��%�%,Ui�0���[�Ժ��'�`�ݼ��I,�,���{J.��^�LEq�`���ҳFf��cש������R��2�I\�*�c"��nc��l@�:;�x�%�V0��w[���3���CRH�����C�o�<膬SC��&�®�I�L�s��ݯ����1�,V=e�`�ayY��uC�SY<NIt���6�:"���X�˓Kם���d�yJ70������c����oHU
̽5b���kaV�f��J�%����0(�e1�ܜ�����1RF���d(�"ad;[��QWuή�7~Ts).���wɭ�y ��ƫ�\x���N��>�l:�s���α�Z�N����@ڱg����%��4�)7��h�y�wR#ch�eD�M�,ق-��c��b����<+�RޱG3")=J��kX���BCΫ�8��m�T�f\�};\�g��H����gA�N����l`���ONM�O ������<�S�]qx�"M���l��;�ν��ɪ���m�Y1>�[��32o΄�'IK������=�aV#ŷ2R&/jɛ����k3�����&T--�sD��Ŝ�*.���2�J�Y���2�{�l,��������C �Uiĥp\k8��}xWt�u;�9D/9'2H��ځ��l�Æ�4ô��θǍ��_&q��7y�Pљ `mk׀w�}&)A��O �x��d���P�a�����U3H,ҡ�?��ѕԸ�6�t�r�sQ��"��),u�'!,���ǘ8���=�X��)9���Z��R�-t�*�ME��U$#���[���T��lvt�/�ė�|pm��#)��V�G�����vJ�n9ɩ�TdJ�-��K���3gE�;-
K�ŒwZ�A�P�|�6_/4��\�I��2��5�-�[���K��ާ.���-ҋ �tȷV�d�@�,!���w:n²�ޥ������h=ݝC:_W]ܭ�Q���{�$#�o�W3k�\5pm����v<y-Gה�k�}$��hڱ�M�9�X{�N�����1�&]�#%��;�_ �,��j�)3���S��z��_�T�wó�;V��g������Mx�_a
��6�K�Itm��#�vK�b��Ʋ6����IJaYu�]�S@��M�1��S�3VM֎��o	�l5���ڙ������]�.;f̶�i�R�8�bռ��nʇc�S��k�l5�����C�����Q� ��O/i��$��37/]�<
���"ʫ�|��njL��r�:�ݥ}���e��:N���'v�8;x�\�]��T��[sfno�V�dT]r`nʨ5M�wx�U�sDY��r.���4R�>k�%u�-�8M�l�R��b��c�w�u�Ү��0G�sf��WGo�(\�!޼�7�2�r�b��E�>Y�G��0�z\�A���t.��[4c��I,g�	-�=��vVF�!����f�R�z�赳g3٨�c�t��E	�z���x�x��<�����S������5�q6*r�gU���7���ʥ�w"�jP����:���Z�2ɇ(Q�s�M�
vUE΢��ۚ���l#S}�Y��37���3�juK\p�A��+n�����.*K��30��0ǨS)�F�B�I�	仧�tk�Bį9i̔��r��b8���F�]�Y��v��fjp �.I�T�ۑs��Ij6kz��]�>o]�xW>Vt *�>}YC���5�w��owzY�z�� u���]%_.�|8�
�D�U�+u*![A��G9��p��WFZ�|ܛYe�:�62����6_�7ןl�N�d�݉rRj9��p\�q��2��U�gF�6�(
Q�]��Sj�4����������tm\�q�o���T�sl���3�bY�λKr��lƔ9qa��h���L�l�Yw�W�(BFW��NGV�����Fر�]Iti���6�^B.H�c�I��,+t3����.��y�}6Th�����+[P2A[��N�:y7q(E["�Bj�K0ѭ��z:��y�\2E)�ѽ�m#\��:���T1
AP���Y�L�3i��M(�V:�F��
����N���*�h�#OA��cr&�rI��˻�s�l�y7^A�7��&e�߂�C�_N�.hfG�u�Rh��ً�q���̗tvJk*�mؼ��2��5$)��:ΏN���T�����aT�7��u�`q��JԨ4��x��r�$��Q�Lj���o�R�z� �/B��"w�ĉ-��,<y�ތ�F>��gP�F?���2�E�䴏�W�^h�R�9w��.u"2�ɻ����%D9�e�Yw[���&㘗*8��J��F�o��'����y]���ӥ��Pf�u7��lGi�up.�P�خ�|�k��o�K���c�ojT�Ӷ�36W{��}����AA�띘:��3Gº�4>���`ͫ�G]�M]NnafR���۝kQ��ň��L��ӣu*'a��u�F��Y�z&��u��X��oe�+�.(�#h��Jveӗ�]K��\��ޮ�X����t7����V���\b��,��P�-Y%�y[�b�6%u7����)�w��.1���խ��IX3i�Ռ"��ΥA���W�CـZ�f�n���ԫwms�{���:w��튼ۘ�k���V��15�>���N��Yo�-��RU+�,�(qfV=��$( Zuf�R+N�|�X�͖�ᄇ}��{�b�]�3$�K;o>�7,�0���<����e��yΕ��d�����|$�gS��^-[Hm�].��v�Y��K�%.������9+�"��|r��PII{����y�4T��IE}s��.��gX�qۡ���&��3.l&�}�֙|Kpg"o~Y��E��mӍ̂	E���Æ�ӹ�%�h�yָ�+��3��5ng;k"�C.6�Зhҙ��qtz�刍tĺ�-&2�I��e��N����ށ�	�&>�p�dz�����z� �ۚ�����a�YPG�2n�wu�[@u�7M/j�AG�j��S�!�s-l57�i�G]�}�Q���<���7-�ܖ��4
��ǁn֌���d����s��s::�0����tʋ~�9��ܫ�m����c�Z�����:��gm���d�]��#3S�&Y�lJ�D���&}���M^�S�t���${�V-دv\�����۷Q������n��K�Ο$�'p�0�:7��3Ӻ��%�T�r��;�3��b3�P��`���+^1�&��EI(��
9}b�5��6�{[x������{|��)ʱ]ȓ�%�52Q��6�)6.��N�t�����
�m���tN9R-qɛ'gEY8�3r�%܈w*T�-(`�de̝�Sr����BJכ���1&�B6c�6��R_l/�H����o�l������������{����������O�������ތN�1EYؿh֭�35}Ҁ�L��<��6(�g���� �V�m��J�w�y���#�+{��h<t�G�������2��e
"�I"IdB������{&�ڰ!������ݣ1�Wb���@�w�Xܷ!��Pku-���ư��M�6��l
d��Uk�E��2�X�Μd�[W�w�l����^vq`]�VMa��pCtX'�Gu���r�w[�BH].R�My�)�0�vܱί)�f�<�s�F��j��!�V�h��)o*[�{�8��4�][��q̠�so��N�C$Q��S@�k���5��i�
W˃�.��dϢ9]���]�E�3o�U���W�� ����nѩ�{YQA�.��j��[괩��$�W��yE��.�4��5�)')˥K �|�d넌n#Zղw�'#D���'<K�M_U��śЪ�TY���Hő�Ύ�,�oW@cQ�1Һ�rO
]z.oP�����:�k璋k�٩ܠ:e�wp$C�F1�-�2ARtn�n��	:�|�42�j�*d�Ī�b�Fspu��W�ƞY�dr�b���Ϋۖ�e2�f����/��5@��cy���]��"����/�r��GS�\Iw��d�'�mJ*ڴ��!]�w����Ṇ��qr�7t�hʲ��٘�F��%��1�glG���w4i�ح�N�%#��ML��4�?q�o���BpTT�ԭ̓q�6\�q輠2.%�Z�uwQ�u��)�v���� iIt�bwL��&vs�]���܃杽��ĉ�]>ؤ�3��q�x���g5�A�nSѠ��qΚwwBvB|��a:mØ)S9����n�r8Y�hܺ|����SǼPǋh���������U�q�i̲�fw)����s�ך��uD�3��)ff�t(��Y�))Y�^�[�c�%$�ʎ�Mqf�͵v�䀹4�Z�'63�o��X�G/�s�3jO6���P�c�"6�݆�T"[������]S��bzN�2���q]Dk͈^��׭��L9�ݕ�%'[	�,����yy���\	i���'<�K4;�\��=�ܜ����\"�=�N�V*ƻa\�}�o�S:s|M��{�_c�i���*\�t�˼�rhg�2駽,薺[C��)f���h8���;��z�7��Qѡ�b�S����oNwEp�ڕk�YiL�u�w�-��EZ�ѾVr�f�����u@��|3r�xTg�\e�)0��v�ʾ��c� ��q�v��vP��C�b4͕�����5�$GL4H�ћt�]�;���c����W:H�Q�$��k{��a���N�6�&q{�0K��oe'%:��M��7�?�ѓ+m�
���ڛ�y�S	����{��J�ζYi�.��ϫhX��@�ЎA|������'c)Д2-}�z�thz6�r�\����y\_>�%c��س�+����|"�F�A3�[]9Z���P��b'!����嗱mlIc�V�c:�ltH�۰ �X�ǰ���i��'J�+���E8,+\#���i�j��㇦�:r��um�j�LI2��S�SY\�%�G+�ZjU�-��#0�]A�~�6VP���L�I ѩ�4%���7HȲd�D9��tJJ��z�[k�ʌ:�(�Ӭ�h�ʳܴ:j�ε(֠���{�|;�5�����1d1cݴ��uh�8��<N����9;��^TCN�;{���JS�٨-a�^��UD.�M��zQnZ�Q�|�^��4s�:�nZ��L��+H�;kK�K՝a.V;X����[���@lm��oP�$�z�n�]��P�n���~��1e�A���h����k��l�#d�O�nJ��Mu�?Z�:ȉ@�_8.$^ �ɑ���Ex��ب��#V�͔��n�+�]�ٱu�xX���M��t�Y�X ��Y���+�(�b���/�֜r�Ra�,b���F�=Ի�����ۮ��ۂ2�u�C�tܴ���H�.fJ��'���f`�u�&�uV5eV �Z�R���k�Z����W�a��R�L:�e���9�n��S9�=a)M���S��AM�T�T�p��/ys�����<��7yݎK�hLr��}%tIvh��7�俕۬���h�ր��f��D���V��/.fB�b0^)Wql��.e�!<���1�n62��ʎڭ�9\y���[���J��
g���N\iI#Uݗ. /Rͼ*�$�L&*�e[�g�	W1"U����ͽ��ܾ�t�g�ۖ#�w.�]�&'Yi[�CKa
GU���PR��m��&ݚ�o
�ϓ��`VAGO )F�p��0�7���<�u^�I��n�X�:VJ���.��֙��CwF�j�Ѯ9/.]J̬�Z�ހr�`O~����}��:�_rP�,Թ�=z�?e:�4&9t2�bFnV�������F����P+Cudk�"p�M�ĉ��8�>��X+�щ'G;na\'$�ƞ̀`���8���3il��ƉW(��2�5}s/P���Y"iz���Z+r��r�5�c@V۽Y
��zn�|�|����2M��$�K�������V�N�Q�rɈaI�f���p�8���+K��u����f"��u�J'K7z<�v��N�Wf3IIQ}���/�, C�:	�k_�P�]ٻV9@.�hE�]�&-ӵ�ON����Jޝy����e�Z��ǜ�Y�j��pL��:^s3����L��FEj�-y�kQ�i["�5��-�LYc��s�oe,:�5o:a:u�ļ!Vgbق_��x� 0��^(�}g7��ң��x��u��U�aٻ��S��xT��p�A�B��\4Т�_f�[Rdj�g��1t)���-�U�n!]�-m\k"�ڳ�LD�X�Ye�)��� �	]��<��t��N{y ���wd���P���]��9g[��-Q��v�'��]�)n>�+�+3%���j
���+eG܂lح��(]�&4.Q,h���8#C9E
���7���Ih�{r�l�L�won���=�æ�N��h��c�v�8��ak��@�CQpbm	&l7l1�^<�wN�	1H���X;0r��w��$tfqp�5y���*��K�Ҿ�U�5s��T���'1�H;�&�L{°t�u7��Ww W����{� E�v������|�4G�t�cY.P�;f��=������K �д�Vsz��Y,�<��4�o��5E'v���Ě����hj�����@IY�Q޵�Q����Ul�܊��$Rb�?wY�K'pE�T®0�M����q��W/,�փ�ƋCa%@^r	�s��5�% c��KI�yչ{ة�ޙf#���?P���9����e�vH���%.���aT�E�������
���X���ų ��@�[/��T[u��#L�v�J0ʺ�N"v�p=M�0��@�
�L�h�˥Y����e�h|+ �pp�|�}yf��E�P�l��k�5�a26rt��2�]rIAf�p��S��׎P�:r`���9f��YĈ��`��A�4���%6�@W2�� �q�����:5��"���-ѥ�}{�	.��%���X6�#�3*u�9��a�{��xK��Ua�񕻖�a(�H�XФ����ݱd^��"�f`/N�3y�M�wX'[�8*��b{�����Oo�Y�����%�ɛ,�U�\�4/��S���P3~��Z����w��\�"�r�+klB�j�;g��wti7|�IQ�a�Ց(��g"�@!����Tso'0��>����n
�ְ��;M�Uum�5�h��3B��-1��"�W��e1��'i>4:\�#b�>���aH�N_RJ@�rѼۥ�@F���&�*k������9-Wp���tW�\�n����v�@�Y6�q���ړ�Z�`@�մ�)��ť��΂yJ>aQ�M5X�(�,����E����'!
E ��̛�"W[�*K��	���l�4��t�뽦� �3l��b�0G�a�-�,��ܾ ��6����v.�lz��2��pؗ?�:�n �݉T��{FX����B�J�D�*��1r��]�հ+76u-R������f��ZI�W�_�X6cH�٨̽��^��R<�*��K)n��{���2:�or�]�h���:-����fb��:��i�M"�i�m:	�u7W�v,W<��#�Vkwhܒ����`��W�5i��p��Y�1��G.���T������2��>rt��.��Wn��ɚl3m��9͘똩*4'6�t�i�}���M�Z���Ҕ���s���6�l�U8s1A=ݮE�:4�}���f�ݧVz����"��C{*����e��=�pi�`Sd�-��2�EԬ	��&0���T�Xj�v1Y@wS�UF��n>�����V�u� ����ٛ�Lv��1}�e�%��)��M�CΥG�@�|t9��:�s-c���V<�4�r`�;y���;d�ʩ�S�F3��f��x��4�q]/��$6S��Zzq��u���[m=��Ŏ�;0��t�m��,Q�������ȣT���m��1^eDH��L��lgr�f���E̽�]�H��^����0t\�16��ɴ�#�YV.8K��4]�yV�t��*р�7U���+=����A�'F�̌����.�m�.3�żԭuy�z�Z�h][��.9@]^X���R�'Ve�i�������W])s'`rU7\��ɝt.���%TO:b�0%��'��6�T����V����s���&�3��a,m��� ��Nl:M^]5�J 7Z������{�$�q�].�]we�5���Yq�ՖBVs��U��� S�_R�����F��Q�r����V3B#6,�V�G����z��LN�T�u��ʏ�
to��[�KYv�Y]�;�n@f�P+Aǃ#��Bz��MVQJ��������:�>���5��/h�r�#�E�Ov��2�{g��F���l��r��}tt�M�t۱$�p���u�XW\�� ���wJ�t���g't714hmۙ�J��ֿ�^andӔ������2�0�s�� �V�*�K�Žt�p4�wG�m#4u��G:J��)4�ѿA�EcuX��ѱ�* �8��/1���v�і7B�2,��p48+ 	�w�VܳV.���+���!���7����B��цkW)Բ�]�Vvj\�i
T�@T뽾��Ar��%�
�%fj�Λy��-[�\ŵ �(Ծ����&lg�R�+F޷W�#5{6�=��$��t�q�+�]#SUp��O��Q�%�?f%�%
�u�m�u��k��Wu����R�Ut�W72�a�N�2�,���N5}:����R�	X��������vTc:�!���C���3]��B_6U�SOId;�����MT0��F��d�nCGn^A���(]�oOEک�(tˤve���󌁦.�@��*,Y"��zv�[!6�o"t6�/���p�O�cAf��&yWl�ՠ�8'GKx�XZ�Ca���nIzk��Ԛ�����qT�v4��]�ߙTc�)�r`'A�:W4�2y�c��h�^maV𖠦�&i푊R��l�6��/n�T�Z��%ݙ\��h
xΦy%�ܵ�V�8P�(��Յ��Y�%RQ���sz�Qv�lj��"��Ȅ�F�n��"�b{B���U��cEW����rl�vf)�j2���������2Π�]����lɷh���GvZ�Q���D$��SC2Jƣ�J�j�'���+-�.��p:z��,��S�[rA���8x��u���Ѳ1��6�sr�L���jqۗ�i����ԧs5�SPD*�vv�	��i���R�/Y����ڿ��Nc��p����pOT��y���2�ш���{��[]Cu���t��r����4U�����O-�r�j�k�1Y��S��g�m�9���T�)�hL��z+���ed�;�22��@�ߠF�e���&�]f�7�c���+mNۋ�v��6}#��� ��5�;T���������]@�mX���]u��^+ŽAt�/k��6݉2%[��Y�<�q�ͥSY�2��u�R�r��=���]D4�a0��]�Xŕw&h��S6�nY:���@s2oQS�d"���/'bnt���R�`�9�A��׀Kg��,�r�4��m��\w��4&���1n�;���Y%a��;���K�l�d��������kaST����ˣ�i�b�Bo�
"��*��Y`.��c���PX�Z� }p�ʔ�;8��\2�zZ]F�L��1��v�����nv�Q�8�rx��}�Uܶ��*=���C��g��ņ&<�mɢ�Tco.�c?���_hz�9{&ʊ�x�_'�#��?���&�������n�ʊ�n�٨H��NdCl�㨃C��:9�M��@�1	]��t�[h;�4�J���b���|/�چ̔BL��}���H�{M�]��Ό����V�0+��.�Ɯ4+�x��dQ�c�]7���or<�3�v�����-�s�1�B,Z7i&
�!G4vcݬ\��t��^�[�ZXRJƚfq��[+��������h����2qY0վ���c��
U1���ό��8�S�cΌ=ϒ����u��c�-H�\�i��50�e�^���;�O,jU�&ep�Y�1�q�eNAk�[��,i����Ɔ�:0b	��!��7m�4�"�n�6��{gerV���Vc��C��(e7�S��q�x�9w��	�`ʕ��t�~c���U�}���D(=��+*6F)��K�m�n'̹]})��㾥� 8�n�V�Ͷ�y3->�9v���+�2�ّ%�GY2���u�ݜ�D��m�8�a�V�Zx�i�;�D=���-rTzҳ����5��)�NV��ܽh��D:�5W҂���2GJ�r��h��n�-�9J���TU�m���du��\����;J�f��{go�3�PO����>�gl�� ��Vq����b��L��O+����:�ڭC��C�����"�{Q�wG�Ek�;[�ˌˢZhJ��>��V�o-�9R�Tl�w�ev7�iK��	�A[�s�����4�Ҭ�]��B�������y�k�XR�Q.���b�H�g#�D(�M���8�֌�JwY����oc���ݏP7l	�ή��Na	Bt��h�ʖ�����U��ӏd�t��s�>�ͷ ��ʂ�p��zE�)ɔ�����Փr�disn�D���7^wf��Bn�-�]f�71�.!������H͊7���ɝ$�B(����+$P�7G�#�)��
�d6��b�Ȯ�:N��ge�:�!.p��|�d�F�e�n���c�䭏C}l���_a���D��Fql�N:��w@J�w�c�e�T��pAi��K4L�U����}n��I�x�۳����3B۱�}�; .b!W.��S�5�0w;�.w
���m�B��9|P�	u�^Cǜ'���fU$`�r�fj:Np�x�RUH�ui�fr��&EFtP�9EU�8�+���55:iUHVfhaպ��EJNe�*�!�JI�ns^.�R�UM��-,�����s�rL$ȲJJ9�Hb"QW�n%ʆ���:s+".Vu�""Rn�����Sj"jz���I-sH�UfRS��"n�8G�$�p�W�J�"��p8�V+5G<��qW�:$N�]\��L�D긳���P)		D΢U��&�$�Kj�,��BB��,�)VU�Tn�*�!��:�*%h�IҬ�Dʹ���F8ܩ�2兤Y,$;�ʴ���N\�e�I-:Q���fFċ�Zekj9\�8��D�! �KȒ�E �(����n�����S.���ugU��!0r�u�2� ��:��f�;��X�8�
�����+1�[u��-K�kO_��΄�t	DW��P�P#p�:�Q��3\%��u���GO{Qp�G����%��A��N"Ғ���7�~Goj�������V5yL3�k�����`O�1� O^�I�M�i�:I��h��t_С�U�K�+�h����[^�צ05�+�a�yS�[W<�p�p잟C�����H[>�j=�IR��x���T0ug��_e.�tX�{*#��,$��Mp�7Z������d9��Z��n�x�5��ݺ�D�덭w�w�l�s��M�����wEr�Ѓ�]l�6%.�?�����b����ش9�ɩy"J�i��L�p1�(2{}F�b��^G���|��5!��N%Bn �rT{��naT��'V�_��}3x6�����HfZ�L-�tW?CC�G���@��Z�u�]r�9��Y�R���V����jܜ&�3���zK�Ȇ�2KT�sb���Z�ԹNT��ݳ��5A����Mu��/�0X:V����L*�ƽ����֙^o��L{�z�U3o*��<9h*У��hr)l��#�����ۼ�Z����t�y(��HVJ���Pz\'�]��}�/ h�R�����l�t��A/�����R5��V��;S7mi���W9�i&�B��:厚���tZ�R�����7����t���%�wU��kd
|}P9�#CKT�D�Ei`)�Q4��w{�74���]�X�:��w!Fb�s�&u�Y�C��l7d�u�륦���ק��,�:��Qa��9A��9��� �팅 d�������dL��թQ��!�d�4,��0��y.w�m(��e�ybn$}�.P��">!� Eԛ���^W*p׀JJ%f�^�\S�OVNH�Y��8�l��֞-K�
;����-���p�a�C�6�u�2t�XZ*'��n���I��wA9�z ��!$�V�S��]>���v��S�<TU%�o���G7!iO0��u�q#{��x+A2j'*]pCܤhma�}MN�EfB��=.�p���d�ϒ�v6�����Y���S�8�wf��z%h�{�v����9�+�_�k��UЁ�$f��37�s�s:�(�e�ϋ���"��x��{8>���{[V�^%w)��[��(Q���KI���Fb�B@)0�xLfP�Õ�>�� ,e����k�D�i��Wbݦ��+92x>[\��AL����Fߟuk����1�{�`�\�0�.���k3��9��oױ[k�"����.���Z�D�u�4Ձ3:s���}\.+�ʽ����g+@�)ؒ԰���c�vl���"��0tӆM�����5�"��g6�R��LtF�,� +|�f�Ho<�h�No���m6�y󕁑/δ+���u|�4���T����T죱��5B�d�oRQ;SBw_�>�w�O��˩H�{�j;��(M���X�5�
S6��{s����T��f�t�,ʤ�*.j�x��eڝb%�0�����Yt��${��٨�k��v :A�r5�7�P��+.)�<zf�>�t�g�hC `�#�`���^I��棰ky���}�e�P��	��nť>*Kw�B�3k�ȼ���3�����D���V���ǭ��7� �*�O[�SW�<��C��G��n�]��R"�������%[ې�᭠v$S�K �n��T9�QS�ӄ��$&5���(��]�\�wF��µн+S�"�{�E�����{�G\&q�lA�r��'�U��+�C�BE*�]�/X��y�,u.�/IU�h����"�K���	'b���#�J�ظ�x(�����sޫ@��(m'�hSF�6�%���JO���[�j_�ei���@e��n=�+���Wl-��eowN��
m�K<1vfK�K�B�m�T�ű�V���XӼ��,¶��4�yD$��n;��i��
���%R1^rp>A���݀u4����qZ�J-w���<����0�Ԫ��9�))���bUS��s [U�qH�b"��/J���p�>�XO1��X���됺�w½���~B��u]�nc>��X��z�#m���U�䣧$ho�H*�j�/��b�X���U�/�t����<{9�ר�܅�J�E>\��^��ˏv)��
���;,#8��B�`���Y���	�|.�o�C5�-���)!-y1E���kY�j��٨��0�|.���K�!O�=����y+��M뼇�V��0��xS�E�#~�i��Fc{>o9��8|�	d�u�����5��� o�Sfn$!����S�a�w���}2�])��`�[�-h�"-Uw#��s�65�#�D�:"(Q�9THɻ�g2`�Ko:u��s��ľ��S|��tޒ��%7~�]�.�H2�(�.Il'��b��Yln���]�����BB;��/�J���i�zL|���"�U��Z�O�� 6.��V	w�s+�G�*A6#��u�)U��7�����O"�+�����~Yu{� \�@��`e9Z�=~߭Tү�]��������n��{���LvS�N��]�V���p���b��d�}�>���m�]��xo����m��7+�j�u��_pp�/d��i�;�v�[/��Z�Y'���g	׳+�������2.y>)�@��N�"%.���&�\ �I����h��^hɆ�qQב�+����B�Uo�P�� ots���A��.�����K�4f�}u�w5����bڹϞ�=��9y�?rFܩQ���ȝ`,b��V�)�v8n�y�y���<.�yн���pu�����M�x��.\�t$����s%���ኲ��͘��W�]��u�j�[Bϱӥ��9R�xEd��N�}�����hF�w�m4�����{KWBfz\=�;�C��c�~
�x�`�г����j܌z�J���v�O�0jl�����.��m�ԧ�߰mp7�9��!9,�\+B�6�m�_sV�1��Z�B�ɾ-e.*+)��T��8��
��I��-�鐶nZ�BJ�֤*xnF���"��}�\Q�Sn.�����z���s[w�v��ӭ`�w��a�(V���!�ڵH�kgj~⽚�L�S�n�}�xZ6������ �.�s�ry���N�b���5�{���5��=���`KF���Ҳ��n񗹾��a�ƌ��ӈ��z���7R)�w����un�n"�W�H���7��=°�d����ۀ���zYpAۙ�X��aF^T���w-�	Z�4f��l^���:iD;�s��C%Z=~��s�kDM��m� ���`���N�d���L�)1g/
��XX99F��c��Z�q�>ja��|��g(�{���Qhh+Tm��Fs��ٽ�^����|��C�=V��ڐ:�o!/�8�Qg$):RV���f�d]R�/]�Fe=5��rG7ܔU���ѳsVJ�F����Þ��#��7ǬN��	�
��ȍ�Ht���V��$}�>��5㿪�ӓ;9�\�!�P�9�:!�)�q7A���/ֽG#~���W\��
{�5\k�~Y�LJ�wF��v���~���z�u�|�(�x_
q���������^�Z�9��� �ld)�c]QYλ]�Ww�����jkn��бb��ǯ_OI+i\�®���ͬ?P��L��@B�b,�Or@̇�\�il���&\�jN������̇�[�4p���V֮'�@��~�=%��=.���j����fo*��ϓULb����6�d�uS�E�8BS���nU=t�]ԤtYz�!M�z��V$4�oqW�J��1��q4���(v����$D˼J�{ط��=�'���2�A�]��ib{љ���_t݆�
U8vQ3�S��7۪����e-mqɥG�1;�U�ln����s���b�����Hi9:��#�#C�}��6��sR77�-�ܔO>^�T+���#]�F�䥗y��"^~�-�}��W:6n;�#x)s�.\�K�rw$B�w���y�����b�xt���V����N�]k���2��� Cj<��#p�)��uL�u�V�vX���vuj�#OȾRWn�CԼ�ƻt�������S�(�M�%�$߆V䢞zs��S���o%��S{�8��z�ޅ�k�.����D� �2p?P�i�E��0�D4��ȡ5��}J�R�brt��ǟ9Y��� זI��tz���%ړ�o�/�$�[p�+j�*�Mo���yۑ��%��>o'���o���+������.�����=�^�rH|
�LS���k�����]���.�c�Y�
�>�۪��y��I���{xAX=�<��;H��$d��=3s�����5�Ѝf���i�Տpb���l�(\;뎐��{r�Lh'u�TQ�[U�=�6�n���h�J��fł}OU=}�Q.P�FbG#�ϯ��*�vf��t��z��Vt7>t6�p���ΆA�8�p&��hZ
�9���j�<�Z92l8f ��q�k:GZ(9M[�f��/
�n}�̹-ޭ�Q�jZT�'et�[�9�nmu��]y&sOdM�pq�����q)�`����Ik�{'P~<|�[�eM������Z��mڈ���M��U�}��Hn��󮽑���	�rBz�[�T=�>H����iT��9l��&JR7���62"xȎH۠[�3q�k�!}3p�p�O
P\k����$t�wD��l�c��557����4�gȻ�"�E��x������(Z�M$�jY0''�,T7��7���l-������
/�{�)ϊy�0��Ta�s E��׀��{S�E�ӅL�O�n]H�t�7;P�DM����/]�l����}�xU�9��q�q�����V��-U:+\Et�w�!��*a�q�c|l����B5�'B`�r/�IL���X�"�fQ�K�cۊ�U~���϶XF`c�S��+��`�x�,��JtO)�5j��ۤ�r������r�Ѕr��ώCW�}v#d�0a��N���-�]u)�:�=%_S��aN|/�Q��ԦTuC�Hs
C�v�[tf7��BG��h�N�)�FV��*:4J�J!RI���6���?�$�Bѱ�:n+�p�-��>Yڍ?s���A���|+h���&+��k}-,b���f)I��ǹlˠX�s[�3}W��Ǣ:/����J뵦�7O+ͳ�����Q��ֽ:��O=C:��cw�Tf/�r��ur�O;�el�s��;�w�F��X�x�Z�6l��㒭 '%�]�(-����yf�RB�@�g2`�Ko:w�f�Αs
�d���d�%�%"��������99@�!��������qٹwK���� G����XP^�=o2{U��=ڏ���#��zkB_7�?�d�@j#���AR	��ri~Uj�E�5 Ŷ�{�8VE�	
���	�x�	܇V�u\�"�m�]/2KUה�'���/Y	�IVj�_�R�Ɛ����+yܼf�j�lQ7��o�:��L��ʢ����y*���__���ɩ���Oo�S�����ir�]5�����0~�M<7m5�=<��W,~��+=<&�Ϧ���.��e""��R�\��\$���\uN�a
rr�1�iF%2u���4���2��+�DEG����u��:�K��G�S�`L0Vt� �]��i)��#�d��t�x�(tv.��������X��g��!�/u�"�j;,��MR��ǒvEW
���늺4q̀��[�ool�sJù�oH��0M�웧��Z>��S���1PD�i������Wi�6]s�l!���o�8	 �Lvi���nBK�x�:�b�8�,͆l#Bq�0cY9���SNىis�M��Տv[����Y�@z˨P�-��ubYf�V�F��?pUs=�>��jW��e�W�Ҝ|�� ��4��Ӌ>�Z�R��|��t�[7�G�	*TZ�#g).ىp�k-O�D�<u�����IȺ�\��֦s��r��k!�l}N������ְ��p�PWr�k4����p蕛ߊ�
�n��<6_ <��������y|:�˼u4M	�(X��$�S��Q�����jr8���E}as�����ت��CX�c���$�f��3uV��nadW���X�[-��k�0�wŕ��T�{J�]@�gѳ���r7����9yМK6�GL9x��Bb3�jܝ���9I�i}��&4�
���ʚ�c���(�C�D\�88a��\"����i�0W�/�5� �X:Um<�EL0�h�ù����).��*�Eg�Sc�]w�;u�t���Z����?m��0�=���q���ծ��L��,=�#��4WBEķܤ������FW��|�89��vH�}�ih�۪13�g�O�4�G4=����)�6
Q�*�`ϖ��S+s�v���ܮ�Ƽ��J��|�%[g���1�@�D��H���T[�7��Gc"(�"y��u�i�s��s�$�P�.��x�^ż���.��vkC�������.oXÜSJ�m�[\n&��r\�Q��6�IV\r�ߥ�go�9eC��T"�h��כ�ɝ�JyF���؋�2���>��=yKU
_5�Cp��Մ�@���`��i���[*�\���J�I��R��Rі���XzB�m6�`�wr�l<%B��5�҆${z��T5��?�IZ�LV�t� ����]�j^�W�']q�}{c*?���9E���r�!!}N�:��X\�U�"���)譵���U=_����L��]jS�CD���t���[;tJ&��s����W}��ܦ�2)ԏ�r�%y�1� 2`�Y�J쩳r�r= R��M��ԬM1�"�3>���Hl���M*�5�Y�֮kb��9B��]s�
؟b��E�P$�3ZA�x��ymM����v`)*oI�ͫ��i�ՙ�C����%
��Dm�hQ	m��T�#lY{ג���\dv�
�V ӭLt&�m������$��z��1�uL��+9>w����du֑��W����Gv.�C�dW��!2�q<ي�4R���{`�Q�&��ׂL� 0�^������Ԉg�zu2�	|w74�-�����؆�9O�n������c���\6<"�̱n�"x�u��*R��+��sX��Md������|6�9-;Ε�5�\��n���/Aqe��s(�k�������z�;��Q�LJ�Aah��^S�l1Ǒ]W�.���y݉�_7r�W���E��"���1�m#.�AERNb�*m
�+pڐ5#(�N�[����T�K�6���n��y�6�
��u	�V��ۋ'd5;d��8�$�g;I��o3kX�YF�]�J��8_ou�k�s�WI�`�{{N���[�\}�)RJ+w�#�V蒭C��{���)v�����s���{�"tɠLFtX�����f�Z�N��T��0u�R�Ǯ���J�kGMm����Sh��åkXK��{��;m��ܢs!�)��1<)h���Ԃɔr-�qd�v�J��������(n�Yq�hN`{�Eí�u�j�a��-!]ִc�*v�kO��96��d���I�Yk�S<�"7�������8>(:���|jf|��߳�tpdL[�.��u;�L�+a���˃�Xgj��Z�7|X�����M��#D�M��k�0,�knX��]8r��ة<�H�\��[��^W9�

��α�X�H�g�f-
�<oWqJ��Bun��Pu`�,��g �ثUH�H֍тv�2�;3]v	/4hKj�J+��Wsk� ʱ�Vȶ�Զ��(���*l�<��;�d:�A��	 W��L�Eg$���	���RDB���$����\d�Yg�Ô�"BH����+$�.hD��rb%��W(\��y�A&�9s��29]2L��4Ij�$P��٫���꘡t*���B��gB՝5a)"t��E)h�Q%#,,�h(�u�QE�pc�.�(Kd��a�ʍ"̒��e��"Q�VjQ�K3�I+eIR���"�h�C�JE�-!��\EiU)R�J��	QQ*")�N����	DᐒU�b'I.����+�eKU�&TZ�ќ�����\�� ��iHX��%F�p�(�#���Y�BDB̍4�,)X��j�q����5 �̺Jlˤ�sp�f��#�35Kia�it-4�K���mӭ-R�+� k/����7�f�ɺg���.���?tg �Oz�9މQ�D�FVc-�<3a8�l\Dm"��� 杽�gUlo5=n�Iv����w��g�͎��aT��E	<C��!V˧z���Q��ۉ���u����n�����O�ױ��`�0�G�o?|�t� }I;<�޶����>�����_�le��vVf��2}�C$�r^$z���n'=��{1۾�U�C���0���4o^9w����y�����#�:�����N&����x�|@���tG�$��<�|����1�Y-Z]��*��	�ɏ�H��9q�˓��v���z����z���s�ޡ:v�S��p7�N��;{�7Hq�!��@��������'��w���	> �k��$�dyJ @ȍX���j�Ue=�����_������
�V)w��N���{�o�|L*��|�t��N�<�^F�'�����ͽN�N$�����7HN�[�ݷ��#��g�� �jϽ� |NUſ��t���nl� �a�����z9{�|��{��~w��o���>�i�&��ǟ�����x��?y�G��q0��}뭔P�8���y�^�.���|<������C>J>����Q���^���]Ƞ�����,t�N���I�ʐ$8�	��<q�w��w�<v�x��i;?|�x�o�n'�8��'�o}#�v������}�޶���x���;W��w�������Uo=����V�?>��-C��!DY��t��8���7�q��~�t�U�8�?�?��a�>�I�����;9��;��忐���7��!:vU�D H��F����1h{�>�'�����~���۹<�,�Ғ��f"���.����۴��>�<��}qҸ~?��>'ht���w�q�C��8t�]����#�x�i�]��|C���I��\���N?�<�q:�{c�f2k<����y�V<����1`�:��t��x�M��s�i0��v��|<�x������c�w�i����}���Wn��&��x������ӼM����GN���~wø�;q��p����Ɩ�3~팻�ipK������(��!��ϼ���eӼ~\��O��N;w��;����7�w��aT���n{����}w�����n����;t��]��8o�t�ۉ�I�M�>���}�gL:�g=㶔i6��h�	��v־�yudͳ�o� +��"������.�*!#���Gw.�3W���y�R�i�zI��$���q�P{38��1r�q��鲫sVu�\�v�u�k�:�CΝ��զP�K����óV�6�$�G��o"�}�}O���8��:����:L/�{��Ѻx���>��ݦ�|~��v�]�X>oz��=q��7�q���z��<����>&?;�,�}C���ϨG�di����l��pp�������8��v��,;)�|@>������o�~|�m��n�w�:q��~��[x�w��bO~M��&<v��|�O�|� �:�ԸN5/u��d���?��aOuhI����<�ϱ����vr� x���G��q	>o�p��ߓ�>c����i���o���z?���@�/:������w�|���~�|����= �e���������S~���w�~Ou������P��'I��?u����n�=O��I��e�u���ݿ]��C�s����ny���ݦ~v��｛��4\��!�G�G��uUV��%%@{�Wv�8�y�7�v�]�<w�{&���v�s���F:M!?S���~F't�� �n>'H�t�Q�x����i0��G�A۾�\���8;���鏌�� �[�hs8���1|����};�v���z	�
��=�ݾ8�;޹���}O]����>�n�v�{z��o�N��펾F$�N�#��ۏ<��?9�t����|�q����1�ŃU���\���$R��t�O�����|�7��8������9��x�����	8�]����?u�;�t�=��&����$���u��8�}O��s�}Iĝ�n���q�����1S�_u������G��{h�TR�wHq0�|C�ާn�v�;���:wN���s!~���;���ۤ�;���1��z���k��㎝�q0�|�=O�8��y���S��y��D���~���ݖ��y���>s�?�q�ۉ��������z���0���瑾!���x~v�]��w��|ǉ�z���O�s
o��݇��t|L)�B~����'Σ�^{�ܭ�zN����i����f*��]���>��$��i��yӿ���������;\��n;��'���N��O�>]p���8�S����?�?�㏛��c� �/������> z���_뾷�n&�	�>�<�z��A�7���Z﷮ʉN��R��FW����^c���p���ᰫ��Z����+��O�+��Vd�n��cy�3�%V�k��`�':��z{�&�t�E���L3Jۘ��)b��m���@k+7dVrY-SȻ\���
��u�]&rq�#�^�}4��7�Ͽ��v��Q�N{�v�8�<~����v����iӎ�J��?��o��?�vW>F'~C�q>��}N��~wo�v�]�v�s�n����	��b�U-5;��"��) Wr(_�?���Ow��u��Rq��:�z�;q7�#�¾[}N~��F��i���������o��pv�v����7�\��w�I�wo�����������kf��F$í���Nk��}~8�����;�N���q�P�s� �]�P����v�}�����_Sq�ۉ�ww.��۟��`��
�����c~C�
=�n�W;_�=NLT���O�����z��#ݡ��Kt�=o��ݿ&�	�Ǵt�+�M��x�;t���M�z��m��:B���z�Q�>_{�.��T<����q޻\�;��v��O�-�$����}���}A�EL}�������s�v�{����)��4��hq����$��x�� ~Iݸ�G:��n&�	��������>�������#_}�;w�i����]�\.���������Ǯ%w���>���Ǧ*b�� �Ù���^x��}�������ON]!����aO_�|wN��!�C�+�	7׭�)��ޡ�8�v�ĝ���I����WHq0��o���>&���_׾ǽ�}��G��t�-	2-	_X�9Y_\g>���=ĝ��:wn�����n!~����y�\
o]������:������qߓ�����q��>;�]&vQNQ�~C�������>&����]�T���~��K�4��X�o퟿~{���
���_�mߑ���o����q]������q$��������ݦ�	���:W�ϣݸ��`��t�ڭ�'I�	�;TC��#ʳ�;�j"����k�3>�3B�ď^ ��{��MH�G�F�'���z7��0����׽c���q�Gަ��?����9�~��=��� q';�uݼv�n����r�5�����^�>�&�G�_�*k�����<8��i7��Ӆ��7�����qǎ%P
o���C�Ͽ�7��!��~��!�������޻�8����:W�N;<����a�o��
b��>�
�b��)��K=�5���x����F;�7|�uf���md��x��i�T|����UA�p�b��i�Zz��l�0N��n�[J�<��(5�7v�wC,f��u:��$�����u;�5����Ȑ��-u�e΂��ūP�%�,�++[M�Zq<���	�5��{j[��r��_�բ�1��w����
�c����n! q/o�'N���|��'c������s��7�^�{��Ҹ���ϼ�7�_�z{�=M����q���bw�S�8���J�#����%��J%��D���L��T'�v�z�~��t��I��Aw����c�~����>�^��;���u�~v⻧|߿p;@�$��翼���&�	��ͺN+�B��y�u�z�L��w ��v��w�Sӳ��1Z>�ު��~v�oϯ�����j���׷.㴨u��y�8�vV�Q��'�����N���~q�}C�8���9��ަ��:O��x|L>A&_�>�\�v��0y}�֔Vz��s~�������N�M�����k�@�ۉ�BI�������n��!������t��q7����j��'��w��M�������=wh}C�q����U1��sJ&7�����?����Oޘ�O�?l�s���ю���'|�n��0������|O��n }�ގ�N$��ۏ��s�&��g�8��7�$�7�9����t���9($;~t��ۉ�B���[�U�{�:�ΟqX������1���7�/��w�;�z���w��}��:>����^���4>c�C�����E�F�PV�т����t��6ȉ��U���3�O�˪��sݰ�i��s�c�w��wu�"�$N�J�u[,�3�L���TC���ݑ
~����_�r��8��|lO�w��.�8C������ ��?r^��ߩ4q���$џm����l7rtD���[�N�v�h<W<�)U��.�\�_��u��������e�2�q&H��ѯi��4K')�5똅޻]�n�;���jؖ�細e))+�^��&�	�.������a��3k'��j*�2�e��öM3��z��;�Xh��T�X�:��OCl�KX37U�綕��=�����9��mR�=�AgD�q�\����d}4sr�F�%(>�̃�%���^��LA���,pm��KOLip��J-�uΩ�k9����9P\E�h����*jkQX�֨0�؉�=oNB��AD܂-�_q����|ը]���f���c�[�
l}����n������K�$9��?f�3�	�QU��v���n�(4�pЉ��&J��F<-��RqZ+���<���x�>�qpH��5n=M%J���~B%3��5i��d�������	�(*�i�a�|5Y�|�J@Œ�R�c����Y2:zC���0n�V�a��B�[��6+ ��a�+����_\�٨�	�0td5Ź�3��lʪT+ >��?Py�[f��"d����Ҥ{$�1�75=�l6i�����M����6�d��ws ��C�-sŏl��b��;��������8�}���A\@���Ҟa�ξ`\c�9;�Mf_s=(�D��RSC�!�)����Q���p�?=�[�,��X��H|��Oby3)��ئ�bI�X2�yn���s0EB͛�@�/�e��xۧs��<"����˾e���ԓ(����w9[4��W��X����9F3j6�9Sq��1��  �c�OkJS��/��α2;�+M���u��+�Z�r�կ�nwV?������y�p��dύ���J��U�7 5�9��Y!T�s䅊���A6X����0Ͻ��_FՆ����F�_r�[���T�F����cf{;��:�C�L˄����P�Lb�ĕ�������\���Ҁ��ū�j�@��]�gx�z����<��cR�Y!��J��cϜ����k!Mƚ�9�v *���s�/ݚ��� �f���5ITdw4"�;�dO;r1�KCa0U����oTa�v������Ʋ�*`��~D ���x4��nc\n��9�E㟱�v�vD��&�����2�$�Xu$,�E�
�\M˚!��
S5 �'��G����78����.���)��o>gx��U�s�8f�����ѯX�Z� ��Ƃ��Z@�峞��������F�-l~ֽ]�i�K���I#]D�[�SH �H��"���W�N�woE#�UFq@��6JR��&cx鯜$�!�����F|��3��`R�4��d�ŕ�"Z��Z���t��C)���Z���3����J=j����A�;��^�q��IP>�+��2�*|0i�Ӻ��7\t=o�n�x1Eo��v�vQ�*�v_[)Ӆ٤q�������[4�I�HEnF�h�,�&�7Q��ܼ�'Y}|��;u��W�C�.�M��D�i1�tX��"���$q�lA�+�U��!}3j�"��2�8�j�Oٌ;��7A�Mf��P �N�rxFK�GȻ��Ⱥp�x(bu���٨f㺏q6��S7�f�^:N�/�@��WڪQr�2낌���=���U9V�p��r�=��C������ K�y`������N���n����yf�\+ۓo�)M򚁻���]���6�g��ƧR��9�.#�t��ՊP�1P,o�����_����}��E�.J(B��B!�a�;(z�}�^sTq�G�k�!���T�Mh}��j�b]�f���q�}�B����h����3�%~�+����y�!>���Ve�K/�0��"ޏ��;�a��KF:	}�乜�~cڰu)���b�*,9�0�.���x�Nѱ�E��w�؃�t��/O�T<-��N>c�e	�c�����<�)E����!u�E6M,)*H.͓�T�7*��	��� '������ ��^݊�y�J�(���D^l� �ʴ;^�,���(�ʻ=�;�{Z�������m恞孥�D����h9�r�k;���e��H�}�����$��21�kw��-4�̊���jEΆL!Y��v����vg"y;r�J�=
 s��c4������嘉F��j�^�3P�rX���τ�vrL��=�Z��	� b���k��e��k����^E`q7�_����#�R���5�9/�|'^��:��TU;�8s&yV��t����\I�U��"'�>Y�F�8���2%���Ы�U"c��r�q��<��o�B,%�^���]K�a�.�}P�l}9��N�6nw�6Z��h�ҭBt�d/��
��~��5@�W9��p��)�ϝ��#�T린1=W��6@�8XՍv.i(����U��t�i\��	V��٬�<��]������Q�[q'�W�$�8:l��W}����FJ�GiX]P!�R���\��^<u)���ө������ᝄ����eͷNg�ؕד�C��4����BCRM�����__���Ӳ��E*���)���:o;.BM�3;�Yp��U�K��5´f<|+���	X5��Iw3e�n�ܺ��e��9l�G�γ8
���q|�,�#\��<�������h�/Yj�P<m�]I��qíΗǅv��d*�2��P����ǋ4����'�ᦫ�9��M��{w�G=[a�X]j t�x$��-w/������"2-s�#[���'u[ۆ��D��n_(kR{�U�W�uI��ҕ
B���F�������]m��"h���S7��Ý�k!�lS�`�*U�<3q)���[my{_�j�8�����e
��
�;P�+�A�l�6=#�^in	��^2w�H^�}.+��i���O"�>�`߀n|3�B����l�����-�-��L��&~q+M	����Q�N`��f\�����캝̤ �$��)_ئ�N7[̓���a��#����~�����r�|�!1M[���[� V���
��U���ݞ���rh
�U~���^[j�\x0�oc#a�26za�=7
H��5��)<�4�9r������@� �r�+>�I�Uk;��93��%��ا9�"_]�\��h�VQUW?k�]0᥊FNdy2W�!���o;]ާ�o:3�]��<�|F�.o�-4��3���cd�l�3[�dM1�B(��;��f?F�ܧ~]�1�U���m�um���J*�ge�w,S����K�7}3�ELKvG�	�')u�
���mm^�3�AV��y�E�Bh���]kϓǮ`�9R��;�gg���ۀ�y;c��#�ve�non�Ů
6) �s�r�3��:e���݁��������wv��,�n�Z���]���Am�᝱L�ϓ�����t�p�Y�QK��}��
�%@�#/��|��7�\0-�fC؆-�ɕ1�;
�P�4���Lc��HP�\�á�c�(�J��t�M�%���L����5bo&��̗���ȋ ِ蹜Y3�E�\q�9��P��֯n`|>��c��ҸZ9�Jy�F�:��q��H�jHg욖�s!�Ҧsx4;EhϘ���`BN�C�Q���i	�zzU�u�d]弁|Y�i���'�Z�$F�����FNķ*ΥU�O�R��V����T�˻o���x�X���������7e�ϋ���ɿ�72�p��X@j����&a�kF�JY��\.����Y�,Y%���(��J|�س~�!wZ�����,h� �2p����]�w�7����r(���j�yQN%d�,�*,3я>r�2#{>k!M����M�zp՚���9���T	�Uc�KF����Uu��#O���t'���u�э�al[y�6�Bq���z���䇸K��+�FK���K�f��`�U �EM$^9��ju��(ھ��)�^��N�e�n�Ѩ�H��(� DK��z��Yq���C]h��c��w���wj��ݷ����6X'��fڶ���&���l$�޵�ێ$��,��LN�j�=.0�f���_� f���;����a5_�:�����}��}9�F4���N��<�SwCk�$mgU;�8�
jpvZc�2/�#�f�)W7��E6՜jo ��oL%��R�(��L�	�M�R�
�mfA��ao�M��ؼ��wu��1�m�,���k�|�j;�i��AA»L�CZ������]W}}H[x��
ZV(iq����ܒ>tU���*wˬ��Mtkq0�p/9nI��oTS�2�4d:j�C6��̺��a2+-[.��+�.��E�^DT:.]̬�NW�AC�h̝Dd������Jrs/Μ( ����)�Vӳ-7�C)n�ݵe`k2�0@7��@��s��;}F�dZ�Eӧp\½�P\Y���ki��؍�|BO..�8d�lb.�_5�e��\2�W
ύ楸�˚*E�*�����C8@�S���V*���nM�RjK]孮�-�GNm;��ُ�*I;Xz���s���w!�e�-F�ݹ��7��>�Aa�u�D��;�����=�9Ý�yw��ZanLl��e���0E`vgCٽ@m�����*;�����urK����Ϯ��ԝDq���4�ȝ��z/nvh;`;}Ί':-98�f��O0�(�)�����mVt�����g�NU��JY������yM�7����ed@�Û�etSzK^�����*��uKd 5ѵt�}��L��v"_su���C����X�WrӋ.j��б��
?��x�p}CE�]�P���$�ӡ�:�\�@�K�%�*R�v�&ջ�
4^�5��;^�Hí�MI��w�������__R岞��=f�a����X�R����2��+�ׁ�M�-��������3۸,�u]t��eF�6���w��l=�J�а��5�%��F:r���ܽU)��%Fc��۲≫�c4͕�d�����sQŢ5ocJAal�#��1�te�K�94�a���x*��:��U۷Eg=����j�@,g��I7��n�B���@��L�k��3����y�۸��s���Ib��{9�[I��6�l�w5��8,��c4'�m*��uY�SR�p[E�ݧ&.:����ʵ���i�OMHΛ)� �aۍ�7.�R��6c����j���jP�N�ʶ� �������βF���1Q�@�z6���\Ch3y�>�O:��#
ރ���y�;S���nx�d�P�/T�D��MU����$e+ͻ��6vkq�:"��p6i|�`犢�g�t���
��έ��ҟ<U���Z�ĳ���ѨU�f
8�Nt��I����E��wy���y�^��8z=JG���0Q�@�|�Q�S.��huJ�+$�T�B��"�eD�K�����Bڅ�&,3W�4�ԱM5,�0�V���ই6Z�s���ƫi���,�	M�I�4�E$�0�DSiih�FQ��Q%����N��iZ*(��npi�+��S���)t˒]Q!RA-i)�٨�Dh����M��4Ū���"�Q��J��%��S���T�0ّ9H��.�H���"!$JR�l�p�S�L�.T�YF��u���ZZ�D4(�"�$�Ie�T��$$R3��&"V��\��QH�ƪDePiV���T�I:T��j�Q�+(V��e�TBI$�	K�E�kR�(����D�b5IC�]ŤI̔Z�%Q�YRaJm��;���,�A�"��ht�L��CCjE����Φ�9�M�"�H��L�(6t�uJ5��4(�"��.J���ӡI-D�f�����q8�Y�*ґ��W9�8��Ȗ����*�T��B��PF����=:ø�FveZ�PUl��Ӽs�	Yu��,u	�*�����P���x�dS�P���J���yl�2���_�#��!f�Қ}�MD��|I��I֠db�@OI1#iř�qM��70\͎�1���������G��3P�JU��0�P66�KP�fy0�e*�6D����N���ݳ�I\� ��$��{��h}q{Ng��i/��1yZ��T\A2�T��&n�mM�2ʕ'I&o9bX�Nu�z�v~2x�:����U�⊝�&y�	��������:�W�bPu��{80"d}+��45`b{�|o
w'��C��N��5GL��P�F��K�n�����%�(P��c�$1jL`RxA!h0��.Y���Oh�<����QiN#��uJx�
9���K,���Є��i���������׋%g)OE�[��#�v�TC�!�x�g�`��[@���n'jɮ��cpl�0��O8�7����IC2�����uN`Ƨr�-��z�������7���U�5��Жc�'��w8��`�}M��Îbe�	_Ȍ�����2�Q+W��J,.�.�ę�'��:R��b��]*,w��J&�Y�k�'k�{y�4��oyצ��3jƳ��=Wt�����8��7�T�=M��\��|犹����-Tެ�yHm�ƹm��%��:�����о�[P�5����n�{�r���������%L��j�[=[Uâ�@!�:�+��0��k�q����F˗�)��E��5�)��2^�No�/��.g�_1�B�G^껖��FŻL*ͭ����rm5��F	���	��PG���U�-."���6�y1�g��OEzR�懯��ss}�½"�n+�{i:� ʇ�$]/o&1�{G1��d���Rn����%�.e�mv�:���Vt�3P�_P��ϟ��g$kZ��O��4�@SGw�Wᶼ�bΑ��ndR6���T���j�.����Z����,�j {Vr˕�wV�·�1�:Z&�\�FL[Py����5cY�)�F|����7B`�E��2ԁԼW�L�G��:�ѫ��yY�~�bxK�PR`�L�}P�[�7����6`S��]���5�t�QO�/�t��҇���|����	��9��p��/>tg�Hە6t�۸hbފ4�=����g����0) �3��A<�	����fF��xA��t�<pJc5�y9'�r*f��k�t��N��G��kF��v��T.b_�-W�;�d��o,0JFe_F���5&�ةSs/PҜ�1Q������5�/����#�_A���M��l���l�K���ۧ�3ei���sT��;�6���}s�ꪯ���'oQeD�	3�#�X��l�S�/f��;ʈ������B=j�v� ���
���2��$��
n�7��-��5WAhs2��t3��r^��4�1?.�Qua��bI:[��b��<��;�ó��H*e
ջ͇Sy�];�����T^�KROإwe�S���Y1�®���򸬵;�r� �!0����h�����"�����⥤�Vb��Ѧ�YT.�!PӬӣ�U�&�`i�S'9��;N�C�V��R�x�+�q���ұ�Am^Ok
�۷�JQ��b���N�/���pa��U/D�9�|Vo$��5�_���x>���!�Ȼ���6�x	6�}���
Ú# ��U'����mƴ���C������y��[*��+�y��ܥ��!�k�0��w�\����N�^�}Եr'�(F1s%�k�d-�����/_\&!E5nN�[}'>��E	�R�2�O#�s��d��	/�W|�ByV�v�9ώT-74�����q;0�V�֎�ת�b�?l�XUu��s�aR?;�50�ʍ�Rz���Y�v<[8_���z�w��ᘫn���1�e�SZNP��\Ů'�r�������=;F��§�[.��g�-�z�?�&��g���G#�n��R��T`Mݷ��FƩF�x������G�ٹ�B�l�(��⤫P8"p����9:��􍸋����p�ɝ�K�$o��yv�'�(ĭY������6<a�P0"s
&����K}�N+E:��E���(j�姙=�ZH��7����25��F�y�@�~�A݀��yѐ��0��U�����[·���pZ}Mm]�4�X�];@F1,M�L�w�A�HX-����yYE��l�>�^����e"�9L���*�p۳!��2 �5�*���q?��^���<��aTJ������ճ{.Jc	�F$�>�M\	��j�y9wsbm�)��4��[�j�����P�uG
cE�5�~������Ҹ_���-)�����+�G�մ�sQՑ#���^
�E�A�vѨ;z�XM9��Ύ"���WH�҉z/�㋚*lQ�<jxF����y��������ްd5��u� p���xz��˙�ӽ��f�g����ֱ[�b3���xk&��̺����\̣�_{�ɹ�'�U�&��r�u��8���}���=�����L�a`�Z�w.�R��o�LY� /<eY;��eKr�c�yw��h��՘��ߧh��oU�Z��֖9u0TgT�}[�J<�W�n�c�*2��n��gt��fZY���u�O����2�xflW^�݌?y7t�6��>��{�*@.]ت���k�.���,���+gE7&�.�V�p���YՊ��
��@�9v\���σ"7��R���UWD��n'+�WU��]5'��H4��J��7�Č���Z�,�v�c�����0��1�z����_),��<=^
�x�.�9�7Tl��wn��YQsW�s�5V��q]�l3Γ�IWM^��\6�;):���0��RzKf$`[c1g]E=�;�]��ø�:�)ʫ��n��O��j�H�J=��6A��A��i�	_ �iyѓ3�4&p�Q�k%@��xؿ�������o �B��Gt7jI7�Tu��'�$y:� 4]H�q��)�Ϲ,�n�F|�s��izk䓴�f
u�M�ȇY0!ʍ�v��0ԎP�IT�a���@2"Jb��#����O�	t2�3s�U�6`��ү�k8��l�}����Ƅ*��^��R�^:�����ip�]�y�t � 
��37wK��/&B��pT��ݪת�m�l�
��w�$6J�Rrx�vY��w��t��m=�4�C_qS^L��}�ѻ��y�^
cw��!��1]���ˡ-9K�n,Ю�O�iJ%��^��u�8�v����KFᮻ1w'��� /sj��;a��í�z5�-���K�P=c܁Fj6:�P�R�{�M��R�(��<�s-�I+�K�NeL&%��́p�l���p`q���$>_g��%ϗ�aQ 6�_��nBTR����X�f�9脮�ƧR�NX8Uw��U����b�7Ŋ��fAߟ_�Y/ݛ����/,�e]AP:=I��Îv$K�.���.d~}�qe@��<�H���2��ʹl���Eb�P�91Q�(y�j�l2��0�1�s��|Woo+Vs,�r�Ww9�<��G�39�*49�5_=Cg~�j�߇R�Y=p�-*,9)'tls��;.r��y��
\��\�W��^���t<3旅8��s��ք��ۍv����[�*�L���f	�_[�-h�".ۤ20D�+�xo������S/w�%M&;{0��i�J&���6�2`��a��s�����u��g$-b�Z��O¯0�ͼ���w�/ts^�~�����۵��}ιs��#�S��>Ȑ����'g��?IU1_�*~�`ɹ{2[�eY�]�&��-��c�]�@3���c]y���m�7c�>���i]�Յp�M����4K�ؗG�z�c�f>n3oPk���r�)qE�{�40��d��2��f�� ��fi��;'R��+h����6Z�L�����_d���s�� /�#�/�*��C]Ǯ^O�ȼ�!N����J��Ǔ�E��$��ՕEӢ�	&t'N��RW���)0�7�#���̝�o�#z�����`�#����h�ԒQr�VMT������#��_s��wژ��o�xL��=u�肤�mqɇ*xvv�-% ���*K3�b%��U˝'�r2�%[�p�F"��v�S)���u�G�[�(QS�8%NC��7v9.�O�Πc�N��ũ\��X�.t���ڬ��Y]���9�8yPg�"7�����r����C��7ә��W^NK���`�l���ľM�ؼ\���p~(�6��c�*�2���c��J�� =e�oF�D�o��7��Z�ҕ���ŀ���K�a͹�9h�F�Li���z#q|�wq�vC�"���;�ч���`���5Ƹz�K��R���^�ۋ�Y�l9�[=�2����Sζ�rBƪ��/{�y1�>�=�O$W��$_��i�N�,�@xj���'�~�M8*���N�u���qa��Ӄ�Ҭ+�*��5���b'黶�"�d��^�f�L�b���[鳉�uQ��D!I�f����NK6S�v"x���\uf�s��(��xos(&�L�"�_,�x�''p�����&t:�"�š?W�W�����.s��
��zg
�[O>����*�4r}fr8��,϶�WR����$��]�Nr���+6zÇ�s<��O�8�	�;\��v�s�->����j�t�8|W9+�2�����ZhH����0�B�d-�K��g���}������'b��Jt�l:/D�<{�7cYS�8�� �(���t��^���W'���6��#bza�OL^v��<�=)��Q�4�Jit���Q��/�i,�����|÷_Q�NL�o*/i��y���s;JL{�LM�����R�����h���<+�"�%��%qZ(�y�<�π�36s�#��w��,b�����;�1)�����A�#vv�TQvl8�U n��$JR2:o[Q���I�2�;@FC�������|��U�A��!m&6T7��;]䄙�J�	q\oldC�L؄��6ʛ��*�6��{�1nfL�!3J�P�=m�T��gh��6�.��욠�U_#�;@ߠDm7����~ڞ����<��̗/\�=��#���*��R��4W���S�1Bm��&(m=<08x�9+"��~ޠ-�(�ܨE���$w��F���up�(U��ܓ^c\7��u�I��W�����|�Sp�`ݮBη�r�9�8�ۃ,'�)�]���o�u�>~�]]����k��������]ړ.�*dd��"�G�Fb�9|�a�E��������t��7���Ӟ5P��n���ҕ���ok�Gw(��3l�զ��f�e�9|k������ԥč�P�A���H�o�4��!��^�R�;�i��������W���e}�@��j�
c���<[ޞ~K��da��y���J�Z�7\�/���C�͟���;��[C*p{�J(��ݶM�O8'�Qگ�R�Sp*� ��)�}�T�\�3�I�߽w��Q�j���s��f�$���56��CTCC>N%d�,�*,3�cϜ�dFhe��5�ϥ��p���D�t��𻈓K�xy���i{U^�0�>�(�NAu��П�5����Z��E$����;��`�`���u~���Tl��v�b*k��toC�sj���e���~;=Fq��c�Y�µ���i�'A�,�C��U�QBk�k���H�{;�)
��#���ʠ�'���C�)W�YR�c`h��Q��(h=pv����q��DL�k[�+˭p,oI��w���Џ����hq��S)��� �j���8���_�����]�W��-_��v.���z�S�5B�q����ܾ��o*޼�N.�.��˾%ݚ�lL]C���(j^��'&�$���UUW�qz)nzt�����b�3.g"���2�S#L7jt���'���H�U�����^)NooQ #�����p�W��DEM/�Ρ'i�6�����3&��dv<`m{��M[��ј�TBh;�"d}-�1pn�<d&O�	t3��ÓO�֫[��D.8^�<�Qu�h_Hy_�hB��U��T�W���hV�y��/��K��Ku�N�)�!IKC��%5#y�}'`P�o�4����>F�{E��u�|��^>��$��]��=�(\	��>�Ȃ�eND�'��\JW�����*-�X)� ��0�zg(l�ݝo�����{r]F���a3�ﻛ��!⷗���*c[Yu���~����_OI�-q���b�j/qe]AP=���ǯ�')+����w�eh�6t�slnlJ�ۧt#�N�� %����訋E��#�"�:�CQa��F�z�ԛ�,��k��{����8�M��V��1���	}��E�ՕF.��u�J��S���[�Q�v�I_��;��4*�nu)w"(�wL�^���ڦ.��kZ���5x/&�B{�9ݑ%q�KU++v.����D��6�EM�YR�dfe�P���B$�CMo{5��I=��ɛ��39n������n���N�ᴐ�h�!wH���'���4�+lfwU�x�±�t�
���7H��)M��iPvX�qk�)V��6o��q�6by�U�МxI���㭘F�����ū
˚B�"H�Nc�/�1�zo
:X"1����\��4�!��݉���Ю�9�u��X,�O��VV%�p��+	��hD+��[tm��A��U.m�5���
����R:���D[
���i����E6E��}��0B���Ԗ�nϤ�s����C{�X�q�U��.+�>��9z �ɓ&�ǹлS�Y4�K� �8RB��v��.��CJCE�'�B|n�P��=�/iK̍�b�c�Y}@�-���d]�(p�仦�P����v[3��11�IclR)]��
���F�;�;��gF��6��L	Q0SfJt�\��}|��oAI˄
<��z��m�hR�v���/�a}k�HS"�|��{��xsy�*�u��G����U�� ��)��>/+_%��6�� ��e��7Z���Xg-���@ؽC3M�9W7F�y�]uS�Ȧ�4]N� f�ĆJ	�{]�X�:hH���(�H��
���V�p��/�y�lW�6;�A��#�o����]t��R[C]d8;x��ծ�ACL�9�&;��[��:9	ʘ�N�
�U�:b�ʉVF.��~U4,Y�R�Wb��;�"K����`��wt��0@�aT��<=����lJ���ػaΒ]��Eo-���n���uȎ
�:�)j�F7�.P�n�w�/vZ	^���Q�W�Ѵ�e06սQݛk`{�3����ڋ�o�x{�]
}'V
1��dʋ��v���;��YT�����1:���egq���p���H��m�X+�[�=��n�m����Y���o#�[*v�h+���{�2_9��R�/�<����U?em?
�R��<�R���·�ƭ��Kn��b��N�HuZNdF��,@��(���&�-��li�=:ZW.���yB)��>�I��cZ9]u+'
Vks������&�,>��3oZ��T��Shf7ܲd���oY�H�C��%�������G�g*�ӱW Z�)�ԭG�0���5���^�1�E@�������<�{[3U��.����+��S9�ymҏ��5 �b�*���,�C N�[��ճKڒ��g�5�	M)wtE�:�X6ݲw�!�Q,�cR�f!Z��r���M�c1emem;ʍ[�)[�k͓v��A6Ӟ'�l�����P�^}�����yc��0�(>'+����n�:t������Vu��'A�;�Fm�0ݼdn��_](�C��1S�(@v\��N��u�ROs��Ѡ �@�E��!dje&dQ�Ĩ��(��rXF��h��ʒ�Z��"EV��TEJ!в�N��Z�,�ғ�a�pK"esY���.bb�Αp���Ej�c �(L�4�K5M���CH�\��ȕ�t��Q$iE�s�9����"�3h�EQ�O#�pIJNY\��L��IL�i�HD�d&&��j�)�Y�eJ&TA�(KD�P�9d��Ra����H��#�5i�j�s�W�R�*Vf�Y�T�s�9DE�H���QU���,�H�Z���D"T�ʑfT��KbdQQ�R�#�DQ&�����U��aR��9�+���*aӛD��EP�bf�+�	$Ұ�%���jQp�5��V�h�"�s��8�֖5�%bek(��r*9�U��J9�k���
IA$��JS����ds-3�Xi]#��IJI�*��b�()��,����,���f��H�e�1ǜ"���S%)S��Ο�Ϧaq�d�"�'i������(1uO���*1�m�W��>R� �P��X�vշ�c�yլ`ѳ�v���U�UDC��Mgij��A��Ͷ���󑫨l]P�
���xe4�)��q�K���j^�Lʹ=:oN���=�nc���ve��ZD#�Ht`������̵�j�ʿL����+o|�&,n��;y�e7�:��9܇�%�|���6���oj�� ����9���%�$��֏�Ĭ�b�`�dR6���T��h#S��>5S��w�*4sz�7&-W��ఙ��M�k®�BAg˯'�Սd^@�	
���[u�,�w'�uu�߻<�M�%Y���l�0�(>�X{�����(Bȸ\l�ߕ�lA��"�����d�S�W{�D{{�;������Z�!l�	�����WyHr���[UX�=�l��(����wb�:�l��χ�ԫ�:N��F]PJ��ᦌD�sSPE3;h�v��iTP�"��[����>���%l�S�/f�ٚN�LT��R�r�N���F�q%tr������P�7���/q��������˖Ù�̮������4T�bܨ@�[����YB���n�b��P��D\X���{�Ѝ�/*�8T{p���n�yL��2[![5H����r_[�gRce��R��p��}��4Z�SrL�k��X�n��w�7�L���̫�iʆ��)ҽ�O�42Y6��3iU������Mf�t��f�S�^�P�ɚaH"<ǘLWY�n��=��R�7~��h�s�YOx4�Y��R�ԥN���5�Z.��Ŀ�U����N��|�}�}(C�*���\b�iV�{JPЭ�}�2�vj��IR�֤*��Ɲ�!�/@��@ˍ%�b�	�\�Y�gYDX&2\W[�s�S�`�?;}�q���Cuƀ�uEW+�x7iC-�5�w�����N{��ݝ�o@B��kaPe��'��߳�x<���_O"�i4h���K}�����C|��6�n�ES&B��Z�U.`��t%p-�,v�}N̹;��D˩�q���h�%Ѹ��.J�'nq��h�I5���	�z b	!Ą-r̅�]���×��!1չ=f��Z��׶t��FbprKITP_�&��`$�Ip��뭥Ƽ5�w�)���V26��#�wo�uoH���d4����RY'!�| �FH ��	�+N���w��s�+���<��)��cE�q-]	�R��Ht5C�^/�וp�t<^�u�@z�t$^]��,��}�w�9�t�z+�Xt���Z'/+½"m׊~h��i*&�N��Ss��]���}Dꉸ��.��#�櫗�k/]���GJ듪fZOiJW��7�����]l�	����M16��rvL���[�s;��TJ�>r���u6���UTD}��h0��B��{��I�V�}���f���X+�B�/V�u1��� �H+�\QG䷪-��{�$��ЏTܥqz�5r&zm&�K��b6X���Ǐ"�@b
���#7��G:"�oס�t&�u�r��Ϝ�2�㊨`mِ�ә��F�Ӱ�[�rq�X�:*OpݴW�i?*v�u|��<豾1�&����Wn1R`P���o\ ���,��k'�Tol�l*���:� Q�cm|)=ga�UE�����=���.�N�7{-�!ѥ}�E)-p�|��<�s��R1u'J|1q�e���^W\4+�:��P�I����bf�Sɨ�פ��������v69;�!o;�j���W�����P2�S3֏+�ú�s}��Ύ!�Ӳ5����u\�u�V�e��.�w�=_̺�Ϡ��Us##'8ݬ��t3�Y�����F}�e�r�!y�;����f��fc"�3B��D��7�uڐ�M�n����Ƥ7t�'p9�z��,�|:�J�X	����+~�Kb��i�ԯ�ż��]���~1L�	R��`,U�{�������Y<�޺�o7vY@/Qn�xt��f�6�i�"��
��-b�iTUfH�j٨�JPMZ��
�_U�Z�܊�䃠[÷��-d�/S��2�,Vͭ�I����}Ir�[��E���!�f�F��4�'GQ0v|������b�.�/��3���\��q�ǐaw=ݭ�&mY��0�}���CWA��,(�zK �#JX��*��* r���ۄN�KQ�=Q�O�݊~f])��X�Ԏ�N�z 0F�\���zK+1"|�:*�re{f��QW6������7f1[G锬hx���W�N�/:KGR�܌:������U2�D�ߐ���.g"���3��m��ўDk��F����!z����v�]��r�{� 4�A��p��}%"*i}�����6WL66u�ȷV
U�9�wٸڿ��Q#�eì��Dd�!�L�L�A��Ba��$qІ�Vd���E���3�M��1Lz��B}���+�C��Q�[졯�r�Y�hV�����>��l��U�8��G(̣�چ�v�Jjw��v�҉�j�|��h�Y��Y�u��S_�H��J��[�P���s>S�AO2�"%1.�ۧ2�[?s����7��B1Ũ��n���dk9vN�.�(� �u�Z��iwˍBﺞICH��E��[+��n8_%����C�'(D:�]���k�e_u���;���]�I�&v�+E�I(��t�[rB��7w�n�O�j�K/^�NH7��ܼݏx�pu'?�_W�U}q��ɬ:��������zvjÞ����}���>^=�Hg�vЧӕ<_h7��}����c� 7�bZcj�F��2�+�6O�m��_P�z%na����7�W.�zZΥ�ut�e@���"�X .tvDTE��%��'�,N�jFB���ws��Ɩ�⒱8d��!r�,Sf�U���0���Uߑ��W)f�u)����<�={����X��p��
F�[��ۣ1���r�r8tØ&�R���c�O_Z�;vT&�%�ls�I�������[.��Ct�4�Ϸ�+4Ӯ�k�L?w���Rg�v3eS�Ȝ�..�X���,Y�
9��vP�<:����>r��-bcQ�Cn�QM3n.*����1X��ߎ�E1�k���R����P�ľ��O�my�;e�'^W��M�/���'r O"8� ����ؚs���];�L�辩u��䡰�'���T�[�dg��ܐ"��t�k��R<%�T�5.�o�f�r�Ό`���x����hN�RY.�	I����-^�|��׳6Pa�n&��}JlZ;[W֧ɋn�U��-�(G��&�ä��R	�6�x뼬�n,�_<[�M>S��fA+��o�����:ƳX]0����������z��s�I ;p}9��z!�F�[n�<ߊI��]P�h�1*�̿h:�w����|P�S�WO�&qʝ�>�\�3�n���������ΐq���Q����B���l�L�o����Ec6��+�rh|��1Nd���ga;�1PB�S��n4�\m�����eMT��\E3}�{*�o\)���:�����e�aL�N%u��̒�g���bK�>�vh��Uͷ�%��u'�1T�+zz��w�}[�4�ے_OgucgK���-}��;+7�j����?V���s�����O���4�I�����	T����F�}4\�MĈ�uCF�S�ⓩr(mC�g[��;OY�n���7��n
��W�ʥ.�9�9m]�(޾+;����瓪���[���g)���::��3-M�%1,�f�ݚK�\ѓNC7�o��Y��5ܘ\[�i��e��}�����w.<D�#K�ں7w���M�w�*w'm1S��=�f�C�����nK���ǔ�a������;��2�ݜ��;�l^�j�;;z�m��i�rY� f�G�p��׷�ѳ�&dvj�2��edɥʏC�͉b���{V�S�	NdsDF�7߾���������w����ne�9�(3}j�\�g���>���)���Ɠ�[���yOk�%���n]|\�J��U����Z��S�]t,��0>��Y�*3[͙]Cһ%srO��$�/�Iuk��
Q顮]����\�.�Fp�4w�gM���ۤ�����x+®Ec\�kN��235���ȕz��_3��I�s�����aL�~K"��ޫ�3��|{��3J�V���9.3�2\0̼�c\��;�l
5$�\��ۛ��M��9J�E0��=XJl�ҹ��-ˍz�U����[��<D�S;�)��	\I���2��%i�^�MX���y�:服���K��u�!����!��<_ARjquļ`�e-t~�]�ڬnF���*=���J.�d������y<��x2�9ɩ�n'u\S� v�Z�ɋ�5Ί''V�c�Ɖ�����ʜ��*޽J#�{o.�7[�V:WxW�h����K���׷�H� (� ̓���/�sU�o������a�(b��� �Q�cI���Ep8WW'�Br�y��qk[j����0��J2!�ʦ�I��ݮ7?}D}��7�\��\TPS������ǉS�N5������x2�N��K��!mvk���o��E��M=��<����S�5�k����7�����t�搕��
�[<�@9S�]el��(0u��r��8�㱛���(�y�)9����8�'l,�n���G8Q�ˈH����f��m��dX)�Y(����[U�(y�D�����M�f��!��`2����=ϭ����[<w"L�9�esZ�2�e	������n�ݺ̇��n��߹�b�{t���!�ks�����5srK�:.���9�ݬ(a�xˢ��%������!��I�5��ft�#;�I\ܥ0�����p29gMfT���}ܭ\�eT	���:d��l6zo���hZ��ާ��Ts���'�W���*G�.��^)�K����4��7�*���4��䨎�x�3��9V-�&�Q�}y�� s�b�]S�Y{[���p�CPf�ws�ݦ�g�O1��9g�cN5)]b��p��@М�u�m��r�A}��p�uz��UβH��o���q��ջr��6��#\���>�����ҹc��S���WE��2��%2���{����2X�3�N��2)�\��IH;;�?��/>Cb����htI{r�^���5�h����o�&�{��!}���̈́��a7�V�:T�D�뗛��2��MY���;[�|m$�Wrp���}#x��b��ወm���{w�D�9"��0�x�;��Z�YR{K�twn�g��ڶҧ��0�#^O'��TT������z)�)D,����7;���f���Ǔ��/���>h�gFn�Y��4x�7�����ٝ�w�};�T�U�Y[qG�r'TTe�ݦ�2ȾZ��R9di��H�G�I�~��BnXN���҆F¥6L�#�w�v���8AJޛl�9�9H�g��8:�ܓ*�"G)��[pDX������:Ҹ�η�qʑ��nV�xa��S,�����R�7^CR�捌�v��B�$�-*�lL��{��0G�Pu�j�Hk�?�2����	����$��z���rn�G�G�N���E�q�G��N��$n&�jOU�u���.[4����3��pI�4hJ1��{?DG��W"�%�5��;���,�X�g���C�oq����쁜NhFf���y���ʝ�q�g�@�U�H���������>}/��J�ǙA�N�ӷ��GQB����ˣ�4%�֮H�"���g���9wFPKx�+�,n^�����9�����8=w"��'�K���b��|JJ9�����F���kX�m�a��%T�Z�A��g��S��{i�t��rX(�a���H���2�r��j�* ������]�&��4-�mt�O:�,���[�eK�L�I9jq�%lRl�!�)��X�9Ӫb�ݖ/��?�e�ۛ��Vo.�^��ՌN-��䐝��w�6�5�&�G�����J���"��'�1T�)XZ�h/�}�R=踵t#��ѭ.�����s���;���x�_A/'{��u6��
`�=V�齈^��`ʍ��y�כz��=���G[�d5`u��0��)�h>
e|�js)�j>
��Nԕ7f[���}�V`��Et;���+�
�ϥѷ��c��ݎP���[A^ *����cxԥ--L��@K�F�W�P���Q�R�Y�y���V���79}o�8;�+�bBJCtfa�
w-:��y�񾺄�����i�.�@꾠{tolF�Rj��]K�ȃOjY�]EFH
��A�kk~�<��G4L����������e̵�s���)���ǭg1Zkh�y+OP�9Sb<��4a.���l2�Ӹ�-�+�Cre�ͭbf�k�V�(�2�-�t�OSz
�qu��e㵄��b��cL��X�mAt�Q�����P����V���"F�h.���kH��U�_2.����Z9%8)�h��#�JQ�c~��y���`�leN�bhS���[:��}�/oN�T��Ӣ�{�5oV>�]b�)(�iQ9w�,m��Z���vܹO���ՄU�R�e�S�Uӣ2��h;vΰ۔��mJCܨ�u�wN�;���``��4m'�2��tt�a����M88ې�n���d�2:��v�֕�-=��9b�M<f�v$t���Ը�V.�&�8���x�����^1%f���Bi	Ɩ�$�ά��acR��i���g'����Y)�[�5����s���KT��f֩"3>���4.���y;X.��56��9���)��2;�X�cM:�WO��/)����)��,��^��� �p�R]��jy۔�[���8<�۱��X������ ���R
�L�5g��"�W���l�ΞYi��*O��Sj'��e���
��$�bE�-�P�E��/�׹[̧�b��
�˴G����.>���g(�/�T�@��Zŧ�"0�(m[���}k�l���vr�����b�����؈�7J��Dn�hp�0WmI,�Z�sv��gE������'!��M���%�:X�#�C���
]zʗq����u�hǭ�iީ3i[�8��7����5q��X*ҥ����o]_cn�|#:Zu��u=ՂN���Fa`c� �JU�#@Ԛ�D1Y�>ɯVf�먃���;ta��*X��M{�uϳ3um��θ"X+,
�׺�	C��ns�;ʑ�!S3��&�e�@�� MrW����w�0��T:�VD�td�^V�/�x�ۿ���k�����6��1P'K�u
��t'$]��Få��N����������.
hYlE��:O]���쎮��n��V����p���Ef�u��q���\�j=�d��b�}���9V��+�0��'%�����]��a7��;*]��(���˶����ؔ��w_c�/-9a�u�(>�݂e�!v�/D�vu���f���Zgv[?)M��1#C.��u��r&���v��}+����we��]�I/�g�	��\�$i�j>��UiF��#Y	P�E�W(!	!:UQ\��GS��]iHs2\l���:��TD�i���B�Rؘr����-B��R��Pd�hk��$$�D��@���F�)��ª���Y����,���j�B�,�Q��F��a�A�db�m":�*Je�hBAU"���"�TUT�"���a%\�YE�C��r��F�$I��,�)�Hr*�����V�E�t�82+��®��A�L\�����˅]2�YQt���yD��5.�E�jJA�*8�^0��r<E��dJ�T��� �J"9A\�"""��x넮Bj���hEeK(�ͤtY�+J.X�f
�(�ЍTD���D�:ˑD9e2�Fl�Er�g:E�G"�PgU�K�R\�<�)6QUUAF�������֡�����l>��o8GY+�@5y��8�d�Jc�\�7�(I�j)�ge2�:��7���_���"#�:]���66���8�3�j��1}\�k8H���Iʪ�͋�������i�v�(�Ӈ�^��������u�)�ۚ�fo��`U���ۜi�z�ҥs]ƨ8���s��9�#���ӣ�Nn�W�]�M��YxZ&�Ȟ�F��%�OSY�����(�e�����9����Gs�9`u�=�:�]n:��R?O7������J���5�ؤ���b~vS_Y���v��D������UT!��ln��d�$��v�~�A��>��W�}�-�%e�?3Pı��%7�C���Ƚu�L�HU�q�Ʈ3��4Y���7;n����P~&�Cꙑ0�nF�)��$�4�c��+_st��7�l6zn1����J��Ǳ���T*��0��_4TES�2�WS/J�ބ�NY���si����#�r���26�5�J�v�.
���rcI���4�u�(�S
��*�����P�A �&��rT�G�M��us{��3�B�\u��$��qOu���T1}tioR��t�ܔ���5�d�����w��q��CZ����UW�:�I��l��!�	��󫏍�Ց�)�*x��m�d=�̺�5x}8�n�I(��اlr�}bx�ۋ���/�5�����ݓW�l�$ީb�n�i)Ã�ȿ��g�î,�#xl���>��E�����Gs^5�g��XJ+��\AN�S�-��i��{�MD�1��U��V	5�J_����{�g��y�μi�S�kc�ɽzL:7���OP6B�C�������^p�����܈<��Yy�T��o���{>g��crۺ�s�3���ׂt�	)D��*�Iw����rs��Q���b)�30N�����S��W,�Up];���h��7*�g=��+�~���B{íK�E��9<�Y7�j>~��,�w��W�G]��Iq<�(3Ԡ zX�@���Sc3����qC����n�{��i��i�����Z�ꀠK(`����[:�uq�[�l_S݁�L�L�Q�����:���m��g�	F��u�խ�W���������1�G#O3��[ԛ�y,��u��N���#l�j]�f���*�w�٬�R���q�;kv�/����'F�)� � �v��}��DGqy�K/y*�w�9Ӫ�[�fZ�����`ƮnIs&�1G']b);�h��L�L���v��'�k\�s�=#mR_-�y�;�4��Tk2�f�o���K]=%�0��\�[�NB�kg�\���ڛ:��O7��7�p����&_�P�YB?wT	���'��uZ��_�Xx���''�N�m�[�)	F[= &j��=��	�	ȺΩ�g�t�s���B�e�~�㔪����`;���<����әjҺ�O�|��$��7M��˗&lZIȸM�<��Q�ĕ=�N.Q�C-��4T��,eeӘ��/�7�#V�t'&�oA{w�N�d󌃬Wi�Z�rɜr�\N긥�|��3�BT�#S�k����'��/o���\�se�����(I�ߵP��?�;���D�u�̟oݞW)�cU�t�m�T�|#$����V{<��v4͕�d���L��ն���^�o��n�0�T3�t(g����xgJ��E���][95tW��Lh�*�g �,���t�u�)5ne���j-4.�ܛ:Q�d�0tD&�`��C/���W�U����~��YAf���~{����ݸ*'ڮ����>��:��<����ݕ̫z�B��6�s���mqƸ����v�ʉn�n��};
�oa{�k��ȭOt+����"��E4�}H�c|�N�$��>�黨58t'�w6���H����;�f�t��e���9�2�@Ψ=��Hc��E���֞��fi��R��uۥ���o_Kx�V������\���Yz`䤊��q7;K�]YWA#�r�T��'��R�M>�f��-�ط��D�%�5(�$�a(�'��5'�z���lE=�|�v��gr�Qj������Z�fs{J����:B�	T~'�|$VP��=�*�+շ�LQ��)����"T���m��LT!(�Kb%_��b�sN�bms�=�ɛ�>}-'��<�i|�2�r�� �J��K�l��vdv%�>����˧t���>�twgg	;�[I:4���V�Ǳm0ٛ�=�:jё����J �8��a�����$�ӫ�����S�u���\*���O-;��F[5�]'F�+J�N:�=ʸ�v��{z��}�I������a¡s)F�¿ʮ2���%;eK�Lش���|Îyl9ȫE�Y�EM���.ؿ5s*��U�n���ug�ˮ>E�MP1��n1Etk����ƺ��z:ܽ���M$k��Ѷv"����������:�n�s	��U�mm�IM
.!q�1�����|��ӌ����y���-�ѥ��fwg�Z�$�6��4ܮ��6��r�����V�Z�]�:T�������-�R~�[;��T^��਷!����C<osٗ�/Uee�V$"�{ǒ��q����̭���3�:����"�E#����Y��M�xq�R�%�����^KVT�a��j��k"u��\[툶���9�wW�<�b�,����K�Xʉ_���P�%J�'Zܧ�ֹ���y��M�o�!���o�5L�|	��ߞ�=������v<����4o�(pj�X[�MzX����n{c���݆oL3OW���6e1��S9�J+p�ue��-���X�U��;KcTr��n��3;�#ܫT� ���#U���ݾ*�܀��x�ڑ���PTO�꘳�I�k\�T���\��W�P-.\�ֹNWW�r�e�_>�����IY����J��:�0�2�{%�c�uv�e)�����lպgr�3�~��n%(�NITlT7�e,��祮��'M�[�C��x�:i9�zb=7��[�k'���u7��:����O���������_)Է�W�4����ƹ��w��228跙�ʱ�7��J$lz�<g���V>{1�ߛ�>r�q�s�ii��{���lts����ZxE@��	j��������zS�u{'ܸݚ��v��TN$�$ؼIȸo�=c�9�!oB�:�:[��Ls�ܮ��č;<TU+����oAN�#S�1���۾x2��&1�=�n���*�l-:��I�Rݸv�{7�Ϋ}	S�N5���޽��x2&Lչ1�_sܞ6QU3���Q;��\M-���/Yf���Iѩ���mv��i�ھұ�3�<c�V��듯���3����e�;o};s��x��0�
�<f{K�\�z�x�uz\�}<�6�@�S�s� �k��ߟWM�4Fق7����Oh�f�r��5�� ���56	�f��hҋ�ꪯ��m�{��]�~y�Nf���ج���NLj���͂�s�y�,�C��������$�{�߆����f�^Z�>�uО����A3ӽ����g7�Ub�mv�MdS;/�9�Ꭹ�";�@�t��������Vd���%�)�u�����췹�r)�rq�����A��@�����V�<E�M��;�f����k>���}�1��9�´P]9��xهڊ�3��N9���D��.���4v�7H�� �ٷ���\��lT��}Π8�M�-n�!��3V铈k=���5c��9"�Vu�l�9�Y*z�!P�����K��K��/u6�� y�t�!�f*UK9gR�2�AŹܞ�M�_�ت��|�Cj��yᯙ�"��p�Xl��C������L��2���}�)W>_��k���Ȑ�[��ktF,�/NB.�NMH�
Y�v��q-3pu�����5+6E�c�<��[��Z�᝟!S����9������2n	YB�AK��òl������)��N�E�sxȺ�9�CW�G{�wKS���]m�������>����Ɽ�Q��Ь�V2��.�$�z���R�����-�X�+�����KR6T�k�yA��}��V�ҍ��)����n_����Dl��,�o-�\��.пn�ʫث���Ř���J�G^|�>�ᎶZ�v���޾J;'\cԼ�sC��T$�oڅ���y<[��GXf�k/J6�>HX�/�ǒ�.��~��ô2��wnʟj��ۚ>��[�'a�w��5S\�!����T���f��Tl�[�"��������Áo�o���_����G<�Pc[�H�9M3�H�c|��8:��� 3|�
���d�$�Ӊ�����z'����L�2�D�[9���ZQD�lkJFqne���Aw	��IZ�by�ϟKz�^�$7����"
}z�&��%7˟�9�K�.d�P%�t8rõk�ƽ����Y��7p��� 'mUe+���R�����=Y�\׎_Rq̡ꏂp^�j�-�zh�0����ۡ�cq��+��T0�Û��v��QuAp����C��4�GWW�V�X��֩D�"�ܯ%J�qhU����^��Q��'�wkz���sg�}_r�;y�*3[ކeu�􍿕%srh�̨�S�i	&�OXۥ���x��5���t��,�5��nt�cs��
�%Q����]9��l�a1i����)Hμp���'4��济�m��1P��5)r��'³z�>�K�o*��}�6���E�a�xƹY/b�!Jkp�����7�/V��tc�AQׁr��G�	N�eK�Lش���C9��5����5X�$�&��L�8��&���D����܍�����E��Պ���_TKL�]
�\�8)W�R{W3���]��F�Y��q��s��j���d���3
g�%�,$�	7ڜ1n�Ҷ���ˎrh?j�I��~�k���B�4���}�PS�&�3�����|��kyܛ�{�ɖ������2$5���d3���j�����I�����Qnv�����D3�nƚV�x�s\UU�!o5:z� �ُ3�ڷ�W�{����Զ'�t��}�JL;q�1�v�E8fK w�A�e�o�W_���tdO�u��sv7��ty���Sd�&X��
Z�f�[��4��\�C�o��� ۼ�˝eq��S�����թB�k�L�S�PyQ%+�����3��(�3`�S��9��-v�؜�c�r��{Yz&U��z�%3�����B V� QwZRMS%�@����s�Ǭnۙ����Ԍ�"�(�$�h~t����7�;Ū�|�t���!��g�lj��"=D{y��� ~V+
�0Os��}�EX����Y)�C2�gϥ�����K�&������#;3@m���p��Ea�1���<�l��B\�ߙ�7XۇIEJys�N\'��'���Ӈ�ʈ�(��ϸ$�P�k�8饌o>�l��7<2v���[j���&��yS���Wn,�c��1;FOI�r��2(�坚�;�Nm%�\q]ШA�q!+��β�Մ�l������u#8kx�I% `pt�xÎx�W.U�"�{��jU��^�3�
Ǌ��DB����a�F��졺��d��?o��9 ��郼�B��Xhаq<��tK�ԴP�րً �:���*�m`鹒13q�@��N��)ua���,��b#c��j�N#���vV�1:�omK�c�.�$S�N�D}$̮uQ[�29*�e29н��`�Uݵ�[Dd�)C�n�CO ��q��`ں�&�� Ђ�{oO^WfP�n�M��Êݳ�� ��,��xEG(v�s��ٕ�(8GZ�H#��1���iV*'����B�o��:!y�3���Bj�:H�D|��hӯ�kܰrW5Ԇ�\ؔX�N�Շ�0�C���јD.kx�F4N;W�<۳GO��X\�S9��Gw:���J���h�2��u��Z���hXJ���1Z�� d��dҡ4^B��ud:��B���9ʅX��d��f��8����YDJ�9 ��Sx8;�f=W)ai�R}����Em��E���T�4s�z��pcw+���U�i��	������L���6�Mva�˔-�h�94�S��U*��M��	��!�eM���d�邖[{(+bT�N1k��w#����wT1U�Z6��iM]�q|"���Ϟ�����,��ܤh��N�C���+�e����N���� `WV�l� ��;���u��J@��q��+����F��f�b��V�w�:S�����<y	Y.2e��t�D���z��X��]����neI��f<��T�5���Ӿ��bۻ-�}�sg��SQ��]3g�s�V��2�2�\������R�V�k�P�WY��:ˡ���@����NmL����s�\�y5��vjVU�)nZY*�`�:��2L�l�qB��߂EB:��z�H��.�Һ,��P��Vޤ�I��]�u�d]8��H�̮��ʰ!A�idz�Kqo��9��:y���o\�"*�4�!�[�nbA+�J⦯�&A�֥J��L[�Xs�>w q.<]ݙŎs�\yC���w�&�rg|D����-ʷ�e��\m�w�|.ֻ���5%�ovIr��-�<J��r�jY8�w$shdޝ��e��Oޕt��ʺò��Ke]a<1�gnM��+�:W,m=�n�����NuJ����M@ۛL:�Os9�ZۄE���6U����i�);O���/o\�.�X�^�
K��܆�[]��(��6�{4���V�q+��B�ha��-�0ƓD��F���\�zN[*���]4u�7����)��e[#�JY�C*�A�,��Y��f'+-U˙*r�n�/_
��Y6wD4��\ƶWI�|i�E7��1꬈8]+ʙ�Ֆ���u�Д��"�p��<�c�1���A��(�k��I2�[�v��v����`��{��g�:	����9#�A�3{z���-i�`�����'���kn��� ���������;�F�r�ډeK9�"+��9T˲��(�2���UY��XR!�**�r
$��NΒ�\Q:ӤQ�N��(��B�(�+��YQ�"#VBIQQQK3��(���Q��Rv�Ts8!L�.U�a(J�S(�TigQ&b$EUr�H䚈Tjr�9�""j	E'��is6[,%IȷG(V��G*� ՕUU�E˓��I2�`a!TG�8Y�ur쬒,����#��P�d���K�U˗)��E���U���\�r$\�G�XQ��e*�����j!�\���H��Z%�*�uC:G�As�˗�͝�<��+�H�����޻��F����ޔ�f8VWy��kVo-���ą�U3N���ٯV���5�F��ad��7��g�r�m�vٟ�}��N4ˀ����.�9	��9�ף�9�!oT/�����6�*�O�W�d���H�]���*�zQ�Y;�N�]��'z�OY�<5����u]i���Z���9|���o��7�Ϋ}	S���߹ܛ�{p�-�0K�=|�;���iJ!f�c������-�ȃ�*/Yx=���,�ԅ�%/�o%g���6^�69eo*�wP���'V�ю�RroIx����_K��IȆ�/��	[�~���c4��J�ͮS��=OYHp��oM�[�ϩ�솹^n�� �]8��(�b���Qg����p�`u��k>�nn!췹�s�k�F��kC4e�s2��~��+y���a)P���o��`�7WS}��[��_[i�|1����Z1�y2�_%N�T���2�t�fD�����R{�5�>�;��B��pB#E�4j�X��!��'~s�-�u0 ��P�� �"���j�ٙ��u�V�u�@	/��	�D����HH1�o:]�+W�5L�}�cV��*�;�8iC�P�A�ˢ��P}�J�� �ZǽZ�	ōv-�S��#�Y��`��]l���zF�����XPt�f��>�(\�տM@�LчL��Zb�<��p�6��GICn��OM�7=n��%�ؗ#��M�^��CQ�G#U�"ڭ(���QW8��,���oa�ٿ�}��	Ti+�z@L�����\ƛ���V���R�f��[�=i-�e�1�Z���Z��htIv�Gt�rs.aK!�Y:Մ�rڼ�}Y��\��3a$��s�[�s�7ƥ�W/ywGmV���:������yu�#x�
v/�N��q<&pX�h�b:�_v�	�¢{�`��7&�\N���b���:��~�<�F��t����M��vi�z!��*��U4J{���D��܈<����xn��g;x�3c���[-=g�O?��t��N��yQ>�k7:�kN��Kx��)+��J���j]=g!���{�6�ݕuK�U���<�#iŜBs��抛]m)y���7Lc��hX T��i�m��h��S�1u�G(��V{"BͭT���sv�eͶ�hxp,Kզ֖6���nL���K����g㛖���G��Ok;r��z���S��-3�E�<)���s3vF�BrC��}~��S�Q5^�J���G"uA�Ny"��SL�sy�Zlv[��Gh�҂���-�u�:�xvէ�����)����ZXa4�S,�΃.N^�qί�-��(嬎λ�Ps*Çf�>ɳa�V���}-�^�5���ט�����(�� g��_As&�/�YA#�,;�V���F0vu�M���Ҽ��+�����z��!�o�w(ܞ�rA��W����k��H��Yͭ�p����Λ�nu�6�~'`@���2�.�IVi�.[��\IA�����m��LT!)�69];��Mk�q���f�ɑ�����Pn���"�D0̼�c\��{�X��B%s9��(ɰ��$x:�Gh�m�.�3b�NYQ�0�u���2��I%����P�	��tb�y���[�S;;|���	#1'$+����[�Ez}���ځz�;����s٤�wǲ^��g�<KRX��V�_t�ҥ��C/~o��b1��wR�ɽ�&3A��Z���_d�/4Kdb�'OwF�Θ�s1qw�U+s%�+�J��BV\�i���eJ.2D8ձ����.��U��I�ϟ�R�|w��M�8Cy؞s���w��oms=�����{�,Zg�P��(`��;"w������O��/\s����q�*��Eҕ2�+�J�gsR��L*{���kyܛ�{֯r����dn���y���f�8���+ni)�<�����Qnv)�9�w���l	�}v'�B�
�\ҕ�ѻ;�o$�0n�(g"uA�g��"���w��Z�-ߗ���Q�wϹ_ѧG\[�l,������	G�ӭ�슍s[Y��繥*�Ŏ����3|v�R�� ����7֠ �/�p���]�K���.W����>L���q��5L�|�P�e�����vbI�s��u�W��k��Ч��]��_[Һm(�$��9��Ua�����:R#�r���|��5p��K�:��z�s��uM\��*j�^:�l�X�g�s9Rtk�c�������}�"jt�O(������_�s�=J�(���4+����s��3|c-��,�����Y���gf/<��N�e:-�1Z����\�,�FWU�_4��Cy�T�9�����W������L�<����+���Z��S���N:id1��[="��֖[�v�(��n��%Q���_Q�c��P��= �ұ��K�����GIb����m>�v�B��"zew�Y�f�s��h��d���=%4g#洵s���B�f^0�B
��=R'�ַ*�]�&m��Ė��,Ɯ���o��^����m��D��v&��Y{Y�i�|�wI�V���^t��U�ˮ�E:1���n'�=��'�u!���W�k�sֽ��N=��b7��μy	S�Nϵ����#c�=-��J'I��nvȜ�qX��h��Duz��
��3#e��#%���ma�z9=�y�j.L�w���?	�W�e�=�:~U&,�[��-<�R���������Ľ9s��;*�$q��S(��}�޼c�*{|2F�t��g���}��ܱ��Pv+y���J\+������'�S���¦�Ф�_5�Z:s�bp�w1hє��y�R6SeJ'��XV�����,�veU�kˬ�r���	Crrg�#���W��^���5 ��(���}�
�u���yM2f��F�qq�@���Tj�zoU#K�G����ه|�ڍnO�e���!����8è @���gn.l�.�򌙶��n�7v	�E������_6�󜗽��#�6r���$�T���p�e�@P%#�,;�k��R{�5��������M�.	#n%7��I.zKF!w���~�1ᵚO�s�d.��I�*l�iT4ϡ��ѓ�;�������A�Ų,�(^_n�J��\1�7�o�1�P\ʧ�V:���/+��7�;�j)V�՝<�7�:�"�fZ��+!���f|�	�U�'Lz��{��{�S�W��V�y}�����i��sp��y+cX�{wwJD)r�L�)L�.;�B�U���F�}Y��y�����ṾMЦ^��9��/�>w7�tKr�8�쬺n�wP0��������uӺ _k�-ʇrm��4����{oh��}JP���x'd�i:���7d�j�).C�Z��S�T��6�$�%n5¥5ǖ����?�u����>ũj�~�j;��G���!}�5P��f�븺zd�x�i��+6��>ǝ�_$������U��AM>y	9[����5��el�O��	�"��;E0��$����ɿ�{y��3+�Օ\�����s��w_%���5�6�E|u��Qnv����]y�5ۣ��ӎ�+�Wg�l��2;��3�N����7	�)�r"��Ȇ�b�B;Qm�'��iH�n/%�r���<��ʓj�3{%��v�OOt����m��v�6��u>�Tfv���"�7�u��*F'��Zm���p�h�37���a�4������Y��]��*%��tU1�d��"C��l�r:�)�0�nZ�����zuZ]7&��̪5o֌���;������/�r�#���>v�_ΙK��s����n*�W+)�ڹ�ga�9DrT	��5Q>��s��囋$ش�)L�D�Xqw)4�_����>�R�zj�O5�]ۚ8s	�U�\[��[*����F�̕�-}A`�;*d�e���������r��:rN�� ��R�K�5	����üt�}�0��u)+&�~���Q����[�Y6�xg;�"r!SK"�x�l�ư�L�}�T�<�ܲ��$6j㋞����^�)oN��L3/!�sJ���"d:�w��k����!L��ϢW:�6�VD��*j
���>��͒u�U��ltsS��Cv);�����E����ͦ��������m�6p�J%��&�n3�9*��B�Xh9���Z�e��hl��7.���Y��Sw�{�p��g�z�58e߼#����Y�_O_�x�
� ��4���k��|VbN)�۷�ټ��g[�J��$��w'^!B�e_=t'����U	����v��.w(�e����oYϾn���y�Eu��PՍ%8�w'����������n��k�:����A�/�%B��̵}×���9&^�\��3ς'��놯����~Eץ&�h:���c�"��hE��
vó�S�W��U᧏�	������M�6�����������2�ֺ>f�c59����;�{�´vO�1���<Fk��t�Zi�)���FL��Ò�J*�����3u�,�n�B�V����$��F����}UQ�7�Ū�rq#��i��g�u���z�q*�|�O%l��2:�M]�Q��J'`S��9<���oO�SL��7'�X%L4c��m��Z�368��VV�¸6n����i=�����_�ri_N�$�.��6�����
ӎv[=[��O��.h��Λ{9�U���1�z��E)��7&����M������̹d�C[�;��ܥk��$�qke(�R�	S��̛�"|id~�3�N���,�]7��Ez8���^1�n!7�n�S=�H&�v@>�f4jG�_]Yg֖$�ޣ�N��=p�a�e�Z��MAS��_N��o�-g��8���I&cX�wdO�Uv���rn9�J�����*y�+���,�M5���eOnB�73(�G��֍��p�����r����b�ҭb��[�瞝�j�N\Ϥ� s��:
��@dJ�]��;��\�Cߢ���4&�<f=4�^��.d��@F��f��*d�H���*S �={ʎWd��W,}ndJ�#�����$�P�%u�D��|��i�ꪪ��2yIv��(��_s?Rݳz�7�Ϋ}	S�N���'&t��蟗�'���bsw��e��%��Xo�+�t�͞W��M�*;��n):E #%���W�5#�����	�~�.�sɅe����P��e!�Z�ܪz�Ck���'h�;pD�*�7
V]��vLr�\Vo8u��'T�nn-�E4�R��O���GTw_H�	f'��e�o�Ri�!��P&��p�s������o[O�Z��ѡ�k��^1�Ƣ�`�S*uĢē�v��w����orK캒�L�̗�[�sK����:��\�z�(���rXv�u_ʓ�P$;���o5q2W^_s�-Q�.�M{��$Uf�/���߭ �6�Mo��j���I��]�>�I�3��7X���J?s�	�_D*2��y&̝�� �ϛ[�ϱް�����.�̺� \]��$���l���.��PT/+�R6�W'Ǭ��▋�v^���v!f���s��R����Fk={�j9��Q���5�A���J��cX �.����]�T�9�7�$�w���*ش��LPy���&
����*:�ЩmdB��%��N���J��t:�N�Z�n�B�0^���Y������S�^m�@�H��@:j�q����uk���G��Ƀe�ƹ]6��v��P�''Ѭ��C[��'MWp��=
Q\��R�{Ki�YJ�������[�+pJb��+'n���/+�,T���͍Kt�gu�[�y����K&q��a7S4z����};]��ǒJIuFx��o1����Qi�����z��x!�n��*,�w4�?x�y�<6w/�lZ�U��0�ew:�����(Cζ��T9&;E#)�F݇w�4Wf*cq�hPw(�q�B:�!�ŨdB�/=̺�lշ�����8���k^ ���v�&
�ƶ��U�E	�vlKz8ٽMF�PuMNN&���V0R�L*�p���h6g�&�/_��%�,>·�����4��\�jN� X���E�kke��n���Scnf��٫�Rl��y}Lⷦ�P�{�,O�Gϵ�T*\�D�>�Ams�ٹX�P=���t��ͦ�ګ4ܭ��6G4��[
�b\�f5��1h���.�N.U�A��[��'nO����p�c��sAm<�S�=/k���ܥrxn,wVEp�m������uo�������={��ͤ�i�b�ƞ�b�Y ;]��t�׽4� ����	�����#�[�ab��p-��ʆ�2�b[�Z�ܛ7-o�.��&�Kg0��C]����)�A�g�YM�9I�TD͡�%�,�X��u�B�\��F���!x�
.�L'(m���zAˑLi�ν�cQVZ6�IV*��e�b��Tg�����=��˚Z�Q��!�=8���H�}��vS��Rۏmt�ּ�)��)�h�S�z͓��ц��AM�[��3sạ��je9��Q@�ޫ��K;��
ƞ2��5N��O��b�Y�z�2+#�Q�f�n�C��9yV;���`R�Wd}2o�����s�f�0Ly�7��Al۵�:㤥�C���].�W��S<��D� �]ev�G�4k!��c��y}ou����JI%�%�hͬ�� Y�"w"{gLM;6Zᗺ,�8N��b�W-�V7����nĺ$���.�M�M�b���o�G��������N4t^_fl�:���CxC��m��2��4Y]����K'���VLr w3S��' �������Be�n��y��|W���3*�ۓ���݆�{����s/�E -���+ǯI��-!}ˎ��bTV^U��o�s���R�N��76a໪�_oT�B��
�P�i\ �Ƅh�DG(���9�W�$(����a�("��!�*e&�A����DX����Ԉ�&ʣT�*g�/B�9yx2�m��*�PPvUE�*�˰�8T8��i�:IEE3
(����\W��UW(����QEV���T��#J8W(+R"�2�"����s���8'�\�F�*.r �QJ�"�E�(�䘩��j�"��UDG'!t*�$��s1r��EW"�x�TT8��TQU^��A�QE�"e�^2<���W�I�'\%�ҧ)�9�D���+�Dh�É��ܭr�NG+�	�(�^R�ED�9��J�3k��e�)��N^(�Z�A�B
�EXduX�U���s�r㸧��ip�Rn0����<bT��ܑ��"������믧e���&ێ�C�vw)�\�6X�g7���H+yq`.��5����].����H��S�UcvK7���U�:9�%6JR3o�CnI���i���ö�!!S*��s�ۺ�:��K�+���|gy"�e��(��P�)�`����]���Y�5�􂣯 .U��7��\��f�I��7����Td���볒�����.OA��v�\_�r��.9�.�q���{eмw�����pY�����x&��5��F��n����q"Kݑi����=I/-���U�7Ɯ�i9\�gӅF��ǻ�םQ���K9������M^u��S�I�[�M���,�ܯ}�هjW��a�⎪t���sg\Q�^@T[���oz�޽�ڭL{�4�U�:�l�b��<�Cw�ƨ8���s�M3���Os�Gb���,�iL������"բ'�FT�k��K4�N����w�%3�K�g�����ʱ(�E���A���=��)�x2�+O��^�zx�~8ϣ"�'�Ւ�t��`pEI�]w�7��ۭ5q��R�}��t���ܩ�hR�v5���[�N�J"ej��V���k��-�"<�*ݻ�;�d�ޥ�%@�빙�؃����H�t���J4̪�oj�jF��J�YB�+q��m3�8�Mɢ�DJ���%�4j�Dѽ �'�)
�n6�T��|Եϥ����iEI'�h(��vpnF��v�%�"��������B�j�3ik=��鸌nv�ҨW*m+n(J׫iB�EDp"~[�7�s޿��'!SK�y�Ͷ�v�^3Q4�)lwQtQ�a𷒛ϭX����1�tr�o�r⹝H��i�lT`J�'�%�_ܶ)�D
�������cX���qM�E�P>�Mޖ��08:L�.5�6*̏��ė�����/ko�����WD�
�Q�[�
V��8��x�ێy��؞�ɾۗ�;��{z�,��#M��v��,����ŉ;�N��nz�On���S�X�x'���'*1]�����E��/t&zl�4��$����U��!sՄ�ShC^�.�=|�z=�>���z3~J�T ��3�9J��#���<�r;��5av�w(��J	n�Y��>B\Hw`Y�kh¶��S_��g(3:�E\�rJ�OwM(̒�B�q�}=�o'�O����N9�u<u���-=�Ԧ����BoN���ݯ���\�QQz����oEMf|fΪ��m=����Q�y�����
��̕p������l�N�:��]��i�Ņ��QR{U�]���)�o�O��ßX�k=��a��u:r�c�;�t�֡k|�!����6�o�-��)��y�����{`�'���QV㋻�N>�sJ>���ϕ��n�췙�r)�ru�T�R5�D��f��:{���r5�v�� �����-[�z�Z`bR������5��Ѭ	;<�a�迥�$�n���A<乣�Γ�i�ͫ��ys�t�6���N��Z�&�;�j�M�p-n���s6�$�s�3s3Nx��t�6�Kd������:�D�����#�__R/w�8��Pmd�}Xv���2�H��E%D����Ayq�u�T��!��W�T��`dNʨQ�V���٩_)�g6y.T��Z�k�nDuJs͈p�wZ��N�EG�*5�ᗏ[Ƹk�΍6�:�L͖r� �
�4)}6T�y��aB��m���%U�n�-�o!�si���v�|��M%OH�����	�ʊ�0w#�S�0%)o[[�=ifZc\�CaR��zAm�ld����<Ō��&�V�ʺ��}"��&lZI�MƳ�9В#���M�))�V^t�[���\�P'w6����]q�,�����m��}/�]c,���i/I��J��9b[rj"q���is��:��5}h���͏u��]�e�Bz�����S����'C��j�'_o�OZ��R>�TO�!�׾�҆ы�$R��	���npY��e�U�+V�����m��{����*-��S�[[��Dc���}Ƅ��S�Ζ(淞Q��=�!�T�}�js��"�g)��ӣ�&-#qdh<�ۯm�oT~��;�nε	d�ܘ[-�6�ȦY-H��ب����U����׺.��&M�5��N��%���OhT2Mq�V�ԍKz\7UKvl��2���w�:}�B���,�`(�U���qAYJ�'��efq�#nk7fђ�1u]s�9cB_X*�'�j�Q���%��Wo:\zis���N�\�JK��GWL���JȠM��`�4z[{�>���n��^@Ǳ��O%%���7�S6d�2eE�(JG�Xj�WL�x"���y�ͪ��������#PK�������JNo�Ko���-:5[w���\s����:�ժd�B�ks���n��%W��e�Nf���ee�8sݔV��f�p���\Iϕ4��7�ߘ후���b�	GiG.��]n�P���k_�&Gø՛e����;�$Zr̴ƹYlf��������5%6�pQ$��P|�����S�T��3a$��a�{z����u���1��^�|݉�.z�B뗕n��}Y���3���f3w�)�׬�e���n9䭻�h�y{q}U�����t��#�K)*���0S�u�bN�58b�Ε��r�����1��df\Ӹ�ԏIS-�0�O������u��j�'�p��u��oh�p����v͎w�;BP��"�z���t�h��i����<�{�8�s˱Hܮ&�c��cg]K�{�N:L�G&Ʉ1Ӄ�cpKe�w�����_]�3x=�`.'&�s��ˊB������w�e�T�!'��7���C. �ݸ��!1�N"�r�5!ļ#��S��QQz��
�s�S�r��t�v�#IP� ����b�\C}]��C܉%�VV�P�D�:��2�u�ޘ״��&U�gH��r�w{�C�>�[wZ����2�߭c�������*ՋkN����f��|�ȦYφq�Jgzu ���R��^�Y���p���k�����[)bҹ�4���&
��
��wE��7�b�X��/$ؼ����ӪߑO�!�k�K���]6�T�����i5�Y1B-���1�-)%f`����D;f��;��4w�gM�7;n��(�
8��IW���f�|�@��k�����8��ND:icϛ� b��ؗ�*���mu�S45ä*�G�'����D�I�/�=�d���Yi�W�T�l��X�G4{�K�a��� A�30���%����W}�X�:B0*|{����{R�{xe%P�@ɻ��i��6�_5,�SR�,�d�-S�9Sԁ٧�t��3��T�ls����5u�Z{��U}sjse��.!�0nBW��W��ωN�v���E7p�zZ������l��s�6)Z �퐝�I��� %;�J��6�*(+�����6/rq�Ī�v&���D����:w��v�լ����ﮟ���s{��f�=���Do?E���zG?^�d{Eh7�>�F���ҕ�zj�Vx��]G8��f.��X�w�6�٧3gӿ7~;�?\�S�>���ϔJ�s���|1ZY���t�<�U�;��C���`
: 3>� \���/�?���m&ïWe�g�6<�s5s�2�7��Sd0$������J%��U�k�����'f)�^'7�U`�>����Cb�q���ṋ��s�U�ex=�U=(�,��v����ut�����=�����W�0�/�d?�~Y}���æ� ����s�-p˽��Zwʗ.G�r�u[��خk�Ϫ�>�H�u�p����-����߅i��H����e�����Dl���ʅs���X�v�:=�qm �Dі� d��1nJ��[hb*`����k����^��r���4�mdݍ��.gv�|r�F�أ������I��Ge�a%�F��N�t�''V��w�u+�i���Úf��ԥ�L�5�oS�A`�����ߎ��Ld<w�mz�=+�}n{Ƈ�(��G�	��~�p�Qýe"T��7�9C����S��H	ΪIV�e�{=��79߳�|���Wlx?Z�d�7�8�%M���%jk�G��<��š1>V*M|�|j���5���<�MOfmxto
�s�s)*=��u�D?Z���'�T曪������5ݙE4=޿���~�1yV�E�,�/�/Ѹ<��������4�x8�������_�s�����@4%�r���ֱ<q��Wy��[ ����*nD6��2=���c�]�=�����:�� ����߯}�'J�x[��Ԩ�5�����n�E���q�"ҧ�|׬O��fP�߬P_?W�O�"]�Eu禣"�Vyp��y�4�J|�=�s������ӱ���_s��6\�뺜~�uAiI/x��f�lR�^�+���l�>�oNN{�u"�4�W���p����)���g��Di��I\�Q4ָ���-��抛�=ʹb���d�~����he��c~6du��-z�����������r
[\2aN�ҟ@�h�w-���u@T|M�O*������1��ȶZ$+��j��;wH�n�QhJjT��;��n�cx`z�JnL��)�Əe�oA����/������Øu�d�p����G�Ar�P�V=8��=U� �q�V�yp|�i�[[Cr98�G����W/Ү�k?F�z�,�<.��:�M���#�N�xx�Wx-�y�����ڮ���9���sO�6>�=��PK��j3���ܰ�����zFD7k��7�[�[�G~��{#F=�֕�0�����67�H�V}4<�Jv��D9Ⱥ� m԰ԟ^Kߧ�~�8�}~����g~'T�&�pK��լ�U{�>g���Zd��ĮIaC�T���Hq̸��������%�Q,�O>��6sRU��cP�����>#~��+'( ���q$y\<��M���+���X���m��2�ֹNU�/�B���}�tv<lO��r��uNY��S3�B\�7^�>MU�c{=�������}W<G��Y���$�/z����T�G�ث�U!��PU�ݫ;v��x����Z<'վ���|==��1�jV��6#c��<�G������ȏ]�Tߢ@��^=}���ʷ�ǣn�84$O������=W�����'Y�s�z��xlG���7���婀i�+%��;�TW-RB7�.��4+����D���#��G���j�2�ѢHE"x��+qm�J����A�*��Q�jvbk�;xk���|�)ض����Ty3��p^S�c�R�����R����os=Qu�5��V�]͌:]���>r=D�S>���,wq�J�ɪ�<�h苦o�3��h���[�y;�O�2�8�4��{}��,��Z�>�1��^�y3oٕ"�0ȩd`��\S7�7����7���[୚�������ZQV��WCѯ�3��{=2G�%��eT��^\��F}�eg�����4U,�/�R��D��[��u�3�9�[�a�s>�����	�����r Ӑ���r����+{s;U��.+1�~������@���4���ӫ�ߛ�Y�}ِG��q�V�bc��Ձ��V~��6_*�O�UW�Ҳ�lt�*��ۙ���������G_��ǽy<\ 	���9���Tp�9�?'?��*���~���k�kEp��g�:��\�xT�^�H���^�"#�y����x{�ڜ�]tF`�	g¡踁F����0㹖��L ��9�י���Q9�R����y�=�s��S�C(�쪝9L E�^�é@'�ذ��z�vZ��}V<I̅�}~����ǎC򭈿;���eD�	B� t���:S��K?~�k4�b����dݸ�#;�Zxd1<'^�W%A�I�>�/m�� P�P�eMY�n��6���c�/�N<(�!NcJ�v������u�h�sF��V��,��u��V�3X�}��C�W���]Nu��{�jv�R7�[���
43V��}jM�j��9��Et�*����k�ߜ�ǈ�)���Ш2�P�f��=�Vob55]s����1n�y_L$���6��:z�Z��N5K��n�*.�/������˼}�gN�j�-�Δ�[����<���|����R��@����a�,S.t��e�Rw�n!�4̚�f�454-P��#�9X�a�Ϸ��o�#VhN>ǌh5�D�O v5Ʋ�	]M/���j˵ ��W�l���V�]墘�`��,<����;���H�&���E�j�����R�'����>�SkR�M]�"룡֬�)����
d7��%�s�4�g���� ����Ve��P}e�BK�K^.�C�A�\�����]]I��K�n�}�jT�Ju;��Ϲ��+���D�r�����2�}OOB��B,�v�nV�n� �t� ǩ��nh!2\�RX�V�r��q�#h���9�@D�i�l�.�fH�oCG	�jI�tȇ��h�%����M˙3*eG�ViZ��ӑ�N���ub��w4�ҹ��w��<��6
��-�K�b;8���%�w����i�_S��:_n�*����+�h�W�P��SY�7y*O\�fS��PF�f�ô�@�*m�V�5ru���:�"�A�og'm��o*�h�;��BXt��.nlvX�V;��Q<ق�vR���+�c�Mf흌d�1�����JEM/��1%f�b�%@R�:���YP �x2�#��dR���mlU{�c}w�A��'V6N��A{n�kk0a��P�V�e�G>����l�Vp�`]�K�4�%7���IW���۔G=�����#&��_�z>G܏��	N[<���`�����A�<JZ� !�v��]��x^l|X�oM�L"�/�K��B[!��w!��s�z�N����y����͎�ݓ�l
�ok���{˱�P���]��!�}�(�c"��Ov�ȫ	
��ʠJU�nR6p�݈�\M��)�y|��s��4��|
�evI�f���a9Qm�<B�%���?=��ӓD��m[_��ֲ���(�ʭ{4Dr�)}�qd���l� 5�+��i(�i�{Ð9
P�wJýu׶���,68]%�t�O�{�c�V�}�����tO-dw ����Q+�&57�(۲'C6�V4u%X�`;2A���"�[R�'m����Kڙ�u�A�rvbA�[')Ʋ������a�V/C�JN���S��2��WyJ���F{���uOP�oE���hE��_�sKD�k6,�����tUÆ�9e5�[�����~���E�"t�_�Q���V�G/Pt�*2�������m<Kr�Q�Ps*I(uNPꇦ�bC�&eL�"r����9wT*�dQ�OOVyʮr�崪�U��Z��q�\�^!
#�Up�WJ��<�:z�U���zE'	�
�t�*
/O���(8�Dr��Ex�q&ȹ\�G&�Q�r�6�J��
��gF���*"2R@���Ԡr�\��k0��D)�8�yTY:��AU�.yJ���uS(���EEQ+�a�ZzN ��Y��%p��H��J�ܸ�#:�e0���Q^�(=0�+���ȎUw(E+q�VG����GW9	�U�*���Wt�z�^ ��(�Z(�4tl^��9a��w����y���{ʪ;w9#[��2sOm�����ފ|�;]ׂ�7Q���N���Óq�!wi0�G5��O�9�c��ݧ<�����x��ʇ�#b<hxr�|�V��$d�/zLz����B���_��s+�L���Nא�#�T3�|6#��Sy��)��ϱ��T8,�}��BY������]��8}E����[�2}"g�١&R�r:RgإO��ܿW���lI�����z������`x��Ddz���(�=�^$ߣ!NK�_e���X'�\�u���*�������hzFπ~�t˷q^u^�Q"[@��3~��,������S3o�T^���L^>([���ɛ�����3����צg���&=�Ӏ5�X`&��+]�|R^V{f�&�В��UG�o�-lo�T�k�q��2�}������z�O�]��ʡf��]����U�û�վ�eI����^]9��������B~�"7���C|=8��vx�O����Ғ��=�����G�ut�^�ӟ,v@;���M�O�����ls���:��	�V�:��J���棽�;��Μ��m֌���T/\Mwu��@�}#��G��w�x���=i�!~������f�<XФ�Jw��o��T�Gr����'����C���{˵��޿���A�VT��v�����9c#�1T�Gh��=�2��O�35R����C��&w�����K����f-�"7���Hw�cm�QE #?yo��S�њg����W_��tn�
���^t�X2��	�wu@�/wK����!ީ��}���>t7�w�lCṋ��r9WP9^OdU=(�-��U$8�]��n�qY�8=쮉> Ӊy=���/��C�{��}ئ��[C�� �2-	��^�1�=����HyM����E�%Q�=s^��}y/bO��2=�<=�~���-���<�V�B=3]=��⣜<�o��V�#ў�#���}!��˥k�an�1���}{=&|���_���q�o}�.��%�RBϡ���(x\!��Nf�$�U$�b�⽟{=�nr�gH���UG�s_,�Un<������jk��P�2�-$�����KߗV���CuTt&�۸�����ի����{֤���X���sL �a	�n�z��Svdu�O�P�⧼�Y��"R��#9�G�T��m��#��7�1��fr=Y�W�h`�lmF)���-��Ƽ���'��層ټ�e�%H���SprY��y����/�m�0%���c������	~�f���ǝ��Zf�<�]����-w����ysǾq�,NE�H'=y���պ���L��Z'Scjl�P��l�s��:�B_r��ag)0]�MG�k��严ˉ��8Ԣmsj�	�d-��j�OW�I��jM�ó�̧�z�d�����1z��2���?,���`��?W�O��<�[��0VR��8Tϣ�ЫpP����״@k�gm׸Z�6��Y�.v�eI�fF�.=wh_��{JWC�j��2C{ӓ��u � �v�����/��1e2<� �����]�O���f��O����>�w�d�m\��6�w�{�+�>�����[�$U��\}j�%�@h�U�3N,�U���F�]@��i��(f�r8vU=њ3�T����7s�.����/�~C����M�.���|
-׼�� ���(gڮ�4�K�qLv���f����Q���r�:3^��:���瞑����[�T}6�7��7�n����1J]�b��Ĉ�B}u�r�H��N܊!�}u^C>8�X{'ג�'�~�8�}~�w*+�sTh����(�^�6g�Ei�U!�`� �
��b�����ra{&r3Q�T֯6���J�}B_z=�s�)�òe�P5rKcɎ��s+�j�B�7�.���R�R���̈́�]��D���W�S)�kw�E���M��u"w�Iī��p68��(�K�=]Ox܆��y�7��sL�����<<%������ctb�9��P-ڍc����]([w]7��7�(<�9+���c���gm��+�B��`�g�ϕ�=�~��G|lO��r���v��H���f|�K���s49�q�)������(����(;��bCa�w�#����S�=V�_ΪC
�Z��&��̳��Y�����S�5]֤d^a�w�QCV�k�cb7��<�G�����ں�O�[ˊ�ي	7�(ϖ
�|��󺄲"M����n��8b�>��X$�Ck=.w����^��^�����{��4�_���j6%٨�!P�D�B��6)�����h��Е��y<零�}MҰGi�{䒐1���\��
������~̩0D��M�c���C��~:��_
ҁ~OB����U�P��=�u��Pȍ~��VD{��=���O��G*�
�l�2V����W�2E��{����1�e2W��yp�~�#y��}C"7�p;���!�V�r��2��|c%{-.�}e }S~��t���<��@�c�?6�<�h��W0�}�d~��G��g$U~����Aj6��	)�b��ᵾ��*竧�6�O@�~��m��w�Ǥ:^�Hq~��I{���״O��켰n�1cۭ�����g"%�Xu�r�λuzk^��.IP�5�w��&�wy�P�Q�P>��
�! �of(��,���B6'�����Kc����s�Iw��ݚ��}�wK���JN�ʛ`J���F���sW�g����^u��$����)}'n�/P��ڝ_%w)���j��;�w3���n<^"摽�޽�+�Ĵ/s�G�ߘ[~�<F�S����0x��P�_�(�:�R��s-�zj]�BiNH�.=�(����9��F�N|���S�[�f���̦ "�/�J��{�\a���gBӏ������WD�/2ğ_�x����\&k��~��Vٕ�0���q��LO�������Җ��}��r꼫Ҳ�0��M�O<F��C���4<�\>��!�.�}�~t�pҬ>�lL�R:g�.��Sa�7]��g�M�ا�~l�@h1�/(_�����ՔUU�z=vD{>����)H���	 /:��XϱJ��_�9��~��xػ���|�'IC.�J���{��Dz�Q]PbИ��h�K�ld���1p\�z����'���xN����z{�Z��+��c������dU��U,�-���k�
���Ҧ|����U�J��C-�����sps��z�G��R=��>s[3�-Ы�L6*���b(g��_~�CMny1�]2���}��f�=�/ %̥��� g-�μb�	\*T-�Et��X�.�L��h���3r�'�bEʑM�#uz4�X=�4��c/7o4OA웪�@cP���&
�8&�(��:�ph��^��'#J&�	� �p�c�}E�M��ca*�׻#���(dk��(d{޹���<�zZF*#H���?�9���.\�ƍ�F^G�ke������~�Q���nC���Do?E��F���w�GLP�kA�Ҧ}�y��Z2<<���=}/>������x۟f�͟N�~;�Lj=�}�P-i��9v�����ޏ+`�y@���f 5���k����Ez�Gj8�ey�C�#@A5���",d��z�z=�>az�x���ڜ�۩�O���&:� ��1Q���d#%Oվ�R䢝h�&���.��9��C~�q���n̥�+�U�}���DU=��v	���j��qRt�(��_��߆G��O����^�|[�L/}~Yw݊o�5�:s�=���>�ck����Q� W��\ �l]RU�w4�!�^Kؓ���X������-�����D�Ϭ\�ܝ6�;�rW�Q�G���Dg�hH7)��Hh9˥k�V����M�^�I��[�q��]�3ڐ-w%5���$�<w���2֨�Ily>%����ow]o��~_��2��5����[;��Y�,^�2�n3��Lm$BY%KY����:@�=!5ѩ�;2�b���1�:��O6�"�*j��8��u!wD�x�/�9F�	U�[�t��n�jaK�p�`���^��IVh��D����9�Z�!�y;�d�����YH��k�VL�ڍ��;�%v1������+G���v�D�/�&'�D8��R�|�x�Lۑ���Ґ��rB��$���w�X���Q��o�bNz��[��	�n��J�����~�kRJ�|�y�d>��r	�7"�6<���7��}2}Y�W��E��H�.�����`�)F��(	�3no_�2z��*nCk=C=���c�]�=������Ǚ�����0U7%)��$�R�7�u�>9��{�V�ƽb}���(F6�����=B#p���C�y��ŕ�w�뎋������;P�D״E�5�ӱ���^�'!�͗(��+�\�Ӯ��|���
�Iީ5^~�L��{ӓ��u"�x!����������YiP
��{�k�t�դ�����3����z��s�O�'�͐F{�y96�w:�q#exg�;�ziP3��n6}�_x��G���=����Hu^���i�� ��d����97{r��+�Ϗ�T���k�����|&�` `u8��W;�Hy����AZ����eWVϷ�Ys?(RD��O��Ƶ�z|]�ҳN��(w(Y|Ep��?*���ʓW���/,�$^�>�MynB&���e�����;�-3�}C��i��v�5�:X��0T� �.Q�ϲ�����@+��pu�&��je�$��^n�o7N��;�~�����/�c	�EӱӐ-��V��2�'�zFCv�="�O�����"�qj|4�m<]�E�Gs��#�ˮ��`$`S��C���!�������"}���s�_��+3O�dߜ瑿0�ԧ�Fp���!�`s&�C�� �뺊Z�M�N+çļǭ�<���aA�{>���o����{����+>���� \*M+��,b�ug��ϱe��<��-���(�{<r/��0<��%���]Od;�.&�HLϕg\�I�j���w���iH���Ӯ�G�/(f�J�Q�W����{�8,�{*{#�lU��qg!\e�mM{�wkׁ���"Ǿ�¸�bj+�̌"���r9�*ԭ�~��xi�0�Tf{�譱N;�O3���׻@�(���|Py"�_��FBG|P��X0��p���ϒX��A�ʣ���D�����}W��G����.:&�㸫�)�95P� ���o�27)�W�%n}�]e�x@5Hw�����B�G�l�ʜ��w�=���w2�wR*`�R����o�w�����m�;׼��� ���V�*��x�GaRU�d�[_hW])�R{�nFՊ�7&*�щj�[H�����(_)=���3�����b�r��aQq��eԣ�.=�i<�>����`J���Ďk�S��n�E�w�7��ꌧj�6䱓7
%`ռx����c/��dx���g�b��~��R���${e���mԋ�^\H�dO�u�ۘ=���ͪ0�j++�W����CC��dg�sr���69��˟�����z}.���U/���������U�H����Ȟ��[Nw�e�Ɵ�F�Yߩ���k~�>�������z9]����w��u/��#�
���,'��������/�9*�_��w�ǧ~�k����_�Xjc�fIx�W���ұ堳W;���ۮ����P��k�9��i�ϊ��3�p���xp{6��G7�Ua�>����#o��:S��9ˮ���	P�\
7>�]��S7�}�Y�Ԅ����w�7ޓw0�w��8��t{����߯اҶ�̣�S���\P^��	G �O���7ޥ��9�^�[��q5�˻��$���~������~W�/å\Z9����{�C�~)I���d�)�N��Pפ�˦2!㼛ƞx��*��=�!��'�?`���)�b݃ҼJ��#���L�X�3_J��XE6�u�
=��7���)�o�m�\]j�S����CG��h��ӆ$\v0�"ʊj엺7����ǦRw�=*3�2�>3�*�*k3-�e�ս!�u�J�Ǫl��_#8G��m��k-��Щ��
X:N�ٽ׎��ȭ�ʇj�ͭ�u4^�NB������o-K5�@�������%W�t�҉S�/AO vz�y9A��e+2>�lВ�P�Y���`Ozυ�.��7ܖw�H���8����}��E����_���K}4@���62SCƑ\m����Vny�7ϊ���ȝg>O��ր�ǅt���Y���{"��U꥟H�l`4%��yt_��x³ЊĊU\Յap�f�1�'7Y���H�ǅ�fO���wN� �����sb�~}g�Ѳ�{�{��ٿ���on�`�T�k�q��2�k��({ީ��w<�6���
�F��P�zӓ�*�^E��ӝ�����2��{����~���meW����ym7ܔw�$w�=�Z3�
4C]�����:r; �6����͟N��/z�1���z���"��G�r]>���y�灏'v�&Ѻ��^a�5�,�}#��<���X�Iֹ5���˽���_��+��>b�'���R�v�u�
��Ǖ�3����y>�PI�\Vs(M�m)��.��!�n�Y��t�?=���,ks����fa����ռ��c�b7�lM�1O�������>3i�s�A����������v�!Nӵ���[�nA��7xt��`6��z�̛q�{F�C[�+5���ې��I��T���B����1��n�R�CXk%r�@�e]�/-Eڤ�ᵖ�.��s��R����$�����hzD/+v�Z��7�b�uR�ܦ,�&��u����^r���ڎ��>�*v����1j��eӷ`��>/N����̨o���LF+s����Uμ����7�d%�qE%d�[z��
�,y��X�Wê֬���*�˺�]s�n��̶跽�04wlvGNe���A�-VO�0j�+a]��Tj�wZ��� �Epyg�M��q���ⶮ閧Jr���R��z.	9q1^����:+5՟	o�6��Z�K�bR��������C��e%h�)�Yp�����z�-����)��s�u�:��,�7잞�ܧ��9�K|d��D�58d�$,\�J��ٶ��J��������ʐ�9j˶�tR��E:�����k"Ji�n���ZZwk�.��]Ml�+s9޾g�S�L�Au�urܥ\�C����,�z��ԛ���c2�r��|U7��7lk@�kˠznʑ����h�}�^u�3,{�+p=��Ifx�W��/<��d���I�]�
�:(K�- ���{2U��qB�=Q�ة�bŔ9��k�u���j�7t���gg]8H���B���z�k�9b�ӧ,w\�>z5Z�9Lo±�l��v�	���r��*tu��2,-Lz�@;K{j��`��/j�9t*�]Z�����]E2CTA�W��M�[��8�^�E�ǜ�ܵ���N��ۄ��2�4�6`V�t9�r�nN�)��ۮ��7�eV��o!�@�����A1�5\l#�p��(_f�\�j�O�U7Y\�?��v�#�0'�#+�Z�1���e �k��ad�<6��;lʳV5ƬN��!g�M���i[���I�t�1���ˎ�b1�(��Zb9|�Nt�F�Kq_q�q�FE�h��h��G)�ƴ�tR�����(�]luk.����ټӹ��卺qY�B��H�Q���M	�B]R׶_^t��R��|�Nv�]��:��򗋊�6K{�>he������2uw�ۅ�5)�3�������D�8�U����Js�
@q����yvN�b��:~�3�}�4�gw���ڥ��9��&Z��u�Y�*wn��`�61\�:C{	g�ғ8s���hrP���Gsw6�ZaXO
%l�|��9��x�}^��jp��=�%3.A�_k{�}����p �"�jn���v��Ѧ#���޺�}��_�PSz�`��A�v2P�$Ȼ��Έ|�o��wL��;���N� �����#�@�����v)Y]�9��n���]OnFqW2�T�0�)AӶnv�S-,��I��y�}�����rU�&�,E����N B���H�+.�;�
�.8�L(���Tp�Av����\���EL�p��Er)��,��L��) �W;�wIq�8d�*
���
�I�Sr����yOL�TȦP��
)%ƙ�ǜ�Q�h��t���8��ÁD���剹�U�r�\WO�e����"���gr������z�w:��UzePD��iU�z��8���p�6��#�C���+�E�.'9�-(��D�g�Yj�*��*��0�8�j��9uGP�r�[�d�AS9#,����EΡgP�\�E�u��N���t�\�8D�d�#��r,�Ye��Ux����)�bp�d�QE\�,�v�9JQ�ƞڝOjن�aq�[�	h�YI�꣮����K���PW�+7��;<N�>l�f�v�]�i��m�Y-'-���#��~57≃j�ע|��5藓޿��/��C�{~Y}�����j%��Tz��	��)�>�=@\ER�sTe�]W�Fw4�Uˋ��W������}�؞��Bs:
���z��ü��8g�+H���23�$�Nf�y9J׆�ۦ1㼛ƽ��'��jz�=�^�k�y椫��ӏ�ޏy�x�u�!-T5|��	� �f���C~����h�57��O�x��g��{&����N�����+��ւ��<��š1>R!���ض=�1dUz���Aj%@|Fo��࡞>Y����:���zԐ$W�B9#�/�\�Q'��b�.�i꺾}�}ϻ����ײ= �{\�q!�7!�cc�i�q�7�2��g��*+=P��=�^�eekk=�^�Đ$'Jm,����S���Spq���� <z������\��Z����Je�ϡV0&��W�<�M��S��s����[#�����p߾�.�_u�=�+v�5���� ��Ji@��dc�&��.)�Ξ�^�k�6�O��H��Ԏ�>#0����\������5�ϼaB�C(z��G_3�$t��g
�:��S��N�y�뫍c|�˥�DF�	�GzM�v��uI���vޜrM�J`6&��s�K�y.��`�ջ�[�9<vt�Ѳ^I΢�_b)���vQ����IE_���$�*u���KޯL��{ӓ�}�R.xq;P���_��
0�Yto����R%Ez���y��}�7=;�w~#~��
{��d{�y9�ͺ���މ+���]zB�k�d(�ǽki�+qz��}�4=�h\��8��W��w�l� ��d����]̀;S&/���N_�:}���:�����x2Ӊ��yاV�<xo������+`�N�,�3�%���o�r0��/a-m~f/�~�S�Y�=#���}�_���7�{�eP�!Wu�����.�#0x�9ؐC��� m԰�W)�?-�{n����h��;�߷�Uc�"}�M�����-������E��Hd``"��V�>���a{�u�-п;�Sߚ|ۉ��W��s��߳��G�5��b|s��>#b����r�� +�T8��Ϛ\G�-;櫖���z,Wp;s"�ǌ�[�~���w�lO�ȏr��ϝۗ�0�|�Xs�Wa�9fh׾��k��# �l=f�J��"�^���U��x=���8��C�*�!l�没�.�,f;��kj�U`2U�/]s�[Xp��f�|�jQ�Y�T�L�:�5�f��Z��n���p���ʻ�;E؃��
��dv�ץ�A��7���p�ڒI2�N�򬗒<F��c�Z�7��a'f�p�6Ug�E~�U!���=u�QMّ�S�s�G �V�lC�cb7��<ƈ�n\"�8�U�p�I(�*�w�v�M������6&�����!c��z�O�<V	=�^����s;~��|�J@��I�c�z������m㸫B��U�4t@f�c�)�V��e���G����B��<��*r!�fT�n������D���+W%�S=�W�כ�(u��[�}m$����e4��r{oҟ�����g���#�����>۩��/��}
�R��f-���+*|����ղ�,�p��dy���ӛ���f���3�����L�_���=�����>�{k�x_�6�����y{~�Ŗ�o~�G�)���k~�>�иLU}7#pU��yGc�����g�~�!����]5��/�9+��s�e~�wP�߯�
�6S\e�t�E��{�M��sP�]T;R5rWs��T����ھN�|��ڐ�C��{�e��I�R�Km�S���zF��߂طjx��+�]�`�	`�z$��1ϰmL�rhP�o��wU֧�R�s�DK��]S��͍Lݻ��^Q0�)����V� 4J�2�M�������Xm'ti���j�"׺_%`��VF-�(�w3s�-��K������zXk���7��y�9�.�����74쭳��{,c�"|��O������j7o�&�ad�	��[���s�^�>���̣�Sݔ�eF�5,@�>>es�C�ǅm��$a�q4�C/2ğ_�o�v��9ʶ/��(eW�\����̱��n���cQR�������U۪n�;�.��x�&�#����C���=QsT���[:�}H��2G�3�p)��J��XE6�9g�c��Sy��)��4�]J�sGr��3��,n_�yP�7����bNPb�	��L���@^u��+�3��G�ɓ�}��+	iE߲vz�Z�G��zO{ֈ�dV)���*��A�~y��ڀ��'^����qB	���i��+>eh�9���z��
����39�dU��U,�-����T���`뭌�=�X�W+�������K#��������{Ԥ{�Nfy��雇��RJ<��T���^Q�O��h>�Z����&�o7/��T�Ϛ�d{_�e�O�P���s'ֻ{4��g�ez�F֛*g�>�7*���\�''ղ��p���g=7����T���"�V�ɳ�7Q �:3>br�(��i��8A��sy�D1E�RU�� �m4�ek�t�K�q��&���u�P�{WQ͝u���`ԤLYZ�k/��v����]�����/_[�T�/k��@����u�)�܂�#�B7��|�}95�i�TLZ�3Q�ևm-O\M���iӗ�v���x����H8�v	��'Jq|��C�����!�j��<J�Y�>>>�����G�*�K�i�(͏9��#~;��'����B��t���6�FGK*��
C^��?�T\���zZ�C.w���rQC�F��37�Y��{�J=�>W�'��#jr;v�w!S� T=��#g��|��#��%�Q�q~�wl`�l�O[��\�	�T[���5��mٔ�֥}ʺ��<�s&��� �/�GE��p��whd�D���k�/"{��1�^7����dq�}')�W L�v(��(��[Cӑ��>��u^U�:�}y/d��#�C��3��;~������Y�JG��YY[+H��B���O�sAR�P�n��x�&��*e��k�����G��{%ϡ�V��#�y%O�v-j��Km>$Ԍ�ow^]#}6:�^8��L�y�R~��Ggi��^����y�+{�Mp�n��ӔS1>]�ī�/�}F��$�u_�֤�7�G���<.
�>Y��-R�א��Z�F��$�޻sVꃡ�x��b܏���IW�s���2g	3�U�m͢/��Tǹ�"8-�@5OՓ�XɊZs3�b��Ʌ9�L��l'���#{YU�B�jv�Ȏ�m���%C?���� �_P��h=MZ��]vf�J-���un�-�C}d�)�^��;����C��̏i���� m~����22�!�sQ�&T�o��؏Uq��F�F|��34��Q[Bz�p|z�G~���`�|��Ld���'~�z��,����!O�<T�����z���]��UCo��gs���6�$�����7�@M� ��P��&�n)��ȍ�h�J�׬O�U7�7>����)% {(G�%��G|�>�z��?�4�j�R�}(`|�:z�{��s��8��1~�]�����=w�����S�k�Ϫ�ޯL���9'�U#�׀W���p����Ac����:���n��1��L���OKӛ����_�X���l�=��Y�S����w=9�[�w�����
#�jǢ��V�Bh{@�x?iŞ��w�[��c���g��{ћu~/5f�`%�)^t���p�U���j|ߒ� *|��G�)կ�~��A(�7����1����<�Th�.}|���mWJ�7��s�5FV]z�Nw>U�:��Ȟy��KTڜ��{w�R��hr=o�-�,�>������<R��"�s�u^C;��s�,L�Ѕ���p���^��������{��\�Z�DnPf�M�P�IA�֮�%~��!���E��ɰ6���ã�f���m�� {�
�\��:�1���Tf��At��+��gbֺ������x��o6|ڦ�D��㇣t�\P���ȟG�}~��z߂ؿZ�)Dt#�Hf 2!�h�niO������������{������e��g�&Ŀ{:w�k��B}���|��A�(�����VQ��#�y-�TO�=�܋�=��2)�x�E㷞���s��3�r��uN^��i�X��fg����W*5��S� �Lϝ\P35>��FM����6yd^}��$6Wx";ޡ�)j{��0]��;޵{�D����dU��B�(+��bj��#��繊(c*ԭ�~��K�M��.���k��2��C�D{��>�߅M���º��$ؚ���X�x�b�>�}�W�=���Z�ݶΖ���O���.v=^X<7�]���c��8�5�[�����B�S�M)�W��p�TW�e_��K�'�}9�2�>m߀���^�>ߥ�t���eH��0ȩdb���O�71���8��>�Qw�7������G�ƽ����yC5��}^��g��K��>ʩ����˼�wc�U{�0�B�bxd��w�3���@��=9�[�a�s>��o��t9�q�u�O;�[5��R���2��"���ǽ��I�Ie�tJ�����V�;�^��<>V�\��R{3&�]���k���b���ٗӋ�q<��v���6�TC_�LD�y��v��u�<��o��-��ۿeKY��Dr[]	����aT�ҏqrM�:t�}�/���[���m9Y=].��;�,�@#x���8�=�S��f_`�)]��sŬ�z;�Y�~�q��1Z3�<:�"��������[c� Z��r4�J,t�fc��[�R�$m7�G��}���?yaB;1(g%�^�A~��t�8}��q�f+ǽ�$�(�s6c��}�ؼ*v��zF�_��-�v����js�]�<Y*�ޑ�XZw��z�EN/�n��=��|�$��,�u���ԥ�}~�>��[fm��-�T��l�Y�ϯ-'�j�G֒����'��	���O�gL��}~��C���p�iߝ�TW������d�3�{6I�J;�w�0�F@��KW>���ӫr��㼛�i������;���4�p今�a��G���D���3�b��J��YSa�����z�ک���i�5���e,�E���/��#��C����g޻bNPb�	��L�[4$���\P�+����Ӟ�� ���Nx��T�;��;�㞓�Z[���@qɮQ����B���Q{�����]��"�P��ʆ���1^�y�ޢF����]�eܛ�S]AJ��>��\�i���t����N�
��:92P.�N�6�Ķ�٩w#�1pUhi��N��܏���ᕜ�"�{,�5�̼R���m�����]��9-�֦�B�O���%Y��������x��&r��;���=�> �?z�ϯ���Q͘��#��|������P��m�V=;\NC�~sQ�!5���z��?�̟9����2>�/v��sp�%)>��D2CB���鼍�^ƥL���d{Z����O�P^�n.�#�n�,m��>��s'a�O���U#��@�Rr}[/.����s�{���nC���yf�yw����ŵ��|���!q�T=��D��?g`3����
4CQ���׸t�,v@;�*\lUŕ7fp�/r��IC=S~�g3gӱ�_��?T��?��$,�gNK�����t�������ey.�gGyv>K;�|,�H�s3y�Y��w��
�zσ����7�ڜ�ݺ�A���>����D鵻��z�#�(x{�/n�d�x���\Չ?R��
u��n̥�>��J�aRڸ�V[��Qf�b-�8_�F*���zn���88�逐,k���aY�FRsX?Tί�m��rnl\�����l��;��T 7�R�sTe�U�:g�r����O�K~����}$J;I~bUհ�M��,-"�&RV��#G��
���:�����M�ig_
�P3�|�p���9��O7��.fXU
�6���� ��d���mӵr�s��]]����p:�V�9Բj���	B6%�ҳ�ϣsouRu�F�TZz��ݧ�9�R����y�~�<�-�V�he'�9"��O��\hC�ߖ̷�LW	�{>9r���o�=K��xͮ�S�Ｇ���ǁ��ǹ
�y9A�< W��D���Q��r2��=��z�R=�+�����3s���:w�ߘ]�c���Z����ϧ(1p���m�����m���V�.�TO���3�U/wC|�-z��N����޵$�z�NG���Ү3ӻz2kk�>�Tk��u�2�Ir+�̌"��5��T���ccb=U�{þ���EEn��x�/+�M�=�,Z�#�@40]~c>�hME?Z�Ŗ�2{�)�x����k=C�^�Q��������}W씥rUiwܢɁ�y#��2�ߴ�Q���\�ێ��[#��3E��f�6����I̡������OyDK�迍zSJ�K ��}(P}�6jr���].����TP��~�zܖ��\��?fT�\����|��' �n�\�
�j6R"�r��(��qY�b*��S#ˠ���ϴ��[���s�O~�f�##�����V&UU�����S��*do r�ƈ�2*t~���%W.4��o�Sn�En�Zٸ�ȹRn�ը��ʼ�!SJĕӏ|�q#�ػ�nE=��d�!7H��N�I������G��d����޼��-[���A|އ[�L�V-Z���"���2���X�%d��n�������wN�-��&S��:7Wb�{N��fjn��ӶvP��r4����b]@%*ot]J	}��s��*wv���q���J[��V"����5K��b���F�e7Wa�v�Y�_gVk���*mA��q4�,T,�g-�J��AdS�1�8Ν�P{3o�'��cR����hv���B��M�XQt�0�/Z�v�o2��yG���S��i�%^���Y�gn���d���Q��\��Z���԰���q2�*D��.���[s��G%2����f���8;����6k��!��+,��(�J�L ��K���?R�d#9���*�Ա�����ۇ!VjGYd�C72��X;�]C؛�����LvNk@�Y��f���27��eM���.<2u�Ae�`]Dy��M����۶�KG1a��F����I1R�EW_L�U���E�4�u3HL:�L�d}��Z�;���ӽG����c6C�%��H
�E���e�vi�[W-Av���բ���Nڕk���_d�b%���>�q���˜2mGY�q�J���4���a�O7��~�S��\���kM�4�)=0�g^7:Ɲ���Im)u��k�-�
�\V��e��/c��I�v�	��9r�i�!���j;�mbtk�%4�(M��� �j,���5�Փ��l���6����6cS|�2ܺ(ժG(B�L�@N����}���Œ��Rܫܘ��;6ly�9�C6�89ĦS�.�V�:�^G>��/7�J��LM�z@�V{�������G��٭�4:ϻy#yh�`sk���Ar㜬�����>�yu�u�o��۽۩� ��1� C�/-�*���1�r�w9ʘ��}�\*�q�s�l�}ph9�	B��設b�&�F��mҼ�}����ۀ��Yk��*&�⹕[��.��m�z|2��G,��zMw��ѹk�lE�������^�bV�8�S�u�sH��#��:��O�9���C��p��
Z[�;gf.6��{�Q+����69�-����ǽ'.6o�m)�;���M�;�B)k=vڦV�]q����WI�&Լ����.����̘�P�O6��r�5��
��z1�|�]Y1sB������K��6���p�N׃P�ZT޹�1��B�*&ֻ�R�PڕhH����b��1aչ�]&��ݗ5�Z�u�����5u��|�SO{+D@�XXbR�V�0R=չ���(w*/�1����9���V��Q��EP��%��"\��,�z*8w�&+��X�w�B��m��$Q1�Kę�^2*���DN���C��
�@�eY�\:w2�Z�PN\vꎜ"
.�%]�*�0�#�ys���N4����P�B�J���<y�Tr�*����:K�6�9�&!�H��(��4�N�Q8�^��QS�W0�+��QȬ�h��BU�TN���Zq<��霪�
�Zr��fd��5f�r���t%KE�8��a帮^0��xÞ2%ˎQDrex&�`W�(�ӝ�$�]CJl���t����V[�GG\�.RK.��3���(��n3�H�9EE�ˑh�9<�����eAh�JJ��	S�.G�s��.�)V�!�"�zx;��x��-s���T�n�u.Y:��%�z�J�C+�H�R�r�<�J��V*���ʙ�R���jV,M��7��]��٨�@�Vmj�YOen�ӽ=i-vq'Ҭ����\��w��3�����;w��ˎg���KphHӭ��O����ϴ��Nӻ��7q�V�yp�v��v������gR��t����aT���Ms�Λ�j������.����:���$�z�M<��S�����w�V<�}�
���6���q���:����k�0_���ܰ��;%�B��sbǞ]�Q���X�H[M�#��~m��;�ab3�[tF`�	`�;H���y7��"��=��v
^�����ejJ'}6;�$�Jߧ�~�/�����[�[~�>[�"ʤ; �P���Dz��-��u��ع�O�����f\W����g��t�׼;Ƅ����|@�e�����;"�����znɿF��G� |*M��ϬW�[��ȯx�E���{��u������+�෌�����V��}�\���{�0���̟U�3R��FM���ICa�E��i��B.{]���U��zY*s���I���+��Hb�	A]zĆ���"����2�J��q`���վ��sE)ۂ<��/�U��Dz�¦�Pb��7�I�5AyU�,v�7j_���V�~�y��Σ�I���M\z	�%�Jy��0����7�
��������ss9��.q�R%\�NL�����<���[�SSk%�F��ׯsθ�Xe��]M�D���&v�A�wSR�povnI���rn���iU'j�`�h��3|��m�z8$�?,����y`���Wx�<wqS�r&��飢�=����w=�<������<�M_�9�'�}9�2�"w�=���y3oٕ"�S �߸ߦ���%��h�K܍�>������ὔ�7��!��{�Ӱ��(k�L��{��=���g�/�Ug����:��!\���{�#�Z��dN��~�}�;)��:
�Fi��z߳�~��P�^���Rgu^�J;�F��'<=�[���'C��=]/"��=�-��4�24���>�C�шN�!��d��!cք1\��f@Y��M7�ߊ�|�����b(=5��t_?��+�x���b¶w��Hw�g�]�N׭{}#��_x-�z�x�yaB3�ݺ�0;�Cۚ�{�y�nmm{՞n9^�+7ŏ@�����s%w�xT�������O����r�.|^���/����U�fM�J}
ćP}�hd���웹������u��g�Ϟ�~�>���d�^U�*�+��w�ƴ�g�s�^ x_�Cر^C �8�cy��������}����4*Q��pz���3&�A=����P^:;Y�	U.���vӋ�l��ڮ1+6�\�ņ�lF�5׃�Ӳ9�
D-���v��U���e��逝Q�$�cG:Z��S��:�+��6�6��/���w%��C�Jm�4�D͂���s��X{j��`@��D���Rü��y�]/�0_ʽ ���tu�?-˦1㼛Ϛy�=r{������'5�E�C !��)��] �+T��|Hտ'C����	�O�Еaצr��}��̝��r��~��c��{�l�T8,���g��&Z� hD��	��˻=o3zdTp�͟�)H����Y��R�c��v=\s�{޴@�z�_�)�)�����ݏ?nj����h��K=@G�+={c=�|<y����eh�8ߞ9�W���º||��39��E��L�`��~,�Z|���[�T�2�5ͻ��hԲ�G������P���jG�</�2|��'] ^����,D�S/�|��
��H7���V��S7�{t�:�!�m{�=���(
���uW��މ�{d���u�`P�{�̗��O�H��^:���n���Mt0G���d%�Y�Z�9	�x�:�E_z�]/C�K0����P��W�A~��g�*V��-�1�>7zD?�Y^띸����3IYK����S��ә�����cy����}גG{:r]�V��ڼ�NXK;��G���y���`�9w�}u@�яV�*�Y��
{`l\5�X(�:����d�5v��&���!x�!����F�A36P�+��I��P�`��ٽ&��{����B]�.s:��y�e�m8����݇Q�x�NH]��}��q~�
����f��|�zfn3���z��g������mNv������i�Cx�_*þU� �Q��WǼ��D����~'�����s!Ң���q�ֶ�ʹ�qt��w>������ϧ���=�e ��7/�hg�)�����'�~���X=bJ���H�'�P�2������:FP��� �)��5F^]W�FDw4�U�u�v�Lj-����+;Ū����\7ާ����
�-�����)���<����Z�e�m?�W9K�\���V=�דx���g�}NuǍ�������- ��2�w�j������Z��-}��^��W���f��gO�W�.<�pY�S\2!۸y�5}��8�Z����FD(�� a�l>(3�qk��vu��{֤���]Ir�Ũ���<ɏ:N�2}�^�T[2�\Bk�ň�"��bࡌ��9�H��^��W��{�=�IFw�����[Ψ��ltBk�~�7�-�d�!O�#�M�0��wTN_���/y�\��6����v�aw�=�u�������v;$yu�H=�RWX�//�Lcy�]�EҲ;r���kE.��	�
��cW�
�T��D�wy�I鷸���T%TY�D�	oK
x�2*�3�++�P��\��Ll��GsrH��wש$�m.����Uw���}3p���\*�zd�:>9��j0��=�NTɯvx�x�^x=�&ħ�wB6���?W�O��l���jȚ�����)�j�2������V�J���}�v���7�9�Y�.u?fT�\��=���>y�r}�R�ا&�ec����zy�R}}5�!Ү��)���VzL�����������|)��$p0�ד>w?M>[��/a��S]�)G�.��_����Οڳ�C�J���)�8�ӿS�� �F�X����v����Q����v��em�5�;"�>/b�쌁t��Ę]���^�Rn{2�og�"���}f���<�����Ġ����|/BZ:���t_���z��z�0(����w�QHw�ez%��Z���?�����ab29m�<Y�;q"�s�Y<�L*��]����펭/�����g\��.�^����'O������_�O��
�"�ۤ3 ���ȓ�z����Zܙ���q�ߎca�QIZ˘*_��;��׼;|lO�{���lVѕ�1���ކc+ò鞙���ȭ���y�s�����YV!�,�[yt_b���}e*��z.�n��v�n)U�;��E��Y��.��v>9ʑ��/�{�D������<��efc�JJp��'3+��je9')7"5���Rh<�����ԾIl����B}�vb�g�{&/���:tv<lO����]��7-���z��P���_�`��S3�W�Kw�Ca���!��,��z�f���8�^5�v6�^n�'IC^`�=T8,���n~q��6W(B:�|џ>�¤b�������K_��ovWp��^8KJ*���6q�o�8�Q�1�� �޻�uA��u�I�5�\�o���E������������C���NCk=.w���}U���D��qWS�rj�{|��a>@ق��j�LG�����j��O�������eKn��!��q�)�Ԇ�V�u;�����Z��H��2m�&�G}�^`����m��?;���3��{=2G���
��M{wV��i¤O�~�Ɓ~_���o�_��*Z��!�L�ӛ������\�T��2�NXe���qj�zg�z=�p;���#�U�i�B�ӕ�=]/>��Od,�@#c�?e�p���l���*����2���Fz������Y�|}�g߿g��h�Cë�*��A�k�E�;���g��em�B��A�Lч�vz�*���Jz.[�(U=�	�=�G��}�V$(<QYt�T1��;�Q�@�N���rl��*���Qť<�nJq2{ҳAS���By��|�n��7�!�u҉Z�ܩ)Vvsc��}eJʝݮ7/���2��A�7�Z�������k���_��ǽy<|���̪А`w`�z|[��[�1�1�ī��>�V�72��O[��\�xT�[^�Hؿ[�[�O����.�"~���v�}?+]��YxR�ȍ��nZ�C 㹖�$��,�u���ў�>{�S�W��,�����8F��q�-rQ�3�/n���Q qA�X�p�G�6M0�e�Cؓ��<=���p����՛��Y�JG��UƜ�}[fVD�\*��9���yuMקan]1����75�˭�ono�W��f����sܲ߅k>��Q3>])��ҩxV|E6��7.�U幊TrD�*���8mM����-�cC��pY��@���lC��(��� T�9~�$����D�KRJ��,�[�
2�!�b�;����ޮ9�>�G��G���1A���O�����M�W�_T9���M "�����9^CǢ�/!��L�7�v=^��<+��?z�eg���Z�+d�@�&��UF���*R Б�^��4:�BY���G&o�=���R=s��{ph��n��O�6� �҅@Nμ�8ڃr���N�Ftu�[��U��=ӻ=I{;��=;�U�X�Q���F)�h䭻�|:���֧N�[[5�+���c��k�n�VJ�%qɻ���0"����h/ymn乖��e@2��7���|юI(��ݵ�����&��3p*��|l�3}7��k���J�׻#ݜ@�q�����J6�IH��Ԑ1��2}�����eP"5�iI��l��\:r;�M�~|s����;�1�(g�Ǚ��:�����P��z$��;�`�G�Q�螾�\پ`�
��{�J䭞}�V@;o��ә��n����O��^HY�Μ�y�Z:X��9̭��<���Wˎ�נT�;׶��u�7�s3y�Y��{�^�sнy<FǑ�5��4:�r��l���䔣����We�^��h��%�n8�y��J�t)�c�ۙxLp��3��x��f���=���Ch^OeS�|(�,�/�ha�q>cA�D�����ٿsY���T��+�)U��=�a��o�#�ǥ�f�F�I��\?:	h�'�*�[~sN�p���gٛ�w�P���fԌ�u�p߽�~b/�#�`V� tR���!���;Z�'DU_�}K���{�U��̪���z�m�_��yO��x����<�N�C�kT{W�-�+�<9P`�|.'0�m��Vd��i�B����]��M�+���`�S�5⺍�H8l��J����,�\�%������>�κ�y�^�p�s��5��A�\��ڳ]�8NYy҂ 4�b�+@�wz��k�z7	��zKj���Nd����O�Δ��3��%��N�+��{L����߼����V8,�u����׵���������H��,z8LO���15<쁆�x>sQ�/��,��_���]~@��jH��
��5χ�v�j����T��vf��AU�3-ՏP���� �h{ST�q�����"�r���>�%�`:=�7�3�{�f|/º!� ��M���S���t�����.6/jD���ц�f���+'��s�>����ڗʾn�K��ɏs�HƮX�67����:>9W;�suw��M�J��,�>�/X�?+�a��2!��}�K��^�@ZN�3���)�_t㥇<Vzȁ�og݊�E�rr��s��2�5���Y�W�A�=���>۩�:'�Ofʽ�8����%CP���ݡ�t]�/�<�
�I��9���n��o��s�Oc�� �ۆQһ���ȇ�R��)��v�w#��W*�r�����Qk�*V7|�Vb�N�;�p*���z�^�X�I��-���f��;
Z��*�ϗRa|�􈨌R=�-T��8 �Y7���q �`H�^ِ�s� �T����*.�(q�[��d'd��n���n2w�<� .H�ͣ/yEA&�7�nܣ"�a;)�:���<Y+w�8�j�8��������۶8T)NǝN�0�����	�u��9��c��oG !���b��W�D_����<���^M�WO|�C� �6&��Ϯ�c�_���ȧ��-rQX�����=���xzEz��Qmdq�{�rۢ3�,�Nv���c�W�uʗ"���41�b��{'ג�^�)���=���^�>*ip��!������t�h��vz�y(� /£X�^�4C�9��!bܘ[>����G�5��b|s�{���a����7M` fׅw�<��S�3� e�Q�X����2���㗓��GK9��{��u�8��3A	��j�z.Fg�㯊�𖇡%u=�.&�IT��P�3פ����o$��<�-.�/�}���q>W>�uZB#��pY��	��[q�C�J
��&����2���]¨��کʌǞ/����pz6�:��!���c��G��~�@>���uA�B�6'�D�t&�f���R�o:���e���{���|��K�+=U���D�<wp�97�ǈ�`�ʲ����9�����g��onz<=U!�\2�K�N�M�	+`=b���W3�>�#cm�����6���1���m�m��m�m�m�cm�M������m�o��m�o�m�m���l��m�m��m�m�ɶ�1���l�F�`���m�m���l���l���l����1��&�`�����`����l��b��L���N��O4� � ���fO� Ċ�� �ADT�]��*���Um���%UPI))*��)UIb�%A*��$�)"֊IP��!�M3a����5������[RkVem�,l�ɲ}�vl�U�mZ��m��Y�6�*���e��:�j6f�C�#*�,QIV���%��kT��v����U��I��U�ͱ�kmU�UfZƃi�,$m5Z�f�΢Ͷ��T���V�[6��JbQ�m��(��6m�jA����ݛj2�z֥m�л��  7�+�K�\:�r�@:����=�����[i���U=�s�\��Wu^�:��w���=ٽ�TT�^/{ 5�r=z�S�Vr[�WT��̶�i�el�QAfY�o� 7x��R�{=^ҭ���9�\�F��ފk��,z(��(��DwmƎ�4h����������F�QGϫ�Q@ P=��ǣ袊(�F��ӎ�
  (ދ�ɖj^۶ն����Z;x  <�� >�=ݮ�n�uGKn��頷�����u����(νp�or�ν^=(����W=���뫷g��=ڊ����T��U�{m{b���+n�vY��  }�B'�S�����z��3�wCZ m)��P���ǧJkm�{����h�5˝���\�=�^��]!�v�bM ��ZŶ��'mhk�=�u�  o}��k�����Ӷ�lܞ�u��v���;�F��d���kӶ�^;�FJW�O#�*[\��4�m��ב�E�:�un�1�=Z�&��i����Z��s����  o5���n�/y<z@{Ƚ���[S�r�U��G�q��j�t����GGF��s�צ�+U���ҁC������Y)[�`*n�X޳J�N�����h��*��k�  �^��47m�����b��׳p�QM-װ����5�,�v��C�EMǧw�ݻcZ:gw�x=w���'{��B��]ԫi;�R֋u.%ݸ��z�IS6�� 3aj�2T֛�  >��a��U��:ӡ��}�OyB��]��{xz��P3��ݳ�A�u^�U]Ygx�zU:�۱9T(h/#��U�Y�˚{�w��m���E6�B���յ�[m+M��  .��5�����w���5U�lN�j:uа;t�Q@Ӵîn��I���=)/Mokkz�=������M:�%n�g@�L�i�-��)CN����K3�9���Ѥ�L�  �{�Y�K�V���4z�������U,�ή��*л�����z=¯j)B��sאhPw�{��.����omx׫m:��Cuwn��K_ 5O�Lʤ�A�� Oh�JRP S�dOUT�a  S�A)U��O�jzj����� �%0eT(L�x���?�������G�����w��Dϲ<�t^7<���u�޺���g]{�;��AQw�� ���QS�AQ�D��* �� (����k��fg��xw�k���,c�S�>ʚol�2�8eB���M�f=�L'�Z�g�鋺@Ȇ��-�u�ӂ�#���ɣ�,��Ԩ`��63*T��{�,m�Ǎ��y��|��Tj��N�[Q��Y�J�b:[�<�)�J ���M]ʙ��d���;�2��jf��⁍�KVՕgtF#v��XԨ��f����0�8��Z� G�Q�g:��jڡ��Z�͓r�t=�6�6e���[����B��q���0 ��횔�2�V5�<5iȕ$1Px˦p�����:�;������0	�˖�r�x_b��4�D���Ў|���� έ�7s�"v�,7un�c�ƢtY�����n�ݽ��,B�c��ݼԞ�;J5t����5LCVli{ne��; �Y��!���-f��5D���Qۓ�C�t�z�A��u̔n�N^� 7�l�(�vbւ�i[�2��ڋv��%���U��ŭ֩�Hif��1�[T�aR\���W4��冖�[��m�ʖ!�*��h���Y�CHa�Ʉ(��{&Z�|+T�֠y��*aY����W�iӣ��^F�+D��,֋���^KK${BB���z�.�ѷE��vְ�=45���*Y��Of�U����܍�࠘�D�;&��r"pEn�Z�T4[�J�kk*��K�ա�'zk6�͔U�,a���R�X��*ur����<�!S���"W�T�3Nj��8��B
LJ�e'%�ķk%�E+�M���vaB͢�+�+��v+E�PAL�v0eo�#���YF�{ZImm7�����ƪC.�]�GX�V�6)/��{.�[�鄐e�Dn�M�	̨SR+l�VW̼E��[U 1f�wp[ՃZ��eZ��mc�XD�bL%p�P-�n�:���4�{��+��B�b�n�ӎ�۬{HH郎�:j�����$�MV�ܔ����;��OP7��G���ev7u�cb�{I��'�g��F7�N�s-��uF&�K�[����Vr�J!oh�h�P�Zr�B�l)��Zr����J!���ɤ+�jywYq$����yZ6��LQ�,Ke�4j�5(kߕ�+Ղ�:�d��v���4lq� R��/ �7Bv�n|����dX^7��~ÚQ��UZ��1bj�[��3V�,�R��J�)Wi-d^']�%jw(\��,kX`e�%��͆�t���:�3H�%��R�C��7i[ň*UӬ�c^�n\:��V�(��耞d��N<)Q��dO1 ,;��)$hw`kVfZ
��$5�l�#h���7A��V�w�T��^�B-6��L�p����f�g�I̬���Y�VC�gCV���Bሃ�eF+4�6��
w4�OI�y��`d���:.�P�gub�S]H�Q�6ށ% u-v�L����bd�vr�S`��x�/�r�����sl9OC��N��N��Qp�5_m!�:���MEjڗ-�,�7�[b�: �7(�ͺ&�%2T��]���p���M��VX��r�
Ё�$68J~��yR���8e�C�O��.�1J�VU�]IX���Ӛc0$,;����f�ګ��ˀ�AZ9l�ߖY�CS����C���`�P��B`�6�=e^�j[)^݂�;%�g�B�a�t�������#[l�%�]wrR��eU����. �y�n旹�$&;��	�n}�����@��J��Glِ�S��I��Mm�'�Vm�B�2��
g%A�mܰm�v�뫡���HQyW�$��3� ���� ��3pYLPF�Ym
(�e��%Zu�Mҍ�u�Í�ŕ��y[eR�������TÊ���ge�����969�D;���H�������A9L]���v����r�(��BPp,���`�3#�0���x����wT,bu�(+n�v�)��Ys)�إ���A��բ���m�W����
�@+s��0�� v��*��a��5�ܔ�Cbv%��ɪa�QR�V��]\/\���6��J����~PZQ�0\��Z���(V��V��s��R)��v�E2$���l�Swd3S^���{��P���wْ��d���:f����XN�h�QL�J��R���Y����WWu�n�5C",�ʻr��`�h wh]��Wre�eP�Z�F�Xu��t)+h%Sm��b�����/�Z��U�X�������&t���(�˨C;�\�q���/X{)1��v�Q���.[6���͆��ì�:���y"K2`s�(4/4T�	ݪ�I��]ʷ��I�4�c���vfV�;c�[�0����P�/UD�-(fh��W�ޥ�V+t�.=��]ʽ�=�$�5�E*����p*9�=T4*���a,Ŷ&�����f�:�Ķ�67��R!#Vo*��f�j
���e�.����%�� ��P�l��ո���#᠅t᫷%;͑d�(�b7d�ŉN	�6[�aF<�/�toQ��Am\�+o[͎�&THP6��u��f�J��*͖JP�D��9m�S�4���e�Yv���Љ� ���v�D�Z�0���y��u(H�kwK�U�<
������1;A��	w��ijۧyN�],k�c3QP�li����
3m��`���l%�sS��[�C3p�U�u
r��z�xkv@:l�ZH��`�/�ض��eVM�Q�l�u���0ݐ.��aŵ23� �$(&�yI�Q�%��#mI&e0�p�����1OVĀ^J0o���B�	���FT�%��˛ea�s!�X�B�.�@^XlÅ�M	B�D�YQn�ۚ�*&G�ml�g˦h�����S��7�+�Ȩ�yn���7x�7+MH�7��Kg%�%�Y�����s�����[J��"c:r�:���j�@oR��t��7sN��b]�l`��T�B�1��7�KTv�÷GN꽤
Q%B����A�S;�`�6
& �RKҬ�X�m̉��OV�"���ِ��@i�,�d��lf���[Y��"?-�[������7<a+�K�YX�Bv���K(rwKL��9�ع��
�-��TM�%�ض�K_m_�Nl�C�,f�i�i,SR��V�1��Yz!i���X�.�ͽ5�˘����Qj�[�h���V^�T�oItþg�e�Ix�����5���۷�,��_H��n	[������1�[N�X�_�2���U�A��/]��A�z-fn��@c�q�`�TGoEu5Hт��[��ņr�8��	
X	���6��T��׀�˕*ؖ\L}�S���"-$��)VL`8�ݻ�PG()��L�Y��nh�e�C%�Gh�tBm���#%�����S��q4��x�l��J����j�mBᫍ���-g�W�V���˧!ZVb�{V!L��£�2��N}��Ȭ]���ݰoK{GHie��0I���q&M��@�lS�x2�lf��c�Z�x�c{m+�ȱ�S�`�T�*�K��mO��Q��	S�.�Z�&Y�0�t��iK-fQ�$5VjX�y�ّ��]1bh�X����m恔pSxc]�Qm�嬲 d��r�ְ�lò�CX��i�T�xS.�{��ihX����Ѫ��j4�.ɶ�'ymL��F�(h�U�X��3���/�H�54�'��/%0��X�R�H�X�`x��
�3�gܻzN�
�RM�{��4����Xʲ��1�%֗X��^H��N<8��t�� Z/+�s);��3]f���QN��$.��V,3Y"d�4�Ƿ����+�x��m���I�,�̦�D�edF��+�R�%���
�a�Ye:s%h�.������h��j�f6�T]���Z�D�Ғ�	(n��x�j�3XV�m,eق���mU�wB��F^@�l8R�0V���%mk�9X�XCW�j�@
S7Q��Qw�F���E������I�qC�6��9fA��u.�t����JA2�8�Z�m��3�U���|.�MfjF��Q�LR� �N�ES��Ϟh	;i�o�)L�6ƫn�K܂7vmCn�M������e�Y�!��<j6@B�!Y��+r�YX���O�V�	���wK#U
(���L^S�oռb�f�ޅ�Id�oKE��*�mD�!�f��˘�9v@��O^�9B�*@L��$���	�.i2��F��4V�-	���I�Z��@��NAh
a�e�Z�ڶ7�xn`߬嗍�h��϶���֍��H��Ue'tI�����($����nS���ck%2Z%}U���l���5�=���Yt��.����a`�bߖV�]�%A8l<�F��d����j�
dh��t�,d�e=*�eP<@���n�u�C(a���V��h��6�e(yOlV����u5�b�h�m�ٚ�rav��u�1�ɕ�UI�V���U��+��*�FI��X-�b	*�E��l#��q�Y*�ɵ���mdr��X�t�t���͈*��RB��(���m5u� �)�oB��]%�ϩ:�ؤZj%.@�{9O�.������,L�r�k̉��gu	��{���ݺ�s5(���f��NkN�`�9�B�(�NV�vq����������ʑRնhS �xѺ��r)(� ��K^:J��w�h����wH��ռjZ��� $`V:ZX���#Z��.���T��1�ysM�h�F֓�~Ø�&PCTg�ױ8���ehؕ--ڴK��6��Z����k@4����L�&hn�F���r�M�h�i�TU�A��ΊZǫ�uu�7��!�[�$�����1��HĪ�K�(S���5{y�gZU��`J��Xo2�hڇ!8�P��m �����Z�������"�����U�ThS�f,�*��kS/^����7�+�[$�Z�̹E��:F7k���iVi1����ʀiyEЭ�m4��;��T��aς�E
����5bFӳoַ)�-سqCr^[M�o�+�*���;ZZ��ƚQ�A����áh �[���3m��,�3+�N�@�B�J�	�(��A�^�YxڐbYv!@&��/�И��j-�m&¬;��Qa��hƦٛz�3{��mVзn��
SU�(�U��ͣ���n��n*X.XlP8*�w�u搐d�:�jGQ�g��|��Ϋ)a����gD�������c��A�%�AK��L���mnZ;n�Ëf���a&�ӹ�g��i���R�G)��#X�Kt��v�V��B��8��"���X�v��*���*�+�<��T�BT6�n�4@aMK`���U��8���Ot��N%mB�7.!�7u�Q*MH\�B�Y���L<�������]�H!!�\���KiT�\�[Uy�h�2e�M��jyWOsU�Q�T��@�Nǒ�\�w/^��%��fE,TG���c��%*�e�1V�5sA��E���ذ�0��lT�=�b6Uƨ��UeYx2koV�[eQ2+�.l̬��'�{t_��n��*�e֘rRЂڧz�6k7�����n�Y�1[:ռ���������W��s^B�2=Z��k%:Np,v҆�H�������`yf��aؐ��8N,N�*q!���4%:�r����O-��,4Q��X�Nd7R��p��,��![M|`�C��lM�0aո�ƥ"�Ux�\�QH)J���D(M#D"�����eRX�f��d�Y�	���f����N2��Z�nK��њ��\�H\@1JQޜ��CX�m��b���  �R �ԭZLr�	y�/l�8���r�^@���>��6��.��/Sr��T`[aQ��5s)ᄪ-�z� ad̹���9���s)Ժm����V��˗$b��S]�ڎ�X����V��&����`�#�H��r9���-���2�Ή$z^!�)�Z���3]ЋO�u+�ڊ[�$�u�YS3B5�kv�bt�c�MKÅ�5���nD�Y�P�8��4����f�Vb�6� ���%�z.��]���f-`�rв��@��Z�12�m`�L�`�b�2��ke�9s,`EA��%Zr��_�H6ꢥ�����6����f§ɱ�U�"�E��ᔬ�I�j:�M����K2�b�Kdv�̵�c9{s^�1�"�.;�4k�*�t5�t�36[V`*�qcif���u(E%�v�3j�ާu"����9�ڗr3w���K��$x��׼q���!ӻxi��Zjf4��T�eS���Aǯ~�/"�ȊȚ��#[$f�°>핽�Uɡ۠M1n���ŉE�4�R�y������ܩ�]?�RqB���FoZ�ќ�.nh�D��4���)Ey���4s
�&#��}�Z����di�)��c���5��픝��ЧH�-+�t���5�(r�ͅ�b��bݡ����X��5��+�oZ���.��� 2�-��L�.���e�wm+,�M;*|�[3��B�^Q�%�ccQ9���xֹ{@��H��N���r��Fv];hm�t��6 ��P��W��)�OὕAXQv�D��a�v�����KbDQ{���P짯�-D+]���D��uk����U�~]�f\T�W�QTr-�>š+ �c&���e{��
��M.���RY��w3`�5iQƀ�i4lF�L�W@���m����]�I[��뇳��E�c�u����\;�ն٧ޣ,���p��r�^Ri���C��6��Cj6�"GY��\ �!yk���(yV�:m��k8�.�;�T��+�9�5ra�ӥ�39ӏ't5���ù\%��;�#�i0����1f��D购�cL׵ɔd��
�+o�I�S�$��p�2�����'?�[��v@�P��xw��1��z��˨Ƙʑ5u}� �e[̦t�3�'�΢�Y˳�����I�J�o���{YG���ynw��3��ҭ�2GvTN�p��}�賵���R.�C�!a�E��p��%��{[���ōg�2�\�a"h}ŏK�ޯ2���m��W�]��ڭ���vv���|��=�m��Gmѱ2�OsC ��Y�I��ضDt�J���|5ׅ2-ژS��@�l��6eL��X��F��=ח�v��Y(Qy�^���M��Q>i�����*��SkC��v�'09�Vi�)�}L�j�]ݢ����InKCqBW}4�V��.�h�V*D78��p�M��ho�U��hH���鉈o)��1�=\ck�2vVS���
yQ���̗tPUb��x�һ�Jx���އ��繼�\���KB ��s+b����#����St��f���>ڜ�I��{ŋ��)"��78��ƿ��J�*т�CY	'p'��&����`G����7f��kZQ?;���SD�cpq�$mU�i7im��n�wW�b���9�uZfm��c]!�(ЀM[B�Q"`�J�n�7xf�x�I�[i���.͒�ҡ�&�N�K�tA�-�?+;�73�7�
���� �1ֹ�r�	�n�Ƈ��n�7U��_O"�.����nyI>+�Ƈα=�J�榎_vY�;�M@����s�_Aj.�[{q�@����bfa���H�+�0�exb�(cw��k��W����;6�^8Y�.Uؒ�E���3d�uy�^��ݍ�W��eJ"��W�,�V���Mom*�l,����r;����#^Cj��'��,��&�kq��I�t[##���U�V��%g'��w�֗&�)��+���7��[뉧V^��x�K���:�n�2���l�����޻2v�ci^Q�ǫ��3�̇�$�q�Eٞ:el��r���:��s��wI���_V�U�x�"�ݮ�9�[�D�"�pZO	����W�痎��ݾ.�U��V�v{v�)15����
[��yc{��˩A���؈P:���7V�N��G�u�ָD��$Nz7��F���&rY�y'<�^o�o]1$0�>�3�-�	(a������`�uX��nE����;y����л�����W(�����vc�W\�^�kL�����8���nDoEf̘{�r*�u���\s�;�5j���^�����*U�Ok�!��,�5u8��@�s���fܲO�8yIc���Z^�R�L!�P<���@(n]�!1�ݑ�֭l�F��Wz<ط�n,�T�z��M���r�v�o/.�F*B�텹J�J��'������oVF���K2=���@��SnvR}���Qg�u�=J���Bi���p�Q�g1��������z}�Z8ޕ�	��:9]�C��l���n�V�������yn�z�Ve�8V�
F���Z̙���N��H�ի+�PZ�j�N�W��.�_P�����d��]��Zz�ৼuT�Fh|�CR6�O�v���@r��D�w|�o�. �˥KHFa�	�J��'f�Vht�	0ΛS	�Y�h�{b^v� ��.��R�v��A�t���&����u�vuZ�4�l.<Ggu	����d�ۋ`�Y�9��jx�-���'��;[�rXN	�>����<�]� ֵo�W_u�	z����E �,�RH[F�by;E���T��V\�U��RY��eψe��3o(�w'<u�1Y��SZ9sl>�3��p��t�]wcyNА�k�捽}}{p��*�2�.�ū��+}]Hq=\)�.��L�'&��]�ebt����۫mCV��Yyk�Y�)��4rW=m2�x;��!�{�g�ͽ�˻��d}o�r��;��MQ!(!�Z��"�#����B��+��ܖvWi�]����gr$ஓV�;�!��n�3}�3-�Jqy}\,��qZ���mm���(-�oō��*B��kX���c��yʦ������ΓY����.U���&e▯t���>!^59��A���ɠV<K�-���˰�I�U�x��!�F;�����&�B?���}Y�ek�++��]q-�7ud�Dnq]�<����3OtU�Z�����[]ϚKm�;��9�]�W�,ܣ�ӏ�I���S8�x**�ę>������b��~�h�3���f��-�����&��:}�n��lj�Q�N������L���m������Q[R��fD�a^����;!���M"r��6�����V�N�$P{��9���k_Q˽��a>�)��h�.�Lw��P[�����K����S�����[�D2�s���K�w�]a|��u�_w�ad���9�_�/}A=|��1���^��F��y�#��[�A��/���Y�V��끊��X�h�4����A+���\6Ҕ����`a4��z�Y���D���;Xc�G��Qu�iJ�>�k@�j�����+Q3�V�{4�U�MCݜ]�g)$/w����+�r�b�w��%3��wx��#�ڋ��^�Ä���Vk;�����L��.�b�w����k݋��_k�.�0�u���� W���9˖L�k9���JW�L.���W#�����:�-�̭�:������%���t�a�>�A�������0��9=x�vf��i�q���k�]��)+-n�+r�t'�IkV����1S�k��4�MIO��gpy7�
�]7jt^,f�����z`��r��:��9�>se����4���6/2!����A������0���j��b��U�0��X�B�L�ޢl%S�wpSz�����ԒY�[�Lnm^ ��m���pY�8��T>�Y����DT��}�oj`�,�H�1�,b-Vn�3�U R��������}�»jZ���<Hy����mp��T�B�-Q���X8K��Ste����	 m@B.�1|���I9bA}�t]�8��fP{yp�9(��/=��lի%����e~��.����rݭ�v���a��2��\;0��T�ݮ�/Hl�2�iv��&��k�ú�����c��ɶ�mZ��﷪n;{�d����f�k7�J������uj2���L��k�s�фM����P��?�G-����upJ��ҍ�΄�zy����S���Qv���6���ʋ}��pI��=rȡ���s����e��M�TT�VV�+{�qA�SA�����aPx���.V��Tָ��n���h�9v��s�'����:���#�mi�ލ��ر4it�䠨�Z2V�y@V�h��r�N[�C�/�r�z���LˮG��pf��[>�EwѴ=�ݕ���FB�qh�y��Nm>�N��o��� T_sѶJ�O�W�V���ZG�ZFi���fG��[)\�g|��f�����K�E��+�<�U-*��v�m���8�f#��f�"�uax�H�
�&�g�ϴ��+ �S�����3��;d�>���Ă�ï����مv�^���$����7&x�y�wtm��w�+�-4���y}�.+k�sZe*�qT�JCHRe����2�����ޣx�����ܮo�u���u�e�6�;�)˹H�����X�(҆kD^�y��T�vԒ�Y�a�#-�-X4���7���	�zdX*����M�C��)N3˖�ǌ�zL��o�v�z�?i��}ջ�`X5�Ze�Tڃٌw��ڗ5��̧Ӕڬ�^�D͋��y�V�zc�HU2Q�ܓA�:8l�'�I[R�W����^������;�/�HXw3%Z��GD^e*O�<;�nxxٶ�Ւ	8<%����,~��=p��]�r�:܇�W5���ݖ�����OAD^�q�[�=�7��U'w(1�=��/s<K�땯1�"v�䜷��4�G2��񊎬b��:W�Ú�8�qt��S�^��u���L�GIJzQ����z��ϧ����2�~mC�o��3\�ﴝ�j�\��6��T���L�=_�/��?wn���Ӎ�m5��8H^]��d�2���y�|f��ՍAlW�(��|��3 ��䇸Zr�7��812��-��qk����50�|T��zĻ{#'ܻU��z�| �]u�X��;�ՠ�b�&����gL�a)/v��1�%Ӿ�7�̔VlX�^W\Q���Xeӭ� �)���J̔m�������b����)[���9aW���_xݺf ���n�tl�#as�����kj�:��S\�^b�����wvܚ�;<H����Q8��	}��ùԣ�T�$Ft�����WLjJ(�=�*>yP��,�*��_r񻝺�f�y���s�'����s����j\�f�ji�^�feu]4t��<� ų�|�˨CM��C��Z}�n�*jz��ǧ	Bf�L���6r�,���dK���_7��_XmKM\�o[�g��k��!�X�Z��'�Wb��[n\y� c}W
�oT:���m�4zc�i4��t0N]�KwFl�a���]WW���R�oZb<AZӑ.��E#j��(FB�{n����DCFS��(��ů��J!�[�GH>����]on�ǟ� ^==��D羽Ao��b�z=O�avؼ�c6��RG����ɽS�a��n>�k��7&�Ùq��z*����
 c5�e� ���̕U�(���*L���mi-e������J��7l�W7�6���oww,ݕn�=�Wлn��.ٓg*լ-������앯�o����r�ݵ���[2,7�.� �֯#��p]W��H�,���7�t��3z�5�0�p8���mˁoa�M��˺"P��jw{"�Y(��$̗�a4���PH��15�v����$IV:k��Wy�v/�����=�쾻}n����m�c���˽��BԬ��Z���sWWc�6.X���v������:���z,��e���On���
8�
��BHܱ�T+{��7rK�J���6b/p�v ]+7@n#�Qwψ����^Χ{,}�Nm�}�*�O[I�b�Y:��M��9�B�%(r@�	0}�8�һ�:�K%�mS*6�JCim��u3�QI�;��ӎ���a�W�wQ�N`�y�E~/�.�s�R��P��3�`�T�]�6��o�U��l!>�W|�Vtp���32b���m�<��ݬ�ӳ��.ݻ:�^�U�=F*�y��j�5��m��	�.%"32}}Ef�+ո��:p���X�(����<�٠���Xk�Iñ`�͖��I1�Zm4y.礮�I�rz��h|���c�eӱ��˦�sT�/Z�K�>�T��N�߼��,%	|+���i�=H�v������Ă@B���;��U�֧ֈ8�^4���(�OVw,�\�qT^X-Գ�X��3�V4EA����{���Ǧ@V�����t֥SSk��+�;i�׃@�j��
Z&�9Ac��6�=:,I�RE'�~ɲ�A��1^�M	C07Zz��՗|o�B3.$r�)az�Ҁ�+��j����y]��h-]�J��S�ދv�w������
�o��ج��y9s�l=���yiGOh�$��I�K�>�'��m\��3Z���C�I�k���7��pꆴb�zsf�p��9��xٹ�`�U�ވ��W�8��Is�u-�<){X�z#�0��	�m��:�մ:@����WZ�̊A�y|_U�!�S�7��S��M(���S�bܚ%x�+S�J���V��>�S4*��C��B�����pഅ��*�݁9u�׋�ͤ�0fe��4����y�`D�Z�Ki��pgF�թgweU�iRm2���LE�����p"�c��8�0_r��3��t�if�6a�f�?v
A��ڎj���7�4Hk�E:��w�!8u��` ���k���Y��.�{B�Y��*��<.�>�g��8�=�뱡��ͣ���Nnn)��[R��4��]�3'�)K+�W�����f+Wh��� Gu������k�����8��U�-۳�+�����pZ��s�Nu�j�3%�nP���+v�1��'P��Pze������:�I�!�'0��n�e����|���R�}�l��\�uΗ̣"��W�� ��:�YxSW;/ow�{��\�)�wa5�#��h�Mk�C+L�	�#���i]�y��Ϙ�����=��bُ���)R��6�+J��cH�i�_�]J"X�O���M��I J�H��dl�:��OV=5�Q1[�a�휮�g#�.[�pỾ�S�Kj�+4Y"�ڥp��#~{BU�ƆVZ���@�H6�kn�6��~��g���F%�|.����R���������-�?NN���k����~�+[�I2Mu7^{��^���R�K�{�cv�]1��f,H����\+ ��Aw�z�N��ڄ뮄j�GOMΩ�i�.]]�� íCs���I����r5.�[}�yۜ�j����6�����微��ҁ�W>��ҥ#�8�9����=���7|�b}r�{�k�l.����r+SGr|Nl:�&	.����ZH:���M�n�S'n�ޭu��_���PTA^�{�����xs����k����8C���B4��j�m
ܡ���[��u�B�zoA�Ⱥǯ�1���a��H,��:w���B�0ge0��]لè;w]�����\����h�6���EnR��
�!Zx�*�2.ߎYv���\QkzߴR�.��-+Z���:����ں�M
p���upG��On����x��`=�c�ڻ�d�����}��Zg1tĨ��7l#����&�mi�?_Z[��3҇ē�sW.�>����~����n��������/({���$�B���L]�ao�)��#��3�N�!��ʏ�M�XOxn�<]#Mr�4�P�)�+*�[%XO79b���)ǝԫ�&���/j�V_�fb���0�j���Ȧ�tD�n�dљmRyj��w�s�H�8�L�o�e��᜗]�1Vj�Y1�}��XYْM�-1��)�Cz�v��jgUf$��=�����vu�O4K;:�7�w�x�|0�N��%V��!QK����y�msSp�ZIU���X{w���c��Mh���j��©Ԓ^�jU���e��]i*��+$��wc0�Nn�jg`�Z�bfV�".|�f�v:(�H�m���kd%k=���&f����\#��~����CM�Fޗ�D���A��Ϟ�yAYn�9�/1|R�&tƲ-�n|7S���r�N�5����:U�D�\��Q��3�|/"��Rz���Q��ej\�̻T'ϋ��xL�q%Ӹ[�K�vk��0n��#��8`��=\0Ϡ5�/�����<�\�2�ͧCV\x^�qE���M�khک����ǡ��T�w��;X
���a�r�Z�VZs\�h�s�9�i��u�O�7�;Tn�����cH�N���s�2�:�s���*�#��g�fw]$�7�$����p.]��J�/�lH�,�e��1s��)#���d�[D�]���}�!�Eg8�;U3� 4"I9�.v�jr�n�	ϖ�;���f�d}|6u�����!,7�d�g'v�T�(�-��n�h���`ݖGEU�wT�(ܗ�i��t\f��h3s���a#5�ױv�v�|���4�7�A��X3�Q����BJZe��)&-w���6e%֩F+%�\���dE3��3��:"�`'r�ڷ��F�Z{^p�;j�TNf�i���H�H�B� m�5g�YC�y��a�C�������ab=�q��z3�9?q���0|���ng��$�ټ�Ь�+~��qd�/�������	��D�ݝ�r��#r��L�#J�s9r�������q����!��d�5I;�N�Ǚ�o+/fw<Ls�s{�ŝ� �60�����Z;AS��
d���֨�fA��p#����n��\�v��X|3K|U��������jS�,�N��i�"�9s��!��=�*��ِ��r���/YM}*�E]$��cV����Aщ���+�oΒ�<3��<�K�η�h<����s�����g (��k�Z~���$&L�1h�%�5���M��˾C����F`�\a�Q'r���D�x�6S���Ԭ��:����G�Ì�ׯ�����5z�a���w7/n�cI���kk��1�c��/˱������_KYn����ͣkJ$`2�	��v�Z��7B(��B����`�k�b�!l����KՄ]r��U�m��jec��ތ�5�2��\�7��m�;�Β���-U	���3*`��x�98s=-�4����>MkH�7�tkO�+;9�����up�'�Z��a*�hA:!�8�V�nZ��9�yFvWa�Gia��sh���+��'�94���?gj����30k�S'@�Xk�v��Wz�IfYu��q=wy�kj����٠�A��}�:��t��Z�j>W��s����=��h�2�z�V���
�t���bP���x�'��g`]՗��:�g5t'���i�X�͊���V,�O_Q���K��
�gJpЅ�u�(�ƪ�=�n��cg+��K���ϟ�q[&
�"����rs#B{`l��#��4�1��Ȟ	�r�;���PHe�i+�fJ�m�lǆ��@��ɂ�M�R�pb�����68�k,8��A�9M���+X@��Q�k)�\��J8r����C��ى�N��hb3W�� Ȯ�N�ee,v���r�yX(�)���
� ��/���nA�M�h�P}C_E�K�j��[RR�]x̘�ԣ��u{�&�Kk3���{�*n�GL���a��3yŦ�Nen`�{jP�z����uD���{�k���Hc%�8�����O]�:�m.�i���=1v����r^���*áΞ�kY���[�n�vtLJ���)��v�q�ʾ�!K�rZ\�^,S@��WDwK�j�Y����/_`�;�<Ã���ͺvH�	�'��%�|Z��ȑ�hN�1�;�T(P-$�����*��f�^u>d$_(;ǥs�UfFw�����H�ntF����ݝ�3�����C%��z���G9Kw��v9}XK f��u����e��אK�T`Oʰ���@k��ػ)沱�X�峾�ċ�EMj��R>�`���%/��73���/B�v��kn*��X4+65��]T6�b�^��7#䫫0t�Ď���op�m+[�F�}����k\�_PN���2�5��Wjy��%⸅ܰ�6��xG���
bh�;�K|���F��v�ǧz+�h-L<��DS+��ʺ���W�ąlms��0�z���U�%)�`u�F�x��V�X�Lcs�?e��P@�Zu^Eq.����r�^Ώ8`�ܙ܀N]���iOlH�}s�0?��5�[<y5ǖ�^����+�ll��һ����.�r�}�p�5���E�2ys|��4��Z$ԡ>��a�,.�6�5]0]�-�m��#���JĮz�@m[�oF彥��jK��ߖH��]�y����b�+o��4�Q�H[����y{ �yP�:����xsݎq=�1���2l}d���7Br�ͧJZ�5��M�y�zQ�A�Wfn�j�4A]�^�m�D�b�.4��`	֮v�ݸ�ud\a�v[O�{�0�j�o��=�q�!����8{"ް�p���<:�Ƭ�(����l��bw�c�nP��F�����}W���F�ٜ�ԍ.�|��|�jIyȼ��aGF1�_WZ�c	����LW�:"��KG�F�L��=��9�V�80-ާo����Yո�L�}2�q���,�C���;#�>�#_a�19sG�#qY��x6���'7�Le`mQu����[�(ʊ*�Z���A.�Q�c�uΜ�g_��r��Qv�^8���4�(j�~6��9v�ȇ�7V��yܥx14�X�r�71�N��vY��>�2��E"�v�,��(�(ϻ��u�s��OmAz��7������G������1���L��ԫ 1�������5%��W��Y[(N�}��b&����\����J��+L�υ�W��]�Xk*Ȳ&l���S�+wEv������ڛ���,Y��;.*�{\��;jn)T�,�ա�����tL�|���圧k]��v���g'�恮��������KNث6�;Gb�NuɌ����T:�g�ή;�P���~r��<�����TZ�������o:�6L��(�wV�����WYWe�u}���n�M3N�)ܲ]c��S%�� ֻW��c7�ڮnJ�A!Զ�R.�����r�ns%mm�ٙ�),��v�}����`�ʧ_.�V�+����f}}���^�WQ�2�1ܥ�84�3++��G�j��V�����a7���E�^�ym8�髗��`Xxu��U���3^��R}�13���}j���K���NϷ�%���sg!Ԯ�ѡ��w2$z�YU�F��8�F�u�|F���w�$q:z�7ZAM٨2�LY@�e�����[ �%�n�/k(��+47yK�B�c#��X��-~���h4�;9u��s��ZY�'�������v�d�)�`�]�8���ۢ�+�+\8�4���{�h���n'z^�w'�J��[�tY,��ڝ����f�>`n�z�S�Kٍ�q}�l�g���:�o0f��5wZ�$�P��������y�8wnk�n��C+Aݲq�s��2�	�czA��³�u�}wP����V+49=���s�B"�ܻ������E��݊�rt����0��q����F����Ǽ.��_o^� �����8�@ܰ�u��˩�Y	
ޝ�1�q�3�]$g����s���=��ͺwĉ9f�XsA�>yO�<i�K;SY]���D%��C�8M]���\Y8��TcLT�k�+K��铒�O��X���x�܃޳z@��2���3wae \}[��R��[.m֭��h6_>�M-�z1|e�a<(�l�}����[�Ԁ���a��f���wJ�1| �L���sܧ�"s�B��ω#n��z-��2�kU9��ի�m�fX	+��_}Z۝������׎�N���l��<�<�,��*�{7pYt��R�/A�(�h��:.�Jn*r��8h�l\T��3��)��)Rf�^�L�|;^���8X���lx�"��m��hd�kN�N�:Z(�%�|L͐_f��Ǥ�CL�tm����H��&�%K��gD�Ԡj^Ǿ��7Ү�_j�Ƹ�e��N>�0���''���p@6����5��-�K��q�{y�K:vK���@���b'��x��3�iǟ[�ӫ�Y�Vm���Ӣ�k\��V+��V�+c���	��`��-�e����W���p���B��i��w�A2��� ��"�+F0�LsW|���}�4�m�R�(sL�ǚ�j W�D�gڻ&6̭�F�r��j���3���ܬ���0J*c�>�Ly+)J�xp�jL��%@�ڶ���C[���ej��1���!�qX�v��rr�.�J�O`b��C�/�n�)nʘH�����ݶ^@\lQ��lN�[��gv���O;�۳
�0C,ЫgU��aM������-�V÷"!��V���<j�u�Ns�r��_{���x��q�P�<�ӽ�D�%֜�	T珋�3ug�mts44#xE乯����<�]`��V�]`����l�Y��q7���ɗ�0���-S�f&1C�}�wZ�����W�����9��ի���JQ�Nax7w���43S�;��؏	C��j��p��ݨEr��z/'6��Νf'�p�+)SR�ؗ��I��7r��7a�n��Ҥ��+}����Q�e��B������/%���G�.$C����=�&r�|���^��Q�gƥZ��1.On.�Ε²�K�Ձ�M�4b�eT�iX�"V�yu���t���nm2;�v���[:gX|���͡��E
������ҮM����Z:��xWr	�5SiZ����Ot�2��{\�5��}��-�ieЫw�fD��VVG�u>�7�i�b2�Z{��R�D�]/��rr��%ud��e|T�Ʊ�J�� 
�5�rs1=ή�Ef�ґ��g����ګsU:΂�Z<��ws�̯3�x�}������k�R8�_;Ӯ0uhA�Ǫ�^7%�LeF��IȪ=t~܍���6�<3F��*R֮�v[zܜG'W��@�L��=��5{�f�n\�)ƈ=�!^�TՋ�n�}��5��ma���m1��3�Pc1u�OpR�k9�ib��1<r���yZ�[B����\�B���x�u���f���و�{�n���m��С�B�u\H�J<���ޣ9`T��^�\H틕篯��ry�����l��bKN������m��G.@[�f��r�f���P�t�왁�Z�����h�V�q�2���/����,��T���ncd�%i���U��Kv���ͷOR�M��wa��ٗցZf��l<coC��f����kBgq�V2a�W
����0�9�7m'�ڕ\4�.�v�K�nS��i=��>"��
�D����*J��NJ�-��Ѕ6��6�	/`��n��x?{^�#�yv�e�lM�]��Lt�]jk�U g[�4n,]yyx���|��NYV��G���4���AN�NM�<C�=73���p���}�D%
���m�b���g(t+&'v�.�V�Z�RI��@��+b5�(;��:q#7��՞T�wj@���>��8U�}X�8���鳰Z�N�{{~��5Al�ع�m����0	�Q��09`��J�W'���q[ iʍC�Fa������='Z�C���l*m��6��(��K��qT{�z�MY���	u�]��8)�Wl��P�y[�B^�Ķ����2�4�$��z��Z��r>�Gm;��I��J�KåR��W�|�&$V�vz_
��(���ד6�dL`�Ci�ؚͮ{H�]b�e`�3u���M(�7K��y���J݃�I��쪃�Ob����rTS����;2't��o��>i��~�]O���L�}Ȥ7���Ր��N'i�]co�K�����fa���F(Ͷ��#kF���;��0劋�t�{w�7�gmfG&;?H�a.�����2��N��<kM�3�]x�um��p<�K�յ���T�]����YpFF%��Ŵ��\ﮚ�R�Iv�GzE�`�Ă�t8ECh�t�ZWSWjo��C��o����e`���+C�����Gh���ea��C;C�F�v�|G�{����|�}_|����twލ��έ�$�\J8��'�5�ƚ��+4+�r�.c��V�a耑q���$G��;D.�m
�&�m[c�W7MG��l��m�#�K6��rQ�n�ˮx�B;�Sˡ�B�%~�;ۜs�[����f�R�fC��8kg��{�+ E�����@ᇐ�v��fJVwE�W��UI��GlI:�M��*�V��3;��[3wN=Y�|o�OT�n<��F���gS��3�Q2QN��C3��kk9ڝW�ue[��9KT	��i�a��Sn�N��V�V��l�7~R��K�I��x�U����,]L�kCx�j�U�,u%���u��犜O;����-yڳ�h�]�Ul�����tιw�u�u�{[3T�7�U�]\�O ���5ܠȲ��b��[mY�W�,}:�r���ו��i��i��v��}��M=v��8G�)�=�7�t`���i��|��X<,��dMZ.�J1����m�ީ*�x�ݜq*1����qva%  �srl�a���7��Z�6�3�$?����F��׍nn��<�U����Q#k)��-���J6�{˖KG���rm������i��-����U����j��s:S�%�|�eXx��z�����.!0�^ٝ����*�Іk��H231�Y��A[���c�g�u��]w�ޱU%4�_fTS��I��FXTS���3��f3D���QUjr�"cQ��%V�V��(j�")��
��S�SDT��")(�¨��"��&0�21��&�K'"�4ԔTT�����b*�u�5Y�P�5&fVY4QREURCMD5Y9� �JH��d���cU�T�AET�DDMD%&kY��*&�Lb��,"� ���Ud9eE`AVNQ4E��MXf��DP�TPPU1�Q���rɳ,�¤��Ȳ
�����*��5�V����2��2F3(�������,̊��Q�U8�Fa��eQ2YSE��IHE���aU�9Y�PE����d���J#32"��hr&�u�j+ ª()VE-�5*(�}�������{��V+ES����
"\����j���V��ú��հ��mH.�{]N�t�f�A|f\�@Ce�|�W�6ѻ��<�>>�'-�a�c,X2��46��-�*q$xp��),`o�_N���h�4����=�l���-h8ʄJO<���f�'üqj���v�v΅�Ӝ��}��e.�ЇϨ���h����T�2ڌA��W��t^���]�Xϩ^foBM���+��r��v�<���\E�;���$Ta��߄���u��/]S�3����(��,!a��!�V!ֈ�v�&hfd�E���C �5,మ����?B���ӗ������ŧV7���| �9֨/Я�l��y'��E��U��ǌ���d���n},;�ʲ�s`���� U���מ�Mc�]j�U���Q޾�h�>'���5m��w��DɌ8B�x�ړ0R]s���lc�t�A��|ˬ��U��	�'-f�צȤ�^�_��Vx�R$���br���=C>��>�*WB��ޣ�v��>֩�Or攱�k����KmuV(@Bm�p�4�Y�ifZ��>�ά_�Ayh�!���䚬z"|�+��Zí��d����;��l�MV^�`T�r��v��u�*���� ц�bYɜ����|p��
��C]�V���$�k^�{j��{�����rq��s�T�G�:5WHn�0uJh�n�ksB8������|��{���.�{�K�ˍq��Vڈ��xS:���X�Y=�A�:;�*)���Ԝ�y'ҽ�܃��zL�x�5��[I��*��˪#�W[en)��P�������xLr3J�)�{1�����E�f��wkU���b���@�7�|�~���k�>N>k4 u�ٵ�!ƾy��9�w���b"D�.�5����L�h+}t�]+F���=>�җ���4�^�\�,Ƭ�.���o`�Aк�l�s�{�l�U���}Wy�{4�C�޸�3e&��C���=��M,*dmd�=Z��[x=3�Ҟ��[��BD ��9g����2����ܮE픚̎`Fĕ�S��"�.8��+)�H΀��*Qbd���!dW
�g���5ડv`����+w�$�oo���6W-��w$&� ���s�&�`Z:e�C��K�gQ#͜�2I{P��!��cm��1Pt�2Zg�KIX��bK���-^˸+(�v�ƱW9{5{����sMn��F���y9$�H��\/U�s��f�	y��%4�;=��Cv�4�#�<�㢠�v�qU��0Nʑ^&�ܝ������"&�x��y�/���`����{`����dJ9}ANU�-���b�-c��/���Uw�Yo��"TS"0{�o�=�@8� �����u�u�ʛU�n��)k�.3R����^zwM��Ǵ�i�q���o�h�n�Fz.��t�X�^�G\x��X�8�n'��y��	u���1�-�'�ΰ��-���+MlP`��bu-a��z�Ϲ���\�Xrvk�+lU��<%z±z
ʤ��AU��!���5;��6�o������Z���G��F�Ī�2x�xA澎�U����"�O�,����G����(o�zzl!f܂�s���OJQ_�NBarޮނƵ��Aت��L�m��6�qF�]۴.��U���;�O�0l'�M�c���J�=59`�hu�Di'�`�z�24JW8��I��z���C2�ڇ{&O��d�xE�ڳ�t-�چC]g̑s��,��Vw�6�7��B�B�0i)���(t�2��9�sT^�|�Ү��n�{&Drv�5��W�����7���ba�k�t�4G��B������|�yG.`��W��Pd�p��p��ogf>��U�C㸯gu+�n��l]��zɗ�-�b��O��z<�EZ�E����+W[�� �'[��uq㾅��AW�e�c7�	�tջe��{�t���w��d4`�!4��j]�H��hv��]�8�VJ�y�`��j�_r
����K��-�F�WT�H�JM+�du+3�3b��h�h��	�"Z��	�N)�xevo��}�,i�$�kD�&�Cbe$��R/�>���^}w��Վ^e����~,^O�S���yy�����V\P�j�;%"4��a�z�L�<��r{�\NP~탦�03�Su�W�)v�=�,M-� ��s w���`���r�ɨ�F%1P���h#Ez�!�i3T��V���L�#�=n�}���v�������s�+:�.X���/,iϟ��vu{V%M��X�������ł(����xJ�{�;B^�߷�7	�{q��ϩpѣ��"|a>G	����per{���[��3����3��[���c]��S�9�V�|8��� l�y�)E�%	kE:ү�w���M��n��-�O7h��g�-�I�[L����5.j���Qzm5��r�1W�*��tF��@�v��B��	��o�����H�xԉM�Asl9�U&��kڱ�30
�,��<�GC��3�(H�]��71� ɝ��>x��w�p$����"	��N�盃�o�Rs�-�4íٽ\5�ޭ&�2�"w=�0�cNx��G]ٻ��5MN���rN��ڦ�:�w �I4�R�����^��IS����*���5��|�;�-�xv6o�H�xN�������#��wv���2��~[%��G�Ӣ�:�<��J����~~sg	1y絁7��jQ�8瓱�u7�d�a�u�4o(�s�O����^}����C��х�T�����v�r�I��g[����\��*��~�̔�Y�܉�=�{��d7���Z�1�̗s�d!��=:��ޥ�E�,���@�5Iί���}������I^
L��tK�tj��k-���g��}!F�X�]M���O��2ę}1r�k��f$��e��VW���|��Ω�����ν��wt��O9�%��c��X��Bx{/�A!����{������׻�ҷ}�A���8���8���]���N��;~;�aZ���=S(�Y[�u��p��o�,�������� �)w�&A:.{Ȯ>���%����
�GM}���w�*Ƙ�f��ge�K�F���S��v�R��BIM�T������FQ3�[�ʻ{�� ���X]�����͞}���J�'�Z �,���=�ukN�:���~9���=y�g����7�������������@���α�~t��u�>�l����dq���[��qao�^v���M���~�1<=�ֶ��Oi�����;��Z�'/0>�f�ި��4�WX�9Y(���h�>zkֽ[i�l/�̂��͇�XNtσRx���;�x���n�Y�z��s깶���s�/S��˦:�>bC4L��Qj�m�0�5�J.���P�����-��;@(�v�u+�.l�2�xU�Y���AjNci�͆T��rs����ĳ�����x!̛��o�a�}Z���v��w��OxN�y���[�)�\�(J!o�ԲG�a��͵$�8�=B�f����k�.'��1d��r<�쮧S;fRph7�ʼ��DT�4�h=���-������ݟ5/pI/��B�A-�F�W]zVv�����^	�{/���f�<��mB���qn�H�%�T��7����Ɇ
1v�}��SiQ���l�.���q���Iw�i+�L�N���w��*e>W����y6$磶N�"�6;']��$�̈́�lܛI��ǜM�S�S�l�>ieA�6Q7��ƾNu_�n��.3�	&N�Λ��Mv�b�����W�:�m͹u��k=��V)��o���-��ĕ^!�<�vO:}z��fN�m���Ϩ;�`vw�e'yt���݂z?r%v�h���җl�ۙ�	����$ǧA���R�a�~�R�]p�/m�1M���>x�5{{�ꃾ}�\���ǧ �wkge��W��{����dӹ��v��2�}ٷ%oT�%����f��ɻ� �*^uX���!�׻�w*��e$/���`�N�������0V�`'/qlY��Jʣ���������jd�ʚ6����_B�ί`�I��=����%�b_��^w4z��m�}ɿ`��귆���i�^�a-�)�?Z�ݧ�˼m��ry��L��lOQ΁Ǜ���z�2x.��N�����i�c
J��lYcO���8�+ɉ�v
��<ZބMiW_���x���|⻰�O^	�r��nԬ�e�CN�Ӌ�Zf�s��э|YwE����r�r��6�9�p+ٙ�ׯС	�[�;�b����������f�{���G��Z��������@�#�~����?s�M����e��	]�鸢�U6���Ja��H��ϭ��s��ל����]��[���;��_`]����L'c������W��ut�8�:�rs��O�f������p�z�vm����x�As�� �}����϶xJ�~z��ꯩ���%J*�������ϦK�0:vJ�Y�K�U�{Y�;�^��T����I�?O�s��%\p���bI���)�+�g��{)ϫ\���v='T���Wg����	��y1r����^ygj�6:'��-����h�|8�4�yT��Ԟ����4�b�/M��zz��yV[>�-��){��RB6�����뚲�:��Sy͹��p��O>�kX;M�lH-�	��b�OF�|�fQ홹٪�:�f���f1^/f�+5�K�%�u��>7Е��w^SF��p�6K��눐���ɻ� b���\X��}9Z��m��-��M�x��p�ѭ�x���݌�ަ�)�񦓮���	M�iz<To�96S��_t�Mav�N�Kk���o�7�;o�t�]����O���P�m%o���v�+��B�
���>�;��{؟����q��w�_o6�r��^u�b���Ȏ��[�xw�u�f�a�3��b��zgk3�ԝ��T��m��u��8vo{�O���ϓ�W�}�z�[�.�G���E�<5e<}��x�ûu:�.������=kk�-�*��ٿ1'�M2�ɳ[ܗ���73.�#o5��ȋ�Ư!�X�_�2w�/-z���r�5�~��̡�X΍Y�kڧ�G7���p��,�:#x���5�}N����yq���U��ލ��;�0����{�^�e`:��Ӣ�>�:CHc��h<O8�:�=�j���5�u�wI{RVԙ.���;!��O���ŋ�&���}g����m)o�=����{�Kѕ'�X���~�u�M��`�%X��G�:>�M#S�^�wq��24K{���R�xhfee5��F*uhT��j�IfD��ڕ��dfհ��f�W�\k��u;a=ĝ�.r�ʶzMn�n�Ծ���V��k#''�h�5��U$RV�Z����x� ���B���WOsoc�����L�>�����S޹����+��vjrQە�o�t��{��u��o*��ݦ��#!���=b?r�j�q�~��-��wN�;�D�׻O:�7f����[���pkkFJ/'��sg�l�hg6.Lzc9���}�=S>3V���� �Ēˏq�ǯ�z��6���,k����fzߎ������j��0N~6� �^�;�ɍ�T���@��{��+���ܖ#��q��7ҷ����Z&yC��J;�T=%vF<{Ҵ�ꋼh��1w�Õ�_�9y��{5��N=YȾ�.��؍��nי�]�8�Nj�[fA}�ٷ�:3;�eAk]b����)Tǻ�z�#oە|�+:<c8���X�:�6�����g���<��D��M��js~�=�-���N�}R�|5��
\���]��0%�C����!-���%ZΫ�؂�J謓�v%^�����a����sr[ʮ���T�l�K�t��ؙ��֝N�c��^��;Q
}�jV^ub��ҠE.�#�r]���l�c���vW6�w�Q�y��p��4��L�'$5ءO+���@�+ժI�u��w����]�@�;]�4��dbf���	`�����->�|&����P�a+3�u2��d
�3�\���J���1^m�����A×��{��n�4?)}�yO�<$�❣s.�e-���B��
��_s)��҆����d}Ǻ{c�A�Wu��`]�;s<��x(2]�����k��.=�Gc��n��gZ��wNs��#V�/QtK
�[���Xd�[j[o"�#<򐋸gf���8pT���q���B:k�ݮ׫;Xݤ�i>U���#2QP�������e�����ٞ(j��y�f��vm�z�7i��bnt�oY1s,\�r�o]�Y:��J-�i{��橴�X�2R��������e;4����5�,f]��lm?.�f�z[zd!E=i=%R�7s�&�yr4�Eb�K:
���c�=w�̻-���q���`MQ���>/+\g��_JW����Ƕ����'7�{.�j��s*@uh���{�F���{��k��0�����atV���8�k�R�e;�^d۽��K}�As8*���܁�{����.'Vq��9q���<Y�B�:�K#��kG��U�H��/b�t?Pǵ;�d9̠DkW�_a��k4>�����>�{F��u�K�c/k���͞�ON���$E���Hd���o]I�A��)��C�+�D�V�:O��Œ�s��&���2�3K�oBn-�����<���:��4��1��1ݝ�V��d͙Q��+(\+���i��lc�S]_PS#S��ѐ�F����+�e�ke��7X��
�ݓ�3eܝ�_f��kj���ۺ�W���%��)ֺ�	Om�d\�[6ld����կ��D�l�+
0�����['C�v�97\�9�FїXtN7*�M}�V�.,�Z���Y�n{�d�a��zf���թ�pO�^�*@)��k��v�V�̕ϛ�MՓx���M�+˝��Ǝ��a�>��������o2oP��E+g���ָnP���p�Rۗ�;b�q�[u2�bæժ�gE��q�Y£Z�l!�f�{w�X��c�}܏݊5��(aA�pMd9�����y5z�x�n���ꧠ�x:�ݗ�WoS��{2��"�l�O%[�X���ɫ�����Y��P�rhOk��ӒƤaO�^Y�3n���z��ͳ�{�-������O�E�Ë���|Yf	�ŷ�m�m}w���S�U	b����A}��f9Z����ٴM�U[ dV�V'[�+��۴��J�S���x�
�$pMI�R[|(,���$.�Q�B�-O�K�D�?f�.�(�'Y�јk4h�ՓF�
�CY�B��fd�IAe��XQDS,L�#9�P�e�1E4P֧*�d�̩���f!TUf.��fd9aERLDQ$M-%e��dU��E�
ԙSCQREE5���Afa4UU%M��Fa�UALJY��M�YS`�Fd�N�������h��!�����Ya!�`TTQE4e�KEAT9U����d��5M9���a�����&��L�ir\��59��ɣ#"�Ԧ��e!��Э5A��!��d��b4L�I�f�R��ɠ�h(
ZZ��
 ��#� $�'�I '4��W�siӲw���?o�Ӱxv���Cn��<±Ӓ�Hj����b��՗ÅB��ݸwW+=.dӄ͒��Z�sa�l�	�T��rs����Q�Gh,P:敽}�(OS�ݠWޡ���Ю�um���m���A��^[�+w,�J#�$��{7�Ҳ(�u;U�wh���vt�kٹ�T�n<�\�՗:��������~[�9�>vB��<��������z`�k����zu)�zi$ͤy�׶1��^A,J�(k<i9�S���;~\es�ؓ1.���vv>w��
��l։'�K�<'Y�/e&���c���E�i�x��|9���Bk�+�Kbą��|ӱ�q����t�<�r�+]��N���[3f�j?g7 y�[�l�����Ju�b��`�ƯU�#���b��/��w�w;sm�ޝ�u�8g�oxNK�(���k�v�X�S�D^��{!�����V�~��O5����r��߇t�:	s.��JR�E��뻍ԛ�.8|����(=?}����s;)Tp
Yr�'�K��i�յ9=�[�Ci���&ɘ���~��7�쮐c6mW��v=�˙��^N 0ޜ�ܵ�(X]��{;7g!��Oma]W�[7��eɏ���CSm�����o�bB��gǐ��u��}MzJ)����ve��j������g'�W\�l���m����wT�zS��=��	09��ɑ��#���o!cҷ�F�:'<ϲ�'��CӽQ�60[/��F_���L.?w�u�n����!%*��_y7��q>w)z{�=�ƹ?|�C8G��ɵq�f�u�go�q{�lZ[m:˥&�D� ���ܾ%�e�w9o×D�0{�nt{}�hP��rY86c�rZꃰ��B�X꿃醟c<�ۋ~�5]q���"�U��س�cT��71��k��_:�B�D,.}��8�~}�e��Z��nĄ��]�z��cN�$�Փ%ؘf�뗕Bzf�4-,˲)u6�l��)\&j��v.��]����W}=�!�Ol�+�d���]�>�,Kc��w�W�����Hb�v�Tnm{LS�g]`iŘh`�+�/�U�1s΄1jVڴ�c�f���j����]-q�5vH�jj��UwSMj����e�u6
=كv�h
�vu6�}��K���˹٤v�4��;��X�,���|NuJj��Ϡt�݄�#詋���t���/9�=(]x/v옉�]Ol�j߯����_6� uK�������4b�ֳ���^�}�Y�����]��e\�K����r�:�ɏݾ���3�m���n1����o��8>X����U
��q��w�J�r�foQ���oL�����{��[�}<�o���k�s}=�T��!��X9Y:+S֪dX���s���ޝ��]�*wA��-9y��lOw�[ͳ��U%y���������f���.�q},����,w�Õ�X]3���jN���{N���:����ު'}=�f�лyE�u����M᜺a���mOP�>׺eZ�_�WL�V];,.�a-�Pu����=�i�&˟Q����G���߳|���}н�,�GG��isQw��l�~s_{3W{9��b�Z�S��I��;2�A�W�q��Lcx-�'����	����]����
�q�O5����1'g�r�P9�=�\�U`���ϕz	̥��T������Y�x7�I��#F�ӱ��Үﳰ�o*X����8��8��KދU�w8b�T�����o^��p��,�:#x��\�9��?w��:]�W���@�����j��s��ͫ�edλ��m{�\�1�9][uy8��=t+����.ggί;���r_V	��L�v~GO�weS�a�r�j	���,�ʹ�.��*���w��D��`�<78<}�P�w�r����ɶJΚSe_���sc|?�x���������ًA��10z�h�֐�j�����_�	�?�������?=߯O؜�r����w{r�O��O%���J�d����o�￻���{������{���>��;���!Ϸ��7/��tsz!�_����Wr}�.]J���KK��ư7+��t}�Ի?|/=@x�#��#�hN������ܓ�p�{�8��r�����&A�y��R��ގK�)�sA�;���;��&C俏:���r�W~i�%�*U#�~��0|�L*y����]��>���=��=���_d�>{ސ�:�pWf�о��:�z9#�oG%�d\�Op�g ��4���/O���^@u�zO-K컎�y���{��ٚ�<�y�8k�>���G��|���G�����u�?�����.�����9/ ����^��szyJ�>oK����n����[�����j߾�|֏�_趴��Vs*vЦ���=48)���j�� qQ�i���G��<1R��*�b�Ѻ�,�ܙV�S{�jã�)יh��B(�w�QZ�.��Ҕ�f͹o��Wz�}]�e�h�8���6�W���3QVJ�b;�Y�9���]�p��C�_��X����FO%|��:��<����5.����/�n^FOg�t��kzyJ�}��~?}����?_'���w^,�o1���l�_���������]ir^�?`�d?�����?K��X�G�2?u��)]�ZK�)z��C�}Ȍ�@}���+�}��[p������<�w�b��Úѹ~����z>���^��i~��Ӯ��'��NK�7Jw�q�kJ�#�����>���B?�D�[N�I�_�o9ǿ�;�����4�K�?o�9}�;޴�O�˹}��y/�:��G��]ira?f���hf!��qְ���!+�W�Dp��ۿ��t�{����_n��r_�$:|惸K�p<y���y'��z>��r�9�}n��ϭ#��^~��_cz��|���� #�ЀO�ߧ��Ү�%�:�~7����7��9��<��X�G�^Y���ܧ�փ�w/<����C�]���KԽK�x/�����~���D~C�����F!sm>��W��x�" xc�.���!��N��y���1]���}//%=޴H�{�ǒ�#��/��Od?os�_d�ҿs]۾���?2_^�"_��2,����AJ��u��(��r^FK���;���ш�_c��9d.����ܙ}/$���rW�pv�����G��~����8w�s�3d��4����L����<���<���h)]��}ir2G^�2_�%�kp���jGr�w��P�]��y�)���"�k���P���	~�%�]����G��1�����O�~�y�������&A�_`���9����y[�K���}�ɒ�wѬ]����A�����e�G� (�~��a���̭������O)#���3�_+�bM�;�-�+w��d��]1��mH�^�S[-��m�������)K���պ$�G=�����,,�}�b� �7k�l�'��:��3@�a`���+�+��vN9�zYǮt��.��o���'�{�+��~��rNH�9�C�(Ns �_ �o7�2!���O�]��X��+���}��b��7�����,�Oʱ�������}�?�㏸�K��}���I�}��!��/ ���\�����)\�����Bs����2OO��(|���i������{�.|J���5��j}�7��b�w}/��rW�����y)�xy��w'��zC��]�o��9'��G �r?�G%�d�\惻��q�,v�����u8��9��ߺY�>��/��Ҿ��X�u��5��ySӬH�<����M��~�G�Լ���u��:��]���/prN��_�A��`�P��A*tE��Ho���R�)ǟh;��}�������^�����!ט>Y/�w�}�SӬw+�du'$܏�X��pP}柸�����������]�-�������sG��/pv{��~�<���~���1${����/p����I�:�)����Ѭw+�d~:��}�ah�����������~D#�@0�zL��y=;�@�Aѭ���#�>�9.��y��ry{/:�K�_,����C��c%��X�����A��o�Z֩�PJ�ew?r���Ѐ˨7���<�q�{�I�~���Bd ���د$�7������ZW��w�r;�]u��=�ֻ��/�=������^��c}8~�WB���}'��NA�]�F��/�}:���_����w!���i9// ��S%��{����`^�Ի�i^^���u�z�����x��ﴏ�;���9)��9&C����K��XjG�w�>�п]~�r]��vf�K�yy�>ҙ����~��s871v�g�>��z���W<,�Hݞd-�{ދ����\�U)ХZt9����нo�(8����Ǜ����eq�U��-7;�W�≠���Q٦M��#�b򣈒��}�{3�Ml�9����Zեv�Xw{�~��Y��J�
^�u����x���I.�⪠���O���g���%|����.A@�?A��
������F+�;���u#�������'{փ�����z�y�
�tM����>t��Gﰏ�������^���y��]�#��/[�M+�?&�����/#%�������F#�G�{�}��������J\���~������џ�x��0������ۃ����|���z��z��s��_a�|��@����z
p~w֗#!t���~����8>������%x�����T��������>���u�'3�N�~hJ�^����?J������y+���?K�=���4'�}�����=��u��y�`��?�F���?W�,����}���G����!��/��~��Hu���w/ ����/Ru���NA����9+���?K�(Ns �>AN��P�}�J��d�Һ���$��~�?S}��;��䏼ť���`��;�����r����wy/r�>�H}��;~�\���?>oO&���oz9.�		=�ۺ��@���?C_��gﬅ=攤�_��G�@}�.u����KK��<��bnW�����w)��O%�M���c�y'a������̕��߹���3�b?�� ��ȏǻѹw�����d��ބ�<���Z�W���z\������GF�7+����܏��yK�7��t�e*�uvKu_������}�}�/�rN����R>N�ǐ�rS�y��w/�����_����{+�z��%�^F@�y/��X�W���~g=׾����=޵����|!�i�}�e�a�� R�~�@{!�����<�7�#��S���;���hܼ���|:ހ��=��.K܇��>Y/�w/�����ԧ���D����vӍ��R�e4�� c�kP{�<��K�*��n!<;���{HĽ�u��uK,��p�W1��D�[5�]���+�x^�ѹ�V�����N�}���k�w\�e���	R�ɓ��ח�Ap������<;����������p�NG�O����V��y/G�h`ܼ�������3xr?H�O~֞K�1�sF��^��;���?}�|s�b�Z�?X2y�h�#��~���俤���y��z�<����X�����V�r�2��4���do�GrrL���ܜ޴r^y���֯����k�{�/a��J'���g￾���W�?`�>�w��FK���k�O��z5���GA��R?_��I�w9!����<��`w�t�K�;��#��\�����sîw���<���N'5�9}/���u������ZL��o��$��FK�)?�{!��?C������+���7�$6k�gs�w����}���|�8�r�{<}��A����w/R���z�{�Gq��s�B�?�����:���w'��=�r�0��M�}o�˽z}�u�?w�:�_�:�ߎ��G��������)���K�~���h仑�h��=�Խ�sC����;�zG��^������7�K�P:���y/<�ϼ�U)�S��w��7�? (����G�A}��Ss��+���O�瘥����N���{���r�=���\��:��?G|�JrN���)]���������5��ߺ�s����P?^Ð�9`��y��؎��w�wy�+�y��p��'5��7+��u/�yÜ��:��)��<�\;�w���G����2�x�d}��@������\����9Ӓ�kr�//�G�Gp�����켗ry��%n^����?H�rN����]���]��{�}�w�j��;�u�>�yé{��sI�}/�Sѽ�A�s��y'[�K��<�}�K�x��X;��|�]�9.�?=�����ܟ}�{<��#�����γ��V�
~��x���f.�!��c�wf`]2��Gu=�%��K�Ha{R�k�4Rˎe�6d6��1���~�'��N{�&<�֞�oS�X�]Y�2�����c;�n�sN��p#9��wroj�v���/ ��#;�+zz�*X���/����D������c�"�O�h��uގ���G9��7/��sx&Cܾ&���Wrt�w�˹]�{���x��X���>�������k҉M"q�뇛�v��+�C�>o�?K�8}��#��ÐR����pR惸w��sx&Cܾ�ן��u��R���#��#�����.OƿlT��������|~�?I܏����/�n=�HyK�+���}��{�9#��oG%�dO<��;���;�H{/��{޽���ه��߇�%�|G�k�b?�lv|6Ի���G�r��䏑����y��{?�����K���Wg�t/pr�oO#�_'���w�� ~���w��G�ۼ��g�ӿ%�>���>�^C�|��<���K�u�S�ܽGZ�r�FOPr@��z�?K�)z��/�n^FOg�t��
/�g���q��Ύʇ�[[�����,���<��n]˿p|z旒�]�K��!���!����~��ֱ܏�du�{��A�y/_y��}���J�+��&�ػ?W�����f���>��N���b�I������G��h�G��{?u��wZ�K�{)��'%䛃%<�K��XjW�9��>d~�~�k��.�̩�v�7�ؿ�w!�oCC�<�����y'�{���^I۽i�[�r��+������?b�>BPw9.憐�U�}�
~�� �x~Uy��{uoy��nW�7b}�}���K���7�����}�d��|�Gװ�^���4����^�}i���s�&����u�ȏ����Q��Vb��?.þ�?��A��'�9%�:4b��q��O����Z�A�wy)ٽh;�r��9���}���/R���-��}g����a��#b�)�RW����߫:S����,�/�Y1�|���JpOn�7ֶ��-����z�l�����*�Wg���Yڼ�PQ(TCo���]v�w;�ɾ��en�0�}�n�M~�mrkJ�' ���oK�k.N�����Nٻ��n�Lv9'����5��{��w��&H�'�����1�/�RPC�~�/��?=b}�����>�����փ��`���y?q�}�J�a���?w���rx�g�_~>�w�w�u�{�����^��p:�B�KѾ������9�r^FK٬�w�ӣܾ��{�r�]�I�4��/���������>���u�u̿~��|y׿s��qԿ�~繣r���zOR�4� �^~��w�����'�nL���r�r_�a��ܾ��t�ڇ��5�~_s��w�lˮ{�{�͛���)���No�>���o�;���冥�>@{�i2��<�)�<�םh�+�z7ޗ#!u�n�#����2��C��~����{��_�%;5����ߺ�߾��s�=_KܾA��4�n����rW#$���䜑�s���pP��� ܾ�O7�d=�ᾴ���?u��b��љ�9���u��g�a޻�}���z��<��Ɨ�P5��Wѹ=�r�u�Wr�'!�ﴇ�Լ����rW#$������{ǐ�
��4���2O��P�s��������s~�>�}w����K����w��b�wy/�ֱ9+��u�'R�S�uޏ#�����C��.����9'I��r
W#�{��w)��޺����s�Þ߿{���5��N��2Nsz�e���+�z�.]�컎�X�w��=kr>�#�?I����u/!�>{�����нA�>�o���k{?o=���^f���p�7+�o˸�Ns�rr_oa��K��u��C��,�����b>܇��ܯ���X��w�������	 {��ߖ#�r��]����\]A�|����k�9=B���%ߘ�����w{�bH�{���/p����M���Υ�u0}���к��8T�~K1~�H�hiO�� ��V�	���X�/M%��j�Z�K��L]�^��If��%z������]�T/���9�٣�4�o�R����]F�Ygj�V	;W;�_C������h,�u:h��Q��]��V���ޖ���dv����huK3z��4c'˝.��=^}�U��YRR�دxu����K�M��M��zy���F�8&5���du���}ܰj�E�9�";F�p��x'�N��l� ��z+��5x��x/Ao�_�P�wK4�mC����F-���,���u�"Tg�a�Msv�DS��j�$�g Q5}�>��q��'���8=��֢�k��>�^�� �tՇöq���=�K����7�rW�$�$:��Q����I���{�����[��Io00��#d�k40��H�j�#��5�b�sH�Զ?D9�$�L�uI�/�a�:�&��|���#YZ;s�[{�rW����y�B �n��t'�y��!�<��z0]ֆp.x�]%5�̪���^U���[ϝĞ�����݊��+f���w�.!A_a���(ޜ;u�ӈV��݅�#�<�\'�VI��i�RR�y����(��x�K�%�A���CI�h�:��/�m�3�\���$L�JsHx�]��x̢ANWA&����懄eM���*V�q�8&�,E�S�<�\W%e�i�2.r2�A���%�q[f��H���f���iu���I,aQu�b�n���̪������%ttB�cp���ǳFI��j�_}m]2:��^�����Tv�S�nG�s ���r��U>7������6�KK�����&�m�1�}QP��N��Ÿ�RJSͧo�B�mr�����l~63���V���P�_?d���5�]�ӟ�e4����M[�Kr9-���re�恶��7P�Z���P�+)r���Fz��]HoPܾ[U�l/�ȃ9��w��õ�}-Y�ks��G]��^R��Ԙ�:}{��VT�S�o�1N�9�u�HL��%�N/Kܼ��JS��j�-Z���86�����6�jҊ�<X�Ti�������Xz��Kʀ��^�\�i�6�maW�7�5�2@���j3D�q���t�ѥ��֬�������wv*��Cyz�*�W{�KOj���F[�Y,�-,j�:�>ΓKTk�F�;/f�;��{���o��	z9B#�*�=�U�t��lJ!��Y�zVc0}����n�86�A�>�v��I�����=�pl�;Bn�M���y��[�Wo�wWl��Nx�ʗ��ъ2�q=՝X0���;A�9�ii���/�6v���dlv ɷ�<	d�J��A�,�B`&b�\gJ7+��L6�I��ٚ�on̽�N�8.�̍LE�s�SEm�+*���f��YԳhm��n���k�>�;�bR���(�)�Ū���(��!��Ġ� �� ��ȡ�ɤ����L�'*�
��

���G21�%���ȳ�3 (��0�K3&���\�L���1��l��Ġ�0"��&��e�ʩ,��+'1�2 r)�
b
��&���&��,��
�+1p����0��h����hL�,� ��,�)L�,�
��Ƞ2J�(�,1L�"��&�S$�p���c02*�s(��)�31)Ȉr�2(�J( ���,��2����H�%��!r(��2S �(�

p�J��,��2i�)�* ��� 2L�r2
L�,�!(32Z�(,Ƅ�r�ri�r�s0b�~I���RDw7��2�5d���dB6�OܖYP"z����
8��.E�I3��j�s�<wS�� �1k[��[�|tU�W�ם��o���g��B�=�Y���<�d<�q�ѿt�����ԏ$��Z9.�${9�n�{}/�w�ܯ�Z�K��C�}��d������w��^�7����5�w��{���}��}���ԯ�nz?`}�z�A������M˸��x&@r����w'ގK��~��}i_/���Z]��s�?u�~���Y�z����[�j���s09/!�zu�{�~��a�_`��~��~������r�2C����9// ��L��~7ޞ{�����ho��_�?y׼���z~������\W��<��J���K�{)F��w'f`���y�R?C��N�~�>�������<�r���iL��u�~�����:����]��؟m˓���ô��b�9!΀��ut�f2rN#FJ�<4{ozaM�mN�9��&V3����doqs�5у�=�iK��WZ�p�nU/G�\�ϥ_���Jڗ*0:vJ�x�䣝3b���)�>�g���R��S��9�%\x"��!���nX�3˫��9r-��o��&6^X]��S��I���v���,	���u�/+Rev=i�9����}M�~�r��;��ܩ�{ʛsw��K�V>]WFƅ*O6�e 9΀���������k��L���6e��n�7�^�3_�`X�I��c
����5o1�	��Q���~���T����t�y|K����j���SSү�2;i���w��� ����T��[��<.�*�ֻ]�Wui��{�>����n�6�o�C�ls���`��y��n����v;^�<��m�;麳�;�{ۚ��0t�k��͉1�ϧkǣ{)����̭�V�wA\�����s�͟U��:���H��c7=�WzI�Β���ٗXN�}�Qb�=���=�>��c �k�+z*��f矣[ͳ\�	��y��C��TQn{�����xи�f1`w�Õ�XN[�Q� ��ח�,??�C�Ɗ��!��h���`/S3����\7�-�~r�s���~�:��[7s��d�{��C ��]N��`T���1'�l+���]{T.��tV�����ov=3l	gh�/���3���k�C�!�s�Ӏ*�U߱H|��}
����g����\'�o�	gh:!o+�t��>��;����}[�zOuչU��qo�/��ʉ��I.�g]�.�tC�AK<���nǱ�g��Z 8E�_J9O�n�[��(m�Ӥ��S
�H���/��oS˭�����]�'����zh�la�˖o�4�N��7�cy�Z$�oV�u��hé��f�cq������Zkn�ԛ��� Цi��U_}TY��]�l��ou�΅�u��p������5��1��ْ?��A<(�nO>�.d)��s�O}����cs�|��cU�>{Ϊ�֋xs������v�y���k9�\1�ԝ�۫�U�`�g<h�mWS㭓[�W��^��m�.��&p�/r��ν�i���Ǿ�Q�L�)���MI�lH_�g�v;;�2�w�����8���p�/`�����vt��tӮ�bĘ����X�6�����7���ENk=ʓ�O�����n��ڳ����)g˧���O�يu�[��P�z�縈��Bǡ�V��㜫Vuma^�8�mw{Q�t�P[�'��W��?u�b�S'�3�W�i����J�����pV����a�叅;�:�e��@�5��G��N�N�^�i�l/�̃����]0��c{¸S��F��e�-����ݹx��)hnS���zp�;�B��:3\���b�i�9$c�lRN��w�w����E��no��������);����_�f+�v����˦��<��\��B�Չ
�������
������}L��2zq/O�/�'Fd��{j��}G�	ȫ�=Rz�����a�V��݌`��8�ނCs�W�Ό�|�l��������٧z��n���G���|�t�7�o��(L�w�Ny�q}K:%t5�R��i͒������!��q����9�N���k��N���[�~�W²�m�\��նvJ!k,P<��C�|]vt�{7>w=
�=��[���Ha���D����`��a�n����h.}h=��]��\�X��˓BAp��N��<�x����%�Rf�����Ɠ�W�=��~9�Y�^�;��t������eɑ�����֋�I����P�{<O�����OM���}7��PW�k�=��%��&��_�Kbą��wO���¯i�/�x�7�y����S���y}#�!5���&=&�Z���,�;���-��-.�ۈ�9�W�ht��`�`/n����T�S�)Av�p.�D��G�W��}�/X�k�V
/&ԉ>㘏p��un����a�I���7������1�۞�n0�\��S�o1Y!���;rk�'諭��� =�Ox]��q�εs���f��ɗ�F�?oϽV-�,��j�L5�I8�{/M����g������6_��C��r��'�z�I�¨V/������*�~��ٿ��nǻݛ�x��l�	�и�g4y�/t��ؾ힏�&�����ݮ�����Y<�h�`����e�m���Gg�q�YF>m�b���=r�N\��?H絋���Y��8ׯsjK�}�%��s�>s຺�޺�l�|3�c9	s��\g&��/cמ���vV�w�^�zK>�
ˣ�]���䵨��M��L�2<�Yl�Ɛ}:[56�<���^���ӣ�x�Gd���u������K^i�Y�%Bm��Vw=��s���/�s�!ξ���g�N��Jz|���7��xJ�I�/ �&V	�vN�[�\�{~�v�%��VyiY����u���8��������N�U�.�dǚ��]���e�<�"�s��<���.�w���jūe�7˃�[\$ ��z�ݡW3;{`�)�'s��	��T��Q�ݻ솢H ���u0����9�qfB�0��k��ƭ~ ��WW������3����'�l�cbU����K�ϦK����ɮ��~4Ammf��|���
4O��
�[�e��}���<�EOp	h������f�<��7��T�c ��23��=;��@���&��������W��J���=���T �<�<���2�Os�=��<y}$�5'����Qq$���٫��[ìf��s^u�Nu�s����G����l�������cWN�#�(_��7&=1�����6��g���Vf�=��}gv`9'S���Ϧ���:��[�q�Y]��>�w���o=<��|/ںüSG*vl���z��'ƅ�P��c{d+\�����6'��𷻵����ﲮ����9�\�km{n��3l�,w�µ��t���Sw��Ӿ-�:�+�~��ߎl����c�u����hw�]�,?s7�g�Pi�ѡ\�Rit6�+��$0S�A�y>����Qd�Ǣ�U,`��x�Xv�Kf�E*%6ԥ�0��f��ۦ���Z�Tr &��s�^�s��m�����u�C3\Z�+�H��ޫr��Kג=}�����Zy�7:~ ��|��=�g�����>��y������3���_�Wñ��a7Rӻ;.�ǃ��\�6g�os�=�Y�tv���O=�TY[|֫�W��u[S����N��ٳ|������Do)�A���hwO=>�F۷� �}}O�y�5���}�=�.��O�;:$6��Ya��r^Ow *SC�5�t���vt�L�u~������%�SI�/�Պ�_�^|�ʻ�K#Y�t�Ok6'w����%\w�E�O�w��3ݪ�zr��*��u�_E��d���%�S��f���:�w�]w����P�U��}~zt��ݟ5LX���m˩<&W��=�]F�N�վ��kVg^�[�8�K�WGۭ�/��+�ع�b3�I��8�D��{�Ww���Y;g���oW�l�%�_I7�O;����1bLzpt�zE魞���na¥�v�{�%�y3���d0�Z��;ڗq0.�s;�4�w���a����9���, 6:v���i�^'=��^��{)'�ѽ���*p�st�cs�W2��$ӹ��՗˅�׫�`������[��"F[c�ةx!7��Z��o�������_n�h����jg�-�g�?}��c�5���3`Oc�>��ƻ&ȅi��Φ��{��=�V����������'�Wc>�w�E�Ani�c��2��V�.���'wv�{��^��z�/����)��8o.'YuA-��ޯu���W�{5���\���U�:6�;E��2��P�� eɵ����"����3��G7��~Q�2u�Uj���Y���~ah��ٌ���M�Ǡ��o�1!��)�љϘ�W�ϵ�c���{�)�	���<'�>�ޱR������o�S;]䏶1�r9�V�#f��fN��h
WX���<�B���y�c�����췩�x�)�ln�] �Yr�y�D�����}:J=�l��g���o�n��3ُ@�x�E^v���ܾ��Z�7DX�a�ݯ�]��xuD��͠�ﮥ[��Tt��
N�g>�v��>�g>��y{ţ�qeČ����vGO�U�5`	$uo;�=}C�2x�:�|��_n塹^u�3�:��z�#�V��X����vn�C�@�kF�ݷ��}�Z2V-���-)7�����j)µ~��������aa�Fp���%_�R���)3G��tM�<h':��/E��g1A�"��_O�E�����|̱&G
~�!�$��]Gd�B���;ܾٱ#U�t����+ބ�mA%�c����b���oZ�3�Y��ѫ�p�\��`�+3=��wm��ל�q�7��k�zkV�tgGS��0O���ǃ'�tW��qZw�J���ޣ����17ݯ�\���)fG�}��|���ݽ��e���T9�N�/=�-����A��M+�[�*d��_��3=sޏu����ƙ�^�'�m��x&X�7ѱ2���~�f�'�0�\.U��ܚ���[U�g�����\�Ê��Co��n���[g���p��,'.q�:G7�g��u�I`��_03�y>�v��z�mP�m�����.��~29Ӿj?s������e�l=�KB�ZyWM���x��[}���	ۏî�ҥ�D�KK��d��U�*�2�����<��yo���m�.m=x�wF/Ok���6ڪ���8Dw�-h7O��xv��z�G��.�� �m��;P�ϓ��Ύn��� :%��:ܢn���Y���]L�~+���a���O	��g�*�gB�gf�c�r.G;0�m�;A����b��%�뫯�r|E���~�f�ө^���/<߳�e`;�&�D!�X�y�C�q����*u��N��J�=��/Ow�N�9�ԓ.g�����V}� ����,�kڌ����r�ԗ�g33�\���j^'�Z�VӷR`hm,�Ƀ�A�;�z߹�&|��Jl�����}�c��ϥ\x"��3x9Z�������ٴ��>�(��{/��ʱM}{~��t�n�c��N�;~���˽�n���h��z�����^89�=�IG����w��||7'�ݝ{8�`ɠ����^���{j=����H�W��eZ+���+��26�V�}snN�=��3�c�̬��l��+��W���1��k�(�eO˒S�0l}�r�M�D.|���)2ۅ�	 �vQ��e�G6���E�׻;D��D�۟��x!�.{��_pr�Cl>x��2��O�l�m�*!/�!�洛������{s"��u.\�xo�/��D��9�]��{��<��@"�A�P���q��u�=�:�CW�b�COspԨ���2�V�Ŷ�������{D����	�6��\�A�2�q�·M�B˺� 6�����ĳn��%,dk2r�r�l|�喷��B�Uu�f;�\���N�:�T���9�iw�psw�ۜz����{ߏA�WH��GY�Z�o_e,�k�Ŗ���u���s���{��!��@��[�/�a"����U�cM�;�vi�Тw����X�Ơ�˧�4��C�d���[�P��9icӬ���ވ�\7'�<]�bK�,�S��E��p����|�J�s$�v�ƟId������u6b���gWr��?4�q�n.�.�Fgw�:�E�W��7��9'���#щ,�F�x���;w)��[b�ed=6�*KT�:�{�YIڮK�Z��
 ��}t3	������h����ĸ	���J=�O�M��veZ0ȷ��e����9���v�4�L��{1�?$�9��&)���|�}}�Ӷ_�kJ��2\��u���uÙ}�S��`Kq��W�:�,���4���՗�L�'5�h��#�$mmℚgB�/���%��������cN0^�3�wq#��,�;�
�Ww�d4�¬���P��p�� ��^G8�l�w#5ݺ:^�¸�Wt6\B
�f�T�[�����X�Ϋ��a*����`dT��Iq��Evh� ���	��/����oNc�����;Μ���/��N�a�۴{
_3]H�Z�>�|��n"��`���K�;d� 쀿w&�~��o7�=G�u����g�������0��0�׃5nWx/{�E���jm�y�x`�]���4��{�\�ؼ�ͨ������o;����!޺��)wq6&V_��M�����2�R���ߙ�����&�1M����`�)���:���[պ7.�w�F#5��"�=imc���u�}K ,��i��U%J���{�� �Օ�j��>���}�;g�ۢ�tn1��3?R�<rRBV�����y������7"x��W'���\��ΰ��9m�5φ���h�CT�b)���J �I��w���;��2�Sx�*Vٝ��0�Q�75�OquY��_[1 �B��!Q+���6�8h����٨ͫTb�x�s����e!��i�1b��%���A�5��q�ݰ�,#n}	��sy�v�U(9z��2��p[�*VPшrY^����ܙ��'��,ȡ�[�^��]��䯂I���@v��mbw���w�^���tTm��������1+##,���(r��ȡ�)2'1*�
�,�)"Z\�	 h(�s0(1�ƌ̥�3"L�ȡ�*(���l�� &�����1)��3JJ�0��ʃ$ɲ�(�l�2��+ �i+%�L�j���hJ\�1�30������
rJr����\̦�#!�0i�%��2J�,�!)L��R�&����2(�3��1�)����2B��*G �
���32�+ (J2�ZC#���,c"�%�c#%���3,�h2��'"�L��!����r �rh0��,©�2s0(j�Z\����,Ī�����
��@̬31��3�P����0�,0���JZhbk �,���Ȥ)r��̰DGģ����U���wܹ���Am�};yfv�V$^+��%�ʅz9���Y4k5�׻ٻ��0Q^�vW����X�.L3���߳U�Y���2t�ޜK��]�{�!�Y��	�N�Lb�����C�Q���Y%��^�Z�/3��6'��7x�bW�Xۣ�:����r
�!o����a����V�\���C�҂�>��v���=7��)�z���c6ˆ�x�t�BvuQ���ӱ�-���Ϛ��&����gh�u;'�>�Oa�JE���i޴���,�ul�}4�&���Ǧm�,�|��(�~ۺ�C��u��c�5ӷ+ko�f�����L�w�f�`�����U�k��[u��3�=�q�>2q�<��[\W4��ʨ�nmd�o~����;�Z�^�~c����b�7�/�Q�1�T��mq����crk ��7lk>t}�=���]O�%ؘ%dk<s�ө=��>��Ϝ{El����|Ϟ�b�!V��`��N�wr�ڳ%$[�-�X%r�F�p�0J�wn�fշ-��w)ȎJ;�8p�}r����К��?��!Q��t���r�OX㯴)ֳ^����Z��������}&�ę��z5���,�vv�m��W�  ����.Q^��U����'�X������ʺ{C76:ƭo�kW�%��x��q��G�*bą迤�r�κ嵱|{-qꤙ�J���;�\�fTZ���o�i���T�� �=8+�Ϟ��b�i�o�0e�WZ�Jc�x<�Wn��^c�ﻺ�}�4���q�I�Ntm��k��V;���g�4n�����Shx���e�ܙ[�z?k�R]�+&=p��g�t��ٛ~����~�Eƨ�9x�-�z�؟�G�Izre�NG��Y{��yѷ��$7<�o��ՙ�=e�~5��@va&M��E��H�<����FL�s�Ot�,�em����٩m+����w�3�������<c6�':cR{=;ە|����޼8#�9�7M��o�v|���\v8o�Hg�ߛ�1����[�����o��[����#씧+�����̑z1��]/ø�nK��1�*0��?A��~o�St��exM̔D0�b���U�ɏ{�(i��d��� Z~C6��f��[]�L�[�Qt�:���.2Öe��c���T��k�E�-4�N��LT%O�}U_}����]���Q;��>��v(��l�ܞ��T��x����n����<<�-��Yu(�X��!΅�u�����J�k=�Lu*�TM���ɧ��|.N�q�L2���y���B������i�7�'���w���@�����v����\�a�vB�5���=��Ã1yJ�N����sjt�mK�s2��KႤ��a�&��4�!�j��S^��'�K�ɩ�g��3���O�$5���m˩{�۞���c�[珦Q06^Zz��^׭�k�a;�r�3�Aʽ��97r��&,:�%���X�q�w���.�-���s �������ˆ�߽9m�_Vfێ����n�QR���g�j��o�{*��z��}'�A�ҋ�+ˣ�?j��q��ْ��ǻcoe�a�x��i켷��:v�������:<O|o|�w؇�u�ɻ�ëE?��!Ʈ����Gse�x�zz֋��F(�΢�)T��<�K�`�������z�K�ޅw������}͸W�H4;�tܙ+9�p�c��d��jY����m-�lF��s�|����,�~ �����lw��f�����8ϻ�������k�&��V9��^/(c�V��S�w>9F>��L{���r�r�q�Mq�Of��6�������EZr�����ށmi��v�b���=rӗ3�Q�$s{���&��5�#��m�^��o17���\�Ӱ��p_xs;���x��
l�;ٲ�Ys|��|��������X]N�Z����Sfؓ7�en{�n�c���d�"�T�����A,�Gh�b��is���2�K:����Ss������ /�=��߷�m���㻘v���,Wǜ��gQi��W�Aѷ�+��9�y��N���RK�{M�t���72���˧c��9�L��7a	�{ɿ>�J�qVv�/rI}R�%�o��-��Oe͎���J4��]=��л�c���W|"��U|����
�ёb���5)YƐ�����uѡ�v�������	�h㋷��)�"��whv���,�n�+m��ى�\���!d�[����/{����N���Hl���M�����j�k�����l�|.e�s|�4���}_UW�K}W^��Y��·~vJ�e���N��N��wcvA��J�^n�k6���ld���9���S�w�K��e'������[�J�=/.k{-wZW��|����!4= 5�q����z��_aǣ�4S�U뭼��t�w�1��S���z<~��m�}4����ߌg��_aǔ;g&��<79{}�1(V�V�5gE�yյ~Rt����)ѻ痥��9詾W��f�����#��a�d��?gV׶@��	��n2���]�'_z�3��+ⶒ�D�/���!y�}�u5� �_0�I�_��w|=�e��e�@s��g�Ⳕq�|��z�Cl�P�c/�k�U"
��u�EG�Ľ6����5'���|������K�9k��
�����V����H�	�Py6c[ݟ=3nY���Gh�����̹vy��8�j���~�<u�vƇ�}���2��:�CNf��`�ܩ;`��'c�\��@�3�Vf|�.����`�:��ԮŤ/w!�7�Vk�P��C!�ڝ�����zGT��&b刡�I�1�36�����u��Xk��p�?���ݓ�sy�������:��:<���N2�o;ɛ��{(�\z��ڽ�T�y�"}�,P�ʣO��N�-�+�\�g�>ܹ&X�5j�k+���8\�T�K���%��f���t�.�gM�������z�dX�SPd^�.n��̿S�=S�������#Y㫧R{���^v�k�ƍ�=>���Ϛ��J��&�L�a�l�g#��G���n�N`\��%����]�[�����m&�w<ؒ� ��$5
v��va��H��}رgǒ�Щ�N�y���O�a��u����菫b��sJ�T!\��kW}&#�4�!SO\�*Iâʴ}J�3�,�yZ/����ڔ�;�Xx`��2_J���KJƵ,=@��hKt-�脛iI���Ek��,q���~�UYg3�q3��h�.:e�s	�v(�'z��32��G0�'����n��u��[K�t����F+j����/�p�%o�� �r�� :<��j�.΀L��׷(��{qo�iݴ���X+7C���,��kN]�]�)_TPm�]��J��j���A��]y�̟{�K7�ܐm�~׼�*��X&~�m�mͫ��)�\ʖ�)�����������'3b��$}�b�Cڂ�b����>�� ��\�Ȝۚw��G�6�����o��{�+0&8��x��bK�����d��M�v�7�ְg!ܢ��bu-a��z�k�F����(�Bc�Xϳ����H49����\��I܎�a;y(�u�D�=냳�V���K�x�k=��C&�r<�	f�wK�Z�\m���,�o�	>h�
鴢fr���=�,o'h�k���Wn
M��gP����-KA���yJ���E�;�#�g�M^�H���g���%{oN���fzI�=Vg�w)eШ�5�\��KZ�B���v��KY,ʳM�OW�������x`q����L񸃥�L�e˴�x�|�5��
//�fK�o4��i�'�{�I9����ǧ��cHn<�<2KƮ�3}2Ɇ�&�R$�#�����rIY�z��Nt,g+l�qy��ds?	W���
�KZ'�.90T70�4�my]���A��}\�$����k7VC=��Y�qeEbOL��JV�IBj����ͯLZ����-Ӯ6a�mS��1�V��Q7/�Ε��G���:��j��r���N� a}�Tx��9,��'%�w�Cd;�/�nd���o%�b���@�l��ۻ�����q�2G�u��J�<���Y���Biu��a�&��_UU}�;�yg�7����e�J��GY�K�H��f��^��5ً}�-%e�X�1�� ��W���w��ˡ���GK��7^�m�g�}�Y/*�>�^
�E.��|2��b/�'w���gI�z �l�*�,��倱m�M�氣\jV&<k=���i𭢞�ᝇ�9�顫�^G\]�։(i���(ߜx�}�e{�
c�^�[�֕���0�ݯ-���E,�{���vF��Mځ}����g��;�aC~]3�ڞY~�1��W�`����d/�Y��}���4>�j��T-+�3�w����2�É9v3C�^�k�_-��6���}����,��^�I�@���㖷�3�~��*��d�";��F^�br�8�5f��\,���ۋ����=,n
�MYEEb��<�Zf��N$p�����E�F�=a��3s�-�Z���?�>���gc5��eC0VZ��!�I�y�ܵ�4��"����b��ǅ3��FX������m\��w�CɘCG��K0�O����<-�{b���2�S���!j>)��辴�|�7c[��#�G.��Q^	���`8[�fi���l[���;V��Z�zH`����Gշ�g<�c����3����'V5mk�NV{wn�Ოe�"�/���6��o>����g=|t+��ﾪk�z���w����c����3��v"oX��_\j�t�6�c��t��!�'5�+
�.1���;�<`A.��c��jiy�4���,I�=��]p���<	��zB��2v_�'� ��d˸&�#׼�<tmIU�b^^���W�E,��r�T��.���P��o���ϫ�6��i*��t�J�:���z��K�޲w}ˋ�%���A3m#s�:�7����9����"���I
�k��\e��p�uf��J/+#�oݺ*�v&[����Jh�=L�������!����	�H�s��h;*y_ԟ/o��C3~�S�;�$fcq�K9���ߛ�I_�� (��B���4�.�O�Y��8Y�����#�����}�r�y�}8�u�&�~)¼���Om0>�ms"Y�՟G���ڄ-R�%�N���X�^w0)＠�
�2�/	{w}�x�5��lpX�|�cK�ػ�Q�bVD��/{�K�����Z�k�?m��+ypʇ�#���"Ꞿ��ة���y��/tm�ؘ32_#35�0HܟM���1��Fw����e�بS�;hc@Rm��Gh���m��1>ǳ޷QPǃ}�u�t�+���oe�!�`]�.�ju-(3P���0�t���8d��9�nP��Wa�N�Y.<����Z�|��OV�M���� T��3jIgs�ѷ���Wrsl��&�!
�´ݺ��\B��B� �&�#s�'�M�~c�珴�{vv5A�	M�b{nWH��f�$v��^ʃ~��(�p�(������*y{��&8-�v��2��3�HmOз�����Zj�N�;�B�2Jȴo���M�|���įΌS|�F��ڇV�J�3�;5�rWaQ��w�'+Y��	�~��&�ا�3���q�*;0�D�f�4y�ڮ��"jU���6�?`���N�J�ݠk�)��m��Tc�n�o���z��i�\�ǇԸ�Rv��19ת0tO���!��v���rQ+��^
̼����l�9�xz��YMD]y-�]�j���9�����,6m�W%�
]]S=�R�>u�c]�E�l�#�a�}+2
���_#�.�Dÿ$�����/�׼�H�qS�xo˄۔�uᜠ���D��ް��Jȃ�Wl�CP����lL�0�v_V
�n5�X�g"��0����;z��� s[���/+�z��W� FL���.��ǰoT]�hˤ�G�9e_a}وP�3f�g�r;F�{�nq�JH3�R�g(۬��;����X�8d���<���WvY�7�Σ<:�X�7�����b��)�#wk�[�C[��$����M��a���1c�����lv�<J��-�WuΗG5��~&�J'H=}s�~��zt{�_�7B�9F�Uʝ�����3Y��]G�tm�_�ܪ��x�e��jRw��es�u����*�F3�Yp�Z�8��f�L�v�uv���E���ɻ]2��yRv����9鑭u%�x�y�wm���w��/ž�{�w�o�����Z7!�s��:��H��jm�.�c�Y����v���������T5�aU]�)̶��2��<w��)
�yە�h�d�/xh���0��]֛�=+oD�msdъ�3�.!oD</,���f��S�dz��$4Y�l�L���b�Ho.��p��0���DG+*u���2����G�\S��_QW��s壃+��ݻ��;����aT���әז�ֳ��K�%Az������=��0Jã%�Q[�%�n-����+#�\w�F"G��w{�A֜W��R<����iG�h84�7 �s����ݜV���X�9�/����7��faɁ�A^���%N�e���ԟr�w��i�Wq�s�����܉L	�+�\w_�:�΁@y������j�R�&PI���ր���^{:�T�x=�p16�i�C�F״����E�qg}|I�<4{��ؗۻ�P\�sq�~5��嶮9Jnm�F���z�S��V�=
[s��8�cf���և��a��sT�o\��r�{]�����y���+�:��TB�wO&VDv���Ù�p�F�I}��1μ����Q��:��y��)9j�:���}g�%��K6��V�Y��z��Z|y\�d����;K�o-�};�Be%��<̋����->y1��:��J�isT���)�X&[,��v�Ɔ���%���' �9���yM�s/sMj�Ra ���Wt\Yđ�/"y%ƛN
���=�՘+���<x{�k�$�]�u)�U#���:����vp�5��eލVՊA~1�ʍ��j�z��\�_e�SZQ���O�m���bS�~�u���Ny�{oxۤX���䮳����Q�����C��$b\�ڽ�o��kF�w5��[��K�ݎ[����Ӳ<�&Χd���(���/DF�+R��y֩��.���^�����^�*/1<@е|v�Fⱉb#��5��U�J�sS���ʡ��2��),,�0;Q�Pޕ˺��H�o��E�	����%��ҫ�ۆm�n��� ~����
Fl̇!32�p��'#*� ,�̀��Ȋ�(����*��j�
)�2��s12(�Z(���&�%l�"`,̩���$2�2()����"#0Ȝ�#!��+3&�f����2�)hrȉ��s3"�"�
r�2�

�
����L��3
+,�2b(�Z

���)�!�2��Jp��
j,�d��ȡ2�*i���*%2r
���&*H�
2C"�*�"�����*(��2�lƚ(��ƀ����
hJhK0ȋ3,�2ʖ�i��&"�2Z�()

�"��J
h����$2 �(rh��
�3i(Z�ɥ2�3ȣ#,���$������k,,���ٹ(�I'�����lM<��L�X�9�ԞR��֡P��_gv<y͛A��y�~��.W�;�s|6;��c����}�Xٚ%_�ؾ���in��1�T�A��sh��%�G>�w�HG+�{E�Y@W�*�^�����g6�K�D�?#{)��=�,��P��&pXV$���u+��-�}ຆ��F#4�O���^E�̖}���Ϗ*�P��~����:��3s�mP���3}|Na3]2H��-�^�����&o���d���`p�.��g��,�`Ӽ��#�t��tS�.)���<Fjų��ױ0&:%��/:�ٙ�}b��S ��:��,x����8Cby��2��^!���u2=.X�L5�x�-q��h[���B��cf+}�-����Mz(P�4 ;�E���+���s�[ET,R��1\{���O>�2��y�%��-^@^�����c�Q[S��Զy_��+�wL�ȕ�t�C�֠7v*��O�g�/>�\^}r��;�9���ɴ�����z��+r!�� ��6u��~�_�T�u�6)	j\��)����2��s�r�rT�=0Z�}�c[�)�^� ���t4Co7��eT����}(q��Oŝ�^��'tN3b÷�TfaǼ���|��^�a�t�7���\�+[�;�^�e]("�uҋM�}I���z.�W}iD^��62�^���H9ppt4cr�09���|��g������p�ڛ&�����=Z��&x߄��\�F�R�!��%��
:v���NkM�`�.�k[����+����{J*걤X��
��+`d�s�&e�D��<F	)��?����/G��$W=����̎`�_�}ՂJ��]C��xT=I�
N��Xͮ�ko|�"���4�ꯚU�}_g��_��-f ��ɓ�WcN	)Z��k�n�ٮ�'μuw@U,3��M�K��Ҫ�WV*�>��=tb��t���*����x�����d���߁�t�F��0�J�"#�P�>��R����E.�`�C׳Nn�.>�75�k�{� �Q�qm�Jd���v�M�X�|+LR��Գa��ދy�dO�����&��^Wj�L��=(i����ǈ��Բ;��ez᳊�Vb`���z����z��˵^��]k�y�/��/�Y���N����끆2��5�X�^��ɼ�ֵd��X�KFJ�����
�S���B�Φwʗq<j]պ�e�l���b��Q��|��k[��Ӄk��������tF+���W���[Ӓ9^�Z���D1�h�sb$�z���gg*������l��5�r�*[�콐�5&I[��M޴����o#GN�Dʪ;��`/u,��N�`�,����}U�}��G��}���Fఌ41y]ZXcJ-+~�d��5"/hBK�� ��sz�׮mFOݵ�]���v�2�j����ǲ��VF�\��(���)�C�ӉMH�k۞����Ek��z^%�?;�6���jbeCj�j�h3dm.�J�̻��m�O�2�,4tC�?skpp���w��s�4�6��⦦&R=*������M^>zpy��q7�]2-���������������DS��i��\\7��<�7�3u���� p=�2���$ǰ��^�ɩ���T��i[.
�ڛ���
�����8R
�[��	�$����|'���W�X��tڊT>i�//�q^�՛'��E-�r���=DD+/�C� �<(Gt�|9�-+�P�˸{��;h��N�cnd:X��Y��EoG�����4�;%B%'�ZHV�\o�댼��6�Pf��Q��)����&9�V^�Q1�aqW"X���rWޯ�$+���*��R��;NR�-�N�&Kt?n�f��&�5�c���W,��	D���\�:R�2jv����tXWރoU��{��h�s�W�^m٤r�O=�~�8h��o�Q�;��Y�+kg'������>���W틅���s�S{.� Ś=æ��N����U�?����ѐ�����!���v{��鑙�0%�p���X6$4�,,��f��������Yb���ԟGKз�-f<��f�y�E�����XԳ\�9��i�-�Ӏ�Q~:.�u��^��FC�=B
��	�Ep�W	x߇�m�(FP�T�YK~�M�nդ3^)+zxeo�L[v�ƴ���C�V���z����Χ��Go�E�u�/���Ֆ��O:8���
��1�WL��~^J��KH��yz���`�Sf�r����.,�n���&�I�*u��wf9u���'dn櫃�{�!�u�,�5��՗:+4�#�]t���h"�ޜ�i�Z��̿�����c�j��;�ÎY*��pGWF�Y8����=ӳ�T0��:��ļъt�F.mA><�MJ�
��n�k.�]���譳�3܀�<|��`��1%^i!X��`aC<UGf��a���Zs�Z�,=͗nZ(qu���5��b�\\Hf�wf�U�9et�sP�� uuH/.^�ϰv	-z���⪴m�(��8y��$��+�8����7�'�N��u-���yf��\��OF�|�.4r^��*N���7Yr�T'�˕�x�wx����z�d�]O�*1�����X�o6��f�;}�J�UV�n����� >X9{����'٧?d�9Kg�2H~wh�W%���ϨS3Jk��4�o	����V��$CX�o�d:�3<1���F�=4�Q�1p���{w���Y���W�峵n$�ޣ�_ϝ��+0v|�H���"�Gˇe�#�$�=մ�P������j���s�(��fWC��t>����s���+"�Ev�	C�>Pò��{sL��zߓHev�f�0�"�<g'��\ST>߇e-�XN���*���cy�ܧ�c�Ah\�Ww�!hzF�zf�*�y��>�~�;*���}�,��\E���!���+��ݷ�����hz��^�x�˴�-���Wyr&w���0q��ޓ���0�w�	T���M��T��ׯ*nR=7����61_#�[m��%垖�Co:3�V��^֖3�ۆ`N+>>s��Wi�~���`��1�/����^D��xvT���Xge!W��fu+Z��ٙ�;��C��0=�7�,a�0(=�����Kc�!U�5<�=2�T!�)��<����p�o Gf����>m�w�Uў�o��˗]�YjS����b�1�Rn�����p��;\�W�tY�=J�c����H�WVa�r[�����o�T�ˀ[�����S�+����+��UW��)d�l���Z[KR�O�pP��A�c}E�w��/�A�;�ȯ�c�����(9����My眲<CTh@�����M��U�T�}}P�gQ-���(�)�K��;Y)������w�S������X�U|�����/>�\]J���ȑ�����9j��}׌�6rwEK�OC�P���kM�%�Q8�����O]�ٷ�xr���J\�1zd���KX�%_G�v��zMC��9Sl�uHGH`���SfUx�ce�Z9��+���~w5E��*Ds���2q�[3�����,�U��ӵ��f��,�~��>B��o���/5�ds�����ՒT��.-�,�J��^xs=���nF���%u_j_q�g��[�-[\Y��Ɂ�Ev4�>���ô�epp��yHʵj�����&T6&RJ�JE�(��ڠ��dO]����$������&q�w�'xpMU��Α�)y;���E��u+��\�]�4WuA��w��p��k�Sm�{L�����L��J�7�9��7F&�X��P�/��u�U�yk�0��ܗQX�f`�����n�k���H^���^�e�jE϶�iށ�g2s���a�ۉ\�n9z$�c2+���lg��ͪw�kr������K ,G9"�st��6L%_ɘ�6$�I�Ү�h��!\jV;��g��Ŵ�9g�Yf�a�O���BM�1���O���X�plyǈ��԰Gyz�>�}����I��K#���r��y�GĠ�m�4׳*Y�zz�{)C�`At�%��[=�P�㲱���_���ོ�Ǝ>���[�0UC�X�P���>{\Dht]�3���1b(c����~��w�L/�`�aUY��&x���1�4;H��!&�{Lţ��'M��o��5�>m �Xښ�׎YҾ�V�YXf��M=A�=		6�,�q��ϽVz.`.dϔϯ��NEl��o,�PںZ���A�����P٧G�(_b�+3�}W�D�t,�(���=CH��o�>*js)�H� �^{m�p���t��yߙ�U�A��7���\zD�O��o�/�Z���{��G0��n�x��e{پ`@2��A14�iڗ<��kL���'9p�
k��P;~�u����5�����¬[޳�2����b�n��I�"��y�%��2�v�J}n��v�n�F�H8ܧ��ge�ڵR_rgfk����|w���	��^6`V��+C� ��A��c��N�3��Rc[�Eb�T�X��O��an�n���| � c:WH����������ΔJ��f5�P_R�lӊ���A�*f� ���9o|�#~>^���
9�ʘ�xPvZ49�-+�y��=`v�&�����u:y^sʆT�1��ʔ��sG������>D��,P��$0k5ĵ�^��xu�c������d�m�{�3�^Vn�2��/%[D܆���	_z��!���w���QK���(O��^w;<�l�m��=�L���0%c�<���X6$4�.�O�+4B/������唖vgs!~�k'�x^W�����y�v!�>�5,��9���a�r��Mly��p=��/}��G*XX�(��qpu/$��}���g/�8,x�w�n^e=pU{�i�u��K~-b5��iZ0zyptC��gV�����͏+b\�H�}�;�lT�vFk��Ms-�ܲe/+�6K�H���)��y�֙R`�'��ߣ�v�Y`ϋ��,��ى˳����#��S=P�����¨�R���s��b�ʆe;�������F���@c)8��z���4�[Gv�\ҡW=x/Y�0���y�N5�k�Z%ڷBpj����7y˾�Ƿ�`������=s��s9,s�� �ć�ߵ#�K6�N�1B~U�l���%�┒��W?S����|x���)'r�B�gn�5X+K2�;���u,x�ڂ�-�24b��GZߵ-����`�I��"�ACuq�h�ɶ�9T:z���U�NO���K@�X7�v�'ݢ���3�X���Ժ�#on�����MS���<�Zc<��]��B�~�����z����,K45�#��c�\\X(&f:���C���׾�F�сiZX��<|Af�'�>9K>�m;�j䡵��A37)�6z����WZ�Y�J7�?̕Vf	s4�)7%ޛ���Ɓ]@�ɋ��Yp�~93we����l:Ox�}ug��I�6Zh`�X��Y��5R.>2+�jT>ٖH�D�4H=���ј3rf�%EO�cN����Rk2s��T���/��� 0z��B�5H�a��{Y�.����� �XD/��ʤ|/��)�Y��m�L	+��
��1�ϛ���.�T��� ˘��i�Wv�����L>�@TRg�.�,vUτ��0�r���X�k�$�'/.;�c1X���7q=&�r��pA�<��yb��0p$�8�:�h؎pY�B��Z.���u��^D)��	�kv�^������=�ݜ-a���-��"Wyz>B̓^]�)ͼ��{���q>�Q�8�f/�}U@��:�Lp�z��α�K�>]�P�J��D�XyT�I�?7�x|�^Y�:�^MI\��3��l�M�:��re�c���+�֋��Y�m�Jr���4Ay�O�d�)_`W�O}�l��qY��ўCؤu�q�������6�z�u�����D�}��Ɲ�t��0}�!�J�fu;��}�q=X=�5VL�j&^���C.c�vK��B���X�ϒ�?R��*���GL;]�t9}2w3��'�ή��ٶ�Jy�w԰1'���*�a�Y<}���>��3.Y7�}�u�XҊ���v{�d��E��h��1����LVD9 |�%䡿��-��v^;�4�H��A�B��q��h���0x�UE�T�|tmF/�X5�F�!d��C	�3j��{MI��hC�h�����-�	~��Uu����+�_��{�j7�_�)�(!�ʛ��1S�v�����|�WJ9�|Y���/T>o�V8�N~�*r����,�}T*�
8 1zL�¥�&U�)�{�Ci9��te�R�jn5o!W�4�pY�<7�.S�8���aA��y��mwl�o��=��+�.�N|��8T�E��slJ��r��K�j@,�QL኿Y8l�Ʈ�&�_9�Ӯ�z��ًQkݲ#C��7+��
��{b���!�����̗DJǍ�[I���}M�]�f�k�>L��7�����;����?���W�W�^��m��{xћ��"����������ǈ۩]�*�&iРHf6�XuyN��0���(+��v9�0���B|:X���RZ%^k�:�
�#��[�3��`p�Lhl���͛����'l �`���u��n�/FWk��-!�<�c,���݁@t���ۅ}q)p������՜[�)):G������|#7��F`�G1n��ݺ�9y|�SV]-�b�ñˬ"���E�K�vn�cB�.f�'mu��3�6���5�Nu��^��k��9�p���N��W�ɜ�r�=ct�|��w1�i�����r��.�#Y�[3���pw%���\/s���务6��s08����zۤ<��hgf���ȑc��}}�e3'ne��u%OF,������ɬ�݅��Ն��jn��oF�ቶr��\�S]�v2���m�wp,��2e*���!ʗ�E��rT�A�ŝ�C[�r�w$6��[GD��=���̀aAWwv���)�����^��EC�a=Fp���&��CXzo�#���Q��"D��\*��}M�2���=w���R��r�Y�W�����/�E[�v��F�IS���O�9�6�ޏ{�X��ͣ]��f�kyZ�i��\���81�Y���m�)�:�BhV�Z)\�f@� �VV�(畓��������g!-<s���e���ʁᶹl���ڵ�V8,�ER�v�Eb�WaLw��,���f���m7.V=����r�$=��L�j��/l�����8J���vy�����ś��7�;�]c�6��+����qȲ�3��oj�OS\��u��$5�K-.ڏ9��F�>'��n�8YF3�fT�f�W8��oV�8yh�w�Fq�s��+���:��5N��bONd���x���_	[-u�<7�7�EyN5���5�]cwW�u@�y�����V�R�r�g"qԂ������CK�:c`�=���e���Ict���:][�L٩p)�4��3�2�}z��`ek��ɋ�78�9�;٦苠63:j�;Y7�}ϥ{"��
̾�هC��G"A�n{i��0�p7L��؄�VM��@�]��Y�G �N��r�kb{u��.9i� �S+�{q��}l!v�"5�_$�=�W��닲sg�az�f[T�Y7L��jܜ���f�j��x�-�F�����܋L�&[{+|��G����ɥ2bH��*��2�,��j�(��2��r�0�"�L�ɢ��("
���1r"R��Z��
2ʄ�ª�0���0�,̌����2Ƞ�Ȉ��j���"�L�L��̰*��ʃ3*h����Bj����2"*����
��#"$�3,�"��ɳ �����
31���1��G0,�p̨"&i�`�2���
*��"��������,�*���JF��(�����"�e��ɢ �c"�,JJ*)��(*�J(�������&�2�&"�2&�����*(�H�����
�(�
��bbs0�*�Z���*"(���3�j"�f"������������J31���*�"���12�0�J���ʨ���"���,���2J���(��?���s�c=�'�������E���S�D���6A��7&����Ȩ� ��o�Lf>Z�u�Ge_;�������+�_�-��'���$�D>v:+�l<^k��#�5�U���T/V}%L]`�uz2��z��Z'�U��4Y�x�~�;B�WZ��9W<wK �6mw�浻ۉ1{lz�K�	GO{�F��T�\ǫ� ʛd�r��w��^}wG��<��`��5]�q*�,��ν�U���q���>���K��]���E��u*Zkv��޶�Y���vN�c}����gt�V�d���K�Jd���v�N��!\j�c�LG���{PV%������y�^{lc^����t4������6���'jv}j�Tv��JNaT�:�-��`)�z��2%�Я�m���ԫ^��5�֭w���kz�K[G<e��f����p�o��V���,J�B�vז�V��3�h�P�U@u�qgն:#�2�����H�1f��L��a���{^��b�X���`��\�S���#�u �Y��9m��'�{��62\y����P��bf̥�p��
�g,�3~��z�d�ٸn�+<�Vz�zXL��&��E]!yvnW<�	��R/��!��E��epzՙٗ&Lc�+��f�oRm��KS1��[�	שrŠ̕3�2�ӱj�Aḻۙ{׸�}΃<k^�Gp���o�O]ݘ�� �h7�
߆m�^>�zk� ���wOGhݴ�����M��G;��T�L�f��L�m]-B׍l���wvW��W����]�k���v���<��)U�"���Ǫ�����!ؗh��/wy�*��1��w����	B6�H��w.�`��^,�{�،3��Y���L)��՚O[��O[��=��xm3�f��)4l� ����{s&�:�i��hp��{U��z�l�>�=&��4S^�+!�ָ>��֔I&cH���V;P�=R�֣���{+J�y9�Ee�ܫ�|�LB��-o���Ѯt�J��.��{��6����7����椳�u�<K�\\X%���"�g�(Q�o�*r�	o-$5����dl��E�V
.��)�tl��~�q�k�V�Dȡ�«�1�ڋ_duD3}��p���Y�c�:�������J}K��*�!x���\E��NU.�ϸ��2��%�(���VW>j��>�i��}����e3z^E�ո�|�X԰k�±�2]	�?,3U�f`ܧ�[4�XRӪ�8f.}藲}��c��@�f"�z{LS�!=��0��s�������SYq�ق��-��\�w�#u�NW����t��iF���D��0�c�fD�^HsqI'����}]��)꾸&����+x�|��K~��<Xg��`y1�AA�	�Ep�qpy�̆h�]�:���d�mޱ)��u^��8�ȖM����Ӧ����2�#](�-� ��O>��$�����oor�Q|ғ{�E�.X�����2�Ms-���-,Xq*�iik���ou�wLh�M�6�Fy��i��F��f'.��҃�$w;�g��j�C:��e���kWj�<�o����>��"t��=P���-eif];�`U]s)	�}�X�)3�(o�HO�%��#�|5��xR��(�}��%cΌS>�h�eͨp'/�	c�U�Bg�D^M��̅Q�$��-�<CG�v��$W�v�/�x�L/�31n^��6�P�E?a���A�²�`���47�,�Ŕ2�;�}T;�j�[���z�	Q��_'~�oK��|"0xk/���l�Xt�Gi���3�9龾�WX�׻!V�O��
�5&2k��>��4\����y���Grc�j%Ia��X�%uxA)�Yߥ9*#w�V}�O�V�˦7�6��EY[��LLW�j�K�`�#�5W��RV�^c;��.�pٱsQ�4Y�2�)���:����|�Ô�3���9U�DS�6��PӜ�7k����ِ��Z�3� ��������d�4�ﾛ-40G,k��wW����� ����9I�j��!�˻H�%�G�y+2���7��i��9�FEq�+�rCP�{��*�5��%5u�_��D�#cG@H���j�.>wYr��V_mClwL	+T �sSL�(z>^>�7�7�c�J�g�d���e�8�/)�D�5�"����jSP�|Xx`:����,N��[�}ۛ8� ��±��+Ժ#�l�wDa��&ʣʥ��m]���U��d���9[�	�a
�=�@�]pY&�x����z���8v��:|`qp�����m��B8Ƕ�N8�|<=��������Tzj��F��YfW�`Κа��?SD�eܖT��δ�9*���c�(B=���pr��f`�s�����Gp��|ž�T�њ5[��Z���5�暳0Um��$��Cp�`���(���+�.sJ�e�z%_R���A���@�,�xe�G�0�,�İ>2�Z=�b�i�t+��VG7�0Bkv�sѬa}�l�1��2�b��T�E�*�Ͻ�7���'�:��fD�g�]�W�d�r�۞���0KsP<	7a%�;�j�1��=�f�&'D]�,��T`M���Lp��|�:N]`f�ݸ�ֵ��{޺)�k:���J}�; .[=�P�\o��U �����\^\�,�����,�Y)�Xws�Ӧ�ҮH�U�eT��3�jR���(K�6)u.>Kb�ym����o�Q����-ɮ��@%;\r����W��}:���j�����~��\��A>���[J��[�7�Ƒ���\��B�v2��o��}+nqP�:N~���q��Lړ�gW�ɋי���&��hDI(�=�����Ca��]�xK�5�U���x�a2(����Y�z�um�v�-�2xT6&F�JM+��Ԭ�w=1���88Ac{�T�I]�s�En�U�Ӎҵ�$�9g�Cs)%])��+ES4��R�xM��U�#�y�E�1�i+2(^��9%!^�!:Wݹ��l�����r尼΂�u�M1<6VΜx�r�`qx��"�s	V��bCL�}(�[ʱ3�i
���6}�:�r��j����Zx�m�����SΡ��q�9�X^��;DX�Y�'��?Q�#��ck}�G�^GoD�d*�@u�:����Y�Z�� @	D�7��I^��;W;��]W�S,Y��4�]in[��Est�ךX/��]�7��8r�q��a��!�;Z��:�˸aə���RY'nu���ۖ1��%9���߾���⯳��KO�m$ɮ�L�#�}�i�u����d��S��$V=[n�c�����2���)+>3*�V`�gR�����V�t:$�m7G8��-�Dq����bV'���_b��TlU�f�\M�2x�;S�`���%]�ͷ�]p��>9E�eJ�6�ͮU�d�_:⪢��k��(��SH��R���*s}���Yy��/��=>H��R%�n';��T�L�W�9�fU���g ���LJ��ɒ+��Ta�`ʛ����Y���u�m?_���o��	����M��E���S�m�J)0)P�-!�GE�a�[Ɩ�,�M�a���Y˕���c�ޛa<Ds mgL��̉��c#���Q5�JQ+�6�]����z�굧�OGAQ�|p��3�f�d狺��L��v:�;�t�WT�i������ew�vg�߼	��o)q3����h���CGIz�C0Շ6��!A�-\��j{wE�s0Kߖ�BaF��l��Y�oML��!�\��@vA�d6�P{n�)�6�g)�����Q6�������:f�Bq�%��4H�ފ�y��j�a������[��#fS�@���\7f��IfE+���d����սϫ5=�N��3�u�����	k�˕�,P��$3�f�/g���<���pǩ\K��h<���.�f�t�<�w��J��SD솟#��;r��n�GL~�v���+��
�vLDи��w-���/�ݞ�@n���`JǞH��E��z�Le{�/e��§�g��R4h��|����n���ԗ��WvB(���}���s���:2��9X��f�A��Zugt#ɏ�*u��+��ʸ�:������P7�*R�듶��ⴍ~2=x�ɵ�r^�N��sn�V��C�6�;���}�pBZn�׶�y��pg>Ɍ8E��$���5'�oA���n0X`o����W^��&
v��8������Ƭ�G�8���f
s0�å��g�]���=�+�p�MTS�g^�����v����`�+hJ��!�e�pv�e��,˧s�-K���!��TU���~�O�jr���\b[Jm*Ba��f%yъ-�� �����H�;�Sh��Y(�w}��}�G���T3���펱7��%�j�59c�o�ŷz+�:m1 Tu^��+�q�V:����8~���i��Z�:��M�Q!_v<�:Ce�]o�L���KG�|w{�fgv�N�c�!�\E<�������ּZ�M7OP�P��3グ��4A�"uU�RDw��Ϣ��2�E3^����4�R�=��y�s��D���ݭW��E�+��̼we��yi�V�{ܫ���\����S�g�����{��˕���0�P�'��@�ڹ(��X��ӦҼ�႟�t2�5�9A^]k4y����C
�M�1V��X�:�x�p���P��:��l#v������*%e��}���J���T��H�Q�r�޹N
�<1R�[^��8g��$sKJϩH���>V=ܮE�&���lIYp�=Q?<:-k={�QY�>\aۙva��H�)�#��]���;㣕7�ne}�������k ��	�!@<�8i5��Z:o�p�~��3�F,���p�{۞.��Z�v���O�}9֘䴖�()(p/�+Խ�J:��˸gZ6}�	��p��ϵ�RO|�;���y��:�"TS"0y������4���&�xS�����M��
.hS�KF.4�>A����i-��*#V��յ��e�W�e�zD�����wF�# �^�{��4<{��)��L�e��Ȗ��rDV���3��Ү�:P�O��x�'���Tbm�I\�\�ߴӵ*n���8�|cn�I�A�{�W0g�	�i�OS�ך��w�Џ|��>鰠��jY��U\���4�V�Dtzm.��l��������'�Gyvk�5��=���j��w���W����YA���n�9�lPV�3�;��|��~����$�Z���޷G�f��x��2�1x!>�=w��F�]Ckm>3�w��iWn91r�5q̊M�s�ŧO���{�a�����6m+M-4֊��2��T$�"-+r_�yz�d��s|��`����v�5�M�@�'�H�+��Eqt����
�7Y��V�m�t�^���M�c��g"��ҷS���G�:�����+Ի�>��}����,��=���⥬����՞�oN�1W����G\�q��u{�<u �0k䦧�(t��_Zg������u�CH�R>KB��"8q������肷�Vq�����C�"M���A�c}�����j��0k�ү5}<���^�b�۾���KL���/-�D�0o�a�ht�ҿ��J�!�͊��}e��"m/z_��m�9q����Ms<�ŧ��6�[J��K���\ӛ���x��2*�}�ɩ7��{�zҫ�_����ov���wڳ�[�D9�<��]Fnq��],����z��d� ����]�Fd�)Խ�D����΋�4V_���x1����=j|����Ɯ���$�9g�Cs)%])�+������(�WN��[>�)޶׼�ӎYkt����Wl#�씼�<�z�L�3Ԩ�+��������t�wNlc�|/+=�yq���"�k�J��h�
d������X�Yٶ�u�
���h#EW�"��i3���[E=��S��Q�t��plyǈ�X^���E�ЗE��h%�W{�u�:v���V��_f&	�����
I��\�rԫ^�xϸ���^���u3�K��Ho{�n#X�~�1�τT��K��}w��X�P�ݙ�\D\���{�*�a}b�����g ��eǻIS�L\�3�X3�6*«6Z蕏C,�9��zY���b�D�O*�O��!�>-�I�[L�����K����j��cz�ו��SH��|�G\��+�r�ROj�e4����$p=5"Y�ۄZs�O�M�v3[�Z��VZ�-V/l���fA.�|*�w{����"Rh���w�i���g�v#,OX��=�*�y�3�����5d���GjBI��Htڗ���k�]\ݵ7����E�;���{�OM�>�p��ά=�$����OPY�����l�9��r|�d
�x`�­Օ��k�v����a^�%�h��S��X�f�{��x�Q�\���sƊ���R�V���5
#-���m�5; �6kj�a������8G]�/�-�''oS���ƑžܗF�;'{e(����;�(��0�s�3y��٦�s����I\�m]�0,�qx���ڱ��x֧�.�Yo��n�����ו���&
�p��H.e�\�Y5���#�<l�#�u6r�q@�hӕV�?��ogεJ~F��W�}���\j��3����Z�[,�i��	����\���X�(�����u�{O��O���'SVa���K+��؋�=+=3�9��d�X:�a��w9�E�c����<o6�����w{�uqOv*�x%�^yR��k�T��9�~G��6@Um}��7ɓ����}Oyw1֥l�h�˨sXW.����w]$�fU���E&��T�'���Z���"@�3�-h��w�9�N`e'���yV{Dڈ^������[���xo���8�҆6��ya����əg^�p6�����2w^vv�d�Q�:���^l�X���؞����zb�4���r;����x�X��Ӣg����n>�:j���/�r̼ܟ���mZ3�7Q�G]���T��p�gnGϩٗ�,ҵv�Kt�:1f�����R�J��$����βR����J.k�j�R�WJ�Z�t>�wLі�GC��R;��!��9f���E�1��+{�E��E,���ǡ�n�ob���ral볺tc�8bzu�[���;h�qwt�+/������.q�E��c8��:�\Z�^��.��듎��Y"�Y+���Q�km*�C��Z���}+)&*�vf1[�!(P��H]������¸a����m�657�hݛ>ѵxF�)\�PS7�<(��>}����*���|�Ce7rF�%�>y�_�C�V�۶�B��A7��X�*k2�n2n%���5$�݇`���;�L��m�탏J�]%�`�YF�d�����5a�'"�˫	��scg ���C���k�U�ݘ���or�onKw�y75.�Y|_�z�#��q��m̖�tw�8�/	��e`��y���k��G�w׎^�[�%ȉ�\�P.�����W0NOZ�����ʻ����A��ڜ����g@�;3�WY`�M�m���c�'��:,ޏ�l���@�WA}�,IC/��wd��ՈM�_���>��p�-5��5�A�q,Wfi����6�3d`�K���~�ѠG�Qk'3s��0I�����ާ�8��䆸�'ּ�k������k���-�<�d�k��Ko���uxլ�e:�v��ߛ�Ɏ>�ۉů�6O P$"?)ʨ"�*�(�+2�ʦ"H��"��(�2�f��(��J
����(�,j�jJ�#�*c#&J������ �,(�"e��Ls��0������"�����
����2�����&�&���)�b0�j)"j�(�(����"�h(����j%���2���0��2��	���)�)���&� �(�̂� �����%��
���,�
��"�J,�����"���b(�(�����bI�0ʨ���$+(�( �3
',���*(��ș�(���rp���H �����rr(���)����������$���h�,��O(��p7��;{��v_5;�T���8CώEɳ����Μ�:��C&�..	$kH4���}���.�Y�#�>yy��"�V�Gt-���]i�T���4�W�3gZ0�ޱeLޙA幒;�)8,���J��1��C�(����h!ŞH?u�z�^k���	M�
W�~���U���p�GP��v:և�L�wH��(�LƷ�	�{ʃ�^�f"�������[z��� /���//�>�Y��%LB��-h�����t�J�:���)��.�_-��|�p�,'����LƲ^\/�]���P�����	a夆��ŵ~�]/Um�!����)��a�́�.�r�E�?��Z2+0����rCO��Byl/ۣ�ks|y���#DY��M�+����U"<���\E��	O<�Q����t�3����G['�]̌e�4?��k��E��v��$�W���!d�� ��M𘦭Oa��ࠦ��/:�G���ڇE*u�����..�����!�^v'�]�vr��n�i�9\F�(c��I���r^-:l}��}����z���^1	�h�y����_[�f�K�8�`�nz�Y����<bx�+Y���/�U���ˁ;J�}c[�ƱO^.-�zP�Yk���)U�O�K�i��f�ӬCpu}���{�K��|N-������x����]���p�+�͌b^��:3���eӽ�ӿ�Pޣ^�1�[Xd�K�=�{�^}�w�H��`����J��K��Ŷ��}��p�J<)��l�4/{S�0/m���9�,=Bk��S=L�!����w��3}��H��Ղ�����!�e�s��L��V�eӹ�:�<JQٜ-���X�E�
����q�ih�p.�XϧȪ�N�R����D0ʞ� y{n�ei�!�l��D_�3�q��Ojn�c~��|}g�ʠX��]�r�SϞgp5|X��R菺�Mx5��cJk�O�R�y��O�5��G	f�ۻZ�.�X����PL˞�2�Ӝ��{���N��7�d��T0pȟj�c��e�K�h<�{l�Kw4xc�}�=�;�牲�
�,erR�~�F��xwîgcVtܗznd��P!�;IT��Xa��J[�1��Қ�|(S=}�C�M��#�5�Vf�������j=lf^�?��r�l�V>%y�y�p2��HCe.*�'^��_��ȶ$ձ���+"d�/!����+~O{i�[�2�e��2/u.�PL�w-ڶ�H[ͦs��Ɗ��h,a�}�W�P�t�ɠQմ��k�	�M�R@̹s9m,�v⣳]Z�c��(sJg-��n��˨=�׸鵢n*+,� ��!�z�U��.�gh#Ӭ;/9��
$��5$=���ܣC������¶8g��x�:�0�׻f,��t�g-
���u�ҼSҸ���D���Y:lL��>~��9,��͜����_6�������~[v���3��P�JIv�,)(0tIX֢��9��2�e���ikӿd�j��١���Z�ׁ��Y�x{�l!Q�_���y�$��-�^�:�X;:�l��oh�����c�j��)y�ʖ8�*��![�%,x����At�#�yX�]Io
e
��3�:���f�۔t��5g��W�,j��;��ؠ�W;��I��W�L)[��;4����R�bMBL^'�g���<N��aA��ޤ�WB�-����o�F��ީ��*nf��oW���w��Xd[�0�7	G����KG��fJ:x���}-f���E�&蝅`�J(g!;��]��k������O��z���5����ۀ绳�>筍����1uڞ�&W(�U.�Q�l����N��{,Fw�(Uj���� �ؘ��a��w���F���MB�{;fqB~�P��W-��$p!ݡZ�3{���(H��1aD��ٗ���{.YQ���jv�wz$N�T���gV�rz���'�g9��X��B��o�d�r�5NV�5���`�\)`�����g)˚�%y�U���B�o8�u;�,;�*�r���������>���{��h�@�a|�E2�y]I���Qz��r�q$摵59s�=r�7���h�����F�w�0L�a����Α'�/��⿷�l<�v��.`�B��xs��1���Qڴ:r�z�R��|'�9��o醑�:Ri]S#�X!���qv�J}����z��F��(5�:Z���ϥ����ӒR���',�*�I*��"��
��X�,'���;�+���}����r�Xs�ZH8�|"�`䔈�o�)yX.��޴�6�z��~X"|�����t�vR�����ו��3�L������s	V1�o�2M��O�j$߮Z�G�t86��m��.���o����f��
Ҟ��g��v'Ϸ�b�8��u,>��!�ضn䃘�7i=DW�ۯ�,�^�~��k>��+�S9�U�i�	�?y�/�����/a�l�n�X���v�*<x�1/)«�bL�[����̀�h(�=���^��nn�^�4wl�;yVp>������}�>��)�k:���Q�:�Dwtճ̳Xq!�h�f�vC�ވ$�����}û�]�P\۝��ג�iqe>�E�4��v;Z�h��v{L�En��;����~y�|���O[�n��,lX*L��P��y�=��֌ߨث
͖�RV=\��GƋ~���k+��ch���j3k�$��f`���ˌ��AпQzm5W�Qυ1Y�^��˧���N魆&K��vq#�MH�ڄpNv	��I���x�5㞹��*S<��\O=�:';n.B ���)Pٗp64Ұ��3gZ2e`���r5����'�k�	����Z�H�GLM0o万a"9��v;��K�����};�w�Z�v���ƫ�z̦ȷ�ќ�`�h��J#eq��qw��A��s�c~�����؃�����TGB�>է!���M�zw���e�����cYA21�x�8�o�����΍�k������S��íz^_�nU�ᒦ!G&T�0 ���:E�������q�{�Z[���O��g	��@F�B�	�%�������҄���P��X�7s��,�+��+��dƟi�MJ�\'8��@���3\;��;"uT�v�)�{�v�y ��.�����:߀�t����S���b�7E���V���b�eG:���X����:T�����o�VVp�-Cw3�[�J>��`�sm���wR�6��.��NO����:>�K��n���ԉ�qY���*�d�.&�3�A1�]�9�+Eͻ��rum���72CK�����
�w҉�~�Coe�j¦�_)�OO7f�:�K�v՚,��q{Fz���֘Z:�$�W���Ei}v(�t��y��B�����+G%b±�2����`ǋ�;uA~��xe���ʚ�~��/L����8+��v߰�	:�5�c���ƔՑj]�6��87��W�����^Ky�W��N�\�������%b��,x�ړ0R߼�2��/�<�ܲ{��l�}�N.#h�v�L��K�AKH�\G�]Ȭw�Y`�>��U��N]��t��]���q���ʝ��Y�\����شZ��j��KmR�+��lˀ�ݦ�k������B�����֬߷���cn�w�^_����C6�mDP�=LP�����:1E�.�л���gC�bhх�8��hN(f�8h��a<E���1%�Ѥ+\��o��Ю{��<�S�T,�T��:�W<�&/y�ϧ��Y����k�/�X�sꢢh��P�j�o����h�`��fZ������w�Ç�^R�9@hp�:p���)�����'f��k_��e4<�A��.���R�[����Ƕ���U#�_�sۖp}2!�����A���9=�ךꟊ�p����k�W��)ׂ��k�Μ�*��+[��S���,����׮)��d3)BH�]�P|2��8�맜��7���h3����B�e4��2<t�gٷ2j5����38߆Kx��X���=ݦ�[V�\���D�jX)s]�)���ġ�)4�X��+3Ox5sK��yCá	j+�+YXE��)Sp�EE��X����.����R'��Mf���h(�<V/9R�wCО�C���HU0��&]�s��H�GY���5.���^�o4���bIƋ[�W�V����\�|tL���X��0�h����]��w{Y��7��{����X%��@O������.X72�=1�{_+հd=�#���<�{e�9�B�X8f��06�oB?t�R�
�7y�����#��k<��pa��V��V���
1�VW��̦2��c�d.f�=WT���=�ŉ}�s�o<�|��63k#t���q���:pn՗�
�E��K�e�E�v�Ϲ��|<�Ѱ�O`���Wi�#�݄gOS��v"yI��
[�������
��8Րҫ��Q�k��@����1�=�^|�\�g���.�m��4kVe*�xyG���Ӟ"�/�	��";�о�J�{ؤS��.�Օ3Q�����]���t��;뵞ڴ�Ǒ�vA^U�Cj!hbb�v�]��K�	u=J������������9��<|bϽ\��/���<��p�t�~�qz%��$�z�:�sۢ(��cu�37\D�f�'"&2�索��!����AcZύ����K�H�+�=[�5i��Py��x�>�hM����$:�]Dvzș�5�W�.�����t���E���>;�c�葤�K��-��qt�&v���,�FM�Xy�ְ�c�<n)�aUD����|��;)b]�~d0q.j`(s���� ����[p�ߥX�3�X��:뗃7���C���[&r96�c�� ��&�:D�q}hPqo��|��^�:Z���%��r�.v���ݚX��j��IsK��[����ɢȷ,�9WL���:ֱ�^.�+ίk��N�]�̹�b��=KɁ�Ev4����$ʌ�ڸ2m�n��9 ��ӫ3�u���8��r�غ
g�9���na$8�p�p1�G��R�]�zg˴|U��I״��V;���E;�{ނ?wUڜS���N$f��y?��ϵ��,����=��`�]b��M!~�~�o�p���_C{qP�{u"B���}g-�w�����c��n�`36bI֤�s��b4b�)�3����JK����is�{G:�%;���6R���n��)v�gէG���-k�J��h�
d�cղ�`��������x��g��+�ұ������B��c�^�9�<U�
<'�[����~+��1�̮�Ѽ�g�a�I�F�յ�1Z�|�10Mfu�Z|+h�Mu�GV��>�i�NJ]
S9�K�z%�%R��'jyg�p0�z���6����ryx�E��l�y�g�o�o��+��m�9v2P��O;��n>�(RH��ġ0����I���o�>X��vMv�=�0��V�3*�f�.3'�A����i��a�E.�A@�N����eh��Yx^��}��)ċ�R%ۄZs�O��6����4�MW6Cav��PW�}�喢�Ї�I��λ��4��f��E��;�2^0׮X�I�ݛ�Y]��Gd�G����7�\C���J���x��^,�q]�=�)ʸ[�ãhр6�9����y�L�}2��r� ��B�3�F��.�w��xj$h+�^M��<F!��eĦ�٫�$��؉��y3C]�$5"�m�B��ڟ*���s\,�r�G�Yq�н������·�:X
"Jᗷ]r]+F�J�E��F�J�\�D�ז�2цI��;lkV��_��}7�7}v��mƶ����>Z�5�ڟU���=��ؽ��Y3bxS;�@�J%�*��gAJ�����*0��(u��Lj��Aͧ���//�nVr�J��*b�z��0�{�;=����==��´m(+i�uP�����Y;��g�����9��S��������_4m���o������M[�l��"������Qy[�H�+/>U�Lܭ��,�opc���8Q��0:�TD6𚩔��9g��mfHk)rz��,Vssh�P�x�������Q�븠��r�j���&{��pu�C\����p�:��%�6�|��=�X�8M�;|�rX԰l�¿9�3:�<GM�mÀ#��>��}�b:��i�gz;Rh[������^��.w��@}qO�[H�� ����/n��^��5�w�����MQ�+��l��F�n1�|3��Ş��K�[��8��Ǿ�m��6��`]�ª�Q���,�d�*�)��|мC~Ǡ����i}=��WUU�f�"%<Ҍ��|��7�"�p}X͐�WUr&0>X�Te�j�cw[�6٦qUL��=��:C�\~|�Kٷם�˺?G�=�r��6�I�x�}9���y����z�N<�\��V3�׹(:�6֣�@�38X�oȺ��s�%R�.����h�z����,3[�³��]���b��:����$��y7��gYA\�T!��C:Vаy�[ػ����r�P��9�r�d�l��E�q_g�Z߼��d�9�\���G/��S5�.jD1b��K�]�;z�>�ٽ�rf�o�zK֜�E3R;��mw 4|�_)�&���Sx��]��t�ƫ!#3��ᥣ�;}�`M]�Z�� ]\C+м
���;���{�~�o�m�J'Y�I��(J�v�[\�	/�:�4iꢈ��V'�e�Y�`E�Ǵ�_Rr�M2P�ɒf�i�Z9�h�k�u wa�j�c�W�"�O/���={���X���\��Ʒ�����,���+�Ѝ�U�
���%�=of[X�\�:�c�/r
wa-�m�ኘ�uson[w�6pǨ��q��W�E|��g1D�X��U&�z8x�-������U<��F����}��%��:�{ۮ
�I�m���Qt+���j�p�ӑRR����+wS�ꔍ��Y�55.4T�^!{u|�r��n���L��k[y]�!�*�4��k��Cڜ �y3c�h��D�ڜK�A�zT�6[��5m�ŝ\�^K��ڡ�.�K�ovG\���̮p|���OrSi��x�-X";]-�vMe�h��X�}�1�+�X��}Kc�Rv�� `<Zt�|d�W@w �@cOX{��<^�[]�� ��F�~�]�k�#Y�����a����+�<�\����e�|qK�z�>�XqάB�/v�*Eɚl�`M�X&.���tw5p�#+���=��Խ��HL0���g5���{|�;�#�Q�f��p�}%�fiY�����/��b�,�������/_�$E3�d�ev��T�9�Z�=���]�����`��|�^ax(2&[���E��V-;�U�34�.�V�O���<�{�wT���h�]}��!�����R��.�|-Ub
��+rT���r#�WJ��:�͖��Brj��a���c�|�T�|:�,���ԕ�B�.�l�/��pi���ݣ(�,�]�g����B��c��9��r��6�EZ�qp}"j���՚j,IonKtv�<w��ܜ�F���>�n��V���gaad���R�5��ң���c]�C�+l!7ʋ����{բ�}�VXm�V*����ry�B&\�chr�P���"�5�w1+..!a=��ROE $���a� ���T¸��^M�ޔU��̡����)�����Z�٩X$W
��aΜ�Q����\��8�	�������h��sb*�0Ɩ�"d��*�j�
��(��0�̒2�#((��r���������̈���"��"��0��*��L̨�2�rɪBj��*�&��*b��*�**&�H���(�����b32����� �*=���-A��ȍYUUVfELF��effTa5�0&���+Y�fa�33�h5��)�S������f�m`f�+Xc5��+3(����"���̉�M`d�ETT�QT�Q&a�k0b21�(*�Ƞ��j�� ��"�2ƙ��X�E5F��+,(����� �aQDS�L��i�58D�AU:3Y��ʪ&b����+0&��"�&�NM4D�IE4LY��QE:�(f�j4�DV���+Xc�	%���
h�#"��*MfQYe�sS�����+���B��IΊ]�8��9�nvS����@����Y���9���hM��˴e65�vuBI�%�:Wݵ�u��u�5ܨ�p(z�I瓫%g�wz�h��*�GԆ��r��0Bl˔��ǯÄg_xbIgwW<�� c88�=���t��Ţ4]��/a�b�Q���M7���:KՀ��K����2�� ���L|iUF.�ezN%(�q!���2�Z=��'�̼ǘ��)�Stow��#}T��>�j�J+�}��<�N4�Co��֣�:����wm%Oo�oӛn�:Ԡ���λ3��c�[�[,���U��P���ЁQ���`Ej1����_U�oƐ3��`�R��)�e4���dik*��\�8�a��fq�;�y)y�Ӄ�M�+��U֧��_J��#�vЦ{�Q(x	��C#�O�{	w;��e˱�Z��&f�w���0Ư��P�fY,�$��K��N.���M����,��b�{��\�����˥������i�9�ʐ^B�]�^��#�]&v]V�v��q��y�,T����o=#)#çLw[�D��J�+f0rJMp�哦��w|�K��P�4

�!>L=�p+��d���Y�+^x��y�Y��z��EJ�J��
~����̷=f�l��u����^7䲄��}|v.���̥�*���R۷�Wz:�"ޚ��
��n��v��*�ޕŷ"*���u)F�c�`���Փ��	��z,g�������X`��V5���,x�2������欥B���i*W �O��*0��LL���Ə�2��0�c��$X�L��]��G}�GU��Ҳ��+z����ח4�j�,q�Mx�mH��o^</��`N+>,k��^��x���;��FN[M�;%�QC�������1x��ȯ����ؠ6b��N��d<�mw�r��{Jw�S�
W/F��2���Um��P�V2
�U������c�o��:F�k��,w���3!���{Ǉ�m�\*�&��qz%��	��M�<�۸1o��m���=.Y5��\I��&2�索��&|\������
h=@�L�2��s�?O-�����Ľ�5G�Zz�Q�܉�hO,�dNQ��O���ŶK����7,R�v���s=�0�QĢ\	;E1ݗ�x�u-d���]�=�B�D!Q�a�9h�'�ˍ﫲�����v�x� �50P�����.�O.X�3��-#�3�lr�㳩��/��Օ����ïB���:x=�ٶ�3�p�0i��y��9�5n.d
CkR����+�7w��ȪD��7�
_ۼ�l�=B-�r�$� �79�v�4�=]���!���r&fuJ�qs��F�X4Rɗ�|��X�Y��u���Ռ��#t�s� i���$��~��Y�v�� �� xS��W�L�)q�ٸ:�̧����8�Y���ү5�^�T�������0�NY�r�;:����ai�Ԧ�#�z	�f��Ϭ���\Y�KɁ�+��>���%��&
�ZIZ��a��C�r1�o|�Z�ڕ�ȫ��;k�Ot���I.���p�0tIH�D�c�Xo�[�էWHE�նIc�=2尽v�/+=�g��i��-�Y+Bf4N�(�Y������\����h�$͔mo�sk�-W��hx���L�>S���d>�^$��4S<G ������"͗�;Dz�B}�>�-ƿ�:׏�O�o�2k���nXs���z��s:�卋Pe��{���U��L�A���K��x"@�o'}�Ј1�+���ݩۮ���
�>�p�����\L]p{��<a��XUVl��?=��=Щ���w�����uAN�X��N#�o�$�m30S���*y3��L���f���gU�j+�b�-�F-��+�g�W������fk,�g#������Q������q�_��F��g_iN�Ws���b�i���_"�>��O��h��Em��V�������ǭ�;�����%eqqDM���fjj��a�/:�'<�B!�b��j��Z`��4�G zjD��.u�ʏ��k�iC�7.���YeNe���C�+-r�Ї�I���.�<li�=5�֌y�y9�s5�w� ���1������l����<mi����#��˱�N�Y��ͼG�*S���>��ޞ�DQ>�����ծ��=��1��t��"�|C��,��f��ӟe���/ݝ?���-�[
f?a��emyN(���z���Zߟ�3n��(�-��Ol�{���>o�z����}���Aͦ�C�]a��Y��d��QϦTłxPu� �����]J���e�v�4';#��R��˸z�m�]�޲v,��cR��o�s85.�C�����#�����+W~�e,"PC��Hf�\��u�^}w_��~�|��cw��VY�P޶��u�+{�ٙ#�W��en��ܪ"	�8.��I��Ϯ�C�:�.�#3��6�\D躼{3�^�A(2f�5e�bCOR�����f�A�ў��t�ah���]���o�3γ����{��k�<������n�i������.��y�
�51%��pWl������q]&�8{��J��C=�V�vT�s+�c�+}W\�s#c��[����Q���"*�w�BT���ji��cs��D�+��x�z������'t��g�య�dK<,�{�L~APs���եݗ�"�c,Q����t�/H��qޔɗ�-�P֑�k�ǳ�cK&ע���N���}���
���kG�ǮQ{H\��
�nA�|3�߱g��*�x�ߤ�#�<�2�Ms,y�,H>>X��!9�촬زV0R�e7���Lu	�=�g�Eސ^�A!��z��N]*%%���*�5۫w���i��/���$v��t9 ��e�s��-1�ق��!�.׋�T�ќ��yy王���X��v2�ǣ�(�����3�T���R�f�)�^baݩ5�����cC����	��!ΨK���҆l���VW�� �L�Ȅ���s�Mt�TF��X9��R�y��L5�8�d\�CmݭT�2���;ֽO�󃼏PƲ��X��wu�k�]k:z����������(A�sik*� ����~&�+'fP������3,�������z��\�8�k=��
�K��s�imX�gr�c�[��]
I��sCKgft�6=��=V⦒��������AųM5:��v�+�k[y�d��	��/�K�VsC��G�g9�����8�q�v�ǜ���M�r5��&���t��=[����o�6M�6/��n����`�A� ���J�s\�g��ġɲ�C#�5�گf?��v6nxh'hA���vu��9������|����e�ȢH�5��Rqu�es9I����MG�un��w�vL�ؚ�x����?}���!�<1C�˳|�i��Y�&v]s�>�C,c�Tc��[��ʽ�x��L	+T!\���JMpr��U�� ��֧�K50�w�ڀ�%��g=�xg.=j�I.��`Ia�!�(�F��-�~���W��js����þ��ӣ�R�Rc�r߬�ͽ��<'�`˲ +�!IjX�f{�c��T�l�wQז\*��߮e1���
̇��4JU��N�M����m]�E�ҍ�p�$�pM����hٷ����I_��/:�p���7�Qj�;X��Y���/#�� ��/�m̚P_��v�삽r�h�D-�1x;n�������n�O+d	[���ƏeOR��_8��̇�uKz���ێ�U�L?[������V�����`˩GH�T�f���1N�fv�^�T�]/�`���9�r����F�G��a�v�.nԛ�us9�b�i[yM�\e�=�%���7�/x+���>�2��q�9&�Fcz^��nD�"V���Ps�kp������}��lv�op�?�Z=*�0�� ���l�iE� r��`�,kB�a��yT��l5��kro: �D��[X�왃��$$FM.zș�5�P�9�&������i\f�ҮKE���C�
��I4�6��\]'I�)˞0��Z��&:�r�@���T-T��}��j�2G�7�(;R�;�v�x�	/�_]]>��xxmvvOZ�&E#lc���c��L+Y{������>%�+�L�OY0��D���"M������;�΁�n�R�W,}=0٭������������%L]~{!ÂxT7��H��I�{����9�s��wj���#�B���q�����=�v9���$�kFIbr�=��&��u�fA�:ߛŉ(�"��}N����h�E=��Xs�ZJˊ�]�dH�*}&R�w@
�S�B�wi��- z�Q��K�E��u�8���tz��Au���5@��ͻ��~Rs�������@[�zUm�f�m,�����W�爱�{lc^���nU���K^�L�r�Z�[+
�W-`�B���o��-�h�YY2��$L6�Oi�JŽ�xl����쩦��k���^'>Z����^ѭ�N�����3Ĕ�<���f��mK����:���RC��:�����8]Ŏ�#����/���@��v����:ȯ,YPkAg�*�^:O�Y�מlr��{i��R�@ܾl���0L���퍋 ��oe��n�=�*<o��o�z�����`���¶��y����s|�h�g;�i�0z���0V�貜��uJy�;��s���!���;G�[@et��<}WW�ŕեd�zʑ�I�[ĻV;��0��Wɲ�}�7�=�z`b�sc6��ϫ-yYED��?
��b`���G9F�ni��5"�6x�^�귚�r���B}�_�ٷڽ��`Zh3du't�l˸iXzj��Ճ/��i�z���hԎ�<p:��^�NX&R=b]��֚��K�v#���]�@F�5\�e�j����0:�W�t"�˙���������;4Mr-if����d��2�Y}�],��DJ�ܑx:�i�:����Pd�FV	�;|�i�wHoC�Q�^�OE_���٬y,JUqm Y��<��O�]íxK�Ӆ�Y��*bO�x��O'��w�U�U�Ł
eB.q������qn���uɖ���fr/�B)��<�Ш��~뛖�/2�f���{W����S��y�/�h��Q�F���W�yC9�W�ۍ���OK*v�'�bFw)B�ri���\�x�3Jɗ�+�=���K.��>�J�=�BBC%}}pvnd}�	w�z�ؙf4����Wl�պk7��~|��;o�����V��E�A�I!��rV)�x�=����^V���Z�!�v�A�X�q�0f�#��;r��l<&���H�[{�!�\��r/9���;�8��:�s��n�S�L�Q��D���#�VhpzD5αZ�Mp�.Y]:}k��ls�9��Ov{��]�gt��`��ỳ�i�(�_�p�-[̫ۂ�ͯz���w�<����\V3Vg	�c�(*�lV{�e%�8���P�W�iӢo��yҒ�g���.^{dG���Ϗ��k��O�>�p>!Z���A��I�� �K�rq�'S};��V2Ǿ>���n0i���tp�r�/A���Н�g	r��'Aq�����#�g=�c�&�5��n�z����Ŕ��-^!m�p���^��2�����}p12�F`U�άJ�k���GE���8���U�������x�1�&og<w���}�H^�$�
tu'Ǽh�����S;���^� "��J��ّQ8��u����[Xv�y��:�W]�w���Ϯ�#nG~�c�Q*6y�{��u�ə�&i�̔���Ľ�x�Jߤ&O~qXW1k^�_f�z3��u��5)~�y��P�as�D�����Ҩ���ԓ���ZG��k{�w;��ͫŕz��gyAU^/.��u��A��yt�QXϲb����E�f��Բ�`�z�Ϋ˸���a��>8}txK��n�<C]z�چ37�L��z�~��*��ΗJ�D���HvP��f�:��e����Җ�l�9�^��sX57O��]i�Td�9���Ӑ~>0dy�n�;\�:��Q+��r	�߻���i��'�v��[voo��4���Vf�
���E|�}r�ܙd�f�#Z\R..����O�������^4��v*m>K��v�Jȃ��ꐪ:'�Cؙva��H�GZW��_��g���J���M9�՗l�O���֢��W%Bɘ��)5� �����K7*L�V��k����Q�[���Qü@��`ܧ�V��C��줔��rX`ؒ��Je�tg�r�ܑ4�xx<N��~�v�!~�,�z�&w6����^����Ԅ.��`>�wv��?.Z�`��݆�^��g���d�:�ȏ;�N[��Ksn���8W�g�:��b�Q�Y��O^����_[tvE���s;)�E����{Vq�T��J��}�l�`��Ea��;)`uq�)��Mh+��q�����:0�5)[�]r�|�{54Ƌ���U��g�\Z���F��#��ۯ<���m��9���ˏ0�:N^��ɎK�@�
�x{�M���,�Rঌ�7�-#[ɉڛ�hV�PM)�R��Q�t5��̌s��B>�P:&9s��Ù �:{��}Z���`Q#O]�ɲ�~�͇H�@�
�|�>�Y�,�5�O�˛ �}+i^���j�@�ɴVl��ɇ�������ȯ	}��y���vp�K�Tg��kz�$�o�םHm%ڳ��7ͫ�!��,����`����'����^~ӹ���.�"��>��ݻ`ݾ(C}���;q��Օ++dszVu3�g��x����x%I�Ԯh��
6l�W�9��ڰo)�I}6�HQ�/e:q�b�c����%Qe�W�#D��$Q��G��.�������s����P2n[���s��n��e8�;�ɒ�$����;�-�(�7i�k�#����N&����En��sm�D�������a�Ч��9�%�ʹA�xػ�Lk�I��b���z�^ϡ�gV��Cpݸ�I���)f�s-�ݐ��ls��O�T8'�X����źf��\��;�ϯw�t+=�@�s.�j�*���;��T=O�ʌׂ���P��7A,=h=��z�R�o�)r���c匱����s��2�[KT�R��[�Kj^I �$ڛWv	,�J�]+9�r)��28znc��S��Գ	m:I�}�Z0����uk �[2_�@�Wl>����^^[���R�5�7�*��R�d�b�|���+1=}��br���}/��sQq�l�;��lo������-h�?N�]FKCMcd�'f�J��Jdpݸo�&7{ڽ2�)�H����˒/1h�=��i>D�%x�ӷ��~7�nYYF]�ۘ8�si9�T(RH���"V���,�lR�ʭ�����v�^_<��dޔ�B�3n-�.Zz�rz2�%�j�����.T��3�{$�Z!�εd�eM�]?g�ñ�z�!~�þ�G'd�����Y�ئC:Y��A{�T�Z��j��<ϖ��J��N�l�+��6/�mM`��7㯬�8+��K�:�Vv���<�����^�lZF��z"\+`9�K��v�**=�D���v���d3+NVQ^��t�r�I�x�`�=�iqW'oNqC��YL�ಂ	R��H��
�/q����ʛϭ�o0�i�Ӕ�C��V>�T�՘.��]or\zD_�Z��#����*wŨs�o��s�t>V02��mc|�vz����J8����B��Ļ�3�
{��s�8/U��.�k��a�&{��vn.��vt��HH @$Q4gִM�Z�j��	)�&&&��`�������*��j��1�(�����Ց�5�TfTEQ�2�"����*&%�X4Tј�afX�D�E� �b�M�)�*��J,�"b&�&�b����+Pa)AEPQeE�%��)��*�����"���ՑALN� ��"H&�b)��������5e�e�!3��Q�"$�ɪ&�))�2¦&��0���I�T�DE5DَEF`eQATUDDLT�UAETUD�Tc2k0����c�ڰՑAMDQ5A���j*#X�U0�DRDUTD�$ET�%ET13EATj2�)�(��H������5�SjL�*(�("f �bf�$'���Ix�}���R��g�ݜb�z��\}}�Y�^�U1	|�ͽ{�cj�5�~(.������蛐����n��սo;)�d���	 ���v;�bT3k��"xL	�k=�/H�W�㶤^�f�႖,}�����M�;�⚬���o��=�Ӭ�D0L�������1W
e=fT>��~��7�ְt������N�/��S�
�Ɉ!�C>L^ۿa����s��v��bi����7�ᤠ|(P�46z�Qc��WNfCﺥ�P��U��Ax)=�y�W�c�}tL��l�թ�Tʹ���Q=�jlgQ-���(���Wyl�,kV]�%8+�����O�\��z
�Z����euYx)WR���ȑ�8ОY6���;���(���i�RR�yav��<k�pA���,����\���m*��:L�sW�m�<8zҧ�k=J�_�p��d��X}�<񸃥-#��@��0q.je
�/�3���0�tީ�JG�e����;4J��I�3}�\�O[92��f'�D�q|�W�Oa��V�:3����/5ڧ��0k�ү5�^���.�	�O
��GY+���W,}1�$A�u���]��<�LV����k��Q�;[79�bGeӼ�0����~&�=^���K�}�h�'$�_hA�Y���k�{0H�wq��Y����{�����Μ�X�<ϟu�w+��2[�S���ˬ�v��{��d���W"�xef��c�-[\Y�^L�]�2%K�dʌ�kM��/]�o����Vh��K�CҪ�W�|,{
�'0q�ܲMt,�]�d���4���;�b��~_�����|�e؝�����������v�8Rη�d���p+��}�o� �A�\p(��@����NX��EQhB��Ƈ�}��L���QO+xdާ�˥+��}9u5��*+e@Q�:�qaz�Gh�W�C�r�_U{V`L�6G�>G-��oA�9N��/P�f`�����Lz��ş�>6�[K&�ݵ7�Z@1�m@�e��}�]4>踵�UBҿ��6�ِ^�[c��Nfx:��<������X�v�ޞtL�Jt W�D�Xg���r��z.Dp=�0��V�39x�j\�����:_�~��g�X�F5���s�L���/Z�W�e0hvq#���PV_�����u�9!��79����FkyKP�
�\����6GRw�*2�P�����P��V��:�@���c�����}Z�,ͱ����N��x���x�h7{F'K�r%iB��sl��ڻʯE%��5К�*�ĥ�x-Хrl��9����*�Y�wn�W|B���v�����a���2�[X�@�9�-��p�nu��L���.OX�:��O����)�.��kM@m.!���yb���h匯V��ʗ���ʔ�d�'~� �U�O�Y땽���-6%�'�Q
�ڳ�(���=����2� �:�~�x�]��s�+k�qD#�������A����i[8.�W�/�8�;� ��e�uP�HG���a�΃�O�.k�^bC�^��e�5b�WV���ʼ�=�Cne�k�"Ұ)�.�]��;l�����cLƥ]B�+z���7&J�n,xo��\rdIb�wI!��Kir��)�uz�Mp��:&��/=*N���ӭ�x��Kev��ܪ"d�<
�+�-�r!Lz���1�����M��K)op�{:蟤�7��EG>���4�,�;aY��h?��JΎ�s�V<#[)[h�7WZ㙛x�n��;��K ��~s 8f&uGh���ۇ(��#t<�z*����r�n}+�P�ʆ�ۙ쭵q�z��sY6�%������� _�K˜cR����|���ؗJ��Y�~M]޻�����^�:�-j�ΩY7/�M
��7$�Զ�kc��+7�օjR^��}��=ۻ�v҃�V��H�Is}ʜ��wk�zƧ�<��=��E��p�e�N��5L]�=x�T7݁'8�GVZ�kG��>0{~��A�qŞ��d���k+|�k� ;�����$m��+�d�]jөTH�g�#y����<�Bq]���h��̳�:�.*g �2UǺ}��5=�;i��p���Z>6��şR�@�9z����M�g*��b���d^u	�؇~���2��#0.�����^[���x��P���mM7���Fh�`���|���q�X�Y7��s��Ծhx}8������VWb���$��1�δԃY�8s2��ڬ����+>,�SW��J+ϲb�V��xFv�_�N����q�<%@��W���2,��fX�v^;���WZΞ�C����-���C��X��.lߞ��=j�$J�h�(���yB��2�R�~�F�u�îp�f>�1ǚĸ^Mt��5sXxۗzo�[ņ���TK)s]�P�{�Q(R˞�u��0�'�9I��hy�Y�{�T��H�Q�P�	�K6�B�qW�=㮼�o��D�fRf9�;ռ86���Rk.��t
>��xmj|8��2������lz�	�.Y�Ϋ�-�����h��w�--�|�w��I��ܩ�4wQ��^"��^8�¶��,Ie��x��6���"F]p�V�G��\j{<49�>�'wb����g/l��`�`F䬈?Ev�{�Y�C�˳����9�Y�����t�--�g׵���V��Qgt���2f0rJMp������w�>�u+/��;���<���X����A�%����ڇ>���a\�<_���U���in�+��a9�Y�F�'Z6}�	���q1�|�Y�z�4X�c�3��!s�{Y��B7@2���]l��/vH3k��"xL	�s�R���c�d<mlk6^(K��>`��gD�~3>R+>8<��pM���ӻ�б��>J�d^u�'����ǺV�a���"=~>�lL`��bu-a������d�C~�Z�&/L���8�'^͏��czwV��R�g
�	ASVxõ��C�_M������b�;.��\VV�j��9`g��g��7�%�o�,��5	7�D�V=���!0�oWm�%���^%����(xe�~5��a���jc�"�t���No�#�N4'�M�a=�t���Nz��Q���q�P�8���ϊ|���ǂݏI�1-���cM=����ǣ�Y]��2��{�I�(�>��zl�+�����侂�,]�3j��x������`�؜zv�r˼kU�[���{��ˉ���η�^nz�W�.��}oNGB5��]��C�Qi.I�a-�gԫ���3�ܹ�����b]C�=m]��X��6Z/=Z������\�Gmݠ~�8�52�~��N�v�W��|�ݐ�j� ۗښ�C�ī�+*G�h�.iΪ�8n�UMie��r�c��r}��
+{���y��%KlJ���T/V}%M/E�h�Fy�=��β��3"爤c�M+P�J�3��_����z,����x��R��z�l;�h#3 ��F�|
��-�c*m�m�#�ۖ�Y<4{
�/��to��$��`�%h��'�Ԕs2�I,��3�o�t,���J�d�C����E�U�)�.�:e��Y�xL���f�+QX��QqmbCL�t�}o*���� �p��){~Y���*/i�k9�ž�}�;����>+qO	P�W��(��Ȱ�&W��Jݺ�-��J��*�wD��IiYP����fY^�,V�ɮ��h�w�6,@|o��[K>v��߅CǍ��~�{g'@�����V�ϟ/}��,RC�V4]���-S�z�W� ��������;��(��w'V�mK�7�#�\ey�K�y:��Tmn��[0)�]me��tk����b�;��6�������)�9}Ktɪ�sy����[6\;i�gu�wK��F��AC���u�Md��X�Jⅿvd�q/Pؠ�3�BҰ'��ܻy���D:���s��_�t(R�9onКL:V�vMv�{|a'm3�a��5%T�)|-*Uz�O�O�-�����_^�G�(�#l�/������z��+̮s_{��V߫pʏ��;Ĵ��0w�U&�;�f���p���Z�U��
�y�*�ѿP��h�kv�����7}t�P������4Î�����S�L�zĻG��5��s[�1f��;lⓞ�d[U�C�u�4�x��y}�O��?�ߚ�U�_�d3�Y�B�Tz+�zQ���Z�Ae�B�r��\�g#Į-��]eD�V�Y*�.�Z�m���Fw��N��H%&��T�k(&E^��:m5*4ļ���+9],LiG�y�I��s/}#��Q�NԞ#�@�:E�t�x.����.��N��1��xj!��U���`:��PS��Cr\.�Nh�Y���r��)�U�5��X��:$v�q�=���tZ�/L����3�\��J͵K�7�f��	B��l�[��%*�#�:X��w���Ե]vH2�y��\�||/�mv�W0g���V=�d�d5]�f��Y�j�pt��2Só�Q�n�G��������%��������-�Dt�V^EV�8$4��;r��]��T��9Vy�g�'�f_`��c������M�g�hn���W�*9��!��dv��(���v����r�>R��ߎZ�~��V�-�$���]�`�ƥ�
���13� ��m��5�e�*fy�F��8Fr�����^;Ko�j���c�(*�lV{�`�y�iV ��R��V���
����P[v�(Ӧ�6��[H>}���)׌�q�p�|D�o�E�v=�m������w���J6���!C&���ź���7��f�\�SB�ug�a�B<�! w�'�7ևO�MЧ]rA�wU�T:��Z>6��ł���P�/��nua��P�Y�ޟh"d.��`�PbK���]ht��<�q�ڽ���pC{h�R7�	kU�c�s���R��]p��u3�:1E�M�auBԭ� nL�x����K�͵������!�x�>$�'eئ]�+Ag"��'R���옼<��vm;���y�=��;)m>߳[<Ѱ�c�9�)��K���и�H펒��o��ʹ�� �s����a��#~ϢyBƯl��^���w,�4浣������h��ls"�fvV>�԰�*h��W&W+��]�1�˚�Y���;�\�f�&��{vݢ�>�4�Z��X�W��������e�VჁ�]��~�^Z�.Sw����4��q�Z�\"$J�h<��u2�3,e4��2<uB	%c�OR<�N[�<Vq�5�j5�M�w��%�X��� ���Ik�L�����K�VYȝ�S�os��%f�i���Ĭ�=�b�$U���.ɖK6l��L��+�-�O��QywO��Fm�ᲓY��ܕ�S��Hj�PA웘 �N�������
�yG6�"C�b�:�T;嚰��Qgt���2f0s�)5���F7�Z7��Q����"����ߪ+(� V
�c=Nd	o�G?���0��G<'�U3u��s'{�ut=��&�y.�7�>�Fϧڀ�4�*�>Lp_9o�xg۩���q���>��Y�H�1ݻ�}O��
eR��ج*��3k�SZ�w�/�vSല�7��Q��*Dw+ygh�3�����+!7���Cit�"{n�>�l9[{�*�c�%~2�ʕ�!F�xmC(���2��$7�d�����!%r���U z���D�^ڠt�x��F��� �^Z$CO�yV ��v�+��S{�@��z���v���<T[�$�Zc�:��wH`��U�d"R��k8�"����u�N�,�jR7�&�O;O�|�煨�x��l��^�3/�iA��v�� �*ɞmD-:��TǞ�=n�$l��>���]���J��(W݆���Qw��q'.�ީ�⾇�e���V�{���*U���b�Ԙpv���>3䖏G��`^�u�XҊ�EX�ܳ��Jx4�G��[S�;��_��i��\�*���WU���qu*��w"G'��מe��룐LiNq��\��(5T��a�ƻ���G���&���\]'I��oj�Xu~��M�+�j	[|G��F�z��>���҃�s)��Wǈ`�K��sֽّ��o�p����ζ�0;w5xJۇ\T4�Nih�.iΨ���X��`tپ1憤ˇ����k��[��	������y��<%���y�?�^���.��[�&Q�r���CjΦ�tѸ��df7#RR�U2:���د���Z�Ş��Ɂ��ƞ�{s�^ٹ%blg�1V�X�>�9K
�I.���T�"�g�^�t�՝�I#�ŕ�U��ᝠ����=ө^N�MEh�t�WL4FR�nfhjQNV
ӛF�E^��x6�\�(��보��z��s/�󉅝�2K1�Վ�B���b[޽���T�+w��(�Y�e�On�*VH,oq-gv�����QW���oR>�����c�pMVv=��r)���Ie���j��01QQ�soD��n1/@fՐ�[W�Y��ż��mV�[VGvy��w��~�;y������Pm�;Fs���q�vcȋ�4��듟nn@���(/*�g\,Դ�mcx��}��3�U���[d����@���+�O+��+s���R2G]�ziu=՚6Q����_�:�����j3;l�LZ��Dζ�{Gz����2���|�&���tKB���8;�]<�2}+�|8�Ɲ�m��zD�&�Zݝ��
�L�\J�ft41�!��6�iu�/�����o�QDuK=�c��H�v�ό�wfw�¬�,�=�>g*��2�蔎�J�V��K#�"x�e��Km~��s����S�/|��:�I��i�u�����Z��yrD_7�����%�����ǔ��.��L�[�D�ǭþ���ljۜ[R��m�I�zs��قSҳUBEh����K��1n#�@P�������Z�C[Xm0� k<�[�nص�J}k��΅5l�}�����K+*�9�,��*3P�i�F�vc�=�齼c kx�w�,
mF��αMr���y�Q�����}����KNY�ҮYh�T���*���Y�l"�T�t��\j�=��"��Tzz�0�a�2�N�˗��|����.�M/w��.y�l��:�0+�oa	��z�n=
�k�Wt�5�L"�1·c;q
��%,������YP�F=��ۓF\���wϹ\녡z�Mb�Au�Tj�������՜�-]��=���$̭,1zl��>���n��I�ߑok}I�[=�Ù�Ü;�P~h�WvyzZd�����zZ�O�b�Y�d�A%���v��b���h��l#�3"��0�OEl�JY:n|��n��G�G�[�ɸp=��(�U�ܪ;&����ۨ��d��9&�v�lǠ�t_WF��K`��4l�0{��7"�Y	U�2��1}�]�j=�k�
�M}�j���7mٓ{�_`�4[ֿvo+�{��<%C�z����ڦ��F�� ��GN#��5�܍q��8��4 � YY���缺7��l�2ӣp�];�JS��W��8�X{��k�g�ة���\(V67LU�U ��[|1&��R��;u}Y;�j��.��6��hM��`�fw_l�,���6�{�t}�V;�m5u���#�P Fi� �[m�$��9cQ�\�u��+��Ú�3E1��8g1��I��D�H�`�]W%޼W�t�-�7����s��@����(��"�
�ѐWy�3QMD�5Q%Sj2h���YQRZ�
*����$*�b"�j��*��)��f��d��*� *�*�&�̭XQMKI05MY�USKAAQ41PTQ$TS��Y�SLCPEPTT�SQјXkV`DU�Z֌�tfeF̆I�L٘Y�AY!�Te��Df9�2�"b���"�3�����XdLQMQE2�E��!����*����(��"bb""
"�"��3�CPZ�*������j*B��!������¬њd�J�3�"�
))���AKa�YUDM������Z�YP�fbj�*���
�3&H*&��� �J)��&��Z�L4QDS�U4QFI�2P�`�EAUQEA�1TS	�?$�D͓�b�w� ڱ�`Ȅ�.H}�d�o�۴X}</#��d=@ܔ^wrke�Y%B�[����ҳpL��7���.$79fwu�:�C=�U��s�F�`9G��]���i&x�U�ayfWӋo�"{�w��h��,i9R�.�tk��z��Ey�%@��bCL�t�}o*�ϻּ���.X��}{Jk��\$����:��l��z���u�z���ǈ�X^��Gh�ŕѷ�ڽt=$W�����|J�=��o�2k֩��u/��?���������7�r?��.^�hwsسgB��y�"8h�keWj̪�R���]�k�H����S����-!�����N�>���N����=�FٱVY��D��X)֕���*D_�o�$�m32�nxw]�nl��c��[��aqv�Ol���Fl���">�砺��/��$�Ů�;7�ufE�;��J�#�<�I���kyKP�}Yk����6�N��Cc�u��g���٩������`8aqrV&��l�F1=cL8����ƣ3	�3c��{�:�47i���Ns�~�7����H�ۻ�[K�҇	�Q�g�>���o�Z����7ѺǦ��m�'��<��	�w��'�mڋ�;	�G���F�g�L��֯mX��jɆ�'.q��l���_Sk�h8�g�Ih[[R�ݛ�^���=9t����ڂb�n���ޝr��2�'���6���w]w�b���6sx9N�R̷g.e'��6 ��wbWr�N��ʾ���n#�0thf�h���\ǫΫZz�N���\P��p���\�a)C����q-kp�3�t���҉X�f5�"����si�
����U��S�u��6��F	��q�C�S�(�yS	�A��@��H���u��{�@�h����F���3ׁ�ޚ|z�w���T���-h5"PB0��U~�l�ŉ��2���о��>��v^΋^��)L��hȬ����'>���b�D�"xM	�v/L��Vx<��1���V�m�c�ݞ�[�F`���*9��i�Y�v��Vh�2�X�3�mg���u�F��%�i���Ls״��^�����S�(z�M�4M<<}�1K�fy��<c���HC�-�*z���a��ڗ�x��_b���눱��<)��w_�ʍ�7�% n�˒�kN��ۇ �X�t�����c���������#�G�����	/r)�sMٸ:]��:l�湏�����	�՟jԮ,����S~�c��8���(�}��j2�_��}�3"�W[tPMXV�DtK�s��L�](�jƘn�P%㬜�Qmb�n�URm�[ش\���1���?-�pw�Z���;�(,Z֜{����/��U�3MhQ�Qgg�՝}.V��rs���]�,��_����^�3)���}��Mu;j穝��G��zj�Gi
�wnm�߁=�q�,�� !u��v�����b��P��Ho�<Cז��<:�54��m*��t�5���\�B��bW�F(�鸌6\��|���C�ٶ�y�n[���Rf���V���\�<dZUq�uDu�[eag"����Q_�y�LZ�蠂��zfя3���\�lq���֫�u"ŕ�āfn;��;���:���0���o�a��}T��{� ���CV�>+A�]BIvhg�'�\8��싉�8����팮i��><�p�-f��d�7�3��l��o�-���C��B�Y���\�#��}r��ƌ��ӝ
��%ġϦ�M�7���=�����.�2��V �!kFJ���,�~{|��&�4�.��c���^�e&�>�`Fĕ��(s9� ����c���>�i�rʜq{\Gl���4���V(v]e�3~Y�ޥ�����P�bL��{�����X�>�MW:B�ʯҜ�3p[e<�&�R�C��Ƀ�ި7��1����b�&pg�M2�j�x���ц9z2�WJ}ւ]r��F��7�r�ݢ�{SJ�(�;��>���JuG]]�˾�T�vt���}}zs�W=��x.,������z7��vh�0n9�bKڇz�����M-�r<
��x��j��Q����:Ƶ/�u^��/�4u�B�]jڼ/5dG�y&}����,��k^�Y�sd�U��$�.��ߣ�坝u�ք'��`���R򵿄���u0^N���kb�����z��g��g�)w��>ki���.���v~n�o���ԧ�!��e�C�D5&S��.���蠯W���0���]�7���!��w�;����#�����U�y
���`�z�Qc��WNfC�ˬ�R����5�R���w�`bO}xU����g��\q%�ҩ�����j�؏��s{D܋�I=W��`���c����1cZ�mU��^JD����+GO��9�x������zk�υ��C�zR2zv3�	C��8������4�$���ئR�.����x�ޮ�Y	��W����5�Ln_j�ζ���E�Z��y�qK��G]R`<C��������X0�{���Σ����b�9q��c��a��J�c$�0��:�Y,vb�`��EMʹR�c{^y�C��ҭ_<F�1`��-�9(5#\���Q�X�b�2m�Tż�^4��/Wd�Tx�w:�m�mvM��n��[Y��!��n�����K�R��Q�<%s��0��wT��+*�|�����8nŀCC�xk��A��׻��^�GI�=�I���Y8�8�my��=.`��*�Mr�n��jK�^e��U5.X�"=w]�[e{���6s�&F��I�uL����lY��>��b��E�^L"��^�<��&g}��y:z��:R���W	���2�TJE�(���T��觇K-a1^�w���=��^�*�A�ӱ��}%"4��>�w�$��S�k=��_n�]�횶���&잖cn���/�h�\�U�cD�S$�Oe�߸�׌Z��g�9Y=�^=(���zx���M0V���Z��>+�������,/R��=^�
�9�y�#./�˯;�8ORW�O�z��´�Mu�rԵ�?��{\���ζ�#�P��qX�	?x��"���d�'�'!�+�ݔ/Ŋ�Uס��v���S�d�{-�;��k���b��}=�FٱV�-t��z����d�a�����O�e�˳j"5���j����q�a�c��5heegfU�}�h�`���}���P�oBb��Q߹����֕��O}yHjVz=^��TR2z�tq�"�L��AU����f�mH��{$ZA���N�L�:*����2�s�1�E\8��5������i����*t/�E���pS|HVa����������؞�_Z�ߛ�n�Ft5�,na9�'��6���o,�P�
�\����f��O!��iҙ^�f��;�Or���r�Xzj��=C�]~���.3�6�y3c��Pw��V'21g<I�֑��v;[�'�G�G�A���tÞb���i/���݁��}������II�eq��qw��A�\ǩ�染7ܫ׼�?�c�G�]�W�2��9�]N���3n�C�(��3@�</yXm=M���E�{���`�����_SEfs��Ꭶ!FZ��xPw�Fh*�Dq-r��>o�^�9���J���]�=�
m�%�5��uu�.��Jփ�*(!<ZHV�\�Ӯ2Ő�X$��(e^6e^�]���z��>�I�`�h̕��U�NHi�1}�J�!��Њ�I�#�)�=^�v��AK��U�y��0�FwK	p��Y`�z��ټ��}]�譊̥TO�}$m+v�&�KF��k���G���v}��w�%t��d�L�YK��ФΈ�5v����] �u]�~,r��3�s�fIʿ5���0�Ыw�{7"\�L\j�;G��h�_�>rs�;{�L�9ODQV��6�u��2M7��8]�7�bȩ�츱��=i��u��/����VwK�pXW����$O�q�Wq���+6���csn8Fc��|��o��fA9�ze��b�#��k����~��c �2%�mz.K�-:lnc𕖱�~�Ӫ\�zU\|C��Q���LE޼B���f�C��?;����y�e�k��\[����VjԮ$x�,�]�eUEK�]��1��3�T�j΂=�4��2��>����3����X�Z>6���@焬>{��ޛ��:���B|���6�Tݦ�k+O	���ṳ5G�yf��!ٗ�-�Vua��wۮQ�<`P�;��mvR��_����J��X�FΨs��_4<X�μ����t�gj>y�� �C.nd,�a�6�h��D����[��v�p�g���5w���8z�����7���ۊ|a�f}8�dJ(o���.�X����PL��v^;���Y���+p���ǡ�%�xW?uA�o��y��|׭]."D�.�5��Jk���fd�����ݛ�[r�Uo�N�~�e���| �Ͷ����D���K�1������9��ޞ��gݧ��^� ��>�K):F�ܥq ��7�3�ܺ�a����(e]J|�v������-oJ�G�A8ۼ�M�0��m���,��um��3�2�f�,��o°O�[�/_M���<2L�7�2[ņ��_k5�NXO2{�m�ʦ��P˞��96ZhN�K����5����#k&A�ee_�a�|��/^�Nߜ�IԙWK�;��v��O�Rk3��o�+"�Ev�{�Y�k;����8�|5g��"�'XD*��G�y�OV�V�j,��%bJ�/��Wf[�R��x�}���&�`���s�u�g�P����ww��e��|�E]�U���2�����B�, z()�v6$�kR�/.�r�~��3��C�bUx8?.>�D�f��\�o'�<�B�Ǆ��M �.� ��M�v�$��^?5�	�&
��#�>����_���[~����N��%*ǈM���C~];Hک��:�g��wI���!N�Wk۽U�9�W�����bt5nX�Wa�`�܆��fg��b�����Mu���f���H�o2�p�XVׁ1�3��0�=J��u�3��~����� �����P���Δ9�#�����KU*/�Q0�4s�|2]���/ov��{����j��V���z��ݽ7��/�N�*�__;���W=˝]tۗ.��ݶ���/�u���6�HB�X��0b.��W.��6����o�i���a��L���{uH�g{�a�����=�R{U��ʪ�*Q>��&��KeI�)�Gh�~�v;��("؇)�ot5���J�D�>�1���?6:� ,~�渷�W_'.{����4���� �DL��]>:61m���R%��,%�N��/��{���7��}�˧�����x��삔vC��g��[ӵU�\˯DF?��B���E���bћJl�tF��
����|����nA���򘬑�Zl��Qg��ӌ��x��g���l���4#�I�8�����x��S��~�y�?���j��u�g"�;��@�;�fO
���i��&���GR�C;Y�g��Vt�ث��y@y<9�˅cs��^��j�q�V�IBj�.�KZG�O�J�*�S4�^�<���'㓓Z��H�����2(^}�Wl���Bˮ��M�I����������ʷ慼	��j�s����j�=ŎӴܴU�s	V��Hi�o��<�"Ѕr���h�޿�ݷ�)�C᧮ [����pw��2n�����V�f,���-�C ��1��^���$�dd���To�O�)�t�7|:e��'Ob�K71�ڂ>�H����Իi��b�Q�%���ۑ鮒ܷ�cB����jp0)\����n�Q�Y��>-�X��[K�o
tS�>�q�C�y��֌�Բ;Du�>��y�[4$�
�����4@����I�����݆}km0�llY�P{3��#�Z�ׇ:t2����c>�>����a3��+�d����^�X���|�][��8���Y���g���pBb��/y�)E�ڻBjMiZ1�5�a���|��.�V�#�O5� <P�rf�.3'�t/�E�+mFl��h������K�A;���O+�^��ܫI��C����O��`�Nn�ʛ�gc5������!/�6,�0g��w�];��z���c��YӍ4�y��l�FL�������ߦ��ɐ�޷�s�Ӭ<��i�#���]�Ϻ�4��f{��B�'�X&=�W�z�����EM�o<�0�c%=�8d�`[�a�,A�#��ԃ���W��֞�=|��O����<��^s;��Ꜿe�e�lǩ pL�K��B���C���W�PTA_�PTA_� �����
��W��������
��W��* �������Q���+�WTA^�W������TA_삢
�qW����䂢
���
���d�Me�Xf0	@�f�A@��̟\�'�<�R�*��QR�����J���H�UBHJT	UD�B�UT��!T�R�"T�R)	(T�!T�$J��aJ�ۆ��Ul�֥J��AJ	v2*"&ڊ��l��CmI-jR(�"�j��̪T��J!�u{<z�kHU$�	4Xj6�+Z���JJSl�TZ�USl����͠U[5heT�Q�	Z-[ZR&���I*�DHI�ٽ�!J)�7�  ��t�(p�⪚
������:`QU��Y�u��Xv+G.ݳm���WY�������h㩣��)tܪYM6�ݪ��:Ԫ�c�R��T!D�� �6��v�ӻ��u��U�5n�#��f�6m5]�[��˶�u�+t���R��wUV�u:k��WYu��3P�ҹ���k���L��%)k)*E%cj�  :���� ��=�x=
(P zw
�B�
(\���СB�
(P���xP��
(P��7xP�B�CB�(^���B� P k�p�Fׅj{+��k����u.�J亇(]�M��N���UQ�   n����+V�vX�v�5n��kL����ݻW:��U�g�]%m�8a���]�LSVڪ�n��RҮ�nUTEm���ζշ\4��EB�JS,�"JQ��  w{����+�Ws�R�V�v�[�vuR�����*�[R�Mn��+*�R��u��tUu��j�p��*�u.u+fm�#��wsV��V����Ф�QB�kJEU!H�UC�  �뱨]wV���*mt��]vݩ*�����]�tⶻe�.���jr��.��J��L�N�4�-v�S��v��qu�R��f�궤�KuT�;�m��&պiWl�Ђ��  {���mT�ۡ�ӧWe�v�:�ukenκg;b�[���gP[��Ti\���Ͷ[�k5����w)j�Wm*�s���v��wl����E�w;[ԪPU ��vض2*��  �{��Wv����Mʕ��F��;uѵ��R�����i�*��V��+�T��W�5G;�pv꣘gThҬtM�*H"*�U�hҠ��  =�TP:�:멦�9w��Y`�hgf�Z�kQm�F�F*�k��uMU[k���*��ػu�ESGIDTJ��P�R��]�  �Ehy�]TT��gkPn��@)jSU�+UP:weUEJ�������k tc������S�*��h�B)�IIU ��F��S�F� )� �SP� S�	���   i"&ʥMF� G�U
J�-�E���E��ƨD�r< Lo��~��[~ʿ���H@�{�l�(B�r�HH���$��	!I�`ID$ �߹��������ۺX�B쬗���Ŝ��V�skj<V�Z���+2��U�5+
�:+*����I`�r!z�j�*�Z"´�#Q%x�Ѕ(Tˉ:��m�n��e�*,40A�KL�GMX��K��72�b���w��,�F۟Yx�Bo#��2�z�e��{!�2PD��[n�b�WHd�kH1c3[�yvat6zr�����M�L¢%��m�;vA���*��Mթt�ݖ��ַi�p��Y+&��`�ҹX���̕q)w���p�U-f��1�����k�N�|լ�e��J�t��>:V,�y�7j�Bq�Y�Pp��ӿ�	?���]�o�4���U��-<ע\��m���, s.�2&�7�,��M������e'�b$��^=��wLv��Z���v��WH��pe�)"s۷wv�5Ѷ�m1�cUe�pi1Sq����̣�3J*Ɔ�UYe=�h6Ҏ!vN:�ה9yFڊ���w(R����`�3/%���7Ӛ��;B���u͓r���c	�' �����aܩD�k@,��c��jTKm�[���\�Y#���0���˨kb���K­Qݛ�ni�62䆔�ʫ�gmV��,��E�ÌB�g5tШ�ɕ����Mh;�E]�) dr�=�՚Q�hk�	i�Wz���B(n�h`N��39mT#v*ǥP�!O6�i�9�dZ�˰�br�,��ŀ�f�ۥ@8ձ��Hn�iڙ��Gؖѽ���r�l��V� �W�l��Y�iV��̰*��
��PonlP�U�e^�Y���t)^ڣh�/�i��cZ2�~�E�Ťf���C��I���Z�	�Mem� ֌�zŴ�+.�O���pJaFiݑGm�pfp��A550;D)�y���:SoLf;��(�I��23�WKo^k	#���qlF�������U�gR�b\�i7&�����Մ�%!co�f����35�.V���(rHȻg`ڍ��b�~����.F�C�*,�T��75��L�h;�r��d�D�M�נ��m��%V��U*
�n-Z�-�ʻF"�4�N3V֝�w*:qa���\Ol�:~4`��x�:�@�лm[md����w�b�cs��"+%��4����Ɗ�M ��S��w2\��4�V����e*��f\�r��!YY���KN��jTuZ�BTǳT�(�4�(ճGQd�Z	��m����fd{�nB܇/U��+�DVjRc��1������6��t��;�|��W�]���:v�*cX>�T��6'
ܚ&3�� (P�uD�f��Z��^Ff%nd)��{�]F��,"��J����u3w~gHQm
���_@�$��M^
M�2�j���H2�7#�hD5�HL�N���J���p�9Zz��ܖ-�3F�T[��Y�-��7eh9E%[Q��c�U�>i�,��I[O�0du-bV�"��V\�q%Gn��EKupm��&�[�S��nQ�K���N]�C�Ց�d$�fSY�f&(̖s4�8�:����1�`�/2#okM�Ĉ8��Z�>y�PH�c�2m`{��W1����m��F����ǩmh��`z�f�sN���a��n�I�
V���^�m�˱���H¶�8�eɖq'@�j��-��(fPNf	N��jU����c>�Y1,�4��5L����Z��Z�So~4���NcF�Hމ���)c��R&kC۠J;Ikd�%ltUm!XJ�9�u�M��K"�4d��ݩHX�>H��{)�����!L>���X�tv��[�BV�"�V���#�10�'r��s7�u��#hi��R��f�����Yz��'�%jrVL�&��*� zLj�'p�����	�n�JKR�ҺiY���n, �glM5��w��k0����{j���+l��c�J�Xn�;x�ԦUc�v1Ǩ��l�o
����Gq�["���M�oU5��˭��BI�
�H�BB&�:M�5-�ZX���|m�MV�%R���${/l�N,-֍�I���_, ���+`w6Y(��f^x�X�j^h�����(}i�Kb�-�%�{2�lqHI�xe\�W#����@��-���MT�v���+	��Qv��#��qMY�w.H�Sj�y����u�ֆ0A�AWM^b@�R(1�p�Рq��	�0̼�`����s����kE�۫���L�m���Awd$��׵��^��G@;Zި"��e�Fheм�	T �xtێ�q��L�������.�K:����04��lB�Q�x.��Ӱ�2m	��R��.Z-el���n�٬��u�# ��k�Y(fV k�������ŷ��/D�ԲMyZLvD��M#e1aR���NdehU���7B���bi��bXܬ�r�%���p9w>��-IY!R��%���XڂFw+R�c��{�RT����V���4vm*t�|j �T[�2�f�%����u]j �2�ͽK�I��0��t��Cf�	��(=�(�N�ͩ��j외���GJh����rPK
�T��:v�d�]�S51�^��&)�r�ژo� X�)�@C�ں.�M�`n�&�d�3`�ޢ�&�bɎA7D���bԬ� �dcl�� VD` jGY���Ƀ5^=�t`kM;��N���C[�A7g"dk�!�\�[,�I۲-k�)nj6eq\��*o҂;�Vbǅ8���1,���f���,�j�86e+wu�J��R�%�YYkM�Q�O�]ec�t�1��
�f]+�DAdJ(�w8��J�V�L֌G ���H�Y�%�!^�M��Z1XV�i�*E������ÁY��BMKt����6�[j���`���i(),њ��Ѵj[��!Ȝr��1%���"����N�DIa�&ˍ2k:br9t,�k�[b�=_h`��W-�rR���lPq�͹��S~��Q���r��'��t����]e�٘���ͫ*�0���e��xP�*Zۦ��O,����;�Y�,�t�"�M����_e�RK�Z��O4��L�֪�!ue�]n��[BX��&�n�aX�ʘ%���s.�[�p��"0�=ٷkd�R��v�f�:TYm�*kZ�ћqֈ⺛���P:D���n�*4t��J��i�Ȉ�Ċ���6�^��,�٭:���z��u��delCeJ�L����V>5v�V�wZXdA5�TC7c-SZ�:��B�L��=p9.�,+m-��Za�-����a�kj쵗��|��&Ea�A�eIqj5�Z����*ң֎)�R�n��*}2�W�
�wf�6���)V�2]FBHR��ܗ�n��Vɦ�/%����N��U�`z�)Vkt�ݵ��q��Ҽ�'A��u)
�F�Mm�s�V�M�3]Z�y�����H�/����"�SyY���Zm�Yn�
i�ס!z�b�6wilm��=�+`u����ɯ�Uc�(-O-����� P�uQ�$��' 4�e��z��=��Z�zJאͤnÔ舍��a�g�IO����viڙ��KT��s$�q�k��$U�O�w[��2V�j�$LW�y��FB�1�����ۥ�M�Y�M�C/T�urF��,���9z��Bol��W@7B���]i�u��zb�F'��{&�h^��b�K���м�>}��1o��V����E�~���t�;��0	(ՠiO���kC�e]����[[�^<�B��WO]M��j޲
X^�@TtJ�Y�uƷ)��[�-�M�3$+,�ܣ�b��H"D�6���=ڊ�\�k�˸�:5�7�2㙭2G�ZŅ��H������z"���T����ɗ�@M��aD���R�8�S Z�̼�*��όy�Q�5�˱`�vB�ɩT�`.�c��kzkUj���t�i/!�౷��r�Cm��$�з)��ȱ5��A�7&<�H�֟�8��Y�a�Q��y���s2�r�J�0Jy.��C%��b�l�إ&�.:N�yM��4�w*o�\�Qə��V��U͗ʎ6�<P�*�܂���ut�1lY���7������]��{)n��{��5dK�ZKv�b�ʈ��f�8�^-n���5%�.Ї2YOE������֗��#��X����mj��/!�x�V6�@���Op.�W �Y����Ç9B��7��R�[�c��$8��[S0�FS;��
Z��t�E�@Z���[j-?G�l�(h���jd:4Zu�pҙ�ܭ�R�I��Yee]�55�%bו���coM+
�;P[ů
��N������e4��\W�QC_�TUi�d�q�yx�R�m�77i;2:n��hեM����#�M�̩�V����B���8n���F���;��w*�Q̧cN�ث1�nk��e@Mɒ��ġ�z�a���2�Pl�O]Y�R���*�Ч�i�{��0Zkh".�Z��9q4i�%ѭ��R��X7t��� �;;�*��0f!���ַpݤ�V�ĻV��Q-����B�Y,'�B;yk.��i���C��R�Qc 5VT��-i��� )�0qC��Q���{o2�z-�Q ��:�Mn��\�I:͛2��N�͡2�Ф��壎�Yh��i�;�q-��)=^UՖ�ވzT��
��dª�o$�jʬ�b!�U��YdZXm�b��mBUKn����%e���x��ccT�bx�i���O-�j�����l42칉�_��Ya=j���At��������sT�dؐ�Z1�z�J�v;tɦ��ژ#�+K�dlQ��B�3x�8&'x��v)�{��S ��sm�r�tѧ%��mKW�lO��-�w56]�4KA����ƥ��YN�&�[���~���3/4]]e奏^�+AC(4#u1��WDf�H��Z"������ kJ7t�$^�ne�蚔��ּ�*�2��e��+b	MX�
=���ݝ��Ʀ��N�fXy1:�gw�u� ��RrI����J�5�LJ�W�ij8�5#�{e�jGSgaF�7�̠�`m�T�wkp�!�Y����6�V��/��<���octF�f4vE`Ьrk�9.LE:�@a��]��/���ݥu5`n��*���ti����lxƻ2�K5ee�n������H6[�wV�v]�&��*Č�3.U�cnJj�0�լ��rl�YRh �Ud�+h�D֊�K�xئh#!���uZ����\N�ЭE:�GⲲ�:$��������Y���M:a	�4�;��7�m��kX�IV�JY������J���W7�sV9�š%#zEJ�X]Z ��kV3Cݣ��!@=��p��*B��̲��7�W �y�U
��5RSDMj�+�����*2q+�oa�m���嵌4�� g懥�f���A�a�����2��(�ke�d�m5wq$~�/4X��-0C��x�ú��U�y�v���Yw�[J1�
:�;��K.P�m�ۛ$ܩ��@M��b[X�rR"PMB�)��)�e��K{�3[@��n
�d��f6kK�����~r�Sse�,��c@+Iݶn9��Zv��f��h5�<oi�k(�s3-:Z3@dٓ*]&e(*���7r�d�N�h=���Hc��:/a�4���T�7qZլd
��hDjj�*�<��v2e���UĨ=��;��T�s-+�PĮ�3�?�@�.���0) ȳ�-�(լn�zl�3`V]vrJKo����{�%��+tcl��p ���۷�r:�/ܹ��O4d��f�y ��d��A](dݽ��`Pp��[�U�y/Y��S�˺�w���ŵe0IQ�Jut���)*�,�聚b��RE\�T���[�Jh��v�c��x�Èѱz�)-�Q������"j��唆!�v�m2�Z"�.c�WJ�Cq^)pi����e��]�յ���VB�C#U��C��˦Bt��Y�7��ɛt�ƃ1�Z��պ>)������F�B�~{XXYeB��(�`c�MR}k�G�7QR�۷c^� ��P�

�ڻݢ�r�(M�C!�m��\i�-3OJ�Z��ٴN�*8F��L��Ve
�6�˨L���R�c��)�.�0�%JQ��NmJ`n�v1��S�6m8���آ�����{���,�br��HZ�,\�@]ʷ5�	vE�	X�B*�+@J:l
�Xol:S6��0�SW��"A�M�X��Yi��-	�mH�-�(=ev񚼴�*�L�����*d��,8Ug���h��1nH����Q���0�q,��n�S
�ej��\�rCh�z2Jz��;�b��L���`�E�D"J�k*Yշ��"�Y:ȶ���A��z 2�b̛�Nf��/��{j�!2�R�d<2�Y��� Cd͙�[4.
�J�;�IaoD2�n춉 �{6�V�-��;�e�8M�+X����u�Ds0Ǎ�{�T�z�S��+�F�te�)2LTڢ�+x�n�Sf�A݊�n����"�h�y��]���Ӵ�u�SB�n9�T���^���q*J�׊�z��Bf-P�x��6���E@,hv�d"�3:\4�����M�3qL �UjΓ��ۥ���ƬAm�WH�۠ 1�@W�O� 3Fb�j[!�ц;�D*M�[��h]��#�L<����X�u7�E ?<D�Nݽ���V@��h����k�C�nl���F���x�f���-#���1�(��t)�vT9HT���Y}��P��=8����o��v�{�1�*ub�m��M3���f��t�P�Պ�B�L�������8F�]J��yA�+��{�;��Dru]I�jP�(7O�X�e��#2�\}|���K+_
��v�\� ��X�v*�	�c��7;!va]h+N]�	��f�v���ܹx%-ĺ�Ru�=ՐD�_m
<�q�}����!���t5K9*=}���`��}Z�|�3!��C�����/��i3������|�0R�#��ۃ��b,��6�W�Ʌ��[��:{�Es�VSTM0��֫�a�v�֍�P�{�\nK���.��En�Jɕ�/����kh��!�� �9B�d�h񷷛s�3�AB �
�dV���:ZX�!�M�g��R�$��$��oZh.އqƓz�KDZ�뉞2:��J8����)��*�5��n�O�HEw}���+ko;����ku-�.뻬
�)�b{�����R��F�3mI>{}qco�E�k\f��t)�4b#�:�m:+j�u�꽮΋��c�v�C;�Bw�¡���n�4����Y�H�լ�:88��>�l�^�֑��5P�vwQtje_K��r��͌���Z���*���	�f�;�4���#�mGtqƶ�0X�X��'�ǃ��W�\��׺�E��@큏mAJc=�pN<�p���ii2X(8����1�;�M������������w�Ȥ<���8���M�Ȧ>\g,K.	Ҍ���=:M�3_U��4�1�mT�����h$����)�\:�;c��l=��Zn��]u`�X���.�]�\��S.�RTu���/�9d�۾�b=#U.��fֈ��z�ż������� εC�(r�2�U��0�r��O��b�{0��.q&�_s9��k3V;���G��`�"�o+���U1��EӲQmeJ��r��]kq��ꮟ&p�B�,Fĥ�b�Qh<�B9$�n�Y��r��+�H��6�]b�M���Y�΁��v�n���w�8�ۓ��q&�f�_=�5i���A�������]'\�!�"�mfN�2��G�wtN�%��FS�}��!417dq�R�v^��rq��=|0xYN��U���ve<��U�J򤶵�ā�	r}mw�m��,�}9<K�܄�9�-�J��]���������&��X]����o�ufk��N���3�?_�q��,����5=�2�={���$g+!��桝sr�e�-�R�6��p�n3�G\C�9R��UcQ�E?�d��%�2ukf��y.��ru�ƈۺ�\���vaeh��d';e�9�[<�/F��4w(����dy�9N�R:���%eA>�۲(�w�����i�S���)I�l��ӌ�ٝ�D�	�>|�
�(�(�8�]�z \D�gm��������3�R�����c!��� �CK&�Mk�Jû��\��=BЇ��ݒ_��#�3!�V��j���b}��{��(,��,�vaD(�Ẃ]V�hR��ֻS���o�J�m��%��������5�D��Ԩ�8N�,��{�B�Uʾth��lK�1U쨠��-�w�!x�̕��2ػ���G�uk��R	��VԽ���](,�EV�*ur^����s͢���Hhh�bb�ݪi�9.2ޛ׵�N�	!�Mu������va|�ŻX�D����=�A
ݷ�_M����-�+�&�Q����F$j�PveęT�=���.{[P��-6`�b�M���s��r��0���N髗�C�3M;
���=Y��Y�b9p=����)��Ӯ��;o�2<iL��;w�w6�[��J�&��ݲĦ7��7e�a�"��̙���j;�Ut%��Ţ��v�7c����WK嵓 "!ۡ�*˳uu�NcT{���a�⿮gշ.�b�r�MJ�+���ԭ���wns{^rѳ��.&�nN����k/8�(�d7æ%����{p5�G�Ct�12��g;R�=LQ�5L~��nA-�l���hAM(��Y6��.�[96Z�zl2�5�3�����^���{ʣ����=ޝ��6���ݛ[vؾICgc�P��:5��qٷ�p}�%\�Hbl<ݻ{7�����4"G�*`�T¤ge�-θ6n�!����K�4�L0L��ټ�l����Q8�E}�tD��+�6�:��I������ix�	+��ە�)�/�w3Ib1j���E>Ej��PftM��$�GU���oA�[#�A��[C����[��m�/���WWi�tv���nz�����`Ũ�j���B�(&f=8U�3{eu�w�^��~��V���jpӂ�����qI�K��:������Nh��Yz	���]�	�5���vj�E����5]���J��k�[zn��{�$3�.K�modZ�$�"Q:"�ȯ�N����� Qu�j�e 7]0��ʰ���l���.�`&�e����Q!�-���Y��{C����{�� _72���̽t�;�T�g)�j8�K�s��u���TC�&��sQ5��^%F��g�+Wevp�E��V�ٔ�l�w_#�M�z� 6�к�P}5O���ǐ�v���Z2AA��j��a�Ⱥ��V�.Xz������*���?���mHy���rW��Ұ��AŔ�d�1Ù�w�NE�Ŷ���R��zZ#u�۾�n�����:�9�|d@�]��j��K���ζ�gJU�Զ�9����	�bZܫ�0ɯ�ᬖ7Qu'VZ����[�����7���s*/�7��.�5c�[6jwK$o���<%.c0�΀�3��Y�0<�܍p,�u#B5,�v�!�8y1G��7����8�g���YR�V<� ���g�N���e<��F`���b��@�U��q͋�H���2����c� ��m!kP���#.!�#��]��;:�ڛ����/� ���	�JN�PI�D:s�i�<V뮁%�Ĩ�r�[;qb�؆��۝�
�}j� ���i5��<�u��|r��^��\��[�������:��mҌ
PFV4�[���{�JO�f�-h��rĮ�aɫn��{�woGp�r����*	�c�t)��q���v�h���c6}V��C3�Y���P�io,�'b�2��'r�m<S�.ۣ�wU\�ڽJN��o|4�X7�rAw��ڼ<ێU��\�w �{��ŻG�]�QI�3�b89��ui�1�q��'L´ۻǁ���gl+����+ ��B_�x3\�s�cǣɉ�E�o�i��;K��p�뾃��b���Y��L[NO\�H�+n��K�g�@�R��k�U�{��PS&�]vU��w������k�;%����;o�9`<��͚�#���j�I�MSӢ<��;{T����Mw9�ҷ0��޼�HE)R�\gh��.��L���Z�+9�h�"{�Nl����1H���$�3����tȵOFZe��<E���� "!���P�����b�iA���38ᚪ�Kە�\Лe��pۧz���@x�Q��Z��4���	˫l�	\K�̑S�F��=�]���*��*�遜���Sʝ�%]'S�nf���ntTc7��yhN�+��!f�,Z�st�d�����WhRq�@1P�ڽ8�=B+˧}F��0��f�������{7��'pŏ��$=�3A�TEF�]*;��G.��`z�y��8���n��W:{�]�F/�-�ڠt6β��5��lc/�EoU���rћ���G���˦n��8�1��&��#K���'�VR��!���<�5َ�
����2���u�ngZo�P
�s̂��c�9�v��Y$��IO��G��üsIO�.Ժ��6�.��Y�MՅ�A.�ϕ��L�x���X�r��u��ҫv�]�������DP��7c��������,G4�W�z��Ԣ���ߠZ�ƳJ�emy�2��aT�3�v,�}v�t��t�(v仪��[[HwW �˻ǻS�p�ul@��B����آ��^.�sj�X�@PC6�>4�	��\�y�����P%S�P��ύ⼥�������	Nm��>��qý���,b����h�2��n��e�l:ڭe��M�x3�w��V��v�o[���ݛ�εk
}Y�����؍�暘%�W�=��z��a-v�
����dp�%�ܤU�v��n�x ��i9�[e�^LōФ&�f�n��3mb܋�/���G7,}�ؤՇ��$)���11�Y��%a%�	�����ݯm6]`�(��36o�V'�S8p�3�RL)�����DsX{�
����Τ�(�X,M{\����ٱ�6ȡ�t���Enh�͖ xiCor���.�YQ���Wm���=4���Uի�KZ����Qϲ�wv�
�N���P-
��{/G �ʙf�x�=��!.̦ͦ�{�MOE��v����������:�v�fVy쁜]6,�s����p�aFi�j���ǰ��#�`��mm}�;Q��7"���Y�e_-{������:�W���m讗�\�Ƙ�v��uL^� �'3�F�uK`�����mT�51u���e	RnQ�h�ν)�w[�S�Δ����On&oڊ+�k�9T��tR�w&���.��]9臊�Ir��*h�{�1j	��Ը���7� �H�a�]�VR� �j�@�b�K����	��Vp��r�5}W���l#baD�}��wPk{��r�;�7olX���&�R�|�$�n�)0]՗r�����U���TN���K��p��z]������X�j�s:WPV�Wµ�Z�U�T5y�m�Gs7�P�Cz�{9�̬���o)�Zӣ�0WW�Lx:���iJ'�ct��l�Z���E�c��d�T�1$˭ܐX;b)=�y�~�HC�S�y��3��6�h1�	�z��e�m��-{|��Y�X���qU��xy2Φ�[��2���4wf|�m���X�=�a�Պ;3;�K�Y�5�� �Jʍm�;'k9S;ǶÛ�g�z�ӫ5+M=�cv����mE�ll�R���E����m��n�dy��u��<�W^����;ՙ!���)��S�4�H�q蔍���ڠb���U���f�����F֐%>`�T�'WA�J�=>�,4�z�2ŉa���`xn��*L�%f�ռ���Ȏi.R���P�w�+-\;l,��;&����]�md��H dj����2�!���6�w��=��l[[i���<�h;}\p���i�6�[�&�@Wj�Y��B�Փ�F�3f���	l,����@\�:��Մnժֹl���`��a��oz<5.J���8AS�Lܠ�Cg�>�Z[��ϲ���;���뚂K��9U��Î�"���)G�@�ʆV������R��*��u��Sᙓg(:�T�Z���j[��Siٶ#b���Rg���!�1��2p�����M&d���r��4xp��r�H������Du,FJ
������2cnB��gjW(Lok��ƋҴ�XI����������*�FBI7��V��4ܚc�[FT����k�H��u��p��γ�.커��Н�[�b�<�mn�=f���B���y��AJ���}�;�8�]�oxN�{V�{Y-`�X)R(���A�����n�3s���о��j�fg[��]�Ȇ�wr����\3Xל��N��}[����/KR��y���b�a��k��3��'�+흢�8.o�Ыy�W"���s���A�O0�C˹׿�TR����IO|�F����OwO�o��@+���v�<Ӡ�or�t���t��0N�i�1�ʌ?����V2x)�xn���"�.�5�AW�Y���{wi��5���1�f�l�m��;V�l_	�X
����e聚͛P`L��k�2T<�c���]egPp��u��+U�FA��l��a��O��o>Vq�9�cY}��TE���;��P�n��OR�]��k��}���5�C�S�C�(^R��0�3���,S�ٮ܆8��1>ɋ2��`꛽\!	1R5�E��k�H�umAfnh{u�\�e�Z�K���bdT��S�j�K�Jt�^A�[�K0;De��aeo��z�i� �^���/�Nq���Y(�uv t���l�KdrM�nV+lm��)$�O�^�������ļ#���a�6�; 1ϫ[s�P����� ��"�m5��9�Π��{{��\*`�Y|3��hwu�tnu͒�^���ņ��(Y�2t��$˲h��o\�0n���G+��sF�1%:�]��Uf���,�7��2�o���ʒ��T���Gu)��yՎҥ[��|�5K����ZTS+@��M���;m\6&��>��P(o}x
C*����,���u}�E;�|酙��3���2�u��4G�Vc�<��r�3U�g\��%]�RO�"�w���!J����k���pwWZ���R�9����QGU��lm�y��/��`���N�g!9��W�$��֫�>��q��ؿt. �y����{{�ܾF�Z�����IvS�0ǐMՊ�d=�{�rt�;��4Xy�Eݽ�Kփڋ�ݬ"*A�2�x�?xApH�9�ɢ"0Cx���|_t��[���Cm�|��Z��'�T��$�,�/b��l���_Wf�'5��N��RΕ���;�d|�e����>��+���})#�,Ir��ԕ$�V���KR	$/.��ϻyt�Xy1��=����%@'[��S�c��]��7�����������B�;�����u�|�5R���u�{�_����x�B�ݛZ!K]���T��o\�+�����W��E8k��4��*���[PK�x	��(ܱB�z�xm�a����el[2+�C �:�n���R�sѡQ,�g��f���+F�Y(f)q�x�^����ZLN��f�ӗ��7�R��W�M�Sx��F�Y(gУ�k�׿v�">P�B,��ͮ����3#�J�c��	�K����|s�&����Q���D�k1ǖ;��f��38pA7/s5�yC��2�xV�Ѭ��>(	J�lܡg�q)�%Ϋ�(صn���g1ú��b�7\i����i>���B�p���jjtŁw\g�;�� �ݲ�fǙ�;�:4��ₐֲ*�-�L܉
�yWv�`S2ؚx%t����5}8���2��ʎyp	x�ͪ
���zD�RZ�S0�����T��"��V�b,Z�]qD;�w�պNd��aڛ�*KF��&�����f�*ѫ�/ڒ�.vq;��JR53�:�6n�o��M�� �̕����Ңy}��"m)�w..�7y��S��9���X֮�䶷�ޚ��i��lP���_-̧Y\%��p�F价l�
�.��}F^b�C�%��mm���Q" �!�΄>{�6��|y<�н],��@��r�=}�o2f\��pk~���Y����A6���>pb9مؼ2�iY��jp��Fu����G6c;4������+4�5��;q�����Sh�g,�c�_V`�Х$N�c����|�H�}�̆�\�l��a�X4�M�e�t�lpg��u������� Rsǎ�6ur8��C�ǔRQ����,4y���n�R:���5�Zq��W[Z��h˼Q1D�Vs�ʻǪ>XAɷ�n�o�s��b��Y�b�g�o�� ���c�"}}9���y5�Qf�q�Ff� =��Nns�q���n���W�	i1qkH3�ժ��M0{�s�[���]�s�I�wn��(뷉����U�i�{I}S��Y�ēSL�����L��n���a؀[ˀ��*���o�+	�[M/l�|:��$��{��'3W��i�yQV�l!k>a�)<'�Jһ��ޝ8è�-��� �y�I�֊R�"�E)�`3��;��=C�k{�rCZ@D��w�j"ѷ4z��7=���CF)W�x���G�n������wZ���q�Q3M�]��m�O��U>ۺ�oVܺ.S;����[����k`^�5��i���7�6�v:M����S���)}y�����W��޹�񝻫L$��ν�yIFn��go��.��/�fs���	@���|�tV^�x8�*��>��DN*����9���ɱ54��fM������|��|��fMƕ;�����υQ�c�2W�I�~�v���9a8�|���
��w�f�dC����<T��}���D��w�4�Č�of�coK�{s)M���@Wom�l��?���ڄ:���v�n��2�;Y�:�KT�-��Ev�8�0���cP�b@hu�y��&�N���o� #��{��FP-�|��_u&��+]�Ί�E�A٬Ÿ��wP�̏���]+��_]a��[(�b�ƹ�	�wY����P�޸�yOl�u��6�H,�j��	�rV��s>�3B�'Z����M��ʇl���8���e��1��q���3�D�)�.�	��0���u����[�� ����GYA�����;���+�j<�8�H�'n�@���gf9�`Lb��Ӓ�^�p�2����٧��2T�wӹY��K�0.��E��h�I�g$�}vs����X9��N8h�P`�M�xa4�z�v:G����Ն<����ב֖�w9˳�d���@��A����Z�{�a�Tc�L���Z����J8�|�����3�j�:�|���WZop-�3>��M���@�5+5n�Oyi�1��u���w�1��n%qI��Kp�C �m�=��-����b���)���Z7v�Һ��ocd�,K����[!��RK�(.:~�w�륆7�en�ܶ���I��7uF����Y�u@T��G���B�˫$0��ѵYѦ��w;TNc��W�,CQ�C:�	�T���%�hA�x�]�S���Eg����V$�6��l�i�N9&����p.�.f];�`�2��O\WX�h�Ok��[-��m�j���<J�:�6�-2/(�\y֙Z�t�q�2ӧq�`f�^��t>���`!�����Aώ++H7P<����յ|n�1��r����e7}(c߃��Y77}��Ԯ[����-��ގ|��Gy'i����"Uays@�6vM�Y�;�An����z���Y��9���E���x������1�w�x�wW�$��0����K�����H�hgP������<&�;,^�]�c�\R=7�*Z�Z��R|���#6Tq�5{'�0kf�c�����"����κK3+HN��\8�U���?8���j���]���YB
H9c0O\���=�䷲�_e$�ú|�����U�w&��\+S�ب%ݱ���|��ېn��9�um��T=x�a�ﰷY(V�!p�q�f�C�4���	������2+B����Lˡq�E��1�=ۤ.A�;��Y��dq�NPbt����\�>_���{oQ]M��Z��P�����P�&R7y,6�����h��걵.k�7S%���W|F3hO7��
t����{bR�κ���DuaQn �
l�]m��漶vT��_]��Ӳ�F-�ݵ��^VR�k;4�Q8����"CTi\��dc�#f^82�X3f䉺�!C�T+M�i����;�*�k�������9ėd�W��Hq�%ԨV�xQ�HŋUL�:q���kJ����Zv����N�`E��������\�{�.ԥY��QWx��Z�^�У���wQe�?+��B��EM7����9������7J�P.���e�0�c�[W���n��E�a��Җ-9�n���A�}Ǣ�ܬT�R�����"�˙u �bjS��̘�,dͤA�5�e�@u0�3�Z�Qu9���Pj\�Ju�w��A�@��Z$8�d'�=�K[7��p�PTL-'���K&V��B6�i����*cf6.�B<�J����ʆlL�m���mnoJ��]���k:���j4�/N�[���}��Y�g�)����-��Q�on!�
������M\�k��Fn��"5�,��2eY]���'�r`#y��k��FW0V���)Ppw�Z���2�K���]	!=�v�>�ô��ܢ1�3՛j�d�-�c�7��9Y��E�J�-@5���W�	�H�u�%�A��_w�--�te�x5�ӻ$��8u��X4�`#�q���� ��c~;��:�T�:����;�n����Hr�����\�^�n��QK��(���a��hL(n�G;//��	F�Nwec�-`H�uu�n�Zw6n�itb�1�����lm�ږU�5���Ǣ�*���X9r+�ֲ����KLd	���)��s�Q��9��Jo��g��V2�n�kl��vZ���DU��0oU�*�F���f.n�yn�LTvQBZkk{]@�f��
Y`wu������oϊ,�����*T�Fm�Y�0m�-�Y��
d6�dDʛ�zkv��˘}<�8@�o7ZVj�,O��oئ�i�u�<�mj9,!����:�z�O/�f#D{*�v��̔�-���T0�ʻw�co(�,[�\��q���f$�C��R�ڑ1lgd*�wNy���ڼ�Lk�j 'XN�ֽj���ICw����e���7�e�Fֆ����
��L4'>f
���y\1;����vL�{�n�/{��p]���q�cB�u�$aU����^P�b.ڵM�5��p�F��L��3{{ϴfW�Yʸ���o���``\�ǚj���f�o)r�.�[�In��
�Ek7�Ž�rL{\�o$���kp�v��t��4$S��6����dn��B�4=c+	H��'@�V�]���N���! e�+X�"�Z�Q
ٮ���v�H��F��g�T�s]�w̭�Y[Yz���)���:����y��l��YI�T��P+��NA[��I�O�m���)�~kٸ=��	��%���eE�6�Aj�7d�i�vط�y+;o�&�Mդ��`/Wl����|�u%k�,� ˥/v�
�Ң/2��ǹB�N��;*m�[�Tz)�k�3j��J%X:�u�F;fq����nj�Bh}BK��Y)����蕮�f�o-�A�`[ݖF[�J�=B����#[1�A�T�(=��*+�9��3��m��)�ͨ��u[�� ��B�pU�#k�U��d9]�V�o%�I�v��)n�����Իlv^��U�ii�P���[d,ͦ�-R�`�_4icX���J����f�6�5��F���h
Ve>�m�db���C�k�0�9�t���`�[�0��V�����a���D��a��D���L��w�#�nݍ�BT%�7��bn�{;^��<�AM�K�Eˡ����!+�ov�]����h�F����f;[�$Г��w:���6��m�Y}8�+X����pd7�7��G&p��^ax�'M�A�����s9B�'trti^T�[�cx2��2���q7��%�J7x�&޾!�)�ް@�'�0u{��|	,<{G6����Ryv���q��WD_4��'n�Rż�gaButp��f�Hԕ[޶���h_=�B�fqղ��)ի]�������sU��̙�_p\��n��,��(j��K��LL�L���J,0�wN��]��A���j��*Y��I�W��їa�xA�F����j%T���R�0V�2��MmmE9�5+�f���f�Z]�	�S)k�	L�O${}��:p�W�"z,��xD�]��z�rr�����t����2�)2-�X��GS\����=&�aN�F��q��Vi�.��G�.���v�Z���uwO&���-���>鴤����3|�Ov3Μʃ���v��{2�Q�С��*G5<J�[#��HhX��)�Z�� ��5v�t�S����H��܊m�v��j��^7��Ϲ�Mo{:Xt2�*z<���_^�t@�J�Y�Ӵ�cI�䮻 ��ofa�S�	sQ� �XZX����V�7�Uʍi�83��J� R��]�B��`qVs�7�)2�	��:�i�<�j��:;��G�W׹�1�{	��	ڂw���a�лu�P�넨&�����TX��;z5�#��/iά�[�r �����-�&GC���g����z��;�fR�miA�K���ErG��9�/8��.�i	P�y��)����2�~UНԁ���4俞���>g�S\��u��7�̕ͅ
�����ĕ�]�M���W1����G�$�Sv�nw"y,*OELx��xf�����h�e^��2��B��ᨹ�ә6L��8K���.�j Ž�\�ŠB[�he@f[Wrr����m��Yv��7;
��|��x8�k&WS�,���Ót������V�mȝ+��p9�c�=0R�:(X�u�.��J�N��[2���`@�t�S�N�y���;DG��K��]���%J�)CJ�5���F�mTtA��X!�!��a�Ѿ�,��I��P*Z�sa�3��]�ׅ�!�!�������_4Q$��[����w��t�Ճ��q:K��z[S��p���iI��1w�+�DJ�]��G�-��j#(���|5Zsv3'c��U���m(�������Y�N(��3 맵�Iŋ�^ɚ���e�C;H�KP+&ZMr@:��4����A�zzU�+�ZTbJotW�i�ۢ�@�F��G��������k�]Ba|{jj�ψ�U�4����6U�M@��<*rO;t�C8(�� 6�:�!T� �ń7*�9Jm!����j_1Oi�Թ! �y�VWr4�<�ײ7N�T�z������r�o��7�};��f�n;�teb����y�� [Ąu9]Yb����n�+����M�N��c!
�%�N�kMi�kUv��[�	h��։��Tjr�����t����^�n�\�M"�\�k��yDWSz�5Wj��GM{�%�\��׫����V�p�/)�!N�0nS,�ݴ��_^=1iX't�CgJp)AH
�m����Bǆ�_ב8�j*Z�F�:�;yn��j�b�&d5ϳ]%����e�j�d(:yϥ,�z�y�j��7�ۢa�f(-�	]���bWC=; �0��������M�Y�L������r� ˷[������v�__J���4=�,k��;K�?���K�r����"�{�t�;�{��,�Z�1���6����tI t-�9Cr��������x�mrժ�:hZ�E�����hbsj���v�F��S�ٔ�
�Î�ep�X5����; ���u Χa��+䴩%vpad��U�4vapc�H+��;놣}��1�	ڛm��?��u��'��f�8k�0��F�����P
R8�^�s���;�c֮6���&�T.��/����Ⱥ�ѹAV�&"�O��l�����sgbu�J�Gs#��Z�|p�y�bu5�a35�w�:���c�nM���Cp7=~OLs/3�U9�m�x5�[��4���0],�MV9�o�uVƫB��9p�K�lY�u@sg�9��t^��I�$���ɧF�y͐זde��:�ʯP�RDQH�����=��yq�\F����|��%�[��0�F�6�tZ�R�wq���S�׽E���F�Rܰ%��mp��[�t�����t�H�Pu+0�<��IV�{D��I<A���t� z]�O	��E,l&��q��I� Tx��ے���^��l���ү������Q�KI۫Ow�ъ�K�k�Pju��ݤ��t����>����Z鹪��� ���SL�D�3:���>��V��bﯴ���_p�\�O5�2)t�����:�γ�?i<�K�C.��l�\��t���S�s��j�g�!Ưj�L�H7c��ĸ��2���m!���]J��m��ǎ��dvWt՚���
�i�VTP��ф�[�k8��*�����]�͘�k�y�*�N�&̭r����!� �u�Z��E��}��y����F��(.�1y8>�g\1�ɔsö;1q��7F��,�`��w
�	�WPtG�{w�e�7M�ƪ�n��
�~�18X(�ϲM�Doo�o>)�P����+��cSTZ�[�;��2�+R�-@�>���ݼf�#A*��� ����p�P���E�jT��q�ޢ�<5v��˟)�7K5!-�FG���4��m����kWZ��k�B^��;"\ ͒� D�I��]�S*�w9V�� ��V��;��y.���Y��X"�^<V�M�&�/���)���+E�eA��c�Ȣ(��E�V
�E
�mQQ|�fR��1�\T�m�E��:eDMZ�(VVV-k\����TQ����UAK���h�0APDb�+���B������1Ī�-��*��QEbԨ��I�Rڈ"(�4A�*-)k�3-��QU@�TQb���w,�VTZ�cm[�.Z�E-!kT"V��lm��T1��`��r�-5jDfZň�R֕��+(�*�
"�Q-�h���0D[B�.�Aq��IE�\J-j�A�b[*CHQt��Qh�,dQU��i*�����A�"(,r�X�J�R��EPJ%[hۍ�*D-m��նҶZ����K�ȸZLk�QB�X���m�-(�FV�b�[R�5�Yr�����]ؤ�y�5�ٯ$'>ޙ��0�x��G2��ǜo���ߺj���,�bM��U֎Rڬ�S,L�@��y]�l?3����	�<�ȵ\]�˸�^�]s�oh�+�lm����Wqpo����
�v�8j�F�-E�E�u~/R���WVzw��G/ZW&�����y-5�� �ݷ����OL42��z`����KϺ@�X:ɕ���	��O�r�$n"(9�m�b+u���f5E�K�P�޸g�U�l9�5ʧ�����{G6�va�*c;c����t�޶u2�����Mn$�k���S�5�c�賔]�̚|Ȏbk{��^c�x���ر�X>m��NJ��5\������Rb�n��ڙ�J�ςS��M.g��f��a���\�{w*SQuF�s��/t���+t'0��uuo,g��X�;�kv�]�K�[{��]x�����1<V
Q��VUlpi����L�^R�89�(JY/��4lN��m(�meRU��Z��EMq3�,��;���pc>�]HS�Y�P�0��s�fP+����9ը*zXk"�ڻ��u ԭ���р�ъg/rNS�暏��i�7�e����<�-��]�=e�ei	��|rw�3b���J2[�� �ѹ��n�_b޹Z���K|��l�\�cS�4������eX�r9�foY��eȎ�����}JH�[y�M^�QM>5����x�N��U�J�&��d[�aл�j�,���N��Yis��K����nBM�-{��ط���C��8h���	F��97ֺ�o�z�`��������w�\��J>�i�&7�J�}�=�����8�����l�{��[j�����W)@��w��!�"�y-���Պ�v�U��W��bN�G>�i]Y|���l���	AD��+GbR��B�Kmmc��ȍ�(aN�7yX�wT:�M-Xv!؎S1����zQ7V�gn��y�֜�Cr���{mXކ]�qK�'SA41��^�H谯g�QX����`;���� W��Sԍ��J�irN�͍L�M�R��Vk�ŋ�T�t��֒9t��Y\J#����;�������u���DHnԜ����إܒ�*�b��%n�M`C�]7x�J4�knh[����WaU�8wv�]�سy�cdG!11�9�mQ�R�:^T3ˍV��r}y֍�j-߹�cfN������5R����xnX6�Q�q�>�hhuC�*�ܜ۵�3]�kX�U�1J�v��[��n^V�Ǝ��'����ӘU��FEȹΥٌ����clvw0��­5�>+���k�/�W�g[��d�W��^����2y0߾řU%p�v�x˶{[՚��Ҽ��c{'W��Մ�Ĳ���q|(?��y(]S�(%{4�n��)�9٭ќ�˼Tf��nȲ�����C�c���]���M�4ݍ`�˓�٦0�S�'��^�d���j���o���Jc���J�7��S}I��m��e�q[Jʪ/9%|��48�8���s�*�c���0v�RW��A=Q^nr��\/m�Yv��	kQ��}rBU(f��J	ek��k�p��q�B�3�V�Q�}�ع]�������|ifg�j'2^+�lZ�.��.X.�����&�{�m"�"��	귮>��O����JS�ܶTb=�9�ڠ0�i̨LJ��Τ��I����aZҞ����t��R�%'t���_1��ןj���ʩ�*^/�����'�T�Af�XY�^�w[Z�k���^3T�KD�����J�(vuy��6!���G�H�%�]]��� ?�:7�H��:|q#_;��ޮv�ѧ�����(L�t�w;�!1b+�\	��D���6?xξ�,C�e�yj��k�U	�9�45�׸(��iⓙ�ܥ�F�\�n�Z�mr�����s�a�����j�u4U�zj۷������x���Z��2������4������<�ևXE�~������>w�:yU�P׬��is#4�;s�bɭ/Oazri��T�]�)�9�/-���Wl�x1��M`,§'<i�����x˶{r�AݙML�a�5��E��9T�y�+�)F:sr�K�(.�M�Y��v'�'h]՝��]�������?=����7�.� Drt5&�ƀ_o���j����=H�����Y�O^�v$�T�m�^�:��owzEW�JB��Ze��V�er�J	�:�1�:��[z���i���sިMJ�9o�� N�R��,�geu�b?m��s�'�-I�_f�!�1��ֱ=��:�kw"�唾�q�Z�[�vRQB��͜�l��ê��uy������ 7>n�� s;)�{݁��9_B�`Z��oz�K�� ���._��3���rB��_�cC��FL�� [~��w\��w�j��\��,�^ܽ��c�]��'��Cs��I�9�e��@��;�;�S��]�T��,)��3ꠣ�w����ϭ����K8��
v<�-b�zkE	�w�c��{۱��G�����3��q$yIuB�AuCfֽ0��t[�.0�Uf�]C��+Cn?yV��jz�V���( P��)'Wh'Y(X�1�=.A$��}�����K������xw;���@ (��������<�wfTM��^��)�o�ի�)�U0Ψ�y;�>�\��:�'��>P'�0����r�Twj׎���G'65�QӘ��į#�Ƨa���I���R��\���5�h#�]ո��Y%�C��$���&M������ul�E��Y��#�"F�w�w4+�l,���s<WNXb�}\WL��Y}2ک�K�Ѹ��YN}؏b��[��L&��X�t.�mD�i^�	��\���ʳΛ�.K���4��V,]g�样j�����mϹ�C�qPC�L��ڛܪ�a=�N�����]\��W��0�`���꽑���c6K�v���; lL�|o��X������ϋ��i�4����h�ex`���� t2Pm߬g���[�V��sV�v����y.��������g6L�U��CtM@4�X�]�C�{�ժ}ޜ�[���6�e��LB����r�SA�̈́�U��U��/j�^�gD�^�ա�ekŕ��B�Ge
"��&i�i�[�Br�gX��H�R�4�f���ȇ �U���Rbg�F�����оp��!G�/��W)=�����8s���Kh'ՃݞoۻL![��b���	Þ�A
�z&��_ew�~���z���#���\�\�4���M��_��:�I��:���(��]΋���/��bF�[+���7��K��r������lY��^�С�.;M�26��Քp)@=M2�xV)������=�ad��:�ݾ�+�ܥ��<�*��3R���}0��Ϭ��՚�lk�M�N�}��\�U���ʎlf��?+�`��ލ��T�E��s�;���X/($Eg��
��u��8Yݛ�w��>�T�7�+��z���}]�}�3�+<��&dH(Y�<��qQa����H��w���."�5ƪ��Ӟ�J�3���ܟ_�'M��H��(�-���2��C#���˳w��A�L;B���x���
��B�Ցz5�m�:��>�g��`�;5wz̼�㻭�yKaȚ��.hd+��Y�{�s�D�s�$\[���9�Գ�h-n�:D��:�6�1�X"�D��7��Ȩ5\��ݜ5��}y�����K���]hvb�a�s���W��ۗ�gȺ���>4�}�����K1w,�@�71^�Q��әN)ѧq��o�4��IR5MB
umt�b�Y������ �z�{�ZCn��%����d��ݛ/�u�2�3�Ҙ��GC��>):�Z9
����e]k���\n�����%SdI����!�Z�=�Q��C��E�q�E>�������^ȡ��3U�ֳ���[�p�_0<�A�+��p�p�UyB��E��&\[����i��!�}�;u���0�L�y��
�f_���4�z����ںK(�_-F+&�����Ig��Fz�UՃ!U�G��\�5.K�fl�#�y���^-���rujl����^E�Tv1l�]x����X�^t�V�;���mL�I֦�#�\����y�xkB�U�A�(>�"X�9p�o��<���:��Muu~WW��;r��.�J���yF�S"�ԟ�x�l>�u�ˏ���q���N�ϟ���C��K����T�I���s��:�uL\I�n=K�=!�O�ʧ�w�����Пc�5>�nH��*�����]Ŵ�+�4N�q!��M�~J�J��C�.c�\��W�%�b�ݼ���8&p��_��!���B-�*}cL��ѝ��X�2�� �:�d���Wg<����P@�."��<x��Za��%�^Z+6+�د��7Sa������������'�#�d���O�hr$O�Ɖ�?h>�|lz��c��;�[�W�*�V��l�y��AU(p:�Z�@��������ɂ�LZ�+}]�ʷ�@�-ٯ��s��o�z�_f�5�>$�,�r`#�M��hP�<����^!�n`��Ry��Y���"ԛ����c�v�=9��Ĕh�r�x..:�~�`�z;1L���O��Wb�?T��Z O9t�{=���2g����^�7jj��t���y�j9�r�r{��<��X�62d��ৎB+��m�.u��F1�,�(e^�M���CVR��eq"�$���i���w�=Ngw���C~.^)چ8?hLjo~e8k�Z}뾈����aq�c�,��tw��<h�g�d;b�	98�3ѹ�O��Z-	{�,DL㪍�T�N�&z�ޏ]���
5of+��w�yh	��+��4��ɣ��^Q�X%����O��q��o \<\@d<.-˧�iU���W�Kzsx]������^��ʕ�J�Q,\k���e[|�����u+�����F���][��>vV��u�zw�՚�X<�'A}�hbF5ܮ�О̬�b:�+o)�4�6��{d����dA�+�$6�;�{^kpG�:C�@l,f���{O�_���^�h�����T߽�V��ΐ\�b�]��[Z9��K��|�F2���e�J�&��F�����⏹B��ܽ��r�G]����!Va����%�wId�O/=�/x+��:�a���q��%J=Gyی�}n��K/��uZ��t�z~��ü�MG��b`���+P�W��I�&
�^����k��1�l�p��piaeYO2��9�M����n�����r��<ȳ��}���C7�5eM��{�(It�)W���P���_Jyt���=�,�[:t&9#t�Be��enc��qU+g�����"�����Hl+������fSF���]�e�����S���o��v����٬V/�⁀���GWhF�����	�w*���9�R����>��AE��8PO���v6tD�p���M�/E�;8ϡ�^�����-��xce���G6��{�L�~��_bw�2�C��R|9Q�3��U�Ś����Db���,	~��{/�尗2+F%y65;,s�2��U<�#`_����
L����'5�D*c�&�å1v
vr�b����/ʾ__�����g�.�oO����v�S���}ئ5|�����U�=�߲+ۘ�c6K�v���+mY������=5���5ٌ����c6Wm2��}�rư��x����k*i7j�ٍ��o�����U��;0�)�x�k���Q�T��ǨD4��P{ԑj�w5v���}��W*����0ߣ˳�]}s<gk|w��%����Zxd~q�>����Z�"{!^ab~C�;[����G��W��N�r��u�cc<9#�KG���Y�*�����7�>pˤ�u�Ԕ/]|T�xs.�*lc�-9W��e#�V7�������G�rk|79�}3v<��r���"�_�Y|_Q�8�2Kv��;�}� ���E�cb�	Y���ؔ�]}����tu��צѺī,��72a��P�:,��°����in!�.YzS���`��m2̻9��qR���Tջ9h�/������*��;�vn��8�u��#��hi6)�:���0ej�v%�N�4�`��x�1�S���f�9J-Q�v�I�\�D�j��k�Jn.,�-ӱw��%y�j�2� B��w��{�ڼ�g(9]���ʝ.���԰"��Ô �[�+xru��q�}�۹G��[��O�̾�Բ�:�w:���[�����r-�}����c*�gkr	Wʤ����B��/��(�f�^�5����P�#���k1.L9����ҙS���u�
Z�\\]��8-�'�k7�5�_v�4�v�r���(�łe��L&��$p ��_L뤻;[Aǔ�N�v>����u@ܬ��m+9-�����"K!��L�<7����2�QPf����Pܨ�ʔ�:�mm�Y�yI���dΊ��N�7�� ��ޢM�n�v�H��GY�E��]���J$2*��b�,�ti�j�˧�����*�c)��K9��\v�%`)�TAZĬ	��"����ҍS�y���e&0���; �ʸ��z�[�k��݇V8���M�%Hh��Ӣ-�r�\ia��Pu-�w�Fd�Q��J��p��ˍE{���f�)��AWjg(�|{����tM�m�\4�cv[�|;��/��X�gVpR��:�5�e��9j��۵������\wo*���=[�3z��fw�%ɞ�ŕD�)�%�V�����Sf�^ w�a<./$���k�= �e7�SKj�r���Z�KC�Y��͎ L���x�YxS�3���c�*�Z�}gk2T�u���"��]����&��~�R��R]� �yY7�$�Uѓjݽ�M�����j�<�������Hr��b
�9�&_ܲY���ݎ����$����&.�A���E��{7����x$�ūJ�<Y��]\8]N�^�޼��+{��Q�;G�|1G�뵴ลQ1G˸Q�<�w4P��N���P���k2����&}^Cs�؁�\�+	OA<{aW}]��sz�{����/+��(��AVP�bѩ�'Y�m\"�T�Ki�7[x 2]@�vi��fr�-�<^N�3���y����ӛ�!�d��9*���X�tC#�͔�#�c7|ܽ�륑��9krU���D�~�x��aDɽ7�i�4
gk)��ݝwC^3�����fof.i�NuV��tP����[�W*iI2�dK����N��Ⱥҙ�u3p��Ko9L�ڀ����&����fn�G��ʤz�GK�������t��6OH ��DQh�W�˘�:��sG��QV��cb�89iեaT�m�E��Ku�X���ӈ��Z$mcX��m�[+5j�iE+iX"��֖
�ڢ�p��)T*5[+e��2%Z,+���
V��LJ�ՋTW([l��bE"���\�Z��[I��1�2�U��R��"�Z�X6�)V��memYEd�k�ZӚ�)j���9E�XPkDm-�-*�W�SZV���е�X��Z؍R�+S,�*�:�5]�,m*�"1EQ,�J����\p�.+��)��,E@���-t܋rؘ�K�XUf��a��m-b֣Z�sm*"��ښpUe)ejR�
@�6�߼U���v̰�7�B'�ii,�y�{"���/x?(��QkxqnW/��iŮ��_fރ�x�s׶�n��p��u)K�p��8��¼�5#~�bk%���L�X��;q�
̻q�輼�������x��6���y��Prۦ w+J7��>�NO��eyz"%H�n/orY������܇މ+G�Ԍ��)U��gF5y^�^I��ָ��sΜ
)�|�Նʅr�f8�쪿)PjA�yGzu��!+$��_kUyvԲ�9�ߩƢ��V9]��Uu}�>�^�i�,8p0���W$/�Wb��8	�~����b9�T���r�@��v)�C��n��{�B�`Ψ�dv]��>sׯ��SD���.�gS���`��!�Tq�����L�s`SYp�s�d�2)h��ȳV�=�(e:���ܥ|@��ŝ��\9��z���.*=�n��=��$�#¯�a���l�MP�~K)_��Aa���Υ�d��x���Ǔ�6^Ŝ<�0�)�����:��y�G1T ~!����R�����r���"Vftd�B�n����>iwm�����؝��QbЖ*h�������:�]bܼ�Ҵ�s�:%��͕�t일�TrtNl��d� :�"s�����/oz�a�B��vX׊�8�}g��!;�ɢrp�>�u��{ȹ�ǎC��܋�a�9ψb�8�����6>ٚ=W3X%A>)���A�[���0h�{�u�"5��ۄfmT8t�Gp��"�}:hr�"b���R�����Y}����[�=UgC�k���p6�X`d��uS��]����^���]�������MA�±��1>T�.^�D�p������r�ɗ�#&�PW���1s>�#2������=���A�xkB�T�O�H�7�\:��9�u�Gq������g��g�����q��^E�F�S"�jL��.s��"�W���P\��|�.n#�j���Z����궩��B��^Dc���Z�:q�ix����!�V7A��V^#���λ�!��"O��t�*xɊ��2��THg ��5�Z/�Wz�:w��i-���@����p%���8�{��F�r�S���Q:ٕ��T�F��P�o&1���|Hb�tWL�4P�M����Za��%�^�$Vn���ﳼC�O��Ҙ��f���23�lA�i��T����J�� ���-����C�P����9����8�]:��״�N�Κ��׻�q�jc��D=ä������[��ak'*K[��E͋�������Qg-=ZFc]���D��Y�t}�J�f�������C�"}�4H�c��>�|o��4�����G��9���>�&��y��m�Õ�B�Ѣ0�."��7��7��	YM��l��x�R˽��Pc]�=�L�"e0��T-�f	W��|6�o���ax�yL�[(N=�Օ['{H7�
�����9���]�ٜ���,�=�������q2m��I�k�=���B#
~{���y�}���a�7�v��s�X��p�>��'���ȡ]i�7���gsa
T0W�ȳ��W[V;s:V͞�]��,C�v����$��q�o*c��TS�O�t�W�F�"��2(`�䊑�U�r	����o \<�5��f+�n9!�|�N��g�,��>.CP�&j�Ĵr~Qx<|o�U|̡m��I�'}�ާ���Ė�XSo��oY�t����c�6s�����O��

*T�3=9���h��o���{��kh�\��H-�sg Xedu��^#��r�]j�5��x���)<�m��u��;�	���G�݊���G���fn�&��L몿�垞.�٘uZ�K���Ng���H�6�=Z�m,ܱ�W2JBв�Jw�u֋���"�ã��Kf�m	���iΝ�����k4#)ɷ��۷qiH	��0������Qq�S��P+��
�J�s��dJV7Sd%�������G�+����.�(��,תW�{U����ZK�-,�2ۗ��xKG�=��*����.��"��=f�3ꠣ�����>��W���b�ߪB�2� 4k���z����a�;���j�NYf ��`$yH�Ƈ��١2_XG�}�:"��y�\)���U��l����� @�c~R*\h4�S4ڪ]�~#]L��.�g;Ӡ��C�Q=etZ�
+�m��瀣��
�?���1��oޫl��ƹV#��D�d�1�^�^�v�N�^V=�{��꠸�k����j��
T�yO,MW��;}����+Ԉ��9�ٯ��U�W��`jvX�L�l�O'LF�̉�V�*\\�U��N���
��r�=K8�ņ�b�gd���ǋ��˝l1������ޮ-��}9�fm�C�@��U{5`ux����!�����u_acْ�sʹq�I���f��;�� /B��,��r�� Bu�"��$j��gz 9q\e���o ����4K5e$~����Emi�̈�,�D���a���IJ��Z��e>7���Fr��#�o�m�w��������e���̜�R|Gf D��e���NN���5�V׻�	��l�/���S'(}2���Z6)���ZNМ�N �-�)�e��|�w�"Xr��0�������!������P��וc�LT�f���/�g�����~����F�
y�.�U�p)��fŧ�ltg�Pٞ����C�K��w��|�ǫ�4�?}x�1��P�u�bG��V<�r�����NA��lt��Տd�8�a[ٜ���x�<>Xk�#�����"���C%���$_)c�(\k��<��eQăe&��_��=k��̗A�K������\�(н�������r�꣼rh�I��S�N�A�>��G_�w^`r�u�<��#��\��Ae�/�~|������CK|��OD�Z�$w9�-���.:���]U���lu���/���e	�b�x�u�xj�r*,��#���@L�J�prj
U")	PI�v.��_��3�@'��f��uʃ�б��2%��]��P.���w�gr}a�pT�]%�%ȧeC#�oWI]��P�CAoor�}Ǌ��w8g_٣���@�Y��މ�}���C�j^룛#�e]�y��7����åN�'�F���J63(s�P*��6*�3i�����t��j`���;:�b�FV�����2�cm�HЯQ�v2���K�~�.��#a���p/UK����W<Cpk���;8�;0�X��&_���La���qf�}����n7��X2|zI~M>�_p�y������`�����<���B%G��ݏY�
��y�%�5��T��L�]��<tl�����^'~|i�9���'1w,�%T!	j���W��o}���c#zmHݚ��ψb����\x)�s�	ZY2���s��~�]	3���{���f
X���-������[��B}��&V� ���D�1s9������gu�Ϋ��B����_<r�g��;�o�����{�9ۻ������&�lm)<��J�|Eb���g��	�@<u˲�����p�:����.P�T���{h�gc[������W��߈��58��r��r��f�H��9p�Ր-Yk'�vͮ�i-�]?9�7c]�Z��h���X�F�S"K�"���Gn�@GfbW�9�D5�<+i�\���pt�M�v�R�n��m����Ine�mZ!Z5�Sv2^��m����y��Z���eg.�溥){��<��E��d�v1�39.D
Q�W�ϒӋ�c�Rܲ֜g�*��3��)K<��]:Z%vr�^��*��gU�MD�
�^Dgm���Z�ӎ;	x������^t1�MU:����jD�L��H�#���/]Ŵ���BpP���zm��*5+�e2��\�Hx����b�gӱ�B�o\*��ob�|��{����'[2�j��/b��)�·����c]� �x>:H�\D���q��s%�ʩˏ�2+�g׭rX��3���L�%j��]�F��A���R,Dg�O���Y�^Li�C6�=���Ź�q�!����<�C\(��z�O�&}T+��*�n���Z�k^s�10��)NPc]��'W`,�r`"�Κ�4(S��iY=j';���'��ʝ��M�7���i�ꯢܡC�u	�/�3t�>^,x��>���'Ϝ��͠�!�8yN͒n�m��a@7�v��}a�\8Q�˛�U�n�9w��b�{�u�lYdt
�P�YJz��yX��n���,C�Ӱ�V��C4�KLb�|�y#�'ow^	8j
s;�2�}�͚1��a�{�仺�$*�hKmpړgtt�Xە��w��v�_q���.2ճ���*GLPe�P�}����N�4ܝ�n�H�tfT�K��y�/�qԁdL�ؒ�ӓ�"�B�+7�P��,O���Z5a�V�\dp�@�f#gS\���u�t��q�Ip���[��=�{ӽ"�j�Ę9�?(�<|o��yuy�������^��f��̡Ӻ��W���>����Pg�1 ڿ��Y]y����u��n���ׁL�K�C�v�P6�m�u��9�EŇT;%FyWW�ش�}W�Ì���*��܂����S|Ӧ`���jǵ�\F}�W)`p"Սv+d��3[ԣw׶�efE�5�v,�
���h^>8�]0G
�sǂl����r���H����$���:y[Hg	������k#g�a=SP�B�/�n>w�pv�/��E���+�s[��t������#��B�C~0�O)6�W�ມ��'\I�99x���'=|M�0W@�C��-U���'o�v��}��B��"51��	י\�2���4vV�"6X3h]�}�!�+OyM�!����>�ý�U��]W}�=aQ�ԃ���FGd�/+�vV�L�r��x�q�(�3j�1�Jh�3f*4.�y�2E�˓ٶQ��l�B`�wL7�9\S�>Hj��Z{{9�[]93��:}���¾�(����6)Ģ��N�o,�>5k��d'z�+Y��U�*<e����T���JM<�)��@Y�fZZ/�Qy��׶���S ����_`N�L�B���:�y��B���ø��=��׎�} Hَ���S;�݊��^G��S���:�/[5S��J�복�75���.���XoC����>hv.��;9@,Ģ�����x9s�nҮ��y1��gm��s��^Oz����נ��X�>���������sa�fK��|�Qَ��Ӥ���*�X�i��H�X{}{������h�e`�䊜�R{�O�m6�V�ޞ�|t2R�X�%+��1薛��{j_��!7�Lm�X@��O~���jK�zyR^ �]f�-�/c:��o���˹B��x؝��^�L	o�����=��ex@����'�Һ������b�~u�Xhi�7q���{��|�gW����<upK��E=矲l*l{�V�3��_6|��c��__8En15������"�JO:�o$@��z*T�[/��{:ׇ��A:��C������ҍޠ�9����P��:��u1Z[��f���	���Z�P;V����kJ�F���WYm��ug�==�Yd�F�ZI�;��9ǃ'.�e��2�;�l<GDrgYy/�����8�դfn���v�� ��݄���������c_#UPs�;�]N���_xz[��]�淰j��3�^z\D�1������y!�C�=gU5��\]��7���^Np��MQs�Y��j^ggރ'������$m�lK8�h��}�~/$��O�"�[�x�$Gc$��U�7���r*��Ў[�q�grT8���J�Bx��.o�I��[(x,�����h�Ϊ=ʁz�z_O9P ]�;�{Z�)hk���oTnx�j�z�e
�"���]B���7ex�!�uѩ��>�\orz(��̸M���aJ����(�_G�Z�Axs�C�0�>K��/�-B���(��{iec�M���5�Q_���\�+`��[Κ/���R�/�E��JJ��o�I}��ns�.�>`Zf���ۗ��C�Jfr�������ƚ��<��������/	������=��8=�]g%��6�n�Cu���o,�ml���	
~�c�.
�޲��ׯ|)m���c�k`�
�9�iB}�p?���}��Z����VQ�y�9]���?cVz�+�儁����n��>�������,���6��Vٮ�g^`T2�3,X��Ʒ���P�
��ĵ��٪j��E��4���hk�#�߂�"er(+v�z�0~������g!\�Ud�-(���N��i�oUj���C���6ʹ�&`=N�f0lʨ�5��q����k�o�n���n�vl ��7
��e
��i�:���hr�u��,�ȢC[Օ"������ˉa��ٕz��ꛔů>��QDz����^��e�-,���MQY1�޼P5��]��㣤�lRu���5�Mt�0��d� 3��=�Um���7�턫��ރ'@o#��X��l��lu���@�G*ѡ���"�f����&Axf��� kt
������p�Ӧ���=�f�=���z�e9�F�jd�ȫE��}/�f��u��~��MpuBo`��� q�E!�5f��v�YWb��Eu��p;�S׭�'�vjď.���x໊�j��Ǉ1�c��;L�@fH�W)�y��bu 3z�ӿ17B��1C��1��5��5Mu�����G�^��w�ʰ7�MɔoM5Ռ����X���)Vj.�,�;�b[j�\�MS��y[�D=�C�v+[8� �<S��*7KSH?��s[�#�w0*�,�K�^D(�(���tV�BpR���{B�\�\��n:s�;�Յ[�o�D��5�B��k}	 Т�g��=E��em�Ъ��6�u���꼊��P�$��x�g5ϡ�vQ�7i�|�����wP�k2�[��ם�-'K4�)���r�bל踩��!�W:� �DE�xv�)��ݮW�v�|���写�U��wp�^��׹�ZDV뢒�M͟nwv�b�.ȻH+�b�����q�=	�%lk�C]HΔs$�6I���8��v����Y)��<J+�R߲[G'k ��b�������=�TK/��5Ɔ��lXp�|��kB�}&Nm���i�_����u��nu����gb�bH�N�4_�^4$��-�����e��q6o���Ɲ�.�ʙp��o:�$S�;X�"�x��R������ry3�i[4��uFzd@<W�F_�f�</�z�:꘢��9F�r�,��`<��x��R]��ՃA!8���Þ�ǹ &�bF��O1-�Y�؏ ��xmVXO���%���܆�����^�5��b�QV�c�u!M�dC:���r�0�a��-$��8�rV)�Ҷ��?����+�.�n��=�[�KF}�4{/Q8�:��s3RY��]	��Л@���ц��i��XW�����N�#B���3+e�P��N�cWoVX�=li�����q� �n��p�2�˯kn8��S`�G�mŘ�n!n�Ǫ�۝��X�%�����X��(g�����l��:ӆ����Û�e:(�I϶\ԶȆ��ncɆQ��rI����J����"�(�J1l���j��5�Ƙ�Ej"���k+Ѻ�L*R�j�&Z*b�j���[m)J����90R�TkZ��6Ե�E
��j��Y�U:L�KiQ��-)k�ڭ����T�*���K��iF�R��hUKlmlm��3e2�֭�c,Z2�Q,V�)m�\�1Km*U-�J)h�Qml��"���ƍ��-�a�l���X镩fJ�V�c�hնU�k[,��jƴ�V������p��Q[E[V�E�-�����q���-(��e(�bT�Z�aU��lDm�h�ձV��1q�Դ�T�P��j1m��KJ2�RZ5[]a�h�h�E*"���c�YkE�TJ�KJ��hڍ�""�,eYc
5+Fڶ��Q+Z��#����ڪ%U�+KjR���kR��m���q�������KܕnC�.�.K�M{�7�,��9��(tD���҂lն�3|���Lwֆu�J��[ٔ0�?����̔�Z)���/?�}r����eA��V�3l���Bnj,C�8�o�Ve�)�����W6g6���E�ӕ\ja��t���\M��즰s����R��e�YW�M�[�#��|��ޜcx��"���u�{��K+�1�
�SA�)�ie�']9\����g��%�{h���y��q�8��VkȰ��dC�x��0���Y���K��'��x/D/�_U�������I�RY�y���!���~ɯ,�'ua�?s3H%Hr��jɈ
)�}�p>|q�R|��i8�㝤9��>a_Y5�i�e�����擾��s���u��˭���������t��(��YP�%��݁�T+<�I�����aQ`}�٧�8��6�>����ì1�j�8�3�٧��L@^�{�C��V'��|1���ﰜ��Gsy[`q������q�w�G)8�g75�UI�+��Y�g\a�_d5�B��o��h���bA}?f0�bB���$��O��q7��x�~�T�߿o��=y�o�w���}���c@�+ӿd>Cl�VLCô1a\VQt��V��-N8��6j�Lz�Qgb��������/ﷹ>e�!Y������ğ�y��>�ϫ�Tkc���槽��qP=�'�zF���>k�|B��w�6�a�1*�N��1XqƲTR]�QI��8�!�Re��'ua��ݚ@�R�u��J���s��y�'��;���_A�j�}�dQ�&<>�L `�'�}@�}�6Ì+�O{Mm�q��O�w!��PR/Xy{���+*�ϩ�R�*��Xq4�Y�����u�E%B������o~}�o�}1��*;�6Wo)��`�ä�6�D8o�t�p(&g;���5�\6�'��;okv(���*U�u��Z��\�p���s�QΔž���1y�٠�̯C��n)��SfeV���(V�])r��9Eo��8�Gͺi�����:��V�s���.~�����<�|�m��1?�̟�TJ����o��Ld��*(q%w����D�+6���C��6ì+��8����a�s *�1��:��M�N3Qa��+u�����ϻ�tw��K^`�#��P* l8�����1�'��<��u��>���x�a�|���I�+=��^�*,4½Vnw�|I�+&�w&�E��:��1�4����l����Q���w~D��8 D�C�X��0*M���ud���B�P�wI��c=�1����O~�H��ǿ��/�w��&�l;�J���'��Vy��^�TX�n�vUɴ��}��]����Q�A�}�k�>d֬<��T�d����J��֕���+?j�P�z�㜰�va�
���߹�Ă�̕������QAH�'�}�m'U��|�����sZkqeٿ�����<&<6"=���\yG�LH+��g�i�0���s�O�~a��6�}f���*,�
��T���u�c*(x���'ٴ��Y�M�7�;�
��
�{��/�����'t��T�䷾��<�	�d{��`
�>N��6��Rxθ��0>a��
���xΧ�?3�ğ���0��������_Rc15>��CI��,�q�2h��4��Vy�'|�߷}K���������z��+��浩8�O�V{���E��0�����h%z�Q��d����>M�`T��p?n��/�9M0���|������&8��J�A}a�}��{��ߴ����3|�����b��
�W�&0�������Agϓ���6����ȺgRc�C�ٽwgY;�{�ru��=J�û�svu��y�kB�2z����U�����\_yME�k%�k�u�5�~�����zÌ+�;7G�6�Y��&5��E"��d$겠���HVw�`i�a����L�C��>�v�Xbq�O���,8�~�OgT'��y~�k�Ѹ�+�K�I? �za@���=�ׁ�z���a������Q��!X~a]���uI�+9ἓH
�M�<`T�����8�ꐯ�}��8�0��LC�}�&���!�P��*��Pc_�M�Zs�*TU��G�im"Cy�=���;��QT]({/۞ �����;iv���O�m!W�|P�����<u�n�	�y���$ѽR�p2H�dbPQ����X� y$�-�]n��[-�N7H96AV���R���;rʛ���3�����"��{��Y���# O���LCi����g��ùgSI<B�]��
�ﵕY?8��+7�&r�'a���ii^�oZ�g*Ato�ړ���g>��z~���N��f֙���ޘ:}���ﳸa�e'ɷ��H,�N��l=B��w��>|`��d�,�P6��\���'
z}UI����Τǌ8�nͤ���O~uy�=+j�u��]������s��(�=��d�=`q�O̚t�o�I�O��(~��8ϡ��L�2'%VO����C�"#�Q��e��Ѳp�!S��}�o��]�ef!���٭a�x�A�`u�,<���6�8 ~�LC��~d�wD4�W�S;d�8�f���p>��!X|�{�6��I�&,L��ޘ� Aֶ^(��F/o䷳;z(i��Rgf�.�z��`oWL+:���:���c+&!���&��5�ߵ<C��1!��5u%bͧ���ISu
������<H,6��hL8���*��%��߁CF�����Y���Hy�Lq���0�Һa��Qg̕�Ʋq1��Ն��vOYyCٺM0�?e&���:�$i'��m'�T����̓���T<��MT�.G�� �d���G�4�$���Z����z�I��=֧U%0+<>̑t�c�7?^!���4�a��q�@�U`{l�%g��&'Y=q�&�i'�T��g���HVa_=�I�)�<"=�f뚐H�˼��Ϸ�������b;��4�`T�T�n��K�B����>T6��6��ý�i�3��!���H.����*C���E�aXh�z�RW���p<" ��ģ�WK~���
�/v�i�����t1ﺬ��W�<&<.;� uI�p�sl��X
��2Co�C���|퇬/�O��M��&0�6�9v�Y�LM��Ă���0�>�*=��b�/�_Ð�v��~<����_�Jş���@�*O�������� �����x��q'��X)�Y:㿽����<J�=9܆�g̕&�~���OS���m'�~�=q� 
��
����#Ff�^�%Gʬj�mv��=:��ͯ�ĥ��]��u�/���iīi��]��3��k�l�6�m{C0�GL& �Q��V�6���;��!�;�����7n5虌M���0�5�I�m-ʻsL��
90���c�EB��\� �]�V�I$���mל�߲��
|��z��򋤛J�CS38��/�T�T������w%I�b��a�qRW��<��h��I�S��d� �γþ`s��*�;���?[>d���\ehS�/Wۑ�lE�js�y��=ꊍ���4��1�s��a��]5�}��
l��ɧl��(xk0���㿽֦��K�C٘�:�Vu�S���4ͳ�c:��6�A|C�ub�u7�cj��}w3w�b T `
H=��ì<E��Vz}܇h|��N3��6���C5M7���=B��N�B������8��ߝ��8�P{�)8�t����0<g_v<'���w�����f��,zcã�0�;��Si�0�<�{惨TR���d8ʇ��1����k�%b�O����Rb�?�������+'\I��xH<���.�| b�Y%���ob)��en^�����3*�Cx��1�N���i=C�d�{��i
�l>�n{����>N��]��*,�w2/P=q��.a����J���5a��=0�ޝ�OѻY����!�Xz�u[�Lzk�C�m 回~��aR{�x�H}l�O�|͠(�Y>q�;�4��T�^�z�R���ɷ�OuM0<��q��d�QM��E�cº��w���Z����3�}�*	|�t5f�z�V~a��{�6Ρ���b)�_�jO�����a�l:�f�W]�|�C��o�wRx���ɾwo�lI�zgr�l��xLF�߇۟i�߰�VX���o} �� F����̕�UT�������>a{M c3�cu�'i�0�wF������k|�C��ϻd�Y+m4�}����@�LK���v��Z�+0���S�7d��`m��U�N!���CI(���.�q�@ǎ5���2T��(��:����&�T>�&�=ɮR����u:��S���R|�����ݵPJ�m�H�yY��w}��8�����6�{@�3�sP�%I��zgrM3�I\a���)�1��XqH9t~����q�Cz���C�gPPS�����{`x�k�ϸ�U|�z�)XJ��΋������3����;t��
�\a���&��g9n,����޼�X7��@�V��{<����9��U��|/L���y*��=q�ؓ��S�N'i���%��9�GaӴ �X�b)7���=�@�r{f��~jW����ޕ��8g_*[�޸JG���US+�M�d�~�M3+�Ne<��
E�Ms�VmR^�{;�0�P���M$i�C=9�a��I��OP��sT3va���~����>�yƸ���p�V}0 � ~I^ϳ�>d�7�h�|偉<}���l�܁��b°�F�S���f�+�4���+����M���L?gp�a�i1���Φ��k�F�]?X�2^u��_r��P
�r��'�b'�c����X�����@�*G��c7�& /'�٦a^�'\~��4�{E8wY��0����&�̕m'��3h
���N�K�7����Z�M�^��|�C2æ�9HVM�c�O��bCf�'䟜I�TY�&>�q�ך������w��'ɏ�d
ΪJ�7����]����p<x��1�i��{�ü�^�=uo�s>߾����_,���Xm�{��I�m!��;�&�R��0*OP�)Y5��
��Y�=d��f�1��+�L�Р�_���h�VT:�����2z���c�G�n�bC�[��os��Ǧ�8���|��q�E ����a�~C�1��#���4��@�*�_]5:Ɉ
)�h��\�1���i�d�w$�ݚa��@�l�����ǜ{�_v���|�Rϒ��'��8�x���i�8��w��}�+��Gy3������hz�E'{C�~f!��9�)���p�� z��B�]�bLK#£�a�G�w\('#x��v|o����� ��y�Z���8¡���6�z�QgP�~̚@Qz���?w�VI��y��8�����C�Rx�L@���L�'�$�T|9�1�f�F: ��=�>���%��������aM0Ϭ1*N=7v�Y򤮏9�i��k��<z�Hc'��dזq�����fiĩZ~�Y1E8Ϗ{���
�罳I�O�!��!�	��x�<��MTlY������ԩ��3l��;7c�()��2�N�*Iyw�L:�Vk�d8�H,�ny���aQ`oϳO�q�'�m}�^�u�"�s�����y��.
�z��
��۽�'�����(��v�lO�t�'�+��C3��~lo�pn��q�����\x_r[Ѽ΍����5����J,6��!����C��$=ƚ���[���wq�]3����w+9�h�s�ݕ2�.>�6`��1^��:�=�3��}H ��(lmw~��  x�l$�����@��V'��CL�&�쇅���VMU���d٭`
�N!^%dRc:���9HV����h���bAZm�S�p�rM?$�� 8�v�e�4�%o�3�2�l�ҝ���8��8���!�y�&!�(b,4¸�5�.�q
����'a�
���S�TY�ެ4���d�gp�X&�����'̼�+3T�xY/~����S�y���3gRqĞ%��ti � q��wO�T��;�������:�H,�a�]5���Z���M<a�1�-��;�'���J��߾�Ib|q�eJ�y��~�ǽ0 ��N�I�O���eCI�'�}@��a�a^�{�k��,�%v���E"�����O�Cg��)
�
���&�1���gXTRU�Vj>��_#��l�r���s? ��������A�0���d�
��P�o��&�'Y1�娡ĕ�lO��D�+6���y�l:°ٙ���M�Y�N�@URbG��n�7��_�(����#"�_����wyHV�tSL=g���1�a��?!Q|X���b����$�<=��E�'b�ܺI�+<���	Qa�:���|I�+';frDG��Q��x|w!�A܍�N�z{��gwy�~z%v�Qg|�I����i ��j~��'���+�j��wt�N�3��1����O~�H��=��x�H;�{̓��ya�S��� xD{��r�$u#P���]�9��3��d��5��|��0��>� ז~d֬XT%d��c�u��)��²z�Af���x��9a�0��zɰ���l� ��J��y'wE"�.��~��ט�}�>��$�'�ʇ������++<�6ΰ�1 �K���4�XTP󿰚a��LCN��i�Cq�@�*y���:Ɍ6j�ERWi75f�x�}�{�%�.��.���2�r�O1�1��g}��;���g�ϰ6����o�ᴂ�l㏓������*��:�a�?&$�}�<a�1!]�\H,��>E:�$(V,Y���?���1�؆���Y˾����\�efpf��Rgd���x�<��J/��M�Y�^�]व�Z\������\����ux^��Y����\�7�ge��8v�_ Ȁ�扐!U�-��YG�)w�"+�^v��C�[��%WunMF��ܖ�������3�^���I4�g��O���aSF��|�a���N8��{>�@�+�J����:ɴ��Xq6�R~9����~e�����l=a�Ri8���1�� ]��5�\
y�T{��z)�)&1k�
��������ɽa?&�8��0�z�Qd�ءԕ�!��ug9�vs�:�h�a�XsVu��}�kB�3��23�_(�W�\�,<����N�=�S��s�;>�i��+�5�?Si��oT�Y9�PR-`T�VT�_ԅa�~���&0>���3�ugXTS���aS���������8Tc�����U�k�g�T�\xL�w��Aԕ�8Ɍ�Xb(x����Xi'�+1�����B��»Փ�ꓨVs��@URo�1 ���3��|�ꐯ��m�&�u�LA;���8��U�T~������p* �����QH,�&��m�ă��톘�i����'Si=B�]��H
,+�XVO�$�
��Y3�Y8��7��ҽd�kX,�%@Qy��3��5������~�z�H,�>�hwvN2��;����Rq6�s��AgRu��fC�TR
;�����Y�P6��_P��*O�
h����TXk,1��q��{��s"��}��ө��~�@���l{�S���xJ�Y���'۳�����d�)�N8���'�T���n�y܁��W��s�~���g��X�Or��\H)*��Ȥ�R���?~��������y����q����N��eg�c?0���Xu�O7��m �`��CH��*��8i�W��&{�t�C�+�xgrJ��+:͚��{�+��{��?#i1
����o������߿{Η�s�}��t���*�t�1 ��<Ⱥa����]0��1�Y�by7@�VLCG��4�Adѿߵ6�S�bC�2䕋4������1'P���vs�Xm�y����x��}�������Ε<dۉ8��膽�Ɏ3��@�WL6eY�J���k'SXb�d�����
ùI�}��I�9�I�TR
}��']�^�P��xa}��<����͟�m𘈶��n�d������+��L ��q^'op��F�P��.9r��q3$�2_:�>�.�Xy��Ko݇WH!��J���b�SFq�N�A����v�*���sz�\0�x��`���6:�Kz�"ƫ[>�.ھ�d�(Y��1Q��=�x{�o/V�k}߇��La�S��m4�I����S����*,��*$�!���H;�L6}GvaP6��lm�d���'�$��I�*xɳ<�`c�b3?�L ���|ܬ��=�,��޷'����o���(,����AI�M��m$��*o���~a���CL��i'�H���C�bA՛�Qa�Y���g�PlL}���q��O��+sn��i3]�V��=I^��sP6��+<=�ړ��!Xm���hF�u�;�g�J����2Ch=�_���y�����4nܧC�k��f�[�s}�q��ʈ@^جb�B��G��M�!���va�I�����������Ҭ��M���L����C�uD0�"�5t��ϕ���<lF8��|Eu���z͸#�5���c����Ç����Y����j1Oι~��:㤘�y��9]�UdL���LMw�Ϗ�9]@�ҷ�������6k�|i��j��7�?,�1�{�x�y�W�-��P�"T��jӾ?W-7�߈^����C��.�%��=�	�����5w]�q/���(�<�L0/�':�J\D'���ٸ��A\���YV���^d�9O�wv�(���.���_���ɕ�ة_v��ᇢGt}�[��P�CҒw�����l+����s-��VR� ��yM�����k]E��`�&��	�WvCNG+-���L)�q�r�Jl��
���I�V���׶�v��}���GS��V��Ւ)��/�\�B�qٳ9`N���B�Y*鞙�`�TFh[�n�I��(q�y�������ï�ל��Tt��� � S�Q�<� �X�TY|z�w�)��tedSɽ��[�{��{v:;i����_���ē��|)�%ъ���{˷�"߻q[X��� ��u�B���ݣ+���8S�2D,�Ɇ���zn��܆y�]Or�&�u�]c��Gj�};R��T�ы�<P�↳^��O���*��{�z鳭yfz)�e��ǭA���`�N@К��sX"��2N��:��e��b��{�y���������C���5���]�0O�t�]w�����R��G\��˵�rf���n�����4��U�VC�/�{�D�ns�ŇN&)址_t�L��'<�'wywO�˹34��'�))�ݓ=R��(y�m�t�dv$��-�&��}[���l�g�r��Gr�5���H(]�9Q����Xg`��`_R�v��lt����d�=xsIO,	͐]���<[G6\r+E�D׶�ϫ�E�r����U�\A�8`�Ŭعݦ��/N����t��v���6˷��a��^��u��@�嚢�NZ�`<�l[�j�?�
��r����Ԥ��5eљ�K��Lu�m=�L�:�^�j�(�^V����R�!��[������K��	W���o����}��/&W\��|�tt}�^Pq�r���S��6����V���!�Xo�TA��gqi�JY�cWd��&-�Ҡ;�j0�\�����qN��f��>��E�����޼���U������9`QEj�GQU63�ӧ�j�E�又ݯy�A�ũ�ǯ��n�V�O�Dp<}_
p{�[��W׮jǣ�B���}�T=��E]2�/f�9I�~6o����^,oˌHl�Ɇ�Xҙ�
L�O-r�(�N�u�n���t�\8�(x���63����2��8_ڈ�M ��%7��\C�z��WE	�9=���╫�ϗ��:"����bʈ��h��FO�B�Ph����3~݌��j�`u�U�C�]>�ޠs���`�T<u��(&�X��I�@�+4e�{�HL�^ܵ~��B��k`Ŗ���{�ܰ�!��H�[�&\&P�ÚbѺdB�^̍�b�qb����U�],��|pQ.��v��-I�E�9��6��@�@��e-��/��Ŝ��P���%.�?���,1���������bmuu7F���u��K���zi�1���wA5��R.۩o��f��p7�˚��bN��V��ub�Ţ�|f�}v]��we`NH�E�a�V޳SR�;Hld��雤ɥI�xғ.�юH��Ul�aWq�vYIđ �Q�9�ˁNǓ�,����C�(���}wj�.����wn��FN�6��5{2�ɏ 5�[�ޣ3�ϙ2��t�V�c�y�XB�MT����_�{��t���SLއnTɁ�O<�{��Mn�! xR��Xk�zgT��̿zj[����}���pT�W.Lm��EJ�� �]y��p�Ǩ6���,oc����׈m�&Ꚓ�@VvԨ� w貯MOQj���f��������,Y4�����t�8��Xo�TL��pu���j�۩�C��c'_2*)�ю	�jP�V��mY�ӼNH1�n�s��ú���!s�az*Tf�k6n6�h�����]��a��鷻�o;jl�h��v�Ui=�E�ƛC+�3n�=9���y��u���T�WQ�R��[FU��>��t++TU}�M���b��v
�q`�ÔdXm���쏅ki�}�������w��x�`���/�.�[���r�6��@��#97ԛZU3��﷙���bv|��,fh:�ץyɸΑ��\��2Lp��Z��έL��\���|G}����f��5��APO�qQ����q/���os�vn�y�k�/�qn�V�ԥq���31������+z��^������Z��\Ȳ�5�Pv;�ݒ�h�.t5�
R�����W�_3���h�]��p}K+oȮ�֍���b��47�i,��fݼ�T�#��V�_:��u5���*�?,4o8\D������e��X�K)�è{�;g=���Z�^j_�5v��<�t��t+������FJ聃3�w�h}MG�k��mhP`,��Z����KjG��9�XeG��&)}��$8r���=�A8�&	���ھ���)�Ѫŉr�^��~c]��㮒N�/v��Y�W;lv)a���m?�費Xx(����:7�F�Z1^������W7{4�l39���_}�����̝�Y��ި�.�+������Vs�/-lO��[��W]��OP�[Y��1�ң[�:�9���@�b�GS�^4-v-�H�˻�LU����!㒈䭋YN��!Cpe8t1W���99��).�۴���&�]���>�gvWo;<B']`��
ؖԦ�ܔ�5 ;.�1u	��V�Ju����c,f̹��6�M�ݠ+z�,.�ASk��U�݈c���J��W٦VB�]p.�j�K�&:�)XN�9ګ{6U1\�r�����6�g�G�5w'f�E-�.���0�͹'�߽��B)B�0RE*6�kFT�Pr�d��)[T)F��ъ6U�V�Z���T\*[ZD�kU����J�Xc������m��Z�FTJ�*�ܵ\��2�mk-�J��KZ[KjQ(�cX�V�J6�n��J���Ŷ��Q�U�E���5l�-+kej�65�VQ�)(����m*�ʉJ�[U���cuqY���
�6ʥ����R��%KiKK�kEZ�SkUQh�)m-��ŊR��ʍm�
նU�-�m��UV�T��Ӏ��mm��KjʣKZ�aQ�e�IR�����Vѭ-�c[jҖ�m�[R�4�
�QU��[)QQj)
�ڎZ�A-�-hT�iD�[c�(�Z�RZбZ�k[d�1b�i�qmR�ԥ���(����F�-�R�D�F�Kj�E����`��U(�ո�(�U�Ʒ-C--iU[J��F���ETV�([J��ѭ)Z�
�"��*����Uܺq\ъ"��铯�i�3:��R��Y�b<GP� {7����uk�<ޤ�*Л�8�ozK��7������{��Sۏ3Sɜ{�1Qpuzhp�U�q�h����>���/
��縆���㬭��$���g�\U� �7�R�#�7`���qQ��nV�dv����}�K���+�K�tv#��*\��Z�t�;���}>��g�`)ֺ�/�X_]x����z�zn��wkok�.Y�e[�����p�. 2����|z-�w�::E��\���5`�N�u����FKu�j��g��Xʦ���8��;eX)�]��j�8xU�;ϕ�m�ܔ,�7�T�ؽ�u���,�jjk�o���"ǐp��[�	��/̢������XXOG=����bޕ�-)�1�@��x���zׇ��.#H�5
���vU�]ݼW�`���m��%F9�T2$���м|s��,ST`��r�ɤn�v�����8�s��h\�쪘��!��*-�Յ��Zϖ���"�L�MЉ��u�垎"�n>S��{\�F���Ppg>�p?�77�;��&3���\Q�ߗ�a��f�}0H�'X�/ZE���\`�h�e����k-��o�g�tƷ���ėh3�p����IR3�T��^c�M�����V�`������m��s/�S.R�']���������7�[H10P#`�)K�[�5�f��u����=�`p6�ܻȆ�]�� z9r���31�� �*Pc�t(�T��8��&흅~O�Πr|�@����{i��C��\�f+�{.����1C9�`�/Oj���7k����*�G::9�/Ǡ����V/�Q����8u#�D��_�ν��^��Vv����^r��3Q�A��֏��`�:'�U�;�>�YXG�/����LfwXv2K����+��/}�����Ǽ�r:����T�N���~��T��|��+А����x<�)������7�Y**+V-���>�t-�'���u{5��ه"�HP��<�d({}m��Ns9�}�K0�d%.
��i�@� �;y��<26!S�@�_�ɝ�վ�yQ�.���JC#b�ڿ^q)���_�0�,	��_PY.x��ҌK�o5��[&�����=��iq�WJ�}��_�ރ��:p)v�{�1uy7w��mm��a{�x�ɬy*���q��F���y�~ ���n���3)N�dsw��=W�����~X���|�E�<z�;������Pn��:s4�BrŃ��J�g�t豶Z��
�2��U�;3�v�2�uL���_1���5Gxy%�;�W���eԾ��ՙ��TwI����� �3��Nl��s���?�  V[5�{��w�9��>g΂�+�zǎt�����l�/ß~p�J�N0��DIۭV���w4�l�w��f)˽`�V�!�E��U��Jנ�_:�������~K�c�t�U���[X�'^P!���`��0}}A9�unT8��<1������r.%H��`�~�}����͑|Qk�sb2�C�)'׼��,#�����ayp��$nߞ�Q��Yx[^8�m��x����U#�o�cO�������u�x�SnEB/�B9n��o!L��I��!,�u�yw�&-���}����(_�I<�v��X�F+�B,G��N}����;�����s}ʠ]U��b�ܟw7m{��!�\d�Y�ܟ�'V�݄�fosBO;m4���K ��=ψ۝BZ�nY勞���+Y�'����`���Esܝ9�����x9A*�o�}��\�sF���'AV{9<��
j����N�B��r����t��zk��Aa՞���K���[��
�CM�P���Tni���_����������jO^�c뺔�6$�'���8����SP�; "+��`,0�8��%�k/�"��lvfnq�]�:��<�{��v�Ӛ��f�FRD6��<�خ�N!RMԖ��������:�Rj��E�ٱb:��O�_W�W�,�3u���UٍX��h~!�frf�^f+���6�_�h�s���n�L�y��k��v�Z�W���w[��ߘ�J���7�����D|VE®}{#s;C�(�"�CQcc�Wyo�c�_����}���b}�n�N�|]*�(r��S�Xg`��`O�-��A��&�z��n{(3�,(C�����+!1N��b����[�3ZWN��2k1��k�w7���xfo�U;}w���W��o�gs�[o�!1�	4=+*0�eA�z��H3��R*8���;����S^n��ũ��qb':�NyUv�)�V/g���&�[����5؀����^�_ٮ�>�NȆǽY�j�5��9�o���'��� t��O�����<}
p���V������^��j] �>�H;��{��L9x�B�x��5,�3>lY�ᕏ%���}��$#}~����fE���w�u�59�(o;k�e1��F-4��% �ެķ�ʫ\�ޘծ���;k7'��q�[[�(F�ϛϲ^����ϽʅcH���a��|��5f���R�Υ؇�:��������,5`)��U�Cc�k�;�ݲ՝/�W�Q��E�d�=�U�*��oZ_����=+79��}��`O�53�ح�ې��S��905��9�"'�5h�ģ�������"�멒���@�u��/�n�g?B]�w;P�
o{x���4a�vҷ}�{
��%���2��DtըQu�Wr�a���E�:��JG������>��y�H�Ԝ�{T/�``^)�r��r�X_�}�*�h\N}��/�����עܗ�*��J����쫶{����p$Y�(z?��C�;=�-�E������A@ �p[s��_fң�#W���d�s}B��c��W�G~lqdx#u@ھS���M�S�Ϻ�Ե��G�s�G�l?j�`Xݦ!ߵ��-2�}��p5�lMq4+�20���rM'��x)�w��pnΛ*�lo!N��yB�����v�zti�� O��5��b�d���{<��_��c�7���}Jr�cpE�#p�Xzϛ�By�#Vf;z�Uf�52�n��dY��ڵ&(/��BX"�nl�;�i��Ὂ�&����7U���S���prK�W{���䏴�G$~H3�k�W*U��޶B��v2��ǸNLJ���vL�^z[����d�m�]�a)��Q���e��2�)���J@Z���A"�P����\�)�M��,�\���Hq)�+����/.�o� ˅�yۉ���ʨ<�`s�=�U�4G�UC�+�(Eq���h�M�U�q�<t��z\>"�v�V$����E�aB�J�r�*,+�aî�X�U4���ect����KNEC����<�ܶ�gV�=`wP���V�����i��
zc�y5 ���ױ2z���;v��W���!)�)����1��5�"�����S�}ۀ���o3\(�L�c�AfYqq=
1H},C��RK�������|eFiS:���
���?xʺ�V��~�z$L\p4<X��.Ϻ�7�^��{�\$�><����L�������ӌ_��(� X��x�qtV)L����檘g+�ZU��wm�b]ۧa����FK��\�%�2�/��"�T֛��j�cv+�:o�{�]�aK��ˏ=L�5ԙ[�;5%:b6Ë+��w���Da�،=�����6{�]��ٯ,>����~�^^��D�^r6���1͕	�2ܜ�C��>ڇ ٌ݈�I�3-�4�szt���f�K���I��b�6�.��ͺurn{2�yS����ث��xs��M̃@�g���=#��L�_�5�o���ێ�-뾜�5��q+��7qb5��8�訡�B���Ϋ�د'���y�uM��H���j�X����������Ee�t����*27����%9pot��L� ZD<�7��}4v���ȓyyF^������[C�Th&��졐��ڿ^q-�ޯ0�ن�bdtV�^�ޡ-��6���wDoK�y&�i?�F=_x:!���i��E�3�o�8����x�:���^�W�v޾}f�}���{6����c�U�)�|r���3`��^o�0�Y�9]�^��x�iUm%�!)~
��Xg̺	�!�m�������A�l��ύ?8�yJnÎ�ĬFOvr�����E�R�����Mu������F�B��iE�^]�=�5��;W.��nF�J~�4;����Br��w�b�ME���6��nE�S����wzi������6R�P�b��h�RPU~��o�CK�R��W9�,.������k�$�����;q�{�]u�<��@��2�wh$$S�Q�<�5V9\�}������>��C��K�%�P㸙�#@�a�($yx�u�tb��
��m�mu�r[������Ul`^��'��Y�73�Ⱙ�����z�X��Z
⮦=h�7���U��E�����y�+j�YҜ|A��w9N!T��
�qk�y����l�W�g^з�ih��Ӌk3+�Nz;�{�(e���T�����x	-�ںy�ꮅ���p.���ܟXl����"��S��?{� �eUl�~��n����3e�ٮC"�]���9�KC��<�+xG�CY�'��T;u[=24SûՎ��9#c�4���G{�!�Z�b��thQ��kQ�2K���<���
�6��b��� ��Bn䊓�Ɍ��n|}y���qn^*Cj�τ��}[P5L�<��<��t����5\9���c��+������{\�!�0��>!����̳'��۲Ԗo����7_�K�,�t|�){��9�
���ȸU��=�4�����U��y��1�e��\��z}Ţ�g�=���[��_t�B<x|�m3��A�t��c0@�%�����o=�vxGF���1ȧ��Ŵse�7"��Y	��_<	��[D����k�}�6���%�γ[ᢡFuW��������Yװ3����ײY����n���	����*��A�Q���i�]W��y��b��h�����.:+!��vv��n[OQ�ƍ�e�(��g�C�^����rÈA� Aup�;1<d��!�uo[˳*u�rX����-�����8�����lOh�:%{Fj��=׽!u�5���!Ku����������3N���2mFq�5���m�k���}�V�^��aI������Ir�����da'��-��G�*���*��3�ӧ�j�(�b��oyD[��G4�sE��|��~ZV��3J�4�|D����XT���Z�B`����ʣ�ͫ:�<�J�eL���ٱ#ƥ�����Ā���~zWu@4p�Ո�s��yB�̐�6mʁe��u�59�(s��ZA��Ƣ"�"�� r�d:��vNU��yW_f>��B�~0�nK�-	��bʈ��h�a��֪���RRMy��W4sϮ�"�i��>�b�K�-���x�E�Pe�ub%���U�sI_l�Q���nĈ~	��"63��
k�*&(����A>�f�N�8�;�rc$Ƚ��z뽻�h�({�&��R&����R\�	��-�xgjM�E�9��.��Qns%y4��]u��㗽���bE�"��?�lx;:S�ܽ�,򯽛���Z`m��H��N��I,�!@<�Ja��\�p)�la�j�j������z� ջ�9U[7�-��p���
J�E�^���>��힛�=�1).���ͱ�Xv�0�a�'sn�q��0T����Pe����Ж�)��~�!8��(����Q ȋW�M�[��J�cM�y�>�"\9�:uV�Z�6Om�($���w��Vwr��x{���:qs��k��Tg�s�F{zՁcv��~�v��}"�OV@{9Z6����sw�9�ٹ�=�[��,\��3p�Y�Q���`�k���
����{�����Zy�	��{�Ep����[�b@�y���Աq��U�/�]ˢ�=���p-�>vʱ��f��i
6o'��,k��;aS}��f�-I�'��B���nl֑�;h��kd��cv5��L\^iI�tX]�ɒ�͍�6kƽ�G�:C�<�&G��u1=F�{�)�@��׊wwf���^��q��B��!��7˒T��1��6�)³^�"���
�}�`���{"�J�����ʱ�Rw���~l�Sn�ȧ�+��=T�·{d���]׊rGJsQ�Tx�2?2�A~�s�g�+�3���Q5�gd~9TfT�b9�rΎ�^���&\7d��YQqs�УT��8�ޒ�l�$�,:5
⠅�f���c���T.����A_K�MT1q���
�B�uoн=�yi��ˈ��Q�s1���t�># ��xuP�x�d[�I%J�k���f�oD���.�/���#�7Q\������uX��[�S�i��Ve�=���gM����2��Է�x�z3V��E^�&}�b�/%��ę�e�W��`bk,ֿ�� �À�Ė���L�*���.+[`�#��yZ�@����ʌG7��X��Ԧj���]^�p�}���iXr��h\k��b���ZN��Q�	�$=LqF����oVlJm��%jwo��Q�mS�a�R3ia�Jt�snO�Y;]JX�q�]�N�-ѵ��ױ̔Zx~z�;�G#�dd�ڼ�'H���1�3C�
��s��`�m�+\T����f'��{���}ʓ���pG�5�^�j�:t��6-�<�֪H��=y�����Q�	���(լj�����.��Pѫ3:�w"��*Z��h��9�$����] ︍�L�>+V[�ZxM(SϏs����Uo�[}�}�V��6�趣y�˻D.�:�|��޾b��8�q����^ԩ�U�"�ݯl���q���s���yR�C�y��<\�ڳ��H!a��#w�6�o�0h��i�ն6�%;	z�ם$,��u�3	��R;ʘW��1P�F����=��^�r�;�#��Ӱn�wa܃U�X�k�H&��Vr�
�BT��{��U��	&�)�7E��F�.�x�C��AV���Wu�](�7��r*dC�S���b�1I��J�@�q�-wK��xs�&���ok�-��z���fusL5%��Ӷ�fG���+$�[B�j��X��bbIfA�6~s�b��2q�[l��W�3�򲷕#(v�:8��e�Tr*\�����e��r@�+��
@�$-s�d���X+�����t�EL�IS���L�꺌]��m�p�Z���rb�5���;��Kǯl�G/hcv	�Z��+zN�rZ-��� �A�x���OZ�*=�G�-w�X��y��P�p"%�f��|lZfӣg`m0���j�@ǵ�/np��d��3�Co��~�>��ov^'�!s�������!����鬺z���[94�P��7�s��>���&r�sk��%�xd��sk���J��ӝ\�{V���wÄyf!e��Ƕ!��)�c���Wf�#rJ�|ᬑ!�Pƍ'�9qRR$֌ۗ���*WYw������0�'V�rk�������[]j��wJ� �9κKӽ��vՇ|'�7?SGiZ���t��!��˵81,���8-����T�i���k�����'l/>�.��w����U��*"�v&�4�ث˴ë�w��p�`Jb���ݯ�#�P��F'X2ɶ�?9�}=Q�̒mz3^5w�j\�=o^-]���I��P;I����J��v^[�'��kw�HUEE��"��� �*I�>$�) �	 RI"���֖[FUV6�+
�U�V��ڢЧ�`8��4����KU����U-k�T�خ�e�D\�2ե
�e4�S-��Q�X-�33-ĵR��,D-jZ*�.1�DQ�*%-���VV"D�m�ح�U�������(����+J�j�]%fZ6Ԣ)q��E*�Ŋ2�Dh�Ѷ��T���fZ�mZ˖�Z�E��n�r��Q2رe�j*ZUj��F�iV�J�V��j�+E[eKh��*Z��fS(i��#�kmQF�T�[j2�h�m�X�Jڈ�J���2*�j����V�(5n2`��+1����L`Q�m���ؗ4�J�@���QQY�W�V��*�E�A0U&$�*T�X��n�b��b[m�T�#+\��X��Z�*��EIR�AH ��J���J=R��q��X�6�����n�C&�wV�WpI��ƪ��l.�H5S�9=7:�.��b���w9���������)Sn����$����}x{$����i�]}Jн�#t�"�l-���w�]gn���&��^�������q���Y��N��(�<z�u�<^��Dl��^[7��Wo%ܴS��z��5�ԭ�'f��:b6Ë45�h�*@�Q���Ga�(6��Pd~�A��lف�C��T\�s���**M�o��cϰ<�5w��!,����=F�����'���W��.����X�i����/kȲ�|�#����>(.��XS��eI��lXr*��"������gU6'���O�0� F��Y��̬i�иcٔI��sd��39�P��0)+�!����άJƭ%3�G�Ge����6�"�V�.��lXo���Ǫ���W�K�b�5���F�w�$�+D���O{W�'Nx���\�/(�Iש�	�.��l6�b�i�MT9�ڕ����>᪝�h�v�8��Ue�c�������&b����,���jȢZB��ҏC��Z�������
�{շ�G��мU.ܮ͒6�K�7&f�7E7��2�G]P��1���.�(Rͽ���v+����S��!�l|��#.�[e�a\�wu��Bչ�����37X	;6Uν�9>��4@U}����9���C�����^՜9*�+K�  ,�M�pND��H��9`�b�h�L�D������r��E)Ꮰ�m��+/*/qۅ�T��ʽ�H�\B�9'��3��4� �D�{�*1]��Q��LJ��vo��Ї�Ω�/2�ɉ�s����<[��=�#}.8��J�H.H�^��yN)�"��J��vWj�P��V�bo:qF�_�Buy)k��fD�ϠP�:�尰��4���гebVq�7��7�:����n��g�p�w'�'(M�� �p����ܠPVL��'vznj�Lj�s,�b�'c��Q�`p�]�L����a��X��*����E'��d�mV�7��/#S��46:� E^�,�����u�ȑz�s�]Y�ኯ<�!T�?7^�3=r9������|P�y��U�ݜ5�.��^m\W��^KR"�m�̸�]�:K�ײ��foCX�|-8T�Z/�*o�`�D�=�+�Iqv���i����d��8�,9���7g3;S�dhc+�b�,�ܾ�s|�/(�7����9�
����<*�H9�Oml��B��������舩�}yG�5��0JB�q��68������%���od�ûwW���؃��wqwi�-t��z8��14�g �Z3�Z�T�kg��>�^�'���Rh!fhN�U�v�j�vYQ�O+�X��3v��!�[R���<�ӼE�|��f)���1� S+f�sOm1>�[���7K���KNT<�{Ʋ��F�{YS��=Gx�#JoP���nq�.û��l�͝E승Ȝ�>�5��5�<oe�̅;,
��\׌��>K�>�u�O8j.�1C�u��u{5؂st�<�	̼d�H=���G1�QSA�.�i��\9�����5��]��8��nv��pWWF��f�U5�]��L�|��#a�#�T 7��N5�5���;"N���Q�G�����1x�C�J�y3I���h@x�N��AZ�X,���tJ#��?O8S��?b�=N�q!��M�b�������S`C����*@N�}�Mj�WՑ.��9��]s�)Y:�;��C�gmcP�T�����JFW��^��ӽ�׾�j"����5_mi�6g_E�	���8��+�=%�'yѠ�^�+�����׳r�Ɖ����SG��)�c��F��5Es��L�x�E�PH���=�7�w��v�bǌ�q��8��sλ*r3����x� g^n�}����$kek�Omxk8�=��s��Н��Wkd�[�A���XrP+Io
L����dpZ��@�I�^;�:��&dY�.
�N;�ɵ�m���N��T��ȅ��oT��4)�o
��s�qt��?W�}��Mor����mX�rX��uLhp����b�O�P��ޮ�!��E�C�a>�u�y��7���3/�p4v����5Z)�ܨ5Qx��Ld�6݃c8�Rw{%�c(�����-�L��Hfz�s�g(1q%#~�?��J	�Y
���p͔��ʮ� �o�=���Z�0-;�Ks������~)_G~n�!��1�ℰ���-^���R���� �߼ߕK��v��X�`s;7Odw�OV@{5�5͢6�ԶV ��ޮ}oV��_�2Ot���'#�������p�q���Z�	����{҄��ۓy(��_�Y*O1\�_�B�^��8eb���������_��=��ÁoY��\��������R�3��V��w=��E�-J���!��r�{B^���:��EzW�zs �i]�ņ);�S�필s��$=k�+Z��:C�<�,p�L��V�VF�K��W�r�p�}˖wT�UnT��_��-&C��鸻�W�ҽA���p>0 ^T��<R�Zr���OP��MjQ��;W��qDX����ǋ)v���Q˷�r�K*�r��9�܍[T�s42�:��=>y�JyI2����_휭�p:�L��oxI�|�������, z�_9�XjT��F����]�7�Φ@�sy�0ܫh��?U}�W÷�9��N� |+k�L➊�}jٞsn[�c=2;�d[��ȧ��V�>�L�<���	J{�;���ͿmfW_�����;Pr�ϥ���NǸ�}bb�k��eG֏m{=�gbt��-!��KB�K�6����ϗ;]��ٻ+:�}�u���r�j���;_v�(�
���T<���~K%����z�{ݪ[��`�*�����,^۶�k��Ջڿ��	aP���"�t��Դ-���TI�Nٮ��Ծu0θ�S>�.�qr�[/>_B��[Xg���Kܼ=�(Z�c�ꎖ��y��=cT2k��[�٩NX���X��d<
�s�+��t�n�\7����5G1d]g[�ܨ���S�QPS@��tX�땝�}AS�1��BS�~��vԂtP���N��E�r2�����; ��ɓ��+��G�7ӹ!��z�X����X]��a�Ɲ#��%�+z�Þξ{[n���\�ˀ�V��._ӓ��<�� �|Q�v��s�ےڭ��̢�PQ�"8�)m��"dI��k^����P%�Q�ܴ˂�%k��*��j��4��T3D
��U�-p�t+aZ��A�P��]�BOL�6�<�ٔ���_^�����
��U��|�ި��WPY&�3xXs�P���Y�P�TL�e���{ܲ�o����jyj[�D(|�!
�2+�}׹�ݬa��!�:VW�㘋�;�[E��2�]��ieq[|�_k���Q�&aJl�.Ru�i���gX��6�E-�F�C���̉F�mAv��� �*ׁ�^�[�C�:���	˯��~N�y�tڞU]y��1����|r�ұ͍��B��4)b��ܭ(޺/�'/:jܬ���*N>�;Of馋�|��8l�u.��b�R�\R�8>�E�E�<����(����	hU~�2�z��9�`Vo�Y=_d���E4(���;`7���(�:���PT�.��҆�{N��*�\�����N�%,.;i�F�b�UpԐ��ҚxwH��wFf�7��b�w��k.�=/et�]X.��>����aX��
��ͩ���ˌ�q_�������B������5*��"ǣ�B`��-X}�g��T#�SkW��^�j�`�^Z�^���W���=�[��K�mJ�	�b.1�����\{�ty� �܀�t�ї2
'�4,(�I�/���7���{;��x:1�m�����<��j�7,S�$+��Tt��ucݛ0}��N��t��6��*�Γ�n��е�+O����܄#��e�����Ahd;H:TT_k.���]^��*m:�-p�7�ף=�vk��͓���e��1jO	�h�sb��
�U�FCs�}EM�E�T"���癴TؓR�{��C�R��6��U��MP��T��w-��?�2_��*�S�1xed�$�x\�És�;z��rm!~t�b�Y���L�:��4K�xV�>�ݛ�0\�lVʎuv�=����rH�~�v��N�Cϻ�!2�\
��GW�@�J0�C�����Y#K/����n�i�;�*���Br�,C�� ���6U�·"�E\�On�E�2g��x���Y�ί�}A=Trֵ��
3����Qr�|\[���Yװ,I�';+�7J��oFw58yM[����*�@4�J��o��s�d�=�^n���c��3���;�����'�z�z��<��&F��<F?P��:�!�[�3��*��ΫN��쌣q\\��%U�MZP.��#Z�����g�8㴼S�h`cB�j�}S��[�� o���Q��ѽ�U�gu�c,P���*���aJm���we9g�t�H䮳��O����-�H��.RC� �Vmw�M�;;������vp�:��	���<N,�Ý�V��Τ{Qn�
�Vm�t�5��vvh�U�	jS��ԣ���-�K��nVF@����3����(W���}��-LEmMx��q�K�ٹ[Y�]ҭ�}�}Z�E��u8�/�6�@�]_��N�}���63����2��0k��d��U�N<l����o�aqpLo�����BSqe��6����mFÞ�r�a�^�{=�����?��Z#<���A���g�=}���!A��n��B���"V���O�� c�ӂ$�8�9�T1���	��E�^�w,{���[>���2�{��#1{���$�Y���=4��h�+){ą�!�=�M)[���.�����փrX�\b��8[�P����,������P���N����w�Jkn�6�w9��/��ΰ�D�0�>���\8V��7������]w������f9G��R��Y`K�Շ$n+{Q�U-8|j�����;[e�=Y��M���q��l�����|�L�aC'�MH�.�NC8r�lg��.�^�S���{N�!��i���vC��V�� �e=��
�w��E�w5���,���m��������}%^l]g���+.n�� �����&� �[��d}���y��s�N"��q/%urWEj����2� �FV�9��	��{k69��m%���F����4��+V3[ڜ�ٺpS���P�%V�*���qJׄ��A�K�-7����eY�3��~��޻9'f���E����|]��8����pL@(���

=�-�\B�v�p �u;�-�b3uZռ=V�[�$ԐR���,uJ�c���6J֦y�L
C�@FJʅԮ{����%�s���Qu7��.# �)�T�B�鸸sc
��2��ۻ�OZf��Ӵ�J�5�qpZ��6�t&h	*�$�w��E�E��u�Z�+����"���ȧ�ꍃ�kڒy���GI�ʽn�0J�R�0�AG��u���8-��Q�������馎N#W`c�o�[�a�z�R~�:��x�K���B�K�6�0��c�v�b���c�|��a�<z�����r1�5��@���*$E!0��H����O%����8�3k��ӫ���ToB�c]WN:���wW�Dq�P��$|���b�6��O�:���r[�Q� P�C�>������P\e�������!�yCb�[�;�������5\�^g$�8W7)��%�:�`��nn-:���z�{7m��P.k�-��,�Pĺ��a��q� ��ej2�h)Ή��Wo$n�pTP��*TV�͑u�8����p�n�Z�]l	m�}|Q�$�U�]��"������or��ٹ������Q�C1+x��z��,k��6u6�s�|E�6
`{�S�W���4�F�6/�y���9c!��Ș�����.*7ם��s��Sʊ�@�u5�'U���Y9��뫚c+�4�)��dd7��dP��ca�pW�K�3���F�xkg25Y�mL|���L��)�u	�){ċ�VR�^<~S3ޡã�V_^tEbQ����{��g�#�����63�&봟�1��&�p��w�	!��nay�,鍗�bX�A�w�Nl��o��6:0�6f��Ț�N4�j
���;�p�����׋+$:��Ϭ���B���<�g��d' �Y�61��.y�d�J5=y�׭��Aܨ���tJ�#=n���
_���fb����iۏ8ΛSf��w;<=��Uk�&�(����� ����^�oP��}��)�q&��pAr2�]Ȼ�I�y�n��qWG�D+��`gҞ^�`<q���RPU~��o�CKC粫o����8�� �۫��n�U��B!�\�������������HaB�"�;��ZYR_2�T�6C�t6�[�땲��ʖ6��'qD��:0n&���b���Or;L��Ky�(v�lHە�pvU�h�U���)u�;��1(�Y�n
W}��VK»��wV\��Ԗ���ja�gGZjQ��Fh�k�_X�����1��1��=�M�������WJ��������w�-�.�)���kK{6�>S";ի�a{+WY��5n�ե���#U��ї��+w���N�3U[�:�cU-�N���,�y����M�lR�Sn�I��[u����2�%
ݴ����U��Q5a�b���T��YJ��'GM���,U�����E��cFo+̏)��x�V�������k�Q	���!.Ʀ�tUy�̫
<&]���lP��(�[�����.��a����874$IO}�Y>c�������*�,U���u��'�!�de$�^U���\n�4�o�}@���y�����g"З �C]���\x�=αC�'���͋VL8�=W�p�ݱ-!��j���t7�.F�wEZF^��5��r��\�)���=/h����`��XKN�

�i�i���{9�ú��n-g0����r�c�b�N��=m]�`�h7�B�:*b�/9�V��bdF��Jf��&p�,�M���+6��<��dS;Bb�����g����F���9�&r{��D��HAv�ݹ3�Դ*:3*�*'��,�M���ϱ]]8��i��8B��Bʁ�S8�b�!	��q�Ύ������D#ko����v�v��c�J��#�ߝa�9+�a^�)z����b�.<��r���۶H�E�w�Z�d����AZ`��|�Ɛ'Włh�cq���R��8��K�E���U�چ����(p:�5��#Q�%$��̩��R�uÜ�R��H���s@��rU�M�;Êj���n,LV��;[��M�V�2gt;K�ȸ��g��c69�t��|��}�h�ac�m����=���pN/8�/5]&6K���@�n���p���x�)!SKA�W0��t�w��.eN�����t�5�m&&{���Y�|U����X�<D�jB��p9����k��f�g[}�E��W2�J�[}D�ptW��n-�Q�d��F^$hB�a}��Wq�6�F�R��8����KR� �;�('hڽj�����Ťi�X�������^n�ް6SBf>n���er�,u��Hg|6�za�□W;�}' ��wv^��Źfc�ICe֣�;U�zq���'4�2����^��"%����*vC��,%����Jdn��٦�|R�ᴕs��M��,�����ܸ����$v�U�0o%#�#K�i�&��{��������j[��kb�%s�՘��w��5��Q(�1�cQ�feʂ"�8#���U\j[�����cr�X��R,[Kh#YDb�VT�aQb��ED�*�SL*
�5X-[c[VQU��*��*���� ��1EeER,�B�e�QM5MR�QTb���DX��j媢���Fµ���P̔�*,PU0X��*1��Qt��CH6�֨��X�*ȱV,T-l�F"�Eb�F(J�*1�E����U5����H�XV.��*���Ud֨`�*P��#mTV٤0f5���U��F0F,b1Tc� ����R"���E`�$TUQXe�,����[i(�Ո���Fj�%DHe�(,U2�b�*�#Uk"0b�:�ce(�U���X�Ԫ�Kcj�U��Z""�m����EP�k*��J�Z�Vز�e� ��U�F����)D��������t	mĹw!�ݙ1�k�N&)�,<Z��)����]�m�L�N�U)�Atf��Y��P�(VO_��6����;�=����=;�ո��4{"w�㈪B�Ar}J��SM`1u��y19��
²�[��UQ��juy(x�&}#@���!ԏ-0��D�k�.�A���Q�ׯ�X��͡v�B=j�(�[}Zb疾�ݰ���"��wk��8(-��%V�����H�����y?����=Ց~��B�Y
��O���K�*��]k]e^��4s����=��"k�4� Q����**��q�LB.�]L6�yF�|ٷL:��d�uDm�țL$A�!�C��TU�D��ܾ�ͫ��Z��WL�	�䝹��۔���n���:��ύ5_h�*�~!����hWI.�yA�&�|�O�2���ws풤>ta�9ψb�����vj��.����t={�+��l�S�G�	����g.��et�%)��t1���*uO+�+q��[�}��8q���ȯ���l*�#����Cش;����LC�@w!��]����W�;�4X���fr��+v3��R�6�
w�5W��n��Š$z��׮gU�����r���uu���n�n����9�n��M4���xIw�o4Nl޽&M<��o{jN�&4:LR<|��x*�T��txg)"���ʆ�z4V^�i�k�M�隰�����{j�s��}�칧�k�ҿ���0'��L���E�(���n^�Ź�:wx�3��VE'�t=u����A�a�xkB���=�J���R��긎�_{�b����O��m����5aLQD�ɑ�/$�x�0���B�̋�*�+�1��f�3��[�5Rnj�8�b����,���L�FR���Ɔ4 <v��G�U?i��R�q�ɥ����K��P����85V9ģ'��
�zn,Q�R�+��ˌU�޶J�}�}�����g&�U�k�<��!�)S�i�X���X��P�0��۾���nox{ǩ�aq��ĸPO�o���:.BSqe��6��W����\#vf��9���_:4��O��"}�m2Eb��ݮ�н�0&\<u"0s$��ǲ����s�&�@NV�>(9�B	8�h����x�{�*���[Ȑ�=8��>��6���/wuq��4{����aX<r��/a�����T8Mob� I�	sJ��^|;���>��������uϭ���� on�3��q�~X��;���H�{L!�}���o#��f�N_1'R&��ꚮ|F^\S]�*��W炱��v�����28�Z#+wNp��w1��꠽��/���\�I�E�9�!��{~n��9��$!g����\�iX��=�e����xN/��z�N�1��	�M�ٴT5�*�.�����8Z��v/t�*��D�a>Z�9ص�{�s�O����A^���ꛍ�ۯFo[��t����1~o}���gZ#Go�7_/=���
~�P���
��qt�X}��V�,n���. 2��Z��P^eSԯk�/�����6x�%֡�>"��We-g%��L���_pZo��ռp��Q´�(��\ҭ��y���W�bv��<:Vjqg���/����~Ļ�
|B	��ٖ��+=ו��,̀�Hb9�P��l�edu�F�H�Jͮ�b���G���z"*j5]�{uo��E`��P�u�Uˈ�P|��p�rq��Pȝ��D̻�q�d���w��t_Da�STzU/E"�����r�@�xu���=�.�6�$��{�y�>�)���^}be����v�0�B�Y�wQ~�;PK��QA�a��W☭�<y���h��ITf�3ٝ��� t:<ɝ�}S�&o>q���ޝYAv�fmLI[��5��� �����U�ں�ך$�Jok��o*��;��>�(��5iR��D`iq���H��&�_:�:�Q�+u��ee�&�s��9���/�MG��[�&���r�f ������~<��0ߕ����!Fݢ�w-:Ù��D¹.����`�A���E
�/~R$O.H������w�h8�� ��=�~�̱G�K�ڰo1�����e����Q��B���)��ܳ���WJ�LΉ�5��,��>���sUL�cо7�'_�_.2��k��lt]/��֥�؎�hŢO`�6����[��C3���1+���P�qz�L������1�8��{Gq��+j���'u�hG�+Ma҈��S����o6動;O��{��������@&��eG��e;g݊aZ~&�oiW,X��=�^|���S#ק���~��g2���CX��b\禵u^����DYvWv�0ߑ3�=$ܚ��U�*ͫ�En����1-r[�؄�
�Óن�bdt>��N�9�`�깚>�F2|+�2�W��1������������M�eR�����:p�}���^�XJ����ီg]{�@	q�x�㘶���һ{�j�)�3lZ��R|Ժ��i6����k���6:rzi�T2;���FX�O�=�7۾)���l.����N�����4-e�݆���&�Z&Q(�!k��6�����/u6:�(,Ғ�O%������SH�o��XY@�b�`�sN����BS�4�w�>.�!9Y�606�E!�m/.Gg��ï�{v��F/E���ptP@�� �T��
X�.�=��S�z��'n=۹nz6��gg!��n�R)k��B����(y��]�kB���o�4�x�~;�C�&�{�1r8n��6��I�.���\�"�� #�`��u#��}RPT/���S�wZ(Ln������YӁE2ϒ��Q,.����n�P�B��}����tAsQ�T��e���"�9�_���Ӝ��f����*������3�4�@�W�6���z�v��杓΁���z��_N��(V]�+�ܟ_�'(M��H�}S;��>�\`��[|��禍4��E+�gU↰�y�j��[�k�6�ۖy�	�܆�gl9s=;/�
������T5�0���6/}�� ��\��2�Z���"�MMt~�Z�!�3���Ҭ���@�>"����ݜ5�.��}y�q�|{[����=�e��^�h�� �TY��)6��S`�oa�K��v�5��
�E�w���Y{����,�f�[���gN�z�d����u ���ge�$�W[\�(��Ew_v�>�٭���f��Y��Vg+B��=�Q�C[�
}҇_	ə/M^��!ـ!7����x�r��|����m�"�h��{!�rp���������
D�}�lث�Q#���dgZ|]+{�+G!�Nm�ݚ�į|C8���vj��:9�Ԑ4K�G
�;wq���b;o�8f�ꞁ0v_e(�Js#a�O݇��ٰ��bU{-���3y%��|!}���·z!ǃ��&����Ҫ�^���w!���]�w���W�3�j��κ�r�~���+<Ǚ�����ֻ��p�p�:��:ƣn^�Ź��N�}�_������)l����	ڮ�>Ʌ�W.�Ө�ї����E�o�rs�1�R��]��\�yɫ�+�;����`�בgѽ�ȿ��_x��r;b�!�u�o��d�Q�{���Թ]�K�u[T�)��b��Z��x+e�c�d���C�;ك�S�fS5W��S�uܑdMˎ�ziN�Z���(�����F+ji^5.��X�6�����+��l@4i 0�
.��
���m��.T��E2!ζeE�|r���87�fx=}����bd«J�D��F95w4kQg]�쥍yX��D�q�u��0ʵ�5-��P�8#���}A�R�on�V<U�����1{b�l����6��:y+��rսY����ո{.k��'k��Lz�ϕb7z֚�Z�KsN�+{����ԝ�a����������z!U�!�j#V�(DK�0�mi�6g_E�BEe����_T�(��n���Y&�[n�,r"EyTG��Ems��2Eb������cн�&�n���=���m�f5ϸ�,�`\�f�����U��X��Lhp�>Y,U��jtv+���.��ݩ��M�eߗG��������q@#����
ǃ�T�E�2��#��s��D���yQ��yu�y�[�~�\c��T?w*g�Npyq%#���5
���i��V�2k���1G�S��l�f��^;�Wm�g>��8p7�+Da��1!C�S�������lJ�
�d;�رA�q[��*��������U��v���:�	xz橸�'�-7��ݣ�F�3��[���K9�9n60����cr��Z�����w>=��_�2���l���PnA��8:&σ�o�>��O(�7xO���z�4��|�a�>vʽ�O��-�9��$G�����-�t��ks��M<�S+5iW�n�6���y�Z)����J�Q�Lz:�eݲa��Sq�)���G��y�H�� ���E��z�8�d|�K�7V��7�E�s(���J��qHF�-+���]�݉���R�2�Z�,�m�9n���oN����v9�=���i�3��!�n�H-�y6r���2:�#}����&��o���v*0$�G�C����Ǡ�:w׮�W���P|��p�i2$*1�:��;q]������{2��Æ�p=2�0����{�,ޔY����:�wteT:*+n���g�t݊�e.�a{�������p��s!G��;����[9����{���Y��+��mvP���db��',�A��q%��U
�����t(��s���N�8��gU6�=��H�4�%Æ�߅������E\���x-���#ǃF��fb#n8���U��W�A~�D8�j��}<�(-q�]Y�wW�F���+�i��^�|N��^x�5�ް"��lg���"7O)�j��voTS��N�O�±.,O<	P�趕*�lJ�KM�:��;�}<~����C�����CJ��I��c��l2^��+�;5%:b6Rj��Y����緷��)�zY�F,4;j�b�\Y��ɂ�l��/y��+���筿�4JOC�{њ�ɛ%*Ŏ���fŭ�)���ң(1�� ��j���\!�yb��3��R�G���;p�t���ڱ�e�f]���15�.f�}�ԅk<e���v	zv�=:�����������}_.~Qq���"�����V���,d ��+$��
�X��%�������|�������6LÍy��'V|�����ܽ�,�8:U�u`J��_7a�*��"���Ɲ��+�����T�k�ns�{|�ؕ�����T6}Ad��sd���s44:tQ�W�u��gz�fmH��e$f��Ҁ�ю�s�+��s����X4]}�U������ ���Iu��?�^1�:�[Xe���P�%6�):�4	�s�FF4oUj�7��=cny,�e�.�z�(6b�CE8i��h���!���q�E�����z%�;�����Ty����U\B����y��Aw�L@��ZQ�ޠ���	�8s�������grW<��&�Vv���dh���C�=gU ��|��jF��Z����]��+��b�x����ϟJbT%-L�1���E4��.:�Ou5����+�yf�޻��hNK��q�s�Uc�QO�L�/��'W����hH�/�9��J����~�6����PR�qҲ��3L��0#,�2>��;t�uӻvݟh�Fx�i\���1��k���s{D�wI]�vY���6�t���r2n��ka;,ح���n�\����������;�zfc�D��Uy$�\b�m.�BJ񃙜������!߁��h����~�W�����Q/=��,�=��Q������6��fg�w(תR�V +B�}�>�L�b��vW�=�#@�{�L��Cw���(��\���(G-r��oE���瀭_`k<�xuCN��-����U7=</���s��`+q�]�2��������AA�7 sX"��E5_@�+��W�W!/���1w/�%j����u|5�K��;r�m�E�
�<��S59����V��>4�h�*�~!���䆏x��V���A���{���`m�{�jF��6%s�r�a٬�y���&�4K�Rb�>36�gM>��^zr��6��X�]&�>�t1����+fÐ{(Ň�D�%1��{�s)�����-U��C��'+3�M�~��(C���,C�� ��ۺ�RY��d�[%��t���H��D]aLk1|���T����O�P�u�����5r��(x�J�zg5F�n��5%�j�U�{u{5�클dT�R�_ԫH�7�\(}��5<�-o��	әz�"�
�'�ܙm���,T�&�o*e!ފQZ�����O���Q��{)��-;l_Ij�(�v.^�='����j��(�zX�S�"h�|�X�GZ}��ż���B=eﺲ�ɛ�0�&`��q8�������"'W>�v-o�j���t���=�Sgk�`Vp��-����Vec\��n���T����@�\o{6O!t%WUB�ӭ�Z�<�"��r�����(��룄ob�p������lҝ���l���2�@���R�'���Dxᦻ������Շ���P�?;����ӂwj�;;@l1�9��|����T`��47e�.�Σ��� ~�����Av�9��]�J�
j�'N��޽N�ј����	[n�;���q\q�o��׋�9�����sM��ƭ�#4�i�+�M3fF��LL��ċ�X����� �uq	�O]��|�
|�f[���\�G�[����'o�� Yv������WMu���>�:Gk�����-��8�ʜi]�q�Y�N�Oi���u����U����&�GR�f:05���(�wr˔����q�[V��A�����N�mZ��|C��K�1]�k-pxfۉ�G�=�ɗq�!J�,aJ)�fn�AOrl�fQ�۠��+_d][%�ܥ
v��"�y��!�qR�qۆGIڢCk�ŧ�)�q__>yJ�6ڃ�V��2�����Oe%�m�	�2mk�hY����!���V!L�Ը����M�u�k�����
�U�����d�rc���Ο"���Z�6����!��h�u���=n��B��e(�:]���7�ū��a��&b�{+�l���&�<�aZ��H�eCX��=�l�w�<K&��})n���(�5����Be^��vBA��Y���}m�\z��v9]l�/b��{Sk0A��P9���,r�3�7C�ˡ���_*�Eu�hm2.�qS�U'4�z�|}��2HV8vcمŰ�}��ը�A�-d�ǻH��f�V@��[1̥�%K쵙�҅�1���2���5�x���O)Vt(���g�֧_R�0�����T�]��-�Ê!��IQ�	�tq��������|�:K����OlXK�JSe��8ǡ���V�y���Z��W��Ey���lӤtf�V���j޳X�:a��(b6�n�Y�4�;n?�
����Zĥu��[]�+���Yk�D'�-
f��TZ�,�� �$�^w���3-��().�k"U�`����򶀉3Z�[۟s�ym&�sRVE�������2Ϯ�cEP�d}Re�=Ct�2���}�q�r﫝�Z25Uj�\-��fʠ��1eE4�O��d9@VQ�՛haj�i�����|-t:�N���g��ض۶�f�j'����$�,�I ��� ~$�R����KB�B�"�
"+R����"A�NC`�����ADEkQd*Ս�Rҫ"1L�(��Ub��U5�Kf��FH��Ab
�����E"����Uԋ
�Q��
�R�1,�T��Q�#@�QEQLq�1d��(��dQDՕ�EEUQAf�d-�*�Ub�H��(��AD��L
�"(�D��PX,��hb`�D����X,DF��E������ QDQX4*�@�b�Yr+`
)T�((H�������P-�ɤ*̤,EX�����UXehE0��"0��T���(�D���E")*W��1T��X�dXQ���
("�ڪ
(#!X�5�����1��*i��P(,bH�H"
�ղ,(�*�~��>�<�>�y�}��r�ڗʡ�K�{&��S��'�|l�/�/A��P���`�6h3z`�y�o!�e���X	���y�{�=��5t�9�7���(h��"s��U]�ȇ�x���܎� ;+m^��5��+�����U,gU�O|���b|�cۆgê��bGN8��Y������z\�b��� �s�6�@���`���D�zx����X=r�3��Cs���Ń�+z05���W��
w|̜�_�~^=_6:B�o\*��o����B.���9��(#�lʋZf:ڧ5�t]O����n�[1�!�(|H�ǘ\D���|863^����{�C]��[��=�]Yp޵�����Q7S�(*��o�EMs��2B�p����9��tj�Liյt�[���u(V����}os�T\P2a=�>Y.�D���9:}���N��ba���=
5���Zܝ\I������G�6�hP�������5�7\�y��ݵ�sEM]`�q�ޢ��a�7WPS�4yP�n��>u����+Į�'
&���tQ�8g6sv�F�
^�v��xom����>��r��ju��E�oZ��ܾW��O�=�{�ɰw�r�/��v�^:��ЩCK�u��ɷR�Z�$��kx��P�uoLzƋ���;L}o�J1[��˼\�C�cC�et�YҜ�ٚ7�#�!}���d����q��.���K��&�V�N�.�{��v�(������Wё�Y�P묂�����S��*��>?k�b�vJ���$*���#�2���uhqʏ�'�ֱI}�̓�pha�`�����Fr�)�^:�}v��j\��zr-�y�TXj��N��^�A�L�[^Uo��╯	�M���+�ģ�Y�X��[�+9����=Ό8��>vW��#�ɣ�4��L�"}u�Y]~��9�:�ƂnI��,~U�=��w��E@����l�[�	��-�\x
�+s�fT�X^��L�h�0��P�܂������G���ç�S�xz;��3�"����;�QnoOF	���An:���9aD�K��[��8WLQ�T�B�]J�X7�r�0+R�v�6\e3�����R�s�<g�^v|_�k>M��n��؇�+����[*	�n*�&U�7O3Z��S�������hgm�a�9�Y�=�q%��O������)df6���=|�^o�K���T��K��RK��Or�~�$�@�a��H��(s�я5+�T~҄�my�;6�ڏ^�M�Fr�3i�
�jNKq��i�}�}��ؽ��'u�� QTS^�����4+sj�ŜsOPz�J��
u�^r���Rl�9��]�oEX��6Ѯg�a�)�`(�^�B�J[x���%#�w���ޔVR	�U��N��R�.��(�Q]������������(�|��y�zK��Sޕ���=]�D��sL�G1|��~��E<V�|oru�T�,.6��H�=��e>�tz�����k���Q�#O�O^B�P��"���={��qz�L��'m[�VA]����-s}���JW�l��
z,��a��;�N�PYˢ��^v,���#�^m�p�������<Ժ��^$����j��K��Ɔ!8{��}��~=û�븎���9\��SIoa�U!	�v -&���2`�^�4�+�Br���){ċ���{g��ˮys��J7/۽�U$'�|ن�bdt>��M�g6L��kC��H��pN�v"��m��/v`�G%X�7�YI���7�����Ӏ]��ض������3B����ۦ1��{��������?*t�7"�NB>�E�DB���.Vx&|]������S����N��7[��J�2�t��z�)��h�ƃ�оp��C�:���	˺I�[.�^#./_���S��D�<5=za����q��KhP��4F��[���&h�i�V3�tC��&�vX6N��=EV�vkت�swr+>�����f��^Ei�[��ZG%�m�(��hj���b�u�7�H��a�9�T�7ȿW���Z��EJ���g���\vd��l�l
0��n��ܭ(��A�u�rш}���δU�䷰j��թy,�Qgicw�����%�P�Z<��jƃC�!9��'�+������l�]�b��T_�a`���~LR�~��c�un7b(i�Da�ǎ�{���-���D�9
�B�/V�k��k\3�}�²�?k���z}����aA�#B����o��^�Ÿ0��@UC�
�h��tG"�X��_Nۥ��wЬS;��Z򧲶����ަ��8�P��Y��b2D,��P�u^(k
㼅�C�d_��BC�Qd1�u�fm��oc�v�ˣ��x
��/���ꆾt� ��QPE��plvuQ�j	x���-�Н��������]Y�����k��?VR�.�~5Ғ����&t����e�Σϰ������6��j/%��Pm���|����qU:8:�+n���p����ub��Xf��&\�.Bݣ��ψb�8���vj�����gi�^�[{n�c�k�z�Wt�h��m`�F��B���|�����r!)��'���U�r��p�:E����It�����d쾾�3��{,l��r�Ǒt�B(y;e��\%,+��r�9輫3�&r���U�����g�>������Ʊ����0kY�S'�K�_�Qo��[6��F�ԓ�nT@��z�jy�E���ΔB����\-�>�'V�$Yw�g!����8�"��qd����T�C�l�ͭ��Qoè(�N��Y������k�[O��%�ے�{7W��g3���禥=�m���E��)�!�u������ Pu�}�TTA���i]�'�X^�ֳ��+�}�,��ch��O�C]��,���ީ�ou2,E�����܎��%�ǆ��@�~N�_�gݥ��k�ϡTD3�҆v�3UO.$��c5�uC7D�Ʀ�W����=�
Un�>�0�[��z�-����!{��/�uD�g=7�x�Gj�o,���޼�j�������|����
��[r6�x���s��P"�B�wW{�ҫ%�VΘ�%�{���T�C}����������צ�fu�A�O��02��z�a9�=�*n(wM�9�Ǻ�6'PB"~ߌ��s�L�vx|�,�z=��Z�zS�t��^���@V�u+*�X=���_M�Ό��j�F��t�7�:;q'΍n��P��]��[�|{���w8_W�3&����ޫ���C�b �7�]	W�y�<�`�HIי���)�R��R�� M�y̓��,�1�tSr�2��EK��M�*\H������-������Z���=��:P�T��t�gbb��=��(
��a��y2�������*���U������1%���a�BӢ�H�*��Jr����s��C�G��S<'8<�,�qz�������r[Y;��.�t4VGDҭs�sd���^2�U�sϬ1r��Խ��/��ׁǗ��蜡����LJ4C�x.!�8�X��5g7}�O�������:C8E�T+�����Vr�{ω���Ǻ~Ū
���+]B���,*�>�t�X})�v�x`̱�6�Y����K��#[�@G�E�MWB�V�uxj��Z���a�Eo�$2xu[�@[^�Ǧ�G�h�A�Y�\"���^k��{�+�MU��J��L��z�Y��8�ѝ<�^�Ӫ�*}��cw�O���~T+���ds�fTAکݳL�qz�y�;Q�Nn��#ز�1�1|�X�4a�+��Q��r�gH�*��-Zv/{U��P��o"h[j�(ᥥ�[P�,����2�Ô��}ك�V%%XuL2f�M�ҵ�v�]�&�/R�ۨR7D6)�I��>�U��A�N4���L�R�r���kB��:w�P�W�M����u��$�;�V��r��8禮�F�v�w� �K��=s�"�skb~"�6p>1�,TzU|��j�Wr���8}jfU�ᚏ�I[��X㼵2��_+�s�����>J0x7PlC��f�qU�f�,j��-3k��9�	ujQ������Nǻ1�)Fi\T)���BY�A�m�Pv�΋zR��ݜ�ۆ��6=蝮:v*�zvw���b�
B�bߔ�n���ЗK�-�79�NR4�.�*�k�����s�V)�C���͝0D8���M5�����=/;}z�������(71|��~��E<2���}��r�X�y��g�uy��y���j�?`�di�V+�*j!=�T�:�+�h�R�,��2��b�g��w,I�������*?a�֦�N��.*�;a���9����6�i�§�3�>U�CΩ�eEBhV�7W���,�B�B�Ç��W�{*>Kɢ��[��"�a��r����g`F�����xF�h�"�tG�ئ�D^�s
�6������T�SAe^驹3��n�uw-��^ޤ��$��2�y�<hm2'�t��m�Bse޹�n�����Ò���Å7qc7:�$�+��)�G5r��P��t) -�SB��zM�UiY��P���S
4�����{m������r�JOwN}C#��ڿ^q)�[���]I��@>U�\�;�Ú�!]��W��}���֡�8XtC+�<m��@5�X���!)P)7}������m�
]�k���7��d��<�W����5�S�"�NB>�E�`��!)��E����f�\&`^M��Q��`�}3�i�Ҵ����l��_h�Ɵ���"��(Q{Eۆ���Y���ٻ��эJ��r����sUŠF��?�Aw�)��ZQ������W]����=W�a�P}/ �r�	qT�gi���ׄX���C�h�:���Ty�f�d᷸_d�!�dI�c62e.�Wݪ���#��m�E`�W���,_�jy��D��
�,���u�
�O��׶�,�9_k�*��w���z�j���v��{�K��J����}6�p*X1$4��i�/yԃy𩜦�i��¢��GrJqww4�_/Wq˷�e]��ʫ�/�	���DH���ܥ}L�w��W�/��Y�r=��ۚ�HCh��Y�j�RםR�j��Q=�Z6q���*z�m\��v+u�Q����0�&���|��ں�&�T2���,DK�G��������;�=�;�mr=q������ő�c{u������B��ʠ4��wRu�Y29Emj=ˮ��=��Yo/k1>}�JF� ���.ˇ8��*����~PӦ0��ʽP��P�����I1���vs�/�Aw�ǹ�QNB��=���z�5B�������z�x�Vj�u�Q�
><5M_P�ھW���p����L���ǧ�s�^[^T��=�
��wп+9�Ơ��6=Z�$�]�~·f��+�ŇN&(�v������w�l��"MG|�~��v�86�^{�X䚝ٸNnR����1�6��a�w��"��
x�0J��뙞>k��3G�2��/��^��d�uL�o�]�/8�{������vGUb�7��zn���=oӷ�a����+
e�|�2��C�kZ+Â�V����mÚ�*�[��U�a�qns�S�C�����������1���TH�{��G�,��gػ���v��4z���x�����lכ�v�睢��Nub�3�5�"�L�2�KQ�vV���j�t۾A�F64�z�5z�s��!�p�#��B�J�y3J�h$�sNܧi1f<�"��5Ƴ7R�}}�w�+�~.�F�5p��FX�1l�]����~v��g��]���aN*�vo��}\�Y(m@�pus쫝���6��j_�F
D=�x��s��3MN|p������_@�rb%�����Y��t�
prPV��=z�-����!cz���?oB���e�l����$�T9k��m�W��x�lv�|��
���r0lە˫�F5�ַ�E������cZԴ�ɵ�\A�(�j"-4��"_z��Q�֘}����63sy��Y���,�.CSq`��9�}�xѿ�PA�O�o�E@4}�X� �TjP�Y��W�9^ɏ?F%N/TW9Y�ˇ��/O�6pD�8�9�T�R.R+_4�:�r==���ָ�^�؄#K��G�{�WJG�xeP��0?"%�?e,�Ĝ���=$��W
1"�x�h�U�X��6��W���9C��uu:Ce��y���np���'w[�����H�Yu�E�����"��P�Wm�`������Ʈx��]�+�.�l��S�_^�:�]-�ŋ��q[��*��>?n�G�k²3�,��t�g�k�����P�}Z�����Ս�i��À�,Շ�X�}z���bJNZ�_��u�.M.�����D�堭�y)���\��N�Ֆk`��ы:��5'�A	;(	��۰�ڟh���+0y4(v�U���ghǻv���}O;��x�u��i|�%�R[@�˽Քw"����G�פXVugK�e�\�K'K+Ⱥv�^��z�צԁ���*�q �T����3W\��]< ��9I��/`�J�CY2���E�>J�\3� �4��9����濗6�j�ЮoIn����++��=v��c�N"AKL@�^���k{њ�vN�[Ž��:]К��_.;Ob���g,7C���Z�z��Xpk�U�x�LD0*��[�^J��2T�⑽ >ܣ"�+���˲r:�!�Q�m�w��B[<	���1��M�[�	S#FjY4p#X�V*v�R�%Cw���!f.���ۧ���Q�zEL�s���K&�v�����i�5%��X��'�ʘe�6{���O`�6�æ����]��m�Z2#HQ�匵>���{�����0b��E'|��i"�
�Ս���դ��U�t�v��Ys׹o�1���1��݉]�0���Y��W����uy�;(��WY��=�
tw��#I�م�&��g����"�;\KoG$vR�I�{�+�\���rw�ukwJOU4&��Ue�B19�GW�-]��n�9.��N��#��8�N���6I�s�2�kWW����3�E��-�G]�7�7Nd��*I���Z��{V��C��y��T���+kt���l~�PH��-SܵrSB݇�e�������7�1�����r&�E�#�gW��A��W@�V�Q����֦�<!3��DOg����*�R��YH+2aFo����\ܨY�g�TMN�q�9
n9�*�6U-����I"���I��3���]��rvP!Xࢳ�I����\1l	q��O�(��Ft:�]�p�N]����a�]��t�.����]���a�mf�/s�vt���5n�p
m�x��j���¢�r����ݻc(`���jn�-=��մ9G3�V��NJ�v.NZ�yD���:|��%[�w\�':�yD���ѡF��ꌬS�H�ٱ�?oS��E�Y�TUE4gaz�@�qjv5K9Ph�Qc��o]n�H����}��e�Ϲ�rN�QY[ܯ C/���/�_+s�mr�+`�(�2b�)�,慫2[ٺX�G��4�+h xL�_1�0�D��zw�gB)�#��
ojy�������+"+����+Fݓ��kI(w�fB�z�+Lv}�`��ؑT+����#�^�So ��m��̠�S=|���^�Z5�����y�ٜp�"�%n5���Ц1uu�E3�V[кa8�)�$G��ځ�N�N�7u}���.{����CɉPPX(��,YH�#�*�$r�++fYTQ@�0Fⲉ
�PX,��(���*�TQEb
(*�¤���JŌr�`(�,TH�%dPUAb����#PUZC-PKB����B,�2E�`,��EEX��b�TbF�҄Ub�AAX.�TER,��QE��R(*��Q\�Y5�h��"$PQH(
"*��$b�*1UX�ԭ�2*�Qm�U��(�H��+"�IDY��A��������"�F�F(��"*�TV$QH����"�"
# ��
�j`������EJ��"�()5lEb���
��#-,R*�\J�V�*����AQ�j�
E�VV*Ȣ���-��X��K�x�vCǪ8��&�jsɝ���nnN���X��{y��R-�h/�%0�7 �(�JA�Mπ��	%���q�����Yُ3�#�:?j`�k���S:=3���W��f��I1����|��bq크s�����C3���g�GD��)��ÁoY�t�F�����tҜ�Գ�R�9ʊ:�|:!�>�ǋ"56jz���E��l�!���w�g Xe~�
�r-鍭ܨ�x);�/������F/�,p��B��jǣ�\B���Ë�m[�^��M�Q���˾ڮ9�½bV����A����|�G<x �Ξd�����=Px���G3�WZ�2@��vdkl�sn���/�g�i��-i���?L�W�I��T�>P�G�z���ϥ���sb/����5��b��,%���r���&8��}���5g�Q���8�z/�U���G)+��GXO���H!(P0R^��'q�������"ma��<�g҄>�i�)��6���OWϲ��wW�GR��H��m�2�!~{�{�0��L�R>]&-�����[�UL��%��N�^�����h��+�1wV���Vb�v���R8Q�!#2��9�\�v}��^�i;��9S��P����̤��7Mڝ���E�Va执P��6�Hf�出M���58C�]'�h YpQ͡�oOMp��16d���i�#��M�ga}N����V�f�$#���m]�Ʉ��p�j��MS|�N�ٛ�c(�Ԧ�uh��^�Z��ֻ�T���t�w>��4
��OC��a�ئ
vr�r���oQ��
ܾ�Ż䳶��i�R/��a��EF��L�n��޿�`z�!T41�wC�n�yr��s[��{#q�`l�ʃct��; ��>y{{��h����y+�����ӳ"����\�+��"��W�Ķ%oW�r}ن�'Cc�����_��a����଀e%�����펩.��;�2	��>e*��u_������ܸ���^�	m��%�a6�G�nv¦�|zkIռ)�|}C��ay>CXe�\w>H�d^I�m��LN��7��˲���!�*α�����z�)����(����0�*�n	�OO2�2��K{wT'3��T�:��C�jȰF�+J/�4bz�"��*#�3��<W�I]���DôȘ7���%�B\D$c�#�6� [��!3���t�)r�5�l�V1K��o�̗1�ơd:�{˳5W�*c��Pq)��5� �;t�A�m��Cb.�ξ��LV��-��U ��ۣ��^t��&\r)א�?b���^�����N����'M���B�(kl����\>~�lޖY�i"Y��zS�����6�H�T�E"$���Tb���yw�pp��#�3�q�CM�0^ՔkԵ���Vr�p�zn�b�AriW��޾S�mȨE��G=n��ɝ'�5�'^f�
�F��(�_ 8�G����yS�cc�o��]���ˣ�Z�<�lN9��i?r3,��G�7l-�!�
b2D,��4uV(k�%�9�`�v��6�efm]c�Z��@~D&}]BZ��nY�yX+��B�A?�i�a��k��>�zn'�͞�E���p���\���9�it}�hO)�S���A{ڇ(��v)�nN�yC1t�δoS�|�mMy>��������k�@�3�&8��Rz�k2��z��f-�3]�{��|��nh<;�R�YL���7�U$�d��2qk}�e�xe68b��X*��[`f��gs��iM.���:�E�e}������ZrkG�e��S�U�ʠi��S��cR��N�N�غ7`;N���9�����Z�R�R�����խ��IVԏ�F]<�q�{���ov��e��0��͎��]�U䞾 +��uQ��z�n���U>�1+$�e�<������N�ʅҖp�`�<���Տr�3a�CkS�n��q����ϕX-OuSW<zKG/bI.�y��g���Ʃ��͢�T�%C�{=*�s����:^�hEl��u�9r�ג���v��~e3�9ٸ����6$Py\)9h�c�U�=Q��ҟD.{���,�,g��r�ݻ�\�b���z��94���o)�O?H�i�=��T�Rkb�1�F>Jå�"8��q��eCZk_r��8?��a����Q֦��W{U�|��ю�#6�Is�ůsg�_��8���0M���/���/�ȁ'��[u��V�b廫)�5#�ac��D�5�:J���x�+
�p>{yҞw(Wv�[}�����'����H)�A�U#Z��S�Ū�GV�=v5�\Fo.��_�4�g�D����x!8:�cr�׫y@{Q��An�¬��'4PS�5�ݎP�ިg�&���-�;��HL�ö����4|Γ��K�H�U�VV�q���ݦ��sl��Y~�~(VMz�/�CT]'b?dvhԓ^O_U}Mk���n_�/dʘw�wfy�L|���Y\���R���%+q�M���Xsݡ�)]��+�a��3v V��L')p���P~5�>��Mv+0�t{�(jv�ļ��H��{�ͫ͢g	��$��U��C.���x)��M<wW�y���lj-��9�y�J�u�ź�]�w�5٣(�#�u����1T�7b�71g1D���<R�Ԓ[�Q|�|톻��m��z�����̨�(@HUMR�<����{X�9��5�/9�v��y�/s��ɧ��4�^U��=��񐩾�]��qܬFA��e�;}���Qn��[�����}{=�q��O@�+��qR���|�-(l��句����5{,7{4݄ݻ��Ya���3M�ys���l.l�횦x��cwB��@��'m�M4%��^��ܱ�`�y3:*kL��g/�?t��SU(>4�����KZ�[Xx\���:��֖�j��v�1]ocSjۇr�6$�R��-*�L�v<oƱa/)�/�owA����t.���nOM��x���Q�=[�Y��eO�3�Y��^B���Z�򦀮/O�����M躥*���<��3[ѓy��D�}���ýB��O'os+��NV��I�Z�o�H���yp��].a]�&�g+ۆ�R~V�_����4��7;izF�&��V��bgxK�7��yr��r�u��W݆ܜi��fzN�����g$�۫".�E:���^.9<ȧ^��"V��&5�9���WT�ó�WUbm-�֝\M;�'o;�!��:N��ky�qU��z��1C�=��:i&9?������|�J�W��S@pQ#CQ=� r{J��oT,hQ��c�����K�c���[��u5�
�F*�x��6	�ba��6v�K���7��R�i�7��~�Sjk�>E��}����\1eE�ށ���;3�Śb��R����ay�Fi>>�OXg�0CJi��6�ٮ���ɝ�ܕ���8��9����������2;0�5��aqU"�g.ݾ��3yk������xj����]�p�٣ц^2�In�6_
��d��Fh&��A��d�E{.�u����4}(F�5<��NJ�eo��d�4zh�5�����Ղ�Ӄey�h�t���Ap��r{J��'�D�@*��T6/v�p�:V��G$�|lkC���5�V�B�yV�%!���
m���z�g�M�'B𡣱�0>�y��m��}�r���'s�/A��J����:߳x�e2�;7]+67�p����H��o��V�ٛ:^�R�If�4��٦�k�!�v,
{g�.��!����s�=����'V�+z(��"���t���]���j���d��ե���������r�@���4Ă�W��ro�uYV��a"5��1��{D�؉�����j�Ib���K	*�r����c����N���@x��^6��R.{��,-ے�	�
GyuzC�EVЖ����WT��G���So�iNy��=����a�g$'�*��P�[o:el���ԗA�J�_=P�ߵ�-/�u�z�{_��Яd��I��j�_�z5�٠sy߹B/\J���h~j�c����yrSp���隘��b��HM����x8�U��~MBu��w=���mxW��^ɪC
ޅ	�m11�=	���}�r\����o�Y�Nv��k�3e����Cq)����\z+o��u�v�B[r�k��܅�W[�+7J�0ѮyΣ�V�{���]�����(��;v9���'��M]O*'�Vj��WVN�D�vV��NM����ѱ�[�Xmέ��r[Vs�5�ϖ�����ӲR3����^�¬U��Ŷilv{����_�Ls9O>���z��cط����pL�����R�x�>�S�C97V^a���mOW+n�5��pk��7�#���J�'jxa�츍hm;N���ی�����E���]�S.s�p7{=y�4:/��51R�sj^�]t�F�NWu���J��6��n��n���E�����­�b��]�db�	�_
t$.�Ԅ�uQ��>��)w@���!�?>^������A�N&��D:�lO�A�z���jOR�^�m�H3��h({�,���u��/:��¹Gћ��(.�v'�Q�ll�X�y<��D�m��ݛ5b|+޾������c� ����x/����xk,*�Ħ`�PZb�1�[#=�E��rne�R�6�݃�^�85��%�zc�N�kN��&\5NOK�z��Cf�H��Ts� �y1���*٫�V�uJ]���˯p�ͮ*w��G$qc�I��[��]���i{Jg�=��X*���(ti�I�N�����Ƥ��Һ�^��V5��Bp$�w�w�7����[Wڈ�.��L�#{��Ts�敬-������A�*L��U˧�oaR2$^�HX�8��[\��P�X	���s5 <���Oݯhz����X�]��>��'7g9Yޞ�����6��Ev��'��*�
�������i������v��٥x����s��5덮�<��N�a��@��4�FQ�����1W�/xj'�t�ؤ^�ڝݱz�o���Xg�0CKK��m�٢8���p�G[�>��Ery0�a���rv���)5�k��{TE��/mFk��u����[^��X���c%ר�~z˿2���xˋ÷��f�J^�/3S^����PҚ�|���~w{�����Q�m늺XH����B`��A+���`ܐ���g��+�/T0�+1������V��J5|8�����SmT峤U�X�6n|��n����y9c�ՙ�u=L[j:�'p\���(;�.2[�Ԁ즯�,7�-�n�C*crM	&Vg(Y����\�)����,g�c��C��+�^��>�G�Z�e��_#�Nci^�c4!����α�qz�Ҙ�0��P_�4�ϯ���b1�7or���]�}W���+�Gշ����:�ٻO���s>�ۖ�/�_N���P�>���]��~	�}ߝ���vں瓧0 �ZR}~���M�dU:��O�{��j���_r��}�=�cYɪ^���}U8X��sZ��g���.f�cX�|�Ts�Һ���Ү-��ܫ��<�`��!+�cC[>8⫍��Tq�X��&{((��;{Y���3�>��;�Eʦ�W�F���W�[����͙��W�w�)k�KN?j�U�\R�N������{�z#�ɉ�D>-�P|z�������<�tU1ln;L�@�m*<��X.��Ť"��(WJ�WG��׃n6\{��녜�8RG�����2`C �Q��uʕx�΅`�Mv���9×}B�Z��)	�M?�;�t7�nl���8������֗R�����°i�n(*5c:�CW;� ���e���j�I�f��7p���IHޜ�(Z�o�B�uJ��=[(쯑su,�Ih~1��U�R6o	u ��pT!(�紷)h��-��a\ ��l�>�V��;�!?A�[0j�n{�/���g	����W!�a*�u9q�)޹�־gl/����(�}o@(*���3��5���ŌgR�+v�"ݭ�+i���I��2��]O%��$�} �vV�3�׹�3�L|���6�u�I���(���s���&�ޢ1k��C����
�"�������]�r#��2�m��ι�,�6{�+��a�F
�m�+�n$�9t�w�f�� �n@��VU�"ٽ���A�á�.+KJ��'V(jh��G�m����޷x�=֫�����t�eu]깑�Bn�Uh�\i7�	�����E7NU��O�W��kT3���N��ƖY�w��ZH&zk�{ǯ�������p�r���P����lt�Ӕ�鎱��#Vay��a���7Cs^-z�X�:(��J�˙w�'T��J;�07ء�}K����1Fyn�k�b��lq'F^n*��p8V��Yٓ��ҝs{�N�Fc�VagnGgjLw͕Bm˼�Y�����8�D���s5�qU�O�'J.�M�ǹ��=ť[Κ��u6�1��Y��P����<���5%}�P58G�5�� �B�f�m���3C�7�m�V��2L�Xէm��Y����� S�M���R�?�K��U�J��[���D���	��j����� ��Wa9&3q��!<���/gN�|{2h�R�m���k��B�Y/sY�<���5���@ݭ�,�k:1��P^Z�����D��Y������U뚶�v��[xU�2�>�D�b�]��<
��ݛb��5\8]�+Px16^!eoa�(��m���;��q�D6��QF�z����w=2^E����YrS�s�gt�Z�w!�tţ��IT��l�.��i�HD`�e���D+n��}��i�WxmZ�s[�ە
V�P��r��d��:��I���r��,��ZЩd4�e^k�|2N��"�V���������˾�.��u)�Mt䝕xy����a�Sm�="ت[&w 1Y�� ��RGK�ܶe��B��s%��8{e��}���^�cޱ3���^���湅��,��q�M��ʡ5���i�6#��n�F��R7xm��7j�p�qp�׶����*��QmpT2��כQv���	J���4���E�h�^Tl���(��i]86k�����a�{�E̚���T&�rIp��T�A�h)UQcC�q�`��E��-��VTEkDDEAEb#YYQH�	l��`�ܸ26ɉ1���`�EE���U�"��H��QQ4�Յ�������T�#(�(���t�F��DUV"��c
�EF�TQ+�kh�+)l�& b
,U�������F��TkPPDUTX$PSEVEUX��S,��1Q[JŌdbV,�`�*�E4�X�UT���5̪��*$UPY�hX�X�����dEM%X��bD��*�F*��Ac ���V*�+�U�
(j�X0�(��,� �r�գ�"bE�*�V�,TT�(���#Xc\J���T
�bԬSU*0�@G�A#�#�A�I����ܕ1z�����-���yju��<t<mkj%�sZ\�q}������S08��|�e���I�lUy]H(�Ia���]Jr���?z��[�p�6���CG$������c׀�$�JG:yU�r���y��v��Ϲ��4��h��N�uz�x���=�u���ʘi;';Eb�M���qlv{��Gfi����e���T�,J��3oj�F{��m�b���;}���L=:8�������}��C�����9�б�Z��y*h,n�b�]S�yw�V���ھio`I�M%m��˜����,ؚ+�8�3�]����X��onJ�纹��׳I��m{X(���v,
{g�.���]�[i���1���wwr#���@�9"���t����Dc��ڶ�V���Bz��̋��oU���m>T�����Z�_ra-j;*I���F�����q�wy^ڨ���k\$��0�+۳%tpWn�N�F�N���U2Ͳ�$�5C��n��v,e��c���b�hӐ^��s�7S��yҡdW>�h�Ew]Xuw�/hZ:pD{.d��g���(�G���_AN ��^"�t��p��H�0��z��K��e2�p�(�s�&L�����=&fg^C(�j�!A7�vĔ��[��]�0�F�؆椰rO�T��
j���o�9 �B
'��~�YS��幖ӱ=�2�^��wj��Ŭ�-�}a�;�����dJu9��v�Q�g'q������ڝ�]~��΃�>�V�4����yGy�W����0�]��c���ܑy֍�v�1A�4��7W�]]gioZ�Ż9����%vJ^T0��
Irt��i��b���t��ťf��s��0�6V�d�3�͎�ӘUպ�Ź���&��U9S�W+�/�報{�iiz{*��_�����0w5�R��s�aT�]'U�6�f_g>G��0����x˰�il��g*��$pyX)1;\�]F�u�V^����Պw]c�u]ײ���v��a�˜����^lv�9@�M�eA�aK_�칧B�@7Z�^��hv�`:�2�O�;O�Cpm]���d�ܳ��c3��wi�YP��}Ñ|�%��N�}P�fԜn��f�v�-��p!���f9ӓ#n��6�r�R�A̫�$Y��! �=��Iit��Ѿڶ�a��A鋦5�Cq�~T�ؖ�e2�b�d��xm`����䶭Q{�CrC�Ԅ���R��Sx:KW��8���*������̛}K�Od���r�(>4�J/��RE�]Z�e�r[�ʬ���[W��	5����R�8��ݬ(&�o��L��j��MU4�zmo8Y��u�W��UXM"9�#��R�^]�]�z�7�GG6δo�+Q��f-�S$F.w����u`��=�~�rBp0 �R�,d�nk��`�c�q��$^2(9 ���(׺����;wJn��=�K�&te���w�dq#�����;��(GlP�&���99.�©fYGw�UU��gB�47S]��d�n���ѱ���:�s�m����#iΒ������}�S�sODlh������1y��oz_W�ebYC��v��XBϫ��5����&zo�u��^��G�cm]1*�C;.Jݶx�o�e����̣���p�]�hr���zZy{Dz�0?n�0���"�A>��h�W��ug���+��[����UX��O���p���{�Y�Qa2��z���<є}�IY���U��l3�������Fk����6��m$sO�0��z{�ɭbF�xR���=�U��[r�`�~��o±Uլ���;Xo.�����f����Cd��x��8e�����d��U�UM���j���]���S�+6�y�s;aSfwö���x��oC�e7b��즬{e��l�mDDX�Fn���15=5�[ݼM};���5u�h�B��}}JgE�.���m�ui%����n���i�Zn{'mtH7+҃�C0�c=w����K��|�����'\5�W�8�8�ջr�X�ი���0�nmb��N��k�8�)�~���9��˿��&��}��\��R����������������ܴH��Z�T��Uc��'��.=��Y\��!?&ELΎ���[k������d�2��+4F�Z��)���ӌV��f�O.0
��%�/w#�]b��u>�Ru�{/YG�����.�n���@�b��6�i� ;a;@=8E���_Q݊��jΘz���h���{*���#�S��b�q�����G�����j�>F�c\k�~����tً�q%�5{g3��j�}}bL��!(xr�١�q��n��]�8kE��/���n��9s�z�h�D=�G)����>�^�����͕�
��	E.SO���K��ބ]�\R��u4C�<j��UJ��K��ݴ��n(2?j{¯3N�u���C�1A�4��G$�]L=���l*K�E�^���#�����R��2����߫����ZӴ��V�����M�s���U'�EA�V��*q蛵��[���@��u-�в&�휖)ܞ%���e��f�r�Y�}�_��:��;��JM;�e����\�]��[ս�>����;.�y2��dYS,-�=ʛkk廯%�v6i�	��'��vn�O'o+�*V{g0�u�/3� ��رJؘ��&8"��[����,/+�ûק�.�����lv�m�A8���pg��}�;��P�
�ӑ�윝�����e�'�$ݮW|��L��Z�c�k��^覃ښ��טD�;�!,z�s:@o������
�o�N�V+�ݔ���o=�M���4�s��p�N�x߻:g��\}kTx��+�(G#�a�1%tPR�|Sx:KW�}����V�daM���\l�ؾRww�]��!�>�bJQGy��]\U��&�X/�z�N�aH��C-{�l���?��Po�[{vh�}t�jD']�&k���6U�;���G\��{��^��{��u�8
:��js�e��KX-+� �F^_Xl��((���#Z�`Y��w�}�9�L:CV��KI��w�8�\�SU��ñ�W(8C��q����ɖ���7�'��%oOx��~��q+y4�9�62�6�C�uj/7kku"T����:%b�
��3��(�����W�jgْ��8�i��Tg�9�I�*W�R�C���{3��v����2������(���j�e�Y^E.d{����y���r�❮����+�M0#���c(֜�U�	e���$�Zç��	�f`�uo\V�")���L��U��v^W@���yCR /2S���U�K��ף-�w�&���^��+ð�#�@�f�:��NaV*��[l]l��c�Z#�f�\��Z�6e���/Oa���Dq�����3;b3�=��=���>�ʞ��p�D�v��x˰�i����j��"G�I�_��T`*�^��rT��k��5��]R�,.�j-�tיM�u�g']�l���p0�ʩ�;�b���c�Ʊ�mr>��Ķ��7zݻ� ��Y�SOyO+{y�.V᭮[�Cr���C}=�p�)��(7ݶ$w3����LPưn1x��K�=��6$��(>�/��<�s3��P^c���v^sس��٪��i�	/kQ�Z�B�F2wϪP\}Tݩ����{ԣ�u��[���!����V�S:��K�·�{�yz��]f�G Dv+�O��j�o�Y^�����[]�-+�/Q	�+�HN��U��#=��oM�կl��ңވc=%�Y�W�f }2 ��U�@��Cĝy�u7�d���(�M����j���������O����5P���}6,��t�[Y ]r-����2)y�e*LZY��#x[]ssYd)�{��e��*��h�w�e�*>:�4�m�D�5�QϬsJ�x�a��g�1ة[�����NnjwdC�N��BU#q(3�o�u�����cP���&��te쑮5·ƂϽ���ܖ�ۣ}֌E�VC=�T���n�V=Of���篹��_qT���Dlh�Wcʼ�6Ll�ʋ��y��9��b�i�6�ؾz�m�<єZ9'Y�WQ鴫��G��޶oZ�m��j{Ř��Jf�������==�ޝ�#�ce�M�3�x�Rd��~ړ[)�+/��5}�7�K|��ԯ.k�Fӳ�Sp�t4���,�R�u�s�/o0{��^���M�]͗M�a���ǝ9����g3��t,CI�W����{���q����n_�6X���|�gI/6�=S��g�s�sÒ�Y�#.hN!E���'������ڀ���r�-��p�r��-����Q��G���5�RA�ka�\�?:�s�:��t�/N)m5t��t�͉��v�7<�S���m��Zu��{8�O[�Ωɦtvm�hh�$&�q��"6Uee��u��AwjGnLC��\�9��g�B�ޓ�&<f�y�jưQ	�����sB�������pN5h�b����9z�Fo:t����غ8�&��^K�؝�{Y��;���>�X��*�(���������	�}�lq��z�	��p"V�⣹�^).O{�K*�������U����v�����������#r�*��KD����kӈ���ƨ�ӓY&z�0`}3QXOO6!�V������N
�ʤkg�:N#��qc��}�x�����K05C;c\3֚'�Ն��S^N��{ӽ�n��	�Z�k�.����l"�D���SBވ���<��W�c�L|����ifi�kx�sw�H�h쥊8$���V��ʇ6K^T*�f�`��
���J�,*��:3�W���sYe�;cäX&��u�Aw��[�ƙ�W�3��2��ܝ׎���VE��"U)5Ce\o6��Ot�����7s0�����j�f�@���9jt�(�ֺ��%��\MHL��a�n���ha����}�fL�[��:=�+�q�3��;�Q�y��乄�jr֦���J��:��NaWX��^g�w0�R���\�Ii�駙q��o-5�X͡�pv_�j�����]�y���v�yҤ]�{)j[�"�4v� 7�b�B�jW�R�젳�U9@&����-e�k��R�
PKbZ��v�e�vny�ҳcE�"	N�F�G>��>�JDs��G����Ķ��7~�
)��:���^�pz����b�N�~�'wi	+��u�7�7�M-`�>���'V�����9I8l{�mܧP���1>(��}k��*�v]�j��T�Gor�k��C8��R���=0I��[{v{0�<t���ŕ}��w�)�T��~�'����J
}�]BC�@�܁"/f�7�ëMnT���w��bNƫ��i]Y|�����H 'P�v����6v
f���W�V�oN�)��`�3}�su�k�)���[[�]��v��K�u��::,e8����/SV��Q5�u��fs��aj��a�
���+�lV	y����Vcxjwj���Tqd�T�ޒ����M���DV75Q�t�h�:�U��� ��f�����#����:�ީS0v�يWN[ؙ�lJX�L����ȴTUj��M�f����� ����gn�p��[R�����A�V��i!B>����$�P�{���0-�I�7���u%�q-Q�xgi���:e���g>VWE����0��eZP]H�t�5�4�6�#B����s�3"�H��Y���"}w��[�S��/S�(ŲS��}:�VNxR~����8�Rw�p:e���j�RW��[]J�eh*Le]�:�t��;�on�t�_8N�<ւ�P*�3�F�]έ>@x��N��G����N'1����EF�L�DP��tƆ�ã��A͵�e�k.inN.Br�N�PlX��6)7%`u��Y֝�燲��kzr�[e���-Y=�z��n��d\��s�f��1�Y���έ6�c�JfV]��ct�BS�m>�Ӆwf�vk��MG�LR���sLa�]�k����uu��n`�c���wLp�3�L�����nڎ������i�(}�]^@igKub���YZA�F۶4r�a;NS�3qV���(1@Q����^�b6���	��hE#Csevۀ0�MMW�&V���T}3��i�:
�w7:�E;�K|'&�mK��8�q�Z�%dw�s�凚r�Sxu�Ok;��GrW7C���u9u��W�b�Y�=�	}Ѥ�7=ᯔ;�����,k5)(.(ԵZuQA�K5x[�f��c�ꮶg)�����zRN�8�F��vf�F%%��'c����HWS8r�,>+o+�[����$�M��8`��9��9��r�Wx���ʜ�o� :������'�ps�ō�R1Fs�_Vc=��r�vT떄����lW�i�(�h�����j���Gr��WA=������[ge�\{�`�]�\:��6Ő5�yG+�1;9�Qn�GGP��D�:��Zz���ݦ�u=�zN��v�eQb�:��6�R%��ܴ��v��N,��u���鮨F�*q�gZ`�i��S'θս8�Jy��wr�{[o�;Ž��p�𩢳.(�����H��ݦtu+Z�s
6�FԳ*�	���6*Y�
���9s��g��qn*9L���|�Y�%�U;GiA�ws��)n@���nF��`�y]_![��Cn���VuV7E�G@�d��l<��t1Csh���dd�y,�E*:U.\��i�|��;�U�X/�c���;9-"�fp�zމ�����;����wG:�ĺ�Tv��@�����Gw�=׺�<}^��eS��i؛sd�~�`�?R�(z�U*�*�Ȱ���d%`�,���(EU"���TX.2�+��DAUEX���X",�QPXċEb�UF5�X��()1DE�MQQc��*��Q��TQT"��4b#,�R�U�"�c(.�� ��,b���(�*PQ`���M$.��#�I�UKj2�R���U�j�F(�
��E�",F(��E�*,X�EFm�UPGmX�ETEU�IX*ň��Ҋ��;eլ�@�D`�(�"�*�(���)dDEDQ����X&6�TUUDX,3,Ȋ����q(��"1bZQ��Eb�%�b�*�h"���ݠ��5Q*TQQV�h[DEH�B���PKJ��PX&���V�bZX�Y�WN+<����Ua���Nlc�!7.�*8��L�6oX���0����ξ�n��b�}oC�Cw�F�;�v���Y�mmgQ�DF��S#{�{Tq����x�O���`C��r��V�P��}�W9kV�Z���gD�r:�Mn6�B.������C@�7Q}Y��mUUf�c������j����1���~���cr@��F�;w��EfiQ���5�����6�Icq|�J�J\�a���.e?�g* ѕ����WO;[���v�|ۗ��s��u:�uʭ��d�����K��i��Hn�	�b5�����c&YU�W�`���glKӺ�+�Ɇ�eQ���r_�Xe�.��n���]�T����Yv���P�}�<+Z�~����X�]S�(.�E�Yw�S.s�y������j݈��Nr��bh<�p�Br���vRW�M�4ݍn���s6���b��4�Jx�B��Cr�>N]�z��ͩܣpr��7�ճW��UP��9ɾ9r�(Ndr��왮�t�MZXր���FkB����յ�;q�����ru׉��¸+�m��i�+HX+�����F�_oIڨ��J�gX�MG�;�HG%�dn�̡Ӆu�$9����aX)�9�%|���|��X��d������A՝��KݎX�(3��R̓����j���֣�>�`B�Gђޘ:�*����jA���o��	�����mU3��&�簈��%*�`#ՕΰU�1�V�p7��=ȼg�N��F�.�mu4�"��ⱬ�r/�d�����q�=KsZ̀�FϷ��5����q�j�z��kD�3�h�4:)j�U�˝�8��j��q����F��qM��B�7�����s��ŭ�B�^N2
��a?F��
��+rc��r��5'JG7c/�+Zp�jv�s�{a���3��N�{�z#z20�gn؃�u�ַu����s�V�u*7�hޢ��p��h�!����C��eu,*�_��<�^t�$8V4��O}�4ߩ�x�-/Oa{Y5�1%(5}r�oqĶw,D�.�
�m![\��A[�:�F$��ӻ9�W���s�U�U�qY�[�8��[��:Ê���r����H�`�r<�"�"j�}�g��WV��c�7�����	]�$R˗����F�v�;�'[��O��B##�i�	ƞ���Ӗ_���{�u�����A��k����_]G���M��i�֪��=�ڣ�1<&1�Üⵔ���{~���k�oq3ܐ�fi~~����9ϓ��X�;�����u������x�3O�wv�مm�ھIo`K�{��v�n3�=�ɪ^x�Ǳ��q����ʪZǗVk9�	��W���NNqM�M5c��D&��K��]��d5�vY�n�A|�q�09M��w��_�Yixs�>�-�v�丮Gc��7��2�|��0*��T�(��$|���~���]��9��2������ʯ�X���0:Gy�	a"*���H��V�j����lDgj�x,޽����$�����G$��J�3�N"Dk�͇�Vg;���ںY��G,x�����y|݈��(!^�CQ�ʟ_c�����Y�#����5�lWl�!�Es�y[v�n\��y�f]�y%x���T�YYV:�.�l�屽�5��OL��9r�gt�4f�$ޢ�zٛ��� �mA�0�5+���(9�SxnL���룂�E*�Z�b�q�G���Q�z���bJ��8��T3֚&Z��"9L��]���[&F�����tw���t6A]4{mX�˽qK�:�ж���3��-UH�n�ޥ�ڷ��7B��k��^P�nH��F���SI���cn6�\:�I������I�s, ��u��nNf�-�f�f����F9�!��i�)�%�7!�T��L�^���ӘU��Sv��qlr��sE�7:#�ݼ���\�.�
io>+���Dq���R��U���H.w7��v5�0�sK8e��ka������oc�٣y�++i84�qm��ݧ���j�9�
�WU�~�A+٦�&˿2�����k�f����yH�E�9�Gr8'# �����vRV6i��-�`���9Qu�9j���~�{=Ο7��Ox7(nP����BA]u� _����X+{����D꜠ξf�9�`�ǣxv�j��dV9V���
�!���n�K ��:��Y-���,�om�S�ىhܥ:v�k�P�C�i�Lх��%�٫E"p�@�lfn�FWeof1gYt�x�g�V>��x�J|/x��P�jq�^����Y����\!w�c���A�Ă��;}k�7�X�we3AM�0�t�_/Ru���"�#�q�7ϨJ	U:�"����wzܧY��]�ζ��}ʬ�S�G\�
}�]BC䙞���ȂM�cݳӮ����+I��ƫ��ZWW��y}c��+{�C��9v��l�Ȃ���:I/t(��/\�`�#_;�wW3�Ţe��p�A�Tt.Q��h{��2!D��Mnu�GT�=���(E޸�ɢ����׸B3�[��6�����]��M<V^P�nM�Z65;}����H�wׅ����K�8?S��ր����4Ǝlw�n��&:��/��%$���XL�,z�m�<;��Gg�,��ƌ���w���!;M'�3of��q��m攇gs��)�/Oa�=��k�뮥��:[|���$>�,d��'o��bkwI�-���;���6m�t��m�V'�٢�KE�Ҳr�ʎ��ژ%ou�w�H�X|�t��
7t`�HՍNu�.]m��������F��Y��ଛ6�/�J;����Js!J��'*��t��F�e���;Xd���=�Ҵ����QR�ܺ�T�t�����$��čO*�eX�U�}���T��I���NҊ��k�	�ͣ��)=c�/Uz&lh���o�O#��J��M�٦�,bfr-�]�����5�[ݼ\��mu��47 6:P�_3�}Jr��"���.�$��RnKw�`�1�W�K�=����r�(>>��q.��%�[��5ݜ�n+7���cU�c�H��G��\+�Dd�|�S�Uu����-�]׎`r��'�P;��-U3�Oɥ�avvڑ(�VҠ���r_���noxy}\�6�vĴLor�Z�i]X/Q�{���NF��u*�&1<��M܆-@�h��%Z�'1���}|Ҵ�@�\zt�nf^���Zm���v��Bp-�T$n)�)�����b$��I'�^�g��D��*?I˓6X�ǝ�n%��jA�+�T�kw؍8��]�͎�+�)aά{{��W�st�#�Q�Q3II4��Ոof�_@�V�z�R�[gDO��,�v_u������e2��;08�%}�u�R���=~mP��v���ۯz�\(���ٍ:X�O!��仔�E�����M ���]��%vd��q�P��e����8�W����7�l��c�1�6�h�j�~�������><_F箺e�	Hj�71����u�G<`���==�'�ګX�y6�:�y�I�5���*��w6�rv�מaUB��<�zhv`������o	9
���7�;bW,�Y�'S���~�ArrCoy6OkEI���9�>�{�|��б
v2�rVv|{��3mw��̙x����rKwn���6�-S>s�����Vv>�)��W�������<e�R��Ǥ�Պ���Ⱦ�'m�KHk�i�>�k���gr��g��N'������tYԦ�����k������n7{�blc�����'����%����o-_i��. 91[|U_^F�tVi� �7���xV/O��P�K��D�]�̄N��iL�a׉�J5|4���L��;ɝ͂�]�H[���
/"|�+���+PyHiLa�j#q��9����S�~��y���=;V���&����C���h���¾�d�c�ݹ!}R�#��K*����rq|}ٖ�n��`!$�ZR�bԹ,�WL�r{k��䐔	�
}�J�����kӈ���sݨt�V���w���~Ά��4���f^_7b4'9o�kr+���k�ƲP��Vb����Q�oT3�D�-Xv;^�S�DF��@���.F-��{���_�}��9��XN�4-�C=Y�]wZoa^���LҒ6_�gT��'.۞��GU7����{�ӬA��CAa�Ш߸�K=�Pړ:�d�����.e?io���M���δ��M.�TU��ؓ�GV;�ۚs
�e?�\2��Wh�o���B� �fa5�ϊ�a����.�r�p�]^6H-�ܯF����\Ŕ���3(Vʞ�RG]��QmU����9���s����.����%W�%����Y��]<�M]$VO.k�RSO�<t�DX��9�^k�^��u�5������W\�b:�m������N)��z���^����g9v��vB10��M��ޭ��f��pyt&/ *n陽�̽0���7Z�;}uK�l����j�e�O��f�mt���a�b{<�fV��<=��U����r�;)+4���MްQM=��;9����pn�w9)+a����hnT��BA]Z��7���=p:EL3��U�qm`�7ИM[�=��6'Æ��e0R�;�`^��틁�R�Ѻ��:���J�	kQݏ�O��C,o�T���uu6hk�}��q�;������U-�Y���P1=�̗)B86\+�R��v�#m�exJd������Һ�˄�����8�o.�9�L�;+l�߽=z��y���)���ϻ]�;cW;XD�K��(�]�&ut�#�2�jYdC �	�ѡ+����T��n�����=҃�x������S�g�ʔ�ҏXgZ��|^L�`�����zi�jh-�m��d��v`�ϓ��1�5(�x�ᔱ��S�����:�Ԩ ӂ,ǽ/���v$�R�����0^̘��*Ӣ�Yg���IY�Ph�}��F�u>�R�Y:��}X�\y��y�Mly�h�?S�Xe�g"�(ъ%��U�{1�7�h�A�.*��c���y�ٳe��01���:O��xZ�M[rs�I�*h7��Թʫ+��=���Zǉ�67KB����øm��y���c��sq6�},p��{;�U�f,њS��}��Mi�݋O�c6����e��!W��7���P3��9�g'r��A��0�h�G��Vn�����Wnb﷞�ڧ�ȝ+*�eجUuO�[ڋw笰7��μ�V��xx��3��z��&���o��A��48��܎͵7
�=�xS��b�I����\���޵a��s��U�y9��j�ި��o��9B�޽Ӧ��\�e�Ϣ�Z�G��+�؈u;����辕�/��z��{�q��\v��}yU���7������\�]7�������$��H@���$ I?���$�$�	'�!$ I?�	!I�$�	'�!$ I?�H@��	!I��$�	'��$ I9H@�XB��H@�XB����$����$��$�	'��$ I?�	!I�	!I���e5�6�	P���!�?���}�����9B��� ��AB�)P�d �"J *�J�RIJ�u�*@"���uJIRUT�T�!J�����h`� �Sjl�#6�!%�V�L�f���m6���TJ8f��V��U�lm5�[Y��2�QTp�l͕�1�٢���2-�-�n  �  f  s���H8۷Mh�T��eQ�f���YbJՍVj
*E����e����Z����-	P�b͚ma)%M7 r�aa������m�5Y*3V��6�aT ��d՛D����36f&��e��f�Q�Q$ r�hm+`��X�XN�p���w"m;a���B�(��f�GN��A֒' �@��4Uk�l:�\�B�l�	R����j��A���F�Ԝ� d�v�-:[8�ˡ�L��    ���T��        �x`�)S�CbhCC&M4�  挘� ���F	� ���T� �h�����挘� ���F	� �i!�	�#I�&��5G�ѡ�hbbO���/��5��_�s�Ξ�+�u��[Ϯ:?.�D�� ����K!5� }������J4H������hh?ќB+&� �D�u� ��d?�@�N!��|���7��������@ �FNo������f�����-nu�e(�����~_���g׳U�-�{���L���&l�z��ͫ�c�j^ּ{����^�O����i��R�x�/^2�KyA^G�2^�d�&
OicB֫z8���<���v�F�㱋-gZDe�ޕ�{[�4�KH�PO(e[�ب�0ݩ�v����H8�:���Y��;yr��u�r�%#�wv��2h��dKc�4ԡ-V={�+$�$uj��L����1=ki��)*��#F�2��3�j�]fU��BՖ��1�C���\W4tX�˲�6�k��P��3v�&%�J�Q�ю���˭����	�I[�������2�S7^���߱S�MU|wm(��ԪBQ{��O�´U�*�o�8ްUF�]�B�z�S#Y�i�6�oq$ѭ�V��k����7#W`�6L���0���K'1F�bL���Jd��E�PK��x&�m�a�6!K5��T�W0c�"%[�1�T/�k6�m�KK���*�k���Q�KN�u�f3���(7&�T�&%ݲ�^�QH*��
ݔ���D��f���O��[9���m^]>u{��1M� ��v�����l��" p�!��Q�ڦNgt���N7��]OR�����XDRN�7G��YJ�tY�
�Te�u��ߒq��n��Xssn�Ʒj��
��'#�GU�ͧ���MOm4��(������-Q��!��m�6����9Fi�J�R�&�Ou!���yl?��2ͳs+n�����v�(J�h�mvv�5&E�����Ά�].$/��Gm��zYA����7�oU�*M����B�����E.�BT�z��� �)��U{��kQ9L0q9��䧭�<@�,���2�gk8��QN��h֚�-Q�1Li�Y�����E��5Ua�
˕��%��u�kumk(57h�ϙ*Sw���0�8��b6쵊���y+tVL(M�����K��s�^`]�dJv������5@�R�6�"V��CE�J;�K��V�Q�1*l�)�b�����Kn��w���)v���u�Q�e,���&��2���utEim�5�i�T�T�n�e]h�u��d%	��ux3&�e3���i@�gi�;��^m왉ҎƐ��4���tTz[�!�����������Uְ֊�6�D�e�;p�;�s6��V���*���0���a"R0���[Ol"M@aÑ��`��g�S찙V-�<��.����TN��Y
��������E������R�>�P��*RM�A�z���6*��u��gN�r��t��'����E��/K��-���CE�Ǯ�MlH���n�d�a��m33�ͳ�{E���4tǉ��Ik��D��ةY�C���� �i��/]X[r��u�4�̼ڲ�lk/d���6���Gc�;��ۣ�vl��u���SI5��Q�Ɗ����ٶpᬥTYVj�k܅^�"�^j����E�֜ܕ+4�Q�:kۛX�;�a�u��ʙ��I:�k,�.�E��mE$��!����f�F�<�Wt�����oqX�Q���B�ǵ#��7j��0��]1WU-XuuTR�V�f)`:V�rV�{-Uʼ|��W�)fb��nR|�����9����svT���UV��c/5����J�B�d�W)AHL+	���M�+�n(3(ňP�����U�����V\��Z�V�DU�i� �'�HX{���`#*k�[���P9+%�)�~�mnPTb�m��ٯ3�N�ňbZSL$PF�0h��h��[yy��
Ϋd��kmk�n�Iڤ�.V��1�f���k�Z�EM7T�ݢ�V�0!���W�OP�u�v�3B��,"�1@��,'37K��V�׷�����{�J�.��1�n���ܬ7u���*9W�.F�k�ڽWVa�����6�F��q:x-0���d;Z^�x��T��@�e�UR���D�&���Gu����fY4�1:�Q���uQ���	.Ci��M�#6�M���)+B�Ǎ�9�z��6��-��
�8�Me3J�k~�*�_�1C�f��i�KT�;[gF6+��-;E��T��Ռ�*�Ϲ���*_d��@�.�R��^Qr�Y�1�e��B�\uj���+.Xd:�2�N�z���*��X�]r9�����է�L<���s3Lj�Y�]�D���;����U��hY�WMf�D�fK���l�b�V�^#l�-]m�V��9�re<�*'Ih������ų&clԦ�yN�߳Uq!�%�vOv��/�QڽH�J�"�ª�ڂ˹w��f�A���p�Y�W�I4�*�bUx�՜�p_:Ѭӕ�HB��^Ԑƍ�8D���-��-�1$�������RjIdA�n��ܹ�\N$�ʛ�*b:.��m���yJfK�!��5�Y��U�d����j���ޡB�^V�(���Kw]��4��;�P�7/�b}��I�+�UJ���Fu�u)�F��@ؚ)�ڢmRnK��SP��M���|�i��Wȑ`�|��Ի��S��[�U�T�VIA]�)f�/*�f�2�o�t�'I㢐|(��;t���p<0ռ-�,�.��;���%����x)����ω��9��������=��uɠ� ���W�H}�x6��kn��yPb�l*�UN��7��]�a��t�0VȪ�Wj`lS�rUV�'-16�]�X���"�5�7Z7,=�L�������R"[�K��o�ЪuL����Z&\��#w��a5�E�_E�
&f�%�1:�4�U��;{ZN�5��hG@�;u��Gg+��i�5����?~G�o�'�}o]�է�A�|4u3Z��u�u����wO���o�&�%��:� �5�r��	�)P2[���M.�ȡ쨥]Z�2�+ܭ�{��޼�z̸m9�ϸԲGa�E��w��u��.�5Lv8�mn��$�i��i�����Zc�2^ک$N�����U�
��q.o�h��Iɽ�<Jr��Q����C51�A����p�颎�S51��纵&NY��V8�lK1u^��v�����[�w�	�"L�\�G)#c:ņ����{s��d|VM熫�Uթo�̭�H_��������4��D���R�̴�ܒJ���K�C�gEѺE=�E
U1g2.m+]�vQ��S"�?b�W��j�{щ�X��Ж�	�9'�)s��c�Q�����Y��#V3N���J��k&��MG�����Ni�r<�+�[�u6�������܊��I����"^=er��R��t�E��/�jA����6�S��!�vN����@
�S( �#X��6��%�P��fV�[�)�j��ط��\�;���̕x��`�7W��5Lw`����X�p�PB���j�'4վՀ�Qo�{O'�v#w+��\=��lnD���8y:z�1���Wfj��ύ�pm<=�J�����	��8e��EQ)�J�+s[*���N�G�Y�A��c�L�+�̨�Ik�g8Z�M�.��Z�q�or�N�9;v�`��h�pCF�`W�l0��x�C��l5�k����G#YQJ8�aO!��2�Q����=|�}(u�`뤸���N�4{��'E��$�W;���ndpv�(RC�]A3�J�o$*�c�6�t��#j�UX�4K��]��i$�9�#tE)��;��6����\rV���S{���δ�տ]]W�t��t�:���aV>�z�Y���w�������c-�ys|��l�I*��͙����5hW���]�(�kg_ �KcJ�g^+��.���[�ȵ.��Eڷ�q�m��o�Z�([�h�|M�$+igL��r$���}e�g�:�!��p�w}[!���P/&c��[lnr�>�һ�7|+h�.�U��H�c�G�W\s�ٻ���v�����d���C G+]j{\3����N!�V��|9�X�r�g+P�ȇ%����zuy5����Y��*�h��ʧbئ�^(c:�WRe]��.���Щ{}��/<r��M^�+s{V�(�j^��Z5T�ɽ["JA�|����������]�����ϜtR}�ud��G���.�p��V��	4��"�d�Q���XV���s�`Q˪B�U�n)�A�g���;�]�q�i*��;VzZ�L�5�]�jE���:�ǜ�ei��i������o-Z�č�K]d75�(��^�2���
�v�x+�1)��n`�i���S�^��G9!�-�� {��W�R��o�L^�ѻ\݂���a��L3v�o��5Z0Y�71,��ٵi.�/���e�Z����D�QJ����-{G�ʽ]�33��yٛ�2�8������V���rW `M�1V�:2󢽥�q,��d^�B����Lm�o{fj�\��d���n��YN�v-���)R�:nE5�Z�[thAlp�Uk���h�/��[s��U�f8y�i�ǹҮ<�efb7����Q��:&�7Z�^S�FeL{��������Oo,�ohDm��TY�d,P���t�×�ww]g+�vծ�G4E.�1�#Ju1k��]�P�%���y�w��&�V�}2k�̺.�;`�tK\ Lt��:�u�a�C��88��a!Eԭcd�yY�wLt,�£b]�AP���DF�����Ai�1Q�0��-�5o`�\8�P5ie�����qH�s�op)N���e�1��^-���@�_�ٗ�\4H�7��L.ICO��ɭgD9Z�ڽ��LUʺ���2e��e�u��4�ű�,�t�[�-��,@��XU9H����ܥ��*5�9vh���nS�kh��L���wr����zs���J���d���8�T��	�E��Uvlѻ{t�����8�3����[��t�Ӆ���:N�h�m�!ju����M9]v�u��������]],����G�	��R��(ѻg�ٛ4Vc��szru��%�;GY��v��[[�!�e��'Ӯ�:	�g�o��'/��!��p�0�S�ޤVTs�-E[{B�w�lޣSn��i��WLo�w$���Qk�FB�����i�&�@�n��gQ[bI2V.�a�g:뛈�F��`(_v��㬹�x�� ���ъ���E��RI�tf'�9��Mʧײ�wnH;Re�u��ܒ5���&��8�w������c�3�x�<�O1��јHUڔ%��ʛٰ���Y�a��0��b}�r�@"��	��n:J�YY�x=������U�Mbu�.�Q��Y5�f ���O-UWgN�r�EJ
Z�����+��L-��)�6�:#6;v�-�$�E$�9$��$�6��|�Ȇm�y,����v�VF�x(̹3C��ӧ!�]g.��ys����y
�K��¶�Gy�U��U(��pf�}�8r�:7��i�-]�q��r��w(���gQ!Qgt۩Q^Ԣ{;����%��Sw���d�\7`�� ��o����1u�͠�-�y`n�a�3f��j�uy(L!��x3Gp{Kv���u#�Z�̡p���,�2if��
��iJ�ɛ�TZ69;���e�W�d�N��ݲV^���4��lv���M�uB1����'���.�n�SoQ��'l�>���_3;�w����u���^����@|�y��r>s���'����� ����u����dUPOg�Q��h{�.k-YX�p��̜�x��W��F��4�v�	��u����J[������;�$%��-���81�˨�2�E�0��u�/�Ԛ�DM�q�� �_M��ѽ;S��#��7��Ԉ_^��w��rLd�쵪��ohԠ�ZiGK�ܻ��{���|N(ɓ�]�.̛�u�񛮦�Y΃j��D�6V�.��(��`�0���@uV�SFa+�j�WM�{6e�]�Zђ�tgGF���!�v�ٽ��P���"�u���ө�ɦ0�%�-�ʸn:om�hWo]�q�֪/	��o.�2�m�[�>�.�cs�.<������iU����ds�j;�Wlm�9T^��%��EgC�v�_T(�ݺ�yk޹R�U��u%ו�]ں��qJK�ݮ���u��!���x'f���ԏ=p��J0r�zl�f�C)���nR����Ѭ�o�2z�2_#[`c��3)����uS\��5�6�f,��Ȼ�n�J'}�88�'�:�kC;SFXQ���W�I�Xً*�ʖ[]*8j�4�f=�>:�a��+<&����]ޭ���������Z�yt9n���>гK�����+�{WǄE�:ܭ.p�ze9o��1�ms����fT4F�I9(�C��y/ᅾ��&T�5��/i��'�b��v�!
̝u�����P�-��7�W+x�T؛�0���hOm���>ݡ<S�ⲥs��<wA]w���Sð��U_3o���AP��k*!�1yّJ��{);��S�6����������.����r�L1+�5P�g4-�K��$A3*m�̑k����;P�ҫ�o�d��ᒭV����T/��I�A29�r�_$�g�p��1��t]�{=��F:����:�s�(+����P�]�7��r�9[���tlޖ�Q!�ZC�@*�K�&ʆ�\�Zf:�"�C��u"9����wH#�x������o�-�\�Q�������t�S9Sg��r�o���v嗶+����w��iR����ʼ��j�����P�Ⱦ�������m�Opێ�-�k(����܇��:�y���K�K�x.Ebq'N�'Z7l��I�.��׻;��1���R�����>�%��<*N�oj���Lv ՎTخ����gU���p:���c�jV�"�N���</4T�e�:s��o�Tl�o�ql�&K�خ�_\|l*Hk5Y��bw/J�ُ5�U�&ɭݛ�����u���Qʬ��lH&�#P�V�wY���.�t,��wb�[��v�� �:��3s't���0=��=����É]e��x*ټ��a+&`;�Mfb�g,մ6_L5�6�]VJ�G�z�e�;�V5ձ%[�ύm%a�m���n�U>X�r𶡃n�PD�[w����y3+&��f�Yj�3��e�I�!���c˝ ����)$ő꣚�Ϻ��,��9�j��a��N5�P?P5���f<3��)-ϊ�7��"�|+*�\�e`�vH9+�T�9��μ�hegFpkW���(V�ٵni�� 6]d�jҫ}��]�z���i+UOE�\����Y�A��³����A�cn��]��@+�H�L�$�G,sx�죝U�kWlgoV�z��K�I>�lKj���wf��\�:�v��khU��M@�\��*|�5���mU]fcI+4~XaԶZ�_�v�nq��Kͨw���o���T����$�q�K�-64� <��f�;�^�ƕ�s�Ss(3U��i<�	��-��S^���Y�I�H&U� ZѩKv=y�6c�qJ��N��4��u�����ܣ49�M�5iS���t��A�5�a��Ӹt�%GJI,�.�pO��S)s�$���Mݎ͎�<�&Ӽ�Mr��N�yI��{�.V��G�C�&&jX9�ܹe��t�yu֣{w�I�e�t]����Zٲ������і����V�^N�#�)뫳���J�pD �mvuN���ؾk&D��Զ���@�٩U�^b�}f��[�v��--ɭ}�P����*Z�/��ߪ�ֹ����8�(�]�sfK�MΗFj��,z��d�!�9:(��ɒ���ڐ�Np�곕s!�j�rT�������]$J���:�qE��̝*�J	�Y7�7��'ۋ9%�nJ3%�x�G!�g@Fe8���8*��ux7\���@ʇ��cl�]�kle���O�9չD�0��H_;0�Q�Ջz�{]�x�ŊM��;�ы����{M^+a���LJ�d�Kd�[
�����M�טr�o0Ɩ����AHm��Ue�/'S�����&R�'2�H6`���q�ɮ�ۡj�*�YUٰ�;�-ܦZ��C�w���sE�	V]�S|��t��(�������D%c�Y�P�X���^Ef>�aظ􂓇j,���g�"�'d���uk.�����V[̲
��2a��5Gt���E4��U��8���j-��q���9>z'�&a��0�4��۬�m.x(�R��b7d�7L�@@�?�L��&S6%ء�t�2��M�v�3:��+U�1�l�t��� ��q�r\�&-ÙT0Qw��%��ԫO>xI?���E�9�bG�ư�)�f�fj�Jh��w0�;qّض7-Y�2���P�pM5`��yA�U�H��UZ��o9U@���XZ���ORTN]-cnл%�kSU�y��P����aTe$h��Π�\��"��C�eY��Ӯ�#gM�Jy²�>�ɔs�='�}  �D"�8󙒼�ꫫ���G��©Mϔ|�>��س�]f�B��ܻH�|G(��0��)�Y�y��0��Wb�����o]���"5���ˬ���0�n�{��コ��Ed���.���Z�Qݥ:W,ߎ�X�cQ��Lo�V��a�#��PQu`Ǜ�6IHS�x9+����X�Z�UkY�:�ZU��p���s%V�'0zO-u�(D-�b�n�vf��4��2��{Ҹv kF�p��a]+(��I!}:4s��r��}�'.f���əZG}��e!-k��,�����aZ5��G뿴U�]*�Q[[:´��2��TG+q�s1���-Y��έpZZ)�V��.�+[TYGV.V��3)�Zc�խL3��	sT0���%�`�w��ۦR��QLr�`��nR�6�.�s,(�Qmpʪ�Ԣ�6�1u�2�)�-�Z[Ki�\�q�iVffK��P�-
���r����Ir�R��."3��Z�@�c�*���-e��Z4pC�:�^��]�O]���Y��M��
�Ld�!|ԝu�}��o��b����w֏��7N����?V�e1��,�.:c$�w�b�C:Eu�F���:�O�ۉ���jjpN��^=P�Y�xE���B�=��/4X��|�v�D�,�Rj��<��3�'
��F���c]����Q�FQ"���Cw}�w�e#�i�/~���Ή�j�qA�>4�m�������.�O:�)���������%t7)n��Ӭ�R�H_Ef����-�Vsf�j$T^�9l�F�P}�5(�4�!�^{�X��xV�j��5p�������7�+�����7s�f���}�>������gz��d�^�l�E��sUUj;H�8n�)S�փ��O��,eC�zy��:�TO�f��o���#GK��^aL>6����{0�����>ؗ+uV��J�y���o����X����!���y�-`���8/���c<�C5Z����CSy�O�4��nw[��c��]�.\�"�,�(� �K:@��\ΠնI��<]��7�@�����}|�&��u|nD�O�e����,�����7��b(�܏Y��6m��;uY����{�)�,St���R�9�<�{��^	���E>�����*ڸ�JbV��Dg���3����8�V+��FT1����b��Zl��ǆMf���[����<*���o�
$�tC�7A�9Y��雛�!*�p���#�Q��a{���3m�L$���b���[W�a�H�]�p�	��}�";�����|�/�s�}؄<6�57�D�h|�ͼ4{�o7ljE���.�U���jАq�h�s�W�ʤ�	�U��I�R��V9�11��P��ץ�9_����G&6�kH�<m�dJu�F��ΰ����P�*�߅U���"��s�f�ln�;�G}%]I��XfѮ��oCNS�@�$tn�0�Ԡ���^�Ώ[�%$Y�%�>��T�י!5���Ԥl|����n�;��mxL�z��l�Ӷ8�=B��4ó�З)C��%�m�TeaN=��w��1��A)����O~�`x�<�/ ��Yw�� ����]� ��;����R-���D��n%#֬v�I�P&]�J%�j�>���!�];ɩ>Gf .H�Ӗ��y7&���Fj+�tUi�r�2��
1� ��|5Ϋx�W�!�	�Z��W�h���f�.�fC��O��n�m��P)����93-؃�9lg�_u�7�S��z��P�3ې+Εg>~H�c���^;������.j:B��k0�H7/x!d�T-^�]��(w�};U�Uf�Gs�o�9�������d����H��H���zW�:*�o5�M̭����La�sh4އg	Ku�ң��-��I~����y8b��!:����S��Z�L���'վe�߃�����b^^���.zXﷻ	�93;����s���G>U�+Ϫ;3��q�=��!�FH�-�̮�s+�mI�T��$%�BTV�x�pH���w`�#s�ս�ud�oU=���o���K����n�9�zvp$n�Ehw5Q�5�f�-�(��n��@��-_J��d�ng���>*Ǻ$��� ��Y�B�ɨ2䋺��{���ˇ����u�o����k׉��Ωj�vK�\Y��\�:qL���XE6�cYy}��Lߛ���km���bbsI�Uʧ�X�i5��q��+��'cz��Nz+�+rΖ�f��f�)~������x<�Szm-M��И�hB�Bn7!M|����{�DZ4+�>
���S#�����k:�]k�Y�M�#JȮ)�[��ئ�	��i)�+Cz���t�γfӫɽ)�f�v�2��D����A���\��|.��&1M'c�@���أ[%՗kp��t�5^�Hމ|�r]�3V7�<��I�#��:lM��J����$H:5/R�����wmL����"�l\Wq���
9)����C�}�r�]�k$;a��n��ާj���M90ol����"ǆ�g��̘j(�Y��Vk�9iɜ�$�������ҋ���mLpmo�u.��Qc}�]
sxEG��tƒ�$���5�4�0a�	МJ�Q;Y=����n�	u���U�'J��Q�ʆ���r�kb��|�u�n�m<�7��n���"����w��ݬg;�s�6�+���4�V����wyթ���(�>ʯ~��G:�Q�����Z￑䣫�F��yv��,5��r�Z)�¥�9�Rb!GF:��u�K_
<��"�w*X�BI;��Sw�]�������:�zփn�S�r��H�oLzA��|���;��\K�Ԡ0N�tk�Mq�����mկ����6�8�3��������oΰ=����1�4aYp^��J��x�|s��2�3��{�dJ.����wg'�+�`�ѩ�7�[�����B��F<=ں������a6�pH��q{ �k6��b�*vu���Nu�;b諍���D���K!����/�O������i��QꆺT����S��=L8˧���qM�t�y���uت�>,u:	�Dk6�����ZpJ�	����k/7��:9���EѽM�;��8쨢����r���?��Xof�q�n�u�ݡ��{�j�>�t*���Zn�%���sOX�,��$�v���hJ��Nv7Ԩ�X�i�)<�wƧP�8آ�뻷���5���ܾ�9�*�Eb8�'�w2�b r,A*(���|k�-˷�9 YٮVj��{V�щY�P�����V�ۈ�����5��uy�F�n�s!s0��4��"TZŨ֊%)���\�-j����ĭs.8�X�-�1D�A_�]Z��0�r�UQX(��X�((�X�-��E\k��UEQDV"���Fڱ�[ձSV�IY,EEU�X-�B�k
''�9��������{���o������r�K��$�^����Xgr��$:����-O&]�
����_��Ku��u��MU��5�C�"��?2�!ghg°��82�ꭓ|���nS�..��u�ǲ�J@�u���|�`��M_v`�ِ�F�sA��j�}ѽ^�,�2YIV�}��
�&hvv�
���&����JʷǷ���0�4#$`po)�4n��+�|�m��v 7{��)9�"0�Ɏ=Q�ȕ%���޺f����F*�c��x�	S}�{ N	7v����sT��SڈJ�uۥ{P��U�9J�7���)��L^�c�DϱUV�^}�/E��w���������5�|�g�oF�畟��t�1jDMG$��D��O7[~Բct{A:Aq``�8�ݛf9#'1��[�v��:�6�ٱ�x7��4[������n�9�n���N�,f�
��. �q3q�(,_����}9s��˳�~>R]���=�ԜJw~巪ˤ�f,5v������tJ2�*�kU䪝qI�X$8.�6��)���� �A�s�ݨ�Xe=鎑��2�݃�5��P��\��`oqߝrw[��rNn��8��Ztr+��ȷB%�;oY��η\����P� xK2���Cr�e
Y�Ҝ)Ұ�_������^��dP�����En���+T�JQŔ��O��U3�ju7�}�&��ҳh�&��h��������a�u��� �]FB�Qm\����	޷W%��p��4S@�Nt�ܭh@R����cX��q�)Z���$��a��q⨵��;�qAC���x!�VxKC��~����] ~�fD�+�-�~>���/_:�J�}�����=��=�\��9���������rj+"H1g\g�Ză5��E�%�A~ˋ��]�V���iۼ�zC-Q'V-	ә[�z����� ��/B���Q}U1���z�,0�/[�ܞڌ�V6�.����Y��3]m.RE=������(mח)����׍xyr��o�ʢ��ZX���s�m�z9#�'�����L�L�����KQ򿛵��>�FJ5Dq��pV�{ir�]e�3��?x�'��ռ�<����yL+U�{�"�i� $���?����[�}WH�jt<��3�[�;���>�S�#+�ǲuΛ܎�N�[���Eo�1M�G�g��G�gk}P=���0oT��3����ĠzPɋ��`���2X/��}�s��إ���Z��zj	أ�ՙ���Ɯ&�
��eur���t�KW�`t9vA�N�!c�y~H��6��x����~��&G�8�UMDY�z+8񐲺��956'p*J�`a~n�C{>ob�غV
�[X��#z�h��/	�FC���Z\� �ww4�0W-oN������^Y��qҡ�kh.~g�v'Q˹�O��C�Q������YT�Ȯv��p�'7;E�ll{�钖��S�����;���+a��L~��	ˏ�z��l�u�}�T'Ժ��K�u��*f?�@ƷW�*�o`���=�{0s����db��G9�� �fH�P	�]�;{��kѱl���D�,<�(Zw�m�ۛ�y�<���� >�v���L6��JD>���j@��7i=�$U@���eM�b�bv�ptQwD&��r0k\�-fwd;���5y�|�Į����n1�ڑ�^޹w�TK������v�VhJ���j0�K�G�/y5ͪq��Y��v���+̜�p���(����u8Jl�d�J��^�
��*97����]Z}���d��=�"m��t��Ƃ��ks��aꞨ�M����[qX�dOV���e����at*���$�u�w�E�7,���v�����m,bb�ݘl3U6��z��꼩�P�VnO�I�a%=�*�b�/E�Էj�t,N����I�'������4_����B���_�Օ\�h�/Mڑ����@�Wci6�����Y�SV�+�M�7�Zn�NPC��ƍv��\��o%:���{p��tY\q��խ������ūu���t�7[�;���ǈ��VN޶-y&��BWݗ^v��.�Mv5W��(��Q~1\�}	GŚ����,k'/���d�I!k�i��H5u�.'�����;K\�W-��kyp�~
��E�]�t�]y��1�P�T��2�G���v�z~�HP\ �{ ���>a����n�p5/_KMu���U�z�Ƹё1|9Qܼ˗�����x�ӣ��..��M��JF�^l�*;����w]%���Ut��'w���L=]ٿ���?U�讕�5pT7�_�� �HrAg'\��d�M*�vb��f�����8^w*xfk#�tJ����f�]e@��8dͺ��%&�h���E�)bh���>��E9�S�k+u,�&�u���O�����Ƅ�#29݂�3��|N7һ�9t�SՅi1ޟ�:�\���^ x3'�����o��c�Bi���p�K)ъ�+��a��7'v����
�b��Y��mn
w�<&��1%p��`!Xʉ����n�vX�d�]����:��jgJ�v5�C�D~�'w5J'���{/M=�r�[%i}�mJԖ��[T�$k��Nd���kj�M<�9dŪF��o�oCx��oh��.LWv��L�'	3��
4�3���n�+/�s�fVBq�n@��F^mJ�ʀ%:��
Dv��7+6�ܧY 9:!�	�C9�o�6����|�ν>A�t�{�UdJ6��ԣ*��V�X���+Q�jF6�VҢ�ũ(T�����(��(�
�E�#�UE2�r�� ���Z��H�X�Ub�B�+*˙�(�\J1�"�AkUYJ����8��c�޾�3�Ӯ���~��o�]��!c�!;NX�Qr)�i���'�����{\V�}���zx�Q�*���C]"޼��7� �S邼b�WghܳkFt�ύe������n9��yW�k�����'�TP�`��=n�x�%�~��a{/2 &��P��-��r������X��T2�k����n���*��!sGm�'Q��N��=��5\_�>cz�F��\5$%;:�����|��gbՅ#h��L���0ě��%���zk�^TWVVq7G���!gy�)�h�I�Դv����z�؋K��3��|F�W��K����B����ن�p�ٹ�l��,֐j��@=Ჶ�7����m^*�s~o��erx�����"�������Ƣ-��a��.b�Xl��(�')�5v@��xJ��b;B|f��T��M�f�Q�|�{�#v���be޽��d�u�&�"֤�9�IeS��{>HI������u{���B,�|+ t���B:��_���ҰHmd8�i�[(��iVs]]��u�����n������1���Tq���`�iZ����wҷ��:�Df��$��U�j*`���k�:�Wa;]��Zi�o
9M�Ԭ���4��^�D=�G��b��Ϣ�:�^3/�3ix�����A)_J#7���tL�9��2;g��}Yo\�̾.Es�<8{�=��.o��׼�h뷧[��Aڅ9U�w����I}�W9�\�����_Ҳ�k����Ӷ�geբG���Y<k#Խ����vj�yG�k���02�#�\R�	�u��Ucޢ�p #���3�?B�{�������镭����(���C��ޢ��n�{�-�ضs�_k�4=���Z�{}l���y<Ң�i^ي8"�V}�[¥c�E 74�{�f�<�N�����w��|6������X�h9)م0"�ơr��L�=KFb>[+��a{�+1�t�Bt�s�a��Pqe�.�^r��[U���wq7D'��i�UqyI">Gz~����N+�V��66t���K���\Ӎ!1�7�XxX�(_�tYݷ�
��B�t��>���A�U�V_Z�ȳЪ+��+t^^���wJ��	cö�%��:�&��J�I��*�Q�0������H��-�������e��Kݲ.����(� �}�#/_�y[3ص�F��
�5�q�4]й�v�ڄ��YQS``�8&0�Z*�4=�)��v��)��Mr����C��wG�l�Q&�+���T�7R-��}bK��o@��[St�K��n26���]kr��Q�5��B��s�FeC���SM����%D_���N��o����=�Yn�pVJE̶�����;���R#N~����L��?W��0n�e�~�A�~\*����ns����x�:io|���ܔ�ӑ�Qmu�U�v�</�* �q��x�o���t��$�r��v
)��p���.j�.���~����K�Ǒ٤���b���>�rF����[d�&noɕ�p}���ron9�����ڮ�/�Uȳ��v���$I^j颯.�IٴO�l9�lIɗ@[5�0��ȩgD����5��NO�}UU���=�)�ܝ��Q����טF�1.�}���{/}��9��zi�}D0�>0�VE�v�P��C��<Cߙ�Z:׻��vR{� �N�$�$��'lĄۤ�|d<�$�=a�,�ߛ��7�o\<HT��I=`tȲ{�XB��:d��8�8�|d m������z��x@�ya�I�=N������N$� xȲ@�C�뾺�|����4�z�1���$�ä57d�����M���I��%�$;=�ق��<��^�{���*��H�|a�C�,��ݐ;C��!��$�'�2N�!�~^�5��7��y}�oi$�!Y'�m�=a� fYP��7�d���{�|9�/����!�q��CĜd%g�Ht�8�Ā��6���� �cʯ���{���I���ڙq�Le�y��NSE�v���D[�y6k����o8���j^��rqRO�W�UV����@ēI!�&�wd���8�l��07�qc�Ha�H�:��|���D!�,�ϥ$:x�q8��Ho�L�,� ��00{Bd�I��ׅ��~��'i�ćL&�B�m�I��O�$�>��Cl�Hx�0ϙ�߽�JȠq�z���d��$�d���$�'L�ɯi!O��0�����y�3�L=a&�ya0�l��CG�H|`t�)�!��N���m> d�|��g^������2t��2t�I'��;H�VI��2Cgt�	��yΝ��u���0�d8��'~Y�e�$���m'L�i ۤ'I��e���|ג,���)�x��C�rZ�'�<��N�N�C��6�6�3}������|�C���'��n��6������ē�I�'}�a��C���x��$:���{��|�C��B|C�C�����BO��m��I��E�l���2z�"#���X��q�X\/ �bz���n��V��x���d4�Bd7�`�g/ ���M�����r�@�?�_U}X��	�$�=O�$8�Ę��2a8æ݆�|��!����I��K�w޳�tf��w$�dǶ�!��d�gā�BbC���Xd� t�|�4�~w�g'����^��I�2O)!�d��L'	�q4�LHq�Rq������=3�^[��u�i�:�:B�2M2o�a:`q����HLd��x�<���o�/R4͡8�a���=d�	�Hx��I���0����&$�d���w��f�׽��I����ċ!���4�2N�s�Hq�q�'!�;��5��3����z��w�&�=2��!�Ei
�z��!�!Y4�6�$��>P�L��	�����i�Hu�N$:I�������N0��gL��$7� �&|�8�]|�oϞ뫞��mI�,<H9d�'L>2N�I�',�H,;d鐬����&�����|��=O��Bb|@;I�� v�=��=B�:H�(��C�IĄ����oI�ߤ�.���JD޼���EX���<\��>���i��~�:��aD�SUt�����q�)�C�{L"� �����M���Bf2���mb͙Z�u᩹+`9��
MX���]�]�,E�(�f�E2�p[�1�kY�U*1Q�;;��W4'��i�橩Q�C�=�l������ُ
��uRnL�h�dH��*���J#{�<�м}Loc�:�ܔ4��n�G���%[=L9[w��]�����K�.�q�B����ԯ&
���]{�J�13DeK�]�8�t�c�۩虺����E�	��Y�)�2QEk��]�guʇ((!���qJLo������I��i
J��¸�׷;Fr�B��M�S+5Ҏ������M\J���]x]�5$u�j�u�YWey���N�� ;��X�HVl�6���2^����K֮[�C.��,ϡ�a`�gP:9f���P�YN�:dfX�� �s�y�aJv%i�-Ut{U���3*`n�'ن�όT��n�gp7d��5�in(Ñ50Ed�0ۂe�b�)ԤZ�kq��:�� ��d��O
;��]?Y�F�)j�
`�X0UTEU��Ń"0��UYQY(�-UTkb���X[U��e�D��ƪ(��@\��QV�Z�cmP�qT�j��X�b[q,V.�4m��*�[���Qʥ�*���R�T�(�@����~~~ID<�n��;l\�T���Y�p�
s��������ߤ����$>'Nϧ�.�;�6����e�ώ7��tFƣ�h����L&��y�P�^����C�R����%��8�����!��a(שឪmd�]'59��mi�[ޱd�Jr��F�wk�Qw�b���,�1�SF��P/����P�qQ'8pqí5`�c"��'qX7ϰ���s�P�賋�)�~s��X�+||�(���ּ���h�c��f����Y�5Α�M��|㘹H�(��W�_}]�����ZPZ�܀�f�ϔ�0! ;�ć�/џ:�궕^w1C]�����r��3k��Pw��_� *ޥ)X�n�@��B�G�U�9�ڟL6"��Ů����0s��lm)�տ?/j=ch��&7�Z�/f�3.�:����O��;���_+�!�Fwq8K�.��2�Pp�#{�D�g�,�Xx_t�17��sJ7�[%���.n
���S�]�N! ͈8�)���ﾪ��﹝ҿoy�0!zW���cG%{�ъ�9����Jl��Л7�v�?dU�+5��L��.�.p�����J*��F(	�q�C0:�n��[N�I�o��|`�=��>�g]��%�C- :���o��?	�R�]���a4��:��[��!�I��%���́�S}� ;�|�)]L$J{^��R���>/ʽ���dѷW��M�[w&�VN��f$a��Sr���'��UU}�$B��,ӝ_D�6/�,ME�3���x�G\���C��;�����#oa���f���Г�n�X:j;b��
yk��N�Z�ծW��6�gV�2u���#�&�롏��HN��=#�M�K�$�%r���6F�O(�~rr��wtoB�
�d�S���	2�앵�Y��c�\(;׹l�KЍ\+�}M�h��U\N�,R�8�"���mQ�f��i�Uq���Ύ��3�cԅrW�� wR�#���9�K���Q]_e�P:��uZ�A/�>'�0��M���>�� ؜t�:���t]y��=��W�$a`�L��Kkj��j˦��˸�M$א��4`u艖�h���c��2�J1�=�]m�n�u��KY�l�$;],�UAѻ�}����S�k�ڷ�P�5.��W8�zM`O���0S5���(>�ly8�7E��M�X�ӕv�Gu�܌"�N7'꯾���)����\��̻�7��:����諌�V�����ѱ�G鶼�AzXS��g��7Y
k�ocr_}�.�y�[����d����,�u9̗��N,�*"\v�`��+S$w�w�����e�Io�lZ�Lg��{�0w�γw��Gk�ٌ4���v	�S�xH�����6�`�t���WW\�E�{���ۺ��a|��?;D�˳�Q3���qL�h%�e򐭎2���W�U}\��V����֪�����K.��áKH�Fr]МX����
�w=K��G)��]���R��n�j{y8�@c��b���.E��|�{
�Yu�S����_��NR�a�u�n�؍o���^{��,{�8��=���
���=�3�vq:���`�S�5c@h.ߣ�s����pyWqϹ�0Ou�HƦ��e�KxI�b��M��crs�\��V�m�B-����ꯪ�e�?w�or�(�j��p�E�@[��"�0��E�<䋾w���ۄ�\5�"A�Gs�L�Pٳ=3�M>��ؙ7Y�}��o�(] eA��dKCB���7fIOs�E���v���H%1�z%J��0��._C�͵�5/g�ۙ�Vǝi��=(l�=t���U���e/JX}�p*��0����2�%/&�ժoa���GwuE������hs�!B�r��E�܎~��ﾪ($x~��=��`��C˂ҙY�A4�@��Q�h�Ԗ���h����ب�3�;/-����M&��pbU�tŘ������w6�j�6v	�8y�X��ݚ��Aեi*�ڂJ/z�=�,��V����B�v_�9������L�L��pZ��Hr�m��h�Օz񳀚{�HEBg�黔���[o�p�ﵫ�՗)�%qz�H:I��1槿�UU�U�/!s�Uƿ'����zҨ�~B��]����d8�ړW��Dt>��=�����x[R�by:�h�_uS�h>ˑȸ)Pg:kؑ�����7YP�u���צ���0�3�x�g��s` �ֵ7��kn�T䩓�h`Sˬ�\��Ho��=~�o�^�<���Bp�#P3M��P0�]چ*P`��H>��\8�sV�C�6��V��f��W�Zi����|	����Y��L�YgK�QB\�Uy���ͱg+(i��4�'���ʺɈ�4�mK;P�ƋٹkP���ca�D�V��r�;z6�IgjI��5;]i%�YԀSoE%��Z�	a⣻d�p����A{���#ib���0�l�ˑ�]by�1(���Q&�3,�(��]����Qw�y�heF�٣Zt�&(�ۻ�vy��w���_]�k���f�[̔�!em���ysg7e��|����~�E����䒃����|㳆��lX���pخ�*D�����Nu��"I��`�J�#�˺������өQ�i<��P�&���δΰ����ޝv�Z�Sk�
��b�|6�.�I���,��oG�E;���h�!�˓`�w]�귕��եhcM
��.F�qY0�u͕�������,*��'>[�M�e��it^D�5ڰ��ϻ���c�u�.˾��I-�O��_\�u�I xX�{]�8�`�:�1���2�5 q�gEzM�MN����u(�V�I��؀�H\'>2�:0id�Ӫy�~y�<�z�_�׏��Ҫ�VҶ�j��12ڍYF��E�-Eh�DBڶ��W*�+�)��ij���m��m˙12�D�e1J���J���J�EKkF�ZW2��J��E[T��e[el[B҅J5˕�[p²���3�mT��\�VLH�E�!1��"5�'�0�Cm3X�\4�)������k�4�6h�2����][J�F��.*87�-���Kk5r�k
��H$A��1�l�g���I��`��:�%���E�Ir*�ﾪ�O(o�hD�Y��M-���5���n�`� �3'{�#]ڔ���QLx������Z��C�^+5p�=Zr��S�.�)���v���א��":n��+9Ov�y)@��:����,uv�E��.oNƩz�̧vm�)kt8���U Y�f�\Ϫ�>���L�Y��`�P���7Ck+���ͥ�6] I��G�����%c��}&?.i&�����;j�;�b���S�-_"Ky_ޏ{�����X�}D����/3;���n��8�f��a|�5��@mq��]�����xR/-W��u$ �.��<i3�N�&��1<s�=��^.+�`0�&���oT��q+��O;����'��[����Gl�vi�s�1իk԰��������q�2·s�M��j.&F�êsn����[��:�:$=�ҝ܍�Y�9^�Z�Pn>�AdMJ�b.x�6���!�gb鰊PX�dң��i��}_}UV8f�����pM@���9��Y23t���#���%^�i|�{�j�������2�9�D��e�ʁv�f�*S��Aⳝ֎�
hoq�[fIp���uRq3�>[�@��1���R��r���^�׮����q$���Hv���
���:�o]���;�/��!� �%ê�h
����d�w��&���J�m�Z��CqN��Qi��2ј�8n$�ԗ����z�gn�?'��@��b��&+��xG���՞J��?_m�U�;z_�]����fn�X��769@U� �-�#cR�zl x��-�	����hё��	m�c�����u���;.l�4�3z{Ҫ�ywZ�R�L�湁U����z�CU��g���!zU�����i�����9�-�-U���O0��ر��m;�uSP"c� lZ�Y}.��s"U䔍��=�oS�cPƛ�������Mp�
��,��Y������[��|�mv��nʽ$��Sg��D�fvz^C����N�`��g]p�O�銎4t� �v���O���	:�)1d�x:/�*�d�X���%Ls�m���>d�<B�c$H��Ö"��z4.��kP!CX]��� ��k�x����D�\\�e]5a �g����vN-(�j�.MT�@�B7I�_\�^����JI����꬜�g(��U���,v�/�Vx�Y�[�.\�A�b�!�-w{k�3(�ݸ''����vj��x�]u����B�aE����j����ڜڶ5=ԑ5۱�2�k�Y��.�5�&�2��8����o^�):*�i5���m��� ~�Z��p�0�Пq;]�
�%o�|}�Gb��[7|nq�˳)��n3#�6薙�Sɹ5�M]�3yN}�U��I���B�~�����yt~�$���DP�e�H���C�G��;+NSl�ѿ^�(���pQ֜��yq�G*/hu49W���zե��R^p�t���׵������v�;�2� �^uݓ�f�i���q�e����[6��]e���"�CH��4��$v�uv�v�''��h��J�]�v��G	���7��g�C�6JŏAˠ��Gr�#�i��LHc�_��X��`��t"p��^��8xn�/�=舞�sG�t���,���m֜%�P��b�}B��=�zn�!o"73\,���pf$N_�Y�އ�����Ѻ�|�:# (���A�,�ͼ5	�#[
�nx��5�����Dt=ی#���n�.���nM��$G ��Rx9x�r;�'�9�M�[yٔ�u+۩��E�1����Gux�spkkG�ߖ疀�ޭ'H>���»�0�Ԛږ�T�-_J���An̢]fWbtI�")��}_}SKelC�7���)��H"��I�ff�_�%.�}~����.Wz뼜�zU�.̙��kC �~�u�M���uҺ~UE��},#�7\َ^}�U*��|(L#�g@���z����v�D��&��Ʌ_�`�N�U�N���+0��jJY�.�H��M��'����x��	�zH�T�`t���q�8S���^:��䞒���+�c��[�v�d8\����E���ﾬ�Yޞ�Ev׬@�~Z����<
M�]�fL���a��"�W�.uuAg���͵�yW��)�*aK�yH>��h{�90�� �ל�C������}{ɿu4�n_��]N�k/60D�wZw�q(]�;x�[���ՄOAG�eY�Y�)����z��UMVT'�S'Z�p�������CU��<�珽�{W�Q Z3�����
������L�T��a�}�{:��Y�i�B��.��V��)�{y�[�G��q{�A�^�cr��p�U.��r�ر����;�U�}d�p�z�v�U.��f�B�!oj��&�W9Gw��m��.����������V3)`Ü댈�L���f����}������2�i����A�S̭�\�4���M#r�uy@�pܮ����#Ի��4k�ƞ�Y�h��N��Z����QڋV�ck\��nr�j�U�����:�U�k���a�t5574^o	F#Nr��L���A�0eJ㵽�:�����|(��Z&V.�n�O�-��q纕ugt��%�&8��˾��ɝ��־��{2p;Ƞ��";4�v�Y��hU<�m�ީmu��� �O�^�@̔�7�����N��[�B�H�5�i,�ي�
�Ր��6:�S������
����*Es�[��J�3`Sx�)����h��2Aý�at%jj�"dޝ�?���
�ߙ�&����j)�*�mQIIV/d�������bU2򒩀nE��cU�[׫���-L�I!%�K��[���ufe�q��Dk�b9l+u���a�Y�sY��TƵ�ԭ��+V�Qm�Q�aG#�VkKr(֮��E��4B�qYX(%��Tr���c�4,�m�VZD�UTթ��4�Q�*���lR�t��b���J����ٌ�Ҙ�\��n�cm�J8�ıUPU������Q�+1�q("���bY��e4��̶]Y���naKeJe31��U�)WYr�N�J�[W�m���P�,F�4�QTKh�0���[Q113�3��;��/����F��SU�
�}3c�!)9?���<G����>��H��89]_=��	p�����R*�[�P�C*
�F���+� ؚ�"��Ɔ���<�����q&0����Y�l���y��޽�y9Ӹ^�8����#�Z�/��"�n3,J(�Y9��GJ���8!>���8�Oy
�:���5���B��	-���ᗸ��n�2�(Q	��%�}|�ǈ][�
Ȗ��y�Vy��~�b�0w��w&���\�͊`
O]�3!h�
2O�_}X�G��ו`�H����D��x�x�K��,���U�V���S4�'������I_�����k%aЎ;�
8�]�βm]ӕwM���^�駮�^��q�^]Q{����8-&� �N�0*��g�M��h6iڰx�`�A=���o2�X��:h�u��c����%�ݱ(tX��ͤ���ύ������>�@�
]v��ѝ:M�Y'�RU�h7l�4̼fD1d�&���	9�ꪫ�	���v��c>tM��α�ƒ<n����]��n򔷇u@�����p��ю�M����� ��|'/�T"v���
��&^=���{G"W���U�z5O$��"��t�WA������]�čջY*�;Ҳww�U)O�,���������r�$F gc&]�Ò3MV�!���i�ՀGoc�p��.�8�(�E�����m�o9�̈4�N&��_}�S/o�>������ܴ���g�G�Z�i�5��ᚲ�J燨j.'�QD�w�af��ħ+x��*��*�E���S}1�LDix�XS��X�#���]���UO,0kƷz�3\.���p��:�/+��4����c�9��ԍ����˕���Xf���ugINan�)FuF�4�^[F�����W��2`���U�ANe�:T��$1�uV���B�8��_W�}��]{?J��g�7t�� W-T�tj"�P�����+���m���fr�l���n�0� ƒF���v���ե|�Y34��A�R�$cn�=UK:.t��1P��{Dk�q¦�+�Ϙ;t�"���vcu)��� �q�;�=\�ZR�D�����~��hpܩ�yѧ;ι��pD�5�N?h�Xd���Kx�*�¯7أ��C_;]���Yg�2��S(�p�[�)�_-bWMh�Qi������M~�+���E�R�"k�����w���#n�$��Hy1�L��pN;x�m�����}��I�c@�T�؄�9�c)���	���ژj�U0�������w}<�WL��<�J�v��;je<To'��l͚=Ux]ΔᴰO�PS�(��q�^��zj\��X��{���jB��չ�����8+�.���T��Q����o#�&��	�<��ܽ�r4㟾��������-����o���S',����^砗�[�c�������f��a`J:
��f�$�V���f\M�1-�%��2;w�ԍO�!(�NtL��w4�`�]�j����l��}D����,�,f�9���(�cw�������SG��;�n�^u��f8�l'�}��:Y��5�`ݕ7\�e]����V�c� j�q�ۗ%U�\����3���95�'p*O�}W����cL��~���J�0j���0]��@�:��B�Yޢ�VBPnwq"`k$���������Nz͖�2D1P�1\,bg����k���:*�
w��E�{���0>�q���������F+I7�tZ�e�%���t�U�_I7#~�>k��;�Sn�-���v�aXɺL5�T��M8)�h$�B���FJ2nМ;��}�UB��9��q�2F�����m?�B��bL��Vw��<��3j���~�xN�!Ȇl-���79��]f-B-��m�#��\�mv��f»���8��E2Vy�ߚ#nm�툷4���_�tb1ɸ4H�٦��9�pl=;����B\ԟZ�_����.��E׈nO�!�hv,�e��S��xڒD��Y����W�v��ar!ͩ.��B,��4rV���B��
���\%�����߸�
��]�,���%�{���;��䟳U'�8��w�qK�}=�C��aa���ڮ���������rDK��WB�u��m\ʏ�}s��:����y
��S2��Cy:�B��o����d�Xc$0�!��*ʠϧ���ŉ�S����װ�S��|��p�X	�ޓ���a(\�ޱ����n�S�Vr]l=�v��h������5��v��
EW�4����2��]i��+,bZ:bU����U^4���j�tv\X2�tyм$��;���;�I-;¨�)�^���m�(3�fX԰VU}/[��;SZ�6F��\G;����t3� �.8�C�E�osDn=D���}!u*��2�b���{y��$
��7��.U��2\�&�VK��2�<�]T�f��{y�˩}�tX�X�,m��-�ڢ�E!�U��mA�c99ԞiR6;1=wR]kpɆ�v̭ ��C�$�P�G�D�em�%C�-�\��ǭ��\�v^�]p�i��,���(�$ܦ���v�p�3xT)G�n��:0����S.��/9�ج5
��f]���Kv�M���◫밷m���w��ts��6l�'R������͘���u�I[NԸ��� z�!����B���݆�_\���c��ɻ�GRv�<<��rݍ�	��>Cx�|m���u��ԑ�	p���ecR]���i';1��Ek}�Z9f�քǙ��/�RX��d�{����J+�HV�$5���
D�6�jZ%i�˓0�R頪�7XS��Z��UV(�Ds3%��9J�J���պ����kTKJ�
�n![m��Y��ȳV�1unkK���%`�F��*bc30E�������S%iuM3����:.j�td��0ոR�jՈ˙�Qլ�Rۊ�mnZ���*9��!�¦�SV���*4ˎ%M5K��k*���J.KR�uG2�
��(�-����e�k3a���M.k
�+ZZE�J���ɨ~�nT���D��ID�)�g6��Rn�N~�����5~Pq�ٻ�#/��35�,Y��)Z�y:��ٞ7�'�|���4ۙ����Z:L��m)7q��c<,9j�i�����ܞ].��o����k*U�o<���bu��M�%U�VZ&S�$T�C��p��f	N�$l�;�����GƦRPt~���e={W�{�pUU���M7��U���6�T/n�W�R\N�y�����o���o�Ǜ+�������9g�E��~�\���,����6�����>���d>�U���b��RKom�͔'�qN�VLy����>�fF(�2u��:�Շ&�:�tLw+Y�&'�ڄ��,���|DW}C|��W���������,�4=��ZUi]!O	:���KS����-ux2E��F�p��z���
�M�h���N�9��MӍ^�U���Ru�h<�Er6�^�b�f�s�W�o��?	�²��wZ2�3C�����<�L���"1�u�\M��������qu�[mb�p�tl�a�=�a��8�:̣�pm�W��r'�qy�ͺ���S�%�j<m��$hP.�U�`��8�9��~$ ���w�\E�O�x�\��`��Z_��<f���Xx߲�҄/2l՛���hy1s��3�a�ӑ_�0��5%։���Zu�%�G��G���r~���6�~�(����}�&= ,���*�r�L\]LzaﯪL/�b��tg���8�N'Fs�0�<a�S�V���b���AI����6w  (ON1�R�VZTe���:�yNUN�ۑy��im��x%�t�/�����}4i��견.�fm�-���z��!l��9BU
1���g�	�[�q��H���׃(ʵ�˼��Љ���W��1��9�Zˍ��Șt��2zR��]���|���J'?}��W$��ٖ?%����i]�L/�h�W��U$���9Q+��W��y�i�EH]zO�ֹ��d,'s]���ޓ����d��;}S�^�)��tk7V&6u�F⌜J�A�$�������<ȑT��L�RR;�(�iݓ�Z}�m骞V�u8G)��US��K&�n�ο^�F�pjT�ۂ��m��:>�	2s
�v,;Pa�<�0i�<��;�[P�O�rAW�mo	w6�\f�;8J{�f�<�n~��DNp;C��&e}�.�&,�����=�N9p�;j�im
���gXsw�����X�㕴瑦ѻ��]<��u�+Q��T4��x\�Q����J��/~^Q���P�������������лK5�+�K�f��]��t� n�4dOn�����C����/�m�u�冼���^
����:���먽v����tƜ8�Tt���z�쮼G��- %�`yC'D�Hю~����*~W�?%[U��N�to����u\�,T�n���`|���ܷ]�q{���Gk���+�3<�.��B�-��X:�u��w��"��{�m�+�/ Ewg�L��̓�\p��}0�o��ho&�+)ኼ�y��l�c�Ї�+5�tB������T�w���P��`���!��]�U)�����7�O���m�����t�A�W����w�^�\\so�ҲR.S��V���=_��߼��O�ϫﾪ�=:��s���2�eGV�_n9��AR�sj������s��9U�W��SX�����E���@��s�J���Xs>�j�<�׻�v�O����XA�ګ<��G��7��C��Q�>d�һ�����������{�b�@��K�N!���s��g]`���N�(�_���ټ�Kk¼Wb���{�L�7�&%�\�+KZ|c�.�C]Ki-��>J��ݓ������UWŀ��������i���4�.���4N�]+�/�Hx�y�:�ưHއ�@���R�9W*n�ye�9��TDj����ޓ�lר^*� Rܾf�`s���H��!	d�{N��J�[�2���~��й)�VDО�v�
N��oM�KI��z>�sS����L��W�:5H*5��teʂ�֫��1�>�FM�wp}[t�+�n%������{*dɴʻ�rt{|�����{%��I?��}�j ��:HY�d���X��$L����:�%�@8�o(׷զl� �M@�9�G�
K'T����	�S٘׵�����3�E�Y�6Z�4�e���%eEq�pu�w���]��S��q����g��u��`ѓ/=��g�t��T��P�I�"�l�Ě�9ٛS0�ܞG}1���>u�՞�G.,�tm`��)����pm>�c]����ڊͲ��%��k�F����{�A�р�q�r��r�h�f�+��,r̜��;�&�պ�������bו�m��I��X�s\!B�cd��i��Ȅ����ŅvS|�tgf�ا�D���\9�:)[䬡6���9U��4����k��C�v���yΥ�Rh�$B��v�k�o�.�T�T�Տ&V�p�k�%է���d��
R�X^���[��V,��8At�3�1�옣N����zNSr��)T�Tx���[Y&>�*Ds%�p�[�vԭ�xb�I �m"e	��Tەk9=��E�>��r�\z�(v
�j��1�\�k�O=z�+��R���5�s\ɷ/�3�>�zw:Ty���n=�ը�xV$E�:sj�3��N��s���kv�X[�^��\n̘�[g;2���t�4����q�y�𭙻�*x�f���O˛��P��&�
�T�[��<�.�mm��2a�"%tfZ�RK��ѽ<��0�*��mȤa���x����.�z�6�ٶ�s�Oz��j�뤦 nQժ��
��YNw:ӋY QD���31�J�\rҥ�7�3�iV����Q��ec��L2R�f�4R�a����fe+Pƥ�e��u��E���-p� ��\����.ffU��ˆb��-��L�aL̪� bTYY1Z5����.[�b�.�ua�Z�Ѻ�
[QL-�ڕ*��c��+J��j�.L-Y�e���f��u�Tծ�f[Sie�k4�8fL��+R�Z6�p˖����UF�	$�h�QC�{����T�El�bdPme�(��J��>����f�g�o��������J��⩭���������H��	��m.z6�ä�1*�60a�oZ73�ewc8y#�z����mvUE��)��j��I�Ϊ�P�jI|��ތ����w6&��l����|�-֗��֚wz�Y>+�#�7������N�f@��;/Kd�/s*��}Y�BB���"��Wu�|u��K��]j�da���LնR�L�ق$�f�着il�¿hc^}��b���cT^L~�i��5l��4}�J2�ml�EW�YZ��nC��&�np�47�Ω���z���r��ګ����}�'�[�_��a�8��ݝ6�gJjr����k+�yj�,7Cc:J��b��^�m�3�8.��)!�[�(���.C�ݙ6�^a��&Ӹq-
�C;���s��G5��h>�O���>NIY�x�������d��3��r��Q��ȜCP�~!�\ˌ���Ϩ�����K�4!���6�h��ʠ��^x v��Vbk(�.�Y�2:�-T����`ړ��Rw�rǧoq�𬧛�?+,(�}~��y��:>'��^�~�C���g����4���Ŝ��+��Tt{�V}�����C0�@���,���FH���/(z6�éat *B�k�=��kՇ��*�ϫ:�N��Uk�}˞��`���x�Z?umjSX�ri���q���7y��)��KC&���6�	{cN6`�h��I�y� �]z���(���ֽD�v�wjn��}�w��)ߖq���Y�Pא
�0�iYճݿmd��h��BȮ@�o��0�&Ue��6�0�/�DcT~�4Q�^#�
ϪvKޛ�c�����k�]�?Us~�嗸��R#|���K�/�L#]��1Ǿ_s]u�LS�//n��=�G)�R�[����tH����di�(�,�a��y�裵*��h�k�4Fj,d�(� �ʙ�Wg��xR�;�Mu�zy�8Rǻ�S׉���s^z�nˑ�
=���$ݱCus�9m���r���k��ɪ�ٻz�Ke�/`h�q�I#���н�Lvҽ���h��������C3�|���'�V�֡�0�dY�d���=�cc�}����~�ۧ�:�^>=�Y�����W�@҈�U�R%z�������G�nuVzU�GG�j Ξ�z��cl��/k}��t�#��Da�����\���"�Sp�����Q��u��]u��}�U�T��� #��{0R㇏����"�0/w]���<�5,����6�1g�4<�8W-����6*͙~��������X?�,Z�52��������ȶ^جO��j�9�P�S0��5e����g{-֞2�Tz��&���%IY�)6|e&CK��MA�6��@���r�\��;����e/��Gr�ZFk�x�=��#N�%�Gi}V��ԅ�Xs�'�~�Cg×yJC��w �i���@�/eUW{=��t5�z�����p0�äY&����m@��!}�ŭc�O�(�B���M�Mxx�F���G��?z�Qw�����}���W�����o.�������4{Y����ٞ}�3��N�8P?T_q��^̩�h�h�^><Mc$!��LF���Q�G>�Q�}���>����6�VW��M�m1�J��sK�n�ہ�E&�F�UǕ��؃e�$�G�����%N�w�=��x����.�^�{�8��q�^��0�0�R�e���iLc�m��3�������'�W?�C��`���-}��QTC�F�Y����a.:<x��v~�r��-���O0�ߴۉR��7�ǜ�k�޶���>�<_�B����k �P�.��ѕ{W��+*6C�*��\fC��gbv��̽1�|��u���E�������Ne9�,TcWѕ��:Ik/2�J���M���9�<�&='^ӽ�zߞ��~��Ǿ^uM>�'�t�<�]Y�=�A��gB�ٸz֥v�C}v�GRcvpo�7w��;���	�w��&p��,�zo���^�
��*94�'�_�A�)���󞘀b����KbOq�K�E�a�\A?^��6E?TG9�%�Z��*��M�{����8{�ӧ��1���] ��y�]^7�v��sV�N{s�zp�C�}د�y�y3 �ER� ��th����~�D0VoS˦R m!�0O�#M>�tX��[��<�g�F�����wӎ;�n<���:l�}����[�|<�����c1[����Xa�`��0��xl;�FV�eA�ʁ70��ƻ.�0M��bˤ;��#�Hd�9ٵ V�7#S�s���Č8ʬ��kP�o;@���\��d�mb�/+ �,�SV�:�N�7�Zn���S+�Y`"�hW!�B�Y�t]���Z׋�|)
!�Mx�,��0��|k�?t�wo��j�ȫ_U�!}�[~ڨ�<�����J�&\<����7F��j���L�p>]:��}C��c�k���M���VOe��ϑ^h�:1.�>?2�XkX�M�f�7���p���@P� =�	�N6o���vx�~��GyV)H��)��ty}}ﮓ�u�<��h���K�3iQ�61��^>(�xчw�+�h:Dֈ�@�q���+��xh��F^{c���λ�N��5���|sb%mg2/��
L�w+x[���'&s��#���B���A�����&TJ����n|�y+|���z�)F�m������.����Wm����5�����z�1vP��#A�㶎w�ӝ%���G9a�V�����sza��G���\��3~Z�6�3���P�����h��<����o�Q)"�)נ����XE"���p����p��B,/Vb�RD"{�rޝ?Q	�,Vg��#�Af�|_��.��L���h�Vℜ�4�ha_��ǎ��Q��2��z�յx��?:��"5A�iC�%���k
xCy �9���2��}th>�S�C:��W#�u6���7_hIQ� z�G2ƃ{w�����R���̈́2�̨B9��N�ZFb�
���e*͆�C"f�%��u��xf�qO���֒���r�8��T ��k7u�8�	�jbW��{�����mdw�B�٧ �2͉j���Ern���l�u����L�:�=��Ѯ����3r��!��Ǘ�R6���䲧,���@"�seA�)rC�gt�U� �7fivE�s;4��E�pdxk��1�[��@�ȭ*��*�e���{��K���9�1'�PЅ]�rX�F):�j��1=��[s';z��|0ջ��c2ЖM9W��';�2aUm�N�nk�7L����*T�Y��D��1EUA�d.9�B񍹕���%ڻu��rܤͰ>�^]��yuu�7��cz�T���{�BN�c]{�_Kȣ����x�*!ֳ���iOs�[�(�jݬ�Zt�{5�y�;C��׻,��ٖ���r}����F�n&�r)�@�ԕu�cnM�D�ѧݶ�5wWcjf%��kӰ+ʥ�VJ�G��-Xa�Y�I4��MU���u���Q�f\�k��s�E��6܌��"LG,ĳ���fSM5s	SI�*�UpX��Yr6��-�S3j��l���ˎX�U.\n6����̦#�TI�ᎳI��:���L���X�q+GJ�L��m�e�\�QQ�\3M��,V�T���TT˃���KK�̕�S%�Z�ȵ[J.Z(�
+m������<������
YaD�7���'	&����<(��~�~��yVn��yP,�B��
�/ۓʺ�[VGk� �A:CQF��<�7c�gn��"j�ћO|l��ۑ�w����{�>k���B͹�RFR��i8���D	E��^w��{߷�c��T����o���;{{E�Oy罺�oޗ�|�h�N<��ݞ�À���<`jZ�{iXDH��I��M�9��D2��0�I�c�tsP�X�6YhQf�k�NQѳvE{��]��X���F4���ȀM�\����Ws+^{h��c��-
:E�z�
,�y�u��'XJs�v� �+˯U�ϔn_h��st5!ɔ ͉���t��N>�sLkRB��u"�:��_�Q���Ӻg(^ﰽ��.b�(e���DPIq�+.�M]�����1�ޟ[�d��9g��(���m�]l\��XDb�k���
�㣗�}��Q�혋U�"�ݙ���c3!e	�Pۿ)�,#��)�n���`����Ǳq��`�l!D�evz����b���]�=	���O����{M=kѽ�op�!ʊ���?^+�8��r��7�/�~�!���t`�s;��ֻNǾ�5���<�5ݯ��'z�����Fϲ� ,kT�=�Ua���̓^�ݣX
ݭu����rl���ñ��&�f�z:�U2�9��&�J!¼��_3t�&Q�@�nc�n�����f.><p�e��"�цU�p��)v�f֙�	�V�ߕ��2�o�<W�Hv���)�Th�8C����7��D3��ָ���B���1py�-�d+���?t5��n�C+��,�F�����MB)��mm��8�R���C�*��h��K��	�]�s��Ŋ{NrQ�h�'g&0E�Շ���f뱖��v����Vk�e��vj���5�=�
T�n��?�9џ%�P�ʭa�a�D��g{��I�R�6�pƬ-�+�]3���EUb���f2pe�g^�x�E�rF���ɥGӕ�At.������W.��oʔ9
���oϻ��"�����#ƹ]"P�a��C�^�zZ=A$��O�h����C.�E3rv��8��4F����DW����۾hVӄ>�/+P�!���#?y�ֳ��v\D�uј*^ҟV�9��:������mF�����Xp�AZ�p9<z{ثڸe�P!�㑰!�@�PÄ2o��{I��c�i����x�h��ƿ�����ҽ~�6|a�cl�N�}�VQ²g�[�}���j��o������t=�|Iz����V��.CSz�΂�	�����y.;��zd�)%�<бu�C�]yOV1g�7��(���U]�G%�������1QaB�a�zt�FW]�U�G�ӧ&^"�s�x���ۦc��Z5z�󝾎��7�v��q����}�ol����=�s.c�,�~�ƂgH��(��놈f��r���}g`@QF�z����*{g��qYn>=E|��7��N�8Q��	�b��+W�#�}S���t��ZN"D�c����^�~���g��WN&�޴q��>>"��k[3ޯ����Yj�#ǋ.,;ZW��D��?z�>���ֳ��n�T
\hc�3]��B��nE*Wl�i���'�zMrZI�cI�@��]t�YRg�Q�ě:s��e��|�Vg�Q�8GK�<л_#f��ㄵ�����]L�#ݏ��b������"��+�I�39f���:c�,�hQ����Y��N�u7+�w�-��C�jF�\��P�_�R�MԳW{ulѳ��h�N�>6a�-#��|��u�;*��iI�m��B����̆�{6E�����"�K� x�ũd��ϥS,��i������Z��+�������N���/o�_�l�e+���	����-^�Ҟ�����Y�u婎
D�!Զ�f&˧>����ͨ�`"}�c��iI3I��uި�>"R�!C�����4�Q�W>�^'��z���M'2�s��t��M������q��=C��)]yOwt�9טm�<�ĦN��q��g�\B,�����(X�{�t�#p��k��ȉ2+����m�t���Z-�,y�h���F 	h�(�����z�:�s(�/r�/����y}gR]��J�7�۶Y�o��KMJb�t���д8�]��dY�y<���7N�c�����w�(̠ER���q9Y�V�C:ED-$h���4�w�ϥM�Dp���:���Ww�#���M ���w��]e{�W%϶���FwG��*�󓙱2\�)&�;!�|x��q�M�ȳda����Ϸ��V�v-�Jߍ�YF��V믹L(� ��W�����r�d��׺�ݕ��&���z��v�~Цj�;��]z������G�*�6|F~2'bcU=�����zraϴT
,�ʹAH���A���=-ZKOv������M�|z�=��W�:�t]^(���Z�kDi���(�u_z���z���G#���%jHa� �:Q�%T����) Lt�r�=��x�����1�4��δX�n�N��5����p�5�+.=9l^��Pq.Ev����bl0�+7_E�8{�N 8.�&���E��7T؝n����|���ϝ��d�h��}e������Fn��ΞjȄ=�6�C�D4�5l��ckrhs�^�Y��\^=�+U���_x���V��;i��z."�� ۃ:���sj��b;�І梪�X�����8�D�bZӤ�>����=��{O-=�0��μÿnӽz���K�N��x�Nl���ǧe����G�D���t&!1�x�e�?YdW!�%��g�5��Ūޭ�)�L(�d�Q�s_��I���|�k#��;Dسq�ի1�o�6YRoW���-�7+P��@��.�8��8�3�U��k���[8��{rd���:gxw���V��ϰ�dmϪ|��h�^>:Mc$��x��r���{�So�m*T�~a���,Z�i��mn�z�O��Y�ߘ�(B�ʈ���ps3�ntH���#�})24�g�_?��"�qn�}:}�/WhqV����B�6Q�����wͮ�O����)Ǜ�J���&��U!��B��c��C�0g2��lܙ�:�,����Am}|j\�<Fձ���3�˔��]�2�2v%ɓ>&&|x����9vwO]C�{uץm/[�{E�s��%��ʆ=Ñ+).�6�:��ܖ�[�F�j�wz�(ڌ�|�}iFi��K�\�A����P�5����Ǽ�޼JA��H:�b������v���R�d양�X��v}�;@ɺ��е%���2��>1KVւ9cя[��=5����lYx tr���+�#u /b��A�vɗ�Eg��V<\��ͮ�`�]	N<��&�!��]��eU\m�w���2�@�	VE����:r�^;ʳ(?�=ה7�H;�o`�C�/K�}DiC%��L�qQL�uK�\*��Z�~[յ�r��$ME���1�.���cK�,z��<T2⛶�"���䂉�B;B��Ú�3�zngSɗ�B���jXq�����P��f�ٜ��J��Cc�MhU�O�YB�"2��+fzx�Y�)�ю��y�6hL�#�����˯����+�x����r�=œ�����Fr����P�6�B�Zݐ�.�K�����(�c�q�YzC]��gC�>v���F�D�)�垚�X�&��F��#�ݑ��.��m9�>�Ε�8��4N�8���ewR�����Нf��י�|9;HҞZ12�FڋZ���L�ڱ����Yp���c�1��nc�LL��s1d�V�j�r��)KZfZ�E.�Ջ4�X4�feɑ�)�[,*[f6�c+h�8��E-E�UT2�U�al�,1 ���.�Ѣ��S32�-��m�r�m3 fZ���ƨࣙ*�uh��[MfC2�5�s)����ў�������Y�5쓭�Sk�YTAH�#�A2�ͯ��k��л�u.��	h]h<���h�ޏN�08д�%�0���]�2k��t��JM�Z�j��n��(�m]�7���:t��\A?w���l�w{�!�	�XGTd�8D�=ha�VUU:�V"�G�u���i��k��������{n�����Q��0��cI�jw�����]��I��y\g����x��o�m�9S%k��LF��n���D+�N�s�06����R��q�r�D����T�ۡ6��O:��|��ս[�F�Jҕ[S7'A��}�����/kL�����S%�4T\���Mqv�4��8�I�ۨ��ۼ��]Ov��/j�}<���.�C��eˤg�-�|jS��]�͑�9W�OT6���Ǎ� @�G/�! -+��[�ڄu�xy_�!�"��4Q���*���9�fy�K�k�9C�V����#s���3���G�+i�k�MR�g]�����s��^�릧O���O\�40߹��5��ٯ�@x�8Fd\�O�ʉ;�9Z�5D{׹^���8�e|A4h���]�Q�1Z>�WuH1�?c�<F���"�#Mr��i��N��֪	w�N����\�r���ݧ(qr��j~��컹/ k.vf�0�&�����\�'a��5��r��KUcԑ�����F���앾��h{���g�堻Af�F��"�
[�z���Ox��H����J�1ֆ�gO@�:ט����vswx��q����_:�pG�d�k=��"�ԙ�D�@x�B��pþ�+�g��,�j��������l��O/s/e�4p����g!�CAa@����[�qi=�������,ȴ�!\��K��_*�m���uו�^>|������k\�oG��έ��٭�w��NSY/O]Y�޺��HsB�@ȫX:tn�c��gk݃�f��z�^!S{�اj���sQ��w��(�Ǧ5زc�Sr���rU6�������e ��Li�{�1�W�*�N�8<t�~XE�n�����,��^cb��W��I��c˘���t�M�!��b����=�Z:��Z<�Fb���ق���QQS��0d�DW5�q�P�h�j�y��~�C|W�V���ܦn�����Y������49i,u�S�0��][���^u�Ȟ&����Ң"���`�k�L�옎
@������c�۾�[�֧�����^�	���O}���,��4|io^�����y���<7���#Ǎ�z����.��͑��^�Us�FȰ�r������%�'I���!Ot^��A��9m�F�]<șI��m�Am���w�,S�]�Vڲ��B��[~��[���f���La~B͑G�?/VAY^��w�W~,�9ih���iz��틹���z��{��o��i�}e�[zx���Wt�5zt���F�X��BL#H�l4�o�*���f��TF��1���>Ś�N0��0����׽��c�E.&/�����?�r���P#��+��Y�H��$_AkL1/=c��Wp1,���"��j&-q�,��Ju[m��\��{�p�<l�!�E!G�dX�\Hψ�^��z󟗂�y7���5�[آݬ�3�(��1x<��RL��R����qL�h%�e򐭎<)G1'�e�VSYJ�g>�7�[}�m(aq��l�aG�i�E��G��w�����҇9Z�Ƴ���G��T��;f{�^e:��Nsxt�y�v�����:v��y�b��֨��+W�y�g�×e�����0��y�x�ŃDM�f�p���w����}�������W�(��{�q��\�۝O �0�9�ՙs��S��q#E �����ރO�׈��\�G>5��w@�6n�mhǇ�S/����G)k�־y�a�g�z_��,]�M�5��
��4(=�YKL&� #�����v�&����˭�2�ki�nKЂ����볯.�˫#j��c�c�>$�U�V���;�����P��t��,iFOg;N�&gH�`�DER'K�-��ܷy�f3����E_i�I��W���]�s�7���0û״���Ίx��on"�j!��k۝�t��Rk⋵���5�6 .ZZy��h��XCi����|���O������w�]'���~�fјn�xҝ�>��9��`Lk�)�ԡ����B쯹�����t��C���K_YDJY㑰��UG&m?]�¼I��}x6�Yj+a��H��x�^���N������ӛ�5L)u9{�"�m���KV.��pY��x�G"r���mm�7�c1� �l�!���N�b�,J��ϼY�\t���!��V1gԁ�U=�W���z��P'�y}QY��V)4!�q`�-�t8:S�����YF��$2���C%3�wӄk�a��qI�%!da|p�;����C>���Q�C1���0�g�,����*�һVh��d
�4A{�H�~���x�s<�#�h��%r�+W�`+�#���OH=��7\����yLT�B�ETçNh�*�l��%��%_�!i��f�b��yx��
��*~�S
�P�]�A�+BrklN'*��)��<G���e�N�:RZ��Y.h�fﯨ�C��y��Muy��k̾�z���ǎڠG��X��5�����񠕟��r�z�Ї�e�j��9;_Y�л���e�]7�oe=�d�G�Z���B�Z��~�׵�&D�.ݒ6��V=�l�W]u^+�4�a�pf�~�_q���f��m!U�d~s�<��a�Q�gO�蠒�fj��۞���]��C�}�:Tx�"a��%lv��T��c�]q
���4�tzp毴�E��ǭL�<�+�_w�U56X���W�*�!U�^L��^���g��d����P�o���E�x�=k�+>�T�_������辺Ro�b���y�=���K�����ZȞޝ+����/���j�i��sÓ=������V�|D�:kW�7����o��O�Q7M��S���fq5��u�<���q��OY�,G��5�5��jT�|�/��;/[�Fw}k���:��cS�т����t�{�<-C����0�T��@Y�3w���f�]����(Զ9�X�p�\_�?B��RIn�!��?#E��S��0z�s��;��t%���&|�*�{���lsT�����~����?�?E+UU�Z cO��0  ���,� ���y?�z�fae~�Jf����kfw�N��nӦI J�DS�P�z	'_ɳ�w�h5,���Z@?v��=0�������}\���|��3�����������3�'_�����<���:<���o�]x@?�O��y��?��9'� ��	<� �O�C�B,,�~G������?@����	�����p>��?Y������O��@ �N����'�?*O�&u�L�?IP���7�__��#�?�/1�����������~��"�?M~���o���� {���/գ�d�M� @	�m�L�d#�P�p����zd�����5���z=?d �9$/�s���i�������MB��>C'�����C���O�~�_�~��%?�f?�m>~ � ?(���'�?|>��q?�O����M���m��P,�'��?��?����'�?�~3����}$��~����t}�� >��Xǿ��g����������8'�p���@������ �O���p��;�L?6�'ׇ݄���3óaI�ܟĜ��I �NNf*�}&L>��;'��� �d�&ΆI��p6Mvy��,O�����2Nr���-���ѽwB��� �O����|�}��  @&���@�8�?\�Y?C�?������ �������}��C�����V?�~�a���������	�d3����w� >��5��d"��C��p�� @'�'�h7�ǣ��h�������>����g���z3d�L�t`�d1�����~�?����?�����ꜝ�a��� >�}����g���ϥ�4r��ԩ�y>�C��{w�n��i��%��xRA� �O������$�_������!  �'�~��8���������Y;o����>�,'���O=���8�.�p�!g�