BZh91AY&SY�QG:�]߀`q����� ����b3                                                @
 
     c�]ﲖ؆��a�Z4h�^@       ` `  ��  @ @                  �v���J� �R%
� )B��"�/�(DD�T�)QP��E��!8�7y��L��BiT��UB%#@���K�C�)^����r�T}9uTp�[�PkK�^���T��ѩ�r4���1.�B.�u�{t@   =�蒒Bo6��x�{�Y�� 9�y�US� �x�h֜���y�zϽ�ȥS���_CC�ΐ����>o���:   ����IA�mPUT*R�DR*]���>�9���:{�<c_|�y�̀}���_ ��|@Ӑ��c �y��g�>����e=� 9���}��  4�������](| >����7�6����s��+�w���s 3��� ��z�O@�9Ǿ�t�b�ѯ�΁>���g�   �؛o�%P �$���%"@.�*_ ��}�Jyƽ����}����x�W��'w|�U;�owA��ѩ�}�@�}s��_B���`�u  �k>IH �=;�Ǿ�� �Gw�iK�Y��=�z�iް>�{� A�T;�)͑�4}�N��T�|�Ҡ    �:y�(�����JT�"�* R�*���P�g���|���W��� �tJB�:�s��B�=���1���<af���w�
����vp�G�0>   ��u������� q�� z��%vx ]�O(�v�����3�ȧ��=�F��K���uBvnf�H   �t�m�A�!U)U	U)�j>��q�`����q4P�{y���[���нj#�nc����0�;֨K����}�y�  ���%;D�}�>F�@��ʕ^ c�a#����@�{ ���xz&>�<�b����cȯ�J��P � �)   �4i0R�`      jx@��P       �Ѫ�1R�`      l��)��       �H�%)(�M4� h�	��oR�PީM12T��h54���2"z'������������K�'��s�^���:�J������I��$�$�?��������Y�D����������i�g�'��S���?'��8@Ad��-���ԀA�VO$��X��dBI!��?������V$��ő�I8�b�LTGT���Db�����*#I��RF,Hő�LT����XŌTœ1c1d�LXœJ�LTœ1S1S�I����c�dŎ�b�*b�*b�*b���bɋ%XŌTŌXŌX�1S1d���,�SI�b��Œb�b��:�,�I�b�)�b�Vb�Œb�,�Œb��LS*�LX�1LSI�b�1LX�uc��1d��LT���$�&*N�b�8�&*LY&,�1d��1N��1d��,b��,�I�b��b��Ւb���b���VI�'Vb�8��$ŌX�1LX�1cU�XŌS1LY&,b��1L^��$�Œb�)�b���$œ���1d��)�$�1LX�1LXŒb�)��Œb�1x�1cIՒb��)���b���$ŌY&,�1LY&,c�I1N,b���b�+�:��8qcŌX�1c&*N���1LX�1S1LS1jɋ$�LY&,�1LT�1d��LSLS1S�1dŌY1cU����,������������S1c1dŌX�LT�LT�\�8��b���b�,b�,��b�,b�,b�,b�,b�*b��J�����������F,b�*b�)����b�,b�*��LTŌXŌTŌV-X�LX�LUV*b�*b�*b�*b�,����YV1SI�b�*b�,b�*b�+�œ�&,b�*bɋ���������&,qS1S1S1S�1eY1S�LXŌXœ1S1SLYV1LY&,b�����&,�$�LTŌTŌY1LY&,UŒb�1LS�1LT�1g1c��)���1c1�Y&,�Y&,�I�b��J��1LS1Rb�,b�VLV*U�T��1I����IVF,LY&,�J��$Œb�1LX�1N����1LSŌSI��-Y&)��,b��,�&,b��,�J�,b�1LSŒb�)���)��,b�*b�1LY&)���,u�GI���,�1LY8��,uc�1S1c8��*uc1c1LXŜV-S:�*b�,�1c�uf,qc1LS1c1L\Y*�)�b�*b�����LXŌY&,b����ELS1LS1SŌX�qX��XŌXŌTŌTŌY��S1c1c1c1c1x�b�*uLT�1SŌX��,qc1S1S�LS1eV,b������)����ŌX�)���)�b�œ1d�ʱ�b�*b�,��*b�-T�I��)��*b�E1c1c1d�1S�ULXb���b�,b�dŎ,b�*b�����b�1cr1S�,b�,b�)�$�1�I*ɋ��bɋ��cJ��$œœŌX�LX�qqc:���������b��b�1c:�,b�,b�,Œ��������b��N�œ�������LXŌY��b�)�&)���*b�-S1c1d��)��b�1c1LS&)1gVLS�b�)�b�,b�/U1c�$œŌXŒb��b�*uLX�1d��YVI���1S1LTŝT�N)���)����8��b�V1c1LXŌYœ1c�����b�Vb�)����)�qcqdŌT꘩�b�,b��LXŌY&,b�,b�)�8�XŎ�b�*b�,b�8�b�,uS1Sœ1g��uc1c1d�1\Y�&*uc1c1S1S1LZ����b�����c���b������œ:��$�1SŌX��,uc1c1S1S����N�b����1SqX��uS1c1SJ��������������՝Y�Y:�����&,b�*b��S������������rJ�������b�,b�,b�W1S1dŌY1S1cN.)�Y&,�1c1eY1S�LXœ�LXŒ��1d���b����Ɋ�Y&,b�*b�,���'Vb�8�,b�ŉ�$�1S�1c'TŒb�)���8�Y&,����LT�1LY&*LT��X☦,b��1LSud�8�LSI�$Ū��ŉ�#&(�%Y�b�1bb����:�☦)���1LY&,b�V,�1d��LS1LS1c��$�I�1d���$ŌY&,b�1qd�b�1S�1LS՘�Œb�1LSI�œI���1LXŌS��,��b�1LX���T�LS1LXŌY&.,�LY&,b�)�b�*uqc�dX�1cŌX�1qb�b���$�1c�udŎ)���*b��)�uqN,b�1LS1d��S�:�LT�1LS1c�1d��ՌS1LS+1LXŌXŒb�,�I���1d��:�LT��,�Ȧ)�$�I��S1d�c�8�*LX��&)1d�D��!�#��A��,�ńb�&,�ňb�*�&*$��I��Hb��$b�RF*C�"1dF,��ISHb�:�1R�1P��1`����'�^�2��� [?���s6]��\��a���.SĶɪwԪ0�^�!�y�7*�˷/h-�X�V��%٣��2����\���n$ݚoh���Ҙ�7u�庳�y&B�"kp��K.���t�3n�:˅]b�F���V��`/V)����7oU�V��7I��ne�4P�Z�)���!� �6��B��5�n����`�o"�Q�U�ZOu�72�I�ww��@���Z��,̶]�ڤpG��4(?\w�-f �Ò��YK��0�QzCin=�)b�]�p+��t/vH̥�(:c,�D�4��b�Mӣgi(��f�"
0:��6K)m��R�l:.S�p3W�ö�L�w&��V)�$e�]ڛ�2�<;��pf7�j��yV��p�V�u�v�m�w��u��Z���#j�y�	ت���7�R�ۭ��ب�Ӗk|�s�
�U��V�*"&e"�����AE�X;��V��ÕQ��j��������5�sr11�;y�-����U�*�՞��i�)
�����*�ұ)�N�		̧!F;Yt�JYf\�F�2��,�ߕ�ڂ��a���Μ��m&��iD��g����*�DndyM�p*̽�e�)�%��$�`�ڪwOsR�0����̺4V)�b��<͌T��M#vo�whԫ؜c$4�������Ab�ۚ�����8횤�j"� 4.��F�e�ө�MTXv]�7E��rFm��U K��׭mAzD�&㨕S�vQ�V&n�nF�ޫkN&*�3����i^����v��h�:܇T��r��@1J�h{�ys����]Vt��찲�e����� 'n�^n��T�F�hn^�Qyz�nno��5-�V^x�Hb�WV����"���5���JYGU���o�h��<˱�CL��Y����U�m4lV�c�X�Q�c`̣��-�Kdf�UV%踆�wW�k��i�`��:��`�^�Ӫ[��-M���T���$\�qX6���,����AR��[�U��5F2�Ds\ �A����SMX�x��(7e�n)3pYAm�u[�0f�Ĳ�ԗx��e��!V #×��ڒ��y��f	�t(eQw�n
t���`�z6ؽ���V:�a��ҭ��:����t�E�����(��Y�Yy�+�n��m]�N���ot^��,�[z��S1�=b꨽ðM��f�Y�:��In��ܸsH�]U�4D�w���`wUM��$�#��w�*��1j�B��R�r�q�BY�uV�T�WSt�$"ٲx��2*���T���ƎbV�n�U����7]ve�Sr��ʩ�9��|�����y`����PZ��Y���ne�ސɐ]%�&z���In�%0�����2��ɷQ4]�&n���f�ʰn�8��^Q+.f�Nii��4wh�"�7z��n�{`�&`��y���.�ʵ���c+a��ڡ�fդ��#y��i����[dU)[��;�N\�TKۨ.�Ѳ���X�[B�kҭ�$�z�+�n��nY؃�q�x�`��6�*��2�正I\i�a�l�@�׵�jf��4Ăص�7{�$�r�wPD�U]ӌ��̄�8�R�ƞe2S�ŅR'ckeT���*���3)�h��QyYY��U*�2�X�2e���j���X�6�Տ]Q�mi{H��p���-Z�Q�̇u��邪��YE���nS�\۵Yd槬L����פ^����j[	]c�o@��Z+\î3,l�K/��������V�8� ���:"1��%��:�yn��m�4��Yj�.���(n�AO�"����*��o����[�񚶮���Xz4��w��#�wM�tt�V�䈘BҪ�s2�a;����CEk�����^�9EUƳd$ڪ$��j�H���ʧ�6��z�J�5]comТ*�V��ZV6��:j���Z�\�l�Tt:��%��!P��1������ݩT���wZ��f��;ץ\�p]ڶ�$��,�ӻZ��ܷ�5��6�	��ec��&7��̡��Pn�n�Um]E�ͫ�74ق����5���a�����
9�Ukv�4�����Ne<Ç0���F���^7��u�{J�&��VF[X�[�U�&�S�NEP̥���j�A�۹��+T3FeҼY�lr�T�ط6��*:��N�h�N^j��r
����1X��nk�[Z�J6O�j���:C-��N��GiT�V�dV�,��e���\w�3	n���]S�-����J�R�Q4�&�/����ҥ��]i�x�hh�X�2��E�J�+�����{(��EՌ`�XN�e-̅T�#pP�\զ��_���5��\`��o`CR*{�腖CZ��TE�ۺ�!r�\2���b�{[�j��F䱳`��[�U����^@M���mԆ�bJ�fn<�jXЅCETY��Z�X��p�j���xq�v����[op�MÃN�B]�w�u#oۈ���ti'dp�-����e,�5/�)ַJ�<�Z372�Z��U�uz�-z0&mv�����k�
�Sm���fP.]�ܷb����f���K�"x��,lU4���[t���֫�vp�R�4�mjlL�/=U�]V�O�]D��ޭ��&��ɭ�V�)�m�&��uTsU:ʫs.�Ʒk �ޤ��C�GUD/\�(���ba$R�{J�C^����S,����[m��c\���ⷵB���=��n�c[W���&���I��9[�lU�0�RU��F��
��q��7�{J�R�
�kC;k1b�����ś�����۵����Gk.��#K\`���6k;o(�mUi�5]�v]���.�݃N�v�(fh����ݬ�
�k��cg1�5�6�!9���&�����k�Ukҵ������N�9Yr�R��dUq��;�&^ë|v��MV���HZLQl���pl�Ugm&^�.f\��2�+9�,���
o4aT���c3t�!LP�� U{F�ck-[��X��+M�5r��57��7t��B�[cBre*��7�t����{3u��F�w���S���9��@�/09Oh2���خ�6���+�I���J��ٞנ�ܺ]^Rթ��6��$�Ct +}�7�8�*�7TN��%J�j�/R�ih��)�2�l-�N%m�X��.���fZͭyT�Å��#g%����++d�w�l���BL��Cn����J�v��������n��q扶$�{V��P�[V쌬C�1�	�fnø�N�՛(�o�ңWxC���&^+�����2��8ff�����r�]�:�˻�P!��l{��ţ��5����47����^d��-SH�	HY�R������#�E��d5�@�k6��m�j^Ԋ^^*��F�I�xkq�˙cS�Y
�mP���tF��ẙ��&��SFR�c0Unݛ�9a�V���jn,��FhܫZ�4��"F]��l�nEnM�-�M�����I�W���D��M�f��+a̦�m���#r����!��"�ܚ7U�z�R�ؽ���3�@��)�UqU?hVC�8��ʤ.j��dZ1X�uU�٦��`�v�a�;Z�Ƌ�f�ƳHN�.�1F*�����H�D©Y��[j��Z����ƅʿ�)��3Ń.��$�Fm�IUatm�xa��2���k�.��ݽ�x!�e���4l���gd9{��ˁ4w0޳�a�WZ�b�:��#|���WU.�wq8����LU��ͻ��w�%�Q�ܩܞ�~��h^[�.�Il�Y��2J��D7b���qlAC6噗B���e�8�˸o��X���J�V\[	�!�Ab�&p���Ө�OUY'u�V�PEX�ݣZ6�V�-�WpQ*�SַJ�ѷ����˺��.������ZB�tEj�P8ic�q-��Y�F`5����ÍVwv��]�*�7��Qz��US�08P��k2+�p�U��r�c��N���iki�`��Sp�i �lvTV�l��4���\eC���;�2=��Y�j9Z�1Uy�M�U7N�k�9�A���T2<�5�]֭u�{U'/f���.�^�f�3%9`�y��#�+�{,l5Cv��t�P��3
ØF�Zo]*��b-��vշ�Z1T�j	.0�o6]n�6����f��m�C/�n�V��Ǚ�]���";{pLĮ�+�s���2����P�;t�Z�$�,K2�Yu{]iu��)��:�ee�+��̬���:&�+يX��fC�-��J������BYɅen7����P���GP�Am\Ws4�hʆSt-:ŒeORGB�wu���e4p��X�oMس<�ɻ��QŠ��,��5guS2�a�z�/6�*��5���2�Ui��B�n��.�Vi�Ֆ)����U�3xq�N���p��rL� x�J��f�wv{wM@�l�4�Tvt����T���ao�5P�T��L�ւ�l���6��jQ�c0��M�5�.�*��r:r"����j�2�ᰬ:�N���^=�7�Q��p,�!f�z���ב���b:��#�C�m�s�kfj�ӻyvz2�w�Lڬո-�ZU���*��4Ucỻ�%	�[�3U�W�[Nݙ~n�Tj�d�na�+ea�	�Wo���ʽ�r桋,B*XVm���h�U�>�eD�e�����W��V�a���U�Mk.�0Ŝ4�X��oc��nz��^�lÝ���I�4w7tG]��U�ov)3r�����ݐ�[X+Z�2����.�~l)���K�p��m��Њ�(���5J����k�(�w�l��[N��3!*;�)�;W�-���N\�[�s6�ѓo|q0�h�YWm'sFJњnj۸�jœ\��z5�kh�)��Ia[�j�=�5�B�"��e���zլ����F�h����mcGRGǙ�0�{�麗��f�9��{$R��BAΉ���죸S0���]�Z�2���V�,���t�gA��Zh�+��Y������&KÌ-:A�k��3/sU�ɻ �7&8:�w�)IQX�o��<(�z�ݹ����k0�i���7�l2�;�r�&ح�Ks�C�1Ī�h*��}W�ח�``�~�KN�k+7kiҖ�����O>Z�rVj�)��)dc�&�f'���g�=�뭵O�ș�A�w-��k%
�L^�r��۷gw��v����m�x�:� �ȏ��"t�l��ZEe��������Ϛ����n��՗�<?%��Wɡ��d�}�:���jC�`^��W˷�ܧY����gD~�2���h�Y�M}KZ��_l��U1_4��t��,R�V�{\n�[9H���į�Q]���)+j[W��{JRMkV6����gDͭ�7\#5����
:jV9l�'}��� ���W�+�[7T��jF�}��.��g�t/�O��k)5L{\��u{GV���1��-h���~�dC��Z�5�K&����͉�#L[uLL�BS`�h��jn)IX��LŢ�k�L�ߏ��_3ݵ}W�h��I�
�˂V�/re���鯢�/���S)yN���S���D\�w���z�Oq��T+��^�ǉ���]�kD�_Z_(�h*%�v�g�q�W�,6��|�L�<�U%'$3�lr���ݬ�\�"έf�ow�[��Y�渪 N�ɛ��S�wo��ZMc�U��:1�﷔eZ|$��bu�<�l��B�J��P���/�/��RF_ݚ��&a�T�Voy�̪0��Ty+]����`ތ��1���2Ⱦ��x.J�V�RᰤZ�St�~���^)�JZ)��Z���c�+��(ҤF(��6��ِ�s6�չ�J��)�ҹW��<�<T_�b={����z�$4ڬά�1>�G�;0Cx�n��y�|�E��F���D���K��}�Z�^������+VUқ�[N���ϖ��*#/q����b�'�0�������f��B�5�^����܇��p��I.�'��Lk�oәJ�g#v����86��}��2'&�d�?~�}�tUd�X�,���֭�Dۼ�������JJ�&&��	b{/B܋.���__�٫�����9`��hg�+���ź�"pݟf`�;;Ҵ��f�[qnK�f.���r��'�(.�ov��]������,s)1fLr��F��Z����Z(�X��bW]������TSy��H҂ɶ��؆M��I%t��ώ�ӭW���ᆰ����#&O��S)Z=ܲ��ψ���ɱ}6�]8��=�^Դ���;R
'����f��2�^Z���:��5�+�\UIen�gv~��~>]\���̎Ո3�K��v�l�x�oڕsj�Nn^�E2 퇮X}��Äأ�Խ�?P��|�k"eu��3�����}s~�߾������s\5�������p���U��{j�V+�WU�F�^�z'�O�]��^���%�RV��Z%�=�Uہ����ݣ;�j����z/9^)�V*��H��<�/���k�s2�]���j�1���ՄU�V�<����5�kpC�����e*��]�ҵLMV[�����M^l�iW0ZGrx�ۆt��v��خ������֤���Ǜ�`{-����SZG��nh�Q,�OqYuZ"k[�ի��&e��ƃ��
<��i�i��7���o��u1+ﾔoc�f�������h���]���̩�]�-ͧ�#ZF��\�������&W��J�C���ix�ك�ۉ,�W���}���h���Vi{6���D��i6��8$�V2U�	HULIO�5U��NmVs��̛i%�Q$J�)���HZ���ԯ��-�����j�����\�/�v;��R�v�*:p�n&��V<}�soۡ����]�Ë���6N,Kn�̹���B>��\n�^��dT�k�f����T6�
�k�(�nc��y��u��&�	-%.����PT1�M��k�����;.��vt����)T�'�$��yB:�w}%3/x�����]�k#d��]Y�ڎ�Ec0C��Z�(��'nJ4Q�2U��K%�%[��M�B>Y�ެ��k�ʫ���j��Vec��]n���Ƈz}����Z43��u�DR��r����$_��-_������o0��?'�I#��	jd-��"KQI	?��I��	��T�Z�@r��A9b"���(()$"��$!YKdH��NXBؑ9dD��H[-!-I$[$�-$��"Zb$�Ör����$I9d"NR!iTE��9a#�ZD����B��$-�ZKR�X��"I9Rr�HZ��!'*I�%�$�"-��l�-BI��� Y �!R��d�-$IjI-���D��	R*I'�����f��Y�O�r�����G�V#��!����ġ�ȨB��KQn�[�K����͜pT�ҳ;�y���%��\Q�Z�6GNx{by������ԛ{ч@�C�-@�(��0��>EX�GJ!�R�b���Xm������_bƆL����L2&�	��&|�AB�0���wWW[J��+,\D��5#��R6��ۡ�}��~�R6>y7������Z#@�CVN`Қ�̪v6�V�����B��Z[]�|�Q����y����e{A�4-�}��c����}��(j)3��Y�-p����Jk9��m�͢e�'І��HQD#a"}u͏�š�� �Q8�Q�a�lA����d^� �H�̈́1��Leؓ���fRe8F*6� [���;{}�g�KĽJ	"d�/R�n� �&��(��$�B�*f�T��È�H�H&$&G"0FXN�:_>��D5��"C-�.[L7t%�{�`�R��m�s�ݧ�߮���THF��Ӿ�"]�Q[�ƪ��!�.�Φo
O��YjUQ�I�V��a$X˪@B�$���u(|l�([����<����x���]jhV�_����]f -Ȑ��}��Un���[

#'�	��0����8�(�u�X�T(6N�b(�d(��S��|Nq�d/B F�d!D5���ϫ���3J�{߇������E�J�q�g�s`�숴��L��D�L6�ְ�Kywf�L�(H����B��Z[]���}���~�>�C|0���7G�]qhhP�4�y�}�n�[i��t�"Rn�d��:(���Ù�fm�k=7hK�Yn$�e!+���{�z���:i\)�r��D��$L��"��th��ٳ��da�'���KP3
 ��u��� �f��2�X���慙\Q�Sna���k��gĖ�P$���P�A��tBd���dMx��t�_ ��`*��:h�EZN����V���Ȕ���XV[
MfL�8
�D�R����0���I�̂�SE1NaL���I(�+�2�⢛mY���p�XID5�SgJ�eډ�f?����n�J--�09�j{hY�ѥy�%m:��qb$2�!�ϸ�M�tX��Ga ��`��c�������N?+o�5
]�	S,!]M]���YL6��K�2_���gy�S�"B/�?�<�$!?���������?�?d$'������?d�������>�O��W�ϡ5�!���W0��B>�3��L���l����S7�`G�I�z+�����X��r�,�]]�ͬY&T�N�Τ�i���+c�t���\R�X����5���󎆷��!�Q�����D5Wˍ�.�:֊�w��m�v)�\ �/�./h�bͩ�m�Œ����d�+8k�ϝΣoIn�ms������I���c�=AɃ��y���m�Xmv��K�9��v���[�b��*��t��e����m�;1�ع����q��}VU�8N�'ut�9�	�lMjxcg.���J;}G9d\�z���1ٚ1����z��a���1]h�І�hih򬮵�Ј�G�I��j��z:�$���+�IqU��t9j�l����l��i�9{�T�6���Wt���.�*s�M�F1�i��N��v�;�k��9�;Q��!ӓ;�:w����Q.��r��-�p�<5U��/���{�"��^�̬H�Q.�O���@���w���I�L5�8ne^�b[SIܪ���e�����V㽠��"$=�_�����ޞ��:���ƵƵ��kZֵ��k�kZֵ�k�kZֵ�k�kZ�5�k^�ֵ�kZֽ5�kXֵ�zkZֵ�kXֵ�k^�ֵֺ�k�ZָƵZֵ�kƵ�kֵ�Mk\kZֵ��j��kZּkU�kZֵ�cZֵ�k^5Zֵ�k_�ֵ�zkZ�5�q�kZ־65�MkZƵ�U�kZֽ��u�kZƵ�k�Z�ֵ�k�Z�kZֵ�j��kZ�ֵ�kZ�Zֵ�{lkZֵ�kƫZֵ�{kZ�Z��u�k�Z׷/���o����{��B�"m��Z����O�.z��X�L�q�lf�4�Y��7u�7L�Ŗk���9�|�.Z�x�Xt�c/t����n�^��w��J����ݬk��5�!��(3	7o[�B�Y9s���,��S׷�+��;�W0i�;�swrmk�����/ml@��6(���U/3\�u�Օ:)In��J�Ksw؎���Zڙ�uA���ד1ޥ��t�p����p.x�n}\��EU�[B�a�Usڼ!�+����{Y]�wq͉���f�z�n=�ӓ�2b����N�ʒ����"���y\��p�q�G�T�wv���\j����˸�b�W��{�/�7����dz���*�hA�a#�ۺ�Y���s��A�̈N�3s,^���x ���rv��q�TX/���ПenA��'����d��΂�/"	�6=�|����!ӟh�˖�5�pMx�Ӿ����"�fH.{ޣ�{�7q�ם�b�XO���D��-t퐥Z��ں�ɝ4h�wc�I©wo.+�VsU�^��N���ҨϦU�ɼ���lkl�����kZ�Ƶ�kZֵ��kZ�ֵ��|kZֵ�U�kZֽ��u�kZֽ��u�kZֵ�q�kZֵ��kZֵ�x�kZֵ�|k\kZ�Zֵ�{kZֵ�mk]zkZ�1�kZ�ֵ���kZ�ֵ���kZ�ֵƵ�kZ��ֵ�kZֶ5�kZ־5�5�kXֵ�zkZ�Zֵ�|lkZֵ�kƫZֵ�{k^�Ƶ�Mk�Zֱ�k�kZֵ�kZֽ��u�kZצ��cZ�ֵ�k�cZֵ�k^5Zָ�|k\w��P����Z�ȝ�/�uI�7Fٕ��1ef�"��uð�{�o^vM�.���ҍ�bU	�z�+5�1+S*
Z�����w\:L�� �nͼ%=T�<Y�񩄅u�-4:�Kk��s*�nn�s�ڤV=�VA��5ݪ�gqI�0^���ËhŪ��mD��'6{kJ>oUT��)�e��$��^$��+����w�*L<�ݲ��Œ�f�ok�ө�$=xn�Y}�'`��h:��pQe�Wb��j�m��c��o�,\�mڳ����t�aVQ��)�Wͷ�]s!��4v $�5�u&]jPh:�Y�{,�SJL�v,:+y�`s.�9��fR��6�P葺�t+�nj���P�0�}���gWnA�������/9a�V�r���';����B�i珮]�"�_^fb���Rj� ����`�y�6�g�ͨ�P�\w������쎺����wq�]�r��]0U�(��lN������R]FRt�Q�hb����"�˼<�k�|����hʪW�|�f��Px ���u췞�X�O��Y�����gs6����V�L�zmkz�P�|2D�Z�B<p������������ֵ�k_ֵָ�k_�kZֵ�x֫Zֵ�k�Ƶ�q�kZ��Ƶ�kZֶ5�kZֵ��kZֵ�kZ�kZֵ��kZֵ�x�ֵ�k�Zֱ�kZֵ��kZֵ��k�kZֵ�k�kZֽ1�k^��ֵֺ�k�Zֵֺ�k�Z�kZֵ�ֵ�k�Z�Zֵ�kZֽ5�q�kZ־65�kZֵ�U�kZֵ�q�kZƵ�k�Z��5�k^=Ƶ�kZ�ƵƵ�kֵ�Mk\kZֵ���k\qƵ��w�kA�����x���+J"��/6�}��vuۺ��B��a��T��vu��6q�o{��S���	uBr�<�qb�݈�6j�FЛ:�h�J�R�vAI�
����;��\E��on�&�U>;I�+Ů&Q��υn�=��+�On�UTێ�oby�vY�R%�M�]����̛%u�m��꽹�o2�vq�5�+����j�IU�+]wI�-�r2�ti� x4̫��͖;�j��²d�!;/�܄N�h9�TbJ���b���&	�kXV�U2/<�N�f;MܣB����b��-�Wuq�lZA�7!'����дk��M�o9س<�>/�#vZ�hV^p�n�|u�Н��Y�ܙ*E�j�أv�ӊc*����O��E%�.��n�V5j�_,+5��-�k.5��ڪ�*9nV�ǈ���ݮ���ڹe���Ʒ�Wm�3�?�g�xD��B����y�nL��k��(n�k�u'��Mt���M�l��Ip33�+N�f^U��Y�E��X��دW	9�MbW[��T,}wH����O&33#��w����><k�Ƶ�k�Zֱ�kZצ��cZֵ�kZצ��u�kZ׶��5�kZ�ƵZֵ�k^5�q�kZ־5�5�kZּ{kZֱ�kZ�ֵ���kZ��ֵ�kZ׍V��kZֵ��kZֵ�lkZֵ�kƫZֵ�k�Z�Zֵ�{kZ�Zֵ�MV����k�kZֽ��ֵ�kZ֫Zֵ�{kZ�Zֵ�MkZƵ�5�kZ��Ƶ�kZֵ��kZֽ��u�kZƵ�k�Z�kZֵ�ֵ�|k�]k�kZ�5�k^��k]qƵ�k]�������=�ϗ̤�-�O��uIh�]����	d�¶���`Ļ`��F�ܭS�uiaS�L���Fe�\-'L��j��[үAleFj�7튈��x�@���V	i:�>�ǸL�i₴�`�ͺ���x�z�Z�Cp"p��Ã/�F!;R�[s��;}��EGV��[�w�.Z��d��x!�M�&��˚h5�b��Hf�7UF���v7\Qɐ�;ni���{*l2V̂ʱ�-JSq�x�gT�U�c~0���I��uۯ���̼�[#��"�l�3O�r��ݦ�,Jt�����<r�s��Q��YrU)˷P�o��oc��:�S�T�m�ᔪ��uL�#:3�fAέ���w0�}�]�ض�4{���鉌=x�3Q"RX�d���อ}����G�p�t69v�y.��2�i�D��r���:�əIX��xf��v��`�dx���;�<%�uCO�������+��pĠ+�u�i�n�2	wo(�v��6Ù�8𗎛����-I/s7�v%���w� �%���U
=y%,3�̦�&`�Y�sVgev7[)sW1�S�Ձ�U9���f3[�2�/sJ*����l��z�M��S�o2N�7�oM4%FC�;��;+�íu��d&�n�u"hY���1��{�g���W#��4��.署F�aXs#Fk[����7Q�^�/V��KUu����a�p��.��v�4��)�=���<N3�c�{Pr�Orn�wO^Z�q�yl�4u�
����TluX� ]t/]��R����������%ȵz� ]2�G���E�Fwvn�
��2�kҝ�Մp���S�y�PJ0n���m��E[N��^�Zb٠�{�����=���0�o��V����_T�3_ݘoh��t�77p�`��� ��']U���pN�!%mvqO,[�X�� ��'[�1kUG��r�=���gwG���Cݚ/;�rg���7��Y�F�lf�xB�y�G��<(%U:wD�Bk�C<'Y�r��B]�笃:�V�5w0Z�b��Y���O:��.�Wڤ0��)�W��3�	M,����Y�˾4@~���ε&o��"�e��ك2!�.9F`����zU>�w%��`xu�&�'A���s�ͺ���vF����qb��%y�M�-:�'.|���l�����[M�ZH��`��r=9*�ټ�J���!T�2��R�Xwz��mXw���VL���0h{[[�u��J�\6�X�_J�o�_w�3������ɽ3Bz57�c�F�iH^��㯌 ����U���e�]~�Wf����5˪:n��^՗�3��u5]�;-�꺰θ0�}{H۳��X��u
�3tn�WV���^ڛ�4-`ܴp��c��j�D���<-U�RիY�3u]8�� m%7d,,V`����� V���������l�uUz)��%��Nݷv��;e�C0�N�;�Z�J&����^��$8�쮚�s.�E�ƨ��֝c8K�uXR/9��#L��d����u{S)��� ���o<��/.�����&�3����TW\�w�aY<��{��[;��e�v�%LhZ �m�D�egb������Um^%���f�:�h��}ZX5{ݴ�]ow^ �R�Z��۽���+[ƳqS�u%����� �j��^;68�ͭ%U�)��]�slj$o��w��;'.nYN^���)ޮ�dәf�o�վ��:Q��W��=�UǵqA�ʙ���@w�O͊ňǅ=7�
-�u���q�[�y���wVڥ	�5���x�yW����\3kgkO�����h����f`����ʼ������������M�V�$ug����i��ʯc4(�zqǸV5N�e>���7���r�d[E����n�J�zws��JR�)Q�vZ��n96ŽU�^���U�^��+=�Ĕu�K���AW��'j7�P_bs�8V�8��=� �"�Y¯.��v�C��{��Y�R��*�Uu�u�V��e׼"Ǳx���{d�.�G䨓��7�T�Je����^�����Q�t�ĺ�Ww^?{1�z��Q���w�qus�3P�j�S�$7�uV�=�uf�-�X�����}~���ۭ�o�N��y�]G��L�-�\���|޳���3�R
_��#�㫹V��i����O9�Wf[LT��T:�'��bï�-;ә,�v@{t�yw����/f[n�J� �ӯe�<��)��;s��ҩ�oAG�Km��;���q;��ݙ��{.ꉼ!�hM�R]���v:�M:R��{t����]�Q�6��J�N�}x��"�1������S{z�o��V�v��#Zf\��X��6����Y�����}�w&���7Z�Ql]"�[ٚ ��Y{�UQ3z�hŝ�/��Y�t;�WLٺ¥���M\)��r���vi˲�FR*�x�;�Yu��ǩ��ϛ�g���������C;���'>�ou���cŕ�܃��9�f���*�T���7��']�8I� ꩻڥm�b����N:TDw�����*ńU�&��]�I'U�ϖ^��i����(Mӓer*���4��7��<�>��6:`�壋���p�"�+s}�'S�#��0o]'�1e�>&�7��rB S��l=V����m����v�ݠu�h�v\��۪����mQșO�U*�:���eմkep.���B$�ط_][^��3ލZZ�7�sv��Eɞ��L�M��֫��ad��n�:��i*������C/�k;��J�{]FR:^nU�YS{�<��2�'fKP�|2U��_wj��CM��ة�"�*�R]{'�ҷd>���\�����h*��p�� ��Mܭ�ͪ�Mb�֏g6��ͱ���h7NWqH���5��mbN��]�b1�:���L��ϴ�,Z.��������ms��v�D𭻬���X;(>�p����y78m��szg\�5�Y:�\���M�c"P��nR�l���5��w"<����a�w�+��םwIa��fÕ�85��V���g`�s+W��W0�ckl���0�;���I�v˺�䯳Y�{���q�&������q�C+��ܺ��xo�
�kH�U� r�p�vVZt�fa쥙���Y.+�\7u��g�]�M;�Y����ē�M�6�oH�.�q{Iخs	�txWm݇{V���c�nn��ҎV��8�ꈺ�f�&����VU�ѻ�-=��K���ܾwUd7���+�M��jS=��q^mo]�skh�L��́���ɘ��a�eM�]�k)L�M��oH�̦QlC/g<θxw3 �W����y]�[{����o��i���˻I��쥖��K��{�.Tsޮla�Y8�
�ĺ��*��,nY/y�Wlzr�eUzV���ʜ�شP�w�U|Vs�X���udom���bv�\�p�R�g����,ҫƫ[��%W�B����/�?��������������bH��������/����Q��O�?�t�@?4)�!ϓ���Y}_�� 0	��K��량���[���}0D�ؒ�i��rj�_v1|�5�<z���xf�D{|��8f/&
λ��I�,~a���@��ڨibq<]��Aȣ�9n�
�f5�%��a�փm�C�X��]K�/6�������mx�E�j3E��B�ΚMsC$Fd��хs�,��
�D�j飛V�7B-�jm#�ULY��lZu�L�aU(�{��k��U� �1M��݉`�6�J�]�z�$.j�kD�����F��(\����7uV�C!�VƴV�i̖���Gv���͗���ă4����m���4���%�G0̲�RRj�i�fQ/S]I�m�\�*�&�Y6q-�T��cM��a,qv̴�e	���i� Rmٌ��Cq��\��l�i֬���c*7B�S2�e�)�GkJ�V�k���a�V���Z-ʛ@�All�m�]A(�����.r�4��7������0���cA"6�&�t��15�2�)6�m�k	hl+J��� ���c.����j.*�P�J�Θ.K�z�-k,4fR�r���L�q�6[-sB9��`8��9ñs��Nٌkb\�4��`u��rh�h@�Ɖ�4ұ�fP�hT�k"�c���˵!����\��Ku��:�%X6\����ƵHi�dD]-��ƹ� �X5	i�����Дj�a�4�8�f�n��b4�me桒�%�)�v7XiiN�%̮���72�t�y&�����6��E�U�͖Ն�9v
�@��4���B�&֌en�c��̊G���mD�d��@s�R�h�]nc1�Ye1.Fۛ
���f4�����"���)4�jh��D�:[8��U.evb�Kc�Dbj�cn����0� �\݂d(�@Ԛ�v�V��Ȓ�H�:�ٛlaMP!�;��V�m�Ss��͛�5���̺�4ΔhJjb�Kb���FbG�2��2Vl�F�ꑪ��]4��M��t1]�x�F�
�tLܒ�&�#�Z�k-s�M��E�e+�cIl���Q��B�K,km�\;T��S+5�7Rir+���Fj!��k��؀�R�W3����Jؚ"<����&�jU���b�Ͳ��\F�inB�b��� �7M`�M�ȋ`D��s��6�[�t	y4�n�)�@й�7\R��#���sM.j��1n�LJðut�[.�(u�Ql��z��+/&&`�+/P#��[k�gX�K1Ake���i ���&6,ڲ�ե�ЄH&���0�kiΡACs��X�Q�ֶ&oSl�J��ՙ�U6��uѲ�	�<M�Kn5��ڹ;r���qLbk�x#�FĴ�F�/*�T�*gi��0�kS�vI�U�!�X5���`Z�[3
ֺ\�C#6Jً�h�aY���{H:�,��5�sJ�VӶ[t��,%��:�&�nx���YaM;��J�TU�Хta���XGZ�lgV=]#,\ԙ�ķ,!�2�!L�S��֋pkPm��1R��-]�s�d�wV�e�eP�&����K��3[.V�9�j�,t�G�m47��,�t-��lP�R)��Vd����:�Wcq	��ح��@�cSR*C%LG1�v#���f���� ��:�퐭�g8��]&�Up�au�6"B%�ҵ�#4!��G�a�r�It\ge��Ώ#P���Yi�݁�-���L]�ۋ*�3�.M1(��mW �I0���.����a.���9(�JԎ��a�	v�k�:jr����ՆP����U���
��V�3`c\��]
l��t���i3Hh�B��\hg�#��cI�p,k+���Dn͂A����Rv�2�b��Y�E�@���Dؖ�c[�;q�8qe�Hf�-�eH�c-����ф�cqqm-�IiJ`8����U��n�F<ʬb��Z�qxuj�4�W��eDLX!�`��z��h�M�L0��#�رU�ISL�nHK�iH�#��؊S&!t#4��dR��#����)m ��f0��-S�YJ�K�Ê�%Łn�\��w-ɦ
lh����k�sX�jʐ�1�ܴ̦۠f%�՚�r���b]i��ج�Lћ�WJ�8]چB�9��Ņ[�p��݆��1�����Mk�v��1�g��m���-�Ê�R�vft�:$baԣi,%�B�V��&ō^��!h��uc��\6���j�f&��+�v�(�ۍT�An��7S!��2]e�יf�)F�����`�ºb��[i�0̕ɐ[��͖ew�f!�䛭m[ʎ�5�����˴�f:���Ѱ�adD-��6ŅlV�v���VP,l�R���f,��lv����:���Ͷa�DA�ll�Fm@�lf����\ Ķ�c�)f���]x�۸5��� L���\�PSj��)�Z@�
���qrVf�6��YiVj��j�c"Fh&4+c,3n@)9�����a�YMԹ[,f
7�2D�T��.��]�;�8%�RmGg�Ѣk[�J�Ƴ5��ZƄ.,4Ƹt��a�l��J���+j��f�n`��N&��،)�6��c#y�^ŭR�@ؠ(i�nWdAe�׬z��תG6am-���[+L��e�5I�t��Վf�+J�����ꕢ���n��hj	rf��*��h�����5[���)��� �K����E� ��+�,�7]q�-,J])��%�-f���Z1 K�8)%ͤ���P�M�cuhbX�9����6�mt���t�s��й�3��R���Uf�	�MM�r�h�
+�ٮ�W�m�R���]Q04���頙��V)*I�l�b��[`:���qvp�e���ڐp�J��6k�+����k�@q���Te)�����XXl5���PU#�[)ne��V��rHYv"��8n�Ka�p�ЦWc�Τktf��`�3]��I�čm�oi��%�k�a��� � n�,�[6�ó�i���4K-�my!f��(j�D��)�p1����fp�̤��ԳM�.�x"���m�J0����`�����ήځ	t)a.��Bh�����MaH�7{:ȱ�L�t[+ں)*����R���-���kcfk!X���awbP�WN��/R��u��h`h,��e���VT��ms,8�W���cΰ3C4�h�Ile̮��kĻ&Ȓ�(���-����)Pk�X��V��큺���7X���.tR�V�f��U��m�JZ�R�0�;���*ٛ�#Y�<Z[5\B�txnvK10�T�tl:���v���Ջ-Չ�ͣ,E��	s�[F��;kb�7CY�c"�l��3q�*Mqkr��"ef��6��FQ$��e�V��N�ƥ��6%�à\8��taZ�#4R1���r��eݣ��h\A�P���ֈ�c�P��[�Ue%��g[����&��Qj2\
�:���y���.Ih�A��9nb�f���;�3YMp��ٌc]5����Ʀ�*%�����2�ˡ&�sn	U�����P�e��\]SXj�sE)laKmn��r�,��y�͗"p��::�e^���qtn�h��L��4��\�`Ɂ�1�0���,8�ne���8vj��\)��mҐX�5�:������lѺ�)e�fl������٭6c��2�U1�Ү��m���7e1��i]� �6(�����o��,!�}Zw2�Q�S�����I���)H���m[i�	���:��(����i��2I8���mPp2�6A��O�
<YCx��O�z�<,�����������C��+2�ե�)�+��:>Y�-�kMW���j�d��F��m26��b�l#�:k�Ȱ��} b"�ҭ�q�qep�>`X7+���!��<JHB�p�r��-�|���-�?3���|h�?��h�����j���Z�cP�m�Z#�I����}u����[>5�Ǐ5��kZֵ�x�kZֱ�=�^��?|�y�qP,,�Z[
���uv��6y<�N��w<�O<xֶ5�kZֵ�U�kZ�qT^��Y�R�U�U�^��E9�rc\�R���	�׏5�=�x��Ǐ�Ƶ�kZּj��kX�/�I=���9��yy�^��Y��p�f�H:��!?S�@&s�߮�L������Ƶ����x��Ǐ>�lkZֵ�kƫZֵ��W錍s+r�ƵW�YEF���2����f����<��jK9N�ؓ�GfX�%(��� D���
I�3h�҂l��1̸�`As.1@P�p5�!#iX�Y�q�P�^��nOq��^���2�edU��a�[2���\�Ę�R�B!�!Q�����b�s݆�-G� ö\��UUar���d��b�i�I �_��nI�J�J����h��L��mSQ�B�K�sr���I&�8 ��N�m/R�IC�D��1]d+�q�Ӥ�aKF��M2����B娱�-��{���06��/GbP����W����Еyb����m)������	��Nf(���.)��3KLJ��."��P���N�.�i�y�͵*"+�2���9,���׭�x4�k�K@�Υ?K���Wβ�(MH�����G��N{�����dwes�ج�=d޶������pS؈��4Xs�D����1��dڸ6Rk-LF��B3,�1�:4�*�-IH8�
撕�&42�JV<*f�T%��kb�����啭ƒطZl-�u5a���/P�
��(�h���[��.���6h�)�xT��\k�i������.�+piZ�.��f��v��X�#�tnى3eƢ�ֵ�#8����YF�۝� ւ�:����l���f�(�+��ep`(��ƺ8IE�Y�t�+��-��&��]���XX��&��D��49��-�����kP��
2�K����EŊ�&h�]���]�5��.�n��lkK��J�W`��a�ܘ�Fk�`��	��h�6f�5���Z�h¦�j�4I��	�2k%mHY�&-�4-���l�)�sd��J��(v�K q�7b�l���Z��0�8�4"2�V$V�[2�ۡ�4l��i���2¬�L�4�!� 	a�]�[r�jRWFǮU�<�<��#�F�"��Ў�-M�L/jb�i6�3.oa�1�2e���8r�EY�
�,�f#����R�ݚ�mR	a�[�̶G[�3P��#`���^ΣeX��,�835Ō�p�E����
,���j�*���\ih��+z(��z�]��'�oR�5�e�t�c`�i�ۦ��u���\Vi��r�`�*Ѯ�e�Y�����
R7:�6���J��G;a6V�1�j�H�})(V�V�d�)��bj]}�XR��3��r1�1���9��}8kB)�b�21[RQ)-m(#Yh��6֖Qh�%���m�,:�zʴ�z��7�K,���"+F��K�0[z�R�����ka-��VP��¶��{ R�/@�lP��p�a(eX+i�dDC�H�Z*R�V��+/������H�@�ǉ ������_m(�t���r
�}峪�'��o��Ȱ�rP��Xx��\�#ǉg�x��� H�F�4�|�5�m�NN
���Q����p8��W���|��/�cm�KDБ.���d���@y��s_i�E3�swu�0a'O���W�w�_��֌���\rJc-�H0�ƫ��B�Mk�[�J΂
�I�}׫D�%����r^(���ޕ��;��m��3'���Ar���݈3Sv�{;"�Ծ������i�bd��i��
�����й���b!�d��m�F6������%��:@9 ͇dϭ斬|�%���=�����ĝ(�����!j"$�������Ey_��,yM=�G��f}��D̓+���h=p�����+m6�W��\$k'���%�UH�e��Z��@�6 �@c�ϙ�/���O�� ��w�Z�E9f�9M�� �	x�^9�H���Hk�s��U�;��3n��[uO�HHv��8RAG�CӞh�gV��̄���#�ӄh ��^;����^��sR�@�E�`�I%��d���Q;�<��<��HU笶���Ɉ�,��>gpI}�����u۟V
t`�6�E� c��Gl&��^�f3 �t!���D&�ٛVU�|���|$1(��'�/��Ow�J�B��E����E<6x_���V�d&�8}�T�� �����j1��_}���|�Mϫ�QD�1 �l���b�8�Ǚ��ll${�fވH_r)%�v���1��쯢$��.�y��oy�a�6b���f;%_K�����f;�7����^]t�_.b��F��eyr�^�v�UT'UTIVJ��t�ݿ3�������&�Ow}��̴���_-�n}��=[unm�����j��@�Ikbu�����]�_����	�ϑH����Î��؜�@���}�9z�e��j@�I��4���x��l�N�y}��:�Q��W�L��[I�����:�he��(ZWc�E�p��T��e%s�4�Z������-�"���Ϲ����i��n��P�'}V�$N]LPPS�r��Zڢ6�$96�!�˼J��"S;�$��+[�$�V� ����Ĳ��e�a7����`Q�����%�9c�8����F���K�c^�1���۞#ii��H/V��(d1C�~��\�*� �JV�?�,�I;��0Ҧ�;�3\� �`�������rlv]�>uOԟ,	P��n�rR�)T���+;�8��}��Z�>��[v�H��0bHyɷ��ݸ+{�{�>c�\��|�$�`}�y�������T�6������D�>�$2�2y��{߿��|�]��գ�pe�#r���fB\KI�UY]tsPǽ���)&��u��|�>'��oLS@٩���z�Lj��Hgϻ�D7��$-�"���{sA ��J�N^�l�X�=<iD���{5 u�	�90��E��	����FbQ6i�_@� )��6<-�����<��eઘ��[ �������s�$'��R�Kכ��УO4�>��,5� ��y�|�fy#��N�>=���`�߸ ~����E2����Q�L�8;ؾ����X�����]��� �P'y��Tg���Z�e�鐾�I��"9���.���[6�^���%ރ;,'�a��$)n�J�5oi�R���	u�t�ya���t�.�#K�-��E�#�Fj���8�;��0����(&���!�ؑF�4�a8�<(�Q�Pƫ��_x���}��'�Y�%��q�h7�Y��ڴB$�{M^7�T��ر4,6#t�fYAM��ip񎕋���h[�MA��p�cb��Ų���R�*-
�lىN��!u�s�Z��N�Bk2���Gy����@��h��Vb�fk��^��2�/M&�Bc]D��.J]kA�B�j�l[s����$1S%�\�9���nK�o3�-��_��� ��� �km>4ɘ��oh�F�|ɠEU1�K��0����%�>;><�l�t����k͹$���ۺ� �ʲb="?����8���[JE��z}�P�'�{�7�//�հEU�w����d>c���!��A�8w�Jh�w�*
J"������q�|/��*��D����D7������#U�<��
�� �ϯ�H5�F��g�G�`$�W˧���Kg	����^K;��^�_ɏ���o3�"�H��+�PUm�ၼJ�K������
��2
P6S9�}��)t%����BX�L�3��6�Z�͓�O�Lڳ����U8�K�+�f5�-�~�đ��+�Pa�7�Nu����{�Dz�$fa8�f	�N�X0Zҷ6�O߼���'}��옩U*���{��㭸H���9���t5�a�3UP�|��(B
P����ii$���Őwz�|J^�l��� 3�^��I_y>l��O��.	R(���2�س��\;��1}c�8�w��b7��F���z`iy�ʼ<�P]�z�f%q�:w�i��A}�Bg�Ȭ߮��-r<���ۚoSC����d�~E���1h##p�"�ߞ�� �4�H�a�F��W8�J1��V1��}�|A�
4�X}�O��� �~_g�A%���#|A�}9��P��,@ݐ	�����c�x�o�uU��o��čԂc�w#ٲ�$�{]�'|<���� ބ�[޿�_�rP�/�q>$��䧐��op����v������i��=b/+�ιD��繐El$N�N��6�\�\e{J�*�&��L����r���*yJ��-�N� F1�1b ��e�1|�A�dηu"][Y������醾p�6?�T��&q�D�grF�	:���xk|�������8��I�{�	R(�׷=G*x�@&oS)Ov�4����M-�M�AݼRe�h��b\j}ԕ=y{F��P�%�)��1�X*d���v�[Uc5+�5i0`������bQ��|s�)�����	m�HÌ�}>-�H m�SjO��^j���I	������N���@wU��ED�B�l&"ښ3خe�a ��?
AVDb��!H#s���������ye��b�	1����%C�B�RԀ$��HB��{н��G����d�lwo[�<�/��C�	T�Aƺ:d�uu��Gn����e�.�p&vڸ�%�53�ž-�L�ܢ)J�5^7;Nur����ͼ�YB�^KB����'�]P��W�w귻��2�Q?�i�D� ć�c�>��]�n�P��C=^@"<ɢ
m�R�ǔ��&,������w���U ��'oE�e��Ba��%�Se�Sٜ�늯T�����۴l��.]eл^]h��|����ڑD�� �3~����~Ht�7�̯��9����P������t��9�.Ch����礟���O�����X��I�����	����3f3��P~u�L�4헟}>�8H7�9o�In{�q��
גߏ�g��~��jAU6HyD�t�H��i���ݙ�*4[�YNG�d��#>|g��t�~y��������b�6��+_�KK�i�g��y�Ӎg�R���xvY�S��������y�+�lG�U�|.�ań5T�h�5�g:��Cz/>.�Cꈣd�q�f��U�.{�q7��{�e�lc��8����XD2f)-�WB�&�"�x3��7@�x#����F_W�����`�c.�J(�I��6mNq�g[fmUL�da �1�/1z�e��e�/��������Z�Mn4sIy0�L��0��&i �.�663[��6�*���6�c"�%�6�iM���f��0;M)�a���Z�h�Kl1�lx�:�-z�ժf���`���\��3���%åHaf.��ԑ[�ِ�B��a���ώU��~c��щI�cM�]��8�F.��C0�l�]���H�����8�˲_㵰B�����sR�>������ ��d	>Ǧ�`�[ِHچB�.w�1����}����E�d��Hi���듟2��Ս��NWɴ�LH���)�M(	�mt�'��&��_^e����R��~�����>H_����%��x�|iо����2og�33|�����D!L���n�	#�k�,��44E�"��!�(K<�T:t<�F�-�.v)*�v�/��ۆwvC�}\�8;KND ��:F�yi�Z��-uf���P���m-�ڰr!�{O_�O6��7�_�"$��r�a�.�:�����Z�K��x@���20
ɼq�̎PW，�^�^_��a}�����"�g�D䊑�ښ������խ��tR+:H�Q�W�IwgV3����޽�,A�c�e�Чأ����dPw�z��B؊L���TF6/:H�ﻠ���ݮ���s��J#i�^�Q�6K^�-�y$�jd@��R<��i���.�k�|%��Kp�~�l��Pc���ͥ�9u[>�-�&6�%M��^y��<�I=����������I ����҈�����`!��&��-mk	\XW�X�]#f�5̮��v\�+ �]Xֈ�T:t5��<��U Cc>��� IUΩb��B==c�~�u���a-bvj�&�g�۲�A������i�^|!J���;C��A��@�AJ�Ty���3`��ze���|}2�����'k3�2�V-*]�Ho�Kӫ��m!���.�K�����d�v�����3Wٯ^x:�{��<��.��D�1^޶3w��u��faݛWc؟6��|q;���c���yRf�ۙx'Lpr����|3��Vz"��^��]�QŊ��*ɜFExO��"���Ӥua<7r��/1�<�^\���۷k:�es��y6��VR۾@�u�V]�=����44[%=����7�wnZ��#{ۮ��mƺ�&�YvЬ���빅Z2��yK���i�޴`�y�9x9!h���U���+.���9G�����7���ѳU�+�{�:n$�s��[P*�����2���������˕��칛6��cڝ��������ѫ��q=O3)ټ����7{����Tw4����̼!�a1s�N�z3�UZY=s2�r�DbO�Wi�.�#2���`��挪ޫݤ�뜯z�v�Mw�n��sK��rK֝���f��+��{�}z���u���b��Z��w&�*�fmV���i�E{㷽��ڣ����ݱ�!�B��a̚έ�/:�Mէ�w.�fp��W[C�������GS�:�˧�m���v�\5�ZT���M�|�}Ɏ#�f
�-�����9�US@ľoC�ұie�U��I���j��h6�H�DĊ:�	�'����׺�3�t��3hva<}A�`;݆���i��n�2��Y���zmV\ԅ�M�@�겳��r�Zm��e�]gNNXR��D�o2���JK�--�Ln[mV���h���j�d�}?L����Ǐ5��cZֵ�kZ��{=�̞΋ЫS�����]E�"��-�-�n���Z�mZ����ߜE��cY^����־G׊���Ǐ��V��kZ׍�kZ�קgg����y;{{b��B����UP�j��CwqF�K��E�n.C:�Og����|x��Ǐ���kZֵ�x�ֽ�̜�[B�2�׵h���'iPyi����f�1UAkQ��9om�����ƽ�q�<x�����꾵�kZ׍�kZ�'�V[l���s�(��IrQ�-8������Z��[J�7b.QK+o�gى�մ��QA��kN����Ly��6�Ѣ5�k�u�-�����\ �%�l,�%,�Qx�Vދ;�K��%��萕���e�+l����B�QJ!cKm�g�_�Yl.@�l����yx||�6ks�K�^��#ҖYm��,z�aj�+N��y�7�e�9�����lUTij-�eܢ��e��f~�.R���F��`����I�I=�ΒzRM݀�;��1b$��s�-��퀙$�fQחOiFڊ r�W{&��(�؟D3�I-�����k�Y^�7�O^O^���^�:�$5S�4�@�V_����ØT�(��I��lO??;2�������ۼ��P��M�O�{�*�2�Sœ�?7�'Րx��9`vD�
�5�Սi������}�濽�w�*j��ԸIkt(��j�v�oΆXU�I�/���p�O��w���7^��̆�ND�$������2$*$��ߛ?D$�`�M���@;���6�Il�?>��T�IͶ��~o>�ݗ;��z�e'���Q���}{�I"w�zF,��p�~w���'œ�LX�)�?;�DB?��ÿ/\��?��8��@�ӷs/�*��$:�����7X�"I=�?y����RN��_߾�~< ��}u<Q���6ΪNo&�~dOR���+L��F3XO#rs|��nn&�od���Ck����~�,���|�H�Y���r�	��[�N�e?O�R꺵�_���U��um����cB|c�8��?�|�/Y
���Y��e^�}�oV8v����ຨ��~>�RYe%�RYbL�b���ﻷ6#P�֌�{_T`N�C���׽��[�@��C�$\rD�1g9Y�'i�B�����Y�>�.��C��'���1?|�Eڦ�n^��F݆j���D0a���t��"����^$��}W> �]�Jd��]*���R�����AFo�3=饼�I*v��>�b yP��o8��;�O�e�0\�Xd3�-�i1-��?G ��9�W[����Tz�)�`�ϖ�_'9�,�U�L�LG]ǉb��\n4�S *w��M��C�K�	.":�Dk��Q��KՍ���ڦ���t�y�^�� ���]K"L��9y��zg����N��lN��l���I[H�X B�%
G�긦2���@}��6�>>�;ij��nz�e���v��^8E7uM01}B��{�k��o�o�nEw��N
�l��]J�24��Rciͺ6��+\uE�����L뒰^3���x<m����>�İ��Y�>����z�����
�P��<�y�x�h��oy4���<Jn�e���u�e�#,ic$���ޜ�LF�	�X��)u]�mJ�76Xf���r5z�s,�b�E褺rc�����۫k5�1[V-�\g`@�-�����֠�eL�3v�Pn��0������l�tv�\�c��Rl�M*��Z�,�0��X��[m�f����7b�D*bٲ�x�I��JW֍Oeq]�٨�,���\5GX�Xg6X�D�ugF�J�����s�v2��_l"O3��] �	io*�]��Ӵ40hgj��K�]3�1��2��\��u�����,���̱jb�Z.oc���ff�ţ�[X��o9 �=�wm�'�ѥ7�W��2ppf��@f]��"#
=T����"I u^��cD�U����	��0��;wG'c<�˒��f?1���ԏp��j�x�Ƴ4�KK� (�]� dő"�DE�Za"����8'���shĹ��MD��%�l���L%���s4ݬ�/��4�����!L@�NVL���- E��ǯv��j�����>ٙ\\[��;�����Sifx	�UY]tT3Z��?}���l*�%\�z8K��#[1�$s;�� -���m�Ψ���s֩��?�7)D��+��q����׾UG=^`w���_}�����U���g�v�s�A�b��}�o.���]���>{��X��y�^�,K�.�~�RN����?��ld�8b��%�4������}��W�2�y�oG����}��u� -���a5@�}�ؓM7r�꯿y��~?O���� 9�U���0o�8j�BAvp��yjd�X���.g��C�7��@�aCČf¹C�h��"���1�F/
��	X�(B�ޙ?m�}��}��(��]���<�I��&���Re�RJ��2��1N�����`�s�?�c\oeG���ƙ��mW��� �����>8����4�8r]�˻���G���+�t �Q�N^2Bf+��fee��l����|����%����	,�װ�����C[_�઎ݿmk34���@a$���T��Y�g��

I8J�����y z���sc3�d���k�� H榆9$���=�Z��c3tl�h ��=�D%O� 8�X�7�I2��2��7�j�e�p~��6p����Z1uYg*��wY�Cr�=p0�F�UA�,��gL�r���g"���e^EqDp�}��~/�<���ߕ���gѾbI����.��V_��a�~|��e�϶����I-�HE��";���7J���d�lw���mc��<DVg4B��#� �Jgzl��"�|�R=��Xc�)irH�5�`$� �钖�3|�}�J@�-��mRg����*�olU�ؘm�a#�R�2��QC0��E�gʇ�>c�j)�[W��\��"<Ŝ���,>�[Ya���,7r1�kh���ȇ��.C��;�]��K��J��N��#�M�54�2��ڛ���|A�T��" |u�Qx�X ]pa Ex�MM�$�%
E��?J�d���s	����X�Pf�Bĵ^&3�mn�:I&���"0RO~c汍��0!��=�ػ;�P���	.ǻ�p��|�P���%{_���c��弝޳��Ve',㵸���4E�M�����:z���F���<��u,���x���:��X�FX�2���_:�M�8��%��5�FRnP�_�� �;��mM��I��,$�>^���YÐn9.5N!��=�%Ӽ<;�w���'e	�󀡴hJ6&���n- ��i�n�cma������!CǼ�P@8���'��z��WC�a]��ưd�Z�A	������j���ꨮ�d�(e]�q6 �	��;���L�@ ��
��̗]S���m��&.��kI%M�8��L%����/T���������� R�����k:�� �@�gLf���D�ACU�����N�"��7�ٻ��eR���nB	���@��堸� L�1=铭ݏY	)'�1a�����;�� kw�ʛ<Z�1p@L���H$c�{@�� ���Kc�^��u�T>_�:ڙ��̱y�o�[�r���b�3���ś��}�����bgnUm<�md~W׸w���Pv��E��)0K�	nTO

"��B��w�y��ˢ���[煪L��:�˽����W�v��ߝ��q��'u��|��l҄����s���^��,"��͍�a�fH���.2����U�c�����6��kD�0�U��:h��O$RR�'�����Ti��ا"�{kn�B��T�0X��U��*�.^W�6�6t�q-vЩ�k�^+b�f!���3F^��A�YO�v�}�f�p9�6����Է:2��U�ѫ(�HM��}���k��mb�so���G��-� 	�A�I1��b�5��X6NZa%�޻$D�$��,B�����	�/y�_�2��i��"���A��ù7�ީR7Q$=��`ń�W-o5nЃ����L]�����̌�xB�L'	&��� ��Z�w6�J8w��[��~��P���@v�����5gs=(" �;�ږ2��Go�,SO���lw�v��o$�'JEX<�$;M�O�T׏u�$0�ᜰ�� hdފc��Ra����I� �8�tr�4�Խ����=|19t%����u��>�F[�9f��i��Yt��x�mnV�R�yMj��__~_�v�`��|T�	؀�ߺ&�&q{����^��q�U/M�G�����+y���- �K�oho�M��~�/~��i�c��|^m��a��tG�;�M�e��o��ʪ�hf��q�o�j��s}��ݑ��x�%%�Y������z�w�t8�+��]���w Hu��M�	|����W�\YȮ,�����z��������A��Y{o�y��LK�l��z��m��,��<<�
*��� ^�!,	��n/(M�`��cS{Ke�����}����]ܻ��:!�<"���;�g�V�W��`���#|<�'�Љ�}�$�w�������{��d4�m�q��ÈJ���.�Y�K8z�2���.y�_�hl��Y��ِ	$�� ���{�bS�������֗�N��{KE�	���j��6Z,*��j�\#V��DK2����	�����4��ź�)�{b3z)��z�7�߻ͬ^�	�~d����߁����o6�!�X�g�x��X�@8�3�˸��`ݙ$�d�u�R	b;zb�}����:C;���4�M��}��&���o���ĝ���9�ꛚ�6u1Uz�+a��G�
��bl^��W�*[Vvһ��yt��Rֹܗ��sFU�ѤGa�4���꜍#,�#2e0�ɅA��`���b�mη��?�L�>gn�`�Xu��u]}B�gu��X6s�V1a�'7�"{�E�޷?��"�>�^${�5�1i�B*"�w@m��@vF]v��F�����@w�������d-b�Ո[W��ކZ8;���N7�x�Շ�ZlY���Dl�4/��[l�a���APM����%�%����x��K�$A';�,yp/�$ <��3,S5� *V��^�3�IC��cn�B����~͘�-�u� H��LҊ�h� 0w~� �;}j�eM`2j�B�$��z��H�I=U���̀�'�����vsr�=�߿����d�k����=-b*����-���'�״:#""!H��۞�[������ƽ��D�h��ZƁ��}���|^GENL.�#�eaܘ�ƍ�[�-dTN��:�sX�r�ۚ��jb���*gu�D��cuK�e�o?d��קN�]t�����9L%�0
�
H�*b� C��,}���L������,=}��� ��y���vߍ ɍ�^��"u�
�3�"����vq����y�!�V�(���c���E0��x�&@�jE���ͭ��G]r��ʲ��>�����d�z��}>�A�r�] v6y���L_g�G���ܦA�M,1�uK<ߜs�������� ���0b��b������.��zg�!���X���`5�)�i���Y��BQ�Xr*)�Ŝ��C��>]�7�TCxv��a �g�Ft-c>g��΄�@��zې�$T,�y\%���������8gr�ӬKx?4�4��T���u��D4`��
��1�VH;>�"!W������J��v�y��M0j߹	i�hp%�Z�z��}�ƀ`��+7�e�z=z��<zb�Ǧ�*���fes��+2��6c5�B�M�+5�{�Үq�G<����q��ڮ�B�ԙOv�k�N[���n�(��vSY����2c�Y]�9m=�7T6m��=��3�����sTΫ۫�9n�N�t�=�s�����V�t,Wt�j���2�>k�&l�dS/����D�H�wP�Q��ö]�7O�*o^�(ݣU-��{ˌUt�(k�gn��łi��T�VFP��+;u��)"�Q����E��M�*��v%r<Z�p[�w��ՓG =37pu�Us17l謥R�Y�|�ZS�r�ɻ�j��WV��5��t��nn��ky[�̵S�:řx6����Y�7N��uJ�5YV��7q�lA���f���O��������)<t�\T�½�*f:Ǡ�R�o�gB�����������o��W��Zlh}��LKj����yl��ےhO�g�pqC�*"�fVR�ֺ�em�ey�yv�n,Y._�]<�2ՖoWڞ���y��a�͟%g�C��޷zC�fU4�U:�1�K��ã �CBQ�h�/�(�#o�}M{�� �c�#WC�-5���*�]�
��>��R4ً�`h(�P��lF�$(F�T%Y>�!�2!6ݷr�9����E�36��,)m���H�V7j���CQ�� hW�&��I��SH��n�6��!�[�#Бn�s1�B�9up��LM�Oy�J=;��<�ïv0�lY��GN�z�7�M`7P�Fz�q�@�v�f,�3�����k�9�Uw�<���=}/���@�7�K}b�}p��~0ƽ�n�+A�E�n��ǉ�;O�7��Rb{�=�v�T�%��]	�
������C
�f�L�B3#hR$��Vи��
��Y�۫���b/�q*��P�,G����_�>��Aw�xE������}2_^֬�ݶ�x�[��BH���X��8���wLY�����{����k�r\�Ye��D��@�,�i�[(�K�9kV�=������w,��Ǐ�_�_U�����k^65��̛ƶ[\'
G/�b�U-�Һ�,mmѕZՊі�q�s�om}k��<x�}x���������Z��ֵ��z��Y�圮^y �9B��-��LT�rk�t`�Җ���A3���ۏ�������Ǐ5������������65�k����l�r|�,ͮfU�b��T�U��V�,Ɍ��2��N�s���u;x�Ǐ>����q����������}{=�̜�[Q��%G",��-��ezj�J�b#l<qS-`�Y��Hv����+-���*�֥*���r��WƵ�q0bcDL��eG�d����� �.҇��=r8��f-eڪ��6C)�,I[U�"�`�ɔ�DE�ƺ�b(,G��
%j��g�Nmrٍ�Y�T�����[fy�3oMr)˘V/^-����:ߩ�B���:�X�S2�񘊪)\����b���3��M���J�b`�M�M6���������W�hڒ�([��B(i�*��tI����H�ny�0��V����B���a�lAs�����P�P���bRa��6�Һ¶�5c�`�� v��F��
���c71Օf��Y\�S���fW��%KK
:1�e,�W�`qev�@.�����6�P&���d�0�E��r�,�C��&��vWU��#Ri��Z)p�;��Q��]��V�(%e�C���Kc���U��
B�u7e3JWjб	j�la2;m%wi���6�h�]GW-�5"�X��Q�a��"%����fd��S5���Kbbku�X��al`���ŭ4-F60�в�m�l2��h�)u��l�$�7A��ڈ���u���L9��@�t���e�b�Th��a2�if��]��V�lk��X�nj^o:n�"L,W�m�A��j����he�����Xu����+��a��L[�!t��0��I����lݑ��5v�ܫu��+���VZ��f��e�X��^��V=����BⱢ�f �6f#����aH�2e���t�[���W4tc���s���$���{.EK@��5%�(�pd����@e^�Cve\�8�%&{-,T%^ԖZ��	R4�F
K�(��L�aY�閛M�m���*��Ak3��H�X�R��]��t�J�-�.�aZ��Uƹ���-�via"F ��ۃ`��l ���[m&��0��� l:&2��cb��Yi�Ҹ��0'w�޼w�i��뽱m�u�u����ö��$;�����]����w2�u�Y��1Aݪ�0�e�Ȅ�\��y��l+�4��̆a]�U�[sZ����s5rZK�9�:6�.nF�����+2fV�]B�
,X��b;.�0�ʶd�i���s�693���7*M5�����Kɣ33l��3F^�+R��_�|y�x���}��z�avCy4K�WC X�&ڰHM�fXl�SQi2�������È���x���V�a	�����}T�Ğ��=1~PDqL��$8��������x�b"��tkK8�v<�H4���NK@�$�v�|T�	=|���ĳ�fE�wM��@��mӏɫD���٭��*�����B w���N�f���5O@M�����z@�54y��Z BgkP�J!�t���TK���諶��xi���bknn2��p���w�K�J���e�`�lgd�Ol����H JS����!H�Ow���C���O����������މk�C�L���"A���?�׏�ީߢN��<}���䜒�>��hev��s��iBR�`���45T�3-�OϿ����.��6�ۙ`O@j$�����$�;�ri{ӯ��y��Vk��S�Ic�Ԉ�L�hxqa�<cd���E�h\�S���r\�?+��=�k�&�/�Z욵�~���&��+�HA�[쇧��N�XE��'S3�a�0a��[��+,%�Ʉ�`,fL$��q]u#�H��G����g�������z�Ͷ�O����&?�lﮰ�o,�L�n�$�I3�致�!��k��R���@�I>�4;��,����h׾@C�t�����S�xs����&���h�sԽIj`�� �wbӄ��W� �PHrOoL����6��H?�T�E]�r6�t�_��t��;k?��0x��א���ґ$��L!��{w�AM�㯺�qU�����W�rs��.�̮K���mX�Yh��@u��/:�LDA#׏ܢ!4(O���|�	L�|�:��e� �Q�	 �뼷�}��X�K`šޭ,]3�Ո"��F�=xs��Gy�gW��U ���2b���mi�e��{����d^=V0h춶��t<D�
"5�Z���4Q$�۫-��� į7�HG�����w�a, 1"<��w?7]#-B�S����oR�}��Ǒ;���-K���$�O���$�u]vNԒ�%�%�u�u�;E�ԝq]u$;`��Il�Gd{�뽩����:�|w�3�?��ɔ3y�i;�x�4�������}����a��ݓ2I�~�� ��Ƈُ��`�+�"t X���#�!7`g�D/�x�I���o2-����7�Ao4�l�@��<Sx9���y�ԧU��{���؆R�{k�,R�,���B�.�"�����~�f˵�K]��U@�H;��1�"��<�F?��f�r�LKC;����̘3�{=3��ۜ��"B���֋l��s�p�z���p4�@�~��N3�� ih�cM��/�6/:�[�Q6F �ݍc�MԎ�z��!y7�n�S �|���PE54
���=� ��ź��� ��n�A�e}�� E��Eژ��A\]k৞���-窻L$gF63���0�X��p�=�Y���.�ߞ1�i��D�푥�ap��������>���rgQ�������:��*�&���޳���=TG��t��U�d�W]��"u�u�#�%��l-���%�3`���M��O���G�1�v@_�A�D��f�'�\�, 	��R'ى �C�����=c�z��F6��6��N�O��˘��4���dbDz�{M����3�nI>Iv?�G�(8��~3�L��^��7�CCyv(�]��������bYkZ�W�r	<8N�P���0��^���`�1�Y�Y�����dW�����x��X1�u�!4(O�G��o�1����h�0�;���<�I��2���\�@'��s6��;臇1
|�ݬ�LＹ��So<�bm�;��gw��N�$�0d�3�:a5�p\�{�@�	DD���[0��9q�s�D����h y��:���U�@�@"{zd�h�=o,�JS���=��6E���*��:�dU�*5�w��}�������HJ�n(E��k/DL�2��	,��Hl	�����a[p*M<y�}����҉���s��I�~�����!���$�u]vN��:��1!
I�{���MS]��[��BS)�ķLR���E�����c�pV��%i�J�t�iY��hj��N�0�.��ZSD�f�V	�`�,�؎�q2R����GBm�i�Hh�YN��&Q͚4�t	k��Pmی�(�,]��.�]7lC��x��[�&�X:�-lskRx'����+�?$�z�Ai�dK�ن��tf5���s��ak6�G*WϿ~����1Pb@���#�๺�H����Ҥ��gMu0nZ�<���#X�jX�A�$��z�x���gh�,��7��t�+u��NtH,ݠ�bw7��@���U�a~�u�<.	3��75��'J�y�'{1I4�9[��yd� �W�zA�=��$R��9	�Ӭ��H�&�	���ت{�F�~����� �꼟7��`wK�Wx�k�?O��`�π�&t��C����/a��<9�Wb�jXH�{��&Q�����C� ��l���3d� s8��һƳb���N#�{лfb#�$�{�&-�ҀSX�%�K�l[`s.�y�\T�&�'��e�O��o����~B$���˽RH �Z\�{�?C�y�LPb���y���0�$��芈P`�1Z��H��7���Di����0C�����H�Xr���Z4O��Tߥ>�r���0�Nu����"8�>�i+<�[H�[jC��=�3����=T���}vBN:��$'W]�GjI:��v�Z�Ж�I-BZIl�h�9�l�����V���w��x�C;y��~�Nǘ�� �x���M]hO7� �M�V��.�h���	�Ք�H��$�8�&���P�4 X�B�[��ֈbHۍ2D5��0�$��:UFjR�W'ۨ��,���=��]�<1W�i6��srt2�}��\�π ����~��{!ny�{��k1�������`�@����w'w!��p�}�-���|7ث3lT�w�'~|=�����#�I�`�#.h��#��EZBhŨE�ނ�!��B����ɳ-{���Z��;c�!m���ũ�5���$y�zFHH�@-x�j�x��R����@T��z��ف� ���1�sT,��'��1A ��|��"�e]�h9���*H�݌���Ѱ-������������+�ٸ"��?��6�g��(��?|jT�ߑ�ڨ��[��//(+ǝ�f��.W,F�+�ѵ�u�o}O�,I�⾻"vĶ	��R�Ԗ���hKD�q]t;BZD�l�-�-�$����o+���zb1��BI-𻀁�$�{x�xO-N��-��6��36��gp���,@{w�g��6�����F����7vŮ���Ä�M� �##�魔�J� X����Nu5[h,h*%,M����8��.�˝>���g�)�m���ck�aZ�]�$�,��n��Qѓ-��i��.����U�Ը�SZ�z{��H�&�	����&��Nd��2/}sc@���Ԓ}p ܂�oA{��!_J�0[?�Pu���F0i�d�Dy�{�yܡ~��g���1�#+*Y�_����Ɇ{�te�����=cL�?�kwIx��$�ن-C�3�c'��ї��r����$mh����9ݒ7�{ۏQ/
<����{|����$�;���gg�z+;k�1���Ǜܞ���n�Pt�[�n�;�����l���Fq���=��e�Z�;��M�{�<��޴��_��兿�?��͝�v�����;b-�����	;,�E�$�Il���o��Z��'V��.'��S �gp1��i%�z�'2y��k�����6�����o(@�4:�O����?ԜC�&���hֳ1]P��aCM��2m����� BPvdxt�:R7���D� �5y#ă���e72gTWHj���UQ���g~u���W�{��{k��$bB���s8�6��D{��[N1�W\x	,m�3g�S8K�KC2���F�Z�oD�c�����CØ��L.�3 �3���Iܪ�zw��hކ	�$w�����$�{��'�a�q}�^#II<F�롯�Ը�O-` ��D]�T����s`M��2Q|�~ʕ�T��]|�
�^Vx�씒����C�PbAl`z8"	 g�B�3�������EҒ�44 A��`��� B���.�A��_t<gR���v�ED�*P�,�d��4�T,�4�1
��E�Z�U���2��ç�T��\4�X���ili�S�
$T~YR
�J���a�|�P�ۦ1�r�^*^V[�vz.Ԗ�	P���"=�����=X�d~��t�ڎ����v��u�u�'W]��"[$����ֿfNKa�s�u��±i�Թ��G%ԂXR��(�3YS�:i���͚�b\"��cK�b���lJ��1�LGB�ՀkZ[��a�Z`rJ�h���n���.�s�K��2�����m!�(E�&��+.]pͶV��i����Rj��p�<����E�%��DV&��]D�6ـ�$e�c7��7� ��?|�$�,Xu�&vw��@��ژ�A�s�RW+�$K���[�;���/��>c�Q����� X '��[�{���+�X�j	�e� H�sDC� ����}�����`H v{7Z�ދO�#�U$x�@p�]ɭ�Qy������:s�444yt24��Є3�o ���C6���1
|L63fZ���r
m�j� ���Z@,�� ����8��.���=]]�ZA>� �m����%$��b6c� )��$=$�Md���4����ȑ�� [x<�����I�<'|xN��&Yn�l�Ͼ����ф�,[�fL���E��b��&EvI�N�S�7�D��BE���~��C��~�0��ozI�m]E�"�vn��B�!�9ÇI���GT�`�v�n�}u>\S���S��b`�vF=u6s�t[�VșWD������g����e�g~#����[E�/w �,
 -��@:I?��u2�u�GW]$q�u�"Gi���߹A"wSKC��{�3�F[�H^��~�U _�v=-��I�J�Q$���=>bvw�s��׽������oon�$�g�жm���'�:q��1���	�AU�h�{u6��2lh� Oz@X���%�#����\=�3�kD�v�gA{��!HMv"&�	�oM� r�7���H���՜��;��H�&�7^!T"�`hҤYV!�����D���	\V		rY�WSEu�AIǷ�"8���u�z��AL��f�z��3�'s��f�}�;]f��@�d��1I!�ּ͑����A�)�$^���L��U����㩌c�Hٙ��l\�E�� y1n��7�U��c���Sv��ke=�cPr�P�c"�1�.�'!$�g�|盟}��������+N��e��om�K)(+�7���t��_?�<~f�x���By]{b��,�w:��!�Q�yi�VuNv���h�Vr��P2úR�J4Q͖��RfG
����E[:P�:�2�e�.n{�������B�s�n2vm����[u�ΡT�n��̺=TŮW�>���u-�T��g7��Or�<�Z/r�DS�b���E:�ϻA�7�^���na��X*Μ[q��zW�yjM��G�q�[bik7Cj�u��n٧�I޺{�����1eym[���u�M���R��2ev��.G��ƁE��]o:W����Y�+��V���T�8hy�
��z�B
q���{y�yu�����T|���;�XUR��Z�[�㼗&VF����s���쮫�WM��j��+Ŗ�d�!0e��e^�Ԋ����N'-J�x��5��\r��՗�nd75;�uޛݳ��ⳙ���Vne��u�[}s.Tu�����ݥ6��tSx��L��=eEsh��ʫy��up�o	����Y�F)�A!tr���S�';�(�ۺ�7u�]�1�7x5��A���(��`Ң�s5�k]��Vƅ8��xD���a��Y��[���^��HK����Yl#e��G�
�uN��8��1��hbb���j���n'8��* �Nբ#�Y��g��s2�)ӮVW�D�o�}�	��}/��2�ᯞ��J�Nm"�Ɠ��
��gͦ<aW��彳�?M/ L�3\دۛ�^c���%�
�\е�_=��M�;�|�ZI qܒ�H]�ܩF�`�hد�EpV�V���fQ����}=���x�Ǐ5��k�k_____^>����}2k��'C�����p�f6P��=��'BBЍU�x�o9.s��N����:��Ǐ��mk\kZֵ����}}}}u����������27zSBX$-�@�9��G���A-髌K)��I��s�������_<cǏ��ֵ���kZ���}}}}u�r���2��S��x�qܢ�1k+�#i�X73�q«mq��}=���sǌx�����Zֵֺ�k�Z�}>�NNs���j�QƉ�o�p���:�S��Zз������$�>�b��E�Z�S74�8��JԵ7��f�s�T�����G�ZZ�@����m�Zԣ��9�0N$�s�Tph��f$�,u��XT]J)�s(S-E���8�Z�9�6�Q��U��$m�3��!X��h�y$�Lh��0SX�UˏyJ�ShWmc��Q�wM͚���!S�x	���]�˔��(�h*"��0W)}�gl���b[rѷ��-��d"&%��a�W0�&Z(���Q\*�;�g�������H~��ۤ�:������:���퀱I$�"�c�����__���{�v�44a��"���mƘ�Q
J��H�[���8�'�yH�;����b@���=��8�x�6���YEڹ�@��>�׽Q�~�!���.�z7ձ'*�w7~�a �s�2� �C� 䵌�3��~�p�B%������|3�4�2��k3�KL�)(��J%�N�-M�`()9�_�gA}��![uzR�qwg��"	&}ɋ)����="�����Z	9�p�`��E���l@�2����e��^ �} F#���H"p�����=�|�z�$;�rV��:!�w�0y�+�6�1ǄY؇�;���]��s��E�[��0X)l���M��
ECt?ݵ% ��,�|�<�,gr	���i�q�V�V�W�v9 ���[���#}�(��nJ"+�æ,�k���n,9�}1��N���*���d|�5�t�Ak�D|P�������&K?RI?^��$�u]u$��$�밓����I�B���IS�g����s����73s0)*Egp	{���;��[�ēv@>�֛c�_�H��q��#��|�R�s�~�OJ-V����L32�
]�-�tB:�s�����$���#b4(+���uʶw �T @�_;�d�Z��Խ*�E��G62ha�^��"�jE��b��*@-�X�O��:|�奋�=X�.ϐ�E�qi�nZ;ޒ$��Q) e�e�<DXN�(����r�8p��7�W��rDUN���H7�g1��L-3�;[ʛ���cL��6!�w����_��&���0 �5��'�p%���]��v���.�LB.�����W頔ɭ�7�Y �JU^�@��L�Aj�jC�h�OwE1c�m�=?L١ur��m�#N|b���n/י������%c��"��t�f�_Ҳ�j���j�c�Ά��>Dq	���$L1�	�>�B��EՅ�K �R�#e\z�_�K�F���X@ �m�y�Y�DQ�	��^�Dq�\v!]u�d�]u�I$�H��"�${�}�_s9{i~Рi�;h;q�5V,1�9�%���ħ#-p�Uc5�D��p�f���m���TDRWh�CBf9�L�f��6��!��Ή�n�z��%hr��]Kb+Fڷd��g�l��溚�)��[�Q��F�f��K	�fi�[T/�:��T���e.�+�
��ͥ��U�7�&P�л%3�T@PA�}�|K�^��S}�=9ŧ;U� ��A�w{]�4��.s75�	#@�z��<�w����NM�F�:hPU�:�a��r��P ��v����4�=�m"m���.~z����cRi��V��-��^}�(��~`o��ͫ���Ko+
Y�@p,�y�9=� ƌ����GC�ϗ�t��D��(?'����K�h��\��q8|�c[jd��S2@#Z,�C�Iކ�`V�c�	�ʈ�^�_1k%�jq����Y� ^K�g�A3��ܟ.+�;�b�m]f�]�ш<��E�Y�{H�#��E���(Q��3��18!�?r�G��)�MfE�G���scB.���Na�^��Þ��L���w��\��0���`z'�&<��������
��*�{�l<=>0��:��چKǛ�c6�k��\v��5���BA�yZ��X���xa!+ �XHq8�� E$��ʇ��؇돮:Gh㎸��8�:�u��%�؂�	XE�HFH)~��o�0���o��}.��,@�D�=�M��� :�������PD(+�<u ����@���A�w��|�B�	|���~�AC>x�k�6
��I�����������_�Ӽґ�m�=�5!�QxZ1 #aХ��l �s%+,iE�Zuji�����5�Q�q�֥�n	��ky��[V$c 	|�0�+�C��������19@�@�Oh[��(�w�|ͯuN?��d�0'��+gkm�-�q)$t7A{��	�{������љ��ߍ�o� ;6�w2$�]<��L�.؇مq�;�1�t���v�,:Sk�2:�+��͆Z�ktr�}��>|���O t3��dZ��˄�[�{&@7��.����|�s)7�Ks<1w�2��ܻ���������}s$�8	�m�����*�цw�ﺘy����)��[͹��
�i 㘂I=޷�����3���,M�v�!���WG3�ء�56.!�+��3F`b�Q�:����Kw��+����X���Ҡ�Z�9��^o6[gl�O�\tJ�:$���W]q�"v�%�%�-"+����p+v�;��/�
e}�Qq
�W�X���w��M������G�Y��?w)�,�6�2��)�.H����_�"���w��	����ч�6l�-��Lhg��V�Oʇ��M�L�/�g�^����B��`B�`	���ѹ8i��G�#���,f��p^Pk�9������l't���g�X�7תGJr�� A���Md����z�n�KHrIk��$�h�ypH�J#���^��b�7\�t(Y
��F]1%3�V�,�o�8���{w��|G<���ʬP`�
!U��x�NxO�Pwޙ���SD	ga��3M��C�^ቅ=�4�Al��'C8�����:Ibw/��*��@�y��p���,�Z2�"������Q��<�^��9{�U��Ow�t��Ѡ^a�6�fU��f�F:<xj۬O?�oA���y(,��d�%C���'믎;+�������'u�bH��I����7$�u�;c]�f��
�|��A���@�G�#o�����g�����K@�	�Ę��#�=�f�o��0��~a���� ���l��)ZJ-��˚&�AX�
��ъm���輂�"!�!y����ۙ,5[I��� v�t�jI%d�{��2�w�$����:IE�M�I�cU�̉H\Vy�WE�jg��%����|Y��.���.�:��DƝ�/d���$U.H�m��Ŝv{�4��E��o-)b�w��������"�$<'��滞ʜ�6/�ֽ��`��^l����{%��8�S���7q��kgtZ~�埬��Hm}���1��x�z�Q ��l��#�v�H�k�����!��=jA,�����@���W�.�W{��U�NO������C�����.����+�ݫ��yV�n�4�y]�������#�+�۵_Z�q0��\U�/
�]Wʞ[�y�Zl�S�+�>���E,'�'t�����ac,�f c YfK3@�̖d!���+Hru��}�m���㫰:l�Y�k��XA�62�
�`"L�3�W[�ka�1
Rm�^r�c5����2[0�ئKZ�m���1�ny
T���õ�F�AcQ[wW4�5�5@f�4�.��P7g;lXKH����d֚U[H�Ԡ�V�:֏���cz��J����C��XA4%�����Vl��7��A���	us\{��c�S�54����y�5�y���td�?\C��47�爌���w�f@$^�73����m�T�g&�Ա�y�9���vuY3��ҳZ��$����}jI��?/@���=G��|q�}���îS�& �{kX��'��s$�zh��| �(����b��8�<��_ScF��8�滦q�hgv�g��[��ު}N�(���~���ޅn<GHxO#21T��h$���3'g���@5{h	$ ��Ҏ���<;�~�P�UA�q���l�I��!Մm��h���*�i��N���1p��P�����ߟ(���_�����=up|��#�ܥ��w 8��^��}O=�J�Mj% �Y܁}r����C�3F��d�T�#z���n�e�+�:�t�4��/E�Au���4/~z*��8�ُ�׃vY�>�H7Nn|س�����놽�7���Hv�%�K0$�8�:�]u�d+���N9'�Ȇ?1���:��?5;�%l\�Cӎ���ɯ}�aD;�)�R��|gg�!gء�������#��d���G|I;}oj:IF�x�\ud�~�=lŵ��`B��!�"i��7Z@�>&+���ˏ%ؒ�q�m���YҬ�aA��e%�ۻ+���������`��K���I��v�VtL7�3��l]��@��9����OF���C���5M�4�fs@��$��Vܚ0�,JYK]��K�al5����{���"�����'�]�y��3�C���kK<��w#7���92�h6�?b��e�')C��$��EE4������إ;�H$grL@,e��A�N��v�⮼���@x	;���"H5T)���b���~�b�#��;3TI������v�Wp�N�W';l�;�-y��u����*����+'W�uf�yǤ��Eb?�kE�JDD|�@ |���� j�;	]u�d�W]q�$��I$΋��ۉ��8}��.�\<E��!z�{�2�u����g�>����;U��HF�s��r��2|j�!��֛��RH��=�~��X[zY���{���� ���E7��I�ӎ=�z4�#�/d=���n�bԆB<�&�.�mMF��3mRҴ�-�KV������,�;if�8i ���`jS;�8p���:ֽQ��x���v@X6^��v���|�y�6>���tOմ�A!��ݚ�$gs�q�dy��WD�����"g���WH@����N�FU@�T"Ij�0��I�7�z���l̎̆(Z��"��c>�I��|I��r��iVM��~M¼�X�&:�.[כ�<I�w�U�=OҾ ��=��ѫV��2V�D8h̬��(�sBQW	����V�:�1�:]_\���\��8��TU%`noCs�Hx��?\k��W]qԊ�;Q]t��/�@���	��;�����L`I;�+�^�D����2�U��S^yb��^�nD�wc���Y]���F�JĖ�c#��K��sq��л@��
v���*��5U��[J�u�[}���w��\����l
c`v�����䏪���?,3���IH6ח��$o���]�a݂�In6����O��ϜK�ǟ|�cwM]�\[K�L�֎��dވgw���.<|��Ko:F_�
��ɱ�"���Y.�%ؓٲ$����F��� ቍ�}��$܃���o�Ju�0��Ya��Ȋ�᯶�<�B����LX_`��;}�ݦ�����6Ϝ1��i;�NPV,T�L�8�^��̣5��4��HΚ��S'Y۟�#�0`�~��ab�5�.�9��������	N�:�oMܕ�����R���s�:o,���v{�-n����ˇs)'��V�#҆��S�J�F��j�RP���z=�*��s"hØl�u�O90N�zby)w���0li7*�0�A8&��k:��ެ+*����v:�4L�{o�n�f����c���^2�,l��O��g�A{꧄�ʘ�<�s(;�͹����N�3�^�U[մN=��b;��]�<�2o^km>��xu]���Sm�U�t�����J雋[83�w�c@�����6���eP[�7��]u�:-��)@���!��/Ṷ�'9n�Lr��r��ߏM{\�rĵ;�e��0E��v�JyU��h���O	�9�s��ʡ��DY���xͼ�D�oM����w(��o��9�7&.��V��/.�.��E^i7�J��u+��p�
��/7}>�k�@����,Nn�y�eK���xc�=���j����nэ��3la;Ll��;��6
[����K��Jdj�ZU��l�h��wӣ��}�)J��Vd�L���
$	$����{�ʻ,O�q��}�Y<�bՓ�^�����I�2�)�I$�-뾯P�Y
���h\ʩ�ːk0�sҏ�h�Jn��lF^y��KNˁ��@�p4�^�o)0�[B��ULDI*7GK��z����{�����3-��7y�mz"����"���#*9��B�U��m�`��.��Րǆ$�uuUN�w�t��A ʢ�+�AUIs�#�*�-sT��$m�As6�OW�zVm͗&ҩ4ƗLa�8n]�;ͤ�z�>oO{Y�e
ͥ2Ԕ#X.& ?}	}��{�9�nO`����3J͍�����.!	[6����f�������kO^\�dB�%0����ݤ�ْ������4I�����j{�gi�+=/���\zl�+x��XE���ƥ^S�8��Z��X�Qr���\�U��Et�l�g9��?>><xǏ5��k]kZֵ�V���Oie�ݳ�;~Ynr��6�
("�˓�^���R�_d�(�Hu�-��=�O������<x����k]kZֵ�W����rpz*=Z�X�ӭ�A�����ǦÔ�޳�5�m.6��J��2�F��f�n����{><x���Ǎ}cZֵֺ�k�Zg�������fʭcJ-�Vmq���*Ԫ���ƔZZ�ڧiFaJU�Z�����}6y;�O'��<}}cZֵ�kZצ�Z׳g8�Z9V�RѢT�r�Q�,hѬ��"`�gY��ƭu��A�im�kK����L���+ݺ㋔F
��n�Rҕ(�km+*QDFXT��n����T)iF���E'��f�L,�\��%�,��V,�J�Į!�9m�ckj�Z��f5�*ҥ*�q�&%e+C[�[�v.�[�Ȧ2�!����AU�6�e����ۘZдh���EX��Ե���6��2��q{���8yj��S���(��*�
(�V��-�&8e.e�uySt���j�r�0�^�W]5΀�ѥM��*ƅ��I������X�e�nb"�\�ltlteWIO��᧭Z[�W�!
i�9d�rJVk��a��d��(Me�R��3+��6h�4\�	3�l��T�.	u��Q6e�ԈSM�+x�M�ֺ�a�����ƺ;
h��j:Q�e��kY���!`��-C �-�0[��,�5]J�Ŷ��]�e��"��,���(����٥FV�!e�2ݔ�E.��L���!�.Ե�˴�%GX5����̬,�Ůں,%�s��Z��14���jP�T���%r���i+�64[��6���Ȭ��L$��h�(�#4#�`G����tثy�1h�Z����M��̛)����N�V�nk
@�Kfp���5�Vj�������mhF�܋�jlR˘��f"��*���],q���xٷ�}@���Jn�1��[`��R��
H.��jb�
M�.i6(���A�-�IA˓7����m#�uGQV�[�+XJF�ۥKn�\�R$���җ[�`��h.�ѱ6���LC9�V����i��6"l��tˍ�tʖj��k0���8s��H�F��e����%Ś��3A����pj�eK@ �f4�0R�X�vP���]s،�q3�S^�`c9f�eĶ)-ƌ��Fj�A�]4��m���#Ia��Gi����`�6.��)HƎ��%��R��f�x���k]X�5Q�\R�c�^��K8��Uk�1t�n��6mSG�ҵ%���A�F�elMn�m�KO�ӧ�߼��toHq��W]qӵq��jI:�!7���꒖��+�uW)�$F9�l�a��/\R�l@ekɴU�,d�D�Ԏ�����^��k�bQceθ��7mVLs6�2�(��EB44CJ VD[/mz�]X�6;Y���eZ8�b��f׌���U�:�@��2�%˥an�Eқ[�)3���r��b��լ)ƙ0K��b�lՙ�s�O���~��w�R%�&�~1�� ���.���*�p<@�WCeBG�!�ʘ�D��}���;�{�9�$T%���i ��o/G�7��H�wg�X�A ���C���3.�wv�z!ô�>��d�'��9��F�gyˀ�ǧo���w����PɊb�w&M����w�W�>NC�xl>�g��[yJ�q- }�!��,��Z�3��()��{=��8695�B�{���Q	#	*�@��������,���'�iĲ�%��9�"D3���3���#�ِcgI�xx��!<p�٫�����kt\Sb\3]��f5�WT�@B�^t����9Aw� l�4ɦw6;a&w �^�wYÐ��^5��̀9����[[4���
I�!x��A ���nC��
���^�x/y=V��a��eb[Sj򰮹0��09/k1�;��VQP���,�1��H�x�q�+����\t��\�@�b��eU�ǒ����������/�gpTb��A��zʲbx�����EBQ>��.�e	 �ٻ���.��M��S�˹��V��4�4�`���@W��I�~��,�^_SI$�9snp��Ɔx�M��z!M�$����;��ɐ@$��y�����#X�U:`��
�M��"�V���k��<�w��s�3��U���8� ��|g�ṽL�+�i�����zg }~#N����%��\��0J��mb�h�\�.J��o(Yl.�.� $\���)�BH�K���P�"��u�c�;��'�I��]��lxV�	^nc��SS@��}>b�����W{_wp���keE�D��w���	=��,�� ����*��a����I�7P�$�	]>���I)��w��;��"�j�~u�1���e��L3zi��]�����Y��2bi�Ws�ũ�uW�f�]�Rڒ��'��D Q�6�ğ��8��D㎸�J�:��C;C`/y0�L����^!��_S =׭���$������>�PD�@zg=�@Iy���2�X�@�]of�
-߽ȍ�?.mL�۠4_�����[�Θ��K3�^W}E��:ua&���&������k��~5=Ub����DՁ,SM5lKd��k�]���Pev��>�?D����3�]���$��� GlދKƦ�E�H����tkK+���"xIHML1TY��{�������%>�o6�I������#��2Fz�x]�3m�����L(T�"��53��3��ҹxɎֺ$����RvL�H���i����=f�s�JI���h�[4�6<��fް[xz;r|��q��%�1{m��p�cO��dm��s�*My��nr�g�ߌFn3t��+>`�	����a��Un�t�yI)�l�+Э��z���7��L�  [���I]u�I�'u�I"�~���� y7ۏQJEBQL�`vw$�ݩ�>��i�b��ޝo
�P�K��N����4�{��a��l � �80�k�P��╌v�`L&l�v�4f�6�G*W��C�}�r6(���R�;�;��S�>gܦL4A�uZF<�a��di��[r�d[:k�xq�9xO��Ǻ�iX�w��n�/	nca��)|%���醗���8�Z�ݬ��ʮ�
u	<-�x>o�l������j���_-��N��E��]��7��Bgp���r�߳���r�9Ao��� D�o�/Ο�ʣ(l�;�݊c!��w�mdt�v�A&��:�bz��eӎ ��BY��H9�\��wI]�z�K[hzguژ)��9nH wtI#}y<�p69.oNV����9�]<s���+�ar��o14r���;,5�J+�F�ه�kL�uK��Nͻ�[*�uy'���{�J��ko.qY��3��wzB�>GТl�@�2�3vj"my�u1e��&��rS�w�x�G��$����0d,�%��,�fHFd�f ����{�䰴#���]s�u�66;!�u�ļ6������[qMAq K���&|c�9{I�Ɖ��d��e�e!�1Yj]��,*q�u51[�� f�Z����f��uc,l3�i*���^�In�	��ظWMGF�!��1�ؙ��Z�����30�nB�ɇ9]��v.���a�8a33&�����$�����/�  A���I2��GWSL�g���^=$���l�&$Q	e���#�Q�����$�]�uW��<��65vﱬ9c������ɣ�k��T03EfD8�.�=���E�L��.��� L���o��؄Iq�41�7�?�����붑.ŝ"+j��Q��J�M��MحQ~=���L�����ω�wlwz���~�����31ம@I ���m'.S������������ʇ�7�x��;&q}ց,A#�M��s�V��9Ő$|."�ZSBznU��V*&��h��� IYb�����d��䗚̄��7b���u6c`*�F,���)��j��R>��V�dsKCJvٴ1�� ��X�g���q�yV��^4@��]ؼ���˪��<�$T%<1��@�k^��_��kX���v���#�z��+oJ���r�^Q1\�jd������v�{y�,���c秾7Ĕ�vͥط^7������o����b|��?t��뎓��q�$���H��XOn����� ט�@--��H�H$R#*�����~����>D�(��,mͨӼ5�A,@���Y̚9����]������54� 3�5���*9�⊑P�������׀!�I�g�^R�δv�IO���n�n��\�� �H@zH=��L�9�i���[�Y�;P�w��呣� �����p����H�m;� �ٽ�㮢58�	D��m].�&ىV�嵍�΄��Q�AѬٲ8�����u'!�(.�<M�LH&�#�m [����oNr���P@K1W�"u�l㛰�'JG6���:I��/c����pvg�X�Td���w����:��3���#:I;���$T%��%�g}nn~����cJ��ai�ew	u����+��bF���Uυ��E+��;.��ۣF��y#b��<�#N�u�$]ta!b�!z޶"�t�'�z{k_��$�u��D���N�8�;$�;C;@ �ng��40q�(!O�����_M�͢5�x�	[<�gi�܁�0��Ƈ r͚o9 {���|ڟE��I	)���8����\C��r�=����C>g��ĕc��^�[���X����L�g�@�L�ݓ:vk�t���<��r��2!�Q#l2kCB�ı�W���v�+i;e�LKs߿�����#�~�Ku�@�/۫��}�\/z�Kj���(T����Rdĉ��a)?�Aw��8���sc��[��z��6w�y�� ����w�&�Y�7r�E5��[�|���w�i����5�4 &>�$\y��O�K,���0���4@ ^rdM3���~�Y�G��-��4��ÿr@_��^�(IR,^��soh�e��Я����\�0 �A>�Y,����A�ϵ���?N��Q�6�^U�u:T�@���i�+>���Ϫ�v�P�s2�Īm�v3��L�����w�ْ������N�+��,N�t������뻾��~~l�����_�h��1�A{xͧ	�g0d�w�M1�yH,-���@�sy;i�d�|k)�{n��~��� �PZj���ں�pi��)�E���؋��B�"���J�0h�t]�;N������~��2H8��gh7���I%�Y�7���^�m�Ǚ�����gg�g��ii�v�̹�$�9���� NX���U=ݷJ>$�Hk����c��� (E�x\g��[��I'��:%~�*�nl��_$F1g'����N���n\/h��wgz̆���& Zw�����Qʛ�Y�kڿ;�M��4�����B��;(���0��_z=3�����������A @��nܒ@������y N{<��{��X�E묭����]��u(Sڤ�vrם�$�4��1e�3�|�f���w�3���U�Һ�Ѭw��+*�=��]܆,�o;;��S��+L��c�F7��Y��f�:$��T���{���<jc-��v�ۼ��G���1�D�x�؍����Q�7�j�ԗ���y��Mm�ʠe�vֻ�Ě��T���s��6��ǧbr�;uؓ��]���<������ O���[��)��̣PˋZ1�U.ر$�i��j�Q®YRm����;]�mh�ܫsW-����-��5GU��S�	(FWl#����L��c��`z�Yp��LXj�t��:��d���@���Is��XCm�����H�g��}t�"����9�m��iؖS
hg�2��Dj�T�6�W���G��O�Rx����A9��3�� ��z͏8��|hhy��ޥfA2�Bi���t���h=S#�T����zІN%�����$�F�L� d�O230C�2�4���羿v�H��w�b�9$�w�@De�)c�Y���š[��]����f]&��CC��t����b"";��Br�Ѡ���.�9w�x�b�}P�,���y�2H/���il��pפ���_�a �>�އp9�k��?]�A���C��j��KE�W�C"}\�2Ȃ.����,�Q��=}��<�Cʄ\���Hl̠��m,�lE �\ˡ
��e���6�(����	BA�O#��CSp|�����a�Њd�ʲ�:Ĺu�t�1�{�(��w��?j��R��Bّ=^Ƹ\��%�.;�"I���|�Xj�yW��U�G�}�P��=7,ƞ��%7�U������J�L���nJ�]��_,��w>��ٟo�����~�?c��a����u�Q�뮤��~{�����^������Lgg��8����b�
b�U��:�Agr����x��]'����2����8FO�}l�twM,����Zͽ|��-��p���Y�:w��P������w�@�U���b�I ��C��'�8j�Y܎��%���Br��1�I;SDy�Bތo��3wz����l��3^��� �A���}�ފu����.!�1@����h�k�.���5��7�r%ʰfTm��ґ��f@A��e�r7��ӫ�|��Loz �3��x��xʚs��:�~�����ߒ �� �_7 RExK��d�|9{�_����T��3�%�m�L��0D���Cy�Lr�b��!���I��/����ZDk�6�_�I̖��߈�ulڗk�j����7v�UJ6����|���a��{2�s�zt�Ɖ���t��ʵ]�7v�)��ڸ[9p�wG���w��K��ƭm�uճ��d����v�[f�OE�/��v�VC�v�G��U3�igq�/�c����18�y�t����̝��es��
����j;��yOj�mv��|��rM���>����7*� �3ko/6��u}x��;-���0C�i��5Y��"�kdh��\�ͣF���Z�WoC��^V����k�����1zl�G�/�i���]3S��:K��V,��7iI�^�F�I��Ʒ���4*n��/^>f�����aӹ�#�whUΝ<R�n����#���wJ��\cE�fT6��!Pj�Z�ھ��Z�U��(en7����uJM�`0R�SH��/r�����B̮�);Ħ�FAt�(�r�k�u�3m,V�u��dW{�.�.����E1V�t�en�X�X�����G���-^��v�wz7�fK�]�Ӊ̱ȡ.���ɟ*fY��<(|q��N��kB���Q�)�N1��d#iX�gp��J)��r�]��x� ��B�(�y{��-��}�����X+���u�2��Q�D �|�;	�F��ʻv�����R5�S|�V���dQB�:�/�Ss��ì�|e�:k֜b�ض�|J��\|�"���)vG1<� �Ԅ$�v�UJ�Fn�K-�ȏ��Tl�{��.�I����'W��9����u>̜�c�����ŀNb_v�Q-��PUQ�J����/ֱ6�)Z*�R;\��>>=5�}{|x���Ǐ��kZֱ�kZ�ֵƵ�Rܲ���I��,Q�5bn��0]nZV�ڵ-��x��6�Z�+*%�r�����믯��<zx����kZ�5�k^�ֱָ��[9d��%�uL�-�N�Л�b(*%���V�Yq)���Z��S�j�*TD�[1��TK=�N��ٓ���x���Ǎ}cZֵ�kZצ��6{6qu��Ŋk+D\Z[�c�h�#��ŭ��dq(V����YYS-ή	��{�����<x���ƾ�ֵ�cZֵ�k�k�%g{��'%��Z�%�(�Y��{�QL�[��
���.P���f7-JΜ�/L��l�a�P�+m�h�`�-�J0��ъ�=���ТTeN�1LK*��)[ZǻEE�+l��z�*�Q`�!QCԮEQb����J�Ѡ���
�j�mE��aZ�s�t���pE����1b�T3,b�V3x���6�D<j�g�"�Z�j�6��L�����b�,Q�(�kk�`�zޚ:���I��T�UW�e��ԼK�[%�ߓ-PH��'�~1؝����X뮓��]B>�{�m� ��S S;���1<�c1� s�t����J��oB9g���b�i3 �<�䷻���2}$ [險�­�Q7�'�@�s�N8�0\�Y ��r�@t�]���w�XKۈ$�OwHƪ7�*R����H�<h�ɵ3AX�6�Ҙՙ������Xi�&��.�s�u��BN;w�r����&��G3�����*7^��Q����z而�W<(�*F���P�	6��Y+�WѷP6c���\���|�v����	&2�`n�J���؇�O��ܷ�U2�c���Eg��(t���E��]<�1���e���{�#~^��,���-.X�or��ݿDq�Rx�$�)f��m�����Ҁ��t�SB���SzX�u�޼o��u��S�ΉX����.���ve�@�[�����w��r������9Z<�G�e9e,�V&�r�[�VD��3Q��~����w2��'�{x�v:�c��t�2d�e�:�~�M�no�[j^�\�;�I�*:�H�?^H]K�9Ӎ"Z����T2��@A �M۫�խ 9vƁ�|���c��Kɟ}��S���,ҥe$��u�Ko��p�uy�����t��Τ��X�iQ&.�ݢ�??>��4nW5�x{�x���c��� ۾o$��=�뺤�[k���g�[{�n��0ְ�I�/��n�]�vE;nO�K	gxg[ޒF8	��.P�m��n�LS�V������S�@����I���xܝU��;�=3�bs@-�Ăw����`Ǚ��(��[��H�BO"��:��b�
��2v��y��RXgqV�ngr��1c=�lҧbG��Z��-�n�C)FF�f�?~����"��į��p#-3�QS,$�8}�xD��� �5W�x�8;���*����7Jf�>QL��V٬�=3P�n�Y�[�]o��]@v��v)Ռ�����k�gh=�B22�ag��Q���+
*���|�. L�Y��,���--�-�2���'��O�v������뮝���=��;��zOZ�K[�,a�hX���Ts��,ٕ�iN�#���e:�`��\ӭ�5�`v��1�����4r�vq��vfy�I[j�+�2�T�$&%�ī�6�P�[�A^�e�	��B���y�5�y����&�Yh�b:e���ĭb\:"Vd��+��ZS/n˸��`ۆ7Dh�aSM	K�	�L�.iS�aA��.h՛���/�V�<��7.CH;�����3��@C�V��Y�,m�TRD;g{50�>c���$�]VqNS�J����s�a-�	3RG�ל��I��z�m��lh�Ɉ 3��i�$VD�+��^1 s^f�����ƕZ$�ބH s8x��p�;;w%x��zg��b�A @�$���0�*��8�h���7�3�/�PɎ3�$�r@�?4;Et���p�Q���8�����:F��;��o��g�����yؘ�ʥ�Sń�� �3�M۽��ӎ����S��o�˦��M�iJi�=���eњ%�E��c}�o�"��)D{�&�љ�a.�[v���I�ޙ3��z�խ�����0�s�"A-6 ��ሁ��{�4W]�DS�j.����V��Y���qk�5��j��J?f��X��*hi���TΤ��s��CуB�b�ys�/@yܶ���>���v:�c�����:�;`��m��������=/���f]x�[�U<���鸕Y9=v����I9����<$�:�,�t�	c��	���Ep�VX�A1�w��R@���5	�0(%�&X��?ߧg/ݰ$���Ҡv���s9!'��=~�&؇ ���k���qx���w	��D�%��ډ�;�
���}���vp)�2�[��ѳ���d�l�x�i����		�˶d�Av���]R��66�RA�F����Z9�e�aؕl;v�j�M��W�i�I	@�q�{����$����GM�$��Ȃv�M+�����M���guX�o����_0����l��������l Kb{7dj 4 ��L�&x-�n���jɱ ��A����x<��'�[1�?v)o3���af���6�Ƕ�L9u|���Ѡ��{S&e�ЍILc�S��Y��#���}a7��
w�ͬ�'~5����_!E���	�{u;u�'c��q�;S���Mc�/�f�v�xb�����/Gp^��S����J/ 5H�Tl�&� �kc$���7���]������Fv{|�uٜ�ꬪ�/��q$ PL�pj�����0� �i/���ln�8r'+&A �gs۩S�:n�L��5N����`G�~�H~ޟI�@u��<k�8�A�鋵������ -)���⮛fkV��1I����1����ab�@)�c}�dl3�$v�`����ݩ�ɖp���@�M�U�*	$��l�WQ6f��ٽp��$n��R<��0+��N3�x�����n�9}.�Q5�
hg���Nk#X�@�}�cɐ��|��ZY�{��AކN�^ǳ�;��,Yt粍;�>�a��0�1-��$����{�}�=v}dUfU�>��/露�^[(��E
48<����pq�X�a�u��*:xS�Iz��a/����&�ɒ��0�dɐ��G�su? A�����#IՏ�C�8ƚ�I|���P�&!�g��;;�k�PǛ�� ;o)�b_�,\�v�]�l ��Jz`=q�^�k��%�#sFbt%؀���[Z�b��bL��\�H@��������O��4t��%�@y�I]�Μv��7u���$Ň� ��}�˽_g9�H#v�� IY�m�-�ꐱ�;V�D�7��$x��y�Sd���r�J
��I=���Gc�.N17�>d���n���v���hf�� H,Ik��-!�^����(�Q���9�kS��K�H,�͙<���Wr������C�h���\��,Fտx<��'�Vb�$c�X^�4��ɹRw�X�$����g��<w${.8�=Ͻ9���큍2�o1�*�˹�V�Vn��s�"��+r��/6�i�L�����T�3M�����nW#"�LѢ�&B��� 8���(�R-��HRr$X4�6��vL�J�8� �L6������=�qd��q�gc��^��f߸x�c��s.����c�Mq 2/mq��5�Yks�
�s4t�&�*�\�pS5k/]^M��Bkrƒ�W��Y������.řFU�H������dImp0G��i���A�.��J�j+\9��d���n���Z��0�ک�j\p�S+hD�eT%ڡ��%�b���,\�,�Q���jXH�r"I��ߢI���������;�k5޼i�cݗ��x
�M��u���{���tL ��ܱ~��D���TC��œ-��JDI�� ��XoB6l��Α=�WS�ٝN�@��jzgX�
)��^L�s}�5��[Q�'��	�9]ސ|�	;�(�Wo�AP�N�UM���2.=lD�r��7��rz��=��	���aMyYK��GBO�5�|�/XJF�f�f���n@��}x���-Z
h��?��8|̀�7uH�P4���Ueܓ��h[���k�@���)Nc]Uf��q�4��;,�lJ�2�J	gr�[_�JEB���uU��̈́1��S@;�<%����Q���]w���K=��v����
O
��)r���r�%ێS���P~����X=���Q��Gz���}֌��q��u]ލV.��b���bğj׼H�e�����u�]����u�]�����^�$� ��ĀL����&|�9z;}3{� \�f�|۝����*�1ًd���yb��w箎/�\v$H��"[�7�n�`��Щv,ݵoW�U��c�<*����?�+���>��̉��;� ��b
���$�t��cz�,��;�v�6���cm�w�m��^g�����M��NY�>�ֈQ��bO����b5κ���ݧQ��Eln�&�0���5�U�ֲ���rZ���=ݮ����߬c� Ded	:ş��d�4�ǡ�T[K;.�؂aML�\���|�����mt��L�Ěgw�/�cR� �\�X�;���b1�5�l��4֩��i�OߢM�ہ����@�$^vψ�9�ײ")�w�jjhs�D�o�%@���C�8�WF�7��T�=�&'�Z�37bF��$�^���{��,k��[钒�),���?��|��@#ϟt0v� �ko�>��ov۽'wD�F�Q�n��{'(ˇ�7�k���r�iq�{���e��#�R�$�����$��>��L\scA��L����:�y���!A�C��L$ky*Q���#�����ØwS����h���f��Y�B�R�f\rZ�]T�͠�
"f�qAI$�(����XSc��C)��8��51��/�<�ռ�nd[�vd�D��k�=�҈�7�L@q�o,k�_(�M,�����b���`x��L3�Wn�Z\��qw,�����qo��ڢ��9滪�Az�y���^ԟ�ޚZ߻uI3�"���BL�����D�q��5h[V�����J��_����`Ks �*3m�'�!n���4��h~dSW\#5�ZqM��k#���ڜ�/1~_|Lœm�h�������>�_��9ї?��Ie��YIe��� a>j���O�n�'wD�F���Rb�}g��M��M�lou$
gl��������᭻�D�ץ7W.>}q�՚
���%���ѕp�,u��e˶omT&Tef��]��� }���� ���j�e������$S�o(,7i�A��NOO�d�,�A��d���3�I҉|�� �&'���ˇ$^6�R�A,@��M����!	wb��e���q�%m�^�� -��gs�<dt�$_6<��&.�Md H:Ŝ��1w�Q'��߹1vb�ۻ���)���!�9�X�-~�ʻ��\;IX�j$g���`�5-3�\ ��M�2;�L5\�O�_��}D��L�O�$Ưn�w��n>��z~����~�0�����s[�H�V� ��ECC �wo!�Dd����'�>8'f7f�5������{�K�W���zB��{y͵)±���GI-딥7�����̀藗7z��e�����E��V�vn�+��U�W��4�v��9�Ҵ^ӳW�r�I�%)+s��o����ML\����W&�ɛWұ9���G��U�z%q\�⻢X�Y�Ww�.�'w�5M`Y��5�J������-�Q���0t�V$�Y��5�(�8v�5����1�C�jG��m��3y�޲�]6��q��7�m�խ<����du��;���ڗwb�Ux��7t��";�
n��U��1߻��V�y#�C0A9v)��<kfYR����5��e/5����E�Q�Q�����ˮ�G��J�SPN�A�k OB�T�ӏ;N�:w���YK��չ��;�|r������Kr|9WSܳW(�`�L\��su�C��A�Q���Eֹt�z���.'��o�.����]�j�>٘s+��������������n�{
ѽ�st����uV���P�w�O(�Q�A�meUWX����n�[�Lu��W�l=8��9���T꨺�̖���)[�	�M-�J{D��]�@�p}سfm�Ŝ�PIyz���n�ontX���%H@M5�+ǈ��`� �S��6�"��ˀ��wM�v��AJp�R�a��`p�P�0�-+o�lF&]�q������sj��X3F�.��K�pP��e�+J�^�V�5�Bh�wr+�����ɧlC�ȥ�1Bƻ��l���h��5F�D�ww^����R��h&=�������ͼSf��͠H$�[��4)bE�6.�~��h���ʡTS�U߶||_^iF$M4n���y�:a�55�^BO���!��HM?B��"S �$ɽ�A�L�K��
�l�"���J4�фC�Y~b>d�pL���NeF%-B�0ˢ��H�%���ݨI\|�� ���ԃO�~��'���e`�pG�Td$J-��nQ.�H,���2'AQG���RDF� �D0�QTL.aG��/iEf2̴-Fe�k�\N�i{y�N���<u�o<x���_]kZֵ�kXֵƵ�S,�9/'��e����`�T2�V6W)EX�Eq�Y��jX�j�D�b�e-N�'�������y<�O�5�ֵ�k^�ֵ�kZ�X�)mb1J���Z�f�R�=Lb�""�Kkź�b ���NO�s�g����y<�N����kZֽ5�kֱֵ�/'o-
�ZELT]eb��(���(��
�T5�R�(��[e��s�c����{x׏=�}}u�kZצ��cZֺ�9/�g&�/I+"#�-0oW�1Y�T��PF��
�����eEJ��w*{P�IEDH((/
U��4�-��(Ф/|H�N�<�q*ԡiF�R��%`�i��)zqq����\±�փ�r��[{ˈ6��Jѭ��2�yg��)�__\�j[i�nX��Se�0����&[h�V��z�m���BY-�	z�D���R��˔��h���QeiU�\ˍ����+YO�qD�SYӉľ��w������ !�Z�I�����.bdp�X`кk��V[ؤ�Ԇ�m�
���&K�%�m�ɳ��L1�bm�m���,1cA��W���]L�ҜYDa	X��v,)�u���\Y���-�9Ak�ۑn��N����p�\Ѱ�
ːѮ�ؘ����lb�Yn�6���,p�j�jZ4�ΰ��W]���� 4��Ý+\�+sK�ެe��L�����l�Sm3�az��z������G
��̵�f2Ll[t�%�^pՍo8٭\��RY�*6-!5�U���"�`q �E�����GE7X���۱��
-���#��t4���\^�X��B4�SW.��Τ�ڃ22�SF�iH[���!#+�۰�as���Z���[`Jˎ ���\�:�n�k�ֆ��1�J���#uWB��4Z��c8ζ�M�l�I���K����
a�!�f��ڴ�� m�X	b�;��V[��]2m�a�������-u�9qy]��e�HD䲹�e�:���;A"nH�K�a��phǙIZ�x���B+������ԚL]4�TKls�a�u=j:�V��庮�J�-,�ѣSv�X:��#6�5,�&�rlU6�Wlg��e֔fՉQcً��Q�ݥ&�YA�v�XjX�X��vԦ��ImB2lan�3d�H���P�	Ie`Q!k�Xnm�Y��e�F�t*�ض�,�j@��mrp,I�X��-&��YG.�\��©}<�o9])���h�e3g��@�~'S�Ie��YIe��#������WQ�:���a2�ҹ�YX��"��[RE��45[���,B0&,���GX���q�e�qnlUŵ��s�J^p����Yu`J�9��j4��]��q5�.s����G�ǽ��v�mq��;�ƀr�[6 M4"`ֶ��å*�00�T��B�
!l%�Z㦵M�,�V�6eF��Ž�9`m�6�3�h̿�>��;�!���$c��YЎ���v&9t�x<a$��^溜�g�dE1q�h&-�/���^,T _[2�����h��ӎ�P=��消4���ő�qUҨ����dg���3׻��I��\0D�KWv�O�l�@���]���^sU<�R��	 ��A�.��yCHsPf�[���@/����f�Eƙ��@3�hx�ɒ%���v8���i�８)t����x�p^z���F�@�>j^���Sx�B��5�3 )��?wc/1d׉μ^y ������I���?,j�9��Ǎ�K��\ͫ�лG%�K���e�%�6������ݵr���送�;>�rX�Lk�@���!���A��� "	�l��w@�!��|�K�x��int:�������c��k+��t���w-���*��C��'7VL|~����L�Z:�eZ�_W�ۯ)�=y�}��ry?�I�%%�RX�N�ŷ�A$�z�y�I�&vr��L	ɣ�0�ɷ�xH$_�&�:����`�����L��$�u��;�I�L�@�Ia��#���g�E=�J
I$�ESeڷ"�v��jI'q�,H��q��3�C�t"b}���{&9[�gk�.�+�v	&wu���wt�+A�Ęe��y�ɡ�����:)�l^�� &.{q�ܝހ���j=�6EY���0s��	B�E4I�D�=�+"v�1׭Į!6H�:8 �H�\���e��`���>��@�@�ı����OzB�{e��[{��D��)I`M� �7���!�$aT�?za�c�U9#dy������˳��w�w�� `�f��������]vl1i���-�;��xk|����@@����M�8��������]���v+yK]dO�H�w8��x��S0IcE��T���}Y�P�.����nG~�:�����=y��ɯ��)���@�r�o}x7�$�Z���X �A�@�>�����b�	3=��c@@���b�8�J@������2�$�'�N��GYË���3�=�9�'�� �AA��R
Dרj��e�X\TB�E%m��6�f��U�i�b��2�l�2pk�rƿ<�>|�q�>Qv��B�H����bLI�������?a=�l/-����Ũ�2K?rY�E��dC�=�/
5�����d���1�]D�w��朔(y-��u_����~��E拻؋Ҧݳ:E��G���(PaH�,��"I���)vp=�wb�_|�g�x���wgr��1�>n��aT�kt��e�^������#�P*��W�ޏ0%��q�kx8����6V?�Q����Nz�׻��^�V�Y�_о��c�MH���h:�ǜ8�L���k������{�̹jmG`�CH�A/���9q����]u:�����������bA>�����;g�6��g`．��/�g^/���P �k��aE	���o �މ�f���z[ !�t��u&�v."=�ы�Dΰ�ev���Ů&���t�0�'k���$𣝸9�ĉ؁y�	�w�㷀@&L�B$�yXv��l��� n�di�׃�J#���ŕx�\����n�A��`$�@��ܑ"�#��	�{��a��� �!�v�!�t�F�E-L�Xm�@o�/��}�X�#.�i�p�el̂�����^��^;����w�0�A������8��ϻ<�cy�	 ���΢��#��X�sw���v��]e��L�=y�ylI�Ӄl?{�J[~0��s&�1���6�)���Gd���Ŝ�DDfJ~��\��[K�{]Fm��Ʊ�$�ڷyH�I�f���\�b��M�[�[_��G�Wèr�f�����C�u�n��l�b�7�n�粈T߫�MYUM���Ũ�Ʈ�_�>jYf�]e��n<���H�c�vO<Y/�Æ]L���������3�y��y�3�y���ϒ��*i~�f�(�S-*�M5��uNŴ�f�YPWƨ��a,�)
�T�M&I��M���-H)`즫Me��;dJ�4�	cl�iYu�q�m�U�6Vl���B�,���j�nP3R�`kj���qڡp�=��Ʀƥ2e	t5�¡�%�µ5�Qk]�ې$��"a]��2fٚ�U�&�]?�K��A�/�ڧU1�z� ;ԑ�p^|q;����v�� A �u���8� �Nn� �P���]c��v��p��>WL���I&�b� �{�O۹[K�	����;�k�ݸ�9J"|N`3�Z1�^J��D�a��W�l���843�D�F�jc�L_ ���oT)$w�&��N< ���w��B�W��
�L�1rI�bv�Of=g*<�p�Gmh��{Ɇ�t5�^þ���)�~���.&��e�{���v��/R@�&��M��9,6;�I�77����i��
9&:�a	��f�M�mf5�&��u�E(AM�p	�������g���b�Ͼ���Ї��˄�	w�p��S2�D�� �}�s&�"�SsC�x�xT ^Z�et��m2$f���ȣ5Be?�*����b��:�9)Xo�l��׹�-N��V�AUG
��S�����Uw��9_���A���w��9�s˳��]�w��~�,���2^�ΒJ���jg�/�[��O�z�#�u6y�@��@��x�$�'�3�(D@��X��ƕ���۫�Z�[I���W�~���Ǎ�����~|L�����u��.7�
j�[˒v���Lm�p�ks]�����궇~�b��yv�x�I*ou��@/
$f�ɒAb]���|��]��_Qɶ8���ߗHI�w�P�e<;��VOߗ���ٌ��`�$Qɠ�֓Kt��X�^k2۴3k�mr�ʍ��Y����;�N��uz'%2gh����7�@,N��y��!��+��l�8c�w�1����m��˻�k\�B��gnh}���KޖX�l
G�R�	y����x�w|����$K�7)�w���'��_|��*��痩�/��N�.���"���..�C�tUM���OB���ٖ�X#8���wNٗ�a��_�Ws���r�y����{���<�ﻳ,$��}Ő�ݷv�P�q�7�׮`�_�eޣ�� w��ƿK� )��_���^}�vq���A���I3lI �7b4a)DH�ݡ IL����';��vF��g��b+�2�6���c�s���������kH����d�κ��6�0â�$��jX�)-��ˍ5#�mk�Z����߽v-�1��/o�P�w DZdI�r���j7zۋ�U�$�.Nu�l A"�]�PaX�Yݹy;K�jia׵'���oB�Es=���A\�q �X9;�<S8r�E��gmu�Q�S�`��Y]����%1��Ë�4�ٰD�39���D *�Yo��<��B�a�pA��T)!q�m��z��[ ��Y�l�e��:���Ke��:�j�p2�t֪_|���"�;����A1�Q�p��H���sD���dN��܎�8r���&-��w!�dd]<�1ݥ�
H���g$	�w|_U�&xz�,[X�ˆ������ߺ����Ϯ��w{9M�i[�]g�Sbۋmu�ǃ��{qӱb�����z�jb�Ӗv��ۥtv�����LX
��T��PR��X��t�őV���1a*V�$��~k$Y�J0'BIP�檪/����e%�RYe"���x�5�C^�7�Pq�"���4������eKdd���w�#�ZE�ؓ�0��h�#��ML��'VC�8~����5�z�Į%�w �� 5.���kp�\;�[T#���2ҫ7���v���]�;sQ|$�x�nB!1rǻ���1�(�~�bQ�L���oܚ��f�a����ڟ���3��z��B��S=��E�c�ܤ8���>�Uz�_���39|���1�(_�å�}� ��n/grL@�{+{���Yݺ�	'����<y�K�<��ᱤ�&"��ǧo��F��;ߙw;S8�B �;�۷��X��Σ�8�c.��.��"��cv�Br
H���}���ke��'̹��jngg��.���v��� ��� Le�3tS#�Y�~8��CӚXN�Q|�K7�1�Bv4�wS�aNW�x���H�Τ�/0�D��$HՍ�j��>y=M�|�ˣ����h�2٣Gٵ��! ���B�+�gX��O�Ú�L�JK,���K,��η{���K�k ;�vyZ�,���h]ZJ��F9��I�B��݊:&[	qFԡ������Yl.�1��du�tQ��ƃ���]%S �IFƱ.;�L嶲��-��f�f)s])h�����Hmuͦ!Y������t4�	�����w������×km�hG�쀻f7 �5D6�QZA�I+v�\B�	9JF��{�dbkR�y��-��+�(P�`��ID�r%U�@��%(�oy�]ɱ��X��m�i���HcK�3��H$0-�OZdዃ0"�j;	�y��T�r���0�c���㢖1�gŴ�GN�g��u�q��\`d�1 V_L� ���$������N˚��q�	������$+��FA$�$6�$�ßw&�qz��N3q��^o9ed�y�c����4�@7��6�&�������q��f�v�r�X��8�͖\��!��y��ᵠ�;k��A��TOW2���8�36\��`nv����aM��p��{�{�
0�/�F)ɒI ^rdE�w`|ݼ����-5��F�ʆ���	���l��ۨH�.��_�?02�<s����C�n�Z�L��)�]W��F��g!|n�g���>��H�3(�,%��4.����Tr�7*�C�/1��_�>���w���Fl���K,��������δ� v���D=,�@��5<�˾Ι����b��.���f�h�R����w$X�3��1�S�I��x�9�����r��m�9��v��xx8<B^��<�&�����>��~U�,��x�J��ʕ���޿�����=斒� ��9��
)��Lbê�X8�	�<}3͐	ʤ��؀{i"I{��vl~�}�i>V�e^���j��(�l!�J�K{V��Ѹ�uX�f������{ٟ'�I�98��aØ��:�N��R1txl��Z��촁,'�P�2�@���_ �"]��l��I�Ow��}�H�@��1�읡�_\0�n�L��}Y���ԟX
+�Z]�A$vwn8J�J^�9��Њb����K@g�P�ۻ�#�o���+���)��wv�p1~�bN�5�M]X�*�j�p۬��+��B����a�Z�:ɺ�'l���!�B��X��qL���$��]ݒ��2��9�g�Iz2�n)���1�M�T5T�C�tyϒ�b��F��XN����I=��%��s��f�@�զ��u�tc��K������佦*�&�Fɴ�E��4�I�\��f��3�ΐ�Z 4���ok!0�fa�r���Lr����yf�ř�̤v�؄��䫫%7y.��R���z_ͣ�=��l��a�3Q�ngbJ��C!�.P��1��[$Y��.���L:��qr�nJ'��mc��A_sv�S��r&���(�#׷�05�S]��T1B��:��c��c*�eK�n֦����B��aL�o-z�=5Yn���a�҆�
�AZ���R���Ս�]u��Uۏo+2��a`���aƗ]g^٭K/�Q���Ү�L\��{~ٺW�(�;y���-��G�[�bnR���n�+*��{����Ҡ�y�9�m��튗;��Dm��w}����|��ϡЏq�=~Z��Z��X��u'�I�d�|�۾��͠{�y"�ô'l:`v�x�wIN\Vf�'iw��R��N�W��<CXE���$�5�f%���a�!�:���x�И����q��#��t�|��(������Ôߨ��R�T�`qK.�I�{5���L۔w=sm��n�mL;����|���ߠ�'�S�V�Ҡ��Mű���h�$�_����u���׏���Ǐ<x���ֵ�zkZ�5�k�c��%Km���ɜmB�)Z��bʕ���5>��
��A*�Y�=�O��<x��Ǐ>>��ֵ�k^�ֵֺ�������w�*v���yŲYyeX��-b�Ku1��iC2�󜮾>>�W��<x�����kZֵ�k�kZ�=K뜲�/8哓�`�1��p���q6��;J���r�휝u����^><x��Ǐ�U�kZֽ��u�kZǯV�rr���r���R�����v�ܻ���򭅴J6�[K�W��jPU��r�KFVV{sV�-�3
=��G�1����k��T�b�[jkUĢ�(��EeelJ�Zc*��mWш���F���F�-ۂ&R���F��*�+��^5έ��mTU���Z�[H�ڠ�9m}�,؞f�3�Pr���)W30�U�X2{�aZ��p�J�ڪ�(t���73�w6RYe%�Y,������ݯ�A��Ze��M������@��TǗ/4]��ՀAy�;��P��;8g�;�O��xc�{���T�>�H �L���L�7%�:��>%y �g��J}�8�v<�Ͷ�ݮyi������=�v=���N8��ד]�7c�{:�j��V����LWj�[3t���u�s��!�$D@��5z�F�Ix\1��1�k��T����D��㷓����(#N�PD�����k�J�b!
�<�!F03�v�rV/�!g�E��t� Ӿ�$���O;�Z7�1lR]�{�{PC�"`��{|<��jb���s��]��h����LE6���ނ9���%���/y�������@ח����r�U����c��2���wj7�T��v���US��U�V��5�+�,�m�dT�`�p�ɏ|�8\=\�ܕ�O�f�O����^��e��Y�ٿ�������&v��<7!a �v�
�v�Je����g��@��@Gg���m�,9NL˚rQ&
����b���� F�[4]fYh��5c"]"�pko��9���n�v�	�w�R)�Ļ��AU��k����,^kI;��-��ww!��΃�$S±��D�ޓ�w[o:Ey��3���L�C8aW$2������o?�w��T	7�6,��B��å$E3�}ؒX�LT�m�S�{�!���T�$\��Uu;�x9�1�A������5sr�g6в%y��ǽ�$�9���� �0Ü޹5�+_,=x�#�j�P��JT�:���{le�+�M\>�]���y��@��54�.�s�ʘ����1wG;}����̨\���GuZ�e~�E;�A�ޢ{woYɊnޫ���>퓆�Wm6�ʬ��hg/����_~��CWP�Z�m�R�|�$4���QX�"�b�R0�=
�
��hB��.����H%̶"�C%�� "��;�n�Kש,���1C޷/]�t늗r����+b +)2���k����R#M����K�%��R�fQ�e����2.���5 �l���b��67������:��[HgL�n�1�)
�Cf�����C���&t�r��ne���9��-e�J&��5������d�r2���u�ť�I�r��==��(�]�ZU�m.�h�4��nc@�2�5v��<�O����Dh)<X{��$gyh�Rm��9ggv�]0Ɔ͈���
�sy��A1��0ϭ5v��	kcKW�"m�����kv� ����H@��\��1g7X4��w�˝mz�K��6E<)�8�|�{�.��sK}a���C8Lu���$�@6�dݽ��;�.,��B�GBv������xF�9}�`X�b��ِK0n�7���?�^�`݊X�q�A�s��_R!���h6���Ɗ�Gջ�-�1��kmx�8��hg������;��9�tp�Jщ���X�ap��i��b�3vb	b���&����4���"!%��oK�P�c���gd-��vy���3j�}��f��^AnoU��{�l ����A47k�OOP��c����ש^d$����i�H7;��JtwNa�U�l_,�͡&"�-=���7m3�2��E�,*�3�}w��ƨ�ˌ�b�AǬ�_��%%�Y,���)���|���0�ś2I���3�1�Tz(��"��1p�k\��"!/SsAۑ!��vd�Av�����{\������48�pw&���]!M�U���E<*� tL,=�q������T��q`	 �a�˖b]���EcS��ч/�3��S�����^b)t�[�=�*$�@�B<�T�[��[�6�K�{kR3�=R��4�ݩKk<T�ސ����87|��7^->�M�w�
<�
XЕՍ���ap"m�YEZCA�����F#��N��;�;�>�C H��4��Щ������ ΒM˫��� ���Ad�A��P�J��a��D[xɘ����d�ë�s�5B��,@ ���Gg���h��. @�'�x�rd3�C���}^�K/����I؍Y>�P���w��{Z`��N�jo��ϋ��d��&r<L^Μ-q���g��ׇ�����s�K),���)+;>yRv�wnqِ���+w��$���sp���]�����덗�lq�pY�D#.�W!�.%���Q��|�a���:t=���)�{�"a1����!���==.��O_1��5��Z�4>����8�^f����$|QA57��3-R[��X�K\ͻljY��u4k�d>}����1�x9�K_B���wt��P�>���͒�Ϟ\�� ��:u��F"G�۽^��0��EUk�lCl��E�R1\��7��Z v�:k��-�t�Hh��R �x%��^��I R���Z���9���RI`������W�ٰ/�Tr$�z�"��@R��6�sx~m��
D�|_i��޿�`��y
�H�gz�� �gnρ ���:0D�wfc8��z�22�ѹ���!�/��Cx;�QY��˦�FmN���8�g��g���|�侾��Ʒ�!�k/���h���g�1���zg��l䤲�K,�Ye���o����8��}y�`���*���7d���U<2�n^��j@�c|��H�; ��ݞ� ���!�r9<,k��r���l�3^�#4��tl�#�7X-*Q�m�fTm�82�-���_��������u5������w2��v�քI����k,	��h^@)f�I�t�a.���0a�I
�
W����5�m�h{��Wx�)u� s��WA�Aƨl3�
c�9��x"�I1�%��'p���1~�ɐ\�>�+v��{o��$�-���x��V�� �}��,��i����X��؇�M�[�t7��:�#&�4lD}�Č<�9��/,�w)Z����,��^� >��;�H\7�n��#�<�+��.ʭf�@���P�m���S�@��ĕ��pN.��f��yY�Mfn��ɠ��BHYEbG}�i��c$��6-
�#�-Y��
�p�h&vT���Nk4۲�+��eˡam��Bw),���),��΋xެM�ܵ�b %������X.�]�mٳ3SE�c:��UI]�ŗ$xS^[�Li�Z3K5Ҫ�VUav�J�K��l�A�4!���j��)bnm.�D�,[\0�m���BP\����k�V X����g9� �lP�G6jUD�$Ƌu5��A�Ф�u��Ձ��U�:ˢ%�2��t�q��pk�vb���ϖ�a�����e��;^�n����7�Mע&,K�3�o��KK=�M�gU�;�@|~���]���D���/ݮl�d���)��x�Y-��#��<�o{b��\T<\���9��N���B��RY5��p�M����c=�H�Dײ�K8���@��
Y�[��F"��OL�=/[��7� �Sq�1�i$OoJ���/q��.��+q��$��^�I$
R37��d�	��@S�w���9O����y�j�L���q�����~���}}���=z��`0	i.8.���P�	��I]��.�)�G,5��`���iU�>����C����I̸1�	����m�7����Q J�쑃�P/��7�� ����~����ijh�R��q�����0,��Թ��cN���4o�n����ƌv����l�U�ZM|o{��K����p^���F���RYe%�RYeX���74@��7�<��n��3��@�wL/@[���Zb���⸇.�ü�������Z�i	����A��g�8FUp�1�ϻc���w ������9r�}�c	tD!���L4�n��>�iP���au9�y�c��]�,���_S���Urs��%��Ә�.����|X����Δ�ro���`�l�A�i����$�{���1ps�7�s����_n�E��*�F��eR�\g��p�:�	�r�P6p��h����~�ʬk#�|����
gv>b�r	b��1��ӯ��]�^���yߒ�+��˿��ya��+iQ �f���<�5�2$m< ��Ь�V��M+�ޠ�݉�I7h�l[�0w+�آ�i\�z��x1�<%�����<�$��HH5� s[`R�|�U�Ē8�m�;����*�\�W0۴�.���<�]zn���ڛ^���ا�pjo3�,���),���p�^P�������6j+�$������Rnh@l�r��s�!�#��RI�-M�u��м�� �8W�35v�|C^��
��ݖ�SĒ/���%0a�nu۬�& [�x�r�;��ɝ�M3���C��rS榄H�� B�3?~?DPEQ�[�Ҏn	\0)�q�hۍ��饌)�I�)�=�2s��m���1�7��Ē��Ah��t�f�����H���c	$�u"݈ܫ����?s[�
��~�����H�����,�����&0��,���o	& w�$���Ͳ�"y���7_Hu*_�S�)�[J�2��_6䉿wx���W���3�1��gq1���X����G_HG�tw�{�2�.@9��$w\�~��Fw�JJg�q�#&�z���T+�|�(h
��f��G.�ٮ4y���N�[ʋˉ��F��G�6�)�O�e%�P,���b�]n�r�f��C�H ����Ћ1�謟s:���E_��e��%u�9����=.���Ŋ�v��;�Ȫ@��)��b���MCZ2:a��#`�k]u�j�씊�u�3/�S��.���\�%��!67�x�|���H<�Oj�$��\7��3�g}l��b<;�����p"�0=r~�������wժp|�t�D��pO�-斀[��{�@���@��FŐH=;[�RI@N�sCkM3��j�\� {��J.���w�T���ݨ"Amb���e�2���NRx�;���{Z&��-��w����#;���~��M��ƪ!�����&�c�NL�����'<�G;���p]١9�a%��t� Ky�vt�HrI޸�1��K����{\D\�7V<�ZL����-��:4����eL%<��̝8U��-e�Bwk��\^�����̳՝2����=��8�ڍ�MO�2��R�,�4�h��d�B��Z�t7��.�	��nU�#�.ѷym=uW���K�u4�]�ԫ��VLy.�/���j�I�ZMo�����G:x�yR�U�֨Us����e)�����eY]���y�u&����;��È̄w6�.�eɅM������}�.���u ���p�q�b��};�;'��,���E���ޞv����b*�y�2�^Y��5Z�)t�/{����.6v���;�k��!��j��崹T�a�݊
k�o�܋;q劶�
ے��4Z���j��X�\й�����j��Z���Ǩ�Ʌ�*����ȳP\a�1$�æ�w/2o0]����ܾ�Cq�]%uk�k8q�mE�o��P��ˮ�C<��ܮ�|v�����rW�^[Ofb�r9b��.��aN�5���׋��[sj�����R�R)�VK�#�-�v���p�#Z����]f��'�/u�l�ٟs��؛����PV�H��,?I R
���_K��-�nk��J��Q�"�2�w�k ��T~�{���\�~U==D,�B�� �A;���$�:
4)TФ�8������u���+nꬂ.�������cIm$#p��[�RT��
~o@���zޭo���05SD�e��D��N�Q&���	�Ҫ���UK��u�2œ�./a��0��W��0*�%U���u��Iu��D�j:��e�~ʲ�4������Cm*M�B,6�r���PϋsiR�JMk�λz��Aa��Z�_�E����F��S8��\փ�B3�T�����MO
5��5����K�齟�\�W1�ͥ��o߿/��1E퀫1��T�ĉ�齭��o{�R�/��R�$O�Ÿ~'�z��hV����DO:UbʨMC#��`��l�|�3f�WiJ��
�E���Yb%.v-�M5����!lX%%eUE�#mF��Ŷ���9*s��M~�W�Ǐ<x�����kZֵ�k�kZ�=-�ﳜ��U�lq1��b,k���(y�E��!f�pE�������}>����Ǐ<k��kZֵ�mk]kg����åj(��Z�1�E�ڶ�%�C��U�eF�ap�����_c��Ǐ<x���Zֵ�k_�ֵ�{��v�e���ʗ�mʊ��kj�-PX卩�3�Z�䯏��}�<x���׏�ֵ�kZ�ֵָ�c���9/�����XS��*m�4c11<Mq�Gm���M���SPG�M���'u���֨���n�mv�E�VcG�Fc��IP�k
���j2�5��J��Y�k�X�c*q̦����+�ȢʵK\fR�z٬��!�u��{n��TzP��a?l�6H]�Y�*��}i���;W�؉����n��sz�v���,f̴h�)��6�W`�n�8�w[��I��ƍ),̷����7R���a#	���P]j��bթpe���ډvLJ�,"�\���
V����z��۵��TnWVʻ
ͳ�l"�q��x����FΥ˚��-��T�1��Sh��]6FT�t-���bh+����bh�3mv�3V�Ъ�끙�6�V�h�;[,�ڶح�:�(�k�0i[�-����v�s6���a.�lK��"�hƋ̮�2!3S��R(7�z���խD�`HlՐ�c�K[���3.�%�lI�+Yc,%���xnrK-����F�u�N
���oUP�:0Չ��F�-�M��AE�.ĥj�c-jlMK;i��%����3���T�x#������vu�5�z�B��T@n���\��ݮeJ��M]�e0�d̼�aS�3D�X��5��f9�K-���.���]���뭁��mCjf1����#uk-�i�����`�v�lX`�*;]̈́!,E�f-��l���γ8�XZVP:V�;CQv
�����^BC]���,,.Պ�8���k.�]�"�Z���35р�,ص��T]5�1�L��r��2���d{1!�U�(��F]k.ĩm�����l�.�,q*V��ZD��k��t�1��Hb��u��ֶ��-LU1fe�B�r�Pt�a����s�������t�V��.ɴ���g�)�M�iZ��e���w9�<���RYe�e�w�k���o]^�t�so���,�}���lJ�.L��� �ʸ�����e`���<�e�x�m)�b�i�ڌhQ�����+`�3�d��4�/2�)vf4͘-
X�5&�i20���Ĩ�\b�2^�lB����tuR�jĉm�J��ͣ�V��	�Z��V�fJ]\��lʹ����/Ӥ������;��ҏ�$�9Y�������ѬSJ�.=W����#ea�w&�vKK��;"�x���Ǜ�Li�D��<�}\�ֲ�b�ǹ@';�Mo|a�z���-�� JPP�#�S1�λ�;�9�8��[����>��)����)���)$�'R(GDG��b�a�e�?) ���X��E���]��״��u���]�O�]��m���$]_4=	[ �(La�������|$�]s>��Iݔ�ig~�R�	3�����X�Z$h6�Ry�)��.L�u��RZJA�K���k�#p뵖Zmg����`�؊[��F����8	�&��C_saxX��3.0�^v�M�����#���=���y�3���֞��{�)E�F"���n���L�\�B��YyWy�j
�s�LSVm�9��\�DX�YǃZ�_�@�j��!�%E3���d��C!�O���WfK	bw܀՝0��CE=\��X��b t�
�L$���G^B�M��E�������A&�xgs���ܷz@�P���z��>��[�vy0�_��Y��9��SтكW1 _�z.j�:I�R(���y�Ґ�U7bbO�er���"ZY�q]hsK<3��#�!ԏ>�[������z��"����U��b�D�e.�7t#V�++�afF������Z��~���_#p'=�2
d�in?6�@�Lc'�C��Hi����xJ�=�L�s7�؏	5�։���i��+g�7���E������neZj�0$�wJEٍ�#�����R���w��M��EbKm�f�u��%P|�T��Ke��:�C:���kY���:�n�땚�� �Ui�7䤧�<�,C!����asٰ$ig����(7�����t�
�y�.Ӗ ��앬|3�0�3�M���㣭�S����� �����(�
>�/�H��K���>C��7����-R1И-�wׇ���N��m�	��jI�D;g5���y����e���i��h<lG;L�|���r�{���I&�9H$ksD����/�.�]�(,������A1����<==�J����jpY3�_��ca����Ms�O���������v�$SNgD808C�UOU�!3�vw=�� ��MF�t$�� <Y���F4&$/��Y���w����4�e5�w��	!)I�c-��������}D�M��1 ��HH&[7�gK߫�<��|;=u>z�ug%�J�{Ҋ6��eDK�ը�WX(K���N� �A�G ��C�h����2��RVOizy��K1���Y��L�/{ν��-{��#��#�"� �����a�!�Y����-��7��] Z����r�g}=y}M�oUX��Ц�kM��M���[l)WlCS#�X1Ch"l��EZ���w���* �!����4��И�����Ӿ.	�.ע��D��od*g���v�9"f)�ܟ~p��j���}�X�O��XK�� \3�����Ҫ��dH�h�&,�F$y�G(g.b3�2�3��gX�r	ؽ����32�����/�%�(_���U�myՠ��	�����]��d��k���	9wJ� P���L1�X�6Vh��n<�܉������r�:�O�����{S���a�F(� ����{��O��2�j�]��J]v�꩟Lm��Է�V�fd7�F��R�P�Hj������V겠�IFW�X����}]P=���@�XW��u���ޮ)�]�#1#1R+���QDS *@�$��T�5x%�����p7	e4͸��tYt�J�j�������eLU�1�[�W4�IkuL�H�fZ�Ѕ- ��š�@�!0R����e@pcI�)��K���d��JuKYSi�g��v-ԂF�Z��I\,;L��]\ٮ�?Od�G{/�)K���L&�]"m�]CWF`lv���:�e�n���ϛ�:�����Y��v�ɯoM����Æ e3�zQ����"Xɮ��/h�
#��[ �}N�g	È,(�� <�Ckx&�a˺B/M�f����E��up���!BI�R5�]w@@�;��)�5�l��<��/zpDN�	�������_���b�F[M��k�d�1B�{t�\��+gO`� �i�9�Y2Q,���&�C���Ͼ�X�e�--m���A�	�J���2Ky�fd�߯}�قc�H)T��AM��>b	��i�p��~��?%����#kĵj��
����A���b��0�u�4%Ɗ+�6�jB�و�j�0BN]��=�S[zm�ω$Pg��vA�sקw��6���0H/�ڹ�F�U���P(O^�;�'[�s�l�O��~������O\(�}}�v�w��ç�%c[�>��{Z	|�*u�yv+��2�K�IO�(@�C|������$c 1#����!7�s$�Ow ��wc�}�"�0>��ku�e��	Q�X������b�U��z�+�E���5Q�#��韷���2I1K�<����X�uѿ���S@��|h]b,��}�^�8����j�mj�n�d��9�$�G�F�@1�<�/ؑ�ъ�Ow:��D�� @{[4�	~���rh�*lR�_}3"1SֽQ�$h"����ƚ�K�aZ)�P�tʲ���L(�y�~���0Kr~7V�X�ى�1��ސ��K�F*�T����'����ȊIP<����;���ѓ`����_3�4���Y�z�g�=+(ڞƇ���.��m���T
߁�yy)jjFؐM�v�����𪯿;��Ay�9ͯ�Z�k[-�������K�[c�m�/���G&ՊN�nDD��ND�dbF2�3��hU���h���L����D;��i}@�P����.(b�SZ�n�,w��A�i�CX�;=5B��Iꮇ1|	�$��F�z�D<A���P����n�Y잻ukC>ٺû�#��[;���#����;��ٓ�����������/8�@�q���Q�f��S���b��&�k�� �\lՌr~}���ho�q����Gyq�6� H�s�ܱ����z!s����4 q�{���b�����w�'|9�� �hz��g5�vy���y鳟��:ْ�2h{0Db���u�b
��Bq?r����=}��t\$�|�3,I�5�!'.�H�ꣁi��-�EY�I�>��H=�u�޵<��/�\���d�y����:ĺ�3�T6q*$�;��&����7\����Ҹw�`��lt@W:EQ��{�9K�t��y7���j�Nݪ�w}պںB[t ��y���̌H�������~��-�E��D]ꝙ ��e���y8ȕ�Z�OM"�Pc�جhhOt�����eB���J,��Q�	J��E�ԙcs��f#A�sҪ� �G�^d ?߮W\5�|�l;Vn�c\��'gJ�����A6���>�rz2"����������e쵕��g�ܤ�l^��"HL�2��������<w�ᯀ��K�S�u�t��M��	�σj�kQ�}�˥mM�GVd��gpv�#^�vob8BN]ґv2�V�5O��l4�V�i�߱��r�D�97�9�V{&D>�w�st��N�+v#� �s&M�g�Ȑw�o�FyMy�I ���p�8r��Rc�����lL�s�=�2ǡ�P�]�V�n���x�۽�꼊�;X�����ۘ��WQ>8�CK˵��yx\{aͭ���f�����+q}I��%�O���>eJz\��ڙ]u��"�L�P�+���0��9�q��� 1#1��%��ŵ/#ZL�,�p�5��b�[M[��%���s6��u�R�<�D�<�r33n,�L�T�@���`�A���9\�M.�6�ĺ�R^ R[�)e�iR5Q�f��i�au.#��	a���)��+��(M��ŻL-�������Оqf��@&�	�l.tH��`��\�-�[n�ډ��)�� (0�9�5���7|.ne�|ޔI$o�0F7���Ex�t�I��K� �߹�RPK�u�,�H2�'���?t�c�^�"��2��G��O���&�)���Ŕ�"�c-�����M&Wz��_�棓�	���no7��zh]"L� ����O@%�)-iGK��,�J�c��Y��$���;�&l޴t�=�W���g�Y��N��I ��9���Z�t"�ӄ�O��ؿs�Bz×	:܍��>mg����/q�6v���ͽT��綊1�&#t�a�.�U�6������c9���܁l��S3���+�8s��m�ޛ�b������M5K�$|�QI]��c�c�'y��>�K�� &>[�l�Q�G�����6�G��Cee��AΩ۔#���J��
�ضov�[nm��;V�����GӊU��S3���o��dK[���%�<P ����x�owt���D��}ĒN�JR06�hY� ���U��3�j���^�K~z�H2�=Y�!��)�E����GFb�4�,KU�rn:�NS8~�px�Y1-�b)�G6��'P%�*�����>3��Re��CП]��;�$�r�b<���Z�L�A��X�cӏ>���4�e@�"!i}�W�h�\���f��
��	mY�H�6�����_�lFBt��R;�]B"��b3:T�a����:ZE�����=�܃Sћ������޷8��N�cP�1rg��
��x����:I0�b:�_V'i{��$	����#��'nd��ṟn<�'��6�iy;��U��%��,�C��fn�V�u��3��*;�Ƈ+8j�z���Σ�\UX�:��6Mi��,d�ئ���ӝ����v�e;\,Q��^�*����V�����S����ᵒ�KSXmJd��F�ja�4Q���z������4h�nF�����+��E;�b��y��3&�#�jgw�vRzl�s:��nbY!�F�ث{7j	�o{�I�YR*G��צkC�%�CH@���}w&�yWh-�ڱ�uA�X��W,�������j��<��|����.uV�uv�8�q�w�
��S7�s���c���5�������|��݈�e�G�%k���������ĺ�
�BH�e����:�w���"nh�W�
�!̼}|��*��t����x�Vf]u[��i4�[E햬�u}a^m�4�^��̞eok���\Q��~ҕX�h���`ܰw6����/��*��^V����.@��6�g�C,S�ܺ������J��vor�ږa�'��9ݭ�K��`�ս4ݡ�85c��;iW\x�y�
b�����;���؞Y��$#�kz���I�8��GH�j��T��M%*��l����l{�����%�cX/:�أ�i��:N5ٶq �Ӽ�T�"}�3:9�H��L��L�$�U�/���E��]ͳ�T�	��	�Ax�^9cڀ!l�7�`���`��/o,��',�kƵ�<|x��Ǐ_[ֵ�k_�ֵ�z�_\�9=���`�cEhۙ��`��wr��g&eؐ1��������������Ƶ�kZ�ƵƵ�k���> [T���4�}��Z$��z����j��wt�8�Yd�����<x�����Ƶ�kZ�ƵƵ�k��[l�����S2��Ic6�n5��9���*�[-�3����c���_c�^<x��ƾ�5�kZֵ�U�kZǿnNs��G�.Z���J�#�L�ʘ�,B7��A Ykwݞ v�.��mV�h�6�����p�����U���E��db����{���\h�ȣd��!(�'�v�j��%�V�W���R����C�!��\�k�TX9J��UeC�j�j�%�+�)�,E:KǬ9�r(�Y��k�b�a�����|��)�N�K��|N������@p�y�onxCK���ֽ�ڄ�w�R�ʣ��.�%���=#g(�o�K�m1Df� H&��І鳾-�i�-���H� �'}[�!��)�Fcc�t�)�� >�B*0v�KԳg�e7CfC�\�XIL����nހ��=���t�q8"�ղ�nݑ�{�98��mk�kGnF!,B������@��������m�^�	��9����V��y�A�n2����О�K��Ё'�}f�����8x�͒�uӠl��^$�@��&�f���[�@ޝ��	'�{�� �ҿlqy#O�-�*r�;<T��T�J�!�w�	c�����L\�v�y��A$�f;��]'O���g�G8y1��涟@rN�&D���]��m�_z�j&3>J}�*s(l���+2�^U@OP}6���ח��W��;������l��JS�%�1�ŋ,Y���~�e\	9��I:N蔨r�v#A�V�ϊ��>����B�?��0�=��3�ow���T�y}ߴ0�A��T��f��TA5��a�I��.n�\ӗ�ї1����������ٵ�������dȱv2ז���= ���NL1��v�tfT�[�a�SG�C�D���Ue�������TOuXD�|�ײ�>mm��I�8��,�A���I���ОJ�6��u�J&y,V���8YS��g�	=���y_�r;��Ie�=�n�(Aӥ|Ķ3�M5�NkE�^�Ci3���Gz�I,I��q9�p�ȥú�^O����H�E� ��;��]'OcUԉL�{5�J��5�G"�c���z	��F����Λ��{�r�L��<ia�GU̝[�dܔ/a��_i��b�k�>�\��4�
��*�Eu=Nd�B�m�(�H�\*2BF�/(av���|f�5�@�YUz�y�7y�����A�c�mV�T����؍u��f�4����:W<CQX��a2��䱵�(�0tڲ�f�˴flĊ��P����ʒ�ame%n��-��$�,b�au��)�h�4�L�M��WDnGv-�uHܶ1�R]����:^ SSZ�,(�
��\A�sk5��L%�H71%k-!-12���r�=��3� �Z4�i�B�� E��$�'t�-��aɠE��gv$C;��@������A��g�7�<`���O媃k?,�H-7��w��c����9��Cx?��D���o�(�M��*֦�fG8�	H�L���$�B	�wؘD�K��\��x�&{.{��MX��P�mVl�s� �J��Td��ЌVR ���xgsҤk8vvwv��ox�K���W�]ϱg:b�"�![�˻����J�N���WRR�c��&�ϭ�$f��K��N3��Q\X�xwJe�0����3ُ΢����*��[��)�����Ś�S5�UuJŌ>V��t�������֠�;�@���认�[�OL�X��q��)B�47{���8�:Ss�N�����e��ʰ�R��>�׽y\Mf����zHW�í����嵻��摅U�wl��#��1���w��/Q�����>4tL	#����������3<I'��`���O�-�j�`���M��K_���<�D��3p�趖x*�9�����Cc!�o�y�~�ʓݾy��o�}>�=$DH(�����L`~�w���)����~���Vu�L�48]��I3�#���R1�]�Li��mg�o�6�T�3�!��[�]2_g�m�	�989��,����+�ffF�P�f�@�yښ-ff����tX��aB ���D¦~h�!��#ѽ21��1�����'��=pYq�Ekc�"Z���|��x���6`��ny�ا����]�S7�	�L���L�A�|rE{�؈�$�;����N��S�s|��;��^�ihg�;s�C����{���k�̲֫y-+-��*�I�;ނT|��vv���EA|�����Y���0](����?$Ւ��UO;��?<rl���.��W&��.]���|r�#!�_9�]��7�-����@�;�U��y�w���S(�n�F1���Wus���Ht��׉,�'\v��ԫ�Q��`ʱ��	:�hF�zd�;�kz)���{�b�����YK�34A�� kV'(ō�kv��Y�h]�9Ѯ`A1�ϣ��v�uI���ƪa�|gS��z�B�\���əpW2M���(%:t�������~h�9S*�x|(�A����j��-!��ɟ�}�^u⣲���--����t�<U&�������r�v����s�]����:q��ܲ&O1�l�vo��:tr��yDD��N�ύ��}�S�A,H�Yd�1wWa������눙�^[R*��8��N�)�u[�f���6��a(%��h�DQ�o���{��?�c �B`��u���Ԫd��dD<?����1��`��\�-��rp���j7�v��p;%k{Ē_��H1rw����/Ӄ}�����`N�*���[N@1�P��\�FQ��##	����O"C��KwRi/��䎫AD���&�B�M���D����+i�N��VE�pxK¿[;�� �j�9�^��|���A ����(cR�Z�2G�p'�� �=�l4�2X�{��(%:t�c�K�?l@D��w��{�wcټ� ��C{�˻���x$����T�=���}վ���� ����"s_���Ր�a�H�m����Ӻr�F�Ё �]��s>3�U�<p�l���*�ឫ�I���;�3䎅�S���\�]�^'���+���o��]lͳ��lcT�	s@��J5��ly7w���� Yו!KՊD5K�!f���j����O���A��ԩ�wf�5i�uA�Hq��e�g�\�=e�[���~b|��9���w�:��1�H`s/C˦-�a�4�tjp:.��
VhkX��B�Շl�hmh�N���ntq��ftH�l"j���u��m��iH�Z�ZPd�3�q:�A�M���/��XK!c�I�H��`R)��x�e��eWl�ju�� - �(q��*Y��X��RP6���6[��,�!Á��#�Ķ钪ͥ��-��X�,����τ���ʈ��b�ZZH�w��ȐI�v~�k�N��96��&�gK�{�5� \D�	<��ԉ/8�ާ�wfyܝ���A��%���������,ײl�#�"�E����0�Nwx����;��Ǯ5⇙�p���Y��T�gih�Mm�h<���MAd���%�A �V���� �ҿg���=�����������A�KV,�y��\�ipX�T�F��u��l^��������IBY���p0����)scxA��){�;{7б���?oH�#�"�3����2}��S'Di.��ߛ�)Mc���H�̱��*j�p摫DQ��^���"�t�.�p���a-��r��`�a��v!CKU��C�����$��Q	�F6����o�J8��3��*��ûR��u�ʊVA}�/o+2�:��w.�^��5toN=�t׈�W���ѻ�~�?Œ���1�>f��9���;��Xmi�gx�I؃�8Muv��$�y���>D�	H���H���Tvą�	/%��P� l��g~g���?�h�$�ն�s�LB������~*$�NO�h�����g3���/��2���4�H�%�;�{w4@Jt�mQ/�� �z�5}ڸ8��o��b֗	�>�$��;Z�'�8w���D���,��~˶�E�����&v����F��.�[�_>�}.�a�]�}ߞh1�j�.kg�'V�M!���Ix����,��Z@Ư"@��u�$S�r�6�7�i��͍ӾR'k�F���8�Ōd�9n��$�l�n���0e���NTDW1����\�	 ��uF�v�G�9I�y�U�ؕ�,�#j��'{E������H�Ⱦ�9[�1���Y�*�
�-�΂��G("|@�ƋK1�c�������*ڿ~�l�:l[-7)�˾�npyJF�<���}��8��leיc�w�(|�^��^C����A�\MH'y��\�����s��&�9�%����9־M����E1���v4hv�Ս/��}W�ϰ��~nG&(r��(Ŷ4�ն:�!kL�������b܏����Ͽ}�2�~z��1�4��_�`1�X����wpO1QNc���'һ2����I{��X1	�@�02��%ƭ�Y�$'�C�89�����8��[}\{Tn6^��H�t�+k;,�3���
��Y�}�y�yc\�Hڴ[?�diTg���>9Q"�����(I��3�]	vc�)����}�s�����}�a&��ėWf�V!H�z��s�=�J�aU�$d#w˧p�x��?nui��ˣ�1��I�><����h�}���$$����$��q7�����-��ic"�R X��V6MV'/ٱ���?MA�m����~#�Ik�rf���qpJ��� �PT��_
]��7�i�gנ�Wk�$�l[kCD<i���(c�����!�l���-~ɟ6��W����:WTK�}�HDgw�����]�5��k8��آ� ���z	�(�����٣�߾�JxIr(�}oH ���ԗ��~0O>�x��޴�� �g��K�&:��$S�r�X0�<��.��lg��I�Ts��3Ҵ�۵y��^)i~m�ܺܯ�A�F6�m�<���w���Cg����Ty("N�ñD�Ȧ(������~^q�@A��H������)��"A����-	$$�8uvR1Č9@�"�b@�b�c �,�*�@�eZ�$��$�,YVX�I$�$�J��1H�$ bB	����%�-Z�K�"�X�i �"�bX�	#�H�(�BU�*�U�*ʱ-Z�Id�V��B�HŌ �!1� �X��R#B0$#�b1��B���Yb�YD�$�,[ȤU�bċ"�T���bŋ !A��R,BD���0$�E"H�c$b�D�RQdT�ȒĖEI,���X�!�$e��D$�,IdX�Ȓ�ȩ%�E�adX�Ȱ�(�,,�,�YT�ȱ%�RK"�ȱ%�RK"�"ĖE�,��YX�Ȣȩ%�bK"��E�,�YY$�*IdIbK"��EI,�Y$�(�,IdXYȰ���d�"K"��EEI,��dQdX�ȱ%�adT�Ȓ�"ȖE�,�"ĖE��Q,�,��YYT�Ȱ�*%�RK"�"ĖE�,�"�Y$�$��,IdYȩ%�Q,�YY$�(�*IdIbK"ĖEI,�Y$�,�dR! !�! ! !�!�! !2*IdX�ȱ%�dK"�Y�! ! ! ! !A��%�%I*��,�H'x�9 K$YY"��"Y"��B%�,�K$T"Y"�D�%�H���;$��ED%�)!,�d��E�(��E�H���ED%�;�"rH���'%�bBY"�IʈrH���E$%�,,[X��H�HK$Y�H���ED'{�$t	bؒ���E�	d�A,�d	d�,�a	d�"�":�$��*;�',Q"YY�,�%H�d["���EH�bKbĄ�E�	d�$��V$�,�ȲHN��vYb�����"�`B��9$YȨ�,Ad["��E� $D�� �H�Y���"ء$�*JZ�D�dI%��($�V� �b�1 �0����IR � ��՟�z�d�����$�Q$�UD$ 
���O��������?�x��?Ο��O������/����� ���և�al�w����ӯ쟟��	�?�'�������I$=x� A�����d��?g$T���4��O�'���?�O�o��	>�K/��ӵd�����'�?��9?���I9��O�'��K��"D�,$���H� ��X���Ab
� YP,RD�Bĕ*%�$�%�RK�T�D�bK�%E�(*IRY"�ĕ$T���%��R%I(�%"Y�$�T,IR��*%I%�*T��,XRJ�YbJ�%*ĖT�Ĩ�KU�X�ʈ����DK`��I$���D�I	l!,��đ$�$%�D�$���U�%�I	e�%��"Ie�	e�"YPIe%J�J��*X"U�	e�b"RP�d�D�K ���T��b$�B�Y�%�
�@� �X���� ��%@�"�$D�A�X��R"�gg��������g�O��$HKBH�l�$��$I%�����I�������%�~��I�6I�������X@A�?��?�����	�?�?�O��K?���oK?ߩ������6O��I��������?��4��,l��'���y2v�Hz�X��) �` Y��B��6O�C��p����O��S'k��{��L�z�v_�?�����S�$���!���}O�����?�O��$�_��L߲9?�I��T���d���#��X@A��?�Y�>O�����?����2o��{����=zvI%�'�9'�O��/�3�'�y�>/P���{�ڲ||��8���$�?,���o����o���$��Y9'﬐�$�/�����O���N$����b��L������� � ���fO� �R     �       
�  �    ( (            �  7R��´kFv�T�5AI"�����(�J)@Ҩ�	P%*�� �"��*+]�*�N̨�m(�DA
T*��        @       (P       �@  
        (      �@rg�r�C�ON@� c�q�ɣ����Ͼ��0)\� �d�i��=��V���$#�   ꏛzh����>L�JR���� �zPRT�4}�E()s4��qI�4PQ����)Ar�iIR�Y�'YJR��e(/�U�)IS�>��� *���5U�eP�   <         {)JR���۔
x��K�(R�R���'E*��w�� y� �S#KՍN&����C�=g�3���� ���|��y�}U(�֭�UU�{�  �����{����� | y����v�{�>����c�@[x 	�Pd|@@���E������UZ���   �        xzS���Kzy����]<@��y����� ��4��6���v���n��|��P]p .�)f=�4<��P�(����  �/��|���{�hS�}����ؾ���gZ�wy�zq��|�Х}� ����Z�����b����s S�J��T��  �        ��7�C�{� �.�(� ؠ2n��v��t�>��G/O z�  �^�C�7B�'����  �}�}�;٧�� `42j@��8�o[N@� �q@R@z�9 �z��#J���
         �AK1������O!�UY�����P �(�rw|�P��@5C!�8 ��9��0}�I!B^ �������������5����9I��h. Q��`zy:=��@t9z����IRM� �)�L���   �{
zj�I � "{R�Ԣ�0�@"��LT�@ 4 I���l�QS�� �����W�_Յ� ��@��3� Aȍ5J�{o_���$�n�?�H@�p@$$?�	!I��	!I�P$�	#		�?�������̧���/_���o�,ۖ�x�#�+�9U��(Y�k�z{�Ҁ
?KV���;�iGm	`����s��c�lW%B��GZ�[���$eͻ���VI�Y3s��%��"�,{�s���p���i�t���f����d�g��C!w��w���+S�i>Ea�u;|�+]�;yW]��zq�����*��>٧��=�`�R�r�Ԛu�Ox��s�[i՜�G�t;ǽ���C�^�M�Y��YJF�}&\[�%�{�P�R���v���Fڰ�t�s�ރg!�7����mՈ�u^�s���Ra	��t35c�TP��
v[غ�ئ��\���h/f����D�-|������nlK4�Xp�2�6�G��n>��p�}k�6��9���N��pZ9�wp�%����*7�d1����i�jg��6(�h T�'S����'����5�85�vp�79+å�)̘�O��*�8��}+۶G�vΝn�����\k,��L����J���I�9����&����^<��B��Z�t��w��G�n� �s�g鰎'�;��h$�t��Q���.,���Ȃr8{���f��%����GT�D������Q�0j�h�ġu��+7ã�˗�n���!j�0巕�P��lk�2aㅁO�� ?����~�_Y4<�n�"�n>-+D.�mx�5����:ê���zX6�f��Z@Æ�7��]��,%���8���8��`�s��Cs��҉���^�<�sq��%���8���\�Yۚ�W�:�_-�WO�:;�����V����N�'-J)��p��F*�a�Z�7mG���E�[��Q��;������OF�y<b�;v��sN(zg�}�p��߃�gY� �Df������R�S-)E����p�6�$�!Q�=��0f�v��v�&v҃i�s�F���7����Q��xJF�;�ok��6�y���n�O<���aF@a >�d��b�?<Sl���J����9f]�s{�ǧ���OQ���;�q������m
�T����غ�8�/̹]\��7&���o4��zX��t�7��wiz��l��G��v�w(<�t�"��8�����NL��޼�R�n�)Ѥ����3w�i �q����=t�
�&��	�V<�w��tm(�{W�tkŹ���%cNs�mSNF�GN�0����)睗k���i����^هd�jG�W�u����9����S�b�K���s�n���#5�̾�4N�z��\dU� �Pہ®��Tˈ�sl�.�.mر)�ڎo>u��
Mkһp؞�L�^.����Ȥǎ
�裀�� W���CQf�-�N^�˙���σ乐����Zqtk��+ l�[Ðv�{x`<�}��	̛����PC�P�4�,�p��&��;{�qU<�|��*��-�z �8rp/)Þ�V9�t�&}u���[�`��ǧ�6[����giVe�9%�𤖶�d%j�6�{��F�L�9E����z���[x1}�z>4����y��7����Z�t1�0ZFE�r�������@<�>|D6_��o�"�>}�[�v�2���D&1V+�fl�鼮��6���������s�$��`Y{���qq�ss�N`Ja��Ϯ�k�wk�ݽrq'S�5���5�E�"�E9�ٝ�ͯ����C�"��fp��T��jb�]�����L"'��(2r�ua�%Ǒa��v��Q�sM�nuC�tqE ��:���Nq�淓9�q�,MEfqċѬ��r�W��q�dpc�1�͇I!luְ�-��]��w#��N��U
W+�9f�.���.G(=%+�s�h]���K$)~�y����2�!�f�������]�d�2�$f��FNH�m%\1!��:V����,��� ��tv"\����*�B5f��"A����o��R������E��LiǼ�N�j�)+[�����6-��X��*ND��6�'۾x���{�^N���U�S�F��,&Me��z��v�s��r�BRv�S�a�v��tmƍc�8Ξ��c�b�آ�|zwf�o�ë{'O�☌�Zu.L��*���;L[�6b�Ɂ�CO'��|�ct�P�	�����J �x[)�N���
�y\K�b��J]h�����*���wjAa�]X����hEuT���B��Y�+�ý���G��h0�Z����i����S�8-�o	i��9b��Y�%���;�'���!��+&��%�0�!N�����شgdU�D�I��ܖQ��a+�{�E����O)� c+��^n��Ք��)�Jw�N:p�����5�z�su!cp��ʜ"��]ϗn�90�)��%�غk8n����8��v�B7&Agݰ*hz��Z���i�i	�J����)�M���zb�������!D'�/�*2�bϔu�f���3�S���sOu��Z�[~�+gp{+d�}��ˢ6�������A���wr?Ky��-�l����3�I��$_8�dq�:t����4��1����&���>��q��Zԯ�wKIِ�7�8����&�;��k���vr��-�w`Q�� �aۮ�A���P]`)���)�msb�����٥����0�f�:�H��2��5��f[�9=:-��{0�J��d�]Ӗ���[�9���'s\R�}���f�Ǹi�v�I�C]�Y�]���Z���2}�msT�V5��E͛L�r��$���\P�5S�:ŢF�6����Qw��93��dC�ϢlZ��{8w�H����C�}�_�c�T԰vu�$ُ�wi؁�4���k����,n�gP�o&�g.Ǔ��҇K�I��קȱ��Θ��f��(����6E�/X�b4�t��g#�8y��q��˄����9՞��bf���m���d@B�	�{13�g7��γD7�ݎ/����жj+Szf��g\�vR�8��S;6�L�ۚ��wm��ٝi!Ȗ,�H�8\�T��0��Swrǡ0a�8��Λ�q�\�,zN�j�u��nqj�d�8�v��c��e})Tojޛ����.�_u�.nn彻��z���i�"\�&�{��׆6WH�[�׽�x�p����ͳ8c��7��_7�;8A���9�]05�sx�zFV-�{�3{�l�7k��n�9�}��1�ٷIī�N���"�;���MSe����eP�!�MƅZ�m��K�6�<��˹
�׹ d��\7/[��m��X+;|sw�}�r{�p�H�gw}ۇf��e
ĘF�s����sy���6�xM������-}�;A��dj�7��1�o��2�E����e�Ae���q�\Y���v��a�v��x(�z�Z�U���p�1}������7���T�:��F���-5^�&�x���ܭ�7@S{�]��Y�~|�yx�5����kN��bO�	ZJ��ocga7�s}��b�տ\ �U�2��ݴ-D��V���-�)�geݭ�bT��6s�N^ J�c79a�{Pvl��+�R��u�˼4<rH�]퇫l
���F��7kwR�� ��n�tٻ�k�FbΘu����s[݇Pv�sQ�F򙦩�-d-�Sp���7��ە�r0�x�L=[c5�z��>w�
d���#��р�f&�ߐ�o��M�·C[0D��s���L)n82�:5q��D���B!�C$�Ly���-(g^�=T��j�����I{�Y�$d��ܸ�z�u�wr����:�HȘOyi��8�E�ف�w�t<�vOо��$�ݝ�m��JDwX˧"��sqnu<b
8�	���Գgpz`H(�@7�kV�.^9�%T+���r�]��b	���+@t׽ר<�ѓŗY�ۓw���ᝡ)�LKol�p�a��v��~�w,�@�`����^s�3q�����u��z�Dn��#�N���NCz����F��7���|��zgB�::�k�|��K3�k+G\X(����Y7ID�����Udܜ寎<��9J�dk�Rc8�z�U���6˷qTC�/��E��q9�λһ���~ ��	�#8��ot�wzgr�q�ۀj�,�Cѫu�ڞ��4��`���m����{2�&i���ch���lL��1��v0�y�ۃL�,�zWlӦ�q�wD-A^j�g`��3y��*_0��u��YI��;��FtF�G��6,U��;���wXk�D�7I�8��?,Oso-/f��K6&��Vn.�F&qg[ؙ�t�/u��3L������{:��:=��s��8n�SM-��˜l����{sx���ik�Ɖh��[�8ga��of��.��c��]�����8��bw�&ͼuriumcX����ܺ������1a�6f��y��x��K�2 :�t*�Z/ ���\��[{�#1q �$��s}f�W�7���pQEC(#��v�Z���yb��v�����y]��"����� O�<Kv�G�����UǓB�U\�4���hzsb;I ��G;MDf�&�r^�J��l�c��2R���9��A� ^Ƹqu�lz{g$�*
=)[�
�&���a�-�Sn��n��)��԰���(s�l@���<��vL��6l�B�������^�@ȴ.��u�g(ъ��tc�sNh�Q��a�s�5�i�fu�4�v�{Fvw�;�e�÷V��jS��*S]인˼���&������se��6��-:�</N��٢����/�6�T9n��m�~��h=P9����g7���DC�x�a@w �f�����n\�m�sx�i�;��t�0M
����l�����e<w�[NM@�7� �UՉLX|{Od��}#p�H���>i��& �g��v+��;P���j�ԥoWt��X���j����Gu���켴u��l��v:�4Kc��r��B���Lr�dh��@!�i�gv���{�i���n]�3fZ%B�9��P��İc'Y�9��C�v��:�҇G��a�.iΪ=�u1�x�m�g=�#ʽ���B/����Fk��T��q$[9ӟ݃k�[d���:g'eW�7x1԰�GiRp{{q���SJ��T��70���[���,\-���ȆX���F�Ks�����<��$+lÐ:N��,=�֝�Ld)�^w͌��/,ᝣ& Q��͛��R����=M�)�ײ��G��+m߄r��:*	���C���vF��V� .�4u�z�m��{.t\�5��e�yr\�ͤ�tl"�sH��n��Ga�ǏTX�=Faz#c.��Ѐ���]�6�h��t�{l'.��WY�>ڱ-����@����`v����M��7N��\ᬶn��m�2$2_np�����Η���#&�}d��^��k�� �=B�kW	�����6�uێ�����=����U�lMx��^�ٛ�j#�wu���3K��8�`sxR�pz!��dz&�N�3��!��s�5��f�͗��ٺ���7�9u�:�U+&Y؉�#h&Qxan�n�܈Q��=�%��	�5��c�t�)�q �q7V���S^3H$����bn�]io�ӢEgvs�Y�`nM�,z��+���׍�1r�;�v�9����j�od�"�x]�>Y�7F�Ѷ��:ނ�[﷨�,�1cd&Y�zʳ�1�C�N��ݯ9����(:���?*�}��{��娓���û�FՈ-��k�,n�!��b��C��Q�]�/��|��G� �o0�[�-����N�Z���(Yx�+W5F2�+��`A�N�6L�6��%U�Ź7 |lW��V�2��H�~��ۜ&�Wr>3�Q+�����R�uo.��qh���SŜ�˰>���-�2v�!d�ňEݴn-�u4�TFZ�U��9Ż6dC{�g��q����4�wpt2�V�c���qiW�DxVW�����^*�yd��y:/9��I��,�k�XA��y�5�GJ>Zz��W�XƼ������$�,��m�*�/�R<&�����y��)����qrl��J�M��0�C^�:v���%=�su��oe%���]�]�b��N��!;�̝�Oc0���+���a�trX��}�#Ʀ���JY����ɝ�k�"_tAc��@;�f�ƴƋ�WT�zf�V��v�]%D�gU$
g�S�:�;tG�����LXy{]=�:;�Eu� BΝ�Q��a�q�'D0��pw�@H�i��U&�-;�<y,�c��l򔻆;����!<���٪!��!�]�&Y�����,_��5l��r��H�yw�w6�ڱ�m���ݺM������O"X��p<��N�tq8�����9r���tq��0=�"�si��vT�hv㣅p�8�ܔ�3����a�z��&��C��N2*�0�t���ww4�Bf������� H�(BI�D� ��EP�E��$�	$RI$*�P(@IH�V T���+ H�d�"� XJ�H�$��$�P! B�!Y"�@�(HT��	 
 �Ad)	 ��b� ��,��!RIE$�HY$
�I"��
d���T�+	%`I*I!)!"�����!!R �P$�d �	 ��a$XBT �XBR,� �) �BAd$�jH,�"�P� �BAd��HBJ���H�I$XAI$���HT��R 
 ��R*���B  BA`
@,�H�O���BC� �$��������:��ƭg9�q�Vn%���6��U���; ����.1��6ok��5v>��{b��t�d���0��S��,�H�h�O�����(�޷��p�/v��<^m�:ߺ�~#o��������eȱY ����F���wb�3DÞSk�թ5�U�O �Y8
8�����sL�_J�Pg�C>�\M�lU���M�{ش�,�i~�D�HԱ�:��h-�ݤ�Z-:K��Dۜd�M�	x�j�F�e�
E�M��zV~!����txb���H�B����ޒ	�.�Jq.��7��"����pO�a��fޘ�x{,��^�:��괮�x�Ӛ�J��u�t`�ۺ�i^8�|u`ҧ��Չ�:���`�ؽƁ�R�l݃�긌�{4�P�Zy�>�Nj�����.���d�!�7���'��;N]�v�Hz�F�{ژF���p'�b·�N��0���ujډ���-�si�wf��be�27�-�}P}7v�#��XI�u82�l�DN)m�A6�]��p�ֵ�n����c7 ^���ׯ�[�'�����h~=�6-X]�0���t��!��C�o5ԃ@�U7�vޏ�_m��۩�7�&�~�����٭�{�DN:"�Y���-[��>���f���@�����+t^��Fo=�^'�	��8U�l���}�+��6-Ldd��HƂ�Oě���R��Ȭz,�&�=v��\E��OM�;x79���{�)�/;�v� u[�rH�7v�T�0���Utp���Wi�g��;�$�������?#�g)k����ֻ�U�F\^;�x�G3�r�u�2��V�9�N��V�R���&�_�>�QC�/֣�q�gvv�s#��G+S���|�.Ej1�}���[���ic���Na��ӀPtkGXVw���}�{w:�� ��}�͕5@��wp3��p�2��'â�={H�MT{r<E��
��/��A
oHO-�0{s�ƋVu��[F�p_1i�}˽�󙻛ݤ4��O�~s��#~��%�W`B=U7Cs�{�������}�D�h�<^*z�nƑɜH���w<0��2�i��1t�� 5�5���9{J�r G�N��v��Fv����z(�>�N�+��k7�]���^w=�$�hr^�<M��ɭ���fY�'��h�(�œ|���<�/#W^5جmċ�{�8\ע;�=�d;��-�tUHW�(A���V��Nd�^���,קs�;�mOP�H|)E�Ṱ<���8��Ն��%q�l���gO��.�&����3�b��-�%�L4oT�{�z<y=`���_'��w�ܞ׶��S�xw]]�H7�����	�w�&�K��Y��.n��+ ;����{\c* �z|Nk�vD��dH� ���}W�����|�zkۦ�dKg��O&S|z2�f�)�4R`���u�/^١���!�/z�2����L����'�疢7YH�h��H��Rɲ�ʄ�'�Ow�,<���#���چo2��١�I�/�c.]Gډ>t[M�7O,z��N��`�����c�l��)%~
k�}dkٰj�=��	��w�R�1���k��Ҋ�9�Јs�wqp"7���'a�
t�3tU��4{�j�X~vbg�ѧ���;ڦ�0 �.�gGvِ���st�^��ܤ4����4羝.��Dܣ ��D�����/e�8A���pz�����C�$�,���dYg�����s��1���9���ˁ�&��Aɾ|	.�Ӣ�}kK<<�\ؼ���<g ަ��;2\n��V�5�+��=���t�h"�g��׳�3��r �Ǵ���`�J�]5g1f(}�ay�V1�+�%h�k�&�c��W��Fؽ� ��(���3�ۻ��@�+�Vg�-������H��wdԃ}���_��bu]K�f�1����\�x3v����d
f�M|��ݦ�_Z0g�)a\��Ȅ�"�P���}Z�>�i��#��y��y�k�P�]� ^�Y��H�ב��y���4���b��6��4�4����:dޔ�=7�)�~�h��縏��׭O<w[$r�W{�ָ�؎Z���0�����_e� gK��n�]܌Ь��y�x��$��*Χl��~�*x�^~^`�8@�ޛ��@ͺ5X9�S�8`:~�>x��e�RA6��������e̒����� Q���u���r/j����VI[sD'sg�oU�A����F���/�k BU���e�U���s���3���K�=�NI6��~Ϋ�ؤ�bЅ��8�l���h���(7�e���P{����`y�t�N��vl�
O���7��������|�yg�|y���
o�-�w2��ō�9e���u�z1���m��@���hB��h8��{H/q���.ɝ;{|���nh�P��Ҽ�$�[�裄�^���q�яg0|�}kW���+���y�7H�9p��n���3���;��mP�L��dҰ\ַ��׬�ή�w/o]�S�}�}���Kr��{�����``:��{t�4���qx�S,��y8�h��A����_,�`y��nr�r.5v�	�x�7�ݘ��;8_h�E��M����*�I��X˻�a��쾓��ǒ���9���f��rڴ������5�����@���n��q��U��IG�X:t���4n������_)$����O�3fQ��7<����;z1��Nv�&1�V=� ��}������|5�8�'N��i�&���un.�P�4H�u��b�t��!q#���
d�%Ǟ 8�µc㗰��;Ԏ�F%תqJ�io�ӧ ��޵�A�Vvgs���Y����$�+���Ш�C���}��d2����ւf��" ��L�;^�鯳i4�ђ�1*��������չO �&�����wA	�Ov��&���tWz�̽��F{�a&%�D/��s�9�E��)���g�{�&T��G�8��źf��x� ��6��z���{�}����vh��S���ک�9�g�2f�/�bh̹w�Ӥ^ӏ���])޺��9��#�ڲ�,�cZ�a�zC���f���yI�G�f���{X��B�wznM�g����MN�_�x�zo2H��}�KQw��B����W=�އ�QJ/�=�M�ၼ}~�xP}�|љ�<q�lN`��X�ħ�[�IT���A�Op�x�J\F�:��0{��&��ټj����`��뻚<�#3��$Y�z]�_����4y{ۍ�����{P>>�����"Ǜ��-�O���L��[e��H>���wO#�#�/Hhh���2ߎ�����m��{)��Ӡ���<�`��X�|y�\"��pv`��@��vxk�>�T��ri]��fU����g�Y�o����2t,e%�7Y��IѲ�����,����=S�a���d�po�=��>rc��g���%�<�M5�Y�9��%ő���5պ�jd۞�OE�cи�{GN*�	�>vOI�p�p{�<�^��Y��̠f�튇p��Ȼ�/��c�l���K���Wn�=&�(���ܷ�^����=vW��LսD���qp#̽�+����Ӏbsm�l��j,A�:�ux��|D�7�m�J�k5Ƙ�s��ȱ@���ݞw}�=��=�-�|�J��4�}�!(؟� �K�<��:.U���M��\��C�޾}�͢�;ҍ�L�ޙ_�Kޙ�D�7�3��*�Uɂ���}��۳�޶�N�+;��8��Y���������^�\Vu�m��|�xG�]n��붪q+۾\r>P�a!gt=���|��/r���t咅������sv���}u�w��DL�nw^�:��٨��a�Hĸ<�ֻ��ߪ��Z�b�n��<9��:�K�c3Y��N����<��5W�'9꽋���l[·U�i׸���l��I�wY��ݫ�w�x8}���whʶ@`������׼+�h}�;�3;��/����wk���b�"����W����
g��W�U�Ɇ�;�8:\��d�ݧ�^`��L����0On�·q�X}��Hq��y���l�����q͵����Sǽ����|1�B`���}k�Z	d�7t=x�s�]��KGk�,BLߧ��ɸ���ӳ:zל{Â�oq��b�F��V�.�(��Uڲ*K�>��"3Q%=�Cu�{ �t�$u��q���t{#�m]�Mz�w����?L�S\Vm�g��������>1��`��K���Ý�}j>�)���Ĺo���\D��N�q�������O��ܺÇ}2J'W��#�Wo�A�q���!+9>��3&��p%��K|�~�97}�,��g��2A�r�gZK7� �<~��.=�wY��V���G:xx�
>;�j���#��Ѭ�p��;9�\���/���ѓ�z�9˜'��;�y���6��������D���P�����I�~�ܥk[#���~���V��3ܻ���
�1h��)�t�_��'�������Y��8�z���c��%�(ޝ|�V�n�Er�p�����2�������ss��˺y�q���؃���y٣�"'���e�Kk���(K�n���W�=}�4K�_gp�ek`ɽ�.�����rc�Lܪ�)6�ݙgf���'�2�= WV�D�L�)T�z��?���on;f�SL�"ׁ��Q%�c@������v��dX^
�3��[9^��l����x����Ǫ�V�6����#�$M�
�J�B����k�����-�o����(��>]8�m��6�N�zLN��(I͙�<l�^L.�C�7�ی�/��]nQ'�J���B���C�M���^��pe{�{�r2%m�r�kZ�/6/29+��7/�./�|������7�j;]�4t�3oW<��Z�:{.���.�},`����<x-ao��������׹=�}ׯs�j�Ƹ�/�]£���+8���ʉ5|���������hUR4��r��gܚ$\����Z�fQ��,E;;�Q��W�7�2��p��YUL�ך��{ON����P�\(㆖�q�T2R�nt�� �٣��u`�dGv2^E0Yx��β���w9�9�cvv���k��,P��I�����W.P���5? 1yl����m�zè-�~�PgPt'�{�pu�;v�%;�#rI]�<��X}�V��񝌮t�{׳�ҷ�]:����r�1�Mجε^k�q�葓Fަo���p�w
�]~��]0�����c��6�ݑ�g���"���g��T��b�6�8y{H��L�rt�M�Z`b쉩?3�ўX�&�	ؕ����w�|]�#��8���z�={�v�2c�v���9 ͹�����z����+�`�o��zחb�ܷ1���M�i=ץ�%
P1Te��v�N�;z)�l��Bo��.��<!�x�V������������k�����9���,��w7�,𝯖���rwH��Ψ�^D�.;�����E!�דF�ob�r5å���Ogc6���э���{=�h��1�~(�B�h���h��!وL�:�z��o6Y��[�z{��[���(��:6�a�넓���۞C���Y���l��5��Y��gg���ޕ�~�GrI���k��Ixz�u�ǎ�{h�W5gwz�M(�U����	t���D�8-�3b�ZFL��o �VƷ6�a�F<���,�`�^&;�冀.�z��JL�u�Ϋ7����wso�� �e�'��tnz���˹W{�4X��Fo2���<��$����-���﷨�[����\и�q�m��p9�	�`m�g��m.��S���O8�{���g��.S������h~�̈��
ȷ�[��䎛�|R�T[#^�Fb^��zB�sk��RY�uS��+�s�h�*`��G�n�-m��,��L/��`էe�a��<���_�e^�x��y�@��g�uIb:>y�>�毟+�H{W���Ď7N<�o>��n�G�\׷�����v>)΀�1�I>�W'�d�¯�T{ >��_���v��Ӕ�k��9Q�y�}����(q�8��o�p*�6�.��N3ƒ|��:=�i��8h���٩��[ݢ�o�\'}y�X�m�h9�r�{�D���=��Ţ�|,V��Ap�=��Yd���l��ջA���W��M�}ݾ�7�]F���T}_w��C��}���~�G�bЦ��$b)�����}F�}��Gx���>�Oq�q�W����u@�x�#̵"@�ѳ��4C��s��pi)��<������-҆=ps��v�7���q�K�=jC�4��Com��=���$Y���uwר��`|{�}�F�=����r���;N�cȽ6��Ͻ2w��V{f97X˓Py�/����rPul��叹����^���\�t��Vʄ�ݬL���Һ�c��X*M�Č�sl���9n�|�4�hK���b>Ct9���ۅ��LY�n(�{h�{ET$ߑ�1�34C}R��}s��3��|��ǽ�ǽ������%��a�{%�Wp��a��^�����k4��4�3����=|�;����z��T{/M�c=�4���C˽6��8�w���˅R�z.��|R��p)�����9���{���{��?�H@�u$�v�n��b�BunF�7V�3�{bv�����3��h��v����rF7g9�v������]���6W�5�d��g�bm���9u��ݠ��Rq.hw!���+�[=m�W&.7+-�ml�Z���"{Z���w>�nyl��b�.%���m�g�G�0�s�;k�=;�ׇ-ԔrC�:	�����vi-vGL���9�������m�2=��fwV��76���kn�[���rNz6�s�V�7cl�%'�y���Ɨe�8W���5�60; c���ێ�n��[��d���4c���N�����r���x����۞�\Λ�}�0����v��d�vw���#=\����hLns��6��ݺ�l7d�y����v]k����N_O-�v��Ů8��y�:��d6�a�cH��:�X�U�����n{�=��w�v���v��n9^��vOn�p��,흝j�֎62!�=�
���:;��g����ܘ�����:�U�����u� �u��;�\ٳ�m�c�p�Bz[�۴���<���=C�S�sG%����x
I����gq�Nq�V�K�n8�8��<�؞���s��ǖm�^�n8�����Z���80�l�d�s�� ���([p˧t��������l�pr��aS��M�\�q"qT=��dw8#+�%�1\���ka�X�[V��rV�4p]����s�ݻɌ31��i�9��ve�;uI�+�&\ti�=TJ�=�{W��й����;[���7n��t�ܜ��#�6{��P=Y:�Ys��$1����w]�u��Y3:��m�
W6��Y�pZ��8qꚓ�Mۮ{6Tw"�ōn�tZۇ��dx�ũ��h؃����5�ݟ=d�2��ݻ]u�`�R]y�]qWO��;�����j���l/�^�U��;u�֋�P�0�u��v�9�%���ɕ5mls��5�[#.��l�[��n�]�l�Gom�pk��޲��l�/c��R;�w:9����s�7V�q����u�Wv���u>D�� �0l�8x��s��]�q^��xv�m�;Dt���r���m�B�su�CKR�r;+ҡl��ܜ�w=��g>݄��q��8���C�-�����^g��\��M��k�:�)�D�\�{=��ܲ&�k��B��S[e�WT�=
��k���N��*�#�r�/��f�u�.[�x�:�BZ�{O;���k��\��]n�w;�r�[�s����4\=�N�z��u7�v�t��$x����n��u9�f�s��ۺ���Ôڎ7j#�k�nɂx�ܡ�,T�qծ��-�kTX�{'m�{VY�e.��8�÷��D��,#�;O��D�V5��W���-�tu��':��`Nբ�1�֒'S���uһ7]ywX3K��#uש]7ۭ�[+�#�x���<���N�DW�����跦�����<��鷈�czM����F�9�"v����Q�6��V���k��c��f����ŕsэ�M���`S�:]*�\`�U��Ls���T�''+��Q��뷪���v�#�]Z��v'T��/Wm��j�[�=�^rvݍkq�kt���Gb�vy�r�����y�.�o�7J�aY��7��{�1���l2r%[���\�S������*b[h��V�'g���|�;c�u�ګ\�K�n6�[vΎ:,#���<�=�sѻF��tuq�<��շF�tc�v�`{`�11��on��k�W�S6�p=[�y�^�Y��=�����`�q��e�c^nC>�zx9�0��/q>�nϖ;����Z��c�k{6�7nI���[qá������v��n��۷�t`���`F�����q�]�F�r�m�ز������nWv�Nru=�<���mc�����N�.��hݫ�jɋ��k3&��mͻH���G]��nm뷡�4z��k�v9��\��l�NO�����y��WA[�QŪ������.�{Q�	���'K2n�Wj�m���q���q�ȣ���M�e�r�)`s�csjoWPm����/<��4�֮m+�;aaN�	��vk�8�Ml����/���s�u�{c���Om�g�ڏnЦ|�8����V��Qs�]Y�jۣ�����n�٢; ��:�ۄ�Q����8�����/7=���lX]��]�8�N�ݺ�ݺSr樼�L��ɛs!�su�x�k\�-*�zp�Y��J�m׮��v7n�^��nV䓭uƎ �e��"��:Ľ���t�ᔽ����hʉn@#��ݒ9�5�k��GH��J�1�:�Ӣ��g�8�nr��g�n��K�ϋ��p��b�˺}+�Y�L�������1G��p�DN�O��Q��z��no*�df�;��;�h�d������[�lg:;��mn7�8u�;����}+\�͸����c>f㣵ӆŉc�+k�N��q1�687e�����:��x�66���;k��r�:��^x�x7e�s�<��ac;����@m���]�kϜk�s��j��t�����\���ի��c�!��t��4�m��Z3���u�R�W��t:-��a�N���'��Gm�;lCq�����2m��C�����׍���;gq�+�.5n�D9S�:�p���<������c���jm�M��u���[�l�mӬG �j4�ɷ�*�:�\�c�n9m�+��<c��<-����g�5s�Ӯ�82]Z-�T�aJ۬t,����ޗ��v㬏V��s:�O���I<�$�b��{3��n'���Ω;.��ѷn#t��̓��p�+�l�1iۛ�{`�u�vo<s�sƑq��5��v�����c�كu�u��6�m�O�y�@�n&�6Mkiū��7cL`�G�m ��g��&S���CѶ,c�O.��<���X���_V�ݱ�&�OJv�\�m��uq��ٮ�w0u�8��y[����N�x�w%���VUu����1�¸ɰ�Km����Ka��Gg"�����竇p�0���J�Äz�B����pj�X[F�q^I�r��1�n}+k�X�G8�X�&qs�d��N����J�L�H�p��oGnv�YH��OT�;�x�K�Q:�q-����t��^���Mc[�ؓ�+ܝ)˽X�9�m�=��sn�h�;�n��wm�nrM�JD�v!u�{<\��u�k��ZFMc��l]m�ܽ[n�Ҷ���	ۗ�[d�+x.UY y���D[��r�YN��Fɺ]��Ub����j'l΄��;t�`C���t�ҹ��q>FG�ph=��nxԮ;rz.{C���X��<��;��.����qW�]$v���ua�]5�<�s���p����ݎ�QÐ�(���9뮎���nݛ=��]97p���/Ki�bW�c���6�`��i�R��ŷCڷ�t�ܷ��=nh�z/+��\�ҐJݝe�ܥ��WG=m���t�
U��r݋/\�:����97@�b�n��9e��-�d/d�5��P]�m��n2v���η=�u�ګ�	�67�ۮ�����<�������k����{��u������%�)qF▹�/��^�'m�{sX̼/�vl�p���sm��1���Џ-ȯ=m���;��q/c�m�y�Y�u�۷J����磲Wk���띋˝Â^�ج��rl���z���n1v��v[Sb⺞��&��w'<!�h�X���w]��s�Y�q���\��}���,�u�6�����wn6�8�5Q����:����ی���y��q���i]�qs�ƷOu�4ۜ�6u���S�z�q7C���.��n��ãI�⮶�b.j�J�t=��e�͆d�]��<@y�N*:w;���vM�U��W@���RG�>^�z|][�v��[���.�p�@mm;��m�'��xgc.`�c8����a���lq��vy���2�t�h��.n8��%9|��e����,҄Q�5�]^�;e��I�n[X��I�LD��/s��۱�`�g�UT%��,%Pvҏ�0qX�!�q���M��nA��8�=�Z�T���M�buJX;u�mv�݈q�g�ycH�7g�@�����x�[�W����8���vMu�{Ut��_6oC�=t�J-�6��qL�v^�I[nd�=�h'3�m�ݹf�p'<���d�6�m��[�e�����^��F_nee=���r۷<�ҽ�⫶0p���p�x�S��,�<V�m�,�=\�#gv�����eֵ׃��A����Ɍ��/9��;���qq��檫�$�Y�ي A��t�n9��.zt��@z�:�h��+G	�s� ͗s��e��8'�xܬ����ۮ�|Ӻ�E��;x�n���=�<<v�����,�k�ˮ6��x���z����.= �!�������h�<�u�r\k/m�ֳ��3�zK��U=���J/6��
✱�Y
;q̒�Ll��ˣ�Yٙʵ�G��6�8�&��vM�����T�]	m��c�d���ݞ�����������o=-�aFh8��m�wU��.�G[V֐�������(*Q��G]��c�2��ռ�=�εj�f2���Z�.g�)��n���;����u܍�ǧ�&�<z��ꋜUћsqۇ����s]�����A�c�c�`xi���v6��n���M���"ҽf{�3p��c�I���\شW>�8웬��aos�l�WV�E�/m�mm�{>k;�@�b
�uۗ�b�<Y�g���N���w���3o��/]cOK����u�Z���T�M�v�:�mjg�*�5TQU�V���TQU�9�B�݆�n���� nq�VQ��h���b[��V���[5�iR�l.�Ҫ���Gl&h�qUnJ�TJ4��ҥ��)n�B�ZZ�;���B�p��aU��\�r4kM�S;%�R��LTv�P�1�0���@P���.�\���i����m]��d�GE��u2kB�X�v+u.��c2ݶm�K���̶�^��t�
�v�����VҬm����S`�P@j6Զ�+Z����(U��kM�lQԶ�Mn�UJ���ij0�K���UsGYsn�Ū-��bƭj�ѭW;���]������6���a�����]Qh��ȋ���ڊֹ�����Ԋ֊uu�p�UU�թZ]K�K��0ɵMmQ�֨�j�(�1��vɄeťڥ�(��ֳ&E.�[J1-����݄���������H�c�=]m��e����V[zlU1v�-�QTm����6��e��b�Z�P�ZR��DL��b7�u�+�V�K-��:�k��au��*(ʴ��uȎ��R�N� ���^���u�]7���\���Ջf�.��hz3�$�A&ݵۋt;���7:	��]�:��bs=���h
�œgv��a�\�\:]�S�a;z�m�p�=����
r�!7�W;�xx�p;o/a�>��<f�s�u���B�l;r�9��h��l�v2Y��s�]n����6u�Ӹ���{n܇����@>C���Xpx�'����N�۵�uy�W��9�)�8㳸��;	۝�VV�]���\�Ӝ���:5�=í���Aظ�%V燎T�΂٘����ڙq�;��΋��n�����]���//u�����7fN���m\f�y[�6,���t���ܥs�5�˶��C㶫l�O���!�Q���rΊ�ժ��p��w-�����O�3ڞ}6}��n�.
�^ӓl_�{�����8�n�����\�y�dml�d�ĮOn|��v��e���5��^|;�ܽ�8^�v���c����c9�_����x��h�-O&�S��۲�݊�Ź{=N:�zt��-��hm�^��]��^���n&��Ǻz$ܛ���cM&��v:�����q{����M��ۉ�7Wg[kv�mu�����\���8���a����-���'�l�<X�Se��{-y��Y�vNwr�y��=U�ڣ�ɸ�ù�5۴�+9�ly�㝻6�Qޣ��-��/	��^��)��In�9#M=��\sm��V��{r�����:���\xˈ�]4�up�	�t�,1kl�GTn˓��Fk���lP�^�iM9�F�U�ҺE�m���q�;xg�����3�=u�6��N/�8��V�&�{L��<rtl�Ł�-p|�_�~v��n�e룎'�t�3�6��r�㊻=�-�9�ⷵڇm���Y�s.��n;�ɧ6��F�9�����E��p�s��n���_(��%�ppv�$���,��`�l�ĩEM�w��z뵞���k�EQ�K���\:�u6����]M.�G%�G1�����DA�<���@��3��G��>OG�p��Q�v�9ϗ���g�QqT�Wk[�]�k�Zb�\��d�J�Z5�;#�e[��E�&�7L]TSj��ۄK���9ҕ��r5��UTk��[vv�.�2&��e��h����.�mک����6DLD���p�N%�?]�$�7�|H$��1&6��vh=P.ki�ʯAu���m����,�9]�H!���LR�]s�@�	.���H7���(WT��ܮ'NۿD&�F�H*�� r���MvӐI {�A�>�S:���]g9$M�S�Hٽ
I�[H�م>;�٪n��C�'�>�`O����O�w:�����YυݢA۽r	�Q�Q�Z$�U�f���@7{�B����l�Z��9�n�H$]������Y}��F��p�
-4K��(��Gn�y��
���|��vV񮻗�a^m����Ϯ*�i��6¬���N�S�I$_nuP��A��&<q͹ �Φ'���$�8J)*��=�6�;n��[���{:x�y�u{�r|�^WD��=��7O^�Oa��?^Rj�z��a�7Y�w{�-�b����5��3y��|pL��}�A�ͩ ��Ϊ$�hu����df���'5ܗ�	(`��b���$�w�:hF�:��������*q�>Wu9H���6$���7 �fp��aRyf��%�� ��ngUu|�*0�-5�$�N�&�`RL7Aa�HGs�g�/��U��L��f���U>��ڠO�>.�����W\�Ib�W/����ʃ�Rq`���$+n��ݼvy�W��a7+���~����8%	i8PK{�ki�$���I%��b�#M�����-).^����Ϊ'�r�i�M6ڄے�m�$�#zy>��ER� �O�����Aw|���<��c�v��ӟ:�[n$��)�b����$���|I ��ݛm���yX���p�-{o�8��s���R�B1��\:/p�qжz����)ȥ%�B�7�:�������5�Y��5{�5�Hw|䝷r_�$��"�C:��/|	=Oz�|H��I��hqԆ�^�WN�%��Ux�4O$Y�e�!����ē�k:ؗˢ#n䲺8x�u��$<�rO���rz��yk���@�)���vHLip"�.nݳ\c���6�W[mRg��ܬ��������p�0�8�^ez���1���W1'u�i���:2f�n9$f9�	CN�Q��r	=�o����W`P ���>>���t�d�G��;m^��i�M6�)���X�N>� �A�麻��k�_d�H/���A�����U�n$��,�b��m�9�g�����2�I>��"|I Wnup�a�J�U�}���(��8�߮9v=�ۢ�%,��_jt�&�N�j�i�����s�'7�5{u^�q��f�2��z��s'6Ɉ���%�[��P)$��D��c3�Y�����ɜ���U�;{�w���I�z� �V�uQ��J�ZPtBۣ��Dy&F��2�9ər���X8���2�\�<���n9��Ͽ��H�H�s�vc�H"�u�$	��T�=�&T���߁��ψ ��9:�Bd�p���$��%n��j��׀�M�� ��Ρ@�Y{�"7;�3^�1�(bm��nh�N��n�:����t8ܘ�ku�$��N��ΑE���	�ᲓjAs���Vi��B�IKi�$�7{6�ĂK��j�n���@�Z�s�r���
p�,�bhx�e��$�ێ|`���mH��A�j��%��h������4q�W�mm)���&t�V6c\�.�7㞺�!�z�8�\3ˠ�8��p,�.��]AE��p	"'EKb-���R�!$4"
i�A���u���Z�lr��ٻW h'�qk��U��[������k�I`:�L\t��P�[$Iq�f�b���Y�q����s���zL��Z6�懪��˹��Fuv���hY���267`�ӹ-�X
�G\ϫ��i5��[vlm���i&��v<;�Lkn{s�]ų��at^�v5�;T���O5ȼ$�Am7.�V�}[5��nzs�u�`�|�v�|л��xҋXu������I"��$�������wns%]�V��[�4�_U� ����*���a���P9َI=�T�]+��b'	��٠A��NeuQ��\�����9^��)�6(��t�����I8�J{.+��O��6����$�y'�P�2�-�Q�\���U���� �(쫚�A}|�A���h\�%��E>ڡ^-v8��M�4�R��$�.�&���^7�H�λ���� ���cr�LM�W�d�����A�4��YU:Ӷ�<��;���fͮ���'sӻ"�~~~���F�u�����5׵D�n�>�kzD��Cx����g2���Iu��mͩ0T()�
0���9��F*�}�fR��-�*�ǖ`}�KcA=r�+5=����n5�;����b�l������~�V��}��J��´��]����> 9|�H6���	h��OnG��]f�ċ0�d�f��+qϏ�g9>��f�*���t	.���A���z"I��8�T������[���e�$���D�A"���f.��`��	&i����J�Za�[�]k�|O���P�v(��N�0뜓�A���^��W�cf��/�#�D��Y�R�����E77F�%�ᰎ-ۧr�ܝ�V��������6Xm4��[��-�$�o�zh���o�@8���A��v��
e�e��'�H��w���*���\�Ēif�$��f��W� �dwd�ҫ�}��^�YT��	(L@PɅ'�q���oP��Ou�@���&�d\��GTS���.e�z�i}^��w�d�,]��z�����;�圩{���m�lu��p?W
����K�=f�cQ���a��o�_9 �FV�U[W � �40\M9���Z���|�OU��4��s�K���3[�,�%�Ϋ��{�Z�.(�Q>;��B�$S�rc:�\ѻ��"椂@���$���$i�9�.yA�s�uf�Oq� ƈ,��i��$m�s��I� �7��.չ��s�s]����T�W�|��ԥCp�l��5:��n�v���A����	���2���i�$]v�P'�+�&I��M�&�� ��'"�#��A#+sj�A�s�H5�Tf"��6��=Yvڅ	��\1U�3Y�DA�_�\��T��\�!kl` ��͡@�.�$���%(ICf�L!���t�rY{	#.�����H"��H���+��Br�Vd�4p��r�'*��^[��Ǹ�X5����g>BhKF*���ǀ�Z;f�7
nH�Ȳ����A��)of��Mݛ)ɣs�G�m�m(~��8��T�$*W�ʸHd]��jtQ�ob�d��)��'� �y�]�|f]\+��a�J8��D���vz�Ѷ���Ch
���;֧���p���s�*��̃�MJ��T���v��Ä��mZI}	FOu�x��I��������x� �A����t��&�0�-�xˮr	-tU���9Q7�@�|i^9������6��3Vjȉ3
�iK���$�nnAɭr	$]��S���NNCB���I���A����m[��[PYpĆ���D�8����ܒ�}��ZQ������T�#~Ic�r	=JKP�i��S���ݮ�G����\��7�lH$��`Nu�U>����l�}�����V`�Ob�mNL�^ܬي�n�4F�1Z�M�Q��º<|�I����G)^�'�Oq�N����N�n�D6�,c��c���jNxqn��NY�U"�n�=nP6E�oM�}w%���͗nچ��O���y�͸��u�w-��v�ю�o[���,b����m���7u׮�K�ٶ�y:��{qA�춸��xJ���v��s�\!��S�p����k�o�\������cՐ���c��\�5p��]�ۑ�����W'��>jŕn�f�c=;�kv0=�Fsn�k��#1��c٣`�ǉiÂ�)��H����&����9�M,�$}���@�(ӕ�&<$���&:�D�Bl��`8��vM����q�mt���4�kH�	��^闢�K���Kw}C��l��9|�E�gU�N�\a��n���$���A���@�]���i&p�s�Z�}ysQ��х,���%ψ>$wnmP$|iv��b֋��l��$f��zu��	�h�y ��ڢ�v�5|۶q�����K���|77:��iv�<��ƧҺ(#��x�:�\&����F�Gם�8��͋�t�gu�p�}��$�qC��$����(�K��9�*l�~K��۴�ٹ��	|��I�ELRB��~쨸VS��~�9��>h�v�#��r^+KR����*���̉��۫8���xM���%���پGj�#��N�}l�,�u��cSlo� ��Ϊ��iv�$�0����K�i����	�6Q��s	"�k�I�K.0�չ7r$F^��M.�>'�w�PSE�S��P3S��,l\eP!wNP��	����I�u}�2N�y-9P$[�p��u$�$�M&���Z�A�x�☫#�$OL�P$)_9>�|���N������y.�X6�<�d�w�sn��96�52�s��X��6��������(T��]�������DS�Wa��o���lwM��b�l�a'	$����>��Ke$�"�����yϡ$壅뽔�g>�� =�V	��nw^�]���՛ ��"�)!Q-�/{j�� �>���I}�+q;+ʹG.�ĕ�$�"�Kˏvʟ�7t;����|�{�7���-c~��)`��}��0����l��0�>�uY�L}��6��x=�}��	ý�O�Ϧ>ߎ�t<��������|�µ�ݟ{������O��=���r�8d�<3�w,H���>��,F��)ޅYω�MN9��y8�o-�7��-}�6ٹ�U$���ث�uM�N�.�f�3�v`���woG]�+�ѡU�Q�e6����i�ju*4H/.w��?�5L>�4ST��=}\�]�w�^Χ&yn<�ǹ:�@^1{�;���C�@�v��H��]������WV����dk���gUq@ʊ��I���Uy/CІ��v�ˮ��9E�z.�[�W��ia�Y=w�K3y$�Q[�v����X=�K��-l���;����!��{�.n%� OyXV���@y�;B��g�#����i�D�w�=4��W��\����,��Ʀi�ɐ/���x���3�O��I��sە��$��Q_O��<�xP����o=�lӹ2y߫�<A:U{��;�k��^>��{^^c��#ǘ��_ݼ��r({��tγ���W�jZ����f���!�r�7ŸÝ�=	��'??f^\
�DZ��]��&z�uv�sv�/�<bN�Ϸ�)�,�6���<�����4ˎ�����ev���KSt���~�p`����v�3VB�,9wi�7�q�q}��s?&@^��^q�`�ۘ�^�U:H��>�mn%���Z�M�no��
�U�V.�Q,X��͋pa�E3��sM[-�����ʡj��b6нk�ik*�J�=9��U�����qeE�]kJ�Q�+cKiJ�[QsVժ�h��mj6���eڬu5��7�e�u��sQL��)A�j[mizK\��-��ѭ�Ֆ��9�֩��+[�SU*ڋ,��+�T�%�*�EbX��mJ�*45�aU�kZ6��-iiTX"4�\�F"�Q����*�)�DFն-m�cJƚ����K[E��52U�keE��Z겕�/T�RīK+�5��FQ�cb�֍l�,�(��5�Q�Q\�m.�Z�\��j[q��-�X�B�T��رm.EE*���M*t*�Q�t��Ƃ/Z�l��cmJ��������m�f[�B��h�u����V��nԭm��m-R�\�Qn�8s\��b�Q(����YQ��Զ��ҴHʈ�V�KZ"�1�m]k�G�2kkk�cPZխ���l�VҠ�ѥ�4V-5���9[l�ڌ\�(��.�"�5�-��ִE,k�n4V����WW�J}�q$�>����͉�I��	@�����˙�C*Tթ���ӪI%X	�u7�k]_��n�|�`Z�A�EaX��A������ٝO�{�4S۸J�{�jc& ���$��ϩ��ogSv�N}펚z�L9�a �Tԭ��E�絷n������<�a1�{v��n��ͷe[6-�����J�J�>��by� kʴ����l<���ۗi��^��@�9ɘO�j��-4����@s}Y�����3{��޴�n�x >|��p�u6���N��Ȥ<���[�@��ը,���-�{�f;:�0�&}��ә�U{� 7=�� 7���>+��AJ��W�ݙ��y3=3� -�S��@m/��{��OT*J�I榿��$��[�B.�G�ẙ����x���Z����Z�m��_pv��,���E�$�ug*b��v/P=+4���uY�'b�EJ-$[π�=||��(���g�ȲD!��-�I�!.���gI<O�;���x�fg$���DGOH�=D������#g��0�?������h ���ߺ�i��T*��z:C�J�������κ�u�6��Ʈ�u�/KR�[�Va�����ny��Q 󪇋�k��Y���w����ul��C�G!����p<�1�d�j��߾��x�:3$ɓ$ɶ�ϨI�(��>��o}��DH�G����fdυ�/��"B<;7��-%B�_>��V��v���u���v�����$a���@G�<�ˀ�,�u��~C�����C�*J�IP�<>���x��<�IP�1��n}É:B��4|��?a,ʄ�ފ�����g��2L��a��n�/[^���<L����u�����2�%���wI��y��ٟ?��	]�� A?!�Ʉ2��������d30̆IR�����	�3{�w��]m�m�[@�YO������ }���__��~I��2M�fw��]�3ę��2d�2m��=��N��+;�H��G;>��G��ӃV��#�"���x���2ۿ�5���F�^��$�{��p�~C�fh̆IP��>�}d@��+^K���$@�0�s��0��fr%K���$�2J�̓8f��������<�rM�b������9��%.������ؽ�s�[m�g�\�}w��Q�L�*�,�ȓ#���,�3����~���(�9��$���E�k��)Ӳ�֜S�[T��B�r\#�$!���رn��2Yv���n�y�]lq���-�|��sv烏<M۳5���8{n�l�U������T�[5/7%�ݞ�t2ԙ�ͱZ��%��2�9��������]g5��`N�on�\���խ�;�������v��Mѳ�s�^�F-ŷm��2wM���V��k�Su�fɍv&X��v�$xf���ck�+������߽����'_$�
�����|��3�d45&K��9�'�*%B�����!SȆC%���������;C�w�{���3���d2J��s�!�q�O?���wY�^�����yy��]�2� "=#�x�鏔��)�����^{���?��L��S&I�I��vq'I�L�3I������!�� A�M�2�q���
��̐9%B�_=��V�z6�������v�!�}���ĝ!RT*J�}����;B��d2J�a���<�n�~���C���f�d�/��p�N�(d�
�������x�	�dǿ���v��֢P�#̋!�g�'��R���=���!RT������8�ԙ�C;��x�IP���C3	��~� Y�ӊ���+���@��>D@@�B�7"HD��]5P�M6�-���C�*��s��|C$چI�>�oL� ���15�]S�<����DL����8��쉒fg$��}������y�2Rd6,7�~��Cĕ
��K�S���D[.ip&P3���0�Y{&�����C��rGm�q�������ϣQ�z�C�?'�7�߸q;C�d�
�Fd3���y��x�IP�h&C>	}��R@��e��{=kn��>�@D��no��ĝ!RT*J�������<O�2c�~�ǧm��n���gI<O0����q�>$�T��?~����_s�)�f�����y�ݩ ����ʌ�%���R�A��Cb͘�u8n�"`��-�ۉ��+|������Sߝ��=K�y�ßRq��!�T+��}�p�
��S��fa7�~��C�=#�@�c�U(#�k���ƶdJ�q�~�s��z�Z�tttn��x���3�~{���d�j%B��~��8�i+�3$Ʉ�2|y��?��ۍE��>G�B#��G���ٟ�ԙ�L��߿}�!���!�ϻ�ջ^��v�uz���;O2o��!J�ޜzOU>G����������x�C&C!��f߿~��!�J�a��*_w>�ė��co'���������$�f{�Ϲ�x�	�d����uy֥�k�ô�!X_�y�8���L�9&C�%���w)8�g���^�J���� |:��x�O�d���}��q��̆IP�a2k�>��;�3���q��Tc�kP�JP� />���F{���-�h��XZ��:�q
�a������2�t��֭��IP�����ψd�P�*������g�2d�2$�~�$zH�Dy;�]�O����������x���!t��m,7����C���!��=+��OH�����2^}"H��wo��ɞ���!����y��3�22���}���f�d����}É8@�=��#��N��0�7ӑ'}�g*f'�d�7���Mף��t��vt��+�s�v��RT?MI�߹�wI�Rd2J�YO��o����~׳�?L�s��{ �3(����j�
�J�f�¦�|�����ίMn��˽-�m�ks.��P�	������s�~�}���L�C3D߿�{�!�<fC3Fd2J��ϸqӴ3������������w��%B���dǛW'���;���P"cP�/�?~� �g�2h&I�M�罜I��L�3G$���������:/������ Fz��ۙ Q������q	C�I�Z� Q%K~��O����2�fC?���8x���{����������*���<��!��a��d����>�ĝ�C$�T�љ����x�&I��yH��>�t��;���-$ˀ�ȫ�!�q62Kg\=C;v�Ml�d�v��������W�Z׭oGǉ:O�f�?}�!�J�#�d0jL���8��^�2%B���~�x�O�d�[�߽�Hx�����v���*&M~���(D|��Ta��h��&*���!�߾���*'?g��S��~�_��>���g3$ɓ$ɦ����ĜN�$��I�����������@�Ȁ�*k#9b�s�7��<C��0�gn�}���L�z�!�y2k���I�+;fC32��������*����g�ߺ��οo�����C���2J�I�M�~�vr�I\̓!_�����i�d�=�N(a��ȈC#�E��_}�2|l�_�_���~g�$�cRd�n�p�e'�Rd3������x�IP�*�&�߽����xs˹Ǐ[��]�y��"����s k`U�"J6r]��R����{+:V	J�B�\6J�j�?j�}Mp�n�ս:�甼�ߧ���T0�7{��qӈfώy�޳ֽt�g��$�W���p?��2M�d�P�/��{�!�Jߗ����������O�2L��y��t�IY�9&f�߿��x���!pRd6�{�!�J�}���ntuH�~��?����z�m黵�&nȻ��]��ƻ6S�ݹ��{u¹n:�~���9�6�o��������É:B��T�
�Ͽs��x�IP�*������ #�w�\�ݲ�<���P�6D�vr�I\̓:3?��������&M��������׭oGg�:O"f�>��g��L�9&C�>^�u�;K���vRq�L�s�w������<C!�!���M��{�!�<����@D﷢8��/���(���D�,�!�c�=�v޷]n������8��_߾����d�
�j�����<O"���G�D8�����/�I�D�34rL��w��<C�I���!�a���y�<IP������)��]x2�~ "�6D���n8���u���z�Fd332��s��<C!�!��d3����v����"��A���I��V����Щ+�̓8f{��9�*y��}�]�zm뤴볤�'�f�>��3�ę�rL���%���t���^��r��?����C>�}�9Щ���a|�߹�;IP�*&�}R$�@� #�jF���!v*Q�s�h�Gxi�%�=5��1�1�~c4�^����XF�(6���(�h�`��]Y�qL���SQ�� �{	/Nd�ӟ������M̀���t��d.�nvw�;���cA���#h��y�Z�ɻ�χ�zz��*+�:��s:E,vv��箰�6�y�e��zf����;��.�]գt���EV��3���ݏ7�ێ��=����\78�q�^��X���խ�n�&�����s���s��ok'm���=Q������pz�b@�u�o�;�r�탡gNʜh�za6��s=���'h2�[�4gX����x��	緤������][N�黼a�C=����;B���2M�f�߽��L�fI��*i����8���G�yUy�0�#�(�}�υ�,(H])2��߾���a��/w��s�uz��u��!�yɻ�p�v!$|�� #��>~�q!d�o��'{��Fx�C&C!������s�v��RT*O57���q'HT��<�K����UE\97{�V=���0��"����"QH�<ȰB>
�:d���
����~��Ý�q��J��D\�k���ڮw蹘7�S�@���L�C0�{�8�l��̆IR����8�a߿��o[��]bpLM$�X(��o�2�2*��H����'F��cP�/���8��gFd�0�&Lm����$�v&I���3w���<C�|w��^?����ma����8���2�xw��ٯ]1��p������'q��*�fC?���8x��^�^'�߷��
��2��y���x9�9�jk���q'gt2J�d����}�9`�G��?W�%]t�I�		���>yK��nօ�s;��@5ug�)���m��T~}��ޭwU귮�S|t���0����q��L���2[����r��6)2��s��v�O�d����u�_d;��$	>����Ϭ����*[���8�i�����ގ��=u��wP�%B����|C$Ơ"=�]�6���H�d8�}C鹓�ƍm��[�:�՗�(9�.Vv0��Ü�D��2G�^�ފÃZ�M�tba�.�F�y�[9�o�<=��G�>��d�3ę
��$�o_��$�v&I���3A�����<C�Rd.��n]֎�ݞT{��=�� Q������unwN�W^��܇hv�d��>���C�30̆f�2��~��!���f˺��� Q%B��T������vwC$��2L�g�>�����L�&�������(Yd_�G�W����n��5�����}�+<�I�Ƥ�o]�p�t���I��*߻�����<C!� D|"��H}�}9_w�{H}`�!�T����ĜB���������u�N�Uo~!�C?~��p<��d�
�J G�/~�`���;Xd��Ϲ�Zs���t���&I�}���$�w$�T��s�~��!��!RT.������ A�iɿ�2���BJB'�v=;�kv�s���Y�Yi�-<pv;����v��!��y�w��ϊ%���G�B�ϸq;C�332�3!��?{�<C$�T�
�o>�����<r���]�d�i�P<�D���@�AA�&s3���s��<L�&��~�կ]U��usMْx�f�>��3���3
#Ȁ�-C�S�d!��DCH��� mI��*�����;B����Y��{���3�d332�����|�w�zT��9ÈD��O���[z:׭��m���!�;��r�Ry�d��3�߾��%|��2%MS[���1:���w�����U}�p�m�c��rdi���n��:�'E�T��熄��;�9���.����{�N�����q'��&f��d+���v�IP�*�a������0�g^���V�t�����n����o�yÉ�;��=�g@$G���|��}�"���L�C&C0������<a��@�#�@Q��#�v�n���x��@̓!_����!�x�&M����7/{��Vގ�t�&a����8�i+<rL�ԙ-�ϸs�I���ߵ��}������!���}�9Щ���a|���8�i*�2%K}��8�bv�a����<��w��ó��v�孴k��p��֪9ՅǯX͸��V�t����A��æm6�i�1�@���D~�����I�C$�P�/����|g�3��d�2L�oy�gq;$ϳ��}	1q�G���n�3�dP<���!�a�����>2�xw�������;�t���5���N��|��?����r��gy�y�$�[�8x��a2&C0����x��r�r%K}��8���$|��7x��f�R�b㽆7���3�"<��릠��ۄPR�,�|�}��g��L��5&K~�9�ID�yG���۱G���*��RT*z!��ɼ��y�<g�2�3!��2k�>��;����{:!�e�YI8Fe��n���c�U
^�2�r�A�(߷&O��$�fI�&I���{É8�IY�rL�y���;C���l�_�s����}�;��wi�G_Rz�;ˎl ��zY�+��B���t�ޞ���{۞��XO��@m�j�;�_/z��{����|N!ԙ��y����!��0�e����[�m�ۭ�܇hv����<���C�332�fC>����<��[=�q��2�7^��|C�9�C$ښ���8���d��2L����r���d����?'!󺬪�S<����Dk��r^ȯh�6��<s��ڻv�ůX�p�/_?�w�g�������'I�f�?�s��|I���d6��o�{Ý�N��Rd3�d3���}�p�
�!������K��a���&���s�x�#2%B��o����(D|��0�i�CN	����D{w�,�� A�Uۻ8��H�f���|g�3��dɒd�~���$�w$�T�������C�<ԙ�&Cu���}�5�p�|��C��a�Ά����Mo]1�wp������'`�hfa��̆y����<C!�!��d3}����7���<��9y�>���_�q�*���2L����$�%s2L�g��~�!�x�&!��ۂ��p� �"=dY�*��d�o_Ds�w��x�Q��""���6)2�2��������C!�_����C�n}���y���V��oӴ:gL�d4&���!^"��-���`�8p�u>R￿��v�I��2M�f����#���{��.��{ďIB#Ȉ�w�$�v�&frL�9����x���!qI��/����!���X>��w�M�
 ��b#R�MzF����3�6�~A�cv�oO9��+nTr2�Z�����J5o��F<}��s=�����v�z5���=L�	��t�����p�C^oE���~��t��.[�f�љ2��}3}�cM-�Q|)�Μwd���Թ�'���͟,osFCz�͌\��?O�
�J� �v����&9|<�k�;"ڼ3��y�:���td��^��t��c�[+x6ߜ��]��;�����U>�y�t�d�=�v�𓵴a�g~��)�[�{���v=].>)���Eӑ:�mef�G�H=7w�^ǽ8�׈�����@&)ry����߆*����˼tNN篧%Ȩ�:6*a7U'tL�2�u��T���h�b�p�X !�.�F��B�,ӆ�~n���C:�Щ�R�$�P��W���8g]�X��)=�*���^M��m|�v[ c*�W�|6b;���#w5������2��|��1{:gn��b�q�Y1u�X|��]�u
��\b��i$�����n�7��c�s�^�S1�	>���>�-�_l6���x�Gl�np�V[Z�o�4'��ۯ�f�.t����'�=�x��w�����+b�s��!�
r���k�|��C�;|2�orx|,�ܽޙ�Fx{�@�����}�(5��\zd����j� �&%��:�������ٛH6�3\��v�i������\i���D�.Sh�~���Y.Nh�u�s�v;�ķ Ш�V������s���IkgNTb�:ڥ[A[Z��`�խk���cm�Ym���R��T�j��ӫ�mQH�e�ږآ-��%r���Ph*[Q���khP���f��
�R��,��5�ӵ)mUZĢ2��U��Q���25�	����K��J+R�Rƨ��K�ږ��(5*Z����u�.�X�YW����R�Vӫ���b���֋�TJ���XŢv� ��j�0Z��F�UP���:�hڍJ�Z���Y[(ƴ\�[ض�R�KKD�h����)Z��-3[�	�T�m]q�Z��h�[Fƕ����iU��k�����m����V����U��ܗF"��ET�V�:�%��fU]vi[cḻbdv�F�A��J�(ĥQb"�����-����mU�rj�"�[h��Z�V�֭��(��kR�:�d�4h�*���4��c[Z;Sڔ-j��ئJ �2���m���k�҈̖���m��U.,���J��k*.e�ɝKh���ۭL�k�(�ӫUT�-�TN��h�*V�ήi\�c�������?���亪0��8:<q;5���XP`�����l�=u�ٓ#Ì)t��7a2�5�M]>�����m�����L��v{u��qg��z�$�wV�a���)˳^��m��n�Ϟ׋Wn����e �g;F�;����U�0s{�](p�nv����D�[e����FL&�ܠn��oa��6C�g�N�9ݍ���;r��o�s�uu��+m�pg[���J�g���`�u�7�[���OGW��V��G�l���.O:����<nd����\���qv��p�]�˫��o=��4�F86�l��^�gqt���F��Dv�"ƍ��S��4.�Y^��3���(G=hn�n{��;[�j�F�[v��{2�n���]�b�W�r;��d3eې�θ6೻!q�SO\y	玄�ͷ�xs�:�2e($\{u�����Ry������h�q��x��6�Ԗ=(�w[u8� n'��盷�9�6�,n0ck�'XI�u�ն�&l�]�@�ya9G���Tm��[���ݰ;a��u�<ẵY��d��9N �������N���ې'�+oq9ق�ݱm<�p�W
M�c�7�w���zSv�y1��Fn���ź�\�9���)�������,p��1�ckY1�u��km���ܸH���4�T+���LT۵�u�:������WSgsa�v�n5�T���ݥ������{\�۰��<:��u��R[��fwk�'\q�i��=^ݼ.-��1����[��Kե��٘�V�v����i�z�Gs��m'[���V�z�ö��=(�S�|X�m̓g��mː���x�3�dO]ry�4��l���>!��u��.w�R�mb0��V�{��;�tKg��[�]���x�\בl��Z8��e�{(��0w:d����[�C�����۟W�.-�c+t�F�9�ۃ۰�U��q�s��c۝Q��GQE7��ww{����kX����be�k��9��\�=���P���Nm۰���S���ձ�q��J`4�����g=��g��`�E��C���t�؁75���0rh�D����'K�:���v��m��;b����6]�Vtp�Ӹpw\��GP�9`����v�v�-\y���d��":�����B���ܛ��V�����m�C�ԗ`�wY��J�u�km���i�Ͱ������m��շQs��i���|! Z��i��<,�D �&�p�w��3!��d3�!�!�T+o���!�@G��ԟ�N���$�A�"H���d��2L�}���r���d�o{��/[��[z;<I�x	�o���8���>E�@��he�/��"H��/r�!�d3��s��
�!�ɐ�fa7����!�<d2J�C���-E�B��dI@G�z{�u�]n�3����8���g����C�*J�I��3�������g3$Ʉ�yR�-:�����B����#HI30䙙Ϟ}�9�*!�_��}�!���tݞ������:(���,� "_�"H�o9(����l�3!����}��8x3�2&C!�!�_�{�!��d�
���D���۠p��~]�2=O�L�g�����<O�2h}��y�������V�vd�!X^{���?>$���I�߽�qϯ��cߺ�:������J�|����;B��2%B���}�8�l�3!�T*	�_~��;C0����5ۿ��6u\�ۮ{��c�`���v�G#��Llr�N��o�g�燿��z�OW���u�C�C>w���x��I��MC0�}�8�3ę�2L�&I��~�q;L�3���Eߎ���$��s�w�9�5&B��\���s�x��!�Ͽ��koF�n��;C��C&�y�É�C�331d��U�'r��G����6�Mw�݅���e��Op����lg@F�1pK��R�=Q-��6w
��8��1,j�f�ě�����x�ȁ��{��<C!���!�i�}��x���d�
�jk���I�t�A^>Dy)
ߔ*����}�]?���N�dǛ�����뮛�m���'I�����߹�xGę�9&C�%���;����\�!���;/�_�O�}^��s���?d2a�fM����q�2%B��ɯ�yÈ�>�.bm6i�14@��`�=�>�>�y��&�g �z� ��P�/;���|g�3��d��&Lm����I�*J�ܓ39����<C��������>���!u&C0�߽�C���v{�~i���i��Hx���������̆ffC?����<g�>�f����Wy�8�$����x��Xx�2MM~��$�;��T*J���޾�<O"t�#��>�ﱳ����/:���#>�ۢ�s4]G'h��᛹-�Lv���իk�&������#���'i�f����x��3�d45&K}��2J�s�q���^@DX ""���k~��Ih��|��C�x3!��2�5��Ȓx� #�/2��Q,2ඡ'PC�9�ߝ}��|C��
������{��C�~���?��L�d�2d�6߻���8���30䙙�����!����@C+>&;\�<6��� a�|��0�n"I�
�,�I�5���N�;C3�fa����{�v�C��d4L�`�/9�}?M*�9i`�boӕ��ߢrcA�.r��+���22.ȟS��c��zO~V�K9�!����^�]2"t�P���UG%��k/��8���a�!�mM��É;;��W�3������P�<OdǛ���l8
C,�2,�|��̟F���yǿ=I�%C�Rd��~p�e'hlRd3��߿u��<�d�d34M���s�x����������Ԃ��2�'LX߼<]��]V�|3>��#�@�'���<	�|���|�����%O"d�1�����N'i�fa�33�����x��Rd*J�x.Ͼ� Y��к����G�K��d���6{Nrok�].�i�5�0�/���;m�IM��;?~OZkz�:Zo����2k���8��Vv3!������{��g�x��RT+7��}��C0T7�3~S����P9�G��I\̓9���'�x�'��^���u�N��2N���7~���g��L�#�@����:x+����$N�����2��q����C�<O�d�d3��}�!�<����d<��;��axO^�C��H�=$>�u�%��^����x��r�>�<��$�T��3�߾��%|�dɒd������K�����q'��33�fg?����x���L�IP��y��s�x��_	{��Ž/][oF�wp���B��$Iig/�eF}R� �� C0̆s�Ρ���L�IP�/�~��C�C0Ð�6��{�$�	(Dn|3�qT���&0�:q��_p���w�$1��Fǵ;�]��PS�s����2�%�vp^U�����/�y��I�W�2L���y�!�x'd����t��oGg�:O0���������2%Kz�����;C}���x<���IP�g����p����IP��o?~��C�x̆f��dɯ^�Èv���n}�q�ܘN�����ۥk���A�}u�pU�����{%ӦN3��tt�Uk�>�����n���^�Uoߐ�J�|����v�I>�2Lj���}�x�8fI�"#ȄO��$zH�G۟W��{���v����o�r!�)2%B��}�!�J�|7���������!�x�M�������љ����'���\�^��m��� p!d3o?{�|Cĕ
��!�cSu���w�%p̓;<�����܃�$y��n"�!҉�QL�{���q�Gę�rL�IR����+�=$�Ȁ���Dss;��˟���'�d2J�f������3���̆C&M���I��߹���=/G]kw]�<a��3�{ϸg����o�P�'�P�0j������&B���$�z�߸q'I�d��G����O��7�:KW�<ar<}��;B��V{������g^}�ӣuN�oZ��<C��C&�{�É�C�fa��̆}�}�x�2�w.�_h���A���U9�$a�9�9���{�$����3$�����<C��>;�t�����<��G:꤂�w�R��墑/�]�P�o\&$��~R<|�5y�3B�D=�{P
F�d���� �o��m�^A��^���v�����z8n�6�I������i�ݐqq��x������t��6;\q�[�[{nB��;Kyw�#�y�\=P��Ŏ�;�BLv5�#Ҩ�:.���uv��3ٲ�z�ۭqMۃ#Z*����W]�.�;�u"#�ݞ���5��%�\���v�=w���f73G`��@�dI��6x]�ޱ���K��ݏAv�܎�g;�G%�2	u�A�z���)�:��E�������C�.�w�w��	�n���8�ę��2Rd�o���t�Cb�!��!���߻��2,k���r��	��]����2���L���8�bq�u��v���c�z�U���xA��O��(�W���[4W<�������Y�L�d�0�&K׽}É2v	�fg$��s���܇�y9I��)2�������C��<�8����poO����n���w����M����8�!Y�3!��2����x�ɐ�h��_}����W�����C�G!�a�d���~��I��+�2L�g�{߹ȜI�[�V��."q(����~!�f̟F]ޠ�l�a�G�Ȉ�y"{���2%B�����p���22̛�~��C�}��߯�������!�=��dɾ���8�i��7����v��������0�r����J�IP�/��}�!�J��������4��]��"�Dy�Ov�I��2L�䙚9��}�x�����L�a|���;IP������s{����pԷ|y������O6�]�6�1�^.�NS���0�E�tS������N��զ�[w���J��y�O��̆IP�����<C�*&C0����x��Q���v5O=���Po�"Rw�d��̓8f|�{�!�$���������=\�oGg�:O"f�>��}f��>^(�"�v��0���e�F\��
SD��(!q~!W%���}{�|�]ՊGk!S��ۤ�Tt��=�V�f`v��L$�z���oOo]� ?�v��}����2��q������t�!�Ʉ2������C�x3!��d2��_�>}��H�pDm�̉#�@���Q&�}^�Uo~!�9�������IP�1�fϽ��|g�2%L�&N���������yϾ8����d*J�9����C�<9I���!���߾���C8��϶����+M�2'��3�$Lت�]56�(�<� |�g���r��&C!�!�m���w�<a��2J�I�7^��I��g�y��:����%x3$�fz����<O"q&!ou[���@�p��#�E��]�l�A�&f�I�Ƥ�z��p�t�-��F1���jƏ"�� "��&�!�T*y�fd�~��C�x3!�T*J��~�$�V�����zy���c�n{����L�]�9���Δ���7[պ�'�4��y��5�����E�u�iF���T+�;��ψt��I������q�3ę��2h&I�n����$�Q�#嵼�:�2=�)��|(���2%B�a���y�<|�2���ǅ:�����[���v�d����N�@Dz}�.6(d�����ϝ����&C$�Vo=�����<r��C$Ʀ�߹É;C7��}�q,��W���Т��E��&\"b������)�� +��X/s�����3��U��11�ϧ8nI�3r�k��?k��k�;mʑ�z��ݓz�j��)Ւl��p-��{��#�I�~�I�;?��"^ǭ"�*�����农��ؔ���(+�D@,�t�^�����dt2eS��Y }�z�\
J�)$D�,s��"D^O8s���zU{��@�餓
3*������W�����?�_�{�����{*��4sB����Vw5ӹ8�=B��#h�qQ��������	!�ٔ����v�(I#쾮cu�3W�+x{�=�t���t�z� Xd�ZP�Q2�u�Q݇�7]�&>}\� �6��e�����e�^2����
sa���)�jB]�G:�P@�Ӯ��~��{�fvV� 	Q������g5���0� ��(N�~z�Ɩ\��0�@�fu] $�g�`��z�T�����u�T>;���	!Uj��og�*�����I�k&`Hˊ��[�:�o_%���vw�L���?�������|�n�f��]0���� ��O�b��%x����)X.�Nۉ�=ަ���f�}���;�&���v���b7!뫬u�4yT�۫��5�<��;���\��{�6��N�b$��`�^N��$�z��.7�t�7�┒>VU�Be�z��F�𕉔Q2���d 5�������x��PG�@z�=c� ��7 ����gi=�x~K��^�	�X�6E3 ׫�"H_~z'ĒGz���W�뼛��� ׳�Ȁ {�M&
� ?&�P��U51��[~��<��wf��Y.}�)	��[�>�z��]Am�����3�XḊ�XX[�R �9p��� �*��+�mmF<�
�W1�$۴�G�F�	�"�nѩu9`�(����:���������H��f����if�A���9�s]���%p2Eol�o��w�~w�� C_{���5�������m�.�p�cY�l/G]�e99�õ�u���:����g�;�����p۬;J�z��lA�b�[�(6���W\�ӰS�p�9}�#����a���$�:�Rm�n���u�v^��g�;��w�U���sOc����[����f;�@籎R�C�'\Y^X�.�o8,���v�v=Tv�0�cʹe����rsr�u%Z����F�u���
���3�瓮�.��; �oK;������?{��ĈU52T:Ksg?�H>ͧ� J ���&36�C.��M�h�}K�	�"s��� =K�j%T�� �=�*�6���TUm��'��9H���	 �z�,D�\��B��#�f�$>��n*)M@LMH7l�d� U�T�IOA0�3�70Y�l`��e�>� oU�a�|"���h����us�W>�U}mD�F�@x�rؐn�X }<�,3���*�N��$�W�I����?�e"�!M W:��%�Ӯ��o�\[��_ۀEMy� @.{WbH1��H����+�޻���mZ=ltu�������c�g���=�uu�>z�ٽge�ܽ|��}��g��&�=�s�t�	%�j�,H��1�1�7�?|?w���>�*��}�P��� �a�Ӷ%��=�؞�o�ǃ��9���Ʋ����[=�Y���Z/�EЛ{r�3��7@�ww�~ďn9��m�q�v�ի�q�V���  LyO�
���"	��$����

u�L�%���<�� |�KR�D#`�m\X| c�����}
���� ���_�" 2�y��ۮ⢔���$���vQ�N\PF/9�F�@]�T� "���  ~�޽y>]��Ý����c����8�n��$��;s�0 ��p�-�D�yOz��[�J��ӬI'�u7꡸�9���v�N�N�u֛���]���\����%ǷJ^��b�-��;_?�~�s�3����>�R�>��p��� ����F^Y�v6�b�'�]yWbH��q!֣Ԧ*j
�	��u6$�3ϻ7	�R�:���� �g���p�������=R����	
����>�/O�8H��Z �ϲ�E��Qu�����<����nѧ�w���_}:�Ϋ�ő��w|\o�=���� ���)���}�wh<OG��I��t{�9���Xr9��t�7�9��>�6����w���Ϊ2{�.w���.g��]�Չnu\���=���2O9�������5��a]�,�V��xd8*�2�����{�sm�E�7��uXf�z+�FO�zs~I|0j�9��o���T+�-�&!�^��w\3�C�0f<Ǐ��p]b�pE���r�6��w�������3��?NXQ����ʯF�jy�K$�Ӵ³�V
�a�1H���F޴vo3�7ca�1K�N\���}0[�o��=�4�劇�f�SS�2��^�xoۉ�>���g��g#��T7�9��=��L�b�ܛ�Z]U1ה�Zޣ�n�b�ih����d~My�����w� @����#���[U�>ߌ��J�4p;{s��^��.2��Sےd(}��X'6���t�pqE�KP�������{�嘆������X�;�G6�j6{ȅ�ۅ;"�,�,9jO6��f���&������n�F��ů���,�W��p�z]��̷�`�L[�<sOd�W����Uy	}Nɷ�x�Fy��qT%>P��Pn
t��Ͱd}K���؞���]���Ij��߰��ʽb�� �]��.������E7�7v�ŋuc��c˗�Q�Uu�h�z�K|����#zg�{��)7L��m�G��ء�2yIR�2��������3,�ȚX7��Ϸss@�wa�ݽ�k`�cX���`��mV�;tR�tT�YX��f�ƶ����EQ��*0f��U�U���mUp�T�U�j1��mJ�l����5��klT��ԫu��є�ZQ�+*�m*�ȵU��A�����* ��m�Ŋ�:J�R�1��V�K���D֥���q�R櫚�X�Fԥ��E��F-V�kDb:�f�U���,:���6�ǡ���@m*0�(��r-b��KJ���R�PX�h��b�����KYUX��+[z�p�)j���-��zJkKj"�Z��`������[m�֢�h���+�u�"�մkX��XT�Y��EP��b"��"��V��eEQR��#E�%b�J*�W4E`��.E
�ԊR�-���-�YYJ�Ym���SZ�����U�QR�mZ�ʂ��m6�h�A����Z-)QRғ5�Q ��[h����"ͩl�_@��D�z���@_���I}ߥ����M-DM)
!D�%�kmV�=��ӹ�/'��@9��o� �w��jk*�7�����(�Ϊ"����2L��l��[  ��R�t❻��DZ����~�� 緥��wz�`�w��Z˓��Vbd�3(�ѓn���<�
�n=^ntu�WS�oi��{�6f���M34o@;s��� �Η�0� �;�UpzU��&�k��J�ΛЕ��?T�!%
n�Wν��+y��T%17]Z�g��O��ggM��H���cW34릪g�$!��z��M
�PP�����K�� 	v��_����6{�W�TN^�h{�[� �]ޫ���v
f �*&���[�9�	{*��OvKbD@ު� /g���=U��pR*�&н9k�<��N�<���t������q�p*�׀T��u]�X��<l����ma[,�ps��ff}���o����ҍ"b�B�K��}a�%����ڏR�};�tL��9�kٷ� ��\X� ����H��ڪ�1���7�(DC��("l�V�&�X��[���vp��k��߿�s��ә&KL{��Y��W _OX�?yQ���	�}����$�=�حw���$���SK�ԣ�#��kw;]���1�� ���U�{<Ę,��t*y�USyG�+¨����IB�o�O�T� ��9>�a��exޟ%� @/w��D e��r�e6Xi�TJ��=rU��ۂs۱ W�U����c��>��ɰw�8�g/�I{}Wk/�)�	�UPAt�Ν�� '��l�Z��Vc��i8^�%`��z�D��#��y�z!�P�z�vƢo���E+�!m����W�fk�wcȏY��L=M���S�����z5���K$'-���$ɨ���4a�"
��E,��u�ο���{w�-�b��b��n�T0��5��p��q�����!� ��1����6*̸�vN֗��&p�����7jܢ��S�!���n�j�z�c���mݻZ�Y����v�M����R�;����c�s���u�1;�kq+mǱ�<k�����Zܷ����t[�����8�*�@/Ѩ(�7(�s��NN�7FD��mك5��v�a��:���5��v����B�.1�8�۵���5`F}���,o��ݿv�"b�T�D��׵K�^m?�|�u7 �1K0��J˜�wz���ߺ��35�LJ��S*d�--o�<�tp���?-�Գ��xo�� D��� ��/�\�������"H��
f����v��1 ��l ɚ�W�$��V��)�D ?wS@{�zUD�TTI3B�n �V����כ��� 	�ʴ�������K��j��=�>��|����!��>�R�S)M$��e8b@%�긱��~�2�U�춟���l wz��J{�ݹ����j����/$��v��&��/c�xթǪ�-Kͱ�ȩR)S�vĢ�����H��om8�$~Χ" ����W�s��蹬���;��$���i8�iF�1T�H"F�w��� Ȏ�n��,��{d�D��/]�TC��8-�X6NL��o��ڲ�^�<����2f����h����f�=��w�F��3��}��{��=����oSI��/�꿬D@p�N�G��YV�{s�萌�nR�P���$��o���@ �w���޼MŌ)G<`� �i� 	=�ٗO:��"ڄ�DT����gu�
���� ��/g���ZmU_-�y^Eݧ�^��`}�u�U)AT��4)v�>�\X@}:��8�5m� ���o�" �^�Uň�2�y�,7"v�Cy9ѦڀQ �n��"`�n�����t�t��.n��Njyg����.���R�S*f�s�{�V�@	n���� ��r�'�>���γ˲�m$H�^�7�O
��������G����ү{*�  ��V	Q��&<��婚�Y9�ά��ZQ�LTUL�7 �r�," �2�� >��UR�-�k���s<eF��$)����*�q�q3�G�$-�wǫ�Gߦx�(Y�HӭnC6 -�ٛ5yD���{�����{�DDG�W6�O3��I�'��1<	��		��US٘��vc�� �q @uN� A�oS6�79�q��$���,�;�QIJ&j��-���@}�O�d�{&�s!n�Ձ��V e�)$��oSI�:{�^���Y�����\�M㶧:nD�W�KG�-�]�v�¦z��ʼ�v�z!B	1�Ͼ���*,-��[�_�a�%�v��$�g���|�Tf_����e�����PC/�|)����&i'/���M�W��]�cZE�\n����� �>˞�)0Y�괘s��.��}�l��1ബA�"C��n�t|	/{:�0Ӥ,����d�:���	g���@{��L��P�H���������XMƲ2���\Y�1����u6@ ��q�B;<�]<�f��T��q��g2��z�����O�A	��UoE������k�.�e�fʤ�	����D}G���a�7A��7)J��SH��H�=��l �m_�e��Yr��g����� o��� �f�]/x��I�[H�Q:��%U�tWo/]�8k;u��z[^�W�G?�o�c*u�O���U%*fj���c�� �v�0�" �{]E�k��3��5y����>/o>���a�s��R��	�/�;� m�W=������Vt:I$�:��	^�U�#�|ㇶr���48�{�?C�����d��`D���� �:��" ���#sݓ�{�V�N��������J�(��a�v���g2���o�$����bIw]+� Y�w)f��4�nR`��� +�Q�LTUL�H�{�U`} �Y��o�>����F���k�M� W���f�t{�7�Ϫb��u����KܔO_^:fnu��U��svɊ�wH;���Q
8��A�K����^E��B���h�3���D}�{�߿���[p�v�q�)���zҝ���5GU�1����m��ܺ�[�<��7�|Em�<|�˵�;n�͗r�>y��gsyۭ���[�LǏ��n�Ȩn;�VۖC`�9l�x&��Dg�l<鰤;ѝ�����n�=w�]K[z��A��:!E��!ڞ�
�t��9�,v7G.5������vN cG��J�s����Wq#&�/=[�����2�z<=^A�%�@\���������~���� �U�U @s���-��.Q�a�=��o� 
�J��p-��$ӄ≗�NFʮT���5w^ծ� ���� ��z�H�)vr;�g��K�Ǆ��h�H��Q2�%��UX$|�:ܐ	w�a��)�9]{^K~ /:�%pY���!���\e�0�&�z"���@�0�rU�,�� Y]T�� D�լI�+��Lj.��=��ˀ>y�\y�JhR�
 %���4~ަ�܋���Ϣ�V�Z;wI+	�N1$�gu^���
q�����P�R�DJS('�.��`ɽuu�c�[�#�sq��a��&���W/7��>Q�LTUA(��ݕI%a9��� ^wSq\����j��{���q��>�kr��5�$	����n�=\�S���d�9{�􇗂���������	&w?62nz�Iwvw�R�������Sy���v�w���ڼ��� >��0 ����n ���}/ݔ^��d���%EED�3SD�l)���^��` N��{�T�Gw���e� }���" �� �?\�)AT��*�]��=H�q�c�8�� �3�u�> ��[� � ������z�����w<��Yy�LTR��3I9`�C_NЯۚf����� ��c� /���@@_OUě�un}����>�j��Myncqr�B�tM�<���ݸ���s��wV�3�]�����Y�����������oU��@�u�z;�Ƿy{�-��G�A{�M��ߔiA!#a�9W �ӷ{j��=��S�t 
�:�� |��$�z{���w���۳�萌��)|MB� H�{�N@ �'��B q�]~�N�{�\���aɱ��/�3T�A�;}��a�21z��!�Vg��^&���t�Z�s��(ճ�j'S�-�i�o�}���we柠� �ަ� 	�s�(���A.a(I�	�W�R���m�����M�D��X �:z�8���q5����ה�q��XT��)&UD�p��)ޝ��zh݀ݜW� �]7��^�Е�)Ξ�
]��ּ�S������C"W;�8ذ�3�q{�M���=ll���g=??y�4�}T�4�����i��;W�$FV�1��=W�.�ڒ�=7�S�%�r��
7�)2%IR�t�7:u�9H�}-��7B�������+� ���$�w$��u���t߲�� �{�8���L�7�q�W Y<�� @k��iR�����݀ U�P���n"C2��_P�DH6��7�x�����^f�� ^3*�( �s 9�����G�&���wd`?�
9�ve:m���{��.<��d�U�3T���v^墇c�ݐC�4H���tX�s+	�� }�E{��z��+gxJ���I*h�-�;s�8 ��_�[�*������{ A�ݩ���/g�� |����f�{�}��8��f�G�a8	�ן>��qvx#�Q�q��[�ܩt�;��wA��������n&�I2�%�@3�W@����!� @���Ҋ�|L���i'>��8}�t"d;�!c���I�1u��BI}w�����ZR��}��I���=c�>=�6�	\GdӞ���/;�ċ�߬>���"�D�i*P��g_�@ ,�t���F{�ooUdn���Up$AY��Ĉ����'k~#H�+������LHe�4���$޴�cS��v�` ��Ss�|�{�.mh.Ξ����&�EL)F̟vKa �Yޫ�;ow�w��oW����{�[ ��}�-ݬ�L��Q9�����~�q[�;KC�7\W#�G����\�k���۳��jW�r���_Cp7����y�6G�y��}��&\nz�S옮m}�ۉvXs�wrn������o���rr%��z�6n_-���gj/��33���tvZ���Ew=����s*\:CI�ڣ�L0a��w����鯶׹R������_Pm�G�y�g�M��-Ǭ�~{�NU�q+6�ؽ9�|���#���2q]Iɔ���c	'��&���9�۷�6ʚ��3���T${�S�{h��Z�v>֚���<+'���G�ܭѪ�N㽘w�]|��_V�m���t�sS,��mT�|VRb��G��oDP��G����,�8B'�^�c	N �T�ݧO�YCŽ3ϡ7��h�I�EA�h��&��^A"狼��;���h2we[��o�wA㾌J:i#�k����G{<�h��Dn��Po�����l*v!�g���#��qA�;���G��o݉�p�z���ҐΪ��PB���O)SZ��He���`Q�ҭBc��K��>�Y�l��~��m��='`���u�ܢ'=<sf������|�x�NM�i�$�@�9��
���%>�S\�|�����M����=|׷n�D��gwZd�j!3i�/5�4�@�Z�
f�C��L�La{#	��93E
7J�n��ÙPT��l�Ȣ,ͅ��y�r�=�;���9��\�>����4r ��F��󞛗\�����v��)j��&i�b3�TQ��e�T�,-�`��KkF�mX��(�*���ͣ.,��`���Qe��Eu��"䕣X
,m�)Yb�(�j��AAV:�kM�9cm)TEED*,
"����E%UEE-,^��N�b�gC����fjĨ�X���X���5A���r5
-�-�Qk)Q�am
�\�V�R�n������6�h�QV��/Z�4� �
�ʬ�6�%[e��J�J�TKJ,[j���*��:�ͅd��`����X�iV��h��UJ)J���Tj�E���Z�%Db����I`kV)X���J�h(-K[Z[R�Vd�fֲ��Qe�VB�*�j�PZ�)j)-l�Ҩ�TUcZ���DU%-
��T�j"������Y+
��dE�*�1��(֕����������d�J�em�DKm��TeZ����V�-�����Z��Ȃ'��瓫��uo[\���njLn9Nݏ6��d�.��zݷn��>��c�8�Smq�ɱ����r�[���7U��v�Wr��n��k������ݺ۪�����]�uN�J��Ur5����gWq����k��b��݋cb�S�$�c��l#ڮ,.�vZ�<�h5�Q͈�,hۛt��K���4�Z9��ԗ6�ήū���w�1����wI�Zm�'E�l�^�F^�K�F��7=�v�ǋ���e�ێ��c=��{5n[ik����y-�,<Q˛�ݤ�/n�Kh�����qqu;�[ű�=G7;��=�>ڰ�����tDg���g�J%�wnY�ViAy�j��X�z�B֞��o5h9�vy�l�����nQ�T���g-n�/F�C�s��㶗���ݱ�q�9���նX�<�7B�9	���1�؍A�=��x�JN��{�֋�\�'%�n��W-�h�0��\���R�Z�&��p�z���̹^��wO]�kϏn9�v�UnM���tn�V��nK���v�m#�kFm�Ź��]�ts��q�K��iM�vԩ;n�}.͖i8^�b�]6��꨹G�Ν�������#��cc�֮a윀Z���	�5q�ݶ��]�����eI���|>A�ڽt�:�˳���|��1�'�7a���s��F'��v�!g��'�oOg��P�C۷*�vk�Q�_.���`��E���m��v�c9�Ȃp��ls���M*t�Z֪���)��]z5�6�G����k���ϓ�1ɲ�n:簗+�6Ms/����t��JyL2Ӌ<u�g.���xsU�=��&��綹���5F"�e���v;�Gn2�U����y�vMط'^��S�mťv�'�)v���:���W1R�=� ��=�i���m;l���ͬ`�;�zy*rvkzwO/7�= S͊nA�yK���X�l����v����}<nˣc.��rkdʛ)�8�4lO^R�6�u&���V�����w���wϛ��tn�66_=/k��>ss����!���c���muh��:�Hb5ƣ�n�n,��=s�k{;n§
kC֛�`��>x�v�&}�e��Y�����q���㱻/ae����.n�w�:�땋�x�i����t�mq����-���t��.ۃ��ז�m\&���D����=e��%� �ͯ+��Yq�ۢ�.���O���-�Z*��Nǐ��=�C��;JN�lx踈��k���Wba�i�A=��ߠ�0�(i�q���uK�RI+7:_� ��V{$�I�������$@\�t� M��L�Q3PI2�%ۈ��J�&Eh[Yc��9����6� �]ުJ�sg<x���9��n�F�Y+͌i�b��H@%��`��%eQ/��Ot���D9��o�%��-�)2%I0A�~'��z��AW߷��oE2�>��Uq @,���o������K}7�-'��L��S`��W` �9���g���Ȭ��w� |�����H���qbH�/����^*�}���ٳ��m��e�tvu�!	�gG�D�����$��ူ�n:��p
k�������7n����A���m?��}Wa @}�Ӏ�]����ѩl����6 $�������c-�m"�)�>&l���H��!s�#��*دb�V��ǉ�yG�I��G&o��:�*��slX�AH@����B*t5�mj��E���b�^¯Nn_�{��٭�T@�� @v��+�~��I=��{�U9vm�I3��� N�	;�J�A:���7�꿢�}��`	9Jw�1y}V����RV�����T����EL��t��z�G>e�K��Ӛ` �gUؒDy��� ?wS�W��F:�Xw�J��e"�HJi*0�ݫO� �u6g��iU)�e�W.�V�U\A�2��@?wSa��*2��Z���E���a�Z$�ڈn& �U1Y8�#I��al��:�i��9c|���7���&I3�=기�>�ǛV��y�Vã��r9�г����ڤ� �ʶ�럒&�AIH�V�}����P��~I{2�, Ϻ�`|���n	8J)p�����+�����þe�u2��&����y�@ ��ӆ$|!�-`����4����ʨ�Ř��9�}�w���1�l�tU���)��G�������u�eꯅ�.�{�ߪ�q5��vX�y53X���~�o� {��I�<��Қ�fR��D�%�3� �[�3���7���r#�� {��0 �Sp�+ޣ��+w����90�����i5�9�{�N!� ��UŚ���r��U�1#o�k��n�` �z�,�V��ߟ߹cM���9'Ge	گC�<��p>��]�sq�!ŷ�V����>�e;f�2�y�] ��M� �U$�3.��1d���i' |>���L����g��, =ժ'ͪEU�lH����	+ުJ�&4�`Kz���un�䉨PRR"S��N!� ���ń�M4f��S�� �� ��z��*^�T�LR�����#�&̟Z.��|�@)��C "+�U\ }��l�+��5�ٰl ����B�*�첶���c������T�B���<�^��T�6m��I��7wGN^�{�0�$h��JA��Gr&���=<~��Dל�ԒCH��I/�w1%��i��<��=��~���n � �*�@_u6z��+}/uz	�R�9x�ҳ�ms��h4؋�E۷<���jy��	��� ���4��[�O�$|	^m]� e�[L
�������3�ٞ�� O6��,����\AN�F�k�B"�nP�(I4�*ʺ؆ |���� ����b��o^M7w=*�3}�Y�yaa}H��n {j��^u8a�*<V�j�nM��{~ ����>2�����՜ϒ&�EB��S`��W����UJӏX	_e_� @�춘 ��r^��e;�K~>�T��-����%��󹐜$���2��=O;�μת��Iu�*�#���lB)l�؉w�.���k�������=ӆ�Y��o�"dz�K��#p�aQD�u���_�`�Ӯ��I�����՗u]<����D�ADDp!�M�ٴ]ض72��!��*%�&'c�7/#��u��6��[���Ysノm�u���ݳ�����Sv��[�vv�h��>�����`,��\�V��K�[ۮ�`ؠr�"��{��xi\a�ղ����Kq��Kkf�W=[�n,��M��M0v�t���x۪IϷ=��u��t�m8�����U��ۤ���ј��ܥ�s�]"�k�+�v���a�~��C!���$���� ��p� �7:��=>����FHwoy�I:���Dz�z�-!D	�iע7���5u%��d�E�گx��^���[I$���l ��b�����ܜf��01��-(���j��7+bKٝO� ?�bcw�<�fp�:�)��,�M\�Y` d!��(TI�N�yR�Wb5�C��8� @ٴ�@'�OJz��� ��M']z@���I)�Sp�S���$�j��)UZ�[o�@n>�I8 �ͦ� ޫ��Ĺ�/���k|�VT� �4U �%*���xz��:�y&�s���YI!G�ȉ*IPTA�����p�,��h$���N �[��� 	=�^��S廊����� ;������VL̤��*�]�}�����_��
=o\��mZ�n�Ӿ��u���G���p$���N̪�j�Z�6��s^�dL2z���G��33��ͻ��   �Φ� >��\X�&!�ьQ����L� �<(�e����e6 DO:�, 	���ތ���󜧫� nm[�"$���,��e4��qE:���{sKܬ��Y@,�ؑ �U%`��k��uc��u}W�
�#H�*"��[�{�� ��S��g]��� ��6 �u\X��ޫpa�����r���B!	�
�PZ��h�runF�A&+�{[���r�7 \󊏿����7�)%0JԮ�k��I=ڻ" ��\ ,���yW�3�}�+{����p�/��8���$�2�(�5��a$������X�ϫ����}�I\�������#}֟vߝ{~�WL̨ER*fJ�v�}긋�Ko�\9,��G`��4�`�G����Y2j��U#!33�VdVMVňo2}�k��m�΃�'��;���	�R��2Z���o ����F}������D  ���X�Y}?��!��J�*	B����LvV2̽}Q�͎����ʻ� ��0 {�OΝ+�Z}�R6p���{�N��,&����9���� �gU�^�EV)w }�ʫ� ��N7" �괽~�zg=*:�������\����W*�dѫn�;V�����q�s<v�x��X�ܜߟ���㾜�wGI7����$��'lȀ ���pM��F��H �{/�|�W�|H�ڄE@"Sa��O�@vu�/>�*�T���L�s�| �z�N���?,0G��-p��)��h���	���@ ��p� ��2H��l\�VYN�~� :�<�H��wSI��2,�Z(�Sgč�^���&?��# ��� 
��~���}�Fz��]�����](C5��Ӷ��J��bzǏ�2U'�Q�j�\~k�͹hC�	�E�޴4�����f׼���dNN^���;j-�����"#oU�zBy�J��*���tý�V��O?U�x�ݚ���o����^�c��73i�� �Oz�Z+��CK�g�~�7��;�F��kn�[�9�ا������v��=���������fS�h6��t@v��r�/fu8� @$���ӓ	}2�N�z��"��7 �F�0TE$��,�U+�����ٳ3���� �u7 I�Uŉ"&saZ)�ʑSO˃�Y�v �l�E@"S`��M��@$�j��	-��^R����WfM`� >=��i8��r& 5G;�BN<Z�	�SK�Cjq�=� ����N!�� �*�Iel��sB�w^S�^m�7����"�*fJ�ۀW���#�����Ne?��U��  Oz�+����M"��Q��oȮk�LNz�X1e���6�T�L��S9�p]U.��)p�=WM��O1w��Bww��^���ƭS�ɱ4��k\��� {¤�d����R�P�/5�*��ֺ0���㞋���2I�uI+v9����u���;��A�&;hun��{!=.5�ܮ�C.�S�PY5ɜZ���1rc:��q�����Ӭs'�>g��[-���*�-����s�iv��Z6�Dz�	ƻc��m�9j��/S�y��Yۀ<NMr����Fu۟=��mۏ8�;�6k�d�q��5�] �km:�{=�tXmy冣�8�<�WO��b#�rkf��)I�����0(��Ac�苾�lH�I��ŀ���0��ٕ"����ӧ�S�$���5��LI��e5'�j�(.��N���@u�]��uz����U� ��z܈����%�8�o:���Io�� ��115DI-�=�J�^O7 %�%����v�/:��>�ݪJ����bq>�\�E$E	M��uo����5�S����a @%U�J� >���8�2��k��v8����A%u�g�i��)"�)��"n��l" ����1lկo�[S^�U$��~�n  ���4FsD�a�[!(E8,��q�>���+��\/ny��`�eK���N��A������"�*fJ��Tk��ov�C  3���^>^�O��y��t#�y��V�"�J*�����o�*����_��W$FY��㇮����n	M[�v�$��?�m�ni[]c�ctE!'�	>��0�o�l���ٺ�9�Vl�W�˽��z��]�����괓��~�� 쫟i+3/��/+b�ξ�����5H�����	����I+^m�Vvv�O��� ��i'�<ަ���QJ)3-,s�͚���p��;�VW*{� `�j~�  t�\siU�};ޥ��i�"'��!AQIBSa�� WӵrV���Dޏ�}�f�զ��l /g���|]��S�;�v��r��T�TH���0���m�&7]:1�	��s�U٘n�v������>���vb�t���a @'���@ �g����O�[����O_���@?wSI�7�dȠ&�T̕����	P�G^<��=�[��V���> }�M� ��ZC잉��m��D �~���J%ELK����a @,s�H@ �]?paC����1b��ve��Ύ>��n�xMv�,�N>�5��4�=�l�y�}׮�v���[��u�W�Ù��S�1=5 �U��p{s�m��n�3���goT�8���C�-��6a�Ǔ��}Ƒg�z:�N�-6W�<�N]�M�������u��R>.�Y�/3Έ9�}��VN�V��b��q���8����w�����5yo���]x�=�bq[D������R�-�qs���9{�+O&���i��x�6Gj`�~�m���Pr�?�^�n���HT+�䑹��Lu�݋J��`�=����+=�/��0v�KP�wM��^ڏwm���n{x܂�����77.{p��9]�<g�Ƹ.k���h��E�N�+r��ߙ�g�[7ሾӍmr�Vq4��S�۱���b@I��Ş�d��z�^8$�.�Nt(;�����:z��p�ɚd���E�6A�W��]��z{9��>�p��0.�y��8j�b�qa�1��x^��f��y=�[��|�r�ޱ�vf�˞�67~�vN,�i�vC��r�����4�}�>[�Z��5Z�F�����A�y�=�=�&����w��ǲvK���꩑a���N�1��+B�������@�]^�B�?vg���s"<��}���"�W�zM�*�g���T�c:����*�Y��w���3 u��W�Т�u`\��;j>E�W]O�U�p�"�ʀ����0��Q�I ���Y9k��)5�!X�mm��i]h�*V���Զ�+-iR�j�-)E�e�A���*X����R(f��V4��b0ZʪV����5-ed�i[j���mZ�����e�Z6���UhR�J!v��h��UV6��`�5���AEԬ�U���"�ň���T*V"U���ceB�k1PR,���4YR����Tj���`�ZZ�e-��c�ҥj��-�B�����֨�j#J[D�QQm��(Ԭ�J��#	U�Z��Q-
�Z-V-b�Yb�mm�֢�D�*[QQ�[*-e$F��
�(UYK*�EU�Զ��K(֪"��#YJѭΉ�j��Dm�Z�QYR�-�����XTDZ�kmm(�R�iKV����H���"����mX�j���Dab�c
[�J6�UAQ����R���իi*���i[�������~ ���� 5�긐�ٻl&�!CS^���y�4��a�K�^n��H�5�P�Wc����!V���tݤ���]7 @�2"&*)R"f[�y;B����:��V��>�g����s�U�  �9W"H1�Sqr�k�u�ҥM�Ȧ�e�&;��O��K�8i'L���m�r�\���??NT��"���{�� �ڹ�uZp�v���S�:�� s�ʳ��RD2S�&\�b#;.f�'��Y��c�" ��m cp��q�V�g7��\���Q�"5J�d���9Ϫ��_m8`�O�j�s���wM,���9W"cޫI�-�$D�}%MMTK� ��[�q�ɝK�J~U=B��!��i�$�g{�~ˑ,�]T�����K��P���y�Cʎ�j���<e˳5Lo���՚�Ǭ�Gɼ���מͰ��=1���3���c����t�A�?��B+��iMJ�(��P;a��N ��mZr_{����N��H���l7���T:��N�U8��ٸ��j����\��b8nC{N �atuqv�|ms0pw�l�fK:"�s���a 	���a7?:�	uWq">�_u7�� QR���@��3�����~x�Dz׿�j��>�m0 �9�-�@y��a�݉�"s5Q{�Y�h"$�&l��0�����` od�z=Ț�*2�;=th$A�2��Dy�V����&`5Jfd������~�w��Z�C��q ��>Ζ� 5�VMf��*���Ʉ��m LM&[��'=�� ��U�I~��VJU�u�� �� ��z�Gx�3ٞ����T�'�k��W`̢GZ���17���D�u�d����S������gg��ǅw18��"��Yy\_�~<�Ą������Z�g���u�:�؜k��lj�����>���îu��t���:���n7-m9��wX�9�8Q�{e����ƭ�́oa-R^d����/2"\i훪����kt[��3�X���n3�R꫎5��9��4'O�<Y=7��`��:��.$�Nˊg�b�n��E��n���k�G��t�K�B˺o]�����ٍp��4�X�]���Gg%6og�E����v�sŴ͎w/X��b�u������jT�EM�/��{{j�L��p�� ��/�݃�ٳZm����^�7 �ϻe���1-B���D��<�����:�_��<ޯD0��l�	%�z�� }u�;�n�u�d����T��%P�͟vK�� ����!�����W�q��V@�� ��"��;�Jf"����v�����tF�g�@���� > �[E� ���5�:��yW�����o�"&����D�)���v�8~���F�k�:��lb<����D�qUz �KG�P����!���.�����'n^(��"2n���=�����]{��sk�Z^d��0���z8	�SI�aS3X�� �{W�	$c޶��tG����^�O�������PW]ziUJ� ��Bv�7;i��^��5ӧ|v/{��.��VnFd�o*�z6ŋs�E�6t���<1A��x�*1]�0�	�ʋ}Õ3Nn��q:N�l���=ά���P@ ��l }���W�f�"M[;-�^��-�@�c�1El�Y�W$��u6 =�������7!��'�z ���JW A�z�}��J*TP��SZ>����ev�$��j�� H�o�m?��s���Q]���c���k5R�3PUL�����a� ��ӈdd�d��+ ��ީ��y��L���m�T�W����>���G�M�PKmǤ��.r[=�n��u�rl�@�$�(D�7��G���fP�l�E��A |�jӀ" �3���̛��!��\P�Z���2�=%E6�e<Q�}s�0��SF�v�{�8� y���  �oSq @s�=S��N���ّ��� <�ɔ�B�Zp v���q> {��$��?hJ=7�O�N�v�o�֑ą.�1���$��bo���`g`i�PW}U�rSԮ6��Ov*v��z�k�A��M$�g��[��bQ����D�n��(�g=�Ĕ����6	w�i�>Ou]zv&r.&� |n�S`DN��/�%P��S`���q�9Cq��sI-��#�}m0H�z�� �=�f��;x	N��7Ɋ:�5��q�p�B..ܑI��k��E���z���|A�A(�<�����AU2J���Co�jӀ ��uM����w^�G���n }�V�_I�0
j�&d�.��P@#�3�^X�@���@$��l 4�U��<��s�ک��O �^Ǡ$����SQN���O���WA��J'*�k��g]5� A�ݦ�� Oɠ>U�Q�Fj��^�Sd�\mӋ�Uj�� �>�HǶ�+ ǽN��gvoѦ �lNS��������<}�ݠ�]C���a��#l�w&�Sj�v�sh�]����)�l���,�	�]�`�����o�~/}��}��vr��q��jk������ ���Ш����nﷴWm���K�ʸ�u[���������5$((%��Pi6�1E�\ƶ^kK ���b����s]�'d*?����޹Ѷ�	Y�}�i�Mʔ�����H�c�r�=�3s���,3*�>�k�}D��
��WW��`.���[�������1 әSA������ݵ�GfsR��K��Ⱀ�x��>$I5 �nM�@@\˷��%c��{ ��*����u6���RU)��ME:q��[{Y|��S|_���ӪW� �e���H=��o]^����B�?�{�k�ͦ�A �2I݄�n�bD��S�[�v�p�*�*��@%]ꤒ�/}��> �{��{�׍~����}0a��ޫ��'LՌ{��ӣ"Z񱜺aϩP�2���)K��7- �U���˳��n��'���xL��D�PÇ�{F���o:f��]�9T�)W1�]v����<��3��y{8�f�d��&��2���Ϟ�dٳ>$����gtrA۴��ӻ#�]=\����Ϝ/2N�S��1�5ӷ\�u�AS�Hݽm��@M�a�����n��-:5`��>n���퇚������lI�Ž��n%6�y���V��)�>[�;����n�k����ZɁ��:�'�lp���n�R����^�rv� ;��57'7����m���D��$��}�v	_�i� " =��oཻ��>����꿬@ݔ�@��Kꉊ� ����uZT���W�Iu:X@y�V��	�u4����Qɶ�+��\�) �ꂪfA����� w��0�J,��_=��@ﺛ�@/o����~<VO@�3f?Z������W`@Wc���=��l�>��:�=����E�����518,$�f���'O��̫L��W���?y�ý���o���L=��n �KN�>p!�30��ʥ2��&(&`�C�:��m�gF8�E�U�'�.�;����֗um�<��??y��H�NEO��[0M��|�� ��6
�^��l�t���$��l�+���IJ�"I�� ��Bgw�����6g�������BbAbe y���fe�ȓN#��ڈ]5I�ߦ�՗q^s�U�����s6�+A���"�}��������V�#�?cD��S�B��f��b}�D,�'�(�
�	M�y�ؑ �ܫ� #=�:Q����ۘx  �{i� ;*購d��������M�8�K��p���ӆ ��eJW�_�y�[@�]�n�^1~$���90��q�V����U(v�Oz�%a{Ӷ9㪕M���ߒπ�+�7  7*�D ]��(0[�ǂ	�l�H8�,W^Fd��:ɧ��ܮ�Nt��e�ܽ?�{��A<l�Bls�M���B$S�hn~��0����*��2�=�����M&�PuM�UT��1QT v�=�:ܐ�q�=y�l�n�k ������~��r#�nz;�k�� ˅p��i)Q$I-�3��(+�O?��w�������n?f��ߎПx�꽽�m�^�$ r�7��O, �ް�Z׻D��=��1ox����(j<=&�`.�F���&��}�?Z��C���UВW������pDT� �)�x��]�l�8ӱO�	++�q@	�X�� {��S7{�5�� A,���N�ߒ,���i"`uz� Km6U���;Q��?��ʛ� ����W�M�s���m���xFp�Ap<�uqEtm��ݒ�D���rg��sۀ�ɚ��n��B�@��4�`&�j*�T���J�������#�=�l2�M̘��4�wWP��O7��^�)�ST�R�����g�)�k�k����t�y�P@$^�s`A�M'�U��D��5K�g���֧[mD �	����[0I'g9�$��u���Ҡ�6��5�  ����!%�QknB�I��Q$(Rr��K�od��"q��H��r ��cy<�$��W<��1Z��cu�qz��狩z�b.F��;[U��J3p��j��l1��:��ѓ��75v��Gn������{�Yӆė4���|O����ﾑ 4��"鬿��I���KeHK*&�cx��!�_U	���K䗴쿦O,�]Ѵ�}�B*E	���'\b۶Mg�U���n�k�ڙ��M�ݾԡ�)y�m%�3�TI#k��$�/WdH �O��(>ܾڢA>;Y�AS}n	�щ�]r�����^�ɗ�'�^P�O�;]�A �oc����#�{9��15���l��	���u�O��vO�� �)g0��]�A;]�H$��d���mD �	�7���t����H!L���Ȓξ���>�3��m�D��rA`����
OTn� �y}B�7��Ľݡ~$��rH$�Gd������$�{<f"��WQ=Ce-�ܺ"�Y�
q�WE_wXC}��{�� ��"�Og"|�Fj��IX�.�:�?=�p$⢐���s|G�l�ő��nq� �����-)m�Z�a���5�u,b�&�����I��_������}�ǒ�G.���޷������ǽ������ٱK��}U�Ǎ�[x��볆����aJ�I�{՚����J��d�V{�h�1����7���g#��tZ�f��J��tC�q�������~Nie`����u�}�n�v�x�<�u��t.���cތ�{G���m�(�Vlri��|���gr�Nv9�f{�����=,�v+6^�Z�BY�<�㇟�z��#x4���2�-{���YG 1�+���Jom5�tonn�=�o�f��~8��{<@�^δq�W��c>>c?r[�l���'1X��"��I�Y��s�!湑�{�1b۲�GCZX����X="�o�5W�^�J�S<�ۏ��U�� �W��J=�s<牃 �1?n�d=��1S*���6�m�NǱ�7\}� ���>��=˼ݶ�y�������љ�ˣp��.��͂{Zg<"~l�gG���-�(P�tF�׆���$6q@^�ou�I�;|:H7ɭX+^�s�y�w���.q��m��hFByw���Y@\E'u�|�m	����_�`�5��6���S���z��r��(5��{���E.ӈ��m����u�X?"��R�h�e�j"�#im�E��b*��FZZRԢ��V�*��x�m-%b�Z[J��ZҭZ��m�KklIm��V���eE�ZR�j "#Q����J�$R��.�Q���Z��QTUPPV��F"�V�h�1��UcZ�R֫�b�)T+b�ʕ���Ec[2lT-J�ձ��Q-
���E�"��Q���E+ZRԢZX�iV6�A��VYZUQ����R֨[B����-�����Z�QE+
�+X��*TX���ĵPE�,�����kEdE�Z+�sQTD�����-lUF����Ԣ��
�T-J6R�+#B��P��+,eVUX�Q�j���Q�UE
�"�B�B��jQb�iݨ���-���kdb��6�EQ�b�*��+,UX�m��PR��ܷ��۱z뮇���k�Xwƫ�s��:5��T�v�x:���pqE:xy�܅z�'����lv����Y݄��el:����y�%��gE���sK�Y�7��ݢ޻˱�����>;֚�؜�fzSCָ�:�H8���;����n.�=�X��qGBs�*�5��n�uԮv����g�h�0��M���a�6�{�Q1&8��و�V3�]]�iN��5�a܎i]�gd��K���N���f��t��g�9q	�6{�tc��kY�Լ(r��-HƳ���D��b�sky���v�����cg�Z�yvKgf����zI��F뵷kOk^�kgVS��TV��]��ݞ9��K�;�:�g��u78]�[���	\S��볎Gv{;��;&���^:���ux^�'�xR�#�Ύ@��W��]�9��	r��g�u��6>|���f�@\BwjM�d໶���{q��K�V�-ю�ˌuɲ�۳�h뗮]�N�Sj�����i�tڱ̲����|r�1�݅��۷���8�0��K��X��F��7'k��ڰN���֧�#�s�h܏Fq@;^�8���Ѷ����g�6��2�N���v�3k�G[=��]y�n|ZĎ�f$�y����g�eA����_E�9˷&:�v��98�]���q;����.��6v�f�k�nvԹL�t���[�#:��a��3mk�h�����ۮ8�}X˓��Y��I�����n���3gkez��(���8�j�F�Ŷ=nt$�y6����b��Lti$�zM��	�VZ7��@��U���۷�w���t��fԕ�X��ֻh�,�/cqÌu<"�(�����:x[����Lq�X'��Y�v6��=�N�u��ls�g���q�9�1p����`����6����>{��^��A�vѵ�g1������j_Mی�+���ۆL�s���v�]��x�\��F�cq��ڵ�n&"ҧ��8��۶�Ō�Ui��{����w&�`3����B;d��ֻn���8q�A�rUV���Gy݄�=hϰ�^�;��d�9�G�����]L�uC����@��Z�[v�.�u��㚱�u���6S�m�v1ǋɎ�p��@�F6�&�ƶ��NU���'�0:�<��r�U���8ħ]a���t
����ܪ��`���ʝ-nqݹ�m�I���ᕶ-�=B�u�!���u'n�줠��7c{b��&.[��S_�����l�F��x��>�|ocrB ��@�3f�b��b ��~�����ԡ�)y�M% ����n��=�LXK��$�řC��[I�����uV�7�q0��j&�T����޿�B_*���i$��R�M9n�>$���;�2f��M�YA6T�9���xhɫ���I���DC����$���O��Q��ʚ�v/�#�U6�h�!pMQ��٢A��|N��ƶ�(ĺV� �k�'Ă|��*�$���0$��+G6xt�gŻm��lι��v�Ys�1�n��b�y�^,�*�v�5"�l�4|�(\�wH^w��(�O���rٞFJ���d�ų��=��fk�ꒉ��.1���/���2��}�~�\��١9���12�WH2�H�Q�A��Fˍ,<���F�vD�Dv���O+�i(�zxTv�ݎf�MI��ڹ���I�<;1�����{��^$�f���'�J��v�2zS�A�^B���Aa8J"|T�uQ����$�":�Ф*�8	��^U	3}�IN�+l����2`�����3�;��|T�Ԋ"wu�$�}���؅���X0\�\�UQ3Z
A&�,��=�b����f��f�1͙ھ�@�;��A��r!��uE������<g2�����A� �s��sѐ�ks�^�=�;Ce��5�р� ��{�ޢO���r$��Vd�
��	W�D�L��N���}Є��B��Z�`��*��E�� �|g>�$�I��r�˜�s�y}}Ѱn���fbJ�`�= �+�p`�M��lMz�ro��#�~Nː��3��g���[��%c=E#j�c�+Nz`1��%�U^���p�C�Q'r���wۿ��r�ܮ`���Q�D��wM+�vz�H �8Ēs1Y�u��&ͪJx�؛ʮrHN�6-2�M�U�W"<��h
���;u�J%V�Ev+� �೯��\�O���|;|w�v��vf2�e8�cn��1ylnq�v�[��J�ۇlW�����e��PI��3�n|A;��DI+6����"-wpRTc��hʜzA=��@��UX�h�EpMQ����_N��6�F_;"I6����9-)�Kry� ��$��D(
<B���Q�!�����\��@9|�} �Vu�P&3:����� �*S��YޫJz��&Z��I[��@�L�s90��Ғ�~�����1z�3��׃Z6���:٩�^lX�&X\��Jޕݕ��[6n�eU���4������b�5��ݸ�"/ڬb�W�m��| �[�2PD��(��T�t�N}�ON>�2�E	 yNϥv��H��b#f���U���j{s��s�Y�Bl��:8�gb�^r��@��\�g���K�bA���>�6�E�ٍ��Z��%=���I+��\$��
���bջ��+#A!g_U15��!6Qe�Rg:�����e�ds�V���U��Q �7�Ę��p�b_56 �t�mD�&d� o{v��N�9 nK���ҽr&gl�$���I&o�����	0�P)�޵���N��B�9��U��7��H7ܮ��h����D[��wT!��p��U�\����y�Ȳ*�!9��^$���$}��'hގj*�D�"���kcw.��4l�2x�Ck��:aL��BFi�.�q�0��϶��MD�a��m�k)����`	��/37���
�{><z���>:��iM&u�`�n:9�`�6��L]b,�
!���g��{v��{�����s֎.�85����ݞ���]��m��]�����;�v������ۮgp�ʩ�ض{��{��#��nݪ�A�u�0�S�̻W<gR:���ݥ����"�r�����f����gOm��ˊ�O^3�6w''CX{vݐ�nV㦗pيY�g�b���Z��k&�힤7<�7�7nw��a� ��U���LR�%P��A�E߹��D��	�$�s�>5R����`}��(g{\�|��bD�i6[-��5\��t�l�5�f��m��$;�ē������v��K��^Kxҋ-�)�&�	�	0�ݧ`|�+��x8��ghs��$�;��O��+;*q��)3K&l����΋x� ��>�+�Y�Jξ���B$�V��K�I�("a�(C���	*��]Uİ�����uâN���|{5\�%f�U�:.v�ł�)���PT�i���Qml�\[� ��n"�nw��s�m���߿`��E�bpn��$�y��$���U�!Mvvp���K�� �A����<nLTLJ�U��w�m=���~�/��,��J3ƬY��sr�H�q�u�-������,g��e�׍���-�F\��e#��Y�{�}�ݢ{27��]t��I�׆A ��P�*�*�Fn:Sm�S}�)5��8����"	 ��٠F7��Eh�3��	����Y��C��Mi)M��AC
A��d�v-2�`I!m�W��w1ؽ �~2�?<��w~�?G+M��$���^��mBJ5�U�����*���}k8J�v	��H$��٠O�7[�B�s\���F��n��"`�J*)�"�gk�:;<�v�s�O�Ez�F�Ν�����s�����B��q�׊HW��^ �w9#���cٻ�\�2���m��39�"��TT&�Ʋ��$�w�8��<�m�y�A *�ڢI��r	!�WLR�}*!�n0��,H�8�!��:�~���\�4���{&yd��,�^���3*�m�����|!�ѻr�U{��_NU�)�<J�j�2w�=&�c�F�>J6.���͞�n���|n���T��PJMCe��5Ցw�*�{nC�ˑ@�<�|A=]�H"�vd��|��C"�.�P���)M��2�� �W1$�=��fp�Z8U�W$��o*�I �g1$�l�b�f/&^�"Tl0B�8�����S�p��m�auv�����ۦWt�<������I�Vb	d��ݚ�>#k���E�v)�Jb	w�����u@�kuωdm H�L�AEB���e� ��75��!UO6������r	�&��K���b����N�>D�AQ(&��g�B�,�2	=԰�vB�Bbwp|H=]�|>6{�C]�%@E�n��9�862n-Y�;(�>[��I;�����󣗖�_?˺�����<�`�λ1�8s���� ~�;9����ň~>���KE
j��V�.�-�"�˘��ٺ���d�Yc�0��y 
,����*��[r�%o^Х}Cf��W6 �v9�$�=�!�J;��pw#�[��C=S�zLku�j��1\���vh�ϫ<ֺön̵�#	0�u]�!	��T0��� �8�d�In�M�Vh�3�,O�ӝ���[M�Rf �L����Q9��<�7Gsz1�xH$*/�O�+���K������hu����H�Bn#�"�H<z�	f_MMV�����n{1�%	,Y�?\���J2sY�MQT�j�_[��z�ĉ�v�F�̩]yTI>7;�j�A��i����!r�A��-�PAO6�D�2s���ռ���iͭ0n���O�$*��E�s�`S�ZnMBPv�XwWf+�a�F�Ap���#+(�M�%�dZ�bپ7�
q�*쫉�[���N'#�G,�O������.�� ��	����u;ll���xլb^�g��<o:���r���;vp�a۫�&׍���c�?=���8��qv��ղ����9�a��1u��;8�x����4N_G+�G&:M���˼�U�7^Wx���ɻz�4�T�۝p;�g���5���EmԏJd*���$�q����tk��ym��ۮ��#�&�,;vیn�R땇r�=/=w\,7Wgm��狓��x��:2e۷l��e��WN�'A��Ͽ��l$0MÈ��4k�|�!f�Т	$��9�5�75N�r���l���9��ݽ��ZJBd#��/��AY�;�Q&�h2H*��h���I1�l�Ui]�Ϫ�km�0Rf �MQ����>��rO�;bot��Ⱦ������yy^���|vt�'�7�P����P�fJ����Fn�PI$��9'ě=�i�_T�w0���>ŻQ��7����W��E���6ˑ�%V�Q ���$�g�d���È��y{O1˲r�NnN�c�m�J�r��˶�-��a"i<��A��d�A<�|H#g9�>'ċ��Aa�O�Dq�f�=}� ��~{�U��,% ���d��\��P��wYҩ�	r���s;ou�2q�Wrm���3�"f�J�웉�y;:z.�-Ƭ治)ڙ%C(✺ݜ��T�ܬ�@�:{\�A =�,���7��r(���j�HBl��C��	� =��ĂVJnN��X$A���ĀI�ݓ�v9[l�BLe�w�b�_{�}]�I7/��FF�)�>+kziM�}0�^@f�<���rI��H�&Ï!B��oe�H++:�]�"�5ћ���A��rIo�X>+kzh�P0nL
0�T��c�t�p�����qٝ�A��:�fq�oC��I���J����Bn�~PT��b@$����A][�G5b�w۬�Z�|O����/����%�
�y]B�������u1 �9ؤ����Q�q����s�׌��e�KLCp�&�h�ܰ@/���Dxzl\�xPCm�՗u9�<x��CCc��!w��㧛�O�f�&]�&�ԇ9=�q��褗�h�vA�|��In�
ւgugrg}=fQ�z�/+�'���f�8v>�Σ�G0��gM���!��ƬY�û���C<�ud�2��y�X=���]O�=���'u���P���Yû��v�JE�K�W ��|
L���o��vb�5kۼ'z9v�0 Y�SB0ɼN*��ʏ �f�d��,�;P�h=�<��5�m֤��=��G�p'����8l����ĳ{T��۽�+�8	����p��m�e�y�]}�w��%�=�}��a�͙��֩�U9�<�T�S�;s�WĎF/&sr���'
>�("�ט��@zfǛ� ǣ�s$�T���֤���۝�?:V���n��J�4p�C	�����v�m��7ݲ�jq�տ�tq�M;m�R��z�y���Oa�'V�T�E�P�)oѿ-���s'b�{��M�{P]�f~�\��~j�%�����^�;��@�h�b����� ~ܑ���d����î�^�$nf�l{4���[ֈ��6;�+�ݹ-x���O5�.������lt������L�!T��<ǫ�!����p��E�^��7s�:�>��p|� ��0�lg�s7{�PI{����p��\4Ku��d*�n�N����ʬ�|:���v
}�O�,t���Oe0[�LUf��P�&��}굑yv��5���ܭ��W�6@�m�TjQE�tتf)ֶ�YF�b�����bݮ(�4kZ"1V(ڴIX�F�5t��h����kKh��m��T+F�S03�,*��Q�Qm��e�m*V6��l
u3���Ueu��XV��� ���eT�ia�K���.*��YJ�`,"�W5-m+lPEV��m�dXQ-�Kj��Ҷ�ҵJ�-����Q)�������B�F�F�\�5��u�TkJ!U(�[Z�2T�5�%�Դ���m�҂�P�t�R��U�Ur"6�%�PR�Ū�Lݵ+�V�R"E*V6�#JVLͭDIj�X��Q`�VV��� �Ѿ��V�W�Q5ĤmSFRr���m����-�(mG�2S�>'��oH�E��+hng^� ==!�U9�ۄ`�Y5F�7j�k�rfm,�Sg�`��	%�f�I6����LM����l�Ap�����MÄ��[��h�m�î޸z��Y�5\�,,o߿��뷚<��x�t�I�/+6k���m�9/#J���Ye�T�?L\%�7��Y9�?�-��D)��߀��[��~�̂���D[�b|w.��^��c`�C��R�q�(b<�p�Pdɭ�DA�|O���SmE@�[ҰHs��^$|m�9�Y|���ᨪ��fr�;�3�q�I;�U4	$��r��e�`^Β��D	&o�ſ�zx��N�~�c��e�'J�q�~,5��^Ǟ���}{�Go77n,3t]t���;����1���\׊.���M�Jh�=z���q�4x틺w�k{z�Ē]�����q�֖�|�x*���R��kF������n���n�X�!�� ����c��ͶP!,d ���o�hQ>[��	�j�7�I��s̡^$��AXi�,� �Rv��|��z��e����A>���A ���5b��Gpޔ��N-�?�)��D)������Հy�w�N觡!~y���9�V�B�;�/�ƘP���p�Pd5�)[�qH>��bA }�̂�ޢm��{�'?��tz����ea+Oe� ����O���T�;�ě�6�/AΘ�:�\���P+w�ț27���]�'��zon#_{gx�"���y��B��3-ʭ���*&I�����Y�z�9���>ej�ԏ)�N��v�����;��b8l��Y��#�Gn<��۞��;;n�C͝�s�5���j�>+�=6ݓ�$ �Ɏy�G���l��X�7o�8�lQn��ջv�x�ޥ�h�����&NiJ�Fh�j�c����Y�;��M���B`��l]�Űy+;�5lH�Ļ]��eݎ�=��u\��7Wj�l�q���"�<�{xq�]r��݄.2�&s�X�5lny��ˊu;v����a!0�� �D��1[y��mSF\gg\�HoU�O��ޡ���,����kH9x�}u9�ۄ`�Y4.��hv�*��¨W!��S�I$���> �=�B�Ί�6�H�d<�y�NΙD�&H*���d@ ����ME�Ĕ#{T˧d۫$@$���H.��SE2�b�K?7���i$R� �52�C�̪$�{��"w+7B�Ho�ڣ(pHL����d�У�H����Ց7t`�)�$�s� �\�mP�-�9���MM����.��E��瞏i㶷g�t�8{��]��ㆳ���K�HD4K[y��!���n[��]��>!��P|H$��a���T��)5o�|��L���x[x�h�pt�rC�7UW:��'M̧������u�Ql@Zֺ��y��3/\�z��C�cWːS;�4TI#܂y���qdQ�Wg�\q�\���	k2�|��䍜��h� ��;���D���I)�MW���Т��9�	ؘt��|YW�Um��%�gME��>$lN`��f��6yk��C4�bI/&ꨂ:�\�Fo,�ù�nj�H�D�WU�o��I8pAAP��x$��r�Dn��3�7TI>8�A �r��� m�T�#)&�ŻH\���z:�vo3�f�	��U�9���j~pg�+֯_�}��:�T�=u���o����U5� �Nw< �V��d��D�d�UxM��$�]��l�Tj�\�>56�̃Zv����D	<�����$@>=�(���\���x���l&�Q�/]��A�œEf�J8�I���T��ԇ)u37V��d߱Y���Tp�[��}�l�?su5��H5ֶ��U|���/+�WF]��m�yR0S�<	$}�|I&��O��m;��HDB������V�ç ���A>'���B�ޣa��\e@�E���y�N�L!7��T)v֙$���=N.��}]���˵�'ă��$G����1��~9������gr!8a�MYk����Y�[u�nLnjD�[��g4���~����`PY����>��s�$�|�o��i��Wz�&2vx��������^v�%C�Be��|a�t�.��(�BʐzE[�|H5ج�>/v�hp�t\��ާ��Y�!	��eU]j�/��GĒ*�jn^ڶ��	7ڮ} �K��fk���m��l�����u�P;ĀW5�	u׵D�Iw���yt���^��}u����>�J羚xA���<x7�ܖ�ő!��ƨG^�9���q���n�=���e��'a�r����Cz�MT��J����e1�[.���H��Ft�m%��Y�۳D����;w�t��Vbg	ŏ��	{��@�K��%����I�Ӝ<b� ����txt=�ɞl])�dgǎ̓pv�9���`'�zu�D&���&u_$��{^��I ��r]#��Y66L࡯�h�I6���'`�I8pAAU��>$;�V��e�W"$�{}TH���r	g��ݸxf�VxA��%DC$��DSκ'�3��H��컎���q
�v[<	��H�|]�9'�vcHBD�d��U@�Z��h�L�T�٠O�y���M�+����8�8|c�ꨐ�jʆ�m��l� �O9$��W0j�;�=�
���$��5��W"prMX��\�UL>��c:�M�Mר�����T����=q49��+�S9�2v���a�~�<F�u����w�}�Į��ϰ���I���0X%�n,���[��v�>�#ՙ�����oT��U�=�zx��ׇ��6�������.���I=vݮ*����s�(0p�#��|�ٻg���'V��/Є�D�iw{v��1llc���yz���˞�;];���Tq��lPm�ƋHmU$z��Ž=����X:���':�:��`ݼݙ�sΰI\��<�i�:�.�6wb6]��ۋJۭ��r{b�ۖWt�G������P�"pApk����A$=�r	${��������U[ݕD�H.����lS�m�DB*���L�rOu�轜�cy��^�9�{�Ȑo�]uON8��k'��I����7}lO�7ڮ`��5����s�� �_o1 �{��A󄘈�IM4�Q�s��}��<`FW[�A$�c� �O���6�V`Z��z`������p,���M0��>��$����_b<.��E�i+ulH��W0$=���,�(f��c���g�prZ�[թ��v���.Ź)��&��Ŷ�������������Wh�Y��5<�ĂO^���ݾ�1F'�\ٗ\ĀI��s�N�	�I���7ݻ#���r���Xu�e2V��,\)���kA&����0Z��.D���rt�H=!���U�?.�@C/kg�w�T+�z.S�xҺJpk�|	�vD�C��T�l	an̘�tM�X�	���T)�V��$���ȇB�p�f^��I��s!��UF,���M�����ot�J�^g1L��C˾�@�]�3��٩�հm��f��!���)��%@)��	3��z�o5:�]׉i�2$��}U�I��_�7|re84���a���p���T�u�vb�m�Oln�n|"!u��S��0�M&]q��r �Kͼ�@��%L+�A����2���DЄPH%��]�d�6�b��^.�$����*�${�I ³�P�3�Λux[��P$���Ȑ_��m|B�� �#�������ܵ�Bֵ����r����^L�n�wm��}-@p�c�s�'���N���<�cy*�S�+22�x�U�W�$}�I���#�!��R��8vĪ�Z����f�A��y-J��W�2D�G��:��Y[)6�i@(*�w��	��r"Z�1�=xJ[}^��5���򹆧�Wr�h�<�F��7�����8���Cv��Z.�����piκ:a��a"!���q�0���H�����-�rI>'7�����YjRf����	�%f�z^�n
@�e4�s@�W>��kQt�zd�ؚ��
>$
��$�W>�A�1%���n�P��jm�&�)ry�$v�\�ĝ�t\&n�=y�7d�Vg9���A�wUT��B�7���_���_�&���� ��Og;>�=�N��4���j�y�e+�g�H@g��PGũ�C�vC4~\��ޔ���.u��r��O�[S�����m��ߑN��p �{�@·�E�L6D"�O�W-�A!�gK9�aq����$���$�w�ȐO���9�1��k�]�0�,�b!�f0\�˽V;5�Bdnv�n��-ӑ]��>�a6�i PR*��x�O����Q�5�^e�I��Y�H'w�Ȃ�	1�iTI����d�tR�n��{������
���;;;����$\��؄���8NQ��fHsݔ(��T�D����I^�|Hwz����jM�mCN���wti5`��v�l�'���7j�${��ߗ~v��s%W�����!BL�P7y�"�{��껩Kj��ɟ@.{rhJ��;��(��7Q!�Fj�ql�S֑�j��J��}�qz�����݊�}���o������7���Nz�Ҵ���=�WQ���G�{�E�徱�l��M�m���\��ק#7.v�_��	�����E."x�����G]��E���n޾5{�)|g�T�-x�{s����a����zH�Z�&�:�W
��g�Z��Y���`���lҤ��7�<���oٺ-pɽ�nk��pE�}�*�-=�i�m�9T�Gp������?h�X�8:��Mw��K��<�wW����td�7ց���E��G���8)p3>�[5�h��p�����lsZ������]F������H{�$ҹͮ{����3\��Y��)��K�@<u��{\������x������y6�?�7���M��m=<b��EvnU��Bg2�D���#���=��������}�:y4�lh�s�3��˳�/O�
��-V�.uP�)�n1�0�1�:�R8R%�9�OzΧa7�V[z#�}`���;�]F�rۏ�{X/Jrj�-|��K�K)׽��Q�K>�Ey�a����;��A���Y�CK���C�:� C��aUu�>�==�������x��|8%�x.o�$Ƅ�ټ8aj�~��6��;��v������]ٱ���{��E�b�=�rm;�y�.*{ǩ.%|�b��]�W�r���K�Y3��D�:��C��4��{R�:���;��9���<�\�AE�L�%�km�V�Gc�f
t=38�J�k.*�s�]j��kb�D�e����)�m��ҩj����֖�9,�lku���qG--���eC#lD�!u��u]I��ڬ̍�3Z���;�=�s�=��=����Q��W2�Z"��j���`ڎ�s�FT��2�l(m�y|8���>�wvJ��k���GQr�S"b�71r�#v�NzZ^��96M��:��fQ�S6W	�c�.�5B�n�U�:�#qAM�ڍ�ZR���TVd,sDb���eL֫���U�v�¨��{��foA�nC9Ej��rIDU�T(�D(Ԩ�ؖ�aR��TZm��F��G]������J\��2�9+PP\�ef�U3qUs�V�5����.{��y�q�u�Dz6T�K���^Gi9������v��������;��j�M˜�����k����S[]���:k;x9۪ί8+�rq��vD�a�]����Q�Ŷ�<�n�6݊z�*���f�ӵ���n����+ϛ��s���wn`��1n�׃q������kNg�i�hu�.8Ɯ(��Cm>IF�뮳]����ݳ{j��b3�rź��n#�M�]7`�!����nԻ= ��r���]�yl,�k�k�����^���\�y��[i�(ug# ]s�����s�,�c3qJs��g������s]�l�B��`�㝠��ݧ�ot�U�(�S����ې�vm���fvq���\cq����x.��uĜ7	z_C�:�2��omvӜ�<��l�h�"�hܙ���r�Msg�s���Ǟ��qίs���8�8}��� ���1�v���s�۞�9�o뎎�X�p�f�9�Ÿ�ݎ�լ[<��s�=��Biwn��qzM���s���x�4Ӷ2Zz�v���>�"�p�7U�'����R��^���)k�(u��+��p�;s�lB�y�[t��D�n�6�^7v��<n�q��m��㣼욣�cp�x�(�bݞ�N0�ܮ2�#���c�9�m�[h���8�+:��m(OV��ׯGg�$q�(��`�Mɧ� 	��s�<����񧉗k΀{
l��nwa��-�c�q�6rv�{��y��AF��\���б�ۜ�u[Or\��ס]�m�n�rrh����X�sюN�&�{m���8��n�k��n.�����3��8)g��\ltrN�2\s�5�ח>ۇQ�ѰNԶ�{3�b�vt6砎�۲��.��
�97F��^�r�=8����u[���;Ob�)�f��S/a�]�l̦S�'�ڂsx�^��1�k�(�n7j�y��4����j�M�c���'��ł9��wN����p�6zʼbI��sF�Bۄ�B�uUM�g�g��9��q��������N��3�uA/ ��tN:ۉ;��덢{/�w2lD<��5�מ8�P��rF�n^�`7��jNh\���ݹ�ϝ.�t�V8Ź���EF�����%#�����gG)�v<v鞮7G]^��l�g.���X���ݸ��>�����wl{[��ē�hC���#յ�Q^y�c�=�3�ѣa���8�ձ�����m+�љ��Lѫ�t���vѲg���?z�5	�ȄT.��'��D�|U�91R�O�L�:�d��=�T	�wB��-��,R|-�^����{���4)����\�mP>W�Ğ�re(긫�q�L�Y�LA���@����� ���O�N)�/��򨭣���u
$��b|:]�l$�M�p�:�=j�J�̚�����MU|I]����s+�DH��?0�]?Y& �뉢�6Ci�Ґgz��	;|�DF��<��'���wgUY�ĀFo+�F������=��$ �`��!0�(�[lpn3��\g�fހnE.�����?f2X��9����z�$�yω�'7�� �t#��N3Q��u"�!gk�vX~M$�dB*��� ��;;�2s��fyd��,$���ԇ�䟹�j���L�:��գ���
eu��9+����h�M���_�Y6�F.��ɝ͒QB��;���A>*���O�o+"A�7��c�F��M�MB

�u<�M������vm���9�No/+�y�`��%%%�-�3=�����ҁ ����A#7�$�=�Qcؾ�����5\�*g�6A&�P�*�U�$�&�䤞nL��<ĂA��s>s��C�*9��ò.������7�v���0GJ|��nV��"uc�(C)����&���	�	����9>��s ���Q��_Of���/@$�y���z�i��AI���uݓ��d�sV���vI$��vd}�|�w�� ���.pwL>X�EB�"�&"P��+���>�gUA��WI��RȞn�.*�Z�%�{ۄKٍ�zM\s�S��o�|��<������/����"��:�n�cgyA��ު�b��wv�I��s.{z�s��m�� ��S�TW[J�
��B"*V�$��٢I_sr���W
bs)k�w(�̋�
!MJR���D����Mٝ�ј���2V9�ɢI�s��l�m�_I.gȘ�h#( m��kv{�96܀�F��81��v]9���~�����I�p�p��9j�=�T|H!��a��3Uw�L��hPp���,�Zp�A�K���t��Q�+w��pI�;}TI!��)M�轲����l�d"HI�Ao��`��R �s�l�B9�͂@%�fP�|����+,0�P�~p�B���f)ԇS�M�I��SD��v�$���n�CI���ީ���
Jv4e���1�4�#�dJ�1tz��]!�};�	՞yu�-Hi��� �-��%��h����7�QM�ے8��{�@�w3}�i��X�Rq��� �yQ�g���ɩ�Iq}�I�'7�ϣT�����ޯ{�Q�a ��x��V��td��� ���3���s[9O�˵?9��8�k������vuJ�S;�gwT�A���=�t`b#-(�J�(P��ROLކ�aCIê�s� ���g.�^���2�@q��O���s�o)�
��4DWj�I�yaL�R-8m)��m�I.e��P[ڞ�$&3�	�������H!LВ�������8Q�_D� ɺ� �H'{]�>%�wW{�hf�w���R	�Ya�ZI�C�b��[0A ������ɣ�X'����	�=z��'�+z����Pf$��A���N.�`m��m�J�A}���L�������{���z�^�ӏ&�f��}��3e�^p��L��nQ"�x"�����w�V^�M������k��ZCW\)��'$��6�ފ�t)�Lp��^�)�'[[��F9�z�19�M�D,^�g����\��ۤ��Dn]��qbunCϮ�:���xlf�
n�Sa�cL=:�E=����&�o��z��^��>s�v�7���彄{qe�&��7]����d�"�l�����L���rqi�g����v��Ɲ�ѣCwm�\�[�@(�ig�+��q:���.�[�ۤ6.6h??>�G3H��������R	$�� �Hy]�F���w��웒����0w�P�~�I%�	�PD�§+��*!��m���,�$N�;2C�ޚ��	CE_6���Yۋ�����#�6Ie2��oꮑ��� �o���v�s��A��s �򷪁3l!?4�nJf3�n\
��N��M���5+$G����&/yvIʈ���f��Js�pk�tQ(�L��+p���4	2wy	�j4�8#U;VX&/�� �U�Q ɽ�*'ν�L���$���m���a��FrKٰ=����C�<v{]�Y�h�N�G0JP�$8F!q���ݚ �_rŕ/�� z�ɀHv~���� ��A2����g��xz
�*�L\=y�Ϊr������x^!G��۴\1}�B:��5�އ�c�bt+xL��Ov��3��m��t��Yn�Q*��'9h�� f9=�D��1{�@"����䊭�rK��d�j'Q|T��
$�';T�	�oi���.s�F�	+����f/�H=����-<%��كZ��$���͖1|j���D�O�;5I޶"�'����ۗ4H�[aL���&��c:ԒO��[�o�[�H�{;�$Fo]P�&/�H$sz�V�8q2��S~���`���K]ᱶ!r��ݶg3�9�wKq�,��*)&+wuÄ`AI��\s�:�L��RA'ٽr$�]��u"/Gv^��캢���$��fX%(M�#��k�7�#Sq4N]F9ˡ@���BA'7��bQ5l3ǱM�'\�W%P�*����I �m�$�h��W�R�뿨Ѽpon�}9y.�p��^�n޾�n�Z1�낰2��H���GVA����g[�R��%Z=F*[׃����sP�	7��%�i��)���>*s��CqH���!��El�h	�}$��kv%�թ��h;ԅ��
�Å	Ü �]��@/j����
�ٵ�nZ�H��r��ު=w��x�&9fX��D�BjH�	d'�Wl�R5���3���Y���3�b7��n^����x�m�ip��� �^�	%�wUq�L�D�\#��I;�n|H�VM8p�)1 �j��gU��5;�g4ٽ�@�H�uϤC�ުo���T��cmq찥�aBL��'k��$�u�TA>ޖ٘o!�TH'��e� ����T	�Ej)���\�:Vu��+��0�3.ܒ	��$�W��dN��2g�Yٛ�������'2�؆�53Tn���A㼝�7���u6WIu�^��b�ɽ�6���ݼ�L��;r.:�Kw�I}�$�D�H�� �ͺ�}9��}{Sy� M��$�o��$f����y5�uF�Ky�Ё%''&��A��	�{$v���N7#�v�.�y�9�t��~����QL�p끞�s�H��{U��f���+q'/$�s ��9��.�J[b&Ii
J|g:܂@9�&o������8K���$�f�������6e�{�uո���P8BO��_N���bHw-S�����tĀH'�����|f���6�9`�P��!��n�n��8v����Hu}�G���=��ē�{��(�;8��}�����K��F,�`*S��'�^)jUF-�@f�_���9xm��L�6���۠��Xɖ�7^ꛝ�@�׾��nfդTA���8x��c�Ɯ�4}"��Y&�,��"��ѝ���#C���׵��מ���>�&퓞l�J��}���fݹ�����i;v,m�.�B2C�:�]--Ƿ4Y@'�w'n}b�-y4WY���i{[����dCŝ���oK��i��nz���٭�ny6Ɨ4o;�ܜ&�l^n�m��v�<�_�<Y�vl�b�5!�n^sxǒ�9#��T�J�Ҭ�lq��{{vꠝ�ѩ5�x��������Q[�����WU`1���];8����� �Q��* �{9=�H��s�	&��D�ckqJ1�W�s��A��rJ��	��)�ч��]������y��݊���f�'ă[��OZy[���+$d&�4L
��p� �^��)�A��rI&��7޽�U�R���$�;��	����r��1�@,������DZ�U1����$<H�ʑ$��A�Sq�6 �s�X�Ya�� �
|z��I �nH6�=*��9I��O�vӐA�vH���֜����~v��őۮ�2�CWnpS�Fr�;��e�mㄌ/x�E��w�"HE��٬I��$�y�����Gi[LI ��9$:��A��j�C�ےf�<:�C�*�XF^�,�HJ5�緂�����.��*V����y�,�ۏ��U@,���l�q�{��򼫞d����4&^=�$��u1 �O��'ʵ�*:�;bs_x��	��	��jQ{v�A'o�d��v779�����rA ���2��!2KA5�R��w8:&�nge����H9�.H>$V�L�I�u�wp����u��3Z��e�(�@���&ֽˋIB��uZ���,K��h�w�u�ݖ���s����s���u���\�t5�&�ݴ.t�lꋴ�Ҧ��7;h�3�}�~w�ی"��.���� ��L�Iz��*&8�[��_k�A$��Ꝕb*8
���$".Ʊ��� �W�3�@$�_9� �=ǲkof��^_	�ZF�!D�u�'�On9$~3ۚ�~�����Z�6Zmx߸/B���V%4vG��h��riCX>�W���Ac^��)q���vu�Sҧ�Vyv���w5s��{A>�Q-���UB�� }��g{m��9�5QJ�6�1����f�zWǬ�����i�ڍrv/��oB_,2	�E�n��{�n�g@������淪Z� a�5ۻ��ĵ��t�g��Rp��/@����S=���$9�{��M�7�Z�����gԻ��=p���2�l"�e��Ԓwy�"}0�.yg��[0���vr�BՠyI�w)2�=�پ�%$pZ��{J:Ӷ�m�1����'��|u�[�oxV!<�Y�.����w���;Wzs���q5�t �y�\i�`�ｊ��1{n����_91���. ���)�[>�7s�^zA�6}�p9+�p��8�.��G�gD�'y�}7�i�����g����Ј��sE�oݳc��{@��� ��z������C��n�s�]'=����U/N���;sӚ~0�:��bo���O���3����y툟L�nh��o�o������z�@��)V~6�_�ڶ��r��S���q\�ZX�4�����n����kN�c��X׈8s�;�ȳ��i���3r,�U���;g>�:U$u{����ƶ`���AL�K[��^�=F�$>�{_�{�*�e��4�z0}<�}=��v�y �������4�r=�D����f����,�Gv�h*�J1��<���W��FZȦa��H��.�k��j��uJ�u�䢎J��m�F�Q�P�e�kY\Th�4j�J�V��M�Tι¶�Q��F�h��l�](�(���]U�6[nV&�V�R�D�ݫ.�U0Ѵ�-ˍ�]wI��բTL]��J��U#hܚ�:�˙[��X�J#�.�[�V����l銰�*릒TQj�Q���M���uN���E���8��͆l[CZ�덭��1n�cj�AYR��lVX�%B��j��1�.ڜQ���ݽ��Y�l�{����Z�L]t�ʊcJ+�յEM���Q��G[0�mmc3D�-Kil��k
f�kLҌ��V�(+v�-��"���u��-YQX�,��Ֆ��ԮiKkMviP�ڙ�(�Z���Vֹ��Tp�\�:�b�iKae,Kf�E-h��m����gV�kG!TE�-U��no_��{;���Â�v��[;�4� �eCP�}v��uk�0��E���A'�z��$��u96��E���yCI�v��2�@��фېg6ܒH9}Lb��p�F��̃�$+����su�$MwSV2�b�n��v�ݙ��u���ۋ���ϵ�^�������d!%	ݛ�#
l�,�;|�Iy�|H�+��I<��F������L��g;\��؃
`�"������_Rg2*��h�	 �f��I5�NA������óS�t97((�8,�`*��M��	Nb)�؎��AY�@$kz�����ZD����V���<f׭[�˘JK��X$�ީ�}��:��OWV�L�K�Ÿ9�zy���%#ȩ�;�]FE\��6Q»��Z�m yh��xd����ĉڑz�HTA3�p�
ۖ$.�؛gE����k�0���6P����뗻��� �o2��A9����+���"��~�"���u�;Q�������r�n��Tv�^������oN�w����L��M��۟�@;{NH �v9�����<dO&��O��ӟ%αԪ��jh��M�}�jrr���;��`�z_ I$���}��2I��s�s6�ws���>ͱ2��CD3����5ے$�WW7Q�'���5]Us���u9H��5=(����`�T1�<���Xv����� �|s��I��y;���=��'C5��I��(���p�3�������Z�7��$���2I ��1e�?��G���N9�>bu��/͇����)f^����E{[̋O˰��ov�p��3��u
n�e^�ǣ24�l�����ۈ��Z���R�����:��7.��3,u�1�ۮU��`J�k�v����� ��l�M����d��K���74k(p\:�k�6�yĈ����|m��6V�k��;�x��v_'H1�1"^�����x�{&w8��]���x��c�X� ��7O���G�l�ܩ�č�3�G�;Y2Q�3��$�;lx����T7s�������kv�3�wnv�x]��v;p�'��~��&_��Cd!�P�=
���I��$@"v��+�n�1uQ@��>>#3�d1�"`��h�����L��_qUM)�Ǉ�U�L��I��s�|-�9�b���;i�4Z�	4�����>�&�A$ݰ���=�v6�M�$6�&|Az�Ϗe�lAJ00�	[���t,����W3�i�n{����$�=����n:gvѣ�F�^�b|���(.Tro\��A��rR�SW�/��ܼ�NrdO���&���}��%+��бY�D���	�x��/N���9ve9�f杻1�=��]��-Au��y��0�L��g�$I� ���$�[�ăf��#b*���A$Nw=w��Kc��e�7��p1�A����bS�X�\��FI,hU�?c���w\n���?0��ء���/�f?No�o���>��K���nvf����{W��'V�OI��;�ĀI��r�ě��U��_�kxD��$۟��> ��$�.M���63(@$��>>��rOS�h�i�%��k�Fea(���$����I#/*}$����7�D���%\˟k(L�(P��!�X�	񮽙{������w�|{�\�	���rA�{}2V�h��,��;�3I��D2��գ
�=��qV��{e�]�Oj�=��l�?>�����`�XV�� �ͧ ���WM]��Q{lېH'�w)��#�a�ACP�e(!�U� ƨc���UOPT�� �3��H$�o9$��$r�i�TN�ER�Q!E6����(J�u�$�x.8s��ސ{�Y�B��̪�]k�	�٦�b{��������(j�/��Հ�.�����jMtx��plk}TF{�(h�5�Ե�}8{����ӐA�"�d�	KpD��$ېzv�"J��z�:+�X#35�$ evO���[|��ǂL1��f�S�h�	�K�4r�@��b���3��`��܉ �@�̙�H=W�MtB��Ê\�i?I/lvcX2f�:�.��av�Lv2]����ؓΜ��E�h�b
)�f!p5׮@$j�dH$��|仍]�\c�	������j�Dƨ��2������RI!h��Oi��ެ��>7W�$��> �-aOo���Op�%���h�J��ْ	=Q�	�Y�0Юv��X$�6^�>�_�p�����@�ZD��]lw�w���j�ĂNM��$���H$�c�V��ܩ��X)u��n�#�k�l���wc�}���K�s,B��Y����O��є�;��Ni�#)���ӎJ76�����B	��nGJۉ$㽔�,Fb�@��':�I3�:'��H9�NN��ɻJ+�����_��:���
Ck�������<��[v+���١��㶙�g+w�����t��LIb��� �f�6$f�H�i���;�2O��[� �\��(�X"!��'z�� �5YI`�ʔ4�H&h�_�;�}hH�S��҈��i �K,�d��'ěΧ �O�k��o+�H>���A ����5ޅ$�H�\%<�+JKq]6#΂Z�'�ݵ"A$�wN��F�
k)P&�^%m�A�i4�:�f�܃��S���&��7x�Ap�x��>$�e9��+zdW�n���V՞
�k+q�J�s���|ޫF����{_*l�R��ߛ'�U�j��~q>̝�g^�_��v�n9@�Ⱦ�s��o�d���bH�q�x;;7/N���\��j��K`��)�^z���(��f��3��]��Y�q�v��g�.�l�-���[v�F�[�n �Mƺe{H��ٷ$[X�ڏ�v�����m6��kG6m-v��.�5�y�2������Cy3�۰;��v۶��׌�jz�9(�m�������O���Y�rc��ۚ�'	a��gs�v����q����ݸ�S�a�9��-ۧsQ��8[��;�Cj 6P�o����{r���I��6�lf�vOm�+����� 6�[E�H6�d�*�ھ��CL@913 H�� �O�/�����`�.^��Ӽ�6E"��)v�� ��w6�Y�t���h���zbIB{ήח�4"��&5@iC(��e+裓7��N����:��$�v{��I[�q#�Ȟ�Y΋+�:�&wi�>�x��M"�p���y�5�����{]g�z�Ċ޹	�����2j�H<LƆ������߾��'X�n�gs#�$fxF���8ܨ��u�rvM�M~����x����/��f�ܒO����d���
F��<�5�=ۯ��@���%.�ڈ��$�G6���j���H��ʭ)sdn(�ΰ�Q���ݘ=޿��
۾���w��6~g���;Y��Y�x��=�%+K�^U؋1���E��$�6�6������RG=��=Z�bԱ;O��	B�Nb����I2k9I �N���t�܅�FfD�A gnuQLU�G[�,"�E�"�RWc��*�9#m��%��+�j�O� ��>W3�8Ll=;~>��:�/a;�i$Q%!"*��6��7�N@3kqP8���uwu@�d�b�H��rVì�;}h��Ő�B%�eWj�ۖ']�u]���
f�;&c��#gAm���ZKA4�E�Px��D�5��	 �{�>gjF:��]UwU H#L�ZvO��KI�C/q���h�s;�ں����/���	tٳ����K��6�a�	6���m��$���9 �GVzƷ�j�]N�B���EK3�xR�V;�C�5�+�C���#�իDJw��<�~���tW5��ѣ5w�/b�u�z���j�O�������ӄ��M��u���1|�@\_i`�.朒	�)��E��U��EML�m.+Ĝ��>��r_�BE�"�Rv��O��gK���nb��U0�1��	{)�>"�s��-��f{l�m@�8�C�@``zk�m�=�p����g��ݱ�N����>��͏԰�DEMk� ��9��{��G�s���S�O{�p`z=��L�i��Q�}��$���j vU`�\��I"�jD�@$^�uP$ѝʧ�4��1k�V�Q"�.P3�nI"�s�
�fLOA0�hd]��$�����Ϊ��6��4�m��M�꼳h�8I���ĂA"�s��$��u��W�����I����iuS ��]N���#�=;��/?o�esV�7�Ŝ��U�]���I���+W|ok\��tӄ�2�&�bk���P�|�9���\A/-��D����	�"�3��$W�LL���\"�w�@e���|�D0�PCm�8X�v�u�;�R����5��vvz������y�n�l�Ā{�:�D�H�s���q�:���[�M}���i����R	�"�d�<m�n�3�n�MHSsSϼH���Ϊ$Au��u����B��x��
I�SH���7��=@:�r	$}*�l*�E���/��tIk9�ûa��%� 7�o��S?h��d$��t�|f���E�S����*������J�Ff
nI6��r	������o*xO�%Ϟ��E��{��B���$�	'� B��P$�	%H@��	!I�`$�	'� IO��$ I?�H@����$��	!I�`$�	'�IJ��$�H@��	!I�p$�	'�@�$��H@��	!I� IO IO��PVI��b�*B�'�v` �������s�qTJ)@P (	 �
 �  �T�@
( (P���
(QT�@
@U
U   �0  ���iZEJ�mB�Z��
PJKg��)P)v:�tҝQ��d�UEQ
ֈ�QI�RIkkQEQZҐl+&� Յ�                                     � U        ��[�ޮ�5痹[��oW�����׷�һ^ �6suu�^c���W��m���ұ� ��w3�5T�ҧ�T�*ZkC�   k��m�Z%� ݚ+��f�\��,��P�N�K{� {ݏNy�UE1{�ͪ/L�Z���X�k*[i�            {�D�iv4}�:W�K����sͥ=��� ��0r��M�t��(R�U'�M*�Ѫ�� �(P���k4(��dS��H�mU%�   R����S��P�K��  �Jc^�*q5B��,����U*�.�� /
UR�e��(U�4�����(��� �]⦆��)��  �        �B�s�׶������R�s���� �tdn����8��}er����� �.��Urлc�l�-����  .W��a��4$+ bB�j�2j�����g�<� � �(�j Ue�1�4�Y�&�o QR�m���           >�^�0��P�#��c����׹y��ҷ� �����������<���=���k� ��i��7z�^!�=&��R�|  ޣ����!�C�< � ��MS�a��qv�iBsm�4:Z�� o zna��*�9�\�Oa��C��1���N��  |        (=��2�n�� s�.a�x�\��h8 :�`�b�:��=�z޲�;�!U�p 8uOox��֚\�t�pE�J$��|  }7��q��ެ�6����� �����l�];˸���-��y��J�� ���\�<��o-\�wP�5馍�8uv�| ��h
J��M  O�bJUM4�&CO�4��M4�Ob�Q������=�'��T� �J=5JJ �)������k�_�������Xy_���Q�Y�n����$�	����$̄ ���$��	!I��$�	"B		��|���gXq�^c���f�pc?����R)bؖN\,���j�d��.���w��C7l�raӻ�m�+�f����I���xwL�&���8�c�բ��!y8=Z��Հ;�Y���1�rV-*�]���X;�딱���VS��Ҿ|��w~�q{��d�6�D@�ŅشQt���\�$;����l��K��_1e�&=��\FB�k��.�ڷ{�YI3��\r�5���0kj��ٖw�ҩwn�K8�gT�G)��7�$��{H����;�I��5�2��I��՞�eל̏�R�w�`��-��E�q�s����M����)��Vn2	QKI
N3co.%�j������x��GŪ�&����K��*��Az�q)-�WҖ��a�gLEa4���]�X��+Y�RhN��J<Ҷ��^ ���r1�
�3fO�,(��r�'����l��A��P�u�č:�=���S�޸BYm`M���œ���^v�'��5w`/�n.�{DQv������H�goR�l�af�Y!�N`�)��Y�t`����o$�ul,KϧPF����nX-DE0gB��JP��L����m*�x�+����`N��C�s��փk�:�m��Im�w���}y���t#��8S�kh��k������ӗ��C��X�E��\'NhMG�ŝ�����ƻ���e��P�fpG5��e���\��Gby9t]�֗���5g=vܸ�����Bq[y)ǝtdw��"�k +$�K�������V���@7��Qs�ڜ�+��9E�u"�*L���n-}�a��F�x�&WS#Ь	�{��m�Y۹P���"f���u�Y��W\���El%ړ�+�.u��4����|�-�Q��H�Ϗ%�n�=b\�D^<�{�u�saB�eb�����n�1��[h��FvԷ2����I�;�5�ҳxۜ�:�-ԩ�x�0w��g6�v�_�]��9(y���|��oܛ�Dg"�0e7�N'�@q��N�1U[�ĲW)�'ь�e�ϖC��n4�c���㣠��e���ք���K8W�\�p5],��S�I�;0OH�N��&�=0p� �r9)��iޝ�����إ�O}�΍j�{�)�wP#.k����5%#/T�$	�r���W�n��X8C"L?]W�v�Z}�G4���ݲ��d[��{1��i�Wii��c\l�X�m$��t�7�$]��P޽*�	n���������x�-*�(Rv.\B���;ؔwBT�3(���ՙ>9ϴdU��Ś �o<��`�0 ���c��5Ը��z=�}qqv�p�� ���L�*�2N�i%}���p������q=�t�L�ND���6n\lS' ��%���R�wSL���t�r!�b�B�]H4bލ� W�ٲ33�eyOK���VYN�#���縣3S��8�uv3����`}�bhE)��Z9�i�j�SK�f����V7n�vgo,�d}"�W��7 ���-�k�T�q.����w,�gk��0f���On/��\�bԧi�`kF�����s0���i�1Α�E��X�� ڨ�s^�+���ǝy@���W{m�{�x��,l�$�r��&�û*#�nr>�(���	�:�ǥ�d����c!ݤ�Ƕ���2�{���3�)ɽ�X�wi�H�v3BG#��J�CJ/���"�3V9�DY^����(:��@Р}�`�=��t�VS��������#�I���E��q⫴>��(��oUlt"��Z�{FՓy�C�y6⺰��g�[�!h�b<W(��]��T�����M��:�&.U��-)�1+���7;k�q��9	�w4q�){jAR7h��p�����GV��ټ\��|s��:���vE��U�/�z|V�ot�=��k�H�ky5u�亦C��;�-�-��j��5m�E`�����mJA�n�r)���*k�.
sDΪ����)dxY*v�3��c��>q����@��pt��`5��TZ�Qg7��
�"��wu�E�S���gC9R��pS��EX����X�4����t�!��¨�ʵG G�kX�2�TqR�KH��B��q��N� �DT!s�a�g=B����,�X�X�G�^b��I��(t�m�R�1�x�p]����f��4җnh.�Yl��|沄/ �f��Z<��V�4(�c�;�<mJ�݅F�έ܂����.ُx�[�юp�-����:�Hi&�R��$��,�9� JܗyKT��=�Oiz�7.u���b!���[�XU�B���x��å��q^���b&�B��{�m�4���D4��GC�%���2:�ӎ�x�j8Nu��u�	EsR�d��j�6�s$�=�m�kiUoWK}�f�!���g7Og��ɱ�P�M5]w*՝�`suj\X��z0���P���BR;q��f��{��ggp,G%Σ� �C�������w���u�����OjRHt��r�Њ�>wC����
HV=Ld�"8ҳV��>��=�ݺ�h*5e��Dc���z��+��윝틦��K�+3 ���o��{O ͙�a�͚op�F�3i�z����Z�}G-�q��En���Fnh�X������5G5F�d�Ær߫C+�m�9XJ� ��6謇5�5��	=d��ȘE[HQv�N��7�P��K���ѻ��	-{��yy��}-aZ�X�i�M��r�(�4�"���c7�ݮp-���oe��ú�� ���c2n�tG����!ס�k����������U���v���z��y,��D���u�E��I��KHEQ�w3czUak�У����7\���[+��$+:@�� ��gX�+��M�N9�`;@t�g�}���°���T��੐q�gA�Ȏ>Z��DQ���q�i����F��;�j�tڱ[�q(i�ښ텋�A��t�N\�s;w�9ڦؾ�%1&J��%9a-�6P4�K��=8@Z�����Z�td�@�5�wU�PdP�/���6�9�	)˹6�B$f$���H��Yyv� -�湙�'!�	�6gqR��ɛ��@q��k�1*ih����4Ӓ�wI�9��M��u�8d'�@�F"D��FmĔ��ˋ<�V�v��4T�5��EW$޾ZjO�	Vno���i5����ۣ�%�h�ɷBq�N�&"��Avn�[X��햶�_I�V��]u��2� ��p;�4�����坽s�ǡ:��:��1���i(�Ю�l�W��0QqE���q[������ ��j��l���K:4t2�{;>�sM���X��vp�4�S4�m���5�)xkN!{����{������)�n�IO���p\D���������6�ie�}�	]�m���*<W.V�;�0�ʁNj��K�r/���< �.�s\�X� ��5�,��V���3^Kil�M;����G]�#^��tv�%��OMǊu���%=�L�)s�v#:���Ү��� g,��,�S�CӃ�=�.�qpl�������{f����7v�$ӱrwDvgr���
Oy	N+�L��	�;^D`��{��j�A�Vh85g݅��٨�ސ,O�)M.$�>=�R��.���mc�Ɇ��ʽY4&x�'h㕎#t��<�{���UgaK	{�ڴ-�c�h�L����=�wf�A+f�!Ge��{z
Rb��]��o.��)5�_�V��;��LBn���>�q>&`�B�l9�i�(�O���R�W��g,`�7V�Cѣ����}��27\��=SH�q��d�a�ݑ��i"���Obsg;�d���8�5�j�7gmC/hC@s��8��X��r��Lt��)�˟@M���p��
���)������g*�,]x�Ԝ��)$�Y̰������0�;��6`�.ڥ���齷V�\����b+7p,k�U��]�� �p��I$�t�R��OSjjT�3*]d��5zp�i�e|�4Y��x�s��d����^
��<m�m�F�� �y��Į��;��3N�i:`�yW��6:JT�^P���%�);��'ǞzH�^v��E$q���<�T���^Y5߸�o����}�ߜ�c�[�)��*�W[�]�^��,钾���M{���.�>�OQm�1n)�8@�7�5e�А˽�,Kr-I���WM/�Ie4`WD�KąGa�Jj5�8�;j�4N=�c�[�H���s��6n^�S���r.m#؞*�=yR&��l�]��c�!���gJ�5:��)n���(Xo�ʲ5V�Y,b�6n
�wD�kUt!N��%r����,a�=l������ض]:�nՍ!'`�U5��	�����ҹ`�D�F%�K\��'a��o]��6Lht�e
`�5��l�Y�D�ѐʥ�%����lUIJ��QY׌j$�'gE�Y):��} P��1�K� )�&]vV�K��*�Өk"���8Y:̑���V��&�G`���Qe�fS��F�H�lN�&��[N�Nu��{��J�VܛwND��:/��6�r�mj]�{����B9�4W{�e�#'��>�/�n�!i��kJB�)�I��Ym\�P�]䮘�܂S�.כ����2]9ڰd�K��d2�-�?ir���<�D�]���;v�ȵF� �V��Й���i�R�P�˨sZ�g��d����JR�5���h�ZAAT�w�j�$0�����Ì4x3]�2������]##̀���$�������V�$0m�miE)��y7t��	K	P���Y��N*���������o\ܫtd�2L��r��Žҡ-�ܹk8;a:ɸ�,�6~��P`�F��� ����
;���9
]&�[��`eVѴ�[�y*U�L��J����N�/tr��l��'1%s^R7)nS�:|ʒ���5E�.�����)r�h`>}����_{�Ӌ�8bI[��
�	38����Tv����BH�1י{_T���y�on�	 ͧ�F�y"�79�n�Fv�ή�0�Yq�ln��g�3�8"���t��Épuk�l�T�I���Ѻ8�+rgw|��.��R���,��K9��p�\���c��ߞ�4Xd��JP�D�wP��C�LP+ǖ�x �i����J7'�ڷD��`�-�&4��g;�x|sk�۸d��]�U�=���	��z#s^�4<rV)ں�q���0�&v�J�Qm�ፊmc���c[��=y�-H�HroCF:VȢM/��n�{ 2V�5[����7���s�L2��f��9�1Ź���3�j�U�IM�3`����G5+ôʒ��Ua{����܏GeDaGF�7T�W������FA�ʈ��:�|C���["��V���O�4X;{
�1�pV-ʮ!����*�y@�mǂ$n��l��l%wi��z if�P��geS:nL��H*^�����cX�ܻ���ب5�7G�Z
f�SF�;�y+[&�7f�^h�S�A�,���[D�K�o";����u���50���8h��+!g1�j�$��֞�"�*��x�ӵdZ��c�7�����,�q��Qe��%�.3C��Lc�wp�Z �L2�rq}�3zcrKr��֌]����C$����˂�9�l�Yoh'9�,|�[Úx�Vy,�g^ˈ-g$�H-3m9Nt����wq�^�D�fZ���>RN�������&����,C���XP�i>
k�_&��0���gE�f���ë�%HƝ��c5�-=_�4c���-2N�+��KօzA�ٲ��>����
��jf˦J�*�R�/~��R7�����7��t8�)݊Ύ�yk��Sn<�d�p�	�aݖD��m.�,�4Ϡs�5�g�V�D���L��^MHp��XM��A�8��"~�=ږ��`�6���"��] Lh��u��N��R ���Z��=㹔\K�r�u��U[�M�:/�L2��Y%,��Yr��R!���5>��d���{�!�v��Cq�cB�5�pr�Մ	b�r�v`���B���e!˚1V�`<�i aY�_.��O���('u��Һ�C{6vD]]�o5�������>�
��β�q��[ڞ2��Ҭ��:�)�S����N��9:�ȵ�k�U� (�Y3(L|���w���������>D�|M��57I��e6��u��`�5r� [��9:A��@�\�e�H���+����]4��F��ʦ�i��T�*\�H������ܔ��*�V��2t��NNh����o��iI��e,CV������.v��ӑ���J�9,���n˔�8\5��4\�Z���������|7��{8�e��(�`V��":����seS@L
F��]&��go/k@�n%�j4�e�	8��Y�:ru3��Z�ǅ�)�D�7i<�&��~����R�{&X�r�)=�jR]n�OpQn �E�l��RN�����=��J!��\&Xlս���Ͽ�g�|I$X
,�H,�J�%a$R� Y E "�$"�BH�E��(+$���I!"��,$a@�� 	!$Y	%d ��$��)$�+$�+	!Y
`P�T�� � �P��%a	��(�$ ���� XH�P�� �$P�"�Y	,�d���Y$VI	Y!%I%a!�@�E�)��	���! ) � $��$  ��I�!�����d���! BE�B�+E	$+ *%d V@T�+
H,��$XB
I �I � �H,���+	*E�I?���BC��$ I?����2���6������n���v�v�i�Q�+�q`����`��K=�qPU�:a�*�n�:U����||�&�lW3\�<��]��;E[��$����g��;���w*�5_/R��b����n_(V�yX(��}�g�y�/�g��s�R�s�:�	��B��L���2T���ظYQ�\��BU�8�(�f�B�|ky.ߒɇP��K)ւ��vz�Vf�����J"9��,�:f�3R��3iJ^ش�L�Ӽw���z��]_i�lC%��[��}";r�G��D(4���Lb��NQ�#�g�����P\�����%�~�و��w�n�I��>����Al��|y�>�Ȝ�ӈ�{�g������-��3�Γ����v1�\(�z�J�DJd�܃��Z*�4���H�k/>g�Mn�4Q�,�0N>��St���^��a81d��χ�|r��K:W�
뒇ϡ�Z[{�,�+�9�v]��:r-��緻��L���q�5r�XwM�i�50���  ��sJ�⻓�T�oL��i��|�֐>9gM.���fr�F�K��5�׽�d5��>Y���E��t\� #�D��Ǚ���ޞ�n��d(��s���w�|�����|�L�;A\�%|�E��xh܆������"Cm\M�>��ҳ��y={n�r�<az1LV�l�F����s�KJ�Z�hտ.��չw������a2ɚ�wi�{#o4�_?�6��]��z�ɬ^���.�ӱ�T�I�qI`���Kʗ"�׺�F-d�Z�3��W�����!K��=-g_m5�ɠO]��<D,�V�R�jyY�I��5p\f�6t%m�W�ٛ���s�́�<����<��,�Smw�]��j��Θnx۱F�8�Y����K9u��O����+�8\�U��B��$�oy�zS�;�޷�M�a^q�V�6�L�sR�n��"�N���f�;���O��Ž�fn�ѡ,UJ�Gu�p���#��CT��s\]0}�yx� ��}}��������[�)��V��i<Rѹ1�4�*���&G�ڒ�n8m�������]�up�U��t��t�e�\�� �,�(M�+�c=��}��%�!6�R�,̇0TUufQ�o*��!ZkC3-dа6S�yh�j��1��=���X7����jVFֈ32I�5����In����yX�=��W��]K�+j
�e�R.[���>W��Z��M�xٳ�e�%K|�/)W�C�E�M9��!Q��h�[���U�.��z��zFp%. ��:�g5�i	^��kͽ����+}1�}g�=��}�9�c��E�2��P�þ��]`"$p��b���;��Kʮo'�[{G�Uڍp:��::��r�z��J�4���Q�a��X��R�>x�ⲢЪ3:�>��l]֐+�f�={��h���#��5��c6<�G�LG�w=��]R�N䂝��Q�w��AFW�kv��މ�+뵎]}:�{Ͻ��"K���#;�|�a�C�.(���dƗ.���e,�ې��[F��g�l�H�F;׶
��h
�G��,���JRo|�-x��G�������{V�.��&l6�b�a��� f�����7�N�E��Gvjg�̐��K����U� *{�OQ���@�,ż4��^�3�ǳlO(:|H̬�7��{��3�98i��ܬ`�omԗ����龬�|�.�{�,J�˹Bz�Z�Y��Ut#��`x��'fj!�-4Vp[�����۞�|���$�k����˶;3�L��gm�e��T��Pw�4E�4�b�o�:53l���3_�uQ&?<:���؉l�p�w���G�.l9���L:��g;�W�d�,8�Z�s�e�`�1q(�1p*��kw1�`$tH�)��Z{~ї������yco�M�S]ܯtfn6�����j����=�M?9N���u2P��߈n�x��lh�3���`�5E�;�������77uf� �VƲ,�0�\}�E���OOa�.p*y_|q!�I���,�/E=]������[��~�]�i�\����A�H����vL*p��0��i�l�P��#�|A�)CE(V�K	��oM�nuN�3��f
��N\���C`��(����m���is#���Q�.�CaJ��s�"7
�>��`=���3����[�{��:U��yMz�� fRT(�;v0(gg��ݖC��3ׯ�鐸7�т@�;Vr�/�������ϲ:�p27;V%*��Vq�X��)���A�5�x-��r|&>�c���+E�j{��@`��Dޮ���vs3���;N)'U��N�s#�6���l��{z�6�nr���5}��eFO@�\^K�\"[H�<�6�w��o�@+i���$��M������	��W[������aY��/��^W��b�,��g����[�iY��M���Np��r��7q��o�CpѲ�ASe<إ�a�ީyrV�w�9v ��\���=�{stX{%��"	�g�E���aqw��Ѹ��~4�@{'�������Od�<��"�����A�}�@ʧ��:8��N�Fm�;[l��O�3��h4`e��f�|�\�f,c�?�΄�{~�rЗ��Ob�	��j��%�=�.��C,�Q����#l�*�dR�Y��K�ɾ��2p6^�u7�vɊʕX�6iy�8<|�͡hgdͥe��*��R�D�&��8߉�_ߟ��Ǜx0T�/��f&�˒O]W�<���͘�-�!NӇ��i�#R�����'	�5��:���UC�n��8jU�9n�
�>�۳���D�K�«��&.uۚ&M�y����F�
�;��O=�7
��Ҿ�u9���\7�M�bwλq��We�� �c|/�К�`��Y��7m[�ײ��X��c,]�Uկ��o���3:q+��qu'\!��v$����y�j3�*�4�w9t0$��$ǝ����8c�1��=��i������;�*yP��z���_E}���*�۷�fl��^�0�Yã]��W���#&��x�$�gq��c�e�3&�ʦ�_]�0\üH}������o{��5f�#��x5U��T���C�W;�O��J��WA�6��6�v�@n�J��Ge�����:��8�N��J��$*��}�ן*�x���=KM_^@�f��.�6�����B�\tf�r,��?sܑRDO�(Cz9��UA�%V��ȟ=���K�AQc���IL�+�a��)��=n��x�\q��7ܵW>ű���J�tA�^�q�bm�����iMz*�9��"�DŢ�6��R��)��X��X�op�+G8����)���>#!�+�:���{�d�;�����{J�au�j빥�o@�^��<��s�`K�/�b���]�a�IP�N�Zj3�v�yHN�φฤ&�{��O��w�Wâ.2�v.�-ڀ�;́൉ܽ�;��sv�s�R`.�W��d��]�JЪ+۽�T��}�EE7��c�;|�Ƥ�eh���]N�!W]�6kӧ0r	pp�W��2��."v�����9��ý�{���6L'Nm��<<���F��B�>^���"lv�_lr���R]#��[�
�$���sv�(L:V��/D���(�tt�77c+C�4���]��ٕ/�g�i�[`�I�S�pF�x\�݌��F��&�<�v�N�,-�3uI;����X�c�{�K]�Ƅrl��5�,������hr�=�gd�ۮL�ۣ��YqP7w�(J�[��2�������oEk��^#����2��㈄�@��tu6Ȅ�.B7cͲ��wg�k9Q$�9J����|;,K�B+���:ټ�Ȇ�K����s��eu�-X=[5�;���OR]�
��}���dsV}����=����_.�Pe#:]��N��b���>ү,� ��~�< Q���\�l�u�<��}E))�Pr B�h�{r�\�Wi�f��6���G�r��t�J����R�\�X�=�\�Q���S��uE�Z+�r��6V}��&#ox�
��d��ע���u	�ğo1iq�qS�5Ou�� �xD}�k�N/��\0�5wԴ�+�K���mU�0���en.�����BvJ��J�u�&Q���
�8N�Ծ��O�x��/�*9j��,�/4⨭�~y�(:�ei���uN���ݛ�اMK��ft�����;�F�y{���{t��t�� ��h�3t��͈ya���6���-y80}}��N���V[���Ҏ㧕X�L��%t�h�X����@�S��%|;�X{KxtX��/�P�ʕ���3�� ��Mn��3�v1�4��������.w[z�`܏��ni�"3�&���ukV���w�	�%1��I�7��=���2R��s�J4d�/w)�d�������t�c�ٞ��ĉ�r��ў�3�z�2���>8�wL�#.�j��o��W���s�hȝ$�1�ͳ�xx�[����Ldmi�˒�T�3�+��7f���܅����H��h�v_ �M��;y�+���t{��d�e��^�������Sz�ɣB�i�Ho 4[D�[sP�� ���E[������ļ�n�r�{#7�E��6�ۗ��R���t�}�OF�x�o���@%�x~ CASKu�Z�1����ș�f��S���@PA�S��Oj�NK�Xp�v���,��Z��/�k��9-7��>��[f���T�3�4)��u;��Kh�{\+d޽U���[��T0S��?1F�o�'�f��>��v��u[����䠌q�֋zc�5
���GqD���� wƮ�	�-�S<{P���>��<Xyt���O  b���:����TH9{��i�Ld����ڛ��﵈;:"�6��tz����1Y�ڒ����nf���t�q����m}�'ig�|�ɫf�G��Irg��Zc<�{(��U3�wT�[�V���t! �$'����_bs7�5�r���e8��;���^\�Y��gI{���զgu�&Z���zAN��[z"���\��>�����r���Vk�`�T���ɐ�v�=>x����/b�u7t�>p�����Ry���	Ѱ>�Y"��/!rv:]��f�S�5��Y�3o�n�X�v��&�+���xc���0&��.���=؏��x�px����r�w:0����fcUDm,ۑ��0� ca���Ƈ��.m�l'�P����G��y�#p�^��#���a<S�s$:1�/csqn�с���q��Ê�W�:�����t��	*���g��7ʱ�4I��s��H
�S��]h�Zǝ)Q�}�<�l7P~�Zq���㉖���l��Ρ�[�0c��to#��U���o�y�|���rX����t�̂��N�ó�� �8BiڙV7�k{���#�.C����xn
��#X�wn(:���dm���g�8����;���E���`�1�߮	蔾�U^x�u�i���"A�{�����-��p�}gEG��"b�Q����uKˍYY.������Yj�uu�|89y���檹�=*Z�^nռ��p�����Ĕ�尛�5�5Ŧ+5���k����瓎�3���N�Vv���k�/�mԲ�3�3�n�'	A�A�@ �{�YQ���yf3e=��x5����׵�ȗk\n���d�n�α�-^՚}��2rDɻx"+M��n_[Ӵ܈��$x�Ń�w���tjg����͙�9��-MW���*��͑��H*�T�mݜ[����.����o#4�����i��ݞ�|���Q�����[����=��Y�aw����G�m��L`VJ:,��u�����sq���ѿ2C
����s��k$����.v�|6�fP�Ɩ��EZ�}!�u��1n^���ި�+�֯��Q�#�Ggs�T{�p�64�2I�aqn�Fc1��h�V&X�H����N���vn��.s�}��OU�,g�3�y�婢��E���+`Y�,���6fzB���[c�7�8��ˢ�>�5�=��lDg]y����B8I:��f�*�b��tt���)��=�t��j�/�͂���8��Y�Iy���-Ga����P�]�.�]�;�w�
N%�k�������;|M�v\K\��C�q�5�j�t.)��t�oc�@�V�p,�'X�;�3#k�w#����6x���e���N�j3��Ld;�p+2�~[�F�f@Z��&���0�їKW��Ѓ�{Jtq�`�WG�����*�)�^Y9vw��9u����O��Y�Yy��N�{�W:�3�#�gD�N�fjzl�w����Q{���E������gD�`�{�N�M�,+ݜ����[w�x�BnV��+��"m��.�zd
�jX�����<���GM�*i�8���5mmt��]J<�SB�O����Ƀ�8>�1:�q�O���Ł��↽�r�%o6�����bmTa>���u�
�����+��ʦC����s�����H���wGIQ�/].�$�����kz�tK�6�T�-�lμ����]s����p.�YSa8��n���E�{��1%m�e��b5�F�=�6n��_n���զ�k��V╋��NޭL�0,�m톣\0�>��wTW�y<q+��ȸ�/�@���ldx�%�%n�H�/0:���Y�Ld��0I�Y18�jq��̦Xql���}2l�+�f9�_l�u�\���a�B���e�ǟπ��<���{������n,�����m4z;n��V���G�Zs�:̇-��k�M��۴��I.7"�S����=F{m�R��ɪһ��x�w�����>����.(Vw=�w�s��.�v'���.���ۧ�ym�#�9ȔݻCǉ��]��b����tXV�tk��FȀ�7F����<n�v8��,��Q�;�۩G��:����5�ug�P�]e�̓rdJ��R��M����X�+8rT�\�y�1���kl�v�d�6�l�0a̬��r�l���m�=�wA�	����0�㳲�ζ�W;V���QݻO=n�l�e$X�X�6o8��t;��=j�b�}N�i��ڙ���l��woS��Hwh{& �Tه!3�s���[r������.ڟ����p��U�S]Z�t���h�[�Wc�i�`<�l�A�����;���|^sѬ�vq�ۡ,NVӹ��|�;���{l�n��{m�tR]���<��Y�[lu�kc��6�t���:����ݫ�Ƹz�Y�:�^�w;��f�g�F,�خ�5ۃ\r��<sl����{H`2Q�l6ml[.�mG��Z޸56ۯ)s#]i��:�x���ɮ��6���3��8�8�;e�peֱ։����,�K�tX9�^��-ꞧ[L���k�����s�q�&8�6�͋V���w\�����AH��&f�����Uѣ������P��m��Z�gGiNn݋2�]uѵ��h�ݶ���3�s�5����۱�7n��0u\;��e�^^�c;���#Ч��jy�;m8td�tm�!۰�9�t�0��ix�!1�n;ڰW<���؝�-�Xy�7lty��7Y��z��IE������֎��I���w5������g:ͨ<�O�r���mpg��D�s�����S
m�6�osۡ SumWX�l�viv��-� �aսy�x�
l�\��Ƹ�ƹ�lgf7lc)q��ptZ���^^`��]��l���N�����ss�Z�l����<\n�3��6�;r��pTey�G�[��9�@��=1�>Ʒ1\��h{-�݇�T��8 Pɀu�j[�S�nD8�sJ�xw(v8�T��N�ۘn�ӳc���x�چݶ��׸ݬ�ٹ6|�F��{4oR�k�;V��<�5�9�
��Vq��[�9�����=F����v�ý\n+�/�Z�ƭe]mc��pdy��-�Y��	�˞�Nwb��	$z���xzq�����Y.v\p�<�l�k�����6a]Ԇ�ڱ��^�e���fw[��3Q�j��D���6�+�p���ݽ]]�;���sn5���#�����}��qv�'��vy�x�Um�����Ðp�[s���f�&����z�	=F{Y�p�]n��������b�n��s�v��q��<���)��s�.N��vl!��õ����s�i}�ك��e��m�d��-��<�vJ�pu6��hO#�r��k��wa�;W�v�vط<m��q�r��xa�6��g�n�m�dÓ��u)�����Fݺsشm�Htp��vmGj�u����FQzW7i0 u��+֒ӻ�Ɠ/8lq��k��V#�k�r�'n^x�dܦ���Vxw�y�ş]�y<���ճ:��=��9��i�v�3���/��/��7�]!8ǰv-��x�O7=���6��kۦ9���9؞��v�79�p�ؽ�&`y��d�ݻ='"m����u��d�����8�yßm6������v��;Ӱ�m7X�4u7[�7Y�V��K׭��۸�dP���+��dޮ��lS���M�z����秞C��k��c��Үݴprv��3&����ӹ4�hy��]��\mĚGG�6{��Ѕ78ᖊ4��Mu����5��g�ݛ> .��La]�8�w7c��c�uvq����ݝ&�#W=��tȓ��gu�{sĻ�⓺�܇��-��#m����t�]e�wN�[u��Lz���z��@��L�x�m&��v�d��ٛv�N�j�<�y�V��n:n��+�kp��w5��۩7�=]�u�7��=��$��r�[0[��"���R,��n9��ҥ[�)��m���rk�I:��^q�,���xv�t�Ϟ�	�krF�����[���F��+;��˚6�{�+�w@��W�C�vs��;`ݮ���{P�<��ʗ�ܨt������ݰ�6nn���m�[v'�������󙫯n�pK%.��m����]Ak�'�칞Kv�n�Þ̓[�6{S�B��vt�`y�F��ٴ[\���,{Yx��s�ŧg�G^�xC]j� e8�'n�b��k�Ÿ������F^f퉤��,��`C1ێ]�wqP��z1WGl:��r������"��)-�Ƕ냏nx�ȝ��������wQ�7�y�˺��.Y��`�6��e'g5��y�Q0�\n��y�M�fݵq���{%S��㨢�v�A��v��v�z�`�Wn(Gfr��E����7G��ϸX|u�l%�5�",���mѪ��2G
��Iڞ]`��򋺞|Ѹn���p���v1�:���Kֻ�.��ny�:C�z��.ՠs;����&:nc��gc"�N�q�vkuv�8���:ȕq��_7oad��c���k��)��h��i���,I���K&�]�n����ʛ�r���X����.{vE�Jn7�xc /;vy�Y���5r�㣶��6c��ѯi�	a
�n�[tպ�m\�c�����Ǳ�lsv$����#��8u̦G2��kl�.B�'V����^w����&�Z��{.��0>n�=�썤L/3�c/XZզu*v�5͸cv"x�B᷈�[XN���{;Ia�J7-L�<S�ٻbp�N�v����萳���Oh����S�d�<���N1vm�.;\q�=��60�y�[�c���o�s���v�;BE�o��Q�<]+�6��^��ͫ�z�2㮺��m����h)mp`n�2����쩱��y������מ����wm�P����m)�����q�7ot/�����]�G[k�vǅ5��D�����m���m�r����s����o;Y�g[��бӎ��f�>}�K�X�,��v'wnp{8�#`献��rn�q�X���X�4]F��FҀ\j4wX�n|�0zcv��:��ͬ���X�Si6:�'�����n�zr{�Le��D��n�tv.�s��sl����n��h[�\���v�N�Wu9�^=�ö�3����2�c��J����9�aL��>yץ,q���PmW�����L���Í�
�u@z9�����ͱ�����5��B�)D���%�����"�g!��
��N�;�f�!(=��x��7$=�L
��%����a�v�=�˶|O.��X���t�������hv�������/Zͷ>K��)!ri�c��b"4�+u���z7<z۝78x{�'�����7g�	�0p
�c�{�V�����nz�;iU�{����>�o',p�[q������<� {��q�+�{g����&����F�ϺZ�{:�G6����9��\���0O<s�ڻf-��'gۜ���qю�{K����_e�Ʈpj���n��P��w�s�s9�X���K������H���˰<tvl�u���玞��
k���]��썹yĕ�:���Xض�������%�q�Nz����{@���`yϲ�;�V�F���M��]�,#mҙ��7on���֢�+m��kP�"��À�j�v:{KJ�����N7i6G���A}�8�cv�Du��x�ݭ�x9��[���ˣ�L=���G��x��V�w[�3�LcAh�!�\v6�t�9����u�t����\��ڭv��n<�K�Ak�݀痥��D�ƹ��o%�w�������N��lloU��K���T���
f��� ��Y�݋1���;e��[��f�n�(�n����ˁv���DRc��u��-���Մ�g33ۯ\IŮ]��ˮ N�-����b�����#;u���og]����y�rn�Y۳)�g����CC�M���ue��S>�NSK��8}ŷs�1�ر���vݮNP���s��<ob�O7dǓ�#�\�p��fN^���]�uWg��/a�u��9��ۥ<Y�3����{�.�ܾy��Z�N;��y9�!��b��;�^y�j�I0l�84=q�X�=\���mn���e�m/rO=v�`q˜�	c��㋷]Գ�����x%z��}d�v�{[s���[���֧.}��8�]g9�W��P:��[Sö�q�5(�+��n������"U��^�yd&]O9�sۧk����k'��v��`q�۳\m:3��rTK��[5�T�-�zVza`�<���&�ћ���ݺ�c��z��j71��N.��^ڹB:��knګ�]ȼpr��n��Y�b���盩=@�B����\�x�6���p��Vd�<k�:�u�/kfR8��o7#<�v�7r����X3u��^㠮z�=��;������n�6vw2+�'Y��cY34;vA�]�M���9Ր]��;]4/��8+<�z�؜%պHٮ�6Zqn�d�����{s����ܱ�w\;M�\hF�y���v�3�y]�[�v�gcg������s�갗��9����u�zy;'h:{W<�l�s��:��^D�q��rC�ƫW89�ׯ"�ٌ�p�je��n�	�C�`���T/ήWCƹ��hv���Juթ��՚+4�w]kM����6����7Qv�ѹ��s��zR₷f��#��B��[��u�]�*�u�T�מ�4�L�H])���mV}�\7j'cVܗ5��k����OvIlV&��g<{�p���G^=��� ��b�b�l�F+F�Uf-0�mJ1�Q(�R�)L��1��5E�D�4+�[b�V�b���"%m�l�8�0Z*�G\Q��m
�Q������(T*V
���ԥR��J��T�XTZ�[nS	iQũl���")*V�F�ۛqh*ڶL8V��h�����Z+--p�ZԴlPQ�[JL�U�*
mAl��1�ڠ�j-�[b-*ъ�!YaF�)q����j��ʍ��V�KD���YR���X�-��(8h�\bTh�[U���,C�#�R�8�6�U+EU[�2�
��ĵ(�jR�����8�vݷq��xw9OK�D�֣F�ZZ1���S����$p{n�;�sm�ڪR��[h��YR�iK?=�{��w󚇍69�m��|�ٹ�cuu��w� ��n��.�4r ��=�s\㝒���ڸ��o�Ogn�l��Q�E�r�nd-����F�Ci��LsZ�s���v8tq��4nND.��ܻV.�6t�n3����e|��!=\B���ՌA\]�{:	�l�ۮ��M���Ua�����!��l��t�28On�N����g�N�U�Z�Ak���nuۦ�xLT�s�\n��NBSY�ا�G$����8��d�1��l]WUyv8�r�t�C���xom�/9��Ͼ\�|7�o���+N�ɵ���w]��v���v�3{8�ެ�]�����X�ua瓎]�v�ϖ���͕��y3&��m�nN��#��]�\�s�	Zu�V��y��
j�(l3�vnݭ�F{q�t��rr\�ln�k��
R^��������.�/���W�#I����m��Y5iУ�v���/6����ݎ'�a�r.M�ܞ���`Mv���qb.�����G\��Jљ�.��*��Ž�ƺ���t!�ܻt\�v��N&dg{n<h��c������M2G�=<b�n*�����Ӏl�u��T��c�
�
Yeƻ�,a�%��x^�d�:׬ /s٩R�y�*�;�U���lJ�Bu=Rc��W��|'l[�rb��ҮM��0smü�"�!{p�����^��o�2u�Rl-<5�7)�/'X.�V��n@�;e����V�6�7g��˲zB�^y�v���ۚm�<���:�f-��a�7 �>r7B�v1����n���w��ʿ4�\;Ŗ�pq;vxq�7��hn#/.�.w�[��F�yPʄ���s�sRq�m�����y�	�D�aC��t��XΒ��3�y>=�_k�}��f��5�ܗt�{����.�z:�um˸��۬(s�r�Uڍtr^����gl�V�+���l�U�-�(Wg*�7Ub&�uS����|k�=�y��KA.�R�Z3�LQ�Ҭ�m��ݗ��om�{9�w�T�y8�����;&ݗ*�l��n�eC�U7m�a1�����'��aW�@xN6v{gp��L�y8ݹ�p��^˸1��q�;g�;v�x6p`y�ۃ>�y��c�����=��l�q��+�O;.ɹ3�r��<=�7�v�ϓr���ax9v��?�����f	z���q��	v�C���w�I�˫)�ܯ��{Ͳ	$����?�׶a
h*&h��F�;�i�&t*��<���O^K`|�������n��{w'�u���9����TD����=t���̯4 3���_]Z��� ��"MzI�*$��E�P��(�f�/{/f�a]l� x�n�@]��p�@#�{n&:vWz�i�����FǓڙ���MP9en�6 �ݮҳ����%f0���h��� f���f,�cEK���?  i�� ��8K/oV�z���ή�v��<ny���ˢ0=�|������1	�K	;q�> 7s+� nokve��}8v����]���DO����M�Ϊ��� �f�h���ݑ�gM=�����`��܆� 8���i<�Y���l��>يh|=7�����x�N�\���k����[�{WC���z�h�]��䩈��2�@vomݐ�Ϊ�gΎ{>�:�P*��&���=�y�6� /7��V j��1Ok2s]ϵ ���3�DF���VW&jTL|U*"J�)���;�`De�טD���v��3$axF��{�������j!P�+z�X$A��y����W�3��d��4�I.��&�D�޺���C�p#3{WA㞉j�	. u�9�R����9.��ў�q����.�n"���~��8��`���[��1��'{�jť�@?�؀ѻ�E��0EMl�I'�{n�>�����D�W�cA���X]���#_��̯p���ۻ����}�>[Z�ةWf���t�Ω�����k�6��_]�" ��ښ^I%;�)X�1�:���[gF����������؎rɹv9�Kn%��kNWϬ��s!�s�Վ`;r[�1'��"�g[c�I��d�m���ݽ��%s~�P*�TMD�8��׮���L��z�p` e7�ŀ��޽rI4;3&��6���7�D���_��v�jg(AJ����|�� ���A�]�"ȁ���M�]��@m�6@fg�5�z�Z^Q���Æ��4�`$D��̺'��qۗ[��Xᒖ�Í'�qֺ9�Z�?w�~�;p�ۦ"j<r'ݹw`� #6������?�x�A���y��4I�g>�_"DO�f
��EMH9���7|�эPRv���\��@Os�K�O��I�k� �O^�`ӷVZ�w]]Gc�`��L�4�Ȉ;^y�G^�y� vT��x���r������>�� �O�����Y�5D� B����7�{x�y>#���$95Z� �7&��$�w����4M�j��W'�%B��gC�$w��uz��\���l/�W>J��e�<�[�4���"	fj��R}3M���%��p'ٔ�`�oܪT
*j�Fѭ�6� A����e[���._�岉��Uh���P`^�c�c]F���t��[q�uS5�0n�f����2S����]�9���܈]Mգ�ݹ��SQV���>*�%ou>~qķ�5Q&� �w�n�[����M��u�L���y�p��D��B&_I0�*
'{.�<Ka>�кQS}SI rj "C�z'L��{Y�^�cw4�a� [`ai�uo�����~�{��`	��}Q��{ӕ����� /w���JqdR�jBT�e
D��W�D؜�sSnR@%��漀 3;���  ݽ�{�!{"qnF��?8.��j�� !L��q�O^�D��	�y9�¥�k���i ���`|��ٖ毅ދ�#Ý�M�܌�,�yI�"��ӗ��O)�{
+��nGFp����u��w�n+�b��|̻T�,#Y�.�XG����N9x�x�	@��ja�:������o1۷d��G�/c�ӷ9�Y�u'n}��m�ĕ��r���Ӡ�[�\h��o.�0p�i�cn�+y�ͯv�2�@�9j��f<V�B��=��4���+��!��U���Zvv�^C��^�u��NûX������|���%�ׄZ���my�-p:86e����f�����;Q�ܝoU�<��WX5�T9'��6�%q{���@�e�aٜs�	$�2y�  �L�s��tVȳ+�-A  H�����5C�">*�%8��裂 Ù�q�&���I$����$��=ϳ@D� {�q��a�F�/c	%�;�B���ҥ��F�I�֗��i2��_w{68�n���" ݽ����T�U*��(�,����[ތ�{ �y݀ |n�ӈ`u���A��}��6ɬ% _s��cm��0P�I[��I%��\��k�1v��}w(6�m�@ �n޹$���$�Ψl��m�ZL �p��f�^xݼ�-��#2�W��+\�N�+�Rn8���owT�R�B����qh��j4I$���PTM[����^�]�wdD�{^�%ꨕT

��$���_ ^��yj�1>̥�c�k*Vd����1�����Lb��0d���㏧��-���:/�ٞ��������� �n��`|w��` �T��tuj�
1޸���Pꈏ��DIM�u>k���y� �W�;n{d$����'Ϧ����Y!AA�	�eR����mx���Ð� ���P�O�~����D������ҷc�F;�@��84XA�PE��)9���� >�n<�SW��֥������^���}wd���?��%Ǥ��
i��l��!�Ny0���8y�{v��V�;jn�ӳ$��}��}�*���7����@^�y��ݾ��~Q��G���3:�d��8.��j��
j�	��ۗjȊ�Ԓ�Q$�y�j
� ������5�u���Uz���U$U�0�2�G�v%�  �?'L�d��Sވ]G���m�ʺW7�k���=�韩~[OM�6�É7�^�}�%,�U����K��Ϭ�s	��}���g�4 ��]�d�f��P��h���;�'��V�{�$��c� ݝ}wa�yY�fu�.iui���ښ4^���$((?A0�*^���V �x����:��������E[�T�)om��7�[��N�2y�;p��)�nٳ��(�:�[�%�$ռ[��k���i"PCw���$�x�(,y�.��!�7��݂�ݼ��ͬ�Ww]������ ��waJ�
ZM!wXE�H�E�5Z�=�-�rN�R��t�;z�� �����٠��.�πR�r��*�"&��;��v�";��@�[���O:�~ ����A�yM0ɭȩ"�AS���}����L~}FP���z��$ ���Dv����ۨ7ؽ�}'7\е��ğ�]��)D�xee���.��;�7YHLW�(i�B�:p��j*��!�x"&��S�!�h͞�3}C�;�h2�Ey����y�{��jJ�^��op{�I� }�3@_�4�����֍o��q�da�"�ŏ	�7���1����A��8,u�<۶9� ����?�~�������շ�X Fu�� @v�y�E)�����N��<�m����3B	���O�ĪNY[�M�>
��&���
�W�U��e�V �yN!������."򼺰�vo%d��fHɥ�"`^��~`ney�A�C/vrj��� :� �3�)u�P�8a��6BAwM�ͪ�׻���> #}��π@v�y�C@��c���\K�t�@�u�y5�'&jAATs�q$^J�{jŭ:��^�\��� G��� ��8` ���w�����aC�����V�'��uc�p7���O]�y�ݰ��*��pۭX���N'�UV�]T�َ�"Fq�A�ӄ�L^�`�������."���;��Q����i�t��J&6պpgt'Jv�I��m�n\��QX���,���4�HZ�n�N���Է)�՘�r�s��v�A�1������kK\<t��%,X0���� ]���r��;�"�|W��۱н{9�Y7�6����=����p�
��j�/n�˗��]q��p�r�Gh+8�u�\���W�뵺��X��Rv�n4Z�D�[\t	u���v�T��ٗ�������]qk����Z� >�5I ק{���}Q���	�8v޹'����j��� �p|a��f7�@!8ݞ��&���yw�^ ����P�۽�q�u� ~��W����Q�
cr��Gwv�z⺥�[]f;]x�j��h�	�{j�@�P��0T�*�[��+&m��� ���I#s{j��ոcu&3�'hlvn�DT\l0�0�F!	y�H�;j�f�gn*Ez{/�Ex��ݵ@��V���]��ؠV̼����2�Ba��=��]�u۷c�x�zR�S��/7����������v&�./�kn������N�[
x�T���bF(���	#3�+£��* �3+(�ϼr=�Y}���zUӏ�N��ٝ�KU`�xrA�]�7'�}��w��ء��A�-�`��V��C��t�{F���.oz��I���^����zW�y[��U )�zj>��� �|u6rD,�꛾�O���lD ��cފ������
��y�I��@�s���ڶ$�7ƚI�Pa��//��ؖ�^����D� �<� &��f��+�LvfW�����A�`�!ùM <��_>
簜O�-�y/��#y��ro�|=�	za��5:�����I��y5ų��+��c۠9�\=,[a�Q���y�=4��UH���:m�p���w"H �]�P9P��q5�Ա��;B�#2��5�I�P� �8$����k����/n�] Bsy�U&�4'9�����΃�������*d�&\�:'&H��e�"���$���F����>�^���.�J��Rձ���q�eܦ�:�sf�A�F,r1�v��UgP�]��ˑ�t�7;ZJ\r�6E�Vf���G��>��G���i��8ߓ��p��$����7�
��51v�3a���[��pQ9}ǌ[4ïfAj�v��=�����_n8w��Ȉ
E��p}ܸ�R�!�.�������D� %�g"V�i�<f�H`3zxg:�"�3����~J*>���r�Ʒ}y��/n�Yw>�hz{"xb�(�!���h��s�~�CۊNZ�^F�>��7ü�FV0ᭋ:&��X�#��j�kmp�f���]�	�����;�Εݛ������s+7*L�����4洫����ώ$r���^��|�Y�Wn�'�xm���-��Q��t��Wӱ�<�����bz����i��]����������)�8L&5:��{I�łj`zOi��Za���A{i�^�3q��z���'���X������i�'�ON�|�%��RY)q_a�9 K˶Q��|�ry/ӷP撦_�d8���a�����Yf=R�0^���bD�z��Ē٩�sUGr���[u����Υ����<�ZvC�\�1�P�p��#]�ٛp�9)I$E���NB7x������<�Ѿ適[�[N%�E�9\���l���)F- ���͓�M!�|�-b��G�r�f��&���Q;W�v��;ޛ*wG�??��K{�t}gϱŭ�'��u��n�K#�����%��J\��S<h�k��w��\s��@��A Q&��U�m��(ť���m�V�6���%�LJ5�JPiJ5��R�F�K[��*�R�EJі؉hX��СX6��ZU�-���J�)mJ�ŭ*Ѭ0�LZ(���H��QTJ���
�Z��+
P���K
�%bȴŦiaKA�Fڪ-j�T�UKE������B�2���-е��D�ؘ�f�͖1�TU+�pԊ�D�E��4�	�XR�l�+�QAjUX�V�Ÿ�
�B�(����B��1J*��������mX��0�TJ�jU�����G6��U�T��ƍ��+��Q�s�Q�Z�V��QeR��ks�8�7)�2��DH�8��sj��#VQ�Ԣ*�*�Q+DX��XUG)\�	�1T�TkX%��(���k�R�Jj��˅I���Z�X���kE�U�R� Ԣ�m!�(�+R�J֍sB�F5��-kh�ĥ���	Z����Z�e*V[b
1���eqVPf��*#00�bTZ�Z��J���e���Ķ�D���`qJԪa�b*��e��kEm�0���Q�EAXԦ����W�s��A��09db!"�Ṗ�����6��*���|�6dH���	��̅��W3T�������bL�I����ؼ ��� �^�z*�s�z��Tq��ӐH�����@;��U����"�����m3��o=��!ݘ�����.v����^w[:��H"� ��[�8r~OE�@��N��6��h;��Tj`e������7j��Ezdsa8a��m$�ul�Ֆ7np���@$��۽�(B%���{*�q�$Ǆ�"�!(pH�]�������H �KRS��I���&�7*�$�۽�^�,�d0�l0�s�:'+�xum���Y5[b�c��W����� w.����]B���@Mݞ�˚�9��®�w�#r��#�ք T\���s]X�ׁk�x?.�����oI�f�s�O���;�rx[記�s`�
���TI#6�@����RT h�^'/�d	�w+�$�]�0+7�:�6�b"<{с��Wn�s�J�]1�c�e�p<����Ǯyx�bx�帋����)s1��+�VvUx���&��.܌��߫jw�{�$
�j>�T�t��ED*���"L�!nԉ>-Uʶ���=�Q�Nd�$�n�Ux�Hr��>4\���������k�[	��[h/r����۹�H/SDD�H��WG-���n�P	�nI��"�!(L�fvfC��2⅑�l��Iq���+��G$�<Z�{EH_Q�*Y$!�.A�� �U��F9��/V����{�\׉�>6��$����v��Um�Yv7�wg���a�9�^���k��z��5*�T]����)�l��"�RyY��Daf�X�go
�R'n���6��y����&�C $1��>x����X�Y_=X%3�\�Ru��c#giQ���nxyk�q�D�1ۍ����wυ�8�u�'#9ݴӧ1=�[���룣[�q�gWn[EÂ��f<)�/[K��t���ya�s����&G{v�"�� =�$����؍���U����O:�a'�c���&n]m�m����k���
��j�Et�����nY.õ\�hݫ�9�.�X��1�,�&��_�Z��j�w�~~��!C3�{�D�3n�I �����_y��F��_#y���l���H�	����5㉣y��wA��xQ�N�ېH'j�*�'j' �DHnv�:���Ш0rQ�D���jF���I�}�+y<8N�"��H�8��ɢZ�6�a�I��ܛ���K3�A�S$�z�2�ĂN��
y��h�#��$T_#`���K���%@W���j}9�� zg�:�r��A���𫱓�2s�9>���*��F�v�K���4$���b=��b4<r��7V��a�HC.�����XL�lN�$�gd�$�۽�@�T-�aq�;�EVvUGdE�A��Q�}�^���,v����3�^���uco�$(�C�,;;/z�*S�Ղ� d���:"�,�&�`e�:��n�
�轢jD)����wd��s{*����~3�TU�w%�DӁ����;��` |=�z$ �U�c������WG��W_UI=��^�V����B$�wh�4z��o��'n��Q?�މ| ��ڛVZ��e���@�\�(m6m����:ڣ�O��=]�6>[����$ 	;�U*�՘7���i�$�6[�
1#�,WJ���.< @�Y7:1������W�s/���~�y��M�K�ٜ��I �wd�$��j�W<<_wop�n��j��I��ʣN���JL&\�����wwM��_NT�ީu3�I"�*�'V�ē��v�t3Q[u��}θ�)'6�� ��f��we
>'���d����Ӽ��I͝��ȣ�kb�w�N���8l���]#�ޣ�j���_��*��ڂg,�!�{/ffB�ͩ���jȘi����'�7{(P �jڸ�	)��M��B����~f�zx��<D��У�|N-��� ������\WX�_<���qdZ�:���4	ݜ~��ɠoz���N�k3T$��쎭���]WI=M�*bا�&?<Z����b�ݺ����m�'Of.��R�9�����Μq�㋹������0�m8�[4Iӵr$�]�"��7�bs�ۛ���ڸ�Uj�a �4���uV�W� �����l��p� ��j�I'j嬨 ��v�ˬ��;���b��'EK,�&���+���(��� �˚{d�� �����w����K�7(zXd10"�_u��r#.�;��ʉ� M�P�r$ ��V�5�X���u49���AOM��ʇ�}Ws�^�M�KL�Y��X9����tC�l��%N�ֳ�H�S�*6V�<�dǖ�I�(C��ܪ�w���lFDWGI5;S�$W���ܪ�$���q`�'/ �D�"�2��Q����9[�C���6�p�n�5��{6�(??���*"i�Q���$��̚���HM��cg�^�W��*_CllB0چm�����ddz�V����ʭ� �GVfUI�z�P �Qv:&�b�nv#�x�1��*h"����[@
���R �'@>i;�����*$�}�uD@Ⴅ�`D@p�eϏ�ɭ��΄��$��4A��]P�EWKP��G��މ 7hN�`e^XD3TT�ez� �Ŧ�
p)�.+v�x�o���x�ȬR{ћ}D�����S�a;���u��{�Mv�pf>���4�A��]n4����M?R�EB��ǢH�L�r�y�V�K�s����돿^�����q�p���ɶ�勘���Z��;�p�ZmmЄ��=s�S*L�vn.x9y��2��rh�۞3���vV�K��3pc�b㣶�hwk�.n�÷9��lݰ��F�Sl�7���O�[u(�6��1�c�Kv*.��[�,���ϱ`�yZ����A��"�!���h���+�<�n]q���S(ٵn�4����+���4"-����n��n�[v�:�Zs�խ��4��Ps��߿~��+>����D�;���@��ȬR�i���Q�V�`��5���y��,�ر���� n��혆�����圿Gd�A&�z�'r+�6��ROO7]~8b�D#�bm$�TI ���|H �sᦊ���	� �ut�;��y�c&)@���o����<���zX�1�(O�y�U�y�I$mv�rޣ�Ԙ�	enP��,�"l���m��^�'���w�Y�j��Z�@��*e��\f��yg�F����^��K�mtQ�z�v������r�v��Èk4�ȱ@"!������	9�� /tHa{^��yA�F�
�:Z� ��Qh�M��F�E��Q �DW���^����l�Τ�J�v�vʥ�֫��|X�j'eұ;�r��+*���9j;�'5}��8ص�X#�Ӷ6��xw�S�$��+����Է�´Ko�Hrߝ�p���@H�j`�z�rh���t�{�劬�H̊��ۜ'Y؄a�Am�����Z�g��2Iv��A�����^M����ԻM_�SW�hSr���J!�\OK��$���3x{��np$]Eb�v�rh�A���5H(=�������K������Z��GP��v ����&:�z�nx�z.Gkml�������޴�<Wk1�;�A� �f��>$_muQ�DK�vj���O�]�T	����DC5@���9��b���ݦ�E;ҥЀI���P�/v��^Q:6�.�*j6��A���!�$a����ʠ>{�?��f�(����m�����T�9���
�Z]���w�y`�����4'���m�k�2���5F�E۝������`$.�u�/y�-�5�+b�j͟��yR���ܚ$���ʟ\:���p�&��hHH)=�	��ۚ�Nn���V"^D��흃��g'<	�����1��{�d���DXt�c""���@$Lu���]���j%����>[��eX�f�^��j���J��B�7����٢6紤k@`�s_���TC$@�i���$��sDn*ôG<"�k������k�==搫�T�I��(	�Yrz���X�W�;�.�7ּǾ��;�* t*�5�)xXY������fF-�j� ̂��(�j�� {�ͧ=G��%���I ��\�$nEbq�p�6�z�&ߺ/����.mJ��kT�P�^��^��ُ׽K�R�yQ!��π�f�5�r�s�5%(�%J�qJ��La.J��j�[�j��^���Wꈭ����;H����Ɲ���}��xy�&vkj����L�D8iTW-�?C�}6�*׎�n�ư=ԕP�X����̪9�iYSq�%�&In���۝�-�j���1qm�KCӳ��ݸuO����I���h!��;ʣ�Gj�RA��o�N�fl�`g޿f�T ���m��M��#]/jp�����뛊�S��B�
������B�W^;�����ٿ@�E�JlX����٠A;ݢ'�F�C��9q�FdV!>$uve�,�J� ���Ͳ��<���}1��ܪ� ���l�r�Q�I�����p� -� �b=Ã
��s�����!)q
��O�e�F�'�
=;�%�P��}�;ɲ��a{{�W�v�y�x;Ak1�ꏁ�5p���SY�{u�`h۪QD��dTTڸF�J����;���s���ą�=-��:v�2<w��6慄ͦ�<�D�h
ͻ�"�"a#��*�X���Kf��r̕��I�p�"�y�bb�n���N�5D�5xj\Lc�w4��=�������oqs�ד���d	ϫ�$���mn�W;Vs�xQ�*j��C���G����ȝ2U�h��7/��=m�� �NO<o��A��Xqmݨ�b4ֆ^����mx\��(�J����4����7�Z�\���/��	�4���J�����?.c|V$ߕŁL�-�\Ҵa�3��:a���6Y[[q�[Y������>�/lFk�}��z����J<u��Nu��y;Y��<�gt[4�4ol̶��輨�n��yG-\;숹|i�!�NF�a�n3��ι�{���B��Pn��[�)��ot�ݲ9��~��A���K�_k�q,�M���aEDġ����0g��t%e`*����&���/�d�Yu��G�n����t��0jZ�EV�ˈ1S�C�';֡BXӜ�+�e�e��Or;n���onV.^J��z���3��Yi��Bs}�%�
��K��y�P�����S��Ԯy|85��O%���G����;�N��+���u�Qk�9�)��f�D��V�K�X:�2��c\s;kw�\��8��t�����h�z@�� ��0Әx���%EV���ԥfR�pV,�mA�"�U��[���,�m�U�E2���j"�m�֣DE-*ʕQP����[-�R�f1VQ�*%-,j%Ac%��R�YV1J��(�Yh�EkQm�Fֶ�F�eU�+.Cҫ*R�X�j(�E[iX6�S-#�UQQc-iV��-)Z���-ŋk��WX�(ҍ�m`�" �KV����*T(6���F�R�KQm[DiU�0RҘj��[VX-�k*�k�*K5Qh�KZ�DR���Z6����E��F%Jʕ�U�YQe��*�+H%k�`�Q��jX�*Z��j)3eE�È�"(��[KR�Ш����
�-�(�m��l�&mK�TPR�Ճh�ت�+*�mF�PDc����Zд�EE`�l�����)�A�QqhU-�����
�b�j��KjĶ�J��*LU�ڌUc[mb��%Q��LP�
�YF1�AT*�2���-*���J%�Qb�#J[H��R�J�f�DX�X,.-��U�,J�(<�����k���r������g�/�
�8��u��m潼�[/�<*�t����%�;�f�m�I=y�i%����ͱ���2\�X�򌌇h0v[��w���C���z�<����$��E=vz�l��#f�NWn!qrF��l���9�%a�)ς&�V���Y#�v���9܄��t��6����Y�B6�u�<��u��ɺ�0��p��v����M��^典(�\4�v0@�λ#N����l����Ѷ������K�zv=�m��[{P���gYe��	�h֝�|d��*�{=�L�c\�N��l����6��G-�ۘn;�mІa_���ݻj1�n��a[$3p:t�^�S�j=�d�����M��ݸ(���}gc"�]�Ԯ��%:T�;1<O[�G�8��"n�`�t�d�>[�d���Z2q{z۝n��6n�n�f�)�.ON���gt�C��W�mW��7�ۄ��ِ|�a�rqQkw���;[���.�[�5��z�Bi0g�<���ݸo+`�W3�S�nޝۤ{���R�{v���X�I�/+9���%�4lf껖��u��+�V˻vy���8:�ܶck�����-\I���'6M���=�s��q�g]���]�nlBu��ԯQ��x0�j���9�8 @Ƕ�a�����hz�[��[��g��ugCv�Z�
��v�m��{I�1͸3n�6	�G�-u��]lij�a�û*��%ͬl�nn�c���'c!��=�:��]����nĀHu]Ӳ<�:=���x�/c�z�*�c��NJݝ<��ϲn�t�<p�S���V��֤��(����^��Az-�n�Ύ^vB��K�
;9<s�BE�=M�f8y�1ûv͔�A9�۝�z.(��e�&��E�=$1>(�ੜ#�v�Z<Ev!��v,qНzy��5�P\�I�:";		De+RVz{k���{mvլ��M�Ě3���{��޾[o��1��n��.gl���4^�cx%U-��(���x5̓�h7�6�������vϗY�0�n��^�v˳y=M)��\Ek��i��5�ݱ���;<4c�Z���Y��8�m��'��������듧��V|�IåSuǂ�&S������-ť�N���unl9�dm����x���I��1m^�qn:��4�mU<y���yݘݲ��Q��b�[��u>t����P ��g��0~L�(p�'?�iH r�o��萮�t�gޞ�:� ���@�Q��Bl8a��O�s��D�l�@�Y�|WnM�A����s�+�>f:V�|����1�1iv���$�r�> :ē��㷷���w�U�A��^D8m��&�e��S�B����0o�zh��{7�k��w"�L������s$��]U�C��wd�UЫ�	P;ފ�8��:�.Ւ�������%B��j����v7^nWt�)��ъF�}"ީD��Ȍ,;�����li�x���e����������lǡpc�}�D�w����H'�r+����)�י	��ͪ�N�vТ"ϝ��ػÄ��<yo�>~���M,������Y��gX��N;/�����)U���g`>]s���%���$���s���K�:v�\�u������$=�����(���{�آ��7��H��+owt��[�c}�7�M�6�a	y�W��;Ud� �f*��s�tHowmxP'qV)$6�d&�A��H�K�j\��+�3A��P�i
�ȬRO���[s*�;�*t"A��|���C`��Y��=�A$�_d�+�2T#�Ĉ�DWU�O�b�I Ƽ�k�3��m��|�JPMUU5USΤN����.�X��G�O2X���s�':9��j���a.�J�DC2��A��DI��ꣳ1�Bf0R�c���>݊� �6�1��#+���I�ھ����0�E��z�@W�~J��[dJO�T������jvE�5!��3@�[RA�ɯ�7�^b5��X�(�Qt��f�i��糳�Ȉ�Q�;NVM`�*;��<q7
t�:��q�;W�2m�n��"ו��?2�3�z2q�폇�  ���	$wEb	���1=8"a�[h/oG*����`y-h��(�n*@P~�������o�k���x���q! ���ɛ�$��٘��
Qï7������>���o݀oLpb���J
��]�3����#M�i*Q�L�D<�-�õ;�B��{B�& �$Dp:���=Yw�D����U��E��..��M6��Y~�wd�UЫ�	������tY<8Z�LJ����>���F;�L�z�e-"8·
!��a����^����(�k����u{��t�H$���$��tМ�e!���D��m;�����������$۹�@�$���RiOi��SoҺ"�6\y��o֍�ZF��x��Yy��ul�0�gg�}��7C�e6��^����--���_�5���	!�H��?mQ>�rÆ ��B||��$��=f�d������H]=<�P�$��~����z_�9�r�0]�γ�]l��ڍKm���Ad��L�NR�ޫ��9��w`\���#����$��Κ$�r�;�ƶ�s��=x{fͯz$>'�{s�Qp�����0�1j��A�0�r"���Ex�O�{9*)�P�]�s��1�ߌZ�
��!%pT1 ��j�T��׉;��c�]=t�X�;�m4�GOn�U>�����_�E��D&���{�-���/7���^J�|�P��|O8�	�y>�jm�'�Qr.@�jl�D�ԶpAH��hP�H��	�<���*�
�<�C)�]��T�g�|�S���.��1!��5�
�w;u�lyKoe�\F�+��G���[��
��]�4yl�Hw�Kst�t�� �����.Tͣ��c�.L^�6��v��
�gi���3�	Q�m��t܊m�N�NSo^K������ۺ9�y��}�\�1�ii�0-��lqsE��n�M;��x�6��6�ؠui�����v�=o[�;O|��.�S�]�>�s��X���p6���^�Sӓ���ɞ�tl��Ƕ�9�wJ�Eضm�=m�Us�n����8����,�v�n%�簩����؄��ۊ�s?߿���ƞ��Q���=���Nj����μ�3[}yиh1[��f�nj.��J�3A-����	�e`��K���� ��t =:����9�cOx�~�Ӎ�.G��DM���E��ںOI�� EtK;)P@xﺕS�C�����Iv1��f�*v�D�W �U��0Er��$�v�2h	7۝TF✠|F�f�$��q	��B0���u�
#{��R�n'�%�{|N�U!>'/3*� o���I�Z�����
H��`Â�`' �]�w&z����J��i��ybX��~��~�t�p��7*DffH�O����bHs��Z���w�(="T �z쌰�\4���TAu�]_;٘� ��?/=A�xΩ�I1��(96xӛ�x
��R5u�ws�/�7�A&<x��79b\z�ٛ�ykRy���{ë�j�ē�neP$��s�A͌�}
�	�;4��ЭÁ�����3�T	 	:y|�yqG��m3(
��*_x�}��(�8D�%C��`�j�{#Tj�΄��^$}��D��Aj�����#3j�)��I\A�A_?*C�]�=�e+�u����w�&�k��%���t��Zf�v������E9�/�P� ,XZD��QQ0�om��t,�=j��p��(9�W���~}����F�kg�'�{����1U�=�(�QF�k���y�D���ίQ��qՒ2��	|:�-��J�Z]eř�N����D�j�D�<�.�߱P����W�n��#�x�#��D�؄\90���aS�kߴ�q%�VJ�ÿc��2lP*Tk�ܹ=�������H�7?�`�N��2�U7/����oG��f��'����G���#/oa-aW�UF�WR裦?g�����������A`HR�����h�R��y�PöJ`v�X����AiDPȲ=�Wd�"x枝���?����S��>��'�+
°��s�����q
����{���������Y4��FT������8�px޼��J��2-ٖ�Xg��t�dx<	 ^��"�!��U;v,l9`T��k|�N T��'�g��$����}���F�uo���I�5�D�HL��D��a6�^a��0WY�OC��ɺ:�e�c'4�����\�oe������§3��h8!ĕ
�YX{�s���,���@����g��쎵�u��y�i
Z~��}�8r�R�l
�~��&n.q���.M�ؓ=��q9++%f?/�]~��.����������IĂ°�)�g��0�c
��
�����G9Y(�����u��dD��#응�Y ![C"">jnrf�����q�4r�RZ���hx"��E ��"sC��$G���q=*P@��߳��H(mD@�~ݑdx�{�b0b���|(G}?d��7�A���*E�I�*Aa��|�0ɱ��@��w����+R����e�����co��u�=�3 _�bL`�\��R�:�^��Z���6�@�ԥx%|	V��S�	L��6<%�R��$B_��!Zk���Pñ�R�7~8�-(� Y��]�,� *Ae��;߻���8�N�7����zN��°��}��6¤�O���G9R%�*~���D�q�1��ϯ����v�c��ړB���鴺6�A�7��h|��o\tZ��r��4~>�\�E�2�Xc�k����!e�-�s��H)l �Y�o� �,����(�)��c�͂k���$6$�T=���H,91�=�o��g,q���paH���@�������U���|C�F�e�������AH)Z3�ߤ~��A{g��l\��>�s0��J\�L�\�1W6Si5�߾�Ă�� ���}��N$�a~r��]�٭s5�x����a�%����d���FVKS��w��֡\$��d��� J�!��������ǻ�^���r]{�����s]ѿҐ� ���w����@��w��u1�ǽ��{���0��R nv�>|�_D�؄�ߡ�B��
�{^�T+%X7��E�}��D�߯s�ɂ��ޢ<	 ƽ��6�X�����')�x"�@�w�������}����6b`�0x����P�u��U�Ȋ�/	=���c���n3�N+�NX�
:S �)�2:3k`(�ʞz�ga	���n��V�W�xxuz�(�0��3˺'bqQ̂����9*xr-rR�M�um�z�E��7��	�ל���u�86s�^t���X���eN�� f�َ�x5n����oa�^L��,ApnW8��+��n2�+̼X5lM�ܛ��T���ܹ�vc��Ya.��wm�^l�uY�>�qvG�][&;g���m���Y��d�t{u��GM�9�T�utqʬ���Y�7i�m�ا<g�:#���n[����N"f���{��$Y VQ���~�q'�+
0��v/g��$yoN�2��'���q���������h�N `�-�J��2-є��c_h?9HYi����/8��=�~)
�h0*_w���N*e���jf�%H���~�XEeȳ�����W�n3�\c.��aSy���r!Ă�YX?}��7���R�k��۳^��oz��`~k�!KO}��h���B����i�`T�����q��
aP�Dzw��FT��:��Ǻ �8��d����tr$�AaF����ۆ�m�Ib%����tq����������œq����;��D�q����\cٹ-q���$��z��B�<	 >�͑V�N��b"������s߻�8�
� VT����CL�%H(T=�~�0�°�����n�_}0) �0b!&��E�䛮1��,�/��=���1k-#�dV�ê��ϧ�,vr��3K�,<§�w}�q$�
�FV}�چ�
Ĩ���ݜH/�}��a�ڮ��;>�<>�Cgo� X�A������چ��
�>�����2\.\]�����>���ed���ԟ��L���M˥��lF�N���U3$��H�U9aͭ���>�Fd����I
���H��-���2��;;��:�/9��I��;��?�q ������I&Щ*{�߻���e>���ѓ�O��׏}�:��G�� �B�WȷFR�t�ii
����to��k�0*s���T��e��~���T����CL�d�PIP�}�~�0�0�(f~;,	Cd��xY�����.�~��?�i2!Y,e`����i�c*J�O~����A`q�
�w��@}�߽��k.q�d��B��{P�AM�'������0�  �#��vȲ,�++%ed��{��ȓ�?����.�a�°�����i�� ����w�8������Xʞ�����y��ஜ���A�4K�)�A���]3n	N�9�'֏3(tc&����?���E�B����}�����!m!m����)
сR
S���l'"G���N57�y���>���>}G�D� "ݻ�,�|/�Kb�L2!�E�T����8�Q
Ƀ�����������6���֎3i�@��߻��5�F�)i���h��:�:��:T��;'�M��B>ߑ��K�4��@���4m: VX�Yc%O����H)�hGY����x�,���\��K]��[��Woj�Q�5�aP�����Ox��(F�ѝ�(dw}.���q�B���Ѿ=O/{�g��L'��4��}ȑ�SaUC셎��7��nggg�{��^!�Ӧe��q�����C\p��)0�����9�Ӯ$�w'N����2�ɖ̗rb1^�0���9G{�� k�W�f�M��Po���9:��j��������r�⏪]gtt��=߰.�ۼ�* W�#3q���?{U��:U���!ݾ�)�1�W�|�^��^U����}o�>N�D��{ȥj֒�dO݇j�����F�=0>���Wr+��]��=�3��jYɇ���\�N��ɠ侂����R�<MS�}97�v�[�O���ܑ�۫���q+�VZcz�x��/��g��}��|��StM���"��#sg]h�J�je�l������{�9;Wܟ�y�a3
˽�P��B��"]��^JI�4:�tlq|��;���,�Oyr�J�Ǘ�P_Y�;��Yv������_�siU�,�=��;�#9u#Ҟn�j���c��Y1[ǭ�oVp���l���у��\�Ԟ�7.1� �W�0�t���9����I��#}���.6��lc��L-���|/���L2�V��9c73�k�^�UB�=9�������7q0T�IWc�w�u����f`}Ȫڀ2�G��)Jy�;����3qǢ� �D�,S�q����'Um�6g5�Q7�> ,X��Qb���k�x��"�	c
¢(Ŭ�����ej��AATŰ���ȰPX��fe0��ͪ[UX���E ��*PU�\YX�-�R� �"��"֢������V*��A������*��k�eIQ��$k()RZR��TDb2
Am�"*ą�TV*��%jVJa�)X6ƥb%V�+�a�g2��E�&Y�p2�KKm�����.0��(�"�0��b��q�a����D�
b�س��`ZPQU�	�ҫ"�D�
�X�q�E������((�X((�ڨ&[�p�kd�Q8�U��R��(Ԣ+-j�UQH����d����j����DU����Q`�ŦR��UQ�q�0�"���)��D�1��Qb�ʕ
�⸨Ȳ��	W*��+5�a�m��-�Qh�c,Kh�ca��QX)X,�ҋ%V*ʣm��2E[jł�
Դ����E��UTQ�������me��EYE�++ ��c�{��I'�%��߻���eH)=߻��6�Ƀ���q��K�d[�L�����~0����Zrb��x@Hx$�wH�B���R������q�+,������8;d����"�@<��H,9�~}��Ÿ�Fcw0�0�����!Ă�YX=���n3l���:��q�}'�q 2 !ϯ(Y��X�i���)
���~�4���Pj3�ov�kXTT�R���"�7�r�Nضa݇�/Wh  2��]��.������m�ܕ�q��a<�]��tq8 VR2T�����q
�������T�N_]�^v��a'S���h�'VJ���;�����8�Ϸ�Ìw7%�3�ctm �q���4��i����Ͽo���wF�)
�Z����h�*Q�w��$7T9��O���#�W�}o�>�/��b�q��q�]�a��O��wAȇ%X?}��6ͲPe@�Ta������7��{����
H[O���@s��JB����������_���&Z�d��F�\��s��{����d�����8D�H)�/}�ۆ�m�IP�{��F���j"aU #�YH~�*;�t��p��F���&i���������}���a,�:d�ź	��6��ر!��^�"���8�����	!=4��Y+*o����@�n8�L��E�4��X>�����!KH[@����򐯱����ϯ`i�)����(�YR��~�4͌�
$�{��F��;���M�}��Ce��"��{.�t��CW��XV���ν�J�������o��\g"a�_Cl<0�����!Ă�YX=���lf�+*A@��w�6��X�x���>�Ԇe�9��@rr�RD/�����l
����ni����2h"���ݲ,� |����c���:��Ӊ�k���	8�XV���y�p��*J!RQ=���8�����VO���v�{�#�5R=�� ���#�c�n1�;8�X8���u�B�B���}���AH/#�:k��y������3s���N�,@���چ����bJ��w�Ѵ�Ý�Z��e���Cm^�G�;�r>��l1���q�H,��tm�d���P/}�{��`Q�>�������w9?k���ԅj�׵;`T�>;���.i��8�g���8�Y�J��Ȍ��dX#�@w_�o;-��^>	����0�aRT*J'��{������S����8	��~���s�{#��ğ���շ.�d��1c5+��j�aʲыL���s ��s�/޻��{��̂�r�-�ɛ��9S�w��B1��ڵ�8KqpY��n-7nԆ�g��nӎB7mi�q�NA#��ε��آ����^����?;���h�����.�*V���Y�j	).lo=F��K͹9Ϗ^�D7e�i6�h��lGm�ʼv�Z���74��{&����1wg���Ɩ����g�עH����1�;A�;C��NOk�����̓��s�]N�Gontv��e}&�y.��������J���e" y�kv��8!E������z�3��R����X?kh6�!m!Ih��{�i�`V�
�����N3�Yu��Y�� ��\��3l� �P�}���+
g�{����G	���r*k?{�q%���{��9��]׵����߿{GY�JʐP,���vq ���w�w@{��i
���K�ǯL����چ����x�ni���\d�M�����8��e���2T���r$�IXQ�a˝�d(��؇՞G�#�@D�v�H,�����>���D�N S���G4�6�(@г�,��_u�~���{}�}�AH(?k�6�^�+FJ{�����
�@��^���3ڿuf�q��8�@D۽�g�ϊ����ˌ��.3���T�����J�d�+��FٶL|���}�c����_s�{g�`Xԅ�������)
�����i�|"�o��tO}�ᦋ D5��=�P�v^��s�^]Au�A��to'4�;��}��N�����|P3���H,�%e*~���$�$������i��&���=���?$�k���H,�ed������� LN�(��d��'��5�����i
ZA	��|}����on��׈��B���zX9���*�Ă)��d��<؉��V�ݢ2v:�D��F-�:�5�����&�lϖV?b�t��<s�HI$���~�o��+Fk�?������r T��?w���l�
����?o�dn�t7�sZ:ã
��v�����1�p�AL�����Q
�c+��ن�6ʁR�o]���Z�g��ǘ�H)i����9H6��?w��;�
��Ӄr��*��]����F�	���o���_��Cl��~��lH,�����H$���<"���|*�sG~��w��x�3�D�;�=dY /_NB�p�.(���Xg�s!��B�B���l�#�����#ບ��J� O�~��{`q8�R�VX�{���c%H(Q~����+���s_\}���\獜�0�cm�nm��l�4�û�)޻i��m��6.��~��Fg�Tv�{���*}�~�AȇQ
�c+���f�+*A@���~��08�=�����߷�WA��ܹ _���E;��;`T����;�SK�7�@�u�4Q#�#쮹���������z�s��G�8�IXQ�a�s�a��*K����ѶN2�X�ɯ}O�X�}kqL{:ހ��&��q��Ìc*cf����rv��������to��G�(�A]���K���hR�v�"�.�x�I��ߟ�.n]��?�����Sӝ�f�l�ٜ�B�R�i��5�Z��N��65
�{�򠭣��{���Z���AH,��jg�%H(߿�wF�q�aLk��1a���˸q �q��h3��k�N~�?�?VJ2�y�~ѱ�d�*J�~��wgk�R��~�t�c��}������B��桤�����+�L�Z�˰0�I���h�q�VJ����Gqk������V�&����70�aRPB�~��q����Q�=߽�G��Y s����&l�$�Б�Q����W�842 (��F��۴a!�&�ę�e�����!�����`�|�(��r"
B������7�HV�*AK>����8�S���Ӝk_�١/�ߵ3q��RT*�}�a�aX^��]���pe��h��*{�����$�
ɞ�;�~��y���m��k���
A@���ݜ`q��S��ߴ���t}�7�����9��COX
���8	�4 �/�{��$Y�R(�S�~��I�*J�����矟�����j����~�*AIS�����N2�J2����h�N d�	�D0��C$D�>�(��� ����1�|��i
Zu���i���`T����l'
�����?jg�G�Q�w��Qv���3ni8i��Y)����T^ܲ[f7ui�s��r�ѯ@�����OG	I�	�/�� 
a�~�mW�����AC�C����Gr0�,Ƽ��p���Ŧ2�a�5�~�I�
�A��߹�F�m�;3��~�9�3��D���o�`q�
ԅ����@m ����*>�R��=�&�Y?B�"`1!���*�����v��q��S��w�;ۦPs�_��߿v��rի��	��=�N VQ���%O��~�ĜB�+V��?n|(G���Xѻ4>�����W#����������D�q�?~�c�Ɍf�pavq�����4�)h��,}�� Oԧ�k��"��x"�|h��}���`q8 T������I�@�"o���E����������ßo��1sK�-�L������t�AH,����J�D z�N������O���A!����9�A��lB��?jH)�ߟ��@a�.��d{���GXk��U���}�k�<��J��S|����N!bJ+�y�P��%B��}��ȳ�������o���|���|��f�G�� ���H���DD2C�'�P5��o���ZB��9�}��HW7'��N�Y�{M=�s���*Ae�~���3c%B��Q{��,�Y�G��˔~[��B;-�Xni��t�yoy㊂Tl2ukR�nُ�/��$R}tc��]!�k.��f���P� �3�d���w��^��:8؀x�`�m�`�l��c�'�N):����[�f�,Ū�5�m��JN(�#����,u�.ݶӧq��(y�k����$�q��1���M�'���=��,V֔�����nn۰���\i�� ˻-�ח�����g�x^�׮!i6D35��O/m�<]r���
`�v������kv��kn��sϥ�c���z"#y�s�a�Ry��=��8���&7Vq������!��|?������!ĕ
�YX=�?h�6�FT
%@��w�vq��k��9��s��i=�o��)���s���l
��]����rѫ��	���߾��Y #�}�}�q5��~�?_{Č�����N!RV�ao}�ۆ�
M�T���ѶNFVKY=q����>��u��#�,�-�D��0`A2(�8�~����B�H[@��wF�)�� �G�#�6�=�g��۵�| �9*X�Yb^���3c%B��"}��,�X>�/oV҈E�j�j
AO{<�A�}Ϳ{w�:I�+%e`��P�&�P*T=��wg|��C��� l|n��s����o2~ B��9�i�`T���L8����p:h޾捧P*Ae*~��dXz�>��[��G�>�w^�c
��RT���d�+%ed��#��G�� [B'�}58���pv���	�u�S�s�ޓ��do]rZ���l`�q3��B�l���H	>⏁�k��HYi
Z;����
B�`V�*_w�w`q8�Sx��u݁Y���jf�*%B�{���a��aDV�6Ɉ,BB�>�"_}����O���W�T�3q��3�W��b���]�맣�ԫ�����Í>����zV�SeN-d�n���T������JUe6��[̘q��-t:�����M0w���4��T
%@���wF���������� Ф+�n���C� S\�I�| �u��y6P(�ˠ0�k�~�G��2VQ����wGq
$�(°�s����)��b�.���$��bs��tq����������pN ^g����w9.2�`A4,�(��rI��G,���<�-�k}���HV�
�K߾�v
A`��y�i��wۻ���I�(��D7���$��}��+��f�.pXm�O{_��q$�VJ2�~��}Gޝ(���3�@�2���`p���-?{���A�(�Ex���'�M��ٙ9�D�&s�^G�cTF�뛠�e���=%�U�z}�]�q��m	j�8l�s��za��L83����>������
�YFJ���w@m$�+
�����4�l*N���~Ͼ�ߎ��0'>�ߴq��� �VT��{�'�����."!�	>�>��|$�ݤ-�1�k�\c�@�5���AH)>�����8�S��%����4��D� <{U���+�_q�R4�|2+
�m�X��3^|,�"%��h��B�Q���}�P�&�R
p������&������k����ɌʚŭM�T�E���F;�V��WK��^àI�?e�X��o��u`�\E���4�n�ƭ	��v���������||���R��{�����؅����4�Q����Ĺ�F�r�'�&���q9���>��k�{�0βVX�S��{��N!D� �����p���*%O��wG=�������]�d���c�F���Dv��l(e�	�g��X9��h6�!B��~��ѾR�'�oq��� �Bw�� Y�J�Yb_��u$6��D=�dx�c{WúpR���i�`A��Ol�z�[n�z��)Ӄb��1h5��V� �E��8�CQ桘'�	���"/쭐-$� �}���i �l�^�ohY�Q�b�!N�1�x��$?��@~� �B����CN�)���W;0fch�'"Os}��� ����<~�}�=�0��5��	8�V�aK�{���laR
J��y�d�+%���Z�����>��5����8�f�鴑P���I�
>ꮐ($-�-�s�s�7�`V�
����׷�߽��m �v%��CL�%Bĕ
���;���1��1��8rB�>|?}�h�K�u��%c��C)?D+%X;߻�l�%e@�P?~��Ѷ�+R�������z��fe��HKJ;����gv�����I�T�`y*���T~��!�\m{%��ݵ��>S���X��$Ьō���GosB?�xG���
��������J^���13��5s�`a6�^��q8 VVJ��S���I�5��z��N0�F��;��0�¤�%Nw��$���R3��dz�@��?I[�tw�@����}�㍋s��������Fp{iޤ�tn�a�!7w��|�(m	�i�|߮a����}������
�K?}�w`q9*c;����d���|��s�CL��P�*���0�V>����#��1��]�H)�����q%B�k~�܋���}ײ�y�wP�'YR
���wg�R������R)
�����e�^5��چ�
s����L.f0f���r$����N T���S���h���X$�+
�}ֱ��~��w�^�{���F%B�������Ad�*AO�{ߴN'�YH�8q��I�
>��@]���銎��G�Hx$����(�x0+FK߽����
����ݟ	>�IV�Y���}� 2<�����0�0�.7��:�6�L�c.��aS��h8!ĖVJ2�{���$�ْ�zy-̽���H{��z��~)�F�-����hNR
Aj�w�A&�|#��Џot\� n�w��\3�e;3e�"��]�%Չ�rN�?ah�ǖ��s��Úh�qUS+�= �`(�� ����I���`�"�G�m^���wv7.wn���5u��:X"\��Ƿ��n��íq���ą�����!A��P�z��'����B]�xN�;�v�{�灻سN�:_ǫ�f9,�
e�r�F�JJ��r�C����P���|Z�n�Z�⬽gM��m;�+���V����f]c�h��:-#;��^X��N����ɑ���F>�6Q��΃:��l�����KY���֛�⛽ˍ�',O!���H[ս���UiN�)��5:�&�5�d��O�@�l�}}��G!��*�庵�C�w�������-z���%:��7R֗7I.���,���2��H���b�Wb��c�:�WU��z�)�wWf,���*!Ǩ��v�>�q⮺b>�kߣvV��R��%ي��T��eVf����>�++-�÷��s.S���@��т����O\N�/_��[Gyɝ�N�I�52��;�
}w��������x.���\O�Ԯ_.�p�AN�o�������jZ��kZ�7(L(n_>͕Q�W�z�kU�=�-Σ�qC 'a��}�;��=�n�s��_�N{�|�s���6�����`1�Z�T���[�c��i�A���C�"Y���+�w�]�f��fO$../�ߌ?v-�a=�dCf�WM}�` `'�2T,AaR��m�*����(���*��!PQ[J���Ŧ��QH��,�*TR(�"�,EJ���*,-J�Jʑ�*B�p�X���3kI�Ve�����jEm$��QB��QJ����eJ�V�J$m*V�Q�cJ�Y�\QIik
����,��0�J�3J,���R�����TQEH�V�+Ukc#b%��m5��Z��B��eQKl[eU�*+mF,UE�T�.��ʳ�Q1JQ�,`�Q��k*EQ�ږ�V[U+QUX���ͫEQ(``a0����Y�B���T2�[[�F(�U
��B��Vң*�
+VDb�DDR�"*��#b�EK�U+�V
��QA`�U�kkE��T`�%\"��V)YJ��QYm*J��q(����T�
VJ��,�X���R��UE��bW3lX�V(�b��Fdm7����>2�,G�	q�^L{,�<����N8`��'c)�8i5�"�\9�a�	9�mK�1ʹ�F�n��:oK��쇝���;V�xz.]=rt;���q���l����cq7ag�km̝�㗘%�͵��6z^ۃ6-��\��}j�]Q���{;qv�<f��vz���u���MJ��|M���#���g� nݘk���9ᱼ�tn�b�n��q�zݓin&��y����|lkwLEu�N��nl��;(u+ɷ/<�:f��������z4�Q�&�\=c�]����Z�s.�ŋ9o;u*u���v�k�z�cb�Ŏy�ob��ѽEy��`H�<���G ��q� .�۟;9��qۺ���t���Zw�,���DKj��i�ն�&��!����sW��v0+�7��_���N�㝋������Q��j�5���W��r�'J��v��;������*�ls���km���yݬ��FG�+�0m��x;�d�;�1s�n{%r���L"X�=�۲ݣ���wg��3�=�6F��9��[�����_Y��q�㣜��58m�UT��tx�c�mۋ�Q�U#�*���R5�����Y5�8�e���-ٸ{�N������<������ч��9�銨�.l����M��ʒ�/i��([�=�y�;ul��;&Ŏ�ų�U��C�G���p��u�v%4l�ͷ\�9�m�s�ݹ��˟;�ʼq;�Wf
�ۨ�c>��\�=*����I�>�9��mg�u���yQ�Ok��g=�\�Ʒ;�b�$.��E��d�Wn����nہ�n�s�J2؏SՎ�s�]5��3Ȱt�э΍�e7]'>lN�^�:8e���g��Xh�s6~+���d39٫q�f��-��e��=Tzx�tj)���6���i3����u=����5k��Q����齺Ë�1��3���.ԛFy�j��i�V�Z�L��ź�3��76�}��:����/���"��G��F�����������{|��ܾ�8��^��gq��$�s�뭕��/!k�����:v�s�9�t7d��滆Lp�I�ݛ(nq��Sې�l��Xy{]�ݍ���p)��Ggy˃����X�����m��v��;����-�m�S;���7�;�Kr������=è�^ٮ۪s�2�n-]�M\q�d�`6�qѮ9(� (�e�l����;�v��n�uW5KtS�#sx����]����\W9���
H��%j.������8�R�r��a?�I���tq9*AH)�����8�T�����w0�
���v� {:��6����FVJ���{�����5�-q���j�����`���A��B����y���}����~ѿ�B�`V�*Y�}���8 V�ﺆ����bJ�}�"~�����|8�#�;���G��1��]Aa�>��}��!ĕ
�_#�˯dW���@�@;peG/�:��s�~��:��A�
ԅ���}���)��h!��u��߾�~ ���2 �4ﯯ$Y������/���Agђ����4r$�IXV�c�wp�AH)7��{���߻�?����Y+*o����q��{ų8��3�d\��ma����� �-���ȫx#x��a?��r�;�Y��T�������AN V��u3l�
$�T>�;�a��a�c{��c��̵n�[�EB���TJ�A@��	���v:�C۬�u*�e�onf�zz�-?������k�����
>��_ݓ@�7�ܓ�G�Ve���쇵pr<o��wU�t,�Dy�!KeX}[�D���T�Twm��#�(���7�i�������"�w�H�<Z���2�^7�^^R��U���q�,-�74�N�����ҿ�I}����{|Εg����ؠ��,k��n�������j�]� ]X	|v��H$����>'ǴZ�\0��Pq������yV�H��ʠH��Q��&�>��f��N��En\�A�}��@	=���c�[8.|�s��Ą+y��	~p��S�TO��{*�����&*<I}����Mx�Gf�Ur�͸�0L�D 3�dGF��-��d�C��M.9`V�(]B�YE��7�J�CNC���s��$Mv�M(zw�T=�o��\��A��f�@R��2n8�E�a�̈[՞A��1=Z�s�⁣�S�A�yB���^�Aӹr��s�R'���'��@f-�!���I��ʢΤOn���WǛ|���[�k#ҋ{nXx�#8?���{z
�aݗr�cZ��͟%�W�v���X�r�=i;��\��{�#��	&��ʢI�~�j+`��pl�	�F�+�`�J/`";�nh��vU	 �U��G�S�N3YT	�^�i���m�譜$�W#p׆�'�|:��EH��z*T ��w�`����N�q��w��0�t��+��6��@ݱ�|���/=�U�=wU��������������B{�y���=�  �yW�x��$Uy�ʕ�\��A���-��&Ilv\�.ڝ$	����A��r	 ���&�%ox��OF��8B�z��$�W"@-�5�^�篗P���{�* O4���,8M�ʐ�ojv�E���N�D�W��j�
���j�{��谠R\.$�Bs-�)�h�/01�m�ǣ.�ȉ�q]��{���C�+�*�*�Vv�8g5��|&����v�:��ꂱ�\�T�V�����+*�E}|�&�&TD}�䏯o&�ۛ���S��
� �'��]��B=���(�笺?3���H!%�PH{uq�T�͓������zlzM������������e6��lVp�}�W"H �켪�E�C%�O��>$!ۅDF%�2�5ӳS���/rQ�B��ؠIr�m@WyH�:����1����Y��K�Cq�-��$	�unMI�,S��b���H�ʷ$�7�2�pn8�Ma�̈[���V�t����3 ��[�@�H;���/����l�	5�IZ� �i4!a�!�v�Gwu�5�-���5ï	�ӒA̮ɢA>=��B�
�h�\R�
�N�����#��9���~�g]�
��� �o�/q8�������LË�{���g;:����k��=�{���$�i�A���!�0&��m��j�����]�71Η��&�u/	�C�u�Z6��=jʾs�i}/�%�w�\Dv����ֻcsB�n�dۢ�]u�o)��V���eQ�q��Fpn���|��N�;6�J�qo�>:���o`�εU�gZ�/m����On�����`pe7^r���`����n�,t���ڜ�^ݸ��'��7�sm�nv��U���m��:z7F���·[nJ�|v�:�ɴ�4��S�go�0#�6� ����rH=u�5�I'ۛ�Tse��[�"#5׈ V�eP%�z"�@�=����iP<���0n��v]x�|;����I�ު�@;���Fm���}o|P��	`�_�-5��t(y�T(��bsZ��N�y�$��ٟ�ͪ�
�)���!�[�F��αSS�����I��٠A3����H�n�$N����@Vn�JFp�3T\w]Q$�ڹ���p�Uv��v&����T��̫rI���!L�:Ѕl$J1�Cʈ�P/A��<n��"�n駝����W���}��=�"0�<���|I��A>#2�όl��u��=��TI>9��TT��5�M�D&��2|�ն0���#T��U�����&o����tD���{���}�!�iz��Rc��m(��t�w*���%���w���fm��ĂA#w直�Fec�J��j�df�{3.+EFk�i�DC"h'��U�Y#�@$�Z�c.���}�S�2��>C�
� � ���n�{mv�9�,:�E�L��U	�w��A��\}��_�]�N��Z�H��I<%�k��$]��z�9�m����%Dt���mc�;��k��r�����o���=;�B�\q�F|�t.%�Z����i��8�ƴ�FL�������3q����=�D�3�$I�뼚s[Ƕ�1QљF��רuc�9�a�B�yGj���T ���-ϳ<�J�ֵ1����:��z�$QsYR�L��f����h�Uu4t@�pl	� �ݩ�H5�{4A��A��$ہ�\���uc��o���ݘ�]ۓ�H��S$�W#��5��:���sZ��Ay�Ä&2��&!<��q�P�f���j^��${k�G�^eQ -��dDC"h �;��������$��̚$}����Έ��p�I��s�B��f`�p���[U�9��B�GS��9hb/��|H���	�{(T�F��Ͽ@��~~��V]q�oN�X��h�5!������f���uc��ve����]�J�K|�8䌽̚�E��P=�c�܅hΗ>$�ٕ@��*�(Ma4!��S��2�ror�����]���%@A��ʅW��y��3�	��BI�ЄA��ۑ��w����	$�D��^Ѳμ�G$K� ��ދ�(�#\�	�j��ډڌ前�����`���P P��M@
�L�Swּ���x=�j�~�d���q�9�����6�%�ݽ��I����췋ɮ(�in���f�{h\弩Ka>���Ӱ�t�c������~�����`��dBmﾊ�I���e�<ʫG{���a����
�މP�H�Ij��bSݗ��eFCf
���l�Zrm 릥J�蹵k��Ǝ�g�3�'����Tr� �L8A[�9<O�����I'1L��i;v�4w<�%@U
��E�V}�Pe���S��>�= ����?F샦$�����ɲI�#{{*�fU�$�]n��YW�R��/BJ"i)�����@S���@	G��������Ѿ$��@�s*ؐu�%D��@ǌ0��w+������)�p��H3w�@Q�$�{�܀I���-��7�r����4,@�plB&�.�� ��̐ �G��/�2E{�ܒ	ٙT�G�]t#��	vl�C`=�r��N�^Lh:2�@��H��ӯ��� ����`��%�"/��U��w�d��Zc�|�����?�L��W���L��;q��ny�ƹ1=l�8�����k���@�9�t	�Ś�n��[a:B9��6���ѻ�i�qvv����v��X흉��p@`S%�㞭�0\�ۈ�3��t'���qιڑ��
޻hH�F9��֡;�v�.�W[pk�yT���i��^���R�N�6��tw5<2A�!�6�ې��G9�,3����z�7!�l��Ʃ����&ض�&�L@l��nfe,nm�
_�����1(h4�~��H�;j�I�O��2�q"zv��,�����@���V�ġ�1aq	�*����jt��*�3�28�V�>��ʠ	�ޚt ����������;�B!��q
�~����̚l���Q��������$nU��w�2��%_%	�"�3T\od�-eT�F� I	�τ�A={�TI>=�ٳ���Gk"�H9���h���ʢ|I��ʥv���k�c�����A��r	�#3�*�'���oeQ1ћ�-�͊�a� ۄZ$?.4�:�Nh;C��V���c<kG\�g��y�7���߼��b0�w��S'�m�d� ���]��v��G��AD�@���5 g�V2"hTU
���mvv�����z�]�[o�Ƶ���z�{M�ܠ^{{rE�*�PY�-�Y&_M���m�Y4�0Ƌ��j�>��#e�x�nd�>$���U[��ܣu�x��s6��.�`̳C(�4R嫕 ��ɠIv"m��ʎ���3g��	��ʯ	��ʢ!v���%�(~M�[ū�����@P�m  �މ| O+/ncr6��:7*�l�qP�0���f��T��P���h���y��6/%@M��H�I��~<�[���_�7L�݃sx�K�9fّ3�6sm׌��=�p�0�v�Qi�1�.�ݼ�^$�wey (����2{P��+7d��J����M44@��Cn	@��"7j}$�ے����ݘ�S~$㙽s@���r	.7�T���G�j�sI{ɜEB6��$�7jؓ~�GF�\y���:�����Y��1�y&�eæ�^����T	�j���ʵ�ɨ����^�11=����iH8��#�#��zH��EZ���y�^*�o��xg1saR���n5���Վ����3���q�sT�7��	�2��J�#b���x��p�ÁrŃ���dz8͔wyI�^T}������X�w���B��m�ʾ�ڑ¹��g�:
��\s�e�Xl�s�ZG.�.��z��0��<ר�j��5$���ƫ�.�t�=��R�4v�(=�\-t�:T5�#5}���}�X�T�kHW;|�O}�;7���������.�z|q	�WY�t�K�=k��R(9�V:�u+�z˜��(j��憶��{{��{ɽQe2���6g{E���	��󰂶{�>��y�� =�02����^��s��<9R���M)�j\�-٧`�}�0{�:��w*���.��7;�&�3�	'gSb�t"c�M��^ܓ�i�;�]�u�����+�t���=x1t��l!fVc�Rh xV���5/f�H�;��S�7�Tȣڵ2��w�_M8���g�vm�wF��1�R�%���^���c±ڗq�^>��^r8�7$�y�Oւ9�氫=8�Eǐ�:{��ue<�g�V�K/�n�c5�msv�x�8n�]q�vj[t���>8��!�k�_vHB�d�v���� ��M�leѥ'N��hAT̛tQ�h]�wJ$��͗-ŬT"�dTUATQDTbņ,YU���
�Kh#E����U�eV̴F ��B�B��
8h����)EW-,EE[J�ES*��J�V1E�-��

��UDV*+0�QUEr�X���eF,b��V6�0�R*�Z�5@PEAEAU��1EDUT�V��т�b���Ċ�F
��UTQQY�"�� �*��F�A"�*1QTQQ�� ��mQPQUH���U�����[lb�b+DA��-*�U�PEFEF��j�TX�c.P������cYE�*�"G(��R�+D��*�����V	R��EX�F2"ְE���ȋA�����#"z�y��P}�sfß���)O��`̳C(�4R�����ŗ���y��^$yVă�Y���=vU��{-�p$�9�B̦b���7�o,	��j{|���'�P�r@Pry��̟q�c=���@P�-�	�BCu��Q�=��v��K�U���Ͷݸ�����i��>��ۡ'�P���nP�	fչ�{�2����7"���M��H�	 �U�$كLZpx�
C�ݪ^j[��Wl�M�>�MlC�> ?'��^�*�	�.�
�]u����R���@�^�Dvԉ�]nMA 6S�T����U�H9�nA�չU�Hy��EB6�s�ѷ������$�nM I'sk���㐯2�LM��7q��D�shk�*��\�{~�R{\�e��H�rU��/z��s>Էni�0WN���і��[Ⱦ��{��>���9��ÂÄ�V��As��/f�S�H| ��7�B����Cso��qV1�����H�����GM�{\^
ɛL�T�˶�k�$9`V�..�x:r�N{;�PXd��ɾL�����Q#�o��-�y����b|I={yB��G�U��/>8oC/��!B��R���o�A>'��*�I �m�P ���˅�z�ă{")�!� ǌ0�϶����A���It��úd�d�A��ꨚ �lCnE@�1�jUj���1=X55P �w?%T Zd��.�\Puzt��uJȽ�|���I" CA��"|w��
 ����@�v��6f���GU�� H$���^7�V����Ok���QO+�,�;FQ��s�ph*��\��)�n�s7���;��oZ�|��k������&{���كv���5xc?*%������DD@`�@�1ے]�m�a�b:���=]<l���=��C����V�s��U^跲u��6�m�S��hR<��tqɢ����K��=���ō�G\i+ܻ�]q��=s�s���	��nwr�|�Cl㛟n��y�k��g��Y�%�tӂ�<�<���d�v�=Q��n��D�m�]�4v�u��{;�ۍ��j�u���.�]�*l�s��v_-%����HE�Z ��[��9��}��q����ݙb��
��iP��?$> 
r�;C_�ށ�4W.�����@�I�����9�����7>;*r@��x+���OWM�˷=8	 �M�_U�"�	8	A��N�;��NX���	}C/��  �S?00�>�`-;�ؐP���@3�S��ˀc�R�ohc��C�/P�@�b��x�YW����NL����"_M��vr��&��<��i$�M;� 2I��ɯ��,�v�%��R�����>�+��L�Y�y�cu�⛲S��mݽ]l;�\�6Y��eg��z�܏Hl=�������7<Ŋ;w�o��꽧j�2	�{o*�;�n��q9����q긒P��qC�$7*��;iU@�κM�[���t�9�ޮ��Kh�A���dY������
�rm�	�ΞW������Qȸ�����;m�Z��*�ؚ
c��}�D�9u\	'�}��D�&�	�\��t'oL��pb����E�|k��k�����5XI"'���I�p'ǻo&� )���$���j�.6������X=�$��d2	���Q �;�޻ɔ�ݴ����.b@$��0ˀc�R�j���u����Ş��,�Љ�[y|H���H;�}^�'�󶜮���(*�������ά�������65뗱�R��<sP�4�UV6�؆�H�{����׷�@�	$;�J����6�z�����T.t� �`^0Э=�n�B�ٗI��d_�>��ʠMCӟ���!L����W��|D6s���
k�kj���}B��B�����`q�{��&y7�9��e�:E�Z5�P�6xA��D6q�9�R�#K����;̦�\d�Le��;���9��wu�O���Ē{6��Ry��Kp�>9{��z��؞dֲ��:���n�h	�>����g*�v�[�&�����$D�\�I��	�f�.��$�2]��cԥ/��y%B�ݾT�p�00;����}�h�J%��J'r�v-���1��q�)�7��L���2��j������l��(�<��A>;�=@Q'��EZ������~��\�e��*�(w��T�R����&� �h^>��W{9eQѼ��nf� �o6z��FdU� ��ˈ�[n�A"/�$��2�Hތ��O��R	;`܎�12���A���T(	-3�Ƥ�!��,QK�sB����?���ϵ zZf�{����ͣ�#	��+���ջ�cuW�*���:�MV��ZkT������D�Q$V���������(im���ɗ�͋E��z6ٍ����g��~� �U�Ry��Ke?(��O/�"����g2G+�]S�@�ڪ�|N���$�7�r���¹W�[��4`�n맒���gD�H�kΦ�Arq�Sd�l�g�d�>�0R��A4�߁q��{U�|+�}5P�7����<�iP���ޑO�S$��#P�7*�&.�=7=�tﶺ��<r�$�{�@�����l�X�"j�lC���Ux��� ��ܚ'Āg&V�֜Dvi �Zʸ�I�u�U�r$���e�I3�{�Z;Q��;MK@�>2jrY$]y�(�ͮ�q��)�؆��yB��Ah�������$��P�P�ʎ�LuP�	��p$��ܪ �I���/{O%�U�>F,4�����k��s��u
���q7Vcn�_n�����̮qOJLMX7����w���E��e�~B9���=&�2L��qֹ��;l��� �c�Xnv9�;(�\-�̚�0�qawen�O����p��+�v.a�tJ�vԹ�6�s��rq�W���jݭ���1֑��� ָ�h��77n�nf�2/]] X��i]��RGtI2p;:]twJZ7n��r	s4	X}�NĖp�0�On�@�1�p�쾨7n6��[h����xm����
]��݈^�uv����s��mtz����3/�����Vڑ�O�~�?>A��"��ͮ�3��W�T��Q��
܉P�$&P&�4p�V��_>�G�\u�X�OK������#<H��j ӗ���3�w�q��ŧuZ�>6��2Kl��){��(���Dg�^g^pA�N8	�ʠI'sk�Q��ٙW�� &�!c��~��n/y"F��H�I=�]B�8�����;|��h����J�"IH�-�i�I�w�T�$�ʹ�fL�(`;�nz½�ۭ�$
�^_R���~��י�`��wW��4۵��@��떉V�g�v�]�|v�[<�h�m���7y
��A�}��� �y��|*����{ ������&Ҡ ����(��2d��C�q'L�O�5��p�n�`�B٤�/nJkOT.[ط���Vb�.�w�g�jb��m+����h2���"鄖��J�ob�Z�~�nh^���k��:*�d�03I�ןxz^����|H�W�@�F,��� �Ɍ�:D)�8K����6`��!mv
�8v�Y$Sq�OK�Ȟ�i���(N,����L��<��>}�������R��x{��(�	�����=��-g��);X�L7� /䮨�M��8 �B;��d�{�^5��|ǲj���*��*����o^����#�
&$�M�K�3��1�8�ݺb�mI����[[����Կ���n�0jl�x�����O���׹#���Q�X%���,on�*�'{@P�7"H��UR*!K|���;[7��p[��o��>:v�$�w�r��V�8�WZN��Q5�d6�-��qy` />�K�*�r^^4�g����l�q^!�C��k�+K�[ڵ|vѵ���G��&�k����-]����Rh�pv�ů1������� �_UĂI��]�Q!�I�
P�p�M���o�E�<���-�e��$���w�@�{6xK��:���);ƍ����L��<��/2��I����E�7����� �/*R����1Y�os���9-X뎶��&pi���d-i�iۄ�3��=Gpf�������\��c=�����,�O���M	7�]C*�rv��[U$���*�!gd�R0jl�d�򪏈u6!�ĠeG�����gĂ)��R�Oܼ�
	x���H�����!��Â!�]U[TH$���D�aq�LZ��Vc;'S�O�޽������z���UURM|T�6=��w��=�Z� "}�4�D�j_�K`�^:Y��M�,�i�m�6�-�.g���4k�.\��m{i���u�s<�ZÑQ�b:O<�[:�1���l�U$�
l�"t<QӔ��de5j���H�� {{v�Xz[�Ԡ$�REHo����t�����p�-~\�oFc���]��|:y��!�F^z�^?\Lm�t����MI'�D��������<�Z�q�����1���O����?�ڭ�?Kg�wnۋ� ���tς K�t����p���:��ݐ ����2v�l%Q�1��۪������ӳ�5��_��`7�|���V �f˞����HI�@�t3	�����q^��3���/<�UA��yUF�/_��� ���� fM����$ML)��D)M�s�ۜ����������N 2o�v�ߊu��O�\�Y��/z��P�j"*����mǭ� _v�=(����~@T�丆�K�o�$J�wnŬ�p�T�]Ř�����uR��#�4�f?�*�a|p�|2��@d�h��<�ܲ�Uz��0�X�=��~��i�e�|��z�Q��bt޾8R�ٽ�WzV)�ҋ|��9.�ه�s��.e�f�+��b�*�m_N��g\�W����4�	�̼{ܙ|���ຍ̡���z��$k���O��e2_d����N��ln*��3�oM��8�.�\�oj͒M@k�����kPr�S�3��pc�������:5�0O�f�!��-�ɀ=WٽP���ս��9�7�oA��k�����:��ESMwVN�F�ȵ;���|q+q�rd���b���Y�V�lw�H1��{m�mA�&ۉć���"���ɏ.��癁���n�h<y���KUB^����j����Xб�"�^�We�y�����h=���S�{̴���+ �ջ���y=�B|Ч�>�r�_���K����j5=���2�>�Pn�z��k跨L��4R�Vf:�NBĄ��1j����L��"F�98�MaG{���������'2j��+�+�G��=�N�[x�c7{;o�o)w�nq��վyoTð�!q�j��ѭ���R������h�s�f{�j*W�w��l��y�+3ɭˊ��K�z�2��C+�Rs���l�Z�wwF�8�o����@l0��&kM�3b�"�����= �Lp�MA�'޹����ذG�gR��9\ÍG��ʫ��C�5Kd�Y'k=vv�T0Ι���b�QU��**+)ENڌTe�UAH���.ڢ(&-AQTAX�V8��l���b�E�EAAQX��8J�QX�*�X*��("ᶅAE�h�D�E-ÅqeQHᢌEQUF"�D�,�+X *�U1h�K"�*
��������EYEUb(Ԩ�$P`��QEADDJ�"�"��±b�����D-�+E�����"���"[F"���"�p�,U��Qc��J�c�P��)��"(��b��(���#+m �E�*DEU�"���ł���TeDEb�U���5(�TEE(�
���AV)�Uf,���og>Bzc&��x�rb��.�w\�d��!�$�9מ`^�k��1ѷq��Pۮ��br[�b���%�.��Rv��ۖ��x�˨��j�\��q<�;��kO�s��9�mǊ��<$b�ԍĜ�ݣ��)���
D���b+�M����Z�aE�['Gn:�p�v3��s�����m�i��1���l���o=X{m|�u�l���;�c��;�Dh-;���ڲv��0v���p{є�&�u�L��a8q�9�pp�9ө� ��������#�5��̗[;����U�W�ō���.J��]�T�uil�;b�ɻM��8Թ�����Nɱ#˫�ˆ�u�l�8��v�\XW'�n=y��͞�yܵ������j6�v݌�t�m��Wdq�p9�ۭk��E��9����C X��ۮ�c�F���lY���]]n�c�
�N]	-����wF�vK,t{/g4�@��
a��m��{sݏ\5ʗ��7|���c/q���c2� ��۝�B����r(�u��u�j��6�Q����g���i�ێ������l���+������2����gRCs����gr�8=�G�=�>���^�\�J;�:9���qȁ���=��u���s�v��i��Q�kq�a���ۆ�#�ku��W9�e87��L���浘D�o[���-6T��ۋ/4pk�sۣ�2�h�a��b��>+��x��.^wv�ѥۗ�x<���WS�Îݜ�VM[��b��=���sng&.MΗ{m�r�;n����]g1�l��p�ͷm���p���� ��v��ls�%ظ[.:��<ۻl-�9rv�s�<3M��sx�mÐ�:o
��s��n��:`�i޷/.��F��;OW[L�b��Ŷ��Y�1��OQ�v�1��Yl���A���n�\�C�MCֺ�n1�e��8��Ke=%�ᛃ\�b��[���!F�^{7�����j{djG3���j��q����M5��M\��_���~n�͘�e��c�øv�v���<�Kuݏ;uu�u`ړ�n݂a��qr�mjݝ�k��V��ѸKv6읰;��ml\W9��[�F�gm�e�����J�#9�uz��k��i�M���N��v3�y�cN
�:���+<��ֺ����<��u����ult͸��i��Ԏ��<xݳ<�V��Ƀa�f����x�N���ݸۮ��^n\���������-Bg�S�ת=(�b kBnݸml�ָ-?����@IJ��*���	;q�Df��j���v����n^n{�s\��±�|�q^LRH�P�d��0#��/�����*�t��37=�e��|�A�^zX�K˻wn�h��L^���n;�霪�H�euMR	�
���V�na����X �K��~��h }�7�Z�]ۛtcz1����p˂L��\�쵶bߣS��tm�� �����,�����z�s�p��O.5`咉��
jaQ
W��Xޫoc�����7����6�1 ^�mݐ �����xd�0EF3�KI�Ã0��[<^��݁���1�����[y,�9z/���B��
�&�&_ǭ�| _vk�`'{%���GO{<^:��/�W�=���� ��ٶ�ҙn2���%EU)m|ocT�Z,���a�W{j.����)8�9ֵd�.k�����Bř�&
�,��|8�2r��p�o�<5��v\ɱ��fZN��S^�(����?�K��1�U  }���ۻ@ d��&��]H�=���wG �r�\j�"T�M'1]��R���qݍS ��\�ђ��ƤJonmشRG��G95(&�("S��5��;=����� ]뿕� ���� ^M㕼��s{f-�#/{�aY����MELD1��Θ�H7�5E��Tum�EnI�u�m݄�	 �;� Hɼrü]�D��^F�A$�eGq]���u�	�9qQ���N5�kF����'MT�{��SS
jaQ
Vq���Հ0�־� ��9aX�;=����e�mm�ڲ:w�Za�ds�T҅E_hv��XMB)��3��p`푯'J�A��v�` >���, m�8����n�N�P��0R��0lD����@g6�$�)1�{�mbZ�G��|F�[���"��B�Zq�䋊���Ó7/FxO0�r:�"��Hڻ�B�E2V�H�@Ά����x ~���	��>�b�"��W�G��\[d��(b��S��u���\�y��DP����|W�x�> ����#bX����1GBIdwlI�
�Dq4 �P�Jr�Zm�A�;w5��m��m��a�O�o}TI$�[��&������tT"Ft���g��i0H��kn�+�{t�8v�uָ�eg�x��qn�hz�a�j^��"*�SQSr+��1�t.j��Mt���9{hut��#�ܣ��r�zo����T��E51P
Sk��ݫ���t�?E�nMq;��@ >Λ�- ����ۿ��/4��q}nm3����SJUB&|�5�\�����X	)~���Lh���6�@.�s��ͻ��g��(�JU�����I��Y��M�~�� �/��of�� d�lϠ��Axx�(��E�	����(P�a!n���}Q{���3ΝO���>��^�Y��wZ�IE��sMM�)��)
��<��S*�b�Xz��$������g��u݇�|���j�ܜ��}�_u��{:ܿ��^�m���0�ؒ!�j���M��Re8)�ƙ(�5fv� ^B�pz��)���kr�<v���?�˃gfhAT�����Lr ���v�;�."���3���f�\�Df�kqj��i)T*��H�0��:&�i�%�(�.�[6I%���ݐ�e��� �\�'����<��cT*���@)^�u=�� a��*`r�l�라�@ �ͻ�"d�l��/c\�U4�QET"e�X��NU����"k�.�ߒ%���T�+�ɼs�z�z<)�fѨ��E��]�)�d])���E(��-����3�f��M�'���P��7{��vA#��e�� W�x�Sؕ't3���2�.�m�(j4�)�u/��'�\�ozث^��!�r���v���D�գ��· PLv�<�N���������nլ)���sc��ۍv�]F��ϙ�l�����V���z����vR����z��۴d�۷'�5��Iq����܋Q���-{c���j��;;���ʹm�Av���q���r��mnɇ;�:ݳ;�M�v�bݻ��CX��Cr���Oc���8:%��3
���p����QۏaF���{yƞ��ûx��e�����-���Av��c��Ҽ��qWQ�y��w���o�8.�Kl�&>
{s����\��U��h�帬��{��w��G9�,���A�dɩAT���´�mP|Oo�2����η�o~�At�l��o��St���)��v�������iLE����0��S�^y� v��Ys��[�����D0�/=-��ځUP���
W��S۷����yX�z��L@|��x��	��a�{�{��vW�sy��k��:T�EP����z��f�Vge�L��-�M[�� ,ɼr�����c:b��n�yws�_Ŀ��x��L�����e��K���>��g[ZP�I�Q[Q��:������U.��R���I�Θ��qy� �ٷv��o�3��GM]�d3�KLh�1T�S�4��������7�w���l����$�Ȫ���T���^YP��h
��<�7(<�|�����Óݴ�K+ ޱ�1�M�7�ܣ���}��˟~����H�;n���J��1�gn"��`�P���' H�啦�j��;wu�� $��9�{�єW�&�w�����@#w�nՂS�[H�b(S4���q\�7���� O�P$ 3wn���>%�����4ĢO��r�D�A�a#35T(�5�y`���O�zoe��ul���r� ٻwdD���i�7�F�ۖ�i�H�d(	�s/=���/nz��qr�[��G�q�)�?;���TQU��G1�j���;]�""�����<u���ݸI$�E�w6��실L�J��&�S�}���^u|<����_~�@�ݝ���|�����H��[
��{;����A1���ixg�{m�E�vs��?�7��g�3u�~��u�s o�$`ݡ(��>��6���֠Z3˘�v�]k� q��.�ww���jZ'+crt���ׯ=Qj�ಸ�q�� �t�m�@2w:[HMd�R��B�%9i�����JfVi ��6I q���@ټs�y���73�r�+����
έ�A1)�TAh8�s�;�LT��`��\���)���� ��� [�x堁[p�yS�����"�=��Z�m�[���/V���mRq���<m����"0D8���[hCm����݀����� �t���y�zflW�Wj&����� FN��L��t"�
�*�-�s�@�~��V��=S}�ی gd�� 3&�x��s���=���a��+�&f�**"j����1I�\Մ ]�<�^=ћi�Hl�l��n����kE����)O��cG�s����8?j̘S�A㽭*bA�^zX	 nfu��,]pC�H�tӓ���7��q��l3��h�Z4Mۡ.��x��D(W5�g�n��}�+2�Ն�̘zz;�����ԡ5ӅJ
�
��'�~��Aۙ��dZ~�ڸ^��@}�����x��	��v���u�����L��Ȑ[���z��]X�I��Ł�-��y競�ai�k����6
e�o/���e"�G��|\�����Έ��λ�
;f�6��=�-2 �/=-.;�D�U*j�P)N:k[ĬE��m��^�fe3� W�x� �g]� ���V�o��Ϊ��Z��9Њ�*(��L�k�@���w`���Ǯ����z��h�B���I��Ͳv���.�0`�/2�"l��� .��s� 2�ՄI�s3n�� H����E���z5x�zXdsE���TR>&��{w:�ȃ��ڊ�'A&"F��x.�m^�W�%���v@�Fmw�yGxYܷ��e?M��ٍ�j�㷺M�]=bP��;�u�ß٫��<HOG}g.C���|�VBכ8"27����7=�3^��'���g7l����k�.��p�Yv�-ѺyV�f�4�6�;���#;d{cF{sp������;�����ݻvI.��p\�"{J$��v��⃱��ú�/۝����x�{7=;�-���Ns�gn�]���r�n�x�(�m�n��w��g���N�t�u�3��}��+Y-�^�����z݉Wplp�dN͸Ů=�H�NuHۏ��]�� !�Ϯ9���vv.�\�,�]��p�9�Ƕmcg�8z1p�I�1��� ����>]uB� ���X|6��¶���T�
�玳�Ej� >�ɲk;�p�6%*�!�:��԰%�tʿMzb��\��^���	 fg]�� ��� ��tMx��~��c���k���Ù(�� R�'^ݸ�6{�D4�d�Y���P⫢��)f�m߭W�k�S���B*����2��z��c��3z��{�{����@�]�i�����˙�D�)�[}�0��������M���ƥ�iy�F�c!���o���"6��� @}���.ɜ����A�b"�1�-��ٍ�=\��:,�!o/6�X�۬����q�O��߸�1������:�X|��<�@n����ݫ�=���Z��E�oWq�rD]�٩�*�(��墴�l4��G_1s;ܰ�P���,`S.Lq�h���p�����n�F�MV��Z:�63���x�rv����8��c�5�o3Vd�ǹ�ّZ=���F�ȃ�ޞ���>ݛ�- �{/b߽.�6"b�.��Ă�\DeR\�z�, �/<�� ;}�7r��7u~��@�]�L� ��9 ���3�R�j��Jl�{w���p����(&��� �&�� �3�(��=�J���9 ��z*�3�"�
�)Tz;N��&�4OI<�(w�->��T�O�k8l >ޛ�1 _fu��2�d��������.z2�un�����\�����[�Y�2���:��v-??����2�lԫ�Ӹ�� ��/<Ҡ�_fu�Ff7���4�.�Dpf������(���>&�5�uڰ�S5��.o��q�祀�_��w�� ����uUslB',FÂS`��
���(�;3]�"���{�Y�MG��O��&d���f9p������C���{����G1MqU��Z��`�k*1���&67�V@�{Ϭ�y�.<(P�.�����˶���V �x�Al��M��ݛ�ڔ���K�-3�E��&iT�Ѷ��'v��]т]��%�9������������¥����/��S*�w}-�ۄ�U}��Z�6Y�X#"��= c�`�*�X�-C�X��ÁG\��VK��ڂ}�m�.lȃ������//.�c��x9����&3P��}�+�jx��>�W+=���s����'�	WXw)�5MG45��p����B�)�������o��(������\j!?Lg._.���	ٯ����[Z��CvX��B����[6Sޠ9�<̶�ڑX���Jm�+�-��$������vt
��{��������+9|�(+�#t{:��鋨�T�M���{Z�Y�Lݽ���*��%g39�2�U�?`Y:�FI�"�X;�;�y����$[3�M�]�gm���_U�����eK�L���]���Մa��Opn��ԝN�=���-�	�	�3)�W�p;<퉆 $�'���	V����4^�G�Q��U����5�f�}�9�l�L���9®�yw}�x����φ�w�L1�3�(�P�'whV�#**�Yt/��:p�y0�����1������._Fc�n�|[锃T��i��Y��& ��ǜ��T����7G|�+{��������89����<�%����E����yu��4�t4ƻ���,EAT�"���1v�*�mR�X�Ub0m���Ub�,V���+E`�������PUTF*�U1J1D���F1b�("��* ���E"�
�(��EQH�E(a���,V�#�X��
(9�����
��e"�X�*��r�7(�nqb��H��Pb�)D�QX� ��Z�X�qeJ��#,X�Qbɔ2�2�Eb�Ub�PPU��RbՈ��"��%DD�m��� �b �Y"�PQEETQPkPe�B""�̥U�D��X(���b�����Qj����,bF���UAH�l���H�#ETP��{�@5޷���_��l�����N �Q�^	rsМ=�<�x�i$Ԫ��- �Wٛw` ���=�CSRq����$�+�p��*5��4؀)M��n���A��:t\uLZn;�կs �.}�b�g]��#'{���e��-f�d�\VI��U"*�J����^������8�hˋ�]���Hte迿�����SJR�&_ǭ� ����v |Y;�-�F�J��j��{�5�C@|��ݻ����"fj�U5J�A&�O�gwni-��7�gz� y��� �� H<�,��5��q3��iW�
pW�1*�����ߒ'�wP�!j��z��Nc�5�}��8�ۛwh��Y�B�F78a���b���47�Ҽ��DU�c�a��N�K` �&���8���oˣf^�@F��hd)��k7q#r�o�BU,a(�iL�{N��K8Q~+o�C[˷y� F��۞�y���vDhI��:�X)�� ���b����q^�L�y樹�����<�bVw7i �F�wK�� 3&���.�ݵK�����(�Q�s^�2�����P�meG�Eh�ثv�@r�O��������W<sߟ����}dA�a�Θ�@fM㘋��^���y#�=�V@�����l>��9ЪiB����F��j��1��e�/���� 4���@ d�9` ����R��������v�2m���= �u�1 �皠�b��T�uTEt���0��IlwtI5䐼�ʂkܧJ�B0ULI��ݷ�JjFuߣ�x_�� �f�� ��ͻ���W����$l�H�����e�ꩂ���U&3|m��v���S�t��<}y5�Iz� ��qZ���!�ӓ���٩E߲��{j�i7Z��a����'�;�rn�=	�־<0���MT���<�iZs��ߞ��b����0��˴N<V��	�!>ٻv=�d�G<�Ir�:����ݶY�;p7��VRݵnv�u���n:�3
�ޭ�;���9q'/��y�V��o=[۲�v� ��xݪŌy��^����kv�j��C�k����r���Xv�x���f� ��d:-c���ݷQ�VT�:�G\h�caݕ���Kх�B�nX�v; 'L�*��pz�n�5IV�Ǟ��>|��o�^z7Ou�n���m�6��u��hl{ �=i�l�� =�sg��b
��S0F���Ϙ	iy� "OϽ9�Dɛ�hcj��Ei~$���,/}!9PL�*��Jm�{w��
��6��F�mݔ� ��- }۷jȈ랏z���呭�ɿ�}�ds��iB�J����=o����wa���u70�z:��}7� d�9` ���v�O�eLL�UJ���T�	7��^��w���7g�  >��ۻ ���nn)Y��h:5���$���M/�ݶ��A�w4��z�n�t?|����A�������l**�s�Ҽ�\�'���uK���
p���'u.��Sh����Q4�)Q�pj:�`��(UKH�-�� H3�u݀�����K�E��ߥu�ۗ� |wv�݄�T�2����AF�<��H%�z��ʨ�u����B�k�Ta��8�1�&2����;OT+.��nX�ܹIsuu0�op�M����E�Ю��^z,�y�jm�g{�@�{wn�"-;�-4RP��v]h}}a�d��Y&lʪT�)�y���ȃ��{�� L�^�{�j�����h ���w�����;�y�yB���,$}�rW�&y�2;0�g��"v[�`�.���=�iufѴ�����N�צLL�UJ���T���S> 3K�:*���|��Z���wv��#N�D?�[���$�o��V��R&"�H4�-\v^0�����������ֳ�wn��9�W����契*�!K�o�q��>;��> �7�Xv��\޿�[��nҲ ��C��-U1S4�B�Lei��5��ٻ�����^+"�wK�hKqZ��=�������}Z
��@λ`���L�9 ���A�^y�"@Q��0z���Q��߆�]9��_f;��&KǏ�RJ��f�J�U:L4�P���NL�����՗uJZ.�Y���Q�ݾɵ�^ɕ�x^H��� �7K�K�[�	ɂf��T�)������UU���ޝ~� ���t�9h�;3��O�����n�zb�y8�ȪK�8v�5
�-�[VĚ%��N�S��ܢL��f��#�3�ҳb}���sF�?�]h����Z��웡�\�������^�n�����[Q�u?>���8j��k���A'v:g�qy�ٙ�v)����� ���O�<�ث"&�D�cG�s�Ղ���ޟV\�V��|�@|d�9h ٙ�Y!��X���okZ��H��~��e��Ɉ�T���m��nf�:���RD{��/@��&��Hٙ�X*��ؒd
%R��Ê�xU[0�����P �]ٛwh����u��մy׳c�8vT_����[�����K�bÄ���K:o+�u��^�����V��zKP�Q�w���2��aӻ���&��vy$1��E�m@uHL�J��y�����F����>��@
�k��@��t�?qolU+��e-�	e�� 7�|C \\9�s����:^��m��rg]:��xϔ̿�����TUD)&�B��������_fs� �N��a�y���{jI���ٝv�=4�T�5UR�"j�6oe �%2v{a�5��}��]M��%�λ� ;�-2�}�mT�n�/���g�cW0����!I���uڲ ;��Dws��]�����v��|����LS�kJ�U3S
�x��w<C+��*�Y=���$�=�D�	��>` �g�e���˕Ӷ �w>�;=����(�SdG]�b$���I��&�mfӦ,׌}Ͷ�~IydolU"�K۹�D�zD�̓�W��S=���<���rϧ�����׮,�����d�H�R���{�p�_p�^�9Ξ	^��]�F��e��������xH� ��.{c�tg����T����c��q�d�vc͗��N[�6E�]vi���tϜ�G�v{;%����%0�ݔX�z���{�c�zӱ�;�b����0��[�Θ�m'8-1��k;��Wb�v����kPz�p��z���wb����ȇg���\�#���N3�ۑ�۴�k��-��[��x�զG1����oΟ;x�W..��a�S�el�P�h	x��)�0��15�x&�I��<8��������ok���A��^����G�Z�ɷ����ڲ �;�_����EUQT�T��o�k��Y�u���/�1���l�l����i vu�u��˽�a��O�`���UU*l$�N ���  Y���F�v�V7�� v�h�" �w3���B�D��Lg�s�{!�fy�` ��������ٙ�˳���ܜ�BIcwj������,D7	DU&4W=�� Aۙ��"r�l�n����v�� Y�X�� #s3��2��]���x=��! ��i66���n7[a",g38�Kv�����k�Ֆ$�}�����`"�U2!i�u>���>ܜ�R �g]�G�{�ys�{]�L�ٕ�h�^2��&��T�)�u=�q$�O-���>qdg:���uY��W�=X�!���ie֖a�_U�֝�B�^k�Je����!ҮTY�x3Z�t�fW:
����Re(zb~�J=e�����}���`$nfu�VA�D��.�6��b����C�%�<��)���v��ǽ�������� vec� �λ�G�=��j�����S������Kɛ[�3|�� ��|Ԁy���@��TW�#�u�ޟP�)	 ��R&�욋!H�j"�I��λ�� ��{	Tg6��<�u����^Ҥ�	%���vA�F���u�[<�8��G["@r��}���b������]��9zL��3���%�U5��f��T��Ј�Xr+��H�m�k�"�[��6�2:���%�5��U�	 c�o�{�D��f)R��9N��w��YR�I���ۻ@i��� H���r��c@?o�%UHMAT�
Sg?mݫ"m� �۪�rS��\���ºg�n:w�U	���m�����=u�^��;.�n;��ڎ�As3ٝ�&r�N�Vc&݌=1R+ȃ3:�f���]�uݑm���z�9Ȧ��	�QQ#h�l���w���	�n���l�����ܬc^��VS��:��ݐ�>��j�����W��'>t�ܜ�Rf8�X�z��'�1� lu�I4�wR���=���f�h��]\��֏=�������v�#��v��{�)ELԔooh
ET"�i���uڰHu���w+������dd\yv��ݢ�<��$�^��)�pj��4��:�h6qԯ^Up�y�q`d�t�@n�c� ȿLD�xۺ���Ղ��ڤL@�����ƃ��S;rs�H| j܅%_������Z��{;��go�����h��i@p҆Sa� U.�۽���.�F"5?J 0�c���@fec #�s��:B�`ޡ2:�e\�祪�t&/���w���w�໐�ra͸��/ޗz.�8�H��6���B">�e�M=�ʚ�O����E�� ���0�lc�L�*�6��Ͷ�"�s��~B�lr�ݔ��9l vV2!�>:�:�X�O�b��AJj &�'HW/x�2��h���7�ŎZ�&s��FV����!5QTTIT����TπA���j@ :�:���~��շ�2_�Zd -ܬc@%���T"i1�͞o�I8�ӝ�0�*x��$�{�D0 F��]� A���+����\*��S(�%*�J��:�h��s]� [�Fxמ�^���Aޞ� wd��#os��Egl�L�
Q_Bc+n\���ʧ�;�g���� H.�5�����/U��;��z�z �c@���SSAUR�)^h��$�?*�N���:�<�>�&�1���λV@�6v�[+�Ş^�e�ۆ�K���+V��)��F���t���4������y��{����{��v�����9f���OP}H��z345V�Z���+}�+��Z3yu��f���6u""�����Q�rYͱō:�b��GJ��`�����8[GB�������t̼ȣ���䧻��"�`���Lzȝ�hn)���Ub�1��z��p�y�^3�O�S�!�3�BN.J�a�2#�D��R��S�
��^m\�S�⅚�5#jbP�4�[���@7t��N�ah�/cZN����w=6�zRA�z�xt����%iv?z�F�s�(oթ+����醕f{�����,��bb8wJ/�]��1��*��J��W��g� ��G���:����1�s�96�Td+M�^RX'uf �uwc�B�7H��C�1���^��a��W��8��Q����+Ӊ�
�5Ӯ��S��(�ޏ8d���Ý�I	N�]j+Ӓ]Y��6����$�e��	;���!ЋSxu�E�),�P�����7>֒��z������ �m�[Y[T�׵�;�P���y%0)җ���bbP����y��C|��J�z�d�f��(��j�������mmj���)^ �%���"��h!x�*��o���Ѹ9^����m6fխ�3���wc%�o����fgu�b����5 ԂM��r�3����c5a�}r�	1�c�&A�x�E1���'J�� �����8��E�MͰ1�+!s��;O.
Q35��P�t�r�;���/A]�܁�6ь������� ���Z��,`�kwh�jX����"��W+��TX�U��j���ni��-�1AUJʠƵAX�b�,.)P�����6Qb(�CX��*DjS�c"���*
�[Z�,�c�L0�%��J�[Q!F.-
�EX��h���a�m�f�6b�������Yb�VUTV1n,���2��)�cEE��\S	��J��TjRV(�Q����Zf��qJ1QH�U1kaKTUU�J3-Epe�*5�$Å�(ڍiP�R����T�[j�%�J̲�&T��ƴq��2��m��E��9���ژT��,�UQ�j��������sh�6��-���k��nv�Sѵ�c�����[z:�i3��8����׭jn��{r��9�886-�2��*6���-v�r'��C�!x�ZŹ:37Vs���x{7d�q�vz�������GG=�۳V��q^�g�Y�m�6��v��:ɺ����p���nųv���Í��R�tϩ�kr��|vꃛ(�<���<l�Z�庩L��93�ѓnȑv^�WU���<�v*x#'�م�.�;�':�H���0�����zc�q��woV�E\�e�=vܸ��͞�!��ᝳ��u�2eG\�q�.�PBA�7.ͦ���.�J&��7i��-c�&yy�;`�]��dL�f�;p[�4uiudݲuӸ�ș�6�q�C��q�[���5�����N�Me��":�di�&\�ls��d[��s�ns�q[������h]�{7����@͸�qdc��s�:v�2�p�k��� )��=Y�;j��z�[���4��䣯9��4nё�ێ�����j��	���;tk�nc�9y����ųl�t�����L۷� ˶{ݘᖷ9�n9��Kk�<pi�2���,y�-�ǹ��j�W��;������m�EcXvȼ�Ȝ(���v��v�t�;�6{!�؎��x�8r�6ǟ1�H.�:P�yŷn�OX���\c�����;4��=�mɆ��s�v�v+��xcq&ms�v�����+��A�)�m�v�;�ٍ�n7%m��j2-���[�F63]L;{q�s��J����.-dI���\��
̮��f����<;�K� �Zŉ޶tF�E�rZ�����[Z������W"��c[y�<s��Vw��qi���L�3�+(+�����wd�zKY �M&:�`��u���*v���1�k�v,y��lc������[8�ᷰW�;S�a뵲#ۨ���svC,s]��c�DUڸ����Ai�ȗ;O2����t�k����=��0T��ͦRخZ���8.�g�㬝��7MОQbN�j��m=N��s��l>��:ݠ.�sw(����ļgy�Ws�k[7m;��粛wj�67d�ݷ��z0�z���ö	݇l��<mek<�祸k(��v���u�'g��+�2�`qL�s�}s�QL\�ݷOdG�v}5��g��f;��]6]��	���h�O8ڃ�9�N|���m�I���v麱˺���}>ܺۻr볋mv\��^����J%�����]pPM���_��t�@��v��-�����-2�>�}<��Oy��{+�I!>��2h��	�USQ%R��v_9b�7��^�;��R�F �'��w ��_�|�}���V`���\%D��&��s�� A�7�X /SͥW�כ�`�5��D@�ھa�*��S(�51PICZ�\�u�������Ft� nV1b����{9ɦI��{n�i���
8��T��"��'�#&�%���	ݬoY/2i���D�mv��`}{u�h=���~�����~��B��0��g�A����r�B�t(�n5�GF�Gl����?�>��M��t�+9Z���l�9q ��|�L֜��t��Ͳ��v�VQ�Q�!�	�S��b� ���d�SnQ�X�׏r�U�).@N�u��S/ۃ��М�w$���OH�c�&Q}O�v%�Ou���s²�����~�Y��,�~�� �]��6�����y�vә�}�y]�>&�͐�UEQ%R��uO[�Fiy�@��&�����vTߵ�D?����Ѳ�K�o�o��*I��A4�ѯ��#�C�Ort�:}�K �f����E�c�~��:��dG�@��6���")MLTPƊ��t"3�|�g��N�RyiF�]���t�9�h__?D���^:��AT�R�n���n���on�5�n����͒LZ0=�?~���@(�*��	�rπ�7K�LD0��m��G�v�^�Cu|6D@�&����qS*��*�Q)���m���FA}O����,�����o��ͦ@�\�]y��^��ґEU"�F��ڠ 7/��D��/E93�V
*&v�:��d�b�C9=��F%j8�VQ�w-ݼ����5�ҧ~J������G�34���eњ_ t�9D^�y�����&�QQUJ���QP�C��Z� �(o�P  W�ʹ 3;j#<�
P�PK<�,�R�*I��A4�Ѯ��� >��k�7��G�5�F	 �%�/�����6@�2s���k�u!�X1|
)���A�һ]Z4U�s��w0�;���s5���.������iJjb���8�6� A�{���a���y�z��oM4VL����ܽm&*/�虈�*R��1�U��Smx����WIo�� ����@,�튤R@�b��6k��2�b���j"������"Sh���""0�֩� �x�V�׻md�9��3�[d��3�}Ӎjj`EU"�F��6�u�>�XmmvO |�+�� �/Q ��"�����E0�`�'Z|�l�wi���$�gu�ʉs�{m��s�7�b���V;�����ϦGdW7g#��w����$�l[�6��L��Ҫ*)UR�0��/� �&���X�ih`i'��D�~2w�}�@vNc��
��f$���ȑ	����Z�q�o�6�36-�&�q�zg#�����RML"	����o� n� d�9�Uu�ϮF}��d�d�
Wa"���A%����A�7��S��@�{�\C.��r� �}2C����ǩ��ʙ��EDJ��ƐiW���#���T ܸW9�t�� 2srZd�fzY;/�a �����r�f�����s�D�⧖"H��`/�4zz!OlPOE�b ٷ��M��	���UR(YJ���V >�ԋ�!�$.
���v��� �\�� ��K�vZ��Ip�Oٗֆ��s�d�����J�T;����'TW����jw��+�G�����*I��N���d��wu�˵�Z����o���'\g������%7;��,�8��f�nK$�xN���4sͲ��;�Ղ��9NL���ۄݣn^[�=���q��r��Lc{c�v�p��뮎���a1��l�g��p��lhz2�{gcs5�x��u�磹�v�nl���{�o�g�6=���&'n��=�4�8lu�3�Sv�&�Ƭo\<q�93�Hwdjw/�Zdu�\��Ȼ<|]0����77g̞;�9׫&��t:n����C�?�>���:�����:�� H/��5@ v�6³:�9��?{�g��C�Ζ�f���VR��J��!M&4{{`�Ni9�����N A�fzZ����@��]i�Q����n��pg��(�A�J��ب ��4���~�T���Ӛ��s�oc�?���&H�ED�_	�4���Sꘉy) �ߚ�@|���n!�>2r�f,�^X�=��y������"�jfb�����׵�m�T�=sS���C/\�r� |wn6�> ���i�s����~~�_]n�W��5ģ��|v���x�9�bm���wA��.��y�2���}��s�\Y3���� �����';%����ڼ���ۖ ��m���!�C��n�R޼�J�O���cX�#�r_l�Z�M�B�cM��l��O�d�L�\E+3ق�Y7��V�j���;�c���\���+f�K�W�T��n!�d�d�@��s3��Q��\��ޖ�}Sd(�4B �Lh��6�F�z�1 $\��=����:�#�����9}-0�{�bp���E�;��ﵚ��g��� �^	 .6�*��+�3*nh�;v�ﹿ�}%�d�(��
�L��Ҧ �g�TOw�5�U�d�|�;��4 �^��� ;'1���휛�<��ÂP%�5�Ѓ�A>=M�
ݖ�˱�ùI�v�v�y�q�;������zy��D��o���D��:b@$��,/Ί����wk���{�L� d��L���!cM�a߰���u����{�4Yv�ژ ��/e�>.�"��&�����s8�^nr'�̰��h�SR��u�T�>�3�*��u��ew�6c�q�S����шu7V�9I�s48��,̬7D�]������Ա�f�:�Y�u|��2���+���ͅ�u�=�� ʾ"#����'���Q*&h�A4��=��J��v
���&� ]ϭ�,��3=- 7{j��Y����a�.�쒢*b�*
(cEp��� A۹�~پ��;qx�K�c ��rЉ=��^�/;��k�4�J\�Q�Cm�7Dj�:8Vb�s3��z��uK���ggVX�=��""
�+�i�u9��,i��w���-e�ؽ4'*�l����ݨ�c�%���&� ������g�ۛ:����ne��. @}�9�XDoci� ���G.��a���3D�SUTD�gx�n� ����� �<�NW����c`|�Y��倀7{��O�$�	����2�����C��B��=��cE|fg�A+����̫�.�#֦u3�C�6�yO��L�ԕ��d*ߒZ��{�P�i��%9���Ӎx�w�8�΍�]��8��A~3yv�1�/Q��Υ��ʜ�sS��r��{�l��D��&�=ݍ�ȁ�޵/V��՚�����P��;.Ej� w�n���\���ccy�$���)���u��, �wM������6m<����|����ؕSJ���9���7w<�$Ԙ�P�.Ʃ����m�D� wv6�}$XvB��
��ȍ���h$P�yƖ�\�p������ܙ��I,�|��pN۪3�SN��q���EI@)^���z;�f��R� �dw����_�qZ\��� }�� �|6�^�T�����&[;��v�����g�E�tn��L Ay7�i$C�3*2C&clFF����5�;s�`�>ؓd�����2�������/y+ՙ4�ێ��rt���s.Y2�O��>�|6@���s�Ͼb;'9|��2��b��(b�Zx���eF�7��kM\�g��-i����q���~�y%q��5Z���L��>^�'��z0�;�Z�!�Jm��^��E�1�\q��\s��>|7��ظ���h���Q����s��Wk^��=s�=�\2t9ٹ�c���1e�B�n�jw �;�����q�n�lt���p��x��y�ډ��<�C^�6i�c�Ț�j��ool�e����}k�w$H8l�)��Z�Wq�"�rbs��<=�B��q����7v
`���멉�Z���^S���γr91�J��^��n����вG�����v���Wi����� �oO0 ��-�'���WQ��Ey��C@�|?�����i�
(���بm��qo=s��ɀD6�F�vNc� Llr�aܺ�r	�{���'��Ķ( 	����PmN�� v�tDW�+�3���I晴I�&?� �\��ܹ�x33*J�R������2g��0s�y�A�d�9` ���wU2e��3�� �}<�4���,��l���C����TI&N�&̜����ch�.�/vZIx�&	��
�{nũ��ErB�2a�����F��c�,��`��Ӷ��k�l���#:ó�-���Ѣ�~���.o�����@���@|��m ϟT��SN�g>dD�o��U�U�h�A5h�oeڰ_9�K�8��0�1���e���������H���hh���8�U���]�0��M�D `l�0��c-���J�����﹘d�*=��O�c�b ����@ ��ۿZ)%E)խ+.O��ؓ^;*�:�*��������j��7��݀@Y�t�{A�'~
����D��" $/���X%$hfB����La�nL���1N|g� �^���A ��w�n�$Iŷ���tnhU6p%Ӻ��U�3QUU��6��_]��{>uy�q�9��h>{������)$F��
[.�e���l�Ӳ��یW,�:��s�.�m�.�8�;e��iˆ��R�Q]�����SS4/���q��d�rl��4I�ϭ/��sd�c�h';.�ကF�vۋ��Q=33IMM�Og� �����=/zz;���I _wmݠ4���C@��=�c��4��
%L��1����� V��גIO���c��d螈9S�Ab%WZP���;��p����H0����o{:�'�{Io�����|������]�*��aͅA��Oh��$ur��6��S�a���re��.�# ��VN8+��
[r�4c��0�<�p���Д��d��yҜ↘BŰU���j;4�r�Jе���b�3��� ��Юn�$�[FnL�kdU���n#f�ʋ��=M��w��8yoG6�w/����l��zc��|�8�֫P��m��C!�{��E�:eLܝ[��e���3p�΢�{cV�{�6*�\j׹t��'�z2�O	=�w��V*|�;$[���ox�&�V�2x>�=�uG�F	B���%��t}{�N���0�����9��8��!���
띃 Mg�b�^��g��{�f�o�bbd�w�}�V	]�(��AR��7 ��������$LL9�t_i=��1����5d:{!�Z��N�ԩ�%Z�w��$��R�mĲY9M�=(��ǩs��y�[�G�xo����~+�+j�U�+O�4⑰��G��q��a�
7J:�/�}.]�/g5��N[����!���n��wPy�e��U3Zn]�;:e�CV��@AfƩY�(t��8bKN���vCV.TŘt�p�-8��ѼV��^<��*��L�M���m�a�
ik��dLD6�GБ`��O$#�,�<�y2PBƫ��d�N�U�����T��LE�pc���ZMS��|�j:
����\�l[DE�	
pMfz�2��A�>4�>8��,ͪ��W	X�֔�iPm*[bV�����J�%KmEamL7�j��kJ4��,֊a0`�V�qJ����AB��Z�մ��k`����
�����V�28�0���Ki��j	Z��c-��--��U��S.-F�m��
�b5q�����p�-Z-V�h�X)�L5%�.i\6�m-�UeKj���p�eVj���kU�+echUUT�PL4-�.���T�T�ڨ�.Y�(�e��(U�F�-�[W.,ba��m�ڈTeV����.��Kh���
�����QZ	YLcib�cV�Q�j�(�R�f�L3c v��=X�n��l+*��ZX�kEkm�lY�S4���V�Z��-^￳����v݁h��[{h䫎OŲ��*hcEk�mv���]�Q����� +7�݂ �z�[@|������GfJ ��eڰR�Y(�_BdG����Aٙ^�ۈ�U�P�b��ooD��MQ�ϭU" ��4*$v��[�QqR��H���E�D6@9�r�2\tr:�m��u��g7GF���m��?~�}?[U�"%\=��� :�� ��������C[�"_��� t�쿘��ASA�L�L����6�_���M؄�(��	0���I'�LЉ$�{����#��O^凧Z��i)��&U6s�L� �̯?�""��L��l�O/uI|��I��PEGb� �!�䡙TV�^����'^O�
�3� "�{l�-u{$ۜ�fyX��o��3�Lr*�̫w��˭�eo�w[���@ϊ��[�8�Ս��ئ�zQ7:��+����d�ZLD$��o����_���`���+�ӈ` ����>�{�F1���a����崂 ����D	۝wg���pA\u� ��6AAy���E��v�ݵtq�o�;Png���˂#�W󿟡���N���a��n5�0��� {��w�8�I�;�xj�dd�U"�[��q߫����"�D��7��v�8w����Ǆg�MD��5I$=��Ey&�tIwd��ruK��M4I1U4-�o��379����66em9�S�Nv�ݙ��{��bԮ�c��0m�䒺z���
�M��
��z"!��;s����A�{W���[�d���$��TѤ���; �"��&�����X 3ok�x�k�v�Ǵ���� ^�u��@��3o�R#��ʷ�"Z<�*Z^����x'�%�LVw:ؗ�v�Ol%��q>��ӷ�Qɸ����O�����ߟ/�۠�ja+v�b����>�u̷q��:����ΞK�k�����a&�+=������f�7���9�m����n�x�t�ļ��gc�;u�3M�gr.��&��ٍ ��}u�g��ݼ���TYy�W��ط/�n���:���x��8�i����O0>9�v��N3eL��s��� �U�
]���'v��n8��u����N�.mq��f4�=uh�7�ZEO:�\��!78���-�]���nէX�����)�D?�{����m�6�d��/���\^oPD�$��h]�B�,�_��I[��BLeh�l�b���mA���v�#'oe�@��&.a#=[�o75�Ob&�^�CiC �A�0���e��>A�^�`��=�0��Ktg��@#;��Ҳ�0��lc�|
L�����a@�#<I�� N������h ;n���	��[�#��I(�˻���`�REULS��}�L�ۜ��@YN�ԑ��޽���I$���دR$��d�	���o�����V�De��0*gn]�y��u���00��3=O�x�n;��a܅����ACG�C2�׷b�+�b�ؚ@$˶��Q5u1Hw�U�K�v��aײ�ǺnbT�%AU'����*�������:O��i��,R��n��}mśN���"�6���ʅE��N���Q�#q�#�������no/b3�=˶�ӷ�� v�y�@|�2�=q5���+)AŃ�Z/�J��n�:A%�/��y���~�Tlu��v� ӷ��s?z�ѸI���<i3���f��u�U�m�TG ��1 ���`"O��O:Q�9���O��z4۟1HS*�h&}��m�`| fnspo�r��3��$�k:[ �y� �^�u߭d�!\Vu�jQ�WG����%۞ݞ5�>np䝝�[;���ہ���Z9���	e���`(m�:���tJI�y���$��Hnh�_���t9q�I�$��󆀮�(�3D|P�K��oB�_
�ލS;}�� >���� "�s��Z@�3)2�!Ν�t���TT#�f fe�h�tĨ" ���j� �E�j�Y�s.&�P[���1���g5X��1tw{�Gs��T]Aｰ-��Rզς�%E���oD���yvk�7����;&.���]z "�s��_�Ie��E*�Q��7��GS�#4�	v7^`A���w����;ڳ���K;pI۬ro�*o�.!�C���K�ݗv>��7��rf��y� �/�9��@6^�14���}�~[�jg��3��^ROj.=��6�E�2��5�z�z٧��9�������u�/S�o�̯DDr��w��4{����N<[r��]4I��[۝wiOH3�m�&)����S>Aɳ��Ξ��{k� {��q�6^�@�#�ܫ��y��@V�J�J��>	�cD�����"=�L@ �N�tϻ5��� wvu�� �{��>���b"��EEPz_�n�8�]8pO�Tz�wf��� K��ۗ���댼��+L��]�@E��\bU!�װʫ��[�;��k,EpLt�y�11���=����.4+�o�WLO�#+^��a_db��@WИ�I���`;2����*�_���o]� /r[ ��r����r=��WT���G	[z^|m��؈D'�G��(s[��<�4�A��8�����' �����z{.����1@�r��={�v*ȯ,&;ט�F��GKܗ��TA1HUu�xM�͙��D��x��~��=�I���|�ۗ���o������e���v��ڐ�86��m���h8~���˯?� ���V��m�;߀����-�ۗ�]J�����i���+o&�ou��I$i�֩��v���@ �ι�,����&N��E�EI��[jQTY[�M� wvs�7�\Zگ{�s�I�%�I}&h zt�l�"�^�x�>^�ބ��_n7�E��Y8�\�E3s����1����ȸ�F��*4�}���f�n���
����-p�G6�*=uu�I2��%m�E�����M��;r��R��+<N��l���Ҷ���]�6��N)όh^m6�Y�Nn2�:�.���yYbU���۴[m�s�5�^C�۳��OZ��e�3�8:�h&�����k۲f瞋k��vs���	˶�p��[][�s�l�`�vmcn�8���ۏ7s���\�tJ K����x��6�Ί���S$8y��[6���!������˫ m��s&��l]��aU��R�I��F�	��i$Ofc�C@ ��]�A5=|�+'�^a�:i� �3<����Y�Q51T�L��W�t�]�^	j�N2F̞}Z�$��4*$�#�O$%7�I^i��y�Z�|�"��ET�7��{M� D^ns��%�r������>��� ���a�Sڦ��⪠%:���[sw޸ޏjͪ�@%5�䖀A�����F��qTx�<�&5 ����4���q
3D|P�:���d� ��l�LLE�$���PQ&����q��i�{3��/o���>Zp��kz�]F���i��֣/�� w6��� �nJb@�x+A�Kn �[K#��v:� 	�g;V  �����:��s�b��'�K�s��i?*:�Bp
~"��n�M$��Ξv4�fZ��N⸙�yU��V]��׈������s�)H&��۸�e��69���{��׳�Ga^୚0�dRp$:�{.{����wh�n�SL� �Uk�Oۏ��6��&��(D�})��ݖ��DGu��>�p��{Y�M�ۈ�H3���i�������4�����Σ�]�g��zM��@Y��������@.��8�ٍ�ʐ#��nҰ�`s������	)���z��������A׷�� dm�U"J��F�<��P���n8�P\ݑ�5���N�E�]�m��ո�]���&�ͷ筰f����H(D4|�3�����ڰx��ng�Dt�i��yն�U���6��o"��������AQT����q B��s_}�1k�8�d ���H�{��&��=蝫jި�|(�G,�
Ҩ�=�b���� Q>�:ζ��V���h5Z����D�7�x�eu���:ל�F{��`:a>TY�A�5�V�k�(��ݸ�F��fVW|�%�Ȉ;3<ဥ�mTM)�P���wM��̚�p��D���$��,�j� ^fW�����ۺ��ٛ�k����OnK`�}�!MTMUE6���l��v����j�ȴ���_O������H����� |-��;�_��u{�����)�ݼQj};����gr��IN\�m������b�*���A�<t�{��@$ݻ�wh(�.����≯O�4��8h�я�	B�)C4�V�eݢxE��Tk����M�*`������j�A��b��ɘ�Ң��W���"�םي��0TU��Y�M��	ov;J��>����t(�k�� Y��p�I%۽�~���)6�"QpL?J�����EL����� ��w^h" ��ۻ@ �̚�ar��Īn�^��>�*Rʼ�θ���aV�/U>�x1�)���7�a~@R� �48��ط�|���MB�&- �����ͥUPU S})������>�rb����$J���ۻE$���ȯR��;�A�~>�XH�� ���>�2b��b�m\�n���h���7���q�~����n9��j�(��F��8����{[�@ 6w2[H/C�rK�� gv��`���C�*>*�%6��zҦ�����k����ί0 wom݀���T��C�9C��f$�ݦ�[+
�)+���]]o��nc�����c{j�GT�3Wg�H����D�p�{�ni#������'P^�s����	wu�-�����f��5�o2[��Gu�4���a �����	;q�>ney�}��ۺV
�fI�I��� �y�I�H@����$��H@��H@�XB�� !$�$�I��$�	'� IO��$ I?��$ I?�H@��H@��	!I�B���$� IO��$ I?���$�hB���IO��$ I?�H@�p	!I���
�2���?��2�� ���9�>�7�`=�h [m�h(Ph�P J��hm��kS@4$ P�VhM��A���N� (^��$���T�@���UB�B���ZJJJ��*��H�JBJJm�H����V�(M��U���QP|                 �                � �   �     E���9��U망��Y��w���l. �)���
J���R.wS��ܝ]X�pP �R�8�r�\Ґ��ҥ�O�   p@�{i�,� ���Gu`��;:iJ�3s t�� � ˨�eC�8� y����IR�c^�   ��  �   (t = �����{� ��CAҳ���k��4��7C[^���{� ���C=�70ʅESl�E|  ��y���z=�=�x  ���=٪.�4��C�T{��@���@�w^Z /2�E"$T��  > �  
      N�{���p ���� x���4 y� {�:=���` z�� x�=ެ��@<8   ����0 �Y��H�$TU� ���0: >g�o0  ��@ v�c� D(�;  �70��</��k��wpʴ�ܵ�6s�ͬ�%HI%/� �   =  (  �ٴ���'uܶ¦�wY��weՕK��u�����m6��dZӝ�ks3�2[��v�]�\�V�iJ���ȡ  �����U�79΋a� �]j�c�ڧ;{��j�7@��gF�W ����wtR{�z*���Hbv5%J��k|    =       އZ��NA���j�;�ڱj���n j���m���ǶN[�l�9�6h�� -��7Lq[u��"-�5E/�  �]�}8��^wP�1� -ڡ��uRڷ!�b�s��*�3��V� κ�n���T[�ĉ��;�7EI���42��!� ���%)P  "~�U(mI( ��E4�@ 4 J~�*��E  4 H�F�)Rjz�`#�?������G�	�N�U�B��?��wU���I_ Y���I[B!#�I_Ȅ��%��$�	&$�BG7�w��*b��+�j��]B;��J�_�����P'���N���E1k,�*�����k~觘�;	lǹ/k����S׸n;߆VK6�H��K��x�U�(�*^�[&Tx��Tr��b�!�rT����.�t�(��CR�b��`��4��f�mⴀՄˀ���[nӹ���a�z���qQp��;w3�ʫH)���+j�+5���	�	就�	��m�}�������]�w��������n�3�m����ՋS3���3�n�6�:˹SYpM�8n�X�f���>ɷB�q�a�Io���x5�X��Jb.�� ���!���
H�"[xӚ�B���]�K!E[q�.�8�J���d��cV\W��g/A��Ը��b#m(6�^��)�DQ�f��)�Ǚ{OU3j���Tڊ��#;�ъ�Z�e�F)��n��
���J����3Lki�+�� ۬���I�����T6�e!U�p~[��Y��z�ۧ(�;�])i{N�#�c�vk]ǖV*,���SLvr�7a���3l���w`�+4M,�l���fLM�f�Xݱ�*�8�Iu�c6���ܔ)D��QJ�����,�Q�KUS�������7MPǫFe����t������N��:u���m���!�u�¶��ϡ�����5Gr8lh�����b�6�i�|�1�"�f̔��WW���l��m�Z��v1c��e��\W]n���C��o6��O[Лg>��S�ѽ�6���m;��a��2L|��&�ʸ�c�{u�mn�2��O�w`44*���b��t��=��w՜nr�����Ckuez�X�6�/%"���=�&�wTF�&
ϧ۔��8�5������rfQ��Yi{�SƮ���Ͳ�Y�L6��XL��ט�� ,�V��33F�5��ua`���P6�g�l)����4��ź��.�,�9Ϯâ����u��������p��)o��O�҅�m���6�*$2��YOϋ�M�;Gw�r�LƎ��vI5����`�2V$(���k
�z���pG�-�oU,�Vӫ��r��6��F�*6)��x��LS�D�݄��MnT�e�� U-��ݣ�vf%�kBl�-�^�!OV�٢U���F��� ��>j�-S�)�v���<�w&0�A/�2�,<2�L��'m�̣V�Yˍ9NJ*�	����'q��y����w�ѭ}�A1m-�Ɗ@�*�ϵ�I�WGkI���ں�Z�P_���tE&a2�Aw��ɓK���eݺ(%E�7J���*�,Ef��OsO��2�͉�.�Uk�V�����[#.LB��|�)�qoBS?���J�����/L�S^�P=ʰ�X��,P�e�.��`�f��ݧh����vlGD���	�I*�T��(a�;�*GZ����)Y���-ʻ��M�(�܎)g@���YN�ӓ2�z�HA6���r��\#|�q�Z��L�Q��t��̵�MOp�S�D��6��Z^�^Y��쵫�A��&H���RƔ0U��oѷ'�P��!�E if3��-��K\�*�]e�k�m�jەf����]<��m�������)4j�Z���6�H1Ak۱�m�fi%�C��eX(�=�u�2��*D�$�ƈ�-`O7t�b�ܸ�;P���@e�[��/)}��f<�S;�K0,�����hݛ�e�ˣt[t��G(X����[��~g#�ga�M�G��[��=�yE�iKx`L��i0f,z�d/�8 ��SNmj��M^+�� 6�ֻ��+F����Z%�͕� ����l��N]�k2�c����e,nbz.�3�i���ףT�[���X4,]&�F�8C������[�N�!t�'o����yklP1m�UԽ22�V�@�V��Y1i�`;�5[�3v�$�k1BP�IZ@��/m�z��-QVneLM]] yC7���Bj��X�QȻՈ*�f�B�R+��&�[W�N�b�j�-xff���]��v�6��F��
W't���o���`�7�so1��f&);��.�4E��'�|�U�y�YA�&��9;FZ�:ml{�%�Ö��.�Kɐ�l�e?��r�E�&��i���a����ڙW-�nc�����Nnݽ��R�N�M�ZEm��#ܢ�̀�ߦ���b6����,�vdG1��Ӹ�ܻ�mQr�ǚY�z��V�h���\��ݽ�R�V\X��z6�R��!7kl�H)���B�;�Ѳ�Kɸ���Nc�2E+kd�¹�W�j�Z3n�)�l��;Ym��Lwn[�/�3�F�&#HػJ�Ȳ��AL���4�+7�c�k���6\�V��51�uP�[�6�k1^��	���	f��%�Ĺ6\q
�웵p�&�Wse��S.�ʛ���.����>	��,��5ذ��r��Z+I;��
Z�9�?:�NVc�ww]-�1��#���(��w��;ݫmm7GC��7.лn�<���.���ڂ��ͭq\&!b򖳖�B����]}v�c��u=�[t���)Qt�X�U�J�[u��9��9Xv�S�Б"T�٦2�-S�e�"��Q(��n9ZB�t��%n��:�A'�.j&�C[(�Ғ���X�/+p͙füڥ�0"�ڍù��2�M�a�z�r:�f��iJ��:Z��Y���tŒ��U�V�'��A��ܧ(]E�m[w�S9���W� Q0D�zp������4���h=�����w �j�
���+6�4��ͽoW��ʼ3�Va�����v�խ�kCf���"HU�D�y �k.�;�Y�Y�\Rj"���i���CX${6fQ��˖5��ê��5Z`mM��ۚktb�t�#6ՍɃo4�C[ݡ�E�=����Q�1mr���nJ֥�s('R��c²����K�f�+Y��J0�H\��X˻��VT����L��J��x��h�f����c��!��L]kmP�ב�r��-\�[+j�����v0<TL԰;� ���&q�io�1�cSne��\�1&:����\YZ�?#�� n-:򣲔ئ˘��z���Ũ���l�%�ɣ�&�9S'�����A�L�S-��E�s�M�fn�2#�>tRn`��<	��s��u�6��c6�hVd����#�va�$����Ks �3#z+ �a�u0�����YK�>�@<��xiD�f*%6��U�H�wS�˗�T�L+�Ӗ۠/�I+�t�h/$f�r#�2�a�3Dr�Y�����pZÖ��j�&]N<�:un�&h6�b�K�Ȉ�7.�*�@:{k�O΅�4���{�nnY�g�f�^�Ŏ�c]b��v�VM����j���͈��]�+�9�����@ݚ�4�sU��m�D���[�b�+J%{Ra��WX07���H���hs�ŕl3m�
�-��Z�*��(�e���1CA�����l,�V��l-��0	�7v��l��Z�[������,ٲk[�L�wJ;p�t&nY�Cכ�D,����[���7xH�Efm�{��fR�P}/u�z1c�˭V���V^m�n�6�{��m
��Q�,��K��o(Њ����=y�ú ��ښ�)�n��2��S(զi^L6]ā�1���K1�5l�Ǧ��Yb�5�����e��xl���J�3֣�s3X%n��/2�K�9��hh]��	�vsj��w�/v��WY�^�	մt�r*D�g �̚Z�亸��o^L
��Vņ���g!��L:�י�.$�x���U/	��mŪf〽e�DV��-�������uZi�V�>�U���/�ZL�=f�㷬i쭻1x]��fԊĂ���z�+(�[rκY���{ôX�H���2�9i���ܣ��)[4Q���Q�Չ�#e�+	����FhZ]�Z�-˥��W�N�I�F4K��ܦ��C�2�3$������qaY�\�Y�B�W/T��c:Pϳm�h��Be�2��F��"ھݙ���A��Uq�Ѣo1.mِ�q��с#N`u�/B���t�U�b��ŗ�e�~�R��5�[��qh�z� �fI�v+���E��.f��-0�՜��c=3p@ݽ�E<.�<�k��L��F����c�r��W��\��c0ZU�7%������ku;B�wJ=��Ae(�n�nX���Ժ	8F�mm��N�un�fRC6��٥Ha#��Ve�L�x��P�Y����r�e�vFȣ�`��/��#!D��ťK��䠻�%;f�/tP���X��ָQ�H"]�Y�:�.�jƊZ��̩-��JJ�P�_۸��Yzt���ʼ�E4�:q�]fn����cq�&l�4��f���y�\w���r�6
E][��%-�Ɩ�&�j�ek@��.��Q�ͭ���rJ[)ۨ�`of�gi�:Y��7k�mXn�J�Xv� ����V��ɸи3A2��a��7��mZH���}��x�vr¥@ڧ���TB߱0M�j�
RI��O �33RC�2���J���W4�) m��r�9,a�vi�x�9ai��%f^�n��ۋQp��˴���ׅ;z�)g"ڙ���K:��w6ap�V� +6w(nT�ܳ�.r<�JDhǥW8��5�mJRf��f
��
�u��B��®��X���v�����^	�ZN�)(��m���&�Q�w%��f%{c%\�d�����W�h:D��N�o!�b�'J�cH��#JW7orK���8�=��RR�L�yJ=�c�~K������2�������{�Y�4*�9z��g��{&c���ݤ o5��pfe�[�n��U�Y��^�,�!C��2-u��t����q^`4�1NJ�a[�KZc7�Z��go��T0�M`9�S���!�#�m]0�1��#3i���vF34V��J�f����K��X�7�������^n`�r�Y��F5�K�\X���rI�˵C���P��^l�0��R��+m�ղY9�+�ͦ��2����ۏ%=����b�Bͥ����wDHmۋI�0��`�T�N���.5rm�s�,|UJ>=.)�rX��mn��Z V"n���%-��N�[ �G1A�����n�C�d'2��`t6#{P�;
�Rl�3l�N� G*�͓���6�.ma8džT��^ql4=���_��R�o���''"��ՠ���2�0�_T�jQM��Z�լ�k����f�퐫h�о��oK`��╹��m��	pЕ� ��/]e��۷�[�/��K�͊�oq^1��+d�c��p-�.fb�ܘ [C	�b|����^��jnڙx˨�2��@�c�|ӻw�ס��9U�X�'�ᆳ
Dl��\C��H5��8�\5���8�p����9>V���iړj�R�(�_B�j͔����r���r�W�iN5�uⶥ�V�G^틵LU��-���x�!M��S�;W-S��v2����tiܺ/�]��@��XKLm���Y����,���h�y��n����:�lb(�+tҒ��"�B�^�f�Y��,��J�2�{��\�7+3q�dΆ*̻�!�j�IN�e1GB �[�|ɶ��,ڲfŴiV��vBh��l��a]��ۻ�4�vb��Z�ʷ��s0%�)P��n��.� ��\�׆�l�
��-j�Y��Y��5�j�R�E a؆�p�w�����ʋ�G�Bf��"�`/^����];��Mջ��ܭ7)��E���dd=x	V�[�ha��K�^)V���w�t�x�� �5�ї��T��%��Zں�wE&f��+�e�ai_j�C�@;�j���N����;�L�4F�u�Z�h���ZDv�H��^�B�ݵŪ�V3z֧����u&B&�c�f̹�%��j��@U��+kUiW����X���N�vh�6�>/A[R�Li�nm�f��e�b��P�u��&���n={�L�d��ڷ��������IeViDBYص�!R���
�dջ�ؾ�g�Yw]��cq�8��ûh7��6���E`�c8��4�W��Ս֊GU����]d5���Ɲ�
��g�t��@Z���Ac��u��}��=�0�oB�Q�řCu[@��5�܂�n���`�F+�m+���i�b�'6�]��7����p��mMFh�̘UkH^�[F�� r�1R��-n��ĵ+D�:5}.��r�U�@\�m�n���v��/&�An��b�]^MJ�e���yiB&A�꩗eh�H��q�7iJݦ�h�Q̺֐���-�f���)�at���[���
:w� 
��%ܘ�	�82� ����v0�ek� ^�/sX@XW�f^b�%ѕx�[��u��`�h
j��X����X�.��ĵ�+N���To7N��m���ѲL����XI�t�M��ku�]-�Eu�U�hn������W�e�@�3v��G6୬u����&�Z�٘��d^]<8b{�b���լJ���w$ǀ���,W�)MT�K[ӭ���h�y!�]���m�uXl2۸�ͻ�<q���e�).\$��ZȜn\�upJ8���ʐ#� �ͥ�.ȱ�����DK�Z\k^�[M^�ʌꕖ��{Q�X����O2�3!\9&��܍`m,�� 2b�5X��/O۹h�7�-u.�Ú��fkX�h.Z5&K��s/Nl�J�V^G�[I5��!�ɻ�E�Y!����kp{|v�����+���7��۶A��Ǥ�[��h��$іPW�
t�1�%Jt���e�L��h��@H�@��I ����� n�*��.�㮲�묮�����:��ˮ�:�㮢�;��.���Ϊ�:�*���������;��+����;��;�躮:�*ꊎ���:�˺쫻�뺻.������.��.�;����:�ʺ�.룫�����������*��캮˫������.�������ˮ����(��讻����;���㺪*�;����벲�J���I B� m$ �쮻;��;�����*����.�諨ꮋ��+������������*���늮�:�.�˫�I! ���IZ������~����?��=�+�>��k��S��0��,K�Q�|��Ϯ�������ڔ�F'&��2���[���O�9LJZΚ3�u-U��X��[���A����m|��(sf���EvIW]�a����sT��X���s�f��wH��E3�-e����(�����]7w��
���n�t:
���&]:��$��BP�S�O�Gl�Y�U����Ab���;���ԭ���2�J;h��T�8.�ˏ8A+r��)_K����z���� �7�G�F�1�H�yYe�Z�ʹM��[D��V�A��\3�1s#�-�l�l��Ü��2��S���`?b��Y������u��V>Q��}t����s�W�ۻ��u�������[�lT(�����5u])��k�[a���s����c�2@�I �m��p}�h� � ��­��r�����v*<t���}[�a�=�e��sC��:�uW-�{}u���đ�3^m�w�t�>�~�_#��4cn�v�^���l��i����c��u�m��.�m�5��8�v�R�,�dΫ�}�Qa��8Ԕ���u�(��:���2N�ye�]���RQ����Da�����m�9�Z����sV)�۬]Rkc��t`*�u�J���m�i��s�21�lB+:�]+l���e�y�Zj��b�5�IY[�>r(���A��x�l�l�Ro��lqoD��ְ���J�����S�`�o3Sj^�sN�R(V���6T�IAR�r�޻Z֝ۂ����#:Zq�v�Ĳ��p]R�4h���f�P�I�&f�}uڷ�S%5aX̕�3��v�es\,U�A�zrSC-�M�7DU�ΏX��U[:��F"���T��^S&�c���Qf��!���#?)���v��k,Gk1:X�Vn�w2�O%��w6���
Np��AW].�r�2��y�7�soi�/*,ٓ�˾T�s�ȟ,�ԫٹ�7�^���X�G����51���7!�P����]�8�p((ܮ�[Z.]f[Y��N�a�0{�t�D���k4��+�������0�q����^��k����oV��²YM\e,�X�s'�Oz�Oњ�89�qW7k�ww�;��06p��XZ����;����h]�iT:�e�_%\�o��炁��Z!AC��{��)KyY�f);��<�Ѹm��\aW��@SwWg5tmA�L]w���ʜlD��E�G:�.f�\I����\����zĘg0X���1��* ��=���,<��*E�;-Ǐ�Xn��#VSo�����qӶ(�4�+즅փ�a6�V5�N��Y`�`��7'[ם:B;4�Ȥ��ܥY2e�է�أnCN�F��=��
#[��2��e�V=?5X�V���c�n��x�b,��v>͢xf3�GX:�^�f�����ZC&P�a�uݷ�
�2�c�oTa�,K8��/;�'�:���-�{,��e٠��������D;��Ep��p7�D%�����[O��]7rV	pb.֚7%��M,��nK�ϵl�v��@k�f��j����N���+xp�&2��;C�ƫ��+^q��bU�YҲJ��
[c����,B�g��̕Ϯ�uP�+fN:�F�fm��㭖�EJvDN��6h3�X�Q%ɷ��7.f�������[��i�c6�=]+��j��Uko8)uI�S�m��Qۊ����Zʼ��WE;�Œմ�k]�z�7/aᕋ.�M۠���%fN������^��.tz6�N�aCs��%���g��X�Z��Yi�Ll�3	��+��*�k�e��c�]�*"��wLLn�������ԥ��]�I�t0�ru�승�rsZ\hfݵv��e<W�Mo���k�t���]�ݹb��:�2.a��vc�j�}�2k|e��r��2���ԥmv�-��L�6*�p<�ݬ�sZ�(�l�^���Y`��d[��5c;k$sn�����zL�\}+*�;�騲�Y�gt�y�TU�v>Vb�ξ|�dYy����IK��/���2v=��=��b���n�ۛ���L�B�8�v��#<��6H�}G:�@�$Z��Wc�:Nw���t&+u�E�M�/6;�%���rޭӫ�Q!�WoU\!�ܛ�N���eeY�ӻΦ��1�F��ۖ�9V6�Þ�7�v�N/�������m 9w���#z	1Z����/&��Y��h�mX��S�Ct�IYg{Q���������X�I�OmWwe��9����@�e�N�]���;e��0�Iůػ�G+%MJ��Dq�(%�t�}��S2	�}հm3T��uf��{7e���Y[�#-+6��c���׮��v;P�c�ʱ�uA�2��e�oؔ��ʹG��-}Ҫ�+oV(-�m�[Y��0"�Z�*�udgK��\�%_rm<o�"�Z�69|���ߐ�yг��F�7qZ��2 �U��v�Pӫ[���t ;Yx�G��k��d�֘GA�a���4�otW[%�#+�ѭ��	�����ltg#�!��%Ey��v��6�����"Jj��絡�Y�Y���v�ҹ��\
�
lH2V�Z��[YL!��7��!�=%�<�>�#Ӗ�;i̫2uu9�%��E�řUhv���lZ�j�Q��PF�O"���ϋے�4��kC�v�����,�X �Ћܦ�F+
�K���R3r�-�*�|]v�gq�B}�U8�y2ՠ���6��	#�ǅ�!��3��������!J�H��X�"ꗮs�:�]��n��@�Ǵ!�7Z�KrAӉ��Jb������B�Ȧ�u���t���=V���R�B�=ڽ*�y�#P�9�U�dG8�ת;��+܃�����k24�А)`�#�H��'vM�v`u��e�1@�p�`�m웆�̻�^B������cLyXq$��򨥌���<ێcuPL��7�.�����q�ʊf�w��YUW����*�+*�J��L2eX��w�lTnI���-�xAw�.�\⮾M�c|E`�ņ����HA5G�{�"��e�ɝy`������#��X��MY/ZX��ε�cbяK����}�p�ۥe��C�h"ڊ��LU#�mlAkS9do�V*��Y])��w)�E��R�Z�C�d���Uǂ�(� ���AZ�.t�V`�Ψwz��}�n�[�+N�*aim�RX�� �[�R��f�ܗt7\mk3�c�>�F�RQ
�%h�.��=���N!K2`W���Ap���ۭ��mB<�]���e36����m�'�UAAN�� z�r��c0�i�o��w�VSFEluoL��i>gz�ʵ�3�q�sp�D�W�,�}�����C&���&'T6���m�w@�/sh��*�>����hJlk���4LZ�hv3����m�չ�f�b��@)�P���kn�؊rt�_(��{%X�ҝ`�e=�D�V���І��k�6�����!t�A��Jݫ������]d2��&��n'�3��P��gr����3rV�ͨE�:�vn��w�&:��A欼�SϝS�K������U���D�����.���<w�`r#�бǱ[`�"�z�����6
�p�ڋm}��L�L�v�����|���j�m�� ����٪��VATցn�m�w3��E$��OI�Y�.V���OK}��)P����ɕ֖̏Re�TAWY�]�	�/xss�=t�w�wh���&q������]JY�=Xӵu�����']��h���D��fu�z�8E{s���J�)d��ew[IȤ=�Tɧ����G+;iT��`���w�P2�Z{o��'9������f\��n�R�UDz1:�ͩ��W��K�+���3��(b�o"��[l�e��zg\��_tȣ�A�8�ul�]���<tU��%8;aR۾��F��!N�q�A�ޓb��e�pO��cv�ڼ�u��_W ���me[㐬Zr�\ǖ�=�U�EZ(.���K5�5A���f���z�n���z)�3���.Xn�'+{"��Ǳ� �M,9�c��u�w
F���Vk�8���lNE%��dV�7�n���J�{γ�n\l���]p��&�p$����7AZ;m#͞	�uK�U��/y-�r��+	H��-�7A�:�.��[]X��Q������F;�ͣ�S�%<����DV�M����r������yo2��ۘ[9���g�=��Y��\bL�B�JoU��-啮�\�=Q�o1�4�n_D�tUc]�X�*�f��T�ư�7�N������*�=��۬E-[Y�ՍO/,� Qg&a�����
���ӝ��Y�C��VQ1#)@��Rޕ)U$�!Y�'/]�k��p�8��Gt��p��y�]��w������\7�Kc:o4�F�����I|z!KM3�d�UX5��%,���2e�w�%�����+��aѩd�r�wz囝A�-ȵ8�՗V�՛����蒶^�!y�;D�(�&:]�)��y��&fi\ޥKx����4��S���-JMTN�:)��l^P��{ـ��a7�.��W#��5a����\��X]�b%��c�/U�#AwK82�X�r��_CڅE/�2��Ň�ʈt�Z�qz���k�Bm��[�ۦ���pi�ҁwLn��	)V��7%N�����l����7� #���a��*ܾ���(m�js/���3�VJ�z����C_V\��T��-
�;;�;��/n���ld����N�u��j�&�������Kxᾼ�eIN.��7-+v�*/�2�v>�͗�(��F|��ٺc�Ԅ..����e���F����/�c�ܳ�a;��������9Vf��m]��W"Yb$�E����̱[{���.����z�Y{Y6V�4[��tl�@q��*T�Ρ>�(j���V�1�ͬ�����l���J�<e����X��m��t�\b���Z�qyA�ނ�̹�i�=��f�6�C�ڻ]���R
�-uV�sa���'�aӋH�eCг9,��[6����è_��Vd<f�_;�8�mv�)'� P��fu�PL����BJ�1.����D:/8\+�A�s��xM��7K���2��j#�ވ	��]�s�I�EF�+�/P�RoQ���{N1n;�f��[�KUxw�I�W��W3[SU���$��%�	KXA���B�KҚn�*
p���������3zJ���9���ۯjJ&e�2��u[�q7bv5`�.���)�d��\��޾�{u;T+�;��ڜ.�j6s0��ӷNGM��m+ח\��K���R�����eq�rm��f�@tY̆�P̼K^�����8�증#JR��q[cD��+�t�K�
JhN`RԮ	�`�Մ	d��͆�����R�n�YA�.�������)���9i��u��)S2F�J0�v!{\G[a^qu�L�N��f�.Fkkݓ�a��d���E !�/9,��7� .�ad3�޻��D�R�Y����x����/��yL�5EnU��=:�SܩTԁ�Wf�����u��8P�w�{�VŢ�I� ����+B�h�J�۝û~�/X/&���h��녹�zzY��h5�h���g�J��G�^W��	�t+�39;یj�4U2�J��6T̷*��֪/�Zn���Ή.4�M�����/��M�\���+��c3�s��̓��e������kpN�,U���M�4�[�)�$E�y9�f�7*-{�,��HD���OW�wk&�R����i��B2���d`���T��+���X�`�
�+�mKh%Fwm���1t�րF��XUi�.��w��*�@dy����*�ge�M�t2���R��Vm�]"��[��ӵ٦�7Y��ت}"��l%Ğ�^u�qޚ�Kx��][�uo��ɫW��l�*���_0j��k���@�)�=V���v s�Z9υ�Cao�}�N�͖��D�O-Wv}I�wX�Y��7�٢�˾LhSnCMK�+I�*�ˆM��`C .�W�#O��ʳ�t�$�;d����a1[��2�+�ea}h�E��v��J��RY��FJ+��[�5�~����3X�c]�8��m�V<�޻+��s,�Mk�ң�vT�;�z�KUީd������{V�,���M�B	z�����p^���VK�-ee9f��xR�7T�ѣK(g�^Gv%u�0X��3ٕ���^-l7י�������[;`f��X~z/S!^6y�k�c.V�������hI�w�Œ���2뮐! Xo�";lL�j7-	��A�v�)Ab�%�º!e^�<�^��|��'xm�\�ɢ,�6��]�w!��S���tZ�Y/n��y�{���m��2+U�4K��AOp�[������vU��`DF��Ԓ��6��m���!hmHd},n�w)<`����"��
�wAwv�U�YZY��Uh�$����PK�ˤщ�͊퇕�b����ԗ,��ĕ"ÝB�6��� �����Ρ��BV%;�p�p\�ݳ)��ݫ7}ՖYҨb���ͱoon<e����㣜�����C ?E��&У�X�轗�10��<�7��]��F��dWq:֊��e$a6�Yp�t�N��(C}ld�T�֢�G��*P�]�Q_qiLr����X��Nc��H�5'�l�P+c(^U��4��1].�Fd�үt�f���6�r���tJ��(t�݄`���[�U�{0e���ӫ�����)x�&P㕖� �,Q{E����V��	�E5m��%���� P$�Va5v�[l��t�U��#W�LM2�$&�wK'+p��H�{���O���ٿ��Y�8�S#�>��IZ]�{���'���;ur�]2]硫�q竫�hW���80�#�p]*֩ͱ��Ϟ�M����;���Gv�eDB9Ʉ��H��,�[������.{�p���+�6����;&�f�ݗ^y�θ����j��m����v^�\�
 �.{p`;r��SKhp�Z;)�nz�,l[n����Ŷ��vV�PQ��n컛[Z ��N�;`xx�,f��ݮ.;sǔ׶\�y�΍W�qΥs��c�S��
'=A�\ad��1׬ĝ4���Ӻ�vi	��v��<����/t5��l�9�޼89��Y�i<r�\ټh�K/g�\4n[&��v8�C[�nzm�3�2rr��-�1ٸ�j�Yu
sd�CGԜ�v�!�=Y�q͔�u��ql�a�6�h��-�m�s#��Sik��m��ʚܛ`6�@��u�n@�]���κ�v�E�3�� =��q ����y)�s�9{S�qVy{d{�sn:��,��nZWۋ1R�bnZ��F�Ѩ�Ҍ�F���=���w	V�;�p����0�f�������ڷm�<\�x:�5Q�V�ٻ8@H��wh�WxzSV떽=�']/�ن�Y��r����3&�Ӻ��R7k�s�t�u�^y}C�D�u�5�=��ݱ�۹�����ɽn8S��3ǅ�ݸ�ls��3���qv�x�:�]�+�5nx��[v�3q϶v�j8�;�ra�K�cX�:ݣ�sڍn�s��;�{z��ԏ;]�����k���G�6ȕe��[i����Kxp�F�펥��t�K�:%OQ�s� -��g�s�s�Og�w�P�q�׎�''�1��x�y�N�N���6N�K]o(�a5�v�X��z���Vvy�[�v;'Its�یqa6�/���[�3ŏoIü�Mv�f�r�n��.#r�����fs̺�2�{,��EPD��E�\p9����ȵ�G�u{����;ݝ�n]l/��$�X�g����=�C�>/+l�u�u����*\���;s�^���O"*���qj��6��.�Ë�c���v����]k�Z�6L���9���j�c�����ksu��%���q���'K4n�<�x��XV��:OX��XӹO.��ǳ;�8��n6=��6�\�tų��NK��U����G����;�y،�ۗY�'O6<r6�(�Tc�l=\9NEQ�n|Hݮ��h�Z�zV��n�<b�.	t<�Ѻ:�ZJޙ������V܋q䶢󳈺�{�r�#��⓪!����7I��6ǰc'���s�bp-�=�N,8�c`���M���s�m��k��r�	Pυ�ĝ�3��\q���tV�1�u�����L�6w���v���Kv۽�u�ƻ9NCK嫛��y�[��nϷvɵ���z�Wv�kqۧ�\n�B��f廔M��rt&��^�F��g�6y)��� n#lٲn:ݻ;,շ:�]���mn���ku@����kq���v9�vF��u��m�����x���l�]U��-�n;���[=�9��y�I���ts=�]�u+���q��z�:V��F��n��F��;�vݻH�n�v��s���n5!�m�]oV����t<n���z�����Ț������=�T�VΉ�8�����v�x1㮶�v��6�gsx;pf����Ecs�q�ZL�^ݠ^����
�Q�N�N���lq���Gkn@��[��sVu�3	��p�<Z9��JuՇ���dOv˸�����P�"�s��\p�y�S��;��c�^x^1Ş,��=vx�_+���Kˠ/R�u�ڱ��-&���0�'[4㋌�m�ϔ{�<���'EG9�q��v�u�e�{:�3��S,�`�Y��n�!C���O��T�������5Wi�u�[�sC۷Oe�;vu����ݷv�P�-�6���䷃a�p��e�yZW�]���&���n���A�,���ݹ����u��Ag����]���\s����Gg�o`�[2{]�7<�����qg���n��٭��̘9vA#fX�@��rO�셵a��8���X�.P{lgB.��=�ӆ����<v�u�ak���=��	����,A�z��Ly��g��^�²�Ֆ�F�#���1����q����z�i���t��qn���؜v�=�ͤlvێ�ۆ�u�Z�%��Q�Y-�cN�6�cs��O�㳷���)�){1��]:-۷)�u��͕f쳈�yD�S�l/�EF�
P�\�Ms�>�G</c�n�r�i8_m�ަ�f���kYNI��rg�n��qۗ�\�lrh2�=q��jD�'V��H�1�;v��[�v5�Z�V|O��P��I(
5D��X�sͲd컫��Zv�hq�Q0=��8�cc,qj8���;Wj�m�̜'&�Ʒ-��8�ļkK��=���6;rs��E#/����8��F�y�3\�Al����_gr>5��a��Ӷ�'��H���a.v�y�����n�m�Yx�����vٍ�<g9;O�j,��;;��=k����==+���Q�qu�m��ü������9]{�i0�xG�ۦ:�ݹ�e���8��FofH����wk��p�r1p��G8ܮ�<7p�g�Φ�<� �����t�a���y6�f���8zS��S�ۧ����k���t���
��f�uZ���<{09��[q��q��ه'dGy��p�q��f��]tKی㜫��{^���&���'n�U�#�n�������c����nM�t�{����ԫ�iV+�[��"������ju�R=���.�0[�]�h�.y��ۧ�[�a:���suю������p�Cm��g[vǷS�O&%�,Bļ��E:#�@�n��������z�z�&���; ���
�ݻ�99랫���m!;�Uu�Z�=#����u���>�n����]�l;�ۍ�و��<ފol�&��6	�:\��9�"s��g9!�燵��b[;�7�����ȡ��>�n^���6��݃i��=Am�;W�M��N�km���다�=:qfv�<]L��\=8�0vɍb���;�1��c��w�&������6Ź:6xw�!��x7
����OQ�y;8��m���;�Nݺ�uP^�حɏk��GH�]�ڶ�q���X��&x�W3�w��r���׈|�C����f�8|t���S|�UN�k���հ�k�U�6��^P\�h������8]���\0W'Qp��i�e�VT鋶�IڹQ���z�ç��q;�H;v����>���6=�Ϯ�&�nk��u�k��󋮝��gɲu���b�=����B\l��۬[9��Y�Om������gV�5�h�m�sf�8���4�s�����c���:NGzOnza��܏%��p.��u�v0��
v��v��̫u�����+�n��M��\=m�V�ECv�����]�q�=��V���Ukd㱤v�l�|\.F���oX�Eѱj�;�K�獭�+�yɉ�m:��We���ip���{2���m]�0��4dH���'(��F�$y�/[Vٙ�Wl�#�^[�x��W]D���=�{7F�Q���;]{�������=�=�):��f�޻gծ�P�a:��ԇm���F4�Xw=��0����B3	�d}s�5�{J/.�v�rY�-�S��N�f�=8G<�</�ٝ�g+��\��f��Nyf���h;u���+�VN��ۀ�[��.�n��8������s��[��-�^�F؝�N�6�t�P�f����Si|�j'��ʌr�F�/\t�lԾ.͡��p�n�����m ��]ۥ�5�`�;�ؚ(#ۖ��=l��:�Փ�,O�nu�ە#�p�m[���zθ�nCg'�e�Y�����9+J&�z��/	;��S5��Mۣ�'v��[�-�[euv���zw�XoYz���^���7e]�������H�����o\�+���V�rg8�����N�0JZ^�,=a}Y7:��%\r��Όw2��Wp(e��Ň�;]c�̙�M�^Mٶ�n�u�V�����n��y��-o��ѣ6�����8*Ltd�3r�z�[�E������o`�@���GfG������z��؀���-�u[��Z���էq��xڃ!�j�xi�W]�X�ȅʉ�*��b��t;v�����I'i6q��n��E�n6'f*���t�͵��,�"��A��;����M��r\�/+cb�`���3����w��3ڣ�u�+�۬��:�8؊.��*�n�m( ���P�5t���+lN�/���)�!��v�=���g���\��̦�鸍��;�b���X��VQ<��<l������b��kW\E��m��N�]s���ym]w\B��Н�v�gfP��ڻ��j�k����������;�5��ʺ.=�_89�ɓ�;f@�܉�]-�m� ���fC7+�+t�Xv��ѭ;(V�K��s�b�=]�FogNG�m�r�β��hS^��gSg���ڍ�m�B��gu��� J������za��Ήz4p7g���ۧÔ��㳴�\q��9�Z�ۙ-�X��&;PA�!D6G[E±�ѱt8��un�j��=��[�����N�\�4���Pm;����":ⳛd���G�q�Oiy<爘��Vcy�e�E�}�s���tWX�ѻ��y�;p[�t�n���(�	v x�ȜdV�9I�wH�0#ۋ�kmq/`�HX7�Y`�8���s�=볳��n6��;��5U�ͣ���<��d]��tu��S�v�<ˎ�j�K��5�I��m�tΈ��,�َ�:��m,�l�]�gd�r3\-߾�#�q��r���m�� pt�r���bt������Vv0�D����H������:�(C�;ͦ����g	�ۧ(�����\lv�ڭ%���)8�6�6�kNAeif6�ݸeh��:� V�����P����xi�	'9,Nۛm�)����޵���D��)%�m�E�ڲ.�8������ͺ(�!�r9 ���"�'���q���);��l��N�N9�NJH�+N�7&hG:\ �t�&M�8$�Jgb\'IfP�9fv�8(ۭ"�� �N8�p#�;�mM�I-���m�igg"e���'fA��� �ka���f�s�(�#���t�;"����m��Fg�8t"G:	!Ӝ����lvQ��ڶ�'&�#��m���}��L� [Y���h��i��9��qۣ>�pu��u�E��g[�=�:�8��;gl���r�ֹ\�\��N;NR8㦶퇠����,���Z'r�W({c��9M�W���/!��tJ�%/A���8��	��svge��u���d�IXy���u���a:^�u˳�[��ۜp9��n}�R�FѼ��[]�"v�[ͷ���ǧ�#�3m�ds���۲�����H��Ӗ֮�۞�yC�ް�G��ܜ�s�+�����qOf:;�_!�6y��kF�nNn�.���vy��/j��;g6L9N�i���=�V�<n�
�FN݁oh՞�mֻO�&����ng�ٵ�m��˃���*nm��v>|����N���uy�m>�=9.�����w��5���r��> �$��g�㮳����B'�g����m�>z;m�2Vg���Km��1������k|�m�=�n�3�C��ӆ�+R�I{mŭ�:��ڡ�m�kv�q�� a,M�r6� ��ֻNʠ�)�k�dE֐;r�� ���5)e�������:aה+n��8�v�v9"�9{
SnV�c؎���-��l��֡�I�w��ЏǇ��A�x��u�x�Q�p���u�=\V8�p�	v���Wn.³��Z��Z�vN�����9y��;�s��#�m�'nc���-��s,�]�C��m��r�T��: Z�Q
݅���PDV=�۶�n1��vuvMgV��B�c����u�&��g�9ݝ���v�<�.W��[�ۍ��bt:of��ƚ�g�/:�g'ݚ+d4��6���Yc��'s� �����i���6բ�����&K�sМ��m=���Ϟ'���A����c���7pۭq�9�9�n���z\]��wϑϾr�-�np<]��gf�'��n�4�F���]s��8�of��]���k�z����p,�{�On/k7������/o`�6�=�`r���v���6l��x=��o&��y�W���Q�^{p��796�`q���W�v������c��'>¾1ʋ�8���g1��{�ٵ�g���޶�v� e���6G��l�\�=���8xvA66p�n�>6rn��'<�vp���-y<z{zZk�x{#���x����۷
����[�3}�~�X�N��EW�"�f��m�܋$�g+�lퟝ�[���r���$��؁��3(4aN�ٞU`M(1lX=C*��i$���^O�5~# ~�R�5��/)�w�)�v͂�HՅw�J}��~�+�@���`�z=���gĖs}x	���⬓f��U�{�Օ�V�vttH��y� �"^8	 ���iװT�-P$��x	:&[JȢ�B�W�����A �?=�p��ݑ~0�E̼$���P ������ʒ��+�// �D�@��{n�ݺ�c�=n�+��Y�w|t]'�<7�����.Tqۄ�u��N�����AM66���D���O^�N�	�}��e�@Ѡ/;�����w�'�3̞��Wm�z�R�ޟ:�����6�p�����{S��MN�l�� ��b�hq/������7[�*�c$u ߬x�<��	s���FV���7��8�1��Xo2��@����l�/�| ����fM�L>�Ó/ĀG�[���~{�������UdVO>ga����v��x�����A��=�A�z�e��^�Ֆ8���S5}���6㖣��������9���mp�"��[�H������=Y���gJ�y�P`_*7aᝮ�y�x�>1��v6�;��v�6ʸ���є��%3{=lhv���E�nk��{�y�i׭>��Sz�u���>Ⱦ�M��M�}�=a��Z�fg�'7����ǈ�v/܎�<^���S��� z��v.{"�{O�[�E�L�V
�8{��0 �O�@P<<�i�(g'��mF��f��ZUN���Y����'g��['g��yꜺyG�X���vƭL�r�������wX��lpi��%��� }���
 y>4����┑:�eR�'�n{4�=�g����[�?��Z���>�瘖�1����d��'vϪ�R�PA���~��$o�ἦ�K��o��z�� �}����wS�!����[7�
�(�+H�s�=�:^^�3��=q�P�
E%RYKk����^g���I��U��>��~�A��H#f/ί��1���H���S� �H>��i>���cE*�	�4����C|�.���o��}�	����O�f_��3i}yrd~������uf�	!D[u�X�����<BxSZ�Z��c`����6��S�GvJ�m�n�U0��V�+�`�YXy���(Q����>��� �n��;͵w����1��W�VA��û�����D���"T����	�tQWКO�у��8�d�'tr`�!;��]���b��J����$J,$,�YF�4��ߌ޹�P?z?n�://}����� �}�G{-�����t����§�8{��#��9M��G��뎹�c�rb7�/Z��˳��se`�M��uqbp�J��}҉�UdVO>s��g�pT 7����e��}Ei��h� ��,���w�� 	��cދ��Wړwu�(��  Wr>�>�=��'��wyP\��G�ƕ��2��zb�X�o���o<qd«���A%�_�P$�9�n����udZ�	!D��ʽv�ˠ���A���.��}��s�׭t*����7����쌻m���Ķ_;��y�&�~9:�������P'��^8	'�I&� ����$�T�P��z����;c:8dj��0Wd�S�p�A�ou]7��.A���;�jK�c����R��Wp���f�_����F�W�;��EB&V#����R�q��u��,9��psF:n�c۷r�D�\��r;�̺R�<k\��=m�۴���qʹ�`6t����c��n�vð��q�vۚ��e�O��۴��=��!�s����̹�ѐ��z�,<�G�eqŎm:[��v�F�p��Vqgmvj�3nۇ�tK�1�a'��u���g���ɝ��c{r[��kn;mGg]��e�ą�ֈܘ拱��g�q���-o�>���( iXm��'�����t�:�{z�d�[����.�Ϳn��g�j�@��5a]�ާ�#1��dA�a�y�I�7�����I���w|�fz���)V/W��0>Í��z7L  ;1|(������Ead�t�4��׀�-Į��WH]� �1��;��ɔ��Mi��m�LT(P����&z�E��e(�n���C�H+H��l��3�_&�\槴ih�--�^��W�� �ǡ@Br�*��{�ӏ�wU�3�j�HX4QJ1�>�㮎�u�N���.�Q���r��O`���~����i*>+2v� ׹��;ؼpy�Sݞ9M�{R�� ��^u/,�� i�A{��TZ_N˂]����ཷ^IY���:т�a���ԝϔ2���n+�>p��G�7;2��9m��<�9ͻ�@R�;�=�tr�THU�t8��!z{��  �aT ',������޿{M`�H4�����\��R%������A ����MƩ�����	/'T ���;VyZ���hVG�q:���;�>K5܆��+�{P��0�#�#3��]d��Y��z�'�ſ%tEZ�B�o�cU`T�|��t)n�?P>�P�ڳ�
;_�@*��_��ٯ�RTn۳�Ia�w[��v�W��O8��y��� ��9���-V_�mS[�m��jwCM=���}}e�+����Xx�q������m��ѩm���X�{�Z��-p�����I��(FG�_�~ {Ϫ�2���~FU V���"�F� ����`�k����E?u���������l�����}"]�Eć�6w��}g���Aj��b]�^V���1��캗]�5�#e�&ReK�#���Z��%��A�������6��H�)��Wx�e����ww� �5V>�>���P��C�5W&剂Et2*�yg���V�	�XXq��{Ѧ>�aUA~�M"}��<��f���NX}}��˨����%vR��;[��g��99co<����4�鎁�WM�s�N�.������y'���6������ ��Ъ�Y�2�cۚ���g{��]���r�)o���]����2�dH$������
�w�� �x�*�'�{jK�g�t�ɶ*Y�>�F¢��IQ�f9�i��9a$�n`ۭV3�t��m�����H �NX
^u/,�����<�%ݫ��},x��F�ti�( >;�<��*@}�Z1O������Յ��������LG���ͫ����"��z;(�L�W�[)V��턼oF;�>����b�>�7`�\�ɯ�y�]|C�g+���L��n�
�_:`�y>Y� �'~�V��E|�:�VH��b��/��m6�n۔����U�=�]�g5!��T��{�heE����n�$����I$�׎ G�W���K��{��H ��w_5�9�b
Q��i�{��v�dr�Fm�sr{�w7��O����|�|G��К|��uJ����W���r�(O­w�c҇��yX��R�8�����m6��wt�?^Ok���5j���I��$���B���"m +�Рx�g?;�+�x_�3�{K�m8�|V=���%|���4�~Ϩ��c���~=�N�{�LK�Ik������̞b"�= �({G�_r&VJ�:�G����<��ןyw~�ب��V�aڿs��;�s}����Z���[UY����Bh5��\��v�P�Q��#UT*U
��b����"��\���tc*;OB]��)����Y����-s�ۮ����;��h���\�÷lloQہ�mWO\e����������D���BE#�i�F���DA��N�_c�]�0d���raq�t3�<�qڽ�c �H=]�ٮ3�qo7j�*��Fwn^k��[�Z����a�rv�:��vO��{��l��4�jˆ�ۋNхU7�D7e�X�u;�q�'�9`+#�~~�yt�M��w;���]޹��j�7�+�����:oWJ��NfC��+��}k�Y���]>� �����jq�k5_Ov��|����.�������������۞���;l�$�����&�d7�n�鷈5�w{��}�>2Nٰ���b����g�����Z�b��Uf��5�]������Ő@ ��7����߯��{�����:�Jf��1�u5j���-oXff���㻱�w���w�|,�@)��� ���ր�߯�F������v��hW}�%��<q-Ӣ磮�v$�mN���v5ۧ��%k?�:i�&�{��^!Y�Uc�k�ss�1 �{�~3 ǧwf�������5�s|�̃lKݻ��n`l�,�,-�ߎ���^�x��a������c�Z���Ap�Ĳ��Ρ1��|��W$S�QT_-NJ��-G��nP�{E��΄�vv)і�~�7�Ag=w�3�lA���A�#ZM{����<��.�c�_?e���2g�}}�`��=�n�@@ 4����H���ߵ{�@ {w�� {�wJϪ�ςGkb+ˁ��oB޸jz������ ɭ�� s�p�@�~מs�w����II��]�b�@9��p��QKSlX�ɸ�Obɑ���$��\o=���xvrniA����ϡ���739���S���$rx���x�ŸL�m]�+'5Z�&�ݭ��� ��>��&�U����̹�0m�����C�W��3��nߺܬb���חT�w�VF�ָX�>ss��@3׽�o-M;��=�k ۞����*=�n��J�uA���X/�ݪ�*��X�nGd�H:Kra���=|�y;�<����d73��+�
w��+h�%�%���Ѡ����~�YCo���=�K
�Ď�m�.�P�S.��4E��C.�E�xAM�8�s�}�a�p!�n.�Dӱ�*�_������oz��( �f��ȩsn������:@tz�����z����ڸ���/H�o�ꊄ�	6�yԂ	���/qч�P�.���V:fw���h|�们�T�H'��=u�����Id��8K��{�Ӽ�78�H�2���C�������:�����(L"��u�:��cK�S�R�9g0��CD�y2����]�Nڷ/�ֻ��_]Y���*d@�	g(���m��
�fZ��{��Q5�gX�,j�[ùH���e��N:+�a;�1[1�^P�X�����S�܈m������sZa��dq�.��98�	�n�5݉eHq�|%�j���SjД��왅�3�����L�)M.��j�.�gB���v�>)���:���ըO�w�L�be˗w�־�S��M�&��+�a�Uk��1�/�F�w8s@�Z���o��v�+�s�S5�i���d
�ù����K��\�b�F�\&M5�q"�.�[��	l���ʼ��P��o �h
�Θm`�j�nt���Ұf	��-��x��k([���sZt/�폶�i!��i�P���+#d�1݊qT�ko���:�b������lǔ�=�&�dn��\�i�\s�E�\g5T3���j��	���ӣ�)�����n���}�����՟}�BY��'M�,�ʷ.N"�(��S�:D�I9,�BR�e��$��r98��!3w'-+s2q�'pHdƣ�Nr9qJ9pt����\���C�H�E"L�0�'$\9I6Ӥ��P� ����N\3mEm�G8fq$Vؑ6�9�[$�S���,�I�p�%���M�\�3Q9K��ۈ̉r�,�!,�せ�[i: )��m@�(�"Ie`�YڳQ)s3�����P�N:R��8��q�%�ͬ�q���	ܔ�v�kr8��C[B�$fK���jD�� �hs�[Y�e֝[Y��BvbA���Єtl6	IB  �pr8�)%B8�8q��cY6��GN��h��X"��*۵�hf�4��u��rw8A ��%4�m��M�Bzոs��G�&��o�����.o;�ӗ�V���&#޾�_?q�.5��OM|��߲�H�]��百{9�'���_jd����i�H�lEyp;�M�@ �7|�{�f���}g�����N�(6Ͻ���1A��3ϴ����@É�{cӆ��Ϟ+g���y�ng����������%�y�QKS@��S'����wF {�������W���ӟd�҃ G����}���ժ��Gkz�f�ر`z�Vm���~95� ]�^��$����� ���7����Jk�S�/���T��X�]��d>���K 9���^u{xo���=� #���d~�����19�*vP�t��Óӑ���r��r� ����,��ww^�������d�Y�9A9��gV_�Y��lK��]\L�Ŝ?�{�r�l W^�V�����+�[�	B�Pծ��r�Z���R+8 ����3\��*�U��f��{1f Ó�_B'���v��k��>#s�sw�7���#s�oǥ��cƟ+҉������v�UZ�-�Ǹ�v�j��pɍ��lv��HQ�У�����I%LE}�A��o>� |�t�`|@�{�i a�{��BpA}~ٜ�w~�������V,Z@Ѫ�r�+$�!C̺g�*K�@���t�� ��,m�<Wy�yql[�9��s.�� 
&��yx	�u|��@�{v=|��Vw�s�oڳZ8����y�$�n�}�d+,��`ݫ��5ߏGy�ѡ�B`E�v�Ł���������^�x��}��jǪ�RQ@���t��$��$ɟ�y4� �ٹ��֛��k^y� Cۑ�����d4�6�ey����]m����IY ��k���s:[�ʵU'n�\B{dR ���IUjj���c���7՗�:؎y�'����{Y��^�[AhDv:��^�Y�4&.��v�=�\�r��vv�oF|uCu�@�1ە5 =.鴝83ۮ�=�g���n��C1�x��=�A������5�V�ۭb��[7�;s�6ùUܙ*��T|m�C�\��yy�x*��+qkp�^��Ө�CY]κ��S�9΄��Y��K�^��y�=���v&nں����v8{M�F�.�R����h�N�u�*�TQ;)%��B9-M@e�7ζ��1Wl����r���|975�s���]L��ֺ�k�uw]�߻!I@~W���H:����w�x��h��vwzF��ܺ��|��r��w9=� ܐӐ��yS~|o������E-La��fNQ��fr{Cm�u��8���×o������J �<�e� Тh�7���E	�P��;�m��Q� =��a��s�YR{�rȋ�W�$���ʪ��*��4�%�1��ز�_=>k���I���rV��S5f�����@w��<σ��z�s�r���9#b���d��.ű���|a9F/l�Ł\������������mnA�[��Ü��� =���� �]�k�0,��5��{;�֐l� F���3=[NU�,����⇾wwz�߬�2x�*Ã�V�&'��RCU��E\읮\y_,��v��K� ���,=x�. �W[w�G�����Ϸ3i�x']QZS�R*��� aUܿ��bo^������~y���ޫ��!�X���'>RA��G��ss8��_<X�c��f�5Þ��@ �k��7� �����H���r�)j������w9��o�������Y>s���� 㻽��{�����|5��f|��z�j�ꤑZ�g�k5�`$�����P~<k�J3���D�*�t���tUꜱU�I�Ӟ�;�z��������c[����l���n��<����p�+jXw����e�L�,�k;;���/�` m����i5y��L�ǆosِb@o���σ1d��$��V��v����W�X��,��ܾzo> <wv7���k�W���S��3{P9��19T+���sY��{[zx������ �t�y}����x5�.�w�r)9�{�j����q��#܍RUjuY���ӷNM-�)'�\ۻ�W���1��e�V��w��W���˜����~y�������w�QN"<��{���u{�ު|����0��ӻ�H;�Of*��'6������ ����(���A�
ޕF�뻫��<�,Q�秲��g}�w���� ���wu�����h|�wo�޾��7cQJ_�"�X5$j��f�Ҝ�B!�cN�l)Uڝ-�(�.{m�ɫS��Ek|z��z~���u@>��}� �!A�ܳ<�z���-��]�/��_Z�A�\�e-�05��ϲ7�s1zk��>f_>%�b ���� u��g�Uw�����ʼ��7L笀I �p܍��^P@����  jZ�rkދy��}��| p��oI ��r{1@\��Yf��Ei�_�����N>��X���=u@�'tg�|�3^y|Jjz�wuR�[�1'{v�Q䧢2����`�35��2,���A��T$�u�S�u����}�U��7��)#���IU&��S�����O��9`����:�aJ�Dz��ɼYs���,Χg3��oR]��#�[�@ �y��ww�����@���r�B`YHN��g</Tx��<óP�;uX�|Gp���Wn:���z����R�7�3�T3�;��@{�מg�=�9�뼅���n��b����� �7�&�N�+[�5�מ`���E÷��f�v� 9��0��7�<��3M�<f���9˪=y�8��,�e�k>ss�0��|�� ֚���Q�L�מ���>=̝̃l^���ً,ت��`ݖ����Z������z�=��@{��I�TO��~�����ᧅQ����:o�r2�#+Nf�����@ {���P�`{����ը��ݻ ��y�U���߻!U��ǧ�cgh�n�J̈́яf�1]��F���&6��������O<+;o���&�W�>��(�^sW�pּ$$_xv��{XG��F��v�{9ɉ3�=�;������;ݶ�Z��w�"ܪm�ӎ�@�ѷq��mm��ɹx[�C�Jy:[�7.N8�؇����Ml]��vx�pU�m���	����r�yD��^
�!����k�s���smӎ�Pss���k��َ�ۍװ}��:�،an��O0<$ok��V�|-��3���Y;P�HK��G8��[�h�X��g���n3��ӱ7v����w�y��WTU�*<��Ws���؃��t���wM�l�Uþ��"�sx7��oسvu�b�qKP ��.�$Oy�}��8{�]�  s��,ϐ ���	�x�(��=sW�����j��c��<�Z�bϖ  �ٻ�� �,<�ohM���緋1  {�tzF���XQ2سY�[չ������}�,� o�t�6#�߮k�����*w*��^̥���k�新���v�"���M�@����n,$��ַ3�ξp}�Y��H9ٺ6��߮��w���{�rj�}E���4Y�R&�Zݥ�cmɶ�kkXN9w@њ�ý�~����S]��V��s��Y� =�n�  .�~�<��C��*w]ssU.�����W�w��k�N��N<�����`���/,�,�z�~�mRr�����JN�͛M�)�Vil����g{}�vp��w9�먑b��Į{�N�S��fR�ϗ�/���ޗ��� �G]�@���o�ݪ5U��y��'3�=��m����U�-@31�r��6 ޹�wg� �N���#��^�ww;!_e���r���XME�����I�=lѾf�����'�o�|rr���A�w]��ҽl8���*��wwz����7�գ*��j�|�Y��� �zk�}�Մ��6h�����|=�Of(1�]x�@wsݻf���*6�*j@?�ZwD�b	`�$�BR�k;�>��z�x���\n�{���µ�l�v[��{��H >볚1 ������f���߹V��eA�����볘<\7�2"�;#+Nf����,��9���kz�^rћ� n�pĀ@.��L�R���{Z,���yn|��i�(�h�q�ă���Y �禞|���FO�o�;�yE�_PIZ������m���q��c�3�Y�n�]
uT��7ٻW:ݡip���Va[���z����'� ;���*�UUz�=�x����3�_�) �9j����Xk=[Է-6k��� x��� �N�
�mN��̻�z�:k2<Gk}�թ�
J���Z�����S�J74�s�_U�>^��r`8^�k����?u��7坓��5�,�Ƿ�8��srq��m�؈ω,v�n&�Y���ϟ>w�6j�k���Z�v:���~a�g�O�Y�����ٯ��,;ǹ��E�|�������b��;�)\���p��To���M���F5�,�6v���� �ƻuF $=���}q��wD�yP��p",��2��k��f�$���� >+�����=:.w����k�1 ��n�}�ƞw⍖��\A���r-o~�>�7o�v�,��������ɧ����#��w��jϒ�mo76��=���L6�6A�kl�<u�e{�6��;����K�F��نZQ-惂ݟ����䖺���<�>����IAȨ�m�v�B��wp~\�j8D
����U߹��� =k� ������^םN���:�o�O�|��wԸ`��;���t��3��[�$��n�=����S��x���������%t|��b�>�� o���\���{F�ff,π@ߍvǤiwOe����n�v�j�������y�o4��> �5�4��������w4�6�.~������~�9Y�g��n��g��>>�34 <��s��{�8��4�����+���(Xݑ��3X{�~*��4f��nS h7�6 �ü̸ {/<dE�㧽�v t;٤�/z4���0�:�y[��s�f�s'�bÇ�U�lx���7�4� ��fe��_t�\>m:a��TZKK\-�{��:��ըZ�Y+K@6�7�f���f�U�Ĳ�kmN����z���w��pّe�<������GÈ�6�!9��j�^:Ye��q펬���R��1����w���w1���=��"u��w#�����ߤ����[�b��2���F��쫂Cp衷u@�^�YNȳH����Uv82��Ѻ�������m�W�B�(W1���pEV��[ͫAq1��wMያ2}/�u&	n��V�k��S��$cMջ/�VS�_`�X�{n��h�;���S���g�e�G��5�s.f��$ve
ϲ˕�F�Xe����ލ��>y��S:_g[��4.�AC�C/.5�E�轼c4u��f�씤ܾ�ivx�x\؃���y5'E�m}�Q��<���h[��h�`7l♘p�� =:�kn�v���H�\w�Γ�'fS��pghq�������T��;��)n���3C&�J����!�R�:�V`g)�;Z�W�}.ZI^D�5̔�dFԬ��z�v�w3�*Af�ޫ�
Ĵpj6j!A�g�B����\�oN�e6��$oo��A��㭁-ޤ��k�
5�v��h��G�L���5ے��Їb�Ƣ�z	{b��E�dA#x���*tt�y�lzj�n��h&��pZ�IK"�T�"0���G����ʟjU��-&`��%d��f���ך�_D"�ma��;����N7-��{���3t�e����m-t�{�U�œ8A� 9��yyk��MnraY���]�iqq61��t�m�ݶ�6ݵ�$��rs�j"�8����r�H(��%m��N���D��eہ��� �BӍ(��۬GD�p��$�+kGE��pH�-��9)9g'i�M)l9Ѷ���mbsn�n��Q"Iܔm�X�Fۋ2�یA:B�:
!���$��Yi#�����'�I�D��B��!8e�)�����w��#�mc�(��9q�JHrI%�h!��:�JP���gu��a�&i	�qNr�0ͻw9S��NHG$���	��ggB�	�:\��%#��A!gZts�lE����!3��."̃�����(��L��I��䕲  �}_�V���졳�S������}v��}��X�-[�r6mDVخ6�b1ۮW�s)(�5��tl�p�mݫ�dVxk p��p��rZ2�s��h[��Y��m�Xxlq��;v[,�̶���:�/���A���k��%�<n���7-g,[qam�yJ�/���7;8�7;N:9����f���x���gۙ�K��'�k����5�����u�N�v�a�nt<��a�áܦ�ѓ���xx֮���λ������zz���.;;n6����/��p�S�����l8^���K���z%.6�ζɲz{�Ϭ݉^B�u�}#�����δGX�m�Nݗ1��DZz��\1J:ڮ�(��D��;���A���Q8�	X�`A6��/M�\��l;
lZ׮����uN�nw���\e:������ɍXї�N�8�R�a7*o6��ݩr�ڞ��ڶ��;Q�;r�Ѷ9zc�EN=��s.��ڽ�A��E،ugu�9���o<�5��:,�ts��X��/i��tkp��^�ƺ�,�6��]�N� �n.���Y��v�ckp�t<��mg�s�����G�1��ƍ��ѹ��]��m�dKv����78L�5��ks�N�]�3Ủ畽z���Mы��l��r�����<����z��9'�����[������=s��5b[)�]��`1��g)���rV��p��Y����[����燷�hN���C˵N�N��pq�X�kkx֑�˱�&ᮗB&��y���|��'m���3��N�7 ����`�� �N ��8��g��a�Ʌ4^in7mq
��'d�[s�Z[��F�N�P��F^�8�k[]�{��W[/g%��^c�Ƿ;`��Zô���:��h��s�6�c$X��7��&N��%˲) �7Ps�N��$lv8��^j�v�)�kp.&�C������Qk�u��09�cuuw䄄��j�4�ӗW�Kw��N��9͍���.�Z�'7�R������E�]<�'T�Î6Yfń;;��8p��S��!�Rv����K�ѭ��3����C8�ܛ��c8.�]S�]�ݮ��c��`���<kmVc���ɹNwW<y���a���kK�ٹ諷m	n�g.�������{'�uW3���V�q�8Y�y9���R۶�5�w|΍�VKo݌��ts����vö9�:�����n���d5�������"��Ts��Cۑ���w\� ��y�0yz���a�ߦ�Ā9ә����lj��I]b5�<b��7��V��= �^��dϐ�sư���<�SOu�7s;՗uj�Jd
��ڳ>t�50 �Ox���L~��3~�gq����� �ޙ��o�9�X��9��W ���#�'f�k����5���|�����b�{]y�~59M�w�W�o�� �5��Ϡx��8�cvFV��a�{\y��|595mHt���t����` {\מb zjrj]�/2����o�Ɏ�b'[��]ga��p[.�ԙm�j�Cb�����HT*	�s8���P�����w[�щ �s\�x� �W�����K�ٞu�rk]Pm�^�z�9��:E@F����Ϫ���/ޡ�>�헓l�\z�<J=��šD{��e�9.��ͦ���g_.��5����{�L��n�Sz��\��94��|�����OW���T�.k��� ��&��s�̳j��=��v�y�*�^6:�#�I]b5��<�@ �٨��_k{��#~�7�^�`	 zjri@H���+b��H�I��׮t޽�n�<w�� i�ϸ6�闰� ���wa�W3Y��8\��y�ǬH�y���r��%Ǉ�N���s#WZ�s݇�P�g���Y�k�0 L��z@��s����]K�׮����Ti�/�*����v��{�r�Ón]��љ�j�;5�[��}���Mb�r�������\y�b�95� ��u�t��*rh��z}�����=4�΍>���v�S�W��.,�9��o���{{�y�� nL��w�����.��9.��\@zw�1t���t9�j���v��7W��r�˂����	}���߮�z��y�����&.љ�4��-�Nw&�U�tˢ���}N�h\ԡ�{�����{��BGs��m����J��WN��+��v�y�<�lu�GP�y����&fT��u�H���M%A ���x�.�f�����^�u[����
��$Q9$Znw�z���k�aw�	��wypbzN�M| ��\ρ��]x�As�c�ߝ׸�ޛip�f"�6�C<�����$�ɖd�u��MZ�^d99z�9�<�r��%�{nz�� �uۋπ�����k��{������nb?,�+t��T֟�;��7.�������6{����r��`$���Ou�b�-���ƟV�ѻk�Ǘ��.` ���6|x��7n�3.zM|�˾\��rkƱ �=��
O���#P����N�ZY��� ޹s >�����2[����1�1n� �u�p�%���z��+����>�k����ܒ�_d�utþ\�50 l\2Һك�x�eCx�ݏ��$��L�<��� 'S���R:�YG�f�xϰ?vG���\�kH���v�z�n�| ��Lm���d}�qd���s7�f������aw(2�c�8��6u����dc����d�#���jXf�<����U��W�As���`w�^3�>���5��Mo��o���f^r� b�kƛ���5��/ä�߃]��*��1Ȩ���5o��LSג�EU >=��y;��ߴ�M\��@.�[␱:BE3Oޝ�Հ�rj���A��Qk���=�����_a����vj��cO�b*j��q���3��&���.wS����`  ��gf ���X�p�7�A�v��3��i����ߞb5nj�7�v��v��ō�}��� �3�_*6þZ[��1�Ϣe�V�V
Y[�OXD�L��r��ܙf�|�->E���{+ҧ��l7�״�yk_c��(^%��?$��d�N��{[�����OzX�j�!�/��]i&��"�G�Xڛv"��g=��pr#�p�N��ܝ�����kq�p@���jw<<��u=n��w9�!ݻkqzד��_ce:��8��y�m�{7�����0�۴�/n@��B��+��Y���8ݛ5pXK�獻j��둖:����w����dXط��M;g�)8�:�:��wYѷں�X�X����۲��Q騬���N:��WJ��(�d��%�<��Z*�uGe?#5�m���zk� |��ky4�glɨC=�k�1 7�ҡ�,VUS��K+���� �]s]T҇.?k.��}vF���y�]��~n��瞖L�wn]��V9RuˏC;#� =�N�@%�;������׳3O\��6�rk�0wڜ́ë�r'FETS5����Ϋ���w<��H��� ,ޯ�π���kg�n�n/��|���Ƹ=���k�Ǘ��� 9�f�}�Ǐ�=���]Ǿ�)'7&� �ս�I�{ATi/sv�ooz�T�I`���9^ۚ� p�pw%���v��퓈�6�x��qi%���é�V9>�O~5�H ��d�Uy�i%��U{�=^|lVC��� �rw��|�j���h���?���f^�;�U��<@X�������@��Xh�k?(��k�Of�aֈT��o C����Lv�q�r���R�z�l��������6�=�ϕ�@}�e��A������ ��=��ͯK��Vy���U��N�A~���� ��V��ird�$o�${�=�m�]潋1 ���� 8;_ιq��wqw٦}�w��&�#`��qf =n*���9�{�@�ܝ�Cϫ�r'FETSZώ��t��U��ܻي��D��ewk���a������ �ssJ��_qUӳ8��gtm�Ke���(2�A6��67XF-��f�c:,��S-����M�պ�xEM[]N=��y7썉9��f�zNnM �ޖ������;��� =�{g���a��V25F���3�J�����}�s~y̚�� 	s��,ρ�<wwK�0�_y�M�R>ɬ��<�2�G>e��<�5�ŋ >㻺���q��Y�/ƽ{�l�	�l�C	2�R�n;�h��l>[�D.s���Eg�1n�w8q��J]wu[��|K�7��g� {���0 ~;��o�X8H��p���+���4�Ky�q�o_s��ŀ�H�e�@|=���
sWW+#�s��� >���8��5eǁ��t��=���G��w�f����j�4����˯��>���*�����u��;&m�W��n���|�����.4l�n��Yޘ4�2�it�x���s�VJ&����9�:*�U���U2�2�U<��l#f��Өyn��  �̺�ë�0EM[]N<��mE���o"�{ʱZآ�󻫰.�qz��H�=��F|�锓�<�s.���=9���c#��H4owJ��7OwS�Ѯ�r�5�wSu  x׮���{��Q�'̭Qϙ~�X��v�w��.��įUr��DЪ�=�F���=�-��.osx>����2Z]d�2�i%��LKg&�+Q�l�J����'Rfl�]�v3�WWYT/"���"'�m���jk.�!���8_^x���Ȫo\��J���uU%�wM�r�����e>��}�-=s�i>�N��v�@ S�̣o����|�fi�=}{ީ�{�������Ӻ#E{�++
���m+vt���6�s��kE���������qk��.��ڝ�P> ;N�P���q��Eֹ�=:�&��d�m�W�0��wv��$
��W���|/4c�B�����;GπH2���$�vs^����[�3��'gn���h6"������g3+`p�1` ���ϛ���{ۧ Ht�27�zs^���y�&9X���s)���i��ָ����S ���o> <k���ׇ�V秓m��٨������8�/�A�ѭzo����QFjk����I�����ߕ���πA���X���(�*{+zw�x�r���fY���lK�P�ܕ�*���V~�'I��D��$Iʫ<�[Y�'s�љ���}���6�J��gvf}�/\�߄�����i�#���+����^ ^����
G�䫄5���[�-�юN�.�+켇�1�Ee�{t0��n�z�f���/X�Vs;��wd����N�I<�S����+�5����E��k���H����Ş���s�ǲ��B�W^{�d!n�<uu��U�v�ܥ�Q��E=Pv���7=���ٚ��$%��5�֍�ݭ�)�O�>:�Ȯg�b�:��N�|]F�n��l��պZC5{��[�uR���Ato���	���>�@ z^٤��%�pN�E�+o��< �>��wu"!�X�d��,?��k� B���F�t��S�l��3 ��{t����GW���xy���wޥC�$�:'eDS5���zf  �^]* ��uٯv�w���l��36����؊����yq�3�G}�����@�s&%���#r�� ���sW�յ��ݜx��Lπ��80�غ�.�ۻW!F���������7����3>�/.��lG��34".��s|���~��N�U%�r���S��䵩�[�fvϣ�'+ӹ�+��_?_����m�@�2s{���|/��x��V��K8��w[���0 ��ҡ����Z����7�y�'�E��Dzv���S�s&�gN�ܴ Z�mg98~t&���x��2Kb���������ǲ��<)�[��-˯��%�޲r��}�9��&��쿬o_ �s3Co��,��s\�{���꼐r0��՗ ��*6��s4  ����zb�g&�n{> ������^p��9%���QT�a����j��z-D�54� ����̸�v{]��Ú�-��ͼĀFC{�T�δ���SWW>A��s3B 8{]����~*<�ތ��9�ԝ�� ����J�^�.������4��;��MU��.KC)�<�+���;v����] 7n��.�<��]�\0�u��d�1J��{sJ�7�y��4 z{]�����9W{��܈��f��8ｙ���̭A��~���{&��v�Ũ]����;Ag�/y�6z_vf �����.�VM�x��T2{62��UVY1�N{�,� <_zi��}&9)���qSr�Q��˔��= YY����]�ȏ5�>�&�2���y�.������'&�;8���lh�\}2d�|n��n�VBI�l�/������M�[�Ӎj��K4P� �٣��]��M�I ���V�,�����L�\�Y=��U-�|�:�zm]Zx�:U,���
qaY�[=����e�ʮ��,)��]���؝T��J�����޵�u*��5mM�R�Mၥ�˟�bFp�h��zk�����뗎��&Ր&�K8�
�����_��զ�G��ܛ�����}�H���0��E���'�����Aܬ�tJ�`�T�g�,��ƫn���Tf��g�A��Rh;UQ*7-�K�K�qYS�-�x�\��Qe�^�I���n�V����|�fZ�k��	��WNH�b��o6�U����Ι��C32��o7�;���j�\���J�����zgI,�oEg<�r��t�:���
�k���D�l��ګ1-VυL햜h��V�ھc].nue�,��WBDE��ŅSV�u&n�7.�-��"e\\qa�e�)ޜ��YDͬ��3
�Ld���:�ovL,[�{�n�Y��e�:.���������c��U�q)��\m�6^T=��$��7��t2>�nIF��Rgb�a��
�o�%�c	�On�&����ﶭA�G2��=��_�:�wK�J�*n�Pԓ�YMJw-�� �	[�O��7�Em饕Q���yZ����y�@u�bK+�/�LD�o%�D�m��c�9p��mX�.(�D�q8�ӉH�*Amc���z�r�<�rr�$���j�:;��rI9vc��ok:����wE8�-���9�D����n�'N86�,R�tJ!	(#�99:/;�j����P��6���J�Q���
��=��{`Q8��h��A'��%�{Ze7b�2�re�';����E�Ͱ�I(m�l�dy^��p":K�����Q.��DD98�9����km�ː��!ͭ{{�GYEDu�!q�&v۴�&���e��(ebpL���Gn�pE^W���UC^� �3{˞*��^�{��t�K��X���#,��Yq����^�4�����kز�����E�]����ɞ�xp��ڻ��둲8�!k��U*��Gg=ɟ` t�`
���<�WP.���UW�+�l���-O^��UP^���ۻ�d~~y��[��@nq\k��'^���\��6���i��D��	�w�y��M�jN�|�fS�o��f}� ��Y�X���8�^�(�l��>�>@v{]��v{͘6J����ˤ�|���;��>W��7�� �{9{ ;�_B���j{u��z�P"�^V���~�bFMg�%� ?��T f���r,߯&$zw]�� ��<wwT����USUUYd��.�;�ط����4����ϰ o�t�6׮m���w��T��z�͠gM���n��f�Yw`3x����f�=�띛����9;,��
���ͼ�����h��w���1�-��w���|�HK-�+��k�=�o*UT]�˻�o������d~S6[4B��y�0{�w_A�קs캫\�8dA��TjH_�c��H���>��w���ú]���0��શ0$����'��Z��J���zw��x�@�ɻ� 	w^��{��*��9f������ ���u��Y����˟�����C��x��5����@/N��H �zw2A�to��R��߉��Bk��HY�hύL����	���� �n�i��������@؏OM�� ��ә���+L�!߬��2kۙ�n�k�A㳓PlA�nwF|�M}���M-�j��nvjj=�A%U5ku�&�5�Of@=�wކg;ٮi�^�%��h���;� ;9�߸��fw�FE=Y�8H<��hp��D�{���c5�xV���d��_��G�6��x[��3^*��yX��ʽt�u��(�@�,����Qʻ��jU6���V�9��^*=�	s�v�P�����,<u/���U�gd�t"d^��6�
�mc���n�	�x۱<ۗ�v��V����	�pvs��s;���vK�ku���Mu��!��G�t�m�i`v��
u�9�l:���v$�-��̻m{n/l���jح�ּ�&�-�糮.(�{:ڞ^.։�q���i�э��� �[c]�{�=v]��3+�8Q�����%J)n�ٹ�� =���� ����d��l9���3��9;7����f}>��p����Uu�{}���/��;3Xrjg� @|���a� ~��=˼��.o{ҷ�sP>��|+>����q �59� m�˘ z3�!g�{���� o^��P`y칉�g����+�R�gƦNCKje�nfe�[�l�5�� ;�e�� zvnk[^���v�K���Fs�3>��ߣ��L-jHf|������҇W}9�ɞ�ٷ���	{޽�> ���1 =;75�(�߯q�[��-u��U�@��!�(;[��#����➵q��.q�ҦR��.ə�u�Tխ�d���'s��� ���wri^\	��g,8��O`� }�u��u���k�"�x��r��6����^M-���i��̧9���l]Fx��+�;آ�mu.&h��T��e�@;�1i��W8����m��2����������fk��?| �k��@$�wt���s��Zn���⾔u�%��#tKU*�q��\�ٜ�����=�����y����w.b@ >+ձ`UA�O��aZ@�z��W�H��8������ԭ�|�wf� ׳F�N�ŵ� ��z�x�9��G	db�03>��n�w2Nw�w���{��@��7���F v�5�Z����A�y��-��а.�Y�hc�5v�Q�T�E�7���n�J
�*FԵʊT�}��}�1T�֤�|�9���� |/�k�������`-0�4���fghR"��o���Kr�i�Z�V����A����M�G�޲�[�qB����� ��Nf(1�$�%�p\9�{�����"	$��q�x׮� ׳�� z�n����^�S>�5�78�e�BZ�����ڴwvY"�N.ڛ�6~�a��c��0��N'r��Ҳ5%��/ua]n�����ꪥ��~�/lo_ z�������e �U*�q�����1�~W�w� =��T�v�� {���w���%^1u��X��:�ej�S�e��59� ���ŇӝKZ=�L�{�n^{sz>,��������ܺ���[��k�&�k�9��5SDeUWa#����y��Ң�u�K�(��Q'K*u�%=�y3��QJ��A���� �OfF��ww~t�������u�׼pWa���&���(�J��kg�w���r����7c�����@|{��uwwg���L������Q����L�֛��l&`k\�ш ~���x��m�sd��w��6#�s��b ﻗ3�7���l��V�-ǁ�]��9�i�s�ڽ�v��H9�N���e:���ָ�)�	��ǉ�����7RNTL��Į�� �wVr�G����_f��'Sa�@���;���(�{;"���b*O�|>�}��'�o�Oي輸�,�0�R�&|��n`of�c�^�Qˋg�ߗu��3��� ��n�;�__��5;��Xup�d�ݼ�����v5]�7�H;u�녧�n�m�w��l<�떧���{��Ĳ6�{�� ~5�4����f�s&�>���ˬ@v{ɜ��
����̱�3���թ�Y�Gy��6 ?w�N������Z�ؿ��F��b*߷ӻ�
r�<�R!��9&g�Of�` �]�����Vǡ_k�ލ����Lρ�<k�=n�m9%�7jn���ק}52=-7�J�߻�k��&}�����,� ���7�V��%Ų!�����Lσ{�̌$���E�;��� �t�[�o43I��� �k^��}5˥F����ϡ�k�f�À�� �����>&��u�e��i�%j�i�k$��uL@A�z�V���jq����Y&�Qܺj_��}��)���~��ٺ>��\�(t�����~o��|[�n��)�8�o`�8˃�9�{;m��"�.�m�p��)wg/��Ƴf�k��ӕ�:��\.�6Fx:���ז{\� �q�v�D���i�s�6G�մv�إj�n����N��&���\v;4b]���gd3s9v��\mκ�+v�/mc9g�Y���4�-��ks��w\N����y�x�Z�������םmɳ���su�Ѱp'�4��� ��7hH)~�F�ӟ����[dp�R����L�f, =������}y�x�o��ֻNs��&` �]*�*7�j���ˈ=�Nb�|p��z����ީ�d��@ �z�| >�Nho>	�sx����&�{���oɛ��
��׃G7c� 7};�@)x���nj���1�@|���uF������:ȣ%���{2K|_.� ў�� e����}~犏��.�`����W`;��zs�NI/�ڝ&�.�;�,�� ��d����r��r�٦��Oz�  =}=�ߏw&��÷	�q���K���_�_ߛ�~d�)a�N��s�W6S�h�·�@�9ԼV�;�߿3ф%��n��5������@����ɘ{��%Z�yn�4�ը!r�@���P>༸�-�Z�K�L�f`{D�/IW)��N�koLˡ�l#����r��^�0������i�bEq�]��{�`�>��df����*X�WPW��.�ֻ�/��z5����|ݽ��Ā�O�ə� �ٽIv/L����=<��ڭ��r�{��ő� ����{�췜oݛ�Ùcm�����1����@.�y3�C��U��n����[��js��wY3A ���f >���c]��}�����N�@\������rf=���@ߍN��r�^�s�";陠7��a�$7�e��zjvk�r gUx�7!�� ��V�
n���q��quv�[�mN��w����?w�$��ݩвk�]ns2 �}�O ���h>���Z>&zfg�`߻���W20���D[��/dm�橏.����A �;���@ �J�x|AfD4�/Ϯ�D��]�U)u0;��� ��5���������WE�{����iޢ7��lt}�o��6�;uiru�?[����c��6��z��|�o7(��з��J��|���o����>��ˬ��5ɪq��L{-��]\A����4�� >�n������$o_ {ڜ�Iﯲ�^ �f�ss�L��UDb5nk�C��ڝ����&7rgw3 ���f��> �9��3%﷭��_�ۇ[u&��F�06뎧�F�kn�X�r��q��Ք�Dȝ���G\�D���2s{��l�8�H =�^a�s]�{y��f���&7�|r��ʛ�ޙ	*N��I5�}����$�W����V�88�3��5�5� #���b�o��޻�:���3'0�W�0��V�%��/�(؃���� u�f�-�Wt�o`��#z ��9����f�#��nzg�v��r��w��`�z�J� ,�0��vs�0��G��*S�>�Ig��?\��%�r����<��q7&��u���[)��+���Y�I��)���j���>�!$-}⪃P���w� {-��>�[�97Ĳ6���x����ߔ������d�`
��uf�A���d��{�fھ��I��dݷ�Z��)�t��v�M��8�u��)��#��Wp�Ѳ�{�gH4Z
���Cۑ� Vy����f�� �J�t��슌Hsz�̆��tA>%*��d�ni�ཾ�=�A��* �4` zs�1�A"�w[�����z���\��I*N�A�3�'�#bA����v��9�H֯�=s�ܜ�sS��g�}��zf��{�KiZ��G���W$��ܧt�΀��d �9��ρ��rIȼ�����>��{��<K���f�#��n�Ow� 6ɪo��9��;݁9��1 g5���riQ���E�/��6���ެ}[]�꾻S�C���K �{��}.V��ܐ�*�_�»\����^���T՗w�fE�:B��3��r���nh�(b��i�vh������}�WF�kZ��;ҟqL
������t�!�:ةήFY�v�v�R�����V�2d����>��A6�Ӣދ�%V����mP�Y�Ղ]fJ��]���
�K��K�ZV�Cj��Ƥdi�%�A�7U����Y����vʬ�yJ+fvZ�T�]�Q�tq�e3�w�#Ʋ_=P2��ئ��tL���N$�+�UG��7��
ړz��[�'����֘�K&�C:wQӆz�FX8�y�nIϜ��ž��.�AI�tX�N��Gil�0U�w:��D��]W5��d�qv���V.�I�1���J�'%�b��ݎ��;;xݍ�e^u��fE1����}y9|y�oٶ/0�:��2���4���Br�*2���U�;'K�۱��͵���m����7�Ϲ��t*�rԫh���jM#-�������7�eJ���릵'25N*�X5n���]��wH��\,�i�B�'c	;d��J��	e�[��T�y�Z��2�t�ۏ&
�_�Օ=�Wr���^`�{���c.;�ZI�]/��5��5�"H��u��^��;ˉ��o\��u�m4����T�rn0�u��O�{���7���<l�;�8���N����}��M,s�g�Sةǧ�uj���a�w�Ej`���.���.]~k3w����R��4�T��ʧB�:AG"��m����%��$K�q�fHYa�vQ�ؒr��rҲP鵧��[�-����m)Hu�ۃ��,�kv�Fnr�J���pr'GBL���nNֲ$��&�����{Z�S��z��{[���(F݅���[m�۳����^��O-٦rd^k���"9�N<-ȳ8fr��m��{d�Y�Yn8BN�mX$� � ������{h�����{�ӛv��"yۍ���G)�d�Ԉ3u����E'9y�s�)I{b�$��9)��on��E&�����w���N���|ڮ��u�GU�v7�obXk���]��lU�n��;n�wS��o=a�{q�;f�v����6v錎9��v���y�pgs��-ۗ� F,�K9|�n�=�O��l��m��G�'7�7nL��cBv��h1shz���]�ݝj�z^0u6������r�]��4d�g�\�.�m����+\:q��
CK[��㧔�ru�­�*ƏY�;kg.����9{A��]�\m�m�M�q8�q���.�|���s�u���%�V& �N�e�A���L�����sC �;�$�wM7l��mϮ*vn9�l.Ѻ{nF{���1��<\Wd܇[j���-,��ҬD6�񣱍�ly�;]�U}�)�v��P�n�����r`�ppwgc�Hj�VHw@�Y��k���X[�-n��α۳��a�uٹ���ƻ/<�Ҝ�vy�����+��;�xY�=q�x훉|=v��э�si��y�ё�q� �� ���p:���؇NӮ�����x���Xヨ��b ��Mѭ�q�5��Ek����S��ks��r箖�/��w;�Q�aΞ/d67�ru�l���#cu7>nzU����/o=<q��nkSo=���Cd�sg�@�ɭ�dU���V�m�R�֝7Hm���f���Q%�����ڥ��V�i��F�P�q��v��c�]�۔�F�(땳��زں�zg�<jF7��Ü�_�������cʻn���M�ֹ�e�;M�w��g�F�;�wg��ց������uǝ��;m�W=[`�a�X3h.R��'Z�q������9�6��V���l�t�a��q�p����qsGka1k����8>|�{
�͇v�f�8@�7\��T6�:v쇆�7nx�y;p��ۋ���o3͹��l�/W9\ی�+�X��$=��61�s���[8���]�2�Mz�&�ٰ��E���KpI��=n[v��z�0snζx�������'��K�Lm,g�:�8�����,{ύ�4�(�1ևv+�L��J�3���0����NL;��y'�˷�ۄc��7V�\.�q��G�z�/Q�cum�a�pt��ݵ��6Mv�9�.#��89�7�Es<��{��l:ג����9vTx��g��v^�˰�<�@ۭ�9׫��xݵ�����>����lb3�%։��P�R؛�%�Qq�:sv2��6�,mp]���cmG��ܥr��A��Vݽ9�;a�W����sv;@tl�v��?����3�Yj���������,�k�0> �&rF�C�� 5��{'�{9�Mb��l��� 3C��J��s�ڷķ��{$Z�u7Ր@ ��zk zɯ�����)�=U�����v�j���D9eB��k�` �x3�J��'Zz2���5��  ��3 @�rj�˞o$%U�W[�f���pw7�=��ߦ��7��X  ��I���{ڝ��d����/�� Rgrf >�n��%��DK���5���=�N�M��]���y�ٯvk �rɥF ��S��B���.�;_DjƇ$�5Y*d$q��Ǡ�n������q��^^�Z��-���-�~�>��3������O24{��ڍ`<b�A�(���3���HP��4Fþ޻�c�aFI��{W���^oS[C9�s�F�F�5F�����l6�������.��WM^��M8�?k��A��BPF,���ѻ�>���ٺ��;��k	���)����~{�N����3Y��*׾�*��g�>z,�,����҇f��oI�f\櫏�/��>���b�)��F(�ۼ��ح�L�Q��j?~��H�t(¢�FC��Q뇾�Q2��F�p����Ԍ����Um�3���4[���5F��a=�����#�#F��k����{\�{|�a掎0����\�h�-���T�Q�0��n��m�2أ'4x��U
r�M�Ō�F��g��z��q��\k��(�Jg��t^�Za%
0�&��9�޾�1�f0�#0��=���F���No��+aM|�a��I��[���ϻ��od%Q��ṋ-�����F�F/�A�(#G�{��Ʊ�;�yﳳ��21FjN�E�[6����Q�8����F0�T²�]���?vY���,�N�@��gd�(�~�w����n-���81���\�w�苕^���\��:�$�F��{�y��m+Q��cJ3�#>���[6�i�b��j0����H��F��h����a��a.�z�N�����0�-�5s�h�-���T�5��GϷ}�1�2أ!��GU9n�.�����#G��wQ�1F��Q�9�ݕ>�׺���譟I�[���(�8�G3���F`�0��#�{�{5cX5F�Q�a�Z��&�V�j^�[f�F����t�wvJ�j��h���__�0�)(#0����f���b�F(ș�5���N�����?��6�0�r�0��W�e�d��\�'\��~��K2�Q��72V����;F�4Ni���{-}�|9�w�b�~db�A�(�����1�B�*P�	)����a�����o�N�UD�F�5�ҍe��e�Vs�w���L)�j0�{���������a#�;~�n�cF0�q�b��\ϴ[�~����alT�Q�8���/�F3[d>��|wET*U�(��Ō)�s}�[\x���Q�R��3�-��W]�wS�8(Ï�G=�k�F0���dL#���sV�lT��0�Fz�@�F,������qjq���k����������-�Ws�qOS. �F�ONv�A�F�3��������n�ե����J=}��<alT�(#Gg}��b��L)������-�ٴ����������ӎ��摌1]
0�*aM�w5l6�h�#�}����%��P�{F0������+aMm��5z��ޡޯ���\aow��FcaF*aM����a�T18�1S=&��l[Z��T��b�ig��}~������pe�FC��T�p�.�cf24v��հ�5�1F�L��EP��Da�|����}���u�}���0��aFF�j��٫a�cQ�j5F*g���-��C�b;�a�m@�W6���m8ҏ����{{�u��ϵ����b���P����{V��(�Q�221FC�z��b��Mm8����n��1�p�����_矯����'5$R���4�ɸ�ze�n��ډ�1��<��t�i��u�0fbiG��ssi6��]�V�X�V��Ϧ�����>uS5�� ߅�+�B�$T���>հǉ�0�N�����c�t]:��)�3Fn�9�ٶa��5���w�5�-������ܿk|������#D��y�a���a��I�h�-�1S�F(�j?߲�_-���_F���YM����D F��W����������g�s��T�"�gr�qv��/�<{�誔�Բ�غ7>�j���(�N1FJg�k�/j��P��h�#������a�#����9��{���#V3��y�a�T���0�#=s_h�+aM9���.�R�[w{��L)߷}�|�BPF.��N��9�4zo�ռk��Q�2#d]��-��S0�*kn?{kH��L+
0�s�e���!�=��/??�iG>߳P���V���1��Fv���ٱ��F��a�Q�~������L�#�F����u����ﵝ�4`��a�J>���[��*{j1G���5�c1��2/�::���S�.�cf24z��j�ʾo~����w��b����Q��(���轅L#0��0�{�����20�#Pgo��[k~�w���)��Fdg�9��c4�4E\��u�rʧa{�h�G�s�h0x�1IA���Oguo��=�=�$����]ǧQ�˿we�[621F��Q�?��֑�(Q�B�IH��;�a�T!n��ś������{Ε�0��O���+�>!<����i=�F�9C:xq��-���ܖ���j�P�o�7nN���꾞̺�{���Mm��ng�� �{�?A�Ħ��]�;d�9WmX��z{rT���ӭ��G�ɡ��q۶��2�l�-Y1��X7F3��a����k�q�Q�zv�=�k>�0�=�F�K��y��8��g=��8��;kYw\q������t�]�<��5�z=k�w/K�p��D�4����Z����uxӵ֌doX�n�,B1۫�+.��؞��{3�PM&'�[�n92���A���v�^Ҳ]�sv��GA7J�-g�R��|�RF�mZ���)���f�}�ͦa���1S
|����0� ��1S
h��wX�18�4z9��u~�������+�r���lV��1S�Q��i�db��ߛ��:�˒�^�1c1��=��k1F��a���k���
��{������S�Da}�oh��L#��0�A��v�1S
?q��@�ټ*�����>�޸�"f�F���G��t�˪����cF'G}�5�m�1d��RPF�w={x5�Q�1S
b�4/�\�j�M�I�.��'H��e4:h(t��f��uH��˿������S#�KiZ������VF^}�w��4ím��1S
~���#l)��SF�;��0ƌa#�#R�\�z-��~������jK��W�*�W�2����#��Q����L�r���w�lQ�24{>��X<b�G�Jg$�z/t-0�/�9|��o�anƈ�8w����#��0�Fs����L)�j0�"dg�}��c4�4{��~P�5�]����J���A��;r��t	Wk�i�G����ؚ�5U%��J5V����}.YT�/�a��8�?k�֑�ń��P����oo�(�Q�2&F(Ƚw��[�l�Q��x�O�w�b�Z{�֑�2P�
b�H�����#���U�#v�vUV�L1���7��l)�5F�\e�oSU�BU�~�z�R��k>�O���R]�Sl�ˡ�m��wE��!N�"hB,r��]���o����.�쩚�vq��V�G�����_���;��Z?5�#0�da"���ی1��SF8�1E(�s��-���T�Q�=O���y�ӽ�o�q�� }��U�:�K��^�1c
h߯y��1F�q�0���;����(�1S
�=����ܞ��<��0�T�����0Ʊ��1S
a�oE��f�F��燍�t��ӱ��a��������q�7Y�����QJѯ_�j<Mcpj1F�L�����b�ldb�G�Pq��sZF0�����8�=�V(�4{W��m�#��r�28Iwul���cf#>���l�0�D�a��?w�֌kF�����\��}����c#�7��wcF8�1S
b���=�ųT��S8�~�}�#�#c��9���~�;U���h]�2X�"���mrݜ={�ؗtn�Y�&Q��~����o|N����wӬQ�4}���F�<b�G�	(Q���轪�H(�8�G}�oh��F���>ޟ��׳os�L-�3��}��ƣ�j0� ��/niV�5ZQ������7,�
�Ͱ�F'G�}�����*aL_k�k&��s�5�Ϗ�M�뚏�X��Q�21Fv}{�lQ�db�@q�5}�}�#S0��Fۿ?v��=o�#�}����F�{����Q]��U[E0�c��_4[6�[�j0�D�a=�֌kF��a#�\�r .�ߥ���/j�ʧ#Ӵ�K�C��h�f�0�dj����=�VCkL���ܥ�suČ�{�i�5��J�+HV�_^��h���a����z-�j�#8�b�Q��}�#�#d�n�WT�B]ݸ^�1c
h߯y��{�s�n�[��	(Q����Э��(�8�#�9��ь)��S0������F���&��g����]j0�T˟_t[��F������uum���0ƌq�w������,%b�PF�v��G�cxg˙w~���y�uy�����3sw�-�3l�Q��b�)��ia��T�F�{[�x4F����'�~�~c��nn�����ť��b��0m��>7G]i�n�lS�R���ߏ�Z������y�go��-�[�j0�A��>�/�0��#��#Dﵾ�0ƌq�h�C�o�~��q�%�^�[ˠ�T�ƣ�e��c1����[����rۅލ�F`������k1F��a7n�6>�hۣl�v��yB���S0�9��v�a��1S
k�k}�a�cQ�b��[|��ֶ[=�_t[�[������l�
��4��[q��v�Im�b��1E(#G޽�Q�X�j1FA��2�~�����^�x[g�Pq�5��e��c.�T(Q��#�����4F�߽�Uȡn�vUV�L1��Fn����G�{޻����|�mA��5�#�}~эca#��#G�{���`8�4A������D|��~O*�U�{&m�׼�:ͬ�Sk%������/��%�f�=S���6FەR͕�׷�8�>�/ҵ�\n�Ǽe����x^�_Ͼ?��?�F(�Q��/�#�-�2��|�n�.���f����3����b1F��Q�1S?N��^�����L��[5��El8�L)��c�L#�0�#Q����[k�#Q��0�#=^�[��F���{yߙ}x���.='�!�P�Tڪ1JA��ms��s�\ Q�[��+mO�ZC.�o����E��T�ц4~q�w̿���-�J�	A=;�j�m��5� ����oe�Fm��5͜�r�&k8������H�t(¡B�$)��ڶ�h�#���S#��wV�I{F0�bFz�y�ٱ���F�ӷxg]F̣�Q�?{W�k[�#0���}߷l1���8�1IG�}�ŵ��N5�絸��s���߲��m�[dU�}#廹��w��1��ן{V�'�Q��a�FrO���B�	(Q�ph�#��/�?2��������0���a������cX5F�Q�aFz���lV7����
�ʹ���Hs�o4�};�}����}��mJ�	A93��x��(�Q�0�*gd��[��*aLT��}�_�F0{�s��}��c�)��U�={�ڶ�0����W"����=�0�`�3w3�-��S0���a���k[�����[20�����h�8�4GF(J=s��l[F�#8�b�&��}�8�����{�~���uߖuQ��m��_���k��靫��M�5&Qo��WT���դ�ݝ�ab�9:����ĴЦ�uݒ�y�_/��7�n��Rz�����xٴ�%�������e�n�l������������3u2��A�.[g�:�s���VEV#7g%��f�[X�!7���j�o< ݈������՝:�w��\m/W7m�����n�m��\��CE����n�]�8��И��2M<�ꇰ{kq��Q��0�چ�p��<=2C�t�1�G<�:�a�e9��݌::�ǝcT7^ljXQ_V6��{^r&���~w��Hy�e/��|�ᑣ/�歬O�Q�(��I�轔-0�TDa�>�1���3u}�g���Z�}����Nw��0Ʊ5F*aL"dg�>ދa�f�F�s}�U#���vT��ю0����0�*aLO�w�c���8�WϾ֟��8�b���Q�r��lVͦF(�q�0��}�iaLT²�M{59�򞾣�W�k��5�x�G�kS$�*��+�^ь4�L#'gsF���L#Q��5�#���cX�0��#20��yG�V�����绦��q�h��#�NO��LV���Q�>��kH�
b�=|��wr;���Fأ>dh�Ͻ�5ϧ�n�;�wU�_cZ�Q��(����b��L)�0�}�y��S0aFA�a�'}�֘cQ}�*g3[���MF�=;��1[
hߧϤ2��q�X^�ة�9��Z��#��)A+�����S׵�9m�����V��'׮l��l�Q�8��<�y�#d�F
a%"u��B�
��U��y��|��X�;$9�sl����:91��x@[����kD�)�\�諣tc��4���ҍL���L�a���a�F��y�5�#��0��#E{~��m�a�g��>�:����_���0��(�L)�����5�c0�9���;vB��wr^�b�0dh��sZa�* QQ�8��a5ź���e[�8`��_7v���e�����9�l։q�Ց�\[EJ�c��x-{�qyv�1C�]Ƌ��ȣ�����\�r���+g��4_��HP���G�����aL��0��#�L�����k�#Q��0���}�׵����VM�E�����p�U#���u/q�4`����Zx�1BPF*aM����Ʊ�8F(����3�C�(����]-�������Q�8�߹�#d�F
0������h�#�4����r���K�1������l�_u����Ok'���L)�F��cX�0��#20�N���L1��#Dq�b��\�z-�k]xɜ����wЦ*F(s�֑�`21FJξ�awu��w��
h���֚��5b�!(Q���轪.y��ޒ7s3�>$l�,�fÛ���aL��0���5N�;�0ưj0�A��0���Ϸ��m3M(�P���)�[��4�X�nWT�{p��A�{8w��{&�uQ��A���Tۭ
����S��:��u��<8�>k>փ��J�%h���֞5�Q���S>�/�St">DiG�~珄�2��Ǯ&.�c�=�kH�(Q�Ja R'7�u��4F�N��UU��T�=�0�ba����l)������Wi󺫭2��>]a��5���0�##��#G�}ة�4`��L��oE�l�b�Q�>s�t�Ut�zέ?w�kH�c#d�s�#�q����\�����{�5m`�5b�$�FzN�E*a��6%W�u�����h̸A����Xsl;<tnwֱf�,v�+L� ��YWn�`���ֲ'�y��a��T|uTĞ�/�1��W�f5�~�{e�ñ�u:Ubj�Fa&XH�;m\T�8�l'n��ƛ��}\I|<\h�{��� η��|�9�i��1J���t�v��ܹ)��#�D�88"T�n�ʝ{�+y���t�R�q���[���Tt8��҅���v���>j�Ky-����c;T�r���P�|�f�wb�
�<ł$��X+���ʨ��,�G���YC�4���Io4���z�*[����+�$�'���߰25])T7,K�t{���Z�7.���-CW$Ν&u���\'jżх�j�sʼţ~���K�B�:��Ҿ���vU�愰�����]��8�v�Kl�ZtU��&����K�o#���ҲWռ&�$�����[b�@���2���'H�]���U�4+�j9\��>�f��Vp
�	�<;)5j�Շ�f�����P�ެ*�uB ���o�[�_����U����\�Z��ǩ��U�)�P�} <��6Lg��\�wc�Vv���G���yuk��j]�Z�_+�n�St�%u<�{�
�yK��V�b|����{�jނl�T���߹͐�U%�{lff���P��r�Qk%���ga/��#3u�g]\l�ͬA���3�b���Y�EW۪�����
�|`�܎C5f�������޵t�:�H+�K�	�O�A)9����VP��8�2ȇN\���i�ڞj)7�z�K�s;�ޛXp�q�bm�3�ݓ��m;μ�Rq	8(��<����{g��w��yiy��{Z��M��{v[[��=�BD�I+4���^v�������N<��� �eڗ^�2�Ns��$����:s0�en�tr��絈�#�B��gy�c��:󱝯&�1Ҋq�c�ٻ��ד޻ܧ&��#{ޒ�s��۽�2�[���#4�6�9i$f�p��u����n��$崛���l�̓���{w�n��ص&dۦݵ�9"�P��m:�/����0�*aL��0�Fz��j�cX5F�j0� ����*�ƴҏ��o�q�
�e �,�����ʟ�`�WI��2����J�%h��=�x�1G�Q���2/]����l�#j�Q�?}�kH�^��ޏ�=��*(�JF��sV�&��8�Oڙr��������al��gnw4[60��j0�F����8��d�!�5?�Pi�T9��sv���4`��	Gn}�ųT��j1G��{��1���ѭ�Lǿg3�3�z��"z�څN[��T]�1�ϣ��a5�T\a�҉]��8�����?#o���;�����<24z��um`�5b� Jg$�z/j����S��G�{��1�3�f���k��>Y�|a��5���m����MF�dg.wz-��SG���v[�%�/[a���G����c���d}�{�o�g��l�~�s������Q�db�����[�l�Q�1SQ8��sZF0�P�
�
0����{��f{V���G_w�S��7q�Uӧ�Ff&����l�0��L)��S��洍����0��#Ek\鎡z�����ía#�#�r�w�ضj�1S�Q�0��{��6�db���g1ʷpu*��T٦,f#F_������}K���4�mX�aLT�I�轔-0��G�0�g����aLT��5v����cCU�N똱������)z����s���Ԧ������8wti�_sݻ��Ԯ�W"�OnLn�9�)���g�j�yS����� q��� Y�G�7�*�դ?�.�{R@��T�\�-�`8�;���F(�b����{V�lT�'������`������b�ldb�A�(�q��洌a��F
a"�z����c0�S�gl�Kۚ�C�G�1���@�HAXE#���AL�Ln	s��r�v��k�L���~~?��W.���alT�I��y��F��a��?}�kFc�20�##�;~�wl1�a7{;���k[�6��ũG.}�-��S=�Q�8���w��1����Wco��*���f1F`�����V�<b�)��s���vo�֨�;]3�9���IB�#0�9�s{F0�c�20�#Pgo�1S
k�#
���}��n�w�f��֋aњa"���l�%�/x�m����Z�#���SG޾wQ�k��F(�21FvsO��}=�r���l)��S5����sZF0�*aXP�	
G��wQ�<h�#���p��U�Oh�1���7�̫�׵����0��j0�A��=o>֌���S��4C��=��0q�h��#3�}��������T�5��G�g5�c0db���9�U���WN��1c0dh��9��<b�D�a%
3�wz/eL%�ݿkGu7w{��t^a�ƈ�8{ﹽ�S1�aF����{Q�5�F����L��oE���0��z����.��]WN�oe����[AwTgy�v��q�Z��o��w��*/;!�O'ڳ�M������˼��f%���뇚��8�������ܶnк��I;%������N>\h�\>{`��
��8��[����s\��]�Ӆn��kv4��+lYmӏ����N;q����mք��v�a�b�d�����p6�.�m��]���^ۈ�}��gp��}�]�N�xE��z�s�z+����zn9�]�y�mk�
����ɵVNz���{L�ᭀ��jK۶�@n���\vr��8�[2�܍�::���L�B;';޿"FQ�T��Ko��N0��ߵ�m�1d��RPF����G�cpj1FD��=w��[�c#j��߹^~z�\�X�ո�Ͻ�#d�F�L*R9�s��1��Gi���
�丬���[3�wz-�0�?Y��~��D�R�s���?�{0~�aD��0���4C�k��a�T��1d��>ދb��b��r��'+���ԕ�V��ִ���#fWޒ�S���W.�m�3;���x��1FP�9'��{T-0�Th�#�N��5c��Rw_#�Φ�dL#����j0Ʊ5F�Q�a�����[�i�h��~�V��q��0�F0�ٿ���f��vo��d��RPF���5�Qƣddb��N�E�[621F��j'��kH�s;{:})�8,aYB�$)��F�4F�s��U\ 섫���c10����f�a�F��a>�5���a���[�ː�骺׉�l4�L�#D�k�n0ƌa#�#�z�w�ط��NQ�8G�{��1���$���o��ד|��Hݶ5�L�;�(�w8��6�mr=.�v�P1�[b![��7��؜�������g�3��j0�5��(��I��+a[(Q�ph�#���oh��aFC����>�}��0�hg�������5��aA�����f�F��s�
�UөVJ�{�1��#�����0�T�R�F���Y��}]�J����E�}�l�P;:M���U����D����641��V�л�����5V^7��;4_"穩��Y�zׂ�%����Mcq��#d�߷�ح�L�Q��j>��֑�)��VP�	�|���Mk�̶^�.����~�ic��F�sz}5�Y!Z�[�,alT����|�L#0���a��5���aF��SC�>ϯ7�m���r�ٙ���*aMq�b�����[֨#8��Q�?s�֑�`21FL�vJʪ��R�H��cf24{5�j5���9]�s�
b��(����[��У�Da>繽�S0aF*aMA����Fֲ�;�����a�*aL1����[���9o�Z�JƯx�m8�>��փ0�QJ���z��G��b�v���w��\�uc����3Rs��l�21F��Q���~洌aLT°T(�@�{��ucƈ�=}��א�����|רH���}eW�cN�&�����%DQȅ�S�D�#��QJk���
(�QB�_�Q����|�l�a���SPj0���5�m�0���aF��k��a��a/��w���i�r��h��A����S���if21FC��7�Q"��1i����?\ޣ��lQ�1S
�j��O�7o���L�b��a��9�w��1�3�dC�5�k��a�`�a�F�v<Ik���"��`��?6xUYWN�Y*��0ƌa�ﵠǌ#���4{��j<�(�j1FG�G��%����9�Kif��ajA�y�������e!vI��ǝ+-X����-�Q��lЁ�e�nn?���.�i�ٱ��5b�D�y��֑�0�(¥
0�R;�s��1�Da���e���U��w�cf0����e�:����WN0��Q�b��ｭ#l)��#0��}����р����J'��Ѧ.s�;��1S�F(�j=f}�#��Q�'{%eU]۩u$w{1�3F�f��F�1F�L$�FW'�ѭ�-0���پ�_{��u�6&��>�>֑��aF*aMFs��cX�a�F�=>ލ1[
h�aW���߽������h�PjR�ܛ&2�8�ڝ�&����u��nۥ�e9v�E۔A�7�}�-\%7de��4��G��u�m�1a(#	A>��6�OQ�2&F(���z4�l)���;���Vg~�����{5�c�( P�	#�k��a���99�F���Sr�h�1��FM��3i��F�Q�k�;��_j��۳�1���h�X�0��#0����;�a�����L�O��L[�u����
���b$�_���{;�1kK�l���{9YN��RN��1c
h���V��Q��aLT����keL$�F��G��eI�_=��̙�:��a�a���s���5F�Q�aFOO��L63L#�s�1�V��R�4����iG{��h/��7���uu+���g����(#����ռ�(�Q�0�*d'/����c#j8�����5�c
��/��(�s6��������jG�={���a���V+*�+n��|�Djn&�w�n7;��՘&Ξ�P�
�S0����ڶ}M�s4��e�rܫe��h��FN�f�3c0�F��L)����X�rf��۝�_a�L�#D5z���р��a��鯴i�z��T�j1G��=��f�(��/2��NC5��սO�0+PR� �N RIqG=���u�oU��,l�p���d�xm���7�I��T��u�3̍��umc�(�N1FJerk��B�	
aM�s��i���0�w������}�c��y��e�9�a�`�a���0�#'f��L63L#D����]��2��4у�#�o�Oc%bވw{�[Gg��[�S
b�c#d'/_l���*k`�j8��e�`e
0�P���e}��������V�6�׾��ݸ]Jn\�m�l)���-�I�iR���wh�l�2�	����6s6��8��_�����G��0�RQ;5�b٪�N&�q���e��1�3��V��շ%��*h�ك#F���[S�u�T�����G�Hk�'{���Z�����b ?���O~]V���:���v��*�'i'E��A�$�b	��`ߦa��=�-��w���q���X�z���������]�!mj��j��#�(�6Qw���{�F2�;1c�����ŏյ����3�'^��N�畷 ̏ s���H<�pr�ܲo.�ne5��������5�zUDV�k��4FȜ$��`l�X��\���v5ͼa.q̯nM��6�gv}m��Q�YR�ZIv���s	���,ڽ�C����<vug\G�u��t�#��� un�8����)�w��Q�tP#��*��c�L��2ղn���N�iS�랺?ύݺ��+��Ľ���p�$��ݵ��t.਴�\�	غ�s����=��s�i� Tn��;%p�k��ݯ��4<k���6� ���>7��N.v޷cV�)������8��V;uMv�ރ��\X  �g�c�SBҕw���`�j�n���n,��8Gn�G�w�0Xc׻���y���A ���x�t��4�~���4��E�;i}wC����Q���̺x������ ^���>U��d�ֲ���׮� m���f7�=���qR![$F`h����Um����߮� rs}���7���oM܁���h�_��`:��K��]^9sOf�` ������V��k~��>�{�ǈ\�ߦ`;��kӜ�ܞ�a�x�j-�(CQ@V����>z]����&M��^ *�#N�-׶o����>�[������q`$���1` ��q}w������
Z���`��=�M74��U���Ec�W���R5�{Q�AYgn!K=���u�쳌�����#���6�v�Ԃ���;ޥR��V���N����B�"	{��ک+WZ���]��ƴK��>s���� �r� ρ�}w���o����IK�=3ޙ�m��˪"���׶�ׅ���w��n ��e�����Q��>g2�lո�۬�Ow��,��ω �H�[��A�g�����<A�>%�{x	_�X*�*�A+����,�G<��ES�<�6��	����$������;<�~#�ƎG��O����}6�ZV�d���n����k��]����/]n6��Ȇ{W�����b Xݓ7���C��t����^��hMEV����*�m�gp����Җ�#,M'O}4%hY#�u�z�׉y��ψ?{��F�e,5cL�_����WF��+)n����I�#� �6!������T{��]8���uY7r����8X�69Gk��l��nnIî(�U�V���Q����WCv����.E�7I�ݎ���$��7,�/ka��n�� �͡���}/�{�C��[���GL�4�=���x*.�9�e�ɛ��O�״��]��H��-ߏ��n���a�;}�vN���ꒆ H���I$�F����˕�ħ���5��ǛU�l�p9�`�����Ɍ�Շ1�3�1�T�T�8_gW=v�"�Dy���Y$��$}��{���S��L�ƭ`%j,�V��n���\�A�.�7@���
R�U�z5�yv��U�{�h�A��`#�5���_{��pY�|�MiKD���=��}��׻�]%N�3��Z{���[� Oc{��=��P�Fd�le�tp�L/_H�AM��L� ם7OĂO��X	$�L�
���G��EB���S�v�>G�o�����O�a`�u�|�$�|^x�&�5���3rJܲ$�'w�L*�x�-�������g�M���7�ҁ\��\�4���U��vsZ�%���&Ը���6(|=��P�A��*���%�R{�~�^8�k7Vh�ٌ�C5�;���&�<o8�������h�tlGe�v����t��X�(Y
xɝ�H?9�o�e`>V=�`/S� �H>�yg�zi�,�VI���7��.��:�Lzؠ ��OB�~�J����-ҡ�r{ف�5+���2��ʼ�<�������r�U�bA��z����o�_4�x�7���R��0�,O��Ͷn:��~��X	$�w2��O���h�;��{��E( �x�*����c(�#���Z���������|�4��vP��x�@|/�VP��z���}�n��!y�~5�.����42;�.q4���fvt��v�ɜ���Ү���t��wl>]9����,ֱ��)����w><8;�
ŜľV�I���0+��S�</V�Q��vm����:�;w]'wso���r�ۧ�Ү�U*U[-c ;We:y�v6s�St�&�-\w8�;�wd�tR�m)��n�k}��0�U\Xݸ���NX^��WkK>�)��֗Y�^�u}Ϯ�u�pu�ΔC�Ct����'�.�7س��Liv�%X:�ޚ[�����+�uC�a|�{��:�5f�ng$:�pܭ����M*��6���#��c���aYE}je4�ζ�x��%��1�Yb����v�`��g����ƚ��"�Q��t��s�=�ܕՖv�e��BY�A\���;��"��g֞n�Yu����j;�����O�������ZS��;8f�rJ
��/U4�"��U������mh���i^끨�v��}�*�)��/s�6�4%@S���:\`�WZ�T0��m�H�����v,���;��Y�3�Žm��/�R��x�m-غE��zu��e��U�n�e�Pl��H>|ɚ�}yB�P���6!+���aW4Z��u�wma�����R�&;z1v�ۍk���$ظ���Զ^�5�u�������A���f�#:����۫s��:���j֮i�/�V8�n��>D��R�j)�e>�ϋ�J���%����Y�������Q_Mv��m@sG����纫v�^��>@�>�ɶG>�-��綗��,k(��ִ�kw[�g��{ڼ�F�u��<�ӏl�7Zq��h6��;2��f3^��g7��@ݮ�b�$��ݥ���W�iOm�Y@�ͺKc�m��f��^���[������!p�v�GgY����7�J��ɶ��<��׽�Me�-2ݶ�7�����2(�8��e[�f͂ٱd'l�;3��6݅m���YGYbE�k+#H����Km�H�m��]5��$�[�(�����vnV���׷m���ݵgi�v��Q�PS7�Kmn�ޔw����rkM�5����{a��넮���	�{�!�z�SD��vvĻ�s�1ʕ��4=[r��ܝ!��6|)��w4�ؖۛ�Ta�����J�N62k��ϊm��K�9L�m�f��_[X�
�k�u�΍�m=�3���qs�oX��{\n4n��s����/7)[���Ǥ�|G;��5��,�u�fH��kI�\mk�;$Ë��5؟<&y���;�s�����u�WU��8���n��3���IĔ�������]�S4�h�0O`�ݣl���9��x�%��q�;�n���'�kX,���*��/��ő⬑���+Z�r��kY.w��'���n��|pR=�����vx��s�\�-ƧIWfz�ş1Xz�c\JS�MF#�aֵ��OG���5��/C\q��O<����&_Om�ul<����-l�U�օ�LrZ=�;]��h�ޱ��e{v˱�Z�d˧=���?��=�I���d��ݎ瓸����`v�nɣ��1����ƎA����[\!�mv׋���,��;NrS��M���〳�»��*��	���m�Tf���v[��m���ذ����v��x�vr�=�2=��b�Z��%���K�9緜k���=8c�|���7���VQ�v:�7Y�س���v�fquֱGltX1v�ݮ�8�	�;k�[5۔,��zB�PX�n�솯V��pjM�&NӮ��F�����ێ5��ζ�cvg�8���Ns���{U��ۀ��Ry��MI7Sg�=��P�m��c[��흩�&��F�ۙ�|e�1��6��^Mn��͞��N���m�r�v������r�1GYu�{��wo'�����E����:��	��tp��P2����}W�vy��9�v����]��X�ݵ��%��-�ึ�GVW�-�֮91�;��ziMkv�l�u�g�s��!7b�ۗ��!�74��@;��2ۛj4v�KmOOm���j$C\�2/n�s�g����/�5�����N=�����^݇p���vf�]b��T=�+ػm3�h�&�u���e��R�n3e�M��Y�hч�k�팕H�r�a�d։�[=V�k���F�l�^���X���F�\�n^�ۍ�a�u�(�q�'��&��# Ѥ7������8Η�h����N�q�����oA3dz��L�	��gV���Ŝ�9�O�<��;�q��)�+�]����������FX:f��氐	 Χ�`�D�k�%�~��z5���2����N�%�y�іs/ �Y��cI�w�m��ZY�$�_�:�H$N�=Y���!�:��8-��څd���F���O|��,���D����\��,�����r�Q�N��S�/8eg��צ�i�,fӘ,�D��I �tR���o��-���i3fa���М����W�����H$��Xk��j;�E��(s�A���@3���c^90�����x�����DYj�RQ3��Q/Nq�������$��"�������~~Ca��3|��}�DA�]7H$�=�`9�������*�g��{�,���ࣇ��O,^��o���p�w�QMܑ�h�	�U�+�eX��ܖ��wqDfTX�vV�Jl�`wR��W�%��]Ps���96�T����ă�.�7�A��,d����>^S�@ǜʥwVMYB�Z"{�H??tC�%�}^�rݯA�Is:f��&{��u�Ԫ�B���7�ټ�����[����'��A �\�,'�;�{�=Si�yWI���dlv���E�]咘\�_ *{�_~��]�x�=T����ӊ�{�ut�ʇ8wD:�XZ
�t��W\gr�ۋVq��!/�ԧҰ���(�����NV]
�j����4i�������$��*@m/3~I��ܑ��������cl�8[�
�i[��!=w�� �N�	��ޘ�M�R�c#����ޞ��ߛ��p�T�kVYb�r�TMEP)/�]<�Ѹ
�v=���AB�N�檨.�)7��s�E�V�z��	H��i�*�]=�|q#�;2b-{�*I�e�n�K�K�[���,��~���]�wVX4EǓװ}V�yz�}s=� �#(IL���}ݾ�V7DyC��^�=�eX�Wdݑy�1P���	��<�=����
�2���EU
 WI�����y�9�w~��MN}h0l�XϜ�vX�d�^��ݸ^|
�K��c�<�������똅U�\z��ذ'�ϷA[�K��4a����蠻Y�� =��>�Br�H �,�9��1���k)�50�^�"����ԩP�퉀�φW����;�ڣh�T��Y�r��>ѧ�A��DB2���`'�Ň�'=��<|��Z�l�O��Yy�(yY�`TG����=��� ��/V<��G��ٯ�z���Ta���	�\�MZ�u�AZS������P��ju*4����0��)�X�/�,'�
���5eB��x��H!�υ7c��k=�+�K�C��lo��{��{Ҏ�~/f��+#d���l�϶�x6��n82k��j�����dv�TR���DBV�٫�7��ZI�hI${��K˙�r�n, �C~}��?���u��U-���ٻ��Lཛྷŧ�S؞e?j&| �}�� ��J�z:��~�/2�w����Q��I��uU{��
�>�i8އ�R��٣A �tXM^ѵF�6�]+Z3�V+>�au��H*䙿D�E���<Q�^�Q{�����(�c=��0.�T���l��H#cŀ�Ƕi���s�?y?y�o���q*�����p�߮�m�2
�;�����q��mC����r��]m�2��9<�'�=�v����)����ubռY�Y;�(S9[o-�@v}h94훫>}y��pdw\1�np����.m �8~Vy��]:�T�vC�ڌFcqo]qv,tR�Z�K�B�n9��U:�ìe���M�}��f�h�oi�]D�uy|��.��c��z�n׆�-���=���2��є��U7���ٌ�E�<n ����x=��f+%{o ���ص��9Ɣ�����ۡx��4���c������v츹����z@Jw���xZ8�����O�
���7aB��ص��O�9�gĂI�kE3�i�^+�绷I ������0��G9�ɽG�Y�������i�{���H>n����Һ�<���F�!VVj�,�ܩ�x'�^��W�6��=���"��lm6e}�M1��94�)�ɢ�[��AQW���{����uZ!���gu�B����
������z�Kx�3W�bo�!x�ila��Y������<3o��*����P~�%�] >��ט��s��h�b�ըu@��#6�.��\�lu�n�E�uWX�T�%C9M���x-
�e]"��ַx	$�w�Dg{�t}�fk�eꙢR��$}�� ����a������Ŋ��n��g��Iw������x��>������k���W�g���:�N�n���sm΢U�WΆ��۲]���I{�|Oĉ���c���i�=��Kȷ���Am�E~��x�p��(M�� ��3lY�t���y�Ϗ�y�n����EI
B�,��w�0u{ۻ2� ��� 
���� ���-�*�^F���P=1U�U҈����1��~}�M=�KLz7�۠t�cC?{����@�{e�$v��> ����#���uG��4Ь�ժ�*�c9�y8ެTQU
��XT壻����eUJ�
��P��?'v&W�^|u�����]�������ovI��	c����{�_
4}OR �����s�: �wn�eg��#ë%���!���E�]]Y�����A���Ag=,`�a�`�H��Ø��WxW�[��Ը��iB����w�W���z�{�����Vz��3�k�KB	pwm�U�kts���`ۗ��̳5�H/t�uS4xOӹ��|�}5��'�����@�ӝ���^�k<os� ����'��^|~�h��~��Ưi ���Q����,�Q���F�{�a ��Xi���H�l���Oγ޼��A�x�ת��G��۞ھ{��� s��\�nS�!�����q�����2vvV1��K_9u�����n�1X��̍�9=y�$�����~}<�Vo{t9=`��ѥE-����5@	>�vl�W�TK�p ����>o~<���	ɱҙ����wvM���Wg�3�Ͷ���m��o��약^���ծ^|I'���O�'p+��7V?^�>��%�+`����3�� �$��	�1���{��cB�<p�ј	�G���oot6!�T�E̊砫vF.��05�kd��3+�K�i���i�bgמ��/1G�B���~.vi��O���/�!4�wH
 E���~�����g |=���c�n�BO8Ud�A+�IF�V�9n�e�#� �p�uQ�q��k�q�P�a�<�q_�����Y5xI��"<�P��F��^{���=��86�ֺ�}ۈ �EU�m�B�%#F���~�`�r�A�8Z~�Zw�I��������v�#��#�����h�ͺuU�Rf'�ܰ��v�$�C7�>��r��� ����M4߳��bo�������Ps�_��y�A|��o�� ��Ѱ �^���w��ִ�'±(
L�4�Vn�$~��ǌ+��V�Ur�O	q'��3�I��v�Ēb�Xm̷�o��	k��1�L��67��h�5����8��t�2��������S�w�k��i�\r]�n��5m�"?g:�n]� q��\�F�M�$���[�\K����9^��X;=cCc6k�gq��SY��;v^�����Ws��v'��jq�{k�N:�w�4��d�\=�����u��ă�r5ɶ��fy=l#ڸF��K����Vx�[���v�|u���Vݠ��v�^��sZu���հ�/�;����P�Z��g�/��;��>1���ڍ� ���/�
ݺ"�+�{��!����wl����GREY�]wg� ����}��g����K�@ #ލ�> x��N&le���f����$v�ۦ�۾EJ��0�a�B�n�TDAe���D�k�ݺMw��=���I�kVeG��P�D�j��U~���G���HG�Ӱ�o�b����T� q���t�QB�I�Ӿ�3����,�K����OůE�%��؍p\���i"�����̻G	À��r������P�N��ߏ�N��
�Z��
����ŇՍb��r��T�	�Fꫲ���n�$�L=�	���B�'Qi��C��8"���J��ػ�������x��^~$�`�{�ʭÙ�^����F�GVIy�'|5��:_�Bk�뛺m7�[@�g��Qn�ƫ�u���ݪ�:��,ҩ�O'֭��,dT�����,�y��;��̳{I��ǽ������zvpŚ��I��Y�y� ���a���>s^��:�j��&묮�,��b��u��ޘ��I&��t���!$����~$�LY�7���B�%�*�w��>���Oo@����H0��� ���}����{=w�iu�Q�T�=贋��l,%hU�~k ����Ѡ�;�-n�޼/P �E
 W��7A�hE���6?�v6zm�Sg�|�6�x��������Wc>��i)p�\_Ϲ�>�2V���'e!]9@z��-�ދ��Y{& (
y��o�]^ef`$}�����.��kU�r�׋��?��A�k~n���a�Q;=��(?X�f�&�e�^!��T ����L
�}9�[����[y]� ���Ʈ���&!Ҋ|XN�^!h��v���U���$޴�`�f����솄��*�v�j�z����aN��+�6a_#�s��N�����4$�n�L��
�
F�lJ�7wq�t��wJ�J��ZVZ�\�N��L�9�_=4�&�X�j�;�v3��.or�ɮV�sܽ�f��Ci���=PKc�b]�1B�]�+�j��\��nŊ��z�L�=�V�<4�W]j3K��9��(��>�^�NV����Zwj��`��հK:n�ْ���x�1R����A;�j�����wYMa�r�&]p:�<�����>5ڰ'h��(T�"Z*�sg/G����cyV��穓|�1�K:o"�w�X���H�7�5�pp]����5���x�:�&=d�u\]g���c�릻�P3y�)pDr�[�n��e�J�;U����˹:�mt�F`ώ�m^��lS�����ArQ��Q��O�P9ݣv��rM��`�4+IGM)�7��KF�&�4te�9]�'�gI32�Z��,:-r��ےu�+��cq}�k��b7�zmf��Y �s���̥MWG3:��*���K7�r����q=Ka��&����_5gE�,0�x�FT��^O��G�㚁�u���-�)�HX�OJ;U>u�;��N��er�T���_˦���r��/gF�s�m8Y��r���lj�m��4p�L����ա�2��K8p�A٪h�TEU$�I$���mFۧmIі�I2N��|��n�����3mYi!Y���C6�m����vlݶ[��g:�F�dn3-����9�Fۍ���-k�����ͻ�[,�IAmi�X��M�ͬێ]�v�vv��3���f�ݶ�u���[Q�g6Y����j��Ee��-h����������mi�-a�q�inw�{n�4�i�k���Vv�3Du��ɵv	�Z��6���u��f�Z,�i���Q�ٶh�=��ݛf�ɶ��h�iim���j&�6��m9#-q@۬Ͷ�XY�Km��a���/{5�n��Mٵ��i�t6���R�k�y�Ѷ��y��c�����U� � ��	�A��/A���{�Y�EIv>�$D���WB��X�'=�X	�ۈа�D�UZ��o�{�������]M�r,�*T G� p^�B���-��C���_�J=���*Kqэ���;-p�Cv..�`z%���[��z�����KY��&(���O� ����0Կ[`l�����g��띚3��7G�Jʺ	^�}���+�h��g��)����H�^�v�$��g�� �^�,>{s9���a�M��g�'"�;_�1>�k�����K�~$�y��B֣�����O�ޝ�b�vi6��^ʓ�� 8E��������N�H4�{F����,a'����,j�E�>4�Y�.Eazi;�p]�2ƚ��(wjL�s�F�d��������h�J�M:�X��N�C��gs���rA��e{�o��9.��B��4R
�w+'Xω�b�NG3�� �d�� �}!]��k��nl�Z��J����pV�8"�YwN�)Ϯ9��\v%u�z:�2�
�z��������uřz���0 ��J��v�J�S6'P/Z�t��7@|Z�b�,��,a�f��H� ��X	�?k�ɯ}$�l�O��$�}, �_xk��ڽ^�Ή�mN�YIc�V�t��>��=�U�����|�5�� ���/	�}&,��&�]�H�{��5�خ�72��#��I2{0a �{��洑���W�(���oϿ{*N�T���n�6�O|������ʟz�x� ({��({[��Pyy��pQ�j�m�+�a*���ovb[�T�TSyY��]�e��׻"�՞���,=h�Hu��$���Tߒ��B���q�xr��V��
�Q��ۄ�{;��B��{Z��W��Yz�p9�3�d6}:������G!��a�U�Q-�m�&�װ���]g<��ǩ�cn�ݐg�:���:vNx.zu�hv5u�Z�m���k,���p
�j��h�.��v۠3�E�MGm�s�a��n0�X�)��u�\�q�I�w8�vx��j5���n"�v�q��l��0GKÆ��ݰ��-�M��e�l������[�u����͹重�jSZzˊ�*�"Ѻ�EM��H-�hP�k~leg��%�=�J�{ ����$�v��$X@��w�o��d��`N�+	T*o&	$���	$y��F�qzzv,W�ۭ��,��7Jͫ ����k�(P���	�ͦ�V߯Q���WI4�^�g����fB��V
�C�<}�*`2��7^�@�w7�L	��3|��L�7�倐��^��we!�:�k�����5w�5���*��I��^�$�7�`:f���<�)/���]�v�Jݮ6���)��1�}pw=� �^�vvr&�!���Q�E)�|�ީ:��1�{�oZω$��t�I��!4Z`Н���+�z|eȰI�D�^������c �{����Ƒ��q|�?Jy}���'8���]�v$��J�H"fV4��t�|P2���f�a�8�E��� &.{L���)��6/+y&*���>��k�� +�|i|.ws�읎{w�rs��aJ�N�ɯ�Nrω��d�a ���6p�^�I�@
�+�+��]�pP$ж�}��ޱ�U}�0�fL�H$��XHOk0c�V]*�䖤GY�-e�9��T��	��ڰ%�<ߧe�ʘ���0z�K�?����%��~�_��2�[�"�Ö6�t���u;��#��^)kN�T�.��#���������3�$3�/w� �)YK�2�[n�_fkZLyZ�M&�o��@v]�9SC��-ze��~Yt���Ljn *�<ʡB���{%��*SMج���H˶կL���Ȫ  �=�ܯ�N�x��q��24�^���\�mE{Ov��
�x/�~�.8��:�OS��ץf�O���w�5��X�b
�/��S��<n޿~&V{�0�;ذ����1T�,�w�޹�"�[���^���O�~��	�s��^��>��gСEM(
������
��WB'�nf1�����������ʀ�o�B�֫�{�l�m�r�.�+��g�Oekq�� *�c%MQYR��EN�T1���6�!�h�uZ+g�3��M�߹@@WO4�IJ��'ssB��u>�5���ω^\*j�]YH�{��_ y���M
�s�P\��>�y*���*\�������(A�\��'yW�_
o�T cӥDs�F]���  �y(|�� >�Ct�l�����[g���|<�( >�2�
�>�����֍�CƄN�Q�%ͬK��B:�˥|�:e�5(���u��V��j�5ټT��oް}�z�^Aw�C/���7j�P@Ø�����C��"f�s8��<���ɫ�k��Kv���7��v��*�^��|����X����3Ë��l�v�Q��Ob�F�#���XX�;jf�'��.|OĀc��ă=��2����M �� ����e�]�F�Q���_
^��~�!�W^8��P�
���O�{������+��ŀ��p���ue#��bk	!�ZI�<���{}w��Я�0H'��gĒg����|z��
���8M9��de�5�}�~���h�H$��0�y��7!�w����3W���o�A�n��(
 {y<�jͿ%K>@TO>��` ��<X�j��-h�ɬ'�=�#&N��G[`��	N�V�a�%a��<���Wm�@�%u��bm��pɮ����v����1�|�A��$�]��5p[96wZ��^��n:.2i��UD:x�2�lqq���i�{W��a�ٰ���p�\�{s�6-���Oqj��vq�희��3�O8�p�I����@�[K��ltV�<p����m�x8�tnЍ���qp����Y�z�G:�/�^�ɏX��>y�M��N-m�5:��4��F�W^�ðb�݋�k�]���u�z� s�Rm�x��;���pH�h^ݘ^��ҫ���ж���K_;�o|�~NJ U:K'�T�� �|��	$O<��}��S՚�_���&�_����-��`�_�5��Ƴ�A�x��9Ӕ��{�@5�C�{QB��*�z���fa��ٗyv�]]$Q����0����j�����N�n& ���(�����rv��7VR?^��&�L"���~�<P ��4��=�j�d����Ծ��92,��2��?!IQ�F���o, � ��Y6�F:�����)� �,�����?n`.u{M\�NV{�\���v[�)Y��v헺_ǗlӼ���������tN��;s7��V�*���ߞ���1@P��P�=�e����;�����$�1�0]Z�h�J�W�?r�}_M��{S�߻�]x�ܱOH���e�7E��V��NN|
5$�s��(�0�q�`Yp���y۷>8�Vo� U���׈$��`�O������=27+�	}�r��n{4�]i_�6��$ж����(���Wj�yS%�\Q?���|���6ɧ�J����6U�>q��}B�}��E\�����	>��-_��,�	熘F��՛@^�+o	 �����>'ד���H$v����B/�w
�V(�p<��8���������9ח����(./B���>���V\�(�*u��ޚϾޖ�cO��������*ǹ�oȯ� +}�R:�jI =i�]��΁ޭo�3�މ�S��(P�~4�E�/rK��1�	8h�wj���Uj�|W��0�H��P@|	�O?cQ�����Z���U�Z�Iǘ)�5[7o�RȻ$���M���I��a�U�1L�~���A��Bk�!�UfU,�ckO��%PY��i1�K�eP P�~(�W����~��^�Zc�SS�����LI$=k  {a���
٪��t�@G�\G07H"���>�k �NY���8�WQ�	��fa �\ְ	>��%�>��~�'��A��8�ut�NiiJ�ᶛ�m�A�x�mi��:ۛQԇ4`N�}��}7�B���YުH +c� ��l_+a�c���w��>�gkXI�,�+�F�Q���Ƹ��k�wvz��$�|�����N@��*H�Y�w���j�F���$݄�o��� Ot*��
��~�VL��`k�T
��c�:U��(�_R�K>8�Ҷ��^ḉ"�bH�9��/���Y;��<-T�����;&NT �O ���'S�y�y\�JɼM�X�f*F�ƝP��k�i�g��7[o�/V{o֨�&�Ԓ�'90O��|�`̾�,���L�I�X�	>�r�A'�=�x���>\��7��Ig0���K֡�u��� 8{s��g��ι�<��\_��x�~�]��?x�6��$��|O��#�f3��r���U3��a�氂g��g�熠WWwuf��ɤ�<�U����o��$<I:��0�G�{0�z�߃�zp��L��T���F��xbְI�ϰ�I.�̒f{'�ȅ��$=�MY�{0���n�FY��I��^!j�i��N�	��� E�U���+Րy���y����j[ۦ��-G-���YE�&�0��� ����*��ψ#�{0O�g��`޾�Ğ�e-so�����۬���{�댝MP�Yp�r��a�U�MΤb�/�s�J�s��Dl��w2�Sb=�:�.R_f
�z�x6܆Zk	��-�E���
��^��@.-oI�T��n����	+`���{>��}�cH݄EZ8xR��=���gd����ZZiJ�sT&?�2tB숟nh{!�/Q�����ʈ7/*<H�*��V�r��u\��V)�R�(�CG�X	os;g1���YUu��4�%���]f��`q^�k��JYq��y`��66��t'vsߍ�l:�������2RP�23v(ZM���=�1ZIb�b��,�U}�V��y�ԩ�譆�i����#�髲b�e��
U�Dv���W9�]�m��J�K� G<y�^F����f�WX�⊡��̬��1ѭ�nժu���جayoK�V��0�r��&�V���)r/,0n�X��\W�v�gW
�9Z���n�'�1ۂ�|Tz�(����N����Ov8:�V��otk"�:��s3x������u�.9��\�N2]
���:>8�6s(TKq�|���;��Cm;�W����RmfSuی���TL��}�ڠV��k�R�l�v���ze ��l5�7�Q�z��Q�
�r0{�1�n��247�9ޞ%�⩏oq�"Qx"�Q]u��U�c"EK$T�u�(�כ����f���0�3!�n��\��L�q��Z�GXr-�1�f���ݼӌ�Q6��[ieR�����S��.��KѠ	�[�;��vΕci��ޕV-0��o>�6�ٶ�����fv�sm�h�km��vԖ�����Z�hu��5�8��k1+vq��"��)�����f�֡m�N��v��g"Z��J_+'�v�5�ۑm�l�f�vջZ�۶�l���!������֭�,��sn���l-&�Y��1��&ݶ��l8��&�֜���Ml�r�`YM�׷oh�[�gL�6�d	�Y����Hr�&6��M�Y7c,vm��8孉�Ֆ�r�96�93F�,��٤��''2�"�8�9��R�Ӷ�Cn�f��)�e����{n��e�Y۴��I
�kS7w2�-khN�c�˳�M�l�e$Zu���6қV��GVKݔ۫ �V �Gge�E����vu�mn�km���6�VۛdT���[d��8��mDY��s��!�[k3��w�����n���7N�Z�Dzܹ{3̰�x#�O����x��n���TF���s���s�a�N�ɔ7<scٹŅ}W]p���	n^���r�=]b�v�����I�Z3��K0��'*q]�����bxqr��Ʈ9�z��;d#=�������.�]�닖�rqq��8�%�/����dG�&&蠅X8(�H�m�=ۤ�Ge��'� ��sg��g��1�>M���r۶�s[h.zM���㛍��s��z۶�oA�qn�w=���=rj��v�գ�{s��ꋝ�N-�@lu�'��i���3�n����Q�˳��I+�G]���b�s��A��u�no*q��#�q�������D|����Q�9���goc���� \2�֯t��N�ŅN���y���XF۞lq;�ٓ��Om���+v��6�1u�n�M�wK۶G,��'[I�/K��i���Jg�\��pg��ޢŵ����ٶ-x1rb^y�īt�'M�������q��g���"��q��۸ͺc�ӓ���׎&4{q�6;[l�8�r���8H�ݱ���ݬz��q:}v�]J=O*6nT,��m������;˝j�c�t���U��F�����R�T;vxwW��F
����T�m��f��	�0뭵�o<#���/cm���Jv٢�4y��.3�S����v���smր����-��-�m��^�j݃4�M���:�㳸!�2.ۗ�_&Tn�7O.Ƈv�u�Srm�k�]��������Ÿk�����V��V�'n�{8��v�e�<���#��= /�v�g�:\z�l�n#vfy�\Ն�Aq�{ ��ے�^n���v�秞Mnt�䝮Mg���O-ݫiW0Tslf��g�;�^��[��v5������v=d��k���]r��vu����'b�t��j�Jp�n�����6��q� �i�n��4h�O8뺭�x܍Uq;��*yJ�'��˃g<;�6�:�	����OB�p	l�D�q�q�cq��tv���ӴM�uny�s���I���wg��k�Os<N�dt��x6F�ݹr��v���ǋ����=��g/.��we�w(��x��:���GZ��ͮ�M��W��Z��N)���1mv��s�q��v�7�۳�uΊ�|�wV{8;uq���,GY�:$lvv��g������g'�rQg5\P�rb�cW����ߍ��k�IY�s�X?|�,$�3�a��'}�[��:(r�+�z�0!VR!]+�|�,��M!W���{p���M�LI�Ȱ�L�40�\l��{�.����a��wwuVm{��y�	 ��k $S{�y{+*��נ�ę���=˦��4ΟX�@�	�뛧�����ٝt�#=٘I$����񞘫�ކ^�l�z���q*�.�x]�d�����,�~=�> ]Љ�t�燾%w���.�B����U�އ)?��ޢA���q�;��r�vyN{�q-۞'��z9go��[9޿/G-���YK竮�K��,��ޙ�	V�l�X�N��9�7u|�ͧ��=N�ܤ ����i_ww�2�v�s=l�qK*��4�At����&�Y�#=Os��V_b�J��Y��6T[�
vvt.Ċݹ��x�+C�$]�9?1� Ը�B�{�@���Ӟ�;o��5X5���e"Ҽ-�XOğI�$ew<���"v���;�	�fE��}�Ș�U���]��A��n�%AVg�{�?6=X	$�߳>�H��h�wFM��H�o.��mq�~��%A��~����m�o۸xz5��Of��xI ��/��-�7�Y�$�$%%��t.�,�P������&�ǷQTj���Y@V�앀��H�y���+�v8[A��5��&��=���m2<���Gp�^�>^�^I�<X	�є�$��+T��=���#U����[���0��7��EQ^v��ّi{*��B_�jf+��&��罚I�̬�^.�R���ѩSPl:�34��&�n�ה˸! �֜JxT��o. e2qd��EQ���vv!l�_c�=c'^��	/�O�~�<�fp���֬,׎o��#��Y�L__lXA��On�Oެ�u�Z�n'��N��}����H�
��O�߷t�@"f5���w]��߭۠H���`�� +�iT+�K�{َ�p�&�Ş<0\ۨ�r]��w�7Wav.����˄�����bݹ�.q�����s���.�M��s���O�ٍa�����1|-�S��$C������������I���R /��zg�/VȒ��	��n�H>�hg��\|f-�3��^&��j�جw��ePK_6>y.( (s�b���o:���{�ﴱ7���ʼi�v��/�ڙ��I�|�.ʱ������KJ��zbNU��$�F�{�=o_m�+gx���zA�8ξB��E�~���ZؼQ�/1������\ǊRLw�S����`p�^�b Ov����7M���<Q�G/�)��o�I6��{��ob�B�1I_��y{Ѻ���GI1�VU�Ӽ�N��['mY���n��z�7,���l�^�dV��7/Ŗ�Gj�E�:����!R7䟹��,i����.�i6��zfr�]%<��0��t�H���mu��J�Z��9�뛺m>f���w�:������ �bư�	3���=M�^���z��x����JŔ��0�um�4�S�#HY��C���� �H-=Y�$��՟~F+�Vg����$���z��)�B�{� �����a�>�����M��J�����$n���y?{ ��J��ePˡ�@P��U
��7Gڵ��ƵU�^����RWn��r���|��:n�z�	��K{Eך�Z�t|J�����e��Yo�P���;���Z���[mh��f�O�ⅎH�pf��޹G�P�ss�v�x{v-v����ۜ����h+�NȘz�zb��荶��Ocv���nZ�GZt3j�[����l	ûu�"s��΃���7h:��}�n�֝��z�nϫ����ă��0;�s�϶�2Ǫ38��]ť��':��w)�|�'�J�I��ձ���^��L���G����g�*
cG�q�cXW�{=n:��&ܷ�ru�Q�r�n��6���>�KU�_R�C�y~$��0�b���|M�K���?g~x��	��`'�V2 �H�O��3>Ÿ�g���=���e�P�D��A�o۠}4{ܶ�WݑD��B�?R���/Mr������X�
��ּ
�Ou�������$�|N�8n������5>�꿉.�ψ"'�n�I �1��YI���x۾̺M�[Ū䢥��9��{2,�\N[�
�����	�4}��5�����NVW��Ї
 :������e�d��������&���ض��u�)\＿~��!~v��~O\�.�$���h?�Ɓw�bs3�٘�Ϛ�n�OۖN�(R��R����XH/G\ug<���+�V�Gq��-����u�3�YkU���c� ���˨��<��"��N��ʴ*�����3M�X-���B�N�P+J [+=/v���k=2�uo��2 �Hן��n���� ���"Z��'�H�7̀��i@u]jl�M���<\1���v�^b�@�m� ��C��b�movL��c�N��wěω̼�yum��4����Ȫ�9�~MT��7���)d�'�A��,7�,�����o�^�:�����J��X��N�w�V�ۧs�1f"v۬�Z���-���Ӻ�|�yOȕ�`�e'�fN�?!Y�	&zf�7��{҃��;tG�c�$MCy*���dh� �cX&�yڽ>�k���7�O� ,��� |;܏ʂ��wH�K�{���M���	�Q�Ɲ)�ߦ�m��A?�!��G����h^�aO#��s�{*�M���Y��X-��3�q����RU�x��;�mh�m��>��:}� �R�c>'��`&ҳV*������m���m��X�j��h�,_��T(WG�o���^e�|l�/	b��#F����6�b�( >=��
��)P��@����G�l?3���B��y(Y"��B˺��:�;�Z�s[z����Ǥ�ָ�R�~~}����Vf,\��y ��60�����gK�I'�����hU���)4�u�bƟ�����g^ٖm�Am�A�ݏ�4>�i�v8nU펨�8M��a� �m�>Ҩ >��6>'�k�̻i{3��@/�,��gc�����u9,iҞ|����G27C<�T &����^獮6�&Sz��樢̩�\��f%��tKB���l����OM����y���i�{��������p��)<1_�*
���}�Cj��[��V���6a*O1���g��g�
�xrR޺h�ֆ�G�wA/�{t�}K]��-��]�}�Ƃ�+�n��g����;�
C����GZ�z�����r+��}�c����<�3�I����z�� �|��7�PC�j|2�&A �����;�l������t��^�,K��੧�i�@Wj�6 <^�*]�':���k-\�{��9Z� t��z����$�G�ŀ�yu��n[�� ���~$�kY�3P�J���}aZ�~����@/����N��|!|U@|;��/�m�;\<	9G�	ݳ�~(U�v��T��y}��LXoS��"U{�����>Ѥ�ń�1g� Iʜ���Ľ��������ݕ�w�دns�l���lrq5s5ssb�P��g,�m�,YՁAd�����}�M�#2)���:�Ĕ� P[�P=�m[�ڻ`fㄣ�f�k�ms��*u�۶��mk���7%�dtq�̬+���M�l�Z8���n����sԽCO��6˲��p�'�����������[s�rhn7tY뮢s9Ŭ�oqU�x�]��u���B�s�R��sh7\��ui0Q�f뮍����;3q�ƹ5��NГ����n']��8��N�ڮ�Q\���]�U���[m-w�h8"����[
�2� g�<��I������g�!�n�<����O6� x�*����P�dX$����C�Vb��*^4�竩��	e�  ���P�:T�R�vߓ^���N��~��%lfg�k��g����h��{�Ӣ�T��IĒ%-��D�ş<m`�DZ�TJF����jc�����4�@
�*@�E�g1}��	T޽�x	�lJ���}aZ�/NL�}�Ѿ��n?p��c�ϯ� ��, ����c�K�|MOtf�>���썊ج���V�GT�I=�J�Ωcn
�"r��Q"-i�S���\��'�zfr-$��쩦�k���,Ja`�Z,�;	/��3/���D٪�@V�z<�i��$�c|9��������XA╆��K��t�+|�����WKƥ�q����ܒjY3��7�q�{�V�[՜b�7�9Wn�.Y�>�>�5*B��0>^P�Or�&�)!U�Fǯ9p$��~�?{Ù��~8�h�B{�_
@W��7�~�笕�j$���Xk��r������~$ݶ��~ْn�O������<�:7�����3�=��t�`�o,�Ѥ���[,#��`�C�s��p�yj� 9w7@}@W����2N��u���p�jL�?�$A-V�[j*pl��f9�'4u��q]�m�~n���y�v�K�������XI'����O��K]��O�T/���|&��a��4�/ �4A���׳� 6��=rz�Q4��N[ɀ<�T 'O�l�^�;Mz��ѯs���T�鞓wI µ�@'�1�?#ݽ��5ep�s�s��6��Rhĳr�>�M�;v��t#ϵ�0Vh4H��5��uVm�v�*�_v��5���b�2�7u���lP�.�k���'^���(uϪQX��u0��<�."�F��+��}��F&).��v�3c�����s�w���`�W�%��yذJ�����<q��)���'{�e�M'w�Mo���U3.�����uņdX���.��Y!�X���C���i��6�[���Ǌ���-�Oj�c[݂��\���Ӻ�te6��y�g 4�[�Z�5OMEX����MC�Ai�;�p�</6�Pg,'5�WwfI�C��l=[|�x��\J�J��z��u�{��!m��-n9��f��[�@=ӮŦ�t��lF���.�aNB��!ix����2�.������	>�qĥi�W`e�O�ǔg[�v��s:��1�����Kc)]N�5N��|r�+ �6`�u�?�������E�z��n�s1rJ��0�y��7/Υ{�xz�E�~Ͱ���]���֫��6XE`��gaI>K"N�ܧ�e��'p9M\��>s2wf;P;���P��������8�uc� 9��Iw�F��N����\*_
q������u��.�{U��5X�z)����w|�\�R�eA`��iW`��+
%�F�ݩ���v�̹,�$����[��\l���;�rdRV�2��b�����K���De�g��r��u�/y<��'��_�����Ow@YCnX����0��*��������߉�4���q%��ZE3f�۰��D�2�ƶt\M�5����2Ӳ�5��\X�sl�1�m#�M����$ҳ�f�1#�8f-�-��kv�ٵ��a`�jK8ʖn3m�DBrB�����m��W�Y����J�m[X 8�nّmd��M��!pt�Gfm��䶴��9�Z6Ӷ�l햠�7"���ݻk:���H#8��f�&k��wYYXVt	dqӡPq�۹F�� 譵f�鰀S7Y���m6�����a8���KK���f�8�;#[q6Ͳ�#4p�6Y0ݷm�)��ԬmmjC�j-B���;ie)4�9;�Y��Y�[���-!�[fX��ݭk2ӑ�v[g9���!�n$B���g"��2KrSn{ޑ=�'(v��m5��Z[Z�"R#�8C[ki�3�ɳ��m��wRiu����4׋��M��.i���ι�뛸�rK��%][�O� �Y{���{܏�7v����\��ck֞���,����l�@U�F�����,O�����3{,z$�Z���6��W��\�y�6.,pv��/�	�=��u8���ȕ���MHB"����u2¸���y'���km6>9��63��Vhor9�*�=d�m"���m|��3�I���-�RK\vJ������6�X�Շ������6�Lw��H>�şL�{o=�ww~�	��� jɫ_$U�=��H$G�  �����r����H$u^��	��,'���F2'IR����/w��있޷�@#�q (wy*@���=�<~ڕr$n�bu�m�G.���
��g��N���$F�k�
��}N�f6��3Q��[�[QΜ1��F�|	����%��*���(�|[�$�{��Cb���Ͱ���	�F��*{Q_ ~$	��l�[���[~�-IF�O�J��/k ����a�]�9{;���k�����/3g�e��RJ���h׷4�k9�U���+�{�Oܲ�Ύ�>,�;܊M���Zl�\DN����4�r�.fҊ�|~��5*U@E�O� w�`[L�G�0�j��7�N]�W��[�+� ����>���\Ƹ� P~�*�}����1�кʼ?b����Ct�n�A�`���7I��ֆ��^��j�ߛd�]7�o�"�@^�3�ɺI!޵��Q�<�گL��.�ϰ��٤��Z�j$���������$�/��bq��*t����G�/]+M�yM9�"і�N��N>�� ��o&�,[�U~��W�<%�ŵ#���'�[�~����W9�AT5;�#v.�S\�2�{U��}�{�F�FS�%�����k/���u��7+˶닪x��5X��6�א��m��Y��m��[Nx�Ѹ�\��c��w%`紷�g�q=�*����Df���um��<S�Nc���/K�{c�ӰLZ '��Ƽ�O�JƦ浗��78㞷"�����p��N�7����qq.�V�xT�����{g�5�lb���$D/�7�rB�DJb��_��I�`y�kZiB)�L
 {�T|�]͊��a��k �����>���,!Z�V�f'���6�b��q�EHey�$��:{t�I����`���o��y-�b�eF�f��{7� �G�E��L����z��A�rn�G�5�ٸ9Z��J�+�*�~8���VW��ZUVEw���Qa?�� �=˕63�O����Ѷ/KH*�ȃ��l�iCӑC�����e��� �ZQ` �?b�x�r�3�S��rr���(ZD
E>�B+cQH���ƀ��krB�8)��Z�	����["-M���7�$��k$���y�үy����w�I-&�D�^��	 h��P�����O�Q�XW��mv_��J�\�~/n�mMq�ND��t��`{+�=��X�9DJ�`�֪u}�&��Ƥe\7g8��:-�A$�nB��G�	}��u�l9�չ�w㙀`#0�v��!_@�EP 6���3�nJ�V��|H�|����O�G�{Ŧ��ʅo}��՟o3.u���� ?jT����������|7ۤ�fin�R���f$��r�6�;�n�a��,���<UB��~UD�鞛�rY^iM8�P�"��xY�y7n��v:E�z9�p^���0��.͎qz���O;yў�M�k�e]�|�A?G����3�w�_S��7��[� ��0g<Xk9�j�����7��װh�\y�����w� �?d$�<�.��R��҄S�"NX �2���98P	�|���,�웹��xO��v?��퉮e��~������0��4\MX��$Rb�kN�q�|�>�qs�B����p��VCf�+�Ȫ>�N���+㙀`#0�v�P�!צ�5d�vk�5Lsk�>�&i$g�����=�^�޻�]&�4��i�F���Z�?��Kϊ�|��k�B��} (���4s��يԮ�Y�Gx�Donm��]���-�a긱s�n8mWGl�^����(�X��������R���i^sw�6�~�n�A�絡��Ty�R�TEA3�aOt�$n��@ص����!��6V�t+��.����}ӟ�/6���'�����X�&��Y�t�#=�Х�J�|0ץ/
]�]e���{������kX	Q/H�E"lR5y���#u��U>�z9�3'7y��	#&�3�I�؇^f3��o�밹$�����>TOs�m��7�M֭�!�A 8����m��;U~�2�t����5+�����Х�;�H[	[T��Q�G�;�{�~�2�����]�Uh��w���b�Ԟ��ڲ}�ZءAG�  ������.��������w�<�>���i�Y;f�xh;j�m�;��_�s1�\5VU�4.��ɛ�4�A��  ����'�}CN���/����&�z�v�6���ܖ��-e�x��.�Ϯ]+�sI���O��` �}J-EU������.�4�_+Uw��q��s�0����U�R>]oz���6/����XO±�$�X�b� �tw���?S|��z���2	/ڗʀ��<����3
�>�@T�^����X�j�n��A?o��j�P��܁׳,~=X	�y�ψ �7��5Q,���̵�c�n>����}�ژ�u,���'��CyR�5זIσ��/�^�Ve��f����M�
���z�ث�X�#�x��_#CV��,Bv�R+Y���"�����nYf謱l����a˵���͸�;,����B���m���g���0���{��\��cc�m�rhvW�2�=��n��|���v �4[���bޚ6��e{�u�p���x��y�2\)�������m{p�䛢D�[.S��Ɲ����ع��O�;��}p�Tg�	����J]U.�w�y9l�2u��f���\z��m JKc�y]�"ʻV����0N�b� $y���6++{d����r�A ��Y��w��P�����?'TZ$.T�hW_,$O�x3�I>o��L[�4���}׹�\m+��9(B�е����$y���I�~.�G����'b��ho��w{lވk%�C�Z�u&���9R9��M���MW���|�f�.�&%yb��P�{�a7��I��8�R�1?{��ķ������||����4~=���}�Wҳ��WL��\u�η�C�M���9;9�gvOU�-�O�׳�HN���TX���:�k������O�����Iӟ�P'�P}�u�n���$�}7~$/{+��ɲڰA�
����S}c�����S:�W�ܒٌ��%�{0r�l�b��$/Ξ^�ب�L�@��C���g�y=]�^%�I�K�T/IB��@P�o�> y>*�Ȝ��I��T5RxX�5a��?G�b�H'��=�d��;ͳLW{ӓ��������*��
Fք�˂�5�p�'���i�O�b�OĘז:۷*��;f?�t~��&�B���]�-��P���:hM'ӷ��E�� '�|�}���{�I��/d�67eo��ĥ�mϗ����������;'5��i������,�En�� Ղl] � y������> ��J����b�t������j|Pz��8��F����C�B�
o����O���>OJ�B�k�L����i��W��݃t�b��ߎ[倐Iּ��H�U	ާ�8����{mY���t�6m���ki>��63͜�:w��QhfV�bQ-�A��ʷx�Ηc8:��=����P��قyE���n��Ήl�I��a?k�	��`�Ud�UX@�)=���'�jnTnu��
xY�@N*B�ޛ<��j��޹� -����e��#�� �t�w���V��p
�9"� o*����'����g�e��)����|)�I=��v⮼��Kn��eݛ�=���4�T��&�N�W�+q���JI���� $��	9��M��\xy���<�|ؚ��~�M٤[��~���!QV\,`�İ��Q�}�Ϊ���+f��G�)�tBA
�X�ڸ�Os�n�@*����a��k���-���g>��^�W�݋"�J�ki�s.5����S�M���ކ4ڧ�<��<�P���_�2�A�l�r�\��⍾�mV H-�k�4[+��xq[+�*+���}�[�!��3p�^*Y	������uZݴ�_6������'�*'jh"��=�g|H#ٱa�b�v�\�x�[� �}�s>m5�gn�����O/O����pi8q�n,޴�z��=���k�Ky�=vu�Hlr^h�e��*YWwT�+Y�|�	>��g���F��,�|�Q�������<�M����PA�Wx�E�nS�����/�I$���ĂA�lX$�%cC�ߨ��r�
���A�$ٴ,�y��O6�U
��@| �;��cUB|^��	#ٱgă��#D$�AU���z���g�v�ԥB��?� W��@ =�=�y<�����`^�~o���d+	X�k���$��_��gse��0�<�� $�ycX	���W����%�"B���B��$�	*�$�Ȅ��%�$�	/��$�Ȅ��%��	!K��$�	/��$�����%�	!J�$�	-�B���$�Ȅ��%��$�	/�!$ I�	!K�IX!$ I��d�Mg��ˈ
A�f�A@��̟\���0      @  � �           @       @     ˼�l :�Uت��͔ Ԩ���t���Q%  (Ԕ�k4�SC[u�Ѫ-j�4:tC]5B�]���                                        (      J��퇾���.�saA!� gp 8��`y�ޘ9=u�.�:� v(��U�C��е�I|   �|̡ꛘ��1p =�����GB��Nm'�tӈ�ۀ��X� 3j9�5ֆ��)������hվ   �      @ Ϣ������*���}uW��î�ϼ �b �ͯm�e�}�w����� �TS6<�a��YuӣUZ>   ��6����j��m�� �T�=eVۛUS �=76�R���UW�;K��w�*T���qbg6�t�֒�D�   �       P <�g�u�-�70j��!҇7 ��6��76���T>��{��}� ��Y���y������ڟ   0�hy@ꎸ 3��GUW�E9ڻa��縺�P�� 8�z.`��B���:R�k Ӟ���4�4�A�ݾ�����O  �          �BR��1��e �iJP}���{� �{igx J

ggK�i@��� �{�>����.}� ^z R���4�iJ\(D��lж��  _0�ǐ w7 ��� 7}� ��  � @27`�r��:��� 4��4��E��  �        �@{{ <��W�@v9 �� ��s r��r�����ָ �Gujˠs*�@��L�  � �v70�u� ���: dB@s��� � 1u�a������� | ��4�* �S�4�R�OS  ���R��� D�2�Q��� �Oښ&*T���C	4�I�B4l����_���^}��5����v�{}�9�Z��$�	&�O��`$�	&��BC�H@�`$�	'��$ I�HH~������������bj�����w�����3ۜ�9�����Kݺ��08�%Ә�)�U�%�Hz��˷��c�p<ܳ�9�1n�c���8Iwn��U��m��T�}}�q�B�a���G�B0r��0��8;���x\z-Z�{qgWB���.� �مGC�;�Kz�E7D�z���"�9����\���&��1p�`���6�H��|u�xp�7i�b�K��\�P����HV�#�G�f�3��Z�
UW Gp��-�^��.���)�ۺ4�\&���ok0o+p�n�TA����@4,��J:H��q	��B3Fv�|0��^��wh�=�_cĬz��ъC.�1a�����
��x�:'-�vq���S��CЭ�֨u	{���	t�<������#����V�r��Go}:oU�*凔�8��q=D�����w��+e�x���;�v0r�OPq�gQϱ=˃�ѣ	]6%�#8�D���2�k�ae�r��ͧTV�薊�{aS��\����Ub� TIW�Op���e�@� �C��������2�n^�]b_
֕7��H�=1f�'{a�i\�Ǯ�4&(A��V��,�;Jԙ8���d�(Xy�-�aع������R��9�Kz�mi�aÎs옻�MB2�蜖陳Od�aZw��:����.]���E'2�]	|	�;���]P���.�,�ǋv�xn`�҆S�ݠ̜�e�X�MO���3\ۜ(�sq��9d�������ɜU����n,���1�iÕ}�/4VIʞ��B½�F��t�qqdh2��4��-.�9���m�gnȎa�;���8�M���XYĻ�̰��$�1�bb���;��r�\C�k�s�NSs�<zs����3�Zs��:���oQ��(�6u��I�vjƁA��/ýĕ����7�$���o���Pif��]��,=���6����l�����[��^T���f��*�3hXFy�gJ�VJ���(����<(�Yw�ٌQ��W>Ԟk{2,�pM��r5��'��r��V�98�v����$�f��ݦ���e��)޲&��=�-}�ȴ�)�۳X��Ӣ�)l%��6iVbZ��,�V@V�Yt���y^�c�:`ӝ�I���*�K�-^ģ����лN���O<�.�%���o8m��M����Q�d�[�H��Z��xH准!720�������Q����p�h��.��<oK����E[��e�ٹ�+5!/1D !�ri�)�x�w�n��7���ӗw5�I�	�C�Cx=�N���U�Qz�zqQ$Ȋ��V�5	p ����L��%�����:�i�Br!]ѯ52�x�8�'v&�����.��;]F�͙Bտش����0�q�2�޹+v,�]�7u`��;��`=U��l�v[؞2gR�W�mįWd쓲*f�9�t]3Fv��#yf��9�F�rV-Ɖ��i������v�{�S�&^t5�3�A(b�ĭW)$a׃N��Y�h�c�Nn�1�0`���:h=�s�D2p��T�K�6s�:oV�U᷏�HQ78Wf�ӉIFh�n�!�����ǖ�6�}��ŷN���v�nƛ��s�lǀ�ځ7C�]<3����4W`�vD�n�1�&M�37�.�\�jeRo#�*�G����(Q!i�Nq?'���I�0�ˊ}�t�^^ �֡jwd�st%@�ӕl��w����Ta� W*<2�D�M,���j��2�˱4_qop��vh�`qCܵ�y�2��Lz���Dx\��fjw�7�_CRG\����5���ݡ[�nQ+y��N� �!���n�\��N�p�9km��M;�<�-սno#�+2�z	�m�\Z�dr�xY�xB �r��3��WB�EȠ�Ɍx����_Q��4�GRw��+G�}��hna��ֻ%�K.��,pƁ���D �c�u��f�؂C�r6��]_:�1#����`��ځ�N<x��ea�*5V�w�w�D6m���iY�5�&��Oh�sP����[���ǫ������8���:Mй��Λ���C�>ġ�4�}fGN�-7�u�$�<����4��68,�<�I����	9��8Os%��R����q5�7�n� f��% F�l1�.滫��z����ak!�rSM��>�����}Ɠ��S��NC�����'��@%�A�fӝڶ�Z��ב��n��5f�q>gSr��1؛Ρ�+�A��Y�
��|i�ǆ��f�()b#{�Ď��Dgr��뇫ȟX�ӟB��@*����J�@��0�$�f��{�]#�OJTV�Ӷ�/u^\�Xw@�=�CӜ0Y�t�t�\F%�8��e� 靇���� �HK���ղ��M�"L��͌��q^E�{V^[�l�v������Ѝ�����х�{U5�s��s�i-	�G1VF�%7��x�U֥�`Q|�C�h-�(8V��e�ظ⹶�c*�ق`kr3�e�����������8-��±ʽV�+�c��ˇ^ǃ�+�7��	�{B7d܄���S\�����h-Bpvoh3$��v����v�y=$G�j�ٝ�F�&7�<yY�@L%� J�Ti�ν,k ����>�b�ϖޘ�E4P�n�
��!��Lasp�d�Q��������G�bx�.�s��E�6`�M޸��Ȩԇf�a��'
�㣶�	�t��7�_^�s�t��;W�~�vk:rчDEj�����͢)�^�S��lX�#Q��B��v�e^^#rR�d�"I�::�ë[�EǓ������Qy�����f�Ta����-�>�a�09��PpŲ�du]D����S��k�z��i#�x1Z_9�JƲ-�EE�]�뽓z]cS-b.Noe��o\�FE�U��ˤ)�0so���h Me����8�qCu�4q/H
[���6���M9Hn�������o�ݸn�E�&N��o>!����E��7&R�ag)]/3���y6C���D��=/_on%�M���h�kg4No[w�
�}׀�:��M��d��ǌn�^�$�l�Qx-���u��d	�0��_.�g����MWnU ���9nn�Dێ��xHH�Ȧ��7ę�ݮW�JOe:`��m|�A���"9V�+�����p���ln���P�`[�	M���ċ�T�l�k�<x��z�u`�N�R�ˡ��f�[�W�p��+s�G �i^��l�S��nѕqG:[3rMT�b��gE�N�C�
��*4ߺL�mn�\C����`if���.;�4p�aѹڝ��q���eC�#����'����"4���ܗ��A1��w5�rߺY�k��(<�N�:��Jŵ��3�g�R����a�ځ�(w#[�'��V]����*'��M��ܟA�!�h��Y-�%YK��Sm�mxͯ�JW��J��}zv��g1a�{ס��뼲���ףe�:^׀����T���F����F�G�V�|�v�;n]R�e�NBB`1��8W��v��8"�o-�~'���ٻFY�|�=q�,����u�E�.�QԹ>)�T7$�9��ٛWE8^w2�Җ���)�g-dă�5���݌�^��y�i�z���.���;4�acCmoW	�*��pf�<�B�u��N,GOv_�i#��H�aoF�F[���N�ӛV��ۯ[�Bm�/zkbf����5"�bs0�]�齧u�q�����ъ�I7^م���d�x��Ni@\9j�6w篖�Gk]{K@̬���p��W�xU����O^3E5G���ir�4�[vk  $�Ws6�۰$��ys����h�X.��.Κ`1L#�懬�_0�ɌhLb81�6��'�v1�u11�S��c(�h<ƴ0�四a���t�.����bE+NhbL��-FJ�7�hN��D;ͽ� �]�=ۀl��I���z,���W�pR6} W��Ytr՛��N��-��z�[�Ȱf�5[q������ܙS��:ԗ���7^;��$�oi��8��G=������I(�-M�#u���v��X��"-c��IkcQ细j�n��U����Z���^R��o=:�O<��ZU��Y�u��h�зFDq���A���Z��ϻbSP�Y��;.pV��f+�6�tY��z7A嫘:d�DnrT����n�;\�5ޒ��f�M�dO����A��`�أ�:w'��7�1���	H'`3�腣����4Y�_�5f�n�$Y��8A�c;P��c���v�Z�V$W��Wr0�����ě�b���7����ja�Nn���ƺ�v���@� t��W�����(�s��8�u��6$���N�X ӽٜWnКw,�=��t�G��]ÅmӅ��+��q�*w乨v�t��J~N2Gr�2+I�w��I��xPd�Ee�#��>26nݍ�	kYݱ���X�J����ۇ��W���|Ӽ�tk��s�.�!��ӓdӏ4ŗ7�v�YĢ�ns{�"^�*0ٵ�5����I�\������u;)��ݝ��ĖH��p�0����]�������x>�	�����67յL�)�Ys�z�?n��xns�(���7KB-��7�s��m�8K��؄5��ȱu�Xq��奎/6�N�t��S��;�^��(w���V�&�(xԭA:n�,-�����1��
�7d��r�ǫ��|ns7t2�Cvo��jYt��5ÖA����9�o�r��r�ۇN%��5�㉱��!����P�7{�3�,���6vm|SI� �����Ӡ�� a����ˑ�jǛ��0	�ك�hT��Vq�ہ���{;*�A��I]f�W��&	3Sj�1l��v-�&��A;/�=]�g1�(|t �N��[(�x`& ��3$�A���Ș�E軪��'~`M#MM�vة]R��ꑉG����A�p͂�N��9��C��Y�-�7�]��z����i�
T��>o:�e^ۡN��Ky����ogNcO��͜����w.���7p׷�B�M�zu����q�d]�7zM]����� ,T���^9P�_R
G7Fl���Ws�C�X�5�e�2�/�{$)f����tA4QTiݏ�h��;9 ����\�u�8�{�Υ�ߢq�egx��&�rSake�Oۻw�Iɒķ;%�����S���4�!;��H�L#�DVI3�<��7�uߊ�f
�� �gpSTŧݜU�{���ș��ٔD������s(�-8n��i��Q�m��sZ��Z� �1�,l< ;�m+D]SjlD�M;0`��jy[p����Gr���Jzy��"t�H=���ya Lμ�>����-cDy�=mb#JsY��k��exvk��[�xT3��۪�7K@�U�m|�+}��e�ƻd���k�vbi��N�I��F����l@���5S�ͺC��٨��NQ�cr��r�F���MIp�UlL����]z���܇hJ=�f��Ś�ߏ�gY�̢u�����l*[F��s�ݡ�\ôP���Q@��2�[��
�W`���ۭ>�א+F0��\�%WN��f�.[D.CC�_"[0���l��^��R>/Aŧ��z�0�T,
-|On��� utΫ���vl�'nu҉TVK��[��9(�a鯔��}�L� �+/�f�����w5����3��b���"�uFw{���U�]�����U����晖]�i���yL�.LY��6s7n�H��
`�3t����)�,X�,�a��,N*���%�ǭ�Gf*�Z7�e�&\鹥췕pU24���6];݂��o��n�9n�N^���R��F��t��(�6qȠ��ݭJ�X�A�-=�y�a��{f�[�D����8w�M��E@8_F3��U�Pt2N�-Q1�����\��u��gKE.�I�I�)�B���~׋:�R���w,c�r�0�*).�A�<�a46D;'kn�OAƸ��Ġ!h�����R�#��]�oq���8�wzDp^X`�wD%l1;s{`��j[�ͫ�3eͩ7ܳÝ�T݃�mwQ9��ő]�M��G$蔋���,��v��{��V�ܐ=�n�V�"#����΄���ζ�>*bI�w�]���zA:?ӡLw
�ӕ���2M�&�1�d������󝼳���]�qm�����ۺ�V#/s�G1�H=l�u�����/-�B��S�%*�V��]�&m����f������G����'�l�w� ���������CFjQ`ߥF���3i�NE�eG�c����a�0k$�Nn��ssn���w��C�	�rb\���vL��q��Ԗ�v��-�'ܺ�SZ�#/f��b��݂�u��^�����Y5a���Iz!�U��)�f�{P{ڰ�UT!�R���v����7�I�̽�8oq�>��z�4A��& �{8{�I9��9{�y�����۞s�bH�HAH
@�X?�I �HJ�H�IYV
�%a!���VB@�dH��P	�!
��B ��$�,	$X@��XABH		Y!�, ���+! � 
I XAB
@P$
�@�$
!+B����@)	$�HH��$�	 T�HE�Y � `B$	XE$���!	$�����
�H@�+$�Y �$I ��,�� �R@���� �!  ��Aa$�d�Ad�H� 
,	"�� R(�HE��� ��B,�d��`@+$��Y aE	$
 
H�!PHHVB�x�HH0$�	'�����W����.�3u�vW��9d~���G
T$u�*a����[��ʱ��o*cw�K����K}E=���Yu~�[T�����)
� ��j�{��H��r�[Z�l���k��!�/!��KqK!+�13�ih����R`E]kobTl��ڙM�D�u�6�tu.+.�N�WsR1$ż�o�Nc�{rg;���g�Z!3�����ئ׫(�=i�{Rɩ�����6m��V����b~zM�1�N�m�o��f�5�-AԔ�>u��7�ǃqd~�����S[>�m/H�镟��=��7'��S�Z*��2@x����3P�AU���|��i���>)k�s����%���?eaJ����j�N�x��k�TN*f�D��ߩ���v�f)i�Ob�w�rQE�V��q�8}�{;؛u�f��z�wL{�e�R�&�7���~ԴL�`�=�=��h�8XO&���y}2j�ywW$��{^�����s���yme�~Vss6vr���+p�y���_d����};=g��MG��;��{�	z�E�Jg�?AQ�2�D�7~z+eߟ{}GB��w��G	%�>�S5������qI��8s�&��
拽����,/m����0L�������E���,���iq���*��-m�������@Uo�=���F�����\yv<��E^��)鷌U��`ɫ��O4�{9��5�xQ�.w�Cq��*3��۴����`�G�����yK�o��_��]�T,�qy��=£e�yȆzt�y�>���Ż\G���p2'�(�veD���r�PUt��\*���C;��]|����c9��}m��|M�O5^Q�M��h\�B�:Yևr��F�id>�V"���2��tZ����ZĦ�%ȓ�)��DRz&��-M�������[�ƴ1A�����ᑙ^�\7�䏺yy��N�#!$�{�q�)���b�9F0�o�ٝ8{<���ܛ|�M���TS�3*��R0�wV�$-f��yDTq8x͆���U�D&��Z'u���ov��y
~���ڜ�pIj��g�o��݋�|�~����>��p�t��w<�K7Q-�h���s�4.�F��DUg�N�)��*�������E�1�ݻ7���-�g4�/	�+	Gb�� \��;|��@��B���x�)�N��G=�E�^���F���k��Y Δa'��#�����uƳ��k9�7A�m]�G���N���������e}��J��!�|�#S��<Y��9��Į��l�ǐ^ˇp.��'�w�����qZ������S���ޚr����!�&+fSvZ��LƇ�Q�X�����Ҫ��G��b���br�e�Jm^�07nL�StUna��q�eI ��;�*�O��Q�g`��f�իo�Z�{f�[�y&Ws�j��ŧ����ŵ��!�(����KsN��[�=��]�o~Zo,��Z���L���Ҧy��9���n���m��F���*��?;���{o^!u��w+B&tE�!�FTDV
%�w�/���`������Og��޵<�vYY�������z����tD*z�ͻ��[�`܅,+�j��Ϟ��<=H���t�Rb��{��>L�!����zm�&u��k��2����o�NV&�u�F��n	�Y)Gޞd+�x���vN�Uܣ;p�4���l(s�8
�ݛ���\�:,�ۮ��ṽ�pF`��hmщq>~�[�-n�/�5w�ө�/׹-�?c�����z���<��Q;6�Mu��z�7B}���`�8�po{
��&Ao���5m�B��1KqmE*��X��Jt��:zu�8kJ�0��Iӎ�hn��9%��t���4�-��J�ٹN uR���;���9C~��C�}��k�_M��gep�V&Fo}�G�
t0�gt�֭V-�Z�!]!`��DzU�v��g���A�w���k}���u�7'֜A\ �-g�=���{u�O��"�~g���T�{�w/{��o��?lP�>Qv��+��D�"�ɣ�{O�S��r�î���=;v�Ij^^��_<O�+�<0�9O�y_>	�D�Mm42�pk�I�z���&����+�}I�ѓl|7��糊U�#-O*g{G�D��j�g�Jtu�ȫ��Z��d\��.F*,J+6�TR�=�M*Z�,���?�2�Y�!=l�q0nM��j���e���G�E"jp���YQ@�^Z�/7&�b�nrd0T�G���g����v.Ci�{/�1K1�ѹ_�On��*��#Bn�z�(��r'�9\]��C��&�m�G�V����+�b�{ch������E��\}�o�	�3���c��haA�j\8X�ّ�R P���x�:8�<#�lk��G��;����<	w�� S��O��m�Rqc���Y�SJ!m~�]Sپ�YP�5�)�I�f�P�$5:iޢc�!���{��P�u75e���g����VS��*o_+�ƭޙ�hX"�:��'�6)���q=�lw3}�>�rt���S�w��P�2{���qx������ӝ�vO�O�x�'��a��׳�Y#6��U{�4Ss�Rf4�;t�� �D;�����N�O��n����plF^]�b������(Eث�0�Q��y�,���X&j�OX2���#��h~¬4z�N3Xa��Z9��u�%��־�z�o9�N�^Q�:�"�>���I!�	��Ɲصr$m㆖n���	��2"�.��2{ӂ��`��L�um^f9�5o-y���e�;ue����L��N��R�XWC�P��`�$���)��@\�`�V�`�<�V�m�I� _]>�un�tI���ތ-�C�����ó���b(�֚I���R����~!nQ!'�����LP��u&��� �ւY����xT��%�/���"��
ͷ�R�1֣�3���0]�G���9���^��}���,;wD ���`�x���V����h�=��Ϡc��	+�g�]�r��r���n^'7O�����ݴ�-d�B���O�{�l��{6�V�2���B��F�
Q��d�v]5bT�������Q��!�p̑�g�ey���F��,����eŽ�U�EH�k�f"�"��4�� 1�	U�31��)=cx��<�����:�r���)�{|vf�|̃ϒ�E����ijG�ǰ��6g4k��lΑnr����0�1U��"ǝ�?vx8m\���{:�x3���\]�7$�=O���V�*���ݎ��Q3.ēY�>�b�e��P���	L��ռ�SlWw*ԑ�C���83N��j�ا��ŠX����^�A{e𗽫��^�;�q�Q2�9��V�fuhΐ�\^N;Y�Xmhȵ �B5����z�nM�&�q u�U��������<uB�M�����/�Ճ��&�`�����bZGW�]�3n?O��3ȵ����8���E�^;�OR���O|wk��k�,�C3�YT0��5bY�_I�&9�7��I�{��pmK���0���^�g��^�������*��.��E�)�x{4��������9�ΠN�y��� ����w�;��X���z�.�ىj{�ĢS[�&��&w{����1���	��ׂ-Y�w�{nz,m.7�7)0���	g�[����y����}�Px��y��X`��H�����#9܀ʊ�̓��Ѫ��b�����\�G��;�X��8*��f���>ޓ�ӽ�k����x����oއ|{�.�F������s�H>�yL�U�^!tMu�suY2�Rf+�=Ђ��J�r�N�C|}���z�����1?wpz�2ϢA�}��o�)YxiT�6����G�*�����7��ޓ|}�̝ത.�0Z�%FK2��+�Fhaq�^��� '���ܮ�o��b�Z'�-4���Ѭ�֠c���נ^�jd�Fcj���8p��e�J�2�s�9A��B�=i�����/��c�{��7�B����X>�i��h�"i�Y����T`�(k��x+T���3��T�G��������%*xǭ�gJg����x��Y���~�i�|�m.]K�;
R͝�|GL�׶���N�Nn�%�_>*�o��=��u?y���f��ga��y��ͳf��q��ý�D1��e8Ux�KG���8��vE�7\��pv�\aoB�.+Yh��r�UH�*Xmee�ê�ֵ��ocwNj��n6ka��!Tz�Fl;�jsn�<���L�Q�}����o��(*ŉ`7.9��D���+�r��q*�����U����3�0:"��t����/D�@Lw�q�b���8�p#d75EA���tl'y����R�]KI7\�+����UXҊDR����t*����3R��]��c�ۆq��@��·F����h��	XssQƴ�d�)�xZ�b�"Zsɤ����Y;���7q�����5�3��ݯ.�VX3ut�9�^�z��O���#>V�v.���-yuP@PB�1;�}��vٳ:�0Φ5�7�f��}2F�� �L�:�_;���0�J_����Q�`�z��.��` ��[{�Zyi�����g\^p�ԛ�GS8f��9�3�q9�{�y^�濒�63Z	���:��-�p?G���ʔ�S�!
��[�0Ika[�*Z�}`�eöy�ǥƶz���om4����\�!<�X��%V�N�_e��.c�\!�@��WFoxH(��qi�ۀ�k��1
O�\W\�h8�`��	C�ē.ی�X��Ggt�<.k��Wl%��<������%��,��	�Ѳ���5�7��9���7B��Ȝ2ɪ,O�&�g�~b���gM�u Oό(T9HV�Ւ��o(@�r�Ijb���N���9���)?Y��_\t�����[�/.�{Y�ɺg�C��am)sj6h8�xM=y��^�.�Y�*JX�r����-���egK�jy�[2^�k���iR6U��$�t)8��.�h�9��	�^P�1v����ǭ�qe˽to���=>���7�ي�=�cç{��.�ދ��V�Z�t�ĶQq0j�.�<�֐�_�s�{f�w��xG��B<�d����Yq���iƹ��tͰS�{s�)�J'U�,�-T�ځǿt�`Z�v��H�w\�u����x��MS&���v��"&gg�n��~҅g�8-7����d�ܤ��N��XH3�W��K�LvyV��� ���<���~$\V�v�`��u�pl)*���К������m�)��qG��v�[�!N`�N���}�+�]4b�����6��I�RO7��K����7լZ��i��Ѵ�T��:�C���N��fsO �:�s�������'������-"��Q�MJ����ͼ�������ڼ���Ӻ�-��"�lJ$����s�XT^Q k��a���{�4t�!/VaRxg'�?-��UE�']�����2U�c���q:�m�{R %xz{k�{�1��j�HݫB��*�,f��U!���w*� ȝ���0R��y�dP��eL�������� �L���ќC4���b�����y9���w�q[n�ݸ�Î=�f�0h#}��7���MK
�U������Ns����t[0lܻ<CG��k��^�V�ޯ9��W��^����z��sŜ�S�Q��K�m�H�#�v�F��W�ʻ}��>�����f�@ĸ�>����3�vTlnV�_%&�?`NULb��������K�m�(8����},���}#DE���b5$i7L�SA���;}w�]J�G5�]��Q�|:k��x�!�W,�y)�i�>�N��������o��IM���N�J��Ӆ���i���O�ރ�Ly������x=�JO�{�eZ��5]H�U[�|Vi0oL(&��&v��7M)�B��{�z�9�5���}g���T�狧H��>�=��v�)�0�ͫ�bW��kl��o��Y���	>��`D��lަ��!�o{�q��7�:p�����A��{����{����
�z��q���F.�'[9�,��;Ȯ��]��4F�m�M]9�SG]�4D�v���OnJk����r��{�r�k睷���e���	��v����C�B�ج�� ���ރof�j���$ؤ�VLu<�⏅�}�Y�;�/��9��%m5��՜4�[�n�q�1"`c4Ě���>�/�b��y���2�a�z\f�Ǚ��z���i���fվ��W�E�"����S��Uor�]��=[{�<�͑j����y��VW�3����]Ԡ��ݑ6�Yp���`�;���{B����!s��
� �fZ��R��ɭ	\RحQ8��F�;��\�'m�'m;4�z���c�q��Ӄ�I�}9|p׮��W��_�������v��"���b��=a�}�z���cx���4�YyX�{���ۻ��e�u��kS�8���仾]Ǯ�h��_����P���{����0�f�P�{^v{)WՕ�^�;$�R�^���.�3�̔Z۝-!5�ZĦ/\Q�P�Hy��R�d���[��� �6��|w!S����;�]���`��;a\N��=��K|*Dg�s{�d�
�z��v�R�n���U��L��Ɲɧ��:�v�S��(�ʽ��W�6V��3���d`p��hlE����)x�8�>��^�L��_݂�{��{pzl�%����#�bѶ�o,��|�=g=۹�<�C�&�|�Oؘ�o������w��7����	!I�$�{���n/0�z�䅶�W�	t��a�OZ9غ{v�֎����3��h�����`F��
�r��6[��b�1��yb_n������u�ûu{Mێ9;<�:�Ӡ�ͻ\<[l��`�p7hMO͇��ň.N�Z�^�=\N�M��<]�2]��<�>*��Z�#���;Op��K��3�c�Y�^�r3��=S��y�U��8���݄|�+��6�<V3�M\r�`s;���4�[���{=��A������L�8�ٟ�nv�:�i.�:�lu���-�<i�8���u�	cj	�M������}�]��`{O]�Zq(�{n�ɲ>�����魜`ݪձP�s��׷l��#����֯ �oc\��ۑ�yRێ!�A�5��|��!y�sH:80v�XMx�!�8���p>u�s�5۱ڣ!�eYK���W��)v�`ź�<�7n9���׷�cv��l7Z�"p'q�ف�n5֛��ɱ�����zX�B�����GXw�>#q�8���흄v1��SsYv�ܥӻ�3���N�:Ʈ��4���BP�ݺ���&�vC�n7n1ܛ�`�ᱼ�^�(�h�1��M���[��^�{f4�\��m�#ώ#C���A��g����]q��w���;sn�`n�k��q�mӫ����.G5�;�y,��<�^�-���l��n�����N�ϑ.=�{�#��ۮ����Δ�ͧ[9[$�[e�����i#z��n�|���6H4���:�݁4�Y]�s�q��-�| +b�j����͌3�8�[�l����[��i��'��۝t&K���� ��u��P��l/<	s���3��6��ܝ��\6�$�۱�]�-��֚�s���ܷM�+���Wr\�GZF;s��ɅP�F��"gm��9q������:C�lg=��ێ�Я��
N<v7X3p�h�[d�����A�Z�9���]D{t��F��x4mW&8���u��O0�vg��{ �M��V��N��쑌��k�ݦ�l�3U�b�*1l���*s�c]�]��ӂ�����mm%����u�B��%7u֮϶�/�a���6+�M�d��I��]��䬜�Ͷ�m�V{zM�n�kgXg6G�S����Q��b��v����5F㋛2B<�Z�����&{Fn<v;[{3����ss��u��lu�vq��v�\�ќ��.#u�*����v��W!����gx�`y���a�Kd��y��N^��q����r:0�[�-�9�ݺ9Y9�nv����k�;pv�m���3F;rf�nۇ&�2i=2�6��/#�^x�l��z��&;;�M���b<k׍\���8e纂���ak��k���x�{"�-�n�׭m��C�8�i�:H.�)p��<]Q�غ��n�L�ldx�[H����u�w]�g��v=�uϷ%�]�-�[��N�A�+���ƞ7$��<�F����om�[�&}c�����'c����H��\�ԩ��m���h۞Ö��٦G��>Z8DNt���p�[�����y���۲]�8�K�V�WIϩz9�au㱣b^��#��{@v���]��Q���mm�\�����t���!�<���l,��B��㚬�b�[{k�j$��q���w&��ܻ��k����<k�si��Tl�ۈ.�q��ײ9{�n������\Ok۟ ]�� Q�]���z��G츳����E���w<[XG;�������GN�;v왳���]eκ�Iz_Xgv׈ՠ�����&90;<�k�5k9 ��b��퇍n#m/l�m�B$�qufaۀ# ����M�Ȼ̄y(��(p`qFd�O[�ke�
N�X�pv�=��v7�:�')��Ń��X��pu���Z䚠n��d{��Eȑ�m��!�Z;vv5Z���Ms�*v0]cv��6���x���c���ݞ�����¢������w\��3��\�og��v�[۝ҧ�ۛ>�8�y���r�ln�-nѵn�!`v����8�R�(�<�ۧqJ���7�6;���uݛ����M��;^v����z�v�uϻ{u�1V.uS��[�1ے#��㳌u(+u�d���tv]Ƭ�1뷉�v�ݠ�[�e��Cn�/;˺#�ܪ���0pth;[��.�1��1�O6�m��m�s�L׍��ݤ���Ǜ7a�&�wq��;]1g�cp�[�	�ڇ�\��BXu�3�vη���^�ݝ��S��N�]�Ϋ{���W����C�c���\��z���w<[��@v��2���f2p0�	�����q��䷶B��Þ�7R��77�����Ǎ�];E؝���/]`�x�s�	;]q�k����ɵԖ\�Tj�/a�5�x����Out��s�m�Gg����ݎu� U�Z�g��Se�6[�9��'�=�"�5�c��pN�q��&C�#�GZ�S��iG��j�8�f&��͡]۳�ڞ2��[u�J�@��n`��;o6q�v�8ɬ�֑���}X�u�ݮI9��t�y1��ԛv�t�x��a�p��9n�5�uƀړ�l9ܽ/]��dJ�Gę2v���v���X�\4B��܈��f휢�1��Wf��fH����8x�\�^���&Hv3����z1�ggY����Y��b��ٱ���@�-���to���e{���7�g�˹�sm��a��ʹ=�v#v��M�w��p�=����
g���t3f8��Nx��t�p=؞�����(]��y������shc�.Ԧ��ݷ��ں7���]
cf��-��sv��sg�vN��c78�=WC�GZv�����n�{�5�ЄO��i.�[��Y����8��Ƭ�z�>9�u�E�����p�v�;=�E�]��bS�!��r��6�W�Z��^z��\k��.�F���=:�����M���n�6W	�ӟkV�:f�`��=n�i�<k4��]��c��ز����!��e1!�\= 0���(�.�����9bc�A��n4�x�FM�t��Ϡ��<�=�������c��f���ۋ����)�v�nq�e�2<��6��u�'�v7t����*gJn�^�ץ7�;���7\s)gusq�����X7۶	x���3�lv�h\�s��ݲh�:�v��#��.�F��L���Y˶��{vCkˊ!�݃���	9m��-��7o;r���.�״����c����7��a࡮�q����;�:�b�n�l[�7j�';���瞻C4�'q����n(�vM�l��v�Eg{[��&��l�v�y���9J��]e����N��uT�������C�د*ݞ�(9�6�36\m��5/W��n��q��)���&�Gms�V����o'�mv��р^er������u)d��c����nm��N�6�.��b���y[�b��S��+����
��U��BH�N�Np.ۣ������Ş�mv�ϴ]\q�j�+���[�rX_E�u6�l	74y�zմ�ɞ��]ms����Ƕճ��Lg���ɓ�����Y66��\��4��nLɝ�ջ��\�r�'�ݒv]�a��n;�'Z;������V��b%5����v.]�n���u�<\8��]e}�q/an]�h�.���˶�M͍���s�nީ���2���m�u�@9�}�m���\-����W-�\�u������&�x�y� �4�;e܌�[N��f�r�,��Y`���alh�m��%�ls���T�Y�tc`�+�,�ݸ�0��pQ�5� wW��3�1��v���ڶĠ=�gD��ܶۅ�4!��В��V���n����DH;;]�zt�Ӕ��Mq���s�8lwDu�tK���s�Gv���I�X*�sv����g����{�k���ƺ���Sc]��'d&�wHp���9�]��z�9�l��vu{g��(��O)hl[�5½�j[8��kp��0�p�����ܳqeӸ�sh�M2�Pn����v5a���) m�;l�z�2��7F�p��9�M֞��i�3�dw.bT���ʃ��Rֳ��c�bȝ�Ӷ$�q9�x�X�0��*O;�ܛOn8Kƫ����]����vW�p�3^�p�;x-�apF�j�ݜ�mj��.w�^��B�uչ�^5ҘM��w<Ǔ�j�sJ8l���6��6�:g�b��l�OIے�n8�=շN�u��{q�:�t��q�T���s�@��y��v}XKԗUr(�Þ���f�\x�j�2;-k���\�s6�n�k:�n���nR#��\n����H��v�y��S��=�۞��і�-�c7`�,�$x캞��]��n��V��4*;a��&N������^wZ��l�;�ayܻN�V룬E8�����$�re'��c��"�۷1����V.ۧvB�GiN�qj�*�l�װ������"��=�8-	uv;A�.rON�U�\�5`�'i�q�ݓj3B��B����㴖.h��$`Sj�5��mɅ;{;-O)1^�m]m�&^�j�Ta����۵�{L� V9H����x��J�q�Gk�Z��uCŝ���6�1P�랸s�㔙�q]$��o[!���z,�ݺ���[��m�{�%-N�W��>9���;w9�YѶ����6�:�%;��j�u۲�r�읲�])Cq��i����yݞ�g̠�o]^y5nc�g]=�[c�K˗�x���F��Y�l��qf��i=�W��n}��ְ����b�]e�z�h�8F뺻�u<�c���S�m�����v$�nrlg�p�K��������\g�g�b�v�\M�x�Q����݋��ַZ�����nˬ.�Cs^��-m���
T���aZ�
ԥZT�TQI[i�Uke����a{nR���ڣR�KUK�̶�aiV,��Z��2��-��U�b��)Pm����V���Lˑ��[`�\qh�ѥ�)iG0�Z�V�iD��-�V����
TJf+\��j*W0���!��!�E�Pm*�A��j����QAT�̨�Lj6����1s�*֥J�h*�2����Y�Ҋ(Ȩ�X�(��`��W3�����[A�Q��-�Dq���U�m�(T���5�A�����mf&*��l�0̱+�F��-V��A���1̤R��[hԢ����bZfX�cZ��¢*��R�2TK(�`�bԲ�FT�m(6[h�°��Q-iaFֱ��TUU�*)�H�F�X��X��!mXVRV6�V����U��ZR�*+m11r�j���YEP����eH�ETmlh��m�%(����������V�q�Y74����Q�^�U���ܷZ��ZV��rU��no[����}5Փa�nMB�!���\81�{<��ǁ�8�;E�:�9��iq�5�D0���&7�捵�=���9��gk\�m��cn:�������v�Z�-)î:�%�w�\�O<�%���7
��m�ݻ7#���]��A0�ק&�rn;��<�>�n������ݹ�Sl����n�b�l�g�@�m��e�a#��ޅ�y�����&�$hф�瞱�;쇛��]p�i�����Ľcg��kb�ZX��G\{sv�v1r����vy���A�s�q�㴛��@[���S���]��]�<�^ �t����]�����wIP��NvnGn�-���pq;cζ��x۶x�;�|q�198�9�+��ݸ�#\s��ʝ��Ǜ������v�����3�wXu��kn�{r25Ӣ��g�-[��K�1�ex��m1�s�"R6���*Ƈ���>r��Ș���-퉻Bݭ�ɵ�{�K��9|�slF�M3�`�ǝzN�l���C�����.]� ���ܜ9���\�8�Y��6�	�.ts\ռ�c���K�xS`ҹ6��Q�]�A��v�7m�G���O�P!��ì��aHd��.u��d��]v�݂=s��mA�dݓ�n��jaO�s������8��v�z�<���:�[׮�G��sm�;k�c�P��O=[l����rܐ779�[���8M�.��
vt�;��a��+� �;�m�c[#��}�l������x�������k]����m����v���|�'�8��Qa���C]���Ml���λS�ǃ�b�jx���]�]^wNuq�@V2Wk9Γ�c��m�u�3
��`�ք�9��fii��Au��D!�ݎ�1�vnŏ1�����o ec) ��\�]����r�n
y��퐛/www]��wo&�ö�ϝ�\�l�pl��#���3��ɎW����pp�;o>E�{s���W
6%2S0n9rjԲ�0��ǹL������v��(�(&�cn�/m��v�0����z˗3��Z��3L-S)KM�v pm�0���r�6�*�Z-U��R���Jp�ɻ�̀���
.�T� �ہ�㝸�y&q��B S���_�?��d�ls'�}o�9w! @)�l ��mJY���u��Bfb��<���� |���b�����\4K�e�/z��\�$s�R��NVć��SU |��n� <�[]������Hs[�iȦĲZ��q ���( ���q��ٵy��ܜ�w=8�6��L�`����Lʵ�s�n-:U�.�l| *�:��0��v u���\�ע��[�� f����6
��fG����vڸ 6�z�K����/;7R�N�J���#�̶��.����Oo��Y�]\X��Ɖ�3D�$A�&�v�w9�(j��<��6��M)J
�i�}q�9�R�T��}f�bD,ܫ�$��z��^���=>A��9�I{��Z�c�KM˙)lzr�� I�������������sD�i�F�0���thӐҢ̭�iʝ��pOxxe�z�F�Oenm������� {r�� D}=bV��f�v���^�/q$	�\4K�e��޻��.�����Ki5샺e>����Ihb��w ��O]ɭv)cD�jY0�Ӱ�����KJ&�/������>O��("6��� |��񵯻'�'�o^�˛�'���*R%L���kӷq! |:�3g��H� ��뛀 +vv�$I%������w����N�3� �$K]z�z-d��>'95���V>�<It����̎%1�7k�D[��q!� FW]#��_u�C�tXY:��� �rz�BF,󑩖�F�L��~��|팙�1�MכW�[@[��� �>n�)7Q�a�c��,��i��r�JVmt�܀^��� �v�vF�NE��Z��)ڙ�2�G������ؘ�7j�{r�K�6*~��?����M��S�����/���&�w3�}���@$G�nO]Ĉ�ϛ�4[��%�D�v.WuK0U�{�O�\�{�>�X A�)����ݔ�Gl�]�bz�=W!�g��a0��L56� ߝE�Z�ʸ�1��,��9 E��ؕ���I%_iݖ�S�o?zu�����13�u�./kv�v�tv�\�p��q�,sv�4��X��4�ο���;�$W�d�:��we;��SR�z}���nI˝�+�K�7P�����S���� /ә�'�ޜ�}  y�5@��v[�� "��w�~�vd�r#�EFf������$t��dO-ܫ� ^���/s�^�	���Iwe��>흃`Ne̹c-\]9~^�.q^�O�=�%���j�4�e��I=��r�8B�,�.�O�׳�͙�j[����az����������<�
�H�����F����x����_���ج���o�}-�h�o���-�	S�\�,�~���OUĄ9�f��̻��7� +��� 3��� @����O�:?B�y�H6P�Ȝ�Ӈ#r�fΫGkO������Y�EA��[��-�??;��m�:i��u����P|	Z�ʸ�I�OQp�uYR�qE������we� ��Y���J�V��z�����^�ՓXȜ�Hjj�^�32�W�=��}���.Ms�3���0į��28��vZ�۸��I�OU�H@���}� @fe� ����b�>j��*e]�+�7�ѵӗ��o��� �{*ℒ!�_X���͹���٪��5��6 ������@�cm�-\]9w �׮���>!O�~^���޷`|�=w" >m-L����V&�'?=�����^�F��V�;h���Y�����t�<���5��z=��nc�#a���ج,��T��5�[���=5u-���f۞=@jy_Z�t���k)��<l�V������~{���voX�mvݎg)�\T����Um�J
6��c����ɺ��q�Ѵ��(�]M�[��G=����K����@���1�v''k�.�	��2%.ˡ:�	�����u��a�����O���nu�㣺�;�=�������k*\��s��7g]v.ú�j�랷rq�ٷ��c�s���wX�u"D<����)�mA.]���@\f����ͪkd��g�k���5;�~���Uݻ� �n��	��cJ��j1v�=�^2IQN�5�~���+>����ۛ����M��kݳ���6߀�)�	��.�U���� ��TT�@o*������I+��3�؈ <�D��1+��r��ӵK{id�(�cȰ�܀"��P� �� |q���ʳ���ё���Nج�Պ|�9��jQ1v
�;U'� r��j:��Ƿ�����O���K�yԈ4��w����F�/�m����;k΋�,�=m�K<��1����r�S�q�9�"7����Sj�njm�?M뜻� 9ڈ� �ս��ڞ�yq%z�����+�x�@i�"�&_Ĺv.WuM{���}��Ov�x�C�熁��0.�u�\��I�ͩ�(�(���[�8]GE��6���7E�[䗋- ���_��ds#�Z�e�C ���IPoe��J߲Z��=�<��D�m��ML(�r���p_�C�ge] �j����<���@��4���`��u�IP��ʂU\Gu۩���\7�� �$�uI#M̷`|�+3+:�̻A��s@A�����G����-v��P�r�긣-�tj�.�UG�|�r��Wܐ�g!��⵮R�	5 ��5=A//(��.�s�9����������S�s�#w���X���2�-J&3���L-�r�X��n��������c�.nܤ����)n�(rԒ�6唷�;�.�K��t.�x�2{�� >Ӳ�+ ��뤬2z�s}���=������ɔ	LL��r�|z�ؐW�W �gn�,�~1yˊ��Q��<���Q�T[ƶ�D��&L��e\�
#��Ì�DW�m)���4:���th��g��:��q��uv��;6���&r�I+���h\D�ȉ7FA5&��D��u��_{�K�� �.��|��n�K�9�;�cu�n)L��>�9뛀 ��m�
X��%]�F��  0|�!Ǣ~UT�{nR� �3�؈���.L���+�P�+�V�
������z�t^��&'nwF��]�nXs-���x1-�X��Ӿ���l �;�ؐ9U ����t�2�o߹��}�r�Np�7�(঍	cM�}�B�3N��ݷ5}^�A$��Y>Q<��!�=$�sŬ�\6$cRK�ۖTo�	B�;�B�@��D����h*�]ĂM��s�O9k��LDH��D�ѱ�1.o�;�=<:|D8�'ĂGD���λS����8^Yf���7�/�K�Pl]�gvXϷ�.����ȝ�''��OI��w����;�����6���֥ұ�R�b�'�f
=�N��b�9NрDMI�)#��&��N�m%��r�8�� �N�[����pt��w������q�����t�n��f�{duͲ������q��֦�
����5��ĝ��\'�0����9�j@5ӊa!	'x�n	�ީ�i>ɯ�9�6K$��1I[�i.��탚�K�<�$�3�l�����N��j/:/��0�B�Ȩ�4bE�e>�t��@�n�W5�b/UG��'��6	�/�<a�5P�SSP�.�ntt�]Jv�e��@�9��>��EQ�s �.3��+g��0dLעjhߞe�@��7�:r�f���k�Wt���y��$S���K�Ê�	���l��`���Nr�k�<�PaM�E������M��`Ӎ֖�
����e@-�M3G�d�to2g��V	�7�
�ch͇�VɈuQ�z8��Y�r��#h�Z:�\��#����9t������8!�Hk��9ۃK��[��ȡZ1\l�Л�w�D����g0;�m�/c�y�N����u��y���o�Z�C��׷1�
rn�bv��v�n�;�L�a�ܽ���Y����=,{�;�;)q�|�-�e�nR�L��QM���q�\&��㴃��X���{���aw:7�2�CfF��u����~�NJ�ΰ9�pv!f*�U��$��"�;13>3PjH�6g�u� ����>輱v�zw5"A&�;�}ZʂH�}ӉfM��$L;��λ�>$ӎw� �]�����9�҉.{:�$q�`I80ᙕ�j�TE������'�ugXD�}N{��'"y�H\�������/9_3���@34MMBE�vؒe�����3��� ��� �N�3�C�l�]��k��?���ɸKb:�^�ŷ-/	;v�st�:��ƌ�fP�`�O����~ð��έ���x�$S��A ��<��0�(�CZ��VBJ���g������\�e�]����Q&iA�Ka߫�{A)y@�wM>0w�o�D��ւ״���Bl֋�0��XY�Dr�FA�8]ѥ'M����+��Y �r,���:&�����J!Cq�32���RW��]b}�y�H�Uow���`�+�uE%�{f�9�lDJr�L;����j���",��Sf�by͓�Ds�_�3�~��wݫn1.�́���B�"��eo_��#������_P�U\o��y͒	�7ڗ��&���>�G��}������W@:�lH�Ƈ�]'ݞ˚\��][~�����n&m��}��t�$�/o�	"�H���uLh�p��j����餻���R
be�H�~]��$�</���Q��FD�M�c�m��[�����N�
=:* ���DRE��tI�H�%�s��,Y�|��I�l2�7n��X��$�<ѧ�j}�Ow�����^�{��L�_j0Ü�W�{\Ǝ�5���}X��2�^)�S��Їt��{�p%n��r��N#Z}
g�H�}|�����#ݾ}1�P�+K����wa�C�0���;n�M�t�cv{���3�n�[��s{R�	6���c�^u��.�@�p�~����*ާ՘��8��k�Qu;�����殷b��t�h~E�o���3��]A��?dxƆ��8׊���l��yU{އۢJ"P�j6qf��3j��՝|u����3y��"�Mބ{�@���&v�tR�h�y{�g�q�f�Ѥ+MZ�ų��<�4W���Y��|q|ow(�����]�璨-�1X�������˹]�Y������iW��HdB�\��*��G��ꀨ�ƶF�FCSZT�1�S�s�[��E�{"�3�����:�M�ZeA��zնy����.������]����=3Y~=��S�V���^݃��j:��ӽ�&��r�3n���T֝HxV|̍𷪋7e��/�.��|O<�U�3њ���Xj
L�qM��7���С�t�0"�i��di��կ�ބDq3������dA�o�(#��4=���o�t�r�D�8\�{n\��"�(�2�$�+E)�M\���"��Jқ��$������T��+o�+��)Xuo�0�	��2�e�J�X���2�((��6��֩i[J�j��*4�V5)l�UuLC��Q�ڨU[`�+Ph�7.emb��Z[*#Z�AQ`�Ub��QJ�UPm*ԪT������lUPE�JV�G���YZ��H���A�Ũ�*-m*(�jU���R(1��QD�-�Z��ej��"�D�A�X���6�¶0��V#-e)X"�(�2��Z*��E�(� �Ƣ�Qq�2���%��Db�+cE�����V1-
��
-��DD�"�ċ-��c��(�ڈ�j�D`�h���1`ʖ(�J�ER�1-�AU-�AJ�ڰE[iZ*�R��-Zƴ�E�P�Ţ�AB�6�"����!iiHU�-��*"��,R�dUb���mPD+DQm�DJ5Qҩm"1UEU����!K(�jUQ�jՒ�X�YclD+k"�ou��z>����U����E1�2L@4�����]�1}YWe�H�k��A ���@�E>��k[T�15��K���D�*G�û���$�O��9������,�h�F�M�A>���� ����m�1s;��M]{x��Ɛ�`_	q�V��-���݀�.�XƆ=�ŊIߤ�-6;�Kwi��ٹV�I�O*�K{9s�����u4�$#^�D��a�4h��&���]8t�s���M��X^�|A�ǩx�+�z�s��s]��)d��|�v�D�J���7�ى/O�toX�	'z���n���D7R�@5��r}9O
�&(Q��+2{L���ė�j��>5ѽ����9�#G�����Q�{��p:Qe���f�'���y�5�-�6��:�d�$���]o���O���ѐhΠ��������s�L���c�.�$�p�u��q�[��T���tc�H �T�AF�"vwqꨗ�xB	��'�!B��Pv��[�R�x,��D��Bs���&�������?KrH�+y'ܑ �N9ܒ	S�V
�C���ݗ3�ļH'ƶ7�I8f%x�3F��Z��gm�^�U��ݍ	'�qP�VOt�$���*��wm�%�ѩKM&�cc��[GeD���j��D�a�BQ8�I�O_�$��Gu���6	M���"$Mzf*��]�t������������B�S 3߯t���j�ݪ1�ڔlo�ӐЂX��6�z��;mx��5W�;��>q9�`	��ԁ�U�*������[Y?��ŷ}4ֆ�6s���(^h���=����f��֖�����'�j�^���8���ៗ�?��n���M��2ͨ�5���;��AAI"O�È�K�d��m�sU���ac�<�枹�����77��#��;/mm��wH�c]�8��C�Ŭ꺔�m�k�ey�ku������z8�|�m��p��;mŘ�s�ʧm���tI֨���S�)�ZCOD6���=x�7' ��هv4���<"�nI���i; O[=q��N;w��v��q�����5��[I9��`;Q9��9��U�L�3�c�;�A�q����l�z�PHv���b�<<���9���S̻����3���H�ڑs��3�F��+�A�#�^̓P�A�&(MI*�y�x��>�5�L^��K��6�ڐ'�ǈ��X��BW�C��B��P4,k�����l O��Ó0���lj�,N�:�O��}� y�L�@R���5p���6P)��%{uK䉌�ԁ��s�6f���:r�_h�@�������±o�����wv` |yF��*2�ӑ�*	�9���H�Wm�(K�%��;����$w�)�fi]%5�u�9���vK0l�u4�k�����-箋sO���b���"�>!�˿.��@�KS��:��Ϋ�����Hպ��#�L���"b�T.�
�̸	�Y��V�3�s��p�e]�8�B�?2��Z���$��ʟ!d�:ݟU^�%aK���5��K�T��B�WOf�$��*��٭�> ��ԁ$������6��[O��B_⭴Bc��)+y�/	��r	Ƴ|���]T0u�hr����PeQ�U&hY�����X��H�fZ����[�s��B�)��'��4�7��UP�Է37i��R��Q��U�xRF>�\�$�P݉� ��^nvb�Fm(���g���gn�z�t񋆺\᷇������ �v��5ЇA�)u��������<�]T}�1$A<�]�O� ��VDv��GN;3o+��^�6�'bo�:SB	b���CY��d��	.�i�\��$T�_$�{_�I�7G]�\�2�#�9��1$R�1`���I'�d� �����r�!�La]��T��V֣�۾�o/lR���~*��m;y��7����G*���?1�9RG�Xc�h��������������^���|T�&7��P�j(EQ)!k��j���)�j�K�{R�$�Ok��t��v{U^+�IL���Ǿ��I2��,Y�߬���lvS� ��pO�g�_���ά�}��Ra
������r=����+��7����M�.Kd��<�6��태�����ߧ�n&�J�?x��زH�{b���v��_�s�m����A�-Ւ��Q�M�5$I�����_v*�0�ğ�NN�Y �=ڐ#�����*a�g��DV�t���4�m��I/��vU�$��wP��#A���<I%�ڿ	{�"����%BNaKIP�;�#��K��D�����~#%���If��9��^���m��M��7v�I
��������^ ��A��2r�؞��
��\*�s�D�FDfv�zL�U��G^�nD�U4L��ehN��MS��:nMɊ�$Uշ��!��~��8�Z�B �c{��>��ԁ �k��=i���?����߶�g�z���y�OWg�xg������ۧ��!��ܷ8��������JF��^7B�r�m	'����)ɋ��ެ��bM�w��H=-�w^�j�55Q5S�4w��(��o'W^���Ƨd�	�{�Af��P&8>���ۃ[�����h�B$MIj���b^^<kz���dN�ս�4T�jD��k�������iݨ���g�����ewu��N�"�
'��'��|E�?8 Af�ҖH��b/]�<x0a�wUи�+W-�u�O�޴�A#����Q<����7��P�db4b��-wl�N�i��Nk�^f�mC"���z'�w���T�%�i�鋖��c�F]����Oy�����٘>�&�ll���yη]=�ݻZzW�B��Vկh��úT^8�^�H�����v�:�tlT;��Y1!�r�nF�2���;��o���l��ۇ���>6{	��/m�w�K�����lv��l��5��ۧȌ
�Z.@6�k����u\k��v�;'�{I�����\S�9�q\���]�qۂ�wC��ˤ��ƣ1�����Z@��PcF��q֫�pu�/i���a�	���T;v�S4hT�}�w�F����$R��Z@�Hu�łQ�sd�
���"�� �2����(2�$UI���E,�d�UM6�	 �O�WuY ��yȰ��,�g�Ψ�ԇ{��3TA�l�䛿�<�t��;�$��K*$�w��Ou��͂|�3Q�EA�5DMEy�f��#T��$��dNl�'���D����q��	�Fv�к�b��4�֫����_>ʿ��Qn.4Xcm�I��sd��9�`�S�9r�����p�|s�pq��<���l��qש�v5����]��7���񵉒�.�W����߽l��5$Lp,�r,��G��z�&3*y�]�4�z�����S�5	|bڲ��	����DE�k.k�<������Ι�k�y��z�vna{�Uy*k�85A�4!m5��p�4^�q�j_Y�r���]r����=9iz�=�=�g6~$�tOt���SԼH%�ybj��C��g.��(�B��31B͔���<��I%��dTvylܢN�� ���"Fod�f��SUU1)G��b���"h��D��e�@��ݴ	$z�c���(�q�eb�	�����4$Lצ����$�H$;}u��hT�Y���߉v�m	����)dm�renFU{6��e�F'�4L�cC�z=\�L�mƛ��2�Ct_q��hM?r�~�CD�����$��}6c���+��)/�^�ډ�WC	Iʑ�D��]uC�m�3d=8���Q�VWj^$��`�ꯥ)��I�م���}��51SP$R@^�4 ���$�W�#�����������;��L��yfI��qW^Bx4������u�jn며̨c�k�ۢه���������  n�OĒ7k� H$>����Y2�*fb��+��z�\��� �Z�v�$so��AQ=���u<��E�Y>繉 K}�ə������H\��d�̷ti��1c��N�X�$�ݺ�1�:	ja̘�Ю���'�
�/n7G0�gn�&mbNܜ�I���a�ܧ�Z�f��?ϫ����?{���$$=��Y �TOl�y{wq��u/��d1�p��0b�ɓIx��,Q�.)�[��z���	٭��>$5۫ ���� �r�o�i�����f�f�sI@j�Ӊ1���x���4>]]�7�U���	$����%L����a�K��%'wۛo9�5�d��s3�>"�w�>!�gE�|OvjF�Y�Z_�c�DED1�f���Y۴tɰ���>����^��6���o���3YrH�"�y��ꢩ��i�K�f>���đm�Ȣe@�H���8���I'��x����IJ��>ɜزJ��V]�)9����1�8܅ ��u��sprɆ�d�w��7c�۵n���9�5�a�{��S/�2�-�;�en:Il���C��kŽ[���>#���$��u��.O�7�-:���N��0�¶;�3PJ�I��݋ ���ԑ>J)�n�nJ���md^R���06�ɫ�,��I\�Z���s�7Q��\�v>qKd�+�
7ݗv��C��a)935g�u�DX��}�e��D�n5ؓ�A+sR�g\Ð���&�;J��a�K��%'W��w	D%�{�]&\��x�U�n� ��/b�8�Ă;��]{҈�<)t�9p�3Z'���F����G��m1��z�hDxF��K�||��~��AN�n*KL5vz�RG���^Em��g��B������Nd��񻇘������;-�[��`Cڝ_wNa:�R�xC��S����!w�;;8������8��o[��OK��r�v�!	��k�y�r�(M���S��`z�TM��%���J ��]�sh��Guf�mP�a�Y<"�Y,Y�`�B5�Q�Aw��gf�S����^{�P�}��8G�Gᣜ��G׳���A�L;Ҏ��J&�7�]�kKx�3�^�t�����XF�,:��BEd*9!�x7w��OV�
S����`&��v��)RVh���\��yS:�<���{���JZx���e�wҬ��ۋo|����w-�:��*V��$�!8o�Q�K�U���ƭF��7�(�ĎS���{�U˳^@Gr7��j\O[���ի�����&	��O���ޏ����3O�����ߘuإT��BR�p�,�����"���%�P&d�H�l��jN1�HP�w�<"�(����liu�xMk=��zd�[I�w��YZĥN�� X"r"�T��r��D�a�{y9t�~���A�"�����*��Łr1T=��gy�X�]��3#��e�}�T�4����Vv�Uvr�X�x���=�Y���\�2!���j��&*Z��9�j%��o���!��E��5��c�i��[����<�MY����۴����!7M�`�GP�H0`�U�U�T�Qeh�mPQKj*�PAFT�ĭ�l���m)hUA-F�h��j�jҕ���!QbU�TQJ�Ub,m��Z�V�
�(��ڢ�F�1cDm�T��* ��X��Db�l��UED@b�iER���*�і��Ҋ�V؍X���iF�Kb�UʌUQ����dV,lj	Qe`����Ĩ���mE��)j�j5����l*�X�F��E+X��1��Z5����b�%cR�`���b�jT��%�Q��"��l�ee[
���kDb"�[+m�j*��*����m�dYm�*Ŵ�QJ�X�H��%�ڍ[YE��c*�AY[Yb֨��Q��"��V���-�*��Q�*,b�A�*�U*5�TQ�%ʣQ
�E,��EJ�R�b0E�֥ZU�T+Ym��*�#���E��*(�XV��ԬE��TX����*�%j��R�J���j������GN�������`��ܓ��Ǝ�1��{]d�.So�7\mM�|�֞ƌo	q@m�!��G�u��2F܉��gv�8ݞ���ԯ�����ۮ�ݹܤ�:�e��P�Xv��Y6�s��^y��k>3�dy�rP���Y���9{q��G6��B��ln����xdn�2K��6z��{�O]�X\��=s�5��G��C���vݎ1z��{M�PSV�*κr�ݏkE�S1����{Pݎ���st���u��9u���5��:���{&<s�-�g���ΞL��7զ��\�6�]��ְ�8v.�=�ŻI{�����V�Z80:�vǲ�cnexuu�n�\��N�۳�������E���W&�c�lC��c�]^���X�Ns��Es�XCK�I�<H鹘�����G6y��Ӷݻ6��.�J��pɴ�j���F�]�nI�kp�}i9{Q�ݢ��0�x��:v6@��.ݮk�=�������@<��4����Ӹ��;��n��3���L��wX�Rl쫨�n���c{<i�V�\ew������@���DY��7t"W�32�ݞ����ᘺ"�#����蓶{"�m���-%J���y�C���ڭ��\؃O�{�۞��e����x{��x�q�q6q�s�ڱ�b1%��d�,�y�=��0k<˓ѝ��W��k� ���us�[�fۭ��SD.rμ��
�gn��s�,l���9sv:���v�Ŕp Q�7l��j۳���F'c��`��Ѷm:��6թ�۶��3�c��/L�G��$�z�z�9��g`Z�l���b�J���%{M�݋Iλp=rbV��khn��OG����d�3�Á��>�R�W�]��);i��ܯcsv��b�#�n\n�p�xP,vU�B�/m�ދ�\5�[mQ�po8��9����\�&�hy뭴�a�ϭɓ�Q�ܳ��9�#Z��[d�5�ӚˣY�@ \�n�F����mg`�sN�<9�lJFB��7��qs=Z�=�;�&�nm�wD��j��A�3���|�u�n�a�s�N����d����9�����.��P�A1ۇ���mӓs�q֞Σ��y��]��=���d|]�n���!���q]��p�nw��]�Si�Azc2\�<�=3���p�����X�Za���<�S+��f��xβ�m�Y3�����mWn�L� \��m�.�Z5����3�4""EL�I� ۆ���ƭxI��Ϋ6F����d�ŒOfrH�3]�
e�$�6䛸P����Վd߭���lnC$�y�"	��,<�x��l8F�����jI��MER��j�	)���x���>*w_U/�/�`@Ҙr�R��ˬ��sզ�
~ڝ��A�N��vg�;��� o'��\(���D.�AT��LI5&b��L�"����>&9��t0!Z�_]�$T�H/F����Ol�4��1>���==�A	h�?�I	)�9�WQ��F�Bz|�yݹ�:ɰM�\�����߯[�;P�[�^�i ����'b{f�A�+d���!��D�@8y;�wM�g	��p+V���q���6��^탵�z��/�	λU	d7����lfi�ۃ��]��x�������=�S~���w78��ՉDP��m�l�s����@&��w��E�~�����ϼ�q��6zڐ�ݲF>�@�צ&�*�bR��ۓ�Gn�Cb���u�p*"��-�$��1؟dOl�F; T�^��=W�qI�	mr�	;P��O�Ot߉��S8����#�E��؂"��SQ&M$g3.����"�LX{p����ANl	�ԍ�U��ݚouC�%),n%�"e
z,v���vζ�q�b7!Z�����r�$�w��}����35dV�g	>#S��$��Hͱ��P�1��&P�:�{K��
X�I��ݭ�K�ܦ�����I���I[N��H�ԉ��PnxY���Q��
'�8ÙnO�{r�$���E� �{�P���NDnu�ݝ��X&������m�����2�KT�w���[��JjT�f�����6e�c'3�կ�g�<M���_x� D���
Y��|�]��]����	��Ilm�7B�71�Fdåuc1����P�/s컄�JqZ����R�L	,n�W�>&�b}&M<�H	 �NH���u�����$����� ����l��˟�������7���(të:�x%y�S�C�7@[s۠���v�׷Q�i�������h+�D���3,Y<��^ �;��Y[��˹�ڶ���Š�:��z�&bJbjdMLD��+1Z�(�����D�'`hMR�I�I�#:������c�6�M�����aw0�K�);��v���BK����N��1�����1t�H{OR$�_��¡J^p!�%�)R�mǔ���m@[D<�V����*:�zOL�G��ݯ�g��#�����c��¼�Z��_�Z��(���ǭR�%}���3���[:3r�Y��ק� ���>�����{B�k�3U5U16��nO�,�s5!l�Gg	����^��J�y5�����-o�&\��jCV9.�C�]J��l��Y����A��T>#�ڐ7\8o8�M��TQ�Đ$���	!GV͕y�!��3M�Hw������X���Q5Bjdɤ�Y�ˢ�Ϯ��u�*�4ܥcH!�ۋ���f�&�?o�������Ƞ�-K�Rէٷs�Y�����L�F�v=�~!B�T��Z�P��.�)`6�'v/���_H��K��� IIΛ���f� �V�ո�Qyn:a300p����y�b�Է%*YIv�ʏC�NN����� �u�lY]t�%�n���O�9T$�Ŋ�!�i���v������K�o��3+�aq���Q]��U�Ӥw�~ zl<�܋|RX�d6/�.�_�����磘���i�MZ�&P�:��m��9�7��
�=g/GGc�hp�78��:{Po����m�UwNa�qY��W;p����|d�<o/�v���vln898x�l��ra����lV��{,�§;�q�ͩw���e+;ϗ\k�Z�y��`�x�v;t[��|g���s��{��<y�����;̓N�`X� �,��ҭ�]��n�!�\�s�����얞֡8L�����&u���������v�j�bW���ې@<];@$�պ��cg�&{�y�A'�+�h�ӑ&""���TQ�ŉ�3U���D�zO�$lel�>���D���R��c�Y��o��`�D�	��&��fX�	*y�I&�S�)ۋ��F�Yle9�<N�f]����Cs09D�i��|=ێ��b��s
���;nl��ݴI>=�o3_oE����a�ɨ����ۗ#D���6���E���gtŜ�
����6I>�oR$���MF!3V�k��S�4��::��G=1q��y��E[��v���3�[������������Ѵ0ӿO��v(�彴	��n/�qE.<Һb�aWM�F�=H��Q5L��MI�G�ܐE����-!N�c\�}�mR}������Vn�����f^Njj�^+��-�bYy|�E@qFS��%b",۹�Ih�����w3_�{�����}@���ׁǾ�q��9..�1���ю��"+�QF�,I|s�݉ �<r�;z�r4��ԉ��n����B�Lq-ʔ��[�ާ'���';U��_%�\TB�}/B�z�;OR��{��V纽	}Cx�$Q-������H �E;��Gc5v�1Gז�|y��$.�q`�Ȃ��k_,�!�}? ����]Kj[�j���n����v8�F^s��M�!J�d����wݭ�cH�N�*�5 I>/���H�M8�r
�u�ɾ���W���(]�mJ��E�CI��Qx�<�����y_�_΀ ��� ���N,�,��n.�1k]��ד���*Y.\���3�?n�k�Q	)]����W��j�0v�V�ra��Ln�@k�~���#��η�����兵�w��T�uס��w�?�	!�#�D˚U�vg�<<=�%[�>������q~'w0$��^��7د�0hnDA��	%d�Œs۶y���{�|���TJȷ䣡6���;�]�ޯ���ʴ�،��ȝk��H$.�p/Ĺ�ԌT�wH���c���U{��v���t��{Am����g����b钚�j+��~�����Lաx�[�$�����Ԉ�z�Ყuǳ�n/�	�����&�Lɒfhi+\�@�.D`q��Er��N���!�n��jwZy�!��]d����T�4(��5Sl�s`����'Ă���U��U���œ�r:�l�	�On��}��u2Y$K%˕7������rӭt��&��آH�oR���-�=<Һ��>����̫6_o{��űa�s���v�kN/�N͚��L��6NgUF�X��+5Z�s!�[�Y�j���xzF�}�����}s�B`ת���Wx	�'�p)uAw=��l�O�s�iB�����Ȫ]�/UW9�R��H[�r��<��z�:�0���KuUí�={pnY:���!�Tf�EI�Y��̺\��$	��_uEF�!E9D��m��$�we����$$n\�3P��Ң�yF]_td�!BoVX$��jD�_E�� 7��^��������$	n5k�w4�;�n�[��q�ކE���A"5� �bQ�HEI�B��U1d_gh�ʻ���NvwX@}�6�X$���[z�n]Hג��$'٩���S4f�MMI��k��>$����P7�N�$T�����[�� ���:�{ۯT]ƶ�٥�'�)[&=�fj�년�w���r�z�G}e���{A�����}�sw�����py�x���@��Wҙ�����\����������a�3ێ*x㥃mm������nN�{i�ޯ0u��lm{�.y�x��*��7Pi�%]��{Uu>����X�T{q�q��ό�����E��c7U��$�[ K�ބֲ��j�q�N ��lܱi�ʤ��8��B�ˡҏk�Ϸ�m���$j3�1�7!{�g���M5�ev����E獬�%n�6�ϧh-��v�q[�FS�li��C���<��/UE���%�H{�$B����N:8lt�E��K��-Ō�$�3F[C�ڍ�����UmN/�mj_(��d�
��1�N-�"�e&L�C�) q.\���D.���|��>qP�������Q$��������7��fL�3@�V��օ��{{5ԬQZ ��$������L>�HR�Nn��"����|V�]Ùڅ.%�)Eo��ω1��c�7z��&�'�WE�><�а	�wn��\X�=�� E#֥�\ �ga���^���n��7q$5�ʆh�r�����*%��S;��_L%ӻ$�!���n0v6���ޘq��-�U�Fa�g�(ꨢ���r��NU���r�wRkF<i�[��qe |�����؟P�là�����k9ٰؖ�S��?M��mo���,�ё;�2�k���{�xxj���$��V	'��n��O �6�d*�ur@�Z$Έ�3Tb�DR@���� ����3ᴨ�ꗮŞ�u~2��`Lښ_%�e�%C6����ēK��������.���	�7b� ��R�$��鐦z::�c��x鄶l/I�&bI��A�V۶	$�s��jN��|H���$usԁ �{�~4���!�l�䟷%�5}���anW�ez-�]]Þ���5����:5��w�Õ څ.%�;�K3i�Is�ʸP�t[��X�`��UՓ�B��H��%�$MD�Q�H�{~�p�A����89;�>'ć/u"A�n��A<�Χ3s\R�%a�g�(ꨣ}�^$�{b��I'�Ao�y��R�F���r�"���rF���O�>z�ذ{5b�ykp�4����8��CYNy����)�sӌ٣V�ǷZg�O\S�ږP3f��v@�G�H�v��ɡ�{��-�;������"E�e1��!n����g����U�[������LM�yh��Ho;�V�uU�Xم���M,sfeޤ��80)p����`@S1:�êǐ�4�eD'unˑ��}���I�����	�mW��h�3���	|8����1-��Y�5j���y`hbZ�7|���q�����v�{��j�����9α�p���d�3hJ�՗%v��y�>G�l��
�㛣�ӯ�U�t����U�£���VI5����s�7!�(M3�IzI��I��N��.1)�y�bژp�t�I'kX!��z��l�ݐ[� u��{�c���g��o������,��򽉋<�pi��GPʑ�<��[�S��;L���G.Wh�=�8���a�����;�D��V"���"|���Zg�����Ϋ�d�^�}�_D7g�i�Gcq�U1�f�����q�/cZ��F�e��)�7���a���
�;j���"rq;�ߝJ��NE9�8�z���n��J�T�"���y�'��B��sF�.�S�t��^#�o�>�Ms|$��]�R�U�szv+w4�Mp����]����S(�݆z��y��� ��7��d��;�֡��=������xdfj���v5�ה�{�0��a�G�|�"��[
 �UY[mEY[**��J��
Z[*(1U�H��b*���*�E�

[AVT��jZ-P�Ub�+*�"F1���2�*�"DU"���AV*��"�Ub��",�R��D��TF1"��-�UQZ�b��*+�*%�D��em���,Q���YZł1��kF�e�cmERZ�QB��@�T#"
��DX�$U#�1ڂ�m*�DjE��[j��X�Ԣ*�QEUQDADj���KlZEDD,EҬATc"*"���%b"��[eKj����*Q*F�-�R�iV�Qm����E�X�-l�*"�VJZ(��Q�(�km",��@Z�Tb�V�m��T1+(��UcZ5*���[l*1Qkc ��P�-�±T`�
��(����T�Z��R���F	hF�ڢ�(��b�حK���-��%eb���Q� �EQ"#"[J��VY�! ��y�|������@��E���w�xLњ��"�!�e���>C����$��6����곑9>���z�/���v���EJ!6�s.$�:�;�F�b��6 1Qi�3��[v���'�:�٘��a�s�(�#�W�n�\�n�r�!1���l�t��u�:�Ne�����-�����L���
��.���Aދw$��No�ii�5���i[Sk��9R���ܕ��٥f
��®]�� �y͸�AG�͂|n��'�;g��̽ �϶D�"�����3)�{~�	�eӱ@�d�峽�|I��Ă (�sd�3"��
�TQ��Ħڊ�ݻr�܌ͼ$��;b���0>�~��E��Ml�ȣ�ꆕ���Ҽݒ�ŭ"������Ê�$�o���>r���y����럖��{pr�#Q�l������H;�X��?D�5QE$̿Q��~�Gk	�TX���N� H���|Iܭ�ӝ���d���UW����|��+��I/)��u���]�K�<k� ۳n��LN��ħ)'��F�!6��r��[e�D�{���(���ݗp�x���P��#!%���A�
���L�iB������^����.��\2A>�uX$�;R$����w�u��m�TL��R�nN�Evu� ��{k��Q8#��i��ZP��<t�"���,�ٕ����n��Fz;{��1���˲I1��y ~3�(�?/ &S>� ���c���B�Um.Đ�lc�L*��E�"�O�y�D���ӇV��窡T}�E�$]Ȭ��hE�iu�kDJ�H�Cv~/�W��{/���^n)�3&6��a�����EL/�� A��z^-2�nf�j�X4�#��c����n;���c��k���c�{�/`%5˷5�B�:��|���V��rz9�/ �M�� �6k�;�֭�T��wmg���V\>y�1�{@�0���ذ���i�bF�Q�q�nT{�]��:K5�[��S�Y�\-�QN�l`ۍ��/a�=\/�u1�v$:9�+��4�]m���y���F��u��D�Jh�&��Y㋞��u��N�ЛG]��}\�:�������{�I�덩��2ŒLwn�^ �ӎ=Z.�����Q
��J(�6
�j[�2K�-ܓ�\_olWa���Y�&9���]Ƕ�~�뼩�֪G�����OH&Q ͡}���w��$���S\���	��^'ėю���	�1@�p7%B��s-�#3s�h��Ng]_�'ď=�����]IvY������jG9���EQQ5Tfm=�$k�wϱD�D4|	�W�A�w ��n7ϟ�7����Y�lXK�Tscu�+:͝��n�G��׬1�X�w�xx�}��}��@ЯUE
�$�$��	ܟ	=��`���Ys�y�ے�D�b^'���#�֠�r���������P�ul�z]Q�Ƿ��c*�8u�Rg��뙘;����57�f���rp��o������C���8,��n�eFL���1s�jqS׊ޱߞ  <'������?dX>__U����miy3õv�M"�$ږ�̄�Q�y%��Jٕ�3�k"��j.��N�<�~$����Q`!�R]�׹��M缵K���3z�Nu�\O��>p��5F�׳�D��|�2$G�����+P�O_��Id�eZ��Û�(���g�LԾ����#6�Y'�;m�bK�{$X�k��>}��{gsעܛ]q��nbz(���;b]���M͹~��zSL�d�d����
!}�[Qd�ӝ�:�4T�g�fT��z�X'A��$ЯUE��$#�7og�5�S��/I����9ڐ$���'��KӲ����Pl9NF�p���v��=/v� ��L��k'c���R�j�U��x��C�f�H0f��~I��68��ɛ��klt�Qx����/۶�%�Њ"m���~��8n����W��}��{�Z��$__�~$�t�ڑT1���-���٪��T�LV\t(� �rq�@�_t��r�:���D��Ӥ{Ћ,d!�JJ���ۿ�#9�X���u��A۬��'Ď��A I}Ӗ#�!����[�2`��MC��1�������oS�ְhי���;�s�!^[�6"D�Mf�MI��nŐH;:��� ��7�>ر�)ܗ��� �{��#;NU��L�D�F{%�-޺�h�O*�E�H:�"I��\�{jQ/q8���ʞU���P��"`תb�;����K��o���oZq.������2^�D��/�FW0�I����"� ���bګ�&�2�{;2�$Ot�E��J�u)�r��5�l�ds�5�ڵ���fȞ��5��m�N+-Z��!�����Q�r��5*i����ѝ�OE�yT�ND���B��I&�u����
����R�ӭ\֛so�9XI ����nGndvr����e,�w2�"A'vX!u���혍렲��5:��0r7,i�6��X����=�n�ͳW`�k]���tuV�ֺ�?�ϼo�}�]�0���H�I·�� �J���6��G8��Q�om���o�T^Iu*Bk�hLԛ_g]�n�:�[9ٶ� ��{"� ���`�cg��H�^�-'���R�jY2�3pq{��Jn��B��]Auę5����'v_�Į��8�D�5�^��7�k�3Y0
ï��&\Z�I$���X$�C��и�pB=��D��^FC��nG�(�{�IAۙVWLWdJ����vp�qł|IYn��y�h�t:��2��pbڲT÷�'6�n3�*j�/&aV�򦻮����GU	�Z��%HR�5���l��F- l�y���>�@���<+��̭�nc��r��; Y���x�÷[��
K��f��vs���N��kn��h������*��묮C`C��5�m����B1ؒ ݍ�:ڛ�y�c�d�ͷ���v;p�"li�c���nF���Q��{1�����m�n�N+sFw;k>�cR��ctn��������^�h���u�=�
���v5���G�d�*G#��Aiy��\����wW!\Wmm/m=�A���5�%�nh����}�MA��m��m�u0�{k�)%���K��c��-�v\e2��ă�|�c���7`*�L�7	Iw]��i#vN��TK��~#]�Y �#������N�,Y�v�ҽ�]Dʐ��#��E�;��I���D�AQN�����
��I}�vU�,��}�ܒ�S5p��Sp]`j��wo��Ԯρ��^'�7��b���|DqT�.�@̈����i:;_����O�ć!|7e{��U���"|Gt<�Ha���N�����/������<�3�^;z�ؙt�nf1�b���i��!"T�CgFpt9NF1�����>"9��>/��
��3YQ�ָ����J������:�4Clj\1M.�n�T+�9/v��Oy7�_��
vܽ��s��S�5�U�T��&f�λ��I��?����_bu]z��}��c�pqI�-:�Ûg��$�Y�@���I�w��iF_}�8�?}v��̔^H�j&)l�'�<�����B�^��ב·�� ��ޙ��C�=�S���mx'�\��
�ɘ���3,=�Ok���1�ėz��$_OdX$�������*2��I��#{ONj�MT���3ю�'Ă˷b�8��+�� 7y�A>/c��J���N��WP���.j�	�H!7$���yu��-qnw��2[�7=��^��O�~�k��k���n�	|�utҸxdm8�l�>��$�Y�z�}�X��#%��A��
 Ξ@`�7�>Z���$��^E�I
:�lI������W섓��P���p�1�mJ�WS$�P+��Qn/W�8�M���8;n{��as��^ƾ���蔧�����?6�0�]�+�rȚ�J=��,}(�f���sf�9DmU{{� WJ��	|�x�꟔Y��in�B�����8���E�Vǉ �E+��O��E=��!�j�М#'��wdo��V$��x�X��Gq�:�z �W�(��Ȝ��𙹥Fnl�H����퓐A���?��Z�5��L��Z�f~� qb�㕽=��Nܽ�n��ڔ�c4O8�+o������Ϋ�L����$�i��&;;lR���B���bG�ŀ���LfE�>+�~t>����	��C����Ŀ#<f�f�wM�I������u;�A�Q9�e���r')���U]ϡ(�v�U��af�`z�&f�%=٨J7ݗ(u���-����]g]�Zx�������3��!gm���xX�׳3�^hv��;��&}���5���_o�ʕ{�7�ǚJ�}��kc{s�N4e���Sx`�&����.�[X��ۺ�����y{��ﾛ$wQ�2�13S"���]��	>��$)�2m�fWJ$���%�P^v]�P���Ly��9vOl�"dh����p�`i�6{r[��.�����65h-|��￼��4&b�g[� �cw��$�/"�Ɋ�Y���Y���1H�fU��ų�H1�nd���w$��v"��iF��	1��aC�&�E:;&���$�#�1�^5mR��'�X��3�侧W��[�(O�7�>���#8b���@�	�-^���6��ݛ��G���$/��Y%��s+.L5�ƒ�ײGm��7���$-ӡni<Ϝg�_X��QHXE��1H��u�A'�X�AG�����!�=dժ�k��8J�ߋ��F�q��o���9�L]9�d���z��J�!���7���x�R=�N��$�}O�4�tb���LO �DC䳏{�gg{�4����(J�Y��GZ�R����U:Y��Lx�G�O%�&�}qz'ѿb+;��C7�F�@��ó�F��OU�1N��f�םg�B�4�A��4w��y��[���j�����'���gK)�ru�4A�ʂ)
���4�I���q9H�ċ�໥D(*c,O�5L��[l�8�
���<��u�zCp��5�	��-��X����NN���Ӊ���·
"������{_�~^4S���Oy���@"gE�&������������R�y�_�Y��ڇ�w��azf�|�p d��>�]ѡn��h�\�9<�N��.`�Fl�A���۪T�D7�:}X��v$��HM7ǖ��yc?6DOL��\���]��c�A��'f`C*�6a����eͦ{��x�4J�'�˥�"=Va�0A��_��K���0�e�yx�ٓ��z�Ӿ�FW<���R՜}�(�Ȥ���(�V_E�K�0#�����5�g[t�Y�b��z+�J��]g�������ǡ{������7��Mb$
��{.�98���G���(W��qw-�1~��i��[����۱vר���jW���G���vbTet�Q;��Ƕ���?G'g2�V3�&L뛽�{\.!����,<�Ө@�!dVp�f�N�5eWwf�e����E�"��J�"��PPX�DV�)�
�Im�h�Q
5X��*E*�"B�b�J�UPX���R�e� �b��ڲ��U�T�#"��EP�mJ� TQAH���H�ʲ����QEb���QX)iV"����*����ҕQD*TTU���R��Qml����Q�iQ�R"E�mB���QkF,QdU�""�+�+�jȨ,TH�YJ�R��Z��	l����E�V�Q"�*ʔV*����[
�J�b���+DbEm�V�F�DQ��bֲ�E��E+X���TD�F*��b�j�TkDETA-�l�­,+(�[QEQB�+�6�eQ�V((�(�U��e(�c�QbQ*�ЩX�DTA@FV��T*�UUX�b�P����"�b�mJ��m��
��~��O8l�는�ǁn��_����WϚ��m�O��'gbc7.��ζ3���u�-���^�T�m��m,�볷�w-�D�y[#�@��9���mv!��>�j�M�"S��������q���j���;5r���(>}��m����2�j�n^r"�q�N@�e�i�^竞�V0<�OU�I��nS�!]`뗝�-<j�u�W-�q=72ۮ��j�e���c*�m�s���Ľ��ƻK�]9�Η�����^Q��|����]��[[�/oc]�^ڃ�i�eڹy�=�:�o<b�mت�Z^꽪z�';o*��6��xM�����]�N����g���#ۍ�l�x�r�]��\��!��q5��q����^r�msU7,�ű�x��.�Q�ĝ�,�����u�;CdmmK�ض��g`�z:t�E������N{8���l|���ϓ@h���,�ͣ5u���m�Af�{� on���c��{rOvϧ�����|���:���iA����q�\�t�p>��2n�Gm�A1��=��Q��:L�6w�������]j���5�a�0Ʈ���!�x|e��A<��ۮ��U�́4Fp�>�ɻ0�r�95���M�&�R��6-��lps3oN���ny� g���k�E�X�{b6���p<>��q�����ҳ���M����A��v�9�Ǯ�n�g�����ú0`�z;[g�zy��sn��^�B��j6ۓmlq�- ,�ݎѲɗ��'i,X�uW��:����Lݗ��]l��:�m�n���9�	�U�p���s=c�\��l���4�ɳ��x:"�b'��T�ܧu��o��K��c�;]�z�rF�n.Kt�2��#ӛ�	]Ƭ<��z�9��t�z��ؘ8��ٻ\%�F�n�(����׷nol½%d�M��!M�0d���@�ǎ�Dˬ�sڸݷ�>�䱻^�3g�����H�d*��im��XW����&�َҜ`�0]����cs�ݦ�Ɗl��	77�)�\rZ��WY���l�C�M��<s��Ht^�O�;��2v�.�Ŷӻ"y��g9�vѶ�1�9�8NQ��������ʧ�-�+,j�ۊ����u�q�����6��vLj�컨�t΋k��olv�x�ѫ�x'gY���V-�!vX���6ǐ%��ۅ��ոõfN^ݹ�ۇ��v�ݺ��\�v�rջ�?_,jT�*�[���2�νq��#��ld�����ebG]bJ�������l��	3�/�y	9�����H
:�D���k��u�^$����[�Lk�Rf"��g�����f����� �y�dX$���$ttM*sQ;D�[���.N	1DS&e�OD�	,�wDy]�*���[�� ���bA�gWO��Y�)'�%���MuQ�\Ľ\��ي��$�}���,�C�յH��V%Oڒ�3d]A��LI�.�j�e�$�m�M��֮�Ep$+��`�|��M��O��jDdvB���m���c!�z���y�nM�����r���GH��[y(CP���~Y���i[�����|����̀O��<�HB�p��a<� �FG[��T�""f�E	3����lc����s�eM�;tD���H˕�3�rM��7��-���/�(^�f�s��&��ř�V���]�N�B\�[���1� �GC��������O��+�emBTy� ��rH8�K���H�ܫ�$�����USۯJ �e���>�H��.N�1DR&e �K��;��h���%�J�@��ԉ$�9��j�1��R:�� �Gx�O�Mx�Q�I�$������B:�+�>��S`�f��A/����\w�������S�E�b��,<-�{ۋ�wk�۵����ϧ��Q�?;��߽c�[�[����ɲ!�m�I/��`ڀsv�{�U[��y1H�̫��S��C�KR�q"�]{*����>�&2��텆�pQ� v�	$�U� �\B��q�vDe����"%11U"����{���I9ʸ$�Vj�F��ω�"n��<�E��-�{U�m��1S�_^3^�F
����	L6b��}���/��FI��y����2��=���yÊ�~��^yo6ar�^���hY���3:��2�@S��wZ�>$@�u��%G_H�6��b�˖�ƻ��/k���(�Bjd̤g�]��˷/z�О��˒ro9 H'�{�,�K賫��{2k/܋T�s=����m{]nL�؝���	�mtv{A�\��m��f(���/� ���<,H/���,A�B���8�kPꋵ٩	��ӗ�G
�*E@4fi"�f]FIpdJB��U]���3=v]�u��A>���d���� ��r�w)�x8V2�D���B����yuu|�,yS�-;�g�28��	
:�l���"R���ÉR]�����q���Jy^p�{g/�	v܋ �=ڢn�����@�Pʭ3�Mx�`S�y�����Ԡ�^���^:���_-�wf����ܼ�l���bܒ�#u:�ٝ��� ��U�:�)0f�S$гg��l����;۲3]���O]q��I򎽛�����M�w�ز���"'�Pc��L��Y���޴��3luœ�������n�=%�b�5&���g�]�>$.݊ S��^+V=��۳�Au�9�;~�|H���F`=�DA��7}x��&��:�oK�����l�HyשyD��K����rd�@�/��C9�B����x�ˢ	+��	��
�AU*WIrϰ8��	���H
��ъ147SK�f����m\oD%
מ_��I�uڂ��*�7��ՙ��2Cۣ1t*"MT�f/<73�^��r�Bʣ��wE�f�H��s`���mA>/�U�b�73f��^�qbe��m��!�������w�~�7��q~���=�W��ZM��2�,B��P'%ȯU����zw��*�)�)����w��=�����o89��5�ƺvݕݬ��i�����1Fͷ[ ���p�8�Cz7e^����"m����K���c��!��\�آ���:<v7���X���g\[����.�ݬd7�]��[�J8q�u�Mk86ǝ��۶����O]�.�śv3ю8�Wڟg[���/cuG]��En}��������Ś
���K�z<�nK]�܎��D�Q��y����Q[��${b������E�r��>������*�T���7b�$맶� �wu"'�܈���Y=���f���־�=��-_B�͠g�Y�t�#O$O��Q'���۩ ��W �U�f�z�9��g	/툀L�kƢ��]�"A>=�*�����1Tk�x^J�	1��g��U�/N!TSF�IVc�{V.�w��	%�l�_)
n��bѱ>1��V�B�I��X@�!LetנIB��X�O�ĭ:�m5�	�!�^�O��b�*;��z�쒫z7�ŖX�3c����[M����Hgc�p�طn��V��#�5c�.&v���}-��T�����|��r��J�� ȋ���&��';���^K�L�I�}3)?�wf5�0��#c��`��n/ܝu�O&X�ٽ�:X���Go��͢�Rx����o��3{�����Z�ў�K��tf�LBB� ��
�j�$�����T}�l�{�.��FGu+@�f���0fR{Y>��j�KќJ��L��[kI��U`��}7�N`<6"<g�^3mWbA��T;Jd�i�`�K��6	 �v퓉]�i� �<�'�厓BU�M �ڜ'��c�K��W���Ρd3��d����@�}���$���I�[!̲@���RK����(u���0��b�y�i�����ߥ��c�P0g�+u`�]6I C�ԍU��ûw�f�:P��{5	FmR����P��J�^�ws������@��VȲ@�ۨ/���zڽ���Ft�52`���&d���$�m�/��o5�]=�2�c��4���XLRW˼�m��9{��Z@װ�<�akz�'��Ps�Ș�+wil;���'�a�-���3W,|�E��q�t�1�n�^��o���*`̥�<��p����d��	���"I�}n��SX�ء~�WM��:	�>3��6<I@=���jNJ�N��o�`��r,@��ԼI'��X�<�Gd�}���|�ΞM��wW'7n����Ks�z�o8�Ӵ�6'����H�,P���)��pB���T���1���$��݋1�׫s��*S$����T�0`ؠn&�uֺ�&Tcx�a��i��I�� O�=ծ�P�Q���OO(�����-�l�]E31j�6�>$�_P�I�*Vx����t��"s�R�K�u`��aEDUL�4,���/ft�\�*v갓K��Av�X�A>P�䌙f�%5[�tԨֶ��:�mX��&���H�y���ڼ���ߔ�a�	쟙���y�P�%�h�vQ��Azh�0sI]��]�1���H��oϷ�}���y5t��֩�H��hX>z���7��`�WvZ�\�B��^�:O����y�]!J:�89�Pqt�ren7g��ϡ��me��a �����kK�z��k�b���/H/o��I$���=�^����+v�� ��ug�厓BU(�Z!�eI�7�s�ne��I#�݋�>$��VH5QU��2����Պ)�R`�ؠ�_,�ڲA>#]�&�ι]�Q�v/�r��
�W:_%{��,���.Y��8S2]�cjl���mm�ү�6�Y��u`�}�p;+�{�0H����aA��T�3$в/��I��A����;������H�۩���M%=�$�49����*s��KSu��>�9z;�2LL7񺨝��a�~�"�Ѡ����I&E�* �`auzh��J�7��~���E�pW-�j��L��1{Y��ظ�m�YC�fj���㵋�U���V;�ud:9�]��:�6�rQ�g=Ri��q������[��Pv��ƶ���7>�������5�ώ�8yWs�h��V�U�Xۘ5�*�{kn#f�"S����9Ӻ�c�=rݣ��f�fۃf6�SP�#a�=�k'!]�z�n5�]^�W����?-���${N
Wñv�@r��N9Y�]����(�[�r�Oέ�����޷[T��3/�:���z�Ő	�5ݺ�8��5b3.@7�����]Y �=� Ϧ�f(��bH��Ʃk��ʙ �Ff�Y$���R"���s<*�U�h$f���hA�� ���#�2ŐI�Ƕ'���as����V	��f\\*q�BI��	p5���v;�Bq��-D�.�U�I�u/	���jZLUU�}�A��V	��J*jj=UF���K��KĒu�Xs.�cw^��3B�U%VI5��"|	��Q�k�S�ӕ%��0�?���{mv������[�[ہ���zћ���:���m��Ͽ���q�fI��^k�$��{h|{�ז9��fM�b��ɭ� �s�KČx������lS7)��P��U;�{{"D��̽������~�m�Sr��d#�}��z�-�����[ ���u�^;�H
�����:��R#��c�,�s ̛؋� xK3��mA���A8�l�ۋ��#u���9� h}5�1F�<I|Gm�_� ��y�Rn꬟vn��!������bj	1F)"���Ȼ����Zտ	%��	$�+jV�Y�?vv�D��f�U"�h@��}C<I=�y��$��-˚rY>��h"|[�W�A'�Os�,�R����~A�3�$B��N�l�Z����tfH���t8q�5j뵮y�3������j=UF�����ܼ�u�X��AS�B�٦��5�|�$u��H[6��neD�N!�sϗIʱ��D�g��B$=��~'ĕ=�~#_Rؖ��*��$���!��ئn�<JQ��U
����t)r$����ؘ΋�j]�8��h+�{fsA���=�h̖ȁ����*;��s|ϸ1�e7��{r�C�ٓ"3��u3'<U�ش��5�K����-�6O���ޞg �F��e���p����������=���٬Ơ�����Ű��o{(�썺��f%z�m87������y�[���1#�|8���{��]��-{|"�p�Ŝ�V�]��Y�4S%�z0kUe;��y����X���.�wl�����ra�;�D~�}��{y�˓�
�՜��&��̼p%�={ڝ�<V<��jdӞQ�n��<���U�{��b�IF�d�4��F��.���|�6o,Eۺ) p�y��������u.}�Qȧ����ͼ���٫�=���\*���ׅ�;���'T��Y�/F����ۖ	3y`�uך�,��R����v���1ə)ÇǾ�.��=_uӞ�E��l���ó۾�v8��T�y%�˭�SS^Y���c��	X���B0Z*2.��u4@�ZC��lj7ĖV��٦BB"v+Ud��3L5�j����JT������ϩӽ�����s���p�ol>�	�̺��؉�x4_��C���ŇVy3�Z�$�+!����Y��}�֬�ޑ`���N�D���*�o�U�5�����U$)Q	���U�(�Y��bY���f���F�l�=���3f5���(��"_������Mb�@��#^�9r�e3����oرz���կ�:���V�L�^�w
(@ �
2Ъ�
�UdTX�Z5*
�U`�cb��-�A""J�E�X�KJ��kE*�5�

*�(�EX���[*TXŭPDQAV�ʋ+�"
%��k-("1����A��UE����X0Db�ImjV��$DE�-���6���Z�1Qb�B6X��ʂ�B��m��k
�T��UVAh���(4���Q�"��E���#bA���((#+E[F�F6�-�k(�kD�J�X��*U`�1B�D*�T#iU���*��"���)E-�*ڠ,�V"#mPQTE���(�*��*�U��4��1�b�5�����b+X�ҔDEc��FV�EJ�Ib�m���ʀ��E`��׾���U�����E�3���$@��k�b��WbF:ݺ,7 �j��>$�T�U�>ݾV�La ��� ��+�^11@���k*ȎǶ��Cw5K���ݿX$�v�D%�ݙp�reTǳ&�6�FJ1���d���g9z�瓎��y����s��<9(�￟�y�	��^�4���� �'��$�R���G��`�ܫ �Ar�Y#y%5��@��$/���>2�N=�q˭U9����H;9�~$�}��$��n�yǳ7�^{ԣrn�s	�Ȣe&,k���o=� ��(o;0':�H��D�;L1��Rj�̤��s�z&M��]u�dI�ڑ$�O����;���X��MX�X�l:yq��g}�ٸ�c{8���=/�t	MxB΂�Z�涳5������Ҝ�eeN���N�e_�<����Mx�Q�]���Й��94�(�(KX'Ĉ[��$y�U��ZZ����{�����=�%G���������6=gs�ٹ���Gg����72���ϧؼ.�i��t��<�I!��^O[�[:Ev�q�5�A��U���6rʲL����=B޶Ɗ���	�gn�	�%��A��Y�(���6a<�ZJ**j=UF�����6��$w�`De�Ms(�L���0��^ ���P�דT i`�e'������������ ��$�����w:����j}�_���Q݋�ğSb�B/z�|C���N��9ךN�sHHv���W�A��,��·�q���_L��{���&���q�"�m�^�:�.��r#����K.����F �������j//
�����	�H�栃f{���j!a�mn���u�`�\67�;7����q٬���m��>޸z6L5�ֹ���!{q��t���`�px޶YyLʝ��n+�G8�v7+ݫ�=O]�n��R�=�uSvJ3�j÷�/5\;m�//=q�N�uպ*���oa�^�X�+��d)��������۝�ӹ��OO72u�����Iݧ�:Īmqv�l�N�p��Y������x%�E��v���,Q2<�A�Mx�Q�VbHO;ud�I*��m�x��e�>3[د�#6�Y#��=F�fb�31���zϏQ�Z�LI6)o+��}b�+�3&��ީ���R�5$��D�`�YB��}�,�TJ�*��@�Gm�Y������kIEDUUQ�ff��sW����׮�p5�U��	W�����z�c�������׀fO&�:HA�`�O�ω1��׌-krt��K����'Ğյd��C�v�_)�������#��rE�����{@U�)��#Gnk���`����l"[�Y�%w̆Sb����k�����c��^5]��<o7"B��w�*�+~�أ�-|�ʙ��������U_N�q��B��E���p5a�-�R���z���J<��6���*���𽌒�hݛ�P՗���a�UN��8�"�t*t�Y�
՛��q>��mYC� I�׊^uh$hhgQ'#��G7p����H�vU���'�جzE>c	� �]V	1��� ۋ&��7	M.��p�hʁ_ؒ�ΨQ�#��@�{yS���ؒF�R�[�v0m|�N2����l(���%W�h�5�@q9�~$�!kԁ$v�j�o���w��DSAE#��!���hyi�q�@j������a�Z�"�k�|������
T��B���P�3w*҄��먯����*���K�&�N��'}Q�TML��es�I����@q��6̽tG�&37R��_�&v�+�5W����v0D׌��W|H$mU�H)����K#M�UDċ����Lq.�KAQs��@{��⫼7.eZ�%�'r�l�\��3��>�3��e`�3�.oN��9���"|Go*�8j«�S	����eVw�[�����A%�T/��r���R�pu��2N�� c��FG7㛸cޓX�㇗L�Q0�k�Q:	�U<H�H=ܪ���o�;��^]�m�����lƹ�;<�pIF4J3���s�����dfb5�BN�-�w%�9p�&Us�fݤF>Ud�I
9t�2�)'8���3����I([�n�K�n�r�J�:T{:�.ĭ��&ȥ���׈ �m<``w����2����T5&�7*f��׉%�-[{5
8�U��\]]��:��;�^�> (��~���"`���6�İ3���QGăݷV	$�����&;�W5ؚ��f�f��p����02�Yu|����B���8)����1ikQz3�>Zv��oM&�lN>��%��j�<w�$�7V
��0"f�2jmx��/�I1����$�Q� �v��b�����0����|"f�ssq�$��S���P2rOXٟ=g�ܨ듗�6,��g+����l�jgn=�E	��%���^��$�}`W����^=���[���u`�_H���U5�5B�EIHWci
1^sb�M>��$Te��>&;�R1�G;�WV�Y75��� �X)RF��T���_�`_��n��੾��Xm��P�ݙqq��NJh�6**LJF{X��ӏ��6O�Ҷ�~�>�P(���~��F�,jBȁ�ݗ`	ޢ�c�sz<�����p���R߽�5�+�3QˮS�'w���Ԃ�Y��S���{8�����e����_���_�R����aRR!RT�{�gR'c+%eO~���@3�D��[����>����q�:#�������N��n��h�C��H����	>˕����}�炘�5�^s7�.v0��73J+N�Njs�/T��sŞ������m�˺9����;&3q	.{k��(�<�w2l�X�n`Bm�k&��t��';kS�J'���ͪ�7V��v{mv�gK��\3��\�,k��zr]�t���[p��wg��d-ɹ:H�ruv��⩖ܯp�=��3۲6}FA��g�nsHdp玀��@f`k���Q�ݏ���j�3/gg��#��F���V��s�0��t�A��9:�!�w^+����>��a�bh��g�Xa����r;H)h����Δ�h��=���`).}���|㿼�9��3=���q��bJ��}���0�
����Jf��4�S�{��'�����^��g�~�i����~f�(ʁD�<���:��X�=���`r�
<	��;H���̤�wك*#54�F�u]��}�}��� VVJ��<���`(q%aXV~��;��~�ߝ����AI�!P3�>����T��FT��{���T��75�r�5k�Wf�×�>�w�}����p�T�%�)-Ϲ���!Z��)��{� �
� VQ;�s��L睼�w��^{�OP�J��~�gXv0�/ۼN�`�6����<��B��uTE����VJ����=���d�|�3�？�
��y���:��-�����ZA��jϹ�ᧃ��>��~r+���7�F�BLp�&b[�8lB`��s����z9��l���7==8
K�j������sp㯀���y�����d��﻽�T*J°�(w>�܆�paR;������}�~>by�����Y++%eO�{�������a�bh��g�:��o͇#�����ў��}�����*�`��$4�s��Rga�]�`���퇧^\T5�.��第�[��(�P�uw9o"�X��O/����k�6q �0+c������
q�+(�Ϲ�ᤂ�"J�.O�����Nv]���'��Ҡ�DMGU�4Ì*{߼�Â%B�R2���Ϸ2q� �g��sZ�T��}۶�YϽ>`v5�Z���}�w�9- Ф+D;�s��I9����֦�htEA@#�����6���?e�yU|L�d��eK����l�r3�����;��l:��I�3+�~�ݝd�9�2����|k����6�YY+*^k��6��^�y�{�����Z�[xm���q�o�����Y+02Ɏ���vw�&�I�]��3�쯶�z�߈��I�^�T�����3��y�͝f��C�`�f!��w�����D��q�&�]���s�l�N$HrBl��;n�q�t�y�q��m��L����x�sc����?�-[��9���
�Y+*_;�{��1&30�1���|����L�f2c�����wX��a�zH��8�Aw �.����S;�w�m����VW��=�gY��1��}�ѾԮT�����0���F���}$	>�靲%e��N���b]}�{��P�f3`��a���ì�%eI��1&8���g��e}����z~9����X�0�H��w�e&Lp�����hֱ4bkYì�N����;���%grɌɖLw��}��,�3I��&3�s��������*f��x�ԫ�'�Q�یJ��!'w��ǘm���s!�{F�jf��Nl�Η�vs=�>{�2�;�T���>Ͳ��1����ȟg����m��b��J���gXy�c���GI��:�ì��3���`�z�|�3�_<��bMG��e��w���Ζq�2�d��LroϽ����'�2b`�&3&S>��6�_�?yw��c+%ea�߿l�6�	1��ϸw-փ5��]�g+�{�:��<f31��YR>_]�|����[��VzO��2$�O��s��:ͲVVJʓ�;��}��'��c%�Y���bg��{��&2c�sߺw<��͹};��X��26y;l���Z9�V��Z���:ݰ�.Sbd����B&F�I(?E/���0���ݝN�1�d�d2Ɏ���vw�d����Lf&g�����Y+*k��7���i��>��vq�d��x�b3���vx�Ȟ3{�����5��E�nl����Ŀ{�{�����ߏ��O_}�`�����q��f2c����o��{��O�10d�fS>��6��Yy,���zS�_����/����g�q�������_er�h\u�u���1�Ͽy���0��1��C�s����3�c1�����w�u��s�����%eI�f$�������,�J��YR��w�m�Ld�G��>
��IG�R�z��'��ܱ�.��t8gD<>��P����f=�;�K'��J��I���?}�reN0�c%efH��}�γ��z:{ݟ�����{������v�\w9N��:�6�Qo���+�Es���:x+�ܳ7�5ٗ����=�I+ͶX7�gF����;���~��>��0f<�<���'��w|���֑�Uxu�a�1���y��3dq��YX>}��9�ΟzU+�7�߉���$��[�v0��F�d���LeK����s,���YX=��6q�z����>���o>��9������/gj�v"�����jrC��A�����}��w�ڼ�����=�������}����dC�Ȇ3��w�m��c�2����q�A1�����<�[t��H�=i�}����K�c&d�>���6�Ld�;���E�n��r�o�u:��}�Χ^�c02=�>Qe�@�9���u�{�y��c>�{L���pI��ɟ��9��VT������8�3�f!���C5��N�&�۷�7��Ɵ{��o��D�4D[��u[�+:�YR��w��<f$��c%e`��l�l�&e�Ɍ������]�������O̬�?2c0�g��{���,���Y\���6u�z���~��/�r�h\u�u��_�����w����������mf2VT�����3��J���c����gv&>�=&O���o��ߖFV����?q���3,����6�1Ͼ_�kZu��3Z�d�tq��<�Χ^�c3,���&;�����O�yϰ�<���4Ϳ�Lf&C>��reNF�Lc1��~��q��b��J���gY�Q�`Ͼ���~{���6+���C����2y�|���,����7��bѽt����Ȣ}'����>'����Kb����Ca��uܩvj��}.[t��y_��i�^ʸ�����!�.��f�fı�s`�aM�l�����r�]��c��SQ/��)���Շ�z��r�H�X�6H�v���l�Oǖ�Y����dZw�-I��m�M��yk�8�X*�n�r�`r�K	�ڙ��I�{�gT�T�[z,:NˮU��l��њv_A�3]����1ǒ�{�+Tг	pѵ�7C!+yo�0Q.��϶���wQ�=�v���w�r:{=��۶���6���o�f�s[��v��9����A��YzU!�N5{di�>���O���VA]rs����́�[N��k`�&�^�=	�9��/{�f���uoY���S��������w�n��Q�t�
�;��^k�0��ǔг�n���4�M~�n�M^�5�>�Ե��}H\��x.���dG����Y���/�[��o�[�t?�>���@/��]�'X���&�C~��S��s�Ҫ���郱���R�)���~��g,��է[�pި5".;���BV5������.��q*iZ����v��� h�k�]��N܋�c���b����Xຍ�W�Y�1']�MvI�4�#�ľ�r�S�ON=�ܔ��������H�{�ǼM�vZf%�u/�<h�
�|�����m�fe�╗/T&�.��"m`�t�2���9����ɍH��֬�QER
AH�����J���X��ITQTb�[Ad��"�AAFШ�T�Ua*,Pcŕ*�V,+Aj��TR��(�TUT��dU�*1UUZ���"�V0����-J�b"�bZ���E�J�V�ADm�b�Vՠ��j
֊���*-�+mVV�PX�(�QE��E�V,��#�E��UFEU�AdU����
�Q���iaF",Z�XW)h�*c@D1(�mZ�`��e`��[YS
�a)QAb����YUQ2��ۋJI���fU1%��"�cK �cLi���,k(Z�U�*��DQO߳f/�u����[2�b}�W%\��Ƙ�&z���s�@B73d���-��H����Pu�Y\u��n.���q��<��)��zK�ٍ��g\�5�w���/mT[{?��n�|�)b��֋�M�ʘ�ú�m�z��å�Sև8���S��������n ��۴%ͻ͙�Y���si��	�g������؉N�p��㴝uɞ8\/`'���ܩvC�}[]g�]�Z�v�]�zh�jءKl�yx�;�N��g8��֋c;����3{=��[:���$U�{8b�h�{�6�F׌<c��=.�/%�|���O�mP����\m�p���<����X62�r�=�q���v� g�[B���=n�շz�>}���7����md��˩;gu�9ܽ�g$�������8�sѶ:;G���l�'.퍔������w�ں�:y��{H^���Z۪m�n))ύ�4�V]�t�Qx0�m�^��3��9�z:�u����0񣸝n-ɱ�;��yJ�U:7gvm�c��G=t�pm�`)�np�{/�d�׳�6�z�8�I��un��^.�۲��ͱ�ʇ���:�nV�^j=�nA���;�ѐ��28�KJ��sn-��wϟ5\���j=�
�ŭ����=4��(��U��݈�����l���i�ƶ��K��D�m$��7m8��y
QKvy��<�k"�l��s�z��Ƣ��:��ۣ��1�Sn���M��C��Wg�q��x�S��^�+�ܺ�|��7̆!�A�z�]����Ɲ����p����x�6�IPl�v����<[�M�E�w�;cW�>y��z�֯k�ƊŃq��N�}�l'mwQX�=G6�Q��,��ɻi�W][V�3��zAs���$�;��x�͌l����;j�ބK\#c����mO1�{\�n�Xݺqr2#�{r_6��|Σ�.�tr1\7-�x�LMv2�x����2�v�kv݄��tu��荜�����X�VW]����'7Vy�/e�;7&��'dJ��[���۷g�S�2�tr�-ە�E�#��E�\uW�_��/���[��3��m�۠3��v�GYꞙ˳�4&.s�1�r�k�d�v#i�v=�.͜E�c�� �6���B��v+iЖ�*K��E�i<�������["ڧX焠�w��).��In�[p��3٢�cg��JtV�g�j6w&�ְ�g.KՎbkq�8nݞz��8.e֑��|�{Q�h�㪿���a�&3���6��YY9�cϽ���,�&e�Ɍ��ɿ~��2x�2bZf��ﾶ�<d�/�{��l�������}���:�=c12s[��7Z��9��y�N���=�g��eg��g>�����>��,�]��6ʇ��a�c1�K��ì��3+*Lw�����N��_	f2gs��ݧ��~N���7�m�&2c��<{�ۍֵn\m�N�A�~�ݝN�Y1��Lfd�~���;�Y<f8��A&3�>�?�w~[���m�9c10a��`�����q��c%ed����vu��<f0��{s�Kn�E�np����b_��{�����߾~殿i�d���̳<����d�VJ��\�߾����'����8Ɍ�~���6̮��~�IYwd�c����γ�Rc10�~�K�\��Srf'cs��l񓬬�������w�m���{ޞo�<��n��y�x�a��a�\�xu�aؘ�I�q��w��{��O,�J��rY��s��x�Ɏ�Ͽ����n>`>)sY9�Z).�sU���E�y�Z:^ݑ7n����������ߵ6&��OY6�0}����zɌ����������'YY++�I�������)���]���������O����1�gP�b�f2W~}�:��<f0ù�N�t�49uW�Y�Jʗ��{G�}�>��w�,J��5Xb���a�;DLR�[5GU2�L\�*um�j#BP����#\]��t�F�MEȁ���z�tPݎ��.{pƕeO���~����{��c&8�Ɏ���vu����&&2c3)�s��g�c.Lf>�}��-�K�C`+����='�B���1U���ḫ೉ц;��}��'YY��3�c1/��{8�3++Lf0옏�g_Ͼ��Ӛ��>�᠉>��A�1���ݞ2y<�.c&e�����᷂c&8~�-�.��r�o�u:8|2>��av2�D��_W���Q�z��W��?l��O�$�c�&33}�Cl���3c1������m���~��Qx>gރ� q��O�i����ɟ�{���%�Y��8Vu�D�b_�}��3`�1�	�co������}�UH��Β��`��yy�"O�&Eo����O��LLq��S7���6��YY++�C���l�6�I����~xf{������9O�[h26p������+c��n��q��G�m�2�e�r�߿�;}�83Jc���1>��y����`�3+*]���r3��J���c�}��:Ͱ�Lf$��w�W�}��z�_9Ͽl�'��c%��1�/=�{��	�������sZӬsU�ָu�l�=��6Q���Dǽ'���������w��sg}�x�pI��Jʙ3���Cl���Lc1��Ͼ�gY�uf!���H���x�A��m�>�>��>?xv��ѡ˪�:ͲVT����x��YY0�1������8Ɍ����zK���	��!N����;��R.=�.A2`�S����򲆂�@�6��B�����ř2�]�^-Z����`��O5T�6s����'ޒ$���d�g?{��l�Le�d�c�߾�gY�Jʝ����Z��u�-y�d�_}�cI�|���U��>��xY�p�3+*_~���g����	��y�:�0�&3+*Lw�{��G4k˯�Tnvq���]Y�����6��^~��Ζ��k.S+�l�N�=��vu:���d�a�Lw�{���ef�ܾ}�����Y��Lf&g�~�!�T����1�����6u�d��v�b�w�{��	�1����s�����~���'zY���m��.l�3{��j�a����\�`�y�������/�c��v��ⳬ>Lf%���q�1&8�d̳?{�8�2VVJ�1�7��{��O�O�$`��~��r��>�>��/�w�g��&2�VV�~�gǱ&3��D��ʙ�1�!�bta��y��<OI��$�O�vQ���G�D>۳��f2VV&3ay��gt�1�bLq߾���<��d�Y���i�6,�1;�#w����}�3�r:kZu�t�Z��m:8���wgS��&2�Vd�&;��}��N��	1��$��"�Lt�:��US��#||$�H�a��`��߼��q��b3�df;�߽��'YXy��ζ��.�.���6âc1/=�{�����n�z��>q�Ɂ�c�����K8Ɍ��ȘɎ�}�:���8Ɍ���/?}��lߏf;������+��J^��N��YK"`82�NU�Q�-������g����wxyxY�ep�9����~�չI�KT	4��ֆ�C�����������c/�����%eN�o~ޙu�]Z��Y��0�}�ݞ'���f3�b^{��pg�g���]׼���<a���a����ì���bLq��]����:��yf2\�313�~���D�����oF�J���(d˙�����-�f��A�*�v��s��8�hgn[��~���˧5�\�W�l���0{��l�tzɌ̲c+%w�{��O�$�c�1���~��T����;w��~8�������_y�ݝg؆3���C�~��_FB�_J��"Z������{���eI��c&s�~N��������c^o��{gY3%�Ɏ&2c���������LLq��)������,�˅���Ny���o�0��Ͼ��q�&3���_b�LҘ�p�1;c��}��:���c2!�ľ���eC��c�;������]���k;��8�Ș�I���J�Ͻ�gY<��d�,�L��L�߷�m�Ld�>���[�U��'�T�z��d�[�0�����>]���OY�,���&?�}�:��WĘ�d���{�y�m�8�����%Ͼv0�:�̹��7���g�}�>�I�o��eG�}�"�RӚ@GH��a��b_���x�I�33,���XY��zr�p٪�>_|~�z΀D�c��y�βu<d���&3)�w��ed��,��pB��>��q�$�I;�}��	T��P[���LFʎ:w��-C�9�W�7����+n��Y�aj�������{�TΝ�cZ�c��7'���B�LlNbBY�f��<�:�zw�ݹ��n��v��m�l�n�c<5w`�,��^��j��(��6yz�-���A�Ч/��[uڶ��g�6����g�ɢ��=�`�ɰ^��z�����Y��KbԎ��9x�q�u�O9x�=���:� ��޷C�.׻v֭�Z疱���](�w�h�4m�,&nP����tq��x��)k��\��Z:��i���[��Y���ẽ������0�<_?�w�u{:.�9o�Y���;���vx�0��C���/��{9�c%ea���^���:�0�c1';�3x.����8�n>}�߶x��VJ��|,��{���1���5�kZ�L�Ͳq:8����F�ޓ���;�Ք��7�����d�+�I��Jʙ���reNF�Lc1�%��}���:�3��}$T+u�}�>�᳽��j[s4k-�³�:��K��op�*N30�1��{���%�Ɏ&2c��Eϵ�~������N�����8Ɍ̦}߷�m��d�VJ�����}���ؓ���ޫ}��3Jc�C����[���6���Ͼ��w����>��I��b_;��p�b�f0Ș�a�����u�d��:8�I�㯽�ݞ2}���]�<�d���e���y��o1�׿e�ֵ���Y�kg6�`��y��׬���&32Ɏ���vw���1�⌬<��xp�i�='�D_}w�g�Ba����f	~��vu�d��u��C����vx���ÿwY�h}��~��Ŷ��7%g���R{��rk��۶��E��	�\�rr�dϳ?h�!�Hĺ9}K���Tļ��px�d����c�y��vβfK1�����߾�gY:�8ɉ�}����
�����}F��~|�1�I�L{��q��gYǢLf&Ns~ޙu�]4�o ������ݝOA���b�>����L��*��=(��E
s�T���Dі-GQt�AoY��?b�(�e�x��I��_�M�Z۬���]���wW���qa~����IyY���Le ���'�|���8�C��J����}���%eI��bLu��{��O,�J��G�j	5[�Y�#6�����}�2Z<��f��iˍ�6������N��LfY1�e�{����O�	1�}�>�3�A}�ymz����V��}3f&1�������q����c1������N����=�/�Z-�֍[np��%eK��7���=��W�v�I��L2�`��y��,�&2�W1�����<d񕒧�2c*]�����o�ÿe�}��}��Led��.���:�=I������}�jf��\�Y�ц?���N��1��c2!�ĺ���r3��<��~;��s]�3��2^s�8u�a��bLf$�~����vv�d���13_~�᷂c&>~��y�k^k�{�����n�9�y���hٕ6t��;yM��鞽ϴ�W������Ь������������Χc�Lfe��dǟ~�G:Y:�d����0�}����S������K�=�*��|ρ���>Gރ� `3�c1矾�����}���WM�]U��m�A1����{�0p�O�v~��ޚ���i?a�5��a`�a���d�VJ�<�ݝd�+%N�Ɍ�)����g�c.Lf?c�w^{��8�>Lf&���KsI]4�n೉���>���ì�dC��1��_{���c%ea���'�{_?o-Jop�^e��3�y5�����]�G;�:k~2T �P�ߗ:/���Ţ\F0�sA�x��'���7p�˭w�|u�0�1��f$�{�:��ٌ�1�R��w�m�1�9��n��F��8��l�N��;�h�p����<�\N^��g�LfL�cϻ��v��c%er$�b]y����VT�}'���a�v.�辛���q|��23{�4u�bu������ֆ�֍[np����ľ{�{�0f2`e�����G;gY3z�������#���&2�W_��G8��2bc���2��~��VJ��&3C������Rc1=�����̞�e;||�]:ۭ)mv�sۛ���0v���y]\�g�	�S`&������-��S5�:�'�~翴u:ì�dC���.�}����1f3`��a��߶u�a�1��w������J�{�2xv�d�,�L�f&o�w�m�c&8{�/��5u��if�\:ɴ�>ߝ���zɌ�,��	���{����޼�y�wG��Ă�IXP��ۆ�laXV��{�i �~�5��������[����_J�'���� lh$��l:&3��7�����2�a�=�G;gY3!f2c�c&==�?w^��o|}�z|��x�&&A�LeKϽ��VJ��d�c�sߴu�z$�bk����4�U���w�N��~��GS�~w����oT�8��C��1���y��l�q��a�c1�}��l�:�YRu�bLw�h�#�/79����s���:����n;x�[�t^9�*�Úw��H��Ȧɛf�L���}�v\>��j�;���u�i]��}~�313[�{��&2c���{u�j7Eэ�6���q��=�gS����g��Dǽ&����=�>��r�ߣO&=��e&3ߟ��m�8���a��dK�~�gY�tC�c1��Fc�}�GXtN�w�n���?�w�\�����5]�h�����o�e{v^�Ay��2َ�4SƓ3X�}��Z������g�D�b^���x�I�33,�����t�����\Ld����:���q��������~g��g�9��l��&2��D/���g�1��~��7ض�iLu�u��c��}���0�1��c9�＾>e�<f���w���1��&3e�}ì��3dq��w��h�'Nٌ�%�ɗ��O���No^?��������W�}���sW4\�)]k�Y4�q����gS�Y1����W}�t/���d�I��zO����S��ȩ�Y��a�T��3c1�����γ��3���C����a�:�a�����R�Z�ܷX�:Ͱ�c1/��{����N��T������}����z��,�&2�W�Ls{�βu:�&&2}�>�0%���,�%����|!z����d���^{��g+*vk�r��4�U�h�y�N�w�ߴu;u���c1f%�Ϸ�m�t����}�f�++K���ì��3c�Ę8���h�'{f2\�c&d,����{����I�� >��dO���a�
.T�������n���l�����R �&Nw�<b�}� �ނ��	�{&}ܒ!��͛J�~�*w3��8�A��a���5�=aɗ��v�ۭ'>��9,�\���r9��팶ו��mNɧ�X���'s�֪{X���c������i�y��d�]P��;s�h�5Ӗ�v�)�9�����6���v�CxM��z�ַ]��U�n7C����͍���ڷOl��۱k�qg�c6+���9�<k�s��힍cNc���%����f.7'8�-gݒ���Vn���G=��	�5g1�=3m�%��d܍�����7/�8H���Z�Х|=���:��c3,���]���퓬���q&3�Ϲ�m�8����?��'r��3�>���qO���}1���}��N2���өmu�5�6Vq����~�����YY?}�ח˯���ǹ���ߝ���u�0�1����ߴq����:�&32���op�9�Led�����ϷoC�w���q�$�be�������:�:�N�}�h�ta�c%ef!�Ŀs���8�C��a������o�m�����Jʓ��1&�?{t��r�d̳?o��ed��v��oY�\�)\��2h�d��m�"v�s88`�ws�}�}~�&32Ɏ��9�'Y�	1��YR����eN0�c%ef%��>��q����W���8>���>��A���>Fcy�w�Z������i�S�}��r<f$��1��>{��9г�ޙGM���z�}��G��I����N�ɉ�����g����s,�ˁd�c�_���g��bfyo�]~�|������۔�/�sʽ�.���e�t:�C7#��gn�)�5Y�������ۧl�ɿ�+=d���8�:�f�fc1/�����c%ea���/�����;�L����i�I����掲q����^�bg��{��Y+��{���]p�m�N�G=���:�zɌ�1�I���e/����T�)t/c���,������7�Ȗ)��Պ�R��Cy;��(����������w�l�w�º��j�@۞�Otd�>��;T��q��y���e~I��"Lf&{���6ʜ�1����Ŀ{��:�3�I��z��Tn�w�ϰ+]�VW�4���~3�ߏ4�[]kMm��a��b^���x�I��c&f0~��9�gY3�d�VJ��y�+߿p�od񕒲�V~2�����s,�˖Lf8���>��q���o߽Os,�q�Lu�u��|$����w(ߏٛ�'���$�O�c1/w{8�3�f3bc1�K��?p�8ðLf2VT�8�߾��Oy���{|�d����f&}�7�m��ɎO>���9��.f��k�Y4������'��&32Ɍ̲cϿ}���u���L�{�9�P:��3�zO���X���A�c11�3�_���γ��C�c1��3}��:à�f0�x�3�>����>|������{R��(s�q�F�y���ͷ1Z8�ݷ<P-��p�n.�����y�Z�#!�?3L>Lf%��oa��1&8�dɖc��}���u�2�d�"c&<��q���}�"�S�|}�}�w���1�c.BɌ�y��3�`�����zff��[pэ�+:�a����N�:�>��I��ݾߚ"SO������}�df3++/��{ì���Ę3dq�}�����rY����?v��&k�����Y�D�zL���� �-�4e���:��翽����&2�Va�Ly��q���bLf8$�bt���M���;��%�b;U�JȥT�KM���5�݃yf�<�V��~�����^�s|�֞�� og��K���n;ۇ�1�J4phJ�lW�Ӌ=�����&��*׹�;3.Y3-R�(�a�:uW��6%DC�At틥�G�V^;8��yy!L^'ק^x�O�n���=��������֮)���,�_J�����Ǻl��E��x7��� ����XЊ�qY���܈ʪs�ˁA��M�9��[Vۙ�sk7^z*�<�؍N��*a϶�D����=r�^Y�sqt�����|I�������vvڇk����R�Qf.��cj����=򝬘7:�Ŏ��A��˼r��4L��:e8�8ʥa���wT^p��3�����_{�;��l�쨨[�
��D�7��n-Dq�0)���f��o,���b.�s���|�~ɑp��D�i���.�E�u-̋�9~��L'9�̄4F:�ZM����op�5�i�d���٫IU�4:$����HA�%;p?/b��{Ӷ�{���X�3��z�.�����Y%	�l	įMb&�I�1KsBx븼�\�OgC�j����[��[<�� ��轫tw���~���e7K�1e���8;\���d���O'���<Z8� ��.%�P��&=��m��i^<�fO���J)�z,!(w@�r�[�N�n��Q,�Q��5m����e��:�o������J����[q?I�����n�m�g��������\��8rwQf��I>�FEUR[A��Y*���EE���F
��8�(m�FکT`�i�W�S"V�1�3[-�)b��R�VbV��*����2*�Z���r1A`�U2��b���E�����ɕ�Z�)PX���EX�kJ�jT�9J,c�Em��LaQ.dp��QjU�Ć$�k0�2�e�AAQ��XTY*�̥b���*,
�#HcR�-�4b4��r� ���֥k�U�bT2Ղ��,J�kV"�*�(�JZ�Kq�E�������*�UPXb�X�
�Kfb�b"(���ł�-(�J1QX
��hV�����}���S��L�`����q�gD1���b�y��h��Y�3;���.�e.����gXu1����������U>>�=fO���}��}��vu�2�d�1�9����'S����1�/����l��������ﵭ{&�Y++�.���γ���:�ޞ�q-r�������>���:�a�c0C��1��������1{����إ��?a�z��8k~C���D�bL�0q�������YY.I��>��A��q�ޙǙ�:HWQ������vX�l=%�4q�ϳ���}g�>4;v�C����<���{u�[���Ǭ��8���y���%gL�c+%y��s�N�c1�������m�80�bg?~;7g>����c4�	{�wgY�JʇA��Cc��{��:�f0������F��k�Y�Jʗ�w{3`8�d��wy�����s��}���%�d̖c&8�Ɏ��u����e_��ZWe��\;��F���<�g��:��d����N%
����Ĉ��T r^�>��=vy��^]�T�Id�i\�P�&%��H�ζ��*=��^I����Ĉ	�7�� {��3��@st����L�1����'�I0i�7"Xj��������6���6ϹƾCnx�ZO`8v�bjt�o�tx��?���|d��B�6Ё���_��P@%�ڤ��d��ڗ��{�wq ����G�-�u��m5Wo�:�܉�Ew��k=��n�S�Ӹ��ꭎvyv펷/�n��$P��Jev�(S$��SӠ�ܻ���k�_P} o�݃���$�W�+�{=�ݝw"  ǭ�u��JNa�.$vY��븠�#+�����\��y�)��� Ǎ� 7�n���׵�/nve+�[��&�1D˂.R[V�A �����  ����s�ܗ{�ڰ ��[IPo���k��h��2��B�{�l���3�o�����P|���� ��A�3��  �ͥ�����"b\��.�V�@	VwU/D/T�y)L]�p V�]�d�]˂����*jhT�Բh��i8�g�Q�=��+_F��s�����wnV��h�1�:{=�=\ܻ{�j2���N좢�K�֓�i4�P��&��N�&j�\�v�U�1�9��k��v6<V�S�����G]k���Aċe�B\�{tE�Nrޭ]��_m®���n��k�q�ɘ�h�]xn��Q����׋���;s������7��m����]\��'m���V�e%{��V�v����,�Zq�qp���ޱb���۶������wfM��͚����5�-v�A/9�9/6�-[���G]�Zt�U���݂n �5m�7����gn9�(@���W��( �ڿ�>�"����z7qMQ��{}Ifc{�" �N�۰n�JI@��(��Z�Ֆmt�f.�׎VU�� ��v�
���+���P�o��|�zt�I�p6�$vY��븠��Ϋ�Ā�"W���cyx� G�p Ww]�X-��$ELЁrI�U�U�ػ̔2���@.۫�����w` ����d�x�yp5����1�U�Kp�L��]���t�%��Q�|_�N��`}�ͷ@
�z�� �������z��TP�E�9���)�L�mvն����V�˃����e�M��Vݖￇ��}��%��R����;���� >m%]�A[޵Ln^G�Yn� �"
�ۿ�>/'�R7(@���s�'H���y��=?��ձF���LѾ9iQJ|���j��Э��zZ��̈���5�P'�����O�n��u;h,&��ç�S����Ϡ�ut� V�]�`>n�1���9�/=��~~�nl$�(�*%;,�����]P|�;��p��F����  W�۔�|�D�IJa�N"Ge����f�O%�|_��`@-zڠ ����ʫ�UWy @��a�*��ӆ(�pE��-�:�  #�*�����>����6���� -�u��ܲ/#�S����m�v.n8g`�q�S�kf��Ë�,�l��ČS]ن��nS)8hU�==�p� ��}A @��up	£qv����I�vĐ���Ҟ�biA1.P�vE�uҰߪ�Ϲ���Y[H ��j���UX�{^�j ��=U0/��RK�@��+�������Ň� z�ٜ�h崽���"����ȼ����V�����=�>�n�9��O�UƆ=��|EAٔ��J���W��fo%�0J��3�T8�g�h���;V� ��� �}�W ,��I"A9Q)�f�?w��&�|�ހ $ݘ��N�J݁ ���������wx[*��p�I;,��z�"� �;j�^�f���*8]u |fe5@�� ��޻�&�"k�ѾG�հ�	�KcV�I՛��Wac���X��M�y�;�H�����wOD�M8b��l������ #��T� "��͇�B����x�������IPo��.�e7-�P�R0��˸a���ݾ1��{([��J�]y�V��޹J�}��3��ow<�@t��X�PLK�!ݑ}�w`a�W��REڜ�]�%��|��J�ZoU�/&�������_��;���� @EV��Ĉ�+g���������U�dr�N��{DN�JZ��Ʃ�d���RnJ�g���[^�;G������ =�c΋�2��p΃�#fz:'0#'Ovj� B��ߤ�
P�@��m�a�$�����P�{��H'׷V i�r�����oB�=/�J{nK��&FNy�ŸIڗnX�������ۗb)cgt�]���W|�"xp�&�D�΂7�� �ݫbD@eu4���5��������Tl�*��A\g\�U�>����1D˂.R]V�A�v�9�x��鼪^������+�I%^�님�ﶶ��+�S��m�P�I���|n]�es��>	Y�'W��5U����"+���}biA1.P�VZ���sq��qn��|fT��" ���j�� �}����".*����^㲥Y~���Z�����P| r�m\P�q��ewQ7�R�wR��\�H�}����@�yLTt����^�y9�<=%kN��k�{��k��{xek�]휁����ޙ;�ӈ�Ip�i�a9powl8�Kɹ�C7��>�힔�&r�n�	�ݯz��X��a�]�,+U��g���ݵB�,�,s;��%ڶ��4m�h1�s�玷��{n!�CǓv�g��R�t��o綅ݶ���lubz6���h��yR��%�n���u���:i������=fx�ձ6M�Ŝ����m���<�T����j�-gu�+�4�,����l������6�ۍ��s���,r�����7���]%ˁ'.]�����)C�vtG��$���@D��S��:�l�V������{�qD���>�#bX�M��r�z�(�����U=�ou�Ā"����7�n��W�f�62���<�Eu�TA���"E
&\s`��ꄈ���u]�|�5�X��O/a��`���n���N�6��m��B%'�
��NZ�OZĪ�g�ܽ���Z��@|�o�݂J�g�N�����[���n�Q�Ҟ�c!A1.P�vZ�ۿ� ��꿤疜��Ϳg�-�ݪj����v �=w$U�镓0��S��BX��H$-n�@�-���wA-��\�s�u�=�z.�htE�n�~��R� g�{���՞ڸ��+���g�z��՗[�M�7P	",�e�!gdo�3 �F(�P�'��=���رm8��n*�O�����p���I�*/w0X����ؖ
=�i�������8"�R0~kd��f�f�]��<�ݴ���x�S���8������=w" .�}��뚦��>��lM8s
\($v\A��븡 +�v�$/L,���z�漼�Nz!��tI*/��Bb<m���"��q1s���o��8�`�^릯�>���p �͎����._�S�D]e��T�fmJO�p>�˹ Ies����R������ ��۸�	est]	T��Jȱ'c5]b�]v�x{kՎ�6�ً�ݛ��9!��SRd�ǻ�
	�r�:�-{v� 
͞��C� 2���Ȉ��v3�u������x����D%3	)O����A7�m��/Wo�� ��`@\�J�Ӯ��S�vF�30
%�@���^��X ���	���4q��V�+�o��ה���WA��a�zM�r�w+���D;�yܔ��1��n�*�m���n�훃64&�@��D�өǖ� �
��]�"H���� �o�eM%��($v\�^�v��e�\�w$���d��D���+i��4��u隫Ȟ�����u���ڿ�"{��D�bb�.&.o�[~u$��U�{7�g�R�ܹ�7�,��� 2���Ioe����J{���{{ӓ=�ܘC���u���s�kF���ۇIt���7.݄�ئx���o������<q��m��_�9bJ�V���oe��G��.��*K��X�� uctA�}�� �b\�w^�����OMvd?es�^N��@V�T	�{.� �&���3������)�����B�-� %]��k� >�ܫ�, �^��_�}�$��z��@�{.� ����L��r'e�^��4�6.��� ��mP$D.�˫�"
ힵ�SWD1�-f_=L:�8�.��aD��2�-���߇�OD�4�"y����wf�8��s�L�D�ڜ�_,՗� �Stu�t��*ZMGb�����U�;Bٳ��}M���MTG���d�舋�<��'7-��VzG73tv���ٽU�`�����j��N��8�N;e5�m��!L��^f�	L60%K��zm��P	G���$�ݞ�")��K�凯�IP�;.� �t\�$���.��9b��#v$���J��P� B��]X V����">+jX��S�E���ԢܐA1.T����۸��vz�$ �0��^Y�[��w��� �̺� +����d�
~R� �����n�\�2�����Wa �^ݫV ����b�^�R��$t�j��D [�ę�0ET�iB�}��J��Z����g��Ο%Ы3�W DVg;I\ |�D�"�h�+�H��;W5�B�5f�͘q������J%�m�S��=�-G�R��b+�^M��q2���;�<R�7�ԇ��ĉ'u��Q�{��9"�$ܨ��7T�,}پ�l�N4$8�!�+ɖ\�W���~z��2��-�(��q�3�w_nu�4�`�۸��}|7��e��]'q`�q����3t�m#&��D]�����`�^M#>�F�MW�D=�io�k��;e߻�y�s�x�˲�˽��/�+n��V�ƕ�S���Y��w�HЀQ�f���V�V^ƺ�8�U v�M�1C7ED�p���Xaܾ��^�'`}��x9���t�j���|;��%����E�
�[�F$����ڰF~���:=G�Cp/K�Ȓ�GU�7ʼ1&�)8�Od+{�i�D7J�����q��t��yJ�+�T����q�<���~�[C8������`ųI�i�'��؈��]8�@����fi�|����<J3�)��<+W�E< �gW�Z��]pa}���Z2�ȼЉ�I�/3����7x�xҡC���A[i��z��72�xE��PݳjE0Zɣ�)�)���a�j���.�W�>0��+�vC��h�����ӫ���N�z� ��3۸�ba��+�|�!b�u��dJ�Yƕs2c^�ӂ_�bD\��2Zu�X̮�p��[.h�������=�s�r�ҷ�_��k��	�T�������ҡV)�DkW�Ub��,E�U`)Qfe\-����,"����R)�-1F,F"*��ʅE8��2��b"��`�U���ej�12.Qab��ab�,���1F�AVbS.eDV�V5�QƊ*����AH��1Gm+m�ej"+hf1+%�ˁE����[(Ԣ�l���m�k`��J�L�K�W-VT)m�J�FEc���ҫl�+DKimQk`�m(�YH��b8���.Sr�Tˈ1rյZض�b֭�X�˃Y���ʷ�Z�h&e�Zւ��Q`�[Z-ZډTe`��)[.7(��V�EX��j�-�h5������.f�U�q�nd��TJ [lV)V��l˽[��5����֬g@F���+�u��sk��p��;�����u��n���]d�7�vN^2�ɅN��f��ܩ�s��<�vY����ٟq�xb��E ܞ!"^Va�vNR�C���ݧ�յ�&}8�l콘��9n˲��W4��Ӷ�G/\z�e�*����#��}\#T�6�8V�p6Ev��us��m���]����8�V<�� |n�������wm"�J=��e�|�V����z1���Yr3�����ݼx2n{0$w]f1׶	+���yܔX���W����lV��N$8�s�¦��JZ����S�9�7�њ�81��8��uL�o^k���{Q�s��"�<.�{q�&�z�6��*�|�XS�F�9��y&�6�j��c�^r����m����U�R��	�ca��5'h]n��q��n���V�6n��<`�hڅ:�#�u͎Nk��������uÜ�_F����غ�҇f��8xJ۳�]$Y�#�������.-pfQ�ݎn�h�9����x�9s�ô;պ��+�u�$8����[�m'9��Ẑ�6�e�۲�hq��Ƶ�[e@ת����9��O�չ-�9��=o�ⶲ��q��n{#։�z���j�-�fB�-FNv�d2v|����z��˜q��s����}��۞�vM�<�������!�m��]�h�s�p���o'\���O��\����l[�çҬq�;lV#�k�ղm�t㍬[W�c��)�f�mÒ{x�ɭ�ڰݷ.��xy.!Wcl�(���W��u���!�8'��8�6�޴�vm@q�J{��A�au��v�m�����H���n���B�l�{m�mqj���q���g�m�v��tv��%�{S�Y��A���]8C]�.�{�W�lq��M�	m���ŷO�Pf�۠�v;H�bc\�h{\X��Ʃ cm[�Άls���� jⵏh;t��ֈ�O.�������7<��^���qXNWm]�{kc;�s�r�F{n���%s��W���tCŊ��{�v�e����%*�q���L��5�^:���qK��l���]n����v�m�8èTzw6x�k��l|\���|v �rqc@i�@�X�.^�g��g0q�guϷ)�Ի��j_$�P!�1nSۤ�5�z�-Õ�.���q��f:ۄ�����K������[�w��)Hg�nK�E�s/�������g_w�۾��wbG�[��+� �">�� 2�찖jj���Z��舋�ԗ�����bb�.R��[~u��s�^�"�e�z���쫋  ���p	%�ͤ��EK�[d��j��Ȩ*"S�0�=z�> �>u� �d��P��0t�  U���W�|�D�QԢ&T�P���G��7���%������ ��j� oe������.*���>��^w��O�[�U\�k� #�r�,�.��F,��%R��j��K�[����Vs$ll�T��ĩ��.�K����z����㍮{{v�r�X	Ƀ=K��y.HΗ?bEbC7P8F���G� ���	w����T�wT�I�swr  Φ���eKr���($t_�G{�w�퉤�3����6-�N軲
��*Y��+mِ�x���Vv\]�X67���M�[�C9FtF�;��gN�Yy�~�s�{j}9���@ |{j�� ��u`D�3�'�qE�����!V�9�C�S#����y��|�쫰�����u�[��z_�o� �;)��@���-%�L9P��	�)����ʗ~�Fl 
�}B@GveU��i�x�u��Ɵ��:��n�"ڔDʗ*Ҋ�ڥ�i�R�N�t��O��[�گ��̪�H+�۶qj�7��ܘ���d)&G
���n�^�<Λr�k[���4o#�9�������Ά�m� �} �5�PQٹWa |WOm��yz��m�Uݾ���i*���ʫ�#bd��M9Sv\GeʸɜU�gjԫ�yA �7.� �;n�b6�+�.}C���N�Pe��SNT�����#�뻋�
�6��`z����ɥ]sQG%[Șe������ɷX:�cg�eK��d^��74G�+:)��K�su{.��H����7{�Vp�f]���4gTf/e�B����� ��J�+N۶*޲�dL�2܊���yɤ߲��{0���v ӽs`��o\�9((�ŗ��+�+Q�FEJ��!0���vĀ¹�2�r6Na�8�D��k}��$m?��4��Ms����=�*q�t�$^B�#�0�χ��v��3z��i_<v�k�Nt�k�۲�����ѭJ"fG*$x��v�,>�W��=5�*��po���ٝt�W��m�0/�˄��6� �w�si)�C���]���u� ��{nn � =\�+�sn���i|��-쎂I��ӕ0'b�_T�� ֶ� 	�����M��" ���v�| z����4܌MGe���;���d���V� � ��i*�wv��u�s(�%*囧���j����	 :Ww�m�G��8޴Ȥ�D�R���U�D+�K--�Z�:g�Ĩ�~�I�zr�B�ӡ����տPDQ�쫱�N�3f�zI��J� �����I{��.�����s.JB"eB�)�r�S؇ݦw���6�9�S��

�����z�����c�͌����p� �Ψ  ��ʫ�+!��c�u}�ATm���| uciT�D[R���ʉ��_v�+���W�U>�_�a��|[M%_���I �ŝ%�:}�G�����\!�
Zp*��[I%��Ϭ> &$�lwҧ{'� @�ͤ���t��܍�I�#NT���Q��t���Q[ @*|� !_�.�� �襯�+k� ��5 V.Ȑ�)�\($vY~�� ��WΕq��VU;�6ojU@-�˫� ��ݚV���E<�nh_�y�|���yAU8�FT�ȥF�����k����Tbxa|�S`}����wN �8����K�@�2����:t+�cQu��]���}�7Z�^9�vp���ve��m`K�Xp�1;���v��H�����)渶�砄�f�ݶ�f�ܼ��{v��x�ʴu�o�#l7nn�;���o�䓆,�t�����i������Upm�W���7l��[�g���;p�Y�h�E뇵��\ֶyk�瞹:��s�k&7`�Z6`5n-�Ӻ��-�w�,v���+�l��is�S���N����������L�"֖o�1"=��J��������O������" �{�.���wCP�p"����w��/c��&�~` �ݗIX>7�ሀ�'I�?zI�d�9��l�2`L�T�1I	�IA$���$�k��^��^�j�d .�˫� ������0KN %]���5yN����힋�w� k�U�X� z������\�"�����&�xՁ�]\;#�*eH��`N�:_VC 4�u�t08z��^S�۫�> �;n� =\�~�h��Y��[ip�PVڑ�ø�i�e�u��n�:6�u�|�L'1��bAk�)�����o�wv]f�_�> ��u4����v1�Ndc}U�H2��d^�sr�r*w ��ڨ�^�D�92�u�/@F��f���-�����x���$&��C��W�Tw=�FU̦t�@�����.�J��U���֑g#�©+o���� �m$�^����V�^��pl�TYP�%�L���h��@$���@��O^U�N/u�^�	Y�r�W���:Ԣ$��$wq�μT��U3���	k;j�$|c�i*#��[ss��3}k� �;�U�]�|)CD��U�+�:���Y�WF��]�t����ۛ��>n�G�ge��oJ�Ǿ�OT|���ú�bdݚN�on��c��tn)����0�.���)d���\����D̀ےbS��|n]�s�T @ge�	��6k���.����v�@|�D�j�D�S��iA#��9{�w�FA7�F�w�y��\0 <����H���t�[�O�s+��̵���a�PH܊���󯢃�=��J����K��<�g{��A��J���3��G��m��~��4g��E�̞���h�z��#`+М!YG{k3T�C�a�Ǫ�X��u.�̨�q�6�^םJ\>n�-�˫�5:�C�	.&fEw��{��[&�P�� �΢(H�쪰V��(�#u�V��F��S�6���n"I�GvE���� �oOP�ߖS{�#jucI����o�� ]��I%�=wW��1��u}c�<�BZ���AI���"V���
���N����v�+�|�UXn��뿿�Ϣ�k�@�bJ�� #sr��� "��YpEF���*�'������N�i$�{2�(���)��dħB���萀k5lO,��`���޶��$-�˫�
ޞ��$�D���ع5��GSo@��]�$�.;,����, 
잫� �N��L�Q�6�|	GoeU� �=w&�\�3r�F�T� ��n���bQ�nmƢT@����  ���$��y�q1,���B�������X��)��4��Z3u����y,��ā�b�;<����%��{�d��"h���#v���s�����|�Τ�+�R�!g�.�� ���T$L�������+ >u{�*3��s�7k}�I���Ձ�};w >m/G��������Һ6"\�U���栊Omc�o�v{5b6���87h������:������A�۸�$��z�� �ϩ��{s0���_]Ձ D{=b�+إy(�3-8@�]��s�� ����ק�4�q��[ @u�ի ����$��~tG��u�����Y��
I-�ħe�=�v��K^��" ���V�s7aӺ��> ��w  ��� �^Ȓ
qTf�1J�ىj���oMl 畹� )�%q �SU F�eT��{��-]���݁�w��Jc��ȭ�����(��U�eL�J�6
����/ <m%P˷���e���V��ڷ��"{B�^y��t��G]�~�i�����6^�3.�`2�үA;�"PR����i����O٦Fy���"��J�m��Z>N3��n1��q0ٌt�u��σb��N�,��L�l-��]�n�<tŷuOF�亇�;��ݽs���q�xۄvՂ5���K��B����շZƺ�3:4 m���ή�����1���c���m���\�v�g��(��CqlكwA���`$��Ӣ��M[�;��u˘H{!{[\pz���L����Ī��xJ�]�g)��qssvl�����Q�M���(��]C������O�˕32-��s��>9��" ���޺��%��}ۺ�=n��9��]��g�J&S�GW���J�^tX#��d���1�@�$|Nu4� �zs���#�T~����\$�)�ų-Ä
U�����	Gf��,H8u�{;f߯׋�@;��;{�I\.�ԅ"���ħe�����&3�{���\��T��� }޺�Ww:�����&ouT�@VkuQ�@�L�
	o�wv @Wg:IE�Ǐ8^�^~����[MP�}up Ww;�	�#�]U��ӫ~�KPE\V�k�`Zg�n:���ի�����N|��\�ې�&\�c��ـJH"W:.\0/�기� >��J���5Ϧ�������d�9�D��]\�Ր9_)��12J^���J �һ�u�*�k!紌�ܥ����dJ��þ1�=�vv.2˸��������Ӫ!I���\z�:�?woOg�'�y8w;�r��N���" �!{w�W D��up	$�7�3�x�&�RG�)O��ߑud^��+��Հ��.ȳ��)ة�h�!^w�� U�ά��'rۆ��*�/��v�#�U]N�Fh}�T�"�z�%pǛ�z5�Q��R�-gm�����
D�i�q)�]����:�"OW�2⒍��V� W�]�����*�<��Y�z2�*�B�!��a�����'����v�ñza�Z�qϷ[\�b��_��~�s�}�9p�dz(˺�����u`D zk�M���˾�(���Y���`�n�W�]532&�eH��n�/Ρ�j���mx��WE��|{��\�X����I�e�UQn�u;�KUV@�|�\L����{����T "��8M]��}̧�F*m�����&.��<<n����\ߵ�&!�[8d��;٫�zo#�<�o���k�#�w�c��~H�Tw�>{��<�q�*�u��n�M��%�l�%�a�-e)"���!����44��3el��n� �8{�]�;�X��P]�K3.^7�t0�p:�!���.��tuDc� �B{u���7;x��n��m�+����ً�$��^v�h=���_��Ŷ-Y��k�K��"7��b�jE��#�E��is\|�̉�w7�uۋ����Ǯ��ْm&����wXv���������<�Z;��ی>BS125����.�z�+$>>IgN�-^�|@+j�vk�H|����o�Κ:�(��{y�:oU�8��z7�4�՚>�]4�*�n�f�ˀI4�:�2��f�Z9_>���ҭkT>����5ǧ�4��w�}۽�(���pqK4�7�����F_^�n��m-���=�,�t�
�*_��-(��c��C��!4����3O�����o�o��J�o�uԱ���Ui�����t>@^Y}�;��Ag0P�Ǟ/o����:����Zb���;2K�۬�X�Q�m����yF,*�^jz�F��.ձ���)i2&������TyM�c�6���3���6VN���1�|�E���ߓ�|�ݘZ.�����[�f��i�d�"�##n�Mb�`KrYp��RN;�E�p��(�����q@�sjJ0�&��^�����9 �=Ю60U��*1*�US0n5�q���Q�.YG*�J�֪�҆\�-CG2�R�k
��)(�*���a�UR6۔�*�ѭ��R�H�V�-""���k�C&Qj����9r
a���P�Um+E�D�PQf%kU��4˙�m3,�Ҡ#J�L�j+�"��-r�cJR��)Y�.fH�4`T�
)R���5� լ��mҒ��`��V�*)�k����s0\V�J�"�Z�Z(T�JZ�
��(�����H�*)m�EF
-cmAZ,�J,X�@�#�«�T�D*Q���Ɋ�m%+r�2��0�kj�j�-k*�֢�mmKV��)���<��m+w���� '9�ؕ{�@�1Ց{�}�"f���J ��W @ J�v�]d[��OR
�=v�����<��.\9%]���T v^���o+m��V�_]Z��w�A$������%M��P�ݞ�7I-�\-��V�V�kZ�-��q�^�lNy��N�UivB`M�g��ЂD������e{]� �{���n�]\K��}��,��w`� ���=� ��D�Q,vY���� ��<�V�2��^�� "�� ��}up U�c*s�}O4꼚s2&�e)l�݂��i*�"�z�X֞�׳�~�	�6��!uo]_����q
&���%(�Υ0�CG)��I�"�u$�z�j�� w;�Nzߠ��Y��e�[�����8Qvi��b�1f昁�;���w��:�����6.���L�&'�VWB� 2���]�3>�d	p�(�wU-��:��k��9f��J�嵛up	��D��m�7s)�Q���fdפ�<C��\�ady�v����[T>�>��b�i��r�NB	V����$uf�+�H��uZ��X���{��y�T� ���uq B�̈́0�"\%6Y������{�N�^�{�����`|� �}��%`����-W9����E�H'-I-$���9��XD ��\ �-��;N�J�_e�V���w�列̊Z�I���`���S[��\1��� []W�XG� ��V� >|�G��u�su��$�d�ل��8�XN��	�^��@ �Ψo�J6=���V���B��]\�?o;�@���?mw���L�*���RX���V=k����]iٓ��^P�����3	VG�.�js��s����VfkZ��2�)UE���� �ƶ��[��c��&I^9���oL��:��k��t���=rK�q��v���vt�U��XU�� gٲ���s�����k�`6��<v��;Dfv��Ʌ;t��5r��!az��d�\��ޭ��tŮjz��ۄ޶6��f'�n�W8�ع��1�i���(8��nM��lZ�瑅�;��	������f��۩*��ݳڻC��6ی�wnӰ��x��Z���n'���s���=��v[�;��_�\ip�'z�k�> �:� �����:=�v�u��]�۫ ��I\��4�m9%]�
�ͪ��WuU*�{ݕ���!�z�_��mst��y����[�^���R�%8%�SE�^�w  �]P� ��B��wUV� ���� ��Ҡ�&I��14I��P�	]��7�d��ǳ  ۽u`| VSU �޺=,z�JD��w�c�%�2e&ڂ�K��^�+}�qg��.|Z���7��$����@�7�����������F�s�Ӧ�z��Eư�S�4�Ѳ�y��������;�xK������?^$�P��{�w` :����+;���߇��w�(�k1݂>�7@Aє�f��.dݑ�κV:�]�°~��W��̇�_&�m�4�H˝,�ߵ��x�w},�S�`>�����槗�n2��o�s��{f�U��\ �����v��Wi^m��f�ݚ�-�=����9� �i*���� ��ڻ�E�3kޟU- z�J�+w������HR0���,��+�ۥ;}�{��. �m:�����ꫀ>���J�ޫ���=���$�n7� �6Ԓ�&��;�]�bD@>�upŉL���E� {T�D *�ۤ���Vzj�����-�7�p��Q��t9�w@��]{esSm�P��<e�ĸ��s��lh�2�mA����QBIE_u]�����`�o݌"�n=������J�.�*�YE��|����J���;����um�Z�pⵗ�D���up�����$��y�n���X�ꮍ��z0;3(Q�"%�L��/ٷq$|{�\@��di{=8��# �������Sҥ��7�;����\ȱ�V��Y��D%�W!��lp���w�I�0T����r�݂1�j��;*�F9J���&��W �=�wp��y2�0ɕ�J�s��^I$�V� #��W��WmZ� %�xK����}9�
�)�_m���sR�!�����y�| =t�gog����ʿ� ,{�V	=�i+� �|�%�7�վ�s^�������3�l�[�ŉ��wM�Q;���6��mˢC�nT'1����sjIjr���~�V s�ڸ�� �}R�.��CLWqO�U��=��l�:�rH�mAO��%޵��S�$^�uT��" �Ϭ� %�תc�s~���ޤ�QE$�|����J�����D�>uI/,�N�nd�G�{2� {;w���jtmI7�d�ˁ2j�^�\�Qk�^G<�Q����X�j����_G�l�����I7���t� /=;ٓ��q�<3�=;�������[��
��KdU��j��4p���w��aNՊZDA�X��L;�|&#���a��5TH�2��,��� r�ڿ�O�S=>��@U��%`/���#��as]�x*��<��9z�"���6(�Q{b�蜶ێ�cu�����B�]@��Cr7�������m�˔����]�H@��L �4��iTK��9�����g�" =/������iK�e����6I�����n�B/�� 9g���@%�� !�f:�^���萍~FE��)���w�q~u> -o��( �7!U]�V��2 �%�} F��`A�*�9_)p�&R�:�={|��o��p�|� Dx�m���:�z��q՛k#a�e-��qV�\eI7�d�ˁ2j�]�wA���~d}�z1�^5����h2N~�g[��  �����w�y�ʼQ�����z{�v�T������j<&�BeZ���V�Pة:�Jo��
�;ԟoN�B�禵��)zpg\���n$����s\s�Y���C�n�6�;/Au]��nNѲv^�q�]��8�����ۧ1@Xy�<�'�6�΋��Gn��' c�`x�-j�$f|����yz�t�ڂ������s��nI�9�!	�u�����w��zb�nM�/\����#k��f:]��\k�;�[/niM8�_GfS|�� ��ދc�p�m�P�P���gwǎqxO=t�<�N3�r�m��e�^7/���-(ݵ�n������Z�O"���3]C��Y��:���+��c�y�".Z��`��FcTJ��{��!��(W=�˹R�4�r&O[�a� q�e��_OUĈ�n ��B�\�)dz7�S-��.]���]Б�ud�\H c%a�Y�_^��$x�u�� WOU�&�C�K�D��M;/�
��$��J������ �2���	,9���8u�J�#��ZbJR��L�k*�k"@ ��Rի�/+ۭ���Ž�� �t��D��X>r�����G���\qRti�X*1��&��s�8�=p*�l�Mm��D��?����s�ՔnK?:^ݻ���z��  0|�%>ޛ�ol�������>D\��'AZ�4)�V{���/ד�|����S�w;$B�`���[�.�Ei��N,�=���O�,�[�Լ�&�L��Z�\��w����ƥ�ܶZ� _N� /�� 3k���֯6'����,�]�#�6�-_�ޜ���� =u@^U�}=�j'־�e��\H� 1�u l_��Z���V����9՟�Z(i��b���S�+� 1�5@|��ٛ�u�n�~�ݨ �*��}ײU0�L�Q6�u�� %k}�t#��-��&/|Ҽ�s�l_7Q �"8�u�ͼ�n�q��ʅ L� ���쳺�:�Eg���ͳ��M��m�����������3P�����g��|	,z�(  #��[����j�l��S*���w��#�x�KbvT�͓*\Jd׾-nu��7>팧��<fW���I*�}���l��]Ӳ�n��#���lCB�V��sȠ�" 9g����uyn���Y.�E[V��qSn5)�放hC��WsȎ����f���������Y�Oݵќ�w�g�)K�XU�\��9ST�{��	y�u ��7�n����-9�p܁Ik;Յt�A�y� ���QA�$}��[� ���\��+x<���P s��0�������4�Y��O��q�V��t��I�!�J�zcg۠����#�[� ��;�VF���*���v^�U[�����&�a3-LO��ӎ�5�qz�[��t%��w"��V9ܲu�����w�ı���
�΢���w�� �;�n -���k��"^7@�,��� ��?�!ÉS2�����]��s���2�+�v,�mz �7��� 
� 3-'*f*k�3~�� ��7�d̎%1��k�n� 
ޞ����۲�DզM??{}�����@�ٖ� ���=��4Kbʻ����g'�~.�;��ͫ������%`@y�n!]fW<���ɮ��۔�&�ÇV�RǑ3�IsQM��&W��_j�������W1�D�Z[<7�Ǚ;�x�j����{mt'�`B���-9��nB����N]Ą ^���=O��n�ᰕ��;� �'�I+�����2�}M�t�I�[310�R4|�W=��(8N���k�dk��<(V ������ԑʗ��]�u	%[��$� �2��D��Uml�qm*Q"-�k�`ֻ$�
a�K%��w ���(���I^ɞ��^�k`��_>��  ���U ����(�����J�5��ʉ�Wpe�z�D�X��	6Ⱥ7�>�5�)� ��v�$I|�C6&�l��Ħ;�-om�����#�M\�Κ�"s'�� ���U �v[�³��]L�����wH���Ƈ0�L���W�uA�,ܫ�&"�o]J�����������`�m?^��l��$�	'��$ I?� �$����$�$�	'��$ I?�B���IO�H@��	!I��IO��$ I?�B��$�	%�$ I9 �$����$�@IO�H@��$�	'�H@�P$�	'`IO�����)��$��3�o�9,����������0�߇��B�  �P 
P)�@ �R�UA@J(
P @I P(�q� #:   (
	
�� �HP$IAI
� AT�*�A@ � ��>�J%@��R"� J)*�) *$�*�QDR% (UP� (/� `U*�J�(�|A�	��+u��F�8 ��Q��F��1
K�(]Ш���R;�U  Q@��  �}΢��ܔ�� �UV��	��
�v�U*���Έ�R7g
%fj@��B�w`�J P�{� �P ((
P
�>��wJL��S�uB��,�T�Y�օ媊S�wB���$`aH��Tyb�AG| �>6�*[�J�q�D��9aTM�ʞ��ܥ� �=�@��+���j;�9UK-UOm�2��P � ��(((*J$�(����(b>ڽ�uJ����UQc��tR�Ȥ���=e�wUS۽oUE\q�(�ۈ��T�'� �Ǔ���qR8rUgI�t���P�nV�tR^�zT�T-�Ԁ�U=���on�T(��  w�*J)���H%I�����r���UR;��QnT��B�j}��1�����/[��*�qTU��N��֫wp� @���(����^ ����� '��
�  4{ �á�� {� q��K������ ����8���^a�� p��>   �說Sl	 *��>��y�s� ��&��>\�"w���@�R*s1QN��T]4��rP;�6�Sw:@ P$W�  �{�qBݝN���sA\�*-�uIwq�P�@�tUww��n����Cu�
}�     S�)J��SA��hF� �4Њ~LBR��B`L� �C`D�2��	J       ��&"� �     �)*SM�  b4  !
�d�b2d�mD�I�d�ѧ��G���O��>����H��Zu�}�K3UoW8�@�� V�e��.�G��?�����	���?�q���!�׃�?�?�?���vA��:0��|��8����э�l�;�L
�60l,G���N�}�4����w���� [�й���(+���V~��}��?�`����1j(D17�w�G��8]ݷy���ul�^�0hdQL���V�fFUM�)qI�^V�BD�f"�2ڱ��F#`�R�ʁ��\YX�~u�H3O�D��x�ȝ^V�;��6���f��^��+��u����#�R=�]nV��f�fr���N�-�#V�zȣ�7ncҭdb����l�i�a�T���L�[&�L�0����<�z��rD�N������;�f�{����;�M�ڦ�9�7NL���H�Y��H�35=f�Hݷ���� [�T��[����1��n�	.�c,5�lџ;D���\�B�LLZ/!d�n2�^:�ѱ�iqX�rllC.jm�Cx�V�y.��[pJp�{b��7�ǥ9�l���OqVV��[OQ�E�gmہ6&�%��#KX�k���#���8�.� r�YH��!{>9�70Z.�fV*vDyx7	.��)�5D&,*�R�ZQ��uu��r٨Yw�ںC�vo5.6˩�ҾKaU�l���kg,�Y�p<
J[+*�f�X�^fPG%�Z;��v��C��M륲sR�w��0��G��e+N�i���{�R����j��yy��fT׊���ZC\����wp�AS�6b�b��di��kc1��/�ss K�nPՔ/3	K,�qѡ�3y��8�j���3`��!��v���ږkBwYuvW�`H�ԡZ��>9��^�da��n���@��x�0m=n�Vn��Җ�hוg[a;�6�.&HTT�j�Ys2�:��,TY�hVAʅV���Y��u�N�4P��I�^���ƧX]��ދMY�8-����V6��!ԩ8�32��zh��4�C��+Ef������d����T�W��׶SӳR���Q6q��9{[��ցY{6��ܲ��ۣ��F0Y(�{�lkGb�mp�wty��k�U��58�� L�7Q����Z�Y�Z��Ú�7K7%���.�׫IMV��2T�Ш�w�7M����ܶ-4� �Yi���sV�8��K%�8Ug�f����ܤ1�
�%]���k.�];K�m�ȶaJZo�r�l�٫T�UA�e���4�el�!=Cff� [��9���ɒc����� �3����t3-;�r���l�[f�k�X��l����6������' 39n�^�۹e6w6V�-��Q6+2�i�Y�z�ɡe�in��{#hU�V��۱��<��6m�j�W�z���!�ذf�/J��lO)	���Ÿ��������3bB�@�1��)�w*�lL�)�V�xU(EY.f먤�t�ѤZ�Ē�r��p53M�C�P曔���8����ssa��oK{A@o�ٌ�Z�6~�"h줤��X��ߋyzs�o���Fd�N`Vy嶥�q�DR��7���m��9����V-���GB�F�R�1Kaؖ�c28Mly�$1d�)�`1!��Y�N��-�((7s6�S6u���N�h� �:N����ES�-9j� ֧���[z�n,��K6E`^�/q�;�ob˰[0sK�ӽ)��0�!6�^Q4�]#�)�v!�D�dHuE�#q�)�J*F`{%�f��kf�u�6���^ɩ�b D�Q2�q�ż�������K6ԗt2�� �j������zk�R�^F� MI��z�X)_���ga�+^�n�w^Ib�{�Ϋ�����Ӹ�&X-�,��U�fd�L��w�4�YYjՑ�(��l�*n]�_L:1����0L8�X���,Wݒe,1�8Sj�cMѺ�˨2�+U����ǎպX�
�@t�Fٻ���r]��̑i�ni�!��vsM�Yq��li�E2�nނ���hO)F�2Q��TҜ��;P��wSҊєN�v���U�Y�l���o@��o䤓w�PJ�6]����k�޴"�Yb�PL˶0�t�W�/a⩎�wm�#q2~ͱPe�`��fݥ�����@��6�(�]�`6dӫt�Y�aT�f�d`׉dڗ�t\W�u�d�7]97#ѩ�0E6f����A�!�1����V��ve���	6��w�em�nc�Y�ꗗ�]�snmYjI�mA��6N�꼊ͩ�,��rX7T�:��&-[����DyR�����X
�-K��Q���L!�m�qk�����wv�ݣ5JX�w �Éj�W`��˳-G�mc��gt�����r�X��Xa�ٍ��zR��r�����-�(�*⻻�U,HՓz��2ι1#yCnґf�&��V
q��Քb���2�S �0�Ь���ٱ�n�P��[�pK/&��RA����B_�k�r��w��)��\�}�Y{�*���k�C0R��N�>�b��t�v0�]ӧJZ:st�2�c�d�q%1}��Y" v�9�R�IRM�H�JY3-7xo!ö��"��^+��˲����M�-���mۺSmjװI@15Kh7D�;a-�-�r֠F�*Q7w%��X,�͟9Z�5$R�N�A�ܿ�ZT(Mr�X�f|��W�U��4]�,��HdAG�jlM�0%��A�V��4,�)0u�b��)6��Z4ᅧ�@n a	I@���MIu0��r.d�-t�`j�/.V:/J�[Gul��Jd{͗p� �ڱ�AvTu�5EY�y���u�3bL	h6X�t��J��q6�9)^�5�3"k�C84����ȫzm[�������76��J�;Cjj-J���2�3).Lz�M�m��wp�+7/0ٹ���R��j��1ҳi[��V=-��f`��봝��m�ĵ����o���:�1�Ƀ�Mb�Y�KT�M{q��mV'�h��cTh9fC�[-D�J�M��ڋ�e�ϘV�C>�P�Ne�!v� #�R�U�ݱϰU�]�J����q�VHn.�1)�����v˜�-hx�䊦䥇tgٻb9
���+)�ާ��hM�Gw+-U�c�ѓ1Yx�&3�rۗA��.k/p�n�//r˽����l��*��cA۴����Z(+x�t��c%3����D��nhߠXi�fB,7f�؉.�^^�ą)�������&1�(��7뛹uz�[�3"�u���Y2�3�^�x�`�S]����/��˵�漹�Q���>�ds@5t�J��/L `�G�+��Smm���wykk��5RiU�����*"�(.3Yvb��SۃV56�Mv�7�^�ܻ`�u�;j�a!b��O e�g�ő�H
6^�m��Pެ�V7b��C&�Ț��ŐA`��d�b$3,�2dq�V���J

�9��{���6�VT��S�p�t���8]K�x�l�O]��v.�&�账��n�c�La�2G��".a`���E%G8n�B���F<���������V���+[ 8s&�00 4�^u�֯v��\Ya�B:��
"�������.�2��#b��E���4���H�F٫��b��i�7�0S�F<��dyk&ẓR%�D�v�Rw�t�ov�m�Q�*���,wv�P�&�y����h�]��L/L���� i����Rr1Y��*
.85�� r�@8�s,mf�^�LS{�Fݲ�^YwD�X4�YF�h�t��y�E�֝����q��g�.�nH���L�AjOR�$A�+p]��6f ��,S���T�,a4�1 �/��'c�݊���:�b��d�7^YحK{n�K�͕�eAX�yYB�N��l�sG
�*L*"�~ʁ7��9�k2�5S���3��.M���ݣWF�El�2�9Y�ZvŐ�ji��.�8w2[w6�ۧx��Y���P.��O���#eQ��S�O�8eg�qݓ������^���,�-��D��=�v�C��XT��6�%��N��ܷV��
w�t��<ѕd��<��eŧ`{k�uq ��.��7M�˶Yq 2�\Kf걛��n�n�-�m�I�6ņ'���J�K��S�E5���ī�R�x4i��[ϒ�0�ڍ;�s�Y��7%��]�mȈ,�"�9�a�ZouO�%[W2�+�N�v\�l���J�Mn��Gf&��?c���2�
c T����1"�(@��;�і��m=��VlKȋ���C�V��ҼD��5b�=�*n�?=��1$�7�n���`SH�J�`B���r���T��ϲŚ�w�V:�2�LŲ�4��\�ݧP��̚�$	�H��"�d�.��c5b��V3v���gLe�!�v��oU�1�M�4D��@�	���yC��/d�ǻs@�ڶ�};*%W��h
!��uh�ˡ*��t�8�uu��C�ƚ�2^��i�ܶh쐛/)`a�44�ҽ�
[I�Z�L;l`�ùM̈�,��Aј�/dy��&#Y$�T�nּ���h^�wE�.�H�ie�*z�6Gq�72;��f�:;�i�nҬ���RŻZ�,�d�i��ڧ�Sw$�8`4���k�œ*����D�!D��v�J��O`Q��A����\�w��X�%^8�}S*"�0�Q�4mc��U�C�'�i��iyP���V�B7� u�#0�J��qbjd45n�lPV��u
����(��V�r^����-���4�Y���"1;�љ�V>�b�#l=2�\�B��� ՘�8����a�j�(]�y�vR)<�L�!qm`�,^oU��m�K4�\r��0N�+$��7��c9�bR1v]�ب�(��Hq�u������WCDe�b��Sy��"'�ǄT#�ُ�لf���qT��I0�f���Yn���Q�PԐ�&�F�<[BJ9�kQ�5��lM̽2V�3)M�ǀ�vt���[�݉@�-�5��b܉KT'"I����7�/$:Й�P�.�f��9���T�lcDf2&4�v�� ��L��f��Z�/a*�����3)���7v�e/�޲�EMI��s^��ܤ0�ѣ�� 5�JN�7b �7k먂̲*��L�Z
#����Y��̬�̥�������.�k
frƵ&i��w7D�7����u*)�C{m����zf]�O,�Xb"�2��l分L`A�XN�Q�H�<�/U�Yf��
KU��"2��Ɏ	�Kby5)&�e���nT�r�̒غf���(�A꽨�S�ʐǬ�L���9��w��i�����f��Y��ҖV;�)��e]d�n�"��E����m�yZ���h��/ ��;�`w��r�.��l��S\�>ʆ�in��\�W�3k�î��o2i��oԅ��V��y�X�CVn
 �:CqC��Z���64)�3q,2�=R��7vɈ� ���H!Qy>7�Ԕ��ӕ�~<߭XS~�u�Y
9m�ӱ����(ɉ��1bi�Blֶv\bbܧCpJ�ܷ�Zvn|���@�jTeD�ּ轁�u���Va�5�Rz��z/>�2�����E4��E��ȯ*�j���v�fd�l[�k3uc���A'+/;�dH�����z��u�ͭEj6���2��a�m��(�a��\\a~- ��9S CE�I�}�Ţ�rX�n��VǴ������Wb}i�s%�A�H!VԼ��Y�����7��ñ	�^���h"�3�Tbd(�c$FM�e��d�U����$�h �dM�0m��e���0n�q
0�"�d�ͥ���Sc�{K96
��W[*+i;c2����b��n��l�2.�-�!��w>T�LԷ\�r�Df�W�O�ɛ�1�h��N�1�gus�g���o8~���?&~��A����,CT��>?UW����H��ꯑp��>g�H����@�BCbHl�M��q�l�0�.�0C�6�\1�i��8�\`]�����c�M��`6��@6	2�
`6؜ I���N0 ��l�P	 �l�C'�N0I�m;`�i��l�Cl�av�v�\m���\����e��60��˃l
api�;cm;a@	�)�.6؜��l.�Apl� e��0.�˱�3�Cl)�P�. 2��Lc��N��c�@*I�#@��?���Ͽ�|z������,?�$�O��W0�$$�}Y�$�}�=ψ���"�	���ᬿ��]_�C���v�����E����Nt�b�7"Y�I���d��p�*�����B�u����*+i�S>u{�0u�o�0�!�v3��=wm�� �r�h�pEґ�^j	ϰC[��[8��nl�?[���(__+�)F�ZJeE�Xxo�6�d�g�t����h�\59����B���2��r.�5;�NZbÝz4)��p].s�`��L!Y�n>�0')�5�[����FB*w���ۮ������YŒ��6/p�yY�9���1���4�o]<˜:��a�x�g2��?^�ڡ��|o��1-{.���i�u+7N���y,=������a�v�W�w���*8z���:�ᗈl��0�e	�.ٱ�[\�J�8�����Lՙ�bٹ-��ai<�yd�)3�5fv/^��l���\wN�]�����,
uo
n�S.�0�U���}N��tT�S��e+Cp��6��'ʺ;��^<��K��M��f0r�39f���Z��Q|�KU�5o];�*��X6d��?u��S�v)�=�(H�D���f��魙	F���vYŅW)f�tt"]=9Q�63P�
�H��Q]��乴��\��9�Ś[�9X�;e]�X4�eؾ�.�Q�i�te]L��N˾U���u�Y�L�p�>����P����wn�p`Qņ]�3-v�3��Q��,�7��ym��*f-Q�VDǭ����W�]Y��%@�����n�
1ӏTI5��J�Mح�b�������~B*[��s�]��af�g^X�&��Sor���l'(lg!�:�Z`m����ۭ�}.Z�J�ҹ�(��24��n�m���u��]�K�1�7UbֵeΈ����sZ i���p;��Gb�]�fT��X�9T�Yk�"��6�|��CG:�΅�b�7�MN��*n
�"�Z������J���h�/V��E�r���י���V��z��2�M�&�	�3�Χ�R��؎�ާ���,��r뵄0�q�}؞���g5+�j�hf�C�Lő�إ�+���(�� 4�p\�%�Z��gZ��Z7�g33��Ul��SU^�#����j쎳]#�
�Yn�1�[�Vc�q��'eD��;4�V��X��-�����.����ɧ[4k-m&��v�S:���s��	��Eͱ��҄�1DgP�,�x���R�,�k��)��gfݨ���=��;x�RN�h:w�c�;��Ȭ�@�鼻-���ŏCv���WM�\�d�*��n�n�LF:��R
��&sw"�->�b�Z�Q�+���2�b_���*��������h�:�}�{�+�p��)�O*���/��V�DK�v:y�k7��F
c[�/��f���.�Z̜rHdϡX��EX[�!�:%�~�;;�p�wm��k���3&B]�)�(�I��ʶ����w��ï�,�dm��O$n$'M�M)ܧ�\�h��5��6��탮_iޙyx��'1B���nr���r2i흽�%�w9���8�s7�LH;�ڀ�z���	�P�,X2!���#/	`�o��ݥ�l쓁�J�����^)�tY�Ec�����]!*oe]��\y�W�C���2�r�R��Tx�:��8�ӹXr�Ֆ^,����v	���~�ٳz�ft�p"r=۱J�.�O�d\ɤ��W5)2��F����Z����ܴά��
�Y�J&I�ͣ��T���i�*��]�G1�i���ɡ�Vsdj��ɸEZ�ʀ]�8"*��AgVa�e����1Wz^S�Y��Tj�ޣP�<j$qah����U�_ҩ��;.�*�wӔ���=.�ܳ�5�:�X�W�o31��CiSk')�fg�y�;�l�>�<�emp�'V�V3��V3�	�[��Gɉ�(����St�����³s.��f��,�T�om�k�D�;j���К�Y� gl ��`\Zy���r�v��×Y��^�-�%闙P]3����B�Q�;;.���EO�]��j�ﴺH g,��3,E9\���p��_	�V��{ʥ�i�}�w(e#AϮҼw�pSE[���K*};*�Ȭ΀wd9����pBd2]������wZ�Y[�z���9*5���v��l�e��BF޻�e���=X5���Ȍ�i�͛j�yj�rFH���m�-t��]L����n����T�c�M�>�+qQS^K=@�Y0P�G73w�_sw*sH��8^n���q�%�l�A=iZ�d;|嫫�WW|.G"�j�;��t�8b��Y�wE�O3lc�\����*a�6���IyȌ�sL��6Zw���d&���8��q݊=V2��u�g6�<���a�%�`ASTѐH��3��@��nvY<��2 j��Z��͐l��V�%��&؎�:S�YY�ы��(��0&ZF&��rl�1V�H���[ج�1��l�LL��p쌚��ܓ�ԍ;��=�&��`�[�i�ăGU����,�>�wzu�3�d�]j�󙹇x�sg���s ��w]���t!]_`4���sr�7���ػL>T�;���C�O;��
b1�6���am��ݷBP��=��ɗ���Enh+�s��b�XcA��x�Ϧ���6�v�ڎ��b8�`h:v�[��\�3C� ���]un�gN��3l�F`8��2�J��|��kؓt��K��5dԴO�`�닫͇u��5�H/d5��C�r�fM[a�Jf)@8���f���sm���ZU��� :�	-���Ɲ.$U������e���:����T�2Ƀw��&���,�\˜���  �$�yf��o�{p$,"x_T�t {�eN�0�5w�u9���eU��WӺq,�k-���ԾCKoS���_*׻M��.��Up��3���3�Q�PjP�����\�V��2N�Ř��G#�J˗y�)�i�	8 �s(����Q[^a'E�CqV���^��7)�cvڍ;q���H�N9�d��L|���q�i�wD�!�-���D�`o��	�W�06���5�+Y�z�۽�:]��y,��u�� ˫s6�y6���Y��#
���ާJ�{t�5n�{nl$M�����x���s��;寥�C����3^'gn��2�x0��$ڨ:�r֠�����W��p�+�4���n�TC�7M� �1b�U�+�r�وo]�+.2�)�jV"�;Mj�+k6�.�_YqU��q�&���E'f�������B8hR�+E��vttZ��22��)�엌4�{�p.�ܭ�\5�}��ݣ�EoE�jL�C�D�!|n��a�Yb��B��������+3�mȱtv.����- �x�vT�ͳ����2i�fݙh�������r�kX�v�P52����lS$h wn�-��b>�U���Q.P�����uy�6��Qw�,�g��P�D����-`��c��.�z�a��2��Hq�
���
��-I%� �D�%�M�ZG�"Czq��z/o��!R�����q��k)_E��G��H�R:��'�R�O��ŉ��F�o@����n2�y��֝�T�k���6�ŵSI�"��ט+$�AˁT�!�֧`�b�e��$���d��x��'WXn��t-�B.���4kuv=YL���fYP;��|&밗`�U�9��T�wTW�2
rl�wܳb����,�P��[��moP��B���ף6������p�O�� G�l"���z �U�z�V�n��i&�q�X,����Q4[⾲>��#h�c(��dej9�����sr�Xxs2������L�V\�Eֺ�X�
6,b�S}r���ޡW�������B��Z��10L�����6v������⇷�WN�J�W:����v��wf�^D�b��E�0��No3��$Y..�
y�ub�Z,qh�\��᮲oz˝YLp'�J�a�e��KWfZgVUCF��HY>rQ8�r��l�͜�T�������U`ƥ�혡�gt<_ݱحނy��u6�6��f\�;VV5B�]l6�[�
��x�U,�(��ŵ׼�Ó]
�/\T�Aj�T��z�ڹ��jY�)GK*�mŐ��׬�ki�Y�Yw�02�m��nV%|U�
+F�@1��F��f��_|�!�vd�3D��r'mZ*:̣�� >1���U�Z��oq���P���&6�v�����!��S}J��n��+��dU�v�L�����r�����ѣȥh<��/5�7��:�Ĩ���]G���ku����Y�sQ\ˈ��]��b��\�5��ͭ�b6V�*� �D5x��C��u��R�Jw<5��[۴Ù�w1�"�zp��8Aw{�"+ux^�ʺ�����f��NGR�vK�1	�4��:EaU�sr��C���{���s�*|�:𮌩�����"�+����0B�I�gfS���i����7�QγS��]����n=m^b�<"/F��[�y/�.�,�˰e��	tz���ά_p���B�M�tE���i�oFw}k:�n������&VG���fڕ���ԥ7U;.��>9V��Al��Rۈ�!��3otoʕu��v_R"ġ���j]�jCܻ3n5��>9�^藒W���O#n����'Zss/�n��|Ku9�(�j�[��s.�yUq�wb�aT��BeP�5F�T<��Sn���q�2�ep�uh��0Aצ�u�Q����y�����w��:郏~ܧ��H2m����ɛ��\]š��d�7;ie�<�&γ�:É�2��*�5��Sͼ��%[�r�,�&c�Ҵ���؅�M�7*��u�Z髉|c�v�+�[-el��.�ަ�S9KY��3n��m\)� m�Vq杫v��S ��i������Vz7rY�EM����)V����	�9\WY:��D�Z�ur�Խ9���nH�R`kmW"��=�:Xu����%s������b��Vw=�w�}*�yS�ɘ$��֞Kl�(
�mK��a�l�5a6�<�4c�er9��#&�Ŏ��ec�EV��&m�
/�OW��O:�J�u��/D�m5O��2��N]��oVK���.]e�N������_A�(И�"��U����;�&��H�΅$p���%��;2n���-�����n��;t�8͂��(m7��S�K�(�괪2B|z�-*�)��+P�9�4l�8^ Vf��Ԩ'U���P�x�Y��d�]�fۼ�!�b��
���8��V�!���-���XsY�p�4,�q��"K�]N�T���d[�E>�`�哣7�x.@��TÂ��dݘ{]d�7]V�lU��nVX���b�X�j�O�KT4;K�L(����,����=��Ҋ�`X�0.U�l
�]gx3��LǊ��T�:�ȵ����5ú�ܽ;�]�O�ͫ�1���Z[z��h#�^]B����e�#q������4O;7q�a�	NC��Y�.�dT�n�꾣�n��F˄8���e�ǯuNכ��ˣ�72!��FXZ�,�J2�xqі��&	�כf霧���rA]�!M���!��O)��ҷaVQX3*拍Ko+�ɕ�W�vHY%���=ȷ��b�+t��μ�٘h�
ɠ�ضi瓷{�#WEʋҮ�o����>�{*Hۓ,�|s6�@F���J
����o8 �ܷm̭�+��*��uu,ھz�r�k�f��b��-ި�j:6��ܰ7/v'Z���=�m۳�\��+.�����ĴP�F�iar�0�=���M�՟��" L�&�� %���A���������j�/D�]�emQ��=#q�c]kCvkf�B�6�;5sF듻�3��j�M�T�խG�Tmg�ƕ�I�tF�rv�9Gh]ڼ[�/m���v}���G���V������Ҹұ��$��# ��F4�4f�M�k��9vݼ�,X^-�����92S�fHDs���Adܖ�y��ܛ�d/f���y���cv��	�s����c[���c���ci&�u<�:L�a����5ۮ����q��XҤr]g�Pj|k-����d��k��n�}+�Z˼[ێ�z�k�m�u��]�¶f�9՛���A��'fv�x��I��Z�m�f�'$�۵Y��D�N:VFbxC�6�u�v�tWV�\k���v̋���N;3�Ϟ�1����D͆(�ܖ��`�n.*��Hqq����8��Ĭ`�7k%R]Z�4&�T��,�is'[��ݻ�%�H���m����G]>���>�F;K��d��q�B]c%����\�,�U[!�
�ժ����7<<񽋇'�\t�u֩�\�Tf�uj@�ҍ�f�-�t!��W@�0�\R͜�\� �Ɯrn�n��kѕfl��`�/�����:�O/1���8�����͍� �h���N�bO$�q�w=rXN���g�,)p�0]<��.��wV�:Ξ����pqu����dS�b�ջ��l�X5ũ�,X3&J&���ܹ�3jF�L�D��k�����Z68���g�c�I9y���F����j0^����V!\� �+e6�%ƻ�0g�uOki����7�qI��f}e�6�X��`["J�,�%��%�mI��ح�=�gn��Q�2��;q���u���,��'��:���ǣ[��ȍ���pv�ݑ!�.�F��T�vKQѕ;7bx�yn�i���ñUkhL5�kv��Z�vݵ�ٛ�,�]57tp�وL\��:8���l��1�ye��!0,����*�H8+�n<&"��n����oQݷhZ�x�L�[�nq�F�*�p]�,;��wg1��*�3�fe�Pt&s���3nM��$�Z�������=R\�8�7�7a3m9�n���J@�[wV���>�XMK�Y
��.�(7�.�Iu#���6Ѷ9#��[��79,���ҕs��kc�9��n,k���:��y`�[p�G���7[1�=�M�Ơ�ٍ��n0E�*�N��:�^XU�;��;��x���l�w�q�.���jT��]���s�i�ȝn8�\���Z-��6�2��	����_v )F���^n��v���ݒ�Z+��lÁDx���I;z�ȥ]ol�u�=�������NIzp��=ͯ��q����ۻ2;�6L<t'HY�do*����X�l#IaU���v#j�&{����nd����!m���{�:�u4[����0��V�kJ 9�t��6��r��`w]r,��<qi2��m;v�NA��l"��onp)�����4�o1�$3balq:,�s��-���(u��=G���k�dqL�X�5Ê�`K��J\�5kB�J�0��J۬Z�VK���Op.��}�v�Z[�Y��1e1�B8��m��s���:�9�����͠�sL��ȡ4B�6���{�2aՉθ4�8��Nl"�A�g�Gv-/l�kFZ-�8�\�(*��/k;D��f.�������Ɏ��ўt�B�9�F���]4.%�`$1F݆[p7����4И���rt
t<۵�Q�p��M�s�袓C;sc	��M��܉�l8Hn.�5�j�-$b�l,x���J�͹��n��kƸ3���$<K�s��9x{l[����.҃*-���BKfc5D5a��5u*LL$�5	X8�M���]ˇ̓��ou�s�3�9������b�Ҷ�ݳm]-��A6�9�5�2<��u[����ȇ=r��@�(zS�O�g��&كW�k��9\u�����:
`����.��A��j.#n��;��z�\��/&�����Xkpfкu�l��젽�V8:Z%��J�]x���L���3CQ`��4�MiQc˙E��I�a�+�I���b����eLۉ޷v�7]���iγ-��s솗S���e��\��P�C��P��j�k��sX2� ��s2+{s��O<�g��+6v�z��痕��v��Iv|���ƭu��2��:�0]D��@���-px�73ژH�C����7[�j䣲�ϰj�kۏ]��u�,@���d㔗��0ɴvs[I��d�e�� �֝]Nm�]6�|\�L9am�hj:^L�t�a��n���۹�n��j1ŷ%���<�ƹ��p��(���<\
g��Vv;!��Cd*�R�"�.sm�] ���Ԧ9j�UCt��<W��x����J�-�x�Fuq���0�jkm���l�]��X0b�=l11�;u��u���ݭp�T�i�
�;�Ō�vz�ۮ�Kc�{&��-s&Cfr5���q<�8mat� ,ƚ�R
r�Eۓ�
�n���N,v�\ms�\���.#0!t�cXb.!�bس0�[��̓ۉ6na�2����]1�i�]�ut{99�u!��&�����%u^XͬB[���]��Ƥv�h�+�J� ̥5"�ܺ��V���[om&�  gS۵�gr��c4I%�ˎ=y��{L�+��k�lc�N;;��9u�&`�J�+�z���/)��M��WW��sf�11�Ì����BR��b��;#+����,v�3Wh:pX0c����ʖ1QbOIj6�ַ)]�\{��26d汁�1t0�.%rMn3�cf\f�@=�c�<6�\��nlޡ��Ȓ
a�f SG��ڶ7���tc1X�J[�:�)�C.���a-�K6�`Q��:�q&��J틻zL=.x�^N���W+7`�Zx�uy�l -Jk)Q���	��g��<i��Jr�\��q�';�X�p�.�6�v��n�rې��Oog��$v��q�ź��v+یR����b�A ���A��=a-s��Z��۱.㋎wo`�<l�o-u��"�4��g��{h�Me�Iv�9���:�}���-z�vyta��m�8#��մ"�Զ��D.�lQ�z^�P� mj�����ާ�rm��[Hb�;n̈́B�3g�y�f��gpic�:��n�̽�s��孲j��z���谮uY�3ah5�����c���[��!g����j뮻K.�97�[�����[z�A�s�Î�r��z�����.�Ħ���1��s�OY �d�Z�ۢ4�9���F�E�Ne��0��"�f3%�նj)� �Hm
>�y�]�64l�K�\��1�[�K���VZ{Zꍓ�wnO$�Y�s�DKvbs]V��s�#��!�nC���<�8�9�k�'�������y�c#���نt�M�e�-�Mˁl,mT���G��ŷ��On��8�q��9�c��VG���+�]d�S\P���J�n��<b���+�6���7��;n^�nf�68Q�n���6Z�uq��v̓$]E��k�����ݺ�����',�ۦ�7�΍�''<�G�P۞+c]�˘�kc���-n<���n΃vX�04�'�\��Ѩ@���ڌvMa���k��r�)���`���-�su���t�/F�r�ݵq��su�.�	]1BmY����I�fzk��ќ�G,��]�ݗ��K��Q���[�J�b��2�
���t��Gu��S�9��%4�i�s��
��N��n*^ss���������;��,q'683����������$�7=��Wb;gK�źk�i�Gm�X�04��v1����ـ,��sksp�KW-4r#���lpƻ&O];�&��\��3!N �.ű��r"4r��e�H[��:�m�n%�gIv��Ӡ����������Ħ���ym�k%0�X3�t8*����y�e�H�7���<�0�4+bR䣞Y6ff��F��qh�=ȧX��1�lF�ha���Xͦ%+�l�[4c�.��u0��mq��A�zLvz�kn.���]����k=I:�9܌���1Q�2:!&%��-��E�D��D�����\�kIa�d��IE�9|P�����C�A�H"#���J�YUr9�UY��'
�+�eA��J9�T*�Tr��97n�'!9DAN��Bt�e��W*��A'2��Q)4ʪ���ĕ
9O�ʊ����ah$]�G8%UHTQ(�����E���r��DL�ȕg.d�Y�(�
/=�̧]�jBI�(�M�MwhQ�]�r"���D�9��QȎr+��W�2"�!ʹ2&�eʉ�:,"��Q�5���?V{�Yt:�uc�C�c֎Pѹx���Yu��G��{T�d�>Ωz�J��M�����N1�-��N�Ɨq\���à��ߎ��:p��xܑ��x�͌�I�ab�܍7g��Dn��Tr��{f9�2;��\�v�ђ�ͱ�7j�
�	���z{v_a��c�,Ħ1�+��N\�,HG��q�̓if֑H�%0�we���c��ywOu��:�#`l@�\PT��kI�Vi��wNk����Fġt#�Rb沎ŗ�X9��+2[��D�SM�u����۷b�Z�����Xk�9]�`�고�\�m2Wu�<��&���\�]�Wi�FL"˃F��#P�+�R[��oc��dF�.�ҵq��\sCJ���\�qX�j�B\�HSf���i�L�*0����&qQِ���Z%�]]4u���`�`ͺܬ�ԉʸ����x��mӪq��;�hIr٢^1k��*,�W�xx�N�/+�kn�3��n��ʹ��-�%��
�mcb�ٹ;dĆ��##��.�
v�E����u?u�3����Q����=C�`��b��j�6�b�-�� pn:�"�1��ד�K����1p&�lh�:�'��8��KJ�f"�ɩ�-�lqj:bm�z;k<��m��|J��Plh͒;������k��릸�I.1vı�	��]c��-��o\���E�2=/����hf�*�B�v��2U�.1�V|7y�魌���v�R�k�9�Q{U�Cm·\]5���D7]*�`�k���\����*�:�n�������l$k�zC��K�ꗻ��x%�����N
IP�V�V�Xb�����nn�w2�(4�"U�����HA����V��	Xȑ���oQ��q�.C�7nxD	�br������U,-Q��X���K��YF�W�-(P�# D�(
F�+D�bA���H(�`��ן/����*�F���6�$O8O�v\��r�e�ݍݐL�@���&%!0'�e1C������n����m| ����C@�%��g߻j.	߬H��U'�t�@L��{�x��B�z� ���Rb0!(�>���W�;�$�FuĒAyt(;���4-�FKi-�}l��q*�&���ˡD��ܿ\-��7�F�D��H-��@��{,aQu���1w
#�
Q�10I���a�e��zWb�3Ne�u�}}~����Z/ٵ��Ewe
���bO_79V
�� '���?��
�A"Wz�=�<�߼�y?(��v��X��34X�:`pa䨮j���m�� �ײn�nGJh+"ɼ������:
z��R�u���=���y݂6b'o�j��$Nb(������Or�/7��$���W�5c'o�( ��t>���k���;��($�IC���(e�x�����8�P��٘ܛ�4
Ϳ���4���_?�K�~�H�� ���.����^�r�$�w]��$�$I���Д�3%��&���3��k4����"&SgW�0��0&��;r�
$wn�� ���t���Ȟ�����,O�9]Y�)U��A?��]!qZЏg	޹b�>6�r��FWD���b���+;u�}A�d�ʄloEc��IN�OO�&�H�M�	��aY�x���i���q͖�t"Rd�iq�T���"�`���NQ�ӂ_"��t�� o���9]�L��DD�2�)��r���7|׉�mвOVĒ>=ٔ;+/0�*���9@,	߬H��U+��eC�2N�i2D�$t�;�H$���{�:�^��w}3�k��n�d�R���\�p���^����T�ݨY���o�잿kk(����y���FWD�A��eQ�b ���WF�ts�v�P������T�Q��HIC��
��=W9����I �lI$����T<���{��@�ـa�$@��3^)�I>$��	�k{��TFTwi ���>$���8���Ʉi��6��D>KjD:� ^����w{ F�!	�1��Q[������6�Ae�DK���R��4�)E��X]U�-��ٙ��Ŗգ.�d��"��U�TB����@������3B<F�D��)�������Z	�4����b>�<ŉM6�Pnm��X��͘�������f��w{���*L��|v��ٙU㽼�J���ǡuT@6���o��G���	�Q&}@ľwd��Ϩoli�̪$���_��׺Ws��W�=9R�F� ��]0	���˳�1I�71	$�nP�|Ok��5��"D�� ��GETGR�E���|Ows�$3���3w��=$�&�}���P����6J��k�Gҵ_fv��)��({}� (g�������s�2�R��Hz�Z���f	��mj܂��}��;*$��i�Ԫ�;\1J�{�:<����Wf�)��CNM�xܙ���W�ؘn�'�t�y�Q�=sm�l[=�����s�d��1t*Z����ơ^���E���k�,�5덝�Aui���l,F:��ֱ]��]�1z��*�Ef�V�D8�]�,�t�yY��qZγ	Ct��\�	��Q��f��c]���WM�CΩ�)�(r��fÙa,e�QtΛ����TB�x��� �>v/��:�U��~Y6�Խ��������y�@ݢ���ʡ�Z�|{�·;z���d�|��X�Nu��`Q�r�!us(�D�Rc�@���fw����uĂI%\-�����c���z�(X$�\I�̝��F�!2����R���K��H>:�$	���7�o��8���b��`� DL��@5�s/1��xܙ6Lv7b�t��'ĝ��[g�X���%�AzHe��,�v����Y��qyv�mnY��LH�3-���d3&�=�n�=jA �F�]Q����l�TUp*���;�L3����)�շ��J��3kD�+�=*b���J�ޱ���׳d�L^����eۭ��Ǵv�د6�jbMT�F`�ͬ����5ؤ�I�˟q��+oC�`����`��K%(����Jg����GL `~yw�*OL�A>��	�����LX�(c�Ak��m�ƽ>�Ӡ �ln� ;;�	vћ�.� W�¨
�[w��F�! z�S����E���̠<s��˪�ݗ`�a�(p0�(Ĉ�>ۏ��ƶD�ygp��[/4!1a������}�\��aMp �ﮨ��{*�.l�{^A�C�B��0�Ճ����4��6�^�����ٗTH;��V�J\5~������������e1@�e�$ߧ*��Aۚ�G�4Zeq��27M��ly��~��U�5���n�2}"�����J玻T�C�>sZ���I�|�=�Q?\����+J�g��U3�.gSS����� +sۗd�ڸ5\٬�Eu�FG)1bD�TI�Q��ud��ڒf�HoH�qg8+.�� 7ݖ,��ړ$����Mp��,��9g<]]=*���&8��6Lv��&���
&�52�!���l��w*�I>��	k{$Bݵk<
�ڠA!�n�$�8�	2D�&��D�K�uG<"�8����:�k�ۻI����� �]�R$�Ј��y��-#���2I��z$ ��t����}K���I$9�a�I$�C�T��2��@�!MM��9��q����tA*u:h�I%�ښ	$��yob�3�k�o�h�螁���z�߼ߛ�����%���k�͕q�)�uCF� ������+;�K��$꛻��=U��		7j��R+J��_���4I�g�%I���^��&�/(���4�-�I4}��!��[��3��$a"�:J��ѰW]�7i�ES*��>�fdLS��Lp�(cϕV�7�i�K��B�H���wa&,}1��{���8$�@?_�lη��!f�PHS�׶Hŧ��vq�-|�{� �� �=��	,e�<!��������$H�2n�(��Os˻%y+��g���S.�H$�GZ�E${;*�#��l�������T��o:��Y�$�u�4�	>ܪ��	wl�RFB�,�F�4n��z�6��#H��Q[���I��b�(�/_�$����I$�n�ݢ�K�i��%�S��wi�
����W����&5�Ujg02�$偑�Ӑ�a�rPQU;Ж�.��:4��['Jʅ{�;rr��"r�����A�xUY�kP�@���UeBV�$�տ�G6bt��Eў]�]7��\m��<nh:��K�lX��wg�HS�K��G�.w�Y�ö2]*���^�����2���6գ�!� �]��tC��듶knǎ��K硞T��ˎk�^�F�I��.[	�)֣-ە���4����=f6�>��&&�@Lh �]35�E]]���%���W�% ���O�_��II+�˻I$���7`$�kw�.��TA$��dc����$h_�K|�H@���q�m�L�$�f�$���>�=	D��.��=�v�3췉ZB�Z���	k�}!$z�L��h������j��D��^]a$;�Z�od�"j��!>��K�}}^��h�{$��7:�ߒI ��r;d<��RK3.��8Nk D̤�����h�Ŷ��4.*ŝ�.��H��:��H$y;M�}X0�X�J����i$.�*κq!͵3��;M9��̎�⮕�������f&7����HI$�߰ʄ�I>����xLc�ʄ����\$�U��Y
�*ҥ!��U�D�I6�Y��m�rS��;6Op����V���Q�t��yf��6��Y��7.Y���N��`����l�0�C�Oj�� $���.Q$�}{dP�c{��hk#Z��^R@�6�z�UN�F�I�;T) �9�b*�=�d(���.}D�<vϲ�%i"$J�*�U��d.ռ���	 �To+��A%�֪�H$�s���5�Pc�m��ji���z����HEZ��g�I�G�̅	?\^�!&��G/�l�	��$���;�܉��v�vA�1k˽P�g��L��N(B�K��L+���ߥ��	fȒ%��'��D�p�ɢ@�n7(��Ye*���wNr�	 Kc�W�)d�*�J�+MB}���H��h���9�5b�H�����D��˻D��4�`Y4͢I��=VB��)U�F_a@I_<�v��K���� �߾|
3���?��h�VX�㩛؈1 �� F���>�v�u��8�w3�oNr�f���R��V�vMv霁�����a���d��i-��v��y�p�Slmk`�ٜ�Z�-�Ui����$bVmMͰ�#�tk,���8]���j�j�AY<�����/M�2�q��W�v�s����Z�z��w��+����O,������J���QM���3��0ܘ;
�ʮ�aӇ�����^�d�I:it��|q�t��v����d��<�v.P�_[��M+��\u^�Z�g
�nc����R��̻=������*Y�e#��d��`PV_m�f�@���2e�;%)|N��!sU�������B)I9yE�NW�Ɍg�'R����2�\n��Щ���n��H����]�m��.R��oR��#�ͤQ�Y����hvch"�8�<)�]������8��/:�Xj3I��C.�.��oS�&��|�-f�,�V�s34_vm:��䏒MZ|��ǛJ�,_.g�j#,[;���]��n�����K;^,U _'�\��֘��47�5����U�je�;#|�u�����9�jwv�V��VHr.��l��d�f�Ӑ�af���{�p�њ�8.���%��Ȟ�y�y{�<w�Ƹ4���0R�9�!khf��zã�׏�ҙ!I�[C�<��UJd$���L�����9:uR*�g((�V��AFa�@��p�r3**�"�2tFS�d��T���DEQ��y�HE�\��T�$�rH��PV�*��T�΄UUʡX��N8W(�M�Q�E��*�T�r(��][(�U���QTQp��\��$U�(�\�AP�"th�X�)"�D���"��e]�k%�B+H����t�F����dsP*��k,����ʳ"���K�s���9p��+�PNy�.}�nxTPQI4��W�]�vDD��n���RNGy$���iw2+w<B(��X9⒁r���#1Sv�(�ث	x�'3=�$nQ��]2 ���!5���H�M�H[]��'z�i��	$��[$�TL����!���_ven�{i�R�I|;󚕥dժ��f�>�!�I?�_a���cޠ�k�'L� ��rHA$��a�%V"w�]�̛��u��R�+�wJ���`�:�'%M��okr�:����h����-�v�o���"P	vvX�@$�HoN��I������\&X[�R($��ˣx�ǀ�B�D�.|}���@���Q�Vb:�$�>ܻ&�K�w�I)���,��.��6�V��O��*BI�'6�� �C���N���o	$�����I��a��O����]aY)U��Bc�g����J'ݠ�(s��v%.�dW֨��^�x��R{%�^�KE%b�[�7:�
��Uu���30Q����Z"ޕ���b���[�"�TB���.*,�w
��K�>����t�@�3)�Lz�*�����I|��({wt>���	/T�]ߒ@$�Y�i$�Pn9}�Z����y�g,=����4
؛$�/]nk��&<��4u�l񠒥V���ZVMZ�(���쐒���n*$�H.wIm@�#4�z2�juۻ���Z�q]��8XRd�
L��>]o�@�(^�u�2�xN�6�I5�yv$���vU��ܹ݃f0��b�"bRWz'�H��I�H^Cmӥ�by>$����J$O�[�V���6�V��O�۬{���\A)qx��I�w@$�K����x�j�L*$�)�BO���tU�e*W~J�"�$�J��W+�!C���eBD�^�% ��̂I>������/��x�gU�/s;Wy�En��O�=o�-��`�{���\`7��ҁ��6�E"�2����S4Ï�+���^z ی^�{z϶�:����ijnk;GKV�l݉q�B۟.�zɺ�Ο\�9��d�(�pv��c�[����l@�zw\��c�]��=���=tۖ�l��{B�[hjy���7�ݷ���J��y�W-���O=��i5w<]6���Vڂ��3�&��Q�n�K��.N3��m.�!��X泺���W����^A"A6��?׸�Mh���TJIw<��%�1��8���o�ڻ�I%�w��&�ĭ+&�U�jO�~{*BK�m�x�o����2�$�$gKO�MOs˱h���#��f+xz��"Q��a��>]o�I {=���s�t��h턐Ix%��H���yW�k��4�`�c�K'��*��_��@z�RI ���v�Ioma��K0*�M�2ix�]����j\'����ݜ4bW�q.����(	[I$��eX� k��BwfV�u��� ��F�LH�i(���2l��a�k����`�i�:9����`0�Дȇ�J�"I$�;b�^��v���g�gsÑ1m���G�r1��I$R�1�3;8v�5�R��!<z}�΍!�ra�\.��T��J����Yw۫6��k��_t�^�䷙�{����C� ���$$�˰�H�b����sJ�̙��V��V��5!/^Ϫ@	>��	$�jݻ׾3�7}�$���IwN�Ic��&H�`D��=;�GY'I%M���䷣q9D�$��<,����$�|�$�֚���Z�D�G���P�~$gKA�[� ���! {����$�O�Z��go������'e���u�f��έh�&G�������UG]3���}���v������������ �I.wI;�q�{�Ǌ�$�O����~� �Z�����	^�U$�šr�8�;���$�H>��'Ā�[dV��w;��BkV���H&п�-��!$�G�[dK$�^��v�8���%G^e�>K�[�<j�m��^Vu�R�������z���9X�_���D�	*O�ͱ����Iy/�;i�]�Y36H�VBQ/�H��������&��ՋH$�H&�(�I.���H�*&sA<B.u����t!��L�&.I��`R^I%��b�5$�NF\l����'�0 %�B�~>���t8=�~��<�vO�c�S�T�r�6���M�gOv��ّ��;YT�R���x�`mX#��ܞ��&�Ib�T)$��yTI�|,5b���TWĚ��жO�hov�Ң��r��s�%g�,X�ض�֗�A$Fڪ	w�UI���6���J3�DBId�W%}�D�=�$ �/����v���+{� :���I��ؕ���H&п�J�O�\/����mW�$�K��U��I��W��T����j�����gzQ�r���}�_��xh,��˿]�+Gc�1�5� �%(f�VP�u��[�F�{����ڪF�S�Wi-U��r����=���rq���ɐ��U$�G��]��Kzwߠo߽�uu�Yw�
�D1��<��6��j��/c�V��\Vn���n+��=zt)N�e�v�I��qU��^Ǻ�*�ܫԊI��ش�q��&T%DK�}��ϡ?���^�/→�3�HI�}��,J�(on8���p��&&"d)15�9߮�@%�7�%%��$����Iy$s˿E��]�BE�����AR�s�/���^f׊��!�I&���d��I���z�[�c �6�G��ϡ���Itm�״�'�at����.�������٫�d���װ��m��|�)�4��&M�3X�3��)/��D�΍JO]�E���om�vM����������O/��ư�^Q4%��\��͚���oH����=�{Uj��\O7��<c��B �C��%�͂�G^Y���d��b�Y�/YH�K4Wr��f�q&
Msa(��;b�ٻp��딓W���Mթ�gE/dw�;UF���M���k�]b\�Xy��jS-��Ơ�ȴU:����&z�h�h�a/v�Z8�@ngUz��퇎�k������_����8nq�J�mݒ��tn*6�It;U^K�h�^{|S�Q���g�$ ������C`�"L\���U$��ll]��h�I$�l�+�I%��I5��ⱊs����ݮ�b��L�)n,-馬ZC�$�m��I@�X	����$�y~�'ĀO��]2V�>�v�%A��	}��#���F��O#�X��%�j�$�H.痻=�g���$���VD���ٵIR�����I3ے�V�Z�"O��p��$�r��A$w��ọ/�e��a"�~$U�+'��$]6ܕY�p�rl�V2���>��M��w<��� O���]2h���$$��u�N��a�����&��D��Dګ!�����g_�J�_n��a��Ǫ�X�kr��4�3^�v��&���\*�D���j���$�;1O���wj��_ZI �q��&�Aw�.�h�7춢�8�r�g�B�]Z�����I�;.��[�[�ÊW���x$JN�$���ݤ1q��&b�7����P΃9�0)W��� �ܪ�	��nQ'�O�ݗ;�S�� Z<�]�}v�$��>'�� Iý�!���:3	~��UI�ǹv��K��"�ȃ-{o�M�K�傍� �v���<��-�l��t�ᗌҷX��.�:m�~y��:mCh��������yUi$��~HM��1_up��q���I$�eش���ȑ ��>.�m�M��.���r�$�$��]�a%�ۑw�H�X}����o�NS=��e mU����{*BI'�}�B$gKƘ��2��`CQ��?:�oP:���Ɯ�DYrP���;I�u��L�o��緰5H\��ԭk7�o�r��G��&�K���d���bh�$@�����=�A�,^�$��|��i%�{=��$<���Y����1��K{tt�ȹ0��"C]��bI�п��"��>��ē=�|I�Mg����&��}{eص=	�al�����:z��mp�i��<sc<���k{�v�$���>���~'6��BRI.�j�+t0��{F�n�Z)$9�ᐓW}�UٵIR�����{X��]Yt�v�;�%n�b�I$�C� :%����4�&�/��RT�h/��-��!$����P�4-ZQj�y���=}��>���2g�DU�DZ�B嶺T��iUQ>��2I$���T�I ��[amv�O�M	�gf��y��7:ޤ��t�ǅ,��E�C��Pd�з�C���ř�݈��#mf���b`�s���E|7	?{jo�cGB��H�'��t�I�����]�n��	+��!&�'װ�$��$���M�,��_�mX�vMI�����΍�Y�(�L�����V.R�~������V�;�w��!$����]2I ��$��u��C��!{��!��TI���T�ͣ�i$� ��O��>� 6Ù��w��BI ��$��nIP�'J�}!��S�~ω7}Ы�j� �JJ2�I$�W�*�$���UN�bI�TV��	!��ڒI;���^�ꁂ$�m���IS���&����$$��˻Ix$�GnE�g7���I��]2}�"%D%D�R���$�v[��]�ju�J��d�G��lo��"�, |�F��>�M�F	�Q��Y��j�=2�VҢ{q�kk*�vD��K�gJ�>�����VˍԘ�Nv��x4kԇjuS2���f�]+j�<�,m�c9�;�eJ���%�Zň�j�a��7-R2N����Tfe�j�S���h�3�=_ ��8dm��
����+�w]A��w�*��׆��s�g!�J��^��c�aś��j�v0���;��6��$�3F[7��\9�$�lV{Yk[�N
����84��1�u+�xӑFN����(���WNV�C)��Wk���ܾw5H��Ab������f_vj�����@��f]�����j�kr&����e��U+��>ZM�2�җ3�1�t�T>��[�)���������7U��L�-ԍ���7S��r�c'aUi�^�]�(ZS�ytn�Ź��ok��V�;Vr�5�Z֌�՝st	�-<F���Ա�[�+�z�ʾ/7�U����fN���`�t�:��k��}ӊ���3nD����w�5%\ne�Ձ�W]_@y���Vc��;(:-�."�̑�	�eMN9��3O�k5Pe��%+\p�ګ=t�'��rr�zcW�Zu��%0��9�t�6�p�|�㚖�T�gN(�α֪��/���os/=�n�!sHmM���8%r���[�"����s�Pz2��X�ZN��;�W��y��2d�OW8�}�w�t�*���:�
bCϟd�Rr��r��r���Gr
"s&S�gw��V�GQ�����#���dP���Tˁ�N�)��O8$���hT�W�S�w��2��:��9����t���v�]�"���C̢rO!���s�o:t���T^��X��s9sR�����2�1W�	�܌���,����'�t����G�)蜏��P�܏S��@)z���&���WL�ddZ`�	'~z�ז�i��m)���:���v;�n1��Yny(�åw���u��.�d����l��:Xb�q��uooi��U)4n����� 鱪M��i���m3c�]��s�n���;q���ަ�v<��Tc7N�χ�@�5 �b�,K�k��3v��\u��"5�i�)�a����3a��帏%cqk�2u�R��C�P�*�����㱨]��:�c=�N��A�Bڱh�cV[lv����<�QQ��t�\r�i�ܗK�.�j�4=�t�y���=i��5θ�k�9t�s��ѭ��k��K���nqb1�Z!eV���蚠����wKˌvu�:���k��ڰ��bL[�n�p�\�-F��,�;���է��\��
�4ɢC��iJ֭���m��y�2&�nN-��c�(���q	���a�]���i&����s8��7'�*@�ݍ��&����GF��r��Ľ�N�d�=%lv������`%�#p]�]H��b�aKE�)�]��
�t��pE��ּ�U�z=�ܳ�k�\���]i��>��S�pg�Η����8�%МM):��l���+�*���������8"QV�+(C8���2�Ԁ�q�1E.+v��dy�8�C�g�mc�v�3�>��b<5u����`�����I3jCY��h�!����nT��x�|s���p��簇7�t�Ӹ{-ڨ���znBn͘�\�#
�,3���y�h�ڣGQnf�v`2U�qV����b�]����R�Zi�"�5��vk���&���lö�N�ځ��@C��p�75������ؐ:ܞJ%0��nŸ|Gn5l�, ����-��Rk��){-�l�2�=ڎUr��Φ�3���pF��pf޷�q���;AwC�&���]��]Ss�Lu���\��.����t�����$Zu��#�q�0����[� �f�F�S�g��Յ��8��/mV�h�W�@�3���~��Y��`�ܭ��b��OT��һ���˳4v�{�hK4c������ ����<DA0:>�i]C�RK�I7�w�X�1�d1"E���- �Sb淎޽�9X��A.�VI!�ݗ!&�^�즷sr3�[�z��I$%.��nIý�!4I�oxk�د�~�
	'��	�>>����j�ڰ�)R��/��;�u�I?�sp�I���$���!�tU�o�a����'��*^Z#dA}W�;P����U'�ˬ�J�V�>'}��wa$ގ�D�k�ڪV}��;שü0kǡ������c�^�E���0�Y�%�ض	v�Gc����Z���0���O�����OĚ$���%��v���Zc�m%���VNV�2� *��m��$�;΋s�]6$D'�]���
3��e���;f�mҖ��Ǐ���jhI�D�f�3��%�N�<mMyN��Z��{޷<��$]����$�?��H���qw,�ǹio9�dJ�D��ޚj���@"3��I$�>�L����k��I$�.�!$�O�[�M,�=v�$���	���PJӉ$�8f���Iډ��	$���i���]qFI�nO\LB�2@)R����t�$�3ے���Փ���䗅t�D�I�j$�k˷���u������)�ڷ؆��y�1�E�;�h�]�5��f.U$�i������.ߊ�4H�;m �+۽�vǧE�H]]Wq�â��� }��'ܲ�v���Q�(���<�'-�>gi�	#��2M����IFڋ���F��LTU���yv@
��\S�u�d�I�{$�&����g6\��P�`��d#1�z�����뺙 ��:�R��E݊��WMIw�GrW�J�4H����!���=께$�I'�ER$�}�]���I�B�jIp�F`��hI$k�I&�W��vA$��Xz�(ј�8R��%]���ۢ}9�j�I�K�����=	ۉ��	 ��]�h��v�RYڳ����"`���,8o͇�1��g��]E'(k���oϟ����u�j�dӸ�
K� ��˻^Iy%�ݱTF�}����'&�d Nwdb_y��6A������2~'|�[]�!H�S ��]�a$v�PIy+�-gd���W��m�&��.iZ�$! ^[�@�[�MIwK�y�}��o��H��rh�G���&Vܼ� ".�\S�}������f�D�<�v�%.{I$�]9w֕;��{���aD3�#��������v��'o��6�=�M�\*�(ًɺ��¾���~H���Wk�7�T9Vh]�#����d ^�L���gOE�tL}�ω$�=�[d�I>Ym����_�ΏK?WZ+��Ղ�5��V���u�g�=l*�+T��Gn�i%h��ߨ��kp�o]RA"OND�Jȴx��iĞ�=�HA�I����=����e|��	�d�R%E�C�ռ�O9�i"PM�U� ye�d'�^�d��r��ތz����6A��߭��$�<���xg -�E�6}�o'ĒG��2I ye��5�YxhI]�!�oN��:�+��H��I$�W.(�I.��t|�*$�s=m�~�뗗dEի�|N�{d���&|I+޶ �ue���{�$�L����׮��ҷ�.>�+ J$���mC����	i���)��H�7GF�U�d�ޥ��s���uy�OZsB�M�Ѹ�қt+����K�P�;�ٻ[T&�\�t�sRv�8���y���ˍ<<`�-Q''g���}��{ �p�Vf�Bx�T�&N���H\�v���G�)ΙH�����!�4p��m-�)�ɩ�]j��]b�ǳ鑋3ۄ$��i����AY��j�ʼ-�Us�c'�U��8��Zf敝�L�����gڱ%]��p>����i$E�l�h������P�{j�Jp+�=��tI����&�Q>�RE R�Q=���%����E��%Gא�%䗒KV[d�$��I*~'��˜�n���q'�O�"�ʮ�R'Z�O���n$���c�(ʊ�' H����PI��%Bo�� �l�h/�	u��.<�f��	����I'�ww�H�lLp�<D�{�*p��[d�b˄j����kvT���#��雪��o["e�%�בU�H'�.�^�b�%�����־�ޙ�����4�6��YßHm�",y{���D3�+�����+n+���x���p-�.�I$w�$�8�t���7H����tle��0!!�w��M���w^Cͥ�A��Yl�]�.��.���<�~��d>��
�Jɫ=��®�.|J�Y|�p�|���V�rk��$�n���Ą��=�g-���r��$�XC�\���h�m"�)`y��I8�$�K�5�U���̍�$�Y��`Y���u��'�����-R�'�L�����锰�KOg� h���O�OĒ}��u�bgkD�>�T6}� 6�ػE|�߭�I?=�О�囋�UomݤJolU$I=�K�8�lV�'������1K�h��0���U#)u<��)k����v�@����Q���[b� ��G{bC�@'��b^�E����y��B$�{�T�ÌɈ�d�1rOK�)$Op��K�Ok����`:$��v��W����X�06';�;Ho#$��ڢ"�O���D�n� �<�g˭<�]��ٮe�^�rb㰎�T]gyW_J�.VS!s3U�wV��BoF<��3�n�Z#a���}�{��ܿ�?h��[tI$���Ve֍�� +w>'��X\�di����Z�MOk���	%��nz�N������D�^�4��i

�R=��d�h������g��|ݶH����Mw�J�-��������-���9NS���-��͸uVe�����ύ�u��{���aQ��@�x���~礪$�	v�UXKn�Q�Xf�9�Or*��$�3��u�Yp�6���BQ/�[��=ة���'��%�QTI�ʿZ+�#o* �!^�ˣ�a��Ɉ�d�1rOK�I$�K����+�tI�4q�11�$I6�*�I�ʻKs��4.�'�w�=�Mmq<�{�&D�͊�H����D���̑cc��4QH���[=���^�L}��v9���B��/��z2E��ʔ��)�{�������䉻دR4�xś�I ˄�~�RI#w��+vp0�0��I$���>�$�{��}�ۯ%	�e�u�e�i]�
�j���716����xX���>�7�=��L���W�I��W�.��K�b�$'�\����[�(��[dGgc���Zl�K�(���2IY����D7���I��I*�?h��ۢ@��K��^2w��������=�R��;��I$��q�!Zĺ�x$�Ak�&�H-튤��8���I�7亜dV�uW$�swv�I ��Uy%�K��vb�OSb�	&�uE�^P�ud�DF��$�"s�L�@����@��(�I;�lI��c����,P޸N�T�dSC�^��i��Mq�L��>S�ms�c���۹O{6��ʍ�Kd�y�X�wP��_�xx��٤T���;u�n}�3�n��U&���9���Wc��!���ب{;d8��s�t�ۢ�nC0q��l�*�m�����j,v(^=P=��;F��B·X9\�n���i�0�͵&��0��<��v�8�s�%�nwP�uuu��=\�S�lO�$��j�g�mk�(����wK��u�\�n��h�f6Y�Kl�k��'7e�n�����A��J�����wh�GERI$�c����
�c�cڄ��Z�sg��+��%;-�~%B�.ל�	$�G=�� '��� ��E/��J{c��	<��	*vR_@��$�	ʉ4��Ac*&˾]8�$�'w��$���|�@�j�HK�۬%:��"Q#=-TH�v�($��˄��������I`qy1�&.I�p�$�;��.��;բ�G��h$�K�c��H�A>컵t��}߿t{������D�p,X�Q�.5Fb��B�]%�Ѕؔº�3u���KWB���=�ר��n�$�w��%�`ui靣�- |Oy�dҘ��V�Kޘޓ��<3R�g7<�������E�\n�;�T��']7y�Ѽ&ܤ~�8r���o^*!X1�)j`�m'(�s+��$�1��	 I'=��	!$����A�o�/�#^7y	5�l�D+J���r;-�h�D��J�� �:xA⸬�K�$��W�W��eѵ���) l���\�f�w��l�I��RA$�ܪ��I��W�U���$�e��γ� l�f�8K^��&���u�W+":(�}�m�&��s�������l�x!��X2�ؿ����V�����N�ƽڛ��Ǭ�s��ti��5�߿���[����d��l�I>��p�D��Zd�w�>�Y��g�Ku�ش�<t" B&"B7D�LIi��]U����U%�Hcܻ$���:I*��d1=��J[%S�
�P*\���l�� ޴ w�ʾ�\������*	�b d�̹���UG.���휲0{Y�e������μ�[�3]z�r|�h%R�����S)|���˥��F���ˍ譱��4�w���72v��D��E��Y��H��|^=�$�46��d���������T�8$���u�e\᝚t�e��:6
��J�z�g$�V�Nl��\ܦ7��{;Ok��.F|ڢ�vhn�q`פ�q��&�Zoi�d\\A���/�'4��<�7�FTa{`�c�d�F�mdz��y���Mvswkr�]�K��`m�_`���.��QQd������T��m��U�F�CK5_ %��o����l���R�40��]��U��!��4��=7�F�ua�-��v�L��>�Ŗ��g��s��
P�E%[�4Y���gD���u,T�ύ�6����n��o�a�p�M�w_�l3{�C��m�Z�u�Ei����n�2���ٷ�O�Gv���eM�B�T���`�:u��ڈ��mj=.�*�_Y�5��vF�nne�gDҰ�r��$��S{��37b`6�7O`o2��WP}�%�7���$�hV�c 0�W6Y����i�n�N-:6�іƘrJL��[yv����nfK�t����/����ᶷ�Zr�������4k�8����e�:�Mt�Ӽv\��>��iv����u�U$>�9T��]�S(BN��z7�ĽK҂#�4�ԡ�
��dA=y��i���p��R>TkTZ�bl>���L�!ĕ(�
C���'V7�*�R�4<��w�prkE��'o'�;&�rb�w9Ar�8Dhh}v��/"
(
C��C�	u#��QjO$��\\#�	Y�H{�!*���d�2�W�c�EM/=̖'^���D�*C�Rr$�	%H���a�$�˗Q>���$�r��H��汜��S��V0I9���&�*�V��L췑�v��$�L��R$J]�I �=��oTf�e$�ǷBQ��*����� ���Ϭ��J�tp@OL�I�� �}�����o�4�䤷��K�4�e΅��T�k�D�0I�R8e�M���{�M�R����]ݯ$�;�I$������P_!sp
��!�4}�ꉕ�b��F�իh�RIR��jqa�Y��I �[�I/$�쨒Izf�E]�h��ƷPb(�.��}�n�d�I���L����ck���Z��i$�2����P�wa]*K��٬xYlr��I$s��M=�lTH�{pv�~�tу��о]�on��Z�e�څ�'fC�ؙ�/�1���(�o�	�j��֎n�ʹ��� ʉ'2�~�I�*_IQ"Ę�k���@%��]���8;E7��$��m�$�D�;t�$���I<��N矽�9)�ڸĺn9��b��c��'Ƕ<��c��뵠��%��y+��@���&?[�@$�c�L����BI���~�{���ĒM���x'���4BBm�eHI�
k���Sy�z_n��Mh�G5� ��{� �%�wN{޹	�/�D�I�TN��$�{rT�s2��3%J�)�a$�:��I����1�B $LD�n�%�P���EO7!� ��2I ���H�I�u��鹀%��&��ue]*K�O{6}R�G�RV�����V�J[��$����'ЃD��Z��t���{�����{��c�~u�\}�v��CSN4tɭ`���;�t�܀x9x��֛�q��@mGǢ]J��u�ӌ��@y�S��WKC{m;�lܛn26���Q�c۵6,<dݜ!9�c�tGHhб��x�1,aq�m�2�6�^;f,r�f[2]����+�$�ً��K�W��kc5���҆���1l�j���vl��k;�$�O:�����Ժ
E���̉)��i㘆�V\�`7CAw���6�`Λ;�|>��T�8���I���cp�D�>�[d��|��h�ݺd�n'@T����IT�>�����a�`�*s�e0(V�F� �m��^�o�J ٴ�(�;'<I����OMNMk�� ����C��@:�K�f��Ҕ��	��:o�z1�>��H#{*Q�c*l� �љB�^a�B"B3@�LI>$�����؈�� ���$�{�����
���s�4�[!Þ���9��dm=��r&@�r�b���(�]
`H*p7y�A��G��oeUx�Bg)� ��m� �u��5o�l�R��cӱ���xgX���k>�P����/K©P��b�ϰ��Ol՟o.��F�)�<�4ۛ�#5�N�`�mi*5&2��{�xUs��|F=� �~Ʃ�z���	8��Ce�R���"���� ��eP�D���[};�(=�h]�m�W��AF�A�+�O%� ������
 o6� 7��kkޞ��(w����x�� ]ZR�� �u걐w1�]�u�R�H�ʪ��u��W�p����LJG3���l�O������^�T��Q�dL���/�_faڢ���HW��u@�D�U��l�]�	]jI$�ꚋ�R��)� ��;��Pp���ts��וT;�uD�,9�w�UYb��)+T�/���t�#3��I��"-�U�ȓ��	5�\��#I�c]�?���9�+� vج�]��؆VPS�0ڼ��'8kΦM�@K�Y�����1���pao���nѴM�R}�NnӖ{x��@���H7�sDj����\Ěxꍎ����$d�R�}ǚdB��޾LW�v�	�n��ysRt��i�ɮ��N���-s�U%͖Ye�f�eS���<�g�H�Č�ލ�"I0"f��r8�	�ŎZ�١�w7@nz*�d
���Uag��@U�h/E�z�� ��@�N�hI�5)Gg9��-	R�k�A�~@fj�_P�]�7� ��� x�J�f�.���J�$�2�DI�o"=&5��'�rO�_W!Owe݊�l����.�d��y���9,���k}��g�E	Kڊ�֜���n�7x�@����#p��3Z��t�����^I���*g^I$��ty�5f5�zwj�iT���?6�Z�]�R�H����N��$���5�nn�����p��tZx����Q�q�5�r����%ڋ��,vn���� �$�ޢO��q �A>�� �OVntp�4r�j�';�|Mˌ�"I0"f���(syE�����c���$��UW������s��m��Ba��dn�`$;r��� �s�{�%Π �t���ڙ@�#n�ҠUX=��\�isE���|H�U@���PO!+D'�֏�qp�1"�ĉ��דD���T��"E�$�$��U����)[5�k: S�.�rT�2/�$*����ㆹ�fObΘ�fZj)�f^��.<���=�{���׳,���m]�M�ʂR�;\�ډۛ��q�Ҝ�Q�)�(�-#A���SjK���!�&Ѹ�u���`u���r	�������Q�6�kh�t�OB�o7GO<��N.N�E����A�%1��n˗tˇl��\x�j��Zn�p^��f��gv��S��g�Tk���ꍑ\۸&�ۃp�2�z��u�n�sAUՎ�4eI .��{�(ݫ�M�[��С�s��D��5�\]���f\�V3�$�k�������$d�����\�+��AΦ�'ݽu@�o{��GU]@�����V�V���� �lL
��-Gt2	mԊ=�sF��`���b r�P����A�UT	=�t(�p8���#�=[5N�eQ��R�\D��H=��N���hW�9�#]"G@�)uD��sD���A�Q7�(
�ѰJ˾vn̒M�E��x�v�;�Ȇ4d#,n�-b룦߾�g��J�$E���3���
���ܬkDvW���*bv�Oz��Dڲ���AZ�ڗ���M���+���8B ��c-3�!�[���o'+=�X��Y�q'=N�ja��:w�Q.<a�����7~M������ݠ(oܦY��5���XAZB�0��h�q$�An�^��1sї��+��� ���u:Yϭ .�'>�s�yQ�[Ñ窼O>�$w���h2|*��u��D���2;b4	5�UA7��BjI׵D�q�	�$�eP��|u�}���{� �G��vi@�9LBWYT�Vvrܚ����]1��w(|_Dش}�������e�@�A#�*�*�w�'���F=�$c��#���Q�ܪ �Z��gM�О�
��Ă	�ʡ@�u9�����:ަ�6QVm*��~��B�1� o�t�_�ɺm�r��U�D���q�7Gt�b��4rbf�K�h��2�����U�֪]��"��3����� �މ${�n��y, �eR��^�>j�K���Dgd	 ��U@��]0;p]i����h:�K9��դ�G�Ъ���!�i�^�w�e�*���΀�z�6r�����8�^*y�8DF�7�:�f#3iiq/+��48l�a]t���ߣ�Q��ӿ�}U� ���yJE���du��JZ���i�̠O��Dr|=��2�k�U�a �kMx��sD��˜o{޺{U�������� &z?Q�>$kAa���4�A������߀F�fҩMu�Tj�N���_�����z��F�TF�
˱��n���s13mX���F�%R��A��|雽��S�pe��;^�q�^�g3��~�3z�q�+תq�KL5�1�P�	}�FM���N˭ܩ���ލ�B��h.��;�� �G����սt�eλ�4�;��t`�e�T�����]�/�2H�5������w"���q'#+�}��נ�s�|H��P�jp���b"�zbH��9
n8��c�<��'�Ē�wyM�qs�7AK��"�{5ӡT*gZ�zA~�^k�2P {�1^�����ѴRV���圆*�wH#g��A7�A�W���<Sk�$��� ��Z�iS�?Z ����ܐ�[�e�A&ۉ$��c�y{1�[3�y���]%KQ�tӳ�W�A��C	�U����C�1B"
�;j��*�MO�Xܤ�z�,:gM���{ݼ7��p�}Y�wQ��Lǀ��B��I9�����C��y�]ne�}��E��PJ=���ju�ƙ�Oq�1� 8ԹG�v"�eH��s5m�0J6t`�}�`KEܵ�QSsf���=[�ӬL:�,xC��(������0)�ܽ���-����Ks���^����j�v'dFf�<�y������옵n
���陲�G���Ş=�^�u�<��Iݬ>D��p,;�u�kF���cW��\މ�#�Be삮R�ug�r�Wجyu՝R�zs����󢦖�$2��6Ⴣ�pZKE!3y��w��ˢ�à[��W�b�圞��}�5�rSe^��8���w�����l�'7�
q�/~�o6��r��bٸ)��fXk�������D"�sGk"a�y֞\����_#����;2+��D�����Â�q���ʕ�4r4�:;e�|��uvIZz�{�Mn�˴���ƑJB��NK����M}�mӄo=�
��+���{�6�X��7�m��ɴ�e��2-Es	��
���Ƹ�ő��
/Z�&�����.B��Bn.1�d����V��1`�s[.�O��%IQ�o��v]�a8��r�Mo*r)��]�����л�xE��W8��v������{����ALYޥ9�<��,�Ep��s��9r���W�8ӧB��:��O!�N�n��:͔�e��&����:���	0�̊�M�H�s�7;�+�9L��i:q�)�'��&Oz���rN\�v=6$QA|�&kԾt����o!��i��
��<��V��NBA#����CT(#�t���ܒDϫκ�O��A/��Nw��a���iʡ�\�p+�)��y��/����)��e��7+ʺu]���S����M�p>�)q��=�t� �.ck�K�������өv��j��L�q60h�s�P���eiŐ+0�;q��;Wn�;8�����1��˦�Zl�b[�4�;e�*5ҩpk]gU�X�z�m����	�5`123^Xs-k�PLm�Ŷ6�k�ܲ�h_i�5�4&�W7I۟��!�2%:���������݀�VC|�8;:��n�m��#��ӝ��Bv��Wbةa�--7B���#f�Bʙ ˎ�s��<�M��A���jum��5���f�y"�Fn��N�^v�����gu��&�tݳ����^]�+��;nW>l�-)s�Қ!0�	]�l�=���s^�{Ւi=����y7�n�'b ���a [{d1Ѻ����Z#<���c����I�w#���s�JN9��v�D4��9��IEYx�%2�
��/G`�s�m����4V+�c��M�.�$#��jg00H�%�LE�CK�3��ˍ�6����D��ϛ���H�u���"����b�
V��K�30=n�<�un�B�c�݌���=vV�]�G&���oZ2�b�&8��Qv݇��,N.pi�恊Tte�n�c@��4B�m�J[����.��q�d��h�=n�l�� ����j��G\�8�LK�-�i˦Bۦ(Lq�W��rz|�\w7*�\k\s��tME�����2���ѥ:w]u���M+D��k�hכ�֜2�yK�E�n^z�T�cU�fmj������f��jz�pnv��n��I�V��a���M˱N%�V	1�f���S�����7XѴ�7c�0x̺�lAs�ѷ'��X�.�$�6�Gfꧫxչ69��g��[կc)��E�X��b:l�`�&S��pF�33�����3�#\�+����#nɸ�C6��L���&�9M�:����G��Z�`̎�ۤ���e�[Tb��l7&V�YC]m&�ۄD�"O;�\Oh�Ѷe�Lݟg��������Z�e|��Q���ۥB�{b����V/7���
'���̘�"*��yC��b����1bkϢ���m  ��������|�n�o��Wh���r� ��iЬ}�tWm����Ay�&�=�怆�I���%E����g����!�H �]�4H$ou��;"cm�wD��y"c"JE%aX5{�:3=�|���>�H�ʪ��T
0���V�v�=�*+m�q�Y�]�/<�5ύ�ܐ�T��,\�|}�wPF���Y৭T ���({ޒ'8�=�N+��S� �N�UQ�8O��0�I0d�6(��'Q9�>؈�r��<;�e��N��I��W=����/�r����Jn՞�&򓬘�����S��sbP����Stj��x����I������';#���!%��cτW��WvY�)WV����Gs�A �u�k�u5���T'����x��@��J ��Z91��F�&�jh�s]�Os���㕈�z���t(��R�(�]��s@��� ��[Bz`����\NU�m�ТA�q>+c��e"��~�� ����͓���Y^L�MVtَ�[f����}~L֩3q��T@'��u���vk��#�_ߝ:;}�3�ߩ-��RPS��Zǡߚ6�� =� �m��]ޫ)e�L1E�e�X�
ʤ�h/&�I�$�IF�J���T�%������$������f9H�<煹����G{1��c�C���U�n
���ɇ�3<�gg^BBO[��&��glg}���Ru�B�uiH=����r��ɤ��ڢA�� ���y'Y�K�����7�OX���%XN��@P}�TT�ri�V���U^$c�� ������{�^C�h�ŉ�4�r�%����y���3R*��gN�}hx|�`�<��Fg@�}�}ݕB"��P�b�rp�+���+5R╫Wh�`���c��u*$ܫ����q$�ݕB��Q���7�V���"E����J
z� �ʪ�B��F���i�q ��*�����$��vL9������'�d�	$os_:�z8�����m[��*Ǉ�ê����2��U3i�MB�ܲ�JT��FF�0[F�yw@��Ru�o���VJ߄�<�<�Y�y�=[.2L�ږ���;��ҹ�}Y�H*2$�u^�A�둰�鱁rq�'b
�Ś���ݧ�SԈ�����L����m4�u����#h�V�r�� �6��w�c�ޡ�=�W���
�i��	��M���r�� ��4r8ԍ��'ăojh�u�ew��.��b�}�_OU.6�nJ�*���Q�$�u�`�T�l
$?kTꀭ��`Vz��"E����O��	KۚKs ��ТI�w4'y��׏}B����}Lvv�c,v4HV� -�����q%���Xi�p�� 	�����
���rԿ^e�H?0�����ᛲ�F�e�Q�r��W�Y�ݝנ馷 /mA�o8ҭ������Ȼ:o2JG2h_�{�pB3�{��6�ҢK3�3,K�������V	H����.�r��56XC,qK��[g��n"�N��6���OJ���C�ܸ�z��bc��r%�Z���vv%��lU��
�IRS3���85�)�&F���\��\�rV��0���+q�3J��Nݧkн-��mQ���5re��h�ݷ��x;��M��|7S/a<iW��LpװzH�D����l�=�� ���_	��r�_��t ��:sF"1d(J`��j>b��k��D|{v�P#yĒ�u%���b�n��)B�Eߏv9�}�� �dC�����L݀P���(
�W1R�j�h)��μ#^�Y���9�Hb�h�I}�$�OvS{���_*�0]�T>�Oԅ����@��PLm��ܥ��+��W��ĂA'�*�o��K���Ϗϐ>�G��#�贄�fb���15�յjz�vB��b�@Q7���FfaI1(qS�4|�ĒH'����+�g�� P��@S�:��Ȋ����[�
���T��9w�P��$��������#"�@���R^V�=�w�����0��
P4�����b������Ӻ��%��I$��ʡ@���}�h�4�p
�Db$*6J���"���]�B� ��$��S]9�$k�O�� �eJ�)'�1*�~=���s.#�}F�8b( >�Ӫ�;ގ]�������8�N��6�QV�V��	��V4���	��� |y�P�I�렍�n4tmKc�	�E
��k�v�iH�=c�{gi�
�+.�T�{���u�D����*�ޘ�>�������#=��Z~T=��1�=�(�
4¿c`WH�8�q�D;7��I$��*�x�u�/O���g�i��/��)(tz�`��<�
Dʮ���uB�U����o*�v�i#yc��3�ħ��R���w8��f����Q�9B�$�;Ƣ���b׻�^��o2�\����|�I@����r�|(}����|��7O6�MMl����PX�b�'j�mc:k9%�I�۠��>ҁ��9Y��	�($ �6�ny���b����pm�1��#
��GM����������vH�y�4Gh�P��f��r�t�b��K�!uf�]IH�?I�پ
f�+!��y�T	$j愙6�A�n���%�Ɖ��0���x{J
���0��wA$���{�5$�T�X9�_]ZRG�� �/�{9���Q����OvP���F�L�V�D�Й�{����FQ����!AY�7�G[�nh79�-��Z�Ci: ��w���$�d��w��Ǝ�YZ��)˧x��� �_mMPx����V�H��F��Y'�u�\��(�\M4�U�E]�X�7��d%�L�&�y�����p���~��:�sr��ݕTzog!,�AH��MU.eP����Tm*J�a{����N�{-��xy�I$Zz��A�ʑF:��x����m/TF�͔�q�| �L��ض'^���H����OvUQ�>Ɖ��J�P�a��1����S6j|H$m��G��\	�B[�Q��(Ή,U����3V�r(�u]j�C�!K�EUD�I=yT+�n�U��o�u���Yl�W��x�ɽΏ�������M+��"�X�(�'�њn�L�]��Zz���� �U����8���{��05e��v��yS�����K��naN�v�Y.���^==��h���5���2�]1�LT�Дu�(sdҳQ���A���_���^�A�y��{��j8���Og�]�/.X�����l�k	�=74cv��Z�k��]�nӵ�z����X�kiiM�yz����S���2t	Iw] �G�0���p}��|�2 ��!���|I�ڡ@�������v�J��h};�q���`�7�Ң�Qc��Xc���I��D����^Vz}������5ݫB�*W`��E��=�� A�=Hnݳ�!�Gf�z�'�{*����*�0.��Gu���o�oQ%kuD�GsʠH$�t^LuA��tⲮk`�T�AAZ�B�������@3��@}�����@��`�J��J[��	�J�Q܎�Zsq�&�!f���� �P��~w���7���f�.ohQ ��D�H=�qFU�f	�]?�����c ��U�	����
gQ^�=<K����],��n�{,�=|�͙�B��W���]�ٹ�l�l����~EA������9Y�I���T	#��A�M�s��7CB�F&V7��	f�I���]g��G�>�����t�)��dD�Tg�"9*�p��jEΉ$���j˴#���	���pB�fE�3�I>=yu�槏n����EA��	 �eЬT�;U<�$` ʛ�		 .��;�����@� �v��g�o{��g�3�	vtO�'z�hS\MS����� ��؞ �}tR��m���h�s�:O�z�@$�{�*�2���r �'���+�>
�Z����� ?>t��S�OV~|�y;?��������8;�,fa�+^t�԰�vuc�uZg�n�wv�WXJ����tJ�|2F���r�9�sE�)��|�6q�z��@8�Q��:����m�H(���z@�ܺ��史\y�k�*t�뚬u�r{N4����op�5j����a���Բ�������V��~cf�ƨ���0/4c3(SJ�LW��R�:p��V!a��4�]j�]dj�r�Ɩ��E���%�ymc�x��͡������(w[�U�8���Y����A����;��򙖙�Rڠ�x�8�ggu���n
+A��r��y���f蔛������WυA�n�uha����]�Zзu����|rd�Gr���5��˃W�>��.�v>7v$������
t̬����VK/�Y�-u��pÙ�m"�ވ��η1�t"v�NeS*U&�����J�@
�4��zk/����$��-�;��z�v'^7��3�AV�vޭ����>٘C,&nƕ�]F����ۆ�	v���C kr� u�������b�y�̶�I�:﬛���]]rfg-$�+ ��kpPs�u>ѐ��novgu�V�Vf%����Gw��\V�
'#��^���AU�3ke�53�K�h���?UBȠI��'��s�Nz�p.�.\.P$�C�Y9��N{�{�=z�"��e�1L�RN\��T�=*.�s��fT��Ӕ�����ad%Vv.�u�G�g�c�kBH�8��e�Փ��Nm�E�@z�W%�z�ەP�����+��H5�SiP�5���H��/$��9P"�{�Nw!�BBr"� �g8\)�.�;�ϐʼ�g������Ƞ�չ�p�����zǝ���ry�T��z�U<�C)�w!�''"t��@V�E"���<�9�ǽ�������<Ƞ)�SPre�v��s0�;r������1��������|q��h���GR�W~=����o�yGϜ	$�{YB��w�F�r�4�^�7�j�)Y��݂�/Nt�	�i�8NyvS���
ǍР7�m�9����L��AR@]�(W5�����[p��F��J�m��.�;]���#~eS[��>���C��` +��ص��z���]!S������
�P"�
���Af�����I>7��@�w�����Y�գ�.�Ȣ]h�$O�)��ۺ	�uB�%��O�`���}��,�g"��"`�Q��{��t���)}GĜͩ�	�Ӝ��#�U���I��A��r�5�~1}���Ӣ�˽�ipej�t���6�_�+ �a�
�Uf��!^o]�0�GsVB7W�_}��Q#�$,���i����TI"��Q$��ReS�\�üF�� �f L�,c\ܾ�[�I(��5����\��~����l��Z}V�7@fz?��(p�B�bpG��� +{���R�X�B��)��b���1�Fp޶(�O���j�R	h���l�k��R�f"AF=�Di�RH$Ⱥ����y��	'��uD�O�g���/��RG�;g`ꞓ�|!�W��KXԒ	=�B�����$�����V+>b�XO�"��?s[�bh��*d<�?5�Cx� �o�i�!�Q��ǎU��J�	)��U�r��[��&�D���y	�MF��C�<:m�X�P����.b*�'���������+a6���qC�8��p��m����)8�חb&�8��69��\�2l\�Z���u%Ȯ�@�����g����\KE��6l������4����4��ؐ����Ю5<�:y6���q�\���#w���gR��&�Vh���:�Snsꭷ(��$�e�"Ts�;f�P�-K����꽧��!���+������ �J*�w��IÜ��|OvUP;��c�ht�K�l�)'�����H��n��bt6o���ul�8_y�	%�jA>$��UI��nhEwe0M�,A�&J3"�J�BA�U�$���e�M+�` C�4���柪���Յv�a�+�z���ע��RRZ4��c���ek؞�������H&��z}Lݞ�t(�A�y@Sp黳:g1]��WJI$�u^��ݔ)��7�:z��SM��y4�X.��ͧ����ɕkGM�	�i��m���<l��lswݞ�i�:��� >��7C�����t�y��S^C�R�b`����B�5|��'03,˴
�Z�cޙ>ߧ��9����@�a@r7�__!�۽�H����l�Y�T�TD�{���$�mР{�ɯ�K��E)�%�����H��n����
��&ee�Ej����(S�: W{���B��,�)2.�QU�l5�n��|	�*�$�t��5��3��TF��0D-r0�Ή/������>�۪ �nUH���b�𣄂�PR�%0�^{A����L��tۮ;NCYr�.u�q�~��Ϲ��n�����1��L
���].�ߢ�]�rf���"�3sg�A0gJ�$�ݏb�J��9w<H%�ʠI#Vr�LΑ]y��f]�W�B�LLv��T8u�$��m�{���&U.J�Ӷ���˷���rݽN�NJ�����kǃ��r��[��n��V-��h5y^X�y4�No�{Օ]�$��^'埊�+V�a�.Ű��s'n�&�K�<0 ������P |:zd"�]O��?(����؁e"R��4�̍ҚJ�* +�z� ��UP�:z:zO��ߺ��>gs�}�Z���+2�j��ӭ�\�7]WSŇ�\�k�}?w=���o�=���ў(
:z6&I�yt��O�q}��y	V�,I"D�آkn��(���=D��r�H$��P��3�+,0�A�DL��9I}uD6�.v;���I>�P�H=}sr0*jB�LLOǻV	��מ%B�&�\׈>}�O#UV�y�L��'&�Kp3��w�*��{�}��q�^����%�4f��pM�T���¾&^U�B�H��/��LPg�oۇ5������j�A���vMx������ϵ��/�Kl�Wh���q�����O�����]��v���_����Ϧ<���.h�O�������*��F�H����_�e�(Z�E��W�l���KU�rdH���>'�z�Q{����W!X�_Z�j�X�D�U`�T	/r��wmw_��A�*�*�=�R*��=f�Z��xߍ{.��Q�1r`U;���#Vr��U�8�H5�Ө`W�B�LLCz�AíH,^M�rN�:����T ��&�5>�:}}<�b;x�$njmj�9�,D��{6����D�q$�U��s1��M]��0%{L�m�G�<p��븛*��U�)uV��\ԏ��v�v�k�\�^6�ٳL����p��V^�X��/�����]���^-��C��q�D󫃞y�\�i�m�Ͱ�F@g�#l���������n��3�̲麳��t�YR�9��w�`֎�$6�W6�4������1�F7�/k�e٪�\⛷.l���3�H�6����k3�a�b룦��=���g�g��	��D	圆���az���3����E��J�G�UA�C]l���95:I7����! �j���u��*���YM��@�P�A㜤B��}�Ș)^0I!��Q��*mP�D�U���h9�B��=s�(�8�BA ��DG<�N؟�΅X�r �!�3�j�A=��P����ֺ`x� (t~le0�u� O��tZ�;�S]���V��:��K[-���wF��Lb`��w�ТFjI$���E������v[JߐX�Ɋ�Z��2Ĥfۼ���2�DGGl���3:�b����~@�(U��o��O���9a�o%���wy�ӫm�U�ui�ʩ�u����X�G���BA'믨P e�3	wV�x��]r��%2�H���� ���$�u�Oc�߈<�)�u�+D�P�D���c�U�:�N	$9�H ��P�_vJ��EܰN*�$��C�$�"U٩ͪ�cx�F�g�4�W�H'��P'��h^�av�y���h�a��p7*��/$򹱶������7s����R;]�����A}9B�$���Fu�*��k��6>�������eX�>���|���ý��b�H'׳�^$�v�UL�Kѽi�/����~]�E$@V-����7��^$ϗT'�4.t��g�{�ו�N�Z��3��6�G�k2@�K��b��j�*��9���Y���*�y$�뺋��s���b͝���ۺ�.�r�����ː�i}�	��Q�$��T�q�m���Ͻ��O�2�����y^��OjJ裓f,�H�Ϊ�{��$��Rmȵ4��5?��/FB�a�`Y�e����u��D-)u�5�4�~��Oa>	�*�5��P=��{T��)��)A�}B�Fg]�T���"&L��҄�۹��p�t�n��>�#Oj��힪���;#�@�L3c��Yy�H5[Q[4n��w�	8��'ƶ�V��^N���*>�+q7TA�r�|O�M��w]np�#
bN�`�׍�W��5ޣk�������'i�2��\�nM�Ӗ�ˢ�v��ѝ�+�:��B�I������}�oﾪ'�G� ��H�U">�(5?%s0�z�=�>k�龡[�";�8�z&��#�.uKQ̉��G��.����0u�X��v�����vLIHHI��uD�9�A$���-|�ڞhƺ�
þ(��$JT�D����nbc��-L�1GĒ�5$��
�q"��0v��7�dѺ�i��� 牊<ϵ����T�*��u�A-f�z몈�20a�����u�5<���"�>3�L�I&�mz�vP�~�8���=Q�I8NՄBHv-���
��t���9���w���sgĒoi�	��񑣎1Wv��{�z�ύ�GLT>�Y�)��6��o^p۽�������	R<����lɃ��]����d��͸xT9�e�YǪ�"�t�F��(�0����ɒ�S,6'7]FỘ�&�P���!���P� �[ĖݦX|�4�FR���J������֥HV�A�̧D�k���;/j8�*(g-Q��r�nBA�7�D�=���e�ê\�*U���p[ǕgXs	6s�Q$g1�r��,��d!ĺl�d�O�pQ�
p51m�9�j���`}���xa��1�;ձ�D4~��iM�\k
6�a����������(���y{9
��)S�������\ϵ�acy�:k��W=:����<U�#ӽ��9�X�pz�Ŋ�����*���ͨ�8_:����WE0i�;�D�J�������Z�ԛh��gk���j���]t��3s61��vȅ��s���3/;�ŝ������5��½c��ޓ,tЊm)�NqK��c�Ձ���ੜ�*n��o9n�;_�:����q�(� 8
5�m��JA�����M*�]��h�uٔU�0�ȊӮ����C�`�v/�y&�H7����Nv��vV���2Tf􋭄2�/7F1�Yd9�>����K���a�Rfr9IY�A$��܊��<�wgq��d5�"�;�o�"�9��M��y�G+����w`����(�ʂ�C�̋�����71P/$�4r�z+��M��bBCr!��s�5G''CiǺ�T�N޻�T^���Nw��r�xM/����`]4����\4@�zvUܓ�ӱ�$9�$�*���A�s�<�np�t�T��R�i�������R��@]8�ȼ� #�F�rJ�C�{�&��^��/=r';ϳ�7\�E�H���Ν����pNʲ�|�А�kcyC��u���@6�L�9��9�s�ݎ̩�\��ie�t��١�k�R�cL�,�e����^�^cth6N=�Cicg�.��=���1���L�z�������3���2�u!(M��ǧ<�ۜ�Pg�&0*�lMa(�,c+R-��f3� \�X�;c1���/h�j��b��j���7@�ل��ke$���-��x�`��h��$g�Y�l$[�+Ю%;�=	����f[%v��q)3E�����|a;]7fp0rB�R{&Z�|�e���헮��H��f7,�/^M�!ͻ�Q�sf���B��b����]��Q�b��;6y��v8'>�m
�\�8�*�9M�X)nY`l�M�[�A���h�d�� -��c3���j3[<�cF�_燐��Ll�c�V��yY9:��p�>v���3�hM�k�G5�4A�4*��	i+��-�>H���_㏎#���l���v���s�$Io6@��ѓ�ËY��I�]ZU��picw0d�s40�	G�����I���]\�M�5�X �-�5v�v��٭:�vṫ�ccK6V�4ɩA,�.<B7n[tz*q��\g���%S���B틨�Δ�.w<x�7`"�^��#��<�-ýmƐ�{Q���r�&��4i1����`l@���^�#�TWH;�]v�\���˹ůn�/:v���[�w�Z엙�Xv���ŨY�ۉ`]�[,\ݥе��4�X�)��l���A-\rP=Fԭ�n��u={!�Vm[���%�N̻���[�k5���z�l��>_Q�2M�/k��Ǟ
�y�y�Qӭ 6;M-s�	��������j��$�ZӢ]yPv�<�mT��]�Y�%��5����`��3���29Yl;�X�RPWaΜnxl�c��"�.�@��1�{NC
��t4Kt#e���K��[�քR�X��Æ�m&K��ݶіv�]I�d�Z��l�Q��ð]�q�'��N�絁X-ۉ���Y�AyGi��(�6�f�K*箠�rv�CJ��,>v;���DE��b������]�E���Kׂ�~t�C�ؘ���&�f�n(	�����(��*��剄���0��`P������{[�J�{��
du�*��Q��.�r�������l|H�-3b�>O�:�os� ��YK! �A��5�㯔���x�j]Mx�y�TH$s�$��V�מ!v�Q�2p0��DE�=|��@$�dؓ�M���	UfU	��=���92�'VMp�F��i Ǡ/I�.����n���/2,K��m���>��,T���	��L|�~2ݷr�"��΀��S�>�/^�6��RR�_/�]�U�}����7ӐKs@ǡ�ō���X�̡�(s��NX2N��p�:�#����R��#�Q�aN��P�׏�r�g������	�� ����(Y��p��rI��x�E/�T��@�K�'ǳ�	i�I��[�q4O�|�'ݝ"A4+��I)�Wf+��ԍ�M�k'��z�I$����+	���0��&Lӎ�'��\�+�j�)�t�'���H5�ҭ�(��������`���0�]YS����4^^�p\���Һ$�Q%���#��eLB�޺�g8I t~lY
̫����({=t�Հy�$��X�l{���qD6�~��Q)� w:D�Iۮ�^5=Rz���)����go"�6��R|� 8��C޻��u���T����a���`,\g7�8�J��,�22DDK[�'"K:U
[p��Q6�C�����sZI#wʕ@P��m/6Q�(D�/,���ٸ�W���1�$�WMx�;�*�2�ɗC��H�x�����dg�@�����n	h�vL��$v�РA#w��w3�-�m@���0e@�s�&("�U��[�M6�M�s����D�v����$�VU|H}�TF;�y^t̉'���㬣��B�	Y2����L׈���Ely�I몼I=��(bxָ�W�sPv�)*Y�C{1��|'���eDۨ���4�P$�vP����H��-T�/b��Ϙ�.��nJ{ۊ�'�H��j˄j�hm4/��@˥��9Y�_gWW��C7�WY2�)D��[�\��jh���j8:eۚ��xy�I�͠(蝪R�H*BBM��A�@�A�j9Fwc��|��Q ��}A��k��:���'(ٞ��<]��^vq�/;]8�!03Yp��m4\w�����aD�J�5/j���@Q$��n�z_=�U˪Č�ʠH��,�!12f�G��?;�Q[���Q� �c�;}t�W�`*�v;|Ҍc�#�a	�z�ТO�s� �Ng]lwT;[y4��J�Հs�Q��XF��ݙ9�·��e
���g�H=u��׼o�o���o�3y�*D*6��R/b� ~t���;6MFK"A"&j��ہ$z몹�H����U��)�����ö���bg+�Lʊ�ЀI[s�7k���l;�%ӗV���j[o���L�rI������5��Q)]��],�㺼b�n6}K*0��ȸuđ�VH޷�bƱ�P�I�V�,It����Պ�l�y�hd+��b&6��j��6���[�`�pT��c�곶 ��s'a���rn:7]mO��ue��.���M���Qk����j]J����%�:�f&ՌNY�n�!�h�Ѥf0��f��M6��/�u�`Mc��V���$H'����k�w>n����7��UO���h��6*���j��{c�{��
��t(w\V\XuU<�K���#&L�\p�;k*���
{��Hy�$A뮡D]Go��2R��� J"`��̀H$����F�eЫ��y�".�L����cH���XF�vb`	��(��XDI�O�:�	>��T�h2�ύ}]�8����g�5A�)EΫlH��v6B)_������10bC�K�2Iu�(�I�oezQ6委Vn��e�R N|��<�������U��!r��0�R�pr:3M]:dK���>~>=l�[��ܫ��r�t�R�iض1�[���6�Qѯ�@�\�����s�67��X�i��o��̷�����
&"U	��������+������NE��C	�1���,ZA{� gQ܃2�P���	#{���Oa�w7�0U�
>�ma�|��2�z����\�N��5����/^��A��\�<��.|}�ջ�/[jGm��ֶ6���Y��A�-�fcccL1�mI ��=䊻J��7�����=�����Hia��p�<盠O{�*y/]�J�
�� #��T�Y��$�z�X��dH$�9��ko�9����=51 ��Fvu߬�K�O���b���Ub�6 C� ������M��F���3Y�^�2ҧm����aT�N����D��'1�$�C(N�Ъ�		N^��66w���e7��َ��J�h�W���D殊|J�=% >����E�.�Y�wT�?L�("�n]݂lZA:�%K�@{�+�����OE�ذH��H ��W�Z���'m�������/R��k���F�cU4�5�5b祭�"�X:ʎ�1"J[���;|Db�$�v窏dG(��%��Uw�_&Hx�E]�Vi�t���/p��C�˓)� ^�� ���@w�~Ujp4��Cs=�!@��(�*v=��z�@�W8̽qG���V�I۞�!���QIP!	4��؋���h�6�$=s�D���A���R�nb����v	(�7/q��L�(DI��B%X$��������k�ͷs�U�Km�|�!-�6�;��~x�n��uW1�� =��g�u��HzǮd���P��P ���v�{R�E=�v\��Ic�db�7��v��i�4cu��+4曙��7]�|��Z��21�q>$ӕ��΅C�q'��-^@���1����BT�2��c�o�z�f��v��I �y.��s�!�ݡ}����Iȩ�0!	Q@�̚$�>v,�I�2J��5ʧ�	�'b�t �{� K�7J�
�()��Ȼ��'Uݻĝ���I��w`�N�ިl�C��Ԏ5whwVi�k�:\
���]N�r���O�7T	$v�l�@|<�УCG��w��q�7�;�����<K����K�(�W��X�@�>���}'��z��9�q��{i����9�����MM�.[5f��V����N�۴��W�����Uς�;�p�����\�&u�vq�kh��ԭ�Ƙ�Y��&����ٙi����4�.V��CJ:jMQT��4ܝvl��Q�&��f�C����4P3����6#����m�͵�<�ghA��E��6s�u��'KkFng��{A�Z�Z1Ƞ;q�r`6�i������\�%\u�K��t�g�d�P��C�:7��~�>y�^>��v,4Ao""
Pbd�����/-B�Pr�� g��
 ym�F�)���]�6efD���=}N��1u���V+�w9���0��|	������@m�m#v���7^�5�Ofq�`�^U����OOD�N�Ve8޸*s�B�K;ҧ%�p��vQT�OZ�
�*�뇛��B�+���I��eNb��k����tA���B0�D;sf`�h݉�lu�Y�v��g�߾}�ūk�<�~��GK�$�{��<g�r9�"f�/�\�������h]� ~z�]BWv��7���.\�ؽ����~�w��[�<�n9zB
�%��I�\A��1�	��7S��)���w��S��d�As� �O}�B�[��	gN:�;��Ӿ�`5��%���l���H�pv�ۆz�X�#v='�*hd��5%D%H ���zc���u��u��EvUQ$�we�]�ӯ/#b��x]�.�՚F�~���*g��aʻj�R����A��T	>}�w`����������mY�:T�v�WPw3���L�Z",s�)=�7�]+��*��?Z� � ��݂j�Ee0=� �/���b�b"Q1�!w:d�3x�}5�$������B�>2w
���'8鵆b@�J�-��N�۰,���w������+C���:�� (����2�N�E��X����-��y0��k	w.�KT��5{#{�\Hm���[Yvf�$/��捰h�ݭMi�"o�4��5[�SwL<-m<����l]��+Sy7!�Ke���W]�m�� ���y�X�\9����W������gP����K�����\W�^}s�+�SK���8�)��v���R���a�����@N-�b��o�1%s��T&��H�[M�U�+LӔI��-�-����[mڗ�{6����3b������mA�ݥ�O�*Uҫoc}MAHEGwzK�H� �	�o���9X�Q���%�G*V��l�L�О@&J��/���5de`S�R��4�����R�+�Aw��u�]��N�����I��K�E
B�]N�rﺹO��eNৰvK �cG/��n'gl�˦�4Ү븭q�������:�q{�"6�̌�0S�v�=�^�G�U���ך�	5�F;[���D�1Ϲ����T��{}�^;����3�̚�,�ѧ)�p����Y���]�&�ٰ=u�N���7�l�j�2�-���+�Z���sA�5�y�30:����G����##�#
a)�܃E�������i���&M;)"�u�ykA:��@�rY��ds��@�q���t�<޴�99�+�
�ry�*�^r�8$��d����=�OK��k��ʹn�tt�r�G��!���#Ƿv�Uw=��I3�{�<����GO��=z�!���a�i7*f<݋�&EMɉ�Gp.Y��;z!�^�eBr��m!#W� �'���v�rF��x�"�Ws�����͔<��wS��^Nxq9c��m5���#��r��'���:���{޹$��<����tˎ������|��	A��s֌y6�P�s̮�=`G(�r5���!���e˱�+ǽ�G���ޤ�dU�|��xf@G���D[���w$ �צ�Es�X���Ԓ� I>�����g�|�þ�q��;珞Ab#�ӿ��Ϯ�~���m�˪$�Ϯ��#�gZ�A�c�PF�8Ù�)�%+���ݒA�U`��c6,q�e�	��wd�s�*5�Ϭ%�ѳ�MBh�D1�	d��H�6��a^�a[��� ۾B�]Y�o�C���	��pH1��FE����WnO�_=���z�t�ՒUI���
O�w%AJkzw��Ն�z�{�dA�iD�~��KF���}�K�������4ً�nU�GTT/1�m\�0��H" w�]�᠌�3ֵ~+���U�z�b^iF�5�{XF�i�0�Q�h��]�`h�>{o[�TH:��F���3>�/��Ϯ�փ-.�F�j4k�0��4����R��[A�8�6{�݁������J\љ)O���v�4#��Xw"d=\ة3�Ӹml����ۆ��7�7���<��;
#2'+F�<	��;��#L�mw|�uEJ�v����qv�Q�l ��c�db�A�����g}�q�M�o�r�1�C҉��۶�Q�l��{�e3-5�ży?�w(݅ ��ʉ�AQ�@B�FFl�5����f!D�
$��R�#������aL._?���pL��	}N�E� G�}�Iz���7�Α�!��aE�=t�6�s��L۪����ز0��u���J5O��������V�'����֘��F�]�)��q��1$=�n��`��AgO]����A���#�Cf�ج�캫�%�,���g�M`iF!���7fX��6�4F�V�U^��}R�FX��1�]{�LCia�������Fe��Ϯ]�S�*��eƌ_��'���^��#�� �殞��Cd`F@߱��e�������4÷Zў�����b��6�0��U��1���zܺ�Aʷ�i�C����0���iA���s���֘�ǽ�M�6SI������4h#�D$=�z��`��h#�=�{XF�� ��kx�G��^N)����6)��q��&-�д�GjV[�
�D{S�s:�:�/�ǘMJ�]�4���n�zy��jyhC�k��Rk56�nm�wb�g�����:3�C)�׍��Q��
�{��%*q۬�bj.^'G8ݔE��f���BF�4�V��+���Q���}����V�nw1�e�Tk�d{:q�:ɇ�i��]#���klyvy��1�G��1!6��6.��3���3=�d�ֶ�F�V��&�[��@�q�����"�m��oY珱b#��g�]�b�4��F(�k�0�)�4F��w��Q�-0�Z�}�j�G=z�/��B4��V3t���iA��6g��,�A���wjU���X���o�q鈄�.��kĽm��	/�O)��Cb5�r��2��F�j3����i��(�Q���㳛��w��=wLCh��=R�U\�XE�ta��a��j4�j4k~��i5�!���w�����Y��i�Ӎq����`a�lCys��0�3L�{�ՕU]I,�h31ۦ�;�wT��ZKlCai�3����Ŗb��4Nw��Q�-#�Q2�ܺiLg>�^2����`D���ٰ0�h��\��%QR�A�1~�0zb"�D$Asܺx�ɛ�}R������s�2�6�4�Q��=�#LCa�(�4]{�M#E��N���R�t��N1�/c�֯m���U�Gn8��q�:ݖU\ן��%�U��,^Fg�S��Q���;�kL�����w�6�է�tы��;��C��,�n4�߽�#L�������VJ*T���0̴�������j4�_�랲���w[oz�gu�?5�-��S�حVb�E��L�F���*9OK�p�7��]β�ޡ��S��]�F�̬�1X��&6�|G���Dh��{̣LCb�҉��۶!���`{��������k�q�h&�>�ݩWl�:h4�G������6"H���v�4�l��{&L���]�c�ֺ����(��w��2�LQ�LQ��~���'8NԬN�e�l[a��v���r�bJ��Ec^�&���������'��I��=��3�]��|�Ƃ4s�װ��L��>gVTuUu$� i�M)���&�j&�a�3�f̦,��j�rz�B���F��c[�4Ŧ�m(ˮr饆���{V,��@��{����{2�n��YWj��.�el�8m+5�M�����ڋ���p��y������߽�e�Ԃ"��r��4�h# 0#!�{8,�5�z�ɛ���*k���aa��1�h��.�0�#D3���r�9*�Q�-#3�r����O��{�uB5������t�@��Ch%�9�h0�؉!�{Vs7�o��2�s�1�o�40#'4��U�ʕ*��4�ۦ�ҍA�A�3�ެ1�m�^^��
��a]u̲?3��A"��ڒۈ��ZV��)�7yWu7���u����㎳���k5�W�i���F��}t��Q��Cgu�X�̴�ɾ[�R��Sh4�G����c/þe��Ch9=��!�4�`FC��X��F�j3����i�5�]��b��Fh�{�M#D/�'jVJ�t2�(�,�#;�n�,2�6��߽�kL
ս�N�g��d�o�!�C�D	�z�0�6!��;�{�F����sT����e�3s�QI����#k��ּ�j�
M��Z n�56�ߞ�]R����?�KU�]5��j(�Q�׵fX��Q�m{��2�1�$����U���m-��owLCia�������S2�C��uu-ܕEKym\h����i鈒�ϸ�U���&�t�7Ƃ1��ްY�j(�L�}��b&(�2����#:�n�8�!��;�)�9V�1hFg�偆�Z�(�h�����Zb�y�o���ý�z�8�A�"Hg[Ձ��؆�Þ���i��ޟ9R�Yr�]<��e4�W릫F�{��kJ0�e�)�,#h��ﻼ�LZa�҃.�릗)���u�N�a�3�cT_����h;���7癝.[.��&��lż9=����V+]
L=��u�M.�����0�g�=&�U���.gM�h���`4��6!�;˧��=W6�\�xfOg�)��w�XfX�m罼#,41F�0�[��FDh�y��bYk����wnV�9�<gs�ݶ먇<E솄�8ql�1uE���������ؼ0��}�,��JF�o��i�����~�1��W��s�Ϊ��划�v���؆��{緄i�l��?j��Uc� i�ij���!��;��#��o�2{]�@Ŗ!�F������2š�bAs~�ia�ҍFo��g�'c��^�M{�ԷrJu-�q��s��!����]<4���Cc�a��~��9[���D4�Q��=�#LCa�(�\߮��џnY�EF9V���m0�ϳ��bG��y̷��K��ҍF��=�i�dh"��LCh0�b;����w��s��pCb�o^��!�[ק*�6�˕t����[iF�J1��u`a�ݾs��OW=ǝ�(h��o��4š�b�#J%��m,5Pj0 ��{z����*w�򩿏ʣ�#h�p"�(t�/9E��[�MbJ��M�7km[�XE���.��<���jd������Ƽ�<�ߩ��e]
�@HQAQ �|m�[�%���D�ڗ�����(t�\V��qE�6z�=���G�q���9۳&�>�jI9�
�f�`�'3���wu)ƻ����]+m�2��!q4l�O.x]���;P�;�J��$a��&�7Gl<��u��ص�$#�"M�\����<��\qW[�n6ڃ��g����F�:����.��jh꺢i�Dۯ'��Ы�u����7�e�� �H�߹v�4Ƃ1�﷬�e0#U�o\��KM��8FXt�1F��}vц���	ꕒ��w�[��wVL2ҍF�Lw��z�s�k�M8�0���m�󘶃4q�l���9��}8!���@y������w#UJ��0Z�f�(�iF!�>ެ1� �=��7oﳬj�ޣ�됓B�%���L.���﷫Fe���ߵutY%UKymAƌ_��ew�z��Cb:H��ػx�Ad;�� e�me�����aþ�y~��\a�(�&����	�4Moq��]'*�Q�-0��s��iF�JF�{����^���w�<�6�KǱlCb�sڰ2�7�{���!��Z�0?����O7���`_W)]p�h�[`��(�tn. z�E����-�%�rr��ùr����<�S�۶�ҍDҌ#g5�XbFZ#G;�o�ط��8sX�oA����붖�(5��wz�dfZ���$�l��Z8��s<�hzb�������j�[����#4��K�@�ņd5ߜ޾Z�Zj��1��!��[��vT��US�d���d��^���{�[��GȘ��5`a��&�j�}��bQ�&Lw-�;��"���#D�l��Y(��yE�da��ve��(�h����`hd`A���u�{����A�Ƃ1C>����9�{xFY���{SN��QvݙL����Xj�u���V��TҌ ����0�� �&��k(���m(3x�a�R���������Q��s����,������.4b��ab5 ��^�V��GY�}�sU^����I�������iF�s�����F�߫j���~Rn)��M��Vu�h�B�����2��:�`�AnL��9ؗ&k������}�NQ�������3a�iA�҃Q���u�e�lCh+~�b@�3~׷:�3ٛ��G�U{�0��g[�p�X���n�QQʧ�Z�P[B6s>Ϯ�s\������0�h��4s��i�bA{�[KF!�5���q�l��V-�A=�r{������t�iƏ{y�C�LTb+��N��	! ����L�a*���}��l��2�1=�/9��5�ۗT�t£ⶕgS�U��H-�δ%���SWD's�q�`F�4�G��o�	�0�Q�h��]�`#D9��+4����-�,#=����}6;�=4bJƣF�y�&����24�붃4q�����X���p�؆��G�u�#L�����q�R��QV;2����uv��jJ1���`a�;[��^{��qd�рh��5�eb��1A�h��m,5Q5����b�fZ��sO��-��,��;��{�;�X�b����^�f�\ԕ��i���w�站�-]lCh��9�e�lG�;߮؆�6a�=�� e�mo�����=�6����޳�#L4���&�~��F��3���5t8��yF���{�0���in�����F=�w��#���b؆�a�"H{�Ձ�0Cq4j�Y���c%׆��H��Zb.I�
.�@�24���m`iF�J0�g�ܑ`�Y�/|:c����L�i䷾��Za�҉��˶���dg��X�3-�I�:�%�Uy�A�=��ꘞ���#Ă$������1�0#5������ҍ������5��&*e�p��v2J����H��}�X'�P�ϴ�u�/(���m]7VN��^�k�r�Oe����q���A�kܻh��'1���L��p��0Őa��vL2҃Q��߽�kLw��y�:α��F��uv�aƂ8�I{��0�7g�"���:��0 Duv'�^�u��;W�x��,Imb��bNGM��\X��Gk��߼:�Uc��m�y�n��ҍF�a�3��l�b�����{��2Ť�D{u���tE�\Y�|�{���'ޠTb23��lY����{�tY%U]m\h����2�h$�2�oRzm�]���G�2Ȼ�� e�`F�J5����4�6LQ�f���8G��ǳ'��>����%xʷ�i�L#=�����Y��;��21�����V<�xմq�lD����&`��6�{���i�뼢�6:u*��3#Jn�vֲV;
�;���J0�Q��ṉe�lCh��{̣LCbKI��붖wZ�&���=:�:�KmF!��^�0�d�M�ͺ�.���:h44w��0��m����h#����1��ޠ�6����5�2̦bG����Q�l#D���	�4u+�u����;�W���X_t�9����>�t�ݺ.��Ύ����B�a�P�P������l�b���5[W�k�}-^��v��O^�Q�.q9	��k)�ѹ�m,���g�l��n�n?.&��gR,�%�E��lw�X�]u+ٵ��<�2dt��Kn��Z�ҭ� �ٖ�$X{q-�S� 9� d������9����D�:α\��&�8,�����ˏl��	{�ekŵG�DN�F%��/QS���¢�F�dp���m;�.ڗӀ��s�H����j���]��Z���A�w#�͠m� ��j̭�wF�rwٔ-�8/D7kw!0èWBfZ|�nej����ݨسPYp�Ō�{;��̀�3�E��ܩ�c�f@1�{J=�5�-d�`��İ+J2scFK��j��B�i�-c)�W/�Jغ�;{Xv��@�1��[b�^m���RAW݇hgq�;�@&���]\Z���G|n�������|������]Y�u1�<�(0�!��Q��3x��t�L��WyЛ�N�\pܻщ=���2o<�q�ٮ游�ƴِ��'�@V�!��{�˻��-|V���&c7X����A�R���Ȍb;ܙ`J��Vj�;d˿��g	��0�>�����=-X�{������)?Gp�

.�{�����eĮ���g���e�=���ޯ;��aBr�򤪃ޏtr��9ە7 �eЋ�Hs���u�
4z{����I�9۫]�wX�
T.˧���<��<�YBq"�R�>�D��<�{ǽ�E���rri�M���wE�g
h�.��f�NWs���L��)�E�Y$\N��T�%EP�T�^I�p��P\��7K"�tɖ����r���RI�S*�dz�ʹw]�t�Sn�o7*i�G2�{�Ay�4���(��y�ziS�'b��*�yܜ�r��L��()�ʵ
���b�\�O*���r�;�r�����WD�XDDTE��*����r��r(���Ĉ������TDh�I
��""���;��NVt���Q(�P�U��S�|�����qc�KҷW����L�'i�^��k��JՋ[�z��^��)������9K*l�9 �;��[��r;;G]ֶ׆c[�����p�
<��絻������]�f�t�zM��5ص��]3]�u[G���B�`zx���v�ۘ�$t]�̒	���X4-����v��s�&D�ꃢxyN�=����ڥ��t�*ڭ^u�;��-^��E�7d���JA�-��WV[3a7v�O3ɹ���n淉�n��c�8̳B�	`��/�v,�b;�a�%j@f�@u6��bָ�m!m�ݱtuk�qؘWh��hY�(����$Ye��v5��v#���J�t\��Z���OgX���|ؕ��P-6,]s�@����(��k��p8�,�7]Bd��G+붳�7nm��*����뉮Gr��Rf�#�ф	�sWA���9��l�cs�e�R��l�Ö�>���Z���!�t벝�tN�۬q]������T�6���F����6oG'��u��^z<p��U�N5읝<�r��v8����X�۔�Q�BΔ6��v���K��&���\���fR��n5v����H�3���E�Lx5�ܲ�cc7[n �.�w]���]8L[KgJp+��cD�qS�5�MP�э��em�	�Mq����@�e��1������v�\����ڋ��D��:G�n���ƹ2��th��d	���\y�|9x�s%�Lj8��}�����Wm�n�Etf�su�W��jY�r:麇�s�Ki^Y�,ӭBhf���+ѣ�a5�����l�s�5s�q��C�u�uD�@W;c56�])���d��.ܦ��YΑ��3�p��C˸�u̝����'��u�r��+̯]��B:U��Gч4�6�lvfݷ7
׻>�qs<'��A l��LpA��;i�l�J�a��M���`�Cݮ\Xg6�̬�Oi�P�%�k�������C����Wb��Pp���,$]]j�DtK�Ypѹ���J���Y�mB�3v��sc�J���w�F���5`a��MF!�k~�0hkL����%�ض����M�}�S�oY�2fn4��;�#L�3�;��UR���,�Қ���J5Q���t|�y]��g�0��Q����y�e�C��;�.�Xj4��`t��\}t�d\=��Y�t�����"&̶�#��;�#,F�I;�.��8�FA��ֵ3�:���b[Q�׹�aa�b� �~��F�ў�=����%��2Ŧ�ƹa���S]��-��J5=�kX4��@����_y0�>1Q�׳`s8�3�gb�A+��0��C2.f�\wWc�R��@�24�����ҍA����ٳ,Y`���n�zo��M�#D߹�eb���%�m,F�MFF{^͋,�A����?������H���`�%�*3hA�f�f�!�"�aD�2�+F�1*I<π���״!�&*1V�?���S
| Ig�@#��e��{j����y��N�-����@�ܻh�Dh��������p��0Ŗ��a�iF�J�	���F?}?V��[nXG*�)�4������OzWuF�_.��}e�:0AO)eA�ѐ/���*���w�_���ob'��#׏s��21�����`q��1�׳`a�lCp��e�aK�fz��q�l��{Ԫ�TU�́�i4�����4��F(�oz�#XF(�Dh�cY�/{��{>�v�FX�0�PaQ���!���b;�fŖe����Mʺ$�Wve��ǻ��j[��9�؎� z׮؆�4�`FE��X,Ck#J5�{��4�=z�7�V��F!��D�}vс�4wۏoUV:R]�#,Za�k�YMF�j4{~�0��3��n��Y	7�b؆�a�"Ho�Ձ��!��G���#L�3z��z_;}�$2]8��.�9Ŝn��%�mF؇�;-L��U�U����~ɮrf��4���!��ҌCf{�Xa�(�6�s��2�1i�b�s�uzց��d�z�m,!�������V�u��wR�%�M�h���`4����=:λ�������;v��G�������2�6�ҍA����#L41Fb�+7s�X�ǎ�h�v��:�#D1���͹pv���1e�f;��da�!��55�{�45�!�"d~��)�v�}/�c9y'��������<�_n{�DX��$��J!EeQ�7Y.^6b��PM�8�Ri�$!�b5�f�����a����4�6h^1׭J���X��f�SY��WE5�:�3���lCg����,�����y�e�I�bJ��]��(�)��z�\��K-F!�׼ز3-���ꮊ��uf�1}�p�"�@�ܻb�q}�+ܣ�A�!�\�l1�4�Pg����Q�b� 4K߮؆Ѯ��nv�1�R��6�Aۂ��oG`cƽ�]'5�.8	�(�W\��~���~f�JK��e�Ʉgq��e0�؆��s�����6!��붃	ƃ�|~���{DxpHm���|(���p�1��v��ݒS�v���7~�kJ5Q���p�Z�vpXf}�Y�,��Q�4F���w�F���F(�4�붖�(5�oϋ��ޙf1��h4��¶ʺv�/:h48��o<�i鈒���lCxh#ٓ��GfV5��1���h���aa��0��4�˶!�r�?Tx�-���#[a�{v��:�=��KMF�MF�c�5�d`FF�߻v�`q���D$;�f���gę�ќ0e"ຍ�ův�2eۉJ:�Ѽ/��y����h�9]�'A�8z��e�db��WM�m�n_����O��w8FY�d鎽j��Ӫ�ِ4�4�s۶��Q�Ҍ 1F{{́��f�|���a��D؆���ụLCb�Ҍ��]���iF���{6,�-������ϲ�]��l��8d�e!ѵl4�sA"k�h]�,��k��v�UU�<؆�^����G�Z~��z�ϸi*�5��AB���?aCj��JAך�u��o\"R�s8��l�	+���쪠|Sj���O��(z�%D�6�N��C��n��P��Q�g9��g�� �ؒA �eMxd�X�"�H���yU���b�{/+�O�TI �M>��H'{��T]6�./�C.]/���E
�'A����
==>�ou_K1yS
�(3t �{�ґ;~t�j�T��ߵ�Gmq��Ж5#ˍ�x��B�"i�U��\��`DL���q0[�&���;ba��goVe|!ƫ��T`�h��k�li���y�F,��uv�nݔG�ҹ%�T��!����Ue���(��lW)/��i��3�;og\���S��[��1����,IKx��3a�%2a��z"g7��dukF\u�<�?���Jbn;�%k4ě��w6��a���i����{��3�S.���pV�W�T77<�&	:��U����zA� �ρ�q �^T׈#����yQ�K��~3�@$�:�Q��%dJ""Tz�OgX�h��T2v�� {�� 2LyZ�#)���L�R�Gs���p��G���=yI�ڪć�}b��a���Dɚ�a���p 7d�{T(y��|���[y��7��3}7�:6F�B�)7g�݀�b@.T�܂:6�ϝ�� ��Ĝ{�굽�ZpLl��FJ��2��3/��\��s��<p��b��������h��4�(Q$�u��>\�A+^�Y0ϷAW���������ذRS����=[|�oS�0o{T&�3���zN6�C^��������u�VZE{lo'\��uF������ì�����U�9�{B�s� ��p]M#�׫c�ɔ (�P��,���$�j��#GsU	����$�ݽ�$W8�En#��o�RP�ՙޔ���'�TI\H$z��ÂrE�Nz`����vK�Э*��6�O�/���'��Zݺ����@P��@C��{K�-���߉C迥���kfٚS:��Ƌ�N�I�4�]Q4�Ʌ3\8��0��)(���8 �q$�|O_]W���\5Nwd^=��wd���]*մ:膂 i0���	T;O��,�(B�m  ��o�Xi��sT�NW��t8"7WH�j�R�y�
�d~�K��M��`	���dA1�.������[}y��p�Mt���s�Jg6P��-2��4��1�$�F�]
#c��� (�P�v��;��.�z@$�q����h	����]���@P՗K��Eh���������ŢS�b2Q>6�$�r(����'����&R�D�1LI!H��*n�
��@c��n��\Vo=����0v��}}t����s@��ά�f�@�U`���2��/,���M��5� B�X�n�;kL��|#�n��gU��Pk��/.0rt��D�����[�^�H7��`X ��&�I/�� ���z���u��F���]J\�D��^�+ѷT�$��]�HYѳ��˼:1�j�N5����=B�
��=�|��]�V������s�vel�V��RV!�ܪz����/{j�@Q�D*=@������tI3jo�b|��P$�ݹ�,Y���`��L���l�7�n��u�zݲu�;1���#���U��"
AR�K���7��	|
A��j�� {ۜ��z�ߠ-�m�2�
�Тo�:Ō��	̠�&E���5����W��`
;���z� :x/;+9Ow9vB��6��ޛ$ ��k�H��6��}t��<۰I ��Hkhz��4�]-��Y�z�L�� Zuwd�|VtH$���#RC3�tUu���F���)Z�p>��鑷�gU��iw$%]{v�q$��^�7��\r�#�4���wa��c��_
հ^�2���y���_//j4qޚ�vk�HV�K�YHc�>7a!i�=�[<�.c��7Yz�JI�@�M��B�k
&4XWS%�#�$�bi�l���!A��\u������q�Ǭ��5���t
���Ս���]������2n-�)��l\�s��n�wvjn!&�����]�Q�KB�eu�Yn�Y��ts�0�m�QCX�@�a,�۶:;!r�XU��Sx5�m^Kb|anS��*��������!DJ�w�K�b�>Y�$�	�uG�f=�w�A��O�$�G}j��8n�/�Rj��TM�Y������$��ĂI���rXЦ���d��@P䔠$�N��h�ӟ΀��m:�z���x�ѱ$���Q�e�Y ĘQvu��&U������Ge�
�n�u�1�DE����$�c�H����w�G���uu���}Z�0U�H$�y�O�zz�s��M�;��d�%$�1
-�"2��-˨i��#ts5��1u�����P�����ӥ�q!� 7��;�Ŧ�ױڠfL~���FID���λ'b�Z�x�<k0F0���K,>�9i�;!h'�|��/�{�N�8mR�����V<�d��"}z�$��N�P$�v�u�>:\G��Z��n%h������`W���@ ��o�oR� ='*��I(��E�*%Q)��\D�@ye
W{TA>7��� ����S���x�}4خ�,�T
nWy��B�r�B���$�c�w��
��O��֨5�������Vu,=�!;��SjAtXh�l-պ��ܨ� 0t��Q!L�k	Ǌ�0���kof�&�� �A���{�<h��Ȣs������@�I]:�p�����ZH�{v,OG��A�۳D5QUF甕$B1��K�vA$d�	�>,|&�~��h��� w,��Q�ϰ�Ow��O_	���v�iF�
ú�S��s����Z��+ь�k�ճ6-핎+m�ݗB�>SN�ꤸ��3*Q+@�!������w���}�����%㑃�pl�7���Tz�߶�{�w-K/�8,�/�KV2��(��+Q.���чtZ�Ϟ�G���݈(��Y���W��Vuw`�� ]�"ͽ�����zmN��`a��O	}r�x�tc������z7ނ�.�j�Ose<ϘY���o7�$T*"�`�������w�EBt�ö`K��N�#Ytge^vK'��W�+�y�0Nwv-eβ�wPߢ���ͳ.08�z���)F�^Q6��Q7�R�t^r��v�vF�t�Â��T���U�J��k��&u�ו}�r�,�W]�jVP��;$;���k=�Q	zqE�R�prܮv�����m�*�e��d�٬��bq<h����YW.�1�#ִ𘘧�F^��2E ��$V�ڱv(N��Rv�udm^ߩ���tҽ��"u�Ƒysk�& ˹�ή��
�4�뽡�7����B��kz��yW��w,�̫��w6�wnۄ��N��Ч�/d����mn�lYɕ�s�a��%�*}�qu�-�O<5Ք�	w�W����Ӛ��\�7��J0E��c1�$�G'8y�I��uNQ�#��A<��I�*��ES�
�s�ETDEU��� ��t�,�"eˁ9�W�$z%2�L��U�G**�����F�\�p�sG8UڥQ-R(��2�:��bx�$��,�"/Z©�]@�]�!�Uq̝R�jD;�⪅Q&QQ%�)��"�Q���+��W�T���)�.E\����R*-C�U��r�8WL�՚�$ij$P,�Ȃt�0��֑8X\����'Vr���.Gt���牤N���=�twrp�Df�Сe��!RJeL8r�#ERڐ��+��ES����^��ɕY$����"��CV�u#�1�����wW�6��{82��ր�� ���B��	^z���M�^�U���\�e�����c�鋜�e�`�k�����B0Ą�%2f�Y�$��k�k��cj����wɂ^�wd�z\	���t����a�I��RQt(�U�N{)P��=]�S��LR[�"�Q�Gc���T����g��ݟGK��{�$d���q3��Pf�ywd���A����R&z�{�;��ؼ�$���A �zcuI~��8o��)�R��.�V�]$�Ԕ:K�L���	��R��ɫo� +�| �����7�"�T�ݗ�
v�,m�OE��� �@��{���|U�g�Ն��v�(&0cmJ�)C��k!]W~f���~�(r��A�����K�����nB=^��]wvZH]!wh<�tz� {��>���Ѧ�I��I�̯W�weX.GK��	��֓M�.56�3F�[���L��p�`N[A9�UЙ��p�h����L���HWvMx��'\;��h���$��z�K,�9V��l܃���c�=Y۴�-@�y��^/����潜�qz3Lkp&{���T&�]�B����`�Q�qQ��a��sʯ�ݗ`���\�J�A$��7{�-����(dZ� ��n]�I ����X2	=W�(�����"��>�S��ϲz$x舏w-�Qd��u^$����O@��-K�up��X*T���<�T�X	|��o�B���F�ќ����0-��X�>���|�n�Hy�D��Gd�v�s��8:�F�]x#ct@L�H��e��`k؊��TJ;<V�s䷬=sٚ��<��f앋e^c�l�*Ĺ��u�Eٹ��.t�ۧ�9��'&��jLe��6��sk���.�hɢ�7Q�U:[u�덪i�1]Q����͹��cdf�ś�v�;D�,x��i�Ov8c�Nj)ݫ@\p:�
<U�5�~��>�-Cv��:=t���I@
�j�z���	�r+��we�'.6�$%!)�4
ΉC���m\�P{dnc��n�Y�OD�NqϢNV��P����%Vޏg��m� $E]��|� {��u ��&[��R2����O�*"�Fa	�lX$��� H=}�jEJ���?/d�^����V�IS��-T+٘�m���__]��GK� ��ʭ���
�í����̳Wd���6�4a*i��[�µHl,�pT�Jv�B�h��s��P��U ���e͓���ŏE
�� �a"��7v��<���J�Ou }�2ൌZY1t�z#��Xݬ.Lݬ�bUuD��-�J=�_,g�Ś��{�j��s���L`�7#��WX�N�eP&:K�����F\tJJDɐs``$}�(�-�YV���z3�9q ���U�P����%W��t�l�M@;W��26$�	�̪��;w���Ld��`��&z���T��"&�{ة�	��cwâ�e��N��.��#w2�H}�����6pW i,Eq�d�zK�{�*��k��K�n�����Ԏ���ϵ���ȉ��]\I>#�2hGwk�!��G��[A�uĒ{M8�&#$��D��x���؜�7�73
LH�	��
��w~$ʁ2Τ���:�\��,h89MLW{{d�i���[�J��g�̐�a�:1]��<-��k��+�xko�w��E)�]
��"�3Q�z�I�X���O�/^P����^\lQ��I��H*�ۛB�{��'���~� �ݡDH��ݓ�A�P�Q������O�9u��T%�d�*�;�N��FmD��1Χ"�b#!�Q7�ز>�k�Ǉ�:�1�����5x�R_+W��nٴP����ؒ4�,m�ծ�gM�����fU�?v6 =� >��v�g�ܛ�f{�����R���E*��J�w�+��y�ܜ`
���� ��B����2��v<�6.�
$]��a��8 �k�	�ޱ{͗"q���wd�ΠW!Dn�Y&�u�y�I���P2m:I}Q>$���Xs*{`��FVV�f����ԸS�V�YQ� �s,��c*^ejM̑�5<i߽껝���[hi5ݷvN\l"Dɚ���M>��qq(�x�]d}�-ݒI�QH
=ϻ�=�^�8U�C��U�>;I�sv�A[��AC�87m�Ll�j	�v����ߔ�ͨ%B;��];	�I�sD�P���l�O�,X$�a��=J�F"`:��Q,m��y�	[�ʼ��	�P$�ފ�reL�=�{ޠ>��AZ��$�@�Z��I�鏀��}'��˅ѓ����
��}~6.� H�E|�^��b�3�=@�݉>#s���H{۷Y�b�Y�y�v(̺U�C�n�Y&Г�o���|{;v��m쉕u�f*$���t ��t�m��jx͞��r�{��g�fJ��Х�&�_j�A������q�ڌ�����RިDe�r:	��j���y�P�*V�B�j�Yek���X���u��Ws7]w,t�v葁�C������5h�ZR[�k��c�%L��6�;WH�6��q�woJ���Q�"q���A��vx�����qö�M\v��q���F�Ѝ�r��ns=������#�h��&`#���R�f�K�Gj��ؼ�t(�rWO�ry��hBb�������������ؒA ���I�v���n�G\��4�T+��u%vغ�HFȕ��,�v*`��pm�$���H{۷dL`c���ϣ��Xfb�\�R0 �LQ��F��ݐH>������jݷB�o{�ׯ����iRIS߃�}�'`m�7���	���݂A�:��S=�� 1�O�_.� H�E|�=}�� G:��=՘���1��I�}�`�A�:u�}��Woz�kz���/O
Ǫ�a:�Yzcv�]>.���1�!ZD��Fװ~>?����C?�Ν�ݱd�9�H=��E�X���u����ۿ��0L�&h�A�K,d�;����<u#�z�V�3&$VU-����j���Р�}Y��ݬv��A-�v/Z$K*�7��A�}�`	=.$x���rPldu�pn�t&��$��T P�]h�	���[ĴSA�=���nݒ�q$���!	�b&���aZPoy� �=�I$��� ��Q/-;���n���$���IS��t�
��Sd5)
>�2��+�j�$�ӱ$�k��ԃ[���}���ƻh�KOO]Եi����#����X˶�������J%D�\��d�GK� ��ު���{˜ 
[h>a®��B�s�~��rGH�3�[��#���MwU
��WA+�=�H�+�z*��H'C9]/���Ͱ+E�K���Gۊ����;��ՓgJO*�T���%���Y�,h�*�6r�x���u��^�huG]
>ˬ�-� {�T(�6�Nc,J���F��u3�Nb����!nĂ|H&�U
�wm���cuo�j(�&$�1@��$�|�l[���Μ�\\O���R(��ݶ��"�\e\�m��ba�H¼��,՗m�ч%���Ŷ1u��＞z�!D����"v8��T�$��ݷ`���!��U�J�  ��鏽|P��AD�� k������i�p�a$�۪�H$��s9�'c/:$����m�X����P�RW���N���t�B��~�`Ou1@���VNV��"Dɑ���v2��#U�B�$�}�`�DgCu.Y�96�g��RH�Tp��7܍F��p���%��)��>#ՙh��6�^k[��-镰�ڴ���l���������hf���y��
��C�ˌ�;,)�� {}�� |/=j�����o|�i�F3�ph�ZE�qs���4s�3����ګ�:�ϧ��a��.~�w�}ul�|���3�A�)���`�̠�P���(*}r���	%R��m����y��	'�7����$��u�_-���c���J$Ϩ��m��	�}�<��uv�$gn��A&3�H�8�Z��D�n�=�n�`T<��B���
��3�k2A�� �=�X�ـa�$@��3E�@�I��B�][�S��1d@X��H3�Aon��C���~ ��~����2(*����ll@����I	 �/�� ����H��D�Ʋ�TBUFiV����?�>���Ō�ѝg�F���ˬh�g)�$CHH�f��>F���_��G��%=��Ʌ1	 �/�bo���=����4�T^��A����c
_AU�l��3��5��_��Ad9����a x(=�`5�+tI �4�����>�?�Ĵ��I �/�-B���!�D��������#�@���?��/�����Po�!A�������~		���$@���������/a"�A�CI��*���
�G��@����`��O�݄��������?��0��~��/ݔ̪����� ��H6}X"�h�*Q�S�7���l?7YII	� �0hK��m�9�ED���R����2P����>��x���B@$▒41�҇��~)}`��>��A|��jA�JcO��踌����"1�|�I�:Y���rJ����=~�?���&��@$�Q&�P0�R>&O���}߂����a�g���"DZH?��'���~�ھ���K	�_z�����K�Y�����Z>G�! ��M=�?O�&��l���P�� �v�H"�)	 HL���$@����Rp�i��pG�P�����o�Lـ�#�a%����@�,�@�S6�]*�	0�3b���	$	�i`���B>��K�ׅw�0�G��Hu$��䁊�$Š1�ͪM���H�qP~��~��:�}iA	 �'`�����TГ���P�ؚ?����_��3�#��>���>�|�P�?h}i|��~�0��ϸG��}뿃G�G�@��G�"����#a�y$@���_<|�������B$����1C�� Q/���Oj���������]Gԃ�`*>"?/�]A����$��3��6P1�$S��~�b���_��σ���#�_�������3t��C�c��W� Y�~�AE�ᯧ���>�2����g�_�GE�4|��5��}{0"�P?�B?o���I ��LK�T�QP4`#��U�~��o�>�I ��}��!�"��C��`�����A�W��V����� ����D#�����Z_�rE8P���