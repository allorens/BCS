BZh91AY&SY&�s֪߀`p���"� ����bA�� �ȥO����H�J�CX��Y� $ٍm��5�R�T�[e�%��������[2�aM�b��ͫmKlB�֤�Z��Q5k_]v���MZڦ��h�S6[hٖ˹�l*֦��֫5ZՒ��V��)-�U�V�mU-�Vmm��֚j�iV��m�kE�b�Qmij�[Kl� �>}�^�6���m����e���+f14�[6mff�Jb���[+e�آ�Vkm�*�6���mK�5km���V��m���# �I��j�V��z�-F��<   �>ն͋���O�X� �)z�q��j�Q֪�av��Zz��{ۮ��v�l��`����罭���n�=�J��m��QZ͵����|   v{�	(r-ʅ���oy8蒨���N=*�{�m��^]Ƕ��Ӯ�����Ul�p�z�V���R�^�
���sN�m��kw�O:���W��W�ٲe4fZ2�bl�4(k�  חڠ*Jo�v�
��Q�yq�M)
W���ެ�7w)��G��J�z�=�*�*V�GxR��9꽸�v����y����֤+��U���=�jj�1��,CM,�Z�f>   	�>��)g>����J����<T���N5�zWMUUU�z�������w��'�4����yB@�q�
"����O<z��lwh��5*����6�[4�[��"4���  {��m����[����E[�qҩzk�V<s�J��[�nm�V�z��*�K�[qITM{^��{�J�ױ炅{k�N�O=J�U'����� �mI[f ȯ�  ���Z5R��痞�x�)U�O{^�+�i����sOJ�7(�-�հǼ�{ԥJ�YM���{R�IU�R���JU���l���g{���B�I^{�k[V�٤d
��Kb�|   ��t��{;����ʕ���{{��R����w����R�M����{uʥIv���R�
U-��S�4vʝ�R����ޝ�^w������S�z���G]z�k��V�UkFUm���VJ�  _>��>�C�Z��t(=9��] G:�k��� i�=@�0��a�F�U���=(��+Ŵ��j4m����� ��p�Z�S��G z�=84w���y )��Êh �ÏA�omp�Az h΀�=�]^�@w+[���(SZ�`*��  x>�-�����T^����@f��D��� ���zU)"�z��E=�7���U����)�>     ��RU(��4� F�E? �)E*C@ i� O��JR�  �  �?�5UP4@�4i�S�T��h   $�D��Ѡ)�D��!�A����ߗ�g�'��~�����۹����sW����T}o~f��/ן\���HBI	'���� �y 	 I�I$�O�		$$��~�?����Ԑ�2�BH���U�BBI	'����$?�HHI;��_���B��0$�`I�D$��$�?tI ~؄����`�����d$� |� |�>F������|� #M"H��$� �B"HȀ���$ |� "@�$����>D���� r$	$9I�IO�! C�H!� H� @�I!��@�Ȅ�@��>F'��HH|�!�!$!�$! � H|��$4BC�H� I�0��$�I>F "�����d$�	4g���`OR���G����T�"�8K�2"��כ�8U^\�Je]�Hd��w70�[*AMRP�J'x���a�b�A-ѷ��1u��7!6�=KU�1�m�uZ����jT7���
�KC��I[M_�2�yj�fʳ�,Ƥ�#����c3N���{V�["Y��(�B�f|��ڙ����B�P��+Y�����i@�ܥJ�8�P�K�9l|�70ۼYZ՘ �˱� ȩ� �	�J��(bth�F�̛!�k`�h�H^�R�Y����8�3e܆������@J8�i,^��EB�ɓd����u(H��$�~GN�U���b��V�ǩ�-1���7�5h���&�[Ā��Vӵ&��e_�Pf�᫵ &+�Yu��m��rU�U೨:-�-���ٕ��/*�B9����&Z�8�or�f{P�E�&�qJ;0]��ի1VݭD���p�t�m�6r�5�y��vٽ�)#a:V�V�.�v�^.�{sPٕ/�x�j�,�I4�Vt=��n��m-fړ+a�Qu��;AX6p㛤��&Í��'"�\'f
jC��¸�K�֍�N���J���s	��\��N��Ǜjnj���:��/E<���]���U�w%*K7BP�ҝ�J��j1�¥��a
Ǘ0'{Z�S�CtE�q�k�x,ܛ��Gykf�P���o4�5N��C{0�tu��w�mV��ާ	r�+�O3EdںY�0�r�=�K(,ʁk{�e�Q����8� Av&���Z�U����Ƈ��S��Ff-�t�.��.��Gr�<R�#�t1�$�h��QZ�ҥ����aW��혤���M(	r;1<2��ܸAڸp� mfS��i=�
�!��ֱ�Y˷[��b4�hA��+j��촞��]�h5� Z�F�P;�p�0��qZ�ǚ���	�f@�9�&moo`��WA��ʗD��̧*x�l�t����C/00.R5&���D0=ͦ�EQj.�����j�U�VjĦ��+D{jj�[b<���'x`,�T5-!���bG���k��j��{�	i�+IkK���"*ܟ/�`a%��z�(?L�F��j���V ��$���m�:���Z��f�{oލ 9fd��W�[i4�r�1��n+�J���Q��p#�����R�1[@�ŶY�e���n	���O���̒��K��u�
?c5�g2���v�/)���<��?���h.A�F��Y��a���]:���H��&��wmm�t��,�;
�KP��e\���7Z]��z&H���d�\��.[�@�ɗ0N���fj�"w[X��J�\�����*�ۙYG^��ಎ�Y�MS�u �Gq��V��2eJ�yL1�ЀA:Y\�W��FT����z�h=DC-���h�m��`�Q\V3N�"^���@\���x"��Gt]5d�MA�6wng�[b�%,��*37p�ͫ29LжݭwX&�� ��^��#��lR� ��챤�,��&�v��oj�1a����i�ݺ��U��Xa7o�����Q�tVS�4�e�:\R�:p�Cqb;��]X�+-��
���ja�m����3�`�6�W�F[�kTp����.ѣ����Q+V�m�n���ޭȜPc�N�Uy{�.�[CF�ՔvIu	9$-4(<ܚځ�i�E�5��9{ǐP�ӷ����e./�nQP���^ӣ3H�l�&�;YSq�Qe��+T��S(k��h8����t`#0[�����P�B��7Z�G@Bd4U����m���/ݯ�?`��)��[��/X���Ô�
�6�'*ӏ&Ī�U�V��T�4����e��i�ئ3���m5�;zr&B�H0nн�~��?��Y.��8\��ҳn�)�Qʂ��X�[vT×H�si��4���5���*�I�c6�c��`HLoMe<�J֪��̢���gC�o!B,��7�hj�J�J�N	ٷ��oC�E4�������Orn^�/K
nG�-F/V��kc�Gr�'�7��K�ùS��t������<`���^�a�Z�7�f8��m��3j�9�..�sT���+˩���z`2 w5؛3s-�5�C�ګ"NV^j
Ňr�{�=
��qL�X���e�[�\'٧���6�]�f�:����ୡ�:I�K�h�ܐ��N���kUWa
�?=G�k�{]�VRz�v@rBmQ������w1 �w���5S)1{������<�Mڈ��X�Vk
��R�bP�B���o&b��+(�Y&Fu!��"S@�;bJ��f���;F��b�;�4�)��5fL���GD�ǂ�:�T��K��h��u�5�Q��PC(-�כ�Q<:A	�-[���wE�!��m}2�V��f2pSG-���=M���*\����6����?Y�a�jb���)���֯]�ڊ}1n�!)e���AX��EZ��8ƍ9��2n�&��RR	Frh
�Ϊ��ւң�-�㴍Mg�4,�t���JIs�2�]O����X�[m�ì�DA8"p 7T�Utl��da�D^�P��
�[���--dt��x��t���:�z7I٨Z7[�*�ԈB�H^Z�[�[JV���b�j�e�{�t�����Q�8����y�),Of��0�Im��$Pzs��6T��*����H/ #R�4�!���j�X�k\���W�iUb�Ʒ'+k/1`b�T͵w�\�v��Suʊ����N����v�+�Y��s�ׁ��i�f˛P�٤$�/��Ͷ���9`=j��-["��e�/e�2���Vda�ۄ��ccnee�o7v����b��ͅ]GAY�kh�h�V�,�-5I���fl��.�<�6������Ac��Qˣ�E1\ijU���t�*1 ѧ���H�%-ʇ(��e�Ym!�VҀ�BlK�$2��9�jC��Il�[a�D(3^RBe�YD�D"�5%=ه9R�0�8d�KU�!T�F�W�,�I�޽f��ZC�B��	*S�yEd�5�y��&����[�Nb�f�3c[K'��E�T]�f��&�R�ɠf;�8��Ӻ��&�����s������kElǛ��
+.�Ak��utiF��[����0�p�ʳi�6�\��5ɷ�m@��ڢ�͸�M@���u��53"��i-&��Yr n��qn��QS^'zU�� 4�Cu�K YI�b���gi�Sn���"Ԍ5l���V��7t`������ǂ��[�A�H����f�,�y!պP��n3�fR��ك3 ���]Ʉd�S$oK��}�0'�6��%M�D�@Ȓ��ݫ��:d7y)]e���+7\9���Yݽs,aT��f�.W -��w���4���Iuc@7���9�Bhi�ͬLӣ��L�i孷3FcQ8�j)j��آD��f+cnޱ�Y�+%p�F��mֽ��I�O�ү7[�:w�y(�vkCa&�����1a���h]D�]��NP0'�����Ӻ�n�[
�{u��V],!7YXI��*�R�Y�L���)5��+�nR���uʂ�u6E,.��2ˆ'���w2��@�����yM�APeX�e�M��.8UeM�h6�m&��I�����U���2=�����ET���˰�4�ff\�˫1�.�4Q�yuyf<�E�26飹�dw+?^�-&�:Fy�n�%�to+tʖ��p�&l���khV\ͭ�ef�O[���-ƪ�����YZщ�t�ܭh��u�!��n,X���.;0���6�ѠD�ŗ6�	K`/7o�(��]�4	Yږ�)�ٗ��L�jģ����S�!b���g)M��p�I�TQ8-%F�㖈�9D�����rI��ʠa/
-�H�m��g-D+��p�U�if�H=z6���j]\��V�ڼ�"�҄�F6�Q���wa飵y��\iî�UKND�[I����BZ;F�K�,]Bu�2�z�f�Ǡ*�E�v��NZ����G"ѦVk>?	�!ot�
v��g(�Te\���׫-)��J]kt��߀{QA�Lz09�j˭h�O!�k�ҕa֋�d�U ���(P�F���b��6֛[���+C��q��\v�/y�ir.��k���.k�L{IL�N�t�Sz��w#7gX�"�2�e3��t�2��_]'�6�%K���8�i�)��C.�[�m���i�bVᣳ�dW���H�GP��00w-�5e֓�\`Y��Z�4�R�=�M�B�bIH;p��h8�XI7I[G%k�3��!X�	T@�ƶ���,�m�6Ь�khکY�/w2LJ�.��)��>.��)f奔�ihH+;�
�w�r��3�՚�U�+1��4Ͳ�H�v�[�ؖ��zfdݩo',:Xef�R�a��l��Pێ^�=V2�֘�R��lg"l'�{���9����M������G9�ksm;����wRAҫQ����;���T�ԏVM�JSAtɤ��f���N&^��,>�W�;2����@�#6�­ 
XX
�&j$b�IN[��e�l���(kb��RL�J).�&�A��t�N��z46T�كm�Z�X�rBi���FmJ�n��H^��^�C����tq�f�PхJu����f]kw ��Vbn�e��}x�Ou�+�[K�Vn��%�X%Kj�y&�)8�V�n�M����^�,˓.�8N����eL[�W�I�!��Za��c®�G�;utg�ʫ� #h[O*Cu�]`�i�4�{�E��ܦ�[���Q���4�l"ާ�j�A��mA/uT�WX�edx7+R��%�+@�1Q@<t��ʁE�kL�h'q�E||Z4����o�jG���Ӵ��P�Rm
zhZ#�s���q���Zor��|�<�Bf��-�o;˕h:!i���0"�S�XT���b���)�&��0�9w
��ܐMmV-�a���Z���G0�,�����1�sv�#��ewI|v�
���<Y��*��>a�܉�9��7�1�َ�r^G�U�]�7/F�q�KV�3Bɴ�,h慶�ܐ��idVMt���T�հb�w��hv��G�e��;C,S;{*x�3�	D�՛h�VF`�HH����m��tm����*�[j��K�����2��9�e-_Qb��7B�̤֮�k�[Y�\��Ɛ�v��i|��hQm��E�+���X1�U/7p)�ԀSq��{�A��h<�)+��So1��2Mz��ͅ^�*,ր'���.V\9�d���/2�q�X.��;�7&�pځQa<l����n�X՜��f�U�wXX�����y��;�mb&�q���,�G��c���ۉvV��5Uެ��˾MWR��(bo��(�:�*V)���ǭ'��I��18�kё��+]nԥ[�308E��Boe�p��MiY{1�n$�3]-.�i��p���sDC :u��N�v�0f��ʾ��0�y�� �#��6��YWi�N��@��Tv޳�c�:q'Z�MIm-�,�St雸o5��Z�\Cp��ز`[f�H�u�i���m�*
[�zn]�K�+N�mL�obv���y&n�5�jҿ���u�cu<�k�7b�*���R�:3����+�c���-^�\�4(��y���^-�y�X�Jӂ�˺���\�vf�Đ#M#����F�D<��@6
�%:-�%:-^���d�4��j8^[{��AU��5w �r5�������{F�]iY��]f�c�v�d����֊�d�v^�(�y��RݩpS�RG[��rҘ��w��vPЅ�S�&�S�)^7�31�*h��,���,{Ch&5�K��4��ɳv��!�Ԛ�2H��\_�p7�~YP��wV�=;��N��EJ�z��d�u����mæ����pTBa!v]����֐��j��^��a���=�a��5{!�f,�5|AχǕ�8�_6s���.�;y�BRA�rLq�l����t*;U��X1���ZrE�Rݲ4���f*�<H�)5���hEJ�n���R��imf];bCC��˵!�A�y
��9l�w&M�n�ֵlt�KaCt�m��D�6�n9cVI,Lt1Sk0h��kI��ʢ�͠2^�0(*ݺ���y@����%��V�
�ܬQ����n�f8��h^�5XK��;�U���x�`�8p]���w ���
	iͱW b FP��Pm]�g��c�(�������"p��B�)W�Lxi��Ͳh�,���Ĺ�(R5}��[|�R�l��g�^]S�`l�-ASp��k��w��OEEj�$B^�ore��t˷J���q���`i�e'Amc<�����1WZ��^���Ʋ��p�}l�VQ(���2L
���t,"�j��%�bH���dē���B�����y2;Ÿ���S��b�m�����5��c �驡m�L�Y��y5�	R�{�u�hf<˺,~��:��iOі7u��ȦO��D����C ����ŷ��yu*X�(���-ql�o;�]`�-�bZ��:�pP��i�ʆ3��Ra٘��ʺ$�-�e�:a׌�e�J&:�B�ѵ��#�R^d��0�˭o5���Д:�Qu��(@K:��nf����еnC��e`3]jd�h��V��0�L�L�
��&lV- Vۻ�Nc�$M�y����A��
�s1�<�e�i8!դj��y��*�2�hQ�ʹ���P3/U�3����l;�ӽ�����flb����"�p�9���s�>6���Z�M�LwU�ƺtB́B���懤�t�̓7V4h#Yl}�|*�&����u��®�dg���ȉ��ylw6C�[�_��wʱ�e�`��zM�,el�,�9�58geeT.����D	}��R�2n"[W��:c��n�C��E���M�V{����_xw��?����k0������%��$��͙�S�A-.0;\�C;�T��u����������.5��!�����em#�7�v����ufC�[:W+���t:}\����Zz���P�s�|�>�a�Зn���Mlp���(�.58Ua��f�;<u�v�<Ͷ�h���]e��5 &9�5���xC��U:K�1ڼ����4eIl��Sn�q6�xd5/e.��-��S�+����'��B_U�]ΙMУ3iv<%}O��w��vYj����]��V���V���t,]%7�U��*���e�ΒjV�:�@$]fsй�X(̲��h�}Y�Gpha���^i��-� #w&���7ֻ:s�����j�N�TA�y
�3GS��E��U��֡���3w�=������t�)n��2�wg��c�<eJ��ԣY�"V����M.)p���Ո�iGh�)��j��a/{R]W))��ǲa��>������5vR��.�2�줛co.T�[�8�Vj.1�PXz���n�|c�S���!��d�Pĝe�eNǮ��N�#����#�'�t�.mƛ�p{�ʼ#�V�8z�u�OL{R�oF�5�F�#�Nw�b޼�[�1��cj[�γ4�ĥ݇���
���U0���׼{ܝ�>��� H��m_o1�6�S�u�شHx��a۶\ii�C1��J:�j%�ѳ�`���a1!x`]6�8����Rj�{K]z�;*±�6�%�O2�J���M��]��ŞU+19���qPb�cr�;�{i��H�w�okޭb��JG���ƚ���%��o U"�LР�]Mʙ���s6�v�	l��_ �}t�l�6��X|z�6�ٵ,�۫�vr�&�Z��U��{�u�4���� /6C3�7xc9beo%]�N��s].ɤ��ʳ��6�p��P�(�IW����9�̭����mt`�٭��ZTP�]ZD�w%Z��铍N�mH;a�J,��z$�up���[d�dV;�N`�.��
��g>�vđ�m����*�����B��Pw���f���H�����ٺ[YŤ�� 2���ي�݁a�b빀ZP������3`ݘ�΢�Fqr6e^G?^�ב���G%�+48
L�^ew1J`�WN�:���!\a�4�n[�6;�p��Db���	*�9P�r��W���]�e��hٙs%�OL��`]ۖ�Wr���Wn��| ����uO���eh�ҝ�^7%K��y����1�����#A��,��rv�.���P��6J��|�7b�;&v�:wX��4��#f�e�J�%>�b�(/_��f�-s�|/7vs^8��=J�]:�M�y����]�mu�9׊�|������i$05�|����|�<5��s����)ھ�,��ǀA�a�xӏ*	�S�ؓ45����GM�4s�j���`�5�:J�\�8��Ţ�8957OZ�Nu�<���gc̡�-x���|��Fo=$�
�Q^�]��܍��f��:�Q�S�;G�T��o�d�k��]�に�P䎓��̾�i�˨���'�S��[��\WxgC��Ym�9����kD�D�\<�ic/{n��ͽ!w7��2�K�ؐ�.�9}��σ����>�SSr�+�/�=�^y����(z8��t�Okik��l���!a�s��NB�uؿ�Tؖm�MQ,m�W__JձI�g6}�b���w�G;:��kK�A$|6�e��0J!ob&C6�)�R�5g5���2۷`Cz�t��|Q�KU.�X4ů%e5�)�On���m�(T]�buw���eQ՛KiΝ�Ƴ,ve</�)ftP���AԙTi�\�G���I�S����bU��t�}$vua���Y+�I�Wu�3I�u��Ч����J����
�VĤO-]�vSKG%8Z�w3wCk7��@�&���MR�Pb�/Z��V��w��_���l�x��µ]��a|�)�}.�V�`�NP4�q�ݴ���� �T�.�*��4��8�t���Wct-�5.��:m�j*�܍�
��f^�0�[��c�p����. [p�[�������KԺ���0I��6�V��w)��)�&�`�>1�\���6��j`���V=� g����-� �{�]d�X���Ğ�*n=���sis���,����y�^��s�^�Ű됳��Ϋ�[�;Xօ1W"q,��������]�$>g��70e�Tx���b�]�O�����f��-4rB;k#��Cj��=םXj����e<��QJ�
�`�#��F5�.�RB�lĨ�g8���	��r�ͭ�Ů�9��I�M�X���Ƭ(����q�H#{�.*���4���m�}1�,�Q��H�u�m\Y�����<�TT��},ek�#.u��n�u�G���-'�e��!_�����/3+En���mjUn�/D�;*���g 2���.���/�~NTj`m�mR�Ļ��/%t���N�uՌxƗ�]!�pcP��!�(��1
��]I��-���_Wc3�ɺn�Uْm�����P�����L)�#��Nᕐ��re��KzzC�֋�5<T*t{�4�X&
�W���*$�׍�Vl��ɡbuˈ��WA/>��=�|�耋�Rn�Z��Q>����3�I�$�t�\��.�d�F��ڻ&��vR�(T�};�m�Dq*������8�;�Y��ъ)[�\�H���:;�w[9�gSÑJ���ԯ��VX�5s��
��
�@��-��͒�u�ˮ�X7zinV9�P���&�U�u*s[1�&�UeG���lOs-��j��[g���n��6,"ꭌ��P���*�iY�f�
����Ӷh�X	��Mp�M���g�� ���K��'���Ky���ka�Oot&H��+lpu�d��X�)�mu4{/5Vbo!�(�[�NŲ����*5X�HԦc�kg	��l�L�员��0;��,�u�ab��ik���:�k=��9sB�R�,�Ncc��Ў�0�')���;neڏ?3]J!-#W�>�X�a�eΫ�l���Y�a)��|�Y�ka9��'�޼��|�8fS�0�� +����U��C �]{�С]M*�7}�����0�@8gA*��u�Zr��2Z��쁭�2�]�&��"��X�G�Y��v�oJ���f���niޝ�T�ԽN�o-�@wS"+�Qѝ��5�W#�;wE9���-ks2e��{(uLɒY�-��;mcD��ER�;Au+\6w�O�\%��(i|���X��k$3���A�Z��R�ZLp�ݬ�ݺ<z��.a��6�\���躻��B�.O�u¨�M���h���я���-��+���K��z�f��n�-R�ܘ-�OUG�H]t��Ҡg�΁8�}�ջ�-%T�%��m���5�&<���ST<��b�O�s���6�٠�]�C#I�#��\�tɦ����P�=k8���C��eq��YQ�r5���P<������ Y�_w҅�MI�9V��8]8T�wt��ȫ�V��+\��Ǆᱦy��v�	��o]���m=YˆJ���5��1!��W'��q��z<YƳ1k\G�>��St�%�ݜg7R�Ow�F�X��N�@n�{n6��F��6v�(F��x�R��9�E(�=!T�����8R����7�Q�V7k��+w:4����g�$
^e��;6��K������ҺۆT��r�ٲ��}t#�l���`�26ܝ�d}3Q7j�-�Ꮠ�)�����,����z�.�I٧6�D� �����ʶ��C��",���z�R�
&K#l3%�:�3��ކ;��m1���N"��Y<j.܏���z��zU�r �i���MV�,?[���O�#��J:U\� �q�k�v��!�!J����պC��}�iyV�w-u���P{;�ϰ�O��LͶ��0�ޝAj�+5�)M�O#A�X:��4�����s�������n��u���]�D�23�ux�P��Q4�U��iY}Ս@'�j�e�{y%�H�e9�������*�U��|c�'S�h=��зQ��i���5����J���Β�pw��*������A�|7$��UЍ�B������4d*g�;�ٮ��.\��A��Aaa��)>���Kܭ�K�Cܫ�ɰG��@��<c�����y�r|�j�Y�PB�f5ޫ��͌G���v5ulq`%�}���s%���}��9y�m�Œ
|�� c��8|�N�:���7�\�o�h]"�fA4V�J���s��;��lh�a�[����e]s��Z���'RY��`�L�ӣYƖ���GT�u0SvJvy�n�\�7�h�7�7;b�J�<�2R�.2V�lP�����p4�b-�m���κ*3lu��֥��C'�lm�Ks��k�����r� �	�e�V3���e`����F� ��n��Ѵn��o���Ĵ���Y�٘��3Gзd�z�i�AJ��iۚ�ڬ�ݎ�@����`��(�輝[�ۀb� �9ʉ��N�fG�Zʺ��U$BZ�:����*��@�r�T������^Π;*�f�]@�8T�m��sxN���r���8k/�mC,bM<���w��+i+Z��*-��3D��ީ,:��6f!ˡ��Y7���'Qջ��M7nIyۅf���q`�ݤ�8f,w�=��?]ː�ε1b"jnK
�+�I[��8ͮPP#�D�+��gN'˯2��pZ3�-���Um0�P�W���V�L��v�4p�A�A��Mm�o�=���Vc4nřtO�E�Pb������H���.����7.<쫥U�7Z-�6I�/��J���o�ȷ�#���Y�fWtbH,f*6�/o^��Y*�i! ��	zw�8-�^	VqP������,>Eֱɡ����%]�R��8B5T쨍2���}'Uެ��Ê�i�pd|��eB��'i�xU���J�][N)��i��6��k����΄Ꝓ���Ģ1�� |�����؍���,���yH����;v��kv��Z1�{t%�繓�
3olK��ER�-��*;�5w:b�4�����Pl{3����ooLO���K����o(=�Duլ�
r�b;g2;��A����^�|�l��F;��ut��nJ��Wp�c�6��{}bݫn܉Lq}
MP"��{f��J;�n��hbǡ��Yj��O�JU����et�g�ֆo�x������F_k��i]�J�!�n�/]C�05
ײ�K��[U�R��-��J���"'@;E���(_7��Ll[���z2�"��t6�r����<[�Y/A4��\\xr\ʽ�c�"]���u6�-��K���X��R_D;N�.���W�U�n��`P���l�v�mK��Uμ6'<��D���̹��H&��b�E�w�cTU-rU�H㧞�}y�"}�K�j����
���r��m����F�9ս�1#Yo]�d+�[Q~����V���6[覵S���ﲙ���q�N�:���t���5�P�~��}D�C�~�2����D�<E�&3%�Dm��&�ٿ��*��f;R]wM������]�ki�pV`�E�q�db����Ӹa�D�t���+���<�K�T\�������4=������ԥpM^����'o7D�\n�gS�ַǴI<;2r��C�����]CQ��k��F�5u�ýuaj��R7}Y�9�s�މ��juN5&�$��4�VM�YM9�gڸw*ײ��Pz��+L{	�2�r6�Of;�\2D�a�'<Z.�!���*t{��t�t�÷���!���
,k���n�6-�貚�{�l��۵��$�D��a�61� j�Uq��jf蓍p�Zz)ܲNj$v���|V�CD��1in5�)�	5��6�$7yu1�v�i0�e�� 4��o]�ߗRY��	.-]M�G���ޭm��b��{kB']v�}u��;P��$|�G��w���b��%�&���L8C�i�T�AD��m͌�6��p0q1�e��M�}pV�t��[��s�X�D@�,�q��׶���*CBM����9sJ�ӕ��2�Ѭ�K�K˳���4�wm ��Gݭ�;8�s��e3(w�0KgT�1K�ub�&pb�B��m w��5��/Fc����~�d�/�ȳs����|6Y���*۳Ɇ�$�i�)�"U�ʂm�&gd��A���E$�2�o9Ч	3w"ڔ�n�4�w99�ཷ�`�s�v��XQ��|5��ү]c�����"���:�n��W ��b<�B�r��ml�x�aG�괋�39��]!vcqa�"�j�M��
�R�+��vI6 `��ipX�r�٤���r�s�'rW��������ȉ�/mփ�k�T�0��u�-��d_+D��w�v��S �H:�)����9:f��/�n���Ü,����u�c�[�k%<S�9a,���{�e�KjoK
�<�WJ�h�Pr�Z�[��U��m�w)Պ2�M�� =$��^�W��>_h��t�
VX�駂ؖ�5��ʥL5/�1A�cr\2����%�e�S{���kE�;gݴ��-�Jt�L�5���%�Q����:N����W"�2js%u��8�b��s�g1'[ɱ�zoW)R�lq�OU�f��y: �}Ox��@�qG+%��}R��%2�r�q�(Ҏ���n�J���[kR�� �5�{�)��Adq˖\�uueu�B�9s����Q�����J���j��9��a�NrZ
T�ƚ���u�dj.ّ'*�ꅦ��d�9$���I$NI&�I'j�s>z���iJ�S�"(��h�`R*D�3]�P �*�솟%KC��9�'����嶬ە����BI�?�_�! $�O���#�}�g���@$	'���|?����G�t����T~��I��?�w3��o9u�Q����ʷ��M�����|L�Yx�w�kc�`���޳�b��;*���M�n���;�K�3J�1P>��D�� "1���Uڷi��vv	S%�U���8;���c��¦��)�2*"`,�Ã.�;�1��sU�|�y)�B`3(���}Et\�����ɘ���nȋ]�N0�R���8�l}	�wèNX���ѝ���KWbnM�i+Ł�n��1-�!�����3�)E�|w���]��Qۃ��Dm �6�����b��	0����8N�V���V��j�M�vT�S(�\`��5]��2�d8Vw.G��ʛ�{C���Z�Au^�늮:y���\!�9@����ӵ�X�;ٺ�.>�z�ǃf��z���i5��g{����șS���א�Y����<c�mk	\�+��˼�� ��d�0Ψ�̥W{��@��p�Mά;]|�m�1ȲV+o�U�>�@9�%�&�v�r�w��#��=����AJ���ʲ�0(Q3�u��7\n�j-M\-
��-�#&s8F�9�:��iQ�jC|W��ͻ��r-��alY���Ӎp�]E���'��`��ǃ�� f'x�b��Sl��Z�-�x�u7NqS˰ʼ�c�"���U��G< ��}	[+�܏�;t�lM����4Kh�Bw<���Kt-�r�R�wӞ��B�&Z�O7�p����C����&1v��m��1\��$���[ӚO}��իɏ3iR��)ؔ�J�{nl�Y	���C�v���*��W-őó.���2hm7J*��R��,���x�`M�7��V�(Yk�Hu���s)���L��e���h�6ڦΉ����&L��+.�+c�JdX���+�0��/z	hEr�Y��Ѷ�d)��T����6�[VL��T|A��L�W}��ҥGS�̇�EծP��f$��V�S!��7���P�sx+�lN��f�!w��-�*ju��#�Պ�޸\Y�#���Wc��V[�}�����	��Ӻ��ۉ���5���/ݒ��C��\t�5�1ԝ�ݻ4Э��4�����m=̽GS����:�]�(�1���]h�9Rc!λbR����S�ѡ]Au��EQ�6%��O�k}9Υ%���@
�,ov!4��Q
٩�	�JL+-Ĝ�ҹ��Sߣ�b!yw���M�]Uokn��%��(S��Y)�GkQ'�5�5V�N�jH��Y�53�����x �31�	Su�D�aқ�l-�׸R�'�i�ذ*����n�,f�]�ٽ7�l�`�Σ�hs�-���s�N�ӭ<�]D�B$�ܺ���ʔ#�2�I��$����ς�>{B4����*�+:b��n��ރ+RV���xS۠ջ�r���`���ۉ�]t��<�u���8����7kJ����tKY�Z#�:}�C��u��l��/$/V�{SR�}$��U��2�����
�m
bR�է�6�Yy�3���zӗ����N�"��$<�ctZ��y��x:6s@T^�cX���[����u�I˝���%u>�X�M�ގ����`l��@�NRD��u/ge:yI�"���e�����a�2�5��V᭕F�0�NQCk���9�J�9m��� �t�h�,.i�tKc.���l�˙h�b�:�P�}������/ ԫ̃�hv��b�ol
\�G���Tk ���UՋ7�ѩs��f���[�N,�a����e��K.�j�\5�ᄀs>���n[=r�Y��x�ks���a;�(,%��ݩ�La�\G�vi�	�O�roV��p�(]����zja��j�����s��eXƴ
�r��}K{�8@:��C^�ck2k����\0o�g�y��2�-r
s)1^7X��T�n��F�wqh
�-�ʗ��xn�f�A��9�V25f�;��73%���A����pȱ�茧r�Jޫu�ԕ7�W5�0�g��w��t�|��)eCc>�zۡ*+���V}����JQ�i#CvD��WF��:����T�n���.���1�5C���S]K6��h����=T�slK&Z�cC�wnݫWgb���D[�)F��G} RB���/^� Y��<y
v���N�5f�N\C����1$-S��g�e
�t9=�!w�BnW8����Or���нsF��X�8�M(�ل��!����ŻX'�Jr)9�e�v�d�m����@�]Օ3�<����6�}�ʹ�w���J�:�+2�:�OJ�h$����ݽ)B�b$�%�͗�̒Յ*d�]�k���XF�%R���Y+��!ˢ��nk69�p����L9|�N	L��fN5����yao�<[��fݵI�vD�V�o���`23E[�VD�2�`�hŪ�k��	�u�Rհv�<�r.�%����ՙТV��bO���
�a8&³3v��:SQ	2��m�����5*�hlW�[�;be�2�kͫ�묥ذfn�R]�8��;e1a9�2�r��;L�s��-X��ج�b���ۘ;�\�"������a��q2�k���i�w38d��/�N�5,^mu��0�k!���֚	����|A.Ifk�Z��~���E=��L7-��Z������/Vd�}�]�|�1رWr*կ�^)}�>bU�f�fR�y�\�_�Nt������K��}��?2uY�A0BoH�:d�[���{��rF����^lf
�:�][����m��=����B��^'��I+6w�^�|��9X �ބ��G��W+K��NQ��NƓ��t�y#��~��ڥ&�fs�Z�7�'{9_6U����.V{P�k���s{Эk�G-gM�|u�3x+|vY*���\�0,BKT&䲶��(ͺ²�O@��U>��*:�%�f�˥�����[[N<�����&;���r�t���݊mS�W���ݐh�B�}���V�I^�.⮺���Ք$k �$�蜳��O�-�q>��:Y�$U�S*J[�+Eu�b��]\^�k�OEG�=�i�W���Tl�̭@�sj�V��k?+�[6I2f	5+���K�.>���ZN�3�	����Vl��3)R��`l��a�7J��*��5
X�F�v7�U9''C�nevn �v�r���h����`�BJ)�T��:�*-�v��e`ݧ�p�0Cn^A6�O/4���jfNx�t��X�t.�>�q�eG�J�ގܥ�7MAt���2u�����x��K3�	j�sJ���}�X�8zɍn�G��,��D����)菲૧�f�`��|gK��:�+0�ut9=���}�h�\�����=zM*@ugmţރ�w[][�����ד����YN����gK�k�45�h�a���*�QJN�p>l.7L݊Uj�.ܓ�
�tz�en=�\R�F]
�'��j<���}�N��ӅIKb�+Y �`��Y�6����3:�!w]��[�5�ݛ�w���Mj��<p���t:� ������M]X�:"M�*����?�Y���,C3-\/��r��X�sa�ۇ-�W�&�l���kB�/q=b[";�¨�sk1(c"�q�Hą_1ppTR#i��_�3XF�r��dR_Eě��v��n�n�{X*�T�᧲n��S.0_1|̡u���Ԯ�bOR�]]c�ʣ"�1E�:��:���{�PՔa��ޘ��ST��M꽱�Z�X�9*oAX��n�����N�m1���ܒ��\��ޛ�`�oX��Qv/A�ɔ��d%��z�
�Y7�EQ�=�`��yFEf��i�ܨ�����g�u+���mB����r���nъEј��j.-�g���B4u���;XK+^��4��>k�z�9���*�uMqc�},�@M�V�z��S��QR����|�sժ��ćuq
!v�fU݌�V����g\t5�̕�m\�\y]6[�E�F�r����z�h�m����8�Y2��'����uK���q��b������rm�6�uͮ"Q 8�h��RW�뱎N��6��.h�Z�R���M�
�:{tOS��RoK�,���p��d��&�j��ǉږ��Y�C��|�F�aO�ᦄ����8go>���oV�{#{�7
�rĊ��tXCh��w���u���$M���D+VB���٭80-'�o3��%�ռ�	D���Y[����R�L�� {�e��*�|�,�n���W��&�frV6�h��F��x[�Y&��^� �Ү����WX�o��S��L2ӭ�,ënuf�/�1�I��;#�e1�U��p��Q�Y�#�ݣ�����-N���Ʃg�;gKsl��n�gP�w�nu�@gԺ�Kk8�Z;�pQU{��j����=�Ӥ�����}Z��GN�֠���Δ5�%u-���X�*��v�	[%Υ�Ư��YV�
��%X�T��O,�U�΢�D���kڕ������]��:n���}XJmfl��IՋ���l���x�}w�5��7��s$v �u�o������蛄������wv����ȍ8^^�"z�sn������L�,z�3�Z���݉���IS��l�qi��VN�!n.�җ�=����Q^�X4>�D�������n@KP�{����\k3�Όr�F/����OJ�W�R�����ƫJ]3��Tt�R�ȯ�V�t��nջ���YZ9�x����L���`�<����ż4�TZ�fJ�ˏH:�pF��k���ϝ�7������X����W	�a�Dq�|#kv�H���b�v�̜6���weZ�8b�%��o}֋��w�Wr���<݇ssh�ȶ�+�ʤ��-'��\3:�����Z��A�X�5�Q;χ_G��W���QA���D���NT��!�Y���6��J"�&޷��>)��:�_ә��+ܑ��$�&_uL	kM�4B�u{��I�;{��ٗ�����H�b�ܻ���b/���e�]6`BcY�nW\vݓ1au>ki2�)��s��P�w�����M�̵`C��DkX��Z:���&�f��o�u(�������ٗ�	:��2<}$	�D��]`��Yp��7�o����h��)T-�YO(;��0\vS�j��T�$��7�J)���9��.������3-�FG*�X�pՑ�Z���:{��ĭK�����i�+3TGFۭ�1�ٛH�,)��r5�`�g�ҭ.�>�QX1̩����3�[��C�V/�j����8H�ra��(7MM[�؄��� |y"�u����8W|6Tȍ��F_3�F�	�m��w��4�G���9c����S�n���u�8:�%R]`��Ts&1G:u]vg+lR��A>�wX�v�~�y��|f�ġ�%ёJ���NY����g\2��]s'JLg]�>�	Ū 芈LAn��#Y(����f�C^W	�K[���v�8��M�{f�t�)3����D���Ӕ�^+F
��9
*N�!�%$�-s"�w��ф���b��+���sL������.h\]�d�L�:���A�v�������JMܮ��ͶM 
�����+��]�5�f=�L�/0����SQ���,�-M�R�$3�Ij�4������e�I7�j�Ŧ	��k=W���+z�[
��m�ӭm�n��ϩ>��܍�n9�Mf�w���J����{}� ��r���-@-��;��k�=�E��5ڼs;�U���'�˦ ���4fL'��#�i8xɮ�Օ��
�bל�A�(]���N`Ee���]+�����,
�B΋1h�:٬�ύ�c�)��hg�TY�۷a�C������þ���Ǝe��TW�̛#[���o��P��5���8ɻ�ʏÎ3[of�&�F��2�aU>��F�-cn���Q��vj���RE�2Q�7�&\Ω[Pf�`W�WD�EÈ�/Z2��[p��1�7��d�NG�4!�We�'ܙ��
�*y��;"��ʧ6�s��oI:%�;2�L<�R�v����+�J���.D��$���+Y�'M�{\�3���)J�EN�Ι�Ɋ�Κ��Q2�/$���5=�=O�qJE�ϗnQ9�KeN`�|*\sC�77]��m�;-I�&^q�.���-��;�/c����T�-����f�#���!���3i.���|b�+n��sfvk����;'*4a��0�����ǴJ�|`��RB-j�h�@�t��� �9ɛ�麛`���6���R���C��{#-��ݼ/V7Y\��N��RsX��y��ˬ���$�����j�@TCv��Ų�)��2լV�U�i�̥LiGdZ8�9lP����-�b�3�����Ν��@�e�}i6�͇oPb�� �q�P�D�����T9t�/��%�'�u��$Y��;��&���U������B�n�F���9�L���|Ӭ�{�Ȩ����C�ܫYTX�s�u�hl�q9-�$z X�i���p�Xt�ۻ��ht��R.����u�v����j�l:mÓ�bf��^u�}}Xm�1I)���>��`���n~KH�I��b̛����bM�w�5��:�䙷Tt�U�,�)'e�{M�+�sSY�Z���1p�g,̦�`7�����B�E5|������*v&n:u"���Z�J��;u���-�ܫC���%ɇ�z.�n?�wKY1Y	?�8�y&����r�w�
�Th�`�"���FgR��V
V/R�SUe�W��B�B��h���1��I��rf��i���.+!�q�pyנ�֚u5�e��(��b�kɕ�4_#E+��5��]܀<7b�[�>�-���Y;+%f�M�Ekӆ��K%m:�6X)��1ocS���|�g�^�����?�����O�C��{�_�'�!��|�������>��~a�~���&�I$T����v��S#��hJs`7u���y�^�ڻ�{��*�r2E������tu��mi$)a+��kUB�^��1�.o�Ԯr���)(L�	��Rs6���<x+��ln�Q�e!�93YKz��z:�ӣ)�H�Ov�#S\{�x��u����_S��&�[���#��m��{��\��6%�_q��8�kx��@ǐ��pا���P�|��wV*[v�doQ��@q&�-�,Rǔ�e�J�(R�y�ۜf�n�S��J�;��"<��"��D�r��]۫��9A-[��z���ӗ�["wws[��|��&�fm�*E@-��.U7.�T;��X���D�]Y��E�oI��0��ws���u�O/eӹ��h�:���9��v���9o�3�q��\um:ə��(��5c��Ta�P:��DD�MZ{]�lX�ks�v���)�״L{%�+J�ۼ��3-�ٝH�C1Tpk&�r�VÃs��r��6�E�j�dx�ebSr̀l�����y�d\�iV���;���7N¢3�P�:.��eZ���Ә;�Zn�/�x�A|�|��k�.T�c4lb3m��r�q�Ɗ;S
r��a_6�.���@lc�똆̙Gb��1�a�s�>�u��)r�;�b��\ܬ7ӣ���[m�͋i9&��>;� U�H���Y$Ю
ΡY�d��������^�� 6���@��I�؆�R�K�i�*d�^��ZZ�|f�a�S�¹`�S�l���8���%�
0�lS�@��d�V;�S#��E"�����-<مJ�kR(�S2�d���R����ZN��-E���kFUV��\�QE�M��M�S"��ʊ{o(��1|�u�[2W>[Yb��K噇/1D-�z��/��9�9�x=��*yl����sl���&jV{sYQ�Pkm
�!����1`�5�JX�[J��,���S
/Z���B�h/�z�>�N��J�rhֲ�彵����,�"�.G<�"��e���T�N-��+TF��̬Q��Z��mm֪�DOTx�R��l��b-J��s`����E�*�zʨs��`����]�*,�R�������U��m��Z�D��ձڢ��U|j#*V�o�Vw��5�%�V	�
&���<h��꿫w�X���rQ��N6�ɼ!L��3��Y�X��ŽZ}W�2Wf��,�u��u�)&�yHW���,\!�HO�y����wuK��)u]���P�eJ�^�1ޏ<������L{3$TI�����e��N���g��9��4�pgO�o'�����FТN	���5�Gl�uqɼ&���g��xq� �glq����5��c'xot�*�_�yWr�������E�?N#d�ޫ��	�ݗ��0.�����N�֠��J�C5���r����;�N~
9���_�gy��t��%��j��xe��m�g��o�SQ��Uc�[�^~��Vd����I��<������p;,f/:�����,�}L��S�_˙��r'����'�V_��� �t��	�G<�j�;��d�Ji��-{-].S���P9�d�9~1}>:��ufe��$g�Q��7��+�<������u��<Y����>��v�b/Ey��	����;~�����b�[sM3yW`J�W�̴�^b�t���S�*��өI�UyG������e>���w��suu����0���Jfp�	P��D�)��N�zd�nRƔ$9�m�{��7���:J�7{9��
�_.x�ȶ�}���T�{ySc��=:G1W~��C�9uE�8)z{;��r��ei5�elx�sn۰�3��ۤl�����t�z��}�,����h���a�|���iι9ï�|OX/t��v��]^�*��Y2z�n�x3'E����&Fwq��p$���E��͍��@�^�����y߫_QO&����-�%xۀ�^����������6ħ����Z�6;�1�=�t&���jFY���'��;�q���z�y%�챚�x�^4�ØO�yG��3~=����*����>Ξ�*C�&�s�/X�Wz�{��oK�����9�M�M�~Ư�OD��'V'��|='Zz�{�Eo�u�{h䝠;&�]q�����6t�W�x!q�G�1]�*�=y~����X�;�>���~�J����yy�1��sĭ1?W�����1Q�F�®ު�"2����u�罽����ԅI��[�n,P+WM�!�m4���;f�罵{�o�Ĳ��&VH��d��`
LX�/�u'Bwk��ck�aF��J��aө1k�:�Ƌ�� ��:^sc[�wYJk/�}�}��� Q��[��74�̿ol��t�C[~������I�޴�z��o�
�zM����E�.~��'���_�ы�>`u�g*ɱ���)]ޓ�����"��pހnǜ�H���3#��'������J�z�}l��+�|0v|�e}���]�\�u��=���۳����Ñ�{G	sGpoN�4��}��84,��q�~�(��~ͽ%8)h�������NΑg���l���2;��,f�M䃞ʃ�Gx`�K|��̷�ܮ��J\^_�!����=5}G������)��L�
������$����-���p{�1A7+���vy�	��g��N�/��YFՎ񺸯�z���SĬ�6����!&f���B4����;���P�\^�H���t�V6nU��|�<����dE�k.��X��,���C��\�>��_b��t�G��}�NVW�&7$��^gN��o�ۑ���E��G�����)�u���c;H�rۿ��y%2���u�SכR�3&��,����B�w)�yR�֗���'f\U���X�U�?��vR�f�����Kʓ5l��䢱�?��Rϩ����H������:�#�v_?d��,��������gsS�9m��}���Fhq�����9l�vP�f���6H렯|��z�V)i#7��7 }���Nՙ;@����f�*��ʿ/t�zwvl���9�{+Ϩ���f�&P�躧�&�录��^���.�2��}��Qn��|�ˡ�eA�Q��|
��Osǁy;�����<1���Z�$�Ea���2���3)��{��}<��q_ �t�ʵ\���r�$����w��_�k�z��ş}dR��G�t���\3�`P�C�_Oe9�o�y�z�v�������!�g� j�Q�y<��-�>df��E`T�/э(6�x�q��n��G5������-����_x����x�Ψ���%G^�o,�:hL�}���6X�V�j�3�������ͮ����[Z�S���z�U{���9u����Y��̎�;1�r��g*����I��A�W�	t���{����r��_l$H����2u2��a}�Jq<[v��i]7�%AdU���/�#�M#6r��l�~�GB���<���Z��W�sc�  ���y��w?���?�AK_R���������+ �?R�^Y�;��^t��b���+Z�b`:�@ci�B���Z^Nm��+���u�Z}(�=Jm\�F��M@��ʜR��{3F��p�����p��:usFA��J���e{�^��ǯP�_�V!95;�=���f����g�ܢ�����ʨ��ޜꧽK+�_g�#�a�=�z�X��c��v۾�.�$v��7Oq]S[C	�� ����n���<����9�%�+]�V����2�Ϛr:��Z�|Z=7=�泸��fN��d�
��՛�g�]p��rs&�<����#�n���:����/���ONe�uތ��ܜmOauu�}�����r��8���f/��!��*�Q���{��X'a�ctAh�e�a�D���6kf�<�5�DO��I�,m������B:��jW���5l�T��_]�4�`{4k�د^����l���� nԶ�{B��&�j!�s.�Z�`JT�l�y�i,�8�v�b���3;�B}q��q��v(�f�vl˟=\n��@eb��b_P`�YS�	�f޴�(�]�����ydr@v��8v�/�گ�O���c'p�h$�����7K���G͝CT׸|�d�/���ο>��r�I����OA��{���+�u��v{[���&u��?��e���Y��LO��;�������o9�S-A�Sκ8�J�Y����}Wo�و'}M�y��p�߹�+2�����x�W�o|�h�O����A�az}g��W��K֩om<�T�����龑����ʙ�e	�O�/�J�2���^P5���=|�s��ypr ���{Ga�x��=bA�2�4{�d8�y�3w G�ݹ扴h�'��1E�����I��NiƋO�)��6l�k�vpR��͙�o�.�\n�ze^tݥ�^�P���r7E1�V�(��єo4�V�^����|K���Q�]yGd6�o˹���+g���R"���7=���w�R���&��	�j��m$k)7����`$��X��e5sb�Z�y��DޭN뛝��_c�#uf9����LE_>�+k��x������ڟ�4�{�-u\�|�Zo��f��ڃ 9�����r�1�};�VfT��Pǳ���߫z��N��>2/����v���HVl�8���_-g<��Р�u�9*z�+~�;�ܵ{I[^v7jo���;>�{��A�=��e>����a��rrx��q���O������A��d���c&�����&j�o���=2��E�=���9��I�}QgO�_׎�o��o\��V�����~����=�K�zL�w���X�8�|;8['�V��`��#�
|�f�/�I�����x�{+��s[q�����H'q�zF�l����}و;������#}[n���߽������0���X�~���� �f`Y&���ko��1��Ūu{���;%v�����>�#���np��'�A1bz]y�]�<&	�m��t�}���2�z6��9$��<�>�;�C���?������d����g5�\���CVeJ:pl�`lk&��)w�u�.
k�I��ɹ���׸�oy��.�.� �H�ui���-��d�Om<�E��鯲�#�'�'>�ᒃ��1��o;�^T�PUi�B���j,��7R�Yx�)'Y�r�%��-,;J9�[��ئ��H��w>�ײs:w��4!�����G� �=��,���C�����B�� o�����R{�Q��N����2��-o�S�#��X�My ��Nf{�8Vr�|�ux����J��KSn	f�vON�C�6����������6�="�sO�k<��;S޵r�{=��;�ɶܾ�㮈��c�$cΞ>=>�L�f�oL��}�[7����[�T��W�L�s=��hu&�r������g��v'��u���$Mo�p/Ӹ#����k9���S��`��v���9u��zcuY�{=u�o��`��'7�{���C��o�v|�5��b�]ɢ_��q=�r�:��m�WP��My�Ms�M�M�L����"8���t������k�~�j>����^�!�S���ɽ���V��j�ݿ��q�oG狆�֖E2�M��!� �kWG���G�Vgj�Y�8{",��ko�%�F��{ݵ�=~�~�f����^t>1���v��+�M'_M�]�D��$	@�A�IR�.���\�J��SFn��\�u�	&�}�FJ�h�YJj���Vt}r:��?|[����x�6�m����x��02��W�Ts�����vb���}]�z�wq��Z�� �X�Ͳy:2�Eg�}��{�V���g��7\���&}�og���Ƈ�S��/���͓��ْӯ�ɵv�ߖﰹl�o���6��q���Ã���(x���b'}��z�4����^�K^|�}6g�Ux��ȴW�o�zU㳶���7�[Υt=Η��"=�闣��*R�~y�t�c�6�ڵ����Vz�z��N1�6����L��GA������^t���ެ}���:cx��k=���#�� �:�]{�{j����Nй����I�����G��y��]��G��d^���&7�~E�Ivϳi��sK�3;�7��D6�K��/-�^��ghY�^h����eCM�@�3�iܬ
{���Zݵ�VHڲ}��T�(��KC���j�J�pn�=���W�V�3�+6�¥em�p1�s�v��$��� u�n:L�Lm���o|�Fu\JfiJL�W�d˃��.�]dX��_��q#GPmM�A�)���qPY�#���N �X��j��Hs-R;�G���ɻ�;g�g�Fv=˗���kՋ�m��q��pnؑ�t��gJ��(`e�ν�o�=S-U�Y��Iس3���Wvhf_���`��`l?K_q��k8=�k'e����ug���~��ySr���(�fKG��kԶ�hd���O˹�ʧ�ҏ���&D~����^BE���ݻ�7��Q`��Q��՗��>��\�П�5�N���^-��4��֊�!���|�5���N������im\���nL������lF�F��3���)��U��[/�ߪ��G�%�L�W>��n�����̿k~޴�:���Z�ص�<�-<Y�Z&O���p]�O�vyg>��C�g�`z�H�g�����T̓(N����q��G����g���/�*&��>���M}��vT��U�Z+�>�����W$1�Eo/*�K� �cWf	�S��
��\��ۥ�0G�Ջ�1L�|^�����t���R���p�&n��u���2^&�G���LÙ�Ch�\�I曥9f=6�����BJjgn����[Z7�`[-J����3QU_I4�gk���� ��V,�Y���Xo��ט��Ϝ5݇4�19���ۚ��w&���|���щ�BeCۨ��Y�f�i^��u������c#V+⵬�3��(�yV��ܺ�������0z�!�1�2�Z�p�1\�8�le�3W��[R��k��ZzYg햣F�ٕ�,Δ�ǧ���!lt <]�Tv1|ӪX x8�e�,kn�[PYZ[�;���oF��hW�DY�*���ǄY]��s+:��<�W�C)q�ټ]���W؞��]؉��b��%/z�˝u���ޤ��;9t�B� �f�R��V�����jE͝���F��Yy�{qV�p(�ԉ�6�cvgm˥y�'I�{6]���)���d���p�j��TpnL8^�v�mn�κ9�n�-ʋ�إ�t������G�N�:4oJ��� Ƿ�|y���5������n��d֥��k&��7z-����W/��/��֜ڏ6�$�kn<��˩��KR�/:�V.�����՛���{Q&g\��W����E��$MW���GR��XYd(Ġ:�e�u)v<���v����)�u��Ɖ�Ժ�Թ�~�U�M��ӊ��tJ�L��t,jM.���.�ʝ��'[2�Y)��.��&�ʰ�cL ���1V�w�:4q3h5cx>�����艓�]i�o{�NL7�7[����q�����eN�2�&�e'Rz����@Ձ�KvZ&��$���KL����Φ�w�p��ӽs`�d%��e^0x�.�Mݐ��ИrX���L�\-�+%��Á�g�7���˱Q���nt�m�ئ�ܴ�n�}"�\i��U�al=r�C��aZA�pP>{[�cOH⻈2U�b���cry�R��iFМ:��:��J��ɲHg]<��à]5�H�6yh�՝�R��
�*���+�@2��	�۝��x�C�6_&����;g�����f�U+,|�a)\��c��G�Gg:��^��(m
�%B��&�8���r��hG��}9V,������$	2��ѭ{��7��V�3�P��/�<׏K`h���/8O6�l�W��ܢ1�5�� �2��r����S3�_Agۣ��,��K�D��ՋEt+�μ���kco�x��
b�ٺ�yk%%�u�r�/Nwtq��}kQ`�(�����1��E��wY3u즭�wAhmX�f@os��r:�[w3�hhJ]�m"6j�Wj���޾(�X-ͣа���ڜ��钲��΋s� ���l*}�o�,K֬U�l����nu��m8�nq�O���P�if�Qh���L��-��6�ƍQ�Ҡũbq��R�B���ȵ���KKkDm�
[X����n5�m�}��kW��aR��YSb�2��+=&As�e[(��
��#2�����VZXT^Y��ETE�K<����2V��rmb�婭�/ms\�u�KJ��)F/ƺ�)��b���F�DQ����T�X�,�T��:�Z��Z6������Y�Q+X�m����z��lV�-E�͈�b>&dP\�Y�6��O�a�:��0��Wd��mZ���W-�e[Y��]aZy�kl[��S�j-ckmA��R�ۄ�+�����Z��a֞'9Nm]b5����1-
�vJZP*�n\pg��J�%���kkQ�|�'9P�U�����є�^s"M�T��v��o
)mכ��j��Ky��֪
��5�*��x2���q�Z��|�y����mh���)�^[��^`����8�R��������.��N1ff�~$
 W�v��}��c��#��k��Ql>�y���^J�l%6�e؇��8����3d��wJ�X�D�`������\v[�#o'd��]�^N�k"��ol�D͙�k�(���(�M+�薒����lު���o&��~M�����v��z�ijIu;�f�ZF	*m8zn�>�n��y�y��'Nk�sO��w�����-����]'���9�>��ݪ��Ɲ��>R�me�[c�
�b��U&=I���������s׋Ӿ�q���}���{�D���Mz�C'�}��S��C��-�7F�Q���|���fT" V�6��R��Hj�Bށ��HYu><�U�!4��8*���%����O�ޥo��G��^�ɷ����	e���SL��@�8K����G���HҾ�Ի&��(L�%�ܪ'��&?tPT·�	���>j�NV����*o��}l�vS�虲��⓲�x�9����g�w֎��~��4_)���ʣ��E�'P���l5�������|c~��5�2���g|ఘ��Ld��ͣ:m�����b�:�O�T���f�1�ur ?
��#�'�G�f~��������}�K����.C�6�ɶ���=�ʥ��^?�W�~,h�I���rsm]�(5�/�kG}|��$l���KԨ���X��Fz�_G�v�ܛ���9iu]���+��/�"�ٓ/�^:��n]׼���cݒ�t�����B���TT�_Fv�ia����6����Y�_M�U^�b^��L�}�W13 �&V���2��i&�pD@���@c�RđC#W�j>�ё��3jY��I�� �# � k+1T(��&b��}#�G�}�D�_v8�712Y����lV�ԏ?��N+�t�������^�l�O�@��ȇ��L(�ZF���	Usc����~��+{d�Ķy�=[>��q����ܼy���_�#��3�\�.�B=�}��R�|o�.0��ؿ��r�� ƛ?8�FE������8������8l)����jI^��W�/iWO�3w�����G͂C�uC�}�+F�d겓�x�wJ�SI��O �Q[�¼�z�|@�1�O.���mL.ag��~�&�Q���H�c���t�Z���~�u��sv�t�	7�ޗ���^/�6N�W��z�/��Q[��Wr_ٗn<{��i�;�j*^`�������g"٧�+�g�fϢ�n�!i�o�W?�c3X���&��q����6NMd���q�Z�A���:��gh��J;c�2d�Kd7������O۹du�7�>��N����au3.`���\�1�e�@Y�/�
��ʱ�5.�-@o�q����W#s��%c��D֚b�.P�g�]thW�״��7�%rP��u� ��裔��3;+u�djT�rU�k��!j=������F�3��V`X�'
4]��0�Ӯ��6�\3��(�uy&>�h�{�֭�O��ⷷ����{��(�����~�􇍖j�^k�1�=5����e�^��N܊¦��r:�J��X��>U�����_��^��{�<��~�=�gJ��E�<B��	O�+���r���]��]t�!��.��n	ˍ{w�q>�� �2�2��H!���;���:K�g�|��n���s�_�ݘ�~���,��z~���2,����y`�5�!7F�ا�.Cw=yO5,OHE�[���-�t{�U&9T�)�L&\C��rP���qi�- h��6��j�c�T�p����s5�U4e�x��
2[����:ҟ'gk�l�E�8�n}Nu��km���Rxn�kBb5��	�E͊�t{;x��:�C���P��Gs��T�qK����Ŵ=��\�ۚ�l��4�a�.�d�_Â�P>j�l˓��yq����cq)1poؤ�m��I�b���&Oo:/V������6���"@����,��S���qKC�ح޵���Ox��eRyO�H�sP&�[F��������?B<����]��nt�%�X{�ynٳ|�l/��8m�۹�7�L��η`L^m;p�r?r�y�H����]*J�*P�R�*�aSkj�k�o�o^�c;[6&�9��w�m��:-����3$�z��
i�rjXTr�PI��8c�]�XT�=��iY�X�_#�P�w�8�g���9�V�[�٭��GEj�Gx[k����j�U�W��]�]7��
��y&9;��s6�-"����(Ͳ�?d5k��7�Z��yg<�B���������"_��޻=�����Z^Jm�ZD�.���y�;���r:�����7]��ޔ���f��yT!�X.f��U+���r�$R���*�V<��[�IɇC�eϴ1Y\=~G�p�H�0�����H�@nW�}�S��*���,��b۸y�B��;�u�R�g�|�}��7?cH���a;��G0����R!w#R*��^�#l�7���31~�aVk�3���`�d�c�MS"�;=�0W�2ڬ�G֧�A����xv+�νnI^7�r��l���jB�f�v/	��n��ן�2N?_�������J®���L��^/�v���}�&]����m�nςi�rGgR��))��R~k����JV?4'�T�e,l*�r����Kep��S�a��,3�c6��e���� _�"�U�ӹ.������b7���%��K{RS�8�|�����q��c��y���s{v��Q���ӽ��i��n���yk��p��y�z�g"�Z���e�[�Z�f@_a�ؑ��z!���ڂ��D,�}��=��yj댁A5��K;."�wF�g��7�_f1�ZN�pô�=��'�tα�6����m��n.�����3�žu�aK�Ѯ���3�g!ހ�g�lU�:}�j٦	�(X'1�@��e��AZ�����߲=��� �.#��=ͬ/��9�Ӗ��`q�Ơxz��Aðز�l-v��gj�\^>�8���]�7��&��/R5�cUWc_�%D���#e�۲�Zkě[ɶ=#Wd�ϼ!3=T��ƶ"��AO^�}ryH~�R1�=��.��_zKg�(Wz��xf�-�[s�s�q���n�1�f�Eo;�h߷��+���m;�x�K�F	Jm8}��}�!M�7.f���]�ˏ��t2P����$I���������sn��2!��N�,V:ѱky�]��"6y瓰�{�Ѻݍq}�"�j� ϰ��~*Ϻ��m�n�5��x&���G2�fHm�'�M������"+��xa/jG���H��)�X�?+ս"ħ�jW:�r����P�&��ɳAYT�k�4]��LE�G�l5V
���}Ғ�ȑR��fO�&��>��K�
���y���ӝ1�OMq����K�5�Eŝ�P�����X;2"��DA�ܣ�2��ױ��=�,��L>�;ƺVL��rγiv�M�d�L��i1���y'C�@�gi9�U��Coz��X ���v�*�xwh��M7�#���'���k��)9[[4��{)X�w5}o��Lۏ��c����/>��-�ڀ�R�CE�a^~R��0���*-98P�Y4�Y\����M��a�Ϗ�wY�ad۫�[���1�����Ǖ�XK�ْ�1�gt��Z�o?�y^�ܴ3���g��m�~j�#-�ۑ�I��6A�=�[�6D'ؤZ�g���nr�h�ڐ�������U�b"䒴���z�ԁ���w�N$�VE������@I|�a������"�%��:26����Cp���M)��,�����)T���F�����歭X��ڕ��ݍ��b�~.����@���O~q���[�M����JJ��#k!� �;�Ƅ�B^{q7������j��2�5�<�=C���N7F�1�d>�U�S�`!=�';�m��Z���H�`|����3RZ�_^��v_=���O
��)�ͯͶ�U]l�W�9��R���j�ݮ�	_J`�ak�^�����J6vF�Oۺ�,?&:;N'�D3��(��pX��R�3����[��eF�j�����=�E�Sҩ8�XrL�į7�4��f��M�z՝�m�eI�Zř���O�}}A�q^,����yM�o�3�C ��{،G�,6���L��}Sl_k��tV@��*���W�UP��"ɣ�'�4	כּ��f]�6�Al��ag�ol&"�[���!5㜫������nн�<0��BN+��Xz�@ud�g�s�my�f�%u��wM��?�$�֜,事����������gy�ÉnC�hu�Ue�c�>�v��S}IGö<�1�KT�!�����M	��.�.!�][$p��%z"��6���SP�w�Ԭb�y����ީ~�S-�x|��3�)��o��<�'l���7+�i��W	��9���>u�\�=�)?Zܡz{���ګ�y������S}-
p���-�����j�,�z�����jeQmr�S��T�k��*u4��U��b��v^P�79.�}JH�UޅJah=�ƃ9����n��42.#T@'�D��>M�΀}�I�$��,�����2.���T<�Xk�St`�.xb�箛r[��.���7<At7�y���e��0���ꤧX���tu�/��L+sh�G<I�,�qX�Q���3���}q����eO9�z��n�k�+4Y-�c���^�wg��_�Bm*�(���ǫ���r�'�&Df�vZ�������E�@�`�#�6�M�zy�(����V�1�q�<Ma�\����<9�l����[KlO�Cw��lQ_7m)x�&i]��Ǽ�NQ�Xw�1c�]wLf�Isj���w��--��݆$�s9�5��M��NZ���.����8��*T8�f�'�Z��~*p��W/,��S<���k2E;µJᨃ]�_ǈ&V����-�;QL�3������XJz29����h��Iky�ѭ|��A���A�Wr��f��V����k	�m�
ϲ}g���lW��-�*k���C_��.]I/y�b�^�{���Oٳ�Z�1�����	�P6�kۭW�#���_�2-.�$��-zs���U�xkb�,��|��7~��Ϧx�[�)uc������C`Fuk>�3,���Ok�:.��x^5�$n�z�0S�{����T����\�d5k�oI��>��&D�c�����h7F0vH��5n/uO6Բ1���槹�7=�T�ɦ����N�ko|=�����<=�\��Pѫ�q%ƼH��!2��>9����o��Z��M���u��k���)����x+i��(�WN&,�뀊�ʯ�~�ɯ�7�V1��������Q+�+��bc�����}.xY��ȑvp�q�Naq�z���U@�G
�4w�Ȣm�?R�ڏ��y��z���y��3��Pd�k�s"��t�q� )
����W��7��3���� ����s��m���Ρ�J^X����8&�	<uÌsZ�ܛڰ�vDy�f �a�k��2|��ͬ7͇|n�M�O�&��<< �i̍~Z0��߁o}�3)��|�S�j�d\�(�7_���H ���/ ��:�5��2���><%�{Az�3��iݮ�}6����K�ߢS�W]&'T�l�\�}��k�,"���O�R�5�4_�k+���@��P�����4�^Cϻ�"ጩ)�TQQ��?7JS�����mޣ2�k�XO�j��3j+����NO�?�z��Ѭ����e_zՄ��Urt�K����Tcf��ʯ×Kf�}¥ws��H�qhX�����N�^��V������a�w V�U���<'��	���9%�sz��9��LX/� (�j�
1q��&��[ҕ����=����^��{��s�[��U�j�5Z�	.ƀ0���|ز�l-v�Ȱ��ռk�\]7��gQ����<�L>����_ˁ�k
�l��n�
Zg��ԉ��'y-_��85�w���z�-[�X6��/a��Q�cT�'b��2�{ｽ�L��!���=�F�V�b�Al�TP·m44����%�����k�������̤�F=�/�d��$ʡ��C�{�f���l� ص�R�K�--��t)D�b|Eҁ�	��t供�e�xw-�̶~�ѷY.�X%7(s�_���*U���%�
�"�e��*����]1f8�gm&#1��8-�m৆�}��%QQ����_UW�^@�v��+�k�/?��q�/M��1�<P��>MF1�{~�������n��Z���6������$I!�WK���y q��eq��T�4ĥk���w[�`�a�n�\��z	USf���-�2yy�6��Ɠk�\_zs�n1J^�-�|�H��)�sjND�qh��#�:��oM|�1j�ŕ�����wT�����f<��q�K�J��\'�r����z�6)�n핐M������&):Oܢ���%�ASe���*��_H̶d,.i��VZ�0�<�b��Mw9K�~��F���ӄx.}�}�5E�'<���tfj�956��TUk�������EB���zJtD�c�Y�s��xK��y�dewN�$;9���F�޸2�:��7��F��{�4/^P�K<����p�bgA�_y3������f�u�Off�6�t���r��r_��̷.�����w�)8�eYav@�VbXs��4�����f��O5��^�Ţ��I������\_,�Kh���)��2"�v2�>>>�o������.���	�64^�;hl�������S� �����Q�����x���&�\�}�j�է��5}�B{�L�f���iж�M�]:�ڻY�g,��+ 4�&fX��؅̔�=��m��t&v�Ge�q5���b���/�����5�][.�f���݄��%jVmm�S��bK>O��[�TG:��ґЬ��xfqz�������\l���93l�^rk/�&�� �s:k'm͓q驩}�ŮD������;���>�Ҽ��t+� ��fQ=[+rc�2��w-�zm=�n�t\f`�uQ�����������u��bMbj��R��U�,�*R�w|s	\ �Tm�:d�FYB�q�[}��r!�t����l9����Pl�It�{�[+����RX�X�xAZ�4	(K��)φϹg;�aN嫈�AZ6���5�7���������l����,R_w6������Kx�|:�t.�p�:3�d�%�Dm��TSf:b���d5��'˟r����WxoR(����DVs��ۜ�-a,.�:D�)�|���4^��ux�-Ϻ�� �|��֭A��#��R=]�<�r�."��G%�ɷt�d�p<�e��X��N��0Y����\�t�9�����k.�&�t�?$d��-��{�E����9a8jTb��cE��N&e�u�o[n����*7v�r�V������݉]�#Y��M��6ѮrHQ�Dk�t��Kko�{��wkZ*K��e��)���{�׾s=wЖ��@ӽn�8օ�p>2Q�&�5���i�ZRMc'���ʊj��������W	���.�f��4�FK��'Ti�p˗�#�+s������M;��&#BZ����C���ݼ+�I�V��zL[J�uf=��
W�����sa�����1�iI|n�f����b�/'4ȾHZ�N�ˠGn��*�W�$�ͨ;r;��k�3.j�IԒ�r��P��f"�_��	�
�,�:������{�9�
�x2�c܎
D��C+^����QF�v��r��M��'%;:��	�&��@r���@^57��q]aayF�G �`�8��}V�L�5@����U��:i�v�V�J�e�x�6|D�֏cQ����GK��r�ۑ��d����m�è�qέ�*Wc(J���a�h��p}2�|�瀻<�����-��p݊y�a2[p���X/T�|m�D�9f`l)�"T����̚��مw��n\\K�/���$*�Y	�ɑ��I�N�39�������SxA�*,J�_wZs�T��F���/����s�'�`�2l:$dV�%�Wj67K�gpo u��ܩA�2Ҩ&�������ע�F��n���dE��m�^	oT���d�Ze�'�5���ʝ��yf�>4H�j�5��b��0,Z�nG��cy�Xz&��RpI���t�zc�őR^>=�Ʉw5�����Ri�z&�1��]ٱ�sg�N}'Ұ�JkTNҌ�F
��*ꥶ��dGn���m����S���ҧ,�o��EY;[X���J�J^^
��͍[^�G7m�8Ŗ�m�(�kUJ�J������
���)kkV�6��F��ڭ*���j����[*U��7���Z�6�R�.nsN9�Xq6[yLkee-9KǑc5FVډU���[j2�ң������(�D<���4Z���歴��mP��UD���J���-檷���*6�R�%���S6�;z��Z[[J�6��*
ݫ��^Z�J�ZR�J�Dn�jmQU�
��DB�����[NYU�֙����q�ED]VԶ�[m�]��`�>������-�w�\ܫB�)m�o�Ab�ET�6��4k-jjF[%�DTDD�]�e����]k�ڋ�5kZږʕ*�:����U�DB�j��u��U)�Q4{k5����F�^Z��u����~N܇�.���5��o�}\��R�Jђ�mmjFfukk����	e]+[�:w*��/X�&<����ԭ��&��xxFɍ����p��/6�|�OI��xл%Ra��y�=z�Ϟ���h;l�ʩD32};=.੻�ޒ�L��k�2[�'�4�+5i�Ck]�Y�3ڶ/�Ԍ�n#��R���o�'}A�Jiu�g��Y} �.Q��SE?��H�����vϴ�T'W�[��x�w����+q��oF�/:Ȟyũ��Ҿ(G�G v����z�%;#s'�7�ǖn��ّP�E��{��X��FA����:ܗ�F(J�~LE�P�9���㜵ׯ#����U.+���;���լ�����S�_���K*ly.����{`x/
�"�^>���~��$F��z��ql��[�j�� ���G��3W�!�=�I3��-��o��3��Қ��1*��^�%"�#��m�p��VT�
�ꕯxaP��)>��yU$��h֙W5}��c������]<��\�)��y(�rq>>27Zc�cR~�2*x+U�l�Տ7$m��Rו,��4{$���1F~��P�-%���ұ�i:W���Y3\�*g}(�]�ʕ1޽��p�I����ndo9ۻ�wq��n�nSc��:�ر�P=S=v���NO��纉�boe���\�u��`�5��\�#�pp��]��9��͌��b��4^�n��=��Rz^㳌=��P��)e�_v�ر׽���=��d��a�ڿ�|�r�"l-��>�n�k��Y��I��t�}�p�tr�.�h'ێu��OO��^)�)�Y��d'�Q��-:L��?H*}��}�~�ꇀ���Mр�����L��7�:�����V^.��@���'vc��=�g,�9ßR��iB�8��2�;�c��]K�=��'g&㺦�y�5D��a��(��Q��t��g�Oc^*���b���K�]��R(��P�̫�b�Tɔ��=�;8ػ�C�����A/�*�s�*�;GT�"u�iMtB�}�qB���yE��w�v��lt����Ē�u˾�BZO�]��cc5	�x�/r�g�MSsP*-�9$�	�i��
�">aY�H�������J�=[f:�P5���}Siō.����jcf4�["�&�G�EBvp��կ�Z�o**��C�fc�q:֚�W�	�wq��<���08��$���}.�pU�����w�fs�t��ם��u4w�B�aԋ����Oznc�n���;��Х�p(aSlQ�gO���6s�22Ֆ����TIR�rY��Pʼ�|k�L�˫�oe����2�;�1��t�})*��llE�����E�N�h͸,��4�ú�j���8�0=����Y�{	ʓ����kc�T� t	�kh�D�]G�t�6��͗&�`���rg�C���΍=�Zm�|~�DKh���|&ME������̶5Y�L��'A�Qi^-��M>~]���(�X2��8u��J#F���Q�+�x�Ξ�L!�`_���w+�-��sh���	rW2vs+b�߫C�wWﶍ)}�7��)�}3mC��x=рc�s��P�V(�a.b{�.;�z�3w��C5q,r�e&���H�w��yR]�R�D��Uy*mڻ�6ͻ3��4�U�n<a��k��E�x�&�%Tǜ�]6�K.��9SqLxN��Vc��텑)�G��м3�qvDLe�C�d���b�*`���� ��I�c/(k���<�î(���xI�-ف��t�`zrE1�+S3c��l��#�9Y�|��q[�s���+��l=����n�eY�X�T|��y�A���Vg��<��WC?N�|J�O��yLW<�8#R�3p�}S���d�7��ŧTm�Wb0��K��6n�t��W%xv4w����{��3"k�7k��������r�u�sd&,���5@/;gL���毫{���� _WCW^:މbbRY\f�1����X�Cep��3�w3D�%LX�t3.|��Ag`4l�F^� /E�N��!�k�
�k6�Qh+�v6-a�HRn��/l��cp:�:ݬO�8Vs�r�3m�����<<����ꪳ�G���F��y*-غKEе^�y��j:=��Ŗl7�im��o�PF%��޾��^p��#Ǽea�/�:�9s�UGv>�+ی*����nz
XtkrĹ��]1�IL+���|�|Vh��W��/]���Z4�R1�|0����"ď)�O��Oz��*�%���w��c9@ga����2i���0#j4Ȅ+y��y��BhnH�;u��=!6�'��� T�vˬ��x@�Y�����(J�(ԕ�y���=�F1�ݯsH�ڨ`���U�
�o'L."r{��/j�k�e�[H]o ��^<9�*��qT�x�d���H�h�}�cQH
�C�g�����{u�N>�'���>��DW?6��^՞��yT���%ɺ����sfR�Syꮮ��9�e�d�j%�i+*�xw���κi�dJ9�h�����3�R���w�T6&;)��1\�َ`����x8伧Z��)9��)��
�ǻ��k�O����~�w������y���U�L�sF�S�z+c9ϵ[9k�O,���|�j�!ܬ0���S�����H�"�ߙ����,2h�]z�j����O���d|OJ���V:;�wV���+�34tm,7�ԁ�Owsu�7mR��􂶱aK��N�7yD��	��g���WX�����c�;F���0,W4/W�;�]N���� x ,^�1��n+����U�-^&�1ο�C=��4�@��kً�Y�i�gi�y]1,D�WgSҧL2w�����&u�/q�K��@����ޖ��O�L-y3��lE&$�d�����\���퓲�3}��]@��;_�x��vԳ��I0U�d�1���
��)���d�`��-�R%>��m�8�r�4����[�g�BU�ش���.����;�'�^cB�1�����#����r�P`U����*��-�hOB�Ϟ�q��v���b8Y�������1#����kJ�PX�0�1�c�y<hu��H���2)�]ACh:1�s1�wOS�N<�tTx�F"�4ʼH�Uѥ�Է)�ZOr��A,�Lt�ΘU<r_"�x]mĮ�\���#d5�c����\��q]�ߞs#a�n{%��9��Lz��;e�\[��d�~ħv�1����xl?�F�K,��yV�o���ut�.bl�7>�g�',:�J������w>gسJ;�Jw�1��e@�#����,��7��~�e5K�ǁ��/x�)�]Y�w=b�����'��%�����ځ����hOwY�v)�dYf�OStW%e��f��cX�cR�$�c�*�0	x�v����zwqb���3���o;y�50��;iI��>�����=�ŕR*�/q��S|s����f�feIB��������B�*v�+��x��7{�*�E��́2߻ύמҁ51�+۪V�� ���|�VP��#b�h\v8.�Cd����m�1��g�
��g���9�)�vr�8�G�n�=�WZ��?<T!���[)q{\r����b����H�'��/Ş��-%���:p�'�j)ժ=���^�SL��W˙>̤��yw,�V�,����+e��KfCd��M�e��ٛkР-��]XF�Hl����s�Dr��2��*}��ݍ�3q��^y��s>�-S7d�ʗ�8���/�f-t.�H��+�[<F�>;�B�=��0��}HX|�bԖo#}�-�u1u%����&��/��[��܊�OM�2㮔�&(�d���&�d;��|��ϫq�jex��(��ɺ5�
��k�T�$���ݜdNqT���;�	�6����ʝ����R�9�N��,S���1a���Z�x��|�^Yg�z�2�䔿G^eVP.�9�����o)����lXm�|6��Q�<��*@�/����pX����E�Q�����0�X�*]�����?Zu��#��S�$�w���?N�����*)ngD��*kGnR\e]]�\]_A�6�h�2�|�R�[�E�Bj� Z��b�o������|�D\�������7�RJ���8do?˾��A�(Gy�_xG�Vk."�2|	�*lOe�(����vW��Nۢ/u镛i��6#I��`��O�`7{V�[�T�z&��1�n
��yfc��F���]���pζ6��|u�ҧ��<L}�3�@[�)*ϮtR7S�wFՋ�ૺ�u�D|Eq���>�(����&�*>��0	���_�����3��:�3�,��}x#�̬]�լ���O��|J	����wO1�I�hj�	�0�
�v-�t�Qv��A�̆R�5����=(��h�O�������l���-�:o��ƌO�v������a�Ͼ	��/)�;�f�DҾ�b,uԦ��F^>'9��C$�O1�"�5�';�:���dd��e�Uc"�P���KAmQ����W�����5J�JOR�ӎ^n_B8:F��|����!��^F�9`��Lw<US"�tSg,��=\��x�I�YI�:��e���+��/h�!%�(LǞ��h�=A�9R/nbS�
�M'�f�?,�0|U���
Cc�
Z��P�^fIQ����K{x�]
�9�;��=�^<���RJ�l<G�պ��Ǎ�}v��r����n+��4ӳ�st�0G����Z"]�}��ne��q2�d�ѽRs��u3���q�o��.��ڜ�m��c��������EFtH���/�}��/�W�U_}�s�''�ɿ��_SO��-�1K��	�	���Gay#���q~4���QI��4�(L�c�ŷ�a>UjƤ��9i��}X��+��o��5�Y?S��Q����$@/q��&wf)Sj#ko����%��Le��~*�洒[+��	�����#Y�7�~�N�콩�^���w�2��HW!Er�n[�$�.k�9:�9���Z̀�y��Q�ӌ��+Fti���Ke피�i7���<����@�����6g���GoY�l�՛�)���	�o}���o��#�~;H�Tɔ�˘�W�>w�C�����}�����r�Y���#2f��1��)�٤վ">kk���s�Yh�ݾ��ˢ��T��%;�"�7hƕ��9Ք���*��\��G��_W�S������!��V�������%��>��uTB��g�>�,x]��}��|�%d�hbf����"%�7cv�\��ʍV��g��Z�+�x�'g��U�v�	�h#.��|QǠ��t���R�t�p%���_�r��+m�~��XW�/�0���ݑSak4�\�YJ|&��ks;y[H@�62�jt��J:6	w�^�M��Sw�V�]�y��ʃ���t��s; Rn���﮻0 ]_1V�sKҎ�C��d��+8�`�wIX�pq�n)�s���m��o�g�7��z"q����'��x�|;�v���R�⊔ͯ^*�/ڲ���\DO=;�z��«b����(�b� ��B^�K���*�+�+^��2j���M�
ʦ�K+Z�T�<5���[��icuO-[y�s�/W������4t$^Z�~�c�N=��s����G�[p��5��'��u?'��C�I��'l�,��>�)xȍ�F��W
ׄ@Y�ځ��ԍ���"�dW��ct덜�=x�P2+$�[c�.q�6���`��Ldu��/�� ��� �Y^�����v�/�ϕ|��}���u�i��H%ի��jD2�ނ�!�	�)���k}:�aj_��j�Kgv8a��Cm<�Y1m���X�ٜ���v�����$�,dY��`��h�؈�s��N.��!��=�Cp�2e��M)�0Ybg���/�ݷU��U&��,<rYۺ��kC �	��0��At_v�����*�[ܞ�l���s+�d�K,3��[�Ѽ���F�CtK�ܴ����4��df���18�#C��2[	��%��r�NV����'��ҙ����\�kyڟo���6o\=L���X�ڼ��u�p|����mV'��M��t��wId���;�����8�s��l�AZ����훫��θܐ��s,�0��$�_,��b����`�օ%"}iی�M��w����c�=� ��o<d��q(��&lR_P���P� 9|�K��!ֹ��r�[:5N쪞^���>��!���+|�k�+��BuȀ��%{!0m?�0���L;�}���/��}x��uM3˃U�ll@�O�'<u֥9�������:ܗ�J���/�Dn`LsRdݞ����~6�
X/D�5��M؏�n�3��}ˉ���%��/�;'ӗ�Mؙ�]�.��ϯf�l�~ܥө��n)R�Խc�j�[A"f�� �'!�B2%���m��-���f�T��J�Ǝi}��iY�M�pq�Ed�	��X���1��QE�(��ߺ�@��C^���8V�ꓺ�{�BjKGrAtc��б�S<���*v��鱜Z��D���
c*���ם���E���ޛ.pmȭ��aqv#Vy��I�]��Q�x���NeL��hu�Y�9�~�
�Ͼd�D}<�L����!m�Ǡ����}�>��i|���R�(�k��~�\�
'�A�@t�/p�f�0���EՂ�Lu�>�f�n��Y�sϏ���=^�o���F��~wa��I{QvKo\O�A�0��+DX�X��z�{�W�Ӓl�gd}p�K49���}k54�ngU�d`rJL.2�����򲻱����\��[޻�����v�F�2���pY�,�m�*ʽ����M�o,�V�a��v���6VSZ���tj�U.[u�ae�)u;8�4MSS��n���7J<���t���o] ��uӠ� ��)W�0q�y�p7��5��wsbY,��.U�/��pt�&�d�yr�:8�S�*�*�z�O/m�E�t����M
��#��`��L�����]�ǻ�?]�v��T֊�D���s�j[X��|h� I��� E���LW���ʌ�zlE+���4�纬X�k�X���m�B����nGS6�GC���A���b�R����e�9��}������ۉ�xqb{U�3��`�VV�rq��#ż���[�� i����a��W�-�k3��tq��U�J	[�r�E�vJñ��06`�u3�.���2q����|%�*���d`u�����T����v#���^��]L�Ò�*�*We��!ҷ��T��(�Je՛{Ω�mAR��!n��<�"��,ݥ���=b�s�Z+,W>�Հ��z��܁.R˛YD��Jҷ�M��ft�:�^Pk�[�&���弰_��=�ʡc�FX�N�Ec#L�\�c����z��>V�Ƀ������)ֳC%��[7RH�}�������+a�zPx&_ ��0rW��ԊAp��7��{�n�T2i������۹��I���&3^+;���hj��	�%���2��P��Mfi)��k�+�$_&�%˻[��u���^-M��N��d���_-�1�|�q�Y͵rgr��6V�E4���%,� +d���Z6��P��.,�[O{A}��YN��[��k���3 ����E7�JDs�j��d��e�ng^m�q�U��1���Io%G]���mt"*u����[!��lp�4���\��ՙS(p���5�gc	r�J;��*��!��{Q�Zhec��;H�~��N� QZ;wY�\T�ݦ���ٻ4��x�;�֦e��]�JM�Y[e�.Jxa�(L�M�^+܁n��-�����V�w�"Suv��]1� ;\+9�l�i҄��8�p��nʉ�j�Q��Ń�3���E�H.�9r��0�1�5�F���s�,^��wk2�-�Qa꒕X�-[����Zp���#0��UEy�Q�H�l�n��ݍٰ�X��Y3��r8�[%��w@{�յqq9�r��w���5�E��N�	�z�V��W$Vb�����R�~
�DZ��K��1N�qvh�<��5�ٳ�L!^ˎ��w�'»�u�֙��ң)�S�cX�Wq�J�-�ޑ"�\;��}]ֶH�f����8�sz�4�&�q�����xZQh���S%-����R�QEQ�.K�8������D�Q5)��F�}܆0X�PS�#jQ^R�h�O)�ߤ��)PTMj���[b�6)X���w�3��j%����*��ŊGsh��
��p�6լ�m���VT�`��	[U��ATU���*f��ra����l�Z�H�DR�X�hӎa֨��<��{��QX�ť��Nڨ��k�6��*2�䨜J/�[ZV��n������5��F�X�X��"'Z���D8�Z��Յ�JW��bыjUu9��YA�mhբ�c*���[UEm�:F��*ł"��Q��`���}6EA*���Y��L�D�AUb/��[N�z�:�J�h��1z�[KR�(�5G�T�4�h�EETgmUV �Tw.�U��U�i���[J�KF)�P`Z���^���r�u*)����jU�J��u�Dyk�2Q��d���U��\�+B�R��;�[�{�ӑ>�P��Z�}�ű�i= �
��B¥��=#N�"ˀb��T1���oj	��p��ks�K:��c�'_"�����ZEG^˟��C�g�^��7'��)�v���6�t�9�ǰ?O7QR��L�GAQ,Z�jYͽQ9��u����&���	���㚠R�Q���ثge�xF��7��;���� `�ݱo*/�Df�%i��PN�$��;9	Z���w-���Vo���oO4/��8��n�R�'+��临T�qC����9�XF���5O�)}qA�Fg'���1���W��[�o/ת��858潊K>P�T��T[>S���
�$�a;�|a�Y;:�T�n�19��Z��]�lYY�E�J*���t|�6p�S�lƙ�l�Gdc޻�k����c4�d�T��H�!NI�"�dG޲��_FHez�ZT��`oL񕾂�uN��,�#ʫ*�&o�N��O7��l\rQ���2�eC�&v/n������.1yP#)�Fb�ooj����Z���d���zD�y���V۫�gg3&K>�ǚ�(�t��@{h��i��[�ƚ�CZ�y��=�hWsDg��Lc��G���������~t���`�9:�����!7�bY:�X��]2�ލEvl�	�J+|!�FS<N�G�v��Dwf����H���<��ɔ�*ʚ�g+S�]s;.4#X��S��j�/u�k��ܗ����j;��^ԋ�v�|.X�tv=c�_}��U}:dJ���?�By���PM�H�z��U�O%�8 �b�y�"��:��rov����ȼ��Ƭ �mm{��4�J�/آYj�����W��]R�����;��u>����;����c�.u�(d�.��WXQ3)��UL��]6ڲ���s�았{W6bv�F8�Y��X���B5>��>k��v��yZ���R��
�m��X����w-�)���4���8�
F!�0[�[�/�yLqyZ�(��E�RS�1�͕s�8&�%���M�����}���|9��9�e@V��Rl6�Y����N����C�28{t�A�7�������B��E�D��u#��/��b)�b�������љ�5�l�d��:�ۛ����v*-mc��`����|�y���\�4�݇ЎN�NlłsO}�Mcp�
w�^���0��+�(冡A����[x��O�~&`f�ّ�}�� �ث��~Xэ�(��e���Y�UA纙:�UҞW9R5�tt�}�L�������^54=ZK�WD{��Ŝ��W�s���A䧽Lp�Ƕ�v�eN�
)���H��|�mJYLՋ���C'kn�-]1_��V�h登�2��7�M�`�����e0��r���νO��n�R\���5��`�v�ѝ6�ප�6og�������������Q���553���i0�=�{��������C��懶�<C�>Ϣ�<�	��0+�az�-�[;���1g�[�)�(=4LAO��N�5c��W�D͙
߁DZH֔O����|#�4�![��4os����#u5�ɻnB�i�5�/'y;b��[<6�P����z_)�+$�@�5

z��c�3\j��0C���v���VB�}�^��,���f�P�l�e����gz_)��}?&"�*bOa3�7U�t�s˸��W�۩��]��z�w�-C'�`�c�Q6�VK����""���x.EZ���x2��3E��d]:�aM0�ʐ��MH8;�is���2i�ɲ��M�VV��m���r��p��y�o�=�M�:&ſ�m��k�HɊ�<�f�5��8��sω�>�r���:�|���v�"߲P�w�Q�,�wG�x��(�+tz$\|��/���O~Ό!�B.:̱u����n���ʾGr�NNlgdKm�7&^�ǲ�>0�)��H��]����׶?>|�m��u��5ͶF�|/m;; �\��*,:�O��*�.�\��J�ƽ��2hDc��\��7���g߆��A���p�[:`�Ar���}���ּ���k<p���w�0j�@r��Q�W�@�̚ �b�F�ގx���%"��9>y�%��W#�Y��+9�:�ŀ�Qۤ�A×�3U�|z̋jt���7�?���� ӽ^����}!��׆->�Ǘn�S,MB�3��}���F��r��x=7:L��7;�g�jDor�5�ݲ��P����ؠKga�/@��iOe,������*��;fS�˂#�L�$�%@�V����]�eM�Ƚ�v8�L6����kg�~���RT������_����D3tOH�v��0P���X����e�2.D�����\AmAt�ٓU�^�!�RvŤM0U�F�禾�Է-�}��ڵ�����v��>��t+W�u(����y	�Cť�zP4�s����A�%�T^%�MA��7�����_t|��Ȥ��,֌�����u�/��P��x���kt�%kH��36�:���!z.4����^��҇j�io��f���3��rw�ǯ�����;��5�K�Yp="*7UCƫ�ׄn��{�:��(!�dKa�כ��kBm�w�^N`��5ͮ��L�D�o.������7	��ǚʛa@n�Z�Z�hS�J�w�KIw7J�5T���%��� ���x���i�L-q���b|TbY��-�nV�NRΗ�Տ�V����^��׃X�ʹ��Q�����9����uGowB\�Yb4;^H3yl��-;�]![�%6t z�jJYr���(.�6�J�LC��7�y����d�	bA �e}��᝷�족� ���&���x��[��� ���񛱡Ϫe�=|Dܯ��V#nj��4KK.�M��^S�ˑXAMY�.ƪ�D}�h�H/����Q��-�U^gћ"ռa[ݵ�ʙ��b�&�[��ϸ��kl^=��6�9eF�{]Ĵ�d���4_<5�K<j4�V=�/.�����F�]ʕ?C�觊e��G���v6����T��-bM9����PՎΨ�Z{T��sҎQ�����"wf8�|uR����v�����r��{˚��e��ҏ�9�?&��ONO��׼y���(��:��)�e��t֚�Mx��ԛ�X-Tv�,�#m)*�j�]�c4��c�u1�Z�bәvxvq�quX��.B���Vr��Fl/ND]v�+�:_/r�Cٽ�H�>��u�a�a����x�W�}��я󩙐c�}3�i֬�%�y���^PM���:UKso)/�� ��6Z��'�c��2���L���W�*ۘ��\5 �f��LcX�y�}&��y�	v43���7�у)渔�PR��� �������5��.���]n����n�%���/b�<�[��v��{1����_-��x2�ٽf,\��n^0�ё�.��/�Q.���T �of���ܛD��,�s��:�m�g*�Q���0C|<=� �w7��'k�����v/�&���`�[4����Lf����M��(�~j�c���
�qK8k��\���k�7��
���W�b.��xj�KT�ρ�^�1�g2<jC��c(_Qg|��¶<A���X�ᶺŹ)�OH~���W���E��$����Ψ��/v�T�-��1�� ����:]6׸����1.�����B����lJX���q�ZX-%�%�m�i����E�ݩmUSk^$%4Z��4��X��ER܅W��A�6_��V%J���':���Y���P�g�q� ����i�X��T�sx�������,]�ʈy��;�{�B]�i��M����ϯ��2wˀ�؍H�4z�mq�%�2��Tȹ��m��ˬ`�~�=&fړJ�Vi㯞��\�B��eٝ)���ؼt{wd):x���NXYU)��E;uK�:U3{�n'��w���ڇ�Ao�o4l���1���<�E�Ժh�/��:�y��ސ�+;uw����ׇ$wGR���5�q�W�_�+3���&t���N@��W��ưvh}w6�:8Ο�$����]�����r�_C���a\\e��]�������
���g�V3�\zV͝w�F����=��Khi�,�(�,`�۝�j;��["���{�f�{���!�\�n����;W��i�z�Iƻ��}1�DsG�������gm����D���ݿ���%�G�y%\��9���B_H�^�V(�$)Wb��6���{�Y�2����ڜ=w�2��K#�T��
8ܶ1NIj\ބr~�	̀��V��g�t���.u����u�*��r�J0./'��3�9e���~�O��ٛ9�Z;;~�L�/=��7���+8��3͉,{APKץ۟�Ǥ���9��е��3�l����[��ݽlU�1S���+�����l�`�� 5��O�9֬�mn�R7�1g�vp1j���(V�U��p��'"�:�
"@�Ѭ�ɦy�fuF�B��U�3��q�8���2c�.١��=��J7�8�ic}����ʆ(J�(��W�2�o)��=���a?��+o�P�a��7�q��͔_s�j�a�vy@Q��|�cӾ�x��ܛA����wUom��E���QQ��*�ۗ�6ò��'d��R���W4�z����Qq�|�r&q���nn�Z�ס�C�t#$S��S�e]���a�5Q,�l�M���b�����K�t��x�b�Z�C��E���ru�#�PS�"T������W�\�v�4�XjK��NN�'QY�pmm�I�MC�������!j�g��hN{'rX.���JSU��.;8IS6gЄvh�&�O�3�o�d�1����{F�}JК�T��NC�H�c'��=��ml�}T��27
�+�'\�[�,Jޔ�K΅��09:����{^�"�hq�Ƕ�VN��l=:��/N��%)f�����9���cnr(���B�2H�!�^��\6A��K�~亅��O��#w�P�m�^�S� =�C�yX\&�d��)M�R͘���̯4����E'��@���(uʺ���_|pF�����/�*[1e���n�\���&l��N�Fla�u�}���j����^g�I'(��7y^����/L��u{ c+qT(ś<U�e*�8���6��Ҟ�,����{ɲ'��b�x�_�v;��)�ΒG���3��1���^y�{�=s�Nq���L2�k:~�:��������?ڣ�dG?��U9��g��>R�3�V 4�`���	q�b��<���ٓ�F]����w�;q�sk�Hϓc��}�J����_-$4�4�*�#
�4Ȁ���o*j�+2�ll�63u^��r7W�<�\�U)pގ"�8�5@oW�BOt\I�2>�5���b�2;܂j�y\��n�L��`k�v�a����m�ō���z�%6��[�>0r'�;��J�������׏��LM���I�UE��)3PQ.̕���T骥H��8�Q�� +FIZ���QD�V`8>4�s#o)�M�ǭ���    ��m3'Y���=������^�L�Y�u֥9�����G��_)�+ۼ��DD1ꌛ�z.WP��{��5z�?�'�(��4�ܴ�V;K�03�-%�;���r�z��F�ӧs}M�K3�#�x�a�QC��S�P!U!���m�c�UC՘A�= T ��o2JM�n}�y݅w���w��;��2l�iG�hDY�M���k*m�n�[q��w���d��j؊�-u�U��\c�W��V;f��?�Bj>�h�F��/R�<��r�h�F��g\l�#n�1BJlk�	�=�QI��]�3�7�*k�Y=M�/��{�[Ņe<r��5Kw�=[��`׿M_ ����?N���8U��V��w�6�,��������	�	i����.�ʲ�d�=	t��HA���C4��(���E��6ȹУ��o��7�hwX�f����J���� V��)Q�\s:b�J9@ʽrє�I�M��9�\�]������)4NwaŊ���g�$<k0�ͩ7G&�q�R)F,�LEel�/��9,\ml`3m�:/�b_1�&��Y�����^=�^���2�
���x����Z.��QlL��b�?`��S�-z���9W�%�c�?�j�^�6��c�orl�0=Oy�}�Cظݞn�>+7Eqk����
�K�%��%��
{�x�����4�g��C�y�����r�*�͉	�~E�ڔ�K������k���b���99"��DC�[r��57p�Pr����ۺ���Bм�fvoO'�_<�+��Z��B�:�9�XA,.w����i�j"y���Q�v�M�=;V��E1��,/̀yX��&2�ϕ2p�s�\�Q6`�ٚC4D	OMOm����#aA�	�Bl7�LN�ON�Z�Нק�60�V6f4�[��NI+ݸb��2����ܤO�+�>���?B<����G2�0�+B�b���ٯo/���{f��sX��u�S��:�)\�n
��}~5��Bbj7�^5�`�|�ی�Mj�سz��(U��+ً��x
�D���x�R2����OH�����~�?}wц�Tk��?^�阤o��ܸ���7J9+M5ٯA����}�4�Pw���	����ލؙڎo?s>�};t�PMn�*���5Mm�(Ah�R�WB��ڱ�I��Q���a�Yҽ�7���Q�\)�A�I^�b�'�>A'�����AN�g*�Gͷ�*4+#\C� ޯo����+޻�V.��~�
,��rfS��]0�
��մ9%S8U]ؘ�7�4�d<YPZ'u��tX��XC]iƊ��1�Y�[��,�:�[u�v�]������1;d�c��Jfr��a�Ÿ(�7;8ò4*퍘��N�ڶ�gvu�u�j�Oi͘Dֶ+��L�ڏW�%����J4�R�/7&7qphc^\�4��Ie
�L��& z�s6j �V½�5o>ӆ]�B�\��L2�N��ӂ�d�:kr�*��,sN�׎NMm.MGX[1Q3]k���Vdヱ�ԕf��X����$Kr���W[ʶg٢�[�Ջ{1��S�ˍ���RT���p�3� � 5��MژҼ�2c�`�2�L&z�-�q��_u���,�b������V��{�3�=�N�zn��6I��1�V"�c������BX.���.G��d�eY�8�lb��qec4��Y�VZ�\���Z��HሞT�-UTcx���ڒ��W��j�R�	�Wu��[�I��[&�"�x�9�Oe���3�T�-���8�Ư��5施'i��h:�V�j�Y���������3���v��mn���ԥg%�3�N<ݑ&�*:��r�{���c�u�y����=�C6����D�)�1oU�ھ��ưm�뺺<jb��ed���IۼSv�4%�u��z�K�vz�j��F�h靎�J�U2eB��e`��<c��G�0W!�k0'oca��y���{��ht��<O'X�A�Xu�����VԷ�@f�ĳ�[���ш����x�P��tl�ER��}R�wӻ%ed�ޚ"/oe�Ն#.�J��5�ȸ�o�ݫ��,Xvr�u�1���R�:-+�{Wr���C�4>q�u�S���ec:eK�س�0_�;+q���Y[���[h1BR�ke_٠|���x�-Yt�����Y�^�QV4Z�+G�������,F�Ԃa���D�Ҩ�cp�w#ckm� ��j�����9.��v���@t�25)���%�!��
���1����x(�T���N�@�x^����2����|��C�G��3o42�!�u�X[>�R�K"�.X/�QV�Z�C'*�d΀ޅ;F1Z;n��"�14���)�k3�`gk7�!��ǥ.��8���|�����Vh��x�`��]��v8k���}k�p춦1�3mu37R��ʶ���"�J�*=/8�:�!�l �ظ��ū�>)����(F���Z1�r���n갎���-�ũRgO;s��������9�^$���;��բܸ��.̆&f��s�[����[�Rܚ��pS%�N��Uw��}D�,t}�7�Y(r�:��J�Й����l�Ab.V�X�	`9�=Ė��M|���
��o�Eb�K�v��XuN�з7T���뜹��m\�P^�C�=�L��L��V"b��D*'q(�M���g�^�u�9��7sS��K�cn.nH�$�>t�u7�m�#S��˵sAs*������J�%J9S",����1�̪���]�����1����\��;��M<�AymJ+'��#Z����,gR��v�Qm�����A֋iDz���V�[Ơ�1�)�W幔D�.h�V(��[mE��h6�֪ƷoZNb�)Z0V�m�ٶPX�����0��6�A�jy��ĵ����QDwm�
���UVM�\*V���m�w�A��ANlc5TA3�Xq�U9IE�4kV�l�^�H�#֨��y�&b���!뗌����j�=��ol�V��#iDԺ��=��"f�m罧����5��{�"�}5Դ��`KV��T����ܹWZ�򙋘�l9ku0"������*���b+�+PQ���6�)��j��f=m��j�v�DX�V�s��*#�Tj68W��yyR�E��kTR��ڊ��.�j��sC�ޞ �i</7%)H�@��:��*�4Vt�(���*Z�V�Y�m����u���zq�fΏ�{�]��6�f#ԧ++;%�Q��Z{nnof ��oc��D	;\?߾�ꯥ�ŏV^��~(�?�%C����	~,�C ���l�X��x��E�.�m�4z�j���-f��)�As�C�k�ͫ4z����b�����c"��9a]tz��TB�}=�-Ȇ%�_���|��ɞ�	 ¿���{Ѝ0>9Hq������N;\S�Ù�.����գ�yR�ߟȀ畟^�7;�԰�CYV19 ���o�����8�Х�����]������W��*4�Qϧ��z���~/|�!}�tk�k�Q��4-�Ϊ�au���s,��l��L�
Ga���o�`��L[�?o<9�뢣Oa��^�Nhʠ�����j*����	�0����j��6m�D���(vF�R=��3V�Rc{8-	��b��#����2G���s	�}�b�R)O(������>�g�Sv
oW*�W[�V�=�LO�r�\k6�>l�����bDu�-[��>��85^���2���e**94lA�76�c�����Q�c~��?-~i#YA2i�K1���,�4��[~N{E�uǙ�f�ͬ�}W����u���w�5J��k�A�Y(C��~��l5x��շWV_*ڏxv�xB5�r�Xr��U&:��-?�b�V�^��W�+�b�.T�kk99��t�R���_��l��s�#Ur�B�g<3q���;g�WOw�O�?ϫ� ����6�['�>?�U����S1��q��č�<�ݏK�?b���	3Q�g�xdZ��5�WJx����t.�q�pe�?q���hf^�.����^"N�y@P1]B~iw�u�9��x�M5�.��\g�{v��"��yUnMcs�W�YR���t�8�����Ј��w����30�+[o��)U�j�@W�=!�	=^�`oV�P7=��� ŨZ�d�����V��V�f����'�{�7�B��uD�G��7jס#0��?k�+�ɤA�	+��Q��K�t�No�dSm�-Q�������I,�)xȍ�F�0�q���<���_�My�60g�L퐪1Q�d��)�9�P������s���ޚ�Q�{�>�Ȋ��M�K�N�W����
�a=��E��:qk����)�s��@��欐i\�c^m���a��"���a�-_)���/	x<�.��xd�6󢝳�[P��e�a���R;pv���[�m�.�ٓ�^�>�4����
�<4'�EH�y�E5v2�r�r�׾\~�P��%5Y��s�1�����2y�5���; .Jĳ�9r�o�Q�oDͲ��
},弧GyOz�b���z'���n�+gYYƛ��T��͈-(}�1.-�h_i㝔��[�����{R��%�r�ժո�۬)�fq�;���¿�W�_}$~+H�������wU����b44��������z�2*��V�uEcB4.�#(=����&Qn.�)��xq�摶׊�0#k!�%�o
���ZdC+b��I�kU�09��1Ll��}��-s���p�C߱�*����	�`p����W�UѦn��j}�⦲��~�`�=�3�V�f�c�;�Jw�H���O!#\�z��P���[7tĴJ��b.Cލ��dn�Ht��u�6��z|I�w�n��~1�4�������n�;�^3C�vW�ǵ%��:xF�o�E?ɫ���Jz+\BWu��C×j;K�{&��㸨���O��7ب\�Ep��F?�㏚�Q����)����-�%e��q���eϧ�:�L��z�WG�9���h3V�>���J7b���e:��4=��4���7"�6�ݰ�k�Z��M7F�9>�Z6�u��R}���m�X�ۗ���˩�'�o���	O��ճ8D��._������w]ӌj;f�catǞ�j)>���
��=�}^dMۣ�n��s�fo"ȱM��Oʯ^ᷦ]
�:B�><���wQ}%ҩjl[�FN�C�f;{�څ��-te�W�rN%�����튠t���4�>�1� �S�dr�WlJ�u6�%=����59��u�7��K�{z�nu�v�H��ﾪ�3���#Hxem����سX�kY5��,�!��S�M��3^�U���e�M�7"M)��v!dm$4��B��~܀C@�2���Q{s2���,���T�l�xm�({�}�c��&���pƧ���5?0���ؠ��/���PA�I�x���;:Y9t���W��gY�a�8����B_<-(V��%G\s1�5M(�\�OZ7ˆ�PΏ!�3�D+�ʴe�;j��FK%�g�H�k�Y�V�`$(�x;9%Xc篎���95}��2���K݉X���Z����еύ~*0���r���9��b�+$���\�#���y�ͺ1���E2���[�I�cs�D��)�=p�T������v��;�z!�Y����~���qr���zD�2}����u�W%�Δ�8�&u��<Ϗ&�Kb},�5�{B�8\�j�0��9p�	�Q�~��P�`8���9,��+1<;��0ƶ6��b��1��vW��n�6�;MX���W��_����8*��[5��*p��5�S��?8�f�xolV�<=� [��4�?&	-��|�����.����yo�H�8���q��4�J�L�띡��]�`VĶr��C޷������x9�U�I�����݌MK�I;r��Q�D=�W�6�C}���7Jc��7��]"�+6We;��w��ۜ�{���9[ӳ$��2��J��s�r{ޅԐ,9�%r�������ky����[n���n'8�~S�s�krt94��d�g��w=�v�]�悯���� d4v-��w���uOi����00qo
kwmc^R4�\�˪�W��T��0�)�����~%m����AnS����yzp�z�RUq�P��a3�^��򂀺}[�~-c�|���*Y9�3��u��omy+�G��p�T�&z�Ti��C���g��%��{�8�&6``�����̈�w�l؛�U�d�5tHȚ[����r֤��0�z�����\��ُ�����تփb� *|�S��9�iJ�M-��V�m���J���R[lq�l����S\��>h�i��lȌ�H�8�<_5+�>��U<+,n��R����QI��j�n�;��a��cYG��)��|��{��g ���t�g������SNv����9w�9{��]��Z��Eb��Lb��pF.:1e�$^�d)�]���� 6��Cf��gO������Z����ب�=�Ў�OtG������̐�-������8`��E��l/�b��L+�����=DǸ%vl�>�
\�M�ټ�r �N�;�^޾Ѡn+�G{z 6b��/�1Bk� E���G�e�Y�c��Xq�Q�X��Y���̗��V	��ľ {�du�T޴W��K8��y��>rcўw�t��ymigz��;���GAcuj�Ir�y�=3��Cz�5��j9��A�2Ѿ�Aé2l�j��SJyGc�Hw���ݒA��.�8mk�<~��U�®&'��e�4+)lͰy��WZ���K�R2ٵ�\h�~���9跌��\�o-u�H��9��Ak�(���F�Bd�奙�GTi��`��v��0h��{�c$�T�^4{���ɴ�]� �l��"Ą�Ӈ1S	�*����n��Xe�2��qU���V\���x��~���Y���(���]���q�=xԺx)�J%�f��.I��X�D�%{��j���1���R"_�麉�cR��zʖO�ͯ@��lŏal\�&`��յ����^��J��0c�rh# S,�>
ʺ�B�kaL�wq�d^�z�}�۩s��l\r����)�`y|�@;��~�Q5"��[ �hzv�c_,ɲ�tv)9os`�N&Ӝ�Su7�v��l�{6��֣�#ZY�;�?)ٜ��޻��fӿ�^�ӊ��8�@���3k=��I=��W�B�Ƕo*m��+�r��Ub�1���
X���{KőAW���z�T�`F�Q�Y0wV���N���T.�T�"v�13X{:�hA;�|�=���*��3->mخ���]5���m����0Oow?����+;I6i������d��2���zO�B����S���O¦|��b�G�[�?}���7�gi��yZrZ�
��A�ޟ���T`����*�,YC���[a���č��\d�A*C8�}�N��J<nq4s��2_bѫ��}ѱ�3��E�/��n��a�\���+H��@K�sЗ��lmЮz�[������g���I3��QL��S�f�r�����r/���^���H�7`����/R�΋�O>t�u:w�:�PcY���亂�v�^=*^Sŭ�=�����=��0#k C�`xT|t�!u�{U���͎)���L���4�ұ��P��Z���#�1�~�~��A�I>�_yݰ>��Ċ���X�0�����g�kǕ����&%<v;��h�4�P(L��.�f�t"�Ø�e�l�r��iw��E���)ý"�<�R�F��o"��V�v�c��G�CvP%;(�L���u-�\}��'tZEs����$���컷�+҇x�5S�ۯ��6�2��s���,���{�X��蔣�9L'�8�k�K1�/t�8N)�(̾\�1�:5��A����r�Sj��΢�4�`��a���SKQҲ�.�ow֩��dO�m]�oI��^�E܏4S�3!w����OK�°�(/��X�L���o��X1�e��8�̥��7NϚ�=����'H�,�ή~x����xz7U�;x�&�ֻ N��ވ�x<-Z���jE�y%��&|2Z��}����_�=�R]�N�����j^����mKܥk�(A�=QI�����ئ6���/�#�?PX1��?�lh��_�ƭ�{�}���|ɿ}�?������L&\��)?X[�/m*�qw�*H��mC�Ӽ����D�깚�m��q���r��U�Z�&�Xs2��x��&��ݯ�fP�Rݩ�]S�Oxzmk��f%w�iĄdQ��B�΃��7�!�o�R���.�<���f7���Lb|�]�ɜ���^	f��1o��
Ò�T|֞�"���R�Q�:�)���F]�K�
-k���,.��%���:wJ�y�HOGC-(��ڄ���>n�]HLi�y��&3x�)3��#uظC�*H7j���FK$�9��zg���D�����!�X[�o�q���g�|��Ji��G��r�z*e��O3��
�tV�#��+�A[w ���3��,υ�0��)e�ya3HS�r8s�lɒ��E�y*�V�շ�մ�[.��-�?�5/2f	���'f0'i�hǕ�#���Ӌ��H �ǵ!�+:��u�tR���	�EZ��sZ��"ˇ����ckL��Xcy1�Ԋ̳ґY2�G�%���8@�������cs���l�>�� ��S0��yc�t��uX��Rc ����MRp�s�\�RH{����;���H>�	�I��@<�aY�M����}�ӦWu͑��ʜ��müZB�>��{�iX�����!���P-BO��@�Z��G��]���3����T�Ϝ�衖2c�,����E琢Ά��=�:N�)v&U-����lQ��z��q��x�/ֵ�J�i�q[+��ƻ|���K(f�DPW,ϡ�]�%������9�GvD�8���"cy�F�wtkr$�45�La��A������ɦ����w�|��G;���}6}�/"5o��S��-,z���)��ܖ�k�SkX��� ��*�V=�X�*�]Jk��F��\c�{�݈�J�0h��a��r�VMx��SlJ�/�v��^_'�|��	��-o�j�s􇧼��⣇�:��T�b���D��T!o%T`�-l�Q�%��)�ʥN��(WE`����l�=�9D���b�g��}E�)v���B4��خ����nHG�l��r�|��E(|��̈́Z~�9W����T%����:�˄>��1��Bm��s~t�<�b:iR���P7�ZDX����z���j��ٸ ���em�6��l٥�'y@s�E�G�۸6�Z>ox)E����x������}�M���ꊾ��_*�<�ؔ酄��1:��drq����d��ڧ�m!�B6g����tW>�	ߡ�懻z����%�혠�`��r|���5G7H��9��B3����Cœ��\瘝T���Dj��g�V�i_�;�J��7Ľ�Ur{�2K��H�z���Ė���qXpF9~����_bП��yB�2nk�L����4E�=�f��tTi��̸�L��=���N�Fu}���Ocj�V!C�ňPl��sxI����;���ײ"_�m�9ˌ��M�|Lwٓ8dfB=:�8u!fB͊9�w��>ݱ
��g�eA�9ډQ�W*o2_�N	���g��t�1>�f�Zg6�6�\�n���εw��+��o|宊ɯ1XLT�0]��ܨ.�X"�F�z �C���ł����k$&M?�=,����}q�Z�3��Yط�~��q��Wq�bl������GAkp�c5Π�c��Oء+68�<s��7�����N�^��ԦxF�a���7cv�\�=�2�=�i�(%$6�2�-�u��D 7���x�}~���n
��+/j��x�j~���qtn���M_j�)�+z���.��$٭r��
���dM�6+�bbG�#��Q�w����U��F�Ŭ;����+[�.�q�!vÝ��4S����bh�Vp*m���v,��w���Պ��W4p=�tAFP����eH˨M]<y2���V�	Vff+:��v����ސ�ơ�,=.�ɬZ�u�����7t��תh�Tl��t�`����jwr�ak#LD�:c���WH㢗d1�ǽ;�F����y�f^�� �j� �>2���9f/&,��'�����Q5|�^e��v��n�W*�S�dsPQb�|,=5�4*_=h�
���Eu�N4�i&�����<���8T��&Ӣ���5�Z����w��V'��G��o0�s��[�uX�u�Ft�wn+%��i	XP�q]�Y�(*��ؕ��0}��>�{7;k\,2��{z���T1<�u�.wr�vT��s���PFB�@)�&����w+i"�
��u@�wAnaR.W�^ga����J���Y/���Tʻ��W\a�I��{���z��#��7�7�i��Nv仗#��FwMի�&��Y�E�7O,�٩��[Y�mt��4c�!��}G��	�m���c.h������Ƌ�-�}v�9�b>��'�ڗ]CU��f��]qʍ6{"�=��_IV���p�9�[��a��P�9��O�!���;=~u�iߐ��:�Y���ҝ�ka*����У�xr������e%{�ܢ��H��Q
J�^ni�c���@Kj*Ka���Mu,q�w�os{�6o!�z�.��^�vG=Qe��u�v��_d����kl���)�� �G�KX3��p�qn��P����L�ȆK�*wfJ��u<*�� ������ښ�������4��l9��F�Zl�භ/��v>p�	n�a�$���xӶ{��wugdY*��iro��HHm�ӌQ��QѼ�Ӻ���m����bo��DP�������|c�=�d�j41��c�R�����,Y9����ѫ��ybi�2�Z�Ul�`��� ֖Q�A�ɋ�<'������k�T*���vB�6�d���
�.�ސ�Ʋɭ��e�15�_5����^9K9�ڴ�W6��A]N拾��h��S�՗��֜��s�儈�Rď=y��u����S���Y��h�%�p��87+�y:�q9[��7���q��z�M��cm�oCɭ�n���q�.�3�z�Ϥ[��.H���MZ���ΰ�k�M�6��` 96��"����*�w|�
�k�*��?�߷�����(y�i�]�K�m�5��$]o㸵���yM�:!��C�#�[�VM�ٹ�AOo�yxf�S^fP�t/���)f�:J�uv)����/6U퇰�-���v�v�;q��Ԓ�,vv��H��p��g��SF��o)���Vڍe-��5���.;�Ze֔�f�)�|��,��)�!���N]�^k*nk�l�5��u���_��fR�yo�WƧm��L�mb0TLªV���e�!�f�-}l�����Kn�p��Y��$rKh��b�6Ǿs��̳%Zʊ��.���(�Q>Z�([}Z��r(��̧��7��J�'�m��X��$FE�KraY�U�V���sB��^5)�zۮ�>s�9eU�+��L��^�\��EL���Gռe�DOiV>Ъ�-b��Q�*kZȶ�*#R�V��ȮK]�dER�JU��E�1�%D�5gR�h��(QTT�޽p�*��kTu��No���/10������8�"ǔ,���K�{�*�k�U
�j)`��w�5�E��QNYrTOv�<�ҍ�`��-����鳭X����T��pS
�Ff��
���c��DLZt�5b�L��[�|ἡUB��PQa��/msY��/T�f��  ����<��M��[X�\uA��L����\N�n�@n�����o��3 ጰ�X'�@�w.?�����^���������5l�k����	��[W�+ul�W�*�IR���N�,�\'�[˴d�y���(��͸��{OB1�9R.�d�e� ��
̼�pxZ�\��~�Y�k*#W;��:i�vs-�\��[6��[;�\��M�l�}@Sy=�R-��=,�|/��U��ͺ�(��>���}Kh[m��5�o�a�$~����3פ�ȿCj���M�b���Ǆ�{���^�aa��.����������l5��NV��ly����7�*����-'��[�}1���|Kג�1�{;�����r�T�@���(t1�ږi1в孓�Y�t�E.��{$��OqOд>.ɯo�]�V�+�2�,�ۦ'�X����'+�y��8���=ݗ�{�g�H�N�E���f(��o�-FW@�?e2�����L����"z����jR�n�����J�c����/������v��82�k����n�)��h��5�Ff�,1yl�B{[z�S\�v��>��k#�D�a�OY�����"��+չ�����{6��(4/�W��f�5�H�lrG� �)۩/�P�]vfʕ���1	��@���R�]�z^��XRb�9�k;:��N�2��7V27J�2��ɼh$$XlG��Ԓ#�ޏ�.��kpoE5j�N5dnf�3�� 8;�����Ǯy�f���q8�H��7��~�%MsQQa�>�I���:��w�p�����Cע�%ݐ�'Z,s��}��+�(Y���w�����}�N��Z���1�\w��{�~��ԕ�@�#��0t�P��mc^=���n��޽�]�5�*��Lj]g�uzpez�n��J��Z���0���t���N���x��wi�ݫ����yɷ�ʵ�`���}MϾϾ�`>���������'��zY��\���(<q-{�h$���^�E�]oX�����	;(��9��ĩA��k����L�%Ki����	K�/�;�_9�-��:Ƹ�]��8���u�c�Ɨ2�,�a�֢�핔+o��0������uC���:4��8���J�)����vx_E����vF�ϫ*u���A�t˟1E'��ܡz�����D(#ghv(�{���՚��G3���;�ѡ4���>�gO�A�c�	>�G�[b���CE���<��S���ꛅ"��$�
�<�T��Wh�4�!�{����eM萤>Dd}�n�ٺ��ٳ(����m�J%c��)����x�YK@V�v��K���8{����`+'�'yړ��}Eϲ<���=���ts��Yo!R�Cs�o^��/�wpH0c6��k6���[Q��Ð�S�.�y.����zLT �#.�l\e�I/�� .6f<5߇���W��=�N�ݩ2�]�d*���\{:b�Q�*��\'�-t���c'�	���H�^�Ly��&\z'��)X���J�6�&��O�H�㚍�Zu�D����87�N�Q.��O"��ч�U�/��%���y�����f~�l&K<��Fk"N=���O���[�������Fq�U|U�q�7������YS��榎m.�����Jn��"2�]r�M׳��7⨂_��jmas�TS.���$⡉#Q�o�fk-=���͗��6���{=��ϫ�����gקJCϛa0p���sL��mZk�Z7^�/U�u�}l�]B�L����u�*��|5�	G�5�r�����Γ��>1�㢝�/_y����_�T�;�f��芎�WR��xBI{�<g垂�reZ��l��q�tV�3Y%;��#�mov��4�n|_\sJ���:�.����c�r����$Ʊ��[���_[�0@]�Z�{���M�ꀄ�f�_�l�2�Ʃ��2נ� �^E�NW�VC��WP�o�]�����{���6��q�-�~T�����-�5���ޱqH���b�0�ާnζ�[��-��rS���Pv���kܺpRv��}�bQq�v�ڦ�\�;�(��Y�O�6݌��<�5�:vEi�Hi��s��>[dV�Kri93��G���E-�Q<?�U�\�:{"�Og�5}����P�RZ��i��UlNr7M�~�!6P��	]
Ǳ�E��_��o��7{��?�?�' A>9끣_�2�`�ex�����P�ͨ�Y��@�bw���9�Z0X�j�ԼM�|�Kj���*I�'�@���O�AcԶ��*zh�ܦ��MFS!3;XN�ڴX��Tȹ��cu���=t��y�ͫ+e����4�F1���m�E�l�ضO�q��z5R�d��SfPޟ�����I�T6�������l���m)��w٣S� s5������EŹ�E>:�O�~���)X���k*>X�z�Oz�2��ג�p�^�舷֩P�����TK���%�E���Q�9�R;^�F3�W���x�yuiZ1*ݝ04Hc\*0�t���S-������J��,����Tsv(F�$����a�6��q�z�R����P���LX,,�
<�"b�"0./'�3���}��ޛ�8[S�`��������0������D;a�e��
��T��T�S��ǋ��=Օƿl��VA��ډЏt%q��;;)�yI�Ͳ�Ct8�
>�u�v��~�{;|���s����Z�)�WyW�w8�Zpe�7�z}��=Fg�&�$�R}i�Xb�^N�5��N�n0�ۻ4��1i�bƦ�сŵ�ۊ�A�mR�����Tge��u���UUc3h�/���aM�Xܧ݌�@|����w�Z�:���6�="�����;���y��p��P~��_w C�x�y]|9H<y�=���ol��D�Z�
"�F��L��2u�1�ºΪ�S�v�xE��T��b�·m5��4��S��Pj%�7�܂�0�G�:�qs�*����jJ�$�AWI�1���(�и��v���f�	I�#.�ڲd-��u�!�H�C���G��v�;�曬g(�+]�_��V�+�}�?_�C�-݆����fdeib5J,��z����.������U#����I^��+v��E탌w�'6��u�)��/4���4>��s��L���Q��I3�b�l[[��~���ۣ�0��5�c�f�S��Sr�@Ў�8伧:�j�NV�y����׵�p�^}͇ea�54�.�q��zvg�\ﬄ��m����=�9�?)T�}ҥk�Qi�]"�Ye[j&�6��WV�T݆�=�z���@����u\��/ג�03;�O�Z�o?|9O+�oH�D ~>���k#R��L���۴�����9%�w&�f*޷�fMb���^�gهv��sr:E�r�Sr�۳�zIC-��;<��lO�a�Rr�y2��}�s���J�:��5�r���u��6�`���%$�I��
�zz��Dl�[
䗹�9͙�����;��{��$Q��1Vc��}!���c� �Ht�O�Oд�a�#o:)چr�jܢ��tq���5l�q�e�����ᛷ�w�Iē��"��g�W�bR!G,�	����8�S;�֘�ϕ��#q:7��F]�M)�.���u�u)T㤑���`�<"<�0�j3\��[�F	}]�:+�Wd%B�;���c��խ�\W(�c����if7D�m�L�i�o�3M�E�{��n�<���R�9F4��Ggd�'`$hcu�4�UW=x����� 8'Ke.)v���Ϯrj.8V���^F���~��>�G��4�r[���rc�f�3D]J��gv^�����{�wZ����������_�߱0x�X��l��^{�Lk�P/]�n]�lA�M�Z~�Ϗ�V���x��P���d�gʛ~�a>��nO~�=ӻ�P�zU��0��e�^��B*;t������R3K�c��J*;c�t����}�O�To)��1�x����^��Xlm�X��wj%T�#+����w>;X�R;#�(���`{=	����]��ݻ��9�({����VT4�EA�R��h�ۚ˫�h���ԧ}�P�(���L_�ck�n�<6�'AB՘]gA��t����z��L��kO\��w���J����TŽ��9�giwS�D-�
I'e�7N�K�͕��;�����?�{�;f����t�5|.7k*m��Z�0����R}���m�X���/�:}G;.eO���������z����w/�<�f~�ܦ��ŉ���a2�QI�mȬЕf��F���
3t��b��/*|���^4w$�Q�t�F�qB9fR,�1j�h������J|�*Ig��n�<w;C.���6���(ncE+HA5Lx=�T���"�h/ٰ	�|�}�lʬ���aƫ-Ti��o���D�^/˟�>�f�nɛɎ�t����ò�7s��׾��:�wD+#v�^:�0�r�LS�uR�bKrsN8>vZP9�R��	����ca��+Z�uOd��CIt/���vH�ƌ8���#�o{gOu��������SHx�Z�+�y�5B��ދ��|ҥe����Ǻg|U(q���׭Gs��
�.(�r��7N�?	�򊧋&�1��О!(�+%���)�o����[�	]C���F)-���Fo3�N'e��+E)��uIV��o8&����z�_V�[&&T��)�Ph���P��ߔ�}��)<"�w�&<�G���,X̚R�Z��?��ݾ��.��<,���U��8ͽރ�e�R��Ga��r��p1)T��+a��-����ۑ�_���Vx�i��_}=�"��K��P�:�m�WӨjۓ:�jW��8r��d���	�&�:����t���n�DNW�n�i�g��-�lK���ͥ@h�.�>���0�+"=v��m]�Z�_��9].����Җ&ʮ
ҷP�kzg��e.�pU����ZØ�@��xx��ݿEUC�S�'
���ƹ����e�;��P�m"�,H*m�O�v�掟JI�w~�L�����Gkw�{�(e\����5�Gw]�5��2����=�X~�;&�:a��+WN�p/���c�#���0{�bR��(Wu�%�_�*�ֱ�	M�	���6�����-*���W\�xO���Ma��{�|�)��0���@[5�W��ЦډR�����MQq7�u1�����N��u��������[Q��%|��T�ԙ�G��H!��Khe9��g���*gKe�,;"&e�?%�m���W��Ɂ^�k��+v`z6�hq�IB�L�xo���Z�ܑ��r�vP���f��yNXP*��f�I���6�xFǚ��I~�7|_g)�"^k��~��=O)h�5�؞���gҮO�Fl�6��)I���򤁪�~��oh]�',/[�I�������G6%[|C�7�̩,��y��
���MaZ����W�u��N��͉�5���Z^-�̯jɔ��cf�]Z��E&m��6z�<�O;��,�[Y6;yO�
����v��Ԧ��[W�-?������;Vf-�[?S��%T��%�D��S��.$����v���/5��-dWv���W�ʒLb����О��yBb�����;��!K��T�A�����ṗs8�Þg3πب�#p���[ld�˾(->��4:׽,F�~�m�J8���F�k�X_P0��iW��w����v5���`6.>P̀���B�Z���h�F�5�����/�W}��,���6��x��[=Y�Ez}����xC;�xg�!0Wt�;���5�����H�)�]��ʁL�k"�:�N�F�
So�g�P"�R#;OT�z	Y����tۮ�,ڼ���8e5K�*+���oǭ3���ӱ��m��H�#�����Ja=�l>�Uue�ëZ�����g�ZK�����9cv�ͻ�0��e�
R�i��ӵ�Ԍ�.*k�pj���%}��_�ۋ��0�����g@ծ��}��٬`lo)�Vμ:kҨi�+[&�"fq|u>���͗��J">�~m��){R5K�'{�&��}�`�iu�;��-��Pvң]zɜ��ݦ�ż��?u>n=���Tq�Z���6G�MTwz�B��\��,�q�ut$�;h[a��_eΉ��ü���,A�v��]^Nm��#���J�Yׄ�^D���n�M�iv�P�/�!��c�ukG����|�	�n���1+^�B����M�	[v݊�Z�-�I�@��|}㾎6�,�v;�Y5/�sª��F8li��ou/��b�Ώr���G�{��U΍���pβt�4�ŔE�&�����Q���%f�����aA�J./�eQ��yN'KGH��+�a��`�tHD����i���1w�p�W���K��Y�s焱��(��;�L����~��ܕrr��Eo31���o�Jݿ@Ǔ��q�`J�ڄ���p��g�}~��gDس6�dMD%QW͋��:%�n�b�[h%��w�Iē*��	��dBy�aG,��B���
��Q��_tR��2��B�{P[S�`����*�Ɗw��F$��`X/������N>�����p3nv7v��1W/Eׅ='��"�*����?p�q��s�7��^+�6�>n�}��ٵCԙ��x�s�����Z��.(��I�Gks`��'a.��o��
g���Оc�%[)�������_l�D�*�"{_R�q���K��v��x�w��0�|��g���t�Y�����v���1��Mqz9�wڗ���2�<�aZ1R��|�:b�V�V]�L�Pn^<����0,M��a;�s���b��b!��LL��]�����k���٭�u5dn�qe ����ؤj�J��9]=��V)n����"�[xs=�é*U�����-��^�j+�a�;J{F��M�z`�j�D/� V,��IR�:.�
�W.u�D����YQ�[Zb�����x�>ݛ+�a+O�wcP���;�v���V��Na�S$�@���5�j���s-*j�+v�]`gyV���Z2݊aʉ��*�Σ�͊��!�71�C�V�5���JF����L[hw*�]��[��8j�H!b'g�tk�R�1g��j<�Y�/8m��"L�S����X]:]e���(V��n�;���tj)e�zLynT�l���F�����Hw�uvW=p:��ǳ�����q���sN�Tv��̭�4JW
�R�[����(Y�����ݕʾĸnJsL��h��g! { ��V"��
���;��V�u�Q뎑�Z����v��UnE�u��f��2�4�o]:Ŗf<V��K�%`�;�Z9|�YS�/�Y����&�逐��r��Dt���Ԁnj�`�W-�.�	��`c�(I:�=�{�e��3ڷ���(�0���wA���������]�&�3��2\�(]r��?�|vS	eګ��n9����7a,�3QN���/�8��j
<�E�+��G�(,E��w���Af0+���Sy�հސ:B������r/A�>����f-�z�f�z�� �(��,�K���>g�ӷ)b�\/E������s,�]��ZРn>��K��M�;7�"��ּ-��;s1���8���*-ak�3Z��sZ8����g�X������Bm�'V,�KU��B�*1rt�l���=�o-n�p�g
�ڰ�fwY���;��\�^���WS6��N���A��˱ Ɩqv_'4�ɜz9W�v�-t;���u�9$�4gM/N]���Or��}�:����5}��H�k��Y�X�
y"쥛�ޣ��}+��-x�z��X ��;��.�S�=Z��9%,k7VXz9���|5�����ެY�]:��<�TḓV�{�d˱�5�rrD3�4��*Hd+ws�T}��)#���:VZ�K�i�X�h!�R��Wf��a5(��	wN���-�8��1ҥ\��ca��˷t�K�+��vP1�
�p��坽Eʙ�TȐrfV�����相�}{+��]Yu�Jr������T�oHG`����k�f>6Ѩ�n�)h��Enq�;���L�v���z���v�Zu����Q���)\�j��ܠQ�its*ܾ��(�+�C�SI���w�owe�˹�S��Ey�`xl�Ǚ���+�J�gM�L#֜�N�_wnfΒ�;r�\�b�);���Ö��1�/]�X��W��^J�ȃ�ʗQvI�ols/Aʼ�'-���$;�W��#��b�q�oy��F�,��Z����_K�[O;fUx����D�N�����rx?HEE��\�ֵ'^�,�+�)j�چb�sP�ȼ�>�^��mM[)�W���*1A��T�5�=&�u6��TC��p�B�)DS�yJ+Ɗn\��Kj��u(�m���3�¼J����81=\yü�3�8Ԫ�h��T��75A��;�)��z�B�ն��SXҫ�u,Q�͐�&EɫE�2"&V�v�UR�n��.�4���X��cFv�u�R�
u���^9�-
״��X�y�9E����,F3PkN[��C�s{M��/-�o6�(���sV���Qƃ�x�%�� �UU/��do����Sy�yҠ�\�Qm�E��&X��wz��r�-R�1]{��1j-kJ�iFǌ�j�,Fq.�<�N
U|���˜�jX�é�Nn����8 k^�[�W��̯��{�<amm�F՜���U���m�
¹*
��_�>R�-W���X}5>����e�.�5R���9r��Z�a��K��V�&�39��Q������p)J�Lr�L&o]��km%GZř�6r�0�__ʴ�x�a��P+��d:w.Z�]��gIa�m�y|��{��/L��'��I��!__��`t��j�v߽�斣�m�ڒ���Bc���+�LMk�oؤ�w��<��ّ�{y�=�忧�q},��w�gx��p�����'T�ʆ(J�Bb-Gʶ|�|���/���#��B��-�b*���{s��}�u�	�zM��.��7�(��<�N?��Eڟ���EF�O�#��5âUbUL�ve�ax^K;��Tw�{.�yA�2W��%���P�#��I~����޴jΤ\�&y�em穓2/�C�}3.`��w�s�ʄC��3e�Ȝ�:.+[%��;\����_>�w�?JO���w��d�7+��c����>�M�����#u����QI����4�&����7��=g9CݝRȏSG�K����Ѩ[�Z�����&�[�s�M��n�{���M��ur;�\��\�焇��%L-�xZd��69��Ƭ]c�1�]Vl\��+�QJ�f�)g��_�����w�u��,����~��]2�2)O�)����b_/���6Xk\w���c�mOo>���Bh��qC�~�(��Q��u1h�����Ը2��6�Zg0�|�	�"7��˫�Jȅz%����:��[P���bY���>�Py��17��X_S?0]MF!N�����ڣ2$K�nBt������]`�I�>��*a69ʼ�GK�]�>�P�Z�d�ǽ���{�&K��<Y�Kw�0-����<���Uz�ч㖫�`�)�g��f�ElB��8��8��
��mYP��,�|m�ˋk9n�/���B�qT�ƭ���w8�N�}L@�.BΫ���xW)]��]� `��!��a�9��V:v�z�	:�jPb���	�?*;ms�o����V�Ҝ�8f���ZH9�`�9�!k���Vo�\�&4:�sn�m+!�\�X\f/]�8U��zh-��vF0Mꆍ���@1ʈx}�"�u��N��>.�	������#[�g��+J��ǉ��3�B�AK�2�j_U�[�w�ܿG��Mh���v��_!Y�_��k�C\/2T��)ܹ
Pn7�6��#6Ο��]�NӲ/�D����]����n�>k{Xp����mق�k����JPn��'MÇ�:�]�-:ś���q��h��S�ߍ��}fS5������lj�����&ّb�*'b��5-�.�؏kw~�3����ƑTnQG���|L_ǿ\��`�_�^��_�/#��:%/sP1>�������*ߛΡk7Q��#�c�WwM�]��G6]{7x�vii���o�&@E#y�N��\BX�wO���P�۝�[�k92zg9j�kU�遜�Ӝe�ԩ���(;�s��F�Y]��4:R�V��yӵQ�����_�_�^C/��1{��Lx��{4$�pf�|y�Ļ�T��Ԩ[�T�cA���ْ��U6M|*��zh��b,����8�Օ6����/!��y�5�A�sW�	\����M�+��)v-�����"����S	�{��n�'����{Vx��XnO�x/��e�9.ŨJ[�d��}��?E�y�*���'�w��^JV?4m`�8��*ާ�xO�xc+B�'$��m� F��W�%���P޾%�F�Urt�K�ݬ7<Mh�X*}�09~��õ�Z��F��,Gܟj��(6��z�2nk�L�u+�nh�[2g����ڨ�0�2��|��[��Q���G5oJ��
>�Aq�3�64Nl? _�����U�m��'w)���E�Z�3W�lZ����p�|ز�̀��o�Vz�����c�\�wc}];z����g����\��i�A3���!��Mz@�r��pF֤M�������gL,���G5�*B�/^��ms~H)�eφ"��B�9��qH(�;�5}[c�
�����Z��|�
�Z񍌽�yұ����6��]���`3��(iW�4Np�>@�8��1s��W:�n��r1Z�e�u-_�o��V��[e�A�!�J
�&S��*��	n_ȕmL턠"�y�ƨ�v\���50��/����R{я)��!� u"��}po�?et�a�ԛ��<��c8M��H��i��ת阝X�ۈ���å7Q�֛'E��P�(/~*���vO�:�͒��|��e׆'���XnO �~W���3�^B#��Ґ�l��O�>A��|�m".zQ�rk�l%ܮ�Sc�	;/�Ȳ�׹�%�]*�k�YH��-�0�궪�-�����^�-x��/�DF�x���N�5b�׻�A��:��1cJ%�e��U6ߊ�ֻ�Վ��և���S�2o���Gll^^;���K\9�v(d��tv��u��s�yO˶E6��yEN7K�-{1�<[�jsr9��M�>���P��VѮ���9��8.eQ��TZrp.�{�P�O�n���4�U_q�4��[/%s��6v}���Y��� �'�㙯�Y������0;y�b�:Ux�}cgU=x�W�7����Hgdc(�HmB}�ah8c�<V�Fd����"��y��5��.��#�)9�G�~}lБۆ6���*ȳ.~9��/�j���so"�fb��N^ţ5�%�?'���qo�I��^"R\1����$-�YY�\٢�,���L��c�ޡ[ӈ-Ɖ*�fXdV-�m��]n҂\��\�g')�mԨ:�䨺hY��#�)�_���	bg1E
R�c��-l]�Kܷ�2�`�q���dgR���f5��V?��M]�z^�˔Ҟ�2q��:�c��J�D݆�<#�v�v%�)��fT�߭_���Y�.�q�g�G�U&�9�9�|�C�����?�(�g��������L�o��V��;�-�f)�9��C�3���thc[dGL��9zaэ�j����Y���~]��e�M����li�u-���7s�kHP��b����9��qf�����^�;���4���P����0�v���}.�ă�^*v34=�Q�&�G���C�Q}�WN�)̈́hގ2��ai^�LE�
������Quiؚ�O4]u�hk�D��o����*�oZ�F��yOk�'za���]8�7�}:��d\���H4�^WkUv6^Y�u/Z�ڳ7h+�jˠ��P�m#"gj�K��&we�]� ���kB�;� ��[w0�~�=�&[�ǆ��>�ݺ�5BǰB����Ee
6�c6�!;>�<r������G��ퟂ�PU�}s��u�%Qg%�>>���1E'��n��H�e��L�4EDOM�ވ�Y-Uɷۧ�mJ�-���IΤh�br��7�
C�[МZ�r� օ����%f��5P���}z���ΌH��R�Z�}s�5�zI���z�0-̀p���ų��H:�R.����N��n����}+�u��ʹ�e���s>��z�E���F6	s�BS�`{�Ι��'}'(��[�N��ˉ����Xf&�給|Q[B���/(m����?R����U@��
��Z9e!�����G_�h�k�>|/me�*W=�S(���Ly� *}��ݍ�$����Ttc��Ō5����n��",]�R��l4�9���H}�)��jSr|sQǷ�x;��	��n��Ub�]C���˱��/0\�p����wU�֞��(���X,�3�%k^*�uI����9�wT��ޮ����1a斬-��%��ef�{³{��ʼ��#���b-ή}���=v��l�R�5�(p�йH�Ä́ņ
�	<���cS�/,�t�YoY:�e�1�;osЩi�7b�o�EOk�\3�
���8g���W�����Y�|D�d��I�d���&�1���չ�n_^�����BE��=��Z؇��[�쁌z��v׏FDO�g�X��tR���'���7Nqk�p�ǲ�e��Y �Ҥf��czg������pS[�����]_V��y�h���݌ƶn���w:�7|�~���~�Y�����]��m��'A�}˕7Y��obp���n]�@����<o&'�&5�;�$�݌p}�P���aPd�:eun��S*��=2���&�e����m�1у+��nn1��]�}�5�<�H���;=�(D�v�^5�U��W����yp5}��2��5y�t�u�p��gve�f(�K"cǕ+��� q��U�Å��wч}�MSCP�	�=%6בi�Mη�0�,�2���n,TVV������ʘh��<|N�?Yt�p�nK}�H4gޥ�,YZg�B�����4�ZVuЮ{���O�!E�NDذ�����}?+�ND��I�cS�
v�!��.s:1�h��r�@�.qD��k�@%yb�TCǕ%؏�%R��Pw���/P䶪x]\�k��'�&��·v�5$��fSĪ�8M��Yu�L����y�+ϱ�������z�c���f�Jv�01��=AUtyX_���y�w�ˤ�=�ڏ�L���v�1�:�.�k�z�e<��pr�n]�i �\_�Ң� u��S�nf��9d�vM;D����k� ���?�o��1�Y7qLqE��_�"�*�:����[L�K������u�1֢���S�RLb�؆�О�7�ٺ�O��Uԁ��KW��S`ӥ�?��0�[�hZX(c��yfh�HɁ��Ezߗ_
��	��m O��ſfuԌ��1��:�܌MS'9��kc��GK�St���s���&�օBs�˰��u4u��hI[�N�L���s��х͠�]h�}Ox�9w�x�}-����z9��=�7p�.��̔���
ך��Q���[�{Æ�M@57�2^��Ml�M�x�9)-�c�+�j�N�f~�>�vu�p�|ز�l�A�VjU/}h�̮��*��K�9O�%�t�3�"�V���Vn@W����e|ޜ���\gf�/yܣ2&���}4��R�^�c�wKs�`	��Ȼ6�r�+�U��|�����v�b��
#�6�T�M?�>,��Q�"���t;i=Ԛ�K���(	��]��`+0W�(O�D�>Aw���@�	1�Q6������߻{�T��/����f��Js�v���	���a��|ȫ�e�u]��q��OK8�	q��MG���jGL`��T׹��E�ݩa��5괥���3k�Q-y�)�H�~mᄽ��UM��靶¬~S�Oj���v����bF�8��ݼ��>x*����/�J��:�V�������3?�x�=GW{����f�S�\!�"jE1��O\��m�n��ب����E6�*o��ee������3ZCΩ�QZ:��z�2 ��x�=��7�A?zO���N1u�v��9�w����w0����e��z�t��1)[Ӭ��ë9�A�F���̟�~�5���_��>ρ���C9F���iN�V����'�
3b�d���P~�����j���ɿ��/�z��G�LS��JR��Y�a�#�*qfT����ӓ�aMY�u�%�:��4��rI*�:���>���`���}��u�\�NxQ���F��̇�0�Ѷ߄.Y!_
�V2���@�	�f����YCT��7�1��!�	�)�1��<vƜ��3���hn��vE)��	���X�>�����mK;�Iē*ȳ��'��dH��Q�Ed�Ir^���rzD�Ǳ��l�/���=g_��\�R�H�d1k��z��LS�U��+��q��%�?s�=sϺyP���L5?�g�>^�q��[^+�x2�i��iK����$q�ݒ�6��<��dek�Jw�27��c�A#B��#C������4;�����/b���]���?^2
,Re�a�ݠb�����{�}���`�(Y��ٻS�7�D�y'lw�EON%ױd\���$k�T�P���?�*ױz�+:]���:�Ȩ�5��d����iyd�5,½�X݄h��A���r��oc�pX���`��Y��H�A��
kб�i�O&2�h��*�^(���'[סn�����g���<S���������w��@Nf+eR����G7%���^��w�f[����p�G�5�k]�D_~��]�}�-Q��0�qj4�����0Y��������<9��f�ݻ���[H!��X�LЇI���v����R������[˜j'^)R��i�w)z��$d�S����i���uV�]�Wm����u����/R-R���M�uԶ}^y�3��⼽��J���C-����;D#��_�ƉnS滀ʺ_��|����muW�R�B�~7*��������v';�qc�^�l���H{�6���!�V�v���Z�;�[oQ��b4����',)%�f�U�^�y��43-�l�!h��5�WZaIڇb3fd��ШUY�E���W4,�Vʳ{P{�j-���5`�qM�r=����=���~R�n._t�B����*�)K�cvB+��.v��A��w36����@}�{��V���WwǞ�V�wg��$�ӑG�i�Ԍ-,��r_���o�p��U�?9�\.����Ƹ���f�>�O������;}��	a�v/��6X�1V_}PYV�.�*��>>��[B�B1PlMW�y+YՔy,�YW(�Q<yU��f t(H��>��Y6��(�����l��]N��*���}v�xlI��G�R�W������n*��l��i-ݼ�9�����A��g�蓴We�l�8�(wct���l�I/.�b3T��Ng��%uY�FlA��\W5��d��%9u��p���9���N��Y���}�+�m��m�)�9a��1C.*��5�Ջ���M���S�W[��y5�������5^;�g+CZ�e�p_-M8\�6�;ݼB9@�8Hk�IUzV��"ٵ.�C����fm�6�Rj6D��^kR2h�L�q�܋VE���j۵} �.�œn�Y:c��vv�[���W�We^u*.����Ē��_L�D-��e<b��Q]|�X�s�M$���٢��G�1�4���W[�ՠn�T�
���CZ@���e���)rO"!������é��k�DX��:z�oCEv5��ULu��kI}C�Z�y�Z�xv���}p��I��A�GXe4mUx.V]��.^;����,�%A)�ְ��-
����Ф�S:�`��:�Q��4mrS{C�.��*���j<Wqɗ�IU�PMo��-N�SH��#��t��xsi�>J�����{���lօj��ѵwj(�~��ã�=W|�+�s��i�[m}�gn����wC����؛�� 0��W#�t1�g�����zB&ȥ�x�7��e����Y���W(�۟A�c  n��-�,���!���Y�u����b�6f#0�7&J�U{���3u��ہ�$s�1ɊD!yv�u�ݔL���	��8����IK+�ǩr�4@�)U�K3;7U8�0N�C�����~}�m�]Sf`���÷����Z�!�;����  T9#��@�9(Y5e�eLڔ�c���2�z�r�bm�-+��#��9�k�`s��U��C.�sFPT�r�a<D���)��h�k IQب[�=])����:��3��z�<���Χ2l��Wez���E�/y���À�i��m�ղX��v�L�$�yQ�%5�>g5,z۩�q���{XYP���G��W�O�r��eCL��=:@3�Ovv�`��E�+N�Sz*2<ݽѲ�gV�u�[>�+��nv�d��/�	mN%��*pç�,'(�7v��t^0P81,E���`ʝ�D�1]Փ���w*��Sb��� �i)z���B��]��Dl�qRwn��J�|���Ist��Y]EK��c1\�E�fEMfgv&��_L��ͺ]]�̬֔���D�n�9�I�T��³R9ܶ�O3(��.f��uWn�z�[�ءt9�Nu�s,�2p3
���->�sK�4.�VD�V앃r����C��5Q�<"�gi��k�A��i8;�)����g%<W ���(]�R��c��>��a�Y�ܜy��K�ޭ�x�	7k2�b�����'	�݋$�H�	�F��F�;�DP�[��S�K��\�r�d�Z��b�\ʽ6LZ�X�euz�Qx�QayE,�h+l�����
ZX�ڌGY�b�P��-u���N��Jֲ"q����^v�X��ņF*��zʙ	m����ӣԨ*��ﻑ�8�V3F(�:�1EouH���A@TL��JiC��H����Tss���E���e�VV�-8��b��h��C2��:��b�]�-k]�����lb�W4�Ƶ���UQ#iYKy���,+*1'-�(�R�s����
�\�^���D�±H(�X�mKj���F��8gix �bZX��:�
6��j:�D:�C_6As
^�ys�6�T�����~7�����d��Ԭ���Q��5Z댊1YnvM��աF%�z����Y`�m>'�9���E��EJ#J�Z�֊�����E��<��,QUb�f�Q���h�B��|�KN�絗ܻ��1��>njUT��7;�:o2��@}o�o8�u%��+�������q�3J�YF�N��x!��)��T�Õ�;�̳�-���� �y��DG;u{��)v[�ip4kQ�@�?x��'Kٯ<�>�;$�.��f����_ƻ���z�N3e�!��؝x�TF���of+�9M#�c�sm��im3��d]��[I�A�gp��3`_+�}���|'[�ͅ���
��W��n��|�]����=,M8�T�&ʯf��f��	)�2ዛ+�����	9������}r�a��f�x�k*cx�K;t��u={�1%�,`�}ܨn	�ݳc9�H�h��GKbg�U5�����ڬ7�Q��ә�-���}֘{�j��Y�ts�b�@�\�V�ح�=f|�pܪ|���H����j0L4P��D��j����H%V������~��=�'���~����I����h��xh;�����lr��F���lރuw��^F�ۭ��63�����'q�,O^�t�iٰ+.��<5ݗ�a�j^Lъu�
= $ �Y��� Ӻ�����#�,�SZ下���Ti�3-u�w�欸�Q���6z�2=��<YJ���[{F����'{Dp�2�Y3�*}�Z��ޘ�����<f�Ӛj��r�0Wf�K�3�TU-%M�Wׯ��߮�/G4Q�5�&8vT�AԆ{���f8-�Y|Y�uqF�B�E��o
}��S����j"򧞛�H��L@��h{X=l<�.u�3|K�N�\��Tʊ�l<&뻈�$��� �~�����<i��}��Ln�1x���7�[^�a�(�ݺ����6�ܱ=v�jf��n;�8k:a��*��\�y��u5E%3���x�� �=��<gx���}�v7Ńۘ(\*ilL�v��ـl�}Y���	��g�d��A��4嬉Qc)�y��|�Z��$�5�_�����d�� �ĊlM�ۏqyU���ͦ�ƛ�!�R6��;rx�Ȋ8V�<s���'����{ݜ��n����W�T�Z�S��lR2<����f�{0�GVwe�B��Sd��y;j�j�����y#���qO�`;����c�^1�18q��y\s:���M同-\鷈�L w8�y"��Ipi3�Q�+��0n-���t5T���Z*[${��[��4��]��I#�ók\�ʓ{ ��eї�`�l,}}h�_Ͼ���zy��;<�uYg�I#h��B�G:c>�'aM���&�w7�]�d��bm�j�q�"��B��L�S�Uu����F3%Y^fǿ5��C�{^/=*U�+z&�{�U�U�[E\�Ku=
k�7�yd�p<M�����9�歏6�ʎ��|�Z� >t���K Y�N)ɫ��҆t;uo&ɽx^�5fČ�T:�4�\�)�E�zզ��4�9G��:"+.�m�")���ϳ��z�l�lĝz��g߇e_��ϺQ֡����bε�m�]�����j�n�+�|��נ҃A��6�[>�4���H�+����c3'vH��Y����G��+�X۲8������Q&��qLZ���*j�+6�T����݄����]�-�G��1��e��'m{�����.�s���b���
S肍L�{cMo"����E-׺����2�`�����|��/��Z)f�K!Q���k"�o�7���ڼ�ĸ[Ə���p%nr�}ڷR$�ZƼ�82�+��Cq�\o�T0�@m*�z����3x�Kv�>*i<yK���JRf��޹W�4����^��dZ���w�ܗ����N�7��s;}���|�W��N���x���j��v�m��w�Y�|�э���B���>61����ç�"h�l��;��!��7��nn���i�ƯX�U��!�KC��I�o��U���k��U�}��1�CV�ݑ�@w�|�[E�-��N3{'o��N����������|�!xk6�Uxnl�qn(�^<��'�0������>����Қ���5Nټ���.O`��T�԰�n�9$��<�(.�eH�?v9�~�,No�,���'���m5/f�]h���7u-���JNp��>�83;I�귍����j�{��F��U���?KR+��P}�k��"����ձ<e�6�I�n^��4�/w������^�U1<�s�c�ݲu���k�`�_����\�`�y.1�Nt��&�� \�%vvť���V�j�	�NA�v5��Z��eP�-+�Kr���,(6C�jž�9�̜
�t�WRS��&���W���s)^r��÷�1����ea�{��y�k�2uD�	[��5ӥՎ�L8\m���-�Y\�_K9��E��>�xj�O�M`�@{CG�{���0���n����3Q��ٲ&���i�2^^�����j�u}��@����]�o��H��-��D���W+bK�����]͓�웧d3�2������Zy�'�z�j�{wyr�����i\Յfj�_aۋ��H$-��7ق|ݼ���=��}V��{�m�}Yw��&=
�ǭ�����b�����ŖX{ԋ[��|�Y3o6���߷S��߸���������q���jշ����g$�nk�{�8�ņ$h�)q)���f�gxV��5�\��~�T<M�O�&d�u�-�|��S3�&�L\Wޱ����#C��k_��@8����v������8Z@��
��c({������o�ơ��>zC�>�=�u�а���[�z�j�䁐ȃ �P� @�:�����qR�4��?}_���m�/dȌ)��_����y�qJ6����L$z���ߥ�:X�����Q��R�=u��G��R� ��wR���Yݏ�Y��,R6_|X�2:w��$��n���R	gg�x����ޗ�ګ��Z���x#�33�'a����F'����Kj(�2�v��R؇P�������UV�ʷJ���V"�.sm�7���:[����T��/���Mn�u�FX����0�F=/9���R�5��g֭�=��d=��4��֞�`���9M[5{����3U�b'Q�A��(�Rv�ZԪ�1[�z���k�t��i�_Su�ݗˍث���(Z�>k"(�q�ǝ+*8�ɴ��@��8��<��j{M��[�=��@m�4�b=^�Wi�.���R�x�ȧ�ʳ\��V��2z,�5q>�t�?&��p["�_iv�8�:�����ni�51YPm���_36�⸥\��1�r�-~���NX�c��ݲ�-٦���CQ�������������A��?���h���x�eZ���$e�U���Z�EwR)��&�/����֛��)h���R��`�ʻ�┟%{�ߕj�������QM\�pqjc#���Xv��#���4���/Ga}7+�����T�$p�I|�J�!�ޮ�
.\R�}�>q
������5uD��/e�p�k�Yә�-���]�� KȢ�[��>,����7����	*Jw�,ugv�t���:$�<Ǥ�Z68�9��G�׮9�Qc��ϫ�=sc���\>߼�M��{�Y;�^Gu�'��l��v��92C�<�3�Y���R6z�<��ܦ7�Xdv3��LJ�O��n!O
꧊ݫ���G���v@>}����9����b!Y�8U�� �uXϘr�b���i�3D��5����T���R6�dy��=�&ͰO����n���#\�a�}�"2֠uK��!�"2O2���v�ʝOe;�,����jesƐ����\a��&vr7@fN*�2k�PN��*����V�-gm��m4#4�lY��A�ע��̮��NM�W���Bª,�%yWs��e9�BE�Ϻ{�K ������[�������_��һp��5�o�1ƙ���9�͇��m ��W�u�^2�w�i�`����j�ܑ-=QMQ�US����k=�b.��Κ=���ޖ�ywr�|��;Yp
��9R䨌ة�l����ҹ���/n��A=]^5zpԿ7*��\�ً�u�3"��X�Ä���b��ك�!��b���U�2���,����x���2�a�B�z�XB�s{�ҟ;���O#z*�%,鷷�+jJ�m�!t+w�fu��՜��Z�d��w���,���cq1.W��π����"�y[�˶k�&:�*m�,�]��W�f$n��4*{�糡�����3��h|�{�qW./� $m���v���d1���Uچn�Ů��!�]�v	��*pv�t�W��㬴+ik��|���kG;���ZK�%�k:�Գ>�@Dc�W���"�f��RݸNfo=�x�x�C���V�-L�}��Hm�(ȃ�k�*���Y�.�E�[���08�Qh�	st�3�
��}��1�m�6"�Y����&��+�U�̱�����_��ܓ����jT!R�2�Ca�8��x��^�"�G3g����2Qu�9	2/�D������S�k��k�s�7~�|Y��Aݹ�ۜ�3�����4j�;v^��t����X�U3.�W�/7/�d��i%��g �ݴ�N��ŧ�C�!�|I �Ҥ���ͩ���k����?z�h��`�/-��Pg���3�2b�y��T*ό>+��;̣�IƮ�����|���&PeY5��E��'PjK�qZ���ɺvl�������:�zhʚ)@��b��k�v۴8pC/"Pĉ��������Gۇv^&��e��<�\F��_�X�p�U��R�a8�J1�-��;w���z��8��m���mMw`1�tW!=����&���G�l`�W�n0��r���ďX�+�T�Us��n�^2���i�ɂ�!v�wU�����-ەĜ��F���l���M���uyʞ���]آ��'�g��T���$n�B���̟Y[|��#,a~����	l*7�d��Y��O>�-G�Ux�~�W�]���w[�����ir�2WX��ꡐ'&9
%���s���"����a��yٴ2:\���q�ұ0��c���m9��v
n�������V�W���^6�(�����5��I�{��Fv:�y2ї�dqc'1_�57I��`�6���zDF�%b��Lə�Ϯ�����$l�y.ԋ����*:R�u��qہk�n�m��l�+R$#yup�x\�1>�v/�d���T�%���	�����km���ʣ>�
�*]�%w"j`�3��9���,�LfmH:
r�H��ulݐ-=t[��0�Ե�=�k/+j�2H�p�\���J���﹛�{�8j;t՗�m.�N��R�)O>r�{˄��A6�~��`�մ%JW1Ǹ`�s�D�9�ڍ�t'��m'���\3�1�B�s|{7���6�z��+3[z}��'�M��L�aA9��D��̸Ye�cG�x��vt6�����L�SŚ�X{���1ŉB��yk7����G��o{��Ȼ�]d�	���)���~a�D�YhFH��c[WQ�۸�;��z���R����:�fջ��Y��pܪ�6[���}�y�Rm��H��q������.�z�����X�����m�fnLL�S�i��f�*��첵�!p�C�,-��I����D�����i�����1��W���i�k�6d�k�Evt^���Hn���ʗv�!�7�Rok<N��ɭ�9���{�Qa���Sl��o�z��GqG�W���g���zﱫ&苁::�~u�m�N��t:�RP�򍄰N�{�0t?H7�Rb��X���;�):;<w/n�w�yRޅ����Չu)����=�v�,�K��祿iGY������LK,��3�d��;�2�bS�Հ�efw]N�`X/[H	���3]����#��B�E�yo������a�����s*zr��k�
��l��aj�L�g>[;HD��9��)3�[4�5��7s%�����=�ƼH�N���l��L����k�v�eI6M�a|;Ʀ��&�eg^�博��K2�V�.����=1�rB�d�c���+0ݱ��W�l�k`�۴�Lx�f�
�ܭ��Mز��)�ntƪ�n���u����Ouj��@�l�r<��
�_RV���:�q�՘��v�=rn��ݡ:e���5$w1)fU�\2�9��J���� Yrm9�c}�R�=�r����M��CEt���橮oR\$�з���L�[��~.�N����%V"�����G��c!�gJm^�1Ԭ��9��QꗎXŖ���N���Y���������f�#��g�^��[�H7Տj!�f���1�w�t��]�]��j=�Yb�X�\��rV:�n`=b���o��TXLڂ�ie���kk��6�2T[qj`���2�;��)�����E��K(��gnEʢ�y1�x�R�,1M���DDm#l�f�_s��'h��^��6�<M�j;�t䩼��,D,�x%��ѭ�*��։�������lv���z�l�r�v^j�:��s�Kv�o���^:�"�וnWd�nDU�����4��x)&).I\5�M[\��-X�3�:����@�j���t��ͮ�^�Z�f:�+^#���Z�Ն�Vd���9��1ٮ�h
q�7}Ͱ����9u^+ꃢ�U_,��DJ��;�kx��QY2Ԩ�[��Nr���q�#��ձY�5��Q��������ER�n<��8��|���o�t�e������6kNҹ��N�/�����Ŗb�8�aD$^�m�ܓYi�*��aLU�X��:3Qa+�L�����H$���f�S�S9�'�t���<�	���c71[I�ڪ`����ŋ@ 8c��բ����z6�>�eL�p3(�`8�@�8-���5!��ruN��mu�*����kJ�y6������L��Qܤy����O��ks{VqYvb�������z�IΥ���[.����������v��#�}X��P�:�M��p��N�T�S�i�P�0�kB'<%6iΜ��ٽ+*�HP�)��I�B����p�Į��>�3D���ױ�1o��f�����V�'FW�#]p�Ζ]�TJNT�R��V<wx�b�̼ޕq�;��)N4b�H���˾ؤVou5ɉ�o���}zjs�9y�����J��5�VE%��J#ĨfVĶ5`���5��b�P���q>�s9omEZ��fU>棯1Mv\��¶�GRQ� �UX(��2UHך���/'�W����R&J�-�f�_O8YmZӍ
������W6VR ��QfNk5�#�mH�(���iG_z�TU��^k���ps�E+X�����3��1��lͱ�M�h񪖍*�Ug[���M�ʍ����F�G���Y|��J%T����̯�x&;l��(��-�-J(q����Ӹ�����U���u��=�W��V�<���юki�Uk�5+Z*2�4E�)�i��'� 4Dd�����]��ĩG_|�N�Wwmm�e���r�P��,}Z��v�Koi(��aG���ү�WZ1T�zZ^ۥ���)S�����bV �Q0��B�L�o� �����G�Ӵ��k�Q�TɵV�['+^.6�n�t������Q��GR�D����̯���S8�sP�J6�UUS��i@
vE��]�kzwrt�����}X�P厔��osm8"�WvӘRy�:� ��q�YD�y\u�b�5�\�4i33j=�j�J����@���A��ޙ��'CԽ�7�4�H�J��]}�����K����2��:W�5JƝP�dej��]ׂ\�>�w0�x�¡_ߟ�Y~��������ְ�m�q/����b�8�ܱ=rƖ���d>�N�X�-|�C��on�T���C^k��g`lf��-Y@�Ϩ������0��\9L9���͎�'8���Z�"fY�V64�7,���nZ�F'<���n�y�H�e'/���;ژ`$�n�n�5�����҈�%�#�R��]UE����n������ ���Y"i���o>��ʹe��CQ3@�1n�:g����=6n'�9�r;O�ޞ1�W@�k�'L��"�&���VF��r����!�c�������}�L�p8y��]nܥՎ��/O�36��ã䈋�^�՗��y�;����Ô('�D���J�u����S+Xz��]�q͇�
�e�m�����������h��w\�����Uu���M_����r�y��gK
�~�.� ��/��f'�Q9RW؇n�E�i^n�o��h<Zk#fn�7���ʃ<񮨧�����S��͎^����6Lε�N �������n����d�O�\悮Nc��e0��3yŅ��{e���D�g��']M��,�B���SK�;@D�5���\U��6�]՚�7��*�(>[���Z�6|E��0V36F��E����i��ǫ�A���h�v�@7Khyv�<ϐ���!j�ܖ8��L+��m�Ӛ�fs4���d�M
֕� +7��m���ǇyB����LJ�ع�./\��|�ڋ�Q>�����P{�#o�$뵶���Ώ5��2�6�nUPl&}��D4&66Ҫ������m��:������v�r�6L�;J6�q�Y�(p�#��#3;����y�y�Lq
� T�M~����7EK���ޞ����>�o6	��|��=������Қ��O��g�o$�Uw������r�~*����ja��9�������k�9)ڒ+.����5d�7����0�g�1ؾfck3&��)�y���'g�ŷ��.��6+N���}�>�*���Jrv�إIƵ�y6�ӣ6=����m8!����=�,f�5|�_sֿ(��|7i��9�S[=�4�*�=�X�*r��Ǌ����93$L��A���I�9=?�-w'�n<�}
����v�N��$��C_���}[$���3������`΁ي{��V���v r�!�[��m7���^��h�����Ƀ�b�ϣJ���C5����4�ź��W�؀U3`�o3��W��՛Ni��7�Z����&����4�(y�9�q#/s	���'x��q:��Ӳ��-jC���T��K$�	�������FtkJ|~���S��"^�jV���o53�?7�`+��������g��W*��d�>飂�N�����ꓶR=@Z��e�%W9�6��hk���$xvId�O��1��uI��B���~�Ýu��7��._0r���i4r��3���P�1�N^�9V\�\��,��ɫ�2�*��+v���ގ�>��;p�벿=}���ok��jxtw@�t��A�p�˶{�%A*Ҭy��]��*�	�-[��W�Z������S�d�B�0���6�$�wW^��Ǐ�&�Ӌ.���!���"��OlO���"5��û�+�tj�lN�7�`��'��<Z�J����MJ4��e��|4���^��v�3X�R���p��]��xx]�q��p����e}����6��>t��Dr�^ݞ�j�n��m���U�6:��'#{7�N�C
%_�vW	7�M�T�����o{dF�n�:���)��ѓyG݂�����37mZ<Ֆ
�>����z�v��o`�nc/��jo-�g��^�����`�YA.{5k���߀%[��:���dٸ� �FEm�T��,|���+7rL��l�u��rۏ5��6CnP��L�ff�7_N�zy6R1�jxmO�,3{O�C�Äwy����0I]���b���OYr�u˿�-Oä5�d6t�8[�lL�3��B3[z�[�5=��i7GKn�LgUwd�"{����M@�(�t�A��i<Y���k6Bn*��>�Uԧ�6�a���#g����N�t�|��k24�w�i����Bqe�}��oq�R�}k'����=�����v�-����r��1XJ��],��b.�Ѷw:m��Kj�u�J���%Az�.���H���w�^>��[��v�L�/zrעm���H-���V�Se��Y]o�P���dU�T�+&5���7���7�fMh�'
�����v��	&���:�^��v��	�}_t\|�� �q��2�����Cz��Q�ݖ�Y2-[�J�N�wvu����mF�ɉ����,~-ydE,9���L%���'W穣!Ok��	���܂~r��Zj�z�D�����v�"�->}K�7A��׋:U�bW7p�K/6�6l���e.����M�������_| ��g��\�;�URx�5��Οi�Mߘ��z���+��"a������N��`֜��αB�m�Fgpǃ�]M�.�J�I����e[��g�u�\>�K,�q[Sn��=M#�3�a���MVv�FhM��^+�e���-jm��M>�{cU�\s��!��e�:�4��;�^�Z���)��2\l�J��UC3oeԆ��=�3Yڻ}�u��46�#�:��Rm;�ڬ�Ov0��;K�~����:*'y���S�a�7{S�1�g�������%�B�E��!Nu`�����Q��Z V��U�t�U���nn4KB7"{�P�6���[��뗐c�12�|2������x+9nǯrtڙ�nZv"�B��<g��1p��,��y��47O*%K������l�N����|��1�#TW�W����Q�.��n��F�gO�`E���8S�n�"�f�
��z�#�B��Y��GHRT�X*SY�u;�:b����y��n��v&���"'2��ݗ�wqgH�<ʊ�v�T�z[��ל��E�{1w:O5�S�Hȉ�T7.��	�Q�P(d�ym:x��º�Y�;s_c��rד细Ω{T���7FGl+��9U�[1��F
��v/ƹ�X&vV��am���䟫wS����i�Z�M�2:Nz��=d���Q'������^8�h�ʯyxʧ�_M5Ϡ����l���y��{|�q�D<Ʒ�Vަ�u2�rʣ�vo|n�Н&!��١;�tϑ�)�4I7�o%�CdFo�9�x���X/+v�+�B�{PiA��Ȩs=y<[m��Uz����!�\�Yp�����D��\l1S������#��g��y�sN�r�wy2�V�Z�  \�enQ&;��\�o�Q/Q�@oY���?w@�
J���ud2 �776��u���W�,gz��#Ҥ���-�Җ�S��Tgk1���g
��q��L�ʢ���qO6P �q�R���:�weϐ7��xUu�&ɹ��ge�S�u��ƀ��iUgi1W+���#��V����f�Cx�<��x��p�q�;v��� Dr53ѱzn��VT��k6�Y�bx��'�������g��Z�g;����ib���5��ѓ�rBz�ގ�������6r��α��O�OIT�{S��hlF"΂��K`��Y����E��EW��t�r|��ǖסR�2ϯ���6d����Z¶V�?$Z(FnȀ��/[��I������;��b��ӭm��dDv�w	�o�?0j�w]ǳdf��ݗ�w:�I�"�-�&�s�bϹwg��{�>O<���@���c_��NY��*]��,<;�����u�L�Nsp8z�u���S�oZ�� �g�:Ż7UH{����M�s�ҳSG)i�i����S��N�r(����W�Z�m��3ys��-�Qn=�Ԇ�2�][V��+2ܿ���W�����:��n�Kվ"��qK�:z:-��=��W;�T�x^6&s6�����|�
�;�U�X�ɺ�b��b��]&�"�ݡY��QS6��m&�QPnړ&�'v>��G$�W��_����4~���U.������Yu���Vux˅U����/�ڲ椶p�֣����V?A�n��`qH�k%]^W+Ȧjk���y�\�:'4s��-M�];e���Q�ZƔ�1�U��۶7��-v6��Аzl��t\l�4c+��R����ݹ,�G��"e��֛8�gF��f;W������;��@AN�v�����_�GG�Zy��BV�q�r6��9�9���w�o�%����-
l���ق-�ޑQ���f�ME欉�ኗ�-+�9,Ś��W�����a�;ieŘu��#f�ZYv�g������Bd���$���H��\�"쒭�q��+t���X�� �!��o):�Fe$�ӣ����4��ɵLZrM�c7Nc���h�p�G&ݗ	y�� @Xdn�������OU"gf�Z��g��;lN^��{G�_���lM�a
`K�kG�n��[+c���L|�K���dB�p�#��	)��n������k�#y\}"����y��Q'*���#��Z�ˮMf��;s�5�Sp�$�9�8V.s����]�	�=��>�kp��c��3f�Hm����s��÷7pV����#e����a^��E��0΃v1�5�I�b�S�ڥ��~�*bl�~��U�Naˢ�\#.����rJ8$���V۶�uc��Ϟ2�~մ,C����Tw����l�F���Vɮ�W�-�*��6�"ͻǔ��Up�`f���)?Z��{�C��u�@s��[а�����ZԪ�'�e��Z�����ws�ݲ�p*8�5������]䤮�z�}Mh���o�$�V���=x�e���i��r]C��͎�M��Z�^����ۅ�j���j�NyM®���בF�=C��1�m��wH�&�OM[+���[�n��U1T����~�����C���99{Q�D���l`�7[]�`G�˝�^Ļ�Xc�0�0{kmcͧ��1[G>]�ʒ3�ݓ��c�g�\����Q���$Fz�/<���d�`*�o��S�o�H�a�}�����ںYi�Т���4.�;��ZuWG�eɠG����r���=z)�n��Dr��Ɛ��c�[�F&q�6+����Ʋ�s,�߻��爼�LBݯLlm�T݈����n�/��cC��ܬ��?|q���17�Y��?6�@���J#ocz�r[�Z��V�뿽8�9ɥ0ތ�&��9U���ّr���~ŝCi���m���~�6EU*�Zu�}�;<l9���q�>��0��.�50j�j�Ei��-۞�#���ґ�=
�GH>u>�m2�l�+"5�,+�<e�m�����nQ���);�������Z���5���+ET�KԶ+DGDً�<2Z�m�"�<�G�1-݇�;���FI�V�;X�N��&=�?cm+��kF�͌��9�T�0"�e���rp�^+	��!�
��h��͌�m�f�M��wFջ�K^�z23 =u,�5?'���e^�U�]�f���幓�;��Z�;}�F�\���YMq�T��pƓ9B�E��>������~ߤN�����^ƻP�.Ip��t]v1�9%oB.]�3yՆ+&]��R+X��n%s�\�Z�3k0��Xvucr�Y�m�t�v�@�����X:�+��.�Ej���3,=yG�^,g6���H�Vr���e.�Ä�&Ӯ�V\�z���+SחPS��Nav������N;�&�F�-��E�Z�+��6j`&^}5e:��6Z%j����������6s�ssY�3]mm �ƀ�b,L��B9�J���_v[w������k� 1�dT6�����������˗P���Ws�tY�n��G�cu��e�>�����ZA:��8��/4ʋe,5;o9H�Z�����h�Ld5Ć��#�x3�ծĹ�u;�35�v^�r��[�j	S5����#t�Q�K3�]�Z�Zz��j=
!n#�/�vlr�)�r�t6�l�T�@�V*���Q���V��W�tض��W��N�y�.,[��\��U�c�.z��rN����#Um,-s��&_1 ԫ��CY�l���:U��77x_?���Ý��`�������z�|Y�E0q��G�֚�W�����ld�b�@Dհ��'gGH�c;�����j���;5*�R�l֤S:Z-��O]n�_I��i�E>4��tp��b�q��L̮�j���2G��V�dU�����	�IՖ��=[�s̱�;D��6X�Q�P�&�9;�o�M�C#u���Z�WR%c���Xuƪ�2�r��b8�'H0�(�]�\��4�	��ڷQ�׭A�T���xN��&*�sC�D�mٴZwW/��s���7�&�7R�)��n�}�jK *�ecn�)-�,�^G�'-]8(mI�g�n�H��tQ7�3l�÷{�;Ey݉Qt��v�:��5�Ȳ�5\M�4`Yz�4E��y�W\���Sh�ɤ�p.��kb�*ۚ�V�i�Q(&�t���0G�-�{EՍ�闍� 2�mF(-�}��I�0�iuN�]����L���D�pY�j<�T��$�wP��\���:}:>ٰ_U܉g ���CovۙSs�� j��O,�3���G���a�]ǄSBS56�9�l3i��uh�}���ȃB'��(�-wr�E�P�'�V_m)�!4i�˝�5�@fVȜSAs{`�|��V�v�t81��X���Ovt��u�N�M�,�%�1uq��h����u��u�e�U�weNuJQ
GR�+����(^.�UY^��	��q)]�ҭn���X�[�6��;�n�s"�c͝oS�KO%��
3`�� �ɏ
w�X��Km�	�RT��v�`M��b��!]��Z�Q�˦�c3�g���u:�Qi��X�T��zD�[V���*��՛��b@D��>���&`���2�ed���a�3�x�n��v� �����;j��,2]���i��U�{㘮�vs�.*��P�B<=�{�ե:gr�i��ۻq7$�:���2@ �5W٘ 
�AV%Gl	֏�DQX�׺�H����6�[��[myK]i^b��/��/.u�B��\�Fŷ��8�����f��g"��K�m]�E��V.�n[G!jR����u[�!y���G��U9Jd7)��+�D�PNS�w��6��V�C֞n��+)ˑ��)3b6�n�u}5r���]Ǽ�`�fj"�Q�-*��m��%�uqo�\��փ�Q~�2ֶ��sUMZ/m�<k�sms�R���2��'0���Tj��7m�
i��H����
��,�h2YU��׉PY}s;�E}k�s���c����8%I����w�O�q!�U���=�q5���(���7�y�/�C�Z�{v���l�r�WyxfEm��,-�QkT=�����(�eb��am���3X(��9�$+8�+��r�3DZ�5̱�TE
%jZ�l&�S�u�V�62��G_��"�E����u�U�-��o�Uf��s��[�U:<&,d���ݽ�����@oRfFu	c>��E�j��c�����NV}�9t5�as��k[��l��K<`���ܗm�G�?N%Fpo�e����\�
h�s*�uƚ�����i��wl)�L�0�[�U�7Kkܭ�N��l�l�I5���bcO>��͑,����B���K��"��<��WNES��U��,�	�	Rڱ��G�����#��̕}Mb�9s�<����v'�=y�>��Q��/O��5�>�,�d�:g���B�"�ӳ픪��LH7I_6͋�D���s�v<�-���Q
 +k�O*�9�~���?r8��+�R���Zk��k��v�4wkx�O��6ϻ׍PF�{#��:#4��(z�]�x�ՙ}3��ė�g4�� �VlG�zT��Ndw�C�p��( �&��u38���Y���Ǔ�:��4:�B�,d1�q����5]��g�+6���W���*ƴw�ǉ8�Lo�|M�>i{����Ԯu�e!�趘শG(`�]&^67==�{̳G �<� ˧���q��+H�$��cI��W��V:w��js;��yԐZ�Ԭb�s_o+�-��W��oC�0�H��,�A�a�G��3|u����X�X�o��f��yǎ���߇Cn�}p֞ ِ"o�{5�7t����>I'�jy{���R)e�Cv�[@#:���lL�����q5�@fRޱ�.�r\=N��rI���Q�C�\�u�.��fC�KY��kh3�+���q����unFo}��\N!jQ@�G�T��T����-��Pܺ�������??�&���8%v/�9���5{���EU�Zr�Uu^{6�qӷsM��٥�"c9�V�{)\���|էM�^�]��)r[7�]Y�[:��	�ʹ���귨>�j���[,A[d_�x��bD2;�{9��$���a"�N0ͣX�v�%��6z�&��?�W�#����v��J�3;���(��m�EUG�tdn�{������{�V���Wמ[���RZO��nB�㷄WH��5��Γ��0
-vd
���W��C�x�"���7���Z{�(���`ZﻘV�V$��ZE��"u�f���2>uJ���&tS�pw\�WE6�	}�1qB�̺׭���ӽ넥�VL(��s$�j�sjT���b���x��4���%A����:����H�N�}Z�=�o|��6�_olkF�i8���z�#�l�/��s4�R�
����Y`�a����A_�<��By�zsg)Y��7S ל��w�ӝ�V�^��
�q������bۭs�������ytb���+]e��Xl���g�;���{s��Yv;z�pA���V�Ƃg϶f�ul��+�,��Ko"rzOR�5�"������3��qP��#�5�}!�!�x}[�޳Q�I�W���~[�VՆ�ʮpލ[�9�f�����U�W���}�wP�C���EM�Y=J���2���x���!�[N�v�B�u6�����T~�ׇ�`�2�n~^��g��0���=�L�\�y%-�U�W�[G��wn�9꼾=��7��f��N&ީ�z�2*�ޕ��(�OY9�Y�ҧ��q9NN����4}����j���z95G�9��V�g��2A�eD5)��*�AX%Թ���"�qN�/�S��;��6iƱ��8�G[?Kչ��Eh�'iN�7(~xR��;���n\����������g��2;��;/����eBW�VUƕ(�8�ہ�.�%�j��=j����{&uY�8�]Խ�Օ�IW�xК����Ks�S��~ޘ����
���Ky(�:�?uK���WY�5��Y� r� ~')���ɨU�ʍ�j� �Sy��4�C�ˍ �N+w$��Ћ���=��c�-/��Ũ��RO5D�pf������S��%c�fU�H�s�Ck.� �D��i�7[;]��Dv�Lnڋ��螲�W��Xʵ^�5��Ry��Ý���$��/��ǡ�}J#tlf��%rmlU����w��ě�O�"��,�u��'�	�KK^�~��o42E���cN�[z�:��enq9�".n����y��Hl?m����� ,)���'Y�ճ�7ڳ�x�1ڒ���
FC�\�X�l�1�&j���N:eO�ï�?V��q�}�����No܎6���rl)����t�o�W�:nr�a�� +�5)V+�;#</�[h0��;y����J���q�}�F�����7Y��YyfYi�9%�R�m��%�s)ME�vv8����o������S�nQ�ѐ۾u��i�03���>*J׏%��MJ"�^��Yu��5��/ձ�
��F�y�kٟ���se��4�\���G��e��+��J�c��!�#�J�,���cs:F�Tw��@�He,� t�\��V�M[~��_t%S�P�M]+3��&�ۉg,�l��L�s�q��㻞놥�v�K+mTB�g���w�Ɣ�2�\�𬨆m5kO�{{��i':���m ��QV�+1�a�If�\i���b�Z"MN��Wn2�:�7�=�s�����H�P9W �-�W�</�[V�ǈ֮G�����:�h?�xF�]^nH�O+t���]Y5�a�,������.ҟFh;���@(Ty�#Lz�u���wJ�
Z���:����RW��ο��=��ʿ�Յ�(G�zD.3q��ݎ��Ԡ�y�X��4�sff7�����'	&ߒƖ����XvY�ॷ��2�Y�`��d��{X�v�5���V�md�SyR��{Jf�2�DF�Z�(�!��<��|�U�<[��-^��c%�I��Q����ɉ^q� m�I3)a{��aբ�ݝ���q�m;�ָ݀��θ�]g�xO$3�K���ed7��5�z:G�͗����+���F
���#���[Φ��׹_im�{z<�;+��+�/z�Qn}}#�[k����B�������ya�b-Σ�Ngý�b:�Q��ތ����SO�&�pk�e�kǑ��^+�<�Ԭ��<�VѴr��9>�I��x[�d���6'��2"���}���GHcŤ4.e;�$�I֝����u��~>U�붭�֞+2"o�{5��wu9%75A�ݷs�Z�Sdwk�l�����(6�[5Ւp�}?	0��Y�����U�S��;X���,�\Əi?O1ɽȡ�dRh.�de�t5�s��
�|4�1����y���8ӝM�)f������M�;j�����^j���k��Vj�3٣���La�c�[�ͅy�����*���J���m�ble,R��u@�e��ι�j��K'�Ųl��M�3���]�-���YL׬!ў]�t�$�%�>[��b��`]X�f]fe�nٰDV5�{*T�F��ܹrQ�dY�+7P�j���=w�;�+g(͙�T�%&��9[tu�j��}\#�VԏMN�@�#�*�]t�S_����0	��l�<7�q�ˏj�PY�;gd�T?�zN��O\����U��̇��0VϬ����;�`�퀏����

|b�닜�W>>�[&��A��yf�~KhG֯�e�"��w�=��wm���$v�!B�Y��{��E�qp
�]Q��C:O,<�su����u�@���~:���̻�I�,#TǯUq}��E����w���{�bHw�ڔ�na6R~�s�u_���M�Y�J9��w�c(�H5o�;c!k��x�o2>n��Nk3�6���搘�9B5�h�4���X���8ݼ���M��46%"�Mʁ�)�i'-�۬[u*����x訊)�{�ԃ���|�[=��`1�غ���īmQ(��P�<*�6��9��LX+)��k5�?`E�a�S���������{�e��m�:�
Q$�;���d�� \�7��}?nBO�e}#w���y¿%8�J"I��	CK�ȌQ%X =/E�O^�A�;���̻�����}�s��˖
�땓ɮ���� }Z�BucE��ˬ�n�D�j�Wg9��⹞
�NR�ٕj�M��Z$��>cy�w���`$1�v��7G&�:l���큽�;�Y
�w<'�*.睲l�l!yu���/#w�b�Hl��
�/et\׽�&=�#<��/c^܍��e���R��l�����>����X�|�Vx�-�����v��$���"��֨�W ��xsL+�P4���Z��:X���cW|8N���!m�M_�bF[3,��K�5��g�o5�U���C�N�����ٜ�ɽ�D��97#�Z�U�H�eR��O%�/��S44JN��
�~�k�j�;�@c���w_oz��O2q��>oQj#4Z���o/[oѬ����'�m���Mˍ6:��	�:�9A��e붹	����z��R��]�)���#s�9+����>Y*�j�!jQ׌��{��X/�gw?���?y�^ލj������T*wZ�h�p�ۍq��:�{���l-���̸߄F����UܖD�ɻ��9�+M���N��j1蚩�3Eں���M�RW1ˬ��P�|��R^V�=Ί6w��qާ�j�6��L{y�CHseOb��ũp*���&)���!S&uLfVt)�޸*e�l.��O2��Ʋ�~#�[���WA�e�`"j��;柆��ɩ����S��א�;ڷ��G\�8����`;/�y��=j�5�%�WMn�3�8�s��anwH�Dv�۪��'�l�l}Y������k������Q���AGA�9�:�������[8�7�V�W��H�b�&)$o�4�ó�8�#���Ű.���lH��qfu�c�}Y�L��� �q�;���0���q#BDd�̯D�8%���P3p�l�+�wcƞ�l<d5*�E򘛩�]�	A��(���]=�<e����k�R��k͇λ�%~�/�a��o񏽏����WZ�F�-YW�������ʭJҪ/
���ϩ�����c;6��Kܼ̥5ӕ~�}�9c�e'N*�J��V{D��<VU�Oo�DD���N�;�������2�'Q�>ɨ5K+yf��&y�d㸀���$�"��D4����y��y�U�O��:�
�}'[�NT@��w�<=.��مa�}G�h��J6+O`�a+���=YֹV�\o�2�n�'��N�u��zRR�ݗ��޽�Γ�XffR�	�4�6��db�p��j'{׋�ޙ�#8ٝ%�}�΀�5ϴv�u��s��7%8/'t�a؅�ՒZ�mfG7��ҍ�W�ό�؂4���j�[�д��?S���;<eO�g/ظq�~�y���"�R����t��o��(5=_���'YI���<�I#wv�/�c�ɨD����Z�e��˙�l�2͆4��$�̮����2��X4�HZ�g;�����)��U�xm�r��^�q�^���nu�����[�|u����E�D)�*��{Wm�:�U�Y}��J:x`�b��ml���D���__�_Zx>��`:u}��Y����p:?���}Um}�v#>$�p4Y��`�תE�f7!��+��b���m3��k/�e��^�h�����cy+^��%�Ή���tZ�jƄl��8[=��궿��'���^���{�����{�I�! ����S��dRB�d @	?��1���<5gd$�H �CȐ$,@�O c 1 1� �  O#$���o	�$�H�$�1qX�I#I$bI�I#�HĒI�I#8���F0�HĒI�I#�HĒI5��K+@ 5�HI%��I$bMf�I$�ВIc	$�I$�� $�1$�F$$���I��F F0�HĒI��F2H� �I$bI�$��I$c$�F0���1��F2I$c!$�d�H�I��F$�H�HI��H1��BF$�B�|����P���� ��ĒH @��������~�_�����������!��?�?w�}�?(?���~�?#�lI!$�������@!!$���BHI��� ��?�?��'��	$$����������a�?d�A��������h�� BH��	@@��BI$d� ?L�$�!I���@� H @B$���O��?9! ��H �E"�$~�{����/������~������߶BHI0~���}��H}����@�oQ??�?	����O�������N~�{I!$����	$$����>���HI5�M�2HI!$�?�?�	�`}`�C��Oa��u�'�8BHI�������!$����!����? ��?z�?0>��a�a��BI	'�����!$��������'�~�C����=�~���_A�~����N���?Q�찠�8����'��C��x@�����
oy ��W��������,��1AY&SYk�D�hY�`P��3'� bI[�!(�Q*E HJ��TR�H�H�RE��J�TAT@��T�H�(��
�*�**��J��BRP����R��UR�UU%$�T%H*"HR����T��	DV�h��R$��6ҍ�T*UB��$��{�
*J)/c**%(D
"B�H*((�% �$�UH��ET��ER�)AQP�B!PJ(BU[eH��  ��PV����iZ��3AF٥�� �jdL
hP�4����T�ڥ`5�ҁXV�m�P�kPiM��YV�-�FR	�U*U"�($I�  j�z(P�B�(3��:CCB�:�(P�B� ܧp�B�
(.ꔶ�h
ՕR��-�e�R�@l�5�)M�6�4 j�Xm5F�b
�H�B�-���   wK�i��M#>�:U i20�-ih6J0*�Zk[*�m�M,�j��j�յ�0���iC$i��Z�kV�!Af�M((��	���V�E
�   }��(�0��J4m��m5�l�mb�m�)��CJV�4��U,+���+R������Xj��bԢ��a��$٪�*TJ���   Y�P(���4
�&
�V���-�"22�PY�
(��CR%��U
����m�T�J*U%UB�A+�  ����ژ(���P*��U��Q�j05��TD)�LTPP�R4����� 
F@�T�H���D�(G    0�TQ̫2������`�m����@�l��(A���I�j�P�L5 Q�`  &�EUA@� �J��   ��  &F    E5  �e �`(   �f��e`  -R����T�H**UR(/   m�  �`�3  j�  F�� M�` �h  mF  M� �
�р�6
��B�$JJ�� q�( �  P�&� �,  �0  & 
�� �
b� khX �"��JT��d ��a%%*h 4 jz�3*� ����R�  �)�$ʠ`&A��&�	��P0<S]�M�5�p�#8��׈�	�L�ɫ��)�>+,����3��mޯ���~�	J���@��$�	$$?R�	'�$I?b�	#@�BC?~��+٠M��k�ZV�/r�c���S����7sV9�:V���n��ǡ�9�ԑ�.��T�)���@�lf�f,��t��f�n�����ذ=C2�i"�#,�[X��t/��MR�9i�m����ջX�W�I[��=����8M8^�W`��w2�=R�xF!R7q�i�2sXd/eYC#��tS�� 2ee�ԄSȄu����y[��hq&��?��z*CB�c�CN��V��Mk�H�>[���3�y����o4Fv�n�::����2UёI��(�+�kL���e�/i�>Z{z5R�Y4)%$���A)v�>�goX�X�8n���@7Ħ��Sn��W!X�*�	r��Y��t@��/��I+h0�'�[f�&Y�p��[��a��K7]8@̘%��Ĥ�9w�QJ� �
2j��7��2jy��ߝ�u(4�ƪ^io6*WM�1]:�.!V&f�Uf3d\�u�(���Ɯ�v��PȚr΃�-F�e�+W[�yT�$�kmk��t�ƫN/���9�6�V�:~��7B�Tb��r�Q�B�8���k{P=�̫�l^
�ޫd�(�1��91�r��K�V����[Knl�c[	;�X�]�a����srmYJ��ORCq�w���t�2���cIZ�&�0*�-��x���Ca#uV��r�愲]�d45Q��X�6]�	���iwW��T�lEo"͘��[�.���i87&�M�Sw$ŸĘ!�����& Д7�DѺm%p� "�'Avd�e�Z���YW�&���I4�cr,u���j�66��0;aT���6�V젝�)�٥r�޹��b{�ܻV���3-$�Y�u6NL�	�^ޫwF<
������h-�@��#��ٟhS�դ�C^�b�l�YDh�*:%g�.�U�M홄n"p\��!�w����р:�R�t��N�j�9Z���n/NJ�Axc
����R�K�ov�AP�Z�CI@������V2��+�Aa���C,��:	(ǹSH�o4u�u�$�$-�����A���Y
��i�-�i560��WR��2��ӏt)Q����J��A ���,Z�nҽ4r�Xu%:Ux��C�E��d[�����n1>���ɧv��0!HG���$pPQ^+������jLi��͹�j��EF)��%{��ZX�b��]�J� ʶ���t�bs�c���[`:�[��⎦��T3��+
�iP�+��T/cx�D�-:�DM�]��b�*�a�
K��#�����{��bU(���Fd�Gf��< ��l5Dk�[7ge��5�J]���)��h[�]
fM0*�!������V�5��c�
��%���E�S�����M����	��$�� �o7Y�V�0�1��fn�5�f�#^�0���T4r^�ȎL˃��J��_ZO�(�iXS7J���X�:$R������5�k-��T#t���ˁm��^�Ѵ^bc5�ՉA%Q �ûD��(���ڲ~9��r@(K���9&e-�	���a*��5<*a��1��'L,�%�i����{�nU��v]0�L��ųX�����F�wW-ZGh�����PG0�j	R�s���6�e��!J*J蝂-�,0���Ȍ�3^��U��K�abm��)����r�1�|�fI�r���9�����Q�&"�f�r��)]�L`@����yݨt�U�Q�K� i�j����{�"�*p�Ŕt
�ܭ�:�6�eE6Ѿ|�=ά�b�Y��B�¶���bM���z��Tʹ-6,;Y�1��N�i��H�ۗrۻ�d�[!��k �ueh�X����K2فV�]8_֜i��[�W�r���o,���q<���`譼��d��cO�a�$ʕ�^�T�P (�啷tm��p�(B!­��ki˙�C��=ݗ�@�Z�ך�J�h��%cos3�*Vl����+tD�%�i4T���Հ���Ԙ��3��s6�4�q=lY�VVӈ�5�	T��P�ɗD�v�j9VV[�I��e����g&��!�,�Vf
U�֔��ܶã ��=�X��'�8���,� Վ� �Zb�Ќ�{�φ��ïV����2�1!�b!�pa;�KTUî�x��	U�V4���̺+.Z"��G ���C Z�ӻ��9Y��Ǒa ��� ��m�kS�%4�j��]ǗZ�]E(�{��㬀���[R��iF�F��5�H�6^��S�J�";)� 3s�`��+(2�+���Qt�Sf�gi��]ޱ��t���kU�H	YB�,Q2��Z6��؉%��Ov�:L�)P�MrcedܡHU���=�T��*z ��Ȥ�� �m �;tn��B3ᙯ�WIS%�*f�-,j)�j����]X$�Թl	�C��? �ZWZNP˺�y��)Ⱅ�V��L���fm,ȶ��#{�T(`�ͺ��LkM�L��0�j������Ŷ[��kOk@:�n�W��DC�r�!VV�`��iJ�W�M���S#vn����[6��u��P�U�,�q�"XQ�sf��zu�Z�SڶK�Y�2�J�����S����&�-^��!�ڌö��
���5���"c��.��գvUX	�u�(RCf�i?��TQ�6�����^)܉ K�����<X� �jƺ7xu7m3p�a�Me�F������U��.�ǘ�n�W�"]����m�6p�ڠP�j�ʚmL�I�F�嬚���`xMD7�m�{�^�F͔���CȢɐ�9-���&�Bd��A�����h���/Jv�0�б%�[�{b�f��,�Ėh�A�:S�E�^��Ґ�n��������@J���&4u!v���5�5�%��uV�iiJU.�]�e��Y�V�;i��0�:-S��/H�a�`dK�n�wCo ����U�X�cQ���������4]=�Ր�T�nX�����m�E�T�@f�>�[�8�58����,Zu��˚���`�� ���*�F���:Or�ň��7C��n 7>�f�%d/U�%�G�¥ME
��5�ӗ��R������_Z&�-�[{�ӿAF@��&V�%��ȥ[9f�M�QM���$���&�ƕ�8��%浛�%/@�^��6�gwd� �O��r�[�Zk"�1�I)�5w��`�zDM��D:skYZ�[����:%�0a����V���m6U�8��x)}�kj�\u:{�݊��o3�F��`�4땑��c	:;��UjV��tcs�#��9D��1eՕAr��	@ж+q;��2�ht�[�yI��iT5j
bZ^8Ȳ��ܭШ0� �3c�����hji��7"i�Zm�5����T��V(�C���m���,)Z0�a�>��j��a���!vj铙qc��t]�17��]ٻu���Q�W��E��q����Kmb�[��T�ں'S��6ط�8h�,��$؎۫f�k�A�j�LM��dZR�4fm���1:{�n[W���1�/d�Gr�pM�K3)���m����y���Q��3B6j9lR���Pdi��Xv��M���zmú�;���/%��k��i��62V2YqT�{CW�sh�������yZF��m�U��]Ӹf�h�WM�t�[v$�4��/�B��A���j�˺X8�e2�̅�k�2�]�P;�(��۠(���&8���V�F0�^�2��2}��2��+r�HP
�ezj��N���A����ٔQt�YX	�3��N\����( �������n�����v��B�bt�ı"�P�s B��n�5��.�A�fJ:E_6�2�lP�r�`j�J��n�GRi�H��$��(m�)]�&�љ �v��� � t�)n-�0�����(E=���
�\�u�^D��X!4����{Z&�Y�oB�`.�Gj�'b
��X4�CB׹���-ͼ�Y3+2�$�f�г�4��B
� l ��=�O�$�	��yB�H����J�ai 	��@dt�j���!�"�I��d�f�@�^�qn,����kj�!sLB�h�/P�y��8�T���n�XZaw�w���d��ˌh�sX�%�.�#nj���(�E��%���v�C��Y0�{����h45+B�`�H��Ő^�Su����r��R�x���U4��7Unf+J��7�K6
TAq���ʺ�)ԗM�J�&:cqĪ�8�[J�f��2n((����Cs5:)e�E�v���a.����@���Q��[$�
��X��-�9x�a��չ�J�)76`��P)X�^=X�u���VѺ����kMm�9Fa�v7I	03�;x�m���r�!sv�r����m��Ǧ��nd�J�.��pD��2�m c����{��*6
�C쩕hm�X�yz�%����pV��D2)A#�LQ*�
ʛu�Ug�s@d�q�:In����8���N�P�+*�l�j҅����˨Y�p�U�3F��Y�p�hِm�)+.�`����nk��u�f�c�X���[o(iB�����[Z��*��i���LA{[�8j2S�q�Z)�hTv�b��g�&Y.��%�U �tYn�e�P�i՚��2�k9��˷Q��&��	m��ɺ�'2���t%�m��M3��E���e�� �Sꂤ
�@G����u��+s^�Y��[��zY�����#¡���!j��i%�<��V9��7 �bԒ�+-:S^�XT�i)
.�e��(�fEV�J\��e�V��L�n���6e`I��aX��(2��ci	V�$chRw�^��a�Q�Թ��Z�],�+b42^ �
H3�HEt��q�d�"YXݣ{T3+,2��j'���,l�+h���ݬ4����eQT���ܔ�GM8ve��}�7�l5�y:��?�`�UV�p^d��	�ӺCvC����ݺ���X��m&N�Y��YH� f@��
8*�RyOi���t��o*�u�fR��V��rcW�֫�wBƕ��9 Xk.���N��q�kPl��a��V�Y	*�(�,��Gt�)Yv��*Q��c�_f���r�N�.�Y�C��&	OZ����)�w>��n7nD�kB֧��;t� Tj�g�e/������ɭӭ���ŎY���[-*׋c�T��rTR�Sm��^��.Z�]A{Hˣ�ث��n����a h&n���
86VˈSs#Ȧ���IB�-�cqlRb�"�n���=�5�`*�B�P9�݋�y	��W/j�{��A�e��uaʶ�A�-���q�kvŭ&�#��,�Wv�5*ݒ�r]feс�{X�34V��h6�,��ŏE
�ܼX_n�e�Y`<-̌1� S�1)����^�R�V��+�5���"��I��́^��چ���t3f�¸ld��rM0B0fj2�:��*1jbW���;K��sY��&�rh�Vm��/W ͦ2�'R�G��u���nK��D-T�Zߕ<��{u�YVn�j<�[�������1=.�F�ݝj���y��۱�wA�z����Z�ߍ�f�d�����E�s0�Z��KV(mi%Ab��ǿHH1ରq�1���Ȟ�K�JE-U����k,�X�����6�-,i�a���;y{4$��xu3{M��Fԓ1��#R�46fC����-D.0��ŉt&�d���iǩ]F���������K�3ʷJt"�xfۆ3R�܉4�M;ϴY)�KIW�����cC*��*IR��BVM,��J֩5�*EX��p��e4�IN��á�XT��dH��6�-���0�[VH�K+3L{�!,�+ [nG&�&��m��mZ��IL���޼+t�g�:pma	Q�Z�ct��,��n�U%�hSd��ӡ ܫZ�A���q]��fس7)���on�[���H��<�m�wZ��n&�ne��m��@QѠ@����-;�F����X�)6�qfPBTf-��v�
�b�t#�eb�%�Ze��z� ����q�]��nce6M�o�i��c3jђ�n�BS1[�V9��*�M<�(IyZއ7'��B���Q*"Kw�����2�m0c`�ŕ�� ްr0>5u�Ռ�L2i��+��̩S<����n\J\yW�#���nI3m,�-�Y��@"��jWF���.`6�v�U�[��X�/3kj�kF�#�����o(T�)�ݺ,X9 �&��U9���el�����2�Vx�,`(��7���4������a���7��� ���h�N�e�����:��L�@�nv��t%��ʗHJ��c�@bN�(��lL�(�u`ү)лM��k^.�Z۲��ʆ�:36��!�S1�:�ڢ��\EBj�E�V5G��Fc���L̢���\�zL[b�7y���"%���ն�Q�YZ���,��2��
�:���O\b���oNhQ���I����r
������ޅ��C(�6�Ti���-b)l�J��5%��1�6
�6]���)a��YVAIA�{�f�R�Xr)W��$�$�(�w@�!d��e$��nJ.�+͹.$F�ͷ�L8�oac8h�6�N�j�2i=��˗����0[Ȳ��㦱;7J�[�ԗ�n34�Q�G շGT͗�U$4����$�y�	ik�6��&���f�}{W�R�(�K��7�f����Jt�$fꎝ�ۏNh�����b1��{���T�%��� �/�&R3QӏpWM�y*](ktv�Y����ord����I
y�˛W�S����t
�ғZ��s��3�ݻ����\S��dЗ.6js�fp�ᝪ���"�<��K{x�#r�D���	��q�i�GQAN��yh��7c�֋��&�t�\U
�X|ֳ(9���"�Ҍ��v�%�U�R���Q$Cc�R� \'+���.�����;*\s3�ryhV���Fu��n��K[�.��X�!��z�B�2��{4yU���s;{�2�E�(Ѽc}�ݻ��T[�{]�#��9\`R�.���f�Z�]4 ��Ж�d���b�3{O�>���ф@�c1i?o:j��5uf�+��Xt���W7S��wq�Lu+�motw��n��ӡ�Fu�#�s9�f� �o�+LwQ���Wu�N�cl+1n�x�7ڍH"S����.^�z�5���<gC&��w�0ZMo&���}�G�o^�O;c�ǡo�l�֨]5�fN2h�o����>�4*�VZ�c���.�'{�MU�9�t)��8�:��/��M֞G�c�j2�����R:q�t����O\�YD��E>Pv�<�1���Zx�g���=�| ��  ��]������7>�X/���U�Hu	��)I�:��v�"
�ޞ�ڊ έ��_9 ����n��R����ò��ok�PM������.x��%;:k9r��Nᔵ��-�ݓz�[�w��*>w� �ti�u�%%҆�R�&�Վ��;�U U�2�І�a�T(S�p����딏�,�Ǝ�7�aÔ�Ư��cr������A�mn1�3ݐ�\8XU���n�f����P��N��.ޭv,�mV
k~̸ﳹl���MZ�����¹a=��ފ:i3a��;�^�ɢV1�l�:�/uT2u+��3�5����%��TՂ10JR��_Y�Qǈ'k�4�U୦�����K$�������I�<��,cS�D�V8O5W�X���4i{�,�r�t�o�PL[7�X�e�i]*�9X⦶�i��׻]��dgbW�����OY�t�`�F��(�(��b}�o�j�H�Y�A��_K��Y��O��� ��vS�w�.mv%PiP�����\kp��Ӻ}JdW�t�G9f{|��ћ�V?]`�Rd���ۭ��	M�
�آ^	Ks���|+�plgWb��+Y��#��2M��ѩ�#\U�9�p��m�����Չ)6��;un�t�7����xH[t�i����ۮ��WN�;���H��������0l�&ގ�T|�E�:ƾ��N�u2f�������nq�a�o��9b����[����j�)���7kn�[EÇ9���U�;mfa�\��\��d̢��x�{��g�{��d�o�=�Bb
2n.�e�:N)�t�����jJ@m`��}/Hb�6�:���%Z�泤���#����(j>z�?wJת_:)��N��к\qru���:�M��|�����
ۼj�
w��a�JK���K�:̠Ce��2�Xok�%�BF]�9�)�"6��kX1�3*`�Vvm�
��'u��M��j0x:���:\��\WB�;��u��ԩ��j
r>��*L���״�T���HY��|�A%9�3	��
2��u�%�TcB�w��u�hNr�;YY�i\��9t(�=��5�e�癖�۸zbmK�Y��v(�T�G1Nug[v"F*D�TָrI�DNiK۝wkѴ՜[��f����1�{m[2YSz��u�wS4HU�'�c��M`�Ad�4��Yܰ<\�:[��n��B6��2�=��R��F��%�yWNgT�ł��+����^G�)��6�v?Gf��k��(���năl���5M[Y�*��l�.l|$OF�_a���G����� k�YR�!g;|WpS��L��s�KY��U�!��li�OT��5^�֊+w�����ʶ_oC�3#���-U�;>��1:έ+�~�iqx����u��,Ybă)#�R���#M��ܖ-#�W*K�wvw��G��O9j쵰a�`��k1��]����±�2��0��i-ġu�IӊЫ�n��o�ل���!��L�52��qo)-��m'L�v6@�8�7a��\�p ��Y;�Xx�4 G�pXz^nų/���mU�I��QN�o�t���ľ�λ���zN���k�$t�4�6nHM�&�w�T5�0_u�fw�'g��N�3���܀ݍUw(*oR4�g2�r�bMJR�u-�d�Ck�`�x��3�'�� ꫻�q�$T��mu+ӨnB���}��#8���*2��#_ȉ��
�o�E, ��"�
�t���J--�Ùu�7�@��9,�x
��%/�9;��3�僶���+`Wie-r��Z�#�w6'�S�2�_L�+������,��+�RS�(�j���wدC	�t�Z�/il�JAN�z��Y�+,�z�����<Rj�:����{F��xb{0���͸�����X�6�9J�R:�H6)��6��*�L��橈9�3Ά���m���&����fQ��;���-�=�l��{��?�\wN��Y�RV�*�a�ݠ�	���e�n�P�F!���Nn�wI+Uw|9�v<�t��n��]l0�,"qEE9؂�j�x�[�љ6���q�%�̒��v�����/��<t]�!���V��u�x8E>陙O�u�M5v�,�H���-]�\�v��Sc}�7'оl��k*n��b�[��V��X��������2�N�_l]�w�����]�'�f�t"V(����7o.4-%Ң��g%";��Z	��T�-:�j]ub͝�Л5�S�����n�C�M�2)�9�m���1YM�_88��[�+;�-��E,F�9*�����XA�{�@+yb��W�'��u)r�O�9s��/FT
<9u�;Q�-o^& `Ӫ%]Ch�^��X� 4�[�����۸�;������n���9�*��'>{���0Y׷�-��l��N�{�R�%�$�nn��+���*�Cz�A�*�J��c(�z)��xt��F[փZ�I�YܵvGMU����`8��0�b�l�u6�u�ӝ�{Z�fwY�ELPS��ʎL�MI�ݭ�&ɫeeÐ�J��N�S�����=t���I�0��ڄ�*��h��Bh�{Lp*�5���4�xث2f"�tC+�9�)�që������9wFJ��h������SY)������Y�m7X�q����I�ke��@��P�=C&�xuT�=Bwό�H3��������;�c���t�43b���������W[l����
ȝ��3;R�eJ6U��@3�Dr�ł��1}i��n�l�hwvTb��Xy䃫q�:�X1�<Z�v�7]��WT�xn.�w@j���>���O��Q�VVJ}��L��e�0�r˫�,c�o��x�r�z��{([�`����zy9���է�QX6h3�耖�+�Y��U�ۇ�;�]MJ���Dꣃi�P����>����N&.��/hNW-�����'u
�j�r���]e'��Q5�ĴMθ�h0��x7+H�����D);�26�L	����7��䵪
\2�ɵ�c�Ԉ �;=��K�Ӧ���@ԭv��O&�}�o�m�twf�;�8�tY� �RuQz��9���`�H�G�ǚ�2��B�/���@�W�Bݬ86��a���	A5�&����鵒�`�Ll�4	�Z� V.B��\:��%��׿����|-B]��uC`�v��D�73:_���YJ�[`��%ʤU��x���n2z����!�p��d�Φ�]fJOg65�0�h��&!qUϡ�`���Q������':߭���1=�7��̖��b����R;0}M�Mބ��:쑏7h+�)W[s�LsbT�d��g$7�K Ɏӥk�V����k�V �s�V2�ӛۉ�a����s�%71��on��Vq� ���s�M��w;�s���s�k��̏��)3�1n�70��ʝt���&���5��9�bz�W�:����]�W`Ա��X��j���ӎ�޽B�H�	X���|S�Ƭ�{��}N��ے<�[��ʭi�S�EN��tf�z.�>J�}�\�R�˛]!�&-	�a)
mN/�8z%n¾ؙ�j��
���[������{\�{[��:.����0��|�|9[��^8���8�������!V3X�.p�]m��o� ��,�n�'f��w�^�\�ʘ�:*��X��v%��
t2�Z����'�LwGw��s��"��������DΎ�t��y�L���A��U�"� v��42`^A���m�%j�M5cwY2�bbݼB��������o&�r���m�KǓ�;�5��E��~��f��A�2�[&Z2H]�D�jo��ۧ!�9L`��EQ�֖�t�BOe���[��1��v�j�u�]��AT��K�s.�0�3l�ѶTԺ�¹�Ѝ.����x�*�4�ː̝�S܅�mma��f��'f��*Te��kU*�%�͝�Z{0��D� ��s�"�k�	8���7ûu����Y�m9��F��W֩�:=����Q]J=F��U�� R��),=N�)��4z�`�'mX�v�FP�����r]ҥv�R�A��e��V�4��
��z����9 j�����4|��i��.��kb�se9�V���y����6:GyXrU� ��B�}ڏI,X��B���i��R�ӭO�X��B�em�"��}[JFv�P�:�\��c���?onlN���ƣo�3��1�`̾�r���1
�LP��h��).8���z﫺vԤ2���h�ҽ�z|E���7x��2��Ȏ��gn�����L�46R�*v��
�=9ݗ�lR�|��=�2�X a�w�*���,��a��@��}�p���]�����0na�T��i�۠ƛ�L9���� Su
�' Y���'�'���c}�6��:aįfoG3Q���
�����A�x�4���,<�֏K4�s���\�����\�/���qa�;dD�]�j�]Ln=v8m�r�_/��ڗ[u�z%�^l�eg+&�⠇<w�+�駥�CF"뫉&h��ʾ��^�ثK,��u�K��=�Сz]��s+������j
�XTx����	e��]P���u����]�ZxT�4JB��Q0yO]EECj��%��ܾA؋Y�
p��m4�0����t�ǵ/{�	�(��V&P�u�c؏.�k;HDd�C;��Pd7���m�b�R���'�����Ӫ4�<�M���{h�l�j�	"�-��q�H���k�x.L]8�u�1Nw� �R�bu.n)��c�Z�aV�%�|�Q�.S.�ݙ�b���$�Q*2�O��hE�{Ҕ��:���{C/���Q��]�/vP�T��rɻI���V�W��JL��MEG�x�6�J[�b)�M�z��OG�`��ݷO7L�oT��9�\h9}����՜�h.�M�e�廝�P�$_/�V���p�Z�hvW �j����W��J� t)��fR���[��U�ˏY��p��/��|��.�DN0(Y�2s7�H��~S {Zj]�T�Xrn��|�qشN�VM<ޚ�L�o�y@X�fJ��}��dd$�8�f�U�9�β��'D�i=�IN�9��B��{�W �Aʒ��N��:�hڲ�Ӭ��H���w��}w���.����=���.���Z\����t��,#=�O]ni ˭X�)Ko��D���e)k���̉g>�
K�J��P��[�o����+�J�3���Re�ścC"vk^Kce�ӣۂtHpg��Mv���ebb��fp�vvt�V_J�D��`����nm��`�7Q�t�1�_\�iben��tkw�N+q�v�O;;s��J2'��9��Y�h�/����8ќ��Vh��4�V.'t���r���@�6�Y1euL���հ~K�(@ͨ0�J���R�tt����1ܜt��L�|�!���Y�y7��;�'Y�kQ>�k�2��s!	�;�����%�V��/y�*�0+��"�b�U���#uj��ݝ.�;�y�9�[lN(mt3N_`0N)�|�Y��n�ܨ�N�ֵ>
�]c�[�u�ZD9oc�-c߳4�3�h����r+��#Si�r,/D�vEned�;!�2�iJP�[(Ȏǿ.Z�c�P��]�Q��n�����Ǻst\�!�'N>�*\{cW+�E�C�S�g�I=VVڬ4�M��붱_1�����;����h���o�L�̡ö��ޖwS�[%)��u�-�����/� 4O�S��n�K��=J��f�L�,�pH�e0�={����`}�3���Ȱ��]]��@��:m{=_����4<z6��g��;�������� ������b���Jܛ�z�.x�
��W!������p���"�N���n�ąnՍ0<ެ��kX!�ͩc�D�K����sy��-ɝ���QJ�t��4��ug.Y�gܺ�ǧm;9V�	�WD����F �r��4�-5D�4�t+qa��C�b���f0�q��!IُF=T�/�,��6ݙ�$�k�nZ�Rغ�BnX��0Vu,��p�z1�6�)�;6�fj�����[�w{���q�n�tE�\��VI���s��Q�w�Q��Yh�E� � �a����٥�{j��\;6B��Sx��f�dw>�m�Jj�X7�f,��P��-!^.���q�c�&���Ýo�4G�L�>�rY�{�<Kb�ټ�e�`,��]�Є�b�m�L�&�"r��+�$���@��%��y�g\8��[����If�Z��*r�\Wi�}���;�[I�Q�46w��a�τ��b��P�(��R�e2����e��G�.�|xv[��
��$��n2�&i��qe�JjXzX�I��ꇆ�1� ����D]�unim��EKc�6�>X�:��� ���w��r��c��:9�V���U�pB��m
��"ݼ}q���)M��n=�8%�hi��!tX�ejg�}I��Ne��vGSf�A�o/�
�'�*��I|�r���٭rƊ{1vWC�PL��t���l{�r�U�-�.a�=�������8���7{ �,�����o%ԍN�hu���V�n�������I���a�u4-ub�#SNJLжU�L>V�CI����oX��(y5��,���ޝ1 �	=���[�{��Mw@�R�hǴ;���Ph��SŮ����©��2n�=BI��(�:���Z�WZ�u�x9�']G�-R����*JnS�J�uM&��.��d�J��<�B!W2�j�#5*](8A�Kp�C5� �Z]���0�.���Y��s��}�v0>��m'�{��˷x�ݛ�L�;A�L4qՇk���;in��dm���	��BD�fҵ7UYԩ��w4��a���:�ql{��g3)�-���;�XY���1E���u���������o��B�v	�s\/6�\�ͭM�X{+��f��r��vT�ˠBao�klC������y�[�.a�Ѻ �ِ�t���Õ�u�}4�4�t�Bzs8Ӱ5x<T�ʷ��n2�]SO����d�����|pC��1��}[P^�1�}��u0�ޭ
w.D����K��e�rb�WbVN��`�A������*�m�{RcPL��3��@��_w� ��lBEP� ut�k[d� �.壱����
�V1}͵�fуꃐ�P�`q��l�oR��*F�q��ܔot	�'Gzd���i��V�V�uu��3!�hۀ���7�4X.�\n�
�vP�p�,�}%���gCDf��C�Wfz~�N�4"x�@.�=��ѱb
��QP��yI���*lLU�� �=�VZ�u����z�-�P; ����̨�Ԡ��A˗��}%�N.h��H`�͕�Qm�eHzr�A/�ƹaӏMJ82��B7F�s��l�܀�炛�ZX�{"C�nX��8n�D�r("05�[Aw:�WM抝s����Vά��*r�3&Z8��I����:�a�����^��
ά��6^�|���ˍ��k��ЎB2�v9��jƾǅMͷM�9W͝�9k炎]�ML஁�r��:�S8U��'�6�囷��erKO*�*�ͤL<�ɧyf+#�D�+|���ˤ�:�VEΣKtrn�*VsW Z#�<�uW���X�7ADRН)j�nS�M���k���GغV��fo.O��O� �i���b3tqK��:L*�[���b�8�t����Kx��3��F�Ƕ��BWw�{�@w8rЦ3����t���ú�Ӝ
ҁY����ͅ�a���;��*t^�:=�SƮ�bܝT�����:�"MG#�Ql��֕��w;+S媶��|uS}M��J��,Ppv{3:���)�u�k�i�ǎ�,<ꯍ�]`��1о� ��=\J��-�w����	,	���w�'L﷨Ig� �V���`'��<_T�U����)R��ts8���J�f�f�[��:���lWV����Pf�zq���<:�^Jf�ԗ��&ogWsd�l�K�-�B4%13#���E�� ��9K��;h���7�3e��5�B��`���p�5�Xc�v/7)P)���ޮ�����t��/z��¬�'��3��og;�wZf2z���:�Tt�1�w[s�'"D�ك9��vh��dGQ��9'��e�O>�cs��X�'�����Z�	)�j�Q������b�V��#��jP)t���=�Y�{�})EG�'Y�x��o�wd��ܡ�n�"�=YY��+<z8\�\�G�>/']��L�kn�����"�\�DҶC�՛z��1����9m^�0tJ�&�6�s��݋^�o���E�\���I�b�q���r`��J�;�J����A(�3V�������/eGm�f��c`��"�O*�/lյ@��9��!�`N��+y;�ݍ���V�!KY�uݜ�K�ٗ�f8"f�5��wK������T�2i����m\( z�VmC�.��u6]�b�Y!z�����)�b�1jm��9����Μ}\
�G��c�^��y9F�Ш5]���ö�=�q�(n�6t�\�N��v��H���\le�nn<�� %�d�O	��uxtl@����x���&��x�WV��6�0�ѓ�]f�.��􄶀\������3-��5�^5G��&j�h7�}Őu��*�K����J�S��n}�^*�ʛ���ԑq҃)X��w��}���u�ևC�!`]4'�{KX�$GY���|Ηʇ=�t�� �JϓV[���
�.��n��MP�,}-��ܠ-����[]sVP�qƀ9��--�{���Wx�T�MU��u�ٸ7S�����k(��N�����P=Ѥ6���{��0up�Z��h���Yx,����Q=�ˎT,�GǴ��[�WY�.��@'�b�]Z���;��J��6.Xͩ����޹ػ쬅*Ug^�L���ԉ m��)���8�"�{d�Ý�]�71l4���%ʻ���e��u�sd{�;`<ڹWƋ����[ҳ�t�Lly0f�.�u;������/�\�*+=)Q�즗L5.M�j�`�.�+�޴�u��l�$Ғ%[,��]k29�2��us[��#߇uu��͙�v��a����`^,��h�.���,>Xթkv)I�ξn�:w>loM6�u�`�*stK6�&5==�+=]��*z�h��Ġ�]g.9��8�-�|嬉VC�C����u���՚s7V�J�u��҂w��u0���hK8,z��Z��[��X��Bx�e�u׫�!6awm�]G\�G;�J���Q١Y5�kX�Z��LB����j�}Ӧ�h�#.����t��F<�ҕf�{]B�9����@�PPj,���u�	�N����I
t�e0FˤUn��8^p$j����Eʴ+	��ÝMq�A�����Ig]�nG�R�uvN��vS���Q��j���+Ui\�KED,���cx�n�/am��4�;
����Wr�V�ۍ�]ѵ����.�-���F��F{n�i&uCN�e,�t����M�d�ܱo��=���e ����L�
��hA1�n�#���r³���) ����r�� ^��e�m��EP�(�J�v�u��Һr5��1��6��	ԍ���G
O/�1���Z���g��H��^q�M��_n�+�m��*u�����О�*�c�US%N�p)M]���v���\�<��n��ձISC��k�\�{��ko\�٪�U���y�-�2���ۄ�xK�L�V�:� 6+�XXսI_41.�4�*|뱄6�y����+/7�s=�M��`⸍\�����]A^.'vE�Hrѻ���w4VE\�E��D+Q}���]]Yx,S,
��ٰ-	�ܪ��/�t���[��\��܃UJBJ�!�����;)�9��f�����r�j����
�.�����T�v�����P���C�^����4֪{ٲ��Y�V�[֬��Fu�����pܾ�Ft���N>�9L��7	qs���Y��4��|6!��ʺ��'.�����'_cvn��-(�:��֜��{6P��d����LSj�F����Y�}Ǖ��"�`�c�h����9p>��j��lCّ?�FJ�dv��O��Mx+3d��NY�|�/�F�uX���m��J+&8�0��W�]J�Qg{F!����ܭ38�8���SX�����q�Ia/lڡ5	�*�|�A�32Q۸@����N��8 )� v똨�����qn�w�M���YB\JN��)�Bʰ��FZU���U�$��bUi�Z�;r�)��;�ޙF*���j�M|�dÖ�d���g^�,П��X�-.��}u�7�^�G�`��<�F���]�����6��u��	���$+�gOs����<s7`(MfEbRO�CSo���,�\Z͜4z�!d��ZYh:&)�8q�o[HV�q%m5�(��0۝�iSˮ�8��[O/�,�䰍I��]>V�BRf�ٸ(�R/v�����sa�L�_U�lj_q�G��Z�J(�;v��;���D��re�9\��S�� ���sr�jv�b��sQ�8mr-pW3�Yu���+Mw>���ggL]ԃ�̰��s�3���΃�޹c�8�V�����\	{x��|�h�H���e�1r�7E*��b2I	�yx�ʵ(.��v:�'lD�8���VŜi�"�+sE;c:�x3���@<���Op���y��������,e�o!�!|����K�H�t��-#qel�{�P���}-����[����[B���O�R�֮}OAY& 3#���0[�n�R?N���w�݄��K���Ү���E�D�sv]���"�]H
��W��^�����¡P�TVK�,ᡄ����v:ae%�b�Pu�=!m�=&��iL��#<9N�݆AȦ�ة]��gY������o(a�������v �L��L�����!�#�Ƌ=L�8�cnK���H���-��ee�uo[��79mJ�5h�u�V&��t� ���B���Y6v�6���Zt�L�� ����f�%�U������1H����Յ�z��k���M�OtD��D�,^,�����|t���2�B�mwu+&h�w]��[c��t�sųp�ĩ�Z�x��â�&��1����꿻��;�w�/sC�|`��m�}8Ղ��O!�j�.o|��ԁ�I^	�DQ�9�^r{e1\_j�:����ZR�<5��
1)�E���H��2��:�E��fkd�»]��b�w�3��'v��0-�Յ�QE�2w�MB�S1[)9�v�
Ω�fq�Y*�'�؆QR��SG]��V�귢1�۶�c�!���ԁh�Bp���Δ���v�=QAWw�wc���я���n�F[�`PP��ӧY87�� � �%{ۮ�܋�<�^`U#Yٴ�[d�	�%ʕ�j���e:y�5}p�K�Nf��+��w!tj�b�k���-WX`��n��B�س+����"0ٱu��-h$Ms�z%,���˾n��P��B>�OjO1Y�.Z�IZ��3C����ש#����w˗�˳�'@p����bc+sz��e`#�1�3�wQ[�$E��$�Z:k���^wYYC�4q�RO�8bS��7�7�	�V�e1)�4��ti��uz�L�*�������R
�rD+*�^��ä��fɮ�	��%8H���ñm!Ǧd���Z)kާ�x��Fʏ6:�c�;��5.	��5[&�͓���UeE�M&����Մ�Y1GO&v�$	nk;8mǋ������a���r�{�3ƙ�u�\n���!h[�!]XSL�[5%�����^T�}����ټn���GR��Wv��5Xۙ� ���T��%7�Z�S
����J�/*���?Cr^VP���1���▨�z* �+n"�s��D����2�]@�Sݺ���v)˃U������ksj8�+x68E䊇|��8L�sE����xA-�e��f��1�����2�R��$f�
4 ��:�tJwo�O+�����<DoX}�o��Xĸ�L��2m�R�.���{o��=Y�6IϸP��B�:�ti�Y��s��d����YӤ�W�����ҩ�w�y�cpu����W>��|����Ej�{���Y4�]&�r�nk���(x�����Q�u@�,�pk`�:⫒r�Y\��E}��lWø�'3��m�Elt�Q�-��e����:�"��q��2뱛�wgd�9g����E���^In�F���Gm��w_#���/����vj��^�v9����w�h�����0���f��U��_Q���]�ʅ��]>��]�I��0IVi���e�w��S��3�k!����c�^���N���-LB��݁�^�P �����B>np�ή��Q�K"�����!-�F�s���9 ���us��Y���B�ϕE�ehj�廬.�yM���Y'�ڣM��w�K^��vX]HR�o8�ˉA�>e���c{B뤑�1.�b0��P4�:]Y�iͰWT�K}4m!��z��+fY�4�.�M��C�iy��x�����'A�J[���8��[�
�p\jd����*�:A,��h�t.�-���j���Y�6&�4c���(�:��x�p̮��#\H9�×ͦ7`�6������S��)�̺p>Ճ0L�6�sS��l���9�:��A�d ;�n�
�-�B�p���Y\��
*Gwx�t�����Y����X������=P3v�d��] �X�Cvb�V`�&��I��T�5yM�VXj�!���ƇN���+����c��ެ+E��d��im�Y��N���;ѣ8b��u�B�' �����VG��=92��yN�./R��H��CvN�Yx�rT)��bPw((�8�+Z��Փ5�/���V�;��qqY]��J���$b(b�g��W_w��.��/�re6{T��$J��j�[��)�5U��O�oU�q�Z�py1p�I���w��#hB�T%�:z��n]M�g"4	�^��i�ʶvw�V����t6oQZ*��}�._�W�_}U�}��﷚�j�,�u�X|ۧ��Y���{�N��/e��Q�]i��][�Yt���٪	�	����%�<�Y�S�.����>��؍:������⛸�-P���-׳�E���)h�P�{F�켻���g��ը7W90�[�Q/�vWge#Jfؽ�ˢ$�#0o#�U��B����%a-�-�V�0C�A�֕s"Wf�O=GeE������+�I��fj<�Δ��w�/�|{��IۚX��Yڬ�ה[4�ϡMc���|�5�;3�2�Y<�O�o=�4���]Uz��<���7U�g�i\)����(��Յ���)[7�^n���4�+���1$Ci0)��wgR�]�45�ƹŜ�zݛ7����<LkS㩛�n)���DAFٝ�jq�ʧv�7#T4^�X��R��]\���F�@���z���Ӣ�W*���T{���oO��TW}i�h8��� K���l��S��V/
�P�Ჯc2f�]�f�Ϋ�,N��=sGP�4���_}��6���S'[��M{�;;��᷽�"T [���b�j��[e�R���;)ݛ��u+�ܥ��yZԷM�d��!n^�س�����������\r�C�	^ͦ�Yg*������C)^��J��-[TH���-���I%��na���=�Wr����xƞ]��u���!:��oA���ͪ��m%����\��o�ֳK����tԫ�MTR��1-2�T" �RQ��lfU�BUd�(��;t)�*̈�FI^��� �J(�4"��Ҕ�J�#0��0̪
T�

r�"��BJ�Y��R(d"���CWZ�*ܠ�*ID��&AnD�y����Y.�T�e[�����T�Mg�^[Y�� K9�)"�&�^�(�DTvۄk�^�QT^��QY D��Έy��մ���Qh���xY��TET�7T���l�QbTA��F���j�zaPQk��^�jD��W1tR
���%]"�<���,�45<�Qu��=�B�,�E<�]T�]S
���B\�	4�/5�ȯSu$�+=L�%#$ə0�	�tQ�)@��+�r�R]<��" 	����u��� w �}�we���s�5fu��rڊ�MwǕa�3����޼�D�P�i��:։D�Y�p6�N�ˬ0��ޥ/ue
"����@�/�4~��환����u���T�P��R�#"�E+�{��4����%���DP�tW�1�-����ݕ��Ȇ�4T2^L�6���Р��S�N� w��뀬�V�'nQ\+�/�"�͎R޵{E˂�a���vv���|ـ�3��-y�(�� u���vV���~���ny���=Шh��H����J�0G=��ԝ5�ܫmm�1s�H�5��
Wot��nv��t��i���� +Φ? �:rE�'���N�m�oW�*�`]��ߍ>���]�\�ǰD*�ߍ��-�ٿ��+\����'L��b���w�%�Ew5)���u�u�PA�v���H���IxY�>gG���|����fK,r1���ǆ :7��h�����bE�J�y4f��&	A�(
�H<!��a3/�e�˵B[�ٴ�Jya.'kF����2�ד)�3�;- ���
�K�T�o�ܝ^�N�;�xV@*1"QX�GB����ip�tW�<�|}�`97��T|��8�܅�(��G�s7��u�Z��,Z������9&��8
�+1F�=�nReuK:��#{H.v�/���Ó����&����70r3�+��I�Q��X���G\$�|x�lt��n_�j��}sF�*N�v@��9NVv�Gj�V:k��dƄM���D.�"U��B��^��ӹ`���1�ٯ�W�ڢ�
T�m�_vLȋ1�����_R�O3Bo#R���G^�TE��}<�'�Z]��p*�@�% �!W�!#?WM
+i�ωH��B5��Q]�ȩ��dK�}��ʸ�v~�ـ
u?FC��j1.)�h��:>+�Y�»�t����Uh%3ʘ��u��79LҮ}��Yz�{ŀk�{�%��QU�v(�S�Ds�[g��S��g�і�;�;���1�&%L��g秢U�I'#�'��<�7k�xO�t�m�)c�&��u殺p�5X�b�;�iՒŇ!N����P�m��M�+X�Æ�_tp�gXO2<Ԣ��<a{����HW��7����ۄ \Xc���`��(H�������6j��	���]�%,u�2��}xb�Gl�zw��a�Y7	�!ŝ[L�t�R��SC����O}��1h��e��e�Uw�͏d�N�b�,�����K��NI"j=M���3y����������/�gd��o�/�lHx��2Dw O^gu�����	��:��J���	�X\K,ӳ��05żǘ����."�����:L(�����y�(Ç�m�a}�Ҷup�@� P�y���4��<g���V�Vϭ{���*����۶��F*T�?kӨ���������Y��7N��8- s�Yx:��®2g\�Ya��O�Z�6j�U��^m��.v��{I��E���޾�Om��
��K\�9)� �oR���.�{ݓn�ȱ!�ʩJr#jx3������K���ꌴ��?\d�!��+)ܾ|�b�[�ge�Uh/�'0��G1Ҹ��:e��%i���zT��C�E)��p�3ju��z��U��W r�`����~B�q��σ��_QLn�Vw�� �����# iT�A��<z��*����~���j"�q{���_@���)�2����x�ٻ���T�wS�^�W�|z!��@�.Txs��G��ԡ\6�,�gV��O[δ�K�W*��]n��1�8WźVC� L)D�5&��O/���}�쩍O{h!��}�W(?�]-1��h�I���[��p'3q�#���|����I\WBaE:�9X�94嫛
��u9�1C�x�b������AGD4��X6��U���k�\��j�T>��e$pi^��+#t-���T߭�9��!M����hb���
\X����������{R|�~Y �����>�[}y�P�1'Vʇ.�����0�*�V.�^wzb�|dy P|���J:ݵ�~��r�
��<0N��F�mP�Y�W3]kz��/��9�� � ?�t�1_�噱���¼��l�G70��o2ئ�]dV�	�z��|�e�R\g��TN|����˙aa"���a�����C�f��Bg{�їoe���	>���؇�Yhj�N7'�D����6x2b�@c�T�!�4#�fS�9_s���:%�܂Q1P2)US��������sh�[���{yr���m1[�Cpuף��,A���١!�ytP.�B�2f8F2�\��f�b �x��s�n�����F;.L`OIW���4q�s@�"�s�f��X�q��+��B1it��c��wL2��P<��#VrɽM��'ٴ�l�Aj#������π�{{$�d��奇��2T�K17[�6��\CP��#�Uy͜/��+' �+ �(� �*���ʘ:}�8�D�F
O���F���N6���q�W%��ޤ��9��a]�t��x(U�����7y����n��.5 ~��7��|�"��桠��.�sh��)����hL I�S��1�{�) ���M��֋z��仹�=�!�Fa�gEIP�vnE�\�K��	��|>��:���v��Q� F����u#
� C�x�a��2;��ԫus������5��F29®g#O�)�!l
�'��=��LO�]�����+K�X�>ܜ�vh��\wA�-l��=W�Ә�x_��qS���5�TF"��b'�U���.~^�+�Օ��*��33�S_"��ȍj�!o��PvX=p��	­c�y��x��oe�(�p.���!�+Nϒ���>׌��U�u��
u[��ᾫdl���9��RW�Q|�4[8,��Y	� a�7����^QnvOiZ]�s&�}/mf�vU�N�oY�o��wU�|:�&~��v�¼��忹�W�b�C��
�u��.Gz(`�2������\G9����T�on��yG�� �$.1�rPpX�*6��H��q�/�ck�{�ƣ���B�_��58�����!3dz�ʹ{̆*z�A�+�軽�u��s�ɋ�UBg��p0N�t;��`T)�"��B�Z6��_��l�,T�V���}:2�T�/u���.�#��bL�ͺ��0����o�q9Cg�?qެX�㙜���f嵧�f�WS��-7C3����Ɂ-�"L����<l��n���f:#�����:�o��ɦ(ܝ+,�B��KY{����p�=Uv�ϑ�=��@���[��q�(�>�t~�N�8�[;��׼ �+v_iVdt'[�=u�[.Z�оz�ixY�����������cx�#�Ցu.7��i�PL+��'=Ձi�j�����cg��٪�Z ��_Q<4�7�*����xW�{iV��'�<�7����_^	�R��l�V�����M���Zit�^t� ZNb��Vw6�o5U�<7yrl���T�pӿ��h����m��p���|�]>��#
�Z��̺g�-�9x�� n��Ǝ&�"�mNpPq��ϳ�:;N㑅�uR�N9�,=���\���v��x}8�I��;��o�c���[pz�\p���q���#j���<����y�yFU|�yx��u!#\d����2��߄���}�*���{�����T��U��[l�ր+�H�K�#).)�<<Ώ�.Yf�
�	 �.�ɽ3G��,i="O�M����]0�As��9����Y�QU�v(�S�Dv��Y�e䋲z�6�
w�<RԐ�y��_#C���f��w�=�K{Z\Ke灝i7��`�L�CLש`۳d*'Nh�ԩy�P���5ڇ�*��{O �v]_S��a��):�+8t�43��5�{Xk^wQu؃�!Ս��YfS�!�t��\��c�rb�W�wv]�uu_\���,63O�>�T��Hc��p�3s����W@>�Sd�D���Lhc�<���	5|�/eFe��a�wt���%��9
b��R"����tA�p�V+w��e��`�\I�:v~��0��zk5�90��S2J�=� ٍ�{��9�>
;((�!����}���ǵ��o�e+�w���7��0K,��0A�.y��[I<����1Ѳ�fr�؍�tO	��-k5,�U	$�g{ue�t,����Մ����M�ш�9�}���yX��".���+����Z��v�&{\�i��51�x@�?[�s�����3w����Q�p"�w�y@p\����]�u��}v�5��/�ۮ>����d�~���4w^;bx��7�Y�Ȃ"Vm؜ך�yx�2,}8n]V�5;œa�r�ȧ�'h1ıcqĽ1m���\��jJ�IoA]�*єX�f6�rM|LF��� ���Ȍ<�ܝpV���"��z�H�}W�)k�xpwK�.��-
iI/��`�ݚ�o�-�OBN���i��aJ�;����������e/�e���՚��5��8�^�W�HP�w����&Ǖ:�N�3��^\n�t�TS�%�Ӂ'cv9±�h>���H�쁁r��`�鯉A,�p=ch�A櫡���ͼ�ym��;=Ϟ-�q��ŏ�߈�]OR��M�J�%Dk�;���W1 "���ϲ4��$C�����=�/N���n�qVgJd3#�7#
�ǖEB�RQ7&4q��D ���`Wa�]Ӛ��/�x�4h�.^���2�'�;>,*sܹ��b:~�� :��x�{s�g��P�����+ϣn||q�[&VZ����p�[#�~�I:�rT����L�p��Æ��p��e��XZ�/a�J:�[��;&�sis�*c|��B�EQ�3�%�Y{��/gz��J�.�xFMౢ <����3ٻP���|w�p�>/k�B�����:��]�.5j{C���9<>��UC�(���˙aa�0�צë����}�)��_=Y�T��UKi��(����:jg_��0�qd�
�1�+��CP0�����-��K�t�7�ryo��S������Sɴt���-Z����N��Y2������Wm�b���f�q'@P �p��k[<-�,K�R�N��7A�8
5��Y#��q#/p�R^��%]�0����
�=�1�q�;�z���[r�:�=�>��\6�ޮ�-n�-���s�����R��#��v���ssXxa0�Z Z�wC\j�b ��}�r{���_"����l�Ҷ���L8��+�Ę�L6pu,�E�m��΅F2ֻ\s�Ρ��0���H�K�x�c�ʻ���\;`�=XJnk�3����ȭ���J}R4婅u�vT�w+-������Y��}Lp��-M�+erk����Ƽ*��<��So�<�N��-R���Y��@��P�"鳑��7M�9B)�;b�鐏TpG���1NP�貲���z�����1*l@������<4m}��F9e�X�P�C%I�fqp����=>��I��>^��E��c�^�k����_O9�G�y<T��#K���i^q�&�IkJ�Y2��غD���2���gC�n�,oҦ���o����[�->r���}v�R%B���PR��ä��rx*T�^3*�Uxn�WZ"������V�m�)�:�55���WnY��X�Sx,�NH�0a�ꢾ�[#_��n���F[|l�n�!֓~���L�v��8s�kӻVWb���m��s,9Z;�;��qc�e��J�����Cz�"S��.hU�n�֦�ֺ�f7n�*n���
���xB�w]ũ8^Eu�X��5^qs'�mҮ�F�ݮ����qZz��J0Y����V��]���#z��`y�Def�����%���+����(C�W��[�	8}d�yLn7:��,�������>O3>��0��fp�7�p�<���4�+�fJ)([��A�3��{�9e�W����:���R�Wt�ׅ�����M�ɡ4�Y��3�~h�nn���< -�#V-ҷ^�w��Z��y,	��M��i��hۑuɮkZ�9�Ե��#2��o+S?PϬ��V�l�������x�2J6WlVW1Ԝ���e�~i{Al�r�w=꼺M3�^?�H��'�8���t����^?jݹ�ӣSxw��};:u�\*wL'	+|r>�<�_=5�P�o�W����� /]B]��ȬF·�S�j�����H�D�V���L��cE#\c/U@G��x� C�UF��iux���;d�d��T,���'5Kg;s�y�M:�"4؎����D�����9�����ٞ�1��Y�V�.�"a[�.9�k��q��7�Wưm�w��0������{X2ڳK�mP
�B��FH���5p��1�gk��LS��� M�}�Z�u�W}�O�H��������V*�]t�N{���Gj�"�z�j�ZZ܈���' :v�Y�cE�t�v��5��2��7cpr9uur����.j���ؙf�5���땰k<3��̳�����˽���w�U��v.���r���J����d.}��I��%tm�W,�g{�:�
�1f�������&�\�]�dtm�ˏ:�О�u.�sr'(���Q��1,��LެV�������m�e$#UgN=T�O��nڬ��N����e��$�}DcKE�q�[YZ:�3�a=��]���Q��8���xP�]k5�1�Fj0 u3Fg;+ ˾�X�"����\U;��U�(��a��-<��$��8�kڳ���v,
TbN�ئX����[Y
��ϏW.؞q�/v���e����U��� �Y�$�u
g��]��V�=���UۚFB�u�ͮ���Tˤ�obATx�+H��F�%7� \���pvќ;��w�n��G�b논�s�?�m��C9Y�L���N2aT�0�����N�UF{;E��]��
TI��]��5v���i�7�[�C2<��w5���G��pJ��<xV;��gs��㲅EQg:�B�cDΒ�<�t��ɶ"��f,x3.WEv��V���zĖ�Q�-C|����כ-�`F����r0���}�M��Q�.�?lʑ��z[ߌ.�%%��G	�A^Ŷv*���I�ξ�8���eN���w��I��p�2���=��pޥY��(N�X�A���	�����n��YM���\<�Vk�kg/)XӓK�����1���2��N��:��a���>��8u�����ӮV*�16���2L���̃��`7py�]���.=b�sH���Q澦F,������K�͊��U�8�4E��K'V��ч� ���[�ػ�8�q�Y`(VL˻ދ��R�{�t9]m��T�F ����1�����9Qzr�*�3]��A�wMH�\��[�����5�sӑ�Ǐ�,I�u2���s��ۃrh�Ɯ}s��rY�tأH�%ô�t)���"SU*�]�/������Rut��3(s�V��͔�E[�f\jGX�m���`Gd�×uiտ���R��+�ۆ�޴����C۵��J�=Ȩ'�WQ�}c;�P�SK�4�yP=ӏl"Q��ui4������b×V,;(��C�[�M�R�|fG�����Px���<v8ͨxf����hc��7��@����1�Z���ghr����W���q�������i^
�z���L4��ɚ���(9�v��A�]l����ːhUx�Qj��4�HJ�&j5����=�8��#j��]���$b��-�6&�̼q�tX|�X�螼}ݕ������K]��P�wQ\E4T��5�����e=2��4�*BWTıC2�I,D<�B*2�qWRK@�D/r+=���4�r.�ٞ�&y�U��� W���^�Q^yUVzz�d�j�QG�yy��jDG�I��D^�RI&a�$��YP���x�aJ��EJ!�v�^̢�4�H�<��
�=W<��
�u�Ġ�+	B�J�(�/)1R�H��˱(9^Rnf�n��	&(I��IDF��`k�V�z�J��[��b�QVa��QQQAI��G��)H!�R.�D�n^�H��i�R/+R�U]�� BD� �]*%3KȨ����J��J��Đ��KC�/35Ң�0�"�� ���\�(�Q"3#ȯ*�7Q=!<f{Up�\"�#��K\�Q��̉CY	EM]G�����/<�
*~�SM!]
�� x >@� >gtdy�K��o-�ɸo�%�)�6\� 	PWv�n��#x�E,��ɷ��ǯ�#w�z�&��%��Es��Q[Gz���ppٹ/[�>>��:��|�Y���b�晄����DI׌�u���Æ!��h3FY�KH.K���N��-��j�Ryn�	u���ޕ�IHJL���z�d�7�V>ŏ���j�T�Ht"��"$2�e
f�+ǳ�02�2S3�\:۔��"u��<�ЫI��[��q��)���<�%���-�C��>O���yH*�̦�߫��^����ʕ,�#7�'`��{�b"�}h=�ٔu�Kd�~��R|�%�I�z���)��J�׵�2�Ц�ᇸ�8�B�l��<d�~��%�����)X�+�c�l���}~t|6��~I��H���`�$�-�W�@�q'ͳ���Pa �OQ�a'��Nc���%��-��nO�,��g]Փ.�Zɓ�-YI+�Kf%�����F�+L�@�P�>/�&k��f�T�{i�,��DX���RM>��q��Հ��`�C/�<��O��Ʉ<�����\��i�a���>�[�a ������l�;�I����U�`2�ail4βж��"�s`U��wz����g�"@m�&��e��m5��Vm% q35�����%�wvB��%]R9ˆu
|����������,)��{�&|�T����ʰ ��B�,E�顡�,�Y{�;��x�[%6��۩��a�m-b�l�e��h��H*�ə��M�i��a����3��<�I�)-��E'P�¾�q����Riz~��X�~��"|����]j�m'37��s��@���Mg,�%$��kS0��>��1t$�L-C�8�M��$u&�xn��Pe �3��|�I��A��a�-�!��z@�S%2��{�ty�k߳�t}׉-�B��y�	�g�W(���2�ZM2_�$��&{�bJi�d�9ZC	l�mY3tZN�N�<�����Jv�����$q���Ǩ�`����1IB��U<��6|J݇��V$��-�ܸi�Ho�w��<���4���3�Z|����^�
�����CI��\)Y�Jd��������/F,�Cm%]Rg%���%@����>;{}��9��:\�җ��x%�h˹ސ�cE%A��Y\ڔ��y�[�C�R3�ܥ�ڎ**�W�0�#$�V&ӄr]�K�ֹ�����q�D�x�2�n�r��u��A�����/wMp��A��yu&	YL�8GB�]�?�^]G�w�汞��C�V����������sY4��f���0�Ro��ɖaM�p�ה:��ө8��Z� [8�hh;�y$O�Rд���R� ��Z0'��Z�n�ǎz�}�I���	l�0���<f�i5ړ�5��RO��4_�N&ejβq$�jC��3L��\�X|>�Ɏ}���^)6J�60��z|�[����ZA}��KI�)D^2q-�L&sS(Jd�`�.|�%�ahZkt�ԕچa�ސ�Az�a]���Z�9e�y�m���~���}�#�
�VM\OK�����4��>�)������}��RS��Ɏф�ϝh�N�e��]�'ϓ3������Q��gZZIL�<�������$aX�y��A|�}�a������p���ٶVm%0��)hq%;M��h�JB��J�����O!L�^nL_l����T�aǎ2]βRN���*C	UN���
m���u��y�Z��=UsV�Ue�>�|����G��"4}i����2�P�����i�P�O�R�0�q�K����M�I�^�:ɤ�B�I��0��I8�*�aL)�*O&b���:��2j��Y�Jk�-��_ya�Q��Ý���C����W�R��W*M��h�؁�:�͡�}g�ɤ�̡�ş6�������䤜B�G�`a�M���S~�!�Jd�;��g\0넖�kB��%r���}6�z}�s7}Y1މ���K����DAz�'�����Z!�لY:�6�O.��0�d�l�۹�!N�fw�y4��L�M����&�FU�6�}�y�0�LQ-E'��M2��DE%�jwjIǬf�Z;W>��h[0���ؠ-�g��5��H,>L�T�(���א�+0������i$����UC	<�!�3/�Vh�$�罳̙�y�l�����>#��b�|������U���5���9�8��2RM3�oRR�\v����Sl�1D�C�Kr�H,�g�͇���SL<�C����[�a�
A|�!�w�i�I>B��`�L�I�)��3���.��aLb�aӯ��S�@q)k�X-*��jZ��],0b�:x�W�9:�gN���b�b�}��Uð��p�;NoZ��'%{�`�ޱ��q��tkz�T���{֢����q,�vd�V!��3Ӳ9_��3�I�%p�D�0DAλa�}R~�;�Hi% y)����,�JC��.�N2Յ!I:�n��SnX�y��M�8��$�����.aY8���k�9��{�R^|���} X�8DH�r�Ѷ@�S%�٧�-�N�RAV|����M!���6Ww�Re��%"�ƙ����R|ɦ������5A�˶!��q�w�3޻���yn���=���b��j�βW��p�&ϻ`aX��F3,�%4���\�'P�u�����2��-�a�H*�综C)hm@��/�B���ƀ�RICDW5~�G/ɭwk+}C��i��1h���z}A��0�fMV�J�m�n���d�P|��vɆy��q���T�B�G}xI��[0�� ZC�l=��|�H,��\�-6����B��aW=՝O6�j�v#�>"#I�-�T��% �o]LT%$�`�L�d��B�M�a��35��B�S
wڇy�!����ϻy|�H��)���C>�8�VnwVL1�����
��@��������
C�=;߱���KH)�n���$�h-��T-Y4����i���9ahJfw�2�,�Ԗ����H*Ρ����(ZAw����x}�����H�4U���x�̎�^�)Ф�,4�g�Pa'P�����+I�)�urRa�����L4ɎQ�L�T�u��D넷	X��ϙ�u��C�u'P�u�{��i>�>c�����OK���]���t����j�Ɛ�H*�����'P��[��!����@�RIO�X8ɤ�B���oI�`)>��L���e��%2�|��a��JCa�:�*O!J�ZǳU�}s��m�9�w��鄝L%����ܘ���KLv����Ag���<�!�����I�R'�^��0�
Af=�bL�y)&�vKx�i<��-��J��]C�a�0��T�-�*�_w�_W��}}�g|��Ihe%$��[�%"�I�U��!\�u��ߨIhW(;u>e;`Rgy�<�'S�i|�"��Rs��>�VM�0�g��2�^�h�ل:ᅠq+������g��3Wh�2b 8ؕr�~o�Zkm�2.�����ETtGےQ�J�`_s��E��m1#�����B�+��Z�`�n�M�od�]d^���9�
r�:S�[7��ނ����<��S�B5�B�h��L� 2"k�}��u��;Y��}�X���*��
�i��c�&P��E�O2_(6��˩:�E��3N��d�O!I��=��`)0·�k�O%�`Rk�y&2_h�
߮e2V�wX�N��>�,]�����G� |GLO4�3̔�f�KCi�Φ���a ���d5FS�Z�\��Ry�l�Ԗ���fӁ۰��Hy��z��:�i:�;�nu&uT�"�w��&W�N�-P��>���O�{��6��L>|o���-��%Py���%*�P��O��q5��i�Hu��j��Ra ����8�B�o�T�e!�|��0�^���M��|�צ��Qw�3|�tߣA� 8�����CI�̖��X[
aJ퓝�$���O3�o2RiIHg�L6�H����Ry
���d.��'P���m&.�R~����(D��,u)<����=佰9��Ǝ�o���I�i9���BՓiL��\�0�]��;�<�fL-G��d�S<�%�{x���AVh����Z����l����u��"��>�����!S��Y�z��A���˔m�7�m��7G\�u+C2����)�%�&�@[?+����H*ɣ�ف%>e�`W��e��2�!l�{��4�H,�5v�)hmB-�AA�F��j�m��06�Y���?!���Q-�Hm=t��%��3��IY�`)���u�̕x�я���RUT��e��2W��	�2�8�+���Ii�[#ݓ�P��AX�=����]
��&�|��9�����i- �w8�3y>B٣%�N2��d1���)3�-�~IhJVB��2Z�C)�+�;�sI<�0�3����aII���|�z�H����9���L��z�{TW�D{�����>�p�+��9�#�?�����\꧞C��k�?]�&�7��>��h�(�6��M�kE��n�7*��g�ty�_���=�|�d6��{�7{G�ɽɻ��}Ĭ@�:�b�{�G��n�L�ʬmJ�U���.�\=x�3���lDʵ|У|���:�Z��\�x"ˠ��{�Ӛz��� y#�A����lsn��:wrӬ%VH��f�x��}U_T8[���;5���OQ������1����������V _�A���/���Myd���}��f��#��O'Dp�{0��N�0V[<�qp�cEB5�2��P댐'���E��"�kM,Ŷ�v��pR�I��x1&d=����8�G|5���Q
���j���M���e�P	F8ȕF�쁽*�q7gY�Q����C~�m_��{N�06:�f[Cyh��ddL �]��`S3���������٢����
���hI�#R�ü�r�dڨY�E)Dn^����ܑ�
4�j:�B���tТ���%#��t헰�rwP�<��=ogV����ƣ��AwXg�ހ"�I!J=&�&P��p�����«n����g�Ϳ��g��7D$�}M�1q�"�䬠:��$�08�ai�=\��+x\�G]�ԟ7u�S�ED>���;acy��Y���٩W@;tI4k2�hci=~�.yFK�EX�}I�]eF_E�&������ud��U�jB�m9N�Y7.P"��fX��#�|�J�e����m�!�df`�5[�V§z�b�Ȳ��ц�'��m�b)$��ǶL?dwA.Tӻ����˚r޾�u�^�C0�����ڙ��ۋ6�,1!�x�+yvM�g#���w�R%ɻ;������3�oS�u}?����m��i�����Evk�+u�3���S���w_��!��=�=f�ȡ\��C�m3���ͯ*B������"]�'Ա�Y��?���<�	�ޙ|;gr�r.�O� ݞЀ� 8�XQ<�!��j�ᨆoL��rí�٦O	�>V�\��J�*g��hw.��J��K���<�؝�m�G^G�{�P������V,r�uÇ$Ό�;+��T�w=�go&uL\D�"�믲�v�����\tX�4�q��-8:�mI�Mg���IqK�[u,���7�C\<3���z:�wJ�V�g��q���b�o��t%��m�)}���n�?s�?;��P�a��o�MgM�,���h��2�Ύ�
�R=f�{�B���7e��W|Ϡ
cQ
gb	��a 
S��ei��]�� �ge�ۮFgF.=P�;���,swP��x�wMA(!�逑�f�3���K1T*�����Omm�5\b���.��7 G#���ݫ�jf� w90F��� ������.��@i泅�iޫjT���%�)��o[=�e^��M5WdW�'PM�Y����hd��`p�V�ǽ�Z'��ڴ��v��H����ީ��F�ws�U�8�4+.�t����z��ؤ��Q��#��br0f�[��>���8�rU�ZC�x����Ǝә�٨x����Ū�j��wDL)�'�R26�7)CN�ue]��t�'�*�q�/Mp��y��B2��N��2��('s7.b8��f��3�q�w�ޠ�����{O���.Y11K�$v�cw��c�H��N����Ԯ�n	n��p.N/�"&Ed�j�l�i����{��v�y�����j/%r�1�ƙ��:������P0U�2L!I��AYv�l@�9<b��r��|gט���v�������s<��譌�T$n��ca̖Q�X>н�%z�#�`{Ip�2����B�^7q�+���΍�9�*�7�,53�j���N��#į��Ơm��_5�p�dō��Qr��Z���H�n%V�����+�k��r5K�a���b<��t��*W���λ]�K����D����.��b�氡p2L1Q�W�X�R� �i���G�3�Ի��¼.zع��:����Aw�A�*���xBo�����ベ��:��L\j"�$ =��ƳOJw{�p�a�dEF�����+�;�x��5 ��&.��j7�`����쳔1����ߏV	R��8E^"�&l�Z.��Ρ�IYR�ѵ����
s��k�k�J$1Sz�K ������mf-3�}�6�=?}U��W�G�:Ӌ���N��v��W_`o����S�xw)T��Vy����<���]����lֺv�-�;J'K�U����<�s�cB��B�U������Ei$`�s�-���凶(C�8��1@�I��A�e����x��j��m�%]�K@���d�Ŝ�矪.�1@3=Oc��^�S����Jv��q������]P�C˺v`��x%ׯ���F|h��*_r���5���)B�a\=W��C��x[{\T��'�F�<:�*�"2��mX����t�=�b�[��|M*����=ƮB2����Q@2��K��us�[N�2�r�4�t؇��U�@+wpF|� �m ;�5>׌��^��Z|��"ԍ��mr�x����"��mu[8[�#�
 �o�I�1��g�6���7(i����Ǹ��y�X=������0ؘU�$�p�R�E���l�e�zr�eb��%fĚr��Y}܁���us��|p=&MGt��<����x[��p����(�e�@.���Mq�(wL�1km��D� /ˊlx�:M���ߍ����%K�� |D:UKJh�.
��u���G-M��S�p���6��B[���ک�78�$��	�#ʸ־�n��c�ď<��<�Vww=ۖ�FB��6��/n�UW�}_�%q#�uw�~������ŏ?���9|�
��p�Ҽ6��!�j���6��a�[�O��!�I���s6��+ޱ�*Z�[]zG��5��R>Φ)�#b���=Ri{��wH����z#�^�5z�U�ajg�f�n���P�!!2���k�<t����{�&��3ݮ�W{���[a|�����p������F��6����,�f7&2N�ڠ��.�e�N���-ȇ_n���������$Ē����:��}2�)���r.�i�u���1\i��Juad��p��e"эw��U@E$"p-"T��{�-�WH���S<�S���d�B+�RN�z�a����y�3�]��oF6��\l��%Q�����T�q9y��	,�nth���s���|�W3�[�5g�mD:wfc�ҔL�J⫨�t��1��y������EG�����U�����H�}Hq�@�Aҙ
Q��b��-������J��_���		QoȌ�W���c-�'�a�x3�+� �!AZo+�'��W�*��4&��㙧l���p�"�x���tV�Y6u3Z3�mb���J��X[�Dg��&���!�$�YϓR���J�7�Q�� �TOPt\�s�J����G�G�OM�E�6�v����M|�}ͷ�D�d>�Sw���tB%OIߢeQ
�[f�l�w�>��@|�/�p�|̶{��#p��1_T7��f�rzVPp�Y&���0e�9�q[�}���X#p뉺b+��!Q������Y�¢�c*1+g&3�~zj"R���HR}�ƺq*ok�NW=Y��`r��:M�l�V9ҏ��U��zo8O��r��#��5����qأ�J�)%�:��j�^D��{���
Ⲟ��u���B L���m����bmQ�P�%l�P#��1 �kE}Q�N�>K�䥎���W�-X	v�]�Dŗ3����js
�Ԁ%�Nr�c�U�P}�b6i��x�k��g�q�R|�nsF�F��vn'f#��:oS�M���}��*W�o*4Tu����ȧP�ԅ��y�e962�j ��d��'��>���K'��Vmi�o��^�P�j�g;|-@�<\�]��P�7�(�Ã��_y]<�GZڊ
�KG��4uG�e���;�P(d�p.:�1˺��8ɫm���u�����P+�$6��o���"�*�%r\�J�F�@��$:�s5�֯����c��}|�\"��fV�c��v&�Xf>�C"tOU3��U᧷ݛ1� Ae��o�|n\ ar4,���c�t�Λ��ˁ<E��q�wب�q�˼�G+evS+ދ4ޖ�s�W�딸�=�v��	*��(h��u»CFI�Xa��:�3*P��X�k���a #�7%��y���rM��b�땮#+����AͷĊW�1ӎᓸe ��q�jZ	��k�dx�&��ܹ�\��.�w�kA���t �f�-}'t���W��e�q$y�x�+���*�d�u�73���1�δԼ��?:�(V�mt�G9����hw� &��kV��P��7ҏYo��rv��z��+*�g_ȧ1��ِ�w6���J�bG��F�Cۜ	?;�ޫe�x":�_r;�F��=��P[q�c��kcN=�Z($�k�t��:k�-�뀽���u;z�2;��u��P`F2��}�/����¥i����Y��dt.��oo"�g�jm�]���n<��s~���̢�mǧ�~>/��.��Y�fJD��˗Yy5��;B��2���fH�3���q�b�VQ���wP����Ȃ�ʜ�Z1E���,r�F�>ZWEcf��Vw+QC���(�,�T�6�&��cmLw�a�3���G��g��� M��%�z9���Κ���`����5^���i!�P��V����Q\ ��0KxG\����\_d��lEs`B�����i<���-���9����m>DЕ�V���Rw���7���29PpU���覠�lN�l�[u�,�kF�V��R���ַht���*A����vX}#z����u5\D|���C6�����"ޕW�sc���/�֟[�>�[lc�S��'lsʇV���8.���%��s
U���]���hQ��5gEY��.��b��WsH
]9��jn�|w*s��@QtjY+��l�c�zB���x}9iГ���-@]X�P�k�E]w�o��c]���΅;`Hu�fX��Z�u�	�II���ꠟ���L�����YiA�K���6�]c�[�s[�u�,�;�A�UF��5�(*�) �06]"h��>{Y�pjT��-��+bT��F�:(��u͕���n'Y������c���vk�e�;Ε>W��]��5�5�z���
��Hw�b��Ȍ�N���<��Lاs)�멊�����S��T��eӣ�|���VT�u�@K�[�B��ձ��_3��d���&�/�.�#˖�Us��Jo|�7��θ�~v���!}�e��Q�u�mމ���C��P�Ր��d���yk�4M���ܨitU�ق�Y-��Q͐�  �Ѥ����mV#l�#�Vad'��b�
]�W�ET��K�+ʳ"#��T��}=rr�Y��T���J)(���t*<��"��sS"���{�Ҩ��y�I�+ܢ#R���̀����(��_D<�f�*��Z��A���f�Q	!9I�R���Uk�.��W���r"��P�y¼� �s�UG��30<�t��\W7<�
������)$�
)Q3<Ш�r�E\�7(�(����Oz�TG<�>I�9�UC4���B�
"�2�/*�*T�����%'�zL��U"��6����gc`�Ha.I*�QQfW��Uyu(��(#���^�}u�J�fF��S
�����Ut�#�)��\��2���hɑPyZ��tܢ"�^D�r�?Z�>曖��y1Ă0]u[�Շ9e�ެQ=��Mn�m�7��b��}`rS���j�}�+8I�P�r�P�?��꯫�	�d�zؼ�(b�?�<���F�!^ө��*��O��f���뎻�ESE�Y}�/���Or���������e>1��J��!����RH�k��Vwl\���$�<��s���Ӗ��]X>���:��"��q,n�0tCqׂ�:������N�����}�w��n�\��.Re��G#B����N�;�rDs72�)鑱f� o9�7�<T���K�E:�o�+/(v>~���.�i3C��*��L�cDp�nFx���<�Ǯ!��Ԯ�˹1�d����R��6������k�����=Nbʜfj%gP����y������=��r�>%�>�ů��/I���]���FXۂ���K�,��r�bea���]�db��\������T�a��v�y����K\+�b)ʓ��mbt���k�ld3"�j@n�{�(d�nO�Pܸ3c�?&��vپ�O\�ױ�*o������A�ڄͷ�lbuE�s��[wp�\�?�c���Y,DL"���C�}������ȅgn��#K:��Su���I|֎�{�S��n��w泱x�f;�o�$��˷���"�Q�k�Q�N�ܴ ������n_TĪ����'�(�WW����i��ǜ��#LT.��3(������Q��S��6䂅��j�~[��T���
�7��-�#Ġ��9�_SYG
qTci������vI1!�у*r�fL���6w�r��,u����xiS��)�;��ș݊�X�F��(e��2�t�
��U�*���-*��@go��b� b� �*�T�nL�C�= �0��p���Y����nLX����]g�������>��#�����S���X����	�w[���p��cg���Ī��=bS�xw)I�K<�+�̌��Q�
Q��$�q�p��)�����c�F;>wLh���YC"Mۅ OTA�\�K/{.�L����;���#�c����#�1@�}p��]6s�?1�o�i�nJ<�nS�8̎�OQ��s�F��[t(�b\�ы�l���&����-S����5�^[;ܳ��}¹@�r̲P�D���������1\��WU�4�5�f�{�;��T{��|,����=��uR�'���Zz�bc�]"b~����R1���s@�����}L@�Ҋ�݇;���9� ���F&4ʑm��^�'ŋ��O9a<�9�2�ʾ�����}�:��b��t��W�5��*}(�S�ܠ�����RF�.$0��wyz�fp]qMVs�1ܑ1��L��q��/��Z;�磌��;о�}=-�l���4�~y�;`
�-��*�$���i�Jّxy�"u��U�fͫ�gx����"a�)��o����e u|�"�� I�7����}]e@���9�ob��l��1Z.�q=;�0�W��ĺ�\rV]�p( b4�;#6���<j˝����/�Ы�	�o�u��l!�f�:�9���_��1h�p��t�{w���e�@`�{��Ӂtl�0�H�|=��<�+S����T�p�ƽn�y�K�7���#F#��S����:ٳ^�|���[�[�a�p0N� C��`E>΂�C�e�����wb#ݸ�(MPs�eϐvXv%u��e#�}�M���s���ߎW����G���gE�m�]�؝2o�b�n{]����z;߶��5�փ�Z%�0�C�tk�QZz�/[[�?8Y0YXH�z�X��F8Ck���(h�{�t��a7C��UY����u�ݹn����V�1o�!���	���}���r��C��'L_�gFȓM[E_�����`լӎƚ�7g8޴����Θ����(��X����'i]�񼌵!�j�(:͸2���/w�P�����R�w�V=�nwj����1��V]�p9:P�GV���.�}~ �{=�}��d\��T;Թ�;��&���}��}Z����|��]3�V�^-b��� ���6tp���[�O���+z����V�]�SW��*�)�  ���q!���D�4T��uN�A0�c����DL|�֊ITE�ڙ�{��k��z�K�>{�+N�%�ya�k�wQ3!)���,9�ci�8
�U����m�]�`嬸�A�t��nP"��
�WT�M
��b�����F�+p��β�z���wI�5\���d�����m+��uP������ )�FC��j1.(�n�[;��H`�<u:ר;�Q٭����ld����5�p�|�q��p����x�g�n��Cꛘ�w���M����G�р_1Q���_�|3��{4�J�������f��!Nw<�B�w@�������)��I����:����C��>N�����E��3��6в���y�܈�ok�_.��Yȉ=>�8��++�'�3��֫z\��:�Vr4 ��p!mU�r�0�S:�u���#�D�NE��̫����ە8%��Or'\V��&�km���x�?X��j-��C�ӊ[kŷ�n]�u_�=����1�O���WPt��c��+R�do]v4��i�����gl��y��()e�[u*[�$�i*�Wa�*To���ԫ��a�e�;�w�ҙ1i�l�<_�_W��W>��QP}�n������[ \	e�I� �U��zh!b���N�%e�8@���/�F�S�����qm����^�k�+���f�:o�N�60Z;��������];�^w<���ak�4�6HyZ�C�tk�����ʢ�|*Q�?�}ܝ�r�V�3�d�^�nj�o��݁g}��gL�n��@q.���-y�����-{�׀��Fe��� �|�ǩi��;xy�S�bk�2��,�dШW��7�3�|NY�����& F��I�8��{��Á��.3\R��§��()�JB�����a ."R��F�S��|�^��^�^�~�l�eg����4�K���E7u	%�wM�4ka���������m"���޾�X!��t48m�3����W����/��Pg%Dl�*zI��ʁCۙ��'w�@���Ttc��GWi���k{z�8������3E�`��r0�����PS���!s��\�ps�< {�L�MI�`�,�뉟�L1��]-1�Ƌwzp�%�ʤ���b���n���¡CZ�X�LPM3�y#���0���tr4C>�w�P����<v߳��3I�\i?3�)��|^��7��@�]�
��ǵ���ߋ��q��1|��r�N�`�Rb3Z�v��kS�!]�BVx+��K������UW�}��_����s>�ɈڎwdY<NR=��(��Qx�T�] �s���q~4 ^��RyK�y�w^��Z=ٮ3+ڇ��5�ƀ�o�����:�o0��yb?p�|��W�x1�_����w�2o+�ئ!7��V]�0���O�hs4:��1f�����=(����%Ժ�[]�k��^�Ng��F�a�\�.?zaؒs�MZ���~-M����WY3���y���j���N��#ĨnO�وs3Y�r�K���X��*Fˌ:L`�ÆTNRq�B:��+�t��Pcc�b9l�:��Zx�g<�V�iNbKD||)���:b�0��>0�Q�(Y0��b b�\��q����؜�)�K�i�� ]��0����������F/0JD�b��*��g�������>{2+��tl�Z�Z�]O�����=/T��>��֏z���-N��|���k8��dp��M�����wn�B�|��d���+/�1���j��nH��.�N�"���;��ts�=.���j]��k�۰z��ь�
ќ���h�w
�ۗ��
}�s9`I���Y9MM��ۘ�m*#��Q9�����%��dT<{;���fuЈŕt�纠��S_>�RνT�|B*7�6��u&\���}U�}M�JI��^)1�y���َ_Y�U��(5�O�E�e��1�q�!�t��[SR622���2�6�4I�UҺ g�(4b��Q
xh���#�N��f�jq%���N�x��z�.��:!��}>T��ֲ�g��ʨc2#e�O:����\�<�n�su��W+6�����s��F�����?��;)R����_3��ej]Ƙ7�E��>��8�7�
M�!��oe�p�U���w�ހ�dP�0J����M}lL<�΢�Xة.j�gbIuYŴwp�3�!0pl7�l�����tC��)9"��7����Q7:�,o:*���y�C����Q�+���71���#+S�f�@4r%��B�IʏX�ott^,M��}�s�d��X+��_^Wʮq��8�3]҃��w~�`#���mq�f0�4�9����S�ue_�l��@k9H��tmp��Wg�Ea�ux��7� �;�:�-��CT�˯:��ҔP�<�:i�U���Θ�a�1�L!�e�B�`�5ڨ`��"��6*l��~"�҈wS{+p)��_l��U��c��q,2ӯ\Kب���NV��=ˊ�u$��y~T����ze���	5��ʵ{�j6w.�U�@*]�5����k����X4��Ѡ���x����8Zn��aw�=������wm�.�d`��G�ꯪ��G����A{�=���p�u�b߳g�?�,;�9H�-dU}bb�W���|�W=�;�૚/����u�?\g:d�1l��;�5��{p?����%��#�ެ�4�|����Uܟ?���ҩ�cx���I�����r1��CE=�<y����1ͽ]����6�44qU�M�w�J�]0Y�惲YXm�L�|E+xs+�uI���Y&�1]i��� O�y����g��YU!�4��q�Z8,l�UZ��L��jS
���xn���x����b��G�È�ߙd�\~"xs]���]��ZWc{���[�mT���{���k7�C�f�p����O4���4����������R���Puvb��dJ���ɚ�F���]�!���r
�:S"�R�G_�
������	
�.�k��Hp{���y�F�b��7q��3e�h)� GE;d:�r0�
2�g��L�/�3��ך4C0Xʃ��Ӹs4�g�����P��7�\As��9+(�#&�fd���ӳrn_=uo��f6�h;��{�:^��6�I�뢇2���8>�XO!}�=8\��'� ��X�V�n}*��w���鏹خ�3nc�Zwp��^a%!N���:�s#m�iAz����G���G�U����p,Y� q�5(FŹ!W�;����\̓>}��e)'�������}�ە��g��� ��c$���혍`�M�l�t������v/dοb�Usѵ�\���<��b,��m�")�����To�"�t<���B�������՝ٱ�Z����+o��� +���
f�I�*6�<�q}u�G�v����Y��ťRA���˽��7)��b�������S ,4�%3I�j��oL��)��b6i{�A�^Z��bc��Zb���r�r�J��׺)��U~2�|�ɥ;d���C���MgdV��a����Z�|��˒�S��y��aW�:�.'U!�u�ZN�6��+�m����RKwehm�@X\fg_�����E��-y@r7�(�Ã��mw��5���C��c�6���MO�u�+�^����Mf��1i���אc���Ǧ��;œ�E�J,����e�z��/F�pA��/J��p��a�RM��Uy���E��AmX�ff=�i��G~�b�P�ϡ��;V_�%˗L.o|Gnv=.�g�'�'b���.�Q�rwnnf��M�kj�-�t�g���7��^��y��Kۣ|'m�:VRm�+9
8.�"�e��(�]��vq��%>��=�>f�'�"��꯫��W/{I�"> R��D�?!V���.���zw5�#���b�IG��Gt��S��
��)t<W{�Ɗ���f�^�쿻e/�7Wϗ���7 G#c��n�H��q{%���8��BW{�`�� 3-{�G�:�����a������U��f˘�4��l{״�˝�,��$���LK�1���]q3Ja���i��cFRN��C�ȳV�1�՚QG����R��V��� ?�x�%��i�J?�����]Q"��S΍5��������b��.O�-j�E�!��=�`�9����(�}V�ï��_f���
�{��Z�7{�^�!K�c�+���A� =
��l@��J�T�Y����P�gwj��-�w�m>;�8A轨L�y��s%�+�C��uP�ඎ])��efջ��%^�=�;�1��+fR5�GS���8�Ck��R��J���g�Pܞ(e����vV���ٗ&�E�(1�*r��2#���qڨs�E�Q�����B�.an�5���R8���]ŗ���[/�+�/H�|`�T-vv]�����v���e��80)[; �(*ti�{vy��Y#H�"v��^U�r�[�N��캎�+/8ŎްA����fdv��<�p!�z@k��u�����qnmg>g��+-f�L�}wv�bfӔ��bٺ�a%�hP�)���l�W�Ի��l�?���<��	.�u�2�R�փǢb޺���+7�=S��$��(nn��b5j�H.�q2��H݇	u�KV>��õ�j�#��k���*넆�oTk|2۱N����h�C"�6�B	��f�m�3����α1���.�H ��e�cZ�Y��k[������!6�}%�̭����1��2'r��P��F��X��׭�xP��2��6����T�|�����A��t�]�s��hP�qj�x�U���fo#���<G:�n\.�¦b�� )
ŭ������)�.B��-v��c�/Up�o@J#�f���x_p��>՚�a�`�mӉ
X��oǰLu�I�
�%���~�it���%=��r҂�+nLkf���xݰ\�{ne�-^��ۣ������� �]��m�稄0�P��aA���K$�k�R��p�Ǩ�ӗm$�ժ�.��j���t�_wTz����D���]�zkrjpmNX p��ôN9�t��1���4���$O��5!��p�N���!�1��E�sҟ�mo%��܊q�:�ӖC�ingV=�H�����k�c��gO\�H:;���kYj���T����(�4�:��m��]-3��mA�޳����)e��B*��_����/ϳ���#qx�\ծހ]v7�{��V:*ع�Ը!�3k�˹�˭�c��:rdWO2�Ao���xk�nu�}��]0���c�h�0�+�V��~�pCz��gg���X�r�a�p'��_�Xۨñ(t|:�g_^t)BF�μn� �+�EM̀��n���7u6r�nb���ox:�S2�#��dT� �	W�n����ɡ5�����W�g����z�$ZU�����i�]Y�Ҳ(ѧ�B�����ŗ�#�]t�kf��PR�r�Z�@��]u�I�f�^�Z۶o��Rɏz�
Ìn&~�H�p�ix^�\n���~y.,�ov������=�+У�mh׺��Ńv|�a0�J|@�`�ޑ3{8%����՝��x�`��]��w��n�"�SJ�O�a���k�@��4o9̷�Q�oi��A�m��k*@��oPŔ^�#�[��qK�^i�7�'d�V�XګC���(334��g�.V�
�yOvt8�*��a�DN�]r��b䰎�����D_�o�����9%@�Co��ϛ��C~E��k�Pj蠍�Q�n��RUEDG�y�Pt\�^egca�A=�EPDQD������G�P^_W.B^M��y�E�Ejꦛ](��T���D�*��B��,-˫R"I(fTS2+��J*�'(��=�Z�m\��Ԑ̽��Q��A��"��Q��
���W����R���G���g�Р䙞�K�2��	��yAU�yrg	]2�/H��%��OO��(��xWD�y%^s.���{Q
+�T��B�**��*�r����M�5���**;ȉ�(32��$�����9
�x^�E^��q��J'����^W�v�	WI/s�L���<��jQj���B�%PU��29�F�EUy��Ԩ/<�	UJ{YU�"#¨�Q�TV
��,b"+��^��G���&*-tjeu.X��.V�I�+�-�
R�y忰����޾9�]�,[au+Y�i�� sO_��>��ʗ�)7���(���o�}}u/�� \7�<+�>U�(���a������S�I��hGRʵ��!.�;���b �)��W(kw\7�kl�`�{�#j&a3C��ܾ�Ҩ�Q��rn���}M.����O�C�h����\s�Ρ�wLm�����
�ٱ3Ƥ���*͔��%�7�nki��� �>*���g>���zy��Jf;+=~��,�S�����9����c�x�3�n̎Ja����*��ƒ}p�t��������ۮ�t�ʩG�[���,��C. �"�E;�EJ*�޿p�ù�����d�.�B�E��!�OdSV��E!���fc2�**O�0w��������y�ÐT��XG��B���Ç[�5E>[_KɌEOk��dak��'��V�����r��������&�dF9�ʣ1��F��z]py����9�V'z����b Z{&@Ze(پ�O�J:�\���VC�Vѿ�L1܄����h����-���B�P�!2D�njf!ҧ�WyZ�>�J�[�����p�5�ϱ51��r����3�sT�/�TcJ���qUw�s`�{�8l�-s��K=v�a��v	;$����w}٤˳�:����,Ƈn�BA��tݜ�0q��{]�%F�=d���W��Zv5�-�* �e̦�ξ�²�n�n��7�~�����R>�:���y^x��eD^Q_Z��Q�/��ٌ��DF�G'f;�7^\��N�oN��P���C��	Β���(G��U��b���3;�t��<��㽕|%��&b�SD���Y�%�O��͙��ah��\=]�1Xb���@^��u�C��O�l&�
�P�W�q��]�hE3ms!�5=y5Xc�TNT!a�C�	À7���\��fwT=�@F�Τ)�"�����o��>����\���W���Cܫw�o��{�L�O5��}"5�nS�q�< ב���V�"n�{;�+D's�C���t�9Qdt8R3e�6�e喳s ��_��O�CW���n��j����}0��?f����I��F��eH�/]>���@!�Áۊ���XP�;�	���Ņ���L�e6z�ǹ6]v�����,S�a�MvR���K�Ip
���2�h�]i!증��TK�O��1�eVoa}�	��Έ�G0���[���6!ۅ���7��Ѣa&��+B����+�f;h1��ZW��4|̠U*��Kt�8wJv�,�k.�dv�J�Y|�KT��$�mf>������'nV7>��3;L9�h5r�(�&����G:R=t���u����v�֍�o�I7|�^N��¬r���U}_Var8��w�0����C�ͼ���f ���l���|��ۧ�HwJoY����>���o8ܥ��U��pL ��{pz�e�	
�w�Q1l�a�)�JQ��P�s�"����Hm��+�jN�1��ohs�G>%���#_0�U�:�L����h���+��=���jW�s�`��E�2���_�N��;%3�v	�4��7�_��"��lnE"�ĳ��w���o��ۄ�
M�]�g�>�ܐ���鏻Uk=��nh�ͧ*���`��MI�ᒳ�Y^�O>�c�7~�Y:8��Q�i��PvT^����Ά�S�y9.gpw�H�x�<<���舨k+�tA���J�g�:8�����7���o>�H����4ZΤ�T0�%,1s�+��g��(H��W���[+���t��G=��X�.e����cv�g�z�a�r��Na�n:��f��H�br�������Ϣ�}gA��ر�5��k�j��vb1��΀ۈ��p0Z;���+��r�Ξwb�h�+ �7�>���.�AQ�
�Rю�5�����h4�.HZ�Mn�s.Fٔ^)�bC��2�{&O�6��Sw[Rs�L3V�wBx�ks'oKo!|���7�sk��p���>	�e^l�o.sb���Nh���@��
�]d~������Y�;��7�����V��"���`���8���H�V�.5�ט���g1��-�=��N�딈gN����������+t���pQW���y�ޫ��=����юΣ������]1��~��>|zr�?T�H��ǭ켩��n˓2��8M~��\�ۥ3���fƁc^m$U}Y*״j�Ch����ٖ� �v����3��
�T'�"�����F�E7u	%�t���W1�umկ06׉�b�,_ ��j.W���Q�U�e"�"�M�u�����Zqܷ3�t�
 ���AW�1"J��.!�n������*��L�.�F�� e�~��~�x����f!ge_�:�r"#X5��V���婆0U�H��z+�-Ɠ�ԻM^*	��=n`;�3=�1-ݐd��p�8����)oM��[92��o��w#�׃��Cn#BN�����Ѩ<ꇕ��8��a�Q�h��hf���Ӱ�^���J�F�:�Y�I��)Xpm�W)"6Ȧ��k�]��}l�i��3�w��P^;�<C�[t0��eL6q���f=vf�(kn�Rd=�eթR���Y:����W#�|g2ӎ��e�(�� �8'vk������� �]o��fZ�I;��?������E���8������d���*ct%�&�oU��yT$p� 	�W��}��vU��9_j\�-/P�q��ڇ���2��ו�^�G�T���9���D�wp���*�ΊץE��5r���\a��c�	aYؓQ~����ٿ�e)���Q�`ku�Q,fވV��C��e5<�/�"(�����[ٕZ|MXc�E�o�ʴ�k�����P�9���(�ւN�eN�[�\�lP��l�9�wk�Y�'LTq�xW�R�}��U�^b*�:��X���]�Y�V@]{�C^�� j_�W89���m�c,�I��3	�ʯ	�tkQ�u��+�fZ�<.��-��1�I��Z�q�|��R�r�?+>��/&u�d��8p#Ʋ��1��ٱ{.&��/� #�]��9����,<7�k��vC�4R��ABٌW�^k3o�\���H�΁�7E	�0�fE(1#8�O�"鳑��7M8G��v�gU��S+_|b<vhG���0�.!��5�v"5�с<u�N��	�K�$/�SV�����d�N{�6h��ȃ�.�f��\��wg%K/���C��Y�;J�&�-&fs�yꝽ�cTݚ�U���R�H������H�s�[�����G{v13���uj^�]����'��3�������]�R�Y�_PM�Ź{3��]���ﾈ��e��.n'�A�zc�����`��r*O0{�����MOQ���{0����e��M�Öޥ��z�k��~ڇ:�ok���r�ʃ��@�{ϕ*�:����[��W׊x�x��77�ғ�����5�\gC�����V"�<(���^<�"�1"IZ{�����՛���S�Y�V�m��c�!�_o&/�&���R:��`���dU �η%F�l+���:$H��V.��\�F��{Ҹ�8�Ɗ���\�l�Cj�h�ᣊ�m�^�C*vo�,�eOe�^��p�-�Ό����Ru��zU$�w혱EClƹ�:�7�Rvl�J$*P��kg���z����@t/�{M3k��\=�Xb���*�R��ʈ�Tq���'�h��B��p�jN���V*}��p���e#Z-ҷ\>������R{*�J�_�:�\XP�y���(jPN�vO�ux�,��-,V��pS�h#AU.��C���*�����%�1�.�g����S9��T>�F�ہ��a�J�qs�1��*.9T�D��ͮ��Gp�+7�'�ԐlŤV�|�4M��mdX��VJ���3�)�&�~�����~]ZY��&=Y�u����z��Oh������9�m�S�.��ur�z�p�g_ŕe������}U�}J%&L�]h��;���̆���"�c.�*�#�Ҭ��o�i�[��񜒰��(\����w�ь�����敟l�"IC�ٔk�J#%b��&JsA�,�9{���X����T�SF��ɍ��J�ڴ��X��4�Mf�kG
�S!��p4�G;�#�#��z]s:6�=�>e鯭^<�>#�e8�D"��;��ᤡ�'N�	)��y�|�#�2���Z(\sj��q=�r�-��`S3��>�(����Κ�U�Fn,�ה4W�5���T�I�9��K�����y�l(X�J�R�j:��ŝko^j�皗�wO�*��Y�G���pJ}¾b�J��&x�����N#7q�f�e�p5oxU�$
(�$��,:������9�i��q�Q�)�����1�/Ҹ�罾�S�ή ��8wXM3���Zz�n��d�#�����֌�����K����&�mR����&����}�_{L�с��7��'l�k�n�e���/D����1*ۙR��N���n��Vk�1!�J�=.]N���g�	��0�ݲ͛\1N&�v@��˪�}�������x�u��\N%���)'m���5b���,�}\8�R�WW5����d��f�]����dI��}_}USs\�=���nz�PV�%�rEBj��k+�
�X��y5��f���W�'않�LS���od��j1of��u��L0E�G:��N9�6~n���k}Q�N���9~�z2�d�~W��]�/g����]7�Ɍ�3������d�'P��P,�C=�C�7Ժ�)܆�3���s��. ǤGƀ��ڵ�引��ɭ�U~-s�7y�%��Ԭ ;���ْ��w�=�2S�Z�V�6'�������aW�:��B8믳mA�إ����С�U�l%��c�xH<{>Ͻ�Θ*
�.�(%�]E^!7�]xjUs˃HV���2�H,��(_{�-�R��yO�����n�?td�?@��So�jw������FѾl��*�_�c�W�.�<����t�.1ĭ1pܱ��W��*cmHU<�X�v�;Ϻz
�����N�Վ�����"�u(pX쿱�)��c2:�{Pp��c&Ӧ�!tQ�Jh�ED��bG�����\h_t�J]w���+x�4ۀ�Ә��J���!:�[��<�^�.gn���֘�F�W[[�O����֟� �]HQ�������D$�٢$>�r?i��d:��n��8���A݃���d�N5����;�˗q�n�w/��.Һ9}L@�-h�V�y���M޿�_}�W�QV�w��b��ǭ�y*#X n�JUܪD�{e��}��z�_M���.�eG<i�J� e[�'	tE;qC ���s��ek����	e_57��u��:�7_��;�;L�AwP݈��&
ި4��]3�hhnZY9�t~���t���認I�_�T5np�= �&
����v��ӌ��g���T����i��������*�P�ʺv�P*�	���im�PXk��i�YPi���u�k5p5�ru������&�ZݱZ'\��ʮ/:�!Ji�*��5}�����/���r��{��(�T�m��N5#��YӚ���*C0c�����`�����#���l[����V+����7|��v3����������eOE0�6��Z[C���$.�o������O$}�uI�X�ˢ�]=���z�˽�-�c>��ۑ��m�Zgcm��O1oiNwe�L�{�
ܨVU<��Y��&�<�yOx�ɫ��"w��')�ff�s%��^4[�o-�W@�@⤨w��V[�5�̚��sb��\����W�e�o=ఞO��T��yN�D���=�;L�3�����|�'��I���着��)>���Hs��j�K���GUb��C\��Q��o�ģBu��$}�y줽CZ��9��;��t����io/.�v�G��&�2Q'�rJ'��ܗ0���9ʹI��-�<��1�,H��lOڍN���E�8�Q����~�0oW�.f\*�YkG����R���v�us�S�9��7R��}�2i�W�ﻞ�J~�����%�e�yf�y��CWK~�c~�'ms��j�֎x�[�(��Ao�Ki��������խB�x�m߾��#�9�H�m-�=N��9����&8J1ۢ�;s�H�f����¼����#Y���*�Ɍ��ոP�
Q�r�^͚2�0,崅�`?��p{-��m�5�\���%G+SpCʚDv��I�G8���<��@o��{<��r�K�Š�w'?|Z��g+d�
.G�j��Swg��5����6�:�4΍����cY=k,��Ɍ�fv�̮�*�V*QD��y����;��	"1!����\�b�@��,q��˵*�۩�'��[8���G+����>=����y���ݙk,}]��]q�s��#�4����CO˺�b70���c7�A���X�� �U������X�3,���Ugj<�D�m��en�u����,��Ot������Fe$�&���	ۙ��L�r��V�{�KX��i*Lދ�pھ�*���Q�{��!<���DP�2�۔0����4!O��\��]AB�W�ń���r�2t�>��f���%3A�N�[�ӫ6��{�ٌ��U����K�7:1{���~���I]ש�;��B�㙚��+=1Tu.r|������Y���v�T�n�F�o�����|6��4�M������lh�&𩗇o+��oE���ݺz�	����|7����v����-7�3.�
]|�<9�!eu��)���ʂ��e�3��.�cdd�ː��nhX��;#̱۷�!�Gs�'r)ˢ���7ad�l�t�Uj�gv(�CɷΓ�̶0�E�H[tu��,+��{�]�:�����8���j5&ϟ�ĺ^�=e��I�xՌ�4�̳w[=��fD������{0��[t�N�z��y���@F��ݷ�K��e��hu���dΣ}h�ik�k���jt&2n�)�&����Kv�Z���9e+v�8zWNu�1���kY=�9DJ��k��:F��ً�s����4u-��;{�7�uv�\Z�&�ݮE�;a�@_����^ {�����l�"8[�:�*dJ�攥�e�Y������쫨�2�V�FR�»^�y��^o`��h�2��>��Zo��D��V�tK������P[b���l/�Bd�&����#�g.Gs��F��fY���)��S0f�W�!�zf�� ����3�47N�c�i̕!Pr�9*`�<fN���I��ZG��y�Y��!����⨾U5.�����%�;���N�+;3s7+�J��>�\Np�3�-��o���i�-���]��l{o6�qr[��Yu2�@ݍ� �,#}�����MҢb�n�1:�n���L�0v���oT1�]v>�Xɇk�[j���{��P��z�m�/V���.��ԡ8�t���/,n�KA�H���F�7��-�|,�`��L��|X �P�}�'Yv	�M=!�����]|������a.L�z�`[��3Д��n���^ր:���K��6"X���q|�#ל�P�/ �>�|`�dɩ۳%�g�F��%��[����ک6�}8a1�k/�Q$�51��j�۳vyj�7�i�	�$4����K���>Y\v����B�>�@�k�H�$5�<�Ӻ�mh��xXh$P{�!��QCģ�"޸�+��*�r�1"�/%�PE&M\��b��S<�d�6��S9Qst���B �®HUJ�2\�bɅ�jQ�b2���H���]]��Y�x��;*Ҽ�2)! �D/��"fOz������i�:ؽ]ryɘ�EEy�X_Ȫ����jP�*`��e$�k����{�Ш�r��$���sȼ��lZ`��$�E�<�.�P�'�����h�2����#�=��L�*
[a\���C�Xا`fFD��!u%�k�m���$�ȍm�"�B��$mO�+ᒦDz=�׈��(�y�,*�+��vdD���Eznk2�"(���t�ƹ�+����	��T��mB����E�H���70�+$&L�Q��č�aW�څq�U5�15w�0,�6
WfV��-���]��]�" �'NJ�5A�wɱ���'3���Ӎ3u��ޒ�ʓ��"#ﾛYh$ݚ�v^����Y��z���l��K�)}qJ�S/�=��ކ��V�(���=����ek�vU��R��%=�/s�l�a�z5�g8�Tش�p��ݯ������ioz��i^�r��v Wy?z�N\��:�[U���O;��ب�o/��j�v�2E|�r�u��p��WǬmKs}J��w9<����&���k{�� -���Lif_m�.��y��R�ֵWɭ���OS�ǪU<���Jx�ʰ�U��5��3��c��j��:��Z�;�Ű�h�w��#�9��q���Yq������M77�L-�P�FF�D��I��ڙ��*o�mx�=ޘV�h�ig��ݼ{��:�L�@��}��5���bN�S���?d��ۆ��v�t���k�R���
�[�)�#������j�g���@�\����3� ��ӹ��)���E>�&r��9o[NoM�@P�K�8+t@�o+f�x�-����X�m��h��iw��l*|J�l��n��T��+F�����5Si�T��u�*S2p��6����3Z-�.Ń�!��UU�۫��>��=�Ӟ��Q��d-wave����}S��h\#�m�NP�����e\������bV�\iOw>Gr�I���6��+ Yy�{�Ҋ�1�e�stBc�[�Vo���ڵ�U�a'Im<Y���8�(�r��6�9@46���iuE�,����T��z�u����4�:��:�!RhmD5��W�����4Z��t�Ʀ�ڝw��o�{��7�������wW��:�q�M�5�[�ï��Fi4�.�u��ʃ��ֺ��ʎ���g8�Tش�p��g4���_m2�Wj.;�-���*�ʈ*��To�-�Tl�|���Bv����Y���r�N$��V����^<%'o$��q����._�k�,����74�d�V�wS��)�}�
�i��>��ۑ�6�:��q؍R��/`~
*�]�Ӊk����>
����Tޥ����sU����Z�g+�x҅��W��~�X/a�;��/��R��3GG
��5^��X�jn�>c���Ot�����RA���|�:��ۤ���I����r�̣.�q�J�r�x����ii�z��]����+P��n�N�'i+=���Ʋ�Mn;z�����>������WLX�$h�������Yažt����|�Kyq��o9Mr�6�л�Q�������)��tf��o�_4���eq�����ߛ^��k��0���b�t>|��2\A��Gt�U.f\*-s�Z:~W�4S����ɧ��c�aI8��ɧL��}��J~����\.����<���=���k1��iɬ�q������;�Q�Oȣ ���+����U����<��3�b{�;�;���ۘi�/��v������D�������~�X�F�w=K��F6C�!�ܚ���d"�9I:p�=���&o� pzz�!s�v���w�\���+Zw�Ǯo��4+��8}e];S�X��s��¸V����@8������(�uy���f���:n��9�)ؼ�y�%=d�+{��/}�L>�R��L��jLR��xh���5i&4���Uk�2���:��xZ�p��v&vu��i>�{&�B�q�P��2���nŷ{�34���Q�ħ���Ob���k��Ǎ�̑��Њ\�E9�ނ-ۅw������otv��{컭���]G�+ӎ�����r���g(���M���S&w�y��B����W��8����s�es�_eDWg;m�-�1J&�#��wm-W	<嵉�O-ho3a���B��h�������P��!k�L�,�yIY�oas���y�p�=ˆ�S]��՛�]�kN�{���X��rkM���j�Y��r�_�Ue�-kn����S]��nJ]jK�\ժ��aP\	́� �q�P~�j+��.��>u[��i��m9ې��u�2v�]��]�o1���j������Z3��껽<��tH�'>ĵ�R���v��[Ni�P��Q��.f\-5vH_VG{U�;�܎���x�PM'���S�j
0#yф��N�����ޗn����U*���֩�Rή��
��*�baz(-돪��o�zo�<�\9.��y��̼�VuL���Kv�Te�9k�up0%g��qV�Ȩ�6*�mͳ@S���k4������l������
�}V�] ~;��v�qY��1j��혖pƆۍq�Դ��	9�גfS�u���W�����4Ru��$�?�z�Yٗ�:m.���[��&��S�f�_f�\ε��ؠC+v�-��b^��n�݈�Trc[�p���֤�j�f�'�%����m_�̀*��/zV�`�xz�k��KtP�s2eom#�Kkqž�Jg�t[�N���2#��+X��y��Š�}��E�=|�=���}�͡i��چv/��J��GY�f��.�&	��_���5z�#Ҍs|WD�v����T)n������˫��-��kj�E��g��8�e��z��oi4�Wד��5�8�Sb������fmW5h�ݷ�OLɍ��a��'��qv����.��=�!���o�?O>�O�:+��c��u܆�w�W7�G`t7>�sԬc}���:�.Y��<��"n{���o�������t�a�댃�W�Pb���N�m'�A��MG��x��B������i#H*��o�P32ph�5�r��*]OG2����Z-�Yث �{�q�;1���z��a�<���:�8)E��K;��(�&��A>��.{����.�!��ev�E�-&�����Ü� gLؕ�����ꯎ�Ι;�������zz�"��vH�>W���L����A��c\�'���JOYw;����>w���1�ݸ�ޣ-�mGf[��k�ul�Cܱ�c��^�E��h�O%�ͥz�n��[��i��I�;o�r�����n	�S0밹�\R��㴟sw�v8�Rn��F�9h�TѼZ����0�!��Et��Xf_�J{�:�v��7X�NǒV9B"�o�w#��bQG�[�Q\�̽)��;�]7ݖ�{�K��;����G?��MCI���:��S$��+i����w���e�s������v'&�b�P�ેAP����.��lv�9CG5�x����L��Q�A��뒲�5N+�M����QX�+��o#���Շ���bu�c�!ņ��Ko-U���|Eꄥ��!p|3~n�N�NE~�:�f�� �E��<�z�٢\���wDn�Ch�����$h���J*k���4�4���#��B˷�S��:�v�MB�]]��[���7Ֆ$��� ��e�cT��&f��gS|�u˥#�Օ��8��G���"���Yyn���UUWӳ�Υ��W�P[~8��ޫ�yu>9�*l\o-hC�\E�2�6jd�K����&�t�_Gih����qM�鶺�����-��1�+1;��m�e�܄����{�j:�eck��78�cnٯ��Ol�O��yJ+�����zg�'ox�[p�6��u}X��TK="D�h�ܷ&��X˗ZW9\��p1�m>���)�ˆ�>��=8�;�+��<�Ź�in�^�;_!Q�W�);)�4��������ʭ�/�l���:ó��,XWq�23\J��J\*�������[�p�J��tL.��Y],WV�y�l����;�AugB\*#1O4��2`��evj��udΠ�{�o���(�ȣ�7�|a)��	���z~4'`F�1!���;mkX{{u���,�p���}n�$8g�oW�9��ñ�[~��흟,�]��FG��@�,��˜}����^˼So!4d:끺�45u-���,�s3��z�|g�
��yuea��踤B^m]p;���v	��U�����c,�-�t��=��#��4;�����W�����v�2o�娦E�����<���Oۺv���q��i�e���o��+��BbZ��8O�E�f�6G~��=WojZ�^p2�'�=�������p��[���p�������|f�Ȑ�fT��굦�k����[v]�}�1���X7��{tt�)��h���]�Q����j�z/S��޹X��թ!%
�����rf�P0R4l�t�+_~�YpZ��������r����+k'^@������3WL�nFra�V(�����E��o�Z��kG�и��U�F��뙨U��^t����N5F*�{Y͊��;5�7�9S�m-�};�/[AZ��R��v���u��&��>!v��^5��n16)�}��w[�ڇ�;�s/L\�E'���q;��*�NT-ko穭�o^�\ĉ�}5V���o����>�9Rm*(s�u��3�k����O=嗌��M�9�]�Y^#�]B,�q���ė۹���F
.v�����@��V��].�j	
��97+�M����n���Z���� h���hb�U,ŷx�BGӺ�V̬nRY��F6��W�1t�a�9��M�}.��s�6])NhbUΥ��]���2�G����E5��D��m�jiN���Pxlk+e&+���YG��������޵2����r�Y�f���ҷ���ӚN��;�(ީs0��K��9�w��흧�:]��Dr}Ɵ�>^����~��7�=���J:i>��+�.컁���Z�C�Fj5�W��]����Sle��6��+��Xq�ֿ�vMh��xf_鴹���j�����wE�]�ݣ��l^��)�+rou>�/�y�tZ�������u�8�q����0��D7��W3|�UG��{����.����}��v�20��T���UӸ
��C�G?^tTR�+��H����^]�F�>���]�o�S�G�MQ�}�� ]�Dc
��*&��5����}[����i՛���@�׮&!*n�.��{u5�X2���pe?������3lr��\݇�����=E�s;l+-��AV�P#����F�z����1��=�6���[u��)]tR ͎���&�wtç�uǟ<;ՌcҮ6�k�p����R��X�PuNb�f�f>�p�j:{�~���S�Ń�R˿AJ���uy9_v��q��oU���u����4z[1ka�ۇL!5A[���_Үb�}ohb�[�n&�[׹u��2���S�zؾ^h�jEsI���m}��FooԖx�;C�O�ٍ7�Pu�:��Qs�k3�.����[Qpo\d�+���kWɻ�jm�N�*wG+j����7S��Ӹ�6�k��gn\j���F��Q��\%��;��ǯǟ��b�՗��O2<~�Om1蒇����T�`V�P����呗ab��ȼKyM�=Vܽ3�s�+��l�����o�%�m���+�N�g���2�1�Y=3�\.t�jK�/��|��Q7_l���i�/�F�P���e���ф��g�݅ٗSm)�"���[*�s�fjN+�A�1��O!U��<* ��	�W+s4'����/�w�
zI.�eo�de5l����J�%o0k�4��������7�蝌�h�*z��RǺ�\��Qk����\Bgoc�62�2�������B_\�;����)����舋�s�x���jj��U��0��2Ҥ��Fs�[mUԒf�:��6����]ʔd��G4�&�J�7\���eWr�zf��u[�S�Vj��D���9�^����;�]L�6r׭�4��]�x���r�.�*��chX3[�,w,���K��n�W;��ަ�7���K%���cU����[��������
�-�CRn���p�$�x��`s�pE&u��Ҽ��>��)#����q�0�\�n��j��/[��]]F�'�����k]we��JC��Ӈd�����n�B������<�vI���8s�V��U*<ǤWR���{z���ed���_	�2�gS�!u��B`
���cq�{���`�X˹g:P�ޢv]����U��y�I��C�wwA��j�E�Q�����[7�.Ch^�H������J���y�̔�j��;�}��)o�cK$x���o�p�9�qV�2�k�Mг�j�N�z�3�����Bc�9`��Fٹ���&��s*1e���cVDcN�W\�gnr�d�f%lv�*,r|����%rd��z]����3��t��yF>����Ƞ;�Sa�w�]¤̕�vc�K���n�3Ms��W1�����8IXn|�¶�=���]qNj�������[�F���}�&�����E�G[�e�Yơ&^��=7��fpA�uA�
��<Af�Eya\�֩��JK��]��]s6�Wsu�ѬXv�&��7��,�}�0T9Ӊ������_9���c���Ί�*O/:��z�b��L�D ����Ñ��{���|X;b�l	x ��\h]�5Ʀ�	S�ɣn;x5��U��5��p�k�˸�X^� �δ`B��؁�G��eҊM��ȩ�K(�&9��6�b<�]y;�oR�c��ԡ�6��ƾ,J�(Btޗ��!!�hmE�G��Yx��Lr[N:�0�ˍ.�V�]6��%V�e��2�g3��IQf�S�˥c�ѓ��j�
���]�sGP��ͱK��y��̱V�㷭s���$u`]YZ��C��Nb�S�L�)r�x�|'�aT� �Id���r��j���G�Q��2��s��}�\��DamdH��mZA�u ��|��خpP<i6�dW�8�w�Vj蒮РӞ}ąe+���H���r��.�)���[$��"]����8ͨ���\�]�3t�!�)��ې��02�$N-Μ�����У�Ց.06S�u[�����U�����a��5Yv�u3\��iݵ��f�!�zv��;�j8E.첳���J�в�I�>ځ� c���4@3��.��wv�7g|��/��[���=%�\WD��;Z�Mvֹ������8��w�Q�J/I���)��Z��$󬻉{%��r��=�/2@���jo&�v.za6]�c1�E:f���g���"���x���Z��6���粦�9y��HQ�h�u12U�EmJeF!썝����Ƿd]r�Y\��KhL�7QL�r���G���z������2)Fݜԙʺ��	Fy�Ģ���t�Y���QCV�Vj�;VzG�*�.��Q��Ut�20$�,�ghC
��0�H�
.{ϟ�ϟ<���2����ɹU�g���Z��Y�ԕֳ�#�)���Ǡ�$�1*�ײ��(��]r��*h��Cb+e����$���F�.�y����3*j^�J'��]�E�mTe4C�FtR��]2/HCr�l{^�=��m��xPyHW�Zb�yU*V&�Be!
TEIrke&�
3)4����N�/"'%o���@���Fn�k����ur8�Re7o.�0�z��GU����h��N�hhY���b�k����ڊ�g��ڇ����s�#~����v�����Y��wT�n���	+z�����W8���x$�osy\�F��Ýݎy_%Gb[�z�*��T�tV��5�1��4���;V����x��i�Ǡ�w'I�|�Zީ���1� [V��V���v�go�C��q*��Ux��0��n5A�*oQGD>�w%��$$��=Y�XQ�AL��P�ۨ/��+��ު����O��s��T�y��]�3Ve�Ws�RZtd����_qKj����ʂ�B��n�ԼH�w�[]~�y��׼䩫�TR�ۻ��������S��c�v�A��[�Q_bP�i�q�fuE�l��@�r�Q���k˽�������nBnMm����W�{��T��l��K�Q)o�'ƫ�45R��k[�5��SZ���ݵ 8J�_t�'�U�<8��m6���=zbU);)���ێ�if���nELՇѴ1	'��h����ʥRT.k�2��[|����2��ו=�YjCc��g������%�i�ԇ�4�N�e@Hr��C�j�f�XѺ�I'N�Ms��Y=}Ҭ �O�'��;'��y=�����OEƶ-u{�S�����O舭U���''d���
cu�9���_J�)p��3�����[�eKJc7@1���i5�5��[���U���)�
�ބ�e�.����[wwc'qɉ����r[�9r�bW	�j�.Q_"�P��T+�+fe���)Z���m�҆�$^ޮO�z�"�BȄ�E���x�QoQ�yC�-�ĵ.�U�9��q]��7���T$�\�� ;L�q�݈Lu�eP�A��S��m�i\�w�}T]��ɨ�����ݝ�N���7_9y&1�����,��M����o�7�Fk��x���Oi�-�Q�pm��D΋���qڡH������v�!��|k�^b�1h3i�ܩuX�F!79�o7����(����|����X����e�Z�����Y8C����n�d��{Gf���{�])C��phf�����es�_eD\�-�֜�^�5(�91_+���ެ���X�{��E)��p{�<>��e�s)�;��My��S�ˈ��H�::å��N��qG�����哸�9�cS�����A@�����ߍ
���k�1\O'G%�sGh���D�
D�ǘr��&�G�1[�MWG/3��}P�|�"˹՝yu��t�슻������^���k��^���c~YoCu��G<F�4l�p�1P�l歫�I�Ӝ֏qK	�}��SH^߆(Ĺ�v&�<O�!^�Cw�8�\��U:����ik���!�2��=cj[���Vq;��W�^�V�y��N1�����c�U'#��Қ�+���=%���Er]���O�#� ����1��N����6��n�ݟ;z���Ag@�v5ԣ��k�;���L���V�>����
ӏ���ȶ��c�Ƶ�nw���{s�ߥy�Z�caY�Ba�.���/�[�ү�k�J����e9J%��ȭޞֽ��z�O=�����Q���{Ձ�(x���uu���x��v#�{��t���pz2�W��|+�6^s�φ.����}��s��<C�m�[��&�f�j��Ԩǻba1�`��i��y��o�"��S�jf�s�F:��=�8�t�8d��"���P�#ie�{n3�wj��5ڻ��so(P��j��i�[3 �iS�1;K��p�]�3� Wø�])v^F�3[��������?>{��M��s�׳�a4�r��ꛫ��˝�论��.�<����c�@�Cy�q�ʏ���Ԋ���X=b�b���l,�8'*�n���rp�*��|n�uã����h�ۼr�� ���]O����\�'v�9�]q��7�����~�ttV՞��]���eL�u����n��ۋ�@��V��O؞�͵�fn9�l��㷮�]��7�G�����s�F>��q6�����4�:��N�R?e&�b�e�3�b���_��8����^��:��e9�[��'��n;]C/1<vV��S�]�pm���*��󟯩U�n���M�6IS'��u��+�����=�z��w�Q�m�������hƺ�<�!��gG��O?VX��:���U�r���m6��dҽW�඾�;?A��"��a��C�xc}�����Ya��K(���;��^8[���e��am7d�Uu�}0�Xv3O+���'f4�uN̽Tt_\+��w|�4����V�
7Պ�QV��ѽW2�v� ӒTl���\=Y��S�͉�":��-��e]��ds����O]M�M}��RW�������ݑ�Z2�����]-�܁������eB�Fw1�,���N����_5�GrX��
i[�y_<gd�;zmigfL��j:y�.
`B�G�s�P;����M|��kM<��Z�\�hiafE��L�(�DΌ%5�!k��.̾)��0�x3'wsJ���T��Z�D�p�)�U�OG�Y��z
���c����{�;��}�#N�4��}N�7�W_{��r�Ü��7�`�2�mȖ�#��<���7L���lr�P�Mꆲ�yU�s�T�e�w3�L�����sV�*��\E�7�A��Ӑ�9�M��\��Ƣ�C��{�8��
����}y����f���r��#��B+.6��Ʃf�ז�_8�q�.��3X�ߋ�8��ޫ�yڟ�p�a ��Q�ܺ���]r������ᡓoe+����ֻQ�6��h��쮚Ls�$��Q��Xʨ�[I��[�^�H�ڱ���q�X_�E�U�m��9�i�v�l��!�"�1l�rC*ք�$\��9��s�jݹ�^�n=�
Vv^�a��QD�=��	2�6�
��[��
z�ǳ���?�}[�v�y�Wg(��n[z����7�Ƀ���'��=�|����<���i�K%�e���s��h?�'۟+ݦ�m�>˚M�B�(��\��ݮ]�I5��QW.'`��Vq����5J�}j0ַ�
dT�)}`<+m�<�����	����3��frW��AOV��-�C�٨�S}\T5A�5�Ѱ��)����%D�¹�KGJ����E^�}�5�W��9V�uSu͕�n��n'WLI3;2�G{Td����>�����ADIIar��^�Sl=�I��7���[��]���b���.�$\K5&�w5}wT�.˸Z�<Jj�w掶�E��<*
�w��%0��l����ރ��Yq�-܄w5&���m&h�����3]�-:D
M{;F(=�ƆؿoFǦX��d�Gj}��/*��	:w�j:?Y;�΅�g��\!��f"vz��Ds��5������n)1"ǘ�Z���)3oEr���N����ak�o���Ճ�+Q�!�w���N��:��b�O+�+�u��ذ���4-X�3'��L�{���L69����ٷm.�jh��.��ǫ_47��Iv0�h�Nt��v��h_���=��{.�*�<6���kύ-��Ψ6��F-sP��}�Yÿ�D��YIЩs���Ѹ�����D5.|�]A[�y���ǹ��=�b;���FJ��Z`qyv������wN
��KV-�z��߯�w�`Uw-{��P]�q8�\s��T�\F���[��q�\.c�̨-g+�SE�ݼ�����l��垛��/�g���W���߽��Ҿ���f�no��i�6O�+�d9G��0����֦�_7��x��\�轙�/0;�S���o������39|B��[8�ڊִ=d�����N��������m��5�m��Wq*.u���J��x�tX0�UnRx�w1Ɨ�_'�鹥W��
����_D����"'W(
�IuY��p�Q��z�I���_c���g|曱Au@�連{��eNjŴ0\c�q�aT
 u`���Ͻ�K��]w�*�LwJ��m>��}	��wO�T��!�@��8�p�ۣ�G����h���^��)�9B���-�W7Op���ӆ��(Y�KS�f�/�"�;����O�ԝ9�J�}���Bo;�r%�]~��f���?+��Ҹ�l.y�1�՜�X�5ˬ6�Y|�x=K��~i��\.t��x���uu�{�\F8�1��7c�+srxV�lU�!�$=���)�V���2�'4��s��;������ә�y����v7�s�*�$��g�`�ܝ��y�V��`3�����x��\�ԓ�5~��48��;1�"ި�Kj�t��gWa2�5��e���9\�ގ�ټ�Zvv�1-�7�UӰ�C�
�Pis��q9�Yog��W~�u�H����ޯ��w�.�}!��<�����Y'5(J��JG�Z�ì��ݮ/1�������7O<\2a��T����,Tr2*�n+D���[C�мt�����}K�_�ʣ7޳�x�T�k ����R������nZ�h�}g#�TR�]=�LR:ñQ1�"�L]�#fF&5>�4����
u����j[s4���z��Q.��A���Zuz����=o����M茬�X�,I��2U�˔2t�3Ƥ���vV3�@��Y��I\$�6�o}���}�.4v*�H�Owz�ޡ��������\�n-������m{ܤ��evk���D�(J��a��է�3m��ަ�����m���d��mJ�V���d����J�;[�5}��vS�p1�m>���%V�:�u��yFt�h�Wf:{�ܮ{��vD�B�/���Qu&����p�+���M&v���f9؅)��B���Y��%C�C�喴t����i-q۳RD�ӓq�UY��T�A�ˤ�W��蔏��.v�wB��2�s�h�]��!:�j��Y9b�oG8�H�<U}s�0��L����-�����®�Ϣ���7��ͧ:��y����[��C�[�����풟=�w�=�>�}�?Mз}U��ї0��9�up�S7�*��&8�jQV����s���o���'ɗ};e��_gЋ�n�$��Cj_�\:	�6�M>৚��Ϸ�#��QZ��n����f^�I��Yz;�pMe�8S��W��Wg5B���}1��R�ce
����uׂ^�q}�l*�G/�'��o���@v�rt�ʹ��g8W+i��4㏯ȭ�zz݅��*�^���bW.0��]`����ۺBL�Ʋ�J}Kq+퀅ˢ%�����������4�2�Pm�t_�O��+����N�.��Z�<dmwa���*ڝA��=4�ؔ�X[xs�^b��{���Q0�7��t\MCR���1�(+��ѩ��V/~�cn���8���7�v�žJf.E]�}5v5#9���{z�Cx��[vu\+=�0*b�Q�f6��S��[�Y��BK`�8��Fu����&�<����T5}5���c2�*��,�h��Omέ������yxB���k��͆�=�o��ieC�t��[�
��ݷ�.�мC��V��q;���WU+�cY6��v��G:Lo�{p;�-R�7��FA�/xԨ1;�T_%Im�p�=ۄa#��}5��AR".��n�ڋw��hX�Q��T�K�_5�G8��3�ÎVM����.e��L>�K��ת��n��#�BJ��s!.�[�D�
B�Ձ)���X�N��*��V���PGU�c)G44���ż┴����D�zW:�nL������ 扦Gi�7#޹6�I�[-+}h�/�Q�/�����Zî�¡7�9����ʹ����Wkօ��XR�)��΃�ͅ;���N�*h�YB�hۥ�N�4�C5��v1s�����e^r9����9X�����Z�|ﻃ5�Ҹ��!��neIw7�9�m��x��,�Pl�[�Β�������pݫ����g��M��Й\M�ζe�K���e�G���j>���nݮ<���;q��n,u�dƊt���K�K��ع�>k��]u��t�p�ƀ���ޚ�ͺ����ۭ�}�j,�O���B���'(j�څe!`,.������� 0�i�Zoq�b�e�;���9l:�>�q�]���v�¨^��n��D�A�axtf��ݫ��:�u$�L�\�L�wgH`k{pZ��\�ʵI���w4s��Rv�p@��/ ��;�0�9�z����oqrtmN&h+���0���D��r�n�,���m96��Yv�Z��k\�@���k�ī|�e�v�WI:
���.����:� ,�(e�F�h�-��wɱ�0��C���}a�X�ڴ)���/A$30�I� ��T�3M��1��zk;���h\�[���LN̠]g1��3]��C�8������s&���MZ���M΃����&��]����;x�+k���Z���$K�(w�ǙN=�'��-�ȣ��mcԕ<��S��kJ�3�RF�b�׵�&�KT��S��7;�\����:͘�*ݬz�M󅕧q�e��=��2���S�j�ӎ|ir�*�WI�'<f.���	���Z'b�K!阃��)q����S#B�
@Tަ)���:�ӨN��.��r�PJ�Axd�����h:���o׋Q���oJ��&�q�cܻ�V,��Jb����}WO[/4���5G��ݫ�7g6�B��V1$]An����5BQڂ�u�v��E��>��*���ʻ�O	8�e]�:8:��*K�-�k8×KO����]�V���4�.�`ӭJs 6�i���S]��q�t����à%f���)j�V,���[��2ku�r�RG*�K=ھV))�w[} ���x�{yY��42vK��w�[��8&�4�'>�R�/���.�n��
�Q�]ם44��S�"���V���qu�1wPi�&��L�quX'N5���W�nP�Y�.���}nrïL�9�qT��/�]�73�5n=�Ή^v�9R�a2gR(��(n?���.r��.�F���)���ȫ�9eͥ���M0-�-9���kP�C⥇�@�8��'xٲ�ԗ]�Щ�a\Z9
�B݃�6�m�EǤ��!:c+�A5Q�ې�m[�:޶�U̷&��OU��P��kZ�4F��52�vi7`������|?��Q��������x�!!D3Ѩ�:R[�y�> n]��QED^� �s��\�FӞ(�TI�
�R��ohG���7�
/��FBDs*J�e)s�j�2eAJ�M�i�P�j�����ħIl��!:AE�;cɲ� �	�Ј�/-t����X}�!JL�<��)uJ���B<�DU72Kr��+B�/�4�FК��g��B��{\n���HE̒�#��ELy�2 �sG��ٽv�z��]2�4�<�3�՛D�M�(���K-U���T���)znL�yE�Jk���#z!Nd�D{+��扅y*E�%�e�=�a^!�W��)S�[$��[�bk+l*jb&�zyTz���=�{d��UCʣ̴K5ݴi!ff�vےMcr�̮��D�T����±+�LP)+E��*![��ŽN$�4�$��t�^��TW���םB3Լ�9�^�*^Iaz�\���5�{nLK*Ԕ%QRJ����m̌W��ʺۆ�fxf_$�%�_#�����3����ώ��2s��Y]�][��V�Wmպڂ�ȗcJ�.�c�	�&�D�˕5�n^qO�b����lSc�V��r��t����?��5�W�QƵq�2i�5�(�@��F��`�|X����>��}r"m�}��x��9��<��Ů�ax,��ã��}���0�C�O�w��P{����5�y�q)�/����cx�k�q�!�oQ������7���/)*9I:v�Q8ڃt��{ZwE�D�[9{_@O1�`�tim���oL��׆����Sg�@�L���q�v��RRU|��k˅�s]�[�k�^b�ǭ�<aC��:����Ϋ�wg�۽R�|6a��
�d~�Ye����ι�r�P(U���}if�qx����p�.�ݝN��ܚ�یӛ*/�f���%��s;���>ſG�~�<�>l\����Ҫc�5�̚ё�Ӻ�D�R��<��]r�b�Y�1E�\�q6��fk��D�7�����Z�.�#�l9/C-�4.��g�y$@���t�(XsT��2*�B��qU�7n{_��+VR�7}L���r'(�T�� ��j��y��e�]��(��a��E}G�mv�g�9���ݼ(��~fm�&���_;�����9���t�ʦ�C}�J���S�nOaݣ]nV�UjU�o����hάou��z`��Q*N���HOLdV�N�S�����W�sŏy^�"������fW=�>
��8ן�"���{I��m5��Ψ�'��KK9�ݼkj'Z#�E���ik�)ɾA�ݘ�q�1w�[k/壦!_l�ri^��W��Y܌�[Ce,���4�wmA��+�`s밹ݥ��v��Ws/4.	:"&�y�z���FX!c�*�EF�Pc�}��s򮄸;�_{��3[*���=p�o:J]��f1֞B��b~Lp����f)��'u=�5h�eU�KsR�ݭ�p���SP��/!9&]y�|U�Q[XY��yot�|��k�����tr�1Tڇ�];
��C���ʓ�\�S������^�Z���S
����'���y]�
��"a��O\z�<&�oE�9����Z�xɕ�1�B,9�='�9V���q:r�;n����w;�Ά�v����w�} n�E��Nuv��֥Ǒ�f�N����_c�x�F=c�>UOby�]����j\*�t�׌���/gz������ʃ��/1��L��ӎx�_���v��kr����3WИܨ/��⺋z��r�����:)S`lk�+���l��u��|�l�Sˆ�vr;J����b�����R �e�x���ٮZu�ڜGw1O-��>ꆯ���H6��1���k�׫{׿�K<������Ӈ�n����y��C��.����0t����%����|u����žu�-���;�\6��v���X��l;og/��Z&�Uom�IlN���/�W%��;��ov�g6����Zf�F�ݍ!�2^�=�p�27�\��.|�\-���}�Ns����"�.t�t��W�4cr���{��Jzds밹ݭ
�QM�"C��:j��>���J�5�Uv�ڂ�U�gE ���ĝC'���Ż����KUo���][YY����妯E�	�5�B2J�m�#z��$�x����ڰ����Q��zoTv3h��.}y��ܕՇtt���M:�����Tپ��o�y��M:F�E��ф���Z����l���v��$�6ֳ��{�j�o�j!N�ph��[�?"�
����z"������⚤����[��w)&6�o�ô�A吮!Մ�	3�������vs.$��l�ͧ��B������|�^޺P�SN�Wd�O�D�"�Pɬ��,k��E����.���oL�-��N�:��J�L�RT���\�{��̷�z �����hS�R��?K_Q��L����U�mbK
Ev5����KV.��#�=��7���s�j�y��Ǐ��r��E��R�ߛ���?=���\�%�8��j�'��@��Q���K�g�O43�R��OS�N{�c=���Q˶������1�kgmv�xoO,�y�b\�M�uY�_\�문���ڗ��.��iu��O9Ջ������{}6�D<\t��LP�<\�Ucr��ʍ��f�����짉a��-��U���+](&���V��U���!�5����3#؝%�O̙Վ���A��V��`�N��얱�8�D.x�-ǃr��E�*N��cc�R�/=��O�nC����cYq���&���Q��e]l�ll��}��-���Z�T\�1Q|�B�L'ΫkyH=�g-Ӭ�|���]k݇�&���+�6�����T\J\*��T;OW7���o��k����{����[m�����A]17�$�\֨�3p��j�_v)�t�Y=1
�����p�v��1N��Q��Ҋܭޠ�3c[[��lv�j���.�S�x�ֺ���s�pԺu{[��k�Z�(�=FC/���S�p?Jחŭ܈Gr�&�ྦྷa�g��X�J:jpn�aX���ݱ��%oTA��lJ���SKC�N�j��[u��*tw!4�j�z+�������L=��pV�4��3�ޙ��k��8�Leo�cb��'e̕��}e];�+c�뢷*s����*��sU���<��1��<Qe�}��B� ��i��+�WV�k�ڠ��-�sx�J����6q��8�b���Fg\>�Q����H-z����]��+{��jK-i�ʥ�iQW�Wd��b�u��i˭x䝷���O���ُ"<o�7u(�B�n��;�S���H\C�^[�Wu�YpZ���S��;����^=�n��V-*t��Ϗo�G�K��C^��CX1L��o\(�R�����]��	����8��bߪ>���u�6��7�e���@�<����Wg�V���}j�8�h����֓b��^���&o+4.KHK�m��w�g�\;r1���{�߈]�U�gy��ǈ5;w�f���V9p;��s�k�[����)���v�A້Q�:�`&��U�|o�� F(�S�u�2R��z��)���*���������j��ge�k�w��Qʗ:M�V��B�?B�=I>wZW�8{��FӦ��:x��n�c��ÝmLv8�ѹS�0�V�ˈK�����Ҩ��q�1�Rp쨻�B���8�w�<���e�0!r�	LWL�9��\�ֵO��s��ћo%>�X=q�=J��v�f������/�|�rjy�ؕ�;#�Nmu��x�ެ��|{q�݇�m�޽�ٝ���v ����l�tuO�[����W=�9��;�(v�n$m�_L7�!בʝ;�ɩg1P�ItÙ#ќdt���u�d��t�h��W�q�*{*�^s�U}5{�m�2K��������OT�Hu7��-�Lpϊޣf�?g5����O�'J~k�W���5���KeTН�W����TA��]��me_�<�o�7����>~���ar���}w	�;IK���'�C�[���|Յ]������ּ�^�l[�Ji^v����wo�^��\�k�b�a���Y�Y�⯎Бh^���~+��`�	S}�	�'B�^��l�o.o:��*��Z6�h]d��h(t��l}OK��xgT�[Xvn*��~�;:���|������M���SmC����$.UG�Z2q�;,���8�ƥyJ�\�O+��ث����ڲ����m]��V6r{+.�žᕔ��ț{ȟJK=���'�}��{��y����[��N��iQ�ֻ5sG	��p���L�uOz�m7;���^��L�q]`_y� >6׹y��7�k�,�4�aӽ�)}�%LE������D�r�N�wk���f�0ު��|�c�}���U�]�V�X�����X-p<fY�����uhI���PJ�B�J-�{y�M��)�U�ui0���nF��K}��x;�E⛖T���xA��G�VmԨ��2/���]CO����1��S�oe��Z�t��p�ah�'�T#�c{~�f}}��)�j���<jq��{�f���y<�_8��V8�����2��Uӝ�ݵ�*zj�����yEs��Y�Iy˙��Wy-�������LS�b���2����]�U�;�v��p��67�7uNve�<����O�4sO!�҄Q�Eo]K�}9O�Q���oC�y����b{s.4��ϑܤ�ڈo����*�����s��aE�z�;�����6U���wo�[�=}�ϣ����6���bg��$v��p}���֦�..@p�ۢ�ѥ���ޙ��h5ܝ'AȎ��t6M�)%�VJ�.�i�;�+X�·* �:��x�~�|��t�V��&ea9��O��yF�m_T�b�+B��A�:��\JF�;����4��r󮵄�t�1�e�I�_RjA�J�]Ք�46]�Ƙ��Wv�m�:�[�隫�M;Q�λ��諃�Wv�d��F�]�K�.7�sr�eމB���^�ާ7���Kw�{��P�j���_ktWeA�u��45��m�2�����Z�g-5�&"������ه��I`Ρ�;ɚ��O`�<�T�X��Q����6�a�,O�yHk�'n�'l��n]��}׶K�7aT�M�;� 5�T$بx�5�Ӽ�?b��C+w�Ϫ�E|��"��Mɴ8�ڬ���D.�[8��Պ�5<�f��3Q[Xwi��(�j����j�n;�אx>㒠��|�|����d8q�s�$`]�˕�=�,�����\��L�c]J�K�wׄ���[�yCUGkpk�o]�Ҽp�qŷ-D��;�%m��"o
��\�ң����s��;�K��������W��K�j⩼��j�����gk1�vk�1�?V̎]wv]��O�1W��錃�*sސ5��]G�/{ٔ䊊���cb�wư����č�r�3(a3�_ڗI�*p�˞�X�gt�.��5��^`���2A�6�?�Kۡ�S��G\�K���_<Fr�e�wY��m5K]�����v���V��4��7�ϛnt���)�����Pfqaf��2s'��p�P+�`{<'��I�s	��H��}^Ӌ���Pt_7^G�y�Yح��N�Sʗ~ɱm��~�3�U�+�+ 	��OKe�z{<&'�j����△^����MB�kv����uU���4����]`����<Ṉ޳6�ܨ]����+3�\���l�H�E����#|�����+���3��y���s��ǰ\�5����;	���6��M��/�f�yv���1~�]>7�>��gK�{3#���Qr��)<}몏l�p��/Iُ_�D�dQ������n�?K�2��Z}d�7���Ω`(�מ� ����:���qS'\5D��5Y�;���%�͘�f����JGn'i��ɭ(g���΀�f���u�/۔��������߿����d~cGn_
�G\\,�n$�>YP��챿n�O��>���c��3ê�3�h�q\�]j����k�^���W�Hh�v��JS�X��tX�}���L�Xl�}��ǲ}������[��F>�s�>���z��K�}�����`�zG[ J�,r3qR�Q�Fq1�BdE�h����`��B�R{�kBʷWFn����w`�D�L�����:p��k0�q"��9�hb�:�U9Jj{N���r��z�R������.��m���X����s�����Q��|��]����,]آ��O��J�o��Yg��#Hy4�e:�O�ڈ��-ᡝ,�K|_*D{�=��1z����닝7�'���m�+�ț@��2���	*vo
� �Q�SaTcv���k����v�}�H�W�u#��-�ۮoW,�dB��X(Tи��zEI�V�1/��cpY���WF�߲�\�
�Գt��#��u�Y�Y��YX{Kn�9u\�V��\���%3��K΄�e���4����H�C����S���q��}okz�m�K����:���v)V�� `V��̻���}Z\�:�9�I�f�̬R̖��`�c��)�gd `]�Q��C��[j2+�aKݠ�� 蛹j�i9Zh�A����Wؒ`H���`YˮhҸ@Z��;��t�-W"��Htx�� ��f�WjVV)�WhB��Ǭ,�K���yh[Z�-�LL];w=O��J��<d4i��H�l$J��H���������ʲ�mQ署�$w�vC����u9}8wov�i��M�%,��Neu��9�D���b�,��;7J20�5�r	1���u��%����{>�H�+���>
=�8J���2]5��.�h�*�d:��ɜ�ю����hJ0QKh�����`�ή`�;6*�e��)����,�W��
7�B�9,��^�������FV�^�ؙB
fx�f9\��^�ӨC�1V�����3@K-THۀ��J�lf�:��T�A��}tZt���u�(C�{"Du��Ѝ���;*��Pׁ u�x1��v�^�f?�h���O�����eX2��e�'��{;u���Ytw:��l7����'Wd�c[�ڻLZbѩ�,�8¬��)A�T�a�<��N>�Tp��ܬ�c�J��'p�4t-ɻ�
��e�g�cZ����������ZPW���K/�*+AK�6�����ŷ�: �Zp0�[y(#Vq	�wA�T:��vG��o��o��{�Pm�7��ֱ�JK'w1����
}���*��f�Wٸ椮�t5hb�to�i	����:����]NǸw}��	b��f�9����Z�D�o&V]ʘqn�������IG�6�k��{*��[o�O���U�{��(�[@fd��p��� �#���wWb˩��L�n���Tۊl+#G��xgs{+��i=�ouG�C�
�K1�{N�	.�[�����Y\���=���7AT���%}&&�b��pM�w��s���G]�Y��8��bg�7G4�2i� ����7��.녙������u*�}tX�a�GȚ�h�ݸ�k��3�O[�g�zGlv9v��� �&4͍l1B���Eg&�����m&Q�Y���i���綕����<M$��4�*G�ع�-۳�����6�١敽���".��kK6"�XEncF�j�ؽz�g�����W���m����(�j�6��J����ѹ�u���d������a�ү]����y�Bݚ�)�̭]���m
.��R�U���Ս�9�.fTjHm���C
�SJ��".�xecN4��#%�ʕ�&�2:k���sh��:�T�ą�$�#k:�Agay�Țfa�H�3���t����p�����QT�6���M��zb&"�����"'RɌ�r��IƜ�<¤C�M,*��Y!t�S����WL�W�\�E#̮�\Vq���"�uh0�┙�^je��-as4L[��B��I�Vz��]fY��#�E=��):�:yxT�؂���X��
B&{��fZ�#��f*IQ""��b�d�)�U�s�t��t�
,D�	=MZ��C�9VҚZJ����U#����i�oޮ>���ە)��.�	uU�F�h����oz:���HJ��K��R۵*Y����2�J�=35�d{�{��@Y�<�g���Q��a���>�#M��@i(�����L����[��m��Y���;�\+O"w%�ڙ�������C������z���gn�op�ɪ���~,����Pz@�u�Q�Q7�|�>�����L^�'���aR��7�{{z��~����<j�����LL7r��|W�a��O��߶�47�'ʤ��Wѻ��(�w���^�o�g=rC,� ��\L��j-	�}>ä�w_��"3X[v{�d�sw��q�}ܭ�<��x��`��z� w��"���k�9�,uE�����{"�N�q��J�v��vT�h�ze�O£��U⏝�r^P޺$�3��χ��U:�Kw�C"U��N�{�3��T\�L�ϫ�T7>�Q���^71~�;rnf=��Loe�}���������L�Oq뉺�Y���d����;��eKO�x<29����3:n�>[�"r��5ྫྷ�ޡ���p��bV��۝�~���K�l֛�u�f�*�_�vW����%��w�s?.�2�v��N�6�6�xr?�x����ԡR�.�T*�I�^,���/�5��դ��ӻ&��&u��휚�ss����N�A�X��53�pd����@�����V.�w�I�.����]d�C�u�O���BRݝl	�#�<���di|n�r��䨎�%���G�kE�zOl��Z;s�纡����\�����Y���|%�����Z�W�v��>�e��+c�ǖ+�p�Eh�Y'N�D��9E���ۇ�,��6�����mO�e�s�k�q���_���l�v�\$o���-��Y(��s��(��B�zhՎ���	����ڱ��;��V�&r'�X�n}~��~>�q���W<��+*q��G�w�.�=>4�&�w\��>�)~6������py�k��zv�;y͹�1�u�wN�f�z����3�ON��`MO#�ovS/#j�z����d������h),�y�S�*�#ه}���Q��)��9���ר�nQ;�x�ϟ\gn�H׋�:,�l�g�In��9�����}މC��D`�z�~o�!\�s27�)�Ez���r���~������Q�u�h����>7��u�RGޜ���	�WN�2T�� ��L����f�vz��I�]z5u�����z
��2�g!L����n����s���%{$��e�Ne�D�s�o�7�)���&}S���.5w���
wE'C�;�f�#���JF�m�E��M)䡫�ƴ}��q��ظ���dJ�[�J�^[ �jng.���p���8��Od7V��m8���[�.�hT[˱�C�[ �hv��ei��A5�\/i�Ss4�_��Vz�[�v�~����3�n9����N�b���f�ޭ��Rшk1g��Z����'�a�Q$>+bn���x�*-Nɥθyk5��U��m�U��;���F1����5�;)�{>���z�*��w�ud�}9��7�x��[}��'ކx����<�`xmQg�C����n�xbH��Ig.e��;P�o7jl�OH��,R��L��=�v�7��y߯���(��W�}�e���h��I㄰���;,b�f�x�z}[��������>�������z�>nw����o�U�[Tp�ˤ���E��o�K\���+̗�
������6/��P�K^�7���mc=�~��#q����;���ٓy�_�ڂ:*��hǷ�IF�튯Td֖.2g|n'] �%/f�s�+ث�<V��=��cs7��y��un{c��j1q�%#q'�O]S L_z����革��ˢ�n4�U�u�q���7ק�μ�z��S��4d{�=p����O�Sq5
�^'c
e�;�y���_��_���$�)ԙ��Sz�ӃC��[�k���װeZ�k��#/��^&;2�Ӓ�_�D��>Uc���#��y5j=5�F�W\�1&bWj��;1�6��u9�7��L��Id���]KY�!L�XUȜ��{h�4m,%�9�p)M��A9۪1Xx�LM�z_9�Qc�Iƿ(;���,����xhs]HSUA��!���w�~� g�X�U��ϳ\�{��~W(:3	�hG�c�,�^����Q�ϩ��o�x��D������nK*�"\����O �8�F'K���DV�
;-��x�}D'�\Q~��=�k�c��S�ي���B{�\y�I��0R<`�t�@gì�S�q��Ǫ=�Ы�U���mqS���K���wg�{k�#.��{ﻳ �r�"n"K�&&��LM>�i�S�|{Y������VBȬQE�=ɚU�$O��;��gz����?	@�L�*���𘦧h�.��#��lmz��;I�PC��+���Mx���v|U``z�����j&X�Y�u�n�#K;G��k�
O����+�l�TZ/O��5��3,�{΀�9�K˸�|Q&���������|�oG$D�k��Y�ܽ#���z�u��"d�Ζ=~�n�{_�����u�z���yG	`fU�Y�g�؋���_��M�p������/��h�q����f����ک�Q��� {��^tx��E����Ѐ�Ì�u�}��f�v�����oj�^\ ���-@���yj꟔���(���fTY;�c|o��\0���
�/n�kw�A@ӫ������M�w���GO����>�V��L���r�`B�e��^�ٲ;r�c�r�_m�Z��G�������o���ք+��	�7'���b��7=5�s�7��Ṫ��G��1PH6W	�R��H��d���go\���?r�l�yܫv������L���5�������v^��ڜ��.0���>���]���u��hp�-��d���Kzn"���w�����j�G�w'H�n};Sވv�"��L�t>��9�T�|��`h�{�g��z�]�ў�p����*�ϖ���Bu~��w��{�#�o���DK��GW��F�S)Y���V�)�,�vbvj�0�2����o=>p� fL��S��o%����B�i�����8�zV�����k'�mA����:���EW��0[5dS>��Kex���|��T�_
	��
��®�6���ZR�!�G����#j=��2 �5
����&��Tb�
�,9KGٟC��n�z����No/��׶�{���;��@�Hf�rCr�0.|Ù�j-	�����5�^�t���}%u�ϵ�ݾ�=��5ϼ�p_z�_�m0V}�^��{,��Q;2�"`1�ِ��ض󢪝1օ���aa�����b�[�s��ή6���u�����*[.�g���ǝ�2�n��)�v	��Z����Д�3)fo։�x�f�W0�X
^oQq	�<�;u3 P��o��� pUui֜��3�+�	b�8Y�r`�T����LZB�������#���~�R.	�5	�Tz��W~8}���;��ߕg�|OKm�fw=>�cb�^zF�M׆�m���P��ީ���o޳Q��Ʀ:#�t<�"^]ǡfO�{ד�7���/���C#�4/<I��Q/ğq���
�wK���Q�끕����Տ���ͷ���Vg��)��.kg�ϣ�}׃�A"��B;�0��R�Ǭ����O��f�:�F��3��:��s�ﷶ���7��v(y���=�qZ;s�纡�mV�!m��)c�}����c�����+9���x�(�y^�/�з�+E��N���3�r�UX;G�E�'#��^�L审���}�^�q;(����~�O��9�ݰ�p����_��(�fIN��&�9);������\6�Xw�;��Ȋڤ�}<���~�q��T|_���F×[Q�T��<��-	@�Q�}��R�����1s�,^��RǮ_��φ��ё�:�S�I��ѹ��Uw��t4�N��ڌ�Q��lL�Q= w�*�S���	�_=���:�>�r�Ez+�ҽ	hH\Nw�6������ӭ���b����Y��������Ƕ6A�CmF'.�*������|:�pE�F�.�i���e�0��Zhs����iZd[�GH�ٺ���_My	 Q��+����E�o.�T�I�]�ڮ�u���:�TR�u���~���PǡOq��:�����5�1P[�M�^/cм�S��)wmUM�w���}��;C>���{����C�z�(�H�JY$6v)M�^��,�������̫����y�(��\U���r=�;�8:�n�\9�%\�����*�u#�xu{6:�^ly��P���2z���{���~����T{�@;�e����@\���3��>SAz��>��z�'�ڒ%�Ã�]{�l3<6����z��c"���L�/^�����u�b�|��Gva&��(�������}q��X��t��=��φ�ϝ���L�M{4c�ՙ�6��л�'���=P�T&%a�/��n����0���z3]p2�Og����v�u!X�#E�	C�uE���u#��nǆ�����%���;n �B�ݨ{���s��b�Uom�f�"�K�|��2g:� ����;����w	�{n�\>����t�̰���'JU�����z/��ێ���}"���y;[6�_����|:���x�<K�q��g\U��t����U�}'����Rx��H'N]��(}D)w`!����X��2f�M�ك��S�sA*�����]e��bgC�M��sr��N*Ӑr��%��a9֍鮛/1J���iSW[@a�z�[}�����4�㉝�T���]Z4�K�������Q�yk���ǐ��i#���d�{�G��H~�x��ǲ�SZ]�O��q:�o�"/X��~�&�zW�>Ds�*�z.��W��{�w��ވ�y��~��_�����~Zx|%����J惘?��x�unϢ������u��Z
@Z+�vW��y�[e��)��� ��S3��+n�<�k���J7��{��.��G�=�~��s�w�>���1��=Q�A�ߢO�SD�0&+���u,��O��^�w���z���u�6r_�ǲ8���}��{����Z�3�9E�d304������7o�<Ww����5Z�י�luG#O=�ȇ�l�������q��x_�䲎l���1ɒnwux��9�O�*P�鑇��N�=�9�K"�_�#�B�g#} lD/��m�2�H�>����C�� z:Y,
=t�Ws���G����3s__.�u9���F(��+����Iy���g����@sͻ��D�I|U�L/W�H����:���v�5�n?rT7N���JY���;�ݦ��EDOu[8}��g>�V �� ��(��|Q����tE5[Ez�_�_���N)G�����aH�l��WR���%���K���|�ܸ��ޘI��"��&�̊���P��V�I��am�٢_��RH��n=�U���$ax6fQNJy���A�]�"�hN�#��n�C�b�z��n��au�����_''���c�ql1��n������޸��]�zF��/Gb����|}G>���n=�5�y�K7�<�K˸��I^$+~;�_��0�g�5����ͭ
���t�oK��t���.=�K�e�'|F����{`s�o���1h�����q��'���N��a��X{�s���gSz� ��Wa(ʐ*T*uo�����#�N]�Ez#��t���{M��;s��\d֔/=5��:��j�;ʦ����+���;���zl��r���o������:��`��q%��ʨxk+i��&w���@�2���O��v��� ד�����n��]�<��]!��<�Rd�$1geE=��똨�D;ʝ}Y��e�C3�^�>e�m�/��w��o�{�����_���p��N���%gzR�u7O����X�2����q�EO5�l�^,[��ߞD����r<S/�{%�V��ݬr�{q��$2L�w�K��,�@��'�WT��9~&�Pl��n�+��h{�71��N��~�y��d�4�����e��Vb]��$�~)�I� k�Qe�{R��z���f���r/{W[\�8��y�m�7�EY��EC�cmT���iA���s �3u�C:�������o�i���V<��ӊ.��s:�(v��ޠ���qĢ�gp��N�/�p����؎Qe���z@�q^�PKe���O���U�cq�@V�����s�D��v���t�>s��O޻yg�q��\LL7Qt��^�gb	h�-�z���*�{���Z{{�;��օ�WSG��@�����n#=�@�lR�x��Xw5B\���yu�m�����g�9��v��a���W�����-�p=Z w�DO��x��a��u��2���}y�����"��ߣ�W�E��y?
��y]���<�DK�{�D�����������gE�J?���"�F��G:��P}�}꜇μyٸ�S����b����M��x���_X��g�~8M3�V�>��R����.�tzMf��fҶ=o�x<�^P��ߛEkB��+�z7�����ՏC�6c{�V9���[��͚�f��3o=s*CO|"�0�]��|Ⳑ��}���uy��t:�幂�|�N
�Iݒ8ra���T?w��vت}B�3��*	t���W��W�F;���~�e�<���t.h���p䤼/�'�V?
���O�&�p�����Qv��J����6�`e�06�A:�E�*Lv�q��N�3R�	j�����.Nڼ*��j�P��n�}4�y}!Ȯ�(�<�
x�_|8�Mr���^K��P��}Ԏ�C��3���+����P|{���	p�wgN��v�1�[���-O�-TՔQ9�ԗ��iR�I06�k����zApF��Z�C�j'��*��.�Q�77�3��n[�SV���x5��aTǖ�b������q��S%ʼ��w	���Q�\���9M8�-m�c�O�{viX�Q��[f���,)�R�g�^�})�i�sw�ߍ��w�]Ə:�!�v��:z�ow���H��_3���M5�����1�y��4�Zڛ򜯔�Ku�&m�i�e��Q^&n���u�dX�7{�8�n����-HMs��6�Q���g=�ۡ����xA����9�r)`��P��3zv�qM�������F�̼LD���:��/�ľ����N�K��v��jl�EY��lDN���gG��,>0Ge5��#H�]� {p�̚qYw�`b
�%BK�Ux���R�d7��N�q��_�2��P_SQ�X�kf�F3Y,�٨3s�$�R��zK�k-��⢫GZ��!�4fWu��Qu�Y�[�e�� @�W���%�p�q�p�j��R6��R�j�����ވ�q���7ʰh	�0�yC�6�"���tk�w݅m���\r��Y��x��޽gy���u�Ub<T�[�k�F
:����FS��Dڶ脦<�e�[��%�0�(�ֻd́8Ue���΅��7�'�0Po���4����{�u���1bͷ�J|f.VPL���ӗN�(i�A|��<7k%,��&%0VZ��'J���P�(L�h�5�f��侔'43����;�ʰn�u7R��]�:�8�C�I��8]���� ��pUy�| W�6�;YN��6��n�ԑ�a��=��,�+)@Zwy�y�O�jU�X����[}�	MК�{깧*�ӃU#���S96�r�c��Hi����|�[s-��y���I��Xŗ;TDڢ��b�Y�M��Eʾ���u
�1��
�Ze���,����g`ɈШ�ohxn\��e�*V�2x��痌�ݫ�9$��@b�D˳d>W o���Z�ĺ���Ғ,���U�D`b�D��:�tJ�nN���Pὲ�ZWT��)�Έ��2�t+�7*�l�o�-�o�e��s�T�Z^êt������K��ɜ�+���f�;�&���{��#x^*x�.�m �;XmKk�X�A#�n�jص�v�<�z�X�v-����fɆ�'�*_]vٮ	'I,6��׽�G�|xj��Z�qW��tʰ��n͒�T(h$�޿^�������{c53�W,C/[s(��2�(��WL74�#k�̥E4�<���4ICt��HJ]\�©,#\��QB:u�"��IY*X�e��$G�������S�b	dB�!"�	&zJj�cN3�Cu�00±t*����	��Xj-mBL��DU*�%R�,�1T��M,�s\ҽ
%�QȲ��"ӹ���E(e�������z�i����]�b*J^��}J<d�zYiD�$ֵ��ɷJ�0�9,Q(�Tf3J�{XG��6h�*j�`�f$�U��VV!.�d?������(a+E���f���W���Ib)�Y=��A0�$�(���RR�4KCW#H��LP�Ȥ>�)-1%��3��K^�dG�iI�_k|��C�>�:ג�s5����
�#��bK��àN�}noS��Tk^j���%+H�^���Bځ�f���N���G�+՞���p����w�jdj������P�p�MN��ݴx�F�'��R��i��}98�AZ��s���j�9<���~�q�t���wOR�.�J]���� vҷ���(��@�j'ҁ�`Y�7�me��D?U\�3���b��ES�ri^l���t8�c�q��c�2&xԩ�uL	����7S.��܏fm��򇣶��yw��>Ztz:yތ��K���{��:��/�¸�B�@�/��"i�D�[�:zf��U�KBU뒯�����,���l��{V����W��Q#zҮfBE����c;���Z�{՛�C��zp{�<����+���^��G�(&s}��N�l9�%_�۽덮�����D�����Z��f��������*�ֱ��9ģ{���dmWc�+˪�������j$���&&�T�3v�|xl>ӹ�p߮:�=�W��)�^v+�$�ϲͩ�����E��g�N�ֽ�EC>%R_M�>���1\rOb�rᇎ�$�2����1�'<�e�� �I퍣[�h��[��TP��d;]z녿i����sh%�-u�}��ʼ�hC�l�|�ݽȕ#M�[wm҉Jպ�]K ڽ�������U{����c�+�彂����,�����zp��!�����\v^N�m^��7������n�Dܬ=.r�O�J���b߹�󝜐=P=�A	��`���7P�'p���t��z.EE`2�&ccr�z7��>��+ޱL_:���9����xbH�^��_�2�m��^;��ת��Z������J�﷧ș�θ����/U��A�_{����z�0�w���:�GS���A�v�ۂ���n��U�������X�ͩp+���ጲ}��~������t����ٴ�\'���G�@�����a�+�|(-r3��z�����>ٶtT�����ϲ�-6�VN�/���Q�kMtdAG��`�7�f!��&����N��o�v6��{�9ƪY�߼��ޜ��\�@>�$v�h���{x�舂�RW���2�Z�?o�����|c�/�Z����+�0wճ��Bn���^��yי폽�������A�茑=5Xޛ��
��L�}�=�z��^�_�{=<���~7/�q��w�;�w����S.R�nK/����;�{>�����k�;���oJc%2��[��?C>����Ӟ8�~�s�y3�,]����N�}�i�Ҹ1v���c�r8����M�]=�G ��,'�pi�ܲ�Tc���Y��[\o9c!�K7Eт�XU��lH6��Ku9ל��:�f����><�<{xf9Gwu!|���y�8?��~�=�Ϊ��+���=㭪��:�W���r6������l��d}N���Ϥ�p`�}q10�EңD�u�����]Lz��ا)�pz����ĜWR������S����3ِC,��*���^��LO�������k�י��ڕ�o7[������Kc�樨�|���z�'��<	-��3�����\��>��f�PɽYkܣV���-�G�F
�O´\C~��r�9�t$�D''�%��\:j�c�\�	�w�Ӯ��;Ѫ����M�������o���Tc^�g!���n�=a�kw�<�q�����z���S�%�Ύ�h�-ͭ�'|k6X�3p�X��ٙ^�.x/)<qy7.�׻���髎��JL]��Ѿ�p��_��B�����'��^N��q�N�ŀ�z��Y;�zb������.� sn�O�ڃO�ي��	�$4sgj.�}���֛�΀�_������og.�X�@yF��$_��O��z�u�e�B����V'0ܗ�ݕP��������,l��A-�^�F���u`�`�s�n�����uf�[e�O�9˹n`s��>�g""\�U��qͱ�;_L��95M�	��GU?�8H���㕊��|_�`��I˝������*Ju�3�}��z���>�?�uP����~�^������ý>�CGG�i��|KvE^�S�'��6!gI�n��L�R������m�Ωy[P���w�����K�}�ˍ�j�g��Q]�^.O����U����Ox͍�PZ��_�<�����D�Tz����������ˣǸzF�P����Q�B�D�u{����늦(/�<+jd{����F|�8ǌ�W.���5N�(q~�>��|n#�~��B9E�����-��Q�[(�
�����7gk�<��+/�!~A��K(ϴP�ws�29�)��������8�B��t�7WJ�Q^��M<�)�G�w�iFt����{=P�=u�h)���u ^����~�"��\�+���x�Cw�W������v�r��z���iV����j=�q�7qq��~8}��Y����6�|��n�53�!ۚ��j�g�o}�j/���S�o�}��u˥ǟ��{f|}���9�J�uov�j��}���kP�P,x�a�Q�1����g��Qs�2)s���n|6����m�u�sхt������zgn7U���G�_f9<럱�呂{�� �s�V����u��^�Lј�V�L��k��i����i�&���7�R�E"���77vV��1!�x�!7o��v�GxjF�ynֿ�嫯{�$�s}J𱏶{��u��I��^�r���Nd�FsǮӒ�����0#����MB>'��������aW���5���J��uU������wy+3�	�����q��{jǰ<�"��U������/^V銋�������ޟf]V�%3����[�ok�S�<�-~TF���]�������/�}��R�^�uq�@q+Q1R�w��[�}��W|r8�������Y��;^�jN?Th�����Z�:v{��^C6����%�y^c��}t]}u����7;,s�z��_��߶q���޸H�ڨ�%;��䜹�w8��!��!�S���U��ɠ����]�r�Gzhm�7���S�|l�����{�~�W/���!��<�����r��}d�S�`��Sn{ŋ��im�>�N�:�I��(��yi�^���=�tz;�y���ϴ���͏=��,���j$��\ES�#�v0�_y11��P}��fo��VW�}���1#'��ў������Y���&Mu*����SD��>�h?f���[���w��o��a�^�{�
5=���l���q�􁃾����䎨wJJ�=�ԡ�t�^J�u���c!%_3���,팜����e�bՂ,�������cRt��ő�oZ��l(��I��p5��R�)�:�)l��]���U��v`Ըi����S����Gz��YڡD���q����f}u8��S�ë���e��8.pu2u�<8KKp���w�R�{����}����*��^�����z��W�܅����TI�2��|w�&� �i���«�EO�s ���������W[�ȃ��%~sGc���k�ԑ9w-��%�EC�rQ$>(��*�&b��u�=�ꇱ=�{���߸?R����2c�u���;>��yYωD��[7P��+���NI�S�׷�p��⓫Ku!k�zF�v�N���X�y�򜗔� z�* ���7P��L-Ǚ�3�]�-��j׺N����j�<2=B|�K>~�������2���(�,v]^W-���=1:1r�G���*����ֲ��f��q��3g\1M������9����^�]���p��(<E���u�v<d��&P�2�/�W�_�TV�J�^�+��U3������TyId�'�"��-��F�\W��l���7D��눝�2�&�����K]��5��_���_�,pq���t�s�n�	煏Gt���)�Q�	`��rl{�*�����d���s�x��.��_�+�ɚLo5�~��L[��p[�!D�O)M��>&;��W�1�u�ɓY{ �R{!�r��M���q��6����vR�,�u���r�d ��v_EO{���7���u�X#�:)��:��D_n�flvw-Jʞ��T�H���^G��<&���L���(�����?n��3�z�խ��Ϻ�Eu���Kn|hﶪ������W��G�����|5|�������2&x��t�cc)�]e������@��^�G���?�~W�����;��{��j��=E���u�a�����w���o�7���:@Ͼ����J�v�\K7����=)dx��:1,�볠Nxy�ؿjPwT��^����@H���*�U
��q7���wQ
�x�%?RF*�m�y�Nޟm�R��i^�}�4���qp�\�/�#똘n���|:͕=���Vw�n�j���yi\֜3Y���b��x����V;�#ř�%�F/l]"b�O��k�~�ڑw��lN������ևq�^e�Ԫ�p�i�~�`
��� �~���|U�����	,H+�5v}����`z.���>���f�}ڼ/�Ds�_�G����*B�I��J�u5s5���Y��3c�o6�T[��Kg�}G"�q����S^�f����s�yw�8����u�^����_s7���o����[��E'a%G׽��#�<�7N
��R�=ū-�Kv�_{�o>��v�$�]�t�u�i�N��;Ð�F4宖k3���f*s�j�fv��{���I��My�UJ4p�9��ݲ��dz,��nn|=q�Z��gu0��qc������Q��O��Q�}��Gk���g��w�gb?2��2�')�ד�O�'Ei�s��u0)FHr���_�c_��B�����{}h�:<kݕQ�p�������ۉڋ��iB��ZF?a\F�a�0��Cފ��A�l\F����ɸ^��"�����j*��7%��dUB�Qx����}�{�Wc]��td�.�G����dCW�1��~&��ϸ���ޏ{-墐��(�g����.^f��>y��j}�Q�����L���	�Ϊ-��Z\Gz_������<7p��B��ؗ'�������<�{�'��( j&X[�@_�<���>�~%�c��>��#ޔ�FO�2µN�بUײ$zx�6�n/���d9Q���;�,H^'�3+�G6�G��ZQ��/:1��Ԋeu�I������:�>�q+�B�󂙣�)�I�[(����6%���kg��j�w��F�7m���lw��>�E��y�K
�%>����.���6\x'�0�h�E��=F�[:�*�68]�:*���DBhg^sy#hj��T�V����8r6�o���p��8�a8﯍8�wh]5�o�%])f�̓���dp�AJ�|�C�����nљ���05�o�.rk�]�=���m�u�	wfT�r3����N�M�-�R����Ke皸o%#�ϥ����@�����&�B�k��WU��s�'��>��ǻH4}j�7�.>�鉧����w�q�~7�k�=/�A��dG�z y�_�#��Zz��^��O�P�70XUj�������_�qߜ�i���.yUx��⇼j�(�I���_l��^3�}�vY&��(�;"j���Q
�}�E.u�9φ�G�f�sܐ!�Fm��VM��Z��;�91��C�r}�_��=%��g��O�T��q]���I��\��]��C���隌�_B��mXb��;�'{ά{�"+��f���WmB��V��=�ҕ��E<�y�)J>�}ҁ��`J�~���M�Q^�]�z+Gx�<KG7|fWm߷�ɚ�*|��^�>����T+�ͪ�k�ý���
�~��Ӭ���/��"������(�Դ8ݣ���{^�f��K$`�5t��i�Ǡx�o�[���]vN3��n�K����9��>��z=�ΟБ�q~V���Zc��W�x[����U�ϛ��d^8l.��p����QeUi���힩���34��!������� �{|���&�[�bv��ґ�L���2�"���#9���E< !%QѬj4p�P�\�z�*py�]�ڊ�v����Kѐr��;��=Vץpy�c�؎`�8���夤鲑��=��{Go���F���X=���~+jPr�B�]���w��.;��<��yϙ����u_\k�Qf9lL�G��SjyQ_	��L�M�E���ܞ�ˮ�\|�y��޽�/N���î]��M�q��U�'��E�%�y�yp��VQ��{.����cU���|Ϸ\i��dd|����F�ׇv���~�D�W��/8�ɻ5���.Č�c��ޙ���tУ�R>��낍<J�׭#������D�3�^��m��vOj��g�l��T�D�AU�P���9��X\s�/��J����Y��<~�5w�u/���7:���@A�BbedG�&˞�.Ke\���}t��{�>��\3<6��T;n�H^�ٮ�=���=Ad�Ҙ�m?L�O� +�{,�ωD��_su�+���U�u�W�Sbe�}��(ί3��зY�7\�:<�5�j_�WNG����M��/��n��ݨ����0����ofﵘ�F�RsK��_7~�O�/U}�1�_Ayv<0�B�(�}�A��<cr��UBL�֒mB���L^�S�}�u}�٥�^�W�	se�r�K9����Ԙ���{�"���ͷ�t����/��/U!�)d#VUJ��8S�E�3˭ݺ��6��We��F�wu�!�%�Z��n�Y��(���շ�L]Q�u�;l�������ͺʍ�5b]�}B�	�0.k.s9
��m6�0��Yo7���E�S�/V�٭��a0w�+V��U�jo,�P1���B�k-Ν�XKD�
R��*'8�t�ef��"9��Ĩ��f�~E+z{�ҡ�k�.s
#�C"�A��N�w5�3W+�����"�şgBK�)�\�$��w�"��x;�^*���������:�]�p �r�}Ȃ8�oU��'h�x��J����0�$m��R���t����5vohI9c�f�w<�!�zs(��.���+��M�mU�;�ty���۝sy'C�H��X`��S���L�kV��N���"�^`�(��vap��ҕڶ�W�����+��;�`Ӿ]#��e�W�ԅ�ǯ΂Jd��}���vM�v�罤M,�|q��܀99�Z�{�`�)񛆟�rau77u�Rou�r��2j�x�Xo���rN��h1��U��mvM̕�"ÁCǬ6yF�8���(V�4eC����[�h����x���bOi����I�N�N�_u��L�:���x1�]Gw9�U���b��̫��p��;^�k%һ�̇�-S]�p���h�w���L��)�Z@��kD�n)Bm]�95�"�Y6.'�f,�mhc�Ww�u'�U��fq׏4��G�_Nd�R�Jt���r����:b�&�#�(f�k�Et�/�sˢ��o+2�C�vQ�"�Д�qn:�A��nɓvsYg��T#B����oWa�iѩ��=Z!��b׽,b�{@l��A���f�[x��4s)0bȜ�i������F7ձ�5q8���t��J�%h5��S�3m�T�yjRIVj��s�|�A�㛼'9OPqpS[$%�����gU�.��uw�i���g�L������w�@�K_1��J�u/���f&�u��ĳ�n�)+#�0l�tp=@�����ܪۤ˭՝��*
��� 
w[�d�[�/�������ͤ�_u-�>x%�qm��U�#X7�־\�����f��%�![ˢ�Ҥ`�`Wh�X�����Mi��ٛ��ܢQ'��t������]�8�K/+��&���$�;t3F�Se.4�^�ݹ��KV��ܵ2$ ➸���\;;(��2�����E0�����	Z�����V�������_̊1�W2ʦ��Z��ى>Niɵ�o:Y�L �Ebc���ٕr����9#چ���w<��4���W6�>�����C{��.vP�;�����c����{�Y��d���k�����H*](a�0�[\��#뫮'�vZ�j`p�����1SzG	qTo-|b��T���1T��f����Ðm(e��9���7vhQe��@!��<־9�h��XZ���V*R�DA	�IAR�ڕ4��R�˾��]s12\Ԋ,��KJ�1P��%�Ȳ�q��KuPI
��E�)�Ԕ��*��-+Qvv�x�B����D��D�2IL�Ũx^jB*N��ig�9��QuЊ�������IfgY>w..�e�f=�y"(I�Y�r^yE�Jy�eR�H%��Q�y�*����Ծֹ;[zڳ�IXENid��0�DvκZHh�Yy�YY�I�6%�jdF`Tb	�^IY�'l;l�	����t�\�O+�2�-CR"E+L-�s ��#n�L�s#K!(���y2�A<�=�HС�"�#�D���])eR1{yc�&�8-������ӭ���D��]O���/v���δ1���K=��9��g_)2�J�{x�K�ڼ�r����f��q�P�g�z7��g:���ۙly������G��2)vg�����ۓ]�������Fl���XZn'g�<l:7==�,yL�ڥ�_F;�x��YD�۵wH�����MTJ�Z$3��۝qV��t�#�Ӡ���%��һg´�9鸌�P�ޮHwYZ��]�Ϻ����l���ڇёq��x<��[���R�e����s�qC<z�S�}���t^z���;\�ć�u�{^W�{-�-��\f	H�D����C��~�늛�����f{%�ޡ�����.W]��GS�o�o�}�u�{~�z������BP��$OM[���^w]�wrr��׳7�7g�MG^T�ܕ��UC�R��=�}^ӛ�L�����n�[��>�R�����3� K�<9����7^�S.�ՉF��K��{�+�܃�,��^��Epmt"=(�=y�@��#P\�+��]
.Z&��c��>�G��#�=S>'�vᨻ�����A�zc�����}#M_��<�r�p`�}q10�D]*5�+�a��x�?�w����K]<�T��r�0�p,�ac���(u^-6�O�i����C�-�j���n��>|������z*�m��ҩ��eڹ��,����r�2���kme������S��	���������kmf��5�T�p��Vөӊor�CC���͛?K���!���v�c�Qr���z�lJ��0�R���v���f\��n�{�z�ل�3��1�z�(gޥW�}��Y��=v@��*>�|Tozg�N{ݘ�ݳ�k|i�p���մo�S)k5�?	�����@y?���^�AZH��#^@��I�ƌ���}:7l̈́;6H]n�M-�h��¾���;k�6o�t�7�u͟-�mڝ�6�rH:S���˒O�����w���6p>���ͦ8��%,z��2<r�˭Wn�7����l�J�ܱ�ު�7�ّ�s�o����G�Ή���q��}�D�߷]~������f_���#9Q>�=����L��sB������q%��;P��+�X��9S���[�^)��tϗ:�j�f��#��i�r<�_�YhP���v~�x�8<���pO�+ޤ�`O$�?U{wє}�ꇝ=G����Ϛ�Y���^%�<Woޭ���1�墐���\f5�&j���j�w��p�g7E���=d���ڠ���w߫�}�2��ˎ�4���@Pxe]ʉ~�԰$SɁ�ǡ�|�Ʀ0��^o����f׫s.�D���ZǼ)�ݠdר��2-5j����ܬ4�+�Oy�����X����_^^mw�Q(�V�p�4wBEZ��;+�^��S:q��^SɮQ��OG+��OY�nN��_?޿��h���%��*�}�`\n�gä�/�a�.�~��UFz�����ZV�T�gi�9�7�F�s�,���%��;�LO�yzN+�R<f���Z7wE��WU�=�Α�F�:�}��]�=���W�b9E��q.��-��Т[(�����6X��|_��"�t7~�*�����A�y����w��#k�W�<%�u�P��}Cޟ���j�f�::��;+7��F<Z��"��A���4-ש#��u ^}��4W��w"��4����9"s�WMnj٬�_�Oa�_M
+���Z;��C��{���~�q�<
��^�Fbѵ�s��W~�*Я���MDχ#q0|=jH�s�w�~;�C��6߅G{ʫ�|��Wx�L	7��|9#�p��;$��	;�O��&�fst�_��!�J�#��W�d3>���4'Ji/%�Оmq��?z������RIA�������CW�m�w>%wgT^�s"��v^�\��D��g�f���|.�;��LΞ�=�Ȁ�"�;�VX=8�����Y�4	Ec{�/��T�F�w���N��#N��L����uu�}A�C���9M��6Lm\�S�ݼ��'m�c!T���+�]A�ǹj�u1h�]3�S�rtsieu��)�AP�J\�� �B�L-!؋To��xU��H.�]x}7.�RN�훜�Iwd�׹��}��=�@�π���g9Ro�'r9�*���	�_w��Φݖ��g�9�P�h���Nz���<7����mV�]/�NF�����N?N��}�pt�{���WhXx��o_<��X�l�Ep�Fd�v�eF���2��\d�\�N�}9�����M{'}�.
Cۻ��۸_�#�������V�t�>6mR���������9ޫ0��C�5|z��-<����}`�Jg��#�=���w�[eJG�%��L	��0k��{y�eW<���H�	^��wl�z������oW��yϙ��W�mի���zǌ-�Qؓ�*n*�Ρ���>��.g�ع�'чYW�����#��}�ё��|{#ޯsT�
p;��rJ�<��z c~[��ݼ�P��k��oR&�
e�C낍C�uǱ�Sg5z+�-��F�z�^�t�z��s�f�������G�دM
�� n7i����F��Wp�֑��G��
��Ӵ-�F�P�Ƿ-܋�L�J����aڙ\����2S���ܧYB����줿j�Mi�6����A�v���S$@���mfyag.�����V>���ӕ���9#��B۵���,��e�`/�zS�-Gq<�FΖ�`jg5��a�sy�]�]��j3�]u䥛�l�KX��ϧ�CD�Vĕ>Bc�A9RN�[7�O����
-�F�8���P�\�M�%�W10�WH��=�!O���/ӛ~��/M,ڞ]�����}	*��==^����z}8����ĢjK�n���x�#`�'���_�8Շ=�}�鄶<k�n=�:-�U����9���]B`�$�>q�a!�h��S�}�ЭWo'��6���)�=�l�>���Ã�Y��G���=��xbHW�������Y�vP4_�gGh4<���P�6���zZ&s����/���(��W��kQ��qћ/�^-��e�S���8o�䣗3���N��a��]���Ǻf�Ζb����z��ޝ��n�K	H��}���5�Q��(x����Co��c/&����6���H���h��Y�k��N�%|���~�{X���Wq���\U��<b�	�$;>]T�Td֖*�����g�ۗw[�Vk����_;�z�t7�Ą�����n��~�Cܤ��BR7%�<�C�w�+�|<�_&)�k�FI�F�֋���s��P��tc9����s�3����5H`߽���G`�U��l����D��c����X���f21�[3 v(�ӓ��jbrʓ�Ч��c�=u4�z�h�v���g`�&�b(�v����	�õ�z��2;Md�d�P��س����}7�3.��XT�u|��p�Qv��!t���nl����8ZL��nϤ�훚�b�_����}U�D��Y����s�2�>�n0�|F��o��vN��'�B�P�F�2���3�w�✁1Mׁ��˸{V%��=�ґ��xڗb�o�<D��{�S�ҦH�Ӝ}�/�����nK* 	.c�׮�Ar�7�Kgq��=�E����5�Գ��w�W��g�cT�g~��k���%�0R>��&��t*	^+Le�mUo�pk�3�ǽ��Aߵ��e�u"�"7����d�2�؀_`��\)��~>���K�5S$ǭun��uRjWD���RG�=J�� ���/~�ߕ�����Ku5y�پW�޼��\ªח��{�=�����O�h�t��&&7'�\.=�W�΀��.�B���<�������(�#ћ%S,r�6��!t_�d�.���q�#�3Z�͕y&S�R����R'�Z>�v�B�s�����ˉ�;��nXW���d��f��d��K8���س�)
�Gm�ԇ;Sry@]��F�Q����U<o�{n��Q���^���t��?�x�~��<&��^�.#p_6"�;�_q�oXwMIoނ��w��S��xLu�,�Wx|ER�wZ�'TM��~z3��,��e�M|{ʬ���oT	�(b
e�6�v���Ȅ����.T�B�Z����FQ�?�a���O3l`�K;�\r�;��d���b�^���2�\�~�k�gZ������ n<��_{��U��1���Ih���C��~73�l=cy��{gyw�J��~�@sϵ_��u~������)Ѿ���X't���K���hd�z��Y��9~��Ó��u�nu���Y����/�>��I��*�9��o�1ޒv_y�JCѹ%�%=;|=Q�����|�ِ���wq�ׯ�s�t��䥣u����}#�i��۸��5�QY�$��&|=qT�����/%3�>�~%�h{��kC��e�8�����wK�H��8۵Q��Yeg� J5= w�������%͡��i������fj��++�6wk��>G8�9�u~��d)��[=K̳��T��}�H�f쫬���ϩv)�=6O�ì���Y
�y��B�{����J������~�dxa�� %/[��`�5��PqGS̖���2`��M�2	�>�}pU7�ٱ��M�x�]���J��y	�+<����u�T='����>G�d3_Z��{A-�F���{��U��ߎmp+�
�APy^�b���۫9��y '��r!�S�zkfsC[�*Q���6��.��K�)����'�~~>��m����v��We+�$o��9II�s����6}`p������$�ʶ�|�e;[�y����G�&�N6Ts�s������dS�r�����Ƕ-Q������9e�o��v�4�����F�+5wzĠ;�g�)��7� *����,x�t�>*�鎸�Q��i�_.u�+n.��?��E�(���u��c��6����s�:R]���4�'�����n�������oD�Q�4��wq8�^��}�y+`�*c��D�$�z�{�*����Bz�����K�|ֽoks���n�Y��}�;��6��y�n3��)���b�QjN}�Dw�uB�}碴f]\e�)v	�h�����1@�c���^�_�mV�]/�N�^ (�~��㌲���}Һa
�ʫ�)�>���G�6�_��:t�/�ge����W��f�vX�k���~�_��F�gp3ʻq_��T� {�}����y⸫�m�7$��q.l��έ<>��~^O[�U�h��'���%���	J���~/�G�{��=�(�_YD�n"\�=2�ȹ�37P��{727@���G�]>���a���Í>g�yי�e{�����罶|adF��5'ȩ��� ׽YF�J;ws��ŕ+�]߰���t���W���.ٴ,l��Ks�i�����|�>���
��V�������\&�ym+}ϸv�.툲�Y2҉����r�=��WU��Mol�95�/��9��B���܇�Z�����}ǆ��Q��&;�i��� z�8�;����ja���3���f���+�|4��A�G�F�W2'�V�1��܌�^g�A(�P"��D�^/낍C�uǱ�Sg>�D�wf������w��@��y�8]��^�>�%.�fCf��B�t���h�q��,�S���r����ī���sɄG��g���\.#+Ղ�s.J�@K�q0Xv�@g����2S�^z���`H�Z�;5��[m���%��iy�7�2�g��OEJ��O�un�A������(��b;��<6����x=��^����?L�w��@�>%_I|U��>��yN}�`y��61�s�I1��F�ޯ"�>f|6�ޫ����_������=p=tA	��}��Yצ�?�V/g��麏nN�nvJ͟q�d7~�O�o�ܳ�r��wc�k>���)����o���8�P�����_�,v����ڇs�~�Ţf�����7�~�TYF���P={�LM9��T���"j+��!<'ð��c.#Ӂ��9]7�/�I�R�������P�G_�^�� ��Z�87�t��agH��3Q����=�͡�W�0W�K49�w钶�G�SOv�����	��<Q����������1G�v�V���3�i��c�M.=�l���P�ck�Km��7���ٹ���l�{ӭ-�ٔ��{�U��]�����9�<}}1;�鿑�=��҆��/b2�B��
ҏ��3R��%��j2��gW��|�������{Y���{��o��\>�<b�	�7%��Ȫc,{��ݠ �t��k�μ�}�4=3�n'U�Ϛ�X��^�"����;��z���l{)��pק�4���(��ͯ����5��ɝ��Em�'�+xc��_����粘�Uv���^����a�)o��p0y�l�sRPJL�"�����AR�p�r_�ǳ���r7ҙJ13Pgg�c<�U���iG��c�r�=�@�Pg��MӐ&)��7��v��J7�;~Y��ˌ�_���O"sק�Nx��N�7�rQ� ;��+�B�.Z&�%�3�%�������]Zy��w��F��ݴ){�ه�U����k����YY(TA����Ң6h�~����ɹKuT����=>�x��ح
��׋�L�F���?zY��c�D�P}���>��mz�v��I������-�F����$x92����n�uD� H���	'� $�ԁ BID	O� BI��$I?�@����H�(�	'� H�b�	'�@�!$�@���$��	O؁ BI�$I?b�	'�@�!$�$��@��p	O�1AY&SY��1�c�_�RY��=�ݐ?���a���^�TT��(
�D
�H�cJU*�l�Z2J%B�UTAUT&Ɣ�$�ZЍ�6"���%*������ɭ` mEm���T0-[mHť�l�QK�e�Z@-f��Y��h�faJ��3m�H���CB�t/3�Ս6�e-Z�Sekf�֙Zՙ�(�k-�5V�ڱ5e���5i��Q�[d�&��f�Fٚf
�+oqݪ��[m���u�ִMl>   �����k�4%ښ��]� �Hv�
v�Mƀ�(�f ��������l��F��(h��c�   ۯ����p)��a���|� : (���
 {�o(�P��\
( �Y�@�� ��p� 	��z�+"�7L��eki�  1��3Uz�V�T
v��ѪfV�P[�� �q�Z�� ��( ���+]ݤ�f͌��Jk@�gx �t�z��.:鵧@v�r�)S]p�nM�;w]�t6�+wb��Y�7v��Ѻ�qV1��ձ�[
B�Z�QWc� �=﫭����͵��t�n�S�]k�R�]ƗZ]�v�j��Uڹ�9�WX�ڬÜq�@v��v��5dۜsm�[vv�ݖݦ쮵�ۜ�l��j��kmu��b�>  �q��p��40��mۺ��QeW6�v�l�[��ݶ��4���v��������T��]v�X�w[�sv�N뜖ܝݍ�Y�.�k	l�2X��Um��x �w�>�X˳��N-���Tu�[Kr�ݺK�Ԭ�]գ�����3w���;9�m�����u�VkV�h�v��mء�gh�h���M��ʭZ*�\�����_]n�VY��:wwR��F�j�U5��'e�n�������r�&����%��9�L��N���iͮ�ݫ��n��j���tƪ�,gwqm���%1�}� >�_&�[lmn�m��!�`�ڴ�:��뭹m6ַvp�꺺:�rܫ��un6��;S���*;�twZML]�sUͮ�gweS���`ʍ[f��ղZ3)� ������۵-WuZ��Ѷ�.+��Z��n�jew:�\�ڝ�l^�嫎���u�-��Nن
�wv�)���k��   � ��*RR4  21����@h     ����IF4��	�i� ��&M�!���       S�IDR���F	�#р�0� Ui114hhLML�~������Z~�������Q����Jq��Yy�
�o���#��,~(������ �
�#e?Ȁ�������?���������l?�=�� ��@�?�J����6H�# �����`}��~��0]����߅�zDDuCo��Z��6w*?����j�4Q.�����"��IC�b���Y23L���m���I�Ȩ�3���mSW+v�wJ]��ML�[�Z��df&�i^Ca��5�VʃC�I&50)��D4m�/Eދ{a��V�	��Q���ԷŠ���ş,whrU��Ǌ���(���l��A;��{��J+eek���d�p3��LP�V��ջ ?���H�f�0�3�V�LU�7��i�VU��ք�VO��Ș��y�qM��KF�ܼ�p:�㉂�� ���TX.��@�c��������JYwB��y2��Um
�O`��Qt^Egv�iז�\�����,T�k%���b�!Q��ΐ��-�ֹy+u�M=�Fʻ9q�M�� ��Q���m˭�R�����:s.R"	yZ��������� �h�y���	��v%�j]]���P�4��j�6j����$V�Wb�l̽��_-�1�%�Iw6��},���18��R���i��QU���L-KFC.��Q�Goe�
6D8�#͈����gG�5��p#�¥�AŢ�SmUԠ`��m*@�ʏmn	�A|E��6�(��iYK鎝&���8^��O�M��Y)��C���cv���<�oi����nhI|�$8�m<G~�C{F�ӌ�R���@ڑ�ig@[��ee;ۦ����P�m�Ǥ]^��t��t	�9�0b�����	ڻO�M-0Udh���M�-ָ�[$��s)P1X�/T���7cli1���y.��r\'l-���{D�^���YpB�i4��7x��ko,jN�c�+l�*�2��Zx�H��^Vdl;�@W����6Es2��K��$����k[i�`7̊V�J�.�j۵����1K�j�lP�<z�Emi��DŔ�j`
�7(l�Y�9v�
[�r=��t��3ZTĦ����,B���r����3VZ	@�kudlO�/4�O
����nC�F!�!��5i=��+�Xi�9G]CA� �A�Y��n�L̓���v�h[)�v�����ܗ�Ȼ�j<i!2$֬�NDu9i��7F��J��(St���z�������j��h-��2��iF[�,��0���Ke�����*l��
��7��D�y����>����4�--�uu�(�J�oFPd�ϲ�ܽ�Ў@V7�Tp4v�����X�9�iG @�4f��I[�͸�nB�a��T�[�1�ֱ��kU͖�E�x��
\�k�ącpQٸ��*��c�!7���?ax�-\�T��J� ��:�����
��6=��ݏP�l�eT�lz�����ɡw����:	��,'@�n��B6e:�#�]٥F���7��Sr�:U��blPR��b�	"TM��i�]�I�Q�� �ڽy@.ݲ���s^�Զ����{�2�t/%m\��[4l�M2A�9��	uPz+/,jJ�5L�2�:яdK�x��zk-%R�A舄Ht�'~y��D�⚚si��S���̱����Ң��k�F�dN\bC������t��
DMw-�����-�8caZ��R��׶���j������	�P�d
n�u����t(�%��8S#�ة�V��`ӥ���p-��y�Ӯ%�YtIq�J����L� ���dԆg��6���їh-�U�ϙ��ř6�B�%�Z"�����`���	ac�(줲�ټ6J��r����z%2��K���J����j��6֌͇-���Yі�n:���״E�Ϣ��jL��C̱k�)�ʈ�ʰL�/�f���� �n5m�틌����j��wA��*�mn���pԤ�����h�Y�kw��m��ٕxp�1�����/De������gp�����Ņ%�eAWb![���.����jZ��ݻ�٧#��L��F�%%����7�@c�Nҭ�E+��v3T�w���Q�D�u�gs&:Od7�һ+(L��� r�T�t��bM��FF��:۩NT�ܩ�6���N�)��$��$q��]qL�4��K�n��(��I�� "����jG2���X]�i�;G�H�J?,��۬���ʥCu�ڎ��E[��3�ԘS��e��91dp�3$��R]m�P���n��;3�ˁO��{��hI�pG]��W�4��1��s�'R8��baY#rcYn%�֊[���>�����ñ\�fAViF�����i|���M9�5��l�9�DZ�f���(ܤ+NJ#(djeܗnE�OwbĆ�9h���Qaպ�Ci�iM���ӆ��!;��n^�ܰb�ݨ�
�Ké흗����Ƣˇ`L�eZø6^֣k��ܦ�Hf�C	6�$6�v^������;P��
�E�A�kcCN�:��b�,�3nff&�e��3-�qi!�Ԋ�K��)���Y!�V��Ѯe�&m���j-z��?1�-��U�wR���@m��Y�FꙠ���7����I�5�w�ER��.�Z�V�NY/Ŧ\�_HE*�̠R�V�̷{�TC��S��qeH7)���\Kkhh��FzV�ٷ�ʒ���[���r��9R;��i��y������ ,�b�C~o":��vT+�M�ѽu�6��.f�xrw@ݸ�ȶ��5mB1��n͒�[����61	��3ڻ��[� %-�K�BX�k1�E�o&�J���&���49�a�Q�)m-85���b��(�К�l�W�Զ��LN.�'Rᙖ�n��=��A$�{W�X��-�F,���&��7`�1%e"+N�$�gN��[��Ggmc{�B̎��e�U�	�T��I^�wT$�4�*:���b���;0
n0�,gn�\A����H(+3]"c%�B���F"R��A��f�;:Z�h�G\�T����V�I[��+J��7
Hi�k�š�M�mDѨ��8�=-F�[���ȩ	������ިU0�F��STl��ު0���!��3N�"�5]�`L5w���X�"�+n�L�"u1�-a`�SR����*�9�5p"Z��r�^�k�[H� �'��
E<��(=*�>n򮬽ٍU�S6���W�-��2�cnIk J^�����7"W�y7�mͨM����R�Ĉ[�VV�A�w ���u�A33AKjL��AJ��
)Nj�1ӥw{x���kB��xh���-3LdH�ˈ���j�b��\��7eX�׵)��N!B"S���k��3I������I�5�9�.]64�ʖ�j؁��M�*d�u슛�"��t%[
�\-YȜ����x��P:�n� �ͫ�I��B�/3Y%�/5�L0�b��2�nZ�<V�a����d@">;y���o]���e�N^cvL��
�u7F�8��"Un+	]f����0j���oG��M�Sdͅ��6SCvIr�P����uh*m쭔0-)��sn�d��O5h��!�'2
 l`�+% ��j����J�͛,����Ͱ�Ap,�n��m^��B�͙4�����iڕx�D5�FD�6l[�8��Tv\�x����	$6�x.���A��f֓H
�7n,.�X�,�p�]����Qb�񂝇�meK�3%�K]_�9g'�ҙp�7%�@7RgJ2�6�F�fK�3k���C�S�E, AX�Z��t��gׂ&�f�c��v��J	��
+�:���sZ8�=ߏ�B�0V��F�|F��BP8��9볐���������\�q�%5��X3O�ۓR{{n�H%]��=�t*x�d�nٷ�T	������n�щs���$H�|����_�m���n�E���Ь٩�Ĭ\�yOB?��؉�Le͚��nL��U�i�CB�S�#\��b�Y9�Y�8w6�'�Ā^��v���P��i@��4���\��9�6
hV�� ���T�bB!�%�����������2'��a3Y#D�V1�*8K����M�,�X�����TNl�T1�/$�5��H�S؄T^�:n��&�7K��yQ�R�{�UE�ʛW��B��fP`O��m�י�e��2�"u�pʘ��&��Y���7�Bi֪���gc�4�$]̶#����J�5�E��Bo&J˄ǭ�jVIL틙�f�li��T*�f٫�6.35�U)_�bY��ʓ=:�X���f�V"�*$���k�=W��[H�C>H^��E!��iK�V�j�dY�An�nmbPb��A�5�ݵv���ˋCU���F�;���B�R��TY��.�̫T7���A�a55�I )d�F嵆n���)�7�o	�I�dt*
[�l����Gn̙4L�2��J��-Cl����AJR&mu7#��xF���[��E1��\������㦆�-c�W�����Ux��2#���X�wsV�2��ç����[�6�X	fg��X�d�W6��M%��uorl�4ڬ�V�e欽�ܵi*�#�e����+�X���:,��זKf��`�cl���^���5��Vڑ^M�4ԤB�Ƌ�c%Ҏ�� lA*Ki;e�WV��TĈ�,�б��Z�&���0�.�(v5�d��Vm���&<QeD(��2;�k,�mI��\�	���D��T�t���+���փm�wG" �[�(DЀ9Pk{���ՠ����F��t�,-�.@��:�V+�G,V��Z�v}P�6��:F�]�8��(+Y1f���u5XP�.ME(�� ��]���� ��}q��MP�[����V,����S�tu֝�Kd�cVV��m��w�+hh���ʘ�򏭬
��8�7X*jٖdڰ��j�	vͅZǘ�[Y���(Yh�k&A�o"7W�8v��N����އ!WO6�VHJ�t�F�ٸ���8Ax~��-����v�Ҽ�@˶��&Skj�:�*Ѱ��F+7I�.�*Њk�n�Gc5שT݉�H���Ztnl��G]�����v�o�К,,����ɺE�:�U�YBT�bv8mj�`��F�g* �fkO2f�f;EkNɎ��MB�=��m+7z�I,PwR%c��i��m����.*ǯ��N�	�9I;�{�^�a-R���x"N����ݵ�ڰDxT��ɀ��(Э�k� X�(�P��X�8*`=�؝Kqaj�8d���Ȃ��oUbsM	��f\w�������<��[�yi]f�k(Q�9��<DJvv�+B:���n�	-t������V��m��u�r����<e��܋Jh�3(�5%�ش)�AS�n�
	��]�pb;�1N�dIX�Qm�Z�����^��bԧ��)\��H��%�y��j��ɊL�����`��#2�܂���fT����2[z0N��l�*(줂.z�N��4��j��㒌�2��Ɇγ�mER)�;w�h�� ������W�b5�X��C�4ҽ�j�9�7HdAͬ��`���1a&��p�"���^n��ޛё��5�3(��h4�n�8��KeZxt=-��%/qǡ��jQ�
vY�ф�ڎH��ĨR �a�gV�s0֕���sd;4NWWC���%�`���8����i4}�+��DJɷM��2�ӻj��V��Wx%�j�B�L&�X�@�h�	�n�i]^��lР1�B�!�%T�rFen�����6�c���	��X	YV�d��#V�bYa��1�x���/7�g2e:"�[����|�ټ ��Ԑeꏝ��b�|1��??�Ϝ�8�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�RI$&�#R��˙7����<�Hv��ԓ�1wc|_b�R���`Z&��<�+:�����(�����,�=�b<4��1e�X���"_�!����{$��[��eG ���u� �]իW��k�N6˕���YP�$�2F@���M㮝��?7/��ͼх>��k{	v%[���1���b`�YX���Z��S���<�v>��}���50�]���fx�/z�}�?�!��u�^7�8|�t�RP�撔B��+6�:2	Y��V^gc��kh�����;	���ΐ���yP�-wE�31��(�"%)�NG�W���w%��]lv#�)��Z75��rt7�]1��{Ie�ں��\=aޤ�q��; �#��:U��[��w3Wg3��_+WwQ�V���&�]+��ڊ�r�;�a�C�(Ǵ�D��ŷI�����6k�N���K�Y[�]<������fj��[�.��<��Ί�㇭J<T�]/eY�j�k��HV��@"r����lZ4x�h�1��Q󵼻GhT�k�Ql^mDb��֨T�3{vc*w�������Љ�q��T�j�b�;�v.wj���k�U��.ٸd4���/Y=�ob��.J2�Y�9"� x���S<sE�;e�^�3]���r����U8����k]�\�>�0vR��reD��#���7E�X���}²W�4���=��Z�~N��O����쭥XE�ᢛ3�H*K���ZZ�{�l7��%���;fR4�'�L�l�х�+�e=���\X�/6�B��Y=��P7n��6��x��7+�Ƅ�^�ݨ�?�2ؠ�<u=yY�*ا���']�0I�UAr��e�D\�	'��n)���������	-�!"���89�ObU�P�1t��;���To�		j\gmP��{7ce���%Al���qh�[@GO2��Vp���hݨ��Ơuw%8�_,�'\�����c�x��y�B���]�k>��eZ)S;mp[� �{S�S_^�)��h��+C"�6�v�(�2�xV�j�h�[O%K�jt��G����U���$���1:���n0�ؤ_��^[x+u����ꋳK5�V
��6��S�ט��W:������]����Wm����P��Leuv�n�Z�+���\�8�n�Y�6�4t����%6�]K��xI|7u�`+ci}v���-S�g�Ȟ�ǖԐTtV6��:�#V��SEn<��W�K[n;��݈n��}u�g<H:B��\+o&y�-����&ܬ�V�n����V���ose:=���8��Q��g,�4X�Nt�9v�J��1�L��lX�Pg.v>M ЙXN��]��S�*֎��͹"�Éѽ�����k-�Z�E�WG�6TZ�%ŴЈ�Xk� ���Z:�U�uz��
�rӜ��H�iNX8��	�r7R���8*+��rT�����卩,֋Ohw�Ή�}�B�:�'n1R/�n��+s�BaW��,���]���e�'��[�tV�"0��v�am;.j1�-�5J! 6�=�dE�u�ა�Œ. ���.�F/�3Dx �{d��)������N�(�v@��y�j�uԒRF�ᬃ�$�h[v(�rw2C����$<�{[%��_[J�i'\�X�U����4�FU\��uf5�����$�zy�K�4�F�{*W<vY����AtuV
oL�_כ�@����]��dn�"D�\Hluj��E�A/x�;��t����z`΀A�.�.���pM���g:g�pK�ـ��q�7JM�<��B�,�B;��<;��G�Ћ8]9wȕ�xĲ�ه�ot�t8.���yq�֔�z��m.��,v�ᖪ1]�mb
ĹNvu�*�N���t��:"s��%\���.�*���ۋo�osɨJǃ9�g.
��a��P阱�y\�ś�-���r�8Ɓ���-o&�Lw��.oL�!�b��z��F!e��C�X�O�Ro)u��0��|咆�VU�F*���.�s/�|�Ϯ�H�ke[�On���.����i�Kivrj޸D��GԶ�f}mw��.�i�ѩVY���b�픙��H���gn��x�&�t�1�\k%�+��L�Z�0$�]�G��+�f��pz��b:�(:R�Y݊�u�o+�b��J���uR�q,�y.�.ݝ�ێ��"��������J�Y�"�]��E(��(�n��:I�l��f���t��^>m��K�qB.� �G{Ce�TWG5�T�둬�V�Xɘ*��w���f|����h�=�Xy72�����*�+�F-H��V[����:v&�*����ȧ��j&�]�<(�D�2�	��d��N=b�]���Ƴ�$��ͥ���n�QՆ�R��׏�W�*�gu��u͋;���w�.RR��wH<��Yy�Gu�:͡+�7���ѣnGiV�*\ks-�"�����%F���'���Zw�֚����MY:lR�)V��F��Zx vo[�8d��B�-Y�z��.hX͘uҠ$.��dK�ᚧd�H�6�,͎>7��SH�շ�����R&�>��*���K����o���s�{�p�rc�|�n��W�l@u����Y�\ �F�il�sX�S��J�u��\mc�<�k��5�C�G��,4������N
K6]�ލ����ky��NCs~\�vw3�\�7[��P�����
��V��Auq����$�����Uj�J������E���~8hxoقu�4����w���Y�uÜ��.x�A�%6����Ae5�pxN'��c��X�u��d�xmW\���m�U�q5�t�v���:�Jc�+�s��Y�ٝVn.��;��i�ҫ���&ņ�zN�����j��Y/c"�V���c#{(�낉c�*L�֊���XCV-�9b.m�w!F���F ��\���Mћ����k����؝Mn
ݔw�cW�_L\sz�-U�Q,i��i�#�ɚ�������ɒu�����GFRY&��F�Ȭж�X|J���^=&D�Ⓧ<ʷ\X����vVuF	l+j�AY�so��'�%^M�=��X��M
>��P�2I,��ePuj�$�m���2W;�����{&��ę�K�fV�⫰�|gB�8Ŵk�]gS@��@��3ثm6�-�w�q�i�M�X�z�mgn�%�.�����Ǒl���p��X{_c�`X�����j%�ѷ����U�	����6FEH-�[��X�xdג�oB��5�w۴wEȖ�-ޱ;�%j��X3n�[�{�P�ە��sqLuo��	m�o��9ή�U�Υ������Q;�@��jV�Uf����+$$�����ݢ����{`Xu z��������&!�����[}�
���D-g;Q�)Kp.��\�=�z*j��H��g�����\`�WZɱx�8�!�W\�*ؒ�.�8���Px��h�w�m��m����n]>d��K	&�H؂w�f�϶��&���aV�m�F�		�'�ԛ�V�zq�%df#G:}�,�@L�Ad����z����v��.oC(�� n�՛t����t�EqZ0@��̵�o� �R>�{�ubZ�wP��'��t�rh|����Z7�]B��l���躕p�Nj�`�`ջ�wh\���"�i��r���u���LI��To����EH��p	�d�pn��K��)����R��X8e� �{�h�5�r�[7���-�:`�Ë�:��Ϲ�����ZѶi�m�NhU96�0� O����wif�[��5��e�v�`F��[\�Z�z����!a�� Yw��;�t����X������&#�nVs :��=��  ��
�J\�돇v-�S wgU�ֹ�p�v���Ν\mU�XF.{��ڷ���L���6^�iA��r�y.�WJYt�B������b��{3�;��ao�V���E.w�b^��ݙ�~s1Ҹ�t֒��a�u��"��'N�{���	�w	���p'J�M*���=�nq}ʐ�b�v�f�b�ÜJi�b�t�/ R.��s}��Y�>b��u��Gl�͐�*�h���^<�PQ�\����D]fTG{6�l��C�w:ǫ�u���ÝJ��l؅�tt������bFNH�P�64$�C���»F��8�<bеѹb�Ҹb{��9��,7�����awW�}�iLo7�%��ݘ��h������@u4g��v���{�s�rm+{Sw:�7�D�n�^���8�W��*5l*tR��o��\5e��E��Xṵ�F�u��� ��h�YXV��EG��j 9{��[̗'�liI�Yxe v��1��(�J�S�W�A��Rz��m����	��ɦ��PdX�������}z�9j|6��?�Q\���.^-xq�hV�ӮJ�J��kccٖ��[]��$���2���� �zq�{ʑ�Ք�h���l��-)I�"���r�N�����:�+ԩ�B�S����7��Pv�+v�T��z�yo'�k`��@� !�����U��m4j�C���u�ˀU�ev����-��K鳹\��L�*��r�fS���[3T�,��8[�U���в��z��[q�{/]0iw���2��=4�sx>�ab�-��R������uӽ�V���bg�Z�l�I��A%&g\�#��\1M�vX���{�$,���t�X�ڮR���0Ӯ��=�-�����rJ�l%[����	�cL壵�)8J(���z�ߦ��Q��ڛ�<�Rڨ��a��N��{'%���mV����gx�X��A��w��ou�Z��p�R"���i�e�nY�N1nw­�Ζh��\K��+gK��'wg���ȫ�pW=���iz�u���	P�������=�Ԧa��MjwՂ�.�ƪ����I�VT�WP���+1)�m��8���Ǔab�Et����G����βeն:

b��nR:p=؆-6ra��})%"Q�[ج��Q������W�V�k��;�9�7��n����}�G�>���j�1��g��B*�o��+�e� dB��IwL�'��^e�v�&���e��}z��<pŔ��3��}2���2�dRe^8����{*�i˖+�7ND��+pn���J:��񈻅�n��kΕ�4\��5#���j�E�OK��HU���0Vs�E&w�\���(Ï���w2 �[���Z��BN' u�S��G&E6�"�9j�&���r���G&�'*99�W�$�_Sշ�dQn���J��/#�v�ȩL����u�]K��;��`V]��2Wv��dvz9�͛�G�G�i�K�̬��`͚��{l������FIJfQ�VWL4�1$�nN��Ժ��҅�'9��%+{`H�i����QZ�����w�H���)ή�b�j����XUvM9�
}ч[�wTػB��=��fPp��iWL���'��6.V���n�]�H�{��a�Çu�#�$�����;yH�\�I���2	ҎG���ك\����Q�}��F5�Vԡ}��2�F�Jj4��9�V�RI�$��ty�.s���Z͎Ar;����y�C+�;N�3S�8�j�I"I$�I$�I$�I%Ux�)�B��sI`���"nQ���(+f�G't�A+�����n'=�ej���ͮ����i��5ٝ�Z�z�z m���V��bw/r��Ŏ��'Ջ�"w{RI$�I$�I/��������ã�?�|�"��$7{o� ���"ؚ?#vD~����|�^�//���>W�*R=����n��7�G��s�RnD���]���j�{��`���1c��Z雷��V#�k�S�h����';J�ڀ,3�J-Y.�Մ��h��:͛�+"��i)��q=��� *����ϔݨ��Q\D�\��R�Vd�aZ���b|6�̡ϥ�;wt�pm<Uf�:n��A��Lc�A5���m���ɫ%�(!�-�{�:MLVT�=�0����ï�J�uз ���Xd�S`�*�T˫�J�C�*�p�c��Ҹ2;'��	��+q��wt'	|X+��C�>��-C��I�wa���5�)� �Oz���z�i�8���n�ið��R��w&Ou4\�cy��qnh��}�@��OfV�$��q�{Z��W4{!��oj��׊-�r���Y����{��K
̽��R��P������k��K�\���	f�; � ��6�!E�]+���N�bo	o�mr��a��[�H�gŬzi�Q�1	
N����]��2� �mc��h��.�U@�찔�|�XQ=w����q:X�m�]���E:�yGi��x�Nck����a,������v����+�J\H�9N��]�S����]��ݢ��nJZ�fR)jrgfЉ�M���:�]\��*�G|�tqԬBy�1" �$�����bv"*�-���2�͑CZᏍ�c���B}i� ��u�U�u{׶�᷷Ygz�z����p�8����ۢ�&�3��ås%��]\�]_�n�Z�f��o:ҭHS� o[9Σ\7�	�KS�<*����\K�n�IԵ�PwC�<�&�4JcbD���29P�&�+�Kk�ɺ��pö�P�;�|Ӈ�B�p�Gy���ް�o5^QQ�(a�J+����)��q�ڬ�7���k :v�Vq�]Ù�K�˯�۝��u���.�X2��U-ܥ�B$�u���wǨf������N����hb(hr�^�WVє�o�\�m`pǖ��-��\W)����j���6�Z�.�DAY��Yۨ�F��}��Go,��S3*@NKVuަ��U {���OD炵s�ԫ��jm�5(��k,��A�.3OJH�R�eWJi!u}t�V[N�r��R��V��Yt�
��+�ّ�[٥��A��%�l�__2�i�\m6�^·�ףNP��\ڐ���|�K�rf�ҧ9m��7r��k!��Wq��]��o<��9��˻�]o<��u�]�Z�b"�fYD���['IQfQ\���"��=�/�&��9��Ws:�)YSsg5��U�kKL��I��9b[�]d�)h+Rʥ�
�p�Hf�28A�;��!k#�����ޙH옥��*elf�e��xSjH6�Ze��=FU�.�I]��bѷ3t��#g�̽q>�摛p�Dqk�1�-���e�t�� ����Q����ab��=9C���R�����l�#:�>�Gk`4�-�'�*Vt@�s���;7��Y����Q��\K(a?p9�$Y܀��)2W �Q��D�3%�^;��W�֒+���J׻V��`˃D�,�L�����k+)��eE��.U�#��Ӡ�Y�,*�*ﲷ{@��.��m�f�<��vJ�
q3�M)�*�*���m�`�-���u��Mn�ȧ�{r���h��t���#p�q�V%�CT�����N���B�u]kX���
F��q���[�j��i\N������EY��(^c�八� &��jJ��%�tVo
�ˤ�l99��N�E�ig]MwԎ�9�/�lO��Gc�uq\�H�K�
:U�J�
�k$�ɝ�1l��Ɉ��S�O-�u�*�:,<�QwfV��LӾ
�SZ�jf�����G�aA\��L��e�R*m$5L8 �ge!�q��)Ӣ�f�Z�B�p�WX�L�O.�G\�wz/�-l�a²��O�i�x7��S��7Ѭ�6��S�(P��3�<o(T'l��W:"��B(��ER�e��s���v�i �E�+#F�)
��V>���wm���\C��+a��#͗O����˝krR����,q�n�g�0��s]��"�Ҩ��9�֦rT��M���l�e5��au��q�hn�}���kb]Ϟ�\Se���m�i�u,�l�V2�̰,R�7�#��
:�\��7�[L���+{Div�Nܣ.tW|^a!`���z捦�Q�jZ�h��Tx�`�z�^ne��W�2^���2d�����Ys�٠���������WL�LMc�N��]⛕���\��s ��]k�)�:����1�d
�0��)�����l8� �8I�uw<D�*Ȣ�������5����R��qڼlu���<\�mP9]
�7Pڭ%3:em�,Y.[Q8�U�(*��v��9�6�Fӡ��C��{tSsr�P���2���;6�5��)6�(U;��kv�!H�G6mu1X���N��ۍUZ��RqW�u�RS/���B��`(.�Q2��:*`&�����/�w��K�7&NM�ɢ�qwz�^��vз`c]��c����H滣.,�o�ި�ٮ��z'���Z�D���P��E+5�moN��/J�-ön�ù2+���*Pvk�������;���ŎoqWYǝ��� BۉWHl���XU.��NMŵ(	AQ��тh��ʃ����k�Ю�1EI^O�(��]K�ܰѼ.0��ⲙq0n����K��/�F�䬾cjW:c�\+)E��k�Pl��e�<�3~5���b�u�ȟL vq��'t*���rCYAfa��G"��֡�Ǣ���D�\����9|ힾ���/CΗ�n)�3sje V��ܥ�f3�����N��ίs+~[Y�':ꇑz�2�"�Z����9^��F]Y��r�G)�B�i�e�j,3�c��'^U��ы���e�P#\�,t#q�. �)e�֖تȸ��2M����md�˛���#��Y�R
KyP��7,Ps�j�V�ۮ�����װ��oV��ChжY']}ꋩ!����M��f�<&�d��h��5��e
��v���{n���C*+q�w���p}�+�V��#�0��,�򍌽{N�`p���寝w;͡Q�>i�	�h�_^�C�%�D�Z~�[6�ۈ�ʢ�7kʍ�ɵ�D��gv�i)�F�!����9m^��˾�E5î�>��3NBd�s@����{�.�ʂ����y��R�1�uE�N�j��7q����Ѧ��&i�:�#V>��u���.t��،�E�e�RV8���>�5�dN��r4�_
��԰N���	���]i!Qd��6VU�'�a
�WS���)d ��_]ޜΕ.�V��ߏЪ�'O�[O{�4�̏j�#�㉃���}�Z��Zo��,T�����&�c�;y�[}1�1ޔc��i�Нn��n$�M����ր�W6qs��z�*!]ۑWSE����Zt+5��7�����L܊�Y�r�rw4
����;N4��rQ�4��;7�-��S��*s
�m3 l��N���X���������s��w��!�&�����v#9��M���AZ��� � �h;�C[m�g3����t��\~/c˝�&����%e5e]�l;�����tE�*3n��Gr�uY	_iۋ�I�E��>�u���l��7"�)j�hV��>|�,�M���d?s���)����R�2��j�}V�y��l�<�%Lj��G�#��i���T�b�3�Ѻ\b���s��vi
\*�H�<�l�L�@L��]����Q"�Af�mX+4�FTs.O@�� ��n���a���̼{EU�=�VL��	R�@a0�	�8�l�A��;�K��*�c#��v1u�q>aE�S���oe��7�&U�.�K~�΄rMZ��9��پ\x�'>�͙Mr�����ڔD�.�)&��3�n��YN��u+طl]p��A�Yn��@\`�����J�N��f-	Y�G[�N��2�s�)�l��@IwL������w*ֺ���kOm��VZ�䕻O�7���C���y[j����0b�r�_]�����i��
�4�}Sf]d:�VPG{9��'��-�b�R9t�z�8�k���+�Jj��ky�	v��5*+�8+na��0*Y]8��l�5����v
8��
"��b�y�^��]D���e��#�y���dܱ���t����m�K&:�F:c�sL�r)O.�s!�f������N*�����ee%a�m��qt�q��ݴ�����X��[v���tmoS�w�E�w�f�X;)r�j�M2m�+P�誳29���w*�jհw5Q<����7�2��:����Ti΋�n��vB��\���7Aފ����f���Z��.ˊS������t��kG;�R��:�uf�յq|�����Ut�o&����)W&R��W.r��>�r���wL�3+,Dͷu,ч*�z�b�B�Z�L:�����yF��f�Ir�����r�1C�]m<�])w絁����~L˫�wΗ ;� ��-NYz�]�O�)1g4��}��u���z�E��6=����ܜ�9�|�R����Q�r���'ED�@�^�e����d�@m����;�H�w]
��L�#udjgU�Ǭ�r9�ܕL��q�۔бcLUהȺ��W�
G���8��-ɶ�+��V��NV���c�@$牅�>�{�
�R��u���ZM];T�IhAȳ-�oKݾ�q�Ѳ6�I#vibf,f�����.��@�V�P��=�k�{�g�Yd[}f���(Ex��4�8:�1Y�6BWy����vu�,z��	�r�Ȅg����:6r���Nˏ�=5"뤏U��Ѷ�:&��NW$�1��Uy�졒��T�S��Yw���\� W����3�S]jX�ʹ�z��9�.�T�\�R{r�M�\]���i�!�(a��2�Z�iV4��N�՘3SdnRl�/�D6�9R�ٷ�YS��t����0Z��� �_)r���-]�f���%.�e����5�B{k�
*VL{;�r� ̣zoec�^��YʸBr� ,+=�ms��!4+`R����]����[p�$p�Yc���+�6v�ݐ:mw�D�n�2�(~\�����2���^�r7x�c��C�P�f��m���p2�]wfn2S͢%\��M͕ej��L�X��[��;����]��E�-S�{���Q�V~�[+
�qY����ؽ�H�o�,��"�k�ʕ�H��wu��MsL�inL�f�����������p�sWI��)'ۭ�Y;{>V��.asU�p��*�X,�<}\�E�k�о�v^�S.���fEud��)��J@ws�].隲V��y��>x��1އYJ�� }�<Bۖ!$N��4a�k�J��[�sWPr2�`ͣ�WDj��sbWlK�����j/��o�l|.cJ��à����1(@����9���I�>���@��ؒ.�L��R�0�EV��=tT���[�-h�e�<2�Z� �r�\��6�^A�.ƣA�j�ۅK��f��7)��C��eQ��۰/mt�	�����,�
�Y["�B%|�d�n�W,��\󈹐��Y�4�Y���YS/>yq>*�X�����ܢ�ɶ*B�%-Z�[7ή��;��t�q}]d����R�p9Af$m�3�I)�\�{V�,��v�>�U�&�O���3��Y"�Q�R���of-�K��u���U��rj��3S�? D@F$I?����&�@9hG��;���ƒI$�I$�IV�h��]��u�rN�nv,�w�v�3:]MA����P�B��.k�*9s8�!{]F��'*�N�_n�ѷkNQ�\e��O�/�x��p��G3��Q5�����*[b��WD��WK�x��'R5�[+IiQk��<���t��f�lG*e֚EЙ�3tI�&=P7��Qy��ʄ�k�|�G}�e��6���9f�a>��՘��BU�ұ�v�R��ڭ��YsI��O�Gd�.��ī��f�־&�)�d,��Jx��G+���be���]��Sލ<w���.�;fŸyq�G�lvC��%��o��*����.5��vؗ<c�;ϰ� r�Fu��.X/pا�VҔ2��:�d�]9lpK���l�sbE����ft�˨���5��3~�`�J]gSV�2�м4���'��(���֥5J=���J�5���;���[���+�����"ᄧ�AI%��Lq��Z����ߟkV�,���X�]^*��ۊ���n%��̜.�C�����*�k����]Os���Ԕ����5ɽ��q�F��빼�B]��72)E���kf�щ�}�
���ܸ^8u���Q��No���nc��k�Gq6���3�}�UcA}�fɪ �������	a������yI>N��e{���j^�=��%�S9��M���Ϟ'�}e1m�:6�(+Ĉ��$���x���rgZ2�[�m�vY���No�x5��ǟ�H�
���dɒ=y�I�#28�Ȣ':���M�
�69�wJ���'��e�>���Ȯ#&ID���!���zG[0����^��x��s�t���w�Iu]$�����>�J,��U���$U��0�I�X��UG��6����1l���5��4;�?W�g�>گ$E��f����=��^ei���גD�M*0���۾~aiU�̼�Z1�K��k5ٶ��yܚ�j
۱����K�vŹ{̸��_�F��)Q��g�h�縒jQe�c�Z��O��a\�U���"�5U�
+2��3��w�?ԯ������o)L��5,F�Q�wQw�Pˮ
�M�6�'�<��C�f	��<j�hݎΐ����ܯ�sV�p�?��ܪ��{��Ʀl^�X��$ꑽY�lֻ���yU9y�����}�f�*�I��`�)���l���R���x�ٜ��z"�l�;x{{��4�o���	B�O��oJ�I�;\���������#[w��&�$���Qg�u�ĔV�E腂q�"�G=^�
|؏o0��v���ป����I�ha	1�^#��E\���.�x
_v_]T��1[8�9*��Y՗�<���bViq�2`��{�"&���:S��v�t�.y��u��SI=-UC�ޞSي����!�##��#�IV�S�M�u���U[��E4�`ali�Ǧ\����¥S:���>�T!5m
��U<���[�L|=�$��RO������!$��)�y����$�!L#��9�@w��lBc;�9̓o����qªi��w|#�
�D=z��>�G[��o�
P�t�P�[ԥNX����=�m4�A�l7�C��9�?����՞��xla��{�PC�/D�Xϒn���vtOWep��#%Ѝt���PČ��.�Cor�U��{�ܺ~p�q�K�
Ge
5��1JQ;����'���7oOI�zC�ȿ�lN'�������h%F�>5n5�i���m,ab�sX�&��*��Ż$F0��I]D	����g.�|���)I�ҔV�K(t�O��L���>g^l���˾�9ܭk6=�)�F{�ЉPة��*3�H�����{��V���߽���©�� �^�˱��ǔ噠VVDI���OE+zt���r��\#��t�F+t\Lȇ]��5r�
�Ë-�\�o��<�	�欙3(C�8�E���0���kA	W]$��ǘ�VTA��i
c�LLFs+.V��rۉ��Ti�����f���N�x/%i��JI;���6���ӂXkMN���/�{[�u��(��8��P��T��|�7�J51w.�Z��B�5��V��}o���j����y16�W`��=�{��d#S'Gq�i:������M������Tde�J���r��rP��Ť��|�h;dB'{�۴��Cԣ�⻟9N[�����Y����(Z{�U���\���뎹�4�txveP�B����A{=*+��N�)�{jg��R��x���gW�%�����J�ޞZX.%�Y
����qJ����S-_�f}\61*�7����ۧK,35L=7�O�xtS�1<��qN��6��V��""��C���Ȕꎬ���Ci�ۉM�N�S�S����������_���ubc�F��Vjլ�|fzr���6��f��M:�E�ͤ�w����3ͳ~<���v�&tгɍ)Ǟ�7z�h��r�W]�^�W��-(�.Y����ńf�
�)Vt��s�s<(%L�ە�6�c]{"�P'�5(��sFc[*�R��"RGo�.jJ[2��G*9t�P<�юq\��.}�몸�^�q��8j��u����cl[�^��O�*ɱJH��^W�G>�h5��:D-�W�=�c�Wp���U	���ͷ84Jy���t�E��e�ݷ>�7n��x�޷9�N����
g�ឞr�<�	�B#:�S�X�y}���r6h�c8����r��9	���	�4n����\���N����xt�N�j�4[�sR�x���1b�.���N�mS�e�\H�&=�T�m�P��ut�ʄ3-�]�U�;��rIį~���My+̗�}�u���#me\�0Q���6�k�S�S���7�O�M����>���F]
��ų�c�z�$�kג�-Ky�^�hו�z�_V,g�jBnҥ3���zt�&4��\T�h����R�V�԰�n�{���o^+�v:�}�z�a��ۺ.[Z��0�H��H���pVM��;E�f�􀽻}�w�\��Y5���j�Q���tu�WpTy��ԓ���ނ\�n'��e���l�#���ʢ��{�'_g@�^nb�+�����,P��b9��d_;vq��F�3]�i�Gz���CTנhX�Ʃ�=Q+�=5�뷉X���.��Ϲ�����]��Y�~��03���)���u�1vƌ��Ʌoe��Ѽ̈́���[ʧ<��V@����lq;�x0kܬКɃ6�lH���}�f�6��_�ÇUX�b.����=GP�����*�����w,���M$i��8C�\���]��b�G3�_�P铺۠\ؘ̈W�Ԟ5Ou�t��]	\<���gL����Bر
[tff�No���aMg_'�nwHѝCt��2q�qW��F�ʐ鶫&���}	��~6�ن_3�C�����[�@ޝ׽,j6�=@S���\3���Y�-Z�L�=ڣ�wH�i�dB,�]����۽#�@�R�X��]�Sf�	�7s֩�Yu��&%�����E�worSX��4��^�d)��r܋��^+Ej+8R�X�����O�7�
�̈́��j�)��+�Ӟ�K�N�`z�̸�Z���w	�G�_W[�S9�^�֭�䝧ˍ;���&k\�1Qm��\��]�l���&ᬬ��W�0� �s�94�঄�f�q����W�Z��d잒SSVbZ�S'7�:�g��S�Hl�g�#9u*ڛX�Bn��)!V3l�%�3�+o�+�2�ʁ�":xR����s�F�r�9�̯g^�r��r�H���2�RF{m
8�B�_NZR�&{�r�糦������ͦX����[�����62�9�*u"�d��T=
��NE���b�����T�$�y�{�N���θ�kLI�5`� �T��]g=�N�0Lܔ���{��� 8v�j����A^l���S��lWoI�)�X���v6��#:V\�T�W:��͉S���b�S����rAa"sTXK�B|p�L__-E�`ҳ�%$m;+vK6�ە���z�;�Ò��SU�3鋑{�{"�xb�RK_+W��3��C�!�#�t-�.��T�v���ن�\�Pf���^�8)'�(JfP�<1Lis(��j�3q�]�I��s�+�y\
�<�RO	L��O,�_v�t��YwI)�w��XQc���y��v50��;-��s0YZˌ�f����1��%1�d)z彸B�;t�xZ5S����_;�9I��X��|_��P��v�[�d!"�[jGk��f�R�y�ݝή~޼���s�@�U�Sy(g�� Zfi���r]�]�ޛ�0�^u�w��g�ڡ��nҹɚ{"��h�w���jk������^<�7YK9��Qg�p���a�[[��a8��� B�"���*����h{�c'D.��k�usLRԅ$�:s����/p��N�VU�'�Z^���S�h��Jh���kC+k��X/�/7mR�D>Md�w]*���o �}�8r6�ꡰ�Zd5n�oT��!��0�W#���T�*7��"���<�F��=������W�E����}~������e:'9�<Ұ�f�|՝U=����0A�� c�t���]�u�MN4���1V��-U��Q����C(\h�<�������7Y����i���	��OBS�*�5�yp�y�Bڐ����Ǫ��y1N��[ʯ	�>�j�u�ħ�����g�<�����fuoq�혹F�z_K�o�5�)�N��387�!sC��mN�A�	�Blצ��+�L��a�.b�d��9�$��.�	t��EV�*���oJ>��(���X5v^���`hi�޷
�B�Kf���8�a�QB�n�O~C����>�ښ�+n�j�3@Hq�[w��~��:s�9,�J�L��DU�.90�\- �5�A�Ş��C�m��	i��r�7�rRG���rJI������!��<V�TU�wsM��\�V�R�zPuu�Nv�)Y���ŃX�U<���S�W]��r��x���w	�
n��)��C-���U���[Q^o����W�[�j���>�;��xect3�41c��(=w�������{�t�� ���*�D1<�L@�"���洹oM���S鞭�œ����:>ѷ FO�)��g{���=���bO_-�wX�<ԛ���k5�vu3���GG��(+�m[�W;�ϩI[���cS�j,�da��b5�~�Q��qN	)�d�=�|�i��{�����^zd�
��n��3҅���;����ʺ"�9n��|���=j���5�!,��}�f�*�I����tI��r>��қ<�VW9b� ͗o&E��X���ۗ�HP�9�+��<�#ta�
�Kn�A�����i*�eޡ��Qʆ����RI��Ź��5�+J��Kn!x2�eͥ�]M��vru�Q�"�犹Hf]2��>p*ԋ�7�t��J�ħ�kt�AYLJg^v�U:�0GH����.d�G�Qm᝖�BD�P���t��rCs�x0��(O#(B�8�F�26o������V�Qu��^���k" TՈ|�HH��A�	�@E^�wZ^����Nr��[B�SvZ5=���"���k��_�����9�,��;lO��y�*f��)�B�tl�%��#��J`C���<�f�
�o��j���6�ݹ�{3A��y±��3�(�����	ɟRtP�����lS���N�w�ob�{�$�N��f��q���٦��Lȼ\cb�usS��y��u*;��d�|₫��6r�F��6�=��?hD{��~[��C謄�횱K��-.�,
���T�+}ǫD�Mz�C���G\�\ڡ�i!\� ��y[:��]��Cև r�/0*c)���6��2����^x!v�Z����S͸���XFY5%s��F��/>�f�W�D�s�e��.�hP]�5%���X8��y6�ri!e:���F��݌�3�Jį_E/���ܹA��>4���4�CMI��/J�:N5,m�j���M%4��L4RL�m�TF�\*AO=�΀��g�K6��2L)ή��ub^����������$�f��pX9e��/h��T�y�fr/���.��rq��k.��O$�6�D�0:�!RZ"冞��v.C��p��Ժ���YÇ;�#���wn�"�N(�\���b�Znl]��4�kkWY^Ӄ�)R���MX�����4e�7//j�-Mo�X�c_\8�%���&�ٛ�Y�$v��n��M3՛��A*	^����j�WMk���M�m��Vc�{h�,3����Vh�ܱK�iAu�gucI,���f�&K�+�VE�	ե�>�)YW:�_]2N�[x�^N��	�Cu=�ʼ�:�����7vi��G0�a�%_㙎��a����K���[ ]�(�A�]��A��z�ɖ��sM_N���Z�M��I$�I$�Im�l}؜ݽ6��&���,�ъ�Y"*��}un�9ۺ�K��jTװ%�c�r]n�.��J�ņ�2���l	��,Y!N�u��E��3��,Y�R�;�摰��%O6Sec%����ml5.�D��jS�}�n����Nd����vWimj���Rk
�9�Ɲo9�s����#/����b�;dYb�T�tCi]ؕr)�lH�
 ^�_�!t�C��.�5bj�m����zn�)Q�>y�^�ƈh��,G�^�ƕ c��zKv�h���Y`����n�L�Lt'�c3qڔAk'
#�����K�́HQ&��Ď!��uW�i�o��Y�ͬn��ǆ��~��;z�w~Kr�A ��V1R���.�:���W���|hc%�~�]E���35���`]��nuQ<�3�!�@`"��$C�G��pIZt�i�y*�;��v��̬=��Ɓ�%���%be�9&❚mctfh��������`��;R�(͈<v���]��,W�kt�ՙ�n˼��N��9Icn�칈���0�I�	�&�}��G"�9���{�9�$�����܍�q�W~���d�߯m��f5���UC34���������;ƞ䇚T��a�D��Χ������dڞ�rm�M�գ)�Wla��0��~���D�~���\�ѱg�T�q�Db�T��Vns	�=�zqe�d�;[��I0���
O̧��]Z�A�{��{VoAj�i-l������$�Qf������}�of����k3�;4h���-d´4�.Jx����EO���<y˽�v7NdV)z۴��_�~&W�
��鳫I��ǅ<����ߗ޻�a6^<�|�5�茘�"��dM)�"o�=?A��Xp������n�z٣7*g!]��i�j�[
��� ��6ٶ<�޴����y�ȿ��<�|_gZ}�Lә5�C�nȺ�7I�q$R�^�ɭx��ѿ[��絜��+�ǽ!����<ʞ�>ǌ�u�a=K�����7̻l�*}%:�Z5k��!ì�۽���x���0���﮳z6�x?�ރ�,5�M�6����>��bzƗ��q�}�"��q���[�;�|�҂� �\�,d-ƹ�q�y!F�K;u`Tr�4�dy�;��aF�U�������mv<�!�Q+r���OR���X7�2�k\nG���K�f}����*��ɥ�~�\��#�������g�&�C�6�L>}�v���3�}��m[�gu}a�r�V��u�~t|����9�=_\��m�'X=��nP�G)���ʽ���5�w���O�YN�͞�~�%QV�Um��o�� ̀~W�+y���7�&�@�76�	�H�/�=�3؟*=��q�/���yq���ޚ��{$G-wdL����ׯ{Z�5I.��H��F\8Ў�:�+h;+�=%n�E��&'+-!Yu�$^}��[���d��ў(�]8����x�G;���3At��ϣ�U�S�MY2�2�p�\��P3b��C#/��s_L}��/�c������S�^|n�X������RW��_d晻��'�U�?=�CG��'f|_�.7FV݃��r{�-ǥ��S�.Ra����os��W��.�[���{H�CVmL"��޵*�#�;L���/od�$;�v��fmGH���״�R;LJH�GL}sa�GxV��~\L�jٖ�^��l!6��~���2���G]��/k~���S^znF�w3�����	��AU�:�m�v�*�'n���U�vzw�_V_��m���,^{��b~��̅²w�*����$ c'���g��<Y��^�J��"�.Z�B���wW��*߫'�/�����3���rQo^_��!j��t��N>a�W��L/���i�{s嘕>jf��<��O�XW&��ϱw�CQ+��
~�=�����޲�O-���WR��m�]��P���<����y
�q����Ȩ�p�Z�'�+���;�Ć��~,9q�G�5"�N؈]����]|< ��1�F��w[�bU�b��?$eyG1�S�*2���'��c�1��bհ(7VC1�ǖ�=<��s�3����Vܗ��.Ĩb��bzʵ��c��	V:�,Ұ��rvk��&��&�͛PNũ����${r�8�F�b�^^m����ڣr���b������ ����̈��j}Roi����K�����t��4�w��&'�ƥJ�e���OG��X��[Þ�j�v+�<���^oy8�I�#�&��l�bo��\a�9�s�^D��Ǻ���s�oFA�p+.F���rUu �[��ܛ��+��5�ܧ�WC�-�<����i��'���Ρr�ۉP0��;���.�Pj�
�U�OKUw8�����v�1�g��	��y{#�h�0��Q�y�׼7�Oj�X�,%��*����]�o���"5�L�1*dS�r��z3R5�n{�>�u�Y��J�5ËW}�U���s�bb%������b��%#��2�fv̊��׽�<O��&t��zء搏	L�_q��m�i�8'!#Q���d�QD�m����V_z�\�D�ʆ��?���8��Ҥ�Õfz�Al��4O;��b9�&(�otj��\�����,Щ�i����T���Ŏ�ڵo9藨lBT��NJH�7{\�R��r+}M�u쥔 (+:���\U^\�S���v�.�mM��\�&Wܣ�P�yǅ��Dk(��:3���N,{������3����ԓ�j|����U���x��ي��a*}�������c���\ߩm@��BB�3+��wR�<ŉ1����M*�;i�M)���$�rںN��zf�\4vUm)X	�D��}6��'#q\�ͥ�ge(^��=�"�)�B�±P�.d��
{�ߠV�T��r�
���0�h�i�A��=2�m��}�yYՀ�[�÷c����լ^'��=��E�$ߨY����=$@�{`�\��Өbڨ9�BE��9Y��[��5�7�z��7|zoX�q�r��בԴC��5�K�@�i���C��_A�$�(Y��=zV��{d�ʊ{��"b��r�T.u�_E��g��b�k7�S�ڑ�Օ|�F.��f�牲w/r�c�ڪ���Hl�k��"O��\�������y�UX;O!�s��
()�&ڇ��Z�޺{y:�����Xj3O��5���g���nI���9�����J��!�:�`:�� v.�Ob��������V�^!�H�ά���� �5I�ҷ�sI虚����s�f��گw<�9j����r��{�)��H"���-�����|z��|Z��"����.`�"�9�_G\�ϳ~V{�c����s~�o�ݓ�3E3���GQ�L�Q^�ݙ*������f���^-��nH���Խ����3�}�7_Ї��U]�trĵ_�{�� ;F�Jn!����z�=������_F�1�Ys�1��*&�Z/��-Hn/��H�����}4Vo|��7�fZ��ʥo=�_A�R3B�&!�c���6ݬ�z�9wk!��)��bD��ؑ�WP�jd]G0�"=G�D�����j�v�;�������W𚍢9�+��_�^�+ɘ����%��v!�8��C۲��s��y�Y �q���X]@���,H��k�e�����s�M�׷I�@dw�y	ͨ�=�9{�ȵ�^D{����C���G1�0�v�6�-ٸ����&b�=��T��qb��1�{��kz躁Q<�	�BE�$SHv/j��@nȷq��D0[�OA{^��S�^�0��J��������Oᶫ~�<�@�>� \[@�h@��=D����D�ڤmj9 �J� �Z��D1����zS��C�{l�G��3}[v1z���_|Į�����#خ7��1q����Ŵ$v��Z�w�H�`ۅ!��jr薜����!�:6������W]���+���ׇB�7;
�\�Z��:��Z�A�\3V��[�l����
�e4z1�!���Ѿ��p��}���12��OFo3-$7T��Z:6俺����`�J���ښ/�5n�U��gHD�����졭v�S��-�d�0<r��u�qn�m����.�z�x��	��zb�6�	�@�eR���H���vԆτ��u�T�?k�v�V�wγ/>���6���;�[T9���!#؇!s�讠Tn�v�E{1]�z.a"Ov�f-U%�v�zP/�e�E����;�j����n�3n������65IȭF�́�SмOA��֨I�}�d_C{�Б[C�h�C5J\�l �J�bMNM�}v�λ�{��튈�-�P����#��-�Rv [X���V�*/��;�.��/a0����nj�譠^�ҏ��k���>xw��,��#�% A �L����Y
�Qy1*a�#�!�R8��_ٳخ�fԾ���Kh��s4��辄�<{=;�����ƹ�{S����㚲s-�`�p�^E2��A3�r���&a =�l�.���©L��[���Eu6�y�H���Y����u�����;efnw�A��a &���)�;�퓸�u/w`�M�rwv7 *��.b�����!x��7�����^-��NWukޱ��ޣ����x�xk�BAs5q}T��C���vT1��7�uDsޡ/3���W��sz\�=�E�u��V���𥳐�-��Kży�7�q�$Wpo��w8j��{T��jø�jv:b��v;{'���@n9��ܲ���k^+x�_����[=��=�r�ds�<)���E��.Z���Ǩ��/�^�+����؆`v	ؗ���޲����q��x_5�Զ�nW��\��
��J�!P�)����Y_�#67�x}N�yE���=��k+8O���a��ɳp�Q��%d]
���{�m��ʼ�#���[u5�	����ӮI�ȃ�F��La����J���)'~�$�dmsۇI�otD���q�>��'>�%D�{bG�]���w	��E�rZ��B_�ew �]�#��T?�?{�����'�w^>�{^B�^n�@w�K虃h�ݬ.�TK��@��i�u	����R�����Z�R�z�xn"�������N�oo�Ѽπ�|>G�{��݄�����#h{Kȗ�h�p����K��	�lv�P[Urؼ�\@r蘘;i�u�Ž�^���k�ͪx[�<j���� ���Bũ�W��1��3�ps}��"��;JZ-I{��*/a!"y��O��*�/�NÇ�m��J�O���-���7�w�($s���9D/jW1;�����W�n��H%�I�9�hHo���D�k֬~�k3��}�vg�ǉ�W}���R;�{!�5=��� ��e9�	3�/�d$OA�Eu��n���b�d��A-�bݱ{v�����~�汮�A�[U�JnP-�%�ۢD�7�-ed�]��V�l�<�kԾ�x�4�����g�5�ڨ<6*
����cw��Q������G���r�@3�I~��zP/�Ԩ/��9D�y�-ʠoE�Rr+h�-�ȏ�����+[�5k�t�+X��wy�w�Z�𽋉'��Pw@�$G�i�C5JsݰT\ŴOr��%@�*#ػ�c�!�� f�B�0v{���{^�Ϸ�bִ��=��tf��.��轄��v6��+x��l����1���CPu/>吨��L�v!c�9�`=�u�jլ��fn�F�u?p��h�jH�j..�K���R���t�f�15OO#�Y=3�*����>BՈv����*bvwwv?W1��{q�3������ɑ�r1M	k�k�A:��![Z�M�"F!��-%����ڒ��xzH �S���8���hZ!�7������]�E�BE�hA�_U�#��~s�����1�1���W�1�Yu�Ƴ�N�׳|祽�׉��)E�{�3�ncV{���А[�V�=��M�;�F�9�z��~#���)�=���"/�5����j߱Z�|�cQ<w�\�}0����j�������/�H���Ǭ����`�,���1q=�/�Q�ȴ��>�������v���g��|3�`;�=��W�j[�Ł3BE�qͩ5�y	�M��[��-~�}T��4��ʤ/F�]�d�}��zׯ��x7��C��<r�M�9u@z8�w����Z;�b���d;0{	���ؼ1��^@-����Y�%���sV���TWۥ�LCq̓�\OG<�$F��ǣ� 疲��Q�0��GQ*�L��<�{Q"�#�=���un�����z��9�p֯���7�{����]-�&' �������c��ۍ��{1�/{e�E�̼��$v�$W�7|W��BW9�z�ɿk�����żH������wT2����,�`��옇�=�oJb:�\-Ob�������.��5�1��ym>�o��ʦ�.U۟|��I��!"�_Z� �]�.
��C�q0�޸��`���b['#�%G�C���ހ����Uwb1��~��)���r.��8/����J�'# �TGV�=���oCȭ��ȦNPH�)ȗ�#ط�����d0~��R_gQ��Հ�s#j��:�cj�Tr�]G&�q�؝����GQ49�r�V�t�6���Q�gtL�>}oz���1���йφ4☯�j�&Kw��OOR��~���ݙ��I��/�k���*b�"� ��ֻ�r����^+���od�{�3�vሻ��v���n����TNBU+ș�@bjڤ7�����#M�`y=���gs[X�@x#�o;UF[�[��n!����`Z/astv(Ho���+�h��=0�킠�j���e=�\�#輌�hj#����9��g�\kǸ���s��h�ME�{&�	D;	;�}���D���sT=�]�QmT�!�� �#�����8'7[+�����Z)�x�#x�-�IȎb_���8NS��؆�˨���H� �9�'�J�8�lz!�QL{�S13	 buΦ�1��c���� H���8��P�:��T �\�}�L9����Spm��w�0}��(��.�Q�z��=�e/�BOs��#zrW����|�����F���x�l)��H�9C��.#���^!w���C	T��+|��/a"�T;�r/����5�����w;�����<�b9�}��ؙ���=���6��R�+��̀�ރQ5����5�q�$Wpu�Y{	��o5���|�~߭�c���*��@5�G�R��z7���z�����;�]_F�;z\DuFA�A*&`Z/��!�����OsY�ݳ�k��9ofO+h>��u�R����=�CE�;�����@yD;E9�ۑZ�~^ďb��FE�q浻k:�-�ױ�s���9������P���7q�+���/*��Ʃ}3�L��C�q=�ݕ9��y�]����u����aw�ON������<z��sj�K�;8	��x�#(��K�Qu#2o�+�Ѷ:q�_fEﰚ���e��ˑjzŪF�]c̏TE�vxZ��W��\]�]�d3�۽��7m�3s���I��W;��u�5]�B��`� �㉷$�*n H,�Ȥ�H$� H�!!!	$	@+Z�{���o� f B!y 29������-@rȷ1��^EŽe�G�Ʊe�L����G�/�XJ��������\�ֱ��y���M_���'"�;����$$W�,r���I�_U,�n"��tyŽa����z��# 3�y�i;������1[���<֬����x�쾁�����>�P=		���UHص�v%A�V��T/�G�b������>�u]���?x#�|�s�|���Ǳ[��nb	���v��8�hH�����P.v��r�UB����Zr./K؆��XϺn���o�_��g{���On�@{OG�oN�s�������޲^.��a=�'��-�#nО�P{T�bq�.�=�X�9ɻ�浬c��oW���J����.�5s�>��:���!"r/�W���Q�����H��bz.!"�)��T�=�	�@�pk�97��g:�1��4�"��^b��A�N�j>/�ȥ�F!� v&uBH��\�"���"��������Y�r�Xz��}���߀� DzL>�>�_F|f�7~�]WM��C��zڣ��,�I�I�8��[�~�0uj����y��!����k䪶Ն:�wUM����;7�X� �����Ó[�?DlLCj+\�޽�EZV��������t���b�Z��v\BƨJ3b�<�2�Z�S]����e�w�	�8�x4	#:������=)o93&=ШVn�bE8&`o^i����sfg6�y�ۓ;o�lG$�x�p�J�����HT�x��ߣ5��<�Q�:��}�i���g>O{��5�TD�	c/V���
�J(�!)_P�ovk�zS�b�'��{\��J�p�.�T`��V�2z�b�u��IZ��fvbɬ�{C�C׷l���:]$�ٹy����\R��Tj���7��$w����27ۡ?^=d��<��O��JN���X|�]{J6jp��H��t�n1��Y�/TJ�ޭ��Ih��c��B�[9��F����J�<}��L���݀\:7X�xE�Ώ&E�ۙ׆�.��)�x9��+Bӱ�2��K��>�R��Ig��n�
I΋�A/;kEoZ�/yX�$�b��[hQ����ﮞ_�;�s�	�i5{)*�9VH�p�õ,��'.���vn���&v�VZ�:�yR:���`WbC\U�Sb��١�i�[�,�62����m��R{��r��S��*	{,�.�Nt���V�?��gw�I$�I$�I-����O���p��v���	Sk1˕�hjTц<�pӔ	;���y��r��à�Ǘ)^�j�o���1Z�����7\�h��;�4��R��K����*QwQ�
�'��JQ���惻�ș��gز�T(ӉGuQ��a(�x�����ʻ.�0���ni����<�F�7 P�^��jx��U��r"�v�PmO�$mؖcj��*P��y�+Zx�7���ᛇ",�����#���;�%]���c2YC�tcYٷ�5��P�6��7��']uҋ�W�gz�#�+�"���4����l����Ztj�:N�u�]fM�<��4k�� �7(e����mR���c0'" ����S���ewK�0/��T��2�-pQ�wV�b��ţ0�f��Q6�����W�r��l�Ѐ�KtU#mh�2�@ѽ
�����IMpJ�:�R$Q����WH�{wR	�MG�5��6B����W`c�w,H��O����jSF]�2{SW�$�x7&i�i�u9(��|2e#$1��	MR��	$�Y��8���=��>r9&�o\mrK{9rK������Y�H��c�= ������S$FM��F���>��H��y�J�ɚ��I}xl��e�!�VT+����>#���R�'�����>6{�J���G�i�[a2Me�Y�qP��7�(�ݵ��t>��[.H�3�F�L\�����g3la��[eݯ����ilG���{F�$ocm�}����E�dhϴk�|%�!ZH��tf�X���r�jMm<��y�.MB�R(�+EB��DVv��(��IO!?�g��\l�ǽ�//*���\�g�"���.���[iO���!�;�U{�ԯ"�{t�M����c�o��{�
��bm��<)&�ʄ�s�[=����#2O��[����yݛoc'�˕��w�[����g��]O�B7=fk}{{x��{,>1��ӎ��F����+��&t��H!��t���.1/6�'N�av��h�m*N�n7�D{�aܕ.�c���ȯ�����G8�N�d��υ�g��ԫ�k��`*
/�v>�Y����NSY;���lDj��|&�Y�N5����,���8���]y!��vciL��"�tep�O�"�k����s�3��a�1��ܽ���3�܈�#�Ho3�mM�S��nU]9�'|�Sln�����ϒhE/�J�0߭ah<�o�Ӳ��ͦW-���[Oצ��P�#�B�0@:��^;-a������%�Awh�~���yC��9�K�:������:L����}���{b�}4��]�s��U�V̷$o�0���Q��R���L���D"��<�P�=�'֣e&�ph�@��v�hn&�r��mT�"����=2ʇS}#����:�;��*Tؚh �o>��]�`T捷Ϛ�M�v4FQ�.�o�R\cf�L�}tt��c�rE7�S7wb�aJ�͡�n%t��u|��eXm�֓��·���=ѷ��j��*7��.� {���aថ{�U;Yn�#|Apt�~Uz�{Qf�Ǽܫ�Mk�%#���f���CU`64�{êp���Ջ������wOl=��o:˫�mB�Ʀ!'e�Q��05��5QO��^a;�1�ޯO`�:��C�b�Gv��OJ�q�`F��NL��bs�=�n�Y[l�7�
i��s��K^���N��|�3�+!k�z�ĔE?`p+'jnf����	���R+�z�5V�Ǘ�Ry����I�Q��PBl�7%��ﳙ�ֶ	%S��.��9>C2�Xr�X���Y!����\�B%3��Աɸ}��#YY��乵L��3q9!55Ƅr���P��[H'�719�`���Q���է���l`R��I��W.�tѻ+�2��O���HS�躆�(of��0 ��.P6��G���$��׿2��i��<�kq�;������qS�dBJj�b��#���뙧f!�Ԡ�o�vq��^�Hc\	WgdjI߿}�=ᛗk[{[Wr{D�_��W�������U4U��,W��u�KR������)���s!,���R�'T��F��fkI�Om���_�`'���TYSk�#�F�zv:����=�/WO<H��8�܂�u+�>�^|�Z�++P�K��ާ˧1R�,t��8)��R�@�+F�2 �ۅ,E��v��ٓhs�	T��
��b�N2&c�8'���c1C���5ۆ%@R��`�$ �S��M���-nE͘����=8�թ�<�w�S����uˬ��:���<��}�yZl;�<2��K��E��[ȼ�M���ӵ�^.��;�ҧu^4�nm��:�ɚnEBT���O#�qMF<S��pu�n���u����S��I����b�G�Y9Q�7C�͊�2��U�D�C�vv`��ŵ���\qLh]�]%#���vZ���ī�F��OM8��M�f�]U�45@�[\���� �w$�>��T~{�<�uk6�ZŢ�1�����U�5Ђ9���j�T���r,7��#��RN<��B�qAU�����H�����c�${;n�v�ا�;�m�a*����ذc4 ��:�sTO�����']�O�d:ICa�j�V<��9ΰs8n�wV&�w��'�`���ޑNz���x�{���>�W5����ՙ�i�h �����
x��N��X��7�s��޺so�%5S+f46̿(C	.1�=t�f�s,�{��r�#�⥎�Tҭ�N`l�e�	�[�'�rW�W��R�̈�y�k'����m�q�CO T�d!.�Ӱ�Bvӎ�r"\QQƄ��A���XT
v(5d�~�e{�N�Z Z�C[�4<�O{Br+��CY��J��풨؎l�u�_�XXS�q�b��ݘ
���<r;����x�J�[��0�$u��t�{�{�ܬ]v����XY��}�J�Q�<�]-@B���v�H|<< �t����jH�4F`�싁�`M���kÐ��L*�V��Y蓞�\���"�G�֨�ߤz\�rݍ�AD;��d���{ �xn��]��_{@5������;��z�?M�s�yV]oJ�ӎ�S^��'ys���`]�~�iBبs[�s+;5�XJ΄桍��s�V-w���uz06��������[�lh�.�S&���#�i��Hд�<w@7YK=V���nm�ir��!>���E\[j���V$s]-��6���Ϧz1�f�v�Z��[����;�'юi�T�=mG�*e�눮]SAH�yx���̧�s��\�a��m@�bX�;Q�{t[QUW]��Ѽ��֥���[��5-�2���Oz��2���'b�!k�gsO�^ݨe*Zt<h,�vc�����iX�}�̘�jأ�X�;k��9՗=�s�c�X*A]�w8������2��<�JS�/LnF�d�7�@�p[��b.ك�c��ߟW�x�������UWR[=�+UG6�e{�p�*z����F-^�G�nOź�~S��t"n}˺��9*��#�
��W��Tղ�s���(ǡs��Ԋ[}��Ի�*�}�۱p�Y}4<�YY�E�U}+���xsF��ȫ���c3T�:�Wr�0���G�M���1�7�ܨVj���mw.����&=�1�h������	�3S�Ls���9�8^�U�yvg]�e�)6��Bt(���HIᦍć��co9�by�������*w^r���P;Mo'��]�����,��[�LSTF�V�Tb����r��8лL�s�v����d<�8�;͹$��ge�}79�CO?���n��]9�)��W?Q:G�Ot��[��Bt�����J1/N-�w�\��� �rt�{OUp���� �G��:�Ǡ}ƴ.ܹ1��,��sR�p�W�����0�:di�w��UR�b�w M�K�В"z�+�*<�R]��xxBﱻ�Uo����˕�݆���	��d�s%�hm�m^����ivܘ�����8���Ü�*�TqJuG|�V�b�&����`H@��zm*z�=ѽ^�W@.�T�\�C��>��%�|��0vc�|�r7˕(��20���$�5�y[<ռC��Q�}B>g|�Q�s�^߱���ι���N�H��FrL��u�����g� ��@U�=S����	_m�-��l�QwI�\��+��|�'�CN���CJ�H��Օ��펃�Sڅݎ�ኻ��z�m�y�)B�p�����/�vx]�J�z����b�)a����*p$��e!
G
�^�.egD��9v��m�̐��f�J�b:[�¢���-3!�2w�u7Y��W���5�&=|φ����l�i�<��� �P���C�*�6�\�����:�=W 2����-��wIńH����c�5u�n����5�.�H�6��_1RL.��8^�8�L������΍�R;ٚ�YA��[Ov��FX4�ViͺY�,��� gu^k0��ɯ����m�!	L$��|nA�(,1�Tn��e<i�}H�G$Θ����:U�.���Gc��״f���Z�sxw���w]�o��vb.�R�tݍ�/[�EJ�%�^���Q��ګUl$���:��L�nEB�eE�ʧIn�9u;ûx�ny�z��-܊�X�A���NJ��wL�Q����׽���"6$\���s��x5=�q��+����x�h�sO�9y=2�b�cf����J�n�}�($������]�}��:E� ]���ޗ�)q��TbV��7�s0���@��*�n9��ᒡ�BR�O���9������N8HI��=�Yː�ZX{�s�\64��(C<��+g���qyY]�z4]]4g��2M'e�\�ĲM���B�ι)�k�#`Y��8&�+�c��%f޴BK`s��2o.���&�t�/:uU
X�J9Io%�{�xx�,ěG3�s�=Φ�uEy�2��1���8��~txLt�7��ΩɊb̫�nWR��lؤ�zR3�p�E�3�S�b*��5��@)ȮUR���T9�Н���	S�ǉ�{s<''My�ˣ�̣}�r�)�F��t5�N���V��n�_v�!p�F��M�+r��ޖ'nM-�m����Y�#�<��QpP�u���V�˕C�[��b��[W����qCN�����c�F6���);WB^�pl���s;ع\̝OcD����=���i��._сGfUd��*��^>�o.4E_1X��_ZJ+<ոt7i�F:��=�L�ֽ�%:��u<����4����ԍ�^<���\��_^-2�s�ށ[k�ͬ6�!%Y��GP[�7�pp�M��aR�y�xARQ,����jv���W���K�Rڝ`��Y�^�;{i%�b�n�͊}QI�-���wl�"���|(�����Iw���;e�&�Ƭ�*�"�Ƭ�"�lԧ�7��rL��Mfs���j���L$�R���m�G��!�+��kJ��Hȷ<�ۑ��v�tV��>����Fv�H-�D����o��yMry!����#OA��%��:uJ�)Ὑr���'�+�h}�Q���Ӫ!�Y��1\�����Ơ�ﻯN�w �Z<���z�ʵE��_r����b)_u�7�F�F�������Y}���e.~����m47mp��4v�(ŵb%�ǵdN:�^u��;�&(��ɮVw%3>B4E��1�^�كޣ�:�|��ێc������F��yas�tE/~���?E�/��HJ�󐑢�҈m]���()󆢽gw���r�є�Sjr��`.uqjq�s9֑��$.e�}{3�J�c�]�(NՌB޻�1������!�mN1R�˱eSva�@L1�ĺ��i����V7�V���ywkx��s.����X�=F(��,��a��Y*'��{��C����/H�{��{I ��Ζ*![r-E�q0�r���r0�r�gJ�*�j���6�F���wn��p��$RM����y}�J"��Q���������`���*�,������a��M��:�uݙ���kw�,����[�����#E��ԁ���K�I��UᏗYѽ�5��E��Q|E�ݦq�dj�.�[srVG��'��%/�\��B�*�T���p1�D �����M��M5KLb�qhq����޸V�F��[QK�Elۻ맋�nEzu�Xq	hov�e	yS�+/j�:R���Kw��9	D�0f����j��R�����h��'�3&�T�k��^��⥷uu��|+X��Ξ�v�p'dM �p���;�h�{�$B���Q�{��S紱ދ{�n�gRI��{0 �ȓGWyu&��:�n�#|�:n�X�d�{����yO���c�-m̮���I$�I$�I%���՝="�N������9��N]n���N�h�"1�Gf���Q��\3�6�]����Б��^����)����l���%Z���ڹcO�J���1;Ki��'a��i70ͼ������e�L].Ժmm���
���� �a4�U���*�����tk�B_�k6嶅��[zuҠ�R��|�^^�c
��9�/�(��w�����93�{a+\���e���	�k��3���FT��Km�*���M��\����Q#+h�������^+�dsˏ��U�w�N��k%�#u����l�e���ķ��YF���D�Z�>�9cE��.��`TWj&��s�+q��6rU�涝���@�����i�`������{����Wщ�}�
��`�ۖ 3��a���y
@�Oe�����n��{>�T�w#J��S�'#��;{��Lu�)	t���Ь{u��Y^��=��d��0����'.C[���r��*G}�;�ؓ�lnI�.U��rJ�z��rIgv%�%��W�͘�]*�T�S�f��	���#����?�gL@�*w�G(�D/J�C�0_�D>�*���^�$j��=q�$	吐"�S�Hd����h�YTzK��]{��f�i&JIy+��f����%��))22#���O"�(�KR�T�9����tQ%]"̬���1D�K�I�<��Y�eN�mk	k��l�׌��D"�%H�.yҘ��Ȧp��IQ��g�z�bmZ뤭`��/H��� ��B��0�]H�g��B��W�'���̼��Լ���nu��P���M�E1s���1m����P�z(�Bt@e�L��S�*�i��U!W+�>W���ad���[�c������9���GT��e]'����bb7�®��(u�t����}�#��J2�ʉ�t\����r�v:��'�����ӱ�<��w����;��J�o��x�2���&n�v*�4���6ugc��`w.��)�]*.,S{^��7��j@�AԺ��#3�O!����[����<��	����b��45ݽ�
��=������,%���E��ݠ�8��'�mϣ'�ױמu�<.��g^�oDeȦ���۵�:7�aZ���-�{�a�l����GF)�)t!q�n���L����b+6%��|�nA����u��V1�x�T!)����y_K��_V�?S�ֆy�� '��+�=�7����@�tp�o3g���5���aK.U�3�;���T��Qv^ۨPЇn�A�[��>y�szp9_:}Esm���:�y˳�C�mq0k�C��/��Q��4�����̵�
�^+�ku�"C��&�$��@;�E�Z��}I����;�t�)+���1eoV��_t����ӼHr"�JO椏�xx�[Z��J�+��������e�G0#{Mu@�"�F	yUCbE%]�c2��SJ��۔�$s�B�K:�@h�^�<�E�/|'a �kܮ%��;-���N�	L�B����'	�����QS�q��z�9x� �t84n�ف�,-&�TgF��k=J�s�4�E\�g(t��`�%��	=�Ӻ���z�s�ZA��N���xĮ}��X�gk8�ڙ��Hn�u*�e�w�:*Gf"�Uo�[��<1uf˕��o��r�j�m[���U/浻r�nג�NM7yQ̦u>��S��+����V�5�>\������Ĵ�h���k�[��랷�[���9�O�[fE��@w9�N<n�_8������V)^iѦx��\gHa�b����;�>~M_��[�{-�`�
4����$m��w�9��c�;I-H6�o@����c��mF���諭��N�x9u"#���k��g�23���p���]rC��W�oy}�x��4�#T��M.=^�j�*of�;�&\���7)t���>��.��t+��[(.�i�S�9��.�k������]NJ��ĎzҸ�8t/(C̃�5��]Z�D����Đ͞Zo}�@j����.��4̀���1�Ľ��I6*�wV��q��@�����U�n+fӘ�C���Py������w"u
�)���\ꄬ3Დqc<��jN�IT`U��b-7s��/D))�*����t�an�1�:k`�:ĮP��%����9�\���	���ұ�E$d�p^��o>�&�N�������;M�����_٤�n���jV$�C��P^�4����W-QʌX���+o�J"���r���T����e���g�A���������zp��j��Ǭ��̝Pc������J�.��s�7u�v���]4t����]�o�����՝���]^����v����|Nu���R§cb{�.�X�.�}Z�e�;����Yݎg��������]]������)�.ʹb|/�ާ#u+���Ŝo���ֹˠ�6NN��[:np�O\ZصN�E�"$��Z�%�0'�z�P��B�C�������:A|�����k*���a�}]��m8r;0
��Q�E!�\��u�Q��k�����eM���9*,�4��'J� �^�|74ԅ���ź&��z�u�ų�c��z��d-:tpP��b���O/7\X�v���L��r��[�V��a��Vl�Q��[��,��<�4Z� 9��wŹ��Β��6�/u4j�j��5)j����o2"� �;�k�ڇlgiӕ�Z��B��S�7�%�֫K	V_���tl��3�'0V�sS�F����8�����ݔ�]k-�`g!pr�(8�ň�35ZRG��}�W�ݗ��vu_�����p8a<��-��jm`��j6]��3Y9�}�o^�z�k�co\%V�= K.eD�O���6��uLAYX����
����x�b�y�����o�{��aۡ
f)K�MF̘q����4N�	{�<���s����뚪6�ޥpʞ��[��8;��I�h�`|Ol4z�J����r�G��mz*�Sy�(W�1�h������\�q[U�{i�wٓ�,v`�K��c揳�=Ԫ>�Z�y�����2vy=����O����چ�n��Uzng¡�<0V7U|�.�)*��O�z}���^�״y֠���n	C�1�}�c�m�rMd̞k��Ar��ya����x�䮬b�;���%ޫ~���}0�����c����`����t*��9=ߊ�(k�o��+F�A���N�|��_m�r��\�e�W+q��S�lu�)�3LSy��G����S&��{.�J[*]2�8�\n%��8�@���4�
����Z�߼=�ym��R��q�>	���_ܷºw��T�v�R��9No�^N���D3��O+��C�>�]W��v˓���Ŋ�/Z�˒/w6s��-�R�L0Su��]��\����f��5]�ɗ�x����p��� �29�r���m��h�l���e�����WO�4�{�{�[L���W�78GP���%&�wѻ}�j�y=%��G�::�O��8s��)���y6�wU�l����>o�e�e�
i�W�3!U���L�vt�'�{wMtYR$Ej
;E�R���#<���F��r�z흼���jH�⨫��Vϡ�V!	A����ƜL�3$�f�PzAdl��\�5^�Oϫ�^Sc����"Mk�R�1��%TY�9v��:��׼�lYuy΍Z�vۥ�.V��L6���9��L�]vV�b�����7Kny3k�v��� ��;��ݬÜ�]9`���wRҦab=�R�[2���k{&/&i�Vp9�	νڧ�^��{UMi�ߚ͹���x��X�5Ⱥi��1���; �:�N�֍y[�o)뼴��,,S��r�����/1�j�y�S"�ٮbE�dU��|�-���
\ve�& ]�/�m���MȎ�B7����=C2�#H_���|���L	�~��wS���S�����l�����=su�=��)��C8�E���V���4�C�C�9�8ʊǺ�7�П�ڤ�8��\E�ک]G�<.�'$�ׯ;9yuM�ofӉe��w�co�\�醙��0é͙��3n�[7�%���/f��Oa��)�NL�R?��q5Ӫ�o��J;�&��72&7n��ޭ�ZY2��X�cv��ܛ��t�!��B]a��������a���V�6Tܕg�nY�{r	��Fy�T�E��7�%1K���>vw�ʋ{�]�v\�y��%������ַ~�1�e���F#�7���T�9��Ww�n����b6�}��Y�������8���~�le�	KxFM��ܮUzj����37�}�]��R���p�U������92�4`w3YI�˦�*~Vw�y❚|t��DGZ��u��Hz�˱�o��:��w�(W�.�	;<7sO���c�W�L����Rfu�R�#!�ye	��e���m���y-,�|j�*�l�W,<[���JuX��6�U��xЬL�S�J�k��x�^��t�M��w*��k�nҌ��=�M	����jFS�7t���wU���^�c�q*��n�Wx�^O<�h�,�w'�-�<�g_w56�^�IÑ؄��G	�r)�K�,FϢJ��m�����U5Yr#{E�kW#l���Q�#�ej9�u���+�Q�q͢{eMJ��0� ����x��ZfP�dp�ƕG��4gU�Kr�w-j�LŻΘ�I�뷜�m����K2�����~����;)�O"d�Y��J�>�|z!�r�P��2��W��'e	�V��1�5������L�����i�l�X��F?��D��{n�a����{�\�x��t�t&4ǝ��bֆNM��֎9Z�T,|����ҙ��qo�9�:g��ʈ�R��¦5�d���n؛R�AS�MG���ai���ڭ��}B�E��^!t1E��0��z�2��>")>�6�7�W���k����J^�Ǝ�	��l�����AQ�+UJVMG�^>M�
�����*/l��9p�(��g�G��`7�S�3���&`6z�2K�ލyV�9y;��
�G���x��/�ʉ7Y��\�w����g���]�\:@XC�W�zf�z�DO}j�m��i���B��D^�(M$�b,51�%$�f�{��$����|�#4L�ȠEp�uĔ8l�e�Hr�����9�����n�R@vhX�����5	������D
����*҄�>�'f��7��5:��W5q��%Zn;��+�v�1�\ba��J�E�utӡ�Y4w��O4�\��IE��֥eUq��.��j�}��a��h��w"�Ӻȼ���C�pU�}u߅�~ܔ\c��ϡ9����M�ړLl�*�]1l�/>��{`x[�^.����Inc�S��{O�yƤ�ܴXl�Ϫf>U�:/��_��`�V&�r�kS�<"S�y:�S�.7.�vg���J�G	,J�E#�c����#�$+T߂�h1��Zo�M��o���s�Aג��ߩR���ڐz���!���Y�GmN�v.S�o��^�N�V%�\6���� ��KD?���3.L]���L&�Q0�¥�un�
�fd~���`�J����%hWN7���谇�ޜ�,��A^������3<��B3�����;�����[�4s29Cj�nF�J�ʌ��fE�ć$�����
��`v4!��,��t�!Ꞿ5��*\�4:f�+�8):�"��0�'þ�E��O�������$��j��Ε���`[�n�ݱ:���)��ɶo--_kޛ{�3�������r��
�SRI��3��P�	��tER�`3�{��A�x�wV��<�:F�ȓ,ᄣ!���iY��br �jQ%I�*�� j�7u]	3l�28Q[���� C�B��cթU�EN���ѱu�}F],�NR>��d�m���>gmˬ�+�m�;D;��-��3C���ı�L�gk�)�&-Sr�7��]�ө�BՇ62��u/��@.N<��|m�����"��z��4h7|�ܩ��:��y9�r]��R�Zܦ��Y��z�4���nZϰ-�p^�i�w$�-��&ҥ�H���"+q�sO#��9u�Qaԡ�
:;B�I%� E�ʌ
�3UEB�m�y��w9	kU��,h����:�Pf*���1ݡ�w:Ɋ ����mc]��V����i˒��Z��ʉtWٔ�^^��=մ��������ſ � iv��j�}�q���fçw�9�X��D�
��g-ա�9N�33b���)Y��[1�j�-0�]g�2�fAqP�ؘ_nP��ʆT���&��%ek<��\������A"��;�W�]�E"��M�E��w:�5Ƀ��i�c���z�=:ng��Tۊ7$�I$�I$�I�.M���*��fev��]�X��9����U�%@Mo/-Z8��ug��Ptӽ�{%��ۘ��|�_g"�N��c��cOcN9��� ,#�ྉb�;cDϹ�<q:=���f�-�j>3�\LBs�jG(؊H`J�Z��f-����]���]N+��1�xD']b�T�3�2�l��J�jE l\�peҶ	�3�諾���Xh������e�j	���ۤ�ȓ,�[JUC9ٓ{b��;����AH �����<��qIT�L�lu����뵑&v�:P�}JR$an��*��m��F�^l�r�ݡ�Y��PB�f�mo.W-��K��L^��ef�	�[�%��W�b�d�ʲ�����h��,���R��9[Ƕ�Hq�u��]�vYx�U䧱��[FR�*а{7����KH��0J�z�B�^���OZ��زC�
�i�1�}j�rRJm�y'p���ӗ��Q�V]�Jn���@owc�N<�,9Mݠ�[�:(.���=���l*�Xo��A��L�u��p��������j�v�b��$�Z��I�����rMI�q����E$�����>�C�T�R�T�#�/J�]ҷ�X�y���"������S��9�TiVzy)/��O���rJ��M< ���O�D�'�ء�a���HV�jg���U���YjI���*�A�Z*EIQ��y*hQ�R+�W!�����J�FNY�HQԮ�x��^X�)��$��Z�H��������C��u�]� �R<5R'�/-GE6B1ʲT�)�4�a�M]4=6e����4�$+�t�"�/W@��IȲA��)ޏb��t�Bk���_ˡ2��%�]�[��b�"��aU++(�;t	�%yy*�i�9njW�QI!%�D�BBR�3�\���]`�$�v�#���U;9�t�ۙwԬ?�W>�a���ec�$a�P)�E]���'o�UUWȩ��=g-PV�?J���ك�_��U���r�����j^��*f��]n뭭�GX�e���K��DA��LK��������X#��s�.�t�8�f�.��Dr�{�%ԣ຋��J��G��>��6%B���s�Ύn�S��gu�m��� ��z����.���U��><ja�]��㼤[�ͮjkl�a� 4�a���������q{ zH���L�;n�;Ѱ�.f�ܼi�����Uu �>zn.e;�4����'B����3�d�mx��b#$�m^�SRȡr����̩�Kq���л�l�BȬ��AQkPC�Y6_eV�.Q�o�� U������:�>kՂ�{/�ײos9��u�s�����:�Uj�*؃Ĺ���r���
�"T��֌۶_���Sy���}
��bBȨ��WWZ>d�(V���a0:^��+� ��dͻ-Z���˙?�����,�M�V�wٔ���߼�]aLN):JX��^��8�ƫ��_�J#����[Ǹ̈́��A��c#d�
�*6���Qd,U,�wdcu�)u�����ME�����9�H�X��������}�_w�Sc7M#���������h,���)U��?*/5!�T�ٽ��'��]1HͰ����Xm�k���yI�b4Y$�3���U���i��Ys���K����:db��Ҹ"m*1t�,����2��^,��!�V��^W]d��[]�����N01�8/�|����!t�{Mз�
�3<�o�jN�'ʋJ�&�/���Av��E�*G>|�U���vh*�<ޭ�7	�t�zzTC�J��Z8O�S^t�ظpi������_�\�%�A����E�(p�	�嘤"C�{X��>�"+%ıtT;��ع<��U4�fc�=fP�>=�	~�pY__��]��b�5�v��~�t}H\˭M���s��܍�b������A����~��6�v�l`���O�ʈw��d�eE����T4�d��^�硎f�;Y>�w��oi�|�Y�}^�O������+�/P���ҙ0f����w7y��Ɣ,��Y=EI�Ti55ܑY�-�����v�u�t*��\n��u"��Ӻ�����V.J}��*�:'�y%� ��Sk���b��~�gzbfP]�<=]� Cڤͥ{o:n^ĵٯɹ�[��/РEHjm������~Z�u��x�ؼ<Ui��3�&%��7������B�~jP(Ӹ�p#,ʡ�+_��f,g^����pq���~��X��N��/7c�ׂo��/S��B+����x㋺=��WzrIi��
T��{�����R���D�N���)��z��St\q�"8�WF��w\�o^*ʵaש*����h5y�vl.��,B`�9H�9qO1����Mf���t^7�^��tJ%�LxT$�z�m�_LWq����S�uc�ޙ5B/*�=󻄿�N�U�t]�	ߏ/���ոȧA�d���G��#�9X�ԍ�F����*|)�K�.P]�/�Y|���s|�J9��Ϛ���Q�0Sq`�t���t[`��k�ɳ�
�kݽy�XֱT�Љ�6�#n����R���l��"zE�[���ns�Yz�N��[�`XE)���}�oK��w�A��zdؔ�������ü�])��Ά�nB��|�[�㳜Onwd�ڱ������qvu�P�`ԑ���4�"��k��VxA��:�O�ʙ�a�
��:=d#=z�u�z<�� ���Vz٦�a1��HZ
u��fp�P��g�ޣ�3sX6=WE�T)�q�"��*�y�,E-�!1�*zL�ї[I�܃�XY��E���\d�p�Wl�B����
�j��>;"��9�w{�,oS�+�ʿBGP��=���)d��G�޿	A]��h8�	zM���N{���[k]�gܠ�\ռ����hηZU��٧rc.*v�Ƭ�v��!�<hf�.6�p�T�^(o���y9�"Ύ�WN�R��-�ܫk���Aa1!���L�x�p�qG@��zy�[�5�v0�=j�e��;����a�94P����$S�Fк����6Ggk���Ƚ�b�![���9���0��X�Z��Z:�(8;�|.���1����Md]U�LC6^�*���Z�q�/�q����#���	]�QW�2l5Z]��ca�����X�*�RܬP��}y�L���sx��..P̠�G��Wtmf��4��q�]�S�odl4����r�9�rRG�U����۾i������tNؾꮈ�8�2'(]��۷�l����>U�Ɗ��ˇ���ۚ�k~�'�}G>�&)}_dQ�3	q�S�g�H?�v�~:�١�&5Vv_GMn��2o68ɭ�=!턬H���#�1t뮼��Kh�F�	�wԆ�돝ٞ���\:/�}
������~��L���&a� <:��=���Y���L�� E!Zʔt,�3�2�.�ҡ�
�����޹w�Oe�2=�F*�`� 	��g�����*(7 �&,9�!��@�NI�K�e:h��7p��|.Q��&E�W)["�2Yn/IB��ݵ9�]|����뮡|��
���� UL����e�ʱڧŐ%A�.6*j⭮|�[����DQ�����ݯ�X��᤿��:�n���Z#����u̳�d�Qx�����3�IHc�i
�%�3����P}�}^0`c�iC����t!��`Ү5��,�y-�4���Y���y���GzoI)mʗ�L�K�>��w3�F�Y��h��3�c5�K]1K}X;x%�L�hI���)k{u�1W<i��o[���k���#�w���m�F������5U��WUGLq�*x���+$ hdi�lJ#W��4��lb+ڞz7��w"��]�lK	�^�ܰk!�d\a\b�G^U��˗�<%a�-�x��>�	�fڭG�����YH�<����^'���Luo��f�����}e�l��G WD�
�]*UaP�����~0m��x{^�	9^����n�[l���4lWN+b���
����>$eGUu+Dg��5�V:��ٸ�b�s�*�f��c�p/�����ŉMޙz�RAfB��v��nN˨�9|�k�ap��{^�Y��'���4�U[ٵ,���]E&Y%ҳ˯Y�^��@3j�Ո�~���E��Z�q��A|u@�9�Pp��_�ݫ��5v��k�~���n����U�t������y����TXb�6;%�>^=�>_c�Oe���+z;� �t}U"�F�\�P5�R���D|oƋ�\Fy\ƕ
�b���Iom�^'��Nt��o�*�\.��_xf�>t�o��m �Ҭu�꽁�2�l�Iˮ��2��xr�}��SgF�:]�[ Yzb��r>��Ho�z��աr�{8w0�or�U���w)^�]�w����-Z��Bv��r7�i��N�5jY�k��Z�c B$:&�WZX�Gr�x�ڇ����)
<}d#�8z�=��{���^����ְN9��s��%̿w��g�C�?Z�N���#���x�畍�	Ϻ\:���%�B��ӲgU�0�ޥ-����]//�4�A�b�Xkn9�V�i��a�[ݤ:4�ż��u�q�}�.�Q��fQ,pU=��}A}2�=W�&z(��ѷ���n*u�\�j�\-�?lY^0@C�֫���Y�O���S��V�Y���<�D7������m�'��,�՝7媙�Sg b&�P�����n1�4����]��̜�E�s�7�x"�U���l��̰�S=s'�zbP��W>ǍzII�v��!�b�h���HױJ6�k�Ez7�
e�Xޞ1A�.8��ނ�t��KPr�E�QW�Q5�˱H��g���cAR������W�cÌTZ�LZ	U�U�,Th� �@�F�{����0���؟e,�0Ȇ��:\�S�r��o}$M����]���*�E��Pf�*��م���eM=�n�4�N�y6!�[�n�q7%:=˃�R����?����n'{ddF���!�.,�>�P$<�p�Q֝��u�*&�;�kn��
`q��\C��bt����2�6��Z�E F��:��NZS���0S��CG�rxR�4|+�w|B��D�7*xݗ,�B��ї����������*��K�]҆P{��*|�DV�4�T׏��/'ܨk��i?_w+	�+�*�c�w���VxA���C�`��?�Ś��r��5�v���
��&�	�2'��e��2��r&#!!��������qM�s�N��� ��/Cb�e���Oy4��H�"�PH�LP��-�^㠝�B��C���3���盧��p$Nb�����8U
@���L����v�<�u�;{=�=Q��']}���bY~����\=��l�Ke����7�D�^a�_�����r�Cӭ�mV�]F��g��f[�+��K7�.$;=꺀�yB��Q��c�
�+U��;I�`�m^���]�%h���aݻ;W�g
�`K=����VG�	8�Ө<��T� �k֪P�R����2[��#H�1��Μ���\�v��NN�������o<���'�T����R�P1��;�0lQ�R�o���0�n=��.�,��3{Rm��5I��hϬ�
\\|)x�X���8Oh�N�^�w W%&-�u<�p�BT�B�x�Bؚ~ V�Z���ʴH���y��7�Y�ܶ�:;՝�Ʃ�!H�����>EA�꼗���a�4:����D�SH<̞����B=�L�����WzK�����m &	��|/��||�H��;��4��MɭՆHa��*ORs4`������>4���B�/��;⾕g4y7�$�<_�W�����W맶�6�3�mU��3"�A>��|5)yڛ�$�z�C��E���*��O�o���WyhTߟ�0P�V+'�=���o(z�I���=&�v�F[��6���U�멥���Ko'/9�.J�L`�uw�(�>&+>D�b	C��� ��*�sP�����k�i�߉�75�]h�њ�eEy�.N1
�w��%kE �^8�*����[�ϴ��[{H���+m������?��_�<ڞd�}h&N�n��*��9�|�dQ��5����`���U�b�ʔ�	�I�W�UgNx��7;�p�(�J�䘵"|�3��>&���r��z�PC��</:���+[|����p0"�N�@�R�"�3rb�9&$v�J0f�@nF_��Z���sn�R���4h�;5~Ã���D�u�=`j$p�`���}�
�>~��_����Ҿ��2{U�7��>�V쪌61:ކlᣭH�F�C<�v����F�<��Y�x�p��ԩS�]AT:y�
�8��az�� ������K�gz��/s�紨�<X'�І�R���`�,���/c�z eDPa��}˘��1�<,z�ꮲ��c?[7������hZƅ�q
��e�����J�5|��`���K��^��o��!"�S��T����9W��o�/2�۹��n�i({W��>��C�Ԭ�Z8Nk�,�@�l� %�*�Poo�AX�3ގ��whTC�ؗ\Q���ΰ������np��:a) �0Y�wU9uZV:�����݄rT���R��
�Y�̩��)�mov,{��V\W���@�4�=�R7�F�UM��G�7��X�dHJ��ޑVSz7��ά&�q��䦘1"tSꫮu�T�{�#m��M,N�A{{Eb�|]�x��P3\��n�Q�g䴸�d�]���ϋJtv�F��WK��ϳT�E�;� �,����x��ђ������j��P�+�j.�9^uй4$�T+���Kz�[�z�l]�q@�3m?� �=��+*XF���.�ʃQP��)�cV��uh����dq�E�VنT���]�mv�/v9:�=�7�R��3r����m�|��	V�i������ wm�MaE�mșMgc[G�WJ��	&�
-(sݫ�^�H�`Nkp��8tV^6i�
�0�(�Z�jK���V6��U9�T������Mr}`�����-��Tɧ6�+T+8��{]��9��4�>-,4�j�v��\T�=���Y�ZJ�L�%�q�>t\�L!�{L9����ǃ����U6�z�����\�z){�X]��J�]�ZImg_9��C���r��v���B_Y��j���Q�V^�n�h�a\N�G9J���U�-Qkf���u�m�$�I$�I$�I&��U�	̜.�s�4S��q�oL�Eě��̽�H�������.RQ�ZyQ���h�xۂ�(����U�m+$�Æb���#�z� 8{ҧr���f��YlpK���WF��y�����$�?��W5���RY&��h��&�����r��nYV�WKwg�a�N4I��Z��N�o��G�]\�UNWf\�y�-nj��8.B/J�gV#�8�3w�ꆸ�H���N�*=E��^�n8��y��|�So!� ��4���uʆ�CPe����Ea���b4�B�f-RK6^�E�C�\2�.�Dڜ6R�6�M�tq~���|�+���+�͟C��8M�|r%�T���W���쒆M�:��NRP���}��^�ѝ��1zI��.�m��)VJ�V�U��L�Y��m�|z:v��	�s*Ě�����5s�h��]���b�J��a
[p��ɩ�Vh��a����0��[��co;fEF�׽j���eb�S�kA�7:i���Ol�*n����%{��U����]L�(A�OLƺ�zU�����j �z���������T����Z9�&U�ΎQ���#}p�.*��ɓ�ؓ�&��tޒv�#�.OT�G"O�RH~��hP��
�C��nV�hAQF�����{���"�g���3��|�=�E}Q�y1I��.ED�rw���#ܢW)'LQ�~}��v��c8E����W���E�d%nW�Y�AEU����Rd^��PO����3
��1p̢���!F�Qg�G�FOh�C��FTQ�f��7<<~�'�
��P�OMʤ](�*
+�A^xxTԠ��½$���¢*/�Ȣ�%R��<L�<ʤ�B�E��%�,�Y����	�Jj�zE�zDO��B�o�W�<�P^$\0���*=�~Ч9��DArS=R�r��'����12JT ��/SsP�WT��{S�)3�=LBL������Ј����_ᴚ�~heGd��[�h�gRW�+��ckV*�ص���̉V6�8+W�k#�F�L��Io��{Vk�u�wC��&�yP�ʖxN�T�E%"�,R����7¹�mrjc��0}����|8��P:xs���`����Z�~|x' �$3�ej׮RqK*��x�]G�������q�����6Q��,��	�~���v����u
=G��Q�a�>�i�<�[�㔽tn�\*�>нIrs;3yG`i��G#�#g�aC68I������M�bg���7��uż*D1Α��_�G�܀���88�פ�j��^=$@]Zy��˨�kչ�2�ᤩ�k�s��>OƮ���T4<zo�w�%W�\M��׽����6�h���ձ�Wlg��A����~�!b�B��~�J*~��̬�bs{���4{�/FUn]E�|/�R%�	�\�Pڙl�cd2J��)��;Ğ���2��U�Ϥ~ز�1�5�)x*�����~X?_P2�^��u�]�v�9���@��mb{�z�UoQ78�O����ݘ�񡦎��[�=cЕ��;���y�;�tW`��vrF�;ȏF����*e��>�ʒp;����%�+,���]�w���5B��cVf�Օ��.,c�K�f���r�^j�6�+�Wg��q�sU�9��"R�(׳��P�,�r�N��k��0�B:����U�f�v+j�)���" ��,�0:��H�i��+�6��D<��:a6i�W��F˼�=�Z`����=]wS	�Ֆ��=���3���3c�'��̫y�G�
c�Ey��K�}(�E�;T.����M�����F��q�iA�6gV%����rkbU\ť!�pD8�~����1Ҋ��R��R��Q��Ou7��o�d�@�����<$�o��#G¸VW|k�D0_)���AX�a�pUz���KӉ���pp���5C(G�z[�A"��,�7ZF�}�d��>��2�җ�X8xW��	X@���ΉX�8#�R������[/�{�o?xo�H�TE�$�{:����f�9;�PA9�ʪ�r:Xг-BY�%��7}e�`釂{�������X��H��)�;��$gT��;�����zV���e]���2f��wH&-��]2�̚�e���+��{X�u�&zX�����!F�1�`�&��j�#�Eӷ��,]
��J��l̸�^�n������yt�3	�A
��(!V)���[�Y^>��,��j�uo9�����:^���$g�/P枺J�����{�h��S�n�l��Ecy��MnaG
B�"lsw���ʝj`Έe�gd襷ΰ)3����͒u����~<�\)�ߗS��}C�&��t��%��N#�y�F�|���)�j�x[�o!��P5��"�͘�6 z���������"����h��t�i�
\�Ī�@�=�Oh�yV㻘����R��P:���D����T����H�<s��n��\���g�Iʸ��Љ�|��K�t����L4ߋ�~<J�L@�Km����M,l��$,H��Wh�)���PY�����%�-S����qT��.�<�z�s���1J"Ȉ���
w�\*���TG�D�:� �i�&j����b��Z�*�E+{^�N
�Зa�gkv�MоW�|�*���q�{���7ӧv4�+��I7b�r�5r[����-Ig���m�v���ML|5�5t�3��$	rX�v(�r�CSFE!��$ܦ�ah�o:��F;�x0�(�u�^��P�ƴeD��w]����*���i��#�?$� �"�����
�xX��a���%�A�؉R�ywSf��Y�v���� [�Q�*��C("�;��L���G����o+�oމي\��a&P�r���]m		`�����G�P�|Mf��.�����H6[M�y��۷Ƕ���W���ڂ�(d�o��� 
�`u΢���fgw�:��y+ޣV���a�ѣ�����i���'�i�����ṅ��7��ZeO{���*訄^�P̙�ɞ͸n�>���X��z���v۱���b��=��(�e�d�ێ�S��tȋ�(Y6y��nQgv%u�T,�yɺ;�R�>]Cf�!P�"+'s:d�<���� ��Ͳ��:�-w�;Z\��/{f|-�Y
�_����x���xR���x�{ޫ2<��y�L`��ݩW��3�����n�-v͌H*ŷm��J�Q�b�UvL�v�-]�G��Ys)f>��f��	R��9)#����m�s.h�⤰n)GM�b��Z>,���m-^��@ꯗ�ᵵ<�S�g�\ۇ�z�d��Xv�;l4���]ĎU��|�U�T*#(4w��y؎;�lt���6��Z_9q޹�5φ��+�qct�b�8�,��Q��D\�.J��U�5�u�t$z���Gw��X�t3��6��U�^���P�S�ϡ�Oa�Gt�`Ȉ��|U�c/��e��I4���Z5����ub�o�X�z�����èa&����:`h�s�� �=t�'��e3���hV���˪��YUo�B]u��)r�\o���?*O_It��s:t�Y�Y�Հ��V�0ljYzT��H\#J;��[����2��o��RsGƞ ���Y�C��}`��(��������.v�jm��5�?S�C���'�@��� ��<&��`E��U��U�~����s��E�D"��ۺ���m��~?h�R:��O�\͊dn��������XZ�~N�����KEW]}a����+���ݴ�N󻂄5�O8��M�E�N�b�*t�gR����Iw�׏w�7qW��Yτ͜���Ӛp̆w6v�-������2��x7r8��{�ͽ*~�A1�֬z�[U�`qyx`��+Բ�Ur乻�גc�ùr���9}ҬV%ZX*�E�E�U�|,T��c��<ur�<7hDdX��-m��a'�d�ID�x�4����C�k�R�UgE>7B���{]�|u����$���{������Y�՝6�S3n�1p+&B6*�L2Ϻz�ξ�>���!%�2�Ҋ��`RɣC����dkx�ڄ:�^{n6��,V*4�	��#C�o�D��z��2�H�RG�]� �󙹾D0��FP:=X�ySHV���R�(z��pЦG��ku�
���ڪ����U�G`26"xB*�P��Ap�u|�:%�=+)��s�˼%0C��!\�h�A�̸����i�(���)f��K"��5��Εҕ���(�F�g#د�Ϲ��[Yo4��,�v�ڝ{P)YׄL`�ijĦ�9�e�2�����2�K��y��o;���˵�v��'R��9\Ø�*(�%<�^j�J��"���R��b�#���b6���g8\�%7����y�������7'~W�}C���'��rcr�!@��8w��T�O
�>T��\*�5ר`4�S�	�ȜZ/o�(��(Y`���0�T��'����T��:ﴭ�ٛ3��r�Z4�MY���d�C �2��^��fJq`�N0�{&��@A��OG�qHq8`>V,ՊB�$���_������M�Ssy�h�Xܮ�]�޶7z���a�=]�x:�X�B�j�@B��\m�Ӈ�!���}Gm�ۇ��M���8����t��@s��A׸"X^��<M<8)������^z8ܛ��Y�����

C�ڢ&���W9�:����9���i<硋4�o,]���X�,���@߷%���.�qof�p����hL�`x3\�#~��͜�~�e�a���)end�X;��y\ʩ��)�|���f�(+n4)K5ef�6҅&މ��:%��
�4č9�,�~��� ǝ�B�������t���0k�����G�F�N%9V�:s�L_J���O90�r�S
��&_,�ӰN�7��;a�����V���x�94EY�.li�\��\���R�t�Z���x�ky7Gz��|9m6��C��/婎�J~�Y^ V� 9�G��/b+0�]��y�{����e��[3�P�PS�u����T�����7�ה%�	���e7�'���D1��M���;����%��**����m��Vؒ�Nz�ʧ�؁�f�
���q���=�������5�u�Ԏ���C5*z�Noj2��	E[�o��3&�!�y�A�T��`��̋��s�
�V�Bͧ�l~����<UC�Pf���,#!����G�č���Yy{����F1t�L�'���@���A(`���~�&��]'Q�mI�^��]K6,*%t7L\�z��u�oO���ϑ�0)G���$�wӗ�K�<@��율/��W���,�I�ˈ�!�[�2/"�)��sk���`��M�2�:������^@r��AUw/ )�����	����c� ܔ���G]�8#���`���/F�Rm��%g4��M��!l�~��GUܷ��d�=0���w�������of�5�r|�ќ�-A������ gS�	כ����U�p�TJ{��AZ2��jK>������qQ�1��2�����x�e��I*}���,���~���\#gFU�v}��-�}�>#�-��[~u�X�xVjR��F8w�_l��81:ރo����9��Ƿn�U(轗��+����N�HW����;��pfsZ ���h��fǵ)����^L�*e*��<=嘆
��r���)$L>�w���n�T{d�1Ǐ5Z�nxC8e_Ps�yCO�$b>KW���P���4c��y�����	o�]�#%{o�IY�Lp�2����
Έ��QV5J�}	�~&1:'���u�������p���ׯ�Fוո��:_�Y��6������i��h���`@~����F�5�C�J�(�q��
z��F��L�W�8E�]����s��Y������L Y(<�Q4��]K:t��jM"�T�7��[W���U�:a�WJ��J��A�t4���/6�0XCÝ5d����ތ����q{�ZP��kF�_�qn�������}bC�Ǖ�����1�I���>�61%�i��跔wspoE	q4-r邒����(�M�o��VH@�2^�T\:;��/�;/z@5�X�����7f"��R�C��B���K�q9]F]GI_.^��P�����yhW�L���q�D�b"�N��E�!�2 %K0�����F��ÈL#�N8�����)��B:�^�;lC*�3�#e���l��J,�u^T����il��>��Z��%�x�j.�j�Ϧ�G΋=C��=�	�a=����v[u���;�����9��X!,fUypT���_cu���ߢ��tײ��~�X3y$���'�Y)�s�%�E1�֬KJ�_�>��½G�>��1�D ������&9V�6�c��zf�����e6eǄ����@��`�UM���.���`)I�tQu�J�j�y��O4]�U�Y��"�{"2C�Ѭ��mbՒ����0llp��>.�|S���cC�3�w���Q��h�e_v��]ͷwLz�Ã�)H��xީQ�,��:E��>�k����R��)trRlcTr݌���t�X�̫��Q���J�*|��A�ul�B-_<�7�t�+x��������,��hl��ʂ�C�Z֫̕�R�|��w�SR�&��6᫚�����:��$k��~��1:fj7}P=m���䩿K�X����}��B2[Ӌ9V���CX�]�M�����=ր�6��p}�,����[/��
�t3]^
�38��a���h���/x�8w�O������/{�Z�b"gJ��>|qɷ|.�u���5�q��'�������.���;�e�_e���9|C�0I�ZIi*2R={-Gv���p�7�r|���i�1Ms4w�+Ch"��*TnV��+��W��Z���HH��k�b��y˗p|*�K̡G���m���ٍ�s��;C F��R�r���_[q�I:���x��%�i�M}-ڋ��H����g(�Y��Oc��0@�u�Ks�����☯�^��ic�p����d�Vl�t����S[�Ь�{ȅu�	vU�ꃍ*c�ص+t:N�E�,�Ћ���=���M�G��_:Xwo�qAA��5{lJ&����u����T{�2�v��N%7�̎�N�ܛѳ��C���ҎI$�I$�I$�cPr˙��C���R`7I����ו�vT� �n���:��=4��K����(��km�.W��uí���*=�P%�x�$�^�����S�O���)�vY���v����2l��Lvl6s�Kj�4"ڸH}��b�7b�IGw.fJ�xz榶�m����@7�k1I;p�Qk�=Zĺ�@�t�t)�ˇU��a�i��,T�7b�p���5�LC�+Ln�tj�
@2\B�X�Lɂ��;��M�<�i@b\�WE`��77n�d��5�f�J�^�+XB;鷊�mª��a��Uu�]IF��+�Ab���n��6���Z���>�l����){g.���b���@����*�^onNZ,E��{�(���S]{p+m�#	��pE�h�N�8�$�lT�}NT�+,��E@a_i]����:�S�椅��������&�}tu�<�r�Y��HmvӁ�V�d�v4m��|y�}�
N��#��gE��LE�|5\I�4��Nv_��툡��d�-v���7��:8@�^��u)�;fMt�M��tMƓMI:�I;���,jF�S��t��U@j?p��_P��J<���"��:x~��e��*d^�$��dD^�Qh���xyJ��p��}��
��A/<�M����*������#�Y���J[�{#�̬�B/�L�^�O�z����/޻$'*�,�"�1=q9��0Kt�t�fى^ԟ2��)�I�!&��A�w�rg�UJ��=��ye��.g�ʆ��i��xFE�L�xP��7z�aBT�+Ցb���?���G��
�+_��χ��o緄G���r�9y՟$�	�D��#�R�Q�a�w�i��H|ｦ5<���J�B�ԕ$#��Šf#�J)��Z\�YR�d��KFE?k*�n�*�Jhc�o�g+ٷ�ι/��<�Z��H�6�����-��1=N�c���o/��C:�o�Fn�yWz��jT]��a})��5\�������V�T��&I��������a#N|�Ӓ~��k��%�蟷WÆY�Q!
ܕt�|�_�P���duN��;�Ԥ������]�t5Ć��bD0K�,DW��B�:SC�tk����0�M������c�I�<0Q|.��B	C(x�������*D��X>���×"X���9�A�X����;P��ۙq�$#M�J*"�
Y��X	x�8[]M��&Qc\�"$٩S�X鲎%5�T�L��"�W�p��y����:]����5-�0?/>������0z%^񐡔���ϝ6��*��ҷ�bqE�"�����S��<.������
/�U��ᇼ��/z��ӹ��{�=Y�X)H�5������F�Ɖ �&=�]��K�ԓw]Kȹ�N:,��<��/��$X"MN�3J닸�cwn��KU[��jk(+����P��dCQU{�!u����֕^B��g��x�ŉN�*�7��`.�[X�����eJs0�Θ�a��.u���ܛ���1�F�W-���,:���X��'[˙��;;�R�3��Lmg2��E�fB���弖}�{�9�����ٺ�أ��h�����ʢ&����{}�:�L�D2�d2'��ъ��h��2�N���P67%�].��
6y-�3~n�w7��u'?^"_��S̠4z�>(b8.s,Z�x�EE�,�qe�!����#6���N�VR0��������q�5I�u��u
�jxB�Ǹ��2����*�럱�)��;G��#�b���wcJ�0N�"8��ؑN	��sL��;ֲt��O&	�H��=����P�*]K�h�FZ��؃}w�(�y�B�E�����+=���!�S���Y?&�|;T��91P�T4���p���f���O�iG),ΰ��f{.��-�jy8଒�̀О�ׇ)$�r�O-��*�@!���������y�_�{_uҾ��p��{�H�b�%��y�NU��P�: }�O�6<��r�A�r���-��k��[Ѕ�z{��ʀ۽yg�ln��ʺ�^p��f�wDl�M�*��r]�c{u��&t�x�@W��e�[C~�[i'�(��z�������8^r���lv1��_tp�@���y�&��9_�۬6�C��ԗ~-�|�atŉ�̓�ܙ�s�,�gҊ&��@ ?�`U(���\�
�#h�n�.�bbB#hU`�J^�˖`�L�����X"���h`c=gۯث�M&�.Gb6eEr�b��j`����WQ�U�^�O{�֯���Z|�.�&��4B�����u����^�돀���]O 
����f��)^�o���YHp!q�5~��?P�6�h��e;5~Ã��D�փ�#X}�9Z���Lkvt���3�~UD�X�Ђx�|kG�qs(1��xE5{����so\�4�7M �"�y;p�T�Erȯ\�B�$ k#O0Ӧ��;X%	3� ~����Iѳ����S��Yoʠ�U�t���İ!�[*�Ϸ��$+=�I��V+�3x�V<!�3���
�Q�؟#��Z����h���m�� �Cӗ���+��<*��h]+��|���HH�Yt��釀�/x☪��11���p���	b�O�>�T�2�HT8�m%��Z��P���m�Q5�)��z5ɬה����(�GrƷ�|����t(P�k;�:��]�oU�S����#���I;��Ss5���.bA�c:�E�{��n�qA�/ج���`�yWB�������wT�P�(*㊺��L|�K�\Q�Sn5��������b����������S�_�u�P�U�;A|O��w���54˰�4ǆ).f^ٞa_[�[�_1V�`�1tP��.bt5L���=CI��Í��ꁄ<:����^D��6��Wǋ;JCJ�I�J]ĉWP�B	R�&�_�ÿg��pHs���9���Ʌ�s�Gޔ|K�8X�DX�	:� C�B +'�=q~y�3��~�������85�G�����`�*Y�l8Ij���Ҳ]O<�i݋���&�_�p�,VR"�ȥ2å �*X(�����Y/9��ۢ�G���h�����+��?�oƕtJ�0;=Zhx��E���-�O�g�&�X�P�-��s��H"�`���n��K�T^^������<е��\��qz ��������׻>q(��Yu�6\Et�^������0gL�i�B���y����ԹI��v�w�vmi��928�������!B��m�RVC&ʛg6�W6�y�J���N�(D��<��2���K��I$���XE��G~���k�4
Q�����E�1��3HC�@B'kfZ�J�f��:B�C$϶(��X�]Oz_F�+�Ժ>`�xa�|�����~zh�|��͆\Fl2��{^S9���㚥��t�n
êˌ޷��R�F��br�#�0�#gԩ�7ᶩD_C6�H�UX}�f�v�n�G]����ƭ���Sk���g�Q�(VJ4��i�c�hb�m�t�Zb&jvS�݋�K�Ln���-L���#��BDh%�,`$i�Oi��:sHS��r=��F�j�mӓK4�z F���`9�"�9H�B�U.���pxl��ɠ�wr'�~���wc��Yx�<k��W1~P:�q��\E�
|��GJ*"�i.E��嶹�w2�N10�(��(0�P{�c��'���h�T��N>J��X�������`׮5����U/��>��<�����s����"=5L2Z ��{4?�U�p���MĈ��wc���c&�eV���]��P�t��t�0�	l�\�o�,�q�nugu�N�ҽ=�dQ��A��M�����{������*WZ���w� !|*�y.��׏��Ԭ�A����N��O
u�c�t,R_{ΰ�^C!�kz%�ԑ�sgV�LjP�H�"ܾ� �Q! {+T*��Ÿ�2��۝��W�N���59�{j!�o���n��fp�P�Y�>Xg�PB�R}�>�$������9ϝwv��Ū�1������1�mԣbi#��/�)�FY�Xb�\�XsLT�\="KT��rh��e�9Hr�49S���ʝL!�{��Y�8�u�l��<)U��/�+���6��c��W�H���]�fs�qN���s�<�b�~�eXޣP{U�;H�W�υbim
Bx�)�Ï[κ��ԟn�s۞b�8�L����<
7�sv���.#tG3F8ZT��Rl^;Ļ�9�h�WK�K#��t+��ר�/婎�`���*O�
ڽ�1evT�����;ڋ'�
��V�'�T,S�L���<%;� ����p�g�;2����t�K�v��eFK4�wI��h9�&CX/fGu�m݋���u_�L!ٱ�x�5U�Ĥh��y�33��K����/8�q�nE:<�::�I�R�^Ɏ''~|"�����ݖ�M,���]T�
��Ⱥ
�n�AG���CHTʺ�@�S>��^2��/�|����o���R���ේ� �*�=7B���y[����a�G�a�t�b�"�ҍ��E�P�tb��3�	�bze,�W��I�ͽ���;�ӱB���4����N_;	�Py�&�fI�n�B�r�����'Zd_��1Aɘ�}GIH��@�>P:�j9f��+{]�z�Vb6�P؅.Y�uX Խ��|�u�K����`"��@��>H��t�+��yDW#�,�t�tTl�ue���#�NU��zO0�ҫb*v��sQ�f�"iW���f��$�TU�ܼ ���2����ޮt֕�%n�J���pȘw��e\�Q²χi��c�#W�8:��D��>��%绸\ܔ�����Dj�C�ʮePdPͪ�o#;�e��(����k�-��S�-N��H]	)�طV�Aՠ�ۢ�dko��S��6����t�^���9%��c��L�Ԃ��$vR̒f����R������U��2���6��
�X�r�7�f�K��+�m�w{�TQ�o:ބ��<�FE�g�:�mN��tȫ�(P�#�u�u�t���>J��$�/�/bO8F�z�61wP�r,��$Ed�o�����V{ݲ����:sI({�3q��x�8�c��p�
����yCn����g���d�f�I=�˵[C���u�x��X�@a� `���t�;��7>@�Q�8��K�th��)�_O�*!�8�ƹfͽ�!ŌA�/ج͸G����ط��_4�!P� �5�ʥ�E����_��X���(��Mye;��)l]�)3����(p��� < d莎�P5���`�ӹ�l�2)i��5Tr{p�P�~�pi\�V��Rʿs�!����$���}`"ǵ��wsN�F�=��e B?*{��!o�fʫ�\OP�}G�J_���:ER$�jh�~�NzZ�2�Q�r���^�P�V�",Fy�d2�/%�|�'�B�~��lGM(s�k�!R���G��=]��,s{Bӣc�=ߖ��珅
��O8��n�[M��/u]�W���DFL"��*c�4lb�s3Wf����:�v��Z��H����!�j'$_{���p�Eɣ�Q1�'#��9���Q���&	~C° ��y;���-̮����,V5]Bx9&���E(�d������|2����-/�����ԴG�`��W
��x���Gw^
G���ۣB�O9�����l?'�A|;7�H"��QbbV9ױ��x��4�{�;�$��Ėv�Yu���(�8W�E�]��V/,C�������~!� �+.A���e=�j̡��Y��5����)������Ѧ��*�,��"|;���E�*8�14�M_K�͔\F�2�Ϙה�`n�鰵S3YS;������MiGIcDM��ꡦ��ڊ(�:g��^��g^�-���H͔!�+�'s�	��K�4�0:E!�"i	kǙ���t�{�m��up#��64��r�r�P��=.�;�u�1��(�k�M!ZЪWw��8(�/�#�q�B��U��Ҭ&Q��2��X�!��:�����[R�9Y���,�J�&®�<�����ɳ���v]�s���.�ȵ����l�YO��T�7u���3��.R飬\�}�7#���o9�A��* ș��!0Q��NT��*�f�\W��	��F��H����/e�b��&��r�����w�}�(�([(��X���sD���f��謢lh,��cP棐�4U~��F%roN��c��v�s'�%����Y�S��3�]Ld3`������nQ'yê#o;�&�������{������<<*uK����P����u�B3�L��}Rg$0{㜥T;�����AT)�@y}�3�O�=�3�y7�ϗMn�P��g!!�^x=�l"xx,J,R���WJ�lA��ݝ�HG��1=>ȩu\@���t�w?h7^�p������p���ѻ�)�>���Ō�fw� [4Xز��7�"�K�Z�ݩ�50v3��Ӵ�C�W;#�����sD���a��z�Y@߷%
l�]N���p���d�YČ�u���9��Z�yn�>{�Z��k{w�}���N�w���HV1�w*7ѡ�A�]�v\���F7xU:ѵ��YZ:w7�P �v OY��fl�Ղd!,����Ʋ���μ#\Z��
3�2�R����2i�eY���>����W{,󚴴�'�L��Tj0�v&����&���z8��}w4��	�/�m�6Rq ��Z�w�TƐT�܏)�8���u��Z��\�5c4�O|b2�=�S;�m��f�[V*��tT�5d���o�J�9z������(��ӤY�e�t&����Z5}o�xo4T\9e�3�T�ݷ�a�7&�0��s$�w��I�7ҔFb��[׼�$�c*�4:��t�����ncP�g�>R�=96�ӯ�-�N����I�L씳t)�#�xyb���vW֍�*����aJLӖ�sn�[O�΀����2e	r`��VJj�G[!�o�x��OY�BT[����L��Ο�>{�a�@�7[s�E켘m���g�ȦV�6q�d�m�P�w9�3�,���^Q�CrI�JU�|ms{D+D�Y�5��6�E���s!�(�SB4hR�����[oT�[]��ć�S}����9ⵜ�"�O�d����;u����ZU<5�ql��-�$�I$�I$�I���`����h����p���s�]8�K�'[��f++�X��f�4bV�V��k-= �?
*:�LN���GK?l��Oj�M��M��������t���޻Kʗ�ܸo��m�,�GQY�5��T��tX-���zp)b[t��,ͧM�c��pi+v9ZoEcb�@#r*��ax���C!�d���`Zs*a
��+s6���1^�b��`���]m��hRTxQ��q@�e�\Ѷ����VF=:B�Z�R<�t7�űB��/�p��<�z�H˻?kU���!����5e�T����#Ǽ<�aN�����7�C%:ЩPˎ�䬆��Ds��0��E�t�cJ�,�[ic����n+q3�>�4=��vheճnj�ա�v�U#�I�"�>;DY`U:�����FW�B��"�=��39<��Gy�a=��Ό#Y�]ß]g[�b$�D�K��+ �}���>�[b�+ϒ�2��Fu]���K��r�-q����Y���{e�7�H�$8n<��ɸ�M�������ӖH��ͩ�����yU!z)'(�,�^�ܹ5T3kfK�b�>vؓ=ޣz$�>����m�{\*<oC�J�^}e�}��3�y2�y.O=?}d��B���$Y1-jm���+0*BK`�P�_�=	ht"�z7��Pu"�:<>�5��{G��`�n���g�V���*�罵�ϑ-t�ȼO�W��b��u*�m	��޻��������$'�ۯ��_&� QyW�z��s�D�J3f�HE���������*��y5O:�ϴ�<z��Bk��y�|�ܢ򬄧���w��Kː�CR��ut��'�AԢ�OB�{��U^�2�ۍ�{��HE����`�ԫ	��]<���n	.IæW1//������efX�IҮ颀8wC��Ы153 D*Z&�_
( �#wR]�3�����<���ڰy����H�X�ϋGh��,�l��M�f�5�#SK���{[fǪ�+����N!
������4.#hd�0u���x�4����a�PA^��.>�t���i�E�ʝ�(_��h[3��v�7�b^��E.�nh5�����k��o��J�Z�?�����M��x"�^��xN�`C���/.%� uq1멬�Bq��Dᎋfv"�!s��&mݶ\������g����\���j�&2� i����|$-z��AN>�j��+[��8h{>U��Цqz8��.���E�T�m+�j}�[J�v�{Yv#>��aU�*�>"�J U�4M<��|�����з3���i������1�'Ƨ��hk��]5ˁ��uNY�5Q�G��Z���^�vye�����5Z�lEuJ!�3`�R�&�*f ��4��q`�E;Y��,#�����L����z��s��n�L&�h��9�g�����*�u��˫�P�ok�<�\�ʼڕ�1а�`0��A�K�ظZ���&�%���|U����*����L�[2B�Rup^e���3�T�s�2��o%�{Z���}�Y܆�?Q�����	�291a߁N�~E�`�u���|%֖�{8s/n'ꚍ�&E��r"�E�%����$�JI}�iK$��1��t��[��z���ZI�V�u�V��v]{ʘ�������+N�5~<'�|��լI98&�2}[���m��dU�4�	U��Q�J���j��>am��SmڋW�-7�>�b�Ps<�>,@Ǵ�(��x˸���#}r�z{
�˭���9u:8�o�)�Qg��Y��wP�r,�X$EK��),WL�lf'����~�L%!è�qę��8��9���͕[!�u\����L��u�+':����i��B}~��<N
��o��G�+O]pn��I�l����^%"�&$H� �,�͊�:j�D#��6�-@�z��O��g��g1�����]��|H�4�:��}���m�=^�_��E�X2S�e?E��q�r�`�0�]�4����V�a��.x������V�z�<9wݸ��|�T���5���\n��ٱ�����ʭ���1�
��y����j�W�gJ貚�朗�6Cz��ԗ|^��o���5ٱ�S�߅PP�U�>���=@F�z|!ӱʍƻg�YY�ݯ�7���Pj�����Q:�`��1~�������5�*�˓�x�����D[x$|-��������6�&gޙP�B	C��N�?5��m�c8�^���Qc�h�r��ˇ�F{���\���)-�u�&�*�|-��p�S%���F���'�!�B�'i�3`��`��sl'�>�洭Љ,wN��h�ZC�P�����G��B>�$���;Pi�*{���ΊNq���}Ψ�DpkX,[�S���s!������)�]Y�HVU^r6�T!U��A���_��'��!>�ln	�)�0�=�J�kq
{7K|v�tC �lym��Z!'<l+�7Qo���X��<1.#vuC���������,&�ʞ9��6C$��jUb��͜���5�mO>��׸����2��z���u��Zo���T%ViV�1ň��[t�ӕ�~q|�w|�5�0"�gj��B��1>:sx#J���lL.�R�Ιܜ��d������D;&:곩Q��7$�IO.N��F��~�*�;6���_�L<<6�j�q�|}�镁���,m��
Z���c�)��Q`[Ei��W��A	B�|��h��Ľ���<=�D�[���y�*�0����Y�1(D"��#���u�D��Q����/�r�o^�*\�da4���>��]��V%^T��]3݃��9���*�b�Y����A�0o%�����]Vт�@3�f�Ѷ}����~a=��^�|n���lz���DE���B�5�@*�o5�+Z9=*�,q<]���*�z(4m�bm;�WZ��3�*F���I ��s��w���^��O�i�.Y��4.0�Kf6(�}2�q��R����K}��.��=�&1�hwƈ�j����a��ibq�ؿM\%�]<�����E�i��A ���w��?�iP�,B@��+Z��ȱu<���MnG�-��/��'%�O���XU��a�5�.���K�K\%;J��:�AɻS��6f0�zof�܏,m�g�j��4f�9����jpP�,��%R��>.ԕ��g0s�nE��������O�B,��Y&w��/9��w��-Z�geN�*�B��z�6[g��V�A��a���H�bCJ^j"�N�f�2�=�{�bL�h3��;�S��K񺘨�8Ybԇ)u�~N� SS�2D�Ƨw�~i��]���ø�G��ɕ�s<��=�(��uf�<l�s�������R*�@�0�(Z>��J���J���U2�x�x\yo2�d�w�9�E�Hh�oڅr8�de�4^>UR&E1CM�P����W9��r���=�[
�x�C��dYЯ�9�v4�OU���c�^b���F'�-w��8@���>�B�*��mR��w��#(H�5�-�u=�yL�cx���������?.%�����\v=m	�D��`<n�-'�=}k^jO� W�E�� EN\#�zxժ�a�/��+8���Gjy8Ҟ�� ��h����M
hHђ>ژ�R�i��η ���V�{t�u5�;���&���v���ym�.���Lu%�U���lU��+��X7����2넧�s�ᢤ«��M���3�j�gu%��^.M��S1�`��:DyР7��s�Qx�?��т�z��:��`�q�u��+V���(�Es�3�œ�(S�Q�A�k���_� vS^M�k7�J�X����(��5�J�����*^^�@x*�:J�UQ��KG3�����8�� ���{+��YpR�y��8���%u]�^����M|�I�zzy��+ȀG�<˫ OE7 ��ŇeȰi��W����#q���U�T-��A�4_�/���96���cʢ�PU]��
�a��i�Y������)�7>���l:��j���L�����������J���ӵ)�'5�M�X|!*�n�*���dVC�j\<oά�𭴥X,�z�>��*��Q����l��8��f��(>�f�B3�;qs][�DM,��s5��<cT��@lׇP�(����-ˣ޺b�Q�J\���s[7xt�x��M�;w���S�9����.�����陗��R�kY�>�z�eq�(�w����rA�!	���o���lN��Q�f)�\dY8pTz�x�T�-Զ�yf^�.:��$�����H�>���R���ɖ�ذ�b)O�,����Ɛ�9��W�ƫ�5q�-����"6b��.x��P:�/���g�i�qhU�߆����Pj�)��ΣV�A}B�mȑg��4&3��i�_K�F�ӦYfKp�'�ͤ�;ެ��bk^yfW&�� ` x��\��s��k�qU+�k�t�,��NJ��j�}C[u�^��9�Gh"| D��?%��z���y��Đ�ʞjȫ�s�>T��:��y�����}
YQs)��̳-�s�'�73�p��
�����
�{��B}���L�NJ0*�Н�E<���$O���Z��w@�iQb
��Pc����p8PȀ|�[�͇j�oy_rI����������ʔ�|,^_X�]C8b};L����n��w���λ��=����q.���b�O��TS��..�GƾG�~O�Fo9�9Q�{�h�|0�8�j}!��KC���'�]��A�r��w�wρ���5�k�^Lk3z��o�`ks3`�f�q2�m%dg�;��8���_^��g2�aѦ���%�R�\5%S=�as/8������b�@��RG��}A.���=��0m���P�tY��2�kX,[�(���]a�����-qu7y�0X���u&�f���m�D���+c]��&yP�TLMĽ�8��_���`lKC"�b�|��Պ���-��ʌ�'D"�&FK}��=q	�
�'[8^T���y!�D�c����+��D�Ž�_q&���pV~^,U���������<,oK.-ף�S86[҄����Y�R��T8`>�{8z��G��Vl �WmIgMgK��Rˉ�1ݓG:�I���$�?U߇�[�@�yx[�X��4�AB �HH���ȱ�$�B�Z��ou-LDPɴ�v�z;@�!a�D�Ԫ�6�>�R2[������Ϩ}���ib���f3 ��i=A�tU=�+���z,Y��=w��2P�C��/������5���ë��WC�^�WJ���R���&յ9�ml|Μ5��Jz�Lj"feKiշKF��*Q'�vm�-�lRT_]��W�uN仡�tr��XulH�̊K�%��Z�A����`i��0�����@cF�n�U�Yϲī����%���������G�L
�ZlOK7`�f���T=�U�<��;�(������i�4]9�U�t�*-B���>>H�p�B�zC�!T읬�M���^��n�q���t0w���r���`�{ ��+2�M��s��(ٓrX�4� Muz] ���!=�7��Ƀ���|%*��T\N���q�~GWZ��:`ʷ�$��D��D{u1b�P�q,؞�%B�=�禜��C`a�H��E�)G\Iz6p��-�"h��m8ʾ���l�u�\�	L!s!�>�R+�K79,�;�˥!�+��|�guwR�5*t�ɣ4���G��ڟ��8˳�J�R�?���>[�~Q�����yl�U�^w^2���*#���U��	�Ƹ{R&E1CJru��M���q#NT��z~r��ӯ"�}�w���'�]0͑b�nߍQy��S=� ���z4�|�7`��,lr{ ���A�T�j�y���K͸�`1-Q���m�O���v��'o+��Y���qvSI<�����Es> w[�}�\..{^��A�[;4]�o2��գ7��:����%�
�? +]�u����V���Ի*��]2\x��^�]|���|r��wpxl0/��	��X�ly��Ǖ :cb�l���9z��w:��~�D���gC����W��ʲ�1J&�&�*�Q���66�V�@~<�f� |j*?]
4L� o�U��~W�ጡ2�G�ދ�3
���fJ��-���9���
y
� R�&�ɯ7T<�-+�S����z{.�l��!T��Glҁa�w�):�"��1A�,�v"�;}�AZ�&����8���l�
D�g(\�T���uJ!��u��=D�*}�	|��=�N��mӱ��$A%�8e�U�In,891a�R,�XAyǶ���R(J��Ԩ�0�)"���%������0_ԫ�M�����}W ��je����+�|^�V��Yu.n�&��b3)��+>t6�d����)α�o�i����c&�w\Xŗ����R��N���P�Ԓ:��1��-��7�v�/e3ϻ����rfn:B��Z��C�ҚH��ʣ:ț{mTyo��rS���e+�q(杤���(ZX�a��t�a�����%g=5���r��ڇx�m�MW.���e�Aw�w<�OS���U�X����6��#}�Q���\�B�I�q�ǻ0�4�Ӂ3@�YV�c�R�,��h�En]����g�ͥlM�E�WԻ�5��D�L�)T��$�1��}]�f��g��`��X/m�Z)��oE��[����u�D Rk�qn[D�Ca�Ʒ� ��A9Uص�rfA�I�+�wJ���b*q�5zA��<�\��Me�ܮcViS��E@V>����9��%>`�l �3��I3.�ӵ��V��|&o���/r]E�+j\9Ju�"�˃�S���tB�u���c�3f���}�2��)��T�ՙaC|O#/�%�ֶ,7���ъ<mr�];��+-w*kj�d��yn.�b[��S����<\n�#3����=�[���1�\�Ӕ�%��q��pu���!��P`'��zu8����Af��V���I$�I$�I$�d��Wn�8�S�&ʑT�k�<Xz���r,�}�Yu��9�*p��������a}{�8��ږ�cW�)��6åښs�^Y�ތo.q+mZp�ڛ�{���B��e�z���I%\L���˜���y:��)&gׅЬ��4+fm�J�,k��͆��H�GN��`PxF�(�]	w���ɵ+vc���	l5��$�e���5Y��� �tY��O��4�Cf���NF�(��E�Y�a���K���n��,LE��_LT{��T�ڤX#Q��p�ڥ#,QS)���qq�k���a|k;�ﺝ��n�4�FFӵ�.�=W�|�� 7�+!T��1a+��2K4���x�\���4a:4�����rp"���+���3�B)n�L���g�ܵCy��9�V�R�T(�n�Tt�zdc���O#2�9�M?=B��ɓ�Gb�eA���*®��V���{�����{Cr���3��-�˒<78c�U�:,Ն
�s'1�����]#��jD�'2$�rk�H�q�ݽ��΍�J��h(��
C��cBE������{�>|�ȝ2���2��v�h_�Q1�i�Q*�FIz�$/R�h��vM�\��#�Z����\�Y�h�����Ţc��].�~����o����]����O��χ>�"״=��W�Y�ڱ9�싕2?1E�K��1bT�B�D�IQ��R�/=����\_7o���P�$�����E;	�)�E2ɤQOy�����F�Tͣ'Z�#�z�ｏ��!�>����AE�����u���}���B�l����l�Z�Z��{���|"x�Ʈ�W���2o�'��J+�EEqB��������½��gk�3ܢ��N���D_��E*�z��N*Um�75
/�+����E��5s*�0�g�E3���b��$��">x^�����PSжe����^�Rѹu߉>��<�ȳ
���މ�����= L�2Ҋ&��~��$�����ɿƼ�	V���ށ�t	�j����.�X�� :�;X�"Qc���C7��7hݝVP�F�u%ߞ��)��lfˌ_� V�u��^�G�]�^^b��E�3f�(w�6��//-��K�������Iu���T�ȫ]8z�Q����T
bX(+��T=K��5v<p�	��c�qs(9�Z<a	^ۦT���e�.���^��}��Q�B���� 0f��-�֧�ȵ�B
!`�!P.eU3v�t�w�1�2���~����H�����4f�(,�c��55�]��IDX~R:�iZPګ�P:�/��~&��!c�W��stj�#J���mdSd���Wj�y�*�T��D��G<]�N��q��,��;��N-�g^�wpn�x1޿b��`�(@��*4�CA��V����W��dH]��=���*����"=����*��Ί���d#A�,�O�r��Z�����J���5�X�.��Z�1�����<�||/�PF|���f�_���7��?e.����!��s�GI&��o�r�A�o@�8r�c%kAp>/[]뇼�q�q�2l����\{4,5�ԗ��������W��n��p��g`k���,�a�A��H-&�!j�"������O4�i�}�t�f>ޠ�bTB��2��jK?<�zš���}����`���}��/�ƒÅPy�)�ܕX_.�*�*�r!�a`x����Ϲ	tl�T�p�t�Aw@����F��9�DW2�8<�]"X���pK�
4=Q�9@׶���_#�ߕ*x�>va��g�#���V�N_�?M�T����pu
c �\��][P�맷c��G^>�iq�*iv7	~�zI���DQ��x���>U�R�=�k@]֨��>����I�i�k�Ll3�P��u1RBqq��2�ӆ�Po�o�!=Ӛݥ.5����zϩ;��]H���~����)��W'[�)�"/�/��D_:�M��=���h��f*���N������u��
���M
%��d����Ijm�j��s�Dq�q�Q눺��N	�E�͍Rˋu�����N��-U�;U�m*����q�)�����A�dvz�9� �԰�%�����-P��xtfH��j^B��ؙ��s��4�I��DsZth���ޢl��y�ٟ&��-�$��n���w�e�\�8����[�w�� �rԵӣ����J*���4���^X��T$n�<pН�B.c��B|����ݬ�]�"f���nv"mJ8Բ8)�G�Ɔ�#7�t\q��}�s��k1��c��^�W�,T��H�^���'V`~74*UC����K
����<�����k=�٣Ϛ�t4�=O��졣�A/�p�.��W��*����b5��ִ�N�qߍye,���$q�߯����v��(J�v�M�;��U��Z��U�]�p}G�xW��0j-�I�*?~^0xJ���:3S߸����*ob��-��Wƻ�y`U)��.�](�5#��<�W���ͷ��5E��3�KcG���>8���>JPc�`��x�#��c?��M���й=��⃞Z� &�ƀ�=J���P_{�ಯ��B���X�y��a��E8T��0k*E�r�<�&X�
	��	9���x�%7)z^����}�g=��>믆�Oܢ�-���<��L��h�/�}2�W�NԺ��&�hNYc,5A0�v\�Y�M���]9^�ɀk{j��{AK�Վ��e��.�l�P���F��Ν��m������|��/y�"p0~VM[.���5�ǆ�S���zIY�m��.����f����ք���dk�W�a�ug��S���y��B���+֣&�g�������0{��y�U�@��-x�8���
�e
N\>9E}�5%���{� �Ǖr��炻�^��i�p�4�@���i�SV�m��$p��.;�Q㣧�;ծ��3�}A��]��r�¶��E��]��v�}V� R�2�׵�
A|rc�VŅ�h����hs'2(OM[WlA�o��\&j��Cc�,�ň�������f<|���ͲɄ���)Q��;g�Z�������xpB�����]Y
Oj/���w1����в+��՘�`��]K���(�L�8Jg+VW��2�z]V�L>Y����E�!��Y��~��&�����8.��q�C��wn]��7�m��Pǜ��0��LXo�#���u�s�/�Y�vߪJ�V s�(�Y~C.*���2.�M޽xv���a-����b�g�ݔ�\�ó��Yu���b��uҝ)E�#��%+�.7����;6�o%�����7����#t��S�@�tҀ�UmGlՙ�,ć$��Q���Fi�ޚռ�.gD~��L�D�"ʸ�*FDl�!7U��"D�f��8����Ԯ��h��>c�T������")X�v@�.��d]�u�����if�
V{-w��ӄI� �Q>uk��Q�>�J�/��I�.`�|o좇�ιu������n���W �Rh9QS��i���*UL��L77UUm�xr�|�)���������,xY*��X^�F}ֈ���B_�b��l����w3U#A�<z��1�U�����Z<a	^�!�
8;gn.cYngR�j6*f9gM��(f�@�	��NJ��\�h��B��/���ˆfsKD�P/K�.а�]����C;xHH�������F�l.>{<�q�.B�j��eB�^�V�V�����Kc�k3��u��"k�熆�.�7x��?o-�]kP�1M����6�}��,K�v�+RT�S�-�&�{�w<�	�(�-��X�H.��r�7����L$M��\s��'�m@�qye���5j�!�:v9%9�d�-s�j�@��%G�$���ꪘ��ѱګ.�úY�5)s:!"F����Ѝ;}.!�,�ݥQ�+j�r}�d��ly�z�a�_Y�����` �
>Q.hh��s���[��^cP�p�
GԽt��)�<����_��p�P�F/ <B�d�����.#��V�w�qX�.���HDDE���'s��3���s�&����S�u*T��X���@i���F�q��J�I�SF0di�UW�z�n�R�d��ŋTQ%�:�ln�P^4@�Y��K��|�~lVMÚ��9�܃����(�����RU���>G���	�C�}(� �|K`�>ٻ�0K^ÔC����x]EV�Xj<U9to�삭n�IE�?gn:�^����Lq@�P�a�ۊ�1bC" W0Y��<j"�� �s�^��\<6�>u{nd3�:Aq����8Ȇ�Y�|�"��ԝ�nS��`zu5��aTM!���n���}��k����+�ל����{+{�g�ʀ�����5��-9.L"��=�f5p"��Y�w�}\d��ے���ׯ��6^��g�sbX�6C��n$[�ޒ�3G��վylR�lq�N����0,��K<3���u��K�j��-鞭֕�JX�<nb��k�e_�?"o޸2�kh`��p�x�##�9���Ow��D���φ��v��z��GR��u
�����u�T�����5ݭr�����*Ԣ��X/ޏGo/޺u��C��O��ԏT��H�N�ݵ*��f�t�D_C6ܢ:6Q^�T��et\i�Y����=��b͚2�v�ͻ\��yE�`~7�Ъ���_��T-�7C����I}�L@��S,����!kLy�+�:������ O4%�ZY���Δ5��Q �jJ9B����\�.��8X�ϒc��E�����Κ�y��Gb�Ȏa�!��a�xt0&w�b,GK7e�5q������N��j����W����4�1�u�w��[K��i�ZY�9U�)�\nD�qE.�j��E!�1b]��<r$������Wh�ݺڗ"�O��$����u��/*i���WK��]�Y�#r?χgN�ށ�'	�D��q�;�y`T�p<h���D0_#㩳W���ۘ��%�Cرb�,|}�u����䮆����/��<
B'��̍a}�ݾ�*����ÉQ�`O��N����Aǳ�b���"7Zr]e����{r�s�=J�ʍ ��-F�j|�<>��@��w�+>����wW:����~�Ҳ͓����:J��8XT�����Ǵ���B��������p$��W�����bW}P�/�*��՟�%�=�^@ݣV���iH�35�Aޣ��eTS�p�{Ve����Y�n0Q�U3�W�7/��'~J�9w����Q�f�.�z�3�����ٝj��󱆬�^>|�W���xo��vg�p���D��{Tl/v_nu֖E�V�9UVt�%���h�D��R�K�l��W|<6Qao�
}.����+�k��� }��r�,�u��۶�S�mȥ6�Eh�|Nq]Ա�bQ�8��H^Kv1���[Jw�$�F%9^f1��Rm�qɬ�ˮ�c�yeʽ3;2�箌,�6�S��$���_�H�����w�o���W;���=�-ji�j� }�.�ؑ9�
$���8⮝(�D�tSE���y��ۏ�]��Z���W�eC5�ġ��L'�ƸU�2�'l�Z�u~o��.�\,W;�.�:%�tz�n��*Kzk~�e�X*UԳ�P�L�8JgU�|ը|��)��b�Lv����̇5x[,t,(xy
/��F���l:R�þ�Y.Ov�ג88ː�]mq���BT��%@�4����Vd_��1NIe��g�/��&��q�B�3�ب}�Dk$p!i�^�bY�/rՉ��t"��m�{�Nfݜ����z�=���%|Ht,A(b7��)Cq�!:�j�d�v����\�C��i�	U*��P�|MhUN]9�����Q���	d�$�Q�rMHmU�:j�AHV�L���tb�))*�c���qn��/B��iks��4�uB�/'%����>�dU�K�I\x�^�.�1|����\��T��$��0\�|���Lb&�`�=�Q�`�Ԥ\���ĳ��*��O�i�W�؜"��n���n=X��ڙ�Z�*#L�.J�6�K�yНna�hŽ��nM�λ�9f����V�-�� ��4�=%!�T0R�.����#X:��^e[���|a�舰��|(i�������gԏ@[�t�S3` w &huq@�p�Z�z3�]�!L�W+�Œ�kgF����\���hCj�A~>��f� *�t�c9���6ɭ͓S�ww%Ce���.�x�����9OS(âԲ�e����w.��ڄ�j��n]�n]"����b��C`@��x{�ek����,���^�ë���C���U���+:��p�Q�: Lt�
ңӔ�m	�{ۘ��y5�q��8�\y0F���×Ze�Eq�
Ie���A��<���5��f�'���]IM>/9WK��dR�s+Iߡxm��9�B?V�j�~�%�O�Y���`�b:Yp!�'=(׌�̖4�=�[.��v�gR�S�}��M
[��j�N�8JO���Å�(.�pT�[

�c���[���>�=M���W�
�z#�N��TF�R�!|z)f������N�5�Ȫ�qc�d�
}-h�eB����e	�hWg�b��P�E�], ���o�96�G�v��Z��Grl��3;w4-����	�:Ur���;�4s�a
{�}ƕ]��u�4�S����l�AD���P�d���8�0nu�)k�N����P4���o̔��}�h�|�Sg&�-^p�x��U�we���/�Q'��Fz#a}7#�A��9!��Mb����u��1q���΃Ej�W*�%qc�� P�~ȹ�RT)
<)����Z�;�M��0*9t�䊈8w�v��7��2��I.vp�&nD<�5��e��9�ϵT����s��Rfu�p�C���] �����F�Ү�Bu�r
d�n�����]+�%�2� �)�z�Lg)������j�mZe-��@�o����ۇwk�E�u��{ZI�"v�1�Ɩ��}���-���v���	\�����mvkBK��%.`�tH'�;��a�����ov�,i�8�6_dU
ҧ6�.�
�]'."�qn���4�y���m���٫n��4�5�f��-���oy��Ҿ�1��t�*�W-e��=0���9D��&���xd�L�<�V�<���9���}����$�I$�I$�Mr:�m�v-����w`4.�&�L��0�m�\�v�B����j��]�Q�;�a��ak��P�>8t��L�ѽ����Y�U���
r��B�b惜[��|u⚨%Ng	T�Z��f��m���F9:ݾ��E���%��KX�fiu7��6r�%�թ8�텕7�ؕ�����xn���jV�p{"���˜s����^�3���������y��Z�WCC�J�sd�W������&�Y
�7�;�PW���qg�,�4ʞ�5�ͦ|�n�������Ƿv��I�%<04��xEun�"��9�V]!�>ٻ�	
n�z^���Wi�������t��������2+�����U�$�)�i=�4���BŮ��T��+������Fc�㽡f �΋�}�J!^�M���B�8���]��\��Sqsn���;5�MIv��s0:ԝ�g����N���s'�|�C�~�}�$-�J����o��yh5l�Ԡ��q�0ɨ�YQ�}{�H��Xd�S�:�Τ08fF\�|�^j�Gq�mH���D��M|��#r&ۑ��!=����L��]/���4H��k&tߌ&zoE����࿗|����y�J4r�=�z$�z}�]���P��؈���$��O׏{�Lf-��R�)��Y5\�n���ش�.���3�;�������퉕�F�nJ���&��>Ҏw��> o��Y�]@�O��c	礮��o���^S#C�X�RL�c��D?~�]hif��G���4��O��_k/��1k��+ۺ'���<y>�7��'���_W����{73���}�-r�(��|�:��|A������y=�ϠV�Y��h�/MIjK��@���R���ѱݕ��>����^Pϵ�^�d'��ަ�٨�(����0�����I>O |��3�����җ4��(���o����>C&B3�4I�Ƽ�~�y7���鶍��<B,�=2!��/���t±9�lSgWr�BEZ�cb�F�Y����5���N���I�Ym�-s�T��NJH�j�����ս�������ahd4΍��Uh�*�Ê�"��(9��!u�֗r��,^�c��Px�@���+�t���d����Y�t�sQt��4�nf	b�^5~:*K �ǨA�����wμ)v"<":)�9���{5Z�L�����3cbJ/�	���)�'�+ڈ!�J�R-�߻�W�0X��nf�P졆�:gne���c�|�v:�V9;�l�w�ԩ*��\w2t4}[������VNXmxh��LZ< ��jmlᔮ�����+z�*�XnQ��/ *�,��(�Eɺ^��,��~ʼ�Io�&z�����=z*}J,�w�y������p��w6d3�bL��L�֯r�Բn�:<����`��T�8W=1	J[2�H���N�!�1K�����R�M��1>�с����Δq烤D�=�2}�UzL����<X�\���r%��Q��P��������~WPs�rm���vVɅtc9^��e�YK&'���]��7�u�䰻7^��Y��W<���	�镸��2��j�gd�E$��עZ���J�M�ӯ��Io�����D�S�'�鳂�Ģ�Ċ�����Y����Pv�2%��Bg\Ɯ�P�ؖ���d� �7Yq<%��4Ni�3�[���J鎢��}l��ܔ�ff�,S�L"@
^�W����<��~�䘰^R���a��~bӰ�b�OB�_t|+E7��
��V�X��l8d�0�H����';v�=P�9n����BC���AU�|�+�!�Ҥ|u^�c�t7޾�S��'YS�V���~>��#)�c�YC�l%��� ��g���x3����Z�?R@vҵ�����B4��T�R���yB��#����Ԟz''�9u�8*
��J�"�*an{z��"͑���&���۽|�����NkJ&��/P��;,p���d�v6p��c�T�E��#tUħ�}�`��>ؐ�SW�w\�o�d]sÆ����|���9~
�ﶰ �ff�;tk�)d��G�W��d�O�T����z8-'6RwΣX�ǲ�3��K�]���^��v��̈����ȔnYno��$�B��EH��c��Iû�Nʖg8܋�%9����/Pt���b�~·�,�o�&-׹W,�<.�b~3�q��z�Ncy�!���oc���,��X])��}�V�&̯�iV:M@Q�/�Z�1YI�$�{�ԑ�+��?R�z�!��Ѱ���^�|��U��;:b�է۝��48ed�C��Ppu~���K=���^�WB�5���gO��Z�M̞�cc͆^��:�T����JO��?_�.��u�9jݷ�H�.jW�	�伈�*�d�x�f�P�q�����'�:�_y?1�RN�_)=��
����S�����C�df�9���Y��Q�g��%2)��6̽�zj���I=�;tr,p���-��E�>����ɋg����b�� P��0Ow�h��q��e[��C���9}��U����ɋ�K����E���M�}�Wf\UѲR�DxT��I�����&#²���*#�9�$0�	��lw��#�Av�+���w���`?d�9r��~��q
I-��6U����j��q���<JD:Ŵ4���ܬ���4�����]�EH.��Zw�E����W�����c���xwsw�D���uw�(!�X"�$O���}���V��^��l�J{��`��o�;�Rn��O�E� wH�1^J\E&Y�!��L�ƋQpAũ˽.�]���՘֠9j������{�h�yQS��i��MȍW}���ӯW+��5Cl�aC��M^d���b����`���۩M�5�k9��3�ُ�'Co*�"�L��p��@��vӸ�x�qf�Om��BfT�,��]x�]b���aB���9S���ԩTˮ����V)�Jg��9�T����w=Z�d��S���࿜��,*~�	��A}2� �⡄�C^�N�%�wj���������ȫ��x鏋)g�q�aѹN1xx�y~��m�/g��Їkip�j�t���w��C`@�t(�A|�x���h�Z���w��R	e�sƆ9f͆�<Q�.�cTq���z�F��*�5�߯V5*U��Ӂ���^tOVv�X7U��!PNG����Z��N��g����۰O`��hݻI.��H{��:_��u�J3�oM�#ڍn����V�#�S����^fm;r�9��9�%nvH�����jA��'�ΨlK��G�[��nTXE[sӼ��o��%���m�C-cݵ��*���6I�"4�����n�SO��*�u�ȥ|��������+x�ؼ��Q��=K��j�]�C�f.!�Qb	�~�S�yE�rխ�OR�X�W�ת�׉��P��| u~�6�At0Di�½�X��Q��K}�ψ��,|V�(�]~h:������`o�����.�i*�Y�}�-��a{�|H+Tc���0v�3$�n۲�p��ٱ����T&e���f�Hg*�z�V
>-�g�O2
0u��g�,�:�؈��H�r��%=�u�� B{�P�5~�������������	{���Ԩ��1�4�f�M�d�*���WlG�,�7L�\KC#Hc��;X��*Ռ�_!{�j{BO9�����-�IQ��6y]�ᓮ���/���˃���	�k{�Q*��GJj�Kw�+1V��f{Fe�O�;̼�SqDs"�k�������[Y˥1{��Α�'Y�8���
ȋ�n���+s,]+G�����9��6=+�z�f���� �x�P�I�ԑ�R]�z{�j�E�E3kb�{ӡƚ�����q�Q^"�&��7�<$�}un���s�YK�-�.)�"y�3���[,�'XU�&�	ڠ̈́P���]�N�~[�76�h(ȸX�."����ʫ�m�i]ʜā]EO��V%��N화}e
�uuNK��'>I�񂜵�"}�T��/d���^������S�!"0��,g�x�@�]�+�+/�A��g7+��a�9V��<�|u�PQ4l�BDhE�&v�F%�A��^7@��U���3��d�\����0�R�!�vύ7G�iVǉ�*��ᕮ�T��L���zxh�*�����8d�T�ȋ"C�&�
�[`GK7�{�W���sybKږQ��&\�jf�S>'Sօ�d��)���~��h�zK���:R�8�����?L�C"�M�%��!8�(R�`ۅjV�x�b��d3��V���ݪ��I�1\F]Fuya�m��9cj�ݪ�a���V����R�,ά���>X����̹��6w��kN8�9�X/2��N�;ʏwS�%���71��8�7~"���2K� ���48)�ɨ�oy�s�f!h�����/?o�|�����\�4ŭP��z׼}�G�8 8U����t��=M���v³)�(�]�D.��:9�N˪�����6=+�1��������Z�	^���ْ.�N� [S�3mL
̲��3�c㏝X��4��Vo��zN����>���crYj,���)y�:l��͆�*$�!fո�j�8����j6�5��4~�(�l�p��JC8qE�Y��m�Ҷ2;�'�^��S�`8ɾ��:j��6X#<-K��(���ŚZ�N8yMUZ��D�Ze��Y�\j�ॻ�<.���Lu����~@TĻ��Ёlo5^��j�z��U�X^�S�Q��Z��)��`�/˃���z�U�	���A�y�,�og���i��/�q�Q(�x�f�P�V�Cjձ��L���w���]�1XRb���q����_�e��IKl�䩻�)v9}� ��<|'��l��TN܍�;ƌ���������V�6﷝񉗙�MA�/7[%,�\��t�jQ��[o��l� s�$�[��rw�Ô�s�nŠ�*_�����ׯ�Ԡ�Vf�l�XS�D��N������Am&�;��u�W'; cYK�w:���晗�Foˌ{5��������@������>�R9�v����u���VhC��m�U:����=���v�t�]3.p�rl ���^}�����-�KMš
xb�#K�Fo��2h%Gs:�sB11�}���"����x,*&fP�!��Q{Ʀ�:K�ؚ���ܵ�u�Y����O�T
vh4n�1�T�����X��Ƴwj;q�c�\���,py��Rx[qw=|:�loD���ǵ8e�e�\%�O��+�������εb	��o��Ĕc�ɸ��M��/��?/��樓�ˆ�	��~N�/1����v�Yu�{%vN
,���\J@-��S6j�e�v8�͵����g�M�1�sR�xN�5�p��Ŋp(W2�WiynU� =f®�@��7/(�s7)#V6�M��<���s�Mi�;�I}�Zd%k�V�+�� ��Q͞�@؋���M������M��O��bq�*�E��vk��'�Gj$��c氽[n����bx�q�tЀ��V{�~��q�;���M�2ڏRT�t�7��b��`h/vr�ӌ�W����ke]Hq��r�i��;u�]S�S��4�<��^���V�r9X`c+ؙ���L��zꩥ�;V���R�6�hŗ�Ut�X�򠂀'AS�(NTוQ���G�9��������滫fz�$��O>�����@��I�4ҾݻȚ���s�����"���w�ӯ0e��E���\�hZۄE=�n��L�cCR,t��=�N��A�L��/���M]�Y=��nRz�Vb�����\��.P/~��P7��T�R��XM���e�G>���}Yl
:�C%`�8f�fR=�cu�ɵҴ��J�a��ob���%F���N�t�bB�Fvv6���IG�z[��~g�4W
�2wS�'rF��L��A;�����sG���ɚ��ĺ�
�H��S)<&���V��w�b������%���o��wM���:��Z��Y;xgo9�w{�K���Uw4����F9�Yp�����]g8��<\�5U֬��۪]��	mEy�U��B����j��x�&rv[������^keS�o�-��;u�P�9�\t�����s�rp�I�bfsZ�ˢ��o������P.x�5]"��K�m.�D1<*5ϫ��w/�ϯ���.�UM�x�N-K�����c�gP���YEK������)��̀��}[�o3�QjI���`��ͺ�R��5�-�j���u\���}�?��$�Ҋ�$�I'�J�D@Fҏ�������"">oG����TƮSZ���/��|�~�1���Hr"�� O�� !X��-f!q���>3��5O�7����0���?������>P9>s��>8�_D�}m�����d1���c豵���_���k��y�6���`�{�cM��D@G�i��?.|/������D� �U��}�)l}������A����2������`���~ߋ��J>�ވ���@�+�l��|d������&>����F�p~pp����Š��k�*�]��q�������)ύ�?�Xf������,���bv�j���6�	�� |EP ����e�N�h�X�V�խ��\���x?����9�+�3��q�>������A��Ɲ������>?R�������G������s��>hF�~���,�P4���O�w�/�����,�Ug�@S�������&~���ĘO�p���l?w��?#?�����t|���?i3O���G����;�!��Gr�����(�D@G�����q?
*R�V읰~��
��&O��P�d�ZI��Cf���O�6?�@FpP���Ϡd07�\-ޤͪT)!���0�,�sG��J��`���.(��~�������������`��� >�?����o��G��:}a��!������������?T X�Q�/�����?��|��������%q�q���;���?�������(���o���C����p���\[6��O���������z�$�?P6>!��ަp�#�l���,��u~?8����~�c?�#�����?w���������"?�}>�������e6C��Q���_�2?
5�澽��A�S���	Q�0_�a�A�������:�}�@G�����2�d?W�ˌ3-.Ȇ5o���k`�|HH�qB��#����w$S�	��