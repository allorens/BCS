BZh91AY&SYO���;ߔpy����߰����  `�����=h���@ ��
�تJ�QUJ��       ((((  >R H�QUUc�  �h�Ҋ$x���Ϸ���u��7�z뷽����]��}�Q��4����VveZwgF֡�;}���gT흱�ބ�4� ���;ꭾ�v�-m����9绷eK�k]��ÏX�@���{��}�sֽ;Ӷ�sV�k��vk+Y9W�K��#������]u������Wu���[wi�:�]ڲ�W�D;�-����9��ow^�Ӯ<s��۽�k��q�7� �{��|�M�u�������m=�Z�y�'�>��o�
6�p���m��-�q���z�t�G��H��/��'=Ǯ{�R��Ν���-������o���ϸ����6޺���V�vڰ�       % ��*@� S��=J�H�4M4ɦ�L L��j����H�`  �  LL	S�) U* & L 	���&j jJ�#��L L���� P�hMɣ=��S��F�I�4�F���HJ�	� `  23Q��/��O�$-����$,}��������DH$tH�DA#�d?�U�n(U�_����҂��C1��I�$�DY5O��S��e�p���  $6!#!:�UUX	� U �C���O��e}�������Q}���:�[�N|9�(�N�mgΩ�|)D�Q(�l�h��e��ң�ȥP�D,[��Ҩ�����<W������=��{Ec�xI�t4�-����[Z!���ֹ�T�ʪl��+Nq;��ra��Rh��>j��@�"1-N���=1%�*�V�]�3e�ctD� �"*����e�F6*�	�zŃ}��Kcz���4]����Yǧ���r�.�[�qMg���+!��CT8���K�l�9-�;��Q�[��E8�k�N�<�=1�OSծMn�e5��e2�t7DB���
�l^��Mcc� �p;���z"���m�`������	�6�����+0q{۫z[�ޘ�ccLq�N8�f2���m�C��+�P�6���(U�cwn.����f81z�_����v�s�ε���x����#X�z:�7x8ў�	�S��FmO+�l�9�88��ǜyoU۴c�k�k��1�=�D�Uָ�u��&;�,S�q]��81�k�j)�C��[2�ৄ�f-*"a�a��rDFK6S�[	�3�-��uNcUej>�3�D�d����ti8u-�R9^2s3	0`.�AA!Q�d�k�y�H��2���i��i�y�a)��4�&ַ�6dD#Sx=q�X:�����E��LC�m�9�[s̘�خ]�y`�V:�����P�M��N#Y�AZ8�T=����N#_�E9-���\-cg�d=l؈���P�_���w��j��S�:��pS<�ۀy�Ǒn"Yq�{���(j��1�C����Y��[n�舉��EÉ�z�/5L^h�q�2"����6����n�z�#���5��\��ǘ8�wn��n$������4��ю"��L����z8!�x�T8M��4k�~���f7v���n-َ+��屽nۦ[�.ƞJh��:��<D؅L�q�c������	���i�i�i�6c�kJ�c���1�������q^�p�(w�M/6RҴ���Ɇ&��u^�=��UVSY�z����)�C��!�
xK�y�b�͈��"!��%�
xL@z �8��m�\DC�2\d8lǉ�8����V�!�˩q��}T�WǙ,F��/u�(�2�y���<��H�+!���N)
)���U�!�ɤLW�u1p�ʭZ1�*t���Da��in)q�]V��3����+4bhİ�i(m2�<�b�V�Y��K�%���<Ũnַ�Zٍ�B�n�x��( M�o�1
��(*#�8��"ر{ؘ�<G¥��d1j1����B��mʕ0�L:B�9�v���E82�LFyz]�b�fc��M���dD{><�ZdF␦آ�B��_Y��+;�"�caZc�9ʫ3�@�G�oS�#j�R�i�����6/yg��j �q(Q�^#�@�\�^B�^Ԙ�>v=��G�da�ƨ��:2�<g^_�W�Y�G���/J#b|!���R�k��"ߑLRdD��XLE���n"��L�
Ѯ�p*D:�qHW,�qH��"�|/�`b�W��b�fc��f�&+D<!������
�B����
���SS��LG���W�k��t�z�X�X��,R�Y�@�ψm
1]Bp�SB��_y%i-���Q*�^l+Af����p�E[:<.lы��`��)�+��}��Z7��-z��X�!:R���T!\�a��D20G�8V�4wwFe6d��#b��ΉȠ���B�B�v�!N�xp��|=�&"�t�q-����E�b<��K-�-�����T�OΖC�,�ӥ�Q[h�d01g��b��\4f:+�Ϩ��Ȉ�,%��؍-�!M�T���.a�f_�����F%�ʢ��+.!����q�,��R�"p�'�y�g�7��)���
~�?ye��*[+��RE%R��4%b�7�
�-8ja��/;A]�0N�X߳S���}�~ŉґD0�kEbe	�ɂ>�(�0��	�2�2S����1z�1H�L50��Ra����50�ַhT��W�g�'�%yz�U6�&,���"�[��-����R8hݘr�p�{'M�bdØa��b�J!5?W±8X-�	��}������u��ByN|ի�7�7ɄC>�-��H~���5�Bы��X����Z�ԿB�b�be|�]kJ���<�)�}?g��D\2b �^�hlG�S��5����&�u�-��-��^xu]��K�۱;gyx�ѹ���o���|{ǰ��L����JڔnQ�+�8�'�m���P||�[U�����&�D�?F�9���l-�%]�_|A/��?�Ͽ��ǲ�D¸���6���	0���a(���G���������ِ�~r�KN~�Ԫ�i(a��P�x= �u�5�KC��薢oU�e0a>�Ϡ��ޯW�E��e��;�R���J�!�.�h�^5�ռi����7<��+#a���H�r��r�b�{���NZ���?r$�S	h�]�waf)���i�N�����q)��`�\l�����C�Rf�ی������w�q�^鏾M]d������Ho商(-�+\��ё5�4���În�C4�� '; �|v�>�郒Խ�5�L�u�G�v��Xq��CҺS>���ԙ��f�aN7y���� ����=�į��̕%��z�O�c�t�:��vsm�w��&r��g|2�O�W���|{��Tm��pZ�v�-��:�GS[��!��dՇ����Y��W=y�~�:�O{}����@mB�3��o�{"%�����̺�]��"��T*i���&����ǘ�����=�]%� �@`ɣt��n��y�Ǚ�9N�z�\5fۥ���3)�6O\˝�F^opNS�Y�jPdl�1ж�P�G$_O{��O<�:����L9������9�'�PIiT�I�B��;5�gf3��M���*�i�aϣ)���6�:Z.�����ڋ���b531�\�W�8��2�ɇz�H}�������q����U�?�O�T�7� ���|�_<ߨd���y�ZK�܁G�b9g��6�����ʌu�p�{[�;$�	��,��=��R�c,o���9�Nl׿�3������[�x�舷�mkw]�Xy"�fu���O�����7�s|x�ョЇׄ�z_ݷ~�+tD١,�w4�s�"��:y�_%��_e�3�O��8�q4T�<]˅Y+P����o\1����S��eT��mD�VR�ee����E�)�*�!�	s�V(�p��h���~ϴ��ٶ��;�Ss<ͻ�'�W�8�id��z���×�{��+*WQNv瞼�K��9g�hňo�Y|G�c�Ь��q�~��Ƶ^"H\|E�ɏ��I|�)�Y�iM����|a^��#!��UD�c�Wļ�\2����rӌ����4��On©햰�.����fLy�t������.�vhD�:K�s4' �}�`�'�W=lϺ�bq��ņ2�Y�2kG�����)�t����:�����wq�1s�ד�e5E4���Y?f��E=�-x����g�5x�^j��������g����9gs�L������G���;.h��Ƕa�ߖ#�sܹ�� �if��g�o��d'����*u�����\���9X��oy(ŀ��O3�j���{i1cx�\�;����,{\%�;��x��3=���Pab���a$�+�9?�l$������t�����)\�q5;g�tٞ>��j�6�������W���+�l��iq����^�~><?t��]�S�n�l|{2���ڍ�%����Z��̻)�L\�݇���#4ZG�ծ��뾽���dn�x�sͭ��¥�*��ybf{%Ų�{ӯlְ��j{s���Z�&3f˴�87��$e��Ӈ����>�4��B�8Y�C��2okl޴���_��ov�R��t�p�7�l�Z�8��6v̷O����q�sfҩ�G�o�U�2�/n�zZ����u"r��r����u��hE�O_f��K������l�}����A���-�}��7�>%��X��&9��ni�B����Q�8���)��p��?"H�	�C��ds2��>4ܼ͍s9����⌯L����U�L�޺;���v��#x��GF����}iK�sV��ُj��w+����P��*~߰�������z�c�����}�=~مq�9su���k��/.鷻�k�B�.���o��ӽ��Fk)��o�'�QЋ���L7���fe�������P�%�
{��h"R&�Iicy]y}����c�������UťG}�t���$��o~�9�3�Ӛ��
V�f�}��c���n6xT8���L"a���Σ���aD2K%6ʧ#�+H����A�1B�0�ݛ~����"R�SF���(�~��i��F�m�6��;�?l���	�ԙ�)�㓶K�Ǭ�<>���4��rƁI���n}bn�f�:�Z��ųp�UcNge���d�re���q��P�{�rlsw�A�F�{3,<+$̢v��{�]V��3�b��y��D����T �a��?jG6�67gۂ��3"gPf^��)(�Om�$�:��%�I�� ���)�>bnp������)�@u3�)_-��]�L¾�I@Ԓ9$��0������{��;�CJ��@��L�&�O��W1��k	�PU��A�Ղג �M�T�3�`�p�h�u�QUk�� ���o�?�	���(����=�pА�O����I�~��%�a ��z4}
(����}E����3V���7`&F���2iB����uA�'��qFe4��D
�m��A��D1�鰑썐����"fY4��h��4���`���W"J�+g�c$���ܦ4�f���gmY��ɝU�G1Y�KI-�4�RZ<F4�+�gن���V�pG�TKř,Zcd�̽�7`��K�Q`�5��n�fg�/���c�8���H`���O��F}ەk	l�	4V����s�hT�K-&KD�BIq�~;�`��4�i��)p�+۠��"�n0��I�b$u��MW�j� �u�>0�s7هQά3j�2��3i4~���L����P�F��/gё���l~OI4�n�9��H�[��2�$�X����Z�g�\��5#02(�=�^���i.9�4kh�TfF[�&~��4Qcq�iN�X�T4A�~K�`�%����fI]T��mk�1t�d�7I����A�Һb4e�h�Ix7�A!�Q*ǄH�(I-���5��ȫ�Fq��	ͨ�-�����Č���3��dg��I�ЊxIu�I�R���I�(M�X�XjÂ�̬��B/ ,F{n�Y������=���i4'm��6���2�έ�A�I�6^�����{�GY�q���&Y
�J�Ԣ1��A���eI[Zgwm6h�X�F͝uX�����_*�$����φ_=��BALU�b])/;���S��ߑ6���">�1NdH����h�p�,7���6�a�"�>x^���e����,�<��>��8M��n@ɓzv�M%�+cM��yu�3Q�
tU���H`��b�ȅBbc|��n�?��|���Ϩ�!V@EA۽>C��Ҡ��2p������l���~G�$� �}R��}��~ϳ���s��� h�  @ �@X 
 �@
 � X0  `@a�r    n��n� H0 4���� �}��/�_K ���<  �� 4B �� ,  H  x ` B 
 � X���{��X J���  �_|�����o�ҙ�  �< H@(l    �  �� �	 $ �  R   *���wt 	 Ҫ�n�� n���������ܚ�}������  `@ �	 ( �ЀD    4`  " 
 �   P� n���n�X $ *��� "����$��H�H  F �  X 
 �x , � h�рh� �<  ,    �<�[����PS�FH�~_|�4��I ( �   �  XP� P   `� 0���  h�b  ��Mݝ�ݐ� �UNї HP��Aܑ�$U��
��O�����$ID�6��o�_���wg��? ���2�����j�ݶ���6��m�lٳn��էo
xxv�[m�n�m��[m�o]�Ҷlٲ�ڴ�n�m�n�m����|�;i(B�b�j�j+B�*^B��Jٳfͫ�m;m��ݶ��m�٣f͛m[x�m��O��>>0�>Ӟ����^���:�ˣ#k%�{1;�)���Vr�~���>Z��ݤ�2o��;ΐ� ��p�D�=�W}����xЋ��i�y��ӽYػ:\�&Z6�-H�.���"��)�BHO�f*cH(��B�<�(k�3C^wVɱv���n6�[mͫ��A6���͎�p�ݒ��h�Y���t��d�����V��\@�Tc
��K	��39_es�V؞u�;T��4�H�U�����xq�g���'t5�.6�۔�[Q���)v�ޱ٢�wnB"y:���*)�	�8|c(�I��$��q����!�5g�"n8B���I14�N_�wxv]Z#�+����yef�"���oR^�wB��K9seYo1�m%'5IF��J�+�%�ۙ��{�|��:�(��{��������c�*'N����{ߦ��(�=;�����~��d��*w���q{��{��o��ϻ��fo��7��$��a�*��q�c����.w�S]fn9��Zm�CB�V�`o��I�n�JbF��`�a�����:��x}i2amO�#��Sd��͈�n#�-��b�'�η���!^$�i?��i�G���HY�x�M"Y�y��%op�c�J�h$r�/��ś�����=�0ܠ}[g�Y ����ղ�sp���9�G�H��������0�UW�m����!�����R�{Roj�Xp�"*��!����҂T4U��C0�Tg�0H��}-]ST�h��]2c�ݗ��)[=��l	�NX�Nn��mD�t�t((����!E��z���Ĭ�
�i�0�KjT�nWF��rY���!�*�=��'P����Ք�����*+9�I)�9K8��;���-:��h]t��J4nV� ��`�UT�Bp7z^��6B�ɿ'S�'Jvc1⪶��1�+-1�uest���.��&��5CL�珮!���0��.��r�Vef5�v��<����,�ۍL%�T�h�K��c�J&��k!��ʝ��X:r_��]-�A�?��J �t�!��Q/I��Y��R?�{�v��(l\���dU�]�a��I�
�'��zYd{*fR��%h9c��_'#4&�I�;n�H2_4JP�)$QtѺ�yD��~�=1��V0n���ST�G%��DTV�
)��\	�����G���y��ۿA���AdA�ZmO�&0�V6˲�E�U#UW�6_��鎝�)�c�Um�Lc�~�򮧷�M&�����P����8f�+��M5@a\IS����2�w���R:��
��ΰr5M*�����S�*P0�l��
D��!�-1�)�v�tՀ�������-�ڶXߜ���c�: ��U]6��N�R�3Y�N�&�aF��Y��*��:qu��8O�ґG�4l�aӦ��y777�'��Vh��d�w$�:2(��y��e����n�j2�R��M��T���s��se+U�X|t�|��,��;>ƽV�ϒ��Ub��"��ᱺj��A8ss�>�{/���{���,�0V
H��MJEQ7J7�TkM�s����0�[3�-�ѹ���v0��zBf�eC'%�¨w�*a�;��W8h��Fá҂�/�:p0�1�X��0�3QD�c(TU��n��hˬ�Yr3����$(ɼ�w�=�G6��璐d�}]�χ�W��Y4�-���˖�-�Sޘ��L��$�J(rڂ����6�ݵ�*�]]�������S�C��Sڠ���'���pp
NV��;��������I���)�,�����2���V%Tݹ.�tҶZ,���m*]�߬s����C��锎�P,(0��K`�a����:�����|5��р}π�ùj,�C�2ra�p��4�;�����P7���0Wzb��2�FĘ�<Jr֚���.��*�Z*1XzaGp~8n)�,�wi�X�s�T�T�D��-�>F0k�#�J*|(�
>�O�8Q\_��.;q���Ǭ⸿/���q~W��L��Z�+�W�W�8|U����h���(G�t�q�/��������x�q���~_��1-_ŜZ����~+�~�R�+���_�
=�s���q�w�fg�����8�.���q1?.Psp'�P��!E���J�������x�x^���zx�=�}m�/<�:q�,�L��x�xxg
��5��{q�W����3�G�Q>P|	c���]�ڿ.�9�FRa3F�'d��-R�K�w�ˑ�V�M"K�0���7����8��p9�ۛ�7�G
�}�6��!��[&+�N3�k�uA	��*D��/����<qo�~���^���L!��������6�fw��7��wuL����o�}ϻ��fygwD{ͥ����fg��>�Ck��wT��-�o��wGww�]u�>�\��)Í4V���\q��Yf£�(��,#$+������D�K�$$O3�-F�2x�c�ͩ�H����+��q��1�L�UZ0�zm(�C)lVr��m(�z��/k⯊.Z/W���n��y��˛�"e;R�l@�4���$�B��%����.�DZ=�����^�'&�F	8	�,B�QbF$��F����?o��j����ۡp��cԀ^ti��,	r�`��,��,�}���juQE	�H����WsN��Ђ�0�&��T4�6�6Ey��~�h�]���63�apa0d;�Z&�ʈ6�%DI�)��B���p�ه��P��ʳ����4֭ƝG��X�*�u{��iq)$I �# �(�nǥ�H�(bM�a�	�JR1���`��g(F�`8%
v#�7ߍN4����.X����<Ye�Y�������t����v;�.�d.��t�Jim�ۦ+&0�������;�N���R�6,c�ed��w���%�H\Rj���c]�X@�ʹ�۬$$$$$�n�L�Ĳ�I�U��μ�umry�}�m��ʜB�*^NK����*�bU�o�4�1�X�yZ�e&���ǂΕ$P�u�K��Rq���#�*̝�f�?�dx~�	���a��Ĉ���qM�"M���C��!F����T�r2�l�K�R��ȍ0��(��ٗi3�N|<��$dH���G
V�ڃ��Pc�_7%�!b��<X�bś#���h6��(���G�mj�wT�Z5������Uum<2��d��12M��.y(����Pa�8l��j0���[ﺜ��u�zm�Q��<W+%�W��lT]ҥ]5�Ȳ��.��Iy��S�e��>9jN�ܒ�Vӣ+��sF�����6��Y,nl��m���8��4�i������i�g�~���՚��9�\�QEh��t���̾v@�nyxZ��,\��)���Gf�6p�����`/p�z�}���Emf��_�L�n���ݮ���i�8k�p0�5�@[,6���	<�֍C�o"f�!:�[�47&\��庁��/��1��_&�����(4P�O@��E)JS�49� )*U��"�,'��xN��ð�������3�B�����E����TSH��5TY��P��y��M{���%!�9rv35%U�0���t.�n֞�%QUU�wt����v�қ8t��l���o�3%r�p��/����.��p��JIʵ�OG�I[Vb���>|�E)N����ԲK�'�yfc�kIdLhb�b�I456��=�n{CL�%kY.t�wn��K7o{�q%�0��5G]Y�J�X:Yr��|%��R4�Ws~���rzO̱�U)m����n��K��N�R����
 (?�͍�$���=p�@�a1ĿS&(��9���t�C��C� �1w�![h����r���<���M�r�^d�D׎
i�ސ�Ӥŋ��u	�!vf������1ٍ�i��i��'3�!��Eh��f�*덧/���T?L<h�Q����Φc*���ܖ�P#�z����=L!�@.�Q3ss@-�Ln��n�S���xtG�c�u���d��p�t����n`��})��R�D��4�����xnwWy�Q� �8 �$��$|���UT�Ӌ�f��4�0�+���`���#����j�LV��ǳЈ��9�~=��m�ve6[����l��i�a.z�%UJ�_4��U�{�gM�y��h�qA��R�P��X\���Dܰ��=��/6��g�5��C�?s���8�O�N�����NAi��K�.�	��M�ZX7�J�+	��ܲt��DL.��ӄ�d�
.��n�v��{��Ⱥ0�a�+LxcoX�4���G��$A21Y��fXI[�,)��;)���QR�!��Ӌ�P	e�z�26X����?RUUT�$�V�n��g������f�tW�]�2�ZéT��kаW�	WӍ>�i���z^��,źw�D�\+d���]Gn��E*�*���¥�
[�N��(�,��Q���D~�GZ�����xWk�q�8�+���6���[c���_ʫ���W���!�z(�z��ҧJ+�>:c���x�|�,��8��3�x�;c�W�z�\Z�]+��bI�d�Y�J�+�3�W���o���k���칞>x׫��y}g�1�mx�q�^>m�7������:^4�f+��׌�x^.=g����{����/<\�x�'f/ū����W�]����N?1\�j�~\=TG�E
%�4o�{+W�~�n��A��w���Cb)��ɦ��e?�f]_lS}H�ۃcc�]�3�Ɠ�o�^�vA<f�~�F�Щq�����yt�k|v���U�[�*��n�{) �A��e�?�<��@��^�^�vp��ª�����۫x��\F�آ�^삲BC�&C �	����q&��q�M+�F��"�5ݙ�a,��?A�X�������+c3�>Ù]�x��M#=�O��f1�*�8�ڄ�:�[C`��56ѢhQ㴠��=p'��G��~��j�ʑrNA�̧��nV��KT��µ�L �(��S�9e�6�����>||<f�B�\0�͛vĜ�Q�Z�`ܛ~$e ���N�mԓ�%ۛs&�0��ݮ�/Q�i��C�x�o���ݛ�柡v�Ӆb��Ln:�i��e܆������Q��V����L�t6�M ��R2�N�y<�7�&&�Գu�
�!B`��c&���u�`��gl�FsB�����* ����qQ~,��R6��t�ٙ���k��{g/k�-I�ȶ��),h��^>yk,�nl�Z�XMe~���y�4�ʖ2�+Y�l�?������}�US3�]ߒs��{���g�9�����wS<��p>��˺���C������C������wU\��p6��ɨK�)��}����Տ�c�٬й���bme�d�u�������N:8���kf"h]�g4��#H[i/�C�{���Ė֮�>��TQb]X*��	��K��0,�q��UU��i�ug|%e�=.�w�Z9Oh�+¢"=�8�ɽ�Q6ٱs3D��(�-�8.g����Q�K��_�b�/��!�Q��kL�M�Kڗ�8�J���$�k^zѸ�������Z�;�;��K�|���z�t�Ҫ^��3GM�
�B'���>��L{~���R�x�R�ӡ�Fuћ\
J5�m�r����J�2�_�s,o��I%��<,�wbe'Q��8/�q8��4��OK+���E�lU��t�Y��xI��Fl�lO9���_܇xC��h�,�-�K���$l�=0�ۖ����UU��|i/�h!�!�DO�OB"S����G6�rCA��r�L^�4����$�3�´��h�]�� ����H@9��L��>i�\�C��=��������mf��,��V���3��,��7���S�������&�m��8wLs��#�8VXr���N��y+r�Up��=g �Uxn�T2��p@�;�a�O#֍�V�Lc�O��c.�OK����(�ny8�I=
�� �S�9.gN�H뤸x�z���BFM�i�F<ز��.]!�]�zHՒ�x�l��e��;{Q#J]!���Ib�)�ݗ,�)8y8r����K�o���9��*�Sn\7�u�9L6��CL���iN�K,�`�<�!D�(���DD����� �K���2�a�"ȟ7m:$�|�6�I��¸�Vt�A8�7Έ��^�ӶO5���7�w�nu��b2���Ct�f�SI��d-lKKi��%��׶chf�2�R���io,ԫmcm�����k)�N�,!�,���m�)�I<�Y���j.�2\ˑ�Y�QdѣLH��̌�����݉�����Ӿ�S��3�@jf�*S�Q�u;�Tt,g���Q��L~�bO��K��9��:�r�xf��2��Gc�8f�g(`�lܔ�ҧ�ǧ+
�1��WŚw�_�ݪ�l����p!��7{�:)4�4�X��e�$���8h�b���&�e��.�ć,c���UO��'���u��I`,1,�Ozn]�Z���R���*��E-�vSe�,nϽ̱Rt�\h��;/��b��_e��~72��0����H��5��=�B�'B��C�L�;��Q�G��]�^�(j�T���	O%t侌:u�6rp���p��I{�m�]�XZ���5!�Z�l���K&������b��[K���l��Μ�.��Oo&�3���a�*n���P ϭŪ�H�7Q�pĺ]�1U%PX	�T*eϣi��#���[�Ħ=V�Ep,�"|Y��J��[mAF65�%���7�c���*�{ ��M0���
���5��I��4V�JQFnz�=�~�����.ڠJ�N��ѕ���O>6zHs _X���nܹӗM�۶��9�ު	S��g�̥a.� �SGf��t'h���K���D( ��!E0x��~�*��H��!U�e�!"��_ņ��Kjl�RN&Da�P_;��o�I�Q�:���I&Ԗ_��)+�n�+[X�l�.4�=��-�BK��c|&䒌5��gR�2�B\l��7�& �/��=��*�(�'�
zd�%�I�痌�d�bm9'�%��!�P�_��-���a�'ۗ`Q����54b�P�!h������(�X�Vn�z6a�J@��NCr���r�33�ǃ���b�8i���V�V}6����]_/{�A����i���	$�Xb�{�y��A��k��� a�e�h�s i2����;i�����`�ü;|�l��N�UwIH\�~Ү��NC���R�d����jm4�T%��90	�T�,F'ٸr�:r�����^-i���~b�[a�����/k����Y�OZ⸮6�+��_+��̶���qj�1_�?�¯���hh�S��?/J�������Z�Y���mx����*?
?Ex(�"?��N;gn3�2�/����|�?3���_�3n��-�6�ϙ��v�m�V׋����z�8�.1���:^.��[��*�WY��}i��OY�yo��zq�/K�[�q�xW���i�:Z�8�Y��mqx�x��+c�DO�6R<�x��f�������3���{�ka�W�$�y5�;;�=����-�����?M��U�K�����WW[<�P^8�>J��O�d��|}�}����H)�6��n]֗���)��w�.�_��C��w{�.���컺�]����ue�W.}����������՗u\��"5��rj�Z8i�Wtu����f��Ϸ/F�}��v5m��rt����@Txm���7%QUT@0�7 l����؄���P�&@�p��UaB�W''�2k)F�@o�?OC�xrTڿ��@|�l�?NK�Zf~�
�;��:��`oo�cM&��̊�����oU�b�z��j����}�B��Аƕ�?��������t��(��e]�M�Kr�����2rl�nx?M��f�O��i�;2���t�<��M�����1N����KX�|�1pN�H�)ސ�f�C��wj5W}���0@��)e4�XV+M���U��FO�~z�ɝ��^�'y�]f[�^I���"�4��9VM���2�`�er�]�Jy1av6C,���4R��Wvh�C���(����h��!�F�V���h	,=h��}�v���L�^�cE��bICX�ejP�T��
.C��VYԮ��e�+�s������M5V�����%��q��0� /6.�uTX�Y��i��W큀�]��:xD��{߉��9ǾǓ'�=��w QS��pX��d�F�X�+��V�*�i�5x^���vl!��PrvQ�ɇG���!�͔�*T�?�T�q06K��to��N8NZ���dw���x>�V���j �����rA�x�7I�8����}i���f��3w�S�@,���(�gnGgo��b�x���W�ﹷ��.E�S��[LE����N�to9Gy�����Ƿ��מh�e�	� ��zC�B�E�>�A��L6q�
+���#�z)���QM��z2ǩ�-��t���O'�$��9Mm�b��Å8��cPs�Z-}�}�a��aX�6��j�����nʶM-����P�@��,ѻ!�����]���͎�R�5aZ*I%����y�)L�<��MhM�a���`dbqE���s���Y����
"B��J5$(t�=:6�ël�|��ߚ���94�+ۀ�lD�af'vz�զ�տ�[�d;����2[�y%ܑs�i��ώ-��<����\�HN1n��#h�hGeL؎-�Ji�#u�p��Y�m]�%�#*�)���ݦLs<i�jϷ(�i��lݖz��u�h�t�;ņ,k\쓩�z1�,�8�:��z0z��(��eCP��&���\�^�۫,U�I!2��)Ļ�u<x�f�/�&~~y����ⰬW��Zz��`�e*/�jq(M3tQ�oZ=�w(F<��9��T􁹝�Oe�S\�te�'I$Npc��mc��&�rb֫Z�x`i�|�p@3�!�ݛ2���j�d���:��ld�e�hۻ�\>9��'�kn����͜�\R�32��f~���x�5Y;rx#԰���&!=R���'�\�0�2H�΁��H~1S�ņ��kAJ=��fN{�TUk@kw$��2y�eJ![1�ל��ɋ�B�{���d�`5ϛ9����ޡ#���Qή99�>�!�2ym\=	0�v�,SmܗI�M�P����9'ǧ����+��K�M�UT����d�T~�'�'��J!�d,Q�x�{���v��sn&�bڄ+~{�{��sF<zn\:��C�"�Ϝ�8��I�O�+e��rW��,>�����Xzz�N���ź����,�]�z�|v������m	2� Yn��aw�8����(�����7��Ǥ�風JO��+�T��L���[]/�x�ǹxǎ1���,��[��m\q�y-�-^-^)����'�_R���[W��:�~^��{�lq\k.��m^�����>��Q�Gb��χC�9E�Y���G'�Trz��!G6C����x�/�n6֗����q����8?�+��yO�%?c���kT?������|�/o���۵x�8Η����q��+��x�1�D����~|P���`H#��`"���?`�ef���U+F*�
љ�t�W�<F�t�X�ŉ���ʑbY䯫1}q%<�)G�-�<�Z��)f]��>.�lj2�Q.Cf>򐯺?H�LMzYxώ�a뻚qJC,6=�Ź�T��6��ӻ���:%�I����	��2��̉�W���{��d�SDܕ�0h2�9�d/jlFI�X�5#*O3a�_0ˉ"�@�X׬�ܮ�߯֬r�k++��!d�� p�Rim�`���b�d͙��'N_�'��3�<�zQ%�,|Q1y��zs�X��~̜X��n>*�7�A���iS��NWR�Iq@�]��V$�'>D�u�,dyqs�$wV3�KJ"����L���T>� YI�[MɽF�_wK�E�Eݖg�-N�v-z�dԾ_=����v%%v{	B�4�H�8
�q�ld�č��b}��P�P��-#�,��&e,B�1?,p��q�Fͭ��ײE:�cF��9�6GC�wt����6�ܤĕX��f�6��r�$ӌ.�M5c!0��w��m~.�wtDk����˻�]����z���s�z���z���s�z���z�.�s�x���z�.�s�x�\��H}S舟J���꫆�%�$*�Bw���-�e���q�F��Ib��0��=(��&��j�;&Ê���o-��m�ԑL�����p�#;�j�Y�Z��R׳fS2�(,�}�� Λ��ICF��d˞�����}3�OO`�����}�X2�X�Wp�%�Q,{�K���6}2��?C�G��ׯ����wL�2|��=�lF5�#οS^}�>���j}9ſ)��aX��Zz"'����~~���k�	�����a�1�a{�/����%�$�t�%��j�KZ���Zᷭ�p�8��٥�����$�ț�7+u_s���݋u��c�>s�(���y'�����g�(���>�0.zfM��۝.�}���vz��1��7.���S�V�%H� t>�$����7L\�2t��.�C�w��sf���V�Qt���a�2|g�6L�'�vd�U]ST7��K���Ֆ6�m�M�NӰ����0��ꪟC�6y.'���s@�.\�����=������%�ӈ�����₊A��QF��}e� 3s�})�X��I�,g��F�}��#?D��2
���I%U|��ܠz�>>To�D�*3����v�TM�a�;$�셏R�F]7�ys1�����țz}��'*d�K2	T�Y�'��OO�a�V�zⱏ��;��YD2�O����44�D,�[nj˅ꀛN	�A�)!��Y2�hj�Cm&���K_ в$���ImՖY���ӗ��/L8��,]�d�/�%��ya��6���j˪�;���s���}t3�70�(:�C�3�pӄ��'�9,>O�6d�M��wd�8�v����t�x@�{=��������Qf�H�o/��)
4Y6��`����x�HR�����H~4$�vg��H�r�?[eɩ����+b%(J?�5!�P.����y��3*��dmƣI�۬�����;5�41.�A�2��n0�t���)�$��y04�"f���+�Y���g"���Mu,�O\<��}�=���:8�8D�#$�i.a��ʗ\�efo���n0�+�<`!��������������� ��L�m e!����&��ν
�U={n&�y-�Ir:0�ߥPy��EF�����İb��t]��4��?uV'�s��0�߀���!��f�R��?yG�v��،�FmMH�r`�I	4D��OŜ�}���ag�OC�%��	��$)'N��C�7|���%^U�xU� ciOS�d�{F0<G�����A�L� ��2����Sq��5M���_!��
��B��?zY�y�w�}��>�K0�HC
x5�����K驳�D۹a�Q��.�xܳdC��`��'�2T��21�b�Uc��1�)�㏧n�f��`�`�6�̼6��8��,.���=�o:�oy)���x[&�Q�B�Y�#�X4KHKHo&����Y���0[o�����/�6
�5�ab�.�Q��%��ԧ%$�`ؑ)�{�r7�\:n�*��^�,0�Ssn��lh�">��/k���-&0^_ٵ�j�Z��v:K;K���-��X�wVvI��P�m�iɔ SO���j�J��6�'

(K(��(����;iZ���jz��,��=T���c�eZ�}~�l�^ p�*�D޸�5*��iۼ���lx�#ul��9�s2I��sϬ�3!r9���t�r�OР�o�-�V�BP�_�Eh��B���@�9L�����u�P�,��,,�҄O��(�(�l�T��ڪ�W�1�qz_���n1��x�+���i�|�����ū�GG��(�0��|(�z*�U�5�_�����v����q\]�ɷ�z�/��e�cZ��^����q��ge�<|���q�x�6�.ק���<^=�\z�>g���ݼcn3k����x�y���:W�/:�1�U�x�\/�����t����~���Q��6?�j�̫�j�Z��3����\i�W����pOT�D𣢊���G���ĳ�+F����~͸B�3l�]�%ʤ�z��__Ci�g���Y��b�Jo}^Ǘ�@f/yߟ���6�:;<m���\���[��>PȒ��7�7E\%�E�?r��k�=�X���fm�⏛��� �<�-{�$�����ɧ>�m�T�p�fK�+��u�����U���\>��������w>���������w>���������w>�������.�w>����ꪬ�㜷�X�1��UvqO�3�J��#��_�t�."kתчp�ڙ2��*m�"�Z��,�ʦ��)
�C ü�>���q�;J?PN��a���lUQc2��X8��X���K/VN�n��v���Wg��j�s-��w�pٰ]-x�ѓiq���~y�r�ɋnI�t���[}sO9����Ah⶜.grHI=Id��:��A�#�SU(�i<`���d�@�O3	p�>�7.�:L���|�P���m��K�cG��1��"Q�a�CNo��R��+����m�K�&"Q	e1d���\�,A#\`���C���M�jp�#Y�b5�$�KL�t�̀Sm��v��[�^��{ X^�)m�e�B�Ic����<�=�$qεVf;�%���l�m~�#��x�Kt�I�-�� m)�$����vnb��.���\�QWaP�:z�fo��n���m���j�5��!��O����������Ռ���kӷ�1�ҫ*�pI⮜��3%����UM4�ڄ!�=O[5zi���ɚ:y�d��:o�L��9תK��c�.^�/|�)�C��=`���O���:��nK�A�s0��	�̪r�<a�WJ�x���L����1�l"����H6�[�S갊���b���t�R�.~�9�.���rp8�4]�_c��x��c�oRI<cnCAȞ�5?K��ɰyF�z��^��M!utv�5�����Ϟ�p����U������0.�n�K�,�>DQbpԆ�;9�Ϯ�j�����dnw��GGjW��U��_8�4��.%���L-�[���ʿ lgй�U@G��K�vQ/~����8�H�(ݹưqKv��)�h�p��_C�t� x�Tw��{�Hxl�|�n�L8�H�O7;��j��זi.X��<��m�m.T�=K�������8#������k5����Q$X�r�Ւ�$�d�UԂJ�E��i9#P@)���~k1>���+�ud!1a��^X⒄5��עw�[�w)�llo-��W��7��#���6�X��/��O<�3��'��P��C�4���_)���BPRK�2�����.�B�@��i4�L��K���1`i�DH�iA����Zݵim�4iJ�Uc��ޏk�E$�T���t�q0��P�i���m��wu$*�����%��U"S����ߡ���C��n��L�h�欺��8vlʰ��ԡ���K��=�@�������$�8��Y���cgJW�qU��_<���q� ��WC@��@�8�Z0�f�hɸ��f�j�>G�D��߇����@����/�r8f"�e��F����rXda�E�b�7�Z��a�����2�J)�󫓩�����J���Xګ��Ώ�YfҒk*��T���u��p�m	N��
M�4]��8c���z?~R���}�GX� �@��m������y[���ntp���t|!�a��WCAF���{��~��d	��uї	���VIAP�q*
pTDEL�'aB����(�ס���P���Q��(�<c-������2|�/��c�q}q�����^/ˋڱ̶����3����g���|��XBh����O�<C'�zM(�]���z�^��iW�W��ʸ�x��28�;gN1ǌ���[Ǭۍ��8�]�O��x�{���|�-q���^.�f�����x�y���:WKƙ�N5W������|i�/�����\gN1���x�1�U�x��8�.qs���Lq���81;KcC�"a�'E��p"�
G�S� ��֤�~��$�7�"{'�z,Q�Pd$\h����������\�sR=SJ���|��^P�k�#��ޔ�dC�FWԆa�%u6�Q��� Lt��K�4�j���5��!Kf�J��*H��G��ն��spv��A�T���L Ui�H�la�B���lЋY��%i͸SRb�����n"�_�g�q"[s�J���'�p���M�����Zr���q{8����=Ǒ�Y���N��7ͫ2Y�n"R;���]9��~��%�*҈9㧴���,e��̪��CƓ
5V� @�R�6|����Q�c��d��}��n����αuM��PRCwR��r���$�e8bc�C���lt��"DH��Ig-jȧw�<ݽ�%#�r�t1o�{����)#l��]�Qĵ�ei�lKD�R�2�0�,c�����q7��7	��s#r^$�ԥ�+��60#H��ț,8�e1�39f{m��b9�����UU�|���}���UYw˹�����37]˹��]��33�|���}��u�]u�8�-�v8�q\Uc��<a��O~lY�4w�:uƼ�JJ2Ҽ�N9��.ɭ��H���%�HT�j�t�.�i����ZxiD�H�KV��HT�Q���)��m[n��stT�s�^jxi:�6�6`��f��j�����&�)�Ѩ22v�Z�<$%�cXNJ��$DXy��9:j}�A��^?v����==a�	�0D�b'����_�i�(.�e��U�dI��ʩT]ɦ̓�i����)&˥HÏ��aHY#���0��В���#������	?f�j�ʫ桇��f5����u(5D�҃����|�~���ں�d� ���GDN#<�u�[)��M�	��<܆1Tc���HO|=������9pzHm��%�&��,P]�Cҏ�_��}6g�7cu��Wm�]�Zth��j{~�̗6T.Y�!h�i��Q��K'�m�r���,_t��i��C{��H�N�r�Ddˤ�h�W9�R�WJ�z���u�y��/]���{��ɋ���HH�����u��$�j��]M*N'��s�ܴ2d�(���(��-]�T6n�G=F���E{�M�����l��+�˧9L��!%bU�ª�e���.�6�1�9�$���S��񍱌m����2�����[��[�&L�QcB'`A�%d涒�ϻ����ZE��<==݄K��m�iX���f&��R�4�d{�e���]�6q�eګ-ܳS���[!��Sb��q��s�ӽZ�勵��ۤ�V�ҕ��Ϡ���Cũg�tFl�,POK�6�\_UI.w'1�����rT�j	G`��bUP5\�ܖ�`�=�4z]ꪓ���Zu-�]��:���%Ν��)����SS�#�����JҞ1�Q�W��4�)��v~�~)�x�z���=i�.Ѥ��Q�狥��e稣��ܐ���	�C>�{�}�.'&�m	'��.���T.{
�*3�&�h�C�P�9
1���t��]��2@�H(�Ex��)�3TnI�MC�np�P��<�5;�=��i�U���|Ѱ����m�g	+	�U|�|i{�nB�u��,���``�v4Vd�S�0��d��$IĖ�{�ɗwS!r4@�FJ(��IWk�FX�f)lʳ2��N���Lz�Xh#F[	α7��r''�{�jJ�v�Z��h��iy���q�s�;��A�O>L�8��y��6*�V2v'&Y�QcC��>���f��lU�c>=��.Q��
n�\�GoΤzx�x��m�c�?^�_��n�٪��Bر)�A>����%�m��/�ˉ�l)��B��6���4��]v��,��Ҷ)8�9͍�1��7��ia��U��	q��l��n���4}�E�\��V�e*u�-Hl�A���U�EFM���(�}�^ˇ`���w�
vx�,K�M|ꆆ�Kf��+Uv�J�ٹ�r�aɉ�1�&����OB"z.��%}��d���K)1��ѝ���~��C��m��Th�ק�y̜/}�5L�<���zx�pOf�<��n�ͱ�o4$u��F�]���߇��)4$&��J.�nl���i8m�krI���4���ᇧm�=<x���W���M��ͮ�w���m)�f͝6m���ǧ��q��q�k��m~v�J��l�i�m��ݶ���!T!yZ��HB�b����6����m�M���fݫf���Ox�o���Fح�6l�j�m6�m�p��������ŗ�]�V���?Ӿ���^꜏;����L���R�MvB��6S^Wi=��t��_���V��v�|��t���կ)�y6Tk�.��!A��D�y���	��4Y�u�c{�5u�G�#Ա�����<93�����7yn���N�IeA�,�J�uꕑ�k�,d���%��{m܂��E@�!���n���(�}t��_8������s}O���ff��s}O���ff��s}O���ff��s}O���ff��s}O���ff��s}M��K�I�M8��8�>�k�}+ɑ����*��;�Y�ɭA�>U �rd9��å���n%
Q��� ϲx�Cy��'�n�ʗVs����M�ޡG/��Gæ��!����UUT�T���T��}�N� ���"l�eQ����ۅ��v�N�zkm����\*a������5,�����������DT����!'a��j�Ӧ���d�>~�]ݗu9;¤�3��MJ	�l�q�2Q�F����UUu�p��-N��dg�}go�T?a��Ꚗw�ya�+�Uq��c|ϯO����VI
qd��$���O}d�],�N�Z�r22��s�vݢ0���J6!0��m�������-�w{�2�L�M�M��Ĳ�ww��FI,�"�eZ��b>2p��U��'v��L���ҍ���Z�EZU�����ڪ*��h�c�#Ӑс¡��?�d�*n=δ�K.{�(��,��>s��g���|߂�\����6����-�0j�s���}�r_;R����~c�r].j��P��ĕ�J.YR�Nx~j����l��5�;(�:v\*��ϼ����WиJ�Qg`��ڤ�Z��UwlE����������HK--:~0���iQ��pnN{^�4r�O@�L�۶�\6@��B�"'�]�4�'��ގ&�8�~��)w��\�*� S�,�P~1~!������
'��g%��7�vt��-���Jf�[���Kkq�h�՚�E+W��F�Ըo��nd�l�$�L6c��	�&Hl콓f�y��T��\I��]9d�A����*��?1�m�?_��[+l��5��T��.Ӓǐ�Y��ĭ��N���]3E�sPͪd.٠�8g���U�d4ƞ�.O���-\��!$�sl&=O=P�&''���0�t�m%�L��j���^�m�׵1U�+�UvǬc`}$����6����}]�l릜Ȟ�}^e�%a5��se�%���V�Il�mg&�ծ��,��l���{;4�v��ń䔬��/��4c�t͐K�ܶZKu$�SS;i����{Fcs;q���mJ[����I���a�t`,m2��Np�����c)���N�;�L�!��,�8tL�����j�$������F�:I�-t%SUEE�-?�`ZN�9���d�]�Ϊx�����+�����z��2-<���쎃Q��{=������ʪ�o�t�߶�TR������dz�UT�Y�6<��U�}����>�
`H��K�C�0��,�)���h���:uܙ5��o�^L����uyݫ�b�JV�U�8QE�oߋ�����V]T�v�<�Og�S�5bܰ]�ʍ���ɮ���i��kn��ʓ��d���٤i�b�!NS}&����iN�cKwe��C^�*r\��*V
�E�/أ&�s��W�WU���|�>ʾ۪���<�C	�Bύτ�[�����6�2��n�����Ͽ�9�U���r�����gt�9(�j�.��g�ԩ��.;}��ɔ��ۄ�	�j����;�EL���6�]�x�8�����8���n�;m�l��6m�lxxxxt��8�\���8���m�v�J��e6�m[m��x���Z�!j���R�B�,B�j���o��v۶�i�+f͛6��:x�׍�|��6�lٳfͶ�m��p��������[h���0�q���*����jN�Jm#a暱��1�ײ G�<V*֗2@�#¿�r/���))�	�n�=����g�a[�H1���a���o�"�9�x�A�a�3f@~<�����H��wH���`�S�0��LƭG�m�5a%��sX��7���ۀ=�������.
t�B�K1�G��}�eL��X.���*tnL���#Lj�i�jKNW��_#�6�OlT�&���d�3a!?��p�]�O��s����gH�X4�ƂS�9�LS�0�֞kd��}�쇹��u�z���\W��X��~/�>Pd!<�oR�Yl�&de��p����}ݧZo<����e�B����h�d%��%�$�$Ac ��j)7�\��`%��e�\��;��>k�۫�����Q��dwst3��Nl�N3�2���$c:�7]�s�y��-�@D��2*�F:9���h_��33?�񫹿�>���]��>���]��.���]��}���33}˹���s�뮺���[�QU\R���1�>��h{*��0�T�~ݩu�)�6g�$�Β<��oe��\[�͚�����t$��[e��JL��Izc���L%��GA�V�0�w�����+6�hK5�+��H�8����ܦ��QI'55�3�z$��I�Q�'��4Z^�/j-W���ϨHm�t�$�c�)�ȧ�S�<:w�̌���6jK��*������x����;��DD�؈�(�Et��<�B��K�H?>$�d��K���⯳7�
*z��N�<0���빽��s����p��sƇ�U��ؕB~��h�Tnpm��>,!�����$R�US_�z=�0*l�pj�:	ED`A0Z߿�ʡ�H�ݰm�g�>
-FK�>U��½�*�ɚQ�z���J�����Oۇ�>�o����Nz�V�.�Fꚪ��y���bl�瀿�Y�WĸzL��!��%(���d��K/Q�$��(�.U��͓b"a@�E �����%y��:B���}����{�_��i�B�/$ۖ�$uU7�kCt5w4���C����2Ί�`��J�Ð�NHZEM#l�S-;���2��Q��Тpô��eܴy�95$r�'�EӅ&6�U�a��U�c���vS���q�����,V�%eȕ��I���!q��rr��GD�F�<��IB8etHbxd�����F�kn�����Yb~�=l��$�~I���l`�4�p�h�s�v�+�p��r���gmل�c��q��.*I(�V����G�S�ҏ�I[G���Cܙ��"�-!�뤐�����Kn�����鹕�À�Rj!B'�A?�=	�=$����	"v ���4vqWr��J:d���ý|����}���(����*��Np�<�O�����#q��8�I�9��nd��a��γj�|Ņ�A��j�R���	M��.nQs�]��Tk'-�t�d��b�"X��(�Ex�z��6�RޛU�kX�	����<hZ����T���ʡ_��x(�;��}��\<����c�ʣg�m�B�d��m�7<NK��(tx�*U�⴪u��{%�*z/��N�jX�,�S�|�<�OS���1�Uq��(���Ey��[1��R���:M�7[0'aR�<,~�T���|BI�?s�>��{���)�)��%d�㑆h܎ٳ�U\V����9<v��/&�垌��)�ҎMl���F�UQc)קI��d�V
4�z��1��ӯ���u���r�7�[h��F�*
2*�ҷ6.��̢ɤ�滲���M�X��k%�޴�U3٤�\Z��K�d�Ót��e��^�l\�V$$��E$:v�)]}wn)��,�m):��k�ҡd�{ROYO��p�3H�!FL���U5JP�l ���v;�����u��j�TsWn��-x��it�Ю�I=��p�p�A:B�'DD����~�Υ�x�/��;��0#?L6|�9_17U�R2��p�{*H�.��CiԿe���!鹓�}
>59ee�u���i$��TV��Ǆ.<>�>>/viW��΀�3Y�j���,r���~?;>=z�xӦ�mv�׍��O]�Ҷl�͛q�m====:x�>q����q^���޻m�lٴٵm���m�m���z��aj+T��BՈZ���Z��Z���ݶ�m6�lٳf�۶��m���;v�m6�1�f͛m[|��!˒ԭ/-KR���oժ|���Bi��}�DFQ\x����E$-������<�qsݑ���Vԛ
b��}�%�S������(̦��R�k�c ����s%�2���7�[Dih����"�p2$P?��u�S���x� G�'j�/�bX�zae�^rl<u�?3�T�|51.���2����7=�I'�a������33���t����33=��O.��·˧�wwL��gC��˻��u�]s�e�G0�UW����N\`3�.4R���55�:(��Tfܪ�V�Ǐx�������)mHE�=��e]�8*C)����mۇ��j�X��e��pE+��8�2,��[������]�i�pDMp��8w�#��������~�pχ�c���-��T�B��.ͫeQ���[Ö����z�z�Ej�N��EW���ӑ��70K�ȮL�ԷC�����1�黶q�Y�EĶ-	����.�p��	�B	�DOi3�p��גҕu,���&�?���ň���IU �`�V��hB�V��Z�\�U�6�5,1,I5AJ���;�2r�Tt��t۩j���=�;��K3���ۉ���t�}삆o��YG�ӧa����o�1/Ut0��e�1ӹ!'SV��D4��84��v�J����B���*�1WuJ�*p硹sI���Y���q%]�ѳ��X�����1�m���}���c����5C'��i�g�&��~���4+�/&��vj���<�ȫ)W���~���>�ZK��W�Z�J�q����R3M�=����ڪ�n9<p.���Q���̏U���itvc1��
6QE�l�i\���t\�%�����}6w����Er�TF�|�������i>�Z&�M0cMj�Cr��HՁ;��DM�P�45����nnQ�C_s��ih7�6%�ӆ�ӯ9B�

4B�O�"C���x%��HIh��l۲�ݻ.��6jh&�;�.����q9!TP��3�[�
߄�o�Z+��g���?_ʒ)���d!>d6����a����\6�Sq�n0ê��ʒ��d��@�b��=��=��3j�/�C�Bb���_�g3&hnY&�7�η�|[�+l���s���l�ZZ���8��w��s�Z���MzՐ�޷�k�ܔY`�*�MQT���q/���1^C��O&҃mG��Rl��*��z#!��Wz�Q��\���.��U?j\���S�P���Bөi�EUQT颽���g9m��|)�1⪻Q�(����CmP�'uϼ�^����:������t��bɆ����I0��UJY��I=t�i�jhk�J�i��BʧZ�1V'���>�n���q�Ĳg8���n�7��Ƃ�S�4t�~UW�?1�]�U��fzNitD���s��$�KǞ*��g�g���Ծ]�cb��Ҙ���mce�[��%%��I=��e0�}S���䠩zٳs�':��N�Ӊt���'t��l�`�p�a�C�tDJr�����Ǫ�t��K��&��g�^j�W+k���D�>p��z��'
y�w�WݘV�pɐ��%CG�_���6����	�l�8�y��o{U��t۔�ۥ�$�� ?�?��$�	�}$�I$�UQ(����Q�G��.�	?���[$!�(���PD"l�����\M���"���D�P}`�,"�RE"�)!H�"�Q�*J��J��*J�*J�*K*K��J,����,�(��R2IY$��(��	(����(�H��J((ְ�I`ɖ0Z3#��Qe(�R2(�X��QR�Z,��1H�E�YE��-(��(��k�Qb��T���YE(��*F%(�E�-(�X��*k�EQb�(�E�-(�E��T��,��r0YEJ,QhQE���g���)j����Ԣ�,��Qb�(��(��*FJ,Qb�5,�EQe(��iHĢ�,Qe`�eQb�(�F���(��,��QE(�E�IeQeK(��E�(��)%�YE�QE�(��Qe)%�YEQE�,��(��,RK(��
,��QeQe)%YE�*Qb�(��(�����,QEQb�(��%Qb��"1(��(��(��(��QE$�X��,���QE�*Qb�YE�*QeX��(�E�IeYEX��(�E�(��YE�X���X��,J,RKYE�YE�Y,T�Rʖ	Č1"F	��$�R��b�(�E�X��(��QI-�YE�X��E�ZIb�E�b�(�(�Ж��ee$���UQhZ�T��*��,�J�T�����R�(��R�RQ,)dR��)d��Y)b�)QD�K%,��K%,R�K���%�Y)b�JX���)d�R�D�K�K��R��)d��K
T���JT��Y)b�JX�Y)b�K%(����K�b�J���Y)b�)J%�TR�*)T���K�Q*R�K�K%,��J�X���b�)d��Y)b�JX��Y(�)b�JX�%,R�*�)aD��JTR�,R�,��JR�%���R�b�)b�J-�b��J��ZZU*(�)b�K�R�,��R�YD�R�,��K�R�,�����,R�K�R�,��K��J%�Y)b�JX���R�,��D�X��Y)R��b���A�!�2#dDF�$�"1Q��"#bH1Ȉ��0U*�Y*EJ�V*�V*�,�EX��*�b��b�"0FD�D`��2#
��d�"�b��Q�H�"�dIH���d�H���"�J���%!RR%"ĊE�ĒR*D�RIH�R,"�JEH�IH�T�E�Q"�dE"�)$R,$�XE"�)"��RI�a;�j���+���ք�2R���(kUF1I	EI	=I_�W������o_.�o��'����(Y�|���Ϭ���������,}i�㯆���?_��L�$>��^�	�{�����Q���?��?�]O�|�O��˿�:|UQ?�~?ݿ~�?o���?���?��!�IQ$�#���J�H�?��O��\�������D�A�#�)�	�q���z3������`��$?8�O�"��Ϡ��~�?������?�)C�B��7�/�f'�L�������5��i�k��u�&�}�C�]f|�~k.��,F�?���獲SA ��HT[���.\)QV�
��"F��dA&�tU
Ԙ�|+pJ�6�M����_��g�n>?@Q ����T�-@���'�$�*�$KET����Y����>��d�����H��O�~�� t?�����#����-2�_ZA�*���k@j�e��ԇ����O�}�����}�:��t;����G�����>����0?��?�|B7��}U�9�;���4~��A�UQ>c����?�d?�������s���ҿ��K��?8��'��p�_��8���EZ�}�!�|ɒ��2��!���*(-}RB-��	��S��q��$	�,�'�l	�pr��e%����d"lp�4}�lF�.Y(��\GUY>G�����o�
��;���oֆ>�*����0��"��'���>6��?��_ǝ�8|���|����'��>���
O��>��џ�ܑ��C����G�����tUTO�J�������_��EU@���n���`��ϴ��O����P��܏�*�$`���F���/$!r�C:?�j� ~r��~^��� n�|y�,~9L������0"�����|��?�JJ��'�|���P���a�����_�Ӵ��D��k%����?Ri����>�� �)����9 '�?����>�M�
��]j���Z\�v�4R}g�����+��)T�d��N�_�~?���"�(H'���