BZh91AY&SYPX5�3ߔpy����߰����  a9��w@  @@S@  �  h�I�M�@ 4�<��  PE*�Z�(I@  ��R  
(��(�R�t�@|6	 � � @�      � :�
 ��:���;2�������n�ׇ�]zʻyƻw�^�(���x	�<��;gm]���C�Kww���ݴ��lyW���b�xnK֭�Ht� �o�hPHE� |7������Vƌ�^�Q��"v�P0��N���{m)��Ɛ�=ޒR������ui�CZWw�Ӻ�oA�l=�hr���zピz:R� we)� ������  �p/�Tم��נ^8
��((�ult�A�ۻ� ��֏E��_p�룾��OG&��6C���N���� y�p��( �
/��v�� z���Ut��tWO�@��)EQ�o�pu��}��V@F���4< < Ϧ�` �x4P���N�d0n�n���N���B� W������Gg�l�(_mC׻�7{e*�7�%�                    �  
 J��47�T�F�����   � � jx@��*4�&&�4� �0b��*F����      i�I4J�F� `  24B� �24�S�1&h�P��I��z���"	�R�"h�2i� � d4��0���'���
��e�E�1nZ��z�����?P7� ��� A �ED@~*�����?�,����� ?(t*f��o��O�?�m�x����������? �f����Q@M9��;�ece���� 8?n�0/r��UPҜkDQ����~�?���W�~?K�����u�����Ӯ�̠�*����c�A|zp����hR�e��Zq;�S��M����H�>�A2���	����BFɣ�MA�K&�s�M��/F�Ci����A�"[���T�m�8�M��<kY%К�5�G1�4t��p,�&�+�I���_[SW����DGMV�����Y���B�&��L9���cw*�;����;Sbu���J�����4�D�H���?�"&�W~��֥|�D�O�0j"<䯑��sR�DG�+��ԫM�D�r��p�W#�H��+���W�4=�[ �6Q�%�DG�({��>����R'�"�V9c����ܮ	��Vķ��-e'�+���H�{)����vW��*��E�DM���1�Xhu��>jR&����舺���\����H��lKy);�8ܤ�ze}_v�"i�Nc+��~�';,�g�D�Lѯ��dd��H'7�\�eP��UK��'2'Y�U:rM�7r��o�:���bw�WN�6��CR�H�K5ȝ���ٳ�eh�t8Hl�A��g��U������>�0y6h��H��ep��Md�9�Y:��Rr���<�G"?t��Ï%a�����%P�I�ڪN�I:q�~�A������Șk�Uq������(_�G�*�f�?a�������Gg�adfY�Ƣ�E�|+����N�2	�Uꨬ�+	��]$��}I>һ�P���Ԯ�%Q%�%�%֕	ؔ�I���(A�bIRIrIu$���5ؕ�%o�ZN��G��;G0���Xh�Ih�"��v��lVqW�R$���z�����zo�-�c/��M��5A�H���x�^�n��>I�)����FP���9>�N��ѽQ&�����I��b&}߳����>ĜÊLN6]�D۲sBu�U�nxmd�#�W	gh�	�P�H�9i:��:<)�5f�K��&a��;�ύ���ޒq6&��$~r�aߺ�����o	Ϸp�K�5�D�9��C�ڨm�)�]��$p��M���w���$���&�h駒	�I��N�)���d��L9��GY&C���ņ���_���|�'�r��n�S!>B��C�w�	e%2M$K+I�!�d��>�"%r� ��1!�'1,L�JHO���$L�dN��ɱ+�q�L��'o��GlLK0o	�鲎��d�G>{"t�����P���p�4p�d�96DL����	Boa�'�d�5��H���xJ7�|���H�BlL&$N��d"$���)Φ	'IbV�"a��6Q����N?pM��R"6YC��:'�ؑ47�Y[H��$Å0�N%�Nk�"f$��8N''�l�#0�4���Ĉ��ᢾ�\�"Z"w�?iNRDG�N��n�8ogi��}�$D�d�65���Ĝ�DD�,��L�oI4si3�;%��	�t'�~���iHa�	�t�F�"kI�D������H��w%d�솉�CT%ĉӨ��c�'��0�D�$&I,��a�t{ʉy:&:#&�w:w����	T�>��lF�9��tl/SCz��:�%�E�J��X�.KD�f��D�K4f�+���'~GM��A
A�L�-�w��q4<��Q&5>�>�uEHj|��N'�&Q����ް���
�ᖂ�i�q����h��D���ò�ac���ca���%Cԡ��92�3=ֽ�d�����7���Y�ʙ����Q:n�����S�ɕR%jCGFn�;�Dy�JNmM��R_.a��u���A.]N��L�jYL6:$��DG�������(�j}�F&���".�a3�#*�o�j"ijQ�F���lDYژ#mM�y>Dd�e:�V�"<��g��Z��	&�3�#�TDs�Z�$��jh�؉��P��DFژp�I'��K�DG�����&*�ɱ�"/j&yS�N���>NuR�u�����w�mJ ��#���[ʔ#2�tN�y:h�}U:#{��c؜rHT�Nu>؏5Q{Q0��TD�� ���U(G[���*t�5(�'ȏuQ�T����#@�ม�?cGɟa<:�0vZ��tF%`��TLܣ�x��IL�h�4��e��mK%��hK4�,���f��D��H�5٣�Dș�F��=m&}éW�����ԍ���YTpѱ���kU���OjP��;,�MD�p�y��F�t��5�YDJ5�������䢲C�t���i/mKd�%%�p�4+R����\>�t��,th�����@�:3�Ҹ`�TFK,��iX;�DG�Dw7ڛ5q*ڔkq/�M�]���_���+Ӆ k��|��߉���r/y��{h�D�LDDDW"��{�wͯ#���5�~���I�c�A�κ�񩖤=M5�k�ױ�c^뼈4�1b<R uDz��׈�㨮�V����G�#�{
^=X�G�#�a�'R�:$�Lv�7���W�����ԗ��8�J�E��H���a����QL��IIv�F��{��#V6�o����}<s�!�[��6W�����{ڈ�Tٌ�R�t�ԭ��l�9|����pf�&�Dl)8�&�QṈ�*j<,&�^.�\��<�ac/��z^�=���!�&#b&���h���MG��[��|t.��=z��Wo#�h��	��i�a��J�B5!#Pܡ�{�����enL�VUNwR���䭓M	�H���?�"&�W~��֥|�D�O�0j"<䯓���\ԤG��J���*��r�8ܤE�\4U�H�R&���2DK�̕��e�DKu)�J}>Ϛ����"q�".�a��%|��R%�nV����-e'�+���H�i�N�+���a��e|���h��D۩H��T��a�����ԤM7)��u+��J���MwR�%���k)8^�_v��w),��H��WM�0��g�D�2�O���)�&��'�pJɜeQ"�W\��9�D�:j�NI���U�<���U'd�j����\7%�K4Du,���'|a~rJ���e�,�x�y{"6��o�j�����l���f�+��"9��D��#�vn���<�NTr&��656���L1�:;�RhzH�����!�Ӭ���Sf�D�������t��Y���P��ڪL3Q�� ���$9�9!����g�����׌gh��)�-�8Y4��Ժ�~:�Q �P.��RO�'�Wq�䮵$��I8����J��Jv��R}㡇�%i%�&���Ev�+�q��!�I���9G0����
:g�8���&E0����I���)�}��z�o�q��}�M�$��C+�	�1Ęn�z���<�.�b�"�"��g�
C
�~x��F�����P�q'G0�:&����3����{h�����!�k�"H������G�G�>!��6h$�4Q\��sr�r��7��ٺ)Q'U��Vn��ٵ�ND,���aM�9,��w��a�&�W���V�y�.Mz�+��K��0�b���x�D����8ᲊ=Q޷g�r�'ut����@.��/S� ��:Q��_6��.�����ą��|UF�.un�4���vc�G-�'��R��񃻟+�-}�A�e[��*!�0>�x����m���&,��.��&�P��U+2���S(��V�����W�}p�fC�ɬ�R����TE"���~�n4p�Ύ��I��J�:?u2q��Qå�)�껺ꌻ�q��ݫ�^(����f,�+O2���[l�L(��d|n�3o���7��%;F�r�q���5��Ӭ7"����:h��fB��9������5��A�Tߋ(��a��V�)Bt�U�Sۚ6d(�¨����BaO�e>�#�
}Un��a����tn��R٦�,�J,�!꤭M��C�5��Cy�U�B�v�H����ً��:�TMm��X�1�nT���ڪ[b`����<(�q�pѢNi^G�x�����Ǐ�(�����'���XW�*��H#�5<fe�o��>��)Lc;�a��ㅱ�υ*qӶܰ�G��2}l{��R4.ˣ~>ʆ2�&`�j���	�eTS��Y��{OL�j�i�t� vg�Y����x�ǧ޳g0���7*�#�t�r��:U���Fݏ�:t��b���t�JQ�ﵮԙ	�FW�}�N����@�P��e8d8i��A��{�^qx ���`p��8����ɯ�^qTt>(���0��i�y��&�N��3�)M�t�Jk:=�<<=@8{姆+4t�J,��m��$���拒k�3FS�(��f�ſ��:��7b�Ə��g	,�I*U]��(p�����XS8SHh�F����^0鲎��s��Ɗ6B�.4G���7�Ŧ�Ѣ#]5�EN�>j������xU���&v�Vt���R�@�$�����<�w�����������s�h��r#g��oO���K�CE�6@�M[g�e�:}
#1f��O�ŏ��8�p�����6Y�Df^^��Y�`���
)�H4
O,�@�z{����t���Ιv�"{�2����3\ ?����(����&'����&-�lfz%�Xxx @��t��m��\�v�jJ����8�+_���!�M(G�O}���= Y������r��<���6Wr�(�
%1i]x�31������e��م���pJ�8@��t�ï���L�e��2����Ȋ�\�:x�����"幌�^�2О����Ə��k�^��@���4�� �|����H@�S���B���	���P@__�>zv���wX�Ǫ� U.�� b4�|a鶣�~�S����F�6����Ҏ�|0�k�,�D|�.��<�v����o~+�h!"���)j��ܔ��]�;D�y�R��i�V�b�O��~������'��;4�@�	l��)�����iG.��YL�"�-�м�Yd�i���/]�6p�$�aJc�,�3��sͬ���=�/M:p��� I[�i۷�#g\w����RVs��ֲ���8�o�����J��h��E��ǈ���qe0R��u�i��<h�0���7pP�z�P��k�Nc��t(��q����a[�{Ҋ,�m7w����$WT�+Kׯ�Ox�pLQ��[e�v�\cl���9M��E����E�j龌�O����z���b��v�Y�s���>yZ�YG"��4�Fa�`Ki��>,�e�,3/n�F��D�h�I�9�4]YGe6�2�hj�<pHY���>&����4Ԋ�Kne��{�Uv!�|p�a��H�G,�o8o�y��?|��45t)y�������(�aT(ݷZ�4{br�t�'���)�?(5f��\U�b��7��v��Å]V��6S�p&Q��A3�]���H�j��3v���և(J���&��|�,����+�i��\���_��I7��r�0/��3��ců>��]�<t򏅤�߂��=Y���윶޽,�eQ����S?_�,ۇ㧗��E�7���Y��\���!𨣷����J]A�[Ww�U�N=<_g,�ڏ�E3��'��(�K���$���Iٮ0��K$�B]��Z�K�u1��,��S���f�.�3�ǫ|��3d�[Cj�#g�8�ㄔI���zh}�(�G� �z|3E�.���ċ�_N;��
xpe4�:2>K�Jzt�$����t�K�KxW�4��t������p`z���xA�4Қp��f�w����/e�(�f�8p�ǌ8p���9�uVY�M�y�l�K0����ϛ0���ɠp�p�>v3����7d����fc�K��Y~��x��%�
�j�8h�FS��tRg��7��Q�S/�2�7�jd*�>|�l�ɳ��2��ݐ��z[�Ӧ �����h���I�e��;u�i���o�m�:Xx��8lѲ�KȀ��a^����:�;��Q��P!/f�}�
t�9$� xl:n��D�g��g�8��g��O�P�y�p�kB~��K���	Q�j��tm���f�k��QU������e�<K��<,�eyf>��ܧF�=QR�M6Q��8a�I�l�e֘s!�k%R7�k�ʴ�,���e�<(��N���J^s�>��o+j�S2#gr:(�E�vh�`Y��-;o�\��L&۽
7es�d��]�y�4�����t���>�5��=��	�_V��!�L=Y�XtZ��k�|�I0�G�s=n�|�gI�{\�8���[6�*ޝ7EYפ8Pʻ��Dz���F,ta���3	��3g#Єl��tE��M�v���Ӆ���z����5��4�nь�GU5!�U@��lݗ�@��Ռ,�.�k�;F�$��tMU��-諻��͞>��.�m���dƤj�1܎3N:����\��V�z��2�l��<qҏWT�������yD�y�a�T�1t�r۶��vj�r�F�a���M�s�w�V�4x�3R4o��0�T�@�����U+�U��]:p	��4t���L����W=�a�(�9�~�wP�^��-���pѠ��Rxf(�h�n��M�"ɑ�f:/c�ק����vwֵ$"?G)�6Yʟ�=݌�Fp�ɵGж�5�I�R�d�(����l�g�"�{�r��M�LNd��h���>���M�ƏY����*2q��N��6l��H�6a�ٶ�f�,�*�$�<�G��L<���L71�
��:}0��m��M����~O��>�T��eW��n�>�CUW5X���n+�A��;���9n���I$���(��ו��zX�uL�ٵ��{�o����?�~��+'��g��F����v���?[�A�|�?-��������c��|����/��v3����F�g6���"�F�U\q@��ii��J12�>�H�y  ���i�E��ҧ)8B�p�3�����y�[E��PH2�V�1P��e0<4^sS~9U�R��
4ܮ�'�jى�*X���E���d�'$1e�:1 檨�����{���>neRkn�6���V���[2��d0>׸�ʡ	��dl��}7X�j�.�-v'KT#��כ�{�4&� ��� LZ 2'p����*��Ŏ�Fnl������{M6�y��A$P�!C0��}j`��*,����؋6���e�q��Pi�x��qB!3�:�������	&���wm�����mCv�*� K��ˢ�(�Ѯֈ���V��-Q3��BT����q]�Qsu)D�#^45� V���SƉ�P�{4I�0�A��֎GumE\y[I�=j�&��@CI�*T�WqfҼ'n�6?��Yz�}�j�+��g
�@��QU�2�P��H���r�Nn5�q�Wǫc���T
㭿.�����S�om[�"iȆ�Ѫ3�j-3�E_R�h��2�b��rUHm!ڄ��Xl�c�����ƣ�4����M&�����Ó�.�õ�#�,M�A���ˮүUv������6��z�Ҏ�К�o,w�]�T
[v�� z�6����bJB�׮�ss�U��a�h]����JmQB%����@\G=�7$�%�1���<ĭ�I�$�!�KS���Q��*��Q�o\�N������P�ι��0����@7�E�8x��]��������� �R�)�9���4	aw�X�`8N�-tz ��#a��$EK����@��ǑĄF�f�;��A���Hv�	}p�M1TD���@���r�;A��O�ԞEY��A�=��X;@�<aT	\��X�I�m��'3̦�q�PR�BKHo/\��Ho)I��1Jw'[�����\�6����~��>��o��|ٸ� {ױ�{�Ä<S�y꬜"?8�<'��?���_��wУ�2ߤ�*���~��������w?c�U⮕W��U^*���WJ���U⸊��������1UU�*���U^�*��t�ګ�].1x�UWUUQUU�*��t�ګ�������ZUmU����J�U�Wv���U]�ګj��[Uv�F�U�Ą�����$B���@�� )A!��@P��H�A��S���0PĔ(jK6 m	�O��W��v�j��[UW��U^+�Uڭ��Ux��U⴬U��W*���U\EUUEUW��Ҫ�V�t��V�U�Ɩ�\X���Uv�j�U^,UUX��Ҵ�U�t��եUUEUW�*�iU^;�w�r IJ!$�#@I � �-�H+�J�!J�"�������I��C�^=f�Uq���1UU�*��*���Uڭ���mU�Wj���UҪ��U^+J��b��"���UU�Ҫ�WJ��[UҪ�ZUW���ޭZ��[UҪ�U\b���*�������UWUUQUU�+A�-
QB�D����EH�9&������=�w�<�������Ux�UUŊ�����1UW�J��ZUW��U^+�Uڭ���m��Uv�UWUUQUU�*��iU^+�V�]�J��U\b��T�iU^����*�*��]*�t��V�U��U\X������>
�!�'p��B�d��H4��3lԃ�r@2:�	F�u ((�bd&B��
�09B�қB�@P����ۼM+���|����Q@& d�����g�~?�����h��?B��Y���p��,M��A8"&$��D؉�L6'N	��� � ��ؚD4"hM�8'��0艂`�'D��e�&	
,����t��A4"pN�`��i-%�a�bY�(�6""`�(Ae��0L0NpNY�6Yf��BhJ�Ȑ�`'�$	� ��D�ӧN�:tDě �"P��:"`��t���AAD�j��x��_韛r���"&~l�s�[M�gV�R�����j�ff�����uƚl���1�͖�t��v��uα��uմvXL���k��*�m\����y�Yf�b���m�e�5�.,�!�j۵v���uMA���è�`�١��ʭ�&� uZKLrfi��X�̽���m�*YelFͦ�v3��K�J�]��\�,wYokf�m<ɋq���&�r�IIm����ٌ�ikc�\����inia8�y��2�K-�If�m���9Bz夵��l��L0�QB]F��0eݹ	����7X��V w��>~w�')J�+-���R>U��P�V�GU����Kf������
�n�&6t4�h,+t�v�:�e5k50b��6,�l�R4I�E��@�*-��t�jW7���f��8>�>�In��M{b]x�6
�Q����/)h�^���ǅ� M�D��jUr���ba[j�� �A�����D1���geXfa�b96���,��G4G�+�ԖQ���hD�w%�]M�iG[�,6ʥ���Œ�t��)c��بz�F[]� ��ͣ�#KK7Y/	��e�.Ҏ#j�F�Қ�����\�:FF���P���3��,m��(,�;v���JК�����m�L�@�v���i�V����]u���`h���k3���k6��b�ky5f��ⅷj���pÜ\�BͰX[*$�Z�
B��2ƶ�7c]��a�
kF�*Ķ�#��5	�$m�3�Lo��rOK�]��)��n�+s�4t�5
ְ6AWYK��^&��.����ֺM�f �՗l�kw[�Hy�SQ�-�\l��L��mB�&�KA�m]i�\u�h9����n�,��׶
͵�ѻm1{��B�l�G-��,��0]*��렦3v����gZ�mv[B����W:(��������&ƕ-%�ն��:GV0����	M�lk�c��Y+/^�L7;m��%�+�v�6���v�k���W|U��-�6�-*@�C��TT�Cf�n�ЍZ�t����i[uĶ�1��X<i�)��Cai�i�a֏/dr��*�i��ചEdm�"S(�U~�^,ʲ5W��>IU�HGaЛc��{7����Ɍ��\C&Ip�m�;=��8[�r�	[�6gО_R R$�ĳk�Q��,�CE��SA��ԅZfk�[m-�Ύ�Ŷ��hB�.��p0b��$� v�`� ]Yr��e����
����٪���a&ԕRP�v���ق���K�4��i�rB��Ò]��*X�.��6�4�97hJ������2���av��D+	�[z��-�K�Z��v������p��Vm�P�B�1�d7WO�z>��q��� ���b��I��c�n��v&^�m+n����ɵr�:�ĺR��[���������j$��q51�з*$���mm�VsvA�ie�!T�l6���++D�յC@ё�8u�+��d7�\9����!7 0[[	r�=l�uQ)�����k���n�.��%vhh��m+u�0�-���7g l��8�v�^Pez����m�"�-����KH������A��L���-��d�[�vƚn*Qv�X�md�eHᶂ��[��0d��n)st���� �-4��K��2�\5e�Y��-�:�iiR���\�k��"P1`��B]V����/�:��MH1c5D]�e�-���i	���q,�y���e�MQæĭ�L�dԿ�Z��eO��� ���{�*���V�����}����UW�*��*�wv�>>>���QUUQU���<| Ҫ��UUTUn����!$�h�4�I4�M<pDrD���a�:p���[jk(U�{wM�n��F�4O-@�-��3�c--	�lK�\lMڼ.�u�ZWZ�0I�e�H�)]-uy��� 6T�[5,CsqΤژ�Z�[��5Q�kl��ѭ�si~}�-��x'%���W�)%ġ��Yl5j���B�:�Fк)3(��ؗj=-�-�6X`X��ob�u�C0+�U�f�W6����y��.��kplu��(�ы.���y��:�m��Pum�vc�r�Sǣ��, ]c2a�`��)�/ KJ��_6�;:�$�JZ5�A�R6���(�e��&�2BYX�ѳR�2�n�8�Y��mw�M-	Ճ�JV�ڔ��cZ��v%��Ql�*��r�{74+��C�)�q�E/��^,�q�"��h&0��v�a*�e�w�7p�0�+m��ٵR��xr*�,36��M�-�f)�(���2M۠d�t�н���o"ݏ�C�\���0h��LHX)�-uuiG
 c�g���5d�*����bx�\VYU׭��#�R�<1�k�'�p�`�D�J!uO܈��yHS|ۃ D�yCRp�B�b�����]���tej]��� �)ӹq7��e�A'Esܥ'�~��!�ƌ4%��~���`�F]�Z�κ�׭Z�6$�I��ġ���$G��)��h�w�e�F�J:��"�x��W3�4�Ў�-�c���D�(5�h�{f&P`�G�V�\�����TEM�'%7m����Ib��2"���խ^Z����ai�l�G�0i�&L�R�����GJՌ ��Y',��8"&	�ćD�tᣔKOUk�1�B��,R��� z��i���)&K�X�&���JN`2���Zlgb�8���5bj����6H{j��k����X<BMz���,�xZ�l5��<C��R�'�cL){��3�|�!t�:�ή�F"P���=m��.#h`U_zU���qgr��y�W��EGN̯Hx��,���(駎0L6$:&C����{!Wv-5>� /1>-cF\OSZ�}ƺ�3�t.#���ڶEOk�U,�B�|�4���S�|����~�F�G�4��eq�&i)'j�"H�G�N�Nt�=F>uU���	˺�w��ۆ�x�"���+E�Qkxk���c!�#x�p
�nN��4tх�a�"`�lHtL0���1%0ՙ}�������2�/B�N�v/<9��9/��S6�<!��y��ʪ(:��X'p-dwVI$�����{�MT�Y�L��|Ԫ��ϫ�2e�eت��\N����=��u��]��ߋ;���7\S�3�z���#Oɯ��D��w����Uρ�)��n+>���	Ã�XPk�u��V�1F��d&9+j�j�^/������Ŵb9r��q���0�-���x��%��m4bT9䧭��┣�-��yDE�(7�n�΍�����9��)#�'��͹'�j�TI���[���LC�=\`�2�Ny�7E��pRE��^f�l��f�3O.������箉P]«�Os�m�K��]Qj�t�8"&	�p:&C�
��p������^� �w= �����f�VG
GXD�LVۃ:�]%�F+��KF�i�b�Y�cm��(�{��
�o���vы���t~�ʆ�S1C�� �B`.�C�	6�h����*��c��"�6�!I�!��h��C����9�0Z0a�D�.!����tК8Y��"`�'�Fa�R��a)s0���A/9AS4O�r� w��`�7B:Z;M�Q�Ƅ[���ϒ�nN@�g`th�7����g`m��<�<0�Ͷ�R-G5u�T�m��Բ&��;�DFF�%��ʐ����!l����X�F�2$���-�a�Y�K�V�}�1O�cci�'�@/rb�A*Ѷ���8H�4��4���p���`�:A0�8h����SE�V�rّ��� "8��BNb� U�`I$+�X���I�b"-���+��+.\N�x�ux�����S���è���#1t��i�J�U��J�C-1n�9��z�_�C�%yJ�Y�Çq
.p.r���pn.+�Y̋WR�1�<��Vo0,��Q'I0�N�8"&	�p��tᣳ]j�T�����E���[!������L��x�W�TUH+r�N�5P���ٔ��3�4�����8�tdv�'"�t [\:�:9gMm�K<z)�&>Y2�\��U�w���[�Xw,?^	���B&���Z��5FUe3t�B�)�q�4�����n�SlP��uGR65Z�6�;@p��sь�DD@J�u��E/x~m�D���.������騕Ƽ�Y^ueJ"�ߕ��!xh��L���Ń9m�F�KzuH��� �s3D��Wa��(�T!������\�)�I�a���V�0x�Ǥ��qx��E��J����G,�Ot@���������8���^h]h�2�t�G�	g�8"&	�p���\Qz��_7\�j��t� 2����8j��ЋG�~Zi�jk�z��8��R���I���6 �!�&�TsQ�D��&H��<P�v�J��b(�i�p3f���UQD��@�s��l7z�z�+�&��b�GV�{�"�ܸ�Uzp:����0�CLh���<�2 �?B
�� t?���ñ�p����0���?����$��M�������8D7�f���H�a�4�M��~���v�p~M�*f�������g!�[Lѭ��:�iD�2�(���G�јi�ѝ�� �ĝ����>��Q�$�x�"x��N�6j��p�4(������z?L"h� �G&�i�Ѭ4�:3Gg��ޏN�5�i����,�lj
����~�F�q����i�dzFh��+G�c���4g�!i�0�7�����y����
4��F|�U5��B>GP��=�^DF�O�xG����1�Z<4���	:>��C��tz?G��3H��$l=#����٣��zx�N�g#�,l�zC6���#̨�
#��0􈽦=#�8H�$�|A- ��vv��}�~��@̥�ź�d��Q#
3_!z���e�S�$�)�!��*,������W[���l�f��ݷw��^~b��/M�te��D��� �̭��v��ћ�Xb�5ʥ��ݢ�
�����5;���q̮��۞�pQ{W�h�K�vhN�u��q:Lv�X�W9��녓�V9¬�9�z+�{z��P҄iW�����g{��ә�%���8G�������������UUTUֽw�eW��k333�Ŋ����ֵ�L��efff{رUWWZ֟d��e�f{��O*����kO�!�0х�x��<'���H&(TDA����*���U[z1n�v�#��U��������^)����q�6ݠ����vT��!��#Zw�5�+���t�7�2ǜZ�~�p�tpJzF��#���LC�b�7�	1�`��Z�����7aL��\�p�8�~�,g�p�\�5P>=B�{�fd�|�щ���6HxH�cwc�O���%�р	��ko+5�u�v��/1�n�=�o�鹪���P�&�L-�)L�оɊ�	),a���.����\�KhV3��#�t�⏏�8t�L:i��3ǆt����kl�� �GT��4�M��L!#��v^��x70����$��J��F��"HD�{$!�MC,�5	m6�a�~f��*���11U� �GW�cC�7�^탢���0Ţ���S�+�zf$T����	yLCcr�0͚t�SD,ɷ�{�y��Pu43F�&D?���P�>�ڋ��&�B[d�)�鋀��NM>����v`��A�/$'[p���*�4���O�d�I�p��âsD������<�W���	zM�D��u$�u�64� ��$�O�4��"`�'Ox�$0��y7�4�L1�HG) o#v�PFE�M��3 ���q]��m�J�K�ǚ���Z����X�e�ck��;MI:���m��m�hC~�e�����T7�w�i�zv����kvR+K�Y�����O�
ܺVY�"�K�W�Q{{VV�Y�Ϟj��ѝZ��4�8�meS]j��
�>	ƿ�����p�Y����e��#�3��ǒ����}�f; ܃��8��$c!1�v�z�>�GG�n�F�L4��'�4�F��l;��n��y�`R8rb8B�a����)LR4��Fvn�Uə�URDT�k�;��(
M����f��-#�	�H[��Sl�ܓ���t/�d	�	�I0B��e��GɆK>�A�h<�@�a��oc%Np^2��!�&�M>Hh�$7c �4c�C��@��B�`��+񥣐K�U
��sy%7��wW���3�+�I*(�G>n�\a9AL8���q�;c�{:zC��LtI���M���~	�pDL��!�` St�D�Y.��A$@�f��u�07#�S�]Ui"	$w{��S��.!.bu����Z�[�5
I��n���cr]�����D���]&�w`ܕ� Hс&���{�UW.�SN.�:;�Ց����{ �A�z޶4��gu<�
^��5����y��<��)l#H�CCh-�3�Y���E��%UعE�Y2�qLYV�@�ݎ�׹��o���s!�8f#��L�֌&u���P�X�nJ]�{.nȞ�hN9I��#遡�ƌG�%�p�x��#�,�J ��C4�&�a�l�?��"t���Q���;�_@�gɔ`��A$@"��cʪ�͓�th5&񄼹���MG=��g�{�i/d/��|�ڭ������u�H�	ӬB��y�6�67C�i8��ƀ3G(j�x4�9���b��C=Kx�#@rC�.)�$���8)!�H���B2*������"T�N^I� �����c���������`0��F����f\ �c�p�y{e�j(��N$p�����t��C�l4��
E�H��b�i<=Q����L#�2F�EẢ��(��N�QHi7x;��7z'[Ԙ�P����0��H��uZ�Pa%%�m��k	��h܍��?Q�l�?Q�0DN�~	F:	?LTX��	3�ڙ,z�c0�Qy�6�m6�hK�d�y��b| ��=��A����9H4Ƥ�0$����x0{O��8T���$�2�o��ha#��C1�
:ՓVj�Mi�$�"H)�����t��i�$8H�04�`pH�8k͓d�I����kHL&���;��K������Ҕ�Bi ���A�c�o�3�D�(�M6[�IjH��"�{�&e�s8%O��c��6Yw��K8�&�kH�)4�񇽖&�d���F1��q���� �,�A�t�Nr`�ϼ�>ZZ�m�$����1qt�#F'�!�&$y��������4lF���hO�g�Â"`��:$0��4`��V�_u���Ê�(p�@g���D9"m�Ғ��%�'g�'|GӔ6״�=qj�0Ov;q��)��VP&	~���b
�8�H$�H�.Zu?��ą���w�1i�݃�����t��ز���=X9�@�n.��w�޸7��-�Χw��o3�w��K�v'U�a��7�XE��413�6ւ�u��Z2�;�E�����|���^J�{7�$�J7$��#��ʮO�R�F��to��; ݗc�i!у��1��|qQ�xh�7�I<R�PG;�fd��4��Ä��vEhЛ��G�;a
�J`A�ܚ�ic@t���l�$� g�u�n$r�0u�
 �1�f30�%�X�߽��{�kmױ�=Ň�)x4��d A6�p@H��u����L^�a�Xv���F̼�0a�����b�p�$�!)�f�%�)M��pY���3t��C�D%P���67V���q�B)*2Y(���(֮H"��%ġ��a�
1�J��87M��G�$�K4���ǎ�<x�����H�~���Rɠ�{{DD@@��A��V�����H&[��O��<'��]�7 ���F���(��#8w-Q���r�z|yxMJ=�j-.�|���h��"H��|P�J�D��y�8�x�(,at�i�����K���j���2�Ȁ��t?�`��қI7J3B��	��:o�	���DB���Bpa	0��G�ICC-"�u�Wh�Z��!#��(�Y
�h�0al;!cV.���v,����f!���*JK���i��>8x�㧏0��:t��Hqq���J"�q�b�'�E��m6�m&����}.�����=5���s��&�\n!�J�Hß(K������-Y
+�La��`		�@WE�"
A���y�b�D�s����#��(a��$�.��)�Ա�ȇ���Y�*$�nq{m���D����Y���D
������E��H�D�Q~��k1p�чHL� ��h�gQ7K���M/��E�4���)�	�{��j��a�T���O�.�܎!˂r����8��Ȕx�C:��գ��RQ(�%�e��ۤKC�E��&�x�f�D��!�(æ��2n$���"�21�����6�m6�hA�C�D�B��Fv8�Ѩ��kbF��bF&=,����䗿|��9�쒕����& ��2&(�L�'h�B2��Zѧ:�9i`�i��0�- !Rg	(�J���vA�|����Y"Ks��Wpt�,a�݂J4j#�����q& pk���0';����j�"�����{�)<����~T�5%�
@�`� ,ӄ�a�P4B% ��'�I�ر�_N��MΎ�6&&�n�*��D#�	1� �e#ȕ�2
�)G�R
0k|3�(�!Q�
ψ���8?���������C�4�=�.\�f��4�e�>F�Oh�=�!i��v\��E�O�^5z^�O��^�G�������zlc��Gc�eA�\�����fAѭ�t�<A&�$��-��4~�Ƒ���~L"�!�G��M �D#Fh�z=�"��-F��Hњ3�N�$P�i���Z5�id=��(z9�F�e��M'Fh��4zi8DA��z9�O�#���4g� ��-:G��3�-,�K"F�#���#Dxh�+��â����*����<�,��̣�<-^��X3F`i��K�;���=�.\�f���M��h�i�OCz?G��8i#�T9��A�X�k���#��#D$� "���o:��%�)U'��4�z�&�w��aX���D�����̆t�&�flm}���M���.zB�!Onm���Y�c�k��0f3T�\���TPJ�\��y�E3Z���p��������<ٕ�瓂*%a�nz�b�BGo�wl�}Tm�����KQ�m��U�����AC�z��\��1fN��rQ[Q�p�As~{s�K]�*f������;:���>���1���s.s�wX:;���2���S5�v,U�O�-�KO�L��m3��mFwƻ.�ZkY�_sSjj�̵��޻}��J�8^a�M��_W_K�#\`��Ǩa�P��aĵ�O2�Ӟ��\kt?�5]H�(4�@/���ż�U�A�@�F���Ѻx�lt�*�il��cRS �b�\��_Af=Hl�plַ�j�[��-/j�b�<�615�fH�M�����i`e�2���R!9/t��c�zgJ{�k{�-�l�03s~�ٻ�wg��*�*�Z�쁙�����������稫�kO�fk33=����{�����ִ�'ٙy��������g�yu�i�@a0ц�0���D�:tHa����zǻ1�N4
A�	�=�MSC�1�X���[�4�9�\.%�+mF�L�`��f-t�Ŭ���&rb%�;Im�,�hKb1&R�8ö&�I����J7D<`UQD4�Cƛ��ֵ�5�m.�PKpVu��1,�$>�7��Z�Y1�f�eP.&���Mccv����bR�36.�%���Bj�v֔&�\̌��Y���8Xŭ�cб��o[n�[[)c)��ъر��2�,0�JKeKF��f��I��]�e6���,̺�k�e���Qڗk�ƫ�]�t��5AnF�V���u���3v��2���n�D�]f�lD��P�Iv� �LT�\R�[�x��1�I�)�����|a����(�����̢6*Q��Y������`�k,�ۦ�˘	:��2mBJY��pq6d_�ѥ�Y�^�a��Ы�¶�=��p����MO����R�&dr�?-�Ŕ��RQJd��0�0�(����Z���6�E*��(�R9�ꐡ�L=���G�61��R��SF��(``��^�1,G10��i�CD�BP0�4�Ah87(���,��߬��B\<��uU(z��z|]#zPPо��ur��">9�U�@`h���I6�ͼ�*����tۇc�CbWi9�щ�a��&�,�K����q��T��y��jG��U2���HY�Z�;��*��A��:'p���Z�G�Pc��)�H�����L$��Ϗ�<x�:tHa�:x��d�錃�S(��Ŷ`tc�1&�����X���U��lcGD��@��R�JH�F�xx�1�h��5�n�ACC��2"���j|� �"f��qQNˢ|vM��t�y|�.4p���A��;o��ѕr�ц����cF��k��}�s3�P�f�P��|9-3�ZlA���9M�؛��$����y��3P��h"[oB#����T�������,!U/2F֜$��L.�0 j (�R��qT#�6}(�_F�)0�,!p��o���F��L���]�;$�‥ բQ�=�Х����bGХ0 ��8I�'�Ş>8x�㧏0��:tf`���l�ȆܰO��S��f+d�^FE�ż���pc�1&��ޡ�+���#|��LM�,74a�:$sc�I���l��0���:Dh��P��0��1Y�%���,lv��4���lCP耉t�h$����n�3a!	�0`_o�a؂ZSʒ&e��U26����i�9�ݠ��ې祒9c%��R%s�B�oj�$(5{&�%Hm���$���hݟ]�m��fZ6��6H���"v7����z\�1p�y.��h�b�XH¸�$2���]�<��$Gd;��Q���n��`i�S g���DNQF,D����^0��T�%�"�����]L�
��83i&�<~<"`��:$0�<t��R>f;wue�Ye�a	�M�n�$���Bd�!&A�K&H<��0�B=sߕ�WQ�3�y�����i(���<q0?6�FL���F�30�N�#����ü�gxxGn��16�D���I���;&%q�������3SD⃽n��H}�_gs�S�K���0���@j:'#rgw}��t�8L3ϝ>"�H��H}�r��D���l�6A�)��|�Q��Q(��8�#D) �򤱡��IRp�r� �:��o87c����d�6e0��#bv#c�F��{��xk�(�E���Љ�����&�0��:tf`�;q2y̼F0��K��`�|uZFaNI槼�X�͎��ݘM��7%k� ���Ȋ7�U@D*oD/J1�c�@S)����S���T�E���iѧ�v0�nG���w�δv��'o:��VGӺ�gzcip��2�'7]�Z0:���h��^ٛ�.ʽ�V
��<�e���l=�j��Պ��X����5�������;�ͯ�.�am4TӴ|5�gJ��׮F���y�CR�<4�0�|���m�U����J6���8d�(`0���B�GĖ3P�b �Ѕr@Ɣ!�=��7tp�&��6|��qB��ѢM���������`�|T#�j��L�Cb�E_y@C}5shCi8�1W�\:q���/���J��#	iBa��F�Bm&�tp�#�� ���L�{�jQH�/E" cKP�?�-��VԖ]K����o�n�<�[���\�o�k��ȥa���"�Zjx�)0��
%Do��h�DL����
 ��L$��g��<x��ǌ0�Ν��5�xn�f�m�զ����1�bMQ(��nR��4j�A*��+%�P�L��e�SGR��$�/ /��4�ۯ�Wpګ���5.�����ɬ87�#:���<Z L���n�Wb�é��)2ARd�{��R��5�����gݔ(a�n�,5@Q����v@�\>D��Lp���<��������a��ա� a�w��C�j""	�;���A��Q~~��s�1�M��q-Q(��h�p��Q�D."H��Rys��C|�Ds�}���/q�;)q+taI��P�CD�VB5B��Ơ(�H,����M�����&�ӢC!�����T=q<���1�bM	/�4�I#9k��Լ�,�F+�(	�
.�8i���!�X�SF}�'�mJIFR��o��P�ta�x�T<B5qWT#���*E�&-B�cBU3���9# ����n"f��(�Q�]P�i�(��n�\ �9�N��L �Fj�DIs�X��'�+t'Ħ;������r\��ţQ�B8�۝����s��4��!�%D.�2bI՘�ԚAҏ���t���Z>��0������pٙz���E�����kI2Q����g�08J:J8�-�R�+�1�(h�|����&Y$,���x��~<"`��:$0�<��N68�X�(�厫Y&�4���0������<�L�xlvi7 ����r���?h�~��҈K��%���r:������ݖ����b�~\]YB����|D!(�Q���'/.,�<p,�<w���H�CA
L82���BRP�G�eͱ�Q/FW��ԃbSG\i����D%�Uqcn(o�DD3$�$�,<4���A	g�QItv�if�6�M(A�'��D�ĺ$p�9��~���7��3��Elplrơ(4N1�=��Ń_;��ҝvLc��aF��!��:h�6x�8x�"'N�#F�0|u.X溮�p�o��V-�n��,�%�*�ZN��nJf�z�ElM�(�|wn4cI�BM�p�yOF"�(����/�WZ���O�S�*���2��W�Å�+��^$t�D<���ْ������sx�S�|��	�&�p�9���I�P�ݡs�-Ţn������A�?LqP��^�L�eȍ�����B�'�DM�B#��'�j:'�M�+|a�L�(�h�؈��ml���pƘ�$�Ùz}4�;�#=t��A���ջ����8�)*�k��h�Q ipe[��)d���l�%�������:<u�"0��I�$�HI�"$6IzN��%�X�S.:�6� �b�'m!&&��120���0h��C�M�l
H�^��>P+w]�D|C>uUN��;S55EO�LP����)B.H!|����P����J´��G���<8��h�yAt@��4@��Y��g�?<xL�W�]]B�|����J7Z�mJ�EMU[�Z���c�$З�is��O�)]�z!�8�e�L�U�
H;�H�JJ�lhiZg��a-�"#0�S�<��DL͖��G7>�E�Ebn��A��K.�ӣn]��5����P@Җ�������Q���x�@h\ ��y,��~\K�(aBʕ� j� �IR�(k�E���;�DK��,
$c!6Ҏ/<^fLSs�q�H<�8Ɗ(���jo�<R'p�j<3�K�R��R4><$(a�_+D��D ��i�Yf�&@t�5��D%C�I�Gfp҂Z%e�SG� �84|5E�Q�
�Y�2�#�D?�g�X��zl�#GcӤh��zY�R?�ψ�������>���߇�������h�k̒<�
#A���њ2�Z:�������Fh�kG��ΚAњ?i�:= �O��zx��|F��z|A��h�i�z<F�ǣ�H�H�Hӄi$h�f�G�@�f�G�H�z3K#G��0��c�8C4��4x3K ���;oH��$�4��i:=,������xY=����H���4l��F��x�N�pzr��K#K!Q&�����4�oH��� z2-W�DyXa�h�'��E�nZ8јB���>���<t��#Gc�zY0=4�6�N�G�H���o[~�On7#�,d�S{3B�+�#�<(�(�	܏I�F�rB>*t����6���Nw�����0�,��vU�v��-����c�T����C;n�FКǸ�Y�����b�qnJea��Gaܷ�/$ӄ22<n>������Oڍ\��Y��۩u��j
�^��]�8�+�j3!�bP̒��9��F�$��N�Q�R�<��Ti�gsO�W��\�wި}u�?�sy�o�s��{��ww��w׭i�O�fk33�⴪��{����Z�ffk33�⮕W��^��Z׹�������t��X����^�a,��,��<p��0DN�a���*Tc�BG��2
!ƮE�8��� +gN���:�7��M�N�0��Fd<(�O�	E<S�"����ۣd�9#�Z��A�$�_N���EJ-@YP�}�S�p���d)+������k޾Mv��|�m���A�R��$��9t�$ ���(caC!��N�G��p�ؓ�+�G�l� �D64v�#�̻���r1'2hz�<\��f�6R%0(a�oҋ��5'J��p��M)VI Xõ��gf8`j�)�q29"�}�D�Q	�����Z82ư����Q�ə���3��!5��uP�
0g
,�J>>,�㆚x��ǌ0�Ν��pT0lDL̴�K)���e�f��D�'����(�n�0�6H�A��Q$!���񹸽O�.!5rD}�b��*7'��:�'ȕB."��m�X�0d��*����`cn�<qӄ���p��"LR�%{����-H@H�Bd"�mz%�QJQf�&��S��:2|ڐ�St��1F�B�,�BS#1J�J(�mw��JF��8� g��GN"Ѫ�gS�4�8#w�k���F�Ep�XA��(�G�<if�<xL�`a�:x�w���d5$�g�
o�����ӽ���Uv"��[V]�����Y���'�)�^� ��<R�3�J$�3�PQlQ��n��U��i��i���e�-C�}�*}ΏJ/׽:U=�/�Z�պ6��9Z�VK��|��VMLw]uu�k�acH�L^���]�]�*띜�Tn�5^�1F�,��Z��Ų�6�����a��/0��������W҆��&Q)4f*^R�^P�0��'z��	q�T��<n*'PU��1|����l�È�ԪP1���DG����̜nM�R�#�lcK�#�AG��oG��p����U�V�����Y�!CE�m"i}�k�L��"�W0�r���$1���)N��h��<
W�Qf�R��&U�@P�ޝ����R7l����DP�U�|����5�l��i�:M�#�؈��]j��#C��8����%a4�B������?ç�0DN��ӣ0ӄ6�<b���-6K��AD�y�D}I�yA��� զE�E���2�9+�aè��0�~��Bqґ��#8�����\+�uE/�#�JjW~le�C@bÔ���v��'&1E�Tbra'����^�E"ז"��i�Tq�vו#��B2���7��"�����Qijݤ�������bF�&a��Mh4K��%dDD�����5f}^ipc� �謔Z10!R����Uu�!�v���0�e.#����,��4���0����4Ӧ�<a�ӣ0|6���;(篥瑻�����L��Q�޶�i��x����~WX�ꦊ���ۢ�b>k�!-<�f&3�W�T|�E@8X�8�D	��lw���P��_�O���ӄ&�D ���2��K�h�����`���`l0�Iߧ)�R*iUP����Ť��8��*�u��h��˴�Pi*��8��JN��8B#��#�z�Ӆ���
(Tʔtjq�0��D��80٘�vL���4�9�l�73�'�訴�,Fɹ�I�h� z�Q��@0��x�Op�Ӈ�ç�0���00�<9>�0�ŞF�<&��	H�t��W�fa��f&�OdzI�չ�iu�'W�J�a����1Q����n~^,x�F!-B�z���I��u�l��*�u^���1J0<3�(��<��\)G�_A�4qG�Hf��D��`�AJ6Z!`�'�4+�~��spILBN�=�5���R�(�9D��mp��u�4p�4Q�.�(�
��aC(%Ih��I��nDG8�E!&1��J8i�uB���P�I�K:x��:x���!���{�����r��j)!��8�\f��l��m�U�0�"Qʘ��7�'S{�h7cm�,�q��m���=Ӽt��4�Z��DMv7V�������Lɶů��c1Y�7]1�+��WsBƳ����30Ѧ2�`��O*l�B����y|F�.���Q�]J
�J�BA|/ߍ~��yZ�A��ѥ�>$,f(E�ad��O�u�ρ��*��$��=`���uM�A�m�i�M,��f+F�'L6�����Q�%ߑ��j|��!D�a�K�xV��V3�!�U[����N#x�|D�<�V�#��+�-N��u%���o��'��61�p��0�1����1J�l�-�a��>$��>0�M<i��::3��D�S�'2#+e��Jө�$1�{֛j"�Dh����H+��r��Yk��G�7�O���{�їM����-�9m�s�s�	�����d�wT���a�J!�l}���w��R���nG�EC,��=s5!
��Gy!#c��d��%��%���j'Э|����<a%-�A�W�bⰁ����#(�qw��*�����RrS���鋕�X���p<AdI�OÇ�?4�Ox�4h#�פ������կ��I�Ix B�l���`6�8��*ۻ�.̌��5B�a�
´޴�H��M�&5���Y���SD�l��$8�k�pᎈ%�>7CML dlR�G���o���>�1�AL�%�ͯ���F�1������J/�۷�F���2�A���5ft�p(��Ci��Z�ixq<BBr�7h����	 �i���ᆚi�O0��p��LgG�b�E$�tձ�����QDB d*GN�Y��X� v0�Z>C%a�x�?�(gi��m��"Xۢ�@���Ɂ'��[�ԪȘ�i��.u��tf��gG�B1b=E���uC����C��������SI��~��w�o���O�9h�h�B�cVp�h����V2Q���q�(�܇�sS��F0����DZ ��(�#�2���x��іi������HѳH��;.4��N����EF�#G�/H�����a�ތ�l7�H7�7�pj�#�f�4�mh��h���4f�$/7DkvB�pg� ��O�|a�:?��|Aњ?��.�A�����<C4�h���#O����t=����G:4�:=�����}����i5���њa3A����FB����\> ��;����cg�|ii=�N�N�M"c��i=�F�NN����4g�#G�4�#�Z6Y;�AF�M����9���� � z1���ʬ*�
'ʏ+Fh�'��E���p3F�ѐ/%�����4�::4�3G�6�����za�ޏƐi�٧H7�7�pe�G�փ<��:<2/
#DnO�c$d���';�G�im���"�9y��oF��샚����r��i�`�Ё)�)J'�$i�'��,���k*f�������`�*r������Ϗ��|6�ʿ��ã�X��9�ie�&U���!�r�@���avz�鳣@茄���i;z�t��n�L���жb�r�M�@OTt]F�/Ho�A�mY�|��f66�U�Fc,�M�XGGF;�+�W*'U׆i�}�kvV�&,�zQrꔱQ�@Ӥ�3q]o͙�4��ǅ�T����Qu�Z�J�)ᓫ&�mK�K*�Ǐw�bm���m��ok)qPS-�XyQ���ڨ���H(��	x�G�ƚ��KMuK1JLCG��Y�����F�ı�a�^�AM=s~ײ�=��7tr�K,�}�S� \L6W`3n�-�=Mn�R0��$�d5$o)||�[�뻶�?��������ݥUⴿ��߷�������t��V���߷�������[Uv�/���o333y������Z[���g�a��0���8tᦘi��4��0g�T͖P�[�Hhݪ11��$�s"91e&����4l,5W6�o\���v�R�ki+͹dIv1���Ү-!��4�[�.,�j����v�J%�S-��r@�Sn7;jަ�&{:̗��LŅ�Mb0b�Ԙa�U6Һ�3���`h���B	%`:l�ca.xy6�6��4f�ah�P��1C��jQ�u��5��1ζU��):��d���*�0�ˠu��� L����i���Yqq�&PRѧVVYK���# I4�)�̴q��6G1���K��z�a-"6:̤�0#�i�ͪ��a�;R^u�d�e/j�@�7H#n-��af������L�VVK��Jٹu�"0��G^�C�u6)�W[+K|m6�m6�4-NP�q��.�{ŋ7^�BB"rĪ7����n��wF=L&��Ppf����G�ɐ��b[t.Ձ/	<D��7�C}�umۻ��:�������)�@�Ep�V
��fL�V+�h(d�d2��>�|�FG�^��p���Ö���}"����F�%R�Q�Pc�K:|A�:G� $g���E"HgU�P��۽f40q����1KDޗ��j���k~6��)��C�w�T>9�	E-{!Zק�����c(4J ���M��h�:@Ht�$,���0ᦘi��4��`�.�}3���P�۪ވ7Q������"<)$��"c-������sq�~����jU
��| ��I.��|uM���}ӡR>�PP�Wֺ���8�1X@˂H���a�y�0�;���A�Dl��
o�3%R���^uq\��D+��m��ԛRTPn�{�Z�m�꬞���6?�
_"���1�nJ,���a(~M�aPe���e"W�B�{�������b�p���� �
8I�<|a��x�O`a�8W��h�X�+������j߼m6�l��@ƻe@���B>��:w��Y�����j<�����Ϊ2���FAyn>ؘ��R��A8���E�Z�gz�uܲ�F�s.���wI+�r�7h`�������&~G�&}���/#f���"TFD+#�)f��4��8n�T_�2��8��i��o�X��d��IUN
f	PX�O߼3����֊̚�m{��fgc�2ЇYK��F����2O��i'Ɯ8x��M4�0��p����T�n\b����v���m6�m�Kc�f��#jG�hh�gJ]E�*����%�Rh��vX����`����di�����F`��+X|Iu��V��.t�o�$g��ӆZ%8x��$f�MT��e���Xe��#�-�EH��� >�w���UT���������R��$�OFA����8����Ģ��J8�Z,5t�{/���ŗ�3�`p4$��(�G�4Ӈ�0�M<i��00��*�y��33�u3g��9%u�\0�[P�$(;ƥR�>���䁶�n��WF�KHʠ�m�G/�֛i��x���x>4��\�_�IAE��E��[��85��N�yX�K�����ف�+/�#W��3��`�X3���2=ȼ����b:�|�u�#�с�rG^�����P���(d��t���hk��i���CE�*��,F|��|J�}O�)�n-p�՝)��;��pф�BӦ#�=�}X�a�	^��Bߥ���<�	��JB8TsWT�»7kj��Y�CV�9�WUP�!���Na)C�����g�r��u���Z�-X鈣��,���!%�G�0�8|i��i�M<a�����~bV�+�U�
b��m&k��6�l��@�M~Q�!q� c�m����Oȩ��1��C7�	(Ld��O�N����:��!�D�Uf���o�뵈�  gL<kE��7���H�V=�!#8�2��"U͞&��hZ�<��pn�WܑA2f$�ȣ�hZ�Q����R��X�~��6�3�r��r<z�X�e"��(,a�|�j9��<|�#�)Ht ��(ҍ(��Æ�i��4��`�fc�E7ql��PRudθ���6�m6�4+����m��4�q�GV�z9�t���ܒ�X��n��:�:>����	1ںHӰ��DGPח��,g�f/��F�~oc��Y~ɋ��|����1�gF|�j��Jrq
�(f"K������2U^���|������a#3g""B\ȸB#���ф#��($e�>7�WN��&�
��ǎ�"C�%���(Ҏ�p��i��4�3�[��;��f�H�6�Ո$�H%�����cn�౺��}���B�83�KtR�5~�V߈���i�6�a	C�U�L<�qs��8���a����Fn���4��p��#��	L��a$� (g�]�Bn>GhxU}$�u�]2d�e�g~��q���cgq؎����q��C�K�����)(gJ<Q�<i��4�Oi�1���΂�ܫ㊷��8)7�*lG�!�Z*[�d��0��j�X��	�c���T`�,p�M��M��b	 �	/2�[���C���]j��IA�&a`�f0j�Sxu�nL3�n�[�+��-�q��k*kY&A�Vҵ"�++u��'m(�������H7m�{�aj�8����H ��XR:�Zf�����RR5=��p��|�Ã#���S
��Du{�؎"��鋈��,!oc��3��2(�@�*��Š���ĸ������á�:ڊ��43��aѨ"��f-3�s�
g��\I�
m��q6�iM���v�BMjT�ɪ.���8�P��L:1��p�C��sʒ7�D4y�rצpD%����3H,�J0��O0�4�ƚx��@ځ����32��1d2KK�8�mDA����I(�W����ϻ)ch��`H�l��.�$�HT2�����_� �""9j�Z ����~.��x.xt|�-��L\^�8��L ,g_)C����y"*b@6H�f�(Vj<��^�pV1����פ�a�WQ�Fc�����E�TA'�HX�Q_L8p��#iyG���yi$�bY�Y����%�:"tЂ$�D8"`���8lM�P�!B �"Q]�,M	b&ı8'D�0��0L�:a��8&8hAB"l�O<%�t<x��<%�����'�,K4a�"%�ق\��d��Ȉ�DLb"a�6pؖA,M<I�I��A�[Z4p4��	�ĂpHt鳇	��� ��6&����"'D�6YB �A,�QD<~Y���w�P?�K[�,JZ�W�����M-K6����`|s�*��t5k�j �j�U��n����~z�ivu.x8�F��᱉Q��JY��U%���L��R�j�HO\��ۺ2:�V*ɖ��4��y6Ӽ}�����5�]�k@��5��J������:z����i1�KI!^oa�~��g>N��	뾫�r�6F֐�4����uw*����{�y�Fw��Xzp#��͑�ݛ�Yo7�����wUmUڴ�����337��Z�j�ե�n�י����z�[Uv���ۿk3339���Wj����ۿh�!�a��,�:i��i�M<a���'���-�����m��&�o��&������5�[m>�b�Q�~,�8Oη6���HA�U^�znrc���#N��@�F��/O�?.����^&�T�%���Y�:�q�5qEM��D�|���d�kŢ|�wPȂ
�eB���Gl>�5F�&��Aj!��A'O�P3�|��.0�~~s�P�/~[�F����բ���GIGW���
l:3�I\-|R%A�2�8Ye(���|a��x�Oa�0��eL��h�j��'�i�<�<���	���y&�m��&����{��ՇDā%�g�"$#O�<j ዧ����-5��-!FD��㏾�j547U�Z�;�MG"��S��?+3~�3�h��,�A���Q�tp�I����L��^
���H�����b/�<H1�cc~�Cnb%���nH�5y�c�l��|��I�V�B:n�8`@�9ʎc�B0$���<���c(�R� y����a,�J4��>0�M<i��0��A�/�>u��ʉ�������[�x��9&r�pXF�e�QD��vX�ջLO��A$^����ʿ���aJ��>��wOwK;�����]��/�^�sj����/d�tp�bv�Bm���Zr�Q���R`퀗u�K����==x�-��Z�K��c4GFJ!\E��7=�0�w�����q�Z;=�y�[uk�d83ɣ�M�aD|�M�EA~p�m�]������*I�͛}�|y���Q����f\�Q�2N#���>A�f��>���Ã�>,�<lrs�L7���D�S)��B�#m�6c�q\k�޷&����̏����⤪7�ؐJ<a%�t�4�M4�0�`��s�(BF�h�$�=�i�" ��AjWҵ1�0"��E��`6e�wM�t���mѤ0�	:�_5�LUJ�&���'����#3<�����K��z�0C �����?#S� �m����%�D�-8�Rz����b۾�*&auB�$>�`�u%@`��o�F�uFprb;�WN@aH��t82z�m=ll�W�&��$g(�K0���a��4�ƚx��^&��Ι��bJ
��&��rJ` b�����m��&�)��ss��F�(���8��<H�h��Q'�}�+F)Fj1G����"���cG�(z�4 ��g�暸Sh(�Y]e�6�mL����ξQ��Rj�e�����$��qZ������y΢vW��0�A�Ƽ���L�
O�>R%w��ĲX��*Қ��u:�j���8�\8̅����3�Y%�(馘|a��i�M<a�������/��Q-2���#��4�M�����PZ�a\��, ��y��Dt���V����YG*U؂�)�?�r1�c1�b�.���\���0(��O�ʿ"Q�@`�oHD#���>�)�GEu>�JP#y�����d>#�w�g�����������D����<�	-�Z���A'�w��È#�X��DGit֎"F2�6�����`p��Ag	,ҏ>0��4�ƚx��^���7%��J+��x�ɖ���e���h�uVM��6iKS��di������ʅ+����m��&�ߋ�]͏�z����s&���[�L������<܇�#[2��}��/NU��(��fޚ��N�hチm�*�깚f4B�r �%��H%�Ҏ`�Ȉ0�����v�Gë
���8��o�8�%�ޔb�P}���|5j��IT6�PR< bp��>F��{�����qT��$U�V�u�4�=\-uH`urE�0�@AE.h�d/�}�ۂ b��hQ�ZR�`��%��dx�ؘ���o�|�ڂ��=�2��y� !||>����ʿ�5a&��c	$fp�K4�Ǎ0��4�ƚx��=�Gf<�h�����)�[��D�.֒��å�,Ԓ��7����U�羗�Ĺ��r|�q%	qOR�K'b��L��2"�A��>\C��:��E���B	#>ESv�>T2�Yѩ��0ߖ-��{�u���-�1�T�"[��µ.KIF�wD*�+���V{� �{����j0�a�,�J1�����$˧ɂe`a�Q�F4�;1��	@D@� �I,|a��i�M<a��*slq,��*.�A$A%���q#�������J8�A򂑋��L$��W�+`��sRx�i�����Cm1���'��(,�%&��$ ̋S?��n�qSP�ƱB��^/E��S�6�Q�\-0���Tp�	R�0�iQ��Dy����nu��'� �6s�a�UL6JUN�?�0�0����WL��gYIgJ>:i��a��x�Oa�0��*oڏq��8�3cAP�,�1և�*G[|�"�"!{�i����0o�Q�KÁ ��kMM�_)8��u����O���×r��=ײA�Ė��f3Dl1:}൴��d�uSg#x��Z�>6�5h��\������0EJ����^����� �K:x��feDA�c��N�I��yI��98u�M%�x���Q:�}��">F����4<1���J�h�]:YD���Ŗ~ �"&�DD�N� �D�8"`�鳆�(ACB ��Q�,M	b&�N�`�pâtD�0N��M�Ή�e�DK:"&Q��К<l���<'�<_	��ĳGMAB"'L4 �Kb"tN�&�DÂl�,�YBhJ��(��'�tD�
JBA!� �0ÇN�<xO(A�f	���"'G�؛4P� � ��B�{�O���D��A�]�n�U����q����h�:ޖ��V᷎�f���D��U���aįrTˌ����۪sS�x���*"
��X.�9��^�֝��<��7i߻*���$~�8�`e�ۃ9����Mz�2�ci�!��L� חgf4���M�Н���v��9T�ВU3K�������V���L37s6��jўr/Y?î�R�T�A"��|���>A$�q*9�<�1���2�	�3΅j��6ܠ��2��IX܂�MkWv"0��[R�Ւ$�$�Q�
Hm�4M���Ri�Hu>��8�V�h����ˁP�[x墭��ѭQ��mj�.�W�L��JKIo�yjQ�,����oX/�����]c��Ќ-���JBTkVb�("����l�y�h�ﳺ�w���SYǼqҪ�V�t���ߵ�����{J��[U�w�ߵ�����{J��[U�w~�Q�����{J��[U�w~�W�C
0�F�,�<t馚x�Oa�0���� �K����~�L�6��V��DZ9	�m�v�l��x,
�ZJ���R��m��Yo\�e5��R�s�\�ok�cMV;,i�0�F�va�����8�kv�ǎ*�SK���˜P� ���TUV���-���U
�D#�.�nѡ�F،˄r��k���b�^��n	�J^�H�Kb\a�ե���!��kt�@J���m�\;��|h>󅫭9v)�J|mi���_FYeas�.ڶC2�a��q�����63e�-T6���+K+�GJ�m2-yq�,7�CǗ�f��!�P֚M�ٔ�Ɨ�	�e�Fڄ�yK��5��!{S��%�ef�E��B��G8��"��X,�z�H$�K�v���/�⚱ǋ���Ws�!�+{��ʨ��wXs3���{�T�ݕ�N���*k��;��ڱt�v �w[���5�z%Ӥ|�p�5�0ul��s5b�Y�<V�ձJ��$Tb;��{�(_�����,2D��֏�Wk��@Ə�#8X/Sm: �Qb��2g*��a�����K���A5�w�F�3����3/���4q�^�C��̳���m��\�C���X@p���_�ܧ��8_ؽi ڴ�B�A�F�]]�G���Ϛ;�艟pcϐÇ�I�$��x��i��4�38z+�3_8Cd�2��Z�������2�VZrϏըfa��f&���hb��0�>�5�6�1a��H�!4凛g& g�	ki%���Ȗx��㈄y�u��K& ���+�C���hY��_ˈ��d��rꦩ{[:s���X|���>>(aE#>0�q4���PQ`��SN����� ��|����r$�g�3�t��
4���:i��4���s;v�!m��V
�Ty$A$^ӑ���3P�����_$���:gU�[M� ��Ԙq|�)	J�9z�|Z~7����S�p���{(g�BH�����pz����Q#�-�aeNH�D�i�|�t�hR�� �����{h(��(���RQ�HI9޶�'�)4�YA�tm�߭�ܽ���ݺ�E��kz����'G������|1I4�(g<t��
4���t�Oi�38NzQ��0ۈarE�Zm����ò1��wq�*ˤļ�R�ک�A�At6�ҿy�uR���0�{Zu#�O��H�8M�o�	wf!TE/]�m�O5W	�l��h�xZ�G��t�A�[oQ}r�E���}��
�s���p�]��ݲ�#�-ٕU�]UGt�,D�{� ,QAÂ��㯖(Gl�Lh�"Bχ��~����tR��y����$Ӆ<i�Ƙt�Oi�L�G�Bs��X����P�U�%i�����{6���i~=��p�Z��s0K���X8go�˦�l�K�
���7��q�r�U���,k�gns}k&v5PV�"3���哶α������Y�S�^����ޮC*�,�㎭���nRɎ�1��R0W�Ǆ�_Cu��!���[Gj�]9���ҍ��c{�:u��=��\7k���hƺQ��\��U������8�R8i���6��ۙ���;��OH�7)����+X`Y�˜E�A`u^��[g[Mx<AgW�n�w"Â�G!�b1{���D50 �n���b>��ߘ�V`� �d�I��ǌ4Ӧi�M<a�a��cy$$ٱ%d��K��'�3�30��Ç���$�[-���Iᴬ�ӏ)���uVc��gI�z�LGR��xJB����4��qRK��+�Z�"�J0�I(���P�Q�x��nO��+�a�8�%������F�]���f�ļƈ�cf.�H� ��q�-����qS#���D,%R���h���<@�0�Q���2�F`p�� 鄜$�O|i�4�0�0���aF���<A$A%����T�M������p%D���IR+Gh�J�Q�'��s��N�l�e#�$%�~���˞��H'	$	��Z�!�8����iHh�Ǟ��4��(Xjэ�[���$��(GO�������4$��z'�N8��N�q5LGL*���<q��+��R<�b:x�4Z<b/��3Y�	0�����tӦ�4��:38�Z HCb
�w���qD"
S�"�,����₊A�}B2g14%�yW>yF�#Tu�ہ̐�;�.���0_�_j�]Va��6I�e�fF��A�ٿh(��JȃE�>P�Qam������Q�40��z �dG��؈��	�ag�U����5��u�⃤qp���D1�c#�X`|4j<�p��:J�f����3�Y'�8x�L>4�M<i��:tfp�Kܯ`V��"vk.��'��<j�̪���Q�" 7��P0U�)�I�7kb�W�h���$�H$�b������|7h����pmf&���e+z��9ۈ�r��;]�.��Aq�J�c&���1-�������V8��9O��,0tUW����z������'�Q�۳P�`�ט�._*7�U�+#�x��&���0��ƶ���U�i��(��Qަ�BR�h�r/K�Ԛﾑ�1��±�lţ���z`R��ȟqv h�]�=��m��#U"�&qӨ_��8���J��L�|�I/-q^�t?[�N.�:����6�,f�a��$醚a�M0�ƚxçDra�lo�HU,[˖k9�cn� ��"�D�Q�4�_�R�":�<b�<.�.g�~wwuT�Ò��KmA�G
�,k�
N^(�tJ�o�.CV`̅\�A%��M�S����p~��s�յ*Ӟ,C9E�[��D6/��t�qS����LUqH���#�Hnm��1 �V��>L�
�Fj�)È�|��pӄ�$؛,�e�~��"X���'JD�X��:tL:lD��(AA6 ��Qf�BhD؉�:u��f	�`�&	�`�!�4tN�(D�"X����Y0J(M�'�|i��<i��i&i��	,��&�:"t�� ��&	��:&�͉bY��4%	BP�A��� �(M	N ����gN0��!�ǋ< �0DD�6&� � �'�!M�G���`�D��Y�����6ɸ��[������u\�Yqnnf��*�!�t�li�JMW]꘷n_`R3���A�	Iu�cn��h;����;[�c�'�j�4��׆�K��C���f��]��j��hbܜ{s��-N���&+C�\����,�xK|]K���v���Μm�e���k�AJ����ʫ�t����oՙ����z�U�Un���Vfffg}�UW��U���zffffwޥUx��[�����a�0��	:I��a��4�Oi���q�;cM��M�O��̸��t�=�D̐g����.���4`�.���}�qt�C6��|���2eU�=@�u_w�����}�b�6Ϛp������͍�g���W
����їd7$�a�PÊ<#����g}}�'@��1njS�x�2��>D�@�kzt�Q��+#�C[
|Z��ޅ3H��I�Oi�t�<i��:tf�������%��e�FB��Px���њ)�s��M��Q�E�c�ё�DuI��Ջ��4�j��b9�6F*~�s³�""��D�����K��=G��ժ��ѝo�+��D��1�;��h���,ӡ"��G�.��C���L����V�][�]Uڿþ�~�}|�����fZ>GD��#�!�Β�G����a<[���*�2M8��#��I�&�i�Ɲ4�Oi���q�m0T�/�.�U`�WF��Rm���A5�pF�8Ԫ�^�Ec�������:݈eТؾ.���\��I�Ix}�{�卪��u�F��8�ϯm|9�ܾ�(�몥L�Rf�^��뺪�d�hF��m^�W��Q���o<�$32��L9u�:�1j��#&@z�cxh�!�;ȧ�A5�YN�:�K�n=f/"����֜�W��GB陱9�˟^,�5'���;�pȘ���q�sW�%ܤq��)�X5pj�ì00�q{4ƌF����ρ���2; �U��i��}� �����Q Ϥ8��ѯ�p�J����®L4x��0N���<p�<'L0���/���L��(11|�{Z�,��i��i������@��/�w���z�4��dV��LȢ�5{��>����_w:�s��2�FG�Z��Z�{����5�<p8v�D/�H��&zd�"��#� ��+ȗ�b>�����=�đR�7͟(�-�וQ�bvd�{�&-�JqG�uD�`qp+�7ўm�ώ� ����v��J)u���SzI��i��4馘x|>0h�F�dҦ��J�=��H6�o� �?���`Ǝ�8��F ֵ�1CIy>�Lx�
N(7n"�G���Q-P?6)B:��V�4����	E$�?�i"�G�D�|�2\DT#��a�`�^GH&_+G~�º:*"ш��|�
���lah�Q+Yӧ>��PB�'2k��<�XΑ��I�O�>0�N�i��4�N�hVM̉_H0Tj
a�Tt�>1DAgN��� p��0!^#˯S!j�W�%�����4�/�j����y���m��.��6����+8�`���p ϑ�}leZB-�m'H�!>Qgh�q�!����e�D1���>P���\���SQ�K|u��'�D/CZ�M>L�ψ㡋���U����$��"��'Ěi��t�L<i��:tgH�z��q�0O2@ƹ-T�5��MkN	�YG Z����x�DR@�ئ6��i.��4h�����r���Sn�V
8�0ZG���	 ��ו�����ƫ	��f��RuP�zo�]�ޥ���}���:�,��4�޶�,�9@�v��dc}�2��e�gaW�a^���i�֖r]K[uwUM �2���F�Ft�����b���i����%刂��F�  ��:�|�%v��s9��l#Q��񍺟���ςU�C��%#�7b���N�]]Z���H�&",$$Շ!�5Nb���>A�m�62Ⱦ$�YW;|9vO8�}�I��)�>��Rh����Y#8F7��a�O�>4馘x�Ot�Α��k��`�qU5%:dD�7DDB)�ag�X�#1Bkģ�M&�ᰣ��}��g�jׁ���RT��˚���`���c|�h���uGxa0��Ǧv�t�����j��}�y&u��a��|�96�Jf��zm���U�8�3qs�WԡRj���7�R<�^�gC�a��9�Q|K�Lc���H�K��BK�7��I���t�L<i��:tgB�fcY�:�ͥ�-z�"ի0 �F:�o{Zm��m����D9���gE(��h���]"�}$+丮�^]/H�Z ߛm��8Bp_+3�oT;��BY�sV{��G����Z�����~�V/�8Bh'���ϾE#�y��BjQ(�Q&"8��RS���wÈ<[M��y6��"8#Q���Ѣ(w|8t�ͺ�֎3�`��J4ӧ�i�M0�0�ѝ#�Q�t�e�9�&a�)���;�֛i��x�/qUQ��SÈ��z�!?������|�b�GQCq589d1���Z!/)�1�*���ul��|��O����7��:E'�����{��:|�aA�� �몰I�҉�4�]ӈ�,�#��+Ǭ��j�������6!u*G#��9�������Іz�5��������e�iC4<xb"&�DL�"A,DD:&��6&�٢�AA�F��&�M���a�a�â&	�`�DMa!�:p���"""'JI�MB%�������7���Y�"hDDL�	��DK�pD�:&:'N�hBP�%���O�D���АD�hD�t�ӧ�'
D�'�<x��	��"t��bl�B �!�p�> ��x�J��6g���w�2�]�hT7m��mH�� �TɎhRT�l�x��^�],uxrQ��,�y�O�*m��}/��6c���N�'j��3�|��,]UU)[F�͝���B��Ru`�>�s�h}J���T𸛩m���v�&�w��S�c�ax^v_,��N��S�+�쨲(j�̔�c%��Un��vvʻ�����g:g!{u�221:��eMDu��wP!6_�y��5݋w�-�H��a�.��x��3���p���ɝk&M�d�#��ӳR�8�\����(�E�_]f49�&�Ø}5���/-X���-�w|K����	�eM~��즛jk�8��@�-v����U�7Zv�0-���U�e���67����RV]���B:Y���}}�OĚQN���6\mh�G%@��+�`�
�7��������EU^�*�ww��L����g���V�[����fffg��UW�J����������z*��iU����|a�0�F0�<'O0��|>0h�F���1��h�8��/܅if�V�45.
�ב���4��eqgu��ݴ�f�r��K�v]P���Ҽ�3K1k#KH;k��b� �k6�c�TA�k#�h��n��&-u-�LǨk
��k�P��s��5�b�7g�vMys�ml`@%�+�8c���4�uږW )J��S`~|�����*�4x-�y���Z*V��^#ՅP��h�s3w$1	M-�.�3h�4�LB���.��)bSB�&i
5��η�.�h=�t)Ny����4��f�%&j�^�ѥ�7h��m8u�^:�b�mZ6�b�m��-!� ���3U��jY���!�Xk4T��5\A%���M��M�D㿟���j��<FnG~/����w�^�tڱ*p83:��5�W\(p7��A`��T��N����V���ʿS+tkCl���	t�
4�/-��A�6�{.�L{�XQV,�GIH/4,� �Dqa��ے֖~�E�l�p##�Q��&b�
�������˗3)�{�w��(ak��Gz�+OA����j�jJ>G� ԡ6�.̳�сB�����G���O]QԠ�Qs��$\r+�[##Zh�٪��)KHX����(�Z�1'��C>]D�p��,��L(����i�M8x�Ot�Μ$�㶩�XM�n�t(�1{�F1�s����k�|�B)�lZ�ˊ�g�+�nc驙 �5�|���p��kaF���Z �<Z2�7A g���Ě�JZy\��̄����	&<5��6�߱)�j��F����qo���A�,���b>E��p<6��ێ"��G�PI��:^���5a���<�'!�J(e��3�t�J4�i�M,�0�ѝ8I��=�r�����Q,VزL�2<_z @���'$��p��_Z��������#�|m����R�X�)hz��-R��/,f�"���0ux�� ��Y��7�Z��c��Qg�GIm}$q�ӈ�yu}�q�\AIOí4�Ʋ���]k��p��S�Оax�4|,�OHYÇ��I,��p��M4��M<aӣ:p���]�E27wU+� BOG� A���_�u.����(��<B)G��a©�?����`��&�Z5��:*�iM����v�lc�G�E(]���+C�m�ߗ����M�$�1u�I!֙>���8raB:��B;m��p�-vR~�����a:H2�^=�I��F�&�ӧ��3%b0>-��`p38��:� g�I>$��p�M:i��4��:3�	"w=%�>���$�Q����+��]*i��:*��m�˨ǎ�`˺*Z �H�V�BFJʝC�v*d��_.�>b1	hg������ŦG&�f��J��=�a1����$��pn���T+�����[I�:$4�=���ѽ��v����it`!�T�(��ss4�ν�id�]E�����*���Z�����p4Rs�7��~Dϛd����i����-]��2WY�oNZ?EY�'eu�C!�� �:v�+�88x<4��� ň��>n1#�0�K��4��aG	j��+ ԑO��URt�O8bc�����r;���L�(�O�%���L$�G�O�>4馞8i��:tgN;&�1�U��kq�9��?� A�Պ��l0~aH����u6�QJ�!��u:��m��b-/2�#�#x�K��WU��-}�B(�oC�JGR���f_d�dr
�,��)E,��m��gI��5�����DDb{�b�{�Ye�j�(��b㴤�w�"D%�8^^G`�)4i�yX���rE���=w��a&�",hb�8Y�����	�Ǆ�Æ�K[Ff-!��^mj�UF�]�QE'F���ӎΌ/s����lc3��G�g�ǉF"1^
P�v�l�f"�Lh(��)}ӯ�j�A�&?��w#��ܧ�����(��ԟ6um�� h�t(�U��:�'s��+��61:L};yȆ��b����Y��O��� �����a�d�d�$>4��4�<xN�a8h��+'nU]kFd$E@bW���|�m�DY�����XR�l�����dUUESp8&])���L�.����Q�QH����QH�  �Xb�*C�4Xb0^�(�8NO\4_�j�ck��WCl���a�1>�f&X��,����F�iM�2�~W�6�x�L�{=xOCw�(Jx��NMsm����ӄ���-Z0��bp8/��餖I:i�M4馞4᧌:h#F%�Ƥ�HEv�1�]�uNS��S^͍��R��u���ݶ�86����H�T�e���"��X�lnn�� @��C����O�i���5+�!��~㩕�:)�:������69Մi�`��iT�����t�wph�v���"�a��"�G��ǉ&�J(�mF�>�{�&+Ѝ��_��8�<HX��"(T�\�6�"57Ry���L̓270��uv(��{>y4t�gX��8�,:U�}�o��T� %qO�S2��u��HEM�&��:�ٷj95�>�ޅ�|��8�&���+X�h2a�L$�GM4��4�Ɯ4�N�鄛�߰��Ğlllm������d��yq�x�b'���C��C����1��l_PHy`/B�MT��,R�n�E�X`4B:��"�p ���ba�d�?G�����s�GIF#�����}'R%u:�l�RZ�2�6�ҩ�#X�1�ȅ� ��� �>���ԣ�($�=k�1�8x���gM�&�!�Ab"&	�D؉���6&� � �"C�hCF��Љ��q��&�0L�0LDL:A:t��,��"%M	��&�pK��bl�Ŝ!�ǏnO0N �%�bpN�""tÂa��	�e�BP�FO��>A�JBA����N�:t艂p�D�6"tD�<`���<l�G��� �$<x �����k.��k�$}�]^�Ax���`B(�oz��%kNY��أI�Q��c0�x�U�meN(��:���r̤u���^Wb)�B�e�2�������yL����z��������SY�Ƭ�@��O�b'DsD�<�C1t��A�Ij+�t�G�uV����EL�"��a��Aд��FͥkZ��5�a&}���ٝ�1��(�TP3y(e鬖F��w�ǵ/�(VQ{�y��*��iU����fffg����1U����fffg����1U����fffg����1U�����ѝ:I�N�t�4Ӧ�xӆ�0�ѝ0��[G����Ȉ��"d���E.��q���GQÑ)�
'"#U�o�0���DE =`}��)���7��d$�5?61�t�ȲH\b���J���Qjr����^G�yyj8�ut(��!��=虙%�F�:��u�0�
��Gf+o*:�4b���!�hK0����	�g��P��Q^���z�ѓu�My%�� m�D�9���'������{�A��h;A�2$�|�X%�9�iI��Qj�G6`��<B�=_TC�
h$��֣�Tߩ�a�����1�[��Ԣ�X��;��1�FKo��x���PI�m��<E�!"�N�G�M�}��ƺ�p^Mb�Z^D(gNp���	���	�!�M��cO"-q�u�Cf���8�ۙ�n�伙�rb�S�~
["<�T��{B�i�F���V�)���Z<I$�y�쿰WG���>4�v�U�ժ�S��}��gwu��.��f$PɻJ�:��:�µ�5��FR�紵]J����T�$s��Ӕ3k�9�P]T��T��UIJQry*� ~����>K�#��m��(�s�������zO��|�Cۗ3�9�L��E2na�U�p:���#��}
��LS��3��Lu�xs����1��{��Kh��$��h@��+׈��u��IɁ�8H�4��0��O�xӦ�x��<aӣ:a+�}��ƒ�A.���Í ��bؾ� $fj�.�\�J�ٹ5�Ƌh*ꨇS�1��&���-�~Z��;�q1.���YЄR��x��A�z!8Dw�&"7��,��W��% ���0\��^�>6�&16)?�+v��Un�w�:���{���z޶������#���Ckh\k�^�<6~h��<�:A��G��ğaG��><i�M<if�:`�8I���'Z���"$�1�DM:���m��ٌm�����lS\\8�t�#�x��&6�|R�w���yqb�)d��vf���Ev]ߛ������%���x��{�*��n�cE��#5�F�.�D�Qh�{�޵�i��q��L�l``6�O��i�"LC,�\�(8Hϊ$�D�N�<'�����EkȚ�&�{���  ���7���� ө��IgN���d��l|b=տ�����w��[�F�T��l]�ȪޢL-4y�-Vtf�h·H_Q���~���lⅫŢ[�ll��"	X}~��G2�$q�K��,|QWP��KVyD�(t��Ֆ�Q�ނ`�0�v�3$5�{�)h��A#:|I��(��Nx�ƚx�1��,1�W �q�)ՕE���5�pX2O_4|�[�25+&6}�go\�齵�f8�G"�bE�I$����C�ߍP�3��}h�!��ہ"w�-E���s���`y���Yl.������E����`�i�n��D�U�K	��9}�X0���󯜍�
Ւi�S3����?<��@��"�(t��q|�-=�^&��ч�[�W�)��'��a�]�e����5n�T���W`Eå.����F�Œl����G�Is2�5q�u-$��B����0��:����3��܎8�sst��Rx�B8ypFY��\,f$�M(��Ӈǌ<i��$�L�	��&H�DC-��ߌ qT7�r�{�7��:<E�ain�ޣ��#��ؒ��,��!+��@��B�'��m��G�!Ia(�:����-LD1���(���:6�x�<o}�ᣆ!4
A����u*�NU�-6��J%<k:���_�E���7h��Ξ%J�<�a�$�G�ᆥ0�:������ o�̐�܋��D:l��G?��<Q��0f$�x7������q�h�s�(��(MM6�Fbإ��� ���!�4�&в��� ۉ�8��D�#�R!̹6�J�<t�!H�b�kJ-�-'�٥���G�����c����~��	!, �&1���FB�A5�S����W��a%4�"-i]�t��p�X�.)H��l8�& ����:��g��B0��N�[�D�U�2�$�:'���tD�(��!ӆ��'ӗR�\��Ť�� ��qx��,�1����1&a�=j/�o(�����pq�qy��b��OPf��>n""�H-Z,�y�����,�o�����^Dc�"�j5D��D8�qy�m��,�/a;����]�����8듗 ��>_h���>���$��((*��aP?����~�?jt쟴��'�?�Ѣ;qÜ@ArQqM��?���4ÿ�[�(D�	���
i�bH�f �&"	��p&���	�Ba�f��&	��&	�bb`�B`�f	�&	!�$����$�H�$����$�"H��D�DIĐI LDL���LDI�DDđ$B�DLDI�$,1$DIDL,D�D�ID�0�D$ PL3L2�D�$A��KDD�	$@D�ID���D�$ADDD��D�I�DB�D$DKDB�KD�$I$DDLDDI��ID�,DLA$ADD�,DK��KDD�,I��$DDI�DD���,DK�D���D�ID�,D,�@D$DDI��K�D�,DK,DK�D�	,DK�D��D$LDLDI$D@DD�,K1$A0LDB��A11ID��LAD$ADD��LDLB�DLDDD�$$ADD�IB�D�1,DD��DD�1$DL0PD�D�0P�D�D�D�B�F��H�$�"H�$��	""b �	���$���b 	��H��	"b"b�"	"X�X���b"b �"b ����$�!��a	 !��&"`�	 5�C$2@C$C$D���D���IL0�I�I��I�II�$BA$2C0��I`000002! @��0��"�d	�2�	(@�0�!"��0�&"@�?�8	 @��0$�*@����Lb �&!`7�7�G� dH�� a��``IB��@+"��@�02!�	�02	(�0�
0	2�(�2���@$(@Ȱ0�+
�°2,� �d)��2 2(��02,)�P&�`aHF  aVT��`eH��j�RE��`dHFE�� dX���XHR dRA eBQ d  2�RBQ %Q %U !R` E$VE $	T  XF $P$,����J@B0��@B0, @J�Hd���!��2$0����0�2$0$2�Ȑ��C"B��Ȑ���+��2$2�0)
CC(C+��0�0�0$0�)C(C+�0�20���� C
K�&C���1d�1��C�C$1����),1��1��2C�
D2C$1��1��@lB�C�C�C$0C)�2C���B���2��2���)2C�C�C�
D20�2��CC$)2���0�C,)2C�C,1��1
IC,2��C,1��C,1����2C2B�C$0C$0C$2�$0C$�B�C$1��3C0�3
D2C�1��2C�0�������I �A0DA0IA$�LA$��AAL�LL�L0D@���LAA$�AA0A�A�DA�D�ALBФ03@1��D�$�A$@3A0DII@��DA@A�ILA0D@LLAPDL	@I�L@2AILA0D	0D�L�D$�L�I L@L$0 L0I$�@1�@�A$$��LI$�DX�$�2@�$$�,�@�$B�dX	�$�2A$�0�I �0@��03 ��00,�L��030�0303D�	��`&� ���"	���&� $� �`�	�`��&`f`I�"a�`�&	�a	�`���(f	�Bb"b �$�(f	�b���<���c���xЛ�8.)�b�������E &TA���7�q3�K�����q����y�O��S��~�8M~�����>�������7"?���?���n��p`������|w�����&�'���a��c�9�n�}>g�������zt�&���g����� ?���_L�`�����4/��?Z�
?�$��%TP���!K�����c�-���O�����?�I0S��P��v�}�����;?h|�~
'�?�U �?���~��?)$D<	��9 ��|b)���&�?s�(��ڝ)��d���̜��m(�9�q�'Hp�Z���RQ[��~����ӻ����O�r|?�������h�2Ҋ*� ���8� b`(�P!�}TR %
���H���w?B\7�0Q!
B��~�"���W���~
��?&� C " A�" �"E��" Q �D�A�S����} ���O�|A���)��<�`?8?;@�@��b����?R������mr�?X�`����C�J?�������}����tC�>o�x��ݜ� ����[�� ������l?�$�?�>/��ϊ��a��~������UE >t>�Y���j�?������{;y{��>�T�~#�� 	��Ȫ� }��X�P������fS�X�ҟi��O���wW�����:K��L8@�`Q���H)'�4Ɵ�aa�M>5 � �&����w ��	�������������\�C�7C��~�!�:�cBq�؎�	�5�gb~��T �9��O�������~N�TP�~cu��`���?7�	�㶔?���������$��O��>�X�?�>�������ߤ�$\�SI����G����Q�vy�Q@��l�̢g�S@?����ꨠ@�g���~��� �>C���>`����)���'O㑥>\�r�3���D}?�X�[5������0��u�!�@~O���>d�R$<P/������τP��T)���-$����� �p�ј�X���?��@��=����=='��$'�8s�������<?����/��~a�	QG�A��7O�&����O��W�����>��<QG�O����>�͋��q�ˀ�hs��~����1�i��:��!��ߏ���H�

 &�