BZh91AY&SYP�0W�~߀`p���"� ����bE~�   >>}�@j�ٍ !���)6�E*�6j�-V��-�DTB���6*�TA�`��lI�6�+S#&��	
-f�m�U���zu tI��-�UMJn�Uɴ�c`Ŭ��l�bŵ(�[��V�-�l��%�SU�5�k2j�m�5�M�@�Pf2V�-��7�{��4md5���gUU�M��m{��^�h�FU�6fV�Ȋ�m�I��Y���������5ZI��U-�i��V��̐�[�,5�6�j�+V���M��I��   .N��nлk��UR��gCl+��˧F��4�E���k�s�:[�5$��*�0Smm�X���5�ֵtk���D�5$�ֶMj��mmR��  ��@}��W�-��h4�I�p�Z*��;�:iJ���U�AYR�K�ԫ�Dn�ݽ[5�ڥw}��}|�z������Kf�5��|�}�[��*IJ��+UZ	�Z�ڢ�g�  �|�jP�������)�4|�}�_Zo`:鯽�|���w/��z{�TU}�O>�y��"z}Y�sR����=���M2V�{��{�N�V��ݼ�zt֗{&�֤�a��J[,|   gw�_l�2�}��W�ބ�m���z_{�A�Ԧ�����[׍>��J�>�x������s�^���Yw�p������]Ov{�5��kǽ<==2���u�l4�*��mdT7�  ��z�[J���-�@i�z}UkW٦>a�*��j�y��oTocһo=L<��-)�ܧ�jkM��=����R�w����m�hU�^��zjt��QE��l��ѕ�k$�  ��O�z5�SsǞ�{۝4ַ�-޴�wk������4���y�z[h:{���vSn�y���k�J�Q�T����Ǘ�:uv׏,ҽ4罨6���j��`i�SM-f��   ;�[��`�6ڝ��*��Ww{�=�@t׻t����z�*��㊥��{��=���=:ڱ�E�*���9���J]��n��h���]oyF	����&�FF�l�[o�  _�O�}^p� MspP�:Z�ր�NpU�V���{ٻ@�j���n��t �s����)��6�J65%�fo�  ǅR�V��8��{<W h��=j�z���x�*�7r���� f� ��p����mmZ�Hԛb�4X��   n<H���}�N  fu� 0� � p]t��GC��c�P�4�LE�����    ��2��Ph2 �M  �{M�(�@��44�)�1	J��� h    ��$�U` 	�  F��&��4�  44 &�$$Ԇ��'��Q�G���j�S�5��������XF�nϵmm�b��W�[kc�<�p�3��s�{����������� $�@HC�I$�BI��!$���S�p!���?��!�r�BH��tT_�А�BI�!�pd��iHBI�������C�Đ�d��Ic	,d%�$�$�$�ĀX��H$!b,IĐ,B� X��0�!b,@c$�0�,d��,@�@�0�@,H� X� � X�%�$� X�2Ib X�2@��B�$����X� ��X�@��b,`�ĐbI!,`B�	,@�X�HB� �$������a ,dBĄX�B! c	!I X���	X�HB�HX��!���,`@��B@�,`@����$�K� �BK	X�,B� �bI$I$,`bX��B� B�KA�$�!%�IbBX�K	c	,I%�c$�1��X��X� � � ,I%�$���$��1!,d%���P��+;�~��z���=�'������eg�[x+%�����\U7ssol]�L�T	�5A,�cN�!d0(A,��v��8lh�w)+��o]�1+�-T�K�]D�ԨV�>t)UއJ%m;_!�m�S6R8e�;�,G
B��[i0�w:��Z1�e��ˠ�Ù��J����q�CN��Da��{L��A͇S+V�a�VU�7���&>p�0���]+����CA��� ���>�Bmj�j�6j����#N�U+i��ۤ�#?j¥��(�{��)���`6	��[Wx�ǅ�v�3q7�[`��f���vMl$�|j���5;aǦ[�w4*�>N|j���L�]�[@����a�
c0,%pe�mX���z!�% M��GBp��Yo��ۭŕ��g7-9�	b^���R�am�B�֌�|P�Π�Y�����e^�$Y�N�Y��7J�&���w.���$2ӫ!kŎ�wc��»���95Ý�Ak�Y���\m��;Zf�h�hY��WV��Z��)ݺ��TX���M
̓	�ĝ���t
d���A1���gY�vY+i�K6�6�2�o>�i��]j�Ra�:QO�Zx��+��"`�eU�D�rıR�0v�+7Kv���lj��]"i�w7u�f��-�������n'J�Ĺ���ML��m�Z�bٚr�ҦZ�x^*:��Q��������	r�ZۭI�.tk�@Y�}���W�W^=��%�E;�02�� ������:��������)P��Q"�nӖw!Ŗ�r=j�Y�`�ݭ���z��r���,�a��"Lˑ)dh9@E#����-���;Q�i�h��PЃ�4�-�����!峒PܫOv�C!G`�/�F~r�nk��b�1�U��A^k+h��KD6��/kj�!J���d��xa3hB�le̫T^$m�'7p�]'L��%-&ed��00�5&��Ж0=ͦ�K�{e�p�R�: ����Z4��������`B�`k&cD���
#n���N��v4$p虍湮&�զ��������z\���dRr}CD�I���Y���^KG�z�x�p�a����$k�o
���f��I�oN�eZ��fk���q�%Xp詹���U�֊��J-j�K��b�ë8�{���	��x��#XV?�"ۦ2��n�����~3Bzf��3dy��l�9mc���*��
laѡ��.��83lԧI�K/$`dT�i;��ԯKy��Ӂ�dnڱ,`��֥ik/"�2G��Z')I0�E��ǐ^��y���'��Z�H/d��:̨���f�&���g�*^.�VF��vyO
�0Q�2\T�N��X(V^a��id��x:��F��b)zI�Z�h2�3�wᮈ�ݗ�`�G!Ŧ��Y/so T�@\���]���`���N�:m�-���}��!�����:h��5�-�HЊK{,a���JML.V�k�p���������uin�=1-�Є7�q�fEPa²��V4f���3n�(���5��k�	���B����eiF�4�Ʒq�n,�R�$M��+4��.����,'xM�6��慮5��jf�=	���:Yb�GW.��[zш�A�\׹N[�a�u(U��ɻ�/hh�v���2N6ʱ����@[L*�1,Y����qc7t��[W-Ce���7�e�$b�״����oRj<�Z���ij���v��ua���T
�f +vPV���((���utt!�hݲ�K�
:�maxಕ�	�0ݍ�,'hZ�m<�U�d�n��-Ո��/m���c^�Nmgs]�51\�V�칌�b�6��+��R["�����e��^D��p��hf��ћ���+)��S��YW�z��3�Q���tm�q[��p捼�u�e�xi���`���z���M�Zj52�6�I[�u�:u��:-C��Z-�ҶlF���[�rliB��Z��Bښ��]����íf�2�o�gr�,�f:x̆+k���<`���V��a��nd�l�K�wV�2�jmL�i�ܬTN:s%=�֩��݃�����72'F�d-�Ugm:ɇc�1�����p���a��4<��ES��'٧F5�m+HDhY�{s[�ୡ�:I�"��гrC�Ll&E��v��ʨ���~׆lz)f�QnR�׋&@rBU�����ᖀ'��Ĵ��s��*Ͳ�x�-�_��E�47�pf�b�S�7hS3j���e�<�q�v0*�.��kge��t��u	+3!�r��a�4�8&2ޛ�B��;UY{��Z��Ʉ�t�氌.�@�̣�1�U�h�n�(�oj��j�XBŲ4X�������wE�Gs$O?^Yܱ�y��Md��}�w��
qҹQDbL�~��w���*�ub�
zj<���kZ9�.}1�v�y3r
e�x�Tƻ�eC�Rm+Z��լ�9�Yy��s��$<�]:e�wWM�;��B�,0C��7T�s�ܬ�k2�K'S�'�QYc�����Cq7ī�ia$��
*�P4F�!n��b�ݷa�G+(�ˠ�X�ұ�k(���-��Զ�����b^��N2�S-�%=�E��&��ڢT�q���lf�ٻs:wQ,��#��A�ske�f${d�"� �Y�pH����q�Ԋ�E���B!l�	��P3�����sY�őG�bX4d�xh��y�Ʌ˳� m��X� {��"�)��]��B�ֲ��m0y6U�,����F��u��5a��au���!(��-V��0�q3���^��ʱج�$�-7Э��ʑ�Jm�J�Yk7;-= .�H�Dg��\tâv��&f�nij�f&�+E�TF�A�$�l���I���f�;�޶6�,����L�К*��i�M�X�&���8���ki����wb̭K[KBJD��2�E�̙x5���KE���n�9h�E��	� �����!a��s%�l8jM�l��R;���D@o&a� syp��+6���6�[r�ux�-�g\o&9���x�So6��z��FM1�G/];��U��xm��M��<;��Ϧ�>5z(s^,�S�(!p�q�kP�
�:����q�U�b�Z(��(�ɩ�{y�M���Խ
]k654�@�_�;!%��nZӦ�@�K�TA�{�7w�����d���ݩM�/f��:�&�Z&�÷,��t�n�4�H��d���R�(;OL�<�"�`�tG(m��mbq:����8 �hI��fU�t�k���@*�2�o�B�H��3���`O�5�Y�{J�'-�ii�񖴬�Rd�U�V�N�ج�L�n=��ݚ�Y���5(^�[�*��Ǜ�-k���q%�Z�%XA��i9z����,F�����W��ј�[��rⴚ.]�6��2�"�6�5�c��8免xn�h��jߖ�2�|���Ԛ�Jf�tDPք��AW�ޕ���5� �XՅRۥF�a���q�S]=Z��z�V��Fq�Ը�Ո^J�i��cH{C6
L��!����7*�'�uʂ����"�đ�b.o%���11�,�#vB�9�%�޼�V��bȊ�.'$���Rch�ɇF��2$�Ħڍ�wxjfit^X�ب�\���&�|�G���͉h��2T�Z�4R��J��̱�GY��LYWi,t�fa�Y*��2�K�/>
Cd͓]7�f��b�����V�����Ƀ/q�@uԂ�o�x6��M�Y��Q��R�ґ�^-:��jV��)��F�-���mh�`/7W�Qo���M䳵�8nSCf-�f٤%�f�R���X1`w�J��6Z/qKn���Xcn�׎+ U�r�8�$q���6	dÉL@���b�ܭ�/+�y�@�T.�3Y��ѵֶ���m�ۭ��$�n����GRS��H�:/2���^�[R��e���tە�z�ƴ!@���Uf�%�J��D�R �M%��t���E�ģ�S�iD����S��z��W��4�	�z`����r�6�v�����n�n�pmP��o�kE�5��F>5B�AR�^�Z�Y�t,���ĵS���Z� �{Hc���Ǫ=є���mHMnD�O���ޔ�|�
����kq*��%dM�A�o]�m�I���.��2�[n��֦��4��]f�N�fV@�No76l�b�w�/U��F�� @F%n;1�fKQ����A�/�;`:����܋���R�'oS@B���Ep2F�u^���"j�3.Q;�q�iYYm���P٦�$VRx[�F�g(Y/󫧢�-�i�Tb�����(Ōܹ��w��J��	�fY�v�4F�7#x*՝Keźq=�}�� �ˈ���]m:�FR^ n�R�Dҁ�kl��ǻN,VNY�⡛x��z�-��ԫ��k�U�]��R͈㴅�ٺc{a��@$F��$�FhR�^T����YstUjJ�*�z�=�Z�k�ܭ�]��sk.SAtɫ���Vm�ɔ��ȃꔱ�'f.��T�V^�&nX�CJ�l���l���]7IŁ`Ɂ"�C�CR� E�2�6n�����z�9-�Z�=
��tރC���Z�A�ɥ���F۳6�S�۩#�ҥŲ�e�n�=R�'�Ô4a�J�L�-�E�ԣḃ��	Y��Z%f��k��X�k�P��?.�_=�3��,'�m�V��ވUn�]T��Rd*�œMcfRf����nC�A^�f]Y<6����J���t��݃���*�=�)�k�����[T�kv�*�	j�R�+k�:�Rv���nSw[�SU�n��$��nV��k6kn
4q�ə�`�`��1᧔MM4Иs�a�5��� 7Vb��&X)hm[`�z�@Ǝ=Xym�e��y��;�Im>c�(ZfՂw�8�)R�A���D�f�S���J�+Z =b��۸�3�ġ��2Ғ	��`q5z2�˺�����*�����;/7��|z��u���s.��E�H�؟;b�c�:�������ر�nE��7B1I;��F�q����Fh��Oe㳚/U���`he�F^��YUP[��h�/�Т	i����٬U��4��h$+^m�q�9��d�z���F)�SN�9T�����:�K�1�)Ďg�W���a���Ǒ*͎��耫1d�6a�OB�Ϸ����}J��W��b�V�o&��9�v$���1;ܧF��-�@�9�A��������j�����T��`�e���՗+9�[��L�4Q��`�-�*��Ņn�,(\���&�.Z�p]k�Qܥͽ��6���X𤳖�㸰���#kt]�Je��Z��ڬ5����H��౏�@Jl���P�u�f��D%�g0��wY��i����dohJ�[�*�v�fXz���/�+!|(���-5��&j��EZW1��M� t�˷Y��0ek6�ܚ�dѺ5-��L3-J�7�g6��ec*�am͋)�"���pl9z���;��{�U�☰#Z��޲�f�т�Ғ3m��2�=4�0�ޥ�B�r�����V�#ڙD���cҋ�3vA��aڼ?��zwm�+��^�"���㈉�ݦ�̽7av��#��t.B��#!sh��-f�<�F:M�V��Ul*saٚk.�����T���PFf��&B��B#Ԝ
;�s#ј!="���+"[��غ��H��V�V���>�Z�S��i,8�'�	�aԶDl1>m��J̘Ňt�Y�Q5qANeIn����e�y%��{Q3���^9��v��eV��ej�"��akQ�x2�MApjvJ�(&j�ɳvC��\�y�$�t��_ؠoo~��FTJ�����M��7�mև�9�0)ZV,�[���.ąB�^ŵ�Y�v�%uv�Z�y�7m�{���il�JC2�0�B
�|f]iY��\�����4].�t%]�qI1ǹ�)zw�]F1�<9��ʧ��v��/l��u1���O%3IzE�I����.T�"^��2R�6haU2d��Xh�Am�f��r#l�<{��b�W:�Kpif�鶝���`b[ʽ66�n8��I��e�w�4@e��Rm�Q�	���ƨ�"��T�L��n�x);�ȵ6�r�����-��S͠��c2�$�W���� 袅����j]X����+sP� f�G-)z,�mMS)JzoubL7�]=��E�	���Y��梯0��|�D�%�lOfe�ńb�`���#.n���V�T�6A�੸l��F%ņފ���Ib-����>[����;�SYy�V6�	i:��X�����eK�P�l87w!�Z&P�z��4���r���´�?�Dn��s6�F�N�����儋`�)�;ձ��T���o�&ʙz��M< 0�VX���)ԥ_p)��p�8�u�e�ub��aZ�-T�dU(�[�ҕYDY"=:2����70� llɆf*��Ӽ���V�軇n�XͱBY�7�S6G��/Z�WkC
����+(\kt7r��R�2�A�F�t��6T�Z�+-����.�2Z�@�ES��3S�t��[�� ٨R��7Aьm�	z]M�.�G1�����i�A�q*��T������օ7�'�7h�)=Y��/�������'z�мKo4`�zS���N'�7^F�hc��Gd<���+j�6NE�I�Q���������
~t��?���5�B��/-̥��j��+��s�IJ�_W�S���E�%m�b��b1t�k�Q����ro�0�k.�S��E��9u��W��Yi]�ޛ�=�d�j��4����U4��f�S����67G�^����J��.���,���Y���y�ӕ�&�ןk���|��� �Y�}9���Uo�~�>�ݽ����5�y��r�%�X�A�3�-Iy���6�>�F������r�5��pGџ��kiI^m����sw-��9��wMi�p�7�,Ѧ%32�qW���D�x� �3rP�nwu쇈�;���/�:�:c]�r�ޤ`��RN�n8O&��e�]eeݞ:���tݗ��T�0�/m��	�A^�gA�n�k7qH�W՛OwM�0������ά����*�R�<{���׏4��a��U|v�Sj 5�'	�N '���ː�/�4�U�w�i���\�_cv���#��:cp#[��L����P�޶��%�<r��+��ʘr���-�Z��:J���e�೶�Z���8�1�d{-����%"�G�%Zy�����YaJc��r��^K������w��Ɍ	��7��c���S�W"uǙ�Qr���v0�ΠNʜ!/�ݷ�V3fL��r��yo��2��{�釽���W�s�5��P�WXӢ��3'2q��06TU�s�&����g�+��ޏ�YD�ՀX�{ˀ�����#�!n�gvk=���o;L�\۳��@%8<�����"�e�<�9�6�t��I�oԥ�qT ��4�e���X��Z�- ��K��ʛ\)��{/D���(u&\wl�����Y�t�0��L�,ߺ��1��Ŭ��\�U�7�܋r[�bH��q�I<�6T]R�:V�]X/l���-vo.�ʃ:�|�s<�͖�A�#�|����OB�r���#�YN�ܠ�]))L%���D.�����ȅ�dX��/��e&vem��ǰ�Q�G�묒���1[�ޡY`�c�U���MW`�\W�0�Pˌ3[,Y}����AY��޻�ѧPJγY�+R�Z^!��pf��($���k[��6n���5k
V�mtw`�l��.X�x!{�m�-@�;��+k�i��k�ḎQ�G�Is��Xu�l�dV$ޔ���Y ��%͝�fa�g�.��}��5����s�~�u�Mp����?m���Bl�u��gw%����x�\9�B�s4�,��,]�]�]�6�pol�9�V��_\4/.W��2�o&k�3Zy�c��Ci�K̮�*�h���t��z�q�p��^�lHjO��� wU A���If��g[�!C2�e�xjd��C�K�^�Q���ZMKۉ+33Tc��N��٠�]0�ڲ�㫦����Ӑ�k �a.'j�:Y�]��d�_a;�m�C�tzw_"��4�[�ح�2QRR��2�{=s� 5�p��қ�u�N[�R��[��c��J�﹒rp�NYצ�V8�f� W��>|�ع�xk����˛)�]#}�� ���๧T짜
c�0����;�^�M�4r�;�ɗ	�3����Aas�b۬�_&���۽�����ZyE�U�1�ŽRl�u�9��o+/79 ��2��&�(����X�9Y�o^/��B�賓��箵���`c�3'�"W:�}u���
N�Mn %��܆�M�T���f��)��D�D�\<�ic/{n��͸���ǃ�F�*dU�.����d�����KA�q�e�o79eL=��.��^gJDl=v����(1�R{[K^�@�pm^:'S�BE�'$Ϫl�͊Z� ��:t�x�7e��zLD'>.i�����qݫ��;�7�`w[ݱ�P�q`Ýb�F��n��;�l�{�fjkJ�Y��S[�`xu[��O�w׫�P:���[�V�9�4є'��oN�7�7�C�4��H���ԘT)�\���X�ջGs���2��N��8^�]�����������w^彮����'&�h[^޻��d�2�+s����ےi���9�f��*Tۉ
�������&�o��	U����s+-NN�f4C�&)�ʙL�rt��Pcd��r3Kk��lS��Ȃp�r�{%��R�m�Ʒ^dܑM|i[�b&ұt"-fd��3�G�h��*��V�L��!X��[�͸���+��*m��xL��Z��R�J�W�0���t��p�á�֋�ń:�%����Fj9��GzKg:��Ŋ����Z/Vc�	�M��8�4���~�9ｭyb�>��d���H���u��kmB�Z)���:��N�fFrΐ�D9Hv�\�FTY\]�9����6<3\��#*4��wAf>םXiT����Ԭ��e!!�����E���wF&s������!��Ǵ2�s;�jۥ�dA��g;2�x���j���N�=s�Q��f��%���,Nf���Gv���jV��"��ū_D2���9U�N�u�G��M�U��y��o�@Zw$��6�tGq�V�X�[訳ӱ���	-��Q�v	�,����V�%%�á]����/���s���3f�[L_r{��N�ad.|�&�)�=�8�����k7*%�Ȕ5oI3����,�C���vCi2Yh�/�OHt+Щͷ�B�G�4�ǆ��S���5mk-؂��N�ha��e\���N��n66��{͗���r�@ �N$g�^H7(鼾w4EY2+�E��ɢݑe_IW]rQ�:�s��*�-�Y���5o'h��V�Ib��H-x���w[9�gSÒ�HM����`-:�K?*8D6x����חb�w�;bt�u��c3m��.k�t��@Pj�Բ�Ni��me����Uړ�|�5�w;_<���`�`ʋ%�F���[��|V�X��ֈ�2�N�F�#V٣� �Z�7 ��t��h`���}۝q�7�4+q,��(5 ���tZ?6��)�x	��.�LY`�8�ܱ��<�3�K���"�c�ǵoR2�i�[˻s�o"Ղ�P���Gs4��̽���/;�;QP�2�c4�;P�=�
�G��0vq9�+s.�2:�P�*Ӥ3�v�Img��U�]�P\��ec�±�:��C�0r�D^3�Z�>#��f�KC�Fb͏u�����8fS�0�� 7�dzºƾ��!R�S�
���#=�q5�r��M3��NWw����y�w&h4ŻZ���-�$L�y���]c�E�����}��=kg^�M�ӋU,���ncG.��i�m�l�η�G���},A���c�IkZI��U�Ba�d�o��h���
��t2V^p�9�c��1�z�Dk�����%��`r��`������z�˩j������m��:*�*��WU��p갠�4�>|�����]irs��J��f<�F�(��2�N9���+��vn����uz��Yē�Mj�
�L���l�{�'�'�t��Fjv��v�oyr:��,�h����f�1�Vl�������d��v���tЮWn�����9�+׋�����c7�O�eG"��Z�*�3ua�>1n�)@�-���a�n�Õ-�!����I:��.��e�r���\������oK�u����W|�^.�)<�R��+�˱���.�f���eI���+]��$�P��M��&DnH�9�wWOw��\a���Qd��r�h�h��"љ@�7V�����3^���="�.���y��M�yE��t(���
�ј���Tڝ��g,��Wu��+;TN��WŦ�����\��T��:�vl\�\�<��N�� cI&��sͲ;��cJY|�\���y���B���׍����	��̈p�%[�(=GX2Hvqv)�1�x3:�
'��v4�]�x���oC�O7lbx�;',�'=
���7���zV2�ejwBL�aQ�J����Z�4�Z���P��p{̻쇸� �VV3�	�7E�h'�������k�&��6�G> ml����4{o ,<�yȌ��v$(L�̄ab�u˻8�	�+�ԝ��V��+2uٱ�p��1�W(QGh��7�.����b�)ۼ�9�R���pɝM9��0�]���WP�C�>1ѓ��;j��v9�7����gm�(�}8�,s��ü'�`7S�f�agA���To����R �mس�0h�m����U\<����c���glZ��r] ��Q�jT�5��t�5� �6\{+^QŪ��+�r� :Զ�]{V�����#������7B�.��P jT@�����s1����+����<ř�1�y ��&���j��ٰtg�o_p��gu��\�j��̂h�w�t�el��˼Ӽ����qxٮ��fWS\�[jR.�^�J�Sx^���;�J
� ���r�ǁ�pK���s��%_�ͪ4q��$�]૧�2�:��4S�$ �n�	�p���%�6�ۣ�lS�f����V��������<���lfT���ړ�Gk'��ے������,��gM�b\�f<	P8�xj�Tꑫ��#+���(a��7�Ĕ$d���'��mu�a(0ǛO�C��Ԋ�[����gQ�y:��� �� �9�D%:��%h�U>Z�!im���{[�5)��z��}�5�[���P���N击.]o��A9{$����M5��w&�Xc33sc37�Ǹq�e���@�w�p���M�Sp*d��R˙4t�d��t�񵺆nn���C�9�n�x�`
/5��=C�ɒ��B���\MM3-a�'RX�\�]B�(þ/B%G�ia�So�)��y�ޗ/��m�M�i�MK��V���<���XN�F��*�0V�d��	��]������2��n\mMI�sCκ`�mo2�l�t�ոzڑ괗9W[w���6Q=!�z��o�-pJ��̘��6�lu6���R,�w+IJi�vpK]��ˡk�wP؃�d�W�Mi&Bl�v�WYI�dmӊ���c_Iՙ����*�i�r�|��"U�e��U�DTOk(��˒�Aƒ��F+�����P}O����F>��ͬx�Z:E�.���Z��)�`h��yۡ�'j����c�n�u�kK�Ѵ(��q�d.pA`ƍ���V��!�8_���9���Hm�%�f�����ٲ'fFv��f��!q�V�j��m�x�1�UmN״�4L�ky��	�M���5��r���¥�d܉�d�f�ۢ�r]�C��f�/�viTE�ڝ>�@̛���<�V�uϬ1��*���NoD�g-X����Gd� �rg+�%�������k�sp޽�+�|N8����Ԉ]�MT�1�4���F(_V�X���뫘�N�c��bY-M3�Wqʽ���<�̬�AiS�A.fM\�v�u�dz�o7vv5Mf@�ن��ړ:+��q|�Ś�g7�~� �n��d]R���m��,T���^¶�����9	J����B���HC<���^�)N�8��]>Y�,�,Aq߄�j�����WX�b�P�w#;�#QkW"�هUQ�́i�ϻVrGi�e�0q'�f法�7jm�`���,�+X��g f^r:�V��{s�T���Uo�.'zEL���&7M�-��f.��;J��7�p�S�RewM��<���\l���G) �eF���1���#���� �֡v��J�<)~ꋖx{}���ɬ�lv6�Wv��6FO��XATN]��j�ǻc��0D�b�Ue:�PTbGs�ws1�����7����a<��gQ�}\���r�b�B��w1}�k��6��:��.a+���re=}�;ܕe�v�#Z��7l�mi%U�;ά��2%iۙvg2��Í��[�KViMth�x���[!j��

!����n�6^�N�[�Ź�67J�-�hoFQ���C��	&닊��a�wi��˖�R�sl�u��lw���CD��Ne�m��
��$�'X�s%hz�Ӭт+�9��4��o%�~��#'	}Ǳ�o��u�7�[j�2F�Ԙ�o�^�g�*�g�h�>r����@���2�F��Lv/��<8B�ii�
�OUX�o�Sc<FV �.�&<�}T���
�ۙ[/�ge���� ��!B%�`y���Z�n,]�n�aN�yϣc�X6M����!���q���XC,ݝO	���]4��roD��V0�9_8���|OJXrC��@�dm+ƺ��P^��%���V> I����Uį�jE���YOE֤a��m��٧���K����{o3��L�C��o��}C{0�]8 ��+�Ԥ���dѸ�����i٘��STw�Oo;��y������9�j�)����G�u�ډ�ۇ��]��mG��ml���B�������22��!����~ꂲTAe�"��}�ϰ(��0�z�R�4��s�Q�{rw%�:�����V�/7m�8���Y�݊Lju	�
��/i�W1�����5tP�/D�錒���u���ׂ�Oc����쥰n����T�N`�R(�_	�pw�Sz!js̫R�P�^�S5�vV�+��a��]�t����.��6)�cv� ��f��'��g�$��hVY�Ns0c���=����*6a*^�ɐL�{�f&i8e�M陽�Zh��cHI"�4'JT5���ޒeZ�����2��l�:,����'H⭊k����N�f��h�\�Jc� :�167*��Ivr�:�� .�Q�3;y��Y��%0�r��*�K�Q�U�R���mnau�֨T����VN�.x�9���L乸,���c��v�bp��J���X�5�t,�j1"-��	R���H�_VV�cQv�r���wnWn��G$rI$�9$��9$��I4�b���t�w����t�!�щH�㪧)�Kq�(��KkMCN�2C�Ȍ����P�!��*���©����F�UQ$�� .�8h
(��	Ϝ9oN�=�����5�v㿾I �I?W�?��� @ ���G����� �I	?͈�>��w�������F��%*���Uݟ�0���l+@�^�o@ɒ.��.�u�OM��y۶�7���j�e�`2����8�k�`gv�3����f�L��`˷oQ�帓���U�	�p����G-��n�KcQoN�����)Ҵ1��x9Á����sV��e0�ỨM	��y�t\�����M�cVV��^a��E1L�K@��]u����Ȱ.0�W�6R-��%V�F�܌�W�SYY��ଜ���lu�QA���j�v(TV�M�v���CHas�zJ�\�B��$7w/e���M=���',���a3-�rmL4�.c��\�S̓����g- �1%5�.�(�u;}�XS����Ҏ�b�}�b]��JESx�̹��7]���7�_u��ٺ�klAn�zLxt���8���l�@�q��a��kX�Rh���X�T�Ԑ-���a�R�᫽�_X&��W!���V�\v��ۘ伕���r�-�����+/�����vD3.������U���B2��B].�&�%\d�l�z6�KۘVa;�hb�ࢹB�Lgnh��e��qq)����v�����ɔ�"��8�wk2�!3�L���NoH	f��jY��j�]�|CЯ'a�V��n��5��ʇcBKD+��Բ9vx@��tl�L|Ɗc�n��[���>�w����o����{���o����{���w���'ɧ��|�&�i�r3��>O���>O���>K��}>�O�����}>O�����|6ң�K���t��œ:R��_<���Gul��y��	�Jy�:��\�l�Z����������V�1unl9��w��X͛Ǐ3j���Д֛��2����VN���2"���qd��K��
(^=��wX�:������-gi��
�,g���k��kXY��h��s���'q� 2|Ƨt����V=r��G3 ����J���1:=8l�u|y��|�4erN�d�e~�b�u@�I$z-*�©�(��F�%Kbr�ee	��S�-��׌�[���n�q��B�&���a��mno��g�����^�9�84�X�p��]EV���Q�՚-u,��/���V[��m�~ƒȷL�:)V���YQ&���vP�t�`���VT�(�8�
]u���%�m���[h�=CS'`�����i4�^��e
7���I��[zxgQ6uX�(��8��r)0u%���ٵ�>_9ΡԎ�РC��2']v�6P�U���r�ˬ�:���)���r�Ʋ��K�_UE��Ro��V��t�l-M�u��ͺ�3�ՇrK��G���4s�����
�s��a���Uoz���n(�t�n�¬@*<ס�n�/�	���-гl'҄��{/��y� e>9ҥW�ؠ�q3Q�yw�&���*{]�oQ.����]=�\q���I`��;�NY���R��=�Kp��A�j^�/+5�XB�tw���}>�_����z}��w����{��w����{���t��|�'&�i�|�%�'��|�'��z�'��_�����}>�/�����}>Y�O)V^V��rp�X�E�օ���1�9�!�-�u%B��L��pY ���瘦��/��x��N��Sxڮ�N�ҕ���]����%	і�Y{��=f�Nt�U��vc����n�rԻ�����'w�5Zxm�������9sur�_q��,m����mѾ�����$x �U�N�bC.��u�g�b2b���r�Dk�B�#�)�M�v��R�M�fh�N�}{ۂ�9J�Z:���V�儹��qJ�k1Z�lN�BM��B��L.ΫK�'pG�=��¸���2(���C��ۈDƝ�Ջ6�ᮋ��j�!8�QKF]`c!L��w՗�F�,�!z�r gФ#��Ϟ���bV�B����m��-!C;s�Ey�La��-�O�@�����l���]���w+碡(�F����6F]�{NҮ�Y�c-c��N��}˜c]>���qm5�/�]f������*a6���ؕ��T�$��]҂��!w*eal=��๦�b|dօ�v{{���d���=ǵ7	�s^�>�}�"�W�����_>�*��ÃaQ�w
}q}/#��v��X�6n�C1W_=�Е-Vcr�ϻ�C�%\��H��F�m�N7�[�auLtƽ��.�d�f��níu�U�XxaH͔8=��*'׼�\�m�7s,Y�bɫ���7�u��5��]�̺˭j���Ly��<y�%=�uGh�����N�=AYn�A�0��Ӏ���0Q����[��0��s�Z�qt��k٠��ٝ�P�ɷ��"x�b]�p`���<琭�6�=���NjG�%���[;���Uw�m#s9����si��Y����'�^,�+�V�O� [R���%z7�r�v���(��z�Z��.T��	}�k��.Cp�m�Z3����ag�[�Г-ty���
=R���A9��g2p:Ef"���r���Kr�vjN��Թ�n�8�g��2i���[f�����RR;%�n�J�����JTwo�×�ګ�y���b�^4$�	Y�AxN	��fn��`a�r��t��_L�ꆴMJ�b��V���V;�泵�]�iqF�X�lް�����\��-8m_C}c��t<��W�,��b�#`�2ʀ��h�3����'eG׶�ܤxԄ��:��"Z��Bk��-� �k�GP8�8�ᬆ�+����U��o��p����╧~���oC�2�n&�Mm��ᥚHU��L�ӵ�����������:����R�6�. ���pJ[��U�V�o����cdz^���WP��􊃦A��`�޷�c�}����c�+�q螜j�B0T�[����a}��Uə�+�r�8���Y	]M�ٕ3
� ���Q�@�NfXճ����s�9M�dnr�C ���G�9��r����M�������K�n�8ں��]^J7��z��̵���	�uv��4n�s��,o|_X� `�Ra�^Fm-ʵˈ�G3|�s5c�w7iU�}���:�b���ۍ��u�m&�n�́��Y���V�۾HP���JK/���h�B����{dm���r[PX�k�n��a��S�k�_����7�E��k�q�L�*�cEs��^E}\^�k���_��hf�Өһ1H�L��'G���R�g�U׳d�$�6�ngv]�B��Y�&���~��5�׺��T���FS�ʤ�މ�Z=x�V]`|����d���et����r�ʢj�n���N��Anb��T98,�@ʌm&5S�� 0G���X�/�&,�bm��@)8�����_r�qd���'��+p|��d�^��o��ޛ���GY�r�:�,������V�=r� ���S.�k�̮��8:akWV�+#���tb��)菱AJ��8ܼm�0����`�YW��J�������Vk��`�VJ;�an��c��t�4�����k�<k�9y��B��د'*���*����oC����o����Ljl����C�b�M0���\R� ,���'��һs��I��0�n�!7��d�U!�\1H]�z�)qi#$�'-��q��d� ���(p �:������ڈ*j�@�'V$�N��l�ܰ��x1k�H�$��w��u\wo`Ѯl"�$���7d؛7;mh�n[�"dF�0�g6�
���yk#a�l��n�	��ЦnvqR�/K�#XR��d�K�eڄ�J���]�̄s�7X�N��
r�n�W��]�T*�]/����nk|� V��1t�B�T��Cf�'P��Z�U�4 �iSUC8\ޫv8�t�GYn����1�]A�JU)ѷ`���ݩY����n+�np�4;��(=-�d%���+,���HL.;xr�Z�7�XӴ9�n�*jf9��Ty����4R-�ʒ�ŐŦ�e��p�.��،Q4Z럸�Q����;Yǃ^Ì�9z/�[El�����m)�:��ŵDI�&�+p=iN�YѸ�Žf�>\�j�Tv���+"��i1+3,�%E�-�N������e�d�\9e6�A�B��u�5�m������ba@�C�R�oˁ�6J���Ml���DjO+�B`�l�MX'\���K��������A����mY�)��[����lg��U������J���"���ۻ���ʧ
�L�����V� ��3^s�D���aM���٧�s�V�Sz�C�Q,�<Ȱ`��)��4Z���;z�s7e�7�p�n(�S��E6�%Z��娠
"ol0�0S�Q5�1�Nb��@�뷷8eM)�=j��7e����u�>[h�]��7�ND��^ԭ��.#N���	���I��\[��JU ���j��o�褐݈�"��K�;z�Vo�}�����֎+�Lc;������HHo|�f/����*�v5H��@��ࣗ����U���۝���A�+[�z�<�i��u(���ᚥ��A,�$<�յ7�%��&�u*��pk7��}�\�uԣ��jZ���V�%��ur�L�K��-g�HXb�i룯U�E'x��s�:����o�o&�T%m�����ȼ���6G7�@�M��Pl�fZ.�4��q�O�i�\�7��s$hA��aq��i����ɷ��(�s�Kҫ��V�ɽ0	��闉�G�5�-ZW]��Y�`f;
����N-]�St�A�9��X�0m@5�W[����$_S�z;�C���W{�r��a�Ӑ����:�
)�T���\s��9�=��8���F�	��@u%�x�֛���d�N��%�ӡ͹W�B�40i�$�ګҳ�&�,�3�9lee:�:lb]O�A;�SnŬ�t�"�t������v��+F�[�DMʃ�r,Q�e��R6�z �iÙ8mcD
�ݔ��G��j���}]O
�܏�3�M:�'1�S�VL6�CM͹)��agl��3׃�Y-؝;�����v�}E��[/��3��®-�eWl��)\�:"�&+���!݅�'Ә��dg6 .���P�e��P[���Y�%P�ݡw3���$��2��Kh�7:>�GJ�n��-��fY��7S��ZP��?�t`J�����!���V��;���������ۍ���E�F��ćb������v��%]�m��Y��-�/r��
&����H0�|N� xٛ�£�R}{� w�c���)V����p��
�������f�w	�׵��:d���dduֺ��c���r�����Au� ���<T��.�We�O7}�ME�>'i��H�uE��$�GkQiئ�n%Z*}R���g����腬u��@U�_C�:��Q"|ڰMꡙN�_ovX��ĸ��f�푉����
�P�cvk�N�����y�l�B�e���A�9�HU���"�Hw�Ҕ�'Nff:�k��s�^=�;1�9Ө:|پ�U��[.)6c�ܢ��1i�����"{e(&\�)E-՝109L��⇅�Yʯ;��w�u�5�0*L�b�X�N^��f�c^W	�E{�Z [�۝v�6�t�Y��h��������5�b�7�Rw)��	%������9��b�w�w}2��L�_�7770�R�0Ě��Z*���o()j,[5`��D��{dm'��wal��L[�Yk2�^a�+���Z�l�E�-�ɨF�091�yZ_K$j����E��O��&n+��<+(r�zѭdJ�ͤ4�5�]1��l>W�F�֛��[���*4���l�ѫ��X�������@0m��H�ٷ|k�ԗd�";��aS��15�1�qd�:��gk@�8a�Tô,��wAj4F�{K�_
,ؑ}A��(e́�%<��vTP���O1魮��K�:4�����;�EZ�H�-��,����O��($ou�v�E��v�f%Tw�!PP�5�ľ��d&�~��5$����4d�P]Q�m��p c@�P�n7����k���0x�v�n�=K(q�bs:��k0�`�ȵِ���G�l,�X��S�����yt$�ۓ1��@�wO7n����7Nj�μ5�ޒt���z%V��V]m�xěx�ތ��6�e�νbn$���Z��n�Q�.�g�Du�B���y�I/���ģI�j�c76�0̍P
u��{[�F]om�N��mf��d�8��\ӨṼ�5�Ku�(����X����f1Xkf	���&�5.,�|9:̑�ٰ�?��w
�t�:��;h���*.1�32�(�΂u�˵��1ܨu̷.�DI-gP,nѠ��L�N����̱���ۉ��Vj�);#	(�f2���:t='5�.�;Jd�9ӥ� ��q=b�5wQ^�d��V�Ħ꾾"����� �j�M�)��c)�"��D��W�OcЦ�2P�4��Nelk��I�=�:�bw.����hmH�(��Jg�.b�@i�Uè7���P�&HG�9�s$��[F�^�����c�$�L1�w.-�0Æ�g7g�(������нf�N}��9X\�����H�墥h�t08("4A��˻�<��Sa�:��Uk����I��wN�����f�Cղ�W��q��H�ff�HŦ2v��#�f!$o��r�&io�Y�[�d�ӐQ�9�W$�:��b�hꔓ��z�[b׮�]����H�,��W��Vs�$"�F�\6�S��>��6�:��)ԗ7V*עT�	�ˮ8�ˎ;Yr�^�7����'6����t�aX--��-����k��7�M�Uu�J�U۱���;�}�������:�����֎��#$��IK5ɛ�u�o%��������s��lb��հG�,�io�����qW�<���+����%hIHÍ��.���H�ӷ�Fq�(�tڔ��"gPӣ]C���F����d�3bI������������O�C��}�_��!���/��4u��b� ��5���_��)��du�]V%9���Y1�y����I,{�FmL�2K��A��
��;XI�I��=�����>b5/��Wo^C�guVA)G�Y�R<���Y�����EXg�H`{�X3O�AX��ӎ�g��]n��ѽ�w�	�ؐ;*�3���K[y2�p�+�����N�:�5�q��X��3������ۢ�v�h��\�%e�����w�Z��m�dD*��8���D0�i��U�X�:�S/�����}��l�)�b�W��`EFs1�Bb�f�1�v4	L�Zp��Zݩ$z�,j����k�f�`�6�/nL�1U-U)�j����<�6:�J���p��!�RU��P_)`�[m��:q|k]4oR�U���n��o��^(5T��u�3����6���.��ˁԬ�YQ4Ei�k{e���X�j�Ը�������̩`����ħ�Vڴ���>����V�H�Ԩ`8D�{J�#ƦR��fs\\�����f×d��6�XU8������tI�w��g���6���c����܂���5�[�w�+�z"�+����ќ�,f�����xx��f'���}:�Ӡ61���L��&Q�k��ol���;d�LjW�.\F�t�4�ӣ��3[m�;�rMp�7+fX��y���c�q3�^g�fT+#O[!�(-��\X@m���q��*MiJ�j6�4Yg'g�����'ZZ�|f��!��`Vi�6y��":�v��Q���:�������S��2Vy֩���QH�-����O6aR��'�aL�ɓ+˵IP��Rw��j,�,��Zʪ�=뚊(���Y鵪dZ�E=7U*��u�[2T3�k#l\�(�K�3^b6��lQb�QD�r��*yl�����.�ĭJ�Nk*:�B#[hW9���f��-)b�m*#X����L(��B�h/Z��{�:�5*ɢ,�yomC�;���E�dQ��9�x͋-��R���pAj6�Jŕ�o)s+k*��#h6��UF
"x���ʕ[ej"�,E�Z�l�T�Qs
���xʨs��`����]�*,�R����Ö�YX�U|�X�3�
�yj�yJ�֢2�iV�
���a�+�Zq�*'�_!�e؀N��Q�n�gs��4j�i�2m�w*�z�'��Ie�U�Zǣ�#��b�3��KPC�ܺF�C��=��o�r�I\~��T|.Cz���S+�9iw�Rφ����嬜Gո|��_M�x���o��k7����&�c���z����m��c��ꡊ����&=���:��#��پ������2ō��h섙�s�K������S ����d����Wq��]�\$6�\Wd�K���Ǯ���E���:�����ur���k�\{Z]<�WM��w�|��;�'��WJv:� �k�r=�3=#�elT]_d��K����h��cՄ�<a���JW��{����f����!ޕ�Yᴩ��r�ž�:��ٞϗ1�Z�O?O��ON��k�ڨ���=���+Vx�ɨ�L������!~��R�'r�����A�ӗ���M�VfZ*rGX3P��� 坮�*���'f/ŋݦ������O�K������c[��#�^c�)vj*Mm��̻��Y�ėa+��j�h��O�,�F�#� ��Kx���0�F��x���ܰӷ���%1:�@�����)��N��H��q#y�tZ�w�[ �+.n�u7�ȽUϫ�of�h;��'N�影Ӥp�Vg����=��T��ˬ���/�g�*d���w����JAʽ���~��2r�ڸ~)�)������D�i���; ���Ѿ}v�드:����!��eŃ�"�`��e�v�nN�������mõ�[�'5�-�.ll6@g�`��1 ���y�V�����gΓ�c�띅),:^�����"߈��n\�����yRn���j{�*���2�w�N~̣�ٵ%)��A�7 >�e-7��2�^5�����=Td�r�.��)����ee��+�yq{|2��+�s}��X�ޘ��=	Xǭ�C�����߳�JY����̥�)�J��������]Wb���}閾�<�������C�;����童?7�z��c϶�����k�^�wC�c"��7�[�y����i�Gf�
I�ײ���4ox:u��罼x��V�u!�u��u�/,S�=�]������[V�v���Č��䆌Z��Ԝ�v�7-s�lf��u�5��ˆ,Lm�=eө
�s�:)��vk��X:����X�r�r7sY|#����t����� �I�n<h1��~�$ٝ� ��nT1}}�4���%+�bh����	M��R�/*�?`5'����Ћ�w}��*3{}�+�]�8]��ڿ,�oK7�n���8�����a���q�}fXGރ����
}f����`_G~qf?L�Çs��}��n`�֧��=�Գ��{���eS��f���yC�U�w�+�>�FF�L�xނ�,�Ed�n�9d��{T�{����B~�E����*z>�o�3����Y8�Y]<k�c^g�`�z'��5}C���je�O�nB@�`u��.�R���=�Rx�q�u7:���R��{|�b� �����D��́<f��}��u��,k�i�����v:�Ү�4����}��OU�y/+Ѳ/1�[Y���X|�\�/�G�ӳ=fK-�x�r�y <��<\9�#+�GԨ�9f)�ݬm�fH�^6��&�Ν��>'T��e�?-��K���ENŚC�G�t����n������-盭����2!�̴� 
�M:L��š���'�dT_Z�Ū��Ҹ��c7�Ψ�L5!հ�%]A���#��g��^}�»0�6�-x���'�����VH�o{��3���d����uދ�藲����Ic�X�������b��IeR�gԜ���P�9]��Y��	ܽ�k&l���m7O`�ZXm��{ygM�W�P���Ć�g�������v���}&"��,!��⦎ʥO߳L`ݵ�n>��@V�S~��==<�N<�Lg�_j~�+��PDo���j�ey�M���m�����:ė������\���9Xd��E�w���0K��a���9>�;��C��:�A���`�Y�/��O�[��n{ֺ?k��~���>�~��U_P�����[���:̽�6���mҔ�������9�s\Ϩ��q�:�۞�oG�<_��Ӓ6�T~z�&J����#���}��$�qc�G�Zb:ns��9�3B����XBu�mؼ��)j�U�S��QYcm�x��7���%����jeI�˺.�w^�%���[{�<z�[�A�ő�X핣{zm��'N&V�)�
YM�2��Η:`P��1X9�����`��F�����x�gqH���S
}�J@�m��]�5񛄟�>@��\��z�k��#�5P8�}[������n5V��-��D��|}���Cr�<���c�k`���Y�z�!�o5�[v��^�UN>�wS�@������3�t�T�?K�+N̹\��=,莦�c��øQ֐L����1��� <f_L<����Þ��s���Pw����6�i_����A�.���C@VºC`~�ǝ�՛�g��1z�R|Tf[�5�0�����=��/j��3�9ٗ�d��b�r�m5�ݯz��YYjiސ	�hsٮk;�=Vd� r��ᵫx8�i�g�\���I̕!��WG]�6V���y���Y����a#�jy.�=�L*����x���ގ/��Z��<m~��m{ۂ�![�_�9V	�(�C��F�/;`�&N��[Y�:�y�T�]��e�׷���Hx:�X#��܇�1��n��A�I���O�H췳o_hnŚ�n���=���5�-����E�3���k�d9�1�[��$eetyAX����=�������q�Q�w��'�W���Ģ��w3�ݎ�
������֜���.���#���z�9ыލ����fN���I��-�ge��؂�cT(���$�����3����@�y�~�����u���n�ە��q��0\����#snc �e������9�g���O;�����7&w��o�������}W?Vc��U��M�y��pv繅tNu|kϗ�w��g�����ߌ���!V��AO���Ǎf��f�K{hy���2�Ǻo�}f�;F�2��O�3�J���W�Z������W=�ݗ'-���E�Xtv�ǋH��$=���o`Bǹk��a�����\����\F(�3b���{h7vo7�E�~�|��j�	='�VM�y��ݞ���r���9}T%͖���]xc�μ�^y?TV��x;7�4�,����U�hl�*���w2��kg�Sޥn!��H�y7�%���ٳ]��X�<�b�f
U���@ѻI�܍ڣ�j��ZʽM�c�Vڕ�>a���T#�;y����*��A�r����=����8����۔�~�p�#]��{�:�	W�x�;�$�dX�r'�50��sTƉW:E���]�:��gw<7��V���N�~�/��j�^�.��Gf�,�!L�+�j^��eOUv^��E�ޘ�̜u��s���������Ej���^������~�yE��Ky���-ULk�3�u��T�Ƚ�^{�������{���=��]S��<�?v��TG����#�[����U�d?[C��"�z�f��OPn<i��]S��{���.��=��^�P�b5����FrSʭϖ�y�$��jzx��d[�6^�Gnii��l��H'pע�K*����9�o�ǜ��ո�2y����v�����n�����'q�cM������W����/DKu��R�՞�o׼���\���}����^�o��ly�8lֆ����xL.���a�1��O@˝����ה,�l��@���h�;bi>+ �=��{ꌨ���܆�J��
�,7o�4�xr��p}'`s%�]u&�����=Z����j��ˁ�B�	Xɸ����Kئw����Lһ����*o�������*ܜ��)b�O�5��mʕ, �Fm���h�Q�gu*�P*I�2��Im3R��o��nlSNIH_����3��'b���"r}P-�N4j�0�hH��j���7_��Y�h�o�X�����]K�Oj�K4����@���������`Z�M=�G��į�@��Jb���I9sV잜q_�6���z���	�?W�:��E��ϔ�@z���\�����=���5Hll}�5����{	�O�Eϰ�4�x�k�bZ$Wo)���M-���=�~>7�m��ܮ^����⟗���Ǿ�W��=�In��%��Ix:�o�2_S�P^z�<�ҽ�P�9C���3\��W����a��5Ǵ�"�����v�n��?U��iJW���d���]���缧@)�[7�׾�y�z�:����1�v�����%+�7�)H3�m?qҵ��g���T��ej|�Q
�om}�{#ͻ����M�o�~��W�1�u����J7�DR�-����h� n㽾�w���G�H���Y�8{%�Z�W��"����{ݵ�y{u���˵�~nP⠍b~���N]I��{9Ǒ{m%`+U�t����u�[ݐ�Y�s���y᧗}��lz�q�W�#3������}�:����o+��\�Q���3�y����ݪ�eOB�y���OR��n���w��I=Q���O�U/���ɐ&m�Vp)z�����f�g7��n���L{|��k�y��5S��y�w�sd�)E�f'^��ʩ���ߖ�s>�$�^��o����cȍd+B�6�O��@o��/g�z�{-g�>��3U�*#�W�{���<�w����g�ˀ��i{(R�3C���?ut�ߙӔ�/�Lŋ��U��Q�d�r��w�6�����C�D�6��w����<�7��I=������9�GS2A��A�c�l2���;ɺ2�.��\�şI�Yt��3�^]����K��nw;�cx���h�u��{���
fwu{��;�.g�@��{cI��g�y�rx���NЪ���K�N��.�γ5*{��c	$m"}��_T�\�e�a�ץ��q���
%T�M�Mvt����7�V8Jd#�KF;�A�gi��C��qTgm�Е��]�t:Q��H���@%�9�(�_	7G]tx�x���V%�)�UÀ��i��=��w>N�;${��I�D%�n�Nj��k���Rerg����|g�C��t�G^����M8��87P�����)���p�װN�Տ�P�ޓ��7����+��j���gS\�;|,��~��gxR����f�����D�����s߲oa�s��'�Q���b�cU�Vd�i����Y�}=(y��WC�^l���k0�f�m����=Գ�߽J��/��%�1��:�jzC^��D=kN�"���{<�>��{���r��=���OC׌Ù���@�=T���c�2�4�~s����n9z�-��z��f���K�N�y̬��Ǐ����bg��ob^��^ޭuⵅ<��ezQ���`Bܼ�^�)�<|�>��k�؏�z�H{g����c�j!����L��Ǫ�wh��������e�H��[���[S�`����`�S�Ƒ��	H�7{���t�E�ᬕ2�m�n�޼�_=y���u���S1�3X�+�nQ] �O��i^=ݓ�6~��on=��;�v^��G�2,�f��v�[��n��"W9.�iUs�1�W
���o��t����4�Eh'�1^=��܋X2gP�
���
ck���u]���Q�D�,�vٷ�G	z�p�l�5"(q�a�ܳzk�Srj8rjܘ��%�ݬ��|��ov��z+G3{�Z�s���IF|�b��ig���6!��e?W�Ȃ�2�7��`�2�X���P޷�+L��{�2Ù�E嫎�u�jIh遂��b�
ux�T�ħV���5���Ѐ��E�nm��nmV!�
&��pdܦ�zw�5H5m7uJ�M٣kz�\�n�.�Jr|c�%S�L���t��_;Wň�;r؋.,z�@��(k���v���$y�2vW`�";y�5��d��K�-�o1����;�&2~u����luѹ8��V�����6� +)Kt�J:��١�fĞT�w7t�X�urw�5����	����:o�K�*Q���Wllئh�w�9���(�y��+�>͡@���3��/�[�<�N�e���*��BA.t���Ӻ��&��c�ot�C��7���^4.v�^ӫ�u�7]�_lTc���y3�@8*+�/3]��j;��O��D�u�g�^�\�;�R���i�M�B+~�4VE�\���a�����zڪZh�k۬�ot�µ
�REj����/kSϴ��f��V�l��4eYy�ծ֤��\�� ���ܾ��&��A��h9ÖRK�ݴh����`=���u-�|���P8u�L.@�����p��4�e\�N��i����[b�ŗH��tNz�cG >�����+:Պ�u�7z'���3!.>)c�;wj���X���e�:�L7�s,�/| 6����jv���4
�|��J$�{��rfʎ��E��S�ʸl��2��:�>��絹s�#��d�5������b���[͒�fᫍ؜9�t��Ե�v��Yju*F�X4s\�ն9m���P�N�@�S.�kC�]�����9�����қ/��C��=�Ɛ���a�T����@HϜH�6����A�{�@����["�w!���9˖��W����E��b�4	GL�N�k�t]
��+T/jLܦ@S�LٓT��ї���.n�l�KYܢ1�5���C�u�W:@�u�s���3��4�F�T�M�����:���5�aw!�d���eʵ
����g�.�E��l3��T���޵
 ���ʌ��l�F�����Z��qQ�4OU��^(��*�{���!����{&�W+"硣��C���{ӓWC�к��u����&--�T�O��b�2����ڷ;)����6L6Fs�nvc�f^m�-��W�0�`��	�-DQ�*>�3�X��Msj�h�X�m*Z�'k6���y>����_X�P�}Y���Y�x����F�����-OL�n5z׶�҈���kVZ�T�vVP���{��D�+��JVzL��8ʶQKj;�FeaX�P�SJ�K
��6������iu.�L���rffnڋ2^�湬��V���)���MuxS˴8"�keV���KNl*f,W�W*^Y�l�KK(�[�mh��,�����m����z��lV�-E�͈�b>&9�Vd�����]J�s��[��-��ik+oR��YV�L#�*Ӵ��ſ�YX��Pb����}R���G��Qx�0�O��6��6�s�a�%�_n�D`W�ˎ❦����
[Z5��־_��d���毜�����mj�\�sx�4[n���-��d���mj��h�^b��Q]R�B�x����痌��5(S����w,��D��R��'��_H޹uU>��fpH�#�@�;>�]��cW{���k�	�A�}��:�VWt�v��ts.����Y�HM����t�tR1'�WҾ�"߲��.6��1s�T:�\����'�~����4PJ�5�y�(���(�N-�䴕wH�Ϋf�UUf�y6>;�hhގo��ϔc3b��q�%�x�;qg����~�N���O�ۆyt^e�dt\;���?��[�;�l�Ck�It�g#�G���3*���n�h����Av��¸b��7�I�Rs=�~���?�}u���樂F��@��E�|�5���6�Y���O���9�q�� �wYc#lMS�<rJ���g����*J�������<��e���YW@����wk����S�#�?�z���]M{�K&�
�[h%�Z���1�g�@��%f���(7ԀF�{��~ɩ��0��r������	�AP/
ހ&+�<��)9[[7���{��!��]�N�{�f��N�i��k7{ퟭ�Z;`m�#��|��W���\Xs*����]B��U�֢nr^&�h`����֬�K�߽��g��c�}0�,��29�Ft�;O���tł*���6
�y�l݆:.�D�N��QD�����þ��t!�|�:�?�O�ʿ�e����h�����A0��<Z��;�oy�7�2"��-�/��;�̾�AEe��9��[wD���-x;԰��v u��rC�{�2Q9�Y ]p/9�f	9�T���T}ے��/NRip�rUӼ���gF6�iy����6�<o�G:�o ��iR\ͧ��I2��S��u�" l��!�o�RđC#W�j>��K�޺����$��lF��/&9�nL��`T��Gf��x?����CB]"nbM4[�ۍ������S	�y.�c��!��\JY���R��#��@TSW��?9\�$��*#�x�$V��a�l�Bz�}q^����q^j�m~��f��is�l�6�(���WP��[�}�q��n���#����h����H=�K��Q�zb���� �c~�p�N	�[{J�~)��g�wf*>`0Hu��d{>Tz�1sYC�I��w&9�l���'�j���Ma^j=b>�}�'�~��6�P������c�d�c�n��1��A�	w-L�ĿA��[pc��O|�A�&���_�D��A15E�����-�g����2&�klŤ˘���Tw	�$��z��7���[4�%u���B�c��ѥўU��Ţ���1�����@��#����Y(j ��z�Pe/~N�j,3�~���zZL�:��z��{�%��x���v�U����]P)Tm���u�/w�s��A��f(��+(V�*�Ի�j��ƾ5mm��,R���+) ��˿Zн}�G�R�����s��ϳ��'K�U�����U�M�RM�JE}�	�k�R�o6QM��C��Ea�t(<� C�fp,c���os+}gv+h�i�[�e���ޘ~�f �Zf��Ί*�(l���Ǥ<l�U(��Xn��A�ml�.z����v�V7�+���U�R�x�y��0^��1A���4�N42L��fo)ӬY��n���S���et���'2�����Au�pN\k۾�i�� �|xbv{$�Lk�Q|�%ݻBu�&�p�­��^{�:>ePzv��P�W��a�/]1���-�<F4æ\��.Cw=yO5,OHE�[���-�t{�U&9T�)�L&\C��rP���>|ZG5�H w��׶k2zs�g~9���%�3^EQ�F\W�Z�a`�$7pztC�h@�m�v��N�|h���Rxn�kBb5��	�M���G�=����Jm���j;�e�)�aqk�%��Ŵ=��\�ۚ�l��4�a�$��������z�Pc�[�����7��Q�� [6�U�$��[��L�<lÑA�9Aq� s�*�2|�	�����%��:�s\R�c�߉�c�6�J�~_�8���x�D��`㈌+��197ƾ�����>���L�|��2L��UP60O�(���Ѵ�7{]nhz�m5�^m���;���^�HM���a �*KM@w����ܤ�gl�#�wÂ�ԓ�os��t�i0��@�aA��mgǢ���ΐ�6�Wa��M<<��j����[���y�-E��t�"Q�],��Q|~#c�P�X��H%�5 ��K��"$J�.)���"�a|̼}A��.�1?]�FwW2t�')��ASlQ�gO^��U-��czߔp~~���3y��e���� !5�7_n��CV�n�>*m�ZD�.���y�;�[��������I�G|W�s�
���!Sܸ�3Mժ��kg�M)HLht+\'�;	麦��Ց;�x����Ft�6$�	-υB1��P
�VMo���*���,��b۸y�'���G[u./kݦ���k(UZʈy��E���#vg�h;5["�.c�/_���f-�3�eUN��[[��;�*gSp�P�ɔ�p��E�.�m��X�J�Ɂ��醕|M�~D]Ĩ���^���Ww[j�(2�9A�4�.��9`T�m��UZ���I�����|j.-�Z"�w(5YI^A��j�͞樒�̧km{v|N+��;8ڗiIOn���_�G7RR���80��)caT��o=�C��B�x�@?5zz_��v*��|KׄQ*��Oqz����|����kЖ�JY���T��WVWG]OK[8��c�1K`�?���͏!@���=_�|sa�����b����Ԧ�A�%ȍ�n�mX�}+Q�����!�!כpe�P�.�9�,�ػ�=��x�W�5�l��c�s��3�to6�=�x;x3{�w["V��[#��U��,I3�7��!���#o�~2�ޝ�T[�:ԲL9�ֶ6&�����7Li���Ij<�.�Y��CA=�,������<xt�U��kw��U�N��4G?:{�X_W�s)�,}?�Ua�� G�̃��z�Z�L��ܑ���y���㋣3t�*}��&��/R5�cU}�c�L�GdtP5�u O��LB@b�����7�D�qw9���H�U�����eC�����dc.{s]��(Ur�3��ٗh��ٍ�cX'u���"ڛci����
��f�43�4�09N�~/�(�H�%M��[/��!�2:��4���֗�I�$�s����&y6jiX��������7��m%(6��X�u�T�2�#u�=��|���{m@�ݺ|���O�b"��!e�o�N/�]nY��~�W��	q��el̐�[��%�^�,�m��0��;m��7��� ��X�
~W�zE�O"�2�t��B���^�Mi�f������ֻ�!�\:��@YN�`��`o��EϽw�~;B�9�?��fƶ�Ɵw6[�|��X�>8�tނ�͡��Og�7�RW���f��6�hn䳂[zU�>� Ǳ��`*cd�X��\�N[&)g1d�2���04��![�D�w�o�&�X[eE��g�	�y��goy��Z�s*��ݣ�4���GD�r^~u�F���l	lҦ�쨶�}͇�W=�*�n�īl�����W�yQn���m��/��
��\1�'�Qi�����ɦ���.�m�0��||����&�\�����������Ŀ��H�?w%E�9������ܴ3���g��m|��o�Z������#�y��-������-3����?����T/��ͩ�	uJ*�rIrۙA�l�[c֡�+H�~�=��/�E��ч�+�����Z)�h���k\2�m�LC���,��}<\�������Y$d�hhu�D(��
�~�ԭC��cj��_��eŧ~P'<J��l�hOi���ޚ��M���vR���,���GD߭婖v7:�`ݝ&��a�g������N7F�1�d>�U�S�3�)��9�Q���O�����6@���|MRc�a���/���E�ӽ3�|0��9U[��Κ�r'}f�O�0���I�E@ �i��Bc��@���_n��t�i�һlB���@�/AB*@��Is��ʫ޸�����l�G����i�T���Q�y&!)a޾i�X��M앚��1�;J&��33S���U��Pyeý4�\�����Z�.,�%�IW+yų�B�w��4Ln���9�㺳����PH�B�<��<�<&R��$�h�˿�e��oTx��7E���������@��M!5f~�U�l���?{�Y̗7����X.����Փ��_�Ι��-�>J��=��C��C�F��'�1�k���n�cw{��х�ķ!ݴ:��j�캁��4�eC�X�ę�O�B~�F�_tP����v���k>�B��ի��-�6ޮb�6%+G:��<�ZYB��*��n.���e
x:����ff��hd���;��]N��-�M�`	�=�b�O�nE`i�;�j��1{z�*�8��2*��g��x>�3��gnY��T1m�A��ʢ�:崧��&�+�ʝM8��hoX�z��7�̈�*",� ~�,U����]� x�^���t���bF֛�>�@>̤��2��*}��W�����s�_��DOȰ���7L�e��G��{��{(���
K�ڞCφv���y9O�]K����vcGHqVM���`�z�ܭt��\ar1ʆ0}���2;)E�p7pk�r�ݒ���� ��r$�,������>�~��S���y��(��y��<e9��u���ɅҘkQL켽�5u]�ڼ@�x�j���37.����@�)�u�8Lin\�T��,��0���w_�7WL�H9�|�-�!5���ǝk�wf��Ͼ���_U�r"B(���׿�������{_��M��NZ���.��{�vg�J�@,ڄ�-Gs��8\p����~e!�5��:�Y��㈁nJ��1 I��S'���S.��,<O{UB��d3ڬ�osC2IO|��˴�~s~ҫ��j����V��W��}��u�D����	G���`s%�5�a{���xhP�����T���W�����5���$Ԗc"�Pq�Da�%����C8#�<�g	o�Z�׺�aK]�d: b����v�q>����UI�9�gu��w�g�e[LO��{s'23��{�Ţ�:��+fI��wAN��:�h"�,ISlQ�`=�}t���`Kdt-��+��3/T{������#�Y���־��R����,a�!��i�VC��oj��9�7��5�ʽ�w��G�#G6��.y�@Y��H�Sn��}�Ό��x��	�ݱ�N�5��n���)��e��cH�۔�ʒ��f.�YDt_���Ǿ���Z�ޕXǗ;k�.���D���L^�D�͹�������t��%�&��$CǠ�3䋀C�(b�pB��ͳbP�i����\Y��W�Q�CKB�V�-��]�l;[���brۧj����+a�v'G�f5w�������=�%�=jP���:����3v�hx���95��3{Qf��	V�הxI���6��n�p��6��>M����_�#��XD)`# FH�X#�{���~��ý~��G�>����U)�g�U2.pk��Sl$��b��_[�����pc&����n�j����*��iݮ�}6����K�ߢQ� �b��LN����8��.XE?+��j,�p�oX�h�e�����nj� �P�	���}�ieINҕq��-�Y��iPIgTT��K�0��3Wq��6�s���S���a���D���W-��r�Q*�:w%�d���n �a׮��=YU�E��j8�Dj(�r��o�u!g��x�YԪZGw3<nD.k�yj�	�@��5Bd�3�L��R�m��x<�C���D���]/}�۞\	�!r��m�i8k�¶W���<�ȵ^f��U�^$\�ý���� kC��]���]�A�4l���ᅡ�k�y���7`3;��L�q�ɀ���ק�ܳ�j��x�2���>��&:\��Gn9�݁BB�/C���r�c��F�o��
wHȱ�f��z� m�����w���v�	������~9�|�b'=v؆�wa�n��-�KH���c���)�տ�s-@pj�4-Su��ట���v��t�w��Ǧ�UK�e�}�Mf�f��F����Λ�ݳ
diƔ`�c��̳K�)9W��}���AJÒ�Ɏ�S(8NS8o]t(���I�b5��^>�e]j���w�]��=�~�}��#1�P��H�d�1 P�X��ks���S\`�Hs�Xk��.���^x{�Gq_�V��YK+�ye�=��:�f)a;møH�CR��a�;��@�]?�T��I����v��q~�crV0&��Eɻw��U6k�^�HR��'��[��V��[�#��$F�[^IN�'�j�dG��B2E2�mO�ȗOh��#�:��zh�狠ŧKV
ʦ�,�k�ʶ��_D�;ݻ����(�]�}8oQ�;���-7gh.���@���?r�NV���M�������}#2ِ ��5������7�=���G�ܢ��ӽ.�Y/�W7��P��0���ӓ�]B��35q����Z�**����z�-�W9/[��ό,G&�H��k޸�h�θgj�Qkw�@���B+e�":��7��F��{�`"��ec��f�
Ѵ=�?�3�x��L�v�4b�+vm7[��fj3i�M�m�)m�%� ���T�X��瞎��F�P8#����6��{ޭ��z".	��[�e�g���^���+��=%�����=c���TM�ZI�d��� ���~��#~@;lh[�걳��kN�O�n��q\�'�N.��X��{s4x靽�<���磞|����I� <F��]��"�Wy�L8Mn力)�r�����N�ٝ&�ÙW|���S[�s��q�z�aݖ���f�����#w��"�7��v�9+R��p��ĥ���|��-4j��]�V��
���]�{�5��|a�{@�N���TM性�K� ����sd��TԾ)ŮD�#S];��wn>��a<᫨���̢z�V��4b"Q!�L��IJ�b�x&�wB[Iu�]�G���Iߒ]Զ$ifXs��[�`X(��C7R\s	�Iu �cw��'Q��U8�^���2B9,i1gE|RG"��j��5%�Fo݌.ڹR5l$�a�Dx+ppu��V��Ϻ��A�s��ނ�Q�TP��UKŧ&V
l�~T7X����І-&;���뽄�s&n�c��(�� ���.�����*�y��r*�KY{�r���>\��a\��U�FT����ty���<�Z�"a���Vs�T�p��Zޘ�ҳe�&���q�����H�%���C��ٹp�eҫ�E�&�L�J'ΦQ���X4)�-�|&�7��R�OE�"��)�wݺ	6�~��&	I�\��Q�#�2qpۺ2�2�����%f�}Z-u[�кn�����/7m�	��f���+%;5�I�t@ᆺ��������3y̚eoa{���D5sc���~6튽!;���:{}�|�{.��ދ,�/d*=q�B(��ݦ�-�/���{d��,8�m��A��s�����0E���#ǜ� ��%z������n�۸�$�ԵW4�e�L�B+Ko}!ŧg`��S{�eb�]�\U�9�	��ΨS�a�|xV�~ChE�f�܋�]�`�._I;'+D.�
���6�T���S����w�uƻJ��Ez8�Ƴ6���Lu:�	bt%�p��^V�YK��6���lP>�g֯z��������.�����PJ���1�[�q�Ϯ��\�i���:!�8-�%M]�]xcC.��������o�C�9g �}0O�d�>�yo9���+�.�F)�\�Wl�d���U��c����׮�c���[���U��u;rY��m�X}���SB��v9g�k�rŰqu��|������kV��k2��J��3.��o�cp]��{V�=}�Q��!u�)���0�Ø�t��	��/��N�ve� �uj��a��)3���<�Xa��Mm�fs��b�e[�%���]w΅k��_v;&N�]�v/,6��"�ޝ�J��a����gpK U���N��8d���vF������lV�XlC��;�t]�]F�0u�y�N�虼�L�L��V:�*x��pb�Ś=�D<7!�=�Vt92���w/C�%�c��Ә�&�wLǦ<�5b�]�l)�x4�a�y�ͦ��|��v�H��S	�O�����%pJ�T�*�+���x��j4�R�n({OUw�ml��Do�y�h9=�'64m�\���ad�mb�������#�+�VkK|���^lj��J�(nۋyf�[{��kE*u*
++#�T*sS��4�z������ը���Ѫ*6�J����b�X�,��R�����6�V�M�T�����ӎk�VM��SҡKNR��X�Q:�Z�U���[j2�Ҽ{ǆ:ִb�p�5Z���v�sk,֣ݳ��u��J�3+�U��6�amKy�-]��r�쉋(�r�}�fѧ�������]�mh+����^ژJ�ZRĕ
�(ݲ�ۺ��aQxZ#�aS<�8&��X�4�v��ex3��*"궥�J�l;Nb�VU��984TWYm֞p��7/�pZ%�ط�P�"��&A��lq���k��*�ƹ�bZPQ���Û�VZ��#8$�3�ɯ%�᜗.k[R�R��9x�ɜL��\ �!�9����yms���X�)�x��o!T湨���b�+�T���
V�o���pχ�d�JK}\�u��Fs�T�kj�8mS�Eѽ��Xq�S�:�Vl���d��$>B���>������ݽ�Ϳ�?(�X+,@P# ( �������{2��i�i����y���zO>3ƅ�*����	�ֶ|��'�A�~��-�gӏ�d�����14�����Ǡ?��A�<*Lu�,���F��M{TJ�[q��U��}Q;�%4:���a�0��� X_D�!ąq�Z`s#�{Ub���ﱡ`r	�΁�4�Ar��XR����"�"m��f�NM�P� Xs�_ץ���2�.�ɍ#r.��(�w&�6�SQ����#���מ���ȉQ�#�qm��e�O�	��6�*'�����^>�� �&mtY���yͻ�\������AaX�Df����~�q�<d��]OR��-���t�CP��C�cr�o"�τ$���(t�g��z��q3A�S]�F%\���d�UDub�Sȫ���JV��C�(���Y�X�WY�6�L֥�b�á�ǫ�X�����$�C\ɘ�e!��1�Qܓ{����!�S�Z�cdX�y�#l�^!_oe2%�G���o��5�/|P�xX�����>�v��@���1�R�W�ٵ}�4��=wof8cj=���12�vN�7<�g��Ͳ�>�<J��s���g�@k��/&[Y��u��7�l�j+����*C\�w��;���Y	k�__8�@���B|5�kl��J�x*���G��m������I"F ����I"�o�a�y�����x�%�N)��D�|9O�6ؼu�r7G,������_2D�R��.B~݀C5��0�*U���� \`Y��d'�Q��-:��"�C���*���f�c�����Ƒ�s�\�&�y\e��?@�8��s�A��u�+���d9L=ggF�iىM`D�Ȯ|Yݏ��KT��{�����kuLĽc�?f��[�2u��\��3.�y��	]l��"��q9�8����V;;0�dls*���2e1��t{����*�?��q�����ҫ�>����t�U>}�f�[�0��Ig@����� '�s3��E2��-��y�%f�y,���,����j(��Q��@OU6����H=�	����
��'���4�:$9�z�ܧ�l�Q��?>R�O�m8��1���}z�RZ���h�ͥ���������έ~�ճyQPw�r��:q�Zi~`�9e;���c��k��x��b����T����ܣz�\�����;uV�h�|�!�é齔�����c��{�
w/c�J��P¦�4�6Ο|��w�D��V[+\翷�
PL�j�a��>�Sa�d���*0�X۩n�J�oBP�}CI{:�)�c`7y��9��g5�D�P#�1Z+j}�'4� ��l��4�#R������{g+R�o-�2P'���ɐ��p��U�5��{,�O�|ݿd��,��,�Y���������9h)��>?|"%�s��Y�1R���ۚz��٫�>�����(��/܈Ʀ�?.���u�Zb�~�#Q"�ʑs���W��xԘ�R6��1��T�׈Bm"Z�.J�FN���m���Y����;��e�&��[[X{3mC��x=рc�s�eJub���V'�"�'��7y[ T1sW�(m�g:�Ey�R9����=>&��Aٹ=���@�O�w�J� �m0���7+=PD썯Gm�����Ss�t�m,���M�@�#�k�Jj�t?M<R��7/c����"`[,z�4'�=�H���S�Wx�yߪL�yC]�p?ng/ԅ6&�֑�J]�T���C &�/���p|��S�p��"p�� �C�=�U������>���ʟ���?�~Zk�C_1nv}0ޢKȃ�Ur}�s�b�����1�޾Uq֜�g+O$��
��9���ޘ���TZ��'}�2B�� 4���f_�dMr��pca �sr�P����Gk��cAap���}�|�#\㧆��՞wa�)�,g��#�Au�)ܤ�u�;dF����/E^���U�^�f�!6�aA��+���9�e�	��P��5���k��U�5�gg/#���.-���n]+��%�^��#f�%�:�����ٜ+9�<�����y�Ϟ�{����@X�1��	EE!��~z�����-M�j����݋��]U�w�q�֢E˱.���ߦF���!��9�Vu dA=���ޑ����γQf�����Z�m���?m����k��H'G@z:���Ꚋ_V��֒���xZ��"w�9�|jȲ�v�l����s��3"��)�O��Oz��*�%���w��c90Q�7&N0|�,�=�ƄC=�٬[�f��<�[�k�^��8�����~�o <��Ë���8�V��2N �g�xhNS��c��s@�ʨ`��VU�
�k�:aq�ܝ�{T��^�.��B����3�I��D�j(f���������>��/C�g�m��g�Ua��L2x�%)�9Uך���⋈�iw���|ǐ�H��� �\��j�w6e!-U07�njFe�d�j%�i+*�x+�j�b����n�ngv�ߚ�3���s�z��1�^��vkN`����x8伧Z��)9��)��
�ǻ��k�O�֢������V��]oC��-���9Q>	�FdZ�o�Di�=.�f�]����R5,a�Ĭ�y�����u�m�c��j�Rg�dd��d���xj��[����6֘�ڔfR4��z���ȩ]����>�W{�Ŗ�ݨ{w�z}%��C]��sS���(�ܖ�k
s;_j콑m"���}�����d������S�6����{����𰑉
!��I@�8tn���n1������j��s�_�!��`��} A�O����,�4�3��<���"b+���S�;��C{P�@��:���%�+�ЪD7qZZ#���R�74��&m툤Ę��c�6�X˚"�8]�v@�U-Z�Iu��{���tkk}u�di%@8# x��;�nN(�h�򾭞n\�R%>��m�8�r�4��>�,���&���#&�
a�Y3�Ĵ��\wE�b}�<;�B2=K�r^ZAff1��л%Ra���	�Z���3\���?���/Ӯ5l��Zj�-,0�4����i���ꍳ�i�FE1�k�(mF!�f1N�m�fo�K�i�� hD�h�D���c�Y��X��C�����r,u�w��ׯ��xF|�VС�yA���ԡaE�!|�{M}0X�W ]]^칗�uW��M7�����yxlAs�5{I�DTo�����^	��2N�0���ȈQ�"�P�5�!�j�^!]��rE��}uw^C�w���nX}���~����/q|KV$�}���B�H�!~ �1��.��/����1)t{ V$��F�?�xlM�o����Wޒ��,�ܸJVn�x<��L�P�SEj�EtZ�v�im�6�,�����{^��oiz7J+/��]�<fz_���׷����׽�ׯ�9o�$>��H������< ��W��	""b���S|s����f�feIB�����6���/����;^���ѭ�ժ(&u>�B#��ETE���Q��*�m�{��~�2���4�+z��؇�aq�D��-��xu�sf��¡;��K��Ԩ)�&5�c�Sc_��˞�εe~x�C#���R������Y�.Ƭ�avH���/�<x��p�A�֢�Z���Ɏ�n�4�-�|�O�)>�]�(U�/(m���|mwِ�"|�C�u;vf��([-R���!��ن5��n�<�'�e��T�dyY�rf�"��|s��R�z�����̉Ώ�v�Ȁ���p3E�fv٘3���wJc��.���vtkiٌ�քN<I�dcX6+��T�J��7
���D�cm-	��>�y��OM�2㮔�=ķD�\SG�_uZ�Nk���A���[��LF�5L�Non}��D�Jm��P�j�`��-��,��0�1J9�.3��{��ʼ�=�+��K_=�_�{�2��=��[̹�%/�יU��z�k�t�N��&C'}=�͙ ;}<)��Hz��%rk��b. ���[�h�wP:�ZeB+�]z'��Lz>�ba��Ɏ�-H�~�o�����TS=,m;tn�ܵ���>4�;�0���%r���*[s�m��L��m�����������o7��=��]��!7|���2�"�j9��MSkP��]zS8ns�Y���:o�6E��O�cx��wz�-Mk���1��L��<���'��g0N�F���/�{���oAU��i�3;�M�����j�Dqx�,+n�n֠: g���6{��>�T��sr��D������]ѵb��*�]|c�0�ے":q���)�
�m{j�N�v�N���mE���6�����ɿL�^�]��~��}�+�5ѭ]Mð�}�%;�;�OWwUj� a�6�6[b銢2�=r�:1�C���uZ0g��Q;(�u�R.~��8|�Uc��I�{���h�_��?Vw�N�u�x��Gdb��t+U�	з(�1��&��>Z��chSQ�n��0(�����8�Y6�Yr�XЋfR��K@v�7�����s�o�띛1����Qn�y�}Ng	J��Q�F]�`�u�#u��D̦;�*��r�)��]c��``�h��Ҭ��[x36,���ӌ���l�0z�A�����H���NXX*�7qSM��N?0|}F5V0W��UwKS��.��	2Th=�R��@�<�3e��
���ݝ³(���z����̵f�vb��J.�[���m�P��p&�j�]/h�]�3��źO^��	�ީ9���; .��߬�85�̺}�Ea����IR-UL+�m��YFpg����� }�I �I Aa	�ׯ�=}s��G�Կ����3�vcϢ:hN������<���6���Ғ��E'�0�ܡ2�n��͌L�V;۝��q��p�����M9�]_�����C����)\w<&�ɝيTڈ���m��	rPx�m����$��FB�^��+DXͱS-��1����V	
m�E��#wq[c!�L4�p2W(�届`��j�m��z&4��P�yn?����
���R���-��R�ɤdޛ����}�(�{�J��R5UkW�k�c�3�Ѱ��ޚ<B��]Q�:E�E)�ؽDq�5k����`�[7�����w�0v�Mz@�rѾ��OWmj9J���A�ہ���	���Ǉ�L'��
�_��ۘ��ӂ-c&��E�7�O�����u�%o���u�^�;B�d�;��0ϱ���|𓞿e{��H��5f��*_�l7�^s@���x���\�ZIG�L��Ƅ���c'��HQ�*�]����^�}O$��v�.Љ�h#.��|QǠ��t���zw�C����
.�|��v{Xr��_��{^Y)G�m-t=��G���͕�i�����;�H<'_)YΆ�%�����^��5BC6<z�Sq��N����u��K�wp�>mr�� S��/x'�i��X婟�����A�7$9|(����lu{�v��ؕucj���B�@�@�w���{��=}w����^�o�uc�1>�*X�	�|U�6_�e;	�(���zw��!��V�᥁VY�ձ���B^�K���*�+�+^��2j���M�
ʦ�K+Z�T�<5���M�/+�f<|�q��|��lֆ+d�PM��v:$��1I�>QḮz���#Z�BxPn�S�x{d9d�zq��~�/��:J�~��#��f��� ]�|`jr�C�:#T
94I�t'�r�>����sW�<^�
��w�� �Z���?-�|K��E����<��
;w�Q|��̃��[��OݪA.�\�P3��+|x��'�*���k�^~Z��f3PW�7_�0�6�Q���������k�Y������B�pF	u���60�3*%mq-0��K�>����j��&^�˔Ҝ�� �|��I�j�H�~�2�z���kv�s0^y��& �O�}ۋtGD�L5lO��=����q��W
8�`�Xg����,�P?>�,�J�P`���xW�&6�)�Rz��C�tbq�F�1`���OJ8�z�ו%�N���s����k6uH2Ӌ0�����?fF�k��ݮ�h9�����B:��A��.�TSݎj&˳u�̓��m�t>���f�uM�Kq��bn\��ped�bvF�+;�C�]���Hu|�%	Q��vļ��t��;/�p��G�*)���>��������7��3{�{���r����؃��t�4;���^$$�y���Y��`���}ޕ$��֦T�-��`���id�UV�^��Nj��t��U���d�ꂠa_����T9���gB����m]SL��ԙ����;�i���aw�2���X�J�gB';
��&�ae�1׉2n�Qw��m��^��l/~��9�(Ne��1�`a�|�-��2�|K�_[����n��Շ��s׆��пÅ��JT��/X⚷a�&aދ����lA�|�j�w|���K[���1{��N��c�����w���M��K������	��T����c4��������Ms�gkZ���,j�6P��a,��r��:��ڀ�O�At���j��j�=���-J�b�e�1��nmk��S�"��x�M�86�V�J����.cS.��m��@�:G߁�<Oq�݉PDY�X2iC���V�}�&�#���e%G�ql^=C�]Fk�ܜ��$��J�&θ�"L3��街��`y�h4�� �{��7a�\�<B.��c�p���5Ctm͘�:�}�|�Pc��&'Eݺ���̬�˜*�p�R���-꼥��k��eKQ����>��2���Pf�t�O֔�,�Vwv��A������J�F=&��۳�(7��9m=�)㖅u���x�ndj��2I�P������7[N,��˗�{8ku�U�>�[�' �5Ѭ�T�nV�Z9��T����ۚ�mN���vYڻ���
����8��NT�8�S��ʅ���f��xUy�^�˼����оcB����ؤK��>o�)����.Ճ�sq[u���9�2X�E]Lܑ�� �L ����4%\M��,���g7fѢn1�\�ډ�Y.4v�cls�����O.w-A��z�=a۶:<�U�¨_M�d���C �-�ۏ�N�O;���mrulN2J�pu���T��}q�]BcW�Ιǔ�i)[��om��{k�@iv���={��[�PhLo�ػb�����Î��_^����tL�[[Af����̕�#.��H��A�1aS��}�7�[�tSB��pn�0<H����*r�`�v�W�^\q=F���P���n�baJ㜎ۊ�V��Q*�a4.�C���{��R�4��-n��3}����d�.�6��&���������l
��ni��)�ͣ@9�K��sI�=:�yOP�����̾ou^�aݸ8M�3�A�c�845�+f]s��Te�u��[m�k�'�ܖ�rm�t�Q��h�^��8i�:!�Ɖ���&f��Z<�<��pi��Jʛ��d[�;�ى&��z��eg�|�b�/%;Zpb��k�Gw��Vj�P�x��k�,t�w �]����G~�W+�4	e)䓉�q�kǦ=em�Fm8�:t_iG_-��s!q���ݩ3�����N+s%�8z9�q��3t6n���\�T
^�����WtVo)V�Ȧ���s/1�N�;�+6�hf�K9�6��&��@�3�j���׌c]H�J��F�Ẇt�3���e�7��uu&��m`�_^PUsP��6qv�(���gख़(�&�ͨ�-f��}-N�w�3��u:t�:�gmq�Y�L�&aݚm2������N9�^<JM�[��y%2 9("�=�f�kt˶�񮭹V�},��\Jz�y�]�]��t�o,d!dV�pN�3Bg3�D�EPÔQ�|Ƹ���A�J�K��!Di�;�Ș9Ǝ��P������&�-�Q�%*�ETZ��bf��j�V_Kj��1nf&<�����imm�|&b׳�r��Lsq�`��8\�<u}��SLɗ�4c��J�h�z48��w%�m<�?��{4��zx��O��ոq�w��h��#�5�ٳ��"�/z�j)Y�r}u�u<�ִM��L�>yz�qfG����$�zD�mu�;�:��l�N;vt�e��w�SL��\m&]�-�y�|��Z+*sT�y�-�.�jf��kEQ�/���^�s�yja�����Q�圞�����|ސ�"��+|����cF,�(�iy�����1��7��{J���5Q峃yl��jsR+�bR�����;;<�W��:�ᨚ�V�G�(���Lŋ��UU��jc� �V���
�sfNۖ-�®tAV;knQV.�r��k��E�h��[e*֊EQ�V(Z4�y��*<J�ݱ�|�z��gZ�ť�)媌^5��melTee�^�:�^�����E��p+ETW�b���%�X�X��"'��"�GĨ��PXڡmR��1�hł5*��;�a�,G��mV��-V1�j�j�-�����^<��"��ؠ���c*"�����<6G�A2��v,���ގL�D�b���F��l|���0���N�X��涖�,Q�j��T�4�y�F"��"�h�TTyۅ��m��o|��56-J�KF)����-_M_[i�)Ԩ�����ԫ���u�Dyk�2Q��d���U�����L0Lu(�d۞�Y=��w�M��������\����/��|�Y���Dr]�{qU��I��Z%������5'���#�)i˙������B�@# �ק����u�ߡ��K���ǔ�;�y�^L:b���Jc�����Z�&[����	��;ю淂�x#L�pR���)��0qz��=��U{�peG0+c[z]���[� a��h�w�m��%Ex������ ���l��BC����������*�8���N��ub���9\`��%Ţ����y�`�YƊ��;�_>��>��G�j�����8����p}\�-aߡƭo/oU��5��Q��Bz�����ȃދ`I �y��?�~i�w�3T]
���`br'{H�x�i�*�5�@93���1�o\k����jKW��IQ� �$9ٙ�wy^uժ���:7��ss�j$�pD��>���`�@00��� �������=�Z�[�vn$��ey��o��tly�fO3�a���h�n����Ӂ��Ǡ�3��^T�]�{�W�Nm(`�)�}zهbmfgB>�������x�<L+����d{FfVv��Rt��BG;�i��*��7�d7��z�#�4s��8r��A�O�q�n�ϼ������c�e_�>���⑝�¢�ͮ�ލE�0~�������Jc�ۺ�<R��#N�B7F��E��P�יY���l<�O�vCŀ�W/�yV�5��z/Mh��7"���w�}�j\u�k4�G6��އ�����������a�{�x4wK�e��S~ ��*	���T�u��*n�n3ex�p����'��r?�N6��W��:޽�Zi��,_�D�Փm� %yb�TCز^��nͬ�M�Nֳe�-���;b�6�l�B^��(d�.��WXQ3)��UL��]6ڲ���s��3�22���b�8����AW.�^��>k��v��yZ���R��
�m��X������:(װ��8�%͌�Q�<*	�<��c:�0�����|`t��N����r".k2Z����+y헻L�6+~4��2���{)'�ѷ��_�3��'�UKz+\*��,�,�H�N���^k���t����_\1�q��8�Q�?�!�>"��z�v\��oϲ �h����	PԻ��ԪZ��@�QEGϞ|��Q�0N�Lh'���I��"{A2i�_^{�t"拉2΋�!�މnܨ�;�X�Z�3T�֡Ů]�r4t�=�^:���DeS�K��������q@q�9f��ژ�1�g���t�l�,���F���؝��M���G���V̧�N�
�|k#���!8�Ki���93�bA�Gm_a���H����T�n�imy���t((���gwi;�&��z\���ֹ��3஛�{ՙ7�	B�د6�a:E���������j|�+�;wm�z �ఖvޥ�0o�{���!!�I0�O=_��{�}~?{�	��폲";��>c�a�HoHj���hY��k�w�r��g�&�х��Yк�0�4'��BB5W�{�����"�=b9pB~�w<*L_4��}�nP�h�/�i�&z��Li�qy;������u��Ls�3�}I��2N �k��PS��c)��U����=�˵lgj�s�/kj��Y��٦� �!vK��:�I��M��*'�QA��x��F(�×qۓZ*�	�SQ�3j���1> Z�O��f�*�mά�a#uNDEoV�\�����eM�f�k��(�u���yRzɩwM.p3]M>�Y6X�����־��9B�1�V�]�q���L��P>�Vn~;pe7�$n��b�*:�[�]f㌳�m�g:�{�J�~�F�t8پ�7M��Ԓ�Ƕ~�3c>8�9����Ɖ�rFWֶ����"��Z�;j%�n����U�8�Zrp�c;"Xko��2�v=���M?#>kr� �|�T�e��	�;��C3m�4+�{i�� u*�PQa�R}��T	u��wzUІ5�~��B#2�z7���|bٸ�t��/u�#���i�=h1�����4�Q��Ob'�y��L��t�	L���r-e��D��p�U�Y�*hi�0��2J��;er�흓b68��I�������`�wb�Ӯ��f�������a����{�x��󑪥�)��1i��<�vr�bj9�'S�F.25�#�x<�;� Ϭ5��{�CВ��:�R�y�S�rn�O?b�-��ɗ�r�4����[���Ɗw�Ww�B�0!���yt[©�-' L��xC���_�=k�N�c���l-�hOV�|��M=��<������y�>NFi4ݐF�#�@���@D/����7�;��$\��/p;\&2��ڂ��&�^�ֽ�`@�d�j�$Yp���=g�I�#:�w�g�__�h�e�j��bv��ܴE��1Q��V���`Y����N03����Ļ	�k+m
1{.���2~_n��sO���E@�o��rT5d��*'�-�/ǆ�󵴇_!ӲXH1l���ȗm���~f�>�[4�����u����=}�8����~/��s�/�.�.���-��lŒxF껇�s��R�PFD��3�͑�&'�|5��mn��$��ġu\)��D���x�ws��%;�S�AN�ۗ����h��M��PD�ҳ",U���E4�ܳoɈ-U��8Im�d��K6��ى�5s-ަ�L��%-��U����7��oع�mM�h!�=��S�ui]��owE�Ue�v�����D�������ڱٛP 92+ץ��Z�W�T��0��U��ߞ�q��}�x}� ��II������!�,l����v��6�ZB˗��w�d�z���`��*��f�*P�ث�S��Yq�Qh�kY�&������{�Q�qeȬ!*�qv5eC	��;.��m���iƯ	r���ow����x·�ki�3�XŨGI���es�%>D���Ae��WK}g	�n�73�XMh�< \��΂5�=��A�kv�#h��J���tS�2����Y�rf�bc�h�k*=��6$�hU�M��Ƥ��Ve�����i0&a1N]T�G<�<ݫl���`��5������j����U��)[�[��7�`���J$W2u��S��[f.�5�6[<t��iO�_%su���v@�8A,	`��+O
�^Ne��᝼pdeQ�	�F�q�S�I���"x��t��0�r�O��G;���q��W��\A,/��mo�/Y�ۍ6�T	��s8F�j�2[ךOX��]�^gE,��7��8����Pt�w!�`�\��r��^Q8i�*��6��;m\5 Lf��LcX�y�}&��y�	v43�39s�����bi��P�^&��f�k�dTX�3�]���u����-E!���{S�M�����\�۟[�u�R�r�겤��x̾�m�3d:s�pKDe�H���;[��rm �.`��l�u��x�����S��}���~�	�����;2r#�q;]���e�K�}a6��C�l	�`�q��o�G��uL�i_t��^Yq'����3�ޖ	��9P�؅���_���g �~�r}y�Ơ����T�j�l#et��<9y�HC=,�3e�˶6��3e�?k��Y�s�,���ov������p�g�~��u��qpt��\�.�k�ZD�.��}t���bp��W�Vh<~�Q5�!i,�/�oKL��.6�Kh��Z�!)��٥]
ǽX�*��<<��v`�e��f�
�g��w����nu�B!�)�d׵�L�ƿ����4��-�om�,]�ʈy��;�{�K��C�n�j�=H��vjcn��\�2A�[@�tIaD̦;�U2.p.y��.��e�����jM+UY���z�Qs�sq[�E��3�-{b�A�G*E��Jr�ʩM�j)۪]��*���7�����覬��,�[���GK�;����y@�q�\mK����q�s���m�t��u㪸��rѵ˳���ri��
���#Giw�Q��V�Q�閼�b�ށ��`�G���뻹.r�������q���쿭�Y	��Wm�wǊ�uڬ��X�����gfy�ֈ�ņ��B�-�X��T�r.���Z�)���g[��{Ղ�[����{=�כ�6���u�-��Wu�wq��sX3�{Q[������~����]}��_���x<�c�q�I�f����Kȏ��n��}.��ⓨ�>g��ㄘ�������.ڽ�
�P��:�c)KQ��c{��ĪX㍅
�n[*�O�M�n�y�w�Lh+·��1��nW'�v{c2��.$�<*L�9��ܧ���Z2�j��R8�kqj�cGl�gb�o҄�G��;�ψ8k�����A��_Io�E�grvcF|uv�L��=z�Hح�gz�޶*���ʅ��C�pf�[Ͱ�o	��	
0�3c������.�u�@��a���ۍη�,�r_���]%y*`kh�V8Jg������c�!��C5����l&��ʎ��5�u�A��i����
6/��b��<�S7d� u�>҂g����y�r�,�%��Y��C)l�[3&a�n�hJl�e�[O�[�y�u	�sӾ�x��ܛA����w7om:�p"�0�%�\azʹ���M�섦���< ��d�U�6^��a#\D6�'\��yx�}ۛ��V��u�{�㌋�"��Ԃ�k*�煏� ɨZ�d�c�eQ�C����u��o�z��׌��x�Z�J��/����ԏ�P��.T�'i<��a���d��Ŗ7;���N��<�nI���e<nG���30�ӹ�ی�V��3�U>���%V@�\����ͳ�Q��ĉ�4<[�ut�7�{�y�� �a� �ѹ��R�&��5�Gղ��1�#��m�#�]ڭ@Mx���so�����pÅ�[Җ�yՄ�09:����{^�"�hq�Ǳ��s�j�.�/������[��0;]q�m�E]9��2H�!�^��\6A��K�~亅�,�a�D���e�g�a"
i���O�p������e)��Y���ٕ�t�\"���������dz�],�`i��w�jk}�Yr���f~�5I~ѿ��#(~
t~�C�����j7r��1��#�}m�$r�1�$�$�K6������U^�q��j�ܙӽ*��n�G��yr3=���-�p9�������,f{Ͳ�,��4�$�?%�_.[ƾ�3��ߩ럣8нT�aF���ì]=\�N���9�Ds�矀ޚ��{g��82�@1�P��2��/�"�u��S�=�9�e��x����;q�sk�Hϓc��}�J�碢�Br��ٲ<i"M��Q0]�{��T�;�Kœj�ڽe�b�Z��1�#�=˹d��.y(�Q'��$��{㜞�ʾR���X:�Ѩ����!q<
���DZ}�y��,[�V �39ֵ��퇄�Q�U􊡻���C�cz��9�6�i
��l�0�����䂧MU*E��/*u�$��̕���:��$�7��;���ҝHA�������>� =��{���^i�fV�����h��u��ۯ��������ȉAr��E�'��.�wyA�dEU��i�!���H�P�_�bۋ����2)�}���g����/1�ߐ5^�r�(�϶�fs�tD�Q��	>�U���y��\�jy��-��߶��Ԫ��� ��*m
E��%&�nYw����[Wý-%��&z%k����[Q��O�U�/��&{������z):�ga��c���e��ȜЍc
j�[�(��H��l]�)q?Li�i�f�zB��w6�����6�s��)���&\�����,����X�����vF�����-��:t4!�y3v���,�z�4�����U��
Sgʼ����+��k��߱�.��,W����ॸ��.�ʲ�d�=	t��HA���C4��(���E��6ȹУ�
�����'m����n+䌨��q��Lz�_"��C�n��2���r�5},D�T���sR�л����\Rh����ϕ�q�|���Z��$�5R��%1�*�41N]�&'_��!�c'gN��ǅޙߘ�'��N�x/�C�_����y�N�+�11$��KOYV���q顯�qr�W��/�O���T �˾V.Y�f�I�K+��d6�=���c�7e�V��b�ܛ}�h�ΨN�}3�AZ�j�{I�]����[����y��y���{�r�*�͉	�~E�ڔ�K������`��ƳG��[�LF�5	�)��{�en˪Aʻڗ�n�~�.�B�U�qٽ<���Gq��9�1OG��"	�2& }G���y��ʛ"x�
Q"��݇�����վ!QLz:K�`�V;5I����u&��y�^U�A�@�:�U�w�����>ڭ�Q��F��\Mf�.i��T[��k�&[�����UR���캶�>���N�^���|I�@�g��ٯ��V>��npf��wÔ_[�[5�����o{y�k7��tYW,��A���<-�)�s|b��y��0�E�h�n��'�_}83�O��V�h�t���CRH"Gt��L�:z0��ð�����W�k�~ǆtS_|��C]V3mM-���%����C�0Cm"`�_��Ƃ�w�L�ѣ���9^�Y��6�h����sy����N�(�[�ʭ��MS[o�Z&��ƼUЬ{��iKr�:$� P�gA��<g�=�pj�Ŭr�*g���W�``ɋ�Si*Y:����6���Vl]�,��^�&�H������Qf[���)��L/x�ҝ	������8�jR�h��,Ɩ�f��:� ����ܲ��f$r��:(����m���S1�אW77��� �|X)Bye�r���t78��dU�c����N���ݰl[og"i^��E�ר^��s��Z�u����\�)Ѡ4w���x���І���!��Pon-8강ԓ�W�z�M�Eͬ�la$L�(�����06:�Li�ZiXY�֋�Tk-�wfu�i�	��L�LmR]��Go<̤ŧKd�Z�w���++yV��ۥA��u�K��S���v�wo��Y��c�p�3�� 5��M�x��1`<x�,py'
*��������Ùw�x�q����GG;�X�b{О��N4�e`��Z U�Χd�X7����,ьX��V$�Wu�LvjG���ԛ��.R��b�6(�q\�k�9V��D*t���U�n��y�klAvS�ef�b�e���6��I��
�M�BK���8�������������Iո�Ƴ��0Z����@�k�n��>���
��;Cgz�:V���9�[��]��&N�(�\l�3�7��ٖeGX<�rv7�_#��1s�l���k���Q�������pc�m:2���ٱēRTҎjͧ��j�l�f����`4�˽�Ժa�y���-Uj��1F���՞VK��]B�R�ڜ��{2��U�X��4�j�a�e2�:.�YE� �W��L��7`�֙n����XzU'1��vX�i�h��e�]q�Q(�_G-�P%���9�nh]&��K�,�)a��d��=�[�|�U`Ĺ���ʹ�+�=�o �����S���ec:eE@v�EMk3u�n�qb0h��b�YGnƾB�q��Z�S���yLW��KU��kN1�'�k��j�j�M����+a�'X�.	����ۦ����	���q�r�C��̸-6u�qe�����,�-�"�CPJ��֝��͖x\o�at��M#%�Z�,8e8�]�x9>�6P�Q�A��v�H���=Fﱏx��H�y�.F�ڱ�:�ԠcIiu�N�uњE_nV�(2JiA�zphM�D��lm,��z;�A6�V��E��0�X�%�|ѣ�Wva�b�ĵ\\�͚}���lơvUڄ��&T%��*>��	�FlF���jڲU���D�+re��`[�lt��d؎�]��˘�8t�yTE�[[��h�J�:�����5}ɨn�󱬤�k��;�����_�/�!��Ҥ�	���\7��ɷ�֩��;k�ˤ���J�����7��^��{B��L��H{4e^d�E+t"��eۚ�Ғ҂�,�V�9����Y:�mG��y��M�s�u��`���R��� "=�D����T����V��!.O"Q �U�Ŏ����*H杫�:�ȯ
]#�ȹ�#�Ռ���,V���@�NAV	��CRIq@��T���E\�\ʥ---j+R��R�Tȋ-/ݼj(�ӌ�����^�vy>���}��g��R���fF�C	�M�oI^�R����5���_)c:��۷��mUF.j������;<�4[J#ֈn�U���� �}�9J�ne9K�m+am����R�kkUc[��'1V�V�m�ٶPX�����0��J �5<�]bZ�Ǎ��(�;�݅^R䪫&�+DDo6��7:؍J�w9���Q�uAx�*�����v��sV�l�\�"��Z��b�L��#Sl��^2�ڗݪ0�k彲�[�2F҉�u��4z%�D�B��{N%m��*kUm��V>��ZP�0%�Qb�ύ�<k�c��ܹWZ�򙋘�l9ku0"������*���b+�+PQK]�QOwkU#)�ܽs�W�҈��֔s��*#�Tj69^Z]��K��-�QJ��j*"��\�+Q�sZ��QD�ֵEj/ã��:xn���������zX�sb�C��XL����oLY�M�v����NQ��@Ud���&��B�u�1�s/��}n>nv������O�a >�W�k9�w�!�h���mQ���!��w��8!�&!7�UL��]6�"h�;�չ��^\8S�:�Qy0*�\3cX޹v�pYs茂��P}�T��w��u���!Q������Ɯ��x�ޯ���;���rH�'>&��\�;	��\m�3��<��9T�qn�����<�E����E'ֽ1ʹT�~/�<�й��?ލ������,�>��o3**ێ��p�(n*��^�� ��饺s�t�ᯱ�Mg H_<�
G�]q��Ք�]3(�%�?��wq^�|E6m��X#��kk:�KW�@�Q^*9��y�~?i��0N�������)k���	�=�q�/�3ń��6hlo)���t���j��R8�oy��M��$x�mr�u���/�F�B�O�& N���"t��4����:�ϲ;����a�.�B���U��z�C���׷j/`�.~H�xED#��*&�6��ߪ��Ór�:�x��τ�}�z߸M͠X��5;�dX�)�O^s�k��v�l�BCJ�-,���kVߓ�ڃ���K��%漍�/ިώ㭶�5i�q����]%����Z���p����Ε�P���kxF��0�W�3��o`��u7��uZ蜢9^>(-�$�ch�p�{��K;k:�Y�fa
���d��Y�GY��Pf<c�بUm����}���o0����:��E�M~|�4���3u��[Ih
�N�.�ʿr�i�$�O���������m�t��\\��Bj1�,n��_��l�6��!cr�g��|fƿRgD���=&�3��4�\�:�q�A��\K(P��Q�U�5�	�Q^�YR��*L������rDT.�<�-����Y�o5��[��AG�P{�����O�Ufb�-D�m�afmk�V3YU�l�k����w�1�`����G��`o�#i�l�[@�<{�v�膒�L�}1����A����E6�J�_��y��9��˼�+4'���f��_�y/�����׫�m�ჯ�
��ƪ4��L�v)�Rs�,�{Ae[j&�%ο��3�0�)���=	�Ό�N�����.�K�3+�N���Ins�QI�s��@��欐i\�c^m���a��"���lh�j�OW�)xP���r�1i��M#oS�r�bj{��Q�F�[5#�v��:`MFM�R̲Z�6;�na���
�<4'�EH�y�E5v2�r�4�(���]�3��z�HaM��U��<��h�~d�Yw���-�᝝HV����F�5��U�{��0��z	I�aW��8��G9�bP�]a��8^g��A�:�1���aQV��u�p���{Sq���cV��{ f��N����������=�O���@�`IY?�܁}:�����E;��lvc1�sO��^y�{��_=GB��L:���n��b���(�\���8�q��j��8#��xK_?�1^Ǥ赪�Z��ꋌ�1��7�����ΧS�c~�h?T��z*,4'�]�hD�k�sIm�
˷��9�rn��v)�E��z<���8Xs�C��nj7�De|�k�Tr��ƾ�$�QP0����7Ь'V��{"����c��C�J����s~���s�U�;�z���� b-�T���U���=�M�w5�ؘ����H��Tg��(��@�L���$8�XP����f]V�F�N�&�������.!��9Q�ᚧ�g�}�.2
}��c�m�Y@樜b1�eϧ�:�zX�\n�����m���*�B{��J��&©�>uG�G�*��?]dw̧*m��^�Ѕ��i�7����ѷE�c�V��핔+m���/#��SF6O����uI5����Z"�������Z�w]ӌj;f�catǞ�j)>���
��q�.V�c)����P0ֵoN�є O�K^�OLT+���|x�B
U/�]Ese�m:�2����v7jf�z���k�I8A�9����h�4��w2��{��w��j��;�f*�S��SkL���"MN}5�k;׽�㢺*+4T��̾�o��=��x{��G*Hj��_q�[kMk&����E��"����&���c*�mr�2�����]cN���/�q�O�"D%&�w-G@^ޘ~�r������2����l6���6�`�k�M�V�f��ޕ�y̘�Lj5�a|�L���|7�p���p�a@���;:Y9t���W��g~�@sv7Am@�Z�G4;��m�&ƠX݉P��3�v٘��c.:���yz��
��p�ڤ�����a���8+����&0-@�<��PX���95}��2���K݉X�;�j\vިOB�w>5����5�ʇ��?&42��O�ȝ�'���c�&[�3άTS)=E�D�V7<����cA���b��^Mq7��M��zVjȹ[�knzy�O�!睠���f��.i�u~7<��&o^�:���gǓU%�B�`��=�gu�=����y�wT��kT^�N��Q��xVцu���}��Yڧ��/!<@�o�x�+O���,��)u~�
��o���DH��Y%=붸�^d�x�+v�������VҰ>N��<��h��*mA�������Ŀ7��o��m�/��/�(}oo�@�ُ�E+�z�F-�5�	�7I�m�K��n����z�f��iuԓ��V23M���ޛ�pgE�7J�2o	W,.�L�vWy�g^�\7nsF@g��� �ox �%�T�������|�w��� �K�E��ճ����(��~�֯��tb��c�Jw�W�YݓZ��%���{k�S�����Amc�Tʑi������]�
0G��2���k��?eP���v~Ƽ�iԸ-S�Ul��Ʃ��aBSESӀ����eN9��*n�n3eUqd��zp�z�RUq�P����q:�(	O�v�ŬtH�k�d��Κeֶ���W�,�
�;0��v���vn5޺�{�~�0O�@��_��f�oF�!>���mۭg�)���ن���[5q\��bYz¹�.^C���=���+�2��rF���S��9�iJ�M-��V�m���J�����c��e����qg��S�i�_����8?�P�>n�zA�]�`��v�򐬱�����K�[�TS�E'汪9��JV?5�P3�!:�O��m����wpMS��}h��`�Z�����޹oP�r�P����	tp���XՃ����TQ���.��:ww/��}xgݨ_�zD��tl�nz�[YԪZ�N5�IQ�v(���R�O�����^�5_��̐����Plc���{�;a_[Z�s���}E�Y���h�{Q>��yǨV徝��F��}�w�{o`��G�w�v]�0E!BU�F"-5�.���~��t}�cN�v�L�V6�j�&v_`q�s�/�+��">��0����9s��Z�����~���&=�y�M^��֐6w���+Ltt7V���2;��U�SI�1��N<�)n-P��p�c�a��#S�Q$i�5f���ڄ7O���T�$rjxh��諮���Pm��+�z�k�pe/@����O�ny�t |j,�-�;/ӽ��Ũc�Xm0o:s]�$h`Q�����}�^�@\3�
�%���~���:P�/,es-��3�ڄfB��Nvn	j���<r�� ���Ay�,�t�0b�>�^�q�1�����Ϯ�W��K8�N+&��&���P�7xӴRR�m#.��J6j}�%��}MIS>�K���Zf��C�^S�~�M>��OBj=�[�XìjS^�eK'�	JfנU�6bǰ�&�؜�=@�FE��!�5��j�+��|�H��&O�����ЫZ�A�.��g�����gr��\ůz�[�k��Li�-�9��7������1�A�����F5��Q<�.ѧGb���6�N V':�Lh.�ǻJq�^����g���'~V+�#uN�k,��+ߨ^�Վ��(�)�����o>������Y�@�/pa��t2��/��YxIv�<V�_W7��F)u��훕=�xC��6�t�n�xգ+s`x8�xzE��qX��#�e˓mZy�9.{V�ە/j�a8�6��u��Mqȶ��QϘ'������ �=�����+Tب7|;�K�\_�ʮ�I�?q�^�ʶ�����O��>�����{��Μ�=���KC�~�c
�/�7���?rTZØ��E'�¨��e�+�li���[9�?u:��rid���(�V�F�\�ݤ��q�;Ssӣu�^�2f5�H=՛�<�K�fG�(ĞɎ��+t�I�w���V�H�r�;�LK3���TP��u�-6�%6�W��t��?w��}_r�H�K 0�|Dϼ�)��(g,�ޡu7���J��E�u���zSBz�����5�j��8#��,���u�P��|j!�`���m3�B�S=<5M>�CW�ԩq��P�61�U<���Br�@ z��E��wV�}[���ؙOB��]VG�ϻU�b���qx�w��4A��(:�P��K�������B��l�r�A�ן`;G�AO@H~b�fӶۛc��g�C>y˷�r�����D�mA��i�c����-/�2N`!�9�@��D�g�V0/ݙ�3������r���U}�������绮�����Jnf�eL����� �p��w8N6�f.
�卙ed�t�+ch>y��QV���	ri�ɳ-���jbSt�>9Y�Xyة�&eBb}k3+zM��7$glj�g%�y�;\;ɛV������tH�D�=��x �����N&�cG2�o�ѐsm��]�j��(�*��ߋ�s\cb��#u]÷�rnMk�F�J͈���0��peC��l��m�F)��R6x����b��R�]-��}c
�}v�S8d��t�ݷ��%����4j<�'�+(V�6�[Bۗ���v]@4cd���𴆉{q~i6��vι�����^~5�S�9�65	�=�O���J�\]�ʆ/!�Pǧ��8E�*eQ7z�f�[x�Ɯhe��zܳG�Uk�GI��̢��*|��-�kǥ��7��jwF�Ҽ�K��.�K�ǒ�/!@���<1���/��i��J��3�L�˟e��_s51t':�`2g&�zW�Y����mN�Dc��y��E��j0�2r�Pz���F]�K�
-k���,=K�wwޮ���n]��.PD��k��m}%1���a��VgI�_k>�T�0.��7b�C��q>7j���FK$���j���D�'�秨ޮ-���&���dS�fp�SNW�<�3����P���].�iGs��g��r���3���X����<�>!-ӈ銵7��e)�2&�xACyKB�t�~��{ك�SE㴥:��V�J^v9�4�c��-���L8;U9ݥQ��)w�f����{�m	�_c[J��Χ`�(,T��ֵ=1���p�AZ&i�Dl��`�:R�R��f6����S:���`1�!�����=}_ǕI	��0f���z��]K�v��[�I�cs�I���s=ГT��L[9v�wqi��i����,������������;~�u��vV�r�F��F"�����KY��B�D�	���z��%|���<ă^yO��,+n��Z�� �?>Q�'3z(e��m-'��+L�Ep.3�x	ݪ�:�%�@�턾��:����=^�f����g������jv1K���&�N���`��ZU����~�LF��3M��y���jFj�uEYE~}�4+e+�2���]1�LqP�u{H��Ր��r����N�˞%�Vj�kS�С�cNJF(זB.6ބ�۪֩��\��Z�%4U���WB��jƑT�<=�mQM����d�E�8U6���Q�b�k��aM�*�!�i�_��7��st�ތ�,]}^�<���t��%鯉�vjc��\�|ƀC`��GD�L�[*�:~��]���g1�T�4��Q�m���T^L
�h���n]�&\�g�/�����Tg��gbf̦^c�N�dc:z�e���k*��-0��]���7���W7t~t���4R�/�ݻpr��<|��vyQ�b�ʾަ]�j��95�+�K�r60R�N�6��k��v�n�3��d�y��"�dh��ۦ����������$�|�G����0��]&'T�l��N>؝,�T<����v`~�#����=>����<m�6({\�{;���[�b��\s�U���b��X��A)X��%@r����x��1���b��P�._G�OsR�~h�l}��+�T7����J�O~
q}As���Mq�OI�4�)����ORqi�@��N����e[��0�W-�7��r�,^67�W<5]!����Z��\`s*2 z���A���m٦\޹?c��󚸯^Ͳs�1�^����X�_۵Z*7G��\�L`�;�~���7ƣ3�;#���Z�3����p�k�ϝ�����~��xV�zRQk��`d�]Yn��6����V\֜�A�d���n�|�u�/��jw�
5�`������D����A2q�??N�!��)�l��uwb�{���Ω���]���@n�v�Ӵ���l�h;���*`���'C��XǪ\�߫��s��E�1<�EM+�E�Ӧc빒'3z�T��;_z",Ϻ�	 ���Mo�e�z��n�c��[��v��jHN�Ώ ���Qj���[�M��- ���m�4|;��h|�˳�veʰ��������޸����xg:��X�C�A8���Ý��&h�2�ZL�vy1��8
t�>z��!A�z�\�V�+8ҔA��6]sG���Eի��᎕��,!����f!Z���5؃����Me��o
���aĥ\F�m�@�j�:�*Z�F���/6�Q0��#LK1���t+���+hfE÷�r�k�%�nQ���:�����.δ!�i
�akg<��F"�I��<���]{b{��*4�ݩQ+}|T#��D-w�p�hy�[V)ɯP=u�.�(����t)'v��,ps�M�N4<��m:�9�\�*�*O��}�n�gHv��d7�����P�˝ɒ3����Y�J�JG �1�&	tA�ՃY�o0��N]q����=��b����stJ�&fe�Z�J!]�5��pq��d,� �)3{B/Ȗ�+phmQ���Ak+Ggi�Ɛ��_=J!D򽓪fB��|�xQ��n�RRab,w1R���$������[j���Y
+]�ԭ��c��fL��fF7FV,��hs�z��2���N�J�1��՗O�ֳ�^h�:U�(�b��ɛݏ�aώ���p��΍Z�n����0�q)�v�eZ��x��,�(n�ns����s��s_a<ﺯ����M׍�|����6�;�=m]+Ӿ�}^��Kz͒�l0�Vhn�)J���rC�������L�zܠ�.o�@��k)T���#dbu���J`]�]���T].�v ��F�N3	�v�Z�.Kw����"��X�,q�#ظ��t�w��>�M�T�8�r�X=��b̃
��]�Q�2=�ã��3�H 2B�?jV��9�pk�o6�kJo^v��	(j�ֱAM��ެr�Gy���-Ǫ"�:0�$��c-<c���X6Dea�\�û����:�ۥ3��UL7�r��}7u����)�-�]z���7h�Tz��.%j:X�Ȓ���WNˠ�Ӳ �Ͳs�=����Cy�6uk��:�
��Q��$��@�;20"�@ຸ1��5�,���5|x���d�Q�5/;VJ�n� ��=�`˧X�j��V�LK{'�A�J���6�itG	u��+	�{|Q�5��5�ǭ9�Y�J�ϫ���H�9�;K��q}M�q�ì0U���K���Nzk���N�Ҝ��k�6�|u�������ٚ�m���iy˸CսDO�Zu��#��}6��[�&ͤF�9�6�D� rm�E=s;P���́j۾,����߷��+Ƿ9�_�8���kS'c`Mv�2.��ҵ��V��+޻�"PpHt�s3Hld�r��tl�t)��W���۷����%K��g6�z�O��z�n��َH�i��;�H����I�ǵ"䞾lx���־]��56����Vڍe-��5�[D�.9�Ze֔���S�����uewx�M����=O'���J��=]�^k*nk�l�5��u��ֿ	�J�媽jrج����i��|�'g�`��0����m�(��f�-}l�����Kn�p��Y��$rKh�b�6ǝ�K�fJ��9h]���Q�}Z�([|�\�Q�N�yj䨲q����8��
�Dd^4�&�%Z5j^>nhSv�Ƣ���u���w�,���_�U`���k�Ԩ����Q��2��"'��*�������SZ�E�QQ����)�����DU*T�_�19�g�Q�1YĽ�A�(QTT�z�UW�֨�Qh�ה��V��&�U2��l�"�P�.K�^��a"�I^�P�T8R�S��*g0��Ҋ)�.J�����Q��������<l�V#)j�[*u�R��D��P�͘�x��X��mb-��UAu((���/-sPcݰyB����x�{�u�lR�ެr��^��f�N.���[���o1u�R-���{C}�|��|>
�����q��?���9b��B��������u��j���*�YP��J�̞rt�}B�aN��}>��R"�m��r���A�����FH�Y0
}��� 煮��������5s�J!� ����`72ڕ�ju��P�^.�|=#�1d�+�C��5�Jq����jj�W�����{�Rt�3,�|�b�W7W���|nO���~�/��|'m�V����|��{|3�S#�A�s�QpΠ�����&���
���{�/o�%k�қ)��e�Ae��ܫ`��O�6��p��ާgi�_%e��"��zO��T	zX��C�f�.Z�0ʅ���y�qІ����	Y�RWi���1���"b���GK�貏n���b�ɚnŢ�r��۫Xk����ԊE�zB,xk�ܠ�|��A�g�Q��������5!�k���rZK��Je�ϣ�)�(tY$d�Y|Z�	��_u���[2&�)ũ�3�P���۶�xn]��K^[:>x�5��Wb>��`�;?\�FB�W �ʚ�1$��뻳4=���3xo@�l�.!a0�)�9#�u�iԋ��w_Gݙ��c2�F!)A�J�JU�D]�X�j���hM�c�<z�8�i]��`є����L�i\��F\q��%f`�5���%j�M[����ot�W��N+v/7��oxyZՀ�� �q���}�C���N741��4�	S\�TXhNY�h g���5y�sd��Ki�r跴]��'Z,s�#�g�X�`���/n�c��6�qF(Lצ�a�(�z�>�g�gx��p`�}�@����c>;���i���aw�q�l|ʬ��%��e���e�8�6_�d�tTNY�O��Њ�O�G���q��}�9���og��x�S�'��e�w��=��]}��OЌ���DܶP�"Z��It����ޱ�3wEJvQw�r!׉R�u�ת)���n��%����g�AI_��X7п:�|�_:ˋ���Ӌ��{���4���fc^��l��[~F��5�/"��\�.������{�.~�ܵ�c�?(����YS��GD��%�-s�)?_��ԕf���v
!A;C�@��ܥ=άә�=�~���YxpE�(A��L���}&���}*<�����̆��;�yoD�Ҝy�;��Qg	�n�@Z��@�]�$�/��i�R�ۙ�]D��#��$"�t�����v}�I*Mك�xJr�;]0�X۵����E.r�h������'yKo�}�)�5����g�|&����0)�+�ѽdu	�wtܖl���s;�����WV0�q���a�w��.��*o;k�멑�v�M���Y'@������Us�G&Xӑ������{��P��<+�$�J,f�:��2��r�.)�몉s�<�Lm��E��eJc��a2��q����!A����Z�U���|zǦn.�ܴ�p���-j§g�(�@n'�UzhÊ ���Q��`c<DkVV���t&K?==��Ȁ�f�]����[�����6��Fq�U|U�q�7������YS��榎m.�����W��x,$N־���n_sQ߆~+-}�^!���*)�GIoqPđ�ǫY� |��͌�\��	/+f��[�@��������E��?LA���JC��Ykc5�`����1k^��ix�괽�>+^G&W��z$�Q� �`h��ށ�6g�D~i�vz����9���,�cV\�F�9(qgŎ�g�1@.uLW�} ��Bd%�!}"'ҧ���)�&����Wv��4�ne��S��n�b�������hρf�Q��)"��ͷ�K�4�
};/�r���_��&��n+��=�W�:�
�kȴ�����p����M�K�6�brm�'����㲻Y`َn��l�5���o�A�9��EYh}=Zt�m�$�tR^�q҃f��wik��ҷ}��>ݗ�G{���7�3�\��ֱ����Y�vv�Y:�H�i��aY7�R��E�U�{���)wS=�3OFS�ٰ�c� �~ �ߨ�|}��Ҕ�_x3�r�!T��p�dm�[���s_�M����WB��jƑ]�Q���Mp~��f���.,�6m���8�2��`�ex��{i^6���Q,�6.3Ё���I��s:�`&�ϝ�����x�z�9�a�=&��0<<�r��h-���Xm�wv&������'p�mZ,qr�d\�F���T�=�e�_['��7�1���b�4�<컓]���v�}�d�7��AףU.vO	�*�7v��igQ�0����F?(^��#H�K�	��1j��:�	
��^sHy �\[�TS㨤���9�����bT���x2�F���vD��t6����֩P���<2��Pސ/�z>i�*�=�K��Ԏ׭Q�΅�Dg%���e�hīvt��!�1p�0t��oW�L�N���u*����Q�ء�އ�M�ڂt�pմ��I�T�0Tdv`�_9?w��S�ƄP�f�Y����]����h��L�z����7��E�����z�������64�ށA����υ�c�}	�[$0s��u;������Џt]��k���j��|���7B�;d�Q��*�����15d�
�,y��P��p*����9S��t& ���,7J�;[��t�nu����'XqZcs0Wb�"Ѷ"-My�mŴ{���.+ܲ1R�mws�8*�K�\|�[�>y��� �s�v8O����
m:��>�g�z���ק�nZ��v�3N�D}��F��}�W�[�N:�g��C�����p��غ�i�Ōo���jw����"(��#	"��(�T94T�����%����2�<�.1�1ٰ�v؆��v������CSiØ�L϶]�0�G�T����3ě�.A�L�'?yT���c'�,�۶lo�	p%$2���jɐ���u�+lh���{���$`�~����9�TN�j(L/-f���t��0�Ԧ�eC'���i*�N(QFfFV� �T��N���&��v(���zw��!���W4�eԂ�kv��E탌w�'6��u�)��/4��$75��ɶ�VU1J��.�w���1����@B���<�7�[=��	Rw�Ś�V�!��蓎K�s�F���lw��x��{]����vV�SIr�7������z0d�w�BWK�Vl��=�9�?)T�}ҥk�Qi�]"��U�֢nr^ 1~����r�tC��z��0�I��#���\s4^�;;H�J�_��EE�����T���T�y����Y�\j�2��#_��rDZRm�2�y>32n����Ńč�DU�g���܋{&n��X��F�����<��lO�q�̭ف�,x7R���b�bU�>�;��q[�R�W`�����J�m��v��(�bu��N�CGow�[٘����Ӽ߀�� o0���B�����7�'����1}@��}B'�*����y�N�3��P&�G3����阕�H����p��6ׇ����w�3�i�A�K利��*)9�"y�	n���6��(3�Ee���N���{*їGnSJ{	��x9}��*&�U�FO�dZ���5&t�"��Sx��d���ˮ�sE�B�;���c��խ�\W(�c����ػ��X:��gx��t;�w�O}�����*�픸�Q�)�����Y3���	�x��U�^*,C��0���	��N���6��[W9./��"bl�ٛK>^1���'{Pghc�N��k^E�:�����ü��Do8Qo�����ฆ�F���d�h�f�3ۛ~�1��G�'ї�^<����s#M��D��޹���+��I?k+�$�L"����_��FfMC)�Vf��f�U����go2��k��ь�⮝�QoM�����jj7�*���~��3��w�%�2�o��i�;���]��UP�-B��%4� �P]7��w��/�J=Q��-��>䇼ᐥ �����Y�nӤ-:9x{�Ov�b����^�u���]_	B[��;Ϯ�-a=#�e$����%�ʬ�7�9Vr��Y~/��U<Pg�ÁDt�j���u%Ӷ���f��{+�8����+�:�)�!kh@��I�+������o���m�w��`����7��B�Z��&�
��W¢�殦�P�ޕ�c ��ئ�ط(V��x)��b6W;:Q��򟙬�en@�7��y׭`�~��@��Sf�V<�ؓ	�=�O�nEf��5ł5���WO����o76�ǐ����c��62L�9fR,�1j�h������J|�*Ig��n�<w;C.���6���(z�ţ�!9�X~�,U���d��7���-�U�Y�#�VZ����V�r�^)�?`*}��Pݓ7���F�╉r�zc�n��W��S<�����dn�ϐ�㪓
�U<�>K�Nȣ�Y�0�5�0mV�M��)���n��Z!�Ek^��5i.��Rz�"�_0��U�/�Y��o�9��yg�-���-��Ň��I�ūWs�N.k�|}h�<��G�g|U(q���׭Gs��
�.(�r��7N�?	��R�&�q���>!)���
�	��:*=�z��);�[�	]C������ӊ����6�z�޽��5}"Gq�p�3\q��]0�@}k깦LzT�hL�5�m�������ݎ���	�|�ǈ���ФQbM	Z��?�~��LB�p�m���Ä�5n����J�wUKZ��h:R��-�l��Hc���ѹ����Q��L'6�9Þ��M�].vr̡Dt52m�Өm�:��
�٨`2�x.��ƕ���}_�����y��aOx��*Br�7?�4ֳ�����D��`㐈¾/��97Ƥ�pD��1��/b'SU���b�͗�S�=@�����/9��H�� ��K�0"�Nv9��'nq�0'̂Y��e��b��/2z^�t�^�B��H� ��>Fm�=t���7k�5`72rm5�w���y�����,?G��e���c �!�-/ ]Y�L0�8�]�ϊ���vMM27�#d��P�?4�۪����T��0��Ri�1HMܪD���y:x�T�岷�^�ow���]헝�:SmBu3�x(Mn����)�v%K'�Oۓ]5E��c�F�#xv7���/���8>��z�������d�wl���L��v��H!��Khe9��g*`�"�t�]�ò ��fX��]6�K.��x�����uqA�|hn]�&\��.3�Uu�orYj;rF*�û(Ud�O`��,(R�������8�bL�X|E`�d����s�R5y����>�NS�28'[E0p�/�=�ɜpsJ�>=����t�'YJ�ϕj��#�r�`V�$m��^�fS���[*��;�
�^,�ƋT��x��a�E���n�+{����xZ�Ϫ>Џ�4���'|h�|��S�&��rf� Qy0z�O43cܼ�[��*kw3���ޙ��f�{�M�N��wL���g��D'֩�ms^Ȗ]��[��"IU��i�]��R;]ou4q�������@���l��r����W�V�$��qS#'.��Xܡ�Ŗ�s7h\��Xu"��ڕ]����`����;C�+����`��ɗ�㟢��#gz��`�7�m�P|�Z�F�k�X_P0��iW��w����v4a�sg� G5�|��v�"�C1��k��vP���M:*G{��f��<L������� q�l��k����L�/N�A�����YLl$\����:�X��E�u����i=9�@�[vFv>�t�z	X���\�s|Y�y�5��p�j�TW�ٲ���;�S�Xc�h�,H�%ÿ6R�x2n^^c��Z8�xd���1����~��c�2}͙�0ۼe�
R�i�����dA�Ww��l�dD��o����=KMG*K~�����(�o�U)��ے����)�Vμ:kҨi�+[&�"#;���b����w�H��c�"'�k�)�4O��v������@�YB��:�������G�����㬡P���(>�[�6O��_c�j��*�:I��K�5�(�i�ĭ�0�m�ݬ&Й4 -����,­d쏝�A�v��� �7X���Nm�}��r���]W���坘����v�s��F�8n��ObM֏��7� /���H+m���#�� ɨZ�d�`��mخu����xiᑆkk�7#��jq�N�YQy��f(�v�l�vltJǰ;���|�Si���Kd��� �b�yn�����L�"ؓD�N�f��(�}j�Y��84|��P~R���T��4#s����+'���c6�7 ��Fv���h�nr���o?�u���-�����վ%���v�JKW��\��zO�L�M�-�8yK]��c&��'nGGT�A��w�ȟ��:K���?�o�Gs���ƚ��"j!*��l\&��.Stx��A.��ø48�����o&:�J�5&q�Ll���XW<o]����]�
�H[![�����-��0Yb�s>�����sđ����|D��Ur�������|۽�ݧ��CU��t='��"�*��-�hO^���Q<��;/l��8;k��#�,�5����YV,eDf�g#����^�b���Dv�07l_�b����P�7��~�3�S�hO1ƒ�����B�9xD�02@�q >L\Lg�-}g�P�~whu��e;�,7G��H��Y$w4��$�c?c��l
�����.���q;gM���EK[ �x���H\*Gh��ܘ��2�H�Bh�q���p��x��h�;��4�4w���aˈ�d��|j-Gf��Q���Q6\X��$�!�|�g�<��|�os�o����%�c������d�2�v� ��nv�)�� ͡-�Si��
ʑ^p밊;W��J���Z�7Y2uim+"�G�mh��6��'
����\�h�\�s�߆SS�qv���[�f��)婊��z��;j�e�#�]�0��cqc�Z14)�*[��]L��tSc�04��WԫM����s3C�Gfn3Q�'.L���)�Ve>��w�Å:�mv])VQ��z���1)���k.���q��Ώ>����r�]>� M)�Ӿ��1^�Y��jG6VrS0ƣ���P�7�uq�z��n-}�R�"�&���PCK���nV`ЯM�-<"ƙWt�fK���з~��_Uř][����c��}a����8�!�t��Ę�;�J���MG�:��2��c7������]�һ�c5V��YN�o1�dk�Áh��u�Ya�܎ s�H�JF�������wׅ#PS� 9��7B���k����v����U1��B�[�:�P��\��և+�z}�<p8E纎�#'��ʶ���'ï�l�����P�U�Ky�����!Nr���n�5a&��鵍(.��f��n�'N��i�<�;v=�X����,�K@��4�l���S�l�8��@n��xq���Hډ�62v�~ʧ��K8�B����{�f=ԝ�� '2�^�w]Go�PY�������hX��ս�Z����oZ�zld�6j���Z�M4�ㅺ�&ո�D*��� q��Җ�k�OF�t^`L��UsrI:�4�j��ux��'J�����M��
'���Q���(�a؝zζ��/:V�P}���(L�Z��J�}G2��7����F�5�.�q���yNI7��Ơ�d[\�[ܫ��d��78=�s��U�T����n�8��+w"�O�զܼ�E?�Q�����M�G���{{s�nIW��v����/�w���CvI���Q=]:Y1�gqP��xoy�s�$1o��vC?\��������#/n���>ۨ�HF��}c��T�q��֞Ż�����'ly��+�AN;̓�mraU ��CWA�9賦�WZ\ޱ�&k�+b�Ո˵��
��{z���Pĭ�Mh�Ξ��gZޟ�^�nJ�X �ۉe�QtȨ麾{ͅM@k@�α���n;lPHX�+����2qs�[=�y��<�@���ֻ�#���Z�o����e�Vz:MP�����=�bp:V)���N7EY�e��쎲G�mV4Za���,-'u�`RW8�J=6�;C�9��#�ݤ��1��1Z�_DQ!'�:���+��u���V;,c�3r١�.}�1��b�r�H-�̻���-:���ظ�8�Ǽ�j\�ʽ����iF�]��Zے��{>-���eW�*1D�N5���㓯����q.I�k'Y���v}�''g�_-)j�چb�sP�ȶ�G�+T���esm��J�J1FzJ-�c�Df�OS���*�u<ѥ�u(�R��)���Kj��'�6ъ��YP��++
3-�q�'����&L��5*�"��Y��b��+z��
'��V�m�`��iUԺ�(�͐��\��^�DD����*�Ucm��E�ƔVУ.,�m,g-��( �*��5e�Z��V^R��<��U����,�,g(5����o)��E�m���2�j���hTF惔JT��d����x��Aik�E3��9���rUE��W2e�9g7��E��T���.�����m��c�d5K#8�W�L)U5ݹ�ƥ�8�d�ˮsCk��8 k^��-y��X���8񅵶�Vr�V
�e�T+
�d+S�=r���K|�^�`R�a����e�j�T���r�ղ���]J�+}�8���8�W�eF�sF��9��(z�1˕0��v�����k��h�blE�%�ţ*����;�+�]��gH������'k��Or�����p��]����HOWo6[4[����7���G6�{<��΄|��K}I���0�z�_��k#G�۫����{z?׿��r����\k�w(�zx�}$t	���hn4�;�	��~Y���v{�c�8����F��T;%�g6va;\����&1[ˀ�O��&#���1�ĺ��ƈZ��At&O|���gP�Տ8𕜖cV��{�0�8��;��Tw�{.�yA��At�;��~��4"=qYg+��؇�9X���B]�*��:�WX��w�s�ʄC��3e�Ȝ�:.+[%�//��^��n/��(�?H���ڱ��@�??��&�|y�����m�)�
�b��~���nP��I!A�k�.//7z��j�y�B'ֈ{Ax}��\�L�E�f�[j��`��E��Ic��G����N�D�,i��[�/��yCn8����L��a{�Xx�����'�;𼌽]	�����í�6��&��-���S�f�m�L�LW?6[��cL:eʢ�=�|~�̂��ѻ�v��/����`a� S�U+\��n*��l�D��m p�o��p/K�u���B����k|b{.���=Uмߥ�����-R��d�^�q������q�W
u�� x�w0Q��]3\�ʻ��N0���	au=�/*+�t�d��{��C�b �� Џ�����(�)����tI���}�!{��C6��--�|z��-m�{��O�߼�����j��T�gR��Lm�yO �y^�4a�x��,�F��y;[>�����e��D��cW�a��9*o���q�8�bc,����T{�8ЬU(q�za9�S��s��rz�L`����.���Y������ �i�q��!�6r�}_%�僩A���T���J��FV?kq�X�s�CE,��,�7� �Gr��z�_P��Lhu*����VC�ؕ�;��ޭL��GTj�h�`/��phy��,!�T4E�`�ȫh��k
��j�j1�`gQ���Ls�b�����p�?^@��G��=�)��d���خ�lff�j)��/���E�J��r�ˑЛ҃q�0��!�t���U�v��|����.�c����=Q�SQf���nԳ���,a��T��g$N.��Fu���[.��{:<��!�/(� �
V�Ƅ�槝��n���cU�$�P�!6̋�p��S���鵄k���?��a�R�=���۔�����f~]��A��U��8�V�����*�'Ѫ�cJp�Y�H���R��o�FhYb���W�M�����|H�bvV�i���X!���p��:�IC�,NѰ��jF�]��3��0:s.֫v'����P�ֶ�M��`+y�s�Wѽ��j{_JF�>��t�Tnh��������0ڋ�F$�|�L^�t�;6���ˋ��6g��zh��f�$�����2�j,�US`��«*禋 ��*��s�.�mYSl
z�����_aFw��ɣr�bI����<�8D��r��QƑ{�Jr���۽�^7^t�s`L[r�5�Y��a�>��W������(An��G�����a�4���s���G7W����X"�&oJQ���5�����9�]A�<�"�P`���D��ت�ļ��J�N��}Q[���T�����|��*.��_��/��:Ɖ����0�\E��m�˪m�RZ��J囚1�̙�F2�n���D�L-P�-�
`�֘v����wf���Kd`��
�uX��p���Ṓq�r�Oˠ�Y�����ѝ�z�_]֋=�E|5��yQ^����S�˳����j�ֽ��]C���=h&|q���d>ѩ��#{��Q�F$<�S�_ye��ԝ��e����!F�NCc���#�˟E�z�R0(�N���.�Y�SDEu��~�Z�~��p+1m������,=(���×��p����mu�9IcMΥ�s�@��
��f_=2�O�v�MB�B�����Jǟ�?����x�ߕ��V��4�3j���1���e����M�.i��іv)G=��y�ދz��{��%h�,*����8��{/������1�ϵ�����;�m�ZGǋMO6�WL��ƾ�G�߲����,5d�J�P\y�&O}2O�:��n	��F��_�Z��w��]=�e5���h_��Y!�{�]����C��v;i���ac`v��)��7&��(��]����b��rv_��P0�����R=xf�Z$��ݙr�]��/O'1ɮi���D�9���ƬC��{���飯��1i�ɲ��*�o�ek]���xj��D�{g�B;�y����FL�oF�p{B�̻�C`<.��V#�N��b��}O)�vȦ��o(���}E�f0'�t��ǥFWMjv��&I���lkZ kOLq�u�n7���rp.�{�P�O�n���4�U_q�4��[/%s��6v}���Y��� �'�㙯�Y������0Q��ş,6�B��ܛ)o=��΂Ŕ:�]cA�#lf:䧦����LF{L�wO�((��kpZyM�	��|��,�ܤ� ek�t༆�=�#I*�'��&;�ן��sfy���&&����v�����.�bg����V�0�]e���7i^8Q��\ٷ��/����;�P��X1��NWL�v���\�҅�\�=�'7�n;����Wd�h����wǹ� w;����_���L�[y��-*�����drKM��=��͹c�mJ����+w K~�3��\���Q���1����ٷDF��Q���.�V�/s��ڵ��E׋�>;��i�[�{Θ�x�&z<�~>��5���G��;a����1c��&yc��`�'��ܨK<�:�X.g�����8���U��ݥ�1�����������/�@���w+�}%�Hu�wc�{Ui	�Y������1ꍯu�[����kf�����2N:*��jKU�P���lne}�r34=�Q�&�G���L����	�
Uވ�0{�y�_.>�0I�bj��ȉ�:���<��v&���]o�1�M<f�z؍b����qP����v�b�]���wU����yח�"�Hx�F7po�d���/M@�7]~����O���p2�LH�|b}$��Jԍ�*�\�ep�+ua�^oN?|��kj!W@��B��̺�
��`�K�/)���m��w��^S�Ѥ;Zg]:.6�+�\��?L���\ɚ����%5��a1�1E'��#1r�����L�.���.M�D��&��=W�*\6P�z����o����թ4�O\�aQ;yr�ώA|����[Z:>�niyYtz;���h���vN@_=or�&�І�/t�Ɵ�����L��\�ʠ�[s�c�\�x7�~#���'sF_z^!Y���1���m�%���Fdi���-^��7M�ٽ���m�����y�i�VЫ}���~啲��}w��̑0T�=	r�8!���N��P�!��2|�^���T�w�E�'�c��S�~�`OK���Xxg����\�_Vs'�ib��8R������O�|#��Bf�a ��ܟԦG�9��R��Q��cm�9��`��	��F�$�w��hKƷT�LK�G<u�Q"�8чe��FK%���	[l��e7g/C5u��̘����J~ �B`N���.Lq���b�gjvoO'�j;�U�EP�h=L�b���y��� ��t�<�=���\A'弮G�/E�:gYo_��C-��i�xӗ/�<Bmј�˓�k$�)ڡ��/�8��,.��
�������\����Ȭ{����ÝX�����L�י���cƟV���?��b#��'|�控�/����/Ub���J�`a���Kjh{`��,�3��G8Z�����w���IUI�9�gu��wc͞�O(���+z8�-e鐏+ћ���98R����Џ����휳�;�w���z/�\��Sms�7���x��l��{G��ir�;םXI��1�<>����ʥ6�L�\��ќ����jr���� ��B�K6��Wp�;�2��+���\��B���g��	��^��\^d)|˲t5�bJ�`��f�ӕ׍�B���lu�0��,��o����H���`D�����>�ڦ��{�=6בi�Mη�0�,�2�Y\NZ�\r��A}ﮙ�eF^��Ev�5��Z� Z�����%T��P��E�+L��]X3��g��}�t+��a��۔���%������W���z-8*r'ŚN��`S���p��3�^6��s9S uK8�Y��ʱ�TC~�G�n�#>6K�<l��ǖ)�0���s)�����d�d��9����ĖL�c��S"���.���� U�:��;�0𓌷��$���f��>��Z��V�W�Uњ!��O��:#�t����B�|3L���舆"�j"]Rؚ#ZL��b��[��k�-!�4���TS�E'���ۙ���Y<]�G�N�2��zL��!@���R"!>�=�ջ4�[{�/B(����ɝ�5�6����iO>�j��f=o��&���!��'�F��z6w ���l�,�;E�a���L�+hiҝ����3��cn���%ࡍwE���7fL�ݔs׾�pT�h�՘�>��X�J]�,֫�m���#n.�˖����E��f���ۨih����-��z(�=z�浝�ۣ��������ZL����]����uyӿ�|����x`��S�|��0OG7�n=�ATG?�0O�^�ϼ�E9|ǡ�r� ^\e��̗�5S[!�i^6JKj���Z�S��֯qk�cF71�Dh�C�`��B�����]ױ 5S����g��<n6vcjٶo�}�cݳ:T��H�ᱰF+�'^����Qj�Y���ƦmM��'���
�^�a������acf��BޠE �i<�i�6�Vi�{�V�}�@"jD]�@\y�&��&=�Z��¢�;6ݩ�C`�7N�l`�9w���uޡ��,c�ű�����-5��'��r��3˙���#�>G�y�m�e��;�\?��b�ω�����<WvҺ�C���=r���	��,b��|�J���߾�����T׹��E�ݩa��5괥������)�wDDŵ䖉'�m�'���?I�p����n�g1��H6���z�o,vu8�peM`a�d�U̲��+M�tĜG��w�gѧd��R^%kv�z�C`�hDN�5�P@�[@��'^ɊN��QI��l�m�T�=������R���Sr��:��{e�,68,s����+��~��eH�8KaW��gp��1�vt���� sts!tfV۩Y����J�xd�F��ʶ�
ѷ�	?�=�q���>�E�z�ɹf���R˅���Ii\�2�-�Z{�����Ռ���~o 	5�����ɵr�����4y��<�BM��Q��#��0�(%G�n��-Y�u�%�9��4��vI&��M�ۜg�)����/������~���:.��<΢<!�C�&7�wH����q��F������g�0�dAg��-�L�0ki���F��1�^4�:q�r�~�H�h3���;,��.�^w�2��"�ɹ8m�ޏ�o~��&$N�r�XܵcSd�|��<�����|�/M/	�:WĄ^l���S=��To"�s#+1�Lv��[�g�����Bް�����A|g41~�]��7i�mWh���<��/&�9�7vO+7�g2 ��>��(�9�b1�
��������k�]U�XTLm7h6D�N��ŵFAydt6q�� ��a{%=.z[�I���z棵~���9���Z����H�m3��hBh��ݲ:�����H����f�5rӝLGEW��v�˝�/^����gB�߹̈́]�'K{p璠g%��Bf;� $����J�?e[N���J�� �m6�v�q�}�u%C�x�3�Ot�}�%wc�ǚu�$����O[������g^�7����u'F�]}����}�M��!��X�Lк�H�ڤ<k�x�Aw�X�20��v�C�k�*^��5��/\�}$���r���v��3��׎���3�X7ay�l����ԋUs��H����-�W���E���79�����I��MosMTk�_k[���x�nS滀ʺ]�KTy9Sq��꯴��\;�x��Jhv�X�9�g�rw����*�T���m����[��"��$��	{��t�0F�����d�0)%�f�U�^�y��43,����_��ӢS��Ћ�jd��~�׮D;3d�����e�"��fh�U���O�=α���'�TFog8wJ��^�SEE�ٸ��Zv��J�4��n�RQ{�^X�!s��-� �u��ޥ�}�t�<hn�Z���<�r�P+�<V9%��8Ȗ��N&���2Co]�!w��� ~�|l��K|�woz��>������Ҽu$��J�ѻvF��}c���f����FӸ��d_+���|�V)݆�p|79�fe┨���t��&�N�����-vJ��/a<HO(��,�H�'1�M��R�z�H�9+a�BMo��۫��������n]M��.u�۵�&��*M�����m]��}C�P�n��ܗ[)�92�y����jݩ\��rΈ��%���3v��-��G��OC��}N��Dإ���]-�/nn.	�9��7V�r�KG`OM�왭n*(��ra���<=+.�G����x�08�Y���v�qX������2B���T�zR\4YjEn�B�v��6v�IO;��i�_vd�֞���&�p�Ŏ3[��D!��M�*��|f\:ZO^F�.�r*������G`����g_m7��]�Fr��x�a3w
��P]��"�v������l�F��B?����7�U�8i;���k�+tE��������p�_]��C��i�X&��O�)�2��$鵯f9DrI�+Q��`W7q�����⬨�'l�Ӵ$:,�f�1�G@���6�],
V$7p���>��b��b#Umִ��p��&��ES�� vy��v�fs�����ti����ֹ>啗�Rc=<�}j��,P��E>�g5�x�ua�ͦ.}w �_is�����v�5��Ԝݕi+�/�Զp���R]o-B9�r;�F,�����=J쎜���:�V_�
�w랋@`�R�����I�[���X�{�C�-4��d�X7jS�o��of1I�Q㋦o]��|�A��[RbJT���,��t��
p�؃����	G�-�^���)xX�uA��rk|��D�'e�yٻt�`�)�k;����n;%rI�ʍ��q��.��[8��ҫ$����5�D�$"��u�(9������k�Y���CK1��m'�mb#(�s��	Ǝ
bd�5j�wzp�-� 0�Jo.�xZ2�T6*���ּ�Rq�J�J�=H��qz��2b�o%��MWS(
��ȅ����Ɗ��ھ��/�%0�4r�:Jj5N|�ԋ��N�]]�mE��.��԰��#��U´]('u�9�n�e�CE�(�m��$���m��tdy��F�k9��M�w�{>����^h��.9�*��8f3S��c�D�'Cn�.�:�� Q�d�U�;��RR�ut�9��ʼ��ɝ��T3�����,V�d�Bi`�[�2��m♕��ͩGy%o&�|J5���b,���Tq%"�u�Jw�%A�sl������ip����vJ�k+��'�����49�V5̖�!����Գ\8�7uyW�u�oJT-+0��G+5���Қjċ+޺�n�nD�����\RD�:�ѻs�h�����h��#Fѵ�j�6c�.�Z�[p`ʦٲ�/F�Ĥ����Xd!�r�0�GW&���IJ�M�I�n�d�H��~'�yK��jc��c)ͥ�q�vJ���X��T�YW�ɋSkl���/��'��N��#X^�K<�mm�R��!KK�Q���2lTJy����r[i�\׉Z�DN5�<a{�ɧ������@�P�b�#Q`�2�B[l�*9���*
�-;��yN �Lъ δE�@QD�<��Pu��J�%4���X�PQ�v��lRf*Vq�YY[�}Zq-��+��m��eKj���f+E�b�Ƶڹ��+��-��2����DL���UQ#iYKy���,+*1'-�<)E�k7o9e�+yr�z�"�,��mRV[h��s��/�KB�x�TAFҟV��C��5��)y�kl.�j�S\�~7�����d��Ԭ���Q��5Z댊1YnvM�1�e�B�K�_/,�Ki�<��J$Q�(��Di[+XZ�QTGP�,x��-VQb��S5���-����u��q9�>�����}75e@n��Y���wGM�U������	ID��J邱�{�tN0��DQ�K�*w�����/0�� �v��T�:�*�����>ޏ>��[��ЙZ��Қw[�d�@ѭFa�a���N���֩�t��+s@���ţ͉L��"�i���	K/bu��Q'gͽ����4�=�aͷPn���Ϝk��vr%m$jE>̵^֗��쮟�Z�y�T
y�_Z���@*�2_Ca�[wa���Gv�U��5;��^#��D��u�=x� �)�2ዚE�ם����i�cJ�=��'%�H�l�eLbOj��3)�٤ĔB|����r��&�v�i�x��#�ݠnө-��(1T�fǣ���j�߹Fc�N&����8;U�	�XE�/���nq�V�ح�=f|�pܪ|���H����j0L4�Z'8u���+����J�I�9o�O�4�V��s�x=Ϥ���$���h��xh;�����lr��F���亳�����W���꥚����Ʌ��I���c�ofּdTO�X����Ԋ�x���JhU�f�u�u4��'�̓�A��-��ta��;�}�+�mny}�+�M'bdw��s_VG�+!�P��18cܨ�(ң�W-͡Rf� ƀ�ێ�c�H��>�glp�����lݝ�T��f��>\�Ǚ����KISz����w뷋��z&�f	��/P@�u!��>&َo�_h\Q�и��|}[n��V�l���������b�M��a�ނߟZ�/|K�N�\��uU(����n���rO\�ܠ
��:����ʠ���>�[�&7R��P����<0�xn�Y�� ăkaQ]���if�rm�p�t8�X�S�\�y��u5E%3���x�� �=�M9�w�K���cq�X=����r����wl1j�����՝�ذ��ny�A��4��NZȕ2�����E�=r@x�X�U�Q
̋c�l���QM����[q�/*�7�6��n8�4+Ψl4��v��!Y�
��1��nӍ���V�vu��Փ���� r�t���v�dy��!%"&�P����ιO���Mwu�s���5�\�|��|7���W���>�y�/�fB������<��mM�`���p����r�M8y�L7ċn-�Mf:d ���o=��B�)3��m�Z���;q�����dHs��`�$#ܘ1WM�/���Bf�����:>�1�Xv�{��9k�zy��86��7�� �F׺���۔��kL�(�֨XbH�������ռq�[n���E���
��S+T��t���[ke=ؗ�O,UG6���d�K,V�M�*�l,��
�R���ʩ��}�����o�y���%]��^��VǛj��Z�2�"֙�|�9{	e2I�95s;�P·n���7�؆�ؑ�ʇW��\�)�E�zզ��4�9G��:"+)^�!�4UuY��7�땲	�[ՠ,�|k=_���j�Ѯp�ػV�u����y��H��^V킻g���z(4��a��}i��1b��W7�=I"����P[�1I���~��U\l�G9�w�0,-��6�0MndΪ�W]ݡ�MI�E��ʓ6U�����r�P+��'�}��N�tZ�^�(�w'�c?2�nW.�s���0R�Djg���7��ayԊ[�t9Oy�eZ�!NU���",_e4���t�E�q�^��z����GE=�oո=U����;��?�^�KS�vf�(���Q�܍o�#}�&��UE��7�i	u��3Cx�u�
h9L/Ე��k�����ӵ���ᴫ�^�R�Nǝc$ɍ����8o���v���P���A�2 ��*��X֮�:���j���q�3������{6n�^��o�.�ts06#"�g���B�(���Csrn�r��T�>��?�x���4!�Z�1��;���*��ܞ�|��u/�9�3Hj��:T{{q���Ŵ_*2ܭ�t6��D����hj��Cj,77]ݍ�&R9��[�e���Q�y��O�a[=x�(��gB�Q&�¸�خ�ށ)����"mU��,&��I<2A�9Au�(p�F����C�Ibsxe�`���-y>�i�%���KD���-���JNp��>�8gi=�V�T|;�Uov3�٣�5���jE`�����u�\7d@9�{Y�_)it��V��*ɳr�\��ʄ��0��=A�\��%�E�1��ݲu���k�`�_����\�`�y.1�Nt��&�� \�%v��e�W?.U=�B�M�;�^��&���,=�S3�� �3"3U�v���1�7P^�)�O�a�v�B���KSxl(�|r����OR2����rF���l
��+/��6�nl��Q�yy�.�6:(��������O�M`�@{Z>��ͨ�x1�U�^{v����޹���l�X�m��//Z���}�d:��� z�X�.ѷ�W��PP����mut���%��������vMӲ�`v\f�c�<��=t�X(��=A��]���C��Ve\�gj.�	e ��`�7o;o;�zOG�8�]��O��N3)w7�wQv���҉�}t.�O>8��+z�kc"����K&m��{�+v&�E��|�P\����I �}̤��Z��T��#��[�xq�8���@f���B�>u�e�
�p�Pk+��/݊���i�[$̙n�ݥ��j�j�ؚ��
$�l���b�$<0c��_@�[ s�[��p��Ǭ+<ƃ)ʲe;���n��2��Q�NC����k	��Y�:��䁐ȃ �P��lg��+~d�u�ᗹ��?~]����O�b0��5~����y�f�A���h�3��_|�å���.��h�s�g-PQ�;n@^d\/gu];��"�qS�T���}�a��N���ĕ���eujV���>�d}�g��~�6/�O)&��u��/L�v�3Y�wm%�|U�J�v��ԗ��Y�1����[��� WD�у)�H�SE�m�F�?�C��<`��\��v6��'r�4�Q�����[�����^ԶR���m3�VM��O*2W~L�b~,��[���z���u�w����b'Q�A��(�Rv�ZԪ�1[�z���k�t��i�_Su�ݜ�݋��q]b����"�)<yҲ����@�T
���<Sˋf��T�*ᕺ��8ۤ�4�b=^�Wi�.���R�x�"�*�r�hg�Zz��� ����k���g��l��}�� ��Zr��6���Жʃm}�������*�G��n��`e��{�pc�i�~^�~~t��!��Y:�B �nh��g�������p���Ğj��{k���*�oOy9d�f�1V�QKǼ��v�^��NA�n��6�0�$�7C��m�}��F"�Tʁ�{�|�ex�"�j���S|�%�ôl[�����L+_CѰ����Mt�S��EL�@��jL�W�Y�z���\�%\��<D�E��gJ(���qS�~��S�c�ץ\-���{/P+����NK$�`O�uI�C}�� ����/��hq����}|�/@���8����n���YOHi3����?�ϫ�����͔��} @��Y;�^Gu�'��l��f5����:�T��`���RY���Ổ��س����Q>O���<+��+v��f������;$>����e���g�1��*�0;1�����+�(�Z4���"r{��Q�`8���5��:��إ�#�|��EH
k0���[L�iy�n��j0ܾΑ��^sy���<��˭�*u=��d��7<�L�x��T�\a��&vr7@fN*�2k�P(I
�Su��N+w�����O���l�,ׅ��k��R�We�Jrh����jQg�+ʻ�F�(��滃]]�y���ͦ;-V��l�-pq)������?�^�;�w
�	d9=�P$�k6�z���W�^��x��i����d_�KrD��E5F�UN��%�5��1}�gM�����i5q�w.�g�
��� ��is�.J�͊���ۋ�Ε�o�@�Q��[���E��C7�T��M�9.�)��pvw��ׯ��nC-�;��R�f��z�[���f�{�����j�7��	��ޣm���D74d��N�
Âzt��)�w��D�Jb����n��6�ou�C��Z�9�����̻	�~E�o�l�VLuT�fY�-��&�H�y2'��糡�����3��h|�{�qW./� $ohGhm��Ci�Z��7vn-u���{�Ln�S�����
�U��`�,jl�j���Z9�eoE!F��D�45��D"f#�ɨ	����v=ȬY��Էn�ٛ�v�c��y��[l�2����!���"a�d�~�_�dv��9o�h�c������7H�= �g��P��h�b.��R�j���㢩�S�F��K�rOXk����4e��3��g�1�d�#o��N��CIw��l�PTvu9��{����r�W�K���nka���r����Y��A���ۜ�
tԈ�]C(7v���t����X�U3.�W�/7/D��֞-6�9y�a�h�pD�]n-=�ys�H��� �|g�&mL�uc\l5�C�Z�-��
z�{K�pg�\�3�2�x��Ӌ�ד��iu3ǩe9���w�9R��V��,� X�'�'U�"�����.l�}�n�DA|�]8����b��wE��E����A�fq*�=o��?�W]���xm���&��e�'���di�-f����'2��˖H�
YN����Cz4��h�iޓ�}�68�����5݀ƺC�
Ed��5jS5��.%� I�h5ϕ}$v$z�)\��ҫ��u"�HwM�L���o~�����J�k���4�M�+��v��6��U��*z�۱�w9���k~�>�h#�۷�2О�Y���/g~�2�W�}����£yFM�mk>
P��Efn���q�=�tWTp�W�&y-��ld�����C NLr/5�ᑵДv;G�)��>�;1ˍ�OH��^n<�:V&�:ls��M�;w��Dk�R}*Fm�0�3�0-��w(�����5��I�{��Fv:�y2ї�dqc'1_�57I��`�6���zGL�uQy�3<�`C�͝=3�Fĝ�Uo%ڑy���
Ll���O���5�FwoX��Q$Cc';�c��k��P��n�- �VN?@z�EM�}��hh��)���Uύ���F2�쬍��In�9����u9��ͩ1I��M��Ҟ��x���r�6r���=��᭨;��#� ��]�T���5�Iw����'�MY}6������)���6N[q�y��v��DFC=t=�m�JR��=�ۘ�2 v)�h�n�?n���� qW�t�]oWǳxO	p�GCfI����eg�/i�P�܊�)�DU䞌�����ݱv���ͣ����F@k&@�a�<᪫�̗��N,H��g��y��q�x���g�
��4ө�Ka�����}f��#�j�48��"	ƶ��q�q�w���Ϩ��	Y[`uD��M�ʌ�;�o5����׫J����b�i���Nv���.qz�������w����L�ɉ��u�1l��Tv��FЅ�$Y���&R�ҩ�7��=�瓚�2��Rk	���SOQݬj|��:���]���F����r�ݵe�����N�=���&�$�W#��E�{�9M�#�پQ�����:q��y�0���h���v�5��`�!IW9�i���Y7�}%�ީI�QҨ���)N#K�'G����Ğp�T�q�C�iǋ2Vs��93Q�*�T@w�aiGF��r��%�,�FENC��R�V\���Q�&H.�V������@&@�Q���Ek���������ܸƊ��I�J]4�=�ȲSJ��0r�)����%�anH��-�j~6�Z�#�Y��uY�Z�zV�ƶ̏�q�qn=�c^]���ѻ@��2��6�*ǽ���RM�{����Mc���X�ihڅƍ�{���#����5�q] N[M���)ޮ���Xf��{ �Pm�lTǎ�}��ާR��M*5!Z�S�!�[�WE%���f�B9����KD�d�V���}q�F��S�<����KY����y�J�k���;u��۫us�ͲޝI%)�V<�����]Z��`���s>��%�B"���u�V6�u5��;^k;�W|��{��ʘ�{��?�Bn��������.��GG:>Ư��6ݭ�c���6_�WZް�^�˙}���^�W!ѳ��k��wJ���X�xZ�Yd�E���5�}5�4�ԫr�ɣ9[ZӅ��n�$��pt���y
�9��s�tX�mu�������ޭ�[�c��QnE�؎5G�������XSͻ)�5yF�=}�թ�:�6ʻ)��Z��'h�w�U�986hX��6��z(n��uh��kx�p&�z7�3�p���&���ae����mр'�a�φ�p3qު�xGh�=[Q�_�Ykt�H��9mr4��v�5�W�܈,��p�pa��wrΊI�^�����X�����T�s,g���;�_'R���ۭr�l�,��홷��Vd���eY��(k�+�R̝�!o�0q\�\��m�T��u�ۗ�(�S�Z� s��diή�b鮉�3�Y��(��Lc;���i�(U��t�X�d���[W�6��T�7{���˩�L�x;Gf��,�u��Nq�3��EK<3�BҵٱZ;��Xi�*��ќ���L���O4�[��wY�vh���<�3�D�re��盱���ù�2H�]��C[ر��1�`�蹡���a�M�ث���!�D�-P�`�ӗ�M�MR1%:�[��
��촁�
YCgP����}M�ZD���溧!�>b��;ڏsT"��^Z�\R�q�Ʊ�y�qW`!���r�[fN�K`�[e�y|:���8���DYછ�:*��޼� �:�6)Μ��i��fgq`v����j.�=�/�@���uo�I�cN���W�l�ɭ���[V)��ѕ�h�(MgDYR�3�edy��<Z���k)$S�G�-'��uon�
E�n���E�7SQ�t;ݾ�;N&���0B�Sp����?�='��[�u�VE%��J#ĨfVĶ5`�{�'�]K��B���'�94�����a��g���Y��ePX�n�ź�����m(���*$A���QS���U#^j�����<��|t��{˟�"d���8&`�5��-�yqZ����%�!Ʈl�H��mE�9�P֨���"Ԣ�"=�}�UE^P*��k�ӳ�QFJ�.ajs~�x���o6f�Ϧ��Z4��U����M�ʕDN�kTz�Ŗ�^b�T���5_��������Qح-J(q�����������U����Db���\[˱[T�ss#F9���TA�2dԭh��X4E�)���785��U��^����޻u�J�v.k��a]͵����Z�D5��,|�<uۭ-���0���b�W�X�+h�S��i{n�7w���DD�P�^*=�oo9�<��rn�
yn����:,5�mF�S&�[�MZ��խ�.�>j��b>i�[J��Rښ�2��5��ų��ZQ�AI$�E~i I�h_�nLh;ۻ�w�HIy�[��җ7���N_fvf.L��,�mݵ�oQ�8��\5�O�*ă�h�z'j=�+J4GU�֬={ͭ��^�L>ᓡ�TŞ3�4�H�J��:z�g�>��-��>ܓ�"n�uŸ�����dej��]ׂ\�>�W�uM�m��|�����:֝����_��|m���9���T^��¢��'�m}ɷ�>�N�X�-}g��|����y�~���������9��s^'�ST�����S8jkva�a��y�'	i�dY��2&c��+\��s�=�S��cmY��Q�=�"Lx�H�?H�o�w?��'�i�fa�[��Q�Y�N3;T��vLfd���"7��{�g@@~�k9�����s�+F�[1Nh�54�ע�:z;eȃ��:�Cj�KX��Izu#a�Hx�o��܆u�|���M������������d�<��%nܥՎ��1�O�ԃ�f܉�6R���9#��U���r�E����z���U;���V�*5)�Q����
v�rIO�wד ��a��y"�7���[�;�VQL.���@��s���ofu��|v����gU�׭�fʳRYY�_n�!%4��Ǐ��l��1�7_Z;ٚ:�\�]QN �zW��wv9�?��a�d��_6 ������]7uu�K$
~@��4rs�)��WY��,-~��._�עM3�ߓ��̆Uc+�M,����(���vr�@��.m���5NoU�U���u%��Z�G�V�3q��7_�-\e^SL�6=_j��'�r�[C����6d)�D?�Z��%�,<�*���sA ��.����+������j!�������Ͳ�^q*8�@)�;]*�4N���Ee��)�WRF�A����5��ly��������B�	�C�>xȸ��J�v�n����p�ܯ�5�ogK��r{�%���
f�o4j��n��޼3~�Ej�u�B��9���">\�/��7��v�6ϻ�͂|�7ˤGj5��eD�n��5�g�o$�Uw������r�~*�χ{Q�,��?}���-{9��m��*~r��LEd�F�d�r	y�h.fcw��F&)�y���[G�����[~Żt��m�����vqJ�l���܉�.t�*�Lͫ6����{Qk�9J�E��Ds�WLl�Yϭܠ��[u�Wg=� L��V�N�\���xYU�r^��đ;֩4��Hߪ��]�r��Koi��2�C8a�`�p�ء���]>����dV��ֺ�>�}�5t�S�u����9I�ڭ�(m7���^����ξ�̘=b�ϣJ���CL����-�8�:�n��`���]5Qt���4Mk�<�z^6�ZW]j�����ys��F^�4�N�r/f�um-�d7����Hs����i�(eMmIh�TgF�����/�k�Ù(;����ټ��l����܆��w��-I��O����֫�p�*��Ei��R=@Z��V�5)��j߯v���m,wdSC2IsM���xd��G�����.��qH��]{q69V�մ���&u���F?	��'*˛k�;�,��ɫ�2�5�R�lq[*���*�;q�e�V�i1�U�������P�nЎ�hb8���;IIN�G�J��C�-㓗<�7koV���u�Y�u���>S��r�3IP�����Y��e���݁S$���k�j�;�]�)�4�)rI��0�
��_r��WK��Q���3B�ܵB��5t[E��8�jr�X3��b��E�uգ��Wo�<.�8�k�8v�n{������ge��u�#V�{vL�W|y�6FS�*ӛ9�27�xD�0�U��v*m8ͭ�!���D�ډ���XR1�� �o�����p0�^;�{��9�8��\�zxo0�#�#���E�'�^Z���ۥ莋��V8��	s���~�ۓ�:��g㛆��Yom������
�ܘ���m�G	�n<�b�m��)���ֆ���'p��l�c��sj}Y�����y���y����$��%�o�)�q㽇����
;0;�ퟠ�P5�L�3��R"���v�bz��i7GKnݜSvDez���/k>�w��������C�4!Zx�6.95�x����֯7)ㄝi�<��1��Z���iԁ��Y�e-\��oT���hN'�[.���3��\�)m�r���3�ȩ�3O�|	�6���(�i,���d��=��hޖ�;�I�F��7��5����a�%q�Q�O��)����1Wl��W9�/�F��3�vn�b��س1C0و�c�5r��0]a׊��њ�U����a�&�BlSVl-��p.o�|��i�  Wf�c\���OR��x{ �<`�$��~��C��M�а�����Z����ޥU�B��:���cj5�LH�e�,����RÞ}�$�Y��]Ad�[�m�ll�]w��w�����W��$cG3W�/��#>mK�7A��׋:U�bW7p�K/6�6l���Gu\O�M˽Ô��V���gFW�PL��KA�Oob�꽟��_uW���ewO�W>��"�|�\Y��� ᴉ[S�b��M�(���r˩�%�I\��v��U����vc\>�K,��v����>S9���ff�.�eB�ܲ�?��5�lާ�olc����~�$4��!��C�Vzgcc:���W���4SL3�d����z��f��}���r�
f�hn�_G�d2M����3�I��7j�=|$a���^7oX���Q;�$dʝ�������F}a�v`n-����Ȭ���m:�o*�.��)o�� *�.ʊ�+W\��{��C��F�s���S�EK�\�4毂����/���V��j�sˊ�\��[�e�[HEhs `mL<��V�t�D�w���ʽ�Ƥ������3�q"��¾>���N£A��R:��hu\ޘ�S�l��y3H����QHjGr̍�6@nG��X*U��Så�Px��at�����O�ۜ��ֹȸ�.���̗�n�d���|�B�h�N��(u��9Ŷ�A��.�I��E�T��722�a8���G�ʬ.PVˑ�;�+gk����"��� =\o��h��*Yb��<�@�J��UjV�s����P��z��J��@���8��������� Ơ7CL��6��>t��K:z�;z�N=\}��rw�݊�����V�V�g�_M5Ϡ��\FK�-ǚ�׷�K�c[���+oSa:�B9e�@g�����04'v��#�S^h�od�K�Mf��Ȍ>�fp�=��"���`�ueGR���Ȩu=y<[m��Uz���!�����[��5���H�������H��5r:��e��4c�Gn�.T%6�=�^p 1MQ'��pvt#x��%5��N��1o��F�u@�/�i��a�-$�Vο���n�f�:T�.�����)j:	hj�9��?�mq5�-����;��#2,�R��n�Υ�d��j��r|�ds�}U]tI�n~�o��bT�t�\g�m*��&*�)n�����9Zq�Y�\�}�~je���m͘[�BF��n�݁Ȭ$��L�mĳ���]dOW?%]{����Sl�y�=��C�]1؍d�td�ܐ�������h�le4ٺ�7�����T��ӿcr3Bɭ��I���D�����QS㚜��=t�7��zc!���1���ɑ�62�l��~H�P�ݑtz�te�#��u��z-Ɔ��V��?N���t:#W<Ǚ�O�ۆ��D�b��h`�v^}��P	!��Z���Ўp�[n��OVE[J�͓�ѳN	4�;�ߤl��.*��wT��5���I�	�r��6��y*+�*oZ�� �h���s��T��3�5�YF���R�p�3}�D��Ν��Q9 q����U@-�~�okz�)�"�{���eֺ���3��ذo2�3:������,�|D9���������x�趏w��}�����cZ#��zB-��[�-�^�7Q�\�����1���]((w/e�I�T��R��w�f���?��ˇ������{w�����'�V�[�+��۫�\*�T�ܹ~V՗5%���ɛQ��l�ө��wB�8�M�����yU�3S]5�3�J�p�H���R=��6�t��;Eo��#La��lo�Z�m��� �ّ���|0h��*`3�H��qe�h��$L��ݚ�g���؛�jѹ]�k�vj����6�O���c���2xu���B\�q�r6��9�9���w�o�%����-Sd�fv�oL>�w+�mv�P����'��*^ܴ���^9��v���2���Aa�;ieŘu��#d�ݥ�o�z*j�E숎���ܱg �{�HL���V����n[��w�]{{���h��@����z0m9M�t��R��$�ٖ3t�;���Drm�p�A0�f@��ȱ}��?a�c���e�Ij{�~\��}�{�7�x}�~lV���F
�:��1�cy�13{=�"c��;������	q�F�9 N�`���7C]�ˍ��}"��U���Q'+,r�6�Ń�d��'��SxӺ�h��&��)dՐԢ�E�bF�o3�7��M���Lc��wP؛!��k2���u�bʱ}[��St��H�p�9�����^�������f��
za��w_�16l?\p�ɍ�m�.���p����/x�G��Z�j�v�.�t�)��Cvz�r�!���T�����l�F���V��@�{�����m�o�$*k9Up�`f���iI���u���N�rP��x��,%�c���q������Yڅ���޼�w8;!��U��ദ��F�g��7�IO�Qo�R���M���j�u=�e2��4�b9.��WY�d�l��r�Ft�f��xھor^�X��)�UW#{�"�Lz�)��,�W�z.�&��	�x\h��W�!����f�qݒM��Cut��v�aO,�����8���q�=u9
�/y;�Xc�ʮ�q�PV?P����֠��F�fC�t�u��OLL�dr<�k7�1�g=����}��ś���������:!�CF�5��8��$�ni}yzl���cl�
���D�ٜ����o]����B�x�v�2��;e�ٔ;4'�Xz�S��S�a�goL?�mU�$Ԓ/%C���hLlm���=�:��p� �����O	��C��m���Rl��ͽ :&b5(�����Y��$�{��)�﮺33��uc��ũ�=O�i�h�p
0#lȹZ�w?bΡ�4�S�]�6���?T"��Zӭ����a����[�]���f�"�-��ꦚ���7�i��s�����ґ��U:A��Ci�6`h
�F=U�
�Of�kh�w�y�Fb�Tvdv�m��N׷��G:sƋ�O���}g��&]װT��2Z��͹�@�1犾�K3!��-)�y��N�ʝcLL{v~*�r��[�X�/��M�.�FZίw'
�Ⱎ|� �������8v6��3d��wJջ�K^������e����LĲ�P*�.�3MCs]WeN(b-c���#j.|Iʬ���M�@{�cA�D��.��������ݍ�Qű�m�qI%�{.I�m���w
�E�u�z�'Fݙ��H-w]��\��$qu��$$�Dl�-�3��l�I�oEb�_te,�+f�u�5�Y��se����"�Lw4UH�����p���Ǎu8��C.��ޣ�8�H�7cF��4db��ɲ���|��M]��Q��U���-N���dşM���t��M'�`�`�4���e��YºJسl43'���%̜��K0_0)gub��8�lsM�|.��� c�dT*���Ն�nto�2���� �¯�u�y���P\�g*���:��8N��Ȯź��o`�E���H���yH�bʕ���u�T����wi����5�-0��e���];&鮻�I̛�n���ܨ]5��&�`���p�.����fR�K\wZ]����Kh��LS��yЦ����k��1p�Ұ �UT7-
A���j�r�s'^�z�7��u��NS�[�d�v�Lk�wM��b��j��w+�;�̤s�7�`O��%��o��޼���{}|�&ɼ�:��a�Wo\�=�L}�G��5�d�xY�'MM��
�&���D��Y��0u�ȷMa�.y�Z�tO2��PO��vr�pn��5�6&}��b��*��]b�7��
�p9�LC]+:�ڝ�`Ô�S��e�)-!���2V�|��1<@W{2��;ɨ��$�Vw�uݷ'�a���Ҹ�����x�3E���l�M:Wf�(`Xܿ�35Lo�[R�*�Iׄ��nMrm�؀v��P�w���8��e��#�f�}����p3���de���xwt9�z��/�5�v���ws{����w #s4�y'�{�*���+���Z����W�qP"��`�c��B�[�+�8xj�fp�i�ɥ��a|6e=�"r���:�e���+x	q�S��A�^�t8Z�\WfXvv�����Av�r�����T��6K�U�^uv �Hk����7vʃ/�r��W�t� 6�ٲ�2D�퇻p���neMΏ8���v�"\��Y� �����X��R;9��O7l�=e�Y���ށ���:�F�+�*�ۅ�Ict�nִ���v�}�hѦ{�C]�Ł�Xk%�sAs{`�I�Ӳox5b��M,E�n�vtۅnr��=�F��h����2��mA�1\�X[�ƒ�3[X�oX᝗HjW�н��Ά�
�V�8K�Z��+�zV-��W9�R��!��k�z���G �vv=O 33���M��bV�HY	�.�9-�j�ڒ�ok�w7�K�wB@���ԍ�)�����;�]N�Tv�,�K����mfq��7]����_�X'��xr�&ʵ�&�2����pN�g_'T*wv�K�7Р;Ky�%�])�3�`S`�X��VR�<�[*X�\2B�G���t��L�*��ݍ�f�w_u�?�	?�"IA �	*�U�Q�u�ƣV*5��*��6��v��G���X"�J��'g��z�|��sR��kA�ӏ\�Fŷ�Ǌ����ݵ�L�_.��WYDYYE`�w-��'���y<�!jR�n��ޕ���=�9�{i�S��Cr�Q/2��b�r��9y��Z֫^!�kN��+)ˑ��)3b6�n�M_M\�g���y�.����E���ZUej�UTKN����F*��E�����mB���^[2u�W�͵΍J*N�UX�2�U-*�V��-qM3Z�8����B�AH�B�'5�T_9��)j�k�s8ŏvmAd�-.)򐦫^j��8��(>�������ڕ[~���NZ��)��V։`�lQj
��NI�l���V,�V�[nJ�1E������
�ʬ
׎yʤ�S�A���D�K[D��i�u�V�4T�E+�V��Ȭ]���d�� ��o=�n�jm���*U:p��j!f<{�RX�]�TbF5\�?Rw�pZ�������{j<���ʽw��w}ΆǮ��V��c���ܗm�G�?N%Fpo�e����\�)��̪��j��9���Q�4��S��av$�x��n�׹[�ِٚ�:�k��d���}='�"Y!3'օi��PnH��O+v�X��2:�s�x�z�{� ���?h=,,��J�G�Mk�˝q�(�~۱<�-�bC��'I�qw��X��$1Οs�����N϶R��a1 �%w��{5�[Ϳ�c$���'쨯mEw[]��3Y�Ù���ϓ� _=��G������{�9��[��|u��}�އ������F��-"��'kݔ��7}�;(lI}&sḬ	�f��y�t�Ndw�C�p��( �&��u38���Oi��>1������T2��"5[wecO5]�fy��o�x�p��Ћ*`r�H��wn�7�>&�r���ʹTq���m_E��Mn�@�
�讐�n��{�݇ Vv��uFvb<<vʛWd�%4	i:ً2J��`�ɹ��u�Xz���qJ.�[���©f���1aϭ����!#���pp�k��O��""�d1���y�~ Nu�:c;�?~�!��Zx�f@��U�y�_�n�$��5<���Щ��c��Z-��B�[u6&|��Zʸ��3)oX�{�.�W]9$���r(���.|�ݗKQ��!����GN ��nB1�gK�{a��܌��ur��B� ���r��;j�m������˟��6�5�s��k�ӭ,ƅ{�W;�r+ū�*�Jӕx
���ٷU�����l�V�,i���K�J�дd����:h?d��:�qK�ٽ
���տ�3��8�|��8]�����C�2T�E��x�ojD2;�{9��$���a"�N0ͣX�v�%��6z�(4����Yb8.�i͗h��l�3���Ԣԝ��U�ё�A��	�"���Px�����u����=4:|�#r��"�Ff��%�t�TQ(ۮ���N�?��~�3맟'�j�z<.B��^3�B]����p���=�=�Y�{d�d���Q��)�^.������okXr'k ��u2�t�8�5e��|����e�7s)S��g
��\�(l�o�}-�괪ۚ�Х��z�d�� y�)���a|�"����|+oV5���3���/������x�'㙦p"�O��㺲�+��M�F���p�i�x��[�v>����U��胾�ޜ�Z�"�ԄǷ�'�[��i،1F��!f�vz�=�`�#���H�Z�,[�9�)�؊�k�m��3ۜ��˱��ۂPm�ڷ�4>}�0�/�ql�~�͎w���2Ǜ��ɺ~�t:L��T#���@�_H~�d^!a���\s�5;��$��	��6DE[��6�\���8�i�n���7��5wL"��`N��v����X���b싸x��Ћ�d6�-������B�u6�QZ.�WN:�A����ۊ���7�kn+��5(�+�/$��
����h�N�ا=W\w���鶴Ӊ��@{����Â��m�
��ƖNq�yt��h\NS��h=s�i�x�v�*9^�M�i�}�5��O���#H\�RnN��zS�V*�,��U3�mD99e��:�u�z����u���1��ML.�c�wcf��@i�I���g%M���6�i��!�2�K��fP=ǻCJ��q��y���J+@���mL�3�(��7�y��zl9�$�MwR��VWM�>*�/Y���Ks�
�OEU��A��|l���=<󝅮+��*oU�wME�{������`dk2j}Mb]6� �Sy��4�C�ˍ �N+w$��Ћ���=��c�-/�����)$�D�����Uy������J|�ݕ��~��ʶ�n{�me�踓xZb���b���S�����'��U⻖2�[6\�銓��(��n7��N�U?}x��Q�c7��+�x���l0���Mu���C�`�X�'�,�%���t?dy��"�gʁ��]��u�BM�-����D\��1�}`�d��4�~>�aaw>#�@XS���}ZZ-[>�pɣ�w�tv���4���W4V6:C�pɚ��-��S�_N~�9ǚ�5�5W�[^`�m��s�Z[��,�a�4�w��k�^\�\�:ȼ#	.��;�T\o�\���ϥ����؋�T�ƻD쎤(a��{tJZ7#�qy �'$�+$�ȅ��ӵ�Pk?���G�7�W�Pj���7(�KhH1�:��ܳlk`�%k,�Z]5(].�qÁ�����3=�'�����9������]^�-;ɠ%���+���j�o,�ۍ+=�������5*��^.M����Q�g��)!��K�[P������oY�j��S�n�+��Ty��[_J��r�����Y�,-�:*\�\e9x���x읠R��U���jdE��1��ҹ9�YQ�j֞q�{��i':̝�qV�	=�AV�(f:�7�,�K�4��]kDGMN��Wn2�:�7�=��ט�Yi�'�tZ�Upq������<*�ǈ֮G�����:�h?�xF�]^nH�O+t���]Y5�a�P��}b���z���:�Lo�3��!�i�T.�v��R;�q-I`�O}��3"\�П+n�ܐ�@l��ݕ�s�!Y����p�ߎ�KȎ����31�-x�>�8I6��4�X��ò͟-�.Q5F{�<sǶ�^�:)Wl���y��<h�*o*GKͥ�yL\B�Ř�VGRg���3YH�r������P9�8̘��H�6�U%�QC3GV1�^���ukvq*�c��r�Mfe�["��{"���%��-C�g�g�2�.�ٹ7���ԧdtz��[(\�`����<�m���in�{��֖� w��ρ��⹫������_H�����+��/�<{�e��Xo؋s��S���j����u���)���<z)���d85�)>�] ���{)�oi�2pU���[޼{��j���|Ү^�)P��D ��d@*
���huA�M B�K��2A���i�n��,G]�����[�j���i�B�"&�W�/lfb~⛃�g��"�A������#t΢����En��=��}ɻ��a��{Jbh�X�"���VE���� ���^[Y�9�L���jf\���y�a��y��(�Ӎ9�ْ��i9XP/H�{�M�:��U ��+�TQw���Y�{4c����4�}�u�����R���Yy)U�zͺlM���jU�
��e��ι�j��K'�Ųl��M�3���]�-���YL�m�/��;�ט���Ӝ���i�z�)剘�k��9��S(�X&�s��5�r\��"hf��Ϋ]�˥���f��ӈ����C���z5�lPi:�fNjrT�+�>�L���Շuҝ�\׆5P-�"��]��{-�0vd��pl��Y��_�̋�{F�����U��̇��0�lzȭ�-��2��D�b��Ք\4z־��k��{��OM�5q�,�O�m�����Z���'�b2n ����]�Gi",����!��vls/��oXC���������!�\�����y��_�wb��lw��P7��ꪌ�5�Wmz�tʒ�v�(�M����ܞm�|V� �1��;)����p���*���#��-I�6�O�7�!FEgu�:��繤&5NP�z�3�<�zx/zs7o({@�Sl�M�H���r�m�}�GI�g���p�U�U��7�&?ʲ?~��} �������!�̈
��k��Z��baR��/O
�M�1�l�
�`����u��wXg�&�up�ї۽�h���-+�b{��~d�|�P�
�i��B��x�C?�;��{Rs�֦h��=N�a�W"-y�0�]sH]޿,~znb�����u�n�費�6d�
3S8���7Ӧ��8l\t�F�m`&���;S(ݽ�d=4��g@^e�J�c�����]�nL�۸���x�Z���LwiYq���c(�_M�D<w{�d���`V�ws $]��}�8��c���xwt��|LPI�Z�m;@�N�e��F٦��%�z�*ֲ�{Ӎx�x��	��@�;|����V�j�3�1<M\�o/23�{�%�_�S�Ǵӹ���oi�tJ���U[�K���g櫇	ڸ��D-��ͷx;a����Trl�Z�Xsϱ�"_��P�ӷ��p�+�g%�ov�2z�M��V�y/Q�;؍N���.�%�>�S&mA�_Մ0yX*�u�W�s��]jCU��5)�N���`?6�����`�"�o�w�>�m�ˍ6:��	�:�9A��e붹�M����Fʕ��u�N�e'����\�'�=a��T�W�	���������5WN�.߀�p����DBީ��m�][�T*wZ�h�p�ۍq��:�{��Sam��e���C�׽U�����vv,��OTwf�f��8W;]����d�Qv������,�̣[B�=��u��S��N��fJದ��n~�W(w[o*��u�)]V��R@�j]afX��y]Eܜ�u=P�(�	��r�*�ٚ���F�)���u����}�}��t6Z6�&�����i�oN���;ٰ���o4�(�����Y���[���/8�R�����飭�fvG{�l-�.���ػuVÁ�d�͔,���Ww��Օs�y����}M �����H�l�q��ҭ�E�2",�����=�L$�{��i����,�T�C��,1���'My�b�^u�g�� �����w}֝��a���}�F����^�VpK��ؠf�n��W�Z�Ǎ=��x�jU>��17S�9��G�Q���GR�Y�b�ﶛa������ͥ��I��o�R>�Oʤ���裦�������o-O=�=�}�*�+J��*�V[>�\*��G����B�pb��gwc�*�����r�.�0N�U���O���:��x�͆fG��3F�#"ZȍƊ��ح�2�'Q�>ɨ5K7����LH0�U�&�0uS:J�xR�(L��y�:6�2���C}���Pv���k��W�a�,���������n�G��4}{�Ԡ����:���	�o�t�������������M��ViI�k�[�L�[K�UwO���b�c;c���S���QϷ���&���خ�5�p⸆⊰^N�Vñ�.�$����"�oFA�L���-�i��S�=]�|:����j�QP��L�ٗ�t����?9�r�Awh�����t��o��(5=_���'YI���<�I��w{x?(�$v3;@��e���AG(�2�g#��=�䑙��#3�O�ys)[����@Z��9�����S��W�lֲi�Z��$�>��0��d�x���ya���L)�*��{Wm�:�P�/��iGOL[z���I${��ۖ��#g�'������_ ��A�'�.�tpQ/�@J�u�֌���p4Y��`�׫�C7wZ��y��E�[�t6��뵗�l�/U��wi��Aey+^��%�Ή���tZ�jƄl����l,�(s�����￿���W����r�BI��	'��S��dRB�BHI$'�P�(u�<�:$aD! H�ȁ$)B �� 	 �	 		 c�,HC� FzMȱ�c@�B X�N0!%" b�  �� 0�Iy�� -��I&ؚI$��F0�d�l��$�Ns�ВIi)$�$@ !$�"I$�$�$@ 2H�� ��$�$d�H���D�$�$d ��I$�H���D��I  �,$�$I$�#$�D���$d ��I!$�#$�D��I2I$B$�H���D��I$�H��I"D "I$�H�	���d��#$ 	I ���?�<B�?��� A�I P!�����������������?����������O�����?i����@��O������IBI���BHI���Є@?�'�����8�BI���>�?�9��~��t=��?�C� ��?`~��L��@$�! R! P� �! H!# �$" a@ d$$� I$dd�HȒI#"I$��$�,$�E$�D �H ?\I	!P���)�`Q��������$P$�H�� �	���߾�_`���?�9!��z��BHI0
��}��!��v�g�������~��BHI>���?o�s���I	$$��$���I��~��$��$���&�$$��x�����t�X(P� ���}�u�S���!	$$���?���_��$��~�� �z�ߏ�~g��A�C���?������%���O?d?�����O������	��hy�C����{��=��>|e��:BHI:����e� �!�?w�0��>��>�������
}�$�!$����Ͼ��~�?l?�1AY&SY8���cـ`P��3'� bI�=�QJ�E"	
���T����UE	
�R��HJ�R��H���*@�����D�)�T�T$����TI))֒*JH
D6b��RHQD�
�Q*����Eh�(�"J��m(�U@��5*�
AJ�QG{J*�D��PP�IE��
���J�T��Q$�U	�JJ�T�DB$�QQP)BET"���e��U   ;q�Ղvk���i��Zr�b�eݺ�+l47aΕ`)����q2��ںnݪM�J��u�R�N�q\렣�j�UVU�i��CrT	 �J���	%^   �
 �BCCB�:w
(P�d=
7��(HP�B�
.�7�B�
*��%m4K��U��ڝq3[jU�Fd�AT�݇.wwT��`��mV�U���H�U �`A   3][b�U4��-�JQ�،,�nƴ[3 [:�ֶ&�ݴ��ݷT�]:�k��'n��;e�u\�m����ӫk�(�T��EET�H�!W�  ��5F����²z�WUa[�ݛ��bMm۸
i��C[a��)�wa]�کr�4:V�PH�mQ��*E�Ԫ��[IH�(��T��At�  �Q@����PKP�

�e�TmC
J�Hh� 1�Z��ʚ�CR��U
���)Dm�T�J*T�U"PR�   muR���*��k(��V*��C
���J��H*�Z��(�*�ڠ�
��ʄ�UPZҔ*�R�!�   8QF4�J�E�`�cC2X(Q�5+E[i�i���*����
��Y&  b`  &T� �E*��
��   ����Pj�d�hEF� �`(ʘ
B��J mP�h �KK4
 R��b*��!!(J)U�  �  � 2 ذ    ��( ��  �������� 
Q�  P���QR�$E!�  X�  �5��c
 ��kF�ŀ@m����  �0�T��
 ,L
 �"��JT��d ��a%%* d ��x�i�� )� ��A� hb'� U)�#@�JD2�Sj`�4�F��&gI&��� =�0DX�<��$P-^�"i�4�	ӽ>����{��o{��~x��������������o��6m���1�v�����>ߕ��?���]iZ���4i���=NXr�m7sV9�:V���n��ǣ��^���em��2��l��WI,��t��f�n�����ذ=C1IIQd���XE;�x�
j�����N�l-,� ���ƺ��JݵI�ͥ���i��
�� f������1
���#N�
�!{*�����w2@d��;��7��k	w�����Mٺ#n�T��
ǲ�	{AZQ5�e"H�n<.@υ�j��=��ڭ����
��(�WFE&����f٭2�i�����hm���J�dФ��כ���gD�%��a��xp�����n+�Mi��
�v%��B��Ul�h	L�5l(�-���Ab�J�%I��Ǚ�oi��� �c-�v�ǌͥ���	�fL�x�R]���(�r��a	�5R�\���5<�M��应rcU-9�6*WM�1]:�.!V&f�Uf3d"��QQ7Q�83V�e`��4� Z�j˴V��j�
Ib�,��z�,{�ϲ�(�)�G��f�Uu��b.�+j*�����!�w^c�8�IW�ؼ��V�Q�ctrc��*f_ʷ5��=v"�[sd��I�嫺�B���P��ڲ�/����x2����Tv���"U�%jX���4����u�;�m���Z���A2�K���Ɔ�6�Z�f˳!16��M!���5�-���A���vkr����m'��)��n䘷�6��@�	�t%��4n��I\,0P��.̖l��W�k*��֗�RI&��nE���6p\�mCv��ޒ]�pa����Au��Ѽe� ҹ{o\��1��n]�+uV�n���J��:�'&}���oU��F�i�	+@�[&�5hGY��>Ц	��IĆ���R�R���TtJ����U�M홄n"p\��!�w����р:�R�t��N�j�9Z���nHC�k\3�7E��5V�Lf�훡t�����mA�ծ�e]�W��U*:f�Ygt Q�r��x�h(��(IfH[�'�%-F�Sh���
2�,�[�( �jlaa�����eiɧ�,R�5*3Ԃr��X��ݥzh�Z��Jt��mԇ���ȶ-OU�Ә�b}�,��N��`B��M�4Hࠢ��n�����jLi��͹�j��EF)��%{��ZX�b��]�J� ʶ���t�bs�c���[`:�[��⎦��T3��+
���tT4��$�!��6ΚcM[��7�ItBɊ�9��).
��[Kn����[̣W{�*=�Y���-�
f�TF�%�vvZ��[����� �6�U�5Цd��K"<a�m�%la�Y��;`�Y2	x�7.M`�͊����`��(�6ED������5
��f2�[Z�t)�#5Q�n�D�ehժ���<�ɂ�yp}t�IP� k�I�R�
ƕ�3t�!�lU���E,�,
��e�Z��a���»�p#-�#v�Cb��6��Lf�Z�($�$xwjI�i��h��'㛌�$�� I���mI�[[F�s"yl�ŗ3X������t��2^6�Z�W�F�XA'e�D�:l[5�A���A�l7urդv�z/l�:�s۩!q�^�R�s���6�e��!J*J蝂-�,0���Ȍ�3^��U��K�abm��)����r�1�|V��bܩe�d�b�'/Te���XК��R�ʘ�.�Q-@�7�P莬2�8bX�OkV�$G�p�����S�F,���U��hX��։�[*)������u`�c��@�B���fb͉6��E뫵S*�L��Xv�0c�����#����.�w(ɸ�CoN�F���-���x�Y��
�������H\��:�:ͺz�v��;�� ������ViI�V4�H&�BL�X%�UJ��
�nY[wF���	�"*�a]F��F���Vm�d鹖͋���;Le��d�m�f|s%J͓P���n��9�6�Q`cEK,�]X,]�I�Z��2�ͲMh�O[d������5��f�CU*!T;2e�:%ݨ�U��SI��e����g&��!�,�Vf
U�֔��ܶã ��=�X��'�9�憗���
cԝ�e@q��:-��g�f�da׫F�|Kp���1��80��%�*��q<qSrU���+L�kf]�-i
ۣ�PRB�0-W�i݉Om��j�Ȱ��PV( ��m�kS�%4�j��]ǗZ�]E(�{��㬀���[R��+�#kd��$BwD]��\�)�%d��Ā��~0f
��z�]�Z^��t)�u3��n��X�B�X��&�ݓ���F�5&���.� �$�.<1=۰�}3H�B�!4-�x�edܡHU���=�T��*z ��I9PA��A�$v��f:.)P�g�3^;��84�4KT�DZX�S��Y�բ:��IE�r�ʇ�~AP������tJ�	jS�a%�V��L���fm,ȶ��#{�T(#Q�u�֚��{�`$+z�;��OJV��-�y5���c7p+�֢!q���n+�f+��5(I�6���o[8���nKz��L�Zf�)u��׸֑,(ʹ�w`�:�@��[%�ݙH%T�b���)��A�[b��m凐��Fa�xsD�\���2�
����H�jѻ*�ͺ�)!��մ��|*(�d����áF)܉ K�����<X� �jƺ7xu7m3p�a�Me�F����J-W�d�ScH	�tj%^ �v�������j�C!�/*i�3'����j�0V���4�f���%{6R���"�&C��ۊ�&�Bd��A�����h���/Jv�0�б%�[�{b�f��,�Ėh�A�:S�E�^��Ґ�n��������@J���&;�лb��ݚ��L:�w4��*�S.�2�Ā��+F�4�t�	��Ǒ�p����H�R{��IڎB��Wub`5�G���"��t�#VB�aS��b�^�����v�-Ri�D�1n`h���ΰb��A7T��h�*�[wc)i;�;5M�F)�����j�/s��ͦ��K_1��%d/U�%�G�¥ME
�7`-9z	�(��8i�����`�Hs��/t���Aѐ&퉕�Iyz�)V�Y��n�Sin���&�:I���z�N&6�y�f�ǉK�+FGW�*͡��3@5��ܬ㖚ȣLl�Ѧ��/H��v�(�Nb�k+An��e�h���CjLlEGn�(핡慫�M�B7�<z
_n�ڷW=�n�ZL���#Fe�u˚u���I��Ԃ�R��$��h���u�l��HŗVU�~��%@a���� ʵ��5n��&#�-�Pը)�-ix�"�ڏr�B��p͎��c�VcI����P܉��i�P�#�/Lq��b��;/Fٻ���Q�s��V�-��oBf��9���9�0}����R3sԩA�U���m,Y��V�n"-RhT��$��ſ��D�gmd�&�v�X�6#XE��Ujbow-�"ҕ�3mm]ɉ��Krڽ8F	�{%�;��n�Y�M�lG���̥U2��!�ѳQ�b���f"�#M�z÷�*l����n���n�y.��s\��Hm^)����ˊ��ݰ����흄]&�8o6����[X�8�W�eo�O^���:#�GA�D�!IZf�Hh4[{sqV��y%�*���i�����=t�E2T�Q�v6��4D�v�
4�6I�!�⺕�ь=�����̟CFi���t
ܱ�/YEޚ��Ӣ0�Pc5<#ve]2�V*Lõ�)S�,e0j�'�u�b��M�`Mc�th�k1:qbX�t(l��!kp7M��y�O �3%#��t�Ҋ����7�J�L�����QkL]6씮�]h̐f�{V�݀G 	:C���U�N�Z"���˅A.j:��"
�Ws,��q��ҽ�B,�7�@�Q#�p�VyD,v���k��`D��n,���zi3t�YؚQ�`�6uz�'�n�t��\��	�T$A��v�f���ٍF� 2	�r����!�"�I��d�f�@�^�qn,����kj�!sLB�h�/P�y��8�T���n�XZaw�w���d��ˌh�sX�%�.�#nj���(�E��%���v�C��Y0�{����h45+B�`�H��Ő^�Su����r��R�x���U4��7Unf+J��7�K6
TAq���ʺ�)ԗM�J�']1��U{T-�t�St�7F^]X������"�f��QC�E0�j����@���Q��[$�
��HW�[�,r���Q��s0�RLق�E@�bUx�c�֦/)[F�,[����5�L�����Q$$���m�)���ʌ�m��i�T^j:�i�Mml��2��]`�����e��@�I�ݰ�i�TlV��S*��t�����KQ�55��-n�dR�Gv��U��6�L�Ϧ��-���t��-��qd��$VUf��Pե̪��˨Y�p�U�3F��Y�p�4l�6ؔ��R0Q�l �75�ں�3r��b,R�yGU-��4�AɅԘ�[Z��*��i���LA{[�d5)ָ�­ƿ�*;n1R��3���NR�W4�EI�������3(ZG��M4��n�[5��leۨ�@	�Ad���Zd�h��@^�:ɶ��&���w���ɲ�y�H��uAR|��#��M�:�㕹�Q���a��sV=,�yb��ލ��P�QK�R�ݴ��ZS+�˛�e1jI ו��)�v��*|���w��Km3"�m%.����۫zc�J7WR^2�$��0�z�Ye1���W�1�);֯A�D0�(�j\��-K.�\�/ {$ͤ"�tw9��%�V7h������Z��f�Ię��K8v�)WR��ɵ6��ED��JX#��;2�_>ʛ�6����Z��0i��+V�/2@
F�izCvC����ݺ���X��m&LM���u�!vټ1���pe+��[)���t��o*�u�fR��V��rcW�֫�wBƕ��9 Xk.���N��q�kPl��a��V��i������j�p�9H�gkjkۨo���ӫdh�i��ݚL��{#��S4�}��n܉`օ�Os v� �ն���_9? %ՓZ�[u�+u���딶^*׋c�T��rTR�Sm��^��.Z�]A{Hˣ�ث��n����a h&n���
86VˈSs#Ȧ���IB�-�cqlRb�"�kl-Ol{Zj;"�U���sQ�md$S�1\��J%�V=�B�mՇ�m��n[�5����ZM�G�Y����jU�%"��ˣ��������[ݠ�4���=*'r�1a}����e��20Ƥ�Oħۛ[�IzUK�Z�@�b ��+���&��6{J�[j�#�͚�
᱓$�4������p�n�ũ�^:��.�g9�ufc��Aɢ�Y��x"� �m1��:�b<7��h.�U�Rhuk~T�%���f��
�yV�;;+]u�bz]L��vta�pVڒ��Z�nǑ�1�әk�5�Pͺ�s1R9�!`��©k��),eX�����f���!�ǂ���3�V3�S"{��A,;�)�V�*Sݬ�c�{�3t۠���͇�� D���Г�Q����-6	RLǷ��J P�ٙf�d��6,Hˡ5+'V�N=J�5��bj�3�/���7*�(Ћe�n�yKCr$ӰM4�>�d�-%\J�H7/�%��l�%JF�)Y4�KQ+Z��\�b�QïM��J��C��C����ȑW�mf[u����9)rf:n��Eաt1�ȴ��Xv^d��F��-U�$�VJr�^�:p3�86����Y1�z�Fc7v*��4��ZZiА �U�ڊA���q]��fس7)���^�`���e�y��t��M���h�/qf���@�����ZwA�p�o��b��Rm �̠���[���^x��Gd��tK���7v��
MeM��̻�����l���N
�I�f�;�%��l��b��s%fU�yhP��nOYf��+H,3!D\��-�������u��1��(SVH�z�����փV3m1��wW*+יR�yI'MRܸ6���~G3-^ܒf�X#�[z�s�E���AQ�Ƌ������)��NØ�/3kj�kF�#�����o(T�)�{tX�rA�M5"�sq���م3��z%��e<�*��X�QLzooU�i;75;����>oS!�Q׺�	:LQ���f��m21��Y�ݳv�KmǕ.����Ǫ�ĝ^Q�ؘlP34�,��^S�v�wRּ.�Z۲��ʆ�:36��!�S1�:�ڢ��\EBj�E�V5G��Fc���L̢���\�zLZ<n�)�?jDKYae�mң.��K��Y0eu�;6�����ޜТ757$�#+Ֆ�/U*#���4��Qtm��wmư�U���J�*h2<Ԗ�Ǌ��+�v�
�`��Lv�eXQ%--K�aȤM^+(�w�l�Q����������V��(�8�6丑[6�M0⭽�M� ᣴ� ];ݫ�ɤ�ڛ.^ʖ�[L�o"��G5�ٺU��Ƥ��q��ҏh.[tuL�zURCJ��*A���H#0--p��f��$�_��/�j��_e�y�F��v6��N����Qӷ[q���ё�F2bbc��Or�X���$��� "��\!��Fj:q�
�O%A��n��k8��ۍ�L���SP	!O;9sj�J|��=�Q�RbKT�Nurf}��s6�;ˊs�����Nw��\3�Vv��S'�v	oodn]h��{!!]6�6h�()��o-�F�`��:�u�D�b�늡[k ��e2�9�X�Q�����꼗�]{��$�lt�T����b<=e�U�b{\eK�fs�O-
��عDg^��X4���Վ+�/��.)�g�cG�]���W3��s.�]����7�}۱�\%E��'��2>��ӕ�V(b�Z,VhU���B�-	i�I�x�.�7��O1��ؙmD mf3����QVjb����@��:�
��q���!i��wm���T��X�t3"c(α�uNevٺ�+������p�>U�z����f-�o��Q�@�u�R����рoSF���\{���dڽ���&I��ҙ{/�CH�M��)�lu��^���j���Y�d�&����}L-��f�Z
�Xl{X�E�D�w)�ʵg4��=�\g�Q:%�;i����v�FK�z�\�� !�gL_.D�ε�K�S�m��3݅��Fx�+cݗ�]@ �nUܽ�(;MsW�"+ ��!��*�I�1vE)#&�c�l�l� �]������������O��J�)K�h�;!�����u��Z�;ݜ��珑9�S����.ߤ�KQAnBѮ��7���{����}�	�R�^]h��8��k]e�f����k�8]`NޕMhCi0檺��w֜�]6�jG�d�����^��+�_q���3+,f��gu��]ݵ��p�[vC�mp�aWC�Z�����z�ιCi�<��ծ�Œ���\:�*���˺ޞ{���]h\8-�������ك$�v]i3a��;�1M�7Y�XQ���Ǒ^y|��淏s�͉A%�w	S*B�f<��ڮ��f�@0�v�S}��T��÷��m�X �2����]��bGT�g����5;dMv8O5W�c豙�L�n3�K�;|z�:V��x�Tݮ��qE@u]�
�gV%�iT^�I�*�����2� _vf>�7];VL�,ˠ��ǆ�K��Y��O���_��ZJw�.mv%Pi@��I�"�,bܮ����S"����K9V{=r6�o.�xR+kun�8sy��M;`*�b��N�d|�v��Žd��yX�+Y��#��2M���ѩ�#\U�ivB#Gq�I�������jĔ�\[�:�U���x�ov�.���=6��a.��|��/��b�u>� 0�j�V���o�4�3s���CDt��g{������#��@�rݓ�+��u���l!���j�|�k3��e<6[]������*U�����gl��W����F���Ԃ_D�n���}yF�F�����[g-㕝����O�^��c[i��baM���泤(W*8�nhcQ��nv���K�|�;��!"�-�*ҽ�eK=�'_ZB���v<-u�ے�6�Ge;�ذ�%��w���� �u�i<��.���F5�H˺�4�>�FЕmk;����Vt�Te�(N��'+��ƣ��|/�'X�Ŕ0�OVa��Z�; ��AN`���R^�0vu�B���X�r��K�q�Js�fwfe�3��K�5���о��`���ք�+���ޙ��#��.������F���������j^
͆��D��:"t�������;�/c�\����Җ/�:����M�Ev�1����b)�e��7l��HM��;��$*��x�t٢�2PY4�/:Vw,�[8����M�6f�[��p���wIt�:�Y�o7�5t!ޡu�%�W;�_k1��-���+;���$�Y�1�v5�ȨZ�d� �&���q�9u[u�FV�Y�d���T+�7P���ލ�XV��U��]����Wʆɥ��Q�77�z���Đ�y���Ӑ��C�j,�PkA[� f���u�ѽ8�����9����'e_
��i��qHB	�����S�K��a��e2��mBn��n7rX��;�M��ݝ�	{GM˹+_A��6��f�.�^p��{\-ɼ+gX�4i�?s)c�B�J���W�9�|��%=���2g�4)�'v���^�Y������zYj��2�-���Q�����ȸ�������f��#�mEX��"B���zgk�è�9}C��i��h�3y{���!6l��#�`u!�[�ܸ^[}�����΁�P܀ݍUs�Tޤi��e���M�9}�L���6�^�w��>`���o:U��l��F�V(&\q'C��톁��\ 룉t΅���0)V3��X
�b������6pÚ�9�Xc}_#�˗���bR�3��x8E�moYbV����Z�+���G&�l�U��U87��w�Wq���Y�#��9
&����]�3���k� h��+�k��[;�S�:��3��CBՠ\/x�!���� �7�����y���w˱\�q��v���8�%v�$�ßm
�H���U��8y�g)<��:M�Ʉ,̣w�w���[l{J�&��3J �*X��D�����t��n�Q``�ͭ�\��bX�d��Gt��WwÝ>z�_�w���]l0�,"qEE9ب*V�7�e�-�m��[��-�":u�>1Pk"����E�2E�N�����p�}�32�Pn����Х�;	@�"w���+�i�ouL��,ܜB�=��U������l��V�={�w3�����2D;�YW۷�Q�iL�-a��!�xVo7B%b�ݡ��oQSv��AR�]*)>їg���C�-�_*#�/(d�ԭ>�V�ٮR����*�uȎ_<3���
WJkZ[w{yLVS}��.b��
��m�z7K��I���+�a�U�G�T "��-l�z��]B������D'7H(^��xr�2t�ͬ��m��pL9��r���u>62�!��m�Kl�oe�0c�F_' 渫�����[��g^���8"ޕ�k]���ęm����v�Z�*�%,7j�*�J��c(�z)��xt��F[փZ�I�Yܿ��5V";������_�����u�Nw�j���af1AN��*92��w|^Z��Rl��V\9
ĩ$��9˭�z�#��.��a#6���v��j�(q�4@��8c�P�m�xݼlP��\�]�QUԻ%K���p���"~�:R�MZ�Z7)6�Cvr����Ҩ(S;���Vh�M�6}����y�wMVYWF��(�C�وٝ}Ti����<��A��<��D�ώ>wP�Ck��hf�D*��$�������2>�YX:�;�]FgjT�BL�EV�.��r�� G*m�����L=�u�e�C��A�1�J��u�u!��^A��:�C�.�&�|�������U�p�u'�>#�����<J��O�u���,�f�YurŌz�����UoRPoe|5, 1����O#�1U����+�s=��sK3�ʱ�p�1x���W��b�Tpm>�1�:���Z���ݚ%�	������X��\�\�]�묤�]j&��������[��i2�Xۈ�"'{&F��a73�F󠂖ܖ�ACk�^�6�xڑ ��g�It:t�Ԟh�����Q)��/��� ����c��n�0dJN�#�Z��'6���7i��8�T�R�y�T���sh*��[���<�3���(&�d�w<��6�Y��	���F�=ד�CK^@
��^U��QY����������hK��B.�l��܈���gK���K)V�lX��T����M�OTâu0��6�U̝���+��I��Ƽ�d�.*��!��3
64���D�[������'�f�ٙ�޹L^���y*Gfϩ��НA`Ч]�1��t%*�nv��lJ�̑����)`�1�t��vC��vtv�vJ��np��]�s{q;�2�]��{Ħ�7�m��tj�0��_.u ���܂��vNs����|�v>y����&tf-�&�|�S��xZ�5�&��v';OU`J��V��k����1R��mXYþzqݛר^)�+���O�z�Ցot=�/�޽{rG�+a�WB��U�1�s��ٺ.�яE�4��Y��K��^9sk�9�dš#z%!M���g@Ģ��W�;cQ��X;8kuP����y�ok��kr��Eз�;fs����g+s��#C�����}G��X��d*�k��뭣}-��R�������d�֛.����+��S�E\۫.İN�Q��Q\w���	����r�t�$SR�߷4��{h��ٮ��=i���Q>VJ���P���L��9==���d�\���n�&@��L[��]�_^[������[�;-��bX�t�w��Ⱥ]��������1�T+d��FI���M��[t�5�)����2z��x.�s�I�s�c�t�1}���Y�Ρ�K�{B�*���wB�b�Նm�6ʚ�Z�W;������/�YC �yr���b���ͭ�5xl��CU���8J���mj�U ����KOft���u_ma�A'�}wf�wn��98�1��2\�j��3'G�X���*+�G��v*��
[��%��ö�;�ƏQ���n�����{x�@\�K�T��
WH6s�՜�٦�:�]��^��=ug [c6_XxƏ�y�� 1�eԂb�-lT`�l�5���xo3;������H�+J����(R�Q�%�@�HX٭"U��Cxu��k{�W��d^_ϫiH���'[�Y�t�g��͉�4��m��x=�8� Y��r�T�![ ����m��%��1XX�o]�wNڔ�ZcsX��W�Cψ�x��&�Y�S������U�v�ɔƆ�\�Nݝ�6�WG�;��]ϒ��`��&_k 3��Pa�\��,2����v�Y�ٚK��u�Ҧ�3��-#\�t�v��:�|`
n�]��;^�$���`[�Z�o���F�8�L ������j9�ARP�و;Of���5凝���f��x6��+��\:�+�%�X.,;l��+��\A��Ǯ��.X+���R�n�OD�+͑��d�\T炮�t}4���hh�]uq$�7�W�u��[ie��#p.��x���/K���esrp@}��-AWk
�]!�A,���ˡ�����>� +�Q�O
��C@�W��z*&)먨�mQ6Ģ6�[��;k<��N �����2�n�Ҙ���b2�;Ev���.�{��Mgi茞�gp^�����M��U�*R5�����;zuF�'�ɠ39^�m-��^�$Xŵ�N>���p/ɋ���&)��` �
Y,N���e4��}S�X�*�D���j8���e��;�W����j%FW	��t����tozR��U�=Ohe��5�j<������J�]��Y7i2r������"
�)A�������F�	Ks�E#�8i�P��I��L\6�۶���ꔀ<��7��/�yC[�Z��m�ɠ��ܷs�j����ԟ�x+Z����M\�@�5j�i\Q@�7~��T�w8
�Yq�0q�t�ӏ����h���<tNf�=po�`kMK�ʞ�M���n;��YJɠ���XQ_i�-�O(��]�o��쌄����*�!����^�Ԥ蕡'�B	)�2��HPz/`�*�h9RU���c]GB��V[�u��	U�N��o��u�C�ۼ�w� �'��Y�א8�K�`q[�n�{d'$F��e�"i���qDm�)q8YJZ�c�s"YϨB���:&{�����e>��AR���9�hqf��ȝ�Zג���p�����꼩�A����YX���x�;]��8U�҆i�(>�$�6��}k�/�z��"Lv ���9nZAؙ[��i1���S���{��������R���|��bZ6�poe4g&�U��$2�3�������8\�hw&M�VLY]S&�;�l��J3j�'R���T��58*5��w',���S+9�k��m^M��x�����p�O���oL��=��Be�3�Fos��C�FU�m��{ʀeL
��vȲ����U=)��Z��gK�N�^ml���ӊ]�ӗ��r�5�f*[�7*3����5�O��WX���]j��[��X���$��Z-�{�6��9ǈ��n���$]�[�Y(ƈk���R�:-��2#��˖�C��"�WgT{-��&,q������7�d	ӏ�k�J�������a�����OG����+Ddq��W�Ly�>�(��1q�-'x��;3(p�u�+7�����V�J`�]l�xD���f����T�5��嶏FƁ�R�rY��4K9�.�L4�^����m��:��,=,�Wl)�=C�΄�^�EE������1��i��t1�+�f�H$���;�X��|��&����1B�<U�B:���a�*k��Bӻ13ۧ�![�cL7�:�t��k�jX�/Q9��8�&�\�p�8rgk$vR��+mM"�]Y˖E��6�.�Cq��N�GմBy��,g���р<��d{�*KFMQ!�;�]
�Xoz��j뙌>�hwÈRvcяU:��+���fv	!��ۃ��DAԶ.���:1��K0r(ތ{aM��G)�͡Y��@�i������j'�r[��}W1���u<=\��j�]��{��VZ/�|;�9�k�bl6iwھ.�͐�����+}ټ�ϬA�{R��V�Y��=8T#5KHE���p9\C5��	�v���[����S*�\�d��Oع�o-�|/�*��A�Q�5rIps������w�����m�����1��w�߿_珏��~|�>�������Z��*r�\Wi�}���;�[I�Q�46w��a�τ��b��P�(��R��S ]���e��G�.�|xv[��
��$��m�+u|��[R���-x�S�jtR��l �t�]M9��e�V�A��,t���E���os�_E�X�%�t��Ưv�h����B�-ȶ]����j����Mcxݦ,��p�m��4��DngoVoR$t��fJ�"�//�
�'�e^+)|{��T>�S�5,�z��v�+N�Y��C��}�B2�������t��9���Γw�
bɻ�K�Ʋ<�K��%7�gZ�t�xP1��.��M&b9�`�d�k�iB�rP`:f��z��a�O啔�z���@�ɭf�f�̝����I�%���ޛ�e�+��v&�Fяhw�|7n��/f>�V����©��3dZ��I3{e����cc^4�Z��U���1���.Z�y[5nT�>ܧ�*�(˲i.y���M��9�� ��"q��q��5(8A�Kp�C5� �Z]��Z	!W�!��m(���c7�V6�u�N��7B��v���h��o.���o9�5��sHf�u�y��XSqEU�J�@Q�wsJ��a���:�ql{��g3)�-���;�XY���1KWX�:wXE��n���c�F��:����y����mjh�����]��&�\��w݁)w@�����TK��k��	o0���F�@7fCUҥ㴢���0��2�X������WvC�^O<�r���Sq��]SMV;f���(g6~���Ǳp�bŝYP^�_F��%���³z� )ܹ���ɵ%�Ѳ�91V��+'Gǝ�̖*��Ⱦ�1���D��e��떧v�����t��p(+�����r�{��`����G�+�X��6�M�F[�B�Bu�ǎ�-�S4T��q��ܔot	�'GXw���یӼ��J(6��e���4u�@�Ea'y3E��U���e	�w/E�����
T}1tT���vj��T����B'�D�ޏ� ����uꡧ�� 9/Tؘ�1v�{e/f#|cֱm*���x���vc�.I���A˗��}%�N:e�ˤ0w$f�E�!�!��qἼ/%�N=5(��jiF��wd9�`�8Kbq炛�:��(����rƇy�u o��A�������Y��۬lW�S;�2�֐^��r*�8񰺏)Y�6q;��F-�Ɛ�@�㍼@8�u�����\�T�Y�E��W�/�q\�z����D�_6vL寞
9wU53��m���jx�yt�	���f��7�\��ʤ�C6���J=;�1Y�&9[��6�7Vu,���in�MۥJZ�\h�����k����̖0]e� @��:@pv�:�4ؙ �Ý�}��b�XS���T\�>��>x����[���9��.�4��
���ywئ� }Xx%�
|z����xOc�J;���b��nY�fs�}�#��rWXw]�Zs�ZP+>W5A����,>��S)t5�#!�{qԭWX�J�ުT�ӑ���j9j�b���d���b=��r�YF޾:�����f%p��(8;�ٙ԰���w�b��+t�� f�1�T�'J���mq�E�)��U�Qm�����,�I`Mo��ڧ}:����q9ƞD��I�(�7C�g*��ej��r�y�:9Y��g��V6�7�r�w$��p\�+�y��ZA�9�5�އ���y)�R^J���s$řhP��gK�%13#��	��իC��/��]j����[]t,=B����p$k�a��ؼܥ@�dJB;z�dj�*��S\����}W�qc;&�yI`ǽ��欇�n`�#��A'Os�u��9Rr$L=�3�-7f���I�n�CNEI�)�^I��0�l���P`SztՠZ�K/�3���m�<o-u'�@i��
]7��xk�h^�JQQ�[�P�fn�6��m����4���U!ǫ+:]g�G��[i7�>/s��XWNPX�wv�7���(���E�N^���rs4NE@�W��(�݌�f�6�t��݋^�o���E�\���I�b�q���YwRVa���ޥ�v�s��Nq5jP������/eGm�f��beAyW�{f��.��N��u�[��%ݍ�s���B��9����)s{0_^��o��	�kE��ky�	�7Gک�&��Rsі6Y�:��u��(enV�X#(H�J�H6�T�u�f��43.sE��5�U�8����2�����$��W�S]���ö�=�q�(n�6t�\�N��v��H��o�&�[�����K�[�A<����6�6	�p�w�<�[[�B����u7ҍmM��*�d�WY�ˬ�!-��v�7����[��t��x�W�Q�"ɚ����<Aק��.f7��+�N����x��*nK�RDa�J��h��W��s9�PZú!`]4'�{KX�$GY���΅ʇ=G�$)�c��Cuk�ܺWj��$�OT����_��O�ڶ��VP�&h]���=�	�P4�[%7V���46n�T�n"��:�����-zj��	l��z7�)qa��pB��r���@�wL�9��&��#E�!{O�u��u�q"�>�y�-5կ�K#�aIT���Sf��qf��#CἯ�U��J��>�d�����V�2�n��N$H���4Nv.���oedR��!B\����[��:ѹ�2=ҝ�m\��E���x��YԺc�6<�3~��r��|���*����91������y��qb�&9�Un����\�������f����V�K;��WZ̎oL�i�\��tH����]`��fsݢ��ξ*��,��E���L��%��ИJ,jԵ�]u�w�Ӹ��czi�����.e*ّ6tA����|Vz�yT��W��A<��%+.+����%Y���ڥ�����U�����gX	-('x��S�߆���ǡ
��]u���D'�1���S:�	���m��:ར9ޚ�.��{�P�,�ڵ��-ak&!c5WKN�2T��G�{F�i�be9�WU���;�0�[Qe�?�����N���Orդ�:K2�#e�*�����o����A
�~5��S\cPm��bY�E|ۑ��9W �z�j�l]�+lǭ�:��U�s�E͘!����P�����h#(��S�F.1���LIPX�]��.�-���F��3�/�����ּ���J�X�nTަA����{�}��P��2	�#0s4+8U�ƕ� ��2���8�ڲlބEX) ^��e�m�5��Y4f�K�ۥt�$k��8\��=W�	�Ի�uխ1p��;�i<X�xB���v=�:g]��[�9�ʕζ�ۦ�(.����О�*�9;T�IS��
SWk%@%	�6��w��ϸѳ�ulRT���Z��;���[z�|��©U���i��Uc���rq�3�[`� �DخXacV�%|�ĺ�Ҝ������>U�!릜�����me)}��{֪�#]F¾�gr�簓{��3��L�ۮ�뭷|�!Z������iڻ�Z��KB�t�'r�v,��L4�s�N�}fmvR��֗t6�IXB�7t�1qgg�Yl(*˝ݝ�� Ȗ���pV�>��Qf��D��n�-8����V��}K�]�6��u>�ȭ���Y甌�O���9�4p��ڗ/4��۽z��Z��"�M��(�\iK��l C+u�y\tR�|��XJ���������D���N*�ǳen�I��4�j�F����Y�}Ǖ��"�`�c�h�S��}ݸ��t؆!�6���Pl��_)���fl�7�$)xz�2��D��l[d��{w���Ɏ;(�-��eJ�Qg{V]�W��nV��yМia�)�l�N�Vo
�8�����mP���n���6l�Ғڌ��jƗ��N��8 )� v똨������ۋu;��l������Rud1M�!*�;څ�B�Y)�Y�'I4��wB�j����/��P��b��haa���e�,;_:Aν�Y�?���ZZ]����o:�r�R��ߘy�pW2�+���ooX3`�OZ7_"�$^�Gn��
�jw`�mt蔓I�il��V%$�_T56���޲�Uŧ\�TO�RC-���8���.�6�In�ժ�Z��7�J��+��L	Ʊ��ܖ�3X�����f�wwC4f�w�`�oy����}L��H}�A�j�(����㵀��j	����r��.��/���P�݉�l��\Ĩ�0"z�vμE��6�hY
�]ϲ0.�Ǔu �3,'b����mHA�t�������ד(#G��p%��De�ᢅ#�Du2���h��Z;�g�l�C`1�,�6�$��*+9�`27�Xk
�$Zenh�lgR�o�cU|uH���)�� sz��7��"�r�P�����-�n���T���%�H�[])^�T,�D_K�:���(�<E��5��%��r|����s��c2C�iގ��o���H�:��� J�D�ظ����g�R�J�'��it��R�Ak�����ޫ*���uq�˭�
�B�QY.,����xn�{���FQѸ=G)� �7!�*�n�Gz�SegH�S��wa�r)��*Wp=��f�� i�6��g}x���k:�݈9�%-;���>D8������S5�3�ےโjK8`��1m@��+-󻷭�N�����i�_ɚ�ރZn��0�H^�y+#�:�6���SV�t��}rM<qk�
���a�Y���A�
,C$�����b���R��w� y)�	7zH��%��jr�|ʾ�q[e����
���Ԭ����v��m����G����G��m�����r�L��|�B�_��P��;ї���/�1�l�}8Ղ��O!�j�.o��Ht����E�C�5�!7�S������*ܫJ\ǆ���B�%;�����sN��j��2b6��X��l���Wk���YS�gQ�=��e��oM(���������&�w)������]gV�՜oA�J�K�:�����#sj�=V�F2�v�c,q�6R}����ֈ��'Mw�)h'9��f�Q�*����w���1���-���ul

!��t�'��$��A�Fs��i�I\��o�6\�[��,�J�7j��ĕm�B�_v+��j䂻k�����u�Άݐ����fWo�[��D�d8-�Y�ւD�=�N�ӹ\e޷}���IVw�̈́<��-V�c�jc���u�C�Tٙ��P�G-��vs�I�(a��_ؘ��޺<�X��n��x ]�n����}���GMs������ƍHe>`�N�`��堦�.������m��+{B������z5�M5�ڐV3�!YW��|"�B]�oUh�(�D������Ǧd��բ���yǊ�l��;&�s��წe�w1h��ν��Z
������]#Ѷ����&(������-�gg��v��5[\L �q=@Gϯ72;���6.�K���=�yޱ
�f�٩/���7��:�g"�����l�*Z�O���q��wjj��3RA�N=�I|� ��gf#Ŭ��^&T�;!�~���jk��A,��8��8ފ�=��I�V����D�ƐY&R+�J{�Y�KS�N\�tV�o�+��5q���8E䊇|��8L�sE����xA-�e���ٜ1��yP
]� f�
4 ��:�tJwo�O+�����<DoXy�jƪؗ���qZ��{F�!Yp1�]�u.�{�ϸP��B�:�ti�Y��s��d�utU��M��Mh�wiT�;뽛m�הp`Pb7pr�\H��r������S�m�����i�/�����`.�z��� �M�u@�,�ss��<�j�I��er�@�7��_㠜�vx6ᢶ��b(͖�Z2���ߝM��P�8�qu��»��<���p����{&���N6�l�`b��=A�� ����rr���뜃���V7��N�3滔��D�Wo�BS���ePޮ_Q���]�ʭ]"��>���W҆ՅY2������t�fp��d:�z��3����S�Q�/.��%w�)�2ŎyB��"p�c+���t�0bV3������J�ѹ\�18N@,�;�\���8z��[;��r�w|��8ևׯv �zm����B�_5�*iG;,)HR�o8�ˉA�>e���c{B뤑�1.�b0��P4�:]Yw+7l�:��MHw4��^��h(v�tj&��!˴��M<Sv�}ՙ�t���p�#��`�Q6mƁ	V�GsF$��(mL ͫT�lȷ��VՀ��қZ���}�F�us�{�eu��q�A�.�m1���m��,R���Wn�8���R:��B7��T��[��X��k/���@v�ݖ�[�����ʲ>D�De���N{Z��N�s>]�Q����*ܳ� 7n����Q8P"QoU�;H�rV��vFܤ��j򛬬��lC[���t�y]QiR�Y���>Jn=�´[�&K׊���_*8��H �*+9�9�z�P�6�;��C���*��>�Ց�OJ�[lVA2�3�ZB���i��v��t+/��SuĠ�P|�c�U}����|��b���ĩo\VEv��X��葈����B�,i]}���lJϸ��ɔ��yS�w�*K��}lr��4�<�V��>��YV-ǽkE�y�ĸ��W6�3cN�v+!����/9��`q�k��mёdǋzVQT0�vw�V�:��Cf������B��y���7����ѷQR�5��km���v�g��1�m:�,����Fu��������]g�T�@(=ǄK�yL�p�`]�a!�}���V��}����n��8��YŤNʏ��E���b��Pu��i��˻�Dy�ǈ7W91pێ�r\��ʼL�^�P��`��m�b��>��N���E���,[�I�-��s"Wf����eC/W���	�Tp6�Q8`b\��;�����wV�rn�C�m�D6�9pU3A�Ц��s�2�Jk�vg0ev�y��;9�7�媴+��͊�fouZP���ݜSF��<nF>^>���[[7�^n��3*EN��2�?�� �m&;:����ޥ8�zhk�s�9���6ook�x,�֧�S7�[��Dm��6�\�wkcr5CE�Ŏ)\��˚X�n� a/�]�e�N�[C-�e9׮��k���~�B����yf�N'��$m���
{m��p:Ԓ�i�9u}�B��K�Y�,�v��|���؛�g�h�Ô{9���F�U��c��rT��r'gu<�6��DCJ�x�!��[#�P�s�l�
B2Է'e;�c6���|�5�w x���֥�h��%�9r�&Ŝ/�������`�B�^�H��m6��9W�-�����J�68�Ux`d�mQ Nv�_[Y$��-��s�|�8]�r�V�yw�XI��WP����U�f��6��մ����\�?����~�����6�,�]s1-2�*D�(��n��eX�%Vw$�̜�hS9\C2#�9Ҧ��$�*\��ЊB.��D�Ù�"�D�̪
T���T��I	+-r�	H����%��]MʶPU�'Q-���%�	���+%�F�TJ&U�dA��Ȫ�N��.T���-��.�xe�s�	˚�At)F�EG��֥t"��UQC��²@�wr�չ��:�aQh���Aj\�������J��S��ʋ!Q��)��X]0�(��ºe����Y�E ��t�D�š��R�PEKp�9��̰E�@���tuB�,�E9R�R�h��Td����j�Q�
���ԓD��I���bd�9���Hd#E"�
йuYV��g:H�d����L�����ݺ-�bC5fu��h�\&��<���v8%���|;����y��p�v�\#����;�.�<��;z���9�(�!���a��.�l�5�2Uu���O�p��R�#"�R�w;��<Ń\ �y"�6�nW���UǦ�Y<�嵛gA�]ʰ:�KT4Jڼ������Gw�^���Mk��s?Tϥ���۔W
�8k��ȯ�3c���T�2����K{Z��.1�����
6g>Z�+"Q�� �9%q��"�[O&�R3��4�mk�{�P�3��5s��0���29�G��鯞�X�kl�����Dp���pPr�{�ӧ�git��i���� +Φ? �:�����8P������5���e�`�^JΝ��]�\�ǰD*�ߍ�
붭�ٿ��+\����'L��b���w�%�Ew5)�����C�R�;�W�w'Mϒ�|Ώ?����W���̐1񌤝�<1�S�Et���l/�P��4�j�,�b��`ը�}J/��LM���L��qCu���-� ��X�<���� ��Zr�H�ɍ�q��U��ZZ�y��*k7��N�Bǉ�+po
�F$J#+��Pڻܭ"�Hڢ�y�����i��G�9S���\��nTp�3{IQ���.rũ�+X}k���w�+�R�f(����(L3�������&��f�]�`I����Q�ݓSU[��9g:�]	�!�UH넓Ϗ�����m��p�[���a�Iߎ��G)���r�u�X,�t�q�ɍ�9Έ]DD�u���j��q=�r�-��c:q���⪵��a��ܝ���$6��j�t����=�.8H��n�:�P"�-����85J��Q[�*�@�B�s#�Txf�я
��+��]�6��\Ҩ���BdT��2%�T>�X���}[� �~��T9Z�K��th��:>^�F�vW����<�/��Q�s�wygM^��mB^֢�����$�J*��
sȎtkl��h�=�g�і�;ùj:�c�abT��>=�c>�%Ҷ`l42�5��x��~;�5e	}ygyn���B�FJ&�LLGl��Y,Xr�|کP�m��M�z�y@�2T��/u���G��W��'�/}��=��
Ⲽ����X��������3|��e��#��!��s�W��n��@��3�f��yK�~(Q�Q�g�z�Fe�p��Y��u�V&��u4;y�������h�_[�^5Px,��ID�H�*����B�K���9$���e7����r��#=b��
�h������P��)ؓ��ٯ�#�z�;���ՀLLA�t�U����m��G�r�f%�Yx�+�CY���&wl}eb<�a���iL�ݴ���4a��e�@X{�L��|�p������^�,UW�+�����5�����;:�d��(�G���̔�`���"�������Q;*�&u�M�t���-[�5}*Շ�/6�?��}�;`��L�:,n���_��(񂠭��(Jo�7�Ժ�uwm�̉;�g"ć*�)ȍ���LH[v�?g1/�c�\j{�2��,�q�c���`Ll��r��]򥻱�v\EV�1R��pC	]Ts+�#�X�x�V�����MO>�R���ɪ�<�
�1o$*��b7�&R�&�2�D�?!Q������p����7p�;�� XR�\]�2���;j�-�6P�<�1ǥn��f��j�7�&}}�Fw�&�Ԙ�Ǿ��	��.;��oN
�v�Cs0B��\��� �/i�B�m�,�\3�n
z�u��]���TU��tn�¾;�Q��0$��j��ίL`TB��ʵf�ʌ-�ŝw�۔���u���!���;R�1��Nf�%�GSwd
����]#�{k�:����^�Z�5�.��S�-39ǋ*�#�d���t@sAI�J��6��U���k�\��j�T>��e$pi^��+#t-���Q�-�)�t�3tK�8T<�hb���
\X��������U�ړ��^OK�$Tb�7xJ�
�ul�r�OM�s����#eZ�r�.���o�&���ْkԋo���j[/��bT6�ܬ��I���Y�����^S[ �﫵5�[Da������sɵ.����^y��5P��"�Zc���_8f��Y��wU�-����2�XXH�+>��vrvw6P�s����F�e��i���BO�g 6!�VZ�E���_@����F&��-�|.U�+z�ߩu����:%�V\�7���H�Z�r���L�P�K��P-���,Y�A��b���jJ�E�̜;��.�	sˢ�w4��1�1�-��;5SC�O�dq�l׼���̎�J��fZ* ޯi]]��Л;��C,���i��7��4#�KKF8[�t�(�����0%e���M��%�D�덑=$!�vk�3��9�n�2SU����N�*]%�����XʤEM�ǷHh���8_+dVN@-tV�Q�>u�N�ӕ0t�8qp�j�y�Ϣ�0����N6���q�W%��ޤ��9��(i�\���*�o�@����j����K@`�ԁ����.�X��/��"�eh�U5�P�(%�*{�X�&^�o�c���R�)�ޏS.a��K��#�f�tT�gf�Q�,G:Fb�|z�:��n�P���;c��E@8(; oK�T�3�3���3o#::�an�pW����&�;H�}�s9~�L�a��%�#��l=h[�ݫ.�ص��5ݚ/�WÐza[,%U�4�5�{\T�i`yU���(�J�櫱�ů��X�~����@)V�|���~�o_�Sj�!p�hEe��ހ�*�>˷�K��IF�<��� ]A X������<'��Xk�2V�\)�ox<��v��1K��!��l_j����"��),�Υ"�ʆ�y?�\4�'�d�X]�S6�}/mf�vU�Jg6�I$�:]����� q��,W
�8k���Q_���AK�g�3<�衃���PV�f}q�</��d�u̷Rꂉ��H-���}\�*��nD��b�[]�:�ƣ���B�_��58����9Q�#��G��b��DR�^��ۇ[kD�K(ݸ�P�Y�,\��]�:�
nH�����mV��}��39K�9�w,{�:��h���,y�Z�H:܏\�Qm���gS��K����ٞ;/qt���;�t}J՜��=S�m�<S7:����Zn�g�${�nol�$9���q6Jm7}}�3���R�[��id�nN��rE!m����Ҕu(m�%鿤�)g�_X����V�l�mJ jϺ��ӤN#����6x̕�/��k�P�n��׾�l�j���e���3����u_�����G��"�\o�	2Ӟ��W��N{��6P{6]��+���dg>�R��Pa�n�����H	��w	F��1�΀��ԗTW:��NB��e2����l�5�i�=>�@-.� +Β����wj*��M+�w|���ɳ�D7�R�N�we���wM�/�«w��F�+b�Y�Z���L�Y&t�-�]���y��`J�6��M��J5�wW��Z�.��4ݻ�)w�C��j_gI�ۦ���e{��K�wY���SѴW��t�6���Yq�B�=Ǜ�@��B&ͺ��}��͌��� ��?]`��F���2�v{�H�o�~ba��Ha�=�JOy�*Pz*��-�
��@���\׷%��jh��b�ϯtU#x�n�97�h��ō'�I����M���t8���+(�o�P��L���G�#�p��/$]���34iߨ�KRC��@G��Y|�x>b��(k������-�iq-��u������L�CLש`۳d*'Nh��h�C���r��5z72�� !ιS:�n颓��1ӇK�C>MӾҔ�wQu؃�!Ս��YfS� 8x��yȣ���^+������y}]�CNd�4lf��}JWd�1H��	S71m�ω{0�c(yZ%�ƵʺvLJo�[�	5|�/eFe��X#�eqʬ�/��)���	1Me|�� �p�q����<��z����`p0���$+��a��\�� jYL0�+d�C���f7���Y�����H����_Srt����{\�^���VR��x<�S��v����An��ݥ���RE�^c�e��(>���4����2���{�*���]�������a.�㻭�|tb=�~��>]qWUӽ�pZ@�YجX�~G5��-?�3�����L�Q���8��?[�s�����Ъ��������Y4��#ϯ(�Sp�^��e{8wG����A&^�|�=OTPV2Z?\Cj�;��1<b��,�dA+��Nk�Z���S>�7.�@���,�� ���E<�;A�%��%�nX��Z�SRT��\��q
�e&����S_��a %)�r#2�'�:{{k��p@�XC3i��)k�xpwK�.��-
iI/��`Ř��^}�n�a �6ӽ�i�_*���x�AX)�R��vY��Y���Y��Î��Qw;HP����{T�?N�3��^\n�t�TS�%�Ӂ'cv9±�h>���H6����3����B�x�bZ1ǥ�鈆��<�t48x����-��'g��Ż���6v�,	�pU��q	�A
��o邂���|a���VÒ!�wX��M���^ur7[��3�2�Û��\c�"��R���1�L�! TB��z	ݺ�<�'�T�V,J<��_�a��I�ϋ
��w.fu����� >^'���g8�{�P��������å����i�B���3.��3����ϋT��yctɃ����:s2��/r��>�KA%�;)G]��a��,E�b�^S�~��?	�f�-����Cf�ok��� ���,h��U�[66�M�q�=�
�B|^�x�.�\��É��ܰ��W���UQ�����@YG��ḛ�ܘb��a��V��>���sW����e�*f���䫞�Пyv��ݕ��n��%�d�
�1�+��CP0��謫�YSغ��6&�͑�\F�`u�b)�ޖ��tf��ў.��ĕH���[�T`� ���+�����g�l�N�pg����|*S�E ����i&�tsy.$e�JK�ßD��F����Uǲ��ܮ3��xxݽ'"(�p������Z�1��uYi�30N�˜���p-�SM�R;tw�J�� �a��@���4�oU4c(��o/�Ae���T�t��R�EBҰɇ�p�q�5�w�R�d\϶K[T�v��ϝBc�a��*'�q���$/�V����Xz7(�;H�w(��Vy���ȭ���J}R4婅u�vT�w+-������Y��}Lp��-NQ�
@��3�k��(
SFY�U�}���bv�)j��VBͼ��*��M��?1�n1�Ni��uPE\!'$���(q�YYA�k�x������K�(��0�fG?�_rv��p�YF�#EC�b��%0W�jm\�ոݎ���c���#�t��.�m0���y�>ϼ��O�lx�7U�C�ݷ۰������7m�ƃ;Ak��0.1��Pw��e��T������
}WS��ʹ�+�gq���H�ڱ�R�~�� -;lLLR��7�ݸ�5EG'z��:�����vSԟ{��4@� F�ŀ:��dRrD	�oT��l�O<E�����g�o�͚a��$:�/P��]h��l���k.��Y�b�F�Q6�`8i4fEZ;����t��2�ӥ\y�a�Wn!�p)ψ��U�n�֦�ֺ�f7n�����w{&�T���5w�w��y������<H{n�w"5N�w��wu�Ê�{��rQ��Πg_'ڴ�ٛ��7�(��$FVky8q��[���+����(C�W��[�	8}d�yLn7:��,�������>O3>��0��fp�7�p�<���4�+�fJ)([��A�=�W���3,��o��)Խ|
��p
����/|�WƮ���ɡ4�Y��3�~h�nn���< -�#V-ҷ^�w��Z��y,	��M��i��hۑuɮ|��b�a�êC|��H����`�A���g�pB�u�H@[��v~�N�%+�++��fq�v[W旴���/��s�N�ˤу>���Ԉ�xC�*���K��H�����ۜ:1�7�xwӳ�X�§t�p���#�0��u��\���Ѹ@#(�F�	�uݷ]�;�G�S�j��ݳ	��ua�,�-��0ާkQ�`�7��L�#���0�B�������vɸ�a��UHn���������<�Ҧ�}�lG��T�"C�y�gs�Z\ARl�I�z,�+rY0�֊ڿ���8��_JD�33��$���ݫ�Z��2ڳK�mP
�B��FH���5p��1�gk��LS��� M�������x��v�ȑ9w7-)ii�U:�����հ�ռE���Ֆ���oN t펳*ƋX�d�i�8ճ�2��7cpr9uur��싴�nQ_k�e�W��֪�|�CsG[��fY�U	R�]����O;�*�ۻfbh9w�k�%Bt�n2>���uW��6�Z���dJ�ms�kw���	n�K.�2:6�eǝV�Oa���E���t��(�͘�j傦oV+h��MBeb�6ﲒ����R'�CX�mV_Z��j�˲�Ǔo�Q��vd��VB�έ��O|��l�*�v��%|:�+�Z�u�gQ��Lу���2�V4�-m5�N��j �=�+���c�,�[ʘ�s?J��oT׵gaD>:�X����L�kW $-���ۙ��]�<�8l���dhe�}�����wf�e��;t����L���˱�j�ǰ֖n��B�u�ͮ���Tˤ�obATx�+JG[P.�*�Z��3x6�4�{�{w�n��G�b논�s�?�m��C9Y�L���N2aT�0������ǥ�Q���Dg"�e�r5E�S	�ǀ��L�U���-�ޡ��W{wWsZɈ�}W��ǅc�(�w9<�!���q���y+nY|JǬ˧gM�}�+1c��r�+���B��}��-Z���93c�6[ji�J���˹]�ƾ�&�ը��i�tN��z[ߌ.�%%��G	�A^Ŷv*���I�ξ�8���eN������Q �Fe�ij{�+��J.�wHP��u����e�nWNU�me6��pi��ͽ��t4����S���r����ێ3�]�Q<l3���V�r%�j��V�r�*��1&���c���6�E�%
�TS�T9:��akP��v]����21<��aU��.Ի��,���K.�T9T=S^�-��b�e���wݖ�n�/��#r� )�W�M�ph��mv*h���(�v���>ݽY�v'"���U�>*f�u2�zιG���7��Nzf\��:X�T�e�F�*=����o�8��"�&�4����d�*2.��s)��{5p�7Z�q��c3iV��_m�F�ڻr�4JdU��eƤu��ؽ�NFvMl8�,�[��QᤷvlD,��I�+/�T1=�]nd�C�\��|�u��3�U1�4��I���8��%��V�I��p0��ϰ�,9ubñ��P��;q��٥)w��dy8H?xu^���:3�c�ڇ�n	yI�<ޣq�t�X�S���޶v�.j���72wE���2�O���x+1�D;��	0��#k&h7׌W��N�[���j�X���n^RyS�2bB�e�BL�keJ+�,{�q��B�=�d�z��W��m��밐Y�����jė[@r{�΢y�]�]�}A*X��fh�d�������)������>���=��:eP�U�!+J+�3.t��C��EFAuX�RK��j!vEgD�3flJ�A�]�L
�TRt��p�Ds6T��EUYӬ�d��2�9.w:9�G,�)+R"��I"��3�')Y���0��J!���̠��C�r"%Y˔J-8�RJiPT�t.Y���F��%��3R����	&(I�	.V��a� �D:���UQKj�b�QVa��QQQM:�G#QJB�ȩ��2+�u�jH���z�AU�A*�.�B�蘰�D �Z�T��#����:�W:�EEĐ����J�2MiQT�Tr�AWL#!g"�����W*�6*�(N9��XF+Bt#�L:Z��%*,Ȕ5�J*uh�9G�g��+�?(�M!ZTN������/���ןߐoJ��e��\���iHd�s�8�&��s�o��oh���_96��}of�	�{2�j��]�tW9���w��;���uvt�K��u�]�/�)������0�z+dM���w�o ���!�>'������ra}���������F�C�ğP����������]��@�$���߇��߈��H��	������j�T�Ht��rr�-&��n���>�=;�i޾���>��L.���$>��7�~�\
o��9���<}8'O�?S�]�97�A����r�����u�� >��������yp�=��R��3��ÿ���w'�=&P}��Ǥ|~&�og}�����	9�M���{M����W��� ����z�c��['�s�܁�'��G��.ܛ��z��%p.;_������;?;�������������_��}$?zy7�~'?K�����7����o�&q�}���7�'��Ͼz��������o�;o���:w��������oG�r�M|���u�a~'��c>���DCD�}�:���,�����Y۾��c�|D}��~�� �����C����9�O���o��P�|󷮎L.�q�|�ǯ�������<������{��6��	�������q"$}�1��F��{�~������|������~8��>�#������oJ����z�����S�nOT��Mu!�����7�'��|��s�����������}�{���$8} ����E�>�>�
p�[�z��1<�9!�d�s�#�|D�����Dx�����nw�?��~����I�S}O[�����&���]��ې�����=&�BN|C��)�!8�_�>y��M�	=�}��ǧ�['�s��}j܆�h����j~�����]��������!~{�i�+�w�����MϷ�!���ɿ�#�����>�A�0��~p~��ߨI����q�C������NӤ�����)�N��������`�$DH������w���n~}�����ۿ����7 ~$��|�ͦw����{C��oǕ��G&���v���<��!�4�'�~X������~A���n��x�?���_��)�9��V�<�`�>c��3��L�����������';{��n��'���>��i�P�q'����i����ؕߩ�o���x�&���v�g�o�x��k�=ymɿ���,���?����(�a�is�J^����ͣ.�3zC��3EesjRZ���k������s�j*��ÊQwj��er��6�#��R��j��ư�vm�X��	�r��6��	����4Z�
뻡�e�.�R`���S�t �#��l�8�����[r?}��$D`����<���|L/������oi!�]���P�0�������������>�'�������9��;��>��}C�av���!���8?��H.���>���dЯH^�����b>#�����?So�>��ro-�8���zM�]����xo���>;&�>X�C�뽻���>8�v�?]�������%p�{s=>P-��G�DH��i��M�	(��������=z���;N���o��7?\r�� 9���=c��{C�a~'�Ϝz��܁�_w������;����������������yq3�����r�!�`��D�ｾ͸�c�C�i����|��_a�<M���M�:L"o��z�K�;L���#�|Cӿ�rr��;��7������\8������{L/ջ�߽�����_>7Y��]�^iIz�x^k��3�mM�Z~8���HH~&����яI��;�y�ͽw�1�|O�8��|@�ts������W�叨x�P��9�A>�>c�B$}h�s�W5n)EV[�����_z�} }"#G�#۳�"�
�߾��]���v��n�H.�~&��|O~!'���~|v���'I���Ǥ�$�֣�N'��o����܁�'�z=��x�&���}��{�j:����ng5=T���!�W���U[~;�~ϟ�`��^C���>����]�}��&��p{;�x���o�$�}��x�߉�|}�Ͽ�c�$���z�zw��r�c��M~���߻�|��������d�z&����3}�G��=����&�1��"����3��r;{yߧ�v�o�O�[��>���w�o����v��<L-q���#}|w�|<��
)�����7�s��~{5;�bN=c7�������""G�>�NO�@s�;�O�s��������nC����<Wx�w����=!�4�'�~�c����C��^�o�O��8����������7�N>���̔<�M_�vL�%Ax]O� ���C۾���a|�c�I����o#x��?S�}N}'����w����C�
{q�܇�x�8�?,s�Ă�w�z���=�}I7����}���TG�}<i�+���ԥy٧��{H%-u ��P��K\T���3���!��N��ө�ErX��i9�p� 9Ɯ*�ӛ�)a=��d�b{�3��1vn��oV��*������8�s�;2u��������,w�&��z8} �G׎b(}}��������H{M }I��}���v��O�w[;�Ą��巴�}8$?�}y=�����aw�����o��>��r����A�}�#�}�b��KϞ����0��~��������Ǵ�8���w��n~�����aW~���}�7�=��~��1'�?HRE�����'&�������������~���4}DC�=��RLg��Zޠ���P��f(}榇�}�񏘡�'����\�����ޝ��dߧ߽�!���|q�ߟ~�c�s����~��?P�0��ߟ�c�r�r��;�C��׬�}I����~������������ws�c��i��1h�"#D{�1d����x��k�������]�P���?ߜo��I���}�����*����7�������������}��OI�ސ�=��9?��������}{XV�ugS;ڴ������"$}�?n�� �����XP?�M�<=ǉ��v��P�{�x��	ޯ������c���hzM ~�߿;���EӴ��;����ܮ��=�M���m����SEz l�ʬ�������D1�{����i�>'&�o��4����9ǳ����M��0������?�N9�N���ǧ���7?P����I�]�]���7�90����������|v�-{=�3�1Ƴ#����D{�",@F�;��|BO�n��W�����O�������;y�;z�[������s�aW'!��w���2��?���=|����0�㾡��{�OK���]���t������0Dh��U>���$��������>8�w�}G�RC�4�={��v�����?<	=+�M��|��ӵ����u���N?_�����I��� G�fW���b�X�5v����P��x�����=�$<C�ry��]������Q��!�>!��<��T�]!���w���<g�����[{@��o����9�v��S���W�|�C>�>�9�H�39�����^�߁'!�4�O����E�o���ߨ_�>8�~~�rnB���[�������?�q����|NL?��|�o����`��?{�U��'���I��������>��~��}>���~�zW	�&"��W.�W����9�Sv�Z{}j��:#��(ҥ}��/����x6����T{�G`�!]�ܖ��I��w]�m�{'�7���)�̀���:S����}|mh/�q� h����;�#]D.x F���̐ b��ꯉμ�Gk1���!�>��?E���@��Py�������}v��?s����x���w������7�$�����oj�Sx���_�o��������:���y��4/�,or�1��nDUʿ�}�����z��^��0����������]�Ou�!���s�S�<��&;�zq�>!�ra|=w�>���;�[s����Oa�� |I�=�~���|v���Ͼ�|M��8<������ɕ�S��T$�D��}��>�?X��N�~�OϿ�~&s����>����ҡ�u�M�?S�'�-�8$>!�������<L.����ސ�OHs��9S}t��~��&��{�������M嘢�f�,�F�#����߿<�����nL�x9��W�����o�I O���=m'�94���}Ov�t��e7�/�o��x�7�/������ć�����ߩ�s����I�VNǱ�%��^�4w��p����������9]�w����&�ǣ|���{w��� {>�����t�����<Ǵ=�w����wF�97��s�9ۿ��q����"���|v�|@�B�eVoާ�3��˔
��o�� |
oo��H�1�w������ۼ���;�v���}���߉�]���8�M?]ɇ��������s�����1�=�x�a����?�_�ʄ�a�/ծ0�X`m���F�o���������r�H~'ށ�ۓ}w�w�~&�S�O[���=;��p{<��H|MV�>^���������H~�ڦ�BW�}��x���9���}�N ��}����>�Y{�o��BP;Ѣ$F���~�����>��Ώ�����������0=�@�,�
��rE�{H@Y}�b�Rxo�-Χ�B�~Ǘ1+e����1����}-W:���x}����@�I������귚�
>�w���5��W��Ȏ��Ip��S:=�K��h�^J%1��kׯ|���h�ڛܛ��Y	��J�	��*���[fvq�̜��ԩ�XH��2��ѭ�ќw؏3b&U�����ɉ�f34�� �9^Mz�w`��ՉX�	�Z�8�$�`ۘ+w�aӺ�:�Ud�9Fk7����U�C����_�����z�e�.�!��?_G��'Nz� ��xh9�7��x{i�,��ޗ��%+�G/b�L�f7<���e���&4T#\c/�U��x�?�Z]b+���owk@�' u/���'��fC�i��㌴pg�\)�9�5�;�����y���ѳ���P	*�WK�tq���p�d9�կE+s����ڿ�5���f`lu(̷�cT��1N��FD�	�ݬ��k��FI��kvh��=������}�Լ����r�dڨY�E)Dn^����ܑ�
4t���C1�b3�B��xr ���Ӷ^�2��Bp����=�[���w�f=�`=�ހ"�I ��I���8@�����\"t^�=2�B�n�;y���m���9 ���b���9K1�Zs�ϵ	d�T�2��2�g��k��Ds܎n�5n�q�$:1�~�YLnGCyM�Y���٩Sa���eq�ׄO<�F�jUޤ�vϭՎu�^�,�J�p�
������NDӡVM˔��Y�&8�*����~�w2�y �kY���ק�T�T�W�[�:0Ф�uM��lE$��C8�ɇᬎ�%ʀ:v6�k�CTCv���B0s����Y�}��Ȯ]��hr�w�p·�3���L�Dvv���D�7gW�}_U){{ܺS�u}?����m��i�����Evk�+u�3���S���w_�������K"�r�9�0���wyR?���<��9>���̿k��V+ߣ����öq�+�"��}�%I��'��5F�pڬ�v�C7b���[�L��|�p�����T���\�O��-�M�T���b� �c��yh��&Έ�/���q�fۮ9&te9+XJ�n�
{4��L꘸��A�:�총�n!�&W7Kw���Z pu�ڒ�I�����"�){+n��|�����k��&w���G].�PJ�l����c�����J{9Ж�읒��1�ݮ~�~wGB�^é�� �w�&��
�]�xU4XΙcgGE ��@���ov�]�a�졷���"V�^�]���j7_(�6�^�jk�=`���u����Ǫgv��r����$�|]5���\�0<ֆs�"W�1T*�����Omm�5\b���.��7 G#���ݫ�m�A
 	d�#X���@C�T��r��:O5�/�N�[R��V�(|�L�j`Ǚ;�T�J.��,��\�ټǇ�*W�Դ2@�08a�Lc�ϭ�Nm[opd>�m�����:=�%w:�[���B��H������Zm�Ky�S�7�2�R����W���T:�V�i����b��;Nf�f��W���8 �+��1J�I�T���]�ӭ�YW/�y�ByR�����0��1����!�eS�PN�n\�p:(�ZGwR�ޫ�C�q ������4���B��]��6��a|��g7�5+��Gv�\�_8DL����eL|�|Oa�|���o0���vMF!��c�3�8�:������P0U�2L!I��AYv�l@�9<i�<2��ϯ1�^/a���)G�!u��ys;�[��H�7۸ƹ��2��/zI^����X�\6̤k����gu@����<���R�랩۬����}�b&�;���<J��<j����YGLX�;O��*����-�d��Uh�ɡ���q��s��R��uG}���,:�cc};�m]l�:{c�D�x8�P<a������&���(\�Wъ@�p���,@�V���$}w�^bC
]�f�#��˭��(Ի��jiWx����}�<���^�qׅfBb�Q)!���5�x֫���X;"*5����3z�M�]�5 ��&.��j7�`����츨(cW/%���;9�p��E�L�Bٹ�JTB�=��i��e�Y�9#s����[�jm��4�ќ��f3jN��=x��(Zgv�xm�z~��ﾯ���y�=�5^��1�<��p����	Ỉ-N��ܥRQY�]osϨnX��YqO
٭t��[�v�N�ܫ�;;�y��R��Wօb�5d�5��:�%��u����i����!ŜE[��x�$�������r�T5V�vM"�i�L@��7/s���&b�fz��Z(8�=Ƨb#]wR*���#㥳����䇗t��v8����C�^�0{�G���R��=� s=d#R��¸z�騇1�����t!dO.��xur�c��F]c��*�ϗ[(ӑR���>&�S8=f��\q��7j���\'ë�B�u��˕q���8����[��3�Y� ��d��1�R��7����*��26s��ˑ�r:�p�����l�n���(X��E'$@��A��گ��pb��;�l{�.��Ń�r���+�5'm�����z;5��.{�-�vQ�ˉ�!�F8\��h�Q�ﻐ#\_Wήq���ɨ����_9��S�S�ύ��Q� ˔�]��]� ��\"Pb��	�� ^��"�:����z��@�֏AMd��7}�L�:t����n\;2�����Z��p���M�m��b�KsTQ�U2F�;�M�UƵ�Z7ZrJ1�bG�_]�+ �����C�!R�d��)D|7����.ޫ+vd�'���V����lX��+S�����G��+�aN�!�j��6��a�[��}�u]��R����Zدz�B`�kqmu�c����H�:�P�䍊����#_��Wt���޻f�#�^�5z�%ajg�f�n���I@NȄ��[0�v���I�)q�����o�=�炻������7>K��Hh���20d�A��}�yep�1��1�\��H�F2�'o�C��ξ�5�9CC��z#dI�%W1bu�#���4W_NE�� <θ�ݪf��	��uad��p��e"эw��U@E$"p-"T��{�Km���q9 FT�?T�97<��eT�ӯ����q�;����C����.�W�э����0�mC�Tj 䁽U: BNE�enBK$E[�/�m_��hD�<U���:DMYǲ�Q��09�������WQ�<�a�*_��h@Nr���U^�G�5V�YIO�.1�(:S"��f�`#�w�6�s�!~IX<t�����!���Dd¾^H��n<sk��9\�ȁ

�t���l��Ytؚfc�8��Mvl�m�sOE�i�Є�-�JQ\� �5{V�!������ɻ��1$�+9�j\��R���To��/���2\��������>�������Ӗw?i������(�L�Ӏ�n�J���D�"�t�&�
��[��Z��E��ρHC�P��C}Lm'�e��j�8�X����ؘ��I���y�M�ql�y�\���6�f҉��ĭ��ϙ�騉R�x��
O����w�H���'�(��K�����cG:M�l�V9�^����
�M�	�B�3Dp��cz��n;t�BL?�[�n���@��ǿ{~8��++�]瞂�����Z�x�굕}��^��ɒ�K�(��D�����'L�%�rR�]f��햬�F.�"b˙�^�b�59�K��@�'#��Z�0��@X{�N���+\,�=�So˽<�ȺSͧ���ǕK���=n�;d��h�����¡�}1V�EG\�v~ )~~���޸w���0[���'\��#�#����N�7<�ӂ��P�+�	���I����j���E��-j����TU���D����G��k�
�KG��4u}e���;�P(d�p.:�1˺��8ɫm���u�����P+�$6��o���"�*�%r\�J�F�@��$:�s5�֯����c��}|�\"��fV�c��s����@�/E�9�+C����w91� Ae��o�|n\ ar4,���c�t�Λ��ˁ7�r�vޝw����ep��l�us�ދ4ޖ�s�W�딸�=�v��	*��(h��u»CFI�X`��:�3*P��X�k���a )�7%��y���rM��b�땮!Wv�s11�!�n�oF��qUg�q�jZ	��k�dx�&��ܹ�\��.�w�kA���t �f�-}'t���W��e�q$y�x�+���*�d�u�73���1�δԼ��?:�(V�mt�G9����hw� &��kV�����Y����m'�M�(ұb�Vu��s�*-��sjqj:T��$xj�l�=����y��^K�#���#��kN#ٙ���}8��4��U��Nf��I�ڰ��17�f>��^9u�V���nU�.҃1���X�}'^^�+OG�u��.GB���f�)&~֦���/���G7᪰���<�/�z}����-�]�� vd�L�\�u��YI��+�c*��d��1�롭7�!���E��`�u	a��l�*ܩ��ʽ]ܜ"�'*th��p�V6l�B:�P�;3
�<�/��	�yѼ�6��}�c<j�{��{�n�ٺP�����MQ,�/����� 3U��Φ�u�oj�n)����:1C�@�69�v�gL����\�Ђ��5}��O�l1�d������Q�Q4%A2U��+x����֌�/�x�#�]�ܓpg={Hv�M���+n�%���v̭��J�kmb�$P��}�C%c�vX}4���3˺�u��q�Sk�#{�.��z�
3[�	��������U���>���w���!Y��׬]E6�K�
�Q��5��+e�HУ�2jΊ�1w֜R}��iK�8��B����ۛv2�]�B�N&���kZ����x}9iГ���-@]X�ο�+QW]�D�v���m�s3�N�!.�2��գ��xNrJL��w�	������J���U��Ծ.pz �iu�; պw5��\R��t�Ta;�1�P|B����	!�b�U�R��������mh*]��f�R��@�S�6T��j�M��f�B�7���U�����ٯq�:>�T�\TN9v^�ה���˚@+��!�du�2_"2�:�G��|.�3b�̧S��+�ֵNc�S�՗N�u�c%YR���.�oE
�VǮG�|���k��8�������.[U��6�_K� ��k��L�`����!}�e��Q�u�mމ���C��P�Ր��d���yk�4M���ܨitU�ق�Y-��Q͐�  �X�Q��.�A^(G.Dp���d'+��){�W"9S�!R��TdQ˔�����L�R̕�R�:��EDI4*9(����L��+��D��y%�E:�]�G5*�r� "-7�"��9DWȇ+���Y��Z����VR�AHL���*L��EV�E��+���y��x�<+��E��r*"�L<���5�Dj�bf�G
��UH��RI�(�D��DS,�U�&ˁ�.UEr�N�"�9�|IșP�F�AUJ�\(9�Y�Qr��J�PU'Q#�(��!��,�W*��[�Aa9�;�
��Y$�eDD\�3*J�\�J8r(#�T
."�J�^fF��)¦JA^�^�H�J��,��a�U$�G'"��k���:���y�(Z��Ri�j���H#�}o�3�'j�����'E�s약.)r���X=Rd�&sF��u�;#v-�����U}�}SS�gW�ؼ�(b�?���G댃$C��UH	���,��0�ڮGk��v���Q�cVg���'51��J�������e��Wz��Lm�9�*�־�iw=&����Ju�G�7�_�՜6j����Pוp��Y^��������&��"�	M|N��TK��k�Q!;k�u.Vh)2�z���}��r�i��"9���X��؄ꠎ��(��Z�W�	�s�N�[����:�_��7}�����wft�C1�8t7#
�yd)���#�.�g1�Jh��O�ю�*�ȿ�*�>��kF�����-~U+I:]z��g��͐��L��*#^�E�)d�j$�(���Qx�O���{]i\2Q��X���,��r�bea���]�db��\��<�y�*�uIvJQ�l��~�8�F!����M�,�7�����`y���̈b���-�`��,@!�<b��h��s������Wf��=s^�䩮�B�Q}�A�ڄͷ�lbuE�s��[wp�\�?�c���Y,DL"�ƃ�^���������ȅgn��#K:��Su��:�N_5����i��hw����^-�������r��u���Dn�UC�(�'9ܺBW���]�}S�����'�(�WW����i����৸j��Py([P5��=�����꩛�S��6䂅��j�~[��T�EI�鈛�w[�G�Pg;k�k(�N*�����{'���y��LHp4`ʜ��?*,M��#\��K��wC�\���w�x�5Vcu�ڻҟ��mBl׫���픫�U��ZU���@�Τg}����܃���S��2�|��;h��uò�Adr��TZ�b5cJ����x:�_]<��<2U����a����V9p#t�q����sZ/��~>�'�%W�a���Z�#ùH��'\�@¼��ʼ���ʢI��w	����\�7�9�c��tƋ�+Ŕ.��1Y+�_�`����mɡ#����z��}��W�|��LP<k�\<�M��O�n��(EC�v�t�U�ܦ7�Hng{8����*���<�3��AăF/�GW�xh��O0�N����at�{�v���i
]0E�ɦJG7蘟����y���+��
�꿦����D��K�<,�j��^��g��l]���pU'ˉ���rR�[�K�pz��^����o"nE�8�t�׍Ȇw?0sA���,�Li�"b%��`�<����k=���{4M�%��$��3z_u��������!�fU��|��J�_J3��3v�/��Wx�c�r\(H`��:������⚬*�(c�"cEv�]H��^+c��w?�}UU��w�}��z[���}6i���e�� �"��"�c�Q+O�L��"��D�kn��͛V%4�����1�&b������-��P�W��)9"�cz���o}���T	mg�<����/��X6���6���DU�$/�X��\�J j��9V��[�~�(.vw{���B�R'����z�४�x���+�O�iѡ���on���SM�@-5Ϲ�4�]/дwM>ύ]�u�)���T�Y}wݾ5�uS��K�k�rr�����G���N]�
Քp�����8eD�Be�B�`�=�@�����}��wFV���]r�Ou�v�/�¨{���m�bWXY�R=g�t��(lW:�y)Ιӳ�[���*agE�m�]�؝2�|��u=�e�^���p@�fu��qG�3
4:'F�U���������s=I��\�!���ۇ��4T=�:{H0����:ռC����Kw{N�@���	F�[0�<��%��۔���`�:b��6���Ո"�+h���h�mos�f�v4֡���٩�o	��1gmH�� ����H��c�[�/o��J��RcJ�bO���@���v	���DK���Q��9��a���}�v��i�&�E�G�W��"��'�� <׳�7�-fE�8�H���c�kk����ﾭ^���z��P�g�V�^-b��� ���6tp���������r�;��E;Q�E�˺���LT�E�㸍�^��U*@޺�F��C���Nr�"&>V�E����q�3����ױ���0�V|�bV��0Kv�Μf���F`�	L���<�aω���zp,ś�h������Zˍ�I��([ `��uH	�P����WM	��s��j�UͲ��Ț{�����'������Si\Uê��>���׽0Nz2P�yj1.(��^�{��H���S�mz���dƂUg��9 ���&+�m\1�9�f��% swD�+�۽mP���3�d�K��M�A�öYR��p��G�կ\]`���MIS717?>,Ӽ@�)���ZW��22K����2��t���n�s�,l�҆�{ʬ����E��3��6в���y�ؓ�|k��A��*�@�ϼ�$+���	�%���u����}өEg #@/'�Q]'!����L ���<��9:�2���3��*pK��&��N(����M���N�@���b�U����X\/N*��[���W����m���Lz�.d���]5��!Jԥ��]�-�ok6s�{�]8@��V��+���$2RU�b�U�eם�I�ewo��E��M��ҙ1i�l�<_�}��}U\�V��*����y���`�,�i9�Zv�u�d-R�o�\���T�ͥU��/�F�Q����؞�~��V���و�mt����l�-�n��M_���];�^w���j݅�����-#�j��Ѯ'gҭ,򨳘�R�y�s��!�ei�c8�LE�v��O���c����U
��K\�8�qW�M����GZ�Lt����n�#2�R됦]!�R�) v������Le��Y��L6'd݆<z#R���VǶ�[y���6F�M�ƞ#�$�fP�q���^=<�ALbRM|LF��)W5e���t5f�9���
�]�������0����}���M�CjJ+���<04ka�������;�?;Ͻ}�C���hp�2g���dCrr7��ђ�ƷU,͸���5Yu���3��N�Ё��Ԩ�� ���1u��޴�.f�n �L�s#�����oqH��sj^Z<���שU�	w����\lT0ٵ��k�*Rs�|a��v�9�Nb�������U�W�^U�֧V1�L���^H鵼�<P���h�}~ލ���"���~�W��N��I���Hd����&�ɼ�]��v@(;�֣][@h�[| ���ϓ�2w��:������kZ�I
���\'�]4�H�g~���>��	%�*�}������r��=)G�:��ҧ��W��3B�c�')y�y�׬F,V�vk�����(�@=^T�x,��}>Q�l�y��S���+��<��w<�����۾��mئ!7��V]�0��'�s�2Z�Q8���`*ڤZ��z���]�w��� �Օ	����1��q�,�`nfuɲ���͉'=4ѻX���{�jm�=U��ɘo�,X��L橈�T�s��*��6�b��h�غ�]7��XHJ�����(p���\dЎ����q:�s����f��gw�ǫ;��8�1%���>��m1H��HBB�͔,�a�11\.yc���HilNI��봆t��b��2΍�����m�b��$S�IWx��k<D����y�ّe�Ѳ�jik�u?k/�lF�t��S_�>��֏z���-N��|���)��4be&��,�1pGk}B�}�p�)��
��<�v;�4Z��A�t�e�I�WY��~�n�rG�ճmI��ܖ������� ���3SCøV6ܽ�S�[��M��b��jl�9��ڝ]C՚mH��4���ǹ�ZE�Ϟ#;��U�*ڟl�o���M|��eK:�QS����v��|s9ԙs_�U_}_SM)&g�x��]�Ϣ��5�"��ȫ�LP<k�\0���٘ct�(E9�l^%�5#tl����p����@�v@�t��E����GTB�&�;H�8S��Y�ڜIy7�����q�(C�n��0�H��1?)��5�=�6UC�,*y���nh�;�-z��1�8�VmWu��ON�y�M&a��呺\���t4ƃ?���K�Hu��w��w��Y��Rny��{Ãt�����!���̂Ab8D�Oa��@v��U�j��z��h�7:���곋h؎��v�L�[9�8r6 ]�,�NH�0a��qz�V�ʤab���nr���!�_VɨҴ�7�S))"2�;6nTG"^]�*$����v�GE��ڼwާ96K���:1���|�����35�(;Z�w�f4���\~��;�+c�����l�ʿ|2ٳ�r��4����F��:����Sn'B*wu�[���S(_.���cJP1\!zO{�b����9��c���v�M'Y�YRz#�{	7#�$S�`ة� ]���J!�M����IܥX5�o�8�u�v*3wz����hd�r�`�I9y_�,�{��^�`�=B@Mm%2�m���n e_u<f^�g]բ����� ʱ�h�l�q<gtBrRp�-7V������{��wNUk�t;�˗s�20R�#�_U}U�#�x��������wȈ��8P��oٳ�ݖ���������LY�
������絇a��sE�8�_.�g��L�f-���|!��X�n��@�\��Y�pA{Փ�;8f����Uܟ?����\7��N�KK��-�t�wE����:�2�;��6�v��3����U�V�7����2�0�LW9��VnS)E+xs�w��^����6���L_�$	�t�>�@Q�rl�B�*�;����8�G��λŏ����jS
���4Ug7<��d�jk�5�-Ҽ���]p����t"�3v\��S�7�t��V�Nn�'�_��}�9��a�WgN3_�䌓�+��1G�,"�^�r�җ�$�Uw����V�~���#R�R�]�!���r
�:S"�n��Y����BFz��&���Z�pR�xp�Gw���mM�\k�L�wZ
r����#��� Q��=�d�x�ٜ�5�V�7r�b׆|{����^B�5	1_S}P��8������22ne����vb�M�箭�T"l�ҭr�:�K�]�;Fѹ#7]9�����])9����'�=��"���pv�d:hn)�Z�Gױ[��b��h͹���[�[�/0���X�ڝ}9���4��Y�_��꯾;���S�i��d_�,�f���<��a��;Ml_h�\0
���>)HY=M����;��m���l�ǤC7\ �Q.5��<C.�ʌ
�'`!����N@�۹����'���lE���@����w�WB��?^D`�y��ąq����Y)MF�k�K8��[ۄ ��K\$��=�@f�g�1c�/����.Ӓ�mr��iT�c19o�{O�)��b��{-��`��d�ai=T4����@Xu[�K�Z�����ה���r�g�K����W�ֽ�O�*���,m�N�,E3����&Y��3�vs�;U"�^>	WA��ĩ�A<�氫ɝs��1A�_e��oi2����ܕ$�vV��d��fu�.�<e
��K^P��
*����]�u�m�Y}=�*����@����G:U�G�W
h�0��ًM�~��&>=5T����,��.jQeD���-�{Օ�z7k��X�x�V��nXۅW|�Ґ�h��u?!���<�kV"��1�V.ٙ�s|}�߹�93�j�՗�r���kx��ggc��� @�zbz�v.�!X���'v��n>��4���[4��*���y��b�	�W�͗�;�W�W����Y��Y2�s�a��u׻��꒟V^��3j��}�W���b<}�&x����Hk/r%q�
���u/Kӹ�Y/�1gd���B�{��j=7܊]q-�����<�-�,m�k�������9�����p[�R+��^�	��܃Y��`��C�e�|���Us/�`�;�m&n =n��v�6\ƈ�s	�[��95���$#��B�w�09�lV0����v�JN|���!���8����,ո�i�f�Q빎`���,����2�{_�<���1�E�iS�t����̾�&�Jog���ŮR0\��Z�V�*C�"b��[�`-.��J:�U�����1�٧�{mX����z���y���j�N"����6��]Pa�M��<c	A�����QC�J��7��NRGאz�=�f��c��ڄͷ�l'2Y⾔>�?7U�h�%ҝ�Wo^<��'oT�$���۟�1\@�
�gh�U�A��!�P�A�N�8���<P˛�/2�Wmwhq�Al��rl�Y1��2�)�";nX�7��9�X�5�1>��#u��f�(�PZ�}�#��;n�U�X;fӔ�wd8kGM.����ȝ(��{;�n����'+g`%N�4�n�<ދ$i�dN�5+ʾ�X�}����ݗQݡ�e�������X�G,ٙ�x�<��t�^��$S=g0��2�[�Yϙ��oA
�A�A��}wv�bfӔ��bٺ�a%�hP�)���l�W�Ի��z'o���<��	.�u�2�R�փǢb޺���+7�=S��$��(nn��b5j�H.�q2��H݇	u�KV>��õ�j�#��k���*널���[�݊wpoV3GJY��O�6�h��ɘ�^Ǖvu���ܛ��t�@� &'�;-hC��6�Z�]mE��i	�K�/Veh��E��(�a�;��҅�6o��_^�l��[�ڃ��]��cZ�T�\����H��z2E��X�W
��CX���s�[��Q�ˀ��c"��T�W��!X��V���%4�Y�%��㳌|����m�	Dx�ֵ�:a�ڳ]�;�-�q!KÜ���	��b©=AT���x�ۭ.�m�S��G-()ұ��4ƶoh�����Ƕ�]b��nH-�;;��)� 4q���૱�-�\����L(1�Q"�d�B{�V� N���zr��ڵB��ս�Y���R����{)5Q7��.�W|h��y586�, �U[��'�:|��w�#�=��d�m�He��,Ӯ�:�}�l���y\���[�g!Ƿ"�~Ϋ���Z[�Տj�R.�% �3���D�3Y��"���9Z�Z���ڃ�<����gS��X���%�~N�/� �,0��˴wZ���_�����+���P�dVx.�s&��ck�(�b���*���I�u�̴�_E��лx���*�g�@ܘg�2�M��:3��0��^'�H5��A�\uq�YŹgڥ|�pw8~�pCz��-n&y�����S^gρQ,�5�q�Uv ��u�ξ��B�$j���%�خ762���PD#M��M���ۘ��,0����̲H���-V�*�Mޔ��Y4 F�յ�PU}�{y�θ5�H��5uo[b�ĺ���dQ�Oz����ӡ�/0GV��R��m��2�n�(�ցj��Ғ5$������l�9-ҥ��h��L������𽎸�+%���\X;�흃=;{W�Gh�ѯuṋ��(�a,���L���"f�(pK���07�;/:�T&���2�k�ݜ&EV��(����j�.�C�h�s�o�����9h��Y*�T�3�ޡ�(��Gp������ oTN�!�+P��V�oݠPffi[N�h\�?�����q�Uf,�t��R������a��7�%9"�,���	���"rJ�������w�!��z�Pj�A�2��B)*�"�#��(���g:̬��p�A�"�"(��N|�h��;�G9Ap��I�	��*��.DV�T�u�N�U&B]0��ӡS����u"$��0*��Ȯ�T�"�bD�*���-K7P��/Z��r��ux��ҹ�QP�*.w�*:Q\�3ѕ��49��wZfgT�%��Ni�EY�r�*��r�s�V��V�H��KSQ$�.D|�p�D�x��<���s��W�$[C8�%EUY%U�\���YN�p�jAUTTT{�95J�fY4�(����s�V��(:�w��yBu���:��Q�8j$�dt�:g,�:�f�/�.t8�UPU�Xj<g<�F�E/.�s��UR�u½B"8Uz�EEr�ep�0+�D�~~��/?��G���&*-f�WR䱭;Z5��:����)C����V����v�����S��W�X���NG�a�o��W�}UR��&����������bȼ���5���G�{gʸE��ZU��_/��9��e�#�eZ�sS��Q��	��1 _�t+�5���5�Q��R=&,F�L�f�QA�}�U�γ��!�B������:ۿ���e����>unC�co�W`��W͉�5%�1Vl��n�.ټ{s[H}nc�A��R۸L�Қ��O2���L�eKR���9B����k�Nk�k+�����%�y�.֪�"��ȫSI���E�g#O�n���t�o�1)��w;r7�P�U��{�p ��7�)�
*P�Q�H4c4��S�D�D�x��ݕU݅U=�M[���@o��������%�0y�T��ֲ���7G�xN���u�Iwi��j�|�������:����0U'ˉ������V�.&��pz��t�̈�49Tf4ޭ������])(>2#`s�`�N�yw*f��ِ�O�����3��xXn(���J�7��Cw���Ɋ�m�[8[�#�� k�z�#�H�jv�M*|��j�J��I��{� ��"� ���"�O皦3qcn_^���6u�j���j�i]��*��l�V/vg���cX��g�܌8�NƤ��^�us���kq��`�qtcC�k! �W:n�b�"�R����.;[�8�/I�A�p;էcY��B�P��\�h��|+(���ozꪯ���'�0�u*�*��~c+輢:��[&�K��cťDF�G'f;�7^\��N�on��R�����%e�P�!������3#fw��A�y���9���9���)M��W��g��?_���U�#p��\=]�1Xb��X�&�A*hE>U���*�@\���܎�V)������Oi��1�*'*�������mv�ސ$��{�V��q�H
(SrE�	�!ڭo���Qp;����o�3��W13x$�m�˷ђ#\F�;7S�yN��i� �
>x疻���n����[0@���W��=���y�M3hne�^����f1���9�*�e����L0��ه~�(h�a�����f#3e��Ep�0b�\�F��7��A�r�m�o'V'�Cr�H�l��N��p���q���A��S�e���K��
��N�d�BL�{;�樗��U�c<ʬ�����e���ai��s��O��\+%u.e��lo̲k��Vy��B��k��ʳ��F�0SOr��h˫�&<ʶ�H�r�G�|�#)��V��]�8b���BZ�K ��6�/��ohF^0��-X��oqK�ؒ5r�(�Z�Z�ʎuJ���ov.`�X���7a�8�h�V�$2H_K��]@�U�_��꯫��.G���H\U����m�݇��0�n�C��u1_T@�#0N�*��L��r�|��n)�}v_��
���\p�P��qoe��ҙ�3p�Ɯ��������\�wv��/6��=��{��|�|�iTW|�2��R�u��}DV�3۫�֥{�=�Ŧ��K�C@�-�1x���@����6�����b�.q'��cq�e�����/R��F���V��O��ʮó�
u<��᲏;z�달UμU�>�?�q6����%g@��T�}���W���K�rF�y���A�Qxb5��>���
u�'%����coG������47mG�|�`B��O�O��,��[K��JWwT��'�7v˶m1���H��`	�JXb�9��q���u$SX+�d魉��L�:|������\�
���]}Qy1��e3ӽL ���d�&�Ì�u|]x�(w Wj������Ϣ�}gA��,v�|���=ے�f#�],m�jvɸ-����ǧ�3��ؿ?J�6�ꏭt��2�0�%-�cQ��1+����K����O3�y]�0W��g��­�ۙ>X���M�mI皘f������Ky��y�
�O�ͮ��S��?D�']�y��y��͊��9�;w��T+up��}U�W��m���7`��V+��舻1yX!���'g�>U��q��_K��531�����yU�@uʒ(��>��t�w?����>n��@q.�*����]�U�쾝I�{�����h�gQ��T��yO���錸ol����݆=DjO�{Á{Ŷ=o�)&e^p��Sz�Y�Jg1]��fƁc^V�AQ5WՒ�{F�41��r{^[�q]�}e�L���+{p��E�!q�%�܍v�n��RQQ�')�4�u�IA�FK�;%��a����Cg���\^�낍DIWɔ�dH�q6���$t�i�W�� 8�:� �r`��똑%K��7v�f��wft�Rr#m�	�2�?m�z<E��������No�"-я�J��=&��,z�wC2oEEr�i9�K��⠜����s3�3���Y gȮ<k������_-��~�A��x�ps��v��Hm�b�`�Iճ��59&,Q�� t�eiw7P�C3�p�D�Ӱ�^���J�F�:�Y�I��)Xpm�W)"6Ȧ�蹼�76����"g�<��H��wjx�P��aW2ʘl�u�R�z"��DP�� ��y��)n�{]LN�G�1WO�WU���y��s,��&Q+�@	Jp6N0���2r��Lu���j�$�\����覆�>�ޞ��\>0<		u������BX��a���X�BG�'�y��_'eY������2��7)��~O}s*]y]��$z�N���%�����VNtV�*.na��{-�K��&��?lǆ³�&<.��X�N����(yL�N��E�=n��%�Û�
��v̦��E�E/��6����s���j�-�|.U�+]E��Ϸ9�s��X�(�1ւN�eO6[�\�lmש,>ª�l�����ڂ�!��l�W����*ү1N�
�����Iv�gEYu�]z���-�|b�\���o5�Q��R=&,F�D�&f��� ��j��3��<����!��Eem��hRb��\r:�5Ա����ڽ��/&u�d��8p#Ʋ�&{|ۛ��k�2���WD-���})���K��������P�c�	u�k�Ư����H�΁�7E4���ȥ$gI���]6r4����9W����U��S+_}�����@f��ê<�P�����؈��F��=:�Sl'},7T��yMZƮ[k�0�縃f����:r�i���Ȟ����F��S,�C��qV���39�<�N����n�J����Y)WGy�ŕ���d�U�a�(�n�#�u-����o�����t��+�������]�R�Y�_PM�Źz�WN�r2O��#ﾉ������U�wC�f�&�Sf�q�j���%�����G��8T��n��d�s]6�[z���Ѯq�j�<-��*s\���}�ʎ�@��YS�Gx
�*CXqrx}`{,CxF7�gJNϾ�wM\�+�����Pϝ*��@������fY�d�;���L�j�ň�ש��Ճ+z���i�7n8�!������mH�
 ���ER,�#�lNp���gD�<j��?`˖��9�/a�3�cEBRDe.w6n!�@4Xp�T�:X���n��Uo>�U �T����y@�[��K~	��'[���Ww�3�U=�����Iٲm(�16a��,�v�77K�W�d�H�AO��T�qXb���*�R��ʈ�TqU�w�����d!�V�p�jO��V*�ol���e#Z-�u���<0 ����_;�sťR/�V.,(SrF��b���d�x�,��>��9E�C�
�v��F!W׵�o�,��u�?^'L�"����|"���3��+�K}�T(;��Ɏ���QtZn����c-,���w	��z��|�I����Mk��Y>�U��0w�
}	�_�)�c��z��ɷ���'q��A��/Y��o0��]@#�zM>�S�.��ur�z�p�w�I�K8 ����}U�}J%&L�]h�W��V��C�W�f1���c���VcsS��4�-����IXyZ�B��'1.\��c9�4z�+��� D��q.�wUZH��a2y�Ĳ���l7��b㯳�R!M��&4T3\c5Lw�$	�_N��e1S���O!d̆a��)�X��ϱ�u���������x���P���U���A0�!<�8b�$t��A����E{�O<\sj��q=�r�-��c��_w�����Z��e<���^Q�
��93f�oRˎ*:�9�l(X�J�St�%���[�9��X�٬�2�k������ˍ�-ҫH�(f��qNf<^V����'���3|���8,|�f@� 
�$��,:���ϯtUy��H�l�G����ǧ��]_R�T�g(�P�쳒Jܠ9ú�_�%%]�e(�T�#�l?N����p���x�{~P�0���N8�����"��y}�2�(=\�&���혍`�M�B������P^�Y<��̨��Cq�YI�7`�+5����^�.�P\ٳ�n��<a�e�6�b�M��%��U�����-)Y۠���A��Ki�D�e��ՊT-��Y.������c:�r'�.M����YӦ<#Z�2L���i?���着nk�g���j��+8+rŒŹ
��5@����p�H#5��`��{���	�%Mu7qN-���;�F-���Y��ɇ	KN#���������^F��V�9nv���<�^	�{���WQ��/';S���&�6.S��!Ř����]�.�
w!������}	P�v�Ê��;q��Q��=�ls�͌�7�w�ZMk�ߨw\���U���[��VOa��D/Z���zon�-z1�������.�n7k��������PU�*.+Z���5�F���yc۾���]�)����N�>Om{��߮����4�ԋ�c�b[W�*U�0r�?�;�!�'pS�z[ˌp�n{_%V���m�S��*�nH'�Թ��f�C�K/�Z:R��IC��_[���<����!A�oh��i�p
���l5Q.f %��;�}�J}!���N�`0-6@�欆�:�V/6���z&ׯ˙�[�yz���1Ѣ�T�Y0oތ�ֽ� b��(�sŌ�.�q&Qu��ݞb��8'^�uE����Gt{�fLub8�s�ftv�φvvw��H���vZY��][f�����a:��I����ﾪ�J����h�WS���YWڃ	LWL���.��Mk�2�mX��N�eG<i�J� e[�'	tE;�6
���9�V���t%��%M���t��ν���}N��7]�Sv'��	���'��L�Z��N~����.��o�QU�����j����CD�Z�q�-�MoU��S��I��,ם��M�r�s��A�RU6���t�+�UJы��f-�Ca��g�'-����K�Ey�},o���>�W�h_Кkv�h�yrj�*���S�)M?�]�毾>X1�E�^NT^/q��j��ۂ�jGl#r��5=)���J׾�/7��k~���Ъ�.$(��v��r�\'i�槛����ON���},���S�L4ͼ����s���+-�ʞH�H�αe�E��{Y�M�x�nB��n�m���X�u���ۋ��b�Ҝ�ˌ�:�+R�P�����d�G��y��C��N]ӖÓ��33T9��ݯ-�7�۫�o��8�*���Ֆ���*u͆��Wd���n���;g^0;7�*�Q��v*%ݼ)���fɝE�Vw;�)>�&O꯾���-�;w���Z��������ŭ↸5���ݔ��F.��s�H���+�Iz��7s�gv��{�'��Kyx�wc���=�y6�TU�.V�{�-�q�i�郑���I��eL�}���$N m߆����잾�.���6��q�.�B連z��s0�V�G������y�foL��<�c�K=Ku-qؗ��&�%pͲ�K4�S�t������y��6��]-�%������[���Z9�Un�Ҕz��Ζ�ݷ�{����Z�K��>ۿ}["F�H����a����b�g���/����#}�W�O�+�+]��5����@�����p��D���l��4eN`X�Ɛ���/ �������<3��r�������!�M";p��ۣ��u�r
�x�y�
��c=�e��wΥ��,c�9��.�9['4`QpZ=�P:��FMݞ� d֜<�;`ۊ�L�����-;C�b �p�%>�VK����ev�W��P0j�&oc�}�n�4�I���n���/Ac�6ZPp�M���yz�U���]Tr��������hט�1Mٖ����ܧU��:���>0�@��;��4���lV#s	X@��3zdޕ�M��g��}�$������N�|�:#�b`�*��G�ȗm�<���u�"�}E����{���2`�c(̤�廇���g�|>�Ў�lw
W��H	Xݱ{@�"�I��t�W�\��:�8tD'�0����\R�r����V��)�+���+�(]��u���{ڡ�S&N��g׺�����h2	�c�x:ufÑ�o`u;1�Yj��������R��B�)���Wt��;��B�q��FV��1Tu.r|������Y���v�T�n�F�o�����|6��4�M������lh�&����p����E-tBe�Kkf�p�#�_�k�$4]���u6KM�Lˮ��_ �yi�{�!�]})�``"2��!GlL��˦��;�a�Y;���#�ۚ&����,v��s���&�܊r諫���Y)�!��3Z����*�rm���-�L*�w�F�E�1�
����WgN�l;�����}0ڍI�����1.�׽CYr;��)M"�U&��#uUI3�m�pܴ�4���wA��!��.ө^��^au3��7�m�Ű+Y{��em1��o�í-wMrt�N��M�<��T��j���:��(f-Y`1ƺs�I��6��Z���	�"T�x�\�#�j��ZW:K�i��GR�L�y��ټ��q��Dv�n�"���k����:��
`�Z�u�Ν��L��J�攥�e�U�n����}��Uʄun�%�wTUm�j��|��F�x��u�J���3{��!��y��uz�*�M���;�r�����2%ʍ!2nKQh���3�#��b1�ژt;�yqM
��� Y�jHį�ڃ�0���=�8�[� Q�4�J��9g�0W3'MRt��ͭ�LY�ެ�M.�gE�t-��M!(])����v�Yٛ��^
U�Y�
�s�Y�.�m
t7��11_i�-���]��l{o6�qr[��Yu2�@ݍ� �,#}����@MҢb�n�1:�n���L�0v���oT1�]v>�Xɇk�[j��{��P��z�m�/V���g&�ԡ8�t���/,n�KA�H���nb������lr)��o� ���C��H�e�'�4�⮜z��Iu��CtN&�%��35ꑁow,�GBR[�fvxi�Z ��t.pT6<x؉bۃ��̏^ryB����E񂥓&�n̖1�z-\�v�f�]�g���R&0m<�p�(c��i�D�����rn���D�u�~�VŻ*�gKj���E�j�:r���n�b}n�(��lHjy��u�����ኂW�a�Ъ��xJ1B�[�r�Z%UL�#9�9r]ܠ�L�B=sv�'�g*��w��)���(�hAɅ^HWT��g7'Bԣ���r��p����Z�S��G��ǄܫJ��"����n9��.#�;���򞻋��ONbIωp��*�^:��rJ��OS)$�Y)Y<y��D�(��%w<u�������eNI��^���'���R֚�h�|�xO.�G(s�)wp�'<.(bS�;�{��G���(���^����Q�s���R�A��N;y+��S"$y�k�<<�E9ϏvXT'��-̈��1g"�lu̱"(KZ�7\u��p)��t'q�*����X9�XPT_"E���vaUY!99���sbF�_U�7P�.z+���~�;�����e���J�.��J�gs ���i��8�!��t�Aa�T�|���bs;��8�7]L0s�KpC�UU��M��n�r��/K7�<��f���=�R��C�z����d���^�a�CRޣoB�ht�۩�oV��PW`�P���R�)�I{�Cgk�{Ѯ�9�ڦŧ�����|篪�^eu��N&5i^�r��v Wy?z��؎Q���U���O;��ب�o/��j�v�2E|�K;���qae|z�Է7Ԫ�:6�\U��M�����%@@o�t��hif_m�.��y��R�ֵVy5��<��a���J����IO�V�j��&�[Fs��v�Gc]J��c"�rضM���dy'>�=I���N�����M77�L-�P�FF�D��I��ڙ��sx�{h+ı��·�G�K>N��ݥ)�q�U��P�����0���U��t�����&g��&�<O;��&��/���ſ��"8M��YmVB���#8Eh�2����.4�a�Ja��QO�ɜ�i���{�E��� (l�Ɯ� R����]�Ӗ��-�ǫ"��C��tC ��w
����<���:��t�	����1��U6�EL`�w]B�3'
<snQ=����u�s�n�b�?UUW�I�5v�}k��1���Nk�B�vf_OZ7��:	�}.�+o.y,[��Ƕ�g�y;�P�Bj+��[�p̿����cb{�����^b��t�����h�w��������+��ǝՓc�R[Oo!z��,�9܄�}����@46���iuE�,����N��N�;[���WZ\^p2��G*��T����S�
��b��4Z��t�Ʀ��«�z{���~7�������wW��:�q�M�5�[�ï��Fi4�.�u��ʃ��ֺ��ʎ���g8�Tش�p��g4���_mc���iq�Al��P�fTAV�*�}�o��gTk�}i�;u��p��w%�;w���=ީ���Rv�KKG{Y<B��ֺ�,��Ʀ�9��J�a.u>�b�'ې�v����[�zk�繽�Uc\7�sǩ�l~�k����>
����Tޥ��J���>��w�X��*�e6���~�X/a�;��/��R��3GG
��5^��X�jn�>c��Z�v��
��m]���ﲻi������@����Ŕe��8IA��S�@��{�K��u��"" T�C�V5�9;蝤��;�Ʋ�Mn;z�����>������WLX�$h�zΩ�\"k,8�ΖRw�O��o.1��m�)�W��ݚs�:�t;]��9��0���÷�
�k/壦�w�[y�n��qy=[�f�X�b�w�p{�̗�Є�ᐕ}.f\*-s�N�}�L�ޓf�>F��no� �KB�Rq��N�l��]�%?WL�O�]ojkf�l��IӴ�c+�ӓYR�'CY�(w��-؟�J<.
�1�b����U����<��3�b{�;ú����;����i�����n����0V�|k��V2��Â�.����/��f�Kv�ʄ��$��jY���4&9H t;qd�U{:�u���J���i߱�������r�����jrk.p5xRF��O����
��+r�7W����Fj�j/S����)��l���^I)�&A[�G�{�Zk۞k���c+܍>��4`j�	+Y8�+����\�5�i�m���gQ�2���o*VoK̭�J�PMMR��b�;�4���Q�ħ���X��c	�ί,��%���t"�<��S��������֦N��2�|�����]G�+ӎ�����r���g(���M���S&w�y��B�����3��Uy����Z��kj��ڠ���ۜZ�&*b�M<GEF��Z�y�6�6)��l>���[�k�fQV��U���+�='+�k-��q�-䕝�:��w�Cܸm�5�������1֓��*od�{iJ>��p/)k�Ϝ7�E{8�j5\��ן{�����ؚ ���Z�y�����w��֫��.��>u[��i��m9ۗsyצ�m$�X����4v8�z5Ԩ��Fwr�Ww���m�B�Nqw?p�kq��ݼki�7|l%b���s0�k�M�˴<a.��Z��2׊��i8��e�R�sP�P#�Q���N�����ޗm�[��]S���z�<JY���{�^8�V�LR�z������p���֫��%�1�9��Ժ���Rݢ�x�Z��B���D��Pu-�� 4�lfk��K����-��{�*�˾Q o�/��������{���u�ug��ڢ��;f%�1����:����A'1��C���}��>���W�_Sf�u��I���ϑ��ٗ�:m.���[��&��Qv,���e��=��³!��Q� bV��b{��eG&5������jK���9q4��vk��]OF?�l	��	�ޕ�X&�<��r��bK3�{��z��T�z'E���/(�"9����]����ŀ�}i�E(=|�=��Չ
���I0���]�x�\6v�\;C�л4�&�~��t�뼏J1���X��G5��Ku�9ĆCC��˫��eF��j�E��g��8�e�������^���r��Ƽ���lZx�5�����[�����h���S���6O�*	���{U���9���_��r�jW5�]��=��]�o�zEs~&�m��Oe�my�>�~��rO�<��n���+c夤�緺�,�}��� ���jT�j��v��CA��[��v���`���w'��� �s���@���� ��]ʍ]�=GG2����Z-�Yث �{�q�;1�ٝ�5�1�v���������9�2�W5������('���E�r��ޢA�D3�̮Ш�e��`p�:<�s����V��_}U����'x�t���|�O_�^���|���P�A���P�q�s����IC�)�K.�p޸�'����\F8[���e��am�S#c{l:�i�][8(<Urƕ���Y�}G���⧒��ҽq۷Qڇ-�q�W�t���}���w>��;*T���.v��78�B}�ޅ��I��5H墠]SE�q]�3;�k%�]0��ٗ�6Ҟ�Χ]��E��?ӱ䕎P������X�R� �&��[�a<��˦���z�w0'u ��p�H��ީ�i3PU�T7`Jc���%m0��F�O2Ǚ"kr�t�mvV����M�$�T6���V�*��µѥ�7m��(h��⧋��<{S�J˸�8�!7k��@V�
����.j�a��0�X�E�iU���,5n
[yj��Fk�j/T%-�s��>�7u7]�s���Z{]P�}�����&�N�T�4K� qPN��hb�`�ݳw�#@e��ZQS]�7��]�/�Q*�����N]�����Փ��j���c���o*��e�o2u���w�Ʃ+�L�G�Φ�<�JGS�+��qwV�iC�E�$xY�YSw��(�����OY�J4"������q]E�W��8�|s�Tظ�ZЇԸ�reTl��5��(��nl��v��.��Ys�Qo�b�z�뫬�`�Q����p6��2��B}�WN�����z-����<_�b�G��v箜<載�_+܍M��o��]-��OI�7�m��՞�f�i��>��2�Ŗ��W;:�\kO�;{Jv#^�EW�Q{�o�e��(y;y�������TE�U��N�|�4�{��v|�LE*�Yӏhh�x����tܔ,+���%�K�_5������E�c��&Rڬ��+�Jy�A�dd��wI�q���J6,�K�Df.{��*��Hg2�5OR���gPz��7���2_���r�\��+�`'�pe��Н��Ҍti���=����ޖu8w�Sq���b)!�~+��1�~����/ggË3�k%���oB%��
<==C����x ��:ZJ���u�(��]�[w��c5/��0龾*�{=�N�����S���X�6`��ż*ċ_/�V2�rј'N��0+ka�;)���u�[��$��DC�9�~O-E2/�U��a�W��~�ӻ���̶ym��=��@vپ����X����|�/T�
�l��{�5*{�'��@evN'��Z�*9I:w�}pUè��wO���K&%�0�e��$��ǥgU�8������p�M�7X��蛌�/Ƕ���=���e�E�*�{����黷�V<ƢujE�IB��5wy\�����)�;
��߼�\��8c������{���א6p,!,c���8ۑ���y�����pqn����+[=mh�V�t�wQ�[1n�U��^t����N5F*�q�͊ykE׼ߦ��mO����q�� �mj�u)�s��u��&��>!v��^5���$ا����n�j��:z]S�;�o�,�I�n�<����N�ʽS�Z���kq�פ1"s�MU�C��S�Nu��^�wTd�+x��U�Ui;)����
�x���.����.�y5|q���ė۹���F
.v����:�_6�l�[��
��wkUئ�F�t�	
�\��-wMvovG4\��S�1\*�bۼS!��u੓k\���F6��W�1t�a�9��M�}.��s�6])NhbUΥ�ӱ�X��2�G����E5��D��m�jiN��3�%�~O;�{���r�9�����
��3���jv\,����y/㺕�}�o���w��W���Q.f\:�`C�ԝG1N���=���GK�٨�M+�ꏗ��������������i�nĸ����kU����\2]���ݾ�;�c�c.)�pGQ_*�Xq�ֿ�vMh��xf_鴹���j�����wE�]�ݣ��lF�v[����7���|�{ͫ��otV�6�ۮQ��ӌ���\�ƀ�!������2�r�l����K�n��[�oy�_h�MC�*��`O!�C��:*)v��i�ic��.�c{�����|�B8�9�=o�������u�]�rvA�}Bs����oo^�Y�n�p/���7q�qpƇK۩�����nc�)�� �����c���������=E�s;l+-�g<�`�7�\v�n��L	�Oo{s�ʍ���6���[u��)]tRA�Ի�;@���鄺N����z��zu���\��'���!��=X������N�|9p�h�t���Wħ#�x�����u�������\k��q7��	�����vuU=-�����]&�8T�T��_u�*�.qW���(�����l(��ڑ+��2����˞��l_/4[5"���`t7>�sԪ#2K�|������y5PPs���=�6�;B�p���[Qpo\d�+���kV97V�M�ɱ�DJ��ڧj9�M��;��5����gۗ�uFAᑯ"Tr=	r���T�k�y�ﱚ�{���w�|�K��3�q�����|�O[@5��#.�No���o)���ۗ�w.w%q�͞�q�n;v�z2[��<���Sék�P�LGtjY=3�\.t�jK�/�����nuaߚؖehK֧�w���YV!��	Mt��k��/�)��ӑEv�ȱJ�9Ff�⺔�p3��[�4��]�ϫ�����ۈ����1���OI ��c��9��즭��[��)^D��pƒ���0�ݽ���}��-�%AoQ��X�X�c��&�j��hW�������i:�!C{��%P����G.��
g8Af���"����^#e4�ڀ�ڨ�Ut�<��H�iR`j#9ҭ��
*�I3y��6����]ʔd��G4�&�J�7\���eWr�zf��u[�S�Vj��D���9�^����;�]L��9k����sᮏl�z�e��l�igK�ʯ�������'fse��7\	���GoS{��Dܥ��GZ�1��ogu�-�L�F���vt�!�7]Zˉ8r�{�T\09ʸ(�	:��i^Zx�WE���Kxn8��uO�L�me5YP��xn.��l�|P�}�����U!����òH�]2U������կzZ7$`|jؚ�8�`ڻ�R��zEu(��׷�����VNqZo@���q�+�uj�\�t& �-_F7�Qz9�p'yw,�J��N�#��� j��A�3)4��z����9�MVh��2��#�kf�%�mة9�?sBS	T�!:ْ��R��r#o��-�lid�oӕ��7*���S�v�pM])�o\&wP��(CLt,�h�7:�Y��]neF# L��[�jȌi����L��Sc�Ė�mr��'�@j(/+rW&Jq��ݽߺ9�i�M��c��/�L<���l>n��T�����u�	w��-�D�\�sU�n�u�y�V� 0��n�U�)�R�c��U��tkwۜp�/��Ӷ2Ԉ�(�wl�k8�$��u���̍�38 �:�N�����0�*;���H� ��Bm%�����b�Tr뙶2����R÷i4�Vgq6Z�jг39�+�Z�XĠ����=��EC�'�7�n��V ���CB��������WD��,ػk`)x 1���Z�{@ǝٺ��x;��"�v�t�ж�#�`v�����h���a�v�HxNӦV�QI�ۙ7�e��7��[Oek��"�au��]lv�Z�4ç�q;�1+��9	�z^v�T�5���*E�͂���jc��qԁ�>\j��<*+�x��w�2�c�G���t$���)��ұ�eh��wQ5K�
�C���`=�g�����wbf�}����ч���^�z���O2ʺ;�'1O�ɦl��sA��>�0��j���Ԭ#w,�����p��-������z��{�k%#Q[Y%�K2��Ԃr����b��@���^Q�+v����%]�@/�<8��
�Wݻ��ё��Ϧ]�SsE(�I]�D�I�'$&p�Qs��̺�f��CvSi� t`eH�[�9K�=�1�G�"\`l�P�����%�K5�(6�����˰������	1W���̾�Ǣ��<w�C�G�ݖVrT>�[�BR�3��PlZ���	l�D:��K�wa�svt���_S:K��V�'�]YN�u�c�S����ⷅ(�
�����֞��j���ؑrGwdyK���P�9FH#˗��U��N�{�:a;��&9�a�5i[��'
"/���Kή���;��<��;��˜���
3-�ݩ�����9Q�w#s�Y.�q<�Yn�W���.�Ns6���<��K#��+���^ty/=ȥ۞jNyW��+0�s�%���Qs�u�E���ՠ�\�̪�Zy\�wp�V��F���{��C�UIF$Y���Ἴ||sW�� ��PHErvUG����U�-N�.e:���=b�X�A$�1*�ל�R��B���S���C���YZ�N��F�-�Fl���S�t�Q8u��(�e���:!��碗�y��ȺB(�q�^M�)<��.�
R+�Zb�r�T�L41B��B"����uܢ$��Fe&�虎y7L�2W{����������75�����v��n�]Fal�e�b��y����ye�N�I᫦����;n�����7�v����;��H�xz���֕��i���P݁)�9͡����㋦�y/��9=峧S��v�VW�QĘ�mC���t<����M`d��"Ʊjv�����c�Ӹ����̅���y.���,e,N�qij/��ؗ�����)v�{Qu�7���7����w;��[�g�t�Q�
6�)���+��A}�q]G��U��Gj|n3�LZ����wŮ���3�l�@w]���v��"�~�)mT7�<����m��8�٣u��X�v���W*���]1si�st�_ͮ���~�V�J�m��'��.y��i�q�fuE�l��@�u!��z���ѯ��{�g�\�nMm����W�{��T��yM�t����B|j�l�A�����7�k%&��[x1�j@p������׀7h���U�ƷD��b���YI�O����vcK6��GKr*f�>���I??['�i���f.}X��\�6euk���˿^T�N��R@}]�xۜet�ܹ-SN��=��:q@Ѱ/J�R�lN��+�	l\���r���@,�����U=�9�*y�P�k���z7Eƶ-u{�S�����G�Uk�jg�����'�)����#]}(�\+���7z~V��RҘ��e�q�Ml�d���}�Uo�ź�{l%�(�H����
�\�;���M�]�,�=�y�;��G<%p�v�qr��rʱ	mA��+�B|x�V��n[e���焉��ޏ���ȼв!8�Qf����
�+��s�� 0ڇ�lj���T��̄���ʄ�����i���:����/-���uS��m�i\�w�}T]��f�/y�*�J��'SP�����1�~��pK�u����n�����Q��%.^ͮ�z��(۸6�o�gE��w8�P�LRpQ�o��>�p�2�=�.���;{��uX��	��{y�'f�@]�'6���g5.�
��~�,��X1�z�Y��B���ʊ�}wjg_����Et��\���ͯr���֏E�q*�f��=�MJ5NLW����7�*;E�ː���s�����bcr;M��go���2�Ӹ-י�u=��($�s��:[���.�z�x�^Y;�3���w*�ʽa�}��>F5�w9�Mr<�����W�)�a�̛fH6�C�n��ƫ����n>�r5�L���J"�5.��~�!\��yR��l�'ތ}�2�c~YoCu��G5�i;yRZB��y�kj��|֏+̛�N\��uY�_Q�s��M�x�nB�چ�&qh�y\�u)=7�M.t(s����Xږ�/�U�L���=��Z���ojq�ͅU	�۪����Қ�+���=%���W%�<���=0L���1��N����6��n�ݟ;z���Ag@�v5Ԩ1)1Q��T�jH;gJb�-���z�?�w�"��Y�#�e�ߺa/�ȁ��R�u�=c�5
̂�Eٜv�E�#�s8Ǜ;���qڮ1�S���yK_vj�����t��J�W��3f7z�>v����ή�� �o}n�tJ�|b�c)O���i�[�Jk��w�]��9������z�o^Jsʷ	���m�A�6o>��	f�G�+�����f��6~���Z���呎��1O~>�!�<�Fȼ�s�T-��Yxl��tL=������#s�(P��j�q�=K*�]8�tbv���ڻ4gGw���*U�!�6���]Ns �Mt�S��k �̋�痯g\�iT�?WՇMGӧ�	[��\y
�ua1� ��Kom<3��n2�S̒��Sϟ#adq�9T�v��s�Ӈ�T���	�:�
�_AޛE.��l�FחM��<K��s���۸�!TC�v��v���:���-{k��{T��n�<�} :�����4ꉅj���ڞ�ͷ�fn9�l�'䟋�}wy�-�~1�J�R��q6�����4�:�ܻx���)5��,����������_ҮnqWٌ�(�����o65B��z)��u����ٮz�������ճ�
�����|f��	���&�C�*d��֥|���ry���s^-�T��k�\��	���:V�#�-U:+	*�nN1�3:�9u�|��5{�mm8ɥz���m}pvbF����:��:��p�����]CO��k/-�m�2�񰶛�qnÃ�+��I��s5<��U�m@�GAu�¼Wwg2��;����.R�����\ƪ��zP�NIQ�s%g":�s2�
�^$GC��º�+[��8l)�H}t��.���m}��RW�������ݑ�Z2�����]-�܁������eB��/er�H�Ǚ��W�|�-�c�)�n5�|�x�鵤M��3�=�B��fK��@��<c�Ҁ�ݭ0��k�/�Zi�Uf���CCH�2-�:f��U�kh�SS2�����F���`��icm1��Úʗ�ZȀ��nEb�(T�F;ٲ�sJ��V��sI������7)�6��w�x�������1�>+xJsyv
)�܉jM<.yF�ϩ60��dr�P�Mꆲ �@?G!�����*�1������8�/�G�ŀ�j|�=�rj5r�+�����{ˆ(��
����}y����f��Ꝟ��Oeκ�k�M�΅�3��z�y#�����z-���>(5>7����SF���ucw���u��zY��k+̼�6UCih��]��)�G�ET���I�.u���6=+U\+i2}~���{V9`>"��;�~�x�h}Ų��ı�2\a12�����L[!�ʵ�?�)��i�]�׺��fnM���R�oB�`�;,G�qw�&Z&��[�xg��1N�ǳ���?�}[�G�򕦹�)�P�1n�巪���{cz��ck��IKX~ɼQ]�u�}n�td���U�Ύc\�M���s�{�ݭ��`��r�ŧ�7�����$����YE�9�~��[���}W�����+�EN�� xV��K���zJ�5��3��frW��AOV��-�C�٨!�u��q�4��.k��am�(S#c]DJ��W5ih�V����"�j��Ӹ�Iށ��#v��A�s�q˨I�ٕr;ڣ'(��ߡ���!�~������5�au6�����n��e9Fc�K%��"<]H��jM��j���]�p�:x��9���m�*�v&�����{���i0�,N��-w��+V\ٗVjM�=2�L�w_7c&k�gsc,��Z�ٝGPF�ؿoFǦX��Y�K���[]��N���Ώ�N��s�e�r�C-u�\ɬܪ����)�M���#������n�p�DL��\�'���m����i�y6zz�ל���X�B�^���lo9M���X�'���U��7�d\��1�y�R��`|0i�ot_2���1t�{6�]��Z�Z�Wgb�h�恦�ri.�M)ΐT������ݷi�R܁YUў@Oɍ��Ɩ����T�{6�y�ϸ�)�t�@O�r��T���Lh�V�;\��� /��+pO:�[x�5p'��@�r�|��T��L�/.յ!p�|6~n�¡Y��`jź�[����n��
��zު�'�ˎs�J���kZ
�i<�P�\�1�PZ�"WN��on�OI�8|�;M��%�}}9��댾h+���ov�}}4�-Ҿ���f�no��i�6O�+�d9G1�ǧb�<�sSb��ˆ����i����V.`w�e^;��:�Jwҳ�8�������Zև��6����հ���R �󍷴�-�אzJ�%EεQ|�-����a:
�ܤ�%��c�/��O��sJ�{>;�Ѯ��P~���D��W	.�#��:㶏W�>|K�p�q���w��W�ݷ/;��mY��Ƶ,*�D�"�y����c2�ˮ�EP^��V*WR����d�򻧰�eXӠMvS�Y�m�ڇ#��Z��4Y�o/P���IWg�ۧkwWW>p��W�D��ދ޽�j��c��g�7�WA?ORt�*����Q	�s�~���}��.��Uq�y4�F�<Ә�LS=â{:�=`�nH��\��b���c���o�:X��Jw�c�k�r��/R쥋�b۩��K��+2ul:��1�k���,.̸����.���<�h�q3�4�h�l6��(D]�Ź��WP�<(��g�`����I���n�t�
���O��'��89��J�5�
��n�LpȂ�� �zU�� C���Jy�/Mgx9;6o;֝��LK}�t�+��µ�\��.�sf���{��n:�$g=��ݾ�}���s����ܽ��]k}c'���%Bƥ#�-^�7�Z���E/
�l�Q)Sw��\6i��?Ia�D��2_��Z�=E_-��h^:|�bz�j�u^����l_���S���}K$�����y��cV��*�CYą����Ը�Ok�����ok)Z{(�dl�h�Ƨ�&��RN�r���Kng|�I~���S<z�A���Zuz����=o����M茬�X��'�J�yr�N�Fxԓvv���b�(X�>��+��F���X[*oN�w?�U��A�ޣ����;�N-��|��&��=5�S_A~ٙ�䫓5:��"�l+Xfơ�3gsM���z��Y��;[o��~T&��:�W���ܳ�o����˚���'g�;��ci���oi*��
�~T'R�{�:��A����7�߱Ш��TE�U��.��Ѹ<�_�e|�����VXP�u��u�<���XV�2��ި�3.|�Z���ͤ��n�I�NM�MUf�SuO.��mp!)��c�]��֎�[�f\N`�+�d'[m_1',W���nQwkj%5�?��.̮ݦ��';h�	��\ݮ��{��P�S�4u��B�v"~�� ��'?W%�tj�1�r���9�]����G*�B-��W0��9�up�S7�*��&8\��3�*��%;s�}q.�ݩ>L��d{�\���-�й1;�j_�[���$N�$���۩�zg����(�LS�D����/�	��P�����ƻ)�i+��(�Լ0�rc����ƚ�y[.�1\��޽|7�y]��	�(��+#����*+6�z�����l�M8���r+ i�6'p�8��,�*�X���%ŷ�H��YZ��;���*gk:����L7ˢ%�����������4�2�Pm�wgט�ޙ�X�^�p�Hڭi��#^핃}8�F���`�KS�.�vL9ί1T^=�|b�	S{�'E��5+���R���8��L�b���6�
죊�ޫ�y�j|[�b�U�'�WasR3��Ƿ�d7����gU±s�3�Y��g�3 [��ɩ��}��-�|������ا��q�ꆯ������fWÍ�9_��{�:�0�1ۼ��,�(_lc�c\�.l5��s}��K*�ۥ4j�U�n��w����b�<���D�r�:�_�����㷴z9�,��U���K�7��FA�/xԨ1;�T_%Im�p�=ۄa#��}5��AR".��n�ڋw��hX�Q��Q���U�X�s��ޛ�7�w�z�[T�#�#3iԮ1�����w��V!)	W�.d%��#kb�ȖaHU�%83 �՜���)ѝ�W�*��Le(�Ɔ�w7��R��7�H�oJ�Y�@�ɀ�Ct�c�B����4���4�[����[��I�e�o��%��9�e�}�q��KXu�8T&��?����H�f��]�Z~aKl�ӻ;J�a=���K+4��Z��TF&X�㳠č9P�b�]�\�4u0~�W��guw8�V5��m�7A֦�;���n��#�Hm���R]���rer�-�:T V볤�i�ľj�r�\7j������Z����+����̳ip�z��H���mA�]m۵ǀ�wZOG��B8���h�@빨��봺9#U�v_t�W'���g�Tդ��f�1R+s�R�s�G5�v�-
�;#�����j�����csS��˜ �:�m���ݶO>��Z�~��{�羀�#�À�(�ҵ��QkVF�dM�r��)�w��Y��\�n� ���̇vq4�����u���t�m^iD�w4s��Rv�p@��)������|x�M��35���ѵ:Mf_c��ч��z \&ۗ�tcu�e��kiɷ������%[Z�H�e�{\�%X��(� �I�V�'�v^4��0`�YC.:5�@�nw;�M�����gn�#C�ˆ�<�0��e�$�f�:��J��i��&Zi��ħ����H���.P*hZ݀v�m����WL����[7.���fZ�6��w�Aț�[]|M�;���V ���Ҷ�\
�.�bD�"�|y�t���z�B�l�;f�=J��W��-i[�t�*H�lWC �:�M���k2(8�Znw,��{Xu�1U�X�f��+N���G\{��e�6��j�Ӓo�.QEY�J�e���ˣ������t�6�B1Ӆ:q�@#�͏�.-˂����u�Yg]�Z����?��*� %�������ߙ�{w|�L���ҭ�	�\��.��EX,V�����xb��6��4�fͬ�Q<�H�!�Sk1�"�w��h���"��t���inڅo:}m�Ta:o�@��V)"��Uޣ���;{��ļ��aF��9q���jr|��.W��i�]`��Z��8@mn�m+x�����8<A�ޝW���r�F��R*s=X@��o!ok�ɭ׬˚I��,�m�`������ ���x�{yY�p�l�*���b�U!�4Ѥ�8��B��x��ݡh�!PV,a&�Vw'�[A��10�n��mJ�������L�H<����8N�k1毂ܡ�6��]k�����^�Jsf�}�1[�oZ]�ո��:%y�@X�K*�	}X0T�P�[1d\���]8�+S ёWf"r˛K'OP�`[jZs5X֡D��K2��q��NN�dq�.���SP¸�rj��c��N���EǤ��!:c+�A5Q�ې�m[�:޶�U̷&��OU��P��kZ�4F��52�vi7`��ӡRWPρ�F�DT7�;�y��bC�E�¤����/q���*"�y稜��Gt�$UD�P�E(�y��G�TJ���8Q|�9#��eI[���纺��NT�d���P������H�B���K�8�!4
*��("3=�x��H��H�f�F�rց�y\>yp���R�0�\�)j�Ҳ5�DESfIl�,JдR�.����KB���fE
E�c��LTJܐ*9�%��;����<nFD��Ew7���X^��(�M�(L�OW7D�M]�Fwt��CsȽ"������l��r�+�Ju��;�!ȅ3%� �ܯ#�4L+��Y�Y�]'��42J�e*yz�I�]����n�S���ӐEGS��xy��w'�01UU�D�[ww��3Q=��$�ʣ2�h\��PJ�
LS
Į �b�IZ.�pTB�y���)�I8a�A%��ӹt:�EEwy�׏P��\�y�C.Iau�Y��뎴Ewd�X�V��*��U�����̌W�<�̫�v���(���sk_�ݜ͔�;,���W,���.��I+g�����mACdK��Ks����O�n�ʉ��7/8�ױ[�|�6)��+OP�b��6������	�J���n5��q�N����U�Kh�E!��hΣg2����B_û.��_kj%5u;4sqk�݊E@up����z�q[�yVnk1�5�{U�}��^��Y�Ħx��<F2���b��6ü&
ޣKj-��&�=ێ+)*9I:v�Q9m�9j�g%��t_(DLU��_@O1�`��̣��e.^ͮ�}�<�ϩ(I=z���I��Fd�_'��r�h���sZ6{J]�y��מ0�����cQ�'�@��_ؔ�v�T����n�¡Y��Yk(㽳�z�
c���ZY��^5�9�)i�x�\46_vu:�S��nS4�c�z�k�OrXO�3�^�s��k�c9�tjl\����Ҫc�5�̚�v'�Ww%J��ʂ�u˹��Ug��s���O홮�U���.����8pb;�K��k���Y�ÞI"/{�]4
.U�_*3"�*�wX�v��t/=�����S~�_ޏ�9�x�q�F�5U�<��Lz�
Ӧ�l��A{���ҕ���-���s�OOv�Ud�&���ȴ5(-�v�mv���_cj%9�7��x�-�o��-'�7������ʹ�՛��:mՍ�L�j%A�֫�䐞�ȭ�)�(�����j����4�:E��ٳ�̮{�&|?nu���t�RB��g!߫���b�$���ig8{��mA��PKDrȲy�{�N@οN%���U�2�ۗ���~Z:b��G&���q�1ܥ��1�lm%��,��Gv�Jb�f>���\��j:�w2�B���"k���������X��V�+B�1�~�V���{�:��K�ɚ�=�L	�2���C�A���:��U�Oԥ�Wm|al�0+9�]��պ}��>�Sd~����T�>����N@�Ɖ��	[�^qyQ7��&q<��`Yx\E���f���LU6���WN°'�뢵��ZP3¥/���:����&hW�V���=`�qW2��n�¢7�8b�:�<��ZT4�7��S�K������7�PL����[q��O�Is�[��;�Ά�v����w�;I��e�s��ݾ�.<�sN���8?|b���#?v�ʩ�O:
�66��p�R��;^3���d����� Jg7*>���xn�0kwKN9�.�C����;�m.�ZvPS/��_Bcr��ʃ��-��ʎ:�_8�M�����9�]]֊@#��-��yp�N�Gih��k8�\|�~8��<��t�ڹ�5�N�v�#�UI={�|ڞ�k�c�7%qh�o~[�5�kս�ߊm��Z�VN�m	��5V8��S�or��t����A�+��z�a��[���]�TY|��[I�t�cYp�k���g�#VݝuN��mr�R/�h�U��s�%���9�3�r��i󿸦�6������Zf�F�]��Y��a�C�1����~	p���h�og��s�]�{b,�YLwO0��x�F7-�q�W�F$��G>�������kΟ�,�=R��˯h��KT�3\%Wiͨ/8�]VtP`��û�u��98m�D�-��-ǒZ��=�T�>�����R�7�ws]l�-E,[�M;
���!+�;I�au�c�*>	���ި:�f�{x6^�nq���8�c��E�"i֦N��f������A��y4���eX���%\n�o��e�n�5�l\ي���5L7�5�[�4sw�؟�J<.
�	芘�z�{g�j�@?�s��Y���$����8v��<��:���&t�����g7a���K��ϼ�~��Z]�V�����VުP�SN�V�N��2�LoZ�d��ME�؛�^�/z����[��,~�N��A�9	U"�Y��Z�N�VvUL=*
n�u�`LktV��E.�+�S����k4�Y��kU����aH�ƺCB�:a��j�汷QvW��[�Qy9���R��/�g(��\o(�-���\.!�����J�����cd�>��27z�dG��]��.���C<�/mt��N{�c=���:=�5oa����<��=�A/w�▛�aXqM#|qG+:�.!&�C��Uf7]�����D#���ub㭰��0��^�M�T8����oc��7�w@�X�.�#	{4��uN�e<K�c�n�N���Z�A0���];@����M_m�g_-��q�����;$��ɝX�)_I�uk��������k���:�B�R�x7-��jq���n瑾w6کPkZ�8���e_ڥPƲ���}�x������fu{����F3U�|��yPZ�T\�1Q|�B�L'ΫkyH>�n�*͕�	\ֽ�{��oiMr��am��ٖ��q�{�m�;Xy.�-��-����j�������U�6��3_t�Q����k��SҨj�Z����|�F=|�_�GLB��)�\7���LS�i�eX��(����6���lv�j���.�S�x�ֺ���s�pԇ@�FLyoQz���q�u�<}��5ܾzR�ya�e�qYP�]p_S��3���t$$ֵ����A�}���k�/��^tX�+�"�9;o�[�f���#��r!4�j�z+���������9k�Kj�:�韱c��4��J��cb��'e̕��}e];�+c�뢷6��m��}�{7P>����6见�,;��8����7�`o�.�j�a�@#G[���\��@nV+f�:��&����l�9�jR�����[���D�C\��p��֙��XF�|5vI)V,�L����7gm�x��齶cȌ$��:����.�����:�����>0��wQ��r4=�ߑ%,�?0�o�����+ד�yˍ�r���7m��p�׵���Iy�_�����X�뭩3�z��7�Qs�V�+��Q���q��6��7�e��@�s����jR�pk���[�ڪ�.�!{h.�ǧ����C�U�[�paZ���V;����2��x�}÷#m�w������5X�w��{�&7�N�c���w=��5���
{�����%F��D�	��Uz��� �QiN�ָ�J�)꿴���wd;{P��_���r�/L��Hמ8EMs��?�y��B�?B�=I>wZW�8{��FӦ��:x��n�c��ÝmLv?�tnT���U����7;��4�1��\b�d�T�Ң�
�biN�k�+���y,*�	eJb�g�Ϯ��v��x��C���������X��FOR�v������3��w��Ʒ>���lv%iB���k��̷Ժ�����n4�W�-���Zw�9��֖n�]�������( ����q*��9y'p�%�Mč�����:�9S�p�5,�*�.�s$z3��n��ζ,��n�m����'���y��U�H�)���0L���Q{�%�[|��M4�Sy
�݊E��]�al��[���$-�/'�ƽǜ�;�Ƙͅ��.��
���Lp�/z�-�������Z��N|�{k�0��rs���sК�z��R��	����n���5f��;Z�	{�o�)�x.V}�O�������v��Z{��Z�b��WP{��7W����ʋ8�7�%M�)�¾�����WR����R��*��Z7�u����
<�h�[S�����3��f��C:O�ggU�7�^�~�7�5jm��q�5Y�.ڣ�8��joX��z's��E\-y<�sSb������C�rW��m���*@^�~�Vak�w)u��̗�Yj��vuVZM��SM}����u�CJ��A��i�
۳Y��6Xe��{��i�y��j����g����ȼ`�9]��iK&���z��sH�;��b���T�Z��ȺXʐ�3 ՟�����;���I�S�1�F�B�f�D�fp���z
���Tn4$��s�%E�b'ZZ�y�M��B��i�5�{�=��5��֛�o��W����4R��fj�l�gv9�,+y��Q;�d_%K(���;�-e�c���j�ˉȵ9N�Pn9�v��q��B:67��s?�Vg5��}���y9^�2"���~����ƾ�ݯ1��eX�S�Ԫ'�9�g�}<f[�+�|R̚G���▴���{���
��1N���aTk+�	LEt�J��c��Hga���w}W"F�N�3����i�;JG��ut	.x�[�/F�ךu�qI�^����j�_�VRLmD7���͕q��v��9��0��=X����j����A�IWƷj-5�g�X��ⲾԬ��bg��$v���<�`ާ��M���t^�4���[�?b�g�:�AȎ��t6M�)%�VJ�.�AƞS���5��+r���җ��O���{��ʞ�N ]0��>R]�q�|-Sh9���b�y���t�q)��붣�\c.���a7]*u�u�t�Ԛ�}�ue/M�l�a#�P۷���:�[��N벵�[���O<f���]�-���w�.��i�A�{��z%�^��;�*����\�Apȇ�L���Ǟ��w��˙ai���2�=�}�M��	_���T=�:}|�ѥ�7��*#�<O�q�%G��5�늶�Εd��Y��ڛ͢=�o��b��;�#b�}C}9�S���~�6����G�TO���xv4�j@��9z����''wT������DOs�%�w���7^�"�������v�dG�8<��+.��V���Ж�F.3�n$�'�"��&����L�>ȭ������7���7+ެ�����Emaݦw����Gexu��c7پ�Y�%I	N�Ck���w�۸~<���B��Z$`}�ϕ�=��=��砰��޶8Z�W�r�=�C5_@<zn�ܠu}�N�+<r�8�*����<}�uǱ�Sg7�<{��z�Lq�(�@ 6G��y� C&���^v�P{	y<��>�F�S�W��ٌ��_3��0�W�܋�z�������y�(W�}��f:�-=艉����Q���� �ZsS�k�*��\�1�}��N{�����~��{2���QWS��m�R\)�TTy�^�[ZX�y���QT�b�����^{�,��d笂� ��wA�q�i�j^�ʘXF�:�]_��s�#��\�L���J������I�rk;}��]Y�J���ͷ:�RwX���ف�knu�38��M�	9���bHVd
���q'���L'QH��}^ӛ>�;��|�yu�ygb��M:}O*]�&Ŷ�s��0ϕV �<�����$�Q�����b~��hޗ�݈��^Up�1n�b��sΪ�C3f���<������Bd�;2�z��c�r�vz�J�4�ϑs;���m#�mi�>�|�����+���3��y���s��ǰ\�5����;	���6��M��/�y;��/w|���t����#3q�,z��̏g��E�'<�����=�Q�q�̽'f=��EdI������n�?K�2��Z}d�7���Ω`/�^{c��=\S��,W2u�TL	�U�ev�������>�IH���1�5��:����~�5߼H�nS�z���_k�w��Wߒ�l2?1���/�]��.	�7^,����7�ک��@�����r��xu@_f{��+���P5�>�|+�v�Z
����\2�JzKzn���Wp�&uϬ6g���c�>�_w��nӵ�EϢ��'��7#��|s�/���/Ã�U���yl�*�����KDF}y�Ǧ�Ȋ	�ѱ��8�}�>�^���օ�n����=����2��8�-ug7]�ta���*a��E3�s.�Ŗu��r�]���4`�]�8�����:�}������!��5��q9Q�7Z�}:�u�S;�lX.��EYZ�Af�v�\��S�F�*�>i�.�uj���[�C:YP���"T��${���z����닝7�'���m�+�ț@��2���	*vo
� �Q�SaTcv���k����v�}�H�W�u#��-�ۮoW,�dB��X(Tи���zEI�V�1/��cpY���WG�o�o.qY�Y�Mo�S:��Ь�:�V�ۮ�]W8գ�h�!f��L�q��8f���1�%��.P뇬�}����yE�[�ޮ[|��.[ѝ}����Tq�0�H���~�ɽ�
���V��+��a5y@F�W��h��:/��6v@��u��;�5��"�����������v����)
��q�}�&�N}���ᆍ+������N(rеr-����f`݃5
�R��Lr�B@Fٷ{vy˥�GF<�-�d�ɦ&.�����Z%
�{�24�v�e6%v�ˤ�Rfpk�Yv�veYU�����C�;ۻ!��M�:���;��[��C��S��x�'2��H̢Msd�fX�m����E�:����U�����zk�=�K���}f���*�
����n�/k�l�Kh�J��wMR鉴%(��sC�`�k�mgW0C��a����]]ږ]�f��启NK$�״��l�h���%�>CIlL�3�X3�[¯]i�!���U������%��$m�`T�B63@�р<���T��¦^VhCp��,P��D���8���vT9G&*��+�y���h���c�*5=k�?���w����lfPO\����v�ߚ�~�Q.�w�J�G"��7�.>]����s8���.A��u��4f+�~�� 5J���),�l�ٮԨk��N�:���7��������� k�T���hU^.*q�Ƹ�P�. ګ���k{�S����i���ș�7)���;����e2�'ea�W;Y��Ÿ�e�Y�O�9k�j�n��(P��ƺ�T)�O��O�cha�1_f㚒�!�0ա��ѾE���oU�t�j'}ֺ.��p��/�����xs�ʵr���L�6����\[�!f���d7�Q�ͮ�����t�z���]��"}z�#�h�̕0NU��Dz���T�N��Q��&j7m�{*m�6���n<3�����g4�ҷ���!څ\��ཧr��A-���I�K��hv_vȞ��E���c�^��T�Jָ&�HL\3l<�I�K<O#�e����C��/�v�$�sE;�魋M���Д{�'G6���m2x{��1��
�(4��.j�e�c:sf�v����c�˶7I�1�vlka����
k�.瓻�G�#���'(�.z������xx��^l/\xM$��4�*G��,��۷<��t�7e�hsJ�ws	(DZ�륛�����uwy���us�G�Ȯ��3wsծF�G�����_*�檏#��k���)�Q�<���:U��WsNF&�[s\2��2�nd]<�
/M�R�U�		��s��MfTjHn��3��z�iW�2"�g�t���/#%�ܩP�t�>2=5�dw<�u��R���$�#�笃H,�����:fa�H�sܥqO5�t�������Twp�]�7wS�Θ���$ʊY�DOR��3�)�2O<�9�KC��	�ª:"K��R��^#�]۞NUܖA"�̯P����u"�j�8Qx�&j�52�%T]0��Mq<UR�(��L����9�\�2By܏9�锞��N\*y����%҅!;D'�s-i����f*IQ"�h���ĲC�U�y�m��-9��bX�u5u����ʼ�,��T�Bu�J�zZüT��Ӛ�y���F�m�9����e�PJugh�ʴ�گ� M�Q2����]3.�����3Y2,|b���i
	~�w<?�����/��9��=���i�}H%��@�.n�do��>��_���,���ފ��y�(6^��\߭ |��z�}�����~��H�;v[{�+�h�t���t{�Y�= s��Ш�[(��>rY	�v����/}�����~���\�V2�-�xc��yg�"ba��&3�KZ}~��١�	>U¦�V_F�w���5�wux���5���嚎PG�&@^5��>�a�Z;�����65g���E=R�$�־��>+�a�\{����Y�-��&��ai���T_���9���*��4�gťg�j0����Gt��/M�~�*�|�#��^��'a�&�|8/nZ�ղ^?��HȕC�;S�^����#�>�#^Ϩ�%,stj3y׍�_��ǜ���t@}D��z�_gٕ�������L�Oq뉺�Y���d������=,{����·�=�gM��r+�H������ޡ���p��bV��۝�~���K�l֛�u�f�*�_�vW������$蜩�b]5�W�]p�N�c�}�9ܼ[���jP�yQ�k)m|)�[�����ubdK� )�.4��ˬ��&���*vJj�#��#���Yc��r�L!%Ջ��h˵��7�AY:P��{���ļ�Էg[j��'�x���f�U��� �d�*!W�Ԭگ��S���pgא+���y��.ty���,�z����dam-}+��[H�G�2�Ǖ����и}��\,��n"e���TemÍ��W�Y�r7��յ>���ϡ�]�g��~&�=��=ڽp��<W�<��9d��e�ܣڑ������������KK5TW��7άn7>��K�zv�#Q�b�y�Q�A`5�i���ץ������Z�7�)<υ��/��� �:����:=�>G�^O����T)��I���_u��{_Pf; �>���uL	��G���^F�G�νŌ����{[�ւ��מ��<®=�w�ޯ*a���¸�RH{bk�)�D���>}pQ���#^/`�ٳ5��%�{h�z=���Ϸ�>��#{���/��:P#�2pw���g�>��x���#ׇ�-F5���o�D��v�Q��Izg����<*�~�%�����{�=�ٯvz<�kRGeU`ūg7�=C�T�9���t����n�=]o�>>��Q����e�V꜔O`��<&�~�(:ח������q��&0S�):���7���rR7�o�y!R�P����Z��ٸ��l\g
[g2%I����G ���I) �:o�]|��F�)>����9l0��6
���2�hT[˱�C�[ �hv��ei��A5�\/i�Ss4�_��VR��?l�gFO��B2��s~�Y��/�_�n_�@x�T��b�Y෱s���=�%C�&�^W�����5�|=؍1��\�ߪ������ׇ`�z����N����^�����C�����kNM|���s���I>�3ǯ6w�����j�>�~��� �D]o�|n%�
��\�u����7�I���{�ފ�i3{Q��w�����9����_{�w��Q�qޒ��ÿD챋՚��霾X�}����>�ӵ����z��s�(�W>�~�����ᯑ0��`��}bZ彔y^d�T�d֟^O�
�o�o����L{k�{��n<��)�����fL�jY�v������1��>�E�^�ɭ,\d���N��4��;aϼH�b�x�[���O�-z)�Ӣ���kJ��
4��� !ݏ	��S�:�3�0��ta7z*�:����E������^g�s���2=����,wM�� +�^S/"�O=�U��8�A��Y#vI�S�3�ՙ�
��h
{��W�Sα���O���J7�^&;2�Ӓ�_�D��>Uc���#��y5j=5�F�W\�1&bWj��;1�6��s�)��ʦeI�ul3:�Y�!L�XUȜ��{h�YujL�1�H�6��n��a�16��}�Y^����W�+��;�;}���s]HSUA�� L}9�1����nkz�jf��љ�w����ѓ����[�Ty3�l���=�7ӣޯW�B����@l���Yc���E�1:Z|{蜪rW���8�Q	⨔�]�������tߩ��T������$���
G�ba�U �eN�����T{�W��b��*r��	y��{�W������>��̂*�3hdA-���^���14��� �×�P�s�x;��=Y"�UE��&iW�>�>��W��~���E?	@�L�*�a�	�};Gt�揺�ju��=��8�'�}{{�p���>��ϊ� S��"�9<MD��3a��ͨ]K;G��0��;;mB��ɰ��/�����5�z=�@y�%��{>(�H�1���^�&��@b�"��ŝ_���r��*����sO��=��_�ۻ���c8�>��G�������9���w������ɴHB�}9_���գ��N��q���7�u0*�dx{��^tx��E����Ѐ�ӴF�p������[��Q��VU�u^m^\ ���-@��HEj꟔���(���fTY;�c|o��\0���]j*d�����5��B��7�����$��gf��Ϣ����j�'I�_Q��+ػ6BgnU�u�[��k_TH�Vs؞H�=�9�F�y�Oi�-;1T}��Mi\��ux�^�#ɀb��l����}値B�2}R|��EE|�Na���>슨Xk쭨��Ӿ7����[#��}�0=z�twjr�|����d��>��ï��C�yh�.3$�PKvn"��λ��z��y�0}�ܝ#�����Oz!ڸ�{�1{����*~>]~��^�+��݃�+.�h�_�N�����alߙ�N��s ]�F{�#�o���DK�G�4�����2���i_:�q|�=ݘ�������;y�:��O��'H�:��x�������H��O��>fz�����"yd�{B���G���B9���n��n��zf���g�r	l�o���m�Գ��~v¿ip��̓�7�pMv_;8��CH�^}�$eC��!������7=s0�EңW�aȂZ>��\%K���J��[ns�x�5�&��h{�}~��N��
~�#�P�h��x�Z���}^�^�����J٘��W\\�[=������Q����/�=O� �i���z� �3�d[�<N�L��L=���݋o:+i�h[�?���{�V*5��=O����l�\�� !WwDs=mvN<�t�kv&�N��Mvz�v�\�*�Wz�X��`��l��:�	�>�~�o:�e��hI��.!��WV�i̡��:R��0�.�c���&�I<�d�mF������#	�3�T�5�Tz��W~8}�Ǚ�V����?3�x�[lp3����z�у}UᗛD*�zdTo�|m)zm�5����D{·��KʏB��B>���z�L���ǚ��F��$��(���O����:�s
��=&�\�2���'4<*�;����^�������[>�}k�
(؎����zW~���ZV~`�'��c(XF���s>��s��P=�z�ȟ)#{�˱C��86;�x�A-�ʇ���P�6�KB��RǺ�������^�������{<Nǎ2�Ǖ�ފ�,��ne��,]UX�=2/ٞ���:g-u�G{������@o��Ln?S'��g�}넍�����G���!i�}��g)ש���y���_�/�7�Zc�J�*����{�cq�_�ǟQ�Zv�>�u\]mA�Q�o�-	@�Q�F�(���s�,^�S�ͩA��>>�ё�:�>���N�F櫧*��r�4�N�:���Ʒ�e%��:7�o�&���l&�|��=q�^G�W�Q(����^��w	J��2k��ؐ�N�of�-����� ^	|�����퍐i���Q�˟�e
�oษw;z�_��wѧK���l.n�v�ˠv�v[O{6A�4[��Y����7����b�
;|�a��:��m�ݪ�I7�r]9d���+�j�U�]{���}ǟ�@k��t�W�B����;��ׄLSt��+��z�!�q��.����ҽ����qq��n1��wg�����U@*�% `H�W��a�L�ʖmz�O���e_�z0�^{�
)�Wn�i�zPL������q�UzK�@Z_X�]D�b}y�^ly��P���B�~6��{"�ԯ�|��zt;�e���$�;fy+���&O~��#���J��!#�88����FXۆ�q��R�Lg�}��2g93�^���
�������)�ĺ�}�������&��U����n��6�|�(�J`��DĶ��1�j������;7���� ��ġD�>���ו�ag���i��u'W�\�ݾ�HV%�������o�y�~yv<0�E}�Qˈ�c����̨{��|�ب�[�~Y�H���)�L�Ψ����;����w	�{n����5ޒ�\�N��t�X8*��.����Ӎk���E�:��.r�o�S*NF�`c�_��q%����{��*��Ε�aʵO���W�>���V�A:r败�@����!K���e�/3'wǱ��8��8W4�{y������Q����&q�8t�k�.��\{x�[�R�ps�F����.jc��X:Ѧ���������1+m�r\��q���Qed��z%�����L�b(�<������s�4���劲m�ƣ�a��vH�X��5�e������
]��C�^��~�&�a{��#W��g�t��Փ��;�]��Dv<�S���b0~��|??�<>����{ꡏ���$][�3꾟;ۚγ�kA����[.~F��QJ�@pu�s}�b�&u�em�'�B�rs=�F��Oy�����Ǿ��q�9�;�T{ט����d����鿢j޿t���O��^�w���z���u�6r_�ǲ8���|X�Q��~-իc>S�Y�@00��ޝ��*߼Ŭ�q��}�=�V�{��}���7��D?SgW�x�/�����x_�r�,�O��(�I�nwux��9�O�*@ó"ϧ�N=�d�o��~��g�
�������Pʽ"h�����Fн1��7������LL%U��՞3s__.䳍4J����{��R^o��Y�q��P�M�`�,��U�L/W�H����:Oˎ4��v����o�Kx�S������C��V�e0o�z��]��%Q/�&�1����z���zn�:.r�\�A�Z�0�wR�Pӗ�]X�?�1�>�/c�rPȜ�q㭽0���EB"�@�� :Y��Qўޖ��%���&��Q�|h�:��P��-�w`�GS��v��j�b���7x���n������5�p|�{� T{�(��9<MD��3a��Cu��5W(�z~/�l�s-�k�31���1����@i�5�^�f��t��yw��(ԙ�t퇘9�\sÞ{��4xg�kB��wƳe�36�_��ٗȥ���g�wq퀹ǻ�ϽُG8�g�����NIC*'+��������?����U�{p&�� PҥB�Q��6�[��"<XD�g����~���3�h����Mi�΀�dj��Ms-�&W���wc@��#2��)�h�{)	xTT+�n$�>쪅������N��}�^�[���n�����wB6���M����ϗ��{�Hh�-�Y(����({q�}s(�^T�����C3�^�>e�mB�wq�߭��t��ˍ	{p��N���%gzR�u7O���띷�o���`>��k�p�'�|-����o��z��<S/�{%�V�WZ�X��޴�5|�9*x����'ƾ����0&*W���	�mԏ\7�C،���C��+�~���� �����n�J ��n���m��x�Q'H�E�5�J)�ڒ��[`�����8�N)���f���hM��V`��P� A��U!�e�P-�6�,������v����/s;�oxn5�-�ϗ=X�2�N(�wA��:2�])�A;���Ez�:�˒�F�G�V�=��a�l��9\EW���D��7�h�]��,n=�
�Y@ww�ny���״{�#�����1�G�Y��|nz�f��T`/J���}���O��W��7�yi��F�7v�P��:h��(��X*"�t@��b�@h� /��Xw5ځ�.�M���\�����2����L?y*��:W�>[,�z� �ʈ���&�PZz�W�V��J*����3c�7ѝDR=�~�+�t�^o£��W~8},y������7yw�]C�,Yy�΋̔X-��d�ds����Y�p�S���>ۘ����)N,�$�ɁJ<Uz3�}�XT0�_�M�L����O����d\�y>�Q�t��Ǯ� ��(K�o͢��et��پ��p��c��H��	VH|sgj�2�LU��M����ͼ��H��9�d��ӾqY�pپ�������Ν
�{ۘ(g��8+�'H�70��F{��{�vO�lU>�[��x���{J��j� *1߯����(���q����B���Y'N�L��3�AbLO��ث���5��.�gb�ҥ��3�Xf����-��/+6�JNNfEy�jWWrv��WNcUʇgsu�c��8�t�
x�_|8�Mr���^AKl���;��;G���%�9+��5p��>=�X[��w���Qc�v�ح�Aq�4.�������E3J��I���^��Gh���6wB���Q=�x�WV�tz�������kr�r������� ��n�bOl!���5Ӆq�ʘ�.U�4�u�X��v�)A tӋ��ޖx���0%X=ꕸ�̕��aOb4[�b��o�Ei�d�����˸��\� �w���1'OZ����Vi۫�t�I����A���e'�h/���7�9_)���L�R�k
��q<Ј����mH���2w�⩻�(R*��!5·�ky����|�Ѹa�[44~@[� �2t2['9�@%#��JP�oN�N)�X���hѹ��I��4�S��81/�fa퓯�ꝭ��&V(�Q��������Q�M`0H�0Wr�!3&�VA�����n�4vXGR����wR��!�N�t�����5	��������[5��1��e&�A���%�:�m��^��XAo�'Z:�7a��2���R��r���|���+!��u����U�tR�;��TĢ����KU��v�R�KfW8:�Mܷ�A����e�E_px��
�
�1%���M.����9��z��4���)��x��>�x�@�u�x7����։�m�7z�3YoV�s	dL+� ���3e摔��N�|F���_f��팻��M�����fݣ�4,�1�+y�J/���K7���8�`]ke`�gAq�媲Xy��LJh��jݺU�p�49J�ʗ��W�L�ۅ}k�r�`AU�#��V౽�c�j!���z���8%k\\�B���|�eJ�f�`���e9��	��p��h�`}yR��u���,��u[�	M����}H��]��e`�{��6�r�c��Hi���9?���mʷ��M�I��Xŗ;TDڢ��b�Y�M��Eʾ���u
�1��
�Pu�t!
Y)-�I�����Ql�g7w:�Y����5ix�a]�,��a8��w�_(�vl����d�=�6RYX�Z�"��RE��;j�h�UȒ�gY��R���S]@*7�TJ��69��Q&U��}f�^-�-�{6�Q�g>�M���:�I]���:�%�A��B��Xk3I�q�{\M=�i��/aC��U�R��L���6�����,�;��-���k`r���ZI��͓HOT���\[Y�°\�l����ˈ�SJ �,w�ۙf�<�軺4Y�7,��O�?��㚙�VX�]wىA
�2�(��V�l�Cu�̥E4�9UKP�%��+I!)j�L*��5�p�C���)T�����%���I�HRUZ��)�q�!B��P��t��9����E�2T��
šV�D�G �:8�p�]wP�*��MK��U���*�"	��,�i]
%�(�U.��ي�(�C#C3QKP5,:$����+y[�b*J]5��(㒡���J$�']u����Ң%O%���aC�VθGS�����%����KJՕVV!-2=�M�������L�#3T��D��S"�yċ� �XD�E$.�)`�%��#H������H|��%�$��f!IX���9�.���gT;���Z�@���������;�y]�T��2w��i�V!���N��5�w�/�����t/�;�#�F��n���g�����p����Q��~'�ӌ�(��)���۔t��]Q�����T�1dfNN�PVdz��L/�r9�����~����Z]���gΦJ+�ݕ�����V�YEa#Q>�]S�x��2�m.ː�#�Pv6|΃�x{X�K}����4�����CM�x�;��u�D���T�S~��|M�˸{w�s6�,��=�7�˽��I�ӣ����do�_����n!��b��d|��`	���noOT߻*��P)hJ�rU���Q{�Y���A�Z���z�^ܖS�CsD�l��*}~�3�;�{iȽ���!��8���^��(���\U�:��r=��s}��N�l{�^��7۽덮��K�:�
�}0P��-� �F��]/���n⯽k���J7��#��f���yuV�y��=�^'��I�;q10�D]"f������Zw!cn���#�J�0�E<���w����Y�6<�"����^L����:׳|J&��*���}q��b�����n�0��H�O!a��M�Bq��P"��s� �k��/5Zj��۪�i[���!wd1HV�#][�/w�z��q�宵o�]�I�r���O.ȵlg#M�[wmҘ��޶WR�N�݆��V�E�6Xj�]לM�R�����ڮ�z"*���1�V���C;AZ8����<,����Y���cK�&����\9a�̟L�=�����v<�d��@�Q&�2����d�]�����E�訬^d�lnV�G=��ﺐ�^v+�������c�;F���r�&X�3ax�G��^�G-^������J�﷧ș�θ~7�f_�|�TZ��U�}���G��s�n;�Q�C#��qw��;^��\�s�7	E�*����ٿ�e�)�ڗ�Z�~�d����������6tGW���hJ��l�>ä�IE��c0Ε�>�s����|:����m��\޻>��Kg�(����۝qF�2 ���pyݙ�/�ǭ �	��v��ߑ�k�.�ݬ�-����XN~�=����Z;�������<��1q�R7%�=3�c��:ϩ�l�����f��C��t����F����{�y����^q���>�9Dl�SQ%�SsP��W�QڼhWmOfj��{�9~�=��e�uT?�_������v>�I}=��a������r���ષw'6�޽�tt��
ޔ�Je���~��G����s�i~���#����ib� C3�lM��V+����k�X=�=%`B�磿�a�H��8��nY`�1�w�p
,�g-�7����n���=��Am,*��6$zM���^��9��8�$!5�|y�x���r���B��X��@P+ś���٣�+�t+��o%�3����:�r��c���Ǉi巶1�~��<Y�v[��|:}%����&&��Th������̇������+�����|�P�I�u(>�<=����7���3ِE�f� �z�&&���>�i�Z;�/k�����ڕ�o7[������Kc�樨�
���z�]�����ؙ��sk��}�;��z�׹F�9��������O¸\G���G���l�v(�D?ID��ɮ5u;j�(O��ۮ��;Ѫ��E��5����n���n�F�k^�Ð��x�7U��5��]lA�.v{ԵEZ�Q4�gGq4|�ևq��3Y����)c��������8��L�VfOcǕy=�L]����vQ���zH�9ӵ�����>����6���X׮�'x/LR�=ٞ����m���{V&�Q���Hl���<��qb�6kM��@w���t��1����]ޱ���ѻW�Hϗ��'<�_�Z.h��N�/�ET<5[P������<]�ʹ5��@�wX8b)���`.j���Y�hi	��i��ܷ0��f�r���N[�Q��3'k�AɃUw8�����*���ǉô�\�t�+�v���G��r���EIN�&a{mu�����йlO���T�r��c���M{'<}�����.�ͤ/0JL���U�;�|�bt�n��L�R������m�Ωy[T9<��r���D{����e�q��w�<��+������7�ܗ`�K�瀞����;�_�)�}t�r"_�ǳOz��~+�{'�/.����uB�{�5F�}�Տ����늦^��(6^���y���#>gC�z����}��P�8��f�Gt�7�\{!��v|�]�[^�D�Q8����������}y���v�� �إ�g�(z;����\s|�~���;�p��zfCwT���XT��B�T{{ƔgKJ;�G����=����ґ^�R��w"���y ����d��7z�z��X:�s/T�z��z
U�@�s:!�x�{��Uǫ���������dm�
��S�'a�q��y��-����p�>�&��_Q����ӊU><�&;�3��>�����%e ���}9x�팸՞��f�#�t�h�>(Ա��z�u+L��;���7f�n��E�����;��,����r�\�C�ry�?c)�M �#��A��L�V��u��^�Lј�V�L��k��i����i�&���7�R�E#z�������ݕ�+� i�4�n��w�3Ӟ���[�z�����y�p��sՉ��}�k�ˬgrM�@z��������2�v�f�Gb�"�9r��$�#�{	��L>Y[��O�I��:�.�=Uy�H�S����%fyA>�pzPwg��ڱ�(�+�%a�/���B��n�w��!�cG�ޟf]V�%3����[�ok�S�<�TZ��TGW��]�����7�:n|���X��n�>� �j&�[���ލ>��y+�9|�M�_��=�'b+ӍI�ꁦ���\B���k$����Myڌ>�sX�Q�y��a�K�emǯ'���g�o��ׯ��o�8�v��\$|�TW�)�CĎy ������(yvIMʜ��VMixN�c�{��9顷߯��F����l���Go޻�[���r���l=>�������_YD�n}8\U0&�X�����ۤ}��:�I��(��yi�^���=�tz;�y�؏e{��U��m�Y(�I�*o�G��aL�
�bc�Ԡ$�W.��Cެ�E�=�H��z�g��v���}�b�ڧP��!��:x� <��9Knו�+=��}�Y{��(�<�\{"�6r#}�=��0w����2!NQe�����)�sC�U����Z���+��I��{Ѕ������L�LZ�E��w:���ljN����:��]]���4��F�Wz�S�u�R� �i��Y_lI���=M�	E9|ldp�N�����OA(;���[�g�S�j�%<,:�uG`IDF��ռ/�:-����.>�4(�R�2|��\^%QZ�֑~��S;�8&"���!��"U���K�s�Q�d��]70Xuj�Qs�s �]/�ǵ����u��>��QW�1�v<A�:���M�9w,3ބ�Ȩ�T�Hh���1N{�F�JӰ��\E.��;��~��K��/,ɏA���L��tq�d	s�Q$6V��>���14�mg�v��ն����N�-ԅ���ڹ:/��~8|�yNK�����LOQ2����^V酸�<�sK��z�B��I����G�cd:�2Y����ŭ�s(�^���e��rڝ��+����*����x��{Q����ޟ"f�θ~7�f_�/UQϼ����=��p��(<E�^<���c�Oz"e�q;,e�c��������c�g#Kb�?o��x�RY7I��3�{��ѪB����:n>g�������;Le�MiW��Zms�ޜ�S�ׯ��O���88���:p�9ַA������wWqj�E=�:a,�nK��T�a�,lFL�� c��ǎQ{7f߮+�ɚLo5�~����֢H�Z'���Z����p���\\�5���
aA�'��*�d�{Z7n�a��}�7e,"ȧQ�ΫOr�dd%x�[渽�;nP��n.�TqN�;8z��.�of�����[���gx����T�H���^G��<:��v�g��F/��)�𞸪�㊥����ҹ�SȮ�X{)mύ��BVz��܇޿qȏs�3޹���4g���AdlL�C	H62�b�{���� z�@��|�]��ȗ�q��a[�L��{=�p�v��S�Y���o㟐χ<J<�);�����_�K��#�}�7^�S.���L�?+�`��q��{\����*���<���R���{Ez:�x��5���׮�Ar�7�Ǚ�}D*�����V:�y�ē���c��DW��Gt�5~�\<��+�Xό�\��ut���V.W�d>�Y�ٻ��Jgo=�sZp�g�W���c#ޔ\���V;�"�,� ���/l]"k}3�������ʔ9i<m������}q��ަ���U����d{נ;�fA�P5/�����I`�A\ɪ��ej�=�9G�[=��{M���Z���r=>�'n!R '�F?Id�����s5���Y��3c�o6�U�d֟i��J_���m��7���#�/\����p�?~[��1�L�e�3y�M�;}�<�R�t��(�;	*>��;=�wL�b�;*��O�r��aR�K\i�8v1��f�� ��v1�x9ֵ�MWTni�],�guh-�f�T�^�����Y��iE�>�g��j�%8J5��%���dz,�/,���ς�ͭ�w�k;��fq=_?fdy'T}(S��e��s�D�yd����S>�븟)6v#��/ND�3�;^�'t��tV��?���u�)F�s��߯�1��	w!U��FF���9tx׻*�\y�1}�=��v�v���{��5�c���n��k3��=�`>�V���u~����L���~��4t<��p�N鸉/�ET<5��z���w�U[�n�td�;2]DN�}�_��dk�����9�^���-墐��(����!ke�-�G�&�Cs�ա[��kƖc���kݴ��U��=>��K��Tų��^xn���![�>��5����3�h��@�����늦�z���)��}t�K����O�������d��c,+�f��EC�
�D�O}�{q��e����Q= w���G���F� �ͩ��?ZQ��/:1��Ԋeu�I�����z�;�>�q+�B��q.��9L�N�D�a^/`{#�}gJ�{=�^���_x��n�-{���AZw�$c~�dz�*�w�!�ۉ��U*1��l��O�*a��
�I����)��Y;0����g��0�!43�9�<��3���ԏmf�)�}c��D�� �	�}|i��+�F.���љ��gm^��˗=�B5�`��>\D;�jjKv��|����z8���7+ʻ�{3	T۾���̩d*QL�nコ��W���%���\KyI})�R�o��p�W�z|j��]X��N����>����A��Wy�q�gM
/����~�P�o�׮+���Tmp+"=���]��w�bӭs�Y�z�\ܟL��n`�:�DM9�;��wN|�^��o��g�W��-�I�7x��}&�;y}�{�x\�x���d�gĢ>+bn���Q�V��wǲ�6����n{�?h͵��ɳ�Q<gb}�&=��yNO�����jd��K���n����.�|:Mk�w�.��!�U���F_/��^�6��/���<���n�{� ������WmB��V���p�9}�LuH�h��R���g��(�� ԯ��/U����eء~z+Gx�7�-��]�m�O�k#����z��&ϳ�P�#6�M���5_���~'�YG#�2'M�:�T6�hU3��Z��������׿�ٔP1�\�B�/�kki �s�2�:D�,�g[��.�A���s�z������Ez;��Y#p��p�CۓZ]��3����I���U�ϛ�����f���9'�(ފ��xk����9���>�{�7��*a�y|���&�[�bv��ғO�`�p�k�q@J鑜��y�������5�l���	��|�,ޤ��olv��]��Ĭ�G��d����9_�OU��\m��v#�3�-�;�i)�l�vOq�^Ǒ���o����Լ�[��KK=�,k��0o��R���;�c�
��
�GG����G���U��~�>1�be<������>&�����MeE�
���Oz]�y^G�>���F�Ӫ=���Wh1�)��;K�Q�����˅�2�Z���z���j�������(���폙�{�#gkû~t	~�_������m�VM٬%�v$gs�-�A(-7]4(�ԁ���/�\i�Wn�i���"���D�3�^��m��vK\��3��k���ٸ�,:�T(��9��X\w~�~>Ī):�����3g\ŀ�g��վ��f���Ҳ#������[=s���&���a��2���
�m���k��gu<��PY3��=�O�9��
��� 3�Q;_su�+���U�u�W�Sbe�}��(ί3���u�cu����5�j_�WNG����*l�(�|}su��E5E{�y�[<�vn�Y��k�'C��	П^�,��@�/���^
!x�o"#�~��9�x��}Ъ����&u.�-���u=�اQ��͚�Cc�\�B�ܧ��i���u&.��^��4��:sm�%a�C���~��DHnA�YՕR�:�N��y�Ĳ�wn��ͥ`�f�5Q���m	�	�u�ͅ(��)͢e����;T��������}�z!��k]9�S��ʍ�5b]�}B�	�0.k.s9
�˕�����9٢�v��ɇ����`�3lV�{L���Y��ccy���Z�;ʰ����OjTNq�����KFDsY�Q�����V��y�C��,\4�G*4�D5샆{ >�j�wUе�a�Y����Ibr�8{�dӁ'��+]��5�V�L����\n��ا  ��-'܈#���^obqF��g��ԫ������wZ�w�.Ω��>f��A�y)���TNÙSJU�T��+�+9ܒ�ج��u��]�un�ι����$_N��ov)�TE&vK5�X�'fmur/0X�d�;0��M��J�[W,5f����:��lN�4�H�,�bD��G�!nq�������8�e_t��G�ݓx]�9�iK(_k�w �2�eN�n��b��=�y��I��7d�*=#&����[�'$��f�A
5Y��6�d��[2,8<z�`7�jӋ����mA�FT;/���[;r�n��Dc��=�ާoM'�;:�}��34�;���u���Vs�͊�+2�DccT�{��X��z���΀�����H����c�t�@h����]���[;�����@Z�^q���6.'�f,�mhc�Ww�u'�U��fq׏4��G�_Nd�R�Jt��lJEj��}v�/&`y�A���Et�/�sˢ��o+2�C�vQ�-=�5�����C �C7dɻ9������(U����ݩ�í͡E��cH@�1lX󥌷���M�1��ux�������ץ\ˢ-�Q�U���E����&�'��N��$j\�����y 38k32���E��:v�5b�.��K��[���W�V�3��!w���Z߹o�+��N�RR]�h�(��)�+��|��17ۮ�8fwmޅ%d)�d����@7_'O��V�&]n��9PU�0��. 
w[�d�[�/��񹫲�'7OVe+G��.-��������<����9N�	�K�B��EO�H0�����n��Na!:��{�h2SŦ�D�WQ��2�#�]ts��=,<�������d������kھ���w�s����ߒ	�j
dH�=q��7H�vvQ3e!5uĊ:a#5iv�����#g;a&�_h�j+�eSW�S��Vlğ'4��Ʒ��¦y[��1�`a�ʹq�s��0t˗�w���[0j��\����Z����E�a�#yQ����kt1��q�=٬�r�RU�5�P�Z�Z$�
�C-�K�WhO����ݖ�����D�5r�Tޑ�\U�E�M��Z�߉��5]i���m��a�҆]c�Nswf�\���c����5�Ԁ�(ʒ�DA	�IAR�n�N��4�j�^����-f$bd�R(��P��iZ�*e�ӑe��Eؖ�A$*��QNc�)KL�*,�����=�N&���T�"O���H�$���P�sRRj�C��us��#E����djb
V˥�����šY|�c��rDP�>\��!ȹ�(��S��Y	dif\��]��B�/�u�u�7�s�IXEL�����D{��KIkK(5+"-$з7ȵ2 �
�A3+�VDjb{�{��G���ui�e�r�̸QZ��D�Jah�\�iڢ:���:ej�#K!(��Ez���+��"����I�����])eBF/b�k6z�}�(�N}Zzu�c#b��ۋ�]O���/v���δ1���K=��9��g_)2�J�{x�K�ڼ�r��k�a�`�&��<�č�h�Ψ~>��[~�>,��#�y�s"�%��?��kp�;�ε~W��<�?L���Nφx�tnz{6X�ϵK��w���V��5�j���o�};�=��0�HgO��:�{l�GǧA�CK�5�vυi�r7�q���}��(�sYZ��]�Ϻ����]�㒨�}�x°w�x|�����&��q�;�Nr.(a��:��$�/%�t<��z5<����$?k�#��u��hvym�b�0JF�$�'�����w\+��s�uj��-�����ɟ2�u�O�S�o�o�}�u�{~�z������BP��$OM[���^w[ۻ��]�����>�j8
�������q������Je-�_�ujض����=���N:&ǐ�l�.�������Mׁ��˷�bQ�i��R��^�G��w �/yW�z\]�J>�^{(+2�P���+��]
.Z&��c��>�}��e﮿��_�����I���U�A��^��u����j�n��x�zK`�z�ba���Q��^++�4+�����Tem<�T��r�0�p,�ac���(u^-6�O��U33u�p�M_|�-���ϒ�8Z����EVM��zU#<L�W>�⥐Y����[}��.n�5I�����:���N@l4��
����ش���*s�Ws�+i���7�V�����%b�k��ýwu�W�z�2ǰ���<��m�@\���Q0�޶t�˘�Xm�oz���d�3��1�z�(gޥW�}��Y��=w?���e�Py��9�vb��uZ��}�&&)umҙ��j��'G{ʯ�{���3�^�AZH��#^@��I�ƌ���}:7l̈́;6H]n�Mf���(<=�vj��7�:ț�:�ϖݡ�Sq����:S���˒O�����w���6p>���ͦ8��%,z��2<r�˭Wn�7����l�J�ܱ�ު�7�ّ�s�o����G�Ή���q��? �7����J�M���
Oe���F��C�L��sB����������V=�#KA��}�rV�Q����lL�s�9����#��i�r<�_�YhP�����,�nK�������6wU{wє}�ꇝ=G����Ϛ�Y���^%�<Woޭ���1�墐���\f5�&j���j�w��p�g7E���=d���ڠ���w߫�}�2��ˎ�15�w @�7�3��,	�`o��_Y��?
�g*ƺL�A<�z�ƨ�}R�k�X�tN%��7�ܡu٫�_r��4��=�f�2
������K�o&����غ�jL�_	�}�V�o���W�7��΃�F�uה�k�C�������F�Uor�݁o��r�(��d	@��튦�z��n�gä�/�a�.�~��UFyU�TeZҷ؊�8sO�ϑ���6��e�l�(��޸�`O�<�'
���h~)���N2F|>��y�w������8=��w���n_�=��c�ĺ#��+�B�l�v�ۛ��b���~���������w�Hw�o�2=�L_���{_���������z�Ah������}W4���F~�����,���yd���A���4-ש#��u ^}��4W��w"�ޯ�!��T��]]5��f�=~�<H��}4(���	h��5�׽�dVz���ǜ�*ǽz u�F�W�5��^繋�����I���Zn&��IN{N�~9��L�6߅G{ʫ�|��Wy�0$�fx��U��{p쓗 $�>�|T���|U��g��ei���kò�5�'��R��M%��ͮ71��P������I(2U��8��j�6�;�������B��~j�/L�\w��>�6�w�U��p�A�{�gOG�Տd@yDQ�+ė�nv�{8k�踙]D�+�~���Z73��v��wN�;n� P��%�
�:��\!Y���/L�1�r)Z{�v�*�=-�FVZ�|��u�媝�ţ�tɐ�S�]�K+��W\YO4��:����Av�D�ZC��/8��C>�vo�_aΛ�Z�'}�ǅ�ͬ翧�������@�π���g:��'>�w!?eP��C�8+���9�۲�Z�Ns�~ц%㜜���K�xn1uG��ڭ6�_���~ Tc�_����Qϼ���vu��� �'����J��z�t������,줸_���r�J�V�tR�/����ߠ���k�8��	pRUX�
��/������Y���k���ñ����՚ǰ���N�L�Oz�l�s��ί��]إǚ�6;�o��L��D{'�߽���l���H���늦���N�N����o}i�O<���Wk����~�����ޯ3�~�3��x۫WY��[��'�T�U09�C;��|�❴�=�D�0�*�����s�|O�z27�/�d{���j�c�Nq�C�P���Do�w����P��k��oR&�
e�C낍C�uǱ�Sg5z+�-��F�z�^�t�YF{ª����~,ߠ܁���W��An�7���luG#P�+��u�H��#�Ʌ]��]c�h�l{r�ȸ^�������aժ�Eϑ̀XZs!u?����Tl�����3���*,����KlM��wc����U/&�_��e�kڬ}����+{��rG������n}Q�n��0��=)ʖ���R6t�;Qa�r���sy�]�]��j3�Ep[V�%�2��ݝ�8-��%��$��p�	ʒt讥�x|vwģ���dF�`��T�s�-����D�S��ѐ}+N�^��w#�9�3Zif���԰��>��IT�q�����Ͻ3���ǽ�@�>%R_su�+���q<�|�2��Ƭ9��r�vG�1����m����)ȗ8=c�D�<	/O�m�HiZ*���wB�]��o{��Zcا���^�U�W��>�^
������wT<�$+�{�o�Ug��@x�~�����;�f�C�����h�Ψ~+�̿^�,��y\>ɭF���Fl�ṫ�Vt�3�r���(���-7�Ӳ�x�{7�|r4����X�=��ީ���i������R!�,�}�!��&�5�2��Bg��g�{�Ef��'´��C�"�����9f�'-;�p~������k�r=��7��+���g�Z�;��gˢ���ɭ,UY�wb�9ѷ.��t�8׌mD�v=^��}�B}����Hu�m��RQ���)��\��;ʕ�>B�0�V��d�Dn�h�ɝ�9[u	��F3�z��:�=���o������~��a�n��fO�$k1�r~1�gy�d�u{R3ح��;'8�`��w��_�]��M|M�V�����Ţ1�O�=��ܘz����۬Zj�T<6Ű�vު�L��Y��(,7�Q珎־Ǘ�E�y��eڼ���v@��mE�c���ң��ݹ�X�S.�͹|���7N�Oz~�S-�T?��Eg�޿i����}���J;�Օ���H[��٦U�@�Ft��Qbb��y)�p��J-�T{��#S~��.�Lߜx����*�u�L��8��_�_��!NQe��ǤW^��D��,y���B�|������R�����^�%��S����<Fw��G�\�>`�]�10�E��PJ�Xjc:�v����85��ݙ����U �����2����s��]�{2�,��h��p����ly���T�1�][�#fyt����ޤ��z�_�A�u�^�=X�+�&��)�XН�X���a�\ªח����e��4��Ϸ�^����D&O¸\{ʯ�"��]`V�Ε����S�7�,���=�Q52�+3a�͒E��MF���mj���c5�\�W��e=�+.�}��"|���nd-8M|�����c�n&�q�Z���3Q�O��%,x�˸Sb�`�*���R�M��w�}�G҆G�T��`yG�?�zrO�ӳ���kG�'Ei8��qC/�ӂ��)ߐ� xLm���i��=Q�5�{/�VS�=iՀ��۸�����b�_��� K3y�A��_^�#�w[��x���D}̀yڑwm��ꭍ�`�S@u�k3+��DR���5���mbLEɆ����ݙ�G��d�����������l�v7�������t����}�ʱW�t�x��%���7���;�����SU����({�kM���>�~����C�K�|�F���P[�py`��S=.�cDM��w޾:�g�_��p��Ƿu��t����c���K�ϫ|Rs�W��8=�nF�/1ޙ��}��u(yF�t�,��Q��F+�{�3���fBf�y���^�qϽ��_w����*o:�H�G����+�mVl�*���\U0&/�p�2S>���~��c�������~N,�}z}��R;��6�Tm�VYY J5= w�������%͡��i������fj��++�6wk��>G8�9�u~��d)��u��F���"��_��c��u�F�ͦ�z�b���d��:�܏u��瞾.���D�=�{�����G�)�� 7;��x��yj�F�#[��tL��� �#���S{�������ߨ��G��B��>���F{�:
A�>��>G�d3_Z��{A-�F���{��U��ߎmp+�
�AP~�O�zq�W��n�Y�W�<%�N[�<��47qVJt��p4��:��V�ة`�u%0c�>��/��ԙ��ݲ�HŶ�
����}�W�u
q��L;�����wc�Fڴ��;*�	�ɔ<�oa��{�D��8^��݈ٺ�0�;�ȫuNT��aq��Ǫ-QN{N���Ӑ�^���.a��KtIL���k��Ww�J�v}���~R��{,�ǉgL��n����s{��?�#D���Ιt^B�����z��:}�j6����/�t<���=��iOa!��D�CY;�����J�ۓMo�w�U�'�{��3}Hy9�|t=q�Β>��	�j�"~���K�|����Z����*���?V#�
�Ԟ�� f�:���_�/U���TG{�T(g߼�]�t���!K�H��D���4Oي�ڏa�}Q�ͪ�k���ҫ����r<q�_���o�WL!1�4j�kO������ͭ��N�%����c/+n�Y����Z�#_�ė�8ѱ��\�ŜW�n��)���guGq�x�*��gL��Fa�����έ<>��~U)g�gfd��B|�j�]�Д��9����дz��#ڲ�5��JF�%��,���c1�u �����s#tX�T}����Oz�8��p(��y���W��:�q��m�Y�2�I�*c�w��5�VFѫ�7�6�r�,�_�mb��������]���|ھ��yv͡cr��n|MNz��GYײ{V18P��ҷ�Ľ\���7{�iX��}õ�wi��p$��*/��-��.eu]
�Mol�95�/�x��FN�f�=r�4_V�S�<5^���	1���J��]�8�`6?w��=�~�.�Ō�~��覊�=<p��Q葥D�̉���f�b�#%W����Ji� ȯz�8����P��q�g��Ϸ�>پ�4{< �ꥐ#+u�=��=���C�� �栝��M
-��%����D��Lk�Wq���'ר��{�5�&q�Gw�p����џzg�]�Nn&���@���B�~+�T�>�	+[f��W�km��};ģ��/=tF�n��D��Z=s�jȚs����Ѹ�]~7J_���)?.�A������{*�1:~�>6�{0�N|J&������}W��,���
lc�羒c��J��ǲ>FXۆ����W�<�{�}.pz�z�*���䳯M~�p�^�N��uܝ�
�앧�}W_��O�o�ܳ�r��wc�k>���*���ώ�-^���,��2�m���ݨw9��9Z&j/n��y���E�n��yu���=W=������̻��죇�(�>�N�q������~*NF�`O�(򜺛3Pz�r��f�I��|�M�;�+��:Fnњ��5��"v��B�W�0W�K49�w钶�G�SOv�����	��<Q��������2V�17�p�NV���3�h�꾐Vp��f�.�b�\Fd[�;�:��Ц��U���N��#fS���o@���ޭ�yS����jΛ��n}(i�b�#*�+��(���5+�].��+zp~�ȱ�����{Y���]���\U��<b�	�7%��Ȫc,{������⼽�U��m���7���g�{,vk�x�~�^G�΍�^�뎿-|(�y�5���n���J2?si�^���5��ɝ��V��xR��;Z���j�x�{)��Whh�f��'}�̜�K��ځ��g�dK���Rf]�`\d��k�~9/������9�L�
�����;>��w�*���C��溘��c�%T�;�tX�����Je�ڱ(����dz[{.2�~�V�A<��^�A9�r<V�M:�ߺr�>�g����t+��n2X�;b^�L{�[�<&������_x��ٻhR����
���}#M}~�p�#�^%��0[:`�{t���!�m�z�r[���7g���{�x�7�hU�v�X�~�g�4��������L�����`�>�qd���^c��]i11���%����:���&Y��=�ށn�'��6m���6m���������6�1�cm�������6���6��ll���l���l���1��|c`���1�cmc6��l���c����1���c`������o��6m���1��Cc`����1����d�Md8վ�qI~HAd����v@�����
�ޅ(HP P ()@ ��

��T�P( ( �R�@��*�PT( R�H��8�T�U%T(�"D�J� )	UPUR((P
�U$�R 
"P!%!T�B�s�UR��$ERQ(�J������(EEBR@P�	@)EPD�*)IQ%!�R����D��ʪR*��  �  �QTs�h4� �`��a� Ͷ�
 f2@ЍU�@��QU$)V�P(G   ��P(!P 6� c 8]\���@��tP(�
;qqJ(R������ ��`̠
 �XQE(�M�"�U �	�� � c���-� ���ڬJ�3(H� !�M�c@h"х�I�I"�e�� �  �(*��� �B��Q"D��hh+i�EJA�cZ�Ն�Y�
K*�ږֶ��TEV���D�J  n�Z��T#i�)I�fګQZ����T����ʥ6-��2Ƴ�F1�eUH�mm��m�Fj�l�Z�2�Š�ٍR�"���$�T)�  ����Sk��-Kj�4��,mh�[h�-������F�e$�6�m�[kV��lj��f�VB�k	�2�aM��I���  �5�US4�Zͱ&�ZVڲZ+I�cm���P���Z�i�cB��kC�ڬE��V�5K �F�P�đJ�Z¨	G  �[�v4���M5I��mV�[-h�l�UA��mV�e�ƻ��F�ƣBUM�Vj�m��5T�*�jʵ�����eDJ�
   vK�*��6��UFU���mb��[F��j��0�j��S�4VXm��h�0F�ՕH-F��E2�%R�kY�P(��H��D-����j�3[`�*h���ʕZVԒ6���kU� ��ڦ���X��i�Q�,*�kYB�R3 P��   ��RT�F # � L &"���)A��0��2b Њ��̩� �@42 &@ �~%J)L@��M0F� EB22&M���6����3
m��H���T� 	�0  *���$T�1M6��M4�`�2�$�5�"q�k�A��P�
 ��?X�����A)�!DA��8�ϧ����?J�!�C��l� ��0��EGL#D�*��@��EF�y�t鵊����^[0Di#�KK9�\ba,�Y$���{�Q�~�#R��Ĩ ��5^V�2�kú�*�^q�h���j`�1�3�[}D
���;��&xc���a!a@���C5]��,�X��XfB�5�[.�5vsc�f�vq!GDyyp� 3�ʖ\8��A��V�L�B|Z1SSk$�൴3��}I�[{�i�{o�A�,��Aqި�с����kl-�*��L�j��Tz�Q�>���AX���ߖ����k���U)k�D+6�nR	Ϧ��\	h{Y�u�mHm�	X��PP�Jb�J"�(1	Wl�j3gn��v���H"�A��Ү�ͦ�'Y�~�N�1.��ͼi%���4x�z���:�E�kX��h�S��8N�>����V�:kV*KG�)aҫ(U�y��E�w��-���ZŅuzj�7���Qme�s�4ŗr�!h��͖�X)쵗[��57n�-#���#���Yf��7;�S]��9�z�"�Y<�,0���j����f���4M�����A�l+�ih�l���kL&�x��n-�����H��R	����2���|�v��wD��d%{Im�h��m�v�]?�S��ԝ�J�_��w�d 7���6�
p�:���𲈳����m����g����l#a�[ ��I���U�6-���n�Ve\��	�vP_)�܎����P�K�N�x�cM��;�|]YAT�d���h��@1���qٖ�FL���#{�%�+wM�yO߰VV�Gj\&�t�:WqV�t��P���Tvv�fe�RK���V=�:����#�Ԃ�gc[ذ�;J��E�ݺi`Wb���S76@��\x�'U	yN���KZ�en]�U�� �n 渲�a¢�VN���\�'qi�SK�b�.7�9%˘�^��C[�^K�Z���f)���9�p&ef\�-d��KZ���j�(o�Ĕ���N�tQ��8JK{yn�y�6��HkԞ,� \��JI �ӷ�ި����WM�[`)w�@(�O7C�=�Wsh@%C���7P]5�;�Z�~�Nm�,�1��w��.�JDm��34�S
V�W%ٸvQ�2��M8���񶐬54�����u`*���q4ј�0x��>��]�9-����.<����ݗS�]���Ԛ�v��Gؙ�`��0�f�9�P8�t��]�n[�dŕ�룸h=�Le7pɖ�6��D&L�����+��W*�]@J�Y�p��Im����[M��K*:�M��W� he�?�Kw��ƠϭQ��ʌ�Z�-X�ݕ�ЁOp^eVݬ��&�ɺ[9`%x�b$�[�PoY�Y�>�/
�OBٶ�Z����o@u��LeG)�lX�%e�e����a�Z��su�̱meK��M�!Ҁ�LA�漋��׈mFo!uv�IٳMY�"h%�cU���j�v�j�t���f�:�׿I:)���Vb;�{�y)�����S��GݷD�!�7m"��N�����,U��P��2���ڵ"7s�Su�U�Ae�ұshe������j�N	1Px*���)I�e��A�y�����WU�/1�Q���0��fV���^�ɴ���c�BƸٺl�v��=�tS��-\gj�����]�T������Z��Xn�q@n4� ����ce�����;��RA}���C�A�)�+jI�
�B��w��`���ҙ��7+/[�V��@�t�poiޅ����u�d��e��k�d×�@kD�j�7z����R5.�J6�u:Ɍ�Љ怭�^�Vb�H�f=�#�A0�wSoI���si+��a+U"�I��YYMP�:��JW�Y�>E�^��O5����b��l,�{�Q�t�-T6�}��T٤��r������[:�&��GdC[2�$r��,�ԎE�Mᣫ�JKJ�3�����&��'���9�&��F��;��ُPb7K����Lܕv�\0�ed+Ec9fhE+�k5���6���o�kh%��w�뛚�Y$5.���btT�[z�&4�YRe��]D�mb)H��$�e9LݭyEQ'͆#����۲�F�/(^ned��ʰc.�cb(-&�U����N�V�n]Z�ʻ:�m�%�V�.9wul���l��C(�v�h�$���]�V�+q�ӓ1�'c`�����A�L\Ī�X��@*�a��XN���u�2*�0���*�V�.DQ���Aߵ��.Q��?���yr��ywIc�U��Y3�����5�+J��ݝ�m�Gu0]�W�H,,4�7�1�{:���ݛ�,��F��x�����k}V�\>8�n�+gp�)Yu�;ћ����Φ������J�f��z��9&��xkE;F�*��V�8y4wF�O�Qթ�
����j�u��Pu�Iu��۳ep����^s�C�?���%hjH����n�sQ�[����Go����'�pm��e?��6��!�-$Ǘ�b�͖����s���j��DgV<9��Op+H66�}�)�KJxRK{E,�h%���]��tN�#�5�/8il�C������+�㻋��-[xj���*�Q�-*ř�V�" X!�Fb�B����ƴ��D�_"un� NѧU�eŵQiOa�kͼ_n�J���)G���+&��3䨇���٭�V�M4�F�>ϱk�T�!]�U�u�[Q�EM�uwNU�ov��Lܨ�����v#�e��N+h����`f4�o�e�����Z@�4����W����xbÖ	܁���&[�&a���&�H�fV(:#4م�Y*Gf���Jd�+EX��wj�@�)�B,a��X[����8�e8�U��`k�E,���<{�`��E(n=��y)�Բ#Θ�.-S��v�1y�*�G�㠒h��mV��׬@^#&i4���Ѻݫ�Ea˴�b��e��JPf��C���Yo.P�Fв�`��b�
mh�u�&K����+N�&�������Y���6���Xi�b�6Q�n�%��܉�d0��^��܆Xp�jlEb8�;x��&��'e�����骀��A��MYȅ����jhւ5Ǧէ��a�u�ᣬ��Hm:�7VVL���aFab��ֶf�o:^�3�F��{�셑�֖HᤶVV�.ڢ�R�.ܫ�Or��6��4���jhjX��{̕�1e"h�t��$x)�3]КRP�E���yMŶ���,�2�0uXx.�ld�ز�v�]�8$	U�U"��Y�,ԛ�Kڰ��5{�u,+-��ve]*}Z6�ݴ!Ǜ��7��/u�)��b����Ա���F�Ji-X�[Dև�AAa�mI�e� �7��l��mb���^�wy�DձF��m9�hP�J{>���&�C�D��|�n�8��K�M�56�+ʌhkr�E^^�n�IZE%�B�@�vY��.�1�6�ږ�b�qP̰E���kwCFf���̈́�Y���#dD+hh��v�cPH r�֔E�l����c��,�ѕ��"&�a�����F:z��*��	J�,1*Q�B�����j-.ƛ)��k;���&�:�Aҭ�9k�k�����k�]�E���J�8�0*.�b���B�D��Y���}ɻ���4��x���e��
��H���b�3�yzL��T~x0�mKv5d��OT;����=]f�;j�9t2�!���s���b�n�]�N�\�޻U�v�	�wW j=Y*�<����U��2��R�	p�D�{�-���7eށ��8Q��֪�����t��g<�k(��YEZ��3 .�p�X�jj���9���U�Z6�&�5�qSу/6�^g��T:+���hʧ��P����&�j�^]!7@!���LP��7��@ޟ�R�[��J�v.�2h��(U��I	�"�M�>�I"��_H����+��
\7x����Fb���c]<�*�q;�J	����@��ɹ���m����:f����*@��
�m�XF=�d1[p�è��N�܂���ݩ�A�>�z��<���,i���Ь�M��|���CP���P���O yAQ�IGy
a]��a���pAQ�wǯofd�w`4�V�T�	nQTM��V�{E��=�2�u�'���/.����M e<�ݍ�2�IW@���V��0���k���|+,�����/�άVi�,c�ɧkm(h�2��f��>T�nӭu�ʡ��V4�HJ�Ar�Q09u!M6km��b,���X���'�H��x0�Y`�f���l���d2@��i��_���7��SN�^C綁�0�ڴU%D���1N��-�k)t/�ʛ��4mnY���M*��:�+�zFq�qt�HZG�C�;1%QY��Q8�莱䗸]�r*���0�>�:�0�����}�]�� �
s��m�� S˰.KSU����V
�o3w���T�P�(�ڋx�{(걙�����R��(���f�r�k[���L������Y��ˎ��ն�Y�t�ռ`�V���ʌm�O" ���Vd�ˠ�6��v����W"KX�7���� -���] �υ�u���ݩJ���M7��u^������Y�/��ob�*�\��L�4�5I㊵d�]9�D�h�f
 H51��a,�ݰ���N�n��Yzi��C�����-S��6��X�˻Q���R��������-2��`Sڃn͂�j�˃���^J���۵��P��(`�r(���D��Z�4b�H�yX������o#�6ޒC�U�;�]a�]X�7Ն�M��'Hh�tk�Lhz��@�Юq�թ[F���w��v����jn1�jbG-oa���p�H��k8c�6�X���/F7�(6ef�� �/��y�7(-]�Cv��Z�ऍ=�A'G3T�)�̻8$��o(\Ym�� P���Evt��;P�\�f�򐣯o��Aܬ���HC�e��1�{Y��VPF2Tyyc)L�U,�,�مſ	�)��)�Cu{�����U���-�	�p�0��,Q�^�b)���t�6��U����Xv�muv�f�a4n@�"�Zb��ڒ��C5�٭���x5��7���oaTq��.� ���E�u�
����H�=J�nʺ[��zb�	�Y-��P�;�<��q����M�\Wu��m�^m4dǃw`�f$J���a���J9���/U[����S�Bb���$�;0l	`���ӱ�:Q���dZ�̨zoE0+�
��b"��2��U�ih6���3�G8�e�����kh�/1�F�YG5���5���zu��;��_%�l��r��;B��{��;Dm8r�+8�([GCACv N�B�Ax���ĥ$0͕�r��Mڙo�U���8���7����kۺ
�����L����G3����6�%�Ր�kM]��<�����
˥7YD���>݆�ݼʕ����\��xR�VØH�yA��N�t�6����&�8���h�n�9��E�3i�xwWmi8e�K�k���"�-����7��+y����,Ox�<Me�и�+%�dK�[�F��xҰ0�Z�^冘����q�D�D��nl�k7A�&��.VU��n袠�h-Ӓ2m��mD���d;Ws��K�4CW����0�[�ɣ��w^V�
@�n�ŀFMҼ9�<Uz�v��]f�s��}y�%�o�F.�Z����oq��	�Z��5
#j�&�M��	�7)��ѨV)F���/�ja0 �i��4�Ocr���é��4({�!�t�d�N��=f�b��Xop��O+W���tJ.���FFF�&]c#2N0�-kN%)j�6��r��@��)�C��\ucb�k����ɲCY����|o|6*I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�JI$�I%�fƤ��2l�>Fk���f5$;���ͳ�
qJc6����^}�YU���Fl�)St5����<4���u\D�Y���_��$���I�7Ҋ�Āz�t�3x�Z$̬X���6ȁCw�k��j	�/]](ҹ�;�1̦�]�x����|#k6�w/���O!���H=���xT�Oij�ɼ�d:���f��&t�K�Ն��=��*^��{�}�w�.k�s<wWH>���,j������1��aT+*������[9�r79�M�V���5`öNq]�S���8�����2�\;5$����G$ʕ���32�p��կ��c�;y�uن�Jf����6��K��9Y]޴���s�܏m`��R;ԐNt��N�c!�9�:�P��DI���x�G���^���<�p�s���RWJjQ�JܧQ��]�����[�V�XMn�HT��-��v�Xq�9�ᇱS�	�J�k��'[rPG	���]�`ծ��7�Cڹ|�N��W��ԫ6��3:T�3d��Q#u�I%���66^�Yuf�5p�x�]�u#�����T%���ӂU�3z������Z���5ڸIU�%��+c�Z=P�/�	�"��$�kJ��㮣(�I\��pٺ�|�G���yͮU�h0�{T �v�ppd���P��	�0�s��:i�Gy���^ĎQN��ؖ�3bV��Nܣc��jvÆ�Uǔ!�����X5�"�&][�5���E�V��R��� �>��Z�R��T&�k��2f�w2E-bͅM�!�;umP�
��ۤi�OR�j��ڜ-�y.*߹���0�X5=�:⣹W��-L�W�s(jz�s{�c@�ժ�Ⱥ���,t$c;�uE��.n1AV�=�w0�ӥ,�Ѡ@�u�f�vV��9PtZH�b[���g�I�y]�p�Y�ٗ+����b��%tl,@�� OD�Y��T����m�+��p�[y�xu��LS#��N�U��i��3��*w�wz�dWS4��vK#:V����hȵV��kC�7i���{�q��
�>��N=V�f��аOm�;����+J��4B�ze��R=-�׳�]A�WpU��Wcb�qk�������OeH���e_�Mw�T�����L�S���]���a��v�)0VL��XrԪ1y�@��4�Ž]zf��
���]��.N�
�IE��Ғ��P���Y�TVf�H�,ӜL���L&��=�0��!#&,�t��ެ����<���rg ͂��l��0�N�~���y�]ث�'VH��:�3I�H�EnLWjس�=R�Z!�"UE�L��NY�kc� �ś6�.��9��ti�;��bQ����3v1���V{��un6mǝG��+�0@"����"���[�K�����Pw����Ι1�Wk���{�h��W�wU]�N��5��v����c-�b�E�W=��L[�8qV�x/��u`ʰ4�@'Z�B%LGK����<|-�[���6H�s�Uu�M�`���9m'�C%y��˦3yО�aޓ㢝(K�M�,��L���#U��
�l���� ����'���ww�2�=���̉P vvF���2����rƻ�QɠF���|0s��yv�d��)��,�r�Hb]w��ְF�;��)�mD#�:)���G�ԒRW���bS����*��	�̷Y����f[��0��4�WXa:(%�ER`ǣb���ҿ�>�����,�M�sON��4k[ͭ�v�g[kU�?1�iV�o�l��oq�g>_r��X��
"������o��K��Dr�vJs���T�>�4� ;32#[Y"!n����J���-w�C`��rWIN�sKb�H�Y��B�efL;�<��t�2�̋$K6=be�̹g�"�^���d���k�;Cs�e^+�p���ٹ.b���ը,%8t�R�"Hq��l� ��1偺�hq��sb������؅A�����"�KX �4fA��:�mԫ�8upۘ6�ZxT������k�c�3� b�u4na�ԋ|z��]��Ox�{Pq�1�&'���蛮{H��@���=a�2�R��W.�Tu�&`%���[s졲,Ww]Ե�lH�]O��Gr�G8Z&F�9z���w�`�1,��f>�w�V�H4�`ĪѰ��i�[�8\ ٫�'gn���M]uܸ45q姥�R�ݐ�����ۋb ��F�C��H4���a:��t�!��JE�w�r�t+��ITf�i�K����们���/u�-�bY�����I�	�ʷ�b�%�2��e�#�n,躽葸�4]��O��:�2];�u:խ_6HAUڥ	�+(卢�ʮ��ӰrD='��6MW7��l��%�M+p�6wr�7B�S�9L��ec�+����[��1����8u���,YeZg��\�I��Y{�;�t&��\'��.p�8�-�{V��IB�+1�	K3;i��:i3^�5� �������^vNi�싷�|�3iE�<�4�^-�*�z��>o��4�Q��V(V�k.�'uP}��q7�Q��74f���y�5^��>�)���L0R���ΰ5�j�R����C��HJ��ݞ�i����6�:Tw��v�ؘw	���]�t�zom��w*6n��l6�a�t�Ys���m�.��DsM�aB��C0c�������;�jU�6��&�5k=r�� ]Һ�һ�zKZ�P�6�ۺ1��)��z��Mqw�v-g:��A1ʄ��u��EVe��v�ۮ*�1]\M�l�ٓ��〵�;s�F�o���R�Jg�}�A759����v��iV*+�^�K�+��t���f����ր��e�v�ڦU��ߜܢ&���t��ƪv|�JkqU������{a�Œ��u/��T�0�7F�V��j�t�<�xF*����D�ܮ�;5ju���['q]�gx޻��T[0���]zBW��w�Ŕr����!'[f/jrm�}����9��xwI�i�p���Z&�k��n��>�l-\:���Ƌa8y���QU�4q�����W��Fⶾ���ev�׷|ʝ���Ѣ���|d��M����e�M�^��wW�ަfݯ����2lH�R��X��� 9J�;�Zj1v�X�P���4t[g3�q]u�͝�d�Mk5�pQ�"���Ce�Il�ڠ�;��x۩�S�E�z*ﴋ:)5F�$�#�v�ۊ����-֛������Mp�� ����n����Y��)������ޭ=�I�L�u����mۊ�.�6 �l�͇��s"y��[Î��v���q6����%(u8|�u]w1��;wL��vm�"\n��bn�r��h�A�Ɏ��gd�P|�읪k�fw0�QL�����F�{ζwK���kV�� 9:�+�*ˬ�c5��]��ɱ1$��a{Z�>BU�6�ȭ���7�w�ff:�K�'g¹Ĭ����w#�v�|Z�ժ�Κ*��ܺd��L8��������*�J$�m����iP1�ٗ%_�NX��ͦ�n�޾ճ�T��VN@F������Z�Wa�&bgb}��R����:��JJ�Qa�|m����Os��]K�/m�՘��c� g��d���a�z�=�x�o�e�Y�9�X�ee���$͕h������kw�@V2�J�����K�wt8��`�W���εԢ3W�]C��vXn�$���* Q��n��.���:�����9[X���ȶ�Ә�:�m�W�^����k.�q��ʣBm1��֊Z�A�H!α�t[W@�X�����j>:l]p�0��t���1���u���f�����3�bV#z�*L��LMo�ok}���o ��6��mGƲ�]}�tL�`�fL��sT�>�ܥ��6'{A�<7��s�)��
W8 =2�F��1�.p�ǽ����/�r�� ]�;�ujza�x�
[cQ}�Eyqn�}6����ݾ�ֆ��rS���S�eJ��B�X���GTvm�RX�5�V�xN	�i�̹��su�ȭ:k��$m�uU���L2�E��ޭ\M_K�`�k�q5�++ {���$�T������#�7Ħ�LK]�Ľuto7  �a<��)¦fH{:�&M�����&��r���o�A�i�m���%Gm��<���z�.���ŧ�H��Ln�K|Lt���BU�\�+ԥ�N��t����ޱ�X���m����d��m \�{pZ�G/�q�a�yݺWrq86̳������2A`�7�]��p�/�q�ve�]o/7s��h�]�f�]�O��r�C3B���n�(J�NaS���Lh��c�+�v��(U�힐 �7he�J��#b�*�rz �W=�H�3ۤ�K��n�M�A��Q͕�C(b�2��R��oVSm�޲������Y�#�d&j"�cj�kO�o�+S����Kٯ�OoXƅu�_9+�*5ӛM�Yg%`Cd���M��=����C|3��sm8����Z�S����Y+j�ĺzv��R���iLJ�4#սSp�k��j�A�Y�j���b%�w�Ga�ѽ�X����]éʑ�i7�X���K:��Yf�F#<,��b����7	��s�ufm�gM�7�4�o)@�̳�#��8Gie�A�9�z'�k���7jv��}Q�wZ�pt�����m���OUqc4r�v;\�c�"*�r�˅'���	)7NMB1���S��[������-�k5J�M���**@��Dm��tv|�֟A���x�	4�pݦ�I�xrX����ԝY�N!+�SO���Du+����Z�����֝oh�_7n����Ju�d39C�@0V\�Q�v7x(�I7e��%�݇+̥�ŧD�r��!��O±��2�ѝn$e�ѵ�̡�'��6�kl;�\_l)�C�$�sL%�;z����������a��q닪�`�Pb�=%H�	$�T+FJ(iv-���&޲w���Y^�*-R�t��L���;z�.u{tv�!|(g<��#�0��v��ۓo�����FZ�.��V/��Ό��Y�+��̏6�x[���PJ�M3�A�Tf��a�;��9dq P��c$�Y�-� lB��Ie;�B#�FZmrv����jʅ�|���9�ob����l�Ǉ�\�v)6�\Y]p�l�Uе�S��{�{f�F$K��QЕ��"$am��Ƶ�2�'�cH�A�5b�j��zff�B�FA�A��")3��n�i�Q�n���hH%��k�(�	ڄ��@�9EC��89^͊u�`t�*�72��2K%U��ʎB�,�A0����6(��D��IS�-�so�䊔��9��r��w�N�шK�;ˮ�3Y]��p�6��Nأ1G�u���skpv\ӓX���gm��UrJSv�I[FmҔē���yئV_��{w���v���H�i����ծu-Kt����IM�M����W��!B����\rVQh�8-2c�''w)�QA�e��_��Tf�Ҷ'��62W1d�o8��}�T�r�G�����2��̒���R>�$Rn�\�W��;vt��O��
ꏣ	Ԩ�÷�����Pí�;[#R�5M�=X�RH\I5 1�n���q�&-��#ÜJr��%���/��n�ri��RI$�I$�I$�I$�I7x��=���	[&�7#�Dܫ���h,wSc��KA,έ��y��j�]+�-e=�5�ʅu9�WGt���9��(�Y�^=E9��QtO&v��k��"oks���ڒI$�I$�IW����Q�F4i#^u�Ưj ��$���vPDu^�D�������=}Y�V+jԓ���� p���;�u�ٺX�޼���[|��`|N�-l���������j�/8=���w�NxBխ��*Kk zo5��1)K�ô����u':[�,��t�IM.v{o%�\�|��#ϝ����Iq�O1�;�$Mm=�'%�\�21���gu͡�|�����&'j��Λ��kh3ӓ�PMpe�ǖ/5���X��
u��<�����U'V�H�����q�e$��k��q�6".�Q�A`ӭ%�\��ηW��n����4�w�3R:�t����}/E�ĺ�����.��g:�fBv�uOZ")��O�
��a�7��	pSyu�,��h������w[�z��{��k���Hs:l����n��Ic�qŝS ��|k��R��gKZ�Z��U�n���#R+�o�re��t�P�j�-��������'�FN��B����]�ggT����$�vx΂�Դe�um9.��~���j|Y�x��n-0M������wwq��G%g%��@���w����ۛ��nH�V��:[��mG��d阠��v�xz,�,���}��N��X��!�Yp��S����H�7N�v�*r�LÀEJ�{/�X\�ݢ�g'&��&�^�(�9���9�n���%����gi���q8�7��d���,�Œ���k"�J��v���Zg�u�N�2���]�A�9,]�N@j��u�[�T\5�tx�5���p�8��e��Q�nK5/9�pJj���&R��R�Ui�7�e���X�����n _66]�P,i�2C�k�XwgW\�|2���B�)*C{\��m%h��ô�32�ێ��T����D���,���P�;��9g���K4Yލb��BMn�K�ǹ���+sK>\N:�����˩y�Zvɑ����j��H.�"���p��	/��]\�`kF�əNح�m+����Y��5�x��$�[�P������m�hps*gYX�ٮ��S��ɂٹ�M���Q�=�,��L8��-��x�\�\��+V�LY�7�K�<7d�8��)�T�d�l]�M�\�nU {��
ʑ��k�n�76�+kQާXj螴k�Jc�:̤�6�j���Xr��n4�iY��B���JIL�]2C�wb:�dpy��w�d�`���"�r�N�J��޸i�䕳o����4�&���vow���}�R�ɻɵ��棴�x2;�lA��
�<F��'���4�:��Y�R���e��M��戂$�X�k&GR��&:�,�q���+ʭ�ͤ;�f'QѦ���WKk�Pz�V�ט��WY��na�YuЙ�b
-�Rᢴ�i�'u��&��k�h�i-�G
��I\��1���{�o7����x�6¡"e�z�a�\9Q��I�Z��;��͵}���y���s��b^�;�f���g��IA�vV�Dݽ:�4��"`v�W��u�S��-���K�mX30�9V�u�k���/M(X.�p���;AWch)X�R�6m]7�����ۺ��{�i(	Z`�J��W�v���ŷ{�:�j�F4�\�^�<ʈ͡���7� m3Z#K;2+��ÝyQ���t�ڮ�!�P�r΍W�fEM�9���5�Y7��;��&���)��p����k4�)�lm�����G���+\Qr��oܵ�ڬ�wȈ��!�n�)X+��^�5����F���r����ݻ�`�����qj�bi�^�A$��j�6�Qx��3u�c7�h :
�s��^_4� ��gӵ�q���	���-9S�W��y�]�H��f`��\��G:}�Y��[iD���L�Vl��-f��>�rr�,�{��l���!��ͅ����ʜ5�Tz���\��j���l���h�[uuw�kuSi!�l�h��ͤ:`j5��{XQ��`� J��H$�J{���J�^r���\ �T�x���n;�ӭ�"������qʛ %�;�������DZ1��f�U�*�u�m���;uj����|��dM �Z��b�i�V�U"*�lPӻ�O����T���#1Yn�3�5�8fΫ�֍5[|�C��%hό��`櫲}ɠ�E��ұ3{[ٔ�sV=EVTzfu�{}J��p`�:b��>�wa~�]qpb3p��Q\lwt�Qr�9u����>{�[62���
:髶�����]�+s�Xv5�'G�U��{���1��-t�C��&=�]���[�.dy���s�}Q�����OtT.it������:��w�A�=�p�"I�J�+��O:mm���;��3yۀ̉BaΫ�k�V�ʳ�m�+y.��f'g>�PI�I>wh��lQu����2D�$���̭\!�Y U��9f�<e�[�(Y��)_S��B�c&3K�Å��Ɯw���v���E�Qg\齊1:����܀�Ht��q��)eY�n����9�괛T�O2��wf쵧r���uA[��YKB���q�&�
���J��)-��n�kX D�-F��}΀�Eh���8�9N��9�H���ܱi�{��4X�.LY���`�C {c�4��t���N�p�Η�QѬ��F���hS(�0�d� �QJ�z�\a��gZ����^S�f^[['*n��͝���:V�"�5���[צ�V�5���=2Z�Ǖg�3�5����*oVV�AQ�k�]%֎ջ��TB���ը$����?q��L]�4S;�8ڳ���f��T�X)�$�.@y�gA�c� a\"���m:��@��!�ܙ�wS������bLd'9lLͰ�̕���8���ot��F��6�]�n��Z��Ը�����4"��#Gv�s�gfu����^/�.���}�wr��I��	i���l�Җ�V����_J����,Ws��s�lA�E��!�G�,��	t� �ִ�pkU��nR�ΗR�kΙ}�G�)�N&�Qh�"ޢs@v����K ��\��L� ��s��T���>��NrF��[H)|�����-���(8Er�X�^vQ���ό��φ�O~;���ξ��/fB���A�de>�ft����:z�i#F�K�-�{Aص�`7�).��c;��,�N
��Q��)���������QxGl��h�2��mD���'���hUͰD��Mh`Fir��tz�3����\�n�]Qν�ښ���<G��f$F�(��C:ܩ�s�[a��r�TpL�]'@z뉻%�ὕ��Ws�'F*E�Id��/�.eEbL�}w}n��o$W	�f�h�R�.&���U�\�J�;p�}w���֮�^ŻV���hƔ47��\�9��nv=�/k�I�l�2��A�[0hu9�{Y�=�PpZ{F�N�v��'�}�B��rW�-P�O��r��Y��E^J|L�O��}Yt���Π+k	�Z�17�*Tj��m����ˇ��]�kkεq�qi�hC������7i��v�� ��sN�1�Y��L��{b�MZ1+��iЭ��m͆����0�ά��h
��ޭɉ�&�Kn���3O(ч7;�:�%80%Ol𬡻�΀�:��9�������u���olrʏ9�rYkBh֑:������]j52�3-w\���@,DRe	�(t���.���W�4"�_��]��A5zWl�ںj't�'\ն��"�޾�Ҷ�J�]�����i�o�]��(�����Ye]cr݀�<���v;(�ӱe�^Zb7�쾕�k�#a�^(���]l��L�[��y�n�^GA�1�ҙ��GK/�ժýK�LQ�M���Hi
\����}͒I�H���jD���C�y��H�m��r�S�4�
9Y%��$��Ø
��*{(�){��	ؘᵳ0�a24#n뛷\(H3uB���J�BC.&܈c�!���N�{�+	�t�.+�V�J����k��X��7��C9q�5&M�/-�v��.tL�̭�4b�\��v�"�N9u���[N���Y�w`�"����v	��㢎"u@o��������ҵ�ZÇ{C(_0͂�&�`D�vܕ�]���.��Ct�,�[��eU�Եd�K&U�h��oP7ˉN��v1��6}�9�B��[�56��x�nk{)��z���ѡ�s77�q+�"z�� ��Ӫ�Hܥ�Ղ[���`H�B�5�D��@�m��ה8bl�Qs)�w���˳Yz��k�'Y[[kt$%
9�Eqws��z|fEʺ�43�����Ӱ4ɛG�#
�7���S.�kD`�t�uϯ$�&Jȥ=�Z]���vVa����ܼ�`�
�tk1���U����#[g���ڛ�U���73E"u:�䨬�[KS����L�8S�/+�*��s��)yU[��P�+ �t�S4��\g_@Om�i���Uָ������DCF\|���IB-u�:P������Z�b�u0a�BA8z�1woy^����W��B�V42/�Vٔkc���y�R��Ma*�(a�6l#����N��)�nV���7����K�̜�XjL`4y����]t��得	4,+;	�ЙXۙ��E�(�i�R�YϞU�Rn��~L�J.����8�	�<[��Z�,�>ә��}��B���:��u!��DJ�{aR�H�4f;m7չ{WAu2�oj�xR�r^=�S�mdZp��{H��V,�dwݭ�}҅u�j2�����V�췹�s�-�E@m�n����[{M ê�]����ڙ�R="bٷ��5e�E���m���:��ڦ%&ڊ���ѝ�
�R�s�uii�g#)$���2E��r�H����B5�eF�d6uu�8ۢ��+=B���6~m�}��3���a
NF��P���.I`ܱ��
�60�K4�XM�g*f���s	����b��`�BY��9c{+q�F,=&����s����uwR`�(��u��*�+�PG��zfK�+�v���9`
�3-�j^���]�	uu7^-=4t.�]r�Y�u0�؍�6Y��xl!�J��ޡ8�3�27Y�Zv���P�!��%���g:}[z��.��Ѳ��4\�����H2�[*d�e����'ji�vMl�g8N㒮�i����W��:��u�T�ս�W��:S*����Q�h�.�֊}���� U�Z��m���]�������!�Չ
O��ͨ�%|�3�>�dʒw����vۗ�����SA�\�RL�Ϛԉǭ����Ug���eJ�-ڮ�ͶJw�C�}M]�N��c�%�ΘF�A� CY��ua�루䈣5��>��;bG�#�me��w�ѻ|e�� Z���ބD��}�ch�U,����I2Ю��^��M���4���̮�Ŗ�jf�i�����B�y����v��s�d�um��9h`q��^�:���zo�2�4mrΕ
�j��W�gZHͬ�efs���}[j���\�$[j��WnV����;��.���-���������0��,�/��۫7F�Q4gS�K���6�h�e��!�Db��o5)�ae2��_k��[x �0�ݢL�1>�w��h�oF�)L���si4���M"� ��H���K�a-R2m��U�:#_:� r����"�D��vv�Eot]=���م�8��=�:�w�G�VQ�*wtOi��/����U�d��3�f�( A»"-B��z�ԧ=�ُi������X���aw]��aÖjvo�r8GJ���(h�}�m͝����e.\�c�.���	�P�Q{uh�X8��2
{���ceDp�ffu��-JSU�
)dbm
B�N���uԆ��9v1�:�%������3\���]y���F���`Ҿؠ ��A��5-�h��Z��I� ���Y����I$�I$���UȘ�bȲ�"��7��Û}��
�V�i�S�oTǝ�< U�]KY��7{���r�ĝ[*�舎w��m��9a�Ր� �0�XʋhrG�6�����yu�F+������]Ѷ��#�SM��+j�Y}ni��<��B�O%u�[]+���j.gf\���3gP�v�l�����t6�;��wjN���nP�/Q���ӻ趷'Q<n|��mqVTo�@�_R	��qC�H�ڕ�U�F�������5Л�)��˵��Pi^�F�mμ}�J�\�D<ۓ.�J���}�cnd�5vw,O;Zv�Z&��w\�,��6�0�e�V{0�Go:s}kWE�",5�4�v12)f�5|Y�� �6̡�4��1��\�ӭ4e��fU�)�c�\�
��_67UÎ
=W	J�+F���!�;V�I���kt�)Q��I���?CNwJ�0e0v;����߬��^q���h#�^c(4if_F�AY��;v��V���O��I%v��b��شwU�b����M�K��Q%��1nj�2P�ȫ���Ջ��m� �M�''[���wU��7>�����ӵ\xvT �97�$� MǪ�o@�e�Y�g^M�U�7#�����8jsݖ�z�hnd��_7ه�rD�P�\��nk)�$�^�q��rO�}uŗl�kZ͙rЭe��,��8��̹H�
�*(m$�LVkZ˫��ƌ�1(��1�i3*s.:f&2�w��f-�L�Q��\V��J�Lѭ�(*�c�,�r�[���Y�Z%q¤o��eӃ���t��AX�������5SF�ơ��DH�8\�3)���0G[%Us*�
�M�.u�W
bbUwZ4�U�2VTr�4r�:u�U��dX¹��8��V�k)R�l�]8z�j�TjZ\a��[m
��˅EQ�,�p�BԡZ�ҵ�*���3Y�#e��ˋ�6��9��v�W��2ۤ�,�S>���t+�U���ˌ�J.)]emTh�\��n�Z-��5�X�nSJ�!��p�e�9�̕��4�L��+ms&��I���LĮf"�5p����SmEr�Kl���Ƴ�iE���m�!F�J�L�E*Ѧ��e1��mh�..UQŬF4���Km��EkUr�Ƴ?��n�suq��;�lTэQ�yQ��ܢd���u�5�����!��i����&@6Rת'#r���.�%�?د� �0�7��L*�k�!{�R7����,>�w[���r�����}�f�*�I���pG^��c�j��ۦ�V�ڬ}W�c�k�=�=�J�U��l��!n��c7�W$��.gf|sx_`x�����Sb�yE��(�Ӻ��J+y"�B�8���$�89���S��{y��맶�/Y܈����޹��j����qW��F�D��m�/�/��\f���W��T^����b�G�+4��0zʽΑMU��)��;|�r�<�|���=��i'���|{��{1T8�p��3dw_$q�*ڪ{ca	�n��w*�u|�ۛj�`ali�Ǧ\����¥S:���>�T!5m
��U<���[�>�.�u}�W��f#j���~	'<��b��и�v�l�׼\�$��l�q�u�sa�V%׳��Z��4���GD*QX|����+E���pR�<�e
�Ɣ�V�f˹Vx�&���[��e�.��E<;��ri�M�ͮ=��1�b)w�&���y;���x��u��VeЍt���PČ��.�Cor�U��{�ܺ~p�q�K���^2���¼"5S���u:&/���v����69�ݵ��ogC�o���� �Q�O�[�yZ8ؗ�!�C8�_\�/"�9kB��ZKaq�k�!�����c�]�|�]�TR�N;�(��P��w*�]1�|�כ9��72�w+Z��S�z,����/2�y[�n3�ne7�}&�ش��+m<������u�@���|�VGX��E�X״�\�+kb���g���<~���P!2�G!��p�V踙��U>j���[ֹt�L-�y��Y2fP��q`���kf�U�^�8�*��M�S&`�}YVĵ�6@v��%���n���t��oS�V�нlݽ��X�њ�Yx��BSj��v����4�^�����[�d���q�sV�B�w\q�P�Ch�B�o#(���WQ.	Z]i����]���
�$�Փ��k�\���=@=��r�`�Q�l��v](�	��ی�H�T��l��lL��'Ԣ�#-�T�+��ے�p}�-'��FE� �"Ⱦ���i�@ǩܷ�|�u����'�M���^�9B�ݺ���]R�\�c��{M<�T"Ц�4�^���z��bW2�����]�nq��ݪ��iFFS�h`�L�t�&9n�ֶ��Qc�R׎)V�}W>B*b���ϫ��%Y��ޛ�t�c�f�������%>
m��($�S����{թ�Ȉ���z�%���.!���h��SiS���F�*��c��Ak�k��f�IU�*�P;��wX�m\A���V�\S�\6��&�]�Ɏ��Q;ۅ�>Ѿx���u�N��ٍ	Z����)x+�Z
��:�e�6�ea�F5�am��C�6����_n���M��xPJ��\�`d����ڭ�s���6TeJl��<f�"�J\�z\�:T3�?$2�]ƌs����_|Tn=���l��!��ׯ���ۼg�u�+g֕dإ$Hm��1:�-������^t�Q��]ÛyT&�}�ͷ84Jy���t�E��e��q�s�v�@7�m�s����ګٰ�|���)����0��"3�%0�卷���(w#f��3�	��7*�C��;� �p�F�ͷ �U)�/�:zƎ��ÉG0F35>�2�Է�(G�<LDX���w{��[T�}�;��u>y�"��]6��lGk�c�è�眒Zs*�:��k�^J�%��`]v�1��YW/�e�덧������k7��S�Sac��O�-⑁�B�71l��랸I<����%KRċ���kF���ך�޽��+9�{,ᒅx���]���{R��c42d]�)U��Ĭ�s=cA��Ɏ��pr\�E����6I�|s����Ӥ��OSo)_Jfӂ��;<2�s{��/Wv��rkakS���a#�x�cutG"B�(;�����2v<�c�3�v����3�Z�Qn���/��[�/71o�HOE�(F�1	���2/����j�{V���Tw��{5Amz��\j�s���s�].�x���\��\��1��]���h��7磕@�v;�S]=P땘ժ8�N\�,�򞃉W&?B59�~IT+�E�t��v3`�ݻ��^�f��L�+bE��wU��[6)�p-�o��É*�n1Q���+f6H��_H�R/�c�WM&���y�#Owa��Z��0��\�b8�����_Z�L������&�rU;p1��/y�F]�=��T#K�k�(�!K`Ό������)������3�n���fB8N*�U��19R6����M���3�Cl��Ǖ�}�_[��V�9@�d|fW�Z��:]�m����1ޅ`0����7`�z����-G +zQ�F��{��A�J倜+2,�=1��>��Y}I���Rղ'#�_gv�%5�PhlcLPN��n��Yz�)�t�Gb������D�9��F��B�.�3a'����|z��碒퓷�3.?�Q�?��;���k��}�g9k�Ws:��s��7�һA!N�rf��C�Ѽ̅�y����F�qh�n[{�-��p����h�3��ɤ74&�7�������ꞙ���;U�V��^�E[�	ٌ�Q�E!�I�Č�ԫjmc9	�/����Xͳ����ĭ�d<�H�R;*\���uK�.w��Gu�˜�2��{���=�y"�V�zT�G�ҴN�燤�%�t��y�/}�rض�XjH�u;c(ϥ�{�,~̱xnm���Tk���x��ǛW�ȴ���Wr��R���G���x�Q���efaݾ�d 1��K����<�ӽ��w\��8���SV<��ܖ����r'����S3��y`�F7�Q�O7��7Ѷ~��e,.mr ;�a�j&wk���KY�2�N9 ����B���O�o�c�ݫ�Q��"RF���L�x�앳G���*Bvq�2����%LV���,�$��qNP�<��Ƙ��жp�+��S�xM�3�;f�r�A�.�{Tञ@�)�B��1�̣9�R�k(y(�Ni�=���!v�J �I<%3�C�<��}����e�$���2�aE�k'e�CA��¯�j��ek.3�s;���;���S���t9������I�h�N��|�d�'��bRM�~��B+e�ʹn������m���@3b�ncݶ��us������
 �ʨ�"�ȹC=�	�3NVӒ�����Q�:�pk��,�>n�+v��L���w�Ek�6x5�S\�.�x�%ȧ������Y�Մ"�>�ՐJ�}[[�]��=y�,S/�O2�ϧ�ɏw���a(���]�!I3�-�]oj�w���J�̤�������C�>�S�%: ����\NC\��K��_��9 K�7�ˢ���Rp�m��CaV��j.�<ީwT&C����{�J���F򰡛�г�v�xu)�S�����Pg=�m�����b�t>N�݀G�kaC�}�՝U=;X!�s4�U�oD<���W�ҽ��O�skK��Q^�u~p���Cl�h�<�������7Y����i���	��OBS�*�5ſ40�{ж�}�s��7�FLS�����mO�Z��h�)�&��5eA��j,mg�w�4J�!��\�����nl)���k\S��A�fporB�k�ڝ���N�ٯM�NV��7��	ЬJ9V�)I����/��dn>�:"�x��]Aܷ�c������'��2�:���[�`oҩЊ�3[�r�3Xz�(EY�Sϐ�.Ľ���en*
7b��$8����~��B�s@{˛�EԺ۱X��z��c-�h/���X�W��є9&�J�ވR�>��Tq�I��E��[�l��5��/YqW�O�������+�J���j!'��4�K�����޹O�]v�1�k)�ww�'D)��w���K���S��T;�	mEy�ZVJ�^�Un1��x���D>��ᕍ��H�Ŏ�������3�wǠ9�����;xt���\�1td�Lns;���6���O�z�^�=�-n�
�Pá��rd�:���L&w��:o�ٹ���$��ܷu��=۱N�ځ�V!Q�E9��۞#&[V������RV��g��Z�=Yd.����u������cZ�2�y�����W�s0���vJ�u����J�` ��O{����tEdr�w���˨z�9�k$BY]�"����U�q8��ڮΪ��N,C�
��Y�p�W^����Q�/�-T-'�oBu�^�G�F���U�:%��:�m��]��ݬ�m�b[2�aU�K�C2v=w�*I7T��M��<��SZ��qѸ���\����ӥ|��Q�"�/U%�ʰ7�����zes#��+�Ҭ�)�Zǝ9PVS�ם��N�E��0a,�K� �����[xge���*<�n�k�z�ι���ȡ<�����\�پ�S�
ryZqE�S�U{7˭���SV!�!#pZe�'{�2i�iz�o�9˫�l!pw�LHI�h��0`{����5 ��O�yo�0��U�s&���'���S�ޕ3όm�!o:6g����0!�V��t3g�e���õTׂǛmn���ٚB��V$�&q��<���93�N�VСy�͊|�F�J��:�#�M	�ȓF��Yt9{�l��Y�����+�b��/G{7�'�	��m��9J��W��l�;�sHm&{�(q�|#��@2yL3�t�}��ųV)eOPt���XQ��Ż��_�E�X7�)M��?.��e_9ڋj�f$���h��k���9GUr�q��9oC�1���v�a&;d�%A*:͵�%�b�keJ˙�ݩ]u�b&��*V,i��o7Y�D�/�[p��+��0�Re���5����^Ԯ`�6�X��V?�qm����in⹐�χY���ƟN�F��7*��N�Z^�5hj�Ð�n����#;��;w&j��k[�zV�m��g \ճ�܊I͛&�pі�e`�˳��Ч�}���́�1\-���
Qy]�uk9.eMr�(��r���D��E�e]"���1"��:mn��`y�%p iۃ$�y-��+�4!�nr�/�&���/�3m$���u[W��+�
�zU��M�E`����~Ӄ�)R���n+t�O�<��؞�˙K�2���]L����H���[k�L�ݡ#�YӸé�f������t��Q�,���3��SCsj�,��_b��a��X��Z9��J�0QK��gVF��B�Ӭ�,�À宼��J�XƥІ��g
Yk!�Xr���(w-���|�������U�M3�#N��qdjy�����K�\��A�'E%P���H��0�V����-�>W�:���t#�p�o^�sVp���䵤��$�I$�I$����ٔ��μ|n�d8ŐH�i5qd������'���N�ꙓ����6魴�\pQ:�m�P�ڮյy۵1k���6���s��}��e���_
9���pt���6P�s���B�/!,[�ӭܜk��g]R��ޥl�+h�"�r���^*��dzԒ����x]K����`���+@,���̢�삮΢��:�TD����'JGHW���(�ojωѕ��oWB��)��o�̼@R��|����1q[������0;�G	ì�ڊ!��wA�D]�����H��u۫�A'C�`[/!�ȝ�a<�F1n��IB^�j�B�(���6��)U2�0����aE<�a�����\�ulb%���6Or��*�.+���܁�`��ƅ�_��u�]�G���ݥ�v5���*i���A �	�GV��W�N���v�%WG1��H���=��s�@l%J��t;�սxS�(�h�[�Cb"�	�a����v���5�lL��܄�����a�R�e���z�un�*L��ܚ�ۏ����O�M�9�;�(�R'
q�F��ܒC;��܍�?}���?�o��bֱ_��,r�1��֙i�5�ʪ�5��M%gɭjc�&��	FR�R�uprҕ����1�_-BQLh��Y��k*.&d�[+-�b�h����\2�t�QGt̪�����j���0��*��A��U(ȫ[h�ֳK\..��˖����+D��n`�v�4�*�s*	��ۼ�����m(ڗ.c��kUۧ+P��k�h�Bc��ʦ���2�iuM3�\��0m2��ˆU�KFй�V��)kR��J�TT�t&�eW5�ɆJ�QZZ*�2d�5~��UVxZ���nem�Ķ��0SMwO2<�՚i�f,4�t�V؎�W
��̸��L¢f���oM�2�˃��*�U0s%Ue�m1�SBنE2����e�+L.�� �-�33�i5��R�p��i"�E��wJ�Se�9r�k3Ekk�L�2�S2b.\��Sp�KU�e�Vܺ2�b��[��&ٗ[�q\h�y��U54�Mc��ю�f;h��uMkX�hݵs3�muR�)j�V�-���3̥�ۼ���m+���`̥�Y�.7T��h?l��PF�j��3-Z%P[|ޝk
ˆU���T�(�B�@�=�Gs�u�9ڳƆ�d�5�P��]��8�͒��ii�Z^�֜;��y}��|I�L�W[���|�(��VI����cUh�ʚ.q��U�	r?Y?���yl߹���T�dQ޷����g�&�C�6�L>}�v���3�}��m[�gu}a�[��<����0��h,�|�W�5=|���j���7(|#����C�������B�O2~��AV>���ɡ[�9U�����|�>�>���D�~W�6��i�]��ژ�
�+�]R�|���)�ܾ8��4��l�2w������5ܑ3�{W^��hV��$�re#0>	���6!duzV�v$W+�Q��ȵ;�����e�+.��Ͻ�a�u��ȫ�U�FC��z��W��-�S4HkL�9�^;Փ-3 !G
���U6(��22�k�5������:x��^L);5����e���[�Z�%M��Ni��/�~�]s�ۄ4p}�vg�r_�6*�V݃��r{�-θ��5�%&�1���t8�j�'�Ux�7yԮJ��m�,�OR��vky�'2Nm��ƺ6�u+���ϩ�H=q)#���Y:_;´�K��`mV̷J�M�a	��];�íp�L�o����W�Gۛ���:��R�K+�<'׉W�꩷!ڸ����z��W���߆��/��6��n��ed��ҭTDg'E�Or�u3'�<�ߵ�>N1��N���T�!1r��EP/��N�V�Y?y|}�hϑ�߭X��z��$�9U@eS��jq�z�&~�ba}>�O�۟,ĩ�P�7����*xmB¹7ϕN}�����^/��S�i�=��o���ym���r�6�.��(Y
�Ɯ��gƁ�+���C���v*#\9�֩������NĄ�$5��g}��
��r�)�xԋ�=b!v��Yu���x�}���n��V͊RD�����1:�.�4n2���'����`��`Pn��{ǖ0=�M[��jd����'wM�v��{��|Zy&�:�:J��%xU��=;��o�nK�+�ӧT����/�od}��8���T���y+����]��,Y��� 8ŭ&�s"/�Z�T��y34���ps�%��"]�E퉉䱩R�Dbh��齖/�Ö��Z�S�^i��x2ˊ���V����}P6<7�M�p��7G5�`իș=Ϲ��7z�ތ���V\��+x���{ܮR�;#
ם�t�<�e|���;9�ć��{y�"�@u[qf�	33N�u�˫��B�s�c���]�>00(�]��yQ��p��uc��mqś��uz��g��������[QM⡡ܜ�yQ����N"#_d�s�E>�,^'�5#^V����YA��Į��\8�w���X�~�=�&"XɊhm�f/�rR:m�
�-R٪Ź׭�ޭ�9j�U�m\d�搏	L�_q��m��z�Z�WǩV�s�����v��R��V.�|�f螙VUdUS�f�Gr_���q��ߓ���D�V�԰GI�"!J�[�;p�� ���/��*:�	!�S:sW�]IՋ��g!�	R��
RG��y��"v�Z�Sn��Ա���c��F.p)��c7(��u��)�7fǊ�uK����t��*�϶���癹�����kv���ڜ��m�ו>��`�&8wnfu�w�9���/���;IX�ɋ]�8�{�����
M�$/c2�owu ���cЭ�=��U�v�4�S���䐮�����}��g/�F�`h�<0�#�=�B!�
��j[�r7Ϭ�Z�vR����+ҙ��)+��A��৸��k5N���.�������3߲VI�yN�6����xɖ��̐�%a�Qa:ɇ�,4���ٙ	�xɯ�2J��������wܻ�M����߾��xHt�0��x�2M�Y>E��H��a��� ��`u��B~垠xɖ�ݰJ����'5?X>�Dwo�?�����/�����i��:~�����	�>Bl�!�N�7��N��.���N'��wVI�y�d:��Y��m����d
��=�߯ފ��E|�>B��3#��^���a��7�%	ZQ7�7I��(vD�]-�]�G�d66�#�����m�x��_ז9Zv����kmW\�	�����\\\�爉�*�}�p5,�۫�g�S[N�z�Y&�F��}	U�p�
����OY�׹@8����$�<�I�u	�o�4��M���N��<Bm��{���L�a����|�eh	0�g竗Lwn|(�G������(O�$�>d�8�ƨOP�&�����'�o�N�qOz���}���{��Vs�ϫ>߹�ڻ�)�������CϿa�����g9�z�9��"�.�z��N��y�!�dԻ慒~I��8�I�t�d�=���>着�����%����I 3�\@�x~`~gr�^���������ԓ����OOS��!Xz�2u����}������=�<�Yn�s�c�>�I���:���4yI>a��o�!���5��x�	ĞO� ~g��9x�+�5�ϙ'���,��Ć�ϒi�D������S���s5���3�k������rI����I�d�>2q��$5<��m�x��C��~g�N2(f�1�?�z�a������xx�]�k���?���&*g�d��@���MM��I>d��|�q�!���{C�'����~�����0�n����I�7�ˑ7ww�'��zz�a���(�N��OȲ[�N[&��̚���B|�ٜ�m�I��ROY2N3�����'9������߿{�t�k��i>CH��I�d�;��VL<�
,��k�Y9l&e8��O��@:���!>`o�M=Bp�£�}��\���h�����u�v�}��m�m��������Cl���ré4Ɉ��k�!�J��{��:�\,֒W����O5d��M�/s������B�� B��ߺ���*3�Ѝ������cz�f�sR�C�d�f6+��y��q�%�`�W+�6���9�җ�S#JW1$;�,�p1�&|r�Ħ˃JT�S�ZǊ*$��L�&ǜnC�9��)3�����:}d<g��M���$�+?!�I=;܆�<T�yaԞ2b,��@�|��'�?"��	�̰?>G�z3�U*���ݸ����f^}�Q�Μ�?2��2L7`,�����I������N;��u��X�y�2[a���@�k�9a:�z?��K��Z~�HJ+%�G����2 $���%fk�	�!����aﴂ�2u8�,�O߹��Y&'S�-���`TcPM�}~S^�5����a�y�a=d���M>�:��	�xɣ�`���6�2M0��gR~���&�8���I�L���LAUƔ|�c_Gn|�<;��}����!�:a����VO��n~��<B|��	��w̜d���Y:�P��l���@��i:��w���;�u��緩/��W�� �>g�\z����2NSim4�~�+	��P�@�r��=a4�xì���'Y'�2c�d=�vVu}j�]f�r����Y��ݡ���P���Zw�	����2݄�����:���ß���T5��2N>���H~a�M!�}��4�M����Uԧ�	-�4~ 	>��"��ԟ�;l��~a���u?v�S�'�;�I��''~���~q'��x�d�Lg���f�y�s�����2i�3���4ɾ�d��k�N2O�ǶN2r�=�	��=x�c!���5�����?3�'��$�f![�오n�3��5���O�'�}�2>K�<Hje���V2��'�M��	�_Y9l����I�N0<C�0�u?�Hq	�3�'g�_o�k�7�����j�]aW�˲]�&��R|�������VC7������s581EE��f��9ï�h�����/l�d^���k������Ĩ�]Mn7w���=[S3/5��>���t+���8�_	R�rwR]��I�˝�}p�\��DM��!�����aXk��g'���,��B,�OY8�<2�q��$��>d�l'���N���~�q �����߹|ڻ�u��x	#�]|@���||0����a'�+Oy��qr�'�P�>I�'m��h q&���I��Q|<�������N�oo�Ѽπ�<`q�d�g���+	����l�r��2c>~;��+{�Y'��)?$�o=d��6Z�>bã��x.��N��d��{�|�u��@6��<`d�8�>g~�x�2M�~��m��@���J���q
���E��Ogh�~����\���{����O��L��4�Rx���H��~`wtx��<�3���<a���Y3��}�4d��C9aԞ>��H�r<	��b��FU�w���|�M�尟�k |��dѫ'י!�!��I���ré6�Y'�T�?d:�q7~�u'��3̲>麖j�����J���y�zb �G�9����3�v�a>�2�W����IY�P�$=퓬�gl<�	G��3����!�A�PW��ws����,�����q'�M��J��&[��C\��$�&��)4�I4ZL�'�a�$�q��	��d�����f�,u��Ue��}�χ�Ͻe{�0���ϐ�,&��Y���}�`VO1�~�T�C�IXN2~�I�=B|��Bmk���vq�s��Y�ם����ǲ~gN���i��,��m'Y8���q���ݒi�>�C�����y��Rz針� V=�d8��@�a̋{��±s5fn�B�u?p���^�)/q�9��OiwD[��>y��FUо�Q���V虇q>��b��
-�(�Eb�������^.���C�Xg�`l��qN	]��z.�9rs�D+��	��$b^T3$�\u�v=Id� ����N6?�xI|�9�u�z����'��O�uO�P=I�N�o�	�S_}�����l:�i�!�����:a�{�~d����Ǐ��k�8g{��B~@�݁�M3�oVC�dѿrq���g��:�I�=�����~@�-6r�x�������I��ϔ�����
ghM�}mf.kn5gޓ��:s��I�s�M3ąa���g��Ɂ�b�=I�}�8�	����O�;l��ì&�d>Hq6���d,��߇j���,�zφwH�~d;��$�2ɩ��C�|�'���a�d�2�������
�s$�{�l�yyDx
��2y�����*+����N>��d:}�̟̇���!ϯ��C�o2O�F�N2x����Rq��}֤� g��?p�k�Z�[���1�>k$��'Xm?06g�`q'�Y��a,��z��O�y�d����M�~֡?0�o�|�qeOQB,�'�:ɿ��s�o^���w�����u� �&��d�����m�$�c'�z��i�3�,
�~�����'�����8��1>O�
�2O��@����a,�������Ү~Ɉ�:[��?ZE�Y=��!8���d6�a8�j�m��4g'�l�_h��}�N0=f�7�d�!�LB}n�7�M:\��>�Q�lx�H�x�'��w/�?[&�I�Rm���8����!��C�x������2�@g���W�❥��cqV��>d;5�C�ORb,ٯ�'P��F�'|�'�a=��*~d��'�Rm{B|�zn���k�	�M'ى�S�+��۠��#.��v�TxM�ف)kk��̙B�ޣtz'��|�	�+�w@�|;p5�!��ζ5*����O:^��K���N\>��ls^3�Pj���j�u��X�3���7j��"q�X�%�Ǽ g����G�oF��
��}�Y��?�����|=�b�h6��u&�c���a�6�>a�
�RN[�J���Y>�M�G�Vw1u��t�;��Te����{�}���<I���d�h�N2����N'��Y<E�����2e���$:�Xh���1a��	�3!6�;���f�7����Y%g���<��z��q'�����/E'S��2V��`u��Bo�� zɖ��`x��3��RN2}�wˮ��޽Ͽ~ߜ���w�1��t�	�u�^X|�x�[���BnY�d�g�䞲u'Qd�I���܇wd�f��:���A9��"H�s��}}X��B��,
���8���'��	֠2y��u�x�a�N��O_�1��Y?{@�'Ru�������j�4�N��}�I���69NN���3>��� {�0=I�Hw��C��P�`x}I�=d�8�P������:���qY&���'d��O�2v���}�~��;�?k�a1�L��a<a���8�������?0��w�O'?~ȡ5C��u�Cɫ!�d�(�O�=�rN"�h����o�������>DxG� i��ӧ�C�Y���ש'�y��OY��I:�a�Y6�z�1I�m!Xx�2u��,̝I۾����7���;��Y&$����N>2q'-��'Y4�O?Y�3ϵ�רN$X�l���|�+&��8�=Jœ�m!����|���o�߽��>ך��&�4��!�O�jo�$��̓�d�;���<Hl��I�����$>��ϐ�d�9�Y�='��L�{�|}D��t�~1w1�)ʕ�ꫴ�ח��r��̰��pѱ�l[ݲ��w����N�ׁ�<ɾ_6�i���8=�f��j�\��݆*����\U�p/��G�1�v3#-� SQa嵽Ü���si�7�F�(4oQ9y�ܒ��xq  H�(�(
E�E���Qb��

���|s���P�#J�Y�M�|����2h�5�'̛��0�f��I���	�~"������P�G��}ʟ8��϶���so��}&�|Ɍ��'�V>�E�qQd�,�[�N�"��'�7�Z�����oRN'��'�<�{��H�݈}�>﹊ߟ@����>	&��M��:��1��%C��E�qr�'�a0�qԟ5&�� �
��a>`f��m��h�~����WU��H�c��>g�}7>g�}~p�I��捤=f�<�2I�LE�����T7;E�u&r�'��f^ |�IG޺�y��ž������_]}m������ŝBq�g4��x�g����I7��4��7�!Ԟ�b,�RIRq��N0�}E����v��in���s����i��$�|*==a+3��A:�4�Y'�v��N��z�=B�G��A�Y&�0�&�`w�Cl��|w�C�|��+��gn������#���b���� �O�q�Vtט�C\�Ӭ��{H(c'SG)"����E�q=���'��b��������#�~�0@���F�|#>3\�?J����d!��']��a��|�nRM��,�۹��躥W����\�Y%x1 ��s]����V���U6�kW�6��`vd�o����|���GdU<�Q�k���lLBJ�l̡N%�;9��2Π�e-t5�Ur��յ������h�F�V-*s̳#��]�m�� MA�9]��C���r1�}Y/{���N3��i�7C|����pH[���-��f�Ϥg��$뗛��4_i��뱵�[�7-��br��W�|�������W)�1^���;V!�����Z���]cJS�V���Պ�S�uv�$��o+��N-��K{(�GG^r�.9�Ջҭ��D��x,J�y�j/��t!�sg\�О����<Ya�u8f>-��]Ɖ��V,���.w�2͍��s��2t5n�7I�<;�k�x�<6l"�c�=�F�Vm�7ֺK�^K��H��gfq��Ԕ�fA	zƺ�@���AB�W
��vάT5�ǈs����,�݂���Bt��Q�s����Ց��񮳈N�wN!�16�&Z�'t�����[y�;:
�Д(��
f����p@��V	RM�(�u抳�N��2�d��RZ��7�wu�RU�["E"%�ۡ�R�_i)^�83m0XX{#-�r�M����z`��ڡhZ��rΜ��X=0��N���gyca>�l�
��S�xh�����˽�
n!����wD���$�I$�I$�qr�j�O�Kv�.�7�oIyu�-][R��*�Ê,��pӴ	;/.a�)��%�RA(G�d�u�nUϏhޚ��:
-�`�Y�ƺ�[�6�i����i�Eq�������ԗ|\��w~yn�`���*�F��qU��M����`�>`���H���Cqf���N�)�r3T�7B��jX�7���Y���7Hޢ�qZ��ʘP$���r��VJ4hTU�ڧ��ˉ�61��MZ;}wn�5�}�M�C'әÞ���p^h��}y9&�,2��2�l']+���K�9�g�$lHB���56'���]��!�kNQ�!�p}3�Q���KT0��xѮȑ�B��D꼊�VAK��f�vŽ���6ҮŅU��dq��emN��ij�;E_Ț뻊F��v�ax>�nI5�9�/㸣���l��F5�]�8��0*�f7C��S�%�]r���]_-j^	Q���$�n��zlnM� �
��P��r��]������ �4u)ZM��a
k8�0��z�4��F\�{�6��2	MR��	$�ZLn4�P�$��k.G$����H�q�?�?����2�b��Ř&��q.��-jP�&SW4�u�t�Q��*(�3WLª����2\�wL��F��1l)GR�T-�p���e6�˅�(�eF����hhҫg���ck�������q���L�f��7Y3,��r��02����K��)�[ZX�����isks\2.\�\�w���B�Q �5f��MD�F�T�@��飤��i��c��]��.���*R��(�WlZm��e,Q�je̬fZ,v�&Z0�.Z�*��[E�Vҕ�ܪ\�F?���+�0��L��}��,X�2�X�3r��%`�Z�e�s*8W�3�]9"�(ͥZ�E�k%UJ�hֶ��5��y�h�U��������T+m��ո������jWY����-w�91��5�&�E�nar٫p[s��\���pr��չDleƶ�۪fk4U޵�GF��}UT���k\���C�vmAɩ���*��܌L�ʉө�o�M[w�Rr���ގ�Ko�T�ar���S� x�s�$�fO�9�l���u�y�����c��N�?t��5����V�F�~��o5����^<m�pz�)U��M(�e��g�)��p|��1_6�m'֑C5���E�ט��5�c��ƫsr��PΨr"8H�r!��m�7�N�U�huUt�;����67UU[�yY�g�� o�!bK���=X�qhf^'h�3��o��.��p��4��hR������J����r�INB�FfvszFu��\�-.���q�J(Bż�[ÞkK~M_xy��b����U�V̷$o�0ߛq8+���6Z�w"u�	�r(Z�Ó�Q��]84	O \��W;J�7f9en6�w�ct�Ş�eC�����}aL��i[Ⱦ�n{:�L�RZ�;
���;Z�>k�6���t�c[+2[y��5��5�b6<+��(HH䯥^�W}�k�iU��qĲ��N���AB;X�9����r���ƴҜ%9��u%߼=� ,��֤_Th�ڞ.��!�|p�������`���y��{^<�ژ=h`J�����ϸNɚ�7*�k1Z���o:˫�mB�Ʀ!'e�Q��0:����B*���T��e�̑�w܃Ǧ\�{%�����<-+���=��92�I�Τ�!���uem�.T�4(e�k�ϻU,uz[�52�*_=����Z�q%O�
�ڛ����s�nq�Ԋ��uN�����'����봟�Iuy	����2���fsZ�$�Owܺ���˩a�Yc���'d�6�G�r)����{�u��>�i҇�ZE�N��s�9%�D��ЎVթ�AqeZ��ӓKx��3� �U�Ö=o#!2��ddt�Ѭ���no\4R:���ߓ�_lM��%Vhs��ѴP�c1�]B���ҚÆ���~$��6}�0qǵǦ`5��}V��wA�R�Y=ܜ���y���I�}�Y���D'����b��6�i��;tee.Ԗ~��3r�kouov�%���7�{���x��ڒm�<��|��Z��.y�}�(2����S[MD�BY];��N8�m�]�꯷z�}��'u���W��m6�;�6�<�aʞ�l��o����%�� L�e�a�gc�C�}��(^�d�=-�|�s,��JN�s��y)�
�±Tis"�R�Y��oZ��0Ƈ;A��Ho0�ǝ�	8�4�� �h�Z��[1���f�J������)M߰Bq��I٦���Y��"��GGe��)S�&�LQ�뼘��wNV{�]e�3���K�9������n�۔������䭆�^O���j�i��u��M#��*wU�Kv�ڹ��)X����T! U��E���<S�ۖ:"dgl�ר���x��Ru�rvX����aUt�(q�A[cX��"�h������96����۔��qq����,3M�;'tc�o�y{O�}�W����3CQ�����y.�{����w$�>��T~{�<�uk6�ZŢ�1�����U�5Ђ9���j�T���r,7��#��RN<��B�qAU����X�b_R��Qlr��cGmҮޑ�mXJ{m#
F��*�\��9P	*�r
UH�`F��N����t�)tF��aC��
s�`�p���M��n;�O��_
�"������{�52�S����jpE���U1��;{˅�u�1�[\��q
��z�:]��6��SU2�cCl�?)���,me'[��m��Ϣ����R�,F�ԩ�[2���H�a����-든�Qs#�;3�]�0�������/XU�۰���@�L�B]��a����D����	��2�M��F���P} ig�(�}���f2v�l�3D��7�1G-�-�5�����.�/o6W�� ��������-n��8+���˒Zy,�8���Ts��v$tU�39�'���s^��d�~�Y?Jҧ���v�n{��C�{�x{�u���$~#0NvE��0&�Tӵ���A��T�WJ- 2��F��Y�<�X����E�������P��nJ�^OF��r�u=��_�^Č熂F�kω��`m_TR�k*�ެO�|m����U�[�Ҽ�t�T׭=I�\��f_���P���5.�ex@�ܯqR���b�L^��$2��馽& ���3R�J�i��:g���Ohs��g$hZr;�w���`��&]Ոƻw5�ID1�*Dl��ٚCdS}X��t�.R۬J�>���ݘ,ۻw�Qޭ�����܈���4�Ϫy���ԕ2���W.���i��}���S�����o��ච*��:�ض�Ч�=�{���o�q�s�HGU'�p��hau2R��3��诧8�ݫy����M��fNޔ1�;7N��#=ݙ)/Y�aV�;ŝ�M���V�9soz����jU{;rM/E��m�K�gB~�>�op)���t�9�;}q�3ge�
A����Tr��o%�xx{� ����-�A��o�[}j�{V��mT �/sA
E˴ź�f-^�G�Nܟ�u@��մ�D�����0�ق��Hm�����v���#�ӗ�~�f=Gm�R��6��iV�݋�t���������J.
���]>��[Ú4��E]�m���Y�b��A��"=�o���O��nTx��Q6����X5�Ǳ�"�w-��8>�;&jw��v�>�0�׊�t�.�뺬��&�N���	<4Ѹ�����m�=�O1=W��\?eN���X��ء�c����ګ����%����}��j����ʌR6�W�\��i��s��T;̇���j���K��o\u�]�Z:d����{�<$^7Y��ޢ3�!��	4���ݻ�c�qN��8�k��\0���a�^:�q���n.��\y����nI�я�nr]Z�W�:m�p���x�0fi�Y��*�F��)H�M��%�pI
>TJ��R�?��}^µ���]U�+���+��y_J���n� J4���ڽ9���1o[���q�K�7�K�9�CnDd�#\�;F�Mu����d��zm*z�=ѽ^�W@.�T�������Z�./v��O�Z���}���(��20�C�SݓP�ƕ�l�V�.�@~�P�s]=P��t��VN�[���J�:]#S��3�����w�1�� ѫ��A�p����i��9������]妕�x�+���f?@c	��9�iU��Z��Z���vjaP���;�
�gsȻ�i��������b[u@����uvU+M�s�#��쥇�'`���7	��)+�z4���K(��j����2C���*���lF�
�v(4n���+�mO#���0A���V�B��c�]�w�*9��6�Onʰw��������DB��})=��l�JR�d��sٽ�d��w�mܴ��J�kL�T���n��(�v����Q[-��RM�Q��H���\�΍��6�	FR�;���A]O�'2%�!E�1�sn�jK>�����W��7p2k襇���oBB��	:<�m
eU��Oh�R��3�MW�'��b��S���g��^7|��xw���w]�o�U��E��WBn����E�w��(�]!��Ԟ��1�{Uj���ܵ[��^R�ɑMȨC:"쨾�T�-֧.�xwo��7�]^���^kh3�݉�P[��J;�wQT���Լ$C�ċ��C�{����5Wep����M�i�/'�X�SN�k��w�m4���v�ԐdO���W٪�4�.����]���ޗ�)q��TbV��7�s0���@��*�n9�R� ��wP'{���l��rTE8HI��=�Yː�ZX{�s�\64���7����[<\��Tj?Um.�Woo�1�lSܶڻO���sk��hvY���Α���L�@��
]f�MI����3_��/��������6r��K���xF��o��Ĺ/�z'���.��38��1�Y�8��~txLt�7��ΩɊc��M\�r���lؤ�zR3�Ô4�&�ij�%�Orez��t8�*~T����vR��ք��eeQ̄-��ռ}��*�t�^Ȏ.e�)Ho�5���Jt��|�����}�dh��q�=7�\�!�A�oK�&�趉��zP���Vy(�(w����m\�T:�:�)��{[��p74��h�O��X8濨����љ^�A�&�%�������4H�hP�S��k֞�j���vf]���*��^>�o.4E_1X��_ZJ+<ոt7i�F:��=�L�ֽ�%:��u<����4����ԍ�^<���݊�V��_^EF�r.�wZ�F�ð�i.�y�S��q�[�X�c��lj�g9T�dZd�J%�g1�A�@f�/7&��N.�V�5���s���jDc�1�[���y^
�GI�u������U�ԫo��
�7u%�xx{����{ɽ�Ֆ��W#Q�ՂvdW����F���I��Y��睉�շ���I8�A�@ۘ��CdW3��
�q#"��OnDVb��o�E!���l{��IQm]*�*�.v�l����'�2x�­o`u��z�¸\��O�^�g{2�W'<&O�ɴ>ڨ�\���.�g{���U	t�pp�?-.:�۾�:�܈:Y�p��4�����_N��B�E�н��⟶ғ���QV�XG��C̎�픹����g��[��⭮�p#C�:,��.�t�PQ��:���ӺRKjZ{һ���f�6<t?���[{�u���Yuʸz��A`)�4nL�<'DR��-җ�Q���jE¯V��z��[���e��ȑ�6�p;9�S̴�����L�t/�ST�'�4[����ۥ�X+H.j�mN{�N�d��r����#��6s�:����V��M���&�B>q#IY��Ƅ�X;�X��95��Y�]�ʆ�
Ȅ�m�8>[��>y�����Ǚ�^莻�`v)�l�Sn� W;�
:)�#v�n8�kmJ�\͓���t��K���ڳ
`3D��d��Yd:�3�t��$����U�B��n�5��q�:%��<�g�y617YѮ4���T�����]ٙt���y��1~r�ʬ�}鲰��\��z�� �-�t`*���o.�46#3��`��6o@ʽ�(Fdve��{i,�Y�Z4�I��sl�5�-�"��j��D��M��n����;+�j�\c�pq��{����]cA�Ǐ���Iҝ��4��0㴬���h>4��:�z��,B�������8Yk�&�K�)Bdv����݅c/�k��MY@�Ʈ�RMk�ȕ*�j�_
�9���'�2��]�	�-flC.�5@��R��|ѻ�7�m[5V�;Q]�ɕ���l\�6��Ln�.Uޞ�;#��#s\�J�<B���nY��ܸy�S#�`�9z��}acδ�I$�I$�I$�3�����UI���ԫ�����.��o��K�.���X�Q�V�޻�r4�qSF4���ޫ�f4fs����1XZ�넸�#��mĻ8�J�W\ȷ{R{zu5Hjնw�:�]Дb�n���/�ܠ��rc)Hή��n<r�n\ �h���)L�������e
��eY�Ԍ,Tޭ�u� ޭ5����/ō��'uw��3Μ-.��ށ�+Kd�M��x�V.�� +����Rt��՚�܉v;6������1�m./j�mu]�z�oXY�|���GLW:*n�n�5��Cݒ���6���)^Aje�(����&J$�k=;����v�M���d�5�:�%=�.C�H�G�yOt9�IH�\�F
oyV�YSt@ۦ�� ��,W@&�b8� ^�q?V�Z���6r��v�2�t�LY��Ҥk�P"���g��:���3.�A����R甎�=�ɦ�&���{�5��D�K�9��ȡP�J��٤��'�ܒE�9����|�nIfG$����аr�]`���¹�ګ��ֶ�ģ�m5Q�ʊ	jӔ�+B�QPSMQ�-(����e�B�j ��,�e�(�֬��F�q���J�hV-B�R��*�chڋm+imV�R�j"��P�V�����j[h�VU�ʘٍ���=J�VDJ�j5�����D��mQ�ھ\r���))iR�*-j�kf�kmY��pb�����T�q̹n̰���j]���(�-��.[.U0�k1��+EJ��1���+Yi�+��*�Kr�9F�T*.RxⱆZ:J+���.Z�R�q1J����ѭbZy�`�Z֬`��E���.��_�X�����fkۃ���~��;�7�Nζ�K�8U�B��e;f�B�H����N��ܩ�s����'8emr�K>�������Z�a��Q�7����#�LF�xU�=%��	�Y55R�\G;��e1����C)��� v:��'����툝˺.�;����+x<k������ޔ��f��b��N|�{3gVv<��r���܁����)��\���5#��#�4��䧐��̋��.��s�Ys-��	C$
hk�{Z�{gs�9��XKU�>�w@7�AbqA�O�۟FO
�c�<�nx][Jν�ވˑM��k�toVµ���P[P6�2*Ú���IԎ�S�R�B�"�u�K���������	l�n����$���5"��#�qP���z�Y�}.r�|7z�9��ފ��:}oK/ӂ��םՋ�t��v3g���5���aK&�OC�5����R�-Dw;KC�ky��}��OM�w�{���ΟQ\�j�X����!�Cw2�	{��Q���K,�u�OU齓zQ�A��mQk&<ѕ&�]���.�(ɪ2U�m��3���V��@�Cn���R�+U9\�]�l���]O5 U��)=�$����mj�{��*����˷�lR�p/ɛ~�Ìz:���TR*ҝ���D�n���O�M*k�nS���!
xa,-�v�g��e7�O/ؿ*��y��ge�Xi�!)�B�±[`��0Z�wݼ�*p�`�N<�X�!��	��Ѹ2f�c����Ѯ5���R��M*W)��)�!	A�b�N���f	��Ē}�ۧ������Į}��X�gk8�٪�M>Cw��V�-+��:*G^"�Uo�[��<1uf˕��o��r�j�m[���U/浻r�nג�NM7yQ̦u>��S��+����V�5�>\������Ĵ�h���k�[��랷�[���9�O�[fE��@w9�N<n�_8������>��G�<$����p�f�:`d,J8��s���/������=��̙�=]vz+�vF�q��uٺ�C�d����o��GC������F����������܇��H��=B5Mp�L��(�t���V����I�]�w���ڵ�\فy0���>��K�W�ڬJ�٬퉗&�^r�CqUU���ױ�BAH#����i�S�9��&햶^P�zz�;��䮊`\�H����:tb�J�w�PO5cꔆ�{q��d�C���s�z�]���.��4́��|���K��t�b�gujq��-T3�����U�n+fӘ�l)��
:y:�74�*#�c<�]�ƕOS�7K�/�MŌ�O Y�;��%Q�W������xZE� `�1�C57��!�n��-�9�Ml�X���d�s0�<+���1�7�:V0C�`���޼3�-r���O|7�>�_o���FhO��˧�6�È�,S����ILm�A���x5�W�N��G*�Ce֬n!tEA7E[��[��ʔI�-7T���0q���W<~W������ε��f�U8�|���15��^qf�T���3T%��ͼRM��*`'K�ȿ�}^��㚳��9˫�}q�����i;8���0з���1Z�����H�-J[����������17I���s<-=��.oύ�����,����)O�vU��x����9�^��,�>q��2/�nA�n�a��c���c���lb�a��QV$��W��sB}�z�f�l��o�2;��gԟV$g5ڣ�v=��eS��V�7/���m�GfY<*1Ȥ6k��/+G3C&�:�R�ݗ^���J�j��_�[r
�����6ϫ��q�[����2/��}��nb�tpP�B--�8�-���u���� �7�z�)VJ��p"yTR[P��.��|�b�o�Y�}�E�X���<�e����6��d×{�O�-]f�D�9)�����v"��V��ڗ�v�+��zƌb�<���M�s���L)���i)�f�kS�'��{�n��5�Mժz�m+}e�'�t�.����iC +44�6oV��sybRG�������O^6��#������!%gX��QM��mF˼}fk'2o����/Wmv�`��Ġ���g�	ę���}Z��vΩ�++>}9�S��2#���?w���.���4X����������lɇ�\sD�0���YpZg<���;m����m��QQ����
��C�������F����G�D��}�W+4y��ע�z�7�r�z��[��S�Y�=b����\�3ދ��q��2GuS�Ƕ���2�5��z��J=�y����h���--ۖ��C�Y*�73�Pޞ+��[�S�f��=
����w�]��<�PBl�7��Q���>�ܶ��&�fO	����OM���mybp�0!�r8+�)m���U7�E�xf�ا��좦�NrA�~�v�>]�Pw�G'��B���;1��҈�H#�M"�R'}��5�λvM�v�z�uG��XȮ���:���qw�v՛���-1i5�#�BR�P̾i`E鰫���ˣ��8��^�D))�ĵ%��=�ym��R��q�?	���q�\��[�];��|�v)PZ�7�ү'wP�u"�@�����|g���ﺢN':_�j���f�X�]�֔�
�=��/z9WGg��+]n36�I��NL���UN__;��R�W{<+}oy<~�<=-����/�K/ydإ��7��8a=zltQ��r�DZ�f�3�s˹�}zoJ�u&��'qS=�=(���^i���?qΞ/��f�/d_L��3�ݗ8)��^�̄!V淾�3}��P�=��5�eH��(�!Kcw��;����P]������I� `�Us�`*��6�X�%S8�N&r���{��/���z��\ӥ]r�
'kL�^m�p�j��>�� 6��c�f�	0��rx2��N������m!���T���q�c�3{S�s3���#t��C6�WjK�� ����Z���f�=C�縔�L˔�B�Z$��Ϋ����L^L�ڬ�s��{�O�r;�����Ϳ5�sa��:��r{*x�y�ُD^e�@�J�o[Ez�s�o)뼴��,,S��r�����/1�j�y�S"�ٮbE�dU��|�-��|�K�̻D�����|ʹ������F�� Rg�bF@�K��)��gQg�9�hOS��!��ۣ����B5�|��v�;��V�nɚT�rTe3�p��hg�Lj��[i������i�y�TV=ԑ������-5�RW�4�y`h�f@;�*�����9��69��7N%�ז��i���sk�g1���0�w�Su��{��ٌ��zd�Y\�k.�O�rg��r����&�s��,g�Q�wJ��7�{�i[*d�yyPm<g�D��r�����";���Xm�f�*y��8�Z���.*�>T�ʊ��;r����tc��ԏ��V��u�;A�J�Dw�ʷ��u$e��^��}�{��b�����'�bC�OmQq"�zʪl��X����ɋ�طRûXz�i��r1�0S��͂ ���W��.�b@��o!��/���~���}�)G�1���&b��X�ʔ�W�S��mu���D��mr�%E?)�B��'Ym�1Y�����Vg�����#���.dƨvUoc*�t���̐�Y;^�[��A
���7���&�f//L�n�_�O C�O>���_+�R�9���]K��<w�h5!�6�}���Y1���=B�^]����#����e���=]jUcWK͚��2��h�=����rθ�W�`�v�,�.4�Q��S�4-����q��ˊu��p'K�̷uY��Y��󜘧r�:*6�p�q�6�b|�4L����$��ѧ�����'��Gڼ��&x/:\3ԩh��Eu�
UO�V��/)GW�^쬇��,A�7qQ�߰&1�r*�����r��EeͮBӚ��f��pU���U��S����R�e������Cn9�@l�=��Ҩ��4�Q��BJ��n.�郩!�>x�����zL��q���>����3��x�`b�:a�Jlʲ
���;��˝#��R#A.a륽1�^�ev./i�c������8��!�np��|���q[�
��W�������/v`�}*8+�y�\�x��PZ89��`ۦ�J5�Ս�M��k�{â��]>�M)�]���Hu�xϡN�^#��ib�(0�j�ҹA»�U�8�	�i���ڭ��}B�E��o���,�0�M"�!�+csnh������7���y�����x�2��,
�>t"�Vֿ҄���l�vxV�U�B=��~���9�(�U��='Ǽ���x�Es�7�#TD=~�ȇ	�X.m����D��wJ��!_w�Uf��t��v'����/.���Vt��������xz6*���0gշH�y4��ޡL@�/S&�w��ȓ*9%N�#�v:9bIFr��_c�a�=)*�]
ax��aC�k�WUL�eE�+0�[r7ȅ�F� ��:^R��k��1�e�҃�:���*%��>tL���-���d�]�Q�x���r���RY<�՝����YGB������]"h�ޥ��j�����V�S��7��$�����,����I΂��w?I�1U�@M�,�"Nڑ�2��K(ܔ\c��ϡ9��q'�9.�7Բm�3�����_{���S�ͳ�fF����G�p��v�9u;{�OC
��R5ƛ|��=��r��f�X������=-g<�>^�˫ݙ�{�Ұ��K��Hǭ����r�y�H�
�7�ƚGdlV��jy��=�㫢�aג���R���f�6,�=��)�k�Y��S���x�N��r�x�8OF�2g�6�Q�>�w�g+C<�C�'��bMܓG |��;���`8}D�+M`�*]@��t��n����~˃E*7�ۭ��e8߸��f-�-oRȣ��T°:$^����CM�R�Zx/����r�����;eo$����M��)*g*2�U��ׁu�(Q�h�G�0�:= ��4,ћo.��C�=W�������J�+�8):�"��0Y1��])�j�7"V7}9X�y�"�ށ�aCq�$����ΰ��GV�a�k/�X$�N���*�l��A�Xy��4�^<��«����S��ߚ��ZU���;QT�`��uo�<q�Q��<�:F�n��6t�u�j�q^���؃;]�6��(T@b��,�U�I�G��Y{���!< �́W4R��z�k;]\��Id��KC#aR3�gI'cխ�e�b��[�6n]��6�zu�(&:�I}��r���ski��L�ѭ���"ቬB(��WԾ�-�����!��
��@%���V�F��2w$��eM)��C����ֻ��*8�<��}q�8�}����w��{٬�)#u'R�j�o!�^G����i��oU�:ݕ������w^	0mV�C1�#���a����Zz�r"N�!9�p9B+�۫u��D1.�W��|,�c�mE�2��+	�{�e�-R�Z���e��ý~��`�xy��;�'�� 4�IԆ̈́���waȞ�wx����t0y0�d������ų��E��������R=��#�OM�O����	�P#h�a}�@��ԹR�R�d���4������:�6ud�	�=�.t��2�,�J�f�%wJ����ٶ�����s�Va��Fft�_E�I$�I$�I$�N��ĮJ�*u�j���MG��U��{ۗӶ��y�a=nj�R��.�RZN��A�O8Q|vgP<:4�޺�չ����:ȜC��n������� l#4���j�h�"w�)X��w���V|k�+��Fn�SP�gŬ�5|1u��P�S3�Փ���:#i��U|_\�kF��:�	]�8��ˤʘ4b�؆�y)M�7��܌�yJ�h��u?�iLGp�kF�q��9);{�2ɥ����z�t���A��J`��O���:����m%S�1f�0q��1lIۦ���{�V��#��^̥ԵIqh�s�������62��a��m�(����ђ͠�6����ݭ��6)�v�Y4-%�ٔ��m^�,����;R��N��K�f���/UZ�b�ᜎ�����b����X��nZ'����E-��dO���c��D�+Y�h;R��]�Y�;�d�,� (I)�>�n!7L-8w�+�ں���S�.ͮ<�88�wt��O�b����cF��u+����`p$��r���NVKA����o.^*��٨��'�$�N&9�܎I�>N7�3"�}��~����e)m���ՔF�KUm�J��
�����
Z�F�m����f��PQ�+YX�R�r���=��%U�Z�6���[KX#-�E��f�Z��iY��V��V���U�Z�V��+�eKmDA2�[Kj*UF�֬AKkh-Q�)Ker؆���Z�-,����Z�YXZ6U�J�%-mZT�R�U����)��1��\�Ep���J�b�(�ʂ�j0m��{p�b�IK[�S�R��
E��U��J�emB�ƭ��Lɍ��J+���T���[(%2ܩF�Z�1��~J��5��4��fJ�(�e\��W�(��)uLK�pY���|��J#D,��+ET2�B�j�ms%ťV,Kh����T�����V1F
���"�#�f���?}�知�\6����^�$�֪.��k�na���f �cW`�f	qT
D%����Ԑ�*���IN+��{���Pb?�%��Cc����u�����<�ѯ5/bn�3]�.�u������Z����;�E/� �cB���ϭ ��yɊ@.E�;{7;2�#���_3V�I{�r�{���h�.���%R��o���޲o�`{X�^O+�9�
�����Y@�@�}Z�pt����*��ja�]��㼤[�ͮjkl�c���\�^>K�r��0�G�
�2���F���r��fN�CSu��A��h�kg^�3ڝ���2�(�/�����j��;bv����9�9K"��/  w#O2�[�-��o#B�Y"�8v�E�A�d�}m�bm<�A��UCc�[�G�y�W�E>z����:�p��{*e�q��~P�h�K:��'zׇ�uf�n�n�le6,	�mw��������}����B�Z��*U�N�#8���8�<6���o����bF4��8�.�,(��)ԋ�x�ٕ!�9=�yV�nS{��y������:�m�@9�,s������U�5���t��z�f��j�9j�G�}6�fL�0g�8tQ[7�y!{�����[�r��{�и�}ϞT����H����ɣ�Q�z}�`,�Ѻ�*�V��sC���4*��7��D���EtP�#6��$Z}a�8e����TAf��@ ��sQ�������~.��w�z�L�R�WM�B�.���8�!U���'�#kH�m;����W"}J�e�
�|;i�����k�OݲR�/B�-�
���gn����K�������)�h��ʋ+G#>�1@m+F;4V����_1��Ok��嫉}IW=����|n����À�N���j������ُz� �+�l����(���1HD�\&��3�}�Av�W�z���N��w��}�#�PG��p�g�+����b#��j�_�l��{����u����X�u{�;��_�Aq>��i9ȊÔ��XT4}�uzIw�u��=Y�<�1�FR�t�f�c Q[�hS��0FIk/��
R�ɏ��}:�Y:�}S�Ww�	<��9���P�6����F��5t��6�ӳ��OQwq��^�Z�\�|s���&���3��FZ��Ѽ�������}���+�?J�R�N��o����=��/� x�mr6҂i�<>��U~���o���5�{��Գ�靹��`���~e�s�{�+��J>
|eP�ES���PҲ]�y��U�=��MH� ���On�Y�~�<
z;�Y����F#uAХ�<�Z���|����~�.?fe�tCqբQr���=�=�S2�Vx=��ܼ�v�s\q�W#�wwn�F�,�C#X�y�H���G S/b�O���bDp6���¹���m��YV��bdt�����G������kDVĻ��%{J킍���ca_)Ŏ�Ȏ�./�Yf�7N�C�k!�fn2�q+�Wo<ɮ�=��*W�ЕK�L��ߍv}Դ*<�q3���A���zȧA�<b[|<�e�ؤfB�xrW�oU��8��`rt����%O�����3ۉ,���Y$����Jr�h~����(w2�x�U��@Viۦ�j����/���*��Z5f��o����o�{$���.��ni�N��j_E`�űP�V�nha��S�Z�[q���*أϮN�H2"�`��m-�+��2��Y|�ܖ�쥅=�D�B�}���-q9��ꯨ���o&Ihr��H��>��Q��X�9�����0y�����6���v��)�?-�O��&������U�C��J�����\<|&�x�x�^0`�J,R�H5�A
�G�W[~=�%���& U�OL,��R-nBO�{�c:P�ۡ��E��4���n+�h�~8Ya@b�E�����1Wל�;�҈�7�逕�eKQe�̏0V>U-xuK�;B\�-i+�{q޵�w]r��U��sV�0l
6Wj�^{�FJ�U�'Ⅳp�VX�"�q�9�]��iO�ˋ
��
F��=�v+�X9��o�K����V���nU���c������md�b�F�J8��uc�<�-��C��l��[���o��
UHS0���(Dqgm	O�
�Q��e�PV�U���u��X��V���Oj7���P�r'L�X:�Z89��J^\K�4Ƈ5l>���D��R��B�*amkX��k�q��1� �G����H6��yO��zx�����O
�7_��ۓ�GO8��t*��	9��족%.mBtn�P���}H� fP�r�5iC�\v�;t��6PC���.�x{��s��/�,O�*��7[�`��R�
��>-|'%���>�kD��yq�����ߩ���Q϶I�_W�GtL�]�^���t+E�(��xF�}�r���:���yS&�c���s��JċJ�ڌ��
�r�~B�M�2����3�s��D���:�,�_C�.�*�����W�'ZdX�H�C&a� <7�]<�t�.ɧ�tT	=�4����1����ΰ�G�.�Wj�(��J��K��On'6�Vd
�����V φ�&xK��2��r�bÛPr��1]{�c��C��f���t��B�"��L�ȮR"�E�d��X�P�뷷oVr�p��Eg0��(����
�]�~�-V�u��X8:�\/�Un*|YkFʇb��*��ϵ�ˬ̈́E<�.}�N�\|0����V�P[V���/�d�Qx��9ͮg���P�(f7�%���=���'y^W��{�1��·�>�m�.[P@�������,ӧ7�^{zy��^�fRɵkH��o�'V ��0�]"��td0[�k�Z}���M9����$�s��*^�����f��z�P�ͺ�Q�z�7�r:່Ueñ�!�{��5U��WUGLq�*x���+$ k�y�����=u���l܌��/Ǻ1�K��5�z����7�cyz����lv�+N�?�箱���Ki+:��Θ�f^�2�V#��!�B��x>:���x��>%}1Վ��n.oz^'�iⵌ�1� WD�\��*U�Z��t�q�:2r�x{<w�������Į�~��S������]�%�`��Zʔ4Rms�5�V:��ٸ�b�s�*�f��c�p/�����ŉMޙz��Dh!��7�rv]E���^����������Ε��ʫ�]�̊}ʚ<�l*W����z����}���F�_-X8��A|qhb��Ѩ,���P�u������j\�e�pN9�W�l�&uU�8J�yp\g�y�S��TX�[�|�g���y��I��}�P�]7ǈ���DR��@�X8N��j>+ƌ�o��#v�
0iv_����o{WK�1̴2�S���i׹Y�����>��S��
�e=�&ft��A��!G2qp�N�� ��w�jt1�:����@�8]j-��fs[%��9�vN\G�B	a�mt���2���]�w����-Z��Bv��r7�i��N�5jY�k��Z�c B$:&�B��3�Dn^ˊ��е��lRx��� 8p�{�ɕ�
�-x|kb#��)���+��q����Y�G�p'��ԯ[u�0�=SU�灉�7k�p��^}bðr���e��:��}�v������-��O�7�6���һЫN��^��-��un�Of;�#��>�#4G]��(���D�����xz�*�}��k̬�~_!9J筤{WJ�m*{Ӂ�0k��,�Y�O�h���.��Io�(�ٗ�˪/���b}�r���<�8�Ze�ٺ�QP��[u�#��Ь�U��.�Ȼ���L��4X�=CzQǁ�.�uX}�f�],��3�2z0צ%I�s�xפ��'nɲ� i����T��Q��]�+ѽH�S/b����q����#�`��:���J��⃨����`<�So�|n5����%�r�ya�m�Չ��A*���hU��d2����R�;�h�k3���ٶ���";���.��77��$M��KF���k��Pokte_.3����w%��{wh�x�(1�ǒ��IN����!��wu%���-.��w�FDfQ�2��,0.��H7N3�j���ټ���0ӝ��J]iy~L4ˈ���bxϡN�p��
ɪ
 ����U��!s�Ͻq	^%W�T�Ld"~��	؁"V���wg���O��-�)vA,�T8�Z�x����>�����MY�`��K�.r\�R���n���;Ѥ?eZ�`
3�ue������x�E���)3�Kj��w���i�=С܍2Y,��2� �΅^�~2��koʑ7[�B��a�ќ3�5�t���hEe��x=��x,(�HRV-?5��i�y�%��#S'
кƼ�10�B1�z�;�Z���2���]�8g��=�eЦ~~��8<=�Ona�$+77�؄2�슰�a�^iV�KQa���M�vZ�eq�������>�����ۜ���q�}4�G��^�PX������ߵ�0�"%��R5�=*硳s8:M�Y��7��VT�:���5��%g_@�p={����i��j٨ql[��o����*�M���k'>j��B�JZ]Y����:+���ܸ�N���3M�<�:���?�����.E�y	DOʩ�(͞66P��c�+�w�`أ��)5a��{+NL�^\<<N�bM����?R��=B���9�5�Q��u�8�Ab����
���z�z�А�.LuD�pu=J���]����{)�kg�ja{�T!��v��ެ�5Oȹ
F��%G;�Ä��\�uf���j�}�H9��wvzx��"Ա�wꗄ[�Y��k�8�^�:	=��t#޵T��\ڇ[�R��ٚ^p������$0�s�'�Jţ��J�}�?]
o��w���cx������Ql��#u�R�=�ԥ;��3s��U9W��!B��當��J^v��l��0�F���B�Q����ʰ=I���mw�M������r�#�9^<��z�Y��@{n�;b[�r���VK�k½(y���i�n&L�oa^p��R��5�N�<6�_+����L�c���~����9~u�`����(�0�ʹ���F��^&��l�U�.3�:�M�]�{r2�2NMØ6G� ���=��yW�z�B���`zd�y��Yi��p��ܯ��'G�vY�a2rVb�YT����re�G*��f��z�کx��T��B���*���b�Ɵ1��#��@��NI�P�'�C<�q�3ܤD����%���Ĺ��l�ko����Y��jY$SAD�� ���N&r��Us��m{����}�3�<:�ڀ���X��>K�*��� �Dp�ls�3�mY|�m�u�1��W�3&B"oj��1G��%�l��=�߇4/L�/йG�:��m��iw��
cL��"*�/$ hdi�l*�q��ȂbzkK���Ԗ�j����C� 
���*�ѫBx�ۦ��1Qj:"�8��TE1\��1ڳ6�^Ŗ:����+�q鸟��|"���u-�/ҫ���٪R�
j��S��FڔU��V(�:ląε��J�B��Fq��Z<�=�.�h.9��%�k�7����WY�؀��rˊ��yr� 	W[V�� �o��9Si�\��
�c�P��:��v����M��s�^��UY�&w���7���~�4m�q�*�tV�������Z��l�e���s+q������o:pUsT�[��,����@��֭T��gCzʬ�ĀZT$�}�N�`�)��a�3@�U���Қb�W|)����B��;�9y���Y1V�x�\*5�2^�v�Xn�4i��X^�W�+�i�����+B��)e#��}�f��F����|rA[Ȃ�g!q<�ʏun1�
�a3�k�BG!�Y��+4���OKE`���N���{c��7����ni�q�!�i��*[������KQ��ٜȱ)wE���XظbōܹSl����y����л�y躓��Vf�.U�Z����HҲ�u`d�/[��@�Du��aj��d�nt�vG�yk�v%�$�0Q�1�p^�Y>B�Q`B�m��1e�}u���r����v��y��V˭�z�Z+fܙ�k{�@����\A��[��kzq��YB��p��*٬����8��Ӿ�
�ۜ֭�y7\S(��5�$��ģ���#�E�a�mA/�w���[�S�ږ(�Gl���\�;V��,.�Y�	�ʉ%�}9��7�apfJ9��ļ�Иr�1ek���J<�J�r�h�y�[�1�F�h�Y�ګk�+/,���u8��I$�I$�I9DEdR�v�(��d�ͭ�w8���"�Y�k?n۱�V7e��@���7��J��92�'m�h �
F�{YLѬV�;{}9~1%[w�D���{ԩE!g�j�޼�� XM�	����!Օx���Y��t���.0��6az��^�4B��'����ްe��E�m�xDH�m؉]�ۻHu�\�KN�w�5G��d�ʭS�wraz�f��v��qM�w�m�c7T��Rm{Y�h�T⒨Zϭ���L��z\�]rf�/玤�eb���s�����u�A��!�o
ۣ�ɪ�-l�OI9y|����p���GveU# n�u�Ո���`����ob��h�����p��/z)h��{[yx�����M���9���1��;����q��XbM��'�����kR�ڳQr�{^�QCo�#-|{]Dͬ0�*�
�MO����Y)���n����chM�q��r��������F��Ȩ �m8f��;�D�ʾr��}�79�1f��BĜ֙�_�O�ҕ�SA[�ѝ+١z�;W(@_Y�0�q��$�����w�խ%�D�헳/�έ��g+�/zԞSw�U�Av������܊�x�l*tIƓNI�$<܎H�|�j9fE$�a���� �Q��G(Z���5�AQF����e�g�TPEA1������������t1F+S-��"�D\�CIE�+Q�D��*J�Ҟ�y���̣�a����"�mEb��s*(�kP�؋Z�QUA��)mQJ�Y�UPM�V�b5��j,�E�(��mE��>e0A5���3�)��#m��t��cYSt��V��eelU)eQ�(��AX���Z���଩V�H0TEE�[kQE-�m�U+XV��ƪ��h������խm�ܨ��P`��-m�,��TD�t�!�Z�mVe�R���*.�DF�m�6yj(�.%�e�FE�ԬʔQZV��T��(*�-iR6��-���2�1J��ZQ+Q�]``
�t(UV�֪�4�4�? c9 �]0a]��S��.��hV�|�҆n⾏�^e�7��s.�Nhi�KM�ɝ]�-� ��uf��N�t��DQ&b`5���F�]�ۮ`S�Tє�d3q�W:m�MLv%�`��3��D(EF�_ ����[>)�,�.��T]��&��X���C�Vª|�׉u�R�u�:J^X���?��Ъ\`��/m�Nه�Y���D
��x�OL8�NDH��mU/tc}[�x���{ wJ��뀋���
�y��L�,� �Hu�od+8w;V�ź��"�H�ں���_rʏP��w�}��-x}����,������SfG5��Nt5���Ps��iM8Ut�� �C�Ԛ)�DP|�w�x����(o{sT ��PzRPg�xXʷ��0�Q�0W�S��ӷ]�N�Y����Ǿ	�@횦�eh�g�fD�Yg�70��,�cd2LN:[�N2yZ�g��oR?7�O.��Az�t�C����~XO.����T�vԗ%h���E9�d����ʴ�V��*�2�Ɵnni\8��m�і�d��4<T:����׼�2m_U�����Mۭ]�+1���rvڛ�ɟs*�p<��m�����w*hXK���UW�_�*\z��Vf�Օ��.,c�K�f�yq�x�Ga������G��Ǹ���^g:�JS��t����nQi�a�{XRR�GX�=j�����m[�2��/��A�%��S0:�ϩP�7<Et��臑X�L&�5j���w�����*7@i�괫�"�JGp����C~heeS����g�����c��+����ADgG|�p2!N��Y�|�:%>k!��\ �4�3����O1�n�{��[XZ��-)�#�!�M�HU�Q�S�D\)f�f�(���'���\��΂QaC-�s]鬵B�C®��y�!���v=��D�J�|�Y�ByR�7b�%��~W���=�҅���xG΂4Ej� 5��������/y�g����ұ�½L�mY���҉x�83�wB�~��,��]z7���{�	����,�'��G��������yQ%f��uw�Ǥ40��enbvL6r�ܕ"�gD���<�l~�7?h�6<��{�+l9S̷)�*KD}�Z�qskw�^�w��]�bE�H&#���nj���S6VQ��hyO:OP虭D~]��ú��Dz�\���<o�2��6s��V\u�c�R]��C�I��`��Rр�Yap�T�_b�G��G}q.��`��[Uc����n�s������#eh$_�^����K�"��n3ݓE�vsf�j+��Jks
8Rl�c���\�T�SF��@M�,�+M�1�CY+F�
m�̒t���x,�Sſ.�q|��8N\U�H�A,轚q#�25����aL�P�w3���3y�%XZ��0���Sؠ;�[�}�7�˚�����P�W���4:�(�Ӯ)��ދ��U�W-m,�ջ����P�'
D����T�����������K�9;���Jp�6�3���~v�h�Uʰѱ���tp�<_	�ī4ƇzI-���~��oM�ش�tw��b����uf���c�7��^�}�gd�}WV���L�z�A^�5�;,[�d)��e�ţ�J����Z��B��|-�`U(�2#~��o(W_"�QХ�Z�]��r�*^<`�3Cd����ṁ|��;�YTu��\ve�Sy}r�s9��o;�h��(�W�����,�xx-��ԙܩ����F��B�p�ā.C�u���ThjhȠ�3��#�Mt��4�au]ȂC6k	d���U��g��5��R|j{�M�چS�8G�����柒\,.؊��F��k��g�D�c}k��yV�Z�.�l�Q1�c��7J@�ʣbT2G����3��Z��Ƈ���vZq�q3���ճr{���=w�+ �R�q!�oܼK����N��E<t8+��=ǎ��M��W6����*�=N�f�C��S�@�� ��îc�J0f�'YA�c��'b}��ك�դ���X���	�`�y�V�G�-�m�ꉕ����B�Od�WjC"�g��n�eϻ��E��9�n����$��הF`����Y�U~�e��n���T������|1T�2�a�j�*�[Ս��ʔ���7άW:�T]��X�Դ9���> Ac����/�\�=��OK���"�o�yfb�(s�~���%�p<�F7:��	�!�&3/gs���L`��ݬ��N����������n�FJ�qwn��3),�`��2���Yvc�����[��"o!�	R�ۅ)#�W����m�s.h��I`�R����+�}ra���Bx���#�G9�,�-�d��ߨV��ðG/B�$r�U7�J�UB����+��(��"��{�ӲkK�.!��8�ƹf͇�K{����:����<"��^Tz���淎�������Pq!(��ۋ��r�F�{b�J����\bފJr9�7��L<�(����DFdDp���kC^�����k����w:��>��k��,��r�x�A`��	AY<li���p�vׇJjY#G���pN=VS;*�օj����I�]*�T|�Iu�R�~����q�?-��;]�Bh���˟N`�l��R�Y�`�RȀkҥ��"B�Q�OL8�r �������=��ڝ�=%��p*���~��o?�� _�x��k�!�m��ov���sQPn�C�:d:�*,����x�x�N�"�3�b��O�|�LꞧY�&���aW9�V��V�T�y�;�����=Yp�ݝx+�n��L؆�z<м燒۬�gZw�/jd���a���{�i��ˬ��Ϋ�xa���ʆP���7Z��]�u���M�U��bb�|&l�^	�?�xe��z�O��B������������MɅh����jbfˠ��yN����2(�+dYT''2sw��$��Xy.[���_t��V�Cb3=�U��\��������:�K^���2�jH{�{�U�6��;����;��ՠ�C��;����h��A��{�HzZ�e�M��n���w��ˋ�k�f�7O#�>u�m�a�"nd�F�P�':�'2a���H�Aݲ��O �uVÚ6�{e\	���<7�]��
NGS�FbL��"�@Ӆ3�#C�o�D��z��+�h�k�]#�^{yy�wP��ʎ�8=V�ySHV���=<��m�!�u�kuӒ�<Lm���/�u\Dv �	Sip�@q��Ap�u9�tJ6SY�]:�:z5���L�-��*��GL<ˈ�c�q�
t���)f��K=F3h�ĺ�#P�гP�t��׆�&D<���ڸ�sJ�l�Һ�ȷ�V�u����޼n�.�J�ΰ���{�
��I|4�*yķ2�{�Ȁ��v݃�w}LJ]p�t󚣧q�\.bz#x�<jE�əJYɫ$�2�U�j��G	�S��`�}uѬzd�r�q�����Gg���n�c��O϶�&�?Z�P"��Ƞ�ʓ��WW�S��d�KX]�T"·g�Տ]k~�҅�)�Ԩ�u�؝�y��c�>�*,~���gEg��V@���ug~�����'���l��p<E-���ogqy�xb���J��Mh!t�FÉq^�38~����y=4뾫�����$�5���˴��g���b�
A�Š�O��=i��MQ/�6��p'�A��o��d�C���P������{�!t�֛��ӳb�4�����j���u)ˬ�҃�a���q�I����Ev�{�(�p�>�����\6vq���/U���8���,��X]yu;�{"����W9�X���W��Dt�נ�<����#h]RQ��l��6\�##o�`����{,E֪d�C�8;�\��U�p�D�[�R&���=p�Y<�{\-S�z}� ��r��2��6A�A}��l�勎���.�0�wY�>�q�n��d�r�M�{���	�i�&+�L{�7/s�VN�ǲ�⠽�"�)"ٸ^���nq7v��d�{�/i��������WcM#�+ӳE�x	�Uu�c;�ݜ�%�%݄d��y�{����e��[3�:8�"�A]ZY�՘��݃��.�:SZ]����|yU�=Qb놣�"yS���]��.��uj�]�~� ��$�P����2-�+Q�<��Yb:�d(w�dQJ&a/tI3�^��#�<��B���C5*z�Noj2��	E[�o��3&�!�y�A�T��`��̋��s�
�V�Bͧ�j� ��O��`�=Zt��F�I�Di��4�[]wŶ���<�oi%�p/xkJذ����w~ˠ1�l����B���ΰ����u�f��r�˔'7���6�vD�J0Xa/]Fa�:�� ��mgS���w+5�x��9P����B��"�j 4׼�K���.���|�K.��+�ks��R�%�g0uz���j�:��=!� %,�)�7&(s� v^!H��3����7�<�&��{aǧ`�Y�W��������"�4g�Vս�9�oR ���}�����(N���m��P�V:�S��5��H<�M9 �7�R�����]�6�����+FVR�Ig��uVv�N*;f>�FW�P�b�,�^�%O���E��g	^�P� Բ6��H��߫��S>X6X#���<1w��|wk�t.���*��N������x�:��p< ��]md>��7<�)�^�O묠���8�C��ր5�����ڹ=3:f��Ui�β�;6=�o�V1���< RR����z��Jt��	��a�j�~��#'=�e�ӎ�[$Z>K��Դ� �u�/}��w^���6)�_�xi/1T0nk��t*�QJ�U�J�}��߉�7�7�)�Qf�f�>�8�����s��	^YX�� 3=�.��%��w\�:馏J�&��is]4:Ī⎨��^���HO�kn���{��p(�"x��ZE���C�][��d�h=�j쩗�Q�QuI�(��+��u��CmV���]*�m*f~^���Լ�q�|�8�1l�t�����=�W��+^EA[�m�9�m��{�W[O�	�����XS�.���/�؏����Umm�h8ZwSq41f�J]m�̵j]�F�gkd�&M���<��(tZ�ĉ�6�b�K���lZ�tݘ�4~9JE�bM�u%HQ�#�'���t:H��G�z�w�ۛ��4_��|�Z�xQ�}�R��z��4��k_���^�ũyɄ�B:�^�;lC*�3�#e���l��J,�!��U�pDT�����t�U=Ip�4c�¼�.7��,�Q�Ç�p���vO�cק䣧n���{��1�`�8z"�`Q�Ni���A�;.R��^S^��~R�o,i/3[l�9���vE1�Ơؔ�~V�`>>ez��+�}���D�8Aio���+�`�Ry����1�'Y��W��*�]��,�s�FT�r�T����s�SZx0�$Ϻ(���V5t��O��.�*�,�ƑJ=�!���rm��j�XM�sΘ668���e�^��θuS^՗�N�=B��F��k	䗭��y#��ڊ,�+�7�TEoK8�Αng�������������)������-��6-�7�
�ɇP"�j�v�v�W�'�q,����e�:Š�C�e��b YX�X�Q{�*U�k�{S�n��ht�p�
���ŜK��.��]���������8nN4�h���u:��u���h\N����d�d�A�m̺�����xz��&vW7v�v�M�ڔ�n��ʶU�i���Eu�݌w#F����p� �l�v�2캳�򥂯Fg��0,쩿\	Hq[�s/o�t���p3l�"�L��P1�2�d2�듳�tr��u*�@�t��9��Z׽��j�jȺuʜ�2�kS�^Q��C�<;�̄�IU�J�t�b*�oh���7'������qNu|u,C�Xfw4{�1͊�2�k"�f�R�wA=�;g%��3�2����X�D��z��ʊ��Gu��	�w�6u*�ź6�n��ۓ;�*$ʰW'.�Z7}��ҋ�r'o��$Q�X�G(�Y�sn\�Ɂ�t��V���s����5�s�4�� �8C��fn��ɽP$�JRPܸ�u5���^��D-w�V��S��h�Eu >Z�s�Ba`h��R�ley��5��3Snu�9:�[]N6�1CZՇ�L�m0��͕���bgl�q�VN��gFD��h�Ն>�ۧ�7@�su��I$�I$�I'F�+s�s;���e�� �	_fp-��w]����Ũj�1���W뗧*pÛ���!�<@*�"�r��1M�X����l��.���%j�rGKq�BPw1;���}��o0������$�9]I���w��]YЋ�%�wgU<�$A:����j�.�W�=]����@*�c���4U��A��`�X�3e�T*R�gZ=��N�l�V$��P
#f]]AghV����j���l,a��2�.�٤�*r$;�������KOX���4P�ׅ*+9��a�M�Į�..��$�.�dj��Z�/��j���͞�����21yyL��h���z�x��j8��`�h+!@4[��.�{ZO�w����0X���x����w�SG; X�*��ջ���.��p�J�d��c2��.�,V#&˷@a_�ܬ�IŷO\�I	�����>�$�G`�ү����e��q��+�rP�;1m3e�g�
N��E�����1�T���5&V�i\*�=C�;R��-��#�)7o5��X,��J}���g:@��\17M5$9���rDV�#Q�S�>���-|�"��'���X�j(.�V貍[S)U1E*F�C�""�Z� �Q-�VED�_#WXb�+���V1��6�+X��"
*ҕq�r���DI��j�-W���j[h�k���eį�,յ��z��J�QDUkJ�
�Y��*�[�+��iU�jm�E4��Z�Aq
�Km��:����[E�l5�i,k�b���̬�*�j,�����&�٫��B�Qun"
imb�PL&MZ��rŢ��m�v��ƣK��hA�����EX��*lM*&TFKj�*Zk[4�kKjԣ�7��2�>�©UDE�
����C�A��"��*�pZ�mˉ��r��{n*�l�UYmS(���5�+1��X���L��m�qP�E�ܦ���ݎjw���4���v�C�-�x�U���q]ѣ�������H�=�����ىƱ��jqpf�0J�So����ӟ��v�K��{kS�^%"l��'��"�t��5����H�P�;�N��ۦs�h^&��u�Tw���bCt\i�"%Ɩ"�S$i�=��X����P�z�gt�{���q֤�T��v«&eC(x���(��rT�C�}/5�Ů�Ǚ����4A�^@��FW�k�~o���ƻ����1~�,�B�,�P�-�������PS�P��Z:V�8_rv[�H���+����`B�.3���ܖZ������b�`�����:σ��H��J��P�3�p�t���UDa��Was�'X�OҔ&�����<;\)�Z�`
3�c 첎�u����&���28�/W1��MX�,q6N#��v�:^�7BѤ�DD��wejR�������5�r�+�.*��h!R� �-'���ĸc�w�.rZ��MsSYAX�����t��vO��P��B���7��U,����}M��Ǐ3��ŏv��@�R��I�9�^�╬0�A]wul�W���K�8�)W�����k�-�G4��`�(ȝqE�Mzt���i���ڶ�(�v��o%�{���n�kx��n��(�<�</6���@p����j�����uN��>�������b���-����o%���EŪ��K�y��Kkr+<�q�U���r�y1�v���H�-�xVD�C���j�*/U�dk�/�'p�}�ȱ�[�ͽ�Ք�?.�/��Y��P�H�4�2�P�Qo�t+�{��:9���qn��!گk,���(,T>��i@�����txeOR��eź����ߖ>0���h�	xW�����-
B�W*�F�X:�%���\5kZ�㲄�Ԯ�Zy7	D0D�2)J�k���Z*��*�,%�ƎP������/w�~�J9In�	�!r����(�vXU��7��Lܹ���S(-��=��4�[m�*U>�C2k�\F���k���y�0��>�Jv�e��
�@;�Urbf/7���~��B�Ձ���߄�ڃx�Ej�e!�3eѬj[|�,�����y�r�M��f��X�7B�w[(�r9t���%�{@�I�`|�~9�P-���B|��s3|w�N�q���
�fb�sx�T�A�u�Ă��/�&�ݽ�A�s�N�i6�C��ԗ~[��7mo�s����� �����+�h h�g�:J65�k�4���2�-���ŗ)�@���R�&\�@be�B/aűb�e�t41���s��Ր�����faI2��9y1a���50nLSR࿫��*�/��e�����n�>ՙw�[ A��P���)%�u�$4f��rLJ�Au�J�G���?o��B��B�0���S�u�3�UYb�I+�]EP��SR,�ۭ#X|����4�c�Q�=�fA�.������hX�?�h��}u��w��R��ǍYپ�J2{�Q�Q~C�Mc.���?��:r�ug���	5(�R�is���3w�L?��A)�Y��,�mSiVV�#�[�hڮ��o���� �Y�aI��V��xY9V<!�3���
�Q�؟LeC7;,ʛ�'���n�r�t�_)q�,�����=���!��!R]����U*���;��:�-� ���O�|��.�\S)�7�+-L"n�-K�4<i-��rAKC��6��*�f�!�@V1��ojL��Z����=�{	�������/#�;,u������z����;�c�9��ӱ�!��Qfkw/(\ă��tr�*#��9�5J<�T6�g�e��b��Q�����=�
�dt�(p2�z�T���ͧ��7�mƸ�\6�X�V��r|�R[R��j)����,�b8�Fg�sK�hi�zWY�~��]f��-�t�wu��*���.�1��N���47�.��ڞx8�_ ��[>C�
ޢ��''�@��%�x-�^�v�*ٞ�*B�lC,12�L��S�7\�Qm�q9�Og=��nu�4!�� ��GfӴYb0$��h!��p�6�~�|�[��e���=�G���qo�N<�]p��-0���%���f�ػ��o u�g
p"�e"+��T�ʲ��@yr���"��r߳}�g�Џ����e5c��J~Q(לK�AePgM�!����#2j8�<|��$�,
Y�l_��}b�Pc�A�(;ָXʷ��0�QU�Z��y��3]E��˭h��|�@׹'^W�+�Wݵ���O�^G����V� �N�kׅ�h3�/�7�[桤T��QБ���6��NM�5H�2��*�:�K8����'J�����N�����Ʈ�=�%^u&�����9��I%�Uj�,l
;����^{]i�R��h5.�� 1��~����>�]f��ǉ{�{�I��=Z|:���}��:�Ucqu=�}`�P:�3G���vU̸�\�������Q�nx�e�f�.�G��3����Gy��t��XuYq����>
]H٘NU`��l��3��6�(�۰"�Ua���=��q�	�=��wuÝ��/WJx:|��`��dƑH@Ӈ���1�41J6�:D-15;)�Dn�ݻ\�1�����2�,>t�[��	����LHd���=����m!O7�|��Y��-�NM,Ӆ�8}g��Z(��.���<3��y`���<:fT)���$L�zr��`�U5�tV�37
o�F}Ƶ��+�z"�?HU�'���QuR�"�ur�]��˶��R>|%x�K�Pa�Z=�1��ث�B�C#���!���uB-��t��|;�>�y\z�\�"σ��a"ǵ/x��,e�VXZ �G�-���������_��TޤGX���eVb�m�iC�PV��AS9�-C�ۗ}w�^�3N�}Yܶ���֞�7n�LH�E����V�#�YY�s(�����\�{o%��:��u:���#��ف��	:g�;\)�1o��%��������0���~���f�[2�,�:�����8\�5DA��>�kA
�����d�q���[�}t�_kSS�������S��C�v'��]./����T�O�x��J�S&�4s�M,��λ�{x��B��DX��	J^�6�v$��9��<6��r��0ĺ�d4�����)<zD��{��Cb�,r��-�"hr��W9�:�24C0�t����QC��G�*��U\�.�kèd<<o��K��<�g��kr+z@�M�NW+}o������:6M������Q����K{uЭ��d�p�Kր�N�]�����K���l�A�
��$cbF��@���I�h]RµI�x��h�Y�%].�,��V�9ЮƚGe�سD��<z��}�R�l�je��{�_V��R�E�õ�+�u�lS�M����,�O1�:���}��Q*���4u�o'v��E�&���t��,Zen��Q���0ej�Ѭ�I�^X$.�ĥui���sw�D�H۬�۷�\@��}�C�:�I_t�}�Aٮ'!�������uś�����tmS&�g�݌�Cp�5��p�<J�5��ҥ���8]�Y�YX�9��O����k�ꬱn,
f��Ŏ���P�~�w�A[�}�kS9O�i�)�b�"����B�m�9Q{'بE%L�B{X��K1kґ�hs�����������[�����E-�Sʸ*��X�'�X+�!z}�y�=����\�@a�w�=I֙�t�P>�p���֋e�-��N�@�C�u�z�Vb6�P؅.Y�uX�^¥>~:�%�����tW� m}Gϒ6��$�����DW#��@,.�U	��((��7&)t�� �#
'ǶƉb*v��sQ�f�"iW���f��)%�!��K$�qRc�9&^��5��ֻ3��]g�0XT��w�[����|=OP���\|0����D��H�4]h�'�^R�Ƴ���r/��2(f�p7������{"Ƿ}^������źv�0'LP�He��-�` ��h���'t�Eu��wW� ����,�}�Ғ��Kk\Y(M�������b�}m�Vj���+)"�ee3X,����(AٶPT"֪�J�ވR�?�i����@�w��|7�oBq�M�@�"�3�P��MU�dU�(��:ٺ��z:
��Ɵ%U}U���'�#@=u���l�B�"�p��Zh׭	�;8����1r��3���I��-���)�c�3�j�k�#:[��~P���|*�d���.�'��S��u%�1H���\Ed
=�(;쁱d�be<���.��!mT|�fW.j��Z�P#�nj���g�X�,ٷ�$r��.�a\�.���\_��i!aP� ��̧C�z�˭<R�q^�#6��!�(���Ix�sjR�t��20�/=�@ ۍ=B6`q�v�,:w<m��E-2���,kt��_B)M�Q�l*{��=��z��|pq��@a�鸇�	.�[�����`c��B�����)��dH�!D6!�bD˝2�:�-	n���i4�����d)8�������8b�ҴYb3�K"�R��!C�W�����2�a����ɩ���)��S/���-s��ã*>�/笊G�q�ź����7�3A5�5b2[�)6�l��nm��.p��H��#j8��i�
@9����]l��#� P���/��<�����Ԣ<Q�JΌ�jP��ў$��s�
� �d�hR���j�H��A��}[EV<Bb�&���]����}d�5��X(����ɍ�]s.!��Tkb#��j�ϒ�_���x�ĩ��ڄ'l�C�De���t�'�f�cL��n���n{aSb,m�:��q�o�y�Zrz�`�����=�8�G
�Ȳ�U���O�0�C��\�D�<xR�G�{�1�}���\��:�Q���v����\{��0d�V	fq��-��,�Q�9��:j�X4l��7��|Ƽ�st�8�|�L�T��-��j�F�Q�X�*k[��e��X���������oS:�QnfϚFl��=5ks����Y�7;_�K�ZCN�H���G'ԫx�0:����b�m�5<%�Y��ov��73l�Յ���~�<b�t\q�x�c�M{��+�
�U�N]��G�q�1��^�d��A��,��kX�d���v�^xWT��VŘ�y[���^�x���Z;��{:���[���-v�,�s2u��ժ�Z��Q�[{s?���t#l,L)a����T��B���hA�;��[�
���+��+ �V�	hz�� �^�p]��M�H�����ۋ���B�ڃ|��04�s.#�$#I�l�+yco���;�j �F�?K4/�ȡ&�ӣ�T�0�4M��\*Q����.X�yݭ��^�Lh���Y�S��1�Q�g�P�)<걿x׸�t*��k$�����̸�*��AQ�+�D��������������YgrR�+�������%MЇ��4�� �2�o��AT)�J����;:/�O�iY�����o>]5�E@~�����:��0"xx�m)
A��G��R�y��j��72z�c�ka�H�"��Dja�u�����#e���/����m���h�X���2a�4Qތl�cb�,b�߶d��/en�皘=ӳW����%�����vF���$�Csג���(�Se��wȳ�G�k�V��=[�4We5v6�V��%��\[z��ױ'/ڼ)j�uw^7پ�=ǂ|F�
̖���*�hn�pQ5�nS�f�;��uëcж�K{����>vk���O-e��]��׭mAFm����1����u�p�2��mXI]s�I�_=Ņ��>xvf�Z!�a��%���8��v�Ib�%��	���6�[�l>�u����������5��n���m��
�Xޮ���}gl��ydn�"/#�o~24*q��T�5	����o�wm ҤM�HVC�R��m�{)a�!ݴ�j����tW���LWXbm�oo7�DA[Wi����R<H���������:�<�I֛2�W5WP�9�TH.���ʴhrîP2��7��%c�5�NZ�{; ��y.ҝi���&%�;)opS��#��ej���0$��� �ô�6aKv��S/%mF�<1���W �@�(QR��{pQ�d��1��y���՟@�i�݌��_�0m�L�vI|[3me�Q�Vz�ۼ�
ې���C����4-W���<K��#XN�4#��{�+��`j�"�U�f�Qݛ�%��by�q:F�53s,�(�2�C4hS����z�� gl[V`���݄K�h���3#ȩ��Fr�3�]"�lB;t(P����O�iqRI$�I$�I$�dc�.�
��a�����O�\/.�Vfԗ�n�2�������8�0n��8�Dҍj�i�_O]M�7������~&<�&H���%�%m3!�F��^̸Qʆ����$�!�̫Zʵeu�҄B���]&�WF�I
AVo�_��;CN�S
��{R�,76�h�/j����3u�GP��V.��3���2�4Hs<NeX&�vm�z^�me#��X#2.��-��l�ײ�If�Ʉ��GMT�8�M��+�1�5�k+Pzb�[Ä+atBr����n	Cq��(�wn�e�5#�C�5X*�Z���?[P�v��<.�]̛�Y�4��XubW�ɲhY���8z���Y��Y9���2J <\���M�V�`�$���qӮf�ǲ]�F1R�K,�iΫ���S����yT5��AY*�����vjjͣu/O<*�+u����b{H�lC	�w �La\Qo%���8���.]�k�]>
�݁�#��c`ՐR�كt�}% eweŢ>� ��d\��ٮ�bX�o���o`�lH��'!M��mH�E$�܎C
�Q�������}����U����5K�|��g�C���g�GN�Mt�f1�V��T����f�ffM`�-�Ta����m�����7��5��I�3Ibi���%��kV`�"�̳7�7��E͔ޔ1���T�K�r���L�Y��Z�(�4:�t�f��kx�Y�L�e-ˆ4�*��k2�i�%�b�-Ƣº�WT�:�(,����*���Or��j�TW,�hm�M�z̗z«��aAE�*�K�7Flq�Q.�Q��ƥf~���bk������I��9m�eDj�-
&_tSH��Skl�,U�U42��5K�U��T�V*�4�ʃ��D�E���2i�UYQ|@��Yʌ�n҈��J
����01j�U]� �H__�>�3&���EU���qd��;�xL�2��
T�*&p�B	��C��u54�]͊��s�( �#wR]�e�>i��޸K"���� 8*����m�<+3������.T�vm�Q��;g�m${U�ۋ,Sd>��Po���������P�
�G���۞>�7�0�\\�v�9�F�?,Tۻh!�Bvh�~<Y�lH�
��fTީ�{�Y"Pʮ�N}�����[��8*C/�%�(J��5�{^���b�#��X��	vi�����]��C����X:eV%��q���&mݶ\���p����r\���kDꍦ.b ���a��n��<N?h��Ͻݯ;�E���MT=�*��P�qf�>'x����x�[3b��{iX޻S���Tc���˳��ոl�7�b'�S��w�W��y-揝�x(z�Iy�Tɴɛ��}n��]�8���ވ�����#���,�F��F�[,�h���s#����+����j��U���D0�lj^�إL���f���>'A�Gӯ8=\2a���"{{v-��9�v��ׄ�#1��ӽcHm��N��� �u��[Z����h���f�a�����{������iT�3~�e�GC*��6�fC7%t�-�I�A����b��yF�vGV�����H���<��ܤ��<Q�����	�3�LXw�S��ߔA/ܼK�>�Lt��:�U��f &E��r"�E�%����$�JI}��g���3�]�e����"��Ù����,"�u�*b��c�W_5�<'����Y6�&�;>��u`��[�+K�_�d�t2eW�am��SmڋW�-2� }���X��z',A�$1�G���ۋ����8w�LW��!<��I�S�S��j�"�%3g��[сwP�r,����9bn���Eg��}����TQ@�y<I�ds�`(G=x4�&�^�sW>b�"��rǺ�C�����穇=KC��:b��9���壟֯q�8ᢺ�h�����ٻ�����Uw�R�
#�7��R�����p͸f�P�S��35����3�Vo*;�����!�W�N���#~��dZ�<��g�j<s���}N��V��=�4�:����b�t4�7��I�V�̒��Ф��<��^��ջ4��
�VSskd�Gdټ���v�k�]���NULf� P����6ܭEd��c����{��jr�'����V�H�y��k,T)�ri?U`�����Pp	�Ψ�?/���Thn5�86�����|���P������Q��'�8�`ֿK4�q.4��0V��!*�ܐ����ן�X�o���%�x�9U�7He>Lw�+ĿX9�����'F�W1<e��
�h܈��\<<�ϗ�F�┖�:�GX���9ƩL8�;\qx?���t|,K�W	C�hs�ʇ�sШ�" Տ����a�i#�񣾙<*P��S!>�A���;Pi�*{���ΊNtX�}μ)u�<�M`d�-S�s!������)�]Y�HVU^r7^�ʆ�Y�SA��_��'�d��u��fp>9\.V�q��/z�c)y��5�C��m�
�9�
�T[�"tB2E� �t-܃v�(��:u6�F�`���<w*��:XG�h��t���{�DF�s�.��Ř��4�鹤�:��uӭ�9��˚�K�|����kc�Mm��WNW���������yuw9ޕ������.[�m���&e�&w�ʃ��Eή����Ϭ�ԃ�V�XiT@�qѬ�J��z�r.���7��P��=*(sX�M�K6g�oS.0M������G��z�9�m赨,��H���]6d3�d�FO��M�K���e�E�4�qF���\)�n�������*�����4U�}G��5�5�4Cgx�^��:�;����h� �͂��ܸo�#.����Dq.4��<]�#�P�Ņ�C���k"d���p�8�v�=��r_ueՒ�k_�����tK����o����[�'���~��4zg���U��R�z�\�px�ֽ#U�q=S��K�*!GJ6���
�P�k���
U7z`w9���ǻb���q�o;��HI=�9��w+`�>^P��u�؎��'�g����7m��7lQ��[ƴ��f7��Z��Dx�CB�������2�����V��3�=8�u���rR�|;��o��|�<
b���ڠ(�%��ȱ+|���Me���N�'��w����l�UeD���WB@k���ic�V�Y!�r�N�.����ם8F�{X8�{|�ڛʮ.hpݾ�9ծ�=��!KҶ�\J[R�93o�I!֖�v��>2�^���}:�T��[�A9�HTS��f6Yf
��G?��ǣ��FH}s��zž{�U��`�0x�3��җ�����l�X��?z�>*۞�w�w���Z��mŎɢ�l�e�RK��슿'Y)�'3�����'�?4�2fX�<J��~��Rϼp�2�x{����\�aO^v"�/�;P@��׭�q� |q�B��>���)О=A����}௖rXb>S�qݱ��m����p���U���v5��S��[8и@��'��rv�a<Pw~��׬xm=^�<*����t�0m��ǥRZ<16�����ˋ�x�O�?�^���r�V��h��K���©ѭUn�)f�к��<�{1�u�}f���(�p�ӕ��"���Cp8���tKؗ9-&üx�,w�?v�t�U{�4] \�k1�7`�\t��g�X\�t��N�e����2��t+��d���쫼ߥh�C���� ��d��}��h��/�ʒể���"������3-so*o]�N���Mp�OFv�l�b���[�:�a�޾�s8��]^��j<�,�	�\����?�Z�=X����:ct��{���	�b�7��^�q�ᛨ�#����Q��9�|�j��/�Q���4gc�1�H(纈p�^n�:��?>��k�t�sY�:U��.owyDly��P,4�����8g3���p��ۓ>¿���T�9��Q�c�x����h's׻[�w�� ����B��ʥ������?Q��H�����}��2аEyZ!�m�P��)��%1a�r,jE����U�Fe��[*��x����(8w�U��>v�R��RcҨ��Z��9�^ V8Gۚz�gٮ1[�.��;�.S~�OO�FYu�*L�������u:���wPQ9�z��ua�]n�P'Y�[���Jq�:�k¶%��^�%�{�����#P�Uq���0X�W��<��b6<矆��}l8W3\�;���5H�hd�xup���]oB��Y3��t�kҶ��.�^�Ræc��ڣ�j��=�km�i��'+4*=C=�zv���u�����Y<���7�U�y��n����U�S�/����Qn(�;�i�r-������*Er]�=�Svc��BI)PW�ĵ%�x �G�(�N��ŗ�v���C�+�>�"CC�x�csY:C��yB"F�w�ߊm�#f.��`�4j�O啰ˈ�oH��OAV[<�=N�5s]�}�l�d<��U�ةT�#|gQ��_K�F�ӦYfN�(СGKQp��bcqUe�/����(�AB�|�\���؎=�qû��ibt�,��NJ��j�}H�Ze��1CU�z��G� :9�G���C��˿o�$/.��=6�W�y�F�*d�ev�)�M���#L����2�=��e��w;��v`�8h��:"�h���ʧsbJ�)����)�K$�7<^Qo[=�=$O��Ph����x*t`�Z-Z6��p1�ʆD�R��l;US{���U;�D1�$u`���.!FS�={H��poƯ�v����F���w7��L���F6�����j�]u%X�ZH���E;|)������ѯ�y?���e�n��y���8a�����vw�7���䘅�	�Rv����d������koд�� %G��u)���NI�y����^iْ����wɗ��U+Q��s(fUx+�.֋꺰�kn�H����N�>:����0D�QI����G���w{bƎ��X��Y��:�ֈ�u��K��/fl����'�96܋�۝��z��*���c�6K�a{Q]*]�>�����A��/:�������su��ܚb,laWO��:�V9;�-��ڌ�'D"�&FK}��=q	�SG����+��^T�c�
C��N�c�����]�J&Vv�qiD@�,J3g���DU>��*���xxJ�^3��O=�v�SVP��=O��J���G�Y��)���2�1$��P:k;=w�g��4��l��ԺO4��
#�IxT�q������X��i�p��G������=Sy�8������]��wqZ:��YO�l�����%��GB�lu:KjV��؃-D�w���G�>������
�����l.�����k�B��)V�6���lәGC�o�"ƎGY����[!}3z[7ƹ�ᤁ����b��86�yxeJRH��;�32������9��t�����MP��a<�r��[��B5�G:�6��PStg%Ȧ�mwU�7�g���[�n֐������ܓ��T����9O�o�'*4���,چt_M��d ���+9�����+�q�Y��+�Wt�!9pj��W
3~_n�R���e^P��p��ug��\�z>�y�]�ݾ���n�0J{�T|�F��Z��K�|q"t�º��᪽ �kǝ��}9���툊�J.f�a�r��AS8�'����s��Q�yv��6dܖ49��& `jA;�HZS��=�"xx}G�m+�t���5��F�)�l���N�2��-C�e�i�ٝ�*���&M��u�����9��؂&�<4@�)�aC�6p�^��DM �=0"-�W����`��6%��D*������O�q��G�܆])E���:���;���S��<qd��[T2��,Ϟm[�QB�"�P"�m���:r�o/q�]S�h�l����A�!nM���J�D�p��MP�(qNN����of�����������с4�ȁ��+���PY�.�fȱb7oƨ��ٵ�g5���Wu$ѤT��D���9�p
��9Aӛ��;��a�:=���&l�q.Q%�����'��<�� Ƀo+��Y���qvSI<�������3����������}^��:�����z��D��~�~]����Ը:�@SӒ�7^�)Y��
̊���],���o&�1?^�.j�G�,LuD�xZ�w��D+"�8�T7Bz�FD�=��O���ם��w��!��a0D�;B,Z�x�Ǉ�b�;�v(5�P{"��r���j�o�?Q�
��%�|����&x3M���O����;hM���|b>���}����WX϶��g�PZxx~b��P��8^��� �/&�pa2+�7o��s�{��R����ԯ{��nw�
���.��,�v"�H�ض�e�bhoi�s�_9̺ ��<�S����2?:�_��
����n�bB�`�Ύ̥�����Kg�EZ�%�(�#��m�ր���.�J��P�d����fwpyݜNQ6=�Q�x��{ʊ�o��ǃ�cIj	y�)�c��[��E���:���a�Ң�t�`pߚ�k>�FMC��"�j}C�st�v�Mu�;m�٩+~t:�wz͗��]kٰ�g��!5}ܬ�/��f�uZ�!:�<�A_i$��-��%�h�]�ۦ��;,�}����w����b��@��h��*���Ș�5Z�>/������Q])njZ�RK����+z|��N���դ7�`W�j�5�k^�N��y$�"���a�u�k��Z�p�Χ5˸f�	ր��j��"���Ho��=P޶+�C�I:�2��f$ot,f��t����=�j]�0�1쎶�i.f��ģ�h��:�v�ك+n���[G/�n�K����ۮ"'�*iR�� x��V�oX���N���RR�.V@�-��dK{��t]�޳���mr������X�6BSnJT�N�5S�H���s���9$��ܺ�1Yz�J�x�UV��rc8�fp���(7�M�id7J�Kś��PY�<2���`��|�֙�@��S�.v���4�`�͙q�6-t&��{�-;t�`�ǀ�Wq�x-3��v|��:,�b�1�u\�;�*+�x�s�F��p��fH�r�bI`�y�Nm��}Xrٛ� ͼ۬ɛ��d�u�7N�R\�V&�/A�Б$;8r��������5�-�+fjrI$�I$�I$�t��T{��|"��qH�k�2���{��}xu$���n�M�,U�H�s�	�'|��R�������=+"�W:6� ���J2�0�szt�j������Q�i�^�n��s4*;��^&#a$��'v�X��[{S/���"�>Xe
�)�B��`�	8����e+�5��uʔ��	�n�qP�[SuF�+��+E�p�W
�Җ,e�֍��	R�4�	��I3q�NDو�]�H�%c���1V9\��[Y6Ύxt'Bp��k˶R��U"��'�g2*Wp�DAP�C nR�,�U���0��WݒwS�+��y���qX�ړ�4;S���u�^�J����ap�[˭�!,M�3�������ʕ�v��"�n��u�ݯ�^}I1nԩW�V뇋ˊ�s�09ӵ�V��
;��ڹR���wTټ�\7L�����e\�Q��['^����5�jV���ۑ�`Y�������$�G�6�o}YnH���u�.`1o-�*Z�.9��^Z�1Ȍ�2�R'�9�'#��[$�7mH��[���eeWt.�.�kEc��r�e���iM���Sn���IZ�`��S32fR���a��;��Leb��T�P�L���2��2���r��4:\LV��V�Wz�Z\��J�MsVU�Q��[ur��4��U��e34�t�i�C��*-��2b.�WH\h�-¸혋���i.��ϵ�O���`�c��1��ZbUF�[U�]3l�Z��]�f� ����W5��eMm�kI��5ui������3YL��k[�ė.1���s�k��!�M�Y�f�D���ģ�]�c��Sl,��c������K��m�޵�n��Dѳ�W`�mj�&~�4�P�+�QQ\--��(*ʆ8��Vi�n9�5�E�Y\�0�h��:ʊ[bԢf��*Bڪ(��h��j���ՑTE���liQTщ�(�cF�ն�ailZ�D6���O5Lݡk(��k0AՃjʕK�ȹh�Į� ��E�MZ��4�R���Q��L�ʁZ����e���y����*�30��s5���J�kQSw����&��./5v�[��5Š`��^�f�0y�㴴w8JsG$�����+O���$���nLPޘ3�d>��GD��Pr�Q�@躆�(wB������ޞ����!��g���n�c"�dV6%8����J��e�J�m/�G1���\�ܡ�������X��z<���j"Utx!�;q~\�|7ml�j0�+�����\VзZ�ú�6-j��e/J	.o��c�������7���"�f�$�ґ�P=v3@�k"�Π����'�znf��������G�+
:�<h[�U��e�X�R�+}Ֆ���s=Py���zv=Jjn�{�=Qd�ιVb�P!Dm�7��R�4��Y���Y��!�t���u�Wf�T�r�#�t=C���Q����W/Xua�$V)��w�*�w��Y}ҡ��ܒ#ܞ�r�L������d#A�
Q$�+�0��`;��qKjǊ�C_�k��H]k��b,%=q=��3��Y�Vÿ|���7lhY�4�P$1�5������t��s�뤓p���^ �-���^^��Ll�h"/�����K>n�������a3r>��u�.�	4�?����^nD)#^����Z���֘ܝ�N��0� ���I�n��Q�v��9سJ���y��F峱Jtd�R�ѕ��RY��{7�Z	�w�1�j?:)�:/ﱮ�E�N��5�u>�n�߶f���M�v�����K�澚%ѲURՃ���D�pN��֋e��j��xxa���(Ȗm���!"ȫ��֨�^�0��Oʕ;\4l��u�n߁�L
�k�ߨ�/� ���?>\���q�lHx�1��OƗVV�pe��������/m}GGP����
�H�ﶚ��0�%xn��];����Lj���T͉(tQ:��!8���N^��Q'��#6B����۞�?M���Ua��R7�4�_�0�+��Gc����w��bٞоq�:Uؽ���~�4pxR�;Y�@��;/��Y���XG�E���Ӯ���m4Vy{�wvw���LB#�f�(迡�q����v�����Rˋu����͔����;��z���~���ڬ�]�c�ECV����r�ӝ \"�E�:R�C�W�v�63�k;���e��Zg��}x+p���1z��N�W�x{�L���\�sw�Ո��L��qfݮF7�B���BP��Ky.�< 9ܵ-t��r7�R����8�pז*fU	�O4'f����&��>jDs��k+rș��"����R�5,�
z��q��H���nDq�9�õ��k����/]+�:���������z�C�����V�ۃ�n��w�����MTE�<�5�<�����Ɠ���s|",h�X�}=�nL��*1@U����9��%��K]��N�1ӥD�K7�D-��4%J;c�Ȣ;���U�%�5o�'<OK�\Q\k½��Z�(�~
yxAc���a`��o�_q�ߋ��~��""z��]�yXU���F���6MO��Ć�>\)������w+/l��9����W_�k��oۦ��a7���AS9���/|��ߔ����k��O] J�md��y�8f*Qf��Ym%��W�����b��1ʭh!�U+�{�ר�.��#Ssq�Ș�g���M݅���b��ҭx�|6~��o�D�����ǘ�:���u���k�u�<������V���3FD�H��Cf�{�\��r�3@�Q��ŻΆ�.R�1��7���YX}DJң�i#ŵm������|���VTF0��*"�2���{-����y�ą(I͌z6��F	k��b��`�cw3�"6�u�|%#��T��x���Йk��赓6��B�^e�qՌ�W�s���KO�Y�_��S'�Vo.>/��ĻR�����Ү*2l�
C(��Xk���.67���mo����Ҏ���5o��J�G	,(`����::x������V�5ה���	�]��hCW��xz�T��,�- �g���zj�X3��蘗a�ǅPc=zm�����$NdP��(X��zܣV�D.Y\ 2�ߟ�������$��n�gw��g��:O��\)Q�t9P����|%'��Â�S���<}ks���^ws�jQ� `�;0��ѫ�9�~�~&xNiu1����𡗿/:މ��7�9���7m\��L�E54���U_����(���^Or/Y��ml)��n�8v��<�^�QV�V�N���F�?^_�k,l�=D�m` z_z��a�c�J���]�������>��+w��5��`��p����u�ZQ2N��W�7$ye쥜�� ��ys��V����������G�H�9;��=�4�5�[Q��5fE��1"%�
��>Z3MF�yټ�K(��X�]Q�N��k�Y8�
�y���>��r�"�לA�1K���٢�ʝ���cI�EO�"4-�L8@�.��d]�u���CsV+f3��^'�
���tlC�2�"��*���Γ�\���Ϯ����.�x-ԋ+���n���Y �M���eZ��J���_��U3K����i�g7[v^\��>Jk,�a�'�_[4l�pUW�*�{��ȥ�X�_�_�a�U��,�yӍ��f�4"F�G!��U[�б>�����]{Q][�!��e��K]�ة�|�62�P��!�&zE8E*�7�\�h��B��/���ˆfsKD�P/K�6�t��}<hZ�em2Hґ�P�V3D3YRn�y��{ǭC�S/ӎ�C.�e�i�aͥ������^'4���p�n�[�T�M{l_L46�I9�;��+����}�ʠ˰�:�3�Z�s�}�n{�Z������W8Ls��cR\�X���X5 ��P�0��xAZ�7a��c���q���S2^�����ټ;"�ͫZ$0�Ě�΢��=4A��"UY[��� W{o�6;Ue��wK:F�.bG@�$H��xcZ�o��#z喛��9emS�O�V�A��K8���./c%ՐA�|�\�ё�4�gK���X�Ǩ�Ɋ���/a�r:�ڂ9>�y˭2�;�/T�<=A�5s�2A�c<�L�<�m~���B�
z�DDXJz�w<S0k_��'��G�{�N�ԩR�@Bƚ8)�EZ<A��oCg*���|�5�B�	�s$�O{}泺�����=���88Z�� 5�24^^��6O �KV� o��MM^B��i�F��C�J�h�:2��>.��;</����t|�C��&6[s��t�	k�p��xx@.^�QT��Mӻ�Ne^}�`�]��Q�����v�{��GGP��yؕ�x��U�P���<j"�� �s�^��\<6�>u{nd3�:Aq����8Ȇ��_��E1\�5F�n]?xu��X�'yCRhh�/Qø�we&y��<�)v��KL��y��N������/�����'���s/��rd�b��}Wn�9p+Hv-�I������J۵�&����6^��g�sbX�6C��l����M&�ų��R�1AO=�.f]A	T+����B��\���԰�I��.�j��-�W݉Q�ɤ���#(u��YK���+�V2�Ǵ0xxq�^�=b58�����v�W��75z���ޢ���W���B�i�O]b&�s���wk\�2��!����(�UXFo�J�,�v(m9=jvi�	�>�%f�8�{�jU�7��B�Z���m�Dtl��ʩ�%��zкg��B�K�y35oN^�A���v�U����gہV���9/����b�*ct;���ԐW�E��lw�/S��B;�}
ź������� o�E�s��M�{��t��U=l�ݣt%Z<L+���>N����\�5n����?V����ilUC2�2c���8`L�V�J:�$^���[��4TT���t�T+����Ê����R�˿��w��*��nQ	7"ʽQL��FK����H�&^�w����gS���,����3�a�s5v�Gg%�'4���Jά��3%-=#r?��=�)˹|$�/�����2�d.�W/�P�i|��&Ά�M/{=�m!kv_i�V�b�|}�ue�����a.^�x:Ŏ'&��̸������*o"&`�K,8��f���15�Z{�(_�XE���E�o�j��=�~ܭ}�E��F���^'q���͘b9A"=����y����{R���e��GJ'�n�B��ӃΒ� T��[i�a������z'M^�ܐ$�AY���]t��,�R�ʜ3����)����^&6�K!�Y���R?M�g`>���ɷ�9\S�Q�jE��!�6��
���pȗY�+3	��T7U'u�j�`!�ち�,�Se���F�{H��p��N��۬����W �*$�uD��f�xPdp"Kf=�6'���ڇ�p3�ײn�A
3uhu���
]HS0�94U��,��m�#�J��)Di��N��elO��l�V2Y����I�<iyM�6��CC�U�].Խ��s5�X�Hm�ُ��"cJ�HU�JMė�4f�&���e��Es뚰�;*%�s�U���/:We�l�ra���YX�Zg׳�T�a�EƮwu%�x{�)�M�F��ܪ:�J��<P�'G㣣��xR3�*���į��m�w}8����Z23�.�B��6O��p�h�NC�"š��|"��鋄�b�5���٨Ih�����v�Gt3��3�P�L�,�w�1���)~\z)�sl{{b��̇��#,v����(p}D
48/V�,������?{=`�{*�U���	S�� i]�FN�ȿS�K> x{���f����z7:�&pz�O�QQ�<��F�6�yW:R%�Јnf����HA�3n�Lgc{Z`���<���%��>$:h������b��1ҳ;:Iq���cw�G֪����u%��PeV򢋳��3��ˢ������w(��y��� ƪP8j�HVr��m���D�ZR$T	�Ǘ�V��A�^�}8���.�0��ui�k���d�pU~�A_ldR��ƒ��K_���@|ǭՌ��*]}.�Ϩ1�!�WY63X���*�5��{��:���-�j��S��b�������و��/�rs�o飱M��P�Ӹ�IZ�P3)�t!�6�길��G۽��G�J�Ae_��[�g� [w��8���|P�N�}B	��f�r�q�%nw��1ڈ����P��I�{��z��#�P�7����	�B�P*�6�ތ��u�g��\x�,��X�8�"���\�V	�`C*r�<}C>�^ ���H�sǁ�m�[�&2�u.���f��}��+��j����g�n�&&��Բ�e����w.��ڄ�j��n]٦��)G<
P�)�T6
>'�]#~3��ʚ�O��#�h8��n_"����l��b��Y|�1z�N�!�J�N���&����+Ȉ��K�f����sɂ7����/:+�P�D���M����I��[[WIq��<zv�p���B��]�Sy�&}�Y[>�~a��Y�2�zz�=|��S�Ӏ�b�p!�'=(׆!~4u�Y�.�[񓺰m[*O��9�;�\`f���B(�~�J7-h�+���e�,:f���EL?��Y�ܗe�L�A��9�NN�$�0
��N�q<O�U�b�tC� ��ie�a���B�W�yw�(V��W*��e-�hN��̲+Vv,:������m��Y��nt)��2��jt̛u�p���:�v���[Ij��F�����QU�lU�&�r^=0V����iT�[}�����*�+���jJ�Bdu�����wGiǷ���mc�fł�U�Gt�2�+E�+���ݩ����LY�j�v�֫��8�iD��F;1^�����z���9��G�˭�ь�4iM0p��u���jX�y���e����eKHU�O"]W Ń8J�w�e�b��D.St����d�I=��(�m�o@ycK�im�Ǉ�Sb�uh)]��<��WF]|����9K�ӮP�&Ju˘�H˱P��P:>W}-SYb�U�T ��vis�dXSJ�wPb�5�C*&R�]0���.NI,��w]�-��\����oj�].�`��9��Ol�2u�n���ţ��u�⤭��b}���z�V�r����=3�nV�7O#�R�%�cj���=u|h�X�ХϮ��
-��3�]�(U���9�y�&��L������$i�mG����oCx%5��欹RB뮸a�Z�Y��a����+�;l)㘬�[�S����ά�&��s�k�MےI$�I$�I$�#�͠�WU�l,Q@�ʺQl��C7�ާ�VҾc2���>.Y�קgj��Y�Y��b���/��'-�x��gZ�\_ 6�"�dUu�P��Wp���:*�gdY���]늀�5k�������)��N���*���qL7Ζ��:��o�^��\�c곴��"��^�*�A��!�xn�����ڒK�v�ʘ��ge����\0PV��q3C��S��`���;�q4:Y�7[\���s38���X�ҋ|��j
"Ù�F��E�U$=]�mk��غK�X��S=�,�8�'��=�Am�أ]��+-8^E����F[VA7��\Ê�,�v���7�,g5΍C��ں/�C#��(���3&P�ٸ�P�&iN�I�Q�ܦ��t�̀��J5E�V{4n�����̡fCa݌Y��9٠U�o�Q:~�&�`�J5}��f�޵�m�y7v�*8�Yhd�6���)F���QP�����N���s'�|�C�~�}�j�2%1�l�7��wj3��+�,��{���[Qɇ;\�m�[rp��ӑi�48w#�2�f�Gq�ڑ<�͉9���$�țnG$���Vz��aZ��ʿ:b��EY�n&9[�D�V��qX��w���1�3UF�,FE��La�WYr٦.�Z�Aq���,�Tr�WwF����ZcK��څ��b��aq2���ˉ�L�*��k*[i�a\ݘ:�ʹ�2��f����"[�e2��U��X��2f\eAW-�]�ۆ	�T�oVf��k�1Ff\*
T��X�%dJ�R?h2X�h�1",M.�����f&,��-�IJ�v�i7�7Ywjk�..����|3�1���0M���E�6�������eP��ڻCHi�貺B�����a�*冽�iPq�J��1�9��Gm�]	m-̒���u����B�uw�[��m�1E\�T4�)r�2�TZ!�8�L@�jc�M}���6���-Z?�̾�v�,�-����)�dm*i0˦Or�L�,�̦c(�
"֠>�b�]�Y�,�塲z��BYӷƚWC��v�f�"(�j�{mF�dtp�v�n6�X+%JOD)H��z�Zz���?�q�~���i@�]e,'C~Gſ*vx_�E���Q}�iw.��ȳz�vT��ߜxX���_�EV �V�<syQ�#��ƋQ��4���^��_v���P��=�c��xR�Dxm#����%c�i�V[���m<�u�ynׇR����=�0_ül�p0+�k �hy�}L����^�V�ULV2%��ua��gne���c�|�v:�V9;�l�w�Ԫ��|���8�C�D�2��Y�xm#5=������C�4z�q�M�X/�:jb���K�W,7(�ŗf��/><e
��~��h��^��u�s�[��w��:�p��(�~�ב����aLD�ِ�	�2
e30dWZ��kRə9��{n�"�nz:�é�҆�f]	�R\a�٤!ڦ)s�q}��jVɲ�'�Z06�}]YҎ<t����闑`4����E�(�ؗ^'�ǹJ6�L^y�#"������"�	M�z�O-t�j�C�Pհ1�X�c�V�M]ܘwe�7�����{D4��Dr�/Z������k"�F���6�nU�fm�NA���u�w�+ZsjH�|�O_� �~���TR�\=>$V������}q��[�|&�fvZj�J�W��}n�O��p42�>\<O�p!�l>��-e�&2Wm��+��iOo�wVNm�gEj5�	�Ƴմ��:�x�G��3����s�& .�f�y�<�����m�U��"�J5"C��D��V�X��l8f�T��H���Ǽ��R8]q�-j��I���������"���YY~���h��/���0��/�S�-�����B������殇x��/܂<5�y�j�e��=�Ǣ�?RP�F�t����\s�!U�*7ԫ�Oi����2��crɋ3O�rxk�@EЃ�E��HIX���\ϼ}�f���p�=YH@;��~�QL�b���h����89�N8@�_��˱���;��,�)��%<�m�ɰ�����S��v��"tÆa��G���u��^;vr~w�VO_�wa+N:5�Ka<�Gh����>�Go�����ЋM���sn�]*��&l���w�䙊�6�Y�6�XzlW��nģs-��Z:��ݘ�sEZ����m␂H�D�S:\nE��%MOa��A�}h?�)�{�{mw�[D!މ�u�uo
�����dw|g��/[�XvD0D�{�eE���Hg�6B̛3�V�c��2�-a���#���m��\��u�P�;��:6Wkܯ�q�
���ggL[���s�z��C��P�(w�KGSԴ8�����Pק)B���43��l�Y�w24��VoG 1�:�\�̊�G��L��u<�9����Ppu|�yz����Re_4�����#�JilOF�����q�h�NC�%,Z�|%/.����̩=R��P����Q�Ҵ�wι���&xD�5���G��o�:f�FflD\��|t!c�_�{%wBT�~���8k��y
Q��~wc{��C@�����u��c}8��a@�W{Q�ӫ2,S�`f�{	v0�g�v��l ��Q��ʈ���L���o:�uu�7t TG�y�(m�3����W��,%#/
 ������˲%�Ud�s�y5��w^b%��3�[�����6��,��o��81���.�ml�*ܰ{7j�7V��CEwB�d$� �ۋ/��5gv��sybRG��>���?�Iگ��A����<N�(�#��cC��w�]b\�c�\O\;��;���:P���)�H�d�+�K����4+��>��X�4c���<�z�Km�$7M��%N�@��R�!�&3���v���#,�yV!�m�ފ{V{;z$�gV����C������0Ŭ�f_L��PF�a����a��YοF}[1���m�PdPɟ��qn�T���%��� b���:ɼ�V��6��K�y�p;1�#c�M|0K~�N�d j�BfĊp���l��^�n�����'0 Y}btϯ'M���F���V�^͖I���E���.�6ޞ%H�r���Wz��6�ʙnq���������L:3i����k��؆z���X�ާ�旷��c��,�~�}��_ӛ>��)�bW����.��3Ԧ�v�u�ș;�X�<hc�l�nQQ��g�e�lX�R�����T��e䛾�qӮʗW/I�j�8BY2'�cV��l�o�Lנ�[NX3cP�;	���.��Al�g��y힇�i۝�1퐸��#�v�%#r�㌷��uu�;wdf�ɷ+V�.,e�&�+��H�rjJ�[@~��ѱ.�!Qn(c���=ɬga�w�B�M§wU���z%�r�͛��( uD�����<��M?|��T}b��V�����	B��gW���3��Wo������|
a�\�|�p9k��elZj�^LW����Fj�$�lр��"[���q�
<%��*v�l��Ař��K{�]8�����F��F�E�RȀh*���l���S�k�i�Ȓ�@�~���;�0e�3�b��9x]	^> //먪����!��k4�M�~��^i�پt��°Q�y���Q��8���XE�ׅ.�G��T�shZ[��;��� C}��=s�O[u�0���P�X{�P}�d���XU�T}���y�׼�z�
��+)(/֪����C,E�!��,�ub���Vh��9���}�'���>��b�*�0Wu��#��#�����a H���������BB��l}����o);m�fv�?!�e��
ܵ����2)3���w���M��crv[��3,�⍥�E���&+l�F�U���n�Z*Te�w���f���k:��ˮ)bR{;R]����i�7��g媬Z]Ozt8��c�k����?./�Q��[[B�_][�{����R�p��t��{L���pw�X/��t�Rvi����R(]�s�ڽ���]Nw�}��}��#�P(��\EoK-�/�V���һ�9�b����D�X&|nBzn��-
�u�N�y눯n�3��k��;�	�Fs��[�/���L@�ʲ�=G��&�`�+ҸТt��.7�������y��m�sTyV��蠢(w�o�#��
tx�g�4r:χ�J�
�Tg�Ys[�isn�E��[��b�]!�Z��GN�T3�Z�h_M��a� �ph��xAc�b��)���}S�7",8��#����V�X���ĺ�欼�D����l���8Z���ı�Wy`T�>P���~^�`A��ve�y���͆�r������7C"�M�%��!8�(R�aL�N_V���j�$u��W$��R;Ǖ,�D���v�Uͳ*�櫅�ӫGRmVc�XXV�T|V'����ȩ���[�R|�)ǲ��os�l孭w���׮;w�{��Y����U�ouw$��Q��71��8�7~"���3���@�[\�^��
f��uo����,]������d�G�;(�/����LE�A
��O�E�]j��$�oC�"2�j�i��7{�!�
�>�l�]w����zpsJ�.�0?-���S�.��}ǒi�L�H�׏09�B��w�SܮҞ�B��xp�>H�m�"KM/XUy싽�މ 3��T��lnK-E��]E/=��M����V�e{d�d,ڷMT����F���TF�/֥^͞.-V��p�#�Y��m�Ҷ2;�'�^��S�`8ɾ��:j��6X#<-K��(���ŚZ�N8yMUZ��D�Ze�޵���V_^��8J�.�X�薏	�:2y[ir0����U�m�Hv�ʬ/y�i�¨�r�u%*[d�Ch�6ypu<����	�a���/W~οy���n�}�pn��V'	��p�h�NC�:�c�݁)�1��ϯ��/[gT�n�G<O�;���ۊ�I)Y��>J����}  k��;����e]�opNz��u��xߓ�@t�f/�� ����ݥ����.�<�w�m��������.:�r��}�<o0b�L��@�4'`b�����I��3�U��t(�9�vM��[u�����L��U�tGQ\���e.5��r�TW�fq��Cr��p��.�Ab.��.d�k�O���j݄�f�:��lTuHҳB�;mr�Ԩ��Ѧ=�_���>I�{ͮ��wN ��򽽓�ZcqT��ہš
xb�#K�Fo��V�w�]�y\
;�q�%��O|3�
����!�b�T^񩾁�\���wG>�[���Տ�
x8� S�A��1�[�1ac8��0M�R[mD�t$������c�����ۋ��<:�loD���ǵ8e�e�\%�O��+�������εb	��o��Ĕc�ɸ��M��&�X����ڕemuM��a�B{V�ÛE���@f�$@cU7:J;Qm%�^��t�3�{�2�^]���x���֫t���Sw�r�ԥ�TCqK<�e��0Թ��J������P�,����&�ӻtn�J��=�0u#8JSM����羏��Й�?|����v��L�i��U�k9#�V���^�-g��T�7��k��V,N8W!U���8�]#����j $���{���)�Z�N;΂�6�Dp��/�z*���<q�շY#v)�����FoP���v��^�����E]���:ʺ��c�����v���7��*�G���ץ3u�k�%8C�^�]�_���T<�co�ٕ��e3ˍ�F,�xҫ��,�yXA@+8�s��[N�����M��6WO[]�^��k��g���H��i+:��R)��"3M��˹�[ړ]9����rR۬)�^`�YPj�xy.D4"����V��s��0Ɔ�X�kz5��<�R��#D_0&�%�.���
�{m#�ׂ���Պ%�XW@��w��n�A[��N�.�h�������.���}Mh0gm]��A*o��Xnv=ڝ.�CNћ[����<[*h앻WR���ekZq\�:ڒԔ|��z��m���\(C���LF ���-2*�.V>�:��~&��H�`K���[�l!#��LD��yԫ�;�k^���n���X�*v�wt۹�C��>�IE���v�gw�T��ύ�WsO�	]��s���մ+-yκ�p9]�*x��j��Yc��T�u}䶢��*��!EE�M솫^Jǋ�g'e�M�̞9��U8v���{`.�4��:r�����X�s^��6�6J[�W�.]�}�'F2�sƑ��6"^�h9u"!���Q�@��ܾ�>�v�ظoiTE4sm�/_6��om�1�3�@�b#T�q�믡�� U"M� ߩ�+�(���#A���T�U]\�0ʆ�L)�g*��L��Q����"�LLDDDDG�L�"4�9|�/�%GKY= ���L��Ig	Չ%o5��R�+�B�	$  
�����J�Q�Q����/�鄺����62�����!@A� b5FFϴ�����CsL9>�K����Pް�G��7�� ���#����#�6$��`���h���^�}� G�7EDPތBJ��i��^i�Cx����zX�媘�4ϩ̳ٛ�$�� �������q�"M��f#@Kph@]�d��2�6H�=�ڐ,�U�L���Cm��p[y�8�u�G���r }���("1��Dr���K�E�ExB(���PC&+�V(M��!f�����n,���M'� �#��^�����ۍ�u>'�RC��.)P���%r3گ��W���N�����M]��"6�e�,Qv��3������B�d���}�GB�������_���DY6���<]x��tԇ2�||�c��� ��{c�]c�}f�&8�q�T�E����G1EF�Q�D}���}���LJ��4P:8�	�X|˟ނ
���DD����!3�0PD`��#c�o���̊hБzLL�x�t%���i	2�`Z�q�H{ʢ"94��qᐻ�z��#�q�������OCߨ&���>&�p�c�(	ˎ��Yc�u�B6��O�LBz��!�6%>;�y*�Q��m��ڃ�$����R;�_K�Xš�z'���'�yy�Mi����ա/d����$��@Qi'�p6�^r_����=~>�9h���s���#ǰ�X2�oޑL�K�$�k��h�6����KE��Kۤ6@� ��,�`؃�:=�n�3D{q�6$º�}r7mf.��B��,]3 �� ��/v�H�����w$S�	��N0