BZh91AY&SY`��F�b_�`q����� ����bE��   }�ǍV�UR���f��hm2�Kf�)����Y�%�m�UVm����J��QCZ�kI�ɐ�В�(��T%R5��m��6a��mv�ګf�Z�k���Y��6����ٲ��Z�6ڕkiJ�"$lٲKjiF�T��&�k��-)6�U�jֶ�iZ(�S&����'Fm%�����:���k"ۣ���6b�Vִ���l��Қfa*���#3#Vi	b�eklYb��ki�Ҳ2©��A[1Z*CP�U��y�V�U)�    ;����;V����ޭ��۠6ú������s0�k�j�:�tt�B]Uֶ���ifwU��&�T�Q�v���t���M���YJ��F�m�{�   �״[j�*o���֙T�5y�.z�)���JJJ�d��x�ꥭ��)*��+W^�zU�U���(�kޥ�H�(U+�{�*QT+���If��3ml��dԏ�   �����jRKｭ��vҕ������\�T�)��{��]��^�O��J�SϾ�y$���m�c�kn�^���UU;e.�x�P�R��ܽ��n�q�Km����2�͌�!)�  ��*R��Z�;���%U{eY��xP�I)�����@��瓻ڻikR��p�٤��vz}������WxJ�
�����(�oz��R��]�V��VL�Kmm��j�  �;��"A_C����$���K��C��r�u*�JP�{]�m:{s��{�w�U"�]��ǅJ�E@lvʽ��n���(TWyʐP$w��U���L�F�MZ�mπ  =�2Z+�w���jQS���z�l�1Cz�x��T�î�JT��]׭ǅ�hz�׶�eH�.����x׮�*�����H�I�pP�R�9=��Z��Ai�6�f�2ma�  :�ϱQ���
�y��Y�'�����n릩IV�����J�-w��xP�ܭ�/v꒭��9m�Z�U-�p��ל7[jhq꼚�VͲj�dٛdٵ5[Y�  g���V����zz7�j� u�:b��h/#����[w����ЁcA�]�^��W��۪�[�m35a�ղ�[E����  �o�T}3�V����F��zx�{+��{\��c�z^���zz�UFڊ��U��n�4x��oJܪ�M���\�Tw���e�Sh�I���Z4k-|   n�:�֊�)�
g��P�E�x����Àz)�{��T�lp�:t7����8������j�/� �  L�%U4M   b ��1JQU@�h  !����R       E?	�)UOP�       �?!0�T�&�hA�A4�$�J)4�bi�2M�M�� d4������F��9?��)��w_b�ݟ[5��/���ߏ�����6�OǾq��� �}������m����cm���N4�������������l�6��!�)U_������6�����;c�������������pc�g Y�k �vÝ�� Y�L�mgm��k&��6�l��Lk!����m��;md6�m��;��� Y ,��6�p@����Y��WcY��k!�ɌY�k&��mgY��CY9�8ɶ��,�v�0Y�eȚ� ��5� �Ll��;�&D��,�����Yc�D�Y���6J8�`��l�`œ80`,�	��&��" `���	D �`�v0bɶ�$L� c;
`Y C�0k&�!�!��86����Y6�p����m�� ,������82�Y6 ,�&����d�Y6�q��d��5�mgY�k;ɍd6�Y��8Őœbɲ�D,�k!��md6����iH��A��ߘ
4@���������}�b�4�/0u�$��4��[�PHr7lQ�o���Z}�m=��.��ݍ"�U���޼�Y� ژ���+ƛn�3��頠�yx�7K�,�e�2*;�*Հ�s]��r�72� [od�٧�q5�Vʹ�u ���+��:�@kx�mԱysoool�X�E�F%% $k�G>��R�Y���HQ+�E�
h^��[��n����4�w��Z]�ݏ@��ŋ7(� Ke�ASsif�^��XC+�V���B��j��R$�[�7�4
Z�P{xD���Sp�^Ex]Yb�I��XBf�q�(,�[���Wh:֯1:��{�Bl���+�!�*B�3f@	wY��*е-.�"�(��N���뼗&֒Xu�Q�1��/.�h�A4�m3�E���1���\&*:�.a�j�G��ۓa��9a*̱���-ȩ�2Ф�ٲ�~�h
Y�&�c4�[*!����n(�k,Th�]�Xo0�2��W�`݃6��摔����qc*�X�5^�Ϣ��V�]aM ;ܖ��Rս3]�����cJ-.6Kݺ�W[��DaMR,cc�7w�-u)e֭"Y�6�t�.��3r�q��N����X�A$��w  ����J9����t2ҵ3���T��<:�)����\ܖ2�[٥֋1V��a�ѵ���/эhP�$��Qt�/��N�~8�"�v�x�v�]�Ҵ8!
L&V�E�&r����%C�1�K"���T����n���I�Ne����[��un�QC�#`��xlRU��^��f^�-Z����%��̺�vVZ7���R3[x��0r��RE�B�����їC[|���,wE0�V�m$m���!�y-�����lM���#CmCA�ܭ+56��i3hSݥx�}aeE�svḓz�4�{,��]f��a��)��5�S��)� Y�񼱩Y�z,���Z���0]1tl���[˛/Q�M�	����^�u(��e��9�s�![��k���N:r�`����/e�K2��uB�۷�&rB\�Y[�kqw΅S�@� [bӾ�.�EL|e�3�V`�>�2B�!m���G����rG)`�W�4`�v�2��q;�&ɠ�A
��_�����e, �Z�������Heb��ڭ�to.���n��R8&��<f��N�	�.���6�.����[p�4��2n3)E�WsU7Rf��@!5xo�W�SO\�zkt�g2��K-�u��I)%�V:�tE/6�]�&���c��s��M�M�}�wB��2�7KPX�BK�C��;�Sw�v��:��(��+75�b���j�x�X�mIzQ�͢Z03�f��CU*�X �륶����m斖+z���U���Ū��ގ���F姀�!�*����2�y1�юV��߀r]e��h�72;.�!�s-�$Ӭ��`"Y[�d�n桉 E�&3]��1��IV�5�V̋�A�w�Y�&� p�z�^ՊkU,{����6mc��VdhM��+�1nc������x0(����Yu���*p���a{�:wS��.�-��%e
��n����Y�/6�r�F��i�IL��jű����̦��+�t�6�56��,��kjjM�M��w;����b4�5�E�#a}� .���d�f'�B�mAu����L0擬Qgvƪ��k�%P�e�L�YB�&�5s���{��K@����x����ؙܬ[y�PRъ�ll)��-؊�:@�p��g&��x1�ŢV˔�Z&jlM��en޵+v(˨��x��.�M0��^^�b�HVD����lh:\zҔ٢�6���I|Ϊeե�c�ݍ��F�&����b�l8���,e7�u�k,�CO�Vtjlm�"f�>bf��7�����{b�
b�[�rfVd5��m�ܓ71�L��t�m!K+)��W�WV��n(M�1�]ݼ�ZI�tB��p!���]�*�A�6orXmPssEdq'�KaB�zZ�EQ�o��KV��ѡ�ɧu�HE�wj���O�r�+�$����
É��E��7f�y�9�abJ�Kۣ>W�k9e��Y�˭�fSɸ�7w%�dԊE�f�Y:6��MR���u���D���y�ɺĉ��,m��1�v��:�He�����`Z)1�!��_!X�����on�r�v:O�1�����W��k�^*)ֱ����� � 4-�c*��1���陲��V�3����5�@x��w��5����iؔ��*I�SG�^l��
�*7QDm=!eZ�ݸ��5�e-tl6�1 �z&+b��m�DN�OK�W{`�! ��X�n&�]Q0hLe<�gV�.��޷�e!P��U��74\Ɍ3����8(��2aa��==b7�ij���vn̓6�[��i�eU��/m4�Uܑ�K�e]�F���Be7E�ܺu��	ߕb��[hC����Z�1�Ek��L���.��7@[u��ꫭb��τb�hbr�jK ̖�c۳h�3빴º�Y$T�YHc�����Eљ0V�3Po3eL�ln��ek2��馋���w)�T�)Kh�
L�,���������X�t�]M�Zn�-$��4��'4X��m�4��ز�6��+\� �ˌ�x�m�&]�5a��m�4R5�ݬZ ܸ�Ӌ!zf�=$P��ʽ���R-dM�zI��̛��#ƶR�Op`��.�SA�x�ⱴ��*��F�j�	a�$���@��)Z��T���m�E<Cˈ�6ؼ%(��!������/VC�M�Z�N�� ���Pa�ؑ;�A0NI�r^ǳQ`n�
�U�n�R�[x��!��-�A�:��m�2����:�T�Q�uz�U�Iso��u�k�MlǪ���n��w3rk�[�ڵ�P���koq	�ɯY������)
�tV*�Pf���R,ŵnU��-�� X.8Vl�t5v�v��U��zV���"gv���$siV�B1+tչ�`����yu�Y���fӌ��w�l;H]��@<ӡ
�57"���3Sz\43v��<�mk�t&�:Bn`�FƑx��ٵ���76<K&�In���Y����D�t�9��t= cx�E��2�Q�0��Iӕb	m��Xǩ6�ޖ�L�%[��4c�Xm�V*�J���:1,�y��f�u-�[�Шn d�N������fA{�3
�{�18��E諴v��&#��.���d�M�z�!gU�«5v���q&��Ma�+4	AKD�
���ܹ{�������7��+�M�=�ӮM�w�"dR!lX��kv4f�éhp��D6Y���m����u�Z
5�4���85���Y���)7b�ELl3�֡�n��ӣ0��SH`�s$�Q����Z���bH�e�Ao��/�)�lcy�ZH��kOt�{�;�3��KE�f�[�h��z��Rl���ӷw��7BǓ
Ui٫�F=�2*�Xcљ0L��b�7V t�3��1�l�u=�@'KZ+8Z��%`cq`�����V֓	˨��,�gvj�T±6���o(B�c���v��lY�ǀ�qљ��h�(���H��Ff�o�>1��Ip�Y���e<4G�)�I-'l��.y��vu}�.rٔ���|	�a��q\*�Ř�42�U������h���A�U��}�h��4�[n��H)hB�E�=<�+l7E�޳W�sX�;F�y�v;{�2[`��QQk�-լ���[�4�܅͹��4*X�����{��t���oN
kw&�L�I6�76��,b�×F��e��gαV�K��:��2R�^pԂM�u6��L!)]^��� 񵉔�+DV0�l�"�.��v E
�V�;�j�pS:�P��J�1�X�7���RD145eJ��JP` �z�f�*�ucu�SU��;yfe�n���^T̡2���O(�fr(�H[����*:^�%Ƕ��+Ua1#�0����0�[�v��ert&�h<���cv0��%mZ�L�Z�����7F�/�V+ME��C�\��3CƬQ�4�i�ƣ��J�Ò	JQS�O(bN8��<)iX�R�bb�<�i	y���[ub���B}{Zj��ٷs]�ݲ��+0}nTie^��84�b�jf8VSe;�F��kJ���`d�0�4P�XŘ��/,�O#'�����0*7��6�1�$��:&�uPYx��}�3Z��=�R��Ӭj�%X����Vd�B�y��/b�U�5PnLЍoՄ���tu������е0E��6�V�C	�n�*�k�ծ�ǉX;5��ݛMӍ^�U���e,�keY�lTSM�g7T�32%���f�w-jtȺ�)엊�k�^��kb�y��d���dS1N�:����o)���ʅ�
:ݚ�U��qY	1W�x����"���0��ǟa���@Aܫ(�E�j8�1x��x�obu�7��$oQ��X
���n1jL�m�n،���C٘�u�[K)"tp�l:�����amfeؘ�* /tlǍ�u0-����2�ǵeD�993[��6�ܲH�8B����Rֶ�=�45"����)˽!��Qۅ����N�&(ώ
9��\߯J�#	Z�f l��y�3W�,��=F	[JWMdc&�V�Y�q�x�{���u2�i4s��13u��Ib���m�R��Κ׏d��5���	+m-��B��:r�v ��`o���v��x@�ioKm����K�_Z��:����ih�E⺱�c�y�r�V��A0�2��ō���!*�ZA[���\�{4P��)>T�G���Yv����TЎ��t���+S$�������RU��y���ӿ�ؠ�l�.���٢2�+f<r썓+�a7�6����C��%fM��n�S�� �n�j0�����'�ea��J���n����YTf�m}qAG2��ՠՍ�Q�)$� �ڽx�{l��QX��tH��T�cj^3��7ʻ�Xf�,�je	�^L.��-�m�f�QF�mZۡe�[�!ޕ�`RKp0��l�{:�g[�Uts6lj��Y�Tʋ)zsdp���Z�ݛ����b��Aj7zV��srL(�Z����o$�[�v�6))3kj`�H!�Ի;��3"�PʕM�.�$�j=��F*�����PIL�����.�*+CB9�LV�H;d1m�̧�1�d�0f�v'��m��]�(��w�jXn����)����c@[-C�NZZtM���X�1��n9��(����^�;E�6	�>#�F���P��4���w�Gi���J�kbъ@��7�V�Xl����LJ�E�0	����oT�*����%nY��-�ڵ�1�k\�1\I�E�t"�YN-M���u��mѬDd����U�̶���T�7C�X�n����[�B�07I�Ӵ�va�K�x	��E�0eQc�4�"m�DP+��*�A��k]m��*��v\�o[t�%Ǝ^�O�-�Y�����8qҚ�Sp��)z��q�m��m3�<I�!jv�Z-�f�Gt�B�Տu;��W�^zjV��Vu?�iI�nd�Z�;Z�D������M]�Ȩ�Õ��܅��Ҕ�y�w ��T� cIl�KAb.����R�[�^�v�3`X+K����RS�(���\�U��[z���0�j�S���i�3CE��u�Q=(/�#�Wn�]d˄9GSXͫ�E}[{���*�M�c�x�
 ��(�B��n7n��T�R�kiPе�K�`�+3Njn=Bo��
�-��Hڋ%@�[*gp$\$=9����&:�Go7[Uu���jJ��:�cץ�9.2�$K6�n�Yp��.2��%Z��w�f�E�yP��ˏ^Ioq��IS2�#&j�k,��.`� %c�j%b�q�(������{�i�1ʺ��kfed�I}eo�6�9�
�!T��v|�U�ڦT��ձ	Jf(�6��Y������"6��ҝnG�]��fSnVƷe)z����d�x2x��U�5*�H��H5R�6Y���mb���0��@��w3��-��D=I�[oM4K��ꙏkl�R�ef$>Ň�'M�W̎Ť��!Ύh��F�Y���%�NZ�բ�,�&�@�e;��7GdO �7�G�elE�4ɓiS��E��Z��;	7�B��د+ �5�[̰�+/2<�����KmK�6�,��&�趩MZ���@��m�Wq%��B���I�h��{���,13��0��Zp-���r^�Dh���0�N��S��%3� �/&�p�z�f�D�V�]�Ѷ�eHtF�n���a�x���%]�$����O��bm]��sh�:�S�X5���ɘ]꥕˫��t��������kx%�=?h�<_gph�H��c���1-cr*��5z$BD]�4�[H�m-6wd����*�igҵ�t6�ؠ� ��b�)s��Z�F�-�脫H�W�t6�Ey�YZl�ZI0i�Ŷ���egخ�^۔�.���/��Z�+^;n�gj�,dU�ڂj�;a�tѓ~ͼ�4��~�4j�&�N�"�R�YY����5�q+�X�*������Ov��S#W1��b�]e�X�*�ҳ-�,X���5�������b�j��Yy��L�iSj���ЬC5�.i��@K*b
#���+r�$�l�YXi����u&C �m�I:�GެY�K�&���2�a1�܏mf����1hW�3�r�i�d/
�0��Q���V����4N��Cдr�HZ"��v��<���l@ �#�U���,�Fi�Я��D3���c=�a4��dٲS!�/�ė;�ى���*�x-�HDX求�{K�ܝ�ႉU�P�����?���M� ����0���J_��3����}`�DV��� -ޕ�Ц�]�-8T���]��y�b����VB雽9Oki�#V� .�iS�<�k\R�n�g�~w��e�Z�l�y��<��λs�l��ko�ȅ�Z4O�r�i��E�̀"�n'���/��B�'bE>�n���(k�8�[9hk=��Y]Ew�;�pf�R�֢��+���y��v�bNNtpQw�R�+����F��dPC{lV(�\upY7	R����vf�B+S��k���|j�.�\���%�<P�(�KB����YOc�r�	�$4'�'Bլ/�kЃ�V��YC7L���.�^��H S,W�}�n�W\3u�od���v�ñT�`P�ݻ�r.*���2�E�׻����7JNW�jW��(_]���9����D�vG[����F 8bj`�gL�����-8���^s�
�����X����3�)��zT�7O��\O`ݰ^M��*}�;����W'O����j�R��*w�����<7y�5G5#(��9������!�*�p��Y��R]�9L����n�)>�kT����X5�K�yZ֊&����3stŹ|鮩�2�t!c�&J��F���L̓1[#b}g�E���]uB��T���9�o4[5���Hf־�#_=�	�OR.ԋ����x�y�����8�f�(�C1W=�o�4ʳn��&��T4��B��Vm�&��hU��ڟ�
�o&�^R����݊�V@��J_7�bU�r8*���a�P�Y��k�}F�m/��(bY�E�i�c-��cn��V����ͬ2��_Lq�3�O�$��Y���?s��N,�)��.b�[A��_VW"-˻#cD̸�K�ɚ�w������4�;,�֠r��T�u=��]�6K�sU�koFATg�i�97�7���A�5[)Q��
V�6h�.�m�İ`����\�؃���1[\�v������PZ�1mp��+�>�u��ŗ:!y�G^�
��4V�oB�PǬ=ѳrh�ϐ���Ǻ��x{�!��ȥ%��Y`���fUΪӋ��MS�q�S{z!ugJ�)2��4LQ�A��-rV;��^6ޝծ��m��]�|kYP3uۘh��Vɳ%M��U#�g0�z��D�bTPYK�<���/��#�_ek3Vo+�{l֭�fmB+N�ss׺��֖��/c;R�Xj����]b%�C3�M6v�M!,�sZ�J��]6e�CNOM+�L;r���(:Q=���-��kk��p���k�ECe�I�9�U�E�����쮧�1n�(�xMS.��W^��ݖ�R���'�@E�VJN]��pπX�<݈9)����Ƚ���C�p�«��Vdtb�]����IJ�wt`޽#�&�x��4pͭ�7�,K�K���W�&c؂��n�u��sxX�E�
�I w]�3�ouӌM�0��aDs���broU�OEk����]�L�B����ys �̤˳A�� �ݚ�.��Pn����kxؔ.R��BwR�SP����9����R�/�5W��x���w=�L%C>Z���OV�!r[{sm��ho{�ǌ�.ж��nu�����xn\��u��܇Yv����5��͙���섞��]��PI�Y�:��c���؜��Za��L�3Y �q�uQ<�D)�:�V�ޙ�����h�{q��k�%]s��vC�U;�F8 fnF���+d�oAͨ6�|�y�c=������%�n5ۤQ �)�8l���������K�ҝ��T�i��.���,B��գ7tӦ�m؈�a8����V�|�10�P�K��F/�ބ�4��)]v����z�8�}v��o��������[��k[(�so��\��-r��҈��כ�q�3
����n�n�&F�2b�}��œ���%�RnrؚnEs릺�<�KtSO��XD5�>R���"�ψ�Ǫ[��ڨ�
�W�W�N��^�T�v�Z��h���X��I&Ӯ�M�w�2�T�bꎩ�*��c��t�j�r���k��;��9Ѽr���ѳQ\%�s	J�2z:=7N��f���S�&9˻y��R�cࢠ�sYҩj|��j�9@�> ��\TgvӤ��|��ԡ�PT�*$N#��m�#��cp�K:��s9<���(��m�9N�<ּ�gJX���nK���ʚ�=�M3��V1=�sG	WݚtbS�|�aj�@�v�^��;.���������<U�.�n�&0Ϙ�S�ʂ�]ԧ6��B�X5��ǰuf��&��V�&�+o(���;������A�#�<lv�=��-G���w�"��_�Ca�G)8Y�=N���6S�����k�ȹ����y@�@[��X;m�|:�kh��^��~즽��廲���6��"w6�,�����.Q�U�,���L7�O9=۔�SXGnHjY���N��X.�g��@�3��;d�,IYr,g��d�]*WhJ�w]��6N&�Ac�łb;9�X���+���e��CN�%Po9k["1��I�c+L��z��*=X�Ȭ�դ�8�����!�<��ʣX��E�%YY�K�&�"a�څ��X�@B�إ���;{�.rK�ݔ�eL��CL���ګ���Wwe0������f����<׬�T�yX&e�h�,.�Lƹ[��J���a\N��P1��U$E![�YE���k��b���B��b����`����^$��:��h�ybt��p-+�d۫�txN��ӻ�ڽ�	���VļS��<��,a�Q}�A�el}�����Yɹh,��l:6e�uo0�],�P�L%Pۡ�ve��i��vVuś�
z�q�t�39\  ی�ЗL���;G�(�<\?n,�=d�̆��׹����E��|�s[�q��֍C�]�T�<���Z��򚴹�Ne������w\���EՖ]���烱�{�cb�7_V��;).5�B�Le'�v�95L2��e�v&�+�b����!�019��AG��k�����S��k��8�޳�:n�7Eu�16�~C�wxR�-���:�7�0B�'hM���eՕ�W0�x�]���h&�ǰRR�B�ƛ�J3'�3�,��h�#�6���٩�8/sh��h�9�ǌ�6�X�)}b�C�������J.�����Nu�U�L�A��z�jC;'L۵v�J�t�t�ԯ���Y�]X)�a�hЗ;�I�Shv]=�Q)N�}�H٧�z�>����^)���!::�tc�DU�#TgCw�%�82�z�4�,h�D6�vw �\�P�}��[�]ek�&�����U&�^�v��gy|����̹�i���`S SuN�q�U�N�N�u|�Eit7&U�����]=jR,lr��:�ö����7D�'�V�)����BI��X�:�ƭ��G Ĭ�k���aD_�+]浞����[R�w-��SN�*qǝ�K���"��j�+!��Q�"���{Ί�F���}����n��y�2��-��e>X.c�iV-)RV�̣S)^��r8'f��Qʕ靓�0%�ͫA]W�%�e���W��J��"z!�߲Cչ��2�Z�m�a񊍱�l֔�$���p�ǯ*1����h�2��@w�xV��V��M�$wokK��GpL�i��qB<YM� ;���7.�p}��us;m���wy	.;틓�lU|���F�w	�o�P�R��Ҟ=;&��	WuνÜD����-����'To3�T�Y r�#��uk��t�M.��P��-����x�{�����Q��ȉ�]b�ʱ����
8ZZTV�X��,N��^�28��Pp	�n]��L�;%.}��taQ�-V��
;Hu�sj
��T�e��W�`�lT��:�
x��e�ɗ|&�� �bQ�͌�� +�c��aFYu�ĭ#��>�
�s,@����=��*;ͼ�y��Ӳ�"2I{v˂����u.f��;����YٗٻYg{Y9<�$Դ��(�o���fhF�ic�n��wK/vvlH��kB[����c�K˴E[��8/9�����Z��-uCX�X�C�8���ĝ��x�G�T9�T�E��X(0#�Tu�\:��B�'�h;���ɣ点��TϦ�;i�I�`�������Rj����Ө�	6%�u0tk�[X�AMΩx�/ ��R3J�V��֫�-�6�c&�r���F���L�5�f� �s,Ir�mq�N��u���K �H`�x�����j�����_��C�0ާ��=�]0l��V���ʷ��jÏ��/+��C0d=�&�Q��������q�+����;�B�*Q�*V�86�%}6�SS�Jr�B��{�i�#�d�n:|"�Y��Ojz�	�4��*Kz�Cl��kna��)\��`�ؐu�-ۡ��� +_ٲCS'|nG�V�Bi�:#��B��:\!�8�Y&�K)l�fo �W0n�m�����P�]���9����Q�ɏ��5
JRc������ZVeFen��u0w�Q4�-�7
z��Ӡ�V�Ē��{�S�+��V>�S4��ݡE4��ӌ"���$���V���,p^������3-�+K��`��x�ݴ0f�� y�t4��pl�p�J�����������u� o:b�T"ܣz��Ї7���Ί��*���&�ۣS��8�����3j�gmX�B�^��K�N�޷��P��yW�V��ux�{)i3u�
��@��N�Sn�k=9[ݲ�1(���Z��u>(-�:@��=���C�Z�vCq�ʊ�+��qne���72l<xJ�gs�v2�kTX��-F�L�����F�_'ֵ�w+xX�B0tWIIچ5�4-H��z�������������d�a<}'Z���M\�E�c;�j�ͽ�&�ss�)#YQ;�|����p�"��=p*p0���V=�c�`:Yr�p�ޡj���Ӓ�';B9�J�	����3(l�z�r�/��5�G����<=�b�i��7�[�{[e�#lAIm��60٫I����)Ht����#ǎ'�fú�u�͢�`0�̭���	��h�j�5��ʁ�[�T����e��ޣ�yY�Hf�_d]ф�V�Ig��kN�l�N�4�Q7+-(8��fC׋�"�AYjR']h�܊�s���1�VOh�6�7�q�Z�76����K2�ȁ�h�N`� #N��d}��:��L>ќ�L]`��*����j�o'�CWh���)]粢��g�]���>j�v����sE�6�ꡘPò�¶�e�۷�+V���&b�+s�2�q�lrӏph�Gcµ�(�n�{[�VkDe�9�H�s����_2F��"�<v<Ur��َ��rFs6���h�,��9�[W��.��@kSAɚ�Q9j�}�o��g'o�>N�ۍ��85���!Y�ٕ',� byR�"4ԓ
!�()���G�,��")�,�n�:8�rC 9ٚ���Ń�Zj��)�e)���\�l r��8�����^ջ&�]�6U�oxP��[eu�[�`�������$ܩ����"ߕ���:m��I��q�u��ɟem�)k;�+A��ɰ&�<s�}2]0��  ��Ok��1��.W	���&d�'AܱᏩG�[��}���8X�k�Cv�j؋�9G����-��׸� �dZ�m�V^��CL:�����+�eSx�D���&��W&��NN��C6���̚,�I�-�k�����DH����W��EV�Faop]n�d��8��<ZKS7��u�|Tέ=�ݑ�i}��]���l�B��ɝ7�56�s��P��@aƻO&���D]I�
<�7��)C%D�0\ V�u�ggc�*@��h�`ܒV�i��-�����ɗ�I/\W���j9���G
s�i[��V���N�3ԍ��Z��bd��A(��f�b��p��#�x��pTej��-5� �e���dNѳҴ��>�P�ʛn�OS���_c�.�߭!�!�4��z"im:�mlen��U2幗sJի1,K�ۓv^ݗ"{*]m��b�Ү���U���^��t.�o���3� �t뻋\.f-0�
Oy�\-c�՗�r����n��ѝLV������/��]aE{k��|�54���Z�k�f�����s�k(�NA����AN׍ɗM|�i$3Ҳ쩦Zzk-ɭV�d�I�]Nf��GwfR��;nY���>l����X��{�-r�!���0��J�j��׳N�Ջ�b��L�
�ں֘��n�ɋ�2���.��WJ�ҟ m#H�Vb�i�Zl�'bTh�S홆�d=[��zSf��8c���]�4ɢ��v�̣S�7mu��n��3s�5�`+�9cn�n�$��Y�yF��LIr{����ﴻ�m����oAHk�r��s�3�ֽ\��4{�AY}m���?
�*����w�y�K��	��+r�H{7���ջ�{Tt�9�)E�&��$ٷ�+���p8:��>Wǟ']����0��]�-5O)XJ,yq�Z�����;I�f�6�ZwW"�$@(��(`[�Q�4�袱)ԮV�u��J7��&�"�����b�	�I��t7�1 *�	&ª8�qͼ�L��S�^���؇te��b!���`;�<����f�I&��2d�I�d�S���"�!QJr�ݕ��y�]��y�V	\��;W6��df�7|��u���Js�8b�OJ�{���}�~��ɂ@���o�`���o��ɏ�m�[��6��v����`6������^�` �������g�c���?``0o����C�������?��?���_���j~O��~_���h�Cgc��0S�Օtނn�<v٠��r�E]�:���mb�T�u��R憬�H[�ܡ,e�;7@c��S	���ff}��;WM�u�:" <s]7Y�K۔)(����Ŝ4ǛJ�v��j��T-�K�w�ѳMZ��S��S�����*�Vuc-���\����ǈ����++T�Y��w�����c�#�M�F�_$���0K#�9[�P�%��7�"�ͻ�Ë�,�v�7�8�� �IZE����e-�U�mT2�ů����4�����u*�����f�w!4��R�>��'/K/�דU�cV�@���w�����ut�[�̝J���y��7�M˷�Ԍ*����v!u��b�;��t0
�3��4:��JZ�ud�	���.�nS�i)�Gk���f��݈L����b���n�[������s/�d�k��N2��,��ayG���#b��J0��d���BuuyjV�ZPťNs9�����9SC���=j���Sr��vfv�9(mLM�{Me=��mu쨜w��GSvu���B�j�1���r���\ב�Ժۆ���Ӛ3�D�V��l���
�i-.C�u˴��QX� �Wf\V
],E#���Xݢ�f���2�'���p��#t��gw���3}�6�[�9��Ț�$���~o����~O�����{���w����{�ޯw����z=w����z;�;���{�^�w��������w�����}>�O����}�+x�j��丕0�N�f��	a�E{�p͢8V�9�&�+s']�V+R؂#c�ް�X1�u�z��X.�#�w0�\j�KGuF.������n�ᝳ;^ܤ�����Ful�y%Z;`53��YJ�ɚ08ή%u�R��W'y�V���/1���b�b�A�㭋�:�>PQ�����ܭ�,��=�š���h��K��u��:�Y3�.�|�FU�k3y��9�_`��@��b7�=i�R�d|4'�9=��5�e��YV����m�ѷ��gSW���s��=�C�!&!�ov�{|��ڔ�f,hH��"N!=����37�;Ǽ�c|8Rċr^uJ���.Rt��d=�Ek3/]_���Y��w}�q?�u��&�ω}κ�f�"��Y��*|�٘&��e=�� �<߰�h�Zi��6ᙦ�j�\gw#c�S�P,e[,?�d`C�Llrek�%�R�o.L\�x�*�����H�Q��ǉ�U�>�ͫ�79��t++�:�Ԥ8�î�v�9Fm&�μ��'��W 㜩�-\�!CW�̴�x9��n�	�J��m�mPz���Hu6cN��jb��6�U��
�rT�����g-+��Xv�܊��7�ֹ�����C��ևkmt�V���]X�Ĭ�����i�:��s{�`�V�+�V͉ZJ|L��yz\��j�S�*�5U��C���Ҿ?o���}>�O���_O�����{���o����{�ޏG����w����{���?����}>�O�����}+���}>�O����S-'N�H�tΆ�G*M���%^�g���vru��%>6�9S�`De ۡ�wÏEl�z��v������g:��YMu�q0Ů����>E�� �O��v���n�R܅�c*�
�Cwg�fMP��tj��璵Y���y*J�ݬ�\�ڂ�_S�PB�W5�PXuݴ�W$*��s�mIءWAgEe}+UP�n�V���R���F�5��T��YCi�"�ioY��&����VR��q�����
U��:gN�tdy��t8��%[�/Gi"]r���ch���q㥘y7ʊ�/h-I��!��9�J Kޓ�r��i���Y�Y�o���0���a=���:�[��ahgI��9,�J�8b�F���hgꝀ��n�U��(��U����63�1�m��s��jJ8T2�4щ՛�g5Wd�朻�QU�}�uM��8��_qb�9l�@jÒ¡]x��%[�%�@���o|�;�r���f��p��ak�n6oH�0�r�^W*�0(��;4(f9X5⿑������nP�z#��C*i��;̜��=�[�����4dN����"nSC�\��%J�+�AX�Οӕй!=����b�3(����{�����ջW7+�2�����oM�#Zf*AT]yK�ݏ^$��Tq��E96�3�gܭ�x���[\���N[9;)w��Vk9��>)*�+2n�6�]��ä-1c�
��,e,��R�]9QB�Yn/��}®,�w��U��v�5��� �v��� /��Q���q'/9�n3:Ё�E<ed����n`�`�M;J�]��B�wɷa�_�9�ME+fI���a��q{�aWA�ߞu��\��f"�)�׊e1'X� [|ݻYE�9��<qE*�]���8L�2KQ;��C�BF���P�4�t�캽�Ӕk]��P�����v�J���V�`�v��D3o{h�����LW)#�Fe_#���fX�m�m�AK}e0�^��z�F%�kd&��W;KK:�Y�n��G���8o��p�}��кG.�����[��!SH�:�����VB�J���h׵�QO�ﻣ��gWP]���b��m��+	]�L��r�U���˝Pd|˙o2l	]w��̨{k��k ]q"���;{�\M8%�^IlNե�w��]CM��K��*�i�n�,�#�ت]3	#+[��m�t����B�98���jT���1d�m��5�����[��CG�l���F��vd���7:E\�4w-�ڃ:t��<���N.S�)�;��c�C�1�
������;�ԝ��y�E�K��A�����=+`���1J��f��4B�3������-�1�-<�i��"VE9�W�2]�_%��
�Ѥ SK��}C�L�uc��u�|E��nv��k�\r+�*5�Ю��P=��7��p��mu���(WS(�S���G���\�],�xLZ�ȍ�z�'�ͫhބ��}�]��51��P�z�������%,�����a��W)+��+e<٠Wm�J���TȮ����S�c�r R�pꗤ��� '���h�Wn�]3���Ƶ�zm����|�R]{n�e�Q#xV,�޵�_�qL�A�6�To�{yV-e9��=qw+�O)s�I�ef:X6F:ȩ;4yګ���2ɢ��W;����E�Qs�6�$���;Z��h�JE%`��KM�rN�t/%\����W0f)b�
a�S$���vc�F�ھp,Ju@�) X�-
b���J Eٺ�%�3,��)�
�(u���b
��s���+�9K �|�$�0�{w !Z���hr�tH����v6�@6����=�/3�Wk�B���;��[�7ݸ��+(V��r��T�vJ���0]8e,M-����u���G�B]n�P�4�G&���]5�覃e�xՒ��ۡo.<�W)�Nq�KU'ZY"N�S��+�;���L��؃�vJ��Q�GK�P{�v�K�P�U��Wu*W]'O��W&�>8�e��k �5��o{V����%��m�#XyD��eM/:0�$�c��̷��ԙNp�h­az3E��<#u�y��`���P�`VH��#u��.or��9VB��A����C�7K�j�Q���-a�+��`�p�U�㹂�j�Z�f���t����IC��y%2�3��9VS"D[o����������q�R罫0��͡��Fnn��oU����|*D��Zw|���q�LIZ� C�ҋ� *j[���.��y��{�K쾚���Ԯ�Mn�M&u�����)�:�h��p��)�*�8vB3^oD$9�d%}�����
-"E���5��0�w���U���$�g1�i(U���5P����4&�x[w�6��EWA�m�ۂ]�ǅm���-�S�F�5ۙԓ�KM�-�O00iu_Յ���[�Uȳe�V贬�;��S!+^��9�7r	7��������2����s�԰��h�v��ࡴ�%�	��:�M�Q��qb���I-y7%�����%ݓ �@J.��kDw3Zy�*��ݱU�m;�MH+e��NW�N��3]�x��˲����E�ʎ��NK,�w��º��Pަr��nF&>FYE�GxͭPɪЧ�o�uI��CE���Ԉ#�S+���+]4~��"�07U�g��g�x=h�':�}Oz����BP�e.�>�U� ��.ӌeĻt� �Y��s#@
�4�p�j�\�-�̽���I�'�)nB�|����t{6��;Yu�@�`l܍�GY��W�������y#�wItAw(kb��/�*w�2��[��:;l�B�x�^�F�Z���»�����[}��44wV����e��vIF��l�#CN�X77�1w����։�|�V���K#�u�)%ι݆�E��@�fZ�ӥ�Y��A-�����m�d��W@i/�	�G��U�vgk�\��,���HF�:�#�3��k�t��%1t����*U�Ǯ�d�K�W]y�������5'j|kÜ�ps�1֜�o�&N}�.�k)LU!�cN\R�����yvol���*�b�ΏPNu���:����(9ZY��.mAt��S�iMՉ���ܗw*�Vu���p6�jt�LBj�\hm2�Ͱ��}��J���:#366���^Sn�u+�i0�3�� �%�+s�;��n^D��WA�;\�[�Au�ˤTsz�ӣw{YG�ZEk΋G5�/kQ�+�@Փ���W
�q���VИ��gHR��ٺ�4nbaw)I�y�m�q�8�yH�<0T;Y3����2P�UV�3���6���/P�Y�w�*���{�ٮ�o@'�X�a˛��͛>��$"���Pռ����[�����'�M��QW��rޅh�؟.A�s�v�uD�����&I����%�P
����^�m[�vd����G#X'u��%R0tB���2�>kzp�D�v��C\���H�ߥ���V�˭�]/	��i����g>Ը���b��\���h蝑^��\	�pJ� kA8Oq649I�� �7��ׁ�W�n��yGI�Y�H��5x>0s�L\�ѕwӻ��"o�����Ik���G�@���Y��H��s L�#�gjyXܲu
U�c�c���
fpPA�*K���}�;{�K6;?u�v^4��"[B��n�I�#m���˽Rrʒ�X��2mFТ�������^�\�rbC��k+k7pZM��9��R�^�`��]cN|6
�QFN���b�p2P�.�f!�F�a��l$&:���ܶBVsf�W�t��DD{wc�6��������t��f��M*짫���imoٺy���Ŕ���ſs��,����G�k�~|F:�v�ə����}���M*�ǮJ�x[�`Y��z��p&��uӕX0��f�.l�A06r.�y�	�Ӂ��n���w�(t�S����D��\�
�y��]���Z�#+]:th��겭䐝�̈́#�V�}�4b@�����`I���:���5�;m<V�Ge�`��*!���lAڨ]���Fƫ�b+��mi&޵!�e-%������/oqɃ�'���_Dݶ52�u����4�[�'���(<)7`m3�8sA�˶.�O� �X;����kD�#���-�K�D�fP����j���������:K8��!�Y%��u�_m�!�;�׹��|J���ڦ�����l�ݥF�^� ����k��V�)�� X�K�y��� ��e�@�"F^�:s��NTٹmM3)���p�eC׏p�'�DK��z��f�X��	���?l�-cC��Y���e�����j�z��3r�IƲ�@��*.��*jn��C��8n3��j}w{��@#�V< �N�k��۷�Rv�7�41;h�}ݠH78�VL�v[�	XIX,s�*�k�م�I�̦F���B�:T{6h`�;n����]����������7�*QNS6B�j�G|벹f�8^Ρ�X2�:��Ɂ��Vj���F�)}1�U���Ǜ��wu�Ji[8W=/6IYw.�ub8W"r��gm���t�B��1��W�eƝhU�wz�L|��v��*�e�}e���̦�8��	5ram����ۚ���%E�\�H�:��#��`��^�[ �5�1;"Ewp@��1��N�4;)�$��f�ueN�D��=��ڴ���8a�|!U�[�A��|D�Qs���o��!���I�P}�J��У���:ޤS��h}�ȁ����y|�V�� �ޫ�\��w]|2�Ւ�@�>Wc�K/�͠�$p��,�� n�3�`���*��v�r�y[S�� ,�	[4�\5=ڏ��<_p��ŵak�L,V^iAөe���i��v0P��4Ѭ5E-�Å�y���T���-wN�j�[��8I�c��Z��ȴ�s/D]S���s�.b����wb�E*��Tqr��+�Apvҹr�١v�6Pn8�V�uq�	���ZiΧ�k�)a�N���YLP*�@3�X��q��I�@�j탆Xw%]m%�Mj�H��[3J�f`�i�u�n��St���{0��P����A�����Yg2�`#�t��ktO��K��6�-��]�3f�O��`����Б���q_h�q(�T��v)d��9S׭�)���C4�״t�o�B��X���z���t"�ZV	�Vw].�!�duه������E���'@N
)�v����Ӿ����eNH��K����\�[2���{4��m�C�r\Нع/����6�]`�YGI�6lh��� �A��j���/7%��a�L�iǽ��*h�O1>�r��1�v ֈ�w=�v�b���z��z^;�'���t*��n>SE�v�ú��׏HwD:�V̺�߲�H��.":�M�8��aQ�������������/�{����������[���7����y��,���v�'��:�x�{�^�<�Eܩ�i�d�E4��;ug��:1�����	��<�t:b�9C)e��@��0c��Z���2��KU��#���*��u���%Ե��˸e���B٥ HXWħ6��;�u[g�h困P�%��N��R՜9m����*�v���e�]j���4�V��6�B,Y���I�w��r����Y��EC��Qm�P��{�d9ǩ���n�+����Fk�4�׫�;4}�Zeek�H//yU��M�\�fGt*�T$�Q�;��cg�|�����+��N�a��V���N,�[�L�/�j�h��2ss�q� �Y���Y�<4�Y¡6Af�=C �
�o*>pu�miIv��4��9*T>wVo�~�oZq�1��k���`k��W6C87�I��>Q�*nR���]�K��-EG�5݈� yY/Y��P��T�)>O34�eJ�&�K��r����͂:�����fK1�֔e=�[�"�f���{
�J܅\b�#\K)��2Q��1��֮�c��wS)�zf[J�uIp����YG�#%��6�+��37t�o�;���.�)4���3�RW���lTmԷ�]��3�;�5ut�n[��ٻȒ\�}��{�`�pV�C}r*}/2��m�ϻ�'D�A�˙�������Y[}ٛ�� ~�E:iR%���Zh:a:�������
G���n�<�^�TL��XhQN��[�M4�4EARf�E�-�RN�E��H�P0I�i~B�
e�I���m���k����~�(�!�F9$7=�VG+��Jw�����T^��{�ۧ�=O�8�Yӟ\����]��}ʚ��3�];�pԋ:�����련��XI{�z�'k���	���������?^���G���z����nD8��}g�9�+Ͻ.�)�QӤ}�*!���%f먺�^���:h�EN���r�-Y��8�Qr�'7I�|�Yv�]��wwO�����	y"n�)�JHnK�d��]�JJ����[�NjJ׎�h��|���J�8�D�L]�ܝ]P�� �&!�,#Yb.���%Q����r���YF���>g���y��{���P����ssh�fQ���Z��75�!)i�\B�U�\�(�n�k�x}��奉�	%P�IʌĥD$Dīd�%V�J�G�^I���=�8E;����w��L�/Q�H-s!�]���";�^t:&��Gu�V�L�wM>�S�Q&�{�=�V[.c�WC1R32O�k'����b�ؾ�L��m�Bŝ�a�"čE6�d�goXRdwE\���˯�o=�|t"��y��bO��T�9���` ���S��B�&J$D�A����< w�n��yt��>�V�y����u�iN��6ؾ�C;*�K,k���v�/7�~um9��ٗ�#8�P� �����c�7Xq��0�o������[������TH�Pέ?eG���ݯ��s��Id��[�y�+y����,N�ջ�.�	k��`	�n���t�0w\s<d�w��ԓ�gV���U[�EN$3.���Y�3҅V��z�]��%�d��W�/S}����W����'�C�ӌ���>��d˙˯9hu���k�����'��v��O���y�l�~���]�1�i(��{s�޽�YދՓ�����y�k�ONֶ���;�WΗ=錭j�{)!�Jw��h��ȴN�Ӌ9/N��C�Cƪy�.��z��.��{(GAm�/6nx��;�m�A�����f$5]=TϽW����^�]�\�����.�'���6FZv"�)@4#�~T�i_/�Ԇ�f��+W����  ��Ah
`J�TV�f�����	W6Ӏhf��}�=��M]��p�W�����R�w٢�0]��a�����+L��fЕ����&��	�!Gw�Aor�1r�	��qG[͟OW_�S��*�n^U�AO�K}ms�o�d�1���}�S}�Xoޜ<q�>�F�9t��젺
�E�W{ؘH+���H���|�NW2k��6�,�=sF[�4v����<��7�hMN>�;��B�r<O�/xiQ���=�3��;<{��u;��cʫle�%��+������^t�'v�����:Nz]GʤM���`���=�yx��߱��O,^�y�3�'�Mǵ��_�h�sOm��Οo�S��w�ƢJ��~����s�J���� �Q���J����R'ٻ~�=^p�G7KN���
��r��+���"[�5a�V����|���G�+7��33Q~�uxݛW���
�ӻ��zmq��/�'�������5>f��>�-�;Yzm�q��5�&�X�z�I:�y��y�}>�<T�1f�cǔ�cP���S�Ht(�7��XZ�ShaLl�u"UAa*��t��-���6r��эl�od�.��Hx�*�z����x����jX��k"��u0�y�7rd�S)�4E�^i��Wp`@z�,�m���&��ΛH���h*s��)�:�W�N���pl�*E$�w�_��C�|� n�Ïc'2�$���͠ ������4Q1t�{ֈ>����	��Jy��X��s�Nz{~�?-����������N�OT{�{�b���S�t�U9�o���Γ��{'�6��XV��%+R�4�{���K�ժ5W�~s��~�D�x��޼V��_!y�y���$[�/k܆��,�J�'è}j����A޿(�����w ���u�����%��s�$1�M3��,f�e�3T���ׅ�������=�sϚ����\|�C[5l̵���/��o3ض�z{OU�x�Rp���h7:�Ԙ��ެ��ܯ��\�%;�)_�y
���O]��|�nH��߸o�Q��Iu�㞉[���6�z����mg�X�_[S��9c��Og_չ�b�s��,�J�ELjfה޸#�k�@10ȵ[�uz�D��\����N:S^w�3Iu�-ĭ�4[�,�N��:�p;eP�jqo~%�]a�a��jgl�8U��ĲVh�%�m`�ۍ��*nL/&Z���t=FQ�f������[���H]��d�9t�O9S�7�;��%C���՝���@/����	Ȳ;���f�˯�{��n]��	�9^�����ثˬe3~u�P�w�ҳ�8�	�Ƚ�lYG��O3ݲ{�{��罓g�����po���X�^C��縷9��0tQYf:���97���Y;��v�X��z���
bnl׃��g*��]�����t���$�;�9�c�;�3<Sqz���yt�W�-{����5��)�׏���=����C;�ݖ�x�t��Ey��r�x����]���kG��{yŪ?F:��N<����սϧ��D���Ǹ����Ȗ��c0�����Gv=V1᧼��[Ч���8��=��rov��#������8{§͞��s7�:�<On�7��N"����go�vs!���n�5�����]���˙6�Z+���F�Zag�G+�����{�ڒ�
�2�y6����휉s��g2��E��a��b5'%�)�{�>����M�w���L��	t=�6�E����������x�o�B�<�M�c�l�H��`�G�2^�ɴ�u�!�V}�"����Q�t��
ZΙ>g��7ʣ6jjh�~8�^�r�<���Q���g�J]#r�]�^Y�z�.�[�c�F��� �.�jy'��3e�}�՟R~��.���F@�����6==���g�(�׽x��ڗX_��3���Z7�Uϳ�+�u~�z�y���9|gy�tFb8O:�Fz����4�{�]�W{՛�.}��_��/b'�Dax�>W�M�>�k�~�%{�{MV#�ON��O|A~��	7Y�Q���>�Vo�������d�/}���^��ob�yj:����Q�;f���������1�F4A���{Fw7���;x�4��xH�u^o��$��嶳�^b�����˃m��מ����E^�S�y|a�9����҆��/�����P���͹'?}o<h���&�Eͮ���uL3�%�,?�3���WY�!�5�]bo!�=��=�t}N(pmmh^��yP4U�]q�/uE��)WK%�)l.��̤*+὇x���Y�0�H��ts�FS$�-�."�`u'R�Sˑk��[�E6��j�wcd�Q�ҩ���\F��i�r�O���/I���y���h�S�O|jV[(Չ{>�Cx��{�O��,՝I�g��c�0����'�}�h�������&m���$����ksV��mzˇJ���V_uv���wNXs�:2��l��w��8�Ծ�z�`_y٫�����Q��o��W�:rz�}!�@�}�:do!J��S��:��9���ʵ�k)�?G�q@���L�'���_��m�U��}fs�C���R�����{��~����yy�~��][�UM��K��Z|O`c&ۤ4v���y�}�@��N#�!�`�~�9�Lj[Z�4��.rr�����o�疛�z�z.���2md�zu����^�4�Z�s�F��k�n��X�S>^۶�A�����AX�Խޛ��P�V�����mii{���T��R�>�3�v�6k���zkr0(�g{�c��	���ގ\�9M�c�f�Dv�M4�B�
��y9�p}�I��tk�Rȉmr?-�������*�,���Xe޶r]�8Cwx��멃��{��Ռt}�_pum1>�d��'.Gɂ}�+ʋlcA���c���/J��K\�;�٭��_U���+�_�{����To�~i�<������ݎpm���!Ѻg��^�<�w��OooI�|`��2z���$��zKʘ<�����3�ǽ���T���z-��T;��硪����>nR��[�O�=-�$�L^�6����Q�y��aV|�MF�p���ۼ{|�x�c'0����'����xޒs�{�Q��Ƭtvݸ�Nc�Z�y�^� q���˃2x�=uݼPuܗOo���Ք�\~������q����k�]�h��/u����7^bτ�x�<��D���ڨߞ�<�ݘ���3��_�?����,�ȹ���zr}^���ה�O(u�9f���b<3��8y��.W��z7��;VNs��&��k{v��Z��O�z݅�ֱ��E	P�ÜVΨ��+�Q)7ĠК}�=^o��z���}���56y7�YD�I�u���%N+b�g��ְ�ہuv���Qe��ʉ�9���-敆�Q�gd��;	���E���N�[��]�7rnu�ւ̫����F�s��tg7���䙗@���#]�)����٩7)|�*+��Fm:C|i�no��+}�������r����M,��S�:\��3�˧yֳ�^� �o���Pr��a�~-�nT�Y��ozqH笡���t�ڞ�T��퀫�ǝmg��_[�=�IǓ�ާ\
#��^.ƨK��/�R��?g^�CcY��r�{�sf�K H���zրb�7t�^�`r���Q����{NI�g���|$�X��w켕���f�n9�2+� ��5�7�N����n���y�;�h��N��g��=<�t���r�y��Gz��wSt�	o�V���3�ý�E{{��ǔ��䁮M0��\��g��N�rHm٨্]w�����w�m�s�Y����CМTg�����qcHw����kV��2�u�v�D���/�ٸ�e�F��N�Ƴ^��1ǈAis{���0�}bv]�J]��&愩�mo �!���ԛ�JĮ��u�[5��r:��Hky�UAV�ك#AT��~��jU�r�nV�B��JHۥ���:(�^���K�-����?+��>;{��^qՎf�y���1>�gVS&��d�:�;e��#�|���Ow�ȼ���}U�*T7;�	����3G�|��Ss��Nz��m9�{��ɏ�7��(�[mO�^�c�:W��Bo���_
���1?j����'���������	AoV.�u��f��ZyI��������V��B��Z}3�j	U�d[a���)���>I�5�7�g�?Z5pӥ2�!W�3C��Z�/6߻z]8����~�a��M�[Md<��b<	�>n��F�gH|v�x�p��0|�1b�*�����M��sè�#H��=Lga���C_�vƩi�Yٽ�����X����˱��B�?���׽K)��^�C{��?t~�A�<Bjް�6����+���W�x�ם厧z�_�2��z��'8������6��>Z���X��!��HHq
{N`p��حYW}|�\��W*($"�_L�#kMm�J�J	�;�e�C���VA��ˍ�r+�W���މ�md&�$;��\�6\:����Ϭ�����U89�5�լMp0�onJh^��;"+A�q���N�o�ޱ0�4��6�Hs-R7�@}y�k�4g��Cݠ*��P{`^r�u����������w�u:�'~΄��W��N��R�t�ǧ�*>)E�̼����y"�Ǎ~�b+���t��g{����<�>�_�'_��jC��f��=��C�e�Ǽ2ݑz1��'�ϴ��h��|�[�,���W�s`1y���/?h�ϫ���\Fuz��z��`�M����ZUr���o���!S����8?���o�Ve����ٺꮘ�}ok/�{�=c#,�W� ���`�g���@���ȿ�u|����y�yU��}t���S��b��Y����/+�fw����y�z�����^����Fܺ^�����<g����eGhժ�w!�����7g���s�2e\�(�Y�AJ�?�������][�|	4Zƶjy���t#,*�c^k2���p���h�n����U�xrvK����6bV����7:�Y�p<qV
'��6	�!=�^����:��±fj�d]G��W]ql���Ds1�]ٺb�Y*�`���]'w��7RR�.���Us�tcP$���[����]�̺�����ׅ�����U�9/�c�gh��blU�Ž��Wj�ss��G��}*ظ�-o⯔�vk���Fei�6�t�Z+�<�z�M��t�_Y���C�l(�/���� ��GFP�ى�J�l�LʐZ9�54������M�eo�Uվ��hX*� ��C\���' Y[wХ��J�	���h�J05Pl�U����Z|[�=җQd䒛�W˗7���KKB�ٹ;4Y�d푞���&+,������m7����і���}n����0<0��l����#IV�V��g,O"����յc��r��[��Xf ]=z՗���[3�4�D�n:ս�����g=ޑ#�Q����*�}��n�8䪱}2�з�0Ks3%cjأ'9�1ݡsDU0I�x�
ɸjbT�JҭԄ���O����Y�/�7-v�N! ���=�� �qnG�(Ñ@V���c���E�ʥ�]�r��j�S�+���@º��>E]����t�j���\Ku-�J�`�+WnI�W]2�q�{��4ս[Z!A��=d�7��M�I|@�� ���[8�:�o�\����R���r��r\�Uo�,B����;��ؿUw�c̆E}G|i�^u	�w5���OjqC�Ƭ��^�5?����}���#/-t����d�EE/��R�N�B���QU��tκ��9Kf��m��S"��-����E	�:�
�c�!��u��n��L���*�=hI�3��u�n�Pg�v36�i��}�r0�F����i����T�Z��[۶��R&5ڐ��R�����e�+k�W�*I�t��9�ٵw$~��FoIVʻ����J�&8���R�q�Y8��`U�
��]�](��w��Ѵ3nPm���QӶ�>�r��;�kl�V��ކ�%n�������q��EqǢc���	ŕʬ=#
�pM��c�,��mg�����1-�"��r�m2Vo�}3&���n��A�V�=S-�uu����T^��9om5.��ul�w�ޫ陂�V�����5�}�3v�-��s�"�͙ ��jWL+���6�s�a��Ԃ�o���y�V%�[��ʚ��wg)�7�c��X��8x��oz��bIVܧ�g�Z�ƆcM<V쳕�ܨ	k�N -��4�2�e�1��A˗+F���XF������Iwog���`fҕ�v�u`�5;}�-
�[�:˲s4��R��v�{\�\N���a�59a�M��3Or��y���6���K�]\�X��ov|26=��rV?x��%I��Dj%_�k��K1:��?[�����J��	�#����y�-1��|ߝ�|�w�P��L$P-J���p����_i���N*y�".����!u�;I']�bDY*Y�뢒�Fd=�����kO�;"�W�f������B�= ��>y9!���⧞�Nxr��4����ÜKNF�4Ϯ:N�w���I�E�u�J蕺��/,ͪ�u�f��<���+�v�U��:"_G<������uİ��[��}���E=��k4ދ��n��2!]�u�W��ja� l��\�I*\���T���[��Ey��DL$�D��<���<��0�%Q>�^OQ��'&=��n�ݺ���C$�*��/"E�RZ,������(F��멪�;���r�'^e�\�z㙦4�=�ӧ��{��9��{*𓓸�i
���{�H�b��KP�<똘�s"*L%,������"u�ڥ�v����u|I��Qד�i�\_	��t��a��c��J��ܱ4L�D�t�y�l:V�)��y�)Z}�����%��&�*n��K��+��z��ͭ��kL�CB�(}}�l2�ɣP�;�����W���<z�|B�,����o������|N�����]&bU*Um�������;�����Oٳ�]����BP��};������I��ǁm�q0ISiù�t�m�@��y�2���y[R�҃s�P�A�M��g�b��7w3ٛԌP�,���?$A���R��K�ی�7�X[�+�̥z\F:�)�E�'���vXțaؔO��!���+������o�{�ǂ�]~��<��3n@DH���R�+�Ԣ�]FM0Yu ��YW@��d0������(ȿg��κ���`�^{4Y��[h���~] k�5�eю��>cs�ԑ�@af�۳���+=y��.u�2���4<z&)9��QI��M��1��|`76����b��t	��;��R_ӹ(�\h0=�:A�����ZQi��j�}jm���99�nջ֢��ke�����oE/3Ű��}0a����2���;�ߠ��|Ⓤk2�t;���vr�G
���c���Y�o{P��YBP=m�C��*��3��dg�J9z�Lf��M���ƴNϽ��鳄�ϑ���t$�b�l��١�0h�E�C}�\�H�ܑ�mW^i-�nK�7�g�n��;��88)�Z/�OJy�4�w0t;�#�iɲ�J��Ċ�o\����X	���d��C�؞f�2���q��;C���:��&�����)=_<ޑ�S^�{s���~�P����� Jy#�J��R���5K���Π��F�n_��s�*~ B��|1W9<f9� OO1�x��.�Y� `��0�њ��*qqa��/��+�ʭ����&��"�L�r5����_D��z�Y�˨�<N ���S�奅p��=�v�S���+۱eߔ��E8�ܳ�B�*���Qa�5ȃ�C9�Y�1�6n��
�z���S��n�5+�zӵ���Ctw��lr��z���3eƸ�3l�OC�z˻��_jۯ^O�+�
�y|�U�t$�VK61�۵����}�r]����N��>�y���d�/{ӄ⒵_ڥ,t	�?}"�.0��Z���}�w��#v:"������-�2��o��3�$��z,���E>�I���L)����{�"���
Yq��7�
���n�/&��5��f���`� ����"OP�6���|�څk�� ��9��｛QN��2FT��m՜���Tu��yud{3����[��+�7�z�ȓv��b�Ң�ZaRk)]E�M�oN��zƓ�]��i�h�c�
y��I�ߞ	�
�+�����i��=mѕ��'^b욁�c������j����G�JE��\j���`�����P2�rk/n6`"f����=/c.]N7|tgj�We������m�H9�ﵞrX�O3�F���������5��t��ml.� ^��|ч(^�J�_����MJ��U�sՍݓڡ��v8������BSe%��u���OW���S��K�C�ӷr�qNdOh|���#���Žt�bX~� ��"y��"U���p=�N����.��E7Ҙ��l��n�}^eǟ��*�,��ȋդ�E��/U	\��^��W��1c&�hh<&���o�upO7)�A��y���K/uF�߹˴-)+�s�r� , l�=������Y���ޙ}qXU0MZ�p��"����
��#ßO��ӤM�>+E<J��:�����؅M��ی��	bb53Bf]/��vq�vJ�.6����~��)���.V���p#V�~=זl��Q]�]l�R��>N	�:׀��㢢���r�x���p	I����S���5˼O>t��+���1ȃ̠O�ioHC!�� ��g�m:�]7�v�4&9t��c��=Y��0����t�\�����'k�NrD⠟H��ȾPKXE��_o;]�w31�"���II��66|{]�5wD-J��GKs ����#��eB��ǫM���3%"�3z���0�W6��r:o�|ʱ���sY?_�F�c�nz��QD��M��6r�a�}��C�e�����w�i���m����0	���*�+�22'hQo������XK�IΣ��@�g��u#K?�[�d��I��J��@� �N�f��ۆ��q!\d�a����u%Ю����r�wC��{� ek,s� ������҃c�����<f `���w�m9�����xME��ݍn�wuSCP���@s�W�ĉ��V��H}�D�7̉��^�r3�wBhݵ} �kƀ��o@e@�3M��Ү�[9MJAeI]
���2��sl�ٙ�Xkz5<�:�����;�
uRVg�|g��|hBEy8+Ed׋PޕX�<J�Nb���Wz�O\�m�r�i������|'̧��j�ƪڟ���P��7_����v������7��+o1�:��l���\��)�Z��	=�G�z�\S�4{M˛�0z�dn5p���������_�c{6��i�^Ø�兕R�� J���Si�5	��¬-�%����e����dn�Ffwv4'b�pF����k�C���j{�<ׂqMiz��r�iΠr*�Ɲ���.���UF��t�SG�""56�&_�"YO�CzGa1B+Ī��A`Y��ùTO��vT��n��Ȟ���s]��J�=�-w�90ILW���&�j���� ,�f7�]F݊uo��4�޲ ���@��$�T�ؕfL���{oWV�9�"v�rG�_�|�����Y;�9���
KS	���hW)j���K;�e.r���'=��U=�
�ZJ>;�������$DC9�2ro1�����v�C�9��QW���M��^`[�t�݆!�3|=(�lsYU��r�_�x�̾?�h��z���]�<�5��s+gl�gU�?�D�6��c�g�Gp�Gyt���@�u?*��>PN���ήk��j�{w�=/:}��ƭ�4y�A�u3��w�LW��d��&��&��|u�y�S�V7sx��$(��2�����h<�#sو�J��(t��UʁDe�����nJ�A��Q��1q88���Pi�hi��MB\g��͔{6�7�m>/�(i0ISi§�S�.��U�tӫ��=�^kI��%`��O��������LpU2g�'�7���X9�g�Yax��ğe����Svv�v�jf�V��K���vE"��ʵmzj>�Pۚ�7����3�jT�Ɗ*����D�o���x�U�s���ܛ"^G�D����*�v�.r#��]A�s�~9�p!�> =��8s������V��&�2j���M�YT�emk]�t�4���'�����0�4��ۻd<���赈·i՟h�0x�v5�}�z��a/r��Q���ǆ?Au�� t.�[�=w~��
z`���7@�hMo`�N��0f�DLnaV���&tͼ���m�,v�ޒ���7�7˘�X�Ew�Ó.�=k����&�\���LO1Ö /h�������K�t����_��"�W�������W��:��P����7��z�����Ix��r�0=�t�����ʠ�%���B���W�9���Tl\Ḹ[R9R�1O�k�i	��a�}���dH�&>���j4��ڂ��s��'QI�f��/����NI��	�'桅�ܐP��7@������sԮL�A{��J3���2`w�\����ݫ���U�C{6�o��5������05$d���
�Z5�B�N��ٝ�N3�����^��t�.SJ{H��:$}b%+��i#�"0N5 Z����1a�#KOT.�0f�d9.�\Yz��d�0�g����>���f�]g!��먍<��#���74�F=fmyԭ��"�ᡂ�1�<��4:�t�C-��g���B]V���U�Y"!,嗼��I$�ċ�vΚ������{��\�ݑ�^;��a�ơ	n��� ��ފ�9�u|N��U�I�A��Q�՜U�D�ݿ�ݽ8��|��t��^F=�ІM�@C�&n��ȝ&
�"M7Qӗ}�u�:���W�bJ�B��7#��in�)��V�S-l��+�A�H���⎥�4���d�;AEk��v�
�"�䭾�ǲJ&Xɪj��םA����G礼��G:L�b�u�rz�y��v{{md dLF��q��'��K P]SU��)c(F/|��D8�=�L[r{�=]Yu�r[6\�`Ȗ'���E�/vsJ�6�X�&~��EK��L�[B>X⾅8��}#�q�E��Y�3'1I�~5)�w$r�5P�,�a��B�5ȓx��'�IAݨG�=B#�<w����	��c�OW<n���ہ��n�*H�]��.ӊ���
����4-��/=��7^v��0����4J�zنnJ�!���%*���O�u8w�1,��&"��)?^,�z�<���QS:��]n-%��/!۸=���m�ՆO2�}j�=��'���:K��g*���6c�	۶���>��%b��_fP��;Y
��J�7p=�Z�+�{W#�����̊�Pu� �;�t��ֿ���e��R^,�܏�E>��z"�i�*�DY�L�Px�sK
~��r-���vp;�׍c�y��e����=�EJ.���ʹ9˵�p��o�V�DY�"袡�75gA��p[1ױ�}�F(]�2a��S�d�����ih�V|7�����*�$���rC3߮�P���9��4�o :�Ⴧ�e?U�f����:�B�'gS�")���G�X�G\ԟ=����ۭЖ<��+Nܻ�%��9�Sfq���X�׫�5���Ί=�Ǫ�=�`wV�����[5�E���"��N��Ts{�}�_����ه��1$�S<zէ ����}�7��
Y6�9����_%:^�0pvζ,U�q�7;'j�#�B��`��<<Θ3C��zf59��e=��[�	�C-)���@�'��g!�2��U6���<��	��vǊj�a�FH��z�r ,>���Ş�S�4���.l�L�]�����r�p�Ƶ�k�5�MIjhJ=_ls��8�>�97ʾ�Z�31�����f�X;�3]a����P/���L��f�]RRu�4bP���"c�dʛn#�Q���c=�jP��M��G���V7c�\��9Zċ�>}>)���>��sG��]��%���,��3���D:��5n/۱�}`wT���AcEA��H��j��Dƞ͒�.T݈�Gygn��Cڦ��HＣ�1�7%�uռ0-/^�c\USc^$�U�	�НƦW ҇Uo�2����f��K�>�B���͕\Y85P@�=�@��\���uq?q��eՔ�n]�SP��Ws�v��uǴ�c��5��Ve���<?����)I�9���Ӑl�o�gr���U?a��/�*𴉐��6��|���gV$��<ʈǆ���(<�j���b�Xy�/kc���Z��Y���cR<�I}+/$�[;�*ٮ��ݨ{FXUpU�Y��ۍ��b>���ҝ�E%aG��׹,��mM��d�T�5e�=N�w��������� ��0��2�Iaɥ׼�}
%0��S-�%Tȹ�jU�o2q����y�(%fw�g�v۝��1ޙ��zwڃ��^̍8zCȎ4���%:a~®��SM�J{o�S�����m��+Pnl�En�g�v��?F(Fږ���m�"��S�<��sV*
���kNO9�Xm��L����o�q�E5����Zt]>CO^&<��������֛%Qǰ�	~Y��gK�[��:7DSܽ���Ɏq�Q�I�F!��;���L��¦NH�u���v7Rw��VKٙ�!�6�>����E�J�����B��(lse@�an�R\o(1��QGA���OL��$�>�cgv�^wm6���s�3�3g�z�D;� a�� �>X�a򠝘�k�%��R�Vg{�9����1�} �Rf�#���ƴ".��sk"�L?D��,��Wy��&�![�(�ge���dwr�G!����*o�`�s�.�<�j��8�]�;�h�O�q���5.0��c�a�^v��5�?_��-��H����j+U��D5��Q�wov3uO�dX,ߠ�R�;�9m�����.ߤn�hvZ1mi�"ӥ6�������Z�Y[ׂƍ�H�BM8�1aRz�*K��n��҄�M����u[�36��;�����J�(V��~?��A�p�s�6\"���=�<8�ۙn�eCg.��+�Ǡ1JXd�܂����T�Y��]}�o&a�m�v����|����'�q�y$�g��
@��&�j��ҁ8��&���5�nMcV��F�:��gg�N����/#�[�+��mz*������8�Dxj��ʡ]��s�ꋑE�G<��Gn&�ӧ*����΁7#jM{�<i�<^7uG=�+��%|�{�^�2��\������ջLS��N�C kU_m��b����ͧZ��n}���u�)Z���I��8 �M��������j����#~X���O�=s�r�[�l;����\ڠ�+��ٱ���X.wd�=��]y�1���?H���yi63׾��m�\|A�E����&鮣�-��֠�V��s����r7F��3Y��hw��UJ�t��Ͼ�j�n��ᦌt��{���tvWr�~�}�/�Í�v�I@+�)䎩Q��J�������`�GI�yN<l/'��"��'��ߍBhO^	t�:���A����%$rFA ���~a#�>X�Y�^��G�w�t0���w�f$��3�	��K�Yj��G�0|D�6�����m��.���-��W3/.$�{]\(���ɔ�S-��� �]f����=�Y�T�w�%k7Je�wN� }�O\�&%Y�*�e/ A�`��\���Ķh�Em�mbܨE?�=۽�	a�xfKy�3+�:��B��B�o����n��`�rP���ĉ�K!���iD�O�s�{N�C?gd��i�o��V��˝��R�</6D��[�-��ג���=�Q���h
E�:���{�8@�%R��Dҫ�%����]��1��V�]-;2�bV�[vk2=o��u��)��ʋ�bԞDZ�w���Fc���U��k݋��v��K�d�m�l�Omsz��#�7��&ABoj�J�v&� n�!��t��3,��PY�a+(��"r�V4�dZ�r�ܢH�[�U���*	��A�,&�����S)��[����][մ�q�hs^T#2w��Smwxc�)��88o6��J��F䛗��7��������� �mZ���|�P'���!�h�L�N���U��<����mFs��,���;;1��6�L#�ǄBǳzi��P
��-�3��Q9���f	#"�Cu%;�K�YL�MS kA�� i]j��39��N-�]� (b�/2�,�:��쾛�g؊��G���ً1��g�\'z,٨�������-bS�Շ`#��ֳ��ǲ5�IV�7kel��� �t�z�ջ��|��{��*��n�9�2�+��NYyQp�F��f�ܽY&\�mE+Y����1����e�F�x�"#xW��K�htc��(��ͬ��CI82Ň\�r�#V�v�wa_o1d�]u'cq��;�(K��,%S��}��t���N t�e������x�;�ȕ��(T��"SS���K���Omv��F�Snۛ�����v!���:aT�r�ۯx�7v�''z��ao����8Ńw��GcĽ}����tVU�;�]l��NQ�����i
S��Os:�������C���:vm�U�[a�������Su��Qu��i��g�LB�{ZB����]I��Ia�����d�ٸr���:��<���+��WVh�Z��o<*xB��9�b�Kg�>���tT�{����R��6����{@Ƞ�4�G�j%�Z�ms��{�kd���hd�V�4lm���/���ۏ%��2��0+�=�"s:�5Tt@�s���lZ9�Yec��Yg��'�pJ��ۺ"�bcQ��2�]M�}4d���]�a�;�'��;�a�&A��thK�Vw��i��	F���L�<�vT;�#�x���z�ԣ����kxd8���{�'}hݶN�6q\� ;�B�&�M�H	��{�nI;7gH+++���O�l�,�D�����YqC�wXl�%x朵ZkW%�ܾ�S�b�N��h�S����$O�����wϩ2O؞�Q�"�R�$��$JD��֖���/J��Bw�.F�^���C;���]��~7��}�u.��S�au#�q1J҉%�9Y���&�۷9eӢY΅i�H��|��w2�������t�Y���<�G��<�3Si��}8��t��)ej���g��e*W��<�����l����C7���F��1-=I��^a�ds��?;�x�EBO�s����=�W!;�9YI�JI#39{�n�J�����I��;��n:NV��{�M
I�*�x�S��y����.Nwƭ_8��p�ԡ�z`��o����>=�eB���{�T�1۹�F��.��^)��_�+����q�-MM�<�� ����^{�3�F���!x����#��y�)D�{ܤ�7�q�^K��ϟ9<�����̢)�����	Y��tw�I#�O�������rYE�rN�C�븺�.�w�9�G�~R>�Kڄr)��7d�E�|�ۓ�x�A�)��'�#)J{��|�ʼ]єK�Æ���ݐ�r����:��]hs����J��m"�wpv;�r)�����nO����&��*�M��~q�!����v2��U��ұ:�EW��d��g)	gS�k`�%���X���]�3��YΖ��pp�QH�J��P�U�ǽ�>��߿o�!�a�Se3�ap(���l.� {�3x �<<����xh0�Z»�aP!�;tj_�|��
z�:xл�L5lsBr͟E�ͣ63�x;k���d�Q�9���H�tb�d��|�K�T����I��<hu��u8��F�1�-4#��UW:��\D÷x��{5}��U�T��p�� ��1���0��.>���c��۠݅�m�X�������}y�4�]�#�Eb�B��j�ZȌ�j�	�t.I��72��"��}��o�Q���웭����Or�o���%5z�,�
�c�D��".-�;ܖ͊���dYg2��/b�j�̍ai�k �"ɞ~�T��$����:��dZ�2����3v틳�ԾK�qm}p
�SP���A��.R� ��x�^{>JJV��شy�x�^�1�
#�Nwkr��ƤUD*P2\�૩�uJ׿a�CнSe�<�D�r�aM�+��QM��<�1s�2R�{ɺ�z��r[���R�q�)��'t�h�t3ڽ�QI�F��N�T�2���4�v�Nͤ&�J�\]�چy˃�{Lz�m�w�S8�-Q07ΰ��ٞ�4ϏX��*��|�{��
�T�J]p;+s����I�sz��yK
߽*��^�Ѝ�ac��II���6�(�v���&+��M�Ⱥᵫ��l<���M��\o3;�w�M�U�'�ʚ�Q�ңq_]�]3��'WCgde��hi�$�?h�v��s�#�s���.l�pl�l�av�0�fھ�P�Z����"o�׵w#1�VB�X��*�D�9V�W��$p$G�`��3h͐DĮ�����'o.rS`�V�)�?`J}�H印js"(s�e�QQe��{s�������;��9���8��R���F��<� ⥗�6q�8v���$mN�����{�.�ޮ����N���v��K�H�?�B�a��(�\��FK%�g�O�C[>��*��N�CO2�k��HI1�q��&#]4A��EG�;8ػ%R���>�Q��� ��� ����zÃL���p�P�Z��D�
+OĖ�W��a��z�V��{A�%`蝇ut���a�q���soW᪶��u=T��L[9z�v�*�w�!����[Q%�Ϥ������|!�;ɳ��R�@��qg�Z��ʸ,:�o�s�G��:#|n�|Ѕ��t�����a�4�vM
�݆=��&w,�>2��z���g��x��01�@J��'cbJ���`��l�H��n]o^�0u���J/��72=�)ܽ�Pn�jF��5��t��)ܱ�Y����y/�9g�~˥t+��Y��I�Қ�+m�����x�e�΋Ժ�H�����fM�:�h��np8Ρ@U�+=��0f��BE`]#[��mZ+Trn�"n�8�V�Q�*f�!ˇ}��g�v��Ҩnf�rl��ػ��՜�ۻ�{�|�o0� �LM�E��M�Lapl��� � Gm����6�����[���q�b���l5�#m��5댜X:n�0L����ߏ�oz�/��ֿΠS6����͇�� ��H����Pl2/L��ˎj��.�ǹT����� ڼ1%��YjŻ�"�	n#:�V=�p����`��X����E.�sʼ�p���54��X�ʍ��~���*9�q,r��7y�_�ݱw�����;�v7j�T]���+��9��ޫ���f\�+�(C�H��v�`]��USs���hy�Y8��Ws�\hE��=�<�H���ۈ�Ⱦ6��d�����%9a`���bub�n��u��M�C��Z�}yv�-�O�݇F�12>�r��#����|�)��|��s�p9�->cN�	�D��%��?X��>ե��EM�H���AE�25[?z%�b�o`	�@�\���`��]��Unv��Vk'�بgG���RV@ϋ�:�Ƒb͐"^[�>&|�I}!�ґ�-gw�aͤY#A��Q��"���=(�}�	͐�`0���#yI�L����sEw]=�mdh�t/�W$5,_��:�u�֟I̲
��#Z@ ԤuZ9F��|�I ��W�.�Ҩ`��k)6��W���J9F�֫7.���)�I�w�rL��,,X���e��r.�Ԓ�9I��&�)��ⷣ&�C���a���o0Ü�aaɶˌ� f��X���rS'����fi��Qn��KE�Y^�y��P$d�0����'zE��ธȋ�U�ưc��q�Ģ�5@Z�[�l�+����]�+����`���#��_���)�=��Ԕ�^=�����C"~��
�|�Z6���m�]"��aÝi>�a8��$��}�%�� ^ػ�����QtB/J&�&`�z8�/�Wٙ���2B67z���t�����6r6V6�PIM�t�P�)a%�W�A�%�5SQg��\��fUCh���ʍ�;�(��\j+��;B]<wW҈�߰k�A=�V�U%���8��V�.�o�����3֖Jq/^d��Y�h���������2x��3'��4o���<�4�^䏼�s��O�
m��]e���n۶��Bqz�y�e]��q�a�5j%�m��� [:j�y6���ql��y�ۻ�jg|�O(j���f��6�t��x8�LSOV5-or(���{9<�:BxǨ�n��N�����/�|�b�񯥹G+���g�H~R���U��T`���bm)F;P̨��Y��)�R�3잳+D�&}���՗k���zj~��O��{nz�]L���nyE���*#(Y�Q��鲑��F1�V-��H� ǘ5s`r�ӗ�A���T�}C4ηq2�J�i��i��:��1[��1���Ҫ��Y�ϫ��]}�_���0.0��( .0` ����=����ԡJ�(��9�_%Z��{VK����Pg��鎂�P��&�(�ọ�
���2V�B��3Z�	�Y���n@���Gt����=�b-�*������,ϯu��{C.�(3`����=}̝��L��7$��'�r��c[�vLwp���O$t��zd/y
u!�ׇ<;9���n�*D���M�z9r�S�H�e���-�|�����Ð�.:��c1��:V0QP�Լ�)�S�<��4.�*�8���c�Y�� �sVlg��7g���Q8nrc/�lq�LDQ1�q�I0Y40�1���<hu�H���2)��Π��)kB]����J��@�������AMWڈ:`$M�+5"o���N�P�$_H��b��(ocմ��f*�ֱcl��\f�կf���j�a��&�\WP��qL(�b��#2=�����pM��{�%d{�R5���ջk����er�jT1ɟ��ߡ���j�JY��'^_��J�`�	���\��B�nn�;z2zR�~�uw^��o'�2mP�d��mǑN��w{?�@�IH~����+߿�b�}��oY�1P4���v����!�y�En���Ѝ�^���v�^їA_�w�Z�xv�:��¼ը�nZ���P�y{��]��89�ɹV$U3��c:�0^u�\P��̶���l����x}���y��xy�x{�����7��^ޮ��TQ�i�*�V������3}��p�L�^9��>�%&��粼3���'��'a>��"=pܤUxDZ�~��y����Jױ�eV����,�[��S޻�l�Fn&3�Fu��(���[urX�**_Gڥ*k����;혖l�&^�Ilnu˺�+.�mވ�-��b�r����n��յ$^C��{o_��N42A�'3ΰ�˵�@�</9�QK^��ѽԋ7D��S�M�b�z�-fP��l*�!FB�r%�
��x��}�~��y�G�k��j;)z�3!�d�c�l�=�n~���_�xuM��:}(��;}c�+��SK�KY�0of���K�:���V��|�)o��C���jÊ�_j�7���Ɣ�a�|�GO��l@^��ǽ�<�Ʌ�ѓ�|�;��9�<�������~�a�f�,s<«;�g�\��8<�f/׏�͕��4T|��CXw�LF-53�ʏ� ��C���)�ß���@X�������<���p�Z��x���ZA%�װ&cS�)��-�<m�a����T�l�`V�-߽�.�O1�VE�>�*�fe�l�<����xيS�2�l;�2+{c����$�*u�F�Ѳ�X�_Ċ���2y�d�W���� 1wo̆��-=Kr�ʒ:[ >��:��[.�f��r�7r�%Zj"{�v��`�]�1�����o0� 7������ y����0���yf�
۷fп�#*2?4V�5M���^�vvT��128kN���vS�����F+�^�8n�����&Ƞ;��*է%P���_.�(��Nr�!E����8�EV�V��A���v�8�ģk�㓗���ة ��9@�*��Y2�3@.�)=PV.��B��f�]�S+�e�����35"&zq�$M\�)�qQ�i�{<��a&k8s� ��L1�����~�}[Wy�t�M�+YQpZdz�Bj=�|w>�ʣظ�-��іe�5�Y��:7=x�mդmJ#�f�c({�cj���w���1�������aQ/��Ӕ�FU�1!SBdU�GO���U7�q�+�,� A=�@��6��C�U��N]!�N���y�S�X�,�)U�~⥓��4˯c{h��c�?~o��8�h	@m�CWj~�)�sf���aM������&�`s�a ���q*�E�Sm��YX�'��x�Iϝ���6WnG3�����B:��g�Y`߷��Z��<��!�g{Um�jN�m�#�8�{�ڪ��4	�p;��/�wu�$�岥�U� wĊ�*�ͮq��QcFt����N�du]W	����tDhpޓ�p>�w�GW���ItW|q�$V�S�B����fZ��S]�:oe��Z�e�ل�=�NeEo}����o7�=������u�����4���[Pw�V�8'D3�p��{���8C�Ny���:_�{���(�=r�a�{xw'x�cq�#P�����<xȈ���'`��zcm�|Eor�-�)F� ����>Fo{F�$�:�2S�go�x�T>��0@=C�J�"~�t�6�q�&��!8q�Mv�q���1�����F�y	�.�zQ���ʁ��]�C(����oAO�ڸ���ʽ�y���;������ֲ�i^޺�}3���(�v���K��ênL�r�ٺN��z�`(O���m!�L�N��e�L����@��3^�jYܵ��E[�ӡ�"�f=��o�3��A�8�&��BC��d���t6�t�����^	!���8�D�U3�\�����P(������J�̙wdJ�-}#�<���H���y���+[�✽�^�(�D������T��#	�P��3�����.���Ϗ����W�h�2y��y�ݛH�wO��Ig9٠��)��+u�"�O��Z�e<�{�!�_���b1��N	�Y��v�	��#�rB�������w��7Es^w/f�������|;�נV-���b�\ec�:"��Fq���:�7w\%��%��}Q̥�]$|{.}+R���Ǜ:Pp�Q���m�3#i�w�&*ws{�x{��0����� f��� M�`��F;"J�v��ü@qҽ������T�x�r��M�h߆<�C�J#�U%�U
�)��Ws�R#������S�*A=�^�PD�,~�MV��L�q-�n�r�ֵю��zN�'���Ϋ�Yc������"��F�b�H��l���wE4������h[tHUl��̺9���2'%K�}�r����6�rT�un�>��樅+�_��R�A^(�3j{R����������V���r�Ǫ�VG������-eO���9{0Q�d��]Q�i��ޤ/{�A��^OݡH<�H�g�s�v�2�0,ך#uK��r��q}:�����9;S+8��}��mC�����1+�c�]�Q���3�y#�Σ�̏L�?8�R/o^�8��/8��R'�Ga�MC�ɗ��)�:F+c�~�
�}�i#��H����~�n��՘l��Z�Q"�uP�:��R�Kz�p�L;�6���>��L�3nH�5��gkՕ�Ƿ\l��a.�d��'<T�W5ƥ���5;;�7�E�/[�xT���n,�	O]��u>vPֱY"+~>���:,X"v�dF�B$�%)��*��<�oq�kh�4	ĥ4yViy�d����w�-V����H^�0R�VL�߻^�*XMǔi��9�pKOt��S��pԋ�8�D:ľ������ }����o7��`<=��k=���u��E�%�q��5ă��}ef�d+sƤ'k�\}}#w]�1[���augV�E�Zޖ��#PO
���^�6\]]3�}>V��UB������8ۣ��>j�9ɗ�s�l�>]�ـ�2l�w��ݷD�(�K�	�6ߥ���j��w΍�ҎyU�����������r��
�>�wq0k2 P֙6�k��Ey��'[q�V�3֢
�xb�﷯Q��N\�U*�
9}r�ꔧ�
��5�����JwO�:�L��\�U�s���� j(Dz�7^��p2�:��UͰ�:�K�a�(�u���EI8�S6M��Z3\B�0�CLB����*l�־:�)�㚯]N�+��}�?P���ke__}��n���f��!��52���Ѧ�`#��҇>��{{�S?��F����Oս�&��#�MA��E�%>D�X���^��+!U�HQ�w!s�h���&=<�mz<\��,Q��[!� e��&��ה^�!2d��E1�)G�����s"6�~�������T��Q[ݒǀC����D^u��m�4�2p%�	�j���Vpћ�	�2�v�0*������+}�go_B��!`��ͷ�-J�w2�O�Θ]�b��qD�3.�rɊ>�����P
���;�J.�f���N,�]�n�m���r�[*�F��Q���9��&N�mvh|���)�r.3��kY[�rs��cP�N�h����u�ё]���*�hj5�V'��e�37����$��9M�yE���5r�D\t�+qr$('�8ۙ�F������[7&]������mMu�V�F�sC�f���1.��3n]����3��S����iy��+ j�+�u;�G�Q����r��{s��ruڻ�|��e��*��m1�c�Ϯ�]��wGW\u,�Q���)nv\�ɂn��݉��y@땐�f3�4r��!I�U}e�K�j3|�u�ș���yn� uZ�0jg��֔�>��6��fj@g#���wmE��Sf��AF[�8�,�����bX�Xgt�:ʻ�����Z��*����G�5K����fpH^,���}�1�ج�8.�7V��������35V7#�F�]� e�4�TYs��ϝ���CZA}�#y�@%u0:$�H2�u�r�wZYC5��Is:��F�m�J[�u��o"Ѱ���{�W*)jG�o5,�)�]�D��o�$VWV ��T��9.dS�Օ��Z��ݠ]g"ڽ�;���:�9]��ri�Rh���Qn�T��n�+D�z��^���: Z�Nw���gvT�x0�r�"��o]$�H��Ӂd˗Xn3)	,T2�p0!&��VM��Zٶ�nWg*Ҟ�p_j���u�,�+nȽM���Y����h�S4oؔx�������k:v3 �r��x��L���K��i�u7_�o'f;���йn�X���Ӭ갯.�c�	����l��ݛ�,,���N�op��}��������`+6�j��#lu^��yS����rﺑ��l](h<|h@� pή�7Gr�hlQ�o2��K;wb�s@��f���WR������)���h�w�e'�EH�.�]�}[��GJ�<p%i�du�l&C�@.��`L'�`ّ��$I�3Fm8w�C���i�p�<��=)uѬ�MXy�e8�-��f�R�m�2���q�wR㠅�,b�Eٖ�(��#��1�>�伝-�܉"f�'{	���V%��	��1��-uۥӷ��ɬ���8pDc��:`Ip�Mj�z-A�]�7[O]ѐ��<sX%»�=y�<�<X���ǉu�̗�R,�P��Rkx�^ڀ�nesY�w\x{����ێU�LF�'}/��/yyȟ�TgϘ�9ɕQ"�S�YWZ�5�&��������`0ef�Ŀ�N�Ӥ������� ?������A�`��U T��>wp�G��|̊"|a}IK.���3�"�7��o���(�9����9^uѹ�~ӗ�CE8���gr�<��ZО����������o�N���ع/�@�)Z���(�J]=w5�S��Z�H�C
���ⴿ`�A|�W\ �����ۜ)�;�e|R9qҷn�%I��9)d\�*�Rr�$%=���d���ʊ-N�����9ȹ�q2"�4Q��܊���sı� �"ʕz�U���VrE��W�/,$�Ng4��wJ���RԵ�an��B�tY{3;B�[IQ�/�{��ȈKA3"Me��|�TW�J�LR�����*
J���TSjaI]|{�wB�҈N^K�a���F�q�b=iu���3���xa���	�56��RM�������F�D$� �DB����z	��>v�jL�˒ |��hR��@����s�Q�t��� �#<ki�0�gQNuXZ;Mb�S��5a�b�����y����o{ޜ·}�@�7�-iᾰV56�����B���2=��^*Y{lN������-b��������qI0�*� �u���0�UjuH�jEP��F�Y�<���m:�=ɟ*+.6r|Ҩ5yv;f����h�;i ��IZ#��_�D��_۝�l]��K���ǡkE=읉ݷ�C2S�L�,%:\V�ft�"���`���`'��c�
�e7'C���ַ�vًZ���o$�z��F��G4]I�mb^��n3�(����>2�юo�Fil�k*4k���9�	|j}�4kԞ�ׄ.���@o�H�*��yM+=���ٞ�R�P�yaǯ�Xu!�V�(�w!�l7�f�T����@�Ĳ�	(��H/;d������=��<�Bk�9	w8׀��B�˅[��<��q6�/����y��چ���Sl�n����&5ң���)��]󵙊a��7v����~���NfJ�����^�:�u�V�S��DO�0��(�a�zgɂ�Ú;�uVĲ���W'�"���?m��d���@b{��[�������I5Z����s�suX��M�yGWbDD&ҋ�1<�j��(mT��SmTvŢK���v�Kn�f�e.О�L=v��e��	���(yZ'ƫ3��K�F�u~�������o7�=��a��`��q+��R��-��ǈ�1��3�H�T1�֨E ��B�ʒ���G�(���_�=_{-���cx��\�K I��t��T�~��i���Y�9��*�̥
|�'��WkjF�?R�3�Mp1�A���L��[�]r44�l��GD��&Y�*�E�j�n�YX�'��M6�v�����j�����4��z��`q�T3#��퐖�2)��R�"�Գ�a��͏@=>[��U{�u��﬜�G�����z�����-��mj������2an�>G��S�k7�����Ǜ�[��n���It�7�R���Πr(�^	G�1��qn\I����֫:CI�uq0��f֚�<� I���Gr}ač�X��j�Z���|^���t�
��_���g�*:>6��3:�=j^')5���RԲ���A�-"�����9����ݐ�����]�G��y8��KXj�(鯣:h׷]sGz����RMV�"����P���ܲ��׍W-NHR\>���,�^Ǥ��[GM��c�l�t�ړ5��Y���ֆ���,�����)j�44*��>���ꂱZ4��Ә�s��p��B�5{�� ��v���઻u�2 Pe\����x�� e����z���:����,>�1���=����.R�kz�V���ޝ���%!fN�SdNY�\G*�z�Y������{�����x��=��aN�SVuP�d��3��a[1�D�/�W�_*�ѵۺ�p�,�O��%y���ez�\◹C3���x.���E����҂nG2%��(_8�H�m��U�i�`��-Z���6�Oi�"k���Yj�c�"��4�Rj�JXe(6�A�����=`�{�����ՉG½ڶ��G��3F���~&<0ru�#�:0������J⟕���vǼ�λ��1�q��w0�u57��X�]�J������O���կ|1�%�ͩ��ʼ�_�]�j5���j�����ΪB�i�����e]~��Ϟ�A�H�K7�]Q�7��գ"��B�,ҜQ����l��w�A8e�.����!S�]	��m];4q���9/x���m�d&d�t}~���� ���x��Ȭ>"˚�'�4��<�����H����&�����yE�O�&���ܩY���_�{R���N0֞7=����g�a0SO��'��i?Dۼc�$�Ʊf�n8(��f��"���)>�%@��im�YB�t����\�ᓜ�ɞ^�g���qyq�a���٦��n�t�p^ݝ������4�nv�����˚�6
7������1<I�!���H���w	6�ld����ԕ��h��nLJZ��]3(����L,�Wi''g�fc�� ���� xy�ɛPir`��z^�n���{9T�q�E�e����l��}~jJ�+��ӽ�ڵc���a��/�hJ���^��~6*D��(�;�z9r�S�	,�O�Љus� ��;�"=v�d�7k����$m*���"X]�-O�ҬR6s�{�Ι�3/?���;�Ɂx������O�ֿ1��!�������x[58����f��ճ|�o7�IH��!u��W̾s��ٛL��.4�L$M�+5#*Þ4%;]k�ok6Hu�q1��l���CY������{9���@�Z���RΥ “b2=���1b�Y���_���(�:���Q:w2>���W�ږ�^7�k�Q�E5CT��J�tuV�� F�o^z��ecC�����r�%.5���k>�"��R��}>I�;|�<���]�C�����Q���X�����X%g�W�������p���t5ȓs9Xo1��.�u�kԓ��A��V�/���EP��z_�:�j�m�yj��~�2��ދ����~-�n.ס=��~g�+!Z�Z)L̕y���N�e�{%F�)���;JB�#v���܄�^'���،&5KEe�엨.��\��ut,'k�PǮ�������뜣k#"�;
�w��ɯ.�h<Q�xz�	\���!��9[ ����O��U}_ϯ���� xxi7�ʍ�C1u>�'r���OE0���H��G������@;�����J_-��)z����~�z��,��y�R~�b��Un��յ$^C��h��gx͚��(+7����vfVV�f�Ӎͱ<���xǏr�b���e߼�0��Yj�F�?=��0���^)�c�ܳ�1)�}C2��7�	�7����鄝Zx�\��J}�)��js"ha�]�
�YY�gp�z�Zj#��栰wVS�F�)
~��dwL3�p*YG�9���YRHa�x髬�=���`�X
�#=s~��אE��`�-W0��nz(����p���b	�"m��Xk�"����`�õ1��9Nv�ݝ�l]�r�a�M�3i�7�8��w(y���S��B���!�z��F�H`�V�Ik5D,k�ϯk1���/si��y�g�[r���opv�=q^Yޘ郆��ˉ$�`P(oHC�3���yL����n���@@��g�۶n�1������\ѯRjK1�� ܐ��nۻt�O��98A��M_�}��_�*�\�C��#3r�f�v����N��T�)�6�WO�[n�����[4�E�c$E+��ƭԶs��jݠx�g0ӡ��nn�����:��ۊ��+$�r�+�(��8�\H|�?���a� ��< �݇"x���rDH���ץ۟XO�=�ƻ6ݧ���?Qx���3H	]&�V�-��'��.��7��೾�(�|sQ��DA�.3�W<ױB��8^��.TC��k��>�3�S�"�^������6�kmLC���{*ME��+�6I������6s�����F�%�� 2w��0��;���s䂰�Ԉ�H��$�-x��q�T%5]בz˼f�Q���=݊ۉٖ�C
�*Ԅ�@%t*׾ǆES˥
@ۏB�4�Q��<n�!����a
ƭnn���3�U�}���V1*?SI��)���Y�.��<<�[㾧�d��]�b��pj5��w�LS�z/�Jz���`ϞH��<E�2���2.sڦۭ\��ݎ���H57i}�ά�o�� 7����u��8�Tx��Dr�^Ø�兀UJn��e�7N��������rq��/{��<��Ɉ��5:!��p���B��z�xW��%�x���N����K;NNĥ6g&�է�i����Z|�"��8
����Z�-����z�'Ӱ��7`}�.�X ��f.[�"������ ���k{Ey�.�x�7|/rnT��d�.�ɼydi�)��Z9��.<���Ѻ�.�e��ඕ�����%�'���s����.�n���<�M]�o��e�ɻ���-��f���^�������� ~��s� ��v�u>e��Hy�Q&T����ߐ���"��ߔA.�z����?9nw^7D����*4��s[[��=���ŝ�;�a���T�Xe55J�����:�.q���J9[ ��P0F�Oמ�-vc�d�%_'*yq��sk��w�Z�{<b�;���#���p�G��>D�Y�3�<��M1(����P�υ�c�y�muk~��v	�g��#$Vo��S��i޸��1�����]" ����_@�!��h���H��\ȦE���h�y�ζ��wV��/ZL�(`���r<�G�Ȅoh(&�2���=+$�K�*�����`��R���}�V�rPH���ދ_��_����5(�q����t���R�)A�+ڠ����^Q� lh3!���9=i�s����5�������rH����ޤ�j��ҁ8�ݼ��Һ̣�Ք+��z1���m��0��*���<JR���	\�e�yH�yQy
�����{�~�2�/Z~��y�E�d�c��SȬ��lwD�{�2j�ɵ+�l��+�k2���9��å�TѮ�U:�X1�U������G�i��[��N:x�Ŗ��5�Xu_�w�����Vmn���<����m���?j^~ڝWk���W}�[�;{��ɍ�9�'K{e�M��M[�r]rV�Ýb��4l%b���������������u����,Vv�k���xi�ؔ�|�]������f>���w��k�KO��8:��VP�ǲ�1�܊9O��x�s��Uy
��" Y�D#�Rܓ�q��\i1���Gq���)Up�����{�s��&��y(���[��cjrr�v=�@3�0r�=~��WWd�����識ά�d�z�
3�fo\5���:�O��J�/id��YP��4�>xk�ح`���������tk��Ҽ2�2#�ʑ��ި4+�/WX��]!��A]�:�����bL5u���x�޽/GC�c�0,�P0��/R���R#� ��Bۋ�~7r�S�$�e�b}n�H�ix���S9x��e�c.���H�X'D���PcS傕j۝4/K�L2gOīv��B~1�w_n��]��=��5����_M肖ȸ$�҅��r�.;LW�=(RjG�*XQ��W����Z��֚�%Us�	G�Mq 鰑7�R2��_HN�xc�Ʃ���¸݌s����h�4���?�hu��t�D�a�b��sB\�v�C���aޤ�N�ǂ;ro*��[�˲��"&�f�6���ɻZ��7��qm�X�1�AL��
���lXB�\g]��[ܬ=s�6�'i�'fÏ!��}+z�Z��*cd�ĝ��j#���O+5a���x�����\u�����n��]�O<��������{�����}���[a6]���_��2��6rw2��ޜK}�/�����~o�� �(���Y��
�ߗ_:=�X��3P!�s�LLx�+��qH�do+�q��5��y�T���q��J�/.T^E����t��?��:aׅ��2Jz��ql�v�C�UC�a0�T ۶���i��!�qU�_e�e��IH�>J�V��>�T��DY�b��殦�-P��
�m�օל�YH2���q�?yU��,�	Ӯ�g��F����;P���ś�Qо��R���8�;�V.�q檍ͷƺ[.0��QI���m�gg���CT0��vF��m��m8�������l+�g�q�
��_��çb�;Y��>$��+^i_P�rr����H]�i��p�٢�n\�2z� �f1�R�ۙ��f��d\�{%uP�n���z�2w����fmm���f��DY�L���BԵ?^�*
���;��[�R�����^�ۙ�S{}�o��y��7�csnrЭ�:���V�VvĨ�0�Uo<�؞EWa�.�֤�OF�F݈�C ���*��#j�P�Y\���U���% ��ŎA�ɬ� R�v͝�&��m��< �{� ~�u(���v�[X[�K+)�"+�Y����i��G��$ǽW�;p�`[#L��}|�����n5V���#9�����U~�����o ��M��{ �����t�L�i-��Xk��d)	&>.0�LF-4�s]ស�o2D(�փ6ɋ;Mr���5x��4㷣S����,%:\P�2_�|9w�( �Z�J��J�0:��oN�פ*)�GOQoW�:�n%&2)�i�P��8{��"�@�=��)�7�o&wNl���0�Z���1c[֬����L�&y�D���愻�Э�Pm\��7x�o��O�GȽ�c9�]��	���>�U�^聄?YxY�ql�j3�������y3g��[wO2N��u�D�����=�t��5�d(�%��E3߀����z��[ݸ�Ke��n�R�!	=6�iͳ��t��iA�k��
ہJj}��dV��G��<�
�5p�LF3���ˍ=
��(k&�Z@)�H�0��nC9Om@FA���w�J���Wm�s�P-4!�.7�\��km(Ah��Ad��XwhT���l�D����2N���*�̼z=��i�Ez��Wu�j�Ч�J�N�؍[#�g� �6.�s� ZXp�{$��~��a]��]����ɲ���)�-����D�V��r�g��ӑën�
ŉh��e�+r�>L^��cջ�r� [ތe�N�u����Z�LF�َ����d:�ʃ[�I���e�>T�u#���FK�ÜҀ��^�[WBtۈ)`^V޾ѣ��JO�c��\�8��2;؟R���5dᄤ))� ɡ�-h.n �;�Ȉ�+���[:z�*�9h*��e��[��,,뾘�|ڏPw����=;�l��Ji=��;�;Iv��+
�LH��ګ�k�̤���t�N�]aյ3rbtr��q�S��=pNxV�47�Pb+{{�d	�G8�[5�3�	ۡz��m1�B��)��+�T#'9I��{�fv:�[t�ߥ�8>'^=���(�p_$���$�K+E���vV�y3��+S¨��i*��{b��yGC87��X���]����ŷ[�n�gn�u�X�̳�{N�X�����$PEɈ�{� (;F�e�n��¯��i쭻[z��Q��7w�P�ڋX�'gn��%6D|4jO^m�_6�c�NM�n�5Ә��mr��
�W��F�i����I�^����w'T�ݬ `���: ���qΘ;#W]�����z�����>=B�cK<��x���;X'�=쉃��&o��S"��L{�vk�-ξUn�y�ꛗ5!-6�8�����OB��M�<����jhq�.^��u�lC��]����Ѱ
�����8�W�~�s�;C�d���o ��7�8�-�:�6�ے����^\[��^ʁ6�&B?�hWn7n\[ש�̽(.�.��9�Ŵt)�4��C2���o	
F�x9��d�y�J��� ����@v[ݩ}#�x����N�Y鮤|�\�ڴ`���o�7�
ùF��������/v%Z-ݸ��q�ٰ���;��7�W*EG���;�q�Ɇ�,@f�.8��!yҭ�v*�VZ[��p�����fgvH7eA�*P#��)o�n#�J���y�WX��<�X��WͶ����%��JQ�����w��:�x����U���^@Bˮ��pNuα�h�.���&����s4�n9�^��64t�cǦN_q�eoH�:�RN.�o��@�S��W ok^�� 1���[u��Y)t�\�b:�s�Z5e�du��m�ЉI��l>�n��d���)}E��������[��>.����$&aqǽG�]7P+AUz-�ə�ݹ@n)b��b�{]��]xU4-]'3`*w��\�����b�%��ԏ�PiVV�U{A��g�&nӐ�+�딣G�?�o&�t���m��B�v�K�$T��Ɔ�SV�`�5L7�gsN,)�JS%�|���sVz��s�O��x�#�s|�,��s��H^�#�|h�;�]����E���e�nQ�Uՠ9�9$��oD��wQY��u�.WA�����4<�����|������܋3"~K{<�eTh�7�C�%�9_����.��\�������P����7��;J��u�S):K�yBs�BB-0���L�I
�[������}uX�FG`x���I����.P�,6�J��8�IY�\H�E	���eY��r�I�&S�}�<#S��P�(�P��Y�S��$���7��y1�g%Y
�JaEPz�Y���v�X�W-$�2�l�DG�)C._������e�J�eUWԧK&�.E�\�$���	�I!j�!V���[�UJXUw$�E��ZlR�B��r�9QQP�nz�R�֝:F��u9�$M���;��+U����s�e�C �$eFd&gI2N��1j���z��*T�W0���+}r�;�IW���N_��㡆֝�������M�H(�����@DSV�Qf1�`�ή6d��}5!eJ����bۨ����K;�̩�j�	��+
,ͫ=�h�5ɘ��noq�YIQ��~H]ϧ���� ߳;l9�o����??Qq7�wr�$%�=7�Q3J%��Թ,�^�4	��l�XH̦G�gˬc����bL$_`��ĹG6v�,��?���Ǯz(%f3�(�L^��!���X{�b�^��?0�hW3�6OF!*��Rש*��d���7Z�p�Ҁ��r��Йܸ�򀯧:(�t�O�^�}�Gw��P)�mx'���i�x���P9 -�Y@���Ma�v����-�n��͌�W�Q���r��#s	�`���߹�qy�@j�+U�#^HBC�.�{*{Ѣq�ZV3m���II�b�M��{\|}��I�p2Sq�^Bk���r�ժ=�و �P�{�.ae����@L��U*uq�Fl�Ѻ�Z�{;�)�<����aU�G1pr���׆��E�8�e�NԌl�Dh1����X-SS��0��!_�^��+��v��3�ig⻔g��b<��5�t�K��mv���"@���(Hq|��?Y��q��5�sv��`+�ǵK3���#T�P�|aϚ��@�5$omA7#�wfP�8l{I��}>hv:����莱HI����K*)��
$V��M�� �sJ]�W����nP���3��]4GbD�L2�ܬ+�7������~�$Wmj� ��,К��>�xtH�V�U�����Wa��aW5�Lt86�8N\��`x������y�=��o�{úqi	[�ɛs�ô�p�7Yx��#���E�~��/�'B�����,)�B�J��!��9�=��]zj1�,�&�̪��n�N�@i�1L1�ڭ�<�t�V�K�ٙ�s�>��g����7SU�@��	��ț`�r���R��)�_�D�W�e;t�¦�(�ՙW�;�ڈa�J�P�v�-��"��T�eVg�v��p�C�yĖq�'�ۧ^���gkl�kA-�k�zu�m�.�k��7#(��o;�(	��kh�LIǍD9f[�qt�em�vڶ�u�y/�ؤSmy7Y�͇��������8F�2t����S4��]���"ސ�Gem8�g�k�J"�^�B��V0֮99@�{.�g�a>��}���MO-ۼ�Fl^�e�|����`e�AGw����8-KWxo��n�n�H��9�51�cqV���y��	bT;U+A�?yA�>��H��47�/�e}�#!Y����{�I��Fܮ{�d(�W����I�I=�9	x�xh/�}�B���"��s���˔e�7�֞R%��*D�VjȢnJ�PY�^��H�[������Ƕa��	����+7�t9�O.�%m̦�;u
-en����=xg}tE@ձrsD^��ы��%p���A,�s�셆��w"�+�q�D��5��Op�H�v_X���yp��9���	m��$Y�{��0 y�� ������?{�����Ѵ	�s� [D���U*u~9���z�EW�i�%��tힸ�=1�7v���i��rr=�3\�lg��vųd��ҁ���L��2��40vn���M'5\EL-��;<������dx뽑ĺ�M�5��I$ܕ������9�"�x�Yϰj�X���α̃��e�۽<�k�fˆ2!��A9�ha;0�f����(�7?d�V�O�/�q��Q�?�-_�g�<P1��tx�-�3`.�*7|vg���:�О���=��~z)���`���
O�~��l,��ڙ8�s�?Q���4�'鬼��9�ȧ�|�����S���W���U*�t�ïu�a�֘/�a�9�\�oUnA�;dI�{b�J}��v#g��({���?]d�|�qͰaV�p�6f�ʫ���wwt�t\��y��y�wB��]a^z-�x���_H[�P7t#)�u]ٱ6�\J[����;4[�%�<��Ô/m*�qw�������|�N��og��28�N�[8VSq�ƁZv��5��\�f��Y�	����Z�X��tn�M�ok���WV��i�JU����Q�ټb���7ku�{��g{Z�}c�wss�$@��Tئq̢�5����-H�D�<�if9E5N��Mw������yy�<�<=���}}�AbXpVx� yY1���Ͼٞ�'�Y�O�61,6s�ĕ�G(øy��)Щ{��wO����^�1�U��Öи�@'�n�|���[M�%��n@�Bx�xX�;���o�E��� �LnDH��vU@Vx��x����@]�F��n.�׻�T]�R�����7���[n]��iI^��DE�����ga{���؞EІ˪7��옵L��M�5|;�d�A+TX_�FK$�9�P�ϭ@�EBBɀX�;EZf:�'�C��ݡK����=A}^�	�b�w*R�l�P�q�����ь\�T9w�@� � �6]��ǚ�=g/;u8��b�9ROGJouX��<��C��D����Lx�\H;ѧ5��ϏMX�b�{W�<�d��$B��_M��zt�>�	1�o�y�^����.5Q2q�s�U/U_���v���M�&�"qR�'>��@J-av"�з8dl@�+=��G_5=ޘR���Q}��(��&�
Z�ĕ��#쏍��D�9��q�* ���=
.2��9����"�9����g=���[P$)�2��f�`0�gjbI�Q����\3@�`9�Vq7B��{r-��d�	����sn�wCo_pM��olb���έY@*��+�`��<��{;����o7� z!��E���3�@��3�Z�/È`�c,s� �>���4t����1xS���~T���u��)Emtȧ���P���ܻhk��P�9�ֱ"o� ���#f�ȓs�\���mZB�D�؀U����ur�ÚW]U��*����P��BԄڒ���p�֌]�[_���&���2�cjJ�-l��n���<��ٯޅ8Ĩf	����Պ���]Т �/�7�Bl���c�;Sz�\�l��pz���kaT</|~���x�X�tjB}q�n�*��qQmJ��ޛF�+�=wu��6ދW��s�gzQ���U������V���Y>�Z�913G.���Y�m��~��OGTٸT9���8o���\c��D3�;+��ii�b��0/V�7S��1�U����\է֟��hs��O�@�Q�'_u��k�N�����ص�^���Bf�pؒ�t�7�	�D����K��D�׭Ql��_�� m���3�T���!���W^�F�1��"_LCn{p�kk:�KW��u�-�X��3�Z#w���n��&�˖!rL�x���t�4`ҫ�
'���v,SJ�:b��S�����ů2�s4H4Y}J�]�7����V�zv�6i,���A�6�W;�o3n��kOL����o,l��ܾ&��-�z�bw;��K
�/���GD�P���Q����{�7�<�a� (}�1Z�}�@��\�?�kU*u3BT�2 �ͯ^�v��Act��P���rwUN�eAPe�:��������B<�� �r"�O�J:��Z��m�Ѓ��׃��~�#�25ݴi���ג��b}dԳ�j�h)t�8!��_@���&/�Z6���^�[�k���l!Q<�սh7\n�F#
UϨ`��Ϛ<�F$��p�0ad�7���u]�&�������f�ov÷�m%�����Ӈ�����T(6`���}�1���W����{���5ʀ��.�s���3&`�k�c��+�rH�9��C�)���!w�ԕ�d�nZ�� �&�@u���|Q�sVF�g9��{�����8��������'0�����wӫ"z;7���QYJ9P��f�]�H榮�C�3����fzsdğOl>�^���Ѿ�L�c��X|�-(9��8�x�J5M�6��Du�P	k[��[ӗ�7I���Wn��N�熨���H�Ԣ��S�%U�"�2>�I+K�p�v���U��LV��}����$2��Kz�@:w]��|�U��*4FZ��זm�:=-�l��֐�#.�Φqf���7]M`�󃣨2�lޮ,]�:��R���e�y��m�H�c��*��V�3]��4��w���Wu,���=
ȶ��p�YU]����y�����{��Ǹʅ|�4���	q��־�ӓ��_U���8�=}���1kZ1��}	�1�
X�Wnق�T�����`e�A��P���>q�8���ڻ�7�7��x�#%�F�"�E?S��r�S#�1sV��,�{T�;z�M7(�L��}ҧ�OU�e��Oo*�o7}����� p�4��%F�*Z�{t+��@���&_��4����D��hS,�t�r# ��z���<��"]��IK���"c�yW�T�|�)V��ޡkV�d�/]�D��۫R�2�	���W��;�"�WQy���\=�%����z26 4���l�gW-�GkU��P��Z]B�X��C��>'5\�:a"nY�C�vCg�K�X�on�Ă����׻�CN�����Ꮐ�x˧����=�G��@~>�R_l��}�W#��[Q�\��g5��D�{#��uZZ�-�'��,ʹ򌙁��E�������6����ԥ}_�����k��Ýs�UGI#�m��5��ܛ�J�S� �w��?O�����t�/�_mZ�p��"��<��-����5VwC��|qś}A�*ok��B�{k]�ʶ+�ɞ�k�����^گd*'xu��������a������e�'>�9���tA��� �նN��4�(q�u���j���o6�I��7,������_}W����%�I�^�T��J���ݳn�͎27�T��ƲU#��܎��ޅ1&k�<�-B�
���Eox�q`<��&�c�IK��PvR����r.Ҟ��}k��Vx/Ô��M��˵�B��r�핯xaP�j)>�K(V�"N<�P�mB/k�n~w�ݧw�|�=9>݃s��ض�����C�.{���{,>�V닿jچ/!�:�F+�ٙ1Z�<�Lձ����cL���=��X���4ZÙ���)�'?0�EY�h�ܚ�r9K��g�x�!FU܉�r�P����r8g�s���rV�|����շ|�*n��^O��5����X��N+�r�ԩDY�	����YjZ�|�*ޖBG��^�.���z���W�'v��T��;�l�
�hW:�RS��HQv��gj`3��S�+{ba/&j���ëe����c:�!��#��x�k�H�n��C�"�!d�q�a,ZV�	Tf̆�*z�\�e8�+��*��u*\e�������g!��Z�:+�$�5�9���B&1�`�Y�a�]P���TziS[��H|�[��o#��4W��/�[����ĥ�q��8��s�CWZo��Xt����T�y�t31�OgM,�*6%�:Bw� ]��|Vob�+�[���][��CuT2�]6���]��'ے��ڭ�ؘ���x/7�o7��=K���z{�߉�Za/��'�F5Bf/V���ll�{	:�ny)1�����MSkP&-���L$���]kieJ��y�ٶA�5 Ҁ�r�=a��$��Tȟi��:E��jrg�%�e֛�ߌ�Ri��Zx��}�/I��?�$"�H�(:�PK^#>��x쁶�l@�+j���DC�U�z����TS�,��_��]�)>PV���A��3B��!SY s^�*9s��LG�j�rG_�tu�I�FjZ��V�"��ltQMHمi��щ�D|�:w��1��s׋Mc7�7��\MG�����F|<2�U�9_k&�ϒ
��H�f���I�4�"=S�Z�z0"ѽU��b�}d"�m�K�jۙ��Ҫ�Z�)��HM�䮅c�խ"��҅3�Cs{��S{�e�^-->-j�>�g�0
�h��i�XĨd�F)�]x��ٕ�=��<�Cj&=y'y^�M���S�P����T�R��@J敋��Ӹ�6'��7fYyz5��>ژ�i>q�w��i����QM�F�I��[<��!Y��J7S�������
�\,{W���8kf��y$h���v�d�F��Ѕ������Oj��A�e*�v��'f�.�^�U�72��.+R��Nj[+�1�f5�'��v5����9�N��bgZ�gV�\N��x�F��*�H��>��|� �o{�y$��*�{����Jt�
�gw�sF�
s��A�ڛ7��!*>�9�9�Z!��%�ks����ߦ��By�[#�b���$���qv/)��ˣ����Z}�����������"ʘ��کTZGd��0��6�׆Dן��&��>�&(A*y9Q�8H�z���~z/�!gA�����-���x0Uj���\sn�Tr������hf8��N���\�W�M�Y�dϦ}���y�-�m�&�T{!I��PcS6%I�#'6�|�km���������j�ݎ���k@����e^0����h[����|�J:��Tԁ�[CM�V��d�u����t�Z�^퍣�F:�<�O�2�@��������.7��qrG'B9}�8�Tɋ���xޚ��q�]����H����!�F4�����Ϛ��E��2!�
	��43�t�n����������F�j̐�ûV۷c8-�D~�N�����}n=UF�;�b�����M�8ʯ(2%�#�A�V]]�Ӫ�!��F9�x�$Y�~2�
���)HT�b�G��p}��2V�W�	�	WmX/���.$�d�V �
�WN�b��xz���#���vҁʛ9�}�v��:k�5B��s#	 �\����c��eVl�S5�� �$���%>@ӓ%7�Hj\*uɥ��F��.��r���-�Yʺ����V�N�����Ym�8ܼ7��bѺݕ���H�r�-yyi�6M=�j;/Z�.�>�m(jhӯ��խ�7�ƭ�t��դs!�^e[�l7�Z}�& u�w�>��C�Ѕ��ԤZ|E�c�m�٧���m0jF�.���Q�{}\�La�S�4�ޒ�!eR��G4�X{��\�z�����*�hwz��ܤ�Ƶïx�&��w���I�m���\��f��;AV';��(�:A�e\L�j��pJi9{\s,����a3�{WV�nX�!��r��T%�7O1��ל=m�J\"<�-��[n��՝eJ����a�/��9W��8��LwU�ڃ9��f���w���s�(�]1IU���+[K8�꜄����<�WI]R#�4v\�z��vZE�S�YuǾCokZF�b\���7o����s�Cw��X���q>��Sr��ꤜԳ��L��Woh��&̥vG���ZDZ̩�i�]Dq�1i�M&�{0����CX����A�S4��z&yV����/�+w6^n�6̹G	�ڻʉ�(7;u=�䲤ڻ/�Pr듰��쾃�,������U��>~7I��Τ6^PJ��a��)��ԭ��@4�mYUH�\w�r�����(X�3ً?����N�Q��Ss�뜒ۂ���钑��Z�rn�M\U
1��"��!�I���:Pn�.�{:�h �*8N��<�S���j��o��͹J:��$5��B�H����cu�L�V�4&�X��ϰjt���¨���N�N�ڶ%v�M��|�/tB-a��0Y2�q���da��v7ں��H�����q��:�^��C��ڷ�.5�d��>��>=��J���u+.�byxgl��1�X�\y`��A�N�Q�T� J�!n_L���D�/`Fe��тt�l�4,V��n�u^���#%!�p�����J��"8@6vd��j�4ʔ5�M�'l/3�ft��n( �uc�C�*�bn�f��5m_u���Oz��㱬�(�����)�vn�n'���˘�؍Y������[��)p��űu��Yj��B�/�Ļ�r�V�a��Xd-��S�ƐjYږ�Y��i��ڳA&�Vٺ�ŉQ�wn�ݬ��>ȸmm�[.Z�x�#w(*Ltѭ��1�Ӂ�^��q�ܙF!�Gz7 ��Qv����F���'�$��V��!�d��+�wJ�.oY��=�I���~~~?O�������8�DQ�Y,�-CA)5�&�K*���gs���@���Sm+o����7��ʧ�hY���.�Ĥ�R�E%I6ReI�e!��RJ��d_�v��������z���Z%EDUa�u�$�TVWe�G	�IR�dȞ�NE!Re*$&V����tMf�R�.UI	d�t��TP��]�޹�e�����1Q�qԪ.uK�)͒j	U�
��4����B�̼��p������Q_uü�SUXDiZI(�3�x�L�*�
M��n��"��T�t�U��8�ݥ�*4��wr5�ui9��rw-��8�#͑��G�VDES�IZ�O<<ڭ��'<��B�8�UU_�;�^"�)��\Lz�����T�YzЈ��AqɈ @@�A&
"+
�+�т���P�IRa���d�:ͪ�=��/kZ��t0��gk����9E��P�z������y��x)luUA��t���N���:� SL\|^%��׹Xö���>Rܦ��%��N��Jv6�Cؽ�9�z��g��L�����#�"uR^�Bڐ���FH�Yu ��U�僜�㡲�a��d-�h�}��ͨ�l63y,5L[���iW<k!�bPh)�HK��zE�����%l��w�ا1�i�b��B➮�X3��汩kxr(�n���0�)�z��>_oE%�j����Mi}x����ذ����q��z���}��9ֽ�n<ֻ�|}�<��a����Kʨlr�D!�5�><ӤB�r�� �k���f�nuC;Ove��*OI� �6��ؖ����)�2���7�*�]�^�y���"���(�T%0xϔ9�P����t�]E<{t�|���(�сsȹ��݋�vy����1?ߣF>�p<��.��y�Zz~T�N~e�
��λ�z3Q�M�<^_D��D�t2-$rb0	Ƒ0�yP��)'�j1��0Or�^��gs,���ư���'L4�#��Zh_A����#�f�Q8�ȵ�*\���w��h���(G��9L�U�f�4�ϛ�6ż�{�Z�8�Y�3����ʘbYW�9��a�������`k����>4M�S�śMе�\�g���k����Ύ`�<n��y�	���=s�5����}s3WU]����� �  n].RL*A�c�c�>��МΧ�#C��ΡR洶��D0�7��������ُ��(!�s^��n�U�48���#�X�`����mމ�a��3e���ǅ6��f�����ݖC)m��P������l��{��E���{�w�y����)
��W�++��m���~Ͱ���P'�nDL��/j�/�.�j��(%"�0�bk=G��v5y]D��^%���]�I;��㉅8�/t�Tܶ��UhSn,������ý��vG�����8�@s~��;�#x5ϒRO��.����X*�E���Iee*��{��̻����ޅ�A�=Z�O�Y]��ܺ�(�yr�l�^����4��%t4�y����j�����4���eN��tĖ�%�.{O%��Ȭ�kuš�.�kz�T�Qf��\kt#6w�N��z/�YB��q3�8x��Wz��a�����&�X�y�Ⱦi�9���ZONM�(��3z���aDQ�w"D>�j���\��H'u��t�i����d��D��-v�On��7H��>
�H��مpn�2+��Ӽ��
�ْj�s J+��p7���=�E�}��!X��	�դ�l=��	�^9�M&��bS����<�%kp�!L[�α_7�u�[*f�m�D��^��i��/���ȷk�����o7�����D�C7Y3�7�8�p���~Kk�B�펹�؉��Β��/V��wUR���*_�Eر&o�Pf�j���f�u[�jK��.�t�8v�9�))"�R���%C;3���9��1�tTSx�Ⱦ�k/k�
��#��x�F�p|V����!�UX�z:ĠUN�������ѻ�olD�b~��#ݜdN*�8�ޞOAdv�~�r�Y�<H;շ��'��_`����>�XόK��P����Iv6z�z�I�cR3��Z)I�mnx�q������ݼN�G��(_C9�U*�����L$@}k깦LhwZ���1�≂��r�]-�&�O5yf4���s-1���(�|69�D#������A^;x�
�w��[�꥘��X�d�⸏��<����ĕ��D}��*p��' ��%?sp�v0B��д�b�:�nl�E��G���b�> �SW���9?�"�<7e,Ǒ총��s���Y�-z�,���>8-i�U�9Z��B���	�J#�u0c��?���������V`�j�U���q]e���!��֮`���$�ɞ̫���z'��+|�8Tq�f�20c�ʗi�c�Qꆭ0慜V�����3v8�u����/�+cp d`q(F��].7{�9U�^���������g���`�o{׺��^*%2���.[�B�-R���U�89���5���������ʊ�vsl�Z�ګ��5	�IY��|eoO�!�U�sn�����x�T1sB��-�Ȝs��~84{�;�s�����ޑ����vT1e�*�Uh��<ҿ@�r|�zg��	�$�Lb������T۫�U2+���޻�!�[/�	�(%f>���t&e�^�!�Q�[����K0����[ջ��]s��(�1Υ��׎W��j�^5	raGf²�_p�9��b��9�m�.C�fs�y��H��4���;�kO��ӵ�^->��EO�`g��ؘ�Ql�`τ��_5�[���Tc��֏dKwb�oga1B	S��
 �GH�T8�Z�f��6e�O�ouc�SY��\C���O�
�7#-�v7Ri����.Ɋ�=~1(�y�*�T�󦽽'8T#ldsg���!I��U*u3R�ᑓ�^>uε��	9ˣ�T�5[���/q�|�~&c��=(�"��0��>U��u_*�Mf/���C�}�k�[��������g�o������)=]K�����h�/w����\=�b���*4���Up���@���h���n%�݊�ɻ4��(r���ݳ��u�I������:��d\ŵ�H�i�������\�u�7��!���1�[�k|<b���Og���d�M}�0R�8k� ���M�`L���.w�3�+ӽ�!��������X��\���	+Ю�S����F�;g3�f�h��v��;�dm���\���Fy��#�ֻݱ�!���;u��9[�E�Ϛ
�uRiM���P�.�T�:�;�i%e<PdN�g�Bj-��O��wj��I�h�$2�r�a�����=�f�E�{s��玔H(��fR�a@�R��"=�J�k�.j��cS^�*Y<SF��fU2�n=���h��$�o�5kv��vG�D�T��T+� 9R.�&�,��Sȭ���R�֢��L�(]��{�M�1�C,�5,�c~+oD������h~�P�u��+HIH�;�UI]z#5!�UY=|�4�Ǩu�m����5E'7�E6ג�ǻ*v��]Q��8S4.��p�[ޙ�b[d��v�헥d����ic�H��J�X�R��(���[ַ׬��NC��8�"�	�B�K����4��b�XO�6g����i1���u�����>�@�oeg33�is�L���D~�C�y�ϟPh��!aO�ξ�;U��wt��)���2��kY���}O��KDҶ���S���a:��NKi����B���|���Y��Rb����-�N��j+��
.[%��6�	����wj���~��UU��=J��pߧ�����"�;Ã�^=	r@��M7��}p�Tkw����;Fk�u`TwK�R:��z�� �ex�~適 p�5�y#�Tn������"���t�B�&�W/7*�n�\�zY�^o��?e�����J�dZH�X	kH�q��Ƨ�z��!߫��v���t�w��V�v�mOAfϮh��y|��4��+O�O�[�nA���a��QX�_�yP�c�'�[iΑg]y(���g�����%�pϏ��6��*1#!fO�����O�Y��=�;@��{Y]f',�0&.��5�ٵ��'�R��|�Q�AZ���p�lO^��������e܌P�;J�˙�>�˯����4��I�%r��
:�E%|�P�6D���ִ`_,w5ļ��A^�bj�7������qWp�&G?R*~��>0����\J/H���/~=L��:��o�'���Ae:��7v��ɘO�
�n3�l����ۼ7eDC���:M"��A���
�=���ڨQ�n��i���"��ޞ��1/+6 ��N!����Ӏ��; �2�Z�(�ћ����U�V�e��Q��Bn>����_�R�w��]�9W6ց]oB�<f���ܮfVɚ��"��lӓ�/zD���E�_|>��{ޞ���*ݒ��ظfv���������R�'^����֢���g��F�\�S���1�8�p^ߥ�,c��}�ߐ���?�u��zɍ�??LJlk�0���I�H�ҫu-3q��Q���]Q�f;��7��(�?V��ߓe	�ˉr�i�Q��ŌB/�G�uᮍ���q�B��sP�s��������*��	2��O��U�<��$�;�i�J/(^1�D?�LL�,�9�v�딞)�?bS�H印js"+V��E�a���vyKS����F<��^񵎷q0��"�:�y��zqΜ�փsRR�+U �,�	P���:��}�f!\vU�r������ס�$Uv2��U�.J4Y-��0�j�
���P��z�^�1�G�{Ea�^�}��*b5�W�`�V*=�;8زT�B��Pӵ���79�P�.V�
�Ωz����~��E��ٶF�b P��d��y=��)9��]��[��u����k�%���M��릓�L���b�/m��<SU���
� -�
A�dL���i�J���������7�!�Q�����i������l�]�4WY��ޮ��F=�Sz��6h\��R����W%��J�z�sټg�.4�a��?��g�S�ɻ��<�إ����!���M�vc���n�#�ƆL3��XK�O�fl\Z�{��h>�y��0���|�H��Nf�-şگ��W�xı���C9S[�	V�kק�SW�Дz���$N*O�Dd_+�Qk��_h�B<-<=���[�kG2 ^l-�#\&C~�h�%'[V.����s|�Kn�����nacmt�cQ?awsзW4�s�c�[��H�!���/��5C]Lj�����&��Ǣ:o������I0^��0*j-dc[-���`�g�h�_`�(Vxk�H)��#B�Y�_A:�~c&%���ao���B�NT_�q�U(i�����Tp�1�8o�j�?���䘇ǥ��[߿c6W��	x��}>5�!�W���5�l׉R�����ߧkH�켍Cum>�����P�2�)V�5P�ԥEکM���h�[@���p�ݬ�نw��[>���}2���Kռ9��l�B��J3"^C��wƁ���+�2��lس���,CE����L�a�xq�B7M�{/)�
T���%V�V���{l.<fLG��=e��H%�~�6.�wl�G����d�x�C�E�4����}6֜���EfK��	��������a��0���1\�e�j����������QBV���7	���<��s��մ�Ӆ��P^F�ݖP�� v��+�\y@�؁�Ž�����8͑��=�7��;+u�@+lbg ��6.�MΉ�����h��}�����.����͘aO���Z���v'j��~��q/"'��/f �\�c�N-UtfE���7}���U�դ���Jz�T��$DC9��NHɷ�6o���MN+�!zV��U�Y���p��x�WdK�;�Ⱦ�r�d� kvo/}*q3_h���;u�
��*�9�N�oa[vޫ��垒����L�X�2]�<��AoHRC�BQ�|��*�B�.����9w��N�(�{m0:}#Ʋ:N�`&}��^:F�I���R�嫵����K<!��e��)���\�ܹC��_��a���s�(�N��x��p�ڠ�(D���9k����%��y�3��f(��ܖk�(^�P����s��޹Gx��������NM�Z��U:�n��V��TX�1>�ԙ����c���h�ʨm�2��ۖ�v�$yW�)�{��$Qa�
{=I��Ic���ϟ SH��O@MG��r@�a�5)����D�e��4[&sx騭�M������4o�R"@yQ5R^�LLf*T̏P�]�i�Vi{����lŶ�XK������X�@]�*���<i܊�̱���a�!ͱy
�L�2���O%��ݚ��u)��+h'un�h�g��Q[u�s#:����H�U���-9��i�k�^�:ⰰ�1�y�N5p��(�����Y��h�=K������a�m�(ۛ��x}�o7��k2�Q�3J��B����xa��yĞ8ۺ�����y6�@����7f�"�3]٩׈�W�Joɫ��u	
CŏvH���b�|�f��N����[W`8Ð�z�RtEq����d��i?����{$�\0`{\��EŹ�G_R�NJ"�@�V���v��'��ײ�ﶱ�&���U���g��Z��&�N��0u��� =��-]���Y���B��{r3X�M���z��`{BV�\�z�	\��3��.ӹʥ���Ca�6g���#5���Q���ٍ7���?}05%ad.�BTn�����
�׻	�X��<�Wj���4��-��#%��'�hD��dZH��`%�"�8�J�U�`a�Q�t���5d?B��礪~%Ra��t�T�'��wMi��7*>Zų�E�}�9oԼ7�L\m㩽~rP3K(;q^Ǣ�mp��1��@K�K"�Ў�*�U75^$֞{fU{s�5ܕos�y�|x$L�]�<�hH]k�\{���crGp/N�L��������-=��	�󋦱�;C�
cy̽�7�w�6�،lx��mk�ׇ5�/u��h�";��w��i<�m �hX5I��B�5)[���뛾�c�>�1;4!֩�����mne�Lr|�q[m�ݭ4c�Ao��	���ط���ᢞʽ�/���{+ieHRW�!��hc Rk3�����3,)����r��7�ES#������;Vb��׶v�I����V����Հ�]t��{��\�P��Ş]�YZ�e���y�B�����y�(�; �5��/=E�T��<]�OP�(�m����nZ���uwu}8�i̫���FD���G2b�_\?L/1��-��.�E���5j3�!z��[�fsX�ZEuևq\������*B�HՔ�cF'��&%��p.-�8���gVH��z��?z��҂���ڸ�Q�׳b#0��Mu�E�8f�l1�R��b-o'-ݕ�q��|'p��s���[�Z+�[�	LF7�oN�w�;�g��E^�^Q�uj�K���!�t��� Gi��z��nG�,p���ؔb3m�>�q-��7�P5ǟen�#�L�[ޒ��5����F��;"g$���R���ISd�ηN$"f\���4�ʝ����J6�X{vq�_U��F����X�4�NU��8�]>��:6M�WR�2�U�Uw�V�#�m[��e타I%=͹��G��abƩ���� �~��G�b�#]-�����J;�����JS���n�>c��{eT�t��{�[���(n�Ѣ`'0=bU�w��f��<A�[�C�f��ձҿ�c��¦56T!.�*p�`岅�L�W 52��s���I�Ĭ�.�S��*�����ȵ��5F�m�f�v�p���U�������f��
�ϛ����i�X"�#�51�LGK���]��yr��_;kT�c�&�ʦ��5.���U�5j�����.�̼��t	]�����{w2�J����\k�8�>yux��;�Ö�p0��4�ݗ�֨��R<�������;���{��u�2}b��O�8�vZHK��)qۄ���	��,�l��8�� 剥Й�r��zuYF����s:uq���̵�C�t뜆�{#֬��9F��-?����k�� ��N@���]7���Q`�c�	X�VqZC��@���Y3v��8��r&��w��#�JA���}3-sb���K*����|�u�q�3���z�_6s7e0�sa�73I��YJ�q��&yee�ˊ�N����k�Ss����QX�� ��P�oWZ� �Z��`�A����#g*��F��6c���j�E2���:¨�����u�݊�����L�ݮD5�s�3V.����^6A��fu�g[?HN7r��O�/�m�+�B�j�����4�z���w��9Y���Md�������;%����K�HG3��d�A��ۊ��.�g��X��\��/���6,���{���UC�i_u҈��]������7���fU)�B%JE�p��*���Zg�G%,)5.�rvU�GS�|���>dQ����|�w��+�T��C�P* ������ԲJ���˪Rs�4�*^�;�j|�8��=k��Xp�i����,�,%�nG���Q�Ĺ�-�]���V��8Z�E�5�*����e�!�����k�{����U������4K�4�vZm3��xDT����9���HHA���]VD�t+�8�!{�y����z�NE}���&r��r����Q
̮�JL��T�sR(��&y$E�*#��'9��
̣�Q���l+����Ys>���eakJ"*�+�XDBj�T+ԯ2��XT�$���K�V���TD^� ��"��٬e��$��-v�L�J{4s`r#8�	^���u�f��2�b����[׹s�C&WL���"))fb��q8��"�I���T�(�1)/ɏ�������_C�d�_�r��?�D!���he[�B�c΃*���ͽ�w���#��'��ʘ�B��莿CK�'��=�����3�{z�59�)��)g#�����"c�Z��Ӳ&,57�
Q�Ռ��qכ�tf�(wG�X^&���S���N�������{ H��S�/q�O8��P�ּ��սP�{�C��UB�L�#�p/\O�Z��T뻣�f����X�O\��f�jӵ���f]�j"��d�O�QˬacT,z� ����W"v�*�{�k6u�W��>�f3��ٹ�c��1���+�}!tJUV#������)�8L&I�lR~��h^�m��q4�<�Lm�w�|��<�G�#��Ǐ��w�٩\ˋb�cj����4Z��ݭ336�4�8�m�4���^J����e�G}��-A����}+�{W#����N<|L��ǽ�*���w�f�yȥ<��\Qx���4S���uM�Ej�~E+(��A�s1pzse��W�/,�w�y1�C��,,�&)��EJ�X��^JV�_�	��uJ��`��P%z~�ǵn^�۵��v��I8�!�SC0�r+W�r�[Cvq�]�we��6)�eJ���H��T\<wGn-�̥|w�qi���m�XP\=�V�rt_��u՞��Ҟ���更3ʼ�Wcv&�&�S2rE��r=�w" a:��
K�P�A�?�>��믾�JC�~).t�a�5��F9�x������U�,��-�˽ZE4|V��"���̺I��[�3��)�y�9�	>�.Z�3����ݜl]��J\m�oT'�Gs���.*��&qŪ�H*��������L	� ��f����*(��l��uX�	I��4�jy�r��w�71u9ۑ�����L�;��夃�qBސ��D� ,���}��Vӭ'=,H6�wǗ��/E*����uh0�a��1k'�x����G������B8�1�"F���{$m-BBQ/�ǃw�h��R����⻐�6ߩ�uII�ė�4"=�w�Bԟ\�� �v`�p�焹����^�qw.}����8�`�LqD��5��&��G=�s|�c4Q���W���O�֨/f�=��m�RQ�.=7,��7_c�Hⷵ�_��L�\�?36{��E~�3�1P=������ʛ�Oߒ?YBy��HM������÷�Q幥�I�0'�=��\J�Ia��|d�|hBL��7�ٰ�ۭ�3�v�l�LXh-��#y�Rދ��޸Wkl\`�C����+P��f�/� �(�k������O�1P�c:=��n�8j�P�{-c�*n�fս�U���S�t+Aӫ�:1�a�y8�U��ך����Ꙉ����������{Jw�8xԡ�I���#4ǰͷ�A+wg�e���s�w�R�j��eX�8땹RlN���Wݚ����E����,%T�9��m��������|�RVs�ݻԵu�҉k63>�^j�έ�4^�Pz8�/a�Jr�ʩM݁%x�~�y�=7C�!8����;m����:�<.��B:zX�;_��s:$-�z���yR������ uC�?&������pb@��]q[ ��Ȉ�Xc�Ź�ė>�T7�����W'��	}P�!��h�e��%�RuL;^��>7\G����t
�C�Ti��_��U��F�f7�>���&�������B{!%	��t���ǥ��Nl��!H��}J�Lԩ8k٨�o��v=ɒTِ�{7ek$�x�`]%�(,�;T���j �����A��"zB�-�)������r�w�=�z�Z?1��mK�1~�gހ���/[�{��>U�V8����i�M��NɣU|�{�[!�zzA�/r����F���,�Wѳ���H�0�<�B��Y�"���7p��ՃKxM&⺽�-9���xG���tg��Nz���g��Y���3f���:�(Ί�M'���]�&͹�Hj��I�~
˜�e�fN��FJA]f)��[�H�R���M�̡o�]�N�][z�l���x`ޔw���~���}��5��7�h�M�@��g�xк���]B7չB���Q=���'��#E��>�u��eu�њ���wG�B����)a���~� ǚ�"z9���=w3���&7�{ȍ�����n���D�3�r��H�#{��T;Қ���(hF�hQ��>U5mn�Ց��EM��2�o]�fz�wT� L7=�2Y��sM��\�j�F�T��WЮԅ�G�EȢ�2b���w�����gWi����4���x�<dS�<oϮ��w6k=�JC�"�����n����݉ڦ3�n%�b#�ݺ��5��}��ltĜr^S�s�QMw���T9͝��j�4�U�\	��o4U�zُ�����	Δrփ[Ѭ8?)EŹ�G_�,��R+H��{1H�� `������a����Ѝ��Md@ɏ��E���&>�N�w[�;���?5!��p�u�MU�C{t�j	P|����t ��7�E����z��:2���-�Q�m�`���b�<��-��ơ�إ����bx�.�1��Q���Ԕ��2��@���k{��i]F��0�+2ȃr�+��"�7c� B�/�i�խ��T�ȴ*�=O9;�W�ب�O�ʱm�	S�Qzأ�4�x,���5�Ssy�����V��k�wq]A:䜝���*V��o�N �tN���b�>�H��5�&��e��2.,<N�o~ }���Ɍ�ւ�����z�-�Ѳ��9r��ϣ���G��D�t6�q,��"T���*/g5i�םᛇ��F���}ױO\��ƅ�*����	�G�}5��i����_H��-�j�KeMZ�"S�h���V�ƕ'`���ی�ʚ��#��`֧��ܺ��t�{&X�a�9s�w3�]-�ͧ`�Lr ل��Ȼ�y��j�X�g�hj�� �;c�+����Q�����97�z�.����V�K:�P(	�Eb��J��yտ��YQ�MD������Z�5F�CI'MT�y�X�Q|�t�m�K4�(��T��@(��@�K�"~��i�����ڕ�:���ͱ�`]nzjŬ!#�q-k��ß��)'{q0����=���V��~��쑡	��<���Hx��e��a���Лp���"M�ư���yBlr'�~[��M0��{@�/b��UDut�Q��Y�X����naP�^S�%�(�*��q�IL��?�>��`�~6}Z�����C�>�K���)����;혖l�&{W �>��<�ߴWJ�&9�~s�2�.{����x�v㼭X.�l�T�T�U�[iV����-K(���V���+CZ���x� ��Wa����]��Ŕ.�jlf�D&�4��S.��������w`�R�J�bǲ�f�lee��fe9R��UCf"gn2;�C��%�2��5s�kྭ�Rwm�N�"=�-��P5���ڝ`Z�z��Y�x`�] ��{S\j/�e)��	�qB��Z̡���=�;�l
�D�9V��\������,�Sj�؞ͭ���	>��^Ne��^���ퟩ��g�T��V�7�ADY�	�����g��>�dl�Ɓ�O�qH��T�S	�5)��x�Jdp?O6�R�⒰�/���F�0��<��m�2��r��V��R6�?H����B�_�i�x�c�ӤM�>+2)��RQ�u���j)�4����3���G�{���N�P͝j��uY[�غ;G�:��oa{;ٳQ�C�=�1��d��( � �	�j�3�}�
(�u�����P�0�r:ޚK�nc�Aw�ݢ7U��n0ǫ�ڣ��}+��@��1@[���ȑa�צ�i�'��Ƨ�YO2��Wͭv�; n,��эo�y�t�]BQ�@�后(	�(VU�W�lo�njf������JH`V_z�}D��V���Wr&�~�k��%%^�h�46<���=,&[KS��ͣ�_��ˤ�y�+����3���2���W+��oP�טi߹�^P-n�v�*+��2��yqۥ�0f]⅍���)�Y�����/a���R��,F	�on�*2Gʊ{�nU�Ϋ��œY�v�o}���� �nj6q-�C�SڅM\�^�q���V�sK�I�x5	$��(ͳ�z4#�\S�k^d�AYoF����a�#�����qg�s3*��G�_s�V�"n�b�)͓��*�S���{�R	���"'뺘1�sEjiY�Ԡ�3�=U���_1,¤��j�M�n�k���Q�DbM-���Q{��O���qd�_
�~Sh�F�����w�_��|,w�@���2p��i�H��/"����.�����]Ьn҅#��z�z �D�j���n%G���;<�{g+���/ݐ9tĖ�&;�d����8��(7�z�:��+'�#;��T'�ɝ��vН�Sg=��"�dK��`?D��]�ܶՙ���G��ݚ[��E���B��f����Q��R�,;����R��>C�u:)��R~k]���>o[s���ޱ=����է�I�����$��mf�vi�S������W'�8蘑�e���=��Ҏ?-_�^Axm�x����I�"Ti"!��
�99n���;�|'{���3dI���W�5"�r5n�Ɋ:�F^�u��ei4"�{F�csR���v��V�窏�G���T'���B��&���6���V�m��)�fX��#�3Cj�'�d���&�ᒦX����al@\�����	1��b�_hؖ;7�����&/s�Mb�j[��5(,V��Z��.�C`1퐠`0� ��U*u3�ػ5uLݎ��FT(�n�t�ǆ��~�s���[<�tr�P�	�֠H�v40nc1[>�<h>�<��uh�?n��HK�%�'�ө�:���MH��da���j�wO�l�t�����H&���Wms�r;M���(������VGX�H�U�~#c�GP��g�cJ~�N)�)2;��6�,z�sk"�P"��ݑ5�l���0dO\�/�x��˺�۽����[z/��2����LZ�{�����p�FT�P�,2�����G5Bj,�������,,���}�r:�;�;z���;gAu�$�8��^�����)c�q�>@���%=�77Y2a9Yٱ���" �b���U�,��͏�\ѿyJPx��$T��T+�!s�귗��s����;-���CN *A�z�o,u�Nl���<Qf�7uG��٧�iᩃb�[61�i�e3��9CZ�cr:��@(	�M��ltĜ{�1I�|���[�G(77k�3'�T+ޒ�{��KRc"�^?�Ӽ�o&&�e9�[�b���δ�E]�T����)��L��͔�D��[H`FB��>�+�׺/N�KA �C^��um��^��k7��\,-�Su��w>�x�v�:3�w.7$��|7���ȭ77�_�3n��"�b��߂Z�#����C5��d�t��vW@4�Mr �پ
/��rP]m�G���E�ˆƷ���I,s�	6��l�ܪg�)�Ǡ��|���.���#n,r����s��(c���=��+�('M��|.�o��>�ON��gU�-�ҩ��bk�'�g�Gz�F�}�]���&����{Q#�Q;��L#H,%r��ޅ=GR�?t�{%x���n���hCe�;;n j͎nǆm�Zf-!�b;�L��U]Њ��@
�"��
�u��'�s�4���!�OD�Ӟ�/!�a�na�^��I��X��G��Zz�u��2�c�ʍ�:r�6L�6�0e��9��L@Vg���] 6������
�Y& �������~���� �
��l2��w��R,\�n�e��,9��۵��5��ӜkN�C�&�}ʝs��x}�b�ABA��~�����h�7M��P�x�f��Ѭl�V�eHƓ�ɑ;�F!��ϺN[v�m�m��5f\ޔh��9��̨8�1:�{iwN���\)����f�91�%�Ϟ�}M�4fNX�Z.e�C!�ed\�A
4�D���}����\7oaC��~��̗��SqHg!@�]�#�Vi�JT�GTt\TM��imT��̝���"m]{p��P��s�B/ߊ���~��������m�53�!���.�L#��'�/MH�Oӵ2Meg7�0��E-��h�h��%�9�S��L�����}n�h�2N9������"�;]�n��Xd֩T�i��'�^VB#�v����M�Ѹ�*����6�0�ɿP}��+U䕺9^�w�қ�St\�+�;Uv#v�/Զd9M� ��"a�Oo4�|�NL���5$Ϙ�&�t�.�z�ͯ��ڋ�=��z��q>�Ò���q=Q=���9H�0:Ӵ�J��U����w'܎*��lwr��c՘�}�Z�Y�g��s��G�{vz�G]��+U��c�����q��w�5��=CƷ|J|:ĀZ5B�K��'� ��TJQ�k�=����j�mj/��ƻtv{�p_i��E�fEH�%���ޤOr���9iVK��"I�|2y��j�y���!�+�5X�dq�C���ژ����O�f��*��,�f�JSx�fM�BqXH}��<�6�E��ݢ�0F�/���+j�ΝѠ�e� y�F��ZO�-�����D35��ۤ #+LT�df��M���4�e�s���&63,ɪ�@E�*�HD�)�P��U�q��p���(fp���!�YoP:����ݓi]3c�m5u�@������-ԑ��RK���*f�0x���G��Y�o!�+2=�D���WN���rU��C���mn�F*�8�Vou����j:�O)u���˶�,Y�WiVJ�6��J�l�{�N.şgn�q���(dP1Dl�����K�3���wd��[���W����[/��o���o�E:QRl�p�t��&�+���6NR�+^�����3�ۂ%8��Z�E�� \3s�*�G�a��1e�cd��*��n��� ��;2�>]��`�ǜ��[�f��3Q�L����'{	ľ�����XG}���T��� ��}kE%�5��/�
qˑ�pU���zi��J�)�fLd֩[���ճv��%*�4��u0��TuM�vo�n�9�CG�A3\��D�t���V�7��F���
�f��
�D���c6�H��Kn��l.Uel�ln������1Ү	�ڴX�= �V	}qd����#�S��
y����MX�X��ĭW%��R��o5ct-	i)�Tg����&T����3�#��
c��&$RZ�T��WQ#n쪀<��Q�*Ń"�h�B�e�\����z|��T�j��E��ߙ+&x���T�gm�̰�*f��&�w:t-�]��K��mÐ=A�-_|��!�4�����PGݵ�=��4v���{:K�5$WT$vn��cЪi�����fئl��E���dMk�-��u��|)����ߛ�����������S}m�x�>X%�;�;��kkU4��u�u=y���̉���'܌`n˴�>�,��-j={�zT�݇�8�@wC뙅��˽��������*�,z��Q��5�p�)0�Y���׵����o	�mS�"շ�X$�kr�j��s7��Mm;ț�����CNj��=\�x޽I�ېu%f��e�ΦMJt6X0A[OF���X�ڭ=*��'G�3~��gc6lRKZS�7��-2�ȆP�.�fӡo:�q�\�m˸��}->�%1��-��m��iD&#@�d���6H�����ͨqp�B�j�v�k�7kB�+����Y��{�7���P�Ou�8�&tb���p /D'sP�:w�ݫn��[�Y�`>΀�+3%1��t�l�y�Qu��4J��P�sN��*t��5��Y���<4݀\a��b-3n-�y�%
��VS]�
�2�Z&(�C�h�drL�mş ]�Ы����ڝ*��;���"���"���D��$\�n�߷}�w����Jar�"�2���Tb]�rZ�D�B�Ĥ��G ���[���}�w��HUf>��B��%S ��D"L��S(�Ȃ#�$��� �2C�:���j��gdUE�ʪ*��"�("�"
#����r##D��h�	+�T#**u��A�纚��Q�B��*"�0�۞eIЈ2B#$�"+�EQ��J�r���TYԇ��(��V*Y�Ir�Dt��Qz;�QL�UJ{�9���jPN]G�Q�E���ʹ���v�Ƞ��A �.D�J5�.�һ.Qr{�AE̋%B�{�dEU���T�_7D�G*��.2*e��'+�9O�9EL��I�@����	4��j��o�켗Y/l'�{i(��x��̪�j��Ib�2t�d�	�a��au�܃��{C^f��������g�����}�t�n>�k�X-�}G�2�ۓ�ϥ{*�~�%^-lfi����K4�����ϣ�'�[��`8�Š6%06��&�`ф�w���I���l��b۷�rp{�Ϗ��C��o��#��&{/)�0e�;�{��1�|0/���>������X�#V����lsMؖǺ��L�m=���)�R"oU{Of&��ד���,@�I���1�î�jx|�ʽ���4�GC�2ʘ§�6n��Fe=f�R
��u�m�(���m��2I�h��GKa�猀�T��f���S��'�J�׳�E5>����5.�oK]����Wjjr��i'm�M�wnU/}G��49�E��خ'g&v��3���L4�PJUjN՛[@�ʯ-�z�[�w�&����(�#Md/3wk{r����D�g69\a%IJՊsFY�V�f=y�V�߻k�����n������ ���r�c!QB�Y�JPK`���w�����+ lgqf��'mgG�wRXe�Y��ƥ��~z���������i�m3��+מ�u��ۺA���x{ $n�mEs�}���}Ҧ���sέ�׻�4\�Tx�m<JDQ]��!�N�8c>o@^�2�=����lP�,C+�z-��v���y����)>["����3t�V��L���c�پQ����e�q�1�����{/b�5.�=���;����ޤ�':��0-�7��Zs=��˾�F�y��mPN����̸8Fl�1<v��ݢ��|y��ge���H���Moz��D�����cۃ��ol�'z���w,��Ц�����������]C��:Xf�ܞ�2K�Xť3����V��I�5ċb}��!��x�j�9	�s*�{:e��l��opd�>���VA=����>�:L�=tGsM�R����x�ӏ��|�j�3�A�6,�-���Q�'�ґ�p2�ll���mn���"{wO��e��q�N��
�.�'�f ��8<��g U��(����u�����gˤ�ܨ��T6�&y��]��N�q�fe o��Y��S��xWvv�״8�����#	�2�{����z"}=�V��2���T���w�zN�ҫ/�)�O:	�FJt���Y��jL������el�I�����EÂh@)��T��s�:��(po�5���4�3w�!G����z�-�� PF�����FN�ϸ�C�d�j�de����>x�fj/�m���CN;�|�.7:V��Wl��q�4P�rC$%S��լ�j<�}Mf@{��3Rʈ��Y�ݨ>\֗�G$���T3�e_ U�9�\�����X����}oa�x���f��d7\6U���=kL�铖=��َ=eV�l��1sR��8X��&�L��h����"oj@e���$���6�i�?j`�����'%�D��z�ëE��g=}B�o�ûYN�r������t�\�k���x3K��&>��{���'��Ζ�O_��ݰ�o\Ӎ���}0�Lpκ�x�F�1җ��l8)L֙� �5�n�}ѽ'x���V9�
5���!�t.*/�<�	����T��MzMn!��m~�~�u����X��r�B[;�	�{f��b/b�� '3O��Z
���AF#�li��EV��U�{�tL�sbj�J�Kơ?+'��٨��;!i���^�C{Gff��L[�7��9�;��[:�6���9�z0r���K{a�-b�"n�Jn7�7��t.%�� ��h_4׼����k1���̋r<��C�V�#�����|����8ֲ^>E�K"��(�� �-�ӣmR��9C@�{fȁ�6��odt�kڃ&|;h1�j����b.���s�:ي���p�`��"H�x6�?}��^���o���l2�p�<xL��@E��*�lə�#Hn�l�:�vv!���-5?�>�k�����G6���xn	Hn�=�����l[ᗓ�>E��Cg܅������\o�M;�ݫ>�&��מ��D�t�M��é���@܂xd�S�1�2mz�sfA���ne]﵁=�J��d�X�4�j�OSD�n-K1�JN�q|��3X���_K�|�&N�|�5�viDճ��7CU"�M�u{b��j�fm�r�tۿt���ܯ/Lv�Y[{afL�岛�FC]��m�6Y�2�W�bs*��wn'����0x&�G�{m*���c��9���3dMɻqӏM&_o�O[�bU9��[ԧ���䀲=ˬ�GEb4�к9��.�K�����`��Q����x�9��{��S�4]�[��'Te�3cp�3!Ê������[�%^��B��˽�Щj����6S�YjeIխۏb6	f"oo�]�g[v>t~�N%���k\�5�0���N풺i� ���l�FJ���vF�u��e�n9�.��o��K�0�j̹���� �5>�<��*��u���6�H�۶��޴�`���Ju9D��t�<F���!wA�ow3z�n��-�F�l� 7oL>��jO@����b�b'~>�[buhӛ��J�(��OO�<5n�}���ih����B�2I��[/9�g��R�[����Zb:n{������8�ŧ���[�*�b�=6#���;���V�i�#�dtv"n���}L��ӥ��q���'�{�}:���kwL;��qM�07�?n-e����Z�A1	�sڱW���ƫ�M�r_<xD�4&�Uѻ��� dJ�H�����ѓ��.p�������v�g�hȌ*}f��2�4�Tf^���s(��{���GKm�*з8�T {�LwC���g�[4��nS��ݩij�gt�1~+��L�u�ڽg'/�u�M�jKܗ��+X�3m���,�El
��ܜK&�V�wfS�6YΚ�(p��ԍ9
gY�]�!��۶���z[���*�>Jrb�n��7)z�Rs-un��,n�r�5�ee���Y�=�y�T��5�h�b��*��g�:�y�<2�r�=�@�Z��,��fU���e��\�c�h�ؤ�9ݘ�%z;[$5�]��#��%�Q�+��l�7i+���*�|e�oF!�1a�u�����f��%ۄ=q������~������3ܖ�ĝeF���޽����v�U�kd[_��/�giv�8��+������)�^���ta�Ȕ�����&[��;�v[q�z�߶ӕX��:�u�fg����n��=��{n6�1���%� �"t��\�Ԗ�ؘ��Y�X�_ZOu�����Z�U�{�~k`1&�͕�����,���b��d@��گE$�/fr�������VNk܎��!��c>���ضy�5f6g�~_j�ǉU�U���UrX�D<�Ѱ�a{)V[���/Y]�@���"o�'M�"ѺU��`�(Zn���W�����1�RG6T�ǹLb�ԟpU��:��Gz��B�0��%��l�nt6,wn�������X��w���0��_�r��|��r��u��{q��>���1��TVjI��5��3W�Օa��� �c�cp��E�1����7����ʅK��Xݘ1�s�M���5�����Y��|�+3�T��+�מAm=$vT.�l�첼��9����(w�3!t�# �*�j�B*bl��ķ^�|����}y#{CX�v���5����B��lЍ2��N�}��`�Ъ򈚙��`�we����9�����6PO�!�LU��R���t���^g<��D(���C&[ae�+�NM΅�/�*�jN�J�(�L����6e�;;rﯺm��v/S�Ė�Ty-S�Ꙟ�����{<� ��{���PP�m������Z�n�V�V�41�Mw�6��KrE6E�̊���7m�������^&�u�4������1���|N���`W=>���t��M0�ڟFMX��%dv;.%eˈ/�w"@�5�SŔ�r�НmSŕ�XB�b�q۩ܠ�V�e��p���M8^X����R�J�t��.���A�MB��Ũ�Z��$Χ}5ϳ�8SX+\v1�X��`1,���H՗l"��O5��,\k�ƾ�ok�=���"�̥n��H���F��l�g�0�PV�}�1�/";[��I�a�]�H���6�D�S���={ag�s�b�V�ɾ�5�,���~\%.q؜����<��{����� n�*Wq��Q�B�-�h��d䰕aM����8DܳI��C��S��#���WFl��"��Y�dݹEw5�\�x�$��g�}Ys��x���a|i��Ð���/س��-�7gE����WK����`�%!����7��VH��:�Һ��'3vC�]��c���}�Gr��8�z�d1���!��}|������o��l�Pmݽ��lWGZ�ⷰt�+hW���b�0�/�/a�=W�\^Mm~�zǾ�?��W�տ$ס�7O��� L�ນS��E1���� ZI��ֻ���~|�����;Mw)y�@��I:T��)�M�'��}�ɗkM�����>���������&�����!t�h{��KM�vV���7��Y���T��.�|S'`Ηe5eXm:�יK�;����������sv� �4�*�Gd��0辛�:v�͵�ʖN�[�s``^y#'�;�fc~�����Om���}%���O�٫�ꉻ���Id۔���崞Z;�"!�'�`��J��ӏ����σ��K�ǘ�H*B*&�:4\�[f���<Q�s~���wf�v�����VeW��+���5֛l�)�f\7I%�LS>�Y;F�u	$鑑�f�A��"oثdR��m���٘p�U��O�.ϸ d�ͅ�ǲ���@�ׂ'y?(���du�ZYҺ�Ƴj��ݕZ�ټ�"���n�
�	�k��}��^�67��iq��]o���Ř�l񑆤��Y�s~���^�nl�f����/�#��GG��EP�=:V"�Ot��i��l��בK�ya^kn�������y�z��(Ԟ��ƚ����p��\�gV�}�Gķ�W�GL�Bۧ�>އ�����Ա�TO�Α(�ǲ�,�vŕC�.�H�+ٌѓ��nkǘ1����W���8R����I9Z�/'�؏!W��gr�g�&aU�7U��
D��sY!ٖ���,X�.����s�r;Yiit[��ߨb<�N��c�F]�ԭ��"� oB��క�T�L���Z���ڽ�=��dX�G�ǭT�$o_%q��1�oaZAE$��V��
NϹ��߉�i'�&�n��>��͠ ��3��[��fV�?���3��s=��q���4�=�}�d!XDSG7n��g�^��b����*/¡����O�ݕ�t�O=�1�'# z���{yB�����׺$i7m2��ڙ�ɟF>��t.�fK�Ȥ��ګZ��4wTV�̄I$���l�z�H�>�x�d���DoQ�Ǆ�."	��-�����	����襉+�C��V[<{e�Ϟ�r�h֚y��!���dYv'{�L6&��.0��,�Z�=c-l��U��l�V؝�UK�1W|��o���א�J�d���؎4	���4��/(�_��=jO��v /��u��FU!��m5ȄWW��p��\9Τ9R��Q�=u����V�װr�)��L۫�r��m���;�wg��WB�1n��W�Ů�X�ÔohJ�7)P�'K�T���
�4�ZӫM٨����c�2�qI:u���/��!uA�T�v9k:�Bfګ�+V9`,�O|����īx,m���y����R�}̲���<��cR����8��]��To���%� ��
b;e�m.C���u�-���b�h���
����Z�<#�����)�txBf���EJ���yǆ�����7N�~��6��,��ͧ��Uq�l��L��i%��`wK���b��(�۬��
�r�
�Y�5��0a�Pc��(��Xt�v;U��^�Ob����a0��Ԭ�����vSH���ӊAi���V�S;N��}եH��٩�ڔ���*]!.�Apv�k���-�%*5�����C��s8w �r��-5S�˻���D�WLL�-�̻��}-U�S^�M��gd�N�l�n����l��]���:�Ƥ��	C:��t=��ζ
JR�nq���W�$�>��"u���].�����7�VK��dN�i�Y*n�[�;�L�ͽ	�&Ů�A���,���b�aҥhf�U���L{�L'�����v�˘)�Wr�����r5�Gw�������6l�y�c����/mgfǲR�c������ZV)1�*�y��F��i��@��h,)���r���`��I"pʟh��S/�waR�Nqi,Й���eج�@�No�ӽ�x,���p)�9+8����Jk����t,�[U��͍fa��>҉�i���{��N(^��m��A`[¸�����j�h�-��֫iid���yA��M+�N�$�c[$�V~� ���Zh����D�V��9m��\�p1��sP]-�7���(2�s,�\�lcS�%Jm4��넝���M�H����5[���L�\$��E�kb.����ygs��^�f�:�ّ���l�T��U*&���{���4wSw]�.�oh�l)���̰�TF���n55'�0MY..����t�{�t��yC�rCr00�Y�\N�O��1\׮S��.{�٫�N��7\@r]u�*��v��j�hvo5G$�r�iUyRμ�s`.��q�b��[P�)�ˣ%ނ!����WwM�y�8���m즳�8�շ_ëÌ3�q��^~I�J��WV�'E���uJ=.���4��OW1�ùC	Z�M�� �}�p���y��n,�U�� c1'��:�nҳ��4K5	�&�
��"���jB����Es5���;��u׏S���r�ԤuN"g�d%�IG^K֜�rwW`�b��Q�0j��rV$�3��ݘ��xE��,�q���us5=J�h@��C�Ej��t���:<j8��]y]d=p8�U�C
����꽸�s!/j��_kN�&��������q|�WĂ>�� '�~�+ED�GNr �ΕG
��{�QTQE�^z���߻}�7ݐ~R��E�"+�e��I,�ֲ�D�L��WR�r �R��w��}�s�L�_�9��E]��$��*�����*��U.TG+�f�ed�9�&l*�R ��"�P�12<��q*]��N�QQ������=�p��ª�R"�#
�u
�̹E��4�$�F�NR�Ԣ��O{�_^NsR4�v99��w<���m��tE̢)��eW*���G.V��87w
�Yr��ÑV����wx"e�%��#8RԢ*�(�Qy�'���R�=s�3���Z�*�O2B�$��p�ݹ9#��*ʢ����}1�ۆ��	Z.�"p�T�ȃS�Nj9��=�nb7R�tx둜�r�H]�X|��N���u�,���ERaĜ2r~��BP%	f�
�vI���.�����ʴ�h�E�����+gW#h㙜�7S��fG$A-V�Z�!yݹ�wʕ���u�3�0Mh�eM���>d
Onh�U��qr>��w��{��w�[+c�gf�c����1��`�t��uB&Cuhk.�t� fJ�jq���
4ሃ���kw��2��)�-�l�������s�0�����@<���,�(ݬ�]3�O�D�����bM��^K�߀p��>�l�HX&c�uMyq��v��w�g�ʄ��F�gf��Ry$Β)�4+h�B�T��gm��{h���-A�/�s�+_N���`��9�5-�c�3��Mi��տ���*�\��L��>�gض;#��M����=]yt��vv�D�:�����c!�|69��,��lƾu����V���ւN��������n��OsX�� ��9�X�N7�5��̀{��0+wW��8P��>���ݧ��4�!^l��i����|��ׂ٪t�b�+��w/�o�n���ܠȢ�yZH�Oq��H�W�b~�H:�*Z�%7���"E�7�}������aL=��Q"��)^+RFy�WG�l
��ڳ�횹t<��w�<:�"�F���R�kݷ��Uت}|�pN7�kT�#���II:�fLJN����g����d�[��Xx`ޔw��A��/�z���2ԧ�r����5+�~C��d%rb�~��f|�� ]i�<�vv�Wz{�w/���P��z�Uy�N���d\��5yv���e�X���SGĪ�G2�9X�t����}Bh���o-Kn'�L2��Ԩ�o__3���N��Y Q��ݹ̝l�r��AK����B�5�r���c2���$�R���%u�{'��׷����	+A��Z�F����GM+�6]�o�ŷ�q�Iu��ڍg�k1�P�z�1���\w����ff��/�o+Mf��F'����a0nR+w�]b�	�6�E��*����ݔ1��f[�p�7�:F}:�P�Em����;
����D]a��2~��X��w͙��OG���%���F�W?L�1�ԿU��'��m�W�-/�!O%'��{����à�mĎ��h��~��K0E��ⶄ��Be�)*y��*/�ܔ�R>H��3(�0!޿��m��׆+�.:�Q�~��|A�.Q���C+=���=��������
������0Y��u>�e2�B��S6Q�w�I΋53�Q��9��Bk\�d'b/^�ۡ�G!T�'�h���x��e�n�9�l�c!��Z|�{��r˟,`M�{���
�/T�n�_p��a2-�[�
��NwΌ��jw�߯ϱ�ư�J��M~���8��_�؂�S[�&��׳[[;9z2�F&�g��=�>���;��9C��Z��$c��a�-f���^c��5�6��٣ǩ�t5�s����RC�N��~���D��Y^.������ĭ{s�S���S�*>�9 ��|ɩ,�-9抋i׶j�Q��P���t�_���Q��+��9���Hwif��.�ʚLB��Z4���ܤ[��cpnz��)ЎX�7�_W���y�i��5�Ϫ �32�x��~�~�O�q��=�E��y0��1���zV풺������W+A��y֜��9}��3�%���u��.���J��U���ZcY�Dϴ��h�`�"ʴU���K7��H_L'_@v���b6��7�&V���������� �<Rk�9�N�`*�hJ\nX�9�k�U�+f�ٗO�`3\����v���9#�ňN���e�*�X��	rAS���&=���P�#ͳ��~f9@F������K�hxkjOcz�3�O^?Q���)�w~9?v�؀^l�Y%�cr)M]?t�¼�S>�\�w.V�/=�;�b|3�A;�,%�F�m��7����[ڎ[JJy�l����9��b2<6�yXue �=��c{�[B8ۚ�[b��cr�DD�B�'6j��I@7�sѰ�[iy��zZ����ջw��)��hkH���iŸe��H�lϢ����~��2����eE�� ����{����Q����k�W��b@��}�᯳o�Lq���6�M��m���F=��='~���nBQ�X�5�0�����uylU�T��87N���-����<���$l�����3�W��ρE�딼��T9����"ⰼn�?*��G��C�}�-��r�o�
�n����:�6	�������k�+�!)��"�h��ɯ6W�ݽ>�uJ#��
ZQ�'��G�7���C�J�9N�H�IyӪB��]�L n�7=Z��sW�:�\�7��a8��9�	���^'�'��Vh���oon�?��(��&M�h���N�y��-l�S�ф��4�ۥv�9y��_�no�m���Q(�@�N�r�k�np�t,�PR(9@���fL��u�X�p�霹��k����KH��C�2���Z-_��w㠙K���=jq��Y;0*�E�e7줊�v�m��,�>�}|��p�:�e;]�4���ڟw&��Y"�=y[ُ>�7>w�r��Y"�@��^�ƪj�N��
������bOPd�%� ��@B.e��G�ř��R��-cV�ʁX��O�i>�S�L<�+�2�5�|�U?h#��ݏ2�7K�v���v�<=���I ���9-8�L�~{����j�>�f�MY�z�9�ȗ-W��k�^L�4�h����#`ׁM$��f_W?r�h�Ξ�ᵂ�� ��z��r�BL5�u���ߚ�O�ޚ�w&�����;;��1�G��9�w��^c�1�Ȁ�ݜ�Yط]���������n������ۗJ�IU�0��E햜�I�*��{F,-��J;��N2�,A8}3*������ήi���;q]Ć곅'��R
r�0����Sr���5{V龉��˫�emj˼.�GL��#�D�Gל釻��Kad9!��t�R6:B�������;4:z���U��x] ;;'�dl�9�5�F�T����ls��J0J��d�W�ue�nB�Ve����}�X�F���fFYp�fDZ�D-6���=���2�~��DO�De�G���P�*:}��\O0����_M��/��,�k�zpzd;�=j���@���]_!ʀ�'rbޝ�n[i��NM�͘m������yXϟ��A����5�����׳.���u�t|����&�2+H�U�
̪+[-���>��h����'��P8��"D^>gS��䂍�L�H����MZ���v��!�k�CDF8�	�uY���氭"�?��p�o�ܑ6�ݴ�WU����w��zC��{P yJ3w}��X^r�4j��|�|��q,��Ѹ��~�5��z"B�Y��tc�/i'�Ve��p�:<-)B�:��c�Jt�qM͒,�Wu�+b��u�7��*l�o.PG�(�<yzo{*�ƈ��Tnb�]��Ag�wq#��V7(e%س�V�ھ�k��tf��-�yړ3/����b�3���v��a��ʓ{_!�����S_����t��>�ݴ�=ۤ�����bn0�ɼf;�&�c��3D��D�������6`�LA��_��M�^M|z�lVfҹ�|��O]ܨ��E��G�?X�6���#��C!��Cǡ�"�4ڰ�;}��yD�Y���Q֕1�j��6�&a�qB._�9���3��}�Q�/�xz��wi��2�c��m���V��3E�x��&����B�"{��F2ё�u��ﰵ�D�O*u��U��e�i�Wf�tsn/=�f;֯�7ʆqwe�n�:�R>���/]��u�k[�yD��y��흠��߶���]W�������8��{}�M�3X���yH�S�݌�	����X�U!�L�'�3�7���A�ܛ}���=i���{�ρ��NO���qU���� ���"���vzh��	����ѥ�A��Ȍt`�ؕ;��[��L=�	�Y}n��;52������"HE���;���Q�@P�=�J��W�z�����x"YG'S2#�C9�v���\�!�G��5:���jә�qTo�<<�~�����ܗqeuz�aUS`�S��]>k���A2���Lf�^h3Վ-���z�8��4�{�%.㊶}J��
�]6�+L}����eB��_yx��nz�q[ŤHט�'���`$�2�Z��������Wv�u�ʘ�ˎ�p]#qG��n�[�i��̔�f3��.r�����ݮ��:,�9tN�I��<ڸ��k�7*<�'�J�&�<�G��B����}ώc�s�J�@/6D,��:��g�k$�n���'U��^9�wmx���� +�ǡ&��R7h���	�w��������ۯ�H��V��k��vn{�9��r0m��-�5X�֤fRTc�n7W�>{c�A2��U��Dc������~��4�k�k�0�f| +3��7�?a������y%�iآ��Q*�tm_x��q��r�/��N��v�WA�ӏϦ
x�s��g���LxS��P�Sf四살d���m3��)^��Z�����օ9�tTU��ƫ2S�9��\�=�\�7��E�\�u6���l-|���1�5�N�8��1&bq@5����.�G�v�{� ��bʟX��f�+t�aA��MN��3Mg����p�i4������^�[�����^�!"����CYp�ۇ���1r�!�9����K+&���\�\
���;UAe��EGC5}�,-iQ9�)b��m��3��p㙴Y/p������ѳ\ʩNr�3q�t,�PS�Pr�6��Vemn����"u��~̥�����U2��I�=iD�؎:#�⤭�w�����/G�����ܑA�n��<��_�n�FZ�9-�g\�%݆K˒�qc8s������s��Y'��J���ُ@��=G�s0�r+�)�d'Pz��;iyk�Z�;�\�H��g�{�ON~�xx��f�x�\�b�ƫ�\��[�^�u��s�<�g����z	Y���f�{����n�I�oe{_An������gX����.e����a[�u�8Q���vq�1���mt7����T�X!��,�j��	��7��х^V>ѧ�:��Ƞ�R;���.���*去)nϵ� ]�b<��J�9WV�ä��Tr��e
�7��H�����l�����r[�,zB��^of�l�Tݽ3���z�XǕ�jT&w_z{�+'XǍ*�}�-�fn�tM>�j�����~m6�Ǝg	�n�`k�9���
�V����՛�F�A-}~����{��,.�F`,3v�Uq��h\���^ɩ�}~�/���}s�����od\�a'Z����)zVpz<���'��dݯv�m�s�C�X���.E�6�E�����\ߦ���ƺ۾��Z��vM�G3!��,Wg�tK��	� �d:W-��Yz'$U��ppT�l�z&�r�:��a&���.�(�OW+�ov�[fƿoI{����|��l�cR�	��c��,�@��W$Iy���:o6�oow.���+)����{���~+�	���#�V5��|>b��u`-�Ø'v]�v�Q���F���=�:1���~��X�i�Ƒ�{��:ǰ8n�ܻ�qj�Kd�1̺QJ�fbY}�6���Z��D���vvYK+`�E�E�aT�!F���}�6�]	�':�Ĺ;솚]��GLt:��m���R�]ykOk;�ް;��"�at���SG)p���'�L��K���=y��uj��^H����m܍.(�����X��ٴ��7��T�yLJ�E�!���;��prlWgBM^�ST��|'!�y�,�.]n  �p�<6�sRwS�3���-]��V$�J�^Ҍ����h�Z˔�����{9M�׌�m��U���񪲶v��Ŝ����Nj�[=N�{�zl�d�T�Y��x+�O`X�MP�d��JQrd��Vv��\�vA鐝<��;�dX"��袝(��H��c*¶�Yy�V�.�����b6��ו��Tp�2���9�n-�����)�L�/#�G��.�v���M�{�\�mèP���v#j㠻�q�/��΄s�[c���Տ�OU{3\�Xle@����Q��׼�>*�M�[�L&�Р޷nq��^�j�λ{\��|��8\�gOgb�K��e�L*R_ 0�x�ʏ�״ �ū���:�
8�T�_���������V���v%b��M��s�;0�Զ��є\wY�u7OP���W/�]͍n���ZXP�lٱ��dPs3o�D*��lIX�fix!zC�r��T��r=���s	eY�1�G3�]�ǲ����_q���C��5�jٜ(3��Rޜ�6�z�	�8��h�2�X���m�X�|���hP5�}�2�F�$�|�
o��a�o!��)�Rھ�ˏ^��ҝu��*/�2�H��`�|:�b.�f�
;�tYF��r�rk��`�))Rm5���!��ʸ�n�lZ���̷�2)l�PKu2)b痂>kEV��XkGR�T`X�,Z� �ݏ;��a�F�a@��%3��iѕ{�CF�ԛX��QJܶs���*�6l��T�4��|cވ�).�Fec�ed���=��`�r�V�/Z*X�=��+��NMtTÒ��j2�7�a�)���LGf�S`h�t��(�ۗ(��+�ŵt�]AtnZ�����)V�z��u��9,^�d� �L�܈G�l�(�U8��/7�bc_
w�^�7'T(Mښ7�wՁּ�V�������� wJ;�&B�u.�JŃ���.sB�Q�9s_=j�}��r)�%5v���Ę�xUe�/5��}N_��Kw0�qu�gQ@ͽ�	t#���m:c�m�l��T՘�����-|�Yk5N׎>̢k�#Mt�.�,�9��n�Q�L�?��A�:���/ϖ�w���š�+�N|���Z��m��5�J}�r�-���#mnj@�1)��ٛ.I���q*πW�3%sr��>��8�sq )S��Ϧ��	�<��#������~��}�rS�WV��2���"#��	9$��Ҫ����Z�x�+%�-���JKt*�w��}�r�*��TUk�}CܶT�A�"��d*'u)��D*��Ԍ�����<�sxm�^z�9�h��t�y]
se�S@#�-�U��%���/WD}���qÅY>w�N�<�Ѕ��6G)w٤dD1��=����$��6GQ
/<q7EZt���n�QT%O%�����8���t��Aj�,����0�Vn���Qir����NbT�{����y�rr]��]>����ĥ��Q�ugԧ�n!䋬���|�v���O�og�� ����G/�1�A(p�JU��~1��9\��OA'%��kH/�ysΏYa���=٢2qOwws�(��NN��V:*!��3jաk��Ǟ"�+p��������E_w���rG�"_��˼����\NV����"��P��ʀaU	`�
�8B��7�]��vl��g^p�S�p�-){�#d���@�b�jM�,L�l���I��z�}; ���l�@b�i�`�޽��jq����r:�D�xM�$Ϙ���)�&�'�mmq�}@�T����&Cp^��Cr�v����@��6ȍԺ�ܒV�V�%u�GZ�j�,]D���Z���Xa�����ygr��d��ѷ��t.%�H�nL�&�4���I�����z�=�Tc46����C�tNz�`���a1 �$͐��cVa���qL՚r�F� �-�����6�!o4�����_M��H�[C�qCC��y���m�R��7�tNvM����m�41\�j�:2a��&�=r���b�fwe���ӱ�t�*c��y�;o0�j{��d�K���'���s�f��=`���-�MA�,xPsDm�NG]�sl�DҚ���ڬhM8�s:�wX���8�E���د#G�^�dV��6���M���ۙ�NT�v�'�;s�t9f &����B��f����^dh��g��E��K:������Y-�*��ԷQ^��I��m��}����m��Іd{jS][yj���]����{��j��E�H������9�~z�moovW����6����|�>faz�-�D+��^}�.��9�oFu�CrXަ�!�`��U��]{2����;�?����+��9��s�Mn��~�F�ky��h �a�܀�SY���/o##�Pΰ�P�h���h�nPO^=��N�����ʍ��P׹�ۓ��v}�>�;.�_��võ�5uێk}�%Ad��w�%wLr�f[���A�}�K�^dn�Y��y�ņ`�m�-�G:9@��_�X��k1��-.��&�"�(}���ޮ�� �*�̇��0V͑[ů{6Ί1��n�V��n�smM[W���Q%�{���8��H����h�+��Χ�H�$L͜�i�/�so�)̯�;s���0��+Iv����t�yO�!�^�"����V�9�a��\Q(߃����|u��HCzl�$f���Ԯ�h���/`�k�b�,w\E�F�:�E<t7���
[��^"X��/(�6A;w���:C��L�\¹_�mugo5Y5z�z�I��������r��Wڎ�T�6ƒc�T⿯�.���7*m��ޞ!��"���;�-=�ǌ�n���u�wi���$&U�]3y��wvg��"Q�F���U�	i�r�@Ѽ�_]�efCT�2k��})��qLGt�����qշ��{���}!R~����z�,vǝY����?[lg�� �i�P#o��|d�Zڬ��i'�
�:��u���;#!��k�u��g��;z���fH}�a�HXg�,�_��/���>7��Y)w��-��>�e�X#z��������<ȼ6}3eV��Ú&	p1#y�M\1�ㅶ�9;^68�k�)�Cl3�y��}������'b�_Sa����x�7�.��ى�V�2F�����%�$�k=�-�%oMx{2q���][q]�Tϫ�/$��ߦ�c�;��`������T~�]�f��b�;�ykI֎R�@�n0�t,�AD��D�،�N�	�f֎��̉s��Tx�<P݀Խr���k�N"��_wKz�*N��.�� �k�DVG��Er�e�<R�2�|�f��8Z%� 
��,/{���|����.���q�<-��^��W�c�/������3�=�D(u9����*ִ�v1}Ye:��:�FT56�Y�{�_lO��G)9��ʵ9�)�;"+���s��J��-T=��pq��)�n��D�z���V�Ӥ��W�4����J�F��Î7A��r���ě14�_��]��~�V��h��n\h2q%��)gT"�Cul����b{�������ˏd?F�w"���sx�׊��w�U�fg+�"źB�����[.�f�~R"�	�N�ᛵѣ��T�r�
3fF�.��^�C�M��S.�<f#Ril��y]��_W�L��]���|�w`���׊�H���������8.V���m��T�M7h���ۻ7D�}~<� A�&Cvx�}q�]���XQS�w�l����}�c�[�zGt�Kb0�rt��� ��@� �1Iג�/�>�w�0�����:�=��'\�W��V��,�^�:w�WS�Mkzf�R�o^R!��i�o3a�=jE�$?J�d|��P]��᫥�ևw[k�A��*�';6t�v�����}��eD2�ޥm�U6�1HI�M�G�ݣ޼cjL�x'�d̩xu��$���9w�����fD�/]`<e"���5���v��h�~�x����̗����>(���fJV̸�1{�e=��v�V�휮l�v^0R���17F��t��F�����5Dvb��<�.��4q�ݙ>&�H��u3�P�R�徛��J�{.�.p*��ORM��;t-"d�*��y]3ƦFC]ǃ��i\�|��6���ƣ�i㷻����z����0��fU��/��Bx�׮�\���
�5�$��^������Go��3y�6��ûY�#.v��mۋ��&�o�m��L��C��7J�nI+e+v�[�����J�4rf��Wi�z�.8n@4�B������z �Z�+b�P2���lESVp�{̬�tB��Ⱥ��zaO�����;�Ƿ�E�����m��mNm�n�����g�y0�l�ϣ\3�P�J���('�yL�玲�/��@/t��k�k��{�vc���
������ ��7���B�#�|��3�b�v���)bwD�1�^�8&&
�c=7�kj{��k��.���yˮdd�;M��7�c(SM5�n��7�v}����t�v��HW�t+�kP��>��?�C��s3����Lj�t���O���]>~'����i�F�=)S)�Xg	A6m5Vf�3mV���XEY4� �)�b���n�Y�l��iq��5Ѐ�'�����.)��<A��b�t^b=�wx�- c_�ީa0�;xj�6���/hl6�}�D+3|�?�ݗ�n�n5�5�e��ǚƆ���� Q� �=Lu6�|x��T>�n�>Q�I����-Ν�팍�D���zFiPsV3#-C���s�S��]7�4��R��¶��/wcfd�w�Py�I57XqU-�x�m�5R���+hDF���e�$��C_t�����9zR�$��� ����ʮ�\\�k]Ñt���R��+�r�6� ��C�mi��=΍�)co٤�^�"�
��8(�� �OA�T2�<��C�:��R8kL�G�R�ֳrY���m*˒Tܷ�ҁ[
�e1@�uϺ��O�[F��Ô�&��cN҉�VŃ\�^����&'�A�鳚��c{O{g2=�i�n���=ւ�s�����i-p���1�$��P���˷�o�1�6X	Dz�qw�Z���\�Ô��£�ۉ4Fv�n�Vw-���ݼ����R��8.�O�]9�`ʆ������[wu�d����[� k�t�I��s�[ $�ю6�g3|E�S���Nq�(��i=ֽ7t�z�[�
�J�wH�m��4;fe�c�T��u��\[���=����w^� ��6Rz�x�G^��KL�Bۤa��e�Fǅ�W{Q�Us}�|?�31���//��;�ܵe%�f�E�v�1���F�E��0��@lJD���nSϷmˮ̃��^_�X���4�T�f6�z�����N�@�g�<����ŝ��wF夎k��[=���'���{�	b�29�̇9�x����v�^*��ǘ�����Ԁ&��q@ד���X�����~�D�?*� ����C��SW?E?��H)�T)nO��Va���n�ڬ�P��Ѧ�+[�z�~�;%t�g#�/ �K	�E{h3��*����%���z���p̼����mԃk�f��*���fB��N�:�Ҏ�v��'���Wy.�p�xc��Ꮶ��>n=�N]�_wq|���1{��R�zYd5�$E�S;�'^]D.��~��9�Fg�sh�����%�U�j���Lϊn$���s��^��g���Z��x%��]�S@xgǡ]x�Nq���I�ǩ�S3��1�6�U!�2�m�(��G296Z�E,472z~EgW����m�4Vj6�R~>��9 ��A*�C)�O���O �ȾS]@�j&�r"��y�S<��]���]��ןq��{��x偛�!�ؚ��5�����f�´ݭ�a���Q�����˶F��:�;f�%�<�����6{��B�rhק�e�w9C��P�Zv�.q��q�jN�8�	3��.�[��6L;�ڬD�sU���YP���/gftU�=wj�y�}��3]�i٘�O����:�3�T�Ƕ7��Oߔ�s���j4+3�b�VZ�i>��3��-�&��ʶ-F{1���k�d��N,����_N����]Qpe��4�ٙSO3��c�b��qe��vo0P��R�>:���lD�����޴��I��nd�fu�B�:Vi#9Q�[U�3�l�64Џ�7)>�{���z�խc��݃y��3��jr��9��]e3Iʲ��݋W��#���޹s�&��vuz1�ȟ(z��L��n�߈!���9ۜ�j)�6�O�Q�7H�:����b��a�6&(c�Wٷ}ǶX�<nH�Q�ډ��X� �$�cT�1�SF���G�������2�@�Nl��q��\�Y�̇�$Q:B��%�UH���cƚ�`͇����LMԈ�9֔��p�}Zv��51G/��ş��n�)&��t��zv*dy�ye�\���ʰҨ�lX�/�B���  �Pq*�%dϖ[<je�滀��hVa����?~-k^¦����y�}?v��VUmx�ʢ��U��c���㎘k�a�{b9�t�5踝�V#,au&Q&�2r$��G1׽L]��@y��Շe
`�h�T����c~[qiM��� `Ǝ�����{�z��ge�u�X�c�W,Y�堡���Y��T"�ӽV��W*bA!��r��؉�]G�jL!���H�#FF�Lgd�U�̕�����/��ʷ�Suɳ���&7(�?��P��Wخ6K���%a����[,͝�-����9w�-N?g��:��V|
�F�	�����H�[�+����/j1P��8���x��Ig���럷��d�F}�PdBz��,��t8�D�wJ�=��$���}���d;�V:zЖ��f,K,��� �]������~�O��i�j����Pgn���[S늗�A��k���~��~NK��+Ñ���u���
���4�Lg��\��#±��d��^w����ê{�wI�q��)$��.j��i�pq��\>_�[������I�fU�og�*�~��	E
�{�6��Y򁻇0�Ǘ���Tr��h{W ۥ����+�(���t�^��p�ת8�0�k�H�t7)F��Du����q�ce�al2��:��|��}���M�����������cm���v 0o����?����?�v _���>�o��L����&q�d�L�g�9�0	���#�d �rl x�ds���s��	��ɜ�c�6���\��8�d0 ���d�� �� vs�3��ɓ g�m�ѐ ����V���wq�m�մ ���m��F 댞�m��2m�  	�m�L� 	���&M��3��ɝ��&v�m�4  �6�dɀ3��ɓm�L��3��d��m�;m�L���m�d 3��dɶ�&p 	� gm�ɓm�L�d6C!��0{8��d��&Ll�����}�!_����@1�l9a����W�����@������u����O�	�����8����o����������?�lm�'���o������1��� cm�� ���@���|?f?�����_ݿ�����o�?�??���a�C����f?@�6��q���_�������-�4ll�l�0�0
l`�D���m��6�8 ��&ö�g;m�q�m�q�m�A�m�d Cm�8 6�d�m�  �6�g& <861����!���������l�c
C]�������@���7����
����x7��?���~�߿��cm��?������߃���yo��?r}?��1������6�?P�8?���7������cm���lm�w���7���>����1���xi��glm�@-����|7�A����?i�N�w���lm��G������?�����o����(�����a�����?�{������������?�cm����~D��lm�p����q���LG���������7�@?_�!�������lm�c� �~��n,�������뾟������~ݿ�6�1���|�H8>{cc�~��?������~���b��L��x�ato
� � ���fO� Đw�{� UUU)UG��l�l�El6iR��U*�J��!E��)��lj%J�PBD�kTUET��
�PEQ!զ��U��U�mhhٲ�&V�l��`�-n�D���FH��K+Z,����)���h�զ����_a�#�j��J{�8͋Y��͕��[�Jse�֘���4�Ƣ����e�E��=��VR
l�Ī�l�Sf�D�6�ֵ��եkm�c6�ً���i-���cXh2��m��7�8͕�ƺ��e�  ������Wu;��^�i��h�s=�=�t�Kw�����Wu駴=6�Y�NqP�h��u;�מ��n�V�k^�zE�]��zW;ݻA�i��{����v�늬�VLl�L[m�Ym��W�  Շ���t: ݆�h/'��� ���C�>��z�44(^����(hhhV����/���S��N��nN��:�g:�w��h�n�=o7�F�N��z���L.��Թ��jn�]��L�Tu�:6ւ�!�RF�   ��B�/�-y������h�+����w��]���Zf����{�^f���{o{X�;Xݷ;mΎ�v�Z������k��[b����z�i[wr�ۋ�m�Zk�(<�`��Ѩ�Z�,�|   �z���5ӷ���w;�:�mwux�֪��u��w�w�s�`�����=��ݴ�Mֱ���k��d��z�tv��w{3�5���C*��{ڶm�i�=R�6-���6mj�����  9��i�(���{h�̬p�;�S��e{5�{q��[UEO^^�6��z��OJ������UM<w�z�B�^9cf��QJy2�5�M��Q��6���  ������oy6��Ůzު�څ������^ڧr�ʪu�]���5��ݳw�;�ƍ7���kZ�����U�6�\�ST��zTSR"�����j�   �}�m�w:�%���J�vޕ�k���מ֨�[������e�Qݫ��=UUsT04 �ˁ@��o����&��k1m���   8�  � (!��JGs� :n7@�Μ@��  9K A|܀U�[�\ �kԉj�-�Z֓Ik_   M�� �y\
 4���������
 o]�� 3Ӝ( CX Bz�:  m��  tZ (Zv�Sf�Z��ٖ�jm�����   7s�P .ݻ�
�v�P �v��7.P@.�n  �m�ZP f�� ۹� �ڮ ��"�ѡ��J&@ �{FRR�@ j��x����h  "��	JT @��U%F� a&R�0�S  O��??���ߦ�sw��}��������tFg,�`�	����V�Vh�e7�������|>����f�������6?���1��3c`�����d�cm����}����}�v,�T��?�f�°|ǳsg2�Y�(QxַN�	nPr�Hm�V�5�L$a���[1;�vh3/^4'��e��+'�eo�����H�bR���9{z�7x���
���Z��l9���v�`9���Y��j웁 ��ڙ2����1͑�j�;q�����PՂ��1���R5�Y���e�K������eks/r:�w��b�(Vf��+
zw)�L�Z��`f�ܖ���[p��dY�nna&��l*�+F�QQ��&�����ՅI^�C 
ͭ1��Q��2Ҭ����յ��yM��,�5�	�;0�+@�`?.ۉ%g��9u+MEVkm;z���ܺAkՁ���g�5�N�j�Ŭ��Dl �"D}��NVC�k#�Ґ�]�a8�x�7ڂ�3(�fR̟+ٗ&a
T���[R���.�b�*�n���F��W#"E�TA��ʓmjw�3TN�y7T�"�G/J��ꥮ,P����	k��+%aL����@�"�b.U���%X�:���+{o���v��̶C�ͭb�T����H=GU�)�c�TXC[aR�e��6T�άpPR�f������E�Oa��*.�2�"�VP��д�X�n�h��cŵ�՜��B��c�/	���E��q��P�Zf!��Z�sRMY9�@�Ӏ��v��vl�n9���T��%��6����"��,�UBf1*^b-�E��N.��7Wf1�U��R��amӷ���S�M�נ ��ͩ�-L�Q��iz�ʑ�SS&����l{��'����"4���-K��&RǸ�ıY�S��j��-Fѣ���
�>.����n���Ә�3i@k�d5p�;�,мV�7�2��r��6�<�r"*�;�u+�0�N�5�u���̦�6�M<_��A����2U�f��&��ʶ��B6��gT�y�eGF�6�Jv�V-!�nh��໒�JݙSnӉ��ܠ��n���ו%^i����>#b>�'̴LZy�i/��a�*;���ʶi��l�B���e�k)`]��&���bb��Z�s4���jJ�p�Z�Y��H�4���	����0Jk����46���ix���8	�3ZI�EAR��kT�b�W��3q�l��#&Ű<��9���Ѹ�.��ŲT�nLv�d�ʡ�Y���%�Ae�GF����TQU����aDpǘA�7O��iּ(b��Z�9H�s0ފKF�C�E�d�z�<O1e��m�X�EJ�جb�j�ڲӴ�^��Y��7�4䤡�$��.��f=ʰ�)�4�[@�j�{N� hڸɘ��>v�5��m��3!B�Z�ʃ���4%�EV)��a�e�ӱwnm�2�W
� Jn���
��Q�)���F���D����!���<A�u�^=��t�
�����}mQR
`�Q͢c��`��Qf�@K�V��3��)Z��l�z�#5!%��1O�୒�π�%��j�̂ʡ��W��
b�\�T�^���F�CxE�ٴ�������%u*\C%K1l[��uj�O�V�:��y)�!YyMGe��\f� խ���J�2��MBbc#Q�R�ۭV���b
�X����I٧�`e�X ��O�ơ{���J��X���c�ۣ�:;fl���[��,k���4�Gur[2A��.����V�66�:�f�uo.����e͒�$������&����,?�1[��^5�f��$�N�#���ڲ*�Ƭ}��nXD9��ۑe)R���� 2�gq�.�@�@*�Yr -M���h��jPյ�
{{ғ2����� �J���#(�Э/I�ˬ�+`�)�8㙔�<td/�*=,��M�)��Њؤ�OEL,�\(�J���ޜwlk�Ր6���lK����[���V�eh��fļE�����h�wB�Fc���8�VC&�tt��Z�:�+z�<�.�7A\�(QJ�%XR�z2��:�L2�2�u�\�X�����a�v����V?���,z�B�AE�a�v�VD�1ޡE�^�̱N��l21��v���$��U��X�%dH)�jP�Yb�2C�^�����(�4ܤ��V�a74m��nR�qi���7tZ]ٷI!�[�x��W6�*�./��a�x�I�JTڳ� �xZouՃ`�Ma�V����Pz1��	*��-B���zUʷw�μ�Sr���eˉK�>FJf�C����[�jhM^L׭��c�1LF�̊�-�MM���ݡt��3(�j ��t:7̚���w�l��hF�X��Fں�(�i�J4�i:f��a�[��-C��e!�jٛ��j�����C�.�a�ݗ@��f�W/fJڻ��6kT�M+�0/]`T\8�F��vd9w`bWh�u���R8ۋ$�h�(]�� �Ȩkv�4!c�CK��81���&�E`��n�J��&#w���Ÿ́�!b=W����G�ݻyj��A'Y�%*
��T�r/��m@�ѼEj�85Z�u�S��d�J���96�=0��Y@�x���࿖�cV:,���Udy1�����7kr[I���S0�\5�YI�46XFVk4�|��nR�W7)!�1'o�z� �7~�b�靽���E�n�L��r�����p@�eӸ˸��"n���lTצ��w�2���٨��1���\Û��z�N'F�Ќ���^ +�qۉ�� k��w "��ņ��[[V�OS�U��W���x�3|�ܨ�G��{RƴX��H�ɡ�����m��ݣiaW1�:.�V�6b�&�wkh���SR�DEk��a=x�R�OkvI��v�]�N��04��6M��0��S���h�ۏ�b&n^�� �ݡN�q��f�Ҝ�ګ�D��� �5��àt�Ή�p��d�ٲfCp���k���:PKZK)i/�\�*�e���cpa�A�dSN[��
9,F*BN\��\�و��872Z+��ѷMhՅ�o�(��YX���&�����n�7]G��b�&��N�J`��a���y�T0��f�[lb���6՚^4��c	WVE�t9�������uel�5-K��yx�e�u.�ɮM
����@��Y� �2@ο�f�(��LZ�A���)�k�
��'6S�	l���V���RĨ/��
C�-$[;mM-�3rk�Mcg�պ���1�/Kǎf��C)M��7-�! �hJ�JݱhfdR�����1{�a���2�<A�l�j^���!Q]M��$�����e�Ր̩.ɟ0O�m��a}�F��H�t]^9D]X���ŒƤ�4�yP��^�F:�&m��#�Z�7b[����N຀I���X��� �C�Hָ�� ,����w�hgD{j�����,�l7��]e�T�;*��{JZ����.�*/v��.@�l��9v��*�V?*Z�#�;��0f��6VJ�bX�'7^5�c��E�ovVts^'h<�vr�%�
�,Vl��2[vv�B� �eм�E�w���
��^��(6
��=�,�T�
V�X�G:�6�:a%�-6-K�����B�Q�-�-�a<*t[G�ƭ
�n9�cvk�u[8[���_wy"��{�yO@H�@�z�4٘��e�M=r�e�sZ[�09�hDu��m���O#��0�u�FIw�T�$������*!
��M�e�Y��}���XM��;�dPn�2�P�K5�5�F�i�����ҎӴ(9Z":���m^l�ٴ��-n��zz���N��z~x-�®��n�r����A��Ŗ-�/+�X��؆<��eA6۬�R� k8��2�F)��䩒-h�3Wm.=���9����NB�5��n�E�$ĵ� (��]K,4���[�����ޑ����V��1RWNf�y�V�[���ш�����N�����Ku�r�v�ֵF�$�ƒD�%M׸�9(jB�E�<�Yxn�+h:јUЪ�61�<d�j�j�B�m;�Z�	��ւ��#q1D)E�x ��`L4N5e�ʄ�͍�G&D�qf��y%���b��Q%.���F�������^Q��*Nbh'u��c؍hȓI��b]MF���!���} ��5����A��{_\��Z[z�9z�<�Bv�1-8^��  O��O���z.ƬĳQk��&&�j�R{LD,��Ы(}�"/bgi⧨��Gd�]J�2��&��OHKr�;��+b�A��a7�A�^c�UJx����ו�:��Qc�t�rfU�f�a^ڒ����2+b�"�[X31����:��f�l���QP$��5�{L�&�R�Z���5�혅�{���f�66V�!6��T���
xe��,�ژ��jY���gr�S�k�r�M�($�u�)�Xˋo0G��x
�Ye�tr ʡ`5J��)B%��x��̔��*�a!��jJ�ް����桵����l=��P��[����,wA�si����SU�J�%w���D�l�šbR��=�YFc�	�47w->� �Y(I���^����Ȓ$(�c1��\��I�ƕ9�lx;�LT�fj�6���om���I (+��)�+6��r�^ڶ�/)��#��9�[��-V�x1��?���kV�T3&�fb���y0.�3;�Y��ʇow�R�CC咲�W�(]�e�$�iˀ^8>v��XnR��:-�@m���u� Z��)TtM�Bj[�mk�x�u�ˑC���iSk�Ő�Y���6���WwV�^��Ui��q���H�r�H�'�.��b�$���-��h��f,�xnS�1�w�7���W����)u�el����[uy=h굘5�GpK�oL��c�K -!u���E��K+*%�
Hk�����E]%F��=���6�
D�֒R�����V�4������h�-�cp\�>�%����Κ&��4�-[[3惱�W5�Y�7t�MՓq�*Z�ێ�'�%[s&�5�Z�F���C���{���n��	�ՏZ�,R�2��,�0�[G�#��cy����~v#8�.��Ԓ�<!oN����H��G�d̀��d�=	�՚[&:�̎X����㢏�d!`�*Y�p�L���[N�-��d1��E��Q߶U�8�:.��Y$��V��pTAa���f�W3C��1���c $��bg���=q���:{X�����L��ݶ�f�hz�n)�V�iQ��3l�F�X��M;�[��%�z�J#q�-U�Gwh�./����@z"v@N6F3�,C+3q�E/�젥ձ�L������*Ճ�˦@ƃ�V��Tȝ��"��u�W����X�V���(�%G,�	�]h��;L��.����P�z6�D�,�;7���"��9n�]�MdN�m[�X�2Σ��с\ ��]��#n�f���������J���%Qh�ȍ�6��J�OF)�ST�+���Ƕ�j�´l�:�+Z�[oql�B_חX�r���5c�1=���3t�ͩx�lw�#c@���D�-+B(�k�ŵ�u���׭�IvqX�^��P[����sE��f��Y&��`e+Ŵ@���˛��x��SJ[OBI��m�a�
��o]n�h�[uGP�V`-cnQf��Qe`����;z1��N^!,��i��6n�t����H�ˤsf��`Ǜ��Xb.Be�G/6#x�KxM��rl��i�P��j�נ�/pP�(()�DWLZ#TXܩ��+1 h�Y��.�n��E�S�e�)#36��f������K��l��K��b������	,CpSs�Y��FV�Z�ѡ9��*.um��Dkd�A5B:*a�k�׺���ݖh �7���4-/5�Z]���@E��H(�p�RF�ݻݻ)d��IrZU-��^��ߖ(m�K.�������Т�d�Y���6�k5���7&4إ�*��mZ���5��P ��������9Ku��ۚ�㙢��д�4*��9uzv�,�w�0�K��6��)���p�>��inZH�YJ��a������[�mS�-TZ�8B%��R'�@��A�&�/w�����bx0�ٳgp�Ly��V���K[a�m�]1S��W��ōDnC����7�`b�Ǐr�i"b�o���hU�-���jJ����i�h;�Pa��2މZ����8,��Z�ʂ6t��Téǋ]�Ud-� ���n,�]�æ�]�( ���Z[�Pi�B+������E]��3/b7�P�ki��	��Q�u��GF��b�U�wo1�Rq�T��!lGsJ��"�-�+~��=yxMZ�*�V�Z�7e�ɲ�I�˭d���Y���ŷV%�IL�i �jBm�����L�a
��U�u&E�Bđԍ�л�r2�n8�(��G�b2�tU���^RA�Ĭ o
4#�7,jkIqc�nP�M��l�X���s1c�(��V�MQ$�ϱ[߅�����C��R�r�Ig�VjjIm=r��MkDN�A滽���4n��QEVq=�%8�%�l+��n�-�c�A/ELotIW,@�+(�]����N���eLn�VE�-<�.�s��% @��j��X���Ek�0T7{,ථ]��$�Lo[�&V��-
������L'E�L�T�q/�Ca�qA�6@�V,�ӹ[c�2�TyR�n`���x��[7���K��잞f{�bm��nY������Z��sx4�f��Sn70�`ٯ�"-s�[̈́n����:9�IT�nX�7rW}��%[=����d���(A�V�̞'C��t=\U_;��6)�mO�h̥�.�K�nk����;�q��@�u������Q�}w�w1�{���w{p�!��$i��w����f��=�C�h�ѭPP���n\�zCHf����t�:�G92bFr'��cܤ=ͱ�k�Jsc�[30ha��W�>��у�#��`�Ip�I���A��l[2j|}���T@W�lg�̺Y�1�\���<[)_s�7�k�.h^��:�2���D�[P1���wX����P ���W�ڜ�C���ӷ1�}��u���2�^��f��Xvr�������0b����.�}7 qǡ��#C׭��(��[V{Z�A]�p�v�{�u7)�A݊7���@��w�
y���Gr{���=��:Qt���s-m5R��]*5�p-��f�X)
1��7��s}Ax��N�5�����M*�!dW[�ǻAG�+�v���ה,��t���}�R�%w����f�d��Umsݧ�}],*�}��������i�v�A,�S�	�����5ۭ�6އ�>�2�Ju/��m��1�׼�)�v-f�T���!���F��Ơо��r̼R�Q܈Zq>C]��L��o��͕y�r�|�VZv��ߞz^�H��A���R�.g yt�Ǆ�vtH����k���9��(�c�&�G�v�
'C���Xs�vQ�\�귺��
ZaO��O޻�T/e�J��A+5��ăj7}Ym3�;�2^�^� �U�[tE�^F�/�SOy�Ħ�v56��҂�ڈs#79���-
�m�.��N_0���x���G��җ�VF��LK�U+˱�4YBrf�[6K��j%-�)�H8w^�y=��l̢�ά+7��z�-�E>Z7Z��2i	��D��#);��\��u��v���I��hk��Z0/x�i�{봑ݖ��1R;a��kXOf&���`+��i�5]c�޽W��!���)�p��t��V�U��Y�6c�g�sJ�o�_f�E�zd���.t��ߖp�v�秺��Ӳ�7j,$�g��"��k)��PX�%�a��J���((���鱧�e{���5�t{R���)*B.�t��	\�ob�A�ȯv�ܭZh�Ͻ����o4= }�f�B�^\�l�]��÷�Vp�Z������=�ī�ܝ�x���o�dB	V�+�J���A��GS�)o[����*��L^��1�o+1ΊY7�f�5��F�[{s%�O6Wi'9��ΖE������:���G�,&U�ږ�j����d|v�k�b;õض���L��k"�'48������M{���u��m^�F�LV㷳,{��s�qm�cwE����.5��z�:���Ç�Bd�>y����xϵ?s>��C#y�+�;��V���Ù���$�*�|Gd�j�H���ww	Q�UNgA �c2!Ţt�'��>/�o*XGu�AZX��+q�oyħہ�(�Z���z� ��<<53"��˚qY�c�y�9�Sjw;c��uR]4��X�U�R������*��{����V�r�+�[�;T���޼��A���9���c��\B��ib�sn�'y�j�[�j�"�b��09ˋ�׆�(��"�A# R�dn��8�9��h����qG��r������T���2K�(\1�3+�+�-�aѽ�)��o8vc7V3$�jX\@E�����|�'�#5�,�o�����;K�EI�w��)�>�v]��S�r ��ƸH;���9�t�j�T��P������CZ7���͚p�)"��4�P�L����KA=|ҁ���5��v��Sg{��j��������mi���.g#���YZdWd'h���H�*���cm��{c{��,�B2�iS+L�5ؠڇ��զ�6���dnT�j\��tS:ǖ��;��i=k���A[��Af�0�Yqo*�ͱ:8!,�t���i͹�����Py����7vY j��;Α�&5c:O��o��t�sb.����\� ̧�7>���r6���hfw9��S9ϙ����a����<�[Z�+�:Z�Nt�5��6����u&ˇ��x��&�V����m��ip����ZN\�_�n���9lP�R��JX�]�td��guٳ�Tm�줹��N$Tz�4;e<!�.vr�x�ű���2��|7��X����^��kqFc����09D�x�1�u���:��F�}:ŪpnY��F�B�[���Y�JZ��?P�\�O����<W]!HP���3o��!�)TO�is�S��c�'e�2�QrM}b����]���@#q���/�]�]Mz��t3��F��RP_����3�Ty��9�����j���!�GZ��&�~|m��ή:�@�9j� *)��2t<��{)-0̅�eݷxO**^GW�ތ]C���e����&�
��U/T+o9k5Uc�lsm�)J�`*����n�-�NrmI��fB��R��"��,���qp9ބv �^^�{�V�f�'l�D��/����iNN�ah�I̞��k�w�R�Ů�5U������P����2�%5s*��Ot��sI�{�Uv4�ג+H��yI������)q�b�m�s���/�������z�/�>s��M*̓x�ׂ���
l�˒��*��R��ǤO���K�O��f?��74�8KHs���g��Ʊ-z5�F?z��OR��FEٚ�XS7�!Q;#°=�[��崋�{-M53�"�{V��i��"�x���ק��Ӻ�eY7��`�9\��ۑ��5�6^�|k�suZ�ͧ�Ho-?,�S�*Yɷ{8�C�܍����
8��N�_Xv\���]�ʧp2h�u�/oU����Z6�}�Q*0(r�qV��7)޾o
u����{�k�*���Z`�����Z��u��yl"y�{4�*�A�����U�`�ou���1�q�h+u�k�)�v��e\�᡹8������R<غ�ۻ[��0΍�}}EF�s�ZW�`��l���9/�76�0��{B!��w�����X�Ks����G�B]�K�qmb���Jhv�3"à]L�����h�O�Ж�ɣ�}Ꮆ
%n���t�{��$ނ��GNEm>�u^uu���ذm]t�.��S�/�Uou�ᾙk��)n�����e[F��rn%������!m{pޒ�F��P�;	D�u�a_=n�,�A�V�ڱR�|qPX�ިE건�GlWP��é��WG���w�t�;�F۽��k��a]5n�<��0c�8�Ք]8	&m�Hs\5}Y��vӤu�@�����X�e�޹�-$d�c�}��vU���*ۗf�,���d��k i�J����YFsWV�Vl�U�H��������\�2Z��-�I�Dƃ��6<����(�L幋��rA�a�t-��)j5H�^K�Ś������j�[��wE����Mޔ�IF���u(��gFk�Y���^������~�eC7P�'C���@]�T��p��e�`{8�9giC���
}��)[:�T+�5�ӵ�Uؖ渻q,�6��h�e8��P�ܼ�{.����e��r��6b����7dŌ��w�:(|0�dMT�Ǹ�f�{C�v�����-91�.������]��R'�V�%�9
�C#�8�r͢���H�86\�}G�����A�U���!ԇ�̔��pϴT��2+�1V��VJK5ג��,�I��tpA�,S��6���No8����s�ΘN�[���/4�g+�u�B��}
,���I
J9wq�����b���j��B5s�z}�D�۵�ת����Gy;�\K*�6��^�0c�Y3���Ѫ���U4�6�S��֪��k�n�3T��`�ق�*��;yl��j�E�Hd�ڜ�{l8����L6o��I:p�Z}3����p�O�I�Zg��|X�3q��rm%笽�)�m��<����$���ו�!�.�v��������UMS�� ��޻�4����}��#[�+�o$��cDf�ܺ�w�'����Z����������'{o�9W�] T��¬}}.�����;��p8B�E��d���Y1�e+F#�tϵ�bu���������sA1Qp�Z�M������h�NoU�YԞ���KJV%�X�xO�7�N�,��|5�����Kz�QCjH���:1���Qip!]G|lp\�-����R��V�n�f�� �M�V:o[������9��Ir��[��3����DgL�ljZ���tv�w^��L~���O��-(s��y�*o�wl��^{�t�: ������<�J�df�l8�l+$��_�%�U�(<��P5���L��@oS�`ޞ�Ǭ>z��׎8�p|ސfC&�ˡY�ƹ�k:�X�!�e����{�6�<��FwM�I��(�7Y/�KwzV}|�Z� ���8����^-ݩ�1;ת�������"�`�G,S�iN��p�W���͘3��s	k
��7]�,=1��f�e�����̑w"R�w��u}��έե#��.}��i���{v�P��:k�x;]mpa��W�I�;�7fetg��XE�����	"xJ�k���0��t?yի�I6Ey/�z���E?���Gs���.ɭ=HY�V�|u�t�N�����t_6�8��>	�(͛;�kL�F3!	��xRھ��׊Su�T�G��$�3ښ'�7[�ĕ�	��d��[B�ҏ�<F�3QY�{�:�b�J֥t�M��[��' 3�׺��p{)�^
��s�,1�*�GV��D�걡�wIAס��L%�\�Q)��#�*f�w* r�ѡ�Ձ��s@�tt����;M釰')�y�rf�e������ҸĽ�zWe���k/T��,ۭgZ���U�|cp�9�up�f��|��.k�,f�;|�>s���}���uކhy�q��tK��#�3��ݹ&T%�yzw���1�ʊ��25�Fj�;x�U�<Y](��vk�V���ī �6������{j���=1�3Ӭ��ֶ�pq��'�	�A����T!Z�
��m�G�0�HN3���� u���'F������^�BQ��Q0(��UN�ԁV�K�:0�����o�;�&�e�yŒ3���8iꀌ��^�e���E=��,f�c��FK=���n�6�p� M�f�u����y��N ��뽴�L+�j/�d���V�Z3�f��^t��H~�3���z���_:^�,��szOD�	h�<F�%��ג��*>��hØ_SGo��*%Ic�������ͣ1*�51[�Q[/�����.����{^}���Y��#���Fe�&�:Q���kV�Sa���7�EU�ݐs:��f@��F�-�"O]��46&+��Erb;�4m����A�۾G*�icS���\�� h�+̾{�󥅔��\iV���co�����y�vJ���`D:��B�kz�3kH��Q�I1���4��כ��8��Ut�ܺ�kC�=`P 4���6���{��Z��-�����:ƃ�s���'n�9�zV��T=m>�4�n[a��%��[I.�(<�XK{��-N(x�J.����}A�\�>Re[����sz�+[����܏m�@�rpO]5n7T���rxݛ^'��Z/_+&Zr�Vb�O-�x��a������f�sO*&�S&���"��FWr{)WA�E4���N����2���Ǟ���X2u�M���f�Jق�G��]0�ܻ6K�]����P#N<Nݔ#�~�v��k�n@��x����H懛�=n�S�g����s�8V�ԛc~�1����1�՛�n�l�0���{E��׷�N�Q�uj�rQ4�Й��q�����Y��Q%9��u�j�J�~֫���u�t��sw{l(�h�B��Q������������-FZX��O���\��{z"3᷃b�r˭��٥t��,պx��wv鱶$T�2�}�֜��1�9N�P�ޝ�(Nn�:[�!�;D�[����)/��.�D����x�)%�Ѿ�;�Xʮ��;ҔN�-�ݔ���*�-��� <�K�ƱWh�kAJ.�u�Dk�B��K��`�w��u�̻N�����"�G&x�hO/3���̉�\������4q��z�捗��o���F�󤊣���^�تV_����Y��խ�0�,p�.와)�����/�s��Ѯp�:u�hcd��L�u\��\].ָf#�dZ�*^�BiK�)(��)vv�C����w3�{�7�"�ϫ��^pq(}u;o�N_y��ނn��:���352��|� ����wz>7�s"S��z��,Amn�'�ws��S��u�V��o���2.�=���=���tə�ǫ�f}N$��W���6��{�O>Κ�vgI�>]'k[�{�V(�!��څ���c:$:�֓wƛ�$�������@�#ܝK��vޘkq�lEZ.������PdL�`�%����gz�X��p�f�9�ޮ,�w˥���D�e��V���GPc+4��]'ٛ�9JEm0]j�xF�]���oV��ތ��j֡짽.������f�+�V�n�uu����v�ԯnt����ݷܶi�1ťf�K�]yS������Q
k7��gBz�����+x�C�"g�=*�fQ\7�46�::�����gV0t�
؝s��u��jw8�a5ܾ|�����ll�c`������翷�����ͻ8��"��2��)���/�o'Ħ�G;�$�Υ�SVA�h���a�O{8m*-nP����N�16�X�ؓff�B�⶛�mvˎmo)�Vwply/EO,g3q's������ˎ��6pm����S\`����
u��"��0Ռ�x6d�bK]�#���P]�����-a��a�͋���G{��&�غ#��՛�]�⬔�k��:�����||�9�оθ��&�/3fr�Jnq�$�Kr�э�AUΤ����}4�1?7�zl�U�+��_g�����kWdg,�M���e����ҝ����o�˛�����(�zh����cbZaH�1��.�S�-�$#u�i�E3�V7Ď5�����1e�e�<�q��C�D�u@wwЩ�#Ʈ���U�����[���-4�-�;{����7�.��W0)N�V��ݢ�5þ.�YrKOyb*`1�Τ�l*pz1j�:*P�wQ���zU:|�1}�qzq|�!��3��|�L���ɁI ��{n�a�x��%��]WY̶̬1��\y��P.ޝ�v��{�b���$+&�s��Lp�ԞJ�� p��ms��!N�n�+��p_v}����g��e�PWs4�ĵ�*��#�R�|Ψ�tk0���O��վ��t��W@�;֙>}D�rz���;�r�BZ��#�儦ŉ�+���e̻��Q����p�7+�t�΂�qn��min�����	���� �h)j���V�n�*����Rզ��ˇǏ�Sm�1|R���gc<c[lB|t�/�c8����Y\�=d
G�����u�p֐7sc���/�5J�Ф�F�k��Z��B��w����3�ي�֘��b�j��8�\�#|Z���/)��v�K3�����y�v�b1So u���Ve�G�q+X\��^���ڡ8�ݣVU)����4���n1k�I�,_A"��t`9W���n��l)v^�G��I�#�P�V���ӧ�V�//^��-tp!�#��e����7{_gfbn+�^�z�&EP��_)qr(�_v��_)��$�!D�n�5]���F������1�-<�C���l�R����n�u�kF�5��X�Q3���#��ЭU��P�����:�G����e��T���yW�gϟJ�t楃D��afq��3���#���\R�ۭ��K7�8�(�;�q���K���N�㸸8"�U��)�u.�9��ވu���fs�vuQ\�K�o,<���kU;�k���_�RۇvGp��a�L�*e8Wl�c��w8�,ih(_|�C'\�ݾ�([*�R!�3&���i-,[b
sj�}��8l8ٵS_��D	P��ꖺF��k`�����k�igz��]L�k��N�ݘ��u��8A6�����O�Xb܊���T&(����,�iw�:h�׊�+
����z����f�K�j��~�}H��ۛJ��L�r�
H�]{�*���қ�L�Z����5����̬廍8t\wZDy���u�a2�i�����(��,�����^}���V����ִбnK�!$��m�X|^^�T5���:�M=2�ͽW���w� ������}}�i����y�}S�8jJ�w���c�[�LO���Aǆ�j2f�%�:�1�7H��A����Qf;��v����K�Z�4NW7��{����<s��V�en����y�T���X�݅e��P�o�-��ާ��\"Qh�RDc��K�^��xfh|�k��4^-�B^����u��]yQ��j�E�۽�Ջ�ۑ��z����b����)]�b�z{����C32�����z@7i�J*�Z�7��=�G�}�۹��k�ͻ|��(�������:C�;ژO|�vb�z/�����)���T�Jj��ǜaH֫�C��j�QH6(�K��Ǣ��S{�j�����8Q��5v���xS�Y��ϸ�)������.�bϑlu:��ø��r���7=�O�W9*1ۍ ��s��q�?,��ù��r�3�#��ӓ�OZ���3+쀋�3{Nü�6e��CCpp8���*Ă6OP�����|��/`#��Rdrf[ws0uN	�}�q���\ޠ��?f%��䗶���8c����{v{F�'M)��3�w8�CZ.V0[���Z�sf�<|�Q�vW;$ה��e]Zt�n9wʋ��wg ��-	B����
��̼V�ŘLJ�Sכ9ʂ��Fy�c�J��m�zx���ކt<;��p6]b���*]�P��Zr��J���6�,`N�@� �pRr��b�d�+H�Q��|�uh��czdp

�Ͷ��P��3��3,te�m��[*]��F����]Y!�e��Ya|{OX���o�7��}��+�{��zJ�g�Ki�����a��\�ޡ>kl����\��%)a�Ӧa��I�{+rkUr�.K'�5��$����%�!���Ѡ�zΪظJ�5�O%h�91���l	Ɔ�q��]��M[D��&TZ "���ע�8�Vu
wR��p�oc��N��-J*��!HG5Gs�+,fjy-�C�3{v�E^}����F�C�	IU���P5�h�d��J�J'cR�{��cc�[}t�v<�r����m��Z�U������>��1�L�m�ٜT���,~�P-���/Y�Ys�%�㾼����[##�aΤ��F��0wZݡ4#bp˧^�����ƙڻ�K�-�z�U궩�oRZa�.���j�喰=��(%>���`��z7�o_2σ��Ć�Ȳ����c������Q��>ɔٵ�ܠ�IjX�B,NME�p]��]���&��M�U3���]��Vb��M8z+�Z��ocv���Ǩ����.��g�MQ|�'_*��n�[�2K��:�/�M&�Rbn�U�c.J��MLq���{��-a��#P�'v-��i�K���[�@�X�z$Qڎ�|��e��k�A��Ri��E˺����J�=�������n�=y�_myU2=���I��9���J,�ffs��瞭���6�V!峻gZ�X4�LUi}�-'�Ί���#J�V��<G�x���mTui>�9z��8z��%4E�!�B�¬�1R�8���W�V�J��;]�j��̼o��t�/������v/s��E�V|��Y���`��4�}��RG8�,��H���x��R��Zh��vd@�*.�yk�su�ǷLZU��L4��*G�7,.�c7'�9�j"��-i��f�hTXp�l��{�kCr��>�M7�B*�h�N�;d�����Z�����,�֦Ӵ����B���n��Q�=�gf%H�W����{���sCqF2S3�X8�U��,�ujAe�{B�lKF���;Uf��� +�詗�CiSc0>=��܏A'����F�vDU4�-�3evQy��a%vVVgз!�M�x���1E��A0�5e��'1��U��B8����
c�zŭcZ���61���#��slu�RB~4w�n��L���`�k�:�� V�� �*ʷ�/ҹ�y�gh�`<���Ry�Y�.+���lu�4���Eޞ��޳��~�a�cc��ﻗ>����N���tj��w^��FL�T)��N΅�%����=�i��sbbӃr�k43--�o�k����s�������0��2���aD�T�u�+i����7�éV.�3��3�Jg-돃Oo����Y��PfNX6Q��'v?�uC >��5��x�+2�������{s��j��R���6��H!�F�Vk5��$�te�c�����4:������}�������8N�]�ϯiW6G3�o��༺Yy�P���-�n�>��M��"���D� �n���s����:v��.�Rad8�6�D���|�IR�{z�#:m�b(\�ڱ��hZ�jn�x�;�+	;b��)=�{�V3����؎f�a��u���nӼN�ֱ;@����>oT!i��+�=���m�o@�(G��q� ��
�ᬸF���#��eg׎^kb�W�or��ω-����5��[VXG�UTsLa�G�>�Srj�HԦi�
�`���zfRia���e^2z_n�+m�Y�;D&\0��v�c2�'=2n)�72g`w��@��d� �H[�Y�U"9:�4s��ا.�� ��Ż�\��/���8v�<�lU��A������0�-W���w�7JU'������\}a����3��΍Ѵt��&�b�vT���
fpD�8����ݙ�)�%�_?Hxh��+Ӈ��L���:ؤ^Ԏ��_V'Ώ%о7ݻG���	#��H�pV({)�yOg��R%�k{[��ݲ��(|���(7z��P������M�d�ZT٪��c�m�C[�YMmb�����S�@{E���c���r��ꁅ�����_M���&E��;�-�*���7I��%ԟw>=�r���o(C�B7c��d[���rT�c��&�2�#���$B�#���tL�J�վ�7���}O�g�O]�^�9X,|.��i=n6|氛yo{�܀�<Ϸ�K��b��Z��/�;c�|���������`[�rg0�F������Aָ6t�֤�E)um��^��E�ʇs׳i|=C⮪_^�"��?J/C:��h#�f�
SO`oQRw+&S[��6T�%��KwC�դ��Ӎ���m��N��a�t(<�CHzŗt�b�>�l
/N����DGL��+���c���T�cm�	$$ǻi>�P���T�M�H�`Tv�~*���;-�%F�G]�O5E�����!e�)��M[�.�8�̦�0�2�cZ�5mu�z���Ǽ���\��3'+F�F�-jh��-��6|�ܵ���\��;:�|<2Yk�ɚ;�-� �|4�s��<���cè�4����'G\�]�H^]u�e�i.n�l���)��ut�{Z��Tb�Vu � ��<�q!Xu^��l��n���Nu�S_��sǲz�H�n�ރ�j9��:��8`,	�������@]=uop���J\�e<���F�
�Ed�{���x��8;W0��%Bu�;}�<�y�.�⛟Ms1ZV����Ս+�=È]�1��]�5wOS���}fD�N���e�������/�j�Иt�iv��X�ҷ4��Y�7�k��ӣZ�Ŏq́��S�i���1�=���^HC��>�-t�:�����9�`ӎ��L~g�{�z���kF����P��1�|���Ū�\�t@]w�`��D,����·hi�)̨����ZzM}��Cj�C��5qP���.cG�sg��1���+��	�sBWLrw\�/�q��9Qt�]�? �ДI������^��E��g�^�����3�<���9u|���;f[4#[��27�Vh�4^Z��%����)�����������Q#��==|Ņ�!#F-��l�J֦V����5j���&���Z�o�c;��,�Fʆ�Y�W�y�.�J�M>��*%���s��U�K�Q	��#�P�cm���3C紲l!^Z�*>r[�x�#i�p�#�㦮����:�*��;)�+�9��i�cS񾏌� �Uׁ*�����fњĉ�!cC���޸�#0ٟ,9��U��yS�\��׀E �\��q�;�ۺޞ5�ÝðV����l�*�'8��6q�}��q�M��D��&�ͺ�l%d0mf#x5fY�ѰpL�� YY�_p�L��y��jhv���
Τ�Xq����f+�6W\�,ky����؜�&/���w�:���G�-tk�Vm�ϐA���+sQ'$}U�#=ҲU>�:(�q�Ay�۱�S>!�mxVOj�_y�c�z�]EGG\F��׳��W1m����\zCZ�v'v���pd���ww{sj����t��Ŋ</���t˥��2!�Y�s��{v�f�5�<��������z���ٴ��=նVb#]�d�,��u{�4�����vљ�ew�ù�)i7�f��c��d��2�[��'ז�J�x�]Y}Ff�m-ʔٜ��+�=���i}S�U�u,��(��u:����������{�����V��Ȼ�S!�j�^�����}Y��e��&�5�cԏ7��Ɣ�	�� ������^���5�0��+̍��m=�o��c�"Ux�Kp`yV�%G;mZu�b�j�Ń���q�*{�z8;�����q����wX��	Q*��Kܨ�)�޻��ģ�a^��B�Z�Xڸ-o<]��}�����55[�ZÔqf�b�*Ĺi�(��[)Px��s>[�pW}�h\�:NoʋCt�����\h� Y5�:�'NK;8p���P�D�+�<�p�YR����t��jmN�Mw���].wK{���\�귮!�k���(��EzwQ�m=ξ�8gy�썽�γJ;	4�9��0޺��m������Li�C6��I8�L�V��P��bJv�N"���s�>U���TC���G����;F]%W�1�CR7�/��5l馉�Z��+���G,�9�rY���,���YZ�_ l�V�vd��3���V�@��A���<���U��k���5�����GW�J_v���/>��q�ʏm�A�oeF�`�3Z�q	�af�ًY���0�B�������X1�8�}{�
�\���;ۻ���NV�@���*�j�r�|�w�4Qڝ�����']���Mڜ�VH�f%�ph�,4Ӈ�e�����AQ��k3�X� N�P�)-��5��Ѯ�$�V�NK�[�^�U+�!���~}���`����� ���Ϟ~���C�H��2�9`��zI�a@�4[�o��#��G���i1+�h���2�}���9`ȝ�w�U%����FT���z���8e1nX��w�.t	�'�S�3�VL�m�ܺJh��
`V�n����r�j�����kF���I}��'�:���Ҩ������auy�RW�78^S�V*L����9/��������9XS�7*�yJO�e�����_5Q���)żFuDx����M���J���Se-U��-�'1���l`y�B��� �睤iy��-t�R8��g�����m�{�4�fI�9�O^����y��|9��X4s��]kA�f�NTl��
���%wb�;���u5V�P�������7gdwX���t8(Z���$���$�o���hަfu|`E�SP���q��rd�׽�MM��>;_4��#i��<a���è�Jc�i�V����$b�Yo�Tj1署�7[�-��g&{��0�^
.��&�v*˭d�W�f���5��5��<,��9���B/���3*.��:�̤��$��11Q�/�Ae�J��k���d�k�����N��W�zEB4�{��}鏵4FEI75W�l ��6�סn`�!*�_Tr�!�{��K�Y2eR�.�E7Vݽ�;3�{aS��o_Nu�ٷʸ��^Z!�_��p��n#��]u��QB�����rW��� Á]�bڽ����v{�e��Z� ��SJ�ZBUE=r���ù���˺]e�9^(��-)i��S�ʊ���=+�����֧���{�����/U*
$%	R,M����V����y	�ET`mP������n�A���=�)�^8�c���$��ԫwbz��ykwst�4�i;����!b���n�Kf����jyf2��-'!rY��y,.�����\����ʭ<�76�\N��wr#��G����s܏ZU�I�٩Ȫ�\��VeQ��FW ����*�R��J�\'P�
�"�-M	�<2�ú9ⴏR�d�#�.s�V9��U,���<:�9TF�N�C�.���t��Te&J��S�G*��Q$n�ȋ��Ns4�9w�E�wTD9�����\��=��B��T��TA��F�j^go%���� ޹��e�"�fA�=Y0�Y�qD_}sev� ��<�)�%�U���ܧ��}�y�1ϕ�F�� N�Io��g������G��xW��T�#D�;r���޾��{n�;՗p��E�\3Y_p�-���爼OT��Ά�-.�W!O}Wafy���Gb��4=n�Z�I�Ĭ �+�xR5��dW��)-��q*�/t{�i�#��{��|��e_�Yy���=��M���{��>@�f�'T}C�C�6��&���RfBn܋;p��~�!�:m�#�8��~5��-C�t���T���L��V���|=;��_�=P��z�"D�T%���JG�\��E���V�ύ�j�[��p[�w#��d��և�>����o� �]u<�<@�����'l.J��銳�71$ѝFh���]���0z��?�H�������c���>�#g��&jO��F�L�] ����&�k��H��ε��t�%�9a�A&Y[T��l�~�dCb�ew�=�9�wg{)��%����e�x��ʑ6�҇�{5�-w��&�5�
�s|��z�X:��]N���ݹ����s����ץ^4��&��Z��7��A�c;�7Q��SW_,���n��AKe�k�#��6���{�2�G����w^ L��?��hK.�"�Ď�[ә���nY�5 �v�0�9/��6������Ѽ���z�ĭi��C�e�<;A���?M,��yFk�D�
����{9^͛��$4�W�����@[����H����h܇Q3�&^C���`��K��V�u��L�i\����]��.��`Hq��_J9ւ/�����.?�h����0]��s+�z�VuQ0{Y�~22�@6���`'�1bM��.���o��9��Z�t�.�H�����퐽[�@��B��X��\4S�G��Tt|s�����!>�+�ƷfJ���&����b�pw��Wz�����6hb&yWʃ���d_�"�!ؾE�Y	U�A��n���s�<�OU�kh{lT�Ȯ��+����ɞ����ɥؽ�!�_®����h=KlV_b��aM��
.JfR��$3�3yߒ��G�8��G�~�����Ai��GG���e��7K�9'�;�7�B"��������L�2K�<�Α��ߜ�eOwv�K�N'�7����s�@c@��� �3��C�Ӌ�w�&�z(����+�j�g��Gԩe���,>�3J�9�k��F��$Ȉ�d7�z�7����� ��K+����Y��	&<��x�i���F3_q��TFĮ����W��Yp�
��.g�=����]�b��N�c+*l-ޭ�/޹ǅ��S��(*΍AԗS���c�t��p��]�EK��i&�bYڶ�Z32��.�=�٠8?�k�ʷ��U�tX�T��N�z�ju��K%i��U�4���r���}��)O+��舻2�+4:Y�1����FuB��Q��n(i�w|ra�R���nAt��0pr=8}�8�1�.)Q��.��r�P�6�%q$��[�Dtܸ[v����F:�.Q��}��f仨{���p���<1�S��k9����bI��k4��!J���Ц���NI�� �O@F�T�z�|�u�B���קq�Zk'(9�Q�@��BP���.��m��;Mz��T�,�K$5�7
gTk}�&{��x�3�4�m.S�_Q,��T���z�)�5��.���KWL���퇠�*���x��.�^w������K���(���,��F���x�{F�9�xV�z�F�ÉK��|UCH�aԺ��OZ&��ir^��g/ꊎf��<��H��u:�RIj��.���'~�ʞ�wh��H�T�DjOLۨ�%b������
X���?�Ӈ>8^厲+�/��,T����ґ��ԟ*L�,N�M�l����9X�H38u᠜��k�N��o�׌��F�]���ނ��z�O����Y���|�f�<��M��+Olw����B�d�wGS9ɛ#���~�,�W̙~٣�����d>˺㍬��SY!�Sa����q��6���*ƿC��7�p���.:&m=w+����6�f��<5�g{Y��	�� ��Ս���{\i=��ڗ@��+fz~oޛ}9����Y��u��'�ŭ�F��T)�NVB��w�4�u����&ܱ���Ly�y^$�;��Fawj����;��W�}+ܴ a�5b�4K�V�\��hQ��A��~!u�_/	3xެ�G]G}p���"��^��9Y����Q�����9��&D����ݪ�d!6�N��>ч`�X}�Uo$���3ǰk�A>�����aҞ��Ϛ���Ī��\t���c-I�H8�a]T>���A��I����Ƙ[L��B�6�����lF/��곘�T������j+�iCΕ|=[-�`G �0��m�� s�� [7 ��'qO��"ŬT����3z�c�t�rk+ �)T� �:�P�:r]�M٭���(�{<:�V�Wbŧ\���{T?�Og`�z��s���_J�y5�ydYG]��]:�
\m��S�Q����h�r���ڕ"�u��ھzŎ��oF��_]��H�)555f gB�����IZ��={r0Wv
r���0���N��Q-�o�g�;q`������ࣞ�>��M<(��0�����<�P��n|l���n/e�l~�؄a���[�s͡�2�ş#��{�^�I�k{��U��w��a�%eki:�rv���O�)B{��;�t����;N�.(��{�P�M.&�<�n^�wn�mҢ��H'���Z�1�oǺ٘��x�uY�+��%գ�B�%�v����	m׻�Eh�7�@{�x*O��2�׆d��0�g~o��r�l��S���ƺ���H�0������)iw��r��"��37�`��K�\<�Љ'��%��ᙂ�� ��e�k����I��v]¼8k�[��W]ea�Ek���=��:��]i~ss>�(��l�Z�˱8��{�7���V��~�b��eu� n-�쓨w�uW"�U�K���w�0�;:�p��h�r;X���r����7���zK|o���zV؆Ǘj�0�,���v�&�g��>m��^�[��7z��iY��������lh^c�m6d.��F�fKd䋻v�=ϒ/�n�v+�������3pM.'������@tW�}#�s��M�v
�.~�҅A:o9���+D�2�>D{�x�E)l`�uok����ؽ��ʀ0�n;Γ2�VX]��Cܗ�mT6+���!�1�:�_�����`�7� �.�z��k=��{^KP��`�xާ�h�IxY�)�u}'�U��n67��\�ed.��8W���Fn��w5���榺��*��ǅ���:v���O��&y�BxC���x��1v��WѸ�g$�a�b)�{e�>cC�cO�(��V��;�S)��_QF��5Mc*����0˻�sg�~���N1<;Ba��c?�
cL(�b\�_�H�E��ݠ��\��N���V�����'�5��@[������>�Z{V䣊�̘!�s�d�����5��{W���E�mg�|~�R���߅�ZKx�$8�x~�?(۹}��l�&}}���syW�:g���Q���b Wʉ{S˨<�;Ͻy�w�5��,BN���7}m�]�<���︨%a$p����:�^�e�a�<~�[�qf*-�fP�kmuV�:��n���/���\90�#�����~4�Uv���N����Jo�����抳:t8���ڬ��:U,�Sm�����&��[B�}��%O�jI�D{����3j�b���h�W�!v�h}�k�0���ujC՟�#d�\Y8`6cX��^.]��<#�������'z�M�o�ζ��l�W�|�kJ��y<�ԧ�9�����=d�屠|l.�z�ΕspR�.�1���7~_U�@K�!������<2㎆���SZSM���0�.;KK8Q�L���C�(��OW�w�jC=dvUc�rTB���梅��=�%R��Cp�y	��l�*��ad��P�ҩ>��	/{�����y.��^\;��g�����Y�8���7�Q�xL�}w}H����幝�v����)ٓ)@*|=1 ��b6h��V�\�xc��M?m�F1l�oT���ʄ��w$�<��ْl��)p��~w����b���툋�+:GG�N�]�sC|�X��y���u7$�溄Qh^ӿ�\�B�m��Fh��<G��lp��;�ң#]�֪��^�=�͏sI���͏Udu���Kλ��g)����S!xF_��}�j�qѮ�]n�s��@��E�0��ڱw�кؚ^�v<�`S L�r`u)�8�0�9����ׁA��1��᧰�V.}AV��ji��%7\�}��{���L �a�؄����Q���y�#�v�ھ��l�]#���h�xp���{�,�t
w
�����B����Q�m.�ö㚗<H�'�5�oգh�!s�O^VI���0�ӛݭ�t2ƕBvp��k���>�+�dRk��U��A�f0�5k�k%n���J��rL��3�� �i�(�D�-��mqW���|���ja{���rSZO�Fx��>�G}}"5sa����*�/�%��J��EL��C�_K�Q��e�K��G�l���I<+�*��D��ǜ���nz��S���HqۡC��@�&Zot�
��O��S�`u<g�Nv�jw��n���WT~b#�&�mS C�Rt��x��G3f�}KBqF�����������v��nU��S�a�`x�=&&�vW�ǆu��6��;bvV��}+if�D�p��y�"�񾩲�h2������mA�|׮�(�#����˔T�/1�K��3z��rÈu.44=t�6�w�1�7Kj�gkK���Äʥo��&���z?~���ļ:̤k�?�Ck�CL���v6�a�ʭ����s8�x :��l��ޙY�ܢC�a�e��w���}s;��k6����/�Y�Y�̣�Ø�������Q�?�p��ٜS�⏱�qc��r����\�ӹ[|����8ē��w=އ*�P��h�0�{�d��{x��ǜ�L��2.�/�rj�����c��Y\��(Ԓ[���*� 1�x��t�K�f����qL]��Z��k�Nτ��C����w���NO�ˍ������2Yv3�v�,�����ǁ�y�JЃ8���Hx�H8�"z5X�ϴ���
�f�Y\5�����C��잺�ԥ�)P!�	�ߠܰ�g�)-.��ܢQ��|�U�x��&��������ӒM�ۼ�f��6u�C�e��wS<e��]j���S<��
�x���轅��Oy*Yۃ]��p�^O[�r�Xt�{W��L�
zz`vZ~��C';�s�k ;��[��na��^����2��n�~�qӍ�m#.�Xg!��T"x�JL��0}��?^�8�џn/R�'������ܣ���:y=�
����f"ʈ�М�5��aƔs�� ���ޞ����y`I������<�S���-�=#�&��:j�#��3��[\K��
 �D	M]�^�B�}o�3��.�᮸S��b����H�&�Zw��.v޾��;�b�$lt0����\H�D9ܫ�w�H��^ҽOT�s1�Λe�^ǵ�J᳨m��x3�Vs�hjW��a�/n�^�����U"Mi�@��X>¸�<�[�O<�Nx�}j�ِ^w[�����>��m��,��:׎n{K�se�8�ֶ��;�xZ٫{PRZp��E�YM���{V��U�v�����n�����d�T�f���e�O܂�r�g����	��ۅp��[���Ӓ��:��2-�-��Wh�L�����=���΢P�:�ƃ	�0�%��@��)>B��g7['].�^��|��#|��"f;�_����`�:^�qR���F����'�o��}k{�ƨ�j��g/����SS>8k.vH��-3s�}� �t�:�!2�i�f����z��|b�W����U��2a\Aw���&q�Ybt��T�q�v}�M��5��z�o:��z�b����o�o�@���δ�����/O�������9Ou��H�Ď��2t���Pfg��\tΟN�|{>�&� �g]��k��0G~���O�FK�U��ve�Hs���a!��t�æ��Y·��ZN+��ݚE��1-���Y[2�-Tѕ��
��8��L���a�fuw,�j�~���j�8��R8׸R����ayҷa@��7́^�.��k�"��zh��s�v��(W_W���&���(��X*�un�C�7�rVٺ�ɸ)G"-���`���K��;��=��󎻸5�=k�&�N�SPu�-i-�$����zW�4|V�!*=�.��u�⤾��XA��\��Q��x#�8~�s����a*b|'���a�ye`5��.��
���^u���0
���t9�M��@�(��T5�-�]���F͸��ʋ����:����p���Z�Zz�^�:��Z������0�v�E��/�u���T���«ZEX�n�"��Õ��J&Ov������-��⾹�U�YŦn���J��o��ާW/"�|4I�{L�kV��s;��ܝ�ݮe��Zb�Lhv߮��4A�G���fc	yf��b�mk��ې_L�2��<|h���v\��"�xh�&�܈��#��<Dy!Ī��X�fu��ݺ��JvS�+Vo�m�c���Q���:a��Ϻ�D�ۙZ��u�;/�8R��V�n̲����'���f�}ț:4TOK7����t7�|;l��
;���٥6&���b\��r�oD(V9�IY�Ŝ�z7��˕0ݸ�)1�o2�(_S�k�c��D��[�&ᛵw6��Q��т�غ��Z��;YX*�"�I"̉��p ]+OЯY�B|"�h[;�Xb&fF�B;T��]��ꟙ����3��3�S�l�<۾Y���la�8�+��'��A��;�j�W�$�Ɋ�B��n��R��[0kݙ�w��Ϗ���J�{^���=�y�~��NB�Yh,�(�XNpG���;[vƬeuK��AZHW-�sg8n�<�N.��ܬ�Z�2�J@��D/Q��-�E��pװ�$��/�M�1�;ss�����<gD�İVl[��A缼��뼖͗�*��o.�ܑ����G�}td4�l�Xb�x �V^�T��^ 4;L�A�b�+���S~z�!��rwfk��[�B�����`du�j��4-�6ԛ�YE�L�ݑ6���j�a�}�{��Lkb�k��]Z"���~�=wL�ܨ�Y����=����� ���ϖ)3�#� ���&�euN�N
[o
�f�0�Xyֺcm�}�����,�b�*�LT8;�8��HϞO�8<7���M�l�=>&�p��ml\���{U �;O8fi�oPz�:�Q��ԄQ7VE%نe�u���y��'_����v.0gϦ<��=ݸ�0�w���
�ߋ�yEm[��D�nd�����R��zL�`�)C+r�:(��tR�*�M�Ch��nE���<('˛%����{>�B��ˋm�U%����0Db�6�F\YC�qV����A�ٗ�󣒰+��s�Z�av�I��p����q�5v���Rq��醎a�>��	Km���GA�R��op�m��H}i�ڤ/�hVn}Z��[��M���٧m>N�w9��uN��{��Ǐ)�hN�9A✵�]&9!��*8Y��6NeВ+քf��kJ���X��԰�rJ�TL���<掬��.�:bQ�t����8�TTN��=A#<�(�����*�d�Ue�u,J�2�dr�u�+吕ܮ�'nK'P�-DPĬ:T��U\�ꨉ�QU(�P%�"s�T�'
B3)5iQ$�N��DUeJ��*b�-VG#�+V�)L�W3� ����dd�u�N��9\I*u#��R�sD��hAgFIJ�)RV�*��]E�T�DL((���ڦ�������+2����D��e���2��-$��.�(���b:��z��I2*9�R)��C����ȕ+s�e���n:�w��3p,m���Ƹ����te�xz�d�k3��kA4w�]��v�����O�WzSF�:s��d:<�e`���X�R�+�4�}ǀ��һ���y��G���n='�~|�;�aT�["o��s����	��<'�|q�90��G�~C�}C�B���$�����)����<��ޕ�H��q鏲\ß����il�k���>�v^�~?����99S~/��ސ���{����w���ό~y��]�?�c�C�S{O'B�7������.	�C��{O.?;�97�A����r����$�����xVw�^��3����=k�AV*�W���[AT�?
�;z�|w�yM�	9���������i_�޸	�!8����~�����z<[�ԟ��>{��ɾ�~��J�&~��b/��l�S���棜�~�c�Y�_��|�}Cۏ�&����w�'}M��z߾v��yL*��{NM�	����Ϗ?�����q��|��|O.ӧ}z�����o��ܮ�_cs�u�0�S۷|C-a��!Oީ�MRⵕ?:�>_=�|��>���o�ݿ<�����P������O�=���90�ӏ?~���n};�a}��<`Dߟ��}����	�����<��rs��|��]�r|C�O}��_>��|?~{���^<�����yT?�I�?x�(yL/�?���ޓH����i���<�~BC�5ԇ����������xpr�_��񼸟����_���Cۺfc�߸�d��3�v���.4/Tĺl����9/�c�>��>�#���ULcۿ����7;���{N��©�'�W�?��L/������{��<�{���S|BN|!�֓}Bq8��|x I�!'���o.<����xC��}^����cݹp�_?�LD	�=?}��7?i7!}���Ӽ+�w�}C����q�r\{y7�}<{��aw���>��~��®�|���S{BM���q�C��G�}��NӤ�>o�ϝ��߯?�?=��ϴ��8�9���������￻zL,��������?�O;��6���ӏ?/HxNv�y]�������s���`�������<{�)���Xj��_xX�������
��{/���}y���7�ӹ�{���,��������N�㓝��.��r!��w�¨|q'�����=&���?�bW{M;y>^�����۽8�P���k�<�-�7�'~Kc{��?��/���[���2Л]f�2�Am$	��Z� �}M�#WȺ���ě�%k*m��~Q�w�7ؽ�zh�AƬ�ME�&�om��,�B�\������F�\�R��.�eo[�7ݬ,�l�K�x�e��K�G�={�w�?>|���Ӄ���q�����0��=x>�zI�w�v���ߝ���zq������P���{N~����w�>;������yL.�;xC����~8�]����1��<|/��'^{������u�ǯ��@���?x�|p(q�����7����o�?�^on�������������6�|�����o��w���}�9���5?}�L}�U��a'��~���ߏ��۹ސ������rohHx�/�o����ϛy@�������s��!�������cϯ��I����o�|�=~��n@����9��;�؏�g��LW���}jl][�(�+�o=�t�g���1\���Oq�B>�11��_ݷ���0�����}|��HI�M���ǉw�i�q�>��<��NC�4���}����粘\|q\q��ɏ�g�}���:-?W�7��ǿ_�~w������i����i<!�4�On>��)�	���}��ɏ)�!;���6��x�!�?�AΜ}~�<�s�;I!�ܯ����<&��S�|u�՟Y�c���!�~h2;B��c�y������>��L.���O�~p~C�aC�{�����H}O�s�����q ���7z���xM���}~��뷤��'���ǔ�$�S��q?~�'�׋)��O��z��xv�~����꼿����z����~�~�-����)����;�^���P����~���<�xC�x��ɾ~���x��M�	=}��xy��r__��xǤ	;y޾����������9T�}HUp������K+]��X����?���������O���>��܁�<���.�Y����u��xO���;��}B�y���������7�~��_�޿G���_|x=�x�����<F�������������w�Ş�z������[��K1(� Q��?ր�n��'�z<^��\{O;ռ~��ra�y��|q�]�4�;����<��4�O��xM�	�<��/1�7�'�������������8��|&���߿��c;K�g]�����z O�?|&���F�7!&��c�I�Ƿ��x���{Nq�=o��]���y�����OV?;�������q ���g��z@��oh^���zy��o�N��'�Ж��4S���WgɅ����s4"e6F}
��5bm8�v�ۺn�Ў���i�f�J��ؚ�5����}7ݺ��c$Ia�(K������yۙO{�K�J*��e����[ٳ��N��K�<WkTfH{'��%}�I��Ϟˉ���m��ϟ~NC�i�O��ݷ�];Hx�#�:��\y��}B�m����>�~y=A�=�����o�߽���=���}������#up1/���)ט��y���^��0��{C�����q��N?o�����M������
aW{Mx>���ސ��_��}��yC�4�П��v�����x�	��'�o�[�v7�'Ӽ���y�S��ǎy��ߟ߿~�78����@�?}�E���ޫ��?|<#�6�	��+����������&�����=��9�\rw���xt�ry�޼�90�}��)�!�����9T?�^X�!�4�'��G�w�~��}��ߟ��~{��&�BC�|C�S�M�߽^���89�|�������ߜo��$��׾�����!*��&�S�{q<���C�s�>�x��|	��]��(� Q*��^?Z�x��>{����7���Ӥ='�9ߏ��Aw���x��~I7���<'��ۓ~B}c�<+�w���}Bq8��=����zM |������"��|�������������7���^ퟞ����3�-�[�W�s��@��?F��1�>�&��M<���9���c���I���L?`?'�ˎ@���G�����C�{���0�������o(ra�}��~v��o���~�_>��	=g�mt�}c&&~����g�G�DyM�	>;z�󼫁M�	���m'�ۂC����;x���-���}��𞷋�aW'o{;˾�L���(|O�s�����׃�aw�~C�W��OUCd��9�OkoV�����|	$~�����roG���>��w�?�������}x������7�$?����U����t�u��ׄ=��8��|'�0��I��]�S~BV>���*��<��3�Y����1�銟�����ǧ��?''���ߝ�=&~O�?;�S�������M�������q ������v��$׸99��ɿ'�9Ӵ��	��>���?@�C�\�p��Hy��ʩ^f���s���M'����E�oޯ	��~���+����4��=���s��!��O�x��M�>�&��|i7��o����׾Wo�x�����0�]�~�^(~|O�S`z��p������������t��rh���%-���[0�Lf���
V����rݜ/��Ť���NW&�4<��P�L/5�WBn`�W��2��ρ�zX�ʅ����y�ˏ���vp�8p�l:Б靝�S9�*�C]%l��܀�6���HJ�\.������Ϟ�l�ý��s����(xL*���y����P�'G?�|��7?�m�<"�����}�yM�	>�����Ҹ��������OA�?&��v�"������~����>r���oD��XS��������_���Ϟ=��aWeǏ~���0�֭���w��x���;�yޣ�}C�������O�zC�;O�>8�w���RC�G�����]�7�'�?y��7�T�P������so��l��f�*�󍘁?9��A�}����=��8����ޓ�;I����w�iP��97�����z�o������'���I�0�ǟ��i�q�ĩ�:C�?�޾q�0�\H/~�֩V���|1i����GML}�`Oޏ~���P����nM����N%}�y>�}BI~y�yۓ��C�����iHx�e7�/v�y\
o�^���ɼ�bC��τ���s�&+���������쿝�����������N���e	�������]��� {>�����:w��n�y�����Uދ���wF�97���Nv�8�@��.ߙ=חi7�$��������?�(��w�vjy�����1���_(�������>&����<'�����^�N��U�����i��L>O~�y���'�9��{�I�0�˿}��r��#�	ğ�#Tn��;(~ڎ���?Bv���T�uE�+�n�����$>'��_��v������ךp)�����]���<�~x�SU���{���L.��?x<��ޕ7�%~~���{Nq�����y}8+�o���������(j�|����h�R�{NL>����_�>?�7z�~|��������q��f<z�\ͪ-P��z��dczNh��"qi�Ĳ瞶�|��1Z�$t>���T�\�y�2����Ξ""���{n-l��Z��a�gM�'��ک�.���ݪ���i8 F�:�xb�K�D�f1�ov�)�q��C��̌Z(�Y=\w3�,���м:XxzP���85M���qa^y;�V_�x9$6�Tt
0�p�MPU}���JTx�d�Ijo�}�k� z���3^��}	�Ꮔ��%gE�w�kn�g5����e=�M�(J˫Rvu�ȺP.���E�̦�n� rgsy�0���%WJ������F5q�:|'m�]�D�%�+s�OW_�/א���k6g��L]���TЇ"&:�����{�r�M������P�t[�e\�G����b7y� ��P�kG
��ʮl���42s�J�CE�L����r�i��v�}ŔS�W�c�u=R�h���j�BɮK��Ƿ+^
O��!7������0�R�My���vak^t�:������,���~mRZ[��}h���!/Į5p�Աp;'b��w���O=7��f�Pk�e']>��Xd��>(�6���f�Onbě[�%y��쇮��7�̯��MM��G1p��H��I#�e�7�e��uL��f m�G���'V�u_k�C	�洫	ĎCt`�_&/�o��uX�����x������RU�u�x�U���#*n�y�VG���"���ɗ�=Lﺟ���Ѩ,|ظWFY���qZ>`[���ٹ|�]%�S�Bb��w��c���G Φg��R��G�Xq���P�K��[/D�w	0n�<�=�xoY�,����=�����x�a������T��wc��(L#0�I�\
(��iOk3mp$���OQ�QC��wa�LXt�ד���Y�|�c��ۑ����b�q�+��I�ŷڼ��Z��޴L�y'����Uo������[Z,[��C����{�����]���+����5��aG�뾖[�����󺥹���h�A><7��``�΁���:^���V+��&-�G��^�p�ԙ���%���7w�����U�L��҆��ă��@Xu[�[TY�5X��,{P��ftj��G���$n#Xϸ)��� �8�v����'�b�ٍ�}CI�U�$2�+E�"k��k��6�٨CK1�(�=���ؓ�!�;l.0pjx�ϲ� \9���V��]���{Ơ�Ϫ�P������N��&�V|�0f�b����顙��	�<�=�ҍM��	����1�>�־��.4D��wl�[�$pB�e	�*�����y$��3�¡�H�{�έ��SBZuܿXW�LӢ�$˯�B��K�b��`qO7�]�uggt�Q�s��j��[l��N���qz�)�괙-�-�!;n�zK�4v�H��z��bX�;�֩�pL	�AC٬�,�R[��*v)J��OX�\R��FpY��u���E�Ml�4zT�*�vfe�5����*�ڦA,���,�"ۧS�����.�:�?j�M��ά��i<'�\WX��/Hss�.�΅D'�]&��0:@ �0$;T�׈�Nҵ+��P�uZ��	'm���r�,ec~��+Fdm&,��Q��Yϔ���zѫwn�%�g�p#Ԩ��t�Ǐ �d���\�y��x�s��J�r���]*�.�����g%��V��,m>�	�v�<�@�M�W���
}B�c�wp�y��(��[�a�Ѯ��ʇ\��=N'll�4A��IvEvʷ�~u<�Vë��\���i_(�:/�a;���g*#����3�[�q, ��K���S�E�n�,�z'p��Y�g���u�ˍ��UƠV��s����5	�a�J��GI��=��RD���R/��Zz�+��,;>n�W�mq�����	/Zig�Q�cW�}G��xr�2�/er��>^�jLGJ�ӞVF�C^Y��vzV>�K��<!:���x^{�Rj3�WDּ�wn4�{Շ�R%������\"����;�g���f�s7�n��ο��t��Ե�盞�2�g�*�B8Q��w�A����t5��W�WY#��b�f��5;4Tҹ1hgJ�M{/�(b7O����S�h�6o�-zu��:�~��-���Dl����|�R����w��*��}��q�
���2��|3x��5���=o;j¶tWG0<E^&�l���i���hz�C}t�u�G�B��`|$*,��=�1gfL�#p)2����"�����츩��ͬL�^�� +e��朰3�]����37`�>͓/��r��v'��d��v��R���r@U�܀Zʰ3�W���(8C�\qͦ�FY��,Fz.a�ڞ
+�9�#.\���j�i��z{ǱS\�(����E5�I�;y|o�F��A�\=ƥ_ 5֮�@�y�2����P�-gb��%j�w*{��X���c�����P��}vo�.�Z�w����Z_�m�uuV������ON�̲�]�6��5s�i$;�9o�P�`z�BΙ�>C<S>��������/t�� *F��=Ż��>�9aҧ�v�v��FʈB	zw>H�炥��x��xf\���~c�|&�����7�e�"ܯ�>�E���;���OXs�q" �;�򯝽��fF*�~e>o���c��40��(=�<��lvL�+��m$��¼8`G&���ϣ�.��b�����cՍU���J����73��U���=�Mz���$��G��uF��Ʒj�sT/�,�.6c�!��(�R��nCM�e.{z
xq��gJę��?��i��}�� ��u�ќDI���w�[*��܎qٮ��[�7޼u�҃��Z9�?r��ׂ*j�m8�nCP�Vq0;;h�G��G��D���� bg���(���f���w
���ɿ�d�:������+6�ʅ�`񣽧�$p������B��W�!�Pg>SS>b���;jɟGH�l*�9$�Tk���ٯ����~��~��U�a����u�@�Z�O<�|/�,���7N��3�w�dc���^��G^x)}��<3p/��t�K��Q��n����H�Rs!���{�ո}U�p�����,�B�P��q�:};mr�h��<V�TM�Kzt��4�׳\zɀ9�ٷ|�:C���~3L�^�.�mh�A�=�z��-<Ù������Kx�^�� ��[�,��#�}T%�l��@�1<;A���XҖ�k�)vgs1yu�p������,�w��,� �%cˢ{��"/Ҵ�����#�����cd�М.��������2߅�ZKx���}}(k�9޷�*P�ߺ�\��*��׭c�l�5#�L�TlIqx<�
��oS�c����+��`��t����-Û�+��^�^~�B]�m���W�-�x��z;�L��!�X��ڋ4I.��t�����05�~!���J�/{�Ӥ�W�<2��P�B�.�y�V�.@:���Y�wt��&�\��.����Y����~����2���+���r:�S�>���YT:(�i]��q$X��F�t�u/U3�XA3 nWUPU~���w*�ܓ���f�n�	��U�����ƥ.V�ݮ�DK�4�qt�3}Q1���O�K�c��wZf��b�u!vP��o�e���wL�-���צ��ށ�M�Ԕ�]���*�N��,av=P�+�(�&f��ԡ�2�������=�p�����A"ܿ���Q�Wy"�gV���Y�<BY��= ��!�H���{�w2���=z��F�x��*@�^�����@����K�~ߊ�{�W��G~��y��9gy�Ոm8V�f��a�@��<�X8��mQ����z�!$Ϣ���i�~C8,f�t���{���sj�n�1A���X����`�X|����ഄt�ǁ��:Y��?g�7��v}*��U+1ƌo[?r�nC�h=Dv����8�ȱb���ۏ}��{e��w�@r7�hz�,��V9Y���}T(�9S��J����9ة;��t ���z�������ʘ�ō�;��w+޵
(r�x�Hn_�,Z�n �}p{���</<Ǆє��25�{��*�}7<��s�Ca5x�{�8�;k��vC��t�D��])Űh>�V�� ���-�=����k7��kV�ʡ�!���]e��
W�kF�jގ捴)��g *5\�o+�y�ʤB޼��OM�'�2�2 \��뗇)�&�������f겔$���v�����t�x@��y7��x����vN�xK�F���:E������XeB��g��.����Iʾ .3-<�D_·�lY���P40�:��Cj�������om�G$����q�=]���!{�2��}A�����n"�[}����d�i�����M�}g����j�k�{ې<.u��.j�+�?{N��,���5�Q�:r����K�k��{:>Tq�)�:QӨ���w�]ODǜ��DW���+���k� �Bps�}=8���w�1��,�|{,aJ�AjtQ�'hPf�����t�r}�ch﷋0���uip>�>컝/A�ѯ��6��w��[�ʷ��F��<����
�2���_2��������8t��!G�����b��(.�[�Z���q�v2���Y0c�S�+�#����(�]�(�\YGm�;e�u���s�V��ڼ��膳�CC�,�烱r��^
q����b,::��o,���w�LP�m)s�:���;�+#�s��l]m�!��Q[��8�[;^7}a7�h=i'3C�-��t�4����B�־�])��AZ0��>ފ���eL�w�ͤ���ǎ^���m�c��3��*�Xr�Ƀv��j����$'݇�04Ջ¨�ﷁ0�;FZ[��J=���c�j�a������"�>����������643�c�N����ws)l������e����.���[u�Ղ�"�k��!�_t&�h+�3k&�aY�"r)�M [�q�w�	(��,R�o@8H��&��;���O�[gXX��=��M�Ep�jK�&�"�&������f�(�M��G�ȱ��p\��u������D`(li��7��Ͳ�7��=�4q���,w�c�jT��s�6�oV�΋{�S�l����f�S" �o��G\Ps"ȅ�ks���˃��Qr	�|��0Z9޽����z�EMLF����2l�i�k1@&vh�W]M�m�4�u9����g�^b-��B	��T�΢�VH����c����3z�2E��ܦ��V��1fۆ�D�A��O�Z�V�@Qr�3�c������Z;���]f�����=��ъ�]H.�ʾ$�ܘ&�&�f�I4�+K����-m�	�]��/N�X�����g�:Z��v2��4�%]E���+���3��c�6$d���v���b��D�ʟ7���Ұ�7�(����Kn�
��_?����T�Q&�I�� �5�|��E���+%QZgI5iQE�EzМ����b��0���C�zUE"�Kj�'-tND��4���s'$�rpu#Α���^��Z�b��U9�(41$����DW$�^�*�H�څ:�EgN�(�b�;�QED�/v�2.�d�%WG'Qb I���3���
Ye["�ı
B�R��i�ܒe��Ad���)�.�20��t�#��lKB��7W0�I �S<��<�OQ�Z9�`DET�h%���V�D�˺H�	E���Eҷs����pQ"�9�u���5(4(�E��fJ�0�I$3)R�t�",�8i&����"����ە��*�+��J�r���$��#�̣��Ј�NF;�l�u<wn�#��a�*�!�ͬ��8eW*$Ú��(*��Rk3+�fB(Z�'=E4DMjF ������ɹ��ި�^�����ꗆ�+W94�Q�*t/7���ߛV�R�g�?r���Y����.}�-S�­CgP�eEO���ﾠ�E���C`��X�kє���@�˪��5���xb�;��*����S�t-�6Uօ��p��Ҷg��:�!"�/�~��A�������e�+�W���^�'�]�3*�/��ݧ�K���� �;��<K�M4�n	�GM��C~������ZKB�:��Ƹɬ�hI|�5���>����5���N_r�JD8��/��:��$��ܘ�CA;�t��%7�Y��(���3ؽ�N&2I�^U����G�t�4r�f�d��M<��}s�r�Η%>�!ۡBK�y��p�+�ܙ������|ת]W�(�nWk�u��:��.xl����� ~��q���u��ک�^×CW���wS�m����NX�u��uu��>4p�b+�\�iI=Sk�xe�щ�)��ik:�)NV�fG����Q�D�����g�	RR�,$�炯�ٻa�=�|{���;򧝙gD����%B��)3�.�Me�9=�0�f̯��\,��$��"%���X����&)�g\<M(�R�%�v��NL��e0]p�vY'�6&L�>CZ[���&#b�+z�Fe�s�ֳ��#��<|���{}�;:�>Ӛ�㫮���}�����`��z?3p�Y̹��+��h�*Eowo��X���hK��G���
�����s�6Wu^˽;Y��¡�"6a�w�pbp8�����[��;�z�b��O>��H3���+~*��\^��!�]ڼJ�Js]#���$��X�lT[�D/��W�&D�
��W����I�ç���;�겨�v���3�C��p�ɋ1A^�5�Uއ�)��8.��+�Wx����D�����ײܥQ_vQ:�������_,�,3�r��
y��M7ǳh�U�I�v�ߨV?muA�.Vt2_o{���Q���D�j�1���:HGe�s�k�����]�g�U��'B�.�9�:���o�{Q��7����p���3��Ȱ���}6�\�ye&��K��qNS:i�L{�6�ۏ}d�6��:'��i�nzD'ϝ���N�/��߷9���[�F\*�L����Z��.ŉЇ��~�?/q�xS�[����k]��d�A�ej�k�zeY�i�|�:o��ce�? �F��.��3a;�W�DN�f۴BP�c.]YQeأƗ�_���
!t\���ͬ<OA���M�u��z�q��[c`O�>��^���H�N���U�"�o_�R���b,���9���I���>�W�
u�O�͏��<4���#���qƭ�U}_UU�3�|���,����٥��K�\��GJ�q��ު%��(*ޛ�/��>'+�k�e�x���:�zA�Q�p�N�E�J�H�|�a'��P��DPTk�5��߾�v}ڔ��U�3��"�S��4�u
9��|5ݞ}D�N��$��rZ��]T27Z�+���+G������N�xaI�^��o��~B���h0�����1���W��7�T�i�I�S3�����=��U��n�::^�q�ѽ�Ҷ�yp��V�Qi��Z���
�o�n�?��XVoy^�^��d[��\��˿.g
�����A���#�WXY�#�}���*��s�y�+��5�w`y����$��M�o<~8ݰ�(n�4zb�_N����&�I�-���M%��˿M����-��m�Ǔ<�ic���B�m���gM�7-j�D�-�k��}-֜�ok�5�8|WK�'�؛�M}�:/�~3P�/*E�>�CM����a���	����7[�ۍa���8ewul�2&��C����*�@����2^ػ��Y�����A�`�ã�{�փ�=w�:i���}��1��`ԩ�k�%�{sx�|���¡��Q���Vnk�1��X1f�o&�2�4���
����l��w�e�B�5 ���
�J��E��r�TŔ��y�,�̇��ad��!6�{��6'R��&�����= �h�N�T�HgRcˣ�������</#$�倯s_N�������ոr�s�9ձ{��T�߅�Z�?-	3�n��Fo�l�ܐ\v��`�
��Y���7�XQ�r��!����k/���Osp��ng�U]�3��o��"sVd_�����+�]��/V���E��tl�N��\4R$�*^W�)�q@�7������}]O`*E���G8��d~��%we���#�P;NF5�ȺlX4	�P����zE��2�C�}X�"���3�N�����Wӑ�5h�!ѴR�����ўl��ä�H�:M�l��X�|1��p�xxy�8��αx��~is�RO3��C���W�p�>����k ��l�G��X���u��?l���<[����'�|�b+܍�&�㧥R{K����,YF���z�h&�p�����K�l�w�-�͆ױ��&��Y�^U�>{]��;��^=h��F&"���Ǣ����� �h�����t��YD�y���6���j���GNt�޲���o'\���;��?����#�|O^&�Eu�tdzf��?x��|�M��mWhc� �sJ�\H[�#
Ct�����d�%��Qů�U��:���8lw�b�>�h����jm-s�t�Mw&-���=��r#:��jv�3�1&~�y�(�ɍ��F������4���îAi�c�b��U���V����P�N�ҕ2�d:��0�"���	�[�,|{6:�s��y����A[��(%�\U��į�����[�:P��?u�
�iz��N���mp�]��H�a��!��@���|:��L����YD�mᬂ:�4����ߒ�^|��~�vKVc���J�Sn����.��]V�˯�B��A��[�W<9����;��.-="(2�g�u��������O>���ZPP�T'��&{/j�fI5�3ˊ�z�Sp~�˹|Ԯ��9H�k�	9^�e��%PE�+�%qG��ò�s�i;�H9>�F�u9�^��;���5�c|��V%P�8��Z�!o\�@�t"�f_��v�� �i8O�r�P����p�J�C��g,s�g��v��冺�)�(��)�]'�Y��bɑ����Dե���.Ow���o�,v�ga*:��^4�����>��"@w�he�I:������%�77ѣ�v���ҹ�qW+�o.WE��z��L��ڊͧ�:gd�o�JW�����కݼ�I�0ݥ��j��o�R|�N���=dQ!�[�lc�wp����y/��St����fӜ�����Y�WT�F&�̷�x�#�U�Oa�(�[�?9刿U�@�$���v�k[�كN9��ߕ�8�虼�}�%��.CL�yW�E�L�@о�U��5�e���>Y�!�*�X�xF�r�Y,��P��8F��!I�裑tx�2�o�,����z|�xI��X�O���+�UJ�I�0Iz�I�uv�j�V%æ<�nUG�����S�ŪjԆeeØ���T7��g?��'_�<�w�qS�;b�9=jtp�n��qg��I�f�3�����G�_�*�p�'g��J�!�v�����Hk�l/}��Rp�0�gf�r��îe����Cن�^�<Fت+�3c�X��^�	�3k�����8�w���l��͓Ӗ��9Sn�<�b3�Z��AՈ��R����ez���������\�c&
�������M��ˇO����Z�Df�&�x
\/Yͫ�~����T�qʖގ��aWQ�$�+���&���C��@�P.;&���}j�iW�4�̷�&����ݹ����Ϭ�+�����r���v�w"
��er��D׫�p%jS�q��XܝCf��9.�]��#��" 7i��%&��ޯ}cI�v!��D��f��c��	���>T�Y�L�S�!������.�,�����U�F�
Ў�3e>�?�.,z��tOXO�����m�2��*�b]�/5����G}ZF���&q��P����`%�v,Z�C��.�;�,�5]�X���13�9=����HK=��է�}V@_S���[Y�(t�[HYw�,�Q�d�ME��s�<���C�S�#�Xx���\��w��O�{MĀ�.�x/�n>����Wi�w%�݆�ti�0a9��ol��:vH��a%���6�"!��Z�ox+����_V���eq�<�*��Ƈ��<�i�tH��jӝD�R^��x�%m����f^�/{�-%���,S�R�p�-����j�aI��}���¥�/� ��R/�)�����Sc'��^�	�+�9YL�3���qS�]p�k��s9`�3k�F�<���Ǻ��y̸5yi�>�!�3ב��h������²����zĽ���A�U+n$��݄	�1�I-ι�E���8�޸�K�ZQ�=��ŀ������l2�}b�N�ǒr,]q�ޟ"�f�@���n�u�r{�UѺ��|��Zn�*8� ��WKA��'u"y�,�]���*�9�\�nb�Ԥ"�X�o^��j��J����f]���T�_}���UǼ�ԗ��7�q>{�(_�P[����; P_�af�.�3Dd�d��YX��]��k���95۵���q/|��G�#�Z,g�C���'�8��]A�W<I���(�z֓8�'�1�l�<�U�%=9f���q���sz�.�}��|�����؎�2�%�%�\�J��B>�b�t�0{�\�kG�6���(��(��>�y��)ߓ˂�k��+h�.��kzR��Ⱦ�FN��O��L[����^a8q+�[Y:5��/�/�vPdk	�ж�ު�� �$g�Yڌ�%k�'Ft�b�V�]'�{U�jZ���c�#>L�s�`�g����뾴-t���c:�x�M#�4OYqQ��+5"#����Ļ��"m[��ζQ��àn�ؒ��xQ�i�r{��#<�G���~���.���*�˅�y�&�{!g����D2n��R�t�l8,d~�ŽX��pu��음������J�Y�8�Q!�o8��u�}*��K��z�:��͛/;|Lf'LEi���B�X Q���բ'.�U|����i�Ǖ,83��[�p�b��4�8��/�n�蚺�0�`7��{��N�/Sx쭜I�鹱u�n���'�u�9oG(��u���qvm�������
��}����C��h(��;>Q�S�Ds5�~Uw�<v�	��5���������^i^����[��U��6�_۶��"iv/}Hi��n�e����b9C�����C9zs�q��4g;��Z%��e&a�=B�Ge!����"q���F��bfX!�4�G0��j����[�*�r�L�P��Jo#x������=v�Vy2%�p�[p�eZg�9gV�R�c4�_��6Ӌ���%��Q/%�{���ą�܀��b6k�z�$l��7u���f��G�O�i�������@dZ�;�js�!��+�,>��(��u���廇/ޯje
a�#!�,V#G2��NJ��5J�7���+�%ȟ+���4m#[Nf�oq�ާf1�϶�0En���9�E^��=�x֎��m��	��en�瓛7�e�3#��7��Za��wX�I�Q}��?M[\.�5���`�
V��2�p���<�N�yj�q¤\��JrN8��:s���PA��T�H�_3Z����j�X@�x��9*ur�8���*��m[��z]�S5�j��uK���t�r���Y|e���$�J��}Y+/I��{[�����{eg��������+汷�����:�__\)j�O6Sf>�h�6�adI˒pC���"��m�G�����پpn��g���,�j~Sp^�3)�t�{4�nCH���f�Ɂ�����7]��<�~�T�����Y�|_(U��)����c˹}:�ܳ�)���d�e���Sj#�J�����s���u�{�	�~�D�9 �{��i����1[|��U1�mV�`�`��(JsO�e� �Sh�雾��e!�PC�}���p�J�C�,��͕=Y��I�B�i�Tڴ�4g��T?�`�TU�G&n+"08+�أm�`EE����T�u'�d���C�yή�╛�"�_x�t~ȵ:3���d�XG��kJ�T�O
���[��c��%x�Q�a�wy�n��FL:��T씈�*D�;&v �}�	> ��K���gr�G�����Б���Պd��^��7�'����qnXqzM�C�]����2U	����|���]��nO]dpc�]�8J#�!I���g+ok6�O���!Z�a�w�4�9G��>�ܛ�qm{�.�ֻ!�dFV&�1�E�o��LV�ࡺ��7���^�zW�O���dzRki'/�{e^��"�t+*�R1�b��h���K��\�w�0�1|����w���ܝf�=nsc�J���J�(�h�7��Y��u'c�z�eĜ�܇^��	d<�U���]wS Wn�Ҋ����#��=��oW7�ɭ����]�'�{�8�:�P�ots&X�<p���ʥCMZs{u֢�:l�@a�����]v<������1lB*��H{fs���Ý�zՐZ�ׄ}@�u�g�e��3����ܬ6]��B#&x��E���w4/7z�p_5����1-�hC��Eb�ׁ��h4����2�1м漧/�Hf+���4�.�����m�-�M�z5�v��Z�Ѭ.��^Q�m�v3z�OwF�� iNq	�ؖ��d����<���
���� �v�[J]�c�G�N��M��Ŀ8��{�l}	�+��=b��\�؄:�0��f��t�|eU���z��
wr��Rͱm��Ï+*����V6w1e��B���6	Kz��Va�܍�N�q�rC�ӓ+3
.���v'����;8Ywǂݍ:8l�ӣ�DD�[�gs ŵ�d�ǃ���� �[D�w"�9[x����^�*2Жh�"�y'b�`���wUu�x����n����ܟE�*��(U���ʹ2w���5y��G�<�2�S`����쥥ak�,�GS��2�)���&MK�"�u>�c)]͹�#9�L���8�F
�3"+{aY�0�x����x� u<�qޝ��a��� ��n��W�7�
���V�Ѹ��u�xu;�0ۧq��+��S���s�;"���!��AZ�V���{+M�b�l	1�� C�\��.ە��if�7�x�U�^���ǵm??f_p�o��G-@&�P�:�'|И�uVĮyLĕ�j%<�Z텘m�4�"�S'��U��9V��4$��i-�n��8LK�ܴ�x1ó; ��F-Ea�*�5�.h�c�еw�n��������|�GE �`�����B۩Q:�k���]]ظ�{�����C��1�����#�i$���Gm�6�J-����rRsI�q���f�j��C3�-b�v�)�*����m�؈���1�lna�2�H,�,���I��݁���X:��
]9�@7]H^��{�M=��v��?,�xU�ntu{� n�(�o4��fs�b�>i�we*���a����ѵ��1� ]��)Z[2�;P���{��!l��<� *��
d�S��n�}h�J��nc�2�a��3Ze;����WҜee�E�<?�X���Y�"�4�w�\~���}|�|x���G�*3,�NT��&��a!���Ȉ*�A�O*�JK��ST�8a(UA�*�)D����]���,$��FВT�H�D
C����L��^����B�,B��MP�'t!�C
��nXU�l嚄�99DN\��s\���a�F!E�"P�12	6f�s�D��b%��V.��t�qD��Y*���Z���9����Q%P�(D�HN�48b�:�r�FI仮�j�E��6D��YUJ�dI�k]�5�#jIY��2"���:nxyb�"�uʀ��L2��ꉊ�{q�T�%Ĳ�ұe�5J��8^b���
T�K���I���QF���=YT�bD:W���T�AHB�JP�U�"I�N��e�hwv��"�N��9�2Q6���L����#wGJT��N��hI�s$��tHԨ����,M0��ܗR����6$ee�v����Urw���D��k}�8X�,.Ĳ�8��c��[�N��]��vo���_)�̫/z�QJ�e�\�8���b]�c�?��U}�PK_C��l�,)��ꩾ}t��b���Hd���\"���*ү^��]���9ZY�}��;m"����9:\ ����ߜ�q쏼��0�k�b�8���8��F��fa�,_N�|�p��$���P�F�v�(�,3�ˇ����M7ǳEW+��uUH髹��dj��։���S�*�9����:�MY��C��u7�?o��ն�~-��\5�Tfv%���x������йbc˚~L�\�αr�Xt�{W��L�+��;By�%Խ·�i�oO�۳�Hg�'z��-2e��f��;ͮ���++wb��������k���ж(ڷu=�w�%��	�xP����it]�����hy1 S#Nng��������Pm��2�:bu.S�^ [M!�
|����ϭi���jevI����.iDBJ�r�[K���VE�XaO$�zǎ�2{ϩ ;
�&m�b���w�^�� ���m{P�wǬ2-����~�%K$sCĞ�1y��Dt��x\�{�_[׺f'�S��"�7�dZ�p����J�LW\T5T5,�Ǭ�p�/M��n��Q�'��*q�s�����P�q)���v�V�!�1V���䠂�0hJ��0D�+��7�%������㋪1)��p��h7:���l\�l��%���꯾���w:йQS�U-K+?��sO�ҿ�=Rׇ:l{��3Ü�򜉑1᯳A�,�'e�%w9��&xK�4 r�\+C��r���+�O�\0��5p��4�5=�|)��:.շX_E�K���j�oo�yKˈ'mwԟ!k)�Fy=���=�:�U����{����-ү�t�A1����1���q����d8jo��2��mW=g��
�{MM,�0�}��ߵ�_Y#�]�l'%�[�Sy�N�ק�6�&�LvMn�A`k.�2A��c���͛��'D���\Ƹ]h���gVu��Ҥ�����.���{��S��f�,��A���x�4�[��N�Nx�����,�3�a�t7��N[���#5_��:A>+3����~��z�^�c �jTO+j�7��c*���t^�{�<G'M��v���F�3��Wv��Yq�re��W�g�Zik�x	T�o��Z�S�WbY��?=�l��Zgnf4{t�D^&%���g�5��~?@��鞪v��w��h��%�ˢzm��c)m�>/�^|r�vv�:zB��Zi��qtUw�<cpݶ5�#5�1��Aw���2�3pP���֍E4D<)%�̾��SE�es(�O����^�u/ii����_�}��z��I)8M�����{=&s"��˽��:��[�8��2�j�j��W~��������B��O�eLǾ]֦�ƶ�}���5��:�y��s\���2R7}b ���A6��q��z�z�C��d�����~Q��_rsi��GM�n��QX|,_�><q���$�a�L�uZ�#/�M�D��8���\�J�⛗��
��kB���;���*岰pU�%T0����\~_S�ŀ�b���|ؿ���r~uX��(KAlm�v^vf�ۄ�ݾ���y`T&�WL��F�|P,dh���W"u�,MZJ8]v�[�������3�KX���B`�~i����8�1�`����R�=/9[�{��a��Rd���B�e� �d��m��i�K�q]����\'���e�vެ��tl[M�eT��[P�ҩv�aBN�X�����R�MR�X:'��۱DԒ�ϗF�$����0��VwzlgVE�(B̭u|]P�ă���/)�U( r�+x�}�:�W�VXz˯��P���h��QƠ�{S,�����!��2��2��s��Z�v0��`�}<��o��!�S�{S�er�#u�!s��;1���xl�r�w�T6����z+{���zXm/Z��o[޻q��d��ѭ��N3=`Kq�J�K��;y�*s �p��b�8���꯾���z����S�_�X��"�ϗ��:e�U�~�jP��/�/���
8��U�Z�AB�)��J�AF�v�Uws��-�2�A[����� ���.�/����m�w��%�˼�{�W��Ӯ����}�%Ʒ~���7�{����_9uXl�[�$~녺Rn��Ǔ���<�p�b�
L�YA���n;qxc3�.�F`�<����{�r����u��<���\om��6���s|&|\��ҙܛh�`9���Ֆ�r�"����ܞ]���&�	x�Ar�����'�f;�yM��M�"5r�^#���^qU�s�Ѿ����`��'�&OR�ި������S�^�u���1Fh�
�%K�+k�K>>s�6�Ե C�}������ȋF�c�J���=%>U�b}G�l��,�¦���<�\�8��&Q{��Cu����1���L	���7��ƘV����*�lsyG7�gt�O��t�DY�ܿE�Jvc�����~U���>-Wi�m���
��Z��̚nn�6v�YG\c�:dɋ,���p]�G��r,�\*���[��c�O�g�t�h�{���:�U��Y�HN)�]��Jo���3s1�ZKi��w���Y����K�V[�k���d<�<�;3vs��j,���GZ�G}V��=6�F���m}�UW�P}���-\��S�q�]0���ɸ���&��^�{����$A��;�t�2.�zo`�Q�4�w�6�a�0i7���.�8��RL�3ΩE���������V`�>�t�����M�Q�0~��9�ì�F�#��������p��_=uN�;�[����s��Z�wFQ��d��Y͸=T�(>5�	~����-�e|�n������c|���xT��%�.ׯ�8�S7o1R�1�:����xz�T�哆�i�½���U��ZU�/�;�E�K;�����ހ�f�����*r�y��ϣ�&���4�F��]�����>�����'��n|굩�w����{<�g�%�v�C����%{���AjP�ֽ;��c�۝γ[3�M:��Wu�0#�W��Lb���sǬ���\kn��0?�n�@w�K9�:�&�}K���z� ���f�π|���\���r��w�T��3ڲX�Rɣ:����=�l��neת�/�b�M7�D�N�w�笖�=LƄ�@k�=�l��j�Xs�wO=|;��.<�ow��G&��+��c�j=��"�Ä*,�r!L����\o���3p���P/S*v�A{%H��"i���m驹�2�ː���p�9r�ù�(�K�����pX��Ξ�g7�t�wr���P���}��@����m�f��R�1��CM���p�JL�_-b�|���q�P����c�u�l��ܾQ���p���)�-V��0��Y�����g��l�Ӓ�*�E��h�n��u�d�7X�KT�!eS�a;Ht�~#�E���=��	����*�q	>[����]s;�RL�=d�O
۽��w|Xd_��^Ӓ;�/GD�a��'��1y�4���;Ѽ��V"A�?��?��:yb9X{������NōM\�@��
퓈�v�-�^�{��I-<�{�D6l����w��sWJtUo-5��P3���pτ���F�>O�יQ
󝡃]۵=�k�K��� q37�3�V"��܊��4J6m���.g2��K�zc��=��-7���C=b!0T�WZ���nz]�����L�Ԝ�5�6��:u2i3q�;� �N�sæ{�o4ѽ�w��X9tG���C�/�g���e�Ɇv��%(�Y��b\�7Z���kg%}�o��	�
lZ�{h�ޘ[���0Y�A��T�߄%e�� �ɓ,�nP[.�f�u+Y�q]]r�J���`��[���*�Ӧ8B����c8^�-����sՋ�i��=����oHJ��ُ�{�e�M�����&ή��)Q[�C�T�-�_��������lc㹛I�ကd�^����<�E~���Ϻ��}.j�Pfbȃ��N�R�UN�cc�ѣ9/c6��L<V�d�����U4!�:/~pz��l��j�2�=z�N��(f�=�8�3�C=��k��,D��%����K�=�/υ �+� �?H��=�t��w���A�����~��>��8��)ڿ��w�s�l�<�����Ӫ��ǂ�gq����<��:<H�+M��G��>���L����s�լ���πwݑ���tu��r���s%��{�;��Qmff�ο?(�w/�7:�F8t��ѱ%����F�7��ۆ�C���s��8��P[�6���Kk3�w�6o½.�E����+�9�$����q�z�bR�ɏ����&���u\x�(e���kq{N-�O��p��mk���ўQod��&��x׷s�z��K>�Wz�l�D�ߐ�_V<�w�S����0�Y0��v������P辚�/yi.-.�ߩ2�����A��#d��.>� y��R������%�5�����o��7�{�s���հ�Kɝ�ؽ(��H�-O���:��}g�C������֞{9e{C/ݺ^���E��Fb�����b��"+�Y�VsK��'��b	Q�p^�s�2ʙ ���W�}�}��J��Yn���K��5�P�J=b�vR:e�<^Z"o�s]��\4�[<;*.h���Fw��ˎvNC�y��E�	���WN���3a�'\宬q�LXT�j/rʛ;i��p5���������v��-˦VˌE���cz�}7��il�a=����z��l7x�K�6�t����o��.!���h��Þ�!%�}��6��m���"��S��k��˝�Tܻv�K�LeM�ӿU(�j�y�(�ޞ�g��#;t�^�db|R��K *�q��z[���ֽUݝK�WyǸ���z�H'^��W�=��k�{�YP�2�:�WW�f'fn_���>g�ְ��;�7�K�6*�襽�xOڀ�Y��nFk�SNn5�wyξ	��������ӛ�g���ol��@�+��k���
��}3��[�Z�wy��a�I(T���q�Iۧ��f̐,LQ(?:K�5�����9�׍IR������l4�W���(�g�o��,o5��QZ��I�G?-�A>�t�o�I������g�{��'��-z蹖<�a.[��	�u�l@����kA$ȩ�~�����u;zS����z.!� ��[b��O��]���ɝh"�+���fI����Ʊ#�.�Wt�2�fA�}�S�}"��1�1)�ڷ͗8]��4E���zUu��s�OsӁo\[eͬ��fw�5&m欫I�mS��Wv},���\ۖ�Mb?}+������{/�W�ܡ���{.��q�>��~�T2d����fX�G���תo��9ݻ��6f.4�Ug�z�6�yb���g��n������x��jq�xn�ìĝ�1�Ѯs�rI�Ͻ�ђ���r��8�õGAE����뾺�{�N��/�Χ�.,o����[Z=�\t�Gض��~�pwz�u�d���)Nkk}PI�~L����y�ƙڅәaƑ�X��ꒇ���<���]ӣ�Q�S��q76[}��jy�a��_��u�ge�'t��~��݂]es<�e��q�+�\)Pיꄴ�h�m\�Q��usH�.�kNO`��V�^��9ǌ͉Jξ��P5�֤x��OD&��g�rC��v��^�MVC>g9�1�wG�ئ�������w��{C��]`�k-������ f���%h����wJ�oJ�ܪ~�m	׼��fH-5trW��9���b��,���K�Zh>ju�8���~ȦQ�{C�S������YM�=�`�b�T�7�n�o��Ζ��6�OMn����쭺��N#9N�x��vR�vD�޺uR�IM�u�T��E/y[�RD�x��������8״�}=m�E�?��_P��fg^{;7��xL���W3]z�',m�7��}(���e���Rev؎}[,q�l�f��U��r��O0��w	���[0�t����h1���jl���;�6����nU��ܬ��L��I���X�a��c�n��q���z5�3Y�A=�
��h���ǒ�y�:6��޽�����,>����+y+��1�a<�^ ��V�ǳ�dU�<*�s�|xʍ
~;'g_�̚hɼ��=�H�0�Bu��7}�>�H�٦�L��!T^]��T޾�ri��\xl����/�'�����aM��<D�y�H*���7).)��W��=���h�Ӛ5��SK��焫�
X]}QvF7��e�>���5LZ��ʷ��"�����~d�Ǘ-S�Gͤ��:�hDU�B�ecR�f����{��Kk��u+�B��+h��kb�����B9��p�=�AX�8Ȋ��e��;��aL���0T��F�ݽ�81��vr�=iX�ʜ���;v���2yY9C�2u�P�S�)}���}B��+����
ո�r�c:��2��E�S���Lo����]���uA�Ӈ�y�!j�	w���T��+[ �}�oF�]��i���a�R���Λ��^��dA�V��qкQԭ���)u�m5���.��9(��r�e��9�qػ��N�Fe[�|;�����i���;�[�>@�������εCx�Hu*��ub��'`q�y�z�}¹eO�n�F%��ֺ����X�iڗ�7-#{k@�D�u����@2_F�Ǻ #B�i��{qhĨ�ݮ̀J))�>�`�q*��V漭���b
�>!���Ci����Bd��֝�sn�����s+p�@�;�mX�{���l��	�θm�3u�s��e6���L��4.��'��NK7N4�FZ���Yot�l���믞sꇩ���MJy���ld����
�cƊ��dO �2�U�m�_Aͻ�R(	.,��Yxi��sv�ozx�uW>h�߸:�ĕ�ZZY�Pe�xU}��s%�<�{|�Z+�7G_�X�v��1�6�ݻ]���G1��6�_���v�#r�N�1�t�h��0EYcN.��,{7l�68<b,�'�t$��VɼY��jѶ�j�k�8%�m5�L���]�kN�?���I*�lI�4���eX�V�Q��)�1g���������ypW�/2[@���dH�Y�up��c���!��fՃ8ͽ�9o�����}�Z]�{776�[I�tEx'4(�`r;2>��'U����9N��ϻie�th�E�[
��	V t�9m����k/c�W}yϐ�i*
Q���g�ؑ�����on����=F65�����B�g:����яb<%�ޘ��o�`-�S�k�6�}E(Bᬼ�
NĶ�X4,}��&�r�^�ܭ�g;�}Z�Wv�=�DZs)�]Uwj�����A���h!y68cF�%h�!���hp����]�y6%�v_h��p_=�qk�z�s}�'Z�C��)iK�ҟmdHgI�����Bu��-
��1t�RX}�/l��f�t�<�K跢��RR��Y&�����{�����*�̕��Na��cͺ��'�(P؃T�bvv��$�N���/H.��8�,�ß5�(��9t�z� �~y�����B4�.�F�1Gw+��*�LÙ�Es/"��`��U��q�*=B��ᲉNV"l��3� ��H�j痐X�VePG=wD��T����d깈n����˓��:Ȩ'D$��/I��f��6s��-��V�i�GJS�&� �S�GrsM��NE9Q!�4�tI4�*ug��C�&TT��wr�Js�E�ww\wZa��H�9z�S�W��8�&�)�!f!(�����E�L̡�.�r�ut��R�$�2,,HԚNI����I''WD���l���D�jE�*��U1Ն�5R�JIe�/0��f�YQUe�!"�eeEb�d��wC�ʖr���В�4L�A�܈<�%N��&�����Uy˝6��Nazt�*�5�0�%���������B<�.y�!�#�t�D�d��O�����]�E��Ҍ�BB5������� ����n(]vi��~ț�/��),_)�{�`1u����t���&�>��A͕�M��>}���(�Gs��>�g�}_}UT�m�v{P;��z��g��@��÷��_���ǴV* ��IW�xn�"\�e�uv��X�r9�c��8��*#����/i��t���ڝ��C���M�\mN��.��<��y���ˎ3�/��zâN��o��K�!AJ6�=��>�~��X3�곱�[E��ͣ}�5�`��s���;q\� ��#��)�Y�ɽ1��y�}v{�{`(.�Խ�nv �I&ϣ�*��Ρ���y���}�.r�->n�6�C��zn���9;-��{5�}���,R����%EV�UTj���4zK���sG��v��ʶ�z�j�2r7�d�x��^�(�77��۝B��}.7��.ӏv�'p,#1�I=�AKS����騦��AW3����]��S�O:R���n�Hl���&���b�X�c�#S�;k�;�;���[���7F���bx<�մ��	�Mm֏�0L�C�#M\��^�t����[�}�3z�+���SNRμ�����)O��g-O��/ �u)���C{�VGq�^���꠺^˫��t6�/~|Gv��/�=����1=ɟ�)�{ͰvSQu$SN�pw2���rI�Ч~z�Bu�􈥹��K���w��/j��ݗ�?O>쉧س�kÜ�=�٦�'�u��*�MY8��F��\f��6�n���g=$Wbp�ܼ]d�3���{>�f3tv�eV�=閺�d}Jl�v�/�q��:e���=xܵ�nr7fQ�D.���t��/˱_Ʊ�TT.-��w+�!8�j������7���gs�B���q���g+/�>;\mι����k��O/b����_]��¶��KhC�T��i��Oz��T��=�S�����8W�������>J[��C����Ë���S������^ښ�sv�aƴ�ܔ��nZʹ�i��==�����k�����WYV�Ri��|�/i�o%>���/�vB��k&jWWBm�P�\!��^�:e&:9���e���l^Õ��ţA�[y����=���T�wӠ3��h��lR���t���B�=��ecy��y�()WY]x$]�l<�9k�a����}G�_�e��OWv��w��wZ6q�Zm����,[�u�� u@}÷5��F֚�BY8�݆�)��\ny���v<�� ��&{�r���â�m0��}����ᾇe��)�7�=�usg�'$�7_o��q�:C���e=�W�\a�i�ypev>":8�R�R鲹��Q���݋$��W�^ix���>|�*/��n�G鄶��\̯��	��"iN�e��΢�zC�iyW����*ޕ�5\<"�R$.�΢�DR׍��B�$�oj��L�c�V��Q�i�.�وc9��#���TBs�|{5�}�����]^~*���kϨ(�;��vU���L����n\�LNn�N�49�>�<3i�l���|���b�,�u���c��V�J��@��n W�]j7�l�+aG\���]Ł���n\�ps�ǻ�������s�]5W�B/��(t)8��^f����_;^�>�Ӵ��^�2�&�GH��2�u�5R��R�����vq�R4����5#l�u=��K���v����d�w׳'�����1s�ߒ\}|Bz�d�M��a��c�L�������o�2�i��o��
�~��G��"#ܾS��Y��D6�D�I�������c����wj�'-��e����4�k�����]�b���������z-������1�	�o])�*��ӎj�,�tiIK���&͸ל-5oa�����q�]�ajR�:ݥ��þ�z��1땛�wH}4��	\}�&��&{��t�ؐ�T�*��[�	�ʷdbg.��z~Z֘��܋o���d.fp+1�4fַ�����v���zAt�V�g���#,���Z�i5�f;�ys��K+d�:��x,��d����2��m|�l�a
n�7�G�s�$�U��/*�7�)��!�ׯ����}�0f�R�|pyǊ*l"	%v>c7w��f
�Ϲ�J���6;�X�TP���o/��ԙ|���#;�������[{t&15e�.oq�=�G糪�3Qj���'�w��/�}���H�h����u僷�\^�Ž'�IU]�T�z�Bz���I}��e�=�h��8u,N�f��X�ؗf��d�1�.:z�]@'+RƩ,�9f>[�|�F��.��Y��䔊���W��T9MzˣWz�FG�|�R�=���:H�;[I��#w�v�陸�M-j��s�68;���gv�
�g1��S��7@��s��_[��-���#��`��ٯ�L�<�6;�>j2b�O��䈿S�Ɠޱoh^��3����e��R�Ν��ŷ㩵�d�~������mX|J�z�{/�o�f;Ȩc¸}j5�:tLV�o��Y\n�ݕ���*Z��x�V_\�:-�I���2�%��2��A�$orJӈm�ڣ�o�<���e)�A��K_���tU}.N����o��k�8K]�����v���-Ke;������������ğ#�!�,�uf�b��������ة�,��֪6n��5vj�Ƈ�gU���VL�\gG<=j��A���5^��Y�����k�~<���lOg�?E}��@ꀺv�@�j���+Nv��jc�ʦ1OH<3T�ۭ"Ƶx�Cp�P������o��S�V�.s/h�)�����qp���^h�����Q��lTJ��n.4gCK�AN]���ᡸV��+8=�"��t���x�Ky��Y7`\9u��:gDLjt\�N�ﾯ�굓�D���=��\�xzku��^�����Z6X­�f��uF2%��ַ�s7Z9{���i��4�o��a?I����h޾�o����n�圬�,q����X~�V����H�����a���,S�Im�+�"N>瑶�s2�����|Oҹ�JR��q�������ӹwcu��dl&򳐞�]��A�������g�8�k�?�K��4Ni��%�����S���_���%����+�f���5W�H�s�5�Ì�TYs�E���*r�[Ԭ_�8�^nb5���[���� �b�~��M��8I�O%�u��w%�kC�N�u��~'����Z�ީ���zн����ݬOI�)Ec)N��F�J��p9 �Q����,�ꬵ�D3̢�i�윎�P~zR���{I�X���E�Υt��̓;�v�]B���^�`?m����5��
Vة�nhf�[�CvLb�-G{y��`R��a��C�v���`բ��U�IG���=J<�J��x7�� �n>W��ѭ��{;�k7�¯1xVM�NTyN
� ���N8of��;�#u�q�\�DD}�/���aI|D׋�6e��o��߲��9��An�8'=��z����-�{�;q]_kZX��5�9�w�Y���R�g�O�cWH�ʽ��O7}��R�|��瓟O(<ͷ�6���UYΠ�+�1�m92�a�\�(�Ӎ��nn�^��77���\a�,d�=Ү�ήVS�G�v��&�S�Kvq��h�>�	��"���#�[�}�<�c������K����=��OZ���=ny��I�f��$ʺ~��2���p_V�"�y���W�=�t�8���n5���-=fSH��evʂB���K��n\w�/����{谷�����7�/J�暙� ����B�L�μW]�+���f864��wr&�	*.��Ю�ٙ}�M_DNk}~�b��ͭl��঻��[̱�<a9�<"*"Ҟ�m�5�OE; ���j^�s�{���閳�y�g��v�u���(�2�Yٓ��ۇ��nA�h�t�Ok��=a�Wuv��32pw��i��hu��Md�G�98�M���Z��ƚ�U��
�b{u�i��$'�Fߤ����6��3}`6�ad��]�!��>��̾t�	M��קVa��Jkm��0�H��w��fW�%�ux	^4�e��r�:/�ֺu8��[�E���RV��P��d;��$kJ���%�ڽg�o<�"r\����e�X�����#,���}���=P��íP����q/w��:�s�3Q�x�{�\�㘮=�]5�7�x\�Y�T��^n�Iכ��nwe��ms6̬�����X�n��/p&%U]�ݮi��33���Ǵs+fW�F�Z��_��mP\v��l^B���WWu��ۧ���'���{�79���vk����V����������*)	��5l��=y�Z�}G��X�j��T�޽>��U��5�ל���<�J��S[F�c��ɧ ��]Q���/����ֵ���Qm�=2zb�T$�{W�$�����3C�PSy]0�lv=�^+L§�ε�z-D�թ5/��p8z��'�#�[���t���4�bfࣶ�=�wV�;�h���e1�3xԌ6�Q��]�1�
�֜�wg_B��r|��p�N:�YV�W|m���nhAS��v��}�h}y��Ay���b��E����Al�#�ױ�C�U}�,��;|�,����{3˴Ŝ�ONF>�P>���H���v���N�����ڶ9sp�����c�JD��z��A�>��w;d�y�:��v�Cow�8��i/���'�w�m"�0��6;۽���;=!�������M��&���䌳��8J�����N]�\���Ju=`����|�m}l��3��g�<����:,��hz 5����rc���#djg�`���=��_{{_\(
{��sw�~��R�ʾȝ[ک컣���ؽ���NHtҏ�+{~��s<��y���p�o7����^�5:19�T�xO3ׁk���8V�q�;5��[�{(�f9��ֲ�Fvg6���W���}�̒n#�qvX�����9��G4��r><q��e�s���QI���{�uF3b��n��.|p��Z��'��1�=!���[j�̐�F�-���MK�N��q[Rn�N��Z��IJ8[zh>h��Q-軸���a���t��6
R(17)��\�99j��;���\�L�����u��v�;dh��z�����jF98횗k:r�7R�������vu����)k���9�Vv���v������<Uv��0UJ��@�b)�of�9}:\{�3F�_��ugR�O��w�{�\#��̬��7�R�<��BZ�z;��7�C�؞ٝ*����};C�G
ݱ�>:_.^�&W�4��'ãO�m{�my�p�K{L+��yϻO+�e#.��N�͓-�HT��a��]��_��1�^@ꁑ�(J�q�pc+-<vs��7���i'pZ!��D��0�_i���E��EB�U��N;��lI��=��'�Y��צG��S���#s�fpNW�\�V���E�w��Xa��5���[��zw�_Oz1GW�0ro���<[9�'��=��G��OO��x�����"=��u}T^�~�نy;�4�d��h%��ln.x�]�tv{3'�i�`}3��>�9_‧��.fO�0�'��I
p3�xI5���>��uzx�|+�����3��bֶ�ں����]L|�BM4���G���GơOX=�k�wL��o�\�Gjihj�[���C%�:]o��恸�;-��;�r\��z��0)��*㽲^::�Y��w�u�ֽ1��9�:���*q����8!��s�u-�����jdʕ�*r;yք��'(*����z�����m��+���tA���<Յ��i�cV���#�r�#�m�㝭Y	�`#x�	�K}���g�oo�4�fbz�R��	<F�� �I�=<4H'-�T<�2k�.���^�F�*hӢeK5�0:�ި�َK!�G�\X�<���%��}���|ćO�Is`o�mQ�۫�{q�۫F�Wo�R�%ˇI���n�q�|e�@�9��f���Q�K�(E�Ռ�C�Y��e<����Qr�nw�l���6n1�zxl�8Rf�*U��������G�V/�Yos⩻����x;hA�ӝ��x��2�v2�%A=9����ڏ��kC���ID�]�VRZ� Sy]:P���q��x�6Q�a �Ϧ��n�L�w��lޓ��j�����%ՄO��q���
��Wq��w��Ka�)�2��n��=��C��nb��5�m%��_���<W�ֺ2�q6팾�iYH�|z�x]���ĩf\�`��]��@-"�b0���[[E��4��d�����=��m m��}�}��92�.��ɬ�ⰶw���R��h�ǘ��;�dU�����9B�T@�C����K9���+�(heQ�t�4%���݄�P��z���ƞ�ާ^z,ڧ��hw�-^o}3M�0��6��&/�൭�|���,����,9Q����[rRH�+]|��b7�i:��ld�(�.�p6�5u�������<K3/1���c�������tT%=��-�DƆ�`�-@)Ƭɵ�i�+� l��X)؜�aw��m$t���v9W�wއŊz����p�w0tÉ�<�]Š븓l�ķ�0N���'��y�MʏxDP�p��1�}GW�x�և]�3w�K�0����&ox�4c��=ZM�7R� Ӯ��]k�����t5�zN`�df����)�X+�$�}�b�x:7��Ry�R�'� �е�1u�maݮn5:�tOa��wn�Y��`�{A����\ĳ"��噜�ndy�гW�$[<#��aR=��ξOV9Q�i_\�^�H9ޢ�}/�Bb�ͳ�joR!�2���>����,��c��6�JW?x l	�P6��;�r)^�t���Rxכ��.)}�>f3�Nt���[��]���eK�Zc�ʤ��t���]WW�{�⮝]��;4s�n*Mt��N�G]�x+�ohq��'}��S6�M�ҭe��Z�4�[�{�ar\2�B�6���ǶN���}5:��>˘t��O۴%$�9�����"9�����vF�8��H���!;S��E9�d�������$D\�b
*��,E�S(�tsu"�VD'"4*8(�Z�,-Md� ��Q(�l�갠��wd�DAsYBf�-9�r��b*k9$�q3L)9�A��QG,��E)r�4NWV*�2�2;�J8rsȺ��U^Hv�E�T�Tp�*�UDjL�Q+�AF���Dj2.kYFgj�0
�PG]��<��S��"���d��J�����E����k*=@�L�]$iZ��Ͳ+2����$�9E\.G)Aj�]:��Iҫ�H�+��՜�,A�I�T"��jc۷/P��]<��<�s�=���zS���At��
��+��9��ry���/ �LV7 �I�ȧefU�q������Чw	�q�چ�}R@��~�|�Lu�1Ox���-��0����n�f]�I �5锲�\�I��jX�\��:ek�&8鎪t4w�Y��ٓ�������9�nԱҏ_�`���Fg��Q�'�۾}�����bW1�Ƿ5��[gUK��o��𥅷��G��Kv��.�8�-��p1��Y����wk����ml��@�]��}�b��1;��?(y%���C��.:qM>����yHwʚ�z��zvT��^���>�{�����I��5ojJ�m��죋��-�I�ɺ�Z�$�¥�*��&���i�O��<n{�3��##X��R�y�nC�޲1#�]�?m+Fs�ܝ$�%�{�I�u.��[��`Z6�p�ŠEꐌ
��譊֧$U'ʧO�=�wo��z�s)���z:��HF��5
�F]�n�ԭN�i�.�ʖ>m� �MJ��b�vh7{�43GGM��2�b�[B�w7�nP�rr��腫]���
�S��z,�:Z���vk�|0s�;o]&�f^4�^��?�oG�8�w�� ��v���>��p�Z�<�A7��=�
�'��7�ǳ����sg�l�㤦Ǯ���<c�Vvvdt�-�Ɔ�)t��b��)�=&a*f�-+���jN{S�.ݡm��%������W��f/�ly��I��Mn9��N�����+4�������ɛ	�_�t�:,�YyL�{%V�Y������<�y���=�Һ�>�	X:�b���3��s�w��,�Fʹ�jp/r���W��^�FI�}���@��f�y,]��Ԟ}w�֮�K�&R��4�V��9ٝ�j�[W��?W�b�bk4b;�\Wy=p��l��K���},v�w�R�:ܼ��31���W��;S�.����D�&�{��N;��+<�0���ݞ���Ѿ#;��Yl��.���<^,o��kg����mOy�s�c).��X����u�5���]b��n_�#���q��88��h7]��
=�{`ԫg��>Ǚ�ζ0N.�YG�2�yKZ����Ef�yn����/t�=)��"��4e��`�9Vbc#n-��\�m-��v��&�A6m9]�� �e.�Y_�UW�#�8JV㾽�.��N1w8⚛V�R��g�-�d��y非��c9�;7���)θ�� ���)F-N�����m��8��:$�u�ܮd�Gd����#}�C���tz���Ur��G�Z�����[~�i^��l�盝�_��M���d����JkWy+�V��D�꾕-{�y����美wE����q��.��e��M�`{���k�[X�xfj���|��өaR\$�1)6��ǝ�=%�u��|poX�W��s�����Cs�7}ڌ��Y�(��-&����"�r�f�0�0��[6��jt�e�����7����eW�����d�&������	>R���VY���m
qےVm%:z��Bޑq�Of}���s��W\5���5�g�ؔ~2ܮ�4��N�A�\+�{�c��<��n,=�=����� xo�Kd�O1��|��Eu�5z�8���zro)����b넫�ث��ZLT.�\d�1���xָ��U?N��5��m����ۓ��Wrvelo:\�'��G\CK;B`��`]�_���覾z�y�6�91T�<ɤ禾zin��x*1c�%Fm���.z*��=s|r����i�7�.�p���g�Y3_r�6��k��(�jK���$�e�*4�Kl=["�W�,,�:.�3�z������{��O��"eZ{���i���I��5��e��-"�Bt�-}e/U�+S��	G)�n�l�ތgY��w��]�ee��6{�
��r�[=�<ݎ�UJ����b����-gB��#9�Ƒ�X��n�F+�\���c=����/뾦�����9�n:�X� ��_�|��pߟ�{xz��>�=�B�|�����-?cO�-���'i������)��ģXY��W���{���s�+�qڈg�;�}�>M�U�o>/8}ං᳉�rq��8{����+�ӝD�7��6u�*��G7��5���iM��E������
�j �[�"�]�r\x*����GaYޭ�m���N�����������5�3l`���9�m�@�./U�[8�H���ٱ����ǅ]��5;��
�+2��K1�-�j���K�q9K3�-���o6��+֔w�D`8�F����}��ī�cni=)��h�(�S�Q���`WB��l��i�굇`"A��ZN�}/�1�-�+u;����������^Z��<�N��օ�L#���}}T��ك��b�/�+�m����Ǉ��4����o��=)Cp���<����s>�(S��>�؜N�;/l�:���s�_��[Le����Kõ�E�ļ�V�F_�p�fm��rM�˂lT3;_	{��7h�G�J�@v�kxd��ɇm���Vs��~�����r��ޚ�d¨g9�K���;��4Z�y"�oX�]��I*���p�ܿ�g;��#�=��oj�m���yL�1s1)�"����x������[O���]�1������v�����l���{;X.�-ߪz�/6�����߇O3}!�ʞ�j���M��cRl���eȴV��n1A`�[|u��n�_{�3�2�j^&wz�U��F��t6j��-�/yTX��W2�u��BYP�Czй.�OV�u߳h��vF�ݪ�s�b�����|�⪇n_U�YC����ٖ�˒�0^���,�;^q3wh$�c��U}nfwj����9�5.�m�;��	��xl=���9�������g2��5�Y27/ 3�3َ�q�㑍�za&���r�m��K�߉�,�F}��sK)���;`׾��Y�Ur�����1Ɇ�!�����Md8`UM{O;9��
R��[�����S��k�\���R�c@�)f��,ʾG��u��o1�+O�TD�k�It�kF(�����lHf��F�����K�4�)r>��ݕL;��ER�̹�9T����s^Y]�f�4�����c���w[�u�M9W-�`I���p�hr��i�n�Y��m�v��-!p�y�3g�':��=|���GQҝ:^ۘ���{it�T�w�����&�����^`'�dO������T�)@�SR���ݲ�ef'���`�Nُ�P�4EA�z���y�����x1b�:��%��:Vp�wW�2�!���GR�� �k_=1z�z�ơ��M�zb^�)�Q�c�3Qr��"0�Z�v0>��1=]c�ۜ�ɍawQ���'_nro	�yV��[��RWi�]��Ѻטq<��$Ļ9*xVk9}*=�F��Mޭ�sc�����٨e�{cٝc�Uy+\�}jK&� �[x���]Y�.�n��ϵ�u�4�]GG���]K�u/����	���n��b�=	��h�ﯜjæ9Ԯ�q��fٕ�y#����2|\/O[���P��2��H��M:o�r�j�|������3��>���Q�+��Y
X��)�vsU����q����M͖{e3��8_�ru��=�:�![��)�<�F)�1��)F#���\��i��V;,Jr%�Ni���o�D��w�A��3�I�A�VF&c.��zakZ�Ѻ����&هP���:{Y{\6�K������{�d����R�Z�䊮m��u�X�8��]ܳ(�%�kcw���}�%]?k��e���\6&=�7	�<�O�;��F����[O��i{+��[a����L%¹8��	�\L���Jc�b���]�x���ras�V�Ȅ�A�w�ӢnS��Ǹ�m�狴�j�bث�)��{ ������>졐qL� �]}�����6�u�*GV��p'$e�F���_u���ϩ���������w��T��|�t�m�r{�0������ԷI����ƍ�t���ah���x\�'fm��c�8��}U<���̘���ZB���Ox�	�[Ѷ+56���U���c~�"}{Ǭ찇:�����/�<s���[s�$�2�Ҡq��ٺ�[��]����op���ڋ��������=��34��������=:�ax�m�X�ͤ�bw�`�<� ��f��=_\��Y���l�8���V��$�8׌�k�uA�{�Yp?��z��i��mɳ�����u�4�F,�Y��ܰ�Υ\cS��[1+$޹�WZG�cQ;��Fe�:�^&5��s8�9�{�+�g�x�v!��V3# �՛}��rs{�کDΗ�N+�/U�{oOڣ]�8�Ź-�鬴�ގ�<>�aZ�Ua�x;Ԓ�k�Z�m+��g8�O��ΥƟy��]jh�t|�������vp����S2���3�72�}���Y��ZF���n�?5|�d�O�	q�T���ꝸK�Fn����\�]�`��(qdT���R�r���W6���>
h�'�7�Bbe�0Z��UU�lL�${|Yw�CU�>QmW����G�Ʒʦ���~��+��r�z,(�u�y��1���Oq[͸��i��rT%�����}�j8�9����m��$�;L�;f'aM��m��RŹ��4�O�b-�p�L�=��\���.ռ���Wr�7�VG5�we���=�݁��"�n/7�Iﯩ�v��L��z�J���G��U���F�8��Q�મj�p�{g��a�]]�a����WP�׀���1�x�/K����\ݲso�h�3uo����~�mX���G��w����/�*����x6��ŻA���.�-V�0�l�Oa<"3�Jzo�. Bu}/��osk�U�	k��I��-ܖj90��� ����ta_ӉN4��wܮsa����|��q�uoL��yc��X�v���u|nڧ(ի�u��f��е��.�ǝ��b�a+���`D��c���Ӱkwc�D�~�Qw��4ѠU�ߋ��mK�5P�s(����(�@��M�.�=���@���7o_W#�|P�����﹣��'���.�<��[�j|��W^�����U��,\�������f���r�RC]���~��c¨gc�Ҍ޷��?zO@���*|u�Q�4�I3�]�{�3�¶6���z��t���ezOQіi��3��u�9���k��ѓ�k�2���l�W�X���@p{+ܐoy.�Iw3�袝)�ӧ�����5��pv1��q�����|�*k����
�1�ֻsŞ�σ���9\�;�s��ء��0Gj��Uعi��T�Q˶������}&�����;ݮݜ���O%ߦ5���&��y�l���L�]�?m+Fq��[��<�}\�ZƝ^c��uf߰nϰ.���LxV�7�o�ٜ�KcTM���"���5���9�����V��:��.������[j١ٛ��;�2�j��.e��g+�.Or�߁���Ԫ����F��}>�ad�l���"f�l�Vt5:�5�
��
�3vr�p�g����J�S��� ��ygU�3�鶰����z��^�X�:
^���*әg�3&V�>���PK�n�j}��k ��t�Օ�n|����@j���G�z�|���{|=�=(���l�h��I��6Y>��d���rgDZ�i!]�\J"�(��3y�2�b>��{1�d�`M�����>���6���/�K��o)���o0��[(@m�u���Ե�;e[�\62��=�"��}ra��t��2�NOI�|r��g�kP�j�]������\u�\���["��6��ʋ3~Z0S�������:�oxR�;w�7*輝\��}:MD��`��d3��l��|Eb�c4tV떩�įN�g l�T'.����g=�}�YB��dX��MF��r}�םX^ ��kec��n�����@峴tډr�ݠ�uk�R*��8��͙&�2k�0vU蕎��3��ǻo�C:�XsGh��u��R���bݎ��Gm	�^�˚��NJ�ЈwZ���.���P�L��8.�W>-�o���D{qW(嵁;�����E�A�n��G|��a���c�F���p
�|+w�mu��]q΀I>�v%ۻm���ajY��fs!7�-՞8T�ʷWV:� ���h�v��X)yݤ����T\\w*Ļ�0�,�_.����N5���-+Τ�	�����B��齘Ub�����ޛv����]��ŕ���=�$�V�g���#]�^�@�Yt�
K�
�;n*%pƫE�W6���c����C���kR��c�m�!*��dT����oLuh���j_v$rڭ�1;��v��>/}TS���<p�F�Tw���Ν^n�2�K�n��8�
���9F]fX!p�8��gk��ӱ�H�XxP%'�n↉R�@a(s��Au'E-�Y�f�˱G�A�Ә"k1n���e
ʛ�ڰ�c��(��Ybl[����}v͒����0��L5������+132.�h��}y�5EJ��+8՚x���v�{VC~<� K������(���{ᨐ��[�vg,������{W^��b�%H�a����P�;��p��:��6棆.�c�F��.m�w�}��ag�o�^l�v�J����Qe��sس%=�5�9`��e�m�'���Z���ᔫ����SgoR)����ގ�<����A�~�j���H�e-ۋmJY�20v_v�K��*�
�Ɔ������kUEw`c�4WV����.�¶��g�!ϴ �v�c|J�(շ����V��5�g���FD��Z�C��7�o%�bp�Jv�<>�@T>O�jb��\vMXc�Eh�c�A�!�z}����a�+R��њFF'}K^�0���"F�.v�������s�%ҵ��9,���|�1���Avdq(c+^���l,��,���#����1R�𦧌�T�*qf���<�^U
!Z�@����Ȏ��b�aj&uXP�5eP$�DPN�A�2%KJ.��4�:4��H������YT)���*�")1�dҠ��ERg���IiJU(Ҩ�eWL�;*��TU�Ѥ%��\�L�BI*&l�$����0$ʴTr2Т���j�&�J�,�"�I˔��j!8Λ4CԜ�B���c(J��Z\/0*����fDȉJ,�hUf�
��J%p�-�b��s�dr�&��RBs��G
��]i�W+�r����(���n����*�:Tr#$�ujt9�����͐G#�e:�&t"��	Ա�r�TQEۜXA8H�
���Ҫ)���rY(%��EQ�\�U�NAFKi � �J#�!ʍB�H�Yd(ڮw*��y��׏^����C��xYk����@���)����CW.���5O���M=���'�$�3�⵭�j�q%Y��gfoV���n:\���Y�Dm�:�>��ñ�	�*�rTO��Po�r5�ʹC�cK�Nb&S�c92��y��3g��Ϋ��5j���kZq�Ř�ഗ.��Z���ن'�_&��f|}�\�;_�:������u�Sx����\����L��J���vھ�x(�Z�,�y3��犽�y��sAk��kngYz+�X��S�8����㼑1!��m�-��]<{o��O\7��OO�]�y����}���ϕ�⊦1ވ5����ک2Q�R�O��S�y�M��X`5���s
�{~D�`�f�--�7��l�e��ˇj�(�[��jz�R~P��ߧ��.��K���h��3I�Ue�s�g�q�sspN���b5�	�`Ɗ�Ȑ�Q��{=w%�ˀ�q�D�Yc��Q��w؛��v�3<���Ui�����j���u5��_qժ���f����,z������#�Wn��;�.��#v{մ6��O3<k4Fj�ۢ��+��T\y-�9����7��%���0�fHe��n��B�t=�wf�OZ�����}t��(�Q]W�C="��(ME/�;�M��=:]�5�o�-��<���1y�����´kj�1���\���I���P]��@��j�$o�d��,=Ԥ�}؜*M��k4�d[{j�*=P���
��:�T`�^'S�G2E�sn);ʏ_'�Ďibp֟�����p2���4w�hU�u*7�M�u���������kb��]��i�܋����I�{��`����OO\��@�k��F�!����y�1+�8�y�O=y���X��۱\JW�R����&��8;��1�/��`}�r���^M�y�����̟b�3�9�������h�"��by�b��V�u����a݃��+���:SDs�/��Pp�Z������j�c��[�ڙ}���>�z��;>���n17�u�=�xO3�^Oe�w�sop����u+g^�塦I��Z�}�<���L�,�m��8k0T�F��Ň�,t����
�0˙�ܥ[�L���Os��sw�A������L��:n#�WZ�4�W����[�nX3E�����W���)Y1L����/�pϗ+Jw��#�7�)7;�S�FLw<րO�E��t�Y*L�a���%��8��*����{��}uWP��W����ڧmü��Nk�:d�/U����Q��u�nOhA�"��5�������t�����x�t�v�e�_�HŐ^��(�S�Zs_���:����$���ͯs�S�3^ힸ&{,#;q\�RV���T���i�|�xn�\�d&��Or�m�:X���*Kt{o���,GMZ:��n�	j3�wح3���>)���-���j�����r�i8n�V�Yħ?]5�cr���V�6y"�^���?D����v��{�^���	bz�On�Ŷ�V�6�bP������G��:��Q��G1��b�x�4m��N�z�);l��Fk��kR���d���}[������C&��N2�Z1�<Wvd�m�	#|���ż}��+ˊ���P���B�K% �j�͗�]�ege��n�������L����4z�2cw�g�/�q���w�j7536>���ˤ�m��*wn�8&w�Z{Vs1�����^7n�q(Q���=�����N�*m��\��Q>G��u}A�zy�o�(�pų%-ÝȫG_�ʾo�_ε�f���hw��Un��_f�����{5�*�na�ې�y�ev�~��yc�YI�=8���ap�5�rv_��HE�����m�:�^��T���F,zb{V��\姗p���d�Ɍ�2E��{�:Ga�]�kn'ᾛE.��2�+���:#��י6�b"%W,��s��{`�[*���G5�AOm��'�~�5��ת����N�8�j��&��)ғ�
�ˍs�W��z�VR�o-��l�[�'Z�ZCIE[��x�y�n3��,��3�ach�- �R���J{r_^�ٻ�1뙹�!{����϶�V���e���&y��Q=<㫹nO:�X�ο��r1��JM��m���k��CKL|Bշ�f���؆���^�Y�C�$p�*���-��k�t:���鑐��� 9ͪB=��ױz�8b�Z��vu���U�Z���jev�y-�|
��OnS�G�GH:&�	�A��f�qp7ۻ�&=�gt��+c`6/;k��@-�'[��bz��S�;��E�Fq>��+PP^��&�l��W��E�U�d�`m|��S
����oΜ��t�zϮ0͎�w���6|�����G������a� tl�hS|o�tx	|��m�3��J�5��"���fip�/�m�.UX�o�x�T��8�u���{�!�����ˎ�xqGWֻ��}���^�W�-���~!��GҺ��������^ϻ(wK�_g��~��/���Y��#,��4fj�L��o���A�sX`;�E���r%�a��Y|���X�`��7K���V�>mř�oBn�ޞ�zŭ��E.��Ow�%��s�Emߪ��(�6^n���]{�n��JЪq(s:k��{�����c�L��XqF���@�<)�9����篝O&�o:˞�5������{1�9T�
�����rKzV�b�}Y&W��d|ڞl��9������w�egBM�]-ڛ;�n�\��rה�/��/9���j�Q�z#�g^ʰi�w\�4�Q�O�<[F���F:�����J[@��#H�i��7�>��ɩ��A(1�����;���|ۚ��l����Χ��q���y�o�K%��v�Tv���2�ϻ�v3��b|j�(�a�]<�4d���GL�;V_y���Ϊ6t��q�β�3�c�q�nL;����P6������r=V�q�e�E�h�#8�2�b1���ܼ�3ѯ_��I(�+�1b�O�^�GsI�/���J3{h��Y����[L�y6^Ӹ��s��9����i��5��Tݎa��;�>����Y�Q�#���m�1����8��n����xq��-�B�8�=BeOݑ;��o/eM�ʷ�jΏF��n �wU�_/s3�#��]�t�2����m��Ř5i���k����c=mWǧ�=�6]����q�N�y���h�{���i'�)�S4yo���G��u}Tzw��~s��)+{����96�Y�=ռQ�A�Z�Z��F+���4�J�{TR1�a�8c�n+�Tz;�k��U�\"�*�����s���թj��=5�v,���X	�2� �x!�����Xhr�-wv�V��Y�0�Z��w��e]3�VPn���ͮ�5f�Y}�cyOhf���{�\�-��p�9�><w(>�:`�}Of���p�O�Z�O`}�B;d���\%�֞B��+�T�I���p�ܢ7B��v�Ǐ2�*7V�2�qe����9�X:�sp�ϔ�4���]w\5�6k�\�*�����$F�zKn'n�
�O)� ���12��X,޵��4��9�������=ҋ���2�_�>�RB�0�����;�e�mm�}Aw����X�����Mܞ�y��o�.�iMS�@�m�f�Ȱ֗��Z�Κ�"ڠ�ߨ��+�S�k�/5<��^���֔���(��U<���k��������8qv�c�z�^��\��ARS��Ed��{N{+������X[mY��݈&{-ڮc=�	n���˦x{� ~^"l�4-�5^��7���Qo6�Ŧl���G��-��}z�n���m��A���Y�߬���9禒�>�Z�d��zo_��-�jw����u�v|2�Y�[C	lU�jϖ��l6g=���W[�����j:H��[C/9��w�p�|sv�+��{�,�עj˷P�˧)Q�X�v<NrF�5���Y��V���l��5��}��E�;�F�_b�������IJ����`u�*oCc���ٗ�t���d��c��r��P���x�-��p0�reↆ�R���:<{�_[���r�{̗��k��*�15�R�}�����G::݊�:��g�G���Qa����0�A�g"�5��Sޔb�����!w�倃t�O��$M�Z�{.���]�}�r������,f��D�cMq/zz���Yc'�fCr{�����\Wvd6N�,�Le�}l����#�"g�s@k��־�ohtԙJ���r��}����\o#8S��O����WA/^>Z���f?P������q�Y�V^�Y##9;JÚ4䅰+%-OˋqH}�m�9V�r��Wy���|�
{h��Ey�'�b�۝�����pM������3}j���)<�v.�o,R�8W<�8,?5�p+�i}C���Yο����kF�wqipډ�vtk�ѝ���2K�&r(3:��q���u��׵
�����M���9�����{�5pU�2�`��J,�&,Ew#��f�{o�������5'�=��=�0�9Z�'s�a�{�~w�B�(̀��=u�=>U]���b�g�Ͻ���<7Ǯ+a�#AYCF��)�O��{/���V���=L��J���	�������zQ�~>�s׈w���C=��#ڈ�p���H�w�?~����+VJoÝZx|'֫|�fh<�]���x	1�w�:�d��^�I}ّ�ڪ�#~]���\C~̚H�8ݹ�=�s�eV���L'��l�9}k@���E�z*<kyq������~>�(���9�߽��"6��]JTb��_#��8ɇ����w���U�W<���A�/�!�R�����R�}9��d:�.'�{�R羶�H��dT����2��(�<����f'����K��2=�\2=�[6�|}9�É�lp�p5�ߕ�v�V^g<��6��K�Ů�U�u��F9��"}�z	�Q~,Ԙ�t=&�/]��y{���WW�#�t>�����j��zV	a`=����g�sF=w������O;��^��
:�V�x�PV�8Vv����C!Is����[�Uq�6��Z"ui�x�l�֬G)�	3-T�=� =����♮�fn��(+�TX���jIK�+U�W\(�����?[`��av&��@������R�Hأ���뷀Hr�N��_�7�k��E����@EE��h��SݿM9�N�������}Q�sl�����6=֚��T��0S�3/Б�5���H���7�zDl[W���ݟJ�;5���:�{0�<�YVϾ�V|1ӹ�,u{3�}X,M�C���=�(˞1��z���~�S������դ痜G��M���"�'�U���3Hc\L{'+ ���J�)�h4iO�WJ���M�e�|�9�}�~�{��G�����{ۙ����w�x[����'���IU��_�5ߖ��S��)hX6k����d.�3q��=:��.FB�b�}�Yba.�s;�m��=D�|)p ��Kc=�m�p�e^�&3�zjw3��\}2�߼���Z�0��Xȧ����5~�^��R�n���5��G��`��?�Unאկ}e;��L��g�G_��]o����n�]�f+��� �
��N�{�yڝ��پ��e��A��aϮ1�V��$n��N�RG��:�v��R���>e���{������?S�vN{�(-!o�~���U�_� s뫊`�{���ȆN}�^�Y� B�I�ƽ#F��J�ߝK�3�T"{�~�*ۛ3]�4ȫ�ʍ�vS�[��>����d\�Ahn�^-���36�/��#Zm�V́0�+�k�	�6�����1j�B�H6U�}�Yj�ok���ծ��TG=��篝���@�̷B�-��^�6���w������,ʺ�>�Im��]�w-l���x6�}Dz�ov�7�wx�o.<H���M�"���u��9�`%�Rj��!<U'��O&6�3�$�C��k���p�|��vZ�V܃�l�L�G8���>Q)N�%3� �t����#�eҊW���j���[S�#�iO�v.�T���Ⱦ�>	^9쾐�������I�����i���9Ԛ�B=�čN�#J����{{���/�0�1j�	���������j��1����9x���(���V��N�8tԻ�y�7��!�v��fѫ4�.�\=��;Ol�>%���`�ΧY�.JD^I�r���62W��MtW\�ћ� `v���!�]���'n����.�c�դ��LԷW:�T%on��a"�+N�xxк��J�͆��Z�.�Do+�kڔ�DhP3�bNA;�����X �-O���C��Oh�ˍ�F��Ӷ���%�[�	�'u���b]؛��Ų*�vMw�}�}H/�op�*�J���ۊv@	|i���o,d�,�gP|p����7�:��j��jojoQƯ1�@��S��l��_Iz��W,w9�����jcH�\y�����Gp`"M2��ڹ�ƅE0���tr-�@�j7�!�ʶJ�ɥɽ����/Ҫ2�[(��18r��b�Vf=�`A����|���r���܌T�N!Y� Tsz�{A����M/���>�"�\�SM��Ԁ�ыl���em�� Aa�=��92���eC[Y_�N��@Yxq�4�>���@n�i�C�-�3[��ʁ!����W���H�"(=PS�e������y�UG�#|r�K3�N��/-�l�&۫��f�g����Z��Q\x�W[�u�0��

�Y���K͡�]m�y�n�ch ��x��xl�,燴���o2��q�WLu7���������dbT�w8_��ԓ��-�2Δ�]sq<Vs�㳕W��f��v��5繁;A�O�K"7c�G�"����e�od^n;�M>δQ�kG��T���&{��zM�<�Z��x��<����+��z�no��ݼ���T�5\E��n�+:d��;��NV����sI�Oi��!�n�2�I����/)gmidW	�XFJ17'Y>���i����0�Cefi�ch<����3�n���r��m��"�=UFt���Sܖ6jg'T�QA׹q8�,�Q��n>˭��EP.�W���!�ZR��
&o��JFXͫ�34��S�&ES���#��+6�RU��N�")��;��+%9����S)�IĊ�(����S3g"�	Άy92�R�T֜�"#E��`PA	Ċ*�.jr&Y��r����%�s9I�9\��DY�u�*1i�D��QF�\����bXj�®ADNeZ���U�*�LBGG,����쪪tY'���'#ħ'<�U�����N(w%�Nl]�9E�E��q*YT�2����rL���LN�
9«�P�ΰ��UT.J�QEz��+,,��*��UU���rN�(�Q�bl��Bfa�Q+�p�
�.G(�9�#6eE$���HRT��WWw����C$�J<'e�!Ri!/ZW
=a�AJ��i�F!DTTr�Y��E��!�C,�x��p��fEE�����|Dh���\�^e�"*d\��I	�Es�$K�7�_��ޯ�Sq_,
��:j�T%5����|#�=��R�)M��f��dvƼ��;��=NbyX���HsF�`ߌnц��`������3c�C���{��do�x44�X�c�� u5��Ú2z���.ߨfo�_�s��ϭ���>`��ؔa?>ȉU��2=��pϽ��\{w<����3��-�eY{ϔM-��>;��S<�����1�y��y�oԿ:r��5�uWF3�Z�}Q<�͜]��	�B��9�`�ɀ��QP��Ո��/Z��4=�ϥ��[b��b���
�@̮��~��t��ǣWZ��=�O1�4'K�,���U2�/⦢���FD �����^:��^�Y{�7�s�Dz^=)۳��R��?L�?{t�͗��+@�s��]��a!�ߊU����>������w����7�q��D�dz���YS+��Mlx*^������<=���:�vyG���]bYEN{+�ܩ�̘���A��gζ+.��%� ����c[��9��-���Pl3mJ1�{,������Y��>�OO�9������a߳���5�7�/��9��ᑊu79臨�=饀��b������������(�is3m珧|ē�3R��e�	k��4�tҏZ��	q��]��ٮ7ʚ)�7퇎˭�ւL�pL2D[ݏ�ח�k=HԮu�u�h3U����E�i����X]r���1��y;2�7�Z-�vf�XGS)����e��c�t�!�v�}$��qj����$(<�]�pw�e^���S����1ޡ�F�CF�263�p�j�-u3���'>�U�Cuǽ8���-�g�f}��C��s���F��Md���S�r��Îŏ�i��S�au5�绲��^��\��r���z������ a{Q����N�G^�zx	��ӛYW�G���|g|��Y��T�|�Wz��|�x�w��vF!p������!@���"��.�=�Fz���9`X2��f�5���O��6��;�j"v���?z��}~�p�m����G���ժ�x�T)��QP~��~����rp�O9���q���J�ٳv��{p�|Z9�ղ#ݡ�Jw�J��}FQ���U��L��_�*-�@��블S�7� X�^Y��^}��{����+��q�o��Ӑ�lJ2%*�e b�W7��R=fV��{=g��*��H���ɬ��c9MƘ~��u���7ޚS{��:�C�7��Q��J��lC/�#.��r�@��Ȑ��j��~~l���^��ȇ��gۦ���A c������_�bC`J���/����%g��&6ϣBKf�>؈���k�s}E$Vk��NU�e����Z���-'J����ƻ���1:f�a`����cr�i�����X�R���=g\��)4��}Uy9Ƽ�Zs�̲�|�	���FiĩU��n#�t���"�k��k:{F�J���~1��[5P|�z���s�Qc������;�I��<��c�xO� 4�� ��q��Q}YB�W�ݑ*��쁒~o�e�*7�t*K>�>��8+6�{��|b%e�p��M��x���2�D#��2}W�����R�{pF���xO�xH�O��!{�3�������lM�PcS��*��̸f3o�.�g��w5CY$�z�ǀ�G3o�������a���Ly�7#���xv�x\	�o���������mw����n��Ujf������u�
C��\Sj�38A������xv��/�g��K�����k�a����9ץk��B�=x�K���{x�ev�΍�-����ƪ��~#ݓO@���s댫���V��w2���d��׼��޷����R�<o�ϐ�T��r7!��5*�-�������}S?	Uig�,wP���dB�{�}�+�-�Uۺw���܇��lv���Q��NϽ�Q�H��{�����v0&��s�|~^�3��=�l�iCX,_)+bNW7�V$���ގn�=(�px�GcƸj@�}[�G�AcB�������>̼�pU���&r�~9m6 nM�`����/悩Z��܎���\7���˟c�'��'x�s��3�r���+�N�Yk��=ߌz��F�Oc����i�.N+�c������;�1aJ�ܥ$ϗG���싵���Y)��Sc�=q('���_������{�f��<}(e�2ؗ��[�>�&.�3�]�L����n��)K�܍w2��`[~)�o���;A�����KХw�>�g|����8�T/\no�=<A��7~�s��jk�w����VB�8�y�ױ��,��6c|%?Fnd	�*�*f|���TT/_��V��� ���O��1ӹ0��y�V��5��˯��X�������g�_��%�GHQT�#U��}5o�lûݯ�]��V�]��v��2}���LCu~=^��v|��fn=�&ӡ�\U9�F\�mB[���X���W{{/�{�����r�ə��~���p_;�c���.���\3�*8/��o딭~��{��_�^�9Z���>��U9�o�v=��c���~�c����3��q��;�f���b����?EN]e�f3����lރ����m��ό9��eH�^��q���u3V_�u�0ԘK%fZ77Wp��!�͉G�_n��ev�5+��RxR���Iԍ�,)-��꽉96�U�!:Tp�2�����찷/���M{���˥���3֟i��Z̳�L��Y��0�R����=.���}{^�3;���W�`����h���SGXKyw�ܽ����=��~�5��3~��7��eO�`U=�s����]��X�T�>���8��W����x�;&=�7��`1A��d]��y{qp}[�v���7Pz,�g��N�:�sr�����=�s۞gg������M�9���rFы
}�w����~��4"oUoz���k���9�Ɵ��|27�߇�||aM�؋��9րZ��% �À��,�{�}�>o�3��N�o����"wְd{��h_��z��s�w)/o��^�&��/=8���]����{���@eЗ��R}J��B��ߩ�V��.~�����m�/E߲�D\(�mL����`��8������˞��Wݠ��%����,b��w�$��ysվDH���P���b.��Cٮ�_�g����_�ke��c��j���S�}|���ԇ�����bs�T��2j�W��Uo����ڭ�������噝Ȼ�w�.�x����]k��)HK�~� ����H�9�\7Tx~J��:���9�Φ�c��\܋[��i�?0�������"0����T�� ˜"�H[���k{}����I�Ś��GD�<��n�����ι�L���)����0��[)�㒦Խ���l���v����*��]=���\��G+RꙜ�KV.Ջ�}���ٴ�;���p��Ǐ��'�7�n|ǫ*e�P�1�8Y�^/'/�7u��Q�u{�+�U����״T���|*z
fn1������V;ۏeg��P��u��Ux�A���o�������5��2�>�k��W��\�o��b�p�=�������^{����bv�b�4�1A�ѵݗ�"�W�f��_Gis3���o��;�v�ҙ�`�Z���~۹�{�&�O�������2�Yp��u�1�w����q0�ev�	��G�N{�s3�������0�|z�vٽ���4'�b��ඝu^�˩{��z�����mL���~���3�����c�1ڌ�m�P��or�������^g�B�ڕyW>��U��)� �����O��V��ôk�����7�4�xVr�^��Wa�=�	��ӥ#��~���w���v�26�K;l�y�����_���d,H��^>�틻��<P�nq��.!�Y�T�����3W\��8tq�����p8�~��WО��G<��ɴ5& {�6�z ��*�j�TU���>ΎQu}�k����cS�9oZ��8\����{�?`�R��K6�8=�ҫ�Vo�Q�#њ�kB�s����jn����w����+��˞�H��꽳՜>S�rs̏���(�<[w�vy"s��{�֝��Cˇ7ղ�nD*�upL��_�*"۴J�yk֤���$u�Una���{��y?1�RC�#ӻ���ٸ����⻙W%*���H�\���B�v�����w>���g��J�q]��C�)Lg�k���5'�z��D�����9_Lm|�{]m��=��B۹�
��dHr��O�?{�)�y@����l���Rz/u�!^�;>�s�<�V��{����EC���6���,{(�Nt��b=�G����y�6kzE�=�=���;�2�ݹS|>ඍ���"����q������s�5��6ed伍d���t��oww���^��J涊
}�$�sJn |<~�p��^�b3��.4d���v^?{����9��r}jW����x�/i3闓Buz�b��i�T/9�����Nq�̛��/=����Yp�>>��L����6c�/�L�P"�C��/G'�EB����|���'�w�_�n��k/(����̬y������{��c�HУ�>���y�*�ͥ�r���ˑ�C�Š�>������.�=-�?z��e��sU��^eI3�	�j�i����Oa��KWb;�oU�zp��=����T�ۃ1��9�m�*�����\xμ#$\U�%e<l%y���R��U{����07+��s�vq;�4�-��$�����n�;h�V0���oY����Z�ر�*���;�����ߥc^>�c+8)0߯�b�q�z��wDu��a��?nޱMn�7>�>Q�z���n�^�]��7~����N�ψu�9��ܞk+k�W��W���Ɵv��0��Tέ�����?eV��O�f����ذ�����I2�yz���r���b�>��$etPr��\)�����;]�m�\4�ff;��_޻�C���1��[Ѿ
{T?OI���ϡV�c��#fw�[��z���z8f�z��=�jFmw�{Q�_���y���X�hlw�f����P4nr�6z����v8��(�@ڙˮ��c�
_�=w2�F�~)��V��9�E�2;�=g#�-^�5|{zz�SR���>���mR�����a�:���j^*S����x�k\�t���Y����u~��e�d��tũ >�EB�q�V��� �̎�>�9���z���WQ�{/�O��t��jφ:�R�&WC��T�HR6*�~���Ϧ��V�^���.��Ջ��*^v{ۤ�{�O��eU@ht�X7��T]G�#�iX׵����u���1$�]{誈<�
*\�����Gy)5VjR����Yi�5���UqZcu�쾩�ѐ�X��w���yQqaRr��3�U��W���;9�?U�R��{^����p�����.x�ʍ�uc�V�#`
>ާ���S��-��U����\s���!��&=���L����+���5����g�s���4�Oٷ��V�{���tcU?���c�kćJw�tT?2c���
�W�ؖ���(�e��<�џPS�+��ܯ�=�[7�b5���幛k=�����X4`��ڣ+�hq^��5p=���w��A���[pH��=���i���~U�����ڒ]h�K'���ɵL���-}��-p����5/T�l#5�Px=�p�^^�\DV�O��Y'����zo���ޙ��&na�� �:���}�vx���=9��jLfPBe͍��zt������ș�Z��n���!\ǲ4�&[&7�|27���|c�������]�+r�z�Gד&�y1?�^���ɛJ���W �Ƴo�">1z�o������#����Ǥ���[�|4>!�g{�]�f��^�t�F#b|b�S�^b{e_h�������xoƝK�y�<<�#��j�^A���%!P9ڹ%ǱT�m�̯wb�{��k�s'����ϐ�/M�K��ל�C����^�|}�Q:�|�혺w�4 �_qQ1�zk��*�;��(z��K�x��wlE9<x~F}ʶ`c.��OU�IEO�ЅqrZ����ę�����[:�y��b�� �!�#���/b����z=��׫A4�Uvm��|�FV��!2k�/!�G�X1��q���ڱ�^��e���7�f���yW����%r9�>G�R]�Hg��jC���D��7���2b�exYUM��u�l���/�ل�+�Y�,OCw�MG�.�0}MPϼ�܇�>���c�����ƀ��b�b�us֯���i.�t�C�Q�h1=�2��?
��yឪs�2�̣�h�^۞������T����P劭�ϳ�%ٯh���[�c�[��fLa�u�5���R��S��|�+�yo�5ރ,`�Ap�q����z}C��u�*�>N�}>������w�,G����������ٟdK�ޚD	|3kn�e�����"��Ԩ5Ϋ��'oPÍ��Dg-X�a�����e�~�ɩ�l�Oxce�����۟i��VA{��o$�1���O{!qs3���G�Z��kC�ױ	U�`x%u��	���H,�A�Ok���hˮIBGm������z�;q�]����>�Nm]�Rv!�y�6����4���
�tf58��V����m�Qm�]���+���`'bˠ���G�t�p�]}�%�&5�I�岀�2�Եk\�F�����oB�_YWz?F3T�ï"^����:�3I\��	G2�X�A]����I��W���,t�Ăwê�ܾ5�H��H����[�q�އ$(��6nNW�f��S���?^5�q=1F�E����rg9�{]~gF+V�g�t�ѓ"W'��^������9�r{;x��y��-�]<sht�b�|��7��b�hLO/�ǻ���ORi	)�eI���txo�l=��A_r!�k�X������G���Y��h~��s�ڰjאR&���曶oga]g�Ʀ^����n�ehRh.8t��Ǵmqj���+5�qc��$M*�ѽ�"&��wAB��"ęcM�9�s��YҴ��ÚSp>�z��ߺ;���J-�z�l,̶z�ˮ�L��k!�k,f����̝Luh^a�	������.��{��X ���RU��8^��%�ݎ���T�p�2p��'d[�2F(��P�\����)M�+$������om���-�6�YdN�%1hzx]���'j�M����Sw�a6;~dƅ�*Q��K`f�{����m��f-$�5xS�K>I�(V}!�tl���U�XSd��Q�02��&(�S�e΋��{`��[������g��=�I]�1�_����l=m���V�+�`��)�n�-U7j"qp�f�mBOP{�!%�E�߽�a5xYnc?RKߝvpy
��2�ާ�A�jĽ ��)�B��!H�{��4�R��֑�����n�|9�3�(b��n�.YuX�9�w�89�S��b�t.!����slK��M"�?�0�Zf3P�����M��y݆�T�5D<�n�2ëQ�'�ӝ�r9�G��g{9���p�@�P�z�V��s/�AZ���S��nеΦ0��*����b�q+Z�e.���rNܡ0_neG�N����Σ2�V��8ƥ� ����;n�N��)>IS�9������U��Qy�%�wH�܁���7_����4D�i�C��][��iD\��oU��`µg�f6`�	_P�p�� {C��(]��V+KΔu3�aٴ�G�&�*��b>P��/T�/�"_]$l�&��n��_���MZ��yT̂3�Zp���Ŗ�,��~t�k��)��Pq��sC3GEj�'iP��F}ǲ�T���E���Zdm�5�yLl���q���t�j��@� �_��r�>�*�]�5K��������x��烺,9DUedIi|]�DR�S��*�Qy	E��p���AJ	U�D�yp��9Ȉ�4wU*9Rt�-e*���6�E	�o�y4�в�J�"���W�Zx��AȾ(W9���
�0������'H"	̢;;sj�"+��]�W
���O2#�,̊�� �͑\�9��|>gUZT��Q�ա�$�����d���kw^ !<6�j%xl�|Vz�C�r��Ƞ��LkPd�,�����bĪ�V�r.<[�Z����%�xI�IR�*�B�����y��#���)Z�$AAG*>(|6|R��.U&��I�'@��y�L��s�$�T"�����W
�<�TDUp�$������x<z���.��\6��I�wio<l��Lͼ�Gqm:O�ڋ��&7.��b�{C�*	l�:�,�������4��lu�/�=�^�m1uѡD���;W��(���a.����5q{rƇq����m���r��O19�յ���K�S�5Yꌧ\�����O��~�W�;F�u�0G�����G���A^�Uc�X�}�k�əHuz��?]����x99U�՟iXD�uR��y�����,�81���]�W7(���|R!��vyX��9\.��Tb.�͎C�l`L<wp�8�N��5�;<�2���[>	�����^���<0��.�%���I�r[K��Kd�̒0�R�9�gǆw���O����A~�ǶB��{���������Q"[����an9�՘}f='����f�K��|;o�W�=��ġpZF(���!��Lg�kf����I���A�v?=��EX��mg������@��*�e� vC��5S�>J⼼V?	�� �~����z�3K� �ɦ�R�+L�嶀��<����� )��ɟ���N?��sުW�~�	��4�b�f� 3��گG]l�^�S;�� /��P�c/�E�[c���S����yG�iG�*L�s�K�WC�Ɖ^�=�P ̐f��7J���e#oK���?Z�����ze��Kv<ׄ��6-��wM&6%�+`X�h��PMHJ�b��y�n���2n�Ҟ֎���xnYې.�n�����#���̞bɗx~�in��q�zFd��샘/�J��s���C�f|�b�Ϯ'�ĉ��E�S��u�/tB1����Ǐ�6�+�v��w�>���ٿ�ȿO:�����&2�}=�؛�z�~�s�`Q��q���㐦�o.U��~�j��IG���>������k��lJ��ү�귍?`���S�|Wުw��>���:�����W��V��h����m8��Z�}3���;�:.7��)�nzO�z@��Aeq���uW�}�@Z��S�+oӆ2�B1��S��V}�Ҍk���6E����L��}ٹ�ٞ��yf�g�}���v��,�����v�/����eV��w3����:D�u�=�q��<�ݼ��Î�����RC|k%[���yqA̚H �w���'*��op����=�=��Y�e�Go�2f;2�o�^C\A��Q��N��_�R�ұɣἥ'^���Q����7 ՞��38� ��p�;�yC����V��[�&)+��U�y�f���K��|ߘ�M�f�y~v�?`��[w�2��1�̄B~F=�+����Pap�u>+���;��ދ�:��ˉm�6 D2����	�/^p�'t(��{��z�En���逦S���c�Ճ�`FS>9Ԇ�z�Mԭ\�]±��m��.b%�u�7v����yl�]Wi؈t��lbM���ۤ6���WڮM�R��Zcj`�8���(]��7�D��b�uL�?_�͇M ~�s�7#["Y��T��6!Ǻ�A̪�=sp��Veve�JY���a�J���ECwՋ��`t�3#]�Y��.j=1=�����+M�{ֻy�/n�>�փ��P�y�`N�]�T�Hhp��H���F@�A��vm���yu$�����f��Δ�a��y�0&���@��U2�H�U������=���]���c�xr��=��߅��ʯ�Dz���d:���a�Ao��W�������{�b�ڭ��	�~��w�w�/���9S�~L���~��"�`-2��n�A�d�۵�[�ߋ�+d���J�P}�>`ѧ(��{>9[�W����N|~~����Puң�v8�����.�:�)�rk�v��Q`#��p�?����^��[��쭛�cv�� �[���>���[�?���feެ�C�}#�qFx���ш}c_���%��*���'6�A�N�{���
R�뱗���Ӝg%��g��m	�/m�/^�w����>ٽ��ɭ�b���U��ۇ��]h~�;'a��������o��:kT[�����ʇ����)�6׭{�ũ�JxPK�㘪	���d�]���^c�������{m_Q��ku�� ]����8�b��釭�����O[�d����K��C([fj��T&j��k�/˂�S8�+DG~�~�qՈ>�K���?n>밸a>��U��W�
Q<W�V6��O4̯C�0�eV��}��W�u�c��p�x-g�7���z|�������ˍgeb���>���9!Ut�|y�f2��Ϳ�~�>ȝ^/�Ǉ����
��؊�oٽY�=�7|?_깘ǎ���� 7қ�
������-��؟�>�U�6ixε�4���cxU-����Q�7���=�T��g�{�Gc�v.T�#w�a p/���ꆇ���=�Tl����ɽnj}�ϥ��49���-��ǧo���H��UKf.Ո��k�����\N�9�������7��e!R�ԐP�֤<�q�gŚ�z�.O��S-�86�^��bcƸ������}7m�Ȁ�����1F=|W�G�o�,��b��dn���wn����\�'o#n�����Hz*N�V&���7$?с+|1��>������1^��=ϴH�
w��Ύ�����4xT.�F�=��/���S�o��ҩΟ�3&0�w�j:�TTI��*�4~�3�LɁ<*�f^vܦ�F�yo4�Yv`c�	�B�-V[M_j9�}���y:;���hnxY }KWp���u��[���>��i¿Ιݾ�,qWx��$��#�2r�o�q>�=��W���]��2,�-�M����.��F��r��s��_/�׷3���������Q�h��~����u�*�Qs�}y[��'�.���^b�7��:Z�Wj���f}(H�����b�ᦶ�{+pC�o�*�������|�69F�ѿt��s.fm�<}9�a�޹���&j|�k'c�C�����ۇ�;��|��c�Y;ո���+����U�~���<|��j�G���\���~w��r��(z3��V/O�z��-m��T��]8r���������>��F5���z��~1�����mt�vg��LUw2ytk��S�>ܡ/A���n���C1�[���f�Ȏ�\�O��پ/�!����*�!��ć�}��W^��p����"9XB�@$z�G�3Q���ʭ~���-G[&]W�A��{���kwN���o>֭����S�cs�{����H_�<��v�k�C���y�d)�T�<w�o:�����Go���I���;9��������ץ��?+w��up���U����Hּ/bZ>���1��k���6=�������z����4��u�ٷ���ȅ[a��%�}ҟ��J��m߶�bpP�S+�Z'�[Jw�]~����/o��p�%��`�kW�;f�_*<̥U�5%λWc��S�xݻz�oQ��]�|��[ޙ��ҳ���aާ9A3�i2��T_s&ʻE�ĵ��tv�y�um�����+W��u��L9c�=E�0�Ga ^m%����ڹ�_����]Ġ�-#y�cc`z�ǢL���=�9y�j6�����S��t��-�Cbfs�{�YUS�א��C��3U��l��|W����3�t��/Ǳ�g˸��ܔ�a��n��Uߨ 2�C�TT/Y���:7ָv�s��ԿyL��:�˸͜V|wRq�׵J��U���|ș�^���6��ۗ�"�ڽ�c]z{��oӴ�J�فf��yh�8�c���t�y����;�*�u���"o��@��(�>9{���W�{�5Z�t��V{.���C�3���=)�צ׮��s>MV�>��ݱ+� v*���D#�i>f}�E��xI���n�6���~�0��nJ�Pc���bx[����Îdum�;��lX�}U��
N�c��c+oh�m9����h�~�L�@�T�6�{ޥ��Nj9���Ey�#A��iҝ5��U�F#+�zF�sެ]^�u��C�H+0=[g�7��9��7_��X�Rk��Oύg�AS��`��Yv�/*�91�[��g�3�J�>˶4��.���R�[V�*t�낕�b��1][QB�6��E�5c�P�W �|o�b���<;�c1�\����\lڥ|���l�*֠�T�) �xoov�S��V�[Cp<�lv��e�p��ԄfෟC�v�:���&����5�磽m�%��c'z�S�[aQ�4�4�.��_؍�W�V>٭U��X�k�w���x�["7>}���_��>�J?S§g�٥=��)W�X��^{kT����6g�iS&#+�gY0�1ߑ�d�����6ߋ�	�0�[���[/�ר������4�2o�
ɞ�1c��߯�0&�l��ϑ�d��=�<;�}�p�����.�&|j�v�뭝��O��x3&|����sM r�����s*�zi�[b�P�69~~<��Tg}�r�������8 68@����K��w�{2��B!�7\Mg��Z��2��5���=>�A���CB1��l��*g>���QP�pm���h�dޠi�]y�3=�>��'֥�z�9�V|<2������1�܊��
F%�=) =��h��W��g�o��O��ұ�/�p���Ӑ���g���j�3+��M�P`dM�Vo���:C,�6o�o���=;�BWD^нG��O�L��~ ���|�C�&�9]2>�<?K���;qG-� ��ͫLĽۯ#�H�t�F���Ս��F��è�|�&.x�^�l�)�.[l���8w�1B�ށ����nI|nM�{�xȨ�{�W�6{�߻o#�.Jb��k��M��Ζm��$�د+xgׯ~���w�	r���	��E9�Q�(�f��1�����I>��̇�ɒ=NewftLˉ�b�x���y��w,��!�.&,�V0~��<�1�k���+tx��z�o��cLg�|��o���u���Y��z���j�T����4|�~�Mv�A��+n�prsj�kC^�>��ɫ�'�;g7ޙ9��e̟�׾t'=�����X�J��{��ad�����x���*�}&cť��}����w��A����Ȏg�B�~><���W�����˦��z�[�9��U{~՞�Ы���dǎUk�di���Du�c��hq�^��]F1�?{^z{���}+3�}�m�m�S��s��jf���#���4{��LzLF�o�ת��wִd?W��~�bx�-�Y������}�z��Ϛ�Y�3H]uL����}u��fږ�F�d�����x�\�^������7]�aO%*�w��E?\x����)ر�3��]����J�x���=�~]e�[���g�o�"��{�e�yM.�8�~0��+��3�n��T�)�f��A�yp�v�����*��T˙�c�����j�\���JӠ�ߏB_x4ë���w��2���`�r�펍���8�y˄69ӗr��շ��^�=i<�LcV������������TFc�[�DƊ�7�j��D����
�n��{�o�L��ݑ���� j̍o 3�ZCeש �~�RG���I�i��Ͻ^����^��>gon�����L�<��l%o˒c��.��{���^���!��̳�5:՟}��ykģ�@���/���)wX�c�f�~����~;<��x6=C�������o�UUz��'�/ѯMq� ���|�����	}����[���Δ̘���?���E��~�̒������j��{s>2��0;��x���e��:5�ȭ����\{2��*�2��+�e��d�	x��ȏ:-yٟdK�&��K��;j�fy~vꂒ*��P��/c�"������x�r��T;�3���5'�f�O��0�lþ�����w�gW�\�}��K��6�A�u{�R��̖}lG�Z�k���x�Զ��_�\W�E6�k�r�ٛ#6��pџ�:M;>�k��n�UkN�#�,ds�����@�����a�c��A��V��k:��^��!�����b�O�*�3�[ꃶ�1�~�=���G��� �"���Q�.&�`�;�C
��{vۭ��e[߅��-�/9̡�◃'Cc+.�gq�z��{��T+��d�Η7�Db���$y}�����	]���Rv�0#�_�.��[���KL��)i_i��o�\9o�Y��B�$�+qc+��SL�{w��� ��p���b!�G��k����M���S���.���'*���I�/6{(R�e�<�y�s:O��B�������nA����X�nC��#b��(yUNf�!�-ϧ����q��fa=���#���Ls�!�c��������)�R�!V�1�❋�:g�����h�%���8�kS3�v� ���블n?,�k�xh�S��C���z�~���{�l>����]�od��ҍz>gt���֤���5��/��1EߊC>~��c=�[(y��]��ߵ5�k�gѝldL���]�Ws,y�;NW��~|��1����z�%�Bߎ���nv�#3���1:���������P�����QP�\A�D[������rU9��1�ב�U����������ݣ�u��U��ؔa�MLۯ ����#F����Qm^�m~�r~��+�6��
s���?W��=�� l�~���\��/WO��2&�NiH��|<b(�>�2�����������;ڧC��g����b�=�a��,�֓>��=��>��������S����yw+k5���at2�d��� ��`���S�dK�ۏ���`�;s��C7^�[!r79"Z�v�-���F�u���`�v��v a�U�9����o`de��Ʒ��5ֹٴ)(ϟ��׉��L���&�ѓ��!�(�g1�f�u�U�F��q�r���w�)��J_�p���d�G�9Ӑ�����q��h8�t,�p��k�f^�!n�I;H�Y�ÁA���[�N�7Q]ȅ�̩���o�U�v�*�@��ov֎���{�9��~���M�Wy�3S�������3�u9
�d���D��Om��pLgkn�Hj�Emgh���kU�ǅ�=��쒪�=�]�1��%���W�P��~�!���7�w���З�\<w����J���9α�Tx͂�!.�>[p�|"��F�W��<[�7����!�ko��û��1LY,�2��A�T`�:;���X�svtQR��Z�y�ٙ�I'0���+D9�V�xAD�Y��7+Y�������N^W�����u8�~��ԕ�7�ۚ+V���&�����m�G�<5������Z�^���v���r���{ۆ\Jw��n{pz ���j��
�k�l�ݞb�|�}L�5z���j6�=;'+%N���I@����#p�P0 $����|����=r��U�c���g�F]���:��H6�(���vD۹b&���ԞM(g�{�bB�<�j�"ژ�e��� (|�9���U�\����%nd��:	!D:���,�x77d���{��d�p�$�ɯ�G��/���['�����=�
y��+�r�<Ϛ��<U���o*�l�|jtG]��.��Z�o�R�.��	��C���;�c�v�u�w v2ԭ��3����.�LZ��ܜ��F����w$
�%��WWϸ��k�7�^��J�<s�m�/�g
�C!u���Z, �+k^
9�:�T�)c�E�4nqO��Òq�-���g��9�u*b��']n��V]�TA� �p�#"��Y�U��58e]\Q�����h��Y��nt�l�Xe��Fż)���vք�C��������&�q����ڲ�>f�m���'Q���鮦lL�J����h웎���}��os|*r����AĔ:7r���\��O��h4h��Kǽ���]�f;�O�[�^�O2���'�B��CiIg��O�$m�}��Z�5�T����Th=�i����B�s75�{��ܣn�a�ܩh��'O[���ݥ�z��R�E��q�S�+��j�M�(P������hMqޚwBή�qd���ܜ�G�;$)]K�J�cئm/��,]g���fXc�r��lEź�1�
3E���;n��Z��qoW�=�em�D��L�S��.����oy[���Ab��"m;��۔�Z����0[�h��?��ަ���-���!#"⦯�1 ��ɮ�f��i�Z� ����1��O��<�}Ϯ�� �o��eȢ��BbB\4B+2��z��NH�Qy����QPQR��I��Qy�*�B%NEQE(��\����-f-�H��f�NB�\���$����8PDʹuA:^��K�IETA۝"�u(��=.�I����B*�JeEU]2
��J�6Z	r��)�u]۔w9�IG1�+�E�$�.�WwtD��@�ȵTwqp�+kRD9&�켹ĉ.U�:�W"5��"��\��]O$�5̽*��S��=B<�p���ֳ:EVG�s��:�(�N�{u�q)U:Ү�S��*.I	dUD^g1H��W�U��Y���"T
u�,�6VN{9��]�縎���=5]wnd�Uh���8�AP��븲�P�aPU�zy��bd�r����S�쫄����Vǯ�g�M��Mլ%�)�w�����b�m��a影��1>z^��;Ӛ���+��Ezw�/�o�m���׏��@j���
=���o�sӿ?]�2:�X�Oۙ�W��������g�^@O�IA��譧8}Y.��_Q�6��U.eF<�zg>��X@#���~|sY�CTn��������5�h0��VɊ�)���0V�v�7�}Χ�G��=���(�?eq�e/*��{�8t�C���%q���W��X<��[���,�=g����q���D֜J���}�Y��x	1����Y;���Og��ɤ��@����6i�ܚƻ}j�-�鑜��2���ҳ <��؎}�z3ʼ���(��\��yM)�:���r=wǼ|�ǝ�ݝZp�y*Ϣ-��I�u��וǟ�=�z27��k`��zM<E���<�E)�%f�z���2��ep�ºg�T�i��9������
�6{�0�X��UN��������>�vq3�m[$L�.T�#~72�@le9����U��My�jv�w���x)�£�m
����t�Lg����w��/���1QP٥C ^���TLɏiV�)Ahǿ�^d	��̹!�JV扈`����`��Y���wX�t��UUb
�G&�x��:��sY�t�R����U�fe��~�磣O��˰�R�5O��dm�w�]�:J�\�u1�Gr-�K�)؃:1�䙵m���`� ᭎�����;W��~�E��L9�m �Ƕ����d��ҙ������v�f��8��xus�;�3�.�>??[c�=jφz�ԅ�ǦY�۹6�4�_�O�tKPv�bzuZV���:����������J�z��^Ɉ���u;��b�fU�0D����c=dWnRԲT�4}U���\���� �����>#z.3p�s��s>B���� c�0����U8��#r��� S��?Q�(���ͯMv��tc�9�~���ˇG���0�q�����&Ks01������;[������"���[~��2�G�,w�7����_��O��� JO������dϡ{^B���#�S�c}�f�?i �zk��44�m�̯pr��(�yY0��.����v���c���g�����w�t'"=������w���}�Y(�����c�T3���7�{�w�4y^\x�c� �ڹ�|��#�F����v�_K���9��jf�&����fw�BCX����g�c��1?eV���i���G[&;>o��3��W�_�3G�{c����b�Em��`��ec�_a7�D���Q��_�R:�U����P���ӳ���Q�W�:��;g�J���	l>l��f˜
��/+'Zo���Haۊl�{esy���ι\NՓK�=��3�R��z|�
�nS��M:�q���-��ݓ��ɣÕ<��b�*G����I�K��a߬ϲ����2���a`��I~��7�%�y�@�%q������2让��3Qu��R��;�>^��^�/��.��ۯ9�}�����U������=�m�#��;���G��z�cѽ���՗��g�w."_�|T��{����Whއ������*=��	�UR��zD��Xb���~��
�9��b<;m����5��]�*{�~���Ґ�G���>�u;��}+�y8�;���>�Az*�V��Nu� ��ȕp�
~��+>�"���"ǎ����[�u����G�9L��w�Ϣ��� t��@��ʱ5n�F�������0�������b�x}�*�-N�3��Gۢ砪��m����.��
��!t�{=bYEN����}*��x��Of���
��ζ��g6�5���r:�u3�lh0A��7�Ӳ�ezz���=i�~F�k�v;rp�,�t��3��/Y�az�1����ٟdD�� =�Y�#�8qW~��~�ɻ_��f�����a�ˠ�f+�U��C����hvm\W�y7�ю�60N&;(:3B�n�{C�Xro����sf��}��Cӫ��vcʜ��0N\��ŀI��^N�7i�������x)�:�����ǧʭ���=�:��F�`�J�.�����D?{����eH��s3M�Ns�T2�E�	����z�������=���4��e�X�:���2=��ͻ�au{�VB�陿�珀��1ýq:3�n������%��VT缣��s�>�G�JK�1b�.�:�k]�x���~�X�~ �c��C�Se��ʟc8�g�����L�~����y`a��=��?n��h{U��;n���3ݑ>Y���]�O���/Ɨ�������^��c�<��2H	�Y#�ۙ�]���Uk�Mb����f�c�{��(r'����2�u[c�}���}~�4�ӑ���cb���
�ۙ���z%Y�oQ>�Uo=|0F����p����N@�3��複g����O
�8�e��u.��ޘ>�LC��mV:ַ�e謙�E�~ ���5��. �q�d�[c"�ߥ����~�_�sX���l���ޏBݮ��3���-�~���7jAͶ��z�P��1G�~)��)T��d%�*�O�vFϔ���Ƨʩ�jD�}G���w7א̐�h�T����RK�ίA�K4����[jY�v�6�ַK)h��X@��In5._���9_�AO�gqqv��2������Gh���E[h����s����ĩW����3G�e7���13Wt�n+�պ�]�G�x�=˯;��Zǐ��	*#�^cvY�V-�����n�mV�~�C٦�l��A�Phq��^�h
�u�9Դk�3�C�����v���ܣ���q��nB�<c�]~�1������[2���L�:���!u�xo����w��7'
�Wՙw�����cϩOt:s�ݚ%�Y��u>�P�|~�˩i�t�������^��/�W���/k|�}��D3���Əh��g��c�}8�v1�S>�u�ϧ -���NT<�k0{ќt�_��S�h�EW��`Q���ݸ����MG�����ߧ���g��÷�//q׳dw;oچ�����Y@�`p>��+A�����d�Yw�t9�?vә�]��L��Zq�ý�f;1�S��؃�����&֘���
|`��)��m��W��M�1����͏{�s^��gR͹'1��>I �z���׼{Q�/��VMn�A��˷9q�z��]�:�//M�]{q.Mp����{S7(�0$�������_���r��\4�1A��dH�&U^lO����lۓeV��i7��U�#���ᑾ���ߏ�ҌS§g�٥qM��2��ߝ�[S���$����x>7jݱ}x��S�i�	>�N����[qh�L�9�E�f��Ĩ�%�̼O�;�{x��V�j�����[�Z�N����ya嵓J�΋��jn ɫ*�!����I3p\�z�;	{�?��F�b�:f��\��)0��ɇ�&|�Wx���}�T�*%�{N�}���j���Ȭ�S4�V��շ~�r��;20���d�[bx����������u{�m��&5�������*�<�D�b�uL�1~72�@��c�s(O3��W�䵾��5�/c���\�c|'3��G�á�BA����ʺ�x,�L>Ey�RO/__#^Dw�;s��4�w�)�~�A�{�O3�́%��zCC�EB���Ϯ��=��WY��=�ތ���������s֬�d/_!���e��	~��/��9����F8�_��>	����V��~��^���g�"=N�|����N���׻��˫uľ����C���<��x�ؕ^нG�r�|��.9��8<�����e��'���_�s����d8��j
��S��?Er�m��eo�^���N}������®NI�s�N���W~:3���z�*S�޻���{c�?0�g�<ƚ���9���[7�cy����v�9�VvU���g3hp�#�r��&������9ڜ1JG`WY$����k*CZ*!�Ҁ�f�k^*;:5���|ڝ94���^�gt�D�'[��q��m5���ՠgP�7��iJ"�m���ݽ��%yػ&1:�p�ߓX�e/���cGr{���s6���NǱڑީc��fh�zF��H�6���\ ��5E�8��{�3�+���y�.>����yМ���h���៙��5^����xؑ�3/����6���?/�D��8���z?=��o����5����^�$�'Tw�S�q߯�2�~cߝ��H�:���C��-�l��1��0�ٷc��کL�Lk^�hq���跼��!刚2�^��U�W����ǃ�߻Y�׈#Β�8�߀S�a��ǧ]��N�f}�^�w�Ԋ	v��:֞�r� �x�X@�<Wy�Y���!q]S=�nf��z�-���_�\獃��\7=ܧF楇�w̳��D�!�c�>�����xǎB��#��v,mL�1w�W��S�.�T���&����Ƿ#|fU�~=5+�v���SK�d{�N���G�!V�y�n��eTK~��wf�^*^�l�Ue�j�� h{3Y�V��b�)���R�ϴ�ٿ��5>3�!C��}ۛ�z9�ܮC���G�8�U3�
9��@��U��/͘���3շ���T���Y�군*:s=-��7S���Ѭf�en:�͇�H�v#�y���NB��մ{���gͬo����Sn�N�������3O�,��f����8ѹ)���t�I�ݹ3,ͥQM�|E��#��Y:u�Ӛ҆�}l���C-����fdA�oˑ�K��1Q���s!?-ù��2���~���{<���������O�G�*�*�J�U�a��6C��Ӟ>�-A����5��p���zh3�Z�[d������=�`�?:�u(w�3�������h�`}o7����������z܋1����������C>~�3e�&��M,_YƸz?J�o��n�w����Z!��o�7�JE/�K��o<}8�v��w�g����>{7�s�ε�:���cܜb�=�V��+n�g6�B��:�m�f\>������2v'�g��5{�F֮�K���̬� `�U)��'~���z�n������{���V�oa�3���O�VU�8~�f9�\W��ð�vyyX:��V�J���X�����bu�W�imߺs�r�\��{ô21O��=��� �d�7nf��x9�OZ���=��{y�ڼ�W�7��w-D�y���_��>� i�1���>تB�yNs��cȭq4&s��I��s�����y)���V��Vn��� ����VN�{�u��!B��,�m��tۮ;T�2�8Φ�8�<�D��{ s��>���u8��Q�	���֬����|���p۳��و�KR��1�W�Nr8
|�D���U��{�}���c6�γn������Ӄ����E49�����v��U��:s��uY[4UH��v��א��3o=(��L�z�L��Ԁ���k1(\A~�ȗ�lg�i���;6;���آ�2C�*'p^�5����O�6�x8��6[��\�t�le4=��@`�%q�ߊ@�,����]^>�z��u��Gs�}�ǧ#�^�̉����e]��u�3>��h̍V���r�]�ǽ�d߲6�e��VW^��V�c�ǷM�v� �4@���D���6k"�)�ێr[�۩>b��?DO�Ӧ#�����U+�A�S�꬏]l�??nT��.��#��e]�� #֕탪�ϢUzt�ݚ-���Dz�ϕc�����.�M���HV`O��=�*�'���Gۃ�F��^�c=}B�C��?s>���~�^�/��g�]2g�[H������V��b}�CF�=�Q��c7n���-J7?�����/]�~���U��fI��#��^��Qݯ~�� c�A?U9Zm9���vk/��f��TWL�����=��
��u��u�i3��	��y1�,�/��J�Po����	�#Z���}�i�2�;���k�\�drz�XZ���.�T�]iY��"�}Ch��}:^�`���-'�y�Ż[�;53{WK�Uӣ�ͽ\@�]�/���v�Ƿg����F����Z����q��P���z���s�U���M�g�.�8�-g����8��{ӛ]*w�� ���?^��b����G+&�@�G�]�ˮ�u�]н;�ݜ Ʊ�->uI��T�>��2�5߼�^ᨻ���§{�z�ɤ�i4��D���V�<�٠/]���ӱ�Zǲ4�	�V^[�?p��O�p��<iaS��A�>�����r�o���>#�V���R<;��:������k�:�����ǲ{��g��l5Jbd����d���<�F��T�v�}���c��V+�{�R�-����x��!�i�dyq�޶o�����7��VT�c��џ!��ϧ":���-���3�����M r���%�ޫ3"&<j�yG���3�7�i4��lC�i��P�gŘw�^ʁ�����J����z}[5咀���m����}Z@��^�gȩ�S���ϩ^�����p'o��霐�_�X��<*�&���+��)�׀E_u�	6�C���K��/W���fz��ll����1���ll��ll�F�����6��ll����1��cc`�����������o��6��ll�}66m�c`���ll����cm�������6��ll����cm�F�����cm���e5�e�xp��!�?���}����ɀ���@I@)�A ($ $��PT���$;��D"T�
P��j)T���R(IR�J�J�P�R�   �5U"�I)H��� ��*�(*@EUH���UD��(*Q)mTD�7�E Ϟ�C`�TfD��3 ����fؠ63ZaT�� 8 3��J���QU��xs�   w;� P�`  �� j���`�� �F�h�< ��%DL��Zh�6j35H�c
��Г1��� � �PWa�Q62��Sm� ����
5�*��ZХ�ӉT�A
H
RE� �5�5{r
��D5Sj)��u�յ5;����CZ���T-�@1el-�c*A`2�	*�Rx ��f\mk٫$�4��5T֚Ѷ�7v��Q�5QR��6�F��v+MY�-+0�% (N� /z��$� �A�f�QU[i5l͙�����b��ZV�ml�X�Mj�XWJ��P�'x ��a��*e�Lm�6k+ ��J�F�Z�U����n�l��ڭ�m��D@ �� wx
ږ�6�6e���2�Z�e-��Qh��2Q#UPT�U� ��
�l��+a�K1�Z�%(A)k*T���Д���}%  ( ���JRPC&���CMC@�{C
R��Bh#A�M44i�ɄQ 4FM2�dȓ�6��Q�
m����TU  z�     ����)�z&M2d� �`b`�I� )Jbaf�4ha �<�:��Y��o�kՍ���t���1lcb�l����QAP>0�9�� ����Pl *"5P(�̀����>������*���A�
��b�TPT0� �B1VPT�p�}Ӧ֪}:��-� �����&��uC^Q0�9I��d��:��~ɰ�/��ᗕ.�!nX�Ğ^+��wb4����g4��B�F��v�D����à-T����7���3n�kF)�+5/^Q�Zˠ�M��{G.�3�/(��n����3X�R�$袊ljI
�6(��w���edWw���U� �n��l�H�
v�r�ۼ ��D=u��ܢ" L�˂�M��CC�P �դB��+�6�n`��Y�:���-w-n�)J��җ�e=
�7(Sڕ��{ݬ?d���Z���ޖ���9%����L�C��X���4+.�fRUf�5����<m�,ɢ�&7�Mf2&%�KQ��U����[aT�X�X�X�n�n��0��c���]j�J5+J��Yj��Bٸ���V`l���R�=ib�(�M��t	��h��Ϋ4��O���#m�V�E�;���/Cw�	A]�ٵ��ʙh�+F�Zѣlr{�mbޫA�E�%Vp/8�jM�h��n�����4����KYMj�7���r�S˹Y�2�WH��v	�k&R�4[ݽB����nܡ�,V����DY��LK9q˷-�x�������{�&m�����Z��C"�Z��WY���K.���ׂ]��D��l�X��r�]�P{e����heXwL/��|찕�=�5���H-��R��]��{zh��ұ����U��i�Z7N��$p���rJ��k���aaD�:"8t^����^6����5i�h�z�/� �)�u^�fS̚!8E��sf!YWJ����6]˒��0e�4}�OukwAM������6|Q��xݜV��$%V�^V�%m �����94����n��{���:��w���u4��& ҹ1颷/h�!��{x�[�7m`0��xt���υ��T�#˦v����U��6%*�ȉ
�1bn�Q���24A�����WI.\_qu����{�k��Z���|���2�ͽ��D���T�T6�wB:���|��^��q��k��uL�[vk�p	>X��/�Ata�G�)a���N�~�Ǌ�4n��u��c�|�S�����l����{��N�vh�T�\:��owd7���;�Ps$xRˢ�+����9�q욫d�ϮWNx�,�W647W�WIV]j�e�荺�D:AU�֬:��ȴL�Q��J�i
K�]l�Y���:A��U�d�H]��BP	dn��+j�:��°7�+��=6�
��(Έқ�xN�G7ϨfY�Y��:�u�{��6��7*�6��n��P%z���z%BaDݻߍ�
Z 4�"Uʰ7M�T`�.+T���f����*�ق2򛧥nnQ��m�Ԧ%�$�kD��!B�4�Û���དྷk���px�tx{���(g�����j�ܬ�㺕)�{�z�]e�
)V��U��д�[1�q+s�������Nm��Q�$c5ύ�9ZA�M]sf-�}.Q�[�U�83s�L�����fV����e"��[��!"� �'Fˠ32���aʺ-^a�Lc����x�V�jj��M�t���N�d�����a��,6-���R���Fȭ�e���ͼ�Hx��m�\�R{i�u̪z�;��x�Y�d_o�h<�
���e�7�g}�Ɂ�1��XaS-�ئJ����	��S��ʙ�-�*]YӮ�3��ph�6U���$u������9X�YD`�o*
���"��`n���0ę�.�{NK�NS�7C4eKI!/vL�xc�[�[��Bĥ��z��d�Jf�N�#X/mG�{�V�zU.)�I����5���H�*��R��!���ۛ���.��*{�a��x���T���p{���]��d40�0�	=zM��YR�8�H��{����/��T� 
��ڸ�_Ѷ0��թ�*0TQ�^V�sh��ӶAXA{O5�ڷpaN�Ы5��P4z�wX��U���U�s�v}zNP��F�'-�i[��q��콫)��)GZ��
 �V�Ժ�K1GWQ��m��*�3lm�M:��6�[ba�jV	�^
ͣ)����ë�b��9��v���:ݑ�n��c0г�QY�򵕆��r4Fq�;�9���4 �gJ���@��v&�Sr'��m����.lXiXK]��jB��Gv�{�%�|�	x��2p���ɳK[��n��A���ԧrѬ���
����Ww���(����0#JR�<�ǃuY��k9�Gs���»�-�V��*�Yl��o̰�1�Vl:�!���p�� f��CTא�D��.��t�i
8J�B<1�Ȑ�6 ^e�U�,d7��bXpiٺ�K�/�� ��g��K�E1�A{��t��.[���,����Wu�h����5��8E�v�S;�m^������d����T�CFTsHt�'�#Ղ2�O�j1Ɏ4�!a���i�Y�ue�����Bn�aIHGB��u>�����̩I����r���+3��b��Z�����
]f���*�ks�M����"ԪMخݎ�3�R�4Ӗwl���"Ǵ6ștŬ�[�A
`	�6H��97��X����i�#:hm4��F̬$��N�ܨw*Sdi�2c͡�Bީ�CsM��emZ)�(�8˗,��06���4�I�&��U����Z �QЭ��vP9�fiAӧ�uѡ#�v�5�n��twCQ��0����h�f��x�Ȅ6��r]�W���n�,,te�m�i��x��q��m'�b��؏4��A��!�e�*�ͺ�7X�Y(A�M6��ݼ�ե�t����W�zh�h�(��y2�ټ�1�lR��Ȕ��W1��Sg��	���-Ty/�Q&L TE> �KuV�\l�an� h;w�ʜ�vp5"�Ռ�s�Ar��A�L���}��4�{͖���+cF�mU��e�d���/%��l�/o���kC9t_m<~��YW��p�Ҟ+B8q}�P�w�^�w���u����Y{�iQ��⫁�-�J�A���^dw�ɷp�s[{�w��i�9��x�ۧ���)X
,�#h�J�st8�Ī
�m���u���á�
��/&�v�Z�W�jbı�6��-�0���ӅtM:���K\�^�.EW{�.��-Z�)[:v��oh�"+���Y).�N���we���vh��Ӆ3,ި��/-�if)���V�Y�:4��,�l��E�o]d��7J���-|�Z_\]����&�֪[�l�=��*W�3t3*j�ܭ���F�{��NG/[�؍B�a
Ewk�cժ����W��ƽNYs0���sK�q�̬�H�@[A��-}|oZE��Ѳ��]��'{�H�E��9��@��2i��hYg&��/,�@1�r31�9h�d�hly���-�jh9G�p�]սu,fn3�/�;��4�G@Q�2��֭C���
ԁd���)�E�.h²Cj�M�2�iY��8U�x����"�m��|H��=�շ�b�)�y�#<d`=�^�ʶv���P�^���`�olm,T4���'������PՠS���3'�A���گ>�S���iFX��-j�j�K�۱3tݼ���S��5���T��S�CIX���B�eR�9�R�ݸ-@w4�ܽ��&k7�����$�m�D���y{��U�D�Se�0��+4��*���b��m��eډ����/!iYhK[�t�'B�ڊ_��Wi���e�D@�-cԎ�tC\�Z̦ku�p�te=���;��KoIn�� "*���P�F�!�ڷB���w���兼�^��K�(!�(�7�2�5�����v
����]ܶGח�I"��u*��_M�3�ɧ�2������XAm4N�1(�i�=u�O�X�tJ�׬�,�ź��^�|Y��7��|m�W�s�����dP{� ViyzU��;��dKV�Q�vK�z�yf����ݧ�m��,�5�lm@ǡR�jе}��R����lK�kE�z��u=�2o��
<@ a����}�q�?j?c㱤ȑ(�.|��>�X��>|��u����+&�T`-�[( ^�]��1uh!�eKr��� �6��z:lEm����8՛�v�E���q)PHˬyx)a㳱9[-=�Ֆj)�*۽t�e˦)�fPy����R�f�؂ɳ{{d�3 �a:�|���fV+XB��1��J5��]i�jK�a<����or���yY��v�K��5�4�\�@�^�%���ͱA�+*��]�D!3<߃�Hݐ�ŨJ�f�U�CxY��mj�#|P\a��'B�e�5���y��Ϡ�]K��2|p̮Y!���D=ݫ�	��k7۩�k��R�	�i��)89j�gƝ$��ۋ���討�҅ҽra|-��N;����ô)3q�ٰ�}6�7}��_J&V���E�xF8������[B=�����������,Z�����aʥ+��)X�iV��W5����V!���_��ܾaߍء-nX��tښ�
��:��n��t�����r��	���f�Cݻ���[�Y1�ٶ5�gl�(X3[Cs����������ܕ�Q�S��։A¾���5���W���θ^��� 4̓����
B�M%���
�͝u1�Р��{G�6�TV2q��،u9�G�{���{ǅ�/d�;���ƴCӱj�OMâi�<u!Q�-��M��9)@�$�phO�j)��9�Pv^�0�@�qg,�Γ�z
�Y�rc�"9�ٹ�o"�N&��Ng��N�Ҳ�a�-w]���J��p>��F��i��1B�LA��gvŇV�
���NN�V��8��9��\]:�����oLֆ�-�$�6Õw��w_-��*i ��heH�b��έ����_ۆ�5b9�ͅY11����6�s��/<3�
w�h��8ֱLJ��䜜Y]��X���F�[����JJ�u��䄁��
�۹wa��^葨���|�̱p���pP}G�#~[�T��>e�����������m�WWDǒ�H����V�Sëq�YOXYX��zG�ܲ��i�V�Z�6�'���ȱ+��(ꓶ���0!N��вш�펿W,�Պt�Q9R�ۧ�h���O�B�I�fQŎ�`cfb�ة���L���nZ�������@b�(�Uw���G-T.�FP��L�2)���G��xs0�	�Y�������T���r�BN��W.!����X�"3�ZJ���Z���W4���xv8���S۞u���U�U��	~(�z�� yLՠ^�C|�R� z��ݛ���z�����s/�.Y��6��mr�Әz�'�gU��a��6*0,��Q�dP�f0���h��+���g�w��4nn�n�+VKb�lb����u��ö���X��SBmr�ݽ�
�
�=�+Y6'+K�2�]f�U�]N�MV���5�]�V�����od���`]"\�����oz��IU�{]ݚ$�Ҷ�U��ҴL��|̢�P/5w���ld`���cW3�=t���"g;w��UB�i��q��"�^ɳ�ɩ@ޅbf��63u�̫�{$��S�k�#QB�E�ܩ��4�Qަ)9v�ҴbZ�ΰN�6�Uu�Wc�� �ի�X�K,��rW^<�X�$�Z�s���Ү�:JV�<�pG��t�od��#k)��T�`ïonv^��m��A:��l��s# 36Ø5�%K]թ6�S'�N�,@!5�;K2���:�=HX�i����k8jSo:�3/�wN{����b�����&қL�����S)^TD�v�:\�AM�fG�H5�<Gs[�Zˊ�q�6
KQ�!t�|�
�,)�l��7�_>�qK9���C�ҹ�g��&���-�7SPln.��C]h�J[]����gX���d�lCk� ��iQ�/�l�.��2�6�d��K�D�r*6�,��(TǓMMOX][Ɍ���,�h,=����\ǧPÂ�mԦ5�PG�Wc1W5������m)���>?7R����$7�����1�&.b���Xkd�>F�μ4�� ���,��hĴ�p�y:n-V�mM5j��z�7z_-T�A˚ԍ���o ��u
ݥj�~)�5�T�ԧ��Dv�F�>�a�����Q�]�5,H�Zj�%v�sm�@����>}�V�lY�GE%:�/$ܔ��ş�+�M�'m��-Y��|u*k�t�L4���!̞ڎ����P��q�Uܡ۾�����As^.��g�h���v����4�m�������6�3���I­�<���������T���8�M�&�9p^ܒ_��Վױ;
 ��й�z}�2{��B4��9uqģE���aV@%�C�\ӵ�0e��-�)�,����ص
K����c��wl�*Wc�捜C�����e��)u1��ƍ��w$bV�������;�&�붆s��lѮ�9��
��6�һ��ᙖ�|��
���܈b暽iH���f�s������K��4��6��c��D�û�YP�D!\�g+�l�K0��[a��{ʑ�EbyӠV�ř9r����)�:̉<.+�im�|.��3�ؚ��.���� `:�6��v4 I�oCyT8L��&���5ΐ�Xbu>Ev���	��WA�J�,�.D+�]���	7*Q�Η1=tƐ�8j:�p4lؙs缅ff|b3����ga�����qI{Mn,�꼁����q�s�G�mt3r��N��+���j��f��q|t���>K��YV]�]A;���a�+���('�u�@�f�c:�X��R�	
A��W�ͪ��׵�{r�ڂ�2E��7����b��5�(3}���_A�t2�)��h0E��h�,;�+�e�{)�aK��U�
��Xȍ����v�y�,;����;Mq�[D��s�/e�����7gA�3t�J��]�Q�F���듳�91�5��:J9��1w2t����,ut�js����T����Wd�q��W:�M���J��� �4���>ܸ�8ۡvP���r���f�"��x�g^�T`�y[��:��;X�-Npp��\''VjEJO�
b�š���U��BV�|^�O����8V�%,����	���'�YV/����6�u�h��v)<��!M�B�U��=P�s�5
��s�.U�3$ci�'Z�0�A�@�S�ܗBp��*0n�
�Y��m�q,p�uQg���ˏA�c�����k� 0�|o:fFxF5(�ї�M�Gz��W�NTk/��H��qJ�pr��F��V ���K���h�Ӷ�;gAu��r�*�oq�雘*�鼊8 F|/��j�ண��ۖ
����ӛtn����2:[�����X�Cx�ήD�X6�H��zsC b.�(�]��V��q�n�C� 뾫����:�Z��Ϧ��ldFU�W݁%n�o�lԩs$���U��BI�R�����mX�	�]�%���*�gs���m�zȾ�Z�T��n�ݣ"A���֧B^an-�Sn�
�slv�Q�Λz��DŻ'iS:̾k��l˸-r��TR�"�Β�V8�@�%���|�F����nnP��|s �sd�]�o#I����q�Ƕd���V�mȄ��v����mT���F��\�F�)$�I$�I$�I$�(�LFJ�rP\2I-�㐸�-�*4>����2n=�]c2�o�U�5ͻ�Hԏ2�N]��)6C"R�6��`n����3{x�j<Q�˝��e����K�yE9�IDS��;2H%鄙$�I"JI$��$�3f0��v�uwM98�k����9�oe垠s#�ð���FS�R�$�.���.̩ұ6�:\�tAeu��6��%�U�	��Q��ֳ�l�T�ݨ����72��j�e�i�{g�y���*�f��9su�D�e��Q�:h�y#��ޚ2.C��6�֮ma�%��#���f)¤��\�#ah�:&)
:���8��Y��o,<�w6�o��ˉY�:�Pr���)gF��X�Y�:���ʒ�nL���^�9DeLr�-�;�TN�z���T@���E���ETwʈ�Ԙ�h
�u�MQ�ޣ;iΕ�3���̢����Q�G��V�Z}�q���-P��n�9��J��C�*�ؾ�N�����ts�h%܊k�I��ׯ���r�U�d�h����b��{��Dh�Wgj��e�ES�n��i�#hu�l6�1|>ɕ|����~ys�o�*�w�\!�ա��p�sC����6�����8�K�KB�tرJ�c��[�C�tQC�"K�����uF	ڮ��ӻNY�on��{xL�^7O/�w�j�_��l�ځr���j�'N����-�F^���Xw ��!-%}S�}Wn]=v��R>&�m�ر�E:�1f�����"���yn�*���$f��-��(��5��^�@�Q��$8=�񙙦^�����U*>��KI�����;��qІ+iq]ԭ;��_PQؓ�Z3��h]c�����҂*��-�ϲc�����Ė폳'V,a�`1%:���!\��ھ{gX���NF�L'̬2>�tQ�N'Yő��^����ب���+�Ww���SR��G9̭��Zp��s�<vQ�2h�aVPc�r�r�;,���sK:hF�}j����զr6 ��n��H��!Zq>�%
��5_1�u��R�rLdWP�F��4�E�Ҡ�ruvZ׀�*�1��:��*�>���5����7��;����B�
 �e��k
��),��%�������y>��9�xZ7�j��
����׵.P����(_D���jY�Z7Z���d}����D�^eKE]՝v.m@��}i��� ol��} X���wk2P6���@*>�zoW:jX,upP���N/b4c�V��\�3�ڱn�!0�k6J6���{�kmT��k�lkЭ8SS+�Re.=#̷֣���8��o���Q����2�XZ�op�i�K�V�� �8��W%�6�ң�5f�n��R��x�y�t��Ц�ޞ�/�Ifj�=t+l�**�g%IT�7�լ�aw]E[�+tj\���C�vʃk]�`Wfh�K��V6�m%��g^�
]�9� �3r��otuu0�m��Aܳ�R+ݮ �Z�WU��x��K�ˮ�+���sN�qo�� �a���0�+/�m(Ri��F�}���w�M�k��[�3����2K�s�ؚ��[��>b�܉��Y�P&4V�{6L��۷ܰ}�oB��]�wõ�An�2�Vh�ۑʗ�ۛ�V��O��jV��b�:��Zh��(�S
��d"N�^Din�}x�i��ua�E��T^��{X���w_�w]�oJOF�71�mYzK��A7\{��k���QCN�6�I�AW׈�M.�T+&�4#F�y׽n��6U��=\��Cj`5���)g��x�"�.��7c�mv5��&�׆�JLW^�E�BQfp,V��m�'Z-_*�>{���XSI���R=�c��p�N�V�sZ0�f�t�A��Ħ#`�M��Vc�������!�V7�������G�Le�a��RН��I�+p<�Mi���׭�i���T�*�-��38�gb� �� ����Ʋ���3�oLT���K�⬁� �}�J5A�gU���c$���� kK;%)������y[�dXk��4��&�����a�:@3�X���K�a�8+���ֈ��y|U��Πx'{��{�`�f�4g
�v��j���P|�,�.sfb!m�*V7׌w)�����J��s��w�p`���IǷ9e�h	��v�5���P���؋�f����ئ�����,�U�֞�-�a���^Ȗ�or��ɕ	�z�u��ʒ�1����5�_�5k)3�`қ2�T;K��TO���g�i;���y��Nt1��x㖃b�Hf�m�J�Λ#��SW�z�*۹+m�^��v�H��[�Uy�q�:#��i�x!��~Q,����uK��.��)mg�An7g�IiWvs��jC��`kI�������5Id�c���w��]��"��f���g+
�ֵ3ǹ��L���H�c��wQ�v��	�ͭ[R�J�z�v�%t�[{v[���ʑ]���y��B:�t]*���)_87o0��rY�ƍ^��*͡�h��M�6'ee
I�|&�.a]�Iv�;�R�W��<;�敶��#�<86��+ ����@-��k�Mr@3�5�|�T+��%�_�&b�b|��B�e���j��Gl�V擖z��u�z5�gAbݤz����2o(�d����[j���R�����r�����C*u۸l���C�����q��\�ܱ�AJ�>�6��jLզ1�k Y[�]�]
-7�y�4�)�ƌ�|6�J�U���ݍ��-Ң�ּ	�H�4wnDsFk��l!�U�s+&���(Щ8断����y#n�+�t�3��1�+$Ԫ��� sJ�h��
�,�m=[9;�C탆���B(��e	V���M\��ȦA	�o��Rv�.���P��(3��9�,��.Z;Fgv�-"w���:��2!*
9A�yj��j�u�$�Td��Ǭd���[��2�0����8�9U�`� ��j¤�:��-�d��8�4]�Y��Mո�Wl�ݷ9<�3)h�v����IKnJ�'�Y$��%�0єoT��w6)rg_p�ɷ���� *oVZ���p�j��&�_)��'H��l�����u˳;8�}��9���yo���8z�}�C�Ǎ� ����`��Jڭ�dT&��p��S��q���$�^����N�%<�;��6�$�k����}B�)i�V��z��'y�tŚ�l���^>��ռd��Q�ִ�0ٝ�i�/7�D�\�v�#��:Azj(R[�NV=�#&=?�������G���a(.8��Py���#��1���MX�����:�����],�}-<��nͺ�q	�Y��w1/2���]��&�p����t鹶�k����onS�wV��U��I�-��>*VR���p� ,�(��°ԧSu�3bB+�҅��eAƕL�;2]ݝ������6�(���Q9���!�…����/Y:�#H�倎�+�)�H3�A���`�9�������(d��gt���!�}�u���z���h�}�(��Ю�V�FX"Ӿ��T�H�Qޭm;؄�dk�c[�m�
��0��pj����n����{�qk�gO_Y}��W�,�{Ǯ�t8)=�%�w]�}cO
�>ܷ� f�O�3�JH!���]��;��z�u��t�t�nS�Oc5�%.�:��u(�gZtik�C���C[!���P�[����7#r��.f2{��=��Ň4�N�o^�麐�#���6of�Td���@���'O>�^3K��&�����D<�j��[�
���m�6�w.#�N:�T�3��O�X� ��Ws�tvݾ��0���+g,�j������:�yq��R��C�G�iE�\I& �b���iV�]�];4���.�dj���#]���r��]WX!,,��ti5��h^Lu.u+�]O.ѫ�Y|i�YRl�|���S�s��ۮ@�-G6KďPQ��1�+�V�q���Ҕa�)���{n��㶉�k;���rG��j�ێf��49[��[Y�y��ѭ�!�hJ�p@¬�pdt\�z�;o�,	3��%�n��6�C���+w�n`�\��+��+J�I ��T˥{�.kLucfț9��]"�ʗ�֓d�����f��K�8[�ާ(��XO>�'t%�6�`�C�`��9�p�'1�3��iq˩���̖k��)��IF8�݀�4ve3��+M��qF�Fm��me2^���[���"��@{gr��`�G5&	�9T:��'r4[�3�Ve��V.��`�ô|ԛ3Jy�����btd+'>���k˺��ͭ9y�&f,�T���RbT����}	�dPn�;t�9��/�
�u��nV�Ew|j�Pv�T~j)�}Zm��Z�yX�l55�
<U]��y�gz���>�	 "���hG�C�݄d�_���s9Ì�rkZ��e�]��Wau&7e�%v����(��p�[g�b��Ԛ�^1Lc3-�W��hn>jp�t�S$�4�x���T�_��d����8�j}���L�Z�����m�f�s]e�-��a^A�%�y���lӾ�9��]�Ir!�"��JԉSd��(�	����}���qvK�m#Ρi��N8���;m�mln��ƻ�Fr�J�
Tl=1'��ۖ��h������#��藻�j�u6Y��Y�K��c#[�GU�Ռ FmŰ=��2��F�Kf����5R]��:��t��ql���Y�usj�Y�<�� ��<3&�d�޷ٜɜ���"��w{`�;Q)zk��bU�y� HǱ�
��-��)Ρ�gY:,Anb��|a��[�:����txn�?��=d@q�:Y�jT��6T<�B���P]D�o��S�뮹/n�8櫗����²׉ʔ��6��/>�GSN��e�fE5*���Z^��8C{��a�Uԫmle�2�w��y��s�>�TQi��4��|�R�qV���S�d�CXi�Ra�i%D0��PV�*��藏_V�s���*p����z�{�IJ	�Ē���(��k=)�咭�ܗU���jVp��]�(��bjU2g���k&�}I�+F\��y.Q�+�UT�<��>U=�����r
O�_{[rr|���2��c���5+���B	�*��Oz��`Rz"�}t��������9�I*����ֱ����3Κ�G'��EPSD�������N��ڿ���/��a ������y9�49�U��-O{J��Y�8��AWir�����x���ɸ�r��L�����bD�ʼfc	ͦNQ�'t�g
+T�������.e�z��zi�G4� �����-� �L�J%�h*��Z�b!��m�L��.��΋ܭ�#.���PV׽+y!�4�A$����5�;�j�m-;��A����R��!�������B�Hq�ؐ�rg�l'ݍ�(U�0�Tq�b�gg\S1��e��Oyf���H��{���1u��c���)���HF�0���Wݦv��=�q�����v���â�6��"���6�"Y��z;{kg�M'�­�w�Q��&6�wc׎uk]z�����q�ٰ���(�����y��Jr7ݹ������x7w��P��j�C�i�{��+�K	Fա�g9V�##�R�1z�H���m�:z�����q=���|ǈ3}��d��ˤ-����鸮ʹ��R3Jo:��;�(a�Z]���n�c�������C����I��d�&�$��o^&�W7��O�%����@�{n��'���Ly�ytg��p�E��QV����'9�"d����L���ouN��vGn��鞸��q�d�5�Y����_`J��Q$Ӭ����u�`�2�<���g�����\�Z�3,k����[Sd�;i�Eѳw��;PXr��e^�˚hR�ڀ�:��qø��fN����R5�5B�wNmE��)ئ��=S����u����J;Va��&�^j�� �I��U�c�񎜢5C�sr+�m]��P�.#��miM�q���|�Z��;[�!����7qOf*��ĺ��is&�B�vn �E���+ �Q�h`P��y�P��n^���flt�.�ۗ1�W�2^��3�(�}��fB�X~�7^�R��o�o�N=���#�=�Ay��Ů��\4WP.�ʸ����vD�o����J�*cu�5�d����*U�n*���1��r�D�ʍg7���ݽ#k��#Æ)��w�&��4+YJg;�ϳ7u�%�$}��L��K�y$ ��|�q>
��9��ֲD��ی4�.(�p*�z7{:�̘�Ey��!�X����{��U�$��I���$s�4^ȧIrYD����f�[�W^~�������P��ju/:]h�nU4��DM��(3�=�Yý��� MR.��x�2�Z�����&m8��AVTdt�-����Vl��󫳫�s�������^�ӣeYE�!Ռŝ��Z[�5����O��x(<���NI#�k
f�>���ö�-s���-�B�u���Ȣ��·<;��]�	�KWb�<�4�����.�v�Y�/\✔ۜJ���t��TLU���j�͒��� ��I���۪�b9�0�/�Db���M�*z1փ}�:���DT��������:��n\����MD�O\m��Gy��`3ڱ���	z�<��U��s���ˣB2M��3�������u��l�q,���g��w.H�k/�x�[F"�h�V��q���h�x�q<pE
��Y�Y�:J	��,�yź���NVE�JTP��!�����l�*4��3�Y���@�L�{e�(�;7��A�4�<��3��ӶΑ�ޥ]I���R�؎h�*WI�k\g-VwJr��r���w���2�-D���d�'̎)�~���E)�*n�U�ۓ@B(�͈Iq�m�����j:��S��yr/�ٽ���]�iZ���;��"���T��������!���T}+�����]yB�����9
̼�Z���x�gt�7rZwݡ��}���M!���ۙ�wlD��(�����~(��,6�<�^H�cT���d�E..�篽Z��k�j^<|�f#5-��2���N�^�e�L7&����PG<F�d��oM�ؖ۞ɇM,�5ݢ�hg؅���/#*%u��Z8���6V��dZ��p��&+��&髻t�=��7�qG�F�N\_>H�,�����G�����QJ�`r�°@�)HӋj��Ҷ��f#V��=W/ݙ�FdTM�E���/�1z3����dz��8{��j�M�5Q�����&X����h�dt��˸��d�WT�5p��og��g!�����Ȣ��U)�o0r�ƛy��nA��Ư�DGd�c:�u�n��qc�qe噤��G�|7�T�"+x^kse>�.�<�XlE����اF�im���ݠ���Z��9W�{���1z^�#q#-�o���s�`�z��7HyJ�)���ॳ4�;u'Wf�PdL5(�#�˓-�������ƶV�8�]�2c��Պ����T(�~�l��0��s#��r�0����u�k&���C�[cw�W�0�۠/l��"���������L��ח�@uV�5!�O{� N���m��$�j-T�kk1L�]��&���觅�m���uE��Q�-�qgnysӹ-V+�n-�C��T8����ȫig��G5]�w{�s�0���E&���G�]In1�}���EqE�@�7Q�5��f�	��*������fu>g�4�3���5�һ+7��ڇ{%X��ףs�ٕ1����q:۽/|��c�#�=��|��`7��Ʌ�X;��2+�̓�aĔ���%-Y�7�E
i�O���s\����C ��>��V�ve�#�WJ�S(�dz�V�n#�"�]����d��^^[5R�d�X��R���J歌�UQ�	F�<�:�_�z�f��uľ�������٨�w�0�t���}�:i`��tV�]qz:-��oT��h͠[IU}���g�؞��t���=N�)勧���#�>�<f`݋��E�ypFcE�b�4'��%����_8�9��Ę8r���e���]m[��u�wv�ͷ�ޝ]b�4Å�Kz��J`���=�sQ�&�s��LU��ļ�:���I�y"�G�p��v����y�{`�yn�2����Q$��cZ�ܼ$���c7n�&�/�[��E�2Z�%8[x�:E�wHQ��y׆�f{�Y9Β�an6+:����V��}��� i��|�����+��+��(�<rS�:��yz�b����̻-4����P���zd{�p ��.nv�V��m�ˋ9�.��Ĭ�2�S����2�藅�53�U���=1��Uܮv���aY.
�(X=P�l���?�����M̸� n-f&��G�6��Ӳ��s?:�U��X��ć`�E]�WR�� L�x���JбN�#WRc�?��&:"�GR4fGLt�Տe��l�%JmR[����/�nw��QF�Dᡣ�����W�=]~���oUm-�ZG:�$�w�N5ݓj%u@N�0��+�Jw)��]2�$���8J��k.�
`�	��jt�"Ks���6�{.Yy��8򯀋I���u������)�!b��`N�f��oj�ٙ���^��;��CW֕X�C,�G8��lXXJL:F��n #9��ټ�E�.V��7�� :��{�b�݃��@o.�� |B��:�����%j��-��N�q4�c}Kj��ܾ�)Ы���i��n^f\�4���u���[E�t�;�9fTZ�4���-gG1]����x��m'z����*j���t�ː�.����^���(ë��pGq_~~���l����8�wM�R�n�t����6q91��Թ��9P<'"�Y�Ye�Ц(۱uj�1��� ��̹�q��I�i!�t3j�v�*�S��@�R�r��Øh;��pU��R�
��N��A�JXH�Qā��\�YV�ŌaE&'��)�ebx�0������}q�%`F���Gu�[y��I��5.�kh�8Z�����N�����Ur'0�C:�2����8�4��k�;`�n��R �J�-ۣyq�������s��i����Z�E.l9{]Gk+����b�©s���̠�t�7�im8)�Z�o�uzV#,�;�1Ь`�ۻ�y[�0��eڶ�;���q�� ��ҕ(ݕ,r��*\�5(Y��!'����+�ܨR8$!���h^��@���e����Wm��|��Z���Ђ-w��,ƥJ��k{�Qy�cg����jEW��l��\�y��7���{=�yOm�}<�{˅h�y��3R�FO���L�?$���R��󱷙Ǵ)��%vd�̤�.����<���nS�Q�}�s:�D��B�������2<�>x��=!�׽7�p�T�^T������J3��yoFz�}�ڗ�<�>�u̫I{bшx�m��Mq�W�4=�ϳp�y�{דޅ�f{N�n���Y��{v�Ir�ћ�*���(M �����+��'�������ԏV�X�"�����1N��	N V�4�z�w���7�m�h9��#H���(���z��ޓ�ٵ���㕱�i�k�1�ݼ<�L^3�L�r��}�q�_rf�X��鯡ٍ�2Q�Sҳ�������To>}�v#d��߉��:�je%�ly�s�Xް�h�⤍�'������&����#��9*�yJ��
����p�YP��xI�k�=�a;��%�B�ݷp)���IZkP����1�`�A髓w���Zv�y]@Tٍ���ם"��ѮdKb⯷A���е����vk�ˬK���<�Mxd#FN`X|�6�5:��X��� �Lr.@k���G��ke_%z3�D��f�mHEۋ�A��
C����%������
uF9Fx���5��2�S���[p3�R{7�7^��f����mn�+.��b��4c��Յ����$�"rf�ޚ�>����8��H뮚��4�L�6�o��}��F�9:��x{����So]�*P;e �˛��r�Y�l�;ˋ�
�*z�Nh�SPw��f+GQu��>g�^6����|@������՞=�5������F	��p����؈Gd���к��� r�6]���R�d"����Y��z����B�͉�����e�,۝��:G'Xਘ$服��nO_-�CØ�#��Y1�|�c�/�e˫����}��ٜi�vr�'�k��
z//������T����݃���}QE�oznT�FT��X���Z���P�B1F�@�;H�aS0�(�Փ�,�8qL�	Y�Qզ�ӱV�	;�/9��{rtՔ���j�s�R�-���bP�#�(�U@�1���C�ݙ2r��~O˻�N�|�M�]]f�aZ��btf�ң�l��l�[}Ӿ�kv���唹d�wS��F��[{2��۲ڽ�k���ZDa�8}}�P��g�y���h|aϘ�ˣQc2�Y�����6��Aan8�Rv���H_q�5��	�
�����ۇ��۽LpF�s���׳8��;�3`默��*���n�^�y�oC.i�_NM�^�Q�Y���'�o ��[(�r��͜��C�k��|*-���tZ�R��Ϻ+��B*�[���g|wkس����z"��*����n��DD���zf�G��ZUd<���'<�q��2'�j��ɖu@d��d���^����7�t���ZL$<�.�$0n��L�� ��X:���NUOP0�$�&M�0�՛�x��s�����'�==P�@�}X���eвt��u�$Ru4�y�Cl�4��P�7��m�ٵ5��׿�m��*nQ�Ɗ���=���Wod�k!v�84��?J/U��5��:.n�,����84�ڗ�KՒɘ(���+I)$���r}���}>�'�Z�6�ԁf��bBi�2d�����	8�aL���I�&�\��[�9�����l�۴<�0��ۢy�a/T(y�Hq�-U$3�X�`q���`)oT%�:�-�g�s�{�xHa�L��@8ì�d��L�
��Hmڤ0��=U �L�m$�N��k[�mY����[߭�e̚�=�u���&P�h'�r��fXm���K�,^��.�(�c�m�i'�����ε�{�!�̘H�.�u�I�T��e����s�,�!s���9A�����`Sl3Yϴ�{����s�����Y!�W��Y&�:�i��]�y��P�d��BݢL��I�|ov�/����5�{�.�<̤�L<Z�4�k��M2W*M �P.�`e L$8�i��!Ć����*����s^�I2�Xt�HI��T$�P4Ɏn�$Q,�$�^�I�����!��o�oW׽�{>��e!�����a��d��6�<��hCi�2)���Bq�ɍX�|�`�H]�`{�ƫ���k{}��]�`g}D��ć�0^�,��:�u��u�`)& ]&Y7j�l$Â�i!��,�_-�}�|���YH������)J�$a>���|�m "�IZ����g0�3�&�4�F�!s�j�O�Vc�t��p9�h�}�G�=�l�9�&=�1}���b�6�u$�څ��q'f����$���L$��)<�5�����͸�������q ��'Y���('�2L�L���j�u���ԇ���9T��s����_V�5[z)4�$�X�-�,�('r��C�2�P�'��[z�:�,��B�@�q�C�mkr���a�6�y������a,˲i����H\K��C�0�S��"���Hz��ί��~zdY �e'q��q��whCL�6��Y�S�@����8��% �It�`r�ώ�׳�z��:��w�$�����8�a	�N!��m	��:̰�� �%�58�0�{ޏ��n��s��۬�(71d0���
�Bm�}T7z \�Ra����k�Hy�a	��U)2��B̚���Đ�h��;YI��h�a����8��Cl&\��a����v�] m�;���;�ߨƽ��{޼�.����
d���$�Lz��m�`h�lL�y&ّ���c�z�/��z�'�+�߽��X�+{ֻ���{�	t���0�CI:ɍ���*E�k8��d�)'XY:�d4��Bm&+����w�o���^v,s������t��7�q����oyL�)�G�]�t�^�Sz�Λ�;.Q\�u�H�����'q�ކ�S�uu�u��B㍹�e��\r݁�u�� u��P�$�],���I������$��Rj�ݢu&02�h����uk��Z����q	ė��Cn�M!f9P&�2�Y��I1TP4��$�%r�i��7��i�qͳ�{\��0݁ԁvu0��	t��&Xm!���x��'x͡
�@�"Ƞi�3��ν|��ŸI�m���a2��T�$�<��I
�Y2�y	�6ɳ�a2,&+oq{e�;�����d�&<Z�8��yZ�&�d��k5!�i�{PC��2Oj�́�T8��&/D��s޽k�7��m'}P7U	kT$�,��I���bCh.M��Q'Xz�4�%�RB�T:�Ԇ1�z��mf���}'Y��8���B�Bɖ���e%=d�z,�(&�d��������u��g<;V���l�����i��"�ޢ@�M��d�),�$�T���d���!Gh�d8µ��m�;oVyl�:��IL�Չ)'�t�@(7S���'6�!� u7M��d��@��r��a%�Ԑ�o�^�޷|{^źB�'��Y �	<���!�m�o��r�C��R]�v�,%3hB�Q8�*��C��?g���_�݉%L�~7��h��bP�\�W+T��2��4>�Z�>��<�h���v��o��m�o\Z:�/���.�K�4aR��\cX�s�����y_!,��d�C�7��N m�%�$��jK�v���q����F�I��<�[���������ַ�Be���E���e�d^ցē��� h�Bm�Kj�.�Ĺ�$�a�:��Y���X3��u�w�ψafK2N�(B�P�d6��2[����m�%��I�E�e�XM��S\�0�_=l�~�ل�	���Hq���I�U%�RB�i!d���0��K��N2u8�3/�o��l���r��{��]��	I.�=�	�B�*H@�2�q�@�I�I��HV�6I�L⤚@�w��Vչ��|��"�<�vM�/��:����2��Lj�8�ުL8��i�RSKSi4�s�:gݽ��{|��I��2�X�m$�m��.���PCL�l&���@�&��!�)��*@�Ӭw~��W-�n���]��'��y�Ij�2����9oTǼP��9;���j�BL׸�/��̻���m3ETy�_�tI/��2��
��|rۡ�������&s���sWwz��,ͳŲ���o�rw
�JS��E��S:�}�R<#�Eaz����b�S
�|���ms'1�2E��_BN����VV�l��ˎ��2�U�͎I�W���S�DrU�Sz�F�U�C�^8 ,6&Nc=�qU�Xj�)I����:�֙��k�i	[xͅ��gGwm\J�x�x��/�N����e��uM]p������6S����qƘ�aΎ�͛�5����º"���w��-o'v�RҨ�yp��6�Xյm�`���d��.G�ƳN���ۄ�k�\>��tJ����^�Q���|�C��P7�]�����ݴ�$�� A�h>�ċ����X!����2M�5�׋yA�Q`�wN؍\�r��V�Vf���%9?U}ZU�M��"f���(�f"έQ��k�k��qu)8ʦ���7��A�i�Ղ;�Gp*%�J}��G���������(��k�,*~��}�ԝe(蘾ݞ"-��Z^jX���;{P
-����:w�ݗD�WjK�מ� �X�rm�
�6�כ�Oh�D�N+�Q7��MV""V�=��N�C����v�;�A��QД\E�|Tr̔!���O+�<���A�㼉ޭi���
���!��F�i\�(���nx}/<W����n�S�3�+��݆�$*vL.�Мz�{�Sɑ ��x�0������\6����W].�&t?�8�ٷ�{��@.)'rW�eCw̓t�Jus���歙�Z1�����M����9&���eìA��3 �L]�  dݧ$��`��vÏH���=�8h�Q�a���Gt{!�n�c/��U�&��DN����V;vɬ�����0�W�[jq��]�����As#:�6�
K)lt�{���oPY�?t7�-��:���Pĸ��nl�������;*�(�uw��r�Wdsz���Iu�V��w6��4c�U:
�"K������+ZC�ӆ�q�s:��#wrJyu|���e��rp*^�xwǤP��ݖFv,�OVuǚ�i��ʳ03���4r�*+���+'��ڽ��l�l޿���LV}��^B�j	��x홉ܘ\��r��t����æ�⡂bʼ�X����JBJx��dc�c�q[�R���R&�#����{�Z��)�X������1��X2�6D�&�9Jf6�]<.�S��`������#�y��41�8D�O�\�ea�Q�`�	�̈+J�Vnq�6QJ�
�:W�F��XnQ0�Q��E�WG)�B��m�'�2�V��ie�]ǡ���UA`�rG@��|恏f˼��؆����HeUֻ�D�N�@�"�l�5l�S��h�1](��SrQ�̔�.K9���QӜ:�֛e���tm���(�@�e�Aٝ!�u�:WY`VE����!Y�)J�c&ʇS�X�4�$\�Y��7.;+�@Dۅ_[�*��E�����W�t.��(~KۡUV�V�7d�[��-�[�\�&M�#���eD����^����R���SޡW�����#���MI��{�fUu<��Ƌ>ݴ5&�ª�
#���f�HIr1���DDA�����4��^�krZغB���%�r\�
����$[�Q��:#!��ڕg&�jrg�6�Uy�u��Ԫ��������?i]Bz�{$���,Ȉ+D���՞�T��Ub
zh��W��5�C��Ь�e8�%�4��b�7�~ku��C+���΅n�Of]�_%�����\0*���,%ܗ/��z �q4�~|p�b��\r��g�G}��C�o,�+��B8u�OՁ?V>�y��w���f�C�ٵ�.��<oL�Z"��X����-y:�K/E�#�O'(�o��T�ϸ�Jd۲��o45KpT�vuѨ��;e�Ď��{~�@6r<Y�	m��x^o�W��6rj����7O��Z�����t{���ӹh�����}�Q�P3V2iu���z�;:�4��(�+��|�񼭜�{�6-�:؁�*վ�kfP�.�u_h���v���w[d�6ε�(���EȲ����O5?xe��QQ�ǵƯ�]'*U�[�z6m.S�����P<G2M���d��{�0[�0-��8~�p�(D�^�J�{e�Ë��XG�N��T.<{�h����ųxʽ�ea�s��1ב���Y�Ǵ�
7�S��Op��J0�R2P9
$άķg()�D�0�P��Xz�`���o�ū�7���.�ó!�JG��w��TV�{���m@��&��e]>F*�t�+�'��o.��ON�:Q��tQs7�����z��(��+r��@�s�;<h�v��\R{�3\i/5^����[C��P��6f_n�*L�f����'Đ��ˌ}��̸��܎�Cd�[3�6Ko%(ʃ0q<ʠ���/*�㛢��֫O4��=���ROy9���0e����w��ˏ��직ƽox�V�⥱�����
����*�����s�����x	DX]�\fj�ȓ�R&J���2#g�ыg�C����r<En�%bt̾jw�r/r(ˣ���@s\y,�n0�J�m��d����(�`O;Y�>��>r*jߟ��j��VXg'�<�
Y��sO��W���,!fX����æTmp��W��Z^�fW��:�r�8���[��v�E�|}�g���L�P-�_����Т1��-���*��,��h�]���ڽ��z-
��b�e����z2��bl��p[�O���K�jH�+�D{ނ��e����{ݰ��[��H�����Xep����HJ��K}���];�.r�9�?,$�^�(�n�P���q�6Tn-��^=DZ�\)苚Q������:�g�2�aJ緎�����|�x_aܘ'p�ٸ��GR���;�nc�6�OI��L�����p���ǯ{|m� ���|[�V�D�l[�G�W,$��l.z��Ӿ�U���X�SC�>�M���Zvr�;3hsm�w�ً#u��ޝv���x%�v٭0���v֭�c��.��]�U"d{O�&f鲎�ڔĊ3T%�h��jew\�j���J͖Eǫ ɇ��`��͢�y"���z"�.�}Ux�͕��Wҙ�kvE�����r|Sr�n;װ2*�S�����؜����w)��zڠ�,�HV yX���W�t\���,�4�=R_f�yʹd9�o��XZX5����AoA+M�����ݭ�[R�� Sgf��#��Z�{�#uV[Ԯ��ӷqUQ�DE���u�㊐�����Yt�E[ޮ��TH1���h-�;�^j���-����EggIѣ��*��f��)�k����t�����o����6�3{ W��QIQ1�z��e�w�j���>E�q�v�Uf�0���.�S�dF��{8�)a��c��H�E}���4�jo�ځ��V��Q���O)W�^"V�J�n�śS�d���3Θ��Q�#@=|�e8ܼqDB9ia�����;�W*��؛RD�s��5���wQ@;Ԕ��$�d^�VK�W����ԧ�{�Q�\�z�C���l��U�D�F���{�x�V���҇xY��$28���5��G<�+�k�=P<�P�C��V^6��:��X��Ԟ��^��Oa�a��w������M���Μ��#�o�\"���2Mj,̍t�y��z]������yʚ̱�aBs��&�ϵv��M��:�x1D�5l|
���!!�[��?W��z!�=�o��Nv���Y\"��2�=��uy�Bzڣؗ=�������/���:��a�uZLĬĜ�~ym\)x�|�G�|�39�1����E��Ϊ�V&+�2i�@e���-�d��}Z(�$`�)G����X\2�-��y�~�����s�f� �v�[�/ˈ��3�I�s���&/�rѯ^��W��/�Fժ�v�;^�B����ƽI�Wc��ԫ��GLN�f�q����-�Y�a\.+:	�1P�9�/C��#_�s�Ӯ�����:�ȶ+lA�ol�'.��;��w��^�8�C����q��s8l�L�v\Bh����SwC��Ҡ;rV���G�S�A]�te]4�ͧ��ɣ�l�k�h՝�x���#��*V��0Z��zyȌ�ȋ�ۓ�-t�S]/l��ؐ9r�h�,��`}Ssm�^�f�AB���'��j;��n����L�:��U�i)�}���a� �������K�O,L<�¬q����<mn7�:�j�5|}2��"�p�#�G���z�'=کo�x���{�N�(�kA灗y��xݺ���w]ev2��gt�1m�ĝ��w��e��3��ԉ<X�<=��;����ktlR"�_���,�C�,�zX���s���eXΎ8��kT��NЃNVoD~ܽ׻��]I��U�n��ov�R������6˩�>�8�OU�Qd��o��iFu�Wʷ���c,Μ���U��̀��}�e�S���6���Mj��p��(�_A�pg=F0&�g�OGt�Zaa՘Jt�z.�O�U�L�K[q��\�8���җ;x{ lU����5d?o���g9J�t�Ty`ɓZ��5=�:B�`���i0�yE9R��H�&�ë����ue��QX�E�E��v��x�`�(���3z8�����I!�n�_xC%n�q��J��[{��
K���WR�����]�)ZO�7��7�6�о6�^��>�R���V[z�(g)?}U_UUB[r{�;����@�mP�v��5��<�9�m�Y�^5�k��Q<D$h\�,Xr/�xc�o�}^r��;��-��,�R�N3x��Y휃�"z��cv����;�Ͼ����n�uE���F��ٲh�=l�4���u>���e]�YZ�����IL���c:۞�]��B�ha�J�I�ͽ�(qh��8X5�ؘ�(@���-�r�G0-�ʱˣ��K�c##M������x�X	x���$ֵS���x��k=_N�n����,�˖U��4�(H����V jl�h���ȵs�q�Uw�ێuť��x���=J��v$���J?J8�/�Z���4\=��fB��k�f�,6)X���n�d��+7��s/HܼY&Y�S݋l+����OvIEbՇ��J9�Bd��j�DHũգ��7�Φ	��mØ�y��q���lf:S0���e�{&��S[��*��.+0��}6a�+:�a��Y�M�/��n�N	jTK�hΏ@����GB�*�v曷�n�I|��;lh�MT�uk��¹���아���$�Vv�۶��$ņ�ݱ)�H� (=���.�c���g�(O��|12�$��3q��{�WV�*�G�VR��=���sR�k%��'#F,�O0��`����j�c�q$���Տ;�
>t"���{������b���������>�g�X��K�f�� �ǐ��a�L�h���t��#v]��9v�dF�
d[� �92+�Y1[r�D�"ÿ��-�gp
���Y-��U�-a�W�3>,E*ɘ�4o2���ȘR%hY��4���3g/��'�E^��8�/ �a���8J�boo% ���ܩe� ���%-n"+Z8=��i��Kt��)-+�d�������3�'&?�ެ槩L�)J����*�4����f�Qq��΄Żҟ�5�:�t���v6ŝ���ݥe���@��W%S-�̩R�F2l���L��ǪI#� �7�[���D������D��]1��߿��Z^F��R�Ċ��0�$�)�3%�H�Q
��2&w��0�)�S�ʑ5\�L��F�&ETZ��l1p��[dy\�*�L7�c�
�<y�H��{�G��%UH��������^r�	�l8�e�in�!�O8ԥ�D��	:�����z��Z_���蚧�!��}c7�C���I�\5-Mr�^��w�v}���0�G�.J"\����`5�a���	M��+}��?'�R�Ɏ��x�q�Z�3
*�8�KO�����h�XUŉrO}�}��PM��d����R���1j�J,�,�ʀsY.]:6iqv�ڮ�j*9#��@�w7<n��~�\n�s�w �!C�[�C����N�������`S���{��s5.N{x��Xf�g\UT<� m%eV��;�H����u�V��۫��s
M�Vf�������}\�V�{dsd�Kz�����}ֱ���;| 9m��OBڻM+Nn�]����ȟ{=��K�P\����} Rz��Q�'8B�#N��Q,T�S�}c�繄��|�L�35�լM�����Հ^|� l�/ean=U��I�os���ٓ[�1،�r�Urt�6l��c�h�����n��}�]a5�W����x+�#q��ﾯ����u7�Ϫ���M����0�{j�.E$�|׈��3tt�9R��v�o?N�W�NV�s�A�!g�Ou��fv8t�)Ӑ�E^�+��V�:bQb���e�,����z8SV+8T�6��q���חqkx��.�C
��ؚg�st
��T�@p��#D�<*W��T�1
;�����!b�-�x�tI���Bqb����Qy�%7�F6��eE�É\��r
�>c$_j΃������f7V�x�AX:����HK.^�^�)�\�e/B�2�=�ب�)�8�}Kt6o7s|o���JB�NO�}_}_T{�{7�+K��l9ʄ������C�Q��zJH��9DL��ڭ�W)�����l����k�XN���6g�D胵��W�n��2{p�̣��=9�\�k�S����.�(o�5���"p%�x�^y¯h�ʮb3��i�����s���r�Y�sk�Ӫ�N���5;��A^�
�Pn�rP
� �,�N�����SkId���W!�'�U�]I�t������z�%Y�y�p�:��:�ޞ%��)0��'��+�J��e�gU�&��K��B�.{z�70�i���.�Q'1Wsʑ�w�U�E��3)K�U�8��\�_z""=#��Ú��rP�F*:	t�4yX�=mf�����MA?5�Հ�.��P6�yZ�:�FzM�X��׉Ҹ�Ƞ�\{-���M��Ő���=X��u2ZW׫"����W��R���k�Vk>��ʽ����y���ؗY��^�!*5r��+7%0�����T=�\����C�#��!�b��9��q��U4�N��Z އ�K3�Sۻ�o��ߎi�X�5n�����CI��yp���ns,����=�����C{{�����;ɴ�ŖTȻ�j��;�Ų3ڷ�����`{ �a�^�7XB�I�9#(�;����ٺjc�[.9���{�7��ۥX�+�ogI��y�9+��]D57�5v�-5U\��݋�,����F�q�Ps8�b\7�<�4�D��ȽY.�;��w*󻸼�qOTc=:�2{����.bn��=Ω�22�G'#�Ḅc��d�`�y-�ܮ�<B��Gc�Z�V���,U`�˹[���t��w]�����7���e,@�~W��*&��1��y[���ba÷�s9���.Z��'G�<(�s��~t�k���<����k��\�w�;բ��(��](�
 8�]�+0Va��|��@
Wb-;e�t�\��^Z�
$� �2jOf�>�4�@�1o�`�n9vU̲�I�!8�[�7OT�l����yD��=�z=J�~le��ܫ���7�V�N�|�>�8�}{�eӒ�Զx���X��g�c6}w�H����D(I�刕�Ⱥb���Oẋ�s~ο.�C4�dnιƵs5ݮ�kk#��9�dۻj3���S�z�^o�Ϗ���8�ۄiQ�#yY���ppfZh�p�rSѻʅ9�˼0uS����D"�
F�i׻��P�Z�b�z�: N�b�����Xz�������㋆��ٳA�b���hi���k�Q"n�6b�����"�k.��D�����4sOs�ߧ��{%z��#���Q.29>�D{ރ'����u��<`A�����L�EWE���D�א"�\��"q�����'��
^[w�*cz��>��U@,U�t�z�ぼ.�ᅑ��tVjs���55��0\�{�gFtU����p4��#k�g>��Ӵ�܆Q
��Ы��er�3Bdn�q�a�ڦ؅�.���fz�v��:�v�2��n�"���W� �ۉ�ͻ����x��Vv<wyۄ��7�
��*SxyV�rj7z�)���#V��(�h�X|�`��Ѯ����(řwݕփ;����v)������;���&Χ�Y�9mn��S'ζ�r�-����7�S����U����R��"=��7o�~�>��#��=�٭u��AA����^����w{�Es��(Y�b��t�5�\E���)��xM���P�.D�Bq4�f�)R�_�Ѳ:�i>uPQh��Z3�'	�B�s{S�}��]Oޡc���	����������������j��1���%jXc+{.�5�{,���1r;B��b�`���s�2&8-.��Y>�C;����P�a�N,le�{NOF�R�K�ަ��
jiP���O�=���1U�k���|ɕ�]o�`�2�|�2�X�~{gE,>0|[X5i��UL@T_y�VL�R�4	�FScg�vp�R���D\���3S�|���r��>n]����m��6Co���A����T9��:D�96�Cbn�4n]9V&p�|�����]�w��TXK�._{ޏz!+��wq1��O�B�Z������t���������r0��z��<�`�T���u���ҥ���a�:6��EJcF˂Q�'FP���q������t�=� �'p�b풛Ӓ�ێXl �-�_	������~�.���W���4s��4X�}���F�-�#B���:���$/�[�Ze_=X@B�h�k0՜@T|�:����jV@��Eˉ�5S^.���R Q�S҄��B�̤��e��P�Zr��T�*���ea�g��a�ŤV�f�q>�Ц�[E9;㎘a��i�Pӡ�������soÃ�҆��4d�Z�~�J��%׸%�a)�rx7`��.Qu�M��ڮ��]W�+/6�Y뽻sW��*W�v� ]j�tj�*d�{`�؇)�5{����!zDɷ�g��@�C�﷯{�q<㜷ô�n��v}��iQ���#��[��re��������K��k��9Y@w��H�DhCe�g��\0V�5��a�����ᢔ0a4h��|���}b2m�L9Q51f��D)g]���\ח{�oԨIj4lNc<�s3���PF�$eCLg�:k��l��<"75����+ٯ�S�Q�0Y84\8�<����=��m@>��g{=�"�|������j�XC��ss1���Qxִ��S����l�f��AD�@q�7Xii^<<�V��Z��*���QR��Z.lTt����40e +w�twhvۙy�h�z�*�,����J�:5�p��� :��3��MS)�lK�j��[3��К���a����O�N��J9}ؔ��/7�<������J�R%�geY���s�\� =��_,�/|����vU��kxG��v'v��$�W[@�F��� l�rlf���=��,�b��w-����"�b�fj���3"��[��沕	ז&�@$F�^��2+T�{W��[��4�B�n��۝w�_2Ti΂�r�A�qr]0w��f�1��tE���Q��Soa LH�b�Ge����\JM'~�)�{c|�3�g3��HѪn�+���w�J�添[;��$�V�b�K�WS4�W��,j�h�	S ̩��j���d��E@�é5MP�m*�T6��ߵ�n{s^��JtEW���^�\R�����\^V�u#�M��uyj�]1��B�a�J�=X�Ú��%R�Q�����zi$����w��.VeJ*m��&�QaTaޛ��6�nޣ� ���iN��Z�ͺ7*a[�\���n��f��!�2��%�o�;�}����w+nh�q��N�([ÆTsGY�.}�뺒 r.mYZ�p�t9���Q�wb8�W���_f,�pN�4ƛw7RD�u�|B+J�}|e���J�B���e��Ω&����7���n�Wo�`�؛���CN�]���G%
9X��w5s�6�YQ�-䬩N���Ȳ�b�R*�[}m�{l8�E��
���pnØ�>�3�#A���o����)Ec{�+�i϶-�PXP�
�����j������mX�zv�%�ʕ+��eS��lJk�H�V��bT��XL�"ff2�o�uL����I��D���@�S/㻳�3��{X%�D���:�-#-��ʰ�;��a0�M׮.r���д��B��G۬L�s��V����UJ���7"s���jIZ��7�q"�*�]sSCs��TDD2���S\�����g;P�Ϸn�x�i��ct�"�57��Q�8����R|��z�[m�aL���H��a�6�f���B���V���i�I���m���G��ߔRr���}p/e�Ǚ�s�Y��Ƣr��T$�R�]�̼쵅ㄷ'���� �Kt�?*�������0�USb6�ȃM�L��S��=�c�ѓ.<O�����R8/r���j��\Ss�[�r�7�E���ƛ���^�W��T]��׆�����Na�y���j�Dm	^5��]z�R%2�ʓ5�x�~�3W���y�}ٲ�� v6�z}���������*`x����m�hW��`����ā�t\ ��3��~G�����o/V�< �4�a�+���Uq��*YP�\�/��u`��򒁍�<=����y��[5�6z/J��f��+>�R�E�N��u����32c+�!��׹>#V��r�ǫ��0h�RV&
#�����Uz97@�,�B�40�Y0t�u�jo�P�����ORU��!.�E���}�EvIǵ~t:�U���B#Ɉ�G��i]��d�)�$<�3Z����ZŜ?'���.������\ �&���}�W�5�]�o��u~�!^�0_R玍��!I���VJ[9���$'�����j}U���=Q���Pօ[��Z�L�o������Ts��σ����������/UyQ�.�Q�e��	���p��"ƳX<��еbT��/�}�¸:GB�j��C����x��r�e9�x�\Z��SN*Nɓ.w���WC��ļV�
-�b�p��~��j���F�\�Z<�:�:��X��� Bx�o�s7�,�v��>Z #����(� �Qњ@�l��[y��O\ǥIr&�FH�١"����O���i���8���n�әNqeN�Y�,8��1Z�����	G�i@=˹J�>I
��W�?�W��_�]��Ps�Z���ٖih����c�KL�k�	wo���������E�m
�~u/P�U�"V�'��K�/��DYv�?�"e��U��GG�������Ճ��Z��co3�'���n�l<%q�(i���z"(V
����X3�a��{��;����G��xX�-��5��д���I�\���z��^s�0E�s��>�f`�}Na:�ɩ�SO!���8��;Ny�1uq�Eza�/+���F���3���ρ����~�n����@Ma5cyd>��-}	����:���љ��g���i������xd~dS��Gr	�ˮ�X�F���[��H�����%��^���n<�`Sؼ*��tk���r�A��gF�>
z�;��8q7�&r<��//U#�S�p�y�ޤf�7;af�(\��i�r/.G[۽Ix����z8���K�g>�eGץQ��$i�?W�������Ϝ]l����j6�RAMʉ2$Ϊ$Q����1<�}���o2�<�ѩ��u�t�D�k��a�30d�o9qU�{ޢ����"�*^|�l��KM���T���ξ���4.:0X�%N>~:DÆ<��0�j���r%0�`*iu3F���ep���4�B���O��d�2�\Y�ux�η�����v�ʢ�ZڤL�0Tg�+�JQh+��9Y�w�ۛDt��42b�F��(�^��<�=~���	�
��T��U��,��g�����
�Ƕ:P	���7Nzl�-���s>i�1�Z�l��4��Z��c����oe0(��\��x�ܿ����U[�"\>�����A���a��Q����Mfۍ��G�&�W(`9��'7��ge8��B�yj��WRQ��VĂS�G2C`�r~�����4��޷fׁ�D?U!W}xB��;ꮑ����~{뎍Qu�6�|����\ݸ̾w�+X���\n+�U�jÛ����<�y[.�H����˕8�\�ӷ����j��P%O3�SQ��{�s��*��Q�k�0x�2s�)S�""t�29�e���=��*,[��
�7���	�}�Y/q���U�w֪ؿ%��"�c�< c��hKU���z/x�ﮍ_��ԅ:�C��2���rg�(H@<���9a�frgB�0
��uε`�.�ʕ3Z�P�>E'�mC�2�[Q3h��k�b(O�®O��;t7��_E¬�=5Y�ā��Z ���xvmi������4��!8Zn"W8k��y�����0���N"����;�b#}��;��qu,�:4_+.$�A9()
�d���8l,�Aͬ�����qNO���s�ι֭��]w���fs6��M�Z�ꊎB�b�	���U�\�ؘ�k���(�bޭ<��ea�gy�<�a�=�n��*��k4����"١j�Ƽ��;���,kVM�x�����pX�V4`�z�B��Fib�,@X�2Ó�V��,�j�ܵQQճ�z���]*�R�b똧uKy�.$�tTAκ�T�C�S�Gx�Rr�@B�4f�ʉi1�e���� �@�u�����t��g
w�-�N�G�pzx��!M�w��n[<B�h�=��v��6e����;�dU�|+@�V�{\��G:���8�QG��S�_�	TEph�*����ԧ���h��yu|�����E{�R��EE�N��r���z| ����0��YS��%<�8=�3���C� j�T=��p1����1�8�����|�����Dw����Á:�3��V
�xs�Yj�@L��z�q$��ա��ك73T�A��:�:�U�WMA�<��gǞ�\�Y�N��W�a�����C�6L�ߑњ@����ެ%�y�����0q(\�P>:-kt�!Z�}�ʣ�Z-|j�u@e��y��Ю<+Ъ&�&�%F��)=���.�\��r��r�����+?hB�0QӃ��^��-�ғTۿP��i����l�m�>��vi�W��
)�_{=}ވ�i��6|<�d
Q��3r	ï�2s�d�3��x���Ɋ��g���^���]O}h�c��G��h
>ܥy�J��0h�ʳF�������L$Y�/�D�Z�q�}$�4��g5����>Wa#��[�-�ԩW,pF�����R�=�o\|¥=�C���x��j��*Q�h�@dыc�Ƨ諭��7'�&��P@����W�3+�V�`�e��f麄���W�0�`����\��a�8�?j��蚃�gi��f���ut� J�1���3����ڿd��[��|��הZSfū��<X���PSh��Y(Ռ�K�ç���Ll�Q���^ןF9>��m]SAM�T������Yg��̓>RXU��C�f��x��P�����|���mj�w٦�C�x*�,R��6����xm�"�Fj���^�=,�	�;xG(p��O�88�P��Z"3�Sn1a����b�.�w{�� �8z}=ʘ"�z��J���v���E����D�?h�q��ƅ��Q3�����zp�=Q�rf���|�j�CL��%�d+/W�$_w%y�㠒�=�u��(P���rZoA���N��$M�?}U�U�8��ү����� �c���=��U_�z`�,��D�P0o�_9. ٹsLO�V�p�";��:r�C�ΩU��>�D�L����*OʱŴ*
�yUκ�Ү�2:ˮ�M븎��2vz�+wF�~���\'��%[��ϲ��yp�f��@XY�D�U�852(g��=���wrOb
��r����6�(k%��t �[�^>͓7���*�<.���5�8N�áZ6����߁�WwK�Vv��x24�1�@��$y�(ג�w���t�����#�ʑud:�jqk�x��Y`b�se�x���ր,Xc��"�����{�	|���gx���Jبz�{�β��k��� �0-�'@ґ��3ec���Q�X�6�l9G��+,�ޡ+���-��|�򾪧��[�L?ɨ�DB��kMEGE�Ut�/nL93s��q|�����2�J�N��!َ��u~��VT[��˛�}�Dw�f�����V�ڀ��M@bk*��a����{P��<+����1�l�lUH�U��FnL}^}�Be��e��=�-�lfm*^��AYW^T�����AP��N�2IKA�x2aވ��5W"q���Ñ6�g&35���L�U~8<+��5b�4�f�8b����� $g�l��C�Ｘ{�h�60:4*�QV&>��zwQѠr��.�[@@}��X��3�
��j�Vi�%~11~���=��^xŪ�P����S�~ѳv�)���O�c���?�]�a~ҫ2�(umJu�_r/k��r&\Y�u��$��!f�˜�'KMN�� ����>
�0.1ݸE����·�2��.���������O����l�f���g%DvA[z[˴y:�:Z5M9��{p� 30����� �W�:�bS:��+F���ufi+3"<��H���$=\�B�4ފ����Z�6⣆��92r�M"��H��V�^iZ9�Gv�:�A6�Z)��]&��\���.7�Egh]DS���4)�&�Xg0&�r�Io,=*��!)Ǖ7-�r#�o�1@*�V�Pu$r��iι�`�S/v聠l�z�*�|[�2�etZ��L�L��<�{SC1�.�����Fzִ76YÛ�ܣ���iQڳ��U��)�[1���}����]�7q]kǟ4��x�ֹ�v���IS�s��Z(,N�k�T�Z��`u�5��'Vm�U�qȦ8yZ�.|Ĺ�)k�k-��D��=��k^pm��7���{0�;�зB�����	g]�ᓸĮ���NY��YWWSHaK���_Wu�\�:�C}/83����(��gK����S�� �u^j�-����׏����ӟv�� &S���НX�s(Sb���]$bb����\��0��{׵g�GNU�2/t��-̵�pߜ��Vj�hU��!�r��,$]�z�a�U�{u�vv(���8�n�>�՗���b�Z��4�h+f�oFEZ���E*��-�Yt�q�tkl*�x�жb>�v�sou��Y�mK����Aii�Yvm�����ޣ���y�+if�����|���%(R	n�`5$7�gI��tv"�Y]J�.�:���.(+ȩ��;wA<�%Iw�LɰY1��"jsRB�6�63:�O��*m��F�I,Qy�~T</f'��h�<U*'�A��İ�H>����OF�n{V�[�����U�z��0��7Om(蜙�EC5K!��ʃ��ɫ�j<����=�z=���[޸�cB)��Zq�Ӓ-뢉d_��^���{��[o�^�v�5Mo�z�+%�Q"�d�ۢI6����*/U�.�C.'�>������lO��.�����7эf��=Ⱦ������(�r�}���4>O'���T�N�ǕWĪ��.GϽ��Ӕs������	�ߟ��?o!!/�mr��f*�wv;���\ns��n�E\h�.�_����M0���33;좖A��S!]:�N�:">��]��(�m�?^��S�Z�|BD�h�C@���ȃ~�}��=�[�+Ǝ�/L-j�5Hm����ٚ2ؽ^x(�Eh"��]ڂ��x�z���Kw�^2X�ܹ��L3^���`���(xh������jV�9���g7/WrΉz4W�7Z%���0�:h���,`]�ul�J4X���u�����bؖ��~�i��{\5Sj�v�8��V�Y�`�P��aqѺPU蠮m�G܂����I��u�p}��ƴ?P��<�UF�ybФ�B���wy"�k�s=8�2[r\��:��F׌����Ճ�@�d�v����1��-:H��*���沸�|�8,aк��m����3{��Y�q�yں�ڮ��Ƿ����Ԉ��*c�W�.(��=J�:x�*�ѳ0����o�x>8��x����ш��úy���=V���� ˿!��;9BTf;���/W.�5����t���u�^���`�Y`ʗ�B�p�vfZv�<M��_��&���Oh��{|�C���L�x-�,ȴ���x�ڍ4}^5b���&��R�j�:������mu����lC4U)156jkffz��289�..����g��C����U��C�EM�He
7��Dt3k�]f�{�0�������l],x���,�J�Lr-��#X�O*
�8�
ok�bÛ�W�!U��I�*jzM�b-)�	/�q6ڠ
�ïyT��h	�]^4d\9��$"���2���j.N=�7��ř��
lb��g�A�:�z�t'x�� �w�����>k'����,s����Z�ial�fJ�Jީwϲ�۳��BF�^z�1�^���UG��۩S?TR!Ҟ��5"˺C�Y"����(�� ����6������O�;�K5A�_�{L̝��/k�N�!����f��:�3*�N�
�Um��S�-ޒ�L(�.p!�zpy֤7��wk�AcD�_n���m�ov����T���jZrv�rv1j�C-s�q;l��&։�J��Ua�;PT�������٘�	{o_i)���0������stph~�I�V8����ü`�6�n���F{�h��8r�W�[�*6`��X4:�`�����P����x�R�k+ 7�>v��+��Y�S'�������:�V��||>��!��`�(C/�j{3;�m��ۙH{�]����]�ޫ��@al�=�����C�����W�gI�ģm��ꪈ^�n�e}p��S��:����T����1��8Xv@�-UP�jQ��&&E;��<�T;d��Ɗ��D`�Mg_����[5��j:0gZ��|L�ݙ�WOK��Adz�X^Q�Ȩ����>�H����=�b��Y�kB�^��t諠a�J�7�j��s�������MXc��P�H�>8S��Q.a�!:bf��ں˜6�7[�][4�`� z�� mi��1�~�����<�Nk\� ��TX�jc���ۨ�- F���1h�&<�������f�����˸Ƀ"c���U0��85X���i�5�X���b%�%x�|t_��:���m!���t�֎>_7�X���bÇ+��!ŷw��+���>��b��-j�W�u ���-G�K��[4�və0�:��W'���5�;�g�^��3p֊@�٧D�Uذ9��E�w��<��}ƵA�k�Uq����v��t-^`LN|�����R��x�3����ǅX��ӣÆq�(3U���ٝq��L;��f.�#_:�<+}j�v�=l�߷٬V c���D��Q�����,V��=hg_�{�����w8�\+٫ T/�;8=f����������RG���e��].�J�B�uft��N��@~A����2]�ګ�Aޤ�ڕ`�VP��V����Uto⬼�oF�r�~�k:,o�A��Y5�u��/����dux�+�=5� K�P��ȊBE�^�{�9�!h��$��7��׆U�(����d�M�ލ�x�V��3}��WĤ]kj5������E�|rg@�C����T���^��%����i%/���B��sf����<6��<��%f&:�+�?hxo��M�f{{��x����كLk���u�.��˄Mջ�Wd+pK�C�����\O'1Ju�n�s-E͸�g����}�v*w*乨��t�%�B6�;���H�B�j����g�����wlvR��Y=ld��]�x�pPi�bT(�ΫH	����]Ω| �tmѫ+�9��vО�؟<ڃ�ƍ#.�^��;5^��w��t�%�c��)k��H������k�Ռ{J�H�\�É��A�<d�t����Ep�f�8�tM���MX�g׮�oX�����8�r3�5Ό�	�B�*� #������r?-�=*v���yd���!:Y�[�![M����T�.1��h�e�#~
��Zm��#⧡�e+�8؏2{9d���5{��:Ӌ,Y�-RC75d]G.NG11{��k�^q����J=�)�����>���W��o���*+\5"U�h�e
yj�&��c�o�g��^8�!t��k_�9������5n�	�qlx�Q���CB6��b� p� �ޒvw���RԔ'Q��}*cn��lD�� �'k7v�3�rdU�0]+��m`!���6Z�L*+��M�Æ���܇FmR�d)�]*�^UϦ"�2���Š+�Z�z\ܩv�1�%҉�-�]LѨ��YJj|v�����
_n�.�W��x:�p|`6@�k�D�v����1�X���їU�}�|j�^��� l�X0:�()��Jsi{�<�����+&���1ΌH��]|!Ob-Ɖ�S)�U�ݽ�A�4j���jK�a�^��F��}q#0c��A;Jh�oq��G�����?ZS�BG`����.��u,��i�.�ɇ�i���KuT;��+qU������OP�+�>�W/{w�r�2p������Pߞ*âvd࠭Z�/���=�"�c=T|�*F�U��WXxk�������\;I������ݨ��..��}���ʜ\.|d��ضq�o,L?:������ۛN��e2��wO�v��5�����{��'�����Z@:~�X-��[C�p���(��h��:��)���:��a��F�"p*�:����	�|)�M�R����C���=0bq��Q]6�G�Zv_)���KC�.D\P��2F�!Ҙb�Htd2!Y*�	�
]����Sd�a�{�Au9-�xD�����F����,���km`����b�޽u���$��K�y,`�h"Ä�'ﾓ'�S�WwG��n��XN;��/,wW��L��L��l��㜥���6�J��I�?
x������@���gy=dR�x�0A��+ X���L�t}h�LG*̙�2���Z3�
w�[PD f�g��M���;!Q���}��֢�2@�*a?�7*׍Bʾ�SS�*�_TX�w3�7��#�	�Y��0 ����cd|<,`�84:0����� U%�n�F�7����	^4p����pჲ�`�b[褞޸+�r��b�Ǧ�A�{�;�N��hU�����f�X���`� X��ī�)��Aێ�1K�1���"���]>5�L^�4sV ���:%g��%���C�fٗ�L�5�Sl���p �eh�Ŵ���[`P�wv�
��+���	�Evl�8C��p���`��u=�:���fH����}_I��ˬ���>�*Ps�R�CU���L֑��F��My.����Ǎ�P$��2d���F����Z���Q��ʍ�/v�n�5��.�J��VPѢW0�����h�����NrK���Q&�|+�h�!���򫡀b`�S�s�8���Qc&dNm�E��s�R���]0Ps�=�4#۩NLʇc� 81����I�i������C����ϻ�+�KJ����+�Dׄ�čQ�sy�ݮ����aT���� ����5�Y�B�Qy�K�j/1I�Y;:�D��8������p�x=2���������^�EB�h�w����籃*��[" �R��[���q���k%
x�#�\q ���F��"i�F�����ӷ����ot#�3z�Vijڜ�PKgw}h�������G�cS�2B>��˦!J��h��g���(�T�܏ �v-��ù�{���2:�}`���noNef�~�w���J���3S�u(@]�������k���M2�ހ��`��`on�F<��m��4��
j�<���e�ngR7��f�pG֒��6�f��ʳ���˩+���(�4_Gz�*��%9�W�Z�zrV`<��fb(�q��_Tl�h���1fe]�-R�5�5 u����*lڔFw�����jY׺v�Tǩ�vp�w��o�x�ehR��r.����3��}.�Z�*ğ�P���a
�d���\���#6��{W��j��]r���f�TN��
�魡�®��>$v��X��6�'�{�)��[ޏ��7��Z�Z��)6L�2��}��F!����K�e|a���a�^H�(�6
�cm�t����]ض(e�����y1|��NUb�q�
W)X��t��$�x������m!(���vk"�6�b�|�య),F��S��.�&�Z^c�
I�O�7C$uYiBr�n��˖��F;-�ԶN3��J�F��R�p�s@cQT���t0�h�-�YAX�d$K��+v�;+%�U)���ܩJXԻt;�v���@�7penf���g��Gu�he��Wc�,Cr�V���
5�m�5����)��x]�Y�,S��hV���l�ԁ�u�@�su�����r�d�Y"��͹�GNaӕ{̓��2ss�r���k9_)��_tw+HfwVCQ�3W�3���+hªTL%�M�kݖR�bG2���ʊn�F��=yU}^�ʎjD!��PN��Яb�Pa���!Yu��e��D����r�/�C�ԺQ�l:�9�OR9����������3�E��"�۲B��ʟ0���w��>�'��&���g��&eC����b^s&�>�{{n�"�}��p�bU�]<��s�\�<R!���G�d�j+m��"�l�lm�g���&O&Ƿ�υo]�]�a�	�{�޲����a�\Ғ"�S�sI�����v�s�j,%(�W��,ZV*(��ox��{�u��|����#���7�:s^��ꇓ�yr�be��恣�J�z���oh��Ūj��QhѺ��#���NW3�k����X�c5et��-,�L���Llƺ2���v�S]��)T�*p+�����Uɪ���*_
��p�s�G�L�hSG���aC�fr{���tT�aP0�$Ռ��zÿm\��1���K���+��Y� ���������)�P*|�/"�#B�� H�F`�����n�7���~����<=d���\�(�Ѹ)c��J*���z�{�e�9�����>�ʬ���.ۙ!��@ >����"��	�h	J+yU���<�Ɗ{�FEr�Q��pP�.f`ɗU�B���*3V���.k�eu�=H/Vsvb�����9	��&��S��u�:J�,}r�m�ڢ���Ûm=�x�~	F{�98r�����Ӕ�}ҝ�\6N���1u5���$�ޘ�t���0�7�u�1�.�M�d��P�D�0�c��b.z`�R�S;a�:��{b�"��^n�3O�5goʧmOs�D��w� ���@K2�Rip�'\�U޷���te�;N.i��h�˞�H6�efA�om�_�ieKĸ���'�׼M��q
�^|�_�ٷ�+��镾�:�ɹّ%��Y�{��Y�j�M��كX48pe��Po�ߦ^�H���A�^^�x��g�A,��,��vi�%i����)���xt��X���^�aa᲍kZ��.'=��U�@e 3Mz�'ǅȼ�{�,�h{���u�������5�K�PD�k�C��Pm���:+Ƭ�X���ʽ�۠య��d�F��[��9y�J���~�;QŽ�uu&(������xM���Iʕt������8�R�r͓�tq�'��L������w-�B��b��gW��ַ��f�%^�udx�2^�=�Ѯ� �K�G�`���]���M�u<.ݶ*��:�v��Y���R�t��>�9�������xp���AV<���1m��k{�so=�rffw�xW�%iyʓ5�BF��X��V��@-?c�ǜ��k�N�^�+�\i�/
����U��A~[J(�}ڜ�*\e��u�%�N�k��1��!�A�ʎ��hN�3Z3L��R�mB�p��C]�PW��4��(u�a>Z<wUcS���N�J��O��y"����&��@~E�@`��{�&w�7�\��V�\ Uث��u��?��i��Ŀ��r�7M��ɚ}�l�KՀ�s�fg��ߋ���Q�]GF=ۧ�1!�l�U^w&R��&5��۝�������-����	��+�l^��W7��ǯo�S�j�̗�+��\,�`�	�7_��n�''ƠP��6c[�5{J`�g4���
g���*�-8 ��`��-=+G�Y�����q��on�?e;ڵ�>�)���3����ӓ������sC� `�zh�y�@��q�V�/L��x��.���Q��չ�"u���1��Z<w�
�X ��
讼���U�P��!����U��ѣ�����[�){���$5��,(5�~5�B^B)I��dL��F^�.��˱�<4+��tK�p_�ǯ��U�;MM��괻O3.K����L���d�(zW*�S���J��l�����76��Nd�7z-�뾺��� f��`y��Vj���ު;f�R͋B���!���R�����]�-̇c���i.��"����ce����2�Q��P�K��\8:Тk�MPh��➗��A��x!ʑ/:�t��:�s�,)�� ������I��2,�����,��/-���2�ڧ��A�PT8U���1>�F:�0o��n��R�3|ڞ+��
^�݀��ʫhU�|�:����=N�L^~��%r��Of�s
رR��t*1�
�0��.���s�t�x��˭5b��Ģl`�56�2�����3�?1p��ʰf�^(/���Z�������F���{�ڗ\[/�cn����aߕPˡD;x(_��o(z�OI�5�l�]7h9N\�m.�rઅ�)-Z7�=q�e^&�e�i{�M�Ď��.�{9���~����5�:�otG�Y=�F�%��gS�[�z�0'@{5^(�fL�8J���yS��a��g�bb����]9hxE�wUޙ\,}z��r�LI��D�f�X�H�>bɄ�j�P؛�J��kqW�S��k'9��J��� *S"�ɑ�B���*;8t���2�B����oyR��N���<xej�GJꋼ[5�Yi��R���VOI5���Lm3=1��ٴlnQE�
���_m*0���b��h�j�xې����!�YiZ��0V߉ʻ��ih�Bx҇ ���X,L�ڽ�z�֭Lk:(��X�H�Ps<+F�7[mDSY����Q��n�����y�BDv���:ЋuSq֍��<Գv�xS3:���2��!�UcYD
�"i`�>�F���7&P�=TI�|rWN7�����I�F(1���X��vzvѹ�{�@I���Uk��fX�w�\N�5j��B�c��rD�s�UUA�i>�7��.��L����=<)���qV�}�vω�{ax����>5��\�K��^S�V�	W��1��٣��3�aos<��Ơ� =�0��tt]9�ᚍ�L32�R�W=%��R���|+*2���A~U�O*P햴{z���(̙���T�J���4jgg�1Ӣ�����m��k�;ªL*���3Ν�G�H�Nf'����� �"��υJ�{wr�|*����W�$6���c����/��ˈP�ʧx<蠰��օظQC·��S�r�Vl{ٜ���(��]n�Lք86~�z�Q���f�U��뛶wy �n,L��
�k,����bZ3ƫq��`�3�S�ge�����_}�g�Z]H@�l2����"��Y)_���ӛ��W$]�y�N�G�����v��q{Vd6q�'着����z��~�ȸAT��Ӏ;�h�ҥ�E7}��Q��!�[�;1Q�[�:![5�Uj�0i0!<lg��X�w�Ͻ���lAc�/�5��:�k�Et3"�B�(�kQ8��rﷸ�<b�b�� ?Z�v2���4-5<�`���3=r����G�\4W ,?r��W<*����fK^����rP��xW]]��.�����*��z�Tŧ�*0��n��u�UEz��W @� }$��棴�طy�����u�0�T�k�v��;�)0���P��o�/L����`H�����|#�c�׸�5Z@5����3���n�Lw��0Vi��`�:%x����g�ه�VE�T5oc7�}��c�[�kMКq�n��0��[W4��t�&3��{W�\�}!(�K��*�峘��m���M��٣̸Sr~��ﾂm���~�b6]��q��CRA� �W-����o�$���C't�;�f���U���
-<kB�#�]p��O\�Z��WBb�����P �����/��c8�kȻ��.�5�V �Q�P�كLy�*�?-��T~�oW�.�#b���]�,0e
C�Ъ&�(P{)V��3y�����gt�Q;��u\�y�#��`�˘�v�觑��s�Q��Û:���#�=!�])�5�Ԝ�]����Ju��-+­j��>��|4h���N1K���Q�K�������5���J@;�AT���W�DK�]i�Qq�zZb��G�·����U��W*j�=�E��՞�`/�f�*J�k�S�ՎY^�C~q��z�ɼJ��Z��f㇠�y$*���Y�z�X�4U9�J{��ԕӉ"�_z=��˻��w/�Y^![���9GC�7�hm� ڰ��1f��7���T�ì��?1k����0�X�B�X��d��.��c�á�b��5����l(	㢲��~�[O(Ù�����)�aH��\���Pƅ1�SZ��R��8*����T��ё�c��7��6�����[��s9��)��mڦه6��U���Z-�l�QY��M�����n�f�7,@�� �%VA�;X=��]�-K�n)^E��Z�4N�*^;C Ӣ���������ً��W2�p�tL8`ї�]�i���:��r��<'*�ȍU7ͻ�r��������FS���S���#G�$Dޛ����{nt�zkރ�ʄU�@��*�q)��>��0U���v�1wC��[��ݻ�lq�uln���M��q�gj�Y��IB�S�Gރ�xcl�єu>Y���9��
ǝ�a�6&��#���!r;n=g���r��g+l�ϴ�7���s1�k&�9/���ܧ�'6n�$�i{X�"!�:�ė�l���ҧ2�4��]�/=��ķ���us�/��i�n��ò�;�����q�tH�ʝa�,T���^��%����¼����\aqM&�g6�5̙10u�ϊOD�"�!	nʼճqWn��Q5�޻�7��z#I�ٱ�z�r��b��j�Mj���Xӳ&��dl�9�#Ƨ�CBڒ�}lCyDb,4x����r��8sj��m����S�r�k]\���գ)wjz7�m�ũm�T݆�
�[�7n�l��,��j�e�w0�q82��f�*BhJ���P���2� ����3Pf_�b�l*�+Z̅QT���4CZh-�"�G,6�p*6��e�����43�@�-1*1R&��h�E�,�9r�ˣB�]�2FV���_~�ۋ"d�<�.�*W����L,���EL<m8�-R�n�Xn��2���WK*ٹE]cK��%a'׸0^��)�qԼ�4�*�I6��[�G	U��~�u���C�V;��x:���(l�3�WYkj
r���m��u�vƍ��}�Q�eb�$cO-jtH>�'0V,�2�`� �TWM�M��PJZ��PݤH��_D&M�;#��B�G�����V�L��S��zlCy������e�(R,Q���-��ɔr|�;?'�r��K}����d���[J����t�^�2}��P��z�tƳ����M*=����Q[X���f�jaD}lFp�5r�dX鞘Q{�uʏ��'�m������Q��x���=\�}���Q�Ɲ���n^D�og@��#�G׼.��e�<�Q<�§:2g�~��Q^Ȧ���״"<��$W�I��(���ъ�E2h�-��0ȏ��{a�� "�&~t�BUG�H�MQH9]�M����^(�۵\l�\r�ƣ��.ld���+�o�r�_��G�g2�n�.9�����m�D�7Ƭ4tS��C�*��,m����X ��z�j*�Ǚ�Eڱ�ѕ�V:)}�hgM_y���p�Q�\��xog9F��+��d���ʶW_�z�W���:���X'�E���Ek̡Hu�}���Vx�0�����P�w� ���Y���TAA�R��7ۖV"\��� ����^�
�&+}^�_](����U���P�S�U���1LR�� K=���B��d�th�P�9~��_;�X9E��S% +vδxR͹��Խ���л�^���/������b�Q��S7�<wd�V�6�Q�� 1����Hր0;0a<���D�����@9���Ox�<f�in��^:���g,��,Ό��;wzN8��{P��P9u7�,��&�+��
�4��)}��T��g���~�SYfT}�N��g�'W�8t9��\O:O�C�X��
L��	�"4��1J%�G�G���͊�P�ճ4i�S5��#PWvڠ$��u����l�h_s,s8*\V0���5��XI�X��7�lcW6�6���5#��'(�<g+��â�VVwN��H�f� K��|=f��9ժ0�B�1�i��J�6nep�\���u��6����.��W���Y��EP�#��+Ѵ�n��o�`�h+�
(㻾��k&��s���'e*����k3;4���D	��P<4<<��m^s���F��s�\����J�PˠZ��Z
J��vM?���5�Ҁ�6]���j>*f�0n-t9t�b��^J�r�v-n�����'�LQ�m]ے,n�)����5c&���j̴�{���!ݸ�an8����?x�m�\��k�.�ʝ�u\2)����Sꤻ �Um����"�˧1���5�a�rW� �-*f����% �~���]¢0{�X�.��V���:���p u�X\ls�v�<�\�8kA�`�5�Ύ�a@��ѭ��=��S"
`�@WPUҕ3��m9�%GO~�3�V<��!p"�P�5��>���U��"<W�P3>ü��7�ւ=^4||���0hYMXd�TqX�g�=�ج*��P�uo9G1<�}�CJ�T��CF�ք+Fᱮ�b:�����_[Bz v^L	��<��n2�ۗ�mJ����i3�T��E0�.z("54���Ppu�h5+Oq���c�k�|�F�����34����	�X5Dڬ�����+�\�l>���i;�l�k��:C����`��k��-t#��Tm�G��.ܟ��$�S۽~��3�5S'D�\)�Z "�CbߗC��
2;�.�bmƲ�Lk�	[^��MOD�(+3���I5(�z����k�<�1�k�]ں0;�]X�tvk	"�qB�o_Y�3��_�6��������-`��.�fo{�uxSҩ��i��{�Z~������0�i�TK���� f͈�S���[7�ҧ�x�ueuN��'e�p 4��e��s�K]C삛��;,�'��;׷�YV���P@Kڂ^߮��6^���.t��T�=�<,W�r���Q�'hV��)�~�Qh�澬�-���qU��V��V:$X�b�ZO�_Q`�r-z:R=�)���Ұݺ�q�J%|�/L�8� �sד���r�j��H]n�	���9V	E@�ٕ�{t\��E"�Ͼ��6^@�s=_77)2�f:L�Pj�ҿ���s:�c%{�̱~�(�|5+~��Ä�Ӥ�O
6e��GO3!K��Pf0 ��	̨rl������F�W�
@�Ϲ+閘���ᔏ��4��������kUj@�΂NKEn�7�,V�ǶT��6�]r�QQ���/V�v"���9ө�0�1ur���b�0cJ���(co�=�I7�P�t�)�c$�r�鼘�p�a�5��6�K���u�CY��=n����;6���o*��\����碰�ot.�U� K���S��ϲ�Pb����Nq1�o����^���#E�KӃ��
٪���b��6��&�Ԛ��șX�meo
�|#ಉ5;�_om^HFe�u�B���umE�Z�i��R��`s���{{� )����1}k��WޏL�ۨR���n�mF�U�&Y�V�Ǉ3��]\PV�}����Ǩx`]����Mhу������廎B�ڬ� �y�p4yO���C|xv|j�L_X����1�F���j�"�\�_��7Ǒ��$�ଦG���50�''�A�����`
}b��!N�m��l���IDÇ{N�:u�H�g�L��>[JLJ�|}f�kU�(!&ݞ����P�B����]q^<>p��#�Ouf�ޞ@e�y���V,a+�*�<+I�ʊ��;v_-DW8�0�f�y0f�)�S38_4���P���EgotF���9���W<*9U�YP�y�zvV	�p#��G�7G��N���A�*�3�jY������(���K����{��ܘi(1�v�L���O\w��/kw�.�d㺥�*Ϧ^�����ov���,A��h�Ǣǃm�G4�eq_a���e��oag~���A��:��C�N/���Ϋm��
�r��l8���C�)����h	�cf�g+3��K��g���e5#'e-.T�e���U������4��x�c�����5F1ך�.N��({�f茐,e�>;6S����mN�|m�Ţ��a�r?:a�M8?><��ޛ�Ϟ��gB��h���	L�����f.w���J�e����q0�=y�6�Z�Zg��}Z�;M�M����{j)���ۮ������L�hV뇯>�;4 �ꗵƧ-.wd�l�I�����c�!ゃQ����#�_��*~�KH�w3#'��s��_fu�3x^5R%}�����R�T��Ǖ  ү[<�2�r�2���Wn�A�xmhr�.Y��.��ԝd��r+��[ֲ,u���|��\��׮d�(�K��)�>nq��)3=��g�@ϸh��Հ*Y�q��^�|�y��f���`��q� YG��֋f�,64�"�x�w^������R�\���5�KFA�3�p8�����5X���f:9�4�1tmtu{ny���U�ª�g!�N��@������C���#�zP/;��
������F�.�����e��&�@�;�V�YyQ���c��7|��݋������
3��ѳ��i�H��g��?V?b0���w�hws�en��}�a�e��TH�(��h�ޖ�ҳ��m�6�}�li`A���4��3]�A��F�;�躺�!�s���J��4��f������I:����0���ﲢn*[�S >�Kz�vd�Dst��Y�癓���,wG5N�j��|.'<�Z��r��U��.4OrLK��ݚc�F�j2/EuF�ͦ�ڧ��ׇ�P�M�t#x��C��LB�v�����OϤ-��EWA��\*n���r�H�U�RC��cU8ם8ܚ����������"���뀪u��G:�i��+�/AY�M
�v�����S7{V{�g��P��\�����"�U��82�f����xX��J�����V̬�3����4N��3Y�%�pৼu7#�ί+5��I�b����p34��k�p����t\���D�l�v�њ�N��vlX���'�:�i '�^�QVxCݴ��r�(�0�4F'\"�sn���E�d^@�d��/��/�͞�p9����Y�^u7�t�;�~;1q�����mDM�Nj��!�d�.]Ne`�^|��HG��=J��'/8��Ȯ�B�kz�=2M�Lf��ؽ�t�(p�{��;P/�_ǔ\�z:bw'{0s�v�YR���^���Ʋg���� 7S	��<jB�T`f�R�|���j�Q�	��iU�S��CUnW+��Yb�`�C�1ۓm2+i�����ä�f�
f�ү�U�t�i]FԜ�ޛ:�4=<\���)�Iӵ�$�9!9`b�X�t�dY8�-�T�F�A�wNfZ���r�6}�Q�B��}]:�}@���N���EmYt��S�cn��$��5}VJ޴�;�0W�1�b�<!�vn��ˆv����e𐷏hm�`�:b��Q�ϸ�JE�{7U��/6dN�dǉVQ�J��Y7r�;� �a�潽o5*O�ܩ-�g�X~�u�����[mϫ9���]�8x��6��ٻ�S�������yD��.���ɵ���K��]𵮎&�/���I�a�K��<s(����:��tx�G뙕�H��LЂus!x���kspaҵS�0�g�iee��a)�*q�]��kt�1�
��>ʓ
�:��96�{{ 7+К<s��g�s�#V�T���W�]K4#Xe�A;#�P�~�FU��D��at%�d ���8�,P�Y�wP՚��4LwPہ�vr�u�A�n�0����V,�b}V�����k��8m�W�,R�ae]�6���%L�rUe���7.a��T���̰HCw{�����ԋ��/���R����Y**Ӡ�z�.�{D�l����. �5�;K��P��q\��\#r�k���.��ߗU�'2٭T��P3���k�,m�x�����f�.�*�\�ʮ�Ї=�s���P����dp,�^�\����� �U}�����1��%f:�+<�b�ͱ
e���Q*a-j�=�ٟ�-*�klhD�tSp�<տ���\���նr��J�������|]}fHg�"h�a�aYTf��0:�+�G�!�ܺo$�*f�dQ.&ZM�Ȥ��m�j̥���;��N~���(��fDUu���#�v���׶p��/*����:3�Wf��ex��=ٹW��>{{�!;u���������hJ��Y�(f�E�C��>s���h�ER����QQp��Ċr�"�B�ڮ����iHN�L�16l�u�BIQ�����)i���o=w�9ֳ���]'���:�s���C��lNss"<G&ͼ�2E7�2_~����Du����5yF�]G,�;�h�*q������{�=A�u�Y����kR5�3�r���tȂ����ʣ���������жݪAf��A�7V����Y�˗�i�l�،ގ9�n�qس5A�&�yӷ�UZ��M�:�lv-{�/:/�D���R��)�F����:9��ݧ�Ve���S�5�u�2s�1]���m��M݅E8�{|H=�պ�bY�Ƞf��=�Y��\�OM"����P�<������{�h���L���x�n+��z��/�5%_8^E�p�N��˚4tGλ/�C$�f�ݛ
N��.�g'�oyŏ�;	Ԉ�f�[���J����l�*G�l���\�rmRQ�ݗ����:�w��6�al_�ʔGY"�ڄ�:��d5�eiyY�Vn��Si:�u�gndɱ��@�r�Jy�g�k�gZ�T�s&/EC���,��`�:qs-��v��u�*"8�V�M����b9�.�w�X���)�"7�W��Z�q��cB����]ѐU��=�^Fإ�y�V�{��s��O\�n��;ƥ�w��}�.{3�ʴ'NTCw�v��}�Ige5}oik/���Q�ד)\w9��AZ�9�wWo>��*����]�ׅ�5�ԝ`5�"�8j�T�$��D�#�aD���3��Gs,���ں�ϟ����������/
3��MBή&��]Zُt�����(���aK���&+Π�?'��^�Vt2�$�q�\���c��IwJG:��l�HC�%�JZ��x��-qe�ÚT��R�fzs��$�3V�/�3�S�u���H��ϑ��J�ChW�u��ø���51Z�^s��p�f�WV����۩��j%�U�ph�훂k�2r	�q�S���):<��(wڝ��]{�V�+qJWh�W�{۱m.�B0��0e��R78�����8,'�S�;~����]1�b"�ۑ��� s	ٖj�W,k�����_)�Ws`��y$d�+��I���#,f�)TN3xtyG5݃��uk���F�L�,�ٖJ�0Oi"�|�YV�Y�zjb�d�z�7�bM�s��:a@Λ�ۻ����^��q���v,�n��{X
f�NUӎ+��Q�N����\Y��l�}�%���M�>r[тᜭ=���n���qM�����6n+�j��X�v�"d)�����m��|bǟ���Is�9=�T��G�D��=q��$��T�8�M�N��s}���+�5N;��~y^fC�+�.�;�N��}�:�\���QWz.F�GV��f5z��7�eNu�KOw$i���$�~�geh��{^#����b���N�ܒ#X�/��Rni'`u�U��d��|��)�l�l�T�C�i�A��E�p99ث{��9~jn_�#�f>LΧ�8�}[�YS����ֶrq��j'������+~�Cޗ�Ù�o�GT�D
�]�Op���wgT�݋���Gx�X�c�[�x�aJ��ʼ�Q2�gF����}��j#I!����7N�)��ƪ��M͝t���������� l9��hڀ�f�b�BbP=݅զ����<���ٵQVd=r�,50'0T��l���w��rۙ�gJT�*����N�
��Wn���IU�8���rՓ���,(b2H�2^���}�>���H>�G6%]k����{ ��^>8�=�/�+`�U�R��f���������O��k	�g�b�ۧ5v�9���}���̞��eW���sa�e�r4�Nf�f+*�W�Q��ώy���nC^3���ETȡ0E�2��7��"�o�i���xqƼUj��U���Y�~3#��U�V��5z�76�L�w,wF#��Y��x�to{eS�8[ɖ��.��}�4�*o���&V�[����gO< �]�^`X��R�n�#��8�,��&��\����>h��5�-=��T�\I�A[o�*tu��@x��Z2
�tVӒ��u�f�M�T�ynv�Zse�
٬]��V�_A��RP[��9���C�a��2��NbU�[ɑp�NҮ����zklF�6&��MW�_�������`�wg^ej�N^��n���u&cV��Η�D���8[�m@r�D������۽#���!��.�&0�姺�#��͋cOt��ky�\��Mj�+��5{%�ff�3����M�L�y3Zr��ɣ"�{�]E�;��[9�m��r*rˑm\}��U��2J�۽hX.5�1��C1�H���t�����=V�sRKG�c�c�TkW^�qg���փE!Y���w�9��%�^�!(Y�8M�d���Y�ZT���sW�R5Z>g�u�D�Q�
�~�-��4b���R�9pN�-L6�f�MmFvt�B�[=�YPw���	��z��}���S��žv/�[�Ұ��"�=�x�S����B��ڡַ�_f�1�;�==��`��kpU�]�:�eo1i���Z-nt�0&p�]j��,dN��0�<�G(�yFِ]�J�ˆ���^Os���;�wy	)Y�Y��jOU_+kt#���	[r�,D��M�8bj0�MH���0�jd�E�d>�������)i,���d�Z^m,C�T�3�+E5p��3���]�!�ϲ�hK�3Uy/�M��u7�� ��o���dq��Unqb�۰�_�]��w����+�p��¨����[�&��"���a֒{��wܚ��\����mξz�@׻��K�;�s49p��Ubs��mT��.�kW�w��1T�n��Q�fïA�L�32��e�x�u��*k)��.��M�x�vF�iV�������>-m�݋�x&X�� H�#L8�������_��8CR�0�s[�ZoC��DfȵN�1#jII��x����F�⊒��n�r�2KSN5�c���0���F$��Ш�үy�r�{�N�oZ�K痙���m�0li� *#��P�g���MLH�=����x�!ͭ��)Q�r���Z$���g{��G�C�9r��wA��y��=b��o)��|S]��=��~Br>���Zx�B���g9�>-g�hխ����>܊���t���Y�Qk���4ۤ�kTtLogI�d4���A�bm��
������!+��J�V�8�����q��Z�����t�J��7�9w%T��˕(tJ��r��f����p�M]I,��.��'�s�9i�F\�ҩ�:H4��l�f��|5͗��螨���p��aT�j���h�Y�r�cZ錬�Y�`Clŷr��ű�V;�8�Y��ӑ�f��.Z̛��I"b�ޭOM���ف�\��6��̨��9m�\�S�{4W�	{�XZ!S˓ٽZ��IĨK�v+��$b��jC�^C$��U���?	�2S��"X����`�Kg:5�)<�^�V.��B��8���`J�Y�`V��f=0��')Z:;|���zCO����>�H����F��o]h��}�_9��ܝ}��Z���d�����;C8��N�2�}��u�<��o(���>��g�
�sܔ(����z.K�Ihf�R&β�v�*N����$��T�D��̦�O��+��}8V#ɔ+�z$�.e�� �}4%Ո�G�vP��
��y�J���w�-��~P\V���p�9� ����Yl̪�s9W��0��P#2�{�p��r��CT�7��Ͷ�WJ1ڴ_:耢�]I/B��b�����+��D�l9;Jr��`�����у����nfI�u}��XqK'q��wXH������͜�ƝvX��%���Qt���e,ӷ�s6
�Ϲ��k��f�Z�g2�l��նD%V�ݽO�ƕ��ؚ�YhML�qf1����Z���`����N38�j��g���A��Cw:Y�F�.�N��!]!rB�G8~U6�]3C�h7�e�<a�˲R��T/����(��LA��v*!��W�^}"(�RWع9T�'�񰨛ش��W5�y�<y�v�jS��mt��5#7�3ޗc�=#	���}����j5�����v{E<��O��{�n=���i�}�.�A;rI/z�����a�k�B����Sȧ�޻���$����YZ*������,�T\Lz�J�TL�R޽�%�S�4C�\�y�}�����~L����\T;FC�s��I��Pd�顇�E��!U�_�U�Ɂ_P��b4ʈ�ib�*��zU^�(���Dny��,�-Q`��K��Je
1U��8z�xJ�����١���*ֱ�_�w��7jٌ�c�8��,}�gl8o��gw+�ޡ+���-�c�fHd���-T��nܻ�_=�gM���{�J�l��lk"�1�z*le�L5���ów�5nky^�u�����#�z+u�Tf��<+'��(��<!�~�h�C�j�<@f����ȫ�ݷ�SZ��_/95n\?=ve4��
vG�8�q��n�(��������k�O�i�s�dX�b��N��͇��N�;��=��
ٱ��%�ݔ=՟w��=��8셠�){J�b�Z�m��k�Z����x��1b�
FBޯE����k}.�%��K9�EN9K�����u��^,aH:n���ڷ�}��s�j��f<{x���s ��y�{�$TM���ۑ����S�^ �6=^���|f�wM?�C�^;�ʝ,����Rg��jHD����z�]Y/�DL�ɧ�|���ݩ�v�+�B�!#�Λ����.�.2=������e���]n��<�}��>S�Y�Z�{�W{�!}��f���0��d��}�v.5�$��76��G2�Cf+6�q�̄�.�k�WC,�P��}�K2�bxP���qشn'.��;���3�L��͡oo"��=��o#WA����" xƖ�ը����uf��2騣������+a])2��ל���]}n�{x/Uy |�c�eG�.�C��H�q�Ŭ��=�D�V�X�u˖E�rKuis�I�����N��ʒ��Q�v��z�yq�jVɦr�6=�^��U��P�庻�e�t��`z]k�Vw��t*�w7����աż�B�	��B�M�q�ӫ�{���I���f�h�:a�M��RO3,�Y�M�����\�ׇ����%���X�7����P��Mq"�$���^��5�W`��kQ�,�39p��.u���ެ�j��=O9Q����]��� ��B���ثuR�%�3!�zv��	S�2�N��#o7nާH.����V�x�xEҖ �)�-����:ձB㋧H����'i�8�1ݾ�k$�ۚ���K��*�I����*��y�}��W4�]MT�ȣG;/7)����*־~��xd��:�U�'1�:�:k�P���O�}��]@�=<�4��Ѹ��;�爮9/q����c�)�뇬E-��k-�����j�s�%�3*c���6��CcT���-����_
����]�D�{���ey�t>�,�����,=��d�|��b�q���̎Z�������MZ�v+.����Y�'/RE�ټ�7�Kz�%m��ӫ;P#�CX��������"�mv�yC9��&�N�cX�:"�aΉ�I�� �W��r�v�5ob�� �ˠgM �9��M�޿ ��{N��:g�����=B���پ����]^Ooy;��i�oTA=���"v���W��[xz���[�"(ˮ��ꦍ7�f��I���y���)�)-7Wզ��nKv�L����i�W�\a9*��y�8��T5�u��ܝSa���WA���A01�3���;���b���Fh��:ҨEwbfl�Л��vn�CV,�+vZ��y~�GʳO�0Vi�����#�q�:�_�J�@�Y�ΨE��%�Ӟ�;�r�h7�1�.��5��[k�h�ut���=�h��.Q6�Cf8�17���Z)��95���a�
�3���q�!�Ҿ�`�f�al-��#3��F �v�4�U<�՛+ϰ�[�(�k���T��\���5�v;���;Κ�sz�ґ����:*��<սuT��QX�O�ٳ<EU�f��T��Q$h��8�����n��=V^?�S�d�->�,��_d�=g<�沊�{V����Aws�["7*)�9�r	h����99���]1&�ߌ[���4��t���>���#j�4x^L��4pƸ>�=@�h$B� �A�Aʩ�x��w���mS<�g[t�b�mk6�2�(b�7��Nۉ厛+"��8q�\�@�����C�Q>Ω&�)u4��j�B��>�rv+8}<��S�}����8ӅȆo�vĈG!�zU���O'k�EFq�+s��r	.�(^��x)N��`��ǇY��c,�E�/n(ce��m�d���a��Z�{ԞD.�u�nמ��\vP$%xzy�Xކ�:�y��=���(X��F���cC����b��6��zq+�PV��y�Wz/gn���kvC�Ҽ���d.*��г�P\,� ��?
�8PZ)����8Q���mB�v�\���9�m�n�*�4�V���p0o�\�7��q�<-;�;E�ܑ)l-��ݚ����q�q�������s1��������\WV���Z��st�1v.t����N��vOx��#+���ղ�=�[6�_=:$ڹ�/1���xk7�\�5������)V83�2���o��,��c�k��ÔH�'iL�B��^��${���r�ɼ2<��[�
#�e�����Ƭ�߫˂[p���I[{Z�(�x빆�>�K�	���=Ry��gX�8�W
��	U�,,}���#xo�ߏo,�F���U�}�5�ݗ�����}+Vs�_���N��5��Ѷ��KQ±�=�Y(�p:ñ��֬v�MedOH���b���P�zxC6���`�=����+غne5����Ӵ�B������
͚��3Q�kg��S22�B�R�s��s���M�B��	ڧ���:���=S۹�|qs�|�D;d��0���o�����t8J5Z�w	oUJަ���Ü�"�8t�.Aw��S��صns,����{�r�f��MtN�u��F`�hԻ�O���!�A�)��kg�sQeݓ%e�5�-��n�슔�%$����7�C{���An��7zחtS���\g�nu2�~X�w����)2l�uKU��Z�^m�&�D�qI�{w��@	%�*�j��A%�yH({�ar��SP&��t<�R���kS�~�f֣a��
��󡵃317�����`���"���g��y����g5.S�ʮ~Q>�6r�5wW��JRl�w#}L'�ő����eD��#��`mj@�k�tFc�w�MZk�"�ap�����4a�B9E^.�UֲẈ<�Čyr����L[��K�]@z/�q�Y�{Q�( ��zy#���v`S4Ur-Bz���(��N��%��MR�j0d��}�z�:�e
��HT�4SJ���aTB$�{�@�*�zK�
�X�8".��K`�Z��l?Wֿ�s/�6�@$���b�(��
%k����U>2��Z�̬�!��g	XP;��x�h��v6�m?T��`���\-m�"����������kۖ3�.�_\*G��15�K���=�L�W��p�T@��T�7���;?�+�7�o���ܞv$�j�?����Y��q�AP1��?j=]��@����h	n-����FF��'��R�ʵ	�T��n��}�c]y������D2�h�m���I�Ux� -^��PC&+�6(M���Jz<�`�&�!����AP57����DͶ�q]Oy��!���k��4�\�y����zx����R0�o�I��C" *�2�(���5ߊӏhl�P�Y=�l�sGB����zp�_��Ĉ�f���;1�tԇB�=����sAP6<c�c�}F�&8�q�t�EӸ�����Q�AP=���}���LJ�A�$h�y8�	�X|K��(*���DD��ƍ�!3� �Bؑ���7�����{6�����������$�e�kƁ!�*��d�9o;N�ܛ�@T���Ձ#c۰�g�P�M������vi@N}��Ue�����z{�1	�OP��ڔ���`�=䠀�GG;m3��b<d�y�}��G�@��_��?�4�2�I��~:bjs�����K�0!��I=]$�ZG��ϻNAk�"O�tG���cC-�m|�vAP;8�]�����<j]1 ��$�fN����A��T�p��İTY�����@T�|��;���y7��*�p�ڐ
�u��ݵ��+�[
t�Δ�t�AXA�$^�:�ӛ���ܑN$/q��