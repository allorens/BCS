BZh91AY&SY0��s�N߀`q���&� ����bI��                /x
Z6����,���1kY�	5M d
m�Գf���µUkY��A��LIT�)f� �����XK5�,m[T2�wvɵ����l�lj��l��e��YKfCU���2��c�i��Bbֵ�P��fʛ[1�6�k&��jh&f�!
��{���[6�n �;l�M(j�U�J�H�x�T�k�v����6pn��i��.�v�ֵY�f�M�l�-���[5IfTV1�i��=���B���*�Є
@�f����l�l����eܷ����h��Nt�k��,M5ӻi�wm.MY������m��dAˏg.�ⒻA�Хhֵ5��k,� >�P�{�v� ���{ϥZP|Ϟo]�B����OT� ׷+�(u�[�<�kp �=�3jp4 �Ӏ���X�4ӎ�wEQ�}wh�]�H�LƑ5��I*�d<��
�7�}�����׻�N�W���}�=5���z��;��m5F�v��}J�P��x��ĩOA����x7j�ڀ�G�]�)U�ٵN��t�C67��﯃�*�/�:[cem��h5�H��JP;��|R$U����^�TE��﯃�}j�J������|����|�((}�}������6� TS��}�v )@����U>��	��ozo��Kv!��Mm�j46�<��$�;מo�)[/|����44��׻*��>�ԛ'�{TW���=����{�4���]�j���z9�{�
����W{����҆��Y��%e��J7�JR������k��6�ܵ��N�z�=�@�;����� ޼�׽ u��]o7� ��z҇�����1"��,��J
A��  ��pz =�n iC�� �4�q��Fݧ �Y���;kXP ��Zp
��h���j��6�k5@��L��|�JP�  f^�u�l�������( 9�@ë� C���D  v��(�
r���5��4�}R�����E��΀ �v�(�㆚ ܺ޼ (�{x��9�p .;�  s�k{� �竸 �Eڱ�E&�֡!���|�TJ����u� ��Y�
4wN� :sv� �n�����G�:������uw �/�   h      ��4�*@� �ѣ S���MT`      jy2
J��@     S�%*�c@'�  FI���%J�d      !R��J����F��Q�M Sd�$�'����o�k�����W5�1?ʷ����Ǻ���s�>�:;���3�����AU����PE\US�0DAW��?��?��8��@AV��U_��U���%O�D_?������3�3�,�����q�1�;le�^�q��c�c�q�n1�����8�1��cx���1�c�q�bq��8�1�c8�1�����3���1�`�0c�1���3���1���3�c�1��8��c1���0c8�7lc3�8��c1��1��0c�1��M���3�c�3��v��1�8�3�c�64�3��8�63�c7�q�c�1�g�1����g�1�g�q�c��1�c�1��1�gx�c8�3�c��8�1��3��8��c��x�0c8�7m��=1��8�1�c8�7�1�`�c�1�gc�1�g�q�c�1�c�c�q�o�8��c0c8�m��3�8�1�c1�c8���1�c�1��q�gxL��3���0cq��c1���1��<lc���3��1�cq�g�q�`�1�g��q�g�q�c�0`�q�c�1�c�q�q�t�3�cc��c�xc8�3�8��1�c���1��1�cq��g��g�q��x�7m���3��8��`�q�g�1�blg�1�g�1�g�8�1��3�c8�1�1�c�0c�1��8���1���q�c�q��1�g1�g�1��x�8�l�8����ccL�c8�1���1�c��1�1��8�1�c8�1��v���0c���m���������������#��#�'����Q����Q�$\`i�q�1�a\e\a�Fe1�q�q�q�q�q�q�	�GSSS�\`^2.00&2�0�2�2�2�3���A��Q�1�1�1�1���T�A�q�q�q�q�q�1�1�`L`aL`eda`d� 1�1�:aeLd\ddde\i�q�1�q�1�1�q�1�q�q�q�q���A�(� � �c �(�(�*c�GG������|`\d2�0�2�0��)����L������)�)��������tȘʘ�8����0�02�2���ʘʝ2�02.2�2�0.2�0�0'1�1�1�1�<eLeLeL`Laaa1��SC �T���C��D���Q�E��Y�1�1�q�q�1�1�q�1�q������1�q�1�q�q�|l`C��c
�
c �
c
c"� �"q�`ad`GSSC�S�������#��#�����eLae`SSS�SS��T���A�A���x�������c"� ��)�SGS�@1�q�LdS�CSW�D����A��T��q�1�q�1�q�q�1�q�q���Q�D��q�q�q�q�q��#����c
�(�
�� L����c Ȇ0>0��*q�L`�A1�N�e�azaLee\a^�GW@� �1�e�GG �U��G�c"0�2�2�2c ̣���+�������"���1��8���1��3��<x����'��7�`�q��i�d�`�c��q�g�q�g���1�3�c3��1��g�c�<q�q�c�g�g<q�`�1��q�g�3�t�0c8�1����Ɍ�0cv�0c'LLc1��1��|`�q�n��q��`�q�{x�8�Lc8Ɍ��n<g�q�g�q��8����0c8��8����3��8��1�g<g�g�q�:`�1�1�g1���g��c�`�1�1�{x`�0t�3��1�1���3��1����v��:g1�c1��`�Lg1��1�d�g�q�c�&q�1�g�q�g�1��{`�Lg1�gy�<c�g1�d�	ǁ��3��3��1ۏd�c�g1��8�0c&2c����LɌ�l�8�3���c8����3��lc2c63��lɍ�1�`�1��f�g8Ɍ�Ɍ��0c0�8Ǎ��g�`�1�lfc�g�q�Ǐ`�q�g�`Ǐ�Lg�3��!�Mˁ��+=��6��Ms��z�)�P��"*�Q������0릖K!��u���nݢ��t�ZPMJ-<B��ܨ���m�p�[���APJ�i��� [����ԙ�Q(�͍�k�3���MQL��/j�[��4*WJ見�m�+][ܦ��F�V����kfP�:�b��J\�q���$\Ǯ� {b�-�P
S��<�*��*-dJqVaN��m�;ޝ3^����� �u��#bj�LR�У���$:jŽnU�����@2��-F�.;N�є�^,n��M��U+Z���hT�i�ӫș���̤/�4%[m����DY�%kK��	��8��F����њ����>�慛��:�$ٳ��.<V�묰��۳ڵ�	���Y�M�h`@��Ɋ�n�yE�vE�e�2�k76AR���0nE�aZ��44溥��D���<_��qӺ�G���n�F�I��q%�U�r�^oav�QB̛inn$��i���r�B�/&
9l�K�z��,��F��mĂ�5�e�4~F3���qLfn��<�;��d��&P����ڻ'$h��ISn�
�;�v���f4�+��D��X�-ݖ���:�[���r�S��m��]���\�
�˷���-հ�ԣ����Q�o4��-ؽ�9�+�ʳ.T�L�⹡�K/��[���!i�DӳmHU!�$�ҫ.�fP�*Ĕ��kr��Sd7VA��˓1�Z7Ψ˺$\�؀���=�[ZbsSӸ��[�۬k">�[�UĲ�\ŷ�`Q�
�9,��r,�j�f��.V)[�ݸ��F��ws]����
�əY�u2�Wr5�!w�=2��eU!�B�2��-u{v��E6��sC����c}�dn�^*Jř7�:*��cH�9`�;2�54{u���J<b����d�U�1�������q��I��R��9������+��S�?2v]��ak�a�e6��m�3۵��^uP��Q,�e�T���t�xuH�{�e�0nH�Ã
��K:�̚�lh^"�x�KJ��
���-=��TRa�GV;&�l)*��h[�8�������V`Z�R� X����,
�A3Q�ݬ��bKy�`ˬ۱�-7D+�^�*0^���8%h�+��ʃenB����̉ ��D����n��If�0��^CJ��E��1B% qbM��&^S*�h'xr��m�2m^���#&-(��^�T��-��xj���Yي��7x�bf�Б���=ښcFOn�и[YUoa;ۤ�$�+2�����m�'SZWw�q��onD�ym2�fj���`���;&X��)����4i�f�b�*M̚�xRͧ�%	X֜�k�SfSחA*�M����p�k2�7.]Ӽ�qY�GZ�U�ȥJ�V�U�a0�2��. �+.򙳅�˴SK3LCVm�q�(L6�c
�e��fkyZ�J�f=���oJS�o~4�Q�j����l�e�tIH`�K��R�y�{���U��[C^˧j�������a̚�РgB�v��ʵ��5��ie�,��TV��[��wERM`�o�L׆���U3��v���h1��]a���y������tP�ɋ=��A�t%R��Q�*�ձL����Z�C�F^�	eYgei�Vݸ�ᅈ�WA�*٤@�Y��D��	���d�S5T��1�G�fa��2JU��J�@��M4��Y���ұ[�֪܃p)�ї��蒷 d�u�y�K��a�̹.�[K��&ZX(�Gn��`B�y�-�k4�N�6�~5�"�4&҃nK�gv���U-�[RKQ��oaؤ��u��(� �Ʀk`��m���r�*nZ�3,���hSЁ���x�%��#�v�ح�����mX�d�VwlR�u���(c��Ј��.»XS���]�ǚ�e��tE-��?4\w	Ī]�Y���55��UC4]�E)�Ax��i�ó�zI��2��ڍ�1���T��Μ��S��:�������f'����z�ee�N�V�n-�6 q=o��j����K5�27)�,3X�DQ_m�Q�X���Gb,��#ӌ��ҰU���uo-V��:Jxr9��Ӊ��u�,ᱚ�v[z�a�XB���k�G[A\��S��
��a�X6���0�*�e|
�{�͛�+dx>Z4�l������F�-����n��f��\&	�;�fm�ڛn�`�ۅA*�4-�M\VM�A�d��F	��4�oh`h�0=���ygm��f���+D�Q�J�X�$o!�p��V'gJ�b��H�r��1m�����ښ̵#�m=��G���IX��a�ch�Em���X(��!Ù0��(�T���h��+��`l^ռ�/�U��M�5M�	#�Mv#�{E0����0��^KK5��W0���e��l�ڛ��[V�D!r�*z^ޫD�wI�촨CZ�Ӕe�j`�C����S�P�JP�[�Dik��Y!F�z
J�VVTY����M\�.���i�J�f
y$��Yj��2A�����N M�W�n�84Yo	����c�u���̘�0��5L
3��݉b�A�؛
�n�I��=T-J8�MZ܌h�AV4p��;�-���Ц����pml����GB�+1���K3mL$�}tl昞�n1��"�M-��<�M%}ef���]`���7T ܼ���^�;�8�iH��J B��̔�6T���[�h�R�-��Y°Kۙ(2N�V������a8��{�K� ���R��(�f���ɭ��SH�`WP�k!I&]��V��d�3fMV&����/�<�Z䱔��"i.k�'^miݳ��zZyb��X�fbq%���Yu3�G*l����[ s!O��-�{J��yI�6,����$�o�W�r$7n�a����X�i��*���Y��s.�]�`���X�MS=;1��̗�F�� V˳����zl���oE]4�d����ܳ5���Wt�n+��(T��fe�a���z/fbXZ�\�]	h\P���i�"���pݢպ�uHҒ�;��!n\��#d�17x�`������Hn7-Yȍ��T��[Q�&���`�/e,�i�
�+�2�����m��E�Iu5ǔiU�Ӥ�D��l�F;i�	͕X(!�
�`��;&���k%X͂�%�^l����/1�@�1������͸țXeeEBl��Yn�jk[�Ԥ�2Q7��)B�m�ߍ�q�sI�h:��&�X�Yn���l^��V(r���v��԰G����IL��8v<�i���'{,�I�t�6c;LC�
�cx�q�,V�U+�Fm�nLN��9p-b+j���u��.�aƘ�����k}���X&ݼ+IY�-S�T$�2�I[L��8��.
���&�z�Z��sCQV�.;���XջE���	���,��kJ8r���F	B��ɱz�+g"�����"ůvQ	�kv�����3H�[kSi+�\H��Ȉ^�6[�^�%�ey̔p���+]�������J��ΒLw1n�$2�^�2��Z
œ����]��Lʱ��9�l'q��ZɬPY�b��]4�%)���ј����^St�c)�V����p�am��ۚ�&\�R2#N�[Y��`�UZ�t�r�L[�ʹޑ�X���6���*���Y���U(�ї����;�UF{��2��9T۸ݫ�Y�C:�vo���Ђ�R�*H��ZR���.&���2��� E�7���	�Wc�w/2�7�5�\f���w,c%�hd0�P+�@�K��X�/V`\E Շ��q��̺_SZo�H@n�PX)<�.��{�ۭ�D������I�j��m��T}t�+.]�7X�KbA��X!bH��.S�w�ۉ"���[�0�4X�r�6'�f'
Y͘7si�X���]���5a���]	r�������a��wz���l:�Ԡ9W�d�z
a��h����jӱ�w���a���0��ka����4�1Xo�o1I��cI�/T9t���6�����s0���wP܀��ÎV\�r���5c��c�p��/NÃ#��$^�C��ͅ鱴!וd�5�՜�Sl�*�;�=qn����66��j��U��Ǘ��æt���p�.����S�pE�W)�H��9���%h�DB�#/Jv&/&�x���Wgt�#-��\�rYϖK#urʛ�Լ�[�I�6&l�K�G2GH��5�El�����Oi9�sjK��?.�d
13Ftj�ӺM<ڂԠ����n�����J)�p��mIf��I� �w6�`-�7u���"�,���N�锺ú�e7bA.�u���/����y�4��ںO@�V��ue�V�G"�U�R�Z*	mER�aȕ�v�vFi��*I���Gn���.�U˶���ۀ��f�P�-��["�r�t�hB��ٳ[���-J��kN��	K�{�P�sl��)��^�^�ݪO��>�E�`�:�ңP�҄:\�رP{���*��A���-ʘ/鸷/d6�6 ��Je'd��ha��ע;�F�3p��4amPn��ʠww��$��GU	������Ѝ=�%f�XR�.�"ݫ��\Lf�t��3�઀T(K����8��!�ͭv����7@�w*�*�tMͺ�ӗvH�Osh4�S.�KW�U�ڔ�7#�Y/L�YY�%rnѵ)c�S6�	�&�V��,�U�lX~Ujl^�rԎ�1��o&��˧�j�`�H[d-:�L(��ʽ���9B�� ��N��B�>.�0�Ǌ^����u�=�ת�aX���O.�L"��k4�f�&ԲM���H�p		�3H�_�K����s�y�r�%(���8���9n�R��6n�kt�be�Cn�:��r�x~S,��3p�FP�`2�,lU4u�i�# �q�t�W!��oO���VΊ��f;�����C+r:eh���Y��^cV��n�E-e����;���&����� ޯ�orm8�+ʉf�ͤ⎋�of�uWl?9��'w�"
UE�u/LÄ�/�Xq���w��f�'Ol��3E��a�6w�T��ڙ�[m��rKy�E��=�/���	�ZoU����+�2a�t�ǔ/���[�L�����1�N�j��R�H E�E23��EԳORyS�����A������a�f=Q�%r���3C�w��G�b�.�M��ڼ��P�����[y/���q�˸tC� 2��6X�լRW�3ʱ��r�!g,�J�Jv��G�F��e�Eҟ_�_`��jv\jR4��J��%,7֦�7��q�p����7䟻o�o��p���驊�sv䴍:�j=���Bq���Hw��u���`�����D^[�6 ��@�����e��ĸM�&�����n�+"�};u����l��ZEx��vQ`܉BF�J�9�̔%YV�.	�,��o4P�m=�ƛ Q�&�ހ��B���.�H6s[�v���J�4�Y�'5��Igo�B6�&o4�MN�S�lf��\�|��.�fi�D��7WGJ���}m�L�]�����N���n���"M$���X'u<�\ōkK��L;�wQɩw�uomlOP�-6�
�%�;�r����e\�^��� *_8��3$���*�] �ruܗ ԻЯ���V�;1���|��f_NK5��X(�{6�FY��{�7p�31m[��1���֢�\�t�Er�v�yvK��δ��mV^�7NDȥ��k�b����qu���]�$^�F,J�<RM��������2+�&�߾�4��[��F��k���N޹�qr���]օ����̮n��92�����jY����!�]�䜭4ta=���\��a��źt�ͧ����{�X\ew��f�l��m�������<�3Υ�f�	�uf��cK��s��P�N��Ct��JZ��akʻ���r���8��6v��
g8�/&�\xB6���Yh��rc����i]-�Iƺf�z2됑a��>4��%<�0�k�&��u�:����Ue�o��`/X'�Y�M��E��2آ~��eM<��5IB�ǻ�8Mp�:��]��lUԴ�ɋ 1Wj0~�؞ꕊ[8���+j������lF+�P��4E�h:��$u�i�띪�b������hv�̣a�I.�SB5hV�w�S!���M��|J�W�c�]��Q=��yn�;���E���a]X�'*�%��px���H��*��6�V��{CE<x�1a^�b囨��;e�g��k�x'*Ͷ�7��+����T��2
���+��7�d�r-nҊ���������I��Ɯ:�tW�)$��Q��X7��=�n�FKc��޼Ƴ=]�uQ#j�+ś�:�S� Ġo�o�d�;oOkNl�O1�X���!ಭc�EQ�^}�TX�)�L���3k�&bY�ؕl�d�|��V	TH��v�z�te�ʒ���*Z��fձL33nK�h�S1C
zvlP�Q՚�c��!0���Hgb���ǚd����ɹ�[x���?&��kn�!ȍj*�*z�;�v�d �i�wA�;����J}������%!�,o�i�V�}F��7�+X�,��,*�^)�<Z�ŏfR������f�g%��a��n'��䙎�<�L�MB�]=Sթ�w��r\��I�$��N�*�zA(2+qHk-����6\�Q�f��	`�Gn$���t�`G���H[o��ҽ\�X�º�vK�������ܶ&uOI�1j8��4@��̅ۢa�j��3t+s��w�qU���dҶl���@�X�q�3LL#M�x��(_�������}��8�e��1�rjSFG�&�镨���_��o��|}� �D�s�����8������U�i�6���S�e沖�GEU&Xa�/{�cc�7L����y-�/�-O^r�Y2�
�Vqy�g;�YX�t�*�upݖr�v�6��ot%�"�9^���չnkZ���J��:Α�N��P��C���}�w[��k����Co��ù�l���i.�98h�,vT:=ܧo,8�Зm.d�eR�A�W�ȏ�Ӹw��wo+�iѭuNWJ����ɢ��E����Ƚ��I��:��j�0Vk�(jW��8�ݾ�|�7[��d��V�W�.:˱��Ī�;�<�佛7���+�W��Ͱ�e�[4�e
6f�(�)�dIՆ�.0�ax{�l���G�/wJMH%�+��;(K3/��{n�@f���;�GmN�9�m�p����K���F�_�K�$���pf�v�m��f�V�TU}fQ�L���c��1�,
�9�����b݁6�]]<��w*�A�b`�H�o����j��4ﻸ�M۳�Y�{�j�ǛX	�b�
C����;�����M��I%8t�����;��Pm�iij�L�zFl>���_�N�Sΐ�2λ��ݸ�T��;���y)+�N��X���m��}�/��a��i;^q3��:�ڶ����ٙ1��̳����t2��1�6�#�}����Q�w�/q�fn�Z��w}�;�K\�Xv��5����7�]qQK"yZ��<�^�H�F�n
V��o��v-=������z�4�o��,u,���Ի�=횯5�]������=�|�wm�6�o,]n�y�����Ԅ_Z�)�{3rg�#*�E� �4���٫EH�.t�<9Z�W���v9a��Й���l��{�!N�Y7Z�k�祁���n��=���{��.��u;9�Yb)����c�b]����p�שox��ze�]uץ�4�Ύ�:��̆���1}Fs�2����J�ptK�ޤ�f!5S����^!�@[N����OF!7���l�pN1�9���eL�W�-�>}�j�T��ԵY����%ݻb�CH\�&n�hʽ�%���ǆ.��ƞɊ��{o�9�����W=��|Ƌ��V�;�O$4؏t����%.���7]N�l��,pK�[�`>�c3E�^����]-5I��=�����χvL[peft�*�-9Y*:ü��!��F݋���[M���ǰd����V��-�˝��/p4��gs�:�S����=bXX(d4�yr�ʅsl;�J܎3[`�R&3k9�'w2���\�A��[�S�mc��\�(K���Gǰ�����ĵ3��Ѧ�
Ñ���ld�Rl6 X+�* ��^a5ُW�M��_`7�Y��%v�0�D��H��
��	�yfb�����%��l��T��Z�!&���Ɲ�S�[Gh�-�f�.��G��R��V�,R�f�6���Ҩ�ӛT�Lc���b��6�p8��"�iYP���{�3�j�F�c��M��9�j����\r������_.�ùDĚ.L��1+���8�.n�G&�W��3�z�_l�Y�ʇ
�m:䂇����q���r��żk]a���[͗3z�1�i�2��8�(���&���p滖�&�2lczK�"�	�x�C�Ku�n���bk/���$��9I!{���@a�"��o�̷�1��0W!��v5y$�9�w�e�5G�����o�r�rnr}���q}�\²��0�'�J�+��q{q��c��aQ�qT1��w��΀m622v2W+�gj�Q�{�}j�C��[��]nlo�J�ht�[�V�[�v�W���u�º@�"h�V0H-�"�ӽ������ݥ�?�1�7�=��Բ��*�f�ۥ���[oQ��Ȟ�f;�U�>�IXb�}b+�$Q�Ó#�8p��w2���^k����we ����{�v��,ܮ=�������pʊ��B#�S�𝝝�W�F��Ր��O�6M�ژf�n$Cr_]��$�(e�y�i(�o�A˱�9W�W�h˧�qv*ِv_1�b]��X����3H������8Ls���˧|5�ǘ)]�Mi���x��f�U}xq)��g!)���ַ��uVV��3���U�(�Z�+�2�.E�E�ՙ~�3�e�����Zس����}��ٸ;3���P��C�
M�}��L�OnLH����D��p}{�b��&����
��s���#����l�����.���fu\�]2�Hs�T��@ْ�����������K<��9+����*�=��˨�5�fAn�r��,r�τ��l����nb�>��[�"vΰ�`�1�8T�#}kvJ�%e[.�Y��F��*#��yEզ��M���w'4��V�X��Ese��^+C�d�j�)����ڄGd$��7'���w+�t�ܛ���������Г����m�NfTX���c{��]�I����7��u��X�:u�u�۳7�11�b�\9微 Y1��:n�����s6���VdM7�t˴��J�N�V-Uk��o�����N��chr�zVi��ۈ�)oX���n�GP*z�/p�d �#���ڍ�<6�.Ԧ��oN�&m�bQ��!�� ��aʤT�R��4��PX�3���|E`��K�������1v�}�u�[Š�K3��0���3�ƞa���ky���;Hvj*vpr;�(�Zńm3t�J���j��wMn�Gn� W2v]K]ഁ�v��[�u�t;c��Z�nv�7t.�#�ҝx���F!���'��76�e5�l)�3�쥷�:�;=�R��wY�t�z�rJr��N����r��f�8�鲩hr�5�nnX��VS��*fm�,�a	���d�2���ގ�9�=D���uIΒښҼW�&���Cwz�gd
�n[v�Z���Q���U���&��y��_�4����:��]�A�A�*<��D�;9wb씹�k�=����h���<{2>A�̭�0��w��kr]�_u�څ��<�O__����x���X+oێ�6�}�Pv��d�rfnj��@�a�����H��"��/��Ɖ�=�+ ��6��uk-h���7��0�s����gyP+	R����7����=S�-9����E�;�2<��9Ĥ����#w�{Y]�{:Q��� �+�(����y��L��Rzz�A�6�н�v8�d�'U���pD+���AS6k���u9�3t�WX��_)����)g1!����!+��ٸpp!i��S��#<��U�f0�:ħ]YVuy�Q�y��v��iT+:�+;��m��{Ii5z$j��7{�>2E�L�,��ܫ�E܄�9(H�j�b��T�!]*�$��Y�@)�Q`��s_�{N�Y/��X$�K����*��Io���G~7�t���E�D*s��ēT���sy��9JkI�a�Kyn5\��D���8<��Cl���	��,�z���+���D:
�]I�:vs˵1����E8t]��vֺgB�t�!��3��ب𜻭�.A�!�����lt�t!Ιk.J'a��f�Cr�M����ei��9^g\�T��3;Zsz=����3����]I��� � ��Aw(Kׂ�>y2����u9�V�IK�fw.;���aTm�Ww&������d�l"E;E����ɺw0�8�Kګ�����\���b���u��|�k�x��q�W�����u6Yb���\%�z�����N���6b]^e�=�}j��+	�����|7�����pp6�� �Tf��=�گ�ؚln�ɬ)��&�jӳ|���Gm���u:�)�3��'���{-p�폛�(E66!:��{WYS��V^)s�S��ҞPl���=2'�&�n$�g;�]�4f'�"$���ğ����q,�A�1A����MԻ5��K��9$�\ﾮ%�'��3�/J�{QJ�Q�7�ycAYɽVM1�`e�E�v��t�K:�Bc�[�-JaN8�1".��u��N��M�P{�7[��[3Li����t���#�p�C�7�(d��]��%Y���t�5���qҚ����RtWN��n�ٵ��f`�t�^�܅A�wȭ�CWr�Z�N�Xe��V�1k�n�׽�w�o����^sskie�C�F-��9#��m�h�0\ewl���U��һH�wQ��0dO������]*��j��<�Dm���0s[+]}�*:��i�=��}�\�m;P��v{�߲����z��B�qa��yܹ]G����$��JA���YН�mMv�������y�v]�Vv�msŷ���Pyw���h�)�u����큨��7�^�f����v��v�r�{GVo^ki녡S\"���Y��r�n3B!��Р�c�s�&1��cr�e�x�>;Xr�|��1���:��\�����h���vMS�r*97���8�m�c��&pg\������e� s��wB�dp��w�e>m]�fͱ]�^ZL����Zk�!��RI.�X˧O��9�u�u,ih{rT\�ݒ��BQ���4����m��ű��gr�SYHu�)ZM�q���q�����i��Y/{+7!N���@2;��5s��]ǹ����#[�9�ɵwB�T*�,Z:�J�\�8��/�T�0m]�.�&�M�ea�%�}A����Е��*��w�!�~T2Nl���&.�5�r؄J�0�.��Wt�Jb�UvU��g��W���N������u�īRFYn��&��Wt�u�����+�<
�<�0��_X��,X���:P�t�ܨ�+�;ct�����n���; y�J���5yw�]��bs⯘�-�����Y�uȘ����1ų�zj_B{�GJA�j:˟o/q���������`[kF���p����n\�V�'	�[|yZ|J�u5�p�5���,oO�`�����լ�S]B�;aİ`��6êØ��:�ֺ7@�@�'9^�&�{`��+rf���8jR��{k�ջl�yF�f!6F�'��'u�9f�=l^:e�,���<F[��/�LR[q�㽦���X.����:��'L���+�#�sܬ��7:����ą������NMM]\�u�L1k6��'7�f�m`��ُ-�N�����h#��`�{"�}hTiǕ����;H2n�����Q�;�<,��f�')wɢ��;�c�s�k\���:��
uc��uo��`�:q6�yr��fL�щ�\O����r���[���k����\�����Td��OED���yˆ�l�;�`����^����̋�V>��J��az;���ت��>Fpu��	j}V�Ȅ���m�z�7E�I���vD
�B�*�ub��@垢�m[�۽Z�-���&@_������m]��*�N@�e�h��!2!f@_b�3.r�}��,����$��(�A�P�J��xr��2=e��4N�F��)�҅x8YiA>��I�ݨ�A��5��Pdx���>i�.�j�X�\�6��m�ю]x�V�;�sN�D0���$��-ѯ6u@��k�l.�>;W{�d�����bQ"0��h��,�2��_F��,Vr7��n�
$P8o*���PY�4Zt�,�r
A�Z.�- �ldb(�mB��#L�׏��
R�~l�l�`�r�viK��Z�F�Ici�O�J
��9�UJ���<���C懤
RR1.n[{���<V�QĞUmvc�b�ʢ�HH%�^��-��Y�(kxÌ��S�́���N�.[�@�^�8RN�U=BA��7Dd���q7�G^��:v"<�:�^��$�r
/�;5�QS%��K���o~��l�5��p��K�e�d�6[Z���F�W~f'Ezȸ.F�UZ�I���V�"��Uj�6Y��j��*)�m��RQl�	�檗�m�U�� ��,�6�j4G��Jc�~<�4����^��Q�PTHB�B[[�~�:ROl�]Z	�),�Mzc�n�AM�2ܫ][�C�7�Vc4��#*L4b�z<짼�I�\Q\Vcڗ�K��Ї�H2r�&�LM��-��k�h$�qC	�I>Z2uq�pU�ۢ��R�F[�`�#uY�j�]����'[a�ب�Sb�X%!k�5D-��\eY��B ��&���Xg[��J���oP�j�v�#�Q"0��kV��\c�s
��'�F�	7�ۙh�C(����%��sm�Wa�}������	r4�2BDa�*�v���O�,���ޞ�U��[��G�B��(W����#�M:�]^xb&�CZ��n�W�jMI�I �Vm:1HqC"�
A���v,I��{]<)�
N@�e�h��!2!f@f�Pp�(i�Q��h��C	��[�9��,H�,@ˈ�T���>l��$�I�F�4�T�&cn7$ֲ�r�Uְ��H@���������I	 �����������A?��o�~A����/ȟ�?�c���:�߭�5�
Si�r�`5����j��t��P�8{�;��*��qP�#f�w�I��PG�~"���-�/�^)ۧZl^c-��ke�Jҿ�sm�'rJUT� w@�n2CK{�d���ѩ��떎���PR� ����e�+;_Go�u4�2zUw:;�٢����Z�W!�UI��b�1Z@�[��)�}�o�ht�h���2M0wږJ�-�ڣ��󑝊����)u�7,��55���
�]�]8�W�ݶ��A�SR��_ 7Bt�T��E�������+m�I���E��]�V�U�>U%���BUR�x�;w��YOS�����&dlˬ���ú&�ǂj��vKJ
��N<Y}�j�,,��]\&vz�9�>�Rv�<o�-O;�l���|�ه&�X3��v��rm5��U�v�J�-НС6茙gH��e(w^�Y[ު|����ΐ3�8]�ʈ��Y#s١-yڑ��h��7K3!}lS�Y�����E`��x��|1�%�g:�L�z �9Ŷ����Z����ve.��:��ק�������~?]u�]q�]zu�]u��]u׷]uק]u�]q�]x뮺뮿u�u�]u�_���뮺뮿]g^�xκ뮿u�]u�]u��]u�]u��u�]u�uק]u�^�u�]|u�u�]u�]u�u�^�u�]u�G]u�]u�㮼u�]u�������z~�_�o�]~:뎺κ뮺��9w�>-�K�;e`v��gM���T;z��`�7�K��TȊ,@�췦���<<*�ɨ���Ҙ��\�ׯF�v(Hɤ��&WV�����h�q��Ϝ ��i:���ůek�I
3T�i�ˡ���k�� T��3cw[aOS74X�#�w�/ ��z[�D�Bden��T��ٮ���E���d�u�Ҽ��`��ךq_�,��Ỳ'<[����ǥbۄ�%�m��dwd͔!�]�i�r��rf6A����g%����݊�􈵪'��G1��P�,��f�rc�z��E�˗	����tP��r��s�j�F�Ͳ8NFn��-Uq֩�d�i�,�*u��#.�ۛXcKx�Mh��#$�1��xn�1d6���m���4�ؓI�f��7Ҭ�ñ;:�#)��/L��,��nX�K+i�]�fWXq��*,��Rt��`�b�v[Yv�(+w3n�U�p�,�x��Ŵ�'�����1�9V�>�{5�{shN�o�`K̕�f\���:i�}j��6XN�g+PY3�.���@������/�C.ߔZ�G�ی�K��Ā����.��Qx���"<�U������ޞ~���뮺뮺�u�u�]u�uק]u�]|u�]{u�]zu�]u�u�^�u�]u�G]u�]u�]tu�{x뮺뎺κ뮺��G]u�]u�]tu�]u�]u��:뮺�:�N���]u�]u��뮺�㮺�ۮ���뮺뮳��뮾?_�ק����~��뮺�믞^�w�����y
%G�q<��#8��WO���y>��{�T�fcԃK٤+퐛7��n!��Z^Ź���-���L��!����dxmmQ����av@Csi�;kH�υ5<�/ą��9�t�{ q����*���V3�<���s'm����2�����$��FD5H�'P�{��%�O����^�8�L���}?vF.!x�Ϻ�X���97�*�>�Z�PB�ց>�\cio�T��6e/qo����� @dwaM^_�e�ё��d��=V�|/��Ԋ��CMz��$/:�n1�"-��k��d3�  �;91�^T�ᙴ2	���v��֩z]��9��5�QG�1�#��
J�:~+.�H�D-��~�h,�O�17M\_�L��+^5b�:ztY0����f�5�Zӕ�{��Bü�ƅ�C�+Ќ>�c�N�0��-xB<<�-�7���谊!�0G��G[&�'�$�۞��y~�^��4����K�:��zy��A�k�qq��5�^Bn]��z"��r�Ł^h%C� ]-,�}�����z�;��ʬ�1{]���0�T�or�.=��\�ϯ���N�����a��2�[d������:��C޸�,��]��U������Θ�V�7n��CI����GE�/;-
�hI�������oT*I�Q�	Tm��|xJQ�z])b�A�U�lN�M�!�e��:f&�Q��㧢i�۹-�ҵL����ov]�`�}uڕ\���{��Ӝ������>����������]u�]u�]u�_����]u�]q�]zu�]u��]u׷]u�^�u�]|u�^:뮺��]g^3����n���]u�]u�뮼u�]u�_���뮺뮺�뮺뮺�u׎��N�뮺�k��뮸뮽:�u�]u�㣮�뮿\~�^?_�����\u�^�u׎�뮸uo^g;��s��y���Y�`�����)�=��&��"�"���j^Ӎ<�oS=9���W���Ц"@��*<}��%KT�?>ز�)1�^�v�ێ�}�}����i�<p�.�z4�ݲNd��!6k��d� >�����Y(Yہ3��\��Ƙ��
���e�w\}�E&��/s��)N4�=)���n�T9��N,�c�IUcs�{Ֆu3
�X���cxJỬ�`[��>��9���ko��[���lJO:��N�Y�}R�C�s�N\��+o��u��������K�ή/gh���7�ސ-)&,���ELU%)�wؑ'��1bB�9�.��R/�'qwt|g.}��:䢦��h�t$8q��y�Ҟ&1��Sˉ=��Y�wb��ѐH¹^XkK�c�2�g��`me�ٖ�hn����;.D��K��R�uE'�:6
>3��!�rU*�z�.IUW��Ҿ� �^XEYw���詔F��߆�Â�b!�f�u5'G���*>o��I�Wqv�R�\�p��޲ATؓA���*V4���8d���FVN��uZ뾲蒰��X�����@�F�T/׻&����k�۽�[1�)6��c`��,1���,���t� n۾���gv�=���Tٹ�]�c;������Ƿ��׎�뮺�����뮺뮺:뮺뮿u㮺뮺㮺�뮺믎��n�뮽�뮺��κ뎺�Ӯ��n�뮾:뮽:뮺뎺��]u�]u��뮺뮺�뮺�ۮ�믎���뮺���^:뮽:뮺뎎�뮺�~�_����~�]u�_�����Ӯ���������;Ͻ[י���$+)��mE�����5�˻<z�/A����K���s��"��j[���TG7�i{Ui4�[�]|-Р��J�Xh'��2����w�����m�UmҞ `�y��Sc��+'X�]��D��F�3gT�o�nn`u��-�w��c^�<K܁L�{ut�*0�#+���g��Eg�\�5`�Vfw�qf_J,"����nS��,Wi�6mg��'��3�.)l:�`b�bb�q��i�)����kiF5vPe�3�#ȼ��]�M����7v�V�q��o)Ps�O��;c+�[�]2J9h�	"���=������M�sׅ�V�t7�8��gim���r�A�jK�ʧ,�}0OV���ѷ��'r���Gd=3y��sh�;�i�W
���^��1Du����z��s�Yk��b�9 �dݟ��V&�9�V,,
#L��Zx%_t�8\*\Ì��s7�!�7�аl	.�6^�b��O�[��\���mk��d����0tUe�Ct&�:��'Kjv�Ӯ�`��ε���a,B#:{�K^|��Nv��}���>��~�����ۮ��n�뮾:�u�]u�㣮�뮺뎺��뮺뮿u㮺뮺㮺�뮺믎��n��뮺�u׎�뮺뎺�Ӯ��n�뮾:뮽:뮺뎺��]u�]u��뮺뮸뮽::κ뮺뮺î��n�뮾:�u�_������~�]u�]tu�]u��]^ �[r��᭝Is��(g]>v����"YV�m�K)�:�F����nA�P놄�n���)A�u��s\���f�V.�ݭ�S$�s�p�si�7̓`,�㡻BCS����שׁ�Y0(a��E"��:0�.�9�2GT/E$;^md��ν��ԞC��+!��13%a����1�������.v���7e�eέYV�N�s�j�8��J�"P�w|sN`@(�;Cܕ�!��b�|�e�m�ƴ�ǢVc\m��ⱄN���ܪ0�B^���>ڳ�f}5^�;p	6�!��0Η,�k�P�91b\%-����+�gm�t�[����T���g�MG�\��NcOX��'H�mMZ�^9*��S;
&g	X*OM�,�x�(�m�b�֦���(wB�Hff� 8(��fWuU�X��RO]:�j��9���#�]r�}m���i�v0銕�<��q�a�T��ulZ�T�w.�yu�Tl��)�J�;$l#��l;�{#p���l;R��:�i�uۨ��,��Kk�VTPޗ��5��1���cCA�����{y2��;���wVz�=��o����������k㮺�ۮ��Ӯ�뮸뮼u�]u�_���뮺뮺�뮺�:뮽���뮺㮺��κ뮿]g]u�]u�㮼u�]u�\u�^�u�]u��]u��]u��]u�\tu�]u�]~:��G]x뮺뮿u�]u�uק^:�n������~�^?_��]u�㣮�뮽��{�3$,��]M��v��QՏ]��+cZ�}N\�O��{H<$���{xg>����sy�vw�ԅ�#�	��ot�2P/ZO�(�^������Ծ�|y�������ة��+*r ��[�G6����M�"ȻJ�=�Ʌ4�Ga���@s3g&�#Y"���s%S��V�*o M\�n�Xz�uS����,�}I����	(���OЈ�#E�5�]�w��ŧ���ܦ/�D,Z7������\�tԳL;W��5��v����'���nU,8������&�x�0�i	�.��;��~O��1�N�w6�[�o�8ٙ���y�k�g��(�"aM�;�~�:��Q�[U5	)t�"A҄2���-h7�����n�&3e�u_tN�n�c$\�>>�]��"�(y�S#��{��m̼�ۊk%�Œs�k��"��f�[�{|.Jд�:Ws�
΂kT�m�P�l�䪋��+��ʙs;�_�s��/��"w�-��aը�Պ������%�Oi�{{�w
��1�1@�hb:��3��Y<���#gKg�N�U��joF^��RF�Ru;�����H�S�B�eY�aV-��ol�u�[��[�׮X��-̺��v��;p=`ř[�;�Zub�rrظWg�eu�l�Dڊn�d�[ۊ�٬��[q�,���3y6��DuU�
��,r���q���/��۫6��3'U丩�/�		�$�[�M-Ҝ7������\��k8�e���0U�W$Vy��[7'];�'����e��(��ԅ�7��s�o{�۲g.i룘,}����9�q+���:dc%S�̓3Jٜ��w�N��z@9�m=�يTS��Z��Y%'�][`���,$.�[�H4]�<�z�wW����3�����L]�R�E�q�>�k:J1��8IV{+!y�I%u��ӝkB�ly� ��e�|���l��MW%O��M�OW��-�����Z��sw ��*r��F檢��T�����2�1b��-�	�7tK5u���u.�9{3"�E?�+ɩ��Jݷ͑,���ª�O١�Z�"�t.환:�8�-3�G��j�W��"H�|1nir�.�l'���ܜ
�dT��z�֢�����M-��n��h�����fq �dj��Hw4��dŏM���)4uV��Mc�XNe�OF����
7#!��$~M�U�q�K���}mt�A�%k#	�
�ϣ�����t���t/��s�-�}O2�8$�\�E[6�f��NCU�K�b��-�|�����r�.�k��j�2V�цl� �Ŋ��V�ym�+:�Ɖ��f��d�O�����7��sfv�������]�,�O��;���ԣ�Ց��-+;&*v�e[��y[r���*u�)��G��V,z�w^�'rg��͙�e�S;���ԲRn�zh��}Cn��ue�9=�0
�Dx9�++Ir	k���hv3WJ��ACeQਸz͌��no<Nn���n�w#�s�ÎAQ�ol�R���eFލ�)���C�x�Ԫ��"W����ԬPͨݹz�8SH�4���b��5�tG��6��ܶ�`V�3j�v�wG��]������6[TC���쇄F���܇YZ��!����J��c�W�hF�j%�ޤj'��f۪s0J:zLW}}jo:�ָ�eή�Ջ{à��7�[��_:�|0���W���%��?oc��V4�w��Y�	�p��1n���gk�R�_F(c\�%,�mnM㹀�����t3g9Wcn�5m��ZP���vZ��a�2�74�-�]y���uk�5J8�7}sW�vr�nx���I��K�A��
�˳hZ|o,����U�E�v�o$,�9�$0�>���m��X.d�Z�I�c�&@����m`1���S[͂�SF��ml���C[�2��2���Ǎ�R�XP̓y���->�����۪ѽ
��r�r�$eLaf&���e�Z(rA��.G|oT��_fM>�q�a�KTdRk��;���[�.\ۈ_'y�pѰT��e�_K���ԡ#�Jʓ�j��N�hW�ݷ�^i��uh*�
v:^d[_t�9ݓq��p^*�1�.U���o��8�C4��9a=h]`���ce����q����(�;���:�t[�)��8>T��V!;�� Y��,1,��u�8�Yj�N�x�rV�9-��Щ��]�
7V\�4��m[j��qG�����^���)�;�2,�y벇���	ʺ�m�������F����%	mN7ծ�Upe7�g���QF�ŢѪ%eKmK[h���������뙭��?�����@���?ϯ��_����z~��߳����#�����n��� ���r�{$�Vq��EK�5q�D�,��.�##,��
+��lvbAX&��Zm�ja:j��:i�i����v����fe��o�z���
����|n2s�ƹCڞ��v�R�Q��m�rc�Ha���YN���;gU+s*�]�oTg�M%QY��Lcq�h��[О�k�����eU���+�b���v)��į!���C<S�7��̆)y�W��vO���申S)�ÍG�W+�&>��v�-S�6Q7�����9\�&l�e�9:&$�.j��redגsQ�S&i��ZH]o��6�hBsxb=�s�!�2�����>��J���Q@@��;6�{5��x":z�U�;�Ɵ��C;�OvoWU�ʥ,\Q��kۛ��!�#���ݩ��K��� 7�$����K��(d̙e��10�#+��i滁i�{6]��1�`=�Q�aNt��m<BD��y���VA�4�}qN/��C���/�3��BT�tl��*#wm;���L��&[u���ɘڄ�䷁�8Mە��1mvǸ!�{��扛י��\E3�X-�I�+��ټ�n)ÔS;&9;���mN�x�(�I0��d�rP�&Ԩ���	Z'Ӫ��s�X$��MU!B��ZIM&�e�R-�l&�2;+ƚՍAyѢ� i5U~=�u+�)ˁ2�T�A��<�$ֺ�J��Z鄢
S=L�_���6W���㥉�$m8�I~F�A:V�h�[�d�MU��@M�� �0YF�N@�	�R+�8nf��%OY�I�{�Ͱ�z�ɖ�Z³H-�La�Wt�HPs��zx�N8�����ۣ��Y�N����`�V�IP�����ϒ�0a����f�z�~i=K wjm�
ш�ƪ
B1Ur�����$�Hvy2.8�}|{{{{t~>��<}6fz��4{5��Ԕ�T*���!@P����U�Ȧ�
���*�$
�a�1�Bb����@PeVEY@����B*���2���đUTRۖ�Db��lQk$��Z�1TX��UTEXEPP���S�s#779>������'_Y�>�Q#����!"#x{i���X�i�Q>�����
*�X�	T��L�m���P�Q���H�,E��b��P�E%�Wzt�J��K23Ss�ɹ�����9>�F2���Ka��J�jF���%��,*]P��-�RuI�v�^$����x����˭h�4��=3�㏯�ooon�����3Ӧ�?$��!��b����g�a6혆�`��+4�a�1���L����2jY���nnjjjt��O���2}��i�T���J�R�YTIU�͸��Q&�̱C�J�QE�ˈb
;�*�-<2�m&$��b����3*��J�U�оᕘe���a�i2��$��Wb�	R
*��*�
��̥咸ʞya�E ��T\I�
�Iw�&%�J��IZ���¢葒���YYR�PPq����4�����^\�JCq��<����i�� �k���8T���l��6͉)q�Iã���Ѣ��!���LH�t��(]�1ѣ��=BT#\��3Ǯ���ml4��;�y���O!�7ޮN�z�O�T�V�M����y���_K*�{��S�ϒ�/K��F�3 ­F��,���fꈝ@��K<��S���� ���voۡ<���+q�l�n,Z����;í���>&�]������U��o�<�I��U�!�jٖ��5��f6ܫc6��Հ��Tk��k<�>�3jhV^�U��oy���Y�[���*�ҷ="�����c�;pu�Ю�@IgE_�ݶ/x��`���7p�ޝ�Sӏ�<��&�=�r�o�|y�;*+�.d+��Kml�+Z�9V����F+����ޓ|��@T�-��z�iz5+�sjw�%�G]
v�X4$�;���{Yox�y��}���x䣷�U+X����O�]
�v󄾗l6*eR���j駪��L��ӫ��R]�n1s��2K��:�"U���5�O\�3��Т��h��2�3������5����>%s�˧ɪ�HN�xq�k$��rShfv5(�5��f��=�2�+gZ<H� x��#]��f�7����F����{..W�Z_a3�{�%�f��ֹ_��Ս;߽}O�~?H�u���dF���%$��k��S�Mnj;��70pg����ϟ(�kb�����h��YwҲ�r�h�(� �@8�j�}jx�Ƅ)}�b;~8CS�E��s�� <,��ޥ�<=u�<�_˸�o�/Y��ek<k�{�~c���Ie���e�BF��g��g/(rj��U�ǐ�A��Uu�Ϧٮ�L��@R[���>�R�m�)$>xU{YsQ��`(��gW�(?�h�Fo%�ݝ�b[����u�2wOd���zHy�&fW�kq9�����V��O$���	��Bv6US�Z�#�͕M�Ky�R��p��a��^�ޕ��@+o]Kz�U-����g�x�t��w�^�m���{�OP���It=Bp�[�&o�g��_��=�y��a�����U�v�[�L���;�5�M��s�8-�'Jzf�W�d�}8F�) �P�h��O���9DT�y����an��{�ۘShxG�0{����ܮ�`�w��@%�}�s�eWg����N[7`�N�����;���o9��W~��2����Bog��f,G*�f�\n:�T��CD��Q��U��f���Z��1�.�%(�$��ݍ���Ĩ��Ԝ���2�StO�ТEF(���^�Y�,H����<Ga��2��b�����8w`�^�;;����W�=ܭ�=~lc��,���}�<�Q{E�_{�m�i�s�e�}ə��^�=��[��{Mzv��<tc�jd�N;�ڳn�#��C��&=�A�9�WJ&��.Ct�R�1K=�G��u3������1O^q�ĉJ*�(Vn��W�Ï
�)�����Z��t�/5��Z��E�B �,��،+rM��ݥ�
>ajѹ�.N(Y�-;:� 0��<��UmN?O��j�7I��!����S(ց!K�	t�>T6��[9�[�����8��)�i�O��b�#�W���n��U�ꪙ��y����������R��Fr�[�Q6�p���LU��Y׏4oXc���ޓ`J�����J$�Ka&�.���}���[ϝ~R?0�]�w�OJ0�0o_-c�O��dm���,_Őu���ѮψH��ڍ�W��69H��x6Q���+���ۻf��]߱[�-����?v���Pj�������)���M�`NV�R�"%SM[nnƹ���{�S�
1�-q�0�� Dǯv�*Y�J�UEH��V��L�Yi7���Ѝg���V����el=�p�!�]�P��x��R���1z|�o+C!IK۶���6%kݙ��.��Ԗ��͔��5�S [~������{��uE��YF��(��zS�Jwc�)n�{dY�Y�65;@B#��uyS굺�]���$"A���Dy4y��lt���M���:�@�}��Bw�z�����;�rۓ��d#�>9v-=!Oj��S��l6�:������}�V�??k��K����Y�PY]����������J���
Zw��.��a]���U�N��{RN�;�^�f����u�0��.�������VX�I������r���u�N��_p׹������y�7�n���S�}�֓dv��߆mbKj�DuL�\*2Ֆ	E ԉ��`ҷS��%��N2��+�2Mk%�����ALH�"~���,�?VӜ|��C�TcfS���T7��o�l�W�}3X�ư�c5�O�)�����E��+vaⅦ���تNa��uCYX���#���Ew�ʖU����m���.���#!�����+� ��-��V�z�۫O������{�����st�������^��A�ٯr�-��M�v��`��t��׽�ǭ6�O�ʝ���S�TYk�0��'?U�m��^�T�6d��K�L�t��a�t������#~���\�=}�v����}~�B�v�H��Wi7���oP5���O�~bM�D;�ܠ��{~FR�T#������@���hm'L�#b�V�����j�h�ф7�0 �!]`�X�T2Qǩݻ�L�ȝ����Xݐ���OzD�2��a����^h�����7.�א� �e�)ꖏ(�c"PJ�ĜB��$[2��Qҳw�����w[�-K�V�����;�'�� %�{.���=L�tc�td���6{'fr��x[��6]���ɂtύ��ו�:�7y�v�Uw&�*��� <��I�@���m��mf�Ϥ\���7ڙNc��� ��3EL)X�6�2�M>鐤�I�$ϯy�ʞ}Ͻ(�y^��cgN�=w$����wSdh��#.-Cܦ�W��ci{�E{a�LwW�j.�v��n�`�8�|C`F��Ɛ:�~Ku^E�=)�6}kR�mB�����H�U��L:��tM?o��t��F������/�.g����&Ȫp��e5�[A� Ad���N{#]�v�x��X�N�;�<u��I;�3^���^�n�/��{�QX>ϲ��o��5ڞ����0(����!�<3�Ы5�y����}6_j��u[$^��[},;��.��	ؘvR�W9FsRF�Q�`�ԋ�N+�"�Y�P��1�
�g�;���s��tN��}�~����oh��bhy�]kz��ы����z<Տ�,̟Nu;3�5|��h(��,&b�K����T�ݣ�LJ�vU�WQ�
	Ԏ�D�bӠ��q(I)"0�[=6�u:��lS(c��ެ9r+򴹮�J������	�l^��8�!�9�(�=�Q��H�n�����W��U�f��F}ίL������go�3��zIǫ���Q�����M�sV��q�Q蝆��9(ѳa-0��I��eB{ݖ�a�:�f5K`�2��ZB�>PΩP{"�n���LZ��A`h�{�\��p0���'a^�\SO��W�	��
&2Y4��m.��H �/�n�Q�B0�!V��򽅗�'�@O�iS�ݷ�����ŉ-wa'%5 ���h�ر��q�7���Z�$GNE�x/{ڧo^����iҌV�S�_+��:>�}q���y�н���9{��Wր�C��9����P/	]��ӹ½����9���$����d5�_x?�9�9n�r����d�H�
��	헍q�U�A��Z"j�n@>�j��\�jТ�)���pZv�D��b�Kl�,h�01+>7�kk�0�U�s�/�SM�J��hM)�[~���K� *\)��ǟ\ޮ���n���R��eNuc �̺!ӟ>y�V*�|�>�i��o�J	k�p˶G0�'َ`�l݁�@�B%>�ի{��>�,1)8��`VIup1C�?�fP�qP����i�K5F6��a0�K�X�*C�٭���{�>�T��`�-����p';���{W������ _ǤsaX�X���V��o��=#�y�v`�����Z2��H�hB�fG��Q�ץ�|e�����"�Q;ibD��e�FJ�ZM�+��b�ZM����� �,���:��C�_LZ��>����o��u�晹�*�8S:�c�ބ�w�S�	�L�<��+e�W�7cyvw��n�"�y���]�z����9B�}����T�Ϗ?�cX�ܽ<�oo��^�."��۞���{���-|6�w�'��Z�ψ���� �\�|���xN�6���f%W5U_}�/n�������&�IڨZ�v��;- Ѱ��iޢ)�ݗ�f�Q�|�J]�:
M�� */.�K;f�e
�O�v��I��d�$Y�$�s�d"�/h���H��G;b�e�РT[ӧgC���}����oo��d52͡�u졒���&q��Q{o����GB0��v�_���NC�٨j�O�(�(�6�r�����u���=�7��vs�&�#F�'_cP����3J�����V
��4�,ha��j1��N,��)��ov �W뵲g=�lk
���� �)�F�WP����������1���ܛ�oӪ�
پ�t�����T�Ws�GǶ�tHƄ_���_`;��Փ�Z��TN��Ϳ���~�q{�))/^H���Z�0�ʑR�e���!�U�@�U~�Г�1$�N��Qj���^4��U��Uו�l��#��M�\|�!��p����<N���9f������V=�k�SפCb\�'��ww�Խ����7��g�z�����t�Yؠ��@���9��ǞjC1�zJd�L�(����r�zB���<��*��5��k(��;xE|��w����2����yr����A'�cy�
{Ӹ�y�\�{�͢�'�KY�:ތ�{y�hI�g:����Mن�C�6�,AT��V+z�/*�;�i��3L<f�;��Fb.�ho����\�W^�7[K�}wZ�}�2��n		?_BZȱY�hS�{%(.����	=D{*��Ԫ�����ßB����{=�z����vn��a��*a�9��]t?ږ:t י`�;���U^ߋ�o���k1��$�W�Jt�4����<<5`@��-�Ns�}u0;�m**0�,�����-?�f�g�b��w/m������6a�e��za��
d����ޖj%^���uX�f9$�nϡf��d�[�eF�|��C!�OK+-]f�����b��~����o���ʟz�9�Ω�k<��W�{>�$��vY]^%� �b���i�gtߥ�s]��;����e�=ڵ�����l��qQ}��~�N��ژ��>�tgf)�`��J�|�P�[o���W��z��F�ٓGqǽ�>���\�N����$�ܼ$�a���Ż4�^;�vJ�����~�������Bf�;�+��6HvʳR���׺#�Sx��Tu�e��`�vl/aC%���w�X��v������do�q��I�l�4�-ؠ���{�r�d���������M�FWSY��WX�甦З�#�p��f�5˸�5��X��-
bs;��i;[w}*������[��Q�;pv������ޝǺYܝ}�+�&5^^PNf�R���v�tݑ©J�-��&NJU���}��wv)a�!��h���l��6S�	hu��.���[�an��C��W�lX<��m�$��ې�>M����������Qb��{��V��8��*���Zӣ�q�����F�7t�WUSL0P:bu���bB��dZ9�D^�3N��n���nbY�9KN:�(�r)��Ԓ�#�&�;u���m>0��I7�9P��z�np��ۯK���C-����9��v�wg)��aS+��͘R[b��ۚlr�uS2��4n�Nh���.�0o;M��EG5��9\o��Vބ���������N;K6�P��l
��'T�[�]��ְ�h�{3������!���g�+�&I��(�GjR7{���v��L5�Q�pX.�e*q��W>zdnZ�ky�Խ���Sܒ����:F �`��6�)�nd���T6����+x"uQ�[6
�DTE��{��J�>��U),��TL[ט2=&[Ԗs�9�
�����&\h��3��/�;��������L�Vك�/y�v���k�\cq-��.�C\��]/,<8�@wi�*�ݗ����j���pȔ���/kw*d9&c�W;������l�N��SbJTCu`Gw��!��M=4�	��]gp�6��:�a��P�^�}Í�ں�#O;L�q��Lwnc�v���Hvn"�d����ٝͷ�\�wm��u[%���"�ܣ�X12"���n���P�ܔ�t�г;W<���i�.��;�өb�Y��9�z�Ӆ����6%���y��]y�A��/���;[-t�3]K1'�H޹�`�YSMqO�A2�m�`�mS��9�8�&&{=�AC$��դ<(v�΃w�to^��W��tEW}�V!����}۩:p�kɞ-Ʒ6��q�5��b����bW֮��gv��|��Pʑ ��Tgwa���u��ut��]I%Q9Ґ���*�6�f��ds
�L߸U���=�vvG�.<�Yٯ-�W8�1A�Y��T����+hv:J2���,j[5=,ۚ�b<�������)�=�4"�=u�WL�5Em����L~Me!R���B�=��55,�r{77555='ӳ�g�̞o��沥��ar��
���f��ѭ�b���LH�wB��,P�gfL��vy>������'ӳ�c>�>>�3>����+"�eE
�FҠ����S��DHr��"�{����ɓr�''�ssSSS�};>�2�w�,���Me�
�PR�eE"��C�ys"ȵX*ŬѴ��1`,>�g����?_���ooo����g�ӟw�� وZ�Om��
ʑˌ�V
Er�Y+;B�<��[���z����ǧ}q�����>����<��z���V�PUdY5�(
���Yr��@�&8�;2dԳ�s��������>��^3��4��_:�TW\��T�Q1+�1���c��-B�֌D*VV��0��+��EŶ��U-
�l}������!Yߖ�Xm�R������hm6��l�f-�T�QJƍPZ�@X��C1gSEAEKb�.�m1+#e%J¦v���¡X���P�b*vԝ��>>��{����o59��5,9�i�8B_d�'��Ӛf��;�m�:�����כ�E��z�)�,��$bF$bF}���n�zp n�N7�|��~��v�wε{H�d�q���G��i�~��|Q dq�7�-z��0b��·�ޖ���9w�@�Q䷂/���c8����"�#QR�����@�dy��cl�
L��B�]$]zG����{y�y0��#����)d�E��fj�X�*Ď�a>%�<��@��}/�
���z�|��r�>^�k���~���~_y �.�g9wY~~N�v��S5���� ��Y ���Z�υ����st�|��C�?������~m�����?�z�x'��p�]n_l���r��8e8t�
�(�W?���� [3�\X��~OL�a�=G��!��a�o��m��E5������ޖ�s>�w��+�nsB`*��@��M'�s۷�z�؁�> 8�Öѐ�3)k�xxfF���;�d>�k�Og��	��G�T �����U^�u͟ �K�P��*m�:rU�<� l�uv@�>�HR�@//���0�<h3>�ۅ3x������*n�VzP�xxw<�Yݵ��<*�����4�>��ǟ���CY~�u����}͟3���������J�B	>�q��YL<�V�.��?q�yx�����δ2�a1a�J}���;����Y����e�Pң�?������/>�큷G.����1��`��
��%[��(�<��)HY˹Ҭ�]d���a�0�3���y�����~�=�驌���<?dh
@4�v��M��3��;7�9���q|<ѻ\Apb'�[�C�If|�u���I�}lz\Cz�攘��ݰ��s�hv�d@CLn�n�Q��;U�Y��<W��*&�I�(����s�p,�0y�&��:�=��N��{|�W�˘��	����������y��3�>`3� ��K�x0��׫�K�f'�F6�/�!�zB��I���#A0ຶ��\��o�8p�IG����j�����}t��ݑ���o\�N�H7�`	%�*�O�,��ދp2�r��w���o8`m��C���g��̻g]N��?h߯6��%���P�����݋������J�F�Z� �N�@�k��1,>��� ��>�?<>	�;��;��D�mS�v)V��Co�� p�p&�K�����3-C�~`hjj�Px�����G�D&n�W%#�z��80)(z���p(�y��sH \�A>o*�Bf�yf𭇯=�	�{��GxӨ�T��l�J�O�v�d0B����Vy��p(�3����ȁ"�x��2db���4e�츘Z��q��b�y�qc�/A�<�N�9Q�;J�p�"�u�M���nq:���R;Wsr���WJ�ˇ˅���/���?��u��K�W0�1�W�,�J7$d��g@�7��&�\$���(:�[�����B�/����)�櫭�k��kmkn2�b���kMtn�	����ϩ,��$>Hy �աv���}��x�duJH�!���v��w9Ckм|���q�QL��Mכ���W'�>��o	�]b&%Te��<y�r/�� 1��Y�A���Y�l>W�0<ѯ=@�@�;[�~��V~C<@��I�:�y�c�lm�l��sn7��~=�Z�<���U5;���c��{���i����	KO;CA����s��1�vv�.�OhF��5b�"���O�	�6� �3��d3`�`����j\�y��C��!�ɽg��.��~CZy�j6�Q��2������2��|-�H������7P�>(�ޞ��o	~s�g G�8�͟A�-�3 ` ��|���#��ɗ��.@ѭ��K#�'��6z15�Y�S������L�~=���Éw4~F*f6O^>�@i~�s��kmK�c��;�«j И�ϩ�es#���p% ih?��55�|}��4L=�R��@�Ȉiǉt��Ȇ@�{����z����E��_i�!`�4����p0��7R�G_�ONX�����������?��3�Z_d.)�_�lͦ��'L?8@6˫�#N9u^�<��9�R��}����Ѳ�륶+�g�x�� u�7��K�ް�b}�ȊoG��3R�g"@��'��	<K҉̝�ݣ��ll��ե�U�Fo<m�Ȩ��Ӏ!~���}�G�
��
��o]��1�.x����T%vis�k�#�Ce�{���`}0*y���Lz3�vZ��"����Q����Y�FR1&YHę��5���$�n�b������c`tF�#���ޟ'�YR�=���7�^�9M��q�MT��T���`��@C 9��;�q���ց����~����荜u��6����s9䋘R�ų]odiO����1���?o��7��冧��4s��ٔ?8!�4��i�#a�v��>g�W��u>�X0���3�f�M9��P=��V} ��l~�ǳ�9�#�M�����Bڼ��q_Z�=�v���nQ��U�%ez��}�ӱp�O�Q��}^�q�S0l	NHE��AD��k\����Vt����}�"�d���G��;� ��7䨁f��sxq��#^L���U�}Y�ҩU�>)ͻ�s�`�3Ӭ=�x��u�Hiȥ��@}�訣��N�E7��S�O��S���沴E�*��z��b/;F���Gīa\��a�q���G�̤��(v0���l O0�Aj Mб]����8t�̫|ٹ>.���s�����/�e��M�>>���a!7��`'҈z��kZ��i��	��s \Ya��#��o?f�>>\%�q�cl���	����w}��!����<w�ޯs����#�i���y�M�b��9�k_p��F�`-=Rhw���M����f�>��h�G��v���<�	��e0It����F@�u΋�<�`�.�<�:���	��<��tp����e.���j���Sk4m0�a/v�KP����HC=����)��Il���=�=ߗ���j���4|ǃ�����>�1����8VT�ǫ#�}- Wl#����ݬ�;���9ѳSw�1ڲGz�&y���V?�7s��l:;<�ME4}�Ϯ�T5���g���ω����̆�тzf�\����ؐ[�Ù�ί8�#���M^`��N���N�Ž��@��#��Q�{/�e�	;�&������}CS ��^�;��A�8��'B�@���sD}P��� 3�(���2"i�ԟ�k�����1����$�Ő;ڢU��Vx�Ͳ@�r��:��K�>�unW@��Sq]�;�G��~4[^�� F�w�D���cՖo�m���_�a^X��0~����KT]�`����u;{=q���aho{����`�4�/�8��Q޾�#�W 9@q���Fޛ�m���r�dw�����ϲ)ޞ�����h{�7[���O���&��M�F��NP=M�ϗ,V�D���2ށӄ[����@%�e� z�(I�����P�;�U���?1*�e��AcCy]�?q3��H���І9=R¹����@�t��At��
B�$_���ٜ�6tFz�ϧ�+K����3�FzfXq��f����Hc�Ʀ#�ۣ)��y�^��s��%�;�&����O}��V���G�f ��}�N%��VҦʯ����{�.|�z��c�Kx�R��O#�23%�i*�w9-��f��ꙹ��>	Ëmlݩ`'���<��Ʉ��5��߽����/�����}�|l�$�vE��R�'|�x��=����o�[zʃ�왷�ҍ��U	�E��\Q���)���_Dz���`�v;�I�"��y݂w:CY�96g$hsX6]q����D�!��xa�������{#o"LܾށQ8`O_�XͰ�O)��ΐ�ӡ�-�ˌ<�]�r�k�Ñ���y�0�Q����&�܆f�O2<cҔ1����v��ˏ�s}[[�9��	9,��Y�jz\ĥ�A�>��l�&Z�7�� ��Y$����I�ݏ.|�.�_1�R���k��d �k�4��EGh-}+����\@7�l�ݬh��Mj�#l=D]��ζ�t��Kt���q�H��������G�zk�uӌ�f������ s�$�	��E_Lw ⾃�x ]z�	a˞}m7�1
< f:�s���bm��USFOE��^6Ĳ���Q����韋y�Vh����s����ȟ�t	�|�R0˵#gz�JD�L��ܴ8M�ÞzQ�g�6L��g���l�]e���v
1_��=lB�{�����
�K8sm�C�ߡ�E�N��Z���*:��u�:��H��)YȒ��}Y��DA��7�2�ߐ,|��	������M�{�/ֻ%k�yW_SyKhufz�\�w|'pۜd|哺-���A�O.��NK�>V*�pS�h�ʡS�6�LI��Q6�a�M�+��#ā����-�ʇ�����,M&A	�E#:�Qu�5C�8��J/��y�t��s�u>�D<=��[�|ؾ;�g���V7{ȷ���a��M�����v)�J�X󍇗h�4�5��s�VZ�dY�j��-J�P82�O�� �g���cb���X.D�B�R����aC�X$��m�en�9硝�^b�;�����~�D���~*��Ǟ��B!���û]�^�*^�L�ǽн��P7�j��a��s�j>�C<pSq>�C���nn�J�,9K�1�c�ֳ�����a��r�E[�ݒ�m�=�0���vF;�*�E�n6�[N��w���l�@>��g{�M!]܉*���l��`i�d���f]P$��#|�{��#��F�VVv�MW�=2���&y�kAZ֓���]��Bz�|��bi��,p=��s�-2�[;���T��M���f���+�4%Dzp���٭R˛���������w����K0��RI^u�����i�����8Ǔ]��6�uH�mL69�^�ý��C�: a�����DD7��8#'���_g�����2C�����q-�R�-u�^oN)v��MVm�5��O��D������3�Z�:�Ծ�%^G���fɯօ�Q�&����+C��y�];=$��][;#��[��s�k�#��#��@���������w�0���5P��_��|�]�� M:�l�^7N�}����K�nC[��E�����ħ��3�fzQoR�G�{�_��CA֛�o7�s���
�D�r�ZTq�qs^[�=ʤj�W�b(��A�IdpM�8�D8k5�w��E����͋ͪ��=��׌96^��1̢�%"������|�$xϣ���̈́e(捔��\����d�2�u�c�330���a�Zi@�H,}S�,Ė��s��J`��ǝp�%k�����<U�a�^�,�/k~_G�H���Υ���xp{�V��dٰ��6a{��u�(�ei�%�p�J�$1��"c�\�d>�@&�vs�A||u�I��c������x���S;�ٕ��py���:�܋x������)�a��:$|a9����&�9�z͹n�,D6_9M����;�| �o���0O�y�іj8�F�X�i�A��j�Q�.9�$�Sз���Heun��%��º!y6�1V�ouT��Z�wm�ސ�Sbh���� ����X�	����e��r�)�}��*I�&��ڍu-��LqQUÈ���%l�S�Wl��G)憷3����C��P���h���rG$��,���e9�Jpe(�rH�6�J���&z��MZ^�����:�k�U	�W�x���y�0�C����<8?p��D2�4���7�Rw8���z��Q����jݺ�k�G�>*�mpL��Bkin�:;��� Aq4�=���ε�kb�A���+VD�~��r��D<��C�v.�i�+[L9mh�&i0��(0�����@�r+�k�:�N���O>��sG��{�ciɎvy0_n��*v{��Ԃ���l�}r_[
�=�om�Q�k���#��j�瞝J'7yRrxsL�ǆ�ws�6��������#���1s�k�gp_���}6�S����G��[Z�9`�DlK�MǏ�ڇC�Z5�;z�wr.j�F��Ʒ<%ϥ���Ն~nֻ��K:X�{ܟ���
{�1T����aHK��8�᭯ͮ6J~[ʨ�{�=���x���{;$�c��m��K��ªZ����3���I�ѓ�F�1,-���C@����ι�9���Mpv��H�!��a�կd��p��|���>?WD'�7p�_�}���Ȏ]��R��`�,L��d0�`G#�_-��]ϮS�a`��$B�<f�Q�׽I�ʹS[F���ye�m��W��E�dؙc2��9ջD1���'K�w��$��A����A����@��a�g�k��ra|�%�]�jus�Ԛ��"�
�op{��gRt�Dģ�ړ��[2�#�f�!��^C+%�����~�����!��0q��퉟CT�"�X���T�,�<�'���|�s��߱v�-�v�9��k��� w����';�c� �k��R��%��X< =��jq&��g��ȗ�7n�S��dO�5�z&�9�嫻AͶ-UH���@�> <D���Ò_��g�F�c�2��g}D5T>b������+�f�v��f�������j$_2�c�%���q�����j ��\�J�w�������ڡ��ŕ��l�k�83J\��Jr��ck _�)���x�z��߹��lk�9� �i�����=�JaL�l����mk�މ�:(٧��{��Mo�ͅ��Ʈdc۴�EC{����2{&]a�j"����I�$���!�`5lA�ɸ��K�@әl��JLA����s�vq�=�E��n���=�^rh,���a����<=��Pq?�M(�R�E{�\���h`���tt݌���o�s��2�S������^���5E>��Om�����69���X;qͻ��TSCT	R�b{g���4�LK�1	���������Vu��~K�Hah$>X������*�v:�ڦk�=��aR��j�5����/]T.$[RM�����Uk����&�=P*UrOAf�Ѳ̴�ܷ�V���V������0�sf]�'�;���"����
ew�H��r�l���bI&u�ʔV�@Bu���p�li�u�x��0kU(�vd��w�/�	�44��z�ߗT.�&��X�e���K%��[(%�e+��/-�c���ac��JṈ����K�B��9$�I.�z�x�/j�ml`Ջw���\3� w:��L�YSo��{ �H�,�v!lN���^V3�[ӷ�j����h�//�ի.��
�{��n�_PD������5&:�Жv���������ak^�:嗡��6�w�^�ys[�w1w-��]b>W�VA�4�"y�{�ŕI����o�z�V]�s)�	%�øe�/s5�bw�B2w]Nw}Qû����']��x�x,WVl˾���Yb��)V��+GX�g8&���O]�CI�ts��q��a���zt��b5Ra�2�5��W�!G���-#tP�॓f���V��g��٥HF�d��aE.o8+;�X��9�XoD�%�8Dz����ٓ��`��\-�3�n��Y������U������@�7�pyt1.�^�ty����ɖ�b��b�3n��Â$yFp��wW!�(�����E���OEte����G�ßc��j��ATB:`�&Q����W �D������8?�!�-���9B��t!?(QH��(��p�S���ݺ�va[G���d�1�����۽BU���0�R���7!7�՘�蝍t��=�n��x��J�겧a&ɫ�Lwڲ�J�.�&&T�d�p�L���^�k�s.���@�-�_K�wlr��(p�b��U��+�k4��`�L5��-M���ǔlp��f������mg;�;:
�����W��u�"U��u�wuK�mXg�ŵ��ʎ��D��]Y}��:��1��jQc��Ec�V�4�V�j�"���pBe�m{s0�aEJ�qb�h^���x�1/{T_kM��6mj YC��
"{ٍ)��8����֯v�h��*6�7���MJry
Ds\&�W/	(ڙ�;;��Pg[�{W�k|jɝ��E��ݪ�{i�O�	oc��Zf���p/3T�v���ϝ'��:�jn��	�q�ڪn
�}��Eߴ�r=�^���'0�WmZ�ΓV�h\Npֺکj[y0�Z2�nܖgwgs���ܲ�f&�2w$����n �
Sz�`WXqt��N��A�-�0V�G�fW>�ir�1nei=G��:����|���Ѿ�r,����[G�_u���י-"�i�d���H�����USDD]k�y`O��#D��D��G�$����5N���e�HjM*0��a�ҒGi��Kr*mRt�Td8`�SLO+RC6ŕB��(�	�#-�
��n�E��TV�11�MTS_b�J���&�q!�dF�"Seo�����Dx2@�eB�b�Cۏ���y;<��M�s���>>?G]}x�O���ǫ�߼� jЩ
�i4��=��;�:���s׷�Ooק~8㏏���ϥ���T�f@�!��r!���]!r��%q��6�ˍE��OOoǧ����||tu�׌����c~���j��0(V�3ۥL`����2�O�e�572vrry<�M�ω��},����`=�;��ԇ������LJ)XT��LVO_�OOn=?_��q���>���x��]�
��>�i�M%@�Օ!����I˓^����������||}}�K,���VV����P���3Z,����Y�s06�fˣVz�7��Ҡx�O���M�q�*
#u�L@�a������#���nЬ+�bcY�*	�D�U�+�H��:��cZ�Cv��]k3�b��f�d/����M��&���(�G�R�	����-�jRY6�K՘��դ��Y�/���;�����%� U��cwyUT_�6����I#-��^o��
�iө���q'� q)R $k%"D+l��b��Oa��I�t,[߅��h-�i���#�äֆ��=�����������4��Iǃ�"��{z5}�QD�, L�j��硍<�rd_;3�g}��C�bˇ(}�}&��o/��	����Fr=斳'�1���ط1�c>ǎL�[I��y(����͊�aP۩�K3��ڞ�.�'\C�a��xph[79�LL/�zfQw�
/��|ǵ��C�raFqzc	U:٫���û̺��䇯&kU1�����!����cLX:�< �[�߱�3�i�a˶�MjFU{�0Aows�znE�q�"Y���Q�%���>�c�=�)����YN��N�H
�'y�w���L|�<�MU8����ݬ�cN #{�������fC�7!|u��Gp��R���=�a�z�T�C00�`�Toԩ�ߕ���{{'&�o�����a'"�N�W*�OYƺi���#���v��I)=?�P�}_��oi��z"�|�k������Y�P�}�H�l����m�͔�C����[��Qi�W�@�W�Yn�z��WȻ�ח.髑����/s�쀃[�ƾEF�qc|;�~|*�5��^Xu���o�N�&`|q�w&EĬ3��xoU���C⼔C����mw��(F�����d�p���6lf�{d��+��m��l�x�R�o��S喫>Z��I��ӵǷ(U�Ky�T�M2
_�x�H	7a�C�I�KR0����Y��L�F�����?[A������fd>=�P�ZĄh�t���'<r&�h�4j�������}���v7m:ָ�����c�`����4{�*WNr�����"��y��n6OmV?@�y�\�<=\s�f[Kzk@����6��6��ur�L�����9ϛ���f��tN�_e��r��7s8u�D8R��ۛE�T1�ڥ����6���Hׇ��_��m�:p�l<�uy��d�ǉ� ������B;�A����"oz7� �cx��O6�Q�(FtD�xg�̍U��_?4�9�y1���5?��y��o��׶�yHC'��ګ�΢Quy�6a�"�tI�6�(k�}�f�jm�NOU�����G{�dUJ�"c1�9-���ŏ�	j��{�S�C��;@$�#�!_nƄ㭪3t���(p�7�gu��ٿsSzTa�iR�C���H�����i[K�� !�q�PY����[���W�2C37�ÝYa��.$�#+^��gҵz�3'�=搚��Y��3G�������� v�a��n��o�c9H7���oɚV{�afzO�sLzD��}N�l���9�Է0-r���z}?�r�̙��1`ͬN�X�-����:s_^&GVGbgn���7��}�F�daG�0���� h���Y[�Q�ʷ2>���C$יu}ٰ?��>�t���H&�]���,�����y��cH�Ӊ�xX �x��C���On�� �R;�q�+/�����xm3#�3�5��P����3��;�N��_6���_>���<��:e%s�D�	�	?��/��ů��޸\SS0k]R���Z����-�KT���}4��	碤W@���O��M�d9���&<dǪ\j�u�8�[�S�'����4h����B4���P%��_���tD
���sGj.Ø��ӽrT$k{���
q}r�d���%v�[k�����|'��sL��h�M�d�t�R�[�?��_g׏�S��������C���y�⢏8]sdss�S�kz�0�Ə���:�3��78L��sG]���%��7��k����y�`D)l����;va������������9���%1��o���ryxa��뛳�=��;ZB�'��ii��
�ӹQ2�.���k٦�{�,���4[�.�T��C8���8@},Ň6�l�x>�Y^�B(���Gl��	��gP����t�sɹ5�i`�]ݼ��/���⧟��u�}G���,HQ�L-��4�	4>���� ���砋c5�x
��tqx���X�X����s��_[�͏�f�s�Lu
�����S4o�6ݼ��zR��@~�z���;j[����Q��F���;:�	\ZGͶa���˭y�9��a��^tP��2��:�n�'����Ӥz��ū����w���Ķ	H�T
F@H��D�T {��??�y��#�	�����T@�k݁��|)���I_.���.��[�s��ė!�R�yX�����Wn�An�nf�y�4�@}��ן�`j~�dos�=���Z҇x"ie�[�n`al�EϺ�@���$�I�M�w����c�ќ�}�����'�I�m�6�q�g�}�)�҉����]�\ �jܞ^!���)b?��_c��C�~��yb{�z����������Po<;�{�{��_���0����"�Q,3�2�z��������~�Wi o�Ȋ���ԯ�>h#���~$s _��:Ac��t���8�@�3Q�%$��LNz=]<s���{��Qv7w������2$�0�V��b'�w�&�w���w�0���v�����mwY�A�xba�a|��ˇ���i>4���zvOz���!�u�_���0;ψt3�mZZ�����	��y��w��G�����>��u�`j�!b��>O��	*{��ݽU���dFv���j^h=�L�VG��9��[3�@�H�s�^ j6b��S�	ۊ9�,i�Iw�ic��ؗ�U#X%�Z7�e7Ќ�u�����5��l�P�P��ty)k崶W=�i
����|M��$�i$!��mAE~��I��\ب��t��6I1�!Ta)4����I�6�t�=�R��܇��rvo{��H��|��Z�Yx����7#�Ni�A|'�(S�y��Ő@���
��zK�W1�֖����$`x�I'%��0܄� �7��VF����@�14����ݳ��u��K.�]�9�`{���;���@5��������va9ߠ���b!U[�m5ˣ'|�ȗf9�ѭ݊s�zȞ��<ٜ�iޥs^5��A�˓���j� N5�G������}��6�����6�4;�����T���6��>!.z|�ӿ�}�4Ta���>g����+��y�����lᬀb��c�F�bm�"m�-�e�K�7>�èˏX�`�cZ���K7R���&�}���m����6Z�L��}Ν�Kiz�M{:4�>�Lj��^?T�z�{��~�����i����,�Ț���Gx IN�H<l'�Ŀ��:P��O4>(�̎�^o6��41�->NX����Ͻ��z�C���M�����^w10�'؇Խ�,��ƦAuk�O�o�?u���� ��^D�y�De�~��z�gݢ$N�ޔE������հ���;"���Xy�[�%������7{�����b7�� ��ֹ��@�a�����>i���Gw��y�8�\�^�XOD�9���L�Ҥx�,�U�Z�$w��A�n�Xx�K��+X?�{�I0�E��I�k�ɏ{ޠ�tų)�/�ʒ��F��B8�-��
7�1�ݻ~��n�C�9ʷ�osr@<�;k/���o��yX�S-�+�Ni��^f3��m�x��a�.a��p��ϩ�����^kѮ E�=����!�`Q�Da�D 
@ �\����{���WX�b*�,�l7*"�.(��|x�F;BvwJ*<�%��j�8q/y�$!��d���P�p(�x�+��Y备�y=l��;0�EG��A:��_����Qu��ɽ�����.�����~��z1�#.����^��W��ߛ�H�"i@(�!��F�Fv�*���Y�����v���0����uY��[p��Z�滭/7���X;$�6y��`S٣��c�l��3y� &�÷��Zag{iH��?[�;�ɴ�ؕ�(�g�������f�ewo�� ��ś�"��y!�C��" &a��h��	B�/J�eB�{u�E��;d�e�����Wk	���㝻�$�2 D�t��W�>����^����7c���s[a�9��a:v��u���E�� �������ͻ�w�9��!�K��y�s6�����
-�N+k��H�u�֨��0��w�jw�/)�:滾�����?�_��Z���&^��!�������ʧ�k]��u�5ڥ�蝹�����ZXeE��8/�{Z��ܫ�+��������2��<�|+(��C���PYX�`�^��J)�?ʃ���ڕ�g�1�ѻ�*�2j�=\^^bKS�ظ<�r�^y�c2���(cH�7���Wqy+2Ж���>v9^�s�;e�
5�b����Wl�7���v�pӢ������J_�x ?� |�� 0�C��80}�C�"!�G�E�iBٷ�	r;�Nf����m���.:j��&��{9�)Ӎ.ˠ4�ك�!�a�EM>� �WL�gL/y��E������ǀ��c#�|�2֠��<Y*s]8%�a8�ܣ�mK0s��ꗾ]�׻�t�z#�� ���/���g�e�L�h���)���G�Pߝ�W6H{*�9�]��n�US�ִw��/�.Cy��}��<��(]�P�|�ľ:Ῠ?� )dV�`x���ٌ̚����|l���C�6I��̏�g��^U�����h�=��H�z�p+��
.����XɍD�"�Àom��v��{�0"+�Ja�S6���i��T8ݕ�mw�H�b�B��+�T<�k�^�������e���2W�b��w��d#�CeCR>�ҲH��ߞ�A��H8�]j�Q���gVD�<��(�?�49v"Y�����0Bow]Ԛa�����<�g�퉣g4q7'�Y�4M�2�#�z{�\y��6�a�^!����W@��4]QI�q�UÉ�f>y�~���Jˬ�Y��"] C��q��[p.&�}{�Ѵ�P��dD��G2�*s���Ӝr{��/-��%E���o�Y9�����6Q�O�+��t�G�.!r�+c@[��[�w���eLsIl���î�#�ڱ7Y��ᒇYX��&؃��m>74�r-��1�+qޝ��v����y盻�_{�=���Ad�H�!��"D � ����~���߯�F��U��Q���:�x/�9��� M���L'S�iL�π�Tof"and�l!��I�Jm�t����>3���6`>91��U?F�^r�4�9���i�� ����䮷Å�H0Q?��}����<�a�n棆�L���ט	)��G��lQ1��/)�5\��΋\������7#�>��q[הte�*
���4�J��a[}���8Q6�؃/GSVi��pm�
�����}^��5�P��ݳ�D���\^�B_�v�<��<c������u���.������׶I����x�>��q��K;ӌ�ٟnÓcm���b/*�Wm/ I�[��Z��9nž�-$�MX�a��a�vDı���^�c�-��k3:��i�w�g�Ki�Q ��
z�,q�����=�����θ2��T���2�7�8IY�.*	�� �R�]� Tn�%`�߽��^�#���onr�_b�X;[�tG޳�F�~�S�ڇ{�tyܿ�d����J�F<��=P��34�� Xf2h�6������F�y)~�&_�<�"n�-���mk���\�
���oE��A�Yx�,��|gً�=�	|qȧ@!1�	P�Z,X�٫�śY���ZwS��|"�sd�1�q�l��"�]�MeX��m뭒��s��P���s\������l���yߗ��&�e������5�pnf��Ą?��H$d$H��P� S�+�O��Q�� ���x .(�ql��Q�qF.	n��j@�\�4�<7�t;���-)��H
�,_��A��hf���m���@��k6Z�M+���;Ǎp���2���IB�~�o��m� O`n�����!d\;ôf�[�γ}wR��ý᧋s8i��d��ό�����8E�q�2w�-L����u��*<Gq��X��ɚ'����]�A�l<;���E�	y'6�q���<�6[i�g���/��ZB�׶�vl�����Z����Z���d�ں�"���KR�ǼD�D8�'����19���l���άp{�i��`���k��ǰ�<x�*�Y����2�M��a?ե��h�d~�B����JZ��Qn�݀ay�'ӓ�{Y��s��f7v� �&-o�a��ႋ�Jq�*#;;�oG{��dy�Ov8}k]�2;�˜���q��%�3* �H��b��K�/ۏw?q�$�F��������������ܡ>�/��H7�[���z's��zZ��U>�;�ָl�Ǜ~��W�yգ�ycM�D;qn��-=��K+�2�y��0/�s
���H'8����E.�����>�%կ�Z醻��X@���Ī*FV�W��;[�^�f��JS����2�J��nݒe�o�"�����]�����h[���y�;6@����n��[Ǚ�MTSFr�T]�Y,�m�c<{iխ��\� td$?��	P�0���U�E82�$�ʣ��H@� 	��y����߾��!��Jp�o@lO��ɀ ��6���{L��8aM���˽��g��.&�K�[٢���w�w� d7�9#`lG�fȌ3�K��KO�5��􆷼g�l�:��ȫ��w�A�'�ϴ��Cx��qh��׵���stF��~D/1�(!�w����x�6�ͬ��yۏ&�^�v2w�R`��m'9��4�wG��o��8��{�9��÷{���G��j=�����I�-o����<��a�0~\��/�(��Y�������M���vVjNG ������li���`�����3�]*5�~VH�^���i7�ۙ��l���s�=oە%ك0nznǩ�9�#"cb�"��o����L�c̗����>{�RxI2����cL=n4gd�f���T?6W\�wE%F�y�-�}J����Lz}c��5��e����
Ż��\�[W��S�7��|~�$5s�y��hs��ꙗf�oUȝ�n�P1D�/�3Yߛ��q_�>��"���(Id���g�z�`/\�4��y����;�G�:��?��U�������<�fXn�C� c��#^䵈�r{�m�孓v;�un�s�#��#�J�ؙ��Wxv��NA�Fz����%�dw�.^ޚ^X�:�b��7��.HT��w�'�{-7�7�9A���63�'C�)��1�hn�m�9�6�]�}��6'v�	zM,L䚻��Vl�U�K�w9v �Vk9)�^�3-g^.�v��wNͼQ���ژ;��˜�n��U�k7m?����
�w7z���M�}75����Lׯ��u{uyi�'ͨ�S;�ʕ���|�!	g[�W/V�n9��1δY�]lٽ��͖����+d��L��r�1}i��f�$ٓ�_	�����8�:�pl9Ǫ��ɴˢ8
圯�ǌ�	��j��a�= Ux"����k5V�f�Y���ى��q�A��j�\��#we@K���ɖ����o�7��wƋx�+S(=���c:u�+xN.�V�r5��F6��@7zc��6�����t<�,�76���#�7���q�庛���i!R���^t짓���:�uE��K�x�*���|�$Cy�J
��&:i5��ϙN��-��L��ffߟm�ήQ�!ruw@�፠�M��ժ\-R]�F� �|�_F�k٣�f�YH�d@}xW�=E��]�YO�����l��J&�z�z`�6v�Q̫Ce�9}]�ȫ��*+��Ř3|_�����]M�%ΛK����`9;Z�j���tո�n���<J�co�֗)wt���m�ٻԦ���L([�:��_-�.�,�F�c��ˬ�;;�Žpz�r�����0�d�B���s�q�uFO':@غYj��k`�Ze1z�ٯQj�҆�!SnCs��� �ɧ\2��Z���{+J]�  ݏ��QF���y�c�f�1C�m܊��%�lP��A7r�f��X��C�.���t�3X��3Y�������]�x�(�	���:���չzi�� D9Fp˹ĢY���y��0�w_�s,���INU(BJ��K�/�a	�Q�Hsi滹��w6�s1���[b��I�MƷ�[ @�b����,�ΔV�nP1Cv;-N����<�� ��j�Lv-۾�'U-{|��)�q1Yҧ9T�+z�%���0�&:�����uF.���,�B��׽� � U�o���8�1���ֵ+����1�9T]�|�k�UĻN�#&E��JP��9/�<����T��ĕ���PY����v�K��٩�O�O�����__^<x��9<��}j��m�*P�{�J��F�9�G������Ƿ����|}__e�Y�ȱh�Xv�*Ŋ*2_l�
��ck<n}����������>>����x�8i�9�Mb��P�2J֊��K���Q�s����==�������|}__^<|�f}f�m@�b`yh�Vyk�*j�Ī�����#7q��}g��^�|~8㏏���3�g�����V�m�ib�Ƹ�A�
�ֹ^�K�C��g�&�'�S����|}_Y����#y���g�����4��XV�9h�fR�3v���L���Wx�Ǯ���A}�i�Nۖ��(��R�%UB�Ҧ8��Vf�".��$�Y�"Q�{��*-c�SWˌ�K�VEa�H�F����rt�KSڬ�ӵˍ��R�!X��{Q���*teӳ�ut1�u}���&v���j�ͩd�� ?pʫ
0���"��`�B(# V~H@�}���j��9��>�&��β.�@c��AY����D4�=�Qbo��utU�nsU|��c�iv��C=����;Sa,�x;�!����n��ۃs\�
9�xc���/���w�7z���w��>E-�/YʐI)���>�z�y�e�P!����Rl����� �ήq]���#�Z�~h�t�ΏZ��s�j�,��]��=���B���(���a��w9l���.��pH4�AfV�G�\�R�T�R*|Γ$X� ӌ��'�d|[��Z���Dl�����QU��y�˻��J?��b}ߨ�`�H��y�vgʃϭ�z߸�`��AU�%�KU֐xvq��^w��@1dw5b��C�g�7EtQ��C� \��6x���i� �նM�݌�щW�=l��>w��p0���?:^U�_�c
X��~����fF�$<WNӑC:ion!�d7�o�EZƖ)�ßW�eQ��!����ܙV�䰨$�4���h�Q��*(Oc$����_r5������Nk� �"�@Iy��1��@dCy�C�y�G�����g�G�~c��ü�皲,nL�����j�9蓏k��H�v�X�'#��Uc������Ȳ�N��'�W���y��[����i��6�o��e�e����fvt�o���ߜ��J������+���0��
�« 0£
��� �$  3˭%|�g���W�C�T.~C�<��dT�(��D'�S6� ��W��2���V��+Z5u�u�Pe��g�`�5�q��6H�	�~�%���`�E#��K1f��[��IL+'U���6�#)�Ӏ��0��)y�G�$�d�^\��`�T	�_��胉��A]�B����aT\�������d�����lԜ�q_L��W�'hx)	|	�[���?E�-(�S5�O�~57[xyZ�yᤁ���,�T9�j�&���ߍ���*鰋�aN;���kɮ���nG+Ɯ���8�c��x��6��G�N4��4�]3����lbg�
==}{�3��U����W�%]R�k?� 8�M���ߌ�vf����Dx�����V�!{�]�[b��H�I��)D�o4��i�`���a��u��>��i�hD��iy�c
�X$%����z_��^���S��;CG23�a�o^e�g��bޝ��Dgu�i��2-O ��z��{&m�m�{�<�%����ut7�����y��lv�a��}j�G��ߎF8]��}���?F��Y�53
{�(O�x4�tT�4�O��\�^tg�=��b�(�raB�%���6�$�4�Y��^`n3��>�;���K,�����-�ӷ�̜�I/F;�M�!Z��y��~�8��h���ȼ�4��]!�m�yί.ToD�n��_t�׭�
�d��jZ����P$9�M���a���e����$���A# AD!��x2�x2�R2,����w�i���<����g6�:e������&�7���8�|-���ώX8���é�B���{UH����u�t�a�����i&�`Ƣ�5REz�v�v9\����!�F�7�x���+ְ�^����qŀF�?w�@>0�ѯ��4�Zg��L�g9�O��La�؜�� �_!�����ı-�B�H/�bFך3�(_\X��N�­�k+���s�x��� ��ts�޿R��^5~�R_�0�D��s����"'���ƨZ��˸W5�����c�57 �聒�H��7�">3��dp"ơǀ퍝���H
�̹k�u����m��pxjfs�06��DW�~A�_D.�����B�d� ��Ƚy:mּ�-�817=���]���ݠ,�t^ʂ��=�o�0�w�;��E4{���!�:���	\��%�C�H��ND�/O9��;n�ڡ}W�߼��C�A�^��dP�#�ODW����8L>�lt�h�7MP�Ӥ����ŉ]\lk�E���RaC���d���ȕ彨c�����6<7��)�1�ۇ�3Nf6�T82���n��Wg[�e��s��2�ɏs4�"y�{|4�����[�m�1Gf�V�V�����n���U�]�#;K/���d�0vr٩ ƞ�W&1qs'�n�΍�_���0/%(^ ��� �h�` �d$��"��}��߿_�_�'����_[��[2�c����7ka�8��%����ȣ�'^z�"XEuB�����N���|�zy�kO6��iÃ�v\�?8��>coE'�c3h�����G�9wy�rf`����oj`�KYq]�$�ti>5D15��7=�^ ��n��	o2�%���4ތbO�r,��!���k���ũt>^����hlLum6��V��^`O��J,�i:e��5C�:!�
��a`>�~�E�˧!rkn�>#+i^-����NpD������;�yL{T�CiI-D��� ��"���͓��Ph�g+~�s|9�KBu� 	9�)LD�{<�Q>�����p;�y��7dA��̠���n�t���;ݏ�j|��E�"���=[x�Q-�)�o���͌s�)�]�~xI���� ����u�x��g_@�>�^��5�_x��'��|9_�к�ȥ6zś��(�s�2~��_��iO��Z�U{h��ߨ`��h�����*h��Y?kUSW�������g���/�ʚ7H�3[.��=������Ӈ�n��Ę�ӛ��ɝ���������r�B�ax��0͵��>���v�u�&�N����}
�/��լ�F���_a����:�k`,c����r���{����a�9
�aC�!A���(pd8#P%����;{���m��7V?�J؄|��^�����/�K|R�|F�ؓ~A>���Ơ��?��bِ㫲�E��:LRxkY�l�R���<k0q�'�}WE����,7�:�Vu�����/�\ڕ|P�WD��v8_'ӧ<�k_y���x�^�s߽��(W5yM܉�kj5n�����|�����ů�|qQN�n?x�1M��m"��4�A��>$�ܮ�Eǒ��w�,�r�bP�C���&�8`C�����|X����=�\��ˋ���Ϲ�]��;�w��;�N�;��L����s-t��c=|�Mx��<	�q>���7�MS�+k�Ʌmti����gx����By%�`�v<" v��v{{mNǻ�_Z�-�~������8</�@l"�f� ^�73����i��y��
!�ZO��'G��c �jj�|��̉m���G8?B O���+)�@�j�g|�Ƀ��m��D0֠7F*f�t�}�����@�_9�A���x�g�5w��4�<2���JwP���x1���hm��G?ջ�`����dY�n>��ݢS�qHt�|N)z��c�]��ѝlV��H}�"(���;�[aչ��2����0V�MQ�p�[�R��oe[��SJgP<ұ,t;����$������	��2�!N*�"�¤0�Zi��s�g�ѕZC�����d|�0�5�Q������ޔ'�{�~����/�_)t�#�u�O�i������<Ͼ0�]0�&���!�8�W���'��1?S�iҺ�a��J��u�
�1$da��h2���¿A��vW�J�4�b�?[�]�<Êϯ�7�k��g�V�e�����߾ט/���w�����L��f�$֯oB�?�+<��E�����Y�-���e��Z����u��R����������O�PZ�����M�Ur5���c���j�Xjf�e�{wpn<pq�c��	�O96gڝ$�}|��n�VT O�*�Z������/�'�βf��e>��qq��4�x���胉�P�J$Cp���x���L_��w'��c��qZM��[�aɲ�1�YK̎a��M��ZzO=KRMO������u���@���&���3{A5���a����`�y�(Ԋچy�S�� ֛́��[@2���;�[a�	�_s�����'M/s&��@?,��߷�N�S� zm�G.�{Bz
؝�[;�w��X�$��k0f����];;(��y�wZ'�g�]�{A��]mYZ�D"�A���2� er��>�ng2j�!�4eo_���r�n7����Յ�Ot��٣~FP
�y4�q/�:��/lY��s9˳�����k}/��٦��$�IT�?	�Ȥ2=�u)��"�@X�Y$���Nv�x�ݸ,�ZX� �y#��ZpۯZߞ�Cs�ꑺ����Y����.0#8���y�2xن�K��[�OtA��jx�#L�`�sγ[Nsʎ��3Xe�h!�	��|{��m�o�f6�30PՍ>���z_����������P�\��F�X��(.3
�����v�U@�o0a��(�fc�Sl)4��=sH||�#�ɟ��K���ZN"L�S��Ѭ��x��&�78�O�k��p#ZE2+�1��AN0��X�-�N�d����M�4�\��Ӭ�>�����ɿ�#�z��ߕ�o��G��(��ņt�W��*!����(>A� ��
�ƹqia�%ጫ��X F�����^<�g�kn1VYg�h"|�k} \��y(�z��x*ݩ^>vi��,0��7I.��WIƟ������+E V�G�~��~!�S�7Ʀ��Ȭ�=�����G<��F�(b-'��t��3t�^G'գ��6�1�W����U�
�(oW�ϼ�c��Q@��o�����"��A��r���<D�����ɺ��]Ǒ�۫sT�\TaRGX�hǋ�1�
#�ֵ�<5�@�i�`��eak���y ���.�#�� ֧˸4�ϓ��q��g1h=���ȣ�V��!��o8���������}T���-�X�؛`��̏� �!�g�'1 0�� �x9��F�j�����Ĩ�TD(e���:"�!P~��yCp�~�l�,\q��?3� �>�4��ڍ9c_,����`b���[�ʷln����ocI'�Y'9�/�Qd�ʧ����L�vƧ؞�ر��N�ͥ"�z����;o�>�3Qg�	;���~7��}��j����{��n�&�	�c��!��-(xm+���K�5�ϲ�A�>kܹq�һ��UvP�@��z��������o��{y���,��';�ϦN(p�ʻ1�����s+#�" �v�{=����sY����mǽ��k��o0�]0L4Cc6�����fn�!�B'?������@ "<�F�͜��'��Y������'y��k!a]!Cq�
䖹��z_�mz^ӌ� 	13�	~�\�����h��f�q��$2�@�F�fg}ɟƺ��Ô�^>�!'���F`�f��kl�ᦛZ!�),�ȶ;���a�?{xt��mr�{�`��t3�[H�
#�Dr�d^�,����ë��k'|�k����EeC�3/�Hsy7���k����ʛ�(�I�f�)PǶ��oX#N����J��IYJ+����4�p���1��zeDO����Ֆ}X���i�n�Yyܥ���d<��lr�.��"�Wb��mM�7bd�u��G�R>�М$I�� ��&~�9�?}�k�h��y���T[ϙ��s}�'�a��u�}�!0gD%�zB��9o�o��g�ϼ��L�-+���s�^3U���}^x��t�T���������~}j�=$�6�oz�L�ny_��}g��jg�ba$���E��c�y� ˘>y����	���af͆����ޖ�^3��0��7�L��kn�w"� ઝ���]������˾=���Z5�4�`�2+HՃ�Y�7���s#�����G��C�F˱�-F��oAsښ��XX\��G$�b�O_��3� ǩ��Y�ek�(u{���_����G:V}^*����-��/1F�������h~��1����q]���d{���?5���	�*�v��A�����!�x�,U��_�w]�e����Á�-��^��^�L+jO'��é���<�
qtq�w3�ߞN�ծL��>m~���M��Ip/8Rׁ�Ưn�!���0>�SPR�\��gVԼU�;b��a4CyS`�]�}לbs�`�����s)�o��DX|�X���hx�Dò����{L�[=n;�z��i������1��N�u����GB�N�]�m$3�V�˽?����ٞ%n�@5�#[͝�����$���s�	R3%l;��4ow��W�:j��n�Ζ9���̓��Mn�?�S$?��9 pnJ�`�H�	K�cj���_߷翷�����P���ɵ4}�{�y�V�3�����ȝ�Wz�x�ȹ���K�nP?=��YMW�������f*��|�����꿄xg�	�O˽��p����}oz�_g<�\��v	�"��l���a��6/D)�	���"'��f�p�uJ�U��Dki�?��p箭�j�����4�Dy��l�I����k}���	�o�:%a��J��b�dΰr��Vc�yK�8La���C��4�k")�G�]�a�8��kb�Q�EY<��f�π|	��l��z�7D��!�'�њ�s~����L��hE�����Q�Mڤ{ņ�g��y�����V��:l���?�~$>��>�E~U�b�g�P��#]����E���?N��:f�����UR�i�0�	X�C�`/����Ԃ}�Q �5L�gށ?�� _b��pOwA���\��!��,�Vě�/#ׁ�O8E醺v�0 %P;@���B�h���g�g������n�G�ǋ�� �ʋ ,�/���r&Bκwm��{��x�/��3�e�������S�t��Fu�͛�2����+U��z��##��H���؏D��qʗ�f�4���r�}LWT���yu5�����v�Q�*��]Vƅ��o��/���z9pKm����&���j�C$�<#�S,<����+�X�x��b��g]c7o����+v�8���Ţ��V����}��N���iq����U�H�B�v����,{|�BL���DiY)5��n��	���6wJj��5rw�J��j�v����L'�b��m,�]j+ �e}o�8�0�ou�Z�nE/�bu�c���н��[�/��;�hoM��X.��X��[h� �O��93r��m>vӹ5�}W:�O���e��ϻrb��:m�H�V
���/��0�����$f��C���Z�\���5�u��oβ�N����go�eqD��f�\�]���M(6�}r��[P�<]�	#�ݩiZ�ǮT
�G�<�����j��gK��Pq>�un�㒐��n�qU^�NLa�6,��xP�8����P&@�2�#W[2�b�"��� ���>j�*⨻����r��[����[�dh:z��ծ���yo>/V[FmӢi�q<W�w���H�=�Ī)���R"�b��m�O���w`Q5q ��"j^WF�"�5Ǣ��ʪ�M�%ܫ<Vu>
w2�\9�:X`�EU>ȃi�r�1���2�XW*���mYg�Sn����A��չy��JUۙ�Ц]��b���wdG-�9�W+o6u��%]ZR-T�9/#)i|�9!�l��Չ��m�1*x�$_�|�4l���g)�n1��d���]"�æ���٦�⏌wQV������,Y/vN���ϻ���,Ɪ&
�qg�ԩ�h��u�9A�8�jɁ˙�P�y�i�"wE��(�nm�77gL�25w@�9F�}O*�7�کf#��p>��A3{��i(nር�ξ}xF�8f��"+�-��7$���ɪ���FH|1�>PU�\�.�y����;!BH�J���m�D�z�.w��a֓������ݿ����������c�^+1�L	L#.���E	|�~|Uɡꋬi�t��e�	e���T�̰qd$��SY�q�]���SU1Gy�q��p�e�d��b�ΨN�-B7���8�gXT�Jx.�J��;kfp�vT�	�-��ǽkfi��̮'Se������k���J=δ��2�{�_��k�:�43 �jۛ�-�¸�c֚4jt�w\7:i��\v1�;+��ۃk�̻}p\�7!nS�*�Z:�c�������-<�J�]}Ń���$��n��a�HS�!�&�v<ݐ�0H�*�0����="�f���6I��Q��8��A�v߮�\��L�d!NE�*gȤ�����(DC��I�h�D�dJ+BF�4��<�H�0Uf�MC� ��^F�!Mn�E�X(&��tbL[X�$8n4�� �ar��,EH�Ջf��
�j��B�]O�̙57<��M�O'�ɹ��������W
JA��莹¢��"�T�q���3&M�O_�����q�u��^;��θ78��ƌ���r�3|�m1�3e���G������������8�:�ϯ����1b��Ь�,4��h�ճ��̙79>������O'���}��ߔO��R[Nn�:AUd]�$������<}g�����_�8㣯�����A�O:%��e2�R�"6��o��((��;�FY�Ss������8�_Y�_}= m��T\�:#��kKT�r�W�z;�1��&�`q
";8������!+TQF��y�Ȉ�̵Klչeb�Rg�2�m�DTA�B�Xq��T�`�d�q+2�Q*Tm�""���R����)��#���p�K��50�(4�8��J����v��d��ɺv��6>�v�%��.g=ޥ�Vj�	;�:t@��zۏ���n�Z�����[l��L4�-��A	M����`N �M�I�E��1��!�~(��!�!��V	r��)�Ͼm��K�x�ӑ"S	u���=W���E{8�-�:r��DMZ�T����}x��+��s������]����c �������6]WSn��ȋ��w��;����#�����{oG3uM��c��o�&�������+�)��o
��ݘ^b���h|��m;�tC�w��N/0f���/ѹ3;�g@s�zy�/ǋNM�U�lh�x��y��'���G�&�Hi��4`8���0�;��/d^1l{�C<0%�P���2g���������3aH�EC�#�I�g��^S�l9߫�C=�C5�s��n�t`Cgó�v/8O��4�?��SL4lx?�a����sW�'zj �ײ͙�Z|s�^�f>%%�p��Av�����6��a��I�js��������z+	�ss�5coT܋*��r�v�;$�XJ�up��>-==e��d�>:�E;Zl�q�p�)�Q}7�k��7�;�������?{��[�vsgܹ&�$gWR@�H482�r��ka�~�5߹�Ri��V�y��G���<�2[D�Ik�����;v�w�V>1�,�}�C�@,>�ӭO�S����i]6^0��&/5����;,%��yC�o	Ǆ���/Klgj��כX������zSy�I
V��Nf�9뜵������H,�����A#$a9D�1�{�~���~���n'1(�ŀ��_l!�葼�N��W�&�i�\j�Mωq�mWMU�@�o(=��ݖ2 j�b�k�@�}��9�+�]��b@K��DI�;�{�^f$�+�ǡ�3�q�Z߹�� K�r�5�,��%�06I%ب���B�I;���f/��Vk����rig���XO���[������[��F=m~!{X
�E8����5r׫5�L�r7�7$Mz���3� �w��y��!�h]�?�����?.��oD#ٌ��Zy0ά�I{�E���^O��ES}�_�"}޼��Q~�c�`}�f{���P[6gY̽�c3Mhu�$��$0hw�瘎�v�����ͧ�}JEt�͟;��\ȻW�g�v~~Zi�)��<&6`�<��v��L�G���͘�dsϵ����8�k#�f�/� mv�z}���j��x�����a�eD�G�{y�;u�h�ǹ��Óܲ�dޒ9s���aeS��{�Y��;�S~�Dx�s<�|��v/�y����Y�:�ǎ�d72>�;ӆ�5�cQ�jĈ�=//p��ۮʺ.��ݞUl�����_�t׽IAF�q^x_����W�.��޾Z��� �&UEOo�.v��iMBJo!9�:��Z���Wô9��Q�ӧe�wF�6��Rt��2�f�\?���FD�F# ��1$0� +��ߟ_���|G&��=�m�6y��g��>n֩�> ��O�G��b�q�����r�l�^�Z^[����M�4�{�h���YC�Y��Fs]4s��e�ќ�2^��Vj��c�>/�ދ��Ĝ�T%8`$�Q�^v1�G�V�|�9��CE��M���L|�Z����VH�kTx^_�SL5�������� |~#>ů/�߯g� ��}w�\�b�Ŏ��bͼ/œ+nx/�#G��,L�������}�_5e�O���r��P_$��LY~Y�U�L�LƎ�`��;�>�2-��Ƴ:��#On�藌��բ�	���\1�x�S�s�,����EV���������i�Dasv�fhP��f����!~��6G���ޯ+���2.�ZHS��߫������g��w��z�Y�S]<}�Qwh.��Ũ�hb�?��$CI����L��=T������:��1�0��qOd�U�ۑ�n��f8�|�"}�@x���ώ��T��ܹ�I9��TyB~�_]a��+��=�v�	��l�ū��wn��v��:�vm�o�.ҭ�\�)N��۵�130�'h���Zzr�h8;r����e�+s��}_��qx12��C��-���#ѽ`*K	"���z9��"�	����'榾ˡ^�P�����y�Sm�
P�8�0i]X���`2}���.O4�c�$�>�i�7��};�uy�n6)�שآH�k.��{���:�@f��+�fy�d/�I�Tl��E�ds_�^[�;u�ÏJ��`l�7���q��ƏL���3;iY`bE3"�6�@���׫�bʛ��[K��+a���ȑ�6��%�Ȅ�N8���i���bCO�rY���:R����dp�,p�.��mc�>�u���#c��oПԄ=��'`p[��\�J7�iU�Og$�NI��E�	��g'��A�4�/�N3޿�`���'�K	��KN�C��;��Ũ<���Pn"��MtL]2�s��Ŕ:���+;�c�xn����rT�ܕ��ጎ�x{�^���8����>h�XC�g��xZB/+�w����b�P����;�?>����[L�*�AT��r�3��n�<�-"����o>�xW����m�~x�]�v��7bi��c�Ֆ���`V�f>���i+�9{�G5E���+u�hVJ���x��	l�8t�`�2c�u}�M�St�9�X뫾t�y[�f>�ʝwݦ�T�	�v��]�"��]�<��rB���2�
"��H�6�!I
��U]]\����u�68��$0�$L���a��V@�ij�/���x\h�bX�bı�}d~f�� �t�u2�kJ�$�CoHG��S�0"w�q��b{�қYo�����Q������- �}�]�+Q<Ÿr����s�(#�����Z�4[���7���H�9)�u��sg-�54�	K��if�����B�^�N3�u�w�=$"2�5���z��p�"o��R��ϔ����W��j�uV��~����z��K�D��R&�^~� V��t�xC��g����;�Y�f���߮o���Fw**=>q��|f/�\��M��!������4�y��F��nJ��mG<y��	D��z=[�"��i�b�5Efv�d%��G��j����Q���\�t
�}���4��͇��gt+l5	� ta���<l��+u��n����x�+9Z@znm���*��3�w�`g���r,׈��#������L��x�n�2��dxc{j�'(C�0`t��팛gv��'��(��Ϝ90Gdi�s>�[y��g��+>�����jeLb���7���|N�ʸL����@^�ռ���)f�|�L��ur��O�w֖;���(�,�tgu�S�&�w`��x*���v�U�������R;N�ܺǮ��[d9�r��q�o���(���?"D�)%#=JD
F� ������{�:�0�^����i���?!�Z�A4��*{;��"�h��ϼ�S'^'Wm���@��L~�JE��`����(�C��dri�G��[K�g��G����wz�%��
l`�ֲ�//�g���z��3�Z�x�|(��e��~��g�ɿ�� w��!���j�{K�H�WW=��� ��lƅnlF�D�Ã��ݖ ���uQ��`��%�ͩ��l�3�V���sz����(r� �l�d�X���-�B���9	m�\�v���/�����;o�<H%*@"}Z@GA�H�����]�������k�.�F�v������q�q�
@��w���r<�qNZ�z/1#�?P��T�\Sf�ixN��"���xZ��b3�Ie(�ds���wŌ��(�$#�$���L,u����[h!�������<柒B���&{ѕ�꣗{���Z��f$���	Q�w�����߼��H�lUl���R��8@���~�!�|�{#��T�밺p��/�)��&K״�R���f����	|&�d�4��a�6����nt��Vr���y�IK�b�Y.�������`\�𸙭J��z
��Zg�����ѧu�e{������jn�'q���v��%�����K�����Y�V�[��**����t�m���+�g�l��'�0��2�a�����ٽh�=���s����#��ͦ}�B���\���w���f}���c�c��W�7q5o�,u{�4���a�4�p~(c����V�� ���(8R�L?l��~����Ǽ�M\x��w��z�t�"�Y{9��?cmw6.o>����v���^���R�S��b%����$��W4ac�6�sG�?�u�[!���Co��0��{T������,ؙ?a����� s}}'�b �����Ŏ�v��l/�T	��(���������̎sm����v��7�؉��gI���辐�hD7��o�މ|����ۙz� �pa�Γ��[�.J,�I�!10�X9��!�_�:Twf�5�]�2�w��)��;�L������i�>�ӑJ�&������!�Dm��nƂ�y�7 ���?����/��D����?/b��O��
H�@@�28�ǹ�t#��.���κ����}p�%�0��>.��v���(7�L�9�(si�ja��*E�>u�������5˝��])#���o�:PSn�����t�.�a���_6�3]�پ K���2*ɛ��.�����;w�gUkR\��c{���v������bI�����z��ѫ�(�3{����vs;a��D-%H�"R��x>�sF��a�f�:���\�E�)�y? �t���~U UhY�Ck�rU.٪���3���m�g��|���7e�&Ʊu�0���M�~b��g�m}� ��l��J����@رHW�в}�#���r?ן���3덩�F��od�k�}᱙���6y���\ƈ`���$���-�2��7�P��.�M�C��`�.[��ǁF6���:�o����}0�ɂ�0�tz�YF˳�I�G?��T�<Һ�E�{˝��<��a����D=$/g�F�c����ǁ)���е�!�7=�y7Pc�Fmr��DS����2�r�o!�D�yC��0׹�p�L3O�77T��Z^D餕�t��D�Mö�N�p'��#�;OF�c��a��C�Dq��3R�q�Yϒ-��s��3�k-a=D�Y]3��P�� �՞U�O�;Ϙ[���C�7t���F��4���n*��	�Xg2�>ֻa+\�Ś�'-�Ń�YCI�m��-��	�	�	Gܘ ]�{Kg��h�HV�T�K��J��˭��%��i���z��/܍e�z̨V��+tH��\�%�\l��J��v��u�7�7Y���Y�
�ʷV�>�ӹ.1��˰�-��`.@#Qk�Ը�d| �Mv(�m*i�b
�D�n��T�neƦR�s��#�%+I��դH�� U�oγ�~��ѫGU�q�������ݯ��5�>��'q����`��a'��i��:_�[>^nUvL�	���W36�i��D@x|5�q `v�ш�vu^�\�B����1���k�U�_%�[�\;�� h[��,���uo���7��h�X|�Y�޼$�4���s0��¡�D=-|�ܤ�[������k�'*�.�zx�"?L1ۮA�˚��[ɑ�tG3��n�rKL�����ZI��#�~����\���ƶ�}
o��T�>��,� ������&�����{ET{����ʧe[�9�
(!=�:rAvF��D�?*g�g��i?�W5��4��?U�|lW׵��w�H�@ws~�07�0X��H���G���Z���1}�(_k2<�e�$��H��4ޟw<�K�m�)Jl�Tγ�^t�"p���M������c�P�Sl�Q�Hg៳�Ri{�?|�w�A���X`(���/�<xZ���O�������P���Cy�a�&�)��Sp���7�t�Ͼ�qV[9��$B�~wC����` M8<P̦P��UM�-9�M��~a��9c��2�U�*��iQ��=Y��ky��1����+���,�m/�z�gͭ�G�7�
C�s�r�ӂe��;�E�Y�19f.�ՙ8>8W��Ldt�I��,�|��i?��D���RZ.������%4k�d^���Gu<Ψ�s�n#��G�E��W?���x_F]�v,��v�z��<0׻#e���~N�?6����X�j3��$│��re:�F!EE�nl��v��E�Q�Թ�^t^��n+�2�����ak1��%��ތH�X�N�c|4#�[?����Q+�9��_�N:��I�UO^t�d��c6]�{��fJ�f���	a�`5���#�X��O��Ƈ�Lؾ~7Mg{v�[�a�8���=�1k9#��'�w���i ��@��1��I��&�i�mo>Er	�N�ّr�sM��{�[;���{��l#�f}��tֆ/��L/�W���|_��8>�/���o
t���g@�^��[jl�+�8�t"A2��D�@'�׉08�Q�+ҩ]� b�����!�<����R��At[H:|`Fs	�%�Q ��sX�ͥ[���M2])��~*�e�������c�z,�Y�l�_9�o����AR�o���=bɊ]��>{Ϻ��ǆ$�dA�U��ө��TqQ8΅�WA�4��yE�C�����e'�=��[���Z'Z	<�.V���*}��LSR|��*�]��Iu��fÛ��c��,�V�\N��<;���>e�B��[��ޫ[��.ǃ�h̻�W	;P�ϧ
�w��'���U�;c�F���f�|*G�]�*[�R��QY��to89��(���)��X��8���z���u�
5:��Ԯ�KH��t�z�|v$U;�������V+e�dK5��1��_ܖ�1Ԝ��:,h�hN��UJ�'�iT7�u�<8fJh��eU(c�z�997�KN��;P�ɶg���!O9�p&jY��\3��*��Zv:�{
��2�2t�+X{E]�5>1ޚe �xھ|�foG�0���}�Z��gN�z��n݌ե�����k!���r�A}�5�#�N�e:��G����*e��I��s���.閔"Uۃ-�� ĳ���)an�R��秜0k�Y���{v�.u�G7�YV�@�J"�TFm�U�4p���;��^�{�=yyD��V��m�ov�]7���kj��l��Pn�� �lK�ꘚuf��e�S�b�vf���u�K�]ƝH4l�� �^��U�R�h�F�6���F9Lٲv�x52����wFuod�E����zA��ƉԺٻ*��Z�;w�\xV[�2cʫ�R"��l�bi+����Me6�f/��l2�y�߮���@��Ğӱ�!�P���M�J<�Wfe��֟d�N��̌է��\�F>��M��ة����d�L����Ў�SJ�a��Y�YPs��V�2AUDV�9,�7�y��uG�/'��E�ۣ�8v�lU����ۤv�5,�u�K�ޑ�M�-Z�bY�C�6��Y6\��w�=��*�C���!��&�ˆnVV�C���	!\�R�ڷ��7z��Y;[%��-]��3 ��o��2��K&�[�GᏵ-��guC��'l�tz�=�I[,J-�X{�m�u��Z����>RԂ
�كd��@�mF�7:�=��"�*H��Z��⌛ vRa��Y�n�gj`��m\��IA���;۳�՞J`�]c�F�r��˦9&�ň���'�'|w��7����,Q�����-WV����A�$ ��e���9�Q��O{vٝ�f����8J� �G�'��k���N��һ�YM��F��o�Ҁ�0�-5Ў��Mm��JΜp���s�8_6\ռOb#O�j �^���z��' �!�<����)�j���tpה�Y�� O{ O�'���z�e]:r
�5"0)�cO������������>���>��]�PX����T���F��ٍW��XTwB�"/gіd���~>>>?q����3��~�]E7����9��f�ՉXb`1Ɗ��e��3&MMϧ�ssss����}}f}}=h;9ģ��W.�$�_���MR��iJ=i�*�,�*XQ<�Fdɩ���������G_Y�_ON�q�6�s��Uv�"�߷jtO���^%�A��T�EEթ��ɓSs�ɹ����>���Ϯ�T�q���p���)Ơ���YL\J���y������U�'Ӳ̚��NM�;?q�>��>��mȚ�{p��E�jP]ӏu
����/�Q/���(�L�!�X��*�F-j.%�/ut�Jݦ5����(�[���
1����*�ER*�Uq����)��Tj-`�Dc*4EE��6�i��mR�0��1�����;�y��邑Zr�#Kt��r�e���Mq;҃��/]5�}گ�_��x��<�"~i>�<������o���?U��h�5?���������Q�I�ndIq5/ɚ�l��7��b��2���'�8Kdό��R�\��G��mU}:�ak|l��6R�.3���o%�������Qfs$N��i2��`6L�;�zh2z��C��]ؼ��k�gsތw9�<ЙMڟ)]7mw�E��nǔ�dўj1�k~zmo~�B6�Խ������E�I�p�{"Sz���ZG6{[�E)�:�Ϡrڛ���Ͷ��w�q�r�B��C7���4)��{�x��C҇���j�)���%�����7�����x,tw�PL8����l��X����E��֌�
���1Q6��;L�-�dC����g>\kr�\;#y>�M>�<� s����뱙)�Z�؞���ι���=I��,kĀ�2,�+!���/���ڳckEp��渜m��0���
x��������O^{�w-�C�Q:�f4f�P�y��tܙ�B��3v�pL�nd{�/����GC��&�U���3�����:��i��pS;ߞ:+�V�7�e�od�r{-Z�ؾG{����V^V/��j�N�\/%��&dL*ۗmk�k��S����g���?��m%��-`��!���Y}8o���.1�E����+Y��h[	K# )4�I�!���|���l�5��yS1潁Sm3�J�[�/K@ƲlG�vDa�ZE�cT����%Y���iI�*G����	��r��4�CIvܛ/b�<���AlցmGAnɳc�L2[��F����tY~�\K�=��͇��� ��*�SE����%#������w}�7ڤ,����ct5��`.O,�[�ؖ�[�N��4�i��iD8[�s���cDc����J ��P��FMtk3@�t���F�u���bF�1�X��\�����w��j�"��|G0�~y|`�s�k;~��>�?Y�g�m���	��;lc�h�ٽ���nuΚ<G��K���0N9���i M2!�0��Z|�����s]��b.��V��]�J�F�&=���EE�ݬ"��:��1������?��@�e#'"�g�@'�gg/���p���4[0���bL�~�i���_C�.x����/o#���]��϶v[���S��jЗ��Q�~�q�z�$���t�O)����X:9^��XL'.c���4��q��cD9.z�a���$�@r�,�#}�Q���Lw�m5�/�q1/Xڮ��&�JO]A�i]�Љ��2����)�pj]��Τ���a8�H
j*�Mre.��֓`��"������Ku9������8��{�8rA%ك�rY�n�m�u�����
ˑ��ڬ���Yg�%��e������@�g��`��w7l��7�3H �#���Ӳ��s����Oa�	��bf��K[��Rb$0�Xx78�o�n�:���ChP��:�X�0���"F��R1��Ϙ@I��c��޷-G/PX]*m̫BnPBh|��oe���|�+��ő�a)?�!1fq���l�u9����C��/���ơ���������.iVC�:�c��.�Y�`�|~���HZ��Os�5��C5��,�?<9$��c�0�aGr��yn�KRĠ�������kש���/@`3��r�@�0��D1��"��k8�U��W�Sռ�p>��2���;_{̃���4&���.��8��V�y4�<3Ur��6F*�ɣ�y��Ar�q,$�#�����X�y�ϸ Oju�Q�m�W��liM~'�y%��d�~�S��o=�i�l����1z,O�	�Mz/h�M����U����͎�q�n�ؽ���Ce=�Z����U[��W\т��@;B���1�U�W��RN86�W��]�8%5�v�`^�]�;�H鵆Zl�4ç`4�W$r5kqG���(2	��)���y�w�������)(V%%H�>�������^]�(�¬�4����,��k��em�Hs�]Ѝ^�@PŐ ��C���u[dL+��6�ԷCC[�4�f޺S/\3.7�"��џ]3S�J�~'E4[��8��<��:i�Qg*�����ȼ�Vԥ1�_u/4U��s��*�Nw1C����:34����R�k���嘱�&`౜�h���
i�֜��2��1s}�IO���H�ov-�[������w*�u��F��Ѧ��w�j F;�Wv��>�!����� ��t۵�q������9ՙ����,��>ۨX��:�K7y�Jl�;��9�4���\�EQ`n,TNǧ@]��2�n]��������#�����gfפ@��"��ؽ����l�Ƨ����V�[��5m��;�����u�.�Pe9���P�������t����X8ebn��*]�ّ���Ӓ�| ]h�'Q��9��k:?+{fb� $L�����Y~?��y'�6�'t+#U@�k�+(����n��kf�
�Aաۭ���-�㦺?=��y��5�'���J��R(L�H�IҒ�AwmH9��O�م��뭍��62��ئ�w)|�vR-������x����^�����ZO�����;C��+�lD�sīx���-Jx����u�za���Z��vϜf��v89g���L��k"�K��q��>b��y�"�	�z$���0m��v@�x��.�ŭE����`ѱ��_zĔ�T��F@/ƛ˞"*f��+^�eI�����E��@YuQ���*:Ƒ�8�o)��k����N���e���on��r����Fbn�\�Z���g���A~�ClN��/+��r�U�/]�XW+!M��3���Q]��-U�ͨ��:є���k�f�^k*�EXoEs��X�H���芖����9U�������FNqz>��O箜���S��cwu�؎f'{�wщ�B�6Sԗ��ɔŖ�cTR��"U���T�8vX�.�L�V�����N9ϻ~'�������{HATԣ��] ��T��z�t�k,�/NG���X1�D�<2��l��{}���R�5v�4_}׾�y�w����e)�T�ZDG��� �5g�y�������*�lz$�~F�����o�wW���-���F�MYn��;{z�>���ԮcG��n0����^��S�����3��5ڕ-�@��X4�9]��I̳7��J[�dȑ� �]��r�и����#�(�Όƽ�W�2�jo[�r,&��n�c�5ر�35&�֦�P<=;���U #��)A��u:X� (V�7�籥;D_�3�ݙ�0w������z��Q:�=w~2�ޓ�s�y	)ǉ/s�ٓ�ѯ"�PgQ��p��iD�(�c�]e�ꤑ�So�ʴ4ٳ��o=l��893��L}VZ�OTI�gf�����tX�}ÓX�/��`�m�r�XpgK���vf��I�j����ZwO{���t�;��A����|P�%��U���-��5��8;&!}��I�]������L�S�.�xP��x�53X��9o�Q����Vme��o^�6A����B�L�� ��]�t�n;�Q�x���w����
\t�*t���R�2��n�g3���U�]��wZ��Z�	M����2�2d@D���A0̈�Ru��0H�H�)G0�)?��h��u����3g���]DKL���e�U?�r�;�="�TZ�msc�+�u �3�ݽ�������P�Lcw��.����!t{t{��UK\���EE��Y�;Kw�qmS�L�[�Atbk!�J�w��}�>� �kٚ�H�f�uT��=o���Q�y�ݕ��'�ز�y�}�r��;��J����e%��7iM?yLW�E��5��'�%���9�d��A�[;m�
�;y�7�g�7�G��s�+�_o�p�gj��j�!/�UW�dh`��k�l��`���}��k���dm����H��ϒ��]�JZ�c�/��G�vl��Ӹ�ۏO.����`Rb��<��Rrx�حv`�m�y9a%	^E�(�����W��G>��a_}�#:*=��]/-���-��vf�1祃�K�.�O�B�;��΢$Ib	8�E�7]�ߔ2��z��D�4�XS��v�R�'�ϸ)֐�g��2X�|ݭ�^
�������C�!���^���2��+.��:�교�uO�:�����}݀�V�>ś%�:>4����.r������x�=j�
4�FT�aY��?{�������7����l� ̌����{+����9�s�[*ug!�>�h�\�3;�cP�O���MċPk�7-"g�R�"���E����k��ףT����P�݉� �vjS_�71-�B��{��~P�,*�V4��I!��h�vF�͒ޯ<fI�}̹�\�������6)~�6I��A��3.�V���U�n}K+?b����N�����E��+�G�L�J͚y���n�楫�D�|H�2���=�}�@󶁉C!l�Y����u\G���y�Fu���3H�7��9�
�>�d^a�����������Q֣�{�N�����w�S~�!���5�^�V.x�k,�y�3^�w���a��wm�%=���Ά���������ѵ|��Nח�h�Yl��@�祏{����;;�7�jcZᯩ�6�,XX�Mu��:��l˹@���|;���&6,MG���ֹ�!Ӊ�Z�����Ӓw|���/�h�λ����%�*Ku�ed��I��tn]�-���Ѽ����4�C{>��\��V�&�5���t!^1�;�KY�2���)($A"��o;���3��7�G�޽��H��}���i��\w2�cX����Ŝ�ju;���Y�}`A���4�v{s���w��y^���:��}�9���昔�6�o�ޒA!�<����uW�Xx����H�\C�i�~������Cq<�9�ޤ'wٛrt$�>_�vQb4�,x���ε�6'u4p+uT�È�������o���ٷ�t`�fYS�k�o�/��Y�;���v����������[���6�c^Lf.3ڌ1��ޡI`�"=j���qz՜�)��h����y8c�9��Ѳ��_���b��Z��Xޙ3�!h��9� ]dՌ�RGDlz��ŗ�|iݫz&`)�b{�[���SM�7��y�,�	`qY�u��*1��y��{�NCb�a3��E٘~�j��*�h�3��y"|���dP|8����V4�
.� �>��Ԓ�}��г�����Q�@d[Iє�ɻ�Z��0~�ݜ� ��&��˘N���ɶ�7l0q[8wArw��ݓ'��]�5���Z�k��"$�ReF�*��<����
�]�����8�>~�}���H���T�b:�v�Sx�����F=Ix��K�:��$~r���@@WIr����x�4��R:�'�UX�ֆ��Gqj5��vvq�*D\9��d�
�lJ���_���WOК0�ڪ�1r�S6�;$�	�iz}��ُ��l4n�]Z�����X�C�A��ȿ���P�>m����6α����3��>�ci� q�3�L�l�����[��\X�渱���W�Πm��zi����[��cyU{��@Y����q�Ӹ��A�U�C�q~�C��0���^vv��q��(�]g=b܉��۹�7q�D����j�?k�����٤��^7^�vr���1a�s��ovr��1!_�����ō����׍����T����=��7`@nN-=ު�_���<�gl�R�8�)/;�����'*�ese4�_pU]��fk���b)akUj����Q�a���Nu%fgwE]mJ<,I}T2��oT����4��<m�چ&xn3s��ߧ��j����{�e����?�r�M��Mb�N�\�8�Ͷ2�{�Õ]0f8�ֻ 鵮NW��H���(�*�Wc�"�_$,D�a�V�,�EWf��l3S��A-�Okm8�e�̓��O�FF��+{;[��t�Sx�����l�;�t��7�����]�K�eM�η}���qn��Aʸґe]v�e�=��or\��P�a�Vp��VM��B�\�6{]���R�Ku�n}���{����X�Cx(�a�R�ǵr�P�tF��RW�uM�o8�gp_JR��9ʱKI�7���MpU.빓u�_N���][�,Z�ݓU��o�=�ܵ�ÎG�p޶����f��yV)��
r���D8:X�dKe	}#F�3���7+�)�K]
�Z�[]�&����s��w)�]k,f�˅�w]�h�ꖩ�@�(���ǫ8X��w.��&��SWV=���9<�wi1s��T���׳n<�T���=�
T+�*��u�U�Y{i�a��1���Z�Y�(5f�p��X캳^L�*/�Ш����[��! {�ym�bb\���]]m�+3ʱ�ɖ]��q��΅���20�"���˖�	uS�v])�<H����q#+�R,Z�v,��WW|e��2�i4ͧp��V��J��|i�B�#eʜ��YwN-g��V乸�r�qD�m��cwsx' �J^sY|��ՁF��U��N�v�����Bn�G�����KUҝWg����j)p΃���pdjl��w��{띢��坼��K0[��u�5��I�{�[e��oܢ�/�Z�[.�:^n[u��4�^�D�#���;��ܨm�˒���IV��]����Z��%�C�#�C�x��.�K�0r�1�_l��!)�p��4�E�Nz]-}�{v����n����ko��ǚ��{��?��ڛ}�OJk���dϖ��5} ݁��+*U��նodR>}L������'+�l}'Vm�ڬ�Z�f޾q�	+�l��L��A%e8O��|�vE��4�l�C��h�sn��Q�����6�3����������˭���DK`��/tQ@1�3oS����8��յo�ma�����wSJ/-6�u����C44z(ՙ�(E|gx�w������T�ջ0f���ù����w2��t�nukw
CwE���T8o`��;->W�fN�bt�ܮ��h�&�2���\LD����̻&Ӫ�:]zy�S"�^�����a!�S��Z�3�}�=(�l�L��N*�ܾLߌ4Q�D�D��j�<������&4Z%�R0����n;�i
�hJW�QhQ�o�yDAX��	�	7��$*5,��7C�i�"��S1�z4�!���N�Z��*=�˸�yy$����H��FD���(�DTX����mQM�]R�DC-h�6�	���u���������g���	��x�+j�%�U�"��Y9�HicP�ա�Q���==��������q�����������%ŧ�E�0ũE�2
�����1Db��FY�_������}_Y�GI"*�EO-���fR�f��=h*( �ʂ�%�Q�}fN�'f��������}>�fN�v��U�`��`���X�-���g" �D�_tfK������Fjd�{{{{{q��}ftڨ("du��]ڂ1`��eE=nZ�1f4PPReO�іd���������}>'���v{�f�mv��X�����-cl���UMT3ETTPU3C�薃DQ|	u��[*1V(�*�**j*���b�T�PC�^�*�]sƱTQ|ՙ�L���"{l��F0X)Z9��J �c��U"0QUb�"��啂 �fY끽��nY}�N]&6�T��O�3[�ȧ4�[�7n��_TA�J`�ip���Q�.��lwP��6�;�:j��J�	@��Hf1(M�`�F�P�0ѓ5�$�E'R�	D�&*&ϻ�F��zt�0?�����{+��P��o�(�I��"�ٛ��f����Cmmk�^�g�ޜ~��5��t���:ˀ�^ޑ�
�0f|����X�GZz��� �)�$��q�\x��%�1�C���A�i岆�#��7��r�rQ�BґKH;�1���5�e�9>�US�lb�(�
�M5l�T����̘�ee�]�_<@,:���b�*/E�5�@Q�Ε��:����g��jq<���0�@J��o-��5�ةS�IDE�%]�1CtLȹ��l�W}�U^ܳjܶ�U1ܖ6�4�!KS��׮�U���U���]�N1{Z�7_y�W�. �;gM�[^�<IbAf��pct����g۽�O鴦�v`Ib3���&.w"�HǞܼ�4�#S��y�_���w۸˝��x;���С����"��߿ZIG�sU�qE����� �8P����W��.��.�f�3���.g���Z� �s}{)�&Cщxfn��� .�bN�u��/��a�N0;�vH/��r�ŶJ�2��g}׋s����a*J���̤l���[��z~��A��6�,���M��}#��Q��bF���ۓ����A�Z�fb[�#����c��lO.������Y�#e٬�����P\C�֊��I����� �(�R;��I�{��y�~��̯�����H=[?\��@���Ο&sǟ+`
����n�9sB��p�H>�wt5��yj�g���V�^7����T�7g�g
� 	>����]��cr�Ur��`�v�+c�u���g!�����]D�>���Xv�\��-�v�"|�%�vz�UV�ў:#�8k��`c���o_&S^��ԭ��1=|Zv���}�DJ�ס�m��K	!����Y}y�}�	��'���E�R�K�>�$F׺'�Zv��gɷ�	���Iu�z{��aL�3�7�?KP˟D�x��Cz/~�~�1J���$��k5dPnmg���?W��^f�M���'}��)�Mg�lU���q�ɘ4�/�P���<����U���s{X��`��ع��M�7ԯ�겛��|�����0R3����Z�7�ps�����1nr�r��?�i��=�+�D_nW�Gwd�ɗ~)��;.9`c��]Ϫ[�TV�ʪ��ڗ�s�e@����L�u�'ݐs�1M泿m7k�=�[u�e-b�sw`v􁞐y��#���7s�_�W^FͳꉬҶf��ˠo���uUC��N'�fG�on��}�hw*ʆG/:E��1�3��X�X�/nዿ��S�p[��G�d�?/c0Y����أ˹F���7a�2޵�*�@h���fc����?�;�~���o�vgh7�]4�σ&(K� P��z}sݪ.�ݨ�wgX�<�]��EmZ���o��׫�_u��J�|�����w����p2��y�V�vvBs5�y����ޯd�1z���BT���$I#��4[�����8�7.3�Kh�h�|��[y��w{�����>γ�[e����~�~9A�����qmh�[ϒ��`�l)u|�Hv;7�ln`\�;�ocN���@z��)��ב�D��'_������Ƿ~�xv<O�V�*F�*�sN
�6�N�w�2F��.��{4���U�e^!>���^K��@�#�)Z�}���@��@K�]e�A�׏6���y�z`�\>]��Fẙ���[Hi�q�4��uůս���
hq�>�e�՗�E�Y'u�'`�f#�n+UyJ�]Qe~|`i8O]��"eokp'�a���������[���T%E���jR��+�<�D�%S}U�s!r�˘�5Pޮ�>�c���W�k,��j�Ƭ�'*f�D�s䱻��}��b �:���ۃ:��v�V�E�1��5K���Cun �����b9�a�n��95���ꊐ�F�H�^�x��Dl1%���j��=�uQ�@l�x��i�'�p@m����5��3��֎��˭^���:��mCͻ}�E��5��eT��A�!'���h|��#�{sPI��_��i��G�r}����>��3z�Y��X#E�&��#/���Z�7��V!�UW2�	�L���o��d�]Q&�3��8!�f�I@"�����A�g�*c�iw�w>ZR.�o}e����l�<qi���a 2�����v��j�^��{�e��%4��/ٛ ��\�o�����!�܍#a�$\f Q���|����wr�ZG$�(���a|'3c#�6�N*Qu������p�!p뚮�ܭ�K������u�c����)������AM�x�t3ߢn��)���A;�(6{{"gҥ�w���~ƽ�>ԕ�I�ޛ��sL&��;��`�C��ۦ���������s�x�f>�{�u��CV@��\ᅱ���r��"���#�WpCFk�z}�i��@]ؐ-c�n��q�j�u���;��z޹�ͽ]�wOq$ud,�ӛF�a���-k*�8�Q�� ��8tK����8�-bt�`1E�GQ�u[�2������UWbQ^Wg��EY��N��)Mf���z�~\�X�:O��}�Z��Zؒ�ܻn\O��i����>n��z.�Sh�k���(�*�m�=3[��25u �#O�P�$��9��Q�n{S�K{�7��?H�7\n1La�/���۠�c�k�wz���7�𽰝-;-^RO��߈�$}�ϑ|�J�*��:=ף���6�+NאE���Umi=e\��B�C����+�齬D���'r�t�F��N���� 8z�b�!�5Ժ�g���I��QCu����Ϊ�;6����i�����sou�]Ub]���.���i�h������Kϻmx�{gm;�R�sE�D��1n���\z��]~��y
��5�1P$�%�&�@��d���j�q0E�G�
XU��:�F�]�1z{�&|�c�Ṕgm��_&*t��p�a��6�tנ2#z#���$t���a_H����L�5�4^�Fk:�u>��d�; q(}����q��g�`ڹ�SF���:lS��,�7?g(�٨�)�$��|p?��3���	��$�d�������S��r"�o�&+5�9l���M����*�[�ql$�r���o:��Gc�ށ�n�m�8��B������k��`l6�����K}�c4'3�+"&-f���y�fفǏe[��lz�{tk���:7q?C�/�g��Gw�=ܮ_�{�[��DA�[�����s"8k�TdmR�G(��z:����)�5����	���Y�vB���ҎpT��	��o$��i�u8�o0wQqpz;G���m�Y����>x�1,<A�Wp٫_�qO�F��}3���^3�{뵜փ��H�2h�[w�;�����󯺂��A}!s���<��]gF��n�r�d�4��u�j�P���D������n(9��Sw��,f�XW�ç��}wA!�R[�I���*���C���j�=7X��E�6|�k�;�[
;�g���8��	U����-z�=�!��ЋgW�{}|`�鹩��ɞ�*��=.��Q[
s�P�^h��5�����۾yw<D�)�݆8ku<Ϭ8�d���Z! շO�|�R^z���G���X�/�b���7.[��x*/dN0�����}��ƪ�Ğ�ֽ���:ؗ�����W!�0�Qٶ�<F� �*�Kt��1W7�q+̓��@�O�ݸ��q°�ϯ<���]����-�.���,�*����nv`�>�dѽFg�q�'د�������i��[��e{��p�y�-6!1k�(�(�>FJ��������0�s����(�=n��}<f�G�u��J�R6{l�g�-t�*0b��h�龓��fX��_xW�$[��yVڅ�;[��nfi��A�|ͣC���`:���5��׳
�{+�P�8H.��@�׻qt�z7otG{u�w�u��	�� �˙;�DGR�wG��U�<��?���������ž��mx�õ�F���G��A�=�l(���df1#��H¯�������ڸ�}ꇡ� �|*�;�M��JW�|u�����R�;;͚��8�]ꁼ���÷�c<��`�א����t�Z�&dbԝ�%����u�]Ǵ		�3ݼ��^ݒ�kx��o�:��"��*,R���u�4v�J{8�o!G��L���TS�#4
趼b��d�t����ވkQ$�xe�݊�w�5��,�N?�pѝ�k��-�=:6�-�y����^˔�J������m
�cN� ��B�����p�,�^&;���}}��eg
r�����A<�t�Gq�@����;�L�C\��v�t���ȑ$�4�.�*@�/�\׽P!�Y|�v�O[{9��Vn�}�?�^'t{�O:Vb݉�.��H��#�jwj�6�)V���H��)�bL���K�)Q�5I�B<x�U�e_�T����Ts�	\�����	��7����=_���A�k���)T��lK����'+.鷌n�����������6�Ӟn��z�� t�Rj֍�����-��@I�'%;�|_�^����X��2��ղ6�yƳI�Y~�X�p�]>ݱ�5�²Yk8l���9��#U�c��2�_����O�/����C*��c�OyG�Ϟ�#v`�L�f�m����-��1~���ֵ��8�Ր��whu�&�r� �46��J��1)�9Y�����nA������	� N���SѨɼ])ޘ����s���|Z9��������Uۀox�����j#�f�}�#�s7��m�wX;vw���S��r�����XJ]d8\��<����>��ȃ�V��m���{�s��O�� h�q;pkbܷ>w
���b�R�{(��̺͸`}�e>��GV^ˠ<�p���¸���5x�z1���݅���W��5�wh0��ك<�3�3��������#�W�䔷}V���q!�o�-�ڭ�������a��o��� y���SE�@8�|�L��J���C`��AX�Yk�9͜nT�����T&������s�Ӎ��Q'����36op�ݓ.ѫ���'7+1�N �wn�:#}Gi���	�9�o^��{n-O��͜wY��ۡ���Y��ie��C<*����z��^�/L�l���:W�oٶ���Sy�;(]O��i����WV@U@W7���m�z�)�yC������Uy�=5ނ�9D�IJH�ߧ�EE�K���W�sk���q*k�8�<xx�^�3��º3sq� ���utuUǒ���w3�b���m��<j���{	�)�>��+��سb��$�]�<�$6���5�Y������z3���|k����03�Oe��#����>���t�����g����Ģ'4mb;$�8�ݯ�<�}�ː �n�:v��[dp�%[�sr����&��
�rNb�5]JuȲ��5��\T��0�rrb�趪�F�'t6�CՖ_ui\��`j⠝��]�ճH�5m�wR��zZqA��r`��o2��Cv�'o1,J���+]q�o� �}��Nn��ks0���@!f�+n�&������hŽ�}���;��{/�h֛g��+Y|�je�W#�����'d�Qaʣ��Ѩ֑�W$Wa�Էr�ڎ��͘c��GH&����WY�z�u��ħ�0�L��
�d����=�Y&Kv��+Eau�SC�{��ɘe2�&z�vU���kԀ˱�ȇnS����'C�V���{�h���Rٕ�3��p���&�Eq�p�/Ն��8�x�ZO
�h��V%���� ����2�V����8�<�y�pV�Ȍz�_p��QM����.vfF�N}S64�p����C83W��������_Wm=Ӡf.(��o�;��i�ho)��]"o����!��|� �&�5G��ok�8�:������)��դv��T�!
�NYԗ:�X�iՠ,�q}ݖw8TΗ%<�xt�Q0e��e��{y̌+8v�}��D�Q�q��f�J�)B���u�p���2-��A��]���|.�#j>$|�א)�@|Ej~�����8E>�ucAdjSV�b��m�kd4�着σ�N���ضv]7ڦouC$�}�u���-[\�7��������PJ��u[�B���I�͔�"�����Le�f7}�i^�C�9]�Ǭ-���z��
��Y]Q����7n��;���α�q�H�&_^]fh͜�̮�ԹQ�T���\��K��8�v���<�E�t�EbP�9��_s����}`ڵ�!�ulVh2J�5��d�UY�\��b��[�f����ofR��Ns��yI^��h���y&gz�gTw��
��<�l����.�t�hrBʍ�O�h�V�p6��<���b*B��YE&y�]U��K�{�_2�{��A�R����P8����ɼ��ݧ2�MZ��]�ʗW��8��t�>�TDE$�x�M��]��c\�v(ĸ_,�����ܻy���1gCWSȶ'P��W�9�.��`��uu���ˡK��b� �HOc5:���$�W,W;D�f+�j�P�D�{/[o�ڂ)�zv�ǯ�+�"�N�nj�]1��®����9�{Wu�:�PYY�:9y!k]n��Ԁ���־J>c;7S#��������owY��y���#�t�'�:_8t㑐NI���ɔ¬	76�]۹���滞�t��Q��(�E#��gm7J,�EUf6"�.C�����q�������㣯���[�4�"s�SɈ�"��YL��}h�ACT��De���}{{{{{q��_Y�6�d�&�n�b��a����ݣQU��TX�T����d���������������۩8}�W%�U_m�飶�㻆
E��&�KJ�ǩB)=�̜q׷��������gC��o�9$B1F+��-/RQD~h�T�ª��>�%���N�MMMML~�G��gT>V�)()"��2��h;�)DPX�P����O���SSSSS���{>�g��G�T'֕>LJZn�}�!�`�>ɩ��1�dXu��F<�ƱE�PPS�Ңδ���`�Z�h`W�A,Y�VE�"ʗ�D�O=���S���f$��Y�f�3Z������c���|E��7�=���LJF�q�a��4( ��y;RH��=r�~�5�xu��8�P���4��ͣ&��n�/�vڈwbM�X�U�`,_��"<7�m=�1��O�u�·�-��c����L�kt3*3c��3�z�D�jdnjx�����m��Vzw��q��d�G�z2��Ζ�/ӳ��Z$N�{���[�#�{�Q� N�BŰ:| �L=�bUf=Vd���Wu��� K�;�V8���������s��s;U(��7ɦ���/8�h�����Ď\\���,�Q�}>�Y�S��ި��e2!�n9C��^�X"+�����Y�<jn�;<�KQ���S����!�g�m�p�<br�ġ|�U\�z=��}� ��jW��t�{aG����s������0��v7�/��j��&�{�L
�2�>�No����3s����;������RS�q��u���wv-f|U��s����d��-P^Y�X�m d��?�@O��.��~�/�v�[:.y��.�ϳ{!K����W]�J�\���K ���Ӯ���mz�-�O�0.6n��ޢ���>dCU�ͱ0�I�v
�;c���ͺ�X���l�Ej�u�����#�{�!�u_Wu"�{�׹�q�B_�4��O*�O>�4��T�>�k�����H~��vBV�)U����5Y��͂�ד�pe�Ӄ������y�7von�Okk,�^y�����g�V����̳e���0�[V���o4f����5�`��Gf�u�r��ʃUn^�D��V�dՙ>]n��V>1\sbw,	��4�h~*,������[}	�_zi�f�?hd҄O�ѽ�`C�� b���+�8/�'�c��z^=LI'Z/7}SZ���6�C؟k���NoS��������^}��H������}��6�?s}�Ou���^c�z���W�#�|Yz%�5t����~O]n�����tntL^4l�FSM,Ψ�U�q�b��
c��e9�)xڃ\��iT���Y�$�A�H����{��k?��Yf�G���y���s+�,Wj��������]�jn�&����9�Bn࣡����2�G�j���w�aiN�b����Fs�ݷØ�Y��:��Q�,4B�['c�3��rR�q���������}��'Nr����Ж�Ýs+�����[����M۝y��CT�'���a���D�i����,��z�o�T��RT"oO��~���yt�5�m�^�p�}����0��������"�H|t��H���*�sl�<��e��nB�LRa^N�,6�欿5����ש��y�^ϥ���{ L�tM����7f ��X�J�i^�N�]�K�ԿU	��C^ h��'��d��s�yQ:�h��΋ױPЭg^��ȚR��:4L�Mz�?Ox�mH�O���'�s���t1&«���Y)VH���S�w'Ʀ��Cu��"}�16xL�hb��]���w����.^��A'm�>�>�P5w���a"��.�wW���m�l�Kz��c�n���ngr��Ḹ�;y���
�b�+:�ocjK3�O��7{�3�-���c� Vlu���N:��C,�KH�lg�z���Z7�5~�C���cO(Gg�+{n�y�~|?*ϴ�ѳ�բ��]D�K�!]o�F��^TXZ��;>H+����N�&����^bpΚ�6C�؏w[Q枨*0zV�"zs��8^�#��Fz"Sׂ��%�v��k�����"�"$I}��}�:���+ˇ���8{��W���q��������u�e8�,!w��ݷ��m[���r��A���^ei�çgT�o�Q��;�*��6�X�̗�r�͂*E΋���)�F^�}a�I��;[����W��鎚�-�훢�8���#l�j �(�C���� 'FM��gO������60�m͗"#���� t����*�zn�ۉ�X_7��:�wf�����k?z�N�T�g�0�>׭�Kt�DH��ޛ�������rY���W���zC�櫬>�ܑ<�T=����_���E�I���؂8� ��v;m��m�N��h���,v�_���Ċ6�(t'�a��"C���%�S���ҳ�\�ͥ�U*��v��"}FP�w�]�n/�z�9����d�ZL�͟^U.ޏJ1ˢk��@i�� �F��Eĺ�Lw+k$����pW�Rí�3�GV�ZʔY�����v��R�k�}2w-��,Yt�7��7kG�\�5�wY����g��k���w��Ni2�e�C0m�Zf1O4�r��8W{�h�9��ȁ�#�@���9׳�F|>����c�r���7U$�@ꫀ&Q:��j3�)�9RfM����Ux�i�h�"����y�wwn�uW��ڝ�y���y�}�Ҩ%���M�����y����#o�@�F>T��Tue,AJm��rS=�1����5�`��������:7���jq0��e��nۘvb]��K������HU�+��-�����p���g%���va���m�W�UO������)ҵ�c=�S1��� �.{:�0S�N�dA�Զc@���c�U@l]��"�6 ��q�3K�F�38�K�~�Ӱ���Z���דw^��Ն��θ��:��cY��&���te\���T>^$�Lm���W���7p�f1��G5Rv1nm�k�;`�[���d:�g���9�Mz�����EGUkSGoh~��(X�Z�
���������n��WOf��#�`��9g��J�X3��N����mc���J�_n��ڝ�3�Ky��p]OKw7*�&���#����[�� �.�/��= g��k�;�^y_����+���~͝Z�=% ��}֫�6::RY�A�>�11fFw7S��i4�n����m�wr\YI�+8	�"8W��47io�{�O4��	8<��eD��a�ѓ5��ېS@(��z;Y�Ҩ��&�:#�r�����}�c#㩨n�g��|�
��=�=Py���)�,ģ�*&2)����75��@�SO��pA����jr{�/{@�.��uݜX*zq���Jջknǰ�P����TqbqMvߔ�V�#	�B�����ճ��P�woiv��`�>�4���wn�����7�h���ݽ�(,v�U���
�[�B/׍@��cE��/�0���r���I���9�F�H�����x��Ħ��}��y>".��x粵����T� �pBɇ��][W��Yֶ�ʪtZ2��D9�����4�*���S?H���D�*j^��Mx�Y�J.;^�R�R��te:~=�_,�br�0-;�o4�RK/����2���ů�"���,rj�芳�Ӭ�|��Uۨ��1�/�l$-�BT�טDI�$�N�*��ݮ���$Rm%��W��W_y����:"��/������"�I��>o\�/�P6-���ʛ��ۜ���zxw�����ݰm�é@TD{��j�v.�w��Q.Kl�c�.�C�������0���[��i��=>����Qf�kd�6��]�x��wY�o0ތ9@��A>-h���fCH^/+��F��<��m���*����1��#F��r[W�י��s!L$��#[)Ns�(a��κo�+}qE�}�jdY�Be	Qok�SѠ������z*j�y�P*"5GH󷷣�ÞTz�<S���kwa�u\)���{�ʧ`j�z^�$��K!�iᥝq�:��&?����r_����S޼>�s������SL�[�$�y��YȂF����uSM��D������&I���=}ʲ�����
����F��K��s;XN OtG�<rm-1��_r�*h���e��f�%��E�.�);N��оI�Ʋ�<��y+r��+��f�u,{���.{ܚ��!ўx��t�`�O	ݡ+ަG#z�L��mu�ǩ���i̹}��>n�j��X^��]�h����G��#�Ā3j�t�+�n_w{���+s��M�H��x����S�э����A���D�0�}�B����{����}�;!�r��d��s��ڷ'���v�,�+�
uI��%u�D�!����.��i�Z��\	��7��N�W�4�7!|#�G'���kz}5��=w$�e�M�k�x�>�X��H�l2�c����m���k׮]To�އ�\�O��������2X�Pd�.�[[�H�΅�2u������۞좛a�D>#���������G���>3�X�n�� ^��t�i˭��R�>��#�nP|�l���k�^�l���7��3;'�d��[�(
��a8��{��rp7$�w��2Yn�5����p-�C-�y�>��e`U���l���zE� ��κ{���ǲ�k�!�.��s��gm���4Հ1�y��n�������=��|_\�W>�e^�2�oR'
=P��sMԩ��K�9[���*��|�-�¯�x��8J_{��Kȏ#���5��۔��A=�Rs���\�v8; �~s팙��#��$�ר� �ʱ��� ��3��3kך�����=�D&�ǚe�R�����9���O��wTC)��u-�(v���8�pS���ש[v�D;��Y�3�J�]>]wޓ�j�1"���Z}�a���&��^��.��.�ŧm4���]�o���1.ޙ�	*����LϽ�̌N���D��CK�B�ݍӺ`���V=�ݠn93��"o']e�}���q�9 ׀����؜˰��N��\tɽh�ξ���om��m�����xU��`����P���W>d[��k��3�_^Q�B�+ෝTz��5���mv�'����A�z�hG�V�*.n���":gy�x�b���סF�8�U���i�~w���n]v�;�ڋj�џD{����a��K�s7:jG�s)3�U�*�l\e&�R���j��ީ��� �:��rE7�I�>���Ss{��p�5��ü��n�_]A;P����#-�a��� �nnl��u����쮉�D�c��c�"J��z2�c����uʨ�f����ۄ��ؖ�4>&���Pf�fYȨ�ݟFg�=���m�,���z���$�n'����h"B�7�N}��O�����s��U�Cke�`�ֈ�ƅ�������c�^�4/]��$��A}!����?U��~��:7�����s �`�p�nq;�����`f|��N��L�����83�����JK8�2���w�.9��J^r��dk$�!\�é8�ob����R�wuת�k`�}�'Â�N)mc��x�����"&�=Nd�>�9��j ���r����K��|er�|gl�nYV�דީr;��l��g���1�,��$�n��y��\t�׮w���4����> S@�$gV��b����B�]�9ш*��_F:Y�pQt����q�}ϰm��M=�3�`�����._;�sKY,R�=y��Ԃ�d`�����n�� �Qשe�y}X���]cz+�⃰b�]��6�l8'u��<�99�4Z�S�,�D|Xvv��ݼ'v9�O���۲u3�C��@���F"k:�p�_wC��^p.���*�����n�}�.��k�xU�xu�䩨�q�ga��t�w��z9*yViP}��6a�!ѱ�i�R�B���g��q��B�ob��ffI�˫	B9>����gf��Ud��� ����i�;r��$b�a=�L�����x�.��;�Z����َ����Z�,��b;��[|�����s[m�g1s8�ms˹��h��u}�Ws��pDB��E�0V�쵰f�-����)L��Yڛ�]-���6u��lpr��gy<��[��u�cy�ۙoWUM�)q���G�*�ngS�cY,F��]Zeܝtّ�IE
?n�*�r;�˾*Tq�u�b�g��Ӭ�7wSw���uF�.�$��k�2��`�sۉ=�S�of���"�̐��M�ܪu�Z��Sy�A�H��6�8	g{b��[��k(R�[�H�4)%��q}f<3*�;Ҹ�ئ����r�w^��n?2#���鿞8�[�3L=
�� k����TI�˶U��D>�**JI wv1���s���3�dim�La��<�
a jW�����fK�I�ڵ�w�sLp���M���h}�YT� ���,�!M�i�s"�B���}�Y�o�Z�!,��
�V,4�P����$��S/�͢>F��$�y��:��ڽ�R���nƈB+�7E$W`���4tS�wvNmp�ɖ2:���D�4b`�k����V�.s�/�u�^i���v� D8��pm�of��bK<�(mh���H3M�cF�b��i�j���e�X�[���	��_s��,�y�k�A�`�DM���B�]�/�8���G�I7�r�r���V�1+=�bT;�e.��zo7h.�7Pu��Vf���aF�|�Wh{��nϛ��$ə�o7�o�;C$5sE�[Wolj���Ln%�v��f\�5���^1���k@�l�A_h���[*�;&M�G~�G���TÖm�sWKM��A'�Y�|'t�M\;��2�%%r�I�xk�/_)0Z���.����]b♰-׃�����o��5�KUӶڊ�S���UWs���+ss:�*�1�!���׮�6ȭ΅5i#pI����:VE�y>ܷ[Btn��t�9	�=��4��UϷ��z�Z�1F�ݣ'<�F��AY���3׻��N��']r�'7�߲��e��ڇ9�v�0�P�IvuE������뚲4~4�B�/�|�|c��һ6�ڏ`��[ND{����op޸�@Ow�E�!c�=<���;2���#*B[e�2��]��!۵30neذD�QN�D�^�E��������B#R.��^&�F��&]��	�E:�,�-�&�-�6�X�]Y-U"����ȯ:���2�a5����/M�(B!N1
-���Q� P�W:Z2��թ�T4v�C-�[W�_�a�ڍF�$h�DS.�j@�E��@�C���$�m'm�Ȳ(�UAQ��,XE�S�(���,���vjjjjjrr|O��c=�C�PQ� T
����� ()̧��V!6\qNωfM�Ϧ�����''I��1weĞS14�n��w RB	�����1Y�B��_�˟L'�{{{{{~����3�F����Ԩ�=feP���\�w�bEr�b$�N,aֲh���O���oooon����Οw���r��E9j�j�QFA]�11�"�&�N�	fMMϦ�����ӓ��}�g���DU{x�>aZ�wf��B�56�a��(�[�b�N̚��MMMMMN�O���1���%���kN��DgiX��@�6���ET�H�ix��`,U<J�A�m@Ϸ���AkPX��U�/�-A@Qߙ��%���m�C-*��Q'�Q@Q�DĘ��ʕ��,bj,F)<H[j� \[U���Dm�Hk,�H��PX���U@UP ��t�62S��`Ba6��t���� w:�O:�Z��w9�-���lWgÂ�Q�9���}ne��T�ݓ�v�y�aյíX�դ��k�.�%"��7T�	"�T�pŬך�7�殟-v?IP�%��a����m�M�P��7<���O{o�\�c��j^��A| �x�Ѷ���b���F�5M`��G�õ��cw�'��z�a�q����s��y����Ջ9�-��hNѠ�KL����wv�b����{���,p���z�Q�׼�bB�d��fi��sb-uMb�P�nہ�&v�CѮv���'��0w�����l
��.��^kOwʤ3�0;�i���d���}}��oY;Wr��x��:��"��u�/�WJ�Ʃ���گuJ�<�Q��Nּ��h�����a��T�y�۽B9I�#w;k��smf���Gz��3�ML/ۦ�L���oS}^���?����iP�[3E��OB��H�"���0�,%s��c6Fr}�*4Zp����*��[�uȬ�3�$	U9~W Z2�����W�r��÷N��W-���[4J�W����΃���<��2�Ff���u-��J��W�E;M�d��d��GZK<����ڰ�H����T��1�|���iγPW	nw �v���ŝ�M759df��l�;c ��yN���=@� H�#����*�xw;�"��4��_7����9�����QL^���;J*�U�x��TZ��C����^7����߳�������_	2�Ѽf_�Qڕ+�7��8���򎷌ʷ�rA�T��hv�Ӳ��	���ݼ��� �j=��'e@U]�%�"�	�2I8��7�����͊:34r�0!��/$�ܞ���T���j���듁9�j٦�g[c��V��H�������bA�o�9���ۘ�x2��Y
Ю�n��p����������I ���Ƈ��;�zw6=�}�����|�;ޙ�Wu7�9��l�jHp����ނ2�N��(����[(D6�ɌQ\Rݍ��\-G�G��N�H���>�@��㋮���'�}���d$��70�����P�� ���(���O���B��s���/BQ}/��"��=���0[T��7D�&j��O�({z�q�ş{�GK�%g���>��]�']� >�W��.�s�v�N�����oj`��:���Z�ܴ�/��c�NA4N��8:.G�k�}�=��ן��%BP�5G�>�ݫQ��ܽ�6�j��l6�W�H����/߅Y�+`�O����j�w���H�c}�߲X�������}��b��(+�\�͚�k���w��X�<v�;�fx�q����4{C�O�xn6u��־gb�x���f�y�����u>�Fi��쌘��.>�W~�����N.�9.X1i�gti.�t�m�܅F�}Q������Y�����6����c�e�Nj@@[��A�N�3
�z6<��b�w����3���,���co���Uݙ~�ζ����3���(`�j�w
���婻�hI�)�j](��JqG�>��Ay�1m�ۓ^�W+�劊�}�<�#���V-�su��k1�:�"!���Y�[��!��aԱ��ptS�E�ws{F,�f��3<��O|�&�U���;되(1v�ܧ�za����A�۫4;2�|�ً�x�s3eA}O�UqC�Iv�����|k/��d�f���-�7���q�c_(�J���˼��jQk�˩�OĹ{��%�� x� >���3��rܾ���܌�����-������U熈�ț5���lf��G'��ײ��ȍc���o^��s����lu�ŷ�.����9��.r� �w��( >^�����Q7��{��~�K��?
[��]iKQ�z��)�sz��ޏ	Q>�/y$�'?����r�^1YR�?�� ��3�J���x?q�M��4;��e��k�_����m�S;��-U��Ä7�������zGd���-���1�w�U7߻��S]�*B���/���ju��������|m���]m�b�]U���Ys��b{юzq�K[�����j��zb��A��^�F�Nyu�`����*�"�F�E�Ϧ��N�Ú�73l���5c��Јw�uͿei�S�M��0c�z�y�f�拭���M�nYnʯϣx��{�`� ��2���c��uZb9(m�X������,VR��r��<����7�_@Wق�ۍ�V(Y}����J-�[�tPQl�X�.�_J��W#�����{M�c
��d͈aC15�YD2�hEƿ;m"J��FĹ�����>ﻝ'�l�6	e�6���egk�~���P�W�A���D���,�}; ��W�z�	�ˋb:�1�<u{�����Ki6+��O>�
w�/	�-n�[k�Gr�.&��d>��3>14����)F�9F�o~��͡[9�l�O���"�8(ToT����fF�7��Uwn7�Ԡl+�����+a�mC�n��f��,d�LWkz��K76L���� V���c{�۴��l�bpL��]D�E�j7-�,���E�<��G�� N�7�������\&�I�j�M;h�3��1���=�;uJ/�DNv�;n��Z6h%$�������wW^6���a�VSI:�=}n-����|^Iv��{�9sPu�9܇��evu0�s���H^8-�0���t��E$���%D�lș�=3���@ǈ7^s�=�0��'��F��}�I�ۚ�8���z��S�s�g���D|��lS�wE/��!]8��%�֕�v�=�����5��}t~�pr���P6�kh�T�u�)�=�K�/7���f�U�Ucx��<H�#�"<E��fhB^g�ۛ��]�_�1�.�����e9��s�7PMJf�!fs�"�$¡TOo���:_�<�v�$��֩����i_������^k ΖȮa2oNs�b}�9 �`%�|!����sZ�V�kU�~�$��L��3��|R�;�c���>�vô{�*q���vy+�@jb�C��5�!���:��:0�߷�TP���s�̴��đ&�'i̈�[8��L�og��@~!�+TT�'���u�_�,p��|��*�%��f ���&�@��4{#�["\6��h{��ט3��U��P-�;�} duL���v:ª��������s����W��V+�����Ml�^1������t�!ӵr�<�Q���mv����(�U�m����
1⡘:|���i[M�kٽݸ����>p��115D�i>9u�[^��I�l��T;G�dR���;W�fXR����o{66��꽸3F�ކ����ӻ��]5F��n��r�]�ϭ��l���"�-۰CC���N����$s��H�� y�b<�x���2�&���b`���1�wʹ�	���#��3������9Y���B���t�h� Pc"�>c�v��*׻�w�bOKnd;�s�u��Mlϖ.����7b/8!�͐	�@ԩ��޶v~�[�r*�_,�p�T����}X�A��A��xŀ����;��c"_�~X�us�ݹτ���-[A���K�ʤhZ���]j���t�mhWpD@���w��{g��F� ٩�;\P�y���8(��U���v���Í:��cƫ�ðal�cW��,�k��)��iݨ����UwsF)_Up����:�@��όf�7G�b*��
�i�?��;�4ݼd���޴ՍE*���v�3C��l�=�d�]�3%�L�erB���B!MD݇��IF������N,����<�l>xy^�҃g[�z�tr��
���]av�?Z���чS;V1���x���\V��gI��jcUN����-����K�7ed�</�I��fM��>�햘�0�ޱ15�C0�뫜�JǷ�t�iw���<����Z�G5��HA�R)��)�#l�V,���c<Ǥ��#JJU�Uw�������n��YԮ�������e]q�K�֪��ށ*:<��<�M:�Dl�ƴ�N a#���v��I��.�E�oXiMzp0�`�.-�su��������5��^���s|3�^5� �A�;��pS�\X��j\UwF,��ϱ6Z�2�?�����m
�R[�M���ؐ͠��َok��1�@��{�4��eFP�Rٵ��/]���1�M�u`�:l�Gz9���Xa뱙+5[u1;7��(O7���Vf��Y��}$v���������`�����8C�
v��;������|5�}�t3�ʔ���w}��wBh�ܳ�Zfr��h���P6���=mD/Q�����g#+6���{��X��Q��������b�Ǔ������V�_KeW�<uG���,�Ov~�9�ڃR��c/�v�0���57b�ݢK�Smf�.Rq*.X����]�z�߱}��_X^Q��AhLA��r^�d-�r�"�`���͵#�a�^J�p�3�%��YZKY1�!�A�Ҹ�M;I�::G�P��[�<��U��V�K��� m"W�TD���]$i��F6ǣ@�T%R��ޣ�]:t6�sU�J�H��C=SV�biD-ٹ�\�wl��ymyG����{��f���'+e���طz��M�;Nza�eLj�w�i�ೲ���tz0ZM׬��Z��ٝ�=m��k�pI��Az����e���:`�-�A�C�+�j�Ƽ��7�٪_6�?@�,���i�{T�V�wd��R��8%�5�3C��'�����0�׵E��bV3�l=k�������2��kXDR����/,�N���.`"���[��x��U���]�H��,ʡ۱�{�� /W��� ��D�~� u`y�C�ʜ�ònFk^k
��Gp[��G?LI7�x��0|Ӝ�藋G�뼳���}�~ܿ�	�:X�<��I.��Ի�4e[���z�J����Ӥl�gXۇjC;چW\�+RN\����6�O��G/u����Y�>���Y��X�Y����~�2�L|�2���]ȣϴl}��l�ƥ���h�?*�U��d�r��IX��5C�r��=�j,�=S���fE����dϖf�p*v����]Y3i�t.�}�5A �v������ͩ�U���J��<H�YUI�[YGJ�7]�BlyN#�/{=��UgH��A���*�>��W��Tl���+�>�ʂ ��w����N-t�gBv
^[��S?0�x�[�S�O�<�aO��[����{f眆 e@�ެ�O4�Mf9���U��e�uvP��n�{]�x����,#gro���wMKD��w#'B�w�=��m���V��퐝�aM~��~��F�����ѝ<چ�_
�8�D�a�z'^Ȇ�8ޞ�Q�U8ϵ��s=�R������d>�}��yU�&�hk�����R��9���li;YX��i�C�2�́13o���`��Z���*@b<�TҾ�l�<��GX�SSQ;#I�O�,u����^�w�����°��^�w[מ�f��љ�ץ��<@��۵�t!����$a��Ĺ.�~����Cs�wz�wozr��i���`(����G�������O �z5�_[�p��^3yOO`#�z����7mu]�8x�hng�`�8w5YtxY5%^"�CSW��׀��P�3ڽԴZ��A�>����T������X������wO�q
�Ud;�rP��ucיm�p3��0��&�}��|{%�:�U��WuwOaY��Bf�]$������֤줦���DZ��w��]R�韒W�{1g1�"�E@e�t�"(S�����˵��m���o�N�Y�s\Jʆ��x�V���'��t{U��O�ޙxm��'PKmZ�(n��o�v���W]cLU�+��a�e��T�P ���R �#Vb�ȺӑD����vF��ws(i�j�K��\�Mt����uKo�t��!&:Rg� �c�&4UX�G8f���+cDÜ��K���7{9�̶�3���6�$�XBW
���ʳ��V<��+뵘�]�x6������ܬ�}�5�ڸ�<­�c��_n�:M/E�Xwlim�A
kdx���	�s)X`_tƦܾ��� @(����9�A&c½N�ko��+fr�]B(�Qڪ�Jn�0�4�T��N��`@E+k�������w�2�ʳe�y-��q���p�*���g`�Ovy����V��\ƕr_s�(^7޼a��Ժڙ�R���_U�,b�qw.�|XQT`�PA��uN����3q�¬�ho��n��Sr����s��S5=�
k�>��`�>gD�f񙫸�_dG�����A¬�w����WX�"S�w���R��^�T���0�3*ܻ2�|�b/6�=(sV�c�1��A3X�C<�8�Y:��Gzsʝ��*���}�卹��:`�d�R���W܌��D�񩲧#��X��緤��3���J(�;o'<ɤ���O�.�A�G�r&��]s�s���A�¤]�+�`��]�1X0���i���sb��\6�Mԥ�u�����,�:<��K�������#d��Һ�Q�VW_���N�����1�:<��I���=
9�7~{�%^ui]�p<�W�c��{�`�!�m[	�	ŵ�0ѐL.�vT�W3B����\+KY�ܦf�,�{���������m��*jQ��l[}�+��b�;j�$�)VB���tN<��l�Is��d)aYg{%��[����L볚�{�*��~skq�mR}]����P�q!�e�ft��f;�����&&�}��k�E7Kޮ��n>�ݷs���{59�����\��Mc�sdkpX6�U�Y��ej�ޱ�J��*)*Uıa�TȢ�w<��w����h�$27�5W\��C��ۮ��������gG�@��C�1U ���gΘ,F"F�*TP*b� V|�<zq������_���}u�׽ǩ��q��b�AE�A$�i1��R,�I줳&���SSSSS���e���=�+�R}�ꤠ�4����Jk`�Z"��E�	fM�g�SSSOn��x���݆�~�r�M/s�u����^@R�Һ��_|{{{{}}g��G�P���:N�R
E��P������S�%a�.��/f��ɹ���������?^:>�i)�(y1���b¡U/�a
�Ҥ��Q��d�yLv�s�Y1��C-�"��z�dQa1�o'Y�P�!X���*"���M2G-d��Ш�g�LB(*�H�T1�0LAT��VCF4���ƾ2��4�$B2%׻��x�n�qa�<Ý�yp�넉E#p꺋�f�k��"�p.��dyo-Z����e�O��ƽ+teY�����{���2�S?��d�2H �WIqr׹yՇSԍ��V?�Ջ�	����v���1AX�d�7�&�������l;i�W�E����ˈ�k�ck��ltܤ��ڹ}�!q��oC�%Q��Yy�>6
������|=�B߯�Hn��mfsg��Z�g��R�۠^[Ļ�;@�"?0׀�7 ���ko0�k'�ĩf͐2;��2���J������箋���g������ዶ�l�G�b�}r���[!Z������Gn���K�_�z�C��ns���u����{skl��M�,��1X��`K,5c�|�f�������,�i�>������~1T�##�����������)�˨Rg&�YG4<�!��CLźX���l��>w#z}�IH�a�CrFo��z�_f����|i)�j�c��H׍�~��`qa��Z��4�2�뼁׬q��;�����:0�X��f��ܺZ>�%�5�iz�XZ�~�N�����j��~����M�j����I]���+E�����oZ,����t��k��"�~���0� x�>��98�\:���P��M�˒�� Ny�z�D/5�ہ۠�§J趟d��uuF�zXg�!/޸���4�m���jܹ�vq��(Ԡ��>�P2ˀe�R͍�V3���)�vJd?[Wi;�~j�<}y=/��E� ��*Η˸�-���t-
6{��ǁ[-{<������6��I�T��EY��{��*��z���T!'<�V��ӈg~����(	T�H�j�����2�v�l/�7%��
�p:��F��0��n�g@ʧ�ݼ�;�硰z.a����o,L��l�Ro�R	����8$L�s��T�P��g,�Olʝ$׸�_5?Gnݑ�7b�Ù�D{} ���z7yo���󵙦.����k��a��d��,���G)�gn��u	b4Ү/f��'��k��X4�Y�ъ�6��6ݥ9��g����>�d~#x�zfVʠ~��~zrk2F��m������R�eݺ�j��NT��bW��(u���ͼF�_L騶)
��Z�Ą�,v�9��?��)b� �C��\�Щa�&�R��v��j����fg
R$Fذ�*��v�0���6xs؞Gd��5�cm�B��8�l�J��)@J�A�x���`<	2a+��2ؠ������);ޯj��Aꑳ}L_T��03 n�a�2DtC�w1��N�'�fY��3�ǯ��V~;��mV���,N��ç�+��{;ɦ�x�-m��������[�W-�t����m2��0L��جoM,qw�2]�x+�z�<�W�ձ}�ri�'LfA��43_�Z�C���K�sRF�|�fT���0U��g���Cg�iQ�^:�,o 6�C�v�=z�2��kt�?~�J�:F,
���o�%$0�v��i���z6�`�큛�������]��V�fns4�^�p� �^��Я�z��%����E�oj8��~��L�e���k�10�MJ��/R�f�YQqGqg���ї�@/j����j�����1��q��f�cH�U{4a=��/
xu:c+Atv���}��z�8y�-<�C�W��Ǜ�����hwL��e��x�s�޿f��HR����y�+M��(��ǆ��oU���Ʈ]�a�m�y�R�h�d�����lL�%m��j�p�O� x�<t[M�N��ژۋ�Uк�h�Xl�)�0<ט�-���^����Ջ�u�u�Uǳ��S�oO�s�΋2M��j�$F��e�JU��{;ݬ.���������w*��H~��!b�^�X/�Z��\�Wn�H��A{����v=���i�{O+;v�RX[�cv�[g"��s's��棏�쑺�4�Z��!CӼ+����L�$���y�y7�9q�j��t�������"5�G��G���L����k_h�NЩ%�&�9�8v�/��۹\�Lz���=1	&�Xo��6Ey�V%�>�����,F[ץ;&Si'����o�H��q�2�S�y�Z��O�G�]�{�T37�}G{ל���?n�s�S�������r�ܥ��-����H*�gO�S���n�s�K1f`:=�G\�QӒY<9SpNĊ����5�_��Nr*�m=��Wo���|�E��wf~�f�רye��oz��K���1��y�|Q'��6Q'�x�0׌]�oC܀��9i�/[�a�r��ۗ���)�ձ�4g<'.�:;��-����&��2<H$2�ֶX��Y�6}��� �ٱ܃+�į9gI��Gk��9�&Ȼ�Sa���[�3؞��\D��TUt������)v{B&*�l���ԪXzm��;�?������>(x��L���^p�*�u��6�t�N�{jUoW��w�Z�����.��[�Q�;3(�\3ֽ
H�4�@vxX����Q��'{D�]-����/*�f��z��3�ؓ� �0CA�[�.U��WVu�_!Y<|��ꆀ��w-r��^E�E�[�k ����w3{2'�lwu����]%���*���A|��0bWxɡ���i����0�2w�(�v�~�o��ޓ�ty#9{�ĭL�	���,�kӒu�����\.�զb�Y�x
��Y�{�z����<ژQ$�����ݬs��S`k/c�_�"�����i�D�c������6�ɩ z���-d��o�5gS��i��j�q]�ϻ��1+G�:���C>����̛�Bv��..ݕ-�϶���f@�{pHq�똜�}Ü�S�A\���2p3a�.�;��Ww��#����l�)�I�Ж�����7�j���jx��X3p�g>)��(�p �N�� wX���1��:/�zx��m׾���Z��O�]���t��6ګ�z�a~�j�Z���y�s��[`C�O��V�u�n�E�{�Z�w`^�s-�G&�+�NZ!�g�2��;]G����E΅b��g%��3�C_a<�Q�9���=q{�.�L�?��م���Q��Y�5����m�pvCe�\�{�gc̻��#=K�tذ��M���n�7�d�P� ;n4�svk� ޝʪ|.]�g���@��U��{������۞��~�a|n���Sq�-S2�z|;����V��Ļ.�J͆���v�WS~O��*�R���|�w]̊�n����E���,N�9�uvmǻ��&ӌc�z���ooD���}�p�nP|�����,�v�����D>0"�"�(͸��/���N��xE��o6��P�e�fs%���\F2�Y�(�p�U�n�|8���"��a�ʸ�����/�b�yNӔ������[*����!%Pa��2�vza+�@�k����(�������R��AU&�
J�Զ}Q��x��	$z��S��W�p14MU��+��<��5T5��qPFX���'��B�#bq���Vc���UV߹+VR�v�<h���S�M2[��`�~�o[5fr�=�N�Ἑ�{�R�l.�ܽ�=ݗ/ŷ# `�N֕f�!-�wș����`�<�[.&�[�m����G�sF����&S�1,E[]��,aZ��^J����3_�!�c�U�q��nռfon�2/k�Џ �<.�w�2a��+��x��4-�7�����ެ�P���캀v�����lz�8<\V�ǡ�l-��ڌ���Kh�B� �}V�L�6�.������^�׮�q�ݶ�k�m��y��צ�w0 ��6"*$4P3��O����{}� �@�#�}x��.��baF�X���|*7�ww7�u����/��XKMk���?�k��e���v�%��B ���JИMAM��r���{�69o�j԰��_2k�J�)���+�Y5_�'^e�r:��u�k�?=�r�z�y��(�}|Q�8����{���M����r�:�ؤc���E�/u�5���� �����L=�I��]�t�R?~��/C>�7a�:�αu��ꜚ��oP1�R]�y��y:;ͭ�5W�&��G��m�h�TU��ɇ�-^�-��cˌ?�%����3�b����P.�\�4!���j|���~6Fy���n�؅�@S �G�H���ud�6s�#��u�U{�f��ڢ�P	U/uo,��ۄ��I����}�!�$j�Pʤ).�3�21*驷ӯ��R���oc9��'��[Lf{�i{�!���X3�19å���n���6�ug{�;�f��2ݛΝ��Cӝw�1��M����ծ��sr����Y�7��˥�޹0�]��j�c���&�9�
���cs����<�y��W��5��ʷ5STO�yy|�,���3��"�����=�" ��I�}���^�*�����F�-<�˩r�=�2a��yƧ'��6��V���Ѫ�LT7�P{�kמ���׾/��t����_p�f�浉Z���.��oW
-}n5DT*4�+)l[l�Ȣ�浤�s�.�=�qN#����Ok��說�[<���_j�c/r�&��q�yIb��xn��<� � G���Y��Fh����D>�@�ȷ8�;K`d�`Gz���ڢ�0�&���klej]ܗT���gF���*P���c�P"�Ɠ2�D<	���g�	��m��3�˓�HI'�Ct|�������HmC��k��ݙ�۞n��]!��h?��W�Oګ�}R�~��Y�ȷ՜li�w��(�$�Q^��߃�l���a�q/Yɓ^z[�&�j|f7��c
�_^�x�R�Qb�����o@�
��7c��#my�O3��}���^��<��0YkX�p��N1O����6z�ʹ5�̾{XM2R9���cg��~�;)�������y�*7�OsV�[��Uuo�� �f�`F�/����w�����ƃdcV��z��y�쩭��{��H2��Xh�_��%ط6���g���~	��z��NȻ���&b�ۗ���}��˙���2�to�7�tNJ�G/�L��cFr�V���-۩ �uQ�wuNԖ�i֒淈���-�����W���'R.�k
ʚϬp<��u������G��ď14򩵫�Kz=Ն�p� ��������7#�;��
E��ԩܵiÝ���B�xS��N�߰��������u�9{gʈn��S*�b-=���Q[�����}	üU�>jp�������[G��P��v��{����??�"�=m�剟O�3��/��S҆UՐ7��k3���]��e��/�������">��S�x�(kSv)�<Ք�D�x�B�v�ɧ��^�U�~Y�Rx���f��P�E��R��K{�Ta��[�>�\��k�6r��v�fs��h��a
�?�,��.y���z�@l٥!�Ȫ�{�G����e��Xh�8y��&�����V�Ц�;����sv�Y9y��[��aAM�Ǿ]�΂��}�+�o����W���O���ʗ���U���EO���Ӏ ���UN.���DL�Nt8y��� ��@��@�"�����"´2+��B�8(�Q�!�XBa	��P BQ B BD 8�O	B$U� BUP����C�H� BP;�8H��!����*�@�0!  �� ��C��!*@���"�@"!�@����B�!��"p$T�P B@�	U$� BA@�%D� �P B@�	DX�����#��������������q8�������*@����(°�H�! 0!
�u�t �������� ������������@�*s�!�R! �	Q�	D�A���A�(BD�8��>A�/���TB�D	�@�HÀ2��~�_���/���?�����������{��� g����Ns��;�s����AW���_�O�A�� "
��O���@��?�_�O����� �*���C��O�{zHy�W�'��/��	��9�?� ��
���UA�T)�
E��E��ZTX��V�X��E�Q`�FYAd�Z)F�bh!FH� X�e�bAfQ� "Ta�b�Fd$eZ�E�X%$X Z��bE�FYdZQ�FE�V�iVFQ�Q�FU�	F� (`YdX�fE� Y�a�bE��e�a�d�dIVeY!X%���E��	VE�XXIIFH@$XdX%X XaY%V���d�a�a�eBE�  % X	H�d$Y	FXIYVXT Y`X$X	FI$XaX	E�F��aRQ�E�VR��E� �I	%Ye Y�	%�hH� X Y�`Q�X�f��Qi�iA�fU�� V�b� �X�ZhV�YQP��Z  �X�D�hAR��T
�  Uy  Ċ�#ï�.��?���DEJE
 P(�G@�����������ðt�|�<�^���?_ۯ�?�O���8�����束�� ]��O�ׯ�>H���� �*�b����� ����$DAW ����4��hx=��p?�����'װ���U�?����� �*�a�(��@����ÿ��������'�~���x��*����������~��aI�/��8~�\����?O��=����$��x �*��I����?�v��A�_����}_�@A����؀����]�<���?T���d�Mg����f�A@��̟\��{�/H���E���PI	R����P��P����*�!BR%
��JJ�*�ER��$�E%�)$%Q%R�B�RA(� �R
D*��� ����(R�$��UBEIPJ%	%@*%�HURR����	ITU
��R"JJ !P�R�@��E*DUEH	UP)TP�TBD�P��J�*(J���@�J��J�$�a�  �$�SF�V�3[V��-��m��E�Ef�B�F��m�#%5�/\.�k3MV�m�١e����UkZV�U5�L�٘�*�**�JIUUO  ���СB��hQ!��E
(P�B��8t*�[MRY�iU�SeI�Fիֲ�U�dV�KZ�!�2�MmJ��i�f��U�EV�T�,�B�
�Q*��
�  Z]L�5�l�3*FŴֲ[,U4ha�D��dh	�(Ԧ�)��5iD�ئ��J�ڭ�٦��RP#*H�(U	
� *�G  ��H�Z��k���5�U���جeT��4�b�LeXԪ�U٦�4�L��	M�֡�T�%"�%(*�G   ��ulI�6-V�k��VJ�vv�����a����iT"��M�fU!�`�]�e��UR��1l�*�ݤR�T$�J�-iU/  gQH�4���o\9YT�.�w"UKX��n�Z��%;�s����D����X uZ�;�B��������9ª*��$UU"D�   ��ҕ-����P;��;5)T7
Ϊ
��:�p*��m�ݳN� �9�T�ۻlӎ0��+�u�]�W:[��J����U$���  p����u9Β����6iQ�.� n��l��F�t�9*��Mʰ�ITuT�ցCv����4��`tZU8�I"�R���(x  ^=U ۵N�*��E�.4.�UQ�4WCF���K��H�7@*J�\����[vH���@��7)n"]e��F�J*�UT��IT�  a碥 /:���v�:*c�AWps��PuV�R�DkwQâ�(÷ ��΀)1����[q3� I� �~@e)J@ �)�IIJ�� 1�L&��	�)� ��54  ��M��C@  BJD2��  =5?#��?O�_�I��&/����J��Т��"ϧv��(�4K?l*;˃⁖�v��_U}�Ԋ��^���_B��*���+��DW�(*"�� 
����Q�����Yr���k8�� hPh�Gr*ݷey�70T��O��j��tj��L���On8��Eն��y)�lR����wu� l �i��H��˽�Cvὦ�JD�m���ְ��-�`nՉ[��1��,nZc���=t6b·v�0�V!�^�ke���`�͚e�� 7s)�׍1;��3��f`���^E3Wrཙ�khۙ���Ʈ�m���MuS�F�E�/h�R�B�n)�#(!�T,���]�*I�W@]:���l1�lZ�i@���g(bm�hch�:�,µ�ۺM<mTk2�y�:R�I���H�4�����a`�I��Yo���m�"�hu���T*+�k:����Dq�F�ѕ�v]z�2�dT;GY{6�h+��OF����E�5g�yV�C�� ��wYw@kSL*JQ��A`]���ĕ��K*a.�F�#��@��9���G5֭��- �P�3:�%���ᔦ��R`�ՎCr�@I#9yS)^�+	J�
7XѦ�]% 7%���{/k���;-�I�r8��!D���d&���Kl\ۧ���j�Xٺ�%�%�	d��r��딆�!��:�K6�&� n��z��k�%�S@�Q�q����B�Ԙ��M���5kA�H�2��%s�Z���� :�%��%5����k�-�)TgiR� ��,��P9��Z��Xݠ�m-w6�A�.�Cѱ&A[�Q�Wj`^����f��.Lʓ4��)P�Me��#)�YA��/6��9u �V�E%Z�I�:��#oz���5�e�R�3ST.�L�5L@iQ�1���WeU�YJ����Uz1�MM�ȩBx$Բ�)��T 1a�V�hoeS�6�&��
N��xӒ�9C-���m�u{f��O�i��9"�\vw74){��0�t5@d�RIJBԡG���KF�âVܫ�-��wY�|�w�^Q�3:[������Y�2�i�.���ӻ�S]��,D�B΢�kq�7x��D��h=W�P�WK.���#�qX����7qK��HJ���[�-H0˛s �q���.�?��/K �ڙ����R�Gt�N��^Lո
h�%�
�v]�����!��P:�bҥW��7�*�ll��4سB�S��l�3i$s(�͢+h�EhF;M\��r��pަ�7�j�R&���n�Nڃ�L��n�%���z��L�f8+h3X*	F^�a��i��;��!��Y{���`+7��ِ�T�h�iȦS��X<���Z2�7*c�Pv#Nm�*��坟c�b��]n��H�,ϥl�sn����m&���)4�fa�,�Ǜp*�a�LѻL���ۀ��Y`���#��X���˂�MkULz�B�F��N�S�^�4�Ʀ�8,����nPh��u�v(�!��{��ۈT�$����--��%��l�ٴXb�R�l�A25y�����X%��B��J�kF#��jZr�{Oc������N�ˬ���p�$&�z�ۙ��Yt��acEj�Y;YyOb���t�'BL�R,Km��2�xn6�@�{s&�yS+h��rXەw[o0�vm&�2E�:jt�f'k[�{��x�.�c0ͼ%�3U��n��13[*��q|�ec�mn:F�]�
�R�M�x3��e	N�Ǒ�̂�K E�8����A��A���hJ6U�kX<� 
')2�zH(��E q��IH�Dۢ�jRеn�eZ�%�Hc8��R��-�(|��5o@�#�ܔ�+1*�dJ�-P؆�f�)l�r7q2#BU���Q<:�FU��L4ʭF�+մFS���"ڎ�;l�;�\u�r�+1Q��&����I��D�����0,?!V^�i�,�n-Aી�)M��^n��uj��A��Q��VKFR���x��]��2�U�4�M�fneن�'Jܳ$�ԪM�X�T����ԓ�8^$^�oo۴���J�ܻ[-mmè��A�)5h%@Q��(-��mn�U��&�!��-�9H��ׂ�T)��#)������v�^�~2L�E�3L��/r�ȑط�AN+9��ʼi]�1xźe���-յ��cf-��
�Ķ*���j苁ܬ=�1)�H�B���[&�� �|,HƭلD��#���e�+.�&��ÖiV+FJ2֒��c$)�P�
�[��6��SeiƝ�V!��Q�Oo*L�*B-}�YGsY��U�u6f�h���ة����me�t�\�u7k)K�����̖��m�ܙGNi�� �-�%*�GA;���h��+#!�<Ug�'�P	����Me�QT�-��hz�V^k6 {P�7��D�eaFnL�z�cV˘ʒnB��`|�Z�����k9|���en�	bSDc-#xb��Վ�������;��J���Ib�DM㙗�sr��=��JMMu��٨�h�[�b�;�h]f�X�5t	�L�w�Y�SN��5\�i�փk1A�������yw%�u�:��Z��z����r�(I�!"�����{+Jo"��T�Mh�!(-�-KX"�V��Fcp<�Ֆ����
k���o72m�%*��9L�ʹ+�7p�Ė�/l�0�q9�Mᣍ�iiʆ��N<���SF��C��N��ILV�0�{I�����I�=*X�5���5j�F(ssMc�qcJ��uI]�1�QYr���a�IFh�{�w�I���)��`M᳑�e�-�Z-[ �������\l��q,BM�2��R�٢�����`ݪ������4��;��U��0�m��ԁ���h�Y]_j��mk;���f��%�[�i��/��8�Y�_`xe)�n�Y{�X.������am�Xݍ�۫�g� �"FS��Q���Z��t7Vmӊ�R�:Y��B0l���6�����Zj�1��R��f�S.彐��!N#p�'pk���y�(��g�b��ul�Ҍ]���4��nA��6PMM4*����ۭW%�+ۉ&�Q	a����|��cf&Z���dm�`��)ܤb���Bֆ�v޽Z�6�&s�Q�iT��-���
�(spQX6�2#m��<�t���"ŘAҊ�����zk!��NU�0m�׉��jƻ��$�1ѠvC46�bz.(��.��;�e�۽�F�sp�Q�T)�8b�CDH:
�d5pєE��R[9$��i�F��$Չ��&�Ȉ�j��Y�u���y�&\.��R�(q��{iÖA�(,���B2��b����A�M�-��-�D&w+A�D�ˑ����Jwc�ڄյ�>VS���+h�*b�I=pѯ.ޚ��I�֎9�-)P�$oٮ������ٔ��,S1i.�ZяF1t�k4�`<B���H�A�%�)cWc�Ce�ek�Qm��1*٢ ����^Rv�e��ŕ�����"�ͭ:n�`k�E��H�)�ic[8�����FH���V�:tб���M�B�˔��f&�=gT��U�L���٭���[Gnc�Pdq<�ڵxU�:r:�-�4GN���}s
s44�vJ��H���Ȟ�
^#��uf�z�7U[S3c��UbԤ1�v6�˗�d9��L
8��u{k헫�WOe).+�S7F��Mj
��.�`3�٣S�4lf	�/m��MY�TN�9LSZov����Xk���q������N��S�@7�h <:R���r#A�A�t�d�Rjm2򣎭�����Mt�֋����\����v��)�Fi��π�Ee#j��G��Ś�e�h�ٗ	@hB���Zn�B]��+W���I�e�F� dq��J<��kq7�8r�VҬ�ԖH� U�)�h@楗B'y������hby�WcXҙ�nD-�֢�l�j�Ө�����A�J�+#�z�~"����*�h��t��h5N��ݽ�[G#"��F�S0a2k���]-z�J���D�P�'v��$A�&^ ��5�<{K V֭t�c�9�'%�����;�6觸�)ڋm�N��-�N:����R�^�1� �2�+�S��v�e�������~2�2-J�R�عF�>̛���,\r��$p�}�̰��J{!i�o!� �:SSڰ��ۗ�n�
���0^%�7SU3JĖ�m�X�qJ�l�B��&���^$��u�
�ou�P�I
�-P*�J^B�Gs/ţ֚63%�RId�u0fnm��5���*;�N�e���`T�v6wJ�Ķ=$[�^�0V�̊�S"ǖ�U�cQgiW���s 'z��a�qޥV�3���,���wwE`�t�Q�Ж�j� ����˺�4���bz�
�c���X�1��t6�6�l��q�l
�4tVU��r���z]��h�Q������L���+[����k��+�b�+[j�e2�cͥ���H�R�`����b�[i�L�q�&�,�w1�Y� �/we���ʳ�L����L(Į*�J��F���$Z�KG"���#q<ڕ1W @��r�7����B�RF&�of��<��؂ c�0���E;z�q-uqj�����.�R����W�emkfEP��a�����qQ:)'[7+�`a�6�2�ɌVJv�3�Tn$ٲ���U+PصPqY�\Lǚ��rk��$L�^LDX/0�Y�mM�1�B�<�m��i������+�Yx�*GdM��˻�]9����4D5�zT�Soc����9��7`������ N�U��9sDT&�*L���Q�8��f�ȨjS"��Lv˼��ܡ�*���6S�-H`�kNbU�V�2���TȠ-�y���m��+#h��Q%��n	�x�rQH�a�s*�ɳY�+.��f-7@��¯^+�:�6�u�䱚XI��5�����g*Ĭ���4�d!PK�h�kUi��SpSp\ݛb�����C���-P��
&&9u�E2r�=.V�/5ԭ��f��ڏC��cǌ@��h��25u�n��Dڦ/FV�w�G�m�����$F�U�-cpP.��
ں�s�І�o%�u�7��0��&taRT��.�j�C��2I�
�#[b&��n4r���l@���$4@�� �˵0�)�j�Of'5\��j��1C�특nڧb�`�[�'�Q�6�iK���.�m��TL��3(�f�����F� b����P�kn
T�[�XD]�s��70�GǛx ��4,�q�E�?0�1��8fl��<R�����7)�%�i�ƀ�5�r���Z)�(���!V�v�C�v!�l&of"j"Ӱ"�[0�4J�t�2�(��Gq�^#�m6��������ō��oE�M�� ���U����0��=m�]\ν+
�)V1Գ�)�R�p֋c�Yv ��^���D���
���ƓWX���J����fXzJ�V5^��(]=*�h�b���ı� V(��߰�^�6�]�4@I(1���d0��
(�n
��2~���`��b3E�(\I�_Pى������?`t�����-�c��o]�.�6M�]�njS�
��tx%�9��@�L��F�eACF�
�(Zm�@�`QGƲne#����J����^�F�l�&/��c־d,̕�@�m��Z䑬;���N�c���z�f*eމi��eڎ��ϞH�u�f��C�^�YxI��+*ըSM�b��X&��^na��� w6�կ+�9p�2KR��(=9��6H�h�Ѱ-���N�w�59�JVT)ͦ�SvTw1�9wG�i2.��i��j�n�Ƴ��l�Yr���cQ�QQ����3)�p��,�_ej��r˧L�y�IE�jhjj�I6�;�0��6fa�P�LCBከ�V��$�Q���U����y�
�]\�YQF�	�EGV������BY�lV�vRVc���D����%����ZYA-T�l?�m&2;*��$E�u�eb�w�;`��Ƕ�B6��v����R���ҐX���*�	(��V&�Ȏ��A`Y�QkP�L�b�*׹y�	o	[Z���YBѧ�*:����i�x��ձo�P4A�ư��MU��wj���Q������@֗�KY���[�Y�s\I���;��`�n�R�f�h��.��nn�5�T��t��f��,�M��b(�=����4�\[tF��j.���Of�Wb���Ӓ�͸��?Y�,(�If��.�a��/FG..����\�5���(*n�,��6����àA2�(ma/��ܙdk��B<8�r�(�R��1Fk*���=Q��Z����n�3����� �SJ�zu�m%�e�I�IG��Ȳ�gpF��Q]ʽ�)���*����������V�.��v勅�HC��ihW,�6t;�L$�\ŷRb%�m�h@��.0�	Z*�V�-�B�⺱*��j�/J2���v)B(��rJ��i��P9�+������jT!�L&���T��X	�5�F��#X��ط-�/��{hR*�`!�jnU�/���r�!t5���b]f�ۨ�� f]ޭ����ʰP�8�,l��f�[�&n������A��n�
p�=�b	V�]aNR&F�i�N�������U\�m*�w�H��R��@2�Տ$��PJ[���������9rkH
�z6�vK��qP�N= %ut��v�o�V��&�X��дh"�5*�J�Vw6�,��hCn�Vj)TX@����B ����ʫ�����-����uI*�/(c��Ғ��z	g^SiM��yC�
�Z�����:�˦.���;�A>�i�m�Y'7:�kGh����7�6=��,�X�u �˰��#{*e�7��iՄOu;��J{*8��Tx�xoxeJ���e����t�Lw�{L�2���V'N�ѥ��0�W��w(�e�s��������^\�Mp�{��:%.�0�4�톦�c_ڍd�}g�����u�lEˋ��:i�
]�rZ
�-�J�^P|)'�lsy}�4�}�ϰ]�8],�z��t=�����T����尾�SsV�e{ɝG�lZ;��)2�Ւ�U��<��s�=rI��MHm�5�C`��eP���y�e���ޖ
���\7}@��-��C�:�O'�:���dGA#�����O#(�ir�Z�6�\=}n1���4��5�S�j��
+]��AVu���
r��LU�z9�v՝Q��.��f��pE+fd��r��?4����ۧa�YK����t&���F�>��o>48��{�o-�wsd���/�d<�m�@m�77oq�ll]�̍Gu�ةZ��*��bѭ@�i�2W�e(z�W��*�4E��jpi�ʴ�D]�=йv0Hn�vQR��J���Mf%�:Y�/j7k�u!D�dڶ ��(wbX�����u��Nކ`� D�r09׽�5y|��+F���[;��E�W�+�n�ɬ�ZV�9�Q����r=�V�����}sZ����.ZL�k�&Q�WOw��QW'w���&��Yo�}����N��$P����V���
�w�nUμ >4ܙ&�R�ѵ��ۋ�7}-���@�X{k]Cf*�Wھ�մ��Z��
��ړ�k:g�Dc�#� *E����4��q
|�847e�%�wS�,��i�p�&����*LG���;+�\�)h�Y{�s`�u�=�����o���v�z��!���l�l,��Y��f$�x��
ӷ�xң����ct�q�����m-���W`S��V9�R���u�d��kR�usl;�y�'�Y��`��vQӛݠ��kUt=�ʇ�z�WH��qLWyp@$�����9e�
�.{emC�TJ���6����6�`ꊶbI��1:�
'`�7/sƵ��Tzi�曷�Ei$�����w�t9݌&[�b� ������U����&h��(��2�l�hF}+��e�
�uDs[;z&�P�,k����:07'\h	YSw�s���CG���Q�u�1
�Y�"�cJ�ݵ8T�x�^mI�.��l`_g]����ޤ܅1Z(e���,cq�G҃�0b��=������մی�uq*P��m���kx��r��; /�}��[�]#���X�ˍU�c*���xE^î�2�ۋ/�+�����t�;N���(�fK�̣f�V�jRXݛ%���W[��1W1�ޖn����v�O�1I20B��-v�P�6�9�-��H'!�Qh�Q�q,&��;K���Sc�C��F0w���a�x&;�w���4����Mt�P���:�N��1D�Q�̷sMؽ"�	�_ʀ�q�ygbG#�n)�q8hښ$t�q��ٸ����PR���$��=��[u�C�,1��5n�� ^���գ��B��T��nU��'��sr��p�5�G{�M�gG�]c4�hEsI��7Z����c+�֢ ��5G��t���
O-S�����yNz��x����︋Y��
��+8�.,�u��6����V�mԗ�v�ʺ�Zi���^�a��=����M]���i�Y�˨1����\�wy��P&��zi�x�X´���%��=�̝$��r�k\j�r���1�
<�[:"�KDt��\�iJ�
{)�B�&�+��ujH�����(�Y��V��X�ӥ�}v`�t�84��V����]HBoZN�T�-�Jݹ��Զrk��5g-�<��PɲhѦ��N�0�KԜ��Ӯ�o��YYӴ�&�/�d�q٣q�$�E����Ի49A�LXZ��cB�{|0�|�*��؃�D�j��5�"eM�}|0ll\�-S�m���wf�s���
.�YjݍX����Ol��5
��t�%�\��1������g%���G��Ud,�`��<�C�:}�kn�;e��2��˵�Ymc��)�.}����������ްz��}�Ѭ��D��_,��,곷1�F�1o���I��n5k�F�̰S�#��ћ�oq��mv�V	�ɳ���6�뛴��o��u�=+�t'(���^��/�7��ܬ�\(�/�~�0P�d�/N���Y��Ҭ>�ͮ1B�	���Ga[��Z-��>��y���k���43Cb�|�A�����t�{�K�p�o�g$�X�%��E��_>�� �P���u�W���t�ֲ����0.��.0k7��u ���,�@�YN k�X�Y�7U�ւ����wU�3C]��s��ѝgv�[���w��ܹ���Y`ݣ�%E����3zo���oWK�75���3�r�J1ɛ%��\n�ý|�k�Is�<�smV�DՍ�HkI��4y^+V��4(�2��Ef*����A�����j�T�f�3ͭ.^nP��M����;y��LcUp�y/���ڬ^rN�An��(��S�j��-\bn�L+�[W[�������Ӵ��udmu���|�w2WT�R�����z�V֚JX�yǷ��E�L��a�]�*sf�T�W���pP������m���8o�B:��e�T�`�zRǄ�]��hS��Y�~Dֶ��=��{:�1�
#�J�t������c�LFh=69�gF9�g�MNR4R0`���sǋ�U���`٥f�7�R�:��Ms3�2\��vm#yW�x˙3� �ͦ���K0�Ւޱ;�њ;�+Xo�b�, �VTA�,�+0��/�=ú|��U�p�m�jѭ=ʗ1Ӌ�k�WV��#ӲX�J�Q���ǽ}[��i�EӁ�����V�Ѝ��X�WV�����I6�C����wJ ���i�%����˖'�e�U�]񳖲�P��F`�Y�*��ûoie*�ʾB��OJy�S	f��]�Ӵ��e�},�aIΞqȁԡ�=�F���6:����,0����*�a�*�s��r��
oqtC���+�K]���Vɫ1[J�
�V�yGd$u�?.�+:���V��}3�IwR�E81��]ve@Vk7L�k��i"��6^h�ٗ\t����ڤ�����|���,��k�]!�^j �lK�1��m�WFv$�J�F4%�	�d��+ӽ0F\v�f���w�l��#��;(X��/&79�n��u��Y\��h-�G�X�E�o]霶�A��R\�;��}��!�y��n_�0_H�Ӡ����jȫrJͧ�X^�s�n�\��8�|x��5�w;�ֲ���9��#��1�E��e9��\sej��5��Q��;����u��>͜��ab��b�l�R�&(O�n��4O|u['3w=�0Hd���l��YSk&���]��۠�+���U�]���or%�]����;�����v}�&j�B�-��ZW]�a�,����͡�+�)w�bt�%�-mJ���nM�ϖ�h��\:`��;�8JWX-�G�6�x]��Y&B�k���NμG�w2����]yJޕ�X׍	��٨���Z��[Cu�|ŷ6c��ţ;Q]�V�5�}�q��ŷ9̭֎����8�.�$� 5u�݂pU�{C�����/���|����o_j�w%��/R�`���ՒT�V��&3^��u��Zkt�[���-�j��Bƪb��X��,gU��ZV/�)1`�-���,��cF�ZeL7bVkYūH=`�b	��N붩Z�p�x	��\�[yc���j<� �qWd9��pa��rX��V�(�]*\���ԃ��*��ִ;|�ZD�r� �ea/++<��Ԭ�;&n���)�Aϔ��jq		IM]p�nm��r�F�.�x���b�R�l^�
9����G�."�=W����-�u7YE���]C������ea;	�u��uL �1�7{���U�CF8;m���@s����j�D�i�ogl�K�{�)"�io�U�5i��{8��d�-�z�/����Cgg!�TB�1S7cY'f�ևM��J�qУ|/{������,����{v�C����C�s`Cݑu�h�[���m�ܩ�A�^]b,�2�X�P�+]�"V��_a��)�TyW�鍥�K�M���d���ɹ��g�kh�l�;��\��[���g,�_ (hѳ32��Y�����;uĸbeF9�U�'9��pyCf>̣]�]�r1���hJ�#X�����Y�e�S�h���n)����:��X.ֲ��k]�2���O�(�ܒ�sK*�E�WB&�lɳk1�Ϩ��x��n����oJ���ȰЖХ�wܘ�_�t�]����˜��Ht.���n�_����Ѡmej[Uԟ��LYD#�-��TۡF-�W�AQ�V���余�]�;,8Fգ�ֆ�a�Q�g�y��ʶ�̠;�b��t�_"��ج�	:&x�g�n����t����lWu���[iC�Y���L���h��S>���}�`�mcb6&�3Ee�v[T9�ܐ`�}����[��k�^�1��fvK̘����Jm=NJ�|,G��[_e���դ�C약u�o�[Н�M���Xֈ	�h��
!}���)��gG�&�����4* _8�q,�k�k��v�sys�@	��ю�^:۲V��H�E�z��w�-�
�
����F�:R$��t�g4���"O�ڻ�s+���+	�D�Ȓ4M��56��v��*�b�3S2��Jg>W
���3z3�u�ʝ���mZ@&CwVq]�g\�d���F�k���[V`ǃ���wIW����,���]N�����|��Ó3��٪}EM]��N�*|��:*���ev.b%`r��XFp��xh�:�_#���`��Wgrj���U��2%�Q���kY����B΢���ǹj3ZA=�N�ф��c7[1m�5>��B��vi����;z��O�%3
[����o9��ҩkV+}��:[X��m��|���o�0tt��r���fe̋_V�=.�֢�2T9P�j험��׳,hRnjW[N��i�TmV��c�+xv�RN��oE��
��W2��ě��8U��ӈc{ǎ]̑>�Gi�!�6�V��&����˽B�H�,�g-�\�A3�1��$��r���R� �]1��Z�]+�_1����:�mb��	��E:-���J�B���s+�*���'Ȍ��r%[2��a�j�d V�ʮ;֗7i6�
y*�.�X��t�v�8DZ��^�w*�ٳ^�#d��w8&.���!��*�<��s�(�kY�s`�]���b��Sv-��N�U�*���5�6U��<M��і{'!E�l�_�W�y1��汼�83���J�غ��ud���e�>��-��Ի`+�gV�5��-��ٸ��)jƲ�d�sx�af����:���޾���}G���H]����T:�U�Ju����}��pl�WE��p]x�ßL{}�{v��7uy;��7��[G�1�}���UХ�18[�;�A@�&:y�Uڷ�V�Z�=�Zƌ9��F�H�%�+�Yϕ��H��z1B�iM��B�=K�o@UH��v� \��ۗ�üc��MO'�ve��d����-�z^��(f�jT"�B�x���j�L
]ުR�]yG�Y��7�٫N(|���ST�|f߈�ž0D5D�1x72���
|��3&������uɡ�>,_TH�J�U�Rto�%]�D=�[n����/f��	�����Ӳ�����7-��ˈ�Ւ-̡y���@T����6�S��j�Yɋ�{�O᤼�Vܽ��z�iX͵Lc��k\�q���'6�u���'qC�;�cΡQ� �B�2��yn�W�in����W��'�N�'��]���AӞ]e�S
yh����$;1�o�9Gi����5�_K���Ǩȕp�3�e[�3�pd�n�#"�.��\0���;�|��+qt���ZT��Û�s����r��{#4e>�N�
����s�Ӝ�uw�Z�uJ�jO;�2u��{n�A��W�a��NMxi��e�G �X�d���pV=J�5�X6M�%Bҍq�,d8��3y�lm0��9\�M���J�p_9�ɽ�6�(]��&��ʻj�_p�l�m)!�E��r���|��:��@�*�[� @'Ո]�)�����w3��Bἴ�s�|�L��g6���?��Ycm�����Yݐ=2�h}�9�Z�W|��B0j���pHv��j)Bmv�z�l�v9.�� (�U�����Xfv�9��g�5r��^_�虨q�0�c(Ә�w0�S�eX�d�\��u�b|��d�`ٿI�`������υ�Ֆθ�s�����1�#������N�s�����V;���<��W�2�C�dX.D��Ś�9���GB��T$�#���+��*��B��-b��ȼ�]�+���� 7Gf;״�IY�� ��8[o/>t��x6ۭ�ݠ�ڐQT�S�Y���`Amh8$��/H�`�n�)g��������v7PN�3le�<�OtKt�v�����dũ�F˛��39�g.�Ö�Y���,;�؏)�c�����s��o�v��Ӥ�>J)��G�J�0�Y ����X$΄Dr�1�p��&D ;�����sM�v9�����P�[Y�	rɫ=�|�c���+�v.ͱ�G�z��p��z�ΰ�co�D�q�I�Cֲ�Q���+V��81.��.���e�՘��G��|(v���T 6�m��\G��;y���6��B���E`�[ЎM��;z��k��� 
��TE{������~����\��V���h�U��uL�5]Y�̜�I]bF�VZPs�O�R���&��)#s*aY���5�l�L��Xk�r�m�]uk�geb����2�����1�M쳠��2 �-9�T��qvzr��n>�:���W8-1
T�*�S�Ϧj�wZ�}���:I��y��Ɓ�5ʽ:�R��}��ǻ�c�λ\Vg���%�4�o\;�+l͜��;d�ܬm[*��z@���t�Ÿ;`|tr��9�����ɏ�K�'7>��yVN;���K�2���an>��x6�'~��0&�R�cf��HzL�밈��r�@Q�2��v�C��Z�V( �+Ǚ��.��2��s�n�F��eGԮ�v2��c^�n�Nf�;'�����ٻm�*`��3�V>i�	zi�n�c&�up�!�Dw6���U[�'C��SJ�uM:!ucu �j�:�d2#�z��ӌB��2��:�T}6]#["�"3�rx�`yX�IAj��o8�Sw�6 �&��xzہq���;Ѕd���OM�׮ճܒ=�9r毻�$�̋V�yZ"]�}�v�7M�B:�U�'/*n����o��iЮKp�vK�Né�=�]a�q�)��:߯e�Z�`�5�4��\�v�5�V#\뭋�j���:u��K�z+�HZ�W�n��[tV�"���� ��XD��Q7�f!�66�9�&�+�|mL�y,6V�t�X�"Ӻ��:�U��N@W	�OOcô���S@�M���}u˾�W]����-�1 &p���^k%5ϗ[����6�5��@��R7���)��hVĨݡbﰬ�Rх��^'x�~������Pl���1�
�¹�������-�&�aʖ/&�*��n*͕�����ˋ�r1��\��Q�]�Y������ {����V̳�i��Lx{o.ܰ�̾:35��yء��,�wJ�;�&0k���xS)�ߺ+Y�\j�51�ۮ:�+Opڕ1�]D�(�8��!7E����Ẕ��]�>)���֠pFA\�AZ/n�hWuy����TÐ�����D\u�Qڷ$tn@�M:�뺲^��*��Q�7@��I�+qS�	�;���gv�p��y�1u�m�lo�#G5��F����\���˛�Vd��s:���֝����iI:�X�:�["�n�ox�%�?HC���b������S�zv#�c&��6r�N����p�WS/�7�G��[b��巏��OT����p�%)J-��b]^p����<lDg]��=l������a7LŻrz�ˎ�#y,ȹ���LNĬ4��|-��o�jU��	9�yV�5P�Q�����[ˏ	�m���,Rc]7mv��ݻ�J��$/VC�����Ψe\6�o�,,��W�����
&����bn!��4N�ײ����]%1Z�&�9�U{9L�78�1π�Nl����,�xT�C᎛�7OQJL������)������,qѴ+8ҵF.:�&�&��厒��/)�ѩf��8'����:�����u��Ld]q�����9ΓA$�Q�Ϻ�&�m��c�&2ph���R��Z��K�0<�4�&��mJ�A#����9e=(��쮫�]L6Z˾�R���$�ha��[X�:|�np���%r�I��]����2�&z��0���צ��Z�pJ
��Û����}��-�H�������Nä�'Ř5��|v�����z�^�'��rIp�L��Cd�-�oa�5.���Ƣ{Ov�6Z��C��lQ�7bh[,����u�	p���͈3��H룙jR�Uј��ت��L��k]]V�V�S^fX.J�¶��A����3����&BZ�(�&d�<A�xg����5�/"hm���UY��v������8@Q�F
���Ƭ5]��9�]�.d巆�u7��%&���;�S�o9�ΠYl���H���{�M[U�� �ѫ{�b�n��r��vU��+߃Vy�.{-�pt��g���z�T3P��Ms=v�k�JMЭv!U�W ��N��(��\�WǤ�������-R�c�{ǇCn�)8��U���u��y[n>mXsE�2���l4*V���c+r���m�$����u���R}��lYF�H�Ǫ�飔�NkIm�E:"Z.��%�V����ǵ�	2�S�M*ty!ʲ���l@�{Ozo6�f�`;Ϣ<�λ��!�W�.���Kα�N�H��`7V7�}�X���̭]�.�
��)z;�-mѩ���_h2վ�5Id�r�wj��Kh��z����Α���+�3�Q��'3U�ib��C����=C������ܝ�)��рa*��Y��A\������bS_wjpVJ���@9ʛ��ṹw]&��S���*nZ�Љ|>Xm�u�t�*η6�͉���Ǐ�n>� ��-5�WC�,8�ݲ{e[Tcڤ��唆��B�oQu�'���W�)��O�~�X��-��*]2Y����̈́�ήQTTS�K�e+������'��	B@�YԴ��1ZJ���l�Ŵ9X�KL��	�sUű�7o��Dc|�-�Y�˼�=YF��N/�j�F31[96R�̵�
<:��m$:�7 6���l�g_n1A������i�8p�l��R���_6�}|&�i�3y;MZ�,��ʲ����&7�����{��Y����'�˖��M.�	��ZS��kPR�8M*��wr��U�`�b�Ven"�s�Hx��[u�fU���I�b� �]�y Y�6�!a=��������,Wn�s��V�d�CCŮ��YC�0T��-����ү!�oh�p��#�}wks[T��������� �gf�Śk8�S�ǀ ��$쨃��-�H����9	�0g8�}�_����L�%�u7w����D��.�W(�+x��N�m�]mq��E��Hpb�������k��:�T�S� ��v��-u��ͭ�8��R�(]-ɋ�G8�*[r��#�/���Liz�c����Uf����/H�v�T���c�V��uǝ��>DTZ�e7��Yi�p�ǒ�򠤹�����5�n����x�e8�6K]�#v1.�^���45��x�1���s&^��Ӹ�� �/��-|۫�yv�ǫo�x���! ctΧϐo:̽b�����iem�>S����/YΣMns.��t�V�����6�υ'���HcM&��V"�W��V�]N۫c:d}�l���#[�ѣGm[:�B̕{�GCq-WY�;��g�ѽ�}���b�y ��q�W�Ћndb��*�r����kMe�c׵g!ޮZ�s�Hf�r�hh�8q�s��4uj�Ny�j���;�x�w�(��Sq]���:�[���xmc�O(���� K#�؞;]$e&`T��]�{�Z���o�ϲud44�s-�7��J)�<)���*�y|5���F6*'N j�@=k�f>� ;%#�{v�3��9ԫ�uVr�0��dӰ]V��a�����@��.��ٵدb��v�����Hn�ӳ�K�瘏S���N�ԍ�쎚�
�q��wu{����^W#��p���[e�m�d<k�Bt�۶9�(����Q�ۯF1c����!���5��T�;9�.������\F�h6v.��YQ���%֕���p�UF6=�|*ˬ�9}"�[��u������J�n��e��+��ZY)oJW�S�`B���}OvV0�fB2�Ι�gP�f�Sݚ��n���U�g�u�q�Y�Y�{]锟 )�]�d��%ʂ,kD��ؠ�WI�F�k�gv��i���똨���s_v�U#W����B��,���v�����[��/M	�g��
^Z+9FQ�}�X��묶��u�������2���K8��&K����T�Gc�C��3(1��j�t0�*�meXи��S���p8�r���&r���Շ]V���Ŀ�x���s7yXi�N뗤+s�wev��]�jP���t	n��2k�Q�2�Y�*SYNof�s���]c��;q��4*e�J;:�ƽ+4c����l|��`�b�$~�q��ЫHpx�&��[��zj X�r�;�ޛ��f����x�%�75���tk�0�H�����P5.�墷�Wg)u�c�{�	��m�����/2���cز�������A,���uι/X&�H�X�l�θ17W�ضKPhh�}�����\&��e�2��o�����t�z�2��[�F$;3�V�55-��K���Ut�@U�R�Z}/ �J+��{ܷ��Xg;��e��Eg<�;S��@��V}{�o	=��k�����u���f�@�<���
j3][Ύ7r��n��	�.�a��L�"�|8����\ܨ.]43�ьѼ�,��P���U�ewa߄��U�����h��݌ ��U�C�c���I�X޲&�Ȼ��7�ao��dV�=�g.έ�0��#�tZ�u�c߻#y�y+O��<�^�Kx\G(�4��e*���]G�*n��^�)nI[|q	S��*�����р�H���Ϣ��*�x
59nc�����-�!����J0�t��R车(�D�.Ʊ���X�v����wt}�)m�#\�TK��P�)bI��K$6�V�**:����|˾t:�-����L�]��V�����f�o�<��{sA4�ތ{3)}78ӹ��un��X���茐V$;����a|�;)=
���m��j>����6�Mէ׶�&�Vk�xdfK�z���ƫ_7F/��@������]��})$��TݭI�ԝ�b�ɲ��[uy�a�f�٣����,���i�b<k��S����ԃdue �<؞�m���K�'{�D��hˮ�u�]!RZL߻o#']ˮ���Bi��Xډ]�.�wțR�s��q���o�R�++�{mC�fSŚh-ucB�\��)��WWk2d�g��6�jX�N6��f^�Z.;��󃦲R��y����E҄U)�w�nK.�iN5���K�2���-l��^�<��>6�9|�H��϶�`v�xe>j���$���í"�����;��.�b�ܥ*�di�R����ͬG]o~�hY����8�����ԉ�
;�븭��Z���2���x�N�]��A����70j���|o�Mިw1�2k����nv��gpZ����Y�V;�_m�[|�=��1g-m�F��k���X�zf�g�ސ��!�ەH�h���UzP[n�F�ac%u�6�R]�J��w��Y�_��`�;�v뫜�(�O&�Uw)�f�Kn��Lu	t;�	ԗ^�n�1o��:�.l�0���;J�s�.ú�B���*����M"7p/mszcS�ۘ2v��u��u�bV�Q����<뀾��nf)5��u�7JC�WfvUʤ�n֗�ٽkU�V�MЭ�E���9���zZ�_JZ���Dp�,�:(���/;���5b�jv�U*�"��k~��p��7�k��L�$
WMwN��E.�`��źۈp��U^�H���/���T��n�E0�LU�v���N��[U�΋,�|cCvbݗ2�4i
��4���cer����A�Kj�v�utW���|�Z�ڶwCkԔ.�Pݮ39e�v*�άZ�+�8ՎA��+y���A���ѻ�-!���{��u�	����VP�i�m������3�&5R��f����K#�&����+}�Z_ �b%b�mf��o�W)Xv�=��΅�h�r��m��ܬ�n4�W������)}�5Y�e�nE%�]�s>�� tT~P�-Kb�,�u۟і؁�e�wM�}3���Y�tŖ�]g%���[J6�3�4�B�V��^]��H�ĩ��u�]Ȅ@+�u���وf�c�m��Z�꒦n�"�{b(N$��G��h4e�5�R&�4lm�
����#�[J�n�:�]��H߳d�����c�!n�
�s�Vt2%�.�ԕ3R�h+G�
�|��=Q�7���v�mS�n��Ƥr�ާ��^Ǭ��`��.�c�29���,�s�7�����1y���:Gv�c�T�� �]�iЏ8���h�U����z�W͍�*�3�!��mRl�}p��5Cv0�ժ�[hv��J���V��R�R�8���:��C���|6�4��J����8M9��m����S�Wp��@�1�=�K��U���Q��hE���ղ�����
l˫6T�:K�l\ꕿ n�Y ���{V;2�Y
:�1 ���M9PT���冲��U�l�v-���|���zή�q%.�zأ���*|
�W;����@��U�r�Q}�ed�l�%M�S�N�:����t�ň��oP���}B��g�wI��Qne;%n`4�4[�wб��2s�dIvok6�fu�ζ�B�Zf�a 7z[����Ѱ��{25�,F�d����M�q�p�+�Z&�K���]%��#&���`�Red�j�z�a�kr�=��-؅,�u��lF�#�:�����Hk%Jڷ5��Z���W3��g��B���0�U�W]��.�;��0{gC[·�n�5�Xu���yK�{%3v�g���]W9�*Vۇa��|&e=՗��oio�oQ�dJ�FŞ8l,���seTGb�oS�zD�op�)�e���1a�X�O���h�`���huݙ��N�TE��������7���:
h�E�j�;y;�䰞÷nƘ; �N�)�������kX�+_��-B�����d�]��@.Z��ﾯ��|�P{�	},cMA.�x����:�է�v#b��swF�i	����\�%K}�Jҝ������j�%���$�sw�
�9܎0�寸+IvT�|��=��ԝW�kuc�]�o�Oೀ;�&X;� �Hnϲ�L�J��-sp0kvZ�<L�ִ�_K�H�3��1K���n���G&#׭�5�	�t��ҰʁA�k�h��n��49�s��t=��ؙ1ke�ۏ�c�%�gKH�ڤ8ʗ��e����O�j�j��p �@y��C��kV"k*c�7�^��cZ5;M�#&̡�.D��}f(T�/r����5ë~c�/��NfL�oQ"�UFS��ͫ`��r��wJ��la��"��K�ٹ�ƺʀ��lf�v:��iVu��H<��a����i}���r���`h�D��vk)�+65d��y8Ҭ�m�ר�K�MM̨)�|���Ef���k��Ŏ����Em��$G<���Q��/D�q�^��T{��/àtD�7��k���We��E��m�%��&Wi`#�C.��fw˺vhb�����7��ELV!Q
M�pQS�3�<�ֲ" ������}��vo��S\'sW�op�Ix(Z��פ��i@���������hT�&aw r�{��ܟds��u�e�/��U�PMl�ӥ�N�2V��	�N�E	���ti4�t��l4�Z��m��-�-�@JPj��N��RWZi:P�z��c�):��))�t�'0h�i��BSMI��V���l�th].���P�"P�T���x��HSJ4,A�]�IM��I����E&��AHi5��ӈ�UJ�I��.�T��u��:(z���+K�i)�4Pt�]4�#M����Hh�i֎�M��
:R��F�(�JMul�x�����t'N�CABQK�AEѦ��e�JQ�I�-HVڊ;n�"��j�`�i(M'Jh��?=޽~�?OWo�+�9^��p�\�.����u��4u
Y�����;��x`Ҿ;6����)�-��u�Y�̘��pՃ�������'���e�0~B�|LKP���]PU�����P:xQ(��t9���]�֗y�#�_��k g�Fg$QB�o�>���Jm���Hs�F����h���W�P�{��G��L��OyY\XU{��*lg���7�}ⰱ�u��hL�w�zϴ�]O-\П���|�؟����(%� P�C�V�-��2�!�f��T����'�����8jP3Y\����R&"�e��sCj����]F����Q�x�'�~��1mA��<< V]����@q�@����J`��'��_s{zT�۝��1��uyԸ#܌E�s���gD;��0��Pj�'�SlͥO�`Ã��y�f*�!yz_�u'[��{����Ö��a��H�V�������*A�ϵ��jk��g�v���Nc"��8^�<k�db��w|��R�,?A^�J��"�~&���ɫ��TuU���z��w���^����|yEV�`O.�f���a�3�8V����ڥg�͏n�7����L>�����ky���������v���|��z=�~�5	�[tgu��+��c,jZiu���]X�����
��ܬ�˻���p�Kl΢���~�[�o����7!�4�$�'�0Pgr���m]fi�+��ʗWQ���h�?5���m�i���ri��T1�%ѯ�R�9w�p\5�-����o�;@����5Ѿ]_WѪ_��0���3�B��U�J���H�z]҃���V��;n�Npf�|;:���0����~ A��y��:�N���twy�u>;�v�O��\j|*��?D�Ş˱d����6a��8�6{�^<�;�H2�}`p��I�$W�Pe���Cn#&#)��x������0�6g$;��뵉���ߙSW�%������M\��y� =Tiu����@��G�[|[$N��GK�k�Z�i!XW����ʘD�������
j���	��C_u�m��֥��hw���5�̴��"F�6:M1��,g%�����VOW��
�~k���AorZ��s='��q������~HV�M���Mj�L �gM� �F)�K�n�C�ۮ��V�vRC�����6(��t,��W��c��J��ë=�c���^����Sf�)aQ��G��c6�#���Y�oK�.Jp�P���3�{oʁx=OH�f��f�jk�v�#�{0	�����̎<7��i^��p4����8_\��Y��aܵ�m���c��n�]�t�l+��l͛3���$B�U���XDk�LRwf�,��^��VV����i�G�Ss�v������i�5(��g��s���ō����U��u���~�w|q�;�8E��4�w��M��*;���'�`��h����aR�,� o���蛠���gS�y�,Ə��n�q|�-�ߗa�����`�}�p5�Z�E�E���ʼ�}P��ݶ�S�~��1a�����ԅc�~<�'\���묟w�|iz���ޗSs���+s��ݢ���|b��`:�{��V�x:��	���p0V��΂��s��%��6U���%�n:��,Z�q�қU1ek��*~��'�qoip���U���o��!��:J��c���X._�ܝ`����jy/ƥV�����j���Nf�Ʉ��vW��)�}P�jr�<�@.�H�B6��p�ՠ�L���P47�OF�3��T��O!;����vl8��T��J�_W[G��J�θWD^��3��ѯ+���f��
�ć�AzB��������͈Uu�7��qc�S���T��WO7F�'�@��.�}.ϥ�NȮ}��y��7˾�Џ��߈͔7ʖ?D�<�\���G[�d̬��qi��p&S�J��(mX��ӝF�� Q��qw��5�jr\fuv�+h1�p.�zjFs�&���\hY.���Ǐ\%r�[o�mG۝�{�ƉI�'@��}�M]��u��{E�bz� �/ˠ�[�^�V�����`t'_@�#vZ���6�r�&�z��+��}��5�6�՞���_u	B�1 s0Y������[RW\>��]4K4պ�O��x�	1�Ĕ�]�oȼ5b��U�.�G��VXT��}N��L�b�T%T��.�	�M�Y.ɓ��ü���x��)��t%ǡGEX5�{��-Qzc_��2�+ǆ#b�Wz��I��C���ᘕ�m�ƌ��}5i����kU�E�#{%��fUJc��Vj=��U�(�+�k��uݲ&{.�O� ��d��>�^s'��Do�ܳ��-S�����_ �h1�^��ΰod5�Q��/iC}�S��s��1���EFGD\�3c�#�$8\���os��\�g�\f��~č���}&�߷�%�>��p�eyϩN딡#x�����<+k91伅�N�hMK\C����˼�SޏG��0^����}*�>�_��?s��^���#E�pe^��� y�ДA�v�EH��e��s즶�OGZ�/�t�{}6�B���3�������e�HV��t9Q#�%�-:���)v���d
f>��I�X��9M��댊�$�Ίj�k���^bڊ^�
*O�p�j#.=;��7�B^�9E*u��q����e��);c�IG{��1�\������\4�,�;����Ym�]�$X�w��1A��W�b�S�~�-��Ӓ�A�)��@F�w;�i�2Sk��zs�G'�����.Z=�?!gˌ( �.��W��&�դ��4�:�S������쑌�_Ů�WC��fD8`��~�WObY�/[Y|cS�}R度��b�g��)��{U�
��8p��]t�c���<k&���~���V�w��!hQ0~����u� %+���_o�UZ�[����1��Q�`��V�D���;㉫�s��g�	��S�!�`ޏȩ��|~`��n߲}�/
*]��RY=����6�iKէ���?��bS�,��|P:�CP_ϒ�ᔽ�����qx��nGx���k�k)��N�51��e��2�4Һ>��=�q�ʇ���Q74���{^��d�> V_���E�.Ujh��偰���_c���-�hgX#*fLƘ��rh����)�np9�;����-�y���>z�J�L�����u|d�~[Q���9�*�ys	r[ǜ��8���vL\.�+��^=��Y�D7}��[6���E�5�Wu��؝n��1Ƶ�X���74q��ϝ�K�/�{Ƀ�vZ�c�-��.�̈́ �QL�����I�jꄬ���t��*�ÍScd������=�ؙ���̊^Hu\�j���X��ւ��Ӷ���[�TX.�
@�-G�����Ԅ/�S80��.�WsU��c<ι��k�p��Aj��NzԯGz��{W��4�k����Y����篅Z݁/�sfp=*v?{xc�c=�_b_�eK�y�v�m!b�n{Ke�P���!��F��1��X�$V�>�VΝط�=[& �:�����V��:��q�����>��{-��/*�֕�O��d�7$�Z�껇�Q�x�~F�,��n�"�Au�l�X85�eo-z,4|�8=�z�}�E*r��K��L�7\n=���O�5[ا蘳��Q3�c�������-�QDr���Ir�磣�f� { *��\:�$7R䋎���B���?Kw� S��9�N�H�HY��
ɝ���כh�N�a�%���ҝ��yr��@Z�����8H�6�X���jW�g�#gw4e���k�J�N�Nk�"� ���hom����+j���V.�Z�/i�h�ߚ�`���p�D�d�H�]嫐{1���O�J��"��zyd����5���\��r�ls����mV�b��-�W���]�L�-���jW`�+`Oor+֢�ŋ�I��/N��Tu
��ʘ�'�f���p3t-�$
�������Oo ��|�I{Äb���V���X�c�������:}�pW���j�7�d��G*�/���-�!�[uI��٧vZ�ay�O�\<4!�+R<C�U�}rխ�9�ཱZ7f���y�5id�W_TBkțR3�O��W��c��K��;=�V> *����1�"�(���Ԧ�M�F ڮ���u�*�׺�ԣ�ٟsƅ���ō���u#��e#�і[���ʕx�c�@Lab��B��!,؍��=X�س{���2[M�O�_����OwL7�4Ə�滁=+�ȸvw�ߟ����+��s�U��5�xG	/�pC�f�>��l��{@D&��Z]��"3b6X�b9u!7
��s�/�k}F����R�[��u��1��:]��w[���K���œ\2�\7ؘ�8)��}�����1��4�򼒌�}4{�{۹/X�}AW�c�e��UvM]�F�[�UZ\+D���YδX�o+O'�IÃ�M�%9�04m��@@�N(�O��{�w�gw7����H�W�.��=QM���SVug%}X���z��^�`�R�,io�{L�{�H)��FI�*�+���k8usc���3�Y�L7��%uWV���B2rܶī��-z���ժ�.��;j�o�$*g^�}��z埳��e��xu�C�?��Ƨխ}l�Z���Z����6Q\31ګ�p'�r��u�gѫq8+���9ڂ��0 w��lS���T�����S�o��Li���2�
��'{
�k�c�@k�;�{G�2��ydT,�TP���`�X@W�c��Vw�;�~�>���!U��^D=(��Cyx�����%S�� zV$��A؜�H��]�Nqp�'�m�N2,:�R�^�g��[i�|��Dk�jNdcR��,L����:eQ����?���Q&�;�#�˶Q�¼�X\�
b�wi��Yf�mvOwE�m��61���^S\���(g�=��s9���t2�WxS��YI��Li�9�f�JVZ�RL�48KuL<G*�����ם�ɏ؉���2r�s�=-�')�j�����4̿��,��y � -,K/fpCW4t��a���7��p\轙f�k�M�5�֖Eb��y@�ʿ!�R��J����+q��]W��c9	f����7�T�3�۞7����U;ڭ�HSgr%����kR�j=���V�32��a�f��s�+�$��.<���gp�o�^�����p�Ѣ���k�G�{:J.W,�jq��q��װºisB��]��|��|/�L:�@_JƇ�k��a��E�W��z9ӛ�b��D���=�4�^|W��5k�n��UǡA�J�e�\�!��՞p?���JJl�l��eT2(��}�2��OUzC���������T�As_GE�� �h�5�+����w4s����sя}=��v�8���|�\�y�����E��U@���+�x���a\S�w�:��W
Η�0�����a�nX�����͎;3�ǎ�:�F2�������gV����]��*[���¶��d;W��Vr��^���xo�X}��2&�e\5q�c���<K��}UA_��i�fs����e^?�W����ê_!��T�&Y����;,�"��^`k����v�H�	K���S(b�<� 7���=5���\�E�{GK(��%B�©��=�~9�.{��Ч�z,Fɯ��Ug���g���/y�$���J�R�Di���	�V�܁pdW\߫�>�k�oƛk0jǠ��5g�u{��Z���C�8���!W�������=�s�����w���T����Ή*yL�V�Au6��wC���'�ɷ�nf�y��2x>�b��Ɍͫ$K�ܫ���T&��MT%�F֎`�P8�Y7�w2�fwu�sE#��Օ�Fw	�*�[���ԈY%�J#V����m7�T]�tx�t)]u8�&�ɸj@�nS�"� ���� ���|��3���~+ޓ);S�Е�"��x�(#2���P���ba8��.�a�y@P�0AD�0�D�r{]��X��*�fFaW���g���V?J𜂪U;���Ⱟ%V!��Q��dȼC|�f��!�Վ�!2�����xQ��^��������9s��b�02h�h^*��c�����-Vz&�����#���N�w�]u��e�#>� q�Ì�fznk�,�=������{�gi�B�{��[�5��lL^8-j�c�"����������ջ��/9��h~���^5�W*��2�ˆ�^�D�����`��ޓ �ķ"sZsA��v��tQ��>�y���~l��7�CW�	�/����R5�1�����h
F�e!�L�fr����W���`��}籋+h
��~��r������ϥa��V���A�u�=����k���P�V�� ���fp�c��h�r��Q|s� e�}���.���,�M-�]����횂�jv�M
��U�C��w��t;v�-)�v�Ѽ��u9�`����͒���*}�R��f�5�Gw��|�V�im��l����p���OG �����p��͡[@^��Y�ư^]�wx�u�X�1�i<���+�悴�Nx��;��8tT�`\4��tU�]�]:)�:���V+v�������V���=�-��3�g��j�|������kU��13��/��y݆��H��F�n���)ѡܾy���V����*#:u���@}9P�zmPϚ��J�]�����>9oEoPѽ׵Ր��%�T�=�"��h�5��Al�d���Uu)�sw�w7A�:9u]H��$��F��<M��7�����m���ۑ�#��p��YI�MVs�l�r�Y|4o�b�*=ٴ�uV�*��F�H��OQ]ӎ���,�z���Y��3n��}��ރ'��V{)��Av���xGL�o��PoRkG|��)e��3M��V�L�t�X
i캹�V��K8zs%g�w���jSC+��i�g��fG^�&3\9Et�y<����G�~���RŠ�\��z5�ܢÖn�*�l��v؆<
��q��$Y�XI�%N��M���.���Y��G�WN"�2ˮ=���*WQv��Q��$������c`��6Iu�i������H�vK9�WZd�#�F�+4����IՎ��ή�"!���KUi�,�.Na�Y�ي�ө��]f�!�z�$NmY]���7���뛻���s���u�� e$�\m�48������ڽ��KxD1S�\h
�2���¸�L���R���Ɲ
��7�`�ǆA$wr�8�I`��{)�QZ���ȹ�m�WpRp���.�X�o<����Il��m%W�M��Ͷ>���Eάd��]�K�N�#���g��*{�Q�M�Q_p(f�\�v8{7�d&
��;�����	ŝ�2;���7F�u����)c���/���X��oo���Wو|�n��s��@VY��n8�!�{V|�P���ݛ�w�p|w!�������j�LPIvwN�Wu�*��d
�K2� �[ɝ���E��S�M�6�؜��7��L��d�u1�N��xpd+���n��+�}����ܡ�����f����LX�����u_dD�u��5����*%��޲�kR�(��N@�ZWc�,ڒ�u+�}�j��}��9����f��Z1]�i�ԅw;z�|!I�m���lv�{��YۖBu���O뻬g֏-��Dűm�Tj��:���l�L�q^[�ZI>��>/]^���{t2��ƪʞKE,�j� c8(l/"L�uuѺ\��e�.�� �s��k7z=n�+���`�',��k�_u��yjhm�i�3K\E��[�mΥ���]�
��:�����}T�[�{��v	b�C�!b�et��
c��C��k����-�V^m*��0;���[{YO�����	�;Ƕv���S�K���@q-%��i{`����i4-%#ЇMwd�Ꞟ;4�D���5ҽv�u]Qv��Ph��$�К%$B��H�È������t���@�Rm�1D�WCGGK�4�4: ���Hf�����ցӤ4�mu�ih������)Kj&�A����P� ևEh�����8�$��MC�:�	CMI�-)B�����)���֎��]#��]:B�m�M=�(��R�I�֗E�lGCK���"{�����j�zh�z�����HuAlPkn�E!I���i:Ovx�֋N�ht:R*�5T�{�����y��y�op��M]�І�j�`x��5:�Ƥ�o%�����Ἶ]=}v�l�+UE�+���J;����>�>��`��
������=o�\C��=��_�����{��������������������C��t��2A�~oU?������>�����z����Ʒ��;`�{���y�\��FLFL��������O���ןd=O������������y<�������*���>G�y{~��<�Hk�=���`������v���|� ����~�P�C���7�84Œ�>�W�gJ����"���}�AO��=/�����4u�ߛ��?e�z����Iw'_�d:?�9���u�C~�4��ߙ��j���~���`����仹[F��c$TI�W��yOz$}�������������~���?c��%Rz���������t�$������=K�O�������_|�ʞ�C���A�������oR���"D���]�1�G��*s����c��������ܾ]R�?�u�O�:�����}�_�z�ϭ�P������>��|�!+���D?������/��
�}�{���!���~ϐtD�9͖�M�����w�\�G�C�?��};������?_9�S�������~ǒ�~�?cA�����'C�~K��Ǟ�Ht!޿�}I���J}�ܽ�T;�� D��P��Q�r��ahHY�d)��ޗ?T� EU ��_TE1UPQ|�l���|��>�����*��=�y���������S��/A�����4u��3@|�'�7��u�C����'�|�t��}~{��>��{G��o>��}��"DH��ޅ�>������x'�!O�|����z�	�$�}���u�^C��Ͽ��)�����O���p�O�����4>��|��������it�������w���v��#����������C�~���k��/y��=�G����@S�.���G���R�w�<�A��#������~ï��~}�����@x}�"p��C芦�(�zu�/�x[������>�#�}#ч���q� 4ih�i�~���~|�PcT$������P�� ����T�å�}�ߑ��_��/~y��(��w���̽A��`_�{1��s�U���v�,��%c����vѲ1$Oi���^u��0]�I�j�4��	�ޢ��\��Gz{�-�2R�u�6�v8�3LL���+�H�&fv��Z�y��uw 0u<��o�3s�;CΊ�T\���x�:5�y���heqw{f�NA���.uOr.�Z�N�g���%�U�U�U���<�~�/!+�����۪}'�^���~~��z��������A�<��5�~�����>O�~|���~ǸJ_���G�!���|��4����">�n�t�x�L�U>�����*�o��p���|?=r�_�=�d�A��N����B|�����Ҿ���>H�~��`����z�>_�|��z��W�>�U��M�5'=b���|��>�"D} y��!�����r�����{>����it�>~z��~���G��'��!�z=� ��k�>��~�����������
}K���>��z���\#��q�6lr����V�+U��B>�B���=�{��h<�_w����z�������%���=��"��uBW�
��q�?`��A��d�y?������~A����>���k�߿�h��
���>���.��>� ��������A�}��?ߜ{���w�Ͼ�	��i��~x���	�|��w:O���_|���.�˪��z�<���߸���J�~{���>I�<����nz�g�_�9���?`�c��za��P������A����_$�S��{���y�=}����}�|�>�����h��o�<���ϙ��������{�����AG�������qr.M�v7�fێ�����<uz����k�^�'��O��=�c�?��%? �y���?c�:C�?cC������K�:�������K��������C�#~w�O�|�O���^���#��vd�O�t�:+��>b ���M�C�>�����P��^���~G����饡����~��=_�~��_����!+���>K��^�G�~?p�?/=}���	]��=������~
���qg;��j��B"DDh��.���'��^4z��O��<ϐ�4�o/]��<��>�y>G�}�_���'�#A���}�h~������Ht�;}���
�����<����,\�� �}�����ߔ%	^�}r|��P�����ɯP|��:_g�w��	g�����߁��Дz}�r~O�:<���~d��
�>A��Ǩ����c�K�"�>��Ö��N�o�(瀀�c,l�9o2z(�T��`�iwy�:�����]�>�9��f�mH�e�!�Y����I�(�ͺߓ�x͔���jK\�+��M�2pr�Ww��A����т�I��J���ݎ�wu3����u�C��I����_�y�����c���|����x~y�}��MRz|�����d=����!���'��~���������������:_����G�"=XQ�s�4ͬ���-�_�|����=����O�t��_a�[�]:��;�����������=C�����EO�}��$��:>K�u�w!C�~O���،>�"!���},���C֑5�ڮ����ޱ�����.�����o�|�����L�M�'�a�Lɋ�p8d���y+�(e6��Kd�e�͹�n��Jf}|�yh�3�n�a�򡕋��W��=����1og��K-K��:>��D���:NO�}���|���cC�+i %G"��7"gc9R�An�֌���A�
7=�CD����'�r*�6d!�����Xa-h⨴5����yW�*�#]�}�5�S�H�.%�>ӊ��\WfU/�o�Ї�3��wУ��������ϯ̇��π�V�?*��4�a.��sZ�u
�b�o-�ԧn��T��-�c��BrDM+v�A�t�����yy��$ﯾ#/�wَ����mp�RZ,QV
uq���W�b�S�i���uˢ�Ĝ�	}�k�V�{|(5�j��t�g׼٧�������u�>�_e*6Z�\���y
y��ܮA\�Kz���&��Q��]Mc����6]������V �	]���n]v�Ԯ�\��@�&�U��{!��շkK`�xwu����o9�����M��+ͱqc�6��g�s����{N�;<mP޹O"�<��4�7�@�?C�2����KGu�H���@�50V,��,^����P`��4�j�r�$	�m�q�2��(�SR)V��K��}���^g�W
}��j5�İ���2�}4��(��X�8����~LW��~����ˉ���J��2BP,]�6��ޕ��&>paLk�F����ܧ@B �������3�|�G'84BZ$�s�{O���~�;�Q�ƙ��O��P���0�n&Y�ULU�T5S�y�=W�#۬|s��H�U�g��#0�F3�����W�j��ח����C�+��r��znO4�G��&�U�Ե�{Y�Y���@����E��j|@�E�.��������R5�ԣ�.{���*��؝�^��Y���{zUǰχ /α�[l����x%$���r��|��+����ň�{0?�������:����<?:�j�U��m��č�L�K$E�|��~�G��4������"� $vs��k�ns:ySw�b�S���ծʊtU��ε�G�ݵ�|�����^{U��C��g���7h ����UvF���e�Yэ�Jr���.���̊7�P[��ڧ^�����A>����S2_"��Dʆ�	�sa�GS�8\>�<n������x��륺ϧ�⯍�i��݋%/rX~u{|�;�Ԙ�<_)�*�1����;�h
E ��e�-uӟ��{~�[o�V�`9�p�ɾ,^L�{?%Q���ۥ�a����W�s6�'bw)K.��t���֬h��������n�z�@�k|T��i�,{�����^Ӝ���gǨL��9v����SMݯ8Z�~
��KW]�~�gP�^��	�-�O�*�a���u������#wL���g�c���+����/``�ŋ���Մ�*��w�b��e��&ҝ����:ȐũZ�ptb��f�n �f`��vҰ��wD
��$KTB�ba�����UOv0�Z�-+{��)���X>��t�ߟ���d��;Ǒ����]�:�n�U�}S<2�\xL�3�<�����{=���>�{�]��k��k�j���|�z���ҀJ��w����lt�jV�\��Ԑ1\<J=wT�+��1T8X�u��+��C�s��`��Iܧ�eD��N�����{�s�%��:d���]�hSM�=��sŹS��__�l�Pe��{M�c_BS�Z�Bx�`��O7�\��L���}Ԓ�k,=�3�Y���#ְ��(��7�]�oP����8kF���������N7�}U����ڵܾ���n�
��MH��5<f�뿭T�]-W��倦�����Pxj\]�B��}4��;�t����2!���~�љx�����s�טT�3��m!��B�T��r���)i�<4��?c�g���.��P?�е�� 6���=��P&�u��q]�z��9l�f���3���X�AR�!��`��0g{�Â�z��"剠h�^�O|�'��b�����c�Q~�b����m\�Hpc��W{2}+ی閸��u�o�E򞓏l��z=X֫}ċK��Ū9��Y���̺z����:���{#���:ˮ�x�}�2���WC8|]���yOI`:�}��&�eTK��Ǵ���C�u�p�h~��\5�Or��1� �S��R��v/����p	�żg֗
�<'�qnn���j��Up�Tp�����Hh���d���x��(�ƞ����l��P̥Y��*`��vw<Ư���ʝ�P��{$ѿ��৖��;PB��BF����*�A	OFT�n]�KT�����Jq�:�e!����Zf��+I�@;;`)��4N�B�`!-a������Kk����o���LV^eby��e��f�r��3:���[@tԞU��f��3^6�w���E8��ԗ\0`� T��m^�oo5���h�'"�z�-�}�\��g�g1�Aά�(M}r�M�guB��|R1��ɶVC�B�z��<<���!�i5��깦��_T�P{�C��lU���%�l�Ю�U��x�Z�(���=�U���f�u���;����Z;��$�,N�H9��2�.�xW��OL:V6:IahX�[�ݡ���vW]����ܼP�[�t�5��Q��¼�p��u�q�Ȭr�'5��/��!&H	�Ǫ�f1�`���R�45�����xZ|��z�Wb�'��s��������� �%��@YV�?RXn"ja�;͒��/*��!ߙk�x�"��㘇�����*��W�����^5��]����HՏkר� �ƻ�y�g���^�����=�u�K��#\�Gª���v��TC�{�_˯nRe)�my�6��wK A^����>εV"��0�^Z�_ /�4=���W<*Y���h��^wsG{�ڭ��wD8Q���q�v�ǡA��~@W:ć	�v�>�^���,q���^��r�����������A���p��7}i>�ˮ�_d��d6�^�^GDjl5����A��VR��[�V>c��z�LZ��-/I��׳hq���5Mn;]m6k��gc�������<�Z�r˂lSx�v�w}G�.�����T1d�}���������{8=�Er"�ӝ^s����9�s�������u0����L�O��a�񬾏���9���������Q�v��1 }:y�w��Hsx��1�U^��p�~�a�g+��<�����=��Bq��Q������G�\��%&�Of��ݏ{���p�EZ��)!�����3����F�L&�<g�6�;k������m��}�����>�b���E�;>�vЯ0�~��&w*���zmt2 ���/��H¬�z�ڸ��B�������$c��b	E��W`������5�����iQ䐆;J�#����e��i�~��*�}��X��Z�tEz��t���]�6���`R�����K�)��7�r���`�����N�n��|��z-�x�<��K{�W�f�-���Ȃb�@�y�͛�r2C Fv��wNL�����x_�,�T��n�;o{ӄ s�y��V3~Y��҃�B����N	g>]T���0;X̿O� ]��xt�V�-��1c�]�D�E�d�"�+�fV�T�։Jq��a��o�
4m���P��o%���ym�l2]o,�xaά����t�OB�
b�R`����b�������ˮ�W��|�T�?p첨.� ��K��.�G6	��1.듳�B�D��|�(�`�=�\N�3���Vlu�<+3�N���Ҽ0�U������^�ۢ����\���qK�l��A^��-CEh�^y+�UZW��0a�|(�ظ+�f\�zKY�O_n�V�M����!㟬��lsY���d�c�{����Ga���z��o�K퍔j�1�o���e�S�j��U��+��Ùa|��z=;�IX��x��i���K�\�i�5�k�\�YY�� b���4��m9C���h�{Yf+V'f�b4��pJ�_{޶U߫�r�O�,?A�|v����
�W�$/�xw�t��$�-�xl8����˧�3q��[��b	6}J�y7�&8<?.��A|s�q�|b�AƉ8�Ȭ�/�ԛ�:���:��vM�踗vfT \k|T��q�㽫힕e����S���͗Wj��:�n������^����l�h;���փ�E��M��n�
=����(��ĩH�5<�h������C�O�5[ا�b�ye^y�M3�N��Ok7+�� ���I�K��`&+�9[D�!Vc�^���i��M�!���1�rˊ�]���\ԜUI���p�6Q���OU[��>�qHcгg\���wx��U�y;v]w��2	��h}���(��1$�����
�u(u ��o꯾��=�߳�2�q,?pR*��Wx��`��xS���_�^dJ�<x:�î�u��s��e<{����~��x��`��������fև�=���]�ϻ�uS�ѻ�Oޫ���^>���AWj}�:ऱ��6�Χ����=e�k
����@}̞.�s+k��MLd*�������0k@&ǥ����Z�t8X�x|-֦O#ʛ�p�X��RÓ����5�/�'(]�KA��CܡM�%V��k�׬�g,:�\<	P�K�Qwu���Z4p}2t�{Q�[$CWWΫ�A:�0ud^�^�u��}>��!]}F�wA�im�nk�kS�����B���U�n>�Ch�yT�R�X} v;2,.Զ�ay��y.���Q��p���c5\�T1,����B��y����Z-��Y�����]��1��k��D���aVNyV�!���k��f��PW9�B��7	�}:��G:V.������f0CF�e`=�쌬Uu�2����HV:�^-�|}��W�>
'�T����mU���u�1��H��Z�Wuʠ��}�S����y��uI��c��b�RǷ/zj��գ�'.�'�����L,�Mԍ��M��ɴ��򳺭��6�a��H�wx���v!Lu��F+;a���ƥ5��m�ްJ���(��8F��5ɢh��s��#w�/�O=�=��1fl0T�Vͥ�╈)�v� ŐG��R�A�﹁#�m�7��Y�K�ve�!��U�fGd.�Z����6�LnRPW4�^a�}��^پZ����
�&Q�HP&�|{�RgA4�]�;��Π�ۓ��	h]u�$�o��)ɾe�*���z�{,8:9��M[w���r��*�ׄ���j��l�#r�;�+]�[ي��8h*_�$[3*SΑ&1��=��}]|��Ee����Y]�m0(��o��QRJC
ˉ�{`�"�������>��Xo3q�	@.Lmap���u"�*��nS��L�K�C���W�{	��fQkc��Π�.sd��V�]%�������5N�n��ǯ5mZ�GT��*d|��x�s��c�.nw[cBm�|��U6�5x;! �Kbŏ�dp=�P�݁�j
�>��Z��)Rn��K�"ibr��}XyikF���e-�h����e�7n���ү�c{�;WK�)���T�YC6���v*��Z��]G�r�E.[u��Ե=1����\�"��V�m���\�M����Ӣ�\�u��ar�eamK���\T҅��02����q�׬��F��-6�z��i�!�[��u�ݸ��š-)
�.�F9��[��S5�q��x�����%�?:xN�#%5H�ˆ��u��ܵH��n�;9!��<�s�8�Q�ݗp�S��f��*����h�m����3Jz����=b�u>��xE���5�k`�5�[W�mDf��V�oj=P�2m�4Y*�mm�c���e/����9X�8{(����]"�IN�������c̒�ץ�ۊGW:�71��9��oht�bWm������(��4��WiVk}aH��QǬ�����{ܶAXjn;İ����R�_e-�rv0<˃���:���"�a�N������̦3-w��/��I�0� ��B��u 7���>�W��$nn�BpXd�9S�t\f�J�{��Ї e�L^�,ryE;��7Z�e\̵��d�9$�9z��GE��Jڧ.�.kD`*�r���n$*T*����9�3M��M�&�FӜe� Ř;{:��e�S��e�d�E�r�.��T;+5i�(T���R�����+�=A�qQ�{�����ݼ�U+1V<��'KC[�Р����z��s�n��e���������6�x���C%Cw)@/�%�ռj�C����N5�>�JU 9xۻ�i�K+o>��J�_soW�A���<QSᩒ�u`U�C��ig>�R_��M%�+[m����RPt�M:�щ�)�KN�PglD�f�v�:�E��V�En��(��%RP�6΃��Z���t(RݓTi4u�����;f�j������k �1�C�5k![`M�$M��E%:4:�˷v��lul1S8�j�Ҷ�q�(�����c������	���)N��%�Z�ĕ����CMض-d�l���];c�Ui�1S��U M݄��+C��`�'lLͷF���&�펇��"u�'mh{��NmI��gA��ER�.�Js��⚮�Ak߾��~z���*#��G�;栺_k�J��hV��&@VU�ы�8�[9�U��]�<�3m;���n�N�����֟磌�{϶{��t���}xfS5^�D��N<����,m�\K������d,�t����v���HA�����`��Y=�_)�sU]���t��l�4�����y��l�N%,ݱ�a^������hp��wP�t�Ep0�L��Nn|�����,�̞�v���YW7#Et�t}���LK�xX�_d�\�e�#��F���^�{lx��2�V���9��Z���WT 56#R<&�[��鄢v�#Dp�RW��m@�e�t3ӂՙ��;XM�``5��j��ˤ��=>�|g=�W�S2!�qj�w��f�:�3�˱�j��C;�;&U?1�RU����X^�+ʗ�d���,:�Rj^�ρC+�0�0�8�SݙL�nZ�λc;8�. ���$����)[7R>մ�u����Ɗ3O
� �xyi�⭱��(8��P�� �v�@�E:�<v�C=����?lYC{�����抵O����N��30��c":d�A�!�n����b��5����ê~��w	��ZV�w`o����y�U��:�o���ɧ��k>�#;Z��V��7[k��-�ꖷ���Ԫ*q[�p��^�]�lH"��t�0f�wll7ڬV���o:�gl��u��\���Y�"�mm��+�ܨI�����E쓧���WՓ];��|f0w�]�znrp&L����.a�WMb gȰY��B)7��⼞<c�ߧ�=~��]�$kG������Bj��i�7T���	��|�&QIغ��/��]���q�r�}�Y�戫�΀�y�>Yj�uW��[R�R (s��MqP�����BI��Ρ�5u�^�'X9g+(�Yne�"(V監��2����_���(Ԅ��^�=���LCD�g����.�?Y���g�=�-��e��v}�>�;�R����b�yc�n_	��/���v�_L�"�M
�<�j�A����	���[ J)�u"���pժ}�_��Z@z>�+�����~���+�Qa��%=u���֪c����0?Ls|�����h���=���IxX�G�8{��1A���������F��v�]	�&�cV����}ջ�~���ѧ�:uW�Ӌ�����q{��/�W�ذ8����f�+�e̞���W{.��������E�86�#�Yk���A��'�9�t�Nj��n�ۛ��U���>��qu�3�L�(,��͜T�z�"�^]Z��\�#}�fUِ8�, dڈ��ݭ���̳ˉ�`�Nʾd�QН3
�XI҇3_(�wn:��]:﹧6���n�	��w�]o.U�
���գ��k�������Mf����������0��[YX<j��r�-6F�F�U?v݉���H�lۊ)��9�b��W
_{���m���*X�`N�ֱ܁A��������W���<y��4\a�L��\@Ϸ�oó)�̮���h>�ڼ�UӮD� |���)~1��O��dB��as��h�����`�G77(eR���OGʯ���2�T��r�8O-�o���ce�EL�T�)·z�e��t��d;�Ѐ3�qm?#Ki�:{�k������lft}���ߺyJ/������\�1�<��Xc�瞗����0v��EO�v��8��{��Oo���W�Y�y�{U<�dx�s�]�^��4З��ώ�ܴ��Oiz�>C�R�ʧ/�)'��ke匨��r������:U�'p�{��׏�{��!{H��||%>pmd��Z�����F}���S�7Ή��ś�U���^T|=��y\��I����J�,�R�+Z[Q�.��$b�w&���fZх�9���G`}�26/:�!F�ٱvY"��wQ�[4Q�Sʝ:��+��X�\��]eݠ{T�ozqV�0������:ֿ�}U�W��[�-=\հw�t�q��Y����ضOWc>�dqҰ�b8����������~^���1�����iQ��=��E�]�����|�[����q'	�����X\��Qy3ts�+��ru&vz3�S��&�����I9����-샽�����}��Vz��&8I����jVys�OU�`�z�߂�������v&��P�4�?��g�h7Jr���Gf�Q�M��¶��s�z�����㫽��}�����&WW����7�5���΃}f��:�s��(3Y��<��=Z��m<��o�.Իs��Î�F8��|����G��_(,uM���W=��E�J6�b���T�K`����j��q�5B����§�贃�N2�j^"��a]����^ld�#2�p�t�7�J��.�1�
�����_n��X}�JƩc�.�W�@u]�piou�����[2:�-�E��K���%J��e-�[��j��c,��b vY�}V��^��G���c��
a:U���%vm��F������
�i~�"#舒�0\ܮ���4�P�y��`�l~ߣ�����W+��p�@�J�WS��6{�6���u7�>�A�}['?�������/�d��I���'Z�P�S>�9G��^=G��c�_P��ʝ���ܥe
ys̨�rp.�z+���8՝��m|d ��>��1�_��4��9e�����?t�I��s�����=�T�Ч7��67�=wW[�3[De6ط�\c���nCNZ�u���w��S�WmҔi{+s\�qn7����\�:��5��ܸmmAt�~X�eB��{ۅ֯s6z-�����㾼ޏh����{J>ڣ:��;���m�a����p��y�nu���ſȚ�ރO�}�\���y<��F��3x�NK���:�?�`T85_!O���<|��=����G�孉\�u˃��|�+ ��������9KD<mD����\7r��ju�]=�+¢$�e�C�^Ia�|�y7;m^#���7q�ң�TR��\Is����GZ���'�r���Ĺ�n�r�@�xZ�l��j��`g�*luovT��������4���e����Z�t
�!Y�ە�[�ũ:��w�����KP6�=A�����ۚ3�ktk�9<�;�����6c�gVd��`�b)��8e�b�y�	<3��9�n�!ky�:��hL[V�=���9[�u,�y@ϼ�~�+	w��B���B-�W0�Q�ڱ��Ε~��Jz1c3�n2o*.�W��3�(;/�UVr���س�A��Q�I��c�$/����
:�N<�z��ʈǎ�T��UD��]����`����n8�c[�r���\�O��}s������.��y��,�|��0u���Ok���<V��{S��hy+��g+���}�le9J{}�TMOsf��xyo��ӌ�'�;Y<��FCSo�W����=��W��L<a�3������!%F��˔�jkr�����\uCY��1[�M
~��W���ާ�6�TC/�;���Ք]x�:o��a�`��:����Ȕ;�Le�u����+5�#k����um xG�b�ƶ����Э���H]q����x޵ݥ�t�om���7q1��DL�AbK;,Z��Z�J(�O磌���(��ޞ{ڻ6��z*ӳ���Y&���:)Uܲ�8������}sn9��+�U�U�΀/���w~�[SfUk�[Gg��{���8ީ�=�=�9�N��|'w>�M3ؗ��W6�ɼ%s>�[T-���tڢ�Y[u�;��k�槕ޔ�����J�e��(�uN{#�9"/>-��
]�EEa����};�j���q��vj�؉�HD�`���b�-���䷔�j�^v��]�w��d�&��N�R����m�Dk�tGP�{qJ)�����l���on��:B��3�9��yï���
�S�Н��l��|���z5�3����%�ʙ}�_���^ҹ�s�h�j��nʢR�K�^8q)�$҇�K�7y�>{�>v3�����9��ڜ�/=�����ƪrY&Z��5��N���^��B�Z�)���M��@H_l��:\�(�[ĭQ0�#ֶ{�;��������}%Y���jz�!7�d���j�y�+;��f]��S��f��ζ�`�6w�Ӧ�c�D3�[��m!ssi���@ѷ���4y��~��X�we�/���6`+��X��ݫ����][޻X�N�I�9v��m�^�;�6��{o��4t�_�5���w�n��x.�Nq�^�Ա�
��ow��+7�[ڞA�C�Oa��Vr[�gzm�~�-C~!r��<v�Prxm.>}�3ף,�hz��L��w����=Ӧ@���j�Q�!|B�=8��Kٔ�x��)U3rLH�lkm�k��&��%"��S�׵Vo���#����ۺR��f�ܻ|�ܫ���Anѿ�%ozÂTG窳��*ߎ�oǺ#��P
^�;��M�؊(�ܹM�-��]趏��t�	t	0���ӝ�w����@��u��D6��q���wO�y����1�M:M�*,.Xc��T��I<���Y�M7���k��U�F���]����O��P��N�Ҟ6�8��P�I��\�Vܢ���F�|���:���j痟��o�I�<!-�ԸWYpi� �R�v�Vs����G�6�Wm�0�09 #�(�\�xSx�bn�zw�˴&�e������zJX2�h�;XGD�[��Q�x.�j�l�v��%&�ڀ�o�m�1o1�K9�x�?�T}D}fp5J;��#�F�0�>�u��k4��{͛���������a\�H�.%���&��K�P���]3���]��g������|�����}4�f��
�n�q�%8Lqm��O�ղ]R���W��R�U���Ox޺7|$q��c�=�=��>~��U�Ư�v� g��{���{�|�� ��N9{��jt[Y�m�&���-�QKYu�p�'�^��l�^�~w�=�k�돯��{�諗�NH�H�ߗ�y�A�>/��_/mU��3C�H������ܺ�R��=T?v��>��H�]G�[�Ꝟ:e�_�8m�/ztd����W5o^`�/0r�J�O}gE��_F����E�/��0�O!�"�k���/O��6���=����0�' µ�Qg�ald9���� �j��O�[��SϗnB���;�����u�+����A//#G�7�\Չ�֚��ؠ�ѥ/�L�;�k�N��Ȋٞҝ�ʸ{�YR�M	l����.f:#1�8&�:�s`]o\51���-U�����+��(q���so����:c�=%3�=����T��䳽Sa��R��EU����MY��&���a+
�A��w��_UU}^����x�qW�k�D{�i�v��iw�?{�n�շ���i�}ԓ��UT��Wܷ����7��U�g���G{>q�)K�&��=��찰�LvB�vՉ�n�y\�N���>D��@}�Qo�����r����5�pO�5�}�'3Z�!���!�&9"/~r�����	���3-gC�=�n��%sҵ?���8]�R(Ҟ�r��N�Z�ya7�K��u��&�V"�C˽���Ԯ��!��9�o�'pf�0�� N���ʃ}�q�5
��H%K����W1��<�|yè�j%�d��>�vHQX��j�!�.G��G��ӏϱ9�
x�0��u�AtYF^��5=&������#������XW�#�����|���=��������˰]�`��]��}÷�zh�}�ȬO�#�Wy���	�R��Aǜ�`Ʉ5<<.�X�}yÃ�qv�d ^�YE}��z3I)v�Kh-�"˸�v��\rD���۽v&ʍ��8/f���l�����2���&[q����J�+6d�9��5L�Ub��rk��q�N����X�AsX�w�C��̦h�@�|��]:T���	��ǝg%+[���dvF�Jĥu�\5�����R�s�h�G{y�(<�%A�ӫ2��d��b�v�	J�Ļ�6R���%M�d$��+j�%�Kz��\�_%��}�#+V��+!hwVrI�)-�)�ٮ���	���eF9����o;XKy�sch��]����s(��G��Ʃt�]-�ײ�;�A{v@0��%2�-�b�7@�64�v���w�(��:O��<Yx�s�]�w���N��φ h��!%v�}$o>wdt�H|Kj��ˮOn]���W�is�|�U�oD]�T���]�y���QAN�ь�WӮJ�hf�!���{�%fNJ�*��`)���Y$s5�g7��q�t���#r�E1���a7��n���_$������wݠt�\:�lN���>-Nn�Nt�s,�r�C��Ԏa����+ݬ��O��I6�m.�,.��`��NcΩ��Z6	���3�V�r{�f����Q�N��n�\��j���`X�:�_*�3���V���--r轂_���d6\��[�m��̢],���n�K���43��[	ݕ�L��*ۏk`ޠ��q�@�t�"��Vu0M[�D��{OI��-6CyJ�LʾR���<�B(df�6��KF6��U��u� 0�t�:��;��S�50�}�kib4�����uٚ�v2h6�˥k���R����/�P���8�"��' -��5���:�W0�ଷ��>��R�ҹ]COp�jES`C���87cC��˥f�*����{@i����K��(�b��`Y�A�T�v�k%�۴9L=ַT�i�!�:hS���U���B�5�Ŷy�n_-�R<o�U��}yۨ�E4��Q:���KW*���}Ý��SV�k��y��˭��, R�X�l2*m�P��oAdN� �^RZ��q�M5���J�fe���I	pқ8B�
Ss8��o[Y�ۣ�؋7�BZ˫��a����c�I+Cg�_�k�+�=�x�c��:�W.����iJW��Nŝ�U��q�h#GJ��;v��&�y��c�%0QggB^g��>�5:.�=ה(ۂ��Ү�e]�bv���X�J��(m +�ڡ�mΝu��6��YK~���Ln�N�^���
Z�kS�ma;�V������k��[G���^7��S/�Ҋ��y5�,�d�PmanL��vtX>����M�sn����v4)?�/��BQ��=�{������h)���]t�%�]����Z��J+Z��)5�DQk-����i�E���C�4[h���Z-d��CF��jB��KkQK3DQ5�5��ZK`�a��`��(�b
h.�"`��z�֪�h�0���M=�t��F�m���tf`��F�la�� ��Uj�&-�cTUQ�6؍b�ABUQDQ:�uF�Z,`�4Q�C�
m��Dh4m��7Y:
��&*" �k���1F�эU��ִ:���"�����E:�6Ɗ6h�[j�����)���UQET@l#M�T�5Q[hѦ$�&jt�P��@�B��������^��f�r��sib��ނ�
ۓ.ƹ��A�X��2�:��v>ưq꬧��&�Iٹ!3ظ\�U�}�}@�f1��w�:�?C\]F5�7*Z��9�:n�֫��Q�(�$ԯ�{��c�U���s�t��O��s�4��rûq�x�{/Ur׀��/:�������^�G�Jsi�-~�:p���y�5^��!�hrW;��7�o"3r{z{Nv���krlb�����_k���J��Mj����@��b��kw�e�i�uq4�V���Dt��������������_vQ���Z��Cž�>��>�����_*9<7��Q�v�ޓ�Sw��	$�Inm�뛦��t�_q���0r�eCޓj�>U�w�>���7Nd�J����9[I��|ֵx�&)�4ܲ�`J��,�2����Վ�%�M�w�O3����ޕ��OÞ�P�@��G�L7��0��Yi]�rFؿyw�8}����O�;�
�#^����ѯ�qԝ��R��[�}r*Y�[��;6_J� >�}ݓ�Ү��,���^��eG3=��3��;���{�d�\һYq�׊��r�А���5���6��ܥYC';�!>֫GF;�pu���i�N��3�p��#׃�-+�����˺�ՠ�����ݷѮ���������d�==�-����o*�噧�l�����1W�{(wz��폒���ؽK�̣'��\�(��q�w��F,sQ�'#�q�v�ݒNEw�tU��k�P�K��W����7ȬK�>z��ʥ޵��P���3���r�KF���L�A���p�^��Ts��E����9��I�j:�7�m�Ẻ��J�R�6⾎�}�R�C}�v���.U�����:�.��\��g��T�|�K��K'P��V�v��x�ڤ��T���q�e��n �rWOޛ�}�-��{X�!{WR�<�R���j�|��J�������g�u�ַ��5�j�N`�C&-+5��V,��\��a d�2�����ic���j�Wr}��t;+������DN�#��=�+��02e$N���{��C��jl�l�_3]������jj����N�ޜ��v�d� ��k'LYI�D|��צ��Ӫ��:������q����_����c4U�:g���!s�mAcd=�l�x�;J�&�uu���۵sj��|Nr�V�jxK`X�j+�E�Offuwsx�����Ǎ9p�V�|��X�{��j�f�{X;p��)$�ﾏ���3���P��N%)gn�S��ڂ麸鄩��áe}�<��05b��+T8�O6�a��5�U��݋ZQ�2i�VͲ�Y[0�Ԅ���G��s�P��*���Y�����5)k���þ�>7���ٞF�Q�$��e���s��C=�M�EwC����3k]�ϐ��^�M��9�O�J�yA~��
�g����f�i�¬�p����l�{orO5��Js��q��r�S/��>*��{IC>K�O՛՝{ �-����B����A�n����*T@2���Y���*�g�;ZW�Ŷ��Jc��qV8.��v�>�L�nؽ�N�n�s��� �^�¸�8���X��{��.����BywM��Oq@�;�n�ؕ�ޝp��W��#���j�ŵ��^�}CWR���=��mQ����4��y�*�MxV���y�fx�8ﺕ�� �c�:�=5�\5U�5�l�}�1g8� BA��>�ۂ���a��M�*�#K��R��}�[dV�'H��p����]��d�v�������ێ{ީ:���]����[f�QP��Ϗ��kƺ�;�M��G����I଀�?�'x�5g�F����Ò�{l�r�םQ�N<���(v��U���w�}By�s���*]�wڟ`�*��p�"abɺ��p̗|�#o�OP�nӻr�K��������]]�ʖ�5�oy�y���t
W�˕mQ��#���U����m�R��m���u5�@�-z>�{=^���n+~4���ߏtߎ����h���vM����_�Oakۣ���N�ϨWr�r�ey�뒃�5�T^ꯋݝ*��2�+��"��F�R�k�YV05�9eɶ]��Z�̀�03��p��w:��.ޫɆ�ru�L�j�=���Pb�:ԫTf�ֱ['c�k�uj�1�wV�}g�hm	��5��¶e�߼6y�E�7#��{��U������/F��^�2�]*J �T�/G%��XY�f>���r	i��T�47��7�:,{�M���u��
��p����w��w��s7�w�N�3-M]R��b���*jO`�u���������Y��G9h�z�,����޸��F�r��_����ﾋ<�=r�ޱ��vL�	cۀ�c�)�bg��;��	��[vI@�i�g�҈�μc]ܩ���8�rp�Ӌ�N~�
x�0�����j��؇@Q))ݳ�9�vU�_�j�����̬�w��z�-��B���Lc./��a���3C��=xg#�!8z�0�Ho�8�y��r]�;|+���?t�J�����=E�c�5��5�r�ȼ�:N�k�:�
!=mzW�8�$��:*�|�&!�1Ι�I꿚���7���77�m��(
�3�\έ3ϵ����R�s��>��\�D������T[�+{��+Az��ͯr�D/i�i���SæO���vH�[=�z,�;��us�R�����Ī�k&c>��*�q���{����+{�l�Bnߖ�=�U�k�
��{��������Y������Q��p��=9p�f��>�&*�)V�k��xw�gK���Q��ޞ�X÷Հ��c��YG�s��.�F��}@�Z��F�j[���ǰ�h�xZ����g�J��:��OTǳO\GF]�ŵ�i2k#���}�W�C�y�V�-K�ͽ��P庎:�	tC*�uNQՑ_].*;���[�|�V;9�K���ݘ�c��(�m�4)����w*���:��y�+Mv�+�'��1���m%[�(��52~���2��>ԭRz:���O	��$�~~���pt;�6��2��s�5;�r�O��Հ�b�z�j���z�N�d�tZ�,����o�\���t�x���I�2������m�|�y?�c)r�k�ʏGv�9��g�./�=����t�z���e�}���<��s�ՠ���8Y�b�u(p]��WW��q/m�z�C�$��ʂ���M⚀�ެ5.^>c��w�*!s�Z��y��qխ:����'/��A�H�3�����>u���sGy�|Qū�{_RʝG�8�I�דOpkl[8F⼋�8'�ѡ��Rx{����ޥ�Rӄ�^���QS5��땚�I�[廂� ���GPL\v��uE���(f�q[���sd ����wM�s���2�$+Z��뫥j�mg,e�=sWW��o�RT�u*,��C�op,�II�uT���e�)A}[�c�|�f53y����}�}�E��w�������m�����/o˩s��V}]<2���������_�Ei�&����W{�񤯻k�������F���=9�&���䳆���eO<�N�I�՞^���q��P��{���}�`�c�ҏ�&�+P�7t>ɓ�\v.k��Nj]��c���]qBʎ����;�b2	���D�2�SK�ތ�{MV��O��ڂ��+�`I�#I�/O66��!|�A���]=AE[G{¾�����}Ϻ�W7�/a�T�ە�m��{۾�V�?Noy�3�\LY�}	��<&J���oW��tW��%{[gf�7����=X}����.[�Q�fe_y��N����=}��Ѩ��:,�������b~j���ByQ66b�!���6j��2ڿ&�`���
{�G=R�=��:����T�q��gV�Д�u���z�4ph�OdI���6
�\�r���6��k�:W�L�V����7��p=ې����/ݬV.�e�4�:P����X�ܝ���fԹ�tA|�D�Z�u4r�Z��,�b]���>��������>�ܟ����=-�7�o$�����E�7��mq�����+'�`��czc��q~X�nq���>�N�i`S���x�r����R��9�XW�#����b���I��v�������2?.�'q���us!��ߎ�)u/k�:����0j^�~�䫫�Y�{���|���F��w+l�QP�v���~(�]G��y���vY��g6�,}S]z{X�k���y�-�ܕ�hy+��l�.9�g|��Sb�{2kW�^���u1��O����;zĪ�M��u����@�����4�w�׋���P�}+v�����Ѯ=������R��.y�ן3�����瓯d<����5VUoE[��;	>�J��]���6��Rp��*v7(�c{��X�==~������o�/��=��/�oT|����-���>����e�3y�A�_�$t-�2o�:��O{7�����vW��8���
6���ں��g��)M��_�CF�x��ޓ�I���p�g�YD�-K�i������ML�i6�7S�zH�����]Ϻ�}��y|�"�}�ޗ���w�����彩�����|��&�.��~�}�HJ��UȚ��4���S�*�I��'N����s[�cgP뎇.P?{��ԯ������{<��=��N�s����e����J]����^�y[rp�݈�HD�`�y��0]ˌպ)�η]�<�y��w1�>퓑i�PS�_>�����	U<VGf>D_U͍�Y��)�I�^�3���Đ2r��2�*��o�|��Ϋ�����]T�^���A�{�=V�O�Xk��]�GVx�s�Y]Lt��O�ꒇ�vvt<�W�Q���l��o�Ǖ��z�(1�ݷ�}yQ�7+ᐾkh��Yo���z��c�4�>?#�w��\=�^�����f�v��J����ƭx���yR��td��,1����V��=���'���E��)��������ҽ�f��{9��W+e����~g�X,�.j�N qu:�PD�'�t��udL���P�O��.�*�ʘ�/-��WBzƙ`��)���)�k*�<WB�;Kw�S|o��O9�����:��y��+�O\�|{���>�Mᗉ�t8k�X�VVC���9��꯾���R��T������d�E�U��}����Q�O]��ڇ�OUf}���2��z�-������<�mQ�~ҕF��|�o�V��"^�W�d�"ε�[�R҇Զ%QW���dSYu���Տ��g86�4H��s��w��v��-�����>�x׫������;<6�tq��9�{m�X�E~����wmS�v�c��N������*�T=�7�VA��Sܽ��"FriL�b�W��^�:��E��ܵ�q{N��n���*s�|`����ܾ]/��nH�����n���U���(j��(�H+���!����u����I�£g�V�g"o�w
��z� ��Ѩ)�,2��i]a5�WN��W����U?m��U��8���3~=����&_eS�N���x&.�}r{.�z�t���w
�+�j�>J����,b�����c��>�{�vem3�<�Shө�
�.�a��� G�Uh�Ԗ[�]�o)��;�񍋫q��)+�ҩ�;V�4)�h�"���f�����i��Y��%#��31��nZJM�T2�t�;�&fl��71Z�t0`xr������ַ��F��C�r��L�ZU���8�.��͔xh����j�7�פ(�X����;_]�F{��(��a񢬅��[;��PP�����3��T*�D-F��i�ld��I(0go+oA�(foQS���]ʗ.kz�uʏ��	�ͮ2���vgY�^	E����h�Wi
� ����k8��u��r��1�q�\��t���ս4֎Nue1C��NM�(ۗ.�|�ږخ�Es���Cw"k)ᠺ ���N����v'qJ����a��2VJ�N�����oW 1��n����]�tP�W1���ٺ��0���J]ǐ�f��yb3�ȕr�r�^e�����ufp��9A@�#�t��gYoE�-�/�;�r�G�ej�����!>�l�oh�9>�-�d�g�(uJb�D��W]�t
��x��)n�9�K[��$�pY`i�*,���ǌj�Z�4���9��E�/)4$�Yy,�yq#С����\��NtC�*A-T`c��(:@M[��!�����4b����^���[-}YC6(t�^�l��4k�r�������[��2�B�Z�n��m���`J��ݺB'��r�U]0�c��S��`������u���J��������IZ���}Σ8 i�V��:���5���)����F�<o�GH0^'҅!��"� ���V�?p��Iciph��s�%Zx�ъ��ҕ�x��²�`;�d���uGC-턏 �{I�Puàv�gRcMd���F�I�0Qy���i�q�gS��_r�}��9�V��;�`hh=O����3�_7y���L:�fV����u�R�����H�x���Ů�t) ���)�O��S���.8���/PIRx�Ήj�R�5��J�5mA�,�c]msF�J�\r�8��'2���3���m�qrn���m�e��CF�5��|��{e8�b��+�b���j���[B�M`�;��ic�A�_
�/rP����U��܀��v�S��(��)�C�����>��wJ�.�;��6�S[�	Ò�R��6ٙ6�Yw3$�o޾��)Q�]�0�5��
���xg�����9���=DH������J�N��	�V f��Uzr��f�.��巘��{��k�4X���X�'��W0�9���B������-%v���T�ĝ��5J���0].�4�۵���7�ɗHb�p�AQ�!^r��  r�|ɔ6Վ����y����U����m1���7c{���`�J�[���'�g:f�]�@k&ck���;$��ԩ���S+f��H�J��}��wJ�U<4�*ujN�u/��c0��4���ӫ�(X�)�Z��֙)bJ���Qu���*����h�(�h�&b4b��M��(�&���F�V������EUm��(��g`�UMQT�Qm��c�آ��AA��M�b�h��ѧl�`���T�AUD���%k3M$�.�Z�D�
�lTh�4�%�1Z�DDM��(�"(љb&�ڱ��mEZ�Av�Ӷ�U;��)"�����
#V5EED5�DUTV٢�L�AA2vuX��M�E�*�PS51v�*����f�Z$��cX)#mIV�DAlj���&	�kTh��"�-�j���"�T3D5�EQ�(�����qc�T�,ME5F�D��M5DED�l��������q6�]����c:���]Fj�g�G~[F>:s�6ڹ%ŽzU�qD���;�
�nWgQ��_�U�W�o5O7ιn��G;�O�%�[�g�^����Eb\~�|ׯ�;E�{e���w	��s�:���U�&2����uO��?4;(�y��\�{�e�S0uuVJ���J�ko'x���\�n^��|=�ܞ-��@֬�g>���E��ˋ�:f�(���^�Բ��^~��w���햸fىI��x��݃,�y2%v���Ɛ���v�ǖ��5[��"��;F�dϷ��z����|����������&n�k�����=I�g�C7|F{�:ū�wuG��(=Y=(��\��gp�������C~"t�����.��{�쉉}I8S9�ϴ���V�\��am&%T)�[�p7�p�}'y�i�fC��Qe����iw\G&������s��7z����f������[�|=ʎw��>��l�����5~�T����������myW��f�m_k�諜K��	�9�b��(S����u^����W��� �o
��jX�Q�M�]D���`̷Ӏ�j��;U�V�lP;Α������Ư�`��f�b��#��:�wK�";���W�e� �ŝ���e,�:ۡ[�"+���=}�DM�����2oÇ:���NT��t�̔#\�~W��މ��ޏ'Y@E�c�gF!���y��B	�½څw3Kieo���蒾�o���$��+ۻ�����U	8U�LR�c�]��=�b�S�e?�w���D���.}�j�t*�օ1	�MB�s
S�q�Jp"�+ܨ�}�K�}�־y���x9T�׵4U-��{�kVLt�?G12�s������q��^�u�?Y�ro�����o�[3���OHu�������6�I�=�ސ�8���IVd�^m�b����10f#��R����i�	�J-]8�����WDDuE��~G��h)u/>��Ρ�x����d��(�J�s�!�k��Vz3�L4��ύ��\�U<���N����$g��{#���eYV�1�����\s�{cuf�-+���{r��yNap�]Y]vhT.�F�֪쮺�d�<�S�研U�����.�C��o���3�c�M�S	� >�.W3ݜ��v��U�Z�;;�iu��7	8�v�s�%���>��2�����
�jԢ�q_;V,��o7��p�B��?}U��ff�jx�添|�oV���yr5���x�>o5,�)9L'����8�T�8:Ƿ����E�Ues�ҕ}���.�I���e����ᨼ�F���/y�o$�S����D�Y<�,��6��]u�kmm��I{�+�9��D����HJ�Wey��~&�W-�nM��V���{������Mgp��]��-eT�6���8�*Ŏ�gk�}�gGK��Ov�)@���噗�X�t5��_�%_>|�[��H�rʱ��ɘ�p7�B�wݻAI=7Kx�NѦy�ڤM���e6�h/vߕ�N:
���5�9�u�@�$�,ޣ�xS����u���4�'�s�>��F��8V�J�cuNAR�����Ќ�����vW��Tj�߰�T��5W���g�s��MF�D_1�;4G���:{9����~�ܕa����"�����GJ�=YDf�'����]�~��[��e��It4����D��;B�ݗ��p��>�]؉��[���5v_�i9�O��L�֩��s]��\��*��o�E�KΩ�^v(2�5Ѯ�r ����7���<�y
���TF�KP�j]u�!G��gW.�zW�}�?4
��{�կ�G�����(xS�~V
j��y�mR� �۞�������|�խ�����_795e��?��-�?#K�/���=���M��&�Q�앏�յmR�C}��2ey	n�a������-KU�޷'��_�b�u�2wTOح��k�e=����a�A�������E7���{��"���c�U���\�D���\8ڐ��%a���6�a�p�ef��W:&'d>ޘ{������^T�h���r�v����{��6/I~~T#�C�&m-�*ӳ������]�ӼVb8Ĺ�ίs����Gl��f�����g骳_*��bЬ9��0J���)ĭ���s�K��>��Ӎ�r���4����CW�8�p�� m������u��t���6��^8ɧH�rʱ�+��V	qW�%n_�s�	�}�Vv�����Gv��d��B�����7ϯ��r/Sn���d6��W;�_MMk}�I�mԗF$,�f7i�O=t)��Z��[�U
Z�B����j݄*s�����M<�֎���ְeb�g.�(�u�l���)8���U��V�aOG[�w*w�T�Ao.�R�����U�����+��O��Ӝ�n{�ym�ӷ��zV^���}9?�����7�I�/��,�W���N~��0/�~�'�zt�Gё�k��?l�?c��O,�=��_���kGE��>�������L�ծ���o�[vLt>�gV�ו�c9_}��/X�x�'�Y);���,��,t��A�t���pV�e����ج�]%�_KD�Z�U{�/��3�%�.�8�u]k��;l��m��g� ���fOeS*OvL���5�H��]�5�
��lճQx��|�^���tj��5U#!-�C�ye�m{;��~(��Խ��N�=��I�C��0O�iڸ���	����T	P�{l��`���=�yo���k��J�+a�Z什7Llz��x��g��ߏ!��M����!v��<�����/��
"Y*支3q7�*�U�T#Q+��-���s����R��PB��E�('�3�o0�9��+=0>'�`�B�t�,�]-ᜄ�3'1��J��VE\�FU�s���bKu���#�2J���pT��Ӵ1J݅���=[:�]��� ��%�$%��{�u9ȳP��ch�+��:��a���
��+�`ݏ�8ž��[�������᧾���n||�n+N��wp-�Ī�R�k۸�2y:������y�旪��yE[���;�����Wuj}��c���t%������>Z������_��:���Ƒ���=�j�k��<�'ԽK�p�n�+���X�Q�:�Y��sj��+��׷�"oz<�R���g�����Su����"Es��E��Ҕy�j�jŕ?C��p-vd'�GZ�$7t�V=����\9u5�Cg�i«v&��!uC1�NϨ�������*��94w.ˍ3������D���:����S1]!�|L���^�/a攚����l�,s��.w3��u[B��d�������o��O�g���R�7;:r�=��Z8��窗 ����d��U*o�OJ�Ӄ��}`���z0^`��v�i�G�2_	�����{%���=%8Cͷ˖jB	W4Z���-I�v�������v�d����m�r����X��&��&ֻ�%��ܐ��R�2�V=��`�}\-�т��G�Q���O��Z}�4�j���μ��e\V�
��X�皯����I�Av���{��f��1��7>� $hz�m{�X��R8��R�����)vtv�^��*�����P߼՝�ܭ�=R�sT��[�����~�	d�)'�X�G<ȭq��7�I��q5��c�`���
���T��<�P�x�[Cɳ{�	�Q�Oo�rڧ�ʝ8oo���9^��^���v{6H���ti׷ݏ��CVD��ɱ΃֣JU�b������o��h�{�W*��T�ݞ��k�b�˅���1MdT]r��ﶒ���w�Y��4u�:��^�	���W�k���xus57�4���=�N��R鍩�r��p�Rq|�����{�m���~�*ȓ�uu�
\k	���w8�}\݋��5i�o� �ڎz:�C�t�Sl*�������ǫ[�]�u�Z�.N�3>�o�o[� ����w)���oi��huk��|���'��v�0�eJ)��Ӡk��mS�7J�Q[�м'O�֎��uĬ�J2�[0��R�Lh�����sh�IM���w~�ꪯL���y�ڽ��3������8�@x6���ÿ�ՠ�gǘj�sCs�="g��ı�b�	s�c�"�d�'w�\ư�z�h�ǜru���p:�4D䣅ۅr�PL�q#�B5�r'C��o�=�Y�9�������fn_�Ym�N��eSY: ���>�����,e.V1w�`]V���ZB�$Vn>ؤ�`���0�{�'��(xS�~R�o:�2�\�T*`���T>����Q�T8��mK��{Ǘ�=�l'�1�z?���<�֘1�#�i(���s=��6�TO��ʭ�>u~�]{�=�d�J8�Bf��Pc��^�Fw��y����_���KP���w>����������y��׹{���OP�\=�r���ߨ��Qʾ��\g.F�<T��κ������ֻ���ZP��VR
�s��]eY�aΔ�v�������"�D;C��$oI��u�u��&ѳC��X����肇��$����k�Zp��*sy"��:S�z�B�>�!�/{z��DD�pg($��=�r�'��I;	�h?>�R��\+�\�d�;ٮPf��������L������/?}�=�Oi���y��8�SMo�ң������nɖ���x0��J��=�-�|����W+�m�p�o�Ց͜����������=b>�
}�;�_r���-Ũ���+�`J�P��C�,y{N�e���f.j���}�j�hOw`rƜV�.�������}�3�f��&u{�����n�W�g��[A�.�.ɸ�Nb�Uj���	CUY����|��Ņ7�'T5Q�5m����M�~�8���#ѷ���bt)��m��f��,N�:6�\�f*>�	T3\�v��0��_Pf0;�P��=�+8	Tpؘ������>�ufDKO�"�^w��o=��[�2E�־Ə��U������LB�&a�}�3M���E�I�zL��ջ�Y;Z\�<Nz���c/[�v�D>�LZ���^X1�фf*����QU��#z��έ��
��D�촬�`�+kc*^�
�:�k��I���4{m։���R��K��wʦq����dwX����m�7�����t`��"`��;HV���p�v�PӚ�����˵7Os"�P/;s�{��!����}V�pW�ܱ>t�-�{�>���{T��|�{�	t7�u�xǵpu���:���\�sUAypf��>˜��c�Q��(�.)t�C_�Ip�v-��s+6�5oj� ������4��]K���+�\���*�f��\�~2[�B��}lo�?{�:�Gq�W{|�ؖ�6�]�==�=�3��zd2������oا�Ӡ�rwT�\�;���������yk'����c8Ǹ9�Dzx���۔|�5U9o�|g�}zTZb� �ٍ'#�	��GZ��ucx�$5��Gt4���E�h�^�z��� ^��3|�+n8'H�[��5���{��{g��\�ּ�纼�(�Vq{}W^���-��|}��c��U�eP}	��4��Jq��@�{�i�qmQ�KϐUj�BQGy��?���J�V�=r�l�ꮸ�,cÁ�0�l�r� ��Z��D��Y�8�6h���C�TZbm-k
�+:Ӡv�aH�=�M���œ,7�tfAX�3���W�{��=��K�VV�{�e�����ɺ{a�U��g$X$��v�C�|�ܬMcv뇞�mX��ݖ�.�=Ƴk�B�M�B�~oP+�BɊ��]=�+/��6Z�[Xz�6t�;�ug$Y9��Zl�ɸ� wxI�b5��*o �*���i!L�;�N��ڦr[�� ��I�2��gXD�v)uݞQ�|�l�4-�α�h��Ȃ)���K�����5�s�|2%n<����]f]2�]n�&���E��i�=*6�B�����ØȞKWq�&�qEv�0�ʱ��od�v���gn�q�=��v�vd�P0n��
]���t�'��w�:�Vs}�����8)n�٢w�K�-en�� �jn���@]�l��f�w����ۺb��=���硚��&���k�F�[n� s��m
�XE]��W"A�t�Hjc�褐��e'��ՍE1��v@1��Z��a�[FfW�x_V�H��Î�����vE���&���W<��G�չ���|���8	9�*98��/+f"�[X�١�3kV%�73"i�'���u$�ˋ�+��)@h][0�-=���S���8��Ջ˹���u^�v���1*�ڜ��*�X���y�t�ɬ=�ň��[�#�(�XsS�6����ʾ�*�4�Oqq�x��$H�vТ�z�RM҇eҌ��un��E5�Þ�N�9E���B]F�Ҙi)�N�JHF�m��T1�KcZ�#�6���^۬`mQ�W|er�8�Z���f���2�Mhm�@۽<�p� ��k�x���\�Lض���δ^-���y�.*>F�mf�V�{ܢ�wdخ�;FVC�kZ��&�%r{H���*,���V����&��jK�ҭ7-�8�NӶ2�.Q�وG]	�� +tM�i��h��c��ְ�39�Փt�&夭��Q�mD�{�����zRkv2c�ۛl�Z�S�f�����`�uuce2C�[�*K��h���n���g+2q�l.7E����F�����ط��qX��푧�n+�6�]p9�Eч�4���]���_�9�؁'6�5�>ȱ�b�(M^O#6��d/���1��7���i����ԫ,��Ğ���������a��V)�,�%kV�HG1_T�=�<X{���2n���wx5��@���y���4���+�z�Uګ��=����6�F�zkyA��e݅�]:�R�9FEa�v�襎f�W�<���Ԩ:�V���9���jo�E����j�Esu�j\w��ޏH_#��vc4s�e�5;(��!TgP��l�
��e%��Ŗ)ov �`��7\�������s����n��������j��Pm��6�UK4A�،��UQ3TCQV���Q-E41t��KcUUTZuD턪-#�)�����bb(�f-�f(�N�-��m��A�d���j��(�)����*���60�vqQTO[����CPTQE�M5EC1T޶J.�z\WZ��Qh��DQVد6�b����h�Ӫ��#�34Wc51�N͍M;���j���QN�S�Ayn��ɮ�rE4QD4��4��y�UAD]h�1Gl�QL�ӊ��`��;gA[������"��"��(�����4EEA��T�QNƫo.�����'LTUv��mMES'����Ҳ�6�k����Gdt6^:�74S�Dw
�����}���t����˃/�!�ѥ�.�TV]=�2s^�No�����,��.������
\67a'
�؊LF5A��F�����h��V�U��������� �}�F�����=_@qΏ8�n�b�3�
Qu��E.l�`<:��`�hW��iuxg9��d��0o�n9�-���P�3�����F��/{Ϩ�ة�j�q5S
���,c���<�c���K�R5u'NRZ�uP��2�5��{d��[��X��>y�{����||aŒv�f��c�Q�X5�^��T[^��R~ұm.��e��׼�n��d(�缍8�N8ϖ.w����Ս�./:����~�����a/������ܼe)�r�~�;|6w�����V����%pl���{��Y�-�V}^�9��ꞌr�~�:p�g��yN5�Jo�ݎ[7��׈W7c�2�T�Y��~�U��a�Έ��c�_nT���{�+m��/ns�o.��{�\TL�uj�.�Ǯ��U�^��Z}ԕr����Fv縵x�a��z�A�;��}�ݼއz�v$�-�e���[\��p��K����\��4�ʴffs��B$�����M�\�m��؜��+���m�K�=�=~�>�u��8�jsO�jTF!)\�MU���[���Gw�����D=�5��h:z����4��w���D����ߡhT��9QVEE�3V�'"��e��^�]����ގm.|�R�Y�o��T`K�0�-ro ��f&�����y��7yr�-�=NOo�;��y��U:��:yl���[�Ր���&6����s��.D��$��;�߯���N[�4�F9��&;�[�=<��B}t�Ϩ�Xk�&�c��*G�~�pχ'	�wۤV��v��n1$�q� C������s�ݓ?rǰ�>�X!D<�u4��ͩ��.�9y��d�ܬ|]*�>fߦ�c%�y?E�\�b�t��sC��=�o�r���#���qn�y�kE>q>R�(��ז׮�x�q7�'�=�ˁq��<��q1i�ٹj��'�o�,��ղ�\ץg"�p���w���7lȕ���@t
a�<6�8�>L�iN��K��v��r�ջMu�o�j؄�Ԭm�W-@�
�[�$�:��Z�O�kv.|���+��]�
�����K:��b��E���-�us�7kq�[�U�eK�����3z֘�k�[���}_P8����]������1=:�#�DƻqP{Qv��}9�m�w"sa�eJ�=T��*9Z�~����_���^���3��*v�ow�_�^MFT��ɼ후�Q�h����"Wm��4��]S���-���ӧ�3���X�%���/RT�/w�!��y�*��в&��Zk�8�,�Z�!�.�6����7���g���x���6#��`�����(��.yew�p�Qd]�����p�]3�����_w=���̮z���?\�[Se>7�����4�;��o�-����8t�}�:M}��/R���ƠW�j��F�����K����)�=�=]���ks��}з�亜��*mf�D����*�p��N.f�x)>��Ϩ��@ʨ:��9���U�^�G_����[�ٗhԮ���(/%�E�˒6�����Jg���ڋ��g"_���;Dkڇ���UW��E,������A_��Y[�����0{����,�f��>�t\L��ӌ!��c�gm�3�1�ml�S���B1ub)���9f�Nob;�o`�B��ޭ�:D宝����F�h�}|̺����kw���훒����i�ןx�����O2��O/X#�X-��H�TCGƥ0�"���Dfu�7�^�ͧ�pΝ�T�+7g��Ï;�b�q�3g��Ǎ�^u�@�Q>D�7���t�KT\Kkb�EEǗ1�k��I�:{��iM�_B�����M{>. �d�C�/�R��wRq��ߒr���i!�����vA��WK�U9��nz}q�U�ϋʱ=�遃����FP������PaY���TvY86�����&z�/�3�"�S�*׹�-�6��o�gq��Y7�`��d:�>B���e篲=�3�t�7�q���\�O"�ճ�&�6�;��Yu;ϱ]���|G��*���zSܡ��	��AprW�P�Q�W �O�o��ڛ��9�6y3ͼ�atCu��ɕ�Z�Ҹ���lx_"�l�ޭ�g޻#k<2%���BY6�8-���}���t��\uxX��ձ9J�5�\<j�1��*��S�����$�ϯ�U��宝��-�ˆ����g���a{>�ٸ�sb�=��퇔Ǯ'�hxb��<
D�԰f��xoN��-����v"EN��鬬|�m�8����x��+z�{�K��}�
�����%��'��m-o*`�{���tZ'>��	uԟ%��xs���?u�G�WG\��ُ�|2���:�-���8�`�C7q�L����{��w�s������@{�=W���2�f�a��>	W�t8�|����F&m�ݥ	X����}��
�ϊρ�^�@79
��O=��O�p�jVvT5�H�,��M璡���|�;�h6੫�wӌ�2:�b#�8h��oߣc%-��w�<x)V�D�F?`�e$�/{u!�^�����ϸ�X-}g�d\9�%���Ey���a�˹��x�NK��N��W{<�7�[�����@,z���z�giL\>=-� ����5�$ �z=1({���Edm5�N{�m��p�����ܑӕ
|O�-�Dg�/Ju>�T/�@���o����yGZ��cO�e��5����S^"��?������/ߑeי��-�����}���n|=�w��D��}d]�z�*���f�<����I���~4��S'�*�x�S0�fI�
[�dۙ(?/]��D򫛏nQ�M��;@��nR�<��*!`_!�>1�8%z��[���Z7����/��|o�N�I��&ߕ5�R}*�m�Y��}G{jD����3UJ�=0ݭ6�!jܮ{�����հ��EU�w��q̓�^��ް(���mM6���an{�P��Q��D�=�2�5��g�ܮo&hk�Z���"퇯o���3%�63v�;�a��0�A.Pr���H���w���ؙ�P�r��VT}�Q�Ԣ�Zc�
S��z�p+�����z{�0{ۖx�ǟ��D���������y���)5쫭�춐S�
��̍��H���L0�ׄ�>���c}�GLy�5���Z���'+�L�ݠ���i����������;�q����m��Ʀe��>���l!3��}��/|F0�n�=�z>^�Nm��G�3�k"��o��^92þub��2�xu3q7�f�iw��j��8{�V�FC[G�g��"��]0N+���=�6��a�_�}�0���\���}y��=�����Ӑ�gL~^V3�Wb"�׹��6F.,�^M�	H���Y�_tO�6Չ�N���r�;�3����M۸u�G�0:o���o힠z�FW��Ϸ-߶�����q�%,��q��n����*�3����q�q��M�=~�q#~����ƃ�v�s�^Tz�.sؔ�47���h����
-΁,z�{�
��F�<t���<����\*�]I��t���(C�q�TH���J��Ǧ�~9��U�/��
��H�s��=��+�Fo/�U!��6��;�̝*[g�����)�B���y'�s�AAGj���y�/�V�l�m������.�Y�O&�/:`	-�m�ա�rŞTMt�^��'V���ׄ3�)|��:o�ZL\<3M�B�]�UԸT]9ut��W���ѩ�fy 3��߲����rª>*�f����#�32�M"���A/}��C����"�U
ն��ꡩ���,\G��u��f��S �]=7 �o������h5��N7�fq��R���o<�Luzd�b��O�5U��w ���,ؿ�z'�<g����j�O��c�Qzg��X%b����v����@�O��ސ����8٩��UL'��tG�����-t粰ײ�w�����f��8��	�;=,e�7�>к��_Ѿ�'�ɰ:u����`Y8;cW>�yk>�Rp����p�c���ܪ=�@�\ux���
f�f�w�}^>9��/�CĖRu��=��>���-�9�Ѓ>�:��U��L\!�>�q��W�f��=(=�i^��w��cѴ��UW��3.xc-���(�{jCy�u�AY��1�ț�&w�\a/�Cu��F�B�ʡBM�����
q	��g�y���,s���^���N%�-��8??a���7���1��Q����q\hy��,cs�z����j����c��z͹t��HZk��U�F�������89ov��C���M��_��k�&��x�C=�Y�0���9�%��gZ&�^�2��
J�a�S5�S����7b��U�8�ӊ�ӯ$ٍon�<ZԤ9$:gu�uJ����V��";�#���᷺��������go��m2WOO�G�uT��+��� ?��Z@�����l���f�MR��2���TG�����_ý��l��U���-[K��T�2�oL�����rћ���������{��s��}@`/��/'�|��D�ԳR��H���X�-����s�46�����m���ڇ�W�P�ϙN��ף�H.���s��(ʜs.H�S��A��돫(��z�^�>G0�/���W�����r���N�o_�������3�7�@+~ˑV�$\*�>5+�z����YF�U��3��{w�Y]��
����H�ʈu5Q]xņg���������@�=j�>\|D�f9��Y4�_�V�j��g'�.
]lm~J��h�G�2�/Mʚ�D� W��R,�x��rrEg��[f~7=�g��n�HaB�\�>���3_m1�Q
�.)UE��>�z�?wc��Q8��
�۵1Z=<����	�6(����=�OT{�v�<�r�N�㳲�	W���L爮v=v��4l�ڨ��rA.�bQ�j��6�������P�!}[Fr���<�r���:%1��8��.�x�����n}�c�U�M�]#{��K.��4�t���)�ܢ��`Yci�i���\��ݶ}�O�{���f�/�WWK�b̭I��q�k�^Ne��'7�P�+��,EU���H����}��_��� m>z��EN��/M蛇[nu��I���Ƌ�Tgtd%{؜�����S0Ɗ�hӅ�3�i��z�7ړ����p���?2eu���4�5�P���:*R=��J���c�S�쇘��U�5�ݷ�: �	�>Ϻd>���I�b]Jg�+ő��X�*��f=�:��1��S��r_��
�KL�ɕ�q�,/g��a���Ǵ�8�S�wHx;��!��C5^������//Q�7���!U���{(˔��L����qΒ7�s��F�������u�W��kG�Ӵ|^|6Ks�Xg�e��'��4���aY^�a�8�{�`������yB�Y���6�e�h�^�hxܹ>_@�!�lĦ{�23g����BTJp�}��dP��>i[s����~���=����o�r<]��咇zb}��	~r��l`��������~+�?�o/����KN�c˺�z�W]L^��R���PU9�I�P�����'��1W���Z�Q��z��W�ۚ7�|;���0��#^��7|\ϯ��"g�ˢ�Y���Z��_�0�\R˨�5$�|F���G�����s\�W��kc�W���Dń|s����Ge�+ф�7���+U�wWSO�a����;	hި}���h`�\�R�l;�^u�.�h`f�'#-d��\��{/���G�)Q�h)D�K��v�Q�Vr��i𸩫[֮�|�+�@v���3w��C5[A�2@���znf�9�]��2�� �ONJ���2�.u2\Uť�+,{@y^ߩ>�A��T�n�5�:�= v2:�\r��ߐ��Q�z���	o|��c�֩���� ��L�.�R�Ԩ~�FMC�;FD�w��w����Tǯ�̔����u|�"�ɩپ�o�}t��Mo��{��z�d�<��o���AG�[��+>Ehj�]G7s�*�g�_u�����H�7Ł?*w���au>���c'ۖl���]�'�0�|�(�Jgi�
���V�J�P�����K�=f�5����G���~\��'�#�Sck˷4���6^�k����^�t����W.˩��S7�z@N��1��z�Rj���u�>ܫW$�Sڽy�����u����J
�ti�é����`\R�)�ɟ�İ����,���\�p��<R�}�8��X�.3د�DyIg���Y��ͫ�_��ɴ����>�?o8^
���<�N�=x�Y��W���O������)�,�=dz�y������Lj�A�����A�6�O��D^Վ���ٶ�s,&��A厇��P��yL�k4B��5s:��Z��=��5���̵>ۨ\�9��ˬ.|�[�M%��P;�GB���ן�Ev����j؄�a#�$#f�v汝C+��;���`�u���H�*��%s7�=����eJj�c
��%=�;8��F����Sב2�����n�s�F���/.�E{l�zaW�.��۴p��l���G�g���p��`��f�ݡ@����K�����Z���9�q�7�d�n*�N�0�}�B�L����Z�͎�0$��N�2���&����^����q��2uaw��j���mwdî�u�v�_^*\U��SU�.���N�0���pΓ:}�����S��˂��4��R�
U��'�F`�l�ӱe]�PE�u%zFKIt���(��.���#f@x%�8_i��(�P>�cD�
ۑ&���U��W{i�.�c�9��I���1-�-���O&��\����<��>j@F�۲f���ML���:Iؠk,�ܾ_Nˎ�\-�Iq��*7"렩f�JU�븚ŭ�^�s��,��4pU`�U��
�S��s��
]=�)��y>r�Yg��mU_z�g�71�yj�Ib�H������FU����� {We �yrU�2��P�r
{\,t �"� �lbV�ɍ)��	�샵�-�k,��`��� V��m_0t3]0���2��\�a���묚�����E��qY��T��#�ɏ4�oe�佋��1q�Xf�����Wv2�ɹ0T�÷j�[�y|���YWj)wC)��r�H��+�����;�W]o/Lͭ�2�Y��c�U�[=�3i�椦k&���F�g�7�`���öu$3���B��"֦a�1cWZ3>b(��e��k�U��6��iŭ�:��nR��Sa��v�d��؍�sVu��$u��;���ںS���s���>s�@��.�<�An0��TR��6�'������v�]i�Z�f�ë���m���]+.��cw���eծ����N)8����ͬ�G��+w:�h]mb���/.�sj����[�i�bv-�FTЗP6V�Y��+Fܦ�����b��%�Ɏ�.�z,L�%��y3*�R�����L١+�%��y���wi��s��ܳa��;����m�b}w��H7nέ�D�F�ъ���XͮǊx��XR�ŝZt�R��k�% �gCAc��
�ڀ��3�ӆ-��S�WE��MP��'	�e�U�+��hq!��V�٫r�i�� �C�vh�Cwt ̆��dRS�5}Iuf�S�b�&�spcVcȫ1��ky�u���#(�&FGvK��C�*V�Q�� {#�C圷j�1�� I�]	���"݂�T9{����V�*�V��{V��V����i1�X����#P襈c���[�6:-}��=jK�q�wy���i��sPeM���h�/!Oe��r��;��u������Z�����j����ji�j"��������tsU1D�Ӫ
)Ѩ#�؊�wMI�;�]'�Eh늪*����h�+���jtV��)��j*�ձ]8���*4���m7��DU7�ד��DDD�����2�cE>l���q4�Pݍ!�q��RPQDEW���Qj�
J&)�������b)*"��D�$MSMDE'���F�A-4��M^X��lđ�V��nڂ	��j�65�*�*�����Eh4�%!UM:1504�gy/�uT�Wy�UPQ�yi����V�1SAW��f����D�%,A�1֢��������T��AE'Z;�cT��g����6��vt��uLM4�]�A�"��{��ߞ�8���輓"o:Ee�5�zGh�
=�y�>�c�B_�F��a����h� =�:v�5�ɽ��{B������6�;��o��r4�{��b5��,����n:�~��UR����ײ�<��Ӕ��ȃn�&�'̫ή�}ǅ�O7�W�~��#ޟ��;�~U��	֖rɵ�cg�}�	y��Ӻ���>j�r��IIc��\:|���u}߀|��נ����`������/1���\·��x}�ck3�V�9��GXQ�K����9}z��^]W�jR�������~�L�yxͅ���G�3.d���	��XT�'����a��^�l�y��5��P�"} z�����ga]. ���SW����pLN�Z��~�ٛ/�վ)��%�)�:����!���1_5U��(
����d_�D�g��~��K�������a�~�=��b���=� ��si�9�񞨚��a�����wT#~�D�Q�C 5�n���:�es�ƍ-rB�.t����_	�x\�G�q�:�Dz��&�Lf@gӦ�g|\�m��cC��h�i�U'ۮ��9�ꇗ=Ek�7����:S���:ʭo���Fo��
��f���楴̕�e*�J�8������{�yN�X���ٵq����z�mA/i�nFOM��*��(T�T�rm�X����d�A\���aNQ]�����o�k����/��|�1`�ka�{�$��<�]tu���)�Y|�m�@��*����/�M
�m���E=�G�.�\/��5Ï�=��H�{}�W�;���&Ttφ�[����u+)��{�/��6:��{�Z��T��6����.��{&Cj�
�]���D�L��+��G퉯m�n��R�����e2���+����%�������Wx���)C�$�Ev��W�~�#�o�3�}ƃj:�ܬ/J��R�w�a?	t<sB���IW��ݏV��;�3z��hr���r�f�%��2ly�Ԡ����N�
��n���N�=�rr�R���YH��9/�p�\r���g���-����i,?�E:��(���Vǟf��Wf��|���w��FGJ5�Inn6d�s�46���� )���~7�0�"���@�}����Cj�J�gǥ�����{,���S�/�:,\lĦ{>��6�޽�@>G0���Wȉ�>Ŋ���_��|ת=s�rzS����D	���� 6k�u�+~��;ϰ�SQo_�^��b;�kw�B��g�6'�ҡP��T���鿥O�{¤����
��}���ճ�ؿRt���99���QG�\qr��'MX���c��HV��>ڷ�0�$�V�fc�Bb�Z���.�x��������Zh�u¬�5|m>�ҫr�3��5��$��noI���=�|\�<W06tz���SD�����H>�����?m�Y���Y}ٹ#�}���O�U��3u�$#�!e=�d�WK���9��2Yk�}�_��T��QU��Zį�_AyV/�,5"kΊ;s�����y+��[xg�}��� U������i�1;�3��~�!z�	n��4�s�D\C��6tj�T�մg1��?B9Hޖ�].�s�YU�ϧ��=��'��%�r�y�)M\=S{7j��.J�"�1��Y(���>�q�O�aU8�o�S�n#��m�����L�G��{VF��z��@w������.>tX�����oԩb������2/�ɝf���h�#�C���P��&��&T�Tf��Q���&f��u!wؽ���{A�Q�}8��
�OL�ɔ���,/d}�a�|���xj�쮗����� .^��{1��>u��N�9RPn\(���`e�d����w�"r�*هe^fkz�ώ_��<����~�Z%��,�Юhi��?Lن�MO���b��p�4��=wc�Qb��ʲ��7�TO�tݩ�����%�a�Q]�V�T�U���k�{q�wK=s�^�<����#�a��G�E`ppj�S���d#��POP��I��2�+v���W��p�X�<�aQ�iؓ�<�Û`�����Ϟ��B}�����k����{�E_�������d���)����S��Ƶ��63�[�����n1֞�l���U�Q����^���#����*-�9(x��*#f%����虎]>��[��ZY�ī�����= �����giLYs��m:�ڨ�|i�3.�ת6��+�X����ݢZ�b�O�V%M�es��'�+=L7
�3>dhs>Bj�L[���f3v<k��@Gv�DӪ�j�4��"��H�<�����>2:|� Gg$�=v�=�P̇�ޜ�+�=r&��C�X&����b���e2)@c�U4� ���[b�x�8}T�eBC=��5Tx�Bfe1p�R�f�D?`�&�T��0�ӝ�+-O!�
��q�'%t�I��t�<P�w~ k�T��}���6�����Oa��	Cn=]~A����S�6k.��߼��	��M!&e3q���W\NA/������������/��kt
s*g�@g��P8���ᷕBm�U�s�F����r�����`�|'�qx���߽�;�{�͵�@Q���lZ��``��Ա.Wm`�i\+x[���9q���A�6�n�o4�\\���s�LGU6t�3�|���A�&�s#����
�P����|㫽� �F�!r�"B��Uݠv��̙"����	�SF�\��<�H��7�i�Ϡ�����`�]�SFL���:�1��i�1*���u��|�oU��;+��l1�s�\g�R6�p2�5Ǘ��f�&|�t�}�	�
�*��*��n:�N��^[�W�;�E��o��v]0N|�p
��܁d�rT	}�E�*��>;=��]m���������<ǐoK��/ȫWV�� :5�@7��͔^�SZ�&�U�����+Of\q�'��<�Wq�����#G�~��D#��,g�D�g4���Fs5�sx�e%�󻡧����6�	��|ʿ�����q�pW���dx�E?g�$t&Q}����r�l���]� p�����W�u;6[W���x%������pR7��>��|���\U��̂*/����O��@�l��1�f=�ÐK��τ��]�>�X�7�VE��-{F/R���g��a�Au��6��\�p�2��5ax���w�2i��sp����~���ݎ��P�u�F��x��P�f�	�:�7j���	;����U�e��*+*����W�t�ouAچ��	Ss�/��*5FN��w�ʅ�^B�8)�]C"����ic�� [Du���J�Q;�������`s�:I�.�y֫X��5t�Vm�8 3���.KV�w.�ۻ��T����wfw�6�wugSy���INț���U���z|&���0�<Hf+��r�ۗ���L>f����G���E�7@�#�
����az=U�^l���O;,�Txq`Z�>���מU��n�Mu{�T�^t�<�G��N�Pj�ax�C͏����!a�:φ�GS~SL�޹������ݱ�O��^o?\��1rWd��o��;sO=����6W�-�3�� 3������ �R�us�3<�=9��ϣΗdy��=S[>�'B��J8���{�W��oK����+� ��8�=�
�mQv|��#}@N�S�6��Y~n�(��H\g��7�_���*�	�o�&���=�O�d����z���%��L�s��G��w��#��Qǒ�nZ�܏{l���Pͺ�a�g��.�z�Ӓ՜\������#�M���|���t�n���,cs�{�7�P��,�G5�����=�Z��h���}����@�+�z2[+vly��R�}�}ǳ]������=�ӔWt-���g�q{�t]8V�GB��d�%�z��{`^\�f���k'�����LDeY�\�>u�l?�!��~,S�1Ωt�� �)q������Z��@_���eF��xr�Ɗ+:�_`e]��98r�ZE��]�2p&��#�r���^;����+%e�j�ut�N�#�k�6��U�'V���^i�#$�]��R�Ԋ[1ӗs|8�.3�����܇���46Ks{2}9������59Y1�yj�9ՂZ���hK��j�yçn����Dy�=tF۪rE���b�f%pܥBUD[v���o���֎�����wӵH�/�ɸ��?]HطU��D���7^c}��ݨ^ /8s��̧���T�g�r$9ʏ+,x��g�'����x�^y^��ay���qf�=�^�zr�?��>G�����)2��q^���)��~��%�k�z�0����.��.垀O��Юr[i�^���5�����-:���>����U""�ǔ�>�Qƚ�t��ݭ���},5��5�f��z��Mn���߶P ؅��^��yb�[��,�='����X���j�n`��2D���r��~1W��k�x��Zh�w�G��S�}���C=���x߈i׃�j��n{�|�C�#�ߠ�K�D]�K��j�lr�5��ǵw~��m \q+�.!3)��8�����L�G���v�ˬ���-�5�S�U��6Z�-`UB�w}ۺc��|u_���۵i�J�S�y�������/�s5��@.tY �G{ˑv���L�Ȧ@μ!�et�-HG��W���ڜZ{W�C�9�x)�7�,���ۼ��+��i<��Y�8����֕FfU���jtNh�k����y���7�262g|o&|�ϣ�C���Q��br�3M�vC��🻢�S�ڼ>QE���kΊ�>��.o�]�*-��"�&S7�,/duXl����}��h�e�tG��&��µIZ�x;�*��G�;�S7���\l
�{l˔�����|�yew��yo�z�%~l�徯-�_��W����\ ���U0*(U{�q����O�<ו��n+�g=>��-���<�#z_3�������uL���uR�t�T��MϬ�[�8^�b��yċ�����*-*�/�x��F����65̹(\W�+��WEI�^C�1���g�J<������;S��3��%#���l�%W�X�ƛ���z�	���;/��7 ,S���Pg�$C�+��ġ0o׏nh�c��,^��>f����Z!����7���ի�z7� 
����D���w~�Z:��DT!�:�Ӓ��I�._�u���s��y�fdY���?����s�9@W�z�L�+�L���X�9Ydo�r �n`�z��q��v�uQ��5���ٚ�f�l���IQx�=�%��0��V,/���n� �#��)�"�QN�h��f\e�����/se����'e����H)NhA��{hQ=�Q�}�7��P���rý�@e���p�\�D�7x��ݍ�f��ȟz/v}�򻭛�uA�|fO�G�Tǲ <�~B���?Y%�����W������T�����ۉL��Kw}����i`OS���c�ީ��Uh���&�7:T�#ӟ"�eo���t������AW�/GUo�l�7�F�o�,.�_�>�L�W[�N��ɨ��8`?`3�ʠ��񧛡l�x8,�����gU���=G�� k���{zX:�	i׸���F܊n��7ch�΍x���}�a�����@�����A��;ef?����i��R��U�y��J�_Q���o��u}��/�]����0��v�Y�N\���U��rȫ��.0�>a�m]'��,UyQ�y�T�K�^��^��!��uj�w�K=��%?����s�W����v=��5�<�ʶZ2<���Q���/�q�z}��߯��ν� -���{ר{k�fֲ�W�c��z���M���l�ͬ������F�޿\v}2��8-Gx�KeF���}��_"�H���t4��66�Bp��{:�^���3���8̵_GdD8>�ʧ]���\
��W�fbQ���f��K���y|/a�^
9�aA1&�e��P����pE촦�+ʴ�rp_b���m�*�Z�t�:��o�m���K����� �6&�5eiY|�hΥ{
�$E[���od�Y9�|�}�����~횏\J��!g����T��W����c���XS��7���a�f�w�ٽ��N(�}�z��}R�!��)�5��-�D���ȊRaVg,�0���P�ת��3�5�V�~ղ�\}�k�x��
| ���E�����*������i$s�R����䮞�������{||Oa��X�w��(�j�>7�����
{>�5�><,�Rgf�ezųڳ_�Z�~ܼu:�W��.P&���T*B�>�����χ� <�+�˩fB���@����������Ƨ�����[��UI!r���vA�U�:]C��T���FϷ�kޫC3i�C3ſ��I��@_P�1�q�V�4��9`��ˋ7���SL�޹�e�M��|"r�����	"���\��62O�Kk���Nz��ۇ]q8s��nR�q�@�_W��KQ�-?���Ԃ�����8ϔ�O��X_��2��/��;GT=�ȫ���O��Z�s�^RW���g���X�{��Lλ�g!�]�y�A�eHo �Ѡ�UX�����f�2qͪ�v�uhwY�cU�{�/���UҒ+�x*�-߫�,Px�gl�Q��ƫ�мl��D����U�u�tD��R��)���X!�̡[�{����А��Y�\�:݌}}Z�b��l��>�)]*����glͨ��s�8L��Xc5�PM�
]��$��z�R��.¡d̋��,�P�wW�9�j��YG�T�c�ۺ�C�˃+f�a[ƒ�#Tzm����.��̬���%m�}f#jd�n�|��=Ì��g.`ƣ'��*�r�VJ�tremu�;۹�A�1�xj*��p�3.�%�f򢍈��^��F���gdC�"�E!<)uw"�*(����O�m�Vn��*ķ7�K(�2�L�ӕ�
�l�.ӹ�N��TWQf��r��F��[q��l��N�R�N:�}Z2�ҫMF��]�� ftq8!����_:�#
�u�3����B)�ɐ��.��CL�WՔ�%J��\����Փ5���+HOvB�Ufs|03Di��"1e��/�^R��O/�d��mMU����.�����/&��(���K4�;o%[ɭa<�3�`[���g�s��8�ӧЁ���WWH����p<ډ�)��R�s��<���}�Zr��;[��\�٨0���ԫ�z騫y��呷G����'V�nc��q�eGIV����{�B���S9/�{O�qK�k�ݥu�d����YW6�fҮ�8��yȮ �G���+��(;o1��y�7�KL�Х���Pg^���2��*f�&��R�qe�e�ѕmT��V�<5��ɦ�jQPy�^�р��Ex9�:3+��XX6��_b�cyCp��J����n�nw��pJ�ge�����;Vryvo(N���e0Zʝ��rM��2�mueYA��hġʺ$LX��t)�I�v�F����]�]M��׮���^�iɓp��_`���w����O��ܭ�a�k�y$�}H��ԫT��͍Ą�YY]��J'e�ڹ�!�C�ݷ��8v���a1�bnV����vd��4�,T��ՒrvVQ{n<����Ǫ=¨��wv���R�/yr�Z��Q�����&�n�9��b�����Q�ȷV]��ؗ��[��|�Y҆R#�Z��
.�I+_|��{�_ U����m�\i�Ջ)[JV�B�a��� �y�A���,��=�Y�U-���a?e���)��<F1�d2��VDo�UrlT��:v\Z��#Wsy�u�g��$VY�j���� rmL�IIN�*������;O]J.X�M�G�/�H���vQ���"�V=��8�Ż���Ӷx+�%�6�K⬬c6���85j����b뫗O�k�r�[�CE=��K�Ct��� ��+�x�V�@��o[�J�iM4��6���l�����Rjp<����8�po�҄>����j�ө���;a����B��D�r����uuWWPP��;`x��&������(Jj��؈)�����ETT��u��Z����1�W�ΧET�ca�61�L�A�hj���/3�����N�)*��*�ݒ�
�d�+Bwb� q����i���#�jB�A�cTkAQ!Al�
Ƴ��-5LE1%3h�2PEHD$Hh렂;b�T:N��ӯ8���M���4��5E	U�h�l���y	�e��DB�QQ)y�QIA@AQ�%QAy�Q2�QDILUS�f�:�d(�i�Hbimhü㪨��!(�"���)��S͂�����������(�Z
#LE,UӐ�Wl��RM��U%P���tEAC�����D�����A���� ו�5C[m۪
�#��I1Tby��]�ǯ޷�={�c�y�{/2Iʭ�p�ƶ�.!	�49ܝ�+�1�9oY�*���>Y�&�96��ǭ}�u$��������yWu����gzc	���!��P�>NUx�x���7�ʏ�o���o�1!��8�S�k{<��Up�KH���G��&Z>Ϻl7}LX����-��}.��t�,��h�^��5Q����|Q���z�×@>�WzD_S��\���l�ɱ�m5H_9�=BT���=�-�Zܾ^�]��3���2=5��?�eG������+��	q{���u���ٺ"Nc{�/���)�>��N�|�|\���̩�]Fy�j%��ِ��{�v6��rK5�w�U�\}���WA����*�Ӡ��`x<��~�L��t<X5�U�.
�O��l~��M~Z�>^����~��=gc����j��_��_���r+�u^���Tc�5/o8lf�)��/�󇎑)�;T*n3�l�@,eB�P��TƜ��ȉ>����E4��dx��K\����u��j�ZU���c��k���FIa|�z���y�͖g1p�M�),C�F�}�#��N'�q3O���_������#�S�|灚��<*!]ׇ\ӗ�=�g��"�ʹ4ؾ�@I��w���3���ѮW[VP�^s�:�4��������^c�cmV[̨r�`�|�Y��آ�^�ʁ+c�^��n�� �m�$��[��۟s��o+\�r��P�vr��Ɋ� 0	��q�]-��e������1�%��i�{�s�(�f��A2T>��ۆ�*�qز��9�=����s�׃�B�0��c"	�^��,'gQ�VM��GB�T'�_Vќ�w�W���ȹ�MW����}=3�_�\N@�^��φ����U�������"}�U��[Y��~�-��	���	\b�q���2���ğ���d�Ec���ۇ�]e�R��O�����:��m=�j{̞������ݑ��c��E�L�7�>E�L����b�T����2L�.y��ހ����u-꼟Eס�¸}L۩�\�G�����ܙL�L���V7<�{?zf��<�O��	�f��6�x?D�C��Np��ӛu,�j2{�@/��3����F�W����#��hn�<�┏�ς��[/����1N�e��-�ǦX����.c_�\��<'���b�P��ny%3�0ߦ�7���G�#G%��>�8=u�C��'���!�lĶ{��ƖH>���5���9��uތρ�|&�_�ڄv_�q(�c����Do�꜔~z������2x2κn�ϒ�n����2��w��b�Y�WZ��7��xħR��nU�a�{te���bno���1��#�Ս�W�M��JaH����PQx�v�sF�����Iy}WԾ9�=�;Tp�cF͜�o�7v>��积�0��z"֥��W�����;p�N��Y��x�V���Տ~	�nù^==]xy>Q�ɪ���]w`�(M�����5�6+������SW��h���û KJ|O�B٤jޟ�n�\(.5 �򢷼C�E�L���̉��b�TG���j�yH�wg�!�:����i  �=|��Ϧſ���r�K|/:}j�{���l~��O�IW ��u�p�����\�N+��5b�����q��N�n"<Hb�:�,[uJ^OeX�,5"|�x�=5���ÅY~�[���g�7��wʷ=c}���N�<fpxN��E�J�629�l�~����]�)ߚ�H
�Gun��>����J�܈ڥ��#�HZfS7:dǫ�&��f&����kʄo����:�Nf�qf/G�c��4�d���u؜��W��,;b�N@�uH���L �O�����K�Ln��^iO���Ӽ���1��V���Ľ���5�חC	����d1��"|.�7qԽj�&⺹�{}>���4��H�*NVz�4
��r*��)����Y虭7�Ŋ��������2C���f�V`�yQ���~)����ܦ}�\�C��Ք�O��=�t��#��f�!�F��}Ɯ��U�Z�;ziA�z�j��
�.Al*|��vWs*�Z�|���>pٺٙò.�"��dH�e���C}Ḛ����5��D/Jev����U��Yޠʾ�Y��إWE�f���t���,��p��m�z��G~��0��;XoK�\s�z}��%߯��{"5����ĉ�"t��>�B��(�7y�i/��Wt6�����G�p�Rɰ�w�J�y
���0�P��=�z5�mitFK�9/����-��F�����n���'̫ή�&}ǅ���R^T�6G�k��u.������/�%}�"�����D��ىA�F���O��� ܵ�����,7���f�\U����Ϲ�|vX.����{6�4W�雁�#�V̀�ӕ�ck�ǹX@~9�"|�LQ0�C���A���-�C�+��L����9���x ���j߬�_*�ʿ�f�x��]Dy�[��*��n�W.��2|�x��|K�Q
�ï��h�/H��W�1RG�W������5����w�ee��E�R����9�+�x�h(4X�*��Q���x�U^�r'�eK�!��&�#y$����#�lJ�zg��ܜ��c����ge����:�Q��,^���Z>6��TF�U��/������s��в`�ĵ��x��.Fi�$�7l�����z���,�N �i�R*��p�w_Eݎ�tQ�2�w+���PԵʾ�D*�b��J�v8����_J'r�>�pŶJ�����aEn	�N�ɺﺚjs�_p�����a��;Cz��W�ᬄih�ņ����ç���-�d��W���W^�15�E3�;C6��?W�v�ϐ�����|�c���b��yU5�A���#�Mv�lK�����b�r˿0{��?|�7�7�^��ΰm��h������}���_~8-o�f*�wΜ�ӛ{����Z�Q�jw�o�S������􁱉�fr:��Y�~�~�Q~u!�.�h+q%;��@tNfZ���{��{{r&�ɝs�K���Cw�z�W��9TrK���ϛV�W�-٦��_�=מ[���}����;�ܼ#~ɴX�ɖ����}Tō���6��D���t9ĝ�n�_�k�}^}w���,��U�V����^3y-������!���/��*̽�Ac�^��X-�u2�#��C��=p��[��{z�<����h��5�qSW
s*;//�,M�C�K�͟:�羠0M{�졎Y������ 7��|'�M�R������۝�ӞM��~5��T;��3p}:\7`x;��e�W�\D�>�c��F�ky
��)����|[��[�eu����j����.+��a~�J�h���;�pJ>�sm�5��2X�@W~��8���l��u#]��ஐ�S�}�z��8�me_Ã0����`�+y��`�u�Y%E{�;�S�#+6�^�n�D���&<Vxc7�˨��¶�%�����~��r	x{�1�(�;/���~�ǕO�FH�"Lɿz⹻�:�ˋПj���3U�{�RM۾�B�=>����T&}��S������Z�+o��˪݆ԅ7y��o��s%Ǻ�	�������RҧkC�c����G���6��,T)����+00 9�`�]�SgʕX�\PՊ3_>t���j�0�B;!e=�vA��c�&���/VS]�\�o��N�ｵ��U)���W/�	����<�ۇ��Zo�N])���a�A�4�wy�s�0����p����el�{&���l�j�T���3�qc\g.Z��ֳ��Xz;=���z�����f�8�^�W��E��xs9���7��<W�dv�������tm����o�<����P�wP�q�W�����q���Aa^�D�OL��}�m���5�e9���󷳋<_��>g>~���EV�t�ȸ���o&|�������_&���:�	ȥ��7������(��D�u��J�yX��dv�S7�s���K�Cc&S8K˪�f�Q|�=���3�Qi$z���<M*;F�=�"L-۾�.m1ҩ�Jt:�S���Z�q7�DMW
�f��gw� j��)
�0ܥ�7�#=G��ORf�d��}7��]W\�ꓘ�.4�]�eGK�^<�e,�5�p�w]�,E�%�X�cR �����=����Ǯ���w�?Q�6�X��W���.2�3i��%�n��7[���XH��+�㔎����o�Å�O���y��.��no�(�>�����#6pg���[=A�.\�1����0���3r��ϼ=v��!8*k�v팏NW���Cg�0v�͉��gJ��\��6��C�����ތ�L�=/�^�B��y�J6��]�c�"�`Jg��(��{]�K�6t@^>�ܥbU|�ڜ������v�]�*�b���ǧ��:��=7\�ڷ�@w�fA��$�B|��bP�dEm����M�>��􎜨�S˧+[~��y��O��3�U	S��.�{2 �����uG�nf�7����!�fR"��\)��t���|����c�����(z<�ѯ��������9@My�Ȼ�t<T#�r!Vm��x��꜃�@�<֕_kR}���3[P�USᜪ���z�����KSC��ȕ�C��W��jf�y�u�.]<e��O��{!H���L���p�"�L��b�o�{�K�W������%t���L������j��*�H^_�a����R�9����a�b�5�pP�=6����]�^��/��w.)ڂ�-}x���b�4�:�Vz9*ɱ�x�J�0֯�����tE��CS�Vp=�P]���M�W[��z�Y]&s��WԒ5�w�z�}x^���eɶF�ʛ�w�ӡ�/�d�⫧*���#�H.����������Iu����Ezb��Í~��:�z���hTV��'�/+=W��>ܞ�q�@�uH��u0fz='E6ڲ�0߸�^�R[����u��r����>�N�����뺡�3�7����rw��۫غ�y�*�#����X�M_��O����c
�CW��ڜ�NUǪ� ���%�$==Y�W#�S[@�4��w�O���G:g��G:�_/Jev��</�j�dw��+}$KP]0O� �9��=���Uv�[W�3�e��7����,��o�+=�/ţ�yO��K�x_�k.YR,��P,?Fz���{����xGޕ@>ʩS���d�>y-�y6Gܫ����|s\��Dn��jUS3S��I�L;�����V%�c۾j���X����C�q��,��,��,Kʷ���w#����}��w��dh�O�C�����D,=�˺/�{o����%�,~�(�W��7h��ҟw���%�񿋝�<��;��dV雁~t<�I~y��)Iy�C��Y%z܏�h!]��պ��8��Mn�{n�ɋ��W�rIb}Z�k��������i�����{�_�K�Q��</_��=�~�&Nr���6�y2wu�*�M���er�ҹĂ�`r��-�)m���\�Vν���fr�Ol�sϏo���^�
��H�s��ʯ ���}o�.@��!�_z��/4*�`�Z�������=5�\-� ��s&�z}� �a�Ba���ϗ��q+�����&k�Q������g�=�uyh�Q��F̂qq�{<��:�J�!�Tz�a�)��~�>4�W��@��*z��ƭqZ�C�8\�o�4ir��H�6p~�q��f���W�<-Hu�E���:��\��E��5s���Z���Y�� �tG��u�b4�t�]>7�����'O�l����e�w�|�������u�/#�c$׼��碻O��8��a�_�5�s�?Z��f3o&_�֗!W[�є�_y��~3q׸�9��z#ݢ�_��O��hҧ�H����{��LJ��л�Uw�{AL)q>a �;] �L�ú��r_���F�=�!���>�f��Cz{}j{�;�X��Ȝ'}1ѓ>Ns���;�x.��F�K�Uj�c.����үZ�Jr*Rz�W��
f�e0�>WzD_���h���|�l7}LX�n�I��<�e��&.3E����[9��n�+p::��IV��N��S�;�w�*�mp]�# ��R����r����ϝ���o��-����ۻ��sq<Oe���g�c�K9��]ݪďf����E^P�z1R��em>���M��ho
z�r�;j��ƚ�����]����6q�����v��s�QeH\+�����/.W��l�ɱ�mfA/Ǯ`/�l
R=����B���Λ<����!���
��6Ks~�p=ʪF�{`^\�ev{���������lv���?{���g��'<<��������@���n����l��s�5)��ћY�X�{Am�+��X�YP�o�a�Q�(�x?T��N���C���WB��u,O����tTy��;�6���p<��D�5����R6K�ro�~��e�O����t^[p<��:�L�$�*����^=�]Dvc��Cb1ϸ�H��*�>1Q�Ԗkn�xǴ8�:�̇�v�L�x�f.DK�/i�7��}�hy�N�K��W��TG��{ר����q���w�_�{�)	��K���{.&_P�>2�w"]�Y�!�����x�p#B,8���_lؿF�;CU:=��Q�/O���c��ɱ4�ŉ��
�ۆ�*�q��vo�],���ey9]��E��Ͼ�`	�S��3�!i�,y<�E��&��
::�>@��w��D�� �xű�E]���E����;�p�Ne�h���vmf㳎����GQ˔s���v�j�_PDmZ�rֳN�N_/�Xv�7�{d!��:�9�żvp;�
�'E�t�Uى`���/guZ�vwa\�H-pB\��ԐQ����F]]�u>�0Ja�\���P8�ge&�29j����.�=�n���R�(��
�`�O��_ٽ'-��sWMV>���Q5i>���0cD������Wa[q��H�o+&MI�HT�p���۲Fv�v˦�h��vFr�kzrq�ʶ�y�Ң�K7!�vY����bL<�
���n�ÿ�|:��F?|+]G���jp`	j�t�f��fۈNH�MC��Y|d��@*��Fc޾�C%iwj3�9˝��]��H�/	�6�MS�.�(��CktQC;d�74V��!@j[� @Z���0pQ����.�c��o��t�mZ��X�z<e9�n]�����}�X��z��stml��Զ��$}:�*�>c�fv��\���2�g���(p����儋7�k-�J�X��|��;[]1���݆-ʛ�ʙ�lu����%��f�6��0Qcks6�s��D�̑
To�������v�#@�̓gR�
�Y�ӻ�-َ���ܘws�k��Ec��ơ�D��Vn���m�<�f�@�6�wI��usV�K�gJa���4Ѓ�ƗM�NM���cN�8ʛp�����q�f'َ����bTrSU�����*�;������}Y��5y�c��&;�q�76^j�2���"�%N�,ihg1n��lN�w)��<T&e�JŔh�,�eK:ũܢѷ,�-l[����i�QHKգ�R*ngXn�N_d�]��/1Λes�Ú���*@�-���B������!-��f��Ԉ)=�q��(uYKX��?��@Aά� �9�eƳ��l�Q��儨���}��A�r���V]���udp��x0:�����'ע��l�S��qޭ�pm�[;����S��c'%�2Ʃ�����q����y�l��6b���X٧!b�Ϋ|�IsC��l���SX�Л�r	�)�7��E���9/g����o�E�<��>uq�sp5��*�Ν�: QVq�aY�4\[���8]�-	��B�%AƄ�}[��}���F��o*�Q�Y�=����IB����Agv�ͬ#�D/���,�G�~�˽� �ŵ��$7e�˴ֺ��Z��ʵq�웯��V�q�ꭺߕg
.�J5���F�m>ތ]u>��,�����ynҲo"X�H�|:P���<��j�J��ˑH!(��{�!���;�%K���KWw<f]pįt�Q&�L"D���xv�SBNѶ�N���w�|�|G�{!݇T�v5$M5@�t�U44R�זZ��O6-Q.�A'T�.�(j���ҕ�h"<�E��Ӥ�����zӪ�'JJ�: ��i����F���R�j��ւ�����v��o.�Ҕ�T�V�$���U1P�h<�"Ѡ�(f��<�#A@�Jy�gITA��4�L�&��ct�b�)�a�e������m�.󃠭i��A���ifX�i�5DTJP���j&��bO �M ttn�K���K����h�]٣�uI@R���%�C�U�4�J	�e(
������BP�4�T!�izt�E4�$vN��B���(
�
�)sň>y���q��QLC�՛ږ�$�T��5*��4��S-����6	�NT�+��vB2�B� r�>��3^�y՛܇W����쇛9[7\񿸸Q	��Y�3��üz����d��j�y�}���2=��Ջ���K��U�+^��&caq���A��z�Lx��3�9�(��MI�x��"n���}�x��}��h�;�:T�{>wbUDgW`3�&l�qn:d>��X�k���;���ң�=���ܱ�~�[ޡ�|�n�2�\߮�%�d�l�;ڃ��.�T��3�͋[�G��_c��=��~7�<2�w��i˒�z�� +����\��oO�d�ir�i����>}�#q�|dF���}^�S[r��Cs�`''F��RPe��g�Hy����q���qv@�ɷ雈ɏ57�P�z�7���9��'E_����In�ģ��k</�bj42/�0u�U20�P�>���v���������82v��~�7t�V����9%E*��9W�'k����ί ����v^���-�ӡo-���(���Q����#�r|�P
�d�s^���KF�1({�+l��m3<Π�.�rc����c5�Y�at.�]'�+�̸�+,#Ċ����j/��-��1�� �b%n�8�k��{�qU�d�f�kE��ٳ/lmu���}ĪC��+-pZ��!;��g­��T뛺]s��C}ǘ��v�t�T�+~�o�"�{Vo�c��6�Uê��lk
]]�	���^6s�79'�*��}o<n&��A������轤F���Kh����#�$Jy�W��ᢡЖ*�Ѩ��zʪ��9@Ty�D�S��L����wnVY��o]Y�]�ȨA�B��+�u�q�C�̆)��r�N���R&�\��%�d�ObS�iz}5��܂�ԼER7�X&�z$|�]�ȓ��_C�T��o��L;�A�f�dm�,��x�j��^�K��D����W�V۔�s��؜+\���q`)u���z`!��;�, g��W2W���ӟkʍ��f�:���V~�A��"֯�`�k�i�@��G��ׄ�L�,��gyGO������t�>��Vy��aF�����N�+#�pp�חB�&w����,L�"���e����'�Hc=�U��^T�����}��l*>PP��NnNVz�4��;�o=�6=K&S����B�i��¿"�"8F�&|���uc|J��C�c��8;�%���Q�y��ɮ�q�q�ؖ�y�}>W8}mn@�K�`��;F�s����=�/E��v�.}�X���^�-�6�-�J��W��_m��&�Vk�}xr�.���2�7쾡���e��B�I'[[��m[�i�T�R<�Z�-D�t(<n�erѻN�˽���r�]�n�9�s4��(�I���VD��K�]�ؔr��,#PO��K�=�5�嫨�ww���9r����=e� =UR1O;�/&�𛌖ʸͬ�/���q�g9����ݷ���=�׆�G���G%�pKGK����K_�س<�)V�x�����ϝ*Tvi!V+����x:ZgC⊟c�=Q~��"�������D��ىA��H�}�ܴwkڃEEJ�z����ר?yW��]^�x�=_��<�]������{��rׁVb�3�X|��׷qMǙ���0�Y&
�%�G��	���U���-ߪ@S%��x�f���۱���Ce��TGz���ɓ_az}�	xk�Ba�z�^�'�x��?NX���bkZ�(��U^�o�T��B��'��Ox,�������@�=-G�j;�c9�q���;$<F/rtF������+(
���fE��D�g�ꮿög0�����E���Q
�d�;�*��½��
�������?+S�~26_UP����9g:ۆ��ih��Xi��Κ�m��{��u�&�m䔯�\� {�>~�S����E�j�m�!{�C�0o�6��n���_lM+wq`	�T�X�Ӻײ'�$=����N��"�ZU\aE��X���W\d7Lb1o
��+�sv��u�o_��'� �L�����Zv��\�{s]���]Ϫ-�ձ@w$.��{y�n�|q�_t��fcƳ�����<�W��ސ19����^O���9�hc�<4�S\��ݽ�h��*���;X��ee�xJ⧢|ǣIr��	�f\;�g>~�hg�QF��������d�w�w*9���5�AX��
�or'	�1ѓ>Ns���v)'*�|�[�+j<��͙	�k�F�8�p��_�Ձl�(9U\��="�m0���M�z}������;��S/��v�go���_����d#�Y�~�)ˠ*�o���2�x���%S�Y[f�sWr�tZ���������W�<��%����8[�T���.k��^{���N���̟��=5z������(�OqL��{�EE��ȸ~�M��%��@OgЭw�`��g1ms�n`Ȃmzv�j��L>��3N���7�xz���9��������Ve~*��0gVw'��	~#�;v������v6�<5�5�Q�_��_��O��*���s�Ub�k�I���@�uB_����X�]Duf;�4.1ϸ�@,e*�}Jc�� ��U�3���[�E�@�[s�0S1���慪y��EDÓ+������1��{��ݯ��Ի��T��1j�^ϟ1�P�B�r��n���e�����gm.���G���$m\��L�S*��������7�����I���F���vb�*�
u��� ��H�ݕ2��70�q����?��R�u����W��T"·��{�ٳ��T.*]is��uqq�d*����޾]�%G�p�~������ S��R*!���ᬄk�Ŕ��qOE�Ee���a��y>zpp��鋈S'�S���\{�C|s�/*��a�^t
����p�Y�%"��kʷ'�}�x\'*��/ǧ��U��qS7�.!*b|n6�i�j�n`��x���`=�ҝ�Գj��9�A�����:�!�9H� �S7�k��	��7^�w��L,���n������]��=���R=�%D��ꈽ�W�p���21��#�Πlb��2����	p9Z��W����O��nr��}�d�r#յ����dm}���:��ϑy�!����I��w�>�|=�����I���g:���ڱ��橛u8˜�]���zh\d�e��x?��f�A�.5f��|�Ǽo���t�wm��]�4mz�p��%�C�@7��6 �kds*|Ϯ%W:)(��ow�yܦo&|9�\�;�t��s�{#}Lp������S�Yy6Kr�GfE�<
��Y�%(q�OyV3�kZ�L��k��(7,ܝ6�r�t�,ŦuO��q�;�^g���Ӆ�ۻ�Y��w\㋏=�:xp4�g(���s;�E[��s�ok�5F�kQ�ި�T�IM��=!<���G�Y�s���jOQ���|� a��0�K��kґ_���NI���Μ���'tx�"R���~��M�(��s������yތρ�P���yM����'k�P�����x��Q���|J����Y�N��b|��Ġ�+l��z�Xӎ��߁c��up���y�D�+�o�u�\��>s9�ʜ.|���׽W2@��ٯ�U������M�>�s����jTWb�N��9�X�l׍�!znT�oِ$���*B���	���|]�����Y�U7�ϽKZ������cE*�B��5��g}w-�T�k&J��`:�Q�eḩ�Z�t��<����pՖF���U�UK�>5� �z����X3�*���w]�%s�Z�}"}�8��A��N�u��T����1�6��;���p��>;"�]��1U{'�;��.��j�|�U�=�Gҙ�s�N �����Oq`Oʝ�j=��g��d�āsU:Ex�o���M[��߫��F��E�X���w��~�A��"֯�`�k�_���+�q�v%E�'�ML-w^�YjV�X��n�7�v5�s�6ŠeO=��!��x��g�e�vK��js86oq�<��X�͋[�Vβu[�11�]C��t��rnP�լX���ݞ��*ʋ�T�=�pR��3EfK�L鮨jM��2�1t�|�gV�Q�A-��йW�V{����e�N|��_zl=�.\=�O�O�]Ĺ��/����0�ǲw��:�.\���� r���xozhl&����^���{��2<�>u�i������z�:��f ŏ3�c��ݹxg��X^:K	�ҙ]����S�{ʋ*�x��h�\N���o��ǻ�������Q��ɴ��W�ٕ�|�Y��{OG�>�}���y>��*�L:��}���<)��G�P��<� ܛG�p�R��w����>�	�G�y�����]��{�4�w�!s�,��eP�=wCo��zpa�HM�O�G 1��j�v��]���x�g�5��5�\H���
C��.Wu*l��%7��2.iUh��v��o���|%�W�=ŋ�v|͟N��׀j3ِE[�n�O�_F̀���0/�(�o�%�>���z;Ѿ{������i�j:]xT�� �������cr-r��~�t�]��0��0nw�Um	�\$��Q���`��	�Q�4j��q+����|�A��qTn!d�m��401�nH'�r�V���[<�sn�R�}Vs�V��2��gAy̫���	�L�Vf37
a�Ũtn��,��g�='n�Ka����wє,�0o8���6j0��J�]�U'\M߮�(\A������ɣ��)���
O�>�^���0 d⮍������9��R�xx��tO���fF}��?�슮�ò6�t�#g�7�zx��`�!ӵV�ݜ�Z��q�~2�&�׃7�f���򼘸~�+h[�<í�k���!a�=����d=ۮ��_w���.}�?G���/��*�t}�w�q����'�YNv�l�F�s; �Y����j���o�y]g|@�tux��	���e�����Ѹ�v��i�O���z�ɾ���u<���H���D�FL���	������P�&g"�����<��`��amӏGh�P�z���y�b�]�����M�ι����s�d7}�P���E��9|o�Qu��|�_���q�����+{P�ì��+��/ܛE�%���M��1���̀0]z���r�
��y�G���KS�}�>0��U�v{U�WKD˕�=�F���W]=�~�T���V�M�3~j��s�{#}@m|�~����U�ƒ���Tv|��hﾅg����_Q�N�]`R��e�#�JAÊ�$�9�{1�i$o��;6u�N����[�����{ru�V�JwwX�$Wٛ˅���z���Ҙ���R�j;��y�O;w�?K����Km�,�m�j�|�S�t����R�֎$�A{�K�EZ���Y�����#7�O�Y=Ņ��6����~�8g�Ճ����;��[�sb���t�e�n���� ڟ+�����3s��ƾ��C��k����=p݁��3�dOy8���k�)��Ԋ�I�(z_���ϕ�ʫn��D�~)`O�=ӵH���ʓ._t(�T�,�Kݙ���R=�����{�M]�� t�v���}�x1H�qQ�6�`�HChx�5�,��~�SH�����n����$�TO����p{�^������k�s����Jۧ��5�S��<*=#�dy���R�G��L�8��_����KL7�ީ�,���ܑ��E��*>��(��)]ׂ$�5�zO�鑞!��P�����}R<W&����evp��Z�����ŕHZƝ=3+�S�7���®�+�=s�j=�X�Eա��@��̓qi�5��f����&r/Ԯ;#�s�XP�iP2�P�m�p�F��s�]�S��t�h�+�y[�X��r�	�>V�ʄ�.J�.mDgU�7Jf-q���4j�7�'�,��jd5I@�Y�幮Уھ�v\�t��/�~�o�=�yW�*���]��V ��X�!�����{H>�S���e(�e�5ά�x�㓱]w4��V8��㖁�[�-k�OD�77�5�a��s2��I�]�>�g��T ���z�&n b�[v�t�?�&e�W��b��idj{[�qȠ;�8rG��v%TFu<2.#&u����-XG�5��&Ǫu�����o_����]O��M�F�~�(���eɶ\�z�@�����P�o}Uù��y�����L��V<��l<�=s�<3�S��v?
�nK��X�e?Ny�J�]x��@�{V��\����,4r/��9H�s��μ4TD��lq�(��FYfy��$����.6���y�ԫ��dM�d���ܨ��x\!��੺�c>�㾡�\_4�����/Ϋ�Wd�����=�z��D��B{�yNwL=��q��#=}XL�3>=N��Hw�O��:A�8�d~�"~wT�l�%�h����E+�;S��3��(����>��&������Z�u�=L�e����@y�;�$�BZ7����B0]��e���U���������rχl.ܲX�F�F���'�mO�w.�&j91Q<d����(���W��
[�����[G�/��m�t�r�i�
Aax�/������s�G�z�N��3��1�ُTqIՃy��.F�B%��WV�hc7��	�zC\쭏!c����Y�${��1���lI���tL���e蒌�438u�w2�^ՙ�hSB�>B�z��L�E;{��!� ��
=�w��!�z�g1��9!������Y�}�o-ބK��r�G��2��/3g�HQ��B�v��ٖ���t݊�����ڎ�J*4�ȶc��;;x�u��vo4w <�A�X����Tn3�2Ү޻:����0Ԓ�V"9t�c-�o�Bd;I+c1sn��V8vPX]��0����;���GDH��O+;+zvЬ2�����G/z�NP�K&p�/^�����%��,�Fl�=�i]����;(P��Q��˰w^����e�q��w,�cshTܪ�x*x:�)]46�Z̥ 9܍�``�&`�o�'x�o(^XBL���Nt!� �JC�]�j��u�����4�4I`<���PJVP����4��r�jԏ*�&�EK���-��E��zڵ��|(Q9˘j��HJ��Tn_P�k��j]��=�=����bm�X��h�4r� �O����ܸK��, ���Ւ�����c=���T�w���[Y��M^��u���n�qq����b��r��y��`Yl#�TuՋB�7����5;9�%��u�j����s���[5c/(Q�k�L�grj��ٷ�|tc!�S�HҼ�>'h�6>�]�)����,�3N+�V��᯶���愾�2��ʀr���%o;">nf;:�9@��
zl4���;��:��ݶ霍���� �l���h��㖊ŗf����-��9�ݕ`�f2{�X5CA����v,�be�����Q��:%��R7�ݛ�� ��+�VrY�"�}��8�F�"LT3�o��^F��A���y�B����/T�����#��:�`�Y���nh ��!Y�˸�z񠆃y]x1����yM<���0�<����eioo��ׯ��I���i���2vQ��s���WW���#�A:��aF�7�H�f�)�cj���K��f��Vk9�8��b{C�Aȹ�C�Y�i]l����%`uh�Zg�;�4G��B��܍�n��b�i��mZij����9�U[*����|0[�ڷk�䲀�o,�W��MX,f�֕�������t�T����/���1>��.�.CV����o��	W^�*�<����M�-�NO\ f�ń�̱Jn����z���,̾6;��˔l����A�K�lV����J-�m��"�4f��q�K�n�I�nr����I9*p�-er=�Y]���g�\�VR���L_L��f蚎��$锨��j�)�`�p|;���wY��iu0R�bmcR�l�;]tm�]�<�h]c71k�khP�莡��s�tf�ֶ��O$m�Z-���[4	��غ�v���}���ȕK�L�n�P�����$`����{/���^횾��˼���46���p��t��r����d��]�ׯ[�����~���M-#%I0���;g��"��C���!ם�"hv3CT4�T�lTAv�T��u���""�J"�����y�4��톨
	��Fڶ�Aшb(
ge��i�iC�(7�2��N�k�	���l�T�+K��*"&�+m��CT��t�DJQE!E.��!@Ĵ�=tOF�.ى�j�ں8����Jt�D�����IAE#F�����i���V��$кB�� ��*������t��)��*ZB��(�B�톂��PP��#���&]:�ĝ�Q]h+݊P���z4�1&��CL�h
�&�����7g��7��.�[�z���Թ�ΗOM,C�<�l�]�xvh�|�~{���
'e���]�R�:����-�.�kR�N��4�g5����}y�s��f�>Y\B�@�9���t�F��1lL��]�;��{���k�D��g��{�_L�=�d]Ð����[^&��sӱ��k�:d�Ӹw8L��q���;0#�I�/mK��3�㶩M_��y7ʉҧ>.�\:�r�U-!�B�Lގ�u�=�^���V,��O!���꧝03ʽ�v�vk~����'P�fpwz�NW����dnOY��H���]w�Vm�r�`_t���z� ^��N���/V�-��({�]� ���wp08�-�qw^��T�����PD�Fz@^���m���Bj���j���������bP����mNN� z��M����k��x�yf�C9�U���܊��+��g�x�t���V)zS+��#�j�\�rx�����m�V�s��G�/|�DS�.��!\���m9�C~�s�G;Xo�/�q۞;,surg�wU�G�9�졞����r�_{)�	̑�<�d�>y-�y6=�ܒ
K�n��ʶ�_QS����OF.2�Cv�G�S#� )=��T�m���K_�غ3ς�~/B9�{�!��g�%��W'{��۷4v)���V�r�� ���９�b�*�r�E�]j���{ד�e���n�w>�\�i�{9��(����]�,�Zi�cq;cy61� �7� ������0�WZ��oEf����Z�z��ݼ�]D^�K��)�\�ۧ=�W���ǅ���Sq�@�E��D����*��x������tcq��#�`!����[��?�~�7>Gw`K��{���G�����g� ��t�����"���z�!��jm~�5���.��U���d@�Y&;GxO�B٤F9�r�π
���Lp��s�-3��(&� yU}j��/�;՘�d�az}� ���P�u�4iz@^9;{�ZG�%ƵܗO��}n��[oȩ�F|x���}O�M�-�O�j�u���z�pTo��],ص��h�ǽ�%�����d��R̋�މ��eV���*���G'�E�������؎ۊ�CG�o'�.ݼ�NuX�-�9I�̘�����#�\:ۆ�9����5�]ؼҌ��=��T}r�M�ST� Tw������_����o���q�o�u��Ј�v�s��i�}��nh*�t�T�Q{[P���+7���x��	�S���ϴ��G݂xb�`�ڻ�F+ܘ�������zx�}*�iS��#+�D�d��oK����g�o�@Jr��S�ɪ�n~����7sT91{]�Ů�-��ט�E`�n�91u5`2�L@Қm�웙z)�Gr�w�U���rtx�wr�]�� 2T�G¤Q�bn�<{p��].uvK�ָ@���WWϵ��a��B��\����jv^�g"�Yv��5��}���7�kF��U�[yq+&u�\dϓ�6��ق�3���P���D̵8goZ���s�u�gҕF\?m�����YL9��ڙ�u�M����;��(S��8��:��v��75�w��B���z���f9�O��r����
���Bͼ��x�1��9Y��{wΰ�4�%��R�}]{�o���~�d1������-����vCǞ�r�חb/���zum��_��O�W]ŋ�Oq�燞o�~�r.>~�Mì]�܏X���Qޝ�7��x��DzdsCn{ۘ ��+&���w�*����A��k�]��O�(��VUW{[��=��I�x�k��WS*۬�_H��@v
�=�cfQg����&�d�Y�B��mx��>�:�=�n��B�!��zn��lEu��c��B���v�o�̈/����]�w�eS��S�鿡@��!��H���7�A�W�8{6pt�qxf=)M�~/cb�w;g)��?Vʦh�ꊇ��J��C9py�5"��e��A��h�ӎ2�	�^�К��#���8�H�9n�{��t���)J�[��j)��2�_VsK�GZ*彥�<���w]��ې(Jڥ��V�p	�d��]��`4%v���BJQ}$��z���ԥ�v��G���Uѷ����v[L#��a�s�g{�>za;�����3_m1�P����L�C�Q�z�l����P��܉�{7Ѫ�W�W� ��ݚ��r��>��!���ŕH_�6zn:�Uz�.�x������V�q��\U`����B��j*�{G���R��is�"����G����`g�qp6��&<ͱ:�i��,���w5�Ӽ�5�}|��x��^����U�1�q�'=1��q��e�5*=�C�߭j�zpUV��(u�e�<��������</��P��N�TEەfE�������˳��=�o���=2=���b�^T��;�?NC�WY��ao��eI�\�z��s3y�]�:�k#t�l^���xT��;�xK�{��es�k�c�>�C�!N�q���s>�k��H�ZS�O����\l
����+ǲe��Q�j9�F�:�kz��Q>^��|��S�:����foyb�|x�zK���j�L�3~�k ^M�L�d�js�a�/RGC��u�8蜰�"e�몿f�ɏ�?}������zKφ��0S;���m������O��󺡯@���F*��$Lϙ��QX2&WP��u��RB�ݻ�{H��>�2�x���G���Ҵ)+�0�540���]�[�T���S8��@!<�xnS��Zo!*J��ium�K�)�ʋY�'��_?j�W��=˅���I��f�:fo)H�t�����&wv����?�d�bt<}�u��ˢ�||'��F�J��8��MϠgW�W�����Uc�>�s�ߩ�C�}1�}>=7πw� EE�0&k�'�-�;/r"��R��1�V�ۙ���y���8l�w`9�,
�l�6}!zJ>tC�d_[��p����m�C�}�,�gr��T����㷙���3)Hr�6�T�����bؐ�������Ǭ�8z}7�wP^�2]*�䚝�W�X�;S!O �6������c8J����;ԫúWu)Ir��3�c�ȝ���x�&t�[�'�2�E���4�L��o!�^�8�X\s���OJJ��z���U>:J�����C�F�����u��b�ZB94��2�Y�Sq�*�o�g���ˋ����e�17���}�*����!]���8������pY��8/�gp�b����}� j��o���V��	ϩ׸�~���e�x�>9��wIP�N�@��|Ixh�6/�/P����Gl�,���9{��3�4ɪbeϰ��{��1�Mz|H�z���4`\慆nfY��^r��f�F0bY,p X?����^�|��$�5�T�W���C���:bt������x����� f�u.�v��B1�5z`K�$����{y�..��J�}RDC��S���&�Jup.�#���,����N��}��ZC�6�鰏y��_={�W�S7�>ǉa��x.<S+_e����Z%�7hl{S�����ϫ�}� K���s�� ��܁e�f��2��\�|�Y��K�X�X~k#D{��4�|{aX������#�Y��@;7�@>�wCO:�,�>��l���0>��]�c�sП�����>�q��~�{=��˓�T঎3<��O��!��C͋�Ay3䟚�f�s�����JG��upw>��ק��dw��y=��hh�3lĠ�m�j�X��pъ{�p�,��	��Y^W��nW�w`=Ǹ�ӳ�o�ޮd^����M�j+¼*͊�YGc��{�+���;�]@�~�����6ȉ1�+\�5�k��qs��z������5�)��WT�4���*��O�� W��*ٛ�cTVНv��FO ��;}�Z�Q9Y�����f��|�xY��vϙ��Ϥ�+��<,Ԧw+�|=�9��#�*�y����!C�ޝ��t{����ĝ���I����|P��Ȑރ��U]�f�ޏf��A[-�т=�,��Xh�뛡| ��';t�ܽ�'�ɼ���V��X�Z�q	�ֹ�_�I�f���(v���R���:{[D6����T�,�	:�52/eFp����Ͳ�j뚙�9�Ku{#���ˍ<�&�ռg�}ˇ��z���\1q
G�2�;�f�U��1qϐ�o�|�n�>�x�`b3ȗ���0�w��X�q�i����3�xL��v=��;��%m�ɸ}�^����o[��������.�^�8/:����+�-32��ә��fs=Ռ��C���z������	b-��G:TjZ$<����n�qs�GV;쉼��MƗ3}3��z�L�ec�������j���zҊ���ڭ��(���e�:�
��ށX��M�ι���&r8�oVN���K���ǀ���;⣷=C�i��Tq��n�F߼�����Pͺ�a�B��*�OH�ɴX@{�`�l��꫇��#�}z])�׾�(M�޾�s�7�W��4���^�p�P�ހ��*GMM�6��[|�v��@�;���O�Xhy��x>s�{#}@m?_�<1N�p��[�Mpb	
O��s+wM�崛������|��˖���>^Wqc�ґP�;�X*ݫ��=��z'��V1��J.f}�72}9�����r� ��U����ݨ�*��2�m��=Y�*�%_����˅S�Z+�{۬�Ǝ��&�H��p�^ʂ┗ݜ<6+��IB`���k�݋(��,�6�'�ܻ[e+RK|X�V���t�+VԲ8�'rܭ]������8��R�8�P��q����s��`a���4I)��pY���"�eIn����Jg�6�����F`�R
 ���~ؕ*��^Ml�v5{��t�3Ro� *���U��I�h���^==$oFc��B�ϸ�/�{�Eyz���|s"{:���Ba�z]zbː�%@�|=t���āJ����h{���>1��,�@dԉ���2���I�G�P�\u1����T=qg�/M���]p�?Y5"��G���>���:�G<�OI�Z�zk4��ܯq�����m1ધ�Y��'��P�/*ǍZ]�2.��H 8�w�!�g�p�F�U!hsn#��&1_��
��%��x��s�u]�霊���n�wZ�o��|�V�-��ȟ`≛�J�YT����T�No���o{.�C������q���zu��^R�p�X�o�	����lC���W����\eq^��}�]��[�H�q�nTNx��3�A��=܆��xWc�C�ߢvp�㧆E�<)0�=��w��OM-�.,��i!ﺼ,&��u>^�:�q���F}�L�:�eΥ�n�٣w&=�l�-�hOW���NXF(eR�#Y���nv��l���ڑ�ˊ����{��zI��zA�e���(w���i.S}c��n�`��}З��\nS�m��Y1�J��sy�kI��]/�U�GtU�V!�3{ �x�Sk����7�u�\��.�R�����fOK1�����hlf�SG��c�*�����כ������$Y��f���ڗ�T��;������˔��EG\�;��$o��.����*'�q^��Ǟ����[����~��O��ޙ@>��\���.ԿY0ڛ��ʇkԑ+�,�+�1f��aok��`o\V͵n�ȃ��.���9޺��'��̀m�I�-���U˼"�%�U��AG��F�ӎ�D�l�{�EF9.��e�P��C��Z0}=���U<v�';&]�4�,u�Nn�u%�x����y��˲UxŎ,t�s��{2_�W2@�PZ5ꨤ<��VR�s�Ǻ�K�ޝ�qn��WTo=>����T)�>-�Dx���S����o<neu�^hP~���˞�XX��B�Pz��YDd���Ҧ��2��2r�낪��Z��#�/^Vn��B�Ϝ��<���W��U�C��DUn�=��������~*�Xϔ����tO��Zg�n鬋����c�t�w:�m��3R&��x�95���7X�NWM�~&M}��TD6�dԃ��� ���U���ܪ�IΑ�c��+M���<ϝ�ro�lY]W�Ky�n{�y��v�����V��`A6��kR��&��*�H[����۔�a���F�Q��VJ�@��a*�N���S(ot�4�w�H6V�aF��v�_;x��smwv��~�8�r\�����%I�~��~TH�0�>��Ӝ�T�e�#�H_�\q2@D�E��<ww���p+����ޜ��*=�!>S[�>,���9�й�]����y�3;*ϼ���
\v�p��N�jG���`	N��m:���x7��|�[����s�ϙ�Ֆw��9溽���]��P��м�����T�6��x.�&�ב�B�[=Ǻ�rv8�-��7�A���*}�+#�q�Tc{�7e
�>ǉa�����CoM����N�j�c���
�^�kh����-At�}*���~{�/&ӛ�,��ʆ�=�a����;�'�\*��[+��ҭ߆GN�G�#}@;>.@z��a�Xɴ|'�!vyNT���j��V%�z��zly\y����-&e��:�`t��I��L�����W��/�g�{0�������_ot�}>e\}�\�W�C!zQsg'�Ҹ��>5�h�}�<\�l�z�'~�Rn��Mމ^��0��x=���ݿ?��_+��<5��A��APO��*"��D_�*"�AQ�*
���PTE� ���*"��PTE� ����AQ�UDW���+�_b��+�_򠨊��DW�T_򠨊����+�������d�Me�D#X+~�Ad����v@������xs�J�H�@�Ȕ�
�D*)D�J�UJP��v5��j���%
����H٪f���ͥI)H�TD�v*$B�%I
�V�,�QZv׀8��j�RE+l�0�H@���@5�d]Tep ;  �  =�챢ZJ���E�J�
��sVSPa-0��l.���
r�� ����P�T\�� �2���c��v�Iv�Hښ((�L�B
P5��2���b��"� ���������[�Zh"	H��i�h�!e1�R�`�FV�mB0���p �Ь�5� ���Mel[4�a�J4�) 8 n*�Ac)-���)�a��٬SL���@�)
��W�Z�U����%ڈ @�
p���´H3ZZ͵��Z��K&�]� ( ��FUIT�P� ��A� E?!�)J�OI���A��aMi��&�&	��0`��5O��ST` i��i��&&R4&�b�h&M#M����S�H$�D�U&��bm4&�bi�M�`����v�V�.'[��蝸K`
?	%��� ;��B4TEA�" 3S�@�ŉl�?ُ��$~���00�Q@%x? ���� 
$#%!Q�{m�YV����Λ.T�C>S%8�3o�C���Ǡ楔�.<=�_~Ӫ]���彛�^��l�n�u����@��)�U`ɶP�kpnm��"L�M��v����qP{���L$��ȑ�z 6Z�!xtnR͢��ZS]�`[��^eňQ��#�D0�S��gE�f�K�V��
��,U�&�"!�+W%����P�U6ܱ�b"E7@U��&t,ߠ�.��-M��×��(��9�(E^�2��.�;M�Z��t2�	Q��Th�������e��af�&ؙF���.��Ïwv9M^-"��- @Ţ\�UҀ�Ӵ"�F�PYgU2`����OF��`ofj�Ӻ#&�,-��mZ�7D�t��J�(i���Iw�-�V��kx*�Oe� FV��vu��u����㭸v�W���m!�v�4ȭ2�ص%Rb���أ�WEEfJu���WUD���PUG���4mҭ�A��*�c��X�䨞�{YV��۴�U�V��J[�Zjmk˙`��X�>��JӸd���� �:3F3�gt���g��QÊ���a�A�q��jXm�n�V�9�kp��t�6���U��0���^@�I:8����Ç3s6�+.(�@	o0
��Qm�V�]L�M?�FK�Q|
w"�dvcn�MT/nɂkƱa��N��4�%�[wA#����Xh[1I��8^���i���6\N�]����EC[b;DM�Bϖ��]�|v�
R��.ܺ�`�X���4SYzn�])���0�KwZݽj���x��p��s����hC�̨���@:CďR����'9��w�k&�D���ö)���U'̜�i�*�ܺe�z�Ĳ�c��]��mړH{�U���)mk��$ғ�g�j�.�@ٱSJ�Ƥ\�@�%F��$-a�F�� �Z�Қ�[�e0���[�`,Jن�Z�Z�P�T35"*�q�w3o� Z��M+9h4�� ���mT31�f5�+ , �]U�%%�A��Kkl�����r���/i�D�*��9uQ�.QPF	"��S�N�[5��hY��ɵn�D�����Њ	L�7]Ų��Y���e(mی*u�l$Dx(2hI�#u��4��0[�^�yp� ,��XÓd4�uM�j�u���R����o[;%��0e�ȡ���ǳk[4�ܒ��@�4�,@�M��ǙD�!��7�[6��ܧ{�B�k˫�L:��`�I�����*�ܬBGX�V$U���X3C�q`�y������Sz�cոff�N���*^яe(�ލ�jd�-i9*�I^n�H�(0��+~E�ʹ���b�vlջ���8��(�ĊWmac2�n�ڗ�v%%z�Z20�LE*��" ���oi-�3��Tʊz֤E�Sd�|�dA�,����.��bV4�!��:ܷ�Z���H 
tK����x��c��^6k*:�i��f�{)4�n�
�_n`�*mS�u��ŭ�T�xn̓E�ո(Uݶ�KSi:�W��cJ�"e]R��v�;���x�BG�9�C4+N���E�U��p! ɎR[��=4vA��i����Q�qZ�Yq�$[aJ3�j���B�ˢ�m�B��%�wT�af%����Q��)��^��WN
Jl�t��C�dm3ed�/�]Ȯ�Kv�=P��^��)�
%���{7`����o0b�ꅷ.�N��;m6+!;�f3�*��lEIU�t�;)^&k~�X�0���2�ئ80�j��GM��IZ�tr�kmJ�Oh×b�5�٦�r�J��s[�Z��{��e�^V:��F���|�&�szMn������1�hS���ķ-L��(��P9���8����U��,�&*�I�0�ST-:Ej��v=pТڼ�Qu d����_�3Ad��O,�s-Hֱ�/ok&������5���S.�e�)8*b�*b��iPG'� �H��0P��.�^��(À�0UZu�m�����5A^�*���\d%��s(�fdю����+1��Df�:ͳWz�6~��i$�B�T{A�����Y"�bb�t�Zw�Y���K��c"Y�M��En6��*��re�ccwWٷ��X���xwv^B��ŰZU�i�Y��A�7r��qu̱%�iR;���djVHC@�q�pv��.��6ō�j�%���n�Z���n�p�h�*�r�#���)��k�&+�n���V�� �M�'q���.�Բ��9u�Ү�\���Mw�nn���}�&iN�n�����;�����(|^�v�l�f͕Y36�K^^� ٨�7��Iz1�p���P-��+Q�ӣ�dy���8��t�:N�v�e��Ki��l���V]*�0i��2���m�dnnMc6�Xy�T�VEj�e\�X���E��5-��*�wt����SئBvi�ձRI��J=�M����D-$�A�h�T���?`o*d�2��VQ��֏�0�[w�N���q�Lى��#Vh�r�l�;e�G�;� �g&�Ĺ���XŻ�ՏM���IF3��⽭�Q�ɢ��M�+X�Qav�LxM�	%����:Dlk̂��8�,�S@ʼ��q�mџr�v�"��/T��q5��Po3]�)� rּۤơ�Y��&�y���F��ń�"�8.�X�.�9�����*@��R�tJ���fj��,��f75�(�R�*���4^*�T�4Z����+��F�����k�e���\Pm@6j
/K��&��[J�b��X2;��{&jD�T�Zf<UDd�"��.�v��cT
���?�����iБ)��ڤui��C���M7��K}~=���W���w�w,��*A�u���i�c5�v��q�a:��#�F�V烷���ɻ�g�{�4��V����(YUʑ�k!�Be�ͮ�`n�^b�7)#�f���;s�+T
�G!�(I��:[x��k�n�N��f?���<�0}h�̍�2Ɗ�Sޘ7p�ƙ�e�=�n�H"���+��^������<g��h�X�b6bN�Ky�R��m��7�E,=��������4H�\CV�je��)�f�����A|{R�sWUS��c�ٰܺ��ֺ��v�����"�Em��t��#���3��"�����݅܃����F�u_Ň9�ޞ"R|k�j���Ng6j�#G!�\�m��U�{o�(��K�[s%�LZ����^_n��Mä,ʕ�-��нVޣ>UF�J�J]���*�%�9&��m��X��i]�9\�uq9�x#A>�^���ꭠ�6��
bq��1od*�r�"Ȩ�W�;G��e��q�(I��6N�(v������o�N��g�����7�Mx��t��\(��,n�Ge�),�����b�/���N����Y&���]�)�s��]Z�ؕ����\�b�s��;��[�[�*J��x{^����˾��T�c�1�9w��viw��\u��54I�
TZ��W%/6��գ���zn\/t�r��t)k�l+yePT��䗵u�n�rY̺��P!�>\.��YhuX­|�m�0z���\�v�o77����5�}�}*���e�h1pdr�P���-�ea��P��Se�U��AU+�u�q،t�sY��|�H�J��U�e㨎�����Ojl��C�0���i��:��[M�CE�r�]��ƍ���MۇJ����5�K�U��pr�(�[�6�-�n
�գ��-]k�>��o)��+�T-s�*�W��v�ؚ)	��ܵe>�����%�6�w��)Y�䎁7}11�±���	f���̐>O9fc:f�[��b�=�9�f��5�<��}���L6g_C��c��Q#p�y92`�;�����:���ԇ!kF�\.�q�ٝ*v�����=�Ȱ}��%wùXF���Q��u������L��j�A�JUU�u�Uz]e]>�6�=.���U����qZ�w;�H��C��9mj��Cs�/@ۧ����W���b���ع7�O�8��!ˣE���W�b9\4�58Ӂ��Z+)0��_oP��QpPZəK7��	���(�ݒ���9q)k�u4����%������5xxs��nJA#ӕ�Yx�K���:	��uՠ�ǃ���c����ܔ�d頄�6�Om.{�1O�%���u	;��U���ȉ���o��k��{�E�pa�qu�z5����:����C�6;���d�Zǻ�Lf�9�jh���lꦌTV�f�x�
�V��-1Zt�ú�c�3�ڶ�l�Ж���[���d���d-B��c8�f�x�
T��?,���j�1e]	����s\�.�4	�p��6R>2*��M��h�u�5^�}��56ε�cfYg�h��Ũń�Yo!��zP�Kol�o�+�_������wiN�\l��Ul ���2��:G_
,��="�%��o����n�2��*3p��YCAz�&5�ޙwBn��SqF/����nv[k k;�b�h���kTR+��X�C�ͻ?j�N�agp�WN�D�/g<��ݾ�/�wB�=
���+-��;��˕w
���Ӕ2ĩ�=Fm����_G�dE٬:vf�E�h�z�G@)|���C�1AAq�����r�>���t��8��ɭl��[m�urj���R�y�2�g�ծf{���5�M�q��z��vP�inulwwFIo^f��-�F+��}�a�n)O����l�j��G�q�.��=�=��%/�-���F�o/|�V�5uN�1�\d��`���R�W����֩1[����1"^�B���s�؅��@ø�o<�VO³Z�����e��8�����Ё�`��k����;�{"b,��}��k�vd4��U�F�t��>wg
�h�[���"�p{�^�[y#���n�fR�cr����Y�*�o6CX{�ۢ��ޱ��_W5[�[�K�u��ٓ���;�Ղ��a�]�^���N�fv�I��[�=ۘY��Q��I*�IeM���;���+C�:��O�˼=C�����9���(VU�փ����k����E����|{h����̙�6��_i�:���y
Eg��n��K=9 ��X���fZm��c���dpWU���$�}T�C}��΂�Qj�&C[�]q��[�:��\'	�g&���W|V��>�&��n����[[�!}����L*�<M/
}��i������^�6]�W��TU�۪�ț"Jn[�HB��}Ll�� i=�k�<��١�c�*m��1O����W��=���M*E�ϻ2�sa��&E@P��l�**ݼ:��4���n�����P.����S�i�.P�,�M��q�lLd�v��=
:(�3���Um.w��P��YnL<�b��ƻF��9��23�T�8P�K �Յ��ugJ�U|r�%jp�f;Au6܊Y����MN\��2]��5�I\�Jm��:e9\غ�s6��Cy��6��fl��r!�ΈI�]1�u����j��ۙ�݅�mK|��;R�yUu�O��d��ykvF�:���*a׃7-�-R�ѬÝqS&C=M՘e޷j���{6�0ה���z�P� ������9Z�D���_1�i�fZ�X��%P��%��w��,���f���o_�c��[��(��\DJ�o*b�Mq6�:��(��:c�4Mdu!&K{M]���!��w�8��H�
��B1ݴ���eP[���y�7DG�K��n��8;Z�/T����#Y%SϏw#i�pM�gC8�u%�ͭ��>���h��'nP���I?&�����eC9�6�rVm�JK�����a�+u�CQ��{w�;n؄&�s]����=����U�1��PW�k۔�Em��w#]��k �MA�9tn�!vT�ܛ�j��i4/6�)����<�fuk�������L��)ʙ��J'o�w�7/4��Ofnd��K%�Ã� d�m���L_X N�4�Cw����S Ǐ��pm�33�J�����+d�9-]��С\ɺ��8��+Y�i��klc�)b�w����37���Oun67����"����$�ѷ)������%��Jo7�7�������/�cr�P���=U�J��<�Оމ��Qx����p����jc����vܝ���U�����DWR��-��I�M��X�����$�d=6���!�oBw�3�6�p����6�>k)�7ۅ,��=�gE	W���^�*�nɋ(J%uP�ɨI{�EJr��"��8���I.)d�s��oM��G^���C��Q�to=.�q�S fm�޺{�a2 2mKs�X=nݦIr�_g,�[��"n>|C��JGu���+&� �b[�rE \�ha����$d�ެ�/1�}Kk�f��%�K�mz�]��
��p�[�:�G��l_#e
��sE�"U3E��������|GBi����x-�c�`��1t!q��#�6��d��G<3q�]�w*��[tr�˟=i��WS�%#ED�.B�e^8s5��a���,�O�i��wG���*��{H8tm�M��ۮ�*S��m�;;o:s+I���Ʈ�k��>n\S&'�>KS�v�-���j7l��XHJݡu�:�l��B��{r�.�|:��'ۇh�H�԰r�m�FQ+�LYZA�Yo|܂�%Z�6
$>.���ڛ�[�
���
�r^�.�e�m«��V	����s&G���*���A��i�7��(":�kU��&�œ�u'{�|�58:���^us
d[�>��{�����cT���A���Đ��ɜ
5I�rӭ6�P}uIXyٔ���fq6��%a���:���Ij}V�����`�.7)s{��\���Z]�A�ŋ y�O��_`�oZA�J�V�A�՝\hC�n�.`�-3ڟu��QHt��_fQ<�����V�2���i�;�N��W��'�K)���3�ƀ#m)E;ľ�����qN{��+�;�m�V��Į�s��6�'��u���Vp#��#j�Bmm�t��&��)5�����k�x�B):�)d���p�+\ǳgTJ�\p�2R�"�;��Yc&l�Zm���ny[���z5Mwέ��*��c*�8�V��g2vM\�̪��BQ8�y㯣cy��m����BB�-f�D���|�1�򈻳R���)7�X��(��n}��e[���}KCd��v��2f�v�U�_I@�-�t3����Dt�O�n���Q��9§Fo�ae�2\�y�s���wM�͊��kn<;�o;��:����HC	)Z���CR�V��T�ǻ��j�F�p��򤞿�����Ku(FU��{9��t�r1�]E���#+U�!6����"����R էY{�Y���(���I�	��1}o��֫i�Ѹ�[�%]��̹5-	���À�j�$0d������6��`�1Z�Z;j���;rX�J�ruz ���ۦ����at\��4��v�oC��7=�:���L����D	��t��$�"W���R*��7(������іE��0��e�*vI�#���R��Xi����^���c�K��qL���w�$�us��k�vdb��W[5l'����7��<�tpUi����qoƕ98��T����ݷ"wZ��S�;U�T�Uo+ws�ƮB���~�Η;B�"�L���~ɅLu(K4�6vv!}�5���-]b'���L����>�wڼ�K�`t��y(���ʍ�9DQ5�u���d:Ө�{��H�+X�.�ً�ۢGt��M9� ݽU���&��,���.��^e��Z/;0dV.	*)�÷�G),�\�XGng�f�\��CE�A$B:�~���hۘ�ج�8.q��q�1ֈnd�ʸ��i��Ĝ����k>m�졵幜.�z��+�q���?Q���{��v�e���wMt���R����N�݌vKq��d��Y�<gd�_���x:Q���Ԟ�Y�X�������uݯ���Q��[�q�f���� ��fe]7��Aț���Ϣ�
C����Ng
и:�b�wӁ��T�F�$�q�j&	lݫۧ��������f��v_��9�F�n}7iW%4Z�{o8�=Q\P��m����|c�w�jw�t��;��_>��f�vXRYV(��"�#]C�e���z���	��AT+�η��[y�3}������oA�i��ʄ:i�>x���!���fΫs,�m�c'�n��6m�/�]jEb�r�^N��i��FEӳE�SSͶQr��o�ԥ��.�ˣ��恬q���j�Xn��KT]�Н��'ͩV��]�O�����WYu�=�A�՜�J��k]V֩��l����b��f��UtE�f��9FL�X�	�C1����=���_��1�o�]�&�vV��:�kGt�(�@�ۼ!��87�oK�Omj�	��׵�r�q>�Uʵ�0d�dGPl���j�Y��ͷs�j��Qgr��7oU�x��r��8��w:�ٰ$��+S֖�KRC�6�Wu^�8��=���zB��0�ةAʜ�u�(�u�
�\��J7�/jy6�"��s\�'@����`2n����&#�n�b��>'^��w�����^�>s�ma=��� ��Mբ�����]���zk"�IM ����9ژH�Le�F���2��Lu��&��ۊ-$
v\2;�\�����Gkg�XhGS3'e�T�<Ð�7�5~Y�v�dwT[�yISV�*����e�Kʲ�QӘCL�7�mN��h�m�0b�f6�q������P�2J��GPR�j�҉j���7�lb�2��M��ejiӤ+4�cX�@kJ։F�PD�u�V��X)��
��1��&��nX
(�ne1�
�)t�Ic��!+f�]�:��-;�\_�F���1MU��\���+3k��6�WÓڲ����uG�Zr/(�5o�+����%�M]A���M]�2y�UszU��n�hmi��@B��|<<̹�_P�ơb�^��;�Ah�լu�b��k^ݮڱ�;���dnk��,/�3s՛���?�Q��A񮝱����Jz}���
��GB�+Wv��Y�W:�
��~X�~7��y��㍆��V~����)U�%��B��>Tu%��J��X��}��v�O���[q�8�t�/��9w���K��>�}s'K9%V�R�,����v\�r�W��v��~j�';fM�6:JN3�c��-ﭽ��7i��=HHV����qsՇrb�^���<��p𰼼i�ad����F�{5*/=}Č��$�����%�h��'��/e�ˍ�]Ky��Qty ��v�¤�N���m�p���AKV�uj����eQ�<�o��Z4�}ˮ�ycP����)���A��0�
��뫇�-�G���̻����l����޸���̦,�^�+�/vpQ�٭qvy;�W3��+ڊ�)M�[�k��W&�%�=ڐ���Kپ�|����C��O�e�ju?hA��Q�������:�0�}�P�Vć�]�����a!-���6C-B{�]=�}�.�Ɯ�COS�-����Mn��j���R�g<'���!~��k�W��. �"��Y[���sH�f�u�5^�Z�5=�i\���[�s�;Ž�%h�B{���^^��n�0m�^I��v�
�o�%T��i�K|��<�^2j�Kozoo��D�Y�ũ%�5�D�o�!����MWUC�Pvp�:Ղ}�r�8QѺc�e׶pgP��_^.Tꓭq�y|�o��T\�;{xs׬6��^���Z�F+�F�V"�؜������]X����ڎC�r=K�;����MH�:jg��f3�ոg�gx3����7�{٧FY��X�� �{P\K[�u����Gֆߵv�,�;]��W����g��8���{6�<�߅zOOHe�hs�%�&g^�#�;QT���\���K�}˾��Ry2�q�ai�'cs��}�����,>2R���D��i����fL䷆m`���j|{����^�yd59�[ʷ�nbOj�4���Y ��u�IU���ow�<k.]�a���r��:w�e?mt��צu��=z�G�z��#Kn�׮z�_�]cC���ז)cxS����>�������W�����&F�H&ޑ�[��r�:f'���Z[6�h�~�"�	��(�㙛��Q��ܶ�\u5��}Ҭ֊�Ŭh�=�.wM�m��*�3s3�TD֐]����p�{۹Ǎ7��݊j�@�ǳ�����u���j����Ց�r�M]�o���.�O�t;b��.I�����h�p9��{Y7<s_n���:��c֙�
��Z���d�n�Cy݂��lA��qfh����8��Hq��mb���U��e�w�00�	�;�G�IeШ�k�KLW�izA���5��şY����t���`�.�8[���{�tB��b��"�5��@�!�B��]HŷHk�0�'7F2a�}^�Fs�T�KG��)����sa�Y��x
ӝ4��w;�&�:W]l_KP�x]&r��>�NЀ�Kx���Mw��Vp�\ţWʽ���y�u�r�'�-��4��,e�K�}Uy��6x�a1�,޿4ٻ�ûP����Ϊ�:e��|���V�����^�����wx��:�l��������_{R�Hyױ��GY���4r��x!��T���7�ޢ*b�/]���T�&�a�;{�QW��m�9&P�4�����~~�*8K�]��^�%v<2ķ_�G�(l�BC��ŧ2Q�nSfE�S�>2�]�̆����7:�ز�D�Va5�[ֻ�J��GCđ��W�6��V��׌�5��ʻyr�o����������E��L�F�o^��g��)k��S[�T赭�z���h�k*ʞ�O�W�f(s��˨p���S�+�N��NOo��9��n��6>],�C��^'�����;+�����H��0�?����������{�b셟���W��s�C�(���|%�X�y��������Dg�e_��~��-�>��nw�n1v]
��\�@�����
�o��5��M��ٻ�y%�o�]1�]��Y-�@������)�mw��^�\u癴�TC�ʵ�Lv�x�9A eV�G���U�ksת�����G0�ޥ�uղ�TZnʾ׹��.e�Z=�蛦��o]�;���΃�&�1]�u�&`�6��uc� ��C=�աʷ��ϕ�s%'&�v��}��el��幋'p�c�,j�veq�Ӿg�UڔX�ل ��p=��hhS`���p�3��'U�L��`5FQ:GK5�����c����@�N3����c���'f�;�f���̓]S�%��~���;���;�uu�*���Y&*.f�mK�����n�����'-���"fK�ꍐIV8g��f�VDRe�#j;lQ�"��-WՉ�A'j��ws0�F���2�f�V�K �U�s	j��D�
bp�F�CC(aWF�;7�c��xC'e�	�X����Ŏ���#�(q�s%�B�3�qc
�:U�dܑL�%)��r�]�шU�Ò�Q���Jn��DҸ%/�K/��ea���;��;�m����G|�PUw���Qa��n�"������O�L��`�B�*�e1���m�h�h�q1QaR�Xi�QE�ui��iU�m��t��+���]h�+�.��)Z�e-�lX,�V��ji3,�U҃mn�j�m�Lb"�q�+Q����-,(V��JR҄�eUբbVT�U��1,a]Z)�*1b���0u���q���`ܥ`���,�&f8 J�;�~��hV���hx�Eٛ������ou2n�K2�h����lj�ͧD�ϖɯ��U�{$�9��:��b��(���I���WG���:���u��U��:��p��s��{� �ox��q��գMeq�ُݷ.��׻���0�G��/��ՙ]#����jX�W�jȻ��� �5�[��ٷ�Y�j��F�ay����x`gl�>^�o;bI;{�4�?g�z�*�\�o%�\;� �33�6ӆ�Ac
e?¶�;���"��:{�W��k�S���?u.�}��՛L5#M�>���6����@=�#�l�gvgx�������s^.�ޱ)���T��{Y�=L�C-��T儴_c���Ｕ_u*���c�d�Úx�g̝ǻ~��l��W��9c���~\�Vd��+j�Ҏ��޻Fʎg=z�J���8Ϫm�u�6�F^������7���u]�,�뽵Z�s�9y��ӧ�Zy�e�����s�G���V�M<jX��|.f����u���|uOP�j��N h�m�A�$'���$7���׾��:����o$:IX|�іHx�B�=́�	�HbBv�I�o)�{��z�t�I�C�E���;��x����a=a�!��\:��]��z�v�=@ě`L��C���׸@���!�v�"��	���Ϲw�w�;$����|��m���>a��$�d;I�M}H���Hy�y�_~/�������ߦ�� ��I&rŐ+$I�
0��+	�Sl��x�:M$:d:��y��]>Co�s N!YP�Y$�>@40�dR�!�]R�<�X����~�:HBt�m��x}I�� o�$)� �L�I6Ȱ0a>`}�>��c�6h�ߗ�#�L����X(Ѫ>a,���U��p�4o��}����51bt1�W_A�>=�6̋X��}�}V+�}�xd��Ha�y@��N��Aa�̳|�|3Ξ�����<C�l��T:Cl�]Y�q�o�$)�c�i�]k����䓤
��|�T6ɴ �6��>�� a��� ��'z5��|뿹ߐ;a=� �"�
�8�� �I>H2��d���@8�k}�^{�rhs�$=���dά�L�ݒ�i|�i�2`b�i$���;�ݾ�_y$;Bx��v�������^XM�q�	;B�'l���o:�O��m�� q���>ghCI=I�CI<d��c k�u�q�y�ԀVN�H9a<`g(OY|�{�B0:I*�N��κ>���!������L	*}h|�d6ȡ{�2x�O��&�������|������!�O���Lax�2C�$���C��y;�ts�_���\�=��S�_�N���w�`S?0���UR+o�/�{���Cw��7�R��)����cW��K��x�]=����5���~�B� `B`�$4������ٮ�9��g�H|�z04�����8��yHt�z�;a�H,��J�����<���/�睆���� f�HOR�v�,S�!�I�!�HVHi'�����{���l�{���>gl���r�z��M2!�$8�`�CG��������.���䇌�d�'�0���8�waā�C�1}P$�Ć��C3g:�z׽��!Ĭ!RC� ��B$6�󬐝���|�;d3��^����뾼$<0�tL���ȡ2���I;M�2u��F�^��k�{	�|��$����M���d��C����d4�|�X���5�{_��浯���B�C���d���4�}N����:a i�Ԑ��t�1�h:�݉�{�{����!�S,���!��!N�t��MR�� ���/�����b��3��,����);+�c��V_Kb\�%ٵ���ׅdW���/R6���X���h��~�C	����̵7n��/,�}�|g���ïi�������U���3����]�k�n�iѪ�ѓ�nZ�.��2V_5��ZMc��ֻ�k}D������@-�j�Ҽ�:�_�+8����Gx]5G������e��1-�u�t��S��$�]5���cW��\H3�.�Z"��Q�Z��wC�Qrt\�6���嬫c��ڻ��nR3"��;9�U����d��8@ ���0t]�ӛ�2r�=�E��[�;�:�kXi�H��\d�8��ԭ��&�	��s\vm+ϼ�����=���9�ғ�Y4�Џ��9�6w���ϙ�w�}wō��23�iP<�αe�k�F��vu-S�S]��I=�������;Cɝ���w��n�Q��ΙDWh*�U�}N��O〷��\gh���e�����W�b���\�}�N����˞���<wa�5�ڷ�u�3�vs�y�Wg^����v����lB;Գkv�=�;��K.�+p�~��g6z����{{�o*x�XJ2����H�Q�u�d��#�ay[���݈SC�\��c��d�fu��-x՛t���hlx(��1
�U��y�}�V����a`�/r���Й��^�>�Dо=�������}��nqx��^|H��en��!�?�_'��K��.����'�T!�����z�p�=N4x��b܏��*������}���`t���F���V��i��w��ۊ�9fj���}MCI����*�n�]ØU�����X�ħ�q`u.8M�o�hOC�-�����lķW�p��KN�+�3w�w�8�'_�4��Cr�����x�_ۻ��#�cǯ�!2ǟ�XF�=��=z?o��A���׫������T<7;�B	׀
"������,����#�8mV~�ɼ=�n���c~��e����	���cvM����V�F'v���\�y�YY+}��z�~�V@����d��SY�⁙w��Fn�j�9<:7�۸-�\��g'�v�~�T��:q<k��~��ߟ�����G��Q�d*:��=q�;z��
f��\h���Q^,N����w����\|����{���)�
y���J�+n��R�T9t4j�M:�3Z������t��
,m��{S�N�ꢞ��UG�UF�FZt���n�m��*�n�-��Y�?]:4���
m�^3]%���31޸oE9Y��;�i���W�iB�T�έ9�Y=����5})o׃hҾj2RW@	I0�ʙq0��Ҫ�w�M�ʖ>�o
^������8���7����Ұ�[�f�]��o��/�����.f0]�A���dQ���Fd˲G����PL���1��'T���-�e�����E��C�vӥ����tR�*&i,����H�q	k0�
"�H���Bو��pd�c���|Ij�D+1�U(�	Q�V�����zK��+�&Ք����J�KK!ڀ�vULc%�+1.��r�)i5����{����^����|� �ݖ+ � yy."�eږ�(*�	�8.�e�șdEF�(a`0,��Q-]��*Q��u��2U�����?w�\�TE�q�R��8ZT�Z7(QÔ��YQb���m�B�j֊ւ���F%�em,P�QIZV�5��a��m���Ҫ��1�bR�R��D����U�j���i��`Œ�B֕�ZY*�e�.��Lj�*E���E���+�H�E*SVQ����)/��z9,�ң��W�r��`��Eo�=�Y�þ���}��J�/�/e���]w7O�D�_����<?6g��_jS�T�W��z�[�/���]���Sv<#�L!�6�G:�v�Vl��<�إ�3������V�ot\�m7�+1
����l����t���7Ϫu��E\k>Ư�-��v����Y"����[�xབྷ+َ��b���C�_L��<ʞPR�8�������__���]R���d[�����oR��{9/�}�UP�_Xޚ=������K����+z����je������I�юy��![]�](��y����i�	��*3��GM�U�r�ǁ���O��u��������`�	�m�32�wgE��nR��y$�z���zcރ� ���LC��@�~�9L����&�c���ȥ�7�������>5��p�9�����~&��Ϲ�<Hm�g{��5��gygw<ӦGkI�9V+���UUUU������}�?׫��ǅ��߯Q����<9�g��d�6u����c=�ܸ��HG�Sl,��Z!u�ãy��!���9Y�,���&��!V�,-�|���A��
`�Z�eIc�
@VpU�^�kU�*L���i���4o �8��wP�׼�_wMh����h֊�XAb�T6���B�x｛����a���QgH�"X �u����cA�/��!���-��JXF,�4'�����㐁�Gx�ǅg��M
���n��X��;�^g�Y�ľ,����\�����+0�;�ތᏘ��6M����B����f�lNm���}_U�ᢸq5��B�~9�����-�8g���a	B�
4q��A�a{�/-�V�(�#�a�f�2>8E�i�
>���؎EDx��6��$�4lm���Ng؟��<>�t����3~LHC���+��7֩<�ʏ��t�W�!L}xt?��4��=ƂM����y]v���>ѡ��(KW�Ku�u���,�	Caa��wJ����b���u�	�K
!�hi�T�b�TM ���tG�����@)�R�1�3z�v�~�[���K��[u�o���������Xo��k��V���S���[�t�m��Ůl���x�}�}U�_��|%�=Ex���=B��:!"
���d���N���"ϱx�~��79�7��,쐦7��S���̎��s���o*�q���Ӵu��8��9!�-�Ѧ*��8kx�,��K��|�"��ț~��N��g)�.��>��}�y���B��kM��,� �؄�v}C	���~"�}���r���#�a�H�B�o�vV^[i�0��FrG��!$x�*c�~�$�R������Bj�*?
.���B����MJ�h����i�,!K��
�:2Ѻ��y��*@L�u���PN�l�e�ЏG���J<!��g,�.j��}R�\��)�oR�^�;���Ӽ�>������_p��-0|h��lW����@�^Ar���7�#��J��n��Hx44���Q��1�L����i؛�Y�^^��r y�,5D3��,͑G�]
��lu�<04~�R��˦�B�4Dy��cK_&����#��|qѓ�x������j�����1�x\BE�!�^K������� (�E~/��<x�R��{V#��i���4��R��->#�몝ݻ,q�AE�DYC���Q�)_޺���7 �s�4����8�
#Ś5�s�}��Y�Λ&V�ė�y]��p(N	�삥{�)S]�n1s��k״m�uk�m�3��6������������W�̣i�?7���?�
�����m"ql������ɝ<E�a��Ǝ��%��0`�Q�őj�5aylm*�vB> �'�[���϶�Dl_���"�Ȃy���`�s�N���8<8m��*,�U �0���v��^o����CDu�Lp��%K'e������;����a�l���H3F���;���(�� �Y�0��Ka�t�;U��w��3�%�x��/��tز8��Z "�Y3�{G���2�|ɭ>:xP���gLk�-��÷���~C%&��R���o1���_��\hh-έˀ�R��ab�grǮj�\��ͬ���������!%����$��{�0�܋3�� ���]�D8Y����0��'�`�Xfz���5K�#�o!E��<h��qz���/ъ�����q�qx�KX�"�K�C9�Xq
4I�/ț>�2!���-����=������Er�Ӟ@i'؇�q�1d9����Ah���ERH{#�#�}�̣�^���\�aG�q~�=1����߲�l>�E�gԸ�5���"G�6j�ǒoZN4t�]ϸ�����#�a�ˈ���V� �C�r�,!�~����W0Ћ�����h��֒�[!��%V���p��B����^Ə|>����"��Ȇe?��;8l�"ʥ��J�H�U�����:ƾĬ����ںhѵ�ܠ��A"iں�	<�b���_.yW�R������U���Z0},�n��9��m��jZ,g��q^)ʈ�'FAZէֽ�z�S=޶*
�~>]�8����@�wh�0���a7lx��8��׏>KR��}�3�C4E�'�a�i�/����
��^��^�>?#��B��m#R���u����b���	�
Zk�W�0!��Q0�5-�9��q�O!��������7�����zz��������PxT�膌u��m�pҧ\�Cv��m��|> y����5��b��
A��e +�z�;��mp�Z��@=B�$(Ȃ�I�nVLǃF����
�]C��
!G�������(M�+m�+�v��^�f�L/����"@��<h��A� �*[�g-���R���1��&��i�x�5�RQ���;=u�j�i��Z���a~6���DWwu��6}�.+n�7�+#���?K7&z�,��<y�վ�H)k�F��5������4W�
�E���I�3<����6w���v�6`��Q���D���7�)��@n]k�[w�T�6�
3Voz�;�	��;&k�������B�Շ����+tpze�]�/�QM���;1�>��Qr�܅t�+Q��M�-��N���uX�q�U�4�;Ǝ�͹�}r�t:����m�lG�kQ��Y��&�v}]�6ؗӆ��uV�ݥ�'�z~�O7]C�L#\[{��HU[��F|i��.�}zC�uQ�%Z}�a��E�U�Ŋ��[�x��u5�r���x]��CY�7>�Y�R'�D�,"ЀfS/C���{-��w6,��X�Jh�r�Ǩ-�y��wF�X��R��+%����OX���l'z���u�Fu�U�Zʺ���UD`�m�RL�ui;�lX5WwIVB���qUn����Gm�Y�d��Ʋ�D�@T���G*�q٬"}u�UՉt*�ʬ��V�5��Z�����E�G.�5m2�m������J�XN�%����i=,���Ԟ�J��o�0���ǎ��i�~�{d��U���aUeVV��ٳ]���F}ݘ�+
��EQDcim�����m�ŀ�E�(�DE�1,Qb�Jµ�Y��2-kXZ��D���ЕEAAKh�U\i��mEE(�(�X�V���ij�Eb �e���-(���b�¢���&8���9ո/8f9?x;���oǤ�C��bL�' �}W����v�t��hd���Ys}�q��=~v~X�����=h�`���9쎃�!u�z�>����N��9}zO��uѰ�X�`l�:n|�SX+�E�>��`
Ȇ�vf��l���r�^ ��;Yn�z��Rp�Y�N��g�<h�s�s_׎�`j
���7P�ecp�!�Y�uC�8Y�E`_bf�8�Ȅ��Ϩ�/z��w3�J�$��0џ��{�Wv{aj�Ah!�dU�8a�AgG- X/�~���	��I�_R��g�5�g;�Ѷ7w_AW\8ӊ4Π�;/���嗐C�f�MfI�!ݢ�p�Or#Pӊβ臝OD��������n���Kc� ȇ-�P#����C��#�Ƭ�l�|����_x�Hn����w���\F�<��`�{�qt$��ǩ�sݧ��[c�x���0��B�*J<��������=���?&�:~���_�g��-_��Die�E%��w���0��(��w�ӫ�mP���9NJ��ShKC�Q`{/W5���n�6o�MNc���.g�Y$S��9z�Z��B��eWvze!`�踰E���C�c(��U�������G�d�UtC������6as��	�s}��ιJ��4׷��8�O5�:�X���90v��V���*뺻4��0x����QI��uԕ�Tf�����5hRD��Y$>���>��Y���#H2�"x���4��C��}�*-�خ���`Q�)�O���7����� b4h�}��� �Z��k�x�[��(
у���5����t�ܱ�~d�}���XR�!�1�P�>b�5�;(�x%��`��\��ތ1��T�|`򎎞:t�K���7��I>!�e��ыO�F�GŤ�՚�:�ߪ���n�Ot�F��I�{2�Et�R�ɭ�%��WkJv������f#�(�m}�:
��1��&��mC}QRg\������z�����h�!`\sP��W����<^��|~�P�B��D}~�ë�o�H�=H1�� �
^4`<G��Zw��[�!Q�=���H��O��Ey6Jb�d�b�w�8�:^�\=�q/�	��\�#ԅF)�<t��\��)��5Q|�Yv���d9[�mi�y�
6|X"�Y���j�3��"�Y�'���~��¨�CLULWK�3L�oT�1���TG��Ԃ#1Q��3gb}��x���I="��I(r���H!�ʱVw�I�j&�����h�(���}���oE���UU_}.����}��8GZ&(���k���#y��K�!D=TwW��P�)��aG��lf:�K"Ȳ!����ccO�G��ʻ��7 �0�{J�0I���u�-]=l!Wg���V���� /��5ݰ#��% �ߴ;q��my䧯Bzg���מ{��>#��Κ	T\a�l�ύ��J���^`�@3)i&��ݴ�G@����s��Da�$G�j�r�{Xc���UԔ����AOŊ�j�	�>6 �4V�U�W�a���E<1�yy��Y��$�*�Gt��yo2��=D7��ee����6��/:�omxm Oj��OE��r�50�.��˦��6�ω$���9�y>9}k>�����G�SN�:2�={o$�r�V�'���B�ñ2��,�?�*����c���0�D�>#��tM(���4�Y���ha~X{��=c�}v��G�}:�?PhC�����o.��]�*6U��14`�6l�,"Z��p:��p�;Ղja�}��n��)#^z{�p@ ����&���h�a�4x!�+WoӢ}���FG Q�����"fߏM�u���"��^�Dq�C9Y"Dh�����E_�O����&�ځ+�iT�g=\�T'�}�U}����v�����#��٬i��g֕y
8B=���E��� �]:/��N��<j��-0EErq���$*�c�����:��!�!�ȠE���½��l-Os��S(�tG
ဆ���W�<�E�!;�n{��^��F���1^HSB�G��}�fߵ�f��@;�m�⎚3m�I�S��h3�7K�t����S�:-��Ű&Qq�^R��4B�ƊB��r�4�/��B��,>~�c�#C<:�Y�������1<B� �_)�����Oάl�9JW�Mmi��NX��^��a�Ɲ&�����צ�Ý�Oy'����)3�p���8I����8~R�6eԛ��3�<x���H�C�Cy�>b�<+�~��K^[��!��k�(m}�1�B��F��eI�{l�������y��?u��!����ʼ_p��� ._x�AQ:�夳X��lS��u���`�뢈B0)VW��v[υ���1 3���\Ja��^72��i�q�,�-x�4l���.�5օEg��L�lώ�!�#�_����̦�:�Zf�E����a͊<-x`7��^*��6�Qcu����IWQ���S�,ngN{�_c���N\�7�+Y���Y�����}������<F�5X���Jzl��M�����B`��%��6s��B���3�-�44S(Tg�.����t��Ue	�4h�f� ��~}1c����O�2��c��FE�4,���N��+q�t�qB���B����o�T�`�*?/"E ң�X_n�C�G����j�E�6�F�}��Ǽ��?[R�5Y��k2�͖t��7���X �E�F4�sv�Y/|�L*�#C��� �5$��k���ʇ�qk� ��x������0��Z�鳌Wy��en�F�Z0�fҎ��:T��V���#�w�<�w:hέ�+u)��>�u� >���g�~�Eg��LS ��)
�g�v�\<��<(��U~>f ?>��Z
c৆:�3�D"(ג"�.;3�zM�`��v���������\=��$?p�%-�N��~�P#�B����V@��e��:�;��E�
�������̠���wg����ˍu[�+�eꆍ�I#/}�9:��a�c��"ʹ6D�vfs�HDa�S�/W�"��b��\�Xo��cM�g��%y�ɿ����� �fΚB�خ�PLzs��G�W+�����uv��}XCB�k� sWsC�,<j��"�jvR����7�f��UW���ɮY[4ٲbY��P�q,_LԤ{��F��D#W�2s��A��dͶGA�����p�*�)z�\K��'�I�N����Ƕ�ற��2u74�[osA�xw4�} �� 2Y�yޙp>���;��K2*I�A�{x>�eds!9ݎC��Cj�['I޼�����{�|�gI�7�nm�҅��xw7j���e�=�^�h��5>7�gZ�6=�=�p�h���oO�sG;uErcbwq���<4u:u��􄀜��Kּ_���f�OvX����/g˼������0�>`sz��yղ!\Z�LuQ��ZN��ܞ�[���B���C����PŇτ��y͵ԏs�� ۸�&;���(M�,6���\T�].'�S.�K��'D;���ic�f����f\�zb����]Ӧ��>�iū7�t�@ut��;��Hji�=ך��V�8�'����Np#v����',Gl˾Y�6��Ҫ�f�-�ꬕ���;�g��YV��doq����cVܷzU;�Z3oWH�m���N����
�\~*ѭL�cEUTG)R,1TQc�q̬����[J����ikAEQUb*�*��+Q�kj����(�UQ�UX��Z(�PF�0Q""(�J�DA��TX�Z1�$I$�A!]VUws�L�� �WO��Ƹ�oV����k:��� ���z�~NS[���Yݳ�f�äS��a���j�^Pg��P�b��:�ȼ~v�f���P��0랖|y�8���6!g?C�O�8�k���g�������Z�_QE4=����O.^}g5B���|x�N���
��Y���+�_-p�����L�=!�:E�eA���3�gq=��|ɟ��|ED�#Zo9��s�;�N�0�B� �E�ȠY�Ʃ��\�1��O�i�҇*����f+,�|;YM){��|��qkVFy3��YHphYt�ew�y���5kV��E6}�Qs�3�h�6z:}�W������[:����;�=�j���9;���蓛oW�UW��t������S�@[}>�YZ�աek�R�Hdu/�J˜��b��r�k��J��v#�أ"�ھ�
��u�j�¼px��Kʷ�uΞ��h���� �J�c_dnώ��♭�s���C��s�LB�����p��X���-��	}K/��G��?���/�"��{i��X��+�E=��z_�5��[f
=�*�of�7HV����^�8xAP����X{�N��vhZ��dQƈC��h��q��H~W��[�F�?+C�Y��Z'� V��#V��;��f�6�`fx*��4H|"t�02m���ӧ����;�H]Qѻ��Y18�O5|���$��^����o�I�9N��a�dR(Vң^�n���*<�/�g�<;MlWN�Q!� ��\�
����]��j�$>0U!Q�tQŔƁ�H����{��q�q�+|=�o�P؅���#6|]c?dZh���&_��[�{����CN����5�4F��3.�\Z��
<ڃ4T+2��>��e�A
���{1��A���4������TLCQ	ٳH�MZ��D���|���HiYX"���C�������v5�+�嬴j}�W1ܝ�3'v ����kwf�ݷ(rs�/�Lή�v�vm�mt�[�wO��ɿ^w�&��Q3�E"&͑��i�~ǍW����r=ֶ׏��A���ȳ����=�~=ٓ�Z�e���µ]�(���;����H��ǊV�g �8a<b��z�%߻��N��@���1�a�M5<��e���Y\�0{�E�ԣX��1�gڴ�{��iP���&�N���D*��g��	� �)��Ց|(�x�D��3����򳦶���]���.e���E�(�(�:��>6��S:��+0�gH��0���hY�{�jh�sQ���vW�l�IE?F'f?cn��(��@>��f�o�z�� �Z}�y�ụw]��z���?W�1x���f�,�N����K�~��Q���<h���S������B��z�~����:-i�:����A��Cb��}��E��w��?yS�V���G�b�#`v�!7�^�̊����!��4ƾ����"�|g3��%Y�֒|I����ldZB.��ygT�Y8�e���!܆�F� Y�����WWz;��*�qz��l.��qo���\�5L���?X,�d_!y��=7������*�n�א"��@i��l�˅�SOBSCך�:��a$��kb�B����C���V�*q蛖�氆�����,&ǻF��.��CA������ꅃF�x���|ED�#Xnl�7���Ś�8�CAA�������C��u�)�Y��шa���C)t�y�,���
�����F��!{��/�ADP��=�oj��4Q�t��F2��4\��6eO�=����I�> CG«�CX�+?	1���ȯeks|�������/�+#���R�U��>�_,?Q���Z��#`�N�$���/aO�W����U�B�ܐ��Obޯ��8�+=9�1�=HW���@�~�}����}����TVAg����>�jM��]uOV3>a��0b�Б�6�F����c2�%&[�U_,0\���4͐?��������U�*�&��A��A����	���jؤ6G�WՇo���l�G�#	�cǨ�oW__����k�?,@V!��D��»�v�@�ڶ8}(`�!�<>���b��
�I�#�J唅�0��^S'�վ�!���:<�L5M� �½,V�髀�=��H�B��1�Z��g��_!B{y�S՞"�,�Eh�<9}��ա5/۾��F��G�~$�1�ؾ�PU���;�qKt�^+�>�k* ��3��^�֙�Ls6����}79�##n�������mG�����6�����~b͙�Q�0�;T�6Ϣrj����
�4V�z<MkC�9y���HQ���Z�Nج���dᇎ�o6�u��~p��4Ə\���VzZ��v���";�,�!4E��v#�ƚu׼�v�z}�ST���ӛ��������^Q�:X&HMB���BΟ� 6���r���-�p�&���Xp��{�0^1g�fk��
6C�{Wdi&5�h��;��{�!^�U��C K�צ�V�����q�b���[��ͥ��f�P��sy��X3��&wCP�A�<�����7����><�{��|O�,�F�DJ�)�<F�5��a�jԼ�*O����z."��x`C�08~��1	qd<*{fU�K���4B�B{+^|��ݽI!)�ʖ�<h��=�,�E���uvE^{��c�#�kÂ��c��Dp��d��εzF����cH�$S�6EZ����40���6r��Րe/���+ήb��s�w���*a�*�����DY��$��f��B)�~�%(P#�'�4Vi�{��ܜuh�� ��!�3��t��]{�1��GU�h5�0�q��pŗ�u��*��n��W�U�X%�JN.]k�l��v�Bo9�3����$K��|M��W�P���É�F�C||?���yj� 0l�4�9���8�Ct�P/�޿��:~f5�_��רw!�1x|m��<�V�9x�!�dy�(����� h��֗�;*h(xU�T�:���B��$�����9��4t�<��J�� ��n$S���8)h\�e���ܨ����3��{���'��uya��/S=KHhWx{l�t�F��p�����\[Z��s|�p�J�o��_uG���8�.@�ǽ�^F��hV����*���]9u�[�Y�!�ƪdё[�7[���˒�,�J1��6cFȬ˹u0��
�FؘY�������]�����}2
��ׂ�ʦ_ �x�
�Q��y�ͱQY�7_N�%vq�h�H�EA�GW�x���sӊY�=0�56��z�L0y�:^o^�Hn�S'+�o�է��V�ĭ�E��L��T{�,��*�Z��x���JNrN���wFL=h;�7`��8E���w�J�p����H�Zz�tn���ث�_o9΋g/�������N3�R��yշ�����ںh�^��jL�D��lJ��B��t�?;ޓo7�9�u���ҍi�kr�%&��x41K�Q�2S:~�,�I�pm�Y�ؓVk���hMu9�:�4��U�\p��3�����z���nC�'��0ɽG����ǹ��}���,��E4WNYu�-�[	�J�Ր�n�b��j��r]�WU�w(n�S

��M
�L�{��o���6H�3�.�ɹ�s
R�ݷ`\��˻�q:͎lc�mX��7�ܸY���:�N��Z}��yٳ�!��U�/��*�=�o_!Ou���[B�Q�C���5��J���j�*���c��!�-�=���-�y���S�E��j#%�1QD�m�X( ��X����(�UQT`� �X�1m�12�TbcUDEQ�dUQ*Q��*���
���2�EX,ƪ����E2��%�b��.R�1,UPEr�b"�(��bD�bc"�3&O����λ��nk:���M�5�<%kLMv��Qk[?��U�c���2�������WK���;8p����1k�F���^͛㦖ƨ�7��n��s��z��>��{��}"���/-]u��kU����S��GW�;8��z��gR{:����
"�F�k�$�lf6rѾd�Ä���W�ޝ�W������yv�4���2���t3�W�݈��<=�t	ί>ܜ#���`"C�����q�J��ь�/:B����~��܋�]������wH������b����2)W?h�+�J/6$ϭI��b�z{5h�W�l�uv�`g�}��!�IƂ��tx�Μ�.D�@�/|>}z_.��HU��u�}����Ǜ致<���+�Jma��աK&�w�禑kCJ?��f���{e���� ƥ�>��dԡ�goA��o8*W���`�^z�3�����'��_r!������JZ�;���f��
�q*/1l�o-������Aoh1y�L�Z�5���͈��}�~��x��Yw{�8����m|[�W�v�ziZ7�j��ky�{An�9�bh釻�Gzpx�����U����4�c�^r{Sx�����ɯo�;X����gƌ��XG�����f�4;"�3�s ��F�6��X����=y@����|#9b.�(i�R��s|��
Sj�<7]����Ņ�P{���}_��+;��{�~��#���){Aq�3�u�ٔ��W����Sӡ}�=n�+θV$u/��a�3>W*˿t�G��׊��FQG�۷�=
����'�����잰�n��F{�����~Kͬ�W�W9�-J�c=ز�w����:s{;hy'��i�E[� ���,MIO^v�ɕ�o�������Џ������y��O���u"D�}�D�#��@��X����
��*t�细E�������7a�5���yO.��_���x��%|"{��o^7i۩���/��b�� �-E�>w�v͞
�%�+�f�j�xasءG��Ǹ��=f��`S}G�<F���c�xmi��\+�խ1����WV%����+\q�Ӻ�-���W������b�?Bw����mz��|��y9ZHy��w���K���tK���J�Od9�ݽ�͎���Y}�r`�5c�w���c��E�~D���O�o<�}�����r~a��V~�ךs�tbS��(�Xz|�θ|�k�~)Kjfuy�^rƟ\�+ry��U@#�Fy[�[M )z�?r���Q�;��C�6p)Qwy��ڙSRL����M����Ѯ�����qً=�w��Yj`����z��eg��o�^��Akqg;#�5�z7<�_L�RLr]�K<>'����"��~ѐ�.�WtW�Am�kS��4Őn�řk9�gI��l�ܪt��] ��f�&���yO���������F��2m�'�!���ܫ����gBm2�{S�s�u.��Qrw�~y�;�^~����=��S�A�I��&z����ħmo�gxc�q%�x�֮�*�U����0:�t�>��6�@���Լ���hҏy�u�e��v�ힿbl�Ww���`[0�Խ��Vp�A�0%ЉJ��#�G�Uv�_K��v�4Q˗��ѓ�{��,�W��|> �7���}���~f��D-�]�R7ˀCm�o<��zǈa8x�mה�!g$��'��.�>;ƺh�aS��ū��ً�����e*��{xf��C�EHj��J��qshM�0l/;뮾�0{�g����)9]�^.�{W���Z� ڔ��?�]2��qؖf�ʗ����O!�]�l�x�J����Q� m�]�dS�����5.����P�ﻭLw,�|5�7�/��`ڴ�^��U�U�gd�� b_�L*���{�����1��WZ�m�!d],3�:,�|xoz��9��x9����=�Vt���<}J�u/�u�����Im�� Z�;�V;}X^	�g�ϯ��õ�66q�w�r�*8�G]�4�]��b�A^�o�5���_F����^�ܗ�W�оcF�����moLdF#�ю��G�Z��:'8o���dn�>v|�����ی�'�=�D�=\�]mn?�����7�d�9����W�4��)��W�Z��U���^ŵ���h���L�I��j]�W-e�����5��C���N�nA]S�)}[���ܞ��}HQnA���z
�'R��d�m]����R:{�k��&.˜B�c󽇶n���¹*wy�J��=��AeN��R��7&_Nu�_[���C���k<T�v�Ef�:*C���2�Uu1�&ܜW ��H�GoOH!��i����bH���I��-���1n�sw��Y����1��5w�u�f��AJ�;AF��Y�����7I�e�;��ʸ{��V���y*h�eiE���*��a�A�!��w����<m���.ѧ��������]�y����ag��xo�+��75:wY��Y����\����:��Qq�͏s�+WDQ�o;&�[�w��jJ�ۥ��֑��DB�ۦ�uX�7{[N�4�XIV�������86[S���\�-���E�2���ZT��X��ãC*��*o;{�Ȯ����S�5&M�G鍻x�3+*��C��hӨ�Q��f]"���_ʕM�-�UM)ʶ(�̥N�w��H��."!��a��LnK�`��"V&����������ƣ��QIb;��oh/^ �AI��H��e]����7�����F���z2��i�X�,a�U�E��wJ*YT%�v}-L �xܔj�e�ϭAe�M�JYD#M�f���R�̰ڣq^4�M��b�ct��21X��U�7��8TUX�NU�mVT���Ǳ+YRQ��jX�U+�LkUPTC-H�n\[m�����AJ����Qˌ������e�,�̲(��R����"-J5����9d�墨�A�!��*�Q`�V.QJ�
�jIR�����
���U-��m�\J"��V6�6�TU�Յ#"��U#�UL����DV+���Z#YR�{�u��NKhfZR��ø����{���Ӵ�.�у�N���JOr���RY֝��~����Gv%�?��p��d#]/��q�`z�|bi�.^ub,+uZ�'��aֲ�Օ����-v���0%��w"$��Ͳ�y��p�Y,Z�z=�W�|8'u�����>�����a �t3k��a�s0;n�ˎfv�&r��qϝ�s˖$�s�C����>�{������������\n1��̽U�@�j�Z}P��Ǭ�:g�������*O���b�	�]����h���\j��s���@}%�}ծ�W�=�y�]��������No�v17�4CB�E���L�$�˥�8�`���ݼ�h���&�'&I�D�^t=�H�Y2ӊ%���L��I��V+��8�Sd�kCnn�=C���4�Kn����Uf躛�&;��S���6y�*�wK/�z-�)���۔��V�I��y�'_16,���Vu��jԻv$6�K�W޾�~?�}��c�$_��<�b���c�n����W�/(5�Ox6�u^���8��@m�rFC��
�t��W���i���G<ػ:q�� V���\k���F=����-�gO�������ܙ>4��:|]v�mh5
�n�$+z��&*�������A�M���?`١�cK����FQ���'���������T
��Kr�#��ꓭa�C:\�k����Y�M]p�9܏v�r.��z��w&�;�:���F�d$�2Q��&� ���Uh$V����BΠ.C����ᏹ
Kt:����h݋zҫ(��YR�y ��\�8�=�Ճ@��4��n@�;���_���.�k���*f�����^�Jt��eE �y��g�fL�݇�
u�GFe>>T�ݴ�u���Qi+X-�y�Y���wF�]%�_N��0G��ՖISQ���}�Gp|��md��붯��=l�QɐWL=�y���v��:��+�캷��n�T�o�v�S�?{m��&���T�6M2@G�1sP49���;��-��%�/�� ﵇��e.=�n'�2��G8�4�6�XU��Bw!q��>���-^  ��8|�>˦H��^�s6p3{T)�����Kn�J�>��2��Χn��HQw�P��g-�v�ۗ�02�]E��;�u��0��n��ዷ���H_���\��6��䝀��-Zw���ot_�W%�	0*�d�]jV/<��ɪ∺Y�3{�jI�<+ҶLðL�7'��Z��uP՚�n������a�M⬾"׮�Wu��JO'�׃2�H0i4�2і���Ú�P���e�Pܙ�g_l>5&��[Z��x�;���Vݯ�g��q�^�I̤7�����2CьŠ`u������6�[��$Wf�����j�����z���U�0�k��0y5xFT櫱�(���;gPv��~13��=�tz*�[�^��^؂�j|�um����J״�h{.3��.���M֓rқ�*Ӿ?N����ٿ���w�,����-����E�����yU��k�N��s��ų�����Gbe
�&.��\��-5 ��FZ���]�s11��6\��e0xh�k���n�9-nN%ָ�R�ۅb}��?2i�qU��\��l�M���W���v�e���k��0������+�v��L��ao��Q��ǩ��\�:{�М��r_��D�����oWKd��o�������W9��3v��|��~,TL��pAA�vF/Qenk��Q�=�j��m�e�X��it��;�pͭ��~�a��\�:�.�m'�i���eo���V?X}�K~��5����-�Eqz�y{��&u��X��R����0��=ْ�H�\��U	�V(����M�����=�n�"��Q�4u���e6�����������*����y8yˡ��6�⨺�'�U��0ߣ|�K��r��u\R
���v��P�'�7���k�^U����\��ʚ׋݉��D�⳻�r�=D�U0G�>u���◣d���D<��x���{�h��~�c�:x���T�}x���Z��x0PS����2�K�k�v¾�\+l׼��^�>�&��N�|8�\�ذΎCM2/��\[���	�ɨ���5u��B����s�N�7b�^.N�pv�Nχ�cJ;�R=ܻ�Z�m������u帟��Ac7��ob�e��tc���u�Z�u����[yQ�P,����}U�n���u~��V��>�t@�<QD&ø�f
ܺ�lnf*y�&0�"���!�f;}�Y�9ݧ���&������ub�&�j�u]`ٸ���/��K�G@!��v�*�:�㹕!D�~ra%��P���r*�xǵ[�=ͯ���x�E"�ể�iնOneM�fh����ޤԺ&�*Q��S5u�T��W� ��*g��%�� �X�sz��u��F�,�MƛV#{L�ή�Xd�k��57�N�w����[�| %��ϝ�e�fr0J�t��+q��o��yn�9txA���-�1V�,q��.ZÀ�]�Z٧��]-�D��� ��wS*K����r��	wX2��*0�7D�uLJ�H�n��XA��,eB%��e<h"��3�$؊�b]�ve��)���6�.�*��6�6�T�.�Ak%�)mT�^`g�t�PY,'0AC	!`8��.�heCl���T6�n}%^8^�mLk����
Q5�1}PS���q"��� n�@�P.��Ma� �%��Y_2�r����&1eXY�'Ec!�jX�PW�и���rb���J�U����0�����A"�
�~IX��b�Gv�r��YrՊֈ�0@��b�b�E��jEQ���6�*#e�qCX�Em�kpj岂�J��eLq�6�*���Z,Y�)K
�
ȕ,r�*&Rb��*Q	YDJ�Y*�R�UJ[+
+m��V����b��VAJ6ՑD@r㈈VKZ���k*T�P+�X("��2�Q~��O7�������F�kT9��ړ{fE�:��\�q��ڣ,1�vֽ��\�i=��tH]?�`�Ӧ�7�������|<B��K�L�"Tw1�ȗx��ǅ_|Y��[��^P^�D��=���r����K����#�^���B�g���Tq��^����V�7S9��o��І;5��F���Kq�:��0}�}�����0m�Z���I��Y��Z�����V�k4����Mh���wLG�n37����7QT<2��E��*ce:����M�U��:cs�~�vF+�f�;�癿a��8�x9�f���.�4%� qJ�j3Ե��^.�U��H��V��Og��	�G]�D�in��Y�&���q�]��dc�d�|���.�C��A�t��Q:���_����f��x���[Q�#�yAu���~M�jv�x�+rŮ����E��k���As��'O�2�놴��a�U}&���ɻbFՂ󍩪� J������O����y���zƙޱ�z߬�H!���]����u�xa4�f��������[@E�V���֎m�ft�ׯ9#�������vfQ�I������n���q�+&�e)�i�>���t��u+jOF��qJ\�|i�W\��N�`�+{�������ex>;�6�N��w=�z�
֠ӕ&�ò��ʅq]��M��^z��`�r�k�ע�Bc��f�̕o����t��w���t�e_���M�l�ED<���`��y�����
�v^�yX�x}O�a�����gm?u�yB!�Mj�	í�*���R��ߧ����ˎߏ��{�9BP��a)�N��jϏ5F�톘���j)��J�[pׯj碵t�O���&�ǯ�v�uμ'��Z�R�'��� ��v;�s܉p=bva	D2�=WWW��YY��{oّGb��,^�2�^ �;�xT+��{�l[��{�=�MY��٦��jC������fG��F����E@Й%�G�3[�zV���b��㵻�jT���l��5%ۡ�d��=K��{�/[��z3S:�½������nVM4�)�he��Q#qi�4��w���UR��<js�R��l���/Мfkc�
]3\��.�I.�Tw,�2v�Y�)�.��]�c�+K��{c�x�yj�Ό�W�.\ �BztR*����
��˥8jk�k�\�	SH{Ƀ��7�疃~۰��|w�S��
������3�pA��q}yll�x�=[<��=�`�
z(�uJ/��n�d�.��O�g*N�{x���������A���g֝;����[&ǛIZ����-p����{E�5�#R�;�F�7יy\�V��<�cjU�9�E*�ϫs�j�.�9JwH/�nj�A��ըS�*3����!�3�淌�s;gH<ڡ�5�:�m9�%(�ע�r������x�z�Q������=~�󓽓�t�w��.^�;�CQP���ZVq�G���	�3/;��9M]/Yx=^�b�;a�̞5ִ|0���^�:{��O���^����r�����V��w�H!ǯ=�DU̬�EҎ��ݦEs�6��:ˬ���7Y<Kvc���[�qi��PU�M���M׬W=���3�뽇N��oV)K6�Z�|묗���y��p��wU�m��[�M���(w�j7�{��>�v�M!�����\��NiT�A���yۙ,{��=�/u�SP4;$7���Jw�8�{�Ð��T�O=�����',��>���_�0x�}�fֺ�Ds��.�m�Y���ʯVYl{	e����ۘ�{;8粴�ۣH�<�W?l�z�t�C��;*�J���Z��J���eoV�}9�bJ��Ed>�Y���-�~�d�ySn��Z���S�ݦ1����Ŋ���=7��T���E��s�K��D�o��W��m�kɏ��\���ɈgQ�ﶧ��W��w���J��Yf�$�εl*o�ǁ\/[��NM��T��笝���.u/�>6{�k�p����l�y,Wn�e��kz�K��$��Bi��o��̾Kٛ��<����7��=�67�y�w�r�,��F}B�筼�릃�~轾oc�ޔ�Hn�)W�F�y0�`�{縉���7��7��z�S�o+�ް:
dVp����6���N�����f��M�{�R虤�#���Q=ۊqe�g6v�b���7+7�O;�,0��쮧��+�A���@]���F��9�<��b�>�;�ymJ˛Y�Po��Mt��ı��
�Lj��«=��n�j��ťvo ��3t����t�{g^ڤ;����)As,h�q]�@�������m�o�M�"�!���76�s�K�7`M��;��(֕ݽA|�6^����9�a[,�6��Js�����
-x�e	'�yG��^����}�w*2*����kw-񴨝�y�.h	���4�Jv�����TV�teaP���6������&N�kT�ƶ��Ugr
���(K�)|��@���l�U�;�⌖ee̵�
�h�Kl�K���@ɯ�Q9u�p'g5�˻���E���0�P�!�������kV�I$��&�����^gk-[�ơI�[V�kA%D�<ݽ���ò�	!\h���M����r���8� �bwn�d�0��b2��B0�6�F���K�YX�U�>��œ�x�TPO�E��j�H�,���(���9��W��gu�V.H!��8,�5�(�(1C&Te9\���ݛ����E �!EE*QIm"�cl*J�h� V�SUJ�Zԅb&$�2��ۖ���Z��Q�"2E�R�D���Ԃ���*((�`c"�e�Qb�V#"�T@U"��V�-�AdPEVEU��
(��*V@X)mE��Q\O��������<�+˴ofӪ�jm��Ӯ�[	�+�W.�W{F���I:�st�ʁ ��P���?i��i^�Ch�����Ǩ[�}}[�}0��LXگVu��K�*��V��7���Pj�w��[c��_��^�9�.����sgF:��ۜ�ʨ�����ͯ`G��
G���c�wZ��n%�t��Ώ.����\*Vì�� ��Fw��J��ӛ��Ķ��r�B���ql����,b#r�l�)T����eM�q=r�.�c�Sɽ��blwj����s��fmݒd�m�S�j�����',4)��k}`��U�z�ֽ���wbk��i��R+0u��|S;ו ������9��y����o�Bt\��cPr�M�
���ǽ���v�c�4��R[��C'b��e��@G��<���ų=4c7��f��0��7oW�y�a�V��+���1oҧ���)ʴ��K-m3~=�s���z�~ll��Sx���:��q?<�[�X|��q���ޭ��	H�k^lIv�� ��gq]e)��]�7{��������2H��`ja��!��Vxeo�]M�{r'��r{�C�>�z�aՒ��ј�W7��a4�n�����[���˼ls5��M�o��SJ�8�9��Ri��|\���5��}�x`���yu�r?�g�>��|i�����{n+z��w�ݻ�Z��}�%�j����4-3�GOĽ�`b]�¥��^��+O�P>��l�]���;z���#�Yæb�z�c�V�{�{^{|5&�'�/0���YO�d����{]A���v�~5�1�MZZ̩���4\�ޛt�t��E�WIL�����Ry�� r��4�G�t���V5�����T%ߛw������t��Pc�
�o����͊�;�`��^�%�i{ӳN��ïw^G�nq=y��y#\���K�|�%՝�-NԌ��wV��z�w��)�K�	B��
�y+����]zqM]k'�����������0�r��޿��a��s�<��~�#`/�p��{x,ڍ��mo���e^�h20���kCN�'^�dovnv�c|����^�>�����:�g
��Q��� �"{M�q�3�x-[�4ȏ��ۀs���%�a�r�2�mv��x���{o-���<�j����j����t��:�)��pv�Yw1hǶ{�Z�2����xw%lYQ��������1��w+С]ط�\Y\Lܽ���������7�*Ĵ7+{A˩�����Hfχ��)Ƴ �7���(,>۽����5{��1²G�UuیpLv�5��;����^o�����Jۮ�����=�����Y��2X��R{�S���y]�������P�vh��s����G3oj�e���n߰�]�8m�Z )އ'��.�{���-}Q��0����=�.�w�.����9,{�g�k������	��r����pʘ:̒d>��#M�i��gc�1N'tW�u�79���X�v{
X`E�=t��0�Q���؅��]tX<D����5�3��5z���s��v�b]S.�'��y���s���"�i��c��c<|S���l#�X�JUffa��ܴ���������Lڝ	ZZ�W�t}t|��*�X*V�]vB,׻LĲ�ޣ�|Ǫ���4�i��v�PJ�x���.�E�nvN�R�t�Y��7�z|8��[�ߔ�n�z��&�<��u���d�ywjA'Y&����7�.���mh ��de�m�
�'	��]��.g�5�\9M�o\ǖ׮�[{ռ�n�8,���HU�il�F�ۥ����9�:x��*����KO�d˷�ҟ����U���ѽM���#�w�1k�}x5&VD��,8�?�;?���+f�٫�����^c������$�	�j�;A��awWח��\�x!c��U�x�^U��b���)�l�p)����<w ���U�H2Z��ڑ�r���x��'�ݸ-���~��ƅzS״|�d���G+LQ]�����XY��^Gz�p��N[u����OB�޻7�o1�}-�`�c3�����ͽ<z�������{3�%��:����Q���W�u��a��ώL�xp������5��g� �f��f�*fr*��=�9KP�zi���!W��}emʎ�S�Vq��i1|GLI�x�:ǘ��9�}�²j�r2�x��}�˚G��D+7��t��5�����X��D/;��~i�!G�_���c4|��ޣ��ߩ�ބul�HM�7�/���Oo4�`JnkTx4�A$'<�:P��]_'ܨڱ�o�&�#��ǶZ��q���J�L������`����BS�hj���V�L�L�{u�Hk��6��[v>�	��Z���2�[d��񵝷x����Y�u��E�aBpY�9
li4v9ӻ$B�Ͷ!EL��z�U�^Rz5�]hv=oh9���ufȉ�NKʅ�s�M��E��9!�`����3�ҭ��:3׶h1�
ܧ�م��\�unA"�����ї.��R�
o�)]��_v.���{Z�&��F�SJ�Lt�9oK��;}��b`1�Yˈ-�Zza���vvN�-&�f���y:%�2���r7�0g��?���\��i� ��
��IеҶ��t�U�8mN�ou֢�a��
	��+Ye��|v<r�1�x-.�'8i��.���ȭ�)��e�\6�m�x�-9����Y�)\�0d�];��l��`�R�����:��=�U�8����<��:�-:�A!���!S!n�yM�D��	�R=0�Սѷ}o�ͭ]Z�x�Q�C4ݠ�6[��}����}ݢ:uڢ�Yz��(v��m��k�>Cb
(
"zʬ �,*J�RQ�J�D�YX��b�Ȳ�V(
Km�kW-Q�j��+�T�TUP��q��J��-Z�5�ʕ��c��H��R)*
,P�%b�Leb�3,�� ��*J�-̨�Xq1���e��b�e�.X,u��e`�!�[�T�9�^�:;�<��]�ꈜW4%	���޸-�U�����-�\�q[i��_4�W��o���3z��]r��ǌ#:��מ^�{.���?5�Lq�]�g�3F�H���e-O�E��Z�9�_z��i�hik�w��A�V�ùl��gt+�E��SG�갵��ȥ������r����R`�[�k�o�+}/����JE�O��=�,����]=�]K ՛7w193ٷ�����t�R��)D��=�EӸN䷢�����^��.������E�Y��AG����ޚ
��ҫ����]~�9��s�� 	wv����� �=C]L�,�����\~dZ�{h���",��[Ӽ/׾Z�֩Cw�;7(�8���'�ǳ��~Qp�o3̃@ⴧn:$�W�dڃp�;QzD_�Mc��=��gj�}]��&��n��Co׋{���-Kk;�<���f�7�tޖ w�:W��{�5�n�������ǩkl]�[�X{z�`*W3M}�]�73���T�u��/�kkeC�5��z&R�z@��m�a=�3zlL��ƌzX�5#�u<��W�U��0UyRst-r�vl�I���9����7���>�h��{��V��	>�3[�oK�j4pOuN�n}bǌ���|;2|�Th5��LC|����}�mi=9�(z������Ԉz�FsޮΘ����R�w�8܏	�-�ȳ�^&ucJ�������u�o{�K�6�<a����J�4@�u�W-���੻�.�
{.Z˛n�@�k�:������jp��im��"GV���W�}Y,z��
E�+'c�������`�
G�`�&
[���k�'�ghI��n���7k�.rN�:�S�oGs���pwj4���#�}Z�Q
|�`ǥj�"�:�����VA[J���Y��,x4ΰ�h�;������YL+ySVV�>����"苗ٝ� T*��'ït��(mb����g2���6il��xW�Y�t�ﶽX���v�*�)�B@->�}�@���֬�y���}�xs=W�E����E	��N�i��%9ƍL�B�V4+���Ag[yf]�Ųj�����>2�o��6�s�j�Fb�=���e��vYo�8^/\깦���l��OX�S^�}�c�
t�细E�yƲn���s�Zdq5|�e`H�4�OQ�rs��͢Eө^q�����/~�-pE���V2�vbΏ`�q��6yN03g�X<_��a�4l��ս�xv��~�*���M��!���}媱�F��OqW���o���e{M�Rm����̭��qe�8��q	ҏ��
��wSR2�{+���5V+�n�}�KN#WO��.����
�����,�c6�~�\��#l��S�E��yU��V?U���x�' ���=�T=�e��f���L
s�����
��齋���{;�s��W��� �v�#�WzIM�y�"8wzy��G.�
����2_�����f��ʓB��� 5ȳ����r�Ƽc�g_s���X퀩�لj�{wW;�-m�K�r�r>�y��hqW�im������+�c$}W���٦�Hvp�$��@�[��ئ��#k��}.Q<��`|~Y{��M��⩾Ժ=0�{3��p��f�c�{��ؔ����[
Oּ�\=ڻ����[�rj�Y&��S�T��7�&�=�Y�}ͧmڹV����t��E�#����K�~�O�{Y*C��6�����F�|�Üy�=B�������)@�%�ߎ<�K�n�3�P��DV�اb���m;����ȸ���t�}3�e��kyV�w��������4�	�g�p�ޝZ��|���#;��]w^�{�}��� ����+z��^�ԡ���J��Y�!��7�HwnS��m��iG��/+��<�_d�N�y�
��G�{y(�����b�[W��W����������,V�-�����g��hMէi��^���˓��EA~��@=�����W_���HS�eR��/#��+�'��]��%;!,l$q�;_/pw
R��$5���u��6Q\�}�����f����y�ǫdG.�������%-W��ՠ���g\�	��|���4+��)z�9�q��Wy��w�/>97��ˬ��0ߝ�w ;��O]C�!O��eo��IWH{	�<���=0N�Ԗ���p�~��	�_�,��V����w{�t�~�������!S�)Z����%@Ď�%@����T�T^��-��,���e5��?�F�5���H����"����s5Ù�;(%6��=!�0?G,���L�P�%�2jl���y���6F��U~�} ���,_9N�Z�7,3���}mk�֖w�-�Q���*L2īuniv
� ?�c�<pΝ]l{  .�  ?�����I,�&_�)�7H7�_���'�I��0��:xjy�D��@��yK�7b r���^3�[2�&E�q� *��z�Vp,�ZP%.��k�i��N�E����>d���0AE=�  ���eLg-(yN�Q@c��h��t�!��L.��K����g�M�VA���ި�`--�SF�M�3|p4I���ҁ�����բ������G���]����� �J� 5�d�&&��5[�?���5��X��t��M���˧e��=dESE����x}ڧ�z8���a�P[���/���1��Ω}�[�D��������R
X��P�� �|S�	�D�K�Ɨ���ɼ��H"��,�� ��,k�DA�f̍�����Z��.�pX*4��O�`���`������2]S�1����)|�A�� ����;7��ڛ� @b�G>�	�Z��	�~9��#���C��:$�9���L|� &F�Z�e��Bx���y�'�ۙpS����tt��H�#�%"J������@/�B݌^�������ǟ�֙�3Pww▪\Caf�<zP�A5�u˞��>�
ۘ��}�?w�_2�CB��U���T0�nܑ=R�d������Z���9Ȼ����Ad�����@@��6 �'���ݻ����M�`�v���Ջ2[�B�O��s�K&��z�̐����n���)�\7h