BZh91AY&SY�Uh�F_�`q���"� ����bM�          �@���,��*���,��c+(	�%�UIm�l��C6�i��	��@�b�Z6`5a�*�&�k�U[0ֶ�UQ��M�k�4PT�2նJ�Z�6�#Ye�(��$�B�%F�5�!-�RͱYj�mh�cY�
4�km6�e�j4�J�5D ��/eV�ɕ�;����6�W �)͉�� �WUSKEZ��K��P6�֨մ�d�ښѶ�XR�eL�V5�F�b�SC&�e�6j���zx�F�jmV� Ҋ(  :h��ڵJ�v�tehжְ-�l���n�Ӵ�U'X��Jvi+�sj�i�;:�Z�cJ�N���H��i%��VT[jj�Kje[kZ�ʔ� =�}־��iM+y]�҃ӥy���)JJ��׼� �o��hU^�k�����)�5��9���9<�٣����� >����[v��]��
��v՛[M-�ilڦ١�[�ϩR�;۫�>)JU}�j�����[3�^^<���<��=Q�ݺ�ݼ��@z�hՓ�|>� ���x��r���}�w��Pt����«�tݷ����Ckͭ���)2��� �4���J� 绯�B��wn����t /b������/����^��Em�_}易����������x��OZv�>�|�������B�v�}�!�K��M[Mil��J+A�@�})J 7�|4[Y��o����+��o��M2�i����{:��.���yӾ�tޔj�[�x��=4���Q��N�}��y��\ ����i̍Q�MkUm���[�J� <��УU�O{��m��ӡd�Ɲ���=�����jb���R�m���t�#�҇9��҇v.�p��i@#���{oLN�&h@r&�S*U�-�(�U6�2|�R ͯo���� �>���ֆ��g@ýx u��v�{ڽL f�R4l=�th��  ;�:͡�2QY�����P y� ��hm�gB��Øʆ��� ��e� .�u@uӀ 6��:�g���U�\�Vڔe�V-�if4���JP �`� �v�@ ���t ]�8���u��p 4w'p+��w@�� �^[� 4�=à�Cڮ�5�F��V�aD��[a�>�)@ y�� 4���AA�K� ��� P8�  0@P�mi��j��A2`P:�� R���P(	  4    !��2�J   @  �~��*IOSjh� 	�  ��d%*��      �*jT��     �JHeM(@d ��$�f��L��a#�4hi�2=M1?��7�?������}����бKK�l}m��Pԇ��;������kw�_T��_������ *�a�'����{�?���(�
�?Ƥ�I��
�
�``EO� 
/���?W���`~��`~��-�Cl
`[����m�l�i4�Cl0m�lb[�6�C6Ķ%�m�lb[�lHĶ�m�[�6Ķ�[�����m�l��-�[Lb[�6���)��-���-�lK`��6�L-�LK`��6Ķ�m�lm�`[���%�m�l`X���-�lK`��6��$e�m�lKb[ؖĶ%�-�1�%�4���m�lKb[alKc��lb[ؖĶ%�-�le0-�l1m�lKb[ضƘ[�:`�ؖ��%�#`[ؖ���-�lb[ؖ�`F%�-�lK`�ؖ����[`��%�-�l`���-�lKb��6Ķ��b[�6���-�lK`FĶ�m�lKb[ؖ����6��ؖ���m�l�L�&��`Ŷl����%�-��-����l
b[`[��ؖ��%�-��ؖ�����%�-�lK`[�F��%��%�-�l`[ؖ���c�Ķ�-�l`�b[e�-���-�lm�l`[���S`[1-��-�lKclKclb[)��-�����clKcl`��J`��� �`�l@m����*���"S��1A�6�� �[b�lm���Zb�lm�-�Q�(6�ؠ� t�[`#LPm���E�6�F� �[b�l m� � [`#lm���A�6�R� �`�0��1� ��@� ���6Ŧ"��R؈逍�T�6�؈� b�l0E�4�؈�K`�l m������銥�D�"6��
[b�l4�m�1� 6�F� �[blm���	�[`�lU-���Q� 6�Rت[bl 4�m�1D�6�R� �Kb�l@m��� 1��Q� ��F�"�[b�lm�6�1P-����(���"F#lm���V���[`#lAm�lQ`lt�J-0P-�-� -�-�-����(�[b�
6�V؀� [`�lAb!LD-���E�[`�lAm�-��#�� [b+lTm���� �� � ��H�B��[b�lm�lQm���T�$`�lUm�-�A�6�V��؊��m���E�*�ض����`��6Ķ%�-�lKm��K`Ŷ-�`�-�`[ؚb[ؖĶ%�m�M����ؖ���-�lKb[��Ķ%�-�lKb[ؖ���Lm�LK`[�Ķ%�-�ld`[�Ķ�-�lb[�Sb[LK`[ؖ��%�-�l-�`[ؖĶ%�-�lK`[�L`���6Ķ%�m�[�6���-�l`�2�6��%�m�lKb[ؖ���L`�lb[ؖ��m0-�l[`�ضĶ&�lJ`�ؖ���m�lM6���6���-�lK`i��)�lK`��6���m��1-�lb��6Ķ��F%�-�lKb[ؖĶ�0m�lK`����%G����(�g0/�mх�Q�MZE���4���EJǙX�F�t�5A:�)���p2C��/5��Yy���tH2&���Ơ$62[�-�ji�dA�niw1$�dml�7VF�C��a��*�䖱IRK[�c۪��֪'r�<D���oQ����7D��ڦ(L��*n�:�7b��	�ܑ�*xr�nь�ʧSw74WUݬN�qQ�(B7u�J	�j���nR�(ñj���*�e��B��0Dm@��A��F���U��i�Wi�̭9�`��?�e�����	�T�I�-�B'�LTL�$��2(���R�#iV�r��F��̽�ʎe�p����uy�|V�:8$�-��=�t&�1��X�D�-�ت�=n�p�Z��I����2�Fȃ�2��[�j�
�����[��P'EVWL�;��n�U0Fs��Qf�}�����%���M���jm^������mV��ˌ�����S46Bջ���:i��p��6v�q�Qk�( {��{1�+�,5s*���s/iRj�b�>�śv�,��k\t�[M�:O]�+,7���K�Qz���wp,l�r��uz�19��T�5LF�Yx��R���2�D�w&�JUz�l�X��am���]����c��T��Uc5	��p�p��2݇���v��ł�+KsF	Y����6�#Ml�w�T"	F�
K-�M�k�3
1Y	�B�̵wT��"㙛5C�X�%㭼s��E�RlPn��ɔ���%��b��ѧ�����K(mCjM�s�U��+>s]�XU���ِe�Ҍ�G1�x��n�8��7�n$�<Ar�]cp%�kW�qwx1K5�N;SEךԂ}b��b�n�fLfm4i���T�h�ņ�W��mْ�ǚ/H 8��}lӬzm��cJ�כ��y47W�QP��%���̼�<�n�m,���h!{E�eu��A#%ivF/Q��Ti���mk�9��E	tqn���KUx#����d�Ar��.\YyM���g0I��V�,�h�3�Fg@ru1ΦV[��c�TZ)M����KsjV&F�ˋk*���#)���n��&�WL����ŧKyU���	��Oj�W�0���]1��Ô�n�Ja@~R��J`5jGn�i����/ݱ�=V�;�����N��V^�&uZ˸�S:�-�i�i՜P��V
�u}���������փܸ�䘝��;�0nR���
!�[l�Ɇ��Z�������(�5x"�Q��مəj�j��Q�m%OKd$,i�XO�BID��1�{+-_,(�»X�׃q��m7�GQ�3F[a�F�XsLf�g7wl�!�ӵ�����P�kx�m0�1s`͠U,v�50�;�-�Ǒ���x��jڭ!9�U]�`��j�Ef횘33V��ބ�n����y���m�-C��k��I�J�ݩa�Sn�S��̻�{�)���$!�FV-J�����Q��]]��j���1h�N'xAt�n�a��Nݰ�!�)٫BJu1[�2)^�b��d���I�Qn�I�D�Ịx1jK	�,�LD�����ؚ{z��'g�)6����;�mV�Jʱ|�>Ɋgq�K3�i���n
��k\�@tV�ԏV,8+1.��E��ur'l6Յx8��+o:�U���{��[ss`*TxH�h��-�/U�QY5�:Xm
��x�8#� [Z�ݶ����\m��짼C�Н#S0\F��M�͔݃0��YM:�N��^�P����&�(
�B-����׵��ł��q:�3Qr��m��bn*������iZ�p�^;�VvM�Z�a!�SV0�CX�R\�XԙqTͲ�;u�ݵ{r滍��\.�k�L�+3f�Kh�7q�;��#�U���ۣ-��m�ph�6��p��ܠ�h̭��ӫMY���Eee���JX4X�dZ����ُ,�L��F
9�Hre~� OA�7n���G�MӪ����P�v�vشI���ڼ����{�V�Xw��q������w��+ͿVޅO2�U�����T;��3S�M.��`��?=�%Ӳ!�ax����;-h�U��Rܥ�V�ܩ�!z�(�n��[J�j�6Tս�`�J�6��V�����ӫGq(�3�3Q�C���B,�AT&0n5��޼�^���̉2/v�Q�2i;%�j����"GZJ��^[��\�Ujkmc��1ળVV\K�'\
�\spU݊Be�{zY�e��7I�c+To��pZ�ҭ�ѣ/Y���Q�{E9��*��dӃ1**���Ԝ��Z󡸫/t�;�֦+��g�黣��R��91M$��
J�B��p���ʊ+z��YB�56�U?���f-Y[�]B7#ͫd���d��v�s�vȈP��i���}3*2�J�%D���U�W�A�-���r�ө�<nF[I⺓MŊ��&6��+`�MV9��x�K�45]�aK�LS�r��)�X��l�z����7P�I���(�r��̆zn�F��x�	n�q�]c�f4�6��Y���Ƣ�*�{b�Ӧf�a�j7��Y�bv��!\�9k���	��]^j�T��۳�BG#݇uU�+ZAb�UhaTڲ+Wn�1�¼$�����֦�O�Z�cW�#�Udh��r���L�$S��)�lJ��D����Y����	N� ^8�������-w0Ѫ�z�9����5��i�8+���'�a�и�A65��V�e4�]fUe8Λ{Xnf�+D��ݎ�eE��4�)'פ�t���A:�˂�
��Ы�0=����J��9{$�I��b�(CU�H��u���t�����,�>��`8A1l)ꮵ�q�A�#�7+:T��*;r�^a�
Ç4j�b5��*2ҽ���M��rk�<�&�1]����waj�Z7@�2o	rk�pJ+3wc�/݌�=��w]!3b"v%�V�x�cr�f�n��t�j���ktGxC�ԙ�aP{@�p��ԕ����<�k)ì���T��ɩ\�w��{��Wu ܻ�{���*�E6��J�,h ���V���h<�,2��m;L�t����B���gt1��r�m���+��a`��	���V����t�0����MeZ���զf0[�Q��|���Y�v��u'�Swh%i�:M�=uNeݡ�.#	s��K�"5��:2�E�m��)d�ӧsd�x��;�Է�J:��y[�qn�-�M����w��
�m;W�B�����ƴ^�\�(U�2�x�cR��n�{�Y,[�fKΘ��*���j��K]�.�o38-vx�����ԭn��totĮ�`5��${��3s�%ا727JA�����75+�j:JևY�h�.��j�VnV1��
ԙ�Dx�b����Z�F�!q���YT�Q��x��4�Ț[��Y٤Q;��<-�h�D�f��� �i�p�R�(��M�fVIR�4�ݝ��X�V!ޜ��uL�x��˂;k&�4��̶��;�F�9T�y���	�uX���7Xv��.��ط����a�J�"��@3J���xP���k�W�^�,)��̆�Rϔ��F�ۡ`�uP��Y���r�ZߘCV�-9+	�Xiؐ�@��Ɂ,��e�x�Ms���x�ۏ��b���a Uo ��-�Ո��] (i����yG2,�JfCACQ�V�������OZ�d:3�2V�Ǒz\��p�76hS58^��pj)EK�ŕ�c`���Vj{Zͫͺ�O]���c6�#M!�%'5i:��^�v!�f��OXÚ)J�+XFf�� �b�3d�U1ƍ����M͹{(�X`���-ȓ�m�m�x�c��s$؅��-��mn�l
��aVh�el�cTۀ�B�L,�^b�&�3E*2`�pۧ��/q���$c��ǈ��m���m
�x嫘�Um�Ɲ��1hs�;��nY��QN��DM�J�m�ZT`I��"��q���j�^U�BUn�)�al����r�1�[Főȱ}Ņ���mf����9���`�qꂰ�<\������mA3Tv�����(�Í0�����9��ӈ�Ue��n�Rk�2�.�2�ȐcC&M�h�Ҳb�J�|k&�Q�ZI���#�ob:���R�J���U0%h�M�H�ȕ��ewfӁ�X�Y5b���u�[�U�ˊ�FQ�c�U�bގ��N���7�W�Hc�R��i�b�]���jm4����M��׆۴�)�%�hM��۬����P�ƪ
����l��ȱ��k��f+�#:2Z��o�՚L0\������f�ַ�#	%�n�Y��O3Ku�(����S�M������V�sO����卩X��x�7���b���ȡ��R�ϯ*ښ�Lko6��C`9��v�h�u�h�Ѹ�lUAK6m��C[
�BG�n����v��R֭�����c�0�sn�#rm7X]�`�aT���X�[y*3�0����)�5��Ä�oCX�];�s]m�������ٻ�(��\!̬Ct�v4!(���Ú*lLa��%�ʞ��7�N�����-;���a�я,����ԊC�1h:�A�!3a^�6�X,.t�qU����P�{�!�gh��f��E�V�ͧ�CN��U{l��q�i(MHo2-×���sp7�I͒��A�K�̦�;��}&�t���y��{�ނZ-X��v��w�R+Z�ؗ;��6m'sբ:t
����f���Ըi�֭%K0�O؞� ׵�[��b�۸��K��D����oowe��+vV3짭^Y7sɡ�i�K�r���]��2�`�.�e�1ؚ��X�V�W^��VL�Pe�j<��]L��x��w7;�nѧ�b���zF�t�7dI��benl�����.�bx�{yYYyv0�ӊY7y��8�s]�J����dK�'�,�g�b��v85�1O�w�]W���ٺ�k�k1;�	� I�l�ē�)�M�<[uC]��^Yr��Sn�wV���e�h*�E�mE�ϹX�»u��KWn���`{��������^��f<K^^��H^QŮ���м��cÆl�MV��,ìީ$ؼ�L,15����b���b�n�R�Ƥ:�S!���ò�ݡ�V�u���ͪ��Dc�ݚ�;2�Sdc,��j�T��5�t��T��CY��ek� �endݧ��݃mǷn�dN^XՉC�J,�	Xܬ@�͘qo�[�ed.�[Ͷ�\�R����T�xN&��jOUT����X�US$��ю��4f�ڽ�+wy�C��ni�6%E(�nb����,�L�1Cjô�WF����ɻhi�*G�:T��U�K�'e�n�q:[�J'赮�:�pI�Sy���������&��o ���z�4�	r ����c 5��E��*�w��P��*Ϊd6�JP�e�T�ޡ�X������L�d��"��e�P`*a��na5#�v��)�-K)퓵X��ƪ��5歇v�2� �)9
̙Oi|MeޕK7�@��e=B�>� /s�5@LIb;�l��*��݆'Y�!NB�cŃ1Ca��Ir�7fFk��Hd�L�:��-��5��\p�٣b�������If��N�)�˷#t�f�\�����eK3��`�ɖ�<�p��rn�����GU@Ґ�x^�;řZ �ɵzj���TW�$�@���f�F&$��⤂v��`ݢ�}X���%ш���^Z�Vɕe�2��2ʒ�Ҭ+2kT*RX�l��ˎ���Z�#'�M�l�:�4]>�t0��K��r�Wq`���Ȟ��jݵ��0e*ݸ�\�m]�e�ct��ņ&�K��ݐ�����.b�.�����J��z1�����!�;��H���{���T�(Q/}"��2��v���x�=�sE���^˴�"Ujq�$lq�֍�r�uZ��]��\�T��z���5غ��qouf���j�&(Vũl�o���Yn�9I⦈;��ov۔�E`�J&�*�-D���l�`���m�g�\Y�,�V+h�UDW1}�&�T2KmV%�c�{��gRi$^9���e���4�wZM�*�}�i�KCU�cM�Y��00����+�v�X	
E�D3i��/�v^���;]��$Q�6u�9KF���tM�7��V⏒��R�"D��*Bsu��V��xI2�ei��gd��ݱ��h�K#�.�Nۛ*�D/��e8��R�K���6�$�.���0��&*�j��v,�>�Q=Wn���VojkQ5�Xt!|�"�2
Ml�Nꦲ�R���s�4�S����177�YU��m%�����恈�ũZE�JC�
��H�A�V%�賄'�cVD�	dJFIĬ��p�H�(ms���$���/M�Z1c����ǫ1[W(� ���<+Դ�̐pm"��#i	�؏;uWgR�R ��B�b�(�]$�����N�8��7U�^i����P9Qu6��{	E�R��1�1��@M8���_>���Ȟl�V�-ib������:���E����ASȯ���h�7B'��اCE�V`���i+��2��	��I�l�1�Y��/�������N&=�
�-Xwj��qP��g���0��Z1dI�jb�rɕ2��$��Z�OVY�r��
����q��i��-$�V��P�j���L���V��:��S�5Z\��iv%�rȥ�����brU��A�[�L5(<K ��+�2魋�OA(j�\�����P�qèҬT�j�Ў���WSD*��\�+��QZ ��5y�ӰY{7�Y�7.jp įf\q�ŕ��޵�fj��j#�3.u�-^m%�cr�tỷ�s������S�c.�-�������ڑ��e��,��B�P;hm+N��oB;�9,�~E<����V���s���V�����-��|���U��ޡ�n�m�>�hy�S��ߏ�a�ʹ����X�"������~_�~/��)���x_Cgv��x�hIpb�ݡ�����/�b�r��>t6�e�y"��Y������[��&6��s�Ju�
jޛm3���U�B|�[���%�Dv���;:��U��\Br�G�-�������Y�x��|yʱ+�����7��T��:�ƓnA�y�������N��`}�q4o}0�e!�(`������f`z��ͷ�%���u�4�9�m�)ŭff�ͷe��r�X�M�b����:<	r�tΑ�˖Kĩ�Ъ+���7tJxn��;��<F�u�����Y���x/7�ڊU��������]g;���맰���nV����M��
�d��u����c�4A{6��r�R�w��^XW�57�^6/����eva��{�I����ƭ�n��]K��f�ه]����`�zR):�����V�(�R��
���|NkFM���,������tuٝ�{^�[�bM,Ѭ-�״ ��(�of������e�1j�ꅖ��'�ݷ�O�F��t��T��}Y�O��V�e㰏1ѹ1V��L�J֌��w�<L��)o}�CeC�z�P$u���(�fL��l�Π�Ͷ�t�mǃB�ض��<,S6,a=r%����u��D���¾�.vr��+X�	�h����$�[ϝ���|k&��R˴��OwZ�9QEV�;��6z�X]��+�lmK�b�e�3���w��V�Mӵ��̪:ά�;h�3-�Γ�V���Eu�X��*]��2����@��fmI[Z16��Ke�N�	N�K�3u0nX�@O:SX�Ƕx{iKJj�7@+���ɛxv��eE�u�7t�r<�)u���p^I��N=�,�mL����2j|m�I����èpT���p�o�Ϫ:׸K �����*s��'M�vŻ�Vrj{Ź�M��ɻ�Æ}�]{,V��ӱ�0vԅ���1k':���8wv��[�%7o:��X�Y�#�1`����X�S�p�����%	X���d(��C=!ݝ�/'k4��k^�ذ�e���tfI�,r�q�,��ض�����ΜǱ�݁�������Ե�E�*&45f�o��f�`�ip56���U\�����ie��Aj��	��u�ف�cFJ�7��]�.�Qν�)⡒��j����A:F�[���"u/a�Y�"0��uu�i=v,.���n�Ի2��W�Z\edhD0e���7��	�7��K$5���JГ����MD�몤ʭņ,=�r�cz88&�z�ɐL7�P��[�&`�).]o$��!���ڑ��d9����LZ|̮w!��Pv'N�g:��\y]��}���8;�X�D� � ��������W� �����x��;�V���޼���+$Q�[��m-�Ӈ\l��O�����Z-��f�t��7��o6��!�r�
j�<��R�)��h5�@z��ާ����1��ѩӾ���m�=�u�z��(�g:m[�ƦgE"��h[���u�O�t����TȒ���qr��w�17��mb�/�VX��v�Jk�&���m��c���)E�.ӛBI�	O��uڮof�<հ�W�����ţn6�a���q��xe��U},F���,b�;��U��I��̻`���V�s'2�0�.�0�a� r��;�89�ŎZ����Y]K/�RL��dnà����Jg&(v
˭ �cU"5`��l�GS�6��253vV�廉mX��S��Pq	#y��+��ה�T,l��]q�I��@���^�%����!��i4�̽�/$,���F��CZ�_�i�xv��EtW�c�O+,�zH��Ovma�������u��H�I�Ҙp�@k���^�l3Wz��?I���ʳ��C$��s�w�(WK���Ωz�d@�W��M�������;kbN�A�]�b��0��U؂Maj,K���w�o*���)�uV�Rc��2v������QTϓ^���T�VG��e�9G�w�e�R˵%�����������U��L�m8w�D�����K_K�ѡ�B�C3D�C�ղ� 4��o��J��y�so9ś����B����n�a�	 �� �U#��Z����6����ꐝ���}�nd���ؙ�H�X�Q�k_�K���f��.dW��n�F
�p}��G��b�(�HˣSGk��p�v��J�qR峎ӄ���@��*`�vEN�����¸p��I�Xqk �*u[s��[��G���*K@�z4E����KɎ�]���Z��n;31�q�����º�Y3��Y#�O��P�b	����N��Y.���4�M6tj�Z��	�����r}�I�b<�Q��$����fqy`\�+{�7�=�B��S$j
�� p���gR�!�n��U2nZ���)I���u��w}�N��r��8���[/0m��x��uc
���B�*Vn�Gow^�jM�law�ϩ\3�=;L�(�
GX]���r����2�]%ݖ�N��D�=N�Gjʫ�xK�[��2��1WJt�Y�׉d��;��z�$�d�,b��u+7F�X齂�@;�&�L�C3��n��s4/"h#}�^�;�.p���v��0��8)�n���a'�W0(�@/#�Z�=�9��3��������t\�)cb\&�fdw�%�A�K#��m��#&���%�K)�;y���f��W@��Q�yR\~̹Ѧ���<x��PV�3�̽Y�����,���s�-o_�����1���qgZ���dv7P;�i]z�Y)Z2X�)T�_`�m���ҭl=ʋR����G�õ�d���{�^CIQ�$��m�:�GY�2�ҭ�
��L�D����;-ZƓ7W�b�%׊͈[rc�qWgA/�;V�]�2�Ӓre_��]0tk��R�T��X��N�팚��8�]%�]���BzV,$��.�i\VAZ���s3����j�wi��}n���1�,ԋ3v�[,l�:��o^v����wYo䶆\� �������F2��@g�䊒ҁ�GY\
�kj�$��*hk8����\(V�ҕ޾6�� �����s9���ʼǃ��U�N�d�����-�ݹ��a3��H�w"���=38�l��s�S�6�Y���fˁ�Rygnj�!W/���p��n����ܑ�9ʵ�h�[�CԆν��]�X<;�Q�
�����nG��P��b��v
��Xx�P�х��rk�Y�G�-��e]9���G{\�]�*@=�3�CI]S�zS��	W�e�׷Bj�q���v�;~Z#��E�����\S���WQ�v��f#�;����ݢ�C7nR���X�ڣ�qg[\E'��u[��zhM�cg	K��f-�J㛼��]n�]p�Oj�{O���FE��M���g�k�d�-a��Ὂ��p<\A���+�b�����N�����R���I5l�{DHn��ʒ��C�<ջ��+����)pyѠ�w9��#���,�tLYkQf6��/��O*�w��Kc���'J�쨶
�'	ɒ��6�΂i���;p^��F��I� �[)v���Y-I�r�7
���M�f��vl7Y�u�(��/�b�B;[�����3gU�/���#m�UK`�be[��Jlfu�}�S��be�.��'4���"X�Km���{�P����3�}������s��\�Sd�n��`�^ƅ��2s�,J�9�8:�x�9t�b�6���o:�|�e�:͉\0�WW���$�.���n.�����Ց
ؒ|��"'�	�K�lw�^���Fq�)�&��Ci䖥���V����+�=d���rt
8;�w�����pp�d@�ܕ/3;U�˘�7��s6�%�)V���t��^��8��㪘*v�*,��F��R_if�\.��{f�ʖ���h��z��$��)���8�`��,��5xl�
;����73P�"a�X��]x�	�-�s��ֶ:;�z���)I�8Z�،��䣚�����hCS��O�$mQf��V3NTw��L����-i�/��ƴ2�����
o���6��)D�V��*��Wh6˸���񖆓(ec6�XE�Y�|�(U;wJv�˻�I6h�/o��:\��k�&�5�c�Q���)jtN�K�����r����ʶ�CC�쫒u�`{�ki�+b]�-���L΢�S�m�6�v��&eᡥ��7E�R]�h�3�쎆�I��\�Y���+>���d�5弼푲{�=S�0v�^�4ze��"f`�Ntb^�M�jW��2�� ���֥gU��7��X�t���W:���sq+�E�4�K�*�[����C�eB��1��ꕵb�ǒ�敁#ҳҽ���w?W��ɨV�!�L�l�T��jo)���%�l]-�W�Xw����ǻi�����\�+��H�o	R���E��72W!&����5����
U�2�9V� �l�
�lDWR�p�h�MJ�q����2E�:�ve�~�`z��,��=�$L���+d����U�\��*t��X�'$-�dt��M�̿gsJ,a�3�'�KtU9Y:.��\��]6�dZ��Kpa��]�:�;��݂hM��r|�7�b���1���b,������˝շNZ�E�B3y[m�x/l(_>�/A��=�%�`�w�=:!� �d�X%6��jV�C:��\H���h3a��k/ҽ�f��yd�Bݯ+�ܲ�H)�?>���h�4i+��lu
�Xjq`�c��v��m�q���\�y��4A�V�fd�u�s�6�u�pͫ�S��}��_CZ(*0��k��.\��n`B�l����v�V&P��d��կO=�s"�bf�'��@<��ꔷ���ep���0-Mp=Hsxő�-��t�r�E\����UT|�ux ��؞9հ��X�:���M�I���1���Y��P�S7�#T]�TGA��;O	�E�͆�Zd��d�ās������k4+����r�ר���pb�ʢ�X��pnҊ�gt����T��gU2f/�8a7]�/rv8X\���y0W"�nM̡y��vjkX�T�6�V��N�v>��w]�-�z�J�43��_4�V�:!E�ףvgdV=�Tr�޵���j����Z�����\ޚo:��o�ֱ⣾}�T59��UB7x<޺ɏ���Ii�5���qr�0s���&����N�o�72��.�����1�]�cԳ����i�1f����:��69��Hn�	�R����ŮW6���%yǺp�.��j�`8�ۢbK��,���X�)n=��JT�I��au���84W/��%P��%	ʝ|{@V��k,��h2p�+(�:�Ҵ�Q��8i��Z˫Ky˼����f�y ��l׍��P#3�*����44�U�}\���v��2(�;�d�f�]̾L��k�:���t��ΕV0�Z�����Y������G��K�G�㝇MX�vږ10i��Ȝ�������d�;c@��w(gJ��m��4\N2����3(�k�|�y��'�%��ħPz��wiSV��ud�0-\ܬ���Mj��EI�Oc�)��݊fӱ�r�E-t_3{qU�:1=bqۥg8�@d��Fmd=O[��K�Co^���1��fkw><X0WIg�\�#{Zyҫ=0�G���>�h�ٺl.γ\jp�[������O#��n�=F�n���X�-�}s{{��P_ly�z�F6�m����O}��4yv��UMtGE��	)a?n��BF��0�/nm�w�Vn8�������r�ӆ�b��
��n�Z��ךj_	��d9$�v��Z�Z�S��p��.�4���;��)��-�usC�:���l�ƀ��sq�'S���;��������rvC�iĦ\h�,=m�B��A
ri��tS�E������'����w �Z�hm� ���3 ���nSeS�����꽿Q�u?{�(XE���I�Ih^�Su�#C���(�V�{���J�E��MA
��1^#�f�c��ĉAYH�@d{�W�TCאЦNG���TL�1�Z�<^"����s�PzFX����iy�Ȋ5ISO�e�5{ً�;��u�I=�c�n{�ɬF<�~��V�#��	��* dB�\}�r&Hh�WńT^���@l��CL??O����Ev���<,��/P���O]1�=�hy��3�D��" McE�C��x�^�e D�>�%g]XO6���[������
"��e�������@�Lݿ��E
ș���G�FC.H�<���ó^�./1�$���$��(/��a��*W��Ξ5Z�>�ꡌ�>�WT���4@;�W�����J�����>2�b�!o�$���D�4D�y^M��>p�E��|q���0�O�?���(�(|�Yߣ�O�?htT���?w�����~u�W���?�~'���9��w�f�؛�*dZ��Vn�A���|����q���][�f+b�j���Oj�6��S޽4���Xq1u���}�'�/��̘�o�����m�j�]���m�v�"�b2�s���-�v
�d�c��\/��(V�gRn�k3EDf��F�^Ĝ�pst^�;ݢ�t<�f��������s\/�)�j�-��Udr�R�%�/�R�ܻR�Q�S�|L뙙�C��	f�4�L�Kz7ϭ����z�ܫ�r5&g�e}��Y�tW��׀D>��< �E�':^aV�-P��֫&�Y]�V��m�kRGъ���]=�I�{��q�tOqS�v�ZSY�l���֜c{�e!�s��EJʥ5��Ѭ�PQ�;�q�!��d��Q�Y�v�
�{�5�n�s� �=�����\]C������&���:92�Ӂ����,O�`�{����aZ	%ۻ-�mн�,��C�;t�ƀ�/��
U�:���"���!o:36p����1�0��g�4)��3RVv��)T�1���K2��em��Nĝ�wSg-�����.U.��LX~��4��+�(��[v�:�[��z���%m��Ɲ���|q�m�qӎ8�>�㏮�q��q�n8�q�qǎ8�8��q�q�q�8�q�q��������q���q�q�88�8�8��q�}q��qӎ8�q�}q�8�8�<q�8�8�<pq�q�q�q��{��>�=����r�Ў�=[n���S��������%�v㽽E(��V����&_�^M�����>ɔ�2ʘ;gfhA&�P���u0�gb�\޵vʴo=ŗ��z+�-��s0��,�����{��b f�|%�S4&RȆ�f��S:�[��� zj�A����*X�u�l�=2r�Z��k�&A/�Y���:VnI�fr,`�7*-[��K�_3��f;��\�p��6 ��`b�]�b>�Ehwu�+����&�9y{.��2��2�9 )���O��ts2�l;|o�y��A�r��D]�ЩS�o	
��D)X�L�m[V^�\��}yi��|�9[�&��!��!خ([�iV$���|-v���M#o[]�9N3i9��9�n(9\�Ѭ��4{��kx�^��s�n$񼬃��\���k�����S���'��.c�;7��q�f��&ή �5B�;�����&�j�^K��K�'�HV�W�s��6z���5�#tJ�<���n(�:)
�}�μ̏�UT��HnY�J'�yTPl��Z��n�ρ�gC)9���q�K�G���ћ��/V��J���5���Et%K�ݏs|מ�����}���֝8<q��q�n8ӎ8�>8�6�8㏎8㍸�:q�q��q�q�v��8�8�8�q�v������ێ8㏎8㎜q�q��i�q�v��8�8���8㏎8�㏎8�㍸�8��8�n8�>8�8�8��>�O��������YS���X�c`�Rݥ�b�쓙A�3s�}�5E�j�-�=�ݪ�	.c����Gu��-����j�S�YO���ˮ�r\!wL�ܴX�յ&h��D�u��1K[�]��!��]�M6i�L�tD:n����}�k!��Ej�n�:�SOl��1�ۣg���Wwie�(�h�%X�[�u6�D5G�i�Ǉ�*&�aӄo#w�(���w� E]o�9a2��\n}v�Q�9A��G{�E!Uq���r抒=�4)叺3����]p�e��
ʗ)�7p�]n�Z�I��9Q[¥\��fU��1w�|�:�vyL�V�,RV����}c���݅�A_;�{�tV:���@7���VA�:�`{֯j�<�'�-l'S����ˡ[H3`��vJ������;�����@��?\��_kҨ;.���k�W8J��R�b�+�s^ pᩍUS����E��mβ�G��I��!R-:��ޅ/�N.JcD�1�����W1��+&+T*��&+���C�в�:�io[4b:���fMݣ��g�7r	ڤ@}�gU�q�����IN�w���'�H|ΑQR�Е+�ɍS��*��B�LQek��qB-+5���*�M<v��q�qǎ8�8�<q�8�8��q�q�|q�m�q��q�|q�t�8㏮8�6�>�c�o���8�i�q�q�q�q�q�qƜq�q�n8�8��q�q�q�n8ӎ8�8��:pq�m�q��q�q��ud�ذo�����4q;���i��>o�Z	���u�O2]��u'J����Ua�bW�E�M�iɦ�4����h�C�:�I��<X��m;X�O�I3��n�f�k����6�`�(f�G6���j�f�6�)�v�:S�������f�4��Png,(Q��+7��Wb�T�-��on�@�7|��D2��Ɏk-�Ũ1Wj�1��vi� ҏz�R���MI��h_�MR��]�9�[Ux��M�ƞ���[5>��[}h���W3Ҷ�$�}| ���Y�wOR��%����h:�.��� 5��/{:�h@�;�>�0"��=��R��1*�q�
�d1�����tH�;h��A7*��@8���a������Md䨓�(P)��}+��I���&t..��Y��ձCIi�wU���
˂�K[xGe+�'[M��Xb������>�fU�Q�*��g1ü���k�f8�Wԗ�-ȓ˝C���;d���,���,����oK��`{�7>����9V�mîK�\c��}�:u+Pk����bֽ�B���@�ku�F�In�
�pK/p���d�1�"n	c:�=������{���U�)�k����3nd�:�%�ok���,GL[{j�\p��Bٱ������j�5H��tNRG����x�><v��8���c�8�8��q�q�pq�q�v�8�8��8�n8�8��8ێ8�8�n�nݻv�8ノ8�8�i�q�}q�8�8ێ8㏎8�q�qǎ8�8�8��8�8���8�>�㎜q�m�W��/˾kA~zݐ���������]`TE���!YGx�9(Ёf�!,C�����wZ�����k޽��wL�ڣ q�lU�e�kɣ�IYܧ�yR��b�V�[���������oew.G�}�,�:�֧:k�l�V���ռ�&˕C��;�ʂԵB:�3.��F[�x�Է��;OEW�n�XcP�Ŗ`܌�\t4%5)õ��S-@C!U�}�t:R�Ժ �@��'J�-�t3�@4����S0r���ՂN�8���gk��`\��DZ� ��I7\�ra�G����pwu��/<��!��ؓ�ǽ�w�2��&q���Q�T�U6��$o�駬V%'PahH�huK'o4���4M�	��*M8ׇ�אYd� �m����d0���l��0��ɟ��;7�=��<W�z�M4�<��@n�5�ynf��y�aV
�Y��B��,]�O����|*�IP��>ʧ�EY�.\�7���(��Zҳ#-����|RJ'���O	�Y�͙7Ȉ�#y���SP��eSC�zn�GK��&G�b.�,���Tޔ0@�o)؎��c�b��V�`����!���p�����^�Uk�n�����ڢ��z)k+��W9:���|��X7B�?[7�#��Cv
}�u�3lkY��k#��F�,aU�3Y� �nrrT{�8�W-%ԏ�7�sgt;�MtԶ,���9X"i����P�T�:����<7��`m駏���9q��鹄�Xd{2�N<�S��/��u�
j�(_|�j�'_K$�zm�ٹwB�L�}�[N��F�7�P/6c9���3�t4���B�5�]B7ϼ5c�DјEwd�H�z��<Y��+U�����?5���zd�+�h���KYk
����Y�S��æ�ge9hh��`�H�|��݁��wV�rSJ6�J󕣷���b�y�����١�C�)x{ri�r f�@nC��޾v"Q��T�E���"�R�J���o
�n��<��9�3��]���:��хn-ˑ��np�7	���{�d��9\�����}�n���	�����8L��|Z�ޡ-��lC����G�(�䔤E|S�{`uл�Z$�LQ9%��O����ibʧ!g�L�R���&Գ���ʀᘞG8����ht'ybm�7�������_!6����}K��@�V=���'"_n[]r+J�5P~gW)�𭥕/���z���n���w=����,c]�Gs��y'ݡ�vYY���ǅ��{{w������w*�?sߑ`�]��A�X���y�\����
?�jU��A�l8�bQ�9����6�׻S+@w{v��_�!�35Xe������V�!�8q���wBI���t��fU.c�����p��L��'�-泹j$�XK4�u[7]��Ŧ7ot�V��1��U��\D�y{���݅���u����MS�U+z��Xn]>C{�fⶹE}V��ab#;�҉ʢpw�q�R�K��8kd7��:g��/���(�D�U�MQ�#�=:���/z��ˏ��Γ�Q�m5����t�0ɘ�5�T�h�d�4�����4y�c2IǮ1)X�J���u��X�YH��ןgB:ja�(v�8��۴��G9�m>���yu=i��u���jp�E�!)�ԩ��"�Nl<��D��b͝}�˭��y�mř\�u��d��-Ynt����+�����ܮϺNʚ��Z�v��qA��b����f�va����⒋&�}��a�B��!kcꂻ:�ٲ#5R���JqRT�4Z�ỊM�������+;u�����b�{�kVmCl#�/�h��e�9�uc���*U�̙&���s�M�T�c]�R��&;^�!Wm����oCwI"S�y�		nC�09V�)��")Y�$s�(����S��0e�`�Յ�#w���Y)�S
����1�����$֧F�awxq]���%��߾�.������miC���5Sec�d֚g-`�]f�ִ�!܄�[U.%��o;�[��M�����V�;�NsΚk��$�QxR׶�8�oC�$#��������vI����u^U&��,�|�477�<cЬ�tzj�k�ƕZ��`2��/�S2R����LA\G")��-Į�Jޢ���8_BGv���%�m�w*jV����_��H�ǚ��v�(ʣ4��O[��vT5+�Sx���`�/+z�Zr�V��2�+]�k���Sx/K:�-�G��Df^��{-�.�^A�-7În9��L�P��"pn7*��ς{\f�	sN۽�eɯ2�]��`g�YD6��O�]2��p�R�C)����NM��,�d�yq(ui�p��9�9-n���f�KԞ!e��A̭ӷad��u%�M�*��j.�R^�8V��x#���V�6���x^�<��M:�h6�2&�WT�pv��:�.at���9uh����7
-7�Ni��(�>ڧ�C��/�MNy�Z�KVd8�ݷ��U#���5u��O<oF�-Z4��^�.��SKY�(^cכ�^'V���3CK�U�;f�QSP�*=��˭���`�U��7��ݑ�71���{{x���.�Ww�bY�ݼ��R�7��1�
���P�T_���]a����6�u6in��2A��(��k-��*̭ao`5:�9�)�c��}Kn�DT���; Ws��D�M7��Ū�VS91�h��=%`;�hgoE�v�a?���76e�ۃ_]��6%LC�Os	f�p}�QWI�j��BGP���;�׃/���j�5	�wL���R{̥�u��i�N"��6��-�\�u.#��աw�l:��}���mT��ڲ5��L�+2��������Pm$��\�=����F��nhi��!	��o�롼�?{���	��-)��<i"ݢ+�q��Q�Jt��;k���&>���na��}�KKSKL�|7�sGF�����=I�D_t<9�2��p��\�Ō+Ui��e&�p+*j������6أ��c[U�Tc�W���=fʃ]���dZ�WNMV��c�I�w�,+놠ܛ�'}g��[�+(S[��6oh{[�U"��ݑB2�IԤ�=�nn�-Nv��� �;�
�ӆLI�N���bC�v�@��bS�ϣ�U˶�u�&Q�yO�k�]�$���=�,��j���ID�ໃ���0O��k��1��Ú���!���d�ob�\up�]؉�B���o:�*�T�Osc��o.�=W�X�.e��4>���8�R�'1��Om��4�{���ۍ��M��
�ٸ�9:�s�mpX:�J�y�m�r���r�}����p����R�}-��Kϋ1�t{\�8����e�׹#��ћ#C��a����(��!��>���o��x%i+�)*��i�.��Q���x:Ml�������(�UT"�t�} Q�����n΄wR{�Ey�Ζs�չ�%[�=M������XK1�¾7cWt˜�.�ǻv�'6�	[{ר��5��T#G$_�`��Ð��N���1J�<�٤�}`��KX�Rŧ{tRxY̎Bf
�t`;�]S&�S�f�Κ��]��\�2����m�J]�xv�AM�)�x�]�;�!J��n
��v��*�.���.��T۽���Ω <����E�3o��Ά�XsP��`D.��ר�����O��J7��ɇM��X�WS��OE��I�*!��B9:�ps�}�|n�`��B:��^�-�&< ����#��z�[,U�,v�N��8�S=}146�$�vR���-Э�P��
�Qn��)%/d��#|�s��u�9�ev�^�SI�{��.�bEIm�Pݚ0�<qr�1��v�,�o�H������$ކ�c��M�Q�h�E>�M^lss.~w$������ډ{u��h�7CcH^�sY�FW����G� U�$�����/�c�ߡ���U\��_�z�j�fH�`H���B��T-��^�O�A@��%2i��be��I4�BY�׊.1
P�IM���1U�Q��.��8�~����d��Q#%��(��"D��q���O�x�'�NT1�p)!	ǭ�iy�wA��4b4}
1����������o�.�+�y��V�o$=�L)�J�E#�]w�a����M33�wˡ}ȺPC�����7Tv+J�>V������f񑎬��!�� ��p�PȻ	�f�:xw]�[Զ��,�C9i�5s�ʆ�У�T��˵}f��D��ke�{�b����)'*�n剙���\�&���H{J�b�Xc���]��Ȁ	�i���?Zp["����V�l�)71��jCO��יݬ�K��DjN
N�W�N�:Ny�7(�t����`�}m1�dMU�Om}a퍼_:z�%�[f��vd'\š�X�5��G���qb�G�3�O��z	�,���މ��V�Y8r�@vZUbΕ�ݚ���W}Y�TXtݥt/�-<R��6]��ɎU�ZAU�����s)9���Ze��le�@�r�:+ݜH�{OHwy���jU���aވTW7�e�R֌�l����~��;��LlsgLF�؅�swof������,ɽ��E�	)�	5�m��7RT���6�&!�rf.��Ǽi����b�Q��)��):�ㇾ��h,u<7&е*��yGw�t���Nt]e��$�a�������9�����䑲
	����.�)Qd6Ce�Ei�C�&j	�c.[
EI�"D��nH���iSA�P���~� Ji��	A�	,�"�$E&���DRHh��1(�P��H��dH��|�i��%(\1��q�)�8ѐe��IMF�!���b�@Sp�a�@L.ѐ�E���Az��а�a�0�C07�m*"�	D&&�,ƛ`�	m#I�ڂMHA�Q�l�#�JFHh��2�rE"."b�$K	�ԁ�R�% ۞D�q)��|(��IETU29��b�(��-H� NP\�"��#Ox��nݻv���o�c��Q�g�N��ɹ0�aUE����Ү8aD��i�6�8�۷nݻv��<�.�}�Ӗ�bWN��.9��r#�(�����v�IEp��/Z���o������۷nݻq��v�T�e�Aru����(T��5�i�;���|��&N�&�SD@�$�t1t�TMݭ,%J�QD
t���׮ݻv�۷o��;�>!��8+XȊ�$P#���a*��@����s��!ʎ)����M I��-�&;�����H�c�7�s[nq8WL��`	'bEP\�r�)�R�����@�i�Qd�ȸ?wp
����l<XrO]w�R�����wnةW|d�V`Pι�V'
�LT��K;��ql#h!�N�s��+QA*��z�/B�]�6�+���H��S�O�Z)���S�Q�+�$f�rN�D����䖎A8�TQN���e ��>���	K��}��>����'��dZkEe�D�s���5:�I�W �K�RIZ,�VQI%E$$QUL�L#��"�PDrò �.ʥ@�8�ȡ �aC�hNAeEAW"͔QT\���
�ӱ�}��$�Q��a򪆐i�|�)F�Fb.(đ�$#c�k�`�#0�s7��y��q)��Z���'�
�n�7[���w\���ܻ�����HP!d��D�Q� �
��	�Kw'u<�C��;ˑㄗ��H���FH��X=�)²�d�o�O^4���-�a����C���������m"���f�'l�e����UJ��8��[���dޭ&���4�>�7�0t<����Qq��)��*�"��%�˙>���$��&���Hjހk������iX�Გ$@��y���51�C��2zL78�wp��]Ȍ[���{�X�rŉ���{�{({ݵ�uN^֛�N^0T�X��z�}�'�㾽9[�1�s�*߈�sE���<�ʰ𮮾~�\�q����,�UmO�>$޹n��~��E
sw�,�ǚ��=��0����K+g��s���~S��إFO���K�wϫ����[=6��!� �۴&}9>�%��ZX����Dg��G=�w��+ry������x{�'!��5������E4��p���Wh�hU��R�����r��[�Di�Uy �T��n<s������˭�&�?iʦ3-�H?D7���ѩ�ԧ��f�茇I2��/�x%ڙU>�{,͖����cD�g!M�X��Z��qL]�!6G����_5~]G+�痿��9����7]6ĿVQ�P.o���
��?lԛ�:b�r�W���]L��?g���{�b��`�#�>��i�.zg�MF�
F�T���t7]r�z��ͫY7o���Ʌ�o��z>;�O���t�!L�����C"x��;�~ף�r��Ƙx��������ox�/����]q�^�i�\����U��}�N|f�s���EO�7�޿
���!��Q�5%������}�����ջk:�x/ޗ�E�Al�z�w��n�켏ó/�s�*��|�H������{z|�n�>�:�i�r?z*�y����|�'ѱޘ�z'��{l������{/t���]d�P������NQ'M��`f{�,`�Q��o���էܟ���W!����&��(M���,�Vݛ:*���b��j�@����"B�z*��yzL]���otv�꺏5Uʾl�D���sS;)���ï�4xc�gvN���8D��}O�®�s�~��9�{�t�xk�������x���+��;����4��~�X����uo�y��O+oű�Z�G�{Ǎ��r�ї�m�@5���W|�o�s��P��Nɵ���'�މ��[:�z�K��;��%���{�~�����Rz*X�v�}�Ͻ���$���9�L��f%ﯦ{�s�k�ѩJ�@�`W�{K�9��{_|)���b�W������>�����3^+���q[YȲ�¾ɳ�b��ȅ%���B����t����T�-sg�>zj�ʡ2�2�㎎�eu˙��RK٫ې�K��]/-��<+��	ɕ�}�S���c�����)0o�fՎ�����OW�0��eͯe���E�͒�u��l�|9-@�P���ц�ve����;�_l
��>��wH�����t��k���&,K��Sk3쩺�J�ѧ��Av�7�!�n�����{<�,6MS��v_o/�Y�74_��m���3ے�+%wK�a�}��띥[�4�{rJ��Bfk��;�>�LRg'_}O�"T��)�=S�zf���V����7��b|�����Șv{���75<�N�^=�.q���~��zϭ�r�
.�'��o�Me
jglվv�J*�C�����3-Le�/�N�i��U��W ������RN���kד��v坠S>��|������ޓ~�r�̞���~� �{f{k��`$�ߛ?��_N���{lN>	���[��|a�jooX����f�g�y�>4�}^�����M�ףe�y ������ƃ14f�����7jZ3��рI'�����y~C2����8��Vf�r���9�m��N^�͏I6w�'u�
��PS�MGYv�H�ߗ�C3W{1��\�p���5�O;z�R�i�y��戃xl�8f=]m���^��zDA���=��v���%oM����[[k䮵�v�c��J��P���-BsDuѡxa�#�Ehm�u]I��;�v�n���f{=޳3ب�D�.�š8U��w����IR:-݆�
h(�N�Ӫۇ�W�ܚ�x䭽=�K�k�&�4�J�׳��B��s�C�U�C�dCǣ��-ͭ���!�|�{��'p�B����DP G�i��}{˷�����@H1AOŗ�?���A{;�/JOshf��:iڋ<٪�V�s�g��$�_�d`��8���}�A��(ΰ�Uy^�t�IV��n����A��0u��P����r��y�Ԟ5��w(���E����[��d+�}i""�bv�SX�@�c{��Z��0x���<@�dt�Y�VxVv��i��.��X��{bB7Q�KG��C�Q"\!�j���f���� T�xq�g�	���y|����Ϣ}��<h�)\�������t*���y��W/9�������$��-UI�ħ�>�l���z��yլ�a��^�?o_غ�{�R�#�u����e,���1�6ڼ��J�~��������k:���S��|�~�L��ȨZ�L+�;�_N���}Sڏ�S�nUw��|<�:�,��]�#(�NU��~9��V�{¨[S�!�2����6x�ѳ-]/��s>��L��A#c{`p;/�o�]�9���[h �L��i��t��؂apy҄�#�3�\���wl��-�X�#��Oz"R�M�U;����<�ɱVA9��Sr=t礃������T�=U�r��M�z8~��g�@�n����7Ě�y���z�G�n@�a����gmzߖ���{\c�5~B���oc�MH���m6�=�hpܦ����s�l��A�uO˽���^f��2���w˽~k�us��-�nw��}���'��=�hp�ڮx��k��}3ҎT��ux�P�x�>����C��x���u�ڵ��n.�<t/p��f�[{�DD}�W˾�y�8������!�v�쉗@�[��,���Ƃ�ӏ���X�w�;뭱�foe��T�o]gbPV_T��V/��o}W!��栘��:��-ch�m�faW���lO}� �Uo��?M�������=�����k�O�,�y-�䟡s-p{�Y@����U��r�9{�<D��,a*{r�g�n���eKήsͿ}�t3��>���g���*+\*����
�|sU��m�@��t�
@=u�V�)�X�f<x�U�U�m��)p�+��.��V򑵓m��:Ŕ⊽)�q�v�<)���jv����j��iV��Ж�z�'n�gW�׽�N=l�Zc��f^�in|j3koŁ�_|�T����U�g�a��?AY�	\p���n׺�M)yo��yf��o�z*���w���{�{jr�|�dk��#�<`�g^	�����95����8����n�����ل�8Ge����"냋=��{�Y�k���*�^�m�$��oOw�����իx��~g=O>��u�[�_�2�=ۆ�V
iOEY�����xzl# I@��,j������M地XC&r�t�73z\�k�3��#k	8��"+5��G��g���fOM���N�͘���l�q�����[�h����T�ߓ��|�	p�{����xmy��^�>u����}���#�^�qq�>���w2�7:|;�I�=�ڶ�|V����6Ȳ�Ok�:�V�9��μ�h�H��'a�i�ґY,:<h�T��qpr��J���=뵾F�싥z���{������I��Y��1Ǚ�-}+*;k^U5��͝���[���܍,�/�̤��ٔ�U2�JKdG��WOV�k�y����~Z�t�/�3H�4&�L�'�EIq����ƅm���eu�!8~sk���Of�fk슟�.�5�MUuht_��g��x�(:���7�P$Ys�n��y7�5��;��O�]tZ�{4��2�cF����i�15S[������䆜dw�Kw��ԗ_>�o�T�{Z47�VѝbQ��X|��57n)�g��I����r�W��\��܄��«y����]o�iS��{3���Hgo0n��Ȭ��3Vw�k�s��'�n�z!��p��b�����8��{��w��|D	�����s{N�ʰ&<��j������L��ӹ����C.�Ӈ��E��K��-�&�A� kj�J�M���otI-��3{k�?�MAh�i���O��O�k/���Y�7�uJ��+˾y\��):D6f��2���BX�.��
,nqa� ��,����m�I��u�Z�/'n��	{��G���8)P�Xy���K��\��5ޣ���Ӥ��p���V]���W^WW@sZ��tz�����t����D+��"�62�N�	��{֯�����nO^U��	y����N���E�T�1����I�[�T�o�R�aOKy�Xz�ǽ­����`�{L|m����������{�w[!?/8~؇��������);�ņx�������^JzL�ׅR�=��w~��v��L���S7��i�\�{&�ʘ������ݻ��s�W���K�w��"=�;��4P ��ϩͧ�5hUܞ����D��\6��fU�'W�b>���UK������zd���h�3+^�>�C�Hd�~�� �#:��Q�%��S����)x�e�ٌ�'�i�ۻ�g�� �1�k��p5���b]�j���.�=;�:��`B�~e@$��>� m�ѭ����0?9��vs���Z��^��%���h��a�����ۻ����3�BX��V�D�*�^Hݩʶ��MX)e��_
v70T\燐1�Q���Iq��m'�1��d;w�c�D�_*U�؇�6���%Au�^g�׫σ�ϲ=����h�YW@,�1�ʋ~�s42�[��Bp��wS�R��d!�����&���Iѿ��j��z������j<#���u�j�_��hYxvL�1���hm�t���������%C`f��ԖR��G}ͷ֔�-;������}�>����ާ-��Xηe����$���+��J�p����o�&~���b�*{�uS���j�?of�9�۬��D9}�y�o�8�W��׾�L�g�T߭����W�5=�{L�e&��2�`�W<��{�=��*Rͷ�<:�gT���Q;[��ހ{v��ַ~����/AC2�(��G�륵�K��8��ـ�=�~�Kc��|3U��M�3��w��d�M.�S�����h
k��ʞ��h!	��//�q���ܡ��@2�#�����N�(��uCigIa��7�=�����>-P�Y���}��	G:ON� =D>��}��Cν�<�_���A�{5g0�gX��6�ѹ�C �5�zӬ��*�����Õ,^���o-��{ASFR$ͻy��K�]�b�R�yXS|�1�m
�1��Y'h[�1QY��\}=Iuym
_9���|�_h�ע5ZJ�E<��6�]��1%[ۻJ!0�=�7o������:X���>�>N3gu����G{Vw�f�O��nP�ͷS-�-Qtƕ�T�p�W3��u^.\�#j;M,�z�2e'�p�[�|��i�`0�W4F�>��;w|e+3z�7��ω�#y���o�:�sU4�i��] (���v';4�ϕ���^�w�:�Ӿ|�fB�J�u9�Er��|�t�_?Oy��uG�se���=�Ѫ.�]D�\�d��+̘�B䒷k3 �����s�����\QǱ�;��N�~yέ���h���:�o�wK���rnB�)f8,Wn��UUӆ��5�s��X��	�/k���'G���N�ҧ)�����|I�)*�ƳwE�p�qvҼ�^�ƃ7�P��8�C��8��5�fqg����܋g9�J����K:�2�H3r�7�e�dV(�]�m���g`��'ne�2�;�86�6�6GC�I��f�I�fݼ���X�ܵ�����5;�	�����=+%�V(A�opɸÏcL�sRUGl�ꫲ�Y�a�rv!���kp'����U{�R��~��H�6�1�~�V�aAT�>�3���H���������>}��^'�:�:������"��n�ʦ�sf3ݷ����tk.�&�A�z����zw�ݕ�(���#&�d����ζ����P:`�l�i$0����W�A���2N�r���u]����6��ա�A�a���Ɖ�������=�Kչ��欘�JQ�zыNrj�xP�Iە��STm�n�f��h]���#N�1�S�XºR�U���A�IG�lt󏸌p4��3���s���I�#\p��2�[��ܹ��k��v�ߵcj��vc�_MG��*�V1���}��X\{w_�%�%f;��tA�%��RT�ڑ����&��MX����]5';1(��ej�[�Zs%�7�9/8&�;�s)�V��^��G����	�X����	�L�����D�˭�V�8EY��4�}��Ko��W�/�E,�ou�4�"f�(!���:��OZ��'-S�6d*�y\�9R����h�l���=K:�t5�f�%],�td�6�R�4'Z���#l����ꎌj�ܗȐ��\֔%�eun��h�vԸg:��O"�F�d����ən)K �:m��(��H����P�aJ�%jH/i��^-��,\bᖿ{h�P~��Q؇NӈqT�'N\���U�G.EvH¨�#%@�i�]�q۷n�<x��ףޝ��5�\���$���K�G9y	J\щ�FR��T�TR���q۷nݻz���|7�"v'
#�E�d�# � Y>&�
��؝%*)t��;v�۷nݸ����;e�p��!;C	�����t�0�):LzIª;(H�� T*�=i�ׯ\z�۷nݻv����)ɨԑ�!I$! ȡ ���.W����H�w'2���U29F�߀��Rj�j$k.G)K*�T!b$]xRr��2�F�����J�a�wU%T.�kN'MS+8R��\��Ԝ��H�!$�N$Sۉ9�8�8�ǜ��N'.�$�f(�?��E&Os�p������z�E�+��T*L�8S()�Q�]�O�H�C�șBQ	QUȥ
UH��aE�L�[4((�"�)$��b��y�����u���ܔٗ�}K�����yu�']"E�Fq9���U8�xbyխdܧP�v�@�1�c罿N��}}4��1��|6[`[cP}oG7�P��6� ����0Q�H��ae��SԹz��m�ʥ�|=��	�<a�d��]1ٰϳ(�[�f�	�'g2Qg��߱�L�V��ַ����b�j��=��8��6ϵ5�g�\_B;�@i�k���lo�?]�Y�v�
�z8d�1����wNd���i�¶���N���&���Af�?����Y�,�t�~�c9��3;�-��w�vJ�^;Z�FgmUU[ŕ	8��ܽE�~���m�OΏ��ʛ�[K�+�X��a�&'n�]0�N,Λ���Gd�M�+� 0����0	�r�4ɒ�
�X���_���Et����FM�c�E�g��[^���ᬶ�\�����鎽,�.��g+ؕf硳�NC�H���^h�tF7 ���QbI���U9pp��}����
��w8��*��IN$�s˨^זU���79��ND�1�����鰽�.!��ϊ����O�3��� K�,e�P�V��b�b)8��k;�-鎪�~x�X�� �{�����CH��@~rg� q��8~79�~k ����+������z��m���w;,-?�26�g�*��ZB�������i:���B�,ʭ���\���ӛ�L�M2 ��I�1���ta��H�蓴���R�]s�-�[����f��օN�E�򸳶�ˣ��f����:j)_y0�� f�:W�]� 5�S1�1�����p@�	�~��i�+c`�?�B/�~�d��#��Ix{���d?G��J�;f9�v����f�7� O_v*��* F6� '�u��@0%眲��tod*]k"���M�~��{�K�vh,J�U��WӬ���ϯ��~����~$�ԡ#W����q��g?ym�*�E{���}`���*1���>�8�=>�(�ǚ:����r�]����)�u�K���}\G����ϼ�;Kј�L����VG�U����V���c�ez��h�rIt+4��gGwaD�l�e�ԛ�>�%����P4��S�}��&��5�Q��xh��5��a�1�V�d+)�=���v걫ϰ3�Q-��~N~w�'�F��^S�oE<�.�6�/b�^!h����� k7?S�}n��bb[��:<ڢD8� W�3��0)�z:�!�ngO�:��=�r6�C�  =��(Ŵ�dޖ,�-���bޯ.��~QP�:a���o�n3���9�29��ԙ��$۹ ��j���^���6�� /�x�zX���턷�/��9�}x���k�P��~,�^yxl61Z˧^SVrN�	�o��L�5/�06��!z�r�n���>��۳h�3�ȇ��� ���u�
��a�^E�=�ÝI���\K)�LJQXWgf�j��Ƨw	����lغ�`S�7J���3V��b�n�>����w������Z�Y�� ���g]V�1�~�������V�5����$�V��|�����*���J�G�qѵkk�&:�����#�M[�[�bb6t�J�m��Í�L"ϰ����vl�~�05�P��cP�\�����u~P���I�n4�2�?�V1	��ʞ��n|ۮ�o+½�n�9K���c�|^� j��C ��4��[\����'��5J���W��v�7����2okr*�^�0�x]zL��^��t��<2��w�
p?�* � ��O]�=3m�C����t��xI5%��y����j�mJ��hi�ٸp+���`hZc�;RC��Yx��� k��~�/C6��|/�.(q��na`�%�/ sO-�K�����ܹޔ,���j©�����uxO��LB	����*=��dV��08a�[:r��ŷ��,'���|Pf)UUWD��� f �>ϓɀ��#<>
~@*���JY>G0��F�_����q/\�vʧ�A
N�$�;^�0q,��d��~��4�~�@u�Da���?��|����2�X5\_M�,�K� ��mi@Z�	�������	���:�J|_Ų]��	��[#��r��ڰ�]j�A}kev1�-��̙�^��'c!2�ݾ��\(5�����-�
;@�)-���f�;{m0��yϿ�u=�1�]~�42(n���%E�;F��w�5��t٠��r
�;+q�N��]r��=�>���U��EoW���e:β��Q���m(kՉ <S3
`0^����<-�R�MA�K;�)�|uB _���BhJ��KC���Ӯܣ\�[�^�����X띋��� �lS���� LIh0%6�$�3�����fv����!�ӽ�|]۫W����6	����pb�C�-�;B����sH�=7��8�C	^)�l��Q�!�r�<��5����x��Qz��ɑ�D9�)�ɀ���&�9"��Q!�_�)W�P��7q!eG��b"�w������b\ST�@*�y�ů��V�����ū ��u�-���{�O���=@s{�z��)c{&!�[�sy4�{��z`-���]~��4] ��Zv�ɞ�KU��u�-���@x��dF1�&���8�6Sl0���K���p��C@5"�D�c9�ץ��&����C���7mG��Ϟ����&��]�{�P�K �m������\[L�p-�jPM�Ǻ�k1�wk��=���Ǚ���kd���z�T�� qz���
�m���p9�8v/]�g��zV����x	��*bɵ��a��vV)O7�����5��*�{
#�m��Ǻ����U���[ǡ�j���O�����v

N=9��ح
��3n��B춰�v��|A,��v��f�b��B��2ҋ���e��c�q�w��&$[��eg�&>t�;�8��٢Ȏ\�L.ϥ�q����e1��)��$}�` ��ރ�%�)@xq�l��������C��6� o_�����-4�y��o:{��מ��!R���Gg�}��_�V?�G�+�$~�4�@�O��K�{��8���#L�8�WF�{�Wu5Y0���}�
����|��]���z3��ޞYgjs��&���^��߀���O5��ǠbI������ޚ{F���9�6�\s+���`���	�o��ިO��V�I�H�?>!�R��Q�ʂ�e��x]K�4mDG�()�e�:W�$]W3�g���6?w��߹)���&佁/A��7"!�����&��V���y�<bl���GM4��[����ybx���߆�4��;_��T{�uļV�A<����M�qx-ZKJ��3���6'�⚳�fA�.n��x��� ���>��)ӑ��/M�����i�n�����>���d���Xh�'�ʋߐ-���a��!�W��[Ս��;^+t�ܹ+��������%4�`uM��� X�{/Bي�	����a����2�h�9d6�a ����>� ��Y2oY[4ڕτ�)��p�́=JϿx��p���Y��?T�����2��i�ퟭ�m�"6����־��*��-�<ces�\����k��>)g+�|ŋG^C�j�����rr���)]wL:Yς�p9N�M	��kBmPޘ�=(m�+��|k�K@�}����o)�8����� /A֍�h˶˱�\�v(�C(��*\G�@LW@�ׂ޶���>�� ���Ȧ))�{��i�=1�������c�ڻ��K��0�s�S ��'�����q@�+�	T��)�M�Vǫ��٠:��K]��^���*�$�OM�W��L�T�`k�?~ڬ"G&��N�׷ �}���n9����R|ܫ��N�j���i�g=�PO�L���0c�L?��D���Bu��C �Zd���|L��"���m��硻v��5��.[���+ݸ���ӛ�ۗ��ԭ�>M����y�s�&����ŷ�2�'ov�Y�q���Ùݘ�7 LQ��.�~�� @�� ����������,Wv���������.����EP�<�W��ք�v���sQv��pp��ݠ9��;�b�Tp~ݞ��8d��t�'=5����</vq�ǀ�	n�� |�&��1M�
-����Ǝ[V�@z[�^�f#��z��X\W�?7����^�Y8�P��?-�q:�U
HS�6�f�Yk�+H6߉_��]y 3�S"j����&X.���>0Ŷz	�Vb{-o�L�y:�P��V_d�q�܊����"T�X%���|�!��,ޗ�8��5�gW�����{)�W������#L B���\|:��3Eޖ��{���������8�q_M�Y�*����3-��h�v�'�l�<�q���)�Pj�!���	�ƒAi�������U�V!EA���Hz=�{j�3����3@������j� 7z�b�{z���*�ju�:z�,5��[c�~�N�Dq�g�W�	�8�܆�v��񛕩�f� ��z;�¹�6�xʗ�f�W^>&i�W@�j����>���N�lw!����{N�6WZ��g�s��U���_�
FeB��S�1p��vn�za��Dx7�7��e�o��Z��;8��v<%
�d�Ǚ�P&~_���@������q�𬰺��5-�xsĴ���h�.OJ���?�=6���nxi��E��F�&��n���<�K2F�k������&=�ﲾ��D3�ܦD��G����f�]���������:�������˗s͂=RX�j�^����v�ظ�EˡC��i���s�^`@�S�P�d3��<�Oϸ��F���s{x��r�\L�tc�,�����j�mɛɊ�J%e�?��p7��޷S$��̟?�3;:\1����GoQgj������ӗ��9����(B��b���v�n1��c3���tOV{�ۡ�c�m�\�B�~.'��������,��U�A���r'���b��ׄ�t5t�E�_m���[\�,ze�`Sq��;x��m�i�v��}����{9_�O�������r�m���^�L������p�\FȈ��&���.{[[��^,+��(|3�f�u��w��3��_�3D�@�P�i�Zi�B�h���U�]�׽�w���ς�0��?LAq"!�]]Ƕ����\��OC�w8�Ia�ӡ�6�Y+9B�E� ��D��s"�A'忓{�~Z"�M��NO7�P��=F;}&��o8r�� ������QS�1�S�_��WM�PE��~������o�lI�����_c���ꯞ�����>Ř5���@��&׌l/ C���
��/B]�����Sk�����0Ϸ����|����]�U�>ɛ�w�}��K�ty��L���|�:n[O�=�rr:�/{Ū�E�'8�#�p� [�|f�,t��a(�5�L�:z륫˿N�J�O��{���c�^�~)ě�gǞ�W���N�[�B���^(�����ؖǹ�/|kY��'�ʼl�5�7�;�/i��&��Ĵkzl����qmT��a)ӯ��'��L��0�%q��o����� 7P3��Pu���t�(�$¾�߭�)��2�g��6�Q�1l�N��=}Vw� <y�]aɤ�`��١,��f�����͜��>����;�[[i{��&Y�*�~���е�!��d5�����ƾ�N��^�ֆ��ʔ�-
�@�/.ngv�l\�o�<r�X�
��HJ��d�oN�#�Ɗ1��y3�8��R��&���iW���FS��l7VandWnb��Fn�ȭ��_U}���[l��ְk[�aCSM�X
��!*"�7Cys7%z�=�0;�x�ߙ^{�S��M�ߕN0)�^C�.)�q��_NE�w{0?FF�J�{�> s
jb9�5n@Eֿ!��OL0���o��m�N6��m��S�mw���W��-��쾙�p�Ź�[>.�?6��L��2���1���z��b~l���x���3O���j]�o8vW�+�t;��ަ
[���M\�zA�����V�'�(�lB����Ib���w74�6p��A�C�3ǡ{��jȀCۡ�1�Qv.��(1�6�5.���!���lW��8��p�c��xx٨i���fd�k��HW8��C��>��`_	r�V��yh�G���h�M�QM�f3�A�Uŝ�@x�F|��3�����W>�o�i�,z���/Z2 cG�zC�>L�(y�v����?}�{��O����^�����A<��G�oC����;����U^���?���^��y��3EXre�!!��^?�1��J�,)]���Ey�ϑ/!��\+YL�7j.=�S�ߝ� �����B�-^����͛�^��dkz�P�P�ӫ�ן$�P껶}��k���} �U0s/$�hg�w��y;�h|9�E���:�Qł��W_nV��,������ �[����=�|��Ϛ�N��^e��T�R��{�SvT��O����/&¹�s��Iݙ�<(?hE$X�@�M4�P@#M%DdAddd�Uqp��j�@{�޸l�{|hw��;�d�W�3�}=>.+7����8�$oٜ���S^4C�R��U�����Xj]r�5��P)߮�ˉ;��&���0;~N!�B�EI����3�[��9��Q�y�v���wC��H�8���O��Q���]��RW�P�;�*���>4mN\��k�Ʌ��u��q�ځ f�z��:j9ɕ��M�\��î����w�~��掼�3��a������#̡��U�HA���rǞ��.�`K=�J��������y������J�Ϸ�;��Ź�&�9�f��� �-�4
�8¼����I��
���-���n�j��;Q�@z���M0�̸�t7c�!��bQ�.��n9��Pf��g��9tk��\+�g��5��ݏ> z�̾b=CZM���7�����8�{���!G;�7�.?��>+��R"yq����oV�^����c��]�Cf ��VX��ԑ�0Ҷ6��T_��`�i_, �g�]_�z���7��l)ל��ɨ���%��k����wq�� �A�����:݄Q�}�O#�X[�_�C�تuÕWR��V���#\���(w6�j�".����"v,�Q��tT��V�Ɓ�v����L�U4�.��f��e
Xl+�T]3�A��JD7(d��b���Y�vؼ��[W��֘�j@a���2��]�q���X�'��o[.��cLS���]&�<D�%�[5�O+�@g��<��.�륓��d̢��&���i�S*q^3��������žGt�B!��2��j�$���}��[�~�g�2�`̫	��6j]�1q�>z�c�89d�w�U��)3���8b]{�&�|FSª�q�'_e����z�J�PǓe�v�R�^g[D˧3�f��Z�l���D%c�L�]@��uGb���.�~����sonK���ٖ�.\�=�3�	X�i�^U���}n�ԒU]'�y���2��抺��-�{6n��j��q�]˓�E�&���
�4��K�#v��2��l��T�bH@�b:-k��%z�����:K�D}ܳ��ޥ+��ERYuj,U~��2���[Q���oa.�9��*�u�CR�K�,6Х�'��M-���t6�Xy�R�r�F�9���,rL^J�kwK/Xe:�pr;�0GK;�N܎�+�gK[�"���#�����T��Ғ��yc�W�6�]*m�ͬ�YE&���iX��a���-���B��Z��4��Cz��ӈV�b�a&������t�V�}߾i[�u묿h�9°c)�O��Ζ�;yJ �V#�3�mow=l��J7:�ŠJ�%o���1����-�v���P율E�$��P���,�ݣ;e#n�L����[�V��f��L��9�7����K�{�Ҧ�HkH�c]5lM$6���� �mV]�a���h�M��-w
��:���fVԱ-�&r�� �W�}�A�Ns���}��3��c����/dP���X̙�R��v��0�z�Ve^�#FYq/���z)0��s�׍hϽ����廨�.���j��wD�&!�<��S[����B���:��Wj�Ks�hhdi�tV9ޚ㵊�V�>��z���n$�
��;	ѵ���f�ܣ+k#ϲ�|��ǅ[]��ر@�7lLd践mgU�ZU��h�V\%�eKצ���0�_.)�n+Nua�SDP\z\,�tOag��+�ډ�h�@�nk.L�"�, 8לM�1+��@q�ǀ��ʺ���uN��ݲ��<����s�fG��^'M����;ǜ�/���zOh��+2�[������;�F�$��}���Xŭ�.�uۭ�1vp�ǜ�hO8�vM�O������TZ�wA��y Z�(:�ˑ٩D鸯s.�ˁ2�*����O���Ku+�D�ԃmv�B0�*���&�t�-��-*81*�1H�*Yj��˧*�=�A�!$d�%e/+0D����M���>�a �}}�/0,#��z����&�5姅I!�j�@��o��|x�Ǐ;v�۷�G��U!UD Huiܛ��m���()���F,�ZBGɩ i�q�ׯ<x��o^��b��Pd*�D�$�Q�,�I���wCJ�8U1�Ҭt�o�8��Ǐ<x���́	2G�bsіp)�¿T"(���P����Ȃ�(*�C���$ ʍTi�]�㷯<x����o�����D_iFT$®QC�N��$���:���p���k$��<�U�E�l�W����	���)�Dj�f�����EȘUSy��x�R�_�}\��!��4�L��}!��Q���u��9C)�	ˎ�p�$�B]�=��������J)̙�*)��.P\��p.$QԶ��Y�ЋP�E]ɉ_x�Bt���=j��t8�v$���1"��.KYa���m4���������eT �!h$d ��4��scN#�a�Z��ι��Nu�N͝|�g�
ru�n�h��\ۏ8�lM��+�(8^�@�eF��u��\��{�zE/:Zx�B��	�~q�<��^r�d��PA�����>o!�<��.|B���bߍ�!�4�4�@�M4�P@v0e�.(`��`����A���UԹ\6��w��5�]g��,��K�2�_8�Ǣ���X��c׿/AU��qWӋ��ggٗƩ��`��O��SEܳ�Z͊co3j����d`43����q��zO>�2$n�N2��j8�9懃:�{��k���߲������g��ֈ8N$T���wi�}"c���t�T5�����&���[��n X�;�c��ss�����|Dl�׸�"w�W��$����>��z���3[g���G7u�9���nQC\��E�R�iE��`Xi�U%��|�r�o�^3�}BW�Ha�ß#�f�la�:���0_����������q��>�Z-�BW^(�;���j�����jd��}�YL�O���>�s�zN-���j]���ϭA��������-�<?F�~�s�=�����]��ڝY��3 w�L�1�N�OL �f�\�X��~>���0��zC8�Q�8���Du���,�~|�ύ��xX�O��3�AAO"n�r����c��9�Ъ��u�R���*ӣ'�a
K&�ă7>_5��R�����B��!9x��C�^B��=��g��X�^�v��>4 �E�L�k�e.�m`;6���K��8��I�`0�{��|ǁ�~���ĵ��WP	���Pա2��yE}��]��X��T�h��3�?qn�K����Y�
�bI�����K���+�7��� H`u�1�h�5�c5D�� d9�/�|��=��܎����{��kǥ��+ܮr^���SH{�h9N5t�j2A�ǹ���C���
���צn��'����Ѽ
�t�,ݍ�3y1C�];5�	t����c�n��r
��=�!�޸*�<�~�£�Kq}���M�;U��o���sC><��*A<)��wy�1,�)s�m�mHM��^����q{�X㊭��d�8bo�T(��+s6l�Q+7�ga�.�C�f�2�e����n��lF�V���6.����	|g�6i�z���[��-s]�/m��ƽ�������Z��o�I���`S�)�����FƊJ�`��p�����k*���c�fm�LB����ώ"���i����Vv���;��=�ʼ��10Ѫ��{����c�K�)��rk�����q�0ǜ3i}�;k�0_����w�R�r���kt�h\�ᴃ2�l$(�&����~ ��X52�~�߲d�ɻ���ƥ��Yf��<�a��컿��q薑o^*1�v.�X���4�f��ｇ� 1�����w�\4S�V�3���J�d�f6�܍�ܾ���c�Aw��(E[�0/;�_�Yط�1A�N=���ds�~�t����[sn��FU@�s�rӶ��)>�`˖[3@N�X�W�|�r�_N�jr�w,7���3����->v���&.��S��AO�x=~�EJi���i��  �
�"2
  w5�w��y�i�b%��F�"���~b��y����Ap%�� -���i�CXƉȹ����i�Ky��:���2a�<6[?53�������Y6�V����C��+[��^�.�C���ݻ��3ۘ���$��R�2�|Yf��\/�_/�tu���5y4)�q.���#W3yd1ygd�i��,#g��6	�Ʃ\���1�l�)i{M��Q��c�ٳ����3Ƿ�L��]@��Zڽ�]T۠�����M��T��@�ȳ1C_�w�lB�|��*)�/���9�����]��j���D�0��33]&�e_��H�E6���tKe��L=�ű�5U�M���yG��-�.h�!�B��g��R��⣘S�׎駭�����:��=���a�k����+߁?-;�ꢏ�����z�Q�T��s�{�&^���p���g���jc}P�cʺ�j_�;�!���z6w=A��{�| E}�4��Q�e���zҒ��0)������`hl�-%���=	�w���T�Ϥ�^��o�t�[m#���hej�w(�zo�*����-DJ���'
�3_<`�n!kڥ��)��K�9-=',u��7�մ�Q���v�����Eu��sF��#r��A��I�(�b�d�{�sˆ�g&ku�<�}@zc���$0�[ִ�1�Z  �� ��<O;���\�[}	M5T����sv1ˋ��/���R'�y��������7U�}����K��G��LS�Ǣ�li��r{�~�B�l��F?���.3�8���~�HN���S��%��KH��dÕ�}��V�Ѯ)��#g��=�A�/խk�����5Y��j���&"�|�z���E}�H�{��K�:@��ݞ��Ɩ���C���6�?�G�����ͭ[�τ�˘�Z�r`r���Trʜ�/�`���{K�##6��A���(CL�`�y�o�����]���%.��~�°;���C�;�U�5Z�Q�2w��ԸJ2'e*��5H�3����W�4�y���BR��׸ĵ�����#Zf"�����H��Y���[6��UW4�/G)�B�T��{�J�ld���`+%O��������Z����`��A�'2-̽B;8��)mB��M��s��s�5��:A,�o��q�dQu~["�))�w��QiM�Jؙ�W�^��X�����d�����-��E��o����N0���>k�R��Jq6��z�w!�\D0�|�ˊ�EȬ��hO����|/j��c:f�M�^�L��Kl��{Wn*mm��S�%��܂B�4�Іύ�>L%F�����J���[�xޛ2��cpWY�2���.����S�.m
��6c/�X*�\���igf7���t��FԂ_��ש����?X�1����v3�6��`ִbCdT��R�PZ� ��xI�8�s"��݃s�����\�N�ChIx��?�-�����k�}Xj'#�+�j}!�2~���d3@�J���meoS��|~�
�Y�;f�V��dcp
���n�7s��a9qI�\�.CsH��K&ي[��K�GN���2D�S�� /K��>��	�W�#]�C�i|���?t��;��/Vqmc��D��}ZE(�{��7d�XW�zF�să�A���\�O-�~���YZ0xt^�t(�zdUj��c�J���_�����|H?~8l���_\6�~y�s5���XMon�������Q�Ǥ���>��I?�g��M4k�C�%l���W���;�2�CV<�Z�Zٰ6�S�"��c#�o�Ķi�;���cGs4l�^�Zf��e:#H���?@�(�%~�=G�X��!�:��~w����v�e	���͋4�5��`�O��y�n�.y�ĪKS��t���C�<����
�5�S�(�P��A��o�~^��0�����v�L��r��d�j}�h�i�$�,5�wU��ʿ
c�/��{����U�xE�Nv�]n�V��ш󷷲;8R�L�!4ދ�y��`W1ّ��Ǭuv�HI�}Ӟ�9�m��2L?ms��u\���LΘ��0>���RX�iv	[���0N'�&W8P�r���Ӄ(w�[`-k N�:�6�e2����1;c. �"H2 ��3�˟>{�O�o^e{�z��w�.���a�tz�b��r�����p����w�����Og��Lx�m�T.�Fm��2�OL!tSH܉�g�>x�k�3Vhy����YO#{�~��g������~szD\�er� ��s�T�)���X<&���~9y��c���ir���ݣ�uɫ�x��dcg~��>�f�r|�_<?�d��4�5��%�\�gYzz ��#�g�l^=y�8��c�N�з�qM>�$O�hƐɖ�f��ݫ��{��/�y��E�G�3w9�׈E���_����5A��f��XT?p-�仦��v��|��S!��Æ�Y���CԠ��&C���!6�T��Q͉?�ۅ�Q���Ћ�f�;��;���:���t)�5[�m�o)�ё;�:\��6��_�2Y ā�"�`t;��Cɞ
ss�鿨�?h�pD4�y麍���O����hUS��;.��x�I����w+c���1��Ge0�&5�3gs���� ��*��ʢ�叏�x�����k���^���a5+�^�r$򉫧�n�N��;�WK��G������W.5��.�j��t6��W���=틅�u�=����X�~�R��Ӄ8ja�a��%�{(�4+b�՚������s_�b��J��������J�1۵$���!�U�cM(%4РT�4��@!QD$A$b0FAVA@E�Y[�~r��󵛔7r�}�0�f��T��L[,����և�'��0����]9|ݒ�ʢ:���FGE��-/Z��0��-U��yy�^�@��L1�؝ٵ�o27��x�ܳ\�u]:�b儋m��3�3 SX���♹��楝�^��ie�W�s��W/bl�3ғ���OC�魙������Xǻ�F�b�4���,�m�+�mF�X'�Y��㖬�w�W_�V'�V�m��j?T��k���e<�Q<�?��F�F��a�_�ۖ�Pn�2'��y]#��p���6c��&|8˧M�T�����A�8&���=��,jAl�d��c߂�y1\�<��N�`	Y�{�F��?��O�h^o䲳5�+�A1g�j �2y�b�����_�A'�ƩC>?#�����w�_ȿv�I�wF<�s7�NRV�P9�v�t��+z{��]�M�P��(�������u��>�sr���|��-�P����-�h���j*z1�XG��]&{Um�M��0ǰ�xa1�]�m�E%�q�z�3v���&������5��*��վU�t��ˆ_V�%+ֆ��>��T�řү]�D pA�����+&��U��387������*��c�z����G�f=�j������;��ח\e�}"���������ֶ18ε��ílQ@�	I$#xx_.�6�|�P�L��5�ޚS�Dڸ	�_t��n*P�5��ӗ�I�1��ʪsӂ&�
k�~Y'҆��w5���y����wO�bs�,�6���<���j��!��2�m���:D���+��;��86/�*:s�2��1��P���I~;���7�.͘�b�j�6��B�29��.�yG7-���@��@f������d��J��,�=ɠ��vwظd�kO�Y�u�l�z�'|pg�]7�4��`׽Zk��Y@�1��������q�3�k��r؞�軻�:�/��)��U�7�3 ���A����:��`ɝӻG�%���Rg=c��#e�-�6ts�ib�t�z;'ɦ�F�u����z�ϱ^�7'�'��w�fY�p�!\�%���wٕ��#L�_2Z-��oU��1��ď�l����ʇ(����������"bە��������#jENK��mku����C�����ð�\�$95.�G"s��
j
͘�=����l�ʟ&�L�����9ʥؑ�jxmh� K�ɋ�]ՙ�``7R�k�Y��rf�8	"�o��g��e�əO���hi�G��X8��q��Ƙ�Ww�.��1<R��̓d"�Q��R��m��^�˷��wvc�EH#o������6�˅u��,ZM�ֶ0N�@\P
 #�G��1�7I����r�7�L�2��R?
������/����>�{?_���yL���Sza��eC	徜y��|/�٪q��Ii�-�s{�����!hLȦ�i���u
�oX�1`'8�d�)mSm�����)�xi�vj-}u��~�����( ;���|]c>f�z�9c�����P�׮���骈u�N�~�}�6���g�{#;�_�ߣ6iߊ��cplcXN(<��&�������}�4�?y���|���P�4#s�1`�z�iQ�.��n9� ���&qe�����sSl�s�K+�z,�Ϳ�oo��h
��˞����F0��%�3��=̖j����"f�p��m���v�]4���s��,��3S�����[����a�"�XFR��#����u���^Z��K�#� ���+�y���2k(�dKǶЉl��w𾭲�1��P�:�sm�3�!��
z���=o���{����F��;>�1͖�8S������ɭ��;[���$?HhgT�\j1�)���dN� S����H}=7�x���[B�Oa�2��˯�j畝h�S�"�`�-��9!�텩�=}����k^��	�$�0�H��6H!�V�F��!�ۯ[U��gm7���JOgC;Htd(��ګMo��R��sק���f�a�����Z~4TP�(SJ�4ЃM4
5 E�$S�ߗ�+��ʹ"��0��i���[@wf�g��vi��ᕿeǑ���ͭح��1YǗ�9�.�6�0�d��9�/�\����`iR���S�5X�;�0`_��E���ұm�����_L��bf����ҁ�] q�a�*���)��E�<���5�;0�%�uۗ��ڰv�M�Q0��߰?���ETi��,��$�Y�b�>&i�W@�j�;ll?6�y�5���#�ܿN ˞�,.`e�D��� � ʀ�hSe�f���d4G@��s�{3�>r�q�XD[�q�m`S��@��yii�:�Q��\��y�X�ڒ^��r�r7�U؁/( j�U?~=������S�4v�ÔW~^�~s����Npd��Y���*̇~�a�(�a97�M�ų|��J(���O�a^Ǧ]E��i�F���O��U0��u/��J��^�%{�&-��1���VЫ}�YyK�^�����4���g)ƹ<E��*9?v�V�m��Bw���������2�%G�����N�ͨ�C�������:���]31�(K_�5�	%��.�'�N	:�(�������|�bEbV�uGENN���b���:-��3��y���f�c�� I`� �
!�p] j-Uoi_�h�Ji�0\w+o��kW+1Qf�^�}611t�q(��@6w�K�o�lyp훦�DŇ�L	ڬx�M�R�`�CZ�'�7�g��42� ����"K�,u�����9
���k��XX����n�D����T��	�sk�����4[�1��s,�cKJ���ǩ5�T�y�w!Y�a6*��v�e����3��������9�s�wi��d��sV���U��q�X����Mw(�ͩ�f��*��4������S�_c8�ȳ�R�en�/�h��Ɠ�]<�w��V����i�1,��wEB��9ܸ�\a����b�D������X�!��]�XM���s^N+���r�<�����y4��Y}������9�؍9y{��@᧛̻��\vwc\�4e�7�)\GP�N[�.�ж�=G����O;jI��j=��z:n��.�&+Sqsi��+xw}n!�Q�Y+��WgY�0\��V��R��w�Y`&.��i�޸��e-��ZU��I���˨��Y�.=;3�WoK������x��j�r^�˅]X]N�Ys�oz�r�zi�O)j:t���pN>;��傻b���rC'��zWn߳`{����"����צ�����~�<~rlT�{�4T��9��;�ة�o/��Z�[�;�cn����p����C�]�\7l�bc��s��������쾐��y��fO��$	jٴ{FodM&�e��l��X�`�cxG�w���p�)��X�[�:��|�u�.�%�ڳ�cS�Ƹ��S�T��)�`B��7csO;��))Q���9n.�sXu"�N�B�5���K��x��U���T���wR�DR�1d��\��9��*H���Te'��Kӵz����&�Lʽh�k}�ɺ�0�5��m����}��}���R��#�]���&�-k���>��-�rj��%:٪q�S�X����H�5&C��P�N�d4�taM:aʛ��tV�F,�[${�8��j3�N�yiڶ���k�����D]���N5�����(V,R�;��:ѝ־_A}�q����]G�)��\��c��Mg�^ŵ�]�c:�2d�W:�D�t����o��v
���ר�,��������Lc�8!����ڸ�ufCr��O	��n*�n7��D��Yz�Rx
Y��D�E�d�1��^d�2Np:�YnJ�/��v��9Wk��NY��:J@�S��|�9d��' ����^u�N$*�֣N�>>���o�Ǐ<x��׮BU$�Q�Bs+R.;;.�A�l����
(i�.����|��~^'��g[���8��׏<x��ׯL� T��e�i����!9����<�����e!��E�kv���<z��Ǐ<z��I
�M�a뗎�w&��7:w��+P|�MMG��M6��8��Ǐ<x��׹$��E���u4FU2QKuw�!�QC�9'&&AE�B��#�DW��>�x� �����rx�OHFw�����C�G�c�;(�;rnWI�	���Aw2*����ƫap��&U'
e�i!	���4�Gt.$�)���@��EG
r.$˵[9\e�ӕ�U��p*�&P��UGAq� NYO�<M!�.��YOI!:h��*���Y3/��ymgw1��X��nVr�kzM��+aU|kt,ɴ��Y�����펆n����;���;��윈� G��h�gZ6�u�I�ce �.ؐQ��Y�V�����t�g��O��L>��Q0��&���Y���~�<�EJ��,�����ݥ��g*h?��.�A\O��߹�.>��<^|�mH¼Q��f�dg�g�B3"��b9���s�L����4�39�Y��DF����hȝQ���(P�qv�G���O]�}=��lq���!SMȝ�cC+��"~@?�ď~T�N�˿g�	�xRgn�E��,�#�fE7;;�vqj��u�W[��}�=o��1LZ��m�����!0W� z����S�=����t�%�b�e����Dt⒎k�����I�dL77��᛽����(�Nt�<U�1�ԣ|�r���xCʄG��'�+=.�"��HQ�q����3JUI��!]3�sK�cn�v�SF%��e���D{�u�f��VZq3q���!_nxC��{ ���|����M��qi���&���$]�
�kZZ��@3��O���U��*S���(u�%�β����߷yۮ^-ف��}z������g�"�����cG>��9_��Oܡ�����7�|��?���=ڕy��<ۉ+��R8%3
o�k	/�Ef�3r�T޽�0՗(<�����p�d��~P����v����T�[c��n�)�X"��R|E�+�<��ӕnU�j�B��({I�[U�ߏl����!�[5�
�(�0;�эkF����A�փ�Y�*"@���;z��0�����%p"��y#�wi�&�Jmw녊B˓ҳ�|j�Û�����
A��<���6��P��%�*q���,]��O"ݙs�z�[�����5���^�q��-he���Y�<(��.g,0lBe�Ʃ�{b�(u�+�&�Ɂ~��yd�|ݻל\�/;�*�]D���a���X���Au�pUD���Um����/�2c�s-��-�nͶCָ��OԀP<�?{�xdф�y�'�s�����p���K4噴q����YyT/w��&��=��z�]O [��<�J�D9�3s8^->}�;fD�WB���%ӿ4�d{�u���P�~\�^��+�!�j�����|�x�����~h�����+�0V�-�м��5?7Z��@�Bde�ͺ�CW�l��F��TZ��F�^,�2�����Θ���p�1͆�}V�y�g�CҎW��5������Z�ˏ���yיA/^�-����01���7�c4��ճ�y�16P�7��M����ғ_��#������ˬ�ڶ��>��o<�6agS�b�=xX�$17&W1N�����M�}��у#4�}��S(Z��+�ѹsG���Yv9	�v8̋�~xz�v:�=c�fFz�<��,��8�X��r�$ec��>�����u§w�]^���߭�kbE3���q�kcNpDB@aD\�|�\��{]��������ns���K;A�ݥ#��oN(�0����T���	��_W��C�1��B�OC�t��Pw�y�fm~/�#1I�.�_+p�R��-���b�9g>�ɶ��ř�d~S�~��H�/��r�ma�&��~�5r���#���fX���A���	��^Y���J8ʜ���޿Ŋu~���\K��L�qz���\}�ŗ��|	�`Z|����?�s���آ[�-����_3���j�tV��IX�n=U�M,�l���ަ�FS0�M��0�G.�����[�v���9�;E"�i/s�srA�au0	y��T�{���b���Y2����`%�*�0Ƚg��j�5���c��8����	��B�{�w�P����on ś�a[�u6�-�HHxXƞ���e!mk�&���z�(V�[)�l��zkg*�9�XN�w8��3&�s3������f�^���`q�t�q+�^p1LkW,�/G��,��
�O��C'�|`ɧ�x�il�3a��!�z�Yx�F/�"���*���7Cl]���:�FEF0ts�h�w�7�R�=n���{�e^y�I��{�x�N�"��M�a���j��u��)FU����E�b�^C�e$�=W�ុ3)zV��|ď	şn26;Z���A.�ORY��%�25�u�V�+J�S��+5�I�B?M �M TB4Ҵ��#�W ��&\on"eL�U|�1o�.���@f̻H�R'z���x�]��č�y����a���a��}А,lD�F,�ʬXi�xZ�]6��-@����{�ɸ�%��b}�KF`�n�v���a��:���k���ÿ�S������S���^�k�2*���}>�hO�Ó� h��sD�%�{՗~R��j��^��0�/��=��^9�f.�o'S�[�c{.�a0֫�/m@{��Ƒ�*���mffl��Ϗ��T*]c�\y$���yȉX�{���A��\T�r�O������A�����0u5����;�b�4�S��/X�Æ��kV�76+3�b�5���Rj 9�gO@s˾�'�͗��n.!����Yw~�
�(�!��+���Y&
[�OO���1{%�٥m�g&a�I�{[�72�1��o�u5v�t*v��_����3��-~̀fԻ@��Q�A!��0�j�7�'�{{��z�rI>���&V!65��o��}%����JTC|��o��;��,y�D�w!�"ڰ̌�z}淓�J��6.�,*�Gi6+S'm>G���/�����6#��Jھ[jo �����f��47yd�����+���]٘��e\�i�=��]�ޝ��	y�e��8V�u�Mܜ�y�������'�%}c�ҕ4�	��� �[bv P�6�.��b�L�-��8t�֘��8�z��ju5ț ^�/ruW���q�Gx��2�^7d��3����s·>��yN��v��Jo]�ʆy˫ơ�����w����n�^������#ҵ�v)��D��	>7�w��K���w�����5�r�71�V��%��<ʋ���7{r;6t3��W�;�g��K�7C$pk.��}��rzb�s�Q��f�m�3y1!Q�[JR]E��;[��X!���XO͍ C�ٯI�Y0L �w��n/��%6�^}�L�[{��G�z��ۄdcCL+�޽�pe�7\�M��c�{F1��{����12%� d��;:f�o�X�D�g�ͬ[��|���~�Q�	_.�S���$����z�t�'�B-��_�{pw2�&�:�qp�͗O^+==�7
��4Lkav������4�C�w�}�Ҹ����yu=���)�6v
���`�.%����ަ|X� ��W�L�a8�{_���K� O\r���1�T���%^���nj�2�:�8<� �<ϯBL�"a��}+򿳮�ԭF��g$��v���������lnq6b�ظ�U�s�wOz�S�����7A}�Y�$�]k9�y�rR��A&2'�c7-����6�W|�tP	s2.�J#�_Z��f��iY���ڮe�o��b�=��=RC�ޓ
;��L���H$i������<����7�
��dG��&a���`f�,��q���]�-�Q�-�OWTd	1D��N�Gu�����|@KJ*��~�~��O�~XmQe=����˰���`�[��Z���N_}�H'"��c�0�7e}�:4�1��0vE@�5r/���"�]�e�����a�L��Cnt1�h����]2 �����d?J;~}�"U��,7�z�T�vlফc|�)C�z~���y�x��$ϧ�+�Э{��y�6���o̙�VQ��VtPx��|��~6����WH�o
���
m��k��N��N���W�.�eo�b���I�C{K�pm���Ǻ�ts�|��/���=S��Y4Z��හ��R�8̱N��ޛlⶻ��?����i��i�����{Ʀ`!{�+� @��.�A`���Ŝ�>J=tD�L/�T�޺�2���
V�Ȓr�5��lh6�@����#	��w��BcY �&C���U�TU����wש��S���C�:�$�5�S�Y�X>�	�1_�����N�GSBg�{���}j�ܢ�|���N+�oNㆯM���d{�rL^
{]���;���:�]':I�Ȇ5�Q@Y[C�7x�*�Ȇ��Ĳ
��/�E^5��[�}ꈓ����2�p�`��Ȩ�R��C])A�ـ��w�i{6�e�w_����cL��Mئ
%T�ue�w�k߲>B?f+CiR�h�h�� � 0�����~��9x����/J��w�%ڮy��o~1.��W'N��u�T�������w/���-pa��A��5��ai|�Qٖ���S/�7�!�Z���	�P*9�lb�hL��ۛCr,��Q�B��D��k<{&�y��a'�/)�T�����MC �(_N���^f��޺�k�ۍf-�Gn�^?�EK���]���(ey�$��m�Ɣ�-��{���5v�����1�\B-�;~�������ꅯ��;lCvlo79`����ˑ��d��L�y�|�<^v~~������������PW�#u�g�L�~?0� .sKTf;6Q����p�/-����O�g������c���a~�\g�s��\�ZbL�*�2�������U��D�ȫ�}���cM���wjN��P]6y_v�����r�}ڨ<	�y�Q�}�^��k���Hr��"�����f5:��8�q�lz�t�y�d��R��f��$n���`5������:�*�v�V���9�^��Mt&ͩ�\WbSU��6���d��[T��=w�?g��D����·N�w'b�fdg�
U��p��<���dd��)�o��m��^�Юf.��f:>̲qB!v���3�}�Ĝˬ��ޣ���z1(�o�(��&�+���K��0�K����˯p)W���D Q߭-hGZƐu�bEb�Ȑ ��r��o>wߞs�����v�3P=� ��o�e
K�����!Ϥ�ߵ��X{��K\�i�=�mr�앸��Z�7�l{kd�H��Lk��|{��,W�q{�j~�"� ����vv%�ud�naFi�tu��`�mm�YV�Z�+��:����q1^*�Na��K��R�"n5���j��)�6��5k��Q��F{Z�T5�����7Pù�v4c��c�=���(�iUΥ�!�y�����q�+v�P ꕯ�_��5��E��(B���1���)D��]��G����ʢ�ߨ�����X"7���S&���dK���Z����X�'����~�r��_פB�m��XA���yN�ا-{�.��:<���=\�\�⓴c�d����C�SH��{q���w������J�
 ���]���O������-�Й��X�v�2wT��q��W�5Y���֞1M�0mlwf���ݭ��O�:���hnR7���#K^�A^�_Ky�z=0XeA��q@'\��+��&>^$3�����x/�^զ0�G1�j^7��[��VԻ���σ�P��qv�JUʛ����٣��+�z���n��o�-)�����r�W{��z�Z�r�6��w���G���r�
@��V��_�qc��4�JSM	M2�$Y�dBAd����{}�7�<�����ݚ�r��<1�-�k�|�)T��1L��]�����FO�gww)�*�?�Yp7^�|O�:xw��|�4{��W0\�=3K,4��n��qk�Zsq��ni���]�
�5�(y��
u�f�)�������҇k�&P�^d��������k3�4rP�s�g$LDI5��C�5���o|F��1V�e��Ԩ��IE5nLٱ�,�vd����ӑ�ߩ�`�f�7r&�J�)�*"�C��4CXN]�~疤� �	��361�]��Ȝ�5xƦ�|e���们7��y�.�2���]6a�SA��o��>�e����(��O�|z�sk4d[s!��N�yƼR�^�x�7}B�rq�����{aي�+v<������9{X �����0�n��C�8`1Aן7�&9?i�i[�=���]�6^=۳�����UxK�o8SU��O>y�Ŵ���5����t�L�2�Hީ-����G��v���Ph�Ҳ��}��~�&�1s��"�Z���ݙ�?=c�x�#���?��G����h6�喗\��{_f{4�ȫ�[��H�^�Q©����Z��Y�]�yz3)�:n��kA|4b�Zճ*�r�:��άx[:�խ�^ɪ�tf��v�����C���������LN�����]��7۽S��$�i���}`-f�hp�[�����ͫ��lڵ}��|���	S�gs�"gΎ����K燪7�F�O�Q�v�.:���uk�wCo�{�!��lOEGs��T��B�X�6�������Q��N�!k�,�ɡ7$��X��.����3��ž�a��n��*����Ce�zb�]�oO��v�G��%��P�?�y׵?���0�����Q�/������s/OFR��Ƴ
�4���m�ʕS���C6[�GS_~�|����G�������զ�B�X:���,��/��]"�<���oeoW� |��Jje<|�b�r��O��2c��b8��h���ߞ������-X]?&��+�w��5!�@����a��L�6���G��1_�Y]�����hU@;���dָ�P���>3�y�n�KH��zn<�WP�va�	�Ķ�G�MӱZ�.��+�1�������MHlSt�O����6K�	���6���9��R�M(@��0�f�_�:� Oò{7v�3x�	j�Փ���&^ӱy�4ԓ�N7�BVl]⬹�C���xK�!�ο����ۖ1���r��):wS@��ZbK+�ᥜ������m��.J��v�Cֳ��S��KF?R��=E&�'*�Q������F���uf���*J�=|�[�2��]y\^uT����<�mcV��֔Ż[6�έ�/`4�0�LRټ"1Z ��VK���g"�����2��ٌf���`t�2ӌ_�{nB�SIlZ�h]q�V%4=�s'�uk�����kEQ��ή;�=��N��g��F.���Z�2�UEN�Q����X�Q�΅u�'�9d��޳�&��6��%P*��M��|�v#k��W�z(4$�b�@��9�쌿�d�U�ٌ�Ǐz������n���$qiaw�>*�ub��&R	[��fh��J�����>/N��n��ֲ�7�S͠\������4VJ����pb����$�G�#9EQ�[��u>�+�bF�x��M����G��ݙ��e�7�$鏶ܸ�3�9UuE�1�W�gl��{���s+F+�����ۛN%%���3��tp�\z��X���4T�F,̻O�u�朜E���e��}��;CO��%�-�ݻ=�9ݟ3�;�g�sRsV朐��EJ�2W]P�X��K�}|i�\[U�au�����0�W�-�9�r�^�r֕�]�W�M����#�y�X�f�v�� ��e̡y���rЖ%�Mk;�"9���zo ��Ph�M���z�IjlYo�XT]����.��J=6̙�o׮�!V���}|t�q`�orȵ��q%J�K؍��c}Y�c}bī�<׍���e����Z֩|���[���ڔ���{�^�,Z�^��m:ɛle�M��ؓ�R,��70+����;�W��KWWZҗF��\_'���=�8+]�m
_Z��`ʩr��f���H����D�x��U�i�w+���@���Ԝ3�X�.t��/�W4]�wN�c��V��'e<�J�:l%'X�j�^շ@��vJ�W��W�`NҶ��Pⲻ5콙�T�{77�hf'�O�h��3B*�I۵p��3s�E�Lr��;K%��ɘMC6�Z���7��'�{:��c}v��q��S�B/dǴ�,���c�k0��b"��jP�����Lźcu��ɖ7:vҒ�Cm6et��;5��ot����!�tR�ͱ���ƒR��n�떯Nɼ4�f5�����'�5ܷ�]n�Z%��=}:^*4�z�$�r�T�#��YmXc���=V��M��}a���6,�5
�*kj�%u�܀v�v�*ؖ�V���E��&󝊅��L-r�������+sO�S�d��ܽ;��z����v_b���Y����i�����!Wu�`gx��o4�q�=u��q��9�>��s/UjcjFє�n+Ghҕ�^v0�ܦ5pq��f�}���o.;y�}���4�6������A%]ڲ���z�<�8ԩ%N����L�(����W��n1��N� ��t�_�"]To��o'���y��k��lтp��0���8P=��B�ˏ�*�@��;|q��O<x��ׯ�|q���hRM�S@��q�#��
)R�1kv���qǎ޼x��Ǐ^��7�e�P�d �F�rsȧ#B�����;s�˰��yݻso�8��o^<x��ǯ\�P���Tӷt�����r�����ג��"���s�5�N�q�<x��Ǐ<z��Z�MA�˪*|I˔*:�<Ƀ�����w ԇQ&\��p�e�CߞvE(�q�����U�3bT�Hek�+
�,�JĞ2�Չ��vU��v�rԞ&��q����ʉ�.��*g�zRNN�r�s��:�v�@I'��&SU����
9�4��pr�k�r��((p��9!E$�ʨ��ɏ������GrN�wA��P��$0�)�!���e��l�'��$���n�t�������},�	Э�1}��d�Ű8��ʦ��ۤ(�6+L�i��РI� �B��BDP�0��#��MC#l��-B̍�)��b!#��HJ��Lq���߭H��ִ;:ыZ��#����gp������c%��Qʲ�/��Z�O�����g�c�xӟƶ.�x@؄˯�S����/Z�����p���	u1W��|���&�T �4�w	��\z44�Z��PKӼLc�m�a2שb;W�Zۨ���Y6��ͶE�hB����˃��[��]m��.��&EZ���B�v� ��N[�I�r�m*�7T�C�綾�4x��'֡&]�b���3�>U������Mh�����6 ���Х��a�9�^= [�G��ְ�s�
ZD��vaW1g.��4�n�[o�CX���|ຎ+�,݈�
`��؅/P��3^�"SԤ]��;�pb��D'E�^L����BgL}v�������ץ~by�K�����/M��J�<�6��XcxJ����'G.�z?�(x��f|�<cX��&���syoϯ�?���ܿx"x��!+~>i��y#����f/�|�ӳd6�a0��D$(��3=�qHѲHҙm��g��c^�B�������u�b�oɅ�s⨇�H�NO��T�\G_�)â�}��`�h��t,6p��%W�f�>�G/���ʇ}6���"��Z��n���@e�f�+�SƷ�~����t��
��>�<mk5Ϫ��igi��:ݗ�h77�H힫v9`�D�е_	W��z���[7+���oQ����xkF��[~��,i� ���� F�*
�� �z���uk<93w��*򭁘`sN�[��X�w<��WK^O�V�� (�3U��";Y��l|U��i��l�����+ɳ��H��̠���c%o|=�~zٻ��<CFL�YW]`����)�<����zg�����>t1xZe3'���!u�0�R���s��oN�"[r��o��]U�biO&)CK�a�FZ-(�KϮ��(V��1cO�Vf	�N�	��]��*6 �(U�7#�1�&E��%փc����"������M�kKDIԲ�Y�[�זEk��`KX�Vk�g�ô
k�e��������Y�UwԻ�����Y���k9�'�����Ӿ3�I�ι��NL��������r��z;���
�^�}�
J��tfVW>ɹL�d�v�W��M�V�;�o"��\M��T��h����[IدK��à�L^%h�}�Y�o�W0>9����1i��+�]��酯����tX�l��X�iq�U.r/2խѨXw�~���|��>�D���=?yB�g�6�VF���)�_��f&�#	ۭq��.���y��7{�;7���y�!��쫣�#��2��+�	�]R��WQ;}�@���=���c�4�v���lǛ�kOWb��V�i��I�{K���R`�B<yY�YGs*[5��܌�2VJ�»U��$���Zӳ���-ki��FA�sU��Ϸ�/浟T}i�5���z.By%�%��@=}i�����
]צEV��8wfL�-Z�#m�1�fW1*;z�����^��������hm���S��q��z�(�"�4�OM�\B�'[�B� ���WPƳѭ$ή�f��H:I&�H���7ޣk�I�k�^��捰�tt��%#f�9B7���c�c�,1̉y�F�:�ߨD���O�L<\�??
?~W��gs�u\��3�|"�8�!��̻[ k�<�{S][��r�Cg��4��R�{|P{����^K9/��H~�R��|�V/��WP��c5�.�r�q>V=�\�mrw�8���mv�Σ��[�wLKy|{�#X�)�++ߓ����n}= cƝ�����L�e\]f�[*�^����wg���F�q=�1[�m�*�J�~��z���e��Şf�{%5�wk{z�jy���a�\&48�
�]X�}q�'���O˨�9D?ּy3_o�Z���	�j�/��l��X�#j$����-y늕
|whg����޼U�,�j�g�����'~����3$u�ʈ�v�
��ݜWI>��eÏ2c���W�W����fT=UI��.���܏J���)
�(�!�~K+������=�Z�WV�X���c�3d�&�,�����TB}��(يA���}W�aw�p���k�`���Z$g��xy���Sb{zʚR��|.>O��$ζ��a�L�`)��{��k���
�2��w#��WsNwW�kT@L�㊋l�I��]������a�3<���Z��>�t���ڻw�8�K��Ӱ�HKO�3����5��%�f�"���FC�y;�#�ҘN�In/��5�Suc6Ưv�V�<�]�[�-��ˋ8���hs��v��C����2:.�]L�̷�G��4 ��˭�`�FM��1 [	��X����C��;F7W��\C�MЫ�/*%Q���K��T(�I�;.�h*{���P���N�~���	�V:7����h��*�pI���w^�`Zl��/.��������9�x4Ɔ4�%���5-~��]�o]����Z�k3!wa����Ї�f~"5f��r��&pݼ���ݮ~X�>g���D`����op�^�����;8֗�d#^��Ȉ��,/��n}4��5�'ۺ�ݧ�FO:�~���ӣ��'�;.���(92�>M�qx�@�T�w�T���v���.�</_���ś$�,�!�?�����g��J�U>���J��}uڰ��ͫ�t�ƫ�����ɍ�'�9Y�/�1�	��HU��a����ǣ�jZ룱�Y0�u[�]�n�};�9��)���n�'���眺�vݡ��H ,�J�w��o���ѝhZ����`,���/��F�Ռ֮����מʼ�l�B�k/j7���zf/���,H*E��J+��-X����#������8�V�k{mFܽ�����l���A��<�_Y�lpcC��\���#��\����#b[JzU�����j���͐MV-�R��EM1J=��&�`#�\=�	����?K�G�V�;X�s��m5Ɇ�R��9�Xc�������P)H�v�)�{�O=q�IU���#�YGY���{������X�Q~��H��ߒ%c�=O�]��^	�ET���0�wַK)������trNR��]cx������t>T3
�Eעli���"����u������v����]8r�����*y��&i���L�Ѽ<P/��P���P��߬K3ǸJm�	� g�(C}���#!1�'��� ��g����b)>5��IJ���@jy�_�1	��U�fV�٦�aXD籄�p�k�)�l�zl�U>wv⫓�Q�n̸�mׄ��k����o4z��1�ˉ 
��J��[����Dm�{�TQk���W�:��}AX��*5���)�3hUxfK����"�J��V������l=��`&�!��*�W����)M1v��Ԧ*�8�n��J�Y�������xU��qu��ַ���$T+��U����:Jg3[Y)�ʂ�,�.'�1[��X�{(�}U�u��k_��~���/!)�1��2$����g�/痄�}}h�'�tO���ʄS�Ƣ�L:Q����7��k��'��M�5�ʲ�y�q)w��A��M{zg�����=p�w���CV
�~�`'�3~�-��ߣ�M�W����rW�n�� ��!ki_Rc|��~�����^ �<���H�3!KĬ&�ۗq҃/(���$�����[���#>ڤ����r��A�=
��*�O�4�؟��3�.�2��ܲ�����H;�9h$%3�?������M#J�Y][�U�w��L'kua�|e=	�&-�X��hp�|bٗA�����cR+b����\�>]7���ܦ(Tm�������w>'y^C�
i��T�
�9�>�k=�o������8,�fO�ץ�,^�ƱS(�õ��*�׎���u���xZ%~��rأrW�i|�	(����I����P��Vf*����\�1�m�v�d�Uz��3&%���8՛� z�x�jr_1�~�m.�[��5�I��7{{|��ͭ���(��Zt��˦���S�׎�=�>�0�m ��R�raW#/��]�_���.}aXK4S[ѻ��Y*�"������o�Ue���Z0Ewrr��|���]A�,��XM��=J�5��]�Q��,��;�)S�[���*�zn�9ʣ��N��Jj�Vf�k&{����PSE4�� S)0�A�;�%Ҿ!�:-�wA�#��R��$})����U����ǀr=2=��*)�dr-���^�6;sڸ�hf��)֠6 r0]�>�U��Y�j3�YZ��]���qX�:�a1«��w֠�4�t�^�7�W9�U�{��Q�-�t�/������|7�
N��
iz��5�
ކSM��D��Z�-���}8�~��@?t@���ƻ��}�T����/�J��g^�"Z��w<X_<0���&]~~R��ό�W�*waΈ��D=O?F-:.09����Y��׻����^���kW|d)������ݮ5�T����mC�Kt�1���JO.�PT�21ҞH��-q�g�dT�ß�ꖯ���9@���w9CU*o�9�����DuB��qH���r�oA�zc�Cc���2%�׹ٰ���۲���C]ٱ|��>��K{ч�&���ԇ��f��טf�l3�y��ҕIoSUm�2�!��� k�*OnR�k�Q,��cg�?@߄��0�bR�1�7���>�  P[�\���-�_�/��p˱�0.q_&{��4�T7inQ�*v��k�;��F�6�[ab���+҅��/ot.ei�X���@xU�s��n�F0p��'��:�gu�0��+�J0�6ss���Wg |�w��h���iB�Ul�e=�3��8�=�ͽ}N�_����������yݛ�fa�W��bb��Y[7�wA�5Ǆ�]9���}u���-����[n���1�����בSى�:����ʚ��7PFD�חM�yە�ˎ�|sq�@��F�k�o�1���!1���ۡ�&��t��Z)�i��8�~zW�~=�a�?���Y-!��|��ZGaP�,����oc+��*U\.���Y�fz.DF'���^�����ÎȤ��\m���5�L0 �K�qs�N;3*��Tx���@SyvE��׶o,�Jq�V�H��I�x�YN�nn�Db�<Be�pTc�e+y��2����S?��|�'
�j�Pɏ1e�5�1I��6c���\��4X�M��'���;G�z�n`;1Oq��@������Q�=)���/p�5�	��t�����r���/c_Q��Xۡ�wE��m���qAJ�hi�Ǣ��;��x��J��cT���-��Y9��_��k�'��Dr���,�Z�a|���<e�3P;D|��X� 4"���ޡ���ϴuگ�^���̥\�
�O���7�l��$��Z�yy��2��%��B�Z������^V�?x�.�=d��'���i��g[a��c"�wknJ����~�a�Īn�z�My*5V�g�J7z�U�ڡV7�U뜰�9������5�*C�.ݴT����v�m8v�;6��J;�]����Dɑ��E�̢���Z=�Ҹv��Z��^Q]9on˽m�]�yޟ���Zŭb֋Z4��b�]Yi����g-}u�|�0�̙���z��!��41��(����T2��>Ex�@j�45�Ŧ�!��������>,��,�c��y�0p���.O�݀�N �g|RXV�zT{���K�����";�L��b��������/hS�|�t��KK��,j����Ȗ=`Oׄ��__�ȫ�1?TJ?�S2�MW=�/]�1���c��gy���Z#�N�3�;������F'��&���뚌n�t5�[�w~��K@�mJ���t������a��6y!�M��I���̓����}u?U$j�+�,e'���@k��캳=ۂ�3����|s���юv�ob�J�ؼx`Zo���U{lP���L�܉���D⹈wܦۮ�z�|u��%�C�
�ý64�k͵0����޸���z )��v/~�d����٬��ar�sfks{*�6��x��d��3���V���:P�O��(	�l������n��[TK�sL��L�ؘ�ݨ��:ںk�Y5<�
^�ځ3k��] ��A�bO���, � �����S΅��'�n��ƘG�tf�=)~����=+RL�J��6P�r��t+fy��՝����J�1��Һ��&�ܠ�T�ZX@^ G(#�:t��5C5�g[m	���F#Dk{�T
ྻ�BV�h���]}u�t��+[{��c�|}���||��'X]�Qţ�U?�؉�L,-WW��TKa
��Sm���[T��IP�aq�i�	��s��έ��M�l����oB�/`�R|k*�������Tc�'���o�)���]c��a�Z�6ɣ�w�c�!T���,C�lҝo_#"4quKŝ;�-/-� �W�ۚ�~w�����:�6�r���-�CC_8P�X/DAm�; TDZ�-5kk��=���sv��� @|�X��0ŕ8s: ��m�k��l?�}�P�r��Λ�J43���Ӭ��5ɍY������{nKJ��!D;�Gy�`�b��n*�G�1�2�آ��[-,�͞�..?��Wj�=fWl��td0���\k�G���!��)^l.6�]�t�ට���m�}�'�w�q�
<4 ����Ezߓ��DX�wG<Q7�B��x��w��3��n�~>��l/'���\j�+�3�����o6��<��ㅏ��!^]Q~T�uD��{��4����g����NFFRڼϘ��~7�
��8�eϤ���,�>j�T>�a�AU���[#��~v�e;l-�*�˅�%��4]8�Vo`�E�<�:�y�%iA>nReg�o�g6S��ŏ��p��b��h�\1��&�������*�5R�;�a�K7|�Q�ȫ�ɦ�n:��r�]l��hɇ�z�oۻԸ�j�;}���esr%�<U.��r�v%Z��[�n�If��+�V6R���+v|�N���,��)p�@tR�T�]^,���R}�_<����ú���l�ۨ�r��&K<�)����P������b����Eˬ�7e�#���\	��zB�U�M�]Qv+���%D�.���hI�;��!ٶq�h{��|�I.�-�r4k����� J5�2z���YGM2��4&�5k}7��u�ftбں��r�t��t�mʚ��X:�Z�%A7�_b��H�����È���Cj=�̻Rr!�S��Vn�VJֆc����N�V���%Gy�"�p���{3_B��%�E�h��e����p���j_�:pU=�c2��ªt���Y��-�v�Bsz�a�j5W�l� 6k�eS�ԙޔ����%���u�^�}���96e�tU���"%����� zͺ�vf�q�vn���n]O\���.z�1!y��Wa����r��N������ݪ�M�y����n�nc��d>��)�yj*Xjuϵ.�p�۹�Ӽ��c���Kl�,�kj�=��J�/G��� ����1��θ��*6��+T�{��F�_�?�_�W�!��H��H+�V��5œ����jA�</�G�˭����Ǘc��%�$Ê�g8FB7)U���3
�U*P�Ҩ`�ӲT�wV��c+[䯣���6�Syv�U�eS֬t+
BJ�w|6�'�Anqk�m���xoDN����n���6�x�^�bNT��A�X��'Q��N�r�x�,ֺ봌�nRkyH1��f,h.�i�x0f�vBqY����3���Q\�`�����yz3j`u0�9uQ�Ls���oZ�a9ۯT��Kàޗa{^��9[�FH�TU���\v�Y�1�m<Z�k��o>���U�ev��	�V�o��={�U ����Ț��)�2��f���Ņ�e�����n]H��c��+J�wM���������r�s�.���1�u��n�Z�<u��)6t�m*\.������Q��Y2�ho6��Ve�\-d��bF�-[|Z{]$��r�R����U'r�Nb���ŎջS��g��O
qf�0m_*w'wU�wjf#�خv��U)��=9�!�n�����r��\��iǇ��x�"!�І���\����ӷ�)��$����H���.����c$0��S��~��B�@#�|Ȉ��ª�BU��v4ӧ<q��o�Ǐ<z��ڢT�O��HJΜ�G"wq՗N��N�;�/ޭ�t�Vu������;z��Ǐ�z�=��HH�Q�ӷ$�s�T	Gp�sGA�:q�q��o^<x��׮N�PǓ*�R�' R@�I Ԩ�@�P�Tz��qǏ=x��Ǐ^�:J���j*{��*H`�Rq�psȳ&!Z�L��#QQ0������t������y*"T2�&fT]�Yr�7YpO$$��UK�H�\�nC�PE	�๑Đ�|t�3�������)3&\���eJ�I'�$�{:����ΙˁI'i*b���l!��6�]t���-��E��%v����c ���\�.��;���u�z�����������|����v��{�S�C���ʥ1�F�u{���g3�9FS4���e7r�m��Y��v�6+溆;�]��&���%^�a�R�1�	��+u8�ow�ӭy��؞�K3o1r!���ne�� ve����5�W�iyoV�0��!�%�ȗ}���
h8��1���dl���n=y;(rg�y��=�E�߼�(C�P�ߞj�L��R?���w��n�d9U�.ؙ��oY���I�h����Q��%�ҩ'�P����yK*�kW#����p�.��i���MoV�<����w~g�ր�Ez�f}�ӡ�����C�@Vn��M\u�J�}�g��o��g�x߼o/s�ܛ��,�~O]0��U�]0����1�x��
VZL+�Z�]���E��~��x��r�e�l�_�X�Wܤ_��=Y���
=�D�Z���ʣU�1sC/�)�/�+�/�H0�R�G��T�")��O��I��Cѽ���vk:�d��5�ք�n=Z8��z�(n��>hnsB6Y����(d��R�X��[�ywnV'�I�ɓ+�s]~2���+�8���;�._z+���!�-�Z��&��T9�Bh��ղop��-e���$�p�2�U��=9�̣y�;��j�%�]*�ι9܆n��X��a팤�3�˗�J�ߑ��SMSLcM9;Ϛ���Bc۳�@k��#�m�'|o��ڼ'������ަkɏ ����'0�GS!��D��tձ�Gw�)ݐ~dL6�B���*�NP��ߋ�	��h���D�>d+�zk�'�a����2I��R9aR��y<�\�2�/ߖ~L�O�X�����������B!��+}mGS-Vb��N���Z�ϱL���｡�i~Y�=>�A�rY��^UM;�|��'���[}&n�w���a8��	��� �	�w]>�^h�j���L��J U�
�����0����Q)?^8|��l���<W޽���5�j}��_s�������@��5󚼾`q>KŨ;��,k^N����ئ�t���c�q���<6YY�]R�9���T)�z��������u���eM	��=z_�F��S]�{1�nE'V�Kk��=���a=�W���é�����
��Y��Qm"K��r� J�>vj����I�=�a�JNؼ}֍/ka�h����]��z!
���B�ѐ�hy�C�j�:d����CO��f�j�ϯI�Nk�!��G{�;k�-��`��!�wXj�nG܇�F���'�^~J���|{�ŵ�b�çEr�V������]��Y:8��-I�`��ڽ�����EۅfK/v��y� ǂ�T�;��5k�q����&�A4��^�����|>
c���H������WNI#���Ir��+	��&q�j-f�{��jٞ$�u>|mx�b��7`��*"G8�y���M��>���ML��Fn5F��x��X�]��w9y���T�N�+7���3᮵pK<n���������}�-��tvN������K�mW0(� �����8��)����+G�a�4��e�s��̗�Oѡ�Q��G��B��r����Tv��Ia8�����7d�6��A���Onb��$ ό���z1���ꨦR#'��5C/�S�ז'���*G6�.���e�+m�Ե2f���^��.�C�t��־���,����S��	�l�6�`U=����g�@�H��D�6'�s���W������l�<}���P���� �ucs����Z�ف@��ql���������9���ȈQ�πm�����oo�Ļ�3J~�)��6�U���	۞���<5�ߙO�,��C����)�%��J�ѭQ&ro��������˓zm=H��g�i���ʀ��KXd��_��iz*=�{R��F_ug�[�������reA���v1���j���,$mQʼw���i������b�&�����W�^�^��}MI���f&9�EiXOie�r�&����S��%;�ivꭷNٖUד=���A�F1�g֊�9�s5ߚ���g�M B~���M4��uj��`�o!5ɹ	�#�({]�2ԩ��f�n��T�Q��0��N��3.��mma�εC�j/��<.=>�r�������%��05���л%�U��eL/͊�6	3K#%����XQ*,�_R��~C�ɦi���ª��]obmy7��t��n����=�zm��N[��O�5�Tc�ީ��]���&�w~�����s3
��;}�.h�k�w��D��\�㜀�;C~�����W1��LB�v_��������#N�:�K���ϛ��s�g��yOm�O��l�h�j�3A�?���z�vڱM_�n�I��˔
UT�I%���>�e�<��!��x]N>�?~4g����R�_}�g o~_n挐�����u�R��>8��,7�	�r�Y��-P��[%���QQ�ء��;ؠ5X�e����1Ԃ��5�ο/k]�/�~@2�|s�)�R�:foM5P�n����Ug���ى�Y�[	�3���>�5�>�PA�p�lakz�Ik�>c��?<5��_܎�͊}�������4�9wdKn�=�9�M4����v�-����'Js��N���$�d
�ׂd���2vΘ��D�gǋim� �6\c8�v��p���\�������Q\1ۼyנ��h84]������w��.q�XՉU�+����O�c �c��3�9y�gK���k�X���~�aS��:w�E\��$N0����|F�g|/;[\*�lG�o,�?�s��qH��-��_����2���1A���b���gZ{Ɖ�
�h���؊�i4O�=;^5�,
1���g�Xh�Ӓ6�ti���f���.�K�9�"y?|~����$��	:�>��G��*9������cl. ��ۙ��Z	�am�8���:y帶Xf���5���we.O�%�ST����SE�T�KJ=c:�O>�p�)b�7�5w���}d��N�ú�"w�m�ʿy�uG�P��߬�����)��''N��Os��>��nne�H+*�������ɣ_��%��1J�Z�c�6i����0��5�	qH�;��aq�̛5ռ���ޏ=��S��at�8��`�=�=6(fb��-8/�����a)l�K�
�S��T�{*am7���M0����&}]���<c��^�Y���>�C'ڸ�k��1)֣��AJ3���6�T9�ަ�+-	iMmO��B�w��������]�Dui�]K������v�7�sy�Z(�Ihj<�{Ýp�TN����l"���J�����w*5u�����9�;�L�E8���YMSڸI���9��V�������Z�̬�&Ǭc�>�\�;�7}:-	7B	�^�}~h�$��	r@��M]��\�v�J�0�$��k��sd瞠�VR�?{���5*��PĞ�l�<.xd�ns���33?i2�{Q�/^�Nnҙ�gf�p֌<yf�������~s��8r��A%��yW���uҷY�;�:�ڨ�gU7q�+�&V����^?m�3�\^琟:H_ǁ:�@�d�=@�\3�w;��O�ޓ�ŭ;�!�{�2t��r�][C��C�	5� q��-��0{�6�Lͩ�눺�n�P���;��������Ǎ�[V��O&�ɌR߲���b�����.�����d<׀9�4Ⱦu��@�f��j+�+��k���|�v��f/#::4ܠ}��eε�t�3�z �~�f{��ƨ
��q���{*��x0ɣJ��=�xP��
n5���h�d�Ey�V���>mQB��:j=�W��Lٛ%��+~嶾"%u��7��G�(A�T4��P�x��t7�5חMü�6�'���3�<�4�����i���{�m��2Emv��ɑa��n�.�!���|�s�df��n��-��M��z�1z>�`Y�,K0�-+�3�l����Ǘ^���S�vHWGmv��]-�p	e0:D�	}��	�h0nK]S�jn,R﷌~F���ՍYmEfX��{������|@��>�]w��v�x��d�f��'��`i�N�G�s�ZGA���ޏ䬫��V߷�e�¹�yP�탥��a �(�5}3ӧyKvy���G�dE{�'�q�5�5S���ϯC�):��A��M[�v�.ڧL�[,�2�Ύ1}J!2��������	���_ּO��ޞ:����)��\1�G&y��i��*Km�}�����ה+z���>��b�3�xs��{�60�CNѪ;��Mۋ�r6�T_e�����,���Ly�(�'͌���]q�5R��������T	�c��r$2�81����S���/�q!-�Qh.^a6q�[�=��d\kCO�)�a!����u?f��r�_��G�1��.���!-��y/7�"�����\�X�6�x�Zyl`,�x�01�d�[��L�����Ҷ��j8��6�b�sv)�P��)6��r��ŕ�Ș�W=W%��Yې�<��$�U��o�q"��������G�&Y�����9)�g���B̉w��;R^|4���3c���ŗ�6X3�x���lo���g��LZD(Ɨ�%���uP5�
���_pN��	32��2X����ǽ9�N�'��U:�dL�ƺ��l<��y�T�-o9�2�k�A��L#�U��})|z�:-�x7��\�{��\ٜ2osr9ڕ$�w��ڹ;ɬ9,�Q�aV����f�e�dV��>>>o7��>�Kz�,Zf6�g��q�������v�d�_�ӳ%�]��l�h�\0�Ӷ�ڍk��;�����1�x3�ב���4������P
�q����*+TK���U��<����y=�Fڷ�]ʹ�k�+�C���c�kǤ�ͯ�t�,O��`�L�:���!�ϯ�DûJ*�^bY�od�y��j�R�f;�>wp"�k�G�~|�=�xg�u=��%Yxڪi�Q�k_�vy�Ԣ;�_��?�U���z�Y�履��Bh&e��Vy��/Y��2V��U����uT�14����׺�DQ�=�_���=,�
i�֡����B:i�g�M��1��6�Y�5e�=�V<�3��������I���#��D�䌊$�6/s�p����'�@��hV�w}G:�dF1�3,���)���a�E�mH��l�d[ǠY�����#+Xr��z��Rs�J�X|G$GoIDP��$X0k���[V�K&�hq�wƠ�i��lm7�Q<��.�(<d˓�s1&�"9���zG5�2��@���z�=��+՛�l?6H	J�ֲ�F���x8�L&�k�����C����׳���Aj���k+��!�/�k�Q�Yv5Q�ĨL�o+�XLE����V�qr�,�r�z"���w65Pk�3�.���C�7��2�ԯJ�FJ�[���cdl�g�W�!rq��1�c�o�����fy����)��jgS����G�sz�<UoyFD�l�m�k�X����#�wo^��M̆�;�)@3�B�'�@���]I��[Y>�F�����"�m7)4e�Tm۬��v�Ƣ�W��S,H2��wf}Ͳ���^� �W�b2)��_��0�g[/5����+�B��甶����ѧ`��t8�4�����8vy���0�����L�*d��4���O�68�>��z;��f��b���?C���-Н^czB\j�3<���L���W�n2o����:u��j�OZ��r|`1�F)>m�m�O���x��u���ⰽ�1a����P���t'8��cٹùd���=ɛPl��:K
M~�q�D��C�A�eG�gD����ą�ni��Qœ>����[x���J���\�(g��V��ِ{��F�� .�-��U���(�Fin|L��|,���w�޸�`�N�Pz�[^ߓĿ�*)��3�v��4�\z�>f�wIlx@��2zF%����H��"@�]����������e��)紾��	y�3YY�{t��1mb�ގ����*5�J
.9t�R�-kR:&�ޕ��3�b��K~���um45u���|�<�z�4Y�]M/`�Ss����03�u�kt�+��n��*	n)�=u�V��Qd�6E�NG�޶�;~�q��l� ^���o7�����؃{�_������}�M�z]2�%@���Y>s��T|A�V������#���7�'K,ֿ*���枯@�Wީ��c��cN�b��vhk�9+�|�C�gk���Q{M������j;Y�z��[��/1t��q�"�C@E��O��z&|�k�3^NT��M��am�r���YQ1ť�}=T7�T�̏T���>��C'ڸ��y��p��7j���j0�����[X��ł92)�w{�ʦ���ޒ)����&�d�+����>r���L�ewDo�x^}�{E�nպY�ݡ�����t>��9b�8�x�����x\����n5�x�y�o��&n�s#�7 d9a�5ry0�2�&�Z������3�6uB㣚B����k[p��Fe/_(��[��}��Nskx�Y�;ٰ�TQ/���V�m��z}	r�M���W[�hY��te����9�q�ٻ]�,ǳ>9���m!���|�(Y����v|��1��{M��d�&���*��c���V
��"4����w)�}u��5�3V���i��B�s6��֡�#.�m�����5��9��KOȗ��4�5u�Bd�vUr����yJn8�
WTO�I5�+XKld�i�ΓX����w���kJ�qu�(ҹ8���.�m�+�$�	�u�Z��\���=��*vU�����r�����h��X�J�l���a�7s��P�l�[j�Tu8�t���wAYR���N������6�ܝz�h"�������f�\̫iI�x��/�ƚ]�Szᡱ�|�����9��'j��Yw\�4:��;�d���Ւ�'H�ض�&:�����qr�*�#���5͗Mfs+.��t�����A� BS�s�f��6Ԭ\rp}�C	u(^.���Lstk���0i����\e�K�j�>��:�(M栻ݓ�1Hj����+8v�͊�i�`�ԏu��.�@�NS�):�/�<`1=��#{ngo�6��L9g8s�;}��=���f���T�Yl�JZ�,]V�1|݉E�DM�
�	�I�"dwٶF�5n�E�ݙ ���a�a���J�v¾�Ȱ����������nl2�oz��9ݛ�;ޱ8U6�w�m��G���j����QVM<&K۷�Ǆ�aݣ9Wx�C@��w���Tog'�j�*�d�Ɂ���f]�$@]���Ԋ&�.��\|�YXze
�<�+_^+\opk$>���u��*
���6�"Z�R��T[k�)İ��YY3١Ʒf�p�Uo=�X���!C��]�����%���GۭYFu�ڽ�؟c���X��,1�*��\J2Q;��7��7V:�$�`i��.�Hw7�������;�)��˜�Y���À��u�#]*,�����jQ�J��ދ4�h��8���z=���Wc��zl�m���ƣ=��r��iڼ����tp14��1�ٔ�85�s<�xEu+�yC�qr��1)CU�ME����b����n>N:��β�K�v4�>Dm��ֹ��1A�=��W\�"�l�Ye>�|�-��jc��Mh7�"�|���=�#��^⌥��[1
f�����uǪ���:Tԕ��4�ב�t�U�k2r}H��1�*�X�5�Wh��S�rg���0]]�|����t2�+�C�KՆV��t�2�\j�\a=�H�S��;�LI�����cl�N�Ǣ]�pk#�"kW(cr�h,����_6"�ΦQ��*ꔸ�G��\2V��)�7�������9�O��A]j�0JcK���X���-T�`��tC3^�.>V�WX�B��uy���/��]\�/�;\s�+�����WS�7'Y���j�}K&�"D���6ʯ(1�ѠO�.N��:SB�(#��L�e�H�>@�a$g��^�dDv�J��A�H�IJ����| |���8��0�z����Q�B���UV��M�v��Ǐ�<x��׹꺫�A��蠭4D�AAW#����;Q4��qǏ;z��Ǐ^����<����i4�>;�L��Qd�O]e�%�d;z�ێ8�Ǐ�x��ǯ^�a٣UDj#Y�e�j�%���t��8�MI�#��A*�mӦ�q�<x��Ǐ=z�:�kP��$�P��D͔vY���]�nK8�c�㓓�.WKZ�����>g�P�Ղv�����|��,�H�.�ܛ�$�nv.�w[���x���sG_dI����N)$�Ri!���"N�Re˳R,���b�	�B�ECy��/ĕT�Ir��z��}����]D�BP �s��3������5��:(��Z�/� �"�D5 ��Ӏ�e�TP܈�)�S^q)�+�j�m�z`�F�w��i3c�H��`�uyLQ�h��-��`�C^0NG��Nyd�.��xj�H�<|�#�jcD�#
7� �������Hy��s�;�����|�w�k9��z���4&~�.��u��dM�rd뻴���G�p���Oc ���?N� ��B��F= r~��&��f��]wDu�Z��r,�����]gCjm]��D�*���i�g<�r���G�����	�V�́��`�T#���ڥ�c�e��7-k�b�������jT���6V@��b�xD��ܦ�˭��!jv�.�1�v�[�� 5������vS��a�g��S;R�W�:�<w݇c$#}Y���}Ut "�U�������E�Ճ95D�2�U
���(�޸I,�N�^5�I�&*:�;(�E�Ӫ��Mw9�6mx9�����>֯[���vY�J���MKÇ[�W��<���/�ʾ�q�F�q��w�����������M>�|�Up�����Hg��wI�c���[�3V�:�S����c;�|��⬬΋���#z����\x�[����O�V	�g͗oSq̗�-Җ0̬a���tU�V=��B�a3W%{W���SY\��ʡ/L�%�i�85ԞWĻz�XS��n���:n�e�;җ_wd�@��
�2���\��#c`��o7[�e>T5}~�J���5��(&;�7d�®�X�w@����������y�s�V��M*��G��dl�M�\g�p�ɞ�u*Ӭ�th,�Y}����}��pA�)�Q�~=S������Ԋ'����(�ؽ�y�B��މv�vg���	���b|ὡ3�8Õ D'v�`em��\�!k�|"�l������1��:�׏�~�h�Ȁ���&Y�>�yh�9S������-m� O5��. C��.4���,�z*g�Yv�b\��q����g]��p��Ц����#�cA���f_�Bx�zi�x
vy6�1Ǭ�9"��0���Էٍ�e��[(�o^�2.i<M^��ﳅ��5�|z(��R"=����Wy��2'�h
���bn]�_M�k�㱆!���5��V�k9`F����J��x�}R�&�2k�_)�57h���qG����O+���o�d����}���I��,O��jU�W7-�P�2��Ԧe����5Jww���b`�bcҺ�s�mv���9o[9()J�k���G5���[]��p �b�z���۬�/y�tk�a�G�*��]�h͙���|��kwƟ�c����6U_q�Uj����^� u�����%^G�}�Z��>׈���ȯ�ϗ�yh��b���l�{��֐1�*���kf�M,�ܰ����p�t�S����}?d�-x9]����Q�W>z���U���[ߚ�2_O�b�����w�g��m���nM%����[���jʑ�ԿG��u��g���u�a���H�M�Z(�/�0��9�[�O��yW*[�fJ$gs
���8��~��߽>���ŷ��,%?P��OBif�M�R0U<N^���b�@vq>Rr��>�״@e��zg�BgI*&9�uvN��rg�=�χ�yu��Erj�q�$L���v�>>���/;?�x>�Ku:�8�(���;M�~[������%��2�0a���t����69Q�ʔ�q��zA�{�aձ��m�f_������s��g�S�M��Y�6����>�[�u,][����%%v��r���X�	�$����7����xv�h8��DaC{���ː�1���:j��2�jmM�&`4��W�ԄuI�j� V�H�n\w'e���gO����{�yyy/////  ����_��ɏ�!kǊ][3��>b��-�}o���+�ת�By�6�����.b���{s;+���-��0ZzT<W*$�WQĽ?mU����U$��<"���X���,@���n�2�(�77�G����趣K �9Z��e/Pɏ���b�-�S��㥬Ϟ�U�߳&�ޤc�[}��Lk��qyF�z��d�r���޽��Wb눜�M'�5�h��4�����a�	Y�5�Y7�W<����f���@�El�i��H��bp�N��tt��U[.����#Q���[e_�:ǎ�m^ފ�n�b�����wm�3fҟR}��s��#F��k!o{8�id�����ȷ�p,D�-�S]wkw �VW��Gw^ ���َ���{|�RM���X[�#n�^Q��/�1y�s���ѫ�Aѹs��A>O��.\Y�G<ʙ$�y�%��Jt�2�+�Ĥ���L�t-)7o�=mgkM���"��S�1��wN�y��ӟfwR���M��%�o��E�������^�T6vZhW�˦�V}�5�t�=��+KT�n��w�1�y�M�.p�G&����tM]�jk\_�1��o�\��YSׯӊgF��;/n���>��������g�ԕ���'��B�}��6�Y�y/��=Bv�*��ö�� �^���3#��/����� ��ș�PE��ce��4�+��o7�������h�99|1�Uֿi��|�2r���fj\�7�:�kMߩ ���Hl0�WH��Ѧ�}�m�y���O��ޤ��#Y�Z��6@n���y�8d^#/����Ÿ���-rA��S���z�G���	�$*ދ��|��ax�Y`P��]v��{�^o}�<�F}�紅>�\=�	X����mL�(�m5;�� ��#z�s�DIWB�@�{'̙�i�rm��v�M7w���PE8�u�bF,��F:��43o"�R��"&v
�n,q1�Ꞡڪ�c��H��v��;Z:���]���<�^����Uu{MsGd���a�׎���m:*i��9ŗ}��*���(}s�O�p �����Ʃ�k�f�O\�E[s����ٙ�F{z�r�sɒ����ͣ���Np��e:����U2�>~ԕ��N���/�+�@����!�����#9����������蟶�ۨ�����)��1��]���~W(��[���om��N͊�z��ݼ���]kO&ZⲂ�������=�r��U�Y��г� �E�3z��0`̙QΟ�Za^o��n�5o=R7�^�[#"���e^Nu'�3� xmf�|�[��F�B�Y|��P����j(��ɱxs7��k��B]��bS8b݆d�����ǕGq�����Yó���y�:o��fS�DÐ�uOlzљ���B����^������ͬ�<�/Agni_"�+�B�7�I����v=��1�DB�LZ�+�J��=��p�u�]oٹn[y���0���ʏ^�7x���q��.�EN>��^4v)=nd�8ݔ���<�>��`;�dil,,$�F2���"^�t���y�
Ԇ�QW�*�6oN�ؐ�d4V�9���o�9���\j��#�~�;򵥹J�%}�H��k|��U&���Fu��9+9w��裨�ۂmf��f��ƝrЃ:�0Mw9�|l������S4���ӵN�;h�-:FX�1����B�z(�gҮ�D�	\���ߓ<���=~1�c�ܭ�2����������;�]��|pi�7ZD.���=�'��t���[�JJ.r0;�-@lɔґx�V/^��J�fk�7=�|l��[Y˽}^w[����:��[���fQ_A����o�������!�cf�����t�3�~�w �B��w���/�2�`�S�yR��t���ӱ�����'7+&�z��c�1I!n^a@� ��	���k��~�{ܷx���<	�7��ȝ��U���Y;:FMFa�x7��K"�Ǥ�xgw������*��W{6%N�����w\��z&�u��Y�K�VH�>7Y;5F�0� �]�g�V���� �
���R�����yY�p��1j��V�Ө��:���SG*2�N�g�M�[����E�8�Tov�����I7�\g.l��x�Y���/��h	�]��zc`R�g�Ѣ;+��r)�M����M�����4w�i���O�RReɫ�oL�k��̻+�HB�
����,��=��,���.�q<�*Ш2����+0T��W�sR�
�ggvd��A,uw���k^��U���i5�����y���*�'l�n����Ȕې�4Ujk��=�0+�.�8�r:����i���z=��'��Bl�mC^� �P;�͹A���<4T���m�m�+xR��I���ȅ?v�����5�eS��O�~����I���s|��N�P�3���7ىW�w�����#�.ze��y8�&��}���!�0fˌ	�WXȪ��1v�j�6i�γݴvb�����+�`Ϻ��P[G��w"x��M�Q��,��#m^�~��AUSNw�Ύo{X�`��U�[�:T�~ቘ/F�Z�ï<�;Xz�57Yܽ�K��<�ǂs�s���}/zÕ��5��b�DT�#zc!Y�Ӻ�P��$�ӑ�]��s���.���K�bR["�'�nR猹��{��|-?{9��~��^�HYPe�+�_���-/g-���?LA���	ݰ�(H��§ ���ֳ�S�)���{n�g�'�fu�ፗ�=�z�O�gt��\:r�V**� Ͻ��bo9K���*�B�O��Z���V�^g֏�4�t��e�o��[L9\�Ÿe#Gw���I{]ec�@��bd0�*���������ǲ��o�ɯps��+7k4��ڨA��-_�y�4+{"C��D�Fbފ	e�0�1��F�<>�g<��.J�{�O{�c�$ِ���L�f�Uw�,���hy�q���:m��/N��Hr�;�m��U؎�SB6�Z\B��6T.���f��A��r�4gK F��<���Kݱ��7~���30ZXȣ��c��]Wx����0*9P���P����
�b��ĚN��_��s�يd{�'�IF��zwzk�z�Cj���]'3������?wyV�ne��'�~�3�Zb�{!�y:]�m��bG�~��vz�;	�m*�m�m�v���"�L�1�����89�]B���-o���������7ݓ�Y�xK`��\
�r���@���p8��ǽ}0
�C=h�J��M�m7�/8qڸ���l���-C)�E�M����88#�}���q��%5cu�+^�[�H��^����0s�ל�l�P����)4��g��;l�nH�ͭ��>�%�| #���ս�l��}�tGosiD�
]r6�U���}|%������;kF���xq�I��{p!�T+�x����������$�ָ��	��Uϖ�$��I��U᩵O�7{e FnD��{���=��e�X`�{[0V֫,�H��3u�z�|��m�$*�R���5=�Ow?KV2����Q3IT^��E�sQ�l��.�;F�tA��|;�.E��K-���Dۙ�#]CL���I�I=77-]f�5�g.㉳w�.�T��l��O�Wz�ȇ�,�L�r���nϛk]��\\�^�)k``�z��SQulh\
XT�{�Vi�X�=�g0ݼ��l�g��ʧB�T���1W�8��j���k�zn�����m?=U^d�dĥI�aA�퐸�Z3���G���-(�o*���8_U�o^����x������J�P�V{�t�Et{�@�\qE�y�L �ՙU���I�3��m��`L��C�t��=��^���yޯ��'��y�y ��K"��ʮ������el����Uͥc���B�xl����֏`غ�g�荫���R�G�lI���ZY{�LU��߀=����`a�ɻǯ��4�!-���L���]�ʜﯪL�D�bj�S*��].�\j1&��BMŕF��ϥ>�z��OP��`=$1�-1�lXn��v�=}�sw_k(}���7_L�wMR�����Kc��
ۗ���ѷ@�=��Ey+H�9kzԥ�A�T�Z���M��ڶrZ�Q��+�RS�&ޮ�9�����5�l��\�	u|ʭd�Dݎ{"YJc�¸,�I�oeWׂ�	�r��񊤓e��
P�󅋌[챔/ik���Ϻ!�wT��C�uw]dl}��MB����dJ�jd�&���O�q��{M�L4�p�k������h��vbܙUJ��s��(�s@�o�d8Jǻ�Baᮓ����Q�z�ܹr�`a��]�K���FV׷�h5{J%�d���Y�мGiY\���{��V�x$�RJ��!Ğ	Rͳ�����:41�4K�K?UC"{E��J�V��NFj�3n�fuo@�D��@�ԍ�Ɯ#��]�t�c4��xZ�;e��'c�k�Ë5��v�R4l��)a�U�y7���xX��<O*�u�BW:b�p{r�y�Kn_�o����61��Kk%Sp�m$�r�Js9f��4�Rcz��[/Y�tls���z�z�*º(��֨f�9&��峝S��.�U솸δ�N޻Z>[(��'��GXӛwFvY�f�So+�-mD��&[���D�
�2�[�'P�M�v���o�Ԙy��.Z�ʛ�<�u2&��8h�:,ˌ_�v���9J�ū�=�ۂ7�8.XΤ(�E_s�8fov�} ��� �!���ط��Nck���E�(��|$YәX�ka�t�l��,s&��蹾�Os;��%��0n���"�UH���	]d�5������\e��N�+�!��fŰя�D���l��bg�u���V_V3Vr�km��|��� ��Z�e3�o�m������K��-�	���A���w��9�_�Z���
�I���V�+��^[���<\Q�<r#[�Z<�	Z��#��D�rc��W0�Kd��J�o�t�ǟ��.�;=��\N!ԍ�F�
\
���a.q�%垜F�Jr��fX�eJ7W��\ۭ�W�ffw7��oy�m�Ќ��A�`e�<-Թ���ü�
�Ղ64��-Ύ�!N�s�yԘ荶;��
���h��r���:�_&�H�R�Xֺ�5�]�4��&��CQ��n.�S�aaw���`��s�TT[����CS�7-�'%fs_:��X�iV��=��.BHw��
?C� �A ������W�L���F��]t���C16wo���o<x�����Ǐ^�XN��$*R�	�WC�<�#�WiT���DHU��|�o{���������Ǐ=z�!!:¥wZ���Jh�V�J���#�:-L[��(�
$�@�4���q�<x���ߛ�~o��|��l"�-��QC���k �IQ��׭��<x�㷯<z�:�
�sT+0�L�Nme4W3K��VԄ��Ljh��Г8EE(m9Qo��Yr�F�.��j�x��"�QH����x�p�0�-�^m�z��I�LR �Ki�!_W�?V���EQ�TO�9T<I�EO ��s�
�a%K���IgTU(��2%͎k@��"((��8K�u�q+鷔���s�.�Dy�Tr���'��~x���~��^�0fr�I;]bq��C�_F��i�kR�ب�t��.�}�^r����y72�z�1�c��k/��W���9�O���5�����s:��
�]SR����c!g(������07�;�����r��|�EQ�����YUz�1��xm���gny_��L�q�ڑˇ��_��g�a̱���zʐ�7M�b��>c�>k��m�ٻ�#u,d4k�������Zv�2�z9��݂d�o��Ӝ�X�ɰ���ց�]E�c�ikK���;;���k�x�j)�Yf���Tե��4 N@n���Y�^�KQ�je��zݖ��5�z���	T���c4������~ͥ�p��-�� ��PX\>��-�ͪl:����R�4�I�6j:g�'p_0p����0��
�X���j�[��3a��g�d����V�\�ݨ=�5}>z���#%QɾSK ���=Ot�%��r�g�2�G�b���V��n,e^ˮ��h��_O��|%�o�]「9����>�J�u�[.����*�� �J�{��ͩy�pa=wC�K�i�Lk�q�5��ןGH�`��
��y� W]�(�\|Ly��ի���%���@�߾?7����d����̨N�M��V_�G���*V�56P�9S{�_Of朞�4����	G���Z����Ih9�ШÕ��M!^���=���d�]�^�N\L�ѽo��,�G�s+����Ǚ}0�j������v�x�K�۱�{uOh:�'��z���/e�������o:�"4V�C4��m��o7��M��x��W����9��7}At8�Nr���1k���ڢ7 ^xa�~��G�Vy�E�<v	�y~��[n��prM�3�����}�����k���_����ߋ�mtT����>��s�K���������ݤG��K� '�%��ًX���3��>۷��_���"���,-��tO�Ir�X��c2��}���Jm�2�:�{�3;M-@]Ё�J[���6x�|�����^�:85�\���c�Mގ[��NB?j��F����m{�i��rnw�~��b�����������+jL��m-c�����*��y(��\��L�X��<\uW�+���Q{�|u�O��]t��8mw��Lż��s�!8]Y
�Za��SR}�������������5y�:�s��R���bռ���Z�dn �s�o��~�tZT�`�e>�<��>��ĽOf��8�\�U��R�э܌@�(,b�-�S�����>p+j��l]���aΧ��{1����H~Uqە.
�T�#_�"�'}�
W�������;渙'��&�M]�nCtT�e�^�%��+]q<���eQ���)_��ol�h�#1���xm�i���G���VL�k�dx��͇��s³o����OQ�:3����n�Y�kn��
��Ag���D�v�SWg��o]�fsv[$�{�N��O5�U�[�����Gup�W��;��7�.%L�[�;f�i�S��&����ͷ�b�`"��Vo����~x���29.���X.O���뢀������R
�'�PB#׶���n�Q���ʷl��y�a��aI�'�<�"����p�o���𓮓��:rS���zθ�r�5��7��4cC!4�ʇ?O�f�WO�n?��%�r��@�V����m��e1Ŭ���ߛM��u�kZ�Wd�������A-���N\���vf��n�v���}�������2����F�E��m��3bdE�42T�Di�*���rz�	�9ѥ�m��k��Y]���w�@vl6���R����R����W���4�0;��&u�3�v���6��گD|�m�0�q�ȼz2�`KwnmOv��'~��m���,�q�FL�ܩ�;h�#۾���m��A3a�4��\�_Rx��ӓꊇ��;��0�n��BzE�gE���3�.��猞U�ݢHj�}ݑJ�_HW�_~9������^�a����F#��ve�槥��C�Q �����|�~�gcʕ�3c����6M���TΘ�7�z{��~�R,���Q_g�>#��}5 )�S��L���5s�4��o�Vy�N����Usf�e�g�Sfuca�Fk\]dCY��0Ӌ4�w�xӏ��fym+�[Y!]\�lc3ȶ[Ƶ���TX�;����O+X�ۢ^�ƻ�ss�������I��b��!�-��f�U��Vr�oJ�2ƴo��{�OO{�.)]���κS3�90����扫��ֲVaX��ɷڊNk��ީ/�I�z��3'�[��c�1�k>����o�@���5#�^׎;f~;+d+7�#�Qc�����u�����f��w�L	�	Q,{9)�x�yo,��nQ6�l�=!mv��D��K�ٰ�L~I� �QHǫ��w�8�ظ�',慹݉g��FJ�ڍ�\5�f{��Y��u�n#9r��i����^�b���n3Xvp���~'l��Q�BvH�l�h���6�����;���).�b&v�:�9h<�DC�\w�=���Z</�®�J�q�mB*�8��;�'w#[j��x�w���@k�/��k�w��rBs��V����߷�Ź�q�
��WNY`6U�����$hϘ�e�rz�l�;��n�3t�2/R�NB�b� ��{ ��z�Kv��2~�*�+?���LL��:`3�3�u+�l��U3�Z[�k$�*�x��)���x�OѦ��U[��[��2�ګX;o�>�-����A9�tvYÕ<�_I���5�A�0�o*��kwm�t�nK/K��.�F�[O�����7y���[��n�8j��U\$~0c�9��o�n*8O��N��:���ᧉ�SOj�Gt�Q5]Wt�c�e�#�8��5MA]O�N�e���Ǭ?+��9���ɫ�eQE�U�gmy�0vbռ�m��W���J���[a������w8T\l��޵��U�Z�kz�	���h�f䪲U\j_�
�u�^y6Xӽy��|�8���-�'!#���+7��4��Uj�s�*���uŞݼv��q���X|d^���j]��z�N��`�
�NܖF3�vb�I+��RX�x�P%�Ȏ���i�K��ny�n��4o:���(Ӌ��;�Y}G����_B}�#󞀚��k�$΋3{�w����z�[�iZ�P֬'Rr56ǷC��j���c\]Ѥw+�nU�Dw-��덫�� �E^2��=W$E
>l����w�ޡ�e5���Δ%�.�3	�N�Rvu��]%�!&��I=�7�����|%n�ԩ� y2�o�����F�&��"�2<[�Q���P�u��0�µ���E9�.�'�����C����Z;��5J��4�6�w#��oz�-�a�I!��|||||}kg��O'��<����*��a[2-��~7��V�泳�7�.VM�x�Y>q��5}�Q��g��k�}�kZ��R����an5O�	�@X[׾ùi�n^O}�s�}߲����paz�/���2U�ϳ�əWX�%W�a��=X�gW?u�>���A{p��-bTA�W��e� a^�/){N���kw�k-\y�n���d�w��Vy+vFY_����!���ڶ��Դ �w�z4���U&ҟd����ym/CH�{��ao��Eer�}x��̂L��2�U	hC�
&(��'!"�,i�O�y�ʃT	��7=��m2�k{̣��M�{d[��mT��k����F�4nS0�f%��@q��`�j��^*|/��Y��[�pb��۫˭�+k���ޣ�r���y�:wp�>�:�d��/��0x����q�PD�����RTO7��jGi��ri��������X�{�0�.=4\Ø���r�P>6��I�#+��¨8��f��G�2��yMdNV2��=��9t�=�T�0���S̍��N�AF*�`��WR������|>ou��36v�F�.u^��8^����;7 F҉���l���fnO#;u�$�z`�H�Ef�
5�(���K�!�ܤq���NiaA�9��UH��'��\��Αq�(��Pnޚ�J���{"��̤R�ǒ⚚b4w�Mj���ڟc��21~;^
��3�Xf}�VU��
��nR��YtX�2X�v��BC}�|��;���F�J���\@�ˀ�;s����M�:������a�=5�ihmL�R̸�Mw���g�ϳ�k����s!���cw�T�`7w��q�ȼF_�����骿f����#��ɬl��h�l��mM�yw-i���|����n�=)��fqT�[�!o ����<}N������5RW�۽�Z�	���֍����-�Yict͌&]����T�!�W�CS�Y�~�~6�_N^{tryv`|�CPM�ӻ8{re٣L�ez�R���y��N�ش�^��;\���U������Ŋg��fS"���0���_Qj�]\{�_1���xұ�7���=��M�x�|}����{���<��&z�.̺��F�φ2��AL��(���*]����3�Kf���|?]�M�oWU��}��j3�NO��*/�j�td�Gvm�r������:����b���D�v��N㩼dd5�m[w��S:�����Zc}��e�����W�u�Q���[zk�=h�c>�چՖvE�k�C�ͻ��Ep}�M>G`k�*��[؏�Ȋ�ٞ��Q��>�B�Y꒧{L�y!��ܾ�⺬�r]�Gz��o�We�6W+c\p�k���꾪H�x��b!��+ӫz��ߝ���k'����`cU��ս����h����~^և�h�`��Y�7�=��F[ݥ�훊��\���;����ŜL{�!['����[K-3�j�,O��Ǐ�����=�L�@P��Wj�2ѽ���F������~,��o~�ί��[o(��j�gjBa��q��k4��$�uo����+r�_�^�����^c���/��E�*Z��}�!᧽��P&(�|:a���ͽU0�7P�T��q�/bo��v1�y}�ؠ���@~F򎸓��zԡ�r��e���75|6C���1�j���q����W;�v���3|y�=N�fh>h�4�uݱ�Go$nU+��=�i�	��#�T��K��Gt!�A9#�u0�ǶGJi��r�kN��a��؀��y��\�C��`�{�v/���1�Ki��Ë�V��d��V���Ԟ�>5Rï���}��H���=y�ﶤ>Ϳ.��c̣q�p��n^���/j[.սN{���e�S4M~�4�nukf�b���S����y��f�����U��N."vX-wcD���#��������VU�X���M��2�f�YٖWG���AuR-~�{�~Xul���z^�X��-�����W.�������ܒ�}��c ��-4VY_Ok���i�A~���7��Ȝ��ѩ���w :9|
��G�s�[iR��k�Cޣ�y|�L{�>]�J�j�0i��["�].�d֨��4j\���8��h�/�^.t��tr�J�jmW@믄]�W�}e3�2����.b�2���J�-Nx�H~��6�o{��,d�C5��T�V�-�"����+X	e�����\�	!فU���9��Y�y��w��u��>Cz�.���sж�
��
V��I�2�H��eJ�m(��L������0M"�A�.ǹH\�|�:�e*���x 4=�2��k�+���@���K�͎��[��v�WΗ �.�s�5+j��uh:�@�#�"���a0͎�=!d�N�� �Dg�+���je��J��}N��c2\�仼)��	f�S�g��]ώ<�r�ReG��V/���'���V��z�U�u6�V�,���l5���-�M�+���7.l�� =���,|:���F%ť ��q���*KAZ�2�6]�WM;3E]��OF�ر)2��iW�r+{�wY��5[�z���J����d��I�y��Y�޺ҬIҊn�m�1�՗},�2���<��*n@&�x&�����dCg7xrCY˺��P�L��3a��$&Cil<1
��48n�z�;
O�Uz��̱p�rAN���7�6��>��o&�.���#T�V$�IXj�w�䱯4h�`��O�[���P{�\�����ٻyݦ��:&�s��Vv�q&I~\��*���(�U�&UF&�v]��6�m�jS�V1n��,�wKLb�ш����,��y�|ߧ�3=��Ӵs�\�y�V�;:Λ��i"�9�[v���,bP,�<���p�A�\Ԟom"mܮ�49�"6�S�hij��{F7Z�a����Zb���ەá�.�`�|���pSr�y�F��iZ{��Vg�k�S�VC�n=%�+�ެA�\���i�1gfqc��dիǒ�3����ͥ��5��M#�j��-��������c���]��qT�Ӹygɧs3"yx���ͩ�$�Ix��DP�wM�}�"�EZD{�[0d��0+Jb���
�+Y�(8w�#9Y�y��盄p ��_׫'�K��q��Z��!�P��dI�-X
Ȟ�K�q���L���J����2>ZVm��F*ci�Z��C6єP#%<$�;�[��:R�]}i��u�Tq�	��2�,ًU��/t�BUY���*��i}���Z�S]vQw�˫���rh�H�pr���n��d�R��v��_m��ܢ�7,���]u��|�37�y�Ν�+Q*��׉���F�=��f�yô�U&�T�hWhJ
QY��ǎ��v6���w`Ht�H�]�W>̕&��xR/�Z��
�"�U�0:�v��v��g�1mx��&�y��Ѯ�&HB���@�,�ڂ�3�vFZ5)<�/���xz^����O�<N�"���"��I)��F&�T�d%�Tۧ���;v�۷������L:�;MH*A>w=tU�2�Qg��B��d��[�]Gtt�:ݾo���q۷nݽv�ǯ^�>M2��
!�E+�J�><�"�G.�I\(.d-�<�Q*u�|�>>��۷n޻v���쑓�	�jj��#��I��t�9r.r�>!�W*5
��I�[��|q۷nݻz��ׯC��5
��|DO:U�:*DfI�f���hp� �(�N(Jh���(���ΜJ�0�}w/dURX����Q����.�!9**"�.X����tp����[i�*�TJ)�T��:J�&EĪ��+��I0��Y�Bh�2��r����8d����33RbB��dU\��Xd��QRh�2P؆�"�b)�W**���T�V�9Q�L,ʲ�*�I��)i!�>�={x�A�E"c�Nʁ�A�a/ �L��4�r����|��6�t�p�&rK0�ֵb��`)�$j
δ\"؆�|�=w��-�z���"v������I6X�PE�J5
a!Bʐ�c$,L-9�8#��%yH�&(�$�8�9��>>>>>>/��g�}���X�� ӷK/Sm�N�g���տ��;�WiJ�Ab8�4e�-�G7�i�e�}B�+Md�
����n(Y�/^K���y�U���|�x�D��eA���3�#�ss�/Rt�Yܨ����rc ϴUa��ϼ���.�k��"[�UL�gEJ�Mqj�q��滭za{�6|x�zg�3��f�0f�ap��jT$��ʀ�r[��p��gq��rb	���m�m�O5w,ӷ�{#}
���ݝ>�&`,3���_4�VY6M��{~]9�g	� ��i����Y�C��%w�l�槽;�[m+;Y���{��#Q�mk�5o��c#��Η�K� ���^kVCv��f��p���)d]��׋B�s*�%n�M2���6>���Xǘɚ|;��Jm䈛�W_J��`][G�r���U��0�Ǩ�B��Xp��۵^1y鬠L�g{��޻�i͜ctMSJ|�TC<�)�b���/vך��E
ו�ڹ���A��ˣe��Xa��+7#�hԝ������}��˾�� Z�3fͺ43��tQ�9f�T
��>>?���H���xuO�5C|{��a�NF�9��s�Ж�<n��n�۪��׻6s)�=����ِT12��l�?{B���/�mV�Mq���%U��Ϊ��QQQ���t��������_�����N=v�TugͲz�d�{�w4r�ܭ�r��v���
�!n`5z�y��V����T3t=ׁ"x�Uyj�Z��V�_T�	��ǀ���+�uO�%Ɏ|�5����&�9"�hj3eos��-��F���c�ӅZ�D؆f ;x3,�ܼ="x��e�6�~�/�:))�[��֑D�>�J�xw4�q�vf����L�����d��u���ŧ*�Y�!�u��뺹Z���|''����h��**a���O9�0LGz#�xM�f�6��T�=/���~�aas�Š`L��=tw�b���*�����+3�Uǝ��`ɸ���T�M�]N����yo���Ny�
�b�3	rK�}��0�5a�j.��x�({1XL3������y[�(�+IŲ����2���F$��u%\�vM�FG�og
��^ƛ�-ɛ��%�Lܤ��9\�����~�����}�t��y��R�4d�;�o}�ễq�"筣�ИL;eR��]�;RD蠽}6j=��C^�4��Kr�T��֧�漮��rb�v�x֞/N0(5oM���i��Д�Uh�N��E�l�;���jg48b�X�]>�����Bx��ã�|[�j;'�PA^�z[�;���;�h�;�;�nȚb�i����f�:`L�y.�&6�R���M2�|n*��?x�o�4���5W൱�z[��Uh���	i�O�ۜ��Ɠ�Y���ӏ�<���%,���]W�۫�]�wj}{\z��et�w)��1��Gm�l;K�Z�9	eqҊ]X¢�ܫbj�K[.�Z�;�����g�CΦ(�k�-0�8�� �憝����Ցl��=�]�ET�H{�GZ�n�WE��G���%XA�X���oL��v�#g�e*ٖ��K�Yr��V��<e���u�l��+�S�0m�3o��1}�腓�K+��2��}���8�Sݻ�]�gf7E�ʥײ�w�!�p��ߥ>�1�y�ؔ������.�d��\�$���>>>>>>s5��؋'k@�o-?7`m��v�E:�ם���# U�/"n���2j��F��q/e�rO�;�N�:��e���������Ä���A�����d�2�аR�������$�=���;��ł��Y6m�l��,�
�z���˭��ܪ�荀5H�VW��\�"_y��O��G�k�B����G0�l�;�r��j�@��&]������dk�K��tN��=�7E�D㦻A�s0oy�˅f��=�o������Ǡ����N*�~��A=��9�7@�R7���v/Ҵ�f+��Wm�7��>���Fު쓳gi�@=�����gmݐc�T՚�.9��a��3v�OM��JڟiC�����.5�T����ܐ�˽Op�~g�ޑ��;�f�U�bj�{���^�1��
c�����˭�mDSO�l��~��Y���&����,+�k�:k}���۬���k��C�GC��Ƀ���z�P2_=R�:������;�!kxVW���ժU���N7K�V+\�k��W^љ�RuVH�w[��܎��޼�V�w�ٮ̮sz�IQ�ƽ����������,{T�����e,��);�,�tќ6�:�m�*� .�m��J���SqJ�ޡ뢺"@q7��&q-��ãp��`2��
��+&�#G{��0��f�Ȭ���[�s���N�dBB���5���:�Aj�V@��l��׎I�[!LZ�Lp��=]wg���zszi�E�
�K���ڀ/��@v8Lx��mÄ(�<�"��k��mX+�RW��e���]��m���vf:��uQ�;4F������+���%Z�p����7��ݒj�����s�jx�]'~�SEꩂ͹���X�)��jv^#�B�V���z:ސCgC�zC�S3�羙³�V���0@<�S�i͘������&k�SC��?�� 5��Mp��<��G�0Ilo�d����j��=~̮�����&��;5\&(v1�� 5��T�{,0�dx�H?�Y�6���h�=o��}�@�2cq��VT_]�Ǝ�1�7έiW�0�Lvڂ��r��y|��9v���8# �����d�ڛ����w��r��z�{�z�c�wbz�W|$��|�*��詐I�vv�d������{��g_-巚�{�0[|g^��3�H�<�8c[f\c��2�~%�iSJۥnҵ���	��Ł�,���Q<�-*2�,t�c2<���g��tĈv�5����a�^{��(l���~�.!H���j�h%z�����j�wU�&���ww5֟��NET�Q�9��Ťy�[K�̌�8O�K	����j?ٹ�⳩/}�_Zk��n��t��J�5doN��%Tr�w��וt��O��}unS<jc�����U�>�"����,5�j��t읢�x�Ѵ|johv*Ī�<U�U���G�i������5�*���{7f��s������g�|No\�7Kk܀���>��aY��z8b�&%�(���'�m;Dz�U��둿�l��*����)���=3͝7n�mQ�k�&�݁�(P{�;9w�oWy-�i�ܟ$ml��Ӻ۹��I����Z5QJ���ͺ�{*��[ߡ-չ6�X���m�D�!�{U%�+nіX�F��>��t�{�=k�~sq�1��:�ٻM��*i�5�mĦ� ճ��s͐h����J�'�Q�}v�;6��#�����������n=�g3�&�o�40\m�=IL���\�%n�ټ���ma���f�6zl����X��,5���}�1#^��E^���~��Z��Ө�+}5]:��ܮT�=|''�M�����(3hp�����Sɥ�����\I1�<��$_���9��z|*t�x�0X{>�r�8���}���V��m�+�%�ix�D�dn�oiʂa����{!�nt��v�T�:�h���>��@=u"ἐ��xЄz�yS�4CwOv��k��Zm�j�=��A.�=鵷G͞��g����	-A3��mn�z����ަ�fK\����,����������,�����F)**��f$�q��F�U�#qM׷�ؙjfC�M=ɑRæ�j�f���Ɏ�M������5ޛ�n�����~��~<�һ2��� �_��Њɜ��m�dUݹ)�9mNkY`��r�����İ9�<���"����]���z��'���O8VZ�m��5-��+h���h����Y��ޔ��sk\�g{j��䥷W.A�+3ed�!O�1�c<�ʿ{��/�ܻ@k��%�]��,̔���ޕ�\.�+���a��z��M]�|*A�p�~�1#_��k��T�hWW:���s��S�)�!��\�c3�e���Z�<?���5%۬��L���(����q	,��y�ۛ�4^r�S�G$>��z%�䷧�}�t�����Y;vh�M�WwRPS��;���:�ս���o��F�NFJg�z<�.�o���,D����$�>`�Y�����A]�p�73�j�U�V�*l^%+�e�2��F/��a��_5-f�,յz�uV�Z�@�Ո��O5Ϩ;�c�Ѡ}�N��s�p6����Wq޹=ۧ��{^Cq����	d[���o�@'[�ޮ��q�ujﷳ��6��ɸ���}�"������=���㌎^/; ����o��Σr�V�p�u��SHY��ٰ����e9HZ}4e�IW�sZ�T]�T˻z5���Bf/�I	�ȝ�u�s���oq�\����R�����[҇��Ҡ{��N,G��MdYsr��n�C{I�����S~)W���|>P�U�g!�e_�?-̖��=�ie���+/i+�����'�>��{Y���͝�z���,/eTy��	���*�����������X�5�I����{��(g;A��Gs�7��Lݒ�TyH�g/r����ϴ�?-}�7x�sT�>y�oS��/>�:���z;OY�և��0��î3�u�V"�]��x�'=sԻ=f����-K�N�ӶK���䕼bl�eC���)�Z:�.;��ڟ��*sk7"��������oC9��*���ez
��o����2	��QQOA�is��u��uUQ7V����"�f��Ò�ϳ�����N'�~�xg�����=;tw{�"�����S4t�ȣr*D�d�Ճ�T3�z�T���;m��մ��f�@[���O���d� z�X�/��Ǯz"-���n�S�4��`<�*�F�v��T6;۔!+���i�^�Z��r5
�r�ˮ�ٴ@�n V�8XB������optp_�8�{���έ/�&�7Jy�|�k �R^�3�b��O���wf���|�*a#j�����.v7���;�U�>O7���%8Ӊ�:��
,��F1�cÝ�fw~����s�k��1�F!�混���{��{�+C�،C"��7"#U��`&�2��,c�ߒ@L�a��a]�;YD���AR�U��z3V���9bc�~m�i�sHI��>ّ\e\  �����t/���k�rk�S����e	݊2�ý��ݑ�E�×i<MC5��8��N2�^��g:���^G���8�E���wU��3]j��m/�ڲ�h�u�����V���P��u�7�̻Y׌���!�>!�h�w���{�l¦�N���_J�T�O�v��{�\B�w2���`�d�r��C�z�tu�䭂���K�$���~��^AH�>�[0�7"�N�\\O���3�������� �w�6Ż���UE�t'MD���q�� v��r��f���i�{-yi�H{�j�erb�G�{GNN݆�s������檣��i���4�	�Զ���dOs6�a�G/����kt\�뫝����G��{�'��s���bF�&:��XY�V�̦�8���PU�m��G��W��.��я^���
:��4���%Gy��d�/}��vW+�@QL<��Z���k���gk��z4�:��e=Cg/{n��:*�/$���U*�e��խ\��;����=̮1^�Y��P�f�	�j��>�3�S���zh��9_۱7����\�yo�R�j�ͪ�D��&Nj\���$Imfn;;8�ӻ��as���t��xc�,��P�\���p�ĵ�7mIP�>�FDt��mrp�f�e�2!����cVo&�����P-k�)��>�Fr�tE�u,������:��'Z!m^ܸ���U.[�MT����ZU��G0�¾h�9�0��U

��|rL�����چ	���хNՠ�]�:z�5��K{
�egj���j�\Gqi�\��|�����un�yH���;0#��ݦ3e�]�WH�r�d���hGj]�A^<�E��Q�T)I�1��WtcLTYqWa����VG��庻Z�36A��؎'��8�뽛�=�E����֋���r�z��Z��O�F�yyMޭ��r���#�Qug)y_DU�W��˼(�*����s�=�՚~��d=E��[\G�8J/D���/BM��#$��S��x�,�H_�,n�:��܈���D](a=�Yt:��ĨTu���M罏ݘ��S�(���bX���Մf�눡X�*�{m���C����#�*���J�9�P���I�)�Y9��=ϯ.�C���Z�:�1*/u՛�$�7Q��,
:�x��Fffڶ�u�n�N;��]"[S&^0e�.}�V"Y�h6+�,��n�jTàc=�pTC���jM��R��kT`�H���K$�륳�RJ�k�o��_[��Ոt%�ұ�VQ��^5w̻��<ނX[�g{��K�rf�Ď���5Ӭr��e�O�h�Wg�qOM9H)g�[�;�ю�j��n�ENi�ѵ;�����Œ��L��zWiJ�_^m��yp�)�0-��[ܳkI�Y��eL�$D���[fn¯V��'��&�Af<f*|�lt���vAl7�1��{�a_L_P�q y�����`�q�4j�q�W��$�3��rixS6Y��w�L����ԙ���Q�	��W+����Y�N�����v�㮝,�Ds�6v�4�6��9�>��fb��p��;��ԱiB��S�mG��eʏV�xܗw֥^8v��q޸��e�{Wq3r��2wS��a�����'iV��|HY�������ӗ�W>�3;xl�JT�Dٕә�pWW�$�s�fLԛ�������}/�
��ܼ"2Ҡ)P�(���Ibʹ�aEDM9+P�,�K$��0�)�ݾ>�v�۷o�ӷ�r��ʪ�0J�rL�BI���$��DE̴�2���0-B�PPA�V�,�|m���nݻv���o^��2I��B�#�%*:��-B��'*�rÉ
*I.*Y���"��v��o��{v�۷n޻z��a'J�%S!(��C(��Ĩ���!g"���
�'8!6!�jaUP�#O^�z��nݻv�ۏ^�D��.Q"Q�QTQUZ'��9�_(L�R"�������$�Z,h��U29r4H�PD\��]H���,�5���V��r�����aI\��%CK�3�$$��,�Ej�"�0��(T���D
(s2TH��6V�aDh�YT\�T˗+�%�rW*�&������04Bg9UE4�S����3��UUǨ�ǌ8QO(�\��U˕:�C9UT$
)�Ć@GΝ��4�R�m��X��"6�ZW,iL3r+㑄���Ӣ��)�ec)X.��:vM�SWi�ڶ�A��坴]�*�'�V����x���[�[-���3�kv5�x1���;�uHmY���6�q��Ėo��n�򧳙�����*�xƭ��61� ���F���%�5Σ�
�|VG�uc��5-�eq������y�J3ݫ�"F�2�WsMrѰ��s����s� �{�:���T���H��/���tG���u��:��u��%�ȸ�J/ذ��Y�T��3U�g�^�|%�'���l����5e��DW�ʴ��vЈ)P���SZ���5�m��K�+3S�������dNO�ٰ���7��Gq��;�;3��q���m��=v7�]z�c��q��a���ͽ�~q�m�M�[\�Mŵ;�������*�����Ϝ^���e	+�{ՙ�%�*UvgR�'F
�g��U���T�,�xk�,	���<��<Z�/.
v��jm�zb�25��t��Z�ز���nwR��wm^Ҩ�b�3�r��-���Qn�ݑ�v�|]-
��q�+��U�x�<h����)Z�aR�n̬��8Ⱥ��.q�w����7����Ƙ���m�q����.��^��j�
XVmEa̟6e�=�\���0܍cWA���6z\��p��ۋ�M�ɻ��a���q5��[��'��׌�[3�3��I�`��jv�Q��=�������5�9`1�*��s7;�nu܉����F�Ct�δ��|
'�t{MO-�;�V�Q��{�U|�Eho�s����=�Z�֑.fR;=r���
^���#+v�f�r�+F�a�j��~<�jPga�u�Q�>���J��ȥamd��5�S�J�9�M��16̮�S�Y.r �'x�H��@2���0�Ţ#w�q�&7�/5���r�cO��~|X�)Z���ϴK*�g%��Bg��b���֩m)���=���ׁ5>
��!�Cy�����c^�ܘ�rz�d��mM�ю����ݫs,�qy�$�U����r��A���m��i�¾_8e_I��r1��s3�_9�7X(v�R�x�WַrY5en��3�qm�p��9lަ6�Z�N���{�4�
�T��t�Z
T�&~��.@��a�Ƴ��-��S��J���p5�g(�9q��K�]��Y���E;VU�w^e9�Q=��b�i}m��:��+��D��?������{Jv����7w؞�Sti�r�\�um��e���/�v7���e>㺲�F!:Dm��r�u����x��k:{%7���������e�0,01�B/�p�y�݃�Y][)W��E�����sAB������r�U�R�}n*��K�{r:��dts�2�W��1��g��$X��j=�"�73��.�L�tUڞ���M�z�0�v�݁�B��Vz��4�4al�Ŋ�����걏��;e?���X��l� 5o���J�Sl���|�O��t�+9�Q'�T�):���i���cz��KgHx�zA�Q�q1��])�Ξ�r(ȅ�"���T#|�DqW�c�ΣO��mܗ޻���	��q���t^72�J�2wU5Ğ;Wɓ�kց��	���=<Zf�ڕ���f,�[��c�`ـ[e��I�o��� ��p����gt��͏�Dp�aY�sȎj�5�j���Cn�Q�Ж�x�se̺E5�j�Si��7�㐥ze�@�݃�/2��j�1q��\SsW�Ʉ��V�r�v�2d�b� �� <����<��8SIF�t�2���P�|>�S�[�ш�Ȯ��#յPڒ��E�y�S��ߞ�H��
ԘQ��Ш�v~��^#}o)ioX*�\���O�q������಍���ʍi�/���d^6�m������j�+�RW��
��Q`���Y�[B!���vJ���޻u�#�Tz2`����ւ|&�2�}G�,l��U�9�ѪoqA9��7�i�:\P�N���j#ҷ&���w,��������ƪʙ�ݾ��<��yۋ���%��:g��n2�w�Zp~�������Kt�  YyC�/ӊ3���,?d6�G��":́o�M��tn6�����rv;iX�z^�ϳ}�9��ހ�m�g�Y�F#0ylny��sS}��douWk�p��Z�)rt��Z�`ʉ,�S�P�nI��5w����/�#b����{樀نs��}��zs�de�^c�.��R?���L�[��3`�q�2�M�ܤe�JَT�n�۾��7���*!}����a�����6D��]��1A�֣>FH���l��]<��#á�HJ/�����O�d���	��]]�6;��j�.�j���>������ ��
���O�ʿ��M�Y�k}]x�w\B�G\_�=%��ڢU@2�/moWtk�2�:�솹����s3�M���"�����Ϲ��5S/n��l{;;�ͺu�N�3���U��R�H;�C]l�>����=��y%��3�ݮ�x�i�T��'��+���O_63���͹ݐ7�TD{�7 �䎹�@�y^�K6�U�^�a����m��Ӎ�y�ψ��;�,�0���	e����ؽ��\U\g��:�|�����W%�ywa�R�0�,W��}�y/+6�Y
���ͼᗳ/�#�����\��(@f��w���m�m�T+���D�m���+W�cח|\]*z�L�X�_�#m�� {r@t��p^�u�!q�q�K|��w�kX9��/�n�۵��������ТЙ�P���>�e��ŧ�Q�`'�	~|�֩�1�l,&�`��3���u�ػ��	�d;���3�:i���7]��/Z:	�+!Z��%�\p,��aA�(����@v��%e+�⣤�#��P�ʴ�r7�,�7y(?��>����������� �o^�X��<�
ɚ��4wkg���"�G�s��v�`cj�}~f���YwUwlr~ ǳ
��@�y����==�1�t�m�\D6�[ej�;��3?��m1`k��R1h�o��7���%�?#�`5�!�<gE��@�!��D+./�e��[,�',��88З��N���q���{�j��o���[��ȅe��X�^�zޯ_v�F5��
(5���hVSH#v�wK gSjh�h���)5�t{��F&K6v��T�gI��<W�Q�[�i�á�˜��Tߵ���Ig��\"r�c�m�ܢ/R�ځh�'7����s�˽X�=���c�w�D��šw�}�����v��Ӂ��9�씩fbQ骰$۫}�J�h|������v������� ���^���q+����� ����Y��v�ƌǟ��_L�퇕cn�����k�틀�鹰L�Lv�w6,�!�,���Ɨg�蛓�6����F�@Ċ���m+
�-�N���?��kn��5�\�			Rn����T���[�x@�����c����.P\�*�H�r��&+���1����H�	���������G�ſ%�|���{;w�Z��#6��K}�n���ΏP}1k�	�u"��Hkp3�K��>�b�³��ʹ=�L�KPћ��l������\�^� ��F@v n�g����Mr�o#{7s�N�OZWy�E�]�$"m:k�6ts�0F�έ�6ؽG�ft�57��4Gu��p~8�+J���U/u
p�:Cn�f�M��!�������޵�FN��_�:OTI���&R0�18i���xԻ�>��Ø{q؀֙v�Fs��1}�_����Q�67ck]kKG���$��T�֛%���<��*f6�EɊ��/���޲�Z�k���t4(w�����QN,�}��όҎD:2 +3w�-b�bc�9�)Ň�Q݇����q��ʰ_r�s���Vǡ��l<�4�[����O.��**2�];�ei�W�ղ�kH�z��Xy���<_�����<ڦ�eP���7w
����6s 7���%=-˙j���f�"y�çnٖN��k��]Ɲo6�4�Y��'F����͛��u�Z����=B7��������0Y�PV	�݋���m�*�_]˙Q�����۝��A��������湜�}�zS�oP�0*��(x;�۴q��He��S�l��лy�T;�
"d�|̮pRR�R�vR�6�R����Hm�,P��ȅ���xa5T}R�`
�%R,�P��,ny�j�(od?mB�^��������PƆ�גy���{��ۮD욭���v���sj�5j��wf���2��}/R}��-v��aS�8������v��~+J[�U^������-��n�۳Y+�9�����2g[�(m�rȽ�n7.�yV�\$ynGy�N_������ݥ�W��E)��e�J1l�#�����GX��9�ʂU�^�"b%Y���\����)�˲�s�-L
Zf�����ak��{�ٽ��w��=[!�H��~�Lz<뗀"�{j}J�	�e�q�r��[l�.�>�^K��pJ�t���L�'+db�0	��QW}/u���-WV�[:�Ur�h�w3:�X�]vfI��x%��6�ه�4���` ��o��&��Zf�uhu���5�jw&�mF6O�c+�ؘ�>�*�-wr�AP�˗7m�6�svu��y��}]��츎p'��U-Ԅp�^DF�z_|Q~GE�ɩ�#�ˉr�xy��Kr�ځ=��#�7��{�ᅻ�&q�H>�.�
ȫ���bx�ռ��ϫsc��WǶ\�1��}��y�?:v�ҝn�\��)˼���L_;f�v�G7����?8j~�����+/>����V���m��p�5�2�wT�-�Z/}�@�k�>�.��D��\C�����k;{':���>��2<ԣ�|dfS;5�X̸�&-��̯�̞��8Z�����x��n��k'�nު���Tꋙ�4�78�]g9�'���#��s?~}������an�~���Ȕ��5�C][����p�K�G{#_|n�<�׻'_����H*���}�1�Gj�V4���[>�V�}�w-|Ghy����$���\ld�T����<�8u�첫�ƏǾ��Q�(�6��\�{��GO�\���Ӷ�+�U�m#��G����oF���4П��H�	/$�Z�6�E$IH!O�b���a&�79��'����q�g���U��Y�ol�:d�YS 8�Lf
mZ��(�������j��� �>v�sf��j|�rNǅ����w��������f�g�~�R���3
�4tleŜ�;�Sf2�H���:�>��pi�sP�Q��[�����_U6��f;,Æі�e��P�;���x�L;��<o'X�{-�E%#�tF \ļ�i�uǤ蝨�s�	���j2���x~U�`;��K���ʨ��ܳӻм��]�xwDotϬ����7��{#N�E=��"l�ɷ]�^����J�,��lB��Q�;�c���%�AW�SIc���he2�������K�ܘiyѸnDoK�k���BG2/{�6CY�}�!�g�m�@J��	����e=���ť�V���f�}:�lg�D>�HmT�5�:@�a�Ȼ� \_)�oT�y���f�������WF:#��5Ѝ�00�@gy���b���g�G����.��PV���(#���O�O�
��dE?}"�A�|=��H�D$b���$B�(�	�FFA��da 0�@`����9ɗ;r�����\��3�.\�3�)���L�1�F*1�db�D ����a�Ep8�&\��m�)��9r��m��#� l���@2 ���VVP`�1�Aa�����\�rc1�������`�Es���"d����1�"��F1`��1�@2�RHP 1�Č��H`0T��U ăH ��0��R @`1�H�R|b�`1�d2&S d2`��AQ���E���!`0Fc#��Xb#`1`0`0 ��`1V`0!#`1F`10Q�h�E��@ 1F�"y �,7�� `;�7l`
ƃ`��`
ƀ0��`�Ј"�@b(�@`��@`�*�@b((�@*� 
����� ����� �@`�(�@b��@`
�@`(�@`��*(@b�����@b��$�@*@`	��(�*@b��� �"@b! `)��(�@b���
��D!
FD"! `	��dB(���@`)��$�"@b��b�����nϿ�b�
�"H�"�Iˁ]�����>�g�?��G��K��������^_�?�$������=��}��dD U�G����~�EQ�D U���?�>0� R�O����s�����" *�矰?G������_pg�L��0�A9`W���?	D�����T$Q!H�T��� H�� EB"�@R H�T"��H	Q"� ��#H+ ��H��HH�H�H,"�Q  �D��B	H"Q"��@R	 HQ ���@�H�D�U!H"��HD�HERE$TH0�d�H�T#bAF@�#B1DaEa	U@�E� ��E@RAU�D�!�DB1! H�D�� I�E/G�J���o���
Ȣ�� � "�>ÀW�����	?�� ����~ϰ( �A�(?���s�y�Y��;_��G����z�~���� ���P����:�U ~�W��?�>�*�-}�:�  ��
~����?Y��NXPPhW���a��~6��V}�����z� ���@=���f���~���C���>���A���@���~!����
 ��}އ�ǈx�_�~A5P���O�������9�����W��i�?������~���_`xx닿���П>��
*������""��S�aǿo_����������e5��d= J�� ?�s2}p$���A����T$T
��ʥJ	E)�TT��T
��TQIDUUR�@�R�������Z0�B�)��Je���d��M��)	m�fl�J���d�l�۹HB�-&��k����lj�m3i��ebM���ڢ��AjaX��-0�i�iN�[K�r�Z��Y[Jh���ml���k2eSV5���m�jL�U�Q��Y�i���3���+e����kZ���D��Y�cf�V�i���U�Ҧ&vgRڭ�4-�   �^�A�V�G�*٭��m�PR���Ͷ�L���@�AM���R�ڶ�k��m�j�&3)M�ۻ�YldH�IΒ+�����EM��Xժնډ��MjW�  w!C��B�
e{p�P�B�
(^��(P�B�
F�^w
k@�X��6�����u�TZ��N���kf�Â�bZi[U-��UYl�[am�V�q�K df��-����mU�  w��:ȓJY��t��2fKRfd��íʀ+kR`�ThИ&�QݥҦ�F�dU�k��U���[f��2�h(�����Yd�-���U��o  wz����ntT��:� �ڥ[;�9Yw:'mU�7N4SB����i�
��(N�q`蒪�eum��u"�v�r[[��`�%�v]e'�  ��"�[yn ��,�i�B���6���Wf�`M�U;�p 	v+PP��������huP('v�(���T
��,��+Zkfd�  ��U�B�� ��.�l4;�c�R%,�p5��p���i�����SXP�*��m;J��˳\ęT!�ش�VɶW� �x��6�n  7m�  �� @V���  v��t  -spFM  	�
 .]��  �U$�[v�U6U5��b�  w� �( W+� G:�  :���@ �ۇ@ ٘  B� 4�pP g� ��"��kT#5��Z��mi� ��T4�ֻ@ mո  �3w  �t�  ;E� �up  :��:� �w  .s.  n�B[e-����[�m�x   �� �J �k� ���h ���  n�n  � ݳ� :�� �\  ����R�! B)�IIR&  4"�&Sjb  ���R�  �{F���T�4 ��O*�@ Ԕ��sG  ��Mc'̔��
��X�d60%��v� ����@�V(UU}�}_W�}|��`(��`  *�
"+��DW�@QX O�������m��'17�v�L&�{�r�J6иe��{r�P��#�	�v��=��"��<�yM)�%Ҽ+�!յnAz5Uú�X{�DR0�ơ$l�j*6�l��Q�x�u��f ����o�_��/Fbh�R��S�]�Y���եP���)lVò'kV�^ԫ ugH[�܄P�a ��B@�^��*k�J��#�Fm�u�Yj�w���D����L�YQ�B��������%�����J�H�����i����,k��̹����2^���L�(<��u��F�>�-wO)�cU� 
��Vԭ�vG5� z�.��7+t��pQh���4�Ko%�n�H��:��WE��Z�,�S!c9�X�Az�L��àfX����6�݁�V�2
�,�y�}{If����keݪz�L�(�Q��L¡z"�=�H��Tʚ�
���yV����$׵�0Լ9�M"��r
*٭�%l
0wT��Q��\ѝvGo���ݜ_\%�m*��UM*[�	+*"�5�2���{(\�sV*� ʆ�͌ݡ&#��ɱ(R�[�6���c�{B�dc����R%�\r����)���'Whe\���ɪӀ��ٻXrl�&�(M0���d�­*�#8�&�zd���o�a��"l���*�S4����a���?Z�a�
,�
���Ѕ�`�J�KD¬�ku.�qV�61��+D�e`�P�,^�@��;pl�>E��Y�ܺ��n�pF8��
�:m���IV�M�B�H��ш�FdՆ���UE��)��H&Ӣ��{�EA�х�-�݌XO(Mj�+u�cp�^�МX*I�K-��)=i��¡GmCp��8\��U`�v�jwr�Im��A�Ե��A*u�H&M��O+E�˰T�/H�+�"�ь��k�9-���J�f���헴Qil�B$b�P��V.������3���8��%�2�ު��=�lP�q%C�G(�!���C��Ť=D�t��fG0n�`�e%����ڠ�bU�b�64��C,�6X7Uϕ�f��[��$���佖����4Rk@�R�W�`hDb	�k�[r�R�XwlRİ+en���XW����)�I�d��P�㤄;B��6Ie77M��N�v�g/i6�pf�4���V�6J��V�'e	T��L�����;�����жRш!b��*��w��^$طg��0H*�����H��
m'�^�/��\)�$�S��Z5���eK�m�i�Wkt����WO�&î�Br�%�	-B�$Ѩ3�ShYq7��+���	�1�Q�d(Rn;�v��z]P�Yp/�i�E���IƎ�z���wF�72�y��fd�Sa�n���:��f��s��3�C_�I��\j��i4a�j��3����R�Fl�F��5���*
�U���ګX{@f[�V�6������%YlQ�H�*��ݹ��|���x6)�5��0[͙WfܧY	D4sQoU���
��Ra)��Vkɔ1�KDhJk
P���T���
�>�'B�F �����S$w&<�cۡH��OXZ�X4����3�I�/F����Z�����9zmҠO��	qk!�T��ֱ� ���c�l�Zhc�i��&Ub�J�w�U�NW���٢��v�8��R�E1Wif��-KN��0�5��6遌���1�m��ݵ3qJ{7z���mJ	���]'�,!F#$XՓ�{ohpJ�I�t�l,fJz� /R�JΛ��htHXV�S��sVe���:��� �8���W���2����M@��j
�$`�:kk܌RǍ�J�l��I��F�[Sa4a 't����r��/ZU �t.��W3i,�ɢ�7�*억��)J����U�N�7-�=���7u���e(XR�^�kb7��Z�1@��&��U�ᴭ��D2�Ut�������ORsTQ'`5��jV}��� r��,�� |κ	�w���JM����u�!s ,�$��ܬ64[fHĉa���Vn*4,���z��/N�ˡX���E�$�lD��R)��(��-��Yט�q�cjէW�*��\e2��7�,ML��**׸p�Ld8R�C]	h�&�������״�J��K�̸�@*d
grM���E�ԩ��wL%Dn�Q�e˸m4N�1�٤�CM�0�{��"����i�.U� +���q!(��m�� �H�۫Z��B�`���f�x�N\�l�N�_�d��%�5����Z9{'z���Ps�ǚĞ!hS��%�v��Vf��7C�5��:�B�����ZܱR:$�Ϋۚ�$0���C)V�h�X��^b'�оi+E���wV�)U�GKoa�Δ)B̵yQdE��Uxû$�7b��� ����lQ���l:�Ww�#��
�֣e)��-;�4�LL��x�� PY��QZ�~�[�^	��������ӵ��@ pY��k�:�nP���7X�H!%�+i�yI�i���ۧ��v\�_`��aBPR��4VP�O7笱��;��Yq�Q�r_��Y�%��7�x�BEX�5`�yY�1�wX5pܽt��V�<I݄�Y�R�K��D�K5�]�b��[+wfL��4ah���FL��ܕ��j=��:��C��W]Z��+��t۹�M@�Q��e���	V��vv��]�A	4ѓ穋�mD��购�b��ҭ�p�Ope�^1eѷ>0�A���֤�Gt����T50�U����
͚-��T4��J��
�a���W����b�c�TW�e�m�m7��q���H�6����C���(cV�f�kFh���G*F�ݥcQ�E���Q6"��r٢c�;@�+3^��	:k5�����Ƙ���6�x����TcVM�1a�(�$Sf��j�EܳpQO>߬%��tF�n�9�V�
Э˓F&v��f�U��cnS62��v�m���O��)��[+F2L��0|Y
𙻰I"����ʴYքj`�E��T�iq/�y���Jt+m㲶֛��`�%���ʹ@Ǭ o&jFdq�
mGPL֭��.����R��AJ�8�'��^��lۏimfJ����K4�mf'N��ۻUi77�F<6ڦ_��kv=ñ4�3-&m�2��Y,+$X	 Qݥv2��YYr^ s\(�uSf%�ͫ�j%�J���̪$Z�U�+I�U�Qc��ڵY�w�ܱM-�R��5퀤��"��4i6�ԝܴc�M"HE�H/M�i��X�4�`�u%�.�����Tj�d6�-��D��u�l��uzEe�D��fCE�� �m[<e�R�����4en�5- j(e9Z@0A���*)T�ѯ�7yLQGrۡBd7�*ш��L|&1v���8Hմ0��������vRZM��<{���a���7jc��T����l5�^����Kg얲F�6FVܳB�h7� 4ѫ*"^Vd�@�7e5,V#)ͺu�!L	v[�yO6��:h"��5@�c˫)�V3#Y��aóe��ķ�N����<xV����('���$Vj���	T7L(�b��'�]]�ce!Y,H�Ȩe������.#�%*	6oۻ�X�X�L-��!���ۙ��2�r��=Ԡ�j"#�G�Jb���D�	�]Jgoh��E�ז/�0�4+Uغ�1S�*<[���BYQ�Z�(��Z&ؙ���b��, ���R.L[k3n�!6���������K�V>�6vS�"}n�
9�h��XV����3��Zq���THh����H�(%+�5���¡�u6��`f�gf��amKV��M�SV֏���v����f��n�f��Z.Lfm�ƀ�ox+e�0���딼emo`��f�����WS1�8�� "����:&��=2&�[��SqM�6�ՉEA{v�J֖�t%����5�����)nٴ��7i��J:�&Z����&��%���@�&�a�s�>؄6��9� �հ���6�$�%c4��+�e*T�,�B���#��u�	;��DZ�4��0�:$"�%v�����]dۥIՓ�B�j��Z7��(+w6�L���q�񚃃rVA�,��(1��`j1�����vakF�rX wO�*Qb��G)R;���z\_4�#{��l�`�Z]�x���ttF,ՖQ���5�#<��w3C�j�a��os.��]�&�5Y.�I�{m�
�o r����̬;���gV�Ӗ���՛�w�I]@����0�y%"��˅����U
��,c�WW����X��jS�d������`m�(�i���s��K%,n� Oi�йkud�4ME/�)��[�.Z�w$*�]G&�0��`=fbɔ�1�Z�ŻV��rJC-2�I�T�G�7U��.�
�sk^���4�����n�ZqǦ�mn��fVI��n\#Xn�������x2̣L��"��yX,�0Co&d��*0.�3C���j�Ȥ�7�����T���*(+v�eFp4m
!ՔsAV�YPx����=�t�C��p�St��ek���b%H��ۙY�����cpJj�ӕ�
5�' 7�7�W�cB-jP�'a�Aٔic���U�FL@�&d	me�DK`A*
��Fb��h��olXX������#�UhR��5��t��@m�dV�S��r�;Z.�]��=��Gwh�Z�b[�7aX�a1
ڀ��ٔ%�PV%4�$��:���Ck洬��-�s�1+]c��.���
�l�\x[�	V����ؽ���'6,��)�m�Q����`�������Hwu��jS�[PA0MҢ)9BB``�҈�뤩9��&�[��t�y���N�	�B20p���k�<7�^N�=�&���9�ջ��l]�l�3K-����D=P�[I�V#kqJ���Z��"pu������F+�1۴>1%d#oYҝ
�p�����K�YK3h�l�C�Praxr�T�!�Z(,��Xop!,Թ,֭���¡e��~���j4�%��9�QD���Gb�J�L����z��Z�
�ȩ���$��E^fa�� J��
&�Q�mksU�Cp�wIT�lش�oq�۳z�i��+PvbJ�i��h��t�̖]�#q����5�5>��k�~d�l�w��mI��-DZ ���J��6�	�%j�PFٵ2�*�X���� ��X�˖vM׹��'�.���b��v�� ��n��e�&�*3d,���qR�RʬS4Z)�B k��m�wpY�M/2Dr����;)L�:a,`�{}���:
"L���
=��{yf��"RlaV.��X�K�Ε�:�o":���$�S�e<��qU��N5�]4ܽ��]A��Z�r�ЃݼX�� �9�^���+��5���qF1KM�3o��1S#^^彀XY$mb{����y����v� ���,ڈc�&at��mŕ��Y3�34�W���(���b�q
U!ܦ�3NՍ#ӻ�wh�Л,}�0cl7���ѻ>T����+���-�i���X��)ں8��wXvc�c.�b�j�!ڛ�5�f�&i�9m�n)��fCm���tfF��סX�\��Ao#Y $��[�jF��h�
7m�g+5Y�&X[���5i($PîKV�̧�7l�ռx���Z.#BM�M�n���0��l&��U��+f�>��E�h�3��9ZRo�S;N5aӚ-���Z�Sٮ%t3FQ���spk5.�n	��jN�\t&]��� �Oj=6E�@|+'��M\+�f�]
�R�e�\36��w[�PFKhL��n�j]��b����:ʡ����gt�,6�E��q塴hʚ�R�*'m�Cenƻoa�ҕ�v6��Mb�ɚ������N+�Z�:y���5%���d�j�d ��G���B��tӔ˵�[t򺸪%cC�7��	��n�e � �+�ڔ�k9p1���S������0��{ԭ�(�-ջ��f�:t������JE1�.���# ���g,�E��+*�(�K2����%����M����j ��[�p��u�;��vB/�06n�3����v֥�[V��uM�SM^�D�0��(�j��
�`(0:�pI-e4EJV2�m;��e�8�õ�K���L�(+�bn�m�(<�ǈ��
���(ɂ�������i]�w����U��Q��ؒck
RQV���mk-@��S���z¬H��9�P�R]�ٽ�**�N�˽:���a�KF^�ѭb��hKV�O�Ǔ7j��J��f\F�!h���8���U��b����ƭ��6��U�췗t��̑4e�/��hR0J��2�s"���Y�K��i�ĭ�%����� $������埮]�D9�P��mS�� �­��[w�%�ӻ�JV���32]2����*�l-�.����w[4��lq����-ɏT�k"�]���a+,<�5�5�o:���[h�lm��խK�(�4I�j�#+N���Lݚ�A�́e���l���J</ ��=��O���à��%�e�ؠ�Z�CUhVkB�Ս/�&��J26)�"ܫ�ݭQYX�f�dy ��^��L��2�w$�U�@:��w��� @+p��2�H���ɕiֺ ,u��J����;�Յ&jd�^nҎ<h�ܼ��-Y���D�wH1,]��ok�a�'>�&���.�pd]!��efyP�{�twEcd���|����E��W-z�cU��1��F֔� nGR;�0pU�� ]�gF�{U�ů`�� �!��$-���g頔��`�����J�%�	�V�v�;�M�K_hq�b�I��C4����ը�2��²��0wN���{9i��m�gm�N���
�m�ƹ�A�R�=�w�n<sG.���hC��u�o$r�6�*�.p�&0v]��oق筹�:}l~��ȢG���N}�nn1)hNwR[$gA��u(bZ�٢��*�Զ�0f�/I��ē1�Y��i蕁,{4Ce��ݵ2� �!}�/{�p�gq�[��B���'�5�{
z�u���U*���oI�:o��n�R���Zv�������8�wQIgDÚh�N��}�HI����nԶVi��o�J��fa�/`΍���zoљ:g��3�wx����H���}��{;_�J���+aJ�R�s8SU.����Z��l�D5�z�bWffjUD��+�I���b�Ր�Q�*	�3�>ݏ�9k��֎��RoU}�)u�z+;�+#Z��<��ʛ�$]s�m,�B�C�o.tnmnc�w�{]fށ�^��1��n�xU�(m���<1
1LҰ��$Z:��ipju�*!�٭�R�!�Ʈ�N��\��X�Z�EqN��^�3���<�YF�{������"^v"WZ��wm*g�' ��|!��Q+c.l��ߚ�[�/��oEdtm1����.P�xeg�)�2ޙ�k�N��"�
���8�XÚ�m���uԱEPd�+Y�7�e�ս-�!���5v�iҠ�y;:-2���[��묊ѝZ-���@���*v�cw'R�g�6!Y��W���-��ƨ��w�������G&l\���×�C9�]�[\��G"�l�5��H�&���@p�붔�T���G��v��͉NĢjv��VNրf����QUҲ�'\19������`��9qA/z{���tO�s����u�8���/D�)/K��}z��s ۨ:�d��ok��ZP�+�g�1=�=+��yl�\�s)������SϜ�]��.���MyV��̓k�x8�\q��t���k��x��w3�_Fb;v�7���u�8v����Xk��;���L�#l> �
p�{�C���X}�
�o
�i-L�]�],
����/���p�6�yi˕{$��e��"���c3�4�Z3�Ԭ]�D�J2��8�
��\D'X�
��k��c1B_;wO���褦n�EU����n�<O�0p/��[|��?U0��Y�D���m�(>�{���Z�6��lu�v�U=S��\����<��Z�{�p�ܴ؂U�;vU����#oN;�s��{X�.�f�8�"kS�&�t��fѹ��!�·	{�+*K��O~����+�c�Y՘,v�|��t4���8AY�*��s|{e�������N�E�<]c�%����5�<�Q�r:���k�ѓ{�:�^���ݾzk$MbTUo8�/fc���$�N�N^�ۺ�*8��L��PȒ��s�Q앎���#+��=��nU���#BN��U�-�}�\��6��,���C0;{ˣy������Օ�hй�\(�����uu�Z� dO->�k/Bu�a�r�h�&�
�4����躗�^	SU�RvRI3�x�{c�������kJs�eƇ19�͎N{3����_0=�L���f�[EƝ��4�sv��WW/��`ų��uv3]�g��H� ����K�C'^�$�a&'K��i���6��W�/n4�yO���f�5�/ ������֥F��+�&�G;����zWb;�Qf4�]���}��eP��
+LK(g8��h^v*�A �:MR���,�O(�w}��+�R�����րXtn<�������8K,�ON�7P�n���r@��MW��2��̮��JFwSכx������������CB���X�0C��۳�q��kl�'>3��JB�r�sV�,�#��ʾtv%�`bs5�RSՁLy��ݶt^��j�`��fۙ�+�$�l�p>G�Ӿ�_�V�Y1��B�)�� �/��B-��N2VN�sa�kt�ü���.V�#�4Fj�r���*pL��q^�
���u�y-�����ecH7Y�c�XZUɣ��09� �ڕ�ط
�b�hw�I�N�
���/����'��Ci��C'��Oe��[@�X��rj�kvU�2�<9�y{�ci��]�^���
����e'�ᡢSOfƥ�����+ܩ?q%fn�������i����K�S���D���;�5�c+#�oȢ����*���_ p/i���b�6E���]�p�Ƿ2��{>s:�0w�����Bhpg��ݖ�n0�s:U�}ß+�8��5k�v��ItO��ͥ�o�#-��8u�!
�]z2eN):�b��0�h旗]��V�&7�]��n�``��샪f!�Qve��
}VUm��*ᫌ�=��V&M�}Hl�*�,B,� ��&���xm�Afe�=EX�Y�ɭXHHNe��s�Vr�`�|�'+}W)�g��	j����%Y��*�:�i�ͬy\Y�z]/qZ�N�tt��/��o���:`��^�(�6Ҿ���v�	�{�ĳr�yL����.��Ǵ�N���K�� J�FҩvS��N���#7��3��Q8�^;�+7�(.RM�2/�[Y/� ��(�W���H�-�*#5�"��ޜ�#��lE�oG�����f�"bM�Q�}x��"����p)�I��`Y;0�;�+�Q#4l�6�9�F�-����4w����G�닞{�w�[���ۚ��|7L��Z����W��E�m�r�F�(�㨞^a{l�`˶��.٬خ�Lk;f�haX@���ڼx��*MY`ˣE��N��.��d���>(A&-�� /z�.Wx��c��V���X���m�:v�٣]تo1R��j��qR���s�`���,{M�[�����#s��p�����n]	b쓕������5��(�S�:�j�=��uEǆ5j9�q�gu��B��B��=��Y�t|i�L�'Z$|*>�Bn�L*q�{+���jx�lu����29u�H~��`j��v&�[:!V/��������y&Y�0�b>��R��{[y�>�%S�ob�.Ӧu�1ֻ�v;��y�$�,��o��[W��J`*��N�{�M��3�:��{�K=lԄNԧ3-�kP���+�e�H4r��{V�� �+6r����մz̝Y��(���¶��+k���q��͕|,qZ�ZŢ�s�]�At�ev����k:�bo�[���8�no/^Y��?=z��2�&�(���6��E�9�t�=���k�S�������K�Mv�_8 S[�g׏''w��v��槦XC6qfR�0GZ�����WZT�2�O{\A@�:[.����Y��6����xQ�z�(�E\"ž�k;���5�0�M��F�c�m>���!�M�f�Rߞ�9:�����(l����n���m�f.�r�{4r[���!�8CZ�Ǿn�M���j��!�7WKv�E��Bx)4{���&�{1���;�U.��z���=���n��z�`K~Ҹm�&^U��uK�4b�7�7��kuMD j:�Q�s��Q�I���z+��Bo_|z,�o洀O�V7y#��V��;���3�,@�y�C����$n�@�Ci�-;ma(��}� �^���I�͜ϻCk��d����w��)�F�W¡ps�y���2��:jS�Ag�z��N��-`lx�I{����hodf��H{�X�ʟc������Q%h�{۾�K��Zϩ�����!�[�N��8���t�[��V�Pڅ�,C��"���лf�7#�)a�k���;�ڝ�b������\ģX�zM��t��Q�����Dv5Y�n�1͗6t�����������s;4��o�H�N=�AC)P�̳oI���V,�;���A�U($�wzW��'.�c9��M�g2�K	3~ؙDpJ�X��s�^ĩ�b%3;�q�,���"�Κ�����r�r�mN�����O1�8{�����='
GF#�4���q���uX�<�ǝ�j�5���S��;9E��Y1���|��e[z��i�٫oft=���������A��>5�����O)��d��\�s�����hZ���c�Z�j�d��B���V��59�c��K�UΧ+֯V�[6�q�Y�M�K������6�{�l�f��Q3���/�h)���,�|�f��9�T�3%sW��X{f�s7�0�NYYa� �����˼��EdB�U*�I5+a�@ ��LD-�/VϦ�Z�l)eՃ՗�'�%q��s1K�[�ns������f+�-we�t3�qMQ�t}����u�J�N�/r��E��2��LJ��F|ેvFپ�b�1����x���;���g^���dR��u��Bn�j��6nNC� ��E'Ol��> X��!:hWm�w�6f����Z���PF9��m�5t�Ϟ]����T��T��qu�ꍋ�7X�ܝoGY���n�j\Ѧ����F��K6ol#DJ���y��֝n��i�fPz�����fpf���H$�nT�����u>K�>���qJ{H-$|�n\�K���Ƥ{ǹW˴�|-��]��=�n^кC����rHa�Ky�}�
��pH��}J�c����(�a�^�@8��W�%��_��3���Lb6�"8�Y�e*�ƀ���̓�^u�'��g�J㒸�d4ꢲpw�숷�1ޠ�\�vws� ZũYN��/@���}��Q*��Ϻ�w��d��� �`��h�%s,^e��ۂ�N�_t�.�MAW5��x�_z��N��h�}�k$�Aʎ-�}i[i�|�j���Aa�[r{p���f���i����vȯ�$�\�ͮY]O���gǕ���\��z��' 5h��[�g5X�+���	$�*��~|�k=��M�X��8{�_$��{Oz`E[ޥ:؛N�;�X�A'kgs��k����|�]Y��l��/2���R����}�{ν�fIR��&�,=5��˾e#V����}���E�-�7}\�M��T�L)�b���u�Zy]��
ի9+{|ܑ*X)�GB>dn,�C�'B���F.�lݢ��|7b�JK�{j�N�-�:����L�[��Y�aG�cjM��N���_r�aZ�=Z�c�T!��T���6�die���\#_��=��͐�T]eb}ֳ��b��Ɔ1�|�V=�9剬LZ߮]!/��U�t,�%�˽���Y�8b�.B���b܋k>�V�*]4l5asv�AT����T��[S�ͺo�������"�͏ �|�<����e�f`A@��<Z+A9.�/�����b���һ����24kwP��n˒��K�7��V(�9f䰚���rtI\���2�w}0\�y�fblsC!����&���f����S��%e��DZ�0���2Vŭ���.����=��9+J�ru�o���|��9���]�f�E�u%�ﻮ-7��|�	̎W&ۏ�íu�4��ٿ<�X�j�j��B>\�
fݹǦ����n�.�m�r���B������lD-��xv�u>j��6���xa�Z�w�c�K��MRt�J2�9OM�ޱ��^=�$�^�Z�yR�q:�Hy�� �K�O�E��p`�ءzWf�H<�v�.C��vf�k =���8^��a\�el^s>�:F���}���f9�d�ӷj- �]�w���R���E
1���q�Wtst6P�5��ov�dW%Vu��*��h`���3�l�Ymw|l-���^*WV�9u�����зX����F-�q�6���A�����	z���u�5?m��{Q�[L����g)��4��e������[�����R�,D��S\�ޡ`utM���7S�G^S��4r]�p�^;�Ro	;������`ȡ��6m�p^���;ّL����a�^c���S�������g_����Ϝs���P8v�L���tv�J��3�S��� ���:�f�!@�^=��~�n����t��i;���d9�n�%1h�ѭ��%ǑGV���\(�ޕm;�D���p��<Oo8ӎ읔��b7���;��H���c/C	�����\�2�
�̣{AHI2�F((ؾ���|�:�RՠY�ݭ�8��}E�.�/�gJR�o+}'ܶ�.�ܫ��:ד���w��!bH��C]�]���K����ASe*�//��`6]�r�mJR��ۙ.�V�����!�eܾo;�ol�e���ǁMX���u�Jۭ�+2��.d��},ZSұ|ޅl*�VQc2��hU�d4�N�^xϞE�F��\~7�N=q����K)`O�WG�S͛F0���.*�.܁��]ޓy�uv�na�}i���*�r�6��?M8|3�;`9�֎y�"�t�4;�|N�j入\Sl���Q1��	:���J�
rӹa��;���Y�])	���s�6��Ҝ��Yg��rxΫ����+�k]���cz�ë�P��%�٘v+G��o\�.��t*`ݗ������{{���e����H��w�����-�]�Z�����.�l��WƖɷX�5-�ڙ�+:�,yy�S���T7k_ݳ:�cip�ȫs���g�j�:����Ի]ܖ���Z���W��a�h:=yxov�{/>�{�T�eX�|y��=n$���� �  
��������޻��~�}�~w|>���?�p,����3zE>��/�d�ab�3,�Lg
�[A<:��4���MvX/u0bޚ]$����kFX�_<P\/�w*BS7� sp��	��|;5�=Ӿ�S�q;�y�.6(��U訶�\�ӏ��7�6�1̘�[xxm��<�v
�B�ΖxU�/f��ɺ	9�(.ۂ0��i�p�mkR����J��Ү�[�㣟ev5θ�v\�&��F�ۨ��K������}��뇷9DݙOD�Gܫ�\�8��m����i��c��[p$�Jx��fsY�ؔW��n6���Px���*�����9�8���"Q�'��������A�ЊN[ŭ+��M�zS[2�m@M��8�|��R����l���C�U�Mo���6��h�n<Mдit�A�G_P��g�z�����pZ�>P+��LZ��^$k����sT����r����gq:�ܗ-�1Ȧ��� �f'9CL��h*�םͭ���U
G7:n��Vrt�'*H��ZLm��Ĺ�<E��NN����Ѣt���s���ޝ:�Vڠ,,a\����T!��B��˟��˫�iV�xv	V�hw!��d���ˌ;̾K�;8�N�_k7Ճu��`��沍�Y�_S5Ӻ���ƻ�������
��u�q���y]tp$�Wh���.@�*o�br��`�xu��bJ�#;�A}�)|V�:ᎄ ��F&��������T��6 � �{�@��L�=V��@^&g5[
-��qź�����	����[��_#�_S׏:�N�����1Z27�}نԮ�m�6�P���en�ժ�z�Z��r+
��ǊM�[�iw,��|9K��M�K���+�q�]�?���ׯ�"�EO����m��I�+�Sӣ�A��<H�VW d�Ϊ�б�+4��!)0i�%���`�����ƙHݖ���{�=��.uGT�]�d�C{[q�.��[lZ�V�<[��[�ew.��'eǖ8�����la�A,,h���M�w^e���3�2�~yM��'n�������0l}�m�N̶,Lh�
W�����*ٻPR6�waF����`0��_��_]� ���z"Ӧw[έ&ɻ�b�q��b�lAt)a^�A��WY��U��M�8�Z���
�"�)5������g��7�7eE��lF�k�s�G��0!�2Q�kf�N�խ=���v)]%��V�b�Lxc�}Rm�v�Dgl�r�d�NN=�{��e���Nm QOo���nj�Pԝ�!�oX�Kk���IFH��%��+�d"���q�/{2�-$V�a�0�Knj8^�����.�*��r�Ã��^�P���θ麸7��Nj�B!�F;��5`�]�j1�L[Գo;�Zu���Cݪ��F��:jS�ں��0u�iv
��1bR�o��0�vN�(B��)�w��۹���gvc�: �,3�����.��2���vF�G=֝ ����t/�v���ĭl���C���N�����Y-��V�Ks�t�͈��������"ɅM�Ci�+WD���+�'�������%AM�~���;�p�����	>�hg����Y���O8��j<@x��\wf�&GBr���-��0Z��6;�i��<�3Pa�t,Y;�X��{���H4VZҫkj�XiK\�;�O��.;��Vvn��/Sw	m�ͲU${�t�D�Ϙ�x�^���au[֚W�l�v�[��/N(w4��hI�d[��q�H�bO��u4`�n��׌�����Cb�r�񋜬��}�y��26�
z��ƒ���Q�<D�#��/VY�"4���A��X�s��CPm
�/��٢p���U�φ�}��te�W�M���w�/�xv��ǖ�`ؒ8���:��Ú0 Yݓ1��9�M-3�K�
�]�\Ɗs���c�e86�4��'��w��6&V]�U��̍jkT�V8�|z�r:�����.���;�v+��.^[hS�33C�	2�h3��Ϯ�
�I}:e{������M�n��G2z�T��k�kb��pc)<xyU�b��\֎6�J���C�0� tQ�)N�����UFTB��f�M���Ԣ;�<Y����f e����kK��ӹ���F�>f��������me��휗�rȕG�s�x��3J�:�%p�X{M�#X��;)��sa%�w�%����ɬ]khR(��p���8ݫ{�5u�&+�����N�+�,���M�E}nR2"���X=�����rۘejd!���pb��P߲c1�לfҢ�t���A�<�ͻ�wG ���D7x�m�'\7VT�;0�.�.lc��섽�ci�\�\	V����ۢ�f6�N�hB	����sVk�켄����Y���K[*'��5蕊rj�=f�ⲝ�iPmt��]-�� �ܫ�ǔze�u��j��hnHC/E���oC2e�7���v�]�0�1B�#�]�����)㝡�ǹ�c�tW\^�j�'L�*�f���lU�̧r)�n�t�1^��{��������h!G����ɇ�+��6'NPC�_^%�������E�3�qu]1�ۯ���h��r-�_u[JvJ�w��`�6�v]Y���3��m�%jҟ��Z��0�L,�F�k�G�cqZ���m�v胛�.Yyb�;1��ox�Q2�K����]r(A�g�Ifq<�t�W�����k18Ѡ/B�A��j��k����/=�_�bB��`�_u����7�z��
瓭�&�r]�Q��t�]�O�y}o,n���0k�Zf�!<�Ɛ�u��ӯ�6wo8C!Eg�p�p]ź��P=�T)l�X.U�� ���`2�u���]����n@��n@���y+%�Z��׳lTHwTۅ��0ӫ�5!�.{�
����>x��$�gg�HZ�@駖^#���ǥ���BJ��T�"w�f$ʙw�e�>�6��CuO6������y�=u2!����~����񼫄�u4�����B�û��*<;)#*�2�'(h�g��b%��)auY���CJ��='�K-���;\/��X�*r��5S��-
K`&?�Rk�风��:AM���P�V�^��S��r��j�̆\�(��4��M޽}�뙼�`��-�r����D0V)BTF���3}f�\5���2a�N�'j�¡�����PUb��WQ`��h��ĥc�w[k�c��܃�b���1��;�2�y����f�OLcJC�}i���Zj�t�h��_nm����k#���*G�ve�X���ə��.S�����vbA?1�$ߛ�b�̽14�m�s���=��,�}%�Yr�+K�C���B�+�`�%�_��+oU�`���7*Jh:��L�M�hY���cC�}֋G�ލj�z(5�΁Wln�Ԏ\�J3X�bb�[��x4o��o&�E�ۚ
�;�+�-5���Z�\Ɋ'j��ݾ�T>�KA��@��N���`�+E	Wbi���Jδ.����[r4֜{�fJ����[h�9��*=z�� ��<��\j�վ�T_>�E�P&+��;9���=TJ���H�sS���W���t����v����N{�z�� Ѭ0k嬎��癵*�q䰥^ݿ�J%z�,�B���T+�x��k��Xk�XE\�(���h� �K�M�5�*��3���s|S� �L��C(mjj�-�.8�C��9�e�O�O�TE��,�������m3yc��w��%q�:ڳL�SN4/#�XqK�QՃ=w3|�=4nU�}�t:��4�<֮�&#:ܣ������.qg#�7Q�M�]���ׇ��z�x� S����N�p�$ �}�qu�#2U����|����TGbB�'����c���l :�����wyX�cj�WU�}0�����p E��E-�9�T�3������6��.P�âm���R+2��VC���B�t�x+��	s{�����+]�/,���e�5�x�o�&{F�ţGqc��ekgy�w����W�yz�����R�f�Ŏ�JcU�2�:(�wf����al�.,߮�㏕%��
G���lZ9�����l�CpH1.;׫N�	lh�/YVp��P�MRv>�	6#wi%Y�6n����t�%#@V��w9r�@��$��b�G@�b�:&�#��]�L��a�0��S�A�*ͦ���ʼ��5��
�}�s��J��7�5t3�.�05RY6��D^������0�)���x +"9�%�Ѽ����{�5'|��t�R`��5��q`��Qe�)lT܆�K�
���~�9N���3�,c�M�[�1��{&wCF��2�ĕ���V��>{�B�x�^ (b�7h�Ž�Ո��ے���_xm+�N��{-b�&�'<߾U�)�:;���ߺ�g}1ö ��j[�'ٳ�p$-�U�?�Mb/^�l��R��.�U�VGϔV��J��9��&��K)}b�����6n̊V��uv戝m�1��	\�N�}�75�"�w�:���u���0#��1&���Wk��B4����g�e�%���Df<9�9����Ɜ�fxa�-P�{Nm����Uo���j����4?��ݮ�#*�ʺ��+�n�&/Y��ڴ����x�����F,���J'������RJ����)7��l����z��z�|.�75F�z�fi���Y��ojJ��#�+��n�ԑ���)$ŨuXC_y���y8_{�o�闬�uk!z�3�����䮡MY#M�Z;���̃#M`W��RW�QP���8���x�L.ʱ�������Twz��Y]�v�ʢ��ㇽ]�Q�]"���^�X\f�X�eV��]
�e=n�
�|�gV�E�7�k%- ǫV�.��7;�o�t�nV�Nb&�l�t�����b�8�-e���Iu�oH>�»��}p�P%-wz宽X.��\e>w/��K��K�]^�!q����0�:R+r���tM��d[-ȱ��(Ĩ#���R��Ђ$������:��i	ǞMr�^fu��}�+w��,����gR��)!ǵQk)���E�Nѩk��ž�N�ly�S���64�J"�-��:�"¶4�c��'.d�?iM��K"P�^���Z�v,�Q�C����m�i5���<������l�Z����o/���9�����Íґ��}���v��fw"=Ŷ� �\C�@�8���gٯ�2�vѰ����!��qwoh.kc�,�;�����ڠ��⃽�tU�k[���J�Q%��Z�	QcV�)YMbBV�,�t������h��rԴ�2d�/]9���g"H�%Nʻ���e�km�M�"�0щ���~�HG[ǳ/��}":�];���:�B�Ƹ[�w���B�,e֭��⊇LԊd}�V��fbf�g����YE�=�v���zse�2
���Ւ�zd'��(�u�_)جq�ɺT��{D�]k���T.�.�n�rh�������.�=Z��ʎ���fQ����w^=�/��K2��5+C�h�@S�y�n��7��h -YNv]�����_kT�WZ�^�y�i"�w|i�R_n�:��3cѻΥ{��z���x��	�.���ԯbwR��s���ጶ� ��r�4���_z��4b���x���49T���m�-��;e��nV#�k׎X�k��.�7���X���|��]2��Sv�7yIP��嫚S�T���
�����s�`>��;5��(���7��s+���f?e�(��iI���Х�:�!s:�v���V"&E������j��S	�ik�҇�㝝����J�P.�/������-]���[�\P'i�˭�TVd[]�����3Z��H�ov�*��E�*�+�d������k�އ(�t�A����x�z��-5y�}wyNƖ�j��x�緇�sVo"s�)o��n��XZNgX�Fa ۾N�� 2F�ы�%0]��]��ǃ3(�X�=%�:��U���Y��܌{.�ܽ3tu�s*��ɍ�]����Q�4�ʗى|If1�l�̫G9P�gYy3V�\nC���X������γ��be�r<u*�ٰ������LPL�ݿ��`Pq1hˤ��+V�W1q���u�eL��#�+���M�Zϰ�,B��
���ˬR��%�Kn��F���ګ��Ƶ%y@YA�9����&�
}8'���d��a�&�����_b������.`F�'m��ǌ��ɸ�@�3#���8lX���;�S jwu��7[]�҃*N���w4l���2�y�0�4-`�\��n���V�#Q��.r��v�[�XW�ޗ0�u��
���o�%]�GSw��<��CSϙ-�
yvY1��R���DH��X�`�ͼ�J��nj٭o�31R���e�כ��<��%t�ݤZ��V�l�v���u�L�&���۹��k�z�C�ND��C�݁���Iw|��-�{aٖH�U[&�n_m,z󦦙��yD��9�v#w0q���8��#m�6�(ɶ��sT���w#b����+PẌ́rI����e��X�
���u�tq�X=
�Z��`�zg"f�F����X�N�t�M����"��E��rmٺƞG�աCq1j�t���}î��X7�{��hW�TQ{��U�;���$T���i7���.��[��>�9��WKkr�._q"��cp.�;x�u����חӎ����I�dpcɒ�=U��
�u]J�PJ�S/x����ōm�	VΨ���.�[�����w�6�{e�-�Nl�1����s�����������˾�'�
�����J��������&(�Z�ǹQ��y��C����W��X�X2�>��S��3e^c���DH<,	���ywQ��mv���IaZ	X,��F��%e����3��f|=Ӵ/�샕Ҋ�&kiR*˳�yOɊ��l���p�w��vp��.�)Ք�o5I���^���P�J��S��v��{���Wwg4C2�'����l�x�Wyj�̵r����Y��>ŹY{��Gx�'�W�P����@*�ۧ}���N��]N�-��`�b֨Y�|�烏��yo��=�� ����vo1ɜԻ%�WN�8��v��r��w�Gh;5p��N몷gLbg���Nr7yL�{Xڙ���+��wQ�d� �H�QpL��q&�>�Or��G��k�\-}���ٺZ{fLb�CC,b��*:��� 5�[�s�'zD"ߎ��
�@9)��dd��!aV��s9�pl�m,ѵ���|Xx=m<�>^Roi>�/�C+mX���-i�701u1X�j���g2c�JclU��S���������N�֐���}�H�B6��p}'.�b�:��O#��Í��:@<4O��,�w�%\3�gk�~�;���}u%��׋���%�j�7)�j�tч�yn�q�;�&�¿��?1�%������#}on�ce���������[��I���
1��D���*b61�Q�5��b�����4b���115�I�PSADLQrIm��p�I�TRL�i2DF��Pm��f)���b6���UFƪf(����h�EU1����֍j�-�kUZ4�F�J
�q�Lj�sEN���Z�KA�
vժ315D�"�*֤��`�c:��)(ѪLZ��h�i�I��v�4[5��*H���k���ƜQ:�N'Pm���"4�A��q�QZ�[&��m;�8�DAshb� ��ګTCF�����a���J(֩�֋cm[A�Q�"Jfjjfb��RE8��#F��l�m�D����bb��
����MV��*�Ui��
Z�60[&�+K��l4%V�JZq�[|���>_�Wٳm�f�,�`��ےnq�<��"ō���ښѣ��[��ٰ���Q�����#��賧h�����n����~x�o�����e"{�
�%�[�_Omh�X�E�}��^S�*S�*�̫�|r����R "�Ϗ��.2<�k�]a�>�tM@��w����B)z�2uu���z���#�F��/c�D	���뿌~�8[�[��E�*�)D<���������f���?g�(6>N�K�~�������b�\B�ud�=x��3�=���9<��BD4�����'�p����DWإ��̌��͘Q����×2b���}�S�ܕ��(��2Ō�b��zi+���a:�b��Wͽ7�#��Y��d��۩�\��_R6}?�u���y�0p������7���}颋�}A��񺽑_eF|%6�1ya}�z�×��a�l�������c5�@�_���z
�
�������*B7�e��'�F.�a6 ;��J�����P׷���l�+=��v��y�tI����tm��g���s��Wy���W�C�)u�e$�_4�/�u�g"�S�$u����y������s�ˎ�XJ��V|�k��'��\Sw�SC�Yi��x{��W�Hh�VE����@���[��(d/lܘ�Xxpn�ڛ̳۵�n��,ܻR���Y�����ʆT�Dv��R��.��T�U�,o>5$�R�Ἤ洩>�Ͳ:�U3+��'�i�g��g��^��Sh�|����J��7���5��Ge�Z���7��&,5�ښ͔"b��B�.�����D �n�C���|{~�Ta����Y��!v�ZD0w�U��}n�]GX8d�I��9#j����1��+Voަ|�Ԁ���5Ơ�δ�CjS�Ä�w26�b�f�*��s�S��r��џ:�^�3@�k�8EE���
H��Qe:&ۃc��Ỳ_ӑ�.9���,Pɘ������9��S�.��\�; uCnȫuP@��hӒ��xT��C������\��t�=df�krzh�te|�T*J���i}�2�+��=����'��h�IA\��8W���s��G����]R��K�1��ic8�(d��+���\U���U O=��9�GVGq��ʚ��a�'�Ny;�\�,�J�]�����U��{f����"��ndC�J]��RX�u{ڷF����5��8�����K5�j� :���}�׀�������)wc�Q]�F,1����]E�v��''A���1�9��@C����ܺ��4+m�jƩK��ڏ��C���󗵶���g�g\n=O����nn܄��t=!�|��_TA�ӳ�ײ���FO6�%��s��^k�*dn��7��H�_}
�����r<��֦0������ ,:ޤp��`���Y֏�Y�~Y�x��6:�J�w�Ғ�;W#�-�n*� �gE����zS�V+����n�±�#�?�vU�L�&j���!�k�5)���e�}�*��r���5�_��(�X��<��;m�f�%<By,�$��<yϧ��D��_ɗ�g�2#kW[g�Q/�aa�ꌸonx�x�� ��#2�L���ª�K�����h�y3T\��iaB��0\=�|c)��j��!�[�ɂj1 ��w�����&ft�����?:���s�xʴ���_�+��8T��ݷt󵝧(�y�;y֓�7�� Pq�*��x��K�(��T{����;�u�f��|~��@;�9e���h���mI��8��Z�*W$���H��"/������9��7%�%�<������c�L"��)��r,���7NJ0�؝�����
7R�"g��y��+-߂��!=��ڪ�SNzm��Un����k��x��+���q��	'�2�N�����2��u��q�(�,�ܼ�X��u�jt0[Ê�h������Q4��/:Y
,;�s����૟$.������]ҳ�y��<J�58S5X.�c�bY:E�e�9{d���޵	���t���Cw��a�c�{�.���@t���p�I�{�I��1X�G8��ьC��%�֣�d��������
�����(V�"�' =W*�P϶._Vu�AӌK>�� [˂�P��uE��uX��O}�X�t3��w:�N��"�U��[���/�s��i�h�]F�}�xT1��;$G���l:��ٸ҇�����`�q�
�GK�r!��E��Mk d$�Q����a�����&0T��.��:�5���w�3���H����o�UTD�K�02S�9��E�xwL\"ᨗ GqHҮ:�u�u��/R����(8͘�X�w�!���hh�hWx+}^�e��dp���9+��gS�7�ٴNYuL`�����:Ks8��c�!V̄2�ҝ�;�71�.)��##�6u�S�z�e�zz��m���pg�p/�F;��<�H�/藆��jUW�����ɽ���O�U��v�[ۤ8J�0]wcB�U_��.�m3 z��>�_��'�aD�Z�zn�\�$��Ұ\f�[�N�ܴ&[�xIj�HՎj6��q;��0�:�,���xrj��]�R�J^�I .��s��S��+tK�kJ��i��_D�*��'4�2��8{���k���,b�a�)u1ܡ����y�Ԥ��t'ʮӃ���b'�)�{*Q��DP�-PfH��U 6չ���Y�X���J5F��4s����4�#=�Di�e�{n����-L���xn̴�ʼ��܋�kX���X{�B�2P���#������`�q��0��	�U,F�^˵]*��a��$C�'B�pJ�q ��/��!p�X����=mހ�U��Q0@��TV������� =�ܖ��I�f��]9�b�p��K����]�<ap����Vו�pQ��E�1�\���2��py}�y_\dy�x��J���"3�QcU�ܾ㱊wq��Z6t��͖��/(��@���:�^c��Ϯ����O=j/Ve��s�Y�I�i��D�gLb�8�����g(
�����ƙ�c4�e�j=ut������7�8S��:��L	��ydWV\E�R�f�����f7�	�91 J�LM)���t;!=<����]C�¬o�^^.V��[���1��:��_��:*�)�L��a�ӻ��g:�,�����/���Cpؤ��uF���:��/�Ax�5��x�U��h�%ц-�O���$ۊI�s͝8���y�Ao�<˶��v��*��X[|��w�;J[q1:n�3���t6R��Q k��;UI+6)Yݺ��o�M���U{p �ϴ\6+]O=�|8~c���`?�����r�_�%�sӛ\ּ��}oC��>�����&-o~Z���x:C�r7 �2��I���
�v��d㸥B�7Z�iLhş:�4�7(h�yS�J8� 9��
�zWJ�K�](z�[��V�P�\�mM���^���ӗ��G��Pg�g��� ����Q�00�K���%�gsk;�o_�!��P���
�U|�Jf��!��pܾ7���|lB����3k!��4/�طC�q��U�LTƀ)EVJ��.6y,��|w"�-廆)h�UIX�L�Y�J�ʔ�;��.1̀�;ک*R�*�ho&T�9�-1(p��{�8��[N��*��ԕq�<1�A��~R��b<i�ob�2�=��Q=�.�����Uɥ�\�����{�f�oT�fXZh����E�C,t+6>���U��9�gl��.���	��c�c'K�U�|�j�S8˓����ol�� 4��G�Q�+�^Y���齆�Z��>O�t�|�m`���X����y�v1��D�Ҏ���h�a�IuZ�K�rf��i��v�lX�f�ķD͠�3&�\�:,뽈'5�R{�6�̖-&ח$vok��wQ|0��Rw��\� �)�g__� U�\6��v�p�}��9��k��:���Y;�p2��T:�*v�2�ύ��=Fa� g�X��&��n�B�RtJqW�5<�����Qhb�B�Hs��f,��º���1!��l[^k�7���.[㶝ϮU�f�UZ�au��k���PxJԏEOL��˯�OK�/��Umѿ}�F��=[��ǵ�/,��YH?���)X� �����,S�M�]̾С�V(�7���B��q�*9ĝ1��u�����g�������̧Rk��A����	�ɾ�	�'��ь��K�{�O>�X�����+%#�B���f1_׽./�5����ngeL=�V��[E�ߌ��ghdRck�P�}�7�ss`�����Z�j��>H�c�#.yem��9���� �3.�����yS�݄o�|c*�?-n49n6�f��}�p]`��<yJn ��	��\!(s�W���c�ާ�%�74�;��v�+y}���1�5�"<ky��W5U�~t"�`O�i}���κa�Z0="X��Û�{�i�076�`Ϸ�V�
�g�Cn��\���$VD�u��Tn:M>Fԗ@WR� K��^����gO�-"0���z�#ΞY��AM凍 �=9�Y���K%���ί��܉������-H�`[�C��os�>K&j�2�mr�-�|���m��H�2��t�s(`���)y9U���򨻒eœ#x˜rT�
V%�*�,	n'��a����h��	x���(i���nd�o�97���u1p���q���ft�7	�p�1��v<�*�R��`�pO��MT+��|��\k:���&�Ƌ㲰��a�ݛd4c�Lt)�eK
[tz���@(����^�����х�F��sd��v�H�R��@�01�	d�*
t��\�ๅ׼.�gpNS�Pd��^�:���XSu�j�?+E�!�F�:AC"7����,���cή�í���+g@�nj�ѱ���(�����W�Y\V{|�+��+�+�V�TB��S!����s�<o�,)��ɣ��L!���������4\�l�D�Q���ucũ�ʡ&e��Y�_S�]�� >��mW�upU&0C��������#w�Ct>�{|�j�W��aٕz�j���\�V���ٞs;�٭`�"��l+�_��e{-X/=j�wZE}&��X.��*k��BƁ�]��bC ���|��S\��tM&��o$-������r+�z�T0����{��㌒�G�XS�ͣ����z�%�E�.�\'b�=�����gm��
��X$*���L;�+ڐ��u��Aᎆp*��s���9и�9c���p:�usg>R��6�AZMv����q+��s�.gx��O�ږ��
^�L���z���8��/�]�>���h�����ϓ��V�� �v�X�s�~zR8\��H�XZ���#Z_5E��]0��u`��F+׈Ώ>y[0O]R�}����;ѫ�|�"@=�A}�u,)���׬r���c��7,EB�v����.�"�|_Pr"�Eċ��.�*���sK"�t1��Ì,uAc���c
���_`zׅz^G���/����7�"��kn_x��� ��$�t���6|����:�k�Q
a��'��N�4ДbT�d�oSh�ܘ��u��vUH�4>9�+�e�
�;������ώ�����#���L���t/�C��z��tC��T��>��Do�];
�>ךp�c2�D��Kq�o�\mI���S�5k8�;\ �0��X)� �7:��ܩ!��l�K�7;�r�*��螁7~ڰҼ9��S�s\�����-M���^\���vj��e1��&��\7�wA�0X�>�ICq�gl{�L��;VPEY͏��f�
�s��q���E�2�6Wr�/��Q|�{�O��땔�����fï�Z9ZD��؋��2�i�~�o��'3�AMF��
b5��>N@|n%�+਀g�9=�݁.�2�~F֗^s5�����{��bz��ܴiI��Q
�}?gLc��8v��ع��m���/�˧7�(VE�M��kѪ	�jY�QX�O9`*�u�Ҽ&s��f�=WⰧ��l׭4߽n�=%���^��$|��ʍ^�,`�5�X�[(	�@��{l�j���I���7��q�i�*Q���Cׂ�\'���*�g%R����[<����}��
S9��)�j������_1�&�fMz9W�}��6����U9n0���v�̾�qo���3XTE���X��Uc�\)`��Þ�`TY�s�a�nPѮ���Ŵ�	U�X�v�n�U3Ҹ��~+%3���IRT�Y�?X�].4�J��)�ƙ��ˏ��,�9"Q蕔�-�\놫�8�S�Z��q��Y�9:��1��V��X�L��G�8��U�a���K�{o�� �~��	2*� 3<݀���=[��������.��h��p��>S/���2�w�,KW<h�Gn�Lnq�b��%W]�b��O�=���>T�y'�����}�r�H�p��iޖ�uˮh�y�Rgh����#�wJMG�Kr�V�Ǩ�Nb��/N!,���.[�Cs> �O���>�82ƫ�
�aVtw`�����u"�]��u[&غ��w�.m���q�~m��.Jh]��I.���w�_*Y"��(E(�v����A���m�,�g���vP��ԟa�����#ߎm�ӚR�K��j�=��u%��G%>w���u�BCYι�1�6dM��P����{y�R����O�{==F`��Y��
b>e�.���A�qך렬�ۮ�A+];��;��&nP��#��8�U�`�-�J���-�Ǡ�d�ܛHZm]��[����[T�o��:/ѡ^�%�`{�w��dMQ&n�����3WM�y7
�t���[q労bN�̧Cz(��N��e����V�@�t9[��f��)�Vb��t
m<�ĥ�oΫ��k�}�lpp�>bԹ�6d�n�:���$���Y���m���f��j����{���v�f3m����W]�1��&��sփ���`:,Z�)OGfw���Ǹl�&n����t�V!�*��dhe�AY��,P�/7��fg9A��Y�VQ�ǽ$���A��o�J�R�=����h���Y�'\�z��d5߈�('�+�H
�U<�R��`&��q�1��ك��S�7V������$�	���7 �Mp3����L��u�堎�;��J�uhd\e���W������U��:�J�+E��&c�WhV�:������k�t��z.ɢ���m�RW�����.<]�:��jG�ۥ �]E^�SƟhm���w��g%W��n�۰����*�ph�� ڗ׽���9SH�W2��OW\���v[�ԯ��ΰ{�n�;~ŢE�M�8_j�u�][�G���H�S���f��psb*ʚ�2a�ܲj�P��X346@���&�3s:��S�A��-�8��7sO-�����y1��iM�\:�*B�z�r��y�1F�D���{�������RH�D��ܮ�Ύ3$$�iIH�3j[-�$�}���w�bT��e9���1�ҝ4�ᘣ$d�N��;�_�ev����Ƿ��`_M��q���e�36��È+�� ���� c>��+S����̻af������l��.���mCG�`�ϭ(zꔙ����Cc��S���a�������-4�g
2훥��|+���Q(��N�1�8�j^L�|���1�ˎ��u��p�5��]N��/��ze�˓�x]45Y䦻�ǫ�{&'ع�2��Uw�����{0��T����H� �YsG<�zà�6BsV�᫃�>�����Wv�*wm5��\�����M�}%�s5�*G�ٓbGIڶ{V{ޮ)�Ix���3ݻPG��*t�)'ܼ�ޫ$Ѥo!{V'^�c�����R����;r�믿z��_cXv1�
�j��j��A��0[(�kJM�)b�-��H`��h��X�""
�46�JSKF�l�EV��Tj�4�DE֨֍:�V� h+Zh�6�Mh4�;b��%4
��PQ3r�D�U40E�-h�4[h���E&����
�A˛1�&�c4h5�Alѭh-�l:�N��!@r72h�hţ4Pѹ���DESATTA�ht�m���b�$6���5Ȉ��N+b��P:�4j h��Mlj��(9��BضD�(�End܍�Ӥ�h��i�*�֥6�T�5�AȤb)b)8N�A�h��N�b�F��	�v�T	QP�GEUt4ĺ4&66ƴ�4���R��HRk1�M�*�X�5;:*�"����j��V����"y&�i}�{��`q/*YVOu�	��>Ӱ}l�c��7z�P�'���@�^����<d���}*��9��w���?�)�����u�K�c�J����y<���x_���?G���Q�>Z��O�w�A��*�h�~}�w	y���n�C�<�"�:����H��JW���7���'��D�+;�C"0D�#�?h�O�wg���sԺ{���On����M���r.T��+�O#�uu!�Hk��u����'���C��9>A���}�]BU��z���Ͻs����깦���M�g�3�B#�b=��O��y/�޹�;��9CﻸK����΀�A��<�]&��!�4��{Ǹ9������/PPy�~<��5HRuy?e�y|����(s��s���O�b����+��\�9���C�����>F��*���~���!ߞw�p� ��N_O|��Gr�������{��_��q꧐�t��A�ב�^c�^�� =�ۮ֧"�3��Y����,}#���o����*B�����$�/���y����g���)�O<�^���:����t�C��<��y���Zc�o~t�h������{��� �|��f᭣[�ݞ��e�8��G�4~�N���	_�����:�>s���u/#����v���`��~���ܐ�C����ܚ��	O�=��nT=��z�B�}!?���`�����;B��Sx�z8	Z�/߿��9I���A��O�� ���|���C���>G�9	^_�:��e����u�4r����i=�mu��5O�>���"��@P��L�����u�h;��˹~��SԺ
#zy��ד�HS���s�?��ܟ���w���?�����S�?n_>��?Gp�O�>�!����/$�A��##���b��>"�Í�&BB���������C��A�ߞ����?������`�Q��y�� >Ǝ�}��ז���>y���r_�*^�޸u ���c�ξ���}��ܝ���@>��
����)���a�fj����+�}���~ꐈ|��/O�/������;�ѥ��=���`��'����?I����z`�	]��޾����:_�w������/?{�@h����GǬ���4����g���_�{��%��X���*y������������diP��(�`�u2	b��/zs�(k#=|P+j�/��Q%S�Mn�Ti��ˤ�7嶛&*�Fڶ�w)�}K�ւ�A��f��<9�٢��A�?��oTB������Nl�Y��k���zs���C�~���u������y/Q��r���^BW�}���������;�� �:�!�9~�<�O�?��{����%/���=A������z��D���}"����Tx��*�Ǯ�y�������~A��'P��t�������|܄�������z����B�|���������)���p��Gӳ�3$�������ٞJ�[PO��J���.����A{�]��r|����{��]=����<��4|����!�w�uP����?c�0}��F����}���O��GQ���H����'�u�թ��9���:��C�_e��Ͻ<�h:�^�>�����)��������9~w��!����Z�����X�<����On��|���~JO�o��`�8x��%��^w�"v�Ƚ�����N�|�I��tu�:���{�������|}��bw�i���Η�y�9��s�N��˨�z���.��*����%|���#��%i:�W��>���1����[��t����)��J~��<�_���������{���K���_�h)����>��u�4v|��^K����}��'q�4>G{����̇/�� ����u/�>���!U#�/Qdy{�4���2�矹��#��^��P��������!�I�rߘ����� �s��C�G$>y�:����h�}��uiG ��}��I������}=ϗP��;>��#�G�}]�^<�s������s�w�]P��_#���'pr@u�����O�u��_c����ɥ��{'��~���}����_�c�J��t~�����u�p��.��G����Ꝙ�&]{�l�}�޼���@h���|]u?��9&�:9	I�>�g��y!.��~������ܞGP{�G���@y�vs�M�k��8~����Oӎ|#��x!B>���t_�uyQ��8}߷��B��ѡ����ΨJ����O��|��?����`��I�N����	O�~����`�r���{=A�:��}�^I��g�?'�w�j>�Q�}�b�n+%��L{۽s�����1�:��A%n��Ζ1��p�M�_W`QP�[�kN�x+�V8嫧�&������SL�W��ⱞSU�B��xry ʠ^+�f]����Y�W-V���fޝ��v��j��@ZΎQu^�A `��#�}�TE��I�?��9�}à���w���t���n��O*O9��}�e����CA�nG����;���쟮��:�K��<�~Ƈ�ny���}w�ރ��ڜ�z���� ��p����1�� ?F���:����<����F�N����އ�;���/>q4up����K�i�'o^����修_zﮐ��}��p|��(��aq%LÒ'�p�������f:��<ܟ%��yuG�����u{=�W����:���y 4o��t��s��#����9	T���9�����l����we� �"!�����'�2��}��^��B �4G��~�B����������_>��z�׷PC��ti??����BU����^��=��+_`:���yI����?��%=��u��A�>��@��Lߌ���Q��Ws��􏈃�}����y��)�}�%��ߘ�;���c_�=��������Ri5�̟�;��t������/$4�u��8�����<���<��A���{��X����l�En���\�W��������C��9	Gϼ��yr#�rOz�ʗ�h��Y���8A�u' <�?_��N���<����K�T���<�C�����ݞ�}�?!��>Q����шS̞�HWk� �⓹��}��pF��~>���B�����ޗ���CA����C��{�K�u�O�w�y\���B#�x?^�p��`��� �:�ԇ�!��D�����B+�i��X�m�D��%Q���'#��r�{���d�O�_~p���C�:����}��}�r:�
�}�;�K��@|y�;��t�<����xO�th��@� >������k��������B>GP��ܐ���A�u�g���S�Q���>G ?����t����ބ��h)��~���y�?p:!��=�>���f����z��9;�;[~䋾W�bG8���+蹆1xP�,`m:H�h*\sO�'��C��]�M�j��k?�,/&�g���X����F�mh�\`+�����|B�'Z5�	�+��9���^����v �(��[Y�є68H˼7Ef�\��S4ɓ���@��Wz���ӝF��H�kRk��6��;��Ȕ���FaSȷsy�i9���:t������$�iw�ٿ�*��Huvu��7<T�ro��0��̋��pn-�_��nj�Al�d��K*�@%q��Pu�t�.WS�v��ÝΚ������@���5�,�"��Uu�GܥDo�_�¥O���a��E��|�n�e>�慍���]xΓ��5�)@�^X�ԁFY�!�z��^��њ�1���g,����)�NB�k2*��"��:w�͞N@|K�{�́�k���1�V	AC���㊔��E�u[-~���������yH�����Wbqg�Cu\&�j������<4��(�[�*����9{L�ه]1�b���V��g%��Z�TEB�s�m���(��y�N�z���F3`e�'�Q9P�YzP��b� �l�'S���O �\9����~���QQ��5���6]��w��^�q�{�GG�������]�s����o�He���!B�|���v�ӵ�Cw�)��-�{��9n0���	�}h�߸�^xx�`>�i]x��ƚ9�N���BZ��3��b(G*�:%/l�j�j�k���飑v�*ܦ� ��E�]��Tp��_-��O_���IX�y�cM��8�qrg��Y{h��6�ɠ��`=��i����9�)^U�q��'�ro_	����y�PSD��7'u�E��2�E�ф-�:�8�7(h�s0�v��͈~�w~GO��6�������׻qN!L���|���Jİ��r�\i��Ѝ񌸄�=q���M-������m-�p�h��f���_�3ꯕi����!�㌽*R��Ƀ�1�2������m�wdH��H>�W�0;R�]5\ zwǞ�>����Bt?s��"Ӈ|�yi��<�`��� )�^d1�^\@�	ʀ�j�X��J���Ʌ�1�
m�BLԴ�t[�A[�P�Um�.��z�F�(�N\�ta<a@��-�U�w�s�R;��ĭpPֻxnf�h����-p�5�������"y�eY��٠o�g��ܼj%dW��=ckR���;�	Xk�W�
v��S8˓��ho(���T+� \w��>g��"T-[+/dO+�HC�˒!���N�n@(e}�.�*wS�?6J5�l��5�m��������@�V�^��r�Տ:��c���S'�!�W'A��fМ�l<�\#.&�K�9�[���0[8�4|K�g{n���z�Z��
��״**�'�$I�a7�yۃR�\�O���>Ko&��ލމ-ٞ+-2����)��y���Ȗ����O�w1����-;R�8��Ic(/�E����/���I@o�+Y���t���jY��U�����p�[�E�)f����]ѻ��p�3NY*D�$Cџ��<iV{n~�{\���iX�~C�J3�]l�Q�v5tmU���b��������������N��f+He�m��LV�eZ�խ(Y=*\B1�i�\�	��1��~���;��:#D��ی;U�V����4��DC��xe�N�C8/U,���hS�c�-/�^��Iʣ/�y����(�ɶ������Tmo.�}u �v�Vg�:Y[hU��7�/��2#{��?^)l�|m�ƹ��� �<�Z���ɺ������`!���	��P�a
%kiaB�g֭��{����a�lr����Y��;�8Y0��_)�5U�>_J�w07��
����-�ԩ���-{�xcڒ�A��cwa�*^\!���w�0[�%��TI�BF-mM�VK��T��������>��j/����'I��Dr7�8�nա��*W��!#pH�����������#Ebw��B���\o�(���3���V��8yuy!��ǛFx�\̭%$�ހ�r�t�����q|���2gyK�x��55�{�7;Y�P�$�5W_jJ=L�`h��Y���Q���"K��&T��t��W94c����}w�}]�洈�\b�F���K�__uB�3��G8�_ތ��o���]5WOSw]M�;�� �xu��%=U��<��_�=�C�U֦2	��M�1&�4㜤o�վjrffʒt%�'쯺l���mD��R��/~0�1�f������C�)�
��F俤��:ѯ�~Y��=�j��u�'��hݞ勄��VN)K�uZ3��D�RB�7@>�*�k8M�&9��Y�c�V�#sj�ӓm��M�m$OB�`������e��2Q����	�`ym7�ba��aa2a��&U%[�ͫ����$�뜳��K���b�|��^*ej d$�Q�'���5�&0OB�����}�s9t�\d��Qs���9��~UQ=O�E�KՕ�N�nr�t�1u������f�R��e*�}��U�S�}+o��@
�Sa�7=���Yw9�J��ϟ#.*�28R�!�m�\Eb::%~2����bC��#��r2Ϲ�"���Đ{/��y5G���-&�,�QV_!fkCS-�ܙX���9:�	��W~����,��kw��Mל����2f��ϪD��6ΩE�rt�>���c�m�kv�)}ݘi���<�]����u�ylڹg��O����=�.�8s9V[��m���U~��m�s/���v'�y�J����,�UXⶳo$u7���#ng��f�L�d;�8\B���Y	QՎ���g����|�$��M��n���\CW=��Bno�YP�r�� h�;M�ܱ�w#c�i]$D��hd�g_�yk�%���m�c�U����0��X��!S��c������	mT6$�����Ȼk��cYy5�x?�������$�%�;f�*�xn���:�^�Y��=����ˌջ��u��]�q�Zb)�raF�荘��*�D���WˀPu}[%	�)����V  r�8�2�/w8΃��
��Ag��}����A`��U�g��[�+֔�tC�	��h]�:�Q�f����ۢxT7�h����
 ���5���
�>>xd���V��m�����Mj�.�+�'�Ø��yXqs�8'�@��t�}7LF�h��s��<��Y�vq���-���1��5"~�0��p����9@I�0ԩ̆3���t�̬"�2��MKSq�`n[�|��(�JZ�mP�$�D5k�y�.U�&��R�Pch�{S�a;P����#���y���!�w������L�;K�ݷՈSE[ u,�,'�2��u������� .��h�bV������Ȉ�]��&|3�b��Ec�w��:�ǅ?��ŝv�l�W��O�o�a�)O����`�Yҷِe��OE��y5��h%\/�}���|�(��pS���FԸZ����N�dQ՘t�ޣ�^���Y��6@�ہ}��+*mQ�u����n�b�p��H����\�]d����z��Z"~|��XϷD��u\sR�gR:+ũ�8�����g�Dt�\��@h���2�;�L!�!�٦��4_���ڔb��3���9�{&���|�\��ڸW�:~���#zd%Ieٽn���~�0�w�m\[�2��Ð�C�冮�me|\Om1�h	��E\�(a1����V�L��d3�n�ǵ�e�ݡyw���.bn��{0�mBb��z@[�X�� Mt�*�6����p��J��8��y��J�SkǡNк�l�Hڇ����W�l����R�`?��������ʳ�eZRBr0h=��ZbP�p�H�Cϒ������f��P�w��S�ǃ)]7]��X�;��S����ox��)_���G&*��U�ÌZ��Ɂ���s��S�y|W�)�;���x!j�/�H=ܩn���nk�8����Q�v"�5�6��<�G'
���i�C�������ϵ'բ�(��O���>���1X-57�No�}�c����L�f�ʭ��4E:�89*�p�2�}�!�����뱋���J�U����Y8�`<���%����)��rW��o�<`l�{!y� 	�� W�/�~��]]�{Զ投qZ;��Ý �= �ϖ�x�7�~|j%J��of������s$pE���V�]�}W�Ā��b�\�G]r��X�|1��4J:C��Tb����y�ķ�I�Yu4,������+��=D��雯�d�W0��ڧA���A�ڪ�`p����R�m�PwE����Yd��!^�Z_γԎ�)y�9:�2�ٿiX�������Cʖ[��n.!W & O������,]��7�N��Dm�J�l�<3h{FE6�Ƨc�U&��1T��c���_hb�	O�6ͳo*4TG<����`�Ҕװ�)��u��0S���eG�lV�y^�S�VGOg�uY�b�����!�� 垊�ƺ�gIn�뎟+�ey۰v�v��%|eU��+#�Dm}��?\cT���"�NԼ
�j�.��z�59�z#��bi!�u���_Z��NpO^�
���߭�Q�XC[�$^3��0E+�]Y@�w@r��hZ��)T@��}�U]j\.�,��^���fذ�}��<<{v�髷�=�z���i�2���������9\<Ƕ©��HmH:\�x��P�4��rí�a��4+&��+7�zh��I�k[)f�Q	,+m�]wB�b�K��WZ�\���X-�8�Q$u��R����!���À6.�ڮ�&h��9�,˗v�,:z�9ܮ؜��cd�E�AC[��-',�q8�,Y�#5��kc�gV���Ź\����J��#A�~Kaxj�_vnOm��4����pyH}.�u��	�O�`0+����gH�X�3���4�5g�����'m�^�eDc�����@�F�a��j��;v;�ەX���26���]�X)��P׭����R�c*Po�#|�S��w��3O&�
��l#8��mc�'7Q3|J���Y�eS����n�	5Ɠ��.��)='X�ԉt�<��r��ssn���bK�8�/'w[�\�/���HЦ�XXk*�v���J6��.�5����"�����pQ3���g�Ӿ�rIӅ��| ����E�������xq�ci�5[�"
����=�B(��5j��̮dY��dq�����lV�>1�9���]l�F�C�u#�J�_gv,�.�U��:7�gCI:1d���%����@hv�#u�\ �}x/�]�Hf�xa:cc&���Y}���`G[�쵂Ԛ��:KR�����46��ڳ�G~z�b���2B܋&���lXZ���Zk���ܺ�K�����n3Ǹ��"��U��7����;��]��g;لh�P1�8�zt9&���ME�$�*ݤ4�9��w4|�8Q����/ 0��&'i�Wr�ܷ��w!ys�d\��oP�4u��y6ӂ{�u�8�-���Q���_�6N�v�K�G;��m�"�u��h$&��S�e�Ntԩ���NX2)t�pS���оG�$`��,m)�b��R��xctR�מc�Vvoo�l�`��q�w�`&����@��jʕ~��f�p�tA�{zA��!Xz��K�k�ut)Q�Pp��J<]3jWVW��h���LcgpҨ3ד�vT؝587/T�3Fh륍�cX��7:�Y�C�D�B��7z����͌��JX���iqb�t8��;}�3yOLu"��;�,@,-`C�w%��Hr�c����\���e��fw-T)Lߍ�ԟ^��&��b�Az�\���ɏp{��/iY����8�,��Q��M&t�l7�5��p3e)�_i<�:-��7�������؍+�������<ԆZ�9�W����d�R03�k����˗�*��Ԩ^��ޡ��\a� ��9ugT*���YVj�3���i=ʞ�̢۠����u5d@S�
u�kN )i(�!4��*X��[b�AN��(���5HP��"6�S��hѪ��5@Pm�4���F�MP��@�i�KM4�K�h��4j��(�:V�
�����M%a�1Q͋j(6�"��(*�&�i���Ѷq�QM1R���QO6bngA�K#���j��C�h�`�e(��)m�اF� (�i�N ���%v�Z(Д�Q�������"���t�h�m��J�����TD�PQ�3V�4P�Pl�II�F��v�bm��!�
�����ѶJ"
�@��-Z�Z��j-��G@SBW#E�4�<�H�k[�[� �$��iH��]]m��ij�&��|�G�N�W.-��;1mL�t�Ľ�ہ���.�#F��GI��'�lw�?v�<�A{���٩��Mr+�����諭6��tz��۳E����E����U���)T�UT�(\d�!W2�=�e��#�������Nf���I��E�P��G&U���/��\��'��@���yo�U�R*���M�=�p�Ʉ����K���bn"z�*�\̻�F�|b����γ�L���,!W�륥VmCF��k�J��[$G2.�Ç\�!��CeDo�6�N�Ay�Ճ�{=��䀐��B���j
�2U�iu;�:_Nc�!q�F�c�#cTY�z��I���}yS�x3�a��	�"�Ș�S`����1p!=�d4zT�$�x���qxWvY�aj�C�����c�<V��0���ྷ�	�ة���p2�0�1G�0��ͪ,������P&+;8��TND��9��2)S7�O�9Y��4��o�`�C������P�V���r5CJ�!p1B�9�r����`0ۊ�b�c��5V�ͨYØӁ�����Ф
�;ݏ0{�)��&��27��60JuL<�hٿމ�2�}^L����J"��C���EA���n�ܭ�?ACO����*��T���d�P�ȷR��u�\��2���n��Bq7�:39��y�o(�il|�$�W�w��O(3aU!�������� �g]�h�\�Ԏ��\?>�7KA�	_`ý�nLsM.����F�c�}��}Dv��e:�<c��:��ǯ����O=�����/��*2g醖\���w�����{�-b^�K�MA�<-�z.U���QXvf)���%UDwn`l.��un1}f���������ȡ�M�pܑ�n\�֫��Y�<i�@_JƇ�}{8�XP�5̘��٭���37j�vCyhu�3Ɯ��}��F��iWicY�	��r.��OQ4��v��s�c+��W�\��}ǘ_?{j[[�V�O3�O�n��Er�ӝI�E�vԞ^�Jg�����<,t���gc��3�;�8ZW�8l'��l�*��)��y��M!4^s����{�ޫ(}�Q����ʅp9RӐ4C�ۖ"�M;a�8G�G�U�h�:y{Wl����u`b�7&H�=L
��84cŌ�i<lƬT�����`����uO7�̵&���OI�E�}�����0���t�	-p����q�i�Z�(�q�s�-
ʜ���:̳�rc�ѿ�bx.Ϣ�DL��Wˈ?Dd5syȬ�fک�&���k����z_%�BIar�.�4�:�92�u�oT��� �^����������cSc4�����OU�b]��Sza��^"�&OT�sP��/�m^6�ݹ�H���ۻ�����q�(uԙ�MN���꯾�����(^�������t}��A�:�[YP�S̖���#}���T�TI{�r]r��{�C]�`��c�>�i�i�7�C P�Xj��D!���?�&+��
��Z�r�����GH�Vk,�4D� V�$&o0;M��`S����#�����ܮST��\��j7N�W�;G��G1�g[�T�x>�ϗ�Q����j�C��*w(�u�s�{��:�+9V�? �{��ň�)\�b*5΃5��,~��*��uY�^�c�!��5�OgS"��Ɍ~��f�������[�,=(t���,AҀɬ��Bu��Қ����F�W�@i��tƅP�/��a��Y[�|ѳ��\6+g���c�����U[xz1�-Gh ,}Z ��}@P�m��N�CW<(k��rʝ:�p!2h�u�Ⱦ�*��W&Oq֎��f r7 �2�W<���ۨZy�4c��;�jB"���G[Xn'n��X�tX-(�v��V���o-¸�%�f�nS:2�Ɗ�7�2����f��>n��[��*���×hm��4��ҲA�ٝժ�R��o� ݾ;0T�;]E]f�&Nd��a�[|����������g�0�}��T43��U3\K���32o}:��t�3F�;�����:�e�f���SWڿ�����>�ʔ䮒�NL	+�H�?��yHA��`*k4�Q{O	UiV�,��o���|���ha�OX�l��ٞ���w��+��h�#j��K�eV1S ���rwU��'�c��}���uu�96��ZW�ѳ��s�w>,�ݼ�2 �_�$h�P�UH�_D�@X���Qp6�wy��+����#���B,gκ�
���Bρ�������2.&��'�D�H�zY���������}���0�T6n�h=����*-�P��$W:,��B���fb���j�*('��Ǚ��Wӑ�5�>��W\!�gY�-;��$+s6����[���E~�ӊQ՜��۪R����H�v��R��D�Tu
�IS>�C����v��$�r#|H���j߇�׽�W5Z2U%uڨ;"��6�ׅm1�P`ja��jt�tngP�trU��o5a��.~Ҷ�n��QR=���'�V+�,�1����_*��漓Z������Ɔ
j��,����D1�X���<ke��f�ǵ�s}�h�M$e��V��y�,�J;�K�Ck�{��m�rQ}$�'.�p�0�q'B�˔0_�/u�L�k��Ʋ6�#(W��n�:��ؕ�)�:�jƏGo��]𜣹6y�;r�N����r��-�9�������͏ަOD��>��>����N��h��\vvx�Yb����.�'��+vh\7:4Z�:b���1���ĽV��ǁu,A8��p�%V���kJ���*h�l�J��_-�qWpF���b�Q��os��C,���cG�q;=*��*�g!�*4����ғ����+{�K�r�3Q��e��UT���6:!��(��5�j����_i{O_ڐ�yͳ��6��i��FQ�y=�خ�Y�k�������{"����*��N<�p�2�o�2�6�u��3?L�r�Ƽ�O�΢���у_za|��Q
��!�M�1��Sr�!m�O�R�MޝF�/V54��{��WL�{��^ҝ�ŕQ��h�7s�}hp�u�\��V|��̠�_K���:���U�n�]����Y�G5J���H���_T$�#�>�+xʿx<���>>�Htot�=��q���q��)�Qe�H	��?/�B�td�5�j���cpx�iQ������ y�D��ng/z��. �0��nEV?R�c�S�b� �gC߹����:���effp�Ǭ!N���w2�q���s};���
�J�W����<��?4hأ�g9;QD�_9!�ϥ��13��u�����Y�޷����>�eb�e�P�xR�*��c6]�8wq���L���H�;�����}�B'ov;�Ok*f��~�_���ꯪ�Lc�^�J�g���UZ��%�Z~d@��ྷ�O�R|�32���7X��Y�-0�"Co�ٕ�C�S�F����*|�e	Z����ZMsx@��`�z6��w4��j�z���B&^V�<#Q��������`e�F�7:V�fV!73Տ�v􆗫���b��ŕ���g�d�Ne�
���މ�2r

�'yo��f��j�d�T;K���2�2�����33�#�n3��3�J1�������a���M���Ql�!`�0O|��\��xW:�ó>�C<�i�uTD�u=s�e�=U�����G�{�Z�^9f���4��gԼ���\���~Të���h{-����藍��#�Gu3uZ {�ct�g�Y|;dp���>ܥu �!U�d�º5]��)���MOP��Pѹ��oNj�c/-�]��'a���*{�#G�������A��I��㖸��[#����j.eG:g�ųm�f;!�1����w=˨~^�{�CmSՋW�e�hR�t���k5�s����][v�;��n�
�ŗ�O��-��Wfd�L�K�z�H�;4@��o�'���Ŷ/��[�s/���Ek@��r��:�5�oZ˂�e�z��P�uq`�$�S��2�. �=�l7��E��UW�}����[����6Ө���sq�*�<�i\a�ҙb�v��ն����!�=�ޣ�:�a�Er�1����hc\�h��xh��v��������#)�g.��^�S_!�Ղ�(z?3��8q�9�Y>I�.g���L1w�JQ{_*A%���L���	D�mo�;�Y�b%:�F;>[8`�K���N���%q��_W/'�E)��ǀ�9-��u��h=p��
�1�A��1�jvI�pخ���j�>�ݳ�В煽su�ƌˁ1�'P�*ڴQ�b
<0�����f�i��G���S��Bqj�U���5�i|p��<@�1��l�'@4K�6�܌�J�/����|��C;=�k�8��°@������/aN�)<<<�t�<j��L�]#8\Έ�싇L8z��f�U�a�_"���D��*�1�/
��EF��f�)1��%�*�KPc*y�w=�ДxW��Z�N�c�vY�R���#���XzP�'F)b�v�ڴ�3��E���t�d7uc�Ξ�ۺl��i��#iV�j<w��^2����5E^��^}k�ӡR��ZA��q�ޡ&���f[o�`��+|�w�P�2���Rܫ#���nCuw.�{��;I�,WN�C��]�v�oo�s�M�iO;���=]��*��2�l�d������˝L��p3�:]��f �M!�{��[�/t�y�g'Ա��U�Y�����5'x�}\�Z=n��ݮ E�2 r6��Cw�)��-���a��:�zI�R�F4�W5oE��9�e;���3Q���o�CZ��h����ҡ�4c�7]�б��y�[�s�LJ �o�,?:�k��}�BD2�y���-�p*�����ȹ}����(ѫ�q�U���ʥ��Q�0&�x����C	��U|�L�pf�)�Ԟ�f�y�y:�/W>aϫ�v�每Ҷ*�Y;��˘�M�� %=[�����T��{:`^[yϓ{ù���kݿ������0ݫ�2aW�=ʀ�d���@��D<����L�s��H��F������w�1(p�{$`��L������%���[6�Gz�O��>�������A}@N'�z�sEB���nt΀B&���$lK3�o%����Ð�QGC��&ۃc�����%a���}Jv��L�.K��:�H�͡�-J����ݾ�����`K����j,���J=��{�>�PBD��t2�˴tW!4�X�fFt]���9:)�9�8���;��/R�ٽZi<O_��k���Ɩ]�b�L��C\2���s�^��>�����T��u;h��T �ϥe��\�v��R��@(eDu
�K�����]��������n_B��z~�>�WA:�0���%sU�"PW\�V�6L!a�Z`�P2�uli|;'���'��2b�t�*bÅS ds�k��g�EY���q������Z�V��rV�A�1c��l!{3h�<�'����xC���"<d^cNE���X�m8�8"3.�y�)�[����R�o���$K,%3����g0Ȩn@�_s�:aj�k���n�du�NΑ�\��r�䮕k����_��/����2/�?p��E��biD��\6�\]P�KnC�p��BFl��:�/T�1Q��� T_RNU��VM\������T6��>�<x!�7�+슦6�V�Ypt�=@.�nr�ֱ�����-��Y���󆑥�v�ꌸMvR?f��%H�M��u�����u{������Y;T��M��,�f��M�)�S��]�v�YT��Ł-V�S��t�
 �R�R�^S�����t s�l��A��!v5����\��h�[���E+٘i���ڼq>S�>-l �XhĜ��/��b���5�b�]N3zޞp�n�O�����>w��	��^�� {���+P��v]i&m?�W�}}UvO9[���~������U�wZ��n�ڇ���Е��诤d�a�5�Wj58�;0sbb�jo�]1[��&�����LS��'�BvE�罜��o3+g���`����Ϯ��x�����ܛ��4'K���^ܨ��:���X���t�CQc�ٰ~��.�ˁލ���S2��8Fz�ַ��[��\Z:ἅV�L+�1]!u}����nMb{���;;WˋO�m&���h�Z��8w�tsu>��Ls�{�����Kze�Jk�K8�g�j�N��Gk5Q������a\Ls�*l����*X!"�#�&x�=�TҸ/+�>���e��N�2�|
�ޚOA`�\�)B�o�l.�}���ά���E��b�3��Qӊ/���w��q���J��ểԸ۞�e�����|�Jŵ�1�ڠ�t�����'�Gml[�������+�p‽[Sr�$fsC����niД�8�^�;/tsCGac�!��z�=wؖ¨g,�/�|_Nf�
X�s�L���m��36!&ЏY�U�`.���W�,��J�yK))���8\A��oqoH���9"�q��u�M�ϖ;�������v��4*��7��޴rֽ+V�shc���KӘn�$m���V��Ĳ&9�m=��ɵu��U�w[�����$�yԚ/WZ�G[0�N�0��f��|[�@Y��q�h�z�P7����ƻ:p��'����IKvG�K�k��ҍ�fh�̹g�R�O;
�/WCZ\Ȋ��ӵG��� ���f�6��
�hZ��t��p`���O�H���l�X{۬-l��t�a�]b�j�^.}�݊Zn{�+�_Y�{-'T��m7�K���;p�S&��~���,fuɕe��[����'���N��Þ��t�
J��%�h�>i��N:>ǧ
���u�{1��2Զ
�[H\u�K�a[��1�Z�#WOk����٩�%��m��G�������i^9wǃ�o�5� j��f�E���eq����e����)dt��}�{R��gmL�9� �38ޝ�#��NU�Y��e6�i�6���Ά�!zZ�#��}Yq�U]���{^��T�w�o���1��`��ke%o�,O�T��]�[��=β:@}���K�`:��ܵ�,�y1�,��
��R]�G�r���cWL��X8E��b�t>��h+��4��*�Kנ@5(���m�L�4+��\�h9*���׃ǹ_I������k��#&�8{r*���I���A���w�E O�=�nVQݔ�2�,�[#Zsjn�l��r�j�1^��i�pX�t�j�@@��#�#{�ؗG�kB��m�c� e�L�����o���Kܙ~��*JcwVt�)S��f����ⲱ�g~h��.�]ۻ۶J|2�*�8K���B_:I��P�k���H>��Tƀ#����/�5)�¢��"�:I�W[�vU�v��� �@�G%��+m�U�v.U�I��m�r�%m�A�"����X�.�:aLNݝ��Wq6��M�k��?O~��>�8�GZs�>ɋ:S�J�J��#v��R(^��f_ 4#Nm�΂���y�w�zY���nF���r	�e�'Hk�Q���Dk�tE��0 �KE�;��5�G�C�7o�mh� r����֥L�7��;mӬC$�n�^+�W�2�ӗ�Q�'�`�48�k!�bщ)���,ىmǚ]jB�,�Y[(�w�+�6��е����wK�zx���	1�Q�0�/07�`jHߞ�қs��G�RV�wOojJ��2j�]5ܻ1�Py!�L�uc���ue4hB ������1��F�1l�F���"*�j����v��)T-	���i�hh����R�@U�(CCE-EJf�JJ��h�5��D�T�E	C��٧Z`��kAb�����I�(֚�b
im���41P�U&�H��Q�TEAKA�CI��m�l�1RP�[jB��)ŧI��Z�F�J��$%�HFƨ2�+J�P��Q-U!CBD�b���*)b))Jt�4klhBIT��Z��'F�и���`���X���A����������6�DR4:DIA��(
�W,�s]��\�쓮`�<=��Pk��[��������$p�,��`��ej�֓�L�������#�}��DD�U�;��5X�?G.p�j[�J�y��j8�O��˩r��Jd�C~p�1[�Cn�s֢b��&��6��c>���ygؕÜ�����{���s\���n�f�gT0��̬��7���QO6��ۍx{�1	T���U�%�}��+Uwd���/3*,�VW;��w��֛��֫]�r87{�Lr���y�Տ`�py�ۚ���XI�ڭT]�C��ޞWZ5�|�^�هz��2��zF���U�-��S(��jn1t�S�Դ��ə\ޜ���룵}
��f��T���D9n�u�����R������W���.����l���[j[Q�u���:�d���N\�W�T�~�/���*zU.��ө�wT�Nlŭ.��_�Bϛ�v*�0�kF��C�s��l�X���Cd�|*פּ�!�ka-�q�f��u|�V�xP�V������*.W[u�:��
p�h��2�KBv��/o;7����тx�A�����2{N-L���d	M�,�*��+v^8�5^��=�����* �=��ʰ�;iʻ���/�L��IJ4�|���V*
�=�f�D���e����b���V��=2?�}U_}V{�W[m�Cmz_m���vx�vu]��Bp�.�s�t��}3}��ch�����X�q��5��R�eT���L�������9�ڕ\_N;�u���E��3�2�o�x�^��b������ٷ���ۉ�Cb�gj!��^�0�����E����Eb'��zy��q�ws��(��.z&#����W�s&��kjy��청v���D��#ܤ�2}�~]K���/�>�����>��ߖ�����D)�h���5K���g4K�[�8��S�<��z���//����\$�j �նά��{�w�tC�~�$:��ֵQgE���;�MF�u�6�Р���b7��g,56�8s�v�V-Ʒ]���J��_w�y?'UZ�:�7���͗	��wݸm�)�W����0�n&���Mw5<���=��HWJ�\G��K�vgee�
6��sr�+)<r����6���`c=�/Xē�t���N�������^�F�^�i�y����b����QX)i�>��>\��̧F^1.���҉��{�{ޣ���x��r�\��2;Z]k:���x��ׯ�Q������V�����S���zIF���O��sq�T�����N�;�	���)ou�����˟E�5��ސ��>/FS�r�*��YB��jZR%_v�2.��M����.���T�[�s�_=�V�0���wֶ��'۵����йZ����U�S�����_d��QZ ����셨�5Q�^	����:B��lFX2�&���n�!Q��S�UB��@kcy�Me���Y�CX�g�/�W�x�ޙ�1c��ҝ�px3�ѫ�E�5���v��I8}eM�����_�n ͼ���`��v��6]�Š7���S���ħ��Ft��&6���aX��p:������Uf�H�k\:kAN33��5��Gl���\k��=̚���^9�`9y�� e���b���Qnr�c��Fr��yۋ]y�Q�޳ꊣe�1�C^���x��<��*P�8�r�S
꺗Ԛ?%�L��}پ��Y��וq�Nd|c��HPWk�b{��&���Q�����ݢ��}��dJ�������Y���6�j�^���"�嘜�t�Ut���� ���eC�r�.�!yulynf��LkA�a?��U4q�(��妺��ʇ�6�aJ���y7Ԫ�*�����5����]�g������"�϶[�km|���%R�H����UtGc��zM�:W���Sb�ŧ�]5�J3o���v�qNso=�K�%���;W���߱�ZWr��v'6ݎ��_V;ك[�^غk�S���q�`iZg�t����7裫��J=d��W)�����m�VJ�{�����xMy�B���]q&�>�����U
u�t�QW*��W.�{.�2(ͯP�+�=p<���؉Z���ˀ�wIn�j�J@�c[]�>���;��#�&�K4Tqf%�-\w/A�[�!���_[�/�U9��Hk�&u���O-�a8{g�k�zS��W�{rQO���r���1�� Q�k0X�.���>�R��ۗ����R�nr(m���20)�0"��I�#Y�9��~��ogj�*��.`+�t5`�� ����)���eN��yQth��h	u��A���X�rI&j�N^�r�z)_@��7�	��Op�bR���~�<��s��?}��}@��ya��C=e�x��g���k��|��p�sv%I�s�����M�f7���+��x؟.����RN�m��(q�4_-WǕ�/- ��
����K<g}�����F/�.6[�6�Q�|���Z��pg&�ӈ��5f.�e�TV�U>ұj�^�}Bi
����U��JsՋ���ӣ^�p��o����s'��/e.�+�=�uy*��MO�f�"w�v�X��B�G9w;	ꯚ�g�\��<��ۏ:$]Ƿܛ���YO�����qʾҲ�57���QO7g�3O�Hiu�wn{/,�՛<�Z�9��F��.U��Ue�=19���5�^���<��/|�o��3�83���/'~�+_jk��J�F��U��y�4�c�4a�O��sЦ�m�M⸀쭿��T��M�J+���]4�����չ�?ݮ0��-�@��B��f��w�G|[9�o���V�v��/aG)ٞf>��ևI�~v5vסw+A���/�(!�\{CH]F�"4��@��$�Gws�����	���JvNLU����wcj��=}�R�=�_}�}Q;5����M�/BC�o9��C��v�Q�.��o�49�g�s��*r����U�;Ro�ܸ&��<Ю1�Ӕcg���uf��R3ʊ��E�2;��s�Ǔ��:�.̄�1ơV7���v&ʘ����b�­jeN<��ح�6K���w��Fk��T���5��#�c�,�b��˽����g��f���ǡ�͌��"�,y�\���o3U��ٮ�����eL�nzV�r�UE�k'�d�C}�yW0�+�f_Wf�Nta�h���Π�yW��%�NGc���-��יV��ǵ�uR�*���]:x�bOj��y;�ԇ��v������u��u�eWoV���#)�i�}�|�v�~�9�r��mE<�K��7�;��|��k�x��V��j6X���Z�ۋ�	���7iu/k�,��Q5���7�P�����*��ި��"�{�)�T�{�(c�wNz��)�VH�R.��u6�.�U�\Ў��1�d�u��I:[(]�*�l ��˫�L��n����d�V����v����h�9
�Jޮ�m`S(y,D�٣�� �J��膀Ë��/��X}���~������~�������Ҳnq�Y�Q�9TwK���;��Kh������������'_�r|sT�`��n+Zȋ8��/��J�Kv&qSYӎ��&_<�{�4�;Q�����:=;�����i|����2>�k)��(]�<������k�c�nѪ�P,v�,e݇*"v%(J��V:�ys� �����}'eV���w���,�����R��*C��L��L�l�^5Ž�Z'��j��K��·zC�w�OSW�9F~N��Hj&Q�U�W[�VG[VA��"�>������ul)�ؽ���:���9t;TZ���f6��ƭ4
�|fB��^�S��7eN���G
�<��5�N�k���f3��"4]����]��_zS��4�eӚ�:u�q�i��8}pUÇ1p�3��A���\�Oa�)^�c���� �����ཤ{ ��������X�-*�B�ػ�,L����,�ٯ�p���j�(��<�����`َ��\��R]�Ô�.��6���W$�k��V��N���"�WfA]����D}����n�,���fe)8�?$�*m�Wݙ�#�m�B�5~�i菤���S�o�7bs�N�:B��M�;�+Z�u��y5w����	=��ѳ�j3Ż��U���bzkTqn�T�bc��$G"�����ͅ)�e
{�W�G`�Y��4�����QS�d��:.�hT�q=�z����G�>37�[�CO�e�g����׃+B'v��<靨-���ל��{���l~r��wb��//�dY��b��Z�q�� �M�{j5���ܖ��m�LwW؄�k�5��
��T[���v~9���Ue��j�J�[�}����T)X���ۈLJopU���&j��gc������͉�ʬ��kf��]�[����{�`��n�򷓣��Uɝ�P����J&�58��qW�4�孑R�k�N�lUסGts@��޷�������f��T\��R2���+��BF��Y������o�e��U��������W�>�(�X��峜��W����R\���7��L�a��G=n�<��vZ_\�3�}|�*�����啬o�yJs�T��0%_@��o�69�`\������V��aָ�ۘ��p��:��u`��)�v'�zU�j�`妅�זf[<�0��>�ż�������୎n�u�I����0�:�fW���-%�o�v)3�l�p�ӯ�Nt:���p���bU3�Hkw�n[8�Eu�%8���XT��رΫΐ�;Y��N_�N;
�e7wKpU�Σ��Ya�����>G�Eq^r��.�|�<X^���7���bV��~���:]q4��me�����E��}���ؠ��ܺ�����4w�n�j��Gv�=��_?U����\t���X��u/>ʴ��T��ڍr�!d�gm�q�S}�Wvr���Θ���(r��t{�í`J�P��Z�έ=�z�~�V�s����g�Esj�!�ױ+��㢵-��-v���fpkSN*]:Sfސ�v�#���~������/*���&�� ��Q��S�B|�Ouqk�*_l�}�s�������\,��M����o9�SL��WQZ��d�ْ]���8ߑq��r\�m6*����u���_����|����W�ܟ�-[D.��;~eeF���9�ۑ�z�if5��k�ݾx�{�o�t/>�o�'�����v���s�=03��m5Ξ��nL��5f;3;=�C����u~�ܶ�"�Vm'�����Ƿ�}0�y�W��Fr��J��T��-��'��8VFo�(�槱vNNU:��
I�/QԮe0���I'÷-Ŧ��r�`J�ж�M}Q'
�&.�z_��b��oOz���d���P���m:F��t��LY�J�]�t���Z�]�xr���{�E�>%����n��+[��G_��*�v%\���6�t��R�GHw#����n"l���	�B��5�?F%ֳ�ٯ�����dŲ�G%;��ۀ��b%��=�b�%��}2�����:�.�ܤm�w����v�&^z'C#�+���+
�{�}~��(Po��S��N�i���Pﯭ��m/�[�����ó��ni�Uԭ@��k�#�qu�������(xa����Vr�v��%�tpm����W2n�������Cy�6A�U�[�d}�MIW�Sκ���s�}M��g����ko4ga���Q)�����Q0��mc�����g-�\����R�H���Ѷ�H7����yNl��WYwH�*��T�D�)U��Z�lgZ��X� ��,����_)ʱ�*P�e�Ҽ���J=s�T8)���Dl����}��79����(��������e���k\q��'�pJ���2�[�:���3�fЈ��1N�g�ĸ���9�r�7j���+�ljiS0�O.U������;<��Sq�nnJHs���5�
/�HM�hf$A�넭2:U(Pɯ�^^�����մ�z��B��N�4�lI��َ�_�bǝ|��e՝�N���l��q��7�qjvE����씣�S��:PVr
�k*a�R[�lZ=B����d�bBN�ZU"H�n��b�=\k���ڟU�k�]�|�qK�7����OD�����eu�ݽ|��e���MV�|��*0�S��GٲN����х|Df;��Q������f`����37���̎Ix)�d����i[rq�W�k�-�NW��r����ȳ��yb�M�D�9}�ky2�R���2Z�����XC=
2�U�%N�݁&�
��DT�+�̳z>���nvg��_M�'��O*՝�K�n�����8ܒ1�ۧ%5�i�.�Nc���a�(�f@������p<:_��+O�pe۱u<ozPp�M
rr���/ �M�;��Q��p9/Rηj��[k~!�?�*.�=����lsMɦf�(�j�*��YY�ox���Zcm�5`�aĮ(A�;&ժU���&4��
�E@a#�^l�2�`2�WtW�\ҽx)�{p�X2�̙�wtp]5��~������;���lJ�����w�1_��]�sz��}AF�3��ʹ�������&L�N'n�<�M�X�Z�*|*+�)���GMD���D�)�I��HX�g:Ս�Xr�O�@��^�rH�ۛ�Y�!�kV��6(lٚ��
	o��֎T׭Awe&v�쑮���{	b/X�t&q���{h�}���b��\{�ղ��������w�ǌ��%�0Ȫ�P��o����V�����*��m]X���n5����Na�����(.���tGm̛��vww]cwUW�w.Gj��!쬼JP�Ӂ�Fr웝�, �|b�Ejڸ)8\��`�������M�j��6�w��"�
�=�A��{d�cs�)i��eط���L))8��`�Qm^�~)�Im4�6��oF	A5}��!Bi\/�����#YLi�����1]g�Lrq�x���v�����Յ=΀�:͓��!�VN��2����WO���F�1�Z�[�Mk�碋�,�p�n��[Qog1�"�R=��
s�Ћ���69T��� )h��F�a�duI4�IIE$H��C��)���h
����h&
�*�(
 ���������)�X�l4�MR�i��h"i�Z��JJ�M:)j����"�("f��$�ZbJi�(j��:I�:�QM,H�kTMAM)MRĔ햀* )�lSEPR�U��*��#IITQi�SElb"*�f�**���)ij�5UKm�j��(� �����%:s1%)AA V'Tb�$�Z��v1C��@lb�&���&��#e)���A�%F��)-�Q�T�*;`�K1�hM���i��hH��B�6���˭�_�}9 ����Z�R뱻{KBM�n-��in ��xusY��@m-�.N�6ȸ���.�h�kG��`?�}�}T*I:�c��V���,n\3����� �����V���:�O-�k��=,D���ΐ��k;_79-X��5�ۨ.;*
��;��ecF.�`�iw�ǯܱ']Lut�^���7ϛ������{Zl�ƽ�����{�ྺ�ί�uV8�Pu�V�T��ͮ���]Y�1C���3��h�겆8������_}s��=�Qʴ����+h��7����5���<�W�6t<��O!�T���?V�QgE���JC	T����Xf�(�ͼ�K��M��kU����1*��H��މ��fV���M�ؐG(a�q��JyoCݸM�)�St��L:�G�m�7!��j-�5��@T=�]7�>����J��H5��i�u��
�OV���=6X)>�1������\S���][�J}��c�\=4�ZZ�,�(��_�z;�*�c������r��K��D2���s��Bݪs��GQ��o��P� �~i�gR$1��}�,�j)���.T}�{������̬ɡ®�v_&�2SQr�E�O����F�+� �w��ﾈ��aN�nT��!ξ9ie>��.˸��4-�Z�f�.�쑹t��z�p�=�*a��Ʈ�fla��п�kˀ�2dk�;�K)�ΝZ��j�E�.�sv2)K1Q�H]�]��+�k���;Цt.�*sBp���ATkU5	�t��M:�bp#�^���^'�݈ͥ�=V�r�l�.⚍Y1!LgHu$��F��q1΁��U+];���r����eZ��Q3��ަTҽ��A��OHQɍC�r�Nڹۘ��$��/tn�����&v����ſ.�����v/Q��$^�NoRƃ���Go��o�αo���#eѾ�+�<��V�����m�^U"��U��P�ur�0�W�{6��;���T5�H\�!{WR��ӤVq{��� �c���SI����k���`굅+s�:�^L_>��#��M�n��3<$��<�7;�z]�[�k����L�\[���r��Y?�jʎDFV������f�^��u�4�������ت7��}�������yݠ��P�.��Ɉ��cWI�⍁NUE���3eA�vH�S�p�~������叅�װ��������i�Ȧ���[�'���vN����E����ν�\��^���#ݤt�|{X�#^s�*�z?�M��z���o @�ǻ�����bg�<�m�5�/�|��m}ڮ�IgѺ�n#��c7!h�藷m¡*��������W�D��)D�rjoMn*I�������F�X-���;�l7ެ�Z|��z9W���|0rۓry����q` ��^��y!=�����O�y���݉�r����`�6Jז�6�^@���������q�n�+iXV�\7��к|�i�j����|8�?�v�F�!W}/ݰ�y������K![�1+�},���3[����|����XSK���F���]�rp�ʜf���ѳź��9�Cӵ��˻�l����Q]�W�R�c)w���lx<|_�R��|K%)�Xw�m+�R��'ƛ��Y*��&OyX��7V��㕌Y�^u�f�n�v3T	�y$����^��9ڈ�G�kW=[�m�6�u	B�i��+J��ҦM�&��v��=9Lc�1�����;k�7����ܮ�K�l_Q���� N��yi���`W��q�������lc��R+�Eb�]��|���^��㪱`Ĳ2�wE���9�N�4�:5��[�ٮ�Aq�Pq]E�Uy9͸N	�'�iA]�2�*q�\�w;q�����2k�խ�y�զ�sS�7��t��S�����Z��+叧j���_=���s�����}zN�+;�����=��-�qʴ����_���y����0�������~�BI� ]%��e����֬rز����sw��ҫ��rot�z��q�/U��=����G�Υ�7�O���}��c�ہ�̪X۫Un;�v�oj�q�V,
Pj�7�J'd�fT��GeoD��<�j�,��=�5_�ZW�yP��Ӕ�S���r����ӓ0{�����y�s��}Wω�zdV�R���	c��(�Br�X����|<jsz�z��㘳mq�:�;˥�̋���{����AI7R�n���ű����P%�՞�<�T�b���X�?Z�Y�g�!��3��1<�������y��n\��9����,W&F�=�D����&wVp!&��7�:.�t�k�����G�٩��fb���\@}�a9��GW7�%�P�:��u���7V��J��'�=�8�CyQ:�̸��d*�a������yN���C6.f�����5Q�5�LE*�B�t�9�/�X��
�*��ʙ��$^��5���6��J�9vV��-WGی��._?����~��"e=)?t\Й�:u;��/����-�j��Ȇ�FEƿw�}x.S�L����l�]�kZ+�AgF��:B�Z��=z��ɩ���TX�*��fșX���n�^��S�n�'+�Z��Ңc�㋍LuC�ɨoUܵp�Q���ͮ �����啴:qv�M�]K�OԲ������z�TU�Z`���Ό螔j�K�V\ڞ�/����B�TB�����Wz�LO
�ꑧ���!*��+�n�c��k
V�0q��k��/�1�gi�`X�:�o`ۊ�-�C>ȑTt+�)���4C�~)W��7��9���)�u�D2���e^��żU��\�o+����p�#I��o )n%�;+��AiWg�e��'])5tℽi���e<͈��J��7]��
�6�_�#��xq�;�Gz�e{S/��=�p���]U�nj'zN"n+:��+:����oB��OO7j�Q�<���{���7���[p�t����Eb�Ur�ˮ��]SMnb���1Xڜ].�7�R��n1����iKce�A9�V8��mě�)�-o�v^���T&7U�ї�����HU���T������5mě��\.������T�[{���髢������4����E��j��-��b%k��,+e2�4h���Gb&2�ާ��Z٧7P�	�,�}�m�oo,�vN˥�Эݝ��:�*ȓ8�\�1ܩ_�8}pUï���j���}�Һ�9�hP���k��V�bF~ǎj#^Om�o�z��;�WƲ�������D�F��wS����yEv�\���U:�:B�Lf�8�m�LV^���ӫ�,:+6���h	�ܸ,%����U���]j�x;�ĵ�n��czKY�Uj�5t�m���Yy�5��S7��p��gݵ�;���O�_�� @�+��ӷq��8]s�'+����Fh�g�]Z]Ƃ���BrUgﾄU �n�fdO�z��+�x��r�=5��Ku�k��ʇ8]YP��beC��<�ٻ�-p��P3+�r9m�N)�b�Խ�O�\��ݭ��ؽ't��yG�=�3��5og�lײ��.qTY�Ð�v/w��ĉ4���Gh��N[��O���ks]�fwF`J�����,���Ap!~����\����-�e򿴭���F4�r��S}�	���
턎+��IZULk[�r�C��E�7�i��y��W=T���Or!r}��6�����<���f���W���&�u�*v��TY�mTi]ִ=�9�(���y�> E}���e2�D��դ�PJrjn1t�n)�4����\of�j&��H�,o�)T6�d@�R,rWls������fv�^�v�;D�}�S�}i�x�U[�
ћW��o֭�8m"��J:�Љ�go��ӎ���d,5�9�k�
FX��Uכ����q5�������q,,89�` �D���5�#A���Լ�9c5�mc���e���Q�dB�ȴ�Ϧuo}۬'�G�LW����#oujl��;�k�"%�33�v�5��دG�	�^s;m��ޝ��ve�K�^���୎��ÿ�]B,��:->���5�!��� =�5;�JX�:,�S�5j�s�-�p��U�Swb�v�Ffy�L-}[4c��ˈ�i�Ŏj5d�]\��p�y�q����j^�Q{�j��s�CҕV�@�C��E?l��Ϊ_���_yV���j����/Iܬw�7���@����
���BYg�{pg}�x�/'*1x����D�jqUgB[U��v�Sn60�L�VF��\vh\v����&����OUE�<)�=�{�h��1TF��������S�_súU�w����-c"�ۙ���<��n�v�Ž�/*�D�+{9	�����Wς:�a���P5�+c�U��㯭�-
�SycO�")�����&���ڎ�uU;/�wbl)�spk_�����4��Sޒͪ����Oev��HwI�Tƶ����&�81.,��Z���֯
�q�l���Χ�]檿�	Pܪ�*5VP+,�^�Y*�"�>���ܨI�ͅ^��e>VrY���fTn���jt�{��E�Ww�$�}X>�s���9(��g�c��P���ҳ�ꯀ���SO�{ŒS=7�v�k�t+םë��r��Ӎ�z��>T.n����vxd]��XW�|���.
�ˇ��[]6����hS��b����W�يct�z)�.��\�󥎾i�o�v�8���n�u�Q�(�\���I��Z���@�{�>�=Aw]�J�t��4�<Я�ĺF�ʗ�0��ó8J���-���%݀����I�ں]�Nc�UAZ݇z9��cx�����q�Ԥȇݦ&P��o�ene��!V}�9Iu��Uw}����&��Y�@U�Z[����*Y�!,���~F��lC>\���^;)?A+
��z���&ł�̸iC�*��Q�\�{�me�x��zDL1?&o��98�]�J�*�4ڭ��u�vƐ�}�g^a��(Ah�)Ӌ�UV�Z���}�k{A��pb6[��
���KV+#\['4]An�i{��Ƀ�ɕ�w��ٗ�ݨ�;��)Fۇ�#��$�ۥEᬮx/-.˝z$�X:�˾��!��S[�nC�gŕBtI7��%����]��WD�\��Io*/���+��p���ˆ�+��Ӛ��GG�����������i+�U�޼���OMj���9�yɾݡcw4*�ĵ�%*��ս/���A�v�)��v�R���,/�6q��^���_ [�\�N�uU���}5po+;��0u�����{��ixØ̚�r:�q)���F�a�Cqc{�������0%�vr�~�C_�H\�ɳƕ�z��+�MXjp�4u֔��m>�oz�d�����%W�_"f��<�����{����겹_Ѫ�iO.��&�ifr��j�]Z�!��N:�vWsq��A�͉��M�.��9n�����n�?�ԣ��^uVg,��:�u�{rnJQ4�����ˋƤ��z`��D��:�
�v)�ui��/��9"*�	���w����%>)���6�Ճ�QT�9��!1��݉�)J1\�U�9i�V���1�3vb@��.������Z�۔��w�ޝ�v�!%�Yc��ξ}��X�sB��
�zLO�9�h����u�q�2�c���u8J�웋�y�gw�,&��2�'`l�0��&&9��.�
�W�gѽ?j�%����x��;�A����/��v\��v�E�]Z�7��CP�Z<fY(R�X릣n��6_-�i�����5�V��@�YlN��@��Túz��^Q��Xۚ��K�ku:���Λ�Y��7���	.�HTN��sya:�EQW>�Ե���T������yAr C6�0�I�*��Tq����К{����,.���0���^���a�YC�1:������r{Ԧ�wЕ�]D�G �R�;�ɶQ�X���w<n��A|���Ɍ�]��]�2sC#��Q:��^��%=u��9+J���-ۧB��#���)ɂ�ոn������0wKn�%���/E���2�N�Gw�N�6:���r�`j�[��$�pn��������2�}��*�4OQ��}�����$�Y�7ٹ׏	P'��Ԗv�~�v�F��_X�h����a��0��9�Z���nl�v/�>*S+2�ӱ���*�� ��T�O���g��-���s.��)�7"�+�:��B5���heة��/T�+�R�7.e��C����s��gOJZ��k�0gP���k�������=��]��C�T�	Y�D]�
�44A���wQ����j�/������&ѝJ�k����3��}��>��s��%]��v������e"煾�a�\��#-Duv�s5���&sf�4��JmՆ�Sx�lǓKa����jHܺ���5�vC2�>�:f{���-��.	�ޞgd��Η�Ct�q��np��[�nD��DlW2U��I�)�<�>�)��cTznXK;1����ʳM�T!�?[M�h���o*ۣd����B+���K(5b8��yL��<6�v��Hjݤ��\�]�~"4�fJf�.�'cH]����z���7SqO�,�YD�DLț��9_g\�y�Xo�m+]��}�խoA!���y!t�jĮ���DB+hTj<n���&�ΚK�bwp�[��yy;��qv "=x"���7�\��d�T���Uw���C��y���<R=���m��*��%{P*	=S�r|MsN�	i�i��)��;��Y����7��
)���yU*R�B�=.
��gN��M�G�O�����U�՘&�QiNک�>�\E���<h�i��)Ұ ��#��;6�k3r�\VB��z�
g��#���WfXgE���7C@�ҞL�N`h�f�P�Y]�]}���5°��"��ulp�����R��h��#����-PPC%m�Z
���M��X��M���4��PQA44�S@D튣N���b+F��ĵF�P��ЅP)��J)6�m�4�:Ck6΂ ���(J
����R*b
*��'F�4.����ڒ���
�i����b�B��&�UQAMMCT1(ht�:4ց��16�i*�]&��ZѤ���������@������A�)i�B&������&�M,�E�P�}���K���#�b�*�j�����Zy.�)��"iJ�"։�����(ZZ]������۾�~������{���Ҵ'Y,
�y����gp��_o����b�9>\|ǳ�Ф^�j����$�U�po+_�.ґ�3������J��u�����*:��4��rZ�.�"�;�ά	l󼰟geRH����a_�ҿ�p�*��Q1S1�3�����_W/ݪe�Bc�|�굦c9�ד!LFt�_%��&�@N���^��im��Xy���l*2�W�x��V�1���T�3�(��C�vt�%�9ˋi���}Cc=[n�7������[K�ƾ�3ޯj�A�~[��^:7�uvn�4������Kjz���eŴo�����<��U�kO0�o��f�����a<j&+m�B]�i��õ���9�Ud\���@B�tsM�+��x�M������gw�*�O}���!�i�`�+��6��{oV9�|��rг~�-��%.3��<=�*�h�K"��7il��F���m�q7��U����Z����y��UB���Ǐe֬��	46���K��߷u�g�T\��6��K��i�LfE_@S���.ĕ7�Y��R�>x���=^�񼱟�UtG"�_g��<��1�OR\Ә��V若��Η[�jNW��eC*�d[˥�fp��JYm�ۤ&c��ʿ�}@�;�o��_�����B͈���M>U{j#U�Wt�o(ყ�uj�ޮ$����q��n�e+���|ʅ����)D�&��M���]�OtN���3���o�jQ�&�%���9mě�ϯ�!��u����X�O亳Cկ��69ؚ�<U�	c�N��T!���3Ooe_Y��5fC{��
�W[|�B��biK0&@����I<���¹��-���ܚ�Ov¹�e��u8l7p�_v+cqL�l���]�on���Q�[yaM<8��+�B��f�x��j��ޜĀyU1��N8Uʜ��4�n�̫[��8��N���N�[��<Q9�V����S���G�|��/���^���V!�,/b��_���J���̰�5:�:qE�g�왆�uF��\vT�G<���*�Y˕^�Hz��m���ɴ#;����j��}O�<�ٙ�㖲��<}G���8���4*�e�Pk��8(6��k��^v?���Ii���8��]%Y��t�r��K���b�w��ݗ��Ӻ��:{w�ƌ���f�Į��T�*�L�	�ݏ���X~�ʥ��Y�U=	�����b�]���1ң�ۅ��T7�5�f��MOp�1m��>��Y�^%��r�'�=ߗR�~*��ϫg<]�=�U�z����x�H福{p�H��J��&g/�^�>��&s5S�:}=�
�/sZ ٕ���P�mŹf��#�q�؊֪��zy�9�kq(��Y>�OwOo�.��xؾ��x]���k��.9�C���i۽��AO��n�r[��97��nn �Z�Q��I��Y��i�f��PIc�='a����F>�x�i\C�ݷ������_�M@b]U�����k�bB,�a�����j���?.�U��R���� �of�#�s����B�'�cj�+g�ᮣr�!k��!=��Ukwގ��ީ�͙f�B��K c��=v�1�>C=��ene�̅Y�{���;�B,�^빊�^RJ��nh����~
����_����>��t�)����1x$h��>���nu��ڵG6����u,K��G˵��N�}�#;w�J	�#�i8�ԫ)������$�ի;�'&~�y�p�l+y������.���Wa��c�uQM�J9�v-Tm��1��T)�q���k*���>��P&9��%�l����q���L̯"5�(����XQ����+�:C���m58����}���c�EY�>��a�ҽEs���.�;M�F��|���X,@s�������f���U聒2��uo]}y9Q��oϨTά���_z���ׇ�O���y��ϵ��O����uE�����q���M�����]�$�&�����{�����ͷ9���J��Xqv����r.X��+�q^��1����o���W�{^��j���y�ؕ��k_��P�q�3���N�˧y��)V����Mt�ބ����:�=i6:Ư0���{;��ex�Y�ݤt�Ƕ��#���o��қ�|l--��7r�ŧ��F�le��ni�X�C#����k�P��SV�Һ��Հ��f�֯W��<0p��>�0�h��[|a�P�[�ʼjF%�u� ��A���3�c��ծC������-k&ߖ��ټz���j�xO��{H*���!�F��H���wRn,��I�1�gL���>��Tf�Ь����Ov�!�͙���Um�ӑO�7�����ݮF����q�A�����I��)D���wV�)���ᑄf@���;]q"[�*�|2b�3M�*0%�-�6�Ȁ�.�?��]�['OV������k�*\��
�54��}ǌO�Yj�%�:Jט���}g�E�pd�O�}��w�ݥacf���TCx&)K1_t��e�۩�]9hѡ��6<�W���Ff���L��r�-p�|� �=�Ӱ`s����f�+��Gf�je6�1��ٯ�����4�"y�8�w��V�8Vr�b���H�>F�]�y�v�eM�j�j-*��ؐ[b/:�e������g.�W��~__f��T=Qh\O�:��j�1�F��M��;-fk�g!�m�7�����C�ɦ�es��NG`�Ys�Qnp�iG �S�y\�D��Hc~5���9<(f��z+�Aq���0��Ζ#��$�P�&�;`vʭǥ�*��v�ŧ|<�h�/z�E�NT���@�>�KS��"lus���W�nK��RwW��E�~�S�!$c�2���6^��b̝Q�r�,�����.�7��/��<�PEC�E�^�����`�Ǣ~�Z��|���m1�_S���ҟ���ܔy�q�9◫:$��N��k�S�ɷN��+�Di[_jo/��=��Wd��IA{��e��px�}�BUC�H�M��YyTY\�5Z�Ҟ\7="�=��K���7�\�W��>��q���1*��o�2�S�{j1�b1I��{Āh�D��ǳ����:R%���`��=�A���}����/^:���jd[��9���m'�s�dӤ��r	E�XE#8��j����t$��Z_>+�������r���O������O\���ӄU7r�s�H�Orˀ�2�'?ww;�+��c���V�Zd�۳j���]�<�����pՑ<�����ɬOv�+����i\��
N�ذ�IIz1M�ۼ�#��t��+���X���b*
�KB�m��^�����W���t���y0�C���v2x�L�|�W��K#7�6�yQ���kp����\�͸ O����}�X`i��m+��tŽ��נλ�$�i�zp�����>����WZ��PK����tR���J��u�m�f�\FXS��,sQ�':����ݛ0�yU䅱�+n�q�J�2�@WΜ��4�lͼʵV�F,�>�&bnh�{�S6��U�7i��aX��z˃�=�;켼|.W5(�yԽ9/��Wv��Kw��V�Η�mɘz&|�V��W-�A�k_��{Θ�^��U�O����c�Pc�D�<p���W�Y��3Lb��庳�C��x�[��=N.qս��Q��켸�Q1Jۛ�6��7���c��V��lvK��\��W�`y_�:��s�_R��8��rЯ"57�|%�"�nYdt{={5�[���2����^v��6�կݴD���O�|n�
gl��ݛ����}�����Ss
l�\���ᰎ�[����V.��]l?S��B���GoS�Or�V����������Af�-
��Bڍ�2�+e:��z�
(W��L��s�TlT�kv���\�cK�p4�X7����܌���e�ܾ:G�d�����q��$�՜n�:��)w���ˮJ��/I�s�R!V��u��5�q�3l���ߒ�]���2�~�F�hS<d�#@u���ː�f�*�NϙG�&��'g�Ucj{�]?S�_4�Mڡ�k-��u�M=R�*j�ա�����1�DM������.�ԋ�I�x�h�)��Ħ����e��k����ƭ�'��.�؀�n����X�U��i��Ն��3{N94.��n�F8�ֈO*'A����ޅx�̇��>�"��'�pp�i�8ٿ��sw���f�oM#~͈m�`��,�J�f!g���`�q.^��@��Uà�'��=!����K5z������sc;%�3���zzB���8_58�Tf�sИ&�*��oMiF3�~�2uMNc2�\e㨼{�A،Q����
�7*u:�wW�U��iW���mBu=B��uGe|q�}�U��F'���#�Gs�,L.S�t�p��Ef��kW,;��^Q�u9��mE��0�F��fFJ�Dev�Se՘�6���'�c7U��L3V!÷�HZh�h��{5��&GZ��(*��J��ئkϑy(�ݻ����y�e�WYZ0@���r��m5�y}��SO���,���.�A���B��5�Nua��7��N�`�'og ��%p�""��3�������R{I13mGh��nQ1K�<��kt���aI��7Gki,}W;i�ZgS�uىd�t�����WR���w��-�|�b܇���1�UG4Fi�w��]c��u�f���Y\�7��O-���֩����t����\�jX�����:P��sp~������]4�G.�Z9GlgU1�x1��&��&����u+K�P���J.��x�k4.��>�ݔbz��Sc]�S�*}j:�9����jQq�.9ie>�����L��x�0-þ�:���:�n5[�I�w�WO��g`�@8O7�7͔��o\�c72�s��ߵkf��§�ĩb����<LB��ޅ}>�m`��d�;%����=�U�!w9Z��Uà�;~1��"t�}���1纯D\��
d���rL�Ƥ��6��%��勴��oSʱ�/�p�����AK1�<'��
Q���V��Ϸ�m
�s�1��|�B�: �x���:�5u�X��B�kE3��>߈zXX��eZ�#�o��'����@n�ZNͦ��˨�7�y8+|����x��;��ͼ���V��,sZ�~Π�M�ԜO�wԌ~P���߳�;5��˜רM���Ux��5h3��U<��e��Nzt*�B̭{��s�±U�X�B��ˊ.�Y�j�-�c]�j.��(Kj����:��ת�>ݛ�`���<�.$(���c�y��Y�O.��8����[ѓ��<���%����y��6}�T���|���V�|y��-��<��q�c�u^^�ݾR�rިk���=��65��WZow)�;��U/I슨���WL\dγy3��}�!��~�i�9�w��F�B�o�FX.���s�m�cY�F���/�W���WIՀ����ɖ�G���qu�*�I�Q�n�ͻ~�ݙ9ﯝ���u[zK=o}r-d`=�E7p*.|���d."=$?B�{g2��7)#7��U��O�q��G��~VT���Cf�=.�}�Sh[���3�B���,Im?~Ya�sJŊ�����E-|�����V�
���p�,vZ���/��EK�n��(�J/9��Ǣ��/L��"����"�͖X�,c�MV5����+���n�&.bv�M�B��,��]�4�L=�2�)hc[������<�.�Η�ٍ�N���,#�]\�F�p�a��|��/��:����
��R;1�h��:�%��\�J��%�۶�މe;����
�C-̭}{Lak�	m��`yٴ��Rv�#��E=͘�o;����9h�'''Γ�:����U��on�
 +���bs�]l��R��f^�m��t·+#3�Ǔ��/�E��m�������>�2�.N���;�r��׼���Qs!ݽˎ��xփZ@��DXJ�gv�Y@�t��M����MK�"]c8��&p��7��4�>�ّn��������{*Ӗ�%�J�������=к�n��ٸ
���XUŒYX"�"�s3o����^Z��v�|vT��A�&�j�\����[�!��Yj e�c���uie���ؠ��
[Y)L��|�/����u���{�@Zq&�$���H����氭��,k���>�'gF�8�Mr��Q�6µ���9�,/����}���S�(ܳV�e;i靯�݇�Mt�`���\u:�kY4ěϳ���MN#nl� ey���D)�h�9mXÝ���Σ�W�(q�����W! ��dZ�Ko �3e��E�T���l4J%����V�O�X����X�G��J�&��m����G���u��z�:�޼����`�o�ᤑ9r�PN�1	HQ��l�pf���f�x��R[>�پ�#�}�Q1.m�|
]6�͈�5��ƅ������!\+V���g��44��r5�[F2��y�&���,9c~g(�R�9���R��*�R}��YV$Y��^��Ó+����M�n�+����@GRH�o�r�u�	���=ب��[u�i�V�e����.���I%���]��#��tk�:�(]
��{vZg���xt9����ve�f�	�\���>�1;�O�,�aS�o�m'�Gk='�u�׏�E���fm��vz_!�l�pA[Oɢ$�#> �.� ��*��za6��Z�?/Oik`ӋϤ���9����]�a8� 6����&.�V+�Vu��ڝj��c�oA���jI�#����x�x��w�H��ӕ�/%�GL�WF��&�5oѝW�ԢE��uΕ�j�ϋ[X�)�Y��Wܪ=p+-�0��h��YJ�}x�5nV��2�ה�H����9Gj�6���օr�':M�p��Py�Fn`bɏ)��x1���
�d��*�\�-Ko�bO{�v�ܧ�-����w	=�S�c˟vr$�)&��bt�:≛���97,��Aҽ�dٝn���[Ky�jNV%�����~㢟�����-�����i����)�d)�b�j��*J
6�D�G$�%%m���)j�ZJ��N������֨�"�
JbJ`���J�d��$�b��h�B�Xh�˄STEQ- A%QG'�ږ�R��M8�B���"
��Z�ht����
*�F�)�R��JJA��"hֹ&b�B!��Z)��唨�������Eڪ(�4TQW-<�M��.5�����RQ��R ���ۖ�d�DE4�T�%�V�M)�1EuQU[��l�jت�))�����(���(��(P>��a��+�ȝ����^���o������r �
:�޸��}�z��;XC}\ݞx�|p���d�JÚ���������/��J�{!��1q���r7�4������Q`@l��^�[��}w���������L�Ç����௧��U�(c�R.s} s��fA%�B.;}��4���͹��t��<'�ݑU���.��	h���=_.�<��"��K�z�x�C���=I��Φ��@��ʪ|� =eD.�v�Ɨ�����>�U�]I@U+��<���v�:�π�6 �D7�������ٴ[��/�G���X^�Q���34ML�ǡ�/2/�d�vz'�}}sf�~�Xd����}@/T����w���տ���ߍ,�~��5��VaŌ�܀���$��8�����]3.c�����ު���<�f��?He�?��S]��G~����������y{�G��Ei��`�mx�Txj�w\����s�~��1���f���75q�5.���W����_�^���l֛�} o����i�2����������A����ʇU��n.�=i�\UX�wi�q��:����{���q�@�q�#�n3��V�g�W��T=j���P�׶�TBQ�kG4�cm;]�Eڞ]�V,���
Q��Vl� ��A�1)�U��[����L�_{��b�<b��魴b{����*��������)ݷh)��R�t@���|/����4�O˳ıH�B%�nr��txq�jf�h���hꨧ#���茹j�s��?/1���գJ������L��&WL����ʹ�EU5�,���n�'>�]S��� ����(��DS���``���b��	Nb��#%�߈w�m�/���ޱ����/�q���:�q��5e���%��j�}�U`~��H�v�bJ����#��B�2e����pv_�z��K�r�G��,��
v]̋���mZ�=�ҏW�߀��Q3�@��)�Y�¨�V�?:a�	H�o�i�z�q�;�]{�:3k��ܻ2�,̝�B���鸃��{�H��+԰���l�J7/��oґ�/�|�Rc���\�s��T�u�+s�X�[XfaŒ�����Q���z��KGw��uC���|��+�y��D�<����W�X j3�dSʧDZ�,����E3�s~�ђ�[3^���=|[��N�|��C�5w&�^>�q�^�"=���������/�g۔G�a�T�q�| �˹�V�+�L�Gd�=�Q
�G��zna�H�J�s�=p��^���Mϑ��X���땗���\)t�;���2��Y�JB���-c��/T�4V*ºuh,'\�:2��9q�����4iv1�_r�{%�nz卸���搳��CU0���)���f�
#�TK��@�(��s�GB��q���OS+=s�3�m1�4K��{#!?P=,}��n �lg�5��ۏVy�>�%t�w�OT-����ͯq�{i�&:�^���.W���މ�+}�%�>�5^�tq`�~�<r��Go�ڇ�=�FmV���zzXU: ���/�W��7g�!Ц���Bx�#��@��O���3�4��;,e�V�+��+����Nn��T��j�.o#|��`?j�&�՞>��z㑸�<W~���=��#յ�������kK�d��|s�3w�ξ�
���=�G���M��iח��w�;���Ǒ�}|�}�IlۧZ
�F��.��ë;wx�f�-�=9�F��L�_\k�8=�>�"�^F�b����ό/H�$��g�dnen8�և�}�<\��=�_�3d����
9S�p���~�����g��̾�(�S~����=Q��s윂Pn&��M7@Z+�ҍ�h�_���N�9�sq�&r�|T�̕KЏC���~��@h�����b���Ϡl����,t�Q��-�
�MO�#j;��[��y:\���m'���o.m�����S��wT٬��aA�R�]�B}��T��]�Gjj-��m�cʋ�d^���'�-��UkP�*w�eG��?X��f4���Ӳۥ���m����GXOF+����@��6�a����5��	��w���q�T��w�tU��ȿ��Iy��!�4��L���]yxV9��BV�Њ��$8]�"����k��9������(�#���Y�\�7��>f�ىA��^p�C�>��d�;g��E��:0�zw���W[��s���>�8~ی��5� 3�T1]�=�}��½+.f�IV��|7xKP��K���7�~�8*�piNo:����s;ܧ Eߠ��5�%)͚���7�Dg����^�WO�T%�S'�rƺ����fj�1�MW��O��
d[>�+(
^�R�\D��d�ҩ����{���f�����R��b*���wlz���p�/UJ"�6|5�����g*l���o�'��t�{�������K�_;�MW�1w;��|�>�q���תQ��۷q�m�6���7��Jq;Le1��)���҄�ܛʹ�y���tV��#T�q`j�p7����`bu�9��{������;~���1���O3B�����A�۲֬�:�,���X��R=��lV��#[�q�e���5Cڭ~�x|Y8wB���tuF�
�L�Z z5�v��kh�F���յ�n�}2$A�*.�I̻OC��-f�ٵx�'�S��:�I�3��j;�xf����t�^�O��}�;}G?�1؛`fJ\;�tsfI6ڴ�h�b�M��h��BN{�{�99tzm��gLz�^g=S�JȪ�i�R��γy3��GT�:�����μ�/T_v\)�b�
n��t���ք�*��DMF1]�q�S7�L��r#�T7��^�}��]��d��9��>�)�)W�Â�X������~�%���r"��4�����s�v�]�^�SBA���ܻ�%>BuO�ym���H�G�ӏ��*=W�W
��p L�zU �UH͊�J���}|�k�w����ע6|��}�~��dyI���5~�p��+�Xâ[6t{��Y�2k��'p�r�;U���U#*"gx�!��k�}<s�^,lm"��x��ˉ&�k%xy���ܝ.�q��<w�\LO����	h��	cԧ���L�y^(����Z�Ƶ�Wd^�z�~�fAn���M�B���1�O�h�i~=�a���>�ۮs��cѢ2(��7&5:Y��⚰<�=5�yPO�.@�����5V�ܢE��Miz}E/r���.�;�W����S���P�oΦ����亭��+��.��x.&n|3cr�6��/j}0-U��K��3n7�m_����Y]�<�`u��W'8#A1=�xzK����e�*a�MeC��G��*(�4&�3<���)�<�L�<�;d4!Uwl�U|jD�ս��_�nV�HI�L��ɨ�[�	dO�����ム뷡�7OA��"�ypғ��>�W�R_�o��x�ʫG��9e���/NO�Q���t�_k�?�+�O�+�����;�u���z�q�q��u���Zj��+4�Y�#��1������k݀���x�م{�W��f�ú���Sb5U��π{>Үk�CFϢ+cG�J����3u�(z;�+E�{��;��ë>��xk+j�z�β=�<1g;aO�D�c��׈y	��v�ס��<���yh�/Գ��T�6�]ø���M����<n�]���l֏o^�-�J֜��>+�=Q�k���w��\�-9��U`޸y~�NՃ�;���vA�}8���z6e�����]zϾ�ޗ��ؿO��u��rۖVF���n%��RɎ>�oS�+�**��[\������E��X�ɖϳ�`v:Z:1��.9��<o�~��%�՞H{
��3��$�����a��z�]�UH��L�QjW����E﯇�����{#}@nC̀\�7q��s}^��Bb�}GҸ�z4���@}2E�*�����f��,��'�6 ��#o��x��/�VP��=��u�t���s,k�{���tL�~�]�<�3���2`�η�Ϻޜ6��3.��h���Mǲ�2��^\ƊCȓ)�;��!�����V纵�$��T����}�E�}Ǌ�$�����S�>�J�wv�#s���~�r-��7�󑤄�z�������Ɨ��E9Hx����o��#:�ާj���<
�z� �3�dT<�tE�/Q�`h+�{謢)�Ӈ��q�KRgN�Y�y��Kj���2�}'!��
����-�zH�UD4{>�e�wC:��s�����Y�.���l�25�g`1j1X�w���1�����C,z�����Qtq��|=���ks�^?���P��_��8����t�cڦ�b��T=qB~�zo�9��Y�Z8�y�B4:n�yC����;�O���R<g�=�7�ͯq���3[L5���'۽!���W��N�e5����M��,߷͍fia}�H�t|�6���}P�6�M�ck� ��o�������MC���=�[�w�����U���uߞ�W��i�X�֍-f����rٿS���^�4��z;|@{>G�׹X��W��<�uj�s�>�G!��o�tuLc����	�&v������}������>���m��@�>~����;���w�w��g$�nE�i\dI;��^C�evp���9��^�!(wZ�&����3h���ۆ`j_�dI%|����oa�v���-[��ae.�"��8�N����x�ˢ�]:���v�e1��?�V��/�5�9+���4�;��d˩r$-G�fřH��>��^~�g��r�b�&u�ɟ"�:d7q���{μ�mϼ\��ǸIh1;�WR�ye��Z�>2a���n��6˛��&*y*/ҙ�X^�vPҽX���>�R���s9���Y.]{�z%e���ToC�Y�2�}�Q�&��+�R�]l�EE�jG_�����ܮ�u9�n-�LM���C��0���C�ǫ��jk.Ypr��L�=��22�%��Qr��T����,ܳۥՋ�ԟF#�\����G!�J<���[��ޯ�I�:'�숩��yC&y�y�X�v�=���4�U�T;�]~��L��G��(�>�u��˒|�Ƽ�L8-\mzruX�:f�����U��)�\�;������U��0��zg'Ӑ��p}ע(ɔ�}���2�2M�u�{$��T'|{'�q����bi��7�û����,Z��7���:ؽ�w�*�ƾ��d&�������
M`��j'���]�����WI�����|0l*(?r���#ל��Ά��g�BJ�hzd_�Ay@W��*Q���[��ӛ�P�����PN�B`��]*Є�q�\1v����1���1�*��m�U���2ъkx<���F�ӸN��e�I흮n���]�i�����/���:u.j�ѧ���8��2~b�
j���ɸǚ$l��OA���2,ZJ����^���3�s�h�e8�>�Wu������|�z��d3��\Gz$���ó��\g�C}b�.��.�_�g	4ې��\��L�q@J�\zṭ�>k�(���ۊ�{l�CǧO�P�X�]Щ��.�g=�ݪgg���e�FJ����M�`mBwiW����)u����_��(�؄�%t=�К�/�N�Gه��9���C+����k�5�T�nu0Zn��l{+GE8�x�ճw���s�
v*P����Ol���M��N�*f=�~�t��L�7�L�'�R������?-���H���~3}�/Ƿ�\y��6=�H,�ti���p795�z��)��&X^;�Y�wwwF)Nz$�/D�+�9�����ʱ_�W2��?Q���Ϩ��7p2��V;Ρ��ÁY~E���q���>���H��>=�7��ߪ�~VT��I� -�SյV{<�zU�ʵYU����*.w�f���Wש�okx���b�n�g����{�GO�{�O�W��Yn�z���L�y/�a�.W�fς����Wx���ԋ��} s���G�{�dx�M.b�V������;M����)@pI� >�6������C2ȓJP9�X�:놥�SQKgRy��n�{t����~{S����Ԡ}��W=���X�� ��-��]�=T��[�=3mY8�����ƴ�ڷ�����(�3w�0<�MG�xO��:'�슬&)����wr��{��Jj򏪨�Xg��=������9���
��j������yC�ߵ];
�����a~=�aٺ�>n|W�(��/���7�~8��� ������^�B�>+�pxe�e�<�����y��X��k7H�+s�&���;���*�G:�7����s檸{���}>���7^	�����%�⯽�2��/!�[LM}�ƙ��ǩ]�5�3����ޙ��򍛏��^����g�)�����s^�;���nDl�y:+M�5����\xo*א3�����Uc��bS��Ϝ��Ȯΐ�d�яsPk�s�8��N�{2}Ņ�Zn5���`J�d
K�~0y�g���̭���?C��Շ5e`��=�+E����9>��V}UFV�;��u��5��H��POzc|�F�Fﺑ��[#��rF�|��8�z=����8_��7	g;�HiS!��Wp��ɝ���k@�w3�>9�u&����|t���~ӑ���}��z�h���<��DSfl WEV ���M�L����4�_�	�Gq=D�J̑=�D�U�*n��[}���2������MǴ�g]�],Jv�>�]���r=hĎ!��Q���rD���y匭'Ҵ΍{�4�f��e�2Ӌ9&���E�u�c";�b���V��(�F��m#��F�.��F�X��^SJ+�4�w����M�AC
_V�zh�I|��;Kf���Y��v�}o�}��if��랪�0:�,V7��ՁT,�����c���ogm=��}e#�Ǻ��݉z�hOV1*�4����)��ԥU�*�@�-=��r}���8���N�UI���e�z���S��
7����jW��[���MU�Д�o
�^��,�S���{��`9�ck�� �ܥ&uj�C�$pp��U�[W�=��ԛaWk5�`��	�=��'Zr���e��8���D�WZ
�F>��P�e�T�Ƌ��pޔ 뛞������:��o3nl8b��Q���aV�v�s�n�!u���ڽ�Yɷ�ﱦl�=�]����8���i���3֛F���bҶa��$7�WÁ;J�r��z�a�yLԌ]tY�+G �I�>w6�[0��|�� 'YN�ϖ�Hc.������ظ�%�h�D�� /k��[�|{;2������ЦG�-���Ϩ���`��
��S�4==��ݗNN�E��rv�${h���pU�ˤ���b=u��9g����f�Q`M7t�БM����j5V[���W|H�C���Xk�Kç�i�T-x�B�s=�,c��[@K�fi8�
�C���a�2ћ�iN��b�Qd�8�Vy8��"����i�r�AW0�6c��q�=�C�p��^κ�E�׸AҰۭJ�Wr��E�/S7���]���)Iy�d=q��w�R��Y�]�i1��̼�#��&���1��+E>��E����vN�\.�v������l��� ���u�_h����#�d=fc�WG���X���V��rK�����I�g-lR����;l��ɉ�(��ř"�sݵiέV�i�9�ٖJ:�0��,r&'���WpVM�I�l��wse=�n�<�Մ���R���ǎ[�o)	����+����\y|�b�R��(Sэ�����x�x��9�±Pg�irrE�lNmPjƚ��DE�S)�͓ 
<�Py�b���a��uоt�E�لVkR,$�6�<YO���W�w6^a���೩L��;~Dy�o�e�:f�S����
{����xt.;�'�&��*�ᮡN�']H�Dĝ!U�}���+t��[IK R�V�\�(^�!N���:h���D�-����Ų*ޫ˔65Z��X���5sj#�����܄姆����B�gNZ���E�5�]Ǳ�Mu�#��GX�F�{k1�U��W�nfZ#�T��!j�K���%�
�(5@�@P�'G-4�[j!h�4�A�� ���ti-�M0E:JJ4�HSMP\�bh*��iLZ���#@m���k`�ӪtQ��kK��nP8�T���h*"��gs���J����mE1P��SHr144D�혇F$���ILܩ�E��!O64:�TT�b"i9r��-1�܎G*"lsjG�:h�KG%�1���&�-X�Q�Z���Ѡ�.ml�l`�-i��bj�l�1�h�j�u�ZհSF��,�٪Z�Ԝ��69�Ψ�F�&����:3��P[4�Q@C�( OĒ(�*����ɂ�m���X1��$b���%���r+��|r�-X{9ΰ&�g֡U&���չ����8vZ�&�6�mnz_Y7�E�{�?FL�����sޗ�ѯzG�U�5%���H�7"���'��v՟�������~�@MO�>G��e���X��h��|=K�{��7����/t��^j'�Tv%Z�>4a��N���dUH��e�Z���6�T�����1q�=�Ƈ 莿*^�.�ex�F��G�A�g�!�"�@i�H�R�KA-fF�5Qu�X4����a�^��p�Uk�}{H���8T_�܇���46O����E�K������W����^�S��Ù���<}]B��x�7<
�z� w�� S�rEB�\���x��Q8fP��	��w}���H��*=4���11����s;��8�h�e��$Z�!��'۩�ohE��}["|�o�?DnQ��#b5�xv@,e*��^���O�c�v$�T��=${A2߽�j�G(�&�{"k.���w>&�\�3_m1�SD�Z�z��O�L�t����;�ͳ����B��ˀ�TK>�&��ۛY��׸����ge�3_��-�%����*���$���|�Iݮ�e]�FR��o��� �`g��1L�X��$�eM�L6D�?ǘ��+��<�i�>�nk�۱\�ޜ�:��2��&;J�R�k�%�u���^�#Ƹ}om��X�MX��uq����(u�9,�j�F��s�S�]������qމ<r��PGnv���t�_f�i��vU�=�����;#=6���,�@�V���N���^���n��	��w�kN�H�g>����[�\���Ҹ|����߲��8�Sq�k�@Oԝg��}�F���qW���ڞ<3յ���󧆽^��&{��۬qz��Az6k�o��L\o�/M��G��?d�u���;g��T>��m�;�v|#�{�M{����ܧ���JENN�6���/��o&|�Ȏ��x���u�{~�W��h�j�6�������i\�O�kܬx��	�z\�.fh	<��̼�a{":�.:i�4��͠%Fd�M�uʏV��Y�w�î%RYX]�ϟ����̰���M��x�ͨh���Ƿ}.���O0������G�O���X+�����r�/ l���2��NE_Kw �|}Y{7y�gu�-������xTy�R+�>������W����s.O�	�:%��v�0�cof�Nm���D�����OV�������g�5}���_�r=3�J9�H��3�dW���5��2�����Q�rsʕOi���l]�h!�KQl9�{�ZFڽ�7R�R�x�3�Z��O���Sٍ��iv�'pc��~u��zy��M�_U��Y�K=��E�m&"�b��n����|9Ya�b�ݍqµ��I�˄�k��q�s�O���'�ݑU��R�gF|}+N�/wz��:�u1o�ޙ�^��#�ݴ�
��T�M�p��qV_�Ǳz� Tz�v��ǖF����>�X�d�^�d�����C�]�����r}*pC��/����	\���n�9+�c�5���z����>���o�;�G�7���Q�ݣ�бD���}��g�/z��n�?�����h�Qz����7j�m{��^� �=�g�R\FG7�g�>���.�XȍUE�z����b�h��蒎\O���b���xl�51t_	y���7[�ZoO�<<����nk|@������ۉ�*8i?P��G�����{���}�O��\d֕d�Zo}#}7X�@�U����n��s�v�<��r�hM_{OS��:d5f��̯N��/O�Rp�ʦ2�&��q�;�z�vz�{s��'�M_�j�w���]�W������%y�v����n�l�K�WET{MF+�.2gY���O:�1�S9\KS��1j5��s��}~�n��ѐ���Z�˔�p79Q�LWzW�Y]��g����N��_kL;5�=R��`�, ��Οn�AԗR'���dv�=w�+J�F��R�	�%�qwwo�=P����׳���a���2)2��/��Z���4��dH�Q4�`�ĪPw�>��%H����7�d76o>�]�7S��`�Ac�,�X��Gϲ���߸��W�v{/���Z�(�,�|��E�Pg��W���Eݍ3����=��s�=�K���{�0�I�����_�_��+�e��������i�'��Z�YGaB����R2�v�
����k6XU}Z��lǼ˥��=��N��H6ǽ�^�W˼�g�%%������FW�+�a��x�Fς����w��H�3�m���g^E,�����UC7�-{�d^���,�t�A�Ua1O��v	kgrcԧ��
��6��{B��)dׯ����d{��ٹq��׍��UE��>��r�LS��;���y\Ǻ2�`-C&dQ��)�֖�#�(��S�mϨvZ O�@����Q�[����$6�r�=6z�}��t��Q�qziP��|��6m?PD���r��S�5>N-]�mT`�*{��}I]w�?F�hW���}��&Mic��2BUS��gޙ���lޤ���+QBg/a]�.���+	��w��[�8?vN��q��3_m0'�\x\j�y������f�fmdZ���ݎc�7T�`�V��k~��z,T2�-��T8�T\���>����Ꝋ�÷��� ����~��f8R��Kru�:ݢtS���\��T;�6-7��Wf���������Ƽ�}��Z,x�H������y�oRWFt�U�^�{�\C�	�7.B;s�.2�Ō�8v5�뎦��d��r/���>�s�YA��)�����S�y�.Y��޻5ߘ��������y��k�z����@��z|��o���[�Cg�h^��X���x�k��Wyhp�-�<�g{�Z4�Ȣ��+�r�r��,]4{�5��}j�eO�K��x�3���}ާ��z�4�~�~�J*�J�M``�s�=p�_�R���1u_��ݸۈɟzc���n�;�����w����X�7"ۖU-�=����Ud���Ū��j>�W��U`MOx���ȱd�g�:�K�h�����=��2�`��Q���oP4ﳜMz���Ͻ���Ϣ�E�L�@�R�]dF�
��Z</��ؾ��{鞫�uRo:���VoѮ���dxaY�y���A�PdET��K��f�5]�tjӓ漖8��9�>�<=
��Οe ^}��b���P�,�z�eO��A 7�Q�����a�=�LN�������rSl������{^��ޜ�g�| y�5�S�/��>,\A�+ǌo�a�~���v�:W��ԧ8w���l��f�;]��!����%εe3h0�R�͑f�[X�,[���^��oT��YA9�ݱ$\﷓�|�ؒ�Ny�WL�֝a]�w�%T-+%{��7X�{���Ŋ8N�T֫:J���u��s3%,]�M�G�Y����O��xLy��e����O�]@;�:~��$d���q�l���
|�~���7(�ei��9��^T&)��Ƨ�S�.v��	���W�ʹ"��������? �Ý�*�F��mf�y>&�\�3�ǵM�F����p5K�3�mz*�s�\��=���
�u�TK��w�z�ۓ�a�O����3_m0��A��E?1��{��Q�.7��{ޙGa{M`��D�8}!�ڇ���P�6�Mc�R+��2n�K�8��Is�u�	�u��zw�^��,���ۡq���p����:3M�챗�=��q���c6�L�S�+{�ў{^�i`k��8��:����t?\r7��>�m�6�Ԏ�S��u�UD�y��ɹB������MiW3�b��HNx���Q��^���;��n�f@��k��y'S>�>jvO�Ͻ[Z
Ȋ�b�X�u��ɟ"�Cwk�82#�u�z� ��A��K���l�	,�{0����{�g�Do�S7.q�9U`MO"��l�;ϩ�c*�y����I�\jM��X�H�QU��j[R�;74��撤9�PsON{y|��M�t*w�o��=W�-֊��Sۋ	��5��Y���Y�U=��:+6��b���RȾJ�N�p2��z��s^��B��.�d`���r�pq�)��esD�9���p$ː伇zտ�?w����S�A������>�d��MF@���
�+��{�Mx�ߦ+t���>d�ǡ2������#oD�wf�EC���+Pe��-�ǦP�ȣ#;lD�:���N���Y��I�YQ�j"��ĿZE��u���'EE��ȿz��^|6Hl��IM0����2�L�f�deO�3� �-9�/ƾX���j�&�_�ǽ#K��Y�_���kuϚuw���yIp:ϣf%�YdM9�Ҵ��TGz�z�u]n`<�zgels�ҧ|���W���fA��sJH
��x��=�����5[F�\��`,b٩,o1�����{�R���g||���@:��z�5]Q�Ϧ���F�i�q������-����>�Ҥ�F}͖T��Dz���>7����.�g�w ^�(�ϫ�vA���9��ܳ�ɪ�J�;��#�=�g̴L��y�Wu�UK!G*��_�tWCTl�z$���i��
2T��e�<�^��zC��hw������{�Uz��75� dw����*+}�}4*}��/Ա=[XT��Ƙ��P�-�u��gC߅e�wSaP��S����sԻ�pHN����f���/ƻ����XS?J�zQ+�ۖ��n���77)�J�;F%:��x���C��=���o	�C���r�i�u�|̛x3{Wq<U���r	��J�)^imَĦ:f�	f�dQ�_��앟��N��t��|+Mƹ������o�>�L�n��>�}�!���g���nL�#;]��B}|�d{D����'
YLed֖.2g|o\����f����7�����i:��ՙ��^��Z:߲��,��/���G�t�ñ����gY�ɟ�-F�Y���l ]�мq�HC�����3�>��{1��A^k��$Pnzj8	��\3+�ɷ��d�k�	g���V}2Ǽs�T;���s�+�-��~\:�laYR�?I�����k������;��ıMm_���{�����-��5Β7�j��G{��7/��qV]2�w��	2�wjr2����g�>�9dUHʕ^�S>f�6XWӡ�~��y<�x��D�1 ����ͨH�̖��c�����}F���m�o��T�7����
�V��{��E���5�VT�ʗ�{��}��0[�j�+�3�fx��}^ӐKGw��f�}<I�{�{NAj�J@�#C�/��p���=��� ��^7��U��>��r�LL?k�,�We3�~�n*sm�=�.y��M�4l��kp�{�r�ѥ9��]�a=�7&k�0b��^�Rg[���rN`\v}������"�`L���u���A�^b������-�&�aչ���Ɋ���x�oo7׮v�(�	����[�4�&�܍1o���>�=�.� ����{��x��5V�)���.��cL�}��Е��r��4�.����	�K�sf���r]V�`y@T/]z��\����كߍ��K�Ǽ��?Vj޶���~4��Ζ4���P������?D�5�S��}S`Nc�qWcN�}424���>=�OW��N���N��z��3[L	���ǅ�y��;�D���V�eQ��bC���Y��G9��y�1��=�O�#�;P��+�X�͚�q�@�\u07�,�?{c$���;��a�h������H�o
н�{OO�aՑUFV�;�WY�1>�N�zk�5�U�q�<�*��o��*׫<z�=�����Z)ǵ,�z�F�9E�Yi�3��E�W��;��w���@L��e��~�i�������z���΢�]O�����'ѓ��s/�ƚ�"� �j���2����Q	M3W���<_��^>�Ы��J'������3;��gݨ�������*���*�ȱq2��s��t�tdF��.:dܷ%cb�j��']txd���u�ZI��Yn�(��P�ʕ���6�Q����(���O�� ^1�^�y;���_S��o=BV0N���N-ُ��Q��nR��a�D�i��S��F��s��l�u�I��:<�K\��]�������^���,�d>���eT����jW��F�
�����8m�Si"Nd�{ay��C+��z
��=��&��d�7�%��;*���E��%z�%����>�����j��Y�ړ���]l1q>t�~�@����~�r��CCd���G=�����Ǽ��#�y֮���W������PԵ~���i�z� �ʈ���S�/�G�ú2ͷ��NUWo`�]����#�NV��3�@vw�&=_7�l��g|}'!��
��� ���7g�ٸ���g�$z:������ܢ=W+L�g|v���j}�1|��R�����e��ӳ�7��N�o�z�
����F���"�"k.��ix|:OF��f�i�W�h�Tz^�F�u�<�А����%@���wP��`ңs��=�]q�ͬ��=���%�����C�5�x�k^�ݓ}�yھꏈ����y��u���lW?EOɜgn'j�uC��Ɔ8�V5�kB��e�g�Ԁ��|��|F}μ
7�ݺ���p��<{=TFi��?	��'��ԭ�������
�R�]��^��W%�@l3:�h��T�-L�<�YևN���Ȳ���w���).؋ܦc�;�u�4J3qg5�ݱ�vyE�i�/O3�h�#G<;�`��̬�kf�k���EmP�jEy�V��o�eZ���n�������r4�Us�o����-��Q��%�]/�_R9N�pnX�,�.iQu�õ�22��y2��������!�H��<�Ut�^����2����ã��}�t4Xj��ti��ؽ�N^�8�{3,�ڏB�1���GP��Ŋ���W{�G�� .��d�f�k��'�XƷ0�N��󱅘U��v�7k:w`�R�D5�rlʘ����b3�u��k,ѩ�AAd۽4f�Gj���47C/P��]�=C�f����+�����	�-6�/N�+fo,yFn^0��On��3j���8@�}C2��ª��U�+R�R�s�C.02uE�6������]�\��hEF�+��T��k�`�pJWF]JǸ���-:�?M��J=��S�zy���T�K37m;�R�7�JDe���0�·�n���9���2����T̗���'{�pU�Y�g�j��ZOeSw"*蚸��7F�ں��I��*��fur�ma7wk.�f}�,|�˵՗�پt�V�u-!��&�`�8��n!�
�Y��������_M�8��cM��:��Y,K�:�k	��E�Q��\jK}�w��%�WӔw�t��u�xRps��7~��1�q/���*�Xn���������������9���ka��6�]f��/Hiy�]y0�طysڎ�����5>���\���33`��v��5^ �{�ɰwػ�������]��?	��TKTT�yʳ�Q5Q-SS�t���X c�
��7���P���ՎhWBZ��l����X�p��X~X�V�}�8$� ^չ/���<���e�J�	�v��en�٫�@`�Q#Wz��J�ҙ�[۰gy���]��7�ў�ԫd��-�E�<���o7�.�����h4�x�m�믖��}��R:�tZ�02C4�-�Yr���Sb�\��8�7n�-+xp��,�dn�MoiF1���;���ά��u�����J�c�g�b{�}����,l������YۀH���];�C���K����Ә�ؾۂ�9�G�ў�l�6�-u�e��v��-�����J��E�=(��g]7�ޗ_u�,!��<-H��:)��L�����/��0;oh�B�6�����aD���]?y��2�E_����<;����M��S��,PY��B��lj�[��3��3Y{����Vm����j=AU�+x�kifY����mP��&�j�����s�K�0Ć*W|.��X��Ѿ�6ბZ5��E��k���sEV�#�q�h�����U�:劋�b��+X�+K���1�m���ڭ�l�SAc�����t��s�1N'F-:�F��s�&-�%:��0r�;\�˔T�1M;ji,f�ZE6�#���D�ɮF.EV��:F�j�Ti��g���MPm�W �	�clQ\���X9b�r�,SA��j��֒jB��ce���(6ŲՌ�:u��X�scXm��gns�MQh��k��V�Ļncѝ�i�skj�t�c\�F��hgZ6B�X�U�c��lVآ����u�u���ߤm�Mj��w	�<lk��:�ޑ=�F�x�pko��5�	��L� I:�R��l��B�m�1ډ�2�f���Z?X��q댔�o�.��@��@Le�{���~��o��G\{�d�]�W��cb�I���fݭT���J���͌���2g}1k���q����n}����S����ň@Oe�����K��B[e�;%���kAYX��x�y3��>E��d7|k�8+1�MR�yua�I̫{��=�w�[v���w�yQ��T��l���2����)�ɖ�uk���V���X5lT���̱Ƕ�{�'�{"��n"^R��o?Q��%���\	n@fcn=�]��dž�;��]�õ���>��N�6�O���}`h����ᐦ�嗿��L�=�ٍ[I�ztG���7����}���j��I���{^F��K��r�����'E_�܏zg�]*��`����f�/�A����~���S#+�U�sai̍��Q�P𤋮���|J7�H�~O����Zr��e���.�@�r�$
���^g ���⫉�s�:2�i܀Xʎ�p��s�^�U�^9w���h�]&�KH�g���.�zk�@�BZ<}u��k	�����q�û���~����C�ٓ|J�؋��ڳ��c�R�S��Ǜn:۽�9� qK���{0(��K%����-Yh������u�Awv���TI�Dt�b2�.
`47/��˥���1�����#k��9#�̪љ.`j�`bguGY0�q8"������'�.Ӹ����E��w�Y9N9�?Y2=�j�r��;'@�@�\K��
d��s��k�|�1^+�������yn�x��nMnG��W��h��P�*5Uo�O��T7��z��4}>��`��Y}��ϧ��g���su���}ʟ���~=U>��TY���z�Q�A<o�;�ϣ���e�e�'�<���,�~�Z�N�Ά=�<��l3;���OveEC��N"]Nx�V�	����l�K�\rP�}�ZU��V�dg���6�����s��{�g�ݛ;�]�uê�ږ~�y�Z_�r
5�cd�ہ���Z�����L>�����u���ȟ!��| �o�ѭ��޺��<��1x��g#�;����=���N��������Q^�[�*�H��G���~ӑ�u�{~�W��u����~��ti�é����`��s+�Ƶ���-��;������L�&s���;��{�|��7���ĥ^VT��!������1kd9�]�J=U����l	�W��7���\�Q��GI��;���k���Uzթ�u���1���ң���#�W)�ٌF��Ά�}��/tmX�b��¯^��D�+�l�=G�q�R�#�8<�����hyJ����2�ه��;=͕Z�M�/���^h����6�r3��x�����Qw7�ݘdg&цQ��w@�Y�uǟ^��֪Ϧ�G9�T��d��K�E�g��l��:�5�M����|��K��fEI�=Xkh.���:�j�t�O��[=��쪑�2�V��x�l�*����j)�u�ڡՏ��UyYc�{�H��5߮��)����o혔dUa11O��r	h�ǒ��-NO�g���l<M��7��~-Uɷ��U���������Q
CsG�GyL�0W��֭��w 6��Q�#�{�L,5	��O��g��DZ W�e��T���:Ӈ���^Z�v;))��!����n�Miz}F�8�4�L:[��É���7e�X�����Ǥ��zw�Ջ���'k��G�rrP�ͭ�����e�35��TB��v��}1z�x��c}C��^ϳ<�=u�W��}cP��>��G����:������>��tV�g�3�m0:}Q�ykԠC�n�F��B�Z���S�����i��EmO~���x3X����A�4�V�� o���B���hf�S�����t���o�5>���{�V��3�O�������ww���1�r��6�� � fzNF!{
)���kv7��-�ϋ���p����Np����a���iw����E�|��}�1�U�p����N؆]��:�t�v����]��,k���F�r|���gqr�3	��/o��kG7Q�I�D����<�B��Q�.�5�g9}I�x���z�+�;�C���[�%���T�A��e"�9�Vi��o��n�o&u��3}2���{
�K�]���6���g{jQQ��gFyE�&O��mW{t��ma��͆�� ��\<%9�ɟ/OQ��i����������Ky^�t�f���u���E��oz�[9��\�SȊ���,^L�}�ΰ;�t�t/Wgz��뎆w�'�;)I*gb}vs���W�d#�Y���>t�(��jW���i��Y�δ�}�ެ�I�=�+��y�l����Q�_�<0���<��[����>Ȫ�b�z��-���:��=j4u�������I�q��8T_�܇���8�|�a#��o��}��eyo*����9�΁1�]��%���=9\
��� �6�ɗDr�F���������oC��|Q���|�M����|��9�5��Q��,��g<}'!V��oL�{��˨U��UN� �5W��#��}//ò7(�W�+L��s�=��[�aן���|?W��(���k���` �ԜB���n��7�	�2����7�xi��.�?c��A���@��&�x`���ٵc�JU���u����Fb�=����!v�Z����MKζ�֧2vv0^!�>Ӑ�We�yٖ۴����V`ʱ}��H�KKw(�a�q���Z��A�@Y��ؕڳc�]T�vO�S�=p�	�z���7>G�k.���>'Y�g%�>AoD�?��������׶N?P닏zF��9�>�* ��X4��#���\{r#k4ü��ps�x��#��-�g�uh~u���,��u�z�=꡴n�����}A�ڇ��~��ٙ��[y�sr���i��<�M�S J�v�ҽ[�1:�<u\�ߟ�V�^ڞ=�N�'�1k���G�}G�n�O��څ�-\�i�����΀��:�V�\r>x�+��D��W�^�iUm�Жԏq�Vւ�������&w��'7d{y��t^����$�9F����W8j�]��B��,)�~��E��*Kg!�ւ�*�	���b�&u�'ȵ2��z�H��=5�[*��F��g��4z�>��+�����r��f��2�*�
<��L���R��7������X��^��$\u?^��#��^�}��ѵ����H�M9�y5�x\֊]��z�w�'w˸��`+=��&}~ڇa:H��w= `�LyNQe���׷��{�w=���%7�=m�a�0�&�jQ�oE��-��4r	8>�N�!��̜	=�6c�X��1�Ǯ٫�F\I�B�#�JY��R��q��b��C���ٲ{ǽ��˸���AGn��ON��s�ݔ[\�9���`��ק�� �/�̌�޸r��VmCF����?cgO���}�S�{$m_���W�jWg�v�<��I^�B���;$��u�s>��3��}��__�|M�(��K�7P��t��n��&u�w�_��~���5xO���6O}N{�FA��;���ޮ���]��7��Te��_���^�ف�k�Ϣ}:����?U� Z�����ɲc���:φ�}�����D	Y@z^���;�h�+���[9}C�r%΁�����5�U)ܚ�����a߳����ͨ�fw�H��L�/
�GS)P�+UQ��@yd��x�mO��/�B�e�q�ULLezc݉������g�omB͗�������~4����UE�������y����[�mڨ����گb���sDx�OP�N����h���l�c�3��~�^��C3� [�T��a��>�NM=�S5���s�:m�P���䡧e��ɭ*�|+M��o��j!;�蹅(,^�w�wfw��}�&��|�"<�n4���AF��1����m,�=h�G�~S�~��J����[��H�;P���-5���9X�2�]�6�tW8θ�j�3�7`��Z7�V�K&���eZ�M�eN��J2u���`b���\���R�w��A���h�d��ȜޛC��f�&WJ�	�������U�^5��{�r��ޝ�|]�T�	^W =�s~F�=:;�t��ym�b���G�wIY�T{Mb�`�n�7���E���ً���ϣfX�Ωw?W���#���W�4c��Ag��S7����Z;���7l�5����G4�7ц|���Ǩ����>�t����v�����g���s����w��^*��ȣ`R�@ȹ�sq�Cjr��p�9H�=���r#\�����2F��h�ǵ���F]]J����Cd{���R�Q)�3Y,*���[fq\c�k$��'�+hW��}�j�������,a�-��������2�V.W�fς��7��9��]���I	�h/O��ǙE��Hү=�W��sp�xO����ePe�y>���2����o)r*����(u9�,\K�s��
Ͻ���g� ���x�T)�g�B�N׻�����`e�Y��'Z��z#7i������K|k����r���R����y^�P��ք�}:o<2���5�g���=�D:�[&���>�q��Ba�.�͛�?PD��~n~���f�^]�?������ oT����1�4��Vzzʀ������m��S,�l�7{α7F�5�>���;2�	�;�������^���o6�x��T��F<֥y�u���89�
P*6�Yr%�lg]�n���}�^���7H.9Y^����d��cL�=�U�+������p�{=�\�Y{1����W	���~�_����]�a�CaY��/�)���8�5��/�^E������ս�2;����5��~��B����/�?c��4����kP���\��#�ގ���p�D^����x�U���G��|2��7�RȪ���y��쩱�3r���+����[^�z�wR<6�_Zu��ztr�=�8g��B��K=Yz�ƃ^Y����h�s#Fz3�p�&u�����lq~���L��b���k�s\����m��JUd{C���o��*g���\;ɔ�.2g�Ӝd7p9߰���K�h��|����b�Յq�*e<��b�܇��Y�"�����EU�1SȊ��"��L�}����i����OV�1����8v��ir�Q��˖a��%Ѩ>tyR.�e���]1_H�M����{'�)��ݜ=�y��%#��k޿dz�J�w6Ksqg�>�"��3�pl>�Y���Ōf����;q��cx�N��XV\���/W�>�)��6���E�t91`���_t�{�d�������Y������ɒ�	/��'�r��nw9��F��p�A]�zZ�p�2V�o0٣Z����a��_L ��p�H)�ɔ���������mG�}u�X����9�H��a_����ϣ��P�eO�����$������Wo\ڟ���Q����9O�d~;��r����s���_ ���#�ʝ��2+��=���Fد*#�Q���{"���s�w>��%����>�f�^>�������[��<p+ڥϓ5^z������$Z�=s���Dz��#c\�d�R�P�-缑���%`�
��91�J�����u %�Q����ˇ�7����8�<��q�?\�]�^��m���4N��j��ȏzA٨�9���� ���	Vn_��]1��0���R�^�Ꚏ�W4�U',�9�kj��W����"�׉�zd`�^�V.#�Q��}AuCt�#a*�R�mH�c>��ü��a3���	W�)/V���w�(�.d{�'�#��(UR=7����v,�9�J�e�+\V������y�α���7�=YU������t�؟O�Uw����7�{�R;�}��pj�c7&��'}1�k��i��O m��d�����x�鹶���0�v��I������f]��o�@e�}�rlQ�"�kH{z�0y����ҹ����2fokT�t�j=a������|�/�h�	��ט!��;����r� ��X�]���m5�*���,coo���@����.��=�Q����f���@Wc��~׮�Ϫ�&.{Ō'Y��.��w_�w�����P^��RGyO�v�>Ҧ������1T�ʜENUXS�1�̢W�����-�ގ�+>��C�Χ���~���:���wH0Q��P�2�[I�@�1MUɱ(�ݾ��R[w�p=�=�*/g�8!q��z��"鳐wkûa�`~�SnJ>o��옪�� ���nnK����:g�i�2.�W�E�/O�6��|a����9���y������gdo?	*n��>�9�'Ѥ��A�<�eL�'�kC�s6_�_uC-�����5�T�;���Э�U�ϔ�i��DLS�rb��>����V1N{�@f��P�N	>UEo�tl�G��
�Ϋ���x�x��]A�g�@�q�A�Ƕ�Y14�����Q��{���r��a���Ew��ϲ�J�sL��@�����{�p����y�5wk*<I�U}����D��1�)I�>����cEB�19ޣ�q	����.�o��B�ԣ;�e?C�xO�d�n�쬽J���\��Bfl�|��r�p�Nw$�-�m����'#�OCO�y��껴k/{�/�us婨���1�k?m�ө�����G����l��R0:/�c��qn_V��D���!�$ѭ�3��=��1zg<�B�-�8&ହ�g#]MZ��GZ��)�g���sE���Y�O%L%ob���,5F��[� �����*(�	˝��w�-P�)���&M���J����f�����T(����#�VU�J�A����7�w/��]����U��b"Z]��\�nQ֋ۉ�`m�i�I��n�XޱRs7w7q�b��n�4KG^���rB�D��\:�L��u��gz�Н���ˮ�Z.0h�t�̎m��5��9���n�Y����@ۉ�pegf����^F��:f��Z�n5N��A�Fu�*�⛺�	B��Xv>��j����k|�u��eMo7<�dF��n��α��V��
��>�ټ���c3�9��%�t�B���/m�״z�e.\���t��m�V�#�٥��]8/`]�y��������*�C;,I���-���}`�]��+�=�њ^zo$r�׶�8n]��Wʖ�J�$�r�����|!��8��3J�c��:Xͫ�7p_U�9��wGR�� #���faz����c�6�e �����g]I���G��\s���K�v�\��x�+�*2v�;:*U{,��&�B�7��^�^A<����?9�\��5E�Y�7]��[���o���o��,y>��b��}���]¬<�j��n-	�
<�A9�ړ�酬GB>gVoh�,���/��D/=��
❰�F�F����}9�C�r�|�}ڗ5��$Z)�4��Ώ��1p�
!��j�ڮU��%�E�X�Y�a�+d�x6�8�Rŀu�\�,�P!Ư�rE]ŵ��C"��� �H.��y����)1dE�|I���-��vrN�>B���� ��Z�V�r�r�q����
�̶�k���G�(ޖFr�bn���;�nWQ�z�<�ɛ�����L_ί�#B��� ��.�LR��[����������ἼD�m�P��Wb1�v�;Z���H�懲֮z�j�V`�Ϻ�-�^◊�;0*�3��p�T�]4D��	�:���g�`��1�]���[W�z(.�xm&.�D'�m�<�S�w��c���������2�<�"m���Ne,m_Aa
�Δ�V,ԗQ��ci���|}ٓ�i�4��nWeǧ �G����}�8;�t+Nfq�/�e����xIB�R{x�^7f骗�IN�����fǎ��\�MSI_>껷���ض��mĺ��֜k8n����)��Ɨ6�}����'xb`���X�.����8-M������@T�S��9��ŎKK�swHH�E��f��3�zb��LK���"iۜ�fg[��}�#$[u�p��huA�e����ᵴlA��s���ƚ��;Q�l颈�i�;h��˗"�+lLm��cUh��bJ�*������1r6�&�'cTUU%ѭb4Q��4cmE:q�T�4Q���j�F�M&�[�"�5m�F�UL�"u�F���b��Y��V���:�6uY�"�[h�rslgPi1��m�b61i-g�$��9�LU�EU�XسP[i�-h�cj�s��ш֨�:Ƣ6���l�6�%UQ[X�խ͋g5UTr4ѣmk�9kk*���m<خmG9��X�U��5E6ؖ5��N�ZM�6�EA���`�l0E�Î���1DmF4s��`�h-֎l�ڭ�I5�H���'ZJ$�����֩��8؈���,ɣ�[Ucc3Պщ�c�f6ME��$�ը��<W�X�ۊ�K�ŝc��]�jp�y�zv]�&s��p}0�$�H���ޚ�ߓU��je\�GSY�r�5����Y6p�f�m��Cu_�M=���Q��3Q�Ư�-��*��������^�7k�S"t�#�Ɋ��R�;����B��s�xj>���NW9]7��<N�GW�=p�ֲ���~�`���iI��r��W�ϓ�3�vQ�� �踟D���Qs�+���r7����S�h�˼{�wZZ���ѽ��逽>�:�c^��lT���g捝ԸL���N�城��/���Xg�*H�ܣ�0�T�ۈ�Z TZ�{���h�z����(�<2�zg0�ʨzF��a��3+�uO�t�v��3�o�>	�uHco���w�}�_��p�����BPW����Ʒ�f��ϲ<��+�/iB�1��=^W���3��/��U���x��{/�uj��l.�g�iZjn���[BO�?5DR�>��ȣ`R�S�Sq�B^����|����e{��u����f�U^�>��b���g!�5΀O*�]K�\��f���:��Z��/Y�.�b�P��
�[1�®�,�n��x�zKtKf���d�ϦW��^7���]W����u�.��q����r��Xԡ�j�����
:F����Z��]g��m-�fM@�Ӆb�	�s�=��f�J��8o!�(q]�:��s74��S�Ul�3C5; 3�u��-;јV�l����!.����L6�S��~��zֺ���(��������5
'�|�A����¯|fGX������۪�9�
9R�Yyޭ .9��èS�b���!����z�y��"��B�TGz�S�Y�r�1g�}�Ji�IϾ��7Z/Jgw>Dw��R}V�|��� .�������?I�HO����;;r'�$G�9��z7(�U��Miz|/�¤y�sf���O�^<2�Cɞ�x�OKc\�O�����uߣ�y��é۫�����N�4��=P���w���D�硡w^��䢏}��s�He���3�5��n�ñg�7�3]4�
��SY�]wG)���]q�ޟTs㓾��ڷ�Æ.;�'���NT<��q@h�j�ܬ����yW�~�;�B��g���ҀF|@P���5^
��e�q���p����z���.�5�ᵑ����S�|+9��)Fת=gWY��H��́��No�kӁ8�,�q��\:UF�O�3�{�{��V�<wʫF������UC�sӱ\F�g�o�~��r��o�ˍ�NCb�g����f֍�CG��f�"Ƈ�,|��z-��-��e�n-,���2�}!���<��Lz�l��^'\Ƚ҂;oW�FR����0^��;��a�@gP申��;��͜1e��s�P��5g1*�N��_��T_m�}t���/�gV������k��$6��`���o�p�#&Y����s��2�����sf1�Uz�S]��6̾Y�m
��c��q=����/7�E3r���U�G�|��cݎ}��pnm����3�A���qџF�=K�G�>�p�������)ٳ�@>ʨ����k,����Ҏn�F��׾�H:�w�.T��^���z�ڏe�!��<&=_�.���X��w5y����zVTU�e�چ�븰_�"��P�o��w"߫�p��)���P:�{�_z«���C{9�Q=�xr	h����$����n#�xz�C��0O>̺u����]���Z�h��
��xq�"��;���9�=�؆��Hȼ������cz��\׮�I�C��;�ʍ�u�"�Q>���ܢ&(��>���/7�;Hݔ�.��`���5k/zD��TP����s�1O�E�9P�6�>���>�v�/���9�ܣܬ��H�����4K�;��?P�~sC}����`ңq>�#���G��l��C���5°���?Nz���z�V+'~�'�ː�r�"�� 򮣔 �N�{B��{�}�����FU��n�����U����Y�'l{m�}�nll�f�������n�u���k#Ǌ�gbM�,��,����p����9��ی�go��x��z�b,���dO���p�s�v@f�j<&:�^���.5�����P�m	�\�,�\o���w£њ{�Q�Ӫ}�w�>���0�/*����qԀ
}1%���|�ݺ�Z���tD�Q�\�27i���������TB�q;,fN�.�����M�ip7��+�~;����ѧ�/X_O�~�G溜����z�W�:p~F���ui�����ʥg��xP�Ep��D�&	�gT��J39�t��~�����~��Ի���v}U7=����Z|)�w����]>S�zy7�F�����9��O�S�WX�dGTf�v�D��⫀����Sx��}>�z��ˌ{�R7�,'������{O����W��c"
��;������F��8�j�O��5b���f�-+}�p���&�x%�Q�}���f�&�S8�}۵9�������yϽ2��D�R������[PѨ��I��9�Q�D��5ޙ�V��=cѪ�����Z$6n ��eL���q��P��O=�2����Ȫ�{�Y��n�A�Gwu�W�G��T~S�Z������[*��O���=jm��ڑ��R�{}���дՋ$��6y���4���_`(��t[؎ ��1�q7��b�LKx��88me��#/n���g�x`��̮��G�O�Q���\���$NM��Q4�c����{ޢ��n�U��&-xO����L�9�ta=�^ʚ{�����������}D;��9��|Nǽ8����1V�āP�KF��=��Ʌ�-�ܞR�v��̪�06��T|�xw`����O�%�qϨyIg ����zj�U)��O�j���y�gH)�������������X��,�Q��><� {���²���{�.�Ne�ӛ
�˻g��}=L{��U�iϷ6��ٵ��3��ƺ�T|o\�2����c��ޖj��3��M��z$���,;��\zp:���q��_i`Oe�#���g�O\�ק�Y���Mf����i����w��n}����>º2|+Mƹ�}g�leȞǟTk��܎��*��z7���g�|�{��fTWo��E|���Nz���ʤ2�&�Ĵ����m��m�ž2w����H�#�B��:��7�#;�Z;��C��x�>2���a=�J��(t�Z�(��[N)n�h����n0���Hco���s��#�~��^�CFG��i����߰'��`d!y�1f�&�����4!7��v�2F�5�B��n��`l8���+��Pt�1��u5mi���!
̥�u�ɉ|��拨s�4%�Ţ��:>��`�t� {H:����z�_R�Rɤ�#J�IV���=ݘ��9����X�A�y�xg�����^)9������#}����dz%*��>����]˽˟D��o��H�@79l	�Uk���	zs��㋤�6'�3^��M^Qc+��ƍ��V�G��~\�<�Hl�:����W(y��C�v�U0��Ӻk���x�/?{��ұ_G}�g���'��5��9�,=�#�&W���Nn��B��?:��7�9�ŏ^�0���z�U{���\�o���]��NnD	�7���q���9��~�e�nӿ}�ܮg �{;����1�my�<�����q�f�e�c�?U{ok��!�g�zH�)��11K�EƟx���g��O���3���.� �]��;k�T�=�������wz�
��Dv_�U�7>ܢ_�d��^��/|�L>^��'��T��eL�G{7|ԓ�6Ͼ�U��t��S]7�#��y6���j6^�'C���;�����W��l<��}��;0�蓧�ު��r��~����3�z��+�B��<-�u{����[�}�[�h����7M��o�|�ܷ`'p�;Τ{��Q�Ԍ�Bl��3�%�Wi��}[o�u��n��M	c�|E�qf��R�8�'"U1�x%@w�}����Y�D�����q��a�w��.�1�dJ'���w)r�dλ�<Pʙ������>��i�d1���
�^.oޚ^�Y����-؝�y����n�~�{q�Z����YC��F���q���4�	{+�>�I����B���Z-{Mt�O�mOY�ci7��?!� }�������W����􁾸��k9����h�'hP�r��3t����u�r��y-�����Z4�Ȣ��V�;�&w�z\��φ�?XnS;�ѫG����&qdz��f��u����mJ7�=�e�:�
Ȫ�&���g\����9��c>��ي�����>xr�ه�O�|kޑ�C�Q����f���n^Ss�b���ϑc/2��k�7����j��*{��{�J�{~8.=���|ϴ�V�b��[�YHfh������ٻ9����=>� yd�*��Q~�\ՠ�q�����z�q����<%��W�Q>�S�����=�\ϲ?ET�;�E����چ�-ZE��_����<������֮A�{���Ƴ�
z�;V�fVϡz )/�gd�����/Ԭ�-͘~*/���K���G�+�S��l%������z�w�&�R�{�T���e�F�+���G�aĭ��j���n�]J��P{K���:O.\'"#���c��
�䶾5��=��{���x��9�OlGz>Ψ8��Zބ#�lv�j��E�y�$��*��Vs�+����Y&}Do��|X��S=7$g��v�� ;+�£ݞc������VֹQ���>��q�7� '�)��H�TCG�}�����1NV��}ǎ_?(��T�:-�u�O��!����=BaW�N��9�)�s�=@��z}$�S�t��<���/������Z=�.�ϐ�>y:\GSJh�*7��dc�P��#'au���J���;4�1�劯3/b��8ǳxc��m{��zx����Wu�j�,��^'�鑞=pՊmL�*�9s�ʦVyv�x鳲�};Q�s�1�ͪӡ���u0��_�9���x7��.2<�Q�����Y�]��{��g�Os$,;��d�B��V��,���\����|��w�+,���V����&&�-#��i����_�l�^ڑ�} ���Lf����}�F��U�b(fA+�]�LM�y�ܰW���i\�S~���q�{خ<��F��t}��'S>c%Ya�����m����G���o�p�yg�l��y2_;����:�=���.iTc�T�Z�S7K��|������Z��'�-����޼~E������;;*��>z���n�d���\F]n����_pĻ>�<h�&�!�F�0Z�֜�rU�����d�x5�A-G�MG:����kW�O!Zq��@<�V,��i����z%3������0R��!�Q�	�ir*틔����|�����?x"X^]O��z3��y�yW���H0;��Ƽj.��؇�2����y_/_����|y5b)z���d�.7��C�.�9��>��c��};̯z���N�v���*.��+ʨx�4�9�L�NE[�j����h��چ����bM��;:���K)�4ϻ�Wu��Q��]�������T��U�sax�FϑSޟ=�4���׾���j*G_����8�:�g|F�~�!ź�%��O����dVYN{�Ef�5��W�Ӭ8l;�==�P�j�jg��\|Z�9�N��=��������1�?nz�ށ�Z$��&=�����_�|1��[!�G�TK�\{ِ���V�KN�]{ϓ�+�5w�XL*�[&���>��0j�,Vj��9��ຠ�}�qӛ�Nj��OlV�!KBӕ���s�J���W�����y��<��u�UK�����<�:.��������r���uZ=��7�8��\�����a�\�tޗ�d֖�B�UZ�j�9�o��8,?s�
�)�Y s����V���G����>���h��]����l2(3K�*��p[�oC2���ܳ]ǆ���7m�. �wũ�Ӕ�ʜ��V����u����%wV�^۹ṱX
�Z���	���qY�9���Z8yW���L��{��}����D��;Le����tV���z���U�#����ù�Џ1�W�*��`5>ޟveE8�mΘ����q��Ië*�ʵ�f�95��L_����[�Ӄк}gY����i���o���y����F1ᗧm��R团��n*o�.��F_q7��5��ɝf��w�WA�Ľ~Ө�����^�c�d�󽘖+]���X<R��>�ғ*}����o�p�6-ς��a`S��g�V7+m�f9���OB����U�я�S�7�E;���r(�\�\�9��,���bx��y��vW\�=f�{	�������9>�J�߆ʔ{=�C�g΀}�UH�偗)3Z�+p-Ҁ�z�7�}X�ܦ�B��Я�~��c�)�9�0�z�q��S^%�����ޠ$CSM@�������/߽���..��.y�͟W���:w�X߽�L�sfpmǩ\H����p�A��De�yX��t��:ŪKA�>�i�R"K�\r	h��	�1ӺP�Rٿ���{"�����#�����
"+����
"+�Q_�����
"+��DW� �"��DE������`DW�DW �"� DW�@Q_�����
"+��(���DE�������d�MfEϾl�~�Ad����v@�����jo��*$U EB�((U

�T(��EJ�
H�  �5�©*DBT%)RJ%P������*�T�*(A%*TD��VW�����$$J�����)JH�QB�D�JJ��*�T�EU;��I	% neDh�L�PmR�
��
H�)�KcT0ڪ�cPk��PR� � ��M-�T2�)�ۛ�M �`  R�0 ��   �B�����Შ��QPU� ���KM���4ͭ�e&��5�m�[j�C3UR�`4m�B��l�	$X�4�l�6�����e�e6JSJ�-MA�XA���kCMIH(��j@��tUT�)*�2F�mXm#3���0�BC3Q��&� BiJRƒ%)�U
(8�uk5��,0� �J���Pa���VZR@��࣭jF��M*J(@QB�����B��lU�R��,օ
kE%mR4k)R٫f��%4J�
�R�X`��H � ���0�h���U���%�dԢ��$�Z�����P � s��j���5�T�Ci�Kk5HV�B�fhe	�BkZjVf���*��8 �Ru�@�aBF��&�)P"���h!�X�F�]�I  ��L*J�Bi�0A�  �bb)႔�C 0� �  U=O�zd�A�  �@��@����F�Pi�d4��JQ4�i��M�05�h<#j�H�
R@�� #� d�M 33t�,]SJI�	1jZX�%�%�V*��Dϩ��G�(��ش��J�K��#Y[�~M��h�Z�#jY�F����/��[���:��0d�d@��0p���*�ĵ��ebY�n� �1o��{7��Ӷ�p���������Ͽ���D�飗;SK]~G����͑�T�?�N'�(%,k�x�JJ��E���k��X2H������*ŢX���"�;i	deef���1��v���W�ٙH��޵��°gQ9|r��ޞ��J��(�sc���*��[ݒ�9y���lQ�4�5�o-�v���n8�;���Y�e�0�d�j�򜭰��R���L�y�*<ʹ���3L8�M��H��N��N�u����n�b��7����:�;k-`yϩ�oM�W���O�=iV�#)㡦�4�#6�Oq�X�V�5\�H��PSh)��mݱ��7RM̺YQfe��|k����7F�L�B�J1iM�与�y��2�]Y��%VU�̢Ӵn���괫)��R:��@�*���v�t�k�T���԰���a��bv�Ts%�Z��5�[���Օ�4�6H�[f�ԤYR����Z�9���v��3��F�Ut��9B��%Q"��	��1R؎��mR��.ZZSX(nX<�kn��z�o�a:,[o1�9mݲ�g��Y��e\'iF.Xr�=�ۖsS��l룳�ω�'giMm,� ���:��v�Y��W��qҵ�6�_a�wEbC�v�w�v���&��x�D�	 �f킝]��}�w�S6��e
�f� �:�k�p�k��m�{��4�E���eU�%�e%U�ŕ�[a�;*�J�4l;=ۖx�F���֍��4n's)F)��ḳ�k�_^��M�a_�X���BTa�C*dF�D�*�#��w�"�Zi`�F�� �QU����#w
�i�9Y6m;��,�%��@������gz���wJ�^�
,Ӂ�[CtI,�#k�5fm�O�6��r8r���1�i�u,3mAkM��2�5���$�r\��3C���c�!�i�㳥E�,NePU��w�bB�,ؙ�
��ܧ������Aƭ$j�r�\�3r\ͣHQ�Mk�Qk�[�ӥ -P���#E�1�fn��6�����Z�'8[���x��������ݛni*7O��uu����,4��ɒkf����ʥw��MX�*1n��T8 R��u�����m�U�w�m[w�n��
�����b�+��Am�:,T�F!Zɖ�;��d��W���Y�M�2�ɗ/p�q]�2��I���(�A�MUr�)m�M�J��V�Į�U�	�0��z�[�N��q��I،:��F�����pM��<�·�����$'rأ�&�B�#V��O-*i�ѷ�V��d��4v�Rن�V�<5x̉-_R��Jnn´��wn���A5��nhNɣ%��&���t;�o�FY2�d���0�v^��L�6V#;N��ow9j-*��j����e��I�e[�����`�i�sh(�A�>�F�]W��lbA�a�� Ρɫ{zRq�P�Sot���n��M�Ďb�L,�j[�u�+a��r�h���&��6��xD���}�Ț�����4UpF0�
���Q"/�9(�^g����ZE���M������(`0�[��%d?�X��z�ݬ���U�%齫?P�]�,�5�$fɖ%´�{Y5��'2��R���C!�PCoY�OF�P���;�0陎S�sX�E������Sj�V+�X�[Z��lA����8K��$�%�ѕ�ݐ�l�Rn��ݕi�0l�H��.v�r�1\�r���Q{5�Ū����m<�}�u1,֊���J���Ӵ�ژ�RzJwj���:'�OhI���h�-"F]\���-�\�>����Ѳ4���geM�еv��3a5�I��䡴�Lރ�Z�N�+��Wؙ���2��l�� �m�ff+��۳5�[���iJl8�,q�23k���7+`z����&�#��V�t�CG�ތ�Y� *��u�,�\D��l�v���cC[�2{:��:�ޫ&�*�u�[��/2L��M��vi�VhC�:�7K%������'��֛«��e�%n�I��*L;�iz���^�	wSzY��Xum�F��;�b�,�Ѣ�nf6B�jPPcf�\�lk�9��&L<6�P���Sʍ�2��p���_c�toZ+祶u�6�f��9u�7AK���,'2NM�(3YW�֫�f�f��M'a֠�Q����5g3R̫a�����UgL�U��<�ÎHm�rť�*�{���S�U
�C��4�vd�UU��',%�6�ȅ�sb�*0c�v��t��5��5Ҹ4[��O��If#�����$�uJ��;�yv���h�I�7�Н��6���흧&*mǹPon��5�/p4��l��5єdGS���<��)��&�3��ۈi� %�֝��ؕ�Zr��.T��\L�Jv���wvtf&��
��]�D�\�̴H��^C2җ��vt�TN�e�uv_i�W�y�G�Z�K��Mp#���层�A����8Q�E�n�fOBr�e���aUn�քX�sV8嵌I[�Kw��W�B%HOv�8!��0^v�"�	ݪ:�҃,a��i���9����ڻ�JM���3�:K�5|�?'��'[]v,�E��Ԙ�Ve-]�"�o�]r}-�[t�<B��ۈ=t,�Y��k[XtqY��|���I`����YT�y���呫U٦�횲\�2�|fQ0U̽J[�T�B��^�G'{�OJwWK��gD4o�t4�n�6�-x�ᑗx�	HZ�sq�Q�W�M5�:ۖa{[H���޺��J�f�Z�h��QDnhɢ��$7j��ך
H�E�DR5J�����RzXy��Y�v�l����TF��6���ߕc�0� ���E��[R�h�2剣Ha���5��5 �,�����e$�qZ����l��VZ�)u['���j�^�l�v��R�D��sPv/H.Z�5�+b��Q��W�O�g ��B��W7k\��)����qr� j�<ѵ�@�f�(�o�N �tn�������ю$����ͩ73l=�t�D1WF�������M���K�H��,��I�9�[zU�����%���7�u����;�^^ౠӷAl�Ia�M�t'fn�<�̳34f�ndJ	G����ae�H �q���lٳhe�cr��F([��*2�֫OԨ'��4�%�x����O��5��TŶ�Y�Gl����N��w°���l����'Q]%��Q���=�u�u�6�k��J���6��۬u0E�jh���b�UةYh�Y-X4��*BV��M�Xm�F��U8,�6��LaZ�ڧ�q��bX�0"^�T��\��<��ө�z�f�Z��v�X�}�'.ea�w�o~Ȳ�՜X5�����CE��
��fW���s*ʋrd�u�[	�Yx�-7\��5ܩ���n�Pb�E,�C�cE�y&��/�8&)*|�{z�a�p���F�Kiܴ�yX�޺�5����z�vo2D2RE��QKl=������ӫ�i��&�0K�ő-��J3V����p^7NR��f�@�+C\a:h5WE�w*ۼ�a��%`��շ����7�RB�^�U�j�t�MY0�%Ƌe�meॷn�wx�P7Sen!���XNfX�4���F3)�uA"�[��bqUV)�O��o��i��V�Q�.��4�B���c2�T����|���Z6��T�q�/��/6�ە8Iץ�u\6��v�=I`�ae`B�kɳ���cl�%�4�MFF�1edܙ��a-���l�z5Е������P��!�i������wy��F��蠻�I��Zx�֒��dm�F��d*[j�q�Ʃ�iwtA��9g-ʪgf�qX���K46��6-���ٛ�+s*J8.<Ld�+vj5�{�떅[�x��;Bݾ%�U�e'�޷&�2��kN�ʠ�/��-u{�T5N������ �� >��J���g�.���aoI���������!��>��*�c:�A�?Z��?LϾm,#8�����������6
�N̩X>��IW���y���^o��7�NU�Y�!��&I$�I$�I$�II$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�K��$�I�$�I$�I�k����2��ut���閁�c,�
���h)-sz���y�;��|�<��)���)��zD��X�cC%�6�ܓ.����sч9��y}7�]�[�g��M���s���CV������4�Z��bw�Z�+Hǡ>N^u���.D�e$1��`���v2y��v�a�Lo�y�7�����B;Jg&yV}�p틣6�����gi�.b���Z�F�%x�M��e�E��;X]�Դu�Gb�k��g��P�qQ8���0>��H�Cp��{��Qr�K�1]�|������"����Q[���[Q8Њ�`έGj�J�2���Z�fT�cBɲ��H��ث�ƛ�2�c2��oY��T����%S�6�mL;����c�&d����:t�.`�k��x�9��7�&E�5�z+�+��T5�<Z.�.%�4ج��lf�ޠ�Y����Md�̥�wb�,UrU�
����Kj��ܩ)�,����Chl/���B:�G5V�M�t��wf�c/	V�X����6X��1ȕ�U���W9�L��D�@�XEީF!sܪǻ�g>B�T�[\:����{zz�X�\#h�T�4@@c�h۶����k!.�޿�ι�3T�4�f�T�unW�_Wx�"��4���)!^]5e�wQ9��jZv`�{j��Y�U>��t-�j��r4�6,r���kU>���L���Fi�*]A�SO��8"g�ŀo�3  �E�q�����.9�Hn�x��eJY	�Zx����#N��K�n���˹�k�"��^Y7/�.�e5/گ#��c�\���f��b�+�������J��1���[`��mK�<�n��VÐ!j���竨�k�m�g{��ӧ9^[q��#���J���mE��8��]骆�u��O4�T����<k���ٌ"���-���:"��"rhE́ �*���/����5eCR�ZEU���2�����:���pS�q�'�5>��44�C��ru�LV�cw����s-�58��r�n\߷����Sv�Ϲ��tE���C.i���I{t�i�c�ق⨐��MX�cXe�+4�ʁ��z���֥7�2��XN�Xj�g#�Rk�[ԣ=zn5w��{�nMӁ��7��I���4��*�!���X�{q:�ꛄc�v q�:�!ep�Y��:�q�m��z0��Q�A���}'Ne�5��ʫ]Y@�l<�]P��S�M���� gv�&Ȣ e�/p�Ǩ�yتm)`�ك)�%�Nщ����ϝ��|f�'~cr�<�Z���hf��X�էFֻ�O��ru�[}H����#�fӤ�7��T\l]ע����c�k���:����_jmb����z�ȭf���5�>���]f���}�z��B�ھ`�W��)D�.U�p鼓"��w��.�q�:�:T�AۤD�P���]e���1ن1�vD�Mrg�=�U���t�f:{�v��r�!�p�a�0c�ͽ�-=�.�Z�q�����׼l�9�4���ݷ�8��ƍ3R�0cA]��[U�(�)�+��ښo���n�u�C>q��4f�����ӌp}�6�ܙЁZ.���p��w���d:�흼uv̷����密J���O\���wA�.,�0����e
�S�Q��̈e����}�4��{+"�i7�S�T�M��N�����s2�G]�7��p�(\�03e_ӴO�Yͼ���9�f�'$�H�uKjY�d3�g���c�٨�l�wfS+[�Uc+��&��FD_Y�븊�N����g�v��XaQ���ࣇH�
��^����+�_��]>evG@�)���K�h�UǱYı�����
�w�R�9)����+�ti�I�i 0�}ו����3xK��wS2��m��mqZ�>��od|�;j鱝��O�Ӑ3� '2���$9r��9dq�Z#����/OoJ}�E�bvS�<��+�"J�h��� ��MN�}��4�+:L�3RSb�h��x�A���|� E٣V��31J���s�b��d�Ɗ��T��\�ŧ�kt*n֬3{C�v�t~�(q��wjt�XH�zo��[�p�2+�a���U������5&���	Iv��}8N5�d�GN*�5��v,=8�GGf��9�v��z�!9
<����L¨_S;�UβV�ޔ���U�Z�hG;]U�~�j):�<U
��﷡�K烴*wL��",�P�Ӻr�xk�M����t9�H�[Z���bҰx��t
u���G�� 7�>�Ֆ��Xz�5��f^�x�ܑ��ViP��e���p�X��W/�N��W�+�m&n�[���rť������Ղ��&�l�ّ
�6�r�����E ₻v�H1�dR����|�Nأ.�r+�4����s�F0_`{6Ż]rMw��	� Ι�ވ��>�ݪd�Wl��\(%k6&�#�zt+���n�Sn)�N�ۣnV�Q�Xp뻘���I8����d�"n��C^�p��%yQ�]�����DdL�U�c��΅KZ���{�^���sJv���i��~�������Sd��E��u`�urt-�)(��嚞��oۖm�F\Q�qܴċn�j$��1n���E㧢�O�70Η2|yhR�4���^���F����(R:�=����l�ǌul��-]h@ؘ�;�u`�o1/kւ�h*�nT�82H�mg
L4�J�En��Y�ݳ�Ӭ3t�RLk"�/P���q��쪕��f��]�9Q�A����y��Bd	C±�����!��ۙ�Vvؾ��-��E��y�&�GR�m�i����S�O/u�ڶ��E���J8j�#�
�t���9�b-L;,G��f\}8��h
����ٷ[�;*�dQÃ)��'5iɧ
w/�U.�:٭�jμ֡p�*�r��4�iz��.��X�m[��k=qkv�����<L�}}�d�r�;��g������b=V�u+a��do��iloCppin	L��sŮ^]�I�n�py(�kUt��ƣ�Ǫ����g�����/(�4-��͂�"��#}G5���J��30����0��[In�E̬[0Qv�V�Tz�s�st˶��=������Zip֚��}5-��� qI��X��7d��oc�/O}�HZ�Pъ����TwM<�B![��G}(U�όÂc-�o�r����B�Zv��5�p�{�@�<�j��dD��|�AM�8�\B��\��|�%�P{���{�)\�kw/���^���{�`y7]eʮMV�8b���N��AQ����:���2V�l�:Va����t�^+ϫj�wn쫻�4�B��q�+X��ӻ*ӜAu���]��A�w���\f��n;amr9T�C2R�J���;U�9B�!�_ΞM���Z����p�2,��F
�X��%���
�;�5[�4m����/�����R�%_������a)������">c:M{�X��hH��$��V+�e�%�H-��v֧��C�M:��#N�8p�ө2�u��!|��W�U�.��9��f�ءZt��5�F�8�b�Lu�����C�r�r�x;�Z��.�}��.(�W�&J���/�V�:M�w��c�l�[wJ�
��!�(x��s5sAJ����3Y�#{��9:V����+z���5u����am.��$���h��y7��&Dn�3�V�7�';�۶�*� ^R�vowZ�0�w����t�p�2�;0l%W^�T�'(�L �$���I0 F �JJ	$� "I)($� ` �$����(�ɱJ!^9F���C��8���eh��V�II<L �?����?�?��u\\y�yj߮۲Ϥ�g<�۵�%�{B���~9���h�=��( �������~w��g�cL�pu�Y�����ט�Ч)���Z/������p_<=���/m}���WJ�Mrk��N��ˣ�p����!��M�:n������0g���#E�3�R��>�g�2y�K��Q�äۉ����sv����+n�c=(�l�N�33Cnn���6���Ya2�8�u�
��VkM�uL�S�U�X� �v�hAv:���&)���K?>���L����������]`�2��%Ϭ��q<y]���:#}���ǔ/���v���@�n��u�-����)�}�E�׆�Qݝ��:�<��T��ÿ-0^�7��Ո:(�q+B��m��0�FɎ�����Up��Syh���.�\����u,ϻ��gU
H�o8��c�f�*�i$F��w&<]y�md`��8#U�C<���4/_[.k?b�z�	S̃i��2v��Ϧ�rl���*j���*���HhPܱ�m���Q��CP㶳Rii�i�i�C�a��.��[�eapCv.pL�\���XO�S�,��7㝷���/�+;z�\��O\��n���.�B旼IB����d�Hw[�u�8�Oi�w�n��:`F�Wp�iG�ۡj�3M]l�-�l�r�'׉'��6��
۸���:��s7f��襲����:8�o��2`&�� l�^f�B�Ў��<�f��w�&B��s`K{ݍXY�F�Ǌ�vZ]��=�ic�6�}8����U��\MD�l�T���H�8��¦�J�yq�kU�-'w�98�\Q���u�&9���saCN�e [����fe�4�`��XG��hv�<���SP��y�����݌�(�ЉL8k4:y����:����>����۸��k���u_T�+Yѹc�����<��ɵ�T����˪�R�;�
����/C�*�a;r8*�,�AX��d��]+rRZ���y+�]8^��0�M�	ޡ�k
��2�{��8s�h�t��UQQ�x���2�Xv�dd��vϺ��;:�I���ZXB�λ�T�<{��R��/�Z/�UIj���f.�zyyȷ2�jm���7v�s�e;��3�E��ZA6'�`�L�39���F�,0iƞ[��zkp�8�l�Ok��GL�i���e�i��"w�`��e�"D���<��8��f.��x�I�gVr����(u潲.�n��*.z�L��_]�H�O��YN��$�Y���۹�,>$_��ǹ�i�tv�cܨn�3�)MY{EV+ί�ηF�rK�`]�7���ز�S��v"v��&�G�l�T{f̩���D��[�#�I�	en���z8S����V^��u�R�	��p��E+?+��q�7�j�%��L�:��=KSQ�M\�9��ɲЖ���e��R�*-��Ҏ'ٺ�B����+6��'�0�P����V;i�Axw���w�,fT��k/��v��R���Rp`L�C�<�a�RXU
uw)GW���������T�:V���k�wNZ֚��[ߖ��H�����@n^n�l:�꽜E�u�|Pג/���ϣ 7.в�W��cZ�X7�հ�37�Z�7_3�1���z�j��OT�E!��૗d]�M�;ZOK���<:���ͬf��.��yuLn[9B7|"��ԡ���	�45�Z�.�u�W�[�/73i�Ġo�T/�d�Ͼ�.����5 0��]�TڟZ�5S���5�V��븣�&�c
@�o6_f/-����K���u͊mH�ZKI�_b�+v�n���7�#Ƭ�k:;z)|sq��E��Lc;��ܱ]8�&hp]�u1eG(Vp@��ѣ�oj7�_E&��;�s&O�4rc�U�.�Y0��d�f�����L�6�;�	7�+��]��h� ����%�Jm<�b��.�fQ3�]����G�~e��;��2c׽J��q\6��;�K��T=lGTFO"�;\����m6�������7�uO p�z�,�7��O^�I>*���Qϭu/��s��/g�v��V��w�T	U�Ԝ�j��
��ݴ���7Ɋkn��VT�z��{w���h�fUѬ�75:���b�]�]�kxS���9,����-Vw�̓9X��R��멘4f�j̠j�͓�9DG�B�_#�yˊRY��v�X��˜(c�iѰI��ƙh�,���x �G�ǹ�NQ�7X�ZJ���Kc�z��V;��Iy�v�h��e��1����fb�}��c31��٬��sEn<�3�Ӿ���eq�g.���m��v�dϴF�C���lVt��`og�ԟ)N�\9��.�6b7Y�]����
ϐC_$(a�oG۳\��e9�9��p�$�l����4���X�և%w`�/��$�c���k!�Y�Vn;ե�\'��̺Ȩ��9CVWa��;�y7�<1U���ġ��;�w�;�e
��A
SM]�V�[zy6��yr��}[I��)�p���{"hw;�d�>�5,�دy��ԀbWL�9�Y��BM4o>���mr:����ٮ<��Vm�8\�>*B7L�N�%*6;��B��;���j��.�b9���d�C�S#+�{3��YN�է�NFZ�'��*�aDͺHoدkp`��鼬�f3OU���D۾��hb,�yi�r�AQ�v��v�5B�f��q�Y��}1�����W\�f�����%�/�ydY�rtӌ��F\ޔh̀Q�%Q̜��J᩵��Ԇ��:�f���c9�osNo^:U5e[wWVsl�z���9�u`y,�t��v�:�K�G��nq�@�tvK�LX�P{��*�"trm=��,�*Q�֙Ɵl�5Tc>���Q����h�	��u]_"k�m^l�YR���*>×���NT����|Z��NA��6�}l�¸��.��"���S#��2�d-r�z-g6^-�Ua͠�~V�v��Ty���WX�:�,�A�����;
���'jx���IH�tW>*n���2�t�ĭ^w!���5�Vz�<w��ʑ�� EC\����Hh�屲m:��UK��)��Dٹz(,ѮS\�f|�*uWcI�SU��9R63F��jfT�3���L��۬y�U����鴌�L����J�r�A9�f�X�<�Lo0y�wӾ�1mv3Y��r9�X�g�T�=yDj�B��lLr������X��s�&+LN����Puݖ��N\L�f_����{s�]ٙu"�'&�f��5�J̺��8������'}�-����7�d���TZ�j�����JS/\�r@y@�Y���5���`vz냩JQ�+�&�B�����
��cY�e�K�go#���<��n=�8�xha�u'��l`���˽#,�z�V���\�.�ńMbW��g �Q��8�H��{�jY!��V�0�^��Nc:Ѵ�\���j+
����7+J2h�z�]�q�2�	o�������ſ�wl����L<�:J�u\Y�ʚ0�:����w�Xk+�ˠ���[���:P�
g^g �	�0�Z��j�3���IM�lw�B�r�d�b��M#�$��\�
TT����fV[�qk+n�.�6i�Rv9�k{.+�\��V��z+��F���T��uj��f�!K��Mb�ɥ%�!vU��6�x&^wgK��7rV��{�0՚Oj��c���+H�8��EzH890�'N�R�N�[��m��bW�B-0�T�P�;]�U�b�0ٵ�x;�ti���{���j�:;q���.��[�{8���jƴ��ne.�i�<0i.�Yk�V���gJf�IZsEaL�m���$|6�D.F]�m��j�j�o��+�?
�F�P�=#h6��_	-弪��F�����#f#3���&bh��p H~�J$�ߺ�6?��w�Ƹ��I$�I$�I$�G*�E�>�H"�%Z���c�˽���s��]���u��V��v��X��cz�P�j��=u�#,��p���βlm�ܸ����RtpP*�s�����9�t�N�W�<Sp�e�3�j��8S[����u��^Ya��M��9|0�뉷��0��`nP��^T��V�0f�ȯ��e�AEd��ͺ��%W,m�t���ۑ�\��˪5�+��}种1	.���s˻qV�,�tLG#3�l��ے�KG��ۮk�*�4�>��Y�s���6ћ|:�k]"E
œlps���[������閚�R�v�qʴ�C�rR��U�%*�-52љ�M����i[ۏ2�edCV�X����g>,@�i�ݍ�{{�#�(��;wo�$�C��@i�:c��Ư���]^IdNE^��Y���wK��V媀�Jݡz-O�p�!5��3YB�T�d��u ���ۧU��L{_e��°��=f������X��YidE�
��S-)�� �����,*��438\����a��U6�0H��D�8�Ld�R��X`�X�l�����*��c-����fZ)l�ĕR�+�2�˔�֮2��C��"���UE�%a�b�8[FT��+Y*�*�0�,��+R
�6�j�"ʺ��
��T++Ri���[j
�YD�����b��%�,�TSܦ�HJ�/)�Pĕ"�(�U**��K[�V�jJ���C�o�gޜ����7Pr �Lڷ���c��ȅ���23/��P�foM�����;�g�H�j�lQ��m�P��0r�[���5���5��3G��ُz^Z[X��NY�L�,좇|L}��df_�¶=��^�Wx8�y�}�2�`m�mhA�?7N<{��N>{�{^��<8F͋% Y�:�
��c��nr�B���e�t�`{ͳ�<�T�3�W����yC�ƴ��w�����h�S*���p�,oI�矯Od�V3��T�V���U�����Q�w��F<�Od�c����=�Gu$%b���}��h]�,�������kit�:'N��&h.bL�Dի׵�*!K:�4��p����
��;���<�_CmPf�S#�g��Ex������F�(U�s�85�9;�NV��j�����i�d	����5&���t#��*��ղ�����ls�[��I��u9��r�8��05���p��ɮ�'����D���|^G=G���桊|&qMTW�{b��L�僉C����+D�ɕW���>g���[Y�9��Tnhm;4&�"�.�Tc;`mG;S�T��W�T���cS�t����2��7��-��P$�
S�'���q[J�Q[����ǹ��J��1�.a�t���sN���f�#йn�[zrK�[�2*}�޹���Z��·�N}Wї%�vVVB�Gj�����jri�I�]�s��Ӂ��0��.�G�I��,`�;F�LK<�vqHe�=�U�;cኟP~uԩ�M�^�h�MG��@y�4��]�0��Z��8�����h��=bI�y���O���V�2����I#8¨�M��	}��Xj.�ޤ��*�i�Y6�Ɲ���g%�\i�Թ�b�2v�=�Śy�x��L�+{W�����3�k9F�.)�V���#��Z������,�j�+���pM����R$$�2�zR�$�����}Gq�HB;\������Y���o��N'{m���Nc��4E�A��ꩵ9H�����m�o��1�DV���F`��0x!v��=n�+Z�^���v�:l�Xg���j�m�A�@]�6�܏]f�.�zj	L���i�]C�D+��PJGA�]��N���Ol��s�.1K��Qb�T�P7]����%ᕭ[���Y~�dY�3�˷1W���[���;JQەnű�����+T��yp��8���t��[s���m����P�¤<}������wh䜔+3�k�O;�6��w�r]Q�:n�wbէ,(V,�w#uC�sTmL]��=�KL��'˗w�o.rt��f]�11��oBX�>�V�R�{�T�w��~X,rs�]���q�o�9H-{��г���<�\�(��&���t����K���彳Ub��{�9�N�[�'!��/������mP��l=�q��ץE���y��;�p� oD{;�n�sQתc���z~w��Vҗ3��}�+B߷J�y�EX��r.��B��2�``�܌xobr�,.���ۭ�-"���/a�S�b���A�+ʶ�K
t��P���d��+l��.G<�\U�^bϯ�s
,Q�F��-u����3�#bJ\5>�bmIj�Y��x�OxlN^*%.<�uݐ���޹�*K��(�kf��7y�-g�s�H�8:y�\�<�'��J�D���:8mj9�X�L-���̘^�g�@n��M�Mב}}����@�N��G�{�N�s���#�B��\�R�3�7y^E�X]���>0َ�7��M����)��ʆ��̮��|&� z��F�[�����N\v1����t�,��h��÷B��P���q����:��7�����2���H<����Z��
��Y!)���t�8�T�}c�ro��#���;���Y�<��*�X\^��ƣAd8|w�d>��H&�s�HI�|+��s��Ǚsf���{Դ�W��wC+n��Xo�� ���"��3�����ؕ7�\�g�,�9e��`��q�7Ͷ;w;2��<�^\5�(Ӿ�Y��Ò��>{�����k���^oM ًԎ����d�$�o��{Q��z�c�Xk:�Va3��A7�i뻤NE�!��θ\�S{,�u�̕� �v���4Z�%\QT�;[/�>{v�:u�5����iƣ�ɿQ�=J���L"'Yݸ�YgoX͡��3 ��xq�GAO^;�3��1�kf��w������+��1�w��
�Uv�=a,�ܧ^r)`l���V�f�!�a���P͍���O;8dm�Mf�Ӈ�m!)%���Au��U��b�~�v�U�)�Ռ:,�uKEwq&q���1�r���Q�w�}�5zP}��^��V"��5x�&P�������1Ow��CJ��nN�U��0��zw`
�B6���� �)۠Ʀ۵a'�ӱ���Ѣ��0�s�X(q1�qy��$8��e�b�I6�4UȞ�IX4�~h���73�q[6�)����Z֯�ќx�k�5��](j}q.�%�ajN��}�q˶4ƌ���=����o$�l#�u0o6z�UOd`�x�Ǽ���?7F�Bz<����ܿeO{��7�=�q��~��p�;�+=�m2�%�7�,biV�	
e�;E��_rr��$�#���%c��Kt�6�߆�ثa]`�'*��-���oqhCq��)��T�*�7��-�c�y]��d�v��ӵ�N�7Kh\�O�ӌoJ>u�hs����q���U����ˍ�0�0M�=��r�=�z^`ހ��Cʯ^TF���������Yc.�m��j�8��z�u�Ï1�:*��v�Ba�Dhf����E�c��GgR�ᙜ�oI	�%��+}\�5�3�Đ��5��#g�����������Q�%1xT�o�W����<:�wӳ��NwU�q���U�s(.�j�kh6���K*b)�����F�iRE~�V�v�N=X���q���1��+��ϫF�ӎ��nvC:�+����ۃ��	2�e�vM�����>}�G������~�۬�eD���W����N�Ǯ�{�I�A�`��y��7&ަ���MkrhB���"���"Z�׭h�w�F���Y�SM�]�6�Ŭ��"�٭[�:��ޱ��]WĊt�+��O�N�^�;�D�+�ǫ��@��:�vjm_<��h�7��K��g@�y����@�+�$7�|q�3<�N�9�_F��h ���M���;��ɺ��j�xln��ȹ�w����$�I!R����yƉv�3L{���7�(fڜ�*��Ĳ3��vCE��뫌��p5y�&7�E��6"�8�1�i�+p��6��	��wv�`�K�P兇���q��T���j�!����Ν��ƱdT��Y�G�g
z��GV�y��]ٽ�Q����*�U����Yԍd.���s�Q(:�f杂�*���j����rb�4��[���0�|��r����]���l�z��O[��i1;2	)�9b��k#����^�!ܰ-���L���H�0rF=3Q��3s޼;D�,l��]�w����Ϯ	��S�{d�t�tt�l��_k��v�d��I���U�eY�9�VB[��(
�e��1�W�^c��
I$�I$�I$�Ij��4�Ld�d+U�wVbG1���l]Z.f'�RɎ�d�1�Q���]�DN��UW���G/&_��w+Cy�
�@`�$��`�X�P��ba.6Yu �Y�%ƍ�,Z`�AJ�A��V��(�E��FPyI�c^bhFCfԆ�-#�L�*�f��ȝ�d<����b��m�F��˗���+2�V@��U��m<ى�ѡ*��Q�%�Nژ
R��6Q�0*�oɊ�,�RKr�˘��`�w-��1��Ry�8���4��m��@Q�/�]�ѡq]ˏ(;y�9Ң�O��h8-�3�����a��E`%�.�$�љ���Qd��~����n�H�HU���;H�P��AZ�Z4XY�b	baE~����T�gjȪ�01\X�h�P�f�K*,XT%�����������1��CYE=d��k6���XJ (
��&2D1&�:v�l*�%d��H�0����Qd3T̲LIF�c%C�CI�
ʁ�b��+D
��*��Vi�LACMjC��LaPPU"����T���*�*���Z�XC2�r�3�s���	3D_�A���p[3�SgG>�tסM��\;��f�Pm��2�Śy�F�JlX��uz�R�;��!O��ᶰ�P��V��oj� ��Ca��3p7�<�����K���s�u��u�8UsC������.�L���kn��J$N��vc��v���|xF����.�}��y���?{���ٻ5l6��6�k[�Y�f�DLO����L���_Z�)PDunO^���aL|���V���*N�5�wL��D3异iyw<��߬�;��qѴ	����.�o_r'�׎s.՟d<���\W�\�v2�p!<�;���O+���ճ���`�\%</��n�ofL��Q������dC�/�˃T��\��땃���!?�-��ls��g?���*�~�ʺ��������û˔#v��=��7�R����@�o�P�'�	������2���eJ&��sɉo<b�ѱ���I�q~���k��Q�/��X!��ך��S7��8��r��!��;�o/�nk��#�/�ɫC��_G�/�/��YO/x����f��7M��]ǫ�zzȯ��j*�����=��;ꏏ˧p�����I���.�DFտ���KF���1����fM�������{-M�e��b�+�����c��kі�t��;M��2D��s�GA1m����o/��	s*Z����%i���9דVV�yJ\w���m|����E�t��p�'a����뛾��� �(ǻ�=ntc��(Ӥɩ����T<�;����]��;���������B.*a�+���f�1yU[m��C���5�א�BR�{yv*��\�4>���z�n��)6�7��ADd��L��~=]J���6Q:���]Jl�#/�pD�1�*U����u�6f�yw�O�:�iLCg�����I�q�2M0ΰ�~o���z��i��C�O�8���:@=OH|ÈbIēL�����7�zd�`vף�}�\����\ѭ���\�7�6��2M�Z)�D�<e�nW���A�v�3��4#�/������"��pOHv;\���a�^���*�x���R"��U�	T�=��1�uxL9�Dd%p|�l�	�@�XCI��CL�����Hv�l��B�̑I:{���]������
*Vw?C��G�1}�=��=N3�'i8��t�P���a��I� ��!�Y�N�:a�l�����_���I��$=���O���;`zΘ2�~S�� k�!�!�y��f��:������w��{����y�0�@�L�$�<d�JɶO��z����`x�SV�=@y}�!�5���g��J�s~}�I<C���C9~@�d�$�'I'lk��i������
��^�����1�S�&Y���(|$�HghOx��`N2,'����M$�htfd��l�u�'�t��T�>O>������H��'�3�T����N�o�<B���@�N�I��x�k~�Vq �G����~��ןo�N08���aS�,!�ai�!��'��G�C�Ok)�C>�'l=d��`v��J�q
Ϸ�y�w�:��<_d4�{3y'$�hbC<����O������ xȡ��&��2)�'Gӗ��}����;�!ۦ���@�)!�,��=I��& x��)=N�Y!�C]ؠx�g���{��=ϫ����z2���zr�c"�*�]�'&���7�L<�QC9b�b����y:]��/��!ZI,[J����\�c/�t|CQj�h�;Ǹ�����z=�9����=���'��:dѪ@醽�;Bu݆$~P4��^D!�v²J�>�� s���־�Y��������XHq�;BV��3�'�t�i&�oz�!�u����'HOY�Ld��t���7_u�\��_C�������6�����=C~��B�<`t��pd6�2f�$��$��u�� ��~3�{5��s�������`C�i i
{g>OY�YP靰���d��C�C��!����l���w�T��_y���H|rɴ�Rm���`x�wǵ�8�x�����yB�{g��4}`bI���~���u���~�C�c��>��R,�����$�$;MwC�'l�z��!�� z��$�1���>��z޷���}�b��$遶�.Y'L��Ƞ2���|�:����ޞ$��|�z�����u�y���y�~g��C�{d�Ʞ8�h垤�Hv��M����6g�'x�0:}��c�>3Q�S���K�o+]�|�}$�̓�|��� ��T;d������i2)'h��	�<���D�����>��38����yLz�c8ϧ)!�l>Hz�֬�!0��x��<�� o�I<|@����M�z<&=����nL�]�"x]}������:Au��b
�`�0�o����׍�m���<1AlK�2X��;'G�����:u�5'��� �M�}��w�۴8�x�L�!�v��&s���'9a���'���{��hH��S�E$��8�~�߰�����ײi��B�B�L���C�_Y'�є����=`h��Ԟ�*C���C]���ٽ7=�f����]�°���6É�Hi3�]`N��>d�H(z���)�]�=d�P���<dP�9�W��=@�y��VLOv�0��铦Me������$�I�>Hv�F�&0;d�O�}Rx�5�ڏ���]������C�(�u@;d�/�'̚-�������z`bH_��hN�M����6��w]߾ϵ���}�潄:O�쀡Oz���d�l>I�`v�����ܓ�q�� m��x�6����ކI��C���I{?,��Чޅ1�i'��a8��v¤�C�@úi��'�|�=Co��%`y����ɓ}}�nz�9h$�����GVC���Bb���@�P�'�'�YXq��!�|=�� ����7׿w�z��Cd�u`$�w�z�|��"�֩6��	=N��$����N�d<Cl�s�w}l��{��~�{$>��I���t$=I�L9OXC}��7d�`u�I�����rwCԁ�u\}տz�G�9����>�,��������tK�k
�x)��~�,U/�0`w&ǻM�,�u���a1��3	�2I�t	�g�^��"��P�y�~x{�v�w޻�}!�<d?'����̇���+o���L��4��u�N�4rȠ�O�����Լ���/����C�|��OhOY�RN���`嘁�'�N$�tԓ��;g�޻������9���|���Hx�t���Cć��������<zH����;��;Bq��E��v�ě1���<�}}�{�~���1$�6�Ğ03�=`|��q>d�z��!�I�
�zwBx���:�� m<B�zf}��y�o�}߆�6ȲCm=-�큮�� �|������������� VC����'�<a�}�����^u�ϰI����Ձ��<`i�I��5�zI;C{�	<`N��:����1ԃֵ��u�}�[��y��Rq���:C���䞧hC�M�$�BI��X����g����	��� )��-�V�w���}�Ϥ����>��zȰ�!��te��z�x��Ĝd���CHi�:�B�����~�g/~�y�}��3�0>�XH������>B��xȰ��p��}d��)�'L��1$�V�z����y�}��C���hi �I��i"��y� ,����'~xuÿ<�̯jz,����Dm˲���� ��)^0�@���\��n�����ޠ�?L��l�&9h���V�W+��8#���O�uq�K�����瘟���zf#��D�DDY��wC9dO׫a���g�����(��pͷ��
�ڸ��_FSySʃӧX@֝�	���B[���p�K��s����g-��Ɓq��FS��L5��S�pJ�N��[��-V_�Z�y�X7����$��D1z?0���G\WBg�S��	���l�F�se�QN�����wt��w>9Q��	��ܙ��s��fk���z��/���ـ�%��U:�� ��9�;}�ξi���(�ê$}"�N��a�y;F�]t��w&	�	�n�%����y%��?�2�y����ߧy�.�J��}k3��}
�bb��ej��D�O�U-�Bf �)fJf̕����{]�z���M<��κ���bv��#1>9�)7F����uO��9)������gH�ؤ�Q��`���� ����=ͥ�����4�K1B"L��/�֮]y���4U�,��>0s�7�݂�䢖���&��b��˄��z% �ϊ��-3}{��L�75�kM��E��o��+F=ov���ⁱS�5�3�C��g�(hÅ@�xf�������|eB���]�"[���u&u�ѥ�KR��Gz�����\(�O]8��J�?�� _;�3=O�m�WFD�����l�\�ڤ�����Y<sR:O��FϽ�@��H@P"�H	"� RP� 
@�E$PR�R,��"���� ���1UU�A`2$�^���{��݃t�қb���^n�Jo������U�"���!^�97?�?�:��0�it`�(ر�s��?���|j�I�
n����la>'��8L��8%rݥD�M/:(���޾�6�#��hL,̼��RIJ_m����D}��#3+�z/UFBj3Q�J[6���������$�Z���D9��+Q����*i�u���rRQ��l�u������5y����$�i,�!�w�I|�}�7u�j�Cqwr`Z�}ZH��|�u�ܭ�֡�*�{E���`A׋f����n�5S
����N �#����Q������@�.H;<��Z�|3�]�ƩՎX�1�x͸�M�}V�q>y��X)=M"Ȇ�����k���Jv�2���V��r�n��z,��g!{�N�}����]ͬ��McKlͮ��t��s$y��I[Ӳ2Z�AYݕ3�VR6{�e5u7D���F)VO���N#˜�7�J�p���SV�^�N ��T�ޏ�ܹ�z:�iX���13˟�ӹy�J�L�MK��h��YZz�������8[�L�q�KfW ��b��g4��][h���0�Yԃ�7�ɵՙ��a�ɸ� �V��R���c�}�\HS���E̕nd��X�0���>�[[��䄃�2%�y�t�ѩ�Pe_p�
�/����/$��q�2Q��N���e뗃$[����2�J�o�I$�I$�I$�I$m�Ѥ���X6_�xa���g,#F�ʪ�[�W��5X�db�U�>�]��upW�)[��f+l�&�
�%��b)��QF�R9�R�`B����92�n,j�jd9Ba���4���˴�D�C�ʰպ�Q��]�`В���ʪ���ZP�yWW]VK��-ϋA:`�ʪ����N]��*��S����&�e
A,�-M)Q�E:��k�M+v��)��R��"�v�+	��yF����#�0�e�Q��0�����f)ID��XyQ�;#���1*��W�Ċ�ڲ!�er�D$w��Չ󥂔���UUɇUUv�T�,�����,�&]��䢯�]��b7��r��,��� V ��s���~���6ʋ_@(œ�b��Z��PQj)ĕ��i��LP�
��eB�%dTd�LC#c����,Y%jH�32���WV��
��T���C2ְ��tɎ0�����&��,��`cL%aR&��Ib�P��J��Vb9�1����'L�Ղ°�"���@$>������"�=�ڛ!��RȻ�f
���E��[���b��I��_}�Dz�k���_Ǝ�z�h�V��S���~��ʧYr��G��#,y�oz6��mf�W�V��V:{n.��t�$V ӸF3V��x¹Yz���J�=�����E���	�]��\ӛ�ɀ��Yp^z��C9D�êV�!�[���\��4���l�uq	,�[UCS-^�����;�ɖ�F*C��%2�t�V#<0�歫�C0�;����Ca�$�8���z�*�XY�I����f��úp�.tϓ�Y^�u���t��ܵ�]���و���;1���s
��[��*>��[+eL>{Kd�Gۚ���5B^݋��ơ�����9��򳿢=�n�\kbK�<��Yؐ���z(�;�1�=��fv�x =��>���l.��Cy�w&��s��U�^�T��9�����Z8�\���캶v B�8bA�@����'���"o�����e��dL�]d��GPǓ�P,�~սټ���2 >Wحdu���ļ�nذ�D��@���Jд�-I�f����W���HeG�㻡-��V���顡����n̽k�z�����JzxƊa�QO1�����`꜂}�D�Z���ܷC3A�k�e�X���`�j3����3��UC'�LV������6o��ŕ|7�M��D
� T��az7�q��+����'�s�O���流gڟ���2bj@��`�V�a�����;�owHnA~�P:�Ъ�D��Y~��7C�y<�}��Y�t-��&X�O�btl5N���)jb����z6�:�v�3HkOZ�gU{�9b��t���j!O]�>�͋�j��̟=F��ۗs��ݨ1���j,;��{��%T1Lz�ֳq��T��CDk���?-}�v����h�mo}�p�:���v;��7ª�
�Z3,�J���Cp2�����X�Rf��y|�5,�1���ǶT�4y���
;��r���"Q�i�tR|���̖3��C�v�=�0�ʪݲ�j%r"�����v�oR��_{ޏG�/P�Rw�]���N����v�"�ҫh��L�<��ݮ�y�է�w<\s���HN<hV�31��Q�/�r�k���s5��;ʥ�q��О��j;(�4�_#apUOM'���6ώ�{F5��%�=;�ɻ��>�a}�����<҅m������MА,+�W9=�ʆ�����u��ݕ���f^�e�j�<�Dq;H�Υ�)����8\'��Ɲ�$劂,��|I�K��nt�Ǧm��/�����s	���fw7��Si0����b�Z�w�fJl�C��|�]5��'f����S���r�K}��b��Ew)f,�Q�����z=�Z�} �\w�G��^��t��m9�|�a�mVg	�w�u��kbbyG��c���VN��xk\((��9�~��ac؜7e���f�τKQ[��
�Y�Co�]Uo0^�+�e'ę!���a�U��ilW����8g��x�R�k�eA�"�ȹh�ԶK���@=�W�&�f/�sѻ����[u`q�V��W
�|#l�5g����X/��{RS�v!��4�u\���셿i�7��|�C�0�gj�t.^������sݷ�5v"<>�+�.P�jQ^	G�Cb�Lj�EcrJ�ۃ6K��LY�^�<�N8/@� �/c�f:�*R��{���Z�9]�W:�1ܥ���\:�g�s���=p�r�J�!ʹ��7p\OOQ�i���Mׯ�t��o���o����{q��
�63�}f/�]k�S�^�� ����m5Ge=j�9»E�yJ7��a$��h���a룑�[�K+.\׬E�&���כa?\S�������_ PW��dc7GD�Y�c�Jo.�L�0�'i ��}i_]�L�Ꚏ2�U
���5bx�� ���6	��Y��������F���#�^h���[��lU������d������s/#�Wt�ss��*NK`}��hHb
��нY)�;޾QA�o�Gq���?z"=�g�u'�����;�-�3�u��n�D�s�����>O�}⳰j7���@�[
����܅ios}��V�^�L/uue�&'��T1���Bo�DrԂa��ɶeD��1U��x�*�l�Z����N�z���t�25Y��@�.��fb~5\�A!:*�<��2F�\�\5�v.��4VE��t�G ^T�N5��J�y<U�Q�/di�A��3}z &d �_s�m���-`ݙ��$�5���8��2&)��Y����n�7��s��(��`�D^�����]G�^L����;8$�yEy�_�.S��y[��kF٫���5�y:�K�Xؑv3���s�`��[�q�˵�4;�Wvss����8p���꯾�������̛������n�MD�`�sz�|�q�D�Y[鞝lҨ~^p "�����m�=ٷ{��L�3*k!a�i��wT��G2�f��љh���)��ˀ��̓��Yk����R�I�w��K�[u���qP���vu��=F�w2�
�:���[����x��*���
�u�n'6�_Q������R���6��d˝��C]i�ݚ�D��JZ"�����K�Ou.�;�T���w���m����ֺ�v����3ve~l�^�zJ(�DL~�|�Ҕ4����{�
�/�ew�4�.Ry���1PV-c7^�(�V�>{ ^��XN�v����C/NefD�^��MN�o[gU��V�<d���{�0gU��&CGh�j�����$�7�,�|7�/F��mGe-�͸�(+\k����;R�{6���z��X5�jk�V�L�,��q��+��FZ�!��̻�������V3檖v3���������>;��WV@|�:Y�׀��'1�e�f��Z6~'�4��-�t�L�C��ڂ�Uh�o�����L��#i|M;���~�6���E�\���ЮŌu�a�]}|���V�dx	EA"����w�6.Niyjp�cz=�؜�+'�Y�Y?MMD��}�T���͵9�Qa�ɶ�-M����ix��׎ơ���4YgHW�u2�nB�\z�����BL�P�ToQ7���0�
+�y̗����Hg��R�U��F+��i���ăBq�tz���{`G��1���}�����g@>����U��C�7�#��A�-�,KUĖ/]��J���\}kH^C���c٪�ugh͢:�A�!�܄�a�V֦2FuQ�}�ؓ��Sb�SL�f��ǹ�|qQ`������φkJ�go;�E���ʘR�z���gM��7x�"��oveyN��BsE����>:x�i��AC�RuX�����g:���opC��yR=��-��j���k�R٥�,��v��l�v鰑�`9Ae�x-�@��S��^f�fHs#?>���Z�z\�&Sw|͔�-����}�E�f�GX�.B�;HXm� ]=������I�����}��w.����@z*�rU�*�'{@�5;�t!ܭ	mr�v�p�sCFKǭ�3�AW.h��t{E��9M2�W�؉��
6��pwc-��wo�%(�ޅB���5HV:��.E y��1f���0M�u��h����17n6�D�=8ؖwǊ����!�Bs宵�s�p�͛f��@z$�`V��4&�����+0ax�Ft�P[�N�_8��Δv���N��Ֆ��t�v�A䑶�B�A�U��3�
�KU�v��*��`�)��]5���(S���"�%�2.��m�<�"r��fK��vu�*���_��u^oIऒI$�I$�I$�屡��h>�C�Y�2��i�Qe�v+>�]�Xm�>���#�1�# ��C�$"P�K-ª�q6�VDvqU��LI�G-fe�`*�K�p��^��838q\����gq�.쇦�
��)����53Uӥ���9l��iݼ��TP����(�R�UY�2�S-F���3aj�EK2Kj �a�
Y��d532��n��f�Y����m�He�"ܵN8�2*�6f<̔�Ʋ�U�q;uE]�̖�SN���JfB+H��D��Z�R\�^��<B�k�B�{ciV{�Z�*�y%�s���}?T�ovUQ�[p��*�J����f+l&ٌs,��RJ�%B�2VJ�$(�,�������ի��C1!Y�f1Cm��$�CT"�-�,+!��	����T�����*�AeBc&k�]d'��	��Ȳ<����s���N��_�� Hv�|�5%p��SB��w�5.B�_֪���L�?Y7���=����j4�B�aןf�|t�<s-�+�}����׏�x�&a;�Y<�0i���*`>���p�8s`TΤ��#/�"5i�2�s��Ԋ�A5Y6�m�\�9�E��@姚Í���Zh�4�ZƖ�׾�Tn���O�������q+i�,���}��;˚GC�B��r��f����'zcd��랣�l��n�p��Ԗ;7�x��>����7�ٮ����죎��*S0؈ �|�v�V��:D�WPU�1��6��E��v�Ll�Vʴ��T�a�/�K0��s��wr^b��O�Alk�0���9�akӥb����c̞�����Â_`El%woN`�n�l03�W�9�ބ�>��E�����M�nt���(t!G�#����)W���>�+%�3~��V��A�პ�S��.bu�X�9x�Ni���U}�h"��#0xI7:��P�5��{X�Z����qyW��J�[Mה��Y���U������2Յ5���<t=V{�c��Dg�?0�60�.����t�I�����{���<x�c���]�hqb�{/.�];WN�ech>��2`�c�h�k���Dq��&|G�q�+��ݜW�R�}�;�n@�n1f���(=��t��'�.e��x����9�f�kB�ț�Wݏ�ʷ"禑�}��k�f�UJT~�ce��=|����,{�a�)zh���^w=�������d~�B�F�������q�ʵ�R�����;г�A<x`�~2�H��;r���*�_�ue�9HV׉����3��ڽ�6眑�'��8�au_\�<=1�\��A��0���Z�����WI�Q�Xj��:I�)�G�X.���٢!v��XZչ�]��us�;�&�p�s���߆����^�S}��rkq������p��!��lT�H]�O�����*{}�]�sò ���/����+.�ه4����٥y&�Y�o�T,R�j�|��O+/:��Q3�r:ke���r��{����;�G���EC�A�¨�n*�}�rM[2�WO�z$�g[�0�����N�J�wN�=��P���'c����d����Ts�2Zn��z��ءpGv��4}|^}��a�,#g<�u�R�v���W�Khf5�s=��V�#L>�>ZO-"�Z��j�q�4����P�c]]V���So]�԰�ݹzƮF΁2�HM�/�$�)ʸ��<͗�����No��?i�O�V�1Le�GR��Q�C�.��Z�ծ�BKO���A '�xH��ʊu�!W�̈�;��J�2keH���0�ל�XT���6j&}J����<`�t'�<hpX^���Fe�O��C��ٕ��N�N:�D��*�񭐕נ[i��2Bl�h�!q1Cc�GH���/�F�n��AE]����q�K�>$]������c���R�&Ӯ�
`$b`�Qoo�K*ܟ{ETs�91�S�f;�"������'�6|��g�g1�U��ё �Ū��3��s]26�q�&a�u�F�[��K�8��*g�&ј(�J�0sto��Z6vc&g��ׂ��&}�������"jhNL��&�_h.v	��ڰ�Ŝ"������|�kO����@���;9�p���a_Q��#�˱�hLJ5b�<T6���]n��afɇB�S^E0���
@�Y�J�[y}n�����l �9ɱ��s~�{������Ѵ&'M�Lw�=�99!��k�?!)@�������|�i�L���y����ṫ��<ni�==KU;e����Taȫ�T����9�m��ea��zX-�s��˝~�Я�rw���5�]8�<JCN���.:�+S
���7�1�lQ��2Y�H��?.8N�|t�e��z�����>X�����'燢f��㥞����j&UZ��׹�:�<9}�Yx�h�����Qq�����[����W���7�T<�=xQw^P�����3n��qv k�[]�������nqm�:^	c�yH��ɳPf�cڲH��3dY�������>�|g/��2U�Ǣ��me�S�4kۈɗ�q��y	�NWp����'1���8Y����2ϊX�ש���W4�.v^�{Բ!J-_o;��TC��ou6;1�M*YMd�@R�֣g�EV��륷��iW]�'O�{�����A���1����G�o�w��f��7f���7qT ���B�Mް���F�1���^w��BQ~;��������õ֬�RVm�/><t��\|�X&W.�t#�p�\F��4���9��Z�駏��=AP�J��Ykw��{/�NL�W1e�3��%F'�EliF����cٗ��߂5-��>�饔v׎���񓺀�+ݿz��V:�h�}��k���կ��yG�1!>�ܹ����r�v�(�����=hx��eG���#H�g���.�D�^� ���!gkⓋ�,PL����@gL:C3�+�k%Y�r����չ5��r~\h�w�VD}Nj�ܚ��{��utn��It�g�e��L�Mݔ�V(��_QfM�����u�ME�V���C�6�l����m�o�H�ː3(i~V~�H��B��v�I�{���vS�3�	��j��J%�0R�c���(�|����=h�TE�˝׾���(�F�V��/��A�
�.:zJ�0��te���x׫huY���^�KI2����f���>����5T8E���y���&~�Pc�4���@�ҕ�'v>i�Nj�zL�o��<F�p�����N\$i˿RN�gV�j�ܭ�����	R��bqW�Ӄ�7Jˠ���ׯ/�n��0���a`4�6���Xf�i�!�������e��I���ig9�������龞4"e���!�n
6�W�h[�1߉}�:n��}�n8&D�u���q����WO	UC~�y�1�6�.u���Vr�OSl3D��{���[��&�w�iGA��G����Ɏڙ��X�Ȝ��}NHˇT'&�#��xȻ�MұD�<�C��H�ON�s�d����g��'t��J�җ<��K�����	�6�"JzD?z����{���&�Z�^>'�LZNsD6�lշ��W��n���n����P:���'��0���ua�6V�5\����<���fN50�c���z�2P#��Yj�N��Y���~kS8}�o)M67(ܷ�w�Sx�gK��z?G���7v����)��sX�Y��~�lc�<3:�t��!�u�(:2����9s9�n�Ƴs �.���[�[,T+�jvr~=�ԷG0���0,�"^?�;���q�d$�g+ϊ[�N�K���lW��|m42 'w��dH_u�[W�sd���Ӥ̖i1�F�e���iL��~�1�(3RA?UW�n##~˺��uؘ��å��,���`�Zp��q�;�7.	yҏl�;mo���Q\��x���s�!�͜x���j���3�4�3|����ၯ��?r����@����a�2J�*��u�é�A煏,$�P�Cǉ��s��ПP*�� �������Jcu
a���8r[�'����{�xV���{�,�/�ޗ��,�����h�H�����yQ��)\s��2'�1���t�a�������w���=����	�Zz��Z>W�	�CX<��<M�2f�^�s!��mv�I��fĊ�8�U�G�n�#dJ�=�P�uvb�����y�a�uQ�~q!ya�S���ݩ����ɬ��zVt��k�y��x8z��In�+Uخ56��vM!��7٥�q�Q�ː� Sw�[Ͳe2+�!��RMI���?W�W�'�����kǱW��ڷ���_O.6QÕO���벤��x�䌤�{ʇ!�^}אa�Lf��o��Ċ���(WJ�6/%��t�e	)�J�/T�I�0����
ˬ���E�8��y)������{3�x]lz-�p����>��f�Y���ނ�!����7�y����N�emJ�{ne8h�<�B�M��2�꜆�,��o��G]�����]�bBůZ�F�J�X�Ǎֽ>��_B��T�/�9Y7��\+�1c�9|�Akӧ��k]�l�O
��j��=i���g{Xc��0�~+;8�W3����+��+-�ճ~՟5ى��y��?<d���+��X��՗��3 �}!YG����rk����$vq�'m���P=�=֩��S�6�.�<4��b0��d�N^^G�8��h{yu���e���Y��A���͒�g �fAɆr�Ԩ���ǝx�[!l���{Ց/��wcgwa{��A;e��h��*�d�[�+��Co�XɶUâ�H����}����Ud���E��J9�3�$�sp�}R�v�p]p/�A���>�y|��3H�jEX���p�%Ƣ;��˄%��!�42U1�}lҵ��e�)|�IR���������tf&R|�x+��ض��os��wh��]�X(�̈�1\q�f�o9v4iV� �͠��;[�Ǵ����볤\������p��b�`(y���sS�]h�s؈���gmݔ
�oa�c� �=y�wj��w2uȀL�7����\�ВI$�I$��I$��3�ץ U�"�'^�tǢk����#Ϯ����v�b+2�v]��{1Q��ºi�4����Zt+*�s��Jsa4k�����Yp	,q�3#ӓo{L�0�˹�Ӈ�n��9���hM�A]��XYW�b,gK��K3T��8��+5-�d|[U|0'��2ob��H�������c�m�ӗk�nƊp��� �of�$�k���:S鑻gB�Ϫh:��ԯOn�v ���%����]�D�άڡZ�s�m��o�k׫����\�ƅ�r��ݫ㕣2U��D���9ݔ �'�(l����.�R�	k��#�y��ډ���.U,��䘩�;���e0��*L����ٸd�Wk�<��;��y��Py �@
I$Q�$Ͽ�U��շ�<���T1Ƥ�oW4q%�U��*��
�hȨ�Zc4㌩��D�i�DQZ�l�T�D����uk�`,10�a�i*M$Y%CN&[ �VVV��0*DM�6�WYka�c=�wkAHm��PY-�nk!�
eB�QB��T3W�&�T�@;LbɌSL��5�	�L`:���	X+1Qs)Z�̄�bq�LjWl̢�ɻC-���Ɉ�ec��*^7�V�~f�x2���u���9˳Z�!+7���W+^�T�Ҿ��t�{=յ@av���b���_:��D�ܹ���ߪ�g���C�h3G�l����'և�견65���grb�]���pe��UUřsvy���
#�����{wFFh���t�5�c�+;�)�A�����W#5�roy�{s�Y~�O;w"t�Q6�a�df��m�20d�gIs'���|�aĊ=�P�|xæ��/�s%��b܂z�<�r�i�Nn\[�h�y�+���p�v�����F��E(��Nm�0Zà���B ��8��؎����`��o�Ʃ3⍬ybeev;��	��5���7�g+�!��W:�P�s���!��)�a�d邼����w]��?uR�i���yt��d�S��YU�:��$���^P�=K?J��w���j�f�9���ɝ���>=�1^p����?���v;�ɼcv�VN��۸q\�����cjeWӐ��M
s�캨���5��@fm��r���'��tա��]���k�(��1ӝ��ۜGR��g-�Bcһ!b�;~~����a�԰�{PIY�Xv�אS=8���|f�n߫{��r�C��O�a�����XQ�|o�q�/W%�o�뭘�7Jz&73�j���M�K�ڳ6_�+;y�H� b��=όi�P�����7U.lƮ� ��U�Io�Ԋ�w0d̪�&eИPn⧍A����Ɍ�JA��l�og���2���qI�tߐ��V����e8,N��[u�卼��Dd���0W��K#���+=ynw��ّ )��K���.v'M����o�I���H��e�@p��\+���yI��&b�ҭܟwlu�Z�8�$\���9\�ܢ�ʯ���7}���v��%,"��ق���ڣ��iB�̒ª����<=��5�ѯ 1�5���o����<�ϯ��d�Z�W�0��/m��&B������9s�Sn����3\�x.en�����~0vl�.�<|t�E��U��g����4�v��/O����EZ��C�"p��Qݸ��	 '�����1QQ0殶t+f��qJ�d�R��9��L+8�t��Ut��MWO��勉N�I��9��<�B��v,6o/��ݳ�oT8D{�8|r���`�h"5W�׏�ig�_V1�����f講η0q�uN+å"�F�P��0����ώ�t�:e�J^�'��1�]� �������}Z��t���;D�N���eT5�b�6��w(�cGGwy%�OND�/Hohl�4��0�6j2��GX(��G�C���~?��º�zC�9��Ԏ���iV���ͬ�Z[�u�^"/�Z}�|��`�-g�5q$i��~U��J9b���~Xm/�հ��m"Qz�5�������C�粷6���r�qY5EbV���)�O*�{Q������y�P1`">�N=�6��ߏ�j��L�Xo]Ա�׼r�s�CX}����ˠ�?]=�\�?��AדⰧ���uy��U�wg���)��P��d�0�Q����i=<B̺ف,�t���X�8ިo�����<!�[��'�[%�e\�/'�<(��p:�L�O�tF����s�o�OL��Ř��;��J0�"7����y�{���{��Q�n�J�͜�HJ�:�\^�"���{���i�����TB����5[�����M���|L�P|iQ˳����7s�@�c5�#h8���G��h4]E��Z�Z��UEA����k�j�fzs֮�S�zOu���X+ҽ�t����D#��*.��|����ZC.�4�������톙��o�������;\0���4��,w<8o;�u��o��zS^_v[��i���<��@?�մ�G�O^�$�ۯ�|a��ᠵ�r�έ�Õ��sS����)X4��oLr6_+#�J|]x֭���Y4ER�E2�� ϔ�N.��=�6Q�����(&y��������x2-5�W�~��|�3��}r����}�GlQ�E�Y|(K��WB]����*"�A�,I�֡*��N��`1�ă/ˏۣ(���\{�:{�2Y��Z}<vN�(�ؾ����ouyJ��,w	��d�	��T��w��VY�On�bM^:,��{O#Df��f��$��  ���}���O��/�~�����"���Du��&�
���cU���N�w���<�'T<tY�x] ���ָ�:�׌Av�Vo��74d�6�s�6��!＾\��0�b§?�������J�W�>�dC�]���ޝ����}\�7̉2�C�9��_l	��f���3���	ێ��J�'�t��%�S2!�y3F̙2����/ˎ�X_ ,��Ɩ	���Up�ݲ��~��2y���=[s�����j�ign��g=�?��R�򥅟j����fW;^��/��/'�yX���[�H�5��ψ�����o�h!Ռ"=��[�~�r�|6�(�Q�^��H������--_����P�V�h0ۻE��,Λ���3�=w�.�^Z��?Y0N\s5V�R�wChʕ*
Ѵٗk�t���[���2.�����v@����4������/9�G�X�pC�k�{���w��ʳs8�?2q?k�'Pä�M��I~�u��uD���++�ON4-3�W�e�$���a{�^۹~unm;��Փj���)\���N9 ���;���g&M1[1�����s�;;�
�V�D43]�hWּv�<lyQ���+�f��^�:h�w����)�1���"Vk���Dg_���'tIdxR������tz��q��~���^�'�6MO	��3�FX�B��NJ6��'�r�&�f����̼d*cdO�ƼP�K�ι�MC��q���N�-*�J�7{K5Q��ӌYs��	�7��y>ͮ<~u^�y��)���8�f�RD��Ҟ����8;��{i-�X�O�v���-b� PL(��X�&7)�2�<o�k�raSK�/�d��@�I�F�+��'U	����?]x�Uӆ2�T���|�[u'�ˏ�3Duzaㄛ��|��Y.rr΅cM�;�B|wӓ����L_P��L0�8}v�Z/�os�VGL+XG�c����cˏ;|���EEE�F�ޫ���*�<��m��;S�7۲��\�ܥ�v��!�N�Y3��ӆ���E���A-'u��y�W�f�o{��'O�W<>�����jU�G�n�,�D�Z�nܗ���b��9�V��y�a|N*6�����饔j!㵕;y���#@�8x�뢕��Jb4�d�SZ(�R�<j,=�y�l�@Z[��^��^P�p�_��`��鲞X�;��
Rjn�L�旣��ݫ��7���1�%��3ʵ,�=�q�$�ywaԡo�hi2�oI�}��U�D:��=׿��	y=پ:���⥾#�7��?�9�d�0���xf;�fo�n��y�8#6jx�[a�8���V�hq�P���3�����j���Gڙ���z`�c-h7K�,՝.
3[IFx/7��o���]WC(���_���7|���U�}ԶIW���;k��x�/j�[׭Y�h�ݕ�X�l4�g�WRvj���;kOz�q���#�iQu��0���"+��\!4<||{�M���Ӣ�3���Q��=�gH������"��Se�@���|����=4�wˏ#��ßT��j����r�3��xբD�t2��s��^C�ˮo���t�ŭ6��y�6p�@��8�4|F�ewWj���e�~:ndŹ�'46u>[��Ak.� 67v����,�Z�wH�N�C�,��Z�%
�b��Uw��,^��we�±c�#������`-�c��P����=�[a��<F6��90�㆑�	�n�ʼ�(%�#mx����[�*�D��'��0�nB��d��+���}Ȟ�v�`о[����Q�&e�v��o���>��ؼE����
�Ƒg�P%J*�L�Q㸃/x#9R�Xgf6��4i�ԆGy�+VG�*x��w^v{r���}�H�f��ˤ=<��R��53¡)�`mh������#��^���n�4Q�Xj��)i'��D4��^�y��'��gsX�Zp�=9�-,��W>wY��r'��q�J�L�L{�|����� ���#�Y����JB���~�g���}HIl�C5邵�]Q6�D:RE	�^��4�t.Kc���vGUu�5yN�6=�st���;V�\ ��e��;	nh__%�H�*=�M�	���4�Vޚ�9ADm����j�Jr��n]:f���д:s�8b��5#�w�ŮU׏��Y7�[ZVu��t�����p��+m�����*�e�E��^�sTe�r�δcP��2��V�����Y�z6w-�N�m���[iПg4p�
���GRY|����}ɦ�H���b�w��ޫ�b��ut���63k��n����s���ü��	��݄�u�]�\v�ڨ#�����^A'Y��U�ı�f�� ��ݏ��S9^Q�r�N"��r����7iR����nLS�l�����n�,=/>q��V�-T��T��{u��k���Q-�g&�:��Jj�fD�}��T�f�K��0���j�:�a�8<ߘ��yW�&�$�I$�I$�I$�HX�f�y*�/2��@�Ph밪;K5�A�UkŌ��Fk�6��3��n�X,�SMc�.���#$nv:�(��A��]i�md�.�a���%ڐ�f���]���4op4fe>�+݃����}Q+CT6:J\�Q�c-�7eh�yR�Tn�D�+�ft��K�G3n�b֬T�QK:5��n@�,:L����]vT�1�no^���RKh�P�@�Х2-'�G���v/H:��+�aJ����8��\�e��_&�tf��.W�^�h��y���p����]��,:��6W#��˕`/�
>�jЭ���͟j�@*f˺
dKei2��ÛL��`�3�1)�34ږp9�Vf�;�.�9���"r���V�a(P&m��d���=9� �k�ѲØ�L�oO;�Y�x�Z��y]Aͪ�q���J���4��_��B!
�@�d�HĒw��j�%I㊐��*)�b��1�B�q1��m"�PYUf�1��6�r�T��hdt43w�-��Qꄮ5��eJ�آؓe(���ݕ��V��P����Vb��%Kh�����ADf8�f�hz��҈bHs�!��*��l��f����B�,ef5X
��b`�#R\�����ي�T�L������_��tnn�<а�����6M�3�V�V�J�0	L����������fg����}>3�5�wat.��1s�8h>ˍ�c`�ʖ3�?��W��R��j+5)�����4X�:�t�OsNUZ�Kʹ�Qڧ��Z��X~f���ώ��Q:+P�룚�a�#Lhc�A�k$'��yx����^l ���֖|l�����R�/�r\���������x��)D�ӈ��̿&;�8��`:J��Hi8mU;��]m�[x��f�|q�[_1S�MZgH>W�`:IX��ϟx��a��bׇ�e+���|�̧�Q~���L�i�޿s��D8�gOj"R�!���Bώ�:<rٻxv�]�ٞ�P�=k��C����H� �9�D��6{ӕY�X�QXO�+v����f�n>���7~��+4�3��r��t^_P=4�xj��5ED��7:;9��x���1AK�8.װ��'?�}���Y�gY��K���-%̔D>]�V�9���ۺٯ�9�ޱp����}s:)�@�b��NP���ÇNrDQ�g]�f���G��E��K��`�æS�T1��x�u��m�c��}����d<Y�͛�?����t��{���du/]���9��XQ�+�r�y�ܔ���d%z�Y�*R榲��zo�^�^ �qةӕ�[/۲*:|r-�_�t��1i�P���M�l���kޫ�.�ńv!-qx��(�ђͩF*e����k�I�����g��|h�b��H�7�<Qg8V�r��}ܝ{��!_]�5��2��w�š�|B&�*�}rz����/�_��F��%΀��#�{r����@b��X��:
�[/.�2rءgY��-�ۜ�Д���)�
e�U�78uvkT��2�`�[��tZ��{l�D�֫�����Ouǻ��}��tG���IW����'��ccp��F���W>�����H��w�u~�{�8<x��D��G����40�凢e���C���W���=��|��H�Ƈ"q��x���H�=m!W�ޓ����*&a��K��l�Y a-�<�=xQ�^A�{�X�޿mSUh4��9x�XK�Υ�e)��w{M�^�K�9]k��D{U��cL>"���֣hqW�%�S���RW�BGy�y1΄���x^�)#��~.��Y����ZdZk��μ�ő�b��빁�U�93P,4\l<D����$Ѯ������Wܷ��t!g֬�ƋJ��e��3<�)Q�+��U�>�z@�ͧFNc��0�Xl�j� }���~1�]Z����mp�!\1������kx��X�T���ꪱ"nNY���[{�,��{G>�=4��Ǎje���gI���6�5����GVR�%��P~u��?��.�i�;%�'��x�>��Ҵ��~z���o�x�������l�QW����E5GNG���]�hx��)�hWV���]
�b�(i|���-�>m�=����?ra��ur�;�7���t�(�Kc \y��=����;Y���N����UC ?)�O���'�����Xо�M������,�e��útԦȧ��ć��]A}�=!gE
R��n>Z�2d���S��NLb��Fz�	ha�u19B�ima�����u�ﲟ���4t�FtR	�ិ��mp�p��.z�ý��]r,�xr$�6�[Y�7��M��8V�ͼt��ӆ�L�}�]t��Q
��0�`�185����GTS�r̷�E+	H�u~���N�;��b�mߞu�n-׫��dc�\�Fo�+7�L$���=�}Zp�l�s�Ct�<���^^�Ъ��sË&g#ML�q��e�u�E92�g]C��ד�UT��A����!#����O8d�gǏo����.����U^�oi�!���f4�?$��.Ȩ|v���b�l�Q��%rkϕ�H#�[ӏ(�X~G�(%t�Г����h=G�j�������:�k܅ֲ{�f`�2׎έ>z��;�m-<��-��l#�iƆj㬑�4jyߚNgoi6<`���4S��I��5)V���˘1<M��� ���N�^"���܁�8�.a��|����ʖNlm��]hX����x>{Qɺ��Y-�!��hD1�n(���WZ;��s��5��x���)�d�j꾌�}�WF���	���{���:MF?Z�q�Ɲz}���p���a�����͋���ު������ǧ�"�����̦(�2���Ī���o�d�ER��hdϔ�q"X�>uԦ2Ek���g�t�7�V;�G��C�Bj��ٟ-03eϢ��%�Htb�!�jtMb�:��8C�#�چ�9�R��n�g~�~m�+�{H����Z���ա�gAG�Ԭ�f�AU�=�i���xQg�}�;��<FLd�-;<��y�"�l�S��T�y��xt���F3#f	lݬ��<6��̫�y{��_C�o�Eb}L>o�xa�XQ�<��@�QȪX�o�9����s{P����N�f �&������+�_ǆ�C��YS �^Nʑ��|yF���>��L��S���Áa�0(k03��/�X�r�I����p��y� ��1jg���f�J�G�N�;��˖�e�3�W
K��{ڰ��ޝ0�/Z���TY���#�kn�'o
�,����w����珈���i���yn�fr �]���W��@���c�<ni�_!hW�^�beNĩRu���Q���J�r%ϝ��DB�\�[~�Z>N��l�ߪ�on�.l���e�9��*jc_Z���H�Sۀ�~�F���;�NOp��yH.>r%���'�?8������>I�v	�*e>���f&�S2KbS,�0K狓��tg���T���C^�V�'�N�`�C]�o�!��j��s��ϲ��yi�^zL
x�Yώx�NJ�4�͝�5��wpf��<|~���c����%�X��^��.�}���wN8�زVn�a�\iY:�1t�{|E�����G

zf��}˾��dMP��0�qk�C��Z#�]�H��l2�Ӻ���@���Wj�n;e(�Xh��xɼ���/$�}�`{�z��Yk��q�]�a��!�����L���jk��מg��[֧��ش�|u�u܅�����u��oeC��1m����O?;�M/�\zq���;V6��X�g*L��Aى��\��72݋S�>�V&Q�&{)�E�j��iƀ?<d�c��p�D��Ѻ���43˅ݠ��ƽF�;�u$(�,ha���4�j���/����EkN�M芈j(q�4�ա!�\z�C�~4:������oi)��ဣچ����p>:hrv1O��̤��Tw�fȀ���:��7�JT��%`k��Y�2�Uot��8��q�7$�gJ�/uj��N�Z\]��A�;�#e�ִ���S�|`�/�}��]�k�;ݛ�����g1|��;���;��n��mκ��z*�����'+�^eE�="������l��Cϟ�⏊2"t�{Z/��"�i��pa|E��=/"_���q�x<�f�ӳ�����e0��D/,=K����w���yn���A�����m[�[��U�f�F�ͧ|�����ݕkyҠ�L��`Q��<pᆎ�=#t�>�dkeQ49��ݨ��Ȟ3�C㜬�.:s���8�3�v���ڑ�!��'��!���ߙ]T+>�ot�و8��[��l��f4	?i^w�Z�YW4�{����erm�W�T����Jy����ʖځ6d�]=r�8ڞg}]���{O�߯6�m�$��1)�"�{W�%:9՛�޽�\�ΜL���t(�^���}�3���9�r��G0Ͱw��� ���\sǝ�Z��A~�]V�ڻ��̝�3F�����`��n�4l騰�;��be#N43P�k$d����Үw������Xh���髋��JT�4�����8�l&�)^�z�ne֑����. �C���O�a6�縑C�v�� �	�cKs������^�|����1K�W^�BLO��ӧ�ֻ<vSi}~Z^S�Rـ�DoO(��Eּ���.mE	&��f�5�o�7.
/X�.�C*�O+tt���������u�:�Ņ�q�;F�ԓgOH���z�c#]�ﱼ�x�w�\#e�8����iG�\�˟m�S���S�0��;,ӑ��}_p���@VnL��S��L�S���l��f벐��ә��^7j݋�(:�*�E���i]u�?nf�,����!�����;|2��^;o/�R��x��ۮp�i"�*�ݭ��kt]�G<����-�IU�u��]�|�+��S$��[��pu���a�Nv�B�={�VTG�Ke���fڐ.ΐ�K9:'Zz��8wU֯�F�Suʬo/���;LL�C)��[��7^��W.��hs�ۏ�nb;;	��O.��Yn�XY�ɸ(; ı���lvW+-c[�X�6���7��0�Pq�Wz/�gb6�X��yIK.�x�
���5��}}	��
�rx�Z��X헲[���ٹ�mIDZǔ.V� [��`��k�`ǜ�l��o/���-������U֜7�`������2��x�F�rI$�I$�I$�H�Vs�eR�pR�j�IaKQ.&~ P�*��HțY�WyG�5���	;'	B�SA�D�b�V^J��3h��Fj�vAD[�������jܔSO-�"�%	��,M��L��
ZITtbti�%�j�t-+�!n_\�I�!Xk�GQv��~×J�I�"T�V�c��~D=}�Ok,����R7*E���NZg"#k:�n�>���$b�ԉ� �[&5E�`e�J�1ēTl8d��(�Ц_+��mڋ(�ur
���<�Z��m��Ẵ��AIEsd�&2]��*�]U;�l�DR�����v��U6n`31��#t]^Q��xe���$�f�2�UA@�VV`�wU�$3%�2T��������۫VhŻ��IAhK�i�EAU`t�
Eu��LZ���TĭV,=a��E��.Ywf*��DQQDf0R�Qexр�����
/��
�P���3$EX��U�i2����0mP��h��fi.%�X��/-�,�j1-�5�1*+(Vn؊[*"���n\��TV%@�DX����U��P4�
����**(�֪$PZ��ˆR��,�PEgW����\�j����S�H���6-��rR]4�C7^j!�c�8$���z��U.4/c��ݮ�kph�A+�:�Q�X��J��8F Ae����1e�W ?Z�Q0��Vt��cOjiv�-���p^,#=��21�f2�`����7=<*���\�;TҐ�t�Iv&oK8~�L]HjV}���B�	aa�Q��e)������YK�.0^O�7G�p���ǔ���Aچ��2������|zvaäX�ańP�{o׾�8�m���_y	J�t�8����v����M�O���!���]���\�����~_Y�i�����6|V=�kgL��#�_3v��=B�]_+��K�>��ٸHjDuɵ/��k�8�m�ӏ6�kjأ�m&�Kt�K޿y�8|-y�=�#��:h����f�L�{��w�+�P^z߻�o/Mlaj%V�<b�m��7���������"F���;Cj�0�ʱ?�2�ǎ�z�0W�k�*�0FU�:����1N߈�j/�8j.7�7R+P����f�y�W��|ge
9i�0�`NZn��ҏR��>"����]��*9`�:�5��fj���N}Ƨ��n򉜽��H�_O:rο�G�C^�B��zk��Z
�>/N���>�-���Q&1�͕(ưل
ܒ�uw{"d��纫����[��(r�P{�ԅ�R��Ә�5�Gs�7R��r,\R�{F[K��]z��{�j+I^<s��wF�<�����-�����G���ΔvU�߹}���C�`>"/��2��K��z�~@���t��V�Y�/b��MO��/�hZ�6��(��{�!��^v3��*����a��`�ڹ�Y+��f���}}5��nJ,�0k�Jci��Y��Ѡ�[̾S�Uȑ*T���D~��;u����vy�&
�g�OhD�ST<<�˪1ŎoL:C4l�ώ�\ge3�AY���Bshib�줆�4�ʃ6�ww)J�����r$c��z��8|hx�]���4�m��u8���qc+j�޽�q��tg�'�e��S73pb�'��8yzڙ.�;燩e[�s�H�=�B��/�}m�h�
�M� �7y�2z�D�U-m��N�I��ܸ}P'��m�O[�ed��16��.H&.>��y �"��e5E�)������j����\|��Ű��~�:��!��5����.���g�������Q�K����f�ǖ�0��4|�����eㆽer��P[\��Z0�mCr,Q�^�6�.�Wk����lV�i�srFjii����|c�����^[�]�Lw�sV�2u�1���Q��9��~��1��]��g�*WC�v��/�Huo��ٜ���+��%�����N\${�Lէ��*��Y�OM��\_�?��gK�t����6u1�ຜ}�`��Ҝ��q��`Փ�2�ޘr�Ɂa�R�����Rf��-��j`{�YF��;��D��xD̏gMΑ��U٫�����ʌrXa��-3oY#L
�1�a#�_q�����}���A��>#M��.<fs�\z�Q�֛��އ_�
�v;��W�g��l.:Z�!�ly��}���x�#I�c��"�ɝ>R�4�GH>^�`�/�����*}���C�|`Z��Ȫ� ��̧�a)*��\���!l/^<w�ٍ�g��\��i��z�:��K�ⓔ�xyI6sO�ӕ���Mp�ʮE��ܝOA|��[�l]��D3����0�u�~��=�:�~�J#����7�*�D0�>�;��7�������n�L�:�Xj�ʓ7!Q���E� +�oz�We�;CK�lD��.#-i/"�r�;P���������=���}�O�˨�&�>�!v�lZ�R��)N#��6���I¸�Nrcf��,^0<E��M;�Εށ�N]�qz<��Pv�:p�Cyq�V�"�����8v-kE�=��3s���j4��U� �1�*���g��KB'��:��n,=c3� ��/(�s��Y3!ю)�y$.����I��b\�+}N����}|��h{C]�9�'�ƈ�u�a���-x�����\o�n�q۸����x_a��{��aXu�X�������#1�8��oV݊=Ԏ�j��ZV�s���UIs�t9p��bc5�3;�Ty4t�n���K�ݽ��,��c�'��h�5u�?�W4����=#Gv?7���[�x�4;�>?kUk�j����u�����n;ۈ�7tD�ꎃFT���"j`���:���[��M�G=�ftFa�O�q�%ȑ�q��[�i^��gM��oo#��ӆR;�y�y�#L�2�9�'�i��$�d�Ӫ��ts�����3�U>3��>H�5�in�b�2�6��7vx�d߀ᱱ#�:�����FrD�w��x���i2g|v�I���<#G-(ĥ!�Դ�>(5�=uoy6�c���t�2�ׇ�f-5�"j}��l�j�h�c���ة����K|r/���H�{(��X��0y�������Fw,GFMͨ|:�����-[��5&mE~�����aΘ����2V��u��n���f֞mM]*���IR��2xk�Pu�N�>N�@����w��z�I��kin�T�b�2X��M�1�|x�Z}�[���4�G��tg��/z�f����+,�V��y���<��Fٚ�R��"�����Q���=ˁ�TYS��|�Kt��+G9���2���b\e\�V�LE��S�83+4m���hس�Gї�h{�^�H�ܵ�����A�6pÃ�ۥ����I����QX�u@� UUGBs���ZOO�"6nXk��������:�щ�.�!�>۫��tў�Y��o�`��p�Fbd��[^,��	
�7����Z��&p��v!�
�6F�zF�~[�}�����kһ9+8ã�i�����ﲾHվك�ף{�r�sjJF�
�M�wzM%�x|�om2�3
uJg
т޸d��|�I��&���^��חX����?��,{�a�)zhʌz���:zޗ��6�x!10Qw?2���}q6UE�#�F{33s����ׯ��3P�A�/S�պ�d�MWi���/�����+x}�!e�����C�Mg���:��W-R�`	3=r�\��g�U2'�\^Ҕ�I4��,a�ђ��.��**�/&���!/ՔHӥ��Ԁ��������3;�S(�9�vd��<lޫ6i��X�wƧ6z�Ay��*g����vt�:_.W�(a�X���M�?Q�;���M�ӧ'=�L��ؙ�Gj}6�˸�� ���� IM��\�Xm{���珋�pƴ�(��0�QPw�gžbffb�G�o�<f!~�%uyK��j�]ݟC�(��OKR߭9RM�i�|9;�9VG2ĭ�$6�2A	��"*hO�������o!�J���$~�zo�|�h��K�V�Q�.Z�/�5d�w�C*�Q�U�v��RVG��W��M#m}	��C��^����*&֑A!Ņ{��:c�������Lo<l�L�CK&'i�)�u3P�ic�Û͛Շ�YJ������/�廕��y��#m}�@�{�?q�\��U�"��ƞatNu�M���G�c��=��|B9��?l{t��i�&��Ӕ�K�� ��⹌���H�3Ա'a��'�X�n���O�H��n��v.8`�[{���e�8�)�.L�ٹ�3��r�\�M
Zvn�X۫�/��.����!V�c�Nhq�9i�����{�'��x ����B9�;�f���G
�mѳH>��� }�+%d!�%Ș����Ӛrp���\�p��k�^̓��\�s�n�L�P�c���f��!Z�nA��^�{&�z�q ��.\�WX5��b^ ��NO�\��f�w:b����)�2�d�h<^;m�������"��eŤz��2�O���X;<�L��ȑ�c�ً긳p�������L��ir-�l��I�kb�TX;¾O�L5��+ޔ0��*��>�s��T�:����E���V�~��ߘs�̧WBS�Ti�L>Gt��TE9B�f]�ȣW$)�R�Z�[�:�N�S��&7z��0�P5;ŕ�5N�9�-��I�{p��Oe� �f~;F��K:��4ťK�kU��jY����5�n��;nӾ��k��{,7�;�,��l��i�ff�m����c4�WXj�8崖��]�Ul���,&޸ۛP����z�)o<\�s#Q#�|/y�mU�*��{FL�*ԡ��â����X%�h|3ge\��L��W��X+"���j�#�;��\4lo$�gQM�۽����!eK|�ַzsqն�!,@�L�ݒ��e�͎��DoUv*�ڛ�~�J�NF������v�֫RP|1b�bG�U�aF��^���:w��Ӂ�jk�{�V����US���2�W��v}����\�>��⣼iV'(���Xu\I��Ǻ�c�F�\��/tڐ��vH5ٚ\�����b˒�f���:�#��9���a�̝�)������Ꚛ��n$�I$�I$�I$�g�r����j���Y��T�;�+8C2���O.E,�br�B�2�A6~T��qP����9mS1F,��3>��wwD�LE���Е0����\�cEQ-��z�X$j��rҰM}JT�a�9Ye�X�aR���@Km�Y�����7u���N$���`�1�fEC+'�H"`w� ��]%g��g$��U�uTRv���mJ$���Z&ٷuT�p�JjLh��4��DmtTy��W�-EWR�Zf�B�$J���̺��$�03lQ�l�upG����͊v.�f%BP��Z.���Q`���7�x%
Y���l5I҅�2U夛*է�ղ�%N�;�E��Ze�`��ݸ��UUe5L�YI�㰩������VfA	 ��D�bb�+jZ���EQX)iEUFe�V�]4P�X�����L�V ��4Ī$Qb�ir�(�Eq,�*�TEf��mh�%)m)YVѭ�J��*-kS+E2�Lm��eE�̈��uM0ƥ�s,��n�`��j �QETm+-
 ����ul�TQ�e�X1�A�"���\a\D����i����j�k������\���8�.8�R�1�T�DX��QU��ڕ��չU�U`�+��e�(��s
�P���8���k1����.��ŋR�[R�#V,rԝ!��,TR,���s�����[����rZn�&5Kzq͒�H�sSœ�S��
��]�h���z����G�w���v��ޔ���֝�����V��j��)ki���ڼ��.+8f�9o��tx���f0��ν\� 	�юoE��i�Xj�z0�NB#��.H&]�ɸx�v&���NF�:� �Tw�sg.y��;ù �[)BG�+)n|s-��V��g�ɛ�7������B*�E訓y4�K�A�$�ncLԜh�+Nk�Q�{&�ZS��9X��-�I��=����fx���\�4[nہ��hPe#��R�_2ra��t��-�wu6����n��� K���d�2���͙�����H_�67�3�V���ý�,݌�YGr��n�����+�ej���^�Aw���0h8��d���j˅�����Y�}L����Q�B���֑��{
�Q,q�ν�`NE�#�����Ŭ��^T��0�@�f��쌘ї�ee������n&y�9�<��f�Z���OX}�>��w<ZzO�1W�:�\_7�Tb׆�E��ɕ�x��Q0�^��
�c����&�r�Y6������y� �u�}����ѾJ]���x���Y1��HXڍ�W�d�6.N���y�TawU*�1������ig�iAj����$sk�A�Ll|��ho.�u�5�m�֤R(���|��2N�Q�ɰ�����Y�Ҙ�@��$�ێ�����ƫ�f�E.��=d�"�F���:T�	�b_��b,;�9�r�^����泺�}��	{��x:��{�o�2&|Y��iwL^¹m���U�g8��PюnP���ZoRM�\�@��ܓule�6󛞬�-�}�Bq�i�2R,�����𙻡J�X��D5���H�`����P�Z�ت}��l����?2�+O*���9G�9cn��݂Vj���'-9����ۥó�K��EFGq3g��m���ӤΧ�l�d,̤�(�,��O�5���gї���wDtY�h��n�2�-�M	\�!��6?:!����gkj��2ս�9]A�؀�6nv,˾A7Ucp�noY�6�^���Y晏n��%�H�s�s	gշ3�T��u�4p�/�N�_�>��m�sd2�^�0��0-#br|g�Ӫ���;z���|Ê-n,G��;b�KUŐ�D���L��d������k�[�	Xe��e�ש�-����-� ��`߳�\v�.����N��{U��;�9�f-��� Ŧf��l��~H���a��N+k�N�˕ܠ����E��Y%T�C�&�Nݓ��y�mV45k�jH�rj'�]���2Q�)�/�]�v7�u�rs�v��y�]4SBg�)j.�
ݡx��'��E���f2!o9��^1OY�h��D8[����`V.�"f�楚�^��n|\7���f�UN����5B�-fs�\�X(\zjNb������)�z�VVp̈́r�]���9�<����-1����V�sf8��5S��"0)��#.'�KxZ
���BzooV���
��ܚ���>J 治%�]�S"�^�M35Xo�#��q�a�v�b\�x��T��sRE���-��rS祭��"�_B��_��c��M�����	E�3${'@��BQ���������W���3U�Qc*��p��ЮV͒!�V
Ŷ�*]��u+u�/f{���n?Fe�t��)��ŝS��`;��Y���C48�W`��R����U�f�"&s$�uǊu�v��*���^5��#꫆k��^�w��Gc�!����~�Q���n
Z�xGe���]�7�k�㝛qu�h��uj���W����y ��$�3�y�6V�b7'�o�zH��ٍ�^z��fѺ�`O��U�o:7s�|F��M.z��\:��c���.T<���`�~�����o��1.AS
n�!y�R�6�9vC�v]r�K��Ǒ|{%y[�߄��Y�4G-Vxׁ�Ǯ\�巑�cJ5�9Vo=�������%�^mŽ#f��8���E���7�W	�{��-Z�Gy�������g��������i��!�����jy���GK;K��bf��:�9)��9�&�yj&�Ag��22:-��������wc׮b�U �1g�VaM&[w�n/X�%�Z�f6�6�k�#��9�R�Sa�����B�:�슙����fg&:_k��^�x]�h�א��}���o��d����>�V7%�{9V�m6�)�~-v�5�Ij�+�i�~�S��5Ppt�!��˻�6�����겄�
#Y4���[$�J���ݚMd���Vd̨d�F����]�s�o8bU}`��']s�N��'"�O�ݨ�Ռ�ż_$,� �Ϻa� Ac����5.Ƈ`w$g72��1��j8%�(�#$�N��䐛዆�k����3�,��n����M>��|Nv��p�A4*ìk���]m%���>�N]��2nf/��y�F�c��������M,�r��[�q,��7����E��^U4��;�7��wj�T�=3P*����*lo����=Y<���]�C-t�`Sg�K(�
IP��g��b:x��^�g0_<��R�6�Q���&{v�n�%.�V�S#=wȫųȌ7�h�痀&�{�\|�g4OM'�q���I���IY�gUќ���<�`�]OL��M��jדԕoKEbe��n�{ -1Z �*7�Ȉ,�t�xy\��j�_�'���S���a`���=`��mȺ�
ql~��������-��2��@��z�x/�h�P�u�N�q��575��l��[���uK�qs�䚽��{);8x1�D����C�<��y?}�1��n[Cwe٪�12Z��d�b}�p��a�jRڹD���M�j�+���#����e�*}�*���ؚn:"雾xԐO��������g�ئ�p!]q�����#w
|��t�^��0N�4� a%��34&�ʹ�`�Ϟ�`�Y[�{ �;���P�º����'!�(��벷�"�M�f�v�do�W��uT�2�<�xbՔ�/v��W��'I��7�B6�DwίF$��ʧ�k���{��j���0���O/ja��ua��6]6�]<S�9Џ{x�ّ|�W~�={���P�x�Z$�1㊪��sW�XȞn����B*y�j���'���)�;���
?�w�K�*S�ź��:�kr�/�� �Vٚm�|ͩD���1!0c���*��O�Y�[Ѫ�Ǵo�a͎�Ƥs��b"^�;�v2�!2�v��U�tC\�P[֌��=�yD���n�����iKɻ�h� l�G�2���m�m.�ߴa�8�P�F�)mSC��� ��u;�ӝ�o��a�l;��i�(�@\lWZ�ʛ�گt��Y%��2`o��>	��ђڳWҼVJ�gy�GED�x�&�T��Y�xtn�;��d@�kc�a�O��*�Yn�p��]ݪ"A������C�5�T38%w��qzo�]#���h`�Fm �i��sZ�\=����'/�)K&Wvv�����ElCw�.�,��^�˷zCC��՜:%�ð_"a|7f�s�i��o���9��*��y�Oo)���!#�]�6�����*���������rI$�I$�I$���������)_p����*���7�m����%�E!�������)2����i���q]��V-�1��Fs�^gȜ�n�Z�r;$�a���U�!d�B`�-�&`�	w0��	�Ta�ٲ̥x�U�WN��%<BX�s)e ���ww�b�7y�l�^R8�$"ą�p�uH�J�-�ʹ2CT);r�Z�>b�@e�K��:�⪠�J��7p�,�s#Y%�����0+��"�JrP��T�60;�Z�*T���չC\��fY�ssVq ��:���QbB��e-
�m��2��C��[`e�I�s���G����c��r�S,������Ur�Q�Q\��UC�b������Ab�T��R����v�&��(��0�j��b�1VZk�(���)J��Wv��Y�,Qb$Qb+*�SxPjX���G�+��E�VcZ�YQ+m,�)ZF�*
2�*��m�Lj�-r�DD�c�LPC��"�Stӎ��A�-*R"���,�U��塅���DV�[J��r�b��h(�J��l�y��J�
D�)�dZ�#�Ī�EUX(��Q�_κ�W�^������k��ri$�a#]_Y�b�	[4BF�:Tw��e��`4��t_["6�U.�B͆�*r6���4�r�����������G�/�oz�b(zb�R���:B�+�n"�z{'�M�0���}bA�Ij/r�`��6��s|^��no?x�,�@�y(�G#cH�u8"�0ז� �0��VjÖ���a�,-Q�����7�G^�,/nw�'�j���K�g+f�3��o�Wf�t�
W�p]$1i��h���}��w�ǁC�M��!��r~w]�F]��x�"���Lj�S�q����U����8���n3���� _Q��lK�(�`�[�E-�M��r�Eb1h7h�ך.	˗�;��1{t�r����yu:�jWp��
��-�+j��;A�9��k3��S���wTq�z��f�ui�9�Ȭ�nЂ ��hl6]�5��3�/��Eҭ:�N�(B(�ʺ�Iӊ��g*�G@ۮѬ�����r���/�Z��cj�خI,a��_x�����'GK���RVi��<[��Y��%B������#��_&̍=�T]�B.�����.�<��i�Ѣ��������<����;ׄ1�lh%M������Ț�;���CqxלT��Յ�5.w ���5�F���]�qU�[�=uW'k^܊�.��`��v}���&�!O{z�cW��u��8�`�^��r�{������cz���[ܮ�U_pĪ�{K��oa�d��M�2��iù�nD0�D�9kWs4d�h6����F���#=\���e�}n����|o���`�s�z���mk\����Y\�a�̈�v@�p����A�[t�An	R������7�.-mA±��Z�D��'b��uÖ1ŉ�g�U����B���	o}���ڵٯ�^��c�8\�Rt�[��sv�̏V��tĳ��`6�u�@9d�Ib��4h�Ç7Ӗ�P��f��ʤ���JQ�
���=��=��#��j�m�.)�2!dI��hڭh�@���|!���Z�'FS;�/1�����闔���L�y�xQY�dtq�ӽ�C��DS}�n��� }��9@��Z�r�KfsN��7�az��9͘ٺ��Q'o-��#N6�a�&	�Үa��*nl��krE�X�*�?#Q�K#zVå���$����ɡU�w2�n)+�j�B�q�x4�ڥ�d��G7����:���|�g40�i,��	�J2@�yR���B�8��Ob�y\�
�6�b�ݹ�QX���N�j'xN�5��ˮX��f�����ju��`����r�"=��]�������#�U��`C<�H��5�5=y\�gWz�kèM���6��^�9\�9��[�dA7��0&�E�(�<y������n�W� ɩ�f��SU��jk\���S���٫}L�j릲�毯 �T�`A����さ��	)�3^�G�"�T����8tҼ��$�/N�s���}��Ց5�k�@0L�d���������m��"t��v�1�F4��x�a.��f��et^�b�,��vT��e_�a�F5�m�q!�ʈL��ܒ�L�D���M��)���ɥ��uIf����M/�U{�[{nc=S4(��
.V�p�֋]j�&���/o��IB;�a>�j�i�ю5��#yj�ѝ��S�������J�*�B7����gp���L��>)��4쇇^k�d�C(��!ba�w���4�D�ݧ1��x� 	p�_��:h�*CS̮n�B��-���Cp,����ņ���Q�Ŵ�Y80�׻S����]:�F�M�n�֬
����'}���y�2�թӚ�guX9&���U�(������)�\|,���{K~�_���Gζ��E��fTݰ���j��gD*��d5QI�&W�S��ѭ*�<�A���J���\���D�oK|e��r3r��?z
�^M��;�$���<켴9�jV$ͬ�Sy�4��b��M���)W���F?f�6�q��v��\��\x��,�yۘ�gw��rW�Λ�zD�Yt1����ϝr�aYA�J�ݜ㎂7x0��M�4��rop,m�޵q�aV���@_]r�E��J�? R�)o����	�^� ��=t��Q��!�'MH��'sط.�#�U���?`�
���<���X���ѷ�ժf-'��}���
�n��(_�V�di���������;e'ټAW}'���9/3f���c�z@Z�(�h�c�t�f���}Y�&�цZ�q�UD�e]Y1x��AuL�>R��\��A���[��84+�ؼ����4K�3�n�ZW�-Ka:7�wK{��c2�,��k�T�9�r�@,��v�(�{b��yw�؄�h�]��%�`���d�����پ��ѐ�cVf��4��W�K:G�;�g�Wb�bj���G�{��cO��~0�͜�������]o�K8�ҳ�"���ę���xf.���/=�[R�zz�.^�-R�+Fa�������5g1l�ka��-%���ڂ�8��l��0ŀut2���S�M�$F����>|ྚ\Ҳ��ଟ�ḉ��{��+��}b8��8��q��W�
�>��w7\$�r~�u�N����L,[_�����V��H$\�}1Vs��L�ֹ3�I��`��f��`���V�0���[������6�����E�ޥY��t�Aᛃ�},W�8[n8�z<��"���r��S�Y�]2vf�q|R%�Ѹ]%3p�@�̪�,�NDe�X.�.̯0@:^]��=}�ؕ����y�t�rj.P
P4���s�
���'wM<���>��#��֘��l��X�K�r���[&8�>��n^b<s����M���cy�91n�8k/Ln\��>���ֿv��W�S��J8t�w*N#�&�c�]��P��#� �'��i�버Jy���Ux$ۼ�rv��>�w'4N>�$L۱&���u�#��KsRq�o.��@�Y'o���/+]bt4±Í�o<&��Ek"r��#y*��f�}��d��%�L��M�6��=C|Z@�FIag^�
�Z�|M�}c�3%b�%uq�trV��zV
���4HRyg�Q��y�έ��1�I�?^�����6on�vlthm�?PW]i���ksTc_�N�GÕ��f��m�(������W3��Wn��@������n���
�B�2���Q$u`œ���a'�O��}�th���<e^ٮ�j�Y��WT�.�p��e<'�+��Y�*���Z���DB�&��J��3^��1n��s�l}�l9�l��+Z���۟1 �\�.���-�& �{�cha�?�8c���U�
�
iI(��U"o�˜UX�y�N�X�/VT{��8q�]��b�R��G��Yxmd��#Z�R�F��:�v����<EI���ok	�$��uc	;Kᥧy����]���-�t�
	����ťj�ٛ[�gf�N�x$a��1<f��]Ѫ��ᙖ�Vs(.���bKof�j�t�Y�v��6���zM]_e}D��j�LRB�I$�I$�I$����A���<�z�ո�.��F�C:	:��SM��	�ˋ�HnN6�v��8����)x����3\=�o�;�^F6�e�u}DIf�|ԉ�h��Ç�딷\;�o�5;��v�s�rƱ�d�?2�[u���O}|�7*uL�s1ۨ�UҾSM��K�.�[��`/t2m�3N��vz�l�Q���0ݳzm�|ˀ��g���y�.ʙ\%i� �g:WQ-�5��z	S����6J�n}�l�sgT8#0���Yֶ�1*f�[��9(U�ś4�a's�(e�t8J��U?]i�u{EЫ>�͈`R�c��>K
�f��xp���=G7c�.v؄��p���v�r�*gR�*K�k�*{Xd�N��lwH&�<�������Hd��m]׌1z��t�+��*��+mq�+W�1��A��¨*���ȼ�1#�v�`�Xhʸ%x�4��Db�E(�VB���EƘ�c�U�Y�(��AUb�PPQWv�
f���Q��PB�FҠ�[*��Ȥm�nfE�cT�,*T+�7��QH�iFEP���PE6�11UH)R�,-�DF`���RJ1H�PY�H��Z�E��H���j� ����b��X�*�V(T��no9��y��^�v �n�]_5Go8�0

�'
���E �[���__kE:?�]҂	D�^{ޗjt�{ژ�!{�%�R���fC�}�/�|�ƫ"w���JŜYZ�J��Z�Y��Q^.U���F�x�W�U�x/Zȝ��5l�_K�I�;�H�6-ղ.�����5U^,����<�Z("�$��t�4Ok�E(���woCr�$��i�Ԙ���P�\A}��Dl3O)��;$z��s�So:�3��6�D��ϫ����6�i,}W�WOL��	ք��^�ƞ�Mx>����^&�{'��s��ޛұu�s&�]8ˏAn���ޏu�x�7�+���^�����$� �:vp��a�*ot��IZ/�)>�����k���U��k��)��wK�1D=Xr���M���CG{0�d[�6�#J�~x*�n�UM���r;�S<E@��yM�3�Z�'u5y):�zeyn�4l�CXUZ��\�q0C��z}X;�>�@Q�-����3z���S4�hX��[�JB,�*�F���i����&�9덇�ghTI ��`{�u��@���5�t����~�oL���i0�1qGt���nJ�K��z�l�;-dmƦ�'�Z�ב��Q��*�%[����C�!C��y8F�jPEHؙ�Q-ڡ]��W[��a��KxT�[�U�_I,�UY4C��=�3�8�[*�s?��6Q�H�9N+����-���wρ!%��shΐ�7B����&�<8��;�S�T)v�[�a.y�\��v���V��KA�:�:m�����&/
 ��N���U|�\�*םe��B;��ot=�UczW��䚅yL�8ù�U���=[���|���hx����A�F�B�׎/n��0��r�Il{���X��c]��-����mE��<�+$��yJ�Y0���Tv�F�ZE����a��p�+��s�(��㗘^������8���R�n ��U�Nd�M��@���W&ώJ�V�Z1�вAA�NBO���I�6������˱Ʒ�B���� #�ys�]$�S�j��x���楑UO����$_:���,��e�������0d��{oh�>��Rq�@��V�n-y��źP
[#�"����9~�t�W�yw��¦�P���{�C��]��.��(0onUwL��LC^ ړi�VOK3�Xr랬� a�6��;W��)�8�_r��"(���MY�j�[Ys��x�GA+F�mc��,�tB
Nm�F+>��=��+���unW�D>N{� �i�X�u���l���-eќ(�\�k5׌�2��u�۽�_�w	�\}�'cj>	���}�+YY�;n�Wz2X.�DT�����Dۥ��s�8bҰ��!�ݻE���뵠�E��P�,���O�+���F�"%T��:��8߹�#b�q���]�*�}j��cE;�^�����q��pD}�tw����5�q>w-.�Q�1y�3��7F$as\��L�qǵ̾T�%~��S8r��o`���h�d\l=q�����i](�d�$��'tnɺ��\�(C�qҧYt;Ӻ.	��Z�<7^P�<��2�*7ꀗ�˛�͊RI�W��]V��;m���Uߍ{��ӝ���}Z��U�Eo��O̷Y�&��D
a����s��PdM7�굉�1�Ӛs����4�<>D���?}��������̋X�0aE�\��8C��'.�!�_2NǧqM\��]�3��MD�O��Fi�C�[HZN�d*]|�.4�co8��\�,i�an�N�sz������x���q����W���<c�9�ddT����tL'�)�"��O�ObS��Bp���F�i���{�ܽ��76��#�z���e��lo>�����r@�}V�?k���EԶ>^����T�������|ra�-�PW	��m[����*��ݕ�Gox��ߨh����9ʤ�Ց�[�M0]��������5�cm[I�t��[v��)[؞Ȉ��	����I�M�:{�E���G>��g&z ���:�u��53O[�:��x/X�ؤ�R����x����nk �t4n^?]r��.^�k;{S~ѻ��T���3m��|�`��ބT�ѧ�E��K�-�)`I@�f��:��4�a�\���o����N����]YO��oMJ�̛ɤƜ� ���⫰�12so9�-��9��3تpE���@ˍ��������|m�ەXk�l��]��KZmm�_�6��eU��t�.w"�.>%��m�~��`o/nPɇ=����EV�[+yo�-t����*�Ĕ�u�qZ��7��B����މٚ�f���*n���x��KW�������|�f�HG!��� jܿX��$�g�����T��e�n8Yè�%,���n_K��5S}�5�E�v��Y5�B=]3ع�����K��i�ټu����U�c֧N��/���D�ۙ������a����=�4�u�X����vP1�ɺ5��w7lֳ���:��E�w��r
X6
�;B�ٽʡF��w�g��ꮃ�TU���;vk##%��x1��ռ�g��Vkk^%"��)�֟ɻPn��x�;��j���7��э�BƎ3nf�O�"�����!�'�s����vћd���g��\V�D��U�68���Rg��7����~9ە���xM���*sk7[�;Q��^ֻ���ZŸ�&�tݳy����-.V!d-���:y@���pie���M�h�	f�<m��P�!�7��:�ߢ�E��W�gx�7K�rlиj���^�#N��3�-�E�k�׼�P[�;qc@�h�eΎ;���x>�]�H�xVtQ��xy��:�M�&��ѷ9z�oHW��'��Ӧq������q��֞Z�l�kD�~�V'�j���' ��h0j!m�⥷H�,�z��Z�-WG���w�����$=v(�8�:�eu�M�,��kk=�̌����w�k���FvY�� E8+��%��jB�i��B���c{aTi��Nɔ������}�8
�DĤ'���t�C��ai��[	,�n�z6��U�t�2��J�=�z�Jbs��E�#�r���Ũ�B&�4�uz�W��.�D z|�
l�p�%&\�Hr�l���O����3����3� �t��XUf���E��sA�|�ᤎ���?;�2m��x��Fy�S{ڲa�+�輶AO��U��j����Jݞ� }C�}�H�>����QgV˩ˈ�D�G�#���@��
��J����U��[ @5�* G��V����7i�ĈΤ����$���&r��a����Ss盖���1ю}��b0�CT����(i��?u�a��Mɸ!UH��X����%��C���3]J��$:!�,�����y5�@�{g.mϝY��n[~�'Ү�v�NI�_V�cV�l���a��C&h�vjI�����v!��3?;%��y����!B8d�{���h9䐁ή�������\�}�1\�w�%^Y���' ��N��ɥj���������_�O��^꾻4~<u8�Q��/e�x����|h�֟=?V���0cWN���>LJ�xZ�7޲����Y��g=_��f�KO�p�O���ۯ����;3l����k׾�������[4�c��eb�ˆ���?^� ��?��&@��:QI6K0���)�Iu56�}w�N�ir�^�F�7��ʸS�%�����y˴��w7q.�{1�E��\�>��.x��>̎۔6�]m�s���o��E�G���7�o�4q�Yh��ִ�:Ӱ��ӓ��W�#��:�]m�Ə��Y��F���SA���i���o�x��3d�����]\��kƯ;��|es:�$@���eniZp��z_��q6��p5c�h:}���Z2�@��`ƣ�D�gڿtX�1���Y奡�h��U���Zw+��c�d�Uɵ4or�$��:���]
�՝z+��9Y��B4Y[4M�0�]�p�M�k�xg��!�V�� 0<�M��I�N��$�0-!���4w2E����@�{U��z��E.�w"f�>OUO�e:�_R����x��8�;S�]�?��]�j���;k�v�>�јj�ǁ='������}Ӯ�����7~���#��vm����,υZhҩ���'	��@�+����Y�����~���8�j���1�W+�Z������p��@��R��?�.,���1������w?w?7��:t2���ߙ���p�s.wB�m��r�#�Ҏ�o��I���Y����s|�Ƿ�h�Q�9vB��������ߧoɺ-�ԼzS�*�@��Y'����Q�WUwg���n��{î��N�:�F���o�O�E�������X�sk��<��f�r��0ȼ�җ�K�]=�5��ܑN$>�p 