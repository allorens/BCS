BZh91AY&SYb7S ��_�py����߰����  `]�� RQ#f��  B�F�,n` ��M(hdn���� 4�=ݥyۤ�%�% zT���G&�64�� � ��N̎@d ��2: ���2n  �2C Р7I�2�)��/iy4}.�W            �=#F�U*�&&�2i� �12h4ba�~�d)*D �h `di���S�"D�@�� 0M   i�j�� F&  ��	�  �D#D��#L�2i�O$ښi��)�m H�i=*��# ML M0�bbuv���{L�Y3f`wACQ1��h �h
�UE���(w�*ϻ���f0�~��@�( ��dP%���iUU`O��AHSq�x�J���>�B��M������ǻ��ۼ}ٵ=>�ss�D�̲�H���q��UͰ���/��}U0�1�����ƕUӪ���9���4�3L�4S[�wK������mo�P�l=����n9[=�1�[�^��E���z9'n��J�
G����H�D�t���UD�A�2`�O%%7U��#q3���9��^*�Vs��-�E�u��F�<��G���ҼU�Rqea�2�{��1�G*WNnlIMJN�M�K�JF�9��½�%��y�OIBT�M�)��ґȍ����l�_�r%zA;������<���ķr����")�Ìì�7+V0��fl�����j�[8Y�2�l�2�P�zY�[���i�<�c�$���'F�#&�D����Rm�Iג��Dr`��Y�e>3�T��gfg�L�5�f�dRi^�z^�O+���5��;�9���K�U�N{�H��{��U���y��w<7r��5�>��s�ܔ����U-�o~�o�m��oW��Z�����,��{��ۻ��{�a�����o[aլ�h!� ��=nMnM�7L�W�������]�<s�z{")��ì!ܓ$�3*�ʪrU�D�NxߺMZoWI��H�Hu0���E
-���/�^�:q(�l�2���!���p��M�Tٱ9"p�= ��V�V�<�g��rk:�<V�k,դddd�N�O%Ğ�mJ�R�ԫJM�"o�+�.z��l�[=�OI��=�l�����!�1��uIFyȝO��-x��憝�&��9S|�x�ɽni���G�mi��=;�鋦O�[��d����'JF�=�9���v5<p�,�D�ʳy!� ȐdG���'��׏AӒ����s�o��3�]Ǫq���8qA�:�q�|o_�D�z�Z��hx��:_K�L�.\Zf�M�:��y3&T�M�o�w3��m��f30�q�B �A��yu�{-�S�����d9��B%��GEi'Jt��8&����KH�V��cD��\�R$������k)xg蟠/М��N}[����-�X��Wy۰�v�cSZ$�-�hԽ_H����	���H���#���j&�D����Ff:�1%��kh�T�Yn5�Ӭ.��R�����a2I�L���<T6��$�����"��8�`��$B����%�7��xp�:VX�e���%-��{�l,����.�|��ШLLV�o��j�i�i�o���n�'i":MsW��d��-!�e{^z�x���n6Yc���ϗ]������k^i�x�f�cߒ��/J<��쪼Y	y�Yl�+)�a��S�h�e=G1���ݽէg�ۀ��.zuk�ug.}�x�v�<A����'Y#4�]�GpD�I�7->!a;y���,)��םF'���9\��l+vn�,��I���i�~�g���ؽ��nvS.yv옍:�D��k&���{V⺹Wus%�Y�ϋv�k����ݬ��]h�6S����G �X����O��a�(��p7�yrR���%a�����v̪��X����T�F���s�Px��_/��܅����З2Y{�O��`�{�M�>.n�$[�Y^�h-�����O;�]v��T�$]����|��V$t��s4n�h���DQ*��b{�I)f#�s�ۡ).�o��JB�X���̸�������wG�ռAt�
������Je��k���q�UU���Um��j,Hձ����Yī!�i�^�t6yθjZ��B��h�4pU!!�D��H���N��N�!� :6�L�7g����o%�+��JF(�,�ɤ���yb�Iq���R�����
b]K�"�2͛���kV;-_2Ev�+��1j�Of�K�z.��nk��y���
�ʙ�1����H]yw�"2�L�^��!�p�4����i{�WM���ٸO���/r�8��5ݽTm0Mf�֩���7�������d������ �,������;�IԵn��Ņ�r����Vg-��Pxm|��Y�^(^5���:>�g�W1�{t�҇E��r$��3��0b�w|��Lx�,��y>Ep{��吧�U���;t��ɳ��k�_vWEY����z왮�U<m�Z���f����L�8���>���~����E×���#q#��p���=�Y����9��y�nw��M6�v�����3jd���)AvPW:/:�$	_c�T��]l���r�Z��nGT*u,��2F�Ba��TEc�4�kN�n֊�MŶ֬���Cܖ��N�f���-��Off`~��\ʌqVWx|��u��+��p�s�m%nO��eb+FH��ɦ0ş1SC����.���Ȭ���do�P����@�mI�%�y_�T���]��r�RU7��a��p��XQ�v������sjݱ)H�V'������f�[¨���bؔQ�ȷ��]��~�q�i��d�1-����cp0HC(��0zV2��l�Jŋ(�\��|k��%h��瘶������;çgM�	�v���r�g�u���Z�l{�XWa�Y��+(Z�UV]!�W�b� "���r�_�����n��Ƣ(���˓�Ӟ1�(�_�M���MO���蝎?.���4n|��UT9R����>g���9WU\b��s�V*��UW�;U\2h�D�j���A��]Q˵v��UUTUy�s���W���1U�i26I���

H)�1X�&�h�5!�@�)�m��گ|���[�9�U�j����dI�x��,P�AC.`u��sZ�h�rf�Z
j��\Uq����*��wj��]����\8�c�g2S�a13	�a��*V����UqWko{w�UUEUUU��HCFMi'f�p5�@�@�Z*js��6���Ҫ�Ux��ۥUUX�����f�
\�U
��$�My�U=nY������UmUn���UUUiU_*�kZ=4�C&��Uh�Ѧw�=UUUU�Ҫ��ݢ����UmUsF�2��޵��Bh�4UcIq!�OO��>�"��T��������u�nv�";�!���0y@D舘%�A�&͉�8lD��pN�l��N'D臄LDDL:t�,J�	�(JB�I�~����-�>�Z����U�N�L�X4F��*��
Tm��e�{%^WL�b�z�x,c�GK<�ۊ�W����ܵ��,�������w\�B�T�Y��K��n5� vJ���ƞ^��oq��D`�	_�z�fЭEdV�䠈<�4(�*I($c��cy�V��}�^�Z�2�}~��&�q�_�o0�n�'b�K�Qϒڠ��w*kbʇ���l�ѩx��xdQc7�	�l��H(1����Ky�b+�Ǝ=ɖ�5�4]������I9�Ϳ�fff`$,���Ē�������Đ������333��333u�:I�����|Ə(�I�"-����\2� 	���-����("j�Mb(��ӧ3C6p�d�ύ&������.">+�1Gˍ����(1_5�(G��㤜
+øTZ�
9��+�W��F,�(YK���vo!�Mk�2=�(�"�I�K
�!��v��Q�+��8��p&�!�r�$�w�p�å�|���a��"8R)>�i%�>�l����ޱ�^| �R����T� �(Mqs%j��#
OK\��1eub5����Y�D�mH�ɪ��8�n��:�
�m�'�g5˘�Z8�P����>4&����iQL�D�W\�mk�Ł]j��A}CT|�PQe`Q�l}�1���O��uP�Sӈ�6�4uJ���L�dO��0ldDC�jA���e>D�jc�t��%qq|�ө,s�O�o�b2\Ka'��iL][۵���|5�b/.`��J��O�>
s���C+�E�_u�l-�D��a��Q��e�}d��V.�65Z,�]8��͵���II�� ���9\��p�c����j`a�$�}�t�Kx�Y��L�Vʀq�(���F��)Z!9�j�#U�ݨ�����Õ=��UY��\�q[�˥�-^Mq+[�?��1��n��QJ���I�xe�7��T�ʤ.�@��o�8o����NF�ZY�$}��Qe�Bc�z=:F�F�F�i:=:F�"!�C4�"�MD����Ѥh�z:�F�#���:;:G�!x���~�|N������<?GN���pg� �rA���a�I1��;�e��g�2���U���fEUn�w1x��ׁy+N��+rO���W��,�⥽-�=�ԣ�i�;뙯��\��}���H��̀x$�$�<H��� �)" I��I�\��(A!����s
�d]��w� �6p�X.�"W�(�����?�B�4О3��9�4o3ʐ�|�XqB��6"�\��N���+eԝ	�p��܌��.�Yg��X� ތ!%I��)Hi\��)�Ҏ}%��0Q�Һ�t�̚�p<�L@dv	�A�|�\T|��	LF��t�Kg��:�&��^�f��gǺ�n���3)����U��.k� �xL�RI-D89$-��M.S�P��_)V�B��Q� Bk�8�
M,��1?#e7ݜ&HVr���eKa�fLHՋ�i#��"��Q'H8Y$���4�)�����ih�XND!ɐ��0��L�K��n����x�rj��n��Ä����ƄP�|�d�Aafm��m˝����Hh��\8J�0ƕ:;��x9�d�e�Ċ#~6q�䚢sH	7e� 5 �#�<��� sd�d90�S��bjSG��~0�'B��Q��b�%4��� �b)�� �qZ*I!�&��#G�6W�&�'\8�h˴6�:2jI�_,_��
\�-d�Z|Ag	>/��ύ7�Ӿ7i.ey�Jd��swc6�×j\9���1�j�
��Ū�K�:��&@�f�"o�d�)�`�w`7�,�&M�0��ST��
MIJM̛6S�A)S(=�[c�;BX�(�[�CRp������S�y�)h��غ�̈́��>5��N0�y0�sE0�~p�5-(F�����ɵ���p�^XZ4�FJhֈ[����
� ��$�Y��󜊙14�J��
uQ`ꔒu�^Q!��3��<�R%uX�ʄPV#�cT|�5H�GU������R�IC$�Y9�o1��IE��6X/�Mmn�,>	e�`q2q��ˤN�Z�p%��!�.J�9AR�G	��6DUKh�!���R\�x�����P�d}M#J=/�i�9���(����#H���F�IF˒
4��GC���8;F�'�H<t�+Ƒ��<p�M ��d|=�q��X��mh�zL=�$i$AG5���\JJ�9)Q�*�3�5=(�Bк�/`�OK�O2ϚqaP�4�4����L]����݂�aǗ�Qfn��ک���.w+�UF+�d�E����Sv�:ؽBɻ�1dR@�p�L������J�yr�^T��>�ն��QI�5�+�{E��Ё�P���5�e�!,����6���W,�����fH�f[�U�Fk�x;�o�6���hT�:�@�}�2�IrPIrPIrPIrPI"I#��7wsEƚ���ı{�l��n�q�	@B@p�;�J�#H!4j�n'lw�9p Cu��q⪌Va1�İA���'�>�������/��,>[ϑA�g�`%&�z�b�#�$=#d`IR�J�¨3[D�!ae=���Š%w�C�]Δz�A�0����71�>/�)D���%�h��²����G!��a�в~��*��	b�� ����#��%.�Hi|�����g�@e��X�Ho	u|�YA������ٚ��i���> �ov#�/�-���M�[@ H�M^�꾤U|�������Ҩ'����g�."���a��$	L4�Dup��8GN#*�>> �����#G�9Q1�sU3��l٫��Ҧ�8Jj)�(�4y��� �C����Ym��+�x�|:�CE|ya��ii��Xqj��#�u���6�(\�����>M��Q'�ǒ	��$7
dm�%64rˀҟ��&��K0��ad��@����Z�ŭ5���8��=	�F%�(>>���|Zj��������)�c�ctu{���yy(��j��J��|V��� ��Y��lJ�||J�吾b�d<S�-^{�y���ZT�|��G��<@M��ڐ�]���AA���]��}Ccv��#��Z8�	V1��⁄�"Uj<��u�3�(T^%��/-�)h��4k����jX���=kʛ@�e��f�T�����<l�cq�*�jE3T�#`;r	�8�
J*R��*�D�8`��]S�BzfG����-ph|,:p�h4������+���?M7*"�Σ��D�|QT�%�g���q�y0e���BĢ�R+P�v����+�=%��f���Ep&����B�2��6�1�R��yWՈ�����O�D'�g�� l������?|Q���Ӥ���j��3Hf����~<M ����<A���3ő���ta;0�9��㧉<i�#�4�oG�|>�GL#"ǣ��2G������a!��������j���ʘ��4�c�R�/�zY�H��nɦ���铦M�xj�_@��o~s�$�I$��$�y$�O$�H$�H$�Ba�p,,Ҋ@/�ѣ/��A�-�O���} �ͦ�%E#_�Pu,�V�8-త��<J�T�p��K>4��ɑ/��m���GCǆ�3����d�ptc�Z4R��Qiu"T�@����҃�z]���'�$�%"|a�H,8h��}Й�%gטb�2\�˝i�{�R��<M�*2�*�R8UWf��1Á�H�V(8��'e|�#}r3�nDD6G��}źp4h�R�ﴃ���	�*�8@p:[n��Q�r��8,�)_#��m���Y!Σ��-(Fu��������GQ�U��@yB��Ʋ �i��i��l��b�J>G�`e���)1������p��$�XY݈"���ř��p�a��D���BӃ|X�ÁI�����mIft�����8�:�R��X�mZ��x�,&t&|u,�9�M>$��Ÿ���WU��X���4i��f�Q�lJq�+X��3��J%.qu�Tj�(�[�iKS/���I�H������_��6�%�����d`������ӑQA�����TtC���pD�b�5�tZ2��yvK:.���7d|��>�x�ױsU�Kc5��ᄮs����E�t�.�#�K:p���?�&YtK�Kp��pG0p3�ΩG�t�+�u��ȣ�+YG'��<���qoHRjpI�>��}p���e��y`jߙh����=)T�4�L��T�&+8r�6�M��'���NqD��5Ջ��ƀ O)���/v�P���^E�(�` ����#Nk��Od�K,��agף�|Lz���,�G�x���f�A=��pCqޭT��a�:�82Ƥ���d���~k��}��YD�-GEFF�DCL�t8|>'G���H���}"�ѳHf��C�I�H(tiii3Fh�>�G���:;:G�����M>#G�4z=<G��������#���0����&�j\I0Q�8��˷����^mTz�:�t�XP^:�j
V�K���c���N�ܫ5n c�F�#��t���^GvKyB:��r��ǙK33+n��ߛ�l������ۗ��N���碼{�-�-�)�ގJ*��N�j�7PQ�B�!�|Eۀe���TjɅ��&��d��۸�MJ�;1�"��˻��:�d�B�%��N��4�mf?�a�Xߍަ���� �bxf+������I#�$p�$�I$�I.J�I$�X"�!`0zv�F�q�)�����70D�K9-*��*�@�� �Nʛl	f�1,Q��bή)+hj�� 	�Ej����M<�r{&*X�:y|A)��ԟJ �B*O��(�<x�WN��Q�6>_"f�j&Hޱ%�Q����IA���8a�A껛\��7��\ ���RZ4���8]�T�h���!4��n=-��*X�%�0�;�dЊ�:Z��j+K�b�p{Qt�h#��C���}���PG*" '�gO�i}$���ڙ& �V�be+(>�()yA���*Y�	Ko|i&�},���i��'��2��l�Q$PQ>�J���*=(ϊ7͸O��;�a�As&*WeEc%t��B�:I	,8mo7���?L/V'��1ȗN.��� �Y"�qE�1�>Kb��S| ��V��#���`�\���8a(�����m��b��R4b�mʱ�>�_>S��08R����:��T�b^��K$�p,�؂�}f)&J��0���!��ɖ|��������m�`يT&���Q&���(Ê�Qپg��n���9GĚI��Y��)~�b1RŊ���F�v���kI;C�2[�B8G֨��tŔX��錅�Ņ�I��hߊZ4Y$�$�`Z�"��j��#W��v�C�r@�q3QoQ�\�ό A-�<R�K��e/�!�E�� �b�h�AH�Pq}-QjX�/~��'$�;Qb�
�1��'Rm4"5B&�cu5 $99\CV�G�(��Z���
G��")xgQ"��Ճ<aZ�i��A���aÃ$�7
ê�4ݟ;���R�Mj��+K�b�6.	���G�p�"_#�6�:Z<�>O�n�j��(jI6H�I%4<ILr�n"�Z1aK�d��/4E|I��m!�T�ѱ�P� v8�� �?Ƒ���'M#���=4�i=$�h�n�F�F����ѭG���vt������<<I��4G�4z?x�O���YnH<9���JЅa1vm{��]��ݻ�U
�#N$��u̧t��wYe��NY��A����l�J���y$�I~I�I$�I$�I$�I�I<"XXY���m7`��ǔ����%� Ϡ�?�E~�ӈ�Qd�m|6/"ΜZ�,��Z���^X�J6ǕQ&��Eiq,W��Lh^,fv�c�*]M/���e!{������8-#`�
>!��I᜵��.�#�R�MAL�ʤ�U�$Yk㋨�8�FAH��Z�p馒t:UGs�pq�&<���V蛰��F�J�G2��ɩ���$��1R$î6˄�Fk��|q�^|��/ǥZ:A�j�(�p }���ι���m�-���o��ID��d�ğ$���`d͈�]��)v�uGQ�m5e�������� {-�l��!�-�ZAָyn)\>�Q�e���> ���Qcyr�y��v&�tD�Y�yY������y����8�_..i��؈�$�j\�hh�zN)2Ֆn#��D�z	V��\,��,,(�c�Q'Q�Aw���ߪ"&ffQK�r�-��c(kQ�n4�*.QF�˂�V"�)D�&R�I��aa��~��������yM�������G]$�Y$v�P~T��
YK*��7������
CEd��6���v&s|&wW`l�^(�J��������u_e�tb�p�$��c�K�t"�y��H�!6uGيWڌ:��_� ֢�d��$����=�"Ӊ�w�Qt��<B�VʽF��68q8g��)�(P��]\0�pp��n��QŴyz�-�eX|>�DF��$)�P�(bKҮ��jڙ���!h�؜1���ۓ��#�\�}g�E��l/��b�!�fCqD��D��h�=p������4�e�F�O&�hǭ�4�6�M���(�4t=8B��$X�"Α���<<�<I��4G���ύ#�����t}� �$�Ó�䍑�VO͵ϊ��k��x�Њݳ"�i��ࡻmV^����0�ݤ���m���F�5�M�Ve��ܔy�x�Xk+2���)�r��P{T��>z��jd��u��e)$y,��D���j�*��D���:�~�=�8�Z���Or&Ց��]6q�
�<vX��t#|�kĢl�'q�L�ZN��7QL�(�TJ5dh��5�I$�I$�I$�I$�I$�I$DP��c/r�QP�1�]�#��"��X���X6D�Uu8؅re��Gs<3��m
�K�F�� �J�e"�U������5��m��(�:�R�ޚ��a_��ۇ����V�g���,��x��%;�\�K�J������Z�M5��!G�!��D�T#��ǵyXӳ~/�R�Qҏ�����������8�q]w�<�Hm��9x���Hȁ�ȵf5ᘳ��| q���������O'T(���P�"rp�(�\�lcd=n`n&�J��`|����|���0%G����cf�%q�,d0����l�QD�W�_�2a1)��r�EQ���J�`�Pr� m) �TP�e����uB���>^T��I,оYBň���_#�֖�y��M�3��C���S.鏮!�!�p\p�,(�n�4T������4bk�gݵʅ����}��ci��D8o���G�x�h��{��� ��
;�����O��+F��=X�����g�-���hӼL�X�=�AF�.��M,�p$����:p�#���JE�+��5,5���G���\�>>T�\�H�r�FPD2j�ʏ�����qNڒ<Pp$��w9Z���ul9�w��C"tTK�h�$����X�jjYg��R�Y�vt�����
#����ˤ��A��i�����Ms�H0���ռ!�>nUl[�RC ��-WkQH�9Z�.��~����"�����C�!J����i��R�gU�>��"�������Y�:=#Ú4�F�4��i<��f��i�Q�Q�ݎ�#K#GC��z3��c�фx}���~:x�7��G����4��a�i����Y� ��~���P?��ڟ8ۣwr|Tք�_4�a�/0��d�5�'f�Tn�[շݣ5*��'���u����ݡ)�4u����	W>^�$�I$�	"�I$�I$�I$�I'�P���A�t�J�Lp�?/�Qh��t�F����,��GY�Y �йa%B��:n���#�_H(���I=f�����Z�cd/5d�����㘉�%�Θ}��GC�ח,�>%�#QU:J�Z8+0�K��y�j+\܊n��Y.!#1�a[�H�DWD�jAؙJ�p�QE"M�d�Y�+�<Nh�_���U/�ʤi�	�.�Ģ,��.�b
��jQ�d���G���N�p,$��zB�4�
���/Y�"����Z��8l�#N"f%X�M��ƚ��Y�:id	+ܑ����!O�����[YR�]r���q��Ue��kȰ_f#��x��1I��������x�l|V��;�׼�-Ho���j�N�}��kQg��L)X�wQ�\>l�]�Y���M>	*��lU1�L��/�H���yV�pW�xՊ�1>�].>��q�����G*"J�����!���_
�}G��c������~�e�]=�+����!G�`��[\R1լD�8	<�肉d���U���Z��ȴ�ߎ.���H�W@��}�x��*��86�����.���bb��ql�o�c���Rx������Z���>_{���wX�J�/��Q�duH­4r��5�b-bT@)qB���Q�Y�
��8Q'�K��(��x�-}+i}p��� �/��K����J���3�]R�:y5!������PqRhk�)���z�e�e�ǣ��I��0�t���D��f��q�F�V�DX��4�4eA��A>���<a>O��xz?��4z=Ƒ���7��Ox�7$xrz���U;��U��;�jM�3d������)5����R��{z�Vd��۴	~ KF՝�b]�PU���-�H�鑡U�q�UvQ�X&(Nm�gW6�����B,*.�;^"Be����UI�<�:�PJ�eF�8r�E��W��fu��甠糰�X�u�M�,2%��T��A��Mc�R�����ML�^ɹ"��V�J�1����*=�X�EcJ�۽��]�C��$�I$�I$�I$�I$�H��I� `0�g��N`�$QU\tQ�T��UO�M��ؔ�/lt����9l��j�/W�e�iJ�+��������q,S����kqj)�G!�M0��I��6kT�l�n���h���p��W�ח�0D�W��}�j����b��T���J&�W:�t���v��1��(c����ц���޶�7M�A4���E�-N]\ϴE�8:S���8a��$��;�65��K��g�Ы�5" �}�t�<�L;�_�E(!|�V��{��xÇ����Ǯj��1��]��q�%׷cr�c-DM�n<��U�ʰ�Dc�8%)�;�2��ھ-m|4b<����=����/)��(bv�p�@.]�_iJ��Ź�<�$��nE��u=_�P��H��X����!�l���3$��gǏ.���g��EC<��јA&�R�BdDNMpm�0����ժ	*I�y�^Q��F�!��/XǞt�A�Mb��kkT�I�4<�<@ײ��k�jqyZi������]�HÝZ�p>��Bk�ն�G���I��(�'�G��ƾ7�7P9�­j�41��3^�cX�8(���GQ�|�Z�E�J	��^7��#�s���
�������GjE>$��qs[���mjcl�J�|�b��L�R�p7S+��f#ʃ��y�]8s�NS81�x�(�?�D舘%�A:A	�bQ�(؉�6%�!��8X�|����O�>DDçKġ>�I�@̩����=ʉ��wVd^L�B�%���["���K��f�k��c�K$�*Ƅ�V�:�ӳ7�\�����R�dT;z]`�3�BWu\XW�t��N�,�cIb*�=��I$�I$�T�\�$��I$�I<"�-p�\�W�U��^�{���I"m��j��,)s�_(F)���^IPb֙�>�Z��ҺX k�K�Z�,���Ƥ+�HKr��봠@��%r��sW����4�Ec:a�NMz��]U���z4������T#N�W�'|qEml�"�E���ܡ3	�4y#j�}DFaǥ@���}��m��G�֍���Ϡ�w��H��H�b�F��ܥ����6��U� ��$����B��G��0���h���
P�:�>+�e�>q.d�a�ǭ�����-��(�p(��'9���Dl�1gvt1�+�&B���&�WD��X��O���1�8���%I����-��z�#��:Ca�4BΡ�n�#��m���T;�d���R��j��>I'��K�"�DSn��s��	ko#ǂĤR�(P��H8�U�;"j� ��#�8�⫮�1���AӉ�1V�)]J(�qO�ސH�M�q4��Dt����>,��JU0C!�Ƚ�w�����:Q��A�k��K��7�ı�E>\<�R�%}h�'ƒPQ����]��̛2�S����^>%yT�8�*8�
�S�͖Y�R����;���fRê���b7�-�+>P2�$���,
�m�ƴ��*����یA�^*	�%��>,�{¾�k��>.Nxf�up�}o��^p~D�%Q%w�UUT ����{ϥ~Ӊ��௬��&J%L�
�h:_��e0Ƙq�]dJ�
P�(J��� �8B`'ip�H�!H@B�)��HA��H�C��)��� BH@0@�JB�J� A"A
@�@� �*A
A
AA*A*Aȁ��J��(A*A
AA�@A�,�B0@0BH�B�#&�+�� �`��B"`��0�$�N$��p�2���8`�`̜L�&$�������L`b	���� 	 	$1ၘ9�9`f ���!��$�"� �&dqa�& ��3�e��("`�1`�`	 8`	��"(��0@� d�& � b�H��	 �`��H	 "
8 $��
�H ("H" ����d��H�"&"	!	�`���Hb&"	 &���!f�H	!	 ��HBa�""$�$�a��" �� �"	!	�b`������f�&�`�Y"!�"a������!�!	 ���$�$�a�B`&�&a�a	���(d�a�Ba�&""�`���� hB@�� a`a`d`e�$	BHR	V	H! ����R		JHH$ ��	`�$ �
`$ *�A A#!���$�&�>�2s�L���l`M��z��0�I �$�k<&:%��c����ï�����_޺�O��k�5�;w�>����k����:��#H�ëQ����gO��Ҟ��鮚���Z��cԟ�����9�C/o�-�s:
������q���}������A�~2EC�D-��?p�����o0�����&0�<'�9�������?�NǗY����Q@P�����yEA��L�׶;W-��.F�(`�'�6_��	����ۤ�� ��m�qv8A�'�|�����ӕ�4�c$�O�^'�����(��y0���
(dȡ�Q�� s00  BP*D*!�� �mՍ�ԇ:a���>=!�C��~���=G Q0A ��� A��h"��$T�� �x�f�yx��	���&�oC���x�<�0r:��`�����h���}�m�ݻ�
�����,�Gܾݿ�}c���z�y�y/P��Q9�cu<�^/�� ���p���H�Gs��َ��=��W��;�Ԋ�`��qپp(�y���OAˑ������`:Ǥ�"���z�@P���W���}��P�d5C��:�D�j���!L��L
(���;j#�匽��'(AE@�����v���+��8�9	�?�a���
l'��&s�C |�T�'w7�;� ��v�q���x�.��(z�SQ>������w��?�ٿ ��δ�re;WAN_ۜ^a��0������7��%Oq������h����'4��#���������� ��s���?�~��"z���aؽ@ue��]��5T�f�#��F�Mi�"�nC�s�\�)/����'��1��	��Q2z�M�.�uA�.~�(
'����=[h���;�zǷ�9�ב� �{��.��<RS䂌p��5T�:�Pr?ڜU:��wB���S�d� �ڼS�?���vNǙ�TE���1<�}������w�/�T���D{SP�@ʜ����{?�]��BA��qL