BZh91AY&SYc�pD�o_�`qc���b� ����b"_          �                            �   @BQT�,  �T�`  �0   @   �                         7�|�)PT���U
PR �@����PU"B$ D%k$���HJE QI(�

 �DAY�I   �Z�R� J
�kϐ���D��@J��Aws�B�+p%��JQww@ݎ�M� w8����	)�U    ^>J( ��� G� ^qQ& �ǰ��y} �I}� :x�yT�� ��- @����/#���   �J� ���(*(��Rݺ$U| c��4���� �� ]��"� 
6���`� .� ˜�(� c����� P |�R@>��}��#����
�� 7a��2 3���<�z�����*� h�� ����1�{� <   ���-� x�@��J(
U �X���v8�@7�����'C����J�����@��c���!݀�w�A^@9� ;�    >})@���@�7�I{�R�}� ��� w�<{h;� ��`z� -� ��B���$2   w�>�WA@�
$
���J�B�T� �����  1� ��R� �� w`�ڀ�`s��GC��:�*�(ݎ@7n�   �O� ��� ��
��r ݃�N�H�� ��, �r(2�����   5�Ғ  ���*RJB��R��> S�Pwn�&�G@Y�*�'S#��t�wEP� ��6    >T� �=��݀�T�X�r݇�A��g@��*��껻�� ��q��         �"`R��4l������ ��'����P      �ʥ(�@     �%H!R�      $�JD�*����     B��iMI5<*xA�ɣ&���2m蟙����?�����?(i(RT]ruy��y�~|F���)��8� �����@U�@EO�D@U��P_�0����?gJ�舀*��:�#�� U񃰕?�QQy�_����&	���?&I��\`1�d1�L��`LqЄ�c�2c3)�2�c!�i�M08ˌ�0�Ì2ˌ�2�2L��c��2���\e4�c�&8�	��e�L��i��q��!�e�\`1�ӎ��	�&2��cL08��)�28��+�2�c��� � c	�aq��	��3�M2���`1��&0�&0�&3�q�L8Ɍ8ɌÌÌ�q�i�1�q�1�1�Lc&�1��1�q�pe�a�e�\e�	��q�q�1�1�d�Ld�d�`�a�1��q�q�1�q�1�:d�a�a�d�fe�\`1�q�q�3�:`�a�d�`�gLc�q�1�1�1�1�d�q��1�q�&1�1�1�q�q�d�a�a�b`�L`�8ɦLa�`�\d�a�N�4Ɍ8Ɍ�Ɍ8��8Ƙ�2c0�2c&2c0�&13�ÌÌ8Ɍ8Ì��Ɍ8Ì8Ìˌ������2c&0�0�&2c&2c&2ccɌ�ˌ8ˌ�Ì�ÌcÌ�Ì8ˌ�Ì8�i�@i�q��d1���&ALdA�Dq�\dWQ� q�\c��q�`GQ� q�\eSL��*i�\dGE�q�L`�fC1�`A�`�Pq�1�	�aGA�q�\`G�q�eq�	�a�Aq�\aE�q�t�Ȏ��q�aQ�Pq�a� 8ʦ��Pq�Ld�A1�dfQ1�Ld� q�`T�@q�q�&U1�LaG�q�A�Dq�]3�"��q�aS�Dq��`�@q�aG�q�`GVaL`A�U1�eG� q�\e1���Pq�\a1�\`�A�Tq�\`WE�Te@�AfG 1�\eD1�\dP�LcL�8� i�Q1�U�@q��AG &aP�`P�\eM2��a�Ed�L`Y�L`P�Uq�C1�C@1�&EeP�eD� d �c ��Gdq��	��@�GLb`�Ce1��\e���Cd1��q�cq��`1��`1��\e1�L����S2c+�`1��L`q��a��i��e��0d1�q���0d1��S`�e1��CLe�Lf`1�Ld1��tޚ������߱�|�;��T��UW�MD�b��4Z.�۫n�RX���[�ܸ�ժ�,�cQ��Kx]#6���S�w`e;�md�lڻ��g3$*��ʸV敹VN�ZY�4xs[8����h[���j�#m-/��d�f�0Yj�V�j�Y�`!P��]jr��H�2����u�=���[�Ks5˪�eMn�S����"�tj<���,������c�_�����Z
C�i&�XDm'�l��]c�KA[x^6���nΚz,�	f�ԧ�Vٷ2�TH*�-��ɍU�����(e !���P���խP[�dј�b`٭.L9Y��
E9�qFi;w�j:��2�^n�h;Zk5Hph��#,ֈKc#Ķ����+���e�1D�Me�b�Z��$=w�7%�q:�����y��F��N��FeY����.��6e+ˬ�R�-�-��A�V[!�fV�`j�
�W���+�/2���wyGt
�X+U���zwlޝ)d.��,���^
X˖�evN���Ien���]`��vPh*8��v��F�	G%��l\sL�2[�f�z�����@�Ÿ�W�X#�(!�KՎ�=��Toffq�5r�f=�{#��1��$�3N�3�n������uPz�v��&&��d6cF��Zl3�e��B�6-�&Â��E�A=�N�p��0�nMmK�N�9uz�����3X7�EF�͹)�b��0<�9l�-��W&�s�b����tL#�e��ci�dO,X�%��(��c��M�ݲ�.�F1�v[�.�ij`ی��M��7t�9XN�vm䗛  k�on�XʙVU�ɗ)�&m�� �TŲ�ǇH�z5�"+w�l��i�3lؐ�m[��R jNP�{g�Ppٻͧz�Ch�cu,>�V�IL`t3NĴ�Е� V�Zs)J@�J*r��2������sV�Ea��,�y�9��ܭ��B-a\�8J�2�b
�QZ��<���l�����w���]Y�!u�Ct�&F�-�jY�Z���ۼ�sP�H��y���Ѡ"�WCeY:Ѵ���YF<7o1��
��N���ׄ,W_�ner{�^���J��yvK3n����%�ǘE�7�v+��WR�\���K��۶�-������4r[>d�ܳ7 h�Pm���7x ݗj,f�y�JQ�ۛ�䗐Ղ�����&Mp�y��B��6����E�C&�vscժ���!�7`��)IY�+4�jn��f��,#[=�鳖N��!����R���%����]�yG6�ˆ������J"�s(Au��D4���T�N��)-�^��wP�<̷{%��5��ñZPup��meʽ�UK���K�ʍS5n�[Z&�Y�j��V��1u��dٹK5��f�F�n�����q*z)ѭҲ�/JW/6��ڙ`U�n���v��ԩ0�I3(��VN��R���׎��xټ˺d��Iu�f=��Ź��&��Aԁ���]�j鑖1�8r����0^�j�0[ʻ���{��eo��͆m�Ȫ�Õy�M�݊[�f��66=��ӵ�w��EQ�f�-����f��j�J���-�H�T�Ӱ�[l�*�l	ub]��tܴ�bolR����Ũ-ʰ2�Ɏ�e��
Zh,j����Q����d�w]��n��pŘ�n��n3/m
�~ƮLǒ�`����p�{0�2�,!R��Rm�7RUa�l� [�Z�e��A�2�<h�on����÷p$�ˤBVM*n���Y�-�*gQ�ܼͲ�^n�b��)؇�.]��SJ����e�̏+N���C���^p��f5m��1�vM_-������/ؖU�V@h�Es/(ܧ`l�4�ٽ̒7a�"Ҷ-��I}�3^]�.�����4ϞjJ�JW{{�Aa�̩2u����w����y
�%�*[�;cV�#�X��	(�	P�&iv�v]f�Ш��^�����n�f4�+b,��.��`�Lb��&�����[SU�Ү�n�A-:Y5�)F��50���m���z�I0P5���J��Y�f��]Ж��&��s3h�~E,���n���-�.��vE[�H]@�2̶����i�����Nˣ�.�F�*)؛K2͋�wX��j�׻���2�I�^�)�1���5JZ����x��tw6E@����.�D0����Tq�2޺�����6V�fkц��ܽՐR�eaW"�6s�c x8�2�롕gv�J͊����V�n���e�Q�ؤ	�,���Z�S&Y2J���H�)�6Ћi�L�p�ߖ	���f�)e)������VT�AP�jh[�!��V%n�_�rG���E�̕��Ȏ��+P��+��+H�>wN��{����c��Ib�$����)�ո2ݣwa��<��1I�xj�&�&�XPm7~Ɖ��-�p�.]wL��t����9mlM9Zf�< �z�S��U�v�	�N͌������"�;�J���jH]��nVPT*�z���{��ͻh�@zJwvx���S�4��"1d76k�f�W�X����{[y�l:f�o:lэ�:5�Z�M��B�jdRa"�Cr��i3z�}2�lc�P�T�y��ٍ�ì:�T4�]ޅ[qIz����]�X�Ck(Z�)�Qm+�5xd*�IYsI��/4��dZ�R�
����4�mk����V�P�e���7=�Tg
F���Ԥ/j=`kX�k�	.*gS���3j�����۴�ɱ!m6L��cVv�VJe+��
l����e<��t�3�]���)E7<m��[u��jۭ���j�#�.��������^�Z��Z�;2��D�OM����l5i�H�����f�V�~ܗ�P�cjɕ.@��f�afS�e:ܒ4@�plf�6��+/oo
�Τ):UH�7���wwww IY�.Rz�&�5n��W�,[��n�(��7���j�lӉ�LM=��OlE�2�J.b����!�m�a�K��w$>,ю�YX&Ѱ�e�8k,�&V�se�*���*�3+̗��J��6��wY�b@	��fO]�C��$#m��´7�ۙ6�ֱ��X��)���]�(+�3.��� )
��͖.�t�2�:R5����-Zi��aY�uw�جlf�de�b�l�ZU�#{n{�ǖ���t��8�طh"�kh�-�;�&�P�z7
��r�m�:��71���U�ic��j6|�neևx^�̭�dy��{�m��::0�5V��i�SVK��h�kbWtp&U0�z��*M�:؞曺�ܽ��P;Ɍ�8����n�6wR�j3����rcl#�.��:ۤ��IXj�K`h�\���ܙr���M6vEⰅ���kE˸̱.]�X�)-���T3��}z�b���{��Ƚ B�������lhmqQ�}�p��}WY ,鸲�uȭ�ZNf)wr�TuV��zj݄.��vi�ţ*n\�H4����౔,��.]������cJ����73%m��+���SnɸE҆��O4��=��x�N}��Lv���F+̻X�j����9r�,ad��'r ��J�4�sP��Zk&�@��pn���)ӖLU�X9�lF��T5=S.dJ=Bm�HK3p�Q�2��&���̢734V�i�l�'r��卨h*�&�8ݙxe�Ǔ`�u�kqlm�*e�Ǥ����N��Ұn���ږ�����gk36eҭ�|#�Ff���8��{l��N��%�GV���M�ƻ�un�3pD�-�5�M�$�9u�&�X��8�lB�8�E�f�V1r�f,�h�{\�bP7�	�"�{�ff:
]����A��Z����WX�w���Q�[(;+N��
���llr�dQb��ŭƓ������B��Qht;�Xpmm��
��Q�������d�1YH���2��1��V��i�	MqŌm輺�͸��iח�;�H��^�����v�#33���ۡ�v�sm,76,ݽ؆�Nf��b��Eޏ���T�B�3r���/2�f��7sbNi���Eu�ji�WN�f�a�=�׆͗�L���D���w4�Ǒj��*U�1�[p���˖�X7�[y7Na��7zh ��ٕ��SB�;�ZN�{(@i�Գ&��t��sn4t'J,˰�l.�)z�9��2�R��i�,9r�@ƚ���1e�;��Q�6�c}Z�`Vmk^��o3.�n˭�mfx.� d��kn���k�l��+(U�S<��1ͽ���%&���e��B�B��U���A�P�	�Fwkaje��7$L#��yV2X�)�N��r�v�B��`��U*0M�S��ri�n,7��1g$����w�M"vb�
��51)1]��Vk�bcn���6�a.�� ��2F����+5J�@1�jl��F�d��K��֨��TT̓N`w��6�Je]%f�x^�D8�MՖ��^D��7�V���ڛ�T�&��ou��*Ȅ�g��*H�"�X��UX���̛��7�eޭVv�37,OnX`�b/wG��b�؆�}���y�dI<�qn:wRY��/M�w��o�����֡:���L!Ӽ��0<��hI�q�n�L]4�
w����d�X朰�u���x���Wĵ�z��{�8tǴ��R�&��� ��X��l<[��H�өV���R�f��j�8(mѧ63i��L��\4�ً��IG�d�I6�JMù��y�Z̥Q�j8p*y��ڵgH�V�w�k2���Xv�&P�'4).ظ��bL"ɖ����WnÖ��"�v� �G�4�-ws�`ƌµ]f�YpV�h�,l��{�宰e��DY���l�MU��v S���]�~}X˳��[CD�1�2 ���sA�x�f�u)B��j{C+4ŚY����7b�u� �vs4�����	U��o��ʙ��=��1����yd^�MP)y� K�����^�/1��1;�)�{e�R·^�;&n�c5	a�BHQ0�읺F��V�U"0,�El[X*�;6.�@m��
ov�*]/)Zr�Ŷ+A��a.��91�WLc�������&�x	:A`¶�s<�T��Yj�m�X+4d9f�E�d�˴+�����Y�[�Lr���x�S�˶VT"�jf�.�Ǻ�%nD�F�"w�ݛi������гlV㻣sl\6�su�`ٽ
fM�!�T�5����Bl� U33ojϦ��4���â�Z`�//^i��ws*�)D	�ł��3�3VKjf]ݺ�ܕ	���d�����#�{�������.�op*�������aX��L���Ncڻ���Re����:F�j(�
̭�kn���vM�����Q$<ԧa�z����i����QN�el,5�ٲS6!D5)��r�`փ�����v2��wp�fd��]i�KR����j.n`��kC�y���`-�EШ�Ć,*�m���i�+6'�͓{�*�ű���idב� ��P6K���,d$%����j�,2����Iz����kkrL3�ܸ����"de���R�stZ�2SF��Z7��>S.+��V6��F<3K���{q�|�
�d��W|6���M�5\�.����E��×v�+H�t�G=�.�����b�b��W�ݽj��-:w6�Zʶ�	�5�
�W��ʻ�����n��E����E:v�&��[BB�bÊ��p衱K�C�+V,�O��+C�5��M5��:������hi	d>����U���W���j+ݱ�mf$+Q�hM��ੴᗎ�42�*D��Fm��[F��[��y��T� �0
r�����X��3V��6l���-aQ�����rTˣ��R����h��ނ�uaR�e
C$��T��X:���r�
��(��s"�
����T��{,Ex�<y33^�d:֤�2�x��vED���D$!T�ɛ���ՓNŗ�-��Z�ш�U���sr��Kw\2X���e��&�R�lz��Y���o`��{MHA�YbnG��qU��k[��^-ݺ�N�d�٥�!��H�t�@�jqݐ4��G��Jn��tVP�]Z����b�'-���F�4%�G�c6+(|S��b7�3:ʲ�V�����'�g����e���'�%2A�Dhׇ��y҄�X��Kz6�Lb�R^$��2�R�|��F�'x��6I�9���ɂ͈{��-(d9��xm��p����rVㅘ]�ua�����4i?E�]���/k���'	�|����|_�fg��3ģw�Jc�t�;4�}�ثh�I1��^�~�$OȻf��-�NiߋG,�*̱��|L,�V�@�`�!�-X��㒊O�N�e\��.��yR\>�rP�Ҵ�^��z�ױ*U�[��6���(�آ���dOB��Wj)o�t�ZQ��2��G3�!#��e�D��3��+���b�)��qg��d|N�4�r�QIJ�V��-Q)n�c�S-����fj�I�J�HD=���KV	c��Z"d�s����č?�_�Әy�?	�p;�K7ȧ�j�ǫ�=	,�.��BN��O�ߴ:��aU���O3�ӈ�#��SI�',N��Ե.�佪�@$k�w=o�2C�d�3��w��R:�?$O#��+Φ��K��?��/�V����$I���h�2��g���W�[J>Gy@'�K��=/��aGpfi�wG�ͭ�r��S8Na���$NP�~�����w����H�%�4��/K�Y���8�:H'�H�p��K�!�ϳ]m�y�^��U�2�A՚�.���!�k|uI��^�J�O$DJzQkAx�pae:)�%@�O
�Wbt���[�Y0�9���k:�2��['�P�=���p��*8哄��ޓrV*
�¸�68�o}fb���9�mĶ���w����7ܑ*�/'q˩�wē���9�C��c<��	xD�X�����!�z(�I$�?��8i�?�#�i<r�$u	wEߪR������˒� �����8��O���(�(- �@� ����4 Ћ@�R��"����"R�"J@�H�B%"�*�P���H�T���J��*4-!B�4��
�
��*�#B �(%"�ҫH	BP	@�B�СH�B�PB��4
�BR��-"� 
J�P% - �P*!B-�P R�!@�P�PS@B��"���(���"SB)B�P�4�*"R4"4��"�B4����3]�q}�I�9�*L���f�Y z�c�� z�:,#ŇV��+vq�2�As� j�<B�(w�+�ܝ��wԇ�}���қ�9��F����ď$pdw=Ǔ��Ǻ�=�\h8�e����|����:��S�qGpj��;� y��B�[�K�����i�
Ԑ$�=!D4%�4h��m}	�N�4�AA�]�:��	��PY�����A���S�D8�L$�`Bfh$���	�� ��¨u��Q܏wb�H{yy	�o�&��3���}�N�$Դ���d�x���
���Z���pq!�z��FF��!�MG�|��|������w�" ������ C���o��S���q�AQ�������]���_D/���?��yw��uh\� �A_+yӞ��β;��N��jА��ˑK�U2s�R'H�����׋_+�Pa��]i�]�/qv)䝛c��F��b��(�/]kr�F	K�T���)�I�4�6��vá�u�
�'����/�N�[����m�&Q�3�R�P�v�S�׳1pʐ#�<]��߆)������(JIru�c�җ맦������*��2��:�Uպlsb �%Z�mgd�U�A�CcQu($otS�u��7�+8WK ݍ���/�E{��b�T2�4��_\Ut��(|���!J� �t��%Ԭ�	܎Y�M�i}d�Mf���}�����.�Vn�<��pr�&nj��8�p��A���$6����m�<���ث:=S_.�6�t�j��U�)�qe'K�t�:��*/�΍�}�l �؇W</�V�l:̓M��v</L��j���t�D�ȆtM���d����7TeN��qνte�d��*�nܹK�=[�[S��`Lm�aٙk2-Fէ�tj'VoQCn��]Fao/�)�[{a\S��zwAೃ��CU��vj"��]b�V<K���Ͱ����.pJK��e�]��3N)���SVB��=Lɰ��������������nݻyv�n�]�ݽ�v�۷������nݻ|v�ݻv��˷nݼ;v�۷�nݻv��۷Nݻv�۷�c�nݻv�۷n�nݻv�۷nݎݻv�۷n;||||y||||v��۷n�]�v�۷nݻv��v�۷nݻv���۷nݻzv�ێ�nݻv��۷n�c�nݻxv�۷nޙ۷nݼ;v�۷�dd�������̮6B[��w�^�eZ;��V�<�N%�]��S���M	Xf�gy����k�u����jTTP�/h�ձ+�cp�Tʅ��){�5�ޚvv��g&y�DtS;W!��5�V,�{�\��� �t'^ڈ��ۋ��<�a%p�X����lm���6(�iQ����G3�w�ջe1=��/��CK��bшxҽy���ng���Y��4�:��}]o�-����������iU��z���R���7�wCt�o3w���3W;5H���	��Ch��t�B{�n�����Ֆn��"h�Ùv���T*V,�9���ʜ�2��l1�Z|���bk#S�w��T�->�6���b���=�u������}���
��:����=nnhD�ל;J��h��y�oEf� ��kV����x��66+������HK�x;�.�n�ӵO���#�7��i�x�l��r��wH���Yu��e�^ɯ���5��|��6�d���md^�4N��#����#֧��y�ݜZ[�:�;�Uβ������̫n����u}u�*�۸�ȉ�2	�^�u�N��ֺ��+7�`�=��]q��q�H��w���ۧ����Ƿon�;v�۷�n�v;v�ێݻyyzyyyv�۷o�흻v�۷nݻgnݻv��ӷn�v�۷n�]�v��۷n�v�۷nޝ�v��nݻv��۷n��v�۷�Ƿ��{{{v�۷�nݸ�۷nݼ�v��÷nݸ�۷nݽ;v�ݻv�۷nݳ�n�;v�۷o���nݻv��ӷn�v;v�۷nޝ�v�۝��o�]�r���|�z3k��L�gkuf� �c������>\�_K�S�J���C�_��:^��-�+�8z���lN�ݴ�R|3u��[4�f�`S'$�ٲ�I��x4�Tb������˒_c*f�~�0��y��u��hdeذM3�G29y���'o&E��Ix7��Eѽ�Y�kE�m�}�t5&���w�/nw�*U�`Ә��w��5v�h��3uP�b��ޠ����*qy;�'Zt$\|V�x%`܊��%ml!n�H�Cp&���u�R^�w��ͫ�F��3�,��{R��7|%����.���2�;�23��vp}�r�_nu
���J�VcE-\1�j��:��.j��`�r�W�3n4��WN ��1y+�0��oK���JY�QT{�B��١ug5p�+�G�X\�V�3�v���e�{�%BX��XoʎcX�ݙ�R�&�������ʗy�.G��N�݄`Ѡoo��ygWz���[�N�1q�{l��:z�74���{�Om�s���[��p��8������t�N���nY�%��[� }���eK/E�euZ;�zfm=�Ţn��PWhλ6Jk��9�Z%�_N��q�G�um��u��O_ g�xY�Vu��n�A�]��[��Y��m��\�����{�~�On�_���n;v�۷n��۶v�۷�o////�]�v��۷n�v�۷nޝ�gnݻv�۷�c�nݻv��۷n�v�۷nޞ��v�nݻv��۷n;v�۷o.ݻ|||||{g��nݻv����۷nݻv���;v�۷nޝ�v�nݻxv�۷o.�nݻv��۷n�]��nݸ�۷n���v�ۦ�����ƶƶM&W�_������f�޴4;�4�� ��a���ؠu약C&sz�]VqcC�����O�U*�Cl��ڛBh<���뙒My�,ct&_c&���8� ��JU�\�G8��y�u5ۡX,�R�w�·�JW[|�
2�=k��.n-�z�X�ĉ 6e_H��x2V4Wʆ�7 �C��ҭX崢�v)�;�S6/# wβ��Ԍ�F�zI�v���v�s1!��}Õvy9�C�o�[ه�iv�=\i�=�GIêzʶd���9����r�I#�DL��T*�����ݩ3-C6�ܒ��ɐ�j�{��|�!��R��$����v���j�s�IV`�"�n��28���S�{��f^�̚kEOb������Xv��������Vw4����Wt;�g�����C6��7g7��:���N�RoOK��3�Z  ��s��d˽\���x���R�ý�w�&���ɭ,�}㺲�t����򞺘�'��%�t�V:�_����YpWb9���{r���*�v��d���G�n+��\�9��c�N��Z�xER�+՗���N��mqhM�'=�[y��3+�������wZ�0,�0�΃u�+��k��b���Y0(+��Z����ʽ��ϙ��P�G;��q��ev�K���=��W�����J�Ւ>�z����r�T���=����oE� ��`������r�^k�۩�t����Ʈ��)zԸ苉�����Qʳh߷l䄅~-ؙ���,ݻ��Vt3��Z� �"��'j�4�B���r�(@Q�D�h����cxn^uХ�d*�5�YyJ�]it��xJ͈S�uY�`Y��B���&�WWv�w<���X1�R�%E���vt��+f�f�={��W�
Nz�H��I�*VG~����q���3\M!���`��Fj�]Y�v�$���JU�|�����U����j�k�1
�uz(��_�۹XИ}F��1�
΁K/�Ӑ݋ѽ��{2�U��wQ�˘ܑ-��k�[[t��,�}V=W��m'�ڽ��WQ�ݭU�#L�'*_/{=ޝ��p[�
�n�M�U�Rj���I������^��7��u,�Y����Ŗ)�FS�I�D�X0�R�Oh��k�u���ղm�,�b����0%u��s��v��B%��8�rՎ�+�M�4�-u%���}s�C�	X{���>��OB� �@;dx�xm�mqzX�Q�=��\)�n��Ku�a�����eG[U[ҳ:Vgu��[]`��m��]�[���rRx��`��y��-�p^��ՃF�(o�o�kgB�I��ܹ��m¸�0ƙ`�1_��|���巚�B���ͬ��|=�Lw��	Բ���@ڇ^������Y����l���R�;�rp�.��+A��Y����e� |'��NZ�Ǉ/�\��СJ��&f�3{a�z�lն���ta}�!�&)ZɃ��j�h�9��F��������yL�yέuY�I�&j@���^��ku�����p��7�Z�S�WD��+1��zJ�B�q�0�7�Y��O�շ�l{Ǧm�����;�ͨGm�7�m9��δ�{Q�s�n�^n�
�woR��B�ѕ�5�׻+�^-������r�,�wU���֕��e]v�K�9�!�з� �VJtK�ֵ<�|5�c��C�U :�Wu��bR��f�Vs�歔љP�e�h��s^�.����{�8Ŝ-��/�z��n
��[p��V�ԧ|;�󐇅m=y�Vھ�{����u6������f�f+�1�Cr�[�0fi��ռ�3�7�� �H�y�9}C]'�	�ʏ*�z�ݺ��uhU�� aB�8`��e�ɉ� ް�p�u7�-i���M�S)�Ga�sY[ˏ��a7�²��]u�^;Z�n�p�A�&3z���*�0���L`��q��m]a�f�d�Ԥ��E�~Z�W#�q�ߙZ���Z�;3��c�-�\�+Fr�{�2�|m��)�����(�����ft�Ǝ���&ۃ6/jJĠڦ�ۺ�y&�����:�xm頠�{b��j|6m�׳�P;9����}��ִnP���{��ջ|�vU�Jg%٭!b�g;�h�b��N�u܍镨��XY�wA�o����F��N�ֵ�}�N�x�y1��עͪ�G�U|6�#ٛdlj���c�3=��y�=��;Pmv��E<י�uq�[����H2�ᡣ�Z�P7�u�X�Uǈ�N�yx�x4�\z�0���UU}՗���I�Q7���Wh
��UTLoHk��u��ʅ>=n�ԹY�Y[�e#�~Ա�̈id�E�s���zD�5"( ��拪��7��.�\E�;�n�4��{+m�ۜ��Q��ʭ�N��t���2=i6��X�hKo�G�vm�V �Ms�-V��`����
i�:Uu�Vɫ+�dtX�̚�{2�������Y%��^�)��4Q�-��,V���U9Y������:�
��wc�����cV���K�Tfe��콻�x�͵CUe 7Fm�p:�����[��jT�A����EѼj�V
K<����u��We{z��,N3���9��Np�`BQ뻮����.���9ò��R;묚�;������w��ܴ��;��m�m���sf���I�rAGY)��OCz�N^���ՅW;9�w��g;���;s5f�:iP{�
�vMÝu7c�[g4�o��t���/m޻�}����xofTAޤ�ͺT�s{1_GKf���|�{ܨ^C���D������7�r���ېR�곚�s9\�Y����k���GcoG=�U���gI������G�3� n���K�Jh�t�_.��0݋+r�[�l[ۖ�.������k���W%6��Wq �RIl3;��T+s
"�Z�wN�ة�Ea	^S�]��Ll���M�;�&�����o>s��m���h�R������L��mvi`�Oc��"�X/�A��V�R������3ksMben�=��oՒ�;ORA�zki��x��b�L�`��u
��Z-JiV��
�o�{��E��ڹ�Ǣk��%<�OvY3yȄS�iP��G�����J������z+�;�����%lНee�T��8��=�����e���'/�4��a�S��Qq��ʺ��}Ȯ�,PS��Uer��w�;-.�]Q��0�T0�'�M��( ��xVպ�O�̫�v�����.ꨊ5rL[Z��^)�0lw���U�h�	��[r�Hup��sx�a�ĳ��8Bt���$0BM�POò�;�A�Y����{wk��s�Vq͒�a����2����{S�(��'����N'�^s��1ʾ�L%WzsI<3hK�(�0<�D�H}Lr�J\�xy̹�u��ɕ��	�a*'{�]W=ɵK�j���I��Kͽ������3|����QY�
�!����v���]f��G�:ݲ��w:�=��f��X�������Θݷ�W=�`l\:NCp��*63yk{V*}B.��)�ܫ��60_up	-��vN=ږvb�4�WE+yص�/7-���}��v撫����k�����[�4e��O��:�,<x�縩U�N�nT�(�ר�^�[�.�uh��vm���R�V�GV�YSl����ж2]fL5��Z8��MJ�ڼ�7cw6�(qs��
�fP\�i��.\�����Ygu���2�V�V��������SM�E�9����yH���A:�uڕ����;�����VZl���(�&�j�3&�6���%�3��0�<�7�� �	7��Tԭɕ+
�fޫ��16�`>[9�ʓ�7/������z-��;+u����#t��	�qwi�Z�\x�b�b�Q�᭘0`ł���\�e�aΤR�;�QŚzH0�y�6E�r���f5�\��I��4:ۢm�.�� �W��|�]���*[w���7v�L��ݦ� ��L)�c[�t�7�R�S�tn�fۖ/c�hR���K��e���[�P�f�е����p^v�j�%�rr��;&'3���:r�±�g���d4�[�R�[<G��j�dˈ�����k��=Ɗ�|��E��YR] o���H/.덥M�,�Fڝ�󷕞�t�-tmf��B�3���-�)=�{{'�亞��5��ì2�jYެ:��%Qaݛ���rq��3������ml%����2�;nU���"�5Ҝd�+y�)|�������,kG��#�wwW;��W��_�f�+ֹ6�p��������+�v�|�Ն]꽓K.Ĭv�gyu�E.�\�x�:�rjԪ0�њ���R���s�ĜYҁ L�Z��|(l5��T;��l4F�}���� p�J���N���m���ڪ٠���y��V��֏@�3�|�'�����g��/`�/ �|�Q�6��e��ö��l��D7�2\�Á�t�΍��n�q5�e��ㄌ=o��G��5�%'TU!�V�{oe���KV3Y��kZ��t���YC�Ev��[���ʐѡ�$ ^ݨފ���ݺ�)�w����4����pk鷔��j��N�.՘v��1�d��M�^8��̗��!9+����prkh<��I��o�a��w�@X/Y	p�jF�^��km-E[Ҹ�n�b��o.��e�/��T�ծ涣�j\R��o�q�%vƯk6��8_9h`�Jķ�)o�rDQ&@�ԑ��.�+s��8���ʬ]f��{6>���)�̧�-)��ѫ9^�s�k�yθ�\o�_����@ �۟������}�*���o���������I��D��^�9�Eƶ?�y瘅��n�,�2f$tf�Z�q���C�o�߇E����Ě�h�OT���O&��7�~y��[��,Śƨ��β�6��3�,�	PnK�Uk?ҿk��Vz��K�tC�ȩ9]���H�غ��	ㅟ�����������l��<<���`:���<���]��6��I�4m�&u۔p���Xx��m�{'S�\-���V�GF�`�#U���KT�����v��R��k+�uٔƩ�QW=���덷�cS��� ]���Q�H�H3']d�ă�5�]�֩@Y%�S1�s�'E�	�qs���5�v�����+�n͆�(���!��i~���~O���< �ѫL�N7\�f]
M�����4�s�5k���^�<=��%N�f�C����CC9�����S:�n-�b��х��m�@�I�u���>֋�z��:� �l$�F�,���\�)����C&(j4�Q�Z�ֶ�F�`Ikzاe��&��Wv-u�ݯ=tZ;%��7P�ИWE!
\�,]e4ף]sN�τ�dm�8�ē3E���f��=61lJqۚ���A�27Qj9 �����$v���ZC�ą:2��%z�9���Z^�sG�ۇu 0�(Aѡ�땋�Ū2u	j��NLs
հ�"�m��%��%Y5�A���Vd��SU�vv����$5�#���P��W���3�>b�ԍ��"�^jJ�,�t�����U�v��܁�R�N�ۊ�Q�@�͌�Ղ��8��A�9�K<)���q��ݻt��:+O�cX0��'[�ó`'�0�ŊRg��Ɔfŉ�Sv�
��v��z��sv����@�ݸ)w=��8��& �Y�{;WXw����<���q��U�S�Dq�ޢ(�Ÿ0�Z�;X�X���[�AwT�Ҕ�ؽB2�L��7M�С��jWB)�#ş�1�K��jxwd#t��H^e+�D�9�Tkn����Eqŭ]]����c��n-�gVINx8����n'8M��l���m�˰*�=���[}|?����'+�z0o
b)%�$SS1nZA��o�����v������["��ui��󋳩F��Z�sűe��e�FXe%Kc,��DV��<��u�#aG��(0-��6SsR�Y���G\Ǌ��)˛��Z�&����hwll%�u;eX�TI\���[�Ɲ�4���i���5�n�]���fw)�2Lbi��l����gf�4����b�up`�4�M�ً)��iQ��1��"^F�|�o,(TMFˬכD�*6�=�V�a�qnl�jF��Xو�:U��ݻW!��i:�X^Ks�X�L=� 4�qN�/Mͱg�x��{:�����Ԇy��v����>;{����$��˧�\6;���yS�pn޼�ٖi�qeHj�m��6d�<�0�*���[F`G�A��'�h�Eq��0]k<�F�T\���g\�GI�M�x�W6[�
�p��X�Gc��ƷGl���
CG��Kky�Z٠�]��[�Ycgt;��;���c�va��G��R\psvD-�Xպ7<a�}���բ��ϱt1�м���NQ5ܖz����P�wK2�`�H�5S0bV�L�I�WIw�ޘ�݌c�o8�'ժ��h�+�u�H�J�(YF��&�5{6d�ǘ�lPt�ƙ�����U��Ǒ�"rc���� ��QNµ�͎��mnN��h1pV��]p�rr嗜�q`��WgV{$ZA�s�v�It!�K\5t��Ik*�h�-���(�n�u\���<��ND밺.y����1Ly�ׯbN�3q��}>x����t;����(yw!�3�=�=��[��u�S�؁{�/6�q�n%Z�έv��6�69�\�7f��'���������7:�N�t���R	;X�в��j[�]�@�m#zٗ�t���E7H�k�tr5H\Fj�VZ���1�vz�q��m��l����bs�$$ֵ�ˡ����/G7lrZ�W'�W�Vix��;n������lx�ݬ3[��շo&���usq��H�Ci��n�rR�w�e�_5��E���5q�]��#��c5.&��j M���L��S۵�n1,;�R���6��@7hL�.u8�r�D��[������L�n9�e�[5,
�5`c	0Q`�;[0��\E㗴S����Cz �VJ;F�f��T'nc�P�2)���hęfˍa��m�O.�հ��ȣohc�L,s5�R�11b�.1.�m��0+`��*��.�6�X��̳��EM��ݺ�L/-��Y�\�!�b	����z|=2Bb6��j����m6��
�٩��t�؎)�4�O\pmûX4��mqZ�����4��A:Į�+���Ol�=�7j�Zֻ�-�a籄9HnqI���=#�����]�E=�Sb��)O�:�jV�n^�P�JzQ��!����|�������)X��^��4<qmC�3m�Y��+�N����+��\GODU�1����sW�KS��5�a�x㫣Sܗ�P�q�m��p��et��ݑǍ�q�[���-�Nuvn���!4ô0�i75	��I�i3Ì�����8���nܨ���K��g����ټ�	TU3`j��l�3�c=�C��(�-to<�,�m���]�Q�*�m�/b���Ux�6b���r>	��٬�`�,Ѕ���:�`�ډ��+�ǎ��Ƙ�ɉ�Rn"�L��cv	M��֚P@�6K����ػN��^x7�!��Ã	N#d��8K�X��[U
Լ��J�GR`lK76����9��p�j�Q�zHUǤ���g���-P��-`����7��M�h� B�Yh���a�H9�%u͒��8�����>;�wݞ9���]n��v�W��<s���^8����L��. L�t��5d-�崕���ٍF�0�M ��u	��xNݻq���ق�������;��:�N`(,k��@�n;��M�ٙ�hPv,CY�]Q��CՎ5�N0n����o�֓ˋ�� ��`o�B�f�ն��n8712=
W��m����|�=�� IL�3���u� �Q�H3$R���K����,�C$!ƗL����q��va]m6�L�d���
��"[��
d���,�6��7i��;Zr�&֡#n��<�366���T.��'Z��j����m	�"\��A��e7����n�I�����n�h�ng7/.W��fۡ�9Ӊ-��#G;fM�/-d����b�9�;:��6�h7V�ƪ,��ű���ئ0�W �[t�̬��CGh]�&�f�0��]Κ4YR�Q�n�ZM�D������~��ŔN@�8�gr]�+�3"��b���r/#���jԻc�ax.������@����9j���N�w�^sOb��Y�pE�m��tE�v��n �c\�r�G�v^����hc�;B��e`G,�ٚT�[���V�C
��Y���F{y�jɝ�zN�S���ay^>��c���㱛OKV�<�n�X,V�ktk=�<te��g�X���Ϯ�,m��e`R�,��*��!F�+,��ב	�����`O͋��θ.{D�'J;D�M���&-�^�!���<�6���B]�Dn�;�����ѽ9�q;�Qԗh���m��^3��뗎̓^	Ɉ�E���f�N�3� ����E�g��Vs�G�����R<N�;�Ÿ㶆U:��mj�������cc�g�1�V9 mH�v����=�����rØXgu�ٱ�!탴�[Y�#Ֆ��DZT��t��y�ۉ�<x��z������]ϲ�
�kOn�X�q�X�W`m��fg�)!��v�	1�*��c�̵��9q<GT��l�s�q�S/\)�w[���j�c�J�+��N��:&:޵m%���+��a-mb�b�d(�ۜe���`\Џ�X�:Թ_����R��S��f;K=H\MI��mu9��1466�Ś������-�Wtk��33!���6%����nsٚ�6:���k{	��cP�:XFP�b��;,�vf�Z�z�^���$"]��D���m�pм;qqV���Wq�E�J��@��٘JH��(U�=����U�M2��Tc�dC0�:��y��n�7P�{p�>���70��v��������[�ve�{<Qۑ^�z�6Wn:N�H{@n�w]�u�	�y��|������Q�Jݷ=��<�q���.c���:V�gpmͨn�Ý���t��&��]�uIb:Ӝ�bڹ	-+ٹ��3h�t]���ցln3�xr�Mb�Q�gD��z�w�$���u���ʝ���mu�']]\c�Nەl��(�G.��ˎHt�cf�f���2�sf�5]����l�����͊[Wĵhכ�6�rG�]N��qC�U��[v#$���ݹy	�۝p1��c�J��iĆk���Wr�n.x�uݵv����s�����+��uׁJ�9⮵�]ՙ��3�n���Y�u��֧U�2�l��WbfR]M5�4�����3JA�]�^�ƙ��P���e�u��!P�kW�B�:TPn?�c3[��P����鯣}��b��[gca�phr�Z 94@���kvۮ=t�m��:���_������S�^�l�%n�Ћ�t[#I����|�/���3��M�Վئˬ�,h�efj��"9|g�ig��N���v�H�q.����ڹ�%Sn��f�vvN�8�jG��%�v���	�;g]$8H"]��(P���y<�b]�3�bݛ�F�����O'����j\�Z��k�ؙ�~�'��_pP�����Z툠��1�	��um�XK5��vQg���490=t�'W��Mw�<�ĉ	o���v%�����>|��|~w�'P��uo�܉
d�:U�r�ȳ��)�b��Q��l���ӷ�g��nݼ<<<<;{gn���"ֵDQ��3PMDYj)��_�'$���`����fxy{v������������n IRP�92BY̊��ԁr"�9'L���DLֲ+S|{{|q��<�=�>�<<<<>�o����j�	��*��D��?i�Z�+���/��9��ҝ��
ws��e�]��,.�%H��w,3U�Vq8��#.芀A�
`J���S��3��N����r��s�vG̝�d�~=�K
@C&������ے�)
�3�1-󃓜
y����3ȧĸ�Eq;)(��3�H��:mS��gq5��E�G	�H��RD��n{2��sdx�~��/�Q2����͒dO�[�ڔ�drIY�fFf��,+����L�Z$�,�q���ӡ������j)b%��D�8�@�J�1��됒���ܝ�w�OgM�P��^q��͘HF�U�)���h���z	���А��up�{�ǯ,�̩!"�
�Y��+��ќ'-�C9'��\C-ٺ���<��q�{�bQ��f&�G_c��xUG�'E���h�]*�0���5';�����6��1+/��ϐ�O/j1���o)kf���F�`�R6KZ@ӯ1���G�ФXA�Ŗ섷@�p�5v9�y����p)uFnKuۂJ�eK:��y��\��7/[��<8EN��3+�[�}�$���U�;�p�4	����]ܯy�t���(^�����GG�Q�x����i㥆}�%n�WLtZ��WG���E��T�?^�<<�z��Ŗb�0�UI+e0��4"�\�+"���� �D�-(��܋�V������6�"�3�ٺ������\��#Є7\9g	�{n��E�����KR�.�-���j�{zC{��l��c+X���gj�{�t�ewr΢���ͅ� �70՗2�m�5�<3��z�D\�:��r�p�-������7��N�m'R��vFKs�i)Ln���@��XjX�uR�肕��^Z���,���iL�u���[��qV���j���sN�WF�욮7]!l��cg=��L\u���ѹ�ŵ6����n��r�v%�;v��;D��u�.��,�=�k:��Z��F��8|��۵�lmq�t�6��d�g�����u�75�����(�T��X/!V�W[��75�3�k���e���f�Bܲ�;=f��Mu����Et3�����Q���)�7Fc���6�U��8��k��C�n7i��ӻ	�\@����`�6���f˞�i����c�����f��Cɓ�ǌ5�J�CV���ŗ/m��o-�]�Nzy:��m�=�%�����!=�Qu�gg�d`��&��v�*�fD����R޺�`sձ3-�l%��	��l�Vf�F�1с�s7a�5��'����h&ǉ��e��^u]�53ڑo:�q��put�}����v��6��X��\m���d��4�k�JǊ��#����v �q͡]�,ؗ���|�rX6����ӻ��B)W�m�iV�"�%��Rۉ�Ȝw9��������Qg����f��c֢6�F��E�,�b���Ij�U�o�n�a+U���R��%��V�a%hf�㸙�sqq��4���Eb���T�t����JUQ��YZ5kJ!R��VZF�C��|��3�[�僥y6�r��x�M�J��=�i�8!�O~���<<'���l��ד�޽��J������$4���M��T��q��߉�\�q�l�\��&��MH���F5�P�A�dƾ�����Ǧ6늘�aR�f��CR
�_Ԓ��.7���'v�~���[>���
eOOo0q_�:��>^�}�j�#�>��'��\��T'���]��*����Y�}|@L��5Q�(�����67vW�%�/b�W����#�S0&gla��b�!�%����[�����Ǡx%���[Ӷ�kV�)c����%5��߿w�K�����ힹ�CZ��O�%��;�o��W>U��ϕH>���2i�2��
��C�i}�j �wq�0���\��p�P�Es�n*�d��"�۠�3NdΫl֪{��im�tirъ��#�faU�d ��F�ӯs���qˠt4����<�mɕf�>l�w�o������qя65p�.�#>����t>l��o+x|t�꫺����T��[$�>K㯯.�Ѹ����z�{��hNxU��*���B���v.��s�7Eǫ$-b���j�>o�]J�Q��-��X.�C����K�J�5'
XUɦ�b�GWjD΄��D�&��'ϛ�T��֢�3�F��Ƶ@�ط���Z�[G��/>% Kw����{�L���w��WC�U��s�ם���¾��C"���}|a[~\i��́��P^�46��d+��>%���%[���Eg [ 
���Q6�����G��u��;M鰛�rw�NYc_�+hA��$�ާ�&�L���S�����x�_�����c�8����L���ʌI����i�"���4�nb1�"U5�l�f��-���j�5S��i��f���g�J��o��ϟ�nwe�Z�H�&Tϛ������K�������zKq�y|g�n��i]�v��Wak#��������R��>l��^����S[9��|C�[oV��=hz���R�.�h�t).|���}�O����v��f}��V}�FkD��E���s^�0lQ����I���EU8[5M���YN�����*?5��_%��۠��}t-�6[���5��}��l-��"R ��_�H��VH��6V��/�W�o������I(ֻ�E����e�Ԭ�K2����]�9;��[�(T��m���s��9��F�Q�>C� :��vt�[5M�o<�������8�bW�.^�}�F}�z6ZgR�A*Y �	L5���"�s\\WP�۱qq��Ǟ�2n��ǭv�V�%s�{���HC?z}g��f��QWr���跗v�?��c��z}�+|9������-3��wF����Y�Ĳ������i�^Ԍ�Ug�>��W���Შa"�e.�nI�*���e%������_՟o�Vi�|[5M��HW�����4���?L����2/*n'rsٗEh�����s+j��l��n�gj��z�z5]U
�S,C��-]c����؜�|���յƛ۪�p
d�桮�)m��
��4Ү�id��o���2�Q�go�k�j;J����׻��&|�!��+�f�\�3�v�M.'Ļ ��� C�E<�K3`��ڔ�"Fs�ͳr����j�swl@�\AP�$�ZC�l�F���`���n�E�7$t�>7�M3�6q�j��-��wAى�;[�7(�l;t�]Պ�=�6�ez�:\�K,�LM��k�ɦ�-��[CB���]����m���=����tF+��r�]{C�C�k��^���*ͮS:�E�{����~�;iJ��5��Q�ƶK�^�uQ�p��K@I@�%y��]�vXޚ��&Ԋ�����ݹ}Y������Z�~��z���C����}���!����c�wݏ1uTǹ�]�wC�t����|d-�;=Ju��R����6+7�^ϥ}u��G��t՞G�d5[ŵ��2�yY����X���}$�ϻ�y������/h��
�Z��o���4z^ 7]�fX<)���k�Ǒ��.��=��%kF�T���=���5����[���?|�|���N�k y�@��a��6��ëR��D�lXoS�`Ġ������RŌ�,X�3��wjp�e߭�j�;�b"��U��
YL7y�6}S�_�CK������W�n�1�����,�%O{AS�{�%M/@/�����.Mkw�hM�=,n�ڎ��W�"�P�tj���J��%0ʽ��Eνx�X���gĖR����i���!��>]�MJ���9�����q�}M�r�Y����)��z�
������F�f���q��C'.�#/2Jѭ�U!2��. ���V?��h�hw�{录M������uJ�n�>��6���d2o����!^`�x6E����؟g�	g��Y��y��o��ƳE�8�P�U(n�&�^��jx�ݿ@��MPZ�y����M����n-�f�CV[xo«���o&W�-�}:}�� ���վ|�6���2T�i���^L�Wg�e4X��������'��_[�ԇ�����Ixk�����!	&���[-�o�l���?��}x�lb�ͤk�\K�>!��i�/#���A(E�&Öj�}��w�>�K��u��EU�6��=�\i^3���#>�i�>�<>l���P�ˋ���b���3��ew-�:t�{'-���N�G���6^],�U�kt�f��$5$��j�<���^9���C^r���U洒DzNՇ�R�gi�0� ^��Y�-q���ºq�JXmT�M�SJ���ײ������S�^�!����z���_o��v����w�Ϫ�����|*C��$��k�C���SζwO*�vϾ}sT��<h�G	�-��-�U�\�"6�oPM��^m��7>��95ל^툺mJ��lT�����ʦ�O�w=Q��4]&N�ҽʦ�d��+�_�>/{���>���I�3S|�T;����V�B�ԡq��Sx`9�w}K��p�\t�)�1:V.j�U�6\8��^C��F�%@��0�U>�Zƒ�T5�7b&t�]�K���'t�|���/��c-����Yە���b�>}��_�dȻK���0�ps&8�KWb�NQ�<����ysz��^^hS����l���Ͼ�_Z튒��]���S�U��k}%�K��c2�Ե ���6r��<(C��"�`æ�W^kFNvKd�O5�p�g͝�'}���Y_TW�8���j�~�G���}M��u�.�`ʭ���zi�7���}�R��:*_)�o���]���6�USf�|��w�q�sy�]�	��3�?=3¸���I]���v0�cϞPݮ�oFop�Dh{�:�5z3�/���jCT���xXΕ�@��܎�ڠ.���O�_O�ش��`�oA��tAȳ[�3��f���PC�;�M�8����+��	��6me,�Rk4+s�L�)n�C��,�:��ku�[݌��K��*�>!�[��S��p�mV���qٳn�g4��nKv���y��jC.i�MX�M�,@�i�:�F$i��z}]�k]���;q&�G�����&�LF.�Q�7^jq�
�t1�����=v�aD�"r!ͬ�h��ͮ����o��>C�+�����SM.�d��B5�K�*%fnil��%ZЉ����ϟn6�o؄�hL���סu9;��w�j�4Mm�쫠!K6R��)��SL�+n2"�V済��R��y�s���ڜ�������s�}����ׂ�)�(^k��-S*�d�6u��n�|:M�-��?��:�7��
�&Sj$��Q;>EYC��V�e
���.�'wخ�Ahh�H]a|P�e�E�Ĩ�KJ��߾�WR}�o�>�zx���݌����}1��4F���'xb�;�~v\�|y�|Ex+/ 7e U��Tcqp7KR;Teti�rئ����&|�=���ܒ"�+q���}mwv�R�>�z�dT�Н����_����.�?lU!������PU��^����-�gp�����y��pV����2�d i�W��uQ�0���:js��fٿ���h���2&P��B�wk}��-d�1	�J���a�h� ������u �j����7v��\�V�]�3�����>����i��)���dUg��@>9��4�^�U<���G~ݯD���
ػ>����M."�5g�V�IH�
����������f�w#�:7��g��B^lᚎR'�73�D���~;hƆl��#�u��a,2�jdʰ �Kr���̓��Z���	�r�.c6���S��;�w�m9ټ���}�o��>^`�zS�T�O�fH�M��nL߳+�4wA�·����y���8�ݪ�9��z}!�l��2f`�0�{��~�2�o{nQPjZ�Eo�Hlӝ\lL��>�J��q���yu�v��/�ݾU��ԯ���VH����r�FN�Nճt���̛�fN�v��j!Ip�
�x���gvz�d�����ǘ_K@����+wlEN���3��H����tT�M	;����T#�k7i<Y�Rʚ���[��u��+�\u����փ�t��]���Z��ޕY�e��[۶�n�u�>̥1!)f.��נ�9tHL��9q;�X�z{W\X�'j�l���U"�+�u�Zk��{E���:�&2�:�M��C����/0U��+�qe��31��r�8N�;gH�D���^_J�Q���U}Z�-]q��֍w��ݰl.��+;p�k���Z��*�z����VF�5�X�4����{Gy��������9��ޠ��+�t��Z�1��֨�冺�;��*��E��s�<w{Z�ֽ8z�b�q�ǩ�{�i��n���b�\��f�G��ol��;�ҽ���+gS�����s�+:���G7{��H�{&�})��c�}N��lu �k����첻�b�nw6�Dl�ɳ�ܼ�n����FfW��v�ݪɝp�f�_a��-"r��%˴�h����X�vp�\��Rܻ��k��e��L��a�Yn�/�^����L2��s���c9�0B��BӝJGG�&K+Qu�v:���w.�)7&+a��hPi����ԇ���>��as.���}��ow�� X�||�h�('4�9��* K�a&!�}��{�#�J~������4��<��.�=|n,��v�EG �eEL���/]��P�Qi�ָ���öyt�OO���������-����I�q�hÝB"����Z��@D��|�G�&�B�N�-LQ=�=��<�=���<<<<>�o�����O��NA�7�E�_��,��wH.TkB����ѡQfk�>�$owo$������;������������������nu�TM?ԕs�U��(���EDW(���w�9�0���>	�e�"��(�W��:E?r�"�M�@�uYO�*���/�!N�A ��"���E�I9Z,"9EȤȪ��}[������OE��������3���烒Ur�}E
��ȹAO;���G���*�:QEED\*�AU��P(����R��?���|����M0�� �;(���TJ��9E}��l�VZ����0�
���(��Y䗩��.W�L�OP'>{;.EL.}ө֞_a�`�5�����[�|��X\Xe�R`��T�Ǚ0�Bw�w�0E�Ǩ�\�l!�/T#uz�g�&���I��s��4���(է"E
�;j�0�A��^ ���A0�#>����������T��r�Mn���y�hU��'���]���8�8c�OdyNL�to�.Us �?����B�˒���cYij�
�b\�,�!�3Z]�X��DxM�6\. �rS�(�T��J��������7U<	r���s����t��Þ<\ES�d*�8&g�C��yA��T m�lp�;�;Q�lЈ�=��r�i.b	�q�Ag;;����cЍ�f�e�,Fb�0��B�5�Xv��|n��dR���̹�`3;�vv��X����?`@9h9
�ES�j����(�P�x��s����l �Zy3��媡�V{nWmwa�����D�a ��T����5귂�&��W�S��{p��tw=^�J׋��nN(i��3��y�
/׸=�2�ip��e`p�o�U檨��p��P�P��ƙr��$�@����,����y�$�����Qay�dh80����	��ԧ� �R'Y�?����]��^��6˭b0P�L;�2�y���>�[���F34/�l~��<͸�\iz�`{r�y��P��ɻ5������;��S$>j ��A�H8�p-&k�${6��v��\����?8��S��f:�`/P� ���I��S*��AcT�Wz5�~W��[ �~eԠ�z�#�m����9��똂@���Z��!p�Jvg�{M��ۇ#|�`Mj�
�$�p��M^5�5}���lt����3�br���5R�s��*���PcT�T����(M0	�Fc�4�����gj{}��������-0s��R^G536��w��1�^2�RN3N�5JUߵl�L�˺�5V"'6�Fg��� O�z�� U �Aj�:v��k�T�bfx7˴�2n3Y���2��uue��3�u|���ٻ���"�b��U��+�³G�[��rb��	�-��ňbˉ)�)�x�*`%��3K�:e��!fh�8 u�m�c	����ѷ"��l� �HT�BRj�V}�5н�)�ce�'��Hu�m���3,�%&��,������y�V��$[qp�ؙ�]ه\�\n�C"�+aAM�[1�[�3,:��Q,�m��a����ŨJ�YV�Y�KQ<�&x�S�)�3Q"u�Y�]/Wb�tn���t��H��?�SmM�Ml�+��-�T�؄tn��̂�
��N�×�EU���_��g���K�3�ݻ:Ϊ/�&w�L筸
t޸�Y>�;����W�`z]���5H��PJbf�!D^v�����@����,�p�9S��^���_i	�����+PG|E�<�c3U����� �偪p�j�9�T���/�!�w/p�����5:���	�A�`r��C��.ݚ�[��j��w3�9M��:aD�І:g��:�/}*w�L�R��3�W�Oʃ6�`ŀ�p
��M&���T�;yU!�+k)�b;��|6��U[9�螱����L&�C��+]����j��.���<������
�òG���ŗiJ�ŷ���n8*�p���UR(�I��l	�����nӐA�,�E����]�2���\F竦�k���^ٹ�+@8on�n�����UЮ����}�5�H'2~����mֳ�b�`kI��o�|Ɲ��������7I�a�X�E��s�X�:����v����Z��!��'C�B L |C�G�����`!�lӨ��W��L�R�5i،��@�P�*,.��y��V�Ni�� U;U!�AN&^���8���^nLv��U�sW���c��k]��&�;ET47I$���a��Y��� rRA�;80���� ܨ�]b���s2jt\X:����f���Y�6�7��7]��-c���n���8"�7׃9���z��� y�ge���+6_��&s�)p ��@;Fk��T��S��^[���O+��%��:�0�W��E��-�pZmCrh�X6���45��ϖ,�Bx�I��Zy�� D[�.Rfz�`�>ތ�y��j󅘅�S�n߸��"!��@[w8r/�9b����'b	�N�e��� ��	f���8>��fӈ�[b�ݵ�s2jy�u�<�z�@�L2�O;���La���=�9�ژ����ir�;����F��.7�k)�&�%2k��ݧ@+�ʛ]YqQ k�OS67������⾱k�ш?�.�G���F״l<l�{��f��I��a�u�Nv�5Vd��w�=��fs�)|a��PFj��9�� ���y��&�t�lf�B����A��)݃����f��]sW����m0r$m_��t^c>!e�g��&�3�e䜂I�"��[@F��:WJ1�����g����o�ξ�̚�`]Cg�3Ÿpj��S��������`Ѣ`
X�9�	��h��!D�L4���&%7U��nX90���"�H$i��v�L�-������vu��z�w��ޟ)�t$��|!	<�zSH� 媓3�d.�h7h9j�J��>�bm0�1�8,�qM��ݍ�z��j�;���+]��U�W����n���XFy��^b5z�N�� �*�P�T���z��6�=���s��4�`��%w��P�R_��xԙ~��(��'�;.q���A�vk�8b*��^T�t��vc���Xbv o��R{v:�mE�ߦ��ѳ�hW_��ү��)|y���S�ۆQg��]W�x���kI�R���&G��Ed˽	q�3|ɋ&Y1dI��4�H�H�"&��o��&580j����A�vR��N��qZ��T_���]K��g3�8����L<ES��I�cO*1�3�>���f"m,�䱬�l�'=���W+�X�Q��{<DA �P�I��9)-�奁=��5n��NXj���oӛ|��7<��ש���B_��(q`[9Ð;�pA�v��BHh9a��&}�,CucdS�v3�r�����Hb>����T�f�;��%��@<2*�܃�Z�@7i��ۈ��DU3����9��gI���A�`k\8�ۇcT�x2�P?7`�!䐷u���8u9T���hu�eod^{.����y�S�;y��襓B�jI{�'L��+����m}��ߛ�Ϣ�^��9j��vO<s�D��
�t%��'؜���T�x�g���#����1��"�����V��m�?>��q�(Y�-.���6�T�B?�ok��6���+&ob��=�(�>�n��4.p�:O�q���>(�},���dԨ�
3	@��w��A��u�k����sv�`�4e�]��L�르�+fP�#�h�֍�L-�E��-H5c�5�6��U���815���0�1�OB<1�W9��VjE��Ke��������� t�����jK���[A�]P ��	�M�i�-ΚjZb��Y�/�v���7� �8�v܎VG��f�qxN���\\�<��nnD���K��^���g���/Q)�m��E�y����u�s2��l5��7J3-GL�Cש��}�82W�`A�&g��i��ۍ����U=tu�fk:�v���j�mm�@FK�ք+]���pϬ��d�X���A�ܧc�Q�@d���u��y��au���Aa~L�-�P��>���3�s� ����pXT�ȪA��:>��6��|�o�S�:+=�B\�� ��gL��P � c!v��2�]ay	kdũ�p��9� 偪p�\���j�벸Vg3��A�b�f>E^��x��^�8,'bq�?�^�@ �T2���q����8=�{˽0mJ��`��"��Ɍ��ȼ���aq<��`����A��w�^��m)ۼW��l���$p�ǈgP�%�d�<\��M�f���i[�$�g`LRE�H9H5R	����i�]w�^z�{�.b��o�ا�-<�5䗞��z��$���bn��`�?m����5��������踽QQ��P�u�ﳷC��Ƴ�/��WG���!���X ���c�����Muq�raBU��$2\n_���h�D��t2
jH!D�H�!N�|(8 ��ى���U_]�³8	!G8$��;��� Eߐ�7W�vv��M�v k�t�+���;��6����"g�C(M�fnd^NU�P���A��sT�;j�<�aIÌ�B&;��V�`�(�,�}bf8c>�R�uZ����nb�s(��m��F3?.b����Ʌڂ��v��i����R=qZ|��KX�B�}��k���y��R�!�[�U;��p��.sG�.<G��A���M]kR�ք�1Ƃ��\�$.�D�M�g�w���,	�NX�vsT��	�O�C�;w��r��#�d^�ysOBf�C��z�`�����.Eū�ɟ�v\���W�8l<C���4��uj���� #&<AmZCM鷤E��N���.R�gv�����Q����v�oo?%�}�3�DfW)fE����V�z;�w�r�9�J}�w����Ro`�j߯� �z��Pgƭ�E?�s��f�3��R��5
4��� ЪP���!�{����k����Z�^g3���@�E���9H5#��T��˯'��N2n�*���<�ۊH � g�Pێ���y3���a�yŅt{ǫن=>�<l��-Z����Q��N9�AuǮ0z�i�d0?��S���=G=Η��t��+Ł�����;�/�׊ D7dQ���}v(٪�ݺ˸�'7��.S� �{R�m�45�ǯ^�������s�n�h�5S��to�V�괸^g3��.�7M�V{w�1f�r�m��b,�aͬ����@Z��+�sf��a,r�g1?xe���W�9| ���
�0pE�KQ}��}�u�:�����	���v���`ib*�j4E�j<�y~�lEƪ|P�v�����h7j��x�&�&L�-��^���8K�}��0<���U;�٭;�z괸^_3�	MX�mm�Y��cF���ǽ7}KX��ƇkNvA� �9��\��pW��|�cۇu��!\uT}&�£(U�>{��σ�ŀCI� �� �*P
*����G?0��_P�޹���1h���ڮ��Ϣ�|J�`A�["�]FwVἙ��90�:dc�sF��̘+��mZ}Iբ�t��]�|.B� �m]���6�cH��j[r.���6����>�6�)��˂���ES�Z��gʟT?i��9:��\e	|��׻��bV�90�0U���q��9�8#�V��<���������¾���ש�+�e�gI����RgÁg��<�M'H�Z���'��D9�N!Ʃ �>]�7�x-�=u�"�r�I�@�<��Z�8�T��
����O$�Zt����n���i�D8��3O��8T��t���&�l�{�-��!�b5x-$k����t���C#�R~�7��X�^p�,�赜�k��W|ι���pA�p����I�f`�0Clĉ�у��h~�jac0�,�{����u;���<��B����^,�e���b����P�ٴ/v�怍�Ԥ�1c��G%^wd���W;������3l�V���P�v"���k���q�u�����;N��ک�E��nY�$6�g�=�]ؘ�chX��{���W&J�OL��͛e��U�Ff3�v��d偅��<1��L��ov�6��h�yn-{J��7ײ�v���t��d�yS�.+���j;�@�ڊ�iݫ��f[����9oA @���Ɉe��ָ���¦Z�P�u+0��ӵ�1v7���"�q6.��qM8wԆ��5-����y�p\u:��k���إ��n��������_}���[S�n+�V����[F�ZvM���'��T��!ѧ4���f�'l�����P��� !��E��!�*���{j-S��*��tU�v\4,�����P�Y9Mţ,�q�JW�̏!O�8X���+��|ޗ:����]]��u���NQ��3k���47����ZT�����PS̾���yeu�T��I����j���4a�9��baf��ѐ�����K�+�c�8Z%�s7�/n���N!u��+o-����tf�4��g��^�On��2�����eb�yC��WY4��TU�)W3;�����rv! 5�rYX3r�&�C��h�����t�+�P����6�f2�>Z��_^ʽn��.K;㋮�;����9�`���E�N��(κ.��Ȉ��AU���.U[P�w���<�/O���o/////����߻���*������R2���r��a�u�p��C�.H�������n�^�^^^^_G�o�^�萣��wZA]uɑC�Z�$�W�v�������뷇����������{�h�KQ��Z4#�;';�D9ȋ��w9'�UU�p����l�8S/K)Q^�k9�B�)�J%]�l�?��r��W
)	��}g��E9�qՔ��E����o�$�*�d'

((���$�&�D_VQ�WP��ؕQG�>⨺^�N��ݧ���|��3P�ȋ��PQ( �q���W0�J
C�������TU�#�Q�n�W/8�p�̢�Np�ZU��Ny����r+��g(uaE��G9�Õs�Ez��.>�Q+��*���wk�>n��c��^��z���bx��k*�0�w���<-<l$l �.%#v�,�*�K�iCh���K�/��b�[��"K��$�s��e�fM���n���Nx��Gn������wl�����#�zD�����{�1��f�܍ݹl�.��pk�ް�L��c������8��ԽѨz�G���|ƌk��۩�a�L��2k�M��M4��	������u��Ꞛ���6<\��Gf8 ��3� ȃa�6�a9���n:�QP��)����on���2gfM�#�nY�)P��Ѻ����(��� Go�p݀Lͤ��8��kv��Qs�D�Y��Uv���n�s������=tB�3����1X��z-��;ú�6�z7">�[���!�#��a�9 #n-{M���[�&�jcJv�Л$뛡v]M�\X������6��eE^r)B�m�I��&w<�%��m�r6n21	�H5�uV[̅rֺ֟=s��k�b��]�0f4.�k���C�cw��~1���7O[��K�;0���+��7�&8�F7v��]��7Yz�A���]�,6��1�..���:�m���n�����h�=#��е��u�����CfH�b[��v����=�"^_�.v�������xַqO%ŨK�i�V�(�bi��\-�(5��n�<�X�8�E����a\�lt��
Q��݄�k�$�5�&����l�-�mtn�ɝ`B;KC�caí��T7N�PGc�u�}LG]���5��=�`�v�6�yp����,� \���ٖ6����,�����N�V�X�/���k��\�B�l�۔��u��gWMy��d��/GX���r��d<'[���o����=�1�$u[l��ɘ�fN�畻4&�[��q�٭;�Sj��J�2���<��X����a)5�)v�OZ��x��Q�^�^��m��q�s�?|q��B�pA�M�@�jT�5����t�����h�`��1 ce0�B!H׷}��Z�,9�0�,� h��*�&��b�D������Ԏ���κ\�c���Yu#�Sv�0h�.m�� ��Q��P���`�X��#L��E㳄�;n^۵��:5:���k�����Ĝx�n4�CV6B"��+KI�vYV��=JGM�L�-�������t&0�&�v�)�SǓ�n���~>{K�����,�>4������%���[6� �3�Pm��:�5c�ik1�+�v�������|�6u�sT�5I�<2��oup�^N_	����c�q�e�A��Hx�T��2�� � �6*w'nI���S�Gs�p��sSG>ћ|O�§��s��>��n&v�=t�����/���o���$�@�A��j�R�<_��G[��O�𜧙�G��:C�;h�p���ک	2Ɲ;K!��u�z����]6M'�kcؤ��O�\n7z�g�'/�<�'P�Dn��T��x$͠�܃�*���T�؊��|���Uӯ�Gc�<���/�§��k��A>�����Ʃ3����2�(!D���NT��J0`D���g�=�����C%vP�;P���l�z����G�q�,`��s4�1�C���x]�K�:��&Ɓ��$��nZoU;85I�-T���Y��̈Ĥ��ߗF�A]�u[6�����wX��n�cr�g��"B���~畻/�$�ᗽ}�
vW�|��	h4�U*�"�'Q��QƵ�Q>��!
���H R ���xv�q9�(ާ�H���7�����*�p ��<	*�+��K�7���C�zA(���2�SB
�=S��oi{��d��/v=S�r��� ��N�L�X��
��1�z�`>�ưz��b5Nf��9�}\�	��ImbD+��Ɏ�LD��B��j�I1��]�8�|���מ�ǌ��E���\���ȜEB���	�ޤU8w���핔��٘����8��LV�'^&n�u:�M3llgZYI�������Y��Tk(���	�A�;N��p�T���L�����=G(t��#oǖ��B��9N��HI�M ݠ������{������n+�Wg5O���7|�pv�A�I�C�E�̇"'r���<AI$��X�kM��N$
�� �Cv��}�����.��X�4v塖�E���(�"G����8���z����)��w��C�[��:�x�������e�^$R��������@z~w魨��_dNg��|A7�;Zuک�5������H�窤�lAk��N�5�L��Y¦}�\�p �RpG��*��Tgϣ�shJ"ӳ�T��CH@�$��(lv�ć~yj,N o��Fj�
Ѣn��C��A��/�9i���=~�|�K|�|��O���4pf��iE��%�Q���FT�-x�ww.�!A�G6t��6�� ��g5H��� �ӫ�����z̏g
th���w�S��?q[V��bݻP�j�
�3�R��O+ͳ���u���{]�eS�g
��ek���ԙ�3��轲O��UaQ��\bPAmb�p�]�)�-8���xǶ|���|+
��K�wpEr�U;�N�Ʃ9
v)�3���5�Q5�9�N&�;w�T���gy�2=|)�W�8#3�u��_P�y��3�XQ��J7}���Ι�Ҁn����Zꇴ�༃K5��o�Xx��z��5/؟v�NG�@�ֳ=U��*&�Cj`�C(��EJ@�������,��vZZ�n �ۇ"�A�ώ����'�g�l���>����t���3h �k�����R����q�1��t�-o�{M�-��4���.x8�bn�� :���bw�-<�����2WhA����Ӛ�¸p��d�����u��R���o��zz!��;y�Kޤ��t������ŧ ���=<�>߶w�����¡s�B��א�z^���])�U6���.��B�*�ñ|����M^~���x|��\��>���+=~|�t�̂Jr7K�T�2J�ӳ��s�� ǜ8y ���XwTI�*�.pA�A�Al�	 ����4�dR����"��ت�q}��9��'��{��Ψ����u�oPpAn�R�0A�|c�8ۿofR	�[�H!��q+��Һ≫:�8�Ef�:�k3�Z}����F�b7VT.7�S�$Ú���<"H|  $��d�CP����
 b��'ϯc�}��:��_^]1,i[�K	c]+��	4��ْ;\M����uK�ϊr�x-�Lq�[�e%˺|�^���tt&.�ڷ�sX���7�&�m������GZ�r��������M��;m,�����&XK��� ۋP
��W�E^nxh{,�j}r�sqEȆ-�{C�Y�)��k��Cܜ7�����AQԄk[�3|�%����ї��ݬB�]��tۭ���&���ɕ%G$�B{��<h|�8 ���+\t¼���;8�����
�_�/�.#E��7��/������������6f@�]�.GW�j�Q��v�U�y _��@����Mp�W|�s��q��T{C�:��]oQ�jKk /��o��	�NA���R!,i/u_lz��uW�k�[��j+"焥�oPpA�R5N�U�[ᣫ�n_ %�s�#�õRg�B��Lw��ٜ�p!�ʂ�:�q�qv��֜�g��K�=����An�!��s�����3����	j���$�w���1v;�x��p�U;�RcB{u{�z�);�n�����
$��nq���;+��V�Њr��9g(��^��N�^XZ�5R�Q�'�N
w����z�.xJ\D��C�����΄1���Ü���U�p�	.3f!DtWd_,ֽ6�&rm�iۣ�Z�4vA��3o��wg/�V�pϲ��)��~�}:e�Ґ�+�����r�(u�cRe��dgt��;����y��#�->��>��!#̀��P	B+@� ����\;U�v���v����~�.��O��D;6(}���&L�S��%
�$o�>�U�]��E�|w���GL��k
���pv�@=s�U�b$�Z� ^���o=��C�/�;S�X��g��'�ǝ����M�xnz��x�!]������q0r�p�ES��R���k�[��ޟH����g�N
�����~��K�'ҝ�f�� ӧT��n�+��ޫe`��%׋�t��Zi��5�V�h6
��v�q���b��BXXz�rs�.R��N3\VX�P&�h��b�8��1ƣ���h#�	�=��ES�T��@�����u�O�F6ҙ�է�E�1�}=Yo<�֠m�sT�ج),�su���L�t;e��Aj�k�ƀ�l˧�0mw_�"���!"���>�׼��5��e�@<
���jb�bSs��`�(��r�YY�n�g9�!|~���W����H��U�
�a�B�H$�4�R �|���=���fs����,�g�9�*N��]�����r`�A�v�C��p���j�5Å]�$��cHf����;���8�8Jػ�X�6Bo+���lD׹;� �u�����VI�M��~����i��F{����w��:7�/j��w�u��0��I���[)4%n5:�CM]��å��a#�~��Ͽ~�	ަ�g.F���+q��Y��o��+���3�&��'�O�=z� "L��m9LQ�N�NA�!	=�V*�x�+�d
���w̗�(�	%�!;ᒄ�Ʋ2�y�V7bjbR�A;i؂.ݜ�媔�]��'w��n_1t�ټ��`A3������ݠ�At�!���"З��N��� 61���8j��26l���ধ3�&�R�¯!���{.�cʼ�e�'�%Oy:Dw�ef0yo�͵���#��(�7����Khߍ��w��2a����j��C���w�S�H� ��b��bH`Sr2@
P�Hu������L��S i3��A���9�C�D��L=�}�j�8�u��k����K��5 ����v,Z�2�l��7����|/�}��?%�>�Y��L�1�`�̽J��[���Z�]���������PO���,���l���cT��Rp3����1�קz��]pp�(>y0�<��C�����d* 8,k�8"�����
o)aL�p�Y6�6���[���ফ3�. �R�s\
�V���ڬ�'�1Z�5y�&����v�C��T�����箲b��Ι�<|+/��d��5`Aj��A�Rgie�n�
��O 'iIN�;y��h1I��ʆ�b3^��+�u�}��j�g��b���C��@v!�ERj�<	&��U�ۉ�5�v�s��}������t��&�8�A���RpA5�+n������2�j�c��7V���Im-r��t�{ÞE�]QD���)l痎����J�9HUg�ɯ�.�Ъ8p�7�����~]���T~��	�ȉ�(�밾��H��Yl#-�e�1n��&���ƛdT���\a�ѓ�"��Z�;uֹ5�WIS�ό5Е���P^.m��r��B���+R�Y�v��k����k�gWZ]qv�5��\T�U�ٔ�틙�q��E���hI�4�	J�bg
Fܐ���4*e�U�]�;v�.��Q/S��W8]<u��y��ƷM�~N����ۨ�`�t�Upk�c�??���#mi��c
�L�-���[��^ݯ>	[�v�8�
�P1Bi�
�j�̂�v�C��p��8�N�
��k/�$=nG�_�����#}�$�3�w��U;9�NCU&�>ݹ|�/Sv��9� �q�T�U����Y\*#���0�9�B26aQ+E�3-p�Y.��T�4 n�SB���p�>����5�D���f�3�9@O�vs����Ʃ8,*�{��Xj���A�v�C�AN�#*ߖ����_2J،I����%���I��X���4y�ڀZ���T��;׭rm�#�s|�t�rk$W�g�����c ���A�5N.�g�$��{��lLpi� #��N�m��I�)��'u�jV̰��	��`̶�^��߿��� ���p�4��z�v�I�j�5�hȴ7:i�pA9ښ�NA7j9��TA�we�.��w��4�)�MfX*��[��,��<�ۅņb���m�7�fާ�7x�q��ɺt7��Eҫ�{��@%�ü~337 0b8�C	�iU)P�B���B�0�_=�w�G?>q�<ϵ����e�%��9���9O5��Ǭb-ݝ�����' �;8�v�Xݧq	s����[S%�'��N�ȩ���+�u��2KPr�R �8I�1�#��u��׻Ha�9�&�U&�Ϻ�n�d�5Y��7*I��AOe�^�Qyňz��8Q)�'�kV��B�n�9�A8�Ĥn��X�P�&�w_u��祗̗8 ��'�
��I��s������m���J��jl�q�����Vx���V[��M�t�!�u	C�^dA�u�֜���Юӱݧ�f�VH�L������D���^�Ǆ(���ES�q�B�)�I�r�L�ޡPr*�;�vɎ���5��Vf�R�qR��k�����p�x���Ln%��ʘ��gm �S��,S�430`?�9\w�)^��:D��������GL̚i��{ ˭���kM�;R�cV���eCF�B����J���D�#�n�4���֫1�8 �3�̚A���[ګs\�;���q�����7�5��:p#����j�7i��m	R��NJ�/w�2�_<�N�咃�����}qSZ����ɕ󔫕$�m�ꬲ��p4� ������۵7J8�:T�Wu�dnh9;Dú-	8�=�{�fd���f�=��v♛�
�u�v�����\ﻝ�<�c��Q��V�nw
�|��n�"vqU���f��Ӯ�w<�l���o<}������Pjv���P_<uո�۫��!,�j�{gU쭣[�u���ѥ��}Pws��96�=��C�+3�0I`�γΦ�\j#��^3À�4ZM���μ��.�껽THc�:���	���I���V���FWs|'7y����>t7qf��v!/^���n��k
�E/+3d�����m]��n�-Ʈ��,ki5Y��`W�C8d�XkK��	������WVN��:xyq��a��yI�3^	M;�w�y�,�8�';ƺ�,�(U��×:��٢o6�_]�G��!�w���/���_h���X=�m��c�o�d��j��zB�G��dϨUi�ESi/�p�/I�]��,�"�S9����8��ؠ��3ua�Yۼ���
4`�7	&����d�Gc���a"��I��f�Mo��ǽ{��~Sv�ܼF�g%L��n<�^j��"H<
�91*��#�D@�ND��BM�g�YوP\����߹�^��^�^^^_G�o���,������\�@I�n��B��G�a^�~��I+��܊v������n��^^^_G�o���(����)P}�'	h�Y�kN�d�W�p�j�QGP��\��T���������������������У�mƪ3Z.t:��0�ǟ�ӟ�/�$P9Ej����/�H�y9z� �7�S��q��x���e��R�c�&S�S
f�<�#�Gt����D�'k�_����"~x��d�좮K�s��\�<R�Q�D�wwy���d����y/>ޘշzf�]D�׏wq�F�C�T�������C��Uȋ��G��;�yAs�о{��FS�tG!%[�|è����~[�ʯ������� )u ����J�)"wp//Ws�kN�Z���+�̩�2�C"0���	PJ   ���v>�w�K/�/��j�y���wby��^!ߗ��=�ZK�c��o1�O�&j�o�?�;�WK����yܵ�K��
HH �l�n�5H80�5S�"��ڰ�l��c���k�ö6ipSU�Η
d*q��.vv1T�2�sº܇�Ɂ���O^�Wl�:�4�3m��f.d�[CNX �Iwu@>�Kh�ZD�R#-Û���"��p�o�W� u�=,�.�:*�s'�b�_!`�8�wxj��Ʃ;A�N�~���n�i��[���lQx�oY\. ��A�d[��CW��C9��gy�8�p��I.7<���*�;*����vy2�z��=�WB�6�py���K�O�8 ���
c%Rql��ol�E.b�Ʌ���7n)��}޼���w�+;K��6�Fou��>�Dy�;��{~ɣ;71������r9����0�L���!=��*�^�+��L8�E�৭�NB�36`�`5
:i��V�B!�;�8ޞϞa�x��<��H>���y���%�R��x��Xø�g�7M�Q�z��.�A�A�`E[��:���X�}^�IR��Ȯ�	��5
t�1n�㇋��ù�����6r@�X쟾oux�;���	�A� m8v"�3�T���*����t��F_�f�P��Mb����NAcT�l�q���1�B�tJ���0���A�p��W�;���;K���܇�W�&p�T{�h�hB،�g�|�T�F28��T��&���=m�����:��3�F=��6�$���U�U!�A�p�2��Uܛw;S(YU��gj�ϓ�6��.���IsA�N�99�r/��fq�Χ-4��0�M�b.�pj��ru�u6����S�U���x]��gi	s��D����I�j��^࠹0�h�;ۈ�^c|b�<��Qv����n"�k#�f��>�t�*6јj�>�o"T�_`Ê��ˀ��bW��P��Hdu+��t�J)ߟ�~�_��m�frYf�b�v�gt�	�b�iS�w9�6)��ݵ�D�:���#T4U%���aC�b�S���k�k�<�r3ji*�v��V�)཮����6t���t�ؼRvzP�u(bű<=����WTiƘr@�3�4�9����L��!�`�=2�����q&�mm���y���x��m�5�X�o�?�O�,�]�7X�lPNp<�Y�-�@��Y�m.���v�y�_��K,��B��U!T(	
;�W���%?~u�I���<^^<&�<�15Ý��T��T�5HA��z^.=/,��v�Ms��w*��ef����t��L���-~�9qiaLc���B�CN�L��p�j�v"�-���t��
���{>}R����8 ��Pr*�;�
�g��r1���<�Q��OW+k�1�R&�;v����^�����&�x��۱1Dg�������|�q���������Eۇ"�*���=�;��Jj��<v].���Iq�I9v�K�j�'���ׄߤm�`<�~������?�\��AF�\ tvM<9�'n(m�4Y$A0D` b��(�ش�nPv �;U =T����t�	��9�BH]g�/��;kPp��؎���ES��T��^jd@'�9�}�iO\�y�'��*qW�vnS��a|�G�g��bR�)a��w�|��n����so���x%]Z�ك��R+Ӣ���f��BA�!��D!�p4jP�MA(PB@-
P��p�_^����3���5�Q�W�ip)qk�[!i5Hdx���^��������-C�k&/v�Ȫp�Zi���Ǫ����{r�`��VrK�oRܛƩ8 �T�c!v��0oX��o��w��~9�F��"*��f���]]O�:��ʰ��)�t�;�J?����[r�	`��eL4MDC�N��<	$kԸ ����ݝ���>�����	����Ε�8���ź�vJ�T'18"fC9�#7��͗���58��۬w�^�W�����A�-X�T��Hyx�2�K�k���VG��l(-�6�bj�gK��`��s��3-��z�����]�pAa9m�p�Eۆɾ�/i_
�]f���8���ep�:���T�����Uk��ZNA�Y���γB������Hx�����]�WG��Q��!.gl�\��[���SI�#�%��O[����S�����'R��7g#���<{σ#ގىSX�Y;���YR3pOrA��x�N�'�Փ�Э���V�&B���;.ћ�L����|F���B
 �����}��=���G�x�b�U�Cz��v��u��Ahg��A�Xk�/I#{��-i7�������j�3u��k����^OLJ�'+z	���b.�/��<�[Y�.�zձ�����~�3|*s��� ׈�p�M;\2n٧��+6fYP���ۓ����c�L�.�4CB#�rp9i���	#���M��xBE�)\A>���2�NE�J�����y�?��z���1��=/��JBH9n���S�`��]�߃����x�&a\�F>���<�m�}�n�˒v/M𩛬ԗRs,P�v�����ώk��`�ּ��M �v�P���x�)�+���*1���������9�B\����|�؊�v"����ND'��Ѹ]�.�� �x���'� �x�SU��t��<\Zm3����g�h������5�,�m7�o� �^Z=�*擟}���r#S���m?��S`�~@�U�l ͤs�x"鳨�y��[:��ֵ�
(�(C�J��h iT(Z��l�>� ����	�A؃T�؊��$|���Ӝ�>�k@�v���'"�����Ip�N;��Ʃ9j�NLB��Ͼ�����%W:�j:���Y�F�k�f�Js&�8��*�[���
��߇�~������ԭ �X�)�ܫή�QW��7HIC��wZ�k�� ���1��v5�g��=:� ��iW\��3�/<L���z�y3o.�>����}5GBK�� ��Bܳ�cT�a��sK�0s��Gx8 � �DӁU�X�N��`'�.zd����v+N�)���1oZ� o8g7i�-v����E􁗈��@��B  ���HKHw����D�W§;|�'C�� )����iϲT�>� z���,wg�;MR�U;;�se�K�ȯ1���=}�;�MGQВ�	�A�۫����ݺ/d7Y��O�]Ħ�S�*�sB����hv�~�f^������]hѵi�5յf��}%=GmM�=S���D��>��3 #��@4�Q5�D�Ou+ZYmI�����n�5�����ŷkOa������ ����,4ZK)+Mn�a�4]�`3:Ql���=�ň�Ulc��1��v���3ԩ�]�&�#�LG$�Қ4�ں��w�W[��E�dJސ99�/n�uٺ��pN6����tکW�z��۹�,�5��qtl�z�:�۹;hŹ��A��&��-�����~��ʹ &���̉�⺞-�ֶ9&1�e�AL�؁�a�~����>��EG�	��r�kx&��f;8��X��R���Iq��r��͸�m����q�˦pj�N���nׁk� ��¢��
;H�p�vn�z�h��U����9�A1ݨ�LG\ܘ��P��N�x�k!v�ݦsv��B��*=ơ��8�r|�����<	p ��@�p�o;��q�p�r{�k��i�10�A�p�]�v�L�U]KT`��U79�. ��NA��Znzc�l5�g�*��!v��9a�k�-{.6���zO\��v���)���뉲��Vv��S@@� ��s�b.ҠIBӴ���O��"�a��X�6�<�x�C���*�8��8o]r[W&0��QIû��"d����-:��7��NEI�xL�yLoO����I5�o���=O��9n���8�ԒJߝ���Х�dw��:�T��ϓ�<�샞R�,�\/���k=w� �Ǉ�����{'س�ץ���Y����%����a�2��/���V���%�`�D ����>"q݌��U���X߲�]NjK�,bӐw���R1(/]m�2�j�A(��Z������6��e�u����u���Vn����UA��;9�NBآ��Sf�&q�vi���I�tL��Lo��WI���	��q �zܧV�+�k9 �8v"����7n�7dǖ�;��z�k�W5��l�땊,we=]NjK�E�,󳚤�ƩL��-���YQ1ԅ�:���.���Լ��[�K�^��ɠ�f��B�K�z��ȇ�B��5��H
�+��7�.��3Y�AH<�M��vk�3��;]hV��S�F�;v��;�Hks܎q�;����rp ά���)��T��:����J9n�!O�X�F��+3B���3�
�<EU�hv��=����T��H�+r~5�wng�'�ĝ/yy��*M��ե`S9|���7�����d�/.���ON�#��5��'��a��%Co>w,Q��)��s�_�' �;;��ɮ�c[8Ġ�iԕ�_g���/�AN�f�7��@�ɬ� ��� ��U}:���']���vq�H/��@��lP�_��HB�@Q�ߩ=��Ͻ�*�O�9�^�F�7h9H�����n��sb�
Tӥ����(:0tn��0��Lkpuk��3S3f����??-
~��DÁ�A�5�U��T������:��Q��jW�2=�Y�W��gSO&�;I�(�����Z��@��}���`�&n�<��z�;��c�ɬ� �	�A�9ÀEW�z�zw<�2�`a��u8 ��N"���� *�ǻ��/WM�O����Ul� ɇ1��9�A�-T☃^q�/C�p�#s�ab<3�y��M5�5�~�Z�\�ߪ3@�w���o$�����I�u:f��q��w�ɑ�PҢը��ܫ|7:�i�k�qԢWW��t).�/��5�9�:�q�������2�� E�!�b�p��˹<&4�#T�A�9,AN�!���Ж�qgo~긽%{+7H)- �s�Y
N�ES�H|\��L�OR�.y:*!DBP�e�9����6w�i��].�ڻK�O^��}�/�ϧ��w�&���)3����^U]瘌�]���Փ=9:�z�ȷ��AT�Ȋwj���gO��>\��!Zgb�V;?L�[����Tg$���-3��gcT�����#�֜hd2�@>�p _����U8����5޾��xyþMUV���+�Y�B\౻A�9��U����NR��d�D�������g3I�mJ��<�et��.�A T��eǲ����n�x��i��
� U �|Ʃ ��}�x�i��^��3�l��r���Tg$���E�#�3�4��R,'0-���y;�L�����Y�+8��P�cۖ�&�J;w��u�Fe�h'P�e��z�=Os�Q����i��ݧ%X4Y�r��w��+6�X/N�bIF7��(�ArǓ�ݜ.&����v��x/����	-J�/��Y]k0r,M����	5�(��-�V��˖x
/g��t�r�_nv�˔x��n�<��(�ܮ���z��<�e�뻈uώ�j�5����6�n��ͩz����K2�l�w��	�l�~��]��Ay��I :2�n�gm��j���^KRA*�ۡ�4ӵ���Mb��4C�o�o�~�Q��K�[��H;���e�f�p:����d��V�c�\��nf�G`ͫy�i�=v�a��h�j��YMT�����K8��f�ǘ��k|G`�7IG������+�l�<�Q��|+�«:���^�H��U�7J�Z��7���t�Gf���u���fb�}I���{��Yf����Ŷ�7X8on��tu^�M[�k{��8�ŵ�I���繒�Ny�uq�ͣ��E��vB��p�%��J8��,vpڭ������Ļ+���چ�����]�gn���[�];6�*Z�fkH���נqwMujɴ��פrc;�˵��a�k�˴Z�L��7	�Ѻ\�[qCK�֩E˃aCf�ճ�v�|�D������oN�4;:�bQ���5�K�N�C�nKc;���G�6F_�b��O�	���������o��	�\/�,�����u>����|xX��J����q���!�5j�vp�H�W �
�"=��2���o��J�W�t��f��N��8�я�����O,�����CSy��m�mf�9i���!�HEr~��<���6�r+Aw�8�!�Y$���w����������������φ���5���</B">�M2�����>	��{�x�s���&����ח�N�Y����_^^�^^]�bĄ(�P8��y��iv:9x����$�A�%򰪼�FT��"�_9,�O7S��U��uP��YM����qz'/l/;���>���9�����~�r)�?x,�I���^y99�3J����z�g���Q7!���(�� ��*�tvTA|�^����y���.�H*��N�����;�Z\T�Ⱦ�W�ӻ�����_!d9��U�J���,��y}ܜ��W<�̃���K{��J�D>}ם����'t�N��
N}�}����˅ܛ�AQ~E�rw{��!2�v��)���l�xK<K��[�Oq�E�3g�>!-�[�a����l�a5m�3D[��W1ԅv&i�8d�b��u��;����ܦ�{<��X�:(	�KP7aB)���t-�P�XƷqmۖU9cx�%����N��ˢ���"W=Ym%�8�k��ͼQ�C����a�c���V7S����n`%���zNI�ዮV��B�wd�jx�e��]�dku��6�P(��8��\tؘFQ�ۘur�N�B���;F�����
m
�z}�lU��ɭZ�B��4��,�@.]qB�42c!H̨�)���as��R�lI��qJ�#ecDk��4��M�=%m�H�CV6��`���СDPM��e��/���y�8�v�c���<kW%�Sc<�x�!�uI]��;+�9��.�X�wd3^�Y\f�"B56JE�\��=��4sh*#����"Q�{]<��Cqťɸ��Yt�nxN ����ny���jX2���A-#��.��q
,��v��˫�l�XMې.ݲf*����l�U��A�ꛂ�l!��%�K��q������ &y}����6*L6�q@nl�A�{>��:�/L��@��tU�!A-�EFK���8�n����}eێ�'�=xo<ے�����RݼE�{o����ε�#���t�ⱀ�J��	;vk�\��s"m���<qC��[8��������:u�s���1:���7���o̓^�=���q]�y.u4h��r�n�g�^9�k�H��X0jĂk�6�e�$l�rl��W��87M�j�A�˪�G�i��$�7���8���x8ysۓ��̲#�N�\u�Cƹj�G�ڼw+�崦�h�X�/�E���:{b�]ձa�s���t[��[�"�{]g"�n��Z9�\�t����?=�=���.�������F�]���i��O|<�hl�G�`��o����KP�|4���Xd&��������6y�$�k�[��O�ߚ�2��GR|U�٫�.	u]-���ځ���U�
p�-�c��½�<l��m<X�C[�>�*����B�*�k!@�����ee�̈r�q�nA;`���pn�ζ�I\&��J���B�����j۔|*�Tsu����G��itN� �A�ݸ�ҥѣ�mOS� ��\ܻ��6�5���%Mt�́�b9&�.��Fl�0��P�����O�6th�搵��FcL����5�K�8���MS'¨ �py_���6�C[<��R�ũ��ޫ{З��t��s���=y���W��� θ�#6]1
��������X�b�GS��C�IT��XĦp{��T�zه|��=�����g�;Ec�5H_��J����`#�Ñ��Ic���LR�ERj����Q�=��]�S�nw/��.8�]=b�����I5I���*b;��1��0t��Prˇc���LR�9�7z����gi	s�V8�!��A*�������`�8��2�9T��`PͿX���F�Z��.>��{rV=dü�Q���������A�-T�7�J1�hݬ�0pnmmE&e��	�A�%y�u��J+�!�3vɜ�J��;�B� ��S�	�Aæ�@"�݌Ӊ>��W�z�T�_�3R\DYj{�(TA�vp5�Ʋ	�bl��Z�S�lO��R�ݻ���u
�P�Õҫ�'�TN��;0��nY��d�P_@Q�-�s�.�cά+��:m�3�G�� 9�Ƙ�wO�[��1X$0� �İ�X5(9uÎ}��ߪ޻Ο/;HK���A�-|�Z[�*"iߞ�����滆k� �N]��p*�����7���n˼ܯ<�Q�A�����! ��� ��*��c[!���~�X��A���tw\SC"�mõ�m�ܘ��S�~��m�q����,�f�;t�`G^�\Zm'�I�T�Aԃ�MRƩ=k�q\=b���{�v��3t���n��y�N1I�k;!�u�fLM]6G���!�ú�
!�C�91�$t�]�F7�����@`���^����x~���F���ɪNXu4��j]�/N��<\�L<�귢��A�Ӿ��0�p�n�r�p�B���b-8ɺ�=��>�`x�A��vv���^��=���M�����)z�M�a�X ���K��y��C��������](>��%��xzr8��b�I`���{Q���C��ay���`�@ȳ�т^L>��ۼ�Y�h�]+�.�h;�ί��5^�.8�����?J!� �	�W��/�z����� ��j�pA�T��U;m;=��F϶�.�ڔ�W���9&��vsx��I�t�����\A���Z|��#af��5�z�mn�pES�� ��8t*�4#�T݂Nӷl��7�˛�ԗ1������!LA��6�r���j��j�Ҳ��%KVɖ��4����b��aڧh]	w����Z,n�hx� �T��̞�޵u��_i	s�q=s��qjq�N8�J���T��Rk�1'�XJ�����Q�x*����̜_O�y��My8�+U!�	�����NX�z� �RH>l�DR�p�S��;�z��)`v�������}�~��Iq�c� �7������Fӳ�� ��[5�2�l!�0!�b�C�ÊY���j��w�2�HK��Z�\f>���|ff��>��U�������B+s�����vK"���ߕD��@��E��?+V�nwP�Y%�B�XaJP�4|O�$2C!�>����tx�Z�Cď�Wi�ݧAk�b*��C���B��$�'���Qs�����Iw�@�Y� @1h8"�
�׶36w<MX�8�|��[�[�7(��<�����:��������F�CXאp|��DS�T�;o��#�zf}�uq���q�)Z=\��Y`�TN߭�T�z�O�6n�T=!��@�Y�:w&[(@.�������\P���!.pMZXE�W�x�w�//0�ܓ=�$����S��Z�����T���2>�^��O��5��	.`A�β��yf���F��1�zL{�n������Ū��g����{�>�ʸ�Ip�A1X��e�/M�N��@�ӐXͧ�]�b7h9k�a��p�rs��S�8Ē[mé���W;�2�HI��1�L��Fc�j������|�����D_��Z�z;�pu6���4EXm�g�#O��Y_�T��,�os�S��;d�&�;8Qv�do��u��{�&��U�O�C2�H:�?R����'��6���f�S1�,��	a�b׀��͗G�:S�Ćr4��S���ܱ�ى���vz�el�7^�׸+f֮ҎNP{#u�zy��뵜�'��G�1AY5�nw�H�1��R� �!f6�z��5��36hD�/ks3G;8>������i����<U�Z;=&q�qł-�زhͨC�/4a�un/�������K��|�x6����_ޭ�an���u	b�����!�v
kY��D;�C�^e�y�o�̤�X���Kf�@7i؂nӌ��F�f�Y]�K��.f�&#��L<��yÃ���I"�ÂMS��9�@F��Z�{ ��|�fk��s����*�5%��jp�f��a��q��HZ7�Q��������"��d�A�5N%����T>�5�����٩��c�f�pI5��X�˳�fSBӾ���a��g�8b�;g�������+��Ip-�A�o���O���=}�ϥ"yb.�:b��e�d]�@�E����#�n�6���G��>��������*�5$�c��qi`�������5��'��
H�Q32�����/)+�>�����n��2�m�߱�=�^���v)��Ѣ��p��k;G]D���}�%��ss���s0(�pAژĘ�gcJ��vWj,n�h�#/Q�rv���eVɪ���'e�̱qˢ����0�|�&��Q͛ݐꫂbOj�r�U��%�T���?�<�����@���n�/9�F�y�\s�}���L>��WA�.�؂�|��k9�B�oyE�&=c;��I~ci spFq��]<7�~��`|or�s�Mt繚�����v#53����j�U/ E�����F-��2]-P���Z��X.�Jέ�U6qe��%ăV��2s�dQ	[��!�C���;m��j��A�N5N<�R}���k�r^��s����WA���Bd�|��[�.
i.��Hi~\�g����ǩ�hQ|zv�c3qY�]�C���h{q��0kdn\�j����^�:�D��R��^��2�B�k����Bc3��z�VJ�O��n3�C���g}�s5^���2��ާ ��MT��*���!)���TqU��#ԃ�Ek����U;)e���8,f�rW8v,*�ۘ�	����C1���%"�uH>(t��n�j��MR���<s��.�9�[�#ʮ�C�$"Ɲ�4�s�r����f�x@���^q����'uu�32���W8�&]��w�\A�g��vr�˚��� �	�!�#g:y9�ж���:_,P;H8$� �T��2P�7.�i{ F^+�S�EC�A�8pI�L�Nϓ^��d��VM�u���#ܜp^����,5k;��K ��b.�H7h;n�9�C��/4�6����5[�:�$vR��<aӀH3h;XW8r*�bU8r��a+_U�l�C��x���	�N��t
u�ƀU��V0b7v��|�h����޲ߞ	�����j����O=�T���Nr����
Y�8��u��63X)�禕 KU �Y
N��T��/��'��u�{���a�;�������ޘ�ɸ�Ip ��>$�ĸ�	At;9�Q>�>]�v�eJƱH ������BR`��=UEš.����k�e=Hܪ|� �p3h;k�9N��;� ��W��!�N.��;�AN�Ы�A7i�v��s~��bߠ�IsX� 5��z�:|��w�Zr9�Q��,�
qvm�9Nbe������N������g��q�����U�e�9��B��b���X�87�CCr�Y�;u!Du�c�Zp౻A����o�+ة�������#f:s��.L����#5���N�T��e�~܇+@���M(�6;`��]�n�Þ;�W����H1�õN�ie�z�w�aY�ڄo�5� �8q��[�z��_Mc����z�"#q�yÚ+%� K��Ů�9�&��A�8#ry��~�;�����v7��6����.����� ����x�/%o�������K�wpA� U8pES� ��g�[@��陯T�߄t��z�;���	�y@ �y�U' �"�U/1S�B�J.�Iΐ���C��0A�1w]����X���/s�bӒD7+]���*�gI�p�k9x��)�УG֜�o��j�D�I����\�<�tuޅ=�ߠ�Iq��A��L`H;j�r��~�����DwoNAJ��3l����^(��$V����Ŭ��K�OH�"���9{uޗ������$�+�����U��`��%	�M\�։�? W�M4�Y��L7q�娢�vMÒ6y�k05ƀ�u�����6n
@Y�qu����qHh��CBc�[+G���Cx�\θ:��&=us�w���f����a�q��MX�+���R�ˆ��I��P����'��#��eSr�uK��[M{:2��sm�0p^��L�60����1��W�I�]4�cҗ��U�d���X~������q.V�@��n��5��k�4%m6�7�~�Q��C���*���DS��r骝��鎜��rK�>�iy��1��NA�vsv�MRvvA��A � �F��P�	��b�3�8<ǵ����S�^ެ~�<��m0�BO8r+ַ�`}���x�9�P�B#�.����`������Y�e�	Y\*��Ц���	.`A'iñ-Ú�� �c��#Ľ��N����;Ƀ�+�j��;՗Q��1Ӟ��vw~ �{ɮmP���Ӳ��s�N�r��Rp	L��1��Q"��t�
c_eNS��w)]W#���H>�pA�A��S�,`���4Ӵ-�lb���39�R�ͧ	E4'Y���&��TK��@�v9��u�Mt65�~~�ߵr�-t�����j��d7i��bi߽
p�9�R�lQ���}�B�U�pr|Ʃ���و8�};U�M٦)��Yb�	�]�3gnfّ��K���c2�wp�b��r���݅����Tu4�4�_f|G~��/B��L7Fed�]�����Z�y�O���2C�/�^;;w˘�7뿽�=��Vz�9%�{���u3��W�f��У�qG���\繞؋��J� ���.�I"��`�H�ؓ�D?Mt=z���\���� ���� ��rH�8v�L��'V�uw�t���\�g>@�v��Gm	J��O��<
\A�ZG�F��R˭N]�ބ$��2P��rN��XҵNI�튇m�ܚ]*c�Պ�5$�{��u��R�<�	�K��n�'l���ǥ�a:�$���s.�\�<$�e:KA�	qi���vs|��~�?��;Z��j���H�q��}����#^��H>����9��?&��~hI�!�����'b	�@97Ϯl�<�hx_y�Oc��ݡ%m����~s̗�R1�J�X�"������;b��̥�g�� �NFbE��	h�b~\_鵺�ݵ0���{7�%1SX)�M;��rl���S�_�����㔶�����me;��u�ǰ�����]��W\�m��2V�V�n��tUΝ�¸^�[.�@KR�U�p����v&��;�u��t���x=x����[5�ۺ��4�y3���v���n��m��l �@���Jw�`-;�Wxh����5c��Qv��*c}D�M���=�SU/�n�kw3*���l�����ѸxX��T'm�3r�J���n���ыm�"�r	̳!�5��;Ժ�h�7Us5�.��$9M��n�o�rf��9vt4y��;6�e���{�L�OR�i�7tLՙ�;�yI�I��,T*��Î�[z�V�l��]�t�ow]<�v��.����t覑��.�<�<�MKbneq��(�#�6�d��(�bu����BNQ�p7,Z�/6�
�m�W�n�* p/*��7��&�T�;m�wA�s㦰���S"�p�i�����T�a���v��V;$��'�Y3\2�-6��rj�(r=of���<�ݵ�WWp�B����ը�ʊ�Iuf��u�WW��کmE%Zu��㵠m��M:3iأ5��j�����p��];A�+�oP'�XiwvA0"��L����2��|o9P��㫬yx���o]u�X��K�hhM+���@L�]0>Y�m�W:��z�cf�\1f������W�{(�c��d|�+�X��rU�z���cĆ�f��j�����;\�����u��b	Wvn� )/�J?��AX�r��U�+HWG�@b���+��Vt����nﯜ|'�8��ߕ�2�9^���y����kt����On��^^^�^_G��}�+_���c�.Q?�|O�O9�z;�e<�����s+����=�t��/On��^^^�^_G������~��}���t��iۦ'�{�AG�d>W"��wMF�Y��ׇ�O�<==�{|}yyx{yy����>�8'ߙ,"s�d*��T}I�{�`b�r��|��"�>{ǆT/\��LĴH��Qy�f�����-v�,��^�����1p����r~�;ͅ�:G�G�"����-�|#�`Dɼے#~���ȸU���t���������y���I֔P��}y�/^�S�K�4�Ш*��u��p�]iEW����~RnQ�Z�w�R֘�{�8��廷�¨�p�1oQ�p���#���zL�r�;���(TQ;u�[��㒅�U}\������VQ^�����TS,%�����t��H%��!�!�i,���Vn8����{9%�0�yӱS,���Nl��8��v5O�z&� w�>^��Ha���^"�9#z2�W	����q��)w�D�r${&��l=�/p4ZcG=n�X� ���Cb�b,�v9���+<���oZ���Tf���׌���;�d�9bA�A�#-ÑT��qC���T�=/)��_��~�itj�Ԙ����6t�6�;bwV9����j�rp�C��M$@� �=F�`�r�;T��h��wF�T�g�{9%�#�Fu^������= A�̄0>��A5��Y0��d��!�*f�rwgg�cG�e�q{w˄�]qz��c�rH2h� ��������̺o62��L����4C���R�1��Û1~�2�0L���u��v��	 �;�>b��8~d.�������v٪��-ܒN�gjTC�޻�gj}�Ӕ��Ip�S��Ǔ��_{`t\+����ୈqr���/���+�F��nR��1��8�Hd1&L/���j-����z��aQe^n����[��mV��;�A��A jd�Ʒ�)���A��d(�@���U8r���k�=f8q�y��3]\U\g1�8&M�XU;;TA��F�Lx���$�D:W��5��c]��v=��l�̴Z�L�U���=��m-b�lys1Fm3ڲݧ4��;E�i�Qbd�w:\\|>�K_�!!D�w$�˂ֻ�d.��ϋG���μ,���u���c+x�/}^�t俳�M�.�1iƩ{ާ����j�#�M��Cƍ �8��:��{\�{:�Uɚ�Ԫ�9��d�pD��U;��KR��02�P�Wg�;�=�BVC�;�R�����'���Њ��l
�n#R�|�Ψ8p�BK�<*S�&�1UN(��xܱ�Pi�59�&��T��G{%����	�N��1ij��k7�G��~�q�{:�o��o�3����������9�xY�W�¬ɛdFz�K���#���2&A3�
aL(`�����޺,��ك�rGm5F�yR٬m�P�
B,�X���ӞF۴b��v����|W=�3m�z�>�tn)H����W�k�!�;+�9�7n9���i/A��.��{v&H�2�t�V"bE��m�9�i.����vI�A�M�X�n�ǅ�8�X��Cb|�r����=�"�!�J6XCW]6�p ���ٴ�J�L������պ��S8-̩V�Bkl��a����¶;wI������F�I��n��`��y��ws��������>��J�3��	��m����Q�j�9�����Wr��nS��5.&�M ߓ��U���
Ux̞��KG:wv�pX���Y��C�7.��5���+�A'M �8r*��E*"=���e_�}�g�=���;����Ư�^ �T���r��U�3p0�m�:%��B.Aav�Onz��ƺ�+��c<2h���yny�����=hx�br��,Sw�"M�z��;uji������I�S�5b���"rw�.�9�����"�>��;ʈ~rkZ��Q)�h@��RF-.m�A8�+�!�Ei��v!!�3̒H%�t�qll�h�;"�ݨ��6��ej�F?��C
��{P<��9�Y�RpA��S�K�j�R�F{�I��<��(/�Zx8 �T��m�V��4D{!#�#Ru��M�����������,ns�ݽ�Y�s�Ql
�x�O�W�'���F@�)�Q�����8f����g���urWq�ܩ8&M1'\8"+=�Qw���ysVC��j�wS�m9ż�Y��u�x��"i̇��P�'"����#��A�9i�� ��Hn��ԍ�5�됣0�r뇏3�4 ���	"�q�6���j�g$�A�N�F�HQϳձ7�G��NA3i1k�!�nЀA�p�͛!^LE���X,��zct�O���[�f�2�p�z(��X�vv-J�{{g���l��J�!�J!�0��.S�������ǧLn��eQ�gh�mv���ϊ�~�����R�o/_E��;�	��N=��.�$OF�M���C�|tt1蕨y�=�����=U ")ݨ�pG������m�K���d8�ʛ��Z�!g��\Ēv��F--T���ѱ�	�#N��C�B�� CT���s#:B�z(�}��љ7���|/��8s����Q#�W�bUח����I��&�*��osÀ���������kXB��.��z�5��:�]a�1|��C10 %�}C�٩����s�8,h�g�N�*~�*���o��o�q���|��Yf�K�;���{�Ѽ�pEpC`�\;� ��x���烒p���o�yd);:b�4h�j�	5�&qWn��ڬ�9]Ӑ����C��rK����-!�Rr3I��:��|}�������G[��)+�l��Ic&�\Dzh�*�.��j��N�$�&�@?k��p*�8�˓{�S'���K��_G�_��)�k���D�aV�ZZ��ZC��ND��>|�9[�1�jr	�Q��*
z�<��V�W2��6Ա�E���/V�yj�zc �wg��T���vv7�!�k�N��ɮ�쬇{�vg�[��	�NA�vpRpE2	Rr*��z�{��f13H9�5H@�̓��Sޕ����g��`j�r1�ׁ$-��;g���k"��8q	lT�[9�XY0e��Yʯ�m�����ϊt���-�z�0D9B���7�C��Y�B�����d5!�(B��{�ƶ2���f�:ev�BeT��T���%1>���Xs��\��,B{�9��?��k�E��B�H[؜��5%�S�ߟi�]G�i4��-��0�l!<V�^���;�g�y��u���E�/�oS�"�"�ñ�vx�w=�|��=�\��;ʖTq�q��r��8 �󁔼U$�U&�ÃR7=x/E�Y���� �#9��eɾ鮯K���sTǍ��Â.�Y~wژ3=�͞���,jq��Zm9��c*��8�)P7�𡿱�Vn����$��k���8sF��@3H=a$�W���Ny<��N�L��wƍtwv�(|�\ 妋��/�3�Q�'�_`��nך�o(&�@���8sF�DynxFПk����u�z}����eҢ�ءX�Ȼw�!b�#�/�J��{L��F�篝\آ;�=������e����յj�#��"Hw�F�B�raɺ/���t+^���o�e�3��.�[�? >C Cγ��g��=�z�4"ͩ��-6�y1m��+T]�������n�Z�]�ӦMqu���#t�����6�WN������af���ܒЭ�"�X����N�7;N�7s��͟�g<�4�p	�gf���-ɫ���C�m���qJe�1۬�`��fǰX���=�����¼9Y��sأO�4nܩ�0�BuMnL�7�Wm�X���[����٥�;v�aI�om.�](�΃��W)n*�b�=��O�{z,�}�����~ӈ��!=Ȟ0vt��t��1X���p�p�pER�0E;�C�k��m�;��d���ΖK��v��6Ё�뺇Gw�	��f7;�2�N�j�W�������#�1IHyԒJW��I�AȫA�I�"��i��F��:��U�����-��X����:��N�� U �d��� |��ڮ����ؔ�O��A���!��W����`�Ȟ2\���Y�/-F�=1)t`�2t�mõ�p�f��
,�r���T<F�R�h��͘u�z�>{5%��rӦAb�<Ъ��LR����������{�=��	J�/��-�Kn<'c�>Kfu�`�r�����c�H$��i���A�"�ÃF��j�;̹7��>������8���r���EɁ�������p��$-Y� ݧ�m���NB���nm,Aw�U���sw(����da6Ƀ+o��,��dt����̾d��wRܜ9�v�۾�^eu��(dY��� ��u9�'�ޡb܎���pEpr�r:�Q�/s�����.��{�>���c'ER�^b"�fr�x9�[�uʮ�d{<�sɰ�ҩӂ	�N��Y�Rd,��B�X9'��;F�cǋ�S��˓y�s��|�3��cFHLb�T��d;�w�=�c�H�d>2�P�1F�9Ր��*s'�ȶ>�Y=#���Q��]�ː�-Ԛ� ��7��])�/e	C�.;�kB���T��è�)h�\�fKKXmbn|����O�l��L���v��4��,)QѻWP�V��>��rK��1��6aAx�cX�r�i�gJA(rWgP|d(w�^�٨�+�>#�Z1�.Fڣ�sk;�s=z�x?�� c��*G���آ��BnPC�G��0U'"��3��Y�{��T�0��HC�ӵ��Z�J��ΰ.��[��k�*���������o�̵j��"=a�YtRҫ�	dV�a����o����ﾡ��Q��G６�W�D�=��1NѧG�U X�􄫷�*�n#��t�w&r�l�������݄����K� �ZpF��]ߨa�Yyf�
���Õ�� 􆐡%�����ksk�����흜[����y�g��l�pl��m�'�l��4����7��X���홈ɣU��in���e��j�ȏ�!J�.�5�qa�v �!�Rb�H&��g��X�(��=�K�+�z��m�ϙ�ƫ<�Ո ��ut*C� ��;2u헮j�1���J�Gu]��݇�|�w�n)���).�BRy�{�s���1d�r�k(9�E������v�.�Q[��kYy�{�늜�w��x;Q�rs�b*�؊TZ�
KD�:q<&4�˘���|o�� ��l�X�>1���<�Qr�!��5�Ԝ^��1��n�f���²���.X�K��門mf�qTӍ��̡�&ާ5lŐ1G$0`�ǋ�v�8d*�8&1B�Â*��ԺtG��"^�w�3gû�#�[��1�Jv �\Z�7��,�ٗ�z��	}�p�8��%$�����c���!�3��c��)\k;�d��� �6���oZ�;4Y�T��Y����wy�g�����~ʸ8D��!d����Yj��J^!�%�"�w�4�'o��\���{�wy-�8�R4h���q����%�և��,�N��p�F�����h�b���U�����S���jwn`s��s!n�k�Y�$�Ӿ���>�l�v�u����z�S��X�8,d���/w����V�7Z�'a�{�$vr(�R��������{�^���{�f�-W a��p�n�cF��S����#���<��c��Z2�б:��ʎ�t�Ut;{�6���ۇP����Ff��n.[gF^^H��:���T�h�I��f^<4�W
yOӊ*7�S�tv�n�q�:��S.���/�+o*�m���WJ��4��\�x ѫ��9St�c+�z�J�ޚ�@rDY����Mf��A��x%Z�Pb��ԧ����B�c��V�E��ӵDخ�ZI����wֱ�E����r�(˭�u�C��ͬ�y�jи)^��ī������6�T��٫����ǽ;z�h�/�V��q��/ y����ڼ�欏ƇQٕc{������V��v�E�¸��HTe,�>e��аo[:���S[w���ĺ)���TƳ��ͣ'��Օc;=
�=隹�)��ݣa�F�w�$�y���o��ބ������0�վ�@9a#�e�ǣq^����7+�8���V�2�g3ݫFU���Z��H���_vn.,�|��WR=�����%vu����-9SoV3`]ws^/m�Z�fX���^N��iqԑ#�t�]Vځb9�nhǮ&��y�}�;[��w1\� Φ �ϖݛ�yؔ�'7���ǘ�1�=`�/^���uʮ�P�c�Itfe#kEJ6p�>��ǲ�W[��o�F;6܌Y;�DΞgp\�Q�4l����f���tmXqwz�J,Z���sHD�v�pJ5�T(�5I��C��&5��`c �:�C
W/��?R��to�;5�f�ՙ#j�k��޲F�^%w����ślm
�@3@Wee�d�:{3�ǽ����QTz@���� tc�vcF#�9v�N��O//on>>������������|i��������?�C�i����l��7ȳ�G�	qoDd�y!$�"��S&M��Z����z}}]>�����DjmZK*k켊���Iʫ�)}�sw'e:)'/D���U|�3׷N��y{z|q����ǧo��uw_hDW{�{�utZe�(��Y�Wf5T%,/u;�Y��Ӿ=�,4%���+�t��
 �@�q��>�9s���ױ�<z���9��s""uq�*�"
Qoq������Ƞ���{���w|�Qm�k�	k=9��!,띡.�l+��$�r"O���%D�9�h����D�V�p�0��|�Y�L�Vr�|���8�t��p�QBt;�w��+�YAQW*�
���9�=�$�ΐE�Ujˑ˲�QE�n�h]	-<��.C�*��=&z]1*Ԩ�i臐�t�@����-���A�I����Tr;��%�"��)��?x��w2痗��/�)��4ub�&�0h�����rt�����:ҊY��m�hnm�=v�-��=t�K��5�/l�]�1�ԏ�������m,p��qʡcg����Ŭ��2����n��n�竵̦9:��m)r�Il]��n����������c`�:P��/i� �I����|��� �Z�ҝ�y�+�W�n.��A�v��#���Y�lc�CT6�0�Eࠒ̝��.��6��`]CZ����&��E���7���X�7���D�i�/&�Y"��{�j�W���bWe��r�xÀ7XN�M���;���ݮ���N�<��.'�j�����k�kY��-Q�i���қ�&ƌXF�	n:����+�˟yi�[|�%���î&�P��*�r�Q-�E�m���{0�ZET�Us(k�z�&�4�cp�9����2<a���㓧/�8���u�GB0��.�I®�j,X���8��pI-e��5.��Mv��]��t���s[�lfx+�V;Nv +\���n�ta��Ӝ2�8�sxG:��d��'ct�ūuvo 8��K)l�b��:��M�����W7n��L�<��"���Ýa��3�D5�F�3���͔��SqF�q���c�-�v9s0�A	5�l�3Vx����mp@�wj������o4��6ص�a�T��b�L�Yx���K�K�����R3D&�GLk��:Y���;Wh���
�u�}Z���J��[t�wu�6u�e�EU��r8�
ѻT\-xt�
W�t0nښjY`��B��ڽ��!�]=�03]n;er�{�e�ݭq��uun�t�۞�t��N�⸹�Y:CY�G�̦��dͭa^��Ʉֱ�S�Vh��y���\U�v,����\��b��Og��i���Ֆ\�i�1`&��+�<h���x���+����d2i�``��_Z�b�����mr͞��ػS`G�D�P�\��fsv�(�B�*.fB��^8�/O*m�ZpI�r{>#]��I���H����SSF�5�y��R`��Г��[���zNx���v�k+Za��Wb/<�U{.7s�4x��#�*�P���qUf���wc�L�4��v��=\�C�p6��D�a����y�YC�����nc��6��m%��s�5㗊N݅e�9.��u���i�/����];5W���D<^��ݏ��gRM���#��Y�$^�M��1F�	�Aȼ�̦��p�-Q���]6���_����s���v �s�,*�z�_y(�1��9�i$���+�Eū!�̪�C�ٝ|�x~��Z��=^�w��C�́q�P�v8v"�h�$��Ɩ���������z���lA�q-k�b	�</�WC�<y����:��X%9�����W�9�L�8�N����L��Aݐ�MF�?*��94�����9���}�랺Wu��x��v ��p*��F��~Ǎ���T�12�O���Ax*!D�I�/i�.�l�����x�R��������|?e�]�v ڲ%�N�b�;^Κ��=~�6�ǃ��vB�'FA�[� j��;� �O,`1�������{��߆R�tE,ó�;��Y�.�VX��{�a�oS��@���W�].���d��R�=s��UYw_��Rf���.�܅����W\v$�����u%ŲS��v��J�?���pb��+1� �$���7��]��� �ER�M�"�:nzz+��uU��@����A�q�*�ih�g��T��F��RH��J�r���	�w ���<jϐ��xZ��NZB�rai���h�҃�@�qb���Hj�Q2e_�H�Z1/�~�������5�Xv$������ �'b�vq,�&��
�J�s�{�h9��������"֡�a�ն��Z�G'Z,�/���I��1�%7K�ub�t���h@$ݡ�qݞ���]Ϯk5���~�����H��BĲ	�\;��ؼ�ߛZ@U�-��[�э`�' �ܞ�GU�!��k�x:\a�c����bZ�E��^���a�;�$����i�i�o1Q��E~k�ߏ�#��|�?	A{���n�;k�&Y�:gf��¯gl��uҺ�궻3��=J�47q 2<�bȰ�ƽ:h�Ѧ�QK�0�x���%umbxͤ��'%;Z����NU+b.�4�qX��ގ��4t�����C��{=�����k�v�A����z�-D o�;�m�g�UJ�y8�g\�R��z���6�ȴ��m��G��etW2��Lt��p��]������'b��:�]��p�:e��!kf�wgb��l���*�dl:�&����7�Q�7u�^J�����n�S g'��N��M9ЛL�&y8 ��^b(Ԅ1H9�&=+Q��L"	��{;}���e��u��x;x��W8r*���<�wlD�ง��v-T��4C�j��Z�H���Ui���I����lW0@�������P��b+�q	�.�����|�Fc�eQ�W<u䮝�O��,FR�DLw.��_З�Ԅ�Y����c�Б�Ո�w��X����J���d�R�ڦ��r����iP���a��֩p#72�MÀ�,��8�v�m��
�)2
�ڍݭ�HO�X���3ӻ���fD]VsI� |h�\��N�R�+��Ϗߓ�ټ{�����zܒ��][4yx]55��S��x,�ؖi�M�z�V[��?:��ϣeU�|��i)8Ν5d�lNu�tW5��T)ٰ�eB1L9�?��R������ÑV��5H�*pD������v�ʹ��t�xͤ��rS�C_;85J^΋���`�^���@�pb�B�Ú���U�^%��N���G�'32�9���>�Z���n�	"���b�&ju�w�c�D�kU�d�p"�x�'��VHى��=�1���0�e�0spA�,\Mv���ÑU9Sr3�����٩�3;���%�<1�-�t�v�>s��T��R�3��_��p^��ۃKc��o{.���%��7F*h�K��ٰVu��S.n�ʾ����Nd;wu����/y-eڈ�w�0��Or��ۖ�>SZ�t��zꃝ�P=w�C�$�<�s
FݒK��,�:a�K���X����5��ה
���q�i�Wmn�F���tJ���,�A�Yq ]m&�ŏ5��if6��:8�WX�ִ��\��ܘ.Ԙ�����Hx�o6�Л%m�R���l�LY���e�s)קq�$�#�n�3A�9�:�;�������z�U��m�^l2�[tqx�z|�>�Q�q��C'߃n�Aԃ��9�Aݔ1z�3;ז�Ә�2j�}�Z�/_^{ǽ�4��CA�;X��I�cc>b��9��Iԍ��GzCk���w��r�'K��p���1 �;)��;��9!,p�[Y��rH9�y����L�N�0<�\�R��y����d�xΤ��Jpx�NC���AcT��4� ���a�����cvJĒ��t�r�yc;�/c{�s=�W�}��m^:`��^��Ӷ}P�w���nd'S8,@��=6�� �nݜ�f�pR�So��u���4d��WR�<���w����C��\�4\��N8f]�eԇ�^r�t([�)B{n��1�w
P��g��d|�w\۴HQ�tf �d��{��g�㧀c�B냵�.-��؊�`�T��ˊ����t�xΤ�������+b�vs��A�@?x�\]���0En�Uۢ�����Ee	�4�rؤ�0V�{
r���6��x��J�
�Ǜ�U�yђ��fn݌c  a�]sӔ�#���3� ���B�÷v��^����M_Y
y���B��!ET޸��U�*Ȓ"ibW��
�$���0�1�N7n�j��@5J�l�}�L�xS�C�7W֡�BPD1�C���N	�A؂*���T�'gJ�W՗�a�H��p�Q܇cT�D}��|��xc�:�nc�����^��/�T���{�9�^�IB�5Z�-��3�������1�����vF��ɪ�c�ڃ�W9.ES�U&��ӎ��������d��e�m�jձ�]rs uhs�ˊ���Bi����^��:�Sp3��2h41�L�n��mY�=�������#�*�mj��Aax��� �U *��A؊�W3�s�A~̎�]�v7��[W��s����m%�A%95��N������K���q���E�xawތb;�5�ׅ��}x��_6��qI�6�~a�(��+�z���u�����Ւ�F>�ռ�5�gÇm�����}�8)�'n�f�e	>�hn����+|ތ�˪�b��	���\�4*�g�g]�.�=���w�;Қ�NA`k��xfн1�3����p)7x���z7�����,��Os��Rt�T�v�p�M8��L]x�t�zj���.y�8���wpA9)� �;85R� �i�Lq�Fȿ^���z�~��~Ϫ�b�C�Z(����`�]��,3g[HL���-C�UB�$�&�o��N5H8 �T�۷�f��_������pb#�c"�_�f�yb=H9���D?Y$��v��0B�bNȽ�`�.gS�LRv����fsM+mt�o,�O�[��(����R�HU~b�/-[�*cɬB؃`�h���:�n�6�P��+
_|;��B������\6q�� �{�x�;7ߘaw���T�H5W3��^�14���at-y�8��:�-5w8�MT[��;�֠��tZ�a�l��_���^VL�:���47�Վ�+�`qay�_��Pxbٛ�˜��_���yV�Wy���̣��̍���޽T6�c2X�# ��upy4�����0���s�^�A��"��R�r��w�3���;X6�;?=_b'�
�qT�}�'��G��h�C��!�hHC�p�{a2$v�n���=n��(���g^�h���}��5R�Uw{�!d.��>G�Ox�j��w��.�E�@��*�ۘ�hMۍl��e��.�
���u4������|����K�L!=��W�HK�%/e_,�T������n�V�ê��s�Ƅ��]yA��Yfp�
�2�1 <����ON׫�,���-7�2�L�w�����d��BR�e��}lК,�� �� U!4��v{f֩U�}޼��U���Y5|�0�M<��l~ߟ�N�~wn_��OmۢԵ���pdk�S��f�ՙ[��u[��Ck�o���uc�+�Ņ]��pX���E���|����35���/:��' � #�l+��ʓ]��a��=z%��`{�碹;L����Z�1�1�6�cbᣎ.�l���>���N�Z� �q��zq��g� <�r!3�Yƃ5ѥW��Ḯy9��E|�����skĻJ`�c7f�v�]qҞ@d������!䩺��<�=���K�`i�v�M����e����i�g��=�Su��(�mU��]A�;Tn�ZmS׽;�yyk۟��j����35u��po۷�|��U�2p�4��"m�ȴ���qU���^��{L�W�>�������O5ų�ꪜձ�O���@t�����'�]�%���Z�=�p_o#/+&��&4���y����T�Mڋ�ko���|r}{��]׋[�^�d�Y�ꬢ/���OL�L�&fn3�'No��Q�.���ᯞ]U3��x�	��1J[̅8U1x]:ד�矾�i������P�ct�pOu ���'[ĕ��R�����xs2M"�ZI5�>�g��f�5Kv�y���/+.��sf#���H�� ���L�v���h)����	�~�%#QV����y��ͅ����_y��z��&���Wm��W/�F��߱�C�`Ê"	�m�7�wo�O0a�ޚ�Q���������aٮ���ѧ$W�coM5�	�hL��.n�v��8�ݽ۝/��U��{ �d!\��Be6��W~���:�g^��ɧ	�{3f���F\�]_s¡o��>��GR�R�U7SL�2�e5�
z3�z1��ųɽ1V�O��^�6�.�x�뙁�1���^y���߿��-3j�9N�˲�#`�6��M� J�E$�xu���Y�ݫ%�e
�mn�}>�r]���>I^E������жmСM���i�q<�'���N����\��茼˻�p-��D�y�]�&�/�P�"�T\��&���"�{c���q7w���-��LLpT�,����J 7��qP���,1�%wy`�]X���a瘕�0i�s�&>�.본�j�!ij$,��wI�ȴo��6ie�
ok�Ǖ���q9�Ǝm�6��P�z`�ecG�;��ə w}d_`.v�.����WvЬ���p�^�8���D�U!�k���ܾ��Z̠��4W��a&���-�*Y��B�au��y9_,���QmI}�,��Zo�����\65�2B�M��m�]S*F����v(��ݥ���8*�(�Q%�z��)5�r�-3o��09
�[I��� �1���S�W/+�îv�u�w�y��߸P�Ei:���h-kI*���Y���V�ݴv޼"��3sJe<�Q/0�y�.6�%KF\�,v�2njl��u��s�>�Dvv�ι����W��oD��[���9�r�
{zO+)ຒ;���g��{b�K+6�s����a���췢>ͧO���VZ�u��W0s�� ��B��#͢�%#�B��76�뫻�+�+�.�YfVRK٫.��W��-�g�m��8��Z����M�'���ܛD� kqb��ÛP�V٫�v��S�%�Y����lţ̶�����oŧ���4����=ι�+2vd^=��J;��������4���]vY�˯��jlJ��/�2[�/��j�Xf�%a���U�]'�:�+��uH��������՞����&�Wt���x�'��D�P��t]סY��?m��̯8>Prw�u�*�ؐie! ;�KPk���;9����ZD���#�!�D�9�
ԸIbX�����<Ip���*�Mm�C�� �ı$���Up��UD�����2o]�B���
��j��ǧ?gO//��><<<8���>�m��H�����	$-�����T��D��\��I+��={q�맇���Ǉ���������`�Qp���U�A�S��\�}��Q��|'�>97�$0DD:VIf?�����u�o�n�^�_G�nٶZ��� Qs�ABdQw���iV�g�aUEr=��e~�'8y�\��?+�$9�")�!(�C �Nv����J��TQ7���X}s�N�y�(���EE��$\�����̈�9T]$���2ږ�SNUTs�8�Q�D��������9j�D��d���Ȏ~;�=B�d�hQ
<�=H*44$�s����hA�QS���EމZ�we��G
e�B�+�!̴�(�P@�+Ew�Q�ؐ�(
9���B�2*"���)!���iݼu�+n^�2���k�;L�v3)�K��y^�� 	��=={�\OTUg��u�!󘺳�N_VF��T�L�&TϞo�Z6a�©�u�T��lF^e����!	�=)�f���q;��6߁��g~��Զ�x���#狖əoI�|]��vyV�ӻ<`� �U��ˉ���uO��o��QK�f�����%����CN���P�Be4w�(m��O�4f�m�k�]U������`/����E��NWF�H[G8�L�Je��~Dy�v7�2��U�����w\�d ��]w ���U8���W\<⎕6��	���sNs�o�*��v��B�To=x)��[�@пDI�����n����x3��l^���V]��f� .w�۫��wmN�_j[�_+����(]��W�O���WR�.�5#u[���'� �.>���w�Y�$������g阙������Uu�{�E`V� �I��Fb�;Z��UvbA���]b�$ѳjЗ|�g��:xno*�Z��U+Y]u2���w�W\�4���v����BmŦ]�|1��$��߄�)�j�T�+P��h�u���|��]m�R�L��zh</M�)����3�
�g�Bc���=`��˷&�j��2[��ΰ�)�ʙ\�*�܊��F��`4����e����2�y���򪬓���{ƽ�I��,%&*gk 윈	Mj2�U��
�"��)wq�@v�T���\߾�"�C{Dǽ`�����O�Vupɭ���n��Hk�����W&���� �o�mv�c]�1n�Os�����M��&��q���P��9z�� ���Wh��sM0X�Α�&��Q4�#-�d�Y��Mr�݊���DT�An��]0����ò.Ƿ3�=c�`T��Nlug��r뫺�n�I`�@��n�t��zN��;��^�׊�"2��CR�/U��{D��pV�����47��6�WD\FF�]�<3me�۷Rrv�af��z�-�J~���@f�k
G6d�9^�v��ή��t[s��P	�u�0s	�Lu)�ʹ���.߮��1�i���Dˁ@o{!�P�$��H .wj��@z�+�=�w�W<�l '��[��6d����6R�*fg��I[Q�מ
2:��d����"u|S(	�[��,j���/c�F�:e\�u��
ߦ���·[�B#�8*�C���ۚ��`.�9��駺r̜�S��yYs�8�zfίUś��yy��9 ��BF@wܻ!4�=Zk����>��A" TD%7v]ߚ��[�g� JC"�p(�܋]�/K��h��vEj��}@\����������f+3Ʋ�/%>xѸ)���n���zX��X� ������u�^�;`$�������**�!xy{^��n�<���X��:g��������ΰ|M����XӞ6c_�	����:�v"�b�¨v�{�2w�&�z���S9���Y�1�6��&4�+���X����#v�(���q��M�r�{��(���Փ1K�p�&tjv2'iw���@�끸	6�xZZ�15V{���B�A��zwWӗj1˷:�l�J����k��|�ʧ�q1�q`��6�4��V�N����٥�Ԁ틩3J������~��3he����ݭ�3�ד9�1�c�ddoU_<�O��U��eSU;;U;��z�{���m�Ygl���<tmF�ɘ�p�7��9�E�8��}�撚e2|-}f(ΈUC��̱gNm�UO�&3�}���ٞ&��wM��]@�T>k06�N2�sϠY.�{�bN��$?��'cs(�$��,�b<7Ɇs���jj��j�~��S�E��^�w��{�r(Y���u���}��\�k&x�Y{T��Q��M���X�o<�@����6n4�wC�*�=�6�4��R�a�M�3%��蜪���U����$!�x(�V���&�%�:�ܒ$��)�Ô�Axu���|��ڹ�J,XL����ӈ׻,��z��y;y�H5Z�`L�vM3X���}W�4�B��{�k6������z��L���.�ݙC[��n*��)����{�>?�C����]�X����d?�T���4٦�����OWg�ݜ-�vJ�\O�{xGi5��j�<ή��x�G��q4����5����˴[%jG����'���0�|�4�L�(3!��+�p��u�5�5��]_u���B������$��g� �"���T���-T�B�6��l
Kʔ�e);[�y>�t?�׷������/@)4�mf���l9��v��\݌&���$ٗd5�|�䏪I�!�\	a	���iߟ�w�d�Q�z��צ�MZ�y
�2��ڴ�^�N&��ݎ���7	�_W���p�UJ�P;۷v��ܛ��U@��"��߳WB}e�����f��{����  ��&SL��<�&����P�����k�{iE���h�x��凭=�*cf����zצg��J��>���6�qڹ\��i�ׯ���w����a�g�`� ��� �]�����g!T�]Q�S-�ev��k%e�P:�eǲu��_s�چ�z���zԜj4b��Qp�]�F����7��ی�7<��kiJ�V̕�Mۊ
۝��������0�j�K�t����ƚ�����GP�u��<\Y6�7"�k������X�[ۤ��Mr�t�0��q�6�Ec��O]��vz�(�c'g����u/��4����u=]� p���)��j�$�vT��>�=�m��E�n��Y��Ժx�y���<
Mn��y6����)�ie��1u���׏j��4����OMV����MQIw�m��H5R�մ�l�fd׳�����J3*��|���A�+!���MU�=�q���L��C�{�w��w�d�Y�9�i�&|�,P�izS��ed	�e4�.Ӝwo�}n�nS�mՑxM\��xN��@g)�3�^�fa�ض��oB�A�kV��ٙ���-�К���;��n�-��KK��!i3��V�:Fo.�`�W^���I�є�g��h�&P�hꇣ�^�x�Z��1��N�:��䗯N�1���]Y�a��,X@�[�=M"�
���ɐ"���_N;�Չ�9����S��z��
�P׽@TcT�	�=��6�؇߫2<t��y8�5�JKZ|�iY����+5D�3Y�Goj$��g�~�N�Y�ۯ�cүf�D�^�kY���kϧ��<��r��8�q���̉�׎����""��=�F�žϼ�~4�RfG�������K)I��T�g��]g���no�=9�zr�<OC;hV�|S)�&�N�n����q�ss�"t{_c�nv��e4�i�2�"ēo +M�}��3��3*k�������@L�u���L�5���7}E	J��4���l\!�&��2�фa�K���e%6��Ԗ��V�hoL�	�w�q������W{�k=�I��g\[ўƆ<�S[U �S}�V��Q�)��g��㜵=g0����S3��$�������2�-�l|=��=��Jo3���]	WW(8%0���6H'=�u7�Wc���:���[�a�Æ�={����V7֫,�����0��Q*�l��$� K]FD��Y��5��� �� L4�6�VJ�� �
��9���裡-���v;�Y�h�^�W�ʣƕy�|N�e!0�f����9�(iQǚ!&���=�Q�Ә���k���"e�pl���1=-d���_�g�4 ]4�,.\@��-�a�0�m	��vrK4t���� B!4� �m�� ��	�嵲��Vfe�v�s{4؎s�J�Um�7�<�i��^$/\�P}�I��w��\�Kz�ۊi��#%UGs�d�q�L��"^`L���� ��'����Z�X�j���Cm�hl�)�P�N��J���{� V��&}��|f�ue�d�k�=�����NS�:|�T�J�^�����}3+����u�w
%WB�e��wDlR�a
���V��w��4�%S�N뙀����ʙ^b%)�Ӣ�k���vC�yI��uog�E��2�DN����EAz�Ҩ��	X�:꼦�QV�pG^y�2ͱ���������|�>R��}n�r(L���圵R�9���+ֲum��<���-0���*�&)�������߭����{ފ�V{��3*��wBot�娝�ك�Y��q��
��a3׺��Gy�^��yI�=�՞�"��S)�̫%"�xF�u]�=/
u-撮=�Ϛ�W:��f�h����*�����7v�^�U\Ug����l��Bg"n՘λ˿eq\�	��`36 k�{{볗�`*��PWGn��۵��4�7x���g坽�[�0l[��ev��6���f]��;�2���jQW^Z�yX�gu������q�@��GX%� bM�`(/J�۽�K�x3��v�+1n���'�Ah�:��Ċ�Xn˂�'����G��v5���~ɤ.�U�j4O��$��-�jh�ˡS)mE`�G��_�_V���s�<�f཭bm7K�6�r�+�.��-�E�0;�=�U�u�ZӴ�Z�������nT�.��#�ՎaЙ{��-��uJ��0Llǧ3����Xpu�9746�r��Z�*^S�"thP޾�ͺ�;{�I"�UЫ���y���xb�4^k�E��k���U�w�lpݎΩ�'��Ս\��B�m_4���u��{�"�A��N��;�Y��1��H����l��;ddi�	R�T7]2u$��k�{Mc�'j�)��ט��ɷf����\V�W�9�`�����3	�o�s������h�+��(z^ �,���ו�$Δ�-�����0n����!�M��Q��Cw ��'�^�z/��=�_n�f�ѫ}�O:��4�ǘ����U�����!�v�Ge�Z�ƪ��Az��=�ǛTt��:G��S/�1���������0��X� �/7�:�n��J�1p��رm��R.5����J��哭^���g5���T�a�]����g؍*�G,�� ��@Ucf�a��}|#=���7����Ϥɹ���|�����6��ټM�累 �K�d_6�$g�AʓeLQT"����[��^�ߏ���>�6V�ANr��9��2��]2.R�����Ȋ2�r�Z}zgO��������������>�ot_RDTQ�#��O��D_S�� ����ˑs�X� ��SƸ{gO��������������}|v�CLoN�(�"����U�"���D�QHI���\��QTL9T\U3!����9W}��D����W9"�)��r9T����.�Up�Ut�
��JL)�һ̎r>dDjEQ=J���R��|N���"d��bD\�(J/2"/'/K�ǃ�*|�r�(��E:���ʨ�".rH�29S�W�W�����Dv}A$D
���eDr�ܽ��Dr�G?�(��Et�p���Ed�*�P��"�U��?�OP�/�����QT�T����<��&mqd�����ք_Z2R[���Զ���/���E��цe�k�C
ڷh��X��uq	���/��8��&)�������s��ê�����vx��t�ڃ>5�r9������%`�5��\�fK��+p��ٯE��p��<�=��4�>(qr�nM�ݸ���t]���ݢXS���ɬūkD�8�׵��6��:67tm��f�l�I�U�od�۶��^�J���q٥%�1��.�N�X爧D0l�ڇk,zї:0�b0s���Ⱥ��#����g�����lk4���+2�-,)��ɴ[��l�L�5n2�V��&�Sr�ݙk���F���:�D�q��<�6[�N8�gT^��(]D��X�,{HVc����O��fZ79���nUts��B�V��@��`���B�je�m�,��.�gxd냚��:+o��@�MeRT��X L6��i�D�m+�8ն`��+�tWZ(]�`���{\��p�%��JXa�5��Vd�q[0T��q`���l)\��1���Ku�03��Ҹ��0#��K�
�h��&����;n�ٲ��s�})vlc����t5B[�h�B�T�{��LҬ+ �Y�.ֲ��Jk���8��y-��늽V�k�Nz��Wn���ݎmP���G6a���u�����b�xrG^5�g���z�N��nnu'*6k)^L��.ܘ���uML�#4����!��B�iظ(s	e��vs�`k`�6&���a΍PQ�j1�8r$;b�n����?n��#��k���4Hˡ��1�a�F95��6(�!fLM�0ݭ��tOVMiQJx�V��Sv�
�v;��eUj��,&H�uڳ)t��,5�NnI�l��ѵ�sd�p�Kjz5�nթrj*,��X���巙�.ſC��>���6���������8.s\�ͦ�P����r䴻��\{�;z�rWki�ui��c�I�y�<�06E��JOh����o3zluۭmFWQ�Zd��=�;]�f�;\J�Y��\Pbm�s3�x�0m���]	�������b�t�j��7�������ސz!��n�EMB��KXz���;����t%�ps���mD�v���a�(MB+�b�DY�ki���3��[���s���k��]�ܜ6�y�:�뭆�8$�q��%/O]���c����c5��#��"������ص'b��e�A�$�_�Rj�j�T�{�\���k�ǳ�6�>�,�ɦ4�օ�4�*�j�=��}`�J��V�n�����f���5�~���n=> :��w����M@��O��W�UuQ�^��˿Np�t&��<��4��Nە��+è�r +��i�7��Ei�[ֿ{=��P��xg�M�(��� y���L̛<$�������xEt�����a������n��"�t�Ζ�1�D'0\�sq��g]f�B�VT�R�<;�D<)�)0��\�˳̦�|�;k��yw��vw�wwz��r3��;� ��T������w��v��%�'`�Z�;O6��v�F-.�;������z���i���͙vFg��^LW��t�\����U�V�/+��oʨ~����7rV��}}�1�=�*��$�㼦�J�ѡ�xU�y������f�mY����ǽ�o���a�����P�&U8H�S��[��;�s9�l�^?��Z��f]�s������g��_w[�+��30��*Zg��]�aM�����7"�=~e����i����ѹ=Y4.|��O����p����!�Զ���������ݮҙ$�O&n�4�o3=S����݅\fs1��\�.{7���ǵ����J�V�i6ۨ�9f]��;ٙw��K�Ba=2D^�D�u66�g���S*e��C�˻�K�U��o8B���wVy^�m;zn���l-eZ��o�[/F������4-ѱ�#�{�xn� ��^N���=Gy���{��&f��ة��x��#R	��L�l�*�u\g+2p*n�B�êَ��`R�= �Q <�����ڮ�
���}4.���eߧ9.Л�R�<��Z����S�D{9?/��)}���G1�wWY��(��W�a�Ƭ)�S�hS;�TDR)$i��
�'��L&VxvȡS�]s^�Q�mc�.�ފ>����6r���T��wt���i�~��8��\���nNc��=戛NN�@���bѮ9��j0�;r��mOq5�8,��fe��r\�[��W*�&Pv�L��J��ϥMz�
�U~�&{���s�̏ "S"�U���׼�w�
}����:�E*�>ו��u�*9����|^��]_Z�Q�tۚ��r]�Z��(K�,���y��<�)��2��Bg��������]���a���9���h�-�	�2�g
;>�P����)�����NS��
�t�g�8����O���t��<L����e���mL�2�g]��}ٙS3��6n�w8S�	�V���ɝ��4�a�t�ߟ�+1��Pv<6�*ewW]L��b=Hv!U���^��o�D�y������&@��m��$�Tq����9�����b��<Ū��S'}��[°"���k�5oNA�yٙS3��=��je�N�g,\&��"�co8ֻqLZ�I�z��o��y�/Hّ7&���g&�p4���O��Oյ;����_x=����tg�v�w̜w;:q�٥��(��9Qʙ.��8r��n��Z��ѣ8]��by�m��P;
�BK�l��eܭs![�R�d4�Wu�����p���cW�Z=��6���$#p7�;�E��4�u���j�w���}�͒ED9���t���㠀�vq�|�5g\b�����#��n�;i��fSҘkK��u' ���Z�S���F��f��gP�u
��kLV��rs��sv9�����f��e��_ϓ�g����:��g\몑n��^9�ь�[h�Z���������/���la&�M2��	�;.��j�Gc�NN���<[4%���ho5:g�2�V�ڗ;�MT]��9v���}ٙS3����O!3�����>�pZ�{�'�L��g Z��׺�P�5�enm���U2��6��U&i�2��d�{��6���5	��S�8���Md��N��.���rLd[�^�oT������D	�L��<���>�7ۙ~����	���`L�����u~�;�?{����\���dR&��i�Zqkv�l��۰��2h��c7�
�&P+�:=<��k��r��{�o���}��mi]�3mT�3����/���N��nc���V_t�D���J	e[�/B��-��%hL�[W*h뙵���nu�sc��	����g�3l�(	�ꜱ�s�����ap�=�T!3�su���S�%$�n��S\�2���"�N�
>��+�eET�%�WK8SL�3:w�{��a�x]!\�v/1R���2���s9R{�%	���e|N.��¾�[����3�۷��K{���wo���'&�ѷ�⒙A�@3^��H�$&�8d�a=�(AN��QcA4���n#c����J]�R�MB]��e������	���er�{��f�TUOb=�U���T�pm6r�ZƩW�$��~K��:0!���u6X�o>�;S�����h�;O�t�t�Xn���>���7��N��%��IQ��{�s1��Ŵ��iW)���ii��%��x&.r������kyĤla�r�O��>��>���'�0��z��N��NM���V�x�
�"��S���/7yF1=��W�Ο��ߏ~�'V�-���k���cԇ({Sn�L�L&�[����K���?��wnU��>_��5�G���u��-�U/q�=�>C�\��%�ܿ�����qi��'/Бb��p���wX�.m����{��rZ�@�Wd�)�nr�j�OS�NNQ������/���d@ �=!���D'���Ub��F��j�̨��x�8y���6�6ST�&�t�>�dG�&�X"���)��o{�w����]K�*<˸F����U��T��Oj)��Z.���Ba0�^�ʱ��g�*�'Ѷ�d����z�b�r�_?-۟2aMR�Lͼ�uw@{��sq��e\���7�$N���8!�s��6.�e'��6��>U92=�pHɂ��.ӓ�A�vQē�w��@]�3Ϛ�'�{�ssn�����Y�9]�#a
�2��i��<��6��?i}�n�C��g]��ev�H�H:G<=��)�6H˻�3� Q�͌�|[>��g����s��=vR=׼.
�{:ZeN"�ey��2��v|�
��e�Ƿr�n���z�rp-nn�j�3�ΝγI<?��)b|��~>�����SL�8���Y=jڏ�u��}��W^]��e���*L�1�UV#y �g�]y1i�'���Nl�;�e#�"PX����D�F�[�m�j�aT����c�i���3]wu����W��'�Ŷ�O)�g@|3��w��ۯ�;� j㢄�� U��QU���f&�]^^]gu��F�f���{uʗS��שZN�� 1�A¾�<8����߫l}�� �=x��B2k!4�MqI���ىl8�����sڗ��7/;�Eb�4��c/W9�l�m�����n;uF�z��Q��+ki���`�+���lKf|�	9��;��!/��*�#j�cK���d�[���t��m���d&4�ɠx�Ua���Z��X�Y�[�E�c��F-�!՚��&��u�[�L�u�׹�~��:˥�g,�i��[nT�v[h�ۨR .f�wOD��S���X�q2n�HzkP��=k�����z��7j}�-u3���i��+��+���ۮ=��Sk�fUzs}4�]��Cp�����9��s�%�Z)6r|(L�Zg��8�����UD�&�$g>F�{�yX���	�<�Tʰ�A��=�#��ƹo*�V���(��W^P=��Vj�7��nY�{��p*�U;���"C��h��No���r��h�è	���u����ܑi@F�kAlm��R�6�+�N�$��d�lG��i<���2�eRߜ�����ٴ]SUӁo*����jZ�Ǜ���\��J���E�ti�=w���w�WB�������0��'�����ҦpTagl.����0���ҝ�i>�30���C��Y˱GfWU�k�X������{�r��=�j��V����~z�*����zø�_���N��h�4J�Bg�&:1�ܧ{���=}1�E���S�L�����ޚ����.naظ��G{q�4귌)ܻ�ܵʛL&g��z��W,u}��������4�%̽�ӷs�Ǉpwp<(�k��8��cJr�(�R��M��.�1uw4!���׹�ol�+�P�~��lԾu����޻1�=�gDʎ�{���M�T�U&-�����V뷪�,n�w��U��\ �CyL�xr�$&�/�dbi �2��S����/���+&��ȍ�o9��]��N��gV��s��� y�u�Oq��ͮ��2�i��Ԩ��PqTE�at ���8��3VU�w/�ЧW���	wB�|nLU��iY�8�Y4����y�Z�N�e��<�O,(�:�FU�˭�2�bfd�5M��%^�.��2�n$ed��m�9�Ӽ�C}��7�v�$TB��(P��a��n�s���X\:]��i�;�j���}�B�K��=ȷ%�F�#^�*2�F^]��iԄ_c�"�Ju}"�W���<�&�}���S��X4���`�u^���<xv�����5Wb}�%��M9�ǹ%�s��ה!���%�ם9ŝ��t�f�]�FV�"�vv��Wx�R;��Uη���2`����f
V�\j᚛=m<����γ@|�P��] �n���(ۣ��j�飑s��5�í蒹�),�����+@�N*���Q�M8��dv��+s�l��Y��9��go���vV���e4ع�m�;�gj9�\4�y\qH�HR�)�ٙ�K!L��vwH=]��b�ڳ��(�V*���Cf�v�p
nڂ���6�E��Q���$���it]�vҵ��j�g�qKn�{y�_p�mT�|l���9¸��%�Dt��kh��[Q��jo��kt����*�%���"�CF�byW܎���񵶄5������WP`�./��e�Y���ج҈�uh�i")�B�P+���B�U\�����P��Ur"#�+��t�Z��;q���/Oo��o�������e�f���"��'
"���r#�ET�'���|g����ׇ����oo���ۺ ��s�(*�����R��zx�r/?׸�0��*�24�QRSY��^��������������}{�٭:*����*�Zr�c"9A¹�+�H��6��d\V$PR�bjT\��$�\rB�t��\�̎EET��ԫ��QȠ�¦wDuer�QRel�8p�-��PTr�(',J�!�%Q�&�Y�W#�Fe%faʠ�P��,R�6�	$!D�Ne�2�:jJ�Q���+�έ"""�����絑Dr,��UD\i\�T)��U�H����%Qʨ㢩���Z��th\��N�EL�R*����"�$$)Q�Ie%�EG(�ar2$���VE�K�艍�����߫]f�m�2��e&,g��@L�N0�^{�뾖�N7�F[5/_	:O������tJiЎ=n���UbƠ6��i��*f���yw��U����}�'������i��"R�'ތ���戦�"�$�Qne��"��pEݵ�"�-j�t�b��n��~��p˵�����n�u�y]���<�I=��s;�扠;�5�(4��m33�۞x���m��r+��������+]��PG���2���ͬ�~'��(������&�B�	A�s���/f���>����FZw���B�JE]��n�ï0rƽP�e\k/J�y]��M����Bמٻ��;H��[ל̷���[��nև�l2���Ub�ܺ��ݶo'h�����uFDhh���.=�(��q�$�'��{�T6a��Pg��ɐ�B|jb�\�^�7��[6��.��O]Yy��{��ZL�	��P�^�i�0i	_"?���\Hu���!��r�X�SFUl�¶�O_=�(��4V41��ҪA�}}�zu�TU^^��~�]A�޶��-Iy��U/Sߴϗ��:�� �c2�i�~��y]��Y.�{Ӛ#��W�j�Zy	n�ammg�f 3&8iY����?���NN]Xfb=��[ԆM.��uƞ3�!��w= w�ܛ�0�C�}W�_x�EU��Z2рf����V;d��D4�x{ɪ��`��F�@+����[��ː�6J�S+��0J��<��R��0,��p����.�����X��Nd�L+����we������L�;(��+�ʅ쇫1(9A���G�0Z7|q�k��PP��c��L�l����rU�$\u�w4*	��P˱�&Ѭ$������Z7����4�1ޙ��Y�ƚ�jj.����T]�ж����6s;��"[\�n8詸�C���k�qlw.1W�)�1�b5�������O�q�&��=IsO�0�n#����a�t]���cэ:4f�#���aK`=a,a��h�F]����Y�Lb]%�evl[6����.��֣ωc��'I�QU
�R��Ra�L��z��垩���G�Dﺄ�E>��z�3�t	�y$���1��=�vs��+�?��ٹW�{�b����-l��G$�f��񴕮۟1g���f��JJe�a���#�9N0@���o�6on;"��Fy5��i7����������T�|�)v@�]�3�=sS��1��J��KUH�/J2��ͬ>^��*�4m�]�����=U��Z+�eL�/>���Ӕ�\M��T�B�$6����&��-1e[����`x\�6��8 �'�}J�d(b��{�q�7����ɟ��zgj�W�N &T�$�z������O����},hu�ԧU��_j�M���gO�����uu�x��7�WLc�FyU���ɋ�y�x�>��83d�� .��y�Y뚞�}ي�p���3���8���Z�z��q3/g�e�^&��r'{�j���E^��E�_X��A��{�~[�-q��  �;W��A��Om���zo��b<�y3Ծ�ø�Ʀ���4b�ml̖>Mv�fϸ��F;ō�ѷ�}sU��1�ɸq5��]�>��*��h�o̱�\lf�m����7P�wF�u��Fa�'$Axu���se&�S>g����cw�G��^^��t�k�v�����n�ʙL&e�Z����t͘��2�v���@�U�r�G�y0�Bf(�쪚˽��x5��f�>lg�P?}�k@��ȨH��%/�o�v2�^2�;GoY��e�����w3�˺S~�7�c�b?V���R�� �3��[t�-�1[@~�0}�޹՞骻ۘ��L@�Ck�iU ���%%�ʢ%���E4ǯz�v����������w�/2�ա� � ׈w���Lo����G���o��9��W�\��q�G�<�5uOO�ί�[�@ů������Mi�nܺ	`酦��.L�lK�+�w�E�^lg�g�t�4�q;Y�Mm��G�v���a���33e ����s�o�q��7����w���+*�kn-�i��l��c6�	�&z�ͷ~��S-q��푞�yƱa���|��L�MT����)",�v��\}�|�����嚤��_��f�BZk�/�d��^���M�d+�b�G�_^�C��MZX�e��ut7���ַ���
��ip�:��P6��߽^�W������]Hd՟���4�>�?}�W��.�rlG6�a�,��9@���ro����`���v��Fւ���v(��9}pHl����g��RAD��$v׹��Be�\�y�=�#(�u,$K�<g"#/���Cbfڪ����'��{�������l]���'���?�x[���d�'k�'P~�hmc�:U3���N�񝯾�������Z���'&Ǵn&�Be4��p�9��p�I�1�V��c=�=�o��#�z�t<�
Jt�71���5���]�T�4ʓT9@�mcwf�}��Uh>��{�S]L���Y���=����"���������މ�[]��C]b�ݵY��q%a�)u��z5�n�v�u�e�~W	�/u�H'�^7�B[�$�=u��ܚk��\�;n�:��� XV�iwX���Ym6�iއ��tn�����ꋞ�^y������'g��e7<On�C��:�=C\������1s�)T&!.��ڳr��㓦�n�9�h���
�64mMr�q��ڑD�˴�Oluz�6���HvtU8ݭ]g.�lK]X�����հ�Q��u����~)���5��t	�.:ƻ���*淤	xd�T$��g^��|m	��D�z��s�$^d�X��̽Oה&T�m5H������xd�/4�5j�{b3�NQ�֏6B�L֕3Ƿ5�I4˶�Je0���}�uW�~���X�p~��|�_��R,��5�럝Ξ�\�L��\��9�+2r�{F�ڼW�Kф��)qm�l��mOت�����
���TFd��Ւ�h��U���Е���'���~zO�6���ICBi��K�B��K��jC�g�k��м���P�}�����6}9��Zӓ��V'���ۑ����;�N)�3/)�?}�迺����uٷ���N��u��1潓����� K/c�!H�9��4�T�{�}��Ƕeu�X���O�Vj�&C�C�a;}C�ݓXh��H��eX�������Cܜ���yT�ffnO'�ny���	�Ւ�h�L[!�v�2��\p�x12��G_�a�W�4������Ϧ����G�Dڷ�2Ez+q�R34�Z�.�]�S �y���3�e�����Qy�bn�yzP��.e���rL��<��_��VjAҚݘ��0�gX�T��w7�f���x���*�s]�m�&P�Z�+b3�'+�K���9���<��j�	��(4�[���#��Ν۩<�+�����^�T�3Ո�4O3ҙ7�v'=��T_��(�NR)WxW&*e��W��TC��y���~�Y'c��Kˬ]c&�_ry:���F_�m�և;�Tϙ,�E�c�rK�߁��,��w�{w�U��S�;Wg�mFfz���y	�3�zjw�Q����mWy�ϋ� &P�y[��9\��m����sƭ�gƻqv�������݄���o��/S���#���v몀�8*O����~������ڑ�l��t&hoN�vΤ;{#�t�B)^F��c�92Էցb2�L�2���
՛����X}d�e?�b����_��rn��HL�1:q��z�,�v8���[�����S�֏sg���;y�5��ja��"9y��"2�iU!TcK�w��r;=/Sd�V*]���m�Q�2��7^<�����i>�ϫZ���լ�R�3����Wg��F�b���)r��%����>���F�d��]���7�vM�;o�A��������՝����]]���s%܃����� 's�I%��@f!�3݉UwG�B����;�>�vz7=8�f1���.4�2�R�{!�S�S�|P$i�O��q��k5[�(�f�W��r���w􃍞���V�y��q7P�r�t�ub=��1���@9]n�>�f݆f�q����? }|k�A������y���[�L�5/z�w"%�	b)&�S(��30�>��[��_���ѝ6Op�TʙBY1�PD>����L<����m؛��jt�u�=���}C1G��<2I�Rl���O~���)νz���y��p�j)���?���[��^5�DW_Ъ(�K��K�%@�t:0:��5���R`yІ�BP!� ��e�HhV�bE�����@�ed�T$!i��	�aBQBD� BD��EMiC@���!�B*��DT�0C �� �5p �!*+J�����WB"��(�!(+J�����CJ��"�����!*+B��@�*���*�"����B�����0���"�!
+@*������!�H*���442����!"+�
����
,3 �!"+B
´0��40��0���2�����,4 4 C@C*�! �@�ʰ�0	(�����D!��i�Hh � ���B@!�d�%�BP hd�U���B!	�$B�H ���� !� ���B@!	W�s����4u~_�
 �H �$ʨD��k��?����?k���3�?>?��?��a��_����+�����_��:����DW�����O�TQ��D@b���>��������P�?��� 
������O��8��C��2v�����y���P~a�-��dPP&  � BY FX �X �U��`BB  $ $eX	 ��d @!eE��X �` !Y	VE� @�d$ �`eYFF@%$Xd	�@�B!BaB!B!B P�B�B P�(QJR�@( T�EX�EhQZQ�@T�QY��g�M(+�TV��AX EbPVaQd�Qa��Y��X�E�X��DV	X!U%�`%Y�h � &�P&  %eX�BU��a FX��`�e��d�I � %�!Y�	�dX�
Utg�-��߫���"
4
�@��H��}�`k�W��}����������DW�h?�?��tП��hi� �n���Ȝ����*�>�?Z~^��'r
 �� 
�����C����~#�"�*����A��C�����h?�5�yO��3��`�" �}���w���������� �y������I���0v:@z��
" ���!�t�I�/�h� ����?��?�x�S�N��Q^S� ��?�� ����ݯ��o��*�(�����������������/��0����d�Mdq�L��Cf�A@��̟\�S|��                              �      � �PB*��T 
P@��@  P  �PPH(J�@R�R�(�  � " @%��*�%
���(R�%%$%DR��!*%�"�T Q*�!J�A*(�@%P�U"�T�)*P_   UBT�T
�H$��h5w�Qn�ǉB�`d)y�Qs 4N�-ހ�<@Wu�DP�)B� q�D{�z�����
HP �W�  ���gAAA^#W{�(<x�� PPS���� �砠��To0�.�����I)V�[�q� ݞ����{9ڡv�DP@��  ;�ʨ��Q*
H�B�T�}5�w�B��y����v�]��=����T#�V�'��� ���U휵JUxUI�*�����^��KhU

D(>  ��i$��jQJ�䔎���]��̶¼�Y*�w��Ē��$��U��B���B��=ǳT�=޼�+N��"�	E( ��R�HJP�J�D"���J���ү-�R��wT����J�r*B0�UY�PU�q$+�QUa��Rr5%W,� �=C���M۪*�: ]�*��"��UJ���$S�UA�zU�UV�被��EU�UR��� (
"|�{
�5B�J*R
J
�$�Rx�L�@V�uD�۪$�۪UpU*�ts%V��%VF�� 9�Up NĀ@�
	 U)� GxA� �<�' lq 709f d.� ]�!\ �b d���` �
(
H�   ԂAIEB����U@� fǐ�@w`�� ��EN �� ̀�70�s ����v0
���(H +�  �y��@��W��>�6>���w 9R� n!A� ���9 .`d�����(5=������4��%*Q�  =�L$�� l� IU4��4i��)*��2@e����J�M4 d�7�����[��?��[�ĒO�$6_O��vç(����9thCo� �!$��� �!$��6?�o��cm� l� $����x�|K+_������W]���VZ��uU�.KG�h]i�vU݊J����֭��Ɂ1�~�	�uH�E,CeZ��:�JU��m@e�͙��!J�\�Pm����5[z�v
���l�t�аmǷ��MJN\kj�75�Y�ߩޜڲ!&�V
ۢ�x$A�^�@�3b"Lj���[;oth��+-�Ja���{O���V�����ʴ,������pU��Ûm����>zIR�E��,�X�)�Km�ej��!�ͻ�pP�*򣂥��f�!{���U�u�;mݡhUK�A����/If�YW�.�7r��qP�ٸǲ��U��A.7F��š��l��N�,ȥlE�daژ�[w�^)b�\����,�7l�i�{�f�F��TEƄ�Í^ja��P���+��e��\r�du��5���o`�I�x\DZMJ*UV"�Q&�!�rG����9�0Ur�F��$ٹ*¯v��Z��Z��ٻ���q�-�ˊ��JܱR��z�!.��h8j��KyK	ȃED�=ƈ;�D������ѮV��J��5!w�Ra�V��O&�O'��nJ�o���{��0�NA-+��۫*�\#2:L��ݹ�f"^��G�3f�m77Dv\N�n��i�wu��j�n��
U�pSz��.��Q��X��e�WH�*���n���D�J^�3N������;9���yN1A��E�l%W���`�i(�m"�1�H�H��7"]G
5nP����f�&�mD)��rˡ�D�َ�6�)Y�P�E�ٚ�`٪�Y�[L���ì91䶖��I;���63\�(����vҵ�/0�X�m�.��0���w2Ї(U��l�tԠoof��p@���U��w�s^�F�m+�qu�B��(��M��e�"6�U�tUU*4)؏��L�����a��lZ���X��n��-��X�mއKKUDe]��t-�9ۥf]�(��̻��`r����T�$�^�[{h��qL�V���whۓ!�@��ڂ���F��YF!��eI��v�d��7���Fde�p�a�l�h͑�ã�e�*.�^&��7�J5��o�Y�$�'ri��\�kL-im��f4��^^�]ƴ[��u]�m3��f�T3sCv+�GKQ��w�7u�tV��.<��"�*.�X(Y�&SՅ^�г2j�u��L����$�K5Nbw6�֢�1	�4��1b��j�-xNXu�7�J��ݸ�,����6��;�o��`�Or�Ь�e�R=܊��ou�9s~�� !�V�،���@h#a�[��`���r
��gXG��=�fG�sdW�6���9.,Z2苎�y+x�#6�{�uVV�T���9�X.���v��mV���f�%�B�
�k����s4�h��\Y�.�d]ʣu�����N˂3Y+$�q6�Z�@�ܼw�����eE����nfP�:�)8�m젫qU�栕�)鬌�w�U���sdR���TA�Ñ���õ58o2���$c�Ayn���;�r��$��a`�w��dƷm�c͏B'vXeЪ	�3HZv�n���ʱ��|��$,B����E^^�6��g^���5���Mz�ջj��a��j��7�55���ٻV��7����J�V��85`&��Z'm�֛�0�Z�w�*��[���kY�\��Uш`T���3T�1��̈́nӔ7@�k+.H��ڽ
�J�$3y��0�Ɇ�����p]�u.�B�A�ܥKҧZf�&+J`7R�M�8���S��gԫ]nV��s2;!i,�Q�4�3T$�6�ҧ���ܷ��Ank��]��gR��m;�	[Iء�5&�YOki�Lu���KE�|��C(;���*�GS���qn�*�̔t$�W�vڻ�34q&�(�T���ܷ[�k��ԗYv�!���^faPj�&ޡy��ZeGF�hV�E+�K��ۢ��ˏ�!mbv�\�IL��wR��]f�@�^����v���'*�ܻ�R5{�UQC���e���A`���NPE��V�f�@Ά"��*�QБn����L�.�͙@���u����%V��Ff\�r�6��D܎!���b��M
wY6�̫ۚ�ͬ�iͨ��U�mMyCo�zڇYCM\,w�
�/onR���d�#�I��U��z��Ӓ�_۴[�U��͕AUb�ܰNmԹ6��,���+2��R�&ൊ���B�v����8�i�h�/^^���ǐۂO3^�V*͇jMR��][���!Z�f��\ٻx�G�m5����۫��e���Н�˧�3��j[3vQ7+N7)�o�f
j��2�]�[z�kr�n�Kڢ�J"\�1�@��Hڬ�+��lV]�c+)ZYNZ	ܻ���q���R0�E�v�UL�t�Y��w�P\�g���r���l�8ɐ�LW��̤*�����n��j��p���L*M�Q*pe������LJ�E��DN�UJ{����%�Aucm�'��ٖN�e��t���"�;R�N[P�x�qh�[`�tKt�[÷�X&bߞ%[d%�/VVVA��"g��D#X�9l�˺O�-7!f��!�Ub��[l)/겪�7��ʶ[��Ѻ7(��A�#7[ٍԫ�[(�F����V)Lݻ�R򓪬�VV)R�Ȫ� ����ٛWA=+oEa�lAM��6����"���1��C��fL{��bg�0�������R�-�lJ�|��D�x���ff�l��n�t�(��7q��w�ȡ�G���ס���,E@�Ŕa�%l���J�["��4�h�j���!Ev���M��&�7
"���v�N|�k0�{v�v���N)��UGu��h�8(j�4�]*�X�c�w5��i����^�����K�*�uy��]n=،g�F \�%k҆�e�"���j���ݰ.]cg5��4VU@�~�U��ܽ��M���!(,�蛇*��r�����4�i�{0c���U�|K�7y[b�ؒO��+���Ӻw�V���U'�.�56#Pѫ�I�n!Knn��g!0�\t�ݴ#(�ۘ��N�o�h%Ku�0F��n]�Bxs,�ܨ*M�˨M�(Ҍ���X���&L��u�)"���9*�:��J���+pbxf[[fL��Q�߮Ȫ̭ME2��X�E�#smLohFZK^T��Y$l���i9f��wY�.��n���߮��U�UuEֽ��6KC,��9��F�k4�{���ʆnR�iQ����˘,�V�L�ǔ	Ӻ�J��1�,Y����ķ7eA���c%�7�
�Mu2���'i]��rU�����K2^e�Ն1��NQM���b͊��h��a��%�&�ֵ��A��!����"�T��Q�e�q����rd��e����Y-?�%�Z9LS̪J}�]�Ԏ�-��4f�z���1m�mٽ0��u[�ki�ȍ �����y�h%t�ʆ�3w[��*BN�s%<��C�@��Se\:�����e#����]�3u5ff]���mlh�UH^+��A�6��Zk$���ْ��*�I�̢�4M��z�,�܏rJś3,*���өe*���;)�c�V���Pu3T!�sY���F�(�kw0�m�%a�&¦�������7�j�&��P'0�H�E������tff�-�*��,�̽�񪭳(�
��d�wy֎(h^ݻ���.��I�sn=	e����އ�0T�.CB�_�Sp�.�Tɰl�{>bn����q�U�������8��t�FU[:un"����.𒓫x%|o����M;Af9i�˻B��{��q�)�۪tq-����ޗR�,��dm����r���&Ycq�L��F��{��J��$Nf�ںc.���\�n��j�E`�<uf%���t�Mz��9�qJ:15zC����VHf�	��/B�1�+.2u%�.�eRU�w�0��K�sj�R�5�0c`��,�'���R�2�޽;���L�9N�SCfkV��$��*h�{���lt��n��)�2��q���W#�m�\�RQ+��'M��*�Z��d�j���${�MZcن^V\���X�i�m��0-�g%I�im��S4�k+VP���ȣ��8�S/6j]ix�V�Ad#��%�7u��yYR��]I�ř0�[���:ؖk#OM7��E����MYu%f�+D3q[�j��;j3,�GtU��I�����7ZN�콪�B��RM�l*�Bx�ژ[�l���z�Ѯa��1%��(�0��hKL��a��ǖ���7�j�l`�=I�Rnc�0���`F�a"�&���(�u���ʚ2��6�xe�qY��W���ۯ�TR�<ё���R�S�٪B��b7�(U�����9{uW��v�흪5H�Z7[��t��!�7�����Ӵ����e��z����)ܬ��ƴX̬ų
sm`�u��m<V��{u�A�&�Y3ɴ%S�d���=[��^��𜩯%ʀ֕t�c��fHB�!E�7I3731	��ϩ˪f�9�s1�T��y'-�҃���U�ͧ�5�$�ͩs,]�8�b�!��XŵR�k*��X]�x�d"���Mnmԭ{�m赘�;�N!�/iK�"�5�a.�m�D.���՗(P��#j=���.�I�A���fG-��Vhn��5/�m�&�������V^l*����
4�:u�e�7�
���ZeWvci��B�7�"V6�V�26�9i-f+;����ɔj�r��m�*�%՝q��9"[j��(X5��S@�b�>����J�e���Ȗ[[�蓉e^n�?^=4fRm�/c/)Ð���ɨ�̈V#��*��f�зM�S(Xt0��6��7xt��2�	�l�u[V�5Z����#fH�p]�ٰ#v�'I8�e�MU���(�YIP��a�����xk6e��)��ѵo,�VȪ[��E��g��n�#������ɷ��5�6�u槵WU���uB�vn�Օ2�*����tiGl�#��ȁ���,�z���cb6�1��̢
%�Y�$�9N�'n廥�W/x1�n�؁��"D]�4Q��wW�fan�Z����Qhfl96�c`{m�y�&kuE�WY�,�ܺ��ٓMZ�?6Y���Ck.�����x؎f9�F��o�d%J[�1I(f�`�eYNq��)/�J�xs���Np�V���>�C�򭭺��K2��ޝ��꼎��($�7Q�ݹU����4���1S����ǵZ�*� �X.��uS^�ܼ�r�j��LV�t���=�&�:yVr��:B�]�m5�2UeA�����v4 ��ڨu�	x����㳴��^a���n2r�Ky2�Vd70n;�gtYY3gچ,i[V*� �,qáʆ�hs2�]�A��F���ּK�z�uw}�Y�V�_^[W��6*�Xݒ�emgΜ�5wĕ4\�{G5��Ҧ��f�*J�m��j�蹭�bU/Y�/&(m��UU^b�K�m8�{�%l[�P�[O,�;D�Z�}ZZ�Vؚ�9�%C^i���J�ʚ�l�D�Xv�$Y%��qU���i�u`�)n+I%eKO42�J�2��Ou���/-��͗�]U���Lϥ̰��(^E��r����騖�[uf�-�{QYl�#ƚML{�BR��j�9�!%8���+��JmY��HY��FDY�z�5&e͘���V��nG��MZ��]�IW�!Y>�Qڷf�.�:��r�S!8�T�Û[Z�,T������Q5iՃ��q�8�8��"޺�R��"�&b�\�>�&�G���ؑm�ʅd���B�ӊ̼��wt��h����mfXl�d��a�X2�.ŲL5_I4�U�[j+)-%�KZv�9g1�DQ��H�mb��7U��Fk��V���j�]��W��2����-p1^h.j�2�
x�Y�e�ʽ��b���B�,��:Y��6o4��M�h�BxwN跹'r&M$��n��Q�;N�ƫ���"u>�vK���`���P7�d��B�V�4hL��t曠�Ɂӯ��tJƬ�[d�S�J�eSp��2U�֐v�X�i�+)-"[oh`2Q�zC:��Y�f|l��6�UM,.P�^��F4�	hj�R�n5�C�F��B����УF�lڰp44ɘ�GV2ɓ�qYv�(U�bM�)=6�ƕ
�+X�L&�x���e��N��-�^�9Yhe����,�5[�����mY�wh�r��ܥW���[W#�y�1�n���7h��c4D��1=�沍��,/^�*��h��c2�M^�����aR�wu�[e���ۥ!�.��tt��|���o��Fk<�ղ�Ѭ����J#jɼ�y.⫆hj��Wq`�HZC`�T�Zlb��"cpl�l�2�������Wta�p+5��T���e�lؖЅLչ�RK�����p��j�F��B�F�BF	�Ҷr�r
&���¶�����1���.�r:;���r,�śv�Nd�n���:6��u�ո2�,�XC
+k75����DwQz��V�ml0��و��K
��-к��tg�h��1]u@�*��A�1���/R�������S.��ͫe��\T�9�0�����[t�A]��?�Zٵ����yi�M�`�YÖ�2��y�����?���ƈ*J�4V<�Z+4��z�)4,���JGA=�˯��N�m���s*ʩ�-��Ħ�1-�OC��a�W�HL�I	��@�l�t���(lOt&��%��+wu�n��Ծ{4��PUM��L�rf��l�n휐<s$֪G+s&el�z�e��ʩ��^�F��Uz+"���	��.5�
U�hCh�#m��eL�y&�䬸r��#�f�m���o��t��q뤥�x�Z�De��UKE'��i�)����-��
��F�R]��;���8��`.����eW��Gk���~� �B@� ����6\c�2��]��
cl�ˍ�����ap �.ˁq��m��l�c*��p (P�2�lˍ���P���c
ll(�v����.� �l���cq� �]���6ˍ����
m�2�M�l�����`S`��P.�l�e�(l(c.� �2��ce��(lc
`�(2��S0��˔P��e�.�(c.��` �P���\l �lap� \l����\]�e�v���\���`P��)��l)��]����P�˃apce�c
� $��� H�W����+X��~�s��uz���)�k���9hDMl�a��"���wM�&��	���]k/3�*�#��h�x�������u"(��{G�)�2Q���ڕ���Ꝗ�Q��
V�Z�(��Uf}
���������0UcA`U�	�CY��n�3�<��=ݷ�EԣyD6�d[{���_��+yeޡ-L}�3͜�ۗXc�fo�3nQ���Q��.w"C��URW�E�L �<�f	��Q��x�F��KL+3xf��T,b���yB��T3�eg��7#�N��g���{�x�G�ovMŊ�u���\��cŧ3��
�g%��YC��gv�+���W͕��K�b�3���W1l�����X��������-
���1`��W�V	ۡ�i�4�AW�,Ѯ�L�V�l�Bŕk���^`�mc[]��N�]�3S)�꽽��²<R#}m�L��˺��5[���G�ƴoh�5;��_9zcne�Y�`7T,�����;6l�&�"��j�a��`ܜ��J6NwӋ�5���欘wQl�Bj`f���!�3�,�1i�8����0�@�w������7:��a�*(�sN]%.�R+cȇ%����ȸ�6�1�щ���С�E�Iǥ�k5�F�{w�iVN���yr��uu���k����x/#mu��s4�֤ZG#	Ck@�zl �M�;͐��f��W|Av�z�V�x)�Z�Z�ݥ{i���9�QaҤ���_n1G���=��q�����F������WËf�z/�1��w���vJ�ܜB�Sraz%��0�+/jД�mV��.�6ؒE�r���y!�FL�Qi���y]Suf���om
��{�Ԭ���g�z���6���Jd�٬WV )�������S��cJc#��?= �1.�5{�P�c�[��Vl�I����G��ȧ5.j��q��UWk���1m>�cbxQ:�Fu��>�d�ۙy�.f�\VJ�r�E���u�e��XnL�������:��)�#-�'!��*y����PL=�W*YB�-r�]wӦ�Y��f��][CC/v���y���.�{��ڽ'�����`޹�{�6���w��C�b���w�lSKKf���+�T���TI[��:���5Z6�n�����i�P*��u�rپT��C`m�u�-�V����}b�[T�o�GK�18��h�E�ʀ�#��i��nd�a���+'X��"��Ҫf�뻢��;�ҹ�A�ܴw��+`ܺ�uD]�
#����.����6�<���V�z���;Hԫ�ɖA�Z�
��\�:������ؚ�Wb�Xz3�8�.�����K���3���4h�Zy�;Q8���{��>��0U
�7rm�K���ʨ$�y��X�B�U��Q;�ʎd�X��̭�yM�>+v����dҗ�l��შY��7B��GS�UVؐV\�-Ѓ=�mU	y��ne�K�.�a�������*�aɁ<��ܧΒ�[^*XZ�����i&oU)�P�ŝ,��u��i�	�覽�nmMZ��7�L�̏��SL�%!Y�x�n5v���W� Z��ż�a�^���e���YT��-ҡ�;���S�tF;�=ɫ�R��Gr��m�tiخ�k@E���n't�Uk�
<��l:�b9�ePti[HX�����W_Ծ����ޝ�S@�ꁓ��ycv�-4^)s�`��A̎�]y��q}�+����b}Q�<Sӻw`U��ۻ�Wiu���kd1|��HFKwogc�+6���bq��C/.�k��y�ҥnag*4���U�&ҋCs�CQ9Z7���;����e�k�n�S�P�{���͋U�f\(4i�ʱ������f?LU%�X��t���]���\0`U�����ign�iSA���3 o\������w1�}�W�[���b�'-��s$�L�FB��T٪2���̪t���Yr[��}rI�ŝ�k(,ko's��n�7WKO'z$�ʊ��T�p�F��B�W��X�i����e�/p۫�I9�	5�}C/;.�9&T��D0��X��,���h�;���)q)0�a�6R�x�����z���#�Q�J,c7��Y��;�F�Wgq��Ir�5�^Ij�zZ� ���/�ڻ9���K����y�o]�2���W�u6��bZ�Rw�9#�\��o	��1-��M ��%
�W)��tL���.�3Υc�c�ʖN�a��r9I>��n:�d�҄D�^C�VCuY�m|LVcJ�Vּo�'n��b����\X��c�K�bQޤ��EU�f��j\eYM�]�oh���3z��wS3�ʠnۋ�۱G|�5ʬ�f�ks[[�zpb[��']:�b��ZUw��K9�Yx�7�ӵv��BeA�ý��m4�rN/r`���Ү���:�b�����N���:���T��+M�+���k0��^ѹ�EGNh4{$#���eEl��~ܽ��b+O����A��+�UEʎtbo(e^�
����:n����k�i�L�|���z�Puµ>��FYFj��Ѭ�V�s�0��ө"�=�M(p��(�����co�9,�.c[z75*��BΧ:����V����+,T�O}�y��0s�MZ6r=4dݹ�ޟw$+>�l&��*ӱ�Y�V�j-n^p"^�����ُ;+GJ�V��I�<��#-����B
P�A��Z�VUԪ�Z��Ƙ�'�/�1.R�-�ŭ��q�{�Nz��r�'7w`�ӯ�^�����H��\��ͼeM1uX��O�x��;P����̬&u�[20nGbUX�W��f]�����U|�To+N���73�-m�w��Q��. Gr�Gk:�NY]w��	�MU�e�n��'�J�T�d�]]���T�7�F������A�����^ee��v�<ʽ�DC��D�u^��.��81p;i��]P��Q�W���er�u�ؤN����4`�o�a�n
���
�t�䫉�uw[�!�C����ډI��7`��¹��񨫞�����]wH;��Nw"��*w0�oD��J�T�F��Uv�u����J2T۬�ո�L/���T�X«���ˈP���!:)�˜��g�R��uaT��ct����=����r��!f7F��I�d�wxr�O��F�꣸OX+ZŰY��������Ƌ�u�ܖ�}ȹ�����n��}�ܶ�]J5��q��i�3l�!N��T3c��eۅ�͊�]��7����3w~$� �v��83l,�]fe
���n�2&s-*�+���2L�C���×�Me)V�մ����s��U��g#��u�r��ى��gu���� Ի�;{��ڳ*�ɰS�f�n��X0Xo�S�x��J�K�<J�h��Vr��J\�Y3t sJN�e��:û��޺'��3,Z��җ��m�=��T��
VP�I�M����+=�/^.��5̾�1W{EU�jܩ���T��s�����,i=���u+��`��w��Ix�^_Ip�j���7�GXff��"�VfK
Ɋ�B⹺���5��YF^l���hJNQ��۝\���<}ۛD͓�L�\����X2:=��kߛYԭ�ޘJo%*�S9Q81Z�u���Rꋑ4�Kwm��[��,Ȇd���O!˧��2��f:�Z3�5�6���?�XF[gx<ʅ��Gk�pf>�ب�B���i�{g�wZ�k��, �n�P��wH��NWN�0�p�F�ޗ�B"_w�M��F]=��g{�38��v�gu���!cD�wu���5�S�-���H����ST�)�IҪv3!�wjț��xEṶ��7g(]�ō�x*�f��.D�`[�u�E:%C����]���w|lA�_Vn��qe]%g*�C+:�B�VP�M���ӂ�����8ᱚ�n�-<�����EǕ���O�-s+�G1��R��3����R��νJP���]l�
�6�����^���y�O��J�F�L�w��n�n���,�v^��,c��ꁄ�J���*�(i ��ݢr-'!U'�UK�W	a)T��	ӑ�i�QP�pヹYZ�=<�4!�૘�WP�T̋��P��l����V��Q�q�[�ۜ��]\;������Id�hӺ�u.���i�+R�R���NdC�
Q��hP�0ͥ[Z�
us��|z(�y��NŧzȬ�@�\�{��_k܇���4��7d�Ww��͒����0�p꣺1'��P���Ŷ�e__X�=��ޗ�t�q����Hݽ���X��^N�e�U�ӕ�z���d4�Ď��q�R��V(�=�ƫ4�Y�/1���d�]���gU:�ȅб�wj�b���"�5����B��[Q�%md�wO��og\���uL`'r;\Ý��͋B\¹>9Kѩ�F�YHP͍��mζ�?�:a
��`�mˎ�L�v�Iu��]��)�It�tv5i����6ë�8�s-Ⱖ((�MT��X�uU���w�b2����霳��&�����Ծ��6{Qu�I�t��T-6�*��Y��vU��7
��5>y����F�����R��uӮi��\ʢ�*���Y��4|����Xtk���eE(��%�
���@��>�6��6˵�Z��[\NK<F�x��d5�nh�z��a�`L:E�9mU�n��I*�
�w��H�;DrW	J붣{N��洶�\�I)�R98.��՗Uf��3���Ύ�kC.NY��Cqf�}5Q��v+��m��3)-�<�U��_d�ȃ�ue.u�o�Tx�؅d"n���4N���m�R啙Vn��P���X��0N�Z%�]>���h���]�L���z��7=��*�ڹ��V}�.'�2���]�����a�׽6[:V�w@��J���Q�Cffu��M#�� �_�Oo�����yً������tߒPj�V����)[.�[����r5�tVmn,L�#v�ԭC]k��2NG�c{��>�i�ͱ/b��Q5n��*���Wʳ!Cw�;%I��jt�vG�q[���K���3
��[�C.���p^e�$�y�I&�U'�X��oPj���3杗|F&e��-O�Z���[]B�؋�y[u[n�Z����
�^<��g)\��72F�ȳ0��2b�;�ٽi��M����ٸ�۱-��3t��2�)z��b��Y��)%n(�tr��I��#}-�������`6�e^��0ܪ'7N;��8܇h�\.�ǌV;��?]mi�܆�9�����YA�-Z�Z1�iL	��7-�6^�;��U�ӭ�N8P,R*��54nk"u�/C�*_guG�7���b�t�0bYt%e�eDZ&�Y��j��Uv&KՌ��Y�ZֺԇlTlżt��V���a���P�YBr���NQ�l�d�r骽x��k�6�]�	 �$9.8i�U֝)+,�9o'SZ�b0H�ݙ��$i�0X ͫ�ྂ5U�ʹ���#[�{)��e!��v�o��c��L�]ӸXQkCj�JGmi�E[�J��Jf�n�}.�d��W3���E�Oa;�΁�$��=��P�n�<H����x"3AߕQ<�}V!��nf�,]��rd���$�9x�P�a<خ��D�um�rF1[�5��1U�3���9:!
b�9�@b�Yֹq5��e�Y�M�R�O���&�@j�y
.i���_q#-a�T�ohKm	���8n+����H;����7�R�6�\��k�����j����E���v���z�Eh*ȇ��Ŝ[�f�'�Q��x�Eb�X�0q���)űk�Dm
����ۙ�[5�U­��1}b3�r̕\��x�Λ7�<�,�4�6�xǶ{���B��^�j�rE�Qf�C��K"���&;�Y�kO����ψov�k�_n&�귎�;'�&�=�m�n�Snξ�عr����w�*W�5����囷����=g,^���P�`�[``�
3��a�#CvL��[�5W+�5������IO��w�
�S���9����qWv"�wxN�^��b��W0͋�7�({��U9!�j֛�B���&oVێJj�h�3�M�LέΒӓw�Es�<v�e��K�1V�A4��ͳ�b1O3l���s&N���T�����WA2���a�����91e�z��͒-Nz2�l���j��9#�a�yu�Ξ���FYm��F��*�6�+Fu�yF�:ѕ�R<����[�*�X�q���1`.+/M豋A| wT]�O�Y�A�n��M��鄥B�[-�-�����y[ӶnVa�X��!�p5t*��6�6���b��S)޺��966�1l��1U��
�6�;L�@�ڗ�^��ڭ�����"UYE�n��:g`�w6�Q%\˾�c']��x��nnS�yMkbC����*�k�K�y,�h�Bu,��z�6���Ī�(�UE�g�h�˪��;.��m,�-�1woUQMP��fKٺ2��X����v)�N�Uo)�t`�;Gc��9�����	��G�JM3�۪�W%���a8j���'Mus����Х���j}�2�]�+������g�L֒��7��Dܭ/��6�7�Yd.ϒ����k*��	�>缪�����P�^�����i�[1�o�7E�+͛S�K��ݒxV+F	Ԟ���S�sPb�uE�X�I��1�雗z�E�X�}Bgb޷���~5��J�3�h���-v\HJ#{ejm�V���Ú%��3-������U��(�r��޷�����^:O�^�ʺ��y�:'^=�L�:�0�l����*�1�{|J��9�Y?M71���d�G�l�ّdm���m��IYH=˸�4���V!�e����͎��72�[�����e�\�^v]�۫����Ӻ�Q*��SܝQN�i�S']S���.�E���Iw$�}}���U��[�䡛�B�Ĳ#�(�(X��J�ءH&e:�5t�)��1����4cDJ�J{J/�ESW�n��ʽ��md9��� ��|;�N�I���~���`f[�ȸ,�kr�Kt���m]Y�\ՠ��;V4�i�X�iF�f/Y�e�Z�P.6�h쑍�&-0�Y��Bɖ��1Z�������&���Gb�`ۭ�hHD��^��׋�.��X�p���{6P���?��y��b���a�I�U�V�T��)L-�5��M�J�w��%��1:Ź��ݰil0)TB�-h�in;g�52B���^񺇈����p��5�0�l�b[z⸃�s�J\+w�4��	��:MQo����X�d�f���&66[�E.�mn�h+0X29n��ˊW����Ǟ]n<�\�L+��������,�bᔱ�"����!sL��f�m�"M٤�鵫#
��-�r������11y���Ȅo�l����SͬVJ�F�{bZ����f7Q�r�M2��Ҵ�J�ᆽt���)�Q�Y��Ԙz�[kl[�=2�ًhB��e�ZF3rMuFa����֋�(X�k&����-��c�\�Db���0eG�F�FĚ�hũ��n	��4\j�6]ckP�k�@�X�K�8YM4c����V��͘���!��*RP�ʗF�\���V;��h�dS���9�bJ1ι�ֲ���]����fVX�s�GJ�U��5�a��%IV�G[liu�9� �X���i�VWCBT�u9����յ�u�*2�A#M�����]�!���Њ˭R�Tm�1��� �t�`�qh.�o*[���ÍbA6�� ��\���k�K�奁B�,mi0٢ͪ̍�^ٙ{2����K#�.xD�t�uѻ&X ��؁��aGLqIgU�m04��GFʮnj ���5�����cUY���9I��j�е��Cf�W�ill���E]�	��ֱc���Ku�k2��Ő�ڹ�u�D(�t�����4q���l��M�ԕZb^-WJJA6!H���u�pmy��q�՚�����-)RKm+�Tl�gJA�d�j�n)V�H���M�D%�[c[�ĪMn��4��qb���m�2�SJ;��4�S����Ԩ�
� fH԰+�	����!ԙZQɢ��V��y�gv��bUq]�B��r^��b��X�e�j��Ҫt��6�H��Lk�Y�X�]"k/M�Bᄻ#Hb��]b��2c���v�0��D�Wf�HMP�Y�m�a�YT��l�	�8֤GMDդ Z��[KF��" m�"]S^,�+��%�G;Y�xX�+��G�Iq��Q�G2;M#T�к�����5v*V1����U�B\ĕ�h��I�<�Y�aC@�nn�FcP��]��bl+���[vpc��m��F��c����t#�P�mr��Y��&�J:`#6���ZT,#�3r��%���XSI`�l[3�ͪ@DK�b�T��f�����SV�b$�vٳ,.CG�t�%�R^,�Z��at��<�m˨7\\h�]�I�FZ��WP�	ڵ�Ѧ�je
��ZP6�^_<���j#6���v�ݫ�`��sf�Z��d��*Lu�QVř��\�6���k�t�O<�����y�*\��u��c�����:S���D��k�f�m��4c���3q�Z@�q��ȶ%��]`L�sQF=� ���;Y���R���h1�L���\Gf�e��10:��]���s���+�-ۖ.�o)����V&i��4R�M��nT�s�X����ͧ�kl|��,KfQ�^f�mL�΄�l�f��CLY��ګ ]K��4a6���Shsq�CSmc��[�Pv�t��BfS���78(���Ě���Vl�Yv����G9ck��%��Kf�۳�0�Y�`@얁����ˍ槔�M��;pk3*��8 �����e�"j2��A�a6K����6��R�LQ����k�Di��̦%cW���Bհ݌�����	t+laB�-��Pcµ�����;Kn�f�7��v�)�r�Z�:���U�<c����Tլ�SkmF�2̡��e���W� ��s.ce�����lش�ʹZ�9B�j6�8�ZJ�u����j9ƌ2��f�]�M5&���4y�pCimq��BѲѥ��01��c��̶�3��g��L�`��ļw36Rc-��p�{qL�M�aWU�!��m��3�.��C�ӭn+Mt�k�M��$�%%��K*M)�⮛&�Ў4eҨ:$�d�ۉ��m&�Ì�Jq"�m�9��3)C]^�Mر ���vJ=�^F�*���8�A��u�G5V�h�)�n���&44�U��͑!m�1��؄s�4h��ml�4�U�43�3E����^!-�'Xk�Xr�ۘ�����m���n3 �Kmj�j���5eS��X��f܃�e����E�[
��P��DJk��1��-ڌ2���.5��n�:%�*M�����4،!4`�ؖ�@�tƴ�f[e��#�$.�J]LY���U
��Yfp݋�͵��e�+
)�e��M���+��1y�b!�.���cZ�.FF'l�-��`Z��]1�)hD�ڀ��4-�f��a��d,%���V��Δ�[t�*`�J�m*�hѬ,�&�IHcFP��,�v�6����#��'\j�fZ��6��i4H��k�*����Ba��,&%�[\�� �5��Mw
�J�#FmR���ZْmW@$	�7ac	qWP��fZ�����4��ba#&L�q66���T��8/8�DcE�Ā���(�3n�]b�t+kn�eĵ�զ!se�b����n��X-��(�d��F&]�I��Ţu�ĉ��I��+
]�p$v�L���l+���6f�1�60��d[J���(󋅱1�m�)������L��1*�0�.6�q^�m�eʹ�:d[,�G5�#��G^G�c�ui�d�X�K2�هka���
�ҭR)�K5
-��k��a�)�s��w=y�iJG���:�l#0�	�n����,�a͠m{L�5Q��Ia(j�Fͭ��<�1amԥ���,�k�b�Q��TL��6�tpR��� R�-�\X�&��4u\Ԇ��&P��ɮ�1PhV���L�F�T�%��g!c�G�0dݛF+�U���,t���F����ٖ�a]a����C�<�]M�m�3��*�&�V�l6,��!Qr
�sjY�;F�ѺT�Ə.,���a �6�jL#+�D�b������u�Ŭ�˅k�c1�.�\���e) &3Fh�'2�\��YB�Wb�4+R��E��ҽe.�^aj1�i�� �K�Ff�`��hQ֙f5�`�踀h�4�[�r�j���N����keGJ�a�9���0̌�IdPu�f�֫�-HQ�b�+]4�]b@u-��%��I�T��J���a�t[f��4��]��L����2Ѳ�Fb#�1�M	��t�f��+��AV;
��(fٮ�,
GF���+o��l�֔�-���R����_<t���lX�W.(�����#��*K�nq5�L��	,#��97,�J�]+)��M7��b3����lee1��їV�/5�m)%Ik���"�,�`����sa6��ZX� ��
Qѡ�[����0)t�X��6�Z���n,����C�C��DN�+w4�B������.�+J��L�
\K[���ͦ�Gk�T�G�Klm3-�q�IH���F�Һ(�T��^�
A"�41�mV<8k^HJ���2��n���r�ڊ5J��\�bg�k��¦�aU�//66��͒jf�5fk0�D�Y^�7��k�Y�#�it�L`ʬ�jn��]��Q�l�rP�:�k\��j@0+�	�*EY�˓M�m:�!�s�0���D]�cq2َ�dڢK�pǬ�0��F�FՋBY3�T�.�h�́v!�����3Fe7K�Q��&Յ��ͼ��,dkae�R%G��zm�E�Z��c\�m!LbZV٥0hPm�,6�����ͬ�"�Y�4t�5��%#k�m	p�ň2��s ��u�c�+t�v�Kk���sH�̒�h0��[�]gE�u�*�]-yT-�D,ae�ueZ䲅�� ˢ�F��e�T������ɰM�[���+t�&�$�t�V� ��|��0����^�U�j�r2��Ԗ`�hDښ��iQ���R��R�Y��u6�FY��pɨv]-��%)t�"���*�up�E��M,v��Fi�>K�y5̲�1�,�,mڱ�1�,-������(�A"U��9Y�;��*-�[30�40�J0�q�ce���Ckv��*�`����0õ�+Im2����Ag[&KH��]�k�cj�8����R��Q��1�m�h;U��5K����<�,��r$Q��h]�h�j0%�c��`�[�r����͈��ݕ�e�"�˭��jX�v����2љ�,�j-�.�°M`$@Z��,�c9���r��am˙����.z�:�,D�ܶ�Ki`Yf�R&�z��Y����n#\ƺ;���aJ�X8.Ж��&R	jYq^�y�&2L˓K@��yn˗r�g8�vՆ�����lw2�]���ԩs��v��]�uB��Hf�0�3���rl�T�Ѵ
 cr\����ya�D�u&��UF]�\��j�[y�2�uH�t�ڣ̋��E(b�e@�M4kjb��0�-.ФJ�dq�.�.ڲ���˭[��2����#kb��S]h&)��ٚ��J���\�t@���Uц�LhͲ�\�L���p2�Զ��VR���:\�J1;b�&v���gJMtMm��n�il�@�8,c�LE�MBҎa��b����5F���4����SFUX:�ţS\�:�,��T,c���3�CjF����k+E��#�f��b�ea��x��U��i�l���l�pBֶm��w�ǒ����$��vK�:�[y�mn��D���+�l�`�ذҭ�VP��O<P��|A��WM�[��4�c�Ih�W�ƫ/�rB�3�J�*��<��\�Knwv��TC$��DQv�i�Xr��;r*��\��äē���Zz�]<��҂�J���rH#��'R��t$�WfdE+EY�d	2�L��q,Σ.9�!:�:���Ң�Ԣc�z��ɛZBK�sҪʓ�ȧwt����y�+�ZȊ��P�N&���9SID���A"�ˮ�����p��UL�-b�Ӥ��h�S*�D�ʪ�N�HHm"� �s���Ĉ�e�v����99�����d�H5+����r�%np��H)<�s���PF�ۑ���]PӲ(����E9�����W�^��L�-b�if'B(=�p�Γ���(��b�EN���AÕ�-PZ��M��t+�9:��WO'9NZGiN�$�G���i��Eյt��"g���lmc��l���ZYq^�2d���Ņ�rfYM��v�u6fG���R�R:�[���GŌ�X���i��!q� ɵ9.6J��Q�r;�m6sn�T4�.��n��J@��:��ƛ<��R�m�v]B��Kqf���@�*Յ�L]2���aF��� ��mb`,@��q�[n���R��0���պ�^������V7-БV�l`RW3ظ�"T�͝�.��9��.���ZU�d�^��n ���ڎ4͑�V�Z1왛Y�f�$d�V(�
5bA�����B��T�`CSC����[��)2mR��Q��Rf�c/\�hu�e�:4}�n<!g�3m��J�l�X�l]�f�v�Ia�%�e�rB�1J'RR�-R��.c��X�F�;�YSR���٥s�t�klM`��VXrP��F�3ۛ�lʺ	Ǝ�i�@I�YYq�a6k��1�]+X����U�	�Ҙ��n�,Z�av����z�K�c6kCL��iS���l�����֊vF(͐N�͋0�b�!e��hMe�]r9*ؗ����b:�F��.�n	7])A�)��u�Lj�Sh��k
�V�XȀg������j��T�5)���cc��9VhKf�T��+a5ulC�vȼPr&�\;G9�D-�,[M�s�,�ղ��k�6+*��X�6��7��fd,�H�&��Q��	�4X=�W:���G���cu�	n�k��h�KK��e�Ux`��Z��e��J��a�)�0sm�X�Vlo.��b��L[�K�-ɮ� F�.k���Ym�����gVfl�9�h�Srf!*=b����ѕEbSke��;Zk��:��JXj0#!�e ŋu�/`���K�CF]�5i��3&�͈R����v��4lK�[-�ˌV��U�i�WL�d.�1ۺI#6@�liZA 5�	���-���Ж��h�V�m�
@Z��GYKJ������H�¬�ӭ��(�jዔ^�0�qͭ���R�%�F��V4�X �eJ�cz�����E��-UU����­8�5�^,��aHǚ�b ���� �4�-�jz�������	HV�2��V�,�5`���׬A.srk2�z�!�2��� y��@����W�H��Wb��&U���_0Iꆶ��9�.���H�O�ȟ$�QJ$�BQ ����+�Q����FbdD�b_��x�J\6�0ޠA� Ij<���w���A@��}{3�}5�
R$�)�J�\ݬv/��i��\qL�4�m�8�Ԋ(�Q$$��w�f���� �s`���n��;ا���u�δ�{ޟv���9��~hO�IТ�H��%B�J�Gts����[�ȧ��K��&{�6�O��?�� �jsY�g�y�2�	�{f��Y��1A\����Z$K�,�+�@�mT��7҄y�/DG�e�׬���4N�z�Ε]�[m�8�D\Q9P2�DeT�Px�PTzAE$�P �H��5�g]:�Uتj��4E��)�HDl�'G�SS�Ө��;�˾�D�����L�g԰^+�p�a^'Z+�l����~]n���n�%�s�eC���#&�<���뤫vq�,���>�܉!q�U2q]E�����ԨQ]A�>:Y���� �:z�������u�S]���co=�@�P$�Q�J}�H�p��O�8�MG)g����yƗX��*�"�n1��,ψ7�8�q��p�yĐAe!%U�	u}��(f�fҎB�<x+ؽ���IV��Oװ8���ǂV'��*Ŋ]��;�/��-�4E0~d�)�w9���h6B�S7fR���Ma��Q����Y���T(�|A!(����T�p��x�	�P���-�Q���>�%O��%%>�ۃ6c1�����S�^=:ZY���E��c�� S� �jE��!%n���	Q^#o$QJ��R�%%4BQ����uNr1����sK�(�>�u�������͎�ut�W1]�弚�j]��\�&��j�Ƚ�U�`R,<��#�gz���w��6V�z��%[��?^�v���ȓ�|��%���K��\h͋3
\H ���v�-�S��k8m�`kޠ|oP`�����ݘ�f�HgǶ:����L�RS@R�>>KI��<W��%��E�*�m7��I�^)C �7R�)O�tԭ6	U|Hh�Gc&�p��l3.e�c��Wj�)@�k��f�F���R8�	�:�H))����r]�-�꤫vq���9��)ox�9W7��$O��O���$�QJ$�BQ���=�a��ŐX7 �G�����u��2��^k^�z�	 ��	�IJl�\w*�w�H�}�3��%	G��*uU���p��cR̊��r"�n1�)Ă1��I�!%"k�2J���U��W� �$�S�JFE���[��IR�ƻ�zy�>�6eu��j���zp����#Ddc�O���3R��ZÑ��ǣF�Lc]��]����e+��Me݄N���tXs��^���ʅ�I��H)*�D��N)�X"�$[yjj��;7�o^��P$|Z�%%5�n���0e-��
�,R�UZ�IFb:n<� ��٣/���qX]5��s�U	���p�Nv�x��|���IP�\�j�S*�E6�c�#�(�t*������q�%	*�|R� ��E�R��T+�h��2n�Υ��T�-���{�A���AjD��#39}Ͻ��ut(�@!�H ��QJ$�BP�
b�D������Slm�`kޠ|mG�P,��%"A�R$;��p�eG9���>IO�:՝�'y�!��{�Etz]����7"�:�E�V����$$�P ��'u�;���My{)'�P�J����ΪZ�g5�^t�oM� %"|BJ��͈�2;Y�� �[�P��j��>�!rmuk���sǠ��������'] RK_b**[��/ ��ެYZ�J�G�H��ڦ�t(���&d���1q���m�WRTå(�DKqq-�ŋ���ʺ�53)�LhQ�ۖ\�$�;��^�1��2���l�������t�&1mW��,R�6ej�VW6�W�c��݈���W�v���v
L��B��.�BKlJ�.�lqXǁ� K��Q�8�
BC\���!(��!aq���)�WL�.����T-lج��3ce��|�=bh��Y��SZũ�0��3)��q ��
J��A*�R��f�� ^'�<��� ��Hx��E���nc`kޯZʟY�thDs�X�DN�ˌ�l����&��fs	�ѓϷ�O��t+�օ�b��-��$WD�%B�J:���tͧ�kA5��8%(RSD�H��x)�9�OVuR�{9�����D5"O���JE�O�!ܧjM
��.�x�H>%᷁�T_q{7�s^�Z� ��],䧣��X#\	 �)�$��>JD�|�S/7�WI���mx�]�rX����q� �]F%"�J'�BQ]2�mgv���q/�}al��h�U�iK�JqcY�2։H;f6�Q	pUٙX�~0���4!ǿ�cߵ4A�R'&lwm-�ꥪ�s[��zE&���C�@��>�	�IW�� ������r0����O�\��3����x��X�T�/L�g���7�3"?!b�B����l������.����90$MN^\�c�{5�s^w�j�	j�RS��AD�ݙ.�D����sz}^J|�>)*���:�`�n��9�g�X�\���q�EtI�@�@J<������@�|ZS^ ���3a�����z��5�ft�{�@���:��j*|�>��P)D�A	D��U�SuF���dbʃՕ1��u�s;����6�H>j��� ��nWT߫�ų�>�� D61�Lh��K�2�b˴am��k�\�Z�&������~�:Yg߬o|�3�T* ��Tc���z�c�t��5�Nen�ClkVA��P;ɐH�L���P$���y@���]���3&lwm-�W�ns[�g	��R$-ݴ3~J���ʤ�@�_0D��;�B��L�F����y6!��s��㥙��1�o��Z>���R��f��9Z�q6���V�0Kvn쇃fF�c"D���zM�BZW�F�Ә�	�P �� KQ��	@�%#�.x`M��!�y��0~��㻴(${bQf3�({M���+�A,��֡�bΨ�q>!%@P>)@�	J�����Μ��v�� mO��,�U�ns[�g	��M �O���JE���k�tz��ᡤAj�
)6&�����[,:�l&�C.�Ĥ]�1��d���>��Y���B�B�J$�BQ#۝����i����l��7V����F�"	�� ��JD�%>�$��F%w(vP��&3�ڛ��:� ��7W<n�᫥w=��~"�'��B�Q��������i�Ex� �R� �׈>J}����G���ڬ[s�߳8O���k�'�G�%�(�ȯR(�Ni�ˀ#'?�V|A�	D�v���6��ˍ��O:�/ O��,Ʉ;N:!2#k��&�ӱW��p�����Z��b4:xh~�#Y��M��o3f�aBكnOFQ&u��H��� h=�h��I�R$��	@��l�����P�@��R�&o������+�A�E�H$%����|���`�!WĖ
	PN�H��kZ%�����6��f�%��_�����=|�{�u������9�r��o�,۬����}&�%9�
*!=��ȓ��||��E(��		D�1������t��wc�Bq#q�|7j�뽛l�����)��dt^M]E�7'��y�+�%O��>!%As�J�1�N5+.f��Z�YAWD��T(�H	D���P'j�F�,��o'`X �n�^���9�r�ko��ٽ����gM }�0z�hD:����|ڑ^)D�Q$�
(w���l��c� D�J��z��5�y6�	�
��A-@��� �)	�Cnc'b3T��� �t[�H^c4��R��6]�Bu��W��42sw뽬�F�4=ہ
�Hu�S�����k8fne��C���#IMc(�v�z͒�vu�]�r���1�:6�P�� �Tr�+��T&#Zi��WW���FU�U�6�,�{ �����@.,�X!�������ƭ0�Ƭ)Ԉ��6;ii)�J�Y�fn�2u���s�e%�&���Df%�`�Ql�kAu�Z�Ʋ��+��^�ƶWQ��gg"4�lD6�ti
2����L����'�|�5�T̪T�l	|���,�jW[���̹��
��]��г3����^�3ݲ����w��B4�f�wQ5���t�8�(��J�e�`9A
�j$�BQ ��
�H>{���,�В��M�Ȝ����,�՛W�߲�O�t��I�Z4�w�Ft�ud��8�G(���P)D�����3B^͞B�v��꼚l�^@Z�%%4)O�W#&!'�g2�[�A���~�����\��tz��z�YA"�$M�8hqԡm>��Ȓ	�>!%U�H ��	�INtv����w8,
P'���^4��V*����ސJΚ�|�X	*sU�����~���*®��ABʦ��lһ��qAH�b��.C[a���,V��w�!	���!oP�R�� ���E���mc꼚l�z]�*�H���@�	�J�4 %"A�R$
Jh���\���˽��f�>�u��ϖWt��խ�/U1���5W��JWO���u9T�]M�ܼ�[PQ��w���pU�a���2����=)��ܹ�n2�U�j�����EtH �
Q��Hr��J$�P�A�A�JJh�R.�[=v"�f�ܬik�x��[�_H&�M5ǂQ�IP�R�"��3��#\��>��		D���}����^M6u��=�3���TQt�����Ma�%"A�Ԧ� �"@>JÕ{{��5髪S�i��E[�Sv�8|Et{51�u0A �ԯ�eFo%�8G�9E͉��u.ٹr;\��c�Gn�% ���4�Ya:j]�uz/��h^��E��oB=�ќ�z�[��ڽ����,��Z��9+ɡ�R$��ψIW�� ��O�G ���|�κ��+�6$�G(��^����y4��G�$��RR��Z��e������g��k����O�J���ŷ�i�G.��n4��֫6��eF1�&�J�U�����Y�uYKMoY�簗�����ˮ�����\q�ڮ�^��2y=i��DEH���l���Ֆ������z���i8k-���<,ŷ�Y�y8�>c���܂�i�8^șn�u�TXc��u��#\�Q�ti&��)�i�y��ژ�a�"��ߨ�Ѣ�c'1�
�m跙�"�{��j�L�{3m���O+]�V5��5���W��SǮeR��y��V����dۻ�
���g:�*�]���7�Ռ�-�v���y�9�7^TTJmH*V���B���L��T�&�mdݠ�e8ʹӫ�%[�LŹ�5W��SSV*Vj�Ǎ�ɡ
�,��O,V�ݪ���R�Xu5a�{�q�X�k�2K%}�+d��14�S鮺�	���ͭ��X��eD�5��̭c�^v�f���)����!�@n��WrU�T��a����W�X��)qʳw������O�a�y�o��9n����֍uu��\�_�'gTRd�Y�xgR7�G'�3�~�q���=t�����F	{�cQ��w''GrẼ��5{Y��92<B������_>JiZ�97�4�q&pŪ0��J��&�Z�*��Kb�grڰ\�����{UYH���+
�W�x],�`���Uڎ,��Mn��f`�FY��Q��g_�ڮV3CcjJmm����ux�+[7D^j#5�^D,��{G��.�#����j2�p��v-�� ��7RUл�ݦ���L�^X�Ld��*�b�2A��� �.:DD�"�ekT��Ny��.x���Q��lJ�*4�OB��M�t�4eeE&��L䨙�T��\ue]�]�;u
�\��
e$���SN��z҈=�X]�L�#�؄�F�B8���Rp�*����ܓ�r��Br�E�X"��'%A<�֑q�&\�;#��ny�.����$����@����9*�UT�k+�vs�;=e7/F'+0)���4$��t�Eq*Adr����h�a�Z�(N®�ˌ.!�8�q:B�q�]8�s[� ��aDr��\nI1u�����ʹARBDWC�ES�I�'qI��
�Bu�2e��!ɖ��t�U��PE2���W�T8�$�s��䳇��99�'&D�U�2$�L���47n�\��
����~�E���I ����RNw5�Re�HRAH+�p- ��a�v�R/^�f�����]�Q
H-����0Ͻp�AH(m�4�Xh������o���^��È�$��>>G�#�a���I �W/�f�e��k>�ܽ�\��A`i����p55D�����I����-4�I�2R�\CI) ������
A@̢�t�mz�H,��_n�Z��{�����k|�w��H,;��;H)
�ܢ��!I����i4�L32�m��
̣I��}������_�g�=�S��J5���t�l��qd�r)���ӴZ�Y�m��k5�U�п�=��~��AIQ
a�z�M�RA@���H,4�W2�ZAH:�fe�i6%n��~��.��Sx �$��I���\��4����bJH,(���6�Xn0���I��$Je.e��D���3,7��@fQiE�����y��h���H)��L;�\4�R
�Q���Cz�}WrK�k^��È�$��>>H)��높
A@���AH)s.����������)����c�=��) ��J_z�Z�) ��35�Re�Q
H,��\ˁh�{�j��s9O�Lt���sX�rm1�$x�$���@{�ZAԢ�Z
��H)��fe�L��I
3(�Aa��$̰�$�}��}�}��Xs�p�'�) �{�ZA`j4�W޸��
A��f\6�]�y�Z�3>��cT���	#��L�J]�p- ������ٮ_��[6���n���\'tF�ܚ���c
�Yw���9��h�|�We����2��^�����8�X2ͼR{ᤂ��?v�I��$JS�T@�JH,32�n�
B��̢�
AH.�ˁ���@��p��`}s���s�-��y��b�W�w���<�\ �̸B����<	�IH s��uG`��s��2fJ��A+4f2�Iz�v#���]֒�fҀ��YSv*�� sTZr�YL��TCBJH,(��P�AH(�ZAO}��[�$X�|��s]��nM���H,=��H)پ}����0
��R
Ay��H)�
a���L�d����E�RAs*���3.d�) �n��.��9y��s��H) ��@� ��w��l�oҒ��љ�}��Sx �$��) ��)��@�5RAa]�jH,60��-&��e��gC%������) ��e���AH(�- ���TH)�f\4�) �B�i ��o[�++���m�}�\�.��V毼8�k��I�|�0��\4�R
���$�H.e@֨��j����d`Rp$� #��?�������q4�gW�I�����JH,9�\4�Xm� }��R&�Ne@��~����s���׾�����i!R�r�H) �����>���5���
| S���L��I
C>�I��
H.e�H)(B�fe�L�e$
̳I �2�w���m׽����|AH<�k�p�Ak����;2��̊���@`Ix�O�2S��hhII��jH,60��-&��Y*2�ʁh�}1hݹ,\k�O��%��A���n͢b9���i6��xH�t��kU���y)֫N��i�h���|��9�g�6��(T�`L6���3B�&���n;)STö�K[�7-��e܂���6m�Y�q���3Q l���P��cKvvQ�f1�&�.sK*0�[��	�V5�aP���J�рʗ6ØZMH˔Ը4ua�2Ģ%�4Jr��hر����6�:�J-�KJR�Ytr
��hb�:y��gX736�Ζ�[4��f"k�#Fe��to��o�}%f-���Ulэ)�6c[���+�2B8�SM�\��i������v�R*�勤��!I��j�ЁL32�m��
!���'¯�/���R�[�;����<	5�0�AI���w�o�~>�|��+���up�'�) �w�- �4�A^����R̸m �`Re�R42R�\C@$��Õ�?p�j�z�^C)���i
H,��_z�Z��s�=����~����ߏ� ��\4�RU�QiAD) �]�@�����3.f�t�z�֙�p�H(\C]�I���W��44�RP�0�p�&�I�,�A`i����F���jG�n|,�r�Ǘ1*f���N>����3��;�->@���d�����4$��»��6�XlaH�ZM!I��R�\@�RAa����
B���_����E��
H-��
j S�ˆ����
d	#�����}��Y������8�O\����Xo;p�'̤���5�Փe}o��H+���
Aa���I �fQi�
H,���2�ZII���m ��3(�����ܭᜯg{��1 �ޮ��S�d�n}�k��$x��$��
B���(���!Is.���3.g) �B�i �߽������s�?�p�ms�(� Wj�c*�plͳ�+3��*��lQT&���Y�����) ����i���H(}�i �44�W2�kTAH4T32ᴂ�J/�_�ՑV�7�l	#���L�=�0���z옻ˁi �����6�XlaH}E�Ѕ$Je.e��D���3.H)�@fQi ����}�n�t{���Y���k��� �8w��q�MΎ���ո"41h7��f+#�Lk&�r����LŸ����CrHI��v�մ昗y57o*����S�0�e�L�%$ ���O����}����V�nb�È��݇�4�R�e�L�e$
;�4�XH+�p2���s��ҡ߾�m �`Rޢ�Q�)���\H)����6�Xm� fQi4!I��K�p-����q�ُ��ӗ�2�p�;i��|9���AH}T�E�J!I���H)�
a��3l��P3(���C
H+�a�H)5���v�g9��u�=���:�H(w,�A`i����Z�
A��f\6�]�]�~�o��������Ϡ~@�(���)��\CI) �֯����[���!���P9�-'D) �P2�޸��JH,32�n�
A@̢��!I��5�
i�fe�L�o~��>�dĂ����4�Xk/���߽���٭������$����A
a��i ����H) �e��5D�R�����{W�����w�=�e���L��A4C,��!7@��Du��S0͗c6챺�*����m��-[0���I'����z2R����4$��}�����q� fQi4�$������w�+3�3ᶾG�>��������7���- ��W���SH�;�3`�I
C2�$��W2��a���Xfe�I �n�����{}��$�H+�\j�)����ᴂ������g��&�O��	#� �<	�x�K�����G{������-&s]_�z����f�H,�K�\@�RAa�ܸi �7T��H:��Z+3P- ��
a��3l��P��4�Xe_i���s�/��lɡ�Cm��N��˪lڼ����7B���9#pYF�s��۰�٣���B��¾u�/Z��*���b�`�v��F�J7W*��u���ͬ�[�9˲����~���A_n��0�AIHS�e�L�����_e�H,4�W2�kTAH4T32ᴂ�`Re���YϷ��W�ϻ&/۸��) ���{P�Aa�����
Ag�A-π� ��x��EfvG�v���H��3��
B����- �Q�]�lT�\l_����J�RS@�� �##+K��S�B�v�e�fq�v�'y����n�R�B՛��t�U�Ĕ8E(�J�4��[R�hF�f���-#��
��#RiPЊ�J��f��U/P ��$S� ����MGf˾S�t:�Y���w�L]f�S\��ܠE�xr�_�T(�H$%Fo���3��l"Q+1�|"�G�\[#�^@�	�A��J2�KE���񼅱�g칐A�sD�H�O��%B�ӌ}�%���Q���<2n���2<%�wU
(���O�IUy�K�2�h �p$���R$T<�w��P�^k�A�sDk=�אp�YW{y��+x�tg�6�L���I�R���F�k�F}��k|���:��7\��CD�En�kQ�Q�����:�$swv��ϳF��j�(�
J���'팏�tU0}M3��j��p͵�-ޠK�A)@�RSD_�������o5Q�E��jf�:eu"�Mp�^j6k2��X@�E��v����e�{��� �(�JFl����#Um[w�}M�*�[>@,���Š�;}B��O�!(�K
P$����R�t��5����4�<k��-��~s���>����푗�)��]{r3�F�H ��P(�HJY�N���Tid�s�f����\ ��H))�%"O��!���y���c� ��zBJ�Ƴa3Ū����܎/�@#WvY��C��"'�V	��Z���G��������2��7Kht����}'x�K2�_���m��w�I�R'�$�]OmV(��mR����{�c�;�S�w+k��Ӯs�b�TWK�����.�{T�M��YC]��*�~+D�Q�n�yN4S�����LL �Y�5Y��SMc�h�GX�a![W���]f���,/m(�G��d���K+�]��kW2c��F���K Ѹ��F5J��fB!Ld��$Gn4ғBE�4�n�煶������]��oC1��\14a��Zsn�`J�\��(&q6�c[�W=]�EI���a,����k��W��E�˩�
\��D��J�WW2�W��~���cAk�t{h���C�*G	h��Β�� 9�R)�$�x�� ���wm
;��H��8�踼u�7mpvC��x�&� q�_9�
R$�)�⒚!����J�kA�
�'��F�������k#����U�l<�����90����JP��O�JhR�r����׫_d˺�wWi�^k�@6��zD��)����QJ$5��)>���cQ� �N�x�A%���w8�8nZ��P �� ���z�H�hs/@�=e��l�{�ޑ���ȪI��d9	N,����UO6S�����M�Gu?�$n�����z��잙�ϟ
�9�!i\h�B�L��h��[�M�����&�*���C�߽������$�!)*-뻅۽�Kw���焉�Li}��Y(R'��ǥ%B�Q��	D�K�9�ʸ�N��f�jݢ�}�ݢ�l���!�p�ꡅ%K���2�-+/��y;��ם�����۱U��y9fP�=
m ���u3:�p���=k�|_D�����U�)�;��w��AyA�Q䔔�1}n���}}2<�� ��H>J=)*
��!�w�,4D�<�)���/�Ӻ�QJ<��	)���]]�3҄\ ��NwM�>�Ǯ�Mvwm�F'�=���F*&�ͻ�A�����"�J$�J'�$��F�#�r�g#D��q<�:�U�9�;���>W�|�	))�%#/̸�t���8�U"U�y#)�$
��q�*�Wn���sեb���R��w��ݚ �ԉ�G�R0��U�����5C����q���a�0�=~�Thy�b)����{�{�.%::��	�W���:<A�MFv��5}�������mt�#z<����"��o�×P�WD�		Đ|��E(�BQC�.�̓g����l�T�9�)yȸ'u::�l5U]>�V_v��W�1[?'����cc��F���Q\�u;u���  {2hcqQy��c-ps�@���$Z� ���J��)�'w2뤞�n��d���`?������9��,�P��q��FVc�U`箷�tyʖ	̫���F�=�"=����*����ة��ڵ�}��{����6�}[�����JGT�;,��U�x>�鮌M�]JK�\LGQ��#YB����MKVR���	a���=��g��Yf.�@��		D�z5�T^8���\ܟmy�C'"z�:��}�@/T� �� �)	IM5��2�(�:�s��V�}�8�$�U|�A#�}�XϊQ��ɋ��!(��S�P0JQ��)H<��CNvo^c�Z�4�#[�>�]>�R'��H���C�(�Fl�>S6�����B��� �����1�L^8����|�8P ہ ���yW��n�9<秉�P��+��Rg��zPShN�V�U��1�u$����l�u�a)�1���×]�7`ykw,�`U��Ҵ�ZJ4?�  7��>���#���w�X��o@��l�w��G��	T��\��N*�q�ؐ9���|A!(�p�LL����R�)�X8%��iK��	J�/7�Q�č	��R�hV�I�(*�*��9d����#u
9�^c��~T�#[��6�bf�Aڷ��A��%���2/���gWq��A(�{�A�#�]��7�-e���3�P?� ��/����D3����?y Og�|D�3�A}$a�z�D�j>�V��̓yU���a@����` �
I*��w�o����ID,M�9�wdMFrW��}ȅO25���wܽ�Wf���~43�B�s�ѦD� B��1FE1�k�yl�!7�}Fs;�nr��%�@�n�K"�٠#vA�u�r�I�g0Q�JY9wU���=��1B>�4�'j#�@�S��)�mZN�Fyn3U�*�f�N@�m�V��BQ2���+���5�[��jؤb{NJ
"T�1Aԍ7N2��I�:����;"��k�yw\�.s	���kg���+�ʳ4�+�V8 �%n�3$ڼn�\�H�Yi����s91;]��*��wsv�w�E��f�&��pݫWdC����9�8aF�X/����-��&��w���lC���;[Ad�Bv��UY)v�|������MEg���=N�K��g���N�/+i<ԜV�Yɠ��Hgz�u�T�O��/.�Vha�6�pݿb�wM�ʨ��ۓ"��H+2�>Y�ݽ�k�7ܳԪ�G����W��4ꔫỊ�M��99�ODҊ]n��oy��;X���Q&1t����e=�h�]������J{pH�*�����M��){��J;�t/�gJ�=a��GeFenVJu��������|�N⻫�g#�����\�M�8v��%��4�����K���x3�^<4sR�r�Bz���p����Z*c-����LfV��:���p_U�"{������R�Ki.���gV�1]+�����
xҨڹ�U6����SZt�XrS�`ܼ&��M�y�]�Ik�q���B���Y܍�WWN��̳b�N���Ma�UW�Ɛ�U¢�aw9u��yу{C]��mAu�fZI�5)�$vb���%#0d�p�S���"3Z/����Ce�p���)�U�j�j��e\�h�\#���wp�G&�m�[J��������G'6瓑AE�-��Μ��L(���G�iP\���ngg��ny�����[��EG��;�I��iD� �^q&D��9�we��w#��d'nqɂx\�*sN]��y�s���w9�k8DȮ����&QNgs"�UΊܪ��TjAEӋ��8�Ȫ��Nr���'qg��]�H�IЋ�B�y�I�9I%NI0їHs�.�q ��W1��҇!��$���d.�Ws����&d��U�'e.�2�]��Yr�t�4�2��� �13�VzĊe9	�
.�)�.ULp�yAzyے\�VU4圻s��˕EӉƝV�E���f��AaM��T�X?;���֓	�]����V��C(�"A��.�ky��f닲��a�b����"a��:��5#c�uՍ�n��+�l�,(�&�lX�����e�*�5m��+qZ�TЌ���\=�і��n6�I�J5�	�f5�&&���u"��c
kZWd��b�K��XS�c��)ji�V��ɣ1�0�T�e4���%5�)��-��U%ِ[[l���L���0!����`�Wb��4 �f�Ḏ�Ye�Ֆ�@�Y�Јˠ+��k)���+�m����q�919�kq+/FR��x��<*�tkoח7��-Zֺ�2�jJ%s	�K.��԰��B�8Һ�
7M�ʰ�uCDm�D+��U�Q�a2-JPP��@�v8����Y����7ZM�h�H�b�3�{1������#v�˰�nķ�I�ӔKW.�@�V��jR�o��j�
�s�˄.f�Ģ)��Kl6[f��xTֲ����7:��v�0L॰�.�����L⭗S��M��]S�4f�8���7L�U�@������SXҮ*e�&e��\d�'�+v�36Q�:��wU�)Q���u�F�u�LWi�#�����tØ��f���2蚍�����3Dţ�%�e�������V��)�GV�H�b�%ɵ�.�ƽ���/��x��<�@ #)�$�{:J�i�-C-�&%j¸5�vk�� �����Sn
CD� �p���[�5+�D�f*�U��.��a��1��8�Eu������2+�k� ���5��*F��4�p��G=�Rk�-l6Ak��$t�����Q6�J[*�5r�өz����ZF�e�f�͖`EFܙ�Ј���!��T��
5a�P����vU�v�i��f�l�L�s�k6��A�h���v�Xh,���s � 57
i��� ���YZ�Лj�n�K�q��c�mH�fں���m�
1�w5��[�*�����Ʊ,�	`�L�r+r��7YX�]�`��W�Ӥ�M#�F�0*�s.5��!�v��)�=ep?���֞Kqؖ^��	+m�m,���$��K�f$f ����h��]Qv�쑄xv,ۥtv@2fLJ����P��
l*I�M*@EG��QR])��q![+ۘ`����vV�����-��#tf`7�1&��q(���k-�V��c��b���#��+s{9_��ߏ��6]�M4`h�S�+�aKn�myIL��J���6�֕���#���L�,g*�9�hW���U��띝����9wz]M���zyh����(�L�
I+�ȃ*]m�gzt��O��5ҽ{��T�!7��6�׈=�$k=E��*f����*�e�4i�*�18�W�؎E��;yA����{1yi�%�@��A�A�����#��r���d��c�s�0~����IB�wG�j�q̓yWb�(����>���k7ؙ�(�%@�d@0a#��S����h�j��/��S̄ߗ@ �s��0���~BI@��ھk��Â����6�3ʦ:�"�v�h�a�c,� �P���E=k�{e
D��0+^���r툼�ϒ�&\z�];��ǈY�����~��� ~H��n��`�Z��GzJ�����d�F���S`~U1�_ghQ�O��˥OЭ���ǖ���tn���zx�Q�p�J�z�0gn7NT�K#���=� g|+�����m`�7��&I���x�FA�P�"�{F��sG&8�+�:�
�@0a��F상�G��FU�[��o�[̔ߗz��:D�lz<F�Я���k��NZL�P�"a�@�'R0�H$i�+V���9v�^�g�o
��^1��4$ �I�!/] A`�@�d��20��uS��F:wB���ڃ��m�$�O�x�7���r�D㝾�5�ǝa���xX4X�"�Z�򴢵�\�l;k�.儢��
%�M�p2�}���� � �BH�#�n�ޙ=ކ�e&��H��zCun���I����(Q�2"�r
}��u`@�D��G�^&2s�lE�|�ϕ�<���"�/{�b�c�'�cZ�� ���`�_$�'��d�l�Ph������]@�]�P:Y�)�;̠�Y7��M�%��G\�t.�H�7��M�T�J׃UV���e�-T^��������WT���<<*t�N�7$�y>���F7��|dL�`�ݠ(tѠwZ6F���o6h��"�r��ry�0��~ހM�#<;OVdFL�G�<FvW�� ��(s2�Ô�Ӟ��
�Va����J���c�'�FH��#x�f�NtN��k�m&�t�J�:!eM��+W�K�C
u�αHub�hU4�Q`w�ؾ��_� ����P������?��%ɩĵ]�_I�}���A��w��"I_P ȃ!0A�{�;Έ��u�D�&�&�r{���y��g�sD3�0~��o�K��v�a������ �2J�|!�:du��P�k��ǋ�"v�>Kdqy�wf�F��U*k�p��>�D���?y/��P�tv?@}�y.d�o�x	Q)��Iwy�J�^(m�.�ua�
�Vz�Z�<��AN��Q3՛���U������W޼h�DT�oG����.z���P�Ld�t�����*&~������|��"IB�D�����tR�\��$Tl�)�J��}��f�bo�#��Έ9���H�����k�ߵ�3B�ۡ[hG[��"�R�(�k��,Eƫm��J�vl���W� OO>}b�I�5W����\�'m�䷫�1�Ղ�C� ��;��da��@�6h��h�8b:�q�^�;:�\�U]���V�ɽO�x0����PD�����xo��F��`W��?�&�2G_"��oe�T���+$Ǿ<ԩ���~���e��������Ѩ�bL���א��q�A��^�zA`SWx����"v�>Kdqy@"�ƭvr*����0�Ѕ�2GD#�3���N�����fB���;��%J�u:}��������
��;�E���VKc�PeK�ծ3$����״��k/j����\rgu�9#b��Sj�̢(S�31�
��io��ӻ�<���KA�l7J�����\$���V��d^���"�փ���T�b�$�6�c-d &iYJ؈�c[���,M,�(�Z��b*�ith�q^��e-�홥+.+)��c�b�)5,&��eh&��4b���eфFW�5��h#ZGHql�/eR��v��T�f.,,G%�A��7I�.iU��(��TU�Q*`��ιK�&����^���.S�04�����gKU�e�M�h�%lhMl�PR�SK��O6��ߞ��o���vA��Y��ޘ�ܜU37���^�ʗ�↏u��P�~���IB����
����^ll�B �G��k�����:OP � �!#��ǵ��Qm#��a���_{9�H�?C�PK��	�D�ߓ=��3h��Ӷ��M�}��H��D�!�IP�{��&U�"B	���?�H�5�'�/�L��bo�G�4r��m^��������
2&$B�#�%
D�"rM��vh0D���.�ТU��:O
�����FH��$AJ�o��=�o�g���eCLf���I�@�Ke5��E%3T��@G.��Ч�?���㥗��3�?!$�Aܞ�`�����I�O�{�E�^�f*ͱ4{\͌q�@�+�H��#d@({���݋��wc���e^#W5�R�3/r;�_C�
�U�^NER3GB�/�&����W��ӵ���,X:ȍ���/��R^>LURſ������G����V;��ܕ󉝝�M��@ �4�� �z*yc�Uv�ߴhw�8Љ�sF��*щ�eM��<�����r�]%[����b��#$t"F�$.3]�m�/�?[��?����(Pw'J������n�R�p ����ׄ]L����?I.�D��B2G�X��r�� �8���v:�3;����SS�g0�?D�"IB�R>�����5W���"�e�ȱ�0�3��0%f�֊%�a��f�`(�5h��E<k�������|�����`�b�ec������ H �FNP���/�����߫��m�M!�����T����<;{i]n�R�w�~B�P�"���2`��e6���� �a�0k�xa�Bz�3Ǒ�n�Uk�y|:�M�ݥ���`����Ћ:�����Ѹ�23m0��ɹ�YAV�R����xr�{+;.����m�>��#	��Ǆx�ݡ@�Ǐ,�����4� �)�(�	iJW��\�̬a��xW�@�F
O(��o�h���u��v���&H���a�����N�G~5�B�������ڭ���W��0�/#�0AC���]�՞$���$�`4�6�6�6��fZ�ܲ�Gj欪)K�"Q+�mZ���_~��g�`�!#��?H�9{��vuo�S+3��� ^�;�������?���}$b�2'� B������Ń�$��WV���k�9��2�/ I�#���=�˪�|����da�������Wǽ{��g�\��g7�ڭ���W�$aDy(Q�0@�$�@�/(T���X���d�D�}�+*]3����to��zXz�s&xd���@��_`�g���օ�J^��g�0�Q��O��=mU�j���׷[g��K�ir�g%���kb�\�v�?]��3(���hyʴS����Fg�G�n�@¼����gֽ˛���<{O�����ag<���x��?ke�D��
�X%��?����&�jśXR�.[l�[� Uq��ҋ�=���1����@/���=ٹ�������Z�"��/*0"p#@��B�Q ��$���0B���O�y>ƫ�$D͚��$�安���m�{�~�_F�B;�P�Y��Y��+���|F����|dLA�]]W����s�3x���x
��	��2GD�W�
�En*2��㎻��}�3���"IB�I�����{[5����<BY�o��3���� ��_P ȃ��?I�g2�|��a�\��[]W�������9��$lG���)��O�J��^�8WR�l3p���*ź7B��M�������3Q�n;C���b��e{8�f���>�OܳF�ވ�"'d���=�<��0�jO�/`� �(�.vp�u%�9�cs�#+�86��K�Kkps��k�ā
�f�M�[�D.Y]R[?�g�,`By��cD�44��K:W��l�^ak��l B2�,��l[Ii�k)Œ�"Am��5�TbB� 8�%E�εIn(�K�+�6ڠ��ڵn�Qq����W[�ָ��Ȭ� ��v�fT#Z��i�mqC
r������&�K���J��\��J�SMb90k�� R�Զ'H*"���_?�_�� �D/����Un��7{��1VH�c����xM�3y� ��$2G@�YC}μq����>��B�y�*o��I:����>�y����F�<�5o/ �dU�
� �#$tA�F��?HŪ���鮫�;��)vkk1����9��"O��|d����޻v����ݯ�X`S������e����=�����8*��VV�<�Q޺�a��$u�/��ت��}%1o�]�(;�{:�?g���7���@#
��/%}"ρL�Ŋ����6��K�Ki6R$a�f�b���k��D���\j�T�ŚO�e�؃ ���:g;�jŶ�����m�zJ]��(�N� ��\g*�s�ѧ��bq�����W���4���ʆ6�U
8Wc�FN�.�TT�<*����[��RmV,Ô�ߧFm1��xF��`���!KEW������	��-����\����|�z��	 �D wvjk�8U�T��
������D#�_%'��A���%�m-tj�:��f�R�q�7�B��O�>#O�v�eAb�i��Nx��6��>ݑ';�Tb�j��mf6�� ��9�7�M�'[�UU�||�<C�B�v&A��~BIB��J���7w���H�n�6vO.p�oq=��y�	̈H�#x^<ń@���T�))���dm��\$�iX�3-�#l�76��0�8q�V|��Nt#y�!�H�~�~�N���)V�uM�]6���z0�j'ֻ4j<�\DN5��y�.&��~gwot�ۚ �>��f�5�U;Y��.�|o�׈ c�>>ޛ}���זwP�s�h���r�ǜ����+S3���׽���cV/��rV�ڑc��Z�ʞUԶtn�)Z���S�vKx���;�of�]���V!/��(����n�t�x�`��gU��U��[�ߊ��F���%K3�ݘf�d^j5��m����R�{Vy�%s�Z�K;��f�̸*Ҫ�'"{.�L���<kC���ǡ���!�i�sW�c�&��B�ћ�
�#(�S���w󡸹S�	�P���M�2��6�`9{kk9W*M�YBnno-���r�V�:Oh�.�gn�KF��Z��}S����o*Ŷz��;8c��^��jXnM�КYQ��b�.�7sm�PKFB[ՔWs5
JY��/k��[�B����y��<Ŧn�MJf��f,t�UͷX��w^m[,�=U���dڡ�
�S*ܦh<xf�C�7�Wy3/F6�v�S�]L��镶$�.N����!�����Rג�`�]a"k������jИ�Ln�vs-Y�����!��~����������~Kb�J��&�:�dt��)�D�5Z�JJ���P��^k�L�6�m;nf;�1��X�w5�P<l�ѷ���si]U�Rij��ad�������a���Mp�P�Pڭ���\��I�v\;^���Y�o/9vK������WJ�J����v�,g=e޳m�Us�"�"���:���Q�+P�Z̥TThHS��\6��Lü+,����fD��GtA���w�������s&6��쥙�+���lg^6�M��bP\�{���kl�IRV#����ҷo4ֻ�-��Թf�1X7�Qn��y �7�u�;1�۔_�@$�
_%A��EǞv+� .��@I���M� ��*�4��L"�)�;�EU
���U�$	PGuaAQ��TN�ke�ʀ�֑E�vQUNdE:uJ.Tv��.U�.I9E��$�SbBB��s8Ŝ<X�\�ei��vS*��u����9E��Q@�2�!��G"�r<��A\��"4��
� -Zd�N�Gr��(��e9��MW!ʓ�;I�=P�,�@P9���(.DU]��$���""r����.P+���*�����Ur�����E��/+"��Q�ZI%y��t�܇;�h\�,���<�U��b���tS�$$w/��3�8qY�����AD�: �#�.M���-�'C�e��>p#��whW���CS]9ٖ�u:����Q�4�V����u2?I/�L!|d����jH󔰹���-��uˮ�v�~Dq�sD�|4�wdO4{��;�Z�tQ���D�2f}TA	���b\�fu��h�an��`���(�
'��#0B[>݌ �F���KDw��^n3�z��U�WP� � ����A����: �9�j��W���6�Kݾ���{s-^�꓎4��dX;��t�s���"8��}���;�>�#��L܋�ي���J�Vgw}�@�~��D0���%
�Ș#گ�ք��t3�Ut(�> ��Z��_I9sy�Ϟ�P>6�O����3���ZB6(˭Áް�.y�˫��i^*��\H�u�zu�+x_u6�#�����:\y�F��(N��.]���{�h�����3����^��%n/Vl��ltγ�.�jN�8�	`�y(Q�0 �zy��Ge�5��A4+�J84���K�7*f唹�U��h�ݮ9��-̻V�PP,�ǵ �?I�@��ݵ7�cꊜ��ߟ@�e���C�^��u/��P�dL�D+�%�k�縍��� #�խ�rK�Nf�>j�� ہ#�Dݒ�<�ѹ�\{�	���#���(2��~ܳ��Ӿ�>�X�RuI�H� �m
�݉ �4ǈ�ڡJ��ʋQ~�9��a>MO�v|�+Yq���*n�~}��9�(^d�9����~�/�ٴ( B�G����]vTb2!�Z���%p�:���|��|m��|ȃ��^#v��/�wt�������Z�3�t�L����kE��{ ��#w%s��M{/�]�ڀ|E:� �C�o�w�����jҧT�P�?���J�A���-HZQ� �P���4Ұ6�/\` �J�KHu�]����v̻G�.r�ds�b�Uգ#u�h��vf�1�w4]��e1�d�(֡m�Z����1�э��@�d�ݣ %�F�����
�"��l[q��\=M�]�tۛMAJ���0�J��s�*b��*��X�Maw#5�A�2�˦����4�g�=�����M��(�K���|�x��r]�BSc��u:�Q�H(º�޿З����{>�'��ݡBV���gNb�I�N^��v�p�/e
bH�$�@�"�Vfl��[�e�L���s��"A}�d,�ƪnw~|o�� ������t0�T���mP��Ո�:Ќ�9��W�bq��͛��<�z�r	%�k2�ǚ�	�|A�d#$T�3�_!_^���|=�Y��  �O�>�ݡ^��jQc:wjN�\p �F�!m�q_}�F&�ϡ�A#�$��a�����w����C�D�]|�%V1�1s���� o�����IB{s*���,�ٔO��T�&��5î��.i���5(عԉ�v�B���n�������H7X������K��e�5}�A\�;+����յ���T}�"s�X�%G����{U~�j�q���U~�$�NX��T��[o�U�1t4[N�ᆳ �Yf�yB#*���OE�ҝ����j�U�n�L���-�������T#>�q�|��mMު��A"7��"��7�s��2'��f���.<g9�؉�X�؋��1Sy/)J*.w~dw��s@�ц~�����2&E����T�z��	�C�~�Ϙ`�&A#
�7�d���d_mpTA�"v׮�K�(�tGj�@�$tA��~�Vl�}�k�����B�3��cc�l�N�\{�`�/6�"`�D6�{3�p��>���$���Tf��r]��Vʬ�v��j�[��DEZMR��T2�}�A�A�2GD#��n�,W,u(�X���w�!��b:��u�l�e��G���I�pO�䅊$�;�g��z|C=���jo2�毻m�X���� d���U��nVA1��̎�?H����$��T�ó�c;�����y�`��Q$К-hRF�)=�S�!������Wn�y������x�\-�Ҧ��/�祂,p<2�Mʾ�ٷh�Ųv3�Ƥ�/�!�^JdL~"D��X�y�)�����D�׈;�'���N�:*.6��@>7�}Ց+sb�;Av(T�6��` �
D���k�5��/��S���o��Yw����@7d�/���F{/q*o1h{�Z��!b�{�b�bk	ZE%fRg���1X3b��8qM
z��-��묲}�ǯ{�/��)禜��0����9���~��"�e'�t�a��ޫN3�囏9A�C[%W~�C�a�F�+΁��s�ڹ�[~} �|�����ј�00����Ⱥ�f�Ԝ�9�$4��Я؟HҞ���,�U�t;x�=�̸t��c��A���d��F� ����s�Fr�3��a��/��J2�������U�+\w� �1�-P=�]�t��c-VR�g�Ȍy9"�L�X^��A���q^�/�W�*�u=�+h�^>�)J��u��wv��$����W��y~�x�G�ۻt;� ��Fߟ�r��'y��BGñ�]��5&�6���7�}A��i�ݡTn���g��y���Y��U$}T��m�R�MG��00`Z�ˣ��S]v�r���,�c���}��4Õeh���\���aձ0�9oQ)`>�h`?B����a��/� �s/5wӾ�LMu?r����[;Ȉ��Uc��xo6�ج�]���:a�뺯r� �a#��BB9`��W����J�������]GG��I+�"�95ְD��w�� �ey(���J��u�l.YWY��j�p7�$c�A��6�U�� da��H$tA����N�S\
[��ܪ�<����HW�k9T����nJ��~"��#�U����ت�Irz�E����(պ�b�F���fR�p��"&5����b�On�po[��7��X^���-�����}��6$�0�E��+�Kvvz0���[k�f��4#.���jR��]4bUZMc�˅k��9�c�eZ��5!�톘f��\[4ʀ�юc�h͘�fk�	eI�����й��cm��TJ�m�
����iuk��`�.l!1T�Bۅ3J%�`Dh^�&"�&�=�fF��m%B�cvf���86i]xɶ���[[GMLF�-��f�=��)e�f�L[�<l6(�ֶ�VR��m�v��봌�I�M�T��g~��>�0�d��۲'������LԛX���@48u���׿{��s�9e��Tg9�r�#�"�9�w������O��qZ�\��nJ�wu��K�m@�A,�wd^���&v���U Og:�3�A|D���޹�9'�+�N��^���&��]��D(@�(P2&�$�_P���]=��?d#�GD#m�;	=Ꙛ����	��.��3Ly�ߏڗ�ͯ�X$B�2J�Ȼ(��Xt�VL�`\���{+�]ԋH�{�z�`�$t21HI�Y�F�g��U�T�J�a����x����a�b"`E4б�fx,��YTa]m�~���Y}}c��>��앨�|�L�r�U�)8�����+���"tb��0A��P"IT	�')$�Y�V�I�e/{6�ea�6����z��H.�)�Ƚ�a����s=P�7���w��v�&�;ӋPw���� <<䏏�l��D��Zrkꊚ����7�4 =� C�2��u��}lq�0AqD��(ȟ�D7Y�{�����
�9�qﶮ�E�s�P � �'�FH�"��J>�4�5�u}o�?�܂�ɴ+RXs�ʩ��V�����썳Usz굞��gA�j�by��759�-�BH�G���}����C��
�g��ԩ�����| ߵ�9��/��*����K,�_�@�6���Hܼ���]��{k�9pDh�R�W$�seH�����'��~{���݉�KRs}����݄C����~��܆8B>�u�F�$2G@�'nVڦ��\��^��'nٿzmR��l���/!@���B�������릹���j'��MN��%�ٯwd�uCzq�� ��n�kuø���b#�oDeP����W��F�n�dC\qٲ��üg
�++7f�Ʈ�ɻ�70}�x :l;*k�S������@��tA�a��K�#�H#"v��\O�P �����Ҕ��{��&��a�p�,�>!�Ȋ�8�s��Bs�J@�$tA����b�Ě�s��7�(vvÞ��<�f��]��!@���@ȟ�z�vP��6�_G��h�ҩW[�l[y͌K�(F��(�Q�cb��k�#u�kbj2��>/��q�՚��_ݚ �ȟ_p�*�ѕ41[Oȉ��oO����P�Q�9�Q�*����TD9n��8��e,��_v�ME�H�����	�2G���m�|�������@���%�IAK陊v;��CFΌź�ָ{���.^ �
��y(Q�0AB�"dc�쑱}��y}v���"\�ջ"@��l(OY쨡��~\#׽4�Y-M�WJ���jnf���QwD�V8��@��ܝ�u(Nr�>�6n�YZ�k^��bխ�.��q2��5���Ēѯ�ȃ��� + �~�}��� dL���s���o�����Ք������{�l����i�q ��2GD���{�=�n�.����XT�*je�`�"�s1��V��V �4��[7P�B�x�B%5�
��ڏ��+�C;o��އx�\[q���0�]f��h�3n��$���%�� 
֔1F��R���9�۲+��
5�=�1[O˄�M@�>�|"����B�tH �� A�IB�2'�J�~�T��\;��zk�麩��}@�����#��20���oY��J�G������/��hP{��ms�\��<��p ���=u|��Ew{B�}��	QG�a"��ۚܭ��ɰK�a�Ȑ��z�eEV���ޟV9}���7�Nࠏ�s�r��ys+�Q�M��Z�d�wVG��9V�^m��n@����^յ����번<��ɮ%t����m��7o*���$��i��)Sw7�Ô�߮gt�����µr��1!�U��ͣkJ��f��Vڔ�;up�3���cՊ[�@��(N�I�� ����u�rnD�#���9��m�Wm<�٥�4&�Peή����]xQ��aIk�k�	V48����r��Qbɧ�.�l�jJ=:��{�`��ƽb��^�nk�O>趚���J�\@�ʶ΅*p�����d�ɣ26D2���h���4"5�P���ad���B����ȝ�s���4]+��YRAw[�1#��t+*Л��1M9��^�Y]l-���]��y���$��B����ޅ��R�g��#�X�dX��)�Ci!D	��7>�f����Sy���V��z��#��/-����)m�b�+CR��/^�2iK	��˝#Q��0R9�v����8C���/s;V�Ud�9��:���)&�v��"���nm	�g��u�UVi��woj'DV�;�ĮWx^�1��pi�tC����4oya[{8r�э���u	=�Ϸ�.�0Q�K.�<��a�}�C�%�'d�wW�:��Z�����^�5F\T���j$,�u�0��%]0����)9b��ö�o[ܰgׯi'���Z0_.b����2�����)��J�-䒠���ʱ�����ܑV���!���^��u*B�qנ��^EpJ��W��/���g!�gT-I��5�'��+���>���!'�:��ē��@疞:�re9�ܮ���@�S��H��L�qՎ���n��8RBBw��\�*�<��ށv뻙y/\��mȎ�NNOU�	��\HU� ��Z��!�e�S^����N�i�l�2�E���"����Ȫs�\��99�\y�u�p��&$����g&��Ԛ�N�!��{V/&1 ���91�tiNL��
(*!*H.�9C�u���͝��2z!DAC��n��:@SKS�{�y�UE2�Qs�ęCϞwVw���1ԇ�P��P����̒N�L��NY�S����-���9>��Pى�K�����W8�#(�.���3�Trݕ��ieSg�Q��6�-��mi�W6�a�qiЛ6���]�����D���n�M˩� D(Tt[-�Zk�]L�"M�9fk6����AV�A�+#5�Yb��Q����W38�ݮF��j����f�bY�l�U��Ķ钺h����L������7�+Cuk.(;CX��a�wJ�)���2Ҕ5��u[��c���&�6Ŕ4t*����� �����	�n��)�鸒�&Ym����C8�&��E���q��m���U�u�:R��.���[�d	�XRZ�t�KP0[��M�k�%�+jb�¼C�ˈ�K]�%Tҫ[Wj�du���]�heBR7K�j,�u��S�r���Ҭ�[&�H\Bƴ��\YU��)H��5�P���e�$I�l�K,{Z��V0Ktm��$�HY�B����HR=��1�2�t�д`4��!�,m��[5�/��{�
$d�X��,6�Թ�.ܪJm��RX��f�Pa9a<<@��,���s^������tHM)����,��1Y�%h$���I�-�f[��k/К�Ҷ՚��mn���7Q	(Fl��p�uPĲ�3���	��dĭ�4�S�VgMж[�2�TH]@
��T�h\�F.	f���M/nj�kX���1ѷJ��������,ښ%ёI�\�n��������1�p�� �E�nC	���t�z�vuDҵ,��h��֑2K��!,�MG%K�]Yn�ɝ.���`��`#.Z.��^����B^U���ݒQ���]����+*��j����bËm�1�Q!�U�:�f��oej���ViL��au���c1��V2��Zif�,��Z����!�1���͹�$ū���\RE���Κm6ӱR�%�*s)ve�)v;:2��J�*�l.���mk4�Zͥܲ	*=�j*��]�:`q)�s]�X*&y�12��5,S0�2��f.uTI�i��Ґ�k��e��wt�<夹+.Q�O��:�!b2l^�eqfk
n5Cn�Zb���#�k��Sk-M�����&YZ��.���E+.�]&��K`���^-�طR��qu4#p�mLǊ&��Ƒ8-�Ij+uLU�m��D���C]f-I�C���]H�H��:�����78�"G;P��[,R1q���Y������*�*n+�4&R-�T�lo�������%Ɇ���M6`�í��f!n�����uhM��iM�=k� qDfРdL�D(u輇�����n�zG=b�y�
�J�a�Я� ��w9�	`���#���.*�F��϶#ǻ�P��s���P�k�n<0����B�2/���Fx�PՈG��@��|a�H��Sp���Ju1�a�G���+i�V9�F8��wd_��H!��y`�<�Q�������5�hWRV��|wdD��{�o�dh.���;�?�Є��H�q��n�rȸٯR�B��8�[�\���NWܼ$B� ����}�4/ש}~�.N�����[������uuC4����Ay��vn���}{��!�嘄=���D�"@�A=g�E�I�t3u�]�=�|A����K�$�_4�j����w��/4�� ���'Nu���,�m��$2t9o*�0N��2�9��㹒R�̶���"�y6~)�es����>~ʸ�O�����?}ګ9u�H�*}��ő ��٨y�sz��V&;�I��[���}��(����ri�t�k�n;�B+��_H����$�AWT#�)���+9A� �t�vD���r	�<�(b����M"Ň��X�s���m�"�AB� �%}"�7W3���τ���i�ݪ��7[��r��� �Ϸvl�$tò�Ѿ����O���+Tb���G���'���]h۩�bK��R8�u�-6bʢF��"��A�a�~���H��Z�oԤ�P�,��q�UY�98x��<-�/٣C��.'Ns�������&�,Wgod�G)P-�p��ʢ�+I�t{s�ՎD���1s��T��0zu}$r!%M*\�B����*�%#����$#N��YA'6p��8(;#*qI����U�-Qξ�D;PQ���;CQh���'����{sV�G�C���9"��Uf�7[����W����ݒ����[����؇��d�zej��t����p� �	�J9�\�nW�@�$`H��� {Y��!���}t�����F�b����z|1�݁��>�qKU����Q��Ld+)R˴S�Xۖc3��dDva3m���UL2�N�TERuy�C7�E���	�y*�d�n�r��b��Wb�ʴnE�H!"�Hf̖\Vd���3m{�g¹C��\7�%���f��U5���B3Ư���)�G �k�M�Q\�hw��N�{MP�{�=��r�	#�g��y���}����
hV�����ݵ�|>�A6���]c-��q+x�yl�I�,c��{�/6
~�O<R�n⚘I�̪n��'�b���w����#��U��m`u0s.�B�(�K�]��{�{�Y��$BH��}$Y�x��^�O����h_+<+�t�k����dn�ݷ�\��������~i�7�]4V��[�wX����l@����J� e�ԫՆ��=�&����N���Shr5C6�{���3/:ڧިbrG"�	<��Ś��6�E�dc�u�'��Um��j�ǆt��e���s��m|�}��}$���iS�X:q�i�,�Ibp�y(wgv>I&U�f1�o�6�����jv����%����E�Z�Gy����bD7`{wdn��1kf�mT�×n�_"r�^���m�$�	7����3�e�%��si
׆˰�d=���m��U�$f�KpfR�2��.�)�x���m�f�H9u���ϵk�2��`�ɮg��Ӻ���i�b+�����%l	X��V�jXᮀA����"@�d��[n��É[�X�E��i5���.�����U,�5�%f����
Q�J@��B�惈��Z�܄˵� kn�ň���166�Y�[Jkz�ڵԄ�f`e��e�%55ņWL����\��ֈ�s\M*�Кda�X�W�����s���[�X�
��7�ߟ>���k[�a�L4i�`��b�残���HiM*Ta��֔�w߿>t� n���������8k��e�A]�ˋ���_	�?������KO��#�U�{�Shpڡ�I=��1�&�5����6��L@tBH��	7ڮ<�D#�N8n�9V��]lb~ۀ1)#�D$"��)W�x�Uݡ�$�׃�u��7Ibp���s{}���۱�"D$�nW��~�jU�@;�m�������ϱǷ`n�Ϯz��~����st��-��E*ie!�Wlm\ c�E�.�3J@�L���H�,�_�ö9*����z���T�����)����ie0R�v�F���Fix_)c���	��Q�V�N�>Y�	Ǧ��ڰr�SAIT��N�`Ë��9'm�"��Z�˱/�q���U���ϫ������|�^��_p�ZX�<���1!�t�s@��¦�����K�Jq��;f�c����cn�N�����ᜤ_I_ޗF�@YU����o�IQy`]������MW+�wڢ�k�J��I/�"�H�Sc;{r�-���r��i��ZX�<����ݰ읛��i>~={K	�gc��C�Ŏ���5�����Ap#���T�$�R.�N��i���<���I����mt2u��5+�7�OEy�ylI$��c��u�˭]�+��	����{o����ܴ�p�n��1�Wp��@�A��۾���E���N^̣Ц��ι�i�W�"*���ז�3v�<̢*�mY�O\��a�
�^�m�gf0�^j�o�+s�5x(uS�� x޶4�=ZX�<��J=y��wwo����q�ݵ`n�mqW-������ޞ�ULy�ӝ;����r!�	#���љp��	v�u㓛yk]ph�$bO��iK|�%�3Xd�2*2��hF
���q�|�f�U�[t�h6��JaI�YB��M�Ѡw�_ct����܃?���s�X�<�j $cMs��<�Nv�{wg۱7�"��&z7�,0����׼�姼J�:��� c��v�g{Z2}����v1" I�є����è0l�O�yt�=ל�������@g)#�J"����apݡ#����ۻ=�7��=a�Z����X�M�+�5Y��y�ڽ�3�6e��a,輗���Z��2�X�k���qn��5}X���&�#&8i_��Q�j:�\���7��"�k��W�c� |����@o����"�I=��8�}sR;����Sf14��l��6)#���;|X�ax"C�m"�q�B�.�7�˛6���^d���]�|�$���?�R!�e�]��g#r��uxq~��w�������s�E��#��.�O#2<��%���쎰��Z�����;6X���*��yK����IH;�u<�ɎÓ�w+�x6cO{�kg�����k�nq�IO�[~ݬ����yK���ֺ�+6+v�+\_K�<�`��c"�}$H������n�_US��L��;��k/8�37v�hQ�,��]�]n�����omù�����}�n�����p:�<V����`���#S��2���Д��C�����4�|���>I'~���o��KΌq�3n���%�u�s5���H���������7�ό.+Z�F�۔	Wsi*=���=i�Z�h��I���	��5M@����q\؉+7��,����d׶�S.�u�Qk�����
�JJcp۲�(M�5�0�7�v�Z�+)�m�MHѻtMQ���W�c(�a���4��.�9��c�XW�����G�3�in蕮�T֥���7X1�)[��0�eb�5a��q��w�G{�{���s��m�t�1�Y��<��;i�Mvu��BI%�"�{�{�`����T%��+.�}<��������p1����huUϷ�����ݡ����neuW��5y��{3vq��6/�#/��	6EXJ�t%n��3�v'V�W��vl�&��kdB�����c���v7`n�%/�s��噔��s��v$�����m}����!�������5V�_*)̛]��^����PɭR;:l��=�D����K�n�@��`�X�y}"�H�Od��{pwe���ڦ�d�j����1��!$H�.U��չO�u�k�����'fk��UX�n�֊T�Ƴ�x֗��A{{�3w,����;�=����(%��U:q�L��'��S�>�N����o~f�Ji�y�ϱ��뫾c���E��y}9L�H����6����\�l�^�v$�����m 3��HĒW�Quz�Lz�F��k�i��֋yz�-w�������Wݨ{d�� $_	'���s��=6:m��Z����G%4���l�������;(��&�T-ۢYM�B�pW$�UsR�G8u�en�%[Mh�,u���A���_�D*���w���q'&^���}mM��^̶�۱����#&���B��df�֙�}h���2����7P�rn,��)���*[��I/�%�_��uJ�Z�{R��vo$lW���!�$g5�V|��7�W39:���兦�׃��}�10$�}���O1�:�|��1A|j�mV��н,SQ�wnb�Bu+��b��iࠫ�����3	Љ�k���,�D�O&)ԑ�O6�����o����2�d5!���]�֞`]��!��[�(55�L�;:���-��1�]�ڑ��Q-ŕ%�v�QǊȪ�9P=s�M܅fCuQě[3��v��L#>���Rݒ��x��3�����1c�w^�đgUM�F6n-����k�suUE-X�{�p�S�Emk+�qU�H�Eh�X:X�U7�����%R�$o^�C�|���ݥ��uXV�;[V�-�A��#N�`�k�r=)7(Юo�gL2�>��T���h��Eg�d��(�"���cD�X��Ia�rv���:t}����[#'v�5Mԅ�hu�m&�7u���T[՝jŉY�#gO;y���˩H$�[݁�{j���ź�]�|kQj��nm�ON�2�kYv�WB�w5��R��hNĦ�͜�#ˬj�TO���]��Q�⾳8ôa�E �Qͫ�Z*�浒�p�E�A���X�=F��+��ۤ��cWf}5���5C{Z1���4�Wm��hu]�:��������\Vt͸��'A$�p&�nꗘ�օ�(Ѭ�
�/m���bfX��y�E�{/N<'�*}��~�[:�,#af�qYɡ�ɩ�S%]p��{ �<��'x��S^�H���ެuYjB��OZ�_e]B�:�ۭP�,��h�P��_?��|��>:%Afyܨu�*::�5��N�y���Q�y: H
�٭�'Kܙ�zs��/�e��
)�����7��s%S��S׮�c��f�s�*������4>NyTp�!q�f�R�L�9<�-=vr���v�)D���N�$خ�Q%:b=e����q�ܹ��{�Z|��:d<���gIusݪ;{��J��G�O��1�<ޔ�TR�˝wsw�`��\h�����,�\Z^��(<�gN�ny�lyNWɤ�
^��ޅ�X�C���=�9�(�RbJ(N|��H]V�#�J��"~��;�J�w.'f�%4��ٲl������"�v}�ݽ��U�c{��ۉ92�N��X����2go)�H��	�k�Z�(]�{\�7A~��Y�7x�{�	#�E�|����g�x&���)�5�v]���G���hi]E�F�UI���e�i�6�#��5}�I`H�a�׫�|b��]���c�9m�d��$�H�B�h���ʹ�}��ȅXv:{��}���/T�|6���I�}ɍԡl._ofK�JIF>>b���G�~����1bL��{7gv�n�����x�]5N��Cޏ�%����|e�]>m��b�n�����iJ뽧�38��&7�T�X���2�Qa��uZ��c���gk����ǴzW�w����zn��Nq淭A�9�߼�/����/�_	#"�̂(��c(���O�ۅ92�>���@I�M̮vÓ�x��o�Map6�W�|�|)lJ����m�[5��S��a��߅�1�_IT���~�q��&[�F\O]�ա�ᘖ܋�#E�v��(�t�{�w�s���c��ֱ�\vꮥ��v)����ߧjǟ����1"Iг>�i�o�㽱�n�����m����	�f�w��I	+�nZ��F�=���(�X�-�[ R˅'	w^p�q�0�I$��E��2�J�I�˷�n��[mp�R(����Ү��n/��7��y�M6hl���%�o!�Uvv������z��4�x]���y�u���8� ���3إ�(�cq�����e_�_����f�+�W	cZ�it�X7kf���T���㉈������nMh潶��a�2��\�v�WF[���Ŗ�	�QN#�ً���e���l��LY	�J�P�$of�Ԙ%`Q:�U�i����f������[kc�\Ej��׫t@��j8�2�V�.�B�0ՙ���ƫi��i��$�����Mq�������4������X/WK5�4bf\�[ml/�1H"�,SF�Ru���_o��%U��������-���jW�8�\_)݉���N�^�5|V��M��]w��e��[ f���>˒��q�>��3�H��	5��a8o�����/o�J�o��|�_�6JG�qo��{�l��>ޏ{v=Wf���/��S���_hwJ�B�M��j�}$`I'z�#)/���x�c��Ҍŉ2� � ��ݍ��6�\���U@�����ѢB@Me9B6������s�Pi��,SF�U�Y^�bt��*ܳ���\kj�e&�����|�y8HĊD"��k4]v�>���0]�_-|�l�(��]�5J[i5���Ri�0�Qk{��T3+����Us)�b��w*�h�[�U��8D��ݑ? <:���諳P�}%�Xjwr�k�+�g!$�4h��7өn����!"O{�n.9Kg��=��b�3w�w��	#!�	#ϸ+U;��:k�EN`��r��[Ws:�]��'�
/-Ǜ{�=����n�JI���ՖhU��wQ�v᧳+T���rF>�����H)�|���|�����Ț��[0�pmlh�U&�n̤&`ɨ%T@�`��&h��W�����I�{⸼���bL��W΄���X� ��y}"�1"���0\�A�-f[��;�S������&Խ�f��Qpk�W������}$bD����E���
جb�o�[ٙ�9$n�bv���m<�X��Wsv���Ym0д�nw��=>�����nǦ���s-jh����4�t��ԭ�Q���q�q��I%/X���Q]�b�9|$�77|x{��ť�2�{v{f�*��*�Qy���$�}"H�����A��lV���y�]-q����M���������Q�<����}�u"�)GXM
�����vp�knÌ#M��D4æҦ�TU:%"�����H�Q��c)V�(��,#�U�@����}$u5V>yxO?�����swǇ��"��������$rB$����d_H���=��h"�}����^��5�w�I���>�ݯn���SX����v�z���62�nR�}����.�fW��
�E`wʬvi���%���^"�xj�rj�^�s3:Zg��+D�N�Xol�d']�:3f�;dNH�2��Mm��/��y���BH�)'����3ޠ��ܸ{ْ+���=� 2G�I��Cbf�2ZD<,w�t�"a;%5�vI����\�2�i2W���SH�S���D$�	�ػ�s�/n�Uov�{���>`����_O)# $O1-�r9��W7���͌Y[��_{nr�H�`$��nU}V����\�}$�OTڡ/�k4�}�r�ԙk��f��_	�RNlwtA�w���$73����B��ʤ��u��wEv��cw��¯}9|��H��I����헗�_�<x�Oj���*c�}�-�2G$5t���N�E?,�Y~w��������]U���fSb�h��sM�Plо�;t�f�r��O>��0Bh檎�uS��Ϳ����wԔmZ�Thn�w�Q!��R]�3t�;a� L�!��:殔��@�,�0TL骎jKm��`�Y��C/d.D��P�t׬��L].(`�Tk�I�%�Y�#��U��b��=i4b���l�t��!�K7.�2˲���MM�ɗ����/����B���#��aX���7��ѵ���Z%v���[Lփt���4���-s1����m��V�	la���4�����&k�j�ږQ�B�f1����� ���E"G�rx��~�/�n��*�+N]�a|��z��{wgv=]"3��q�/zG(�V��.�r.�]&�½�"v���yoՍ�� ;�I�޼{�]@��p���ݕ��*5�ہ�$�$�ߞ�Vs�)���y|$��4v�S��Z�|7`"\��15I�H|��BH��$��wf���
�{ޗo9˵����_l�7v�u>��Pޥ��,��K2� �;ݒ�(����)H�ͥmq�kx��R�MSd�t�z}�Zw���
�kc�p�n��̕�2$Os<����~�BD$����xN��'���N�zv������R�}�8p�.b̓��Aa֊�n��4vU�kvb��z����b�'u��xt�����f��1W�e�l�ǻ�/��J3/��9<}�����KJ�{uӘ7��z��|�~��2�2�����Ȅ�I�{�|����]��d' n����˄svV�F#�����ycg����^�`{�H��1"�����c(�t�fքة��K��nǆ�ę��+P�7\du:�	:	4�u,�%�آE�`��&ACqf�	��s����]=~_k�����[���y�nZ̵m�����1mGf5�=����Up�c�`�.�QQvVOpq��J�1|6�q��d]u�{V��dP��I+�!�0V׽5�s��)�X�u�ټ�\/pl�{{/�*22�'}3��rs�������*��l�ݛJJo*��b N]��'�)bYѦ6�se�����9��)�Ŭ����$��RG�{�l�go2Wz�w��/���v"�)v�ܵ�j�\�Ϭ�N�hemx�z�)	�`H���$�E	ffؽ;p���G����db:��q�q$	[����v��g�}f����&���Ku�nܡ5(ҳ\�����&���j;Cj7	j�/�`֤.ݡ���x��*/�)�Ŭ��E����J�ʶ�ls��I/�#z/��`�w�q��K�|���V��_l��	��u����=�&���_�I7�s���g�;�ѫ)C���#��m��8F�E�j��}~��[�'�P�H��.b�������}����ѩ:.�1S�T���Ꮄ4wEB�K�}W����o�E&@�3F+�$��Wz��=QM5t3��U�l�2�=a���S��f��.�$��y	�G"E���]꺺�/����Os�����3/o�x}~�"�����n_�ʟ�6[e�h�E�B�Vj��6�Û,
�Pc�Q1�*�]��]D���}z�v�h����tZ����x�vM>ϮguȤ_I��-3�����f��P��"��:[��y| �Iu=����{m
�{��_I�{�u�Ӌ���e�y\����V����$���M˟g�=�:�	��"��OQ�y���G_�o�_8��M�!�%	#�E%�r�0����{i����壬����Iǻ�b�I� $߁U���Ky%xrf؂��u�5g�㇖Q8���6�0K�r�p�N�=f��i<�YT(Pݚ,�ڬ�:��Ls�%[������}Ww��g�K=+�mR-X��o�Α[�ho���:���qUb���ț�웯.��X�Y�j<m��S�Z�����O#���u+e���ΡP�.����v����9�޵k:��5�e���9���I��a_���q5��;�w*�ek��>ǻ��,))�YuAܭ9a�(��P���5Sn���ڄue��o���[���Ԁ�P�Vr�9f![Y;d}�.Y�&�f��`\����j�}7�P�uuYx�X���y����^u&����EwZ�+q񎹴w�T�#�qS��c�v��!�e�nV�k/Svr�`*m����R��I�>h+9�w�r�N�r��՛X��-co��YK��9: �e�x*�C�ef��h��ȷ��u�aW#S����L� Mk��f�]�6�\��/2ђD���������b��ؤ��2t[���ŧ���D�8��*�Q�m
Mb0����ro���4q�3���Jvju�S���]�
D`/y�m���!)��۽��V�ڬ{3f�|Tv]"v�P�w5v(��*olaS����)���Շ!ۖST��`��ɡb�����㮂P��m���ԯRq�j;��j��+*�
�t�	��tt�.�T�J܇K*Q�iT�����N���w�8(�p�����W�۞�{�p�3��ȟ�x����|���%��7d�Ju��4,5ᰌMi�q�N��N4�9bh.���bCk����E��t���@�2nO�$-N��	�o:b��6&�1$k�v�\H^r'5�,�C��Giz�C���{��\��(�g�	��V�RI] �U�	�x���#E,.�� �f��5�bc�l��'e����.��91<�*.^^��=r#1
��AE��fe�B�%C���	=[��D���Ɏ���8P0�&' HIzMvMn9&:�����ޖ�0@��IIP�+��] �o>�d�NN��N��+�*�*�[�U.��r��,��@-Ň$ �A�.�T^��^7)��+�-q���r�Tmu
�3��13�At����f	�X@�f �Ժˈ`e3i6�oc([	F�M,�a�67f��c
�*�j��bY	���8�5v�AU�F���K��ԭ�l�Ha���[h�XU�ci�M�����ݜ^i�`ZÛT��]��2�����-J5O�r����ČI���LM(�]�;Tڅ�p��"�Ʊ��u��Øb"�	45#,B-�K���;��c�e��hXJᅒ؄b]3�tM�sm�m���н�vmY�jU�R�p8�7mZ���;�HZ��9�����l��Y��L���-���"͛�mɱ�7!��4i�TiQ�Qĩf����X�`�.�F��Y�j�*Z�B[
����Q��*B=�9�5�$mM�.�3��)3\�9
�ra�+k�J0α�9u�\U�X��̈́u���.x�j�f	�U��I�!�"a`b�:�l��qR���SA���Z������jb�96�3\��w�j4��:�cKV�-Z�.Vީu�cw:ʨ�TMGun���^6L�7��e��� l�+J��Y���q�U�����J��h��,\�K���;H���S\��D��fv�+���P+����#���A&I���Gu#qX6[�i�'3j�ss���ѭ��Ŷ)�l؎e�ư��S-�ⵂ�ա,�L��M+rf�Y����ae�IbU+��5��y�[xr93��+�:b3F�)j�c�R՚�XD�\�Bh1R�6���m�au�n���ry�a5s�����eu-LP32Q
�X׭N��s���{b55.�"�2�<R+��Fi�P����2�%�����;<1m���FqE�kM���qT�U�˳@ג�.����X� CEQ�f����a2�6ˮ���aui�%5SJlb0���ˈ�ڥ��K��٬%t�Bʏ͕��5���+�&R&6���f���KYXຳk�&J�B�:��)z�ve�������/T5�Tr�:g�Wk4z���)e�jNf�b�֥�l�#Sn ��@mݥ%�ЙX+.*�k-�kTCj�09˛����L3V��	�[^� �+V�{s�L;�`��x�bB�R6�
͂[a��W�����tf�D�X,�Q��M��WxL�e�6�j+]nk�-����a۸�W$#��.H��l��h<�6���k��  �$��c�χ֖��*����F]�k �4��\6hfe�tn�Ę71��5�$�{\=�ݑ�j�춲y�o)[zj��7�M��.�@Ώ7wwo�w��oV:��'qgwU�ފ��Σ<�9a�9�������x�9���}�%�щ�	#�Ԡ��zt���w��l��w��$r/�RL���-� ������-U��M�rEf�R������zbp�>�]#�E"�I%L���QΔ�L��}ϸ��f�說��$��JX8^�u������1�nHL�e��{i�	��鈡4�1ܤN��iI US0�l�L����I_	&��*4W���n�-��7$�72}�J�1"���U뻡����0��y���ٻy�.`a��`q����2�,к�sSx��ۨl9s��·{n�|u��y��j��[�kTuv��' ���㞚7%����?�)3��(�����I	c~��ߟc���4k��s�=F�L�	jj�1"��y��ű}$c��Z+����rN=��^}���G[��5r ;d��H��p�9�U&ko�G;PY�����/��")%z�oⲳ|���O��P�ͻK��YT��bk�R@��R����rM^�]�I�M����bE"���p�y��}ƴVi��| |E��0K'`��ٯ�$�$�'畉w���q}����N���b�{��|�7v}��oFKs��U�|�s�$RF$���^��eO
��uյ�w5��\�nPU�}���H��m��v;�.�e��AP�{��K��*���٩���D�u����|��{=Z=�4V�Ƿ�=��с�H�F$(T�꩚㜒M>��S��=��Wiޜ|]�e
�uw��t�f=�ңpu��Ϊ�:/�_I�E&�:�JvtS��|=ػo$������U��0|vK�_����-��"��-̹Qe�2��n,j-j7-f�ʘ�mZ	�H��,���'/���"W���<�B���m��p�:*�3zH-\TydRG��7ȫ}#1��m�U�ἣ��B�]��v9����@��t;u�"!$����+'�ٸ�Ǌ�҃xgm����	$�$�f>�R��1��E٬	���Ź颒��m�z�ϵt�B�{ih��9�L���w0�����������Ab��5+�mw��ɴ3!�S:D���t왣S�Q�\n�W�����	#��ַ�t6#�r�o#���̡X��}-	�KI�T�{�U�y�Q՚7����X�]����e���;`J������(�S����	�I�f�ڥ���x�p�s�&���>��+�۰7vG�^^t'?b��+���|�_�qΞ�E+R���-��f����n��ggM`�LO/��H�/����fo7�{N{çsZ+4���jjH��H���J0�� xSH�7�n�Ә�*�|1�����ۉZ��Z{Y_V���$r!�ISժ�d��3�N<��)Z�M�]�dR/�����Xŕo��&�ǋi�o�6�n�2�:�Z=C���r?��X���9ײ��+��7+��u�A]��kUn�ʐ�^�eК��%���Ɠj���VQX�Z@�kR��Fe�L���	��e�*���lܰvu�X.Ձ�lI���6�Eiڙtsi�a6�$e�0.��R,��u��07X�60��:QCW����K�΃-��&�C9��K�&�"$���U��b�sM.)�ݥE(ke��b���V:��h-W\��r�Q7(���m�vz�)�̦����lnu>z��m��P�!u�6��h�-Qt�IZ�
ۡ��c1�t��UN�H�^^�s\�IV��-=�ӹ�+4����(�X#�}z�f�bD��."��\.�_m!61�3T{�׼o�����}���9<��Jס�^�$�G��I,} �cH��{b����uf��z�{��td_H��0$�u�Y�-S�U���W-�Ac��s�k��W @�eT^�僕<�{��I�	�؂����q��v���noh����I$���)wU�շ�R+>@�F�UTI��5��Z$9,hf�8�����r�����kfC���'� =�ݟn��o-�nj�Ro{�bDc:��Y#1{1:wwlnǫ��R������l�vE�h^����۸7������h���P�T�)�i9Q��E�jL�{�p�y�2�<��J�Ƴ;gVGDP�)����N[��,�Ŷ�I�ӫk���W�/x>��\k�=�3P��H�RG�'n������w�J�S���ƻnoh��ۈ	#/�BH�k����͎��]�<7`U�����{U��������ފ5Ȁ�IbN��⌣1�ne>=j\ۭ�W�W�6I'kT�F��hXN�T␃a��7�H]��7a�iZ���k�lt(C9�b+L�?�W���/��nVH�ϭ��.�7�wxs�RҼ�Z=���]��5"G����;A�lUd���	�/K����]�6��V�OWG��sT���7z1gmAX��	$���*�{�-~tP��n��GE=�ܬ���wQ�p�	i+�.������(3�Q�7v^Ҭ�h��6-��j|�n�Q
�0���=����o��BjI.L2��wSsa~�t}n�n��['��WT��M�ydL���y�s��q���1"d��c��3rd7 I�9�}xe+٤��w����A�eP���!p)�4�$�D:��Z6�ˋ�i����G�Ը��f]������߾��$A߯��4Owm�j�[�<�B����m�|O_��21"/���+˺�a��rm���״�ܛ�^�2G����s���R�(	�y��w�>!(%�W�JF�B�+���.�z��Ӽ2���oG�ݎh����J'���!)��N�K�[Y�j��n� Z� �)Y���OO���l���)
���DR��k�;�v-����]���j�iW`j����������b`+:�k�DT�����BO/KI���l��	����2�����R� ����	@��t��Y���r�P�j�����	}���r�Sh|@���$kR(�������G�g�o��D`�g*b �K�Ys�[e,�E`��̬�[ClRʶՂ$ĺ���]�����ӿQi��SQ�l�������Ϋ;I��<D��
//3ѽ�>��>] $��	(�
)Hw7r�˽���������ߠ��͓W�/�P%��@��D�`�;	}��ߦ>����{A����6���KnV5��z.g��X�ϯ��oGû��A{ H�y�:n�Cn��7Q٦�����MnD��Я�
�]-g�뾫2���r����M�P��}��\6�W��Ă+�4Cn�y�AmЯ���Bc�Pa�P+~��낹��7{�K����C�>�$6�ۑ��H�����&�,�Q˥��C�7t��l�ă�Q�om�ʠ{y�i\�X���w�'>��*\�>�ȵ�+�X�|c��%�M��Dt6J�F���ɮ��1�.���­c&��M����|�؋v�svIZ9�ۮ�%E��P`��LK6�b�[�u&�m[	`ʽ�kWF�YV�ii���]�T����w���Z%cm��:l)�����M�=��ۙ3( �K�@���6�S���]�Gk�
���(b�Wh�8Z]�r�b�)�YXj��:�&-�������	4�\?����L��$n�١c2J�ⲍ-4&q��.2��,I�#��R������>�΅x��ۚ�7yq��>Ϣ�䷣���
�>7�n�����~{��+����^ �"|Cn�m����0j������P�������)\m'��|}���5:��D+�泪~�)�I����@���$6�Qm�|܌ߞT�6����/�����6�d���K��y���� ����t(�@#��np��-w����P+�@-��ۻ���U��/\Sz>��q@�/���8{�����)`�ﾑ$6�P%�4A��	N�u���ԨN�4{��ٝVv������4F�>n3���_o.]�mK�_��% �R��F��%����լ��3%ؘJ��aU6�
Exk���܃v����|܉;ߍ'�Aߓâ�~
\�{�t�__tP�"H����܊ �����#�Һf8�}tE�w�,V^g�|�\��N���F*�7�*��e�K\y�D��c��
�|k��h]��_:y�6]Qm�ں��������}�������o\Sz>��(!|�͹���s4ݎ� �8uȒ+2��@/�� �"A�����O��1Y��}�fR��O����{�ju��<|ۚ!�#)�c�fz	YP0�k�Q|�n���~2��~O���)
��h����mV}��x�yU��E�O�>-���
�������ѱ�8|gM�>\��=�q-����q@��6�A7#n���޷�>{����
�6]s;XH�Y����uձscf2`��r�ء�z�߬!���E�$۪�nEzm޲����2���oG�dP���Okܩ�E��^/�H%�4Cn|�1�#��?Y�}��wҁ�L����O>���â�~
\�����wH�yy7�B�y�H��zJ�4AmТ�O� ۘ��sw���9�_UO9�Kݮ�X7q�Bs�V���ж��Q�掑#!nH�n����Q�u\�a���������i\Q���v�Z�ɑ���C]�5']OAmW\��5L'��Ӹ����X�U]�_rIK��Z�T��u��tY�j��>߲v��Y�����Gz�ԝٗ�ͤ8Ԙ���-��v����}�-w2�D�ݒ���j�0�H���� ��7!�C�QķvͪȜ#t��1�c�آ�0��B�KQ�]WD�}�ǋ�(h�{��	b�S9�B��:o�nM��3�r�괾�2*R��]�ed޾ĕ֬���컷-�Sב�B<�]�\X(�@�Y��(*�o�I�ͬ�.��nSqY�E��
F�.T[ˊI��z�t�b��]�Q�j��o�t�5V��Ih�7��f[�V6�:��yK�����Z{d7XY*�]�I�v����k!k	K�|*�7���,t��Dn��흘��v����6-2ʪ�!"6�бg�Q<m-lA�����v�+���s�c���-�W�r���5g6F+�5P�ݶ�*f���!g�scr&�JT%�Z�bÕY�h�'n0ma����7ϳ,�4su�^�4a��Z0"���QN�P2c`h[��J�ڧC�W{A��8κ�v�n엮q/{��a�ܡ��m�w]�Q�Z�
'U�Rٿ=�ˊ�p�j�v�)��lV�\.���mZ��K�ϝ��Nn�*��e��pa;V��*�vwU���k��[:M�(q
�R��
b{��u���eϛ�ƕ9���A�'(�r��p:aoY^�z�<8�;^��U*E�q9NZ�AG9A^d�y٥p�"�dW9hbϫu�O�ȯ�v�$�bDQz!ȹQQQ:�w����" �Қ\��9E9����H��*e\��U�I�p��$�\��ޱ!����,����,;"���}�2"��z8Nd%��
]®G����9q�H.�㤔y'*��z��AW��*����ܱ
�L��r��:�US�	<������>i$�aP�I��^qLEa�S�Y\z'ޱ�= ��]�_7�EեItҎ��'�b`%O{�*�J�����$8�V�[�N�S����*�P(�6�.�J'��ޝ7�G� AG$��ES�ڝ|��v��w}@��'��^Mϵ�Cn�7J��Hp���34 [�$s��6�T������Ϋ����A�s@b�7�[Sg��sb|A=��@��P%�Cn�ے9�
��}8���"c>]���U���Uo�O}@�o�t�!�U�ۡ�?��=x~���=M��u!-�L���fJ�<-y�̫+�=��0�k�l2bh,�O���Ye����e���
-Ǥ��oyq�����r�������O]]� H��w�|� ۟$��wo@�L�����#�u^=�R��f>��(Ϋ���ޏ�A7�h�NE�u��A��S]��/��@�p$[t(��AȌw�0 C��l��;��ZyZ*����|^}4wH�۟Pmכ� �N��<�)��T(��[sC���7��|3uܶ�ß|(�j����.���~��O5������ v�$���`qs���I�i�';���T�S��ڜ'oP;n�����[��|
寮]HmȠ[sD�I��%t1w��;"o:�	t��;J�)>ޏ|o�� �N�x��A�'�>���_@$���*�M��j͚�c*fKx.������HPИ[�����s�	ﺅx��!�9�h���Fm}���>��r�pto��F�y�O�6D�>W�ŷB�q �[sDS;k[14��zAi��iq����7]�h|9�+`H ��
-���.Ϻn����@�s�Yy����|ۡ�Gݍw�CR���/�Ls퓴�r���|}|�S�@�|ۚ����O~m�>�T(�s@[�>�-��_fh�τ'�^}>���{�+�#1Ϸ�in'�͹��
��d�D-CO5:��_��wm�ß}@��$|�
-��7#�V��~��C��ם2�Q9�k�,�&��fQ����s9M���5r������ߧcy���\1��]}�.�5�s/t2�
����t$Ѱ����� �݅�i��e�T!X-���lni�b[�%��F�іޡAdL9�haY��fЙ1 찵���
[�b�t"2��%��[rU(�yŶ�ܑ�%��5.s3Biv��5��(�fYu�.����7R;]��u�TRj��--�M5b���ذFX�u�Y�B�R��M(�3���)�vl0����5�c�NMr���oY��H(�3+@̈́�Ks,"A�Lh�D�¼���#�D�u^mȯ;֚3���Gi��'��}�?���^I9=����(�G����#An����8I6�L�c�=�5�� Nr�~O7���3EU�!?��>��m����p����}c�ܧ��{����t(��	mɲ��ޕ�l�;e����>��P$G�Р[s^ ��O�mרG[��~��5�Ѵz9^ϰ}�$���t(x�Fz{�ci��'��MO�r��s ���ho�tH ��Mt[� ���
-����߭|�����o��}�������y��#��Cn�����������F�/꾜�j*K���:k��s �+H0��fl��ɊؘR�hM�u�>����W��Т�I�nh}�5���:��C���P���e�>��ܡE/�� �"HmЯ6�����ݿ[�c��su��U�F��]��k3p���$ʳHm������,��:��5���ybS����-��LT��rٱh�d���+�}�(e�ډ�z>ciT�'��}�7�h�NEx���Cx~���� f��_�@����ۡ@�� ��
�}�^�q=;Sʩ��ޱk>��uO���h��"A��ۡ@�C�:�tf��}yݯ'<A����������z�����m�w}^�|�*.{�;Tf�nv�]4AN@m�y�4!�m�%Q��ԓ����.���fz\|�ҩ�O���x�9���P-Ǥ����;>������ѣ!H]�Cp�9+h͹.�SE�q�5�\WH-�����_��~���,�'���O���r&{V��w�-}{�.�����6:��Y�o}:A�|���ۯ7 ��ы�D�mt���m�U���75���x[����i�w}^�|G�ȯܛ�}������~\1@�+�P ���Ȓt+����;9�蹋����NtJ�aJ�,e}��ҩ���3��?y����^��i�6}q5Գ��fJ�'2���Wk1�ٸ�p����ٝ���S�����>�s@�5:�q�͹�ۡA��k��w�}o��7�~s��L�-+駳�gڵ
��J�@���},��}�T��͸�`��W��B�q��4mȢ�B��_}�7ѹ9y�k?u��uմ���H�� �>n�ۚ�2�����p�$���%���Z�f4��p�"���M-�*�mdCDUMb�����P'�����^!�B��mL��|�Ҋ�O����V���GN��_gϾ�R� r��D�Am�ۡ@��I.��Z��χ�/����3صG�OzJϵ����
o�t�!�x�ջ̣w6��P��8�ڣ�u9�mТ�H �ۗ{��7��U�Ѕ�H4uմ���H���'��͹�Cp$۪N�}�q�)��/�� �Ux��C'[{S����5��oG�7�5�>�����lZ܋S��g-i�7���٭�h�c�nl��K�}��;g��[Y 6f��ķv7�K�Q�]��j�+%�a�f؁��"���f�dL++��̉ɹ�t(�	ۯ6��w�!��f܀���}[��_N��3k�+��A��׈#�D�;����wP��m]��2�b�Re"�����|��@��t	GU[3@���3(E�e��1S+�*���F���������g9�U�o�][Hp}�ɽ,d�3���kr$۪���ً\�=��B�Zt(mkl����1Jk+_����'��ԓ�E����]�?VQ�6������?��$6�P-��Aȟ�7�W	���P��ޅ�Z���N�������'�����#An<uh�#�2Qn:S�s����b��7�.��>��	�|Fqi8���B7�4A�D�u^m�G��$6�VQ���`8E}���T>t�5�\}�R������}�^!'"�q$n[뿬�?;�]]��}�,)�Tg^�U���5dkqJj[ţ^#�͉G��=��N���v��4��m��El��#p��i��p�h�'mAK*��b��3ZDt�1i[c�e:�x����U��*�]���yO����iR15������+�s)2�a3��m3Qrld�͢-,�[l!!�6�gTa�HDC��3���$�n��(@eKTl6{S�q�a��%�Jљ���&��R�܍-�\a4MS�W0s�[m�l�vqC&v��C��k~�Ѱ(�˰��R��VYu�^�"\L6k4z�)���u3�fW�^�Ht�-��7"G���_S�ޅ�w��n|'{��q��BɆWr�8G�H���x��B�n$�[sDwn|���>��d<����0�@9�;3��Z�o�^�Hp}�@�� ���6�}���E'd��@�R��$6��ۡw��W�կ�����U�\�E�)Uek�z>}�@��
�� ��!�^�r���.b��;Sn����t(��h|܉��Ծ̽�_k��f��w��@6��ľ��ص�|3�e�B���E��A�mϛr4��B�<���\�WLE��׶���A�|A�B�m��+��L�Q�'�P��g�ˣJ��E�ņ�[��b���6\FZ���%ҿb���9�4 wH���
ݶٯ�还�U�������<���Y�[��u'=�
}B��$�[s��כ�)�
m��$Uѥ�ʯշ��I��r�Y;*��;zfy����AY|�7o.�on�>=N�M�1��,�$M�s��Ŝ}}Z-T���%>��{���2��}�ֱ��'{�@�M}�"|CoZ�u�~���EtzA��>�[�>m��7ս"}�Վb��m�>����A��[sD܀���`'��[�#��u^-���5���J������ �� �׽��/�Y����؟A�9�u@��HۡE�%V��9����.D�s����/~��W��n�'zG���hGt�۟g�t�|m�y�٢bb':��\��3E�殍�k�,avk�r�0��e���3D��A���������	m�}���ſ��5���}C�/�w���t(F)_MR�� ���,����ꮄ������
�k�W�^6k�=C�/_�����	9[�8pځ3"�_iͬ���4Gb��8-�[s@�<܏���>�����R+tDmI҂��y@��ޓ3�$�V�������'f�EeY��;f��9�[�-�bn�a�xv�wCG��r�^fl���⚾W��j�X�߄�}^����t���^!�B�q>#�K���fvϨ_*{�Aۚ�{y9���߆����>�(8F|� �di����{+��$6�W�s@�܉!�Q���7���g(Ww-�:؎�!�5�����M�Mx�t(�A-�������`o\W��|,�t-V�@pQ���ɓc3`�TԮ�lQuvL��#H�7��� ȝ�(�tGr;��^\����89?��C^�9��ط�]��!������n��a��Q��8���X+"A��׼�M��w�-�>�#� ��t(����1�K��� ��x��An@m�ۡ���˹���;{'��o�wd0����M�M�^n m����x��9���qe
?}�D�3�������F�۬N��W|(^}4x�������V2��w�\���e�X��J���^J�K��K젔�P���*�3G-|������&�%:��aP@�T�ɑ��Wh�w�H��|A-��6�W�q��/�A��;��y�֝�Oq߅����ww�?7B�mϫ�ȱ�c�Nx'��$���E!TuUj1Јd�x��[����#k�m�#[˝u�g�{�
jh��Cn}M���/������x�2��^�L�ϝ
+�A���-��>ٮ��bXD���7��x��	��������߷X�τ��
�M{�H!��6Bʚ��z�n������6�P-Ă	m��gW���\��7��Q�k3C���W���G7"�n}A���PM���n��<C�BN}^	�3[�S�5�a�e��z=��3�����~_\�g���ſ��Cn�y�AmכsHY1�#dA���bjdH��o}yz~w��'3�+������@m��<=�8�G(�)��~$�m-�H����%��]C��H��׶"T,�r��Z��Y&
��tt"�)sZ,�c;+������Jǲs�;��;2�(���tG^���y��+rd�[�9�_m���!Hm�Ŧ����}D5��Zw[�u[�`#5�rW֭8�t���ve�u[S,b�C�9�c0Ԩ����l�8Wf⥖��J���̷�����;*<���v��9L()iEd8�)];.���Ǭ�d6��l�Q�d��rj��#*�:4Ⱥ��!�)_5�:ee]�zy�����֞�k��:5b�Hgբn���_'��~I���fNɕ�:���yW&^��(�������$Kr]���`�r�[��r�}�P.�1{��͵�45�S�{Qe��pc�M
Ա��T&j��k*=�#w#��ꮾ̹�<҆�静v�3���U҈���k��o�ɤf�a���E��y�8�6i�}rꮨ����4U�[B����,�%m��R���{�%,�B�(�ќ�5FVf7�i��I�Ś�RLQ��2��O���U[K�ӆ�k/Z�V>�w(De+5��F��4r�lt6wE��*n����QhR�3kn�,;y�2V��XV=�Fg7S�R�^:§���;Ck7-�^���9�*j��islҽʺp�����kv�U�+�,?bչ�Qt7v���s����kU��]U_@E�bT�ٗR�;�F�T�K
uIX�Z��n�^���˰~��b���M��F��U�m��"u-J9��4a�0�4�.
6K�ƱαY.Uu�Z�=�RHr�܏�$�d��V�sRQ:T�bYL`��@JD�;�n����uʈ��Gw7 �q̃R�ZU�� �T�J�'CA9G�I78\���s����d%�Ru"ȪI�+���ӔD�DQ�'$"n�����Q蜈�E\�E�(��j䲹wP�����!Q�)̤��Tj*�#6^���Q�CL��I��r��eȣ�UQE�*����ȋ0�-B砎�9�)�Mj$��Veܩ2Z�΂t�*�EEEE2�NHȊ���X�Bg%\���I�++��r���ȋ�YQ�i˓"�$	�r2ŕ�{�QTd��"�W.G8Ey,�ԺȪ��

�UUr�p�UneW�/Zh�� �LrB/Z�D�Y�2*�(���U\�K2��(�;9	.l��JV�U��Y�R�����iE*J'#��";.PJ�5ZIA�Yz�9�TW+�(!��s����VATjC�88>zޮ����:=l�UCk�nin���;7�(cd��ԇl�t�F\Qwd��A,��kæ��B�1[��ci�-�+o9��fl,I�iNlT�98(��Lf��z��0n�`����x��+[�Iht�w`M]1��Z]o�Sl���L�E�ye.�JS8)j���
�n��Yt��`���0Yl.��F�Y��0�׮�(� Ѥ+a���B]՚3,�s2V0� ��ASA��ll�n�E�RP���,�RY�t���3�\&cȄ�(���a�ƮY�9�2SR�5tMe�:���O�������`��&�ZjX݁����L˓MR�˞U+M2�CZB[C.�)qe�	L5��p�A&��&�,�kl�խ�	#�l�n]���,-�"�G@cx#t�̐�aL�UIcE���0�V���M�E�,��n�Wp\D�b��f�5\f�X&�ʜ�4![44)�0�n.љ�� ���
�I�X#٭V�dlѵ�����JS,&[�n��JU΃���١F��Gm"l�Z٩ѭ���*ʜK`�l��.��5�3pb�����Թ�DG5\�Ֆ�����1-��"]U��+�4�[�g��X���7.����l9M��Xn�������i\��΄qطs�B�l�&\��"%Z�Ee�텈��L6��P�vI�F�Y���c5
Ҙ$�,4�c�C
��M
b�S�cnm?��/���ML�e�;<�cV����CE �Ӊ��d��\h�ư2���.�5�˘\�e`��d�eni��h�h5v�u)ƥ���R�e�ZV%�-eŷ���H�t�0Qn�rX�B,a�.%��Qh�F�,J����5.�mK5l+U!j7���:]bh�a%�qli�̀�nj (9,�&�1d�i�2�/o ��k��y�9�,���g]��WF�]Vl�t3�iج�n���hk��Z�:;�l��&l.4P�6�^e�^ո�)uBa�U4�s����u�[�S2�Υ̭s��:
���t)�-j-��4�.=G����@�]	��0��ˠ��p�
�43�j��[��JV-C;5r��a�QB1`�YFk��io8��K�l)��:a��iA�B͌XYR��9mSkE �,�l��ج
�����$-�m������ZZ�J�E�5�[2��B��!��X�FiW
��+k*kJ(P�o.��ϥ>��e�-,��S� �m.�1��<�q�XfP���6������|s�����I�滖t'5�o��bh|?��n�'�;c�Kn 亅�܉!�"�[s^9��)_�`�A�/�^�/�E��~�����5������ݝ4>Iכ��!qb�Q:(�v��	��B�nh��Z����Bc�/M��%����[�u���*�MGt�!�U�܊-đ���y�g�Îz��_*S�O�nk�ĩc���9�����8�"q��y�*/_�zt|�@m�n}A�Cl������ޙ�گ�w?]w�����]x�{:}I:q ��ۛ�������~���w���䴧6��v.h� 2��cPm5�[1+��[�ұ��s����`~|�B����ۚ ���n*�/O��}���pU�P̟߮������t�� ��Ux��
�n$��4skg�՚���tU���n��'&S�f���%^J�v��Oiі��m̦*p�����N��I��cf�ڋp�\�V��p���>>k��u�&������z>���p$B�B�nH�����'=�$��ǹ� AnD���z�@mЮ�;迾��K��m�]��LUe�����{:k��y��ۚ ��
d\_P���U�A�c�^-����u����?#���/s૾6�� �ͧ��u������,��}B�n$��5�r(��h�(��4ĩ��|K�������z>��	�H+�
-��p+d��%����$t��jc�:,��%fp�DCB2� �����,��B�g��m�sD�D�t+�6�W�+*���Wi��>'5�L��5��DΑ�)��H �ۚ6��	�	��f���/���o��4|�M�v꿶�����n��O}@�O��6�y���&���s���r|�4��9�nF��Iŷ$BO��Zp��~�}���\����:;�F��Y.-QAK���Y���j�E�V�g/�=�[��>R�Av��o�U����F� j�	���5�fk��|��K�A\�P-��r$ۡC.�\�**c������D�����n�$���W��6*����|�:h}���MC�����A?/��Cn��!�B�nbٽ����;3w�r'����mo)�n>
{�@�M A�����۠��w�u��phI���Q���MZسJ�](�t!��5�t��f�mL7k.����}�9�x}μ�g� ���v�.�����z>��|�}7W�(w����@���nD�u^m�>�#�]V�"����	J��u�6*���q� ���@Ru��~0�oѭ�s@���(�	��B�-���]�ʲ��}����Z�Q��cU������} 6�W��t+Ÿ��G��`�VM�Wm
+�H>-���_ �~����z>��/`I�s�ؿ���+([�(l]�&�⮈�Ն9L*��(���>�b�(A����t*h�Iɨ����ػ��g��c�<o�u'�F"�=����S@�;�I�	mϛ��6��UĞ;���Nu#�]g_�ت�k�q�gM��@��s+��s�<զ��i?)Ɓ��Es���{L���Tfٺ�n*;Wk�K�4�%���a�i|���-��|܋޻���_/���)*��&!)|Ԣ�dI��PmЯ�H%�4���ۢ�er'�ZsC��k��e���|�}��B�"�nL��LQ�G�'�e�T����7"Hm�x��8��>�V�S��.��-�Sv�ˣ�}��@�5:[� �ۚ6��$i�b3r���@�7\��N�|܉��ͯ�������	_�W}@�^}4D��1�i�e1�n�z�C�7�ۚ�
��6tm?��r�3��k�o��5�e��|.���w/�@�p'�΅x��7!.���"r����ș�6�Do�]Q�ȓ�ʹ��J�V+�аa����ԛ�B�b��t���F���WT��.��vXrh�s*.�T#�kٺ��+�Z�#
���Yp��\�f�3L���h�!R��m5ä�6ة��d�ݯ)ژt�rl��%۶��DVBJ12�"�M5� J�Ж\�]��(b0�`��쬧�Rˎ%��X��1H6��R��z؛X�6ּ��$�+"$ɍ������uL��Ic��4ʄ�m����s���,b�p$�ʂ�lc�6�c��-��nC����)e�0�Q��J�����x�&�[�J� �,�H��V����'��d|u���!�B�ې�!���;?6*n����7�و�\�*~ �{>���׈m�y�C�ͽ����*f��yO�����߱�,����	_�u�����{�D�b.��<~�������x�7��
��>-��"ֱWݧ����eN]�����;���q���O�s�n@m�6��B�b�W)�AjD��Яt(9Z;��gY��Sv����ǻg���&FF��w����Mu��I�B�[s1���}���5�'������}'sm�����Ϧ��D�۠+�6�jϳ ��xa�`����K :�f
�'�yc�%{Wj唫�.�]M�̒�Bꕻ��!!����B=��ḓ���u!�]WV�|2���w/�\���}�R(Nh� ��^m� C��-��C��J�}�*h5���aJ�����e�t�f>�<�n��.1S!mN�p�gZ�YU��`�
��ϫ��w�)��q����B���ˣ�=�>�jt+Ÿ��nL�0A wj}mh�AN�r(��Cp8|G^�usVoVgo-Ϡ�尕�_�/>� �H�u^mȢ�I�*���D�¾nl%B��=>-��wR�����㗎�ùH��	 ���L��^��Q]�7�\d-����΂�9Cn�n|�6��Ī�?K=�����|��\>hTݽ�t �O���B�q ��/�}W|�%c��5�U��v���b�B`���6��u�#`ư�k�J��R�T�N���_g ;��ۚ܉[��5�nu�'*턯����-��;,��ٽ>�����x��y���nh����;1�YӖ���ĐA���H.���s�^;��@�����ۙN��	�;�X���0P �5�r$u���+v_O:�Y��iF�a@J�&���&����Rd+/��28�wE����긷U�n��g~�p��0U��Щ�{����v�59�q�>i�۪�>��6�����@�A�B�_}4-ȝ߯i�Տ��.��J�
��@��M�igK�c��#�U�����E��	m�x��ۡE�k�p~��C�9��>}_L�m��X�|/����:�n}���9����z�~��~�h^q��kal��h-4u�EK�I�ƙ4�"ЃkG��%ҿ��g�~{��/~d�t+ŷB��?>�=9����ߗG�Vz��t�}o�P)ğ6�ͽ�p'�[�}�!�+߾��M�ޭ�S�s�a+૾	y�� �H�Cn}?{��/E��+��|A�;� ��B�[�۝��ߊȭ������kX�|/�q��|�Р[sD7HmСKo��	�9�).}6A� �]U�ۡ^�9���4.n���>�x�t�9��ro����q���hM����UN\�P(�k1�	h[2�-���.#)3F��gPu2w��Ǚy��8\��n�@CuN(��χ���|A_O�z(�O�!�B�[s1��ӛk&��ȗ�oꩾ���*��*�
��(��A�t�!�U����y�?֯�y_�g�<d�T)Ske�6
���*�4u@�E6����,��:�c�G||�C�ϛ�ۚ��=E��}�U��������%�tr9��E��nD�۪ŷ5�(n�芆�LT��1�_u
����V:��q����B���ˣ�	��A�y�1��6y��Q��/�����m� ��
 ���r}o���i}�SW��Wr�U�W�>��@{�H!�^�6�W�q����6=�B�� �ۚW ����Ͼ*���>_
�>�ʏ�tE�Mhϡ�����l���D�u����܀���c��1����������=9����ߓ��Οjs��	m�{���0�g���Q����5�.��qz��Sٜ���7V��d)b�T��6(��y��E�%٧-K��d:{f�S�;9<�f�q��&6�6��}K^����6JeS,�+Kآ$i�[��4��0e�H[hӍ�t���X�Q��WL�tC3i����+��3l�K.�ы6Ma��DWE7k�Z[k�p���Uu�#�!*�[S7:Y���#I�6qn��]��h���Ha��Űre!0L��VR��P�h���e3ֵq�.!s�eif�[AV�׿W���>jX	�i�Ʈ�vì��0��r閣�56�FU-���_��z�a!���=�B�nh[�#9n8���g�&�[*�
�B�ϖ�i9�|H�s�܍-���[sDG׳9==TQ���D�	���\�������[��|��N8A\�͹�j����郹u���Y
�7"@!�U�t+j�1�/�����>7<ê�G�Uv��Ǿ�����Qn=%�4m����������!}���|AnF|��U<���f�.�+��>��O~(���Tn/��0E������`�n}M�qVk���������gf�3_I�ퟷ�U�����P'	 �μ۝!�<J���=c�������"��\��,����e��kT��m�e�� ���M��A����͎�#��b�)*a]b�j�&��ά�cW]_"s��O�V�s2�	��hc�E����?�V�Y$��pԏ�?LUF�m���,ʮ*�����)d��Ṹ��78����U�]^W�[jS�W��T�d��0�g��5��^����D�|�w��o�f�.�}��o�t���w�Y��J�K��Vg�(������A�n��H ���>̬��y]F���uֵU�������H>�
-��7"|Cn�P��-��}֏U�`R� �]>�ۡ^��=��Vw�Cٻo�q��t���}3����>7�$�s��� �H-��nR����CqI?%���&������OG�;�.|6��P ��h�;�H!�U�t7:i�=	�]���E����QN�d$�!	��[�IT��3��\QA�lm��R���,�\�뿞�?	����
-Đ|[sS�P��}�n|�q��wo�)7�B����rp5B�R�AnD�۠([s�τ�?��eU�\�>�U���}==܎ֿ���V�k��'���rt(��\�ϰ�e}}U��#ǚ� ��H��	6�͹�A�c �w��V��:������:Z6Z}�L�󊭼{Q�+a6�â�����^��U�N���5��
�W�F�Uq�����VU�4���m+6�o:�_rc�-��w;]J+�m�@�uF� 6�����7X�6������gU�|M�ٯ�g0��R�wfd������ή�	��O�wjQ���)��p�geX�Y�R�z�pU��
���o)ǣRS&�U-��ԉ-R�vA���.�(<��:ė�՝)�j�µ���O�J���g7�[-sʧ��̝ #�wX�M˼�5��_1Ûu{ �4�w�)A)�-�lY���.�F7e��˕g,PR�2�[�e7Q"����������z�K�$O˭�ݺe�i=��:
�=����Uݱ;���ݛ1�!(�e7wO��vf�*ShV^<���Uwӎ�Ƀ2q��2�V�q��ف���d�0�����f֪�����Y��#ݓ��5���ӫ=��Ӻ���ʥN�(q�V	�NmK��gW|{3N:��tg3���d�q�wp跬�ۭ��N]T�-=j34]���:��qn��;�3��$� ��y2e��z�R�ub]��%�4�/Q5e\��6���tj��tùcӧN��v�t����R��SkiL ��T��)z��M�U�AZ��H����C6�U�vީmJ��n�wJyn2�X���^�a���:�htXY�.]�PgF��D$ң�Z����7��Jq�:��}��:Z�1���=+.P.l�ن�NS������vR��n�;�a����N�i{)�]��t�17�}ӊޡ҆�{]+n�����};�E	U��Uf���gH�(�QUDswIΔ���Ŧ"9�#�����"��U�;��.fDH�DQkH��ETTW#�W

�"����aE�#�A.S �"�*8Q��Dg"̣%ո{����kEi�*"��TG9]#K��Q\���Y�,�I�*��V��n���!����UI�{��*��RBr"9R�TY49L".�4*�!	!	$�,L�EI.l������W�J�2(��ʳ);C�$'T��:\�\�hP����Q�i2&r(��u(���]t�dQ��Qz-�e\nBG�*U�C��)в�WI"�"�S��@�s��\ʉ��C�(�v�E2�i�r��wdp���*�C�6�	��q�i9�L<��	��9YYv�!"�.\�L�'t�:�v���UCTJd�SU[+�y���9Ǵ��r���o������$����>n�\�}�G�7�
���q�ۚ~k��}W��ϕM���W�����O{�M�?0���^ ��H!�T-��n@m��}�#_z!�
ut7�v����	�sDr��q�[o�����o5���h�PYT�@����.��ȍ�`i� �[�d12V�-5���b�-4\�쯼(�@�ﺼ۝ �܉���N����r���o��F�U}��C���"������mЯ�A��Ƥ��Cu�s�{��ק�UtO�Y�,�E[��}�P'	�.t(۟�]���ϝ|��>0�ߕP'�s@�� ��z�|ۡ��lF���w�/"����͇
������{� �:�q��[sD6�v�A���<Qam���Ȣ�O��|�Bfom�&���}����"-��8���7Ļ��R=&+If��%;�7-[��_K�ړ�G��\,����m$��{�h�4j"9�RU���!�Z]Y������(�H%�4AmР[���.Z�OW�&�)wW�1_g�/��c��>�|q��\�P�>�7"}�TԺ���~���vH6-5�b�fT�i�̱t�,��A��^�1m����Vo�o���?>}����!�U�t(}���.����p���z=�ޕ����UD�C{_WL� ��
��[s^!�T-��B��mL���+:(^�G7f�?t����O��[Q��¯��H���hGt���ð������kב���A�[� ���%���}3�c�;&�;�XWn���}@�����΅x����y�����9t�]�8N��}A�B�z�=7���q�����c�[[�ۗ��Y����\w�>;�Mx��
�I6�P-�ϬF�����~y!)H|�w�~̊M�*�{��]?�|Cn}A�A�8�=d�)�QY�����3���c��g_�t��V�4��.�9���ؑH`�9]F.NMZR���Mf=�s��R�A�J�����q���ڧ4��� ��%��c)x+m��3R<�qf
^��ku���h鐶YoW�����e��T�*�n��@���c�]2�j�E-#��X00�HvD�Զgc�&��Y\����kPa�9�{�^���C�x�)�)�l-I��T��i�29�fc�YIa��j�g�s]4\��qu��I`˻*ؖ
��7������,�R-ij�� �[	�GGKeek	�.�u�be��MuLD�|A��s�s�7�	m�z��Tz�}�|��n���|(B��5��}�0(�����M� ���nh���}Js#�'���D^�W�MЯ�_O�{�\
�����A��@���Qn)o��G�r�U\����ۡ@�����V\gHs��B�����J�kӴ��_�����D���&fh�s3F�2�{���}��^�B�}�ۙ���\+ﵪ�n���� �$f}Y��%{�φx�٠A9Cn�۟Sr$��@�s�7ay��CuW����~��Z�oG��mt� �yЯ�@>m�,����r�b`��`&��P����1-���򌢋�u�Q�J�]�֝SXz��hc�E�<��hs��r'&��_}x��;IK��_P�i>�W�����Ȓ7��
��q�-��.�,54{�DO�ޭ&���J������[|K�z�r�%����Ӭd�p�2b��Y�W��eXq�
�ɵh�n����7���� |��|��_}�+�n�û~�p$��N�ܘt�u�&�����'  B�ר��!����t:������A��~;�N�eV���|A ��A�
�n$��5�u�1��[�3��+���܋���߾�[��ԡ��|��?��EP֦HSd��Lp#�����B�q� �� ��QnV���ڙ]��!}��Z�v8>_
�	�РSs@�܅������	��࿐��M[���q��
j�l5��7��60�eU	��g���������̟[�cn�s����YU���|E��n�n>o&h���T(�Hn|���	=ѹ�U���?p�O�?�O�o�	}��߄f�W���^��h�;�I���!lU������=�/�� ��Qn$�<[s}?M�������Syjv�Oڻ����]�I��>������U'�U���s'c%�c���:g.�Uwz��&� ���n6�^�Ri�Űӵv�|;�ޯc�$rt(�� ����%�R��S��U8AȐG?���ۡ�>���~�7Z�gG� �k���5���俄)�\|3��I���!�B��	 ���
-�����p&�}�+�6x&���o�3R�+�|�=�MGt�����bm���K���L:)���*�L�+�v�V�i�R\f��fG���~�l�/�P��5K�Mu��|�e�;��9��ݓ��hTp��{B��M[�$6�P ��"��/�	�ޚ�;���[^�N�wwg]W�Wć/[�:=�7�4 rt(�%����������ɠB��O�@ۡ^-����[��Eq{s*tS���Z�f��+�|��Nw���y^-��q�#�]������ő��!�@�D�|[s^o�&������ܾ�N8�$>��a�w���۟������J�����yY��y��J�v^����=���]uQ	���l�r�)�Ƿ�E*�*h�)�	���EY�Q0D`�y/�����0��@P>)��7"A��^���퐾o�k���T>���ޏ� �����B�-ĐOw?^Vww��~B�L�@��HR98��Ge����]����حLY��TAG/��ۇ������E�4Cp2,|��?Z߄f��+����_�F{�+>����WHs�6�2� ۜ#�i�5qw����H �����I����_;Yo��W����Ȣە���+�2w�XcH�B�$P<�� �܉!�^���8L|����k�}�o��mPa�z����kz}CyТ�zKn|��ۦ'��VlL -U��:Cp'&�4���7�+V�k�|�|y}4��;�Ν��K���5����B�n'�͹�6�Qn>����q�>^��z�t��;�;������#���y:�۟Sr!��B�������-M+,����)X(�^�b'�����-!C-u/T��h�T��f��+"�4��������1R�"0��[��i
l�h�KHd�2�R�1e�3m&��h��k3���X�T�o,��!��X�5�n�nb4 ��q��f�t&��e6%���i�d�5�@J��f+�1�+&��"�ZJ��V��6i�V�4�k+�`�S�F�J1ee�현�b�h�5,ЍM�
�Mn�r0ҺZ�M*�ekr=kf����aF�L$�T��o�^��>����q�]��h�s�t�1�.��K�FĖ��q����Y��9�^�g޲�33SQ33F��c9�M��|ȧ����b$����S�S�͑���sD6����"���V�Q��?b��D��\�շ�ʡ%�-|/���y}>�wH�������s�������>�#�O|��ۡ^-Ǥ��]�$��&*�}�)�j���>
p$��N�۝�7"Hmרm �.����"|F�>��
�q��M�H�Ȧ��|�@5<�����~����L��y0~��6����I6�Qm���v���g�b=7"~��|����ʔ�Ȧ��G���h����쯏wP4{��'�Ԧj.a�Z��Y�1xȁv�����q��`:�l�XE:��mZ]Q�A�'��>r(� �总[��W�~��������A�{���HO���� �7"Hm׫͹�����Q��/�M{6�,MT��Ԩ�J�"�	g�Y7iK��k�%}����ei¯vP�]�i�jXڡ��UU�ۑN���"3����~�W�:�������E�o���A����B�p��Y�{7h��@�l�#�h
�H ��y�>n޾{��y������*J�&��_/����A�>6�Cn��`#&��؀���D���P�� |[sB�oLUpo}%���������2H�>�/�9��{�h��	���nhCr$�S���7n��~#~��H�;7�|>�G�E�o���MgM�E��Knm}�;���W_[h��H+�-0�4�
�i36�ʋ�9�u�`X�[nk�i~�[��}�f�ߺ� [s^ �"rl.�?m���U�4���}������}E�hqH�Gs�^-�[� �۟dN?0�ԌWp@�R�v�Rj���}%�������8�Iܝy�9�w�u'�>#s���:AnD���P�n��|�wAI��N��ZgG��֖'%�3�j\�0�e��Sf��Eqn�uk���lQ�}��71U�k�Qov��K$�t��u-�����T0ͦ�oG� ����yР[� �[sD6�����k��E�РR�|܉ɰ��?m���U�6�ñ|(��k�[�oW|�	����n�^>|�P-���[s^ ��P-�e.Ϣ>��gu�*���z�ʾ��p���G��$o9m�Cr81��T,r�H��nv�H��-�� Ía���H"[�26�a�EP�J�bu��5�] 6�Cn���E>�S�f�o����C�������Ͼ��� �nh��P>-���~?e��>7�h�;�2l.�?m���[y6���~����}������ɼ���P�
q'��5�n��{m̱�#��`�nlv���eM�8>R>8�O�rt(��AnD�u���O�C?t׈�H�}U�܌�]Q��>�\������k>�� ]��-5�~�}O�^Y�1����)�Bu3꺫����A+�Aۡ��J���N�!�z=1�������.']Y�;�0��d������!6R��tn=��w{8������ ������%�!�B�nc��}�a^H���Η��ҖU�k����������H!�@W�mК���X�g����}���e�e��j��3[�p:l��Һj��s\�4a���,b�:�Ϟ^�>z�!�}�B�q ��ۚ3�W��E|�c��|(�?W��\ �ʅx��k�7 6�g�nh�س��h����΅x����T�}���i���|&��F�@�W�����z|���<G��P �� �u��� ��]|B�N�j����?m����S_��P>?/���>!�U���
��27�63�e�T(�-�����W����l�c��}@�� ����a��I;��/�}C�@m��ۚ�7 6��G�gے����u#vTƽ�T,�I<q�Y�D�|�X!�;�� H���	'� 	! ����clc� l�p���m��o����� �1���o�`��� l���o��	'�$I(@����B$���cm� �1���6m��6�p�o�m��} 6m���
�2��Y��c�������>�������h �              @        |P3�*J$
�� @D�E P���  }*
 
H *� �Q"����U)B�)�� �R��B��
� ��
�D�T� �
$� � ���R�U%�2}� n��j��RX�Ҩ�D�d��ܪ+�wtQu��JB� g�RZO:�wH��R����N�#� �+�zRX�=�w` y��[� r� T)E� ϔ�UE )TU;�Wv���"n�}w�ԩ�	Yʜ��{eQ7��zz��%J�!�tҨ)B�{� ��*SMc�F�FI���P�@nJ�L�$�W,Ht� �(��Ц�5@"R�H(U ��5�Un�B�MP}nmT�o
*rЪ��è�ͨ���wUP�:+R�)e�TUU ��S֫l�������$�ލQK=(��Uu����$��UQn�B�V�)dUn7wI"wn���$ |  �"�
P�@I.�Q�UU�jUVcbJ��r����*M��$���+�IT��CuA;�$)����x ����j���P�w���ê��jBM��Tse%KJ�Q+6������n�=j+��  ��  w��(UUQAJC��U�U�ͤ����I���EG���U]j���AUY����A8�V�7���wH	(
*�  �{��R]�����<wU�W�އ�sjYj��:US��Lw�W{��+����Ww��     ��JR�  �L� �`j��Ȕ�� �    �ʩI�~�P ` �`L ��P%)I�h�2bi�M44�S�)*��S�& ���2�  H��)#@zMShj6Q�����<Ԟ�I��w�}��x��$4��6��,�� HHH���d� B=g�1@�� @��B$$JG�BBD�8��?��O������&��		��� HHH�B�00��،4BBE0����O���~~��m !!" W�.Ty4ԭ8k��A��
޾9��>u�+�op�����^��j�㍦`��T�*�t�D^ԗ*�BQi%A"/�t	���6��-X�V�ՔT�*�]��1#%%r�
V.֭�Dʽ9R�R@ؼ�p�M��n�慶�Zk�;6�V�5�T�?\�fַmP�T�M�i`U�L�����l+%aԝS&l�V^V8�U?��T�1(rU8�w�v�ӇTǸ�w[�6�³i���T�ؽ���m��eЈQu�c^Cea�圄6���*`#]Un��T��W��^ۛu�UV�K{�0��YÔ��ųp#5b�lSÉ�Vc���Q85����ks⬭�I�]�+Ȱ���m��hզ�Ȇ	BJ�*V�C1���j3x���Vnf�k&k
��7���xnS�y)lu�ww�.Zr�4V��K���wb�c%�]����1^�X�Xܭ�FT��L�Ŏ r�t��uP�J�۰��e����c��h���2��`�\���dAYJ�V����U��1ҽ����U��DoU�k^���9b�����dU)�/�I����ya�I4�t����QPᣬӠ�"�Բi���u�Dv�ڧ���f]�[�t4f���7^ns͎�6(�W�q(+i��\
�*ܦ���

����"��EV�F�&U<Q�In�	yA�{ZY�e�۷�ա��UZ��ܖ�Lu�ʎ�ڛ���&��Y�;#�)�2�.KU*�闫5��5h�����%u����+F�A�Qc.��,��c>��E�6P�Z����u����f�l�zfin4��J^YƋ�u�$�T)��A�6ڭ�Eb��;�cg	�D[�r3Lnf��i�!ph���8 5�w@�ɤԉʨ�uUU���.�v/.�˄Ǧ���wŵ��,)Co$7�N槇%�Ta�M�E]�YW�m�[�Lw(R�3/�j1�ә�t�]�n�FP2M��L#Y�Y��S��u<5n�Bn��UV*�.�r�$��VT�[�kr�T��1N�a��&�ɶH۽�+#ڥ;J�M�U�vr�kLm��#�O,�Em�D�51����dș93-:%).h�0�P��y-c�6�]mн36��8A7Zܱ���\��qb�����̔��͠�ۘ�=��h8��#5MZqVD4�!ks0I')*CqWճ��:�� �q;�s&��&�V�7Z�3XQU�������C���2�dzw��J��vR��B����vmFœJ�������ӸUIG�ֺ$c�wp��ΒMkܕN1�����kk.�;�z�X�#l�p��OX?��8e��T�,�Q��k�\3~�YB����"v�Ua�aׯC[��ʓ6�M��i�ݍd����mj��sZס�]-�ۗ���X�ڬ��~'tAU�Wx)a�q:˟%�XHSV꽘*k�C�h�[�ը�����Օ�To/+L��	�.�%��ݗmҤ�,�+wf:�X֨���p9���R� 先;@�ۗujK�����F#i��v�m����.eF�����.ܛ0�o4m 1VH�nĺ,PJ9y)���Ӭr�[���y�W�V�D��W>v�Ii����b��6�X���L�kn���5�x4������ڛF諪H룙��ڹ{�^�ɐ�V�W�V�jݥ{���;T�	����č�]�)��c��8�m�]F� �P9B��P�v(����H[�'��CU���5;�	�f�U�D���v������U�#Ϯ��N�s.Ɯ8��ҵ*b�)�qhӶ�Z�td���%λѝrUT5Qڕ���Q
y�$��T�RV����[q�4�F[Ŧ�Qw��cv���,�������ɦ�jA�0m7����)�Q�HªU�؁�(f��I�h��I�;y�[��Z�1T��wF�9��hEe���U�í
s��v�ЂG0�y��ݷ��(�'+��k�wy5��1zFe�S׆���h��R��"���"��h��-���kI,j�q�ڥ*e'Y$ŉ��MYg`ѷ��IZ+�6��r^K&��G��ho�c�a���ݻ4�1��Mz3X�\.|��ܻ�5IH�d2�:n��#bAWSe	�C�d�	��[��y�X��/���*
��A�e\�q�S%�Rv+fK�8��Wcu�F	�Va&���5zՔ&1z�4�!d#n�M��W��^���"iܨ*���.�v���l��*+��}[6��r+k�wN�Fނ�N��nӧ�\۬�N�V1[r�U`� ��B��k.V˻������"쒴��:6LW�=��#e�b<�[�NJ�{w0�ղ
�ںs����x�����E�6��ݡL�Ȋ0Y�����5[������:`tK�5[S[�'l�k׳g���j�Z�f^�����V*XM%Q�����&��[�+?e�n�겞]]��Z֭:��It��R�֍x]+�XV�6��m氨V|��¢J�Z��Ra�'(����x6�"-�*��7��<k�in�90�d�d�:�Nb�,��2j�ʩ�.��[6h���9����.e]��1A��CCI�����%xl&�F�P�{�p!��+��jK��nZ�V�ubnnAv�;hC�G���p�V��_8�b+Uۂ���v��wx�(6J�U���dX�Mۧ�i�)L��Ju���JaЄ��ڬ�TI��77	7��١J6Ӕ�%���*�.ɔ���qg�Mm�e�u`�V���謲�����UV[x�)hkr�j��^<�p�U�%��e�̳���"J�a��Ss&˅�2�ch9"����f^�ԶX{���f),��U҆����.�$�����;��n��\�m�A�4��Jk%e�M�Q�P8
wnm�]��Ӗ浔u������Ҷ�ޭW�&Q�n�:չ��<�(�kN������$Poj��m*s�*�5�1m����˨^�y�VM�A�X�RP��Q-/kZb񍌽n�.���č[�rǏ.�V%��F�{��o7�ar�u�[L�id���K�[E�A(͓H��l�U���S5G(�h^Lݥ�)�P����q�D���+ �j^�*��t���v�rh��%�qn�cە\H�E\�٩-���>2��n�����p����X�V��,��o�ltԱ��ge��N���6�Y���)��ܷ�V�U�j���',䭉���2q��JRٕ��MG��sF1����B5T�[�1⳿W�-'N�T���U�e%�IY{��8����,�'d�^�b-�%LW�Q�vQ-�e�a
#ǖ�X��ޝ�;�R=�j༖u՘r�G���]�W����E�
��PO��]
���$�'2#qǵN��m�̥�Ǳ�GJ����Sԥ�n���v�l��t��+��ͫ�0�ӛU���[e��0G4��;q���;bֆʛ�L�u��Kr�����&�/M33R����K�@�Ү`�U�&=¥c��Mh��^B�IVF��bD�v��.|��:$&���N���\IV7�u�`�ŌV~p�ܱU�����d�0���Te$����,Bڥ4\�3r���/F'4�4B٩�D�©=YW��R�YkS47%�e[���U!�˺у�%�GA+�@�ٴS�q��:��bV1S��Zz����ș�k#������XP�a���{y2k��4cnmS
'�)���y���܈A�X�n�ˏv��	zB�$CHz�T�Vb� C՚jdӶ�*���aD2e�3.�)J�g�e��yTƲ.c���1�ce������ےAug)8������35f̪z��� ������i���[�aA��:���٨����Gk#[%)��W��wj�cԌ1�(VS�[�F��j��d��Y�F0v�V���ُp����Y�WA�'�]Z_a�.�7��B��K8ۖt��2V]'M9�6�%��m�ݙL5d���f�{�	�����"��d���_�o^�,P�3u۲���M��-�7؆��Ӆ�b]�f�T�ـ�������[p�+F�U�
u�u�nĉ�C�S���w�wV�UF�!U`�h�_[j[ʛ����;pTjT�B�[c($1�h�q�UH��W,��cX*ַR��y��QV.���	`ߩ��3;m�b��]
$M�C�W���a��XYc���@�p�hź�����ܼ����!Gv�Ecywr����Uݰp��T��286���}s5��-x�n
�#iU���Y�D��MZ�ms���y'k��a��.Z�nF5�t��Щ�q�ċ�qf�4�ݦ��i�˒}.��U�2&0�eQ@�����NTx��<�z���bPk��mV�g��J�Q҉�M0i�aͩ�4
�:�Y��"��Ӎ�*�.�I՘�v�A��@�ţb���Y��V:�[)}z�ِn��P�����١�,��V�nT���B�C$V���JK2�������30��/��7[�(d.�l�&u�t�h�Y�G�;�
�T�=�oFn�.��h�V����&&��;c,�#P�^A�e{o%��)L��ۼ�l#5)��u��U	Ain0�l��U:�eZ]m��w
��{yf�Pe��#4'�𪪻����gMՍL���	�U�f�{b�l�D��
�r���r�BuV)��(]bySt'uw��^U��8�LAl�Ӧ��0�Tݑ�+oQ���}��[�0��*+���i�ڣ7.�Y�ek�%�·0;����׈+GV�{��)���g��8�ej4���&iz�͒��T�-ݨ���"�a���7r�EV;ʬ�-��u{5�U]m���L�;SWF)�XQS�HX�+,\Y���*Ji��r�CRK`��R��Z��B�S2`�	y+-�ݽ5���խ���D"Y���Z��],�D��.������Uc
�5��+xF3��i�[�9˻)VN�e��7�fH�m7vk0���d߱S�ə�G����Zڷ���)��0P�.��B�^����*�%`?iŷ��[�W2e�SU9r^&�!��\��2��۸�n�n蠉�V�3�d�*Sö��,�]h����]�ՇmӠf�[ILZ$6!���A��W��*�ͪ�F���c2BZ�n=�mm$�Q�Ky$�X��E��������P�yP�]V�(eUT�j�#��H����R���N	���3�d�đm�:�K��~G��كL���zݶ��x�I$�<�$!y��+��+��;��*�;��:�㫮���:�軮��:��*�ꎺ�誺4��I!6��M� !��Wu]wQWGWtuQq��wu]E�qu�wq]wwt]��t]wwW��U�wTW]u�U�]D]��quq�u�]���u]�IWwEWqWTW]\u�w]�]�Q�W����U��]�u�Q�]�]��wwtU�u�tu]�]wGu�u�wUtWwqHm	%�����Ѿyǲy���� BBDq�g9  G�!Z,� �		���Ǐ{���3Ss���yy�{����x�A�ͺ�SE�ui�b��l�_�����R]�W}QT^�YV�9fH�F�e���㭬�����V6�QD��Uā�ud�y%'uój
��۾.u��%2Z���ȭ��O�n��ʻ��S��b�`*%y}nM�ڱԍ	t*^�� u�uv�lf�ۼi��y�#VsY(����[�p��%5B9
��ԷT�D���;�c��.B*#���4-d:H�Vj]�2��uN�`w7y��F�g&a;+����9��3)�W|�i�a�T��^p}�*�=��W,�q�n��ڹ��a5�M���E4�$O�S��P���g"���M[D��/�:�2�yX2������l��?�\�������R	&�2!�02�ϝ�te	W;�PFꕩ�Ն�P�R�NwI��ŵY�Z���=]��������Vb�����Z�t����X��}"�=T��7\��M�+��d�$�Q6��n�j��V]9psҢ�T@��l��T�S
��Scn�SB�4�i��b�P�WwI�x��RUN���������M]e�Ք]+�y��(Uї-rm�,�[�n�ۊU���Z�-mV�3��4�Ui�r�ԭ��#yP��7a7-��[PQKN�rk�]�wb��UF{1��Ŝw��w a�S�)�ɉ�VڔT��Kفw�ճo��I]�y݆�mޥ�kfU�h��`�	�i]ȴ.���7��*��M�<��
�޷*��Uu����c�^:���wn�v���@�u]���d���Us�6�9�̍�.��`�X�`LnгE{n��7�D��Y-=�W�5ir��*1�-�&�_>���XUU\�gow:�N����Vn�k;ה5c�MrBm���+EU�wgbG�KYt�����N���E7j<�e�Ԋ�wYL�D�Vv��F����|�5]1Bd��	)c�m^q�TBI��9{�X�l�Ne&P҃�|�UZJ�Yìc�iu�[�gJU�}c-���h�n���70�sUC�W�㽼���ܝ]���J+F�t�x��#ʢ�sr�qpjunU�x)8�jC���ω�6w`���C�$.Ƭy�2�]��]��r�^�YR�_M��˪���Cήu]��vR��ŕ�ncQ�tξ��N'��Ӱ���fr���Ju��97�ݽu{YE]�S�L��;�9Rl��{YF�S�]}0�gV��b���`��n��.�Z�!��e���.N/�Y��p�Yܳ�6���{�i�q#���e�p�U�o:SKq�UÓe�b��*�>.@�-VFi�8S�c�-��.�͋���g	��a()��s%%�V�mm١��A�Ñ�����;HӬђP\p��Uέ�hoB�z&Z|���o_]]e̬'�m�eV>v#��d���ٺxs�qL�t��f�G���v0R��֠i>�I�]�,s�#�e�Yt(e�"���٨ݧ��1iH�T���d+ouنC�t�c"^Rz�1��ʐ�D�*&JHj��	dJ���X�0m�n��Z	J+,aB'r�UP��8���sK���wv��/�,���q�Gc�Q�4�Y�m�`�kk,�P�r}��f|�Ar�WYm|��X2�l��J_e�'�b�Fvrf�S������k�:3]Rٮ����&M,�WY�۲��l�gV)�e�MZ�Z&�˺WI��o�w&�2�����ڡ�3��
ܸ��1����5LS[0�P�UA�[���u�c�BCHr�X���r�ٮG#̦�a��[�������fUӅXi'P�vn�^_</;�Qr��³0�R�D&�ou�L�t�;r��d��b���k.O��n�)*�R����բۿ��L�����z�z��	������!L�-�!��R:��o1���\����+\��Hq�e.���n�u�(b�����a͕W{UK/�$j��mrc��MP6kS�̕�&�55r�5N�K�*�0H*�vƝ
i�����U���p,L���3;ź�oe
S-�juC�S瀾݇e���2���S��gn���v^�nj�Ȧd����N��N͕�=�u�h�	�O��G��8*��5� �57���6�ռ�B �s3�uX�!�Z����q��"�*Q7]hn��� �1%&�N�;{�Ӝ�7:ͪ�9�N���CJ�'W�nT/�Y��f�%S������8�TQ`��72�N2LX7���ű���]�P[��#K��poB��E��'_5�m��w{��O

քs5V�{�{���O�����_L�^����};c�bp��e'SkD�d�Yһ�R��(>܌̚n��([4F��f��6�@�#i����ì"�=3�]^��]�.����T�q�m�T�#]VLȆ���UN��ɻ�cr� R1�nU��3ꂍee�}�wiKR�-�a�I7�4��.M�G֐y��u8����ٲ�1M;k�i�����W:^��!H�^��{�C�x��u[���ݮT�B�X/h�lv�|$a������!��i��9;�^*�T�b�Ԁ�J��^<q{Wpm(�7S��/5�(�ג�A�L����S�Ԭ�;u�76S���,Ք�tu���Flt�E��/�k�Q�}w7��}����(���}KwR�2��A8[ttL�����lܬ`b�ѭ�x2�(b�5�l-.Y��,���Գ��+��͕ٜ���w[��7h=�9�˽��Bk3�j�vneԫ�i�e�f�Ҵ=�
�U�#J�D��_�m�4�1+��je����!ul�����!K��ô��%�)+l�ڬ�v�y��Y��C`�;��Tl��m�{�]��wEY�Un���ɲ���}x(S�f�����E����+U�)J�%u�mu�3�2�kQŖļ+�d�ҧhVU�?]ۏ�ֲ�6v2AJ�51Pw��T����
��H�"�l���)�Z�;&`n��!>ٲ�Wc5�x3�p����EayP�N�V2Ѽ����w2��}G� Άl6W�w�ye�(�reZs+s0Y�����e뺱;t��}������|�M����7�m9�Z��������Й��v�P�Y������Y��6�&;{�A�ZX�����\�K�N�����}�l��YWƸDVC�4���4�U���b���B�p�}|yf��r�����9�L�ZX�sK�ګ{Hv*��`�BuT�)a9W���en%ݶ�ڦ��Y��N�a{F[�E��N�/�M뗤G՘��]��/6���v���j�K9�qAjnݼ7�H��Ѝ4IĕuX�p̖�K�̃u �&X�[�����5O:�_U�U�7[�0垭���ݭ8-�N�W��T:�D(���2�Mk�Kn�U�p��ƖЧ���!�׋oK��1�&�E,�A��4�]��<��&�);��E�1��m1���1AM%vt;t�66劥����P�g���u�Ē���'v���D��iQw�*z�Eɝy�f���ꋦi��6�]��օcm�;�,5���w�͙b�u�ٜͭY3iER��\WT�kbM=&fEx�D+3�8��Vm}�þ�y �x��#=-M��h��mt��Nk*����T�)qyɶS̜�53ben^�wVi��]y��4mO�l�%ݳ�f��SWu�buVcx�������j��61��}�6+kb�y�͈�k*�-ц�W
�^u�(�R͸�Z�(��	׽[z��D���T���D����Y՘��ܼ�;]6�_]O2�Ͱ�m��h�f�"0oL۪$�ۺE\3$Q�Ô��9���.��1nݒ�E�Rh(6���7@���w�T�	����C��V;�����/*��77��;ox���/�g����LM��U�L��1V�M���b���j��|�����:vU>�}5u3 ��b�R-8�A��ؖݍ,'�o:�;��ܻm"*����w���,�)�ܻ���N���Y��iyf�mV�`Cm	��s��ګ��[M��P������z���V\�A,�!	��wUW����C�0* �n#�i���fIU�j\��<=��F�m���{t0أHs�#�(Iͫ2��2Ɲ��6�6a�1���RdW36#v*���A�ܭP(��
�i�H��Ÿ�MvVnq.��f��
��\B�� ���كy!���b�1�n�BM3�B��F��ӳ�&MX���K��p����R�T���׏n�������\���Ƴ�n^��}�&f
��w�P֕������_/��ך����S��ںPϷ^����}W�Y���ac�{�J�W�����G\�;�F3�lQI�,ZkM����S�X�+6��Js-;����Y0�EY<}�v�4�M]f�7�%dT��2i+��b�bv�]���Tq���c�$Ùn�=6c��Ab������9�
�׊�fZ�&t�W���F�mK*��ks{*��C7m�iA��Nų�nؠ��qT�������u����*r�Y���׋1a-Wo�ެ�;�܄%�Pֺڝ\�<�G^n)�+�LWJ��}^�2r��J�ӧ��zv̲�ݐ;H��S���լ�c��j�R�c��UT�w7��V���B�q�-�dꫴ�z+��
7v�uF�����Y���嶙�v�Wb�v�*�T�q��a(��mag�:� ������':���SS ЩӮ.�;O.�PبFA�r����LR�S��,!���&�wᤘUFyK���;e�I����ʱ���T#+-���J[��;�A
�+��6b��}|ڼ�M�2*u��.c����w<�QYד�v�9έ�;n�=ɚz4��9�T�5�z7hc9�:�#�bbTBp��M�3�L��������[aY�\-�o�%v��WƤ��xK��w:���uo�fYw�����5�-�-��ܮ�ۘ9NNU�8�e$��׆cKl؇mLʊ����6q#�hK��Ɩm9$��,�+|�����)�$9uRd�u*�@���:ѪgqY�Z��-����PM�e�*��,і;U��NK��uQu�FJ�*�SZw\E(HK�:b�YUb�Q����Y���ˋ��w�w굤��v%��c$Iګ�4N)U˗uoԈ��+��R���\���7��)؇�R�vouy1
.�@�&���o��m2��U:�Fe�r���	�]�t�5Ɲiu���.�|�(:�WU�I�2�(!�B;�LH]�4n�q�o����Γ+s�s�o��FΠ�(fQ�cp�v���%�Q�b�����5�	nޭw�=�� x{�C6��4m�u��D��(ơ��?�n��є�憵3�-6�I�챸�kc����KnJ�!���N���Jd_q�ݹL;f�v�Џ�'�c)'��6�����۴v�`�\� �c+O]�A�mt�$`��jlѸ�:�r&V�n:%7,�}<yM'2�i��ў�㍸ug�u' �'۞�k��2[vcq�a�3�y�N�q�4!�8��$tOk�Um6���ێc]h�F����z�7��n�YJ�PKBj�1544����k����=�ou;��i�W��Rb�Uu��O�<�Pֳ��h~l�e��z�gV���:+-�q�e��t����qm�Vq�sZd�v�n�	�6�(��pp晔֖�=��zJ��v�A۶���PeѮ��-�N��mYk���F����g��q�$U�4ƄB ����BhF#讘�zq�M��Kç�Ź�J���)]*F��4��Bl$��yl�p��u�f/Wm�wKlQx���tYlv�v:	J:4%vkm��R4� n�9��g8���:���7[w2�r�ps�`.�nI�H�ѽ����
v�0ـ���N�e�mZMh��`(�KWT4e�K�-,)�'�uk�6�����gQ�|V,FI�\��tՈ�b �:����`�s��
���탎�v�z㺂�]��Q�c��v;��´y�a�.8��}���u���K�]1�GiE|I��$ۍ�IN'97wi�CC�0�zz�m��n�c�J��b����f��*.̷Jifmg�z��ݤqJ	���[��:��Y��d���k�`0ۊ�71Y�K]�P0U��3��'B�B��z�K��ۡ\ 8m�mh���К�jH��lXXj�k:��Hu%�5�Ĭ9�a`XK5��&�]��p=��F8ە�nʵ݌�1l�q�G��	YkA���M�fÔ�܌q�5 ���wma�mvm\�B��*�G� �x�]ne��+.��.)c��Z�:h1s�k&����#s���[��`��!����ˡld�,�ֱPn%A���p��.)M�SU![rRi�6�[`4���z�9ɤ���8��j�긱����";k��<�=�u�bz��m�tPv��.ҾVQ�]��zz�an6�m�6 �Pc���n��p/ �sV��T)�s����M�������X=��Y�gʃւN�<�j7���ztq���;c79����Ѹ&m��2,���X*�{�����ԡ��t�:h!qqP,�˯��خ�y��'��-hn��Z��k�h�xxdfkt\�j]�B%�X�P���I�#��Z6� ����vS�p3ۏ+Ѭ��S�ƍ�0&(ܡ���r��PԶ�S֞*�ŕ�ݮ^�����[7nMm�8�'n��/A��Oj'X�ڷ;��A�J7=�����k�0c`ݹ�n��Ī����yr�1M0.h�;X��	*Ԇ60t�+�KVb�X���)�]6��k�R9K��i-0͸d�J�i/ n"�鋢:�\�id�Fi��m������h1V�� `����':��j�sҙ�{#��J����]��D�6��4����'P�9&Aی�8��Mv�Jomv�L�y�%) [�Y��Q��2�bRkhmbJ���SZ^�Z�E)��ZX@J�iWe�n3�9�]�xx���һ�̷Ms�Wl�n��|}�#���ۃ����ƍ�\�佐�y���5����K�0�iK�(8�N��Oc�w�Mɸ�.kô۔7�`筯<vB6ii�I��.��R�6x,%ێ8vy�[�7M�]3�����l]]�KGn�to�ӝT��^����ρLy.��#��GpY�f�0\��n٦=t�,*(�iv�f���yA�L�B�XAMt�v�l�6��ǔe�0��A��:�B$�i����K���ư&šYe�ִK)�[	�k��nM#ӷ\��oZ�,�sSZ��c�te���N�$1�V��Mz�<u���[����c�sj��`�6x諈옂�ɶ2���D3�q�&�D�[q���{O�X�v��h�1@�f���Y`鹇� s��I�(;.]x���t�4���w�Y烇��1�W��u<��\���<U��7K%��l;\����iOn��u�-@��[�kq�r�l�#�g�<���`"�H�S��>�s�����\�c�-�U�& �s���k��O�<lٺ�7[y���mq��\C�ˀ�9�n�l/k�����v/%=�G�/[6����g!�"\�u����S�����tƃ�R�G
�Ra��[�#֎<�x9��˅��2��%ځl!��4�Xb��ݺ�7R�5Q�[�ƶ\ch0�r��T�nM��&�n$�޹�'GX^���]�m��z9 6Fc+��2�
RR�h��xA�����-��4�}��Ō��^��v���*����nJ���<�ɀGe��4Ů���٧�?7|�0D�a�p-%��5Ζ«[fC��[�N9�{-�ʋ�f���['o��n�0��{=hμ�͂�����`�l-�|�|��v�u���lG'r$��YK���x�X���Ka͌���H�9�	��a��E�6M[�G5�V��l/�������rR���1:k=^9�H���L��c�8طC�պ�s\����A��$�#D�1h�2Jtpp6��y�pO�ڵBY��G�����m���nk���a�!�,
K�D1�Yź�۫�f�'�8���'<6|��u.t�'n��4W+c]��=Ap��2ۢ�yb�q�-�X��결m��ӫ��q���gn�WBnoJ���L�8fq
l��@B��.��+��e������d�c��Bb��ͱ�"�%�H9ޜ-�����ě��;k[����v֞����֮s�hm7� �mA�L���c�D��Cr��e�<yyџcӁ��M۠�mn��ֹ�5A�y�m��]�n5�m����[\�� ӄ�"�T��5ܮ���G;9�^��A�p��5�Y��Y��gK��!.�,F�Q�t�Ka{\��î��w`V������ώ\�A����X�45���í�k^a���m���]<Yx k�N\b�8��]�ę9�ܜ��r��NĂ\v��0PV����zcq�wC�Sh]����--�6���NǮt蕲�P�j������G'�{pq&"xyF��Tۍm��M]E�u�;+�p�Dηj���m\��<mFoGZn��`�8�˂gs��a���k���5llZP�瘕i)=r$ݸ�v�S��]�u�鶰��o@�C�''i�u-ل*V�vj�P!�� ���#�hqƻ���u�G����ޓ��PX�(��w8�1����3�=���%��F����QL�\��:r{])�<%�.]�}�����iB0㬡�66��D�򻷛����;����Cu��'N���K�
���� 5ٜ��D�۶8˰ܢ�K��㧘�H��H�(`�+,74��C[af���M�=v�<K���m(r��U�W�SkZ��Q���ݬ�uk����f�3F���qj�Ս�m��F8v	�IH������0a[��I���>_>�6̚�V������Z��Q7,ņ��"���h�e���lsR�u��O2X5g��N^ۖ]�2��Y�M�M\�c{�s�^[:��ݖ�h�#�:G��秸+- E�������e���@��u�4E�9��G9!��a�Y��^���<�8���gm�$�5�q3tfH��yĜ,��m���6���jDC�m��rYd�G6+y��;�9{X��r>ڑ{X#Z�NYf��&�n�w�8���� !99ӗ�˶�I�Nw�hL�J���)��m!iH8K-ȕ8Ҳ��p�;m������g^���kti�Ys�qJm���=��9y�sc7պtD1��M�6�,@*>S��&&"h�� ���Lj����I�˭��ݳY{Ѽ[&n*m�+�n6YM��O�@ֳ�yLѰ��zѸ8�i���5��c�q�Aø�^�x�uv���{A��h�Z��6��q{m�J=���`cHp&����6J7e��_f�G[�cv�	�t\nkqe+a���e4�M��v4[�t˗V��ƭuwGYz����U.��Sh�h�ʼ�l�]`��Ik���ٻu�+����q���^�k���G2T eɇ��@l6���]e �<1�X�A��'�P�+w&�x6'�y��fo\�q3q��v��g]��;����{b+�����Y��<y�ܝҷ4<i�p�h�\P���q�!&�K����A���]���v�<�ؼwmi�mv����\��8㠴�=w&1jBj���ٹ!�cUT��	+�=���u�a�&n���2��5jr��X��<��3Yc�7on��4
s�xc�ÓZ� �� v�pM�8�)��b�B;�K%M-�%K�C�L���\��3�u�;�ۮ�. ���\T631�3�F36%Ͱ60YX�
�7/+&���q��[X4�O�
�7N�q��I�`狓��=[d �8�x���c]��Z�.	��+�Aڮ�g�'L����q�����!�Q%�r����!A1��W9qv+���\݇��Ѭh ��M�$� �&��wx��#�Gn��aƼc)(���R���R�K[@P�R(����e����V�,P�� +`���۸=�*��xC�l9��d9^\�a�� ��y^2�TJJV�@��N-��W���������t�p��^���t�]�k6��ڵI����_�Q���ub�*�v��b�����D�dO�����Z�FOLܚT����o���o�ʏiy�E��򻻻��v�	\]�P�[	.3�����w'm�O%����E�{+��m�j�y��
ʻ�T[�;��̯Y𻋺[��]d���Aes�|� ���wO�"�������j;��L9�P)�X�2�B5ҋk�=�}�ν�����zR\d]v�f&�����,�Ǯ�}� ��*��e|2+�Zh;�Jf�,��:�ܬ�%W��g{_�R�*9uQj6�eL���	���w
��Q��otڞ��dy卑SYъ��d ���<-P�T���s}���x������Ц�)
u��-݉�1i�M��(<�l�o�B���y�3��2�d��-�({�����iT���,ݛ�m�Qڟ�l�"\ݍ,f��]�qKk�l[f��p���������u���s|��x��CP��v2��G���F�H�ɩ���W������?y�Z9yW��1|0���a���4,�s��Wt���b��/��9X����ojj���T5�{j �=33=��#�٤�ODN�E�9Y��zU<�yϮ��T�ىԗ�ͫ<����lg[�}�	������t�|.��׵��Ӊ&��SZ'�����w��E�^ǈ�f��:�p}��3��M�0U�W��n�k��ۇ�ze+��8ws뽬z�k�꧜��&6c=��'ً1�}�u5❍�d���\���W�Q��dŹi�i�8qd]��ms�V��;h-l��{��7q����'���w@����H{�q[��=��=	�p�(tM�a��x�����3�:[�N"�s
�U$z���Sس�^�7��)��7����3�3b�k��?y�ܼ��}]��������o$4���_�'`a�f�ט������a�l�cCchp�w)�1��<����e^����e�Uu�lU��u�"���̶�]�����+��ⷝ��C:�e9!x��1̪��{������=.�;*=�]�в�N>��@n0��;�����l��yyd8A��#�-��i�2�g�l[t����Ux��{:+y�q����v�6.�-��-c�����f*���ٺ���18�}�<�"j�͹ʻ�-D�e�+���B!B�}����Zi��WZ^l��Q&7���\��3�&�8��ܱڝ]o=߃�|�����Q�J��/*vl�K�f�����,��n���%9J)%U�W	T��,,�a:�N�n��b�;z�I��F�;V�B�9�2�r�yic-D(n9r���߾���Q�����6.B��;=�Zv5�C[dRqA_w�"=���,�Ԧ��==.�����v[���3c�qd��+�4�b�y�k�[������f��2pܟnǬ�!��<��u|�H��r.g?�C�=d]��(p�Y�����/c�u�B�k���y��t�ٖP�{B��z�,KQww'�=/�itM>�7�ޒt]�l���{HE��H*�PF��T
�M�f�\	���l6ل�	b͆�]R����b��'U������`;n���#���E�b�Sދ�S�<�7�U�<��
�U��,��7I��p��O*n�-;Wf��/���oz��*� �>���a��P�ڮc��geG��qi������}���geީQ÷7ge�-���I�Ϯ��x���FE�f�q�%^�2N~ؾ�z[�-�F�̿�31�Ź�*�����'{�~���߾v�?f/�<N�ѹ����hM�5��Q�����lJ��a!J�]Һsb�X~��^3��p�i��	
��cH�Q뻑v*\�9WQ��7�1=ĭל:�/�'۬��܃#1��{�&Ϯp���^|љd׺�`�d��rɫ�E:3[��;EL�v�7�^�7��Ʈ��]��j]ǘ����	�9��w��ڶ�O[7��g 9���T]���=f��>̊��!U�'d��bha2����g��g՗21�.ЄФ[��n捵��4�Hȑn��y]�^ί:���ޅN�GC����s�s׀a�Y�����݉��-o�ٍ�/g}����3�^_��;O�2��6��]�ڷC��w5��=ĭל\v\���7��g��|�nE���;�]'�7쵐t7��u���`h�4���>u�tvwVǢ��եP�O1�%d���x��m���T�l����>����kA��3وg<�W��$�/����zw<<5�7�Dw�bS�$�W�쫤�X۝ח���Z����m�$����$�]Ѻ���㘆d�y�j�x����wE�u�9���,�D^��QT��t*y�Σ�^u�������]���>�wn�%񽺅N���q+��%�z�.�Ev��|�f�z��x�a�+u�W@�J�n�ܗ���u� ]�����t=}�Orۨ�W��uM�����k$�U�o���f]k<jb�+r�T)p'���|�z�c�L=}������;���F�:�lЁ�P=G�mÙ����t�_X�9�-ۮ�ֹ5�`���$��vxm%6eĻv�ݍ�����;H"�h�4��6�iJGm,�z2 ���;�Ny��<���<p@$�ӱ��s�65�ǻm�e��-F��;��߫��Yp��c�e;k��ӎ:.�]Ł[�Q����P܋��{�S�V7��a_O_[��U�F��Ø�Bd�8��}�=�<��{������y��l-������]���h�[��{<�V�^�M��]G�����nLԥeP�[T�қ�x:��WztM-vh��'[��w Y�)���V���u%����bk���睴�ގ�|{N���f�4ܸս���ax�@k��mv4�Dɪ�dwu�9ڕVv_3|�3����g�s�3b�=K#�Z�t穠y"��0VU��H�!˔nhۥ��mT�Ƶ".�[(�ț���w�
�u��#�W'��g�LwW��aj��s�1ySf��z�[�{Ô�=��d]�ګ�u(�����-G�ŗ۽U����:��u l�q1NR�R�d]���Yu2N�I�8��j����1��p���f^s;�ϱ%H�
�2�b�J`�40X�&�+t�JZ�h�R�K�=��}����Rt��f^T�1�� ]�о��ٮ��b�{���v�|�2��0��<��o��tp�}����l����~U����?,��Z�������S�ܮĹgrLKgT1:����1ڽ������Ue������+?Y�ު,K�\��-_3�nZϸ��U��U�6��(�ӆ�U�yTIZ�ٚ9�&v�й.����Ɍ�Ƌ>1�E�gh���_��㘟��7�Uc"�U#�"\y77kgL1������[D��t��@�N��γV��Yw8Ȇ��6�Jȭ����9W
�\)��Z�SD=Ks:lPJ�N�]�g�gEf��ݡ�2�3\���DMT�q1�,(@1&\�-B:�'��l�f_N2�fuW`�ʻ��<sNmv��d�]��A}z�9��{+cs��f�;�n�bP��I���캙1%f��F����5E��d�D2��Ȳ��X�ver	�:�����2���xmf����u��z�u]X]�p�_fwt��%T�j��7jAP�+v��;�]�i�5Kj��++�0����Z�up9�T�5>b���z����}Z`�Cl�n16fќ��k��Ӱ�D����'T2o^](�n���ǜ�{�Y]���i.ƫ_I{bs�Ga�|V�k���ej�oM��9�r1]B��jr��f�����{	�d���H�X
�I�$�g�{Z�Y��ygyy�$��⭭%�,�	;o<�!�9�l�F���"H�I�<��%m�Ok���[q�/l�{`��m�{�9{gr�,n�-S��u6�/.�{[�BD{imiȉ/krvٖ%'��j�^Y����e�gr �$��=���݀E6{��$�dRk`%�rI�͚(p��:��Y[;r'I��iȒfH�@��]Oθ}]�[��}�qwr��S�ږؼ˽wv�4K��u�}�_G�0صF֐&ky�-�����{�~��לߡ��&���f 31��=�<�(�������m�;0�X��o\AWt�����u���9 f5잶=o�&w;��^�������ffcl����É���h���'O{���;�u�t.�i𻋸��Ⴋ�g]�^��m7�2��2��]+Mkؾ���ܝpz�o+��/0����\}EFd^Q]�m�鎪Ȳ)���
n2��
�V�ٽ�Բ:ʾ
��Cs���&sوfd,V�Ac[�V�<�
��}��A�>�}��$�0����JD��A���6�cr����E7q�ЉF���;��wt��7��_Y��2���<�t��;����Z���n����r�]hy|8kw]�#��{��n�F�Yqvn\�Q՛��	��[�tǺ��ً1|���Q�v���40������c�]�tb��3��c^��n���.�����-dF��kp��5������+P4F�r�^����^�s]Ho��*�=q���r����o�.�n[]诹׻�����o�VÉ�b3�2�!��4nf���PnvXm$G���x��՘�n����;\,�U���*�J�$�F�e�4غ���Cq����$���n�`���qy���0��{O6�.:�=٠�-�{����簜u���H�i�{��~��&�̱K�d�nrX
FhsFY��+(k�Ri�Ԡ2.�]�k3��Cz��}7�xw��b�˘c��ts���Y��2���n�GV(�T��x\�ʥd]�y5Z5I��kyqփ��I�]���J�ߌ!l�Ie�f.�o�h��-���z���vD�і~Vbs3(��ث�Y[���Y��R��\�Ř�~!��d}��sk58`rf���瀈4"·�[O��o{�����ޭ��w\k��l���yww ]��̍��!N���}һ:��P�q伽i�죛6��4�X7w؅R����9u�A�B^,:7Z���h���G��<�}q{�^_�u}c{�0; [q�1�!Z�f/����ݚ��:Ǟy�3}_��_C��fT
��S\����OJ�}��N�$�A6���F��tq����f�
Ovfy�=|����R�y�#:z��4o���%.��w.�dŔ��㖪'�q�u��2���_f,??8=����=~��ht�w�f,̡��_��]P����ɲ߫��rwP�����Ol7w7}�E�����;`j�L�zr))�"�m��h�*v�J��_x������(��cvF�f�.���x{���5�pu�U����dY�]�bJ��W����繡vn���=ぜG�K��e�Ok��@p���)�4!�P
ZUD�{�b��Wy���� 7�iQ�uQ�z�P�@к���@P��0����Y}��5�*ȴ�q1�0ޑnM���Gs[���8q������;�"�U@�*�@^��z}�a�;� 4í�{ۚ���UB �5(M	a4U@�T�%L@c�n����;a4+�)�a����ַΫ�������hCL
����
���p��@����6�Bh7P�&�P�L4�*� �����3��y������o�
� 	h]hF� �T)�aMU-�^9]������ nj �Bª����F���X�����H4#ݟ��_s�����L?�m��*L��7�h��i��dZ(A���Ĺ��Z誵[����_���	x7p�*�2Е1U �
� �o~;�Ѝ�:�x�uΫp������� ��b��6� ˋ��ţ̬jҳB��6	�(t�Ҽ��nk\yX���&g�; ����+��KM��	S�V����M�}@^`:Њ�k<楘�b3 ��.T 
b����RЋ5�nl��]�*��q4,b���BK�]�do�}5��aщ.�KB��,4#f����#m� ����KB��B�ІUJ ��2І�S@p�gvFv>!t]�Ϧ�2qs?x � ��#B5� �@��,�@Ўo\9[齠��*hC+��)�
� ��7��;9�p޷���	a�
��
�d�4�+P��aMU#BUP
F�:�"�U A����]���� 8W���!�G੿��>hh;�)��B$`��
�@g{g���,�ꣁ����:�AUY��$(o-G3�Znm�8j�J��"�/dg�T�0k3�|$��ڷ��nq���\v;�L�N�j��ĳ7h��If�dn�vx�]s���'h{jl=;��9ǆ:�5����T�X�,�����H�!F���-/�\ۭ'78<r� �r�r��Z7W+۬Mb`%e����&+-�+-�	xF[�ܺ�n#a��{�����0�����C:��q)���a@ه�ē)�:��@xhC��KB��%�0�����s��u�t�y�
�[������.�!�!4*�)�UP��L bJ�KB7���:��n�x�!LZ�ћ�	�v��g���t޷�f�BXhPe�PT�3��'y��#@sP�9���2���UJH��[�]C���)�M� 2���q �hC�� ���4U@�Uw�j��f�����0��"F���%�T�����:��u���І0+0
F�21���u��F� KB®�)�P�UB �U(��f3��99͂(h� *�{��e��k|@V! KW�KB��>��� �f��}SSC��FѺ��"���z�U Q���FC#I3�K��A���@)hC;��P�����l���Mc{��u���)��{n���,�!��P�0CMP�*�24%G��|<>�_;ӕ�6f ���*n��yu�Ej��w����rF��T���WF�sx�ƴ�.nO�HB�<<4/�$�q� ���}��^GuӨ�F�1�Y�RІjT��Y�橚B,az�����h3P
ZUD�4��� &������g5��V�=��[��ք1���u�HЪ�	���P4#7�DF��D�w�ƶfq��B!�v�	U����5�������BA�@)hFw}���`q�"�
�`���B ���B����PT��i��������:ί��뮢�Ө�F�6s �hC5D4*�Z�P������Yi֗2�74&$�t�U`b䄸����Wr��I5��7 �4#uD�TДP���;�j��o���ͼ;��l@N�����%)�44T�`�������f�޾!hS�Z�r�'yW}����{��Ѡ�! I۔"X*h+�_7�!�� $h��!�6�UH"ZT!}@���~�^�U~���P+�2(�V	YfĹ5I+��I�OwQ���ëh�Ϊ�W�o�-�����W�}
3�W;�׏@f�Z�q�u�_zu���`g0�$�
�BX
�@K ��_g73Ȥ��І��B%0Zh!�UP3�V���b�Z�P� 	h]hD�۬cyn�� [Ba� *�04!�
�-eBB�� �r�B�����dQ����[�Q�4����]����� ���� b��_�q2,]"��H]�y�LX�&l��7,D�ˢ�j)�䓮�<����'����#u �hUP�c
h�k{�q��T_zu���hG9ݚ�-ð7���>�
� KB
�@K ��@�UB ��S�p�s��!,4�3� ���]�;�Ư�o�
�SB
�:�@Pw4�x�#Cb�jSBBB��$hCL*��u�W3;�A�����������]��hGn4hT 
���;�o;�M
Ƅ5�H"Z�JF�}����U��_zu���B`g0
Z�w}#���9�C�r߁
�"B�]]�S?����٥Rh��Ȼ�8���#U���.�6��ju��b'��g|��H?G���@��� $`��
�#BT�
h7���;�޳~6�g���u��k����[���Ж�@"F�U Jh4��K���"a�E��<#�Һ2��3@�ì�� �ђ�70�]N�$}9'?Y'��%�
� ��6P���]�dt�wN7��oPhE�;}�3�0�7u(D�.H�+� ��pІ0.�
Z�c[|�1��lƅ��І0��<���g��f�ӨTF���)��p�Gj:�A:@��@S � $hCh5�#B.� ]��
� 9}�k��c����s�n���/�401�B�І^�)�]�4!����w#B1��u��@+M��#B� 	hCaw	]�]��r_;������﾿�F�w�@��hkn�A��~e׵����A�ͯL��eOxL���6���h��w����-�^�x���4�hNJ���a������R�����5��FN�<L���(l�s&d����+���Mfc��
*�@�w���n�	ҫ�Y���
�WU�8�>�#)<L��
W�e��3�If7j#MBOu��4�;��%uޑ0�,��Tӳӻz]H���AGxʫ�W]�{�!�G�ѥv��}��j�|����t�]:V�eWW^m��t�H�fgajT�l�WT����[�r;�]�\�;2��pVR+[���6.���R�u\�*)Ҿ����9X#��8A��r�7�(,�n�J@؁:�m�]]5K�Z"����r?ٔf٪��bN�/��j����ɴ�2oe��
	���&�T3�AWۙ����@�NH����{�卮�Y���5%��[ڠ�t�ڽ���ʗ��Xw��Pff��X�!Sz�TGQ�C{.�P��䶗���+mؤAu�s.�a����q(c�R�#KŞ"�Nu�֕�o� �{G ��e��Gof�_e�177�Z)
|�)�T�'{n���7���\��ӵW7���G�olnٛ�nl@Yj���1qU�� G�Ċ$�I�
��Imݢ��~&�m�)ļ��������m��G :s�yk۴��ID$�<{�wۈp�	�Fۜt���;�V�J���:{�HW���z�y�ם��%�9��,�tT�u@Y��n�qՠBYg^v����Ѷt,ŝa9�sns����k8�wyݧy�on𽛎(S�0��H�%�G;�;:PC���e���u�	yvqYV�E"A�Ol%�ݦ�[gI		�;��Nζݗ�qt��n]�r��C�%�im�������W�ҮC��z�6çKKoWnT�����x/��k�������8D�v��p�gp&8����;T�#-f!�Yf֚	+/m�j�
+ˣc��:�m�$��z���M38�vݖ�����s��^��qӕ'e��E˫�n���(6�:�w�qס�ݎța�� �k���^3��Ӽ#s�Oi�N@3B���#t�ұu�k�E�R.,x�L:]x]L��lWmq��pG�1m������VX*��B�u����vOY&�Vz��o�����tV��d��n	@.F�jG�N.=��݌�eN�M��4	����E�"����vF�v���0�5���fҘx)����f�و<<Kb��*�?:��VC�৴nۮ�#N�d���H1�9�dwqs�.�K� ��c7M.,���x%� ��5:�lKѰ�n]�8���zb�M��i+���Ӯۄ�ɞV��B��Vq��n�ץm۷����5��̞+v����: +���f�Y�V�3Y9�]��{u]��lEV�,�׵^�N�VӢ���iu�����x^azN�\���Ks�r�;���$����`M1Ƶ�:�,�;<�X�y�8Q�9ط*q�Fu�n�C:
ل-i�d"����܈�p�k�>|���-��'c*�����	��+⻞�8�ζ#�Le%,9���4Xb]��UϤ��n��6Rm1Ivit�<t�g�ߏ��NI:�Z^��)J��HŰ��8tY�tz䫇3���8��%�s0c.,�K���q���k�<ѹgWh�f�M����v��/��x�������ɕ����fYc���]Af�Kf]�6җ*:�Cjzݲ� J��Y�����C!�����������(��.cS�u�s�5�djs^���[NP`g@����{�>�\'�����];�U���m�ͯ�kB�g���h����Q����ْ`�Q��˜�m��_i�qu<˞�*{�g��Cۑ�2=�h>��ױ�i׳!�v���ewN�^�C�|��������h�m���Er�kGI]���� r���G���^��Y]h�ҩH̛\�M�Wv�َx9���І��Q�Q�29*n떛�|6��u���E�{����i��Q�$�^��}�\��].��#)��vo���Ff,]��r�\��[s�a\�P�_��| ޕ�;c�������;n-�og�`Q�o���(-�և��n�m�I�/�߻��rWi��p��3330c��Z0$&!5��v_�9��	���������M��0�It��Ns��1gt��|�6�~���zW������6�\R.&�����nf�.�ؘBj;k�����zw�;�o}�s�8m6��CUˋ�(���̀3#�":F�w_r0�X}Z�w\��.�3�Б��q��?L�41�����������"�:剣��eۈ�Z!Xk�$��R[w}�yU�q)m��Wl���B��i,��B�u�������<#i����V�z���c��+ٙ�Ss�������K��f@u�w�;���6��:��=�����U�i��k��W�eV���OT�K��݇;��� �H�m���Qyߓ�Lb�krμV:%������p�x.* մ��N����̀3#g����N����7�T�s����@6�h78�k�u����T�u�Ou��M_{�8�o!MV]�T�-��͠����}~�}2���:��-	m�k�Uv�3/ �C��qw�wo���Ҽ+P��}u����^�yfv7HW^�hY�����w1Q̓���ogK����`+�+�nkfbB�B�Cp�u³7y�x#^3}A��aU@UUce�o*��ߏ5]i��uG��2<3��;������$:�\m=���ƛ�]��"XSnSfh��������B{oݗ�|�OA��
���؜�{2d{2^�$���+���Ԥ���|+Pɶ6Y����|�o&۰�6�w\�vw�������>���3"�CWF�����ݠ3)�u�[vN��M���2H�m6����Y��-�ؓ|iSz��{Ӱ�e�X$�6e�<�{KX��u�s��${{��cݗN���:_D��<��t������[�k�m����$��$�҇�l�����%�4G]b�yh]��Xh���l��*:C�ٸ-���^����i�:�]\�8�H���֠��-f WB�m+s@��Q��-��6v�G;J�V&M.��fa��Ƭ�ח�b�m�a�d2����r<u�m��#n�4x��G{�����F�肻p�ᳶ�Ϯ�D��q5j�&�Y]_�����ƾm��~s�يf�羙o�>Z����' �m|�
Q��P�u��5�iW;�U��d��n�e�L*�L:n����10DB�ص�t�7���N�^���A�vwHFJ����fFR[�ˏ]F�j�u@�ܹoBT�y�V��7a� m6�Ex�7�m�s����/v�V�ܞk�͡�u�֮�s~���:�gme�\.c��K	r�����ͤ4��:u��cأّ���\�O�e7���Ux�[�y��m��^.yO�f�n�����{YTʬ��z�j�c���u�U�Ώc��[1�f4M�˲m��k/+|$	 �}}`b�ݾL�u[M�s��d�l��꺭=UI���۶�
}F�՞�����fl�hHݶ�L4oln�:[�e�kyAJ�|�)�o'�;�U*�iz�R��v_6���U۾�n	�o����>�������3#1FHux����Њ��+��"8{*�<��|��WB�5aj��"�恚��m �j���9�]v���{�易r���^́k���҅t�ћ�O.M>S�޷��*/��M��pfN�߉�-	��۬ͺl�
��bT��L���F�ח�;��o��^-�o*z���.�ZյU���e,�j��{����z��[W��Tx>������| �;�o���_@̍�\���J��Wz��e���W��m ����+o�P]�^}�ޕ/�w:���M��h�S���������qu9s����Z7P�-fySB*��~�����d{3-�z�UT�j�K��m5��}U�����dN����7ا����W]����6�h�=�~�N/���m�e�=�N�!K=ޜ�K�νQ}�n�m7N���J�[���ǋkZg�ju��=���ۿ`�9آo�������G&�mE�+��
(�~�d�Dl�Y�j�S��n�8�,�8�u$��j��Ȫ��i��+��ٳ���,}}���ݞ̓�1|�m�gY��`ŋ���Qf�����W�;[c;�m	q]V��J�𘆶�7<���_������k�5Tl��̡��ew%õ5����F���W[��¼��7�[��%��▀ȃh6�~F��H�7q�g�9����=�b8�i��ho_{D�}�L�P3!)M7}�i�o'�;�H#dM�I�Cx�m�������%��#�r�u�ޞ��M��	��}��Z�w���'�
a��VR�=0��`�m�"k;e����E��J��U�P�^�1�,@f��dH�$�99'߼�$ʙ��FQ��jZ9���\a�M]���vm��8��˞���8��#��lɓe��G�b�i]L\ą�xInP���}�������cLr v�4j<�R�Q �3�1�B�-�06�ƱOTv=r�۱�ckфn�c��p<�6+�ᐮ�輪���ܹ�i��q6��F�c�t�c�P��v��$�U��: 3Pm ��s=O}7}�'�-~{�;Χ|�m�m?e��q����\��c]�o'�' љ�z6uEIP6�k�����jj[������]��f�M������h6��*��=�՛�^{z����v��x^!}y��%����͠�`�������'gN�^��6�u�:��9�vW ������$��c�S"4+��L^!AΖ�ez�����hI��������s����#����(�����6��T��Nޚl�lL��*8��3aOwL�&EE�oU&��`آ�%�.R���܅�߇�� }��O�앿n����Uǆ��g�;�x��3�|���m�Tќ�#�p��7�x
k܃k��ͭ�VJ>��]/������Ou��\���ۡ;�L���}�����F稽y�U'u9���=��=����ib�n�B�����l�U]�k�:�5���=�m3:���`#H��Wh����'��hv�Ow_�'s�ν�=��y�A���S�*n�p��n��ֽWê��m�7`և�1�k�����Ǻ��S�ny�1֙���n᜖w5vmc�Уn�4%{L+�ys��JI:OLn)h^��˻�i��b��^�e�3����ˤ�$c¶jE=4eI˽�sKn��u��ɂ��&*��6oqsY�	�����aZ�.Ι���L��홪��Kk��T�6�ږ��;s1cXwt)s-]R�7uj�w�;#�l�d9���:p��ȎBr��v�)Z�����w�$m;��Zuu'xXa�,�T��+Uv_�B+y���:%k���b�T�W,Ȃ[�h:�S�b�J���w�.��������s*�p<V���Mq�*��%�z����f7A�+g*S���:�j��ݻu���z]�<_IY�[lL�5�<z�E6���
�y5���UN��Y�Й����2&)��J�ћ�M͚.���v,�����^Vn5E�!��p`��#��kN�n"��̾���SkY�j���`��͒�rq��;��͐�����xU5�)Oہ�xIYy� ����o77�M4ٗ��;��E�2��K��=QUG�*:ª�oj�
�Vvv���2d�Tv��8�>�.��gv:�ݮ㝛j�[�ykj��-df�q7Z��j���1p6&��8�CJM������:Ƴ*ٿݱ٬��r�
-����ŷjӲ9��;kt��"�oz�{V[�mh�;�"8�{����tq�p���NN�/kgdPq��=�$�͙D���m�%	���jQ�$��w6�N^��[d"N�:;���9"N��;s�lJyŻn��{Z��d���#����8���kϵ����$���&ێ(8'".���8�`}�|�D��Z �NO��bm������-w��ƫw[�5�n���M�@6�k��Od���7��|��:��y<=7\��d�(���H��^��m �l�;:�;��Z�;=f�t��w��n��b��[�a�mY�v:�QI�H��u�He�kD�H�"��W��r؃i��So��^K��'��1����u������Sŭ	q�M��P�l7���znG�$��QPmS�6݀�����ة+����ʉ�z���>�fff`'������_ͩ.�w=ȼ�������[]�~�)��̫�P�'*5tc��aq��v�LLdø��d;x���u0/�x{��.���6�A����mfL����v��+�V-�v��=�.yG��n͛mJ�]s��#��t�����H�	�UF�UN������ُ���\鹾>̞8�������u��h�|���P{U�lv.����g.~���|M�\���h6�o��ChK�U���x{��]��J�Ջ��w�k�����y�i�b��׻�N���\��^T�5ԫ*�;|�_�n�����b�յ�2s��پ�~؃h��<ۦN]G��.�J��������<*;Ug$���!�:w��2�$�uL���9afN�Wu�o2"��&���t��>�l�=m�Xls�=�Z�vRuʲ���+��u#��
&���w5nu��s٫7R�@Q�SV� �C��1�Ѹ��\����Cvv�K�|�,^��9:�z,m�xw>?>	󝑪w�{Bj�^O\�z��-SX�]fv8]��}��l�f)���\]�H�SW��?N}�'���d�v�o���Og���&�{�c��mԧNܚ��l��ُ�󺫝����G�!���MH���t�P333�/�W����oFgG��:��\��3*�]a]��fG��S}�Vb{<&׫�}�Xw�>�����m|o��QF�r����󻫝7<y�A����<�u���M�B�l�i`;�k�ˣ�i��j�Z,�pr�����ᜃi�*���7잮���>��m�֣M��o@ɶ�#c:���DGo���&���޴ɬ�'f��Bet�8#4�Ǯi4�`f�[�����~�U�_k�r����ށ��U���M@6݆�0����Fk��wus��y�M��k�M�4�!�7�v�f���~��N��Q|P�-�Vd��<[ΗG.�T���7�3 fV�U�^�S�=�'�!l�?[s٥Y]\�H�B`5vV�m�aNߤ������%�蓽�j�t��~������}]�hw����v:y=���u�P���6��9�J�-̘�N7���ǟ/�i����+<s�i�)�o+�Q	n73��܅��6��|��J���a���������{��]�����L�+��6�m����{u�O��;ɵ/עO{�������gP�f���a��o�s#R���/h��4K�	��
�5�a�V��u%�Q��U
�**�b�:sql�B[v�5|���Q�j��������׾[��U+��Rq�`�Z���33(f@� �J��E���'w�����}^@w�}X��x����m6�a��&{���1�4T���+W�۶�m�Ӝ1dV��3 e�}	w5R���W�ҬQ�M�w�\&(����;�ԏ{2Wl��u(��f�w�I�YVb�*�;� >�������٧ߥ�r#����w�U����^_w���bR�y�n�B�݋θ0쥵�qN������P������W��f������{4T�	�~�ޤ�e�� �w�m%����������\��Ik��]��Sw����CZm��6{+���T3���ĝ��.�������n�G���T�>v�����ogQ��=��i��:�s������OY����ڷ��+wg8�w�@6|�3J��z�Q���kzL�n�����`m+ʋ2��V�7��0숙WV1�e�	�� ����W�([��zQ5�u�<����ҹ1�@γ&���5�����%���b�ui.��xf�8-n֢R�G7�.��d�ˢ�2a"�At����]2%��8�r�V�{�؋�͆w�<�b����1�v�� zY�=S�3��а��}~����v/4Yә��ݶ�ln*,*r��Lb�\���}��g;���m�����My��}*�Xm|mW��񣰳��q�Nԙ�w���܁����^J-G�#ّ�7�5c�\�:�}�qo[�9�}V��|���s�֓>~*�����׫�묚oVw�T�P7|�4�3W>�k��m|�K�1^�W�M�Q�������M�?�զ\wOi�>��ٶ؉2i���2��3v�5��8���8���ߎ{�}��Ӆσ�k^oD�ct�*�NGlfc����f���1�ǥ�b����EM��FƓ��U��Gvѫ�Y������-n^\��"�����=��: �Vls��&�՜:�јs�i?t�r��m��S�pu��d]㞯#��}Q�h6�Ca�v�[��^!m}�Y�W>5�y��ʬ���u��3#ّ�̭��V��BK�6뼛oS����M��bڻ�6��zUe|�R!Uۨ.-mٻQ۵ͮ�8TBUU�/����Zs������/pͯ��^3��^���m����=ҩU�i�%>���������чѿ-����h�hc��(M�wz����-�f��g;���^�^����+��{��.�=Pb�h�Q�k$Gխ�8,�ˢ�xx��뼜oV}=̌�Y�3�n��K��2!%e�nxB���v��])��2 �m|����g�]~p�b�ul��)ik��5�2d�*zf����	b��Uq3,֭�ـ� ��S�l`M��u?>g@ř^̆�V�/���W��1z�jEZ4m��g�y��[`dK޽����n�{��s���d��՜�A�x��I��+=]=����W;���m��)�]���z�{1;՝���1��}�="���l��gU��w���k�4�[Y����R���Z]"7grCN�wS֨m-Fb�t�Cyh��X�9T/����ùڛM��g��Um���/�pHmo���ܯ6�@7�/i�P�
V(�S�u�D��Ml���x��n����UR7}{��:/�A�t������ ���T�����m6�yi���#iY�P7�;��w\��֕xW��7,9��Ы�o��ƃm��ð>%�!j��]�vw��~&�m��O*&^�/6�m:��^��y�oIޜ��3�n�R��2�fe��u����w�S�K5�|�xr̬��E��1j�f���*�EM3��h�3^�N�)\�����N����dK3��v�owik��{�Y�p\��uf�%Mk:�� ޟm�ዧm�hfƙ�b.����T���lҽ�l�pV�8�%k�E7H�̺����5�1We���6��VwwI�7'\�]7�S���.Y�J��(d�ʜ~w1���L�^�K��U�\�fǳr��W�g�153t�I�����n�ݩ�'F݉��Sȁu{��^홚L˕qDB��M�oD͓7�F=[kd��O�A��so;,�Yv��s�9{����ش������E"=�^.�[�%����7Qj��6ճ,�H �(T�ʆ��d:�^B(z�#y��{tn3u��Z�#yR��)o����������6%s�C]̩J�Wo)��{;�-�7Ume�gkr�1�Ƨ
ݪ̭4�*L��6UK7x��;3�Z�YF�s�q+��9[9��s\q_�9�Q3��Pڜ�����S)�Q�ȭ��uD�#���v�U1�7zJ�[�V�D��]P�Ë~�uoFU���mW-�Ү����������v��3�l#���ܧv3��u~Gۜ�m��� ���;;ο���.N����=�;q�t��bq�o6�kw�׷_7�xv�٭n$�K�lw��z��aXo���%,漩%2�yL�8X���gm���,����������^{k;��);�6����	+m��y�v�k�%���$��
6L���Չ��̅ [yϷ�k��G_mw�D_of�bG�I�!����c��c����xg�[ؕ�����B+m�rt�p\{ڲ�+��99�6�m��&�ȒJ_+��-���i_l��6��Z3>۲�ۓ7fok�y�y�q�io;��=�-4e.ɦ��[f�ҹ�����f�0X�D%q��iLm�1���c�>ő��%�-�*5�r����\n�	����v��!�Y�p5��8����|�E�j��ƅ�{���n�G�b��&�L+I- �Gb�;':��x��9tԣʵQyT�
���ر��av�q�v.�4�n1������o�m�q�{A�p6{E�Ttle�������M:��5�]y��7֍6֤1تy���d���3��n��G�\�ʷX��㲨q�b�E}�:zI�U��\\
���a�=�y[��X�DR<���@��f�x�4���ع���jWi�&!�L�b�,-]���<�h�wX:�%���-n��c����:^�hf�5� l�vln5��tI�2M�0��`l�u�mn���ʡ�9���)3m���l���)�Sk�������X���0K�����u��1�xr�Y.Wv-(��H6N{q.�`��^��#ݛ��q0c���j���-�(�th��&�A�[��w4�ۧ�N㰘��@f-������"h��k�W W0�9�SX�9�N4����=�2�R�$47'i��UF��G=��×�nyosrY�\�=<�z���tQ����0v=)���vk\����w9�Mu�W<�,��2�Hٵ҃�m�Fm���n(=�0�]�q����!�)sv�;���v��5O:��\/j�bz���i{1��΃����؛!F�j�ZrNN�u��R��ڳ4^�ڸI�î����v��0Ji43�Kv���U��^��;�g�8/=�q�m��܁�����N��9q6N9�7��<�kb���k��I�7U�u���vn���\fY6�qӟ!�����������щ��ۈ��X��c�]U���������/U�gfۉ�/6{dpԻ���&d�1T�O[���������o%�;��T.����=��d��:��Z5@Y=����ym=Μ��1G�\<ڮC�i�@�����`T���N���i_xOr���dfG���YQ6�Ԯ�3#� ���.K����Skj�|7s�6�i���ɝ�p�ԅz��/}�<﷛𦧓h7<BZK�h�t{7Yӹ�bǰ�Qq̪$�h���F�Uv�؇4@7:5ٯ�Ԭ֕�Y�a�U��;��y����09�zd�>��v�C�uU)�@��8��V��̗u�F�I)���G��)�D�+'f�gs�R�+��{���
��S��a�	r\2�fG�!¾�[5�,�UC�e����C�.�|�o����o��ɶ�؈���<�*~C��c[��2�ZWê2"JP��87� 9�`6�h6��x�1�P4�����28%ڸe@���nZ���4Mo��vq�=�u�i�a�)ll���L�\���Nu��_6�󽏯ݾ�w[���^���Dx���k��曧g���_�t~����֕p��3z+���*{��>��D0~2+)�]��^P���}�����v��zyͻn�i�QL�\i���/��_m�%����w�>��sI�v������(~���}"�*�p���sm���}�V�Ŵ�sK'r��~���V�Bv/V��	��|D�P2!DH��34�
h��.�m��c�B����A�R$�ٟ�"�o�������)H�m�kce5!���LjX��I����*<�j=#� �Ă;�
e {�G"���3��ܮ:\A�"K��dI!FED;�-m�>!��j����5��d7A��;��mu4yV���?P���
��$@���س^���f'�)��D���H#v=>ݑ'v$�ZCy٢�=}���`�݉���dr+�O�r�O�g����X�U3@��WNr�B���邪f{�.ګ�H��32�d9�/f܈�*p�*�R�b�X���+�U��7�$eܒ��F]�$n�]?C���T@Λ���z�u���xk��0ȨL�L�Y�,НI��c�*�-J2��	-+��V�uh�ml�ڜ�'��H�,�כ����r����OHS�D�8w����C�_H��dTE�Fe���:�� �q"]+B�Es	��^ +�(P2 �2��y}��'�P>/�H;�$�ٟ�r��s���U�m����U���m}_OW�,d_I��:(��V�#5
3U"<����{���S�tI�c�ށ����H;� ���2P�"�>`�����Ԫ��h^c!����A.�����YvFz�H���5�1	p���I{;��`R�C��uL\��q�{&OVv�Y}���>��i�l�I�;��a���-��W6²mZ�y�NIs&�Y�vo#Y��Ҵ���ٜ��sCy��E�M�+AY����ND�^��heҗH�hl���5\�ڶ��nÓ�xMq�܉�^��]҃�e�ݍf޳z���p	ҕ��+,�z�m�ܴܡf��M�����F��z�#N��d�l����h���0b�����_Ǟ|q�z�Y�y|����[ظf�q���)�1����@�W���QP�~2!Do�.����\H �>Q�k��g2���tO��D���Ѩp��[T~�}BJ�E�A���;���1t=�oW���L��SU$��As�Q�rf���^��;���
����ٞ{��r�^m���Ր.m���L2�P �j�D0����}0���5�ˋ�gr�����$[� �3��W�߻��'�u{��Y�ᴭ	�u�M^9�S\�$�+MS5���qD�9G�`�ު��|68.�7���a��j�����	(Q!Gv<�4i��9T�"�3T��}"\�]H)&���W]m�6��f�<��Wu�yk���FGe�����?���H����o׋V�ظf�q�Ց$s��}��W�����j��������FED({uP6���l���= ����"A�����糖졳�ִ|�Q���d�uT�=�����H ���A��n��/w�6��B��
2*(Q&;Թͽ�=R'u�n�<[�����q��j��Ȩ���u���DUR��B�]��6#n�L!Q�Sn,�n����d}��e��O�9�<�x�cV�>mFRzB�"�b��1�����$�ĐN�O�}W�S=}�0{c�WD�U$�w��a>��	n�����;���%̉"��'�=;�$���Po�,w��]��̔�WV���V;���������]ۄ'c�����%e��gn�J�P���l�N�| �=7'y���r��|A6��&РdT Ȩ�(W�X�WW��C�z!G�Q!AD��ϗ#t��S�5�$]�P�ù�NC��U����"����!FDT��h��:���ЧU�Ǫ��+�"���8����v�3,b�Q��M����*�ҵ�7*6aY\d]���^_;g������Z����3���/�X貣�&\ A�P��T~�}&P ȅ3cy�u\��H8�H!�J[�r7m�= �~TAޡ@���.Yy�����3<�A�/�C���ȷ��yK%�l����ݕ{�û�Wو
}B����&Pɽ$��(��D��Hݑ#�d�K�s�cQY�k"A:�%.,���f��]b��n�kiN�]��\El��,VX8'��A�&B���3ՑY7W���S	y)7V�{���n6u�p�deܩWpK.�]��dY��>1���;��>\��{O	��T;���P�k-�״b^�*$��`b�]s�h�ݯ5�=T�5r�w�l��N~�_<	݅3:�}ئ��	��l����cyھ���P�D�@�.*�u�X(�R'ڠOr�Z�eoƢ�=��D��FE�Ȥ�E�G�Q�(����;��ݑ=\jB1��orh�ǲ���<�"J�����aV�^�������@A��'���U�݊k�0�	�AKkdP�WW}"�D4"dT!@#6J�}X{�6㭝��<�W�
���׈?^���H��WbGy�F}Fgrh�ݢn亝X��T�Ų�g2��K���S���>{{���W���8 �t�qv�!ȇ����X�cV�ss�$�:1=q4-8�u����K ��V:��Z��D��& �;3�B��\[��k����k4�$Tԡ�:�]XOm��:��{;ٜ�g���˶�-vd�t��< dy���y7:v����������������e���gb⬣�#��]GY�[˛u��S��$c� �ĐwdOB�R�����Rp�r�:�a5q��۟���_� ��������%��p>]
fPA�b���7�O�`I�����8�V/=�.E�B����(QU|d��o�Iet�'���m}�mQv��"�IT;Vx:YSnn}�,�@P��r�m�*��}~TCI�s���/��=(Q�Q�ED%
E`���G�P>򫻿݋��0�O�@�A�'�v=;�7�����������IJ�WM)u!��;�(\�Xk����*)6�}�A;��P,�ٟ�"@\�֣�s�SJ����XA�B���%}@�$	"�3�
�F)b��+~�t��fh�򬹪��ԝvJړT��I����wQ���P�&���*��t�)�~  ����O�R'�U���\��͐���p���O�ʡGq}_��� �"ܩw�W�˼������ޡ@��(Ⱦ�(	h���Kd��������r��nѶ�&���q �-��0�TA;ʁU}"��_Z
1��,�ej�������t�tI�Ȓ7f|wdOF���~�ݕ���\kJК��1t�#�T`ݕ-��k2ޟr�(��I݉ؗUZ�C�]8����pW���4� ��Q�P �(I�>ݏR�o6��F
��>)ȕ�-A=��W=6׾ �mQ���u&}�ݫ�T�g9Q�@�5RP�dTAW��P���=Xz�3wv�����|y��$�3c��l��2�qB�X&kv!s(�nl���Z���$���u7���T��yR�e�\�ɔz'��Ŝ{���z�0��V���q��y����:�u����R�=H��<e�y�f�;����C�h�q�j��sS9��A���é��f��3�<��9���f�κ�dd�;r6*ܝ"7'1�*4x��dbu�]\'�Q�v�-�᷹��;�U�*��N�RM�߭�ʖ�J���[5��z�	�8̮;8X�8]�����;��Ė����������S:�N5E������xJ��Y�﹍[�h)+w�LAX���q�]�:c�{)��q7�n��vRSɓ9ooATj|j��X�� �D����V/��Cj���ޝ�k�+p'V!�3������#Pn�f�Χ'j�2uu�F�-�X.��֋���b�^劒B�Y��Y4�����u�ws�Uf.�s֞VTN�ֹ� �H�m�v�T�5����V1T�KMbĮF��Ԯ�&|gmGw1����[ֶF^�[�wl��B�t�
�n�z���k�a��4�HU9T����M����O׻�T���ڃ���csZŜ��u��kQ�ۼ���յ��=�}���Si�C�i)sW���G����5���������[�ff�.��ye��.C�\'�L���{m�u�����}`_jn�h�E�{^ɳ²ʜ�T��BP� r��彾����׸^��;/ ��K-���!9XQal%�Y�=緂W��޽y�٥�ɷ[���2p����8#af��if1L��}����n��ٚOm������v�f{�g�c��6-NB��n�5�,:��8%O>ʦ8�Ov;w��9@�*a��!!-H���%�{V�N>�����^���b�c�0Z^[5h-X���Z
�(ZK��x
���Yr�W��)T�������; �:��m�o��q��	L�߈ߍ��McuW&��F<r%���D�+�%
2/�����j�A͡E�	݉uU��K�a�(�&����w�
���"��.P#����w@��]�^<b��A5�$��b�AE��k�V��.�]�U�Wen�l�<op����H�!g����ja�>x�/_���|�l�vD�
��\%<͐�����{J�kRVA�@9��"J�}_�y\�®$�uC��@�vs�x�} ���'��"�����hi#܅��	(P"J���=��.�t�n�>~����A����B�2* � D�Q�7��8>N}���"z)ao��J{{!G	�tH!r�޷w3�`�%d�!;ŵ��^�^��6���xR��KS�R>�P��<�߃o�w{��^x%s#ݟ��p��|ܒ;����]�����'�e�Hʪz6��w�7ޟ;�$oH��2Pڔ�p�(���!HP�����ۮz�s/V�+�u�-ɢ�*�n��O��A��
IB�?IB��f����.�^/*�5皾��(� $X��d@d��^��Z�U���ޑ (���ot���B�����"H��߽����(P7|A��ʈ2W�, ��7k8e��[7�7�����ȨD�(�*�Yf�T"4(�B�2P����������j�j��p3ܨ���$�Ȁ�+��ۺ��A�"�k)v���Q�	��HJ@�|D�3}�ST.��w��ڕV[�Q��F�^ޢi���gU�FL���Du\�zw$m);z�ȩ2�|=�?�}�l�u�j���tb�4����<��u�̹�36���ŏQ]�RB��p۵�Gv��U�E7M͈�U���qM˻6�����^I�HՄ(+4-X2������:��vh2��j��ۇ��j�|g���^���8 ��[/�q��nk���ߩ�����k.����.-�M`Tڅ����q�%���?/�@H���t��98w{�t֟v��!�^У���%&
Ȩ����!�;�8�ϻ`>*�����s��G��۱1�����9�8���IB���J]^"�=��6w�wL�5xP ߕ|Aݠ$���(Q�P!�o�h�R�Z�B�j���E[wst�s�e[��m��Gd(�/p��ꯈ#��$��dTD�	��fc��'t+Y�vv˝F�=Ʈ'����;|A2!X�|&���4+(j��U
Ɠ<�d`=f�6��`�`աwhvWޤ<_ ��Ȩ"�D�<�_L7[�t�هܶ�D\yTo��$�FD�
�I��I��Wu0�/;���w�jI��Z�h����rn�{&@�����@�3.�!c�"3v�����ڑ�J$��$:�IFJ���L5��p(��B��J<pP��Т5��;� nǷ`JZ�{��ip��s��GM��}"E����[�G��[�gE�wdHq+>���� ��Fg8Z�h���Q�}@Ⱦ�(Q�.��7�s�M���\1���m��e��Ǘ��<']w}���Ҍ7 7]iݣ)1ذ��Լ��5�E&�ϻ�2����yg�<��B��&�{��_T�mx��t-��R�g!@�* �$�ȅ=���e8#.�I�!�0���e��AW	��� n��wo�=��'g���v=���I��5ˣ��������S~��iȵy5�[WJ(N�`�2hK����4��e��	�C�^A�5Rk���=��|_^���7��, �@I�@Kf,ѳAJD���|}�"[�;���s��G�=�V�[���q�͍ �{U%
�D(d�_I���	��d#z9����
�A�=)H�$�_(a����3�dUX�TmY8M�Z��F�t��xh]�u
�R7I]^/��TAk��T:�f��s���O
+�V!�A�����2P�D�_H��=T}�����P}'[�Byc�F�8�j�A%"N�m�w�X^l#Ԩ��P3����Fl����3	t.J���*���D��HQ/�C�QUDS��,2/������J�kn�pP��zA6�HO��;����]�$�J^]�.h��2j���**&�YpdLUcJ�5�ok�`��n;�(��6��s#�{�|A9v�wbH݀7w��t��t����Az{�i���^#u
E�"�o3���}?w��KcPn'�Cr���.�V)�5��̣S���A�����Q+>es���*�~��[j A�(����/��}����{�=U�/�y]�X��{��/:A�	�Iݍ�\�fg�� �R���d Ct+��t=e�=���.I:��c�q}�x�wk�|AE�Vgm���`�P$��N�Q+>e.w��*�S�uvN*j"��=!���YȨ�%}"�^�ϼ��7}|kg���{�W~�Nr�_H��+�Ö����x޳j���=�=����ҿIov��*��]��I����]\41�,کGb�������,�g��9�Pg�53Fz�OX�6�W4s�%�����bb���ia��:7F�X�9�#$km��������nx�ٻuA�N�zt�ͧ�ȣ��O5�-簕 n�l�`\X��ܝ��Uzè.�X�ݬO�u�ݵC�s����n9<��t,��Õͦ�����#�����q��>�9��˽��e�	�Gi�D�r���;�FY�$���Nrv��3[CS�so&"�
���?H�%
�/E�j��U��@��V�����M�C�V���=#\��SMF��Dz�
D�wA�J("dTAֳ�2�&䷹'xj�����
2* �B�"J�����3=�1��$s�N��wQX���A9���O1� �ϯ	�%P&D(��d[.��$t�;�^І7��G6WiV%p�M�y8v=�Zӿ��E�`	i�mt�̺Y�i�K�W[��n�������H�"N�zN�HJ�ҬU����	R�fľ�Իut@`�ϹŐwd�	ݏ��-��b��\��R�Q��zjs�6��0-�-an1%!5�jPP-\�")�:ȿ;�Lp^H�'!��'����x�lq��O�)O�`�F�M�`�ܨ����(��,%=^�\��N��ޕ�#SҨ*�S�����'�EDW������P�}��?H��]ު�;�Ħ/ p4�	�s4��h<�܀�("�A��|D�̑u������H�Z统aX��� ��ǧ�Le�����v��������A�E�9�>P�Y�X�،�5�شݥ����C��E���*����#WiT@�6�Fmݬ�v�'"��
EG���� � �wUv�az�Oo��1�㸅�B����'���@�hWǹQ!DIU��J��!Bo�Ǘ�MYj�a�q��e�<B��Uvl"U���D+kn]l4kV-fR��UϦ��q���y��+y���M��}"������/�m���B�[N8��v�������+���$\��"���J�	"�Dr��Ɂ�;��E�ޣ8c�b�!FEDH��x�ܩ�r��I���W�<���c�G�lT��������I���?2�=e��ώ�r�{��o-���8�HS+UzP�9Qȫ�$�ȅپ&���v�b�qĂt�
6��]�5���Jx�D��H��s �XMx8��qd_/�IB���2&6U>~�K��w}Gxc��	�@V���`"D(��u�u�ۏPdHb�O���oWs�
�[5���q$0g�pp���Pl�6y�:��l��'xų�V6�{)����*��N��W��r݉�
7.$Λ�냮N��Q������D�P2.-#��5�e&�퉭\��P8�G�>�>#v=;�*��y}څ1*"H�Sk�i�9�
��Е;&p�Z�U��g|yy�e��X˻Av'ܮ��s�L^w�qn�Z�u��(Q訉�D�Q�Q
����݀��P#rg�)ʷ��k�o-����1P ���D
^K��D_W�	��"�}RP�;��c�g
���B����P ��
IU��'�ȸ��[�I݆�v��s�L^G�@���#.2H�P�֤.�#N�%1�rI�#H�ZR)�][ݮ���kc���H �"N�zN�h�Gj����핐�Jm��v5�Q�p�J�<��3���q|:��]����s�yބ� ǑW���۸ʶ�=�n�6	̛!�vѭ�&f"��R�M6�(9s)��;�uN[�ٷ2���ґL'��u���o�(��st��Ԝ2R����8���cZ�}�$�q�5Ύ757���W�oSh��1�7z[��Vpj	jGqX.�9G6d�c{f�N�ݛ�0�E�zm:����vrUe�+a�rɊ�sn���WϛW���E�e����䳒��"��~�K[���r��<މZk59����V�dmݼw�7�٩:�n��VSZ�ܚ�גĤ,��:M����X̣U�8*���k��T���>�N�m�-&�*�,��uI��s��FVƪ�
F�4�(��QB��gn�n!s��/*�ҧ���*5����<=u$���k��۾�yu��ͮ+kn�����=���;��]�cf�n�xz�e��5��vfL�uu��GT=�ˎm��d2i*�7ק����MVh��C��Z8���:5[��gWWv|�Vb�eG�+���Oe��ت�,Q=�,r֓�p���"P�P*����|��o���f���;-o{�����&ٱnK�_zľ�l�Eb�����ٝ���,���{m�[g��&a��ޞ�n[6��q�FV�VG�kP+-|ޚۯ��f��m3Q`��k/�Ӧس y��m���&d�����=�R�͋n��$�vv����m��!�H+e�qĒM�#K6Ӎ���ʹ�-f�����^��Ym�m�"Kv��6�w���ٳL�bD,0�{Y�[�f��g1�4γm��u����Nۭ�O/{q�D�!5�����m֖sk��z���NR̓k%�-�[��mii�5�]��%	��dl�s���kן�>fo{q/b%uH�c���F���9Y:܈�g���Ƿ:K�x�ӈ9�֠�^X���]��K�0A�4�3m��s�RP�J䴈��l�\n����x��ů9�L�-���a�^6wc�q���sl����^%I��$�A��b��ⓩ.�u�Ŝ�h�Sp�=�:ͮ�}��7����I��f�KTp�=v��8�1��Xr�r��6e�1ڐw<]md�R�ٹ"#���2rf�_Q�45����݋�;B`�۝;��!{mlx�+�m�B�dOOLg-9�c��.�5b��$!����Y�
���O'/n����XǨ3�����wZ�T�)�ZC�iLo麏S�v��8�ؼ�yܴ�r�ez��z�#�U��L;����K�䃍Ҹz�Qq���!�z�;����BT�I5����wݝ��ظw�k���Q85ݮ���{`	�j�yx�P��2�$KV8�`XK�`��F��BZt,5�t<k��Ih���n���1SMi�
%��E%��xn`��C8ף���cP8��V3	�ֶ�έd�JbLݭW]l�ȖIwHoh83���z6�˙��}�a�v��F�i��F6��8�	W��Ԗh[�g�ԜY�Y�����%�3Mv"qv��<�Ѷ�о�����r��D��.ˡ��G��r�=p��Q�v�F���yV�5<]a�^��h��{A�*mKSֺyݱ�E\��=#�7A����p�gvx��ƼR�=�o�o���m�\���/l�&��e��c���%��ƶ�6T�\\KM�瀂6�L1�%�5ІLRڔ�n�JMN�LcW�ۢ��f��#����6��_6ι�i�B$-�,�xd��q�#a������1�]�63s�rt���
�17U�GJ�W~�Aօ_P�dTA��R�w����ȥVVm��r���Q��"|FtzD0Ȁ�}~
K�wn:���ݺ�7��a1y�	� .�n�M��6#֨P#r��N�DH�%W�I@�'չ�ה�k�O-���]ĐBS�ز	݉#vD�|-�q�V�H9���`�7dq����	�\��] �]�q]m�`k���Jd_PE_4"_H��fua�Eb�[c_�q[��o��0Ȩ�%�Q�֞�U(%b���u��^V#����c<3���Uh݌�@��^�`�onyR��4��9��Sjz���P �'���$�A	ܱ�T|��Ī���&�+�^��d�0@���BV���̴�^���w�_9Qg\6j��k��s�G4p5� ����}V�֮FElz\}��l��	�b��P�|��{U D��#���]��V��gpp���>��> �W�/�B"~�����B�� O���Wʗw)�o͎ ���n�;'���J��q����@����
l �b�`gFS}�lMj�+zA�_W��E�IC��v�3'�՘�.��(�ąт�ؚiy��e5�k	��ƌ�iM�����l��y煟n��T��8�1��/8H��*���� ���"|F�{v,��!]SՄ�r'��H毒�|��<G6=�.$F�}"��f�_���Fm
ȅd��VA�샢JQ�n>�1M3;���7s(xMwU�w�����"�ފm�5{8k��/+z.�#u�q���N��V��Z�
ސMtz_H�7f|wdH2*���·�IZrՐ@�B���!�b�8����/;�	��!J�5��?Z�s��dTA�D�Q�}RP�$��VU	�R�!��5|�+R������
�Ⱦ�d]B��Ǹ���I ���ƗXM,�,f��2�l��f�X8����ם�F�>��Yf�q��筈���
ޟ;�-��G)�����v$�wb|D!oc�<�c�n$����8�N ��i��	�@S�
�Ȕoؒ5�~��(��A��%}_H�/�Գ'=���3٫���?[TF���?H��(W���y_@�>�;�U���6����i���U^�3�{/ks��1��}Ye \w3nn֗�Y6��+\�ܗK�;N�m����Æ���}_�(Ȩ�dT�}"k�cJ�]U���\3÷��P'؅�$@�vUA:����҄��5��\�K�������n]nFͽ�����_T�"�D=��{��s3���!������)S�7b�F�� ���'�v)���I�T��@���	]��D��	w'E���$Ȓ	ΏT�(Ⱦ�dL�;���[��c�V�3���7�(���
E@�%
"J���\X1=����={�'���|��x��{�lH#zE�VC�L?ȓ�����H�|dB�nuUV+��YB��橮`�6��z\q�#v}>;�:'���{^����lz�M��炌���j>���]���3
��</1���;z�e���H�k�g�m\��RF�@���7�c����]:,l�Ѻ��A%���79��]b�㷬zO8!�k&�������S���³x�B��t{96864MM]øw�;��`caC��>�o`1�m�;h8�kU�Nv�ܼ�u���AM���x_!��x6]�s�'�x��[NVX�W"T��k-	��݌�եu|������@Ȩ�dU�޽�+����m}�N��4���
����%&H �Ă�8)��@uG���%5}�����;����J$R�n�R��X�ŵ_܅�(���(�<n�����w��@�&��zA�$��@ݹ�P�d_w��M�z/��!�T�/[���S�>� =Pӵ�`g
8�Av�$B��Q!DI�J���^J�r)�v+h�Oݎ>�J�ؒ�xO:��y޳����+]�a�Z���z'v�x�њ�vm�V�E>�N�(��P2/�C���5ͩ��U�V%����	��}��` �ۥX��#k�H���f�-2e�a�k{z�뫳�E2��7��1DMl�&q�R�)�]�����d�ȯka�A�� ',՗����-�s�
#څ"���jN��]�j���쁻��!����v��V��1<FE�&�}��"�AE��]�}�*�{A{>ݑ �X�R�k�S!Lz\q�\��pQ�>)H���bH2W�*�ͱ��Ӿ��qo�<oP�XD�h�]Ӭۡ,�!L��	�Zݻn�7�̡H
�s��J^V&m����7�Ǟ�<��H��ٟnȕ���;�S�wc�z^�Tb���;�Q辠d_H����yc��}v(�r$�X���ͩ���;�Q-[�[���z���ܨ��"E�z��z������MC�3hT��h���g)�XOM�E�����%�S*\|�)���K��N���U6N&l&)���#��;�$�ݙ�d����7Hjg�۲$sV����nv���Q�5����1�b����U}"A���~̋i�N�h���b���HU���A~�$_H�~�5�rҞ�6��*�$�u���)�{A/8*�:Ѻ��U�hE�y|��?H��N�a���LS��Ϻb5ځ�!�sc۰,����Y<��o�]��>;-�WѮ�,k��� D-��n�����8�e� �$��AݟQOc]םhQ�if�u�Cqt�\$]��$�����v,�leS��Q���=����dwb}є��6{�e1O���#�T�9]��|�D:Wg8*CG��q�o�L�t[d5Ө���LiJ��N,4��0�[��:�W�Cf�=����D�@�$B�o�_WQ��zF�U��;J��68����}"�A2$��"��%aUa"iu��"KH%�`�(��+�"��2Tsy�}o�����xt>ݑ#�PŽe���:�ɑ����}�ʁ?P쯤B��P ����2����$ۏI��)-�;�ٴ����l!)�_x���
ȐBs>�U�JE�}%^��5�G$�y<��jz��7ջB��	%
b[ټS��`Y"Jq��:%Z��i��
ߗ�z�SE��r��` �"�7c۰�O�Ϻ�}�ՋX���m1K�n!D7k����#��h�g8�6�-��;(��ͽ�;�]�<�ۋ�]�A�>�̓c�����톄���CN�M�4�J]h����W�3��ps���bu�:ܕC�f��XE��o49(�2NS��r�����j;NP�:.:��Z$�=����h���;"���g�ks�x)��*��A��Fŵ�����j����jZ�f�Z�^�D��.#T$�F�4�t��.��~��.�7m�")�8`�M�T�՛�j�".����_{Pψ�}"�j�,������NX�����d_Q�}&P?"�y���ni��A{BP8�iٗ�S��A5���,������QO�$4j��=��`2*?H��#��W=u/g�{o:f���n!_whQ�QI@I���2/�ψ�}"���~��jz�A7���y,:8b�A3ʈ��}"A���:u�|+x�J�Bu�:���� |���s�!�MJ|��A�����Q�#{8ۇ���psTa�l2���-�3�<������<��3�K8W+��Lb�{V���B�"J�j���a�Q5,��s�W��'l����_	ά2�*��c5/*t,ٸ,I��#���V]e�5/LYf�M#ގ#\zF�|�9���_jz���F�dJ��_�뿥/�0P&rE����&���)�Y<}%��|+=sî�����GrE�O�����;g����P�{U@2*���g���ZcWzA�> ���0o�8��"H؅"���@�<���܎���W�׏�����D�}�qQv�"�	�r�������w�h��v��8qT�y�]�#ł��rX�,��Z�^@�C���z�ݐ�!���u�HwޟodD��s{��j���ݑ'b�� Ȩ�����DwV�/_��RΤƨk H ���MM	�vl++��#�B�3�ꒅ%W�IC ,����o�ky|6sh�lh��֣�c?�5]�d���#mTht��:�6M�՟������[Y��ӹS,�.��ͣ\n����[��z�A��r���)@��շlՋ3�R�D�}r��j����gl�Y��t���٭���xD��5S�ܦ�\A]gi�t����UMmRԫb.R��&��r�:�����5ɼr�X�S8�;�]�����c��Ϥ���ܵW��y�)mI��s��wi�u5]��&�׹Z��Gr�
Xח8=#&�����]�8�Oe]𮶺�7�W�*�v,�
th�,�ۖk��r��r�\�z��84�����"�Ӫ�ܽ�m]H;�2��F�pŷA�vaM�ND=��S�!S��+!qsB�UѺ;k�H)�2�i]�)M�)pkf�,bo�-DL\\:˓1S��,�Snqk뙩W�n-��yب�1uE;f�벆��w��aU�UN�*�c��M��ݏA����VF�C�iX����!I��V ��nS��)��,�y9��r�`���"��c��a�z�]cjFt�.9�ÝMV+gN�<�Q̛ �/1l�TseωH�A?/�_R�,�:4�n�m�m���[v�-�͋������Y��9��׶'����r�����j1!;+n�kb���z�Gg��wG�M��m׽om[&�۴��Ƴ5om��Y���׶��[n��=���ke�F�m�۱�mk(��vL�t�pIb��ڷy�5;-"t�qm�^^��v��Xma8�G�ͻXXn��� �f��t:'fw��,��5mؙ���Dnv�u�Z�{�6��l�yۡH���a�^^r�5	�ma���J*�$H����h%�es���|7:'�����(Ȩ���P��Z�H�{����B�r�A��j��y[�܊|'��'�c��d�f@�f��dTA�Ȩ�%
2&�V/<EXG�P���xU:�Ԙ����Bp$ؐF�_U��ܝ�oF�U2dH��� �z����q<�B��9�y�
����j� >�DIB�"J�ٓ�p���k����zV^���(�T?"�D0��n��b�z�B��C���w!�O��H<�H#v�5�&&\W�\��,����N�H ����p���wp���1�����oP�"�D�f߷��R���tz����s\6�+{�	��%<��@����Vf�Q�%�3f��!b�m���ѣqt}�t��
])���b�%EYS�Q�GA��x%����QU�P �_H��_���Ρ@(5��5�Py��� �������=����tz�]`Kk(\U76n6TKi��U�l�6�@���{U|A}B���}�͓��{7Ԙ�;*Q�
9���;`H�zF�"J�Qܳ�U��澠��j�s\6�+{��kcҔ�v	��b2z�5�r�B�2P�"��2P�Ƿ�ɜ�a�4F��������� ����(Ȩ����<���{�L��d�8UOZ�L%�dxN�dT!��Y>ޠ$C��"JD�M��O�~����|�.Y
�Ƹ�ؒ
S�ؿ	ݎt'�U�Q�߯ME�[Ȥy�����܎#R�j�CUN�H��ZS��/��u�z�ߺ�}�Z���ЂR<�R���{S�l�������:6�����/k������>|�>w^��\k<o7]d��#���f�%&�Xi�tC,&�V��N��n6����4�<^w���v�X�V�%0�Ε��3�g%O@�m����c���N�����]��*���O�[������c+��Hj�G\�l��Aˁ'��Б��2�����#��_�{�͇�#�⃻��5��'��vE��QȃK=���T~�\\��MO,�L%�d:�H;��F�=<���ޡ@���JD�_%�zc�����,SOc\q���"N�I$��=Փw!�����꒾�ы8���y�5�>>��'FOT���"��/�^�_���V,�QzI4U�k�o�
�B� ��(șe��_]�m����?\iq��ż���:�뭫*l��u�bWUiZH��<������m
"E�IC}Z3���}��$T�*���QB3P�_/�"�Qi˱�ڻr�?i~�5�r*���5X�a9��S6�E��U٘MA��q�ݜą�&�1|�H���P�-����z��ѱ���xu`y�A5���F��;�f�W�:D�~TAyP �%
2/�W�{8{wQt��k��k���@�A�"A݉%
"Dg�����ʁ}B��/���P�\x���Q���$��,r�3���\_I�	�
+�<;�h�h5�$���Xخ�p<��D�
r$�*�2P�~���F]uņ7F��k�n�m�׮kx���u��wH��M�WY��/Wջ_H���E��jygJa.�n�q��A�I\��%&}@�"�}X����f�ȟ�GG1��.O&��Q�5�$�D��s\��57��H ��> ���}"����L���D��XLiEH��Kǳ��a.�q�/4O�nG�^FW*�Z�սȭ���%_NLsC�����(�(W�/�_\w���H�_la�}����պ�����] ���/����Pg�=9���݉�"��K��1gΐ��M�����Eڼ?j�"rdT~�9[���{	�7b�v^��#��	�9�<]���6.���}�������<�xq�P���\�+�xu�����ve4�<�	�쒾�}�Ȩ,W�����/Jt0ډ��z������L%���#\�2/^�:�us��B��T	�_H�"�����[hz���ws��W�&��r�E�*IT.������z��i�#v|�{�e��u��z\p",�97�^�A]֬�'A_l�J-]r�d�-E��1=��g�<i9��,83N�=��F��:�Hlv
��Dt+���E��d_P����l���Tc��n�wE�&��3:��` �(9��>���|~�c֒�zg�<��u�xٴ<mF]��]aalW_m�N�I`O�ݙ�ݐy�8�so*��������x���rEDd_I�	�
#rg�2���,3�TA���5��{���$]Bp$�ח��u�� ���g* �(Q�}@Ȩj�~�:]$۪��E�7�񘀩�(F쁻~���S�ݺ̞��-�$j��ݑ0����q���>��#"��&-r�C�5D�yPH��Ar���n&`h�"OS�y��
|$]�@I+�$�����<�7��W�{��S35-UW��ث9��U�I�ا����R0�S�'5S|{z���3�?C`��-�e�s�`4��h1�)v[6��`P#�$έc�!c{n�js6�m͊47�ywe��m&�䷅b�gs]=V֬�C,�J˩Q�YVb��q+t&wY���q��^���m��%���}���n�4�0�1��ڂ2����4@n��ذ�sb����ڒ��f�P�8�����>gN�H ��WI�L�vt6�-�cp(�����JD0Ȩ��_W�����`�s>nm�G3���{	GAۉ�N�FE�</�X=j���B�"J�E�%fC�*����w��i���r����|d�@Ȩ�tt=|%K��F"�t��Y����w*��y���{*M�Ηy�F�v�� nؐA�W�(P"@������w����e�%}J$uȐwbO�c�>9�~�����Jh�lܸ�"Z@t�^x��,��1.מb{�(C�}"���ף\�2_=��E�랕���>Α>#ώ�;�'���e��I�ѥ3�����V$W.�d�f���oY���psfK$�sa�v��TJsY.��v����HW:�̪��[	�m��)wcp�L�3�	�_t_H�|D�+�%��QJ��p�[%�%�(�A�"AݏIݏnߤZ���>2j�D��InȐT��X�׋��w�A5� �[�'�uLB'�W��z�A�P"D(Ȉ;�H���p����������\	 �hP2*��%7OT��@���j��U��u�-m�+u� Mn�f�O�'����y��y,ݑ>;�&>;õ�y/!(�(�{���L����e
>��%���@��]ˉi�;�T0��c�%R��ƻ\&������D�����wH��	�H��`?H���Nϊ�(�!��<f�=���혅���aR����-*�"r`�5�h�APw�9�&zj:�ؗ֨�׏Ka�	W|G(wbH;�$��]4�u���"4(�����������	�T�:�Z�O9�����$�ȅ�W�'�{����0�p}�f5��4���$G9F�z}�7W�y�\٢G4�]�ˡ�
˞*<���j��8*JW[�A���nРdTA ȼr��+�ϴ���u�	��=�$�=#vD��ِN�O�v�T�H��CS>�as�3�����	��r$��Z������ĦV�F�����]�Kw%�e>�&s*Fr���i��� ��;�HIU��9L*�xe�'�*_h�����؞��\�k_n�a.�+�"�.qN�#W��ͩ���U�4+Aa{�w7	@�3{.����T&�t�v��ެX<sUF�
"J�A�QJD�ݼ�������P��<ue(�A�ު����E��\Cf�YV�;w2�=~�ͮ4�)vԄQy�uf�B��L�Mlj�`�=��̷��������K\&��U��3)��]�t������Y��H#.
}�R���3j$�yB1z��־���A*�H �H��
��*�k���'�ĀD�QU|d��{������#�=����_x�/���(�d_I��oz�ЄwG���݁ ����1��	�O��r{]����h�$_W�_H���QJdR���9b���!�*�]�׵s�.��\ n����:p2�IX���꣞E�����+��/ՙ}��J�ݰ�"E��o�+CZ�S�Mt[�HV�w�(�V5Y�o�ާ1��7��d3D�G&�b�����-a��q��R�Ra=�6��U�@��ِ�^��@�+L웦�X�s'ZW}6�,It�j���*��e�v��vyI����eN�����˫��:"�5w9�����-��8��v�u����*iUx���{.�;r�*�>TvK5�͍�Hɷj�am�o�F��=֎��LS�H�j�t�F��J����A�JV��oCs7݅L�s��R��r��־%t��t1b�r��SS�=yA���"�+rTƺ���Y�������r��:�oMwwPQ��ĳ����s4WYW�hF�Tu��F�m)x�u,y�^e*��V�6�T[S��ɹ)5����ŠgguA%;i:)�L���f�V/=]U�Wa��\���7�HP.;|�v[��n�6F�q�m9W4�N�z�L��9.�L#s&��-�����/r�8���r�s�1h"q�4��W���W
�*�������	,^��Ԃ��;�7B�hd�_Y#2�x䳸-����Cm���6�6�H�%�cgaڶ�p�665�@%X�E!$m��n�P$����kD���v9�vBFےۣ6�Bvk,���!a�1��y�bv,f�4'����h�d!:D3E�]�)ɗ��(�l����{ݜ���4�K��r)�%p���k6�rd��';;�.EdݝlŨQ{h�"�Ӆ儑��n��%��Dm�E6:6��{;�=�B���Ѳ�Z���y6쵡��i��q8�"[d��I8㵫kkV;d��l��{E�tM��Kke��pe�ى��H�4�#��ŋ̕�e�9�g	^�ۖٷC���a��Q6�Ƙ�+�r��r� �a��a��W�n��6�h�/9����ݣ�Ϟ��Yͮmwf��x�uׁqӻZ*հ<u���k���Ӑ�#�T�Y�+�u����t�l�]]>�]�� �]Ӛ�d�a�23��:���8���
�v!:x݀C�;=yN��n,=�q�bG�ص]l��4{v�5ؚ�V�uׇ��l�;k�7WV���(kz�Vޙ�暆.h�
̌$�=>E8���tnK��a.L��!�t��e��@���[��|�/ ��G#Mo#����v�xb�FivZ4-qe��[6g(U��B�zr>M܇.�P��Οb]�on��8�<@O)��8���n��z����i�7n��vB�+]�Bp��@]�a���&�%r��\���pԣ�7��ًf��.�-��ΰ�b3�m�`�� � G��X��ՙB�&�ٴ�	�E����٪&���J$�gdl���k�Q�ݖ�]�Mpn�ir�����=�ywj��y*q`6����J�+��p��n�Y�����sX�qa���� �չ����󫙊i��n4�s"B:��1&Ș�hÏ)��������nܡ���8iG�h@x�ķ%T%�m�j.&ݡ�n��!�ۧ�A�=�89�e�眽�3��7����]��ȼ���Ԭ�S^	M���ny��pWc�-�͸����mn���Fv'�]���`��TUf^��K�-�.�qꨢ�t\��v��;O^�PL틣
SmDۏq�R{<[���Q�<�:����{m�����\��ҳKLT
�0uCa�r�Y77��{W'X{M�8� �:��k�<��2t�Y�1�WK�a+E�
�i�!f���ǆf̰f6��l��]>��|~�a�2۔��S9�22��^e4�tЙ�SPj���'��d��|r��v�>e��/c�%[+Z��@-D�Ả��Т��}�P��
#:���pj�
�� �>����b�S��#�. 7�_6���7+�Tz�-[5�f���G�7�}-
#�
���Рm��ͫN��(����wx�dw2�Օ��ԣ�B�1�{P �q ��@��!��fi@̨��w�`�"A�e`�c�s5A�z}GМ��s��<��������>&f�@)��j�lh"av�kX.]t#.��N�}>;�� �mW�ڡ.���OZ��L.���S�s@ �>,��-�����co��|7)y���E\�nC�@���;�r�]���V��5�܂��fwK��r)b�Ƭ,��k��y�=[̧�elpJ$�2=�����&�y�E�}�"|pǈ9�[��긌��e�C��5F��V1�ܒʩ	N��U��:��o�7����d:=�+�ȑ�6Ӿuk�q0�;P��3�My% fX�@̑ ���6���By���W;ñ}�q}@4mQ��}B4�B�J�AmĲܔ�!٭)
]+�h�hY�],�kϾ����#ӑ'Fd��ͳ+�S��}��ڦFhmЯ��B�-|ڲ	mQ>��o�&W�Ǒ݉u7ʟ:�٘�Dqځ$�p�Y1���MO1>ND�-ȟiD6�o+�F�)nߑ��WU��e+�;؝ulǘܤ7Y5~Ô1o=+�8Ys*��<hR�P-l%�ћe-n�aؾ�6��_��k�hz���7`QT�:`��"A{f�����5A�H �DK��ξ�p	��|Z����d{2:�bI"L����}n]�ܴ�� �H#�D�0A�d�Fz̪!w}��B�v�zc��݉/k֌��cfە�&��Y���2�/ԉ#2D����E��+cׅE��md�5�!�-�!��m	#�C|h���f����S����`Br$��u���FQ�)G���@�[^�مjl6k*��}��7���@�hQξf�-Т�w���M�[� ��|r>o��/��d�[A5����p���L�7[�]䥲�|��.{�]E9ڕ�dZ����13�f��E�M��Y]���Ѳ��u.Li5�ĦT7U5RK�����I�nD��������Pw�4c�'"H��<��Ͽ^Ϟ��^��و�Բ��	�"˝&7kٲ��+�F��K�� �����:����;]�m�E�a�Y���4��"J1�B��YDM�����Y ��_�|��i}��M���Ց$a�����@�?lB� 7B�g��}�z����Lw;sT��I�>� �D���Z��҄A(��dH�������l"8�E�	kw��P �B��|���P!����R$�>�(�Y��ݭ�M�����'��E�i{h;�ê�銯��~x�_����V̡�\���B�s����.Ξ�K5�g�̳Ip��g}]YJ*!j���Є
k��<�d��Dn+X;X�b;J�i�@�f�i.Nū-N �t#.���Ŗ[Xm-��D�a�.m�(8�NQe��2���uv�I�٭��v;W=[�hcY���)-���c��502��
/a���X[�W*ɜɠ�1��n7:�o��ϧ�iY��3P�GQf��K��j�M-�u�n����,Y>�@����T8T�s�UA� �Q�ǯ۬�Z��u�[TA-��������wN��*�,��#�ځ$��W���V�X���([�_�W�������-��d�[A5� ��E�G����B��9r��(��9�$۸P���nꃸ���Z�re��3��5|���k�k�ՙ>����g�8��*�,��#�ڀ; Y� ����l���V�X4���D�k����vfq�
:��%ˬ�Z7b�O���<��W����x�������ɝ�uU.���AP ��	mQ	m
���ý|�e�W���wS�7��:�kn�e'����i���^���Ճ����������?=C��1j�yzvs������Q�\�N߸���TA�P!��h�ը�fK�e�wi���>Ɂ��6��P#E��N�'�e�+�B�7�y���ԭ��q �.�a��1Qڨ����([�@E��޳�d���1J�t�(;�>�k�$fK���i�s��׏����)Cj��d�#-"�%�E#�ɘ�f��Ҭ��Nꯈ-|ڰA�S��ƚ��\ D�OL���`��Y@��@��P%��6��޲�`"u}_Bw��^�Ͻ����Z��[LV<�ѡ�4�@�!�Q����2}]dJ�9�B˃U�6��5f쪉�n�Fbw^��{��(`k}����}�P���IB��n�mB�iֹy��M���Cu_�ͫ!����rC����ّ^ �Ȟ������yM����	�Kr��OEv�����P ��-В3*��~�.|H�y}�҇��eԭ�q�TAk���A�}w��j���iң�D��Q)��Mx�b2�7c[v��C�xFYz����"K۸|���˽���Ula�d�F:��A [TA-�g��O��Q��uD��������M���@�A�E�$t�lh9b�s(�ɺ��|�e���{��x�:�ͯOu7u�x�o[T%�@������cp�)Y�fO�j��]ծ]�|'�`�B�PSR髡aٴ�r&r���ی�xb�=K��܊:!��H��T�.*F]�\���ώ@�����_6�X��*��2|���W�Z���r�H ���Vd��'�S�o�ز�ĽWjckƺ즱�h�,nѯ
Ͳ�l���d��`��2��������s�R�=�������X �[TCH�hQ4}��"�w$I{W�wSN�l:��тm �t��_`���wUK��d"ڢ	m�ۼ(�k��/�M�-���Q�@��$�����/�]"A�># C��r�/y��N(�Ww�ڎ�xFQ> ���T� O�$H8Y�ۧ�+�0��=�q����u{a�4}�Fd�|r�����M=ĶE�ո�2��$Ԃ��C<ZU7-�<�۝�n�M-��(_)�fQ�f�:��q�b�7_YF��UѲ��b���Հ�Smn�p`Z\��.#b.ܚ��W��1����n��Î6�$�3�C\����cD���7(�t5��\r���X�j�L�][�L��(��1e�R㷔�n9���ӝ}�����Ok�g�&��������7��fn��pa5F�^��q������0��]L_�%��mQ�����W���	��@���ЎR�D@P:}��̑ ���uj(
ܟ"#����ۭ�[�:��X�)*T(�E�w
����C2}��fHڣ]$ͷY����W�ul��/�Q�|Z���sMm>Z�������� �[^���W���[���
f-�1-�g��
!��K(~n�og�
��޴$oޙ�o��ݽ^���RT*����$��:w�Zy�d��X�!h�K��(-Kj�
P&̄?nP��� [�=/ݛ�n��ح0��w�	��k�Ր@-����]s0���C���7EL�E������e��l=��1�L�N-�h�èp�vҲ5޵�7'.�h�7ںa1� 9H#�D�)L����̯��B�n��G��)�,��1�m��������* ��mY�ڢ@﷍�����Q�t((���<���{A�zOx���b���i�b��ZԿe���3�y��b���x?�bG�+�:^_x��]t7;<M>z_��f��prk* ��[���e���D��"|F@���u&�:��J��B����j�:_g�G�T%�D4�-�$!B	9�;!Ԅp� �\����V��{A_ �>���є�qt�K�� ���X!��@6�f�j3ڪ�2/ �\͆໻Tћw�mYy�Ӝ�yw������:�>Sz�N��ͽ5�����1�TZ�ֻ$��&�����3����Q��,M�왼	cl�ǂ�'��$5v��io�ջ��p���'}U}t��|�տ�ؚy�R�&��Jܛp��v���oVT�n�7�d�GU�)�ډv��)O�"f�4��ϬԵ9�]�RN�(�����*�'F����wnM7˺ �"��/u���r��YGe�gjڼZ�1�vν?a�*��[|@|��V��i���A�]�I=��um���Ia�܄�W�fm�6��u<�v8F_f���]įM��ʉ&����y��m�}zlfn��,�$��iX/��j��֎��n �9&!}�푷�m�h�q3��J��uv�N��q*�{�i���TC��
��#gW�l�)E�W�!������uݨ���CHY�����cÁ��0s8n����iQP���m���m���Y���ꯨJ%<j�+��B�!�a«N��9�iY�W�4	$�3���ofݾ��56��ahk�/gs5�,��m�:�S��sE^�N�(�W�N^LW���3D�ĕ�q'[d^��kw���r	�i�m�� �N�N�-�K����ܳq%���vY6Ե�r9I�-��v���%�k��Y�e��ܽ�����^�����	�vn<זb;-kn�ؤS�m,�D��,7Y��׎�z�ZQ�Z7��v�S�R�E�6��ר�'�Ԭ�m�����6�9�i�y�=�Sۄy�m`�ٜ��&ٶ��w�{�zN�i�jI痬�����R��t�1mc����������9#�3N۰Q��� ���#7Y�N�6�i��Z�u6���I!Gm�ɋY�\�	��֙	�%���ĭ�)ƶ9EĔ��/�����N��yN�Z�B�([�D6�O[+�J8h��$�=9wp�M�WSɕ��w���U&E��_W�b��@��Ck�Hꘋ6OEꨑ�2'��Z���-ڑ[�@�(���W̋0�o۵���M��I٘����H]{"�nc8�ϧ���>9��}��NdN���sq��F�����T�����6Ch���Bnyv�A��}�_ڟp�m�gSɕ���5q$̉�N��,�8�"��}�>�@��8;����R�L�s[ݝC_��C�(����AڠB�Q�:��������گ���#��\kހMT	�]�!hX�h��W�Cj�u�z���l�xo��@��1̷�co�"dv�[��x�]�J��T�Tw"�F���$ːNFd�#0$Ab��p#�}�z�b������M\P �� A-�λ�}0Z�MD��x[��d7:�:�c�i��pc[v���߼#,��2�@A��s]����n\��$O@��wyP~a�������ͫ?6�����Y�sE���1���1�X�yN�V��ϩ6��/r�3hP (��
!���*s�'��R���Lڎj�Ө!�D�U
�����x� �c�%q�*�$�]���/W2�n�h�>&ii�V�@Ǖ�� �j�����@��ߌOkn*�^cv�l>���(}+�l��X���Uz���L��]E�7$79fEY�ժ�X-�ۥ��`e/�$�d��3��`�RW��l�x���e�ƺ���K�6z.g��C�ǲˢ�u�u٦�����m6���:���wG:����Swm9<Wg�-�͗9Un)&Uu��I��N�3��&��7�q��]���:Ku��4qڠ������:�U'M�#���
<+��Ը�m��>��b�K3���4£�h����<K
gG��;�vs��;$���F%��ąc��6�ٴ���i�Ǒ�}E�D4%�(����y�1�{"N;�]X�%̺��рAhQ��㸲}G�kO��̋�����mr�A�f�t\;,oq�0�* {���U2mV��x�x����Rg5
J�|�V�+:�Lڏw�\H ���9�װX9����hP�|��)/Nȿd�eU7+XV��cw�F>�32�d0���u���ؕ&�F��F���F��e�0���<��'-`�.6���,�~/=!{�l��ǟ���C������7j.r� g���v�c��A�RJ���|��ctW*Ü�˛.2X�pq�sf�U���Z�[��;oZ.��$�sS�IQ��e��F�Lq�>� w>c�[��"mG5q> ��dd���f���d� �D�� ��An�|Y�7B��v��M��+����'�eG�
7_Wů�V~*+��Q�
��ڣװdf�����!� A�@��T~5�6#e
6�g�n��ԫ�V_� ���=s��zs�z����}�Ym}@�����8��'���n�qVKt�řX�R-t�w)�7q���D�ݼ�� ��m�)�aZ\�ޑj��f΂t�y
w/���j��|C�\�/���Z�+{ttw7.w�� r_3���Z��%v�(��@�P �� �}_���_OegOT��N�I�1�v���#i����]�+'uhKt7�U�]3`�3YF�+r��T��,��Sb�|��v�U�^?^*#HE�D[_;T�a�¸y!�(�D�Q~�׹��[��ݏI�)�3{�zp�O��[@6���ͮ3v�}��U��t���K����* �5>���7��wJ��δ��¦f��KP��!��f��j�n�y�o����2�>�#��[���il{�d��O%�r��W�j�h/�B��^I�!d�8�2c
��v7x
�����j�YM}�M}G"�Ȓ�d+`��}��PvJ�p�Av��C(���fD�ru�3��J@[~�a��ud4'�����W�ʻ.�z�kF�R���ڷJΟ���l��{�����b�%�zT��ӗʝ=��'&�Um\̚���^?NT|��(�Т����Dz�wjzS8�Ҫ�cw��`�� fX�a�D����������hK(�2��CW3\W�.�Q���²��f�*꺢�	�U��[TA�_L��G�h�q�"y�xZ\��.�Hh"���͡�fO��`"��Y#JD�������{�*� *׾#HE�O<K�E��U,r��(�РY@��zz-}Ώ.ZUZ��n��h�zx���G1QV��3��?6� �ڮ����kC�S#x@>9P$���^M`}��z��s�(���?7@6-��}�&���do��ilqƮ<��#�dB&���Շ�}�5T�=;b�^��_��<g^�5J	�m��d�X�nf>~�ϼ�{��:��c9�a0m�:P�Բ��i�Z�u9�C�lk�Fα��W:�"޲��Nz���q�kkq�aZM!��#R�t��8I�n��;�c�X8Ÿ�V������L�6�cn����(�8BՖ��c��n�y�`�1:�6{/t�lsx!u5�;o���#��w/4M�MK�����؄�f��k��	؅sk�l�"g\>��3|;�kr�-]����G�WŠ�k�������\ҽ�3�T�*���L�)�� � HjD�0�M�{�L��L�L��T�2�e4T,TfsR3�-�f��̶�ilp �����dQ��D2(�s�Ӹ�Q��u��؞«\����@����W"H[>��-� ��E���+lY*|�7�ӽ�b%3ȦF�d��R$�c<�Mw^^|zy�u�jLG@�/k����2�����;T>��w9@�W���o|CA�{����7skc��R��p��[�dp ������m
hx���5x=V-��8o��}�suf�J�3/�@�3�����2��9�5��6����*�qf]N:��¬\���0+�H#3.�ҷ^���r�~�TC?6��Oc��9^�Ǐ�Uo�C�D��ZGj([�_3&B.���>�{ %�3�>={	�sw6�=Ʈ$��s��9�퀼tH ��Q	m
�
,��5�O;afϞ���
�pV7zA4`��3&<���������5��Z���Q˥⮎r��k�X�])m]�6��AȾ�_6��	mY�oI3:�iL���8���A�O�2@̱ ��ϲ�Ʉ�R�����E�^��ؼ~�TA��i�]V+ϔP� cB�-Т�ɾ�=�>Ȅ�*ݏ5z����w;�nݱ��g�"�WwNkQ��D�S�i8������Jn��[
�an���o]���.Ԝ�q[�N]zϭG��$��L�9�����̝���X�]ő뻱wkNh�)ʠO�e���_s���sgVU�[A+�K��`��z�ќ�o(�]݊�����j���}���/9zdފ�.w�Sq�ɱ�>;u뻟]���^���ڸp%���D�g87��G�+G4�q�Qd���b�U0�9]��x�˖���>�����Y|3'��+�.���OfR\�IY����*�MQ�	��G��VF��)q�@��r�q��ů���vL���j3�T(ؽ�zC^U�WdnΚ��nޛ���Yq�	q��sd䮻����Z�2z�%���{�_ݮ��h�;�L���	��RmF�ͶG��~�n�\]ǅ�z���w=-��olHՇ"tz��w"����@.�h���b�wWl�K�܎]w�M�A���>ۀ���wV�f�Y���إ/8C{�U Y��Y�UU,��6��0�O{�=ݕ��{=)�tl,����W������"$czl:�;�)���]���-ky��=g�_��??Y���n�����Uu�$~?�!m !!#�~�n�ԈMFQq�D��z0~X3F8�LHHBR4� cH?�	 ���`S��y���xh+��g�P�2�(���` BBG�17ᅽ�K��|����#��S��/�&�9��rz�jqXE�j�Q�JJ�[�_�BO$�xe^mb��������>��Ƿޟ� ��� ���IA����!		��&�	I�<���G����P/��H?�����{�C�2��K�p|? ���p?(���b�E?SB�F}�F�J
��g�������bQ��`">3Hϧ�}~>Dޟ�>r�T�Q?1����������ǧ�hc� ���/��0m<��F�PI�iD�����G�C����@HH�
b�Y_Dy���Q��?���P����â1���%������B�����]�
��=�� $$g�r����G�{�����G���A���8�ĠV��#�������x�Q�@�E�^���>}
�������� !!#н�����M���<e��ԍ��9H�F��/$�!!#)�� $$~�� ������%�"Ƈ���fB2/�Q�$!!"��D����)R?L�����$$$$1����%�=aA�c��<�L8d!�{�W(*��A�h�F��LjB��HHڐ��ϑ��KԏX �������LC�/��[G�~��>��<�N���y�A?��<b�'��$~g�/o~������}ǥ�}^��  BBG��/<�O7�7�" ����� �� !!"�r�OJO����7������8�B</0Ry��q�X�	J �~�`cJR����b��/��݆k�ƾ��z��~��5%��<��|W�@$$|=Ǭ�o����ϔ{�R43����/08���x����	@~�dK����H���)�}D�J�U�}OB�_��������҆�A����g)҄�4��J���yl��H�w�|կ���"�(H~�\� 