BZh91AY&SY�����_�`q���#� ?���b?��� ;�U��X�U��41}��Z���L�L�I���Q�J�4� �D�@LT���m@���2�A�R!��kL)m����Vkj�XQ6�[���e��i)�fk3L��k+3+fe�m�c*�ДKf��ʵ���jiRZ٦*F�ٶ�-!�-����@c坫EU�5*��*�K365m)1��Vi��j��ٖ�Vm���U�fm�l��U��je��M���iT�S)�,�f��jRɪ-�V5������R�ɢ�+� ��}���9ڀf������Z�xẪ����w=܎��V^�kz�]��nW�[n��e��i�Z��Ų+�����h�[7v�Kh���ٵKV�S�  �|*��3�nJ��J���t��Jo#9J�$��{��@V�W{�xzU"*�s۽SL����)��	���*�%t�q��zJ��<�=C�ZZ�sv���R	t�o�  ��{iT��F���i*REz�*���窥�W��J��Kt����B�ۃ�(-����=RP�N�^�)R�TUwqI^۶�y�Y�mmj�$�E��)��O�  ��R�)=��x�=J��z�t�H(��W���jB�罶��4ҕK�z��T�U)�芗m
y��ޤ�
���m�A)WM+8�zP�ҡ/ux*&-�&�J��ȵ��O�  e���*��|�Е�*���:ԥTR���
��'�;��h�]m�j�R��UGr\V�M)]��JT�T���BjR��=��IZ�N����l�/s��UhѭRھ  i��vЩJ���*UU�R��ޥ*S�֜�R��W�I=�ǏzJ���z�z�*
W��yU)
Uw��r����=�ޅ-4�Vꗰ�U��mM-�m�ڭ�P�  ���j����^J�������R��{����ҕ*�י�JPU^�r�TF��W�IU)S���w�J^�]��{^���JBY�w����=3T�L��ƶ�iTͱG�   �}]P(����PQ��q�-�Gu.� Q����Ǡ=�.z(Ӯ��\��Y���U@������u����\�����j�[R�-�m�h��/�  ����S����V ����)��sm��'�y�j�g�@��f��U �<����Us�8���S�z��(���(٨�[eh�7�  Z�>�mG�J�]�Y�׀����W�M�Ei���g�^zC^�m\h �K�47a��( � (  ���2�*��4�44� �{M�%*�0  M0 �{%*� F�2CB)�&����      �~$����7�h4�0 0I�����O%?M��'�h�S�O���Q��[���4T�sO΢��I\�ҫɥ>�N�.e������n\�.��}�}�}����{�o���cmm���Ccm���|��A�6����=���?���?�����{�?�m���w�eV 6��}3�Y����o?w��}ތ�8M����߈�7��~��7�86��~B�!�����!��{� {������c����C�@��v7��Lm�8�{�l�`Ǹ� <m�m�	��<��=�`��m��0^�7�C�&��|� >c���8� ��`>c���� |������plBm������{���oq6 q����86�{�|�loq67��l{����loq6Ǹ�7��� �q��8 �}��! }��@���|Ϸ�q�ƽf��0r
�0�j����qVV1����I���x=\��FW�f=UY��/���1P�S6���:e�����\�g7�aJw{��@�Ua���� % �ZC-�pE������X�g��NNq�hlìf��K��ms�"w۵뛏���_]�j�b����زYˀL�m�X��=����)VM�Ы.GvЊ�	�Of\��yHVHk��7N;��*O{����b��e�q�4����e6�N��P-x����}������)�)e��i*�o
�X��I#���֦v�G6j'v��wt�wau��\EN�\�V^��V�m[�X�+�*�
�Uu	�r�X�8��R�۷��� �������Rf�L/P)���@P5�Q�D��qВ�7�a��,�2Ar��J�%.}���>wF����εK45���45:I�:U���f�n���p�yo9b��K��D��A�����8�в��<�1�1�v!�F%Dsfhky��8����%�;��Q�2�n�1�\�FY��i�[�h�VV	Q�ka�V�P��5h�u%�J�h
�-���-(�B�X�J�`h�T�ňr�f�n��Ճ��g��D�)�!�skR)JNl�����xv�Ͳ��m˕�	R���F�P�\<`��4n��҂2N�K���yi�tD��]އ�F��ڙHus�qjѼM�0��ۀ�g�ִچ��{K�׵sqվEG�8���'�R�*�Y{�w{v�	�ʏ&�Z�������A��:L�u��v��0Y���G*�h���%x�`9��h��FoUpeÐ�;V�J��`���A��0��j���)�un�T:�f�Uiٷ��Hs��:�@ӡ����c�_Q��ތ2G>P�+ۖ14OQ�l�_-�.�k�M:�MӮ�|���ePӺxgb��B�LǇ��dYh��Р�s%�1^�se��4�x}
g>)W�6m���4�;C�£TqPK)+��X���0�yͶtB�(�SpT�����F���6�S�4�~6hS[V��	�
��E�;@�@mE��ԥ$VH�C+hjU���"7)���z�&u9�v�Pq��W�:М����lEf�ძNY��1���;M:��GPɣ��{!=�q��j��__|{+��/��#� �PA�ob;/5L	�d�Z�ƜC��S�m�I(�̈�d�
�Ċ�pA�7xow%B�p{��c��^�j=�gr[G,�BbN���Գ�
 �ؘ�N���7rͭ�e�Z��ǑB�V��S8�Yù�bы����n֢W�5�v���v�28��ɷ.����M�yY[i֝��3h��Y�m��M���K�g�Q���,�cjə��͆���H�):�2sN�#mrO�x%�73�u�2WRVWXᗟq������Z��˦$��	��W��[�=���ֺ��'�*MU+T@6��d���f��0�²6et���g+�ðC�9���J��T)V��=�PeZ����7[M�{�V�������Wh���1�7����,�G�v-Ǝ!	/n�mԍR����a��'$�&5�nd��ީ��d�a �F��H�5,l��9�U-���kXN��i�X�"в��<�罬�uڢ���5����P8�IUh��J�ۆ]�E�}�ݖE�J�ę��w��k1�ǒ���LET����}*��8��b�&��s�i�1�M�hń�xqIGt�p�����" ��Ι� ��p )�j5�0�ᨸw��L�f��K
��7���j��9�,HE/��#����[�԰�ٷ�5i���xz��[f��rB���o
Ą�(V��42�!���:����xi�}c\v�`7&�X����wW4��U욃���;��M'����~�@�H�)���= Z�����a�X� ���\���v�N�~%��546��}�uD�+�+O)�߷�� ��h1�jף���BTY8�oj�͸)e�>�Z��x�օ8"zk��,ts	��&ڍ�*�V���e�\|�鳅�r4N����d�J�g`
��΃(�_|wI04��A��NP���6�Yj-[̡�����.�)�"pAi)�j-Ø�� 8 vc�hWx�,G���i[Ķ��i��]
Ԛ��4[�,�Z��*w)nӆ*�st�rE�X2Ѯ^����;�GrJ�Cer൅׮l��Ӕ�.�.��E�_��Dړ"�REH#��zC��#�w&,�����E�36u -�8o�DRġ[�4s�O
c��6������ Ф��^a<7���S�u����V덦��6�n���:*	#�f�Z�y���{t�k���J7���Pޘ�\�Y��"3FV��0�a-�n���0ޜ�6b�,���I�"1Z1�"m
%��aO6���t�OcZ��A���/�BY9���e�Ҏ��IM��yE��+�,w(���;�5 ��[���Z��G�R�sd�jU0]�ɇJᯇ	�uw.K_7~h^%�23�;uצ2�!�݊eu��pwWO��tbz�j�X]��}���.x.�n)�\,��C��QS\u*�ް�Ɇ���vx	%nޜr�h�I�kD�`k��M�\"-�4nՑpژ�;��f#z�������dܨc(n�uoe�J׻7^��Q����>��:�̽�^�nhs�P�q����t*����uίGFdJ��8�+*و.��4�u�`H�w++sLŤ)n�G�X!�����ڱ yB�"�M��¾�v��;�i�=o}���;d�d]{�oE(
-.LAk#�@�6�}%�΁���3y�ݽ�D 6nv�.�80{E��s!cc�%5����( �k��U͝��XŸvj4��`o�ݍE���GqV䢷.j��*2隖$w`�(�e��T�yx�3W)�oI�ɒ�Ʌã�f+x����]�Ĉ٢+��kX��D+��e8 ��L�������9L�|���s]�^�ׂ��۴���}����f��Bj�D�<,U��h%4Y���Yݔ,��md���/.
�8�e�jYq��JC�(���fk���ȧJ�-xD�y�u�E��c/QT��g8�)�i����`c7�� _!��8ڐA^�6��'q�q9l�ۂB8E�y�p>[)	��n�&��n-���4�<)wo-���Y�PS�L�@a�4j8Ǵg
��+^E7�ek�m.��'���[w���k`���߮�e(2�jʇ,4t1)n��j�r�s��<�@n�x��pt�Zr�p�(v�}w�S�8�!! &�5�iURQVȅ�4�q�hC�++�4��H0$ݭT �0mwjO@��Wʇ<4�g����7Z*\K�,^ j� �6����&k�J
W!8q�Xͼ)T�J��r�a�b�;����_�e*��1Nɖ�l�J�ÓZ�L�����0������q���N����\�2�YA����6˭Y�b5�8��s�qmְ>�������E��B���� �{�� �6["�,@���-�ϮG1���׆�x�E,Cɕ��a����M��+�A�v^SC������9�
a��Q��D�M7˿H�ǳI��p���{�U�_���`�.�.%�]�m9+�2Pm��0_uǨ�q�s&f���wIܙGb��E�c��Z�7���l����Bbm�dY2��۬� �I��z��̵��V&���*:�A\��=��n��q�I �4�"��+é���Ie�;��b����B�\b]�&�:7.�׌���X��:t��m꒜&=��K�1Jv$8Jחq�<�;Z�	�sS ���b��D�WxFX��.7z�׳UH�b��9��Q&��l��h�<(V]�� ��m���Q�4	�8,�9��^�/U�&�/;��<Mҷ�co��U�����&�;2���pP�(�Z�!����}�ۻyڱmY�u,qB�'�D5�4f�{�ѐ#�u�٦�eɡ�H	�v�3:RR= 	�C��p"�����K��uQ3sQ��t�у����M="�M�}��h����ߚ������
.N+��=Of����p|4NX���,F�K�E��GHM@Fc�[W�F�c{�z��+�4��Pa��[��t�QϺv���ß��H��1��bj,�s(�ڂi<5��o��<�]���W��Y�K�d�O"{6�B9��-�fZv)iL��̏]Df	3s[N�j �B���s��I�9Z�pf�p��Fko����F���K=wFO�zPV�Ů�S��#th�\�d���P��'in�����`��+R���'̓k#l1�F������!z�Z�m��NI�%�w!�S�JS�٬�Ws�ʺ����bEPs5����|]�C�RS뜛}�VԺ�y�q���Q��ӆ��t�.Hj)}N�:��^A1oTsr��Z��(��Z'�;�m�7̲��grc�
c�J��0�j˭��ve��.-�wZ���o�!x5�ޒ?�.R�s����pࣷ��e���8$��RL1��~S^.�Ӛph��1op�R��/����bђ��4`�H�Q�Vw�`9����3j�d\�����,�aU�*6(V57\dKX��ǩ�j ��z.c�5Q�;���ܑvB*�MB�k�keۮ0I��b�G"�Z7�`�����Fͺ�c�n>C�p
����5��r�t��4.����i��4%�z�J&'�9K�(;�uÌ0n%p۹gry�|����A��a��3P����׎�q9}R������r v ,Im�3�)�n[���cnGq�z�*��2b�T�@#����7tlDh��Ն悆5����t6�N�,	�Q�UYN�"�bB��v�6�7GMĄU�u	�� ��r7��-�h�[/���m(5M��u����өFExd�����A����m�P
݁�eֻ֭e���ڎ)�U�N	G7d��
29�a!&��k!fa�l�v�$�N�̧�H&&}�7	v"�>pd�T��@�g|��<�u���׫3�2Ϣ֮a@e҂��[#wP�TR�n&���܊�ф<o��Α�ӎ�7�M��\-9��\�NܚD�(�d�I�����8dr�N��a��H�����d�'�/
G(��sD����J��L�&�q���*W�3A�XD����44́)����ph{p�-<�36U�V�sn�ے�Zt1m=�ͨ�&�+�X2��A���f���/�j|�V���֞��\y�Y�n��J�g~�/��4�M����j�8������#x���b�m©����両ٜ��H�	�{r�pm !�5��T;\�ov��4�"B�]�'Tw. k���(5bUe��+#��L7Z�s ��x��t��7��ZwvH�����m�k*n	«xot���2���AP�/o5JlF�-��Swf�GhZ,!�\���6��ʰ�?tB�i��
�-�m�I�͂�̸"�7{�O$���Pw^���������`�݌lXMKgr�xk
�px:E�+��W��0J����{�9��;q9���v���b	� �G�pH�(��T��ԫ[c �{7R̺{> �8vfc@Ep(�\�zhZ�@�TK��aې,�hԽy�2�*��Ɏ�S�D�	�@�JJe�� ڇ �e�Z�\!v�Gy��#�.�k�k����ue��
��ͭv�0Z0N_QNq���g�.�� �!:�W|��N��7Wr��`�+N(ᨌ��\�d8��y�5k�pF&�=�Q�b��%��[Jf�ySe�e��v�qb�B����
� o���6V\V%������V���||8�f���Aָ�<|��`{ז*�)�N��9�dq��T��d�E�4s�j�r�hZgb�Y�m �fO�Q`���,��e�*=�$�z^��i8���w���jKY%�PT��c�2�Do(�Ә�Rmf��5g"dS�Z�MQJ����w՗kM����i���5:WYP�*N��0�<7Yo"�ю�X��p�X�P��%��|�o-�[�5q��j�e���3w7�m�=ssb�/%���{��&�0Q6>lq��9��΄�uO��`8���S��ٺ�D�F��/N��s(�-��(��yš���+�ܤr����X�(`��9C�b�r�B� �7plb��l�Ϋ:��.��8������V΍w��P�M3��xU^ �ظf��"�Nq%ˍ�⭄MV�ep`�ܩ� J�5�iS�7nP�j��N�ݓX�0���Q��[|�Y�õݚ&0��0�'�+i�¬>U�h�v�U�Þ7�3w�Z���0�O�&ǃ��[�(�]�bM-�xqs	�cf��M�ױh4k$Ѱ۷�m�XE���r�j��ց�����)X�X�0Sǲ۹��-���%�b�Ȧ���@`�P�ٱ���S��f�B�'�g"�GRΏ������+�<�J�"��y�j4-K��[[dm��4%+r]	����-b\
����L�ъH߸�јo�Ӿ�JW^`.�N�f�����$%�Ubto7(��V�+q=�a(I�VT�h�2)W���x��������q�������8���O����D^^����eޣ�u�\���R�Rc<�����{��Z!��`�F)�=�%ښqO�X�"gCcz��.��J�KNs�|	# �TXSHW���<�DY�8�~�z P�!XO���y�*�˷����N=R_:e�+��4{n	Gd�dc�7Ƕ'B��w&2;�R*	�6�Ν��S7����±�f�:�{�/��W\<>��
��"�L�gk�G�;L7HRu���:d*Y�8%7���v�~wD+p�(>�vTf񺽱b��Ap�J�"�Y���gQx�T!���R�D�֩N��uA0;7��t+*l���3j,Ύ�0-�8�K1_>�7�Ӽ�j�NĴŞD��gXr؍�-�0�s�rc�Cɓ��]8��#�#=ݤ]^Y��^�ق^C1����J�_5���t�S܊�s"l��Ҭ��xV�	��*PIa4h%�Zy�E<�3�x�s�w��A�)��Ա#��3�F��7u����Q�/�y�M^�tK}���#Tg/K%�J�]Clp��q$��/z�߬���$�q
�X���ۗ0p��+���E�uͼ�.��Ǻ�	1�ۣj.�-̈́�
�������wt��{13pn\ܽD���&Q���[��a�$��#l�%e��Mq�P�֙�_��5��D�w��̣x7�϶m�>=��W���[����
�(J�,�֋����@<�`XF! ���Ļ���zcC�yUOoP ���i����j�;l񗆣��)W�,�9��̰��j��ݒ��~�@����H�87�0�.��`:fu��Gt���F�ϙ��ʸ@����p��5(�{}"X]��el�Ӎ�y0�IB�Չ��!6�����j�rBS�9Sh�hH/7/�yWD�M�NV+U5�� a��k�Ų4�������i�ʢ�ɩ�	�ES�TWy0�M�R�:���֑�ݔ��3}�{��ޤkÂ �A�S��mN���n��SD��\�4�r����/[�虽>�ǀ�����}�Ņ��e�i�t�P�T��3�v��ڭ�y,�*h깛���A[#�q��0KЯ:Q�3��לJ��اc��Uz��O_�4��2�Cg�#x�2u��`�V�U�nB�V\O���%jU�=�b�cF):��������ɯ��7�.��Ĳ�.�tǰS�l��y��v�EPt�81�LP�y�!F�͇���%5��`�ػ]�����r�2 �=�-}4��w�^M��;��A��VG�Մo���e�2͛�[n^;5t/��� �+������|�[�\�	;�&;2� 
!�Ew{GJ{q�Z�q��7=́��[�3�T��[d�4�f��
�G�{���q��\z`8�O�T��5���ư;.�%�;)�9:�ۛB>V�P�Zj��9�խ��sq�5GY�%����d*�X-��jQhJ��9��ha�1�5������!Cnv9\~�{�t�4e���;p���^�^����C�cyc�ei���Ic����~�F���Mh��,��f,,���q<�{
w�!v�-p�˥i��-i���i"�=�T�D����y��f`��3��|#ս	��{�\��V�l�8F�g-
{��ko�z��k���$�1'X��}!��V��o왖x�0�����C��\+JU��c�����+�Z+k��+��Z�U5̬�B��ë��|[��*'�q�^0:����䷝$���M]���;�*7]��m<N��Ի�p��ێ��h�� ���\�϶�i����y�z�e,`�!����G
|���g �r��
�H��+i�r�,{�%�\s�(�H��A�v�س3x��R��03w�{�p�!�:n��Û6*��I8���)r;;N�WK��'d��
W��=f�+�pVEn���5)0˓y�z�ݰ��]GD�8h�#�c�.`�H�y��C{ã6p�*;e�6	�v� �<��Î��b��mL�#	�;�t�8V�M�nS��[N��T�m��a�����'nE�Vݻ̑���޷+q�t��4��!����D4zv�H^��w��EV�3w�zd�h�;�e^�e��1�u���kaKtww��D���v�|��'`Q��x��3f{6��~4F�%�J;7[1�Y��Rl�<4r�
[�|��n�qvEc�{����-�AtD"��ޡ3�2��e���t�����{�'��x��=��;�˸ d��c���bPk�j2�mC��i��,�ބ*��YɄL�>x�8l�`�æWr�,��7��}�L��aEm��t՜�e���\N.����
�]^�m#�f���`����c}�Q��vo-�,�ʢ�$y���W�U��"{�T[173���Rw��)g��������gh.������[�Ftƫ~���%&��z�h��%��i��=Y-s+�k<;���w�6Ἆ�����Ǚ]�`MÖɣF�=�d�^t2�Sənn �gd;+U�y̝_i킊ۏ�r�g�h��[#�G_V�̓�Dw��{'��!�=�Y3\�I/o����l�����F��ϧs}L�6������v^�2`�wF��d�φNz&�j��z73���%��;G��=�b����u��"�iʙa�����k���P���:��!��E��S8JQ��J����BE���Fkj����%�����2s:����U�5	�e$��*+�==�	3��UH�h�RK58R�-�U�6DlH�o3�K��4oWL6)�g\ƚ���w9�S�3,Ljnpx0�}n���	W�{'�����6�I����76���E�a���2�3re�Ehd%I���[�3K8
�$�Y�8'�h��e^'�v����5<<�w�kC��9I�n���B>��(E�^�$1Ge��a�C�kҊ�h{��8!� ��GA���w���!��>��4���dU���sI�m_��4n/��\}t!��ܔU�d��<"^���R֖%���{f̦�U��`C6���Bܝl��u���Yp_�wW�v�S�I$m���*q��`:¦�iem�2e��)�:�P�0��`�	ƍ8o
C�J��ˡ�����X��裴����䜷���G�z�b�I7�f�d�x�X�mŠ���v��I_<�0�Æ����<��G�;�y�'e;Z�u��M�S���EB��ⶕ�U�Q'A�V0�6l�b�����^6{G�^��δp\���=�f�]�hG��a�vCS僻t�H�r �P�s���>�^*�oG�چ�圣Rp�g��>����oؑtx�;W�j)+�$�e�AP f��ݡ˶���>��1p�u�.�Z�xf�L�lu��_�w�;o+�6�y�<���U��_^; 9gQ������*��U�Jfsv)�.��)�ޘ�]�ˎ�3�uL��P��c�2Ց��؜���^�CA������t�H�ҍY6ʚ�Iԥꭼ.�ډ�*��U��l��:;mp8�jT�eCW���K(u�⺺WAmf�×��4y��F:�j������s;qNl�X�Wr�������=��EF��r{�z���-#��5��L]�ԙ��]l5\�1�ef���^��2��+��*�SU5Z�;�S��s9%�|��6*��Ҁ�Φ��^ѷ5�*�t��23��v�3��D*�ч�_]J��WD��6/tx�ѷ��8�����*Eۼ�g��g�R(��qnG]Wf�ИK��b�s䥱"(4'\�A���rڨ�[�kE��V�x��s���3ؽ(�������mm
���}\L���V�8�]�㳥�Ja���ǣ`�ɁIY:U5b�Md�6,�,���u��s9��f;f���9��#R<�1㓋v>��W��sI�j��:$Mg4{OLs�\vlH���w��H3���Y���۷&��1�ݾ~"sˋ�m��o���ɝv�+���B���0
��p� �~�{�^y���R�{صs� �q�X(=���J��`��gx��ku������r����=�\�j�w�I{����)��[�q�1�����b��=V0e=}��; �RO^�&�æ���������FI,5��xw�V�gk�[�����o8�U4N�����7�y31�y�x�m�a"���3�n�:y�{��q��&V-�HT������G��<�Gn�巯U�N�w"z�@N����	3���m���+�pʑZ����u\��6d�dƤ�����hD�fYN�/.}�r�gR2�}�܎�T�ֶJU�rPgq*�ڻ!��f�D��s�;��� �?cY�^���s�p�Z��K3�H*�:�l�]�Sx^�r[{�]q���P��8���Z|�����Hi��+��1��F��sS�V^ֵ�r�'s��M��l��;�l�i�A���Q�aR���fT< �p�&����\n��<X�>�E��dc{AVS5�ַ�6��C)U�xq��TCi^��XD� �WRY��k]%6�1�ݚ�2�N=۽~�U�4��Q:���8.��,נ�pN�Qj��ቡy��ThC�w�?e��[��ir��LV�c����bZ2�:�I�-���3z*��<�մTX��U�lJQ��=�L�yʝ8�1���T�_7��@�w��|G�>SՃ�L�ͣ7=z ��m�	%����Di�Gn�ӗ2�ʕc��ݲ�<��	49 �]ɺAWfٺ��^���e�1�6�.Ke��Dly��;��t�j���]r��	L�2�ۻ�+>�HB_hOeh��/�ZO�A�z���@��{�uf��C��0T仗s�ͧv6��;��3*=�#y�@�:��dU
���ۓ{f�ª�O��pS�2�&�����T������C$�{A(���������\���=�2���k�Jg2i�Z�y/&��][+��
�SkR��}:��i��H-p�Ė�Уo.��޹���^��n�����қ���\��n�	����'F��ҩ��Y��.���b�<�Z��v9qֹ���;Ml	h)���~�V Q�Ǵ�I/>�НcЩ�(�f��P��
�l4�w��	���krW�k�_�0��nz�yٿY�	S���+�q���u=Df�ז�Vn*dE:�4�)}ʚ�:XU�i�f�g|��ǗOz���ɓ��9�Q�]��ͮIIܘ�S�j����+T����"����G�<�}�I���>�'=#�
S�zi���-g\4�I��z�%w��S�R��
�5���0�����vJ�˩f9ћ��_��W�~M��N��Ņ���z<2ɑ�����O��Ҟ��|�~�3�����YG�F��S�;�D�n����\J�2밇�)���6�:���
�nŖ�ѭ&ad7���*Y����&�+����+������<ڴ�ś-��_~^}��?npH�g�v�O.IܖgP�E���f�s4����`�S,ɥ�5��'���]��&�^xl�n�R��7�)n[.RH�KA %���(v5F��FF�+�j��˝���ʚ��*s�;��,FX6�"o�9��a�RV���.5ׂH�B%�{}� ��x$6v4��;<)�ev(9;@Vһ^|�y�[�x��v�	���q�����(�:��6����ɝ7^L���8ދ�%�R�\���3z�e'��2��8��ݛ�S��������D9��wN�"�H���P1�W���u]�M�����ƞ� ��.�'�8q��H���R��1��I�l�ghuՁ�Xۿ��55�V�IP2��GQh�%1.�3�8���p�vGe.ӵ�蝮����e"�Ad���#��<��.��Y����H�޳B��K�-��x��������Ìt�/�cN�w�o/�R���1�$m� ��;*o̦-tw���h����Y���˽y��M������HG"a�J}٫��e���]�Hi]V�P#��/�uth{ژ^�=pR}tuEN���RK	G�Ξ|Ov�{�%�2
_�^���%5�RX2 ����F�n�g]I�V�&<��E�i��]n��u���z�e���%����!�9kKh�_�js�㒱��"�c(%?W�qT�C�3u"��l#�;S<�'�^�n}{u��4����n���q��W���ֻ�{�xF!w����uR������\�2=����H2�^�}�6Z�ݚm�љ����5�f��)�)��BY���`2��tg��Wmk�^�[��˗xo���ܬ:�PGC:����Q�4`���Y��}�����b���,�)	"�t���2�������L�3�H��O!�HR�ì,�{}�vؙrun����s���
�ї{O�M��ι����SS�&9|�%˚C�3��,��vɀ����f�E���8tc<�@$�#�wok�*e�}��[ۘl�9�뒈t܏�!PQ|��0�o)N.��5��-',��/o%��]95;�w���a�O%�F�"�qj:f�wl	����T�x�F�h�Sa6=�����(��j��o���>���o=�懓�I�|�t#��=����2�t�N+K5CǙ|>.۵y�,#����v��T�μ�&ː�e',�0̢)�ji����]�z�-W�I��d\�\\�to\�f,beҎ�b�Xi��.Bd�l	��iU��9*ʚ�!$�J]��[n����]+U�get�-�r�y�k��o��`o>nn0#��R��Z�t���,��y��kY�̠�.�+p��e���ާ��Չ�Ջ/}ɀ& �Np{~!��O.ZX�i��@��d)�c���n�rbf	>x��T�R����1������0m���O�����?�{�ck�����O��?O�ߝ���?���UƳ�P*_J/)�Lf�o�nK�z���+�U�/��&r�%3Ӏ�w�;	R�W�c[{ͻ֏*���ו1Y����s�p�T�i������kޤf��7�T<��1'ʃG�Z�/�f���cR&WP�G��a$h�{����s~@��#Ƿ�kbu�ݽ���ܭ�̂K�zV�;D^P�Q��u��[�y���\ƳaP1�:����a��̡m�U^X��M4�֯��hc�7�⇊��hht�:G/{S�e��ᐩ����6�X��ʤ������a7�ѩKɒ)Љ�s�٫�d]�C+�I���rEV-�o��
ގY��� ����k��V�il\���pg)�zs*�sT�ɖ�Jߤ�m�jn>�Y�a���0y��S]�C�3�I0�<~��F����C�)шx�u�.m[tʡή:A��d�9%����n�(�6{�)��.Y��	�uԊ��\�<fw%�v�L�6N���f6��D&)�q2�H�]v�$��Le��h�HT�p�~4R�y�o;���o3镌˻K-��C��dK��M޹}7\A#�3sL\f\|�U�-��k�U|�M�S�
<V�of����#.���ۡ���m����4bE[�*�ܛ���A�<�x����s
����"$K�̚�-�Վ�f,Y�n2�����ϙ�»�:Tj�`�ѮO�\=�7b��&;7�y�fL�1,�w�!ۣ�/wf݌H��<%�5�j�xn�ho��E�*r����r�#��aY��Q�*�ͮ1)+n�-N�urO��ڹ�6�fڜ����Ŵ^�[B	�d�NΡ���5t8�1=�.�v�{�]^Bd�N�-�hBK��vf"��+�ӗs���� �V^��%��Yzr�ө�)n�B�ΘJ�Ʈ�3nhMβ�.�8�bT�B�0e>���-�wb&r�~�h�Z֏���C��g��ed��� +0ܭ;�ӺAվ��qyt�;}�M�m�ڻ6`�t�m<��6M�[f��
ܣ�V�I�S��T*��ͤk��˘�7�+VM��*k8��.���]�R��1�d�qfS�m��w�KN��$�X�t:�n���>��2M�Ja�a��<�����؎M�0���IW*��8{<��w���!fK�h����VGv�ޫ�;�u��|��%�%�K�KJ��6uL%<o����wr��L��6n�u+Tt2�ժ.��=��Q��mK�%Iu��n���F���ɓ:�������y�q,���{���/C�f�Y�;p��M)ʗ{��Yr��K���2�kn�S��u��;(&�w	̒vp-�S6n)�[՜Zy�'B���GsUBn�X�ާ��������%ᕙH����rܘ[YKz�^�7GJ��$!�p�ǒ�Qįk{F�&n=8�3��~l���P�Ģ�����TX����1hܙ$~�Gq�kQ�8#�\�D�����f�� @�1�'��Q���(�̝�KZ71�ks��5��\i��n�Q��,���O	��b8}��1]��s�5<|�qخ�dC+�a<W�}sgnB9��*�\e�)��ܠ�T*u;���+�3z�ժZ{$j�Ў�*�VҮ���1�����8�nk�6$�Қ�;f��TX��'Sk��d��fv\��pwv�!�)���"���w�Fr��.!�9�C�:�YS9�dt���[Y���l����8�Sp�����m��~yO�;���T�$���`���"��s����j�>Z]v'EL�6�<��VqF�r�֕�އ*����p�v��������.k�����v�.08�]�����ST��N��ճ�N�vt�����ǡ�qЌ,BW�ٹ�v#��+��|����+��F��4>|�k�k�����Լ�p��I�,L�s� 7�m��zH��r��B���ZGsW;�	���vlo c8>u��ZT��(rq��W�/�7P�.�&z��FJo��sَ�)�X�Ҧ���ޝr�W�0�}��ᷧ��Q;kV�0�%;)�;NS��&9��2E����8s�^�W�}��уmuP	u��8\&�I}���^�tjB�m&mke5�:	p�wG:��Jj���Sƴc)������4�|$ʚ����*�5C��єb!c�������+�xc�����+��)�ua�)y;��.p�}�rN��༡�s�^\]���K3�	�Y��8�nh�'n�3m���q�t�E Z��`pϊΣI�֓;}X���+��B\䷢�n!]T+qXQQǕ��b�Vn�o��:�V0�0��'w�������vt���R�	*�;�\!�M�=K�6c�2��8��"�pV/8��}g�ø}���)h��C�h�1	N�\PWA|�&T��P�Ե���`�Y}���L�iq��sd����"1��'�=�.&81�}ݪ=&[ӻ������J㢄B�y<~h�v��\�n��4WNQ��v�κkf�rH�۔�-�].���i]:נ³��-�2%��=c7ݞ�$[z=�\���!eݎt���)u빭"�JW�v�q���Ԣu����_�m h���ź9�F�����[Dt��=R�����*@-͑^�sM��4ȖN��
�B����^�[Լ!{��*����p<����"��]���v̷�P�/S<�n]j.]c	���v�X�͍i���a�\0�8h�鹹Ft�t2��y&�q][.5��L�g�u�Pb�������)h` tf�k����?_�3;�UA�SylH�͔�Jw;��/v�$����x:|�*�V�Lc��1Y9�BK�Z�:3��ݚ�E;�S�%|Û�*c��ʆL�v�Q��	w��ݻV�OT�s(�H�*�����9��\Ð*�z雂i��3EL�= 4����n�4�t�k�<7O]���78�0�m���VBe�;
��V��A>�>(Rpx�4HW�y�n�!{E|�KΗ|2�� a��>��w�B��`�7|�B�;����v��ܚu��t�����!��׵�ru�eD0�Ug%o�m�-�{���p\���O:*E[�}�K ��}���H0��v�9�+�=�(O�z�0�[�[\��w��.��f��"Rj��W�#ϲ���:���>������؁�Ђ���&��b���W�l�����.ARo`�vu�]���+7m^T�,1<�Xu-�a�@��8�okl"���)"�u����ܕј�d�yL���Z�.���-^n�����T:�e�f�X�^�0[���/3���Ķ� �%}g9�<�9t)�c��ӄ?a��,���]Ke�[���u*Vx1�E��;2��t"��hֹ$l:����@u�O�pU�nZnV!�qj��u�T��T(�A�bs��죮%E�,�i�a硇�c���\��ӫ�W�-�qH�Y�"�aX��I�2
ս�"�z�&� �8@�|��d�'�����_������[���g���%��|�)�s���z�@�
V��Z�#8�u����͙\�q��0�,M���%�,d�^*�,� �: U��{d�y�z�ݱ�P����xKW�]ޏ=�vz�>�V2��#hn;uwc����er�żZw����s}�ь8.*_k�=2処��|���6��LAr��w�cό|���S.y�)��C����G-wxpu�kE��ivnv�e�N"]s��FJ���!���k#OU]\�!Σ�[��(d4(K���h-�Vz%;:�V̥��ͺB�hΣS���~.D��,��Fٹ�OfM��K�җ��V�K�JO���Y;b���v�7�jE���xί��H��Vd6��qY\I	����f�ձ��RRR�L���ܳ�g�� E�d��w�,W]���jtJ�j����F�.}.�:�0����&�4GU�ɂ��;��]�u.�>�Gw��XH �rop�%]ǓT$�ʃ��F�ʀ���瓡���zQjD���G3����F#��~kG�6ric��'.NO�q
wLZ����x op�=�q{�!:Ve[����Y��園�G��������۳*��\׌�3�^CO*+#㷙X�Wi�c]`IG(�I�+���wAYn�������n��(;&�fY��Fq8D�o��y�`Է�w���s�-A�g�W3���-�VOe;�G<���Wn2U�m�C���6��B����gb��dT��雽9�a�w�=W
���c��IP��xS����Ob��)v蘊ޑ�ԊM/$�\=B���_&=��<F�SS��%}�;�$=�A@������`�sps{������ټ�ԓ&�8\���fR�����\��y+{Z�R�.r)=]B��r��U�[:����r��\��z��8���+�++�ʛ��S�
�����g����s:�=\w�<���9�Aǆ\�/2+���A��	8�ϫ�ݖ��DltM�ou�C��J�CJd����4�/V�a|�h�
�B�1G|_*�Iݭ:�vi�(zN�u�iD$�J��t�fF�ݎ�^��5^�o�B�7{f��c�ӭa�}]���/��n���bW�������`a���b��Y�̱µ���8�?(���{W�:ʔ${-� �J͘�kN�8]�őg�6d�&S�]��0آPd��qY���Ύ(,�	��t�����W����ܵ�[N���P��r��q�k,*>2����b;AP�ܟ*���z��{ ��Ut`��,�p�7�I)0���_e��(�%��#4x�|��<���'���@�W��Յ�n�`�x�v��W�ʉ=��c^:�hq�է��r$��2�)�����,�-�����r�{ʦ����:b�C�Py�.�|zѤb��cs�`Ile!1<�ƌ����Wx&ΤxM�j�wy���2Jw!�]�:5��&�����a�;5]75:���v��i��Z8S���j�=����`�����k�ńz�J2.�y��P�e �n�ؾ�f��yp�[��w�W�8�t�ausp5W�:īL��٧B�r:���mu�2� ��+������|/�OV��QF���jH�C;5�]۽Dւ�+�ڻM����P�畖�G��������{˫����I�w�m��$)0w�,�t,J����&2
�)@���­����pd/�1�M^����w�m���f�il��1F\ӽ��ޱ��kz��ے<&ʨ������L1�����ϐ�4Ui�Ɨ�;�ݛ�w��T�$@�t��c^�K�cG�E�O��ʙsB�PU:��uܖ���޸���Y&��<�Y��pB��rG`٫!���0N��z^�[�I7�a�ӭ�(p	_t���,���9Ko�ST�ct�ߟ`�/$�Ч�M��Ma٫���L-
~W��ݏ�������X��ś��]@Q*� yWM̩G6fw,�n;K���|@٢�z�P�6��^.h���]Y:�;���@A�t>]������n�,LPq2�c�3��L��lqډ�y��H��Kj�+<�*�m�8D��N�d��x^�g$ɩ��,1��>�Yhu�[d����B�;[m( ��n�=.s۟\�x	Z��m]e:v�j���.ӷ����s�ZGJC#d���sk���tcç����7��#�z�\�������޼�_%�0�H�7kZZ�Y|dIae�By��/1ïH�q���ܾ��fcy��ކ�9%�mN;Y9��Lٺ߻s�-C��e欘������`�3�4܅�x먲ׇ�<q�|x �zdZ��Mʚx��%���(P���,1�jx���Wm��p|y��A�/[�=��6�"l��V.�c������u��k:|�cُ�:l�9p��kU�"8��C���+o�m��0�(X��ʛ�ef�{% �F��ʼ��3��6��t_I&��j�ώ2�k@.f�գ*Bk��ث��#Q���{����YZ����M�ņ�C�f�x���~�����*��7U�q~>
w��gv�\;[Ǹu�;5Ԣ�n٠�ʅ��\�2RH�Ƭ��W=�/V�1j A��dN��.��ocJ^��"�\;���+�{���b������ļ�:�g�<� �XDٙv���68�N��p��DܥrW^nL
�wy�c�߂ށM]}���5ԣJ#pK�r����`�@�5oTMp9��Gs.�K������
zRp3��V�m.���qi j�NY�⫨eu+�GN��"&Ʒ*Qٴ"�/;�i]].�#��9�9�A�^obkM���NmS���;3�Gm:+izmH��J�Umo)M%���y��O��,�^�ir@�r ?O]��&驵{���	<(�n��ϣ`��Z���m�s���+�K�d��Щ��Tp�ȺN!�z��������x�7�'1iN���.�Bm<�W��^:�R�;�[�ա�a�[�u��D���*�UYk�X+of7J]݁F��d'�r��ڮ�̍�U��>��1	<C3�٧��N= ��m�0��ޤ��)3�6���#�z!�i�|�:9v��9.=�-���>O{췘P4�ClnR�(wE�f����I�Z������ �r�P��"2r̲ґ�:��f_�vu Q�LEV�Z��0��ά閛�Z�](I����l��Ŏ���j�B�Bt�fLl��R�G:�$�
�`F�*��Zt��H=ĺf�x��ʡr��c=
�7X�ߍʵ9Z+`�.�3<ٸ��*�4T��gMv�A:'+� ���+yg<z�۞��� �H���yå�'����}���?{�?/���w�?�����~�����~�����P���4O�\}�Y��a���,��b�ݟA��6��G��$խ�6�F�{��e�Թ<�=eK�ƯQ��V�/_<��&U��$w8�G��9��`�qc\��x5?��]��6Lk	i�h��O���[��t2�	�������P�\�D���U8ܢ�m{���pU�v6P�[b�s��z�,v�rJ^�s��R����ioO@�p��3�+^��N����&���������nS��u7\*�f��L�.��)U��xs	[:��sX��[�4J�[!u�/�J�\ͱrbͶGe@rD~o�n*�ˠ.��N�r鍡*K�Z%�j�ߡ�["�&Ę�!�_����n�}�bkځ�Ӄ:�P��c�z��ƹ�[.j����e�;n��
���)�sH}w�W�����NޗE	�De���$���@��썕'��N �_��ԟP˥��Ʊ��[s�e3;����a�;X�S����a������*��T��ʳB[�Sa{�y*���ڰ��Gy
w������.��7+S����[7�ٚ��(��^�����z�Y:����%t�3��`]�z��C�)ϯ�����C�=˗5�^������B�[�n�u<i�/*��t,T�o��ΠG�v
�u�R�%Լ��9�bi���|0NS�D�N�Vo'ARQFɱ.���kd+ufV���yɤ��3��9�/n���8�K�>d�Ş��|B �Ĝ�AQ�W(���7D'!aK�\F�$�)��DTOL3;"��r��
i��mC"��L(����PfW(�G%�r=AB�r�s��!AQ�����\�ԣ:y#�u��r.s�䨅A�wX\��u«��ES�s�4x�NN�iAAG�dEޒW"�G� �*�p��d"���h�I�r�;�VeE&='� ��UN�z��(*��֌��Y����)ò�*Q��S�d<N�r�����s��]��zqȧ��輧9G"(��뻔QT+J��קeޟB�9DQs���eY!�+��]�&s��Z	B�Y�EȪ����TG�y�y#	A���&]�
������&��򷤲4݆� ��0�L]o.��E���V�}V���{������ZTS���o���S3�����s��P��5Ȭ�I�V��6>���8�V����f/'Y>d��亽[q�,�K�+�}���,��%ю�n��TX�u';{�_����ڊϐ��{>�!�ck�\�RF��gH�^�)s}=�ӣ7�NA�X�x;��zl���nu�I,Ԓ����V�^ܬ��=�^'�k�#ʹ}�+����2��+���Ǜ��xͯy�6?R^�^H�{��l�W��dXB�J$SV6����le����������*��*�{o۹�6�\d/��2/�;e�Bj[�AJ=��n�}H�Sڇ�⾓�7��%{[5��~�t>����`���/$�F��B�`z��EoU,�����j��XF�}�}J����r��K��>��2��
�k"�������ڳҽ��g�T~fÕ�}����/(��^u�vM�{ju�n7�3k����S6Cuuf�b~ޮ�l�mV�V:W�W�*�V9��:�T6�=�7K�%K�Qe�rT4yr.�ƹn�d���;5����E���#�5ս�u���F�I�]�����cn�jqn�ll/T��j4�^ڹ��԰���S5�yZʝ��Rʝ��qy���{1?Q�+���d��P�\�-�4b�8�S9"�u�Gj�w�g��a��W����g�!�+WCC�R�q���ccD�I�7SGY�[d>h9d���}^~e��g�}��71=^ط��Cf�����,����Y�]�5�&�/m_z���<s�I��w�!L~k��� ��[�l���Z�Z*
�/|%�X[[�=�o�g ����j��z<���eNZ�bT�7��s,ٕ�#B�)`����N-��Ux�>��8/b)5J�o�z�3���"gs/L+0@���<<%.�����ۿ;���"ȗj�I�[;�/��~��H��sF\� H�jR�C��
�ŉ}��xȃ�kwo�����]�s�ύy6jN����O����{#s���Dq�uxΛ���"��s�:��yH��ojG����mK�Ew�X��f��m#�r�^��>���G�0!���K�Y$%,Lk+[sM�qp��t�Huտ��<F1����S1zЙ ���7�f�=�f\�}���%gպ�����[&:��b�ϧy�����ү����܇�TU�:d���(w{�7����Ytպ{K27��S^{�M��>�{Y�<�y��)���2M�+��Я;t��t�
�/�d���3i�j�5���p;A�|�oӵ=��Wk��L�6�����O]3:���S|R'���p5��C��^�¹��a����Q�<�z��T�T�K�SD]�t6��Q6Tw��Gb=}丅=h�P������3����,1e��zNx�:�P˼��R��{��שn����TBE���y�U���D�_�Ҽ�CZ{B�J�n�v�m���b�ܐ�hj��T��ݮ��w���B�*�c���5ݮ��y{��RA|y���a��A�����MzoK��*���a�C+�?a�~��{��x+�������V�k�9�4�ӉJO�d.|&����ĂdkB��4wȿd;�R�����l�_.�y���^���<;쪿O�y@J<ܡ�#wuc��+��| �^�w_�0���0%>7}2�t���.� ���;ȱ�<��\A�[�o�}���vo	7c��#�j�~��{|<��Y�x��G'WU��4����Z]\nj�Rp:�O)�޲%{���e�qX�Agu%�Z4�U�jc�\5��^\�Mz��d��{�(j�+<,�B��ѩ#I�)+Ѱ��=o�Yﰚe��<���h�c<#�-܎�8;m%�G.Ci{�]����z<s��O�ɾ��у�������J��krҽ��3���g�=S�sK^p��}7֏ї�;yuҼ�So�ڨt͋�ގ�s�#��9[���s7ސ�z �.��Ut�]y�8j�/��ٮ�9R�K���Ì��[p{����V��K��U���<^�
_\��L�z����m��\-q	��"�z�����{ON�?r�%Z�[�x�ΟX�{���k���{򩾡-9�l����丩��ą�U�m�8�:��|�k�$�8(W��me����w.��;5��J`�3JT�ܩ��7?���W��d˜�\pT�HNe��C���x�=��3��P�Ɛ���n�.J+�Ķ+Bws��X<���C���0y�v��5W��-!�{އq�g	���WY������<r�:Q:6L׳s�9-ѻ�{9�����k�e���1��Ы�N���vf\r�J	z?���Jݡ#�o�����{�s��҉����C���(�z�e�����[�y�J$�f��D�w�����@��	b@���+j���	D�����ux�P�m�(��z���[�����/���T���e�=~��U�2���YcO���Wo�f��}G���ڬXͿW�Ozo��׌���_K��$����{�}��c?qꊪϽKgž�5�GRE.K}3�����U���8�P�=�n}NX5�G�Q|GW�˔�ty�y���v�Av�ٱ�{��Qw���Qr���K$�ݼ�e��7yS�*6wޚ;1ףޭ���K�-���[>5�Ó&!K�Ͻ^��ם��[�_�	�~z�c���~ee�����@�:��Ӿ�9^�Y��%�	�x�PI�3�x�1�0��x���Y��y} �EEV��Etd��.�6102Ȼ �o3{):��+Z(+v�	�c�k��.V]��40�](m��=�����ᾑ=܋�H�Uo7-�.҈^Sv;Հx�)w-��
�N�=B�������j�ӧ}梫^�����z�w��]V[��Gv�Y�|`"��L�U�H��Y�R�^yuﶤ˦*�/D�mc��g�ԏ�jzM����.䇂���zN�\�o�#����b~oT�*�k&M^�>�W��_����W� ȓOc���=��Ķ�����ຄ�J<�I��u�:��K�{$Շf�M�F�OF�ɡ��P�\�l��b'�p!�c{�b�]��u�I�e'�ΦUN���7F�/p��<�B�YCF3`^��|g���s�W�.��ճ��-�&�%`$P��0}k6����=��\��<�����=��L�{��n�b�1�ԏ��+ˌV��ȍ>����d��Չ�V&'u)��]��b�g��:8N��'����ސ���U�9Y�B��G�~&���z����������M#r&i.pu`�XV\��C�{�����洀�G�׋0�l���1-u)�ӕ�Zx�;�T�>�QN���W��k��8y��0`��X����|wyk�Z���K���N|lʿ�D�`������hG�f��@�W�ި+�7&{�K�I;"�~5Iت5��RY��W��*���^���XcB8��T�)/W �D��u�{�ЩZ�>�sݱ.�`�^�9槅�g�G���N�o=������&�IҺ״�Ε��ZO�%|��O�O�1�"n���������t�p3'od�d�[�^i�8�b���f�&̮d���W^yBS�Y�{�<^�����.�v(1�"n5^���z���j�z����8���VC�&�bӈN��=�=��.:����}����s~��V�=cL���6��<���	�k�n���kݹ�s�p��f�^[#/~��2�(@���,��C+`l���35��R���:Ƕ�^���]�)�\�{BY�w�ڰ�³��'��>�ܮ�˵��hЊ0�L��=��dƲ��r=���C{<��sN�#J�;{Kd��Zl���m�yHW���1�x�^q#
�y�C,�L��745Qm�I���3`�J��\gYt^u��ؕ9EZq̾TlqR,\@�y#JN���R�{+�Z�����YʊE������{#�Jٱzf�v��sZR�{���ճ*�>~�S��߫��&��HX�PU|�U\M���P����]���/=��J�k���Ғ�^�q�{եb��d�U�������ծ�S�����<"��eu{�$|�%{�v�ء
��GX'�k��z�fױ��yJ�.ȿ�NX�3�A"�{�U�(�;�p{���JTtwv�����?W���u)]Ine�6̣�����9u�ڻ:�]QN<.�pW�"I�s�@����$�Z�)$cNg������N�lЪ���Y���p���*w���Cs��m%�秶��|<�ib�����q�����g�ЕcD��m������{'S����V�k�^��Y+�s�9��/��rد�Q�����z���)��c>�P鑞�g�	L���g��U�B�h����h�3S^�
��.��猂*�7�s�)]�F�E	&�~�xID��x1�3�����E�r86��1>��y���m���e���5�B-U����Q��I�v��� ���]Q���(Pvgh��
n͆E'Sջ��f��۹���j5�tk�U�F�m�Ѣ�EOz�|VG�ɜ(m��ܵ����U��*�t3�է)�!K֡�C��K�U�
��F���s@��zM�z?>�f��[𖊸L���9��o����%_3B��Hב���/zOW�ޢ��=�`��c��=�\v��X�I�����W����f�$�F����R�<i
K-�K��~�;b�絽�_ފ���̥�>�LU��=�g/N��9(��������b�ՉC�����8;���3���T=WY�yX+���{9	�VRJ���n����A%h{��+��Vѕ`3c��e��Y�V�rT��Oʶ��<|W{�t�^�}�{9���.�_ע�&}�:"�&<��p���$����0f��Ǯп�<��V�Ѩ,?w%c}����`T�u� �!L�:�b���*�˕�7@���,m\R��ʝ��%dH-���g���̋��	/�'�&*"�v\ŀ�b����j7k�Y��N�{+1t���{�1���r���FlZ;�6�����
j��vLԲ��[�����������5f$*P̊Hnp��[b5��wNm2}8c\Ly�*�����O�C����vz������>�sl�jr�Nȭ7�x�yv�(G�R϶mZK�ֳ{�ƕ!YR�>�{��2�+�����w4���>W�R����2�{_��d�l}�j�2&�Ѣ��۬��e��P���Cts�gs1i��^�;�l�=���>p
g��M_��u��m���X��s��]�����?"}퇡�����uY[����Y�j���s;D�]㧥���y�0���h�`�@���*"�qϷ������Hs2W����O�Q�T�c6ob���{�����/��
�%�e�4�:���sz9Lm�؂k&�a�Ѽ�NY�����rQ�԰���|�zH̛o='J.�O.�Gg�~*3T|3({"�;g�E	���2�uu/�b������ڃ��҈�9-�}wa(�c��q�ѭ��c��Pu�)�*S�.���1�5b�rh��F p��{�����q�<��F���������3���_���R1yn\2���,S��
q�/b����gd̽.fZ���V�J��9nf��be%��HM����>q@՜��f��Tf�.�Ԝ�o@%*��*�/�e[1��X-�=��y�����ugκ�r�8�Y�0�;1-G5�x�5� �����<�sOm�
u�N�FiLg&�<��b��ı����2�;y����]ڴ����8�踎�Jӎu��3L��wQ�u��j"p�(���p_Ip��YE��|���s���+�⦯y�P��ݩ�3xA�B����tx�ф������Pᣖ�;�|f��#WCZ�'� �1-#��7.8���������8���p���!�1��|d��u��$٘<�c�0����ԡnicdjW0͒���5h�4c����u��� p�8��rugH�ɴ�esf�_!����N���2�r�ft�"�'��rY�(��
�"�i�eZ8�rȔ�V�� v��rp�31�aB�n��h�uo8Qa��Ŵ��O� � ����v��,E�ع@�=��v��WՔT@����OגW*�ea��m�A�q�͚V�"�{4���I�;���-H j��.ڥqe^*�,�`#���W�p���s	��5V�Ɖ���@�gfR�8jE�O��-�M�@<��{ݜֲ�;�^����ͺ7=^�:�B�n��N8O�ݵ-�JpQjB�k`y+u���s,�$������4�_oVϞ��I%�0.��~���z� t�.���+�Z�|���E�L�v��
A�c�Xh�5�Y����mr���CS�I�w:�����GN�|n-�f�(�y/Nu+�ck�h�R���|Zs�b�Ox�z`@N{<5�m�Z�l��^ܼ��
����z��	CM��l�-e�����ԅt��g+3�F+q�}ڧ��F��}�ׯ���K��w t=�x��֜�;])��%ح�C=�e^}$z��B�b�:�Q�}+Q&q��.�{ԭm�j�'O�e=���X���W��ֳo�Tp�f,c���/�e�s��c{��&L�M�KaO���䥆���kB����2;����YN���G��;Ŕ���+s��`nn#��3�2$�y<�A��[���ϧ�2o�B
�����9u�/����%���#-�Eq	e飴u���}�28����#/6kmbc�$h���#kbϑw��q��xV~4V;J�*`�é��7��A��8Ft�,WH3n�S�Q�bg�U�p�)��E�"�dr���t��{�|�|��]d4/���>���������vn뜈Q׼mN�.��L,�V:��ܤ0]��#�R&tb��=��;1h���G�&i�ƹID���Rv%q���y�M�t��$?�/�ŽG��r�os���0>��=k�18s�W�]�<�ѻ�=+�=?9��%D\�Q3��Ur3�f}Pɘ�\��MԞZ�.�W�!ԱJ�̽��Ȣ*�z��aȉΔw<�wk)�Er�H��Eݹr�z$9\��T��D/���w��QE\�"��&p��E��*+1j==�L�"yFI�����e
��98�p�<vRI30���0��w^=��99�xK(啺hf���>Y�tN�ʧ:w�y�w��D�QU|y{H�1�x;��C�惝˗x�!>8�z�W���^�r�����r��y�U^w��ȒDM�V��]S:RIAEW���Ƞ���r'$yC0�b_T*�$�D���H�A"���V�!Q-�q�����`z=��cL��%�.b ��)1%>���Y�&�v��t�j>�=A�ţxM��r���}^�x��<�z�)��5�-����t��J[͊��4f,< d}}Tjx�Uļ��2Wx�	w����:�*pjr�k6q.�wk?DQ�E�xxC�U"l�9����TJ^뇗�R�F�nW���xyAO�����+������*�-��\��{���dc���5��P�]a��������}כ'�ri��������!v�����$�Y��}_fp��x�Nu���	]bڳw��^��.�d0+z=�~�آ=�ꔘ�z��T��1Q�
��E�lI�w���z���}���r�=��rߡ����ܪ��ڳ��>J�I�RW/J`k�~��MTG��ae`��P�����2���~��D�[���J�r�P�|�.20
�_A�r�x`U�t^�ץ=���Ǧ��%�j	܇����Dv��f{�ܫ[��P��{a��[��Tr`s�ރ���}���� P��}BP�F��{o�T�uQ���O�V9��!�Ji��j��҆z�]E�GFv\x���ϔ��G<0֌B>�p{D�9y}�3��=�AuZ�������OF��f�7�R�1�����pv�i6[�'_C��+��If����C��E|���
������+B��o��c���=Q�2�m	�&���NWNLYX����B������4XL�*�Uw�f�}��٘��V`C8I;�}_4�&y��z���R�_wܩ*9�~H�e�<<��.鿪a�#ă��Ճ�%{]t���=�Y���mo�yWt�g˫����̸�0EͲ
Ь�4+��kM>��5&'6.�Z�ݕ�B�t�<iW}�~��;�S[tW�J�şx��!OxO�8����AV���;���-�Y}�gU�EC��r�f�����?���0q����<=.�'H�E�=������.-yMvWQ]��4xc����lt7�`GJ�u���s��qc�)!���{,�8�UD�)��׷���@��P�`!��Oގ��3�g%m}}?{���i�xy�A�u�ƮS�0���wD��6�TgW�(����?�k�<F��ި��#-���@vv�{r#&|�Ο�A�ٯ�H�OQ���M]V�z�+�b�NF�P(>�m]���n]����ת����r]L9�ϼ��8�T=MD���}Ʋ���P��I�W^�n�1qy�"̪̀�ɍph��װ��^��D�1ӟ%E���/>d��w&3��ʗ�Ǘ��_�K޹`3o�C�����<�x���vr���ڄҾ#��͡��+?�os!��.�w�����Ur�<}ľ�p"�ln�B"����uh)��g�	k^�Ę��1�#��Tho]���m�An���wQ��졑�r�����mqO��_@N���0�Q�p@ʍ8|>=Ӓ�ܼm��܌���c�gs}�s҇s7������\~W����迩}��oA즎�c+a��s��=@�u�z�����d*�sy��}�,u��6B��:��JdX�'��4c��z9d�h�� ����2d���j6E����Ֆ��\|���6z���_���_��{^�` KX�0]�P�A�^�~��V���l?^fMJ/==њ���z+��n1|�;�N����=�%���B
�@.��FlDm�$�%�x�ك��{zИ9,i�����*��3e@8���{uL�gإ��4��mE��qI�1*����a�s�.6>���~�c�Oݨ�x[��z�N'INC�jG>�J�w<��9���zcO{{��	�f��F��#�Wi�����kd,s�v_�����������c�w������͐v_)l}�!'�XDX<D��VX�A=˳9�n����:��{ڇy�5�to0D��K'if6�}���1%j����5��a֨�ܨ����څ��7N��	�5~��t�)�(L&sA��1�J�����S��FxKS�>��ݧ���l�o`�s��x�t*��h�v�vH��U�K,�d�%A�a�\9<S�^W90a��q�3�a� _2�0�С
E�1|kc�+d��:����k�%���ew�fe������{I3ΰ'��hX7��`v�3m�'��%3��45|�Q�~�Z+><��:ϱ���W�Tb�:n��L?���ݖ��wة�%���^G℻��y����u����Xꊘ�ӊOi���wd]/x�Mt^��.v�*b3b�wޑ+z�N,�m�Uq�V�{r�u�}��Cаъ�����S�{��GDs�V<jŹ:<��+)��E�)�.�VMvĬ�6�R��c�J,`�&!xc�{+�h1���<ŸJ�8�Q���av�cے��q|���d;��fȒ�\�I��[�.X����Em@�)�2�>�!��t��q�������:�n_�h�#���x+s�{�3��+/�Y4�ؕ���u�=F�r���T`E�G5e2�����R�ue��?*FUɩ�_H��;�z
b&-����dע��wp�M��tq�{k� ��|Ў]��*��F|�(D>�S�~r.D����d�����gv���^����>��3�˗�#~����H�	2�N:�4�>ڐ}�C�����Tӧ�c��t���9����OB�l����[�]�z9��C��2e>����BU�Jf�i�ș�c�MD��-�>��e龗�S����XChqx�.T���.j���(��
YѺY��!��F,�6b���
;�J������=,�ym��x����('���6>#��/g��1������x��%��WW�ט����rx�#�W��#�j�_��	�k��� ��c	���\b��7�Eo��4ˍ�5��^�:�����6�ŏ?���q{���d�v��ˈd*�X%`CHVj�O֯UmU��{1��pVb��.:y�1����
k�BJB������VB�;L.��b,��lUm�xz�Q��!M�b��ޟ#[�ߒ"�@u%*lI�sW1�:2�}{"��yj��RD�ɓ��k�K*Ǥ�c�Ńu����͜^\\tݬ�Q�n?7�0Z�R&(ި�V���#�s��S��ԢS:YRh`��z�yk�~*O�n�\و�V�=�O�P������-՛$�;�����&{�P�S=`���C�7���xe������M��~��@�[q��U_MP��x��V\����]^����JNO�Xr=�X��;�b�G�c�@�\�z1WD�7UY�6��g��*�r���Va�\fUu/����<�'�����m���Yy��2�xr���@:��Yrbs���E�*zhA���#��g50q�൧4�X*-��ug0އy�݅"�v�>�1�+���ܡ1����"YV�fP���	��0{!�6P˷}=*!Cۯ8&WN���Yr���R&�qƬ�eY��SU>��]���v�])�A޷�4幅4�-�̺�\dew��=&��CX�\P��]�f�yw�|1�~��G��b8��0��ԋ\YnT͹M�����ѽ��)���/iw>ʫ�HS����
_�`�$1�C��H9��B�m��]�X^�r~J��?o�gb��l��k��0��X%+0+q��C�6�шEÃز%����tf�c��s�4��W.��fX�U-,şr����"��Dp�6~!f(h��~�A�{W�P��F:f6в�P�*>��NF`�ANTx5�y6˿��q����2
����j��K�����b�p�s�qJ)u��Y�׾��8�������E�(�����3��guM�,�D�U�l]{����c�8ؿ�WF��5x����!inB�*��8����q�%��d��_�������2�,���E�� 0銏F���=vd��"��|��-�C�a���e^��7.c��/������(����BLhA�bk���m�~���vJ�w��w��Ty-��ZկT�F��Qu��GGM^/(�CW����A�[����b,`����`܈׸QW���bs"��!"�@�^0�c�����>jM��DR�d೰�)9S1)B5p�֩i�^T�f-8��x����S�7��Q ��xq$�����j�i��*U���f՘��1��?o�!IT����鼚D��j��((��ګި���u+s��WD5Qʰ함�<C��\��R�8���olQ^��=�LI\��H�*>t�.ۓ,�J}�}t�wB��� eڰ����~��g�0��p�h�$��C��y�Wz��#p��:·?m����Ǣ�'ag�h��޽��O��=LG�Ӂ*.^4Ay�%�0_e�3�jK�񖡙���[motS��W��{ρ�܏���pG�Q�	�ǹb��~���~��W���G��G�1�����E.wDu9/<2(����ц����=����u����l��{�ʛG��z�X��b=`�#�D,��3�ʸ4z�0�z.�<x�AJ��1�&ě�3�x�3{��~U<mt���R�!fv�ۑ�P��*AQc���s��|�gP|,Y�
�
�(M���5�~oK�H��nŖ��7(Mmפh�	�[V�g7��=9�.}�os6�gE��/.�s2:=��F���#�1gʭl�ęP1�t;A���	�?t��.&����l��|��.�&kպ\ɲ���Z
TG��I��
��_�o�����ez+���w�+���ڷ���Q�/C��؈Af�3,B�!/8	U�ml�k5S]��59�# ��3��5�Z�2�M��}\^]7=y϶t�=�� Z4���)Y/�F��.�r���>�=�Oq�[�@���X'�E���g���#���{#�)�}8�%9��f�9�wv,��]5��6�JD8W���B|���C�;J�}3���X�켏N�wt���v����3�=7��1ʂ"W����
��\G��],�/�Or�̂r�uAqy�F�e��qޜ�u{m��ޛS��{$��6����$�P-BO��XU��~~�D`���O84�n�</sϮ-�o7� W�X�����#CJ�-h���Fj���Z&�:n����n���7!��q�7rvLw��V�6&������^�Ļ��y���-���<�מS1�����]�$1�^�:���뙌3�n2
�a��K�6-0�["~Y#}[����������\?z�Ʋ�H�F%	��
�熚L�װ�^���<Ÿ�|����Ȏ�D��/�IԻӌ/���?nE��/Jf>�5ɎB4*�;�j-��q~�i!��FWE�[;u~˜�n���z������#u��ѹ4�ʤ���P>k�*e��{�U�x�i�}uۮZg�8�em���e���9�Ț�����Ժd+R�*�aD��3$׼3�����S���3;��0�0�ܟ]�^���ru>َ:ӁER�àd4N�,��f�K��K6�њz�,)�3+;n�d�m��}�ҳ�_G�Vwܲ�������nXSPԧ�FwGb
��
f/}aYp5�N��W��{,:����*`z���^�-��^.���.\͵/��a�����e\�恵�p���ܬ2Z���́�{�������-p��۩�y��Ľ�w=;����r�F%�|�T��r��1��.�	O����p��#M�-]d�i�2�N:�atn�7�01㹝WY4%��.�b�{�R�yl!�z����k��ƺ�Pa�W�KTr�]똧��ꢯ.�W
���{��������!ll
�0���6�Ȩd�'�/Q����F�A.��z�pS�>L��d���>5%��	|�Dx)
�ږǯ_���w,߶�N�)_B��/�j:Q�ؘ��j{��ք����)_eW���_:��\P�z���1G͛�s}����-�m�:��֩O�"!nߠ:�	SbHlPb��1jtd���&��"*��u��������j�\�<0l!�Q`�d79�͜^��3�Y3B��[��6�=�8���-�=��}=ȝ�);��V��s0&�-c��.�أ�q`e�Ŭ��������
P�{���{ʙv�����a����ܺ��泣��nc�T]r7�`2�~y�����!}܏���s�s 8���殻T�c���������,R��������C�C�mW�xe����]Ƅ8�����֥�ysf#p����̺ۺ^l�ڼ���Ȅ}F���e�?��i_��!*�����������-��ج��>�蕛/}�=o����{lp<g��,�F�U+�Aƪ6���xU�~Q��_u�K�;����KD�yX`י�3�Ð��7-�\'m���R��RW(�|��V�B��)Ď���}���NxvGe8^Tn/,q˺}*���X0���#w����v��h^��V���ٚ�k{�=üMD�Q�^�g�0��n�.�m��Qr��u��r3����{f���s�$���̌7ju_*�x�����/р�ˊ>�;}��㐍n}NZ�/զﴭ�>q��5���U���'�z������\8=�@�@�#���r;g,��#���J1���5`��R~J���%'/�~HⲈ�m�b��<�x^d@���kĳ�7{%
���X1��l�f�nTy�Fm<g熢7ë&b;��� �	C�A�35����~�@"anP��]�X鳟G��/�_-2WvC���Ѓ%Y�GU̇�s;��f}]��̋���_1�}�hq���&)�����4V͕Ϟ`��j��;N�\uc5���qQ�����J�ܣصk,vO!�{ �]�q�^�c[�^Y�u~]ӂ�<_�ᑱ�=�v�b5,���\��/�ۜﮢs��$���"�|��A
��^�H�ԂsqU��]uf"�JX�W��֝�ݨn�j�V.�Mt��3�^[I��Z��o@�\Vv@�z+}�̳�i���ISP+�mzi����m%�l����{ϯ�9
�ֳd3�W��������Cz;o'� J�@�J�������U�Գ�bH�J�:�k�m����'�8|yL�,�΄$ǉQ�`���y�k:�t�g:��gz�hJ��u��a�v�=6䗀9t�+�ϟd#�[���n��c�i��w��j��JC7�xz]YE	6iSV�t��S��7�i��*����J�84����
����QjEM�L�?J��GY7O��ۚ�<}fe���&i������;g�fI��ih��א�e�&�~�؇���Ɔ�{��E�U�X�M�غ4�3�\��]r�����zpx�5�����50���1c�iz7,^�)`�A�l�Ld�C�>�N������-�v�@��&����S��1`�]3��vܳ�6��[+MoD)��k�7Hfg)�w�P�xa��[����-[���bՐ�c֪�K�᧸�œ�vh��!#ǁ�7`���Z{/Q����6�3��$�|NA�ev�u(S�2=�{1���)�c�zvS���8r��V�Q�Ǘ3�,�޻�=�cm�/`]r_*l���>1�c.��3&����&[u�~��Z�ֶM���|�<��E�ұ�y"z-�A7u��^n6�ꃭ���p]�w���c48	���dx�/���ë KdCc��b�T$��ƃ�՗9��<*ѭ�Q9�|7.��"8��%��>/T3.��:o15oŵ�]v�m(��Q����Ï.u�H�hCڕ���"/�ʥ���pX]�y���cܴ�CJ\����͒����uc3V�L���3�cY#_D����<�&����b�U�^Tr��<�{N�rD�*4m��`�ʋ�wk�y�f�R�|9�y�)"�=�����k�m줮ҍ r�6�Q�O
=f�[�y'������N�Z���;���5��Y]�fT�SkAu/����.��6>��S�:Qru�SCfp�1�X�^�ʔJ�,N&�xR6��+�Y�J�����T�S$�V]>�9��g!�q�*@�ӖX�ˤڂ!L��}���`x�b;NUY�ah,���M�!�i�����fBK�ҹma��������k+Ǳ͝k4�*ޢx�kX���^K/�'sC�j9[S����=�d+G M��K����AVʸ\����
�\�n{"��.^���:�y%�
��-Ԋ����k��D�r5�K���S.�{�\��d˅�'!�Dh`�v��z��Urx��J"*4B>�p���Ts�^I+$�I&F��d��w3�P�	��#�T�y�|�z�_ʧ��<IUj�2�У����$����NS�s�U-g��a��1�+R���ȹ���;˺X�R��奜+AL#�ĚHW(�I9�-@�Nr��$���y�>d��.(�4q4�����\4���L��z��*H����ר�*���N��
��U�ȢqJ�Vi&�J�Q&E&BWH�@p�N����8E9�"P���Ö\���Qˇ.WId�+�UP�8t�(��%r�Ԉ�P�Ur��;���1j��>���,2�[.�	�/)�:b�2YQ֪K�St��
\3*�B�A6vy��S��T�	�����g�"|?O�}����u�Ez�:�W�p�Oj#V�qS[e.��y=Ox���p_�"��=���*�Ԝ�2F��3�=ਧ�ѳ���#<�,����Z[���*��8���������DT{��W�E9���-Y�BA�L�>��CV���u��cu�k*r4���u67w"���\lc7��V�c=;28m�<��%=���BO��b^ގ����;%xw3���u�8����r��ʸ�%��xwD���ɣ�U�%=���LP�#��$(��گD�q��E�ĉʽ�B���R_�Z�>�)lHኘ�wLp>olQ^��$���+�b�NF�Pw0�I��I4���b"���/.mL�:Cx/h��a�ǔ��	���J�3��ʕ�.D���Y�$��u��`��Ll9i��܏�ʋ:}�ذM��8����D�2\yn�v��)�v�g��`�ˠ����d�jeQT =?1����܏���p@ʎ8|�ǺpJ�r�����oR37w:��vO��U�{�Ȣ e9/��E@�����k�!��*�c+a���E�󭍕��v _��Y2�kԬs(5ᚣg2��/^+:��*Ũsn��W[�{����ݹ���R����8����^3H�7|��cqG�
Z�}�&��u;�Ȓ�Υm*�,Nc�|+��k�Ԁ6�}%^ŬA�̛h�N#�Ҷ5ͼ\��K_e�����U}����{[8�}g��~4:���	�!e+�'�S",S�FZ9g��@Ѫ�F�ّ۵"|`�����7xgF���g���u�sB6$����a�+�����o
�Ey_�W�3��~����"�Hmt��T#צ�<�p��-.!z�M�ŗܢ~�;��~dG|�D����9�w��hQY�M�w��h����X��4zV#�1b�[#3��*>��k�`F���ڈ2#NΕ3�Ƣo�[.�v�p��W�(=+�L������7ڬέ�Q��S��0��"W�L����o����p��|9HKcX`_�]B|���C�;J��B��\E�j[�먻}��ª#3�Ԧ+�<Bf�A�byi�+hlI��X|C�\E���M�7-���n$�6���KS��և���F>���1�%qd�w1ah��z���>�.���QPG��/=�<��r�n�U��]���wh�S�DwXHJr�i]B�&��&���G��%#�]�{�<D1�)9o�-ρ5�9;i쑻M�� b��hp����U��`HPژ���H���E=�ᷨK�:}hI�O�{��uu��z��Cr$�ۄs&J�c�<����A�5Ktn����E���W�_m���ƹ��tyֺ�u���������]-]���"���s�b[&'���C�Nzy�3A�:.��_�����|���wÚ��v�}�bh+�`��e{�8��e�b��q���~�T�21���������`V�ͨsf���Hgf��2$��~k�-���ƌ
��C�k�����t�-Ǿ�[}���E<0���?VY��Ə���w��iE�^(���ڄ`U�a������'�|L�e\��zrסΊ����ĭ�gϻ�&]�R�֮��&�`���pS�<���7a�ͨY{�U��,{�Cl?3�����W�94a��.���s!���gv�s!(��1�Pc�٘���'�`����k��e?r�$gz;W���=�Q�R2�޽]eu�Թ����uyw]�Zh`t``�Mx�ѐ4�p��iu �;뒤��Jz:k��R���=d�c�^�nR��� ��a\����x��q��}F�|6��&Re\�%�v���2_]��N[��Gb��LV/�PYh!������Di��}��!q�u.W^]dzct���N|�%9s��?z�8�YR�ÇP�b�M�S.>�G}��Ⱥf8������w�Ut��mh0g)��ޥ�ƨo�Z�3l�z���<e��)�b热e
��+jԥ��3��v.)�犺��2���Uǳ*�飼�sBY�ƅ�/��K�t�8~*��ѡv3�ı�^|��-ϼ�?N�����������>.����v������v�!�Υ_VN��?�q��
�����,�T�i�����y�ۍ`�yF�Ű����#q��4���c4�ZBT~��VB�;L#]�w�����G��z3H�������
�g��}�u���B�� :��TؒؠŎh�a�5�ʝ>Ǣ���Va���m����*��P��F�u����k6q.��Y��1[���n��x�/�{ΰq9Kvb�mu �Oج�&xPS���ϊ�:���$?�ނd�B������ӿ���n[��7mx��q�&�D�m�E���fk�FE)�?����2󰙇�a�=�n������~���Ÿ�|���՗9m_���O�$�Ҝ�L�0�{�cy֜����=�u0/�]�h���5�z#��!)�j[j�:n���O���K�>O�3�emR�I[ڵ��=�j�3���7�(��Q��>X�r��[������q�٫~[�M�ڍ���εj�)r�j�~c2`=�&�!����v�n�X\Yn|����K�1�M�Y�Uu�_�2����+%X\7��՘t�gQ���l.�ȭ���=��cұi�+�����ʜ��N����}_��kb��mR�j�dz�f� ͇z�;�IB�0�9�3;&�	�B-�uZ���2u��$�8���u��Ѧ��~���難v@z{����=�a�S�§���$08p�ȿD��Q�{�����Gi���~�JF�H*�*�����Z��b�}�v�!�ې@!��,2шE�{]��t�C�걨���9��}�F0��F`[mM���k��1{�ʒ����c�C�lb��e�pc����5�*r�4�騱~�v�g�h�gu7=y�Y6�}�0Mxr�7�t(�3u?
�������@���c��'�5;ڬ�ո~S[e.��{�P�Q�a��?,�l/\&|v�n/�k���(���"}aqL`},W�cT��<V��m�	*��Ňǣ����
*f�;���dp�gO�C���b�Zi��[�=t�x[u��=Ex�=��U��\�M��gQ�5�ש�u{J{�	G���>�מ�9+T�<��(L��n���v�U��}�"��j`�yA��F�3��b�Om�J���ptE�F9�������=Zq�Fu�gK��_�c�>���6$����� ���'�F�P��a���ݯ����ۃ ��7��/�����7���]j�b˓m�֙����/��>�R�F�1��)����1}e�e���+���~����
���X��
�a�Q�e��5�{��q�R��`O�_q���u��0F����yI�D������着����Ke,�/�·f�w[�������o�sTp
�×�����U��Tj�+F�����q��eR�j�`�4cr�r|���;<T���,|R��.^4Agѽ�1R��*�����M�V#��[�N�p��k&C]�ԴpfTq����H;�[�"�{,�/n�Ƿ%��F:v܃º��&)�d}�4:0�pB����;G�;˸�O��#���]�~�ǣ�惄�GX.[�ct|�+W��L��L1Ã���d�K�1��~W69CaU�,�[H~���6�����]7'�})�T:/Ϣƕ�zl�aX�4xa�?A+b �{ݑكB��h7�~��x�
[n�^��pF,����B!�5���GKCw�C�V�'{�۴�ˑ*��lU�rG=/��U���e@8���xvᦳ�ذ�.�Y��݋܎^Y�P\A,+;�t_�8G�6:4�ڌǎ���=o�˳/C����I|���|�/Z��e���eç�-����(p��>aWJ:n!��@��K�#�u�sy�SQp�Rp�d��z#8����3Fx̠��M�J�Tg��v	>[.�y����h. �Z�J�ޥu�;�=N%��s&���7�KFqO#֟-�b{qK��-�aK����-����Ч����v�s6]�}��S�]p*<�<�U���r��~����}�}�j��ؽ��{�g�{���;+��A�L�\h}C�"%x+)��vĸ���:�\�o3��dܹ�d;���.'1f�G;��Dn���r�ch��a��}�IZ��%�Q�K=��^݈Q��E���C���u����{{��
�bG��BJt��u��O{�q)�fUZ�᪀��k�]�z"�P�V���jx�͜��F�6&����rCya��H��Z#���;���$��|��~��=�ʝ?*14<)���	NE׽�Y5�R�7������LC�]���Y��8���ݕ�	~�x�E|&��PW�M�B�F#�������7-�l~��1���P����3�PP�ƈ.r���.��#�rjaFxk���
�a���G�xzʌ�
���&{��j8����q˧�4�+��z��R����xJ��:�}J�Cg�k[n�v�r����ŋ^E��x.�nXSPܷ�F�\'k:A�7ʰv�r�/��F���Wf@�<0k',UtR~�LB+bŵ�u:;�\���j�u\3dv�E��v����=��6y��$&���*7E�Ŷ_�� v/r\�����(od:���?X�P&��I1M�¥)����[����l�CjPi�],������Pɕ��b)��'b}���݈m�C��4�������)t�:���R �J��]�_�� ��	W���g߫f��ȅ5"LW�*��_ԅ8����
ťԂ��xU�z�����<����m��ʔ`�w԰�f���>_1�C�f�'.r�ߠ(?-ZFV��X�?a�^4�ݗ^�B�*����ᘽ�S�ڥ��B�������"^���k�c���zNmC��Jm��,+��	u=�N�����ѧê���H}c�PѬ'a森.�}P�^3'�B�}9x����d�.�Q��ڎbq�į�������.!R
;k��Uwˆj�MM��V^߄p\0>��F+Ր�,�a�}��jF��Pڱ��������Z��>�]�H�$_fdT�Fxy�O��cB�B�lV��6�$D-��S�SbKb�����i�؉�~�j���.�_���W�����8)�\1�Q�u���͜^�qq�{���Q��eׁ,D��yӘ������Z�6�ʱD�l��,,��ϊ�:������������y�s��]���{o���!����k�I��9#�ri��ϲ�K5(~��{⼌]���O���3�"q�͚q�y{^kB�M�:x,��Z<n�L��׿������}F��SW��KP5<��Hg����>j@A�tb�]#�6�²�^�s�ԡ/0�d廝�:<׆��{�j�+��&���X��U��_}*Y�`Ǽ�T(��׃���\��?_s���J؎>���'���q�/J����U$����DA��|)DN�̱:&�dM�1�/em��3�D�0�%5� ڳ>�ˌK%I���cxH[f/U��ٞµp�)8�߃q��qYF�ʍ���>�V������7���C�:��&�l�<�q�-g���"d��7��n`;^�R/า��n�޾���9%�~~�>q�
!��'Z�?��!�8/������[�>��I�%�gw��cG��sq~��:��s���%'[�~j�
�X����,(���*��N�jT)q�n��c2_���=�m�6q��u$7]�ܩ*9��1�D>���ߔF̞=;[zW�"������*aOx�AR�P�Z����nTg�j�M�����l�����2#ffb���gNr\�C%@�U�6���y�W��=ܟ}��g�N�_ǳ�h�&ċ��B�bݑx73WJ�ݞ�̂�������ӳz���"ym�!'*�o�W���aI"���7ϟ�zL��'��J泻i�2IMo/]\Q��x�p�ل���:�a���H�o�ɋu��:-�Y��b'��~�N��ZZL��`��#c�/��D-��M���Wӌq����x�`��M>���>�>����}�(��u���tv>q�%Ʃ�(?�2����ӇԶ�=ݙ�q��Pr�E{qT�ҟu�U��1����t�sԄm�:��'���������>�����ns�m��ٯ�����:����9�tI�}���J�<��'����LP�"���\��,EE]vHS�W��>��^�>��M�b�!�o-�)��I��dz�D�̻��f�	��cޮ���>��1�9P�wjH苀������ßGySqȨ{�h�'/�ǒ�C��~�������f�U���j�r���x�|��/���J��TBɍqC�W���-.���_�d�2	���z-G��Uf<_���~`hk���pe>8z�b}�{����Յ#�ٯ��>�r����nF`yFR�}Y~p4:0�@v��*��S�G���^��=�_����ʨ����M	���\��"}J����&�X�L1Ã��/�t�ݲ˻�-�/��c�ǆ�[B�;��nK���5/��e~�i�a���%��*��tkk���8bx���#��ɩ����������r�}��� �J>z�i�E���A��S1�n�p����=����S����m�f������'�$��{�a+*0\��+۝�`g٨��Mf���iG*Jx7m���).�uN�h�G�f:6�R�_L�8�}�N2��͸yt�λH\��ɯ�'��o�=�ϳ��꼧�������_(���+v����陖a��J�(�Ͱ�����vZ�GKíRG�Kр��ɸ��+��@�}� {����}aZ��Wj=x�K�QU���)fH�d�y��F�S�/��Qw�-�zȔr�'>�1��E9�\1�aZ2�Y����L�Y�{.y���Xi�� CW\ܮ�j�Z/�2����3��{[c*Z�4\����2��0��(~�'�ʝ��0ʥU�[�-�Զ�#h�����k���gb�O�Q\:�m�,��˺&
K���z���ل�'$y8f�9}L�ũ��}׷i�ܮ��rjΐ2E��2�G���;�#�J{̜��LE�l%]�ؽ���B�K:�m͢�&�o5���*���i��v/;�����]ۺ�pK���e��C;��4�D���^�NĨbӻq^�4m�F���ۘ�n�s͑�W;��iDg9�xY��Ve�5g�PS�8d�ǵ�;��9�+<�x6�4Ҵ�Yȅ0�(���K]����۳w�rg{�V��j�yi�����)?U ��ϱ%����ޕ]@6�D��g�)��)�ǝ��LL51���GO.#W0���nھ-9���V�4'G/3�&o-��jޚ��F��7|{Gh3�z|󻯝#��Q�Z�N�ٛ����{�kaۭd�lw_�y{7G���%k�j�p�}V[P�/K�\������#��Y@���3e�SztR����N�����c����o;��T�z&�*�Qgj�G�
��8-���x7I%��d��}3eL�\���r��'.51�����wk��F�>��d�vZך�e^���߶Zc&*戩6Xܜ�C��ex�N�w��r�5!�Lؔ�K>����wý:�4���J�#]�7��*1�bW)��F�͜0Zu+f`һN���>�*����J�������*z]���f�K�!�j����uIF䢒�ҍ�xʑ�Y��;�MءhЮ�+G֘o;skwtE�nnl8���C�o���;�7�Q}�7��V{�C�B�� !1�����>��2k�{�I�ٖ�~�)�A��Y�9�Ò݅��s�ӥ#�!��<Wi�h�R�B�ᤙmeeˆT��yE����AR9���p\�\���U�� �]�|U��f��k�;��Y�uң|��Ϲq��e��Ī��7vU���@̒��0�Q��.�L��٣x�E�J�fa�*K�|�]�7y�LjY���.��z�8+PJ'$�p������VY1*�7�B�q�쒠�y'�&W�I%TS4EJ�FEB�B�IT�heoW8S�$�Q�!&��9GȔW
!�L�[˜ri$Y�\�r���%6�ƒL#+R��Da�M���I&L���t��V�$��t� �J�#�iAWi3�P.Z`�\TH���U(Q(B
T�J�i�V�9p�̩�
qYO"�
�PĸY�A����(�2�.�vV���72H�IV�QO�.�� (�SbE$�5D��C�*ЙC�"����J\��\�RǕ�ڪcHNV,�X��!!��)��̄�NRpI*e\�u����QTU���浦����fHq��%�t�[D�:�G�GJ�s*���X&��D*�!��Ȯω�Ij5B�ZG.iA�"�$� 8��{�H��qw.u����Ό΢Df�b
�k��"�#y&�ޅV&W3oV�$�U4K��3�c��S�8�tUK&G��>�,���^H���h��lT��7�\�fŭZ\�O��,���P�Zj�4����6.f�x7;�p�bD��r��Xv�	q�*��Rx��x��ş*��3e��=O"�:&�Ɵe�umR�"x,=�PVA��Vp�c��c畂۫{#�ܾ�󃾨�N�&ɩ�9Y5'6�5w�o9I�]�gݔ#��	lB�¾��6�,
�(鸇��v˴v��1;,�����@�}�d,�9�;.������Λ����R
���5�Z)�ԮMF�K�t]��/�D����s��S�G)x;�#�=�P
Uj`���-�؄v����$�Qj�ѝ�rP_(w��t��b�yq ��
Nn��@���i�(z�	�;�$$���[J�>�����#qn��1��*���NtZf�X%�@��P���r��9�'-u,�}�3:�rϻ��c�^)*��U�\�IF�z}s���T�:�O���܉���}�}��ߍ�A�s��WTFs��{�~�ݝ5z����O7=�r*�^�$D��[�~)���P��>�b1_E��.�,�>����č��fi�"B=��o����+6�-Юf�LS�hEttՑ`ʏ�w9�ť۝�ڭ���W��};5���D����^���v�o^�%�����A(�;ͫ�����B�Ք��y
)�M��vN���~��Y�h9����������F/,�����?�N��]F{C��y����F`]{��5�LS
�
B}����b&�7s���c�c̿������`�ܼn�Sl��+V`z7�A�yLx�Q>��fɏ����}��R�OxN�sCC�;�A��~�]�/Ъ�~4a��e�3��"Ǹ�7A���彙�t��
ؿ�u�T�5'�4�%�B��u;�nT��m�~�:�0��Br����f�O���eQ��~\|�/���.9�2�� ���E��=s��w.7rn���^<��귧|;#Z��BO���> ��6c��ˇ���Di]Jl����v����󷲯�/���q�t�f���B�i�
r�A����/�]k<�=�n}�"���.��w�c#�;��[�ϓ��.q����YU�bOanN��3C*;�D��mZ�4yi�u�'|�!�
�p��������ʨ��Q	*�<��f���3n�O�w!ǅ��V�����_g��p�ڎ՛�!:9E�*?t�a�[�IB�¥�S�bL��Ā5W�t7R8�,�2�����k�R]�͓�Q�Y{5hS���ܔ4�o1�=�|Z�����06�Ty��>f���+6�%0qs���Q��!hM��ߕ0MԵü�NA���"�[!F�
��W}r�8����������aIEn�k޾��n���X-�� � ��#�n���se�DB�7O�:��6&V{�^��������Ӻ��,p��#�J�-�5��S����
Zhz+!�듲R�q�e��4��&�]�5潦�E0;֠2��T�D�m㞊3Q���$<0c�>0�QR�x\p.w
,��e��/�뼃���<��x��C�	�'�m�='&��f�$d#�fa%�,x]��k���
��xe��ལ���-Ǳ+bcUnx[W�.�zH�94�wo����|��޼}��̾iu
cp*�����ؓ���=OSAJ���\5m���uTTҮ.��s�I+�_+Xx	RV(R���M���M����`h�2�qx,q˹R��z�t�����Κ��j�s%p�{|y�FNZ�/��L��ɺq�����6��5�tY�l?K��s����w�IE��,C��:
U�$O��ہY�W�(S7��`9�"�G\�E�b��ٍ��}�z�ʪ��m>9�n��G�n��,gc��@X��~���-����wL���]����8�ۿp�y��RAW4�*�y�l,�z�cם��=�Mr/7h���{F�w(I�6E.���CO��<>������"ygco�����763��sN��bҨ��ao�d;���F�
鸽�����ϳ����:	�MO�DW�#��^�v�u}���Sdc���Ku�%Ϧ}~
��WV��x}Y���Y�F�:�%j����5����cӯ�����`�T���u�*0y�P)��*�����mm���O��~PL���R&8y�t">��T4mv�}�g'H�DcsNr��l=���_ݟ}���ٶ�%t���a��t���4X�A�l�+=r��Lz٨��{�¼��:�'*�=O��xfyd{�a��P~sR)�xQ`P�*=kr�o˸֕ҬwW^�C܎1,�2�$wD�=̞9�������)e���g��k�Wު��y����L��|��W�wZS'yA�������'��i6���'��U����>����C�+`P����>���m^A�6$����b4&��'�m�;��\M�_��Uv�貭p��ѬT_=��I��!�ٳ��`����ÿ>�dx;�q[��D���o��ǒ�������+�����W���G)��=�=LC��j�goi�h�iˤq��m��;��-�c����rj_t&��PǇK=��� �m�p}�<;��N�e�&�8��?s��}�|�N�/�:�5�z)n�
�GV�-Nz峠(�<���s�Dњ�_{��w��V(ӵ$;���ԭ�R�Yw^%F�D��w��}�}��w<9�z��7����h���@옣���T�)�z~|�	�}��]B87e��N�e�.�Ǘ�:L��F�\��/Dc�l�#0
���Ȧ~��ц��������3ʙ�����ߖ��\ƈ��u�ˇ��V&��|�YJ���3욁cG�9w��||#ض}��pO�.C*�z��c��иey����m�9����T:/���a�z��%�����`=^�o�Oͯ�aL�h��7S�;��QR� �Z\B�����-��n�+{���^�y�����ȼ�K�i�ORT� ����68���z��Ħ��I�+�u�{
�YT��ם9����7��2�>*��'`�R�b� �6s�g1����7ᗾ�.=�&�ɱ7��"�׽����=#�:���t��`�MH|Eto�pL�"+�P�o
�n�gٱ�b��U��p��F\Gy��vAZ������ ��3gO��^� ���!'�a92lA����a��}�<@bv��uԷ�q�*SJc~J��ĉ�!p����_m��P���p��^�u�'-�W-=�%q�1��*�xֳvV_c`M�w��P��Th��\;C�n�竳2�%�M�M���˯2�U���k�q�0���.��f���k�1���D8�\����+��Rne��u�+s�)�Q�<v���g���%�}��_UUu�C󃯊����Z�K�6(�s�Y[	!�b}�V!4Gu�����[J�*:�FX�����~��1=ڨv�Ħo��(P�" ��P�=^�U�9�&r��;�ؚ�1Sww^U�잻��8�����a�r?E�2�ʃ�]eK#����Hrr�ӫ�L���/�d�5c*/G���gu�FbY������\���E�9��y�[��1�٣A�2*�F��=�Ŋͯ*��Ή���PD�J����5����4�)�RQ�NL��*c��q$���ަ&��t=���~b/���1nB�s��tiWw@�2��WI�ȩɼrdE�N+�7׵�.�HՅU	��2���G��u�r�!U�r��Fm��MD�|Sg��L���]p�|�<Zǅ���_�J�?q�!�b�^.���Z�3�����x����YN���^dCO���s���O��i��_dр�S�?_Xp����ԋ��n�A��O/\�S���2�z�uS�\dw=;���r��A\����g�������{OyE���H�l~��ΔT�u�w%�/�Sxla{�����k�`_�4 �R��^�M�(�Ă��J�����37���N!��qd��C��Ԕ�Z�c�Fs)e%���)c�[�W]\�o�X�_�%�RvK�N��6�7���9�o�������������Xu?J�}�@1��X?�6U�9�l�ݖ�{��J	尃���6 #�P7{�au�����/��Xss�M��ϭ���	u=�	�S�,�Q����L	^V F��駼L;����W`�%�)��Ll񦉺W:�{@��q� ��+���)f�����;bp��Q���zQ�=W��c��<9�P���꯳���
���5=�)��	?r�Q���ʾZv΍U��]�����!�ؚ^д����c�Y�q�t�䈅{��M��a����焕�K�I\?n�y��8)�����'�H�9�;;9���2�"GK1��y�K����wd���ٰƆ�T���x�A꬚�6S����ß�������ERYP�קÑ�w�̛�Ԑ�w�G&�p��LA@c����׈�=��}f��X3>�����Q�u�솻���w�����������Ÿ�%lC��^l�j���T�ʫ��7Ɗ���ʮv���J���0���ؒ;�a+��GKF�W�|Va��HL�b�OY=���W�'�дD�����5����821�=��ڶ���}�"|�G*��vX����If�lƨ��Hs� ��v6�ʖ`F���1��k�W�Y�xG?|�/M0�f��� g�vL��350mlY�����N�eU}_}_U?e ���O���Ƃ����)8�ߛ�Dׁ��vQcE�F������Ҽd����ޫu����ܟz��1���&@yQ���]@c�5�&>}�M�^�kj`;^P�s��]�7�1����ojC���>uE�~:�e��n���?��H��}�� ��M�yzd���GVNS�p��>�#o���n:�).y�v��Ŏ?5fX]bz�,s1��,^�ub����!l:�6E�up���\v���=�m�6G��l:^�1{�T������<.�ޠ|ו�y�W/yk��t�p'�lT�O3���bՃ	R���ܨ�5k&ٯ�o��y՛�'w�*��=��V�O	�G)Ϫce�<j:t�ڈǟ:��S[d�Z)��;������������q�'쀑��6��>t�ީ�yg�x��|��9�GMS�]���k��퍫#xo��4�ܰR��Rbe1a�F�-3�G��j8�ټc�������>�c�y��GM��E��n��7Q9�$7��V���$� ��'V�ѫ����g$=�x.M�_�����2�D^�22�A��)��[W��Ui�>��c��80 ݡg�lVv��o)^dw���̻x��#���;N���'�����3�� ��g��# P���o5"KN�!osrX(o������T��꯾����R�<���D�t�oc�W��{���Ja:1��ɳ�U�%=�W5�GmQĳ���~B��.��O�9��G��-�1S�LF���MZ*^�0�V<�$���f��2'�jL�}����
non�g ?t��^��#��s��ʘsJ�AV��k�B��%�Z�)���7����%Q�^���`�8sr�bj9.��Z��R"zTc3������~v_۴\�h���K�a񬎹4�>� =?1�`���r>}�q)���Qs39�U^W�Sx�k�܎�˸6��Nېx
���VE2:�P�^��cՊ���9�e�u��HAR�k�ڹ�"���,.,�~SA�xu��V����=�����o�3�Eb�?o�^bG+��O�x�aJ�c��;�ۓ�r����B��cϢ����7��HOk�o<eu�+��;&�P��"�����b�������1e�7n
����Bƽ��۟wn��ʸ,c�2#�H�.��A�s�!q�lq�^�G��>#V�F@2�wkĈ�����3}�ځ0��d���]@��e֍g�+n�A,�x/`�w�5�V�X��f���b�!�W�Bc�β(�b��"ٓ�/1b޹�XX�)����QP�9�4��k�D4�]�\��̳�"���ݡ������{�~|���ͥz�O�o���9��W�v�g�ShPЬ���ƾ;�����y��ݟ0��=�B۶,�W��ا���N���rԇ�V�
pL�
�	����%���dǺ1�qsK���<ƛ��#̨kA�~���� �L�(4��9��J����^�l{��+ڊ93�q���P�8S�_	W{�^�q���pD�{�@[�0�D-����w�j�����,�۵�{�����+)vb#C�Q����"E�E��3Ċ�(MxwXHJr��um���ϼ3�9�s=�hrk��ɞ�	��@��W�>����9�&r�Z�]�3��|�Y%Љ>-��~
_ٹc�%F��2�MOP�☠��	uU�����a��$�T< �숼�ۿk�,����g�X��Ǆ�&VȒ7� ^]��q8�8�_�҃�!�jAPw|f����L��Z����t�-Ǳ+ƈ.p���ϗ^��#əRQ*=9Y��h�ϊ��=��zOB,,�Y^������g�u�.�J�)�Fem����>#E�4`�=ӳ?�~^-ba1�2���VA�z��������2ˇ�&���y�Y��H�ѧC����]�B��Ym�!�e�m�\3v�Ww�u�W�����'��t!Ubm�v�d�s�Z<��8�h9'�n�g �t�r��d�\��9��f�(u�i¡�7����>�X(w���Ͱ����g,e���,7ڼ ��w�{d�}���g0:���Z����W�^����'H��tL�z{}��s���:5ҟ���˩y>�	�H���[�ha��si��s:��`V�rՓ��/'bwN�G*� �6�VfE����'7Y�+�n���{B�]Ŭ����
r�gZ���U�-�t2h���7�v��R���bB��o�R��F�hf��vR7i�Ѣ���.��MJ��͙]rv�*��q����i^<�I	��R��%"��>��qU��L{nM����e����]4�9:��^حv�T]LǶN6�j�z��(����'��`P�+0��iY�GeT��eZg ��z�]ȹ5Yh�ʞC�+B�|F�0&��?(I0P���`ђ�6�D%Ɣ��[��Z��B����A�0)b�����#	��{�Ҙ���x�?L�����=������M�h��{�{�iQ[HN���.l��w�u�cvn�3=����y ;D��CL?w�/���ъ��
�^I�"�W^��������S*]&��o�*�N�*��[�ery�wk�(�Wr�Wr;}��yc/ ǝ�53�D8f�K�q��jo�3~��w-_V�ֻ9�)ݹ�θ+���9�����ŷ��=�Υ�����)M���?w����iՍv�s�
S^��(�o����UX����cV4��>6�����ǵ�e�j�@���,8�e�MVc��7�Naѩ�*'P!�O�X�p�l�:�����v�̊P���m�_����4��C�<`m3� ���_�7�l5˷�FW.gZ��L3o����p����;E��{+r���˂�K���:ۗx^�05�Q쳽L�W�^���K*���<�r��v���ΰ��`o���:�xy�Ϝ��	��=t-'˧gB������:xi�*�q�O�X��(vʾdx�'_:31:Q���~Ƃw�B�]�`���+���M-n�w1_u��@6���蚾s.�3�Mm��qͣ	Q>���7k�3��E҆c�d���wPxG{Z�\�6X+�%�ټ�yR:kl�F��g��s&�Ec���P�K�(E�Ζٳ[5�:͖
[Ϥ�ybF���t:�h]�������T����<�[��8,�U��vou�j��Ӈ�\�]"�N�����q	�(���/9}|/vN��۹�p���(`(���,V��OyW}��J����7'(˭鳰�nM2�~��[#�h�cE`�:�ܽ�b��ۣ�'')ٸԒ_B��'����=��|��8��P���QY�����Gg*J�*T"��QL��(ͅ�n����av$˲���	�"NQ�S�O!	�N�"Jꪓ)3/�H��D8�f)d�;��dr3ZJ�ƙ�NR}�9�Z�
�p�PMU.uc����ys"��*�#����"�2��i����,�I&��^W�B*f����$�'�\��4��V�t�=N]�-��TP��Ⱥr+�xBfA{�;*�Bt��*&U5�.��̌��f����CE%Y�{w�C�dXI}q�^�P�D����<NT���(�TQhȓ�:����]��=۸x�=I9��B"U����d:�y
�'�
uO��n�	)*F�/��//\���.8sBu�Q�Ҙ\�2���$� ��
�IH",:L�e9�k��\�Y*7!"�*.\Nq�Fb ��#��a�.��=�b>�7���ԭiwN@B��#��B�wӐ]� ����,��t�	n� x���s��~�|�۱���fg�fPͽ�ٞ�OW�5RL@C�C]�W�&r{�A�U7(t�%+bn]F���(��u|�W#�'ՎA�u�~�;a�G���}$q�!�b�����Qr�O0�G�'��d�N��~�f|���	�C9�k�->� m?�^/�ɣ�2�_�y����JKd����������ڑ���*��s�ܨH>�S�\��42�W �Ϗ>x�	�+��|⻮`�^�>�J��|o�6פf|�*���wށ������PYh!��?*�˙Õ��(���^���;uq���!�vϠ�[���%9s��??z�9I�+5C�U"�u��5��s!�aЖ&�O�X`
�M�K�]dI��;?y�WՓ���+�1�u*��*�,_
�Ǻbx��AG��%`��ڤ:~�z�C�~�ؘ�^���OԄ���t,Fw,��9ݝb��b�����q0�jg~bT
�>R/�Y�q�t���U�阰K�<ӛŹ��p2����$���Ŏhɏ�X��m���?�=0xR�C���/�L�G7�Q�4TJ���ʓ.��½�Ʋ�=c0�䩸%'�V����o�̈́�$�N�ɞι���
��n�X_sf=�'Ӗ�6�YؗX�3�"<���%	���W0���J��=i2ȾS�pu:�_�r���}����h�TYI"�͝�͗fv�Db�����jdM��y��Jf�+�Hx`�yk���Vp����"��Wu�)}뼂9�b7ʼ���C�&�D�h���94�q�7�.�E�֫6Ok��*e�H诘�sc�������ལ��������5e�}mE�_�m�ӹq�X��2�7(�b�ҝ�	T�5���8#���ག��]�0��\75�i>�~���v��Wx���po)Q��P򔘁����]�g?]~ߢ�^��G�_���&�h�O�;�{���O�,Nչy�}`�}���\�8��]��k&L>�&�"���\�t�s�c1�Y�����Ze��ʨ�O��!��	N)�����p��Q;u�p�����C̪
_��r�ſ�� -�As�]�Z�8뒕c�~�%'S��5fX]b{|��Eֽ{ճ�.�uܕ��D3�)�u:6E���}9��c����[MM����u'��K�L�;c�;�%c�����Ǳ�Ajf?��0)�C���0��H=/�V�����ZdWll�#�N���^9y͉B��ik����^��w���/���^d^�r���3�(+7�^7$a����b�5��������Z�s�S���]a������I�T�$֗B٥;H�Y9� �O�٭�v�WxjeIӤ�g�6�ӝ�����y�����ۙ9���������q�ɘ��(`XCj�ѵڽ�y�ײ�l���H�~7%`�s��1�dϴnUu���^��{E<'���=1�C`�/���ӳz�<�,�5`���F�(�F^�>;�O�/�G?��0'�r�K���	�&U��P�}]�1��{B����������y�lt7�w6�ȸ����0~�C��JdXEb�}�%=�F+ΫwY:�T0�:j�����Dߜ�}��;%{�������#�ҘN�y��j�,d�c���bY�E�z��0^e�{9�u�L$�ьF�DH�1%��9��>�9lH�T�8l���g��¢b6<�Eũ����+�̉7�bJՆ�NC��M͍�ݜ��:Cy㷞�O�+:���"Og_EG�]��hn�5p�b��HΟQ^ג�����K�Ø��Hq����������щ��e{.�/o{z�K���<�ܵ�/>d��vLQ�y�])� =??��7�N3��]P�*�Ƿ�ٔz���8�9.�SNS�1Ӷ���;ՑO���3<����{<��}�s�$���][z}o1�t�*NN��v_��>��:�,�<k.��s �'S�G������P5s{7�n�ׁS9z������x��W�x}�6_pe�y�X�ݧ[�巣f��X.�r�2t=��y��F\2�������ؕ������{�E�ֈdw�a���WQ.,�~SA�x#�%�D,��L�Y�*yP�/=��q�up4l�W��},9��)+h\5�u�6ܜ�yK�*����_��.1�8~�I�_��� K0#!e�R�wI�����b��n��@o߼��Ƚ��|�+0-i�?o�M<9�vߙRD�]5JTn\q ��4z^ ��ś]β�SZ���r��{)�4T�������8B��J	�-�g<B��\w�
��(a9�:o�.||�d�66����Uo�;��Ӏ'INF|-�R�Р���B�<k�}%���Я^�yw�5��,���=�[���[!c�������&n�1ʂ"VD��*s}츆X�W�\%.��'��0�"�m�'�wfA9���n���݂v׆�B5�k��g�A����[�2:���ĕkKK��)�����[/��@����&���xI�w���/��v(C��-h�<�u�&{�c�C��
u
�U{�W��ԙo�H�lif{(ǣ�1����nE�P[�q�M\������ݢ.�6��u�/.RF�c���Z�f�<�ylQ%Ə`۸ek1��JXdgu�R�J��Bn:B���9X���SK��"S�(�*�r�OkjN��o�����7W���J����������[�k��~�5�i'�����,	w���Z�c�O�HbB�AUT{Wo�FDd�F
'��T���˨1��/Nt�	�����~޼�c.�#�����c�|�9V��U໋y�]b��]مհ��㠪L�%A�_cD8��u'�n���l�߹��^I_�2�=B^��`U�w��A��g~XŸAM9|ݨ6��>�z+g�]���t���=`6�.����k��2Gο���)AMB��>�:��f��x�E��c.�v��̺s�6()�ɗ�4�%�B���]IZc}[�NW�-��u�Uޥduߣ�L폶������O���Ñ4|��� 8R8\�ɼ�Ӣ���_A���J��B�s��=;���<CAn[
�����f}t�����q�b����3*�G��<6v{�@p�z�Ԡ2�q�t�A��+�~(eG�*_��]��lo�Q�{#\_W�'�Y�M����!�n�wR�Y�з��O�UA8D�r]�\�<�Sn����<�v}�Υ��+_b��;�h��Z�D�6��Y�KR�&��U]�6nLS�������|�,сp�+3�K<W{g/uپ�z���:����['��{��W9�H�]ޤ������<����m��hL<t������o�����l;�9�g��@�V� ��`Xy�F��d�/]dI��e��u�u*��oޗ�R���>&s/Ʒ"�`�?�� ���>����j�^���|8�9^�������H-���T�>��^?�ǽ�����V>��p��X5�]G	>�Y
qwOmwq�������3�F0z�uI��/����#U�_ZP�M8)���)��>
2�uٺ�ɩV\%�=�}���k6s����=��Eb��xC�v�D��s�:o&��n'E�,�)�}4�[�kdr8z�<0�*V����Sު1�ͳ�<��g�	��;�hǶ~PU3�+<�{r���t�%ա�1���~��-����?_��[�%LC��YsR��9�I���y�]��@;9�Ly=]*�c1P(8#�� w�lhϟ��3�Ñ�]��S�SdaJ��ѽ��v�yu�G�H��q����G�b��/��,!S�5V�#¥�}�A��˛,t���d[��w�2��.1f*\�H�������L��|��]���L�}�~6Dep�|�fLZ6朩~�oD�HM8����>7A�Vg���ž���A�ydN$��d�fѬF6���n�L&��k��~z�~���D��$^���W���
� |�:��,k��}=�����db��'`�2hWʣ��+)d��V���E�U�|��R���QU��#?z��S��qe��.S���YzzA	W��>���Ӑ6����.�YQ��~��O{��%
�E���~������q�)Is�C���N�՘�w��~��G��j�ݦ';�b�-`� \8;�"\����f@[mM�v6I�t�FF����ظ��WKؼ�䗍�����cOt�L9�x�z]*	R�w[r�^��ta~���7���([~��)���Ԧ>w�׾�)v�8_pY�F�l�5;ڬW�.#�2�5�=gQ��tԶ�T��;�nl�u����.t˫ur�	p�rv<�gP�b�����͔7ˌ�S����<yv;���*��8�����|9`���T���ʰ���з�.W����^��f�g������[�n-�*a��!��2-h�R@鼚���ifqJLn�X}W���IH!N$�'+@�{���W���QN���\�O�혤�v�@��������Q)ޱ	H9�Ш���{U��ϻh��tؐ~��q�TD�I�=�e"p��/�7G52�W�4p�>���D)�}zn���Jo\/�,`�nǇ(�.:��5�y`��*�gvlp��p�GCᕹ$2�=�^�eNcǾW�Ayt��|Mp6OGok'7N�o�ڬɭEw�P6�������9�J�ܻG�����+��\I�SW,0��Bh
�[Wk�='Ho/h�U��hj�֧;š�ٯA�C�v�rqиi�ȝ
�'�G�eJ#(�s!=\nϟ���D���6�Y���=�{����u��'�T�?N��y�� �v�\h}��#�eK��O��J>�y�5�|ǫ$x��%���_��0�����1ާ�8nrU[���FHy��܉X��)�}�05n��zbfL��N������;|�4t�+a���q�(8M�`�o��鱻��}F b�n���V��rS)�)�h��6H[B�;�����ܯ!�g)B��ѵ.����f���X�v8��.��d7�b����1xF?rݏ@�����x���RSkm{���ݛ��f����ݷ���H�t�(�F����㔐8��km�|��u��m����:w���^���*����g`Z��V|1J
� �Ь���M��1f�/s���i����4F<տH��O[��'IO���#�`���xL�{'��ˈ﮺c2.�̶乹1�P�Q�V��(�G�;�ƞ'�`W�[��Cow�jUͬ�lv�M�+���T��<Hh��+�(��A���u�Wp��{�:���.�LbrlC������+y\�x����rh9&��!�:Δ�;u���2*��(��9E�u� ����>��������!����D���xi����qp:Z��������3p�����W�<=T�g[��#V�W��(�]��X�"ȣ���	�]?fA���*J�L��-��b�ǽ��b<�V���ُV��xV�'=�I\��P�F�,:���TD���=�3<HuNt'�b�S����u�J4N��lh1���m�'�1Ħw�[��@��P���9���b(�9t,Vp���S��+T��;��PzPR�������~���.]eK=F&�)@�܌�#f/�z񻮯�5���2�c��q�B�a���!������!B|���7�6L�X�7�����7�#�ɠ׏�#��v{��7�S�Е���\඼Fgˮ�(9�N%��o���g����rl)����l���#��@�b�,�ܼn��J����~��a�z�Z]1�r8W�T�ܧ��RL@CiC]�W�*9?w��;��k�ۗ���YY�Tk��Ն�x�D��3�Fm� ��t�����_@�MC|Gb�y�;�X|����˭�/�q��ҟ>��&)�콲��%][�{���Q۶�9�.�Ko�0�yx����:p��a���Jz�u��ǘ�<�uM|�5hoH��]Jӄ�:+�M��c(�ڐ�;�K�:�-K��L�Ҵ�$�����s��b��;�ﾪ��(2*}龗oj}�Q��6ԿGQ�~{ƣ��HzI� ���M���|pY�L�LWw�3�*��ћ�G����w��A^w�9:��tvF���r�e��f5���� q?ʳ���U�[�(+P�4o��i�2�H�]��>�1X��PW;��Ӹ`��;����|��+���	�,���k�/����;g��u���)7,������U�3�n��P�ʻ���c�����8<ԉ��EC&�x]dI��;'�y^{;*{Z���#�/�������.!��#���a;�@t�j�d@k�������~!�4�屙%)��߾�ϋ����߷_���Md����'��;�E�Yg�^nF�n�������~=;߃�!_�t��J[��A��������ڣS��q4�(��һ�JY]������X!�1�]�ܝ��qq�~��b(�V�6͆4s�2&�m�:o&���uU�y_��^�~����WPr`������m�J���N�]�ͳ��lC�F�	�3��F�8��:��Ƽ�}C:u~������=<�@Vg��6q��1��J��/)���O2)8��k$���Ѧ��3��HF�J��Q����x�a�|S��������̥���r]�����.#Ҟ��U�[ݪ�F�i��␢!Yn��c^p;�d�:�e8�5c� c�Ұ�Hx�9�tG��F�k���h��y��/��C�!C�����K��e�s�;,%rk������5b���g:Í�����A�&��b�a������ �۽o����N�n�4[�F��֣��k,h`t�}]7v+.��3q�I��t�pW�1�b��
�L�����ӹW�v_t�4�\gU��]�؅L�3M��m�<�P�`}�x����u�,�2d�;8��-���<\��u�����m�N��S�IJ5���vl�=�ơ�F�%�����=���
�6.����t�_�a�R��tP���;���Hj9Ô��*����v�t|���TbKϑ#�S���]��n3�Jn�懳�ۈ),Pj��f�7d>]�m�����tĵ���h%�e[Bb�����È���4���dJ��M��f\�wpS[i�u5�.b�6H��SQ5�j�z��*r�p���Y.��Ѿ�|#܏�>��Q͢��)2da���-�	&2�8��Z{nE��>��uƂ＼h;:�#d ⎶������e�C�\�ËD�0g�59{q�^a74����)���66듍�]��)�o I�cf�+u���<��5V��ٟ��EE�-��An���A�#�	��\}��qE̬�U��b��[E����m�/�o&0^s��öf>�+�ٛ��%��	O&'Wn���)*c��9�[.��.ȫ]���yo�g"��w��.�s��I���=���η��swQR�%�K.�����*ś#�otW��c�жZ��I�яq�$
�c�L��O��B��Ô�wHl�GB���lѝ0uq�*b�|^�f6f�k#�OQ�����kh�m�ay4���^KL��S �0��n�����N'2����1�v����S9����*�R��F\M$�o�8 ��P0k�p'���G:/V`ɍ�o:e�h�X�!y�R��;'�d��}��NTck#}��\����k���r櫸�:����M�OoĖ]c�(j;gr-��z�=�'C�������u՛ǭ9��2�a>��?˱&�;�<f3s}f�\h'�@/=�ot��ɐ'�:�r}�wd������Uu�q	�p�f�gL᡻���%HR�uϡݤ!�%��өD��9M��vc%<'+�Wn���dٵ��m��1wD�� WL��)j���r�C�as�T�f=L	�-�w>LZ>�{��>M{���V�T�����R�}˻��@˦)�Su��ny�	�&
\z�sx޹����._�:�=���q:z4�\�x���_&��t<�n�ǞA;(��I8*gRo���<�(.	E�*�#��Y�"��;��ɮ��Ԅ�3"�A� r,�.�^�2���d���r��Q^��w;1Qi�� ��MX\�U�G�s��7 �8PMQ9�e]�
�-wf��rr �+ey�	Sq���AX���gr�S(�9ʡ+�e���8$2��@�E�EC��i:�^mʞ�O��L��]dTU��i"nx�A"�*C��J*�t��)+�M��\( 즕48�T���,��e	�$<�*�d�2�[)$��ur�p��Bg5
��W��z�E*�E�N$Y���a��B�p����P!Y��$p�}��Go�o�!��~�F��g��E��cb
CX��-�M�¡�׾w`�0)�wr�ǁ��;�Gω��%���{���}����O�w߿l��48k?�V�xHȬ�߯���[;����s�5+bF�g����2r����ytV���U	^��x	T�Xа�鋰�I���?W���`�,��D�'�P{ݚ�2C���ϛVa�\fUw��ؤ�Q�)8�߾n5^���:�V�6�x��7��8a���r~��+�ϊsi�sҪܼ}`�!�\dOeth�VR�_!����TY��Xj���1�~ͽ_F8�b����+n`;^�R[�炪.S���!��*�'���N�_f.�۷y���~��1_T�W��؎?vߠ����E���\�%�0�wK�X�1qF���������WY5��C�6C��(t��n�O^U�oݬ�f������i�G��6�fMO/W��m\��tJ��}��VQ1���Y�>h���{�#&^V"����0���ZT�-��+۷}P��[�(�:c����Mx[���DhXC�B�H�]���3��'Ӿ�u}�h�g��,�נk
ka��ܺ�=�����t��x4s�������U���W���0�.T��׎�^���okM��AV�Hh�s�ߝB���q�u��A�)8�v�ǟe��{O��b�.q65]�Z�Wx}@ ca:���y/N_���N�)RZH��r9"|��w���R�M�]Ռ��M�RN�d𛂞�������y��'�e��ܶ!{�O-��$�0'����oT���ʨ���ڕ�6�11ѳ�}�H��4:qaپ�~lw��]b:yo�qxw�`���8�t�E��dU�{g����yʻ�����$� �etI�N^��^�W^�ܞ�.�h����uռ��k�&f3�O����./��\%CP~��I�Q����>��M�A�����lD����6���M�`9�䫫�=Hx�T1y'�C���766�vr������؊>|q(F�6�T�+�������x9Y�\:V:���Oʻ'�G�eJ�9F��{��Q�UgeND�����7�G�֡��_N��b�T\�h����qN�ߺ,���?:�,�>�#�hn���S���:��N��W#_]B<#*4�9.��ܶՂղ܌�]~��D�oTB޹����q��y3]��}�G���[.���{�0�_ü����ˇঃ������؋<����ۭ�>^��m��q\��&Dئ��r�}���Q[B��j/�m�0<�����K�">�6wUm�V����F;S�c|9��' |Š�'l�����?g�5������쁄秣�]����`ӊI,���Ww�K�<�)q��,�i�8ڭ.����>�<K�sq�R'�5�Ǆ؀�ݳ�#@�O����l���o�Yп����+��O}�w2Z�*/�v$t�_F?r��O�ݏ��y�M��Χ�8iwov����|���َ��F���2 ri���t���m� K�����Rw��F��n.�D狸�����.�9����{#1&T���ďw���T�+>�(+ ����Jnr;���dυu�o���](�Q��`���G`
z�Jr���+�0�����Oy�G"b�d���Td��\���$!��b��e7�7>��A���������N�W9�ۃ��I^���O�U.���K����������/!����=��F(��^p{�n}u���4�[G��r{�\�Z���D}a֯5��{k3Ď�;��lLuE�|�����Mz�1$�p1۰�}���8����`���u����������16K�V_wx]<�0�}]�F�6&���o,0~i��;������S��4�;	��vy{YL��%���я/M�Au��1����["N��������(��<\z��)��窢������.k0��"�:�� ZP�����u����%��{��/�	k�4��u�E];Ѫ<��D�lq�����׫��U�I��+bm�|�,�kKz<ߛ�������2�e����f�60>�f�A��������~�c��V+还�q~����a����t<Ÿ�|���Db���#,��p��dݸ�~�{�G�^��}�%�\��#��t��?!�w�g��)�.� gF�mO���WvK������I;�>�U% ��?5�{�Lh�P�c+}�û1u!w�
�8��q�ɨ٥<m��]�A���q
��S0�X6h@�M%|�j�k ���}�ފ5W^UG�<ݘan����mJ���j_�����j7�+�*	h��p�MB���w����'�s�Ϯ1n�c��-�����W����ya�����k�!'�[
��3���L�sY��q���tx��˗�o��H�&U��wK���C�0hE��ui[��K�t�K��	�u����x���k�|Td<�����'IN\��J��c��9�}����"��޸�]d	W�$p��f���k�T2n��?͎�������w�}��շ+f��U�v{�ɂwW�Guo���GΟ�^��3�H�C��OܯOt�(�����]�ц�s(4X�E`��V�l2T�����c��N����h�p{���*7tiWP���L9��%%L��CR�.u�q��T��szq�*gr�+0oU�f;��<�4/��k��ҝҐ�p��У;��$��u�{���-��`�5��$r�JT~����S��X�"��C�v\ծ���%V�P��Uz��7�XF��߀H�V��RBTؒ���S�'�ڣS�z�'�¨�ixNYk�Qcå�.�X7Y�q���ุ�?wk1����!�9ڙ�E�����:0Q[>�ׯǝl�?��M![�
�]_�W�7���޻�#�f#|��eр��H[�-��������}�+��Rc���䘠���ک��0Tw�x����q�nFp�PiPʂ�VIx�(�B=9�s�ZW�:�鱒riI�.�H����;���WFI�oR7��<�LB�9�x�:�|���=��p[�mY���q�*���#�"\�3�4,*q�UZ��3Sr��7ĺ��;��y���o��=V��V��}`�?6ˌ�����Օ,���	ҰN>�&��C����qR��q�__kj`=��E�����U)�:�d==��^S=��*�~Ƣ�I�N�����{��ѡ�t-7p�ϲ⏈ӷ͟5˷\�Πz�? EV�{6L�}���	rB���c�ǯ�SW2S�B��>\hN�n�T;�k]����,�	�Vt���ؤ��>� ��;�}���Pp�*FQ�;�L���)��]�fK�)���̗r୼#�P����uƣ�xܾ㒤�-�'jY����|�ʏj��K��w��0*�X��}d!�� lʍ���}g����f-����.�_|&�}5=��q�`��9;���f�{�~H�vQ�1��1@h��������N�s���#�a�lc���7��i{����,3���;�>o�׭�Dݢ�,!�5"mv���Um�k���_T@�~ѵ�K�*������N�Z���^o���U�_Fx4s�«ծ�8���Q����s
Ք㜻�sܷ��!inB�*����������p���o��{�D�ɭ�}=���죶	Zg�o�W������QZ��)\B���^H����Ė��F�/f�;Aj��X�/?z;�P�E�����®"�:�$צM
����'ԗ�g�כī3��{W�1CX�]b�����������[���~fl�g�ރ����Ho�p��#SW���$���+�^I�#X�r��ڒ;�G�����i7}Q/��y�,_���a��ySePp�W�;����YR�����sEF�R��c�ܜ./�죔?k-�Y���/��~�&��B�L�ߜ0*f��k\��^�}��������1zc K�~"�u+zT��̡29���}#
��Ƌ�'u��`�B#~i�Lv���@�&.�K{�|��̈LǴ�͋�fS V���*}���-�wܬ~�&7����a��}&z�����/� �d�}���R�7������F�����%�VG�:�	�|a���G�Ӈ���r:�.�h�yl�#4F��^S?{3IIy�����{���~@�������;z{*���u��ᨐ�6�}i��|7	���WJY~��r�\�M���W�$L�&�h�1^���<~�a%m�@^e��~��-Һő��0�3UV�LuZ�]Ĝ��P�=e����(�o
�*,v(h9��ZόpV�L����n��f�����	��n,���P�k|ȎM"]�T�F���f��(�#���Z~޶&/%飳؏�ǟ*��3L�_C����/�8D���46D+_Q�iǧ�/�A����w���ѯ��b�z�lti�{��:���O[���)�ϭ�Rϰ_EX]׾���\&���(GhK�@���%X��
�o��Oi�t��BϜ����� ��}�삉�뷉V3�C:~.pD�B�x)V��],��ܺE�#�u@2H��:\�q��9ԯ&&���+��f暒��2�,��˛3 <0�ء�;�]��q��'�F����^�5�Q�_㭩�=��~�/rE���!��#Ճ�ڽR}�O����aZp	���曐��`a(��?���ُ�N��w!y�T���\C� %w1ah���x�U��I��"�Z��r�+늋=���¯�u!3s�tN;��q#��:���]a�'��1Һ��h��z�&�l����X���P��� ��15P�O��a���O�k6r����ؚ�RÞo,0~i�	w��G!�]�
u��^?.�S!�۴�s ���:^��/s/�^�����a���T�3�< �	��$�����������qn��&��WJ
����B��B�`�w��^���<Ÿ��8xՋsY���_[�h���ٝŪ�w���^���)����L}�F�^�Q����ɾNDE��uo�df8^���v�{�������d;��f�>^2��C�@k�*��Ǝ^E�\��j7X��9W���_a�ݝp��~��ˁ�nq3��+/�k&�����>���b�x�#�)��5������a�m{�o��.s6Կ}Fx�qR2�6��u����c$�v�1�b`�2��R�DV2�b��A^w�<3\��?w=;���9�B�i�7�aEt���\��H�*}{���bf�:%W[V:�X��p�g������"����CB��2��;���Ӱٺ��mK�ٜ�[oV�t�M�|�������@�+:U��q:�]]�e�Y2KD�Jf��¬:��;\�F����]"�}�6-�����T�}<�����7�����-Y��[�6\����
Z���e\�1��e�	LҘ��𪮾b�Q�����;/�$K��+�/�~"D�� i�����x�@)u���0��y�=|��Q�ד��P�꜌>������䅺� ���P6��C&�x]dI�$�ÈV�dm+�z�y��w���>�ݱ�Z��Q}�0N��(�`��\����P��jU�5�s�rz�7��95Y��
ue�azڞϔ�ք��E�M��VB��*at����P,z"��Y�����w<yo��=��z|�{���B�� :��HK��A�ј���?^����x�w���`�qb����Q\(:0`p��f�!��5�8����#�Y��T�6ͅO� �7�d���ʟ������-C{fb�W�R�L�eH\Y���~��N�񿯤����و���؇Q��a&bM>6���wWe��pǹx�>��>�3Oì��FFjp_��xS��ڽ���ొ�\�o|=Y����y��B����}�H��T�+ҟ)4�p�*�duW�v�T4\}#Y�tI6h�=��-�Ko���!ki<9-���
⬼g4�7PLd%�Q�R�Q�0d��D�;��/ܘkv��3X����Ӆ�Z���Ε{���EGƥ��A{�͛�#��@S�>o�=yX/l�K�vv+����<������Y����eP�IOw�T��}�g��(�W�|ڳ>�ˌϪ��� t�K��̤�k�~3�ao�*�4�g{(D��@��Ɓ޷�4��Un^>�a��q�=��&��|���U՛�{_X/�1����b�L����.,�>
��O�:�e������雜^�7�gU�]p�K�l��h0������~�AS�]�d8�)Is���1���/��x���n�Ա�X~qc�V`U�7 ,�����kF!���S����.���,c�}fp���D���$k��;�b�ܩ*9�~H���!����,���7"b���\
��̟WIq�o�Y]�v������9Q�5k&ߟ�ɛ�"n>�A_�sQؗ�o�g�&��t��+�|R�\/���}ֈǁո~S[g9u�ԍ��S��@H�"����[��P/�]yp<:J|)�D�Q�:8�9���"ym�!/��0|�X|CtT燥�c��}|]�Z1XR52�2+�$8Be<�/���޳keu��m��Dt��|����>���x�bĊ�M7Dl�uNJ�z��%�y����^px͸Y�xt�J^�e�VQ��E�]�Z'c��Jv.��"����u����<&�1������fe�E1�t���I&�nќF	r���]9y� ��:�ÎU�f9�r;�Ŵ����_]#�[yQ��I��hZ��Hm�ݱ��j�p�a��ucs��u�{�}]-)m�ː����U�p�:i�t�#%�a�r�ۻd��yӯgh�����*[=\�"Y/�[]���$'j}�=�"��ۃ���L�X���Q䛦�r�p�:AYv����-{�G*���Ռ�-�!Dm���z�]��p1�"97b1Z��{�lVX�3^vu��r�e��EJyh�f�֡��^���`9K���(�%�D���Xk��-�z�yK���]WX\��Ɋ�7ۺ
(�㼻6(�3�p���ӏKȜ���P+�V�Y��zW�����g�{���,#؁��z$C��wxfWG<B���y�9�6�rcܛ��-3���u/n��Nc9�. ���Ώu'��ڔ����+����A�5���b��K6�)l�1C��I���S�=�"��b7ٝ:;Hu��
(�!L%eXFO�+��z�Ϙ����Jl��}2�i�}#�Ӻ��,wV`c�����Cњ�����֮�?V�
���v�.�lR@F�˭�w4��;���<o��^����L[C����Fd��Vtл|�������k�f<�>�MR6:Q��;���iI^J5�Ar���W@��w;�h�'OЖ�/J�N�c{��h�s�Ծ.5T��T��%)ǐu�����U;P��nt�s�cz� ���b�]4$�y��/M�c�/|��]T���"�H�ݾ� u|ౢ�r�괟J3gr���7��+^��{Lvj�T�S�h6THR=�}���@�� Q��l7��'x��fyP��o�;�D��rg�� r�6Q�|�0ts�XUѣ�c|)�iW5F��'v�����{���Kn�2}�P1.��zt����ں���n���S3�d���V��<rm'N�<�)���֕��y���,��f��Y
�Z�KO������(��Z�V��ܗ����93���w#Ob���
���]�u��z��Z�T�"]Z�O
N�mjysl�7|�g����e���xHdcק�0�Jw	M̱{�[�+���S��O
-W�=�:�o��x��+8N�<� �h��6T�4剎K�����i�9��EG�{h�%�'S瓉��̿�á�}�����9E.pCfH�����3��76��=�U���?=>��A��'ӽ�.Q�9����j
'���Z}�r� �I����=�)�{"�s��rw�8��f�$��us�V�E���v��ew5n�ma��hW�e�������a)��T�v��ozk�,Y]���u<V�__4O���k	�~�zS��E����/1L�JRE��a$F|A ���;IP���%gH�(�r�.A����QWl��"��H�:$��ZĮ!�I�R�M;"L)��I0����NZ��A9"�����Gga��@�PYP7�iܕ�P2��I`v.U�
bȦHK1�RM9AL�
*�9fr�4*�
"#$�\�<��@\+@ͅ\)V]�d���IԼ�M!SRbs�9p��q����l��Ȟ����(���Ar�� *���((�$�F�QTSN\)+��z�˕;.Q���+���0��@�]�qR*	�o^y�NP��Z��Qפ97&�+�[�!<�!s�B�LJ�	F%� � �V��E�Eh�R�ˑQ\��I-���9�.U�E�l.�2f�s2�UYq8�!>7�"yc����};��x��9��&�y�y����:ܡR�[���v�1e�v�
���;!�ga��J�1����?��l���ee�K)���$��9���\I�A�,K�ގ���yn�G�Uw��!�B��+Y�r)W��������8}���J�<��8����P��: �1K���_>�f���^�Y��9�a�;��H8��p[�bM_�O���x�Xa+��Uܴ,��ha�=���� c��Cx/h��L9���� �������UW����	���T^弫�h������Ǣ�'ad.`���85�}1��<�J���[L� ��<���3�~�/ޘ�)v���jW[[���;?j�L��r7M/���2�ܼ�1�v��k
aE��0���;a
T䍕��ȣ�
���pB>ވg���!�WP�ݸurf��;�k�xc=�x�E��=`�k����~Rf}�P/��A�+�T��)!m���|��Ʋ�Nd�U\ON$��x���}�R�Kp����j,sX,�:*�'&�O��A�����=)P�{.=p�$zz��џ?��q�p	�z�M��ۛ�ݨ�vߙ�|9BD���@AY�'��k��0<��`5��h�~�`��%X�5*�IHt�naŠh��bbf���:3�'n�7��I�"�o����G�=��9v��a����%[�I�=��:ݛ��	V�x��2����B��iX���R������kINP��!*�3�nΧ���4�_�u>�U�1��AF�HF�O�1gʭl���*�����)�'`��·�>�
I����K�����%B�E(p~���Ǎ��#܈ǟ:���z�N|�%9-�R����&��C�ؼ���!z�!.���'��8
�o��O_�=�t��}gej>���_F%w��>��#�\Fy���a��T��V���I��],��ܺ~��UF��yJ��r}�W�ـ�^�s7qd���/墤�!�YiX�D}a֨��TD�����x1ˠ�B*s2u�͸$w�Nx'���Y�����a��Oɝ�`����ٶ��(�ʫ�=��a�Ww`sr��9�&�g#>�wi�5�TÒ���,�2���ʖ�xFt?M_u]��0�=��̮��ޡ.��8���tb�zn2����T�<fŽ�2�D���=[�6l�d����{���@�?]�-@W�
��V�����O�����Ǆ<Ÿ�T>�V�շ4g<4����������;��I�&`��h�G��
�C�\���;?)�و���4�A�)\=��uI�]�9�q�+�(烝{p`bm�
�T5z��sIjPJ�1ѣ�sH��b����Gwގb����)ۨ����z�e�}�$��e%)�:�U��v+�ԥ;�j�9���� ;�kz������#�U��}PW�n�4�7j�)�F`��R�r�+�U$�:�������ʗ�=��iݿ]�>��s�p{�?[wm����~�a��p�gH#�̺s�+,@�Mw���KںG�T��)�u��.`z����#Jرl���o��.;����0�{ƣ�ʑ�dF�OZ�~qz��<�� l�9�f�g1�lm�g�K��3�'c���B@>�Sїf�VM@o�ծ�N�Ats�����K��¶8�6\���-ZF`	2�H�]�온�s��CGb�g���,2�J�&��^���C��6~#�����k��!�} �Q��ok߫;!������˹���
������>U��c`Va>5CF��d�#ƬY;&;阼�Gm�ץ��5�w��d��ˈG�X"aZ��H��OR�����O�&�������!v\��F툍^���M}hI��ҕ�-N�|2CGq4�ty̨l��8�6�����!�4Kr/�g����t��DW�}ԟ��ğ�lPb��17\=?�i�X��z0�ma&��YG��U��ץ��/�����i/�m�K���寽�Z'��Pv�5R�b*��z=�ҁ�0����NQ,o�/��זe�9����VNkb c��}�^	e*�?��<�x{�Cְ���l�gn펩�e�2��沐��������z��j�?�S��q4����!�Q&r���IIqq�ݮ�(�pou��=����~1��N��
��)������[�������+�_�?�މͳ�h�Wt�1�c�lA�>��0Q��.��{��f��n��0P�g�A��z������ƺ"[�HS�Sۛ��1���{+bj˜�ڿ@+��Rc��*�c�1Q�ubɻ���9]�7.׫�"X$K���y��'��!)�nx6��ϭ��0Uw���b\��93�X�$�ūD�IN</3�WI�7��{��^`��Y'��-ϥU�o�\6ը0����Yv��G��J���Uow=Y��k{�/��L�}�M���{�p���jH�[�3nSb:�|<�Jsq�<b6{NfJ�F�:�O�prC��Z����}u}�@��f�㐞ymɚ1��^�[�y���Vܟ1a)"���ݱ��>RF��s�B@�w�8��u�h��g+}�����wm�Q=[�<�<׻�b�ܩ*9�21�Dp�7㘑<�P1P�߉m,��Z�m����+�{������r4�hۋF�9�𞃙�c�{���{�k���U�ԗF�@�A�r��ֱF�WG��_�S ��2�'��٩C�(�m�*�3�j��t{�^�fOr���-�g���jr?CPo]#�vi�����awΎ�P̐�gdo�"�����޸�xbKG�𽝮�q�����ܨ�=�*'�>c}�&�nR&�[ �8AS�ܳ\��>�k�R���sޒ�S�v�1����5��yu}{�=�;�?_�CG&RB�8�<�(.�9��e^�`+��غ�lj���C�+x����܅�U���tT9��D_��f�q��j�b��je1a�E�C^����ַ!���q�k|�����Kd�q��K�8c���iq�]2,-�OM��+�36Ċ���QQ7�_��{��;��W&D��٣���w���
^۷L/Zs;�bJ�/ᓱ�O�7�H���x* wΈp�$��S��S�fq{��T�]�6�����*lH8��p[Cňw�J���O{�bJ��r5���*3�.��偋���+L�t�rx�!��^��=�Ý���t.MD���}Ʋ��fk�ٻ���d����"�Ldhq�M���#�t���^X���ۖ�� �� ��8�z�J^������5�{���K����\ə0���j86��S��>�V���G�$��_�zc�Q�eb�����h�0��b��v8"� ]�u�7�ք{�Cv��ut�G�/��e��+/hG73�:+��$]j+0ʙ6ܦ2NI�r���ժ�����Bǵ+v()�!im�[���w,[�[m4�0Q�S��:#r�y�ӂ���������]���?mCG�C�w!��{�P��+a������*���&����{��i�=�B9X������V�|�JdE�a�hs�q����=$z5eE�A�j�AF�z��ۓ�r����#���E�]W�{Uбh�pC�/Q�̑�#l)Q�
&gs�"��>���^-.!z�M���ano��B!�5�
���ٝ�M��1�:�L�o�]OU^xu��\vb������J��Z�[#v������@T}���*8����~�]�����"$!=@�
$)p�8����� u}Hd���S��T���wܯ|�$��b}K2�{ȃ�L���PC�.¡G
�"X��r���zGiP:�a_h;�Ml��;���)��qJf�A}C��A[`BL`����St���	�]UT+�&��WGE�
ݩ�g�k�G�\j;���cv!�l9;�bJ��&8k :����xT�⼡�KV�U�v-���⤋r��]��#��HOِ7B�C���`m�'�?&v��	�>#.&�����E��J�C>{��z��f�9��Y����D�֝8\��j)���sL�8�<��b
>���_@��/x�y�^nڇKRq#�,�Q�o��ݺ��؄�Q���q6�����Z��	-�&L�3���{j�d��
��={��(�c�)9�Ź�5�9�Od��lMA0䷖!�~���.<�Ǟ��v{.���kok�+j�A\4<!�y��:�5�R��!s��=��1��?`Ǽg�r�.���Q�����c�"wh�eѩ~�S��ъ��A�3��YA�ﳃ�Z6q�wFN-�qqTo�pg޽�j]��3>]{�@����r&(0�"�r#U�pɏ���N���t-qS��dv-X*-� �Vƿ�չxݨw���^����RL@C�G�wCj�}3���OTq��_V0�NdHб_��m���W����a��p�gH�5N}�������ʎf}�\uu�<K��)#�p��H^�S{6�@ j6�W�uD{lm�:�:/Tr��eH~��f	����]p2�>5 �&���ǌi�s�퐴��O����).z87J�p�ݮs|`��X�׫"�)skB�A\�k.6`<�\8��7�Di��߄ȯ{��	o�G�\	��<�����g��}Sᘽ�S�ڥ��01�� �g�M�ן_2����Xb��v#?��{�[�y=��r�^V�*�Dt.��i2�jroq��h�j)���=����w<3��/5]�T<��Y�@U��T�ލ�19�y��ӳ��T2T�9� 8詋�gl����xx_H�K���#���=5���.-�G�l��G=}{v?˚<����\�Y�z�o^a�P?��}Ҝ�&�]2�7��!�@l
��'����k��^�Y|2�����u{K��\2�$䍎��9�3�W���W}v\B-߄L7"# AНk2��bȤK�5ꈀ�Kh�q�|�C��B#w��j{�ք�9E�n�}l9:}�;�\HF�d��C��j������h��LJr/�Q�|8׺[�H�W�}Ԥ�9��A���3�2	%������\]_������U�pS��8�Cң�k!��8׶q{���A�]����+pt	{8$n��UK'i��ì@��Soګ�Q)�,�Hx`��ό� �Sk���%,?ٳF��\"&�fA�ٹn#ݴ!�w���G�����L��>bD�������<.A.�l�W�����ܷ������Q��1n=�lp<g��'���q�/}+Ҟ�4��x�&���=��f��D_*���[a�^g��SA�*�n[Up���q�UW�u��W��ú{��L=��w�r�%�%餝�j���o�Q��2�qyc�-Ͼ�V����\d}���q�x� �i뿻��t��e�8On���m����i�d!Th�ޜ�E�ᅚ\��Q�Ŝ��<��2�p�&�=�m(�*��ާ��.ݼAS��/��ʽ;�np���&|��	�
rd���#�>ݧ4v������WRđ/����������0��7�C��f���O�=�&�"��m�#�j9�n[�3nS�FgMS[pMd߲�+�2=q�Y�S������$08p0�>6�t.��m�e�Y��y%��fB�{>�w��6��:[�;	I������r� �Doܰ�Z1�p{z��R�4�Jt�g�1U�򥗞�3��v��g���y�ܩ*9����!��� w�z��5����As�t���X~�A��t.�f
��F5k&���@#�&���H����xu�<�Q�l�_��RD>���������=�Ќx0b���}���>S��M��u�^Aیe_��1EF;̂�.)���VƩϸ�9ⷈ�?���f�������t���]��@l{�)i�o�2b:R�K�)	�&S��C����u��cu�k��}��=cګ�5w ��Y�১Q�5�ש�m�:��%=��pA��xc��Gr��E�����&�=�M�kF��v�������Q����w��Һ�;䎛ɤF�34(k�Qa���qͽX���u2��j2R����/Oj�	qt��[[Rp�P�Z�Z@}]���F�}*v���
�iwf¬Y'W�e�^>on"]��e�P*k��ci�
U�<��r,p��,n��n��|�4;�pN�N�w����8���s�!�9��o+�?7��Of�1KbA�a�qM�5~�>���*���2vO{��9_?��5�{�L�)�V�˝�0߬6���Sv0ySN:���IZ/�;]�eĸ���0k{=�ޕ��M���]ߌ]�ny�+Ϯ9��J�#���M��U$\�����}��py��������&>/�\���\{�ާ�4I��C���v�μξRH�;��{%�{��	n��?W����?{J}�!R~w�\�	�C���b:ݷˣ�z0ʽa�A����=����~BO^���걈f;��<i�cQ|�9��>�����v7��c��ɓK�\Y'Ԓ��X����i����;͒�QV�7�ے�uy�Q�^19����v�n�Z��Bzs��g�xQU�=Ϛ�s�{�y�;+�Ϧ	�μڏ#m.1c�L		�Ѩ��������Q���,1��B����_�+`��yDvT�9$l���7h���y;�guCٵi��t«���L�T��u,ŧr��k��	*b�c7;	����y�8GM`,Y����W�[�/E6���:=���޺�I_EU6�1���vo�d~�	1�5k�3�>i^Y�e.2�����v��r����ш�HQ�^-晩�m�`�s]m�WPu�aH�*h��e:�Xwz��!<�I<���ð�v��3��שnv_�X�����Z	�˞'	mfƲ�Ǵ���؉�Y�o�ΎT([�G�`^M |�5f�D#��k�x63R�ie�̝�Ja�}�0\�МD��r���x��5k��Q���l٧l���r��]Y������!u� ��D[)�RW\@l$��D�KM:�
lYGj��p����QTb������\��ݴvm:�	���NP�����+m�4[���\*����Y��qR��FJ*�^���٭*���딻}�n������ybʼ��K���|��c��B��\B{F�>�.^�8��,�w|�6 �O3}�H��I>�JR�ܽVy�k`J�Q8X��Z�`5r
[���I���8T5�w�u�G�-v�F^k����	����inT����!rdX��t���1 s}�߈8�/�;��=�)|3�����i~sq+��sSݽ�wU�	����W�¹�6\iُ ���x�vZ�9�7tʱ���Qs��n�������W�����杠��|�A�:H�o������r��G��U��E�<9�(!���<���uڀܮ�Ƭwv'+�#5���v<��Xr/[Y�dҼ|A�I6ɇ��*�2`}�`�W)`�EMSJx	w�W,̭��vU����<ȅ�B�3n�	k�X��;�_Q��Ƙ�ԫI�]}��Ӄ}�5�	��4�<������v�$���8d'��UЕ���]�g�&��]X�;{29���`c787cBL�w�$g�{ΰ�*��(���oWݝġ��QQvG:uN�Uv��b㴩i�۹t�(��qj��r�笭��`�0����60:��<N-@�
vd�ke�\T�YS���9Z2	w�@�Rs�$5g7J��LL�w�b䳧���B�}�gά�3 '
��۔���L��ŕ7��#`;Æ����aKg�)���쾣���58NN�fn��f9����^7NE�54���.ڶy ə��;�r-9�6±�Jgwq����EN�VwP�����uҞ�f�q2�v�?g3��Ǭ�|3�4r��;-�ݓ'Jbi�w��wkq��!�&�e'g�\ж�X��+�vɊws��Z��N�Փ]o�\\��ΥG��˥+����9�Le�LͰ��Z��YB����v��M�W�b��w�,��r`��;#9��PmR��w�*w5/{��Н]�i$9c���z顖v�Q�nJcx�ɻ�x��2?|�?"�$�H$$��U��]2�$������9�(��9W$P��:E�����Q�H�'#J��E0��<��*�CK"{;K�(��y�U�"(�.U�#�ȋ�$��.e��"(�Ez ��e�9�<��PU8BI�"��IEʢ��o)� �(����AQY%f��Ш

�Q�O�J����;/$�r{<��\�.\8A�}'7FQ�Uz3�.W�Vdʸrzdr�W�H�����G(s�9˼uS��$�ETg���|q�wn�!0����E֐�XD\�̸��r�<�y0����v������v��Z��	da���\wr*갼�����8���]g"�5x�'8P\���\�r�ī#+�T��N{�1�(�x���t x��=s��Db#�Ǆ|�E��8��E��p*�������Bl�uȻ)�9.���zC�9�(����3��Ȭu�s�³���(I"��TH�wցW�Q� �A ���+wwpc>�f�>^w�9�]]�J���K�mvbYAȸ\ *V!L�ڱd��x�ӟ�G��gL������X
Dh���aMI���w_ψ�DB��@1��h����%���쟺�!�B<�~�-.p��s�V��bB�|��-x�%1|HT���d��l%D�9���!w{�����Jд����Ew���U�D�,�\�pfr���^����U�_H�şw��bܐM��梀Z��+�)��n�^�=����5к�k.Ϗ`�[{����V�B��q�!fBfh��pd��-t�7%���Ͻ⟉҈��6;[{�y0���}��n��Q�8�E%�^�>܌���e��Ha�	G+���ܩf�˗鬛N��*�٪[�Ww�["��V�זeX9X�H{�)��gn��n؟{������<�Ba�M�6~��3���%�9���7v������d��m����X�jEG�'C�\�X]m��M��6դ�?Og\a��Oo"g�k��~��h<�RS9�@�X\�a���pt
��e��	_��ה�u!�f6}�V�eC���M���ڱ�j��b���5j� pcm)]����MآA4;���w��,!�yٓ��6D6��9R�о��:i�}LnO��L�t����>꾵�ˈ�4p5;���¿���v�;���̴�:��·ujq�J��½�mfʥO~<u��+�-�>�斚Z���=����.��~�^�f����]�jM�V���r+�6�g|��cn�=x�Z��!n��+����V�����D綗��y�����_@�@H{׷z�\��(�ᫌx,�<;n��p��Z�H������\�_G�����x���\=��R�N� _?]�?u�
��oǹޟ�*��q	X����B�<���g���ڴ�����׾���k�q�OZr�����N/g9�pt�ۘ���]��h]D�N��U�.���^�7E&���	`��Dy��T�M��*e��e��=�9�t
g�b�6��~Җ�w۾bO*W�u�Ezl��y�U��<������w�ѕ`mā�����°]��wc�/N�����gr��I��ze��N���q=�qN�3��Xx��f�0�e^�-`�㛕5�t��f�Ȏ���&q�d[$���ëQ��̼�R^� :vЈ�/*��[�c�V Ґ��Cc�د�:{����O�m�4+�۪�a[ӳ[�����o��5�iw�Y�{q#���|�P���Q���Z�G7�����~�x^���I�_R�K������*�9�Vl-�MQ&�,O��A�g���7����&R��j٦�3��%g����&v�1{�f=���5z��b)�{Ѕ�]q���I�������H�W�5׽�:�6�O�_цv��1�KclV�v;Н��4��x��W�ͫ���'���ةq:j2>ھ�}�[ �+������Z���eCU��/��u�����3Ij����JV~H�x>�ϣo���q����GcE�I/"U�S�녎,Mwzf�o/�/-$�겞�-�[�O���B�6���<mLLX;�o�2=5]�)�u�"+�ER�{��1�?"�=cL�;E��u��YE����9��j�#y�X�X�"�T�:��˸�#\����Z~�����b9T5r&�>�@�����n8����}�yr�=˖�i�֓S�A0�3(�]�r�ʽ��T�7����7�
y�N'|{���E�ζ-JN���s�������wf,��51u����:��"��<%ׇ�d�yyuq�1A�g3��3���}��~A�W�yX:��{�W���O[{Rb��4��$���_�u�X��ъ��Th���e[��\�÷�T�;{h����K5N�^ڳK��A �>��]FU�THaUhΩ�m���2;x�X��y�u����y�	c�!`&P]���Y+j���������+nv���f�=�>�����xmzǛaba�͖��x�\Q~�g�EK�ڳ��=�"�O���޶�h��?w�������e��7>��d���f�z�f���.8#�)?
�3s����%�y	 [�r;�{;��	���/={{�z�NV�.�u\������!�[7#�\���=Is1&c==�o�����[E�I"~��c������=��Z��)Y���~����Uv�������4?��I`���ϣ��|�8��a�z=?0ǁ4�~�����5;���2�z���mf�k[â����s��x݁IyM�֖CynM��)���
�Q��Oe�x䝡��Ԝ��-��-f��n�TjS:�[�=�_9��~�{�\ ����d�k1v;�O��㈐[�i�f
֏U�5^�ةfy9�]��=H�ퟗ��Sw���}ozv�_U���$�Oy�Rf��^���qđ}����F��[EY�#��ey�p(�E��]�s^��WW]�xU=ƫP̀�B�{�Z�z�
��U޲;�<}γ���l��{�qVk*��(����#��Z/^4;��F�������imm�#��\e�9�R�?Xݱ����o�n��8�!P�(c{$y����'n��������6�,(.:^1�֌>�6�f�Z�ՂQ#�����ş�ݙo��P&l��y/�cylm/g3�V�Ag�U��^ڈ����{�:}z�*��ډ��T&�q�ߵ�ë�{��!i�/���؏Y̬��}����O��^�ӫ:�8�.%��1�n����k��lM��0��P��d*B6<�OVwtp���W��*��O�⟉ҍz�����u�H?�����?����w��'�zmW�bl]{�;�V���s�Ӑf�B�3`���t>��v�t{��B���4�Ÿ�+���1�{5��ʅ%�.�2��KOo`�rv�B�e��gk1:O�$����YD�����N\��cHaޜģ�?j�����ɗe�[P�>�*���F�n�!�x�
��b�:}���_��ⷛg�-��}��c�c�IC��S�Y�
z��*��r��Ǽذ��s������d��X�d�!�ۼ,������ܸ3Q�6c�?�!�������T��j�I&g��i�s�d�e��T��L�,�b�����}���/E;X���i���)��ds���}'�왝[����Bz���m�[�-4�y���c�#>�0ggoO��Yr��K������Y�v���檄�ݦz�,|�\W]]w����G�ܪ��T�wB��?,�#���*5P�^���%���<������;�	=Gq�ⱔ��M,�-X0m��J��p���P�I��烸��ݠsB�j�[ߕ5�)���w�r���+���)!�L��+����o�̥-�d��y"z�ŗ����ӓ�����F�������XB��jt�������/���]Z����owXl�G���2�Z2�b�V󍥈�3!7TW��1�aG�>��{s��O�'��hr��7��ngdɆ-5��P�ޒs�ؖ=����������w�z�#�������z�F������z�nZ/��͌��S����7� g��ctRl'�W�[��zvϐ[�Q�ZE3��xm�LW�b���������4s3�U�{�(^��r�->����g6�cG5@�����q8:�0�^e�.��CރF4M��2��^��M�g0�i��5�iw�Y�`m��Y����l�2��E߳|���W3»[U���?��}jW����2�����򚼣����-�Cup��1m���#�5���/���m[����/��W���Q�N��vǵy<r0PK�,f���B�yu��k �����5x�q�̋��ޗ�ִL�p˗��PC(Kcn��FQލ�J[����J�V�{2���T{�zoR��V���^W�{Ӷ d��BP��2���{�v,�	~��l��k�	N� ��܎��G��A�2WM�W��v�Z"�u��瀁Uz�*�1�wm�����`�y˞_<��o�V�M��v�J+:��e6)���JJ�=f�C���_�(9��\mvGG�=u��wi��2����n�R�2J�=������ӥ����-�.����Ï�+Y���-����g})�Wۯ_���Dw���y�������٬��,��Mw
" �ꪾ�\F��n��s(��a?w7����"�<�9�[*�G�s�}}��~��3���$k]C��Ȳ'��:���=�Sj��9y.�GWA:�.�C7���;�:h�8�Vu����F�5����וQ�]��C3��x-Jy���"}1z:<#*ߖ�ͤ�6����1������䏁_Y[V;�w�E-_Q�t��؜��6�kU8�S�]{�ҟ"��/�T�J��Y=��Tv*���j�p��o��/~�W���a�#e�����g(X#W�5��%�������~m��Ї���k"�Ś�]�����&7ѝW���˽�gX���0'S�x����f����?�����W3>��c�N�#� 4+�7z�{��?6�����I�L3'k}�4u���x� ����W�'�j�Բ��J���GD~��������nT���H�a�b&c��\�-0���/sy:c�� v��{"���^���Qg����~՗}\3��oB�9yfU�8<�0R~H`�h����2
�Cїs��U���{�^U���*N�����2��Aq�qO���=�n��,�I������y}�vt���Y��3���_fm�lS�K�k®6�]�n�w�	1�,S�E%]-��6���qw:��$g_��u,�{�˂yop�(O�zy����Sw�E�ϣ�[ޝ���-����>��5�[柛B��Z>U�;�"�}�<{͒���[��wDI���޹�ŕ�����B��V?�g����dFv�k�*�;�;q�91k4PU~������i^s����8��@�7��HM[>�O���z�<F��G���1���?]�嶭�"!P�
%���R��y����U�Izp��|�MZ�?}~x�S�Z�*�FC:�q�ɝ��_���k�*	�#WM�,��|�;}R�N�9�=]]�忏��F��A�0�B�$��Ug�d5�MÝˑ���/hH�o��YQ�
N�h0�-�&��h*≯CEX��u��R �.�)Rt\���r|�<"�̴m�7V��TJ����W����!��^�Vd{ch/g3�V���%Q]�z�d����ht����/b?���Cީ�L��L��t�3��ٛ�7����D!��i�!dԌO�x�ǆ�M�!�'���Io~�>=����bt�E^��A���<��$4����ô����:���#T07��=��8^~ERg�������e��?8��A�f�O��~�2�m�"�0R��h���[�I��U]�y�k��hY��/�:k	[�e\�"XY��D���8]o���͎b+�-g����a��u4R�Ȧ�"w3|e�ϖ�W�-�_�Y�z�.�'˵lB��\�G����x�V��y
�x#mXI'�����97�O�C �{�|O��l���;��(h���PK�-<7-'��N��6���o����5�*뭫ޟ �����l0Ǫx=��з֊�߾CEaT�ذ4��:��5�>�yc�f�����fb�b�4S�U���E;V>�wh)� 5/V�@C�u�i�B00���Wю�:7���R�Ӵ�P�ኮ�
�����u�1fBUlv�-�.��@V{^�boU�Jǜ��� �����ȝ�f��6q����ZpU^�Skf��қ�%s2����!g�MM=Gv�/jTe��W�S�5�5�WyDh�R�-w4Ceu������a?*cf_1��j���=��~��|�:'����r��^l�̯h���;��R�E��`�W%U��b�w+��w|ֆ>ΧP��7�S`�ȭ�p���vF�ͮ�U����qe9Y���vq��tU��U�u��.����A�vc⺌5���P��	![�؃���&���S{���#��9���@N�U�J��yRO��oR��͹�Z���C;h�����&�X��_i�Eo|��H�4`Po����{��Wwk�7�Ҧ2c����9V�9__Ez��g.Vo�I��ڧ�+Y|��FN;Z�s�Ǩ}�PgD\��6���կ7dwӶ�[�mΗyg��*Sr�r��퍺�F�ۜ����z���]���8�+���VTz�5�������eq2���t�2m����!���U��v¶�:�S��»�C+6��5b;ѵ6�jN����4�-�ŧ[�!�w
N��\t6Hҙ���Ł{<~�a��-~雞J<��ȳH5GV�5n��a�n����y5:��O%�>�Yuy�k�ۻjܖ�:>�΢5i�,C7K�J�6��;����x�c�0��z��R�丞�:�4���t��ˁd�vEq�����D�#w��X���-�Z�S���÷� �{��hn�<4����-�Ki�]�!+VvlnRZ��}�>;�nD�j�z���^�j��F������7f����Rwbj�4��}�R�k <��ҷ+�V�PS4�{=�>W��6�85��y���� c.�M(�N�u�����t+��H��v�g3��r��ۻ���`{L`t�����oB��u�;��	��5(��=|�6��Y����y���8+x&�:�读�ocX����Y˞yY�W�0֠x�Yځ�_l썂��������G<�M�Y��R�ŷ��z��Z!���L�4/e7C��&�m��f7 ��Ogh�N�(܏Y�>�Mp�O��>���&n���f��@�.�{��/i����S���ѹ�U����s፝����e޾�dӗ6�o�3��+9���^�v���d��N�tI*�Qu�Һ���L�⍚�w4�ЋIR��oc���o�w��j�wv�@��(�Cb�z�JׯU�Y�lL�cf�bX�cpnÙ�^� �%v��|�=�f쮥��5R�l6�;[�-����q��-N�-<�����Jo$U�m�*�=�^�+��rU��G�{�]}|;0Y!@�����@#��"�u� ��*�R��X�*�\��C�u9':T�y<�Ǒl��u0�<dENIQQO��9���)��B��̒(����S�B��%s���'�/V�ӧIQ
��:=ZF ��T�K,���PEEʉ�T���QE��U����U\�"4���J�UTTTA�'�B�yB���r
�r
�U,�Q����� � �\���Nt����ES'Yҫ��wE�ꌫ:AL���*���ZQIB��AQL��ȸ��wq��A}R�QE�R4x���\�*��B,����U#�9�6ʮeA�yo<BT�'=X9�+�*R�U޻��"��#�Vt��]�����.�\T��W5
�Y$�2���	]:p���'2"���K�ۄ���_oQ���O&�*�I�E����aj�������nK	�cR)K�w*;�!�6���"��u����)a��H���������4u��;!񺽸Bh�D=Z�a���؞%"\����_�wn���Y�D�#�༶��}0!�]��z����y��O��;ۤ�j���E�c��'��ʠjU} ­�
�3��'b(�Vz{o��R�B\������f���Z�����6��t���n�6�H�w���ZS\T�?buS�={F���c7���Fjw����<,q��e���Ȫ�{]��V�C0��OL�魺=>�4������3�2!��Q Z	XѪ�������p��7AA̸�<"���+|8P���.�����XULg��~��~ҏ\��w�����%Ί�~W{�p���y6�A��DW������8:�������-��G�=\s�,[y��ޗ��M�߳�V
-��7�^U����ݕ�Q��TO�(K�2�7\��Ǿ��ȯV��?�v�F�c+��JQ�n��A���7ם���^�\��s�$�{ën<n���ɹʆ��|��z��-ޮ����<�E��mZ�x�&^X��ā~��k_�pM[��ێ��U���n	��K�hǷ�.�K!���R�K鰬�<������'���;<��0�����zL��S��J�h�+ː�h>�Y7�>�{q�&@J�!�oz3/����n<w�ɞ���f_�<��r&�~�C��_��E�L~�� 
�
.�1�(����&Qm�D�u�v���[;��Bo�?N�bk��t��u���{���$#mX����b=�߰�����웫v��t�xO����/U�_fe����{o�}��CJ��F�]n�����2B$��h��/����=��U�|%/�<}�aȻ�I��������>��hW21ǳ���W��!rww�V6��T����Y��U,$w7��}Ɗ.�ʺ��7��o����3կ�M��������_1ʾ��X���I�~}��>WW]�*�*'�rb��p�p3��ύ�<9'�Ϻ�!�Z���t�0Q\<6v��Ov%�3�X�v�l=��=��0K������~Z0�f=�#+=>� <65<+6a��\�X���D��\�.�O+�@�Ib,�s��f)b���{�6�� �Ƴ9M\��ֱp�P�Q �Cm$��\����Ư��4���Jk��xi����l�W�l���8U�Oi�:�����e֝��ٛ�e�sz:��'E����N��Z-gQ�c�U�ۖ��q��?/F`���K�K��c��;�+;z��Blw$-2�����%J��[� ��*���l�Rt.�e�����6�ቇm�,'����SZw`��VFf{��f�c���q?`yX�{��I��mk�g �=�1�U�"%e!��j�v�j�X�q��,�*00�
O�E�����D�P2���������y��>��+�b�D+��>�X�2�F
��qO�4���8o!-os.���vۯv���Ͱ��mi$L�;�w�]��_XC�S�]�U5Vw�L�n���P�s]��Ζ�Λv������W�J���Dת�gW�X�p�	��X�;d/9��n΢�`�}ozwR�}����;|ח���:9@�A��;��u�~
���6O�Ϫ�(�Z�o��Ī������Y'��:�G�}���Mȁ��D�����*����_>ѧh������~u����%����?�N���� �N��y�x����rK��]��f�Iֺ�B�IT�!M���9��|�z3���hJ����Q.ܱY�iq����{��mNs�'�o���]kV�몷�l,�����lK�y^�UҖ�����J��3�o�6=��D[ݵ�m�������{�		��]�6��ϕbȬ�N3�o�uk�٧�V���u��ןcO�S��������ʔ���숭S��s⵴a���h_�!KEkƈ��D�y�ʘ���7���oiBt%^�f�m�lm/g2��i��*�����z����2b��˫I`W�5��q��:v��mؽ�t(��m���#�S���df���r�^q�T�*��1�gǳ�׻��$���5�i��X~֡�G�z�k�Ns�4��u���>���S�'J�q���jy���G�RF��<N>��ɇe���l_����2��a��HDQ]6(�}�n�������Y!��dW��5��w6�5����Wfxe��9Czi43�-!K'����=4�5��TNn�.h3L�Ul+�X�f�38���#{��S�G`x1��N���5o�82�l�Z�N��W/%��(t�f�"�����OD���ų�[�h� ^�N�+�Y���34[okq�q}(�T7:��${*�b�	�rG]������b�<�y��0ю��K�4�'������Ï�<+s=�ٞ��0��Ku����B�9Z�m���6��f���a��i�Wg���[s�c.w�Pc���AZ�SX�ۖ��
:�L����I���뼊�ƣ#�W����o�<���{m�Eo�P��1�[/�okn���wq��������m'�{Z���q��8ol��y�L�Wq�d$�2Jo�~��S���J�Qy�,�?v��9`��Z���7����wxCH[��|�ȳ�RO���#E����c��W��]�ǆA�hO�Buo'��~���?�H�E��?MqS��s� r� ����d�ׅ�8�E�ŤB���
,hj���|6����Q���=h<֌(��5/׫_�,����`��N�ю��!��a*�a��3_���_ϟdW��0]�޽qŭc�s��W%��I9�)dj���@����6�d8�9_��Ǐ�)�}�e�{�x*����g<tU�p���G�M�Jj�����X�[�R�bj�����ǽ� ����l�����+Tr�K��d��T�������"*q���'.r���ھ�8?���=�-�dS2ªcM�o9��;"i1F�ϻUE�ھ]�{�<�3����5G��eXv:�Bu5����RW���s�Ͼ-�U۶Gz���?g0���������FM@��}S��βu�����ν^�c�l׫o���a�}h�]�r�f
;Եi�N�̷˽�lώFh쯳[z)��f�Ƕ#XL���xĨvWU3������ݓ�P��@�̽y*�E��萻z�Q����'eyr�7&�\�Y�U�nof�f(�$V��m�'��Fq��h��-^&TM���!���J�#p���M|���t�呶�/k◕�j��J8L���t>5��מ��ie�����G���c}g�|�u�<�6�[�]by.ϻ���xdQ���s�W�:#=�j��V�q�7Ǽ���Ϫ�O]��>���6ί{*�ذj�%ڜlp���MP�I1���ݱ,�:5h=E��գFh�1l�헓/�~�T�q�xx8%�l����z��܅��;��9bܺ���הy9�\���s�#�6��q>4�ah��}����]�geV�EY���\q������1(̀���K�,۽g��Q
��s|q�#}�b�����b�z��`3��7��BF�`u����E�I���Fd��?"�Ȗ,��'v�q��ܟ�H�Z��#�w�4tHA��ugX}�ŃD3=��q������<�����l>nW�ю��!���GD�4��vo�q�я0��>��[���w��&;�/bt��I	N~梂�U��*ǩ	�Ḱ�b��LR9�����*�'��+���	��L�k�K��OV�{�X�U�X�\��0e���)߽`��O1g�������l#�&��c�j����3�V�!�j�΄7O��]Q�����<�N�;7�-a����þ�N�@�^��r#�>wܖF�9e�V
�<����v���55Eo�o]y׍�zU/o^(>��@�֕'z����vr$1���lQl@1�2A^��ɺ���[��&_ c��\�G��OC3���^=��
���yf�r]�t u&�+����a#ü��8�1c�CRf<���J Y��y�W�����5��~fM�5 �G�ެ�B%N��@��_'�����[rG�q
Jq�Z��"��I���!fB�t�v�B��h�)$cK�{'�*���(����)���tS����-��[��z����Ci��v�������Oux����h�m�s������0�~�C�ʞ��=���Q|�9��b���`	VK՞�	�D k�g��#�}r�u��h�7��ey�w��ܚ�||;.k�~��9�R��j�e�V����O>G��|��}������٭��V��뾳�͌}�:6�l,#o��oT�Bh5�Mi�1���.QѾ��~��;OO4�ק�qym���a
�}s[�R�dTO��w-��+Y�r��_H\�+�7���҇��_�b�ӥa��B���B|���9�Dڴ��萆������=����R�/����\����yZ'r�7}�I}I/�ᬬ�'Z���s}�b�
�У3t?����}[����U�#�,l}��Y�
c�L����7��3j})�����27���C�X�H�6XB��ָ	�]�b����Lt��qi�W�-�4֓�.�s��U�>��oYә$-���Xi�8u�bT/cJT�GRɤѹ|l��Bx���Is��QS�N�x�{T-��ʱ�ੌX.��'VΏ�_������[蛷�^Q�j�����Z���4�F]����n���˪�J�@ݘ"�z������B���7�L;�g���c�]��-���t�q����A�A|s"������kiޅ����3﹵���	��c,ʩ�a�W�!�e����0������ؿ�<���X�a�M%͡M� Nˆ4�g��F�����}��=`�P}�Ld��B��+]m�����>��:b(�܉���~����2����!��(%��9��߄+��5"ޞ�{G9�5���<�~�l�x#���������~�1�����^��5��|'�R��:���	}��.�=�+�C�6���P<���_�����B]��p�f���=�򝊧>��]+����07�*@𫴢װ�{q�dvDKuǧ�Ч7\���so^�A�'Y���,��c�EEO�'�o�g���A�3�Q[��n��;xQ�q�}��C���}�cC��E�p�Y�����b�j�r�+��+��"J��Ͽ��`yW��n��+zf�Qt��p�Ĝ4����T��ޞVԢ��k	�h���Y�I��nyr�kMN�
It_9�~Т��U�5z����qg�MqNȿ�����p���ڴ�-L�z�b���V��8��+�������,�l>����W��M�>�S���lL��V�����*堯"g��V�qճ�D�w�%W��~�
KuW\�r8
�i��Rl[a��_Gx[ͯ,�|lp�f�8�p`+^��*��T�������z��c�&�xŎj"��֡l�pGu���N7��]�(�/��}v��g6�l�0�[i�C����O-~�ԙG�^9=�V�VT��CnEW�xPzگV�0�&���cv���ߍU�N��Y͎�z�̻98<�0W?c�FM菔����o�ē��U8ow�곝\�$����%�ȑA?X�C��! �A�8x�r.�^q�ym�e���O�y�H��w��rL0�Ʒ8��
�p���.KP�>8s�j��@xA���ǵ�<5BGF���q��	���.�y�.�lɘ�+턵Z�ٗ%�����
�tUNp^s4�s�N�w��sV�.��z.�&�'un0�Чw��7��n����k�퓙w.�n^�l[U��lVo�ӕc>�B�V�}u��_!E�љfz�W���~ �F{}��ٰbR�����
:�]�3Z�����S��Ud�
�y��?K�.ȑyN��z�ã&����呇��M,��W�I6I��rꏲu����N1�=��hǽݳ)�
-��n8�-6ܥ���T`�E�=6�u]v�\��I�K&`hT����Ώ(�9��qi�v����-�%p�r�	�t��vT��k/WB�v,��hjd8Vᏸ�֘�n�!i/n�4�r�۸X:��R�2b����h}�ʺ�F�mIx����u�9C�-j �D����Bf�mX�;$�N��1� ����P2o��[�鯤���^�| ^���w�度k��������#�v��t���)}ZM�*�*}�O�˾rm-��E/p)��@�E�ME�ζ�	��݇��vM[��~�& ���->Y`^��8���/� B�vtc���۝�|uj��eT��ހ�Ev4��-� 6M�Ir7*H֪�٫q�|��ꕸ���䬱<V�����i���Ga�I��g��u��4ǡ��&g`�Od�eh̷ʅ�Ur�f}*�ct�`|5��ջ�N�y3D���E�m���-���^U��<*��B��L3]�W~�=���b��=��fS���a�sl���	���ʳ�ч4��\+��&C�m\�\�N��9Q]HD�u�qvV��{L>�a�]��<��
b������Oj֨��ǒ쎱�����1���^ {o�X2�T��\���R�Ѻ�4u�g1%���j�z�Z�h�v�+�,�6U��nk�����Wf�Ap^#���)#��/���Ӭ�t�����_9:n-��m�Y[��J�jmqz�R�\^��qeu��n�N�S	Q1��3�g�]�F�o����mF��SjPC�n����^���J�\��%w��fzJ�LI+8@s�{r�l�?�c��9����|x��\h�;S����de�)���e>!j9���Y��5ᨅ\	�S�4�֝�+J��9�����W.)Z�ZT�;: �q�w�����/�0yg�2�խנ+ܽI����ܝ-H�����q�˶Y��/�������������O�����I9��gu�]V(�r{+{:������ѱ {���Ia®tA^���ے�]�̺Je�ɎB:��
��2�7w�ͼ�qe�0�"�R�qy1�@�'[�$���`�we��G_ʗo{o���վ����?� f���� `DV���TL����ZҬ������*H�UE\�����Z�e�ND��(�EUȊ��VJo���E\%B����PQ�d��~,�(��,%�ArL���DQ��9Fg ��*��˕E��J�EEAh�Q�Eʊ��"��2�_I�VG �UQR�s$�"�
H4
"���E^q��2
p����C�ۉ�(�^l��UU�Q̎\���e$�C�Y���E*/Ey�AEUU�'�S=\���/R#Թ�P�dB���Q����QEfE\��(���VEPF�"��Z�[�E�p�B��Zd�i;��:˗�QDDy���}#�|��z��{t�ul���vܕ��	��˭A�`�S͍��VT;�U��5�q;�;g��Q��I�쮔���Z�:�s��~��{��-�麟�Fv5PC�7��w�r�|��q�Pr�Ux�L?7�+�����,��{_%��wg��!��5o6����	�C���v{*�y������=�]��nG>t��gw�ћ�ܻ�O��7���b���}�~���`���}���*�f|w&�/^W^���d�p$>��9\�-���QT�Os}�0u��kwT�����Wa�&���2G�06�߄p�c�H֬u���x<Ut�gV/4��u���F���M�"?���5s�|@��h�jv�Gz/�«��K*+��x��ӑ��y.Q��6[t�������6��J��W��q��W�Jw�]o���{���=]堫���y�N�w��}��ߠ��^�XS��5՞��n���	�;�(X]�7��թ���H�nS�Ⱥݸ��{�}�z�M���l�P�C/OMb]�ڋU�{�%Z�W��\�q}��1Yp�D�7ý��o]v^WTP>����O��]�7|�����e8�Э�kp�ª9��)�p�ɰU�׮����b�n�Ywu�dq&v��k=�(h_�����T.�˳���^�6�8�k���DA4�%��]�h!���x�3/�u��YX�>��;�m
�>��g&+�fΔǳ5f�^ =�
�N�Mz,�,e�VTOοC(��;K��>0�^�7���fw8���;�x�5�ZT��ߝg�u�vr���x8����L<���X�.h@Ʉ(n-��[o!Sd6�4�1�������0���Y=��z_���2u��ބ+�M�igKi�S��u�-gn�;�>�f=��{{ggԠ�v�8z���hu���Ge�gQ|�{z7~�;k�kզ���wN��;au�F����'���u���^Z+ϊ�eGl�.��'�|�L���,�v���{�����.�2*�#��f����Vd��92}ro�������^�乡����VX޸$X�x�"�<6*�;LyE٦\�^e�w.�û-��[!��\�@O��!��8�k�9u׵����9�5���,5	��FdW�f�֨K�o�=�8��ox~@�#ua�-`܂�h�5�lc�ɺ���a�\#�I%�~^���/�-
v��3��@��c�q����&���|��͖GΞj�~�9w�ڷ�r�Y�d��D��Xg�j�?�?P=���=���\��q�����yy�Sq��E�b7���&}ں��)X�4(Ѭ�_�ٶ������	Z�AyU�3�U�MNb����:�U����侘!���x���k;�W���3�Gܧ�e��^{��3g�>hX	(���ٹ��aN����g���>�K�Wd�ת+���}��o��J<��P]�74������lJ�f��<\��>>ͻ�^9������&�zojos�/�v->1�/-�g:��^nI�~�S>�T�I���<h*v��{|�{U����djܵ��ϺPǴ.�֎��_+?� _��8��^CůZ�l_g���ϬG0�KIkGfaIp��F�]A�ޚ��K�ى�43�[�4�K��5;Y�Y���jȟC3�ÇW�L7"'�vI��b}\O%��l�,���^�k2�s�+�`VQ8X^��Gk���ǖ��M%:*���B9�bԵ%���w��iB
�ޣ|M�Y}�Kyd9���G�*`xT�nv�s��pC�?z<*�^H��M]�p��ëv?��{��=�q�]�$ jZzt�C��fm���Ѱ�����+n�z�W��h��:m��۽ǽ
6�a���{Q=�\��t��z�f�^��c���~sAcڽ��i[�k��ϣ��N�?<���钰�֙~�����_ok�Rj��)KwVug�Hs����D$9�/meV[:<3�6\	����?W[��W�a���#MxN4+��]ڡW��Oa���o��:��<��ä1��϶����qeS�����A�*7�ښ�V���K�?=���WX6�᱆8v���}p:�ٺ�]��Ɵc�w6�����-J{�h�q��w�X=V���d�������s�ּ6�{?:!&�a��}�oў��Q 1*����wZ=Qm����n�mr�^�1=ɾO��A�xє��1~���#S&�6�&�7�J,$�pjJ6s~3�>�]P>)��z����-`�x5��z�f�V7.��WY�U*
<�8Y|B �or*�!RDn�u�WN�$�N�����gM���n;�A2�v��TWP�_^��e�S鏸��~3��x�����g��+w�<�
'���wެ���,�
�?6�������fn��I��[ن׌e�!���֩�� �V���?�F��A>��vQ���z��쪤�]���̻"�<���;5�ӏt�`@r�e���L���[���ڶi����̿�A3������Qp� ��0v�;�s��Ƅ<qX��?�I'o�l���y����B7�{�-�T�n#r����U
��~n��9��[o �|�夵���#ޛ�s�8zE�o�^�Y���Db��НW��w�{������C��<��˾ڋ���	�em����q��@�;�{;O��Y�#���՞m��u����x����P���h��o���t>j�W�r�>�/��޳�Z(�^3��&��EsU��r}���G=���"G�i�#�B�Cq���򹊦�Tu�R��a返�T�q�U���C�\���;���8��=�&f�R0&~����)��ש�[��k	�#sc|��+9���6����'PJ��ca��tł�e�2����A_�����]�]/��Ir�7/h5l�+f����Y�۶�sT�S9k��zM�O=���̩��}���lK�w���i�\��k��������r���6_��{o�D>��2��&�ީ@���x��-tߏz�otkؙjп�	��xZ�9���x��Z���w ���t:ᛟM�3��y����Bo�!i�o�(;�ƺ�N���ӆV5�re��
�+.�Ϯω�/_�aO'���"/�O��F8^����
ֵ�~q#��'3?�;U������.��i�s5��Oj������ퟂk�.4j�X�a�	N����
Sy~����+�u��93^}q�<!&���U�%vz��3_Y���@��Ƅ��vF��z�8O�����M����w����c�c�"����kER��ՙ��݇��X�A��B��U��vA���vis����jY6ld&��nٓk.U��c��.W��{�s��Pk������bDRr)�҂lᙿV����+�2�]��wx��UÑ�����eL�Ҋ���W�g�x��6�+<8���"=��ԼQ��
=��uf���t�|�s�s�^�FZ�*��e߇�B����T���5�m�&L�\�V.v$��I��(�Wr�t�l}׊����
@�/�oY��_<j׍�u��TE�ۼ�.��_��Ue�o��ޗn�N�=����N��̋��Tf�O��n\K㓽�2O���Ď�̌}Έgua�q�#}��onb�0���m��k���lm�~�o�t�v�h��]6���t^惙�����j���ū�BÉC6�{`P!糹/5�mb]X��Ɇ�=�V;SށM�kh�¹?^�K������_���Y�Xk=��|�JЪ�~�2�8a�>U���/ݞ�e�@w��ג���)���4��"�3�X?L��{��������_ܛ�/�J`�(p��va����u;.�l���߼�}�{����5*��]�/4����6뻫.�h 8~=u����; ,5g��RU�b���o7Q��Ch���<�C�)'��L������)�1�x���-�l(e���yv�W2I�em8��t���9�Y�(Y��BC"��[�:�R�%uǊրn�8���>�b�^Jŏ*�^Z5oEO�j�����DZ�{�Wxj��Q�ڛ�L;,�O�3��2̯.œ~�щW}�_Y/���,(j����l�^��a��m�������M��[U�r~}7�pf�z=�m�w�9�e/[�M����|9����܊�5�ȉ�\�����+���f�,bE~����Sv;!
�䎖�JшMR��^�}ћٶs�RD-�`$�2GGX�2��$ hKOv�0]]ms��}=v����|����O*I�2��#��8ݾ��B���y�.+�5�J�g%p.�<���^s_,{W��+[i ��[W5��d��f�U�5.�u�{�{x�� >�U$~���������M��mc�c������^�W{�u��=!�bu"��m޳]n����s|Bi�F�'q٩S�3�nv�9[���B,r�j��lo�}Ő=�)[���Rh�v1�Eה葮>ǟ;��w�N'8oP}�jkQ����ˣQ-�2�Y���������N��|5�u�Y(�mMpqws1;��-�DRF�c-	1��Mfwd�������;�N֝�k��7��N��z�Ӏ8�Q/��]�$�}=I�/}�!��y ۼ(XĈ����o��pPS*'����W����3�џ�<�~����m�]kF+�"F�O߇u���Ǣ�jL���S辣��z����ct@I�`á��"��i�VXܻ�W�x��2�+����8r�6��}��+��17ܛ?'�X�Q��$u_�?m��f���w{ǧ���1D��}}ޓﹶ0��j���^p ��uYFⷆ.�9��^,0��Cå��S���u�*WC3�Q[6˂H�̜쥾�[�Ю��ʷ�??t�QW���"��Ŵ/�_�X{�������B^޼�P|9�9[d6��j֓�k�vE��("��5h������J����^?��B��_ѭ�Җ�� 6��Y90�~�����z9=��]x�����]���>�[�ގ���9�Q��.|R���=^/cj�f����uPz��R�*�PI=�y_� �g��#H����m�3�}Ȩ��;E�]$����.�S���pX處,�{
�k�[�\����5�YfԾ��nS2�5$�Q͵iRikY��<��i�W�H|rOV����t����Lc��JH��?|�z��̳*D<�~O�v~�_<��ȸ�ɭ]UҖO]�����_ϣ�@�W҆����:������/J�:�c1)�勗� 2l��]������E�cz����W�o����M�䨆<�,^^ػa�/HJ�TB.�#���m!�5�0I��s<.Y��r������>Q��9wK�-���]�o�[2���5�Wc��V(���ܼ#���<����^k�
v�������D:�U�M�2#��/ۆ,dwO�kٸ=m7�;��&~up�a.������Ƕ���I��wFyi�W�Q���c
���y�����M�$����u�6^��ٖ(/{���٧�%X�0V�Ʋ����^@:�֫^F���y��Ph{8.V�����u��#���������?�����^�~)��6����l�����~��X�1���=���d��� #�0#���`O�����86!�Bm���dv�m�;���m�D�m��6�C��țm�8�l�m�D6�"  �6�'����m�Gm���؄6�#��Ȇ�dv�l���"m��wm�!��m�Gm���dv�l�m�D l���"m�`���m���d@ ��dv�l�m�D�m��țm�!�ۣ��m���dM����D6�#��dCm�&�l�m�D��\X2&��� ���C�O�m�}ɰ`�Dc�����?�������������?���?���o�Ѵ?��~���>�������dq��>�cm�>���~���?Pm����=�lm��&�O��7ٍ����q�����Shm����������?����罿����I��`q���߆�;��c�!��v��`� "�gm�l x&m�0!�m�l`��`�6 <��#��ߏ�?��1�P�P�\c?f>F�w��|?�y��ߑ�����鍱�6ߎ�6�y������o�|O�����}���lm���>[����|Pm���clm�I����i����}���8 �cm�d���������7��ǳ��_��x}����n7��m��6ߑ�>�_��clm�/[�R�����}���;��ߛ��y�v�6���~s���6���~�|����(}������q�|߯��,|����������6޲�!�ߜo�q�����7��}��>^��Clm����oE�}7���cm?���{���o���o���d�Mf����Af�A@��̟\��`z(2�6؊�F��J���%a�
BU	)@�J�T

l�l(��@�lԂ�@b�M

h�k@	��ZM4�em6ضŬ�J��/]֍��jV��c%��%��[ZK[5%[hkKb��R�Z�CLM��(P�jhP�"Ԋ�*�=�����V��R�Q�P��&Պ�«"֢Uklj�ME�֕�V��m��m�6���մYkMlH͍5k3e��U��CF�kf����LTM��  n�t��j�f�24��+�M�U45}��[�Tjl[v�.�Q4^��[n�0�5Y5M����r����6�%B�T��[mlR4�+R5dm�cv�  ��
(��CC}�\= � P 4�ۇ�B�
(P���n �СB�
��{�9DtYT�K�\u�� *j�AR��ұMhR��[}t��Z
�t͙���j���V��>   �*��[l�ݥ(R�[l<ٶ%����T֫6�cY���5�Z�Ҷҧ�yyq탪iV���C��m��=�٭[5*X,:kM+]���[w�Z�e����  s������������Fi���SVQ5/��iV���R�-�{=�҅V7����V�uݭ�f�s�`ј��T��i�i˭
핵5UV��  �U 	�QTQB�������l ��gw
�:+3 (Q����Gp �e
Ѳ�á�]m�b�&�ٓ1M-�� ׃E
��(!�, �[7�h�� LY�� kU PZ�AU5whGUk�@i͚ʥ6��`KC�� �
��pP�um�@P]V
�h�T�����`�5LSM�;� �+�4km����)U�'���&�kiU�#6�-�� ���餕�z�Q*�[���Qm�+�w($�+�{�� u��mq��7R�(*�z�<IQK���QTA���RIS9z�j(�ҕM�����  	����u}Ǘmډ]��zPT�I�[�R�U�7)ܪl��㽼�F�f�R�*@����$�+\N�������Jvp�y4V6ڑ��0�3�  �}�MT[�����Q���zDD)c�ooeͩ
����"��/sC�)lח�oJQIQ^8�Rb�.q�8 �v�8z$)T����R� �a "�)IR�h0�O��T��  ���)J0  SzhUJ@ hi"LʩM  ��������?&�nl���?m���r�ܞ�O��9�����<�[�%o�翚y��$�{�}y�p	O�	$$?� BI��	O�@�!$B$���ϻ�gO����j@Y��k����v�i�]ep�j�Vsww����8���:d��;�!MZ/ �v#�2`¦����C̜V�]��s���a)
ҥ��t�r�����^o[�7q�{sWgeX���mÏ�6��n�N%�ۨbɻ�&V-�{u�5Yi��{�bl�M����z2�ͼ���[�^�D]�?�u�nӷk[f����pBv�H5��.�=Պ�u߶�&�JΖ��7j<ӢK�!/�4�Fk�{U�0�j����9���Y�'�p��ҭ���@�78��1�*^��
�C��e���m���܌-����b�,��C����;B-�`��"ca�ٍ�v:ά����^A�$�R΢>�5��3۽��s��1t��5���9SQdu[D�^�N���f�sEe�4f�sI�J��4��րA�nV2x� ���iWs{
���f̤,`l�*CN�ӤI83�(JI��EqL��u��]�����ݥd�4]�rF)��g\�YT�r�"qYz�Vr�o�E��U���6{r��U��}��q����%��9in,%+��:=�7��������8an�{O=m��A�F��ׂ��eЉ{{S�`�#��&�L�<�������������5�ە�)HԄ�-�Kjכ/tWGm�8=ހ�mF�t����W>	��.�( �)n7C2��8��Ή����#��v-�ss�k7�w��c�1nRBK�jn^q꼽X�"F�c�:ff���]����D2V8/3S���@eW8^-���gw+Ρ���`�&��ՙ|�� ��� ��j�Z	�"�-�	�[��O�з��t����;Wz��z�W�,�/RͶV�1����ԖF�s�3Z��K�.rL���Wt�
}����7�{M ����cs������q�"7]��٢��w1j��}����6���w�g;D=cy��'jV��glv%���HY�z��v�Q������<P�t��i� #�Q���e�pQ�a�Nc�K����c'N�kv�$9voϰc��N���-]Y�U��]Goc+q�����q�7�1��f�j�|#�Z���/��w�Q�ۅ)�q��Ҏ:�	x��B���Ra@U��1f�oƷZ�����t��������.륲�k�{��!X�-+�����8un��W�w�b[�z�ۍ��{���8�T���ž�85:a|T�+m��^��"�xo7��Mv�-W�착A�a[���GS��f�Lz쏢f��$��`�[p�����ނ$ة�-��:6�7Aކ�T"�-F�L��(��(i:V�֜ev�括�����k=F���QA"���X��w�Y��(����vC�k:���,#g���Fb�vW#n�j����֝��@���<�	t4)�Dn�[��}�rdUM�
����Qs'�u�V�������j���nj�7gu<J1oxWH�Z[v���|�+X��x�u�jю�X�<�^(�<�;����7A��-���ƻy��t,uc�xk̾`:�Z�j|��H4�f�^:��d�"�J��ݮ�Y:�u�>���Wܧ<����vkPֵ�7-��� �+���U����o<l�>v٦���9g!T�S�`�x�yԙV���<C�`y,n���FxmA����� ��ځ$�(���_I�^�!�ve�,ν��ig�1=%������v��,����"B�Y:�m��|�HgX�pF�ag��a�aov>��\	x��۹�3\a��rV8� U<��7�`#�HG
	�BΗ�[J�[/�b�6�2�P[��"s�G�ִ�)�̡����i3�|;�+i�x��z��nvi�8٥���@ۧb�о�v����bɼ��K�-�(��	oQ�F�mVi�L�tX`jRnkC���@�ި
 T�	�ž���Ziy��Iv ŷv͓%�A^\S��
#^ˆڜ�,�紉�C��1��.i�u��.0=+z�Y��a�7�<5�7Z�[�]-g���-��um�"Ck����� ���8�4Q=�w��A��"{2�<����ݷY���l��Lc��w6�5M^���a��� ƻ�=�ƭQ)n���9�{.v�@�qȣ׼��X%҇3�%vip��tO�v-Z62`T��cvv��x��Ud��W�	�z��y��NL��ק�̰�bIV�ʳ�gi�t�7��s4LCN�2_\�+;nӒm<��2w>�w6�B�9�p0�Ŏ���U�֙U�y\y0�"Vm�NƧv����@�!��>Y��Ȑ�ˠ�^���Zo/��(R}]�Z�FHS��t6&.Ѹ�۵�hZ�=S�&��|�e=�u����wU�_]�!�i���C�<7�ie�-�iR�a��k�ͭ�zu���ʴ�4oU���G-o+LkI��)����l>����»�Ã�q�+��~����b�"3Z}7v�z*�V�Ry8����椉�������}�u��T�S�����@S#�Ů'��\�����T�%6)�	(2�Y���nX��وfvSH��D���]w�x�Dp�U��0hU#��a]�������b��`��2���э���vh��$ۊ���$��z��`�ۺ]�V����� j膷���[a]v��VXv�m�u�Ʈ�h%�������O��n
�Ʊ��o�%�a-<7@$xn:��wh��s��gRZz���`�u��e�Mu�t_fCcKoSX¸���1�7$�,z�� y��^G�W����K�G���BL�F������ޢ+0���8�+N/�C׋�h�����-krtbΓY.�E���܆F8,������wٌ;pk�'��u��Y���!	N�g"moW۔�L5(�e�=�����y7���tb���ζv�����˻t�e�ee-jC\�q�.�����^�h��0�fvW�F+,rڱc��w=�ބ�����x���Uu�t3�MFd!B�	Z	q�����
�k�jse.&��i��sO�����0P㱬<������s[�T�8n��h��Vӿ���A76��5�S�%��*���x��� �8��%M����hG&��څ�ɓ��ܻ�ND�\0�k@��&�1�,k�ϭeX���7��u4��4�a�CF�:���wٺ�O��0
X�D	�-)2����!�u��Ӕ��m&P�� 49�'wK����h�u�ڻ6�.Χ�uՏ+��q3Zn�Y�b�bL<=u���W�뢱.��Y�V�&��I�;8�ݭU���*���������NC�t��n�ʗ|�rR�8�1�Z� F���B��<;(�3#�a�+b��q��ַq� �S/z��-��W#��x{��@���o8�#R�gU��+���]�j�򁺴��~���ª��i��b�Z(�n�u� zPr�U:��6�&�)ko�&-*��t�y�U2q���Ѷ,���e�RŵZu��Phc��^��DK�M}��np��p4\����������s@Z;�����bw��7��cE���g1^N�Ҝ��G'%���S#Py���څ����L�nWBR�n�ՅUէ��aޞ�F�6i�X��v�+53Dݠ��j}ٳ$ː��)�9wU�����m�u���c-����O6��f�ptf��޷�Qm�E/h0)(͹I�sZ� Nm��,-uLc�T�N��i�L!�Xi����'G2�̲��jн������{�Z[q������t՝���.B�
�r	�Wf��W�,:�4�œ������M��=J�ۼ��|����jD�V�>/��狒J�,T.��\��^���U[N��4���5�ɚ���5��cq�q���5C��5�N	<�� �y<�^:
sf����0e_rmiüQ7F�<��ӎG��*�u�-�]������5�%O�ܱ�Ywj�|~�@� �hvҷ�I6{@�1bee�j�.�lސa;9.;�.�40e��5�C��>˃S p3{��׷���t�0݂�F%x p��.����E�-뺲nblQ:	Q	����b�7I�>��i �`$�sj���l��� �oO԰pg.m�h{��I���I2���ǽ1���Y��@��u=+*���A�}K8�V0
Y�5��+IF�ɓ�^�1	��^��vL�/"٤ٰ���=��[�]��z�%Dao���v�n�uio[������VC�a�2:[K�w<��߬$��vv҆�-� �[�\7 \�%�Z��؇f]ӯ��������^h9��V`O3�������N�&�RwxwC�����,�tn��*���u�ֱ"���31�,�I����(ef^S�h�g��&O���)g'h�%f�هA�qh|��M���;ywJ��[��f�Ý��N�R:j��^�Xi�Ŕn�F��1:ã�(4�sdwB�KD��M��XW��)Q�������k���[jt4��BţrukwSOGL'w�t���=+{c-��;�����M��ɛ���;R��uX�F�sGn{8��R�dǱ�8��yU�w��hin�3�L��"��R�i/Yz�7l<�=�A�b��ux�=�[���c�Yz2�3��uj��n�� �4E:��rS��*�y�[喷��5A{�Be��0�ҳ�G}��E��O,ǥ��*��͌@8ijk.�ݘ��x��4#��"���o\w��,u!-�-7��W$�.�}*EU���]���Y�帰���e��L��י�|����W�c�\&�6�1�gV.���[3lYz2s<[˔F�3�u��T�
���5�Z�����N�s�^>�f8��)P*w��2L�����s/�j��%�hx]�I����vD�cS��x]�^ƞE,u����/4�,�">�z(M�Kh�@�n��Ϋ<&v���n�H�j��cf*o$�]WWf+��P���GY�ji^��&��!�6�83����ĝ6kQ�+�i%u�Y%v���-�����[�����VS{B���x��ܑ��IWcoi[vM�#3/,���0���s��ת�@p��OI����uYoNoe9�ks��9e��0��rYs��<X�Gز�k��E��3�2m�o�e�C���Ӡ��Wgjsb���v�t�^m�w5�Zc�\ $�R��9�� ,��tK�+3�x��{羗Ry}vR�v�wW��o�:T�q��#�$��D��:̥�5B�ݒ]�6a��la=8�a�\].^�(R�2����7��H�^ؘU)�Jې\�uE��N���B���yA������6멽��n<������P��$0 G>�oA�L����ԧdO�xجp/��r����&o,�uÚ�O�ꢛ�v,��Z9�ۃ��Ԉ��UU�+��.y�ˠ)9t�@}]�*b�]�i��9$>72����t	EX�R�Wgr���GWWY]�X��㵬O��fN���s�Qg���2���%<�)p�{�XP��)���G,�DE��v����p��{�x�<Eqy���KY��i��E�dLJ��Wt�Zy����C�9Ճ$��K����n������ɧ~�3V@�c#@<I��ԉ�x�V1o=(k,Κx8�F��x�;pY]bcP�q�ǥqAѧƓg���掭T�ئI��V)ZE�l����Ql�ݫ�b������NQz��+!;V�\�T��옗ew7��T�כ�o����"�S�1�O�i"�e��i`�P,��6A�A��6���M�6�z��e�}V�ň�sa�V'_ȣ�^C/��h>�w9��.�o��c�?gIYǬ���� ��[�$�׿�k.�&rD7L�}�Q3]�^pdp�����L��-�+/��&�n��E"��sWjB���hЎ�0�Z8����wS�V�&o<#��
�Cn{ף=ԥ5�'���K��,�ݜq�#γQ��	b@U3�YCT�.�{���C]���Ntڦ��X�\9
ܨ���� ����tM�
3�q�XG(KLt@
�At��M��Dؐ�s�:3�7:24;!�p���2�uդ�{ʬ,F�����&�e��������zw�A�`�wwp�bJu���4��zgVw:�dB�Qq��o	�ڬ�g���:^��w(�e�t�R���]�p��SV�T㓴�j�MT-ظ�ĞA���g>nk6��f���s5�;��gց9nY���Jm+�WKٛ�=��B(��,�mw=[�1��[�ESs�X�󰂣�ɠ-L��bP�q�����ǹ���ח���U�#��ic�����j�'VL�{I}�C�g$��דZ�j����$*Cej�w`�-X�{dR�Z����g<��@��l�J0��(=KF��_S2��<2n�A�{�,�\������{�R���ڏ��M��}u�7� H`sF.�4>|c����`���j���{��s�d�3��������/�ݧT��v�Ƒcu���QE`}�M'�����_9':�z��."�r�娼bF69p`�.�\I5�
X9 ����
��w]�3x���[�ݶw���_�z9�&PV�# yRK��\Ӝ�\�6^�qy�l�:��h���]�Q�$��z��%p|>�k�(�Q�(�8�"躝L�V~�إt�-�;s����TQ]2]�+�U�ݓ���,��;n̮�G�p,Ki3�j��$m<X<��tOk�,�k+׳���0�'���+��S�]��{�׮�(��'_-�3�L]��9w�>��uNn.���'(QJ�d�B:�G�fWc::t��?�yoP�^n�ɂ�hhvy��m�����;���T�rJ������.��^��K�ț|b�*���!�&⨯��G�6��XIA ��s��`K��Ee��4�6���wP7�d�^�4jL���-�+r��u���ڒR��1�1auu�]}t	f<}�+=�d�Zʉ��� ����S.��I3i�^��hP|z�̿��X��,�-)�f�v�.��<i�'G�\�{~�Y|`��c��j�yO	��/��Ӝr�]X��� u���
JF��b>̒�+�g1�O�{*�{��n\ߦȻ�v\�>�h[�&��<��E3���я��e۷B��(nK�]c��]����n%�l�Aվ��l"����qt��S8�kPt��P�����J�N�)̙���k�eh�;(�����������Ѡ��5�ݯ�id�5:yM�C�;�1�xz"����wM�I���h|��}�v�\<ٽ�+B�m!���w��kz�L�5�VxRG�%gcƍxW\�;s�iKz��1a�����2�d���=|Frj��zˉ�t��n���1r�WR����bX��u�\)-Q9Kq�۴��[l2���`��Ţ��֎"Z5��ѩ�H�/��9�;���A/M[rMXd���M��j<Q{aΏ�%��a5rږ�9í�H��^�7���l�đ��@iZ�łī��j�@y5vqnb\�����`@7sj-ĳVt;�m5'�K!�+��9�qvf}ei]�/�l
�����>G��!Yqz���ci��wPs,��8�u��w*+*��]��e୵���s�RY����hWm�W@�gN��LP�w)�AyMY8���Y��иeN�ƥ�g�����	Qvɭ[��!j���p��Ȝ�ɔ+@`��_Nj��L\��Gz�f0�����	�Vc�`w7���zl��ZB�g����ڷ=ڰomx�4kY���D����g��؀��a�ݮBxn�W�G�*J����Ǥ:��3��7�:	��2o'��9���鹹Վ����<��8 xns�nr�v��k����;iw��r��)�΅��摧�g+:Ń�Dq�z�(��zäYظ1#���AX�[pfpX�B.���fp18���|.�	�Sp��4��X�3�
�%�f]��u�8�QӉ|3yv����p^�F���n�噤�X�[YV6g2q֣t�0
�r��<�݃fNӫ��{n;K�kά�q S��8��6��`��[䞵����y�X�L�r�Y�p_p��l�[�E��.}{݇V�z�A�]�y�nTs9�H^Ü�9N�j��&/8	W0i����EoBx�s@���g0W[n�vi��f]�/ 
�k�1�R=m�����x��[-���i�]�H��K�T�w-�d.���*�Y�m^-u���*|P��Af%�2��]+1�1�nn2�<܃�K��3h>���`l��1:޺ut�*J���u��q��l����Uٝ���{���
����3��WC2��lk颇C��Y��]��xA���&��5+�u�}��8�Kޣ;����!͂�D�1*�m�m�����G�����ʹb���̕���5jY���ј-ұn&]����:Ѝ��M#]d�B*�se���Uw�Uݬj���|����K��B�
�/w��kb;GZW$3��\u�馞�lˉ�w�N�ӠuK�"�;�՛�2�!�a�Mׯ�/��Cۣ4��n�O���p��k��'� ��7��C�:��v��l�CH�����x4�tTJ���<mT�w��.��0<�j�EV�o(��n�r珼���>o�����.��ه��.�DPܵL=�0͖Ү��-�(v��%� �z�<N�i�I�]KN�ͧ�z���5W�Vr��P�e��v���t�'�P�q��7��P����}tEv��H�X����[s����`�<l��.�`hde-+�d��.�]��l�ᬜ�i�&u체A����tV�٦d���
��]��VY�#-�	\���X�L��U�wx]�qn�Jm1ۘ٤1]k����\��*�m�Է�3n.��]�u�^;��g�P�U��n>ݥ�n6��Z/DPZ,R�d��`,Ӽ7F����0V���f,�ޞ�k|��eH�!S�l�L;#�;��&����ܜ)�%�D�R��m�)�_IՂ}�ׇ�B.C\�=���e��^��J�d��v4�Z�f�Fp9�x?C���9��]�����.)ca1u�R"����Ⱥ\�ݹ,\\1X��x�ѣk�#�`V�\��r�h�g�4��)�́�f�`�fd��,�ҽ�q۾�;{��4�v=��QQ&�v!i�8���N{l���D�!]Rev�*�o�F�m�Tg:OVҶ]��Z�̼�d�#.��7H�b������N����b�mQ�Y����� cu� C���)��uE\v�h�-K�%���)�hS5e5&�_P$6�ۥ��7�%����(�ݎ �A�*wfƋ4Oy�n�\%u�����K�ٴ��u���=Cc
�]�\��;N���Y��h��̺�Xv�pe�b�9�l4CF�/r��{��1�L;}{
�=+���왴"��Y�(�w��޹_-���7f��qRn-k�E�#�@���2�����k��lZ��h�Y.xo&A��WA�E������+/�E�	�
m�vd!��*uJ���.�u�7�H��#H��>)�h{M;�(_e�"R��6��P�ǵ��t:��n���c!�B�e��ZG$GG�7
�GN`ݳ���EY��E�CB���`���u]��0p��vmڠy�s�^p�=��e���hu����Z�^0��<��2��k.�gݣ�G�[��T�hR
w��x)Q�O�]�ԍA�J=��б��0��
�s;����>���P�l��n���Jb\Ԁ9����0���s�5(^gJ3f@�O5k�����8��z��O_1��C��]f4���r�G���^��˓!Wv�v�-9���Q�#G^�G��\�N�ph�V�qR�'��^C4[Tn�'�menJ��@ޫ愀��=�g\9���ďS�7x<t@}�I��]��m�YX*���!J^u-q���k��oЧ��K�gc�ո����0nV�0�}�S�6f^�]]`����@1S�������f�wLۤ��q���݊a��mP��J9A�ܫ'Wn�M����¬)C�"4�Lt/So"����Hu/���9��\�����֖5Cڤ��^�M��PN�4x������M�8����ą�еNV�t���xD�$+�󥞏�P����!r*��E���OS1�.�Z�G��������Dsi��W������$��#w!��.��ә�MY�3��)M�Ѭ�|msHs|6ZJŎzi��e�h��REN�n��S����oK�fL�h��-�f�<�+}xy7]#y����&8W͐�nlx����LחU��@r�i庽=Z�	E,Y�Q���M�j�v{q׭ҥF�44���l2Q�2� Q�J���P�9�b��3a-T�����`)t|�᥵uՙn�LO�dy`m]m]%�G�Q3�mn��s�e��؇u�ڥ�P槆uÁ/q.G�(_ 2�7I�u�V=�[H�.<��j Ey��)�9 r��m����Pn�s����&��U�:$�v�6!�F�_������������Q�����9]ti����w ��:ESh�B�m��$�]-�r�Xs� ��S�@�H��5!�(��B��IQڬ�m���r�����S��aΰ�L��a\�n�-�B�mr\i��m��Y��u)���U�Hօ��>�m���T3Z���:����[��Q��V��3�Y2n��3dv^;��5E"��lMJd�	����d�Hm�Й��J��~�:��<��g���`(��sZ�ov+RM�`��:��{�����P���(�y�`,L���2�me�$c/�]Z�5)�QrsTo�^(z�ѻ�,m]lr���8�X����߆��;��s�YGP�[�����`d�9��V��<�5�6�n;�V��ٜ��jTA]E��de.:M��D-:K����{�WpS��Ϯ��OU�1�����[?[�K�0k!۽��6��{nԭJ�+|�<�]s��XuǡZ�;���P�F+m�U̒��^՗�l�f����S�x�{�[�+�����΢���NHɻz�6��Wͦ��� �;�m_U�DVq�*&0N9�Wm�)�ЩO�˩N�h���7�ky[U��fӨ�Z��ff.�]#�z�%���V�N�P�.�zG�Ia�,J�z�Ϟ[�ھS����%jݦ�.��)�u��
��YtÂ�P�"�{�Z<��l�}����ނ��kI��PS���+E<7!��NӘ�0ݼ�L�5���\e�AŬ�Ti3y����z�{P�\Ȯ�/�{�!���ѽ�k_k�SOX8�	�},�	::�]޶8�7R���@��ǁ�پ���Xz����sT�̳[��K�����w�:����� 5yu_v�U�������6ԫ���cQI��Je���@p�yKs��w�v˗}1��%��[`�lǂ2�f���:\��	��maz�Ʋ�wn�Ϸd'�7���3/(������=���h���-��������ms�n�>G[��]:�]��_+���������L/&����M� ډȺ+3-�{d�{�k��Q���Zt��7�������] ��Ǧ�v�m$\䱎ۊ�^(��'D��R6����h�4��Ԧ2��O6�@�`c�ד.��&겠J4�s�s��à� �I�1�������%��n�T���2��>T�����%Mn/C�]E\;z�̰^V�#i+�S[�Y��֭ξib9GFlV7cT�0v��w�o�vt�1�Bs�	�bT�A�Ƞh�a��*�!�vKۧV��Kr4��zo�F�A���i��`[s��1]�����D���פ�Yw ��7�<T�ۃ7ά-mq��IC1�\�tB�%����-�ZF�p��b�PyT7�b"�VҶ�
ʱN��4�"c�I>��kW�Y&�2�v n�����&���Q�d��`�3��ª)���W��	ı'al��0%�����Q��G�WYum]�$�j�)e��AZ-����0�c�]+4���-;��ֆ��2˼&����h���WST�@���V�y�[�С�.�'�ш�^5�W��q��کH��\0X[��)�~�y.P�,{�`�$jb� ۖ��hWG��.-%�+ѿc3+uZr�8ҵ|��Φ�W	��XV�/��袅`S�{/�����r��ʸK�YwF�cD�:f<���rY[�\)Kr�jQ&��3RSC"J��#oN�2ٜ,b�+-Ɇ�%X��t̲Z�=H����,��q�CA��WyWv	J���0�{��-�)��'^��w+I��=�$��*ѹQV�t�΂����Mg�ӝ���N?W0'׷���C�-h;�;*�M���Q�ֶ�qQ\y8�պgX�ȶ�k��@&k��^�4H�a<�ʛ��MފX�:&�=x����Ʀ�������V72����p�dЧx-��1 os�nv�#��.TPA��nf���Iٚ�@.�P��@���;�|sq������x9��R.��]f�Dٓ An���ނ��i+�wT��v�bJ\�����wZ��O��Z�ﴦ-^k�Zƒ]����PYK��9�bmN��w���0��xs�Y^^�G�ܫ.���k3L��o�ܳsxuc����3Y��������bV����C�ڱ������S)W�Z��L�w�Y��19W1q����:��õ)�<K����ݵ��u�V��6�OF�ۭ�Q�˦�xw��v�ML�����^3/a��'�Y@���i�Z;�ee����g��C��<ڽ�f�ޞ���X����Zt6*��,�<�4��d�P9��ά�Z���#��Y]����݊�� ^�<���w0ԣ�e����ձ��e�%3����g��\����*�ݥ��Y}P)|˾�&V�R*_�0���˚UҐ�q�����9l3y/0��5����m��lw���O�V�;������Ň+>#�2�x)S�*.VS��p+W���^'*T�9*̆Sb�|[�|!�W9Y�C"�s�Y�7t��_:�G���U���&�Ax�쳳��-،lNz�|[~�=�e�B�0z�jл�=l}j�v �2U�҃WrM��aȞ�^.�+1*R��3�l�+�,��N���u�$��7��$��u���	��733 #x�K����&��h�Yc�ϓ{�89X��4��m�<OlN��tjF26��W�oZ�q�'�\�P�s�C�lEmɨ��S\��s3x˲w=,F�6YND�r�4�!�!ǩ7Rs�b�i���3���L�󩭲xw'j}�L�Y���6,e�w���y�o�F�i��Ye1�6W*�o�R�$C�ae �SϽ�7O~���{�8��������$���G�D}}���(+��#vw�,@ɞ�?���}t!�,1��*��++��7\Yk�܆ �qws\_S�{(Wq331�t}7q�B��9vO!L�K5z�o���cj��6[�"�#�MIci\���L[�qJs]E�Z�n�)��.s]�ɫ�	��_��>C59d�;�k���ц����9�pWt'\ha!|^��C�7�scܦ�CD��-��Z�ܥ�c�3_L������06�y\�S�+�s,��jrJ��,����J���{-L���C6��Lja���/�5�&6�T"���+*!\�<�{�L�!�d\���m���(8Ir^ۻ�eͤ�'��Ju���Ϟ(t<�mlov�9OE!{�벝��e[R���ǆr�6VkV��ZK?)t�� bVVv	���*c��
n�m�&�^��l aT���g|Y�]��W��ó�R�8�hk��j��p�[M�47T�ʹe����*�-2^E��Xom`K�U;h�^�Gr־1��PS��QX�W�2�ͥ\��n�v�u�P*�i��04��϶�,S#ι��W/�=�L�u���N=}�'�T��*�v3�/�G��mE��V��\�ٱ}�c7�m�[F��e��Cr�\+1�[a���v�-su���=��d:��=YZ�ZR*-��u�		L�S��U���C�uuZ�����B�3*����\V)�T�xz�l]WT
�( qܩy�)�[9;)<�{o����{n��iΫ-Tj�d�����O�6u�����)�Ll��Σ���ŷW��L�I>S6l�%Dڳ���l��5BA��)�4��U��L���ع�t�ޕ2�\W�œ9��5t`�ʕ��kW��:�B(*K�r��35CA�[:�=V��eؚ��N����;SPQ܈�6�e(��xVd%��;����:�w(s0�qE�V웽�٫�����1��b��&�fk�6�u�u�m��|uly������ٜ�Z{|���G��2�.��$þ��/��]�lFh��}r�V�1�Z5=�w٤��,yt���X�Fj���c��2u�L騏4�8�%7xV^��p/U]��ܙ��Fj�q��&�{�$�Gx��oX���T���9ʳ�
�Z���7X���F�Lǭ�_'uz�SM����!��cE;��8����gA�`������]W�Q�#H��ͳ�}ꒊW9���	:���G$ ��ѽ�^��[�ь:��JY�\�����QN��v�7:.�Hs�=�����[���CuA�>�[�ː�f����5d
�sh�F6*'33-9��i���ٺaV�����tw0��1�l�AQ�)V�$�P�hW����zH&2���CmX�/k�E��"#x�i5��Jm<؞fV�f,�f�Us,��;ݟ�c��u�؂YN��wq��`���cw���u�0�P����[;���~��j�݀���p����o\2��ݧ��5E�"�)s�Q��G���oQ$���,X���;y������:n�]l�H(>�q�oi�/��>��!Zbx��*���O�Sn���l�!�Ѥ��uJ�Y�3��h'{,�X�f�<M��2̮iѫ�R�7��"����=�PՉc���:�?whv�,�;����5��os��v�nh����鬵BQy{Y��5��6��eK�B[��1j�R���]��Σ:�L8�;�{)���8J5���H�S��-�%NRB���n�������W�f�0���I��J :pm2�͕��}��n���˒�=��mѽ9��iS�:�l,ǁ�^g�(7�rn�hɇL�ea��E�c�jҥ���Xd��iv��+x�Wxo�ܝD���G6�Z�\K�xv�1;��' 7h�[��sh�Esʊ�Y�4Rlj��LB���\%кʋ/^�A
ǎ�{R�u-Iś��Ѻ��J�{z�8�o����&�������lb�1fR��u��@aὗ���Zt.���O�<�2��^f,���&� c3��Loa�ɔq{�rﮬd�����M�{�\�x���	���Gk�?m�J�=�Du\��?(��5�9�o�
�XV�A��MI�H�in�nx����Jj����naF)��OE�w�T�g,�2�8*.šF*B`�v����U5Q9������Bev�|yR�Ww�L�)`������r��fp�
�V�u�5�f�7��م�˫�f�S�Pڼ�:6.��'G�U��XtkX�k�����!�1��k��x�]�evs���Bb�!���Z��_h�[w.!�%-�k�����ٲ�1ep�C:��˷�W(2������B���W�=�J�L\hP5��H��Ӆ�K(j��.9t�n�!�)M�𪠶-�A��д�ڙ��m>z_��b����k��T���$��3</
�(��!��c���n�ۼx �\y�m���^a�bfM��U�S���n������.��q5��'}�Qp�5a���|4���ʔ6�Pk\�LK<0Yh�+�SS���kj���1��N����Ex��WS%�LwY�����9Z���ٖ�l(�>޶1�$)�x=�Ku#��"B��֊��
w��Gj��y2�eѲQPľ��毮�N�k��[0Ty(���K�鈴�N�D�F�ͮŇ��ׁ�"^ݢ�M�J��Q%6,��[І7Ԓ�6C��y�=�ݬ�(p���x���v��t�)�4%挿���N�hCy�;���&at�e�n�la�O`�	\�
�-ظ��^zCzpzh��Y7�uC�u�e��וo0�DS�8���ϝ[�sL�:�m[�K�-�SSwgz�5�@��6]��GFZ����wkhܗ8Fw�� ə��w�]m�սbs���Â�V�j��Ў�7xp�t��7����̥��ŽX�WR��zm+J�-H�{�w����u,���N���jm�L�J�>�k��-����ʁV�q�$��e2�`2��+5�W�tf�����7l�
߀㛻�`8�v��Rr�ut^���O'\٩NԤ�1�3��x7%v���Z�l�LP7�73xՙl��*�|�9�$(��*�[�n}�G�Ϯ���Ӌ"�g�+'�^��&�e4�*[��L��O\�w>B�򅴻4ۙP���zQ���X�vjp���m�ގD�GS�]��f�V��ynh7t�x�tf�����>�N�W���z�o3CTs�F�#'h�˗Q���w�t3,ճ��#y�Vm�ިm�_d���m���繚s�|$��qxԢ/o��kK�	wYה���	=�e҇��c�8p󩫴JDᩲ�+P���k�������E��N����9�i6����x�Ao�N� ����������k.�ƞ�������X�{N��v���1SoN'�E��4W���Zxr�Gk��Eۄ��Plv�L�Y}�p���ܮ����b��-z2�q�a�M@���x�` �G�t�}�)�:�0��� J�e�A�kCm\c���c5oWe3��aj�z�EoKH^L	.�2�yb�}O�g����z�]!�"�Q�s>y٣9˨��g��Zsz�ΐS����-`v$[�ܮ�c�R�vZ�47���N��wG��Lv��u��KBl^Q�]��C�.�:Nw$����1��K{��N޾\&�n]m��w�!N]���O;5n�$��n�Nǣ^�-h�0ᗴ��n+�K�O�>͉`7V&�yq[x.�j�k;�td�����f،��Y&�����S��a>ҹ1���b&�U�B���t�&��dK�s���[c������Xp�Ӷ����"��,)*+��f�o-��єF�kV��w��`��~솎��pWY˾ʗf�y���PXU��[���7��D�����d�"n�q�9�1�m�|�}�חz:`��p��>�ts"S^�ץh��kQ�Añ�2��ZQb�7��+���[���]���˛Dٻ��k��z���h�%��V���T7춻Sg1�S�el�8"GgvuX覬٪�U����ˋ�w}V��h����6���+gc�FNѠi#$�|�;F���y'$��8��8��ȅK4�CA«>�a��ݳ��x͎����Ծ�-����*Ϲ���O�7[WJ��ű��p��xx���_ H��!��7�������)]������e8ʬ�a���ȯ�B�u,��x�*�V<]h��؝�Vj���*;�+ݎ�U��Ur�\@x��u헇y�!��]F�7�������!W\�|���S��Ύ��S��R+�LyN�;M���T*�^�Uw�q]����7��b�1�o:�"��2�<�y��+�ee��}����<Кv���>^����5ts�k��sU]��f�n>GZ��:d�^�h�NѺz�Ʀ�-��+>g2�6�XyO&K�x�jVzr+��/)��y�Y��W���9f;@�2K�4w�aU��d�1ŧ��mv*n)![�K־ԟ��k���^O1�)���!sr��"�y���'T�f՛�x�i�r�D��G������c��c�!�ʅE�QU����VOt�<+��Ѳ���^4�׸�;�ﷻ�-+6u���%q9��{h�K��S#39'�u�$��!� 4�궉�o��#5�58�����vh�	�Q	�����b���Ӱ�sN˧;��Z�멁�w���KUq���@������@͛����4La��)-WT4�[�ێ��Dn�D)#VԘv�nm
3���;���e	��+���)ҙ�:��Q�Z�P�P�p��2%�U���y��]���x�37*�l2z� -SÕ�Ynј�+,	�ps�+A]A��n�{�(�)V���$�h��]@C�;��F����ر.7Es�1�OA|���nlHi�`�`�>NΜ��Y�d�_  E8'��HJ`��}�^H �)	1I�.���R��ؒ:�`V��]���ӐE%��	{̯%�����M�zb�̺ĉ$ز/��.;�3��H��)�����mM}ڈ��Vu�R�6��l��eU�鼕���.,��k��+t�b��;�����w˫�Smvc���e`o��Syפ|�o|�l�B�{/
ϰC���ʌ�p�!�b���t�����EEיm?�ǳ4jfp.��mCF�9}����r�c~m�7|.��U�m>����b���~}Ҟ�1��B�(��?�T�bP�Ϸ�[�(�Я(�*m��ƶ��W�6�*����J?V�C�!���bSB�7E�|D^֩���B*�.�D�{�.��22v6g=0��G��Z4[�ת����ݺ�7�T���h6��{����b\�d�;�U�{E�ɇ!���>b��`Y�Yj_.�7��A��M��y�a\��ӈ�p;Z_ooS}��2�r��@'���x�lQw�[��J��"p��)wnf7Z���)��B����H�ӟ �]cwIҷ����s��̦2�od������<�)�v�;4����T����I��3VP�3oV�P�f�U1R��1Z3�5�����0�.�#֓���:�2$���C3�w$��w|��4x�.�Xb�)K,�����-
�e�� ��x����Q��ｐ��8��ۗXm��Nٶ	��y�c�N�՜�us$�s�m�E+��y�E��	�c8����ʗ���ע���%5����.��@�V,��'a�z�Se���.�K��mڛ
Ω��m]�*��=�尩��)P9�YZ���i�r{���x��<K,^�0I��Y�cL8�e� ���ˢ�S��{�[�6�ڮ��d����aq��������\ؙ�6�T���R�Pٻ݊Z��Zgpвt-�T؎�w;�$�]�t0�˭,��m����Î�Je�Ý6���(ڈL�^a��V�A �ؘ3o\C ��})غ��=��XX���#�R���Y{��vǫ�+��DĂ�쫠/b�&oWI�Lo-ۚ��4�'m5p��-b;����F��C&x�1f��]�2�F�^���"�Ruq[��������Ouˇ)x�o)@�%��Y�*D&w��5����!�d@�p�.xnmfAren����'�L�ӽ|ǀ�!�Ɇ�쥆,j��eR�ŃK��w�Z��w�'�ZY�)� �]�Hlg��8`�.;��R��K^����F)Y2h�؅=�b���"�\�]u-Tv����&^�$���wp%��d�2gJP�ܵ0����H(Ls��k=�pȈo���Y#5������#ա=��Ι
�;j�K�Dy�����C��5��q(��$f4�]�@*HA{w�VZ�\6��OzH������L�j�$'R`�\�^Ю@Vs[@*�J�w��{��`�v����#Ʃrl����YY���:�}Pgy>�Wm�xf��ȶC�
���&Pl�͐��6%�m6 z�hۗ�G��
d0���ʦ�R��3� ���}�R�_U�]K�mCQ��x��]�.�0 �Y�|��WȊ���Y�$�Q�D`��vk�}6��kǹ|��J�2��kw��7G)
>���-��V^�\��r�.FW��b��/e�}��N��� Gh�})v���0Ԣ��@t�����v�L�5mma�:"���{��5��֝U���Z8�kO	�Rz��8�o$J��.8�8Y�����N�������) *�	���[��U���Qvv^q�}$���!4ILr���GT�7�}��y����9��gߏo��$I8?SY�q�ѺV�I�o�݇8`���>ء�Mݳ����c�۴��Ѝ��I>1��X+Sb�5u�F��iw7Ӎ��IcS����B�1u�qV�9ۺ��#���-�D�$�%a!�I�c�Z��<�Z=3(���'�"	RA���߯3��lAr�=���ٗCrPE���LuR��͛��|:��hx��^���ه�*I�0��
�)�(ۇRU(�s/t�ñM3\�wB]WF����gVU���Zݬ8�\�0�����m�}�H2u b���5l��7K�1__R�
W2̡Z��*2��tj h���ӳ�ZJ�:ժ+Wqgi5����fL�&��ż0u����BS5�b1�����h�Wz���v*�/o���x*s88u�8�U}��>��>��m�IL��y*U����+nަ���E��)���o��^�wN��w{�[�Z�K�'v� �"�S���U�O��x4�����d�wB�j���<���'�
�0h�����ܬP�Y�5/��$�m.*�2�Û��ʜD��pbB��8��f�>Z�V�2A^���}v��ox_X����_.x!�n��^�ub��u&@�w��\����d�I �S�k���y��6��뢼���G��4d2�;1l2h�kq�!Y%�>W)<÷%X�k T[��	�.j�ܬ,Di	Su-�v�EDE��EDb������2(��TX�B�H����A��Eb*J�(�+SqX��(��F0T�(��H����\B��f2��TQe�UaYq
�h���PQ�Řʢ*�"�Kh�EE*"Ebb���mU�1QDb���QX��0�b#TYP��*�d1-�TX*�H�-��aX)UUAĪ��Z����1X��e���5QTQEPU)�C-fYEDb���8�0EU��8*�������*�\Ƀ2�TR���X�R�"8�+UEEEAUFEQX�
֪��U���Dm(�&Z*(�R�#�"(�Z��#�#�*(����Lcj��E�X��X�Պ��JbT����+X�Qb�X��(�"���#E�X�R���D�������E�nO��>��g�����I׫�)c�f;q��mښ���jKI8[���r�丈I\�PcnRNS���b��'�����QI��j�F~�x������b��;�3����"�7��_�˨��� p��0��
���t�q�As�u���P�`�4���<��&y�Q�����K.�j�θ�ݹ��継7�{|��/i����m����`�+�M�:�b�:Jǆ_�nq<vƾ�p��5���+X�Ȑ�q�|�.a�C��٩�{Y���l�D�������zn�zq��o��{lΟ�D�4����L
�k>����^��׽��/����ڲ]]�a/A�; fE��k�gHDABE�W�zd����LGc�̌����.%�g��}�md���Ls�`�y�f֎vWN�J�E}a���x4]=�	3����X}�C�r��߭�Ӧh 0le�M,�f띪-������$��zT:֫�˃�A��+��9�Ӥf�-_#�E�VX�z����6���Lu���1�N����}t�1x�19�eB�K�J
/����|�8̋���������m[�/�i`� +��پz�o�1\K5k;��ܡ]R�T�ufT�`Ҿ�Z���b947��+�%����$6���"�}ЭU^�&n�]9<�LSmd�YW�g�s��3�!��.�h�8��;w���2d����0�*2��G��M�R�G)�J�c�)i1.�:��f�ڳm㴲pm���Vk{�+���~^0_��H�N}O�0�tI<T ;��V���lv�cB{vTu(vl�#���L�S����x`�5_��7!��&ۨ:hK?���%MY�b/B��w�|�] 7��5�y�7֫�����_N��ա�9t���c$n-��{U�\���|8��\���4B��#_�$J�tg�Go����h�m�d�l������r-���ŝ0�Z��UB���p(�E>P��"x����jm�y�U�:��S��1[���QLaׇv�"\�����uZ<ɓЛ�9�|��W�L�L#�_a�u�~�s�k>�AVy|�x���ٺ�Ǿ{QgW�"�s�<���ٌ{tn��iXgƘ���3��}@7En^��P��	��>8/�}\L_۲ÿ�h`b��T�߹�!#]|:��P�x��+�4�~�K�W��)�����a�Ț��6KgR tF�b�cQ���fFa�H7jh!U.I�^�8-[{��h^�Nf�Uv����I)�V}$0�4�D��,p*���j�����g�uw:q�K^t�y�M<��{�Q]ѽ!]D5�b��U����웕f����YٹF��xh�j`�%�*����nKU���H��{\#,[ ,�CN-�&�%�͢1ӥg(Ł��{��L,"t�b3K�28e�@7�E�wC�u_PZw+�g��e�%0�+]u������7U���m0Z��}ƀ��O{�ۙ����ev�n�c������{7'ڒLL��:�˩A�k&�6�.Jn�ȇ�_;�k�0Vz���n��5zWx�qu� ���qmj�>^蜕��*f���oh�x�*�H�\폟(Z��v�W��1#��qqj�جZm�8[[$�fX 橑��G��t�p�J�0_�e4a�6w�����%l�޽��y�.�]��2x��.����R�&���Vg���*!k���b���Ŭ{f::wai��<�"hq-��	������ĥZi\^!?g�'��܁�YhG�Ӽ�'d��8����ǀ�z=�V(�@w��Ԇ�&�5A�.sR܎u9}'ӽ�䱊���C�*ˍ,�������8C�d�8�M)���&v���o��ͯ��.��8��I[����!��/\�7�Ha�1�'fM�1�X]&�'��(�W\f��8�;���_����͌Ԫ�喫V�^c�*K0+��sX��q�i �2���p�!�P���i�5�� 3]j7�e/�q���S��3k1�S��W4�זiV�,@�JIU����.ihG�ѮU����{qݺS�d�Fց�X1�J	�'��^@a�uF�T����b�������p!L���P"���Y*0�'F�|���P�@��'�b��T���Q��PW�;��E����ʩ����ؼW�z,�2�y��}	\�K��0��DTad�c��;���y~�)�Z+�)�V����$�x
����9J�,��e�_4y�����z;�r�8i�YG��.�˽9�K�J1��O;��u�Ƚ�s��[ �L�]�u�_ot柝���N��C*���\D�=�m���y������=�e�
4��Je���2����U�b����B�r7jS�UZ�Q��q��.P�%�(�RX��t�ϴ���k��x��G]:��}s�P�9�+h���q���Q��W�s�����Vl|�"R��7z3\L!�d���C�O�x�k����78��a�+Z%д|_$�>݇}�.V�ڽ����? R��/�[�b@��o~巘L�ծ��Y��f�;O��{����Q =ɨ�F*������k��v�����w�4�д�k�eF��S��)����ͦ3ݞ�@X+;�h�'��`���swaB���ا(3Ĺj�[��z��G�y���jQ/{؁#}����U���44�`i+8)��#+ʖ��Ջ�[[�QP�O���4+hlb�)��ٳ!�ɹ��E�nf�8ܑ_7D]9�S��Q����A�|.+\fɊ���w-8%�֣��=��ة�f2͖�}f0CF��dtt��6j~KtG�⥭�^ȋ�2�s�b�G&�.�un@Røs�즺�C!�VY�F2eן�b��{�8�%ó=ח&�d������B�VKF+T�ֵr�z��*d����g;�䣅n�9��D����C��'��p���]]��+�x��u)O!�5=8nf�a�tŻv�u(ǎv�$!�S�Bǵb����=�c�>�;�b��o�l�銤�V�t�ȝ�t �%n���n�3��qX�=�z���K,��,�����`����c:½��*�7Ģ�[7�m��ʘzP�굕���
���P�X6kJ&0B�ga�F���xB���MWY���d��u +q�`����sh�7V7��x�;��������]7u���q��$F��u�^���@1xa���I�����t��_f���wg�4�ꜯ��N��*�+`<u��x�s��mʺ�4İvl�<S8*wFodh����emv�85&!�=Wlggx�}w�Ө���hU�W\�Zܰ��8h�a	��m�hl��GΛ�yrLy.[��0��&�>�Ԯ�V-Z^l���xG^^�Xlf�Z�H"�W\��*Y�,���`��*MV�,�.�}q��E[���u���W��KT�ZV�����s�v�Hˋ�I�G3�U}�a�ZxH(�UP���xU]��X�t�.�ae�ۄ�]/G��K��l�\`$�J ���.����);�I��}�)�-��#g��E	�i���,�.�cj-��M"��t�%fw�[�#mB�S�]����s��2��oj��v��e�6�r�GL����*�����r�`cm\o��g���c�؈�R5���R��u�����/K��wp�A�ZoY�>zo�Ė�K������ݔ!��-&�.��o�\=�#��:���1ˤLMR�!P��.�q��X�I���p
�j�
0�9��5��d��]딏RU�Z5�����E�Nn8�9W&/�Τ
Ȇi�8Z8F�)���D�Q����C�j��h�7j�CTh����q{c���3__ɩ�;�S̙6��9�<�"�7�L#�0���oU�T2��6;ӯ-���Iױ��un4�֐e�R ���[��'/����u�)sJ���N]����k�:E���#8,��	"�f� ��2}aM^�e1+m�����C���f�U-�ӣ�*Eh�Q���vEͲj��u�-6���Y��^����7-͵�^}�m�X+k�;���xE�����/��R*�ъ2,�{�W��G��+�;���u8:��Ã�O������O���T�,�u���*�n��8���{�f��,��~�f�T=6J_�ր��A�Fz�f*Th�L�oGf<IU	��X~z����eT�=��<u��IO2H`�Ƚ1u;��'�粻�O-V[���W5]zG¯��Z��i�S0���Ek�����7O�W��*�͹��y�k�O��l��P�	�ɨnS/��=?w�~=�U�����5��v	"	�p'DU��]bա�o�M�|֏Un7"*#��k�9���m�eg����`,�x���UtܼX�~"���_��B4R�R��vQeQ��|��\>�̇0�m\>�8��YK�gA��F���rwXT�`xQ%T�$�d\t�$n1]Aw�p�q*X�5�у^{����{h:o�6���s��[��W�<c��PJU���Ls+!O�=����r5�n9�N�
�ʻ�J�	n>�z+�^��+9ͧt���Xʿo��E�L�]�,z���]������H˙���V^�Ր��ٸr!���3�� ���"�S;wn���l�Y��U��O���af|�D_>��[o��i���ANj�R4�ɽ�
+�r��}�y��!��3 d�:�'�=+A����)�ll�/tO��5���M����J&o*E}�Ҹ�3�8�kjp�6 �H���� �'<!��ENl��}&�^�,���ptq�_�x���.�&ۘ�2m��V�*\I�44�k��6��7wuh4{�[��Ѩ8�ʍ/�.#T�7��R|fLl4��-��jh���')S��S��*k���n������C+��b��R���:��w��'w"�&B���I5����j4����������{2P0�a�7gh�����kʩ��i���#���c}Ve��<9���K�64�]a���x��u.���8�cD`�)�yV� L�#�;�Z.�!��2ӯ�<�`߮�o�J:X8k��������߹����j�^��u���'K阉�m["U&Y9F-�~����W^F����c4���.ˋ�����R�{��?�����R�%:\��ن"���"�&T�y�
��``�����Oü�`z�#��z�3�L�=zh��=Rź�}Բ�U�Ӕc9^^:S���a�^�s�[���S9�na��&&��ٞjS���-a{Ζ�Gn�l�Q�)��� `#0꛵3WΒ�S��_;}�Z�Ej�81��=6���b$+wjq�hM\�6�R�|V`�)��8&}�������x!�g���[׌c	��T�(Gm���0�T�0l��2g�۪�s�l|�UBsu���&΋�Ϥ�)��gG��-����o�M���խt-(a�N��þ��r�N���<e��,�=�N��y�ϗFp���O�ۙ[~�D�u^�hm�o�A���N�@(*a���	�qb.A:&M���U��ⷕ���Y�6�a���"7��.�p�U�)}(��K̆[Wu������2��=�p.wJ���_-���]6a�l�r�`���UHȮ�<�	�5�6j�F��[�cH�����\�܀��nx}�u0�rՖp��n��f*�k��b���s8ܮU�r�����t��<kG��x�4�8=u�����=G�iS%�&/�4��N67�[��F���B���Ee.��ו�=)!R�O!�G��=��EEr���2��@�cCY47���'��}���e��k��ccd�L�Vr���U
c��J�Z�j2��ne<��s|�.�3��z��Zs�a�Y����.�b���{�ٰS9���t�ĵ%���u.IX�]�GuO���l
БM<v��14�əCUl$d�g`s�I��{WYo���
�`�-�{����W4�Z,e���&sK��e���N�N}��@9s����P�W�VL��!��r�X��l5��j�w�ȴS�4s��|O��}���*a�C��V����qY�2��Υ�2��t��vf�kˀ��=�D���o,�h���r�wۍc g��CY�s[��[�'��3����	�\fon�\�|`�*�*8�>�w�)���ׂ��(cI���L�p˭��r�J[��^;4]�=��:h"|� �� �O����@%���6H3~Ț�+m˩��x�3g�w��~�Kχ�_gm�1�IӴ�x���ֵ^F]E�B�ڽَ�w�o�#�jg69�T���ˇ�	�����ŏGX6Mp������ ��nWbu�r�nT��N���V#�ـ�C,P�\���jK/����8�EX6��ocg�ON�kΚk,�Oi�Fy����=�_K,p��k��D���>��PWu�N�ʃ:�yyk})s8n���2a�"�g���FxB�<4s����+=k�Գ.���#Zi���w���:X�s�#�X9q����c�}��8�&�H�{4iI��%���9�ث�d9` �xz��ת�nl}ή��]��)Õ����U��k�ṑҶ�N�}+���B,�'�:uo�T���;H�y��`�%;��QiT�À��q!�6�D^P�啎�9�2���Cv0Ww��W5��q�e���$�ƺhQq���˪�JN��J�n�2J�{�y���r�z��̬'�9������U 4�ݺi���.�鴦%����Z� ���O�;v�^���4�dۂ!�1�rή�5i��c�s�W�k�ڜ��M4��]2�A�zQ��X*�z�ѓ��H�ꔞ 5_�S�tDUj����M�V.����W�W��Wuc�/kkU�U�v"�
�ㆹ�o�9�輻h� �xu|Sun�ع�K�R�X����C�1M��.j�!'���Go]'k��{x�7j��w3����Fo.��
�B�ZW̚�m�V3k���b�LKyי��-����R�N�!.d����k��>�N�͋�� )N���Fͤ�U�@�����q�J�o��8N]5�n�r�M�̱ۉ��mP��5�@��'���aEɺ���C6�D`�`���硥�So����.>\i=U.�2�9`�����֗(��V���1U����Y�<���M��njtw��q\R���2��(S4��Ԇ1����v&�9ۆ�kܱ[Y����w��-,P$�}ݝ�isv�kH��b����_'�f�� �=g
�΃�/�=��~���o���{�S�=W�g0��2kBI�5pt�僓 Pe�6��e[ͻ�]t��[`�O�m�<n�V�N<�C!��"'��w3|�d	#Yʙ۩�*1$#=Y�f��V��&�4-i괕�8;7g �J�������4�ү��~�zZdw=4;�DE�H}�`�=P�g��ZX��R9��Pի�Yrs��h=ǻ6�t���.��VR���^Jqdە�ǣ�3t�c8�+��F�X�07{1�V���7��}t�
 �^"p��j���Dli��%򻨔�rY-j������*xa����i[/9���T�b�O�yP,��y��#���f޻�U�P�e�Ӻ�x��o�{7Ҽ�&1<UX9�d��J�&�����ˤ����shBc���lb����������sC �)�&�IǙ��:
?h��"�"P�[���b�Kn�P��ˢou����G:��F��yB͊Wu]u�
-c�iC=���!�(^<GN{i0H��U��ݍ<�P.���3u�1M7`�}xO\�ԍ�n�f�T�[����B./*��$��Fi�wlh�Uj�.�W���Ha��~���>�6JJ��m��K�1���ή=������"��Q�uɓAƒ�ţ�ׇ͔:
�&�P�r��4�ۂ��pg)�S;�<�}� [ׯGme*��Yӷ$��5�M۬�*c�7�`R�֊".�AEQA�V��\��%1*֪*�����(�)�1EeJ�UUT�PX�[lH���X�q�X�m��*���A`�ȃ-������Eb*���EVJ"��mX�\e
ƪ.&a���lb�$��R((*�%AE���"�TUP��F-B����VҲ-j�ŋ	��*���b��"��̊+ �*�j���AG(UTEp�Q��J��PAU$m
� ��Z�5*AEk*6�2��c�TJ��EQQjV
#+%�KKAVDb��B�kQJ��LqrŊb��c(1LZX��HT�,�Um����6���0�[W1��a�Z�ZЩ�I�Q*V6ʉhV,�US�ET��QjG�UUҠW���*QP����hj����:j��2�Tm$6��윮�(�-�/>>����ۖ�/bq�jD܌]�+.�]���R��"�} }#�B3�?!�S]��P������HVu����&&$ST��M�I�1�I��2^�~�<��A��d��ŕ��x�='����8�Pߟ#�P�(Tm�4��X����B#���N�ّI�
�ɉ���x�m��P��x��VT��'ŝa���`)9���zɬ�+4]sG�4�I�Ğ}����O��?9�$g�|CC;�m�W,�V����s�DG�|��������ɾ�:�g̗,�Nۤ�B��_m~�~B��(m�)4�3H|�@�0X?�1���u1�2�0Ұ<�q=O�%��7; q��X$��.qq�����"�P�����@�>C�c>�rz��
��s��m&!X�s5�'P��L����M��*|��v���O����_,�����>M'�/�M q(k�z~ޜ�?s?f����d�8��d�l�f+�׺'��N!|�ܲ,�O�0���j~O8���;��?!���u�P�b�<���ot�f>�����&����ɚ��Ou�{&d�rO!V��I	q@G�1&H?��
b��%@�{�u����Sϼ��~d��C�}�i'�Y<u��!Y�K��7�:����J�O��I��5�8���j�R_�~���O��^0&&[Y~S��z��,��E���I<LC�+>La����$gXh��?!������E�zɈxf`q+=d�g�<����N!YY.翻���B��3$�}���xN[��5뾉�����YW=�Cǈ8�g���J��~L�a��+gO,�<M����O>��qf!��fH,����S��H*���?!���Ry�`k��C$��ʀ�����|(�kN��΍VE.�N?$��������Ę��R�?&��y��M�|�O'���z�Xx��yd�1Y?�$�1ĝB���3�?8��4�Si�3ϼé��`�#�,m�����s�M�Wg|�(��z�?�܁�HV|�fwDǬ��ɹ�ri��;I�=<�x�U:�~���ă�?3�iY�%d����O4�?2_0�CN2bb���bO���#��WӂP�0׃�z�n�'U݉��O�]"�M�"�]��t�>O�{|����1.��M4�n�SuYUg.�L��ln�cņؤvN�
�T��b��Sx̉��#2hۓ�`y6��]u��L�Qq� ��B�K1g֘�N)�8\��/�KAt5;s+����O�}D}����a��>v�C�+����&�i�Y����AI�{��:�r���eN���Oɏ{`c8�a��s}èx�P��e��P���=�R.'̘�	�ׇ���X����>��}}�X�'�Ȥ�g��4��8�O�7�jI_�l�x�LM}�5'��!S�>I�<� ��O��S�I�?'��y߾�~k5�w������k>g�bAN���*O�T5�L�&!���VbR��<����:�&�����<d�c?s<Ci/Y<7���ϙ*��.I�Vx�Y��2~C}�q��W���{�<���Z_��4G7%1��hB��^���Y�<q��gSi�|-L1��e��(����˧�i
��Ě}d��?�E�vɜ���/2m ��K�{ݓ�<H;�<�g﷣\�9�]y����Ϗ<�^��f�+��Oɴ�'�3���m'�̘��B��W�����HVi����d���C�Led�8�.�N�T��e9�g��)</�g��I�����|��秺�����y{�Af&�bw��h*H(n}��xÈc'�ɯhT���&w0ɦx�r���i=B���Xk�B����4�����c��m�Hx���#��>�����c/��k.�w���^����4�a�
��~�i'��=I}���L�f!���?!�}�l�4�0>�4��*N�S�@�):�&=N0��*rr�&�$Ӥ�B��Ʋz��3�~���'�������ǿzo��z�����&��%@����c'YY�J��!�/,����2M$�=q'��wA�R�I��X�l�bAw;�8é�t�!���4����׌Ӷ��z~ͽ����?g�����~�O���f�$�L���@���L�K!���Pݳ;I��w�}��'��Y+?k܇i�O\g�}��:�2}=�<H)8�~�rM��HV|^w_}$��"�B���Vǯ=�b���|ͲT���ˌ�]���f�.P���L�cN0ݿ�I�O�yu��z�$�f��M��~C~�̆�B�^��?O����g���2bN�Y���Θ�m�����>����c�8���Pϓ��=���@-���~�TΈG)�[�m��T���W�݆��o9�z��	�h�t�ۼu�J�9��=Yzkh�]�Md���:��{��S�-�kCtA��k���UtΫ%/��U�ٱWÄ�g1�����9�t`q���?k�Vx�P1��ghc�d�z�M��i�V��8����=�<�+>C���e=C��Ag[���3��ɬ��� ��A�4J���r�%�ڻ������ԟ�����5�O:���j�}I�I4���6�W�N&y>��H92m4�̕'�i��Ɍ�񇩉8��'����q�8�N���
�0�g@�q�󪆛�Ŧ��u��>�>�����g|������`VE4y�tq�-�~5̛g�Ǭ���w,�L���� �|�Xk�'�b���LV~d�� �i1�D��/
N��{Z(���:��P��p����a��I�`):͜�m����i
����Y7l�x�C�m������Z�:�U}�i';C�K��hg�1>g7��%H,�����i���@��vX�N���3x�+􏘏���c;-��B�^���,4�Ԭ��j�Y1'���d���Y�^��`q����L�%@����[`�YY+��:�a�Y���4��xD��>%4��}u��>��n�Z�'�n�
ϐ�:t��=LH)���?3l�:�0�
�*'�b�yI�2�Y4�Ĭ���6�i�t����!R
�ɽs�<I� �������`����>xi?sݩ��[�M���;�
~<eg�����b�OS��s�`):�\|5a�����Xm�ϓ?}f3�11�<f̺H*Ȣ�i��x���~���8�&<d��<т>�>�������{F]����u����C
�sߵ&�I�I�s���&+=a�}�h�8�돝��6�HW�y�M�Iʹ1�&&}`l>�ed�����nj�I�VJ���t��|@����W[��g�New@+o��P�~d��������15��8�H,�\�C�=C:sXiYԕ���g��e
�~M��I�J������&$�|��d�k|X(c�B��>��1m흅^b�DP�*N꟞;`�YRr�I��c���y�T��ɈnsߴM�HV|��o��!�:��9���L�8�'�� Ұ��a��!�����g)���|�U1G�`<+��x,��z�&"�3�H��ݬ��ŝ�8fmh�u�jSn��%=k���ҕ_*20���Dp
 ��6����ڕͰiفaY5^��N`��f���S��ۧΚ|'hW���7L�����x�Kye+�:�����e/��pb)U�͝"����{0�����L�e�CI{a����LB�kTϯY>M3l��d�M��eg���i'P��y�}�U������kĝB��8�������Sc�}�=��.��=�����R
�(����6�m�;d�?8���l�i �����ԟ�Ă�����K�M!���Mr�d�f�����Y<=�5�4�Ru
���Rn�n�꫺���5����q��1����}1;d��l�/ri�2[d����P�%ed����b�d����Ĝ��P�l�R�OXg��u'��Af��揘x�!�����ҳ�+��b�}��#�+��j=ᾗ9S^�����t���%gg~�ߖi�y�;������w�u
���ߎXz���%AC��`�YP��4����>Ce��'�ĩ�&n���=�X���$}����@'߼��|��]_�����1���g��膕��Vo�r~Ci��s��x�>�b�y�aXT뤝t�l6�H+�Ρ��M!R~B��ɤ�<I�*�ģ'YSF_�����@��k�=����د|G�X
N9��Rz���<ާ�>q�3����3�:�ÿ{渇�Y<��hP�z�<`_���Cl��Lx�v�i�����{C�=C6r���%�`��4`�jɁFӍ�dn,Q���i����ܤP:�8��g�L��Rq�ky��'���S�f�13��a6�2[d������������u�u����I�(c=O��C~S�#���g<���1i�h���B>�ă�rz��m4�P�u��*J���C(T=�^�̘�Įϼ��&���LC����+%�<��
N�X��u�Ruf�*~7�'�0Y |D{����(]ț^x�b���OɌ?'M��j�R~OS<;��&�����<h2|�������5Z��:�� �)��:f���ޘ�D�jSS�����9_v���(��bO3EG�j���z�EO,�/��K�7�.��ɷ[v;}񦒗�}zo$�%��Z�m
��]4�KP�R�:)��@X�x �,�}:A�/.`�=���M�	�e�1�*؜����/�K�O�ů>��Y��/�b�cw��8�n���dD���f�g�T�\�@ټڨO�Ξ�!��j0����ȉ���(���'I@.�f�<��	Q��V�y�zˮ�3��e�P�[��,�,h�6��\!pM"�P<j���Z�q��Uh�P�=� Hd�0rq��)���[U��;u��C�8`�K]�v��\>�pr�6Ԕ����m3�"bI������艉0��_l�5;������p�M_�^�3f�բ��ݝs^�	��C̏kV<��<�y���Y����1��ʦю��ozyw�b����},�*�?�z�135�58+W B|����G��R=]���MIٙ�ltWr�X����Te�Pɨm���i�8\#�UJ�5(���Bf�O�%��8́Sq�̐݁���Λ�O��;F�����|�I�S̙)�Z�yv8Ex�=9�����E����3�ת�X����g�W����zWU�-����F����P;q��&��e:FmBw���q`0.a����a��q֫��ݔ�����%O��O���#�0��ה�[�Y��E�m��ڷm4���
��!�`u#��wKi ��<.�)��;ՠ}��(p�iv�����`��%���1���y-έ������͍7HG�� 9u!�*�9l͡�l�ƀg��3�&ƪU�cZ�1��խ��$�6�g9S�O����Ƕҳ���u��9����鿉CAˌ�@
�uQbFŔ╴�,�7��-:�b���;��u"��K9T}Ϟ=I)�a}�a��\U�EEFs��{�� +s�Ȕa"Yb�j�Ew݋C�ՈӦa>t����{��]r�HVIH-�ۛ�.+&!3q���&���_m����/�fۨ�zZ82�$�.j�ua}�YD.��\���#0/|ѷ-�5�1�)���]t��s���nS+)�������k��6qBT�A���$�:���L��geU�8��_σ�3�gf��VOc�v/^����W�������OW�P �9�t�$n1]AwM�	*X��o.��N�n��e��s�wt�i6uÞ
�0��rQ���> �w�����P�R��l�u�v�ee�R��U�Zq�Hq7���	�$yK�@�����'�W��|����۞H�N�y����
��I�G>s:!��v����+�6 �H�|jR=[��0���$��,��-[}XF�{n%J`�vew�_i�n���U�<���r�jB��Ӽ~���yۘ��}�)�Ķ����+�r:׋ѵ��w���W{\l�5�^�.����v���̺1&E���M{X�(�9x'�=����h,�g�>��֞QT�X�<&�pE©L��
S:8����ܛ�nc��d�U�J�S2����n�T\md���~�����3�)WK��?������Ƣ��s!2�Ԙ���&ۘ�}�\��x^Lce��ָ�������fs���`�5�s�Kc��ã�^˿���;�^��te�mB����y�8���I?H�#����[@��	��b��wO�e�aϺ�}�L`dF5RdT7l49�5���uLF',N�(-��:�S�	���;��X��br����\��;C�8 �ޔ�����$�S=�u�G�L۬����@�%Y��U3i�C���贆	�n&�����J9���L_5l�I�NE�v�W�q�:!ٌt��ŵB�Mˎ�P�9:�td�ٗGԪNl�Xن"���)�edT���蘻��=)�l�7ѝ/�Q�����B�2��3��X��uRC�	@�_O�#�˼�]mM��{ݕ݊��6���9�)vT�B ��g��p^�|���6>�F�E�z�_��ě�������r�mn��B��W`́�yw\����R�/�'0�~/R�~�}x��{�?_���T$�v�=��rV�[�c��xk�X+"t����۩�%��/N�7���q�m7*��q�FN�|��e�]�zÆ�#�$���X�����j����;�����0�=�7_,.&�G\�Ƹ�J�?A���*6�"����"of+�t�:��GU�������Os��k�!ay�#��TP,�u��N�Dycs�^�g���oIv�e��c�;1�U�ڱ�r�WfY�7�a�ӐܑM�P摞$4t摷4X���E+q�k������W�A�P����[��z;l��-s1���9�T̳��t��ς7���(z�#<�?L�_#�����:��0����]l �TYQٷ�n,ް�����>y+cC!7�����Bu���ta�X֏#o�������}-�b���m�65R����ϳ��9`sϪ, ~�TE.0�`�4��:c�}�i�6��[�8��U�'v3%4���!潾	��+ !Q�ɡ���Lt�z��a��.a��d�����'jsx�⸿���{sa'w�S��zl}��hW3b�h�s�`o,@��A�����ۢ�d1�y�����SJ�V���A�Y���j|�g,���e̬��ǔE���55W��6�[��]2�wn�FS:k�!k���G=�ow=���"Gs�(P�^�I�.�^�3!�X�,���T�Ea��ɼ$;��г����^W9u�����v�	y�e]������iwP>��z����BO�҉��:FNsU�~�<9�(��k>����%ͣ�\��I��s�WZ�7�P8?�ou��u�AuB��]x�NSQ��cc��fD�3YZn��ݳ-h�X���*�=����q'EFnT�(��}�k*����:�Fp?b�Y=�Mw{gj��|�O2E���Qn����\<;)c�v�C.�BN��=�ʏ��^�-�d���'�=��'
5��r𯆈ae��L��T�gӕ��Q1|P$�S�H}�R΍��爀�=���b�Lk�X�4�[�5%������:�t��}����1Z��9��'�xL<��i��ֶ�Y�v��,p��:\T5'J�;S��Z_���{Ǽ5���{�+���@�
H�0��_l�5;������p�t��]����0��˧�鱮;���~tt��~UƇ@	2��i.��o�W��12.&�`E��X�8��ɂ(;���ˤL\35���\�F�0���&�3�:�{�/�^�F����u; G֠b�B�l߼�x��:Y���f#��<�4��`�t��v�9a@0�>��6SUڣ�����t��s��q�[��Ȕ,�̀nYw[��H34�.]'w�s�8'�b���#�)E���iTH�}:��]��.���'���J#5%w:�^3L�
J�=(���BfI�w�x�X<��4D!�W>�-+��Oب�+Or}_ɪ"�O2d��j]��I4�{W�:ue4��q�<"�ؿuR�|+Tc�
����0ECNx�W��fC���]�ň���%$D����;���°ߍ�^렫iW�ྐྵ\L\n��h`bҧ�Ù[�/*UHJ,�bUå�����U��*p�D���s+�j��P�r�δ ��Ir��5��;;t5�oZW�N�]�A�cQ�N���df��:��҉ݳ0��Ū��|yX�nJ|�Wn���?k��>ܷv&-��FR�l�,E��iW��'E^�I�L�|2ҘN��(�}��cT�Yl���\e��7�!#����Y5�9L�߭��u�_͸�Q��Ԝx���as"�;�Z�(JMa�aT	���*�2UH������`2��r�YM��7���+T9��YE�Qb�u�� `�����;�媡+�1�>�����s���yMbس2����j�2&�����߇��n�ھ��̬wn����iZv�"�1�X>Ǹў~E!kt�4��"��H�!ψ_^�#�4㫋G
I�t��^���нf�I�'|Ӊ'�V�m\
]W-!�[���1�e9JQ�s����{mRa'�V���E�V)q�L��(Q�+���^�*�dT:���B)2wfg6lE���X�U�3'R5�vU��p@`ع?��\�G�0�<�"���б��TxoY�~��g5�9��ið,#z'�\��M<-�ȩP��{������c����+�i�b=Y�GZcq�[x'b��w3	�W��)M.p�vftt���4��ʽF���g`��7xj��4���(i��:�I�879i�T5\�!}�cZ㢄�C�H��#]��c�a���\Uj���{j�;�Y����L�j�Ga����UǛ�i�ņ������{e�`T�Y��q o1���*{��G yX������Ģ����5�x�kQ8�f���,�3knѱ�N(�x��k_^TH��L�}��
?'N>�v�=���S+U��7��i�r=\&
�*�v��l��;��X�h@����{n��{������.Q �;��W�����!^���� ��q�����a���A�W��u�ޜx7+�2(l���N�S�5|DW�E<�S�^�����'���\��Z]����k-Z�l^'*n+7{д����$�9��C���;�y<��yѾ!�J�,�t�u�W5N1͆�ۆ���9*��(��^9��*�R����Z|���D6'�F�v;��f\@^Y��&��x��R���̈������}���_� �)��ٗe,��!��Q`��V�8+�7�\�'1�g5R.�����W�"}�seKڂA�>�+�t,`����L	�+@-��b�i���9�Uˍ&z�V�Hƺ�vf0pP������1𛻍S@�6�����:f�o��J�f�3E��������it9��ا	�K3����{w	����6�^D7RF�u�q��nH)F� 6�,�\��u�܈7:U����A�t�����5�v�xr�)N��Օ��di�w�W�I�N0�R��-V氙��b�A;�r��FJ�Z�ͽ��'b"[�мg�{�ab+�OMui��Ҝ�����T&�py3��X�z[9�k^���^.o.��[ȃ�e�r��9
�Y/���b��M�7\���^��z��&�b� �o/vŤg#h�d�n�0�v蝠��,:�$���YcsO:������:A�SU��������o{��6c�(����V}���&+N�� ��et�2�Q$i��TNȕ�����Y{(f�V�����yם�B�vF��u��:��\i���x�Grش����׻2א���gﷵ1�Ȳ(*�$�*),����(+k@A�djTT�m��RbV+mA̸��+m�b�b(�fZ������	-�R�AEUeB�r�TEX�QH�r�[eAd�QAZ�I
)(�EE�e�"ŕ���X��Hc
���0QAA��QE��E�,XTPQjJ�������h�� �PYXX� ��b�()�����[d�"
)Z��8�r�AIZ�,QX����"*ƴE ��,��-��EX�QU[J�J�R�ܸ,X��@��PD0XE�e�U��`��,�(�DH�h)R�D@�U�T��QAZ�*����+"�PR@ET��,�%E "DUI0�[*���c�ZE��bc!�~���P7H{}\ss�5�6��C�8Y�?�F��0U��7�%R�GZ7�;ri�6�Pm�u}�EǃJM�Y��G�\�nN%�(�nT-��g�B8pd�ȃ(	�{�ȸ�H⩂���0�T�"�u\�i��v����ȇ�p���p�S`\�h}�����e�?dSVu�H&o����m�]��S�N���)��熒�f ��Ӂ>H�� AHx}�\+�����=���g��)�=���'�ⷄ��������D9��Z�t���1�|���R�]�V�d�7��R�Ѻ�loIu�7�p�-��%��6˹Ｌ�/�����|�<�I(B	��x+)T1"����V�Nd5�1M'fH�,+���Bo9�����GSU`*�)e��y�1}�Y�X�]h;�ڃ���W �r(���B���=j�$�C�3�r]~�`��*�m�'ΆL.��~�.�u��E���s�#2�'������XX�n���N�3ؼ,/ƐU[�hS�	�;�f*��zY{�"tPî�{����wF3ݻJ����[7�����<�`���/EG~TE�^Y�^ǥ�i���hѶ,2��VZf���52��E[gst���Cv��b�h��:��#u�ث��OX_2��1�����c�����z���]Ġ�r��1�Ŵ�T�oqO���5h��f�
��)杔�0c%ƵN���l۬�u����_��3B�� ����t�U3f�Fi(�1�[%Re�")����Ӛ_]�-��ڡ��	~�)^h���kF�6m�L��O��6��ѕ*�S�.�V6a�����\�{n�eј�湔���l!S��5�6+�NeAn�Z`����+C�
1��l�Ӥ��Ő3%ԮC��dvh��-�ȧ\ό����7���|~�*�����u�M�kݺ��KU!_r�Gf�����z3��a��C�n�zn&�G\�ƣ�$�3>(��rE��O'�J��c;�UE��)SÑ�C1�d���{����,�r {��;�u�:c���XYƹ��"��eZڱ�r)5q6e��p�a���"7�n��sH��-��h����\���W���]-d/�y�´�e���[��{�N�1� ��G�Պ7u�>�b}��O{�Q�[p��s%9�5?(�A�htW*�7��x}�u0��'.r$�������g3I�^Q��@>P���G��}X֏#o�����僧�L��� l�
�jg{K�&p�N�RWGm��7Z�L�k��5�K;z��г�/�X��+����.��m<87oe����T�b��!B��8�fV4�	�O:v��|�*=}Y���ǩg]�����}Y����G��PWS�q���G��\�i�gM��C�qT~��T�y�,y�E�0DTqD�!i��2�^�������ͽ�s���ƌ��q�5��:Urn0��r���mX��^��c�Ϣ��Եu�S��h�.9ʘ���S�5��6��~o���`�m���@r�H}r$�������ڕw�qk��$��ʖ����L�C/���;�3Gm��ʘzP�굕���[9_y,�����|����g�����X���,�7�~�xx���p[�c 9sFi���"v`�̨�w�ܱXu�V7��x�F,�@Ya�2:�L� 1�a� �ҳ��\v&�u�r=Og��k�x�|��4�š��Zn��},��"tTu���v�n��~y��}��Nw���v>�-�*ܦ���_;�����~hv�Cff,��~¯��gHge�ؔ������v`��}�]�χ:zr�ae���3-S����&0k���Rvz�WhP�zA&��5J�X�)��H�ʞ�IgD`�/j��p��~�yW�m�XYHG�u��̳-Ԍ:�LV�nC��H}�=0P��2���q-mh����ug7ÄeK�X�	��T)�ݝ�[y5{��3�q���Y�JS��ԻZX&�����S����Vj�����|����.f
�V�K�B��pu�r�]F�j��������\�r{�~�� ����)���.��.���Z�#3s�3U]sɉ�rR}��[���K>~��
�<_���ϙ	�Hu�w�����Å���]�EJOY}��3$����u�M�Pt�	g�Ƈ�	ZM%�|�����(��Z�5A�F�w��tM�ۂ0W�5hg�]"b������R� B�|���ɿ,��]�G���Xkq�z����:�����U�m��� �h���0���G��F����-��w�z�,,��~���T�gh�j���������x�n����eW��>�kq��E��U��zg�T�"L�¥�����k>j�z���ȸu9�����fF��߰�N��)�^'�s��4�4T-T�
�Bk�lg�q�5{�_ڨ``��s�<�T��v ڧ¦V��9�;w�+:!9��_y�j]&��n��4�s$��Z����뛍.� ?������gQ��Y��hn����b��о0��*�G����]�z�0�;e:r��!㺹�q�Or���W���:�뫺�"1�<p�2��B>'����Z�g�R��'Vs�i�J?q(���ʭ键o2s��T���73��m�e R�՜�0e�S��}�#Kf���u����P�GJ��>�vi�k4T>���ei,��ϝ�qJa�o��ZٸiW��z�B�yJ��k%	,���_%�qUCu�Tw��h�l�Y,�k��_o�[�����m���&q����͙���T�ܒbIc�΅q�T�PW3"61:�X�L��V��2�&#�	Ȑ�y��ڮ�k�f/L��5�9 �0�
��}o���}R�0��_�ׂ�d�z���1��3k���2�nq�j��6��(G	��$�A����E�LԘ(�՞˭(�>Zo�=������=,`n�	��=p��P�T+��rQ��>�(%*�W^�@�򭎾}]Rڂ]lZ7�m}���.��9�|u�ᤦ`��R]2zT �1��8]s�R�U�ꕝ��B��_M�����?_�'��N�8�tCe��a��)M�=ϫ��[�������� D��3d��<��ꔎ�Х3���]nM�s!�s8�y�� 7�V'1���py��=M>I^48��{���U������Jө̆��Rb��}����|�^�)*�(����Ix(�����0��Պ�Y����Io{��ч�/J���i
�m���6�	g���캷W`��g:Ǜ�Y(J��1��6����ZŽ��ʼ˧���\��V��q���S�
n`� �g������WՎY�f��B��n�	�c71��j��ʯݔ(�b���N��~�Vƣ	����S������7��E��S<��#c���1]H5��q�l	K>�����ms���kbOe��Z�+�����/�Sbt�,P8v�}m
xa9B�x�S�w63aO�>��3�P���9�T�h��-��T���L�7_4n9�A������0E�/���O�{$���k��/����NSJ"Q�٘�橁�J��'>���6��F�1��j�����������}���˪K���K�Լ΍j1貵y�,j�"���#b-���9�֌/��sI�7��ۯ<�N��8X�+��-���t>�lb���Ĉ�o�RJ��їUgw�f���C�7)�����(��N�v5�f��_��+���WS���S�њŶ^v��\쏨�UL6�C�a_=��w��q7::�\�(a�N�|P����o�Vd��U�Q�\Jc��wb������PR��"9�f6��Kޙ�
��_D���v���{�Ef�ـ�g�"֌W+WoRC����{8=0�'�E���'.��7{����B�gc���gI֗5���s'�dC#�{L�_Y�0�ՍA-���u�F�U-8�m��(�W�� m����^n�����1;�0H�v������C��+��&�/�/ �PV��3�����VS=���1�r�#��"̥o����U}K�x,�Ns�ˈ��D8�$lJU�2�B3���\;;l��-��0(7-",���wTΌ%�� ��iA����Ҵ�#��ž��7(E��<>�KX�-�<��LK������XjS��l�ξ��Rt�v��s��c"2�C�8R1S�,!��+DOBo�3��P���B�3�~�IS%�r��Q`���� �Zl���x;����ܲةI<� �����$*]tj{lbj�M��������j�g�O}�ǻ{��cO�q&쾓F|�-�pﯸ����)�������É�
T�6>ڇu@��--#f�%�TΊ�Px���1}V<2���x�r�=�?�
�zP�굕��̓�̍�y�,��	T���
�MC1`٨�Ɍ�0����Zo,�#����8���� ��fmk���B�N#�M���1Q�*t�4c�*�B��]x�J1��k6�3CNq>�vh���u��}�ǵ���kU�y��0夞6�{u�a�2�M<��-�-����<�Up��ݻX�c�+�kj�K�]&:�,)7����^�{��|��Pp�n�oFiwKcH�]�[�镇�,�KJHH���D}щsp�MOE�����SN�.�=�J��6�tVnT頉k��`�l	�Zh<�$���P��t�W�y]�����"��n{m��.�1�'��hv�왘��� �һ����e:��wJK�9_)0���$j1+�Q�^4C-��f.Z�;>���x��Һv-[=�<�^�'RZ� ��pW���4�%r���,�1��ӈ����p����<��ڛ�A�5�\`�Q�@b`����gAH��j��v�鯜���Jgs8t'wv:6���ᘷ����������	�:����}F�>�y�ΈFxB7/__M�%���.�j32ꮅ�I���icq��&ۨ:k�,�����t����|���{���=��)�dES��V��²�󞖃.Q0������T���?�GWLA�#0�}o(��,QV����g�>�1_kF�9L2z!�\bXD���U{X�a����ز���nt�әUv{�;��ւ�?vӘ��lx)����j���<ɓp��9�VU��lP�o�s�A>��Q�>�Rv��tD')�h��E�J�,f�<��[����Z�T9���ڸ�O=(�U���C8K�^>��[|�B�	+@��2od�p�k.�/�����Ƌ�u��Rcf�;�m�O;^n犸Ꮏ����,��Y���^V{���$���5|��=��i�q�J꺅����SaU���=OJ	KP���ngzN���tK*�i�<�Z��AVM{���W�(2�maն�n.E�
p]:}�o:�!f��ueX�\�ƔN��߽VNT�����:p���d �~�\lp)��h��@��e�\�s23�n��_��|a9�ET��bm��f��yM^X΍ϟ�]P�'�+�� ���x�U8��&υ\�u^���Z��kl�~�w�-g؝G��6�`��uALx
7]1.@\K,��)�������^eX��ν��5Ў��!�)�>qiQ>a-���Pe�ȧ���t��0XH���Z���:V�v��D�;��_�)��㢏T��:�* � z�[�ʾ�a���avz�Y�pk��W��a9���ht�g�`3�ڸ}�g<~+��>$�* ��$/�J�,`�X[�{}�&�.CS�p�tV�!"�\����h�}�������R�QDÃ��"�ܒBN5��Ad�7�Իֺ�I�ޝj��e|y.�w�t�y�'�����P����4�:��c]t�_t��3��n�Mh1Ŋ����#�[��8]�O���2��M+�v��]����^�z�"�,u�7B+ŒD��!r��}_UUf{�n:SFx�#p��:��B����p�s���Hq6��e	��Һ�w��
j�ô�ou@X�������D��k�+��'Is:!��v���@Tv��ׂo:3<Ni�
��  )�q�)�)���%��cD!;SS{�[i˕�uL�&�*��N$����E*�]x��.��4Ƣ��s!;��V0�ޱ���d���Y�`�+�'ޣ��<0�8��Gր.�Te.�ё����_-"�iZo4���w�_`|�܋	��k�nX#��4��	����]�~���u�2e������3�^���������)�#���3<X�p�v���f�^�qk��s�QM�v>2:�T�_��iV���S+��V�|z�o���:�9��]+�tV�юϡ;՚�������ENq5�zr�y�����[ �L�_ݔ&*�Y��`,�~�t:O�߻,O���*Y����Jt����:2�T�%��l�1�bh^㛒oMC��u�Mc�F�N�m���ťx�p�W��Y�(ΝP#[�����-ٕ,��M�&���b]F+�[Y�ʹ�S$�5%c��`9�]����#�˜rp��I���ɭ���i9YT��v��91�<��=����� lz�eU=��i����~A�Iv؇�8��%�v=�Z��=���t1��m��?,�g5�S �6� L��ٯU�/t���Z�&�S���|.�#�����Yr^���g<lm
/&�KN�w��/lnNܳZp]m�{#jA��`��X&�c���ŏ���0۬WH����7<Y��g%���#\g�%���uu���Q��}a��;�ۤ`ʰ�^��{��畔���lX�u,�]v<�H}���h�l[��Yz���C��r�l<�LF�h-z���{.�w�#�Z��.��'�I����[��Ь�ks"oϥӕ�E�S� ����ۓ�ԩ��P4���QUҷu������
�*��\rs�8���wP�ژ�-�g��+Mkh�n�LR@7Q�����N��r����p)�� �5�.]������ʼ�7y�sk�>�8i6,v�}�i��w!K��6<���ّ]~�JR��r0��'���y�,��g������'�eBS'P[�M��/�Ã�$�3dն�Ls���ٺ5:锾h����r��_1�Z�W/��7�w�����@(ݎ�
��H5Ʉ�4]
���>Y�� �]c����^��#"�^�+�2�6�<q�X;����_�l�E5 �\�m�z�Wn�*�z�����-=���h���%[�{D��{��Ɗ�7��=�t��5˼T��3]n��˭��)(�y�3SP���e���bE+���V���qu���� �Y{���O{�]�D�:��S2���F5�щ�{H���7^�*���C5�:�̒�~.�ToQ疀0Q�
W��cr9܂�˭Π�fj�/�z\��R�&0����f��bW+�X���Y'YL&����a�>|0h^^�4V��W�^&��j\�V;���^Y<��{3�p�a�=��Cq���N�u�Dsޖ��ssاP���W���Iѐ�r�Y�u�p�q|CZg�*��U���pk�f�
�5�|Z�e����]������ɯ*f�y��P��M�����I�j�oD�$�jrT���yZ;�c��b�Y�u���I���6���=��s=��㾼���79n���Smg����DJRl��PxggU�}���=Y!x�Qp��Ψ{�	M �qݹ�r͢b���mu�df8ܨ������$�yy�B�/\����F*�뽷A��ݗ��h�����4�z-��"_U�US�.���;
N��y�NǀȠ�H��:�5e���>
a���U3"YI,j��P��I���[��,�"F�    @
�[m�`��A���@���F
�e�ʕ�h(�b��#"��2���`�QUV"��"��v�Ƴ)EQ@R�,U%�ŬZ��%��b,D�IU��0R*"0��bA���Q
��EPX� �X���AB�*6�aAH��b�EUA[aD(AAb�lTFе(,b6�U-�"�UE%B�H��ذQF��kPKq�Ŋ9IU�J����*���D�Q�iUF[d�Q#i[�E+I�F(����`*��,�BQ��EDP�
Q�����Q+
��I�X�F,UPTH�IF#��H�!Y����X,TRҪ�B�2�B����q�9B��`�k*�%D@X��*V]ie��1i��+��jn�0[��7"�Aj{�����`ͬ�z}��󠛊F�Z�;��NҖ^}�9+.)tg�����Ǘ��^8n�L��R���k�f�|k~�`�t*
��t���Q:�"��ӑ0#�Wd��Gd�U.	�U���7)��u���9�*#=� ʻ����mf���hL��P5��d���Y4(}�[��7z[�!cn�znntu�.O�(��oF*�s�R�F+�o��a�*ֲ�5]�fCY�ɾ�\�0�[9
ݳ���Q����W`j�v�fy�d �ԞL1�)l��=I���2�q�S0�i����m�t��q@����R�#=�������Δd%#�=*x�X O"z�:���e9t7��J�7]�=���f'�ڕ`�xѼ��H��G�ZH#���W*�7 )a�g���Fʆ��o(�̩S��l!�Z��l���PĀu��%]��ӪƴysM�1��u�۽,�����\�RL��R�h9`sȯ�����Bӛ��D�¡���&H��\���W9�6��ۄ#S�c�5W' !�7,,�\/��>�3��H�����-���6f��V�5��G����.�UK��n�j�60X�������1҈Z��݁�ÍoW$0�1Ĳ��5��j��*ީ��`��h{��T�s��f�]^�6�Q\�~,)햌�]b��$���Μ�Ġ��Ԋ�Y�?}_}��}�{���z6%rק�&¸��}�:�"�H����N�NF�@9s����p�]����n��>/��}ln�}��{�e�g~���a�Ř��7��|+&זK�:�U�6F!�,�MW��\s���k4�"|d�gI��k�B�?g�����n�� 6LoWb����t ��C7�f#�p������ڰUL��z�j_�y,�x,$3�X���O���`���v���I;�-��U�i�Y:3ngNŔK@�BXۑ1��"�.���nph���d�)��wc�ܑV���m��W]/>�ݭ!�-��zRk}{����V�6H�}EG�֪#/�Q ��UB�����Yon1q-S���~:dY7�2���{����fV�3���2����\u����2�	�\��h�^��v���n�^J˵Uݼ�����ዂi���$��:y��2���3��}9x�����X�QY��32H��n봎�ԝ*�[0�v�(��ϙ�ji!�]�/g����Yf�+D��,���9��ge:�h�����\����
�5�#,�Y��񠅡�;
̍S��Y���ѝ}4��#�:)��:�h���Ha87�){H�$��p�K���aˑ�x%�K�\��^d׶�����z	=��YHT�z>�>��3d'�9 �q��ͮ1SW���X�n���n�鯂��q��0@�����3�մc����g��7�\F\ƅ��u�U�*95hd9t��f0"i��)Z�����N�D2C�(��O���s�7/~�O=��R=\��F�j2��P�m��3L�z�k�tyVC�0����u�t��}k���z���׶�<��x�7Z�q�O���A��2E)Q[�
P6����V�H!�`u��b��$��0�M�"�����uu�y0����Ksʲ5P�p�Wq\�znO$ai���l�<e��aXn��UB�N�
�GKk��bs��w&t@N���^z�i������&�.!�}���!\�7�ʱ���{N�1!�oޫ'*n����)*d#�C���F��c� �st#��3MOs�P~޴���h���fe��u��r���$%?8U�/�L�@`�i䌥0�!����N��8+f�H����~	^Ԟ�q�:O�_�L,��;�wtn�b7��,��r�}^xm��s)��ʦ��oY#����en��R&�DNV yYhj�6־��/��}���S��e��]�8�u�!��9=V{Sn���!�nf5G:	�3'Iv��}���� ��Ojb:�X�3zsT�ʊ�V�Y�jYU84�uS�I�@�w
��ѱ�z]�x�N�}�}��UV���]�ލ�jo�낽V����4����K��o�U��ȧ���t7���!�4j�=��<��)���q��R�}��J�:(�uN"� ��Pn���r���/�tW:u[wi*NGo��/�޶>����9���6�d�~�#��I�T|w������6}c�w4�ya��<���b8ǽW����\�\��]D*T�*��쎸L�ڕ�f�:�
����W�*����N���)�݆�&ـ2~uHM@��g�7���ICެO��]���f?r�����߄��Wt��:H�pCeC���6�9�p�S��c�.��(Ѓ�s$�7��� ���R�Ѻ�n�1�#�E���A]��&̘O��{[t/ܖi3+�@Q8��QJ��C����cZb�T�33�jv�u�g�!N���L�5&*N̛��#]��4� ]<�����.����F)\l�0��os�X�������6����U��T��GL��*8��q]H8Q/`d�ꑩ�A'�qw���V�ymڊ�� ԕ]]�靎衺(�L7��n�l�f�ɛ����Ls�sڟ�Dl�o��]t��bY������%��nx/c:�k^���bcw��ԝܣGX7ۻ��lPn�:�nw
�q*��$Y�����U^�݊�t�i���tk�P����e������3=�D�`�x�搡�#t�%.��k�/�z��4���wj��[G(ƈ��S9���^t�S����:�TWI�#�'���K���Un����N��e�,�<�ӟT�x�r#fb&��`dJ��&�,�����'w��:3�]C��x|�ҳ�T�Xy9uIA�%�:��gF5�Y2��	��1��}��i�Q��G�Qt=�k�f�����ß
��̨-�3�%�&���i]b���)w��S�-ä"۔�K�����(X�+6����=�C�~�6���v��U��,��TJWbn�dC�0�]��=����j�]���;�Z�ǵ�:ʒL�?A�_jS+TX���J]��!��{D-7�ީ����]�M��wUi�o�I�@�B���	qj���D�2�q�S0�iɩ���J�ĥڛ�<|�u���W�e��:���G>D])�֕<`����oWy/b�[D��x7�{1���|�;;��0X���y[�}Wؾ���R�!�v��kuAZ}��~`OPՔi
��lS�%��J�ʽ�0z=�n�������ח���r^X�u��dg��6��Y%�Ó8WWc:�j�+�XR�3��e�W��� ����� >"�{Vj�UPgd���tf�+����J8��A�P�BG�ɎqW�l䗑0�{��dT^��.�ֆ=�>ʄ��C>rՖp��p��EL�](��3�Oa��NVR�O��
������vt���%q��ԃ��j�1l��R�k���"��S�"8"uJ|U�s���f��a�hZYyQ��v���cj�v������MUɸ��T7,/Սy��қ9LqQ�پzg�T�?(�_�Y�t[��6L��&Ҿ���A�N�N}��\���[��k��)�������]P��VL�b�r�\��n����b���`��@�ޯk�;XCM3�j����V���A嵚i�l�iD�Q���
�,�q'�'�C@�19[�Jܩ������2:�"�\�;�Ս쎭��gN�0e�>|P{\��Z�y��_a�[�3��;w/�)�1|�3#"�w�t��S��Vpwћ��Pə���*Pc�a׬�D���J��2r+] �qwc�ܑ_[���j��ºן6��+/i%��?,��t
��]�7�E��!M�H����QU��e��
�^ǝ����)?Y�9��*�(c���W^��ռ������>Q
��h�/�
��ܦF�u����%9���=L��>��w��֏7ؚ��k}j1������ ��"%w�vc���l���*��0䭎��Q�Į�`�ON�ǵ	�o	4�&RY�I�J��5�Wp��	;S(	���uJţ��%r��r��d�Α�}�U�&���)mGM"��x� ����#�}��Yf�-qW���=I���*f����X��:\W�I҃VC�B:$�7(���>d$ji"��������S���%m�,�q�xEC�\8d:j��sK��w��ð%���*�.*����t:�YGi��$ÝU�m\�p*�W��\��2�D���`D�S�*U8aԒ�m�U:3:��/��B%���0�q'��7�-���1_kF�9L2y�\�i�8uNu��ׁ�{suQ�π�o�O�I�|�]_+SoCϏ[�.��<��zue���s`�[a��H<u�!�打���c�Q&�T<�Q��L�}�륳���װ�<��>�Y���bvr�h��{���z�dk��*�P;p�(֕�pޘ���]X#���pOvU�t���u�p�7��R^��iR'V�K)f��&v�9Y�!��AZ^:�i��J�{�lO�!Hk$ա�Y7,d}�����:�u�0�t�6˗hh���g�%+��4%�Z�qF6Y͛j9�ە��]hPz6�aH`$J��z>�#��uq��h�u�I�����){qڝ!>�?�<vw��7Za;�W�c�q�n!�][w%1Zx�31�_���r�:��C����Bu��3#0���ԋ��uI.D�8oa�]���e��_WVTh$�J�!�'��Hȥ0�6X�[6Ү�k;�����m��y�3�C�9/��w�OI�b����g� �3��P
��Y5�S/��]{FF`s[�c�������2�{�����c�����<<�	h���~j�DEnO?�L^[�7��7�h�\�gD��vˆ�2�)���=9�E.�qu� @�T�o���,{u���`1��FOKѯN=����!�Ч����v�W��1#��I�2��؝nV���4����7�!�Lƣxn�H�R����1��N�s��R�Q(�ͤ�N$�V�=C�B����.���D�����S��Z���N���)����C��`K��MQ(	�׻�:S�����'e� !���A�����?g�[¾��t�d��x���/l��dp-y�k-�uu�>5�ɾ�چѱt�wF��ݠ.�aG�mL�9w�Y���r��b�L�8��,�K��{h1,%s�����W��h�q�K�J����7��d=���wѰ/\�;����5���Y=�t{ﾈ��"������
M��pD)�~�y�5)�� �E3�:JGp�x��5bV���O^��5r����	J9W&ԗ�B��K�Z��2��U��t9�x�+!�i�Y�v�o�KmE�g&�N��V\w:���2c~i;2o��#]¬~�vd��(���O�P���f��W��(\܍��NR[W�uM��N���6���VD��4��Ŭ��pg�Ek��Oy�]�u���i�.��S���{��Z��ݫ/�j�l>j���9�-�ޯ�b�6����+9=���)���|�g��.�zN��̥Ȫ89��ُw��s����*���\���*&>�i���sO\n��yO��U��%Z֖n�S�k�c2�
��w��=����cl��1����뒦�j�E��m6.Z}q+�o�{G3�A�Ds�:�a3����U��Rm@([s�k#���F6:�5��}q/�Y����ǲ�S�~��߰�u�p����e�_fi��`i����v�Ѭ>Av��OK��4���"�
%Wp�I����syr�k/-��[Yٗ8���D0�;�k�r����"�,�����������ϝ��Y�v��2��I����⡓?�>�����m�����Q
�˺��+~�=[����ٽ�{��1��48�ݍ{rsXt�?� �E|8�������٨)<�p��=nО�":Na����f�L���
�|������mo���T9�s�;�aF��x^f����b�F��:W�����Қ̡7��m��u�r�a-��=I嶟�OK�sZ�wCC%J3�ξ��Ϥ�s�	U�x&E`�fME>^��y;=�\��/�������bb9���K
���ڼщ�y���sԴE��L����������}�˄���w�r�(_��^�F�i,N9ؾ���ɪ5�#Q���]K���]�$<��~�c/j��<�sK�����������s��\���z����v:w}��8]"�������m�T.s�fF��.��{���D��a଒�uY���0v��PJ�G��_�n��J̊S�3�Vs�g�E$&"�|��Co����a|v������A��nP�9����(��`�x�����&�u^�k���q�qIB����g,k��!\�Q&o�;q�Z�y̥J�-���(���Jf�N])N��gj���]2���R�D��[Y��r>��B��檀�&|�u���b�<W��Kr��}���l�Ʌ؛R���&"%C�W^������Ob���޻o������@Ǣ�m>����#���%їj��?�g�b�.�*��/�p��9u��:b|�op�M{6�:.�\gy"�uz'S��Đ����^�5*]7Z�oUw;x�Z���VWlm��h�{�-�T�z��Ң�U'h��r��J=���:��ܼ�v�>C���qEY�}�T��8 �7A�;8^�!��x�"�,Z��@I�Rj�c1���)<�K[��񲫾�A����
wF��n�ЛS_.gB���,��7���VK���/��q;/B��'�;k�)�KzŤ-NeSӨ��ȱ}j�Clv�V��
�L�Z�����^��<��K��a�x�	O�vח�{�^4�-�
{��ee4V^����'i�JV��Zn�[��m9J�*�x���oub�Fb�7O�C0���9���'c 0ݘ^��G�o+�,s4Dޝ�Iut)��emE�DhaM4z��cs�v涤ܙò�H���`p"ݓ)�W-�� ��\XYS�ɊL�7�NSHk����f�m�9��Y�lAMk�����P�5)�˥��hg
�k�N���\�6�ą� b����s�T�Z�C/,���ظ32=
���i܉���k�{F�5��)G5�	��܇�&�7�'AvWPϕhr�+.f���Y��8�g$.ݧM�6���9��Y�]���u��Vm
(E��'Y� IJ�Z	�U͡�n�$�$I,�	p���o��F�\W.МW{��6�*J�R������Y/0��۰{#�6��<��n����pɧ��̤�..�����
��I�÷��-3]���gI��Վ�n�.�Z&	�n�H-Nr��T��4���W�.���nE��Ӓ��s��K��r��9K-�6�3T�-ZQGKWN�l�գ��+RR�Z�ަb2��}��2���1}�=OҰ���}A{y�yfc�uY��s{�fJJ��7t��+\"���UcM���@n���`��k����8u۔��#��B�iXٷ}�����{�tDזd����A,�FvbKL�gV�iʽ�t�Ckw�O�D�F%^�3)-��ZW�Y�N������g�Cz���a=�o%ꇋ �y��{m̓��ѫr��;�`�ZVX��M��/����9����|�����
8�J�Pj��ع�kL���|W�
K"��X)�XYl�k"�l�@P"�UL�b�*$Y��0�
�$���
�B�`���kIX�--�j"���\eaR"�F"b�H�-R��q��**ŤD�U�X���V��k"°VJ�b�\	R���A`�PdD�**�"�E*��(*��,+b�r��Y1�DTYYY��`�V�J"�d�b�B�!R�*�b0�(���X9HT���6����ih%)U[hDDAdX ��X�YR�ȫm�*���*
���6���,b"ȤD`�ш�h�Y,��,U� �b�00kU"��e`.!P
��Y�
��Y�H����BEX
TYRb-W�#�f�9��Vv$��DB��Qa庰�W-�����f��%8�����IbIqQ�������3�Ħg ~���>�2�ۦ��K��z���~^�g��ჾR����gUf�*��W�_j��_��N[N�Jl\����H��ᇜ�{ ��� X�2�J3sw�����y]J�K��̹I�q������
߂o�7���mm��	�7J���m���i��ꄮ4�V1�V�{���ϖ�s7�6m�C���ޢ� 6~-�<�j\�뒫�����\\Ձ�)v1�w>��\���q;��oh���06~+����I�b��:�%䰺��������9����m�m����U(w|�
�;��Ғ�1,oC��h��ᘃn��4o4���Z�o�uCb�]��J��~,R����X��sjrG��ڳި�����g5�7��=G-��rj��}�I��5�un 0`�9���[��\o��AhM�B��C^f�»�i�|��*u��a�8i7��zn�Р�����-l8Wv��d�B���v�e}5�6�^aqݷH��V��sC=�ڽW�j�%0���f�k#�.v�Vj� 2�ѫ]��[%uE� K��FގP�x�/Xk���.���Q9�x5/�}��_}7��7:�oR~���Ϻ�ٸ�I���ʎ\�6�21�s��S��4��:�+�NArɞCfN�]��*�?-R���uأ�k�<|=k����#���n5���b5��O����ڭ���Q���0_]�{֖�k��B��A��f�ܝm�'�dc�j�,A�]P3���û;3�Ez5���oz6��o������Ƚ�O��t:�.g���C2j�9�~�ߴ,#<�W/W�e6��h��Fg(�z��e�9	�\�3csG\J蜚�L��圌���ۅϦ�6$��q7�3r�b�%��l��p ��W�%�ơ�1������ �L.�oV�^��.�؃]bz�/�T�ܸ���F��u��}y����TRf9�ul�9:�׀�����^�e8�U9���<e��}q->����v���P`>Y��ߴ�s�n��!�X�{i��w�Q�9�`�B�{���ʺl9�S c�}���t��Y5�˲�^�(����+��x�'ժj#�^�T�6r�%��6r�哒S)o[�Ds7;��!��G��7y19�����X�&�5Ȥ�mkU(�nK��ﾪ��xV��.����e��̮o��=:OE5;��+��*��Yw%<��(k}�����4Ryqc]��s�Y
WI��f�+ 6�scu�N��g�L������f����/��gn|�hh�{��+�MlvsCOl�lٟ�?t%W�-5s�:�o����wM]����k�r��̇9�}Zw7���9�K>T��qԖ�@I�F��T�������˙�-�3�5q�)D����?\�s"`�*��*wƻ��ؤ{7�,w��i{�����_CI�Q	��,����CdZ�6��}�^�� V1/�-\\�s�Dh�~\��U��:5i�5���3��g��,�׸�h^��\��o��P�Te�t�z���^�;�R��8g�#�J���<T()=\#�"��@��gj��U�;4y���e�ru�������t5R��`�y��+ݗ���
�hP��RE�ԋ9�:_u �]>�{ʹ���|���+�86:���$�m"��zS�Շ��y@HA]f�9�W��~���XX@XQ�b;F�����F�g98_Q��W	;����9�n=���Ȓ�����Wae��o8*�F���y<�����t}j������~xeJ��)�j��^�p.�$�;��D=�	|<0�s�\��Q��[�
�UN���CU��%*��ק�@��|�l\KO�"Wf�Θ���H>
��v]����bބ+��C�%87\E���Ҝ%it�6*"�5��i���·;l��{�Ss���.�
L�R�_��JV���ކ���{P�{늫�o6��V��Y�1�y�/�C'��pQP(����*��٨)<�p�މ��\9۪��oo��r�v��R�D
�>~	1ZRV����yۍ��<����]%�wz�=ϛ��b�F����������)��ɝ�"0�%���Ɯ^om�i[9�c;��*Q��9Д�� ��p�VT�۪�����=..�{a����������
�b~�7#�Vtʂ읶i=�:�
�K�`n��f�7����hb��$Dc�]�a�{巐�ce�P����7WQ��L`����Х4v��s&u��o�u�嗨�l��`hU��m����(���2%5��;��mܽٺ��g{h��*����b/\%4�o,��ꪯ�*K�*?P�D���'y���[W���Z.��5	&��]µh	�	�����9�C�`�u\��;�)F��OBj�}i�*�U@��	r���I��c��ʘ}dK]"�����{�
�Q�����ه�`l��8���s��R-p����ڇs:��bE����G��������S����%2	L�:�
��X�LeN���R��c���q�������8��[O�+FcQt��)�]���7ow�g*9ʲ��7���V�Ia&�'v$�j���o�f�&�Ķ���؅�}&��U%Qłf�	�GE`{E\�:�6�MN�KC��m7��SO�6�Ĕ����X��÷��Oo�����N��_��^R��T����v�r]�	mNƚ���t�X��i��oz�P������O�Pr8�[R��Yї��I+a��VD?]�kB�vR�Y[uzhzQ���F�,�̷LK��ؽ�av�CPJMޓ��������
���ӝ'�Vf���⭬�0��xi�
�A�RŽ��pU۳yshQ^-ȗ*k4X�@}�!d� �l~�����c|����f�ѻ�m�kn���[�i(�����������`���n�Oo Vݬn֫���o��k��Ψl\�]_
+��E�ۄ�g!�!`88�!�_|��|��_�ZL^���Cb���K�˫��^�Ͷ����j����[K��}j�\r�4����h���[K6mO���Vê�/B�ʾƖ����oRu�����!�б���Ay�c�ĸ��#9���Q3�l���jn����u�lf�u�Rĉ
�0Ҏl�;7<�=tj"�0k��k�u?k�'�C��å�]�.y��_vi}.g���w-���b��:���U㑵�qY��qk��lL�C��v�����E'��n����u�X���5��u}�3���.��[�S�z.;TU�l`_�Z�������Z.�E���L�E=|���YF�x�<|r�W�/�رK
��X�x(�Ǹ�߅f|F3Ƕ}���!j��J��9�ʎ���<����K���;X�O��N����f�LN�Ktj�B�� ��gUܭM=��ii�`�4K'V%c��˽��]��0�5�}}�|҇,���3,ޡw�z��QՕ�%0���晸��
v&�@=gEe�G��p˄{輘�������3-��_�t�W�֟T�C��O$F��h�T�FR�i�Ȧ�_��5�l^�ʊ@h�`�ڗ#ka���[��CIW>iM�����V5�OYp�|Z{�og��<�U[V�p,+��z��~�j�6'E�컧aWʕM.on�އ��i��m�;MŠA�eʮ��� ���/8֔��*�[�_�\5����~w���w���	�xOk[ﯭ�?�L%����f@[Չ�e�w��>YD�j�=1��6�߫���כL��	C-���3ೖ�N_i�*f';R�n�r�T�㏓c~k"U#<Gy���ڞ�|�ݻ��g�M�n�u�Wx����j|��T�g�-m^?S�}�:�(�Զ�+VpK^<D��]]�4/~Y�L�Y{��k���>\�}̬��t�i���`���u�����T�&��T鋙Z��a���3�W+6�*��;�L�����G�T,��y���&��y �����~�u�y{��[���dǻ���Cθz>�ﾭd�C��1������ֳ���O��I�P��j�>�Dr��'*+I�z��aXX�;�=۹:��U����i�-��s8�	2tw#A]F�)��u�VQ�s��g��V�q���k򗷉�=+*��-|��9k�Y85¹{F��c&󡘪�뒴e�'[��Efٮ.+j��9N�,�E�|��:Q��{��1w�܏b�7XGxtJ�P��<baꉾ���˙�����b�]���[�ٳn�W��e|U�;�)�R�Y�(�vOQ��_T@��I�_-r�6�t�휔qum*�wxV�o���X=u�ru�]](��}nˆ��Ϭ��b�7s����I�6^�TQ�@X[y�������+G7�CV���0�%v�ʛ���sR�f�3z�C�>Q[I+�T���'�fe<�ZTUeU��k����+m�@{x�{��ۼ4�W&��|�9N����_�{)'նh��>��QPnT;��̵�X�w�ۻ�i�)b��}V�	�r��`	�o%bֻ���29�}GMѭ�x��c� M��V%G�sk1+Y�Y����#-��e=z�:.�٣����R�@���邌��)+[[����54&E���m*��ϳAѽ�~�a�F��/��sQ��9}݅�RѰ�o�d�
�[N�%��W��{ݷ�)i[9�1�60����P%%А�{w
���ge��q`3}�J�{�6���\ղ�;x}pW�eM�\+r�Ԑ$�tsI�`����.�P2�.{T�D�[V�:֋O��I�p�b�*�h^<콫s�m�py�9�"~x:A���Ü���O&��㖙6��q��;\���/�5�ǵxe����Y�]�j�̷�S��p2NE>q�t)�5��뭸�ᕍ������� �:�&�W�@��,[�;'��Dk���Rq�\�z��ֲ5����f�P̢��D�"&�:����jV1C��U�k��'춝�M�[��{�Aw�h��m�!�*��^��U�����F��Wl���,��o^������@qE����X�i��^Iz�c�Jx�o���J���Of�">7��?��,�yf����k���>d�K�^6t�A�zFDV�x�k@;�]�hq�~I�	![�S��_|�����9�kuՕ�T5q���L��-��]������
2�Kk�b��޲��]�:�i��ꄯK�lT[M쩔j����s��yr�V���Y=�F�v��O�j=��=��/��ĩWyq�]�$�ͦ�gA�{������->��(t�d�!򯶒{Oco��V�-��q��$���
emM4޾bzվ[f��:{��TH��Dæ�PE�����z͇��cPQ�/
�{��-�k���lV|�u|(ta���zJ���}�}RpwP�)�C;�k�e���׭�ŋ5�]D)wq��q}�yWqtBt#�h�����\�u���}�|ى�}2&���h˫P���D�G�p�����Kf�'�����D,}q�����[�ʹ(��A0�|�
�L�r �W��ݛ�����V��P��p�k�;;��x�XNPi\\����|T�rq5g�;���A+�&»���&�4�m����N]�u�;u�GrSb���!ai��F8q�pG[�&0���e۽FYw�7�sV&˶����h.ݠb9tEK����V鵐P�o���Γ��Z<(ؚ�+S��WNv0S��8��C4���j��CMWu�ӻ�]uG'� �����s��	Cm(�َ�HQ#���yY+G_uL@�����\��4�I��8���L��V��ӑ��Z(slU�E��%Ր�8���ak��i[��Z"�{����{$.�<K��=�Uzni��/����@c~v�^�%(�f,�E���4����w	��ُ���#�4�����5�"��+hw�� ��:�MR��f���]3֪J�P��r	����`Rэfu���s#�Z>�&׻�]`/�a�M�w wϳxS�����4����&��t�G_Rx^"�+���E�L���Èd��81�@VH��]w�^8�h�@7I-�`��]�Z1�S+j6��n����j�̻=�Vl烥cQY#�<]��������>�19��xp��Ӓv�,[{���&�O\��."덎��u�H�!���Rq[δ.�y�&񾂗^S�Q\�[Zr�gd2������̌*#7�gs�8�O:����II��Q�ۂe�Be�����g��PD�2�ʹ��|�Z�]��y���Ǝ�Ʃ��:�fg�ٲD՝ �YƟ^&���t��P!s䃇2d�1w�:;���n9��d�mΩ
9JL����ư2�ؔ�H_q��!���䃂|���
[�ek (U厳�2��PN�E�7��G�������y����[uv�i�.�lKP���U��'+�J�X?�u\���2аV���/uhytIՔ**gq��/�e`ad2ыS�l������`����,��͗�������,��R���f�tLYu��f�&�͹%�9�������B�KYMGB#c[�Zt+Q����m.��(�vsY�(�ة�n��Rq����X�S�ث6e�5L�F�ifԉv��x��5��v��n�Cw��`�7���k��Ԧ��K^���X����J���L�`{���f �.��n�e�L������*V?��C���k���y������m����@Ú�7��6���}�d�rK�������вص��;@nL$�c� �'m
}���;I�En�P{B���[jH��7$z-����M<���a�}�Yץ՛�n��x���E!N��̀6�D6�]w�irr|�"V0�h�k^�ꇛ	�*	R=�� ��כ�ܐ���kZɚ�^���W�V�{)�n`�������wC�)qItX����=j�����o#��a����u����`J���T[��]�p���,��[�2m�х������~&1Ea�<eC�(-j`����̰R��XB�@X,FJ��QJ�T�c� �������W
0L�YZ�����jB�,����I�%��La�Y"Z�j�� X�(�YF�CF)P��IYU �q�c��T�YY%EDU (T,�!*H�
UIF
Ab�X�B�� ,��Ad�mJʈ�"0Y"��(�)(�J�*��VAVJ0h�
���P*A`T�VE��X�h�KZ,�eB��fo�M߱�v��=��b�nѼ�����E"��R��f{7���ya���&N!H�ޝח���%���'�"KG��U|6�E�jm�U�7^��	�5��_Bn5���b5��`��������yZ�����Cr6���{��]X�9:���U�9N���W8i��n�O��% �zXM��y<�m�_nV>e�F'�g������<@tr��n�-�9�e��tf i���3�N[�q
e�9	�]S�0$�&�셙�ڪ���?_Y��C2��|��+nJa^�2��i���}��|���7�߶�zD�̠�	��V�Fө��P���X}n޵ѯ4��G<:�Bi��m���ۇ�?^��@nA�V��=��Lv!��n�II�!�۞�7�cr��k.O��i��og�>��گB�v�O-J��w�E�u�iT�w]a�B�S_.o_�C���my
������d�u��½s���ۃ�`>gBJԆ�%�4Rymc]�>ٞ5~/rz<J�,`�ֳk���[Ĳm���;&��9{�Q��^}��,P��բ�*>|XUW-`�SF i�k����m&�oC�Xk����z�3�6Kx�J�J�i�]�TTr���������.�h��k!u�9:V*5�G��>�9�����c=mP���]0T	h��<�`[��[{q̬�r�P�8��E{�ھ����g�#��	L@`�KE@��2�Ǻ���6��%9�"��s�s[�gp5p�Z�)P�E>�Ů�v����Vs���o^��8{�*�i���l>���&��و�&��ĲY6�:��l�ٸ��z��e�}F�L�Mƻ��c]Z^,{o�꾾J'��]@�»sgSڽ׵��_ܝN��Ԩl�q$1B�U+��^���WY�S�3�yyԹ�}���k��yP8U�O��:Q��ۭ��Q��}Ẽ0ugj��Vh��Y\�ʑ7{8��w��E*�v���z�7�\s����c���s�]�� ns��ņ�"�K�]��G��8��6�pl]�����l�[���fTl�>1ݤ�����SU��2u�J�\�iu���,P�D�jVNQ�j�\ꋁ����Jb6h�ə\����p�%�X 0[xfm9���w
)u�"W�c1��d�y����X�ܽ�5V�ڸ�Y�6����֭ܮʟ�f��g<��Mݥ \�r�;ޫ�����{�-g��h��ϡ�/�ፊ��b�Z}J��}YFҬwF��{2��d��z5<&�ˀ��S���.����O��Pk��oc��=n3e곕\�AJA�QS��¨��\o-�k�q=yG$�5r�+kgy�6K[�EoD�﹁�T�EF�K��:{*%)/465S�v��{s!v8z�<㔥*�P����`$�iI-)�V90# ����ji�V���_r�9��Pع�(�q+�����M������T���c�JA�T-�ۅ-+�g5�gpT41xgw(���{�M����s��'=+�pM��xe%�[/��q�q>��Lvѓ�B|���[�ԃ�U@ۛ��N%�й:�Z.�O��$�}?�WUTܩ�e#}M[REG!�ì����y�/�R�<��當ƍ�8]�,u�v=��V�������$�w3Lz�Ղ�K���刚��X�NL�Ӊ�Uq�'��%�q�']t��K�ѕ�c�����ֺ����l�Wj�u��R�Jkta�^�����H���z^p�hp?"��oQ�ݶ�hiK�Ld����Q���c����(���q��eLk�'����_V�ݿ�W>�f���Sz�m��[�����-8G�F;P�uQ�����1i,�RA�*�I"�-��.%���î7[��+��/VCs�dk��/zͽ�3C���U�0[z:=�{	���˓�fr��ͩM��^-�n�oJ��i��ɗ=������/7d��s������k��晹I�r��Σ�z�㘝 ���Ov�k�wv�{g*)�U����SS��.��n���MWOd>k���x��cKL�"�<�m�t�����ֵ�/��Ff,�sEMЧpʧ�KC�mT�?���zˇ���->�7�_
1�����G�j{��4�$R�te�m,f�T������k����-��1��]���B��UI`��˄u��k�����-�k�!�Φ���W9tI��Ss����'4Y�x�)a��Z�T癇�k:.��4��S]
���w����Cwe�^k��>�u���`juJa�>�}�7cl�w|�.���Ͷ�bQ��dn8Sٔ�籝���C?{l��~���r>���-醵�T]�5��]A^�h%��Et<�j�'�?_�I�9�<�b;���[���;��B�/;`3Q��<cCT���t�G*��4<�kis�V.7��M��n�Sj��t��;�9up��0抈o"~T���9�R������:�ٸ�Iƃ��^*Ns'J�{�D�4�s���pˍj��g����\ܭَ��&�s֤�w8�d����wv�x��.-s���k�u1�Ș�:b�"�QOuy��k���1a'�ۉ�ʷ^r��q���p�[#;��Vn����}[Z��I	�_8���̿���MnV>e�F'�g��t�St*�A�LbY�Ҟ+k���7_43(󑘫�6���e�(������X��mMwR��;�zs�ZO�[�c}NY=U�H|�rwd��q�*�ƅڌj5jS[1��N&�˵�-�͘��9T��F]���W=%!�	�C���W�P\��s���\W١�=�Ҋ�u�����B���g�)��ƛFUs�6�E�ѥ�úK���ӊM�̦4m�/PI3z27%�4ag�`us����0]��r�N־WR.U��0��gU�В���.zԫ$����[�j��R��t^�OB�����M���ٷ^�U{g�j=懨ߥ��Gt�5���P̍��눺���S
�:V5�QX�z���of;l�A�[�G��ĳr���َގ�@���vOK���D*U4��|��c���3��:(�ΐi�y��R��b�K@pq_�kJJ�Pu-�)<�����Qq���3|��آ��V)�}Q�K���%��O5���'�eU�df{�? lDr: n>�Gh�F�K
���߮^V6��pa��5���r����J��m���d)F��9�@����kU�lO:�SSp�hnl����0ӧ�2��j|�8õ�~R�����nL�E�]ՐҋW��+���sN5�z�֦]|�Q�i0Sq��GwU]����$�d��*�9�C����U�Tw�#U�yr^&hi�s����;o��V�*Z2���,��]v�Z�я�w1I��By�iq��>��t��c;��,��<���d^�B,#t�yh#Dnˀ#�|�T�6@���\�oUj���4���g6��O[��|yC���3@�瀔6��|]�(�խӡW���P���_o�;�fbH�2;Юe��1��kh�7Ċ}����.>guj�g�	=��:�%s��W���C���vo��_>�gVh��Y�Zf��aA�Y��ۙ�{I�9���|�9꾎�7\�es��(?+��HHEљ��eP]s���+C��b/�qpRl\�[p�޾͘�g+�c0���"'��Y��\J\@)�*��5х�}&�i�D�͵������e��Ȋy�f�죎+ڂ�A�_mK������u���7���K�\��M%j��f�~{e�06b
p9\mOK�����J��os{�О��E��jc�E{�/zx���U��h��7��*�UR�S}���	��3R�;�����p�WХ*�P����G���W��`�m�������kf�������_u�8�[��nQ�#�}�� @M�5U��'s���:Jנ�{���׹*�{ͅJ�w�ܭ��K��`W�vp���k1��m���E�|��q�ޘ��GJPf�ݨ�Y
y�u�6��U拖KIڶouD��Ʈ���}VR]����F�Htz�)�:�j�1��9b�Ն�7��[Է�n���֘�������r�D�F����9y�T6��y��A�Ϧ��s�	�{�*歗��3�,��5q���"'*w���y��:a� �P6�s�8�ծN�֋�O���M��-cn���Nu����ƧI��(ms+wrw��hvP.zD ��Ƚ��U��AXn�8z�է�n5���ᗴ�o~�g��K��e�����vM����{W����v/$�����'[��<���F�Y��A���)�&P�3��kh$($J�*�q��nW;*^���Z�t:�����e�]Z�<�а�.Q��������9D�[NԦ��o�C���z,��O�0O�M�ˀ�O�̢�,��+n>�����o�f�&ł�Q�{�
=�3���W�І�A�AW ��s9:�-R�F�]��A�vP%R8�k�R$L����V�SY����V���)��/j֮CD�Ѯ|d�V����A��PHl�~�݊�f���<akG\,:O�s�T0qYZ�����[�{"s�`�1�I�����|e���%���$��S�����;�zpJ-&�"�}k��z���Q�*�ּ���!sL���M��7y��o.���z�\�����@�܀܂���u�0f��y�o����N��|���������-�iT
�6���׵\o����%��	��k�o�D�.ƻ>|3�i ���}
z�o�\�3�,P�wLZ.4�Y������ZW�w�[ѽ�(��)W��q7��?)Fx�t!)�h'������oR��6�]sgT��U8��+g�k"~T���y#�7�뜚�f_���կxdbƈ]c��#m>f�|�.5��R��6q�4#�$AQ"l��P�'�=/+�f�Z��S�p��k�=	��j�~�dt����3��K�Z���2|�}Q:�����]X�9:��ᕌ�ߝ�3���w����l��O;��k�mS���ޙ��j׶j����цe��'D�Əc�s%b���N�yd[����)�zG(� v� ��$�VF��G� Y,��;7_��8���t��.��xẆs���/+ܱh��p���qǲ��g8�����%�u�ZE���c�2�.'���Sܛ{���|Ӯ*
ٓ�v���S��ӓmBW85��e훬c2�9���ہ+F\g(�|����6�)��vR��+Qq	�W�v�6bݛ�.­��t��Ĕ�eZ�C|}���a�Y��=���3$D�[q-�{H<��`�JĻ+p��C���=.o!;�.alTsM�So�_f���9_RaW.:*�I�ґ��]�q�\�J��D�
��p5�_<e�i��O���Qq��fxf��QΊ:�0v|�jz\��L��7��ǡ��Ƙ:e��Y�9LM�5k�B��aPGs5�%b���oMAI���F᭧S]���z��k��O�ʕ�(r��Q�-9�෺w��+bl��=�+�.�n�����8�[���r��?(JC �����/*���!�ۗlG��e�89��O��t�
�v��X����M���@x�>'�`z�"��ި!���;o���*����'�<.�Mi�_��,�U#\m���a���;����i��9�@�+�y��n��������M<�e��E�e����VT��RKշ6�jB��<{�H3`+Q5�鑌�ؕ�C8��.�t}u��u��\�6sQy�}S���#�����b�'|1i���𳳸��}P��77kd�dӺ���PQ����|�[ǍL��_R>]�^ZC�h�k�wݴ�2{����xv�
]G�7��V5�������ssgV�`���y�c*d ��Jh�z^�dd�6��Vi�r��PB��Z66���U{��s�b��{ ���D���q�M��j39hC������Bһ�ׁ0=6pR�������f?��*-��We6	�!��6,b=˫f�-#8�B@�a:y��gA+&L�ԇ;�t�81�c2�nk]�9/Q"��l�J�6��']:(��y��2��/�u��X��XŞ!ԭ�3u��5mi�/��^� t�|�SfY��c��)��j������΂.G�*���G��xZ2]CqصD�.�g7E�}V�S��hE�X��\�!K�}��D�(nP���$ݙB�k�3�+\��ߑ��K���52�R��*��%}�`�n_+N,�-��`�$�ĎlO�,^���wc�|��3T�EK�����nD�4���a��Fֶ��ѥ�[*�z���6�Њ᮶��:p�݃��)Φ$�ݹ*����.�r)+:h�N �;�a��/Y���<�����zT-.�����b��IS�|�^#�wȽ�r�l��a�	���:I��in�s�c����B���߰h76e�Ȫ��L�X �ќD��7��p��؊5pn�1��������$�,pz�g8.�F���$#�_�*�.���#����X늧K���)S
ژܡ�oefr��y�f}��]�xv�Z{}.� a/v�6Z�s^`Sa�s#4r�y�{�Q��Z�ev�����.*���1;r����ʽ�J���]R���re�h��V)Ví�b8]<T��fh����H����݈-�؃`,#�Ի��������A�8k/,��&Pd֋ˎ���6���ǁ�b��䷔�fv���x�qU
�L��5�eZ�.yƭ��ٔ����"�ޣ�h'���K<��vf�u �tWnE���32�\�u�"k�º���qJ���w�I5�)t�)Q0�wp\]ڜ�{b�olnX��t���y��/n	�q':���[����A�p�q�M"�yq���6��j\,d&���������s�AB�.l/`�:pG�צQ��g�]��c$��s�Nc�g���px��yWڅ˕t�ԡ��.d_s�s�܂}��n�N�����*�wW�u���aDJ�Qd�VTZԬ�%T��FҲ�J�¢���J�E" ��ȱIY�b�Z֖�T��*�b2�%`�VB��+*�$��i�"ĩ+ �
ZZ���d�b��4�Z��ȵ���0kj�"�
�XQ��Z"°���R1�T��F
4j�R6��0�ep����b&V���X"(#b��
��VT�b�Uh��8�RE����@D��La�	��嘐ĕ�"��Kd
�TXR��
��VKm��°�X+mBV ��H�c�(�X*�
őkmZ��3?k�u��:��=�_�Z�W�v��.����jwq���Yt{&��>'�c��`��h�iV)��z����bɻ����W��n*��2�&����w5�0��	I�QפrYq���X3���,7�7�=�I���ʄ����gw ��=cadvɬ�y}���O�yP˘��Ss�m_ѩmF�]'�k��q�rUո��kR�k��'Xw.^��\v4����/.�N0}��eLa�e�f���S���1%��i��1�[P38�ҵ�繕N6wZ����FTf�
��oe����*��ci��W�؆H�u1Q�}��=��~�>�}��ys��%!�̙ŷ�s�����#u�fT{���;p��9ek��С���ҿ��aQ7�8	6��kk7�6�����%Nn����p�8N��-W�N��v��lW�&�Ĵ���L�[���X�+t��e�����Aղ\�ꄯ�.�����W�u&�;��R^C�q�+U�X
�e]r��z
�{Y4���9+1*XsI˶2;p� \i>^��p���Uh=\�����Gl�QY�^'Y�|ɖ�_L���H�HK1Er�w���ښl;�J�A�1˩���%7`R��D�l�Vs)��>��{��%9�yWѵ=.�*��(��=��V�%�˾�r����{o�X?����7�P(t���*���I8}���#�C{��p�
FV��ŷ��P�-��r��B�O|�k%9�x���E8���s��d���}h�{[֩����}��ί�?C�g��gL᫝������\5��!u���f|�-��Rҿ��k!��M��
�>�Vk[���(���ʆ��M}Թ��C�\�����図�ux�UJ�	��Vc�G� �F'��6;�m���'����E�GE����]����t�*������Z�䎎Cd����Ӽ��i�"Ъ�#׉��s��k�MI�����T�'���������u�
��~ɶ�����~U{Y��N�ָr���w3���9��|G.8\�Qvn>3������}�6Gp�1f���������vqv�1��c�k���Y�����}��'P�DJbზZ�fvW+��^�$Q3����О��v��>m��x��*���wq�R3p�R�KN.�I��;m��R�p���2\��rn�^���N�r�ڙz���]���ݠ���Q�j�	����e��{ f:3u�s��'-��l)x���u۷3SR�$�\_YʎC2�
��>]9:B����i���W:O%;7ӻ�fWh~�x��g���B�[A;/�VAV���SS��<���ʤ��{f�y�7��i�����\A���9QH�<�\����j�B��T��=8�.J�n����ކ���|Z{�މq��\VR��p�)M���7��X>��ؓ�P�ԾO:��y�<��*�ҵ6�ڪ��s�t�?�����Ғ�8�[�P}�G��g�;/k���|Q�<[.{�WT�9�P(l���-y��Gyk��-'��9ú�]̷�qN�>���#��T61�o��B�{5K��Z��%��d����d��Z��smva�o\	3�%K�WcZ�.���|M໙V�ɾ�Vyv����u��$<sdE��	u�\v��)��>n��9gv�W7(�v��h��-`�Y�#4[0l�s����9�JJ'0sU�Yr#��nD�f��˹D��H�����4ͱ_5�*�����h��K�Qk���j'���E��3��r���Z��\�6�;�\k��A�R���6ANÇ���v��	�ͭ���{7�mjz������N�����z�e�2x*;��z�B�cm��n�N�uq��t���'��Y�F���t�����ڜ߾�cal}_@�U�q<�n�j7+�9|I��5��
Y41x�k�8�{����|e����dά��>�����^:f��efc��U��'2�����u�q���]�A��2���<z+�L�7D��}ٚ�KW9����z&-��Ĥؿ��֖oGf�휨�Ta�el�u��c,k��㸜��q��Tԧ	^�
�b���"�}r�6�t��ϸ'n�f�=wX�t%$
f���Fԩ:����\l<_Ci��KO�9����VD���f�ǽ^[���J�l�M:]���G�NN����m��aQ�Ç�8�����hOۅ�&�����_/<�j.�����-�<��w���^��4�뗐!�'�ǥ��E��|z����v+�m�f���Ց��'r�B;juJ�s�`�ar�=/~����J��s{k����x�4�� �o�gy�6K[�l�Q#�9���_w3q�%b��zA'��nv�Rr�۴���ۙk���gS�h�υ���*KE}���1�\��ۛ��RRp���i�y�Y}��8�s��Cb��3GL(J̤�-��H�Rit"��<��VC����I�p�kle���&#<G0d�����1�<���	�Ɨ�(5/�ڟ�}�D�I��P�3M�����y��C�.�2�k~��=�K��^)����6/h�2*�ԷS-=���)C[}�j��o.�0�OGW\8j��CdZ�uq��w"u5�/.�8�ui���X���~����\}��6��\�1�[_Ψ2��?=������~�Ѷ>�/�YG��r���V:���7X�H�u1[.΍�x������Ԕ[ٻ)�#پŜr �O��^����J�X�էxR+0�x�Gz��KT�i`s��úZ�Ӣ;�9�yW�`���혮�r�D�LP�h,�f�le���,�Bی��z����b�V��2$���Epj�8s�))E{�N��s6Tj�J���%�یm�O>�2�o��t6�y1�F��G_���б��x��ޅd��ћ����v�8�)6.%��mo[*�.��������ߠs�n�W�U�ײ�6J��0��ئ�b�ְ�zݣkGq[�Y~;{�`�o\s�:�#j\�P�F�J1���-v_@���#��X���ڽ)�uix�y���Y�U�g��j3���/m>�:�Զ�g^-�dvmL�?�o<����zt6�ٽ�:y�A�>P.Y��v�e��=��O�n�<�
���k��p�(z�<�
R�C�;�ٹ9E7
��wp:�f��1`CZ嵽*}5��h�5�XO�z��f�Jֲ��L��=[����t�EF��d�P��Qi1x���2	�[�X�i��9��G*�KT4}7K��M�=��.hG�+�=W���3�!�އCQy�< K���H�1�7e�54���O�a��c���?������}Ee
�����p5�1���v[�[��m^#���W�Q��Z>��dsS���Ⱥ�Ӷ�Y���sot����d�q[T����w5��2<w�g�K
�<ib��ـy�ۛ��n'ڸ\�\rnFIpoNVT�|��7%>�F�m0��Ь�DLr?@+a��r�vՖ5�B=�M���d�C<�%��q�pr���n5�ʘ�ds�-i�s 9s����N��97Mmή]�w=����I�r�W���X��J�Y�i%������=���i	�M��S6���|:�S���)��>ny�r4U��Qpլ���j�qlמ\Ǩ�� ���/�����E����E=�+멎����:�r���~��lKA$��	�ڸ�><���e}3x�9hLfF,�ܥ֘�H��M�m�Į�W�{g*)�U�:��S��=,�:�V�ҫ�ދק�_��{-=R���q���o�u��cJB�Y�pVT���ܕX�+�_�CY=O�"Z}ޯ����LvZ�����h�ܱuW#�Wm��jLY����Z�̠�hґ�2�We�#��"�ػީq�ͫ�B���|G�pEI�S�߮,��Q���7
�V>��D}K��$���JxBi�� 
F�v�"b!���guD�n��AӧSO�ۇ���z��Z(�[1�VL��3M�P�j������]%��w3ZRW�*�K|j}�[Z�Ż���ő��ۮ(���)]:��������f#�Q�����N<W[3��D��y�e�Ub���ECc&!�3�r�	F��gv�=�ɠ+{K�./����g�?�8g&�5�6m�����R3�8	X�3�˘za�Z6N��g���S���7ӭh�}˙��l��k L�1�u80�on�:�Gr��V8��n{�o��n5-���\Z�
n1�RpBu��3�u˾�*5̢V�"�j��ۛ:��]X��N��8e)|��8lLåS�������c��#�b��#\v�RS�T�VEB.6���*�es�k�]�˙�vn�ʃ�F�f�!W�Y>
���;��q�TE"��/_�����R�����@۴U-Ҧ7��z(�M�;�r���*ئ�
6h/��`�D�������R��/�S��L�}�ۤӻ�5-/�9��L.^f`N�M��䙚���N�㵔�\+G�đ�F�-H"Cu�{�Jx{w�a�������1n��!�C�dNiUҡ�ΛF�B랢;x\M�L���ciou���ʤ@�	��5ۅrݧ�PE��B����\5ip��-���or�}r�5�M�nһ:]R��J�p��9���*V�s�N���c[W��}؅�n�zh.���Eڵ&�
���.��%A�>US��+�*�J�sxg���3$,A"�n���N�^����ޞB�zu����O�A��֔��*0�l���7W��ZB��fh���<�o��:���S�c��ܨ�4$�xm[��4�m���1���񯜾���}��ld�9Fx���%@ee1�ێ
�Y�t����&�ί��ʄ�L^���wG�������,5*��^�CA���I�8$�𽆹�m�v�0įR���r�ww�������F���j����h�����9�:u���#��-7<zl�CX-.���v��O���׻�<^W�o�]��FZ��u/-.�#��βk���3@hS��
PY�k}��e�i��˝�&<�M��ϕ-O3�m��W1֨q��q��n�2�t��@뛕�nq-��KkS.�O��g2��CU>e��T΃ �]���A�tD�"�����+�s����^"7�dZo�w#y�&�2�69�u��ޏw���c� �ޯ��Y4*5�H5���@8�K�
�����\�{���Dq{?�Uu{Q�|�����{~��J�~�=.s�t��*=CT�q�6Q��:AЧ*��ZE�m�]J������rJ�x�ڡ�#.vC�0���q�䁷�YCO����Vwz�~�ܶ;<�<�9��ʁ����U�tIrʕ2���� �^���{>���,b��>�ȳb����Yk�/՗�Q���S�ߏ�wA�/ ��_���r��5�o����~��|p6��T����ݼڿ<�L+O׆�w�/�e)�Yd��|g����Q��@7�}v!����F��سώ�tJdz1D����=����f/�s�D�$�B2�2���*>�l� �'
�c+�|���������::Ag��I���C�茮
�%TB�	RC}�K��5���_-�`?*���8nm���iSÏiVe�� ډ��[�<Ø�;��S�/�w!��I�5�7K��in�3�g���D�.
W]v�j�0���U6�ɕ�oV*&����3��ŷ��Qk=b�� �\ӭ�%���ד^m1R���w�oL�,|x����:k��5 ŋ4)���[2q��lU���w�����sJ���2�d�Z��)�sf����U����.J����ik�Ӗ��:����O�m���!�N]�}�>���ީ�u���v��)+5ԙ�v�2�Cf�p�2�D�o#�s+� ����b�=�E+}��#�懮d~яa��!��U,�n6�K�3���f*T��ڲ�i.�f���� ue��]�<9����э�='�<�"���hK6m�s�7�#�9,�'�i����'	��14_2~���j�Bt�����v����s�
xz��T�j��
�u�|�j5�"3���$����&M��C�d�?�e��w�h�7F�%ҏ#v�8͙s��0�s�2�r�(�Y3ky3�^��V����P�ZUm�]��S����,��Z��DՑU[q�\2��zR�v��'�ˀCA]�\���&��}�| ���ݫ�LAKWJ�����ʺ���I.�w�,��!�Nrtp�S��t�alڣw��o��}t��&֎�Ywu0���q�C6��zvD֭��e����5�׆�S�3��&�跹t�!˃]d�����1"a٧t���[0][��;ޣ���g7��<��{�������%4ʸ���4��`��x��[�na�5��՛z�j44�;ä%��tXݺ��S�ރ�Yr�6��s�v7��B��gc��͔�xIr˔o��V��!��(-�E�U�)��V�t�YZv�|�co��gسo�́ir�t���<N.ehY��"�K��)���r��r�R]�e�0<�N}:c�p��˄i��-��*�,��C�������Gz��fb�s��I�b�<��8���g�"���ۯ=CΎ�L"���V�&��{��_G3��,\�X�aE����z�-��3�ڰ+.[�����X�mA-�/cesR�^�w�Pw&��T�Y���t�j��xwnLck��ЭE��Sd؛�3�gon�g�'�:b-:Gd㵏���N�� ���[:'�^�=��FvS�9���=�j�T	]k�b.�Wuذ7{��[;CA�g�P	��'k�vu�;&�W�����]����C�[>e�K;�C�	�gvrH�t�JRS��]�<�����^���)�qVm�5�l���1q�b�V^�x-��6��)�H��v곯PV�
�l|p���.��.s|�Z�e��d4�nX�˗��$���o���gS2�6�2�fvLxs��g<�c�(i��@k�P�JȲ[dm�`�m��Td\T��XZ��T���V((�E$H���VJ±B �`�QBT[iP��V��RڰU�,Ĭ)�)���T�	RT��ڰ��Y
�"�TVDE
�,����
�d�X�օk%E��J�UPS��Ղ%[J�h�[jʣR�mh�Q%kօ�*�KdP��*J�k[aZ���iT�Pc[j�Z�el�(�b0kEh�RcT��KK 6��Ʊq-����(Q���-�`��d�ʋ
��,�����AB���őB�@D}��6g���߼��Vk�,]IGE�ev��v� l�%�m]����%��7)!"Ҷ�k֕º��m}����^
������`���˥Ō�]����*���^����K=�U#:�.���ͅY;#1��~����S��I������Y��Z�)9�"��;��h����sSkW�1;����b���@J�������E�K�3��W���ϝ0�ӽ~g��Ͻ�_�.jl�O�^��T����{ ,r�!0t�P;��c>��To�W-v�xz��+#A���债��z�ݜp�#'\��jd�3�=>�w T)d�@2��쨨����2���8�,��Y|?6�Q˸��W�-fx'�R}�n�����C���Ԃ�'����x�=;x�x�Vx���.��-��hfGa���C�Ϧ`�8�^���|��WdɨS�Q�ݯT����xb����2���\xdWy_�Z]������+#~�&�[����Fv2^�7R:��a�cvyq�/�<K^��+����Ug���n�+;��_m��u^�c}����^�7&�ɿt5s�X�XCو��d�`09�E��L*Sfǁ΍V���~�Lcˌ�g*�Y&=���|�)�Z��7��88F��ܯ��vC˼[Wdܷq�w� �s�Y��������y���/����IYH����Ml':�ps�-��J[�ޚ�tH3��/�����k��a�cJ_'tw��")V^ ��^/0eN#��z�o��g�zb,������Q_�v�K���=�~�c޼]�ۆ�`F.~�����M?=1���ֳ��Ȩ7"c�zdA�(�!ѶҮ���D��A��:���Fs5��GW��Lӎe��%��v����¡t�nI=�'�P�X3W�
{�&�g��z��UK:��hw��s�t���_�8�;� o��`yE�>��(J����rA�xE�����5��_��y:������,�n޷.�U��D�,u�b���h( yQ����Gۜu:=�BE�>��^�8ٌ�VD�{�O{���*:v[@�C��郥q���0�#�a72�^�3Q���f�ͧ�b�gc�Q�2�9���{��X�_����e�>��NbiL�. ����1+��w���Y>��sE︒�3��Q����*6�o�����,�)?�����lq/��٨���0jGaF���Q��#�X��-G3h�ts3��?ol�-����à;��@f\̏N��C.|H:�ʬU^�ŗ�m�'HzK7薷{}j��� �O8nĽ歆�S�>IE�-T'�6�x�&�Z���X��@���<������j[t��Ժeϥ:B�K�F�nV�b��+�t7Q�(�i5�r�L�p9�z��0�5s)n��/w�BԨ�W�6to�4\���o��W�V��QZ�
�\��*�r�9��{Ϧ`��\�/��7�=AD�xL����s�$}���I��^�ɇ��ab��]|2+�/���j�C�~��e��;��s��^5.g�Ƌ��7T\G�w3gC'�d�V'tù�^��N�=��lxr��9U�{�48s���7�^G"5����M�n�y}��z��&��k7�C�K»���k=t7j�(S���%�� {s��1�W�̿Lw��^��ݓ��nM�,;q/�\J����v�[�{Ѿ��Z�f�F�x��1�����c:O}��|r�}�^:/N�^�������=��NWx��L��>���S\�y�t��v,��u�2���᳴�ȼsaT���ȕ}�1J�~TcОT��Z�ǲ�,\u�z��:,���q��=��6�����.�[ܪ���߶K�2�̐��VK��$��� ��LuL���Zʂ���?����s�7�.���'�GtK�t�<mw���hpD��2N�08{ڧ�r:e���b�{ڮ���� b;��h^ej���o�C����>3{w�A�h�gOSv��J�8����F���a��1�ː���]�Z/z�3��d�q�h��&�^M��\���P2G���jp��:�M&�n���
�}=��;Gw}��&���!�w�9��י^RFq_yIN��eM2 �rʇ�y�۹>��)����n��^��{"%�;��E��l7�<d{�F�ޚfj�(�E ����y+p��Q���>�'�J���H���s���*6���c#ӽ~��L��q�Z�� 2�{��7�K�dz.d�M���㤌�u�he'O�l,z�ܬ��U�0����b�/h��z�Vb���qZ7;�e�Bǣ�D4�8�5��E
]��ϫ]>7�鎸����Vb�Yc蹺}��u�rW�{媙�����w��c�u>(lq8��@�2����1����w�����pTz;g�7�r{�`����O�RTc� ������Y4*5�H5,�P8;��4�3�	~��#B���8�a�=�齬�<�W��k��s�o�����gzrN^�K:4�vH=���q�P�@r�ҕK�EC�pн�g-jG(OA��+�����7��?O��6����X�3G�܎��K�:Z?_ɼ����+R���< ϥ�_�ϫՌ�^��>�غc�3�	�L������\
J*��T=����W���3���z���h}�+����^z��}Ns�u���=���s�ԓ�,��;��$���(Kם�<b	O�"k&�]0�(�55w�i���ӠkUa��%�b��:��n�*�Žʈ�CNs�z1�N��Y;��x�C��\{�@y��W�����楛�tj�.��T����W����ɳ�徼4^��)E��%����S�U�3�@nzqߦ��:^���}��y��>�LC�t�~{A9�?mE,�r�i�'�8Py�j��bJ}��zT���Ǻ�>F؛�����5â�v��$������� �*��J��}�{�VP����K;' ���wG��~늹n���x�>�Y�gT�ni�Ev�VWn{�I#U�����0t�6є&
�x�2�c]r9�Rq�ZF�Rңޓ�)��(�W���/!Ү}}���ȯL�4���|]?Io���u�w`9��89�q�)��G���g�4�z���6M�/��6P��F��.��wO�	�J���Z>����۱B��;������ER�}>u��A�ZK����߽y���O:	���N���2��]��v��V�M��R�do���{5'�mׁ�@�x��X�dY<;�2����g5��t{�1��u�ʘ���`�Be .�^V�/���{"�&�oHyz�|�x�L���1���dT��.�ɕm����Ʈ2y���n	� vR�[&�-ȶ*t-Y�N�}�O�z���������s9ٝȁ���ܥ���%b̾CCcʱ�q��^=g#�_���|����?PM�{ޠ;�*���L�����]��sy����A��Q����q�K;e��.�}Y7#{�VF��G�[���a�S�<%,��,㮼����p�x��_@�a\�fs��t�]�ǟݶ�<1�{��������-j�{U��p�u`cS�>�VB�z�Q��������	�,_�YW�*Ux�L u��1M��M�u�����v��񠚾8�/U�s³�S��d��*�j���ʤ�sjW��=vw�o�� W��?d��/ޓ>�qT�h�ó�$�O���יu�>�/L����z� �9����Ṇ!t1��C!̎ᓿS�e�r�ϫ����ܜ�U�κ���}8�gh�]%�o�8=B]C���R�Bʩfo�O�c�G^Ag����v �,fIPz��NzE�����J~3�E�>9 ��뛿u'���O�1��C��پ�]-ް�l�v�U����38O��,5��3�0�G<��`�2/�[s��G�W�hH}>f˿���iEQۀ10S��15%�#�Q�G]�B���u7u�Ɵ����1�hxZ[t�Z2/�i��	V){do>go��gy��JjW7q�]�_h��@�s�a��h�_E(X�i����N9؄,��q��:�-�+��1�;�Ő�����y�i��z����@�@5�l�郥��ۨ�$@���Dk=k	�$UIe�CA�\M����^v�}���������#k�W�&�S%K��@l�$,�xV��W�m���+���Q�F\���_�vo���{���h8��d>W� :'�/�8����q�A/����U�+���e����~��]��<��3Q������㞟P�8n�t�`F���o�Uֹ�S2=e�H'����{>����9v�9�\�f����)`�����̗��=ݜ�#��
���'�'�2a���.:�_�t�o;�í��.��sӬLs���7�\��ޅ�B�^�7�@����B��N�,�T�j�N�q5��9�H�����Ux;�%������#����������^/c�V
7�4+��q����ʁ��]`1>���FX��`���$�Y4}�tny_���k�P�P��>^����\3���|���gr7xAfH���/Pޅ>�,� �t��
#�<k�qyV���GY�c��o�̊�|�Y.7�#�,�@���kkѭ^�Q�:�1v��U2��gG"�#ѩX�=z.�5�fYŅ�D=W:���73C����Ef�v7Ē�Zu9,u�\� ��XCC�����M�i��NS���I.����e�6�tr7$�0)�▷��с+١+��-{���W��;ixc	p���^�����9�����r�z}~�x�uԘn��s����+���Ӝ����v��Pt�c�g�v��f�_���ޯ�'�|�d��l7���ý��{�dW�ǖ|g8�|�*Q����2�|�����^��YP_
b���ή��*:���f��P�!�x��O��y�����CK$�{v�8�E�U>ۊ3�oލ���o�ɐx�o$D��f��י[TF�~RFTC�a\eM2 ��q��+�v������:L`���x�3�~�3L���s�hl���Y�?����.1��zȞl�O0O]e^�P|��范̎$\�Wc�����;7�\��=�Pqy-�#=����E�k� �s�%��h��2%31�p6����1"�-9���{�F��+r`����¹~��y�;B��Ǆ�8}�7��|б��D��������*;��k���9�>���f�c.�җ�f����w#�ό����w�!� '�u ��8�^��K���9�DE�̗>����o�r�=�.�\�i���iƊ/T��N�H�=�|�:Yԟ$%	ZiKy��ΏS��U�T*�)��,��n0�����,�,>�?�Ÿ]
��w#�8sc/�i����'Q�c<��!S���ۛp���̸6��۫�]<U^��䭎��c�\���7��6�hV���e���X���n�.��99Ø��,��c��;�S�7�{~��N?HT�#}���u�*H�
}��V/M�1,���=�G�/�R��4
�����d���Bxzg��2J�酕��>�%/^׻��?~za�3���9�2�P��fg(�ڕ_��ٖ/;�D���*��5���󃵑��ŭbzuk���Ыx�cʝ7��ݸ�,d����|s�@y��k�c[�p:f.3^��u�ӂ���k��Ms;Ar�^z����Y���/d|g����QGj����\sG��q>�ؙ���V<;3��,�'�)�|n�i���!��'+�|�*Q���<j$��׽�U� Ǟ꜂�v'ɋT��Zr��wL��kN�|�=tI��?7���{px�;|��Y	P��z���ߘ�& ��*@_]?3]��~늿�;��^����O�_�\��w�2=�`Hw;��ܹ����`�A*3�%��7�[,d>��r!ߩ
��z�1�wָ���\�NQ�����A�뙯���Kܱͬ�n�Y��έ�i_,��f�PS\�����Zs�,V�ɋr=�΀c;��]���VL�55�+Wf�.�J�y���]�|=w�C���ヸ�5:�Be�H�K
��ޗd_-e5��u-���M�W[4�攮�س�~}Y����J5����Q%��8��8�x'ʐ�}�wުg"���S�̒�>d[��n#,�|���.B�KGu�0�F���َ��]�F�L�ydHի�%c��f�#���c�҉��˟˩)d�@2��ӷ'�|��2�dg�c�gʏ�e�ב�p�n;�׃�ڟ��^ w�!։���A�,�2ΒrQhz3v��Jǯ|���>�INa����43#��;A�>��\���-���n�޷���Z�+=�k&������O���PrP��ao]><2"���:�<3Y7#k���;M8'����]5=�w0q�T����dYd��C
�Άfs����'���>�YpW��G�:��g�WV���<��z�v���1kw&4=g�0�M�Q���`�	���q��`�^뎺Q���s��dG���}^�g�顚{�xV{*t�ɪ�' /P蛻~å�;Z�M{�O��EN��k�
��쑑N_�'+���r���=��9'h�|�}^=�!¯�u
��&�G�1��(�o?fe�B���Ѱf�p�q�9
�9`2���)9@}���!͎� Xƕuyד��o�s��4�����ܞ����=�}�DEOQ�W&�nDf��G�Z��x~Ȭ��<����3�S�pK!��;���B	:#A�]�"��cj��Ne��)v9;i�UE
b��E[��w>_s�j�F�WwP�b T[\�7��O���Ȟ�
]c�f^ʹ;`�V�W�fU�@�M�����k͏wպ��Wy�3�{�1�ܘ;;x���⢍�هpӖ++@��n��9Sp-���YC3�]����ro��x����<X)��(�?U~-Ι�W��:Wț�M[h�]��}�9�)0�^��\�C�J�u���U�i^}�g�+�w)f�̊7���
}c�D� ��e�^�v�qbǖ�P;��1L�NZS2�>��5Ң8*}��K2��Ȏ���v�e�mVeZA���5�9/p�6���ᒀ�꿏�9�<m�V��4]l��r��)B��`sŌ�	�[[uw��Z�{��6�������/(#N��fƜ�VV�>q��.�1c�֩�Dץj*���E�|��1'�-G39��}�:���r�/b�&�$Tg��Bj�[ǚ={b��}A��d=CE��4	���I}��s/7	�g@�")]'-�Zv��e7��(�!ힽcX���w�Iz���lQ�)�%�����5�-�V�6�n��m��qS���ݮkD�p�"�J�l�lU#r�pi�׆�6. q�oTĦ�u��umu�����W��Y�q"�\��Q�ɥ�.�^7!v�����>�Vr��|yʆ�M�7���|qs�F�pc�k�0I�K�w5ϑF1�F���Y�8�n
@�Z�=Z� ��7	g�:qƗ-4�O%�|�<5\m�];��#�wJ���!&�W��m,��1��vr�w��#��fT��1j�>�"��Va.�ȉwɊD�陳C�_�'�>�tv�	����k|s� ���M4�{z%HL�n�<z�f�RvZC^^h�����t��h�+O/U�3���^Η��uN������AMGx���J3z�����Y�������fV�hK+�A�v���nVh� ,�%'��.�B�%qڷ����l]��]6��1�fH.���H_c�!�4-��u�2�u�u�C��{�w�rU�M0�=J��B�����v�	��&�,z��L���4���!
��yW{&���V!7�B�¿[�?[�����5-,�����(�o��\�wEu#��;�:����kzH� �ͭ�6����DA����X�6/��u�,�x$ں組�����N`\;i��3Y����Ӄ����'2��&b�Й��F5��[Ov-�k��;�U�d=t�|n�����>#�Dѡ@W�E��eb�����i%Ve���X� ���X,���"Ƞ([`�����b��UA�TD+%VJ�QH��d�QR-�X�TFET�	R�����(�d1�*��B�T�"�Uh������jU�+���)ZAkR
(,,P��Eb�dm*Ĭ(�RTZª(���V�T-*1AYmPV4��
�" ���0EUX�X̥Am�X�e���UD���E�TX�RJTmJ��(Ƶ`�b*��֩R�iEQB�%�%jA`�b�
(�b�YR�UDF1E��QB��PF
�E�$X�iDT�a��aD�m�����,X�
���`�T��Z��"��-�Q��V*µ
ʣ��d3Cv�X[��Dޞ�J�R�I�'�0��ά&�X�m�CF���f�zS���]Yu<���3�J��ޫ�D��YY�������]G�]UGk��=ƾ�s#���&i�2����v�Oe�k�9\*\3�{�ok5���fn��T|���_����ς���u�z��s2�kuaױ�f��,��yΪ<��������T�qvȉc��b���P�����X�n�k�>7���b��'~$�E���)ٟ�ff�{Up����,��U��m�qD��Aʠ�AK�"�[s��y�>畄=1��y�7xj}bG�����v���ge��!�郥}�@J�3�be��]�Ş���Uc3���;s�ƭ�(f�x�w����W�-c9��!��{�F׫�Jd�w� 6D�5�r��ቻrr<G�u��t_��Q��>B�n��G�(���7��hm��/�� ��CȬ^�wX�Ta41��O����Ml�����dc��jp[=��n����[#"&%�PomoA���S2*<t��3(8F�e:�43mW��G:|n9��=�����>�.�&�{�3ahh3�'��s��e��>�$�"�U2a��'�X�]Z'\�����v�^,h�߇��g�$۸�h�Z��J��+�������,��_�W����R�^��w6뽬�ؑ]�,XE�~|ɘ��GyK������ǭ����t��׽ 9G`54�suK�_1�ѝX
�ӻ9f<��g$Ak��A'0n��Ju,����z =䵀�M�H(S�k�!�w��5�G�S�U���B��N�w�&�;��V�Ǫ����������޶G:� _�+����:�����{/:.�yk��M߈�V��kf� g�J��F����b��@Ԯ'N}���U�uU�s;��W�v�k����p�:�~�p�:��k��\����1�Qƃ��s8h�<h�=`R�I�r�|NW��7Q�����7�����:Ęy��A~L�5qԇވ�l���@����+솽�e��:�2��}��;*���޸9�ocl��-_H�qZF�kM��A�EA��
��u���m����zh8<n�Pw�b���:��gD��=����ͮgk��C��/r�i�'�8�0�ʘ�U�}C���UKb���Щ����r����m�z�1����z���e����Ҵ�N�`p�c����5�
�~;��'�X�z�@��7� �'�����+|��Gȑne��G�vX�9�ߗ`�W�.�:���K �@�8���r�E���Ӯ"��-�_�����N+|}T��n�lК<�r+��9�9z�)٩�W�M���f�uaZ�7�}��Y�*���G.\�B�e�x�[�"��.�K�-o�&-m��Ʃ]�,�ҥe�q>R�+�R�l�B�?�U	-��Oz��j�^�9��z#�[��큷z�	��_�����Q���P}$L�\qh�bu|�?w9�"�^Kf�5~��}�m۲��|�ݨ�}h�yV�Q�fE|�J���n�DL]:�42):|zc�ޢ2.\��̇%�۝�k�4��#+5-�[%��aө��'�L���Xb��_��k������H�@�V�������N������!�U#��x����o���ީ�mK'�>#�06C�����Y=626��sR6�|��)�w_�u��'�8� 9M��� mB����x��%�qq���ۅ۸g܆*No�����ҽӊ������dܿP�I���-����m�q1&��Y6�x��{X�;��e|j8+�����Y~GK�x�j��}��=�:��'~��x�����s^�goa�R�J���Y��_����:v�����C�����*U~*sfX��< �Ο\ª/6����j���,.U�)�HͭW� )ҋ:<Nf��2�������T���z��ʃB:[U�YQN}��;�;r�i5��|�o�Q�ܨ�"O�L��1�yo	�P�afT�#���ks��;�0��Q4��!�*�Ϊ����%�>�t�(�n߅�[�)���|6��Nu�.��ӛ��90�S0LV&)j��пen�]r��;.$��ewZ�4$�ǥd5�Wr�`��m��\N�̦�J�l�q�r�@:���F�9��X\χU���E8|n�ͧ������B�E�t�ĔV���ٙ8]-�/3e�R#�EНC�o�!��i٠Ag��Hxg��?mE,���YE�~;�b��CU�N�@��x	����-/��-8�oK������ ��W���z�юy���9j%�n&�O������A�>AH��u�x���J=^�#���Ҍ�D��:���M;���;??T��U3�J. 	I7�C�#��S����4M?=���.�б�����_�7d��6z:V�:\���p�1�b$/l�̍��Xj}=�I맚k�w��}y��z����L������*��Q>�d/�{�ު���v�R�:���q;6��ɮ��>00ouzKn|�%�5�h��RA��;>����y���}���TR�������xܚ��g9�_s�2+����m��tځJ�ѧ}B���ޱ�9�C�d��e���
㮽ǆ}\��waO�n7�1�eWI�6�4}75WU'&�~63�
����")N��KV_���gb�6�w�<j����@Tr�����Ѯ1�B0Qĕ�wX��b{��7�ʹ�㊚��&k�Y��i�Ҿ�w�c�-Yb�M�G�e'C+P���ꀗ�d�b�w`݁��g���Ĵ=P1z����$�tb�H���<����z��1�oǽAN��B��W���{�8�U��lFG��Q&E�&�A��}�!|bS���>�Ů�{G�I�x�]Tz��~�l[�w����:>m_n����/�ҏ-<MT�����:�~���Nޞ��F�7�m��r*g���5�/?\����s��C�q�[5�����;�B<��K<}[}�ޏg,���+��jJ7.e#G��d48[�N��������{#%-��.'2Xs�5�ݙ���ޡ�ܖ)N���	"�MF��RQ�oZ�p���/��N	Ѕ/Zر3�w=��j6=�nwjz�F�F����� y:+�x]d�|o��aǪ�>]�7�����9m��j�{���]��m�{��:}0t� yT`O���q�-������Xm��V��p�8��\$z}�^����+~�_��t�:�� ��eߞ��8�z�x�ظ��}H�%���=v(f��{"C�����i���z�����H�"F��0���6�ʃ���(��{k����L��7D��Y� t�ڸPW�!p'r�.a������Wtk!uս������[������_fEε�l��0��UqY�a���Kt>�<�էv�A��*e��s�x�d�Je���|���ܖ�~�'?V~�
S��)��u��B�[�6_����9��yց������ݩ��7�K�f�x��7d��m;�t���_���F�[U�+ޟ"|VXW��N�a�<�^��:�uϘW�u�Lzk�2+�Y��>ȟ/�j�W�l;+Fr�9��U�y���3ה�����^�I����d�,z�D��т_�x�^���"�)W�+U{��ju�z<��?ff��r{�3��z8gП����zed{�@��čw2:4�}a���0��f�Ԝʗ��c��t49��۟܎�����u�x_ݷ���y���Y���7ɠ�s"�6Y:r�≛�����+�mj������C���q_��T���^�U^�2�1�R���o��лݘ�A��q3x��srk�t�:v�"2�=�U3f�'Y:f�8z��~��&�7p�l���8n�*�w]�z���ފ���5��Ȉ�P'=�2S�$F:s�>���xFzW��£M'��ЕFzQC�R�x�����j1�s:v��P�Ŏ���Q��t�\��}��2|�@ڊ��v\쳮�5]"N^W���w�����gwY��G�Ѽ��^q
��V��߻�WW<�2ޑ=Y��KJ�����/4 	��7�tKQ��h�6v��9z6�0��
�>6\���Ȳ�:{Ȁq[�V���s}R� .6cuf.�Q�;U^�9W����V�����$�!�Q�D�$�#�`�S��۟w���}��,SV�GE"�\?�� z\��	������y��7=熄T^Pp縓�WS��ռ�='��^�bܔ��`���s�>�s �!7�"c�]�����>�2�#)�0�SY3����Sy�{.���h�a 75���W��2�^|����~V"Zs�k�-��`7��ʢpk�:csՐ�u�Һ|Gq�3�L�ơABK�
S�ƕ�ᐎq[��[fy�t΅��ɗ�$j�]�=T�͓tK��-}�<c��J�0���"n��d]r�����^�s�7|*��9٬DU(g���_���K4�-��Bǣ�(�x��`�ܧ��7?%����.�t�]*j��5�:;�����~UR;�׉�z|{!� %��AE��!靓���?V��W�{�cB��z!�;\g���q�uƊ��3��W&���s~��p���C]̂�����u��ٷ��7)4'Ĝ�>��ه_uz�Ml�izwK�Փr$n����{�:+�x����3�K�>ڙ���[��v�BcL Df�%^�9���ܕy8Y`9�yI(mD��]�S��fCf�u�39��}�k�U/[�n�Oi�i�[���O�8]�)����4m�+�1ⲳhs�u�x�v�xU��: ]W[�1�|�@ᎳzF������}fɷ�~����z鼿��5�'�}{����u�(Ox���7�b�.�c��^W�������7���"0�DL���C���:2*U~&��,^R�.�$
�[�s
���y�=���ϫՌ�6��Ud/�ҋ3�&�~0&�þ��U�������E�o�W��vqx����~>����	�gk��}xk�j"�O���,-�<���`��`�Q������G��T��?P��P��O�d\g���G�^Y^�<}9\\�ʤ3Πϼ�'o�7!�&K�L��r90��:�����dukN�|�=ovt7��fwi��ˁ���v%�+8�炽 �9Q�	3�,	�@\F�$|25�W�'Zr���g����kK��x��˼���>�������lj<��T��L�P��]�;�!F���i��:�ٶ�*��ݹ�-�G4�4�iq�ӎ	W��D�%��8�#o{.�]={�������oZ��ӽ~�NY2 l�\�o�����;��	�J��y���g��DQ�d�|31\.C�43�e�:R��K�-���x3dL,�r�v��qϪ��%����ը=�ͱ=�^��?;,亷�Hz��3�[v�j#��Y�)���FH1v�*/c�f_G[ڶ��3���RQb�h5�-mMJCO!t*7Gt��=P�>{�F^�0���D�#�t2o� ��lǼ�F��z���/�LR�O����`����~���������fa=�I�n������C�s���~69\����[���9�}R��3)�c"2���'gY�5}�Fs���I����v�4����d�&�Y��d���z���4�h_�7�w�����-���!SĻ����xIٽ�$��F��:��p�͞�dY�Z�����{@V�ٮШ�T�4Ө�on��ng��=�d�~��y]�����j|vE����TI�g�w&����ui����k��Т���Y��S��w>�[ TF��c�S���Y�zhf�ã��R)N`�^�"���F3雽�g��܃�ia�����5�b��Hȧ/ޓ>�z|�pj�о���潗��;o�M���IQ���%	����wtn+g�1z�@�L�Ѽn�!�sV�{�V]r��D�߫��:���u~D�iA��?����2;*��^�>��^g�2�'�^)�f�m��Us��[g7r�~^������%�f�� �ɑg~��a�#��0]��N�#����4��%���f����:u�
��8�Q�b�RP<��]�z�z�,����&VwJ�Ê�[n���J��}mMz��u<ˏ
o�
��(��eһ*5-S����ޟx��;�,�9�
���e� �.+�~�F�a��)��z�� G��߼�e�ϰW�+��C���d�������a���|�@� %鑔;/z�C���*}�[~ǳ�}��#��^�����+|��W�\���rx� y!���E	��W�l��k7����|���g��3L�=�?8{;�5����	l�U��*�gF�������mA�=7�@�jI�\.#�Z>�s���Tm�߯��.3͚)?�c:�S��щ��ww����p��g�?��D��w�y
��9���5pڿI�5�&��V�������ǃ�'��3ß� �4�d �N�fc���ʝ��m��Ϲ��S���)�s�}w��.&���0D��&�pǱ��^��ɂV�'�@��u�zz�&*�l	�;o4���=��7;ʫ�'븸���Y�U��+}����U�T�K=eh[���}O��G1	�Y�1�ܯ�%��r���z!�߯�~����rc�5ҏU��m&����ϞmH��]��-��>7D�zG�r����1�~MtY��H�#31齨�YˬN�YԏoY�[a�wꛩ��Kb��D;������S	��N^!-��lҋjA�fN{L5OJ��Det��]�i|���(jW�@��;�բ��:��Ǫ�ǽk��hw�fsR�˲k1�(����sE�r�:,�{��p�	N�[�(�O,K<Y{@��]z��Z���v��QW�Ս��3e�=*�&��s�#o>���f�v�q�e�f�ӎ�������h�iV��-k�s0q7*��ڍf�9���pg�Ky�A��m;�'-P�;�U��W�q�?q�A"�=����M���`X����Br�� <K:`W�Օw�ˏ��flȺ��o�DJyL��:Ţ��'��`{�X2[�o�+>��Yw���Z�U�Y��C�Jr"����lg6ǅW^��Ƶ�Lb�_K���V�/�U�����D2q� A�8�����"� D����(������}a�K�ܱ��G3T���=��v�3b��\۬@��i�T��ǃHݹ���F_4��1�>{�,x�li�X1'[X8=ک��X�N,�j
ڝ]�e',�Gպ)�0S5t��C��RT	ǋIU�8Y��N�yF��9�wS�q4N���j���z�F�{��8	���e
z�wX�{]W�k�jU�H�j�� 3w9�8kI�qVCt�^��6���m�\�ϯ2���U�vlUk;�D����M:��wd6���G�vN�ۈS��`9[8�d��1|mh�;�y�=vf1YW�jn�����j>�ѧ]x�S0e�_z�ǽ�s��9O�N�d},\tT�s
1gَeop�8L���{�W����|7H~k^��^�ۊw��o�v�K��|JS��k���
֗��K�Cc$,XEc"둼�e�Pb;�$�.�K!f�:��];�0ݸ4ՙ���Z4�_^�˫R	t�-���P��6��qw�)i���qI�,�������o�h�����v�Me�Ǘ����Z����V�H.W [E,��`պ����`�O4�,{��#g�����2c�u�G1����c:���Ҳ�$��Vi�g2�{*JXM�]1o�����5�o���
E}6�1�MK0Vk-k&��ҤZ����+%Lr��� {�՗���v�`�+dB����+�fXZ.ƽ%��5��@�a�;QZ�{���s-I�Lb�r�5�΢K�f�F����$���Xe*�N�kܒ��.$��	
Хkέ�Eުux��A)������5s)oRiU�FN�SM��[�YN��.�7owq�Z=>�V��0᣻r���1�v���U98���,޼z�?�k �Z��>�-�������Ql�,'��X���S.�[���`�:���zl*�|w���;.�J�c��%L����V)XVB�(�2�`� +U`*�J�dX#"���
��AJ�� �1ADJ�Z���`����5�*��A��QH��&%�iek�H,T`�",�QPX�QVH����b���T
ѕ��`���c"�Y�Ī�*��V�V*(�)���R"���"�+
 ,��+QB�)U1L����0(��e���\IE��*�YQX�U��DdTDX�*�Q�l�b*��pPAƠ� �����F
���"1D�S̨*���e(.2�F"����"*��PmTb���[h�TQQQ�qU�X�D�!F��h� ����X�mADD��"�E�ňԭ�E���b)����D�PQV(*��(�� fU�UE���m kg�OpD:�}�~��س�}���r��Y�1/i���ao৻��3"��:����$���Ȧ�i��͹��o�4����꼯�ά'����Zㆥ�:u2���e���B���׳i�PA�`�;ŋME�y��A�=�F���rL�u������*c�����/u%q��4cސ1\m�f_mo�Y��c���Xr��^_c����<��^�·��Ϩ������E;U�J���^@���?2+��x��b�>�2��ڰ|2��������1U�"���>�Ɇ���RJn���J�8����5޺���� �$��.�a���O?���V��!nz�~L>���ٞV!ߘ)bqB] {�J����@[ٺ��n{�� �1<|�� �}sWD���zϤ�>��z �(g�r�^�@��&�DO�;�٧���<GݦC�>���2+;;=���_9�p�@6L��I�~u?��v@�;|�DKNwM��w�s��AA���r��Vbb��_��DmD9�f��(���(*R�����݈u�|�5M��Z�P�����a/���nw���L��C�xǴ��,�{�9����P]�w�{�3O����Ei��R�א.`��5�&%rm��o;���P#�=���fxR,�|�Ky� ���������xz���W�PG����k����/�p>�F�75{�=ہ\�]� W_�!9�*�p��r�(눥�J(��5@E��oQ]FI��1�2)-�X�1����?+~��,�i��б���(��O��D���1����or�y��GY �
��gO�V�i��R���x[�~n�M�{��;ά��u �)d��S�(M��u�����.PA���6G3�C2E���1П���?Pn=����/׿%�V�f��ˍu+�K���\F�].�
W-"����{qiz��5�����X���^�,uX���	l����Я�l���� �o��~�J��~���<���q�����*.ڵ�g\Y��ǣ�W���]���Y���38nr�e��?N�fr��*�t��;�|&;�k���˙�X��< ϧ���r+Ռ��1��uf���T����*��P�`��%*1�����!B�+>���#Mx-�����~�k����U���ڈ�Rx���鹙�@�'�#N�����:1�!��FV4�}��bF�z��3��z�<�+և�����UdIT�T̸����q�d�*b#&EНC�P�����f�y��y!�5���>�D#ܻ���d�^}V���+tbv{�=~�N��n3լ���R�繘]Թx���\"���}��z��m}��N,ᇣQ���(�$ �C������_T���e�p�����Ħ�:+���Ih�/�ON�"w��MNJ�xoꜮ�'��@`l@�R�n�>�O����W;����Ve��vE��;���3F�Փ���Ge|bx��ώ� -2��R�f�8�e���]���q4+cʵ�Zf�}b�U1��{��h�:�6��4"t�����-wdK�5~����Nb��z��T[��kƷ������f�?^���&[@�M4!}�J.�����O�e�c���r�W�_�1��[F����hu��|��������"}��:7s�W���o���i��sS�ly�)��q�p}JܞF���_v��g2w�\m��t�~���e�}C�x=1R����sq�J6'J ��82_W
���_9|y�j<�����+��F�9��ZZ=4L�� j�{n�GdɨS����_�=8��K��j�/>�q�7.����U�^
�Lc�B����ix㉃Vz�Q���}C&�����tg���;5u4S�~#}]5�K�U����ᐝyg�zg�V�^8Ū���J(ȳ���05�i�/��?�
0ھ��:�����̭};í7+=�_�W���k(�t�t����ǉhRӸA��gږ tΙ.͖vq���e0g^���F����W���n;Ÿ�����
��q+r�8r�J��Q���l��57�`��C�x��`��xˮGƕp;���+s��2!׫�����g��3��Ƕ�o>1~tQ+{T+�v������4�K(����?{݋��#"��zNW�1�目�#:l��ݾ���y͚�H�)�>����L��6r\�3����Ʋ��G��L�e��b ����q���b�}[��GY������ѷ�y����.��o�^S*�����o�ߢ��l݊�����gA{�U�Q�;�#��b��9F4���,	ȱuʏ�τ�@S��ձ{������%��S�!���=�]��r@o�<�GN�Y'P1���ñ�v�MyF�C�2,��8�`�W��$\K~���V�Qүҁ�P��+�rQ�I���=�}�x@��=��M���z�Ƣ����_��g'���ޤ8��>��tp�=n4r�(�Վ�LAS�@L�I-�qe��1���Tk~�ˈ>�����P�R�}�FUZ�&���yV�^�fiHƾ5-���DͿZ�+���_��|�F�ҧ(	��)����ӌlOu�:i��m������19�/lKdTJ����F*�gp]��n��L��3I�!F�L�FS}w�<yϗuhv�i��T��r]Jm�V��Y+)j�����X����
޼R'�=3�f�m1�������������ʹ>r|�S%��L��Gδ	sNfB�际�Sc#)�~,eVߟ��^_G�y)��!?���ݺ5\�;����o=J����-�=oC����7�z�L>��0��>+�M������A4FҞ�������놮�1���E�?P����A�U��}�*A���f}�4-8�v���qW>�^�/�=sJ�ND+�#�xhq�{~�W�����U����	Uܺڼ�yQ;��[ �B�g'�<M1�^�2n��R��Q�M���7���!�W����B�jB�<���\j4���9�`��Xz� \_�aT�
#Y:l������2䛁�:��F��*�{8�}�9�{#��r�U�pz�t/���Y�^��>�t<秫��/�^���o����77^Fl�S��ɮg(.����Ɉ��ļ�w�x��_��t��Gx��>T}�gSϸ��8�O�
=����{��T�P�za|�i�<I�v��je^F<	���u�,lZ�r�i�N��=S�����ё�x�G���_����&�������8��A�	�o��@�<���8Tz��e�̓��/�4|�ݸ��8�AɸOƽh�x���=���o������S~H�����ҹsrծ�"<��(Bz������-wD"7�De(�S�vY��w����{F(��M����"o/8����rypT�t�K$���(|��uKe�wp|n+�뉹n���y�5_�e��~���s�`8s�觎�x����;��C���@��x���e����S��z�.^���_�p�օ�i���i�>���^��{�fiL��8(#�"��c��c�Σ���Meb#=�2�4�I�K����/%��M���T̊S%zn ��v:�����������G�̫�3{�V{�(;�r�6��_���㞙��=Q�'�N�
�,��a{�(/��3z����-�c�Վ��El�t�G:c��w#���]ȿ7^'���;ά��R��N�TZ�1��^Wh.ɡ�����ARܜ�,��ם��?mx(~uro�>�xh�^�=��s&�ߵ�ם�=������]@8����k,�1�^���Ȭ���߻�mhA���z�IG���[��*n}������l�|k�:EV_��+��G;��� n&��
�3�d]�����gX��Oz�m-g��q��M3���Nlχ�:�5Yg@�%�-���C<t9b~̱)���S�j����em�c��ײ�����~u��m+�+V����?d�f�t���ϱֽY��z�*���NOx���޻�]�냥�c{�ԑ�s7\���qX�.U@��U�C��Es�����dV336nJ�eWT����%�#�0+��<� ���3�w�{�c{+�:Qf~����S����#W�sN_��w;Ӿ<t{-U�'�kMxR�S�M��}^�ⲝ!�s��:�t�p닑�:�~}q]�xnC�U0`]a����7\��z�C_i����K���/���>�<9r�G!Q��-�����ћ��ޥr&8��Al��C�&G��x�ϣ[����{N{����nF��7~ճ�܍�B˟}]��'+���U
|	=_L�#�Xt����t|n=~��G7�������;<j�{���,� ���p�"�.��Q��<�b�^3|e��!:g�yޅހ�Mz��6��Rӝ���v9�7��6v~mH|��6}0t���ۨ��Ӄ�7�xUQYW��!��RG�2es����z����2^K�7d�me4Є4�����D+`��j�U03<'���U�7�\�_o��s��,#E��lx�Q>~3��q�:�ɯr9w��w�{��Y>�G3 ���%�{��b��2F�˓q���cg}�~����3�wZҘ��Eճ����h������J���AS�²-67����3�X��V�wX�<j�O���2T�U���PWy[.���9��ђ-v�.�R�*���{��s�n���b���v[x�mѬ�<�E���h�}�
����:�+��
��G��L��Y<+�3/��*pVS��Y�m/���_���s��L�Zs3���8��/n1�[k��C�g�auP�v5��{t��Ȯj�.a��Kꍵ����k{[�Vj1�3&�e�3�_1���r~j�Vz�Q�<K^���W���!��F�3G�'�n���R'���=q�w��!:����x�ޫlؑ��S���wQ������Ƃu�=0R0�Y~�u��}���<��ϧY��]◧�,mk�,t���ｿ�Y�����b&��Eڃ�����'�)��@V��$dS��Iϫ��B��'k��Wos�sWj�w}�������;\�|6�e��}����t�g>�� �}>$CT9�9��{���v'�q�q�����E�{m
���:."ܒz�P���u�z��s2ʸ~�=ue_��S�8��O�(ޖT;E���O�=�b��9F4Ȟ���e�0�c���$��>��j>��f˫�x˖��{\�g�=�]��q�Aޘ�GN�Y'k�#%xv�����91�:�B�12���������Y^���Zo��<���y�}��B�t٫��S{�ʋ�X��F$����]�+;ܕ�O��r�Guӫ�bˢp��L���:�j���O�2��>;ef9�d�gvBx-���ε��IFuRY��kfE��{ޝu0|���.%�^����+~�*:U��@ᨇN�G&���F�վ�B����Q=��D�����o�^/v��ny\U������:��C���W��0f�۽���=+��/uV	��2zU����"~�끿�KG�c{�c�$G���vTY3v��u����z}ӵ��{ՠS�fQx�-�zH6�H^����_�8p�����=�Ӿ��Q�,K�/����=%��[%�Õ��:DG��O���{UyR匯v0�ag9���p����Vᑍ������0w��c��W�L�������g�^k�(}D-Ǒ�i�f<��ʽ�����놮�1�'��?P���z���`�Z�#c���efW�	d��c��w5��*�G�ҿ����y~�	羼��h���&N)�������z3r�e�Y6=^�}U�Jxt�ٯ�c��2�e�3>�3W��b��)B�k�t�崲;��o�V �V��i�!Y㛟�_��]�Ϫex�r6e������42+���P��Ӗ%��-���
|8?��]n��gб��������u�`���ޔ��Uc��2�cLE���Y{��t��G5J.�e��M=�n-�N|j���o	�1'�;���"�l��&����[��=m�������b������;�W�k�DN��"�8�d{��B���3�~^��ne��3�_]z����k�`(SR��/���Ҩ��=�O���z��ϩ���Z�U��̉<K�1ީ��G���;��<=�]R�t�L<�>� o���h���=�~+"�Hya���e�و�EL��D���^��}>�M��1�5�H_]S�'iһ�|:�����/�p��n{����WKg/c:�ب��:�L5�*�3�*`\u��>*��{B�9�!����"��+��C�eC�#ς����� � ���q��}45O��Msl�=���ς��͌�S^|�<r�n���>��q��AE�AlD����[��K�cq�����;�u`�z���6}�f�!���نk��#,����%�<��q�#�d���R}W��~ک��	��ʚ{;�_�p������϶_����hl�����t�@����m��Ddx�L7͋��3	V`�K�6Rٵʡֵr�ꈣ�}�[�����ҿĄ$���@!!�	'�H�	'��$I,@����$I?�@���`$�� BI��	O��H��@���$I7��	&@$I,�H�2�	'� H�2�	'� H�R�	'�H�~ H���
�2����XW��������>�������|y(�
P� QI� �   ����	(@����U
H�>�p���I �
�BU
��J�AEx�H0|�V�U[A�l�4l6�b���hw$E(0	�N��06e\  u�  .Y�֭a�mERB��*�ua��im�&���eU6-��U

 M�[dئ���Š�&��T��Tf��j�R P�d�ʍ�Z���B�0��2�fRW;���%'`h� �U,�؁�R*�5R���e�����@F�LfI�"�,(��b�vs��3-Ъ-��*A�"��EQ@�����f�cm��fiT�6a����ȑ*Pp m�5F��ͫ1�i�Q6m���5�%T�1t��)�3h�P�U�2���*׽@�IP � �=�
�)SM4	���a�h1S�)*�h �   Ls���Jh��@��  E?�)R�`4`  �`$@�4	�)��y2OSh�7����S�@%$�4�4&��  ޮ]]�ye�=��٥c�il��H�ل�+�ǌ�"$s?5�#:�I.F:�Z�o�"Gw~�%�V�������_��i����r?j�I�*�	��"E%�6󵄐H��I¤2J�
E�*BHHΤr���N���͟�&EO���ν��=z���[V�Z�j�F�@�"$�A$��I&��$*��E����%UQTy
��_��wd��6�oͶ�i�6�m��㖝�/��+z��0�']�*Xť�d��f�>����W:N9�K�Y)*���m�a˕��T��~>���g�F�J����%��s �Y)��(�^�+*�Ӗ�63P�J�k�(�T�ڕ��/B���ڭ
���!�N�pˬ!�+;�<�Ч�_|�[YǱ�N�o�9�5FR�c5઎�j�K29l?�k%j�.�G(�:��heೂnkR�%1��Hi积^���%��=ϑ.�&� t�Tt�Ķd�L4誄|fe�u4	�Rmc׃si奻L��w�k���Ժ�����p:��f�o6Y�F=5�y��d�rO����{8  |j�����Y5�ɋte
un�������(R0hc��4���f�e͒�Hsn��%�&������nWg_���H5v�ͳ1�$S���/^8�Ь�--A�iH.�����s*}�,��`D#5�lc�m#2���a�0]�˨�d��AMM��Vc��#,ц����4�I�Gv� U3t+x.ͽ`���{�RQ��o�=�E��eͨaB��Ե�G���K�g/%��a��{-���a,cK5v�ؾE`V�V���60�s2��c,� vt^���c�v�P``�El��S䆨1���ˡ��`"�@l�{/W�����-H3(46�M�{�Cj�`���%��J��Yu���I�֜����O74���"����L`Wn�6lc����-+��֯΋��3R����a�y�ޅ��aN*�g�sǻ���6T9���D��R�v�	�q�m�W���^�4��y��72M��b��·.������Y����ZS2P�tnA���mbcq����)��F��$�N��4���dYL㫻3&-[%��/%��8��J���MlB,;{)Z.��
gF��e��.Q�kH��6&7�eӬp14n�ʁ���o �҂p�7z�^+�GEf�f��T�flQ��A���F��G�h���չ�֗�EU�DY�Wn�!KI�x9mdx��9(�\Ax�v,(�7{d�9y�b�5/�D�o(J�p�aE`[j��������+�� �fB!y�{�+Q3/Kd�(ȵ��,���V
O��JVO/��ab�b��V*�fX�G�������p+�n �2R:���ۍ��t����PA�1���K6��+�Ѧ�9� V��h����l��h�U�#��]lu�݊��pL!S��ckAb���NV
wYIѺ�Ų� �V֔��Z�k�J�#6�+*9�
�H�H]����	�L[�̅Ɍ����L.�^5�k�y5��IX��1X���\G���1L���SPD]a'r�h�o�i}��I�hfp
���U��5�nƥ�M`
n�F�ǀV\�A��ȌiO&�(���KwQO�v6�f�|(����@XYB����ac����tj��A�A�X*�+��,��/�����4v��r�[�lL�w'���R�ZՈ@��]�{�s2��l�N�j�Y�Ḧ́.�v��b�U����,È��̽�Y��NS��t#�]n)&	��C1f�k-�~��L��M�U�؈ռ4d�5XDb���Ժ1�Zw�i�d%h��)F`�0^�'����x�E
Ϟ�EԠ�u�N�"�V�*
n�H�GY�)ᙷ��؀o���w~dٶ��WY��=a��#k�>�6Fn#u{P�N����Q9�,�*��*�!l���Z/�ܭǺ�����Hަ>�MN�8AHW��Y�N��N�rb�R�9�/(I���P2�)GW�pYܚ��X
�Ҁ.��UsA�n v�c���+W��%�'�Jw8[2���B4�4d�4;n]m��;�.��Z8Sv���S��ؚx��h<.��H4�bl
�Y�jf9%��mX0�y����YRحY�(�U���.�X��ր�/u��+"�h���Y����	j3*L�i�N�6���1Ք�Oi�以�I�ue��Ks,�-2IHYBa�7#T� �'x{n���eec�dʖ^黶�EXզ�82^�_ ��c�.�:��:v�RӪ������iY���dl-Z��S�Gq|I(��@��/!����7�r��!�B��F��?[�D����it0!���R�[FӬ�Zw�&[��X�$����b���ؓ:�!��)YdYkMm=��`v��p��P�f^�0m͒RA�4��v��1�H� �T�4/w�RZ"�P�B��װU=�6���M݀!8E��Ǻ��H����e�DV�X�h�R�(����{� c3f�,��֭J�Ơ�۱z-�`�ؙ�Y��x�c��Pz�3�Qe$�2��=OHU��&�3[�^
�Uy�5t*�o�xu������ٍ��RVV^auu��"�&��՛VjU��֪d�e �5;��ϕ2��5��\rn����Y4�4��XN[xЛ-�4^�;I3�Z�ͽ& 2��߯p�:N�Ʈw�r���ȭ��Т��&eIqZ����&.�����MM]�,A �N[����nV�X�eZ ��F�����d���n�����xB��ؘ��7J����Bx^�ͅ�"\t���c�����a�q�����ۤu>J?��m~�5�����������بv��yҌ�7r�}�֫U-%��yh�3���&���
��8�4���"ڹ&l��s/�<��P;���fm�)��ɔ8�H�u�"�ݸ��]��a�&;��y�p�5�Y6��U�e�AE0m�k.\�]dO�`�W|�9�|9f�Z��JSTDwM�Uh2��sq�>�t��h&��3��XZF�h�W���q�ț����fՐ�<:j=u��Mr��t��ˢ�������z��(b��S�D�7���Ge� �q콮���e������/�W�����PIo��&�5�3|յ9Y�Z�<5���|A�R�_Qz�k�)�y���vcWH�3u�bؙ��R�T�V�F�k2:��0��w](m"�ٌ�B�b�{3B2�.��Q�:��L^�����tN�8�X%H�b��y�X���kk%��5X��;��� �\�x����Q�"F��ʎ�r��a��|����%�*�/d��ȴֶk+�;���u���T6� 阔�%S����-iO'QT����LF8u>|b*gv�%8��UۥH� �-	^Y�Q�2�]� U��&�F�]��oq���l(详8�o.^1�'�]8�&���i+��⽶{��˜t.S�s�a��K��$t}�Q��pU�+�;!U�����l��+�p�u�3��%	O60��s���0�J-jw�m"{,	��*��9�@�V]�F�6E�}��2�ٰ��.�ݨ��S�ʇF��;15���ɸ�S�B�.�K�.�<�Zz ��4M�o��i��wK7T=��p�'v�ԋ��Nf�`(mR�	���� +���)���\��%��� Lr�]�ټ0� �,�/���Ϋn%��r������ʹ�����;��r���*X�v5��S�y��]X�V���Vx�ِ[ӻ��f��?�̣W;6���n[�I�Q��wD+d���-�}φ,+3�����P�I	�������M[�۷�����]*WC����1N�����cۨ�tk�k�Q%�9��}|�8�A%��C[;��6s
������K������"8�3y��ˣJd����sw��p��G�g39V���q�[*U��9�0mV+������^u�Q�Zetn�U�ò�L�5�����+n���LMb��ҵے�+t�ˤ9�P��aX����Tjݴ�!�1�c����D(�jKefqJ�JSz��ٍ�غ*sy8#�
\\�Z�p�S��c�f�>���P�^n�BZm���Ow����CTB���ć�e\l�?=fK�ыgf�s��(U�N8joA�([�am���L���oݪS��P�m`f=��G']�{K�k�B^aNua��%%�aL1�dD�$�K���zseJ}Lw�Dt�*{4n��.h�����u�T�mP�������[�(��7��Ȗ�vC(Yux/}�3�.�{<^�YB�3���gB���k�%�5Rt��W�H
5�mc�GEj��kv�em�O���<[�;��"����Q���E^�7K��c�Q�yy�:LQ�h�(��0i`Y���rS��#q� k6������hTtCX�:]wV��8�1YH�ho&oD�����zڻ�u!&�c���۠Y���juq!��/bY!��V���Ƣ9��s�R4r�:N�e�ꄸr�^�ʹM1E���EP[.V�r��6奜�Gd��������:$�)9���!2��H��6o^E����r8�l�=�,���j����Kz����aV����Ʋ��)�R��M��3��gA۸�uu@��F�!K���r��{m�E������|
��6�|�.4kf%�ڮTٹ���;v�S�5K.�W#�sy��-32ѩ�̝�9&�wu�Wgn5�.��K!|ڢ7�`m�ZUm۽��'����]l�\�c5H��{y�E���C�'�b��rr��ĠÆ��2��(6�r|i���j�B�g�f巭К��c�DrՎq՚���3<=�q�?G>�FA��٦�y�v���fn�S��P�Q�/�>�+A��S��$J��X4�4��]�`�'M��ܨ�*Y����"p�)��:8��n95�p�ts 3�%-p���������w!%G+,.Qΐw@p�Ih{2e�G4k��F����@I%6�q�;$��{�������r����U�sq�x�:��p�T��hH�#�58��EF���XQ�ѽ\�椒H��rԕ.)PM�˝&f�T�:'$��>�2<�}��$ހ�����{��5��tj�p�.��rrh �$��\�rmegQI�r�[�XAp�R�p5'n�fZ�H"r!�K*J=��Ss�#��ǲU��AaK��`�#�|,����gt�W��u�IG4�$�sq��j^�Fۖ��!Е[a��R���]��S���2gs��t������Yͦ�_1
ޫim8��=ͥi�l�޽6m��f�u���Ŋ,�I���̬�PҁZ��K]Z��*�l�( �F# -&�M��.�X��P �H�2?w�l�W߻s-�L8}�!!#�5��}�kשHٗ.�l�$荜7Z��=������UOL��k��%_�_o{�X�vXՑ�,㻡�4��t�4J�)#�7�m��i��5���U���F��9&Ώ��b;PBh���)����R����h�����냳{]f�X���|��R�څ��݌t�W�h��5�Q�����*4�euY���sl�h��2x�n�\���;ҡ�n�j�&р;�u��U��=`��%6��7�&+l�o��}�c�1-�h�������ua��Y�PT �b����V`���Ek��y`��o+�<�	Z�ʵ��E;�3Gz���U�ϫ���Kʄ�{�-��n�"K�����+�\ι��ppr���]H\k{s�r�#����Nogk;�m
�V�j�I6�j��Fe�H���"Jų������J�m8@���T�`��O�J��/	��aoQٛ1�X�&T˒��mv�L��}wi�h�ŋ�kv$Ă@��k�M�YfY��y�QLe������Ŧ��@7oO«%oMi��U��h�B���m�|j,��{�hh�ٺqWM�y@R�D����	w�n�`�ju��qU�t�dglFh���V���\�צ��<6�F6m�)1�������!JQ٭�W"��9FF<�R&��HGY=���hT����fK5e��e�(�n�+��2!+O�em�sha�Qk�D\�r��t���1T���@��70-�r[��)�Ӌ���B9cg�[�Y�m����O��c��1�R���|
��YKn*�(v �ְZ�g.��iPr�jp�<�i;7�]��'	�!��@v�[Yoj.������ϴw���&.̑��j��ޖo(qz�a+s��՟�N��/Y4X���:^a'vT�I�ڳ�u����M���!ݐӊq5fX�s�p���:�$q��x)3�C����t��c�t]f.�$Ӊرn�^����aU��k��5��ެ�t�J�����j�C�g2�9[�B����(�)��0���^c?`zFP8E��8�hٴp����	��'�;��w���zgXب��+Bڦ��¼QY۰�;hY��f���K&���Th�e�k$�U������mI7�]$�*/�Xˏ�� �m�nPs<���qj�Yh���=��qo��=�N�T�Vd%`�
��������)�7L5�=l�:��;p�6�}�w�QL�ɔV���p],D2��}�Y��w{�V�BԀ&�
�H��D���@���@���&�c�z����=&�q#�h�����rs���,4�!T۵��;� 9ʔ�\.�����S�X�V�J&�X��-��"dXؚ�Eŋ,��;(16��	�󍘺�zr�[����["ۮm���o_V� �O5���[�m��	{���B{7Q�L��{��m2�{m���MI��5f��Rn#Y�
����Zp������Ndf��Z73���lV'�*T{aQ�KT�GY}�z(�s�f�̡$<�lBu��)��4���ݱ��U��zhM;{���s2�T�&���ˉM�x�U����W��H�����yD���Y�Ĩ��4�/�ڣ+@ám�go4�Y�
t>	�Y��6Ay��n��w	G`����[8�ڛD����n�� �b��}�� gg���&��Q��eӰ�e.�5m�>�\;�Y튧w��5,��h�7yr�YRm
5����2�u*TxإȪ��ҫ�A�gzZ� ��[7��e��_,�)�t�v��;e��3��y���H��'�d�9FҘ��=��$H��dm��"�
.�Z���t2+�[���6Ո��H�I���]٬�C��q�s�:J@G}��.��9�m	�3iP?	�_Jͤ��0YH�B�؉��.�y���a��#Vv�sm�qҺ��v{p���J�k�|����ɡ�q4Rx�!ڳpu����[3��U-�D�ʺ;*q�,(j�k��隲��lgL/C+y���óLn�)�kF%u���]e����3!����l�n��%V�[���ٖޢ@srѹݓ4*G;:��M��0���M����A�WIRid�Y�r�d�i�v�-_a&CD1�.�<��V��=@�xu4cW)&w/���Xx$�Sv��%-Aou-�)}���GB�R�gc,��Xb�T7W˒�V����Fm�vg|'^�����7���6'��kNv;&`��[��:�,�Pܽ�e��)++��!7S�m��x>�]�Z��a���LC�1Br�Y��e�cC��}&�:�n�0]��di9�t�,t,�%gi;uv�$K����%�L��Z�*CW[�jCps� ��s5ŧ�N��Cw��`pv�p�{gR��y�8���-��VU�Pc.�Y�|i��ƅ�]���u4�%�o-n�iS�5���έ:&��z��8�O�u_u��HWOF�Y�0f���ٚ�Y�*	\���J�I�����s��,��p��Qh=�j3���D3�1lL���ڇx��5�F���CU��O�U�9ӗ��k]��5�����~�_�PQT5M"U+��W�D��~��eW@����j~������$#�;U��d�����{�ݽ���S�6�|��4Y�լ��;Z	E���Z�ӌ7�Gh�����:�w.��o��%<�Ϡ���K�pε���]4��ኮ�
ȝ��'�-u�gY�V��#�(e3d,@��Ś�Y�f�;�}����4��I�X���=x��t�C|Iv�~�a���)Z�x����]����_Y��7&��=XóJ�)�Ԍ$δ�JNl��G�FI"�I��$�4�S-�.>{
�%/��>/�%z�4((���^�H�Z�;"\�-4���L^dT�fTr��][3-�Z̊`��*�4�PQKH[�Վqd�DiW)�!$� ��!��kp�Sr[%�#�.Ԕ�� ���`Ŗ�^.�EQl�pUO�kkꈟ����s��}o3m9�ĩ���^�c��mF௫�O��ߪ�w����ϕq���ߧc�Bg�-Y6�^cK'l��t��jeF�멭=�����Gۓe{����^��ɖ�q�OĸuV*�ױ�]��o��r-�gq�7��mLt�z�հ���4�рn���-vW�`�����i/7��B���M�*�;p�9���dﮡ��,iW,1�b��x֮�:u�H��Ft��4�g��<_=N���:���2A+�.׈ù´����\����@W�[�!����uF����]������M����we�u�x�0���Z#�e���z�x��䙱L��=�Xg4�oi��"�:�p�{� ����)��u�Ա����c1"�b���+��,�ͧ��6��c�Ƿ �e'�A��dt$���Q;�Vɠ�;s/B�)?Ƌh�����P�Q�b�.��d�����{�L뛛~U6�/+�f9d�\v���99�;��?l�߻z��,3E���=6!*.��{�����ǋ���S{8F^�WV�B�!����jq9��~�/f��s�ÏD�b1㚸�?H�gj�>o�m�����=������Wv D<VE��s�*p`�l�3��T+FD;5�-5��a!U�B�u��/�@�xy��������:���|i����6�4�`0�k+��&�,T�)^�����uʓ{�hV��k��ȋ�zl��C�J��~��K�Rs�R��,��wnE/8�ң���훹��s����#�s�ώ~�e8�z��eg������ë��ϗ������t���^b��i�]�*ib��$��:�`����:�$�$�-�GTdY,A��^x�����p\ق�(� ��>���e�^��x&�+����ݼl:�0ª��mٲ&��	�hK��i�CX�ȳ��rx,N�YM�SiD��`�k��$tH����{}�J�Sg{5�.�g>ÁP�3<�H[�z�嗙Di�W-��\!�L2�*��\m����28S��=0�,e�KaOJ�[j8�29�G�Ưǖ���Ղ:!���a�#ݓA�+�6�jXѢ���+D���rH,#g��mw�3�:��CV$�3�}d�ԙ�s�� gw5tL�
�[ѐ�{����H��th?9@�X'G� ��������_CD#%e�I�Rw�\�M���:�u|�D��YZ�/X3�)�m.�5�a�	m��x�\����{�e���)�I$=&+���
���27xȹ��PJ۔k�BS9��{R�R�Q�D���-�� z��{���u���cEn��갽}2*F�ƺ��nV�70�����~븅!w��������W���m�R�j���]�R-׺<��
}��ֺ�AĿ��"RU����mh��I)N��`pL�-"j�a����ɽ|�l�&�^<\��4��ʺuz�)�A%X�f�I����C���:R��}�3Nf�uf��c;�n�Y��w��yM8��lV}=���y2V,��v�;�NCt����{ -�?_Rx�XmS�S m��<h��\I�Yۢ^�=/��)\�lX��|�҈6��[�DV�z�1���:�Oj��w��d���Y ���a����g0�ZoOm�ζZ�2M�&2���Ĩ��Z�ZH�4l������Xp�<�7��-��l�ٗ�ɢ���,�t.�U�#!3&�.Uz�*�M{jW�z@j�r�����8:7�.^�?v�W�Ԉ����*,r�{�?Q�q��-�)��g�\j��|TW[3A���F������#:u7T(�"�yy�#���[~�1*��8�Q�(e�Y��4p�s��)5�e���\4���C�,�Ο�_L��m�}��$5#x��#�����	�q��K�4xT��XNsp��E�IC=�ޚ�l������gs6[�%���`"��!���f5=��+����R�X|�k��:�WK�L�}��A�
��"M�`�Y(�"]u=��Z��M:����ve����y�kӜ��Pw8���}�ҿ�4��K����to{w����B6��4����1n�9����͡ه�R��n;uק��a+��'�`��f�+[�S�S��\��͊\;�����m�Y�E�;
 �/�@�a���jq�������GL��b��Xl�n6h-n�{I�mg5}�Ӷ�ECp1@p���]K��h� ,�v�81io2�#���܂b'*����"��dV�;:���8J���"yD����v�p-��0B��w�ڌ�b77]`���nMcf����Z8�B���')v������U��S�#��_a5�~�`�mj����3})_C���$�-��Ue���9�+I���	���<�wL]	�T�=��a"��뽨���<m%�b$�����!�ף�4e�"����e_Gѱ�_s���YA%e�����\�XG2���e��q��Us��j�Ǘ��(�{|����Cvq)�j��X�a'��.=P�:�9�\.#�'�F��z����J#ҥG6G�f9"jI��$��#�W����j�r�]c8��������i�`�K)cS		�j-$b��!$F����R�4� ��QTZ,�e��@A1D��J��U�[�E��Z �bDK$�5lK�Ihܲ-*ȑZiS��SpDQ��)cIl0�C*�
$����}���9�oR�|j�]qP�Id�
��=YA6��h�����v�'���v��o�z����1}$��7�n��o��J�K�-�>�~�b��E�.�$��ԯr}�n����~�ua���3 �9�(�j�vMЭy�>�$�_>�Q���зM�៑�f ��߼�U�@f�y�.���/�s>��}�|�;���/-�{�꿻�}�O��~׵�u���"Z�Þ�c�����ӨY$����ގ麲��D�B�����/;�}������`�����xw�w@�a&�i��|���w��[��,=�E<������og�������b�y���]�#͵��oM��\��X
3�������ƽ�%�y���Ӻ�Q�cm�aqG[�g�^�~��ǯĳ�}H�����@�^��R�o~�}�}�����q߻b�;�̮����?y������+OV���n�`���I%}?c�RFjߛbg���!���/�b�}���O_��7W�y�����W�~�\h���ԉ�����#���#��?{}��?j=a�o���ˣ1�n�$�8�[}����@we��`�O{'�q��3m���)��*���c���L�i�5�����M�7�FR�oq��+�����W���;���z4����0���v&Q#][��ϊ^Mw��`#3G(ij��eF�I6��).�����o�M���c��}��ܫ����t��+-|�=|��^|���lU��?�����"K��lU�"�ޡ;���g����&|[��}�`�P�2*�h��:��1��21X��:�O��w���W<����n����P|��4S�|եq�P��W���US��/y�㼢�(�Fڪ��%Q�q(2�j�8J�!�;�UD74
g%R��Uj���װd���r�\���S�d��gm�>ig���/��-���6he��ގw�w}o�J(�փ�J&��Q�*�"Py��G��%�ߥ�V�u��r�����6�m���5UԪ���S�U/v5G����Te
�W�>5��g��҃�}�i���E(��UB�a
�MQ���Ҩ�mmUZJ羾�Ϲޕ䮴
{Р�Gmj��U\j�ڪ�UG�Zh���6�V��3�����j�� |�-���Fq*�!\k�4�Q3 6����B֒�@.��޻�{�ߨ:��+M���U�U��P_aA�0�Q�^@�Ɗ��+mPw����k���A]CmQ��>j��V�ݕTB�y�P�ĠɉUG�%P�B��q�_�^�
��j��P��j���R��"y<�jڪ:�hR�4W;��^s.�Ϻi��r��h� j�5U�1�U��@�Qցh�4�)h�Q���e��1�k��h�U��ǥ�U�G�UmUh-h��q���-}Ԯ=���ˑ�Q#�˗k/�_6��o�)�R����5`ב;�*Ĥ��%F�$��u�W]R����}F��u��U_�hQ|�(u�:�R��J�EWP8�����N�y�*��i�UԬ5A@�5F޵U4q*�5䣉G����G��mD(�q�{��y��Uz�Q���W����Vڣ��Te(>h�!^j�%�!G��G3����!�^j�mU|�U�T" N5Tb��Em+mQ�X�V�GZ�1=��ؿ��9���6��u���QFSᢲ��Zy&aF�+(6�a�G7��������Q�9�TC��!Fg���5UiU�
����+-Ue"m��u��>�7�0�y�Q�+��ZJ�ܢ҂�4Qg��(��6Ī�A5
�cTi�����{�{�Dk��|�Xr��Q�@�iA�9�Pi��B��W���U�MU���:���y<�Xk�U�e��
�h��[h���>k�Q����n���+�gٽꪎ�Q�:�F����	��<�r�4ىG��J��C�G�5TN߉�����M�mY����Z��LV��Z=}X���L�Oޣ��3nZ ���Ӎ��^��w�����>ڪ�!Xj�)���e+��A)���i/�UhԁĠ�5A�g���|�Jrm��%F�����u���%Q�*�� 4V�		EN�F��ם�����i(�%UR�iU�|�j��h���u(8����-V2�ƃ�Y��Ok��yڪ6Х��Ҹ�W��ʪ.]O~���i.�v'G�V��W�#��~m���k����E/��z�Z�+\�� ���[Wg��3CyT��dY�Gn���̌'K8A��3���Y�j�D^w��U�����ӽFY�Hl�*V���+�=���Ԩޝ���ǒ� ���d����Y>��}����ҳ�-���Z����� F�8����c6(Z�
Y��Vs5,-�͌�Ĭ�Ћއ�Z� c��s���*ɂ�5Z)���1r�R��u��c8�����0�7wG���8>~.A�����{����Q���z�y7\�\����c�8y�������:�lOWL�`t2I�jw)�:��Az�����0�v�
���冯pw�=��}�����J8�w��	x�6�Q��m��ͺ�v�\G����o�R�]t[􉦯��6�W`k/
K��U��2�v���X�s��k�r�hl���r�Kɑ9�<2�nAD����uu�̋y;+0�J�K@���N�>�Z�EV�Hx]3y��u��u�X��L�����U�� ^1�8�ji~������?�yT�1��I_��coA������4�W��%�� ���YC�>t��:�(�� ��zd�^�+�!�)�;�q7}�=��ß !}�iC�h:S�by�x�:18>�Y,�]Z�EB�ѳ���Eu)}�I
\Cu��χ�4N���?E�h�7f.�=\�c�#�v6��/����|�x��Z���3��͖+����6��	��_����� +~{7�����z2�nF��3tSױ{��8�F�7��uESA]Ya��W?�!H���yB�ϳ�;�W�%o�1�G�ׅ�L疪_h���ǆ�GRܡ)@��+]��U�����W?	�ɴ��ٟG�]�Rbu�.[�nkt�d�W�|(��]Yy̋';�\r����	�}��㢌H�stB��U���Ǐ�cf��9Q\�'�'nfѺ��`�p`����4��o%���5�eU���szd@s	�w�����.�K6��q�n��>���z�b�&#�� �`~����+�ϖ���~�V�;Ԩn���uSa���J:�Y����ɁZ���K�L�B'fdZ×��,�ʺ��������.��:#:c|��3Wc%f�n����^�V4����)���|冨5�w
�$��,e�i �#����L�٢�A�t����/`�����$ ��۲�۽;R�7���6Eɜp�9�J�ť��>�}Z�=�'�Y��J2����OS�]Y�Da�zT��A�'#��G$MI"q�$��r�2+��t�y��޲���/���2����>��7!cC��$��^)�"E�LbD[m2�4�e�a$Uc$�r�eʒ�F�n�Qp˖�-D��.\��h�+���[x��$���r�ۍܥTbF��]�[HSJ*�JZJETn�V�QwmP�DQ�D��n22$�i-�-�I��,�[kH�G�.�Gn	�$�������(���KNw#`13c�k�g�ߴ	n��?����{�|�}t	�����쐾K�czj�۽,\�z�H*\�X�lZ��t\M(�_�����t�䷪�{�d�>�lt�.��Z&�~H�-�7������܂Z�D�0�L�z���wnl���mL��o����E�,����`ޛ��E)�Bs��v�-
"�g����_�E���vm�/���_-����,�5wX��T�[-o���)�ˣ���ņ\]�;F�� JiO���r1����Fw�.�Da)u:U�����NV��Bs����K[��{+���vX-f�oY�Mr��/r�N�	�=^�}ס�WO��]ى���Gҕ��Vt_����}�5�V��ij�8sov�3���z��|��v�%��}AZ�(�^���e�;E*�]_��ݾ'ÿ��6���-�J��n���b)Y��z{`-Ncp��lh�[+�oo�0̩Y�����M6��\%����?�#ڼ���ŤH�IQ;����=5����t#z�w��.r"�Z�z�*�s��5��'�s.�R�[�ۙ�{(�t�x�
���R�<��Y���d�G=�vE�M��h7��~^�A��>Cf��.��x
~�aGgy@7U��\_���Ϗ�R��m�=:C͘��f��o��H� !�9��Sl@���Ђ�Ժ�9�6�s���i�?φ��@��y�ƞ�p�8��;��`=�8!�Zma�;D]B��t�)`V-��7:/��{�:�����ZM�k�2nP��8�����iqN�Oko_�vG���E��z��i�\�FlEN(m���ǾF��]�$��:�&ӹ��?L�_�w����r�9����o£�̬b?r;��S�)���Y�'��p�麲������W�V�m���ei��k���BnD��c���7�y��e�x�k��q��yW9Ӗ,�Q������g�ڪ�k�x�s�`��zq�qL4+ξ+�! w�x��Q��Ǵԭ�x�IY�;�2�{L��������JGw��>��P��@��F2�:8-����k��_�x������Q\31��غ��r�쩚z��-�L1���+dT�����RO�����[kՇ�?��ڏ?8蛢�w`�yԛR�}!�Rѽ��{�B���_����d��l����ƦX	ϧ��j*��3�o��ϔ���O�cTRݏ����pDiy��U�s�y𮆃��y�v;4�)�=3B��uL��Y��U�2�̜��Uq����]!yCx�9�߹�`P�� ���,��}��M{�w�eCy6wK,(��h-�ɖZ�W��~I������oW|����&�LE�د���9A]'_��fᷧ>�o־3����t#}}���<�H5^�쏮��)mJ����?*;���-�#��W±]������y��f�M��� ~��[Uk��1S�U� �sc�l1U���G�Nauz��^����KLKtdˮ��-���I᠔�7���0mpN��ܹY��������-�����7�懽��[�Dx�W��ǖ�S�x�%���˗]��ז5o�f������{3�X��}�޴�����o� �Ą? �ڔ+U���qq��)�T�X�+:��Q�9��PخF��ֵ]��⻅Fg/[N�.�q#�:R��\>;���ЬC�7�!�[8�e�]G>�n{�ـA��Ѫ�ԗn�Q�v��wv+Ț�hd�jK6��������K�O�g�G�.�^;뢛L�y��V���p�M�dW�RzT�y4�hw���'�=簢�R��}�+S��}{?�>����3�?2/�I%߱`��;�b�nBˋ8s���Sە>$�p=��0�����6���토�8/��\
�~}�=�M*yʵ�����w��c]� ��^'�o�X��nc�s��,ђh����]�r�u��������7vrI�_}_WͶ��������g��f��c�����w1ӗ��3��nI�a�;�����G��}�bCǨ������t��k���ݠ�2��J�Ne�Uw �r-����a{�1��Ro��@�ւ¥�mKj�K����"��PO?J��vp�ѓ��0�X�Ee+�jz��r������bo
0^Wmz�p�lBY����ɱ�ou��Y;>'CB!�z��h�D�fP|�%"�k�(�J/T�Ho�b�ԁ�����B�j���l��C�Yr���TD׋�ج�����?T�"������F�F�է��-��z,�6
1�+��Wڕ�l���|u0e2�rV����<!�P}LӢ8�r�fZ��iZk��Vܫ���ŹI1�#�c깸�n<I���צ����)*upnk�W}���+�5\\(�8Jn��Q¬��S��k9Jw��/d�l�A�u{3s#f�T���٧L:F�t�0�(��nu�ђ�7�w;1�K�&Ѥ�
qeiBX��	�Zр_�$:�î��\�9����8εp���U2d׳Fr�n9�	��Yz����_�/�et�� ��(rYڋK.�g'[��U�pS{�3nd;F��J`�&G/+7�٥f���ޔ,��XE�:wE٣f�Ms���f5��R���	�E���$M�"j9$���u30δ�vDq��m��|�}��z�[����Ew.�bE11�XԖ��-�Y	!1x�`�p�2�n�-�"���c%b��F�$%��Z�Y$FH���H.$�crF ܹwTTmń�F��h�bU�SdX�Z�!m���m\#L�##R�Z�$�b,DL0�&%�kM" �/� � �ik���*5��K��蟃�����{��Pֶ��^T��Jn����m6���P��Z��߶H��{��^p��P����ʽ��{��Z���q�v��Xl�g����,HY�`CHK���k({ �n��	Jh�Fpa���ךj,���^�R�-/���Ν�+�|��l$g�{�
��N%�uxb�{���`Ke8�)*̤+����Q��l���W�'�����[�u���8�4� �S���@q��(�i��e�������'jF����[\)o�3�5H�o F������*��둩���Tx�#�|u�"�^u��,ѣ���?q�)��x���k��W���V=��8���hC[�/d>;\�[��xen<rF��s�qf�=�Z�4���A<�Z�=�+�Q��<���o/V�[�[k*���V��ryǱ��Z��iʗ�Ɛq�n���V�4�D�]������aC��U}_Rm3����,�_�w�(��V�RM������ZX�1s��Iq�|���@�<J��J��g�N�*�NS<�x[m>��!JeY�N�u�{Q��Y,�}=� 3����}�I�y{��vr�ԗ��sjE�����y�^g:�c�u-�5�x'%���ժ����W���,P�/������xU�z�+,V*Fahȣ�� j]ƫ�x�	V%#�Z*7�����M����ɢ�Ŕ���kx�����'}85}�Mtt�_���Ox�o��^�U��o�l���m������{��nX������c�̍��V'��Y�/p����3|��_h�)��i��G�P#�;5q���� ���q5Hފ���ᶰ�eB_d�����bK�,;"��?G%'mU邖aLE;V-�<��Lr��	m��҃���N9?����m��śߍ~���5|��j��X�^<�#�:�������E��[(T��E*�봼E�X�ً���x����K�����e��Fi^/�g�cf� y��Y	̜y��9�ŵ���aȄ��({�9��\��
����&9��!�h}�=�>
���g�}Quk#׿�5�I�8[�*�y�9l �j;��,�F5e�}��\��������m��?O�њi��?r�ER��J=����<������^��E,!A��������~��l����#XT�eOG���eY���I
�\�Ҹ���7 �H��X��3_؜jGu�ii�����&�uJ�iy[��T�#6��H�x�]�Sɚڏ��hVO���缳��������M�#�F�ɧ�c�d�׳�q�qt�Ÿ�|�"�Ű���Gh쁲�Q�ﾪ�����Q����]߷�J��(��O*�F�Pۇ}�.�=O�o!�gk�?��Bc�[�v�����"�M���Q�K���˹*��}�b[~��5�Cu������&�� ��~��D�[b�1�Xf{ԎSQ4I]�'{�A*߄���Y,�珻��ΰ������^��Y�]
ڌ��9��P)	�ZRZmǏ7�[ƴϤ�)��������i�~��}yF�W��o���1����:��ْ^l�A訍����q_L9ͅ[��#����~�\�r�������As�ӎ�ѡV�(��苺�/Aٞg�����B��~�g��GsC}�EC]��d^T�|w77=���f�=��}�w�S�>1{������������J�����ԯx]͗��o��GQ\")W�����(�:�Q4���UU}r//��^�Ev}Ǻk���ў>�/gBB��1+��K��T����r����O�_� �}��ґ��t��뺞ԅL�1˭��<�Ec�^����5z�xp�5��R�h�Ə�v
�93�j��Xu2l�kj�oOy�{�w�r��<5�G�*
��
�X �{}h{��X��x|+˕cԅ1���_�x.5�ּ�@>}{X�U�5kC�^�W�k�S�?g�<��X�c�%]�9E��V�;z��ǠL�;nZ,4����!��K��;�UPW9�w����]F�L%_.��t{���<STe��R�}uB�(��b����j����b�Ǉ�UȾ,բF}��
��PAHo+��l]/e;��x�^呰��wB�eMݭ�5Ď&�	�Xl�Ʊ�nw�N��>¦�<ҪCP�pƧ��{�����]�0�2���8�S�fo�ލ�ԩ�iZ�a<�5ס���Cٽo�5t*��%������Y�`���F�rOvWZ��y�i�e;�����q������԰��y�$a\�Y*�Y�3;�c�%n��K�|�o�l�� "����ck/��	5�11;n���7���ܫV���&�����h�/8Z�N|��@�\���T�d��B�v9�6�
���Z6�ŭ܊�� �:�}:�fYrY�
`�������/����;����W^'���,�M+�C���]�Q\��(��-���i׎�yv���[�Y���w;!��OZ�R��
�� n��=���W�=��;,3���l����S��kp��~bH�r׎��uu�&����DU�����	+:�Yw���6�QPC2�R�=Xa��3�.ql��v��s�-mn���n��Y?��p�G�5x^!��՘{2[`T���eH����{o�T�Rm��������wi��M ��rk�@���h�vS��/3#��Vv�<O4�澙(.�ף��~뢪���e�;%v��t��4�L����8N��V��� eEd�R���	Q�zC�H[�D�rI��vؖc$&Rظ�~8)Lܨ�c-2�H"�ŘH���dnE�H�%C	nj�ŗcKr�pa��K��R-(��BR�#d���J&$�.��B�-j��R�1�ش�[x��p�ZJd�
�	1�\H���%��LB������6�Ɔ�L$0��]8�$��������.� 0F��&*]�݈Պ�]��\��1#v3m�%]��Y�B�"I��ƈ��AqS���k=�I��O����si��&	�I��\�;�
 �7�s�e�bMc�����U�ց���c�I�>c
�G�xxV8����[�b�g��+�~�&��M���a����{�v�4�|�i�����7<�κ��n3+����Q���O��}gɟ,�tV�T�8S5�iz�Ça�����w^+�� �J��<>���eU�־���l�kE� �
��σ([:*��AiU���������*4� h��V�(���¨�eÖ'�뒽�i��ͳx��߾����-�2�Tˠֺ��z�\m��M�Ћ��^�2��<�㜓mF����(�{���x�p�^wu��+Q2��k����8��|�PY[zM�ywF�Ϭ�|�Άǵ�<Hy�0���'�Zק;+������o=��ΕӲN9z����_17�voz1�ZOvu�;���<iW�������7��ǹ{]��p��*�i2�b[Ͻ�ǝg귯�4������!�Z�r����.��]e��k��.;�]JZu(�9����>��j��<�4������Z>�u��eq��X(V㡓P}1��^4�
xtW�Կ~��ըǃ5՚�u'�����S�/ƶ����=�����oY���uoDWQՔ�N}���|�n��W���u����*����X?�3-���R�(Q�I�j���y����k|���f��[��b�_����o�5�����+���+:Fib�U�D�DW�޽ԯ�)F��q�n����5�Ӥۓ�y�;�C-r�E�KN
LѯVC~�Y�p���u���e:�d��/}*������v�#���L�T��ƌrC^3�����sR'�u	�X쭫�^�=���{���1�\|��ǉƳ����O��|=������,l�˗��I9ݽzl"�W��M���.�`�9[&�,�̽�������[g��n������AVq�ܑ�ncݾr(n�������nP�UZ+���:��vW��Z�:D��]嗟Y��X��~�Į�]��X�ƍ��׼���"َ�:��H hP�Q��4xU��}w�8w��!b��(
�i��,PvOg(�j�����=���</ƫT_1WZq{�e��N|n���]��f�];����ޞ���'[O�'$#�ȜIs/�)x����J��)�ަ�"��H!�3�:ư6����κ���:�_Y��Y��-ܻr,) �Ţlʝ��
�h �s�i����U}�:q����w�y���b.T����}�$f�{�]v�#�����W(a<�52Hk^�f�g�m�!��z��5�ͤ7:S����N{w�N�N�ܮ5���ף��*Ç�sw��u��4�������wq�{y�}�<�X�>�OV���J'�_(=��z鎇���*C�X��<)F�u�^�ޛ�lz����\>�~����o�/zJl�cQ�μ�#!q���
c�/kmgw�}34�!��f|���7�׭b�4_����.TS�v��t��\/��ίz���t�R�\�n��2��ʕ1���(�s��;��_��%�4����c��w6p�'y��޷^����i�M�����1ۼm0�cI��p�FiB�^T�@��;�y��5Wȵc�f�}p�]�X;�C]����J�`��R'�AX �������X�}�*^��3��J��X ���z���,�Ri�j��f��y�eq�3�13�^�¡��p��x�;��ݝΥ������u	����J3��|�Gw�Ӯ���B^��� "�ˍ�Պ^*���g�?]�����59|��������2�b��!y�鼜�r�_�Y��n�l�1�6���_W�RE��v�q�~f|��g[�m�?�Ljv��Ϸ�����5_� ��� �_4no?h~��n����0�(j��R�kG�簧��}�{�� �����3^^4��P�����!��M1î�<��Ë�s:�}�o9�-2���or��Yz�N�ϳ��a���4Y��>L�_��(;����*�:2�yr𥆊3K��^���f7܍@E5j���
�[gGњ���{=׷�]p�h֏�C�?�:デߚ��ؕ���_�[��S{�B
�i�+�㛟��C�w`Ӌܱ�!s�����*�]7vSrI��Uo�9���4�S�iZǡ,���^���m!�*�%˫��ϥ��� _���F�'=��gQ��[ď�0��5b 0j�{"�3'� �x}�Eh�
��(T�Cv�L�8p��Π�&�ƶ����֨����C&�\r�q�9��zoF�=Gs���K����)�M[�ʐ���U�x�p������~x�y=�L�[��^	��|BL�K�W�ػ1�]-@��w�����g���5���&�~9��%��&�)�,��}Q8Z������I�FU���'�+:"����UU6�w���/Vq�n]�������Ȝ���w�c�-]���޿�vkP�g�m����5�͘�f�a���_��.��*#cº߱�Q/�v��UHT�����a�J��<�����Ww�q�9E��W]"��-��{��I�)��QV >t)�:~xp����M����f��m
^=ko��i��/ۗ�*q�t�&�u�zz�w5�xx��n,h㦬U�.
�k�{ʰ���}}������y�J��������^��6w<=�^�^��\R�wm��k;������7���I\�} Of���ɆZ���}���W�����ϕ,Ww��uc��<+:�s�Ѻk4���SǨW��~��m��/�̭�KƬAl��?^D��P��p�> �m��6��UO�3�*b���������ܭx�`)�5�q�UzpS��GۺS�ߪ�A�c�� �A���Ϯ}?!HU6j���T� o	�ŷ���
�٪�q2�̢�9��������:�μ�<C��j�����,`�6��o���}�5��<��k݂�2�p2���ٛ�I�ߝf\�}��!�BZ�u��d�VF/Y�[x[YyO��ƺ�V;�+@�V|�����E�(؜8�H�	8s�R����N�Q�33[g��`��v�j��Jv��0Q�
�v�_&��G�2�6�P@��	�;Lj\�����9��݄g��<�-��Dr�\҇��� U���Z�24�l&$����¤w��H�L���[V���pپ��2]�-�.�
���f�(�X�y�m���T����{\�7�B�j�.�Is���y�~�s�~9�`�l�+j����>���g��B����u� �He��wT�\�����2��顨�n74uGB����E�H��۫x5���z�N��<��GqT���*S����tp� ��x&�Y��mgm�N k�c{/~:��U�[�
��6q�cv栍5�6�w�
���_s�X�S�mu�}�l��گ�\�Y��s��w(�L�BƄf[��cq��f��㴩�,�\��'A�G�$��$��r&"�\침*HK����с��޻���@�@
�
-��b�\n]�-��b%a&&G�hU��@��i$o,-��L0m1%�l�b���Iq����1`�c�v�`��%�Y���Ae�3coB�܂3mԒ�j8Zʻ�e�Yn�a�[�K.�n�wd�Ai��2۫KH�1krV%�B�$B���X0dT�KwcJ�.�F��l�\1���$"���!�7r�h\%��qőln�cq1v� �cc$�[����0ƕZkI"*�AY"Ӌ�u��8�v�t�kZ�?6�{���%Z]^0ĩr�(bs�_U}\�֫=t���u�j�d�>v������kפ��^�]�|,UЙNͻ��lu��/��Km=�i�����ܔ^c�d��B���l`�	���=B��M5b�NkXƳ;�gٍ~��W��]�z��Yk=�TٗV,W�?W�i�T�O�*Wy�=�fj�u÷R�ק��/�#Y��h������1U�C��Ӂ�N�P�!שz�滽�������L=��%�;��:�M�{|�L�y	���P�a���?�a����罙��
�@�L�.�[��[籞�ڡ���0㹣9��Tw`ݻJ����,��}��[�7�{��q�����0�0vV�nQR�r�o#�3�Õ�d��S�=CԿe��S��Wg�����°~F��W���C/Ro�o>ν��=M�V�";�]&C��w���s^�.�������M+SЉ�I^Υ���s�{�޻E�ww^K,���&��e��M�*x�z�!�`�����6�kY��`�������h�Eh�T�R������u�� |~8ho�W�\��
��cv��
�_�g�PPw�_�;9{E��~��B���-Q�%���Iyۨ59�]��$��f��ҝ�V�q����}���U�\��:L�/�_����,���\�7����ږkо:.�A��X
��K�/zϙy���ι{�i������ne�N�+a�v��^�D�U�Xb��F���c��TGZ8V3�_�k��}�;�p�5��m��V��|��gs)����i��{����k)�Sn�����8us{��&��͕�C-�,hB��@
�8�v��c|E5�E[�j$#�J�e�w�1��~ɧ��#Z'�_7���B�
��������b�Qb�1\��5��ޝ<B��n�?uԼ���^ō�;����Ŋ���*�!�?�~
�9�s���Hz�Y�	�ޘy�0��[M�MN���d��By��M�w+~�����S;���=�+jƔ�5	�g�Ϛ�����dy.W���1`���;5��`��{�����[�6�M'_=O;�&����3�y�+q�,W�|,xWztN��܅{7���w�쬡�ù�p۷������� c�GE"j�+�i{������b��}c��P��|��Y�C��s]�fNo7Gqp�x:����J�c�D�o�]YW�w�����s�r�x?�f�)ѫ:Θ�a��i�xa�Q���5�@�4�}�
��{��V�b��D���%m2��j�z������k�-X�՛����������U��\xs�E�4�
�����3�6�R�Y5|�*Uک3���C!w�I߮}�`�>�
ѐ�2u3ٴ�\y|��:�{Y̯'_nV���X)x�����߳һmx@EЭ��jǇ�!5��M!���
��cE�*Zk��k:���k׽��3�i��6����̼v��]�	�Z��_gX冮q8�٦���>��+HkW������ss����W�ح��5��Q��`b�Sm%ܻ�g��4�ڦ/q�3�*�j)?��꣜��+H}O{�WsNX�[�1�]�~�s<�Ɗ����1\x�b�?e���pk��u�va&g�!nX�L=��%λ{u��8�޵�v����L�cB��ս��ұ/w�Rυ`�#���g/!�g�,]Q�m��[y��٩1p�s^�����篽����5涙n�1�R�W
�:({ٕ��`��x֏��Gp�ɈNg�׷�mq;�h�z֕���<��5����~��<E�or�׎K�������~Ú=��~ݡ�r1a���Woiz{��ۂ4��]*\īJ�t�X%%6a*6��꯫��k�V�*CW�jC��O��R���S��8W�s��%hz�^�x�k7�x����U�̮�k����{�ب>I�q2r�׽`�	!ha��C\�q�.Ѷf��_{�k�t�Smv��3��ii���$������օ��+
�}�?%=F(<�6=�A�xՉB�9|G��T�+w��n�V�Ԍ�k�٩ćf���
�p�hRg�I�P�T�֎X��9pu�H���ߥ�i��f����~����P/�%�zs��{����Vf���l��G�������n
��"�3nZ $��`���ԓ�Oﾪ�9�k���a>>�k�I�U�n�	��������t�
��,����"� ="!�Q�uS2�῍��w�Y��͕P^?>D`�ɤ)���>�+�����������j.Uf�i�B�W���h�?��w-�W�V��|����ؼ��瑱Lf����)���𫇇�xn��|����n���4�������f�M{�O��g�m� �U��ÅX�~�������Lҳ��
h��wT�f�׮UԿ��>�.�W��r��o�SL�S�ϝ�ӷ�6��X�9��dJlc�Ԭ�i��Șn���Kn}�J��%�O���y�pۿJ��㲸�q����/�����OŊ�4�}z�Y���<�o��W�� ~4�XxxU^��3u�o`��5T��!��� �{N�8<�v���U(Ab��0��ԃg�,u{=�/m�Gyu����<j�P-X����*v.���`P����h����,fӷ�2_Ԅ;��5W��8h.n0��vV����Rz��/��y�S��c��5���|�N�9�a*�$�=5�N��O���7�7o�;��&e,���- �rY<^�E��M�D��)x�$�Q��_W�kjI=������/�1�+�!�$��>�׷~�@�χMg�!�Ы5�㦶j����{X)�+Eh���2���tF���4r��^��+L�dՋ1�:�u�;��|櫭<�k�oK����w�s�I��k��8V�}�i�ɧP��bJ���Lvh�z�.������엜�2s��;�o��8�a�0�{e�e�-����{&}�k|h�E��|t�+��.��=����N-.5��b�|�+!��������4��M^��T&頞؞67`륐����  ��}��p��"�nQ3zRKv��[�0��E[kcV�i��@g��x�L���i�Jt
;6����ÖY�1�*��$�9[ՠ�{H<~�-�^U̗V%)z�z������:-V�u3����L�{��Sj��}]U��gܻ��4��O2����m�7C�A]O��%��7i>yW��A���ą�ˎ��<������x�-�hKMsdQ�ͅ�f�>}Ň��7�-��e<Xv.*�v��Z�b�EMa>�l9��iԶr�08ܦ��<)�8�̹�,�x���B�Z�qȸ��ӣ������5t8k����V�Ӷc�����E��v�Į!{lj4���[-�:�D�nM�'_n7���f�T{��y؆�b�K](o�N�חZ�]8���p�zYV+OW4+��s"\�v��zuw=rs��l��S���T'%��^�Ш�W�N�ho���*ـ���c-�j�>1S���tXl�%�.U�7���7��I�%n8�8���v8:9�[[Q�λ���P�U�A�I+mHƢ�j�Ȅ���&&,�L7�+!�J���0��1%�m�$�RH��k�wwv��7XL*-����n�X��b�H�TK4t�I&>��I�!�Hw!�mҋ��KlQ��v-���p�.B�J%�D���!�Ì2`Xȭ��ZF�^1m+mݸ�0Lq� �6Kax�+,K�K�EE.mW�6V&�Wlėx�����Ym�L㙸��4[�5^ 5j�J��>��������s|�$R���c�?M��������w��w=���t�'u+RDw:Lތ��9}޺mۦ��WMB�lM+^M��7�s����i�z�;8�����8U��tW��P�G�+�h�U���`���k.��o�� h沯mdz�v�6�Nono����J�{�54�eMA��$q�̞�F����S�5���y� ���/��盰[U^8���Z�)�u��G;�?�����u��/ܘ�X�������!+��f���D�sv�&�̲.]s�p���%�������z #�2�(R�����M�m��>W���B�]g���S
ϦG�	.�8)KZ��=v��t������dp�|�0Ps�<��&�c�������^��-Z{4C��o�n{2fxo>Sw1�}�<9��6�x�#(g�U㗻��ȝz�Y�t�S9_�߅й�+�|���&f�S�k.�P���BzI��}�g�=�g��u�a<T���W5fq#V<�yy�q8j��j�f��!�lO>L�x��wܜ�y�e6�c�T�t�3�V�~>���}���ߞ
�^6l]٢y�9
L���
)���$�0t��qA��D��s�>���#���r�[�Ϯ� ���w���+p5ן�!�5�ց��)��DX�<�з����-z�ɔ�׭kr��k��3�o�ҭ�yf��<*x�
��M}�����G�P��iY�2Ǽ~�@��&{�m!��f��+�ئҪ~(T�2��{;d��o]�q������.5:�ZW��j�����y���4~`�8!^�8uQ^y#v�z�;�8�� �����훞�q�o��B��X�����3N�˫W�|���k�#�~�ôW0�l��]1?f��®�� }�zY��HesI� D3*VqE�?���6ۯ]~�ݛt��m�ʖ��R*q}��`���eX�~�`��/��U�5t�ƽ��ؿ����Z9�ji��MRm�j�J޳�ν~M��ݕ�Ӥ��d�	�M�׎�X8ju����w�,V�B��)�?]׺�p�O���y�3ņ$s��P�^ӝGj{a����{lS˪��1Y.wN����C��mg���ux[��A ��xy�E�[�ߍ��Y���O�~���� +���&�b�Aw�#�5�pnsB�!�1�����UU6�7�����x����!��ަ!a^��V���jo����Ҳ=������,�zu+y��-�YDev��܍`��ݝ� �����fZq��p�QD=I)���;0g���<7˿��U�䷕$lg+��
~�Ϲ^�ɽB��г�R
��_ϳh���b��W�a�{��
�8 ��"���ܝ4@yK�"s�X�"�ݫDEt��M�'��}T�l�c�������������=cm}t��q�x
�&�z�:_���P�H�Zr_�ޡw�����޶T���Axv��Eޤ�naբ{d��ȉ�����{١�\%��*�i�wd�W�-�E�|ZN�Iu��]:�H=o/)�&��I�tU�	y}{��J�cu�m�����p-z;�jM���[�8&Lh�74q�+$T��ʕ�NO��4۱��5��	��m��#f�md[��g�-�-{㾁�SP�b�'3G&����׶珪Ot��ZDH�=t�$�by~��(-�'x�+Y�2��އ+kk�yj��\;l���������w0�::Xw:h���5�j�t��f�f���#�e�̮����Z�7-ލOr�}ŶM����Ӣ J���;��Ko����-G?������w�K�~��^�삄�0E��M������`8B};.��=��;��7�W��M��_7�VQ�i�:��!�#v]?>��2�}}��皨�F�ZXo��K.�}@c߲�C��,U�dz'fG&��}�G�s2��Rt�*YZ5,�5���U~�V��t��$��<�kݡi��gh�i+��b�0\�Ip푕���k�yd���#`�E���˕��ӟ��}�Sm5_��w����!5�+��sC�&v�ُ5
X�qԝ3���ﺊ����=�i��.�:P�X-����O��;.�XcHL�ߺ$��{��>���W��h�r�qv���
�{;�\�#�=�Xz�$;�}�$� ������U��������37d���n�Wt:/q��Rn��e�.fa�iWCC%%�X)�����6���/��"²�z?[��JٵG��/�8��x��B������m��=���6�m|�T�E�3�}G_N3E1��Va��S����`ʳ���r.�Y��h�O�=����s�	۹�1z���TG�
����rr�ly��y�=������AU�[�~=cذ`U!�62���uo*fk�a#i�y\
K+��*��{�uI�S�����W�eZQ����.0�c�쉀g!�6A��L��7٩v��/G�����muG�[h�[�v����ۦp558tĊ��z��)�=�x7uú���;(���;����*�P�h�-��L����Ҕ�}cM�R��|�N[{Wn�S��S(�DVٺ��M�sCǠ���,)���ٵnqzI)�S�-�G6��,PG��O;Fm��+�׬B�%��ų����VE����c>���� ���v��i|�P5+)��qm��|u�E[�B�'B���T�p�]�_T8ܓ	8;J ˸XIw\6���"��P4S�}@��Ÿ�[&w"�@���j��U�'����e���3z\UeP�$W"�lG!ˮ�[t�u�	�33{s*�bB��w�X��dn�6���S.�v�=�a4���]g�E<Q�����Ƶ��f�9�u�4�͛F)����P�\��y�HXN�n�X/�ds{�
H3�rH�Ddi���U�G;�,���	H3(o�:OP�HT��%Q����a�rY$��[	n�bXY[,C��Ի��%�1�!���e��.�����mb2�X�!`��e��@�	2Qt�>!E�a�7�Ċ7ڍ�$�$n@k
�����KE�.][�r�[tĺ��X�7tݬ��b+R���v��]�A%��62]�m��-I!$��Kl�EH�TM&��C�L�A>�6�(��a�Z�?M08�%��$����H�,��ݔh"-��{9/R�o�|�ث��5-�)9$����ٟ�+���s9md���!����f׀l3-�����#���*t�b۷5ZeՅ��Cm����p��r�G�A��bǹ[�7�13wA�"���N�6��vF��+s�_�ڳ��A��B�WcIO9aO�H��*�
W���z�j�I8�#{�H-��a�]^�z����ؗ�R�qq=��i�,g��oy�pv��ez��a�r��)��M�ۯǯe�E����������r^�,�d4�+m��7�i�l�r1�qن)��ʝ���[��^��s�޽j9��0{�>��_ǜ&t��+3�3y��z����XuwM�{�]'%;�)T�Hz�|n�2����KS�c��ߛ�w����'�×V����sn����A��%Zj8���8$�B�Gݰ��<B34r����R�jI6�z�����WBv�t�f���P���=E��u�q:5��/?/6���S�c�[9`6��v\K�M�s�{��.�����yf^10�՟���[�]��5�1�]jO_p�v��bW[�tF��LE��^�^_�26�����7]z�����*�e���64�ӷ*Ȳ@ʙ��U�D�rؕji6�q���+�Pe�H>����x6j�:#��O��):z�njћ��r��Cj��������^3�$ `�ֺ�;��?����SM�#��>_;�}b-�[�oñ8�1�U�yE~3�ë�>ʐ�����~1y������ޱ�%�ð�F*ޜ����s!�����]���P��ױ^��^��tv�j@���7���m��:	:��B��J����T5bRY%��qĈ%�:�v� ��mx�*v=�n��-�C{�{���R���s8Յ�ȟt���6�՞�nj�÷gQ��<�ٿ{������*��(�z��gqx���]�h�u��9�����	�� pE9z���^�t;�v�w�GN�֫6MmU�r>�6�62��Np=��Wg_pV�I�D�1pF�뜉u��12KۖH%�z�l7�b�$�����Un�Y�������7��M�ܐW��d>��eFV�ZF�͗ �/����G+z���o$��yMB��#+�9Y�SK�]�^E��[G�ƒm̤}��w<��+���Hv�.��/S�̸�0]�C��y>oA�W�������.'݂�Oߙ�J����w��5���ѷ��?;��0:9P!�{5�����
�^���Z����I�	+���v���"XѺ�,�ަX����wv_A�\x���E��쏷S�·|�{��=T��]��HNv�.���<�z��64NB�H��$q����i�5{IU�=��Ep�����
ϼ{���7.$��:G��v�Sj�_F �/xvU+�v�̦偹b�/�9G�t�cx��\�`E��xl�o��p��r$5�H�0kg�N���/\��IGl�ꍰ���$v�<��$�n֥u�Z���'ҽ�~��t��]w��L�Oj��N�i�f��Jvα�a���Xn�"�'.�7��-�@��3�:q�{*h��ȵ]8�9��0ݕ��._��3[�vC=m	g��4���ǝ�O�8p�Z����\��[t�O�e!@P=��I<�e���E��T��8�(c�u�żkc�����p;͞"��V8;
S��q#��8�V3³ю�*�7�Ě�h�W;<�� L�>7��5�!�'������tHJ�^�q]`����B�;��l��v��冲�8F�����8^y��Y�1`�F�X�/ypsᯨ�TO���x{ӕ�ה����,z'WB�p�=k^�_��b�x�~l��J�&�5����\c���*�!$f��އ�����������w꾢���{_u>@���y��T�X�d�ث;�>�8��=מ��7S��-htr�dH�L�&���E?]���$�(RY�)G��j�v9���#�X>��%l/��+b��#�&������A�]���uԬ��S�𧻓�3ï.��c��3��\�*lʼS_�E��HL����{���,Vd�%�=�q�ٱ�-�7v�#@���L�kqi�I��tZ�)#C5�x��}WJ�`WK��v�[i�q�<�M�p��M�yQ��x\������絷s_�р�zd5�;�wÖv>=�7�ٲ�~xeM�.Y����bL륻�{�s"���P�N m�_�*�`�,jVrvP��N8�o6�������nX�586��D�8^�N����kw�\��=�ɛ�^n��4����S�]���0Iq�EZ�׍�nm̴cu��L[׉�J#�.&Br��ΝǓ�8�>��[�jJ�+f�=yI�w�Sd��_vui[��	���ڏ�NQ����*���Om��ס��C�
ʼ���g(������0���ނ��՗��$��vY(E��s4{��@�M��{)WRl8m�k�}jۭC�rM�V1��҄�{���3IrH̒Dm�蜒�X�'������o���͵ɥ�Km�z��\[�r츑n�n�\`ԑ����-�b���,mq��C�I#.$B��uuj]�mDS�jY��1��Km��[RY��J$�F춡cr�^�$���n�IV4�%��I����ZX��.%�B�.%�km�q-[X��^p7.�m%�ڥ[e�D�m�]$��� �8\��q��mZ�DV1�� �X��1q[H��m%�m��-�*�$�Œ�$�R7 %�wwt�.�]�0�EE/���B��^^�����y6�.ܖ�I |;a�Rq��m�.�?<c�;�vS��k�W�y=�����O:��l��Y���qR������1�IKw�2]����K(�}f�H�iL�q=ܡ��WE�
��P~S��]ҕ�bK/�,�vT�>�qP��0�c��Y@�Pʠ�5���c��O���P�Z9}�R�k�˽�?
�\���,_m�,�o����X>�&��]jEVo��ҳ�-�	$����^���Ȍ��X��p���:�dKd�+�ӱ����6��{����@cT$@e�em�D+�ǲ�l�u���X�XF5F����KZ������_��閾8��⮬~v�ު2���O{W�V�ټ�:/�RՋ����C�g����@_�z/���+��3�ʺ͠Q���`��\��W=��2N�4؂�^hƈ�Pi]3�j7e"��E�u�ܫ���;�z&G6�����=�v?]��h~)���S�
��(�����<��u�F�W.6�7���5yt�XUw���d�<T�]iN+��:W�k��ZiQg�b�K�J�PP�tLYkZ����ⶎP��ۄ(+n���[�tg��M����R�;7�!��HG�}���I��?\Fb�{:�N~��7��-kzjވ���)��)$xz<W��-����ݳX`�n�w緕.����H�����U�/��yϤ��n?u���u$�A�M��olg�7���ŹXcކ�ܤ}�d�PM��X��.8���8�]�5`�YQf�uql�6AYM��^�]Z�����e\
����ˣ��ӟ���w�$���$U>4�9�����fe��c/���v1���`�b�>�\b��6E��WHk�;w+D�I(���%���b�`�������"*k�^��6��{�c�pw7���j���6V�����#����7�Hug�M���c�9]�x&eR��åbş�^��&[�V\|�W}�������[׭e��
�N`yX��(5�%��s�f�:�7^'��[�V��5��=国dV}��Y�i���J{��2Ng/r�7�K����M��P��	�&�Yj8�M-7�|FXF^ٯY���[)��h��S멽�t������f�f��a�/�n�B�퉭������5��*�Ua������yۭ-�wH�ARB.�y��"%ʌ�hY��:X��]"5�{�^�V@�=/&��:gX�R�k�h��z�;��x=��۩�?dl�@�΅�vfm�!����[�ߧn{8p�؃��ae�� >�pm��\�Y��H$}Wt[�[�.���!W�K�ܓ}`d��{6�X�d����fWP�j�}$��AŁ[���CN!�y��t̥Z��o�۽=^�5��r��I;�P?]xD�ǒ(c���Ύ:7W���F/R�&BrS��x��;;Dg�ȓǎf'Y���ՔVkWS� ��r����m^3�QБ�1�9xK�b����P�C�;�R-2H%���H㊕\��/m�$��r���U<U�ߩ��Ӕ�S�_��U�H��/x��k��痍����:{(��n�~���=��2�!iu
v�s��pˮ�$Ĕ�,��e���DN���SA��A�~���������y����x]E��-߬���9b�·���_[��H��胪z[Ӵ�x燼��3��P�9c��AQ�\.��V=���;���nI	$�2�����}��}���C�|���K
巔r�fl�c��w�Vo���6ЎR��(cm>^I
ٕ�z=Z��j �5�]�u��e������#E'14��
>���`���x����F6�t4U�׬۔pؼ���|�u����p;�̒X��;�ЙB;�8���[�4�rX�,8>x����́a\[���Sg���v�GLO*VtE�H1_�����1��'�9C����y����6b��Ԧ�}X��G
�V����7���{k�fث����6"#���Bm�1�d�ȦBfV���սuk�vud-lz��6�;���n�s[�~�
�O��5��L���²�<���v6P$l���='�L1�^i��}~vH^��W�x�eJ\^���?;�o�l�Z�g$�^����\�im֓B��(��V��\\d�c����r�_��x� Uv���P�	�︐٬�޺.�4o�dL2�i� �Ѻ�%l�a��E�C!�w���yE��SN)�!�9�/�XF��S�Μ:���Ț���ug]r�۰Pi���%�Y�h>oGM�����&e1{t������ 2ij-a�N}@,4���@3Gh�WS2�x�ٵ|�K����uf�i�x*y�s�r���]�)JS4�c&W�5��S�/���z�O�t�\�\�ݙ6�N��M���͢��I�4O9�:�G9�ɜa�K���W0�U�%���<�+�`�>�OH"�HO(�h^%�P���5�����ybUr�3Qb�<��L���b2����o^7J#Ϻ�VN�J�/!�s�dT�0��*&���bd=[��ųJ�hb��#"r�^�N�7 �&I"2H�$�eq�F�^*{�l�;��2�>;D���r�sw����őDPF��xYPq	X��-��c�QĂ�Ҍn�wpm0ۆ8�Q0Ғ�)r� 2�,E�ئ&10���lG�ĻeF.U���DLaF��*�H��e��˻-H��1"�dbH(�L2�v\�BL7l-,KKY.ȴ�b�M�*�����-�(�"8Kj��6� ������0�R�d��h���Q*�|�QĚia�����/�`7�U���3s]�*: #~����'ҍo�᭪��FL���0^Y؄�Ã��)���fT�gTˮ5ߴ]xG;sP�~O�zqָ��~2��نu�U^��p�J[����&�hM�a�t�㾋V�ZwME�����Һ��rh�Ȼ��Xީ�����oW-�>���L�۬%<��-�����i��X7q�%K��C�"��ueH��C|M����ǅk��YH����Q/2:�C��Gi��01�L�ɉZ\)P^����+RrT��&k���or��w�i��F�����w��f��H��
"B�i��S���q�3�;W�q-���&,?�EOM�W�s�n��v��ށ����]�W��kk����o7:� �jN�jﷸr�������x�CV%#�Y*7��Jo���oו����/��Ժ���!£߼�ժ�Z_�3����k��cf2�X_�t�a��M�t#kV�i�p��[w��7�a���,,�`�J��^�Y��P�8o�DU±��j2�H^{�FNuk�V"�5�O��v��t�Grx����ƽ�-����7=@�}�*;�M:�M�I���=�۩d�Zu����V�x��l�OV�:婼=�D/ B��Th��=z��Ѹ���E��T)�J���B�b���Bb���;x_�ʤL{��ݤ���7��c�Q�.�w��;E��g_�U�y����*�a9�?]-C����4�$�#Y-&]�xo��}.��}fq%����𙏼,�}�ʾΓf�9�4������[k�q=�ѽ����Ǭ�i�ר�ܬ��I$��P�.�Џ�+��Cyv�F���z��׽�N�^��d*�]]M��{,�
����~BkVv]ּ3=�7��y��.�^��[yv�;�{8!Fd��7Q��9�y.wN3&�5��]��a��>��T�uz��ß�[�}���z|Z�uŽ2m9@<�.S�tў(K�7�*$ԭ`�W�o�H�@�ٍ�}���ua9����o	��`�w��5�@�4�p��\/�A�G����2�w���s�<�Sמ:�Χr��Œc�u���k
h2�/m�qx'i`�sr�����������9]]�2T]Ye{FK�-��^o�*�۲G�*Z���Y����iO�G����;�t3�!�F)��לo�5��9k�B��+�U3�Z��0{��k�b�Y�n���6�
�g�y�k������!-z�L�A��1o�>����s
E^H/7�8?a�5��K½���+���OVN�[��rml�5��H�݇_:*��	��d:+�l��$u�Ԃ@Ȭۏ�z}f?7��%��S?���>�f�!O�&��Ҵ���G�]�B��U�m��d�w7�szs�zc�?^�e���예���p8��g�{۶�k=Δ�=�v5 �w�e�]43�N=-�\��(DR�Xj ht���Dۅ"��mkt��T��ݍb��޴Er'�)0�z��\+�F%z)�(�N�4>�������Ý*�w�(�2�5�4�[;vQ���tF���d�Fu��zt���~&����%�]��F�,�y��̶Q��Z��R��b�z���7B�,�&pF���G����������q�Y��W����]��n,E@��3�pMۖ���Y;�s�\�q��o�þ�o���-SLmjD%c7����s����?E5<����F]�����B��2Vvi�%�sO��>pgT��3��p�9ggL�邮��j��u����2 ���<�<I4y����	C�o=i.^��K���7��M�R��M8���E8_�74�S^+���c�o�2^e��2p،]E���M���0ܹYȖ�H���X��{7��**��Y7�{ә�����{�#�=���x{�`�O���<W}�k�VX�]7��8e_AP-7��*��$j�[#�i���������w!����^(�x���ۈ�.��X_�I
Cln�T|z�$l��U�L��=Y�XZ����?�k���;WX����ը��@�E)EU.�%QT7�|�H����Mi$BF�G�TSZ���`�d%`�e�g!�����b��
Ό�z�!֫J$�I*���U@I� *���UUE�P�
���1�A%�&0fL��QTAU2
(��˵�R�EZQiE�)�l��ZJ���M��Pd?�>��j��� סU*�D������B��P QT- $b�)��O�_�����?�[�<_�J�bl>�T��I��Zs%ౣa���B)�]L�r�#G��Rl�C��B�����f�f���;UAE�5�o��c�k�|�,�@�HH��&q"G7�U!J��];�S��$ڰ�?�?�HrE}1p������e��~.�/�T��q<�����!#C���G��_��iਥJX�i��j�⪨���m�U�J��?��;A�B��W��_/�d/L4�1U&�7�y��]T�(η�^���(�R��^����Y$�H����%F:�Yv4�{1�0@@��
�4=YN ��A �((�blii
&ʕd����k���M1�0G�c~���0�"Q�("5F��T�TD�2J(j�J��s�Cw"tkh�q3�M�F0��R��<��I���f��3'���~��lc�������-u��}�mw%%��D�^XTԼ9��172w#��o~�d���k�zg�ˍ��y=u�|��=ݯ&swy�Ul�9�O%#�;�Mh�8o��2z����N��%�y9��v�W�bQG����jj14.�?q,7y��b��"��4!"E��B"G�<��"�RV/�HꥥU��q��{{%��RjĦ�1bF�!쌛�BFI�8/J*���x�aޅR�p?T���*���TLV���r���F�;t��ۂ��,�I
J?� ��'*����U%�7���EU�A�^��gr�^�-L�(����a���	�.�D�b���I���Q���jH��,0tt�Oߋ�}���⓱7����)�b0$u�N�70����W��Q:�O��Q��L1x�R}2�x�>�޴�"Gc�sŗ':����Z��<��~�k���D�D��3x��.��}��q�o=��n��.ޏ}�Q�ƚ�P5t'������SeU����g����y�7T�R3MR5j��|���/���cԗk`�*�~y�)D��S�:��Eajm��������iљ�Pԣ�2�W���pc��UI���uZ4�d��Sa!��������ʢR$��	?�*��O1q�֍�,H�S�=>N���������'��yqI�bo3���&F8�Ȱ}R��K�]��r8�E>6-�W�(O����o\��w$S�	��| 