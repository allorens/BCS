BZh91AY&SY� ���_�py����߰����  a^         z       ���(�(UED�UBR�P� �
	T��<J(�IJ�%EB � �f��|
��}�=�k�rއ-�z�<k����v���z���[�Wg8 U㧦���"6ʡw���
-� �d!��J��K�
FX)[j6�OT��Z� �������5���VR5�v�ޓ�=�\���tu�wj��/y5��v�����՞�ۮ����ImE��w����U���NY���Sb��6� �,6���J^�Ľ�������ْ��������������T¨y(w^��F��#m�%vݚ]�R��{���v�I���  �	R��#�A׭s/w��;ǧ��{��\��2���[{��]EP�!�zgf�7w�q��r���7Ov���`���u�wWS��x� zUKcު׻W��u�n�]މy��m;k���=�F��9뷽��� x$7Q7k��x�
�b�ەu�Gv��%�.��u��Xo\�|M(    @J%%P (T�@,  ր   �~�jR��&�i��`  OЈ��(=F�2 i��FF&��*{E$
� � bi�  $�A	R�р4�!� `�dHhF��4��&�2�A4z&��iT�	�R�MA�C�0�D�n�P@�*��h� [�_ĺ����
�7Zb>�����(�	� EGx���C�	TQ?��z\QJ������Q|�`@�c�@I!�@nAQ�X�h~�.*��$�A>-�7�G1�&!�I$�I$�S�TT�q?:����g��ُl�����^�jQ��y��fe�8�p�� O!����0cpG�]t($d���F.,oa<�ផ�Fi�u�2�$��
M ci�Yԕ�����t�FMBq����i�8�p�dk!��_0`ǰG�b8�Lj�Id��Ʉ��	�b\s\E�(6�$i3�(��B�JIvDqT�X��}��z����%�5T*(��Bc�����zX�1\Bd��L�u�҅�. qЙ������W��Gȡ��L������Dc��i)b�Y�4i`�.v1�0pQ�0�����bR2I�"I������*	�� v���`��1����;e�bLu����L��B��-±�`V�V!�B���&@ǵJ�!3�,������2FaMQ	�|Ϙ�!2p�B�J�B��1�Bf�g�D8Hi@��"��2�0���4s���4c9�(�8p�ƛ.@���CT&1��wBe���8d��(�[���2c(c݄�hۅ����i���Ơ��$���w�iC���1�N4ӊ��)�(�8�LCţ��d3u�ÒC/S��Y>�ib�4d�4f�0ic��e���(8s�a]�Q�2D�L�#.Y�ǌ�QԢH����3R_?�C��=Lf�!��҂
�E3/Y�4�I'���w�Z��2%'�	�i[P�cW�B�r�c8���2�����cWjL%C�c"y&aD���p����q��!�c�b���	�琙�dd��0Ĭ�c(w��c&:q0��at�`���F$�@�K��8_1�Bc;���5��c��#)��\a����p��Ln�L� Lcʄ�9\a,K�;L��9�L���1�BcHgs!K�E�Lc4i3I8wФd�>_3(e$�0s��ɕ�������!2�Im|�3���SHcD&1���PC��z�c�Z1�
� ��ɐ1�
F1��0d�����g����I�LC8�\XÍEm2�*�D}� �H�")h��Gck$f=P�����H`�i�2��4g�C�ꑃ��� ��c0f>P���C�X�T|�����3�-$�,b1҆1�s�3���mFH�p�����CC5 J�2���O�2�,��c4c��ŕ?/�?���1���:P�1�c8�j cL'�1SQt&h�z��@�gI.P�:L��FE&1=P�kXkdX��##�Q�	����-$��t��g�F�Y#�Q���� c%ʆH�cj �&7J0f9�0X�Q�2]���3y��PƸ�
G�ʏz��ˆ`��}��d�u�я�����"!�A�6�
(��e��J�-���p�ҋ���e��w
"2"I-&YAC�&=�Lz�3�q\V��p���X�	�\D�$�"	��"�1È֙�gR��M0�QI��Ld�)A�	/��bL�7-q�d�D�.�Rd���5���n�3L݈x��D?�`��C d	�Gى���Ez��=������f{l�����3�Պ>`�C�1J���1�[���[qY
,�2���0f���4ñ&��G�S����C�Tac�qG���֣	�v�8�F�dK�1�S0撲�d9P�6�Z��(d�P�?�c�Q&�1�c��/�⏘�ڌ$e�(c֬cB����H�%�H�H�mDf�QM$���37���YIA����,c��	4c��e�j,�j(D��@�֭�F�^��騁�p��h�Q�Iï��;�Q.�%�1����ӹQ��Q�k�!����3�Pǩ�������/�gr��,���I0h�4c�|*,�Ln�(��,v��$d�!G�2�c撣SI1�ߘ�$c!���a��c4�Ցb=_0b8��2�$f�!���,���#�s �	#~Lb)8VH���@�|����H�K��qj�1�����:\.�����Uq��&aڵ҉4�dA���0fJf�C$�(g9�s�1�Q�fҲݑ��P��+� ;P����U�E�5R-%)�wv2^�e�C,�1�& �A�.
OT2�{ma�P�Q\�4�l�C(D:����(����Ĥ\%��i�q��re�u��(�U����D��ˈw�>cX����P.P"���D$�v���ǈL��Ꮧ7�ь�ۈ��b!�3�Ť)�'�2�Y�$�e��V2E_/�<Le6�	�c�Q���H��!�8R1�Q�����6SV��7�>feE�r��4��Q:Q�j��C9�$�����c1�,��Lf9P��3�r�n��K���ʄ	��j�1p�IΔh�r����� �j>�e!�!��C dcQ�S�2�[�ќڎ8e��\3Kڌ����@���!��fH�'jH+����W&a#��8L��(1�	�v��z&6��!Q���H�3n"�2R7�~0i&��y�+��X��a,K���ߜ(dC�,d�ɖ2��3F[�����YC��S4c��X1��lf�I��q#�K��T���YE�J�[4����EO�c-��(c(ߙŏ,q�|���2~��p�9�XS�H�-g�ȑ2K��e2E)��Cf[�ZI���(S���E8Pg�"��k6���. ���PJL/�r�F��KJ���I�S�p��{!&�P��S����n�aƬ�8!v�I�җ��T($�!��21mA��1���)+���U��B�!Ƃ�����w�$���[<�m�{��*�2��%ۯ�/���u������{ٓ۲̛������I����5�Foou���Չr�ȶT>��rz��6W3Tl�v̨Qwr����sw΍Y?- �}�٠�����qU��6o��&�3#���Z}�>�i����dYv�,�K�L�u~7ss�,Y77���5�x���v�u������F_�Û��&u%��nڏ��l�O�ӻr/q+�P��eF��Ŵ�ly]NzT\�:�}���:bg�:��&���wh�Ѫ�K���5?��־,�7���1�ۇ�҇s'��]<y{;5٩)�ne�^ګ/�(�w�B�OǴ��Y�����u�H�b�O(錩Yp�����ܵ�|~�'{�t��~�q3/n�p���3��t�9��S��h��5����$� �l�����M�XX�}��.Ja���M)�[�[��NI�;�돩_!���R�T�}+��\L_^ٛ���+����}�]�T�����컌��"g��������ǆu��������9D�K�SR(��>{&��!#_����H:CcO���9��
N�}���D�����tˮ:of�������e����H�w�����f_���o�Ok{�o=J��ef)qx�]������[}O6zk6�T˩��NGd�qwܶ
]���]���K�9�u�����nk�N�r~����O^���b����y�Y�v�J?��G�,g��A�[��C���E�eBԖ�j&�eNZ�"2��ws.������(��w���t�[\Z�ҁe2˸�͕�W�������47�⧣�enM̺3}�>�d��B�".Vϳw�s����Y�f2g��#nbٛ�����Wf�G��~q޼�YOf.������TT�%[=���C�"zcnsN�?~/�1V}����˯�:m���-�ܙ�����MK����j����L�;�zS3p;�BdO��;=�m���_R��"v�Fî�Q�eZ�ڢ�ט�{�+�����{��Bzos|w��ك�;������3|Dϡ�ϯ�}'��~��c��̏u��4�)�_b&/k�N)Ov�+/jz5XF��Q7��<�v}3li���3�n�,7��6::+���K�ͤ�m���2�����m�)l3%:xtC��{S<L�N����kW�X���/�U7w�.(�������t�g_N�&��;3]�7�kG�t�wg��Z����5�3�y�)�uv�����n�ʜ�"�雲z�]����j�v�l�wMNf����y*� �-t�Պ��
�⧕rJk��w�]qy�����#9K�^��E�����L篬���[K�;�Y�it�woJ�v�Y���F}J�����UN*Y}�%���n+������%DO[^ƻro1Dڮ\�Q�{wi,��땕���I'��SSQ�=��nK%Y�|B��9v7+�i��'�gx��VLRsni��Z��F�ȋm�K��_�O�{]�7�})��g{`=U�9k2�a0����D�Q�Y����<�gދ_~��ѧjƛv^���fljR�C,կr����7�ߕ��Mg�{�9;32\6��@̕��}�Ϟ������g�[R�A]�'��k�釙{�ٻ�/9�:*��o&SSLDOU�t�-�\����R�6�۷70�TE52L�NϽ}޾�2�����������3N�˝�5T��^�ogM���޻KZ��ޑ�MB���=9;*���oj��d���e��\�.�g}����O:�en�����S����lf,:�P�y��#��d͐gvg�����%W_=�r�z�vu�����q��d��{57r:�SGVob���}p���햯�����XZz����Z+f�r}�����n�_+��x�2��]T�\�^�l�es�﷣�F�a�=�ޝ�wݎ/�yM�fo�����=�FU�m���{5f#���w{.ś>立���\��o�U��S1�ՙѐ��nOoN�\������>�v/4̝�EӍ��"l��s9�¯6fdӰ���e�8�g�����n(��û3rE�C���og����2�<o�i���i��^�ۤ ���\2�wݝ�uդm�Z:m���}�A�c_}&��Å����<���'q�|�C����T�цU�Sq�ύ���Pu�ً~���e��O�Y�ӽ��|e�@��LM�z0�df=�Z�4�<��{={�Տ=�̧������a�����ۡ��0�zzv��Ր�{�i[�����qu�ܙ2��Gd7�껇I�1Bh�ǝyp#w��	:O��ű��zhۂ�_hi�{�d��u}���/_Z���ߺ����M��a�ź�����Æ��B&�Q�Qc���u^�{��vt�ע�U)e�W����m5�OF�,��/�ovC.��l�Y�B�1&���d0Y�,k#0ݪy��Fif�w��v{l�尮2U�T����̼�u7�<Z������ޝ��F��yd�{��}����NXv_<�����2&��{$�VW{C��I/G��֣7v ��~m�Kd;O�}dz)U�L���1}���Nᙿm�ܗ×Ұa��7^n僲nN�K�:�]0�>��!J�ٽ�g}$c��¦��N�w1B�˩����J^�{�]̮�j�Ut�Č��vF�e����=�F���w�"�]=�0�뛾����ґ���xx�G{�6�S����~��:��ˁ�����5��{d5`��N�c�{۞�������%>�L����L���ku��Ļ�����ckr��ב{��N���(J�u��ؽ����2�fr����������v��˫�N���"�&���n�f���aW�b�O6�G�=�d����7g�}wd�I�r}�{�}7�%��y_*ƺ��7Tg*��#�{&zf�s�{��6<Y�������Y���=]�N����f.���q=�霵����vo�)eɐ�n�������ی��Ko��:�mL�F�f����}3�̽��˸����`w9�v=���Ni��T�Q��ר��s���������.���]ۓ���E�}7#�>�K��ck��M���Ƨgj�{�Y�5�;��uz熩���,$�;s7�˾r(�����������o��}���B������Q�{�nu�Q*ɍ�f�,���m�w(���՗Ԡ�it>Q}O(���u�ݻ�ݘ�NMN?j��w��N�]�!���RZw����6��-ȫ����ܙF酽zrޛ轚��\��,v䞛%�I>��b\��d��*=0��!]ą��ݡ��Rd$x=00M�<�#�{y�oD��!	�z�F&5V#�}m�gx�ܺїi��ŅD�`Җ1nt�խ�Y5F;N4�Jc4��)��&�ْTؘ�4���ɡc95R��Ul��vX�W�s����V���\8u�b�8Kz�Z�׳������g�r�,��&ʘ� �qʭw�1��s�[�ozE���#�E��4��%,4���$=y
L���ŕ�g���5�{7V�ӵbP�ٵ�����0���Ktayn��mkq�>�d�Ք�(�%��$o�˝YJ����$Y�*�����Z�U�^gs�vdᄑ� ��A��6U-��RƬsy-�B:�*Ց�RIZ��"��K����e�Y]R��Q[+ ��9N[��Ԧ�N�����]�흸!�o�b�~E�U#����շ�d뢬���HBd��eu���gs2�5M�b6uI%{���c��c�X���[v"0�^r�N�W��HVH��_����;�e�*D�s�q�K�LX�tu[�36�5��u���\�I6�ΰd�˟��Ǝ|��}feV>B��-��ȣ"���*����]�������
�\\��J��[5j��b�Z�W4�� %�V���";P�,� �:�&Lqrq_��8�=2鍋�4�y�r3\�k9dT�K�!;~:�T�֨w	�\=M�=UΘ�;iY1ktl�!�|v�Wa�1`�Qư�^�S��G��[�4�)>,|$��b��.��gVCK!`|,lj��ras&;�X��jE�����X�D��~��-]_g��$�܋2����q��h4���-��B���)ڋ&%��A���3v�䰙�w5����Ԍ�͵]1mNCA�!HKlХo�޻���(�d�"���T�*Ơ=z��"���BF�#cjD��P��]33np_kBBw�>�Ք�3��3Ʒ��R�쏭AS6[��qO=�1���!##��(�L�g ��Ƚ';dÝ�KlK�yK9����M�cg7&4��+%f6�ŭ�$�[~��K��c��	e����Mnڭ�Y!��[�#�U\QnJ���8���1}ً5o
@ �!��!<_�ne��[���U�,"�C��^6���dw�\�g�g&a�^a��c_nQP޶�%�7<�xqO�3��+ܸR}�������Wm7"�
�S��<Z�ٴ����G�w�	��}� ޡ� �V��5�14��ݪ,ɢ?��8����'��,sm�����(�&��`��>�,r�Th�p���݇��y]���	 IB0M�ֻM����y�y��m�n[m�m�o[�m�m��m�cm��lm�����ݶ��z��m�nm�m��Ӧ�m��m����m�n[m�m�m��~G�||}�||��[�ۖ�o�m��m���m��6�����7-���r��˻or�n�m�nm��m��6�����m��1���Ѷ�xۖ��\"*�,� H�� ����$|���|۞���ݶ��z�m���6�m�i�۶ۦ�n�n�m�xff[m�M���ܶ�v�t�m��m6�v�t�r�m�m�m����m��r�}��( K���{՞��6��ܺm�x۶ۖ�oM��|��m�nm���m��fdfcm�m��4�m�m�m�m��m��6�۶ۦ�n�n�n[m�cn���G�BH "EdDB,��B���hi�x� �(���o������ ����p.7��c�8�FfC8f�`�`�F�2�I#$�H���@�$cc(����q� ��g3�"�(f�3�H�4d�ec��H d�1�c$c(c��$`�N���ӥ�ɖQ:�:�!�!�1�1�1�g1`����0e��Y#�Lg3�3�Q�8��h�ƌ4ќ3�4gac,C dь�FX�8c�0`����!�0n�[��N�ߪ��Oq����T��L��v�f�Z�RJ��Y���|�$��ȇ�;+���YV:��I��?eŏ>ʽ�ӥ������N���ˮ���%l��[2IXL��Q�2-m���k��acj�hj��betż��rMf>��r�To�O&��w���!�$БM�]�/6����ݠ���_�n�|�����Bjn�<���#��<�&ZN`��(Jp��Z�Jf�"�M�15�q�|�0�8�9ۚ�/VW�cLY�f}�ͺXD�^!I�o��{}�ȝ�@V�)�W����Z,F)i�Ƈ���ʪn���WOn�E7��(�A��J/(�%ή
~S�7�c�쵶H�EZ�m���R��� ���~�.�"YU���"�'�Q�s�{����F�`),de�nIe�0������)cD���T��I{�KQ��ӛD�LЦo��[�I)`�Wk�2_wHv�!Fޚ�8WF�H�z)����	ϫ���#;i�Wj{�©^7rc���f)�s�U��P(�P�JZ��曤�JGK46�d����H�t��חW�D�iv`���Վ� (䎲3��e��^�-�w����xk)iD�!�^s������}>>>��{����������>�=�{��{www��>>�����g�wwq�x�ꪥ���y��<��κ���m�R2N8��3J���%�FC��pJ�'�����d��uK��l�b�n]�UnIk�WIV��F�Ϟ�x�X��R�E�L�lW]���&J���e3�J$y�ޛMf�gp��.��$�ĒIȣF�+aZ�73��!��Hh>�0����d�����,��M��,���z5Q��uk�w��y$M�]9��;릵����;��<>��<�i=Qh�$Ԏ�[��Q�sƮ!�&�
����C������fQƃA�3�x��8�`�H�8���6͔���"eM7K:�ti�}R]��s�+&	,،�,=�U=��fh=8oa�3��u��h���v��R�;����C&%raQ!y4�Z�҅�Nð���s��;�&��^r��"!��s�˕U�G*̷iwLD"� ��(0��X�4�F3�0fd���,���(!��_&r���Vd��Q�_���u��i�w~�޺2q��rQ�;>�%��[ti4����\	с��a�.�^;��']R�9�j����⚆�ta4I�hw�J�1Xp��C�-2���q���淭�'�C�ȣ!�=�6xhgi�4c8�`�H�8���.-���Ҭ���h�4Bi	��ГBv	�<����P5��6��3V���)�ڌ����*B���V�.f�a��5 ΂?s��JX噊Q�g�۠�bl��G����V���zn�1���h�rù�-����Xl@�(g��ar�rNr��+iW���C��(��4f�Ƙ32FI�p�_/#�&��:�dj����"pqZ,����K��I��ݼ��4&�����x��I��R-v��eҒ1���d�E�֦��Pː��+&��i#+mNv���M �PQ��ʬ�`V��mTe�[VN�S��&�Z�%���Vi��=Ka�-�蘬�OF"D��n
?2$Y,�8a���߻��0��ه�e�*>�4a��ɱ�<�������|����ȦbE��e�$��8�N�9������}%6&
l���c���,ea��h�q�����8�N:۬V�ʈ�%�V��{�;Y��*̒��7����)�C�6����t蛛�A81��$�gIXZ����a�ZD�C�YfT���龍�v��פ�H��6�a%<���jC�Rx�*AE�"]����x�4�F3�0fd���,�3m&�p����g�JRa��m[D�l#U��5�C�P�m��"仱�:��F�ܱG9#]��^z�)��Mj����2��á�'�HnEE���k�C.-\C�yʌb�d�y�v�i��<\���>���L4Ï:�i�ic0c$d�qg��|�k@i�8�{�\�j����ǯQ�Y5f�Ǯ���������v��Uc�~u�eK��Nu"$�#����Ny��3�hs���� ���nN�>�;�)���"����GϘ�4mg��)�i[�k�(����4����2o�u�)�4�Ɣp�ƌgX��'b��j�|�Z޼O�D䓶\l��6��d�Rj�d\��*,W!,��h1�K/+�#V�F@�<�0�,.�Vڮ�l��[�D��S�5<By�G����ۛ[F��7l����p飉�����UVi�C�0��=;�R�:�p���YN��MÝ��dcK�!�A�2p2O���ӡ�Z�M�ʲ��a�6"e�k���F{��^�g��
zq�FjIxh�UR>����^y�p�4��1�2N8��`�ˋ$�
�T�}f����g����:x�k�Uϓ4�<���Z�Wr�]DB�x$!��ڤ$8�Y~��9�D��arM��i�l�vI����9� ɉ�8�R
2�ֲ��|xa녰�&NC�b-!��^���f1,&���;�|x�����|t����f���I�p����d��<B6�p��,���0Ӭbi�-<i~=s˷�cɴ��������[K�u��2�N�ίO/�����>y|y>_ͯͯ�/ɇ��+��_�|Ǔ�<ƓɅ�ǘK�-���Ǚ_�k�by~u�<�L�_��i��ז�e�ů))���y"z���yk��%��1'���K�y��<�'�^߮~e�O��O��?0��/O�m���<�<�L�<�����~G^_o:�����:�����u��_�c�uxqo8�'���lZy<���؞x� �Ƒ�a2</�N�Ix�����u�e�W�������@�g��X�a2����.w����"b)�! #n�Dkv�կ������m�zw]���f��s+�n��������X�����y���,�q���ĥ�����ȳ�n�ɼ�b�Y�!Ǎ�l�EmdqCc��Sjwl��N�5rN����f
o_5�о�{��ŏ�S�QDX��gI��s���m�����f�+ӟN5���� y�m�ߤ�|P�]Y�/��B���Tĭ�h�,=��"هꂿo꾥�4��JR���>�������ww�������{wwww��}��{���������ޏ{����ww}��}�,��^q��:��:�O2�2�.�ۯ>>/���>�ֲ涪�2l�I��a62z��d���G���P� ��	�����pL�`����ԩ�N�Y!�}ѥ: f�t`x�BM�"Q%@�0�+ �&��Q,��-	�8!|���[�Z�f��ƕ ��S 2C���R 0��9�)��
#	j�taΊI��6��?%�K��=IE��F��42C^��Ô�hC꾜���������<d�1�J�5���̛��N�D� �6�0�|�2���vS(v����y��_��u�\|�̼��ˎ6�ͼ����/rI%DB�}0X�0��d��P�s� �`�XC(����8"'�����K��QJ��hu��1�JGL��:��N���D}UW��*J.9�dx2C���HdO2��Q6`�&�C��Hx2M�	,A@�DG�E��L!p~�I���M	(�؞O���76%����k2���U#�J� � �d5�ګn�pM�!��$�1�B0�O�N�<��DO̡<dRGTUNp��9�M�VCB	�I�k�K'�!���e��GͿ<����8돖��<�(c0g�=�MZد�&+o�.ݣr�c�&U�6pC*��ݙ�u��d֙]s+a�l�p{�lpm�B�l����M���Z�B�w�_�E���r�R�����dm�Qf�%��t�����*��n
�B��� B�&��K��Icm�mJ#���9ms�g8���Ug����@�t@ў �����J��A`~��[pղ	<�tjNC҈���!:�a->�'NID@��@�d�'�ih�l�B;�>jI���B�hDN�!���@{d��-4!'��<sR}i��$�[TD}T@������,b`{��M0S�X��8~X�����d�~�M4"h�i4�Âd��.a�bؔH�R.��Ԕi�_�KR���%�Am��q��S�t�ѐ��nL�Y�y=0D��b�R��~�~f���]4��m�~q����<�O<�/2뭺�o;z�a&�Ub"�Dd}����D���P��D���D�dPr¦"&�0Od��Z��FJ�	�Ì���!�C�!���&@aD�2�M���Hh>,�I�c�
07 OP�D@��(��2b�B��2�"{���=��Y��%a$�[�N��ꈨ��NA�� w���E8�����:08���7��6a0�OFaDM��#"'LT�� �!�
[
"$��}�#Z3����2BJY�0Ğ�}YO�<���8��u�<��0�̺�n����Yb\wRI%DE?2�=�㓛�FC�����M�4"'�0��D��T����][	�# h���}�iL	��d�hND��톧D�'�Mz2Na�0I��!G�BƇ��X�h���t�b������m-�����|$��9�i'{������L��,;
��'�e����,7������C�7���j�7P�C>�FE&�*`�L$L��"$0��S�rt.X�za20颈�6���L����r�O�4��8���㍺��<��0�̺�n��Ϥ��?R�GV�� \�@>`i\A�J}UV"&FFQ?�'��y��F��v �
�(`h�?b<)XOt�g�9�C�ީ�,l���Z���vK��Vҙ�@�J�L�!y`�D!�!�=Ҧ���r��c]����s��l��A�0Cqc$���A7�dD=Υj��C��z2O�(���҇qd����$��2C�d��i٤��5$c1��I���=�hڣL��'D �'�c\��Y&�?	��@М���#$3IT�i��)�S�-q%�0��YCe�X���YD�'Fԟ0��CT�Iѕ������+F�y��y���u��(��J<P�`�R��TUU*��c��+똃 ejV��xnq��$�B�p��j,��`�cA�ex�*�ٙ��o�o3��|�ه�o�d�9�#�zݫ��Pr�(����cQ�cB����7��JEޛEKk��m�G��/N;���g�a�8��~]S�����1X�iHA!�"��T�$<�� IR�' ��� ���rbO���K�N[sP�S��yL�
0�Q�萬H
�d�2� ҇�	�!@��9�t֜ծ�m!�C�J���[(v�[�a�bJ�E�P0d�Ȫ���(���x {!��4�	:�2ɡ#$Кd��20>��a�q���4n�:)}�/
)�c���k��t��{N]����ɓp�8\��2Ɗ�*r֟W�^6�#x��S�Ǒ�E�&+(�TSչ#$oNUҭ�J<�θ��?8ۮ�[�2��2�.�ۯ99��3˿�UTH~<|�6����wr?Cӄ� ��Tr�>I�,9���Q'�r�ﭮ�H?�K"��6#JA8fv ː�*d?�4&���77� Iܣ�������DCsk��V{��֣�
]�Z��N^�)�<����=������K*5M��}8���7Y�¼E>���i,�#vfS-q��j�Y*����~i�'X�0[��F��m���~q�[uo�0��2�.�ۯ6�=�r��ZvI$�r�>F"��9Ѹ~M���~�}O֒���+}\E�u��]��ܓ,""FZ�!� ��1���l2�"��AM)�KL$GEg�f#j�~Z���iX�DC��9�3f_��8Y�xr�y�3�ܸѹ,���b`�0��)��=���7E#"E�~��0{�4�R����2��f'�SY9Hm�W��V��{�A�!�uqnT���òTKV����?RA�[�_�>~u�iӯ<��a��u��y���y2C;]�Sp�J��4�ˮe\�}ip��j��A��Ja��XT0�3�����Z7!�f+m2��*$�4�kk}Q�FQ^��ϳ�\<�!�m�)���[W1)�]ɘ�j�.f�ܝ�)�3��d.�Z�?U�����8�oi�N[�"�y�2��"n�?�d4Y<���2��������-Z��V��k�����-l�')�GF��a�J���	+��Ue��=�~�nA��E)�R4���g�RW�BI%VgϪ�u�?~8d��zU�L�^.4��\O�ɴ�L�^S��Wl.�Ɨ�����ci�痴�y�	��&i,^�Ő1x�/~e�<�~q~qm�ͯͮ�_����^�_�[�<ǜ^S̯\�/���-�����y��>O'�y�'���y~Z����֞=reh�Hn��*?
?/է�|h����0�&_��y�L<Ǔ�\�ly��x���?/��_�W���?4�g�?8ƞ_�_^_�/�ח�{��6���^=�q����ĳ�2H�и�6��i���y�e�|�y~q~e�S���S���z_2�_��Y�O��i��6����#�G����?4�d�����!������i�_`�d�x��R!nEIa��J�����TP�m��/�w�����k�P)�L�KX,G���n}ډ.��w�T������ly��ș�?����:�M�(7�k��Γz�s�#��+U�s�1��6�u�trb��M�r��VU>��ډ�����1M>���㵫�b��A
�:�nn�kf�T�9�)kʳ%VE%���8��vd�����$ȧ�実BSǣ�gmp�����gy؜U�D6���B*ew��^�e�W����T�+�x��U���٣{�����M�};]ou{.��Rv�Y�3��wY�k\]�-�Ә��dР�H���.(F�j�G���54�wnkZ�A�˭g WnC�p�2���F:b��/n��~9u�]_m���q���޶���+���T��99t��y��>3��zG.U\�S�nc9u�8?��O���2�`�2�&��2�$�����2�ݥ#R1D�3�.�*��c�kU8��շ��՝5^B�h���!��d�ƷmH�t��/�!d�W�M�Z�p&֛M{5����4Yk����ӻC�� �i#����l��A�8�6�-��i+�u�:cճ�Ĵ��n����{e�{1k��,i%���nP����[o#�!ZE%�AJ�Sw��*)��7�P�P�R�A0�~1���~}�ۻ���������}��o}�������mﻻ���>��0f�c8����$�ef���U
Tۆ��U����;׺�E�je�%UڀrFee��Q�h��H5ڸJB�B�i��|���YK	e�MY��Tu�y�ț,.��e%SU���콘�,h-V�	؛r�ݲ�B��;�45 �Ŭ�����[Glcm�r���/	�x|O�֏�w)�f��-Ƙ%5�l?�Obl3$�x�O��p�ш���'�{[�=�(S�����(SM��ᰚBC���=4h�@���{�{�������>i���0�p�˒����W�NS�NX��=?+d�O��X�#5�����y��u�^~q����<I����J�Bʙ��w���*��r��)���<?JK7�;=*��Q>)�òvj�d��~Z�ߩ�����Q�=g�������l�5����i�r���Q�v��*̸�V澔����2t���?uكd��[%f�i� ��8�Wnb
�9>��A�(nB��*�����0t��hS	��
`��!���^6��Xj~���ꮢI9T���>y�_�q��:���y��e�[u�����I��EIA��a�ѡ�UD?�?�hÌ�U���?;M�o�3�3Z����ˍ�T�̖��-󙋗0�y�sT�a���''f� �O|��S뚙��u�b8\޴ࢮ�La�g�@�l�<?Cl���TW�cR�h.�!�v�!���)�/���=QQL�֗���6S��Ɔ�褎��N>�K?4���_�y��t���y�i�]mן>^�u=�UD��>����Λ=TΌ.����d|Q���ϡrSW�k��q��uX�-�6�]:3p�aHI�i4tׁ���C��iY�;��)�Ǔ�9�:x���y��8{4d��0����0�df����k���4h��p	����Q[s3(���%G�g�=\n�y�I"2ɿ����?RS�;ïI�2�ԏ�f�6�������6ӧ^yg�x��3xѫ[)&h���U(�ciO��텔�v��v���Q�ˆ`�Y�:�N5��0�5���Ћ֏�rIKg��*�9eΜ����dB�nѤ�����jr�v��L�D  BZ��5�%�v�'lp�Z�(��
���7�a�h��ِ�W�/��]a�G��b�������C�����}C�!��0?C�g����4i]cuw�v=��)�M�¦������y�o�R�l�CՏ�CZLWs�~]0���4���������Ytب��d�>��->��Id�UIO���>�0�����D	�!�����,c����e�u��y��.1+qRn(�\⪢�����M���T�r>�����c|l��sa�ںk��$[,�f�G=&�+E�u�Z�}MS��lյl�Q�l����V��km0m�)y>U+d�t`���>�|0�y�jK��ǘ�*�qjZ-�mUO��#C��S�P�J���<�����0<2n���;�|��/��m�$�MW��>u��~y���t�-�y�]uj�~]�ͨi�e�M�� J�+��ۦ-�߹�~�qr�p�i���������2�%:���G�w�n��f��1�nz��[�7M)��2����������L�k�I4�1q>>OS��4g�`�_I����N>FVJglST�Ѻ~��ϓK.���U�y���n�մq)�3�N4��xnŴ��
&C����J�`��ߝq矜m�N���y��(c0g�6�!�)��FL/�j��{��!Ϣ��'|��&K�a�^�z�T�b�ܲ��ffffi0QD0�Ð����ô����y���XO��-��9�f���
��鏤�>����g����^	�xk����=4j[V���t����(3W�|�?<�s2��Dm������ ��@e2ɼW�4��8����6ӧ]G�x��1�3Ɲ���S�
��ɕw)�*M��1�Lv���
AޛM�c�X���:��c�P[$O�[�V�k"c�ˀ`��C��X��"G�0X��31�@w�I�  ���!���ex���f8�Je�Z*�#�O	����CxC��!A�C��'x)ǵ��2&x���0y��ۤ�Fit��U�^�Y[�F�~��4�ȉ��Ca4���8�M�ޏ-��'�����Mn�Qw�$��D�l>�~��s9Ι���p������4�]�N7>��4E�x���41U����8����Q�e�Y��Dy�=�2�QQ�D
�(D�I�74ҥv�dޫ�UU�?;�l��3����l�/h�Z&�F"S�܇�!�,0��i�~J�f��J�ֳ2���;�<b$O8�7$�0��E�� �&��I˶+�iY$��K$�ۧi��qt˜^�w{`�S���m�̞~巰ٳ��0��D8L?-�� O�b�g��K�����?�dxL�3ıxdp�Va�P���<��yyN0�0�����o1��fLm<��y���qn<�z�W��a<�u|�]����������~q<����yq۞//\���<Ǔ�<�ϗ��+�̱i�y����Ǚ�obi~O'�_��=�SǗ���\z�yu�jM.4�M�/�[�\��_V�����<�z�������y����x�<���~L��n~i�������_��<���؛{��q8��"��y}y|�K󫯘y�<��|y>����z�G������Xx�zV�N����Q���<�<�FR�i�yo�/�#�O�O���?�	����}��$�n�����㋧$~�N�]�����뛪*�Y=�OLA��^�1�F����ࠟ1���"���P� 	_Tt��Mů�B��c�w���l1ZWi4�:̹�ަ����mƩͩ�-#�As�W�����OcVS"2+k������������www�}��mﻻ���<�m��www{Ǜm���s��=�CO<��y�iӮ��<Q�J��F��L%�W
f�Q^�$�!m��6a�o\K]#Wl1�p����'��C_/O�z�0�C�p�6�������A�s|Qrq�FI�كD�d��߳��q���Z,�zp�
=�R��f��y�۴���鱟C���cl�ψ�r�?{W.��қ��Y+OS8��,4�����t��Ǌ<IG�`�Ou��>�I$��=�Q�;߻�$�{|2��4j&�Y�|��K����emr�d����p�g�:{r~���g cO��孇)��:����'+h�)���7��%LY�2���P�,���C�ӌ�Ja�׆NM@ԟ}5]?-�~x�5�˩)�i��;K;��
��[�6����?>~m�N��<Q�J<3x�W�I�H�!ڋ٫���Q�H̹*��xA�BH�G��J0v�������e�sb8�H�����.&˙�MF�,P@����9H�E9`��8��|x퓊#�� �V���lY��NM��[-1��rF�D(":��U��YZ��~ 	9�M-v�8���%�d�%����Jh��<>�h
z>�NR�[_����ŭ�?+�l�Y�,�1
zf��y�a>�aJ�ks,.�n�;]�M+4���k2H��V֟�WI4�2�SO��{��i�͇b{|�?8"�?����m�Y����S�6���M��=>E�O;ӝr�&0�NS�Y�qן<���t���2���n��fv�x���V�3j��=>�Kko���8o��[��p����!�i`�Zە�p��Á�MA�b��bi�mt��K|��m�]���R�qc��s��"�h�$њ�b:��P��vp��M�l(YX����~�iȑ�7��I�Su��C��2�7��VZ-<=��_߅>����8�κ����t���2���n���b籅�rI$�r��L��l�L�y��6��q�NU�N,����k]�N����dDC�h�*k�!b�*�Z��g�C���$�Eh��q���Eg7.��#��'�׫�B�~ÿ�x���]:Ȼ��F��.�L�W��o�K�9OJ~�u�Y�_�˩ۖ�v�[�N�ە���d���f��^�NS�ԓ��C��~�H���ϟ<�<�N�uy�^a��l���vB=��)����p�:�j>i�/b~�~.�*VQ���h�R�%�鄐SEi�z�����}���a!�Bj�Y�5��e�_l��ߠ��p��2���:l�7�ن��
y��՚|M����&/Z?z����?U[���ێS-+&*�D����ta�i����?8���b��G�<X��N�Z$J#O�;���m��bx,��:�+O{2�����0�u�E8q�G�weӚ����c�+n�6+n�C�����sY!Zkd%���l�AR�mt&�Ix��ei�����`��֣����I�)��I$���ZJĖr�XBrl�1�\0ժ�`l��rtL:oG���7���(�掘hO�w��P���=�qwU�}K�#�rgPY�pNC��E������*f�0��6]!k}U��?l�y'�b�#����@�t�8�+UM��)',����ez��$e��cYSxNS�?�	�)�^�.K�>��#(�ߜq���,`�!�<Q�3x�r�B�<�M�B�˙���
e���7��I$Bq�Sբ�Y���%��|�0돩���j�e���h�i��S�Y�}���4!�Xh�S�2��O��J�͛��0<�C��Ȅ�.��&���,�Ȋv^2�]�Y%'#'����Ξ�$��dR�&ϏMn�S��jf7������a�r�3Y��y���6}I�Yw)���rW���~q��~~q��t�g�x�Ō��4�^�GLR��F�ꪢ����>����ޚ=���\�3%�ì�bȲ~5�C�}����l|��0g;��x}<���v`~ϔ�a�2�V�c�X��)�S��h�s����a�OHɹ����g�0=цE|��٣$��v"�t�Z�Ð��n~��2��n��,����E��1K[+�S�?�X����μ���N�ue�^i��y�q������0	V�j�.��}I$����+/S�t�9�gi��V�h�2}���C���a2K
�F]Z�Z��\)Y��zc��*~C�6d	&K�i��M)�Mѡ�!�"��[n��iX0��t�^�	i�c�&��e[6��d���E�5Q~���G��]=H�T���"����=~[L�	á�@�����q�5i�l�b��n��<�3���3�{�2|t$�ᑢ�a��F�xXG�^^E���Kyp�<���I�c̯O\��y�����t�I:�N'��_[[ΰǝ_��y|i~|��_�^�)���Xx�y~O<��<�<�6���)��������痗��[y�'��y~NI���.<���04���S�X��w�e�|)�|����������y�^�_������̮�\z�yq������w�?4���߱0����c�\�yzy^:��p�(K���g�䨏�S��O9s�1<�'��6�O���e�<�y�N<�\_����|����S���>)~:]	L.ƟO�K��H��~8�ֿ��b��K���Mf�m6+�R�s��sT�ɫ�L��������x������i6;�U$��̎���d���W*u�� �Y@Y[�"�g���7�+��l��G��R-��k�=_�����ԫ��s3��x�]�����l�oE�X8rws�w�۬�SC���]!�+�E�r����T��s���<�YM�:���Muo���vUS��%$]��ʣd���Zs���D,�����X��f4�2�Ĩ\Sl�R	�g��V2�X�IIm�\:��h�K&7��7$ݓF��h�xfb���Vj괲D�ղ�͒2&�lhۖl�F������E�M�h9*�&�Ҫ�[I��uy����a�v���qZ��θ��e��D���[������-��I����L���Վ���5���$"5�.2����6�9�u��Y��mZ\ܛLi�7re���j��$�%Z��LmR��2N
8�����a�T��h22HT�A�[(�-.HKY$m���3�����0�b���A����������߽���o��������m��www{�^m��}����}B<x��1�31�g�x�Ō��4�ԉj�*�)�D�D���kE�$eq��)��+������J^ѱ�#�Te��<�\�&�3
�r��'A�n��tn�ʦK�Lm�Y������*��� ��51�U��^J�k)j[��f�2�Q$�H����7fN�]w)-t���ٌcV�-�[����3��4s��H�&1Q�]6�-���[C*��h��r����l��rrsk�d��9�3��|��"�W�s�]K][M���]τ��-(k���̫�30ƚ̘T��~����C�5�����y�]��+޼LLv�m�<�m??:�ʹ��Qמe�^i��y�k�����Kn����{=&C!���YD�N�8k�Ky��OQnI4j�Oݧk�\�S��;L��~f��I�)�Ϩ�JWG���a��OXI���7�9�R�R]U��(� �9����]�V�����T�h��CSg:S���{
^d�挾.ST��߹"�`�[����c�|����aſ#�4���~m�N���<�̼�m��s�za�h5����{�sG��ԙ;�ND��g������ӆ�o��3Z�|�hl�,���f��9{��"�Ҋ�Nd�)hD��1�>j�S�j��n$r0o��U��<̒6`��q�s���%���z�W_Z�u���SJ�)���]�T�I-��H���j���i�Vۮ??8㭴��Q��y��m�^'���3_a�⪢�<щAZ�e�Oj{�~�d��i�z��k���S)$E�h�WZ(�cĒ�i�����Hy��<h�?/D{*���G����l�%2~?���4�)$�״˜�%�E��R����^#��W����{xg	Yo��CU�?��=�*[{76�N��Sݭ['�Ub7K[-��u�y��1g�<Q�`�}ޅj�ꉧ#	4���i�f���I�(�%P����Ec�0���|eE9k��֛���Jw�k��5h5r�@ BS &�`&V鴘Z�]�a]f�%n�,&�EUcZ�jxt�O8?{�E�Êv���4���]ĒT_#�m��OS�ڛe�N�g���������;��kI��L�oK�1�W�Ja�D�?St�#t��et�W��j�C�u��}Xa�̏�aJ�.	���ۤƅ�d��¢�)����wT�4��*�ER((�X���R��B��R[��:t��~u�jG>~eo<���<�Nuu�^e�[8z|y>ej߲�e8����Jn��6&�'aM��$���wE����̕�J�tԦ_���~F��[��p�ZLֱ�t=�JN迿���Z]0��RY���a���̓'���l�G'�xl�?�]�[[A=�]��F�E	��1�Ȫ��!���:l6�>Y��c�%l��M��=�����ݏr�.�1N�`�~��/�T���4��YG ��<�ʹ��Q�^e�^u��x�^Zi� ���4xa��}eZ&�x�ٽ�V]����n�|(�B�7������˓��(~�l���粛�({�ׇ�1�Ԯl��.���B9��F1�	 qUj�7�"�} �Չo��F�5}L�1R�����_2�D;}__\ˉ���;
j%�����L�ڈ���^~�����
4�8�Y��!��G�<2�=>=Y>Del⪢?}2�gT����-�Ch��ig��Obmw���'u�#$���#��9�~��d�!o�a��~�a
��ψ�9�ާ��#tZ�L�L;Ç�R��܅>ՙ��:�-�8 ��à�4̟����F1�Q����0C��)�t�U�~��~|���8�m8u�uיy��b�����L��������jF��,��2U�̯��c�AkX�T�q%�Ƣ�b�q���Xd��N.��6VH�óno3tź��Ѭs�h�<��Y���*�q�� 	J��в���u`�Z�W#���]�$1	{�������H�mo��޾1x�bN7�q�S�]>kIt���Ѿ��S�EQD>0�?h�;
��~uV�p���	�r)�l�T��A*��6!�a��p������s��K�a�M[P��.	�a�4qo,�51ЇC�0�d>���+R����짇H,��q�8�1�x�G�`��z��C#�Hi!���3OY�фC��Ջ*oVGU~�UT7Ks����u����E��뻷���ͱ,�g��V�s�K��L�����lZ��w:�e�-X7V��ه������e�co� ����3�wl���a����Zt�0ѓAq*j���L��)�Y0��#O�76n�9�sÇ�ӆ� ��vנ���;m1�}�_2��8��~q�{'�y�^u�4�y�F`����2�C8��ќ�1�3��4f�3�,�Fp�!�c0c�Y$��1�1���C�Q��֑գ�N�a�V��:�:��q C�1���c`���^y��y��y��y���FH���шќp�4g1�3��0�
1�d�2ؙ�;D�iƖ3P1�d@�P��p� e�2��DӮJ���tyW�n�����jww�3���/��K��ܹ���N�LP�gӠ�+�n�<�2�7sf'V��1	WrE��AZ�웣&�	|��'onZ�R�J���}	u��c�;�x��K`��DN6Q�托�Z~7=����W5l��\u�gwn�������m���ww{��y��v�����z<�o�}�������4��8�Y��!��Ǌ<3a��S�;�ep�⪢=2n5#�I�����k��E�O�e�h��JWs�!���a�i4`���C��4�P��mk$��@x��m�f���`/���D�W���on�gL[�ӌ5Y�W��h��'n�\��T�i�_B���C�ZLGʺ��
Y �(n���_�|��?6Ӈ]G]a�y��p��w*[@�OZ\י�UU�m�ji�~�zT�V�|�0��`�[�7���ա%�n�ƤZ�i��b�u.�}\���>���̻M�"#壬�`�]y�i�.�[��˻��j��gԶ�R����N�_���130��7a2	D�����Y�_��r�)�f)F[�8��8�m8u�u�y��m���/ߟ�M�P��˘�s�b�-'V��Ew����c#d�H��P0�Q�q�Hj�L�G���UV�L�L�E]2:HL��t� K�>:��P�KJ�	t���%u��mH]�����S�����u�9Kb�=��Q�U�S���(v0��jnAa#%2	�g��[Kd�
r�7W^vL��4�2�E�~�����=^í8��n0}��p��G�]ܖ��i�9�$�L��է�����]�^P�!�����jh���f9��R|(�� ��;���ܕ6�GXe������:�6���2Fx��0e�<u��]��)�a���!�:}ǇrHf�%�p�)�|�R��H�'X'�Xu�>���� ��{�fN�S�$m�a���2ᅧ�K��|^$}'�#�!��Cs]�f���A9�EO���"}!�<!A6��h��Nۉ\��8$��6��~ձ�a�)�mw��b~m��[�>y�~m�;'Q�Xu���N�>=��}lLhAq1�I.�U���p����&h>ק��{�˽��[Y�S��UYj�}H�Y�5?���g�_Q�&�t�q֭nkS5.e�F	E't��MOD�<T�k_�Oޜ;�Z��(��.�4�U)�`�^�5[�ǝ���4��D��~�ٙf[��z��������_M��+^�����8��a�q��8c�H��Λ>05�|��gnd⪢�<��]���g(�F�*M3^��Oҝm9����GJ��%��(�U�1S�p�O�5��"&�p��p�P�6e���<;'�����O�6�5Y�FHFY'\�>�͟TJ�I&�)�NA>���~����;��N��a.V`t�S�?0�~����?Cgg���Y)��f�Z�F[[����8�ac���f�{�؈q30���~��.7��:�o�%��G!���o$/Z��y�ŝ��T�o6FD�ɉ�D�IQx�6�\��,���γ7[0�i�y��KF�yI7-kq(�F�eTVf� ����| �0ب�`���ג��qЬ-��ZI�+r��6�a�φ
��؇;����5���|H�߰���k|�I��^������?7.rp�p݊P4�G�aMʑv�a�)��T�m�43����!Â}:�Caa�t�'Y般MS��ɇ���{��kR�Z�nڼu�	HO~�����y��T��R�L8~����T��۫0�`��3�@�H�xc4��d��[�$��E�� ����=�(g�V�A�וn���aK����aO�t����ˊڿ�������R��4��w+xd:�ᐰB�8������*Sne*����:�[J�,�w�����d���V���ݩ��dҽ�����K�^���hD�h��?'�x�ac8dd��G�3V/��D�	c��uc[Sa� �C�����b�7�R�~5�Aw��������]e��t�?uf��8e���3M��ZfZw�ax�j�Z2-{p#k�+��P�G���z�ȹXm8Ì�b�P�^h���A;�4����Fz��U�{-�[����������Zֵ��hy��짰g��/���������:�N���u�_�y�_4�3Қ��9��!M#PĒ�AUEV2Jʙ�UD<�=Ed�2�U�jO�����k��=(f:>�
F�Wus1Ǔ�F�y5���?9��`�I���yy�ٸd�PL��}94\?8Y�e!G�)�T��'A6'fn~��6";���}�~�WL��_?2G䣮�l6�d���8�G�3��Y�#ͼ�0��G�Z:�8묰e�3Fp3��qf����2�`�0Ɩ�H��c��2�$0`�!���e�c g�0`����$$�� �`�!�!�!�2�c��2�!�g�x����4f���4њ3FI�F��q�8њE(`�1�p�4f���3L8��"A�C �@��!�p��d���jR�QY>�.X�	T�l����B�>�"1ʹ��,��llx��h�2�e_f\��{�rq�6���?H��6�ϺvcSb�;���_L[������B\�q@�&#>x(l��z\1���Wj��Yk���X���^�V�ǄF{n�Y����owJY+)����z���k�H� Ώ	pˍ��f<� Lr�a�Z*�Yl�=�x���2K$ڮf�G^ǖٍ���Z����1��ɱ��#��с�I!"�7h���0��V�����IZ�;���h�A�n6�F �J�:N��b���,��ӑC�P`��u(�6k{��:5v)�2@U�E����U6V��qIr��~�����2H2a��f*HO������œnnj��oQ�l�^���.3'oL̾~����%�1��ª�xr��GI���&�ٔ���h|랍赺R���b[L�LP�##�5غ.��W�������#2��U�i�t&����N]��5E#����s+�[�GGYG�d��T�X)�+AH�J�����K+c�FJZ���q*�	FF���e�p�$M���峎.ĕκ����K�f����R����v��V��o-QT��f
O��}�{���w{��y��v�����{��o�������z|�}ݾ����x�ǉ8��q�� c$g�<1�Y��]~�_))L�T�Ld�Ś�\#2K+5��i&-K�k���\Q�fql�t�Y����FȒLQ��35�\ٮ�]^]�5Ə-Jm.k��M�&eM
���k���$e����� 	9yX(bP'-j��Y��a��m]	�蚇a��xxc%�U�x�'ZDd��'����Q�F��L�?b�'f���F鶜��"&X|~�ŵ�-���D�XY﫚���p������v+m/��xn�=�T�1~՟����LА��4��h2���s�
	D����LW<�~�����O��8�3�@�$����ό>��d�G�b�*�͈KKQVKZ�a�����S�UDv��h��}�L�����s�2d:y
BB��{�h����k�csY���|	`�?L>��h�b��H��5���6�-����')g��=���i����L�EJ�,�� GW����b�8r{����K�3LR����5m�E���׷h�q+�W�=:Ӛ�oq��ς���y��Q<2Fi�8�8d�N<P�<ig�j�l�2�dyT�q��H���R/S���!��;^~mh��b�+�F��kj��k2�Д����ǝ$���lY����
ԇMu��u��.�\�!�[���~6X~A�v�u$(�x�^n�m.�OԺm��t��n[D^��ye�G�BvDWڮ`m��g�K0Z�RS	t��[q�x���0gd�IǋǍ,����o�332냕�U�)��=u�����?C���Du�)0?_�����bSfT�F-��I���'��{�r���}N0�Kԙd�漊y�H��8��҇��r}���Y%#t��a��8�WU�O)ϛ����r�ul价粉�u�E{�y�)�z�����EX�8���ǎ8�8c$�N(�ח����tO"dvYOf*#?I4خ��N9K)Օfp&&ZQE�Ms-����� �vr�R��s��L9�M:��%����z�`TI'�j�n*�*�N,�� J�wM���4"(j�X舋��:5���^���,9�Q4!����ǅ�0�'��O	�K
fCO�O���Uٱ�BO5������)���ϕ8'��a�F��O�쒲���2��߽�|���z����v���m%��I��Wj�:!��}'���jM��������?Sߤ�u��i�Fq�g��'qG�q�O˾���ު�Dg㥙>�����pDMO��6�?C�?~^a舚�<��ǈ����)�OM�C:��yܺ�0�r�^�O�-�~�2#�����U�R�+l���0�W-���a����Xx`�t2C�/�6fZ�8"'��C!���4M�Ӯ��-�|댼㮸�8c$�N(��<iＤ$S:,�����g�X�pw8���?C�h�;>�����]�2捞̆��':���E<��t�M�Ҏ?]cu\���f�j-�����!�y����M���d,��=�����˾l}�Fi�aN;���~}U��]�:�����Dq_��}1��.O���H�A��8�O��xќ1�q'>=<>:|s����Q���
~�$����|�aD�}ഘt�������bA��,���{k[zcnl^�����	i�h�oǹå��|#ʴj���d���|��w�Y�m�_���=_�n�mh�Wꅹ�˽�g�	�~�h�W:��i�Sbj!t>n)��j�/i}�a��|��+��!��i1Y�[O6�O�y�4gd�I�x�ƞ/���^���_(��9��<C��LS3'���l��U�
5	e�u���dM�Z���w�<�.�;a�x�u�c�Z�92q�Ym *�2��#Pj�0��+r7hP�u�+"5>I$���Ԫ���5B���G�X��\C��D� ���M��pЉa����M�ߧ��HC|(��m�����:OǇ�>�a�8gƎzk��5�i�yU1^D�qf�O�w�F�Fi����E��.�ârE�`p�,0M��N{u��#]5ֳ�-�2��z���臾s����W嵆�n��[n�#L�:��f�c8�h��8��8�Ǎ<N��˚-�nk!�J�]k�UV"�V항�%�O8ηLR-�0����&Ɇ���Jh�(�i���U��]}Kq?u�iF7"�P��Ea��YQl%h�%�]K�$i��OSl�����M�I;�SF��Q;N̯w�s�U[|3U��u�V�8g�f�kK	,f@�$��ϙeo<�<�8�H�.�m�M��c8���!�3f�B�(�p�q�RL�H0c�Kc�iC1:u�:�t��0���ӣ��� �1�f�cDt���2�/8��6�ϝlc ь��3M�4f�1���i�8њaaE�&1�`�ƌ��3L8fA �!�Y @��22K$d�����s��2�&��[��j�ɛ1�e�J����G��=�	Ϊ�5J"���MZލqU��V�,��s]�^�e��P�T���*`�����ۜ��'6�2λȎI�{�����3ۖ�d��;�|���;������wJ�JT�ꎭ^�q��39"����<vd�o��}���{ޟ6�wo����{������ww��{��}������0�ǎ,���ƌጓ�8��x�ÔW�*�D�)ɕ~4\�x�Ӥ|�[5֫�Y�}�;��b?6���%a0�O�aa��������=ttX�i���SK8�e�(Ţz�8mS��Љ�q2�䵫���(����G�3��/�O\�&�}�ko���<���~��b�.�e�z��ۮ}&�9V����2�8c8�h��8��8�Ǎ>3f2(k��{LHL��Y4���B8��UV"g������u_#U6z$�+O������^[�e����V1��)Y>�rV�gB����)ޫ�X&��O�B۠�"~�Xw�?U���NCa��X~��K�;���fi�ӢT��.����LP���44�,)�}\e��|�2ˮ�i��q��1�q'q�x���S���I�T��gt*92�e��-+�NZ*����%LV[��<���t��IU,lu�Q����cnDͻ��`�S$ηer��u�� pB{�7��P+Ȯydh�k-������$�n��]qL6��ձ��YJJ�b�}ڗu[6�|��b��;��h��#�m"H�t��͙G)�e0ؔ6wn���xU*\�b�O`����]�qg	�~�3�k�܎[R��BI8w�<���F(D����D�YfxcǍκÌ8ˏ8����J��UU#�ݎ�7s#���=��܆���O�*(w�6R�8MC��nz����_��_�)m�i�i�ySFV��;��޶�=?j���v0�M�؛��򠊪����VR��޺�NkN��:t�C	�Ȋ��nM�M	�<6{�p�0�k�m?i�b��됿�rMUv�}�-��<Y���ƌጓ�8��x�þ��L̦x��G�ٝ<�V�̶�h�Ξ��6<O��!4�}�U�!�b1=�~5�<<T���R������K��hDa�٫�BT�E��q�r�	Hh��7\��[k�#�δ�D�g~�j�#�R-�FQj�n$�Z��4u�m�pF&�%b�o��l���K8g�q�Fp�H�8��xў!�q�˜UX��d��DGOnO�`�O��}�!�{�o��f�;	vq����n	ӾI'����s8N��`�ix�V�t������pMXCl;���o5�]k�ܭU��On���u���%�R:���ǐ�{7'��M�Ap��͈`�R��Ţ�a�~i���\y��'q��R�QDB�j��
�D�	��:Ȣ�W1>G�(*؀� %�T0Dh��eD�"Q�B�+�l��jfM-�p! =�2���X��$��K�LE���)$�0���UV"k9tב�4]a]�TX�nd�m\��>�8s�|��e2�4�����w�0��B�pn��FJQ3$�D���ޏMᲫ�r"X}��v(�D����T�!�Q94'9�����b`&A8'�_{떙�Y�������U�iT<��{z���kD#]��>�&2���yǛe��4��:�ϝq�Xu�q�|�W�,�_e:��J�>�v,�N�L�IQH,	���Q��Xm)�ԖDwQ�a��S�:XR��Ò�D�~J�g�tI�G��r	�5��н����Z&;�S5�m�mF�V��'�>IN&��徭�[�z\?CG�h���/�[��>��֧�?zrz~4a������ƌ጑�qGx��h��[3>L�kWE���UV"nSѲ{0ѡ7<�hK+�OyST2�Õ�[�|�Fj�H�;�D���ai�S1�b�\��ͮ�i��,��7GՃlֻ3~\.Q�l(�:�p;2Hl�=&�	��=F�ҟ���a��:���k�i��\i����4ӭ���g��8�4c$d�Qƞ<i�<�Am�_�h�0����:��I9<�D�g>,09
$~�}2%�d�ز��]n�y�{�ci�ɽ�L<�t�V*��׵��b���ٯ�Y�x�:�/���<�Q0�g!���ṣ��i~m���4�L4��IQx̸�q�-bO���WV��n�뎣�<p���3	0e@�$���$��1��aG��K<x��c8�����X�gH����3K	�D0`�!�ec0c����t����Ӭa[ ��B3D22A�c�ΰ��:˫uיy���<�o<�g4���h��4cđ�8gh�4��XAC�1�X��3�,cBb0�c�(������1�Y#(�|���s�ET�R�jyzB�T�ϟ�2��FMp�,�Kb�n�{f��fRe��=sX�Ν�	�Bs<{�g«l�ʪ��}����1�/����f)s���X��ݹ����c�ˤYx޼��%�6�5Y��h6F�n��e�׃���<�3-b&S��/�ff֜Ɏǒ�~���܉�ܖ�6�����{�mM�o���3Wr��з5�/5�֛��>�xX
 Oc_G�W	�L�����>ۗ�m�8c�b�2�0A޵��O�;�='���]��[/�j��`)"��İ�|���^�k]�v��!�ݞ߽���J�h}&P`n�����Ƈ�ߵD�06��ss��u���ə:y�w\�eS"���Ⱥ�=:tզ�h͏w�y����:U�/���:���:[�7.{��!��XD]�IJ9d�M͋��g0�$����E���6(	�7&�ַp��e+�f+�;���{�ZA�XJ]������N�2��F��RE$�+�8�ɤKL�g+.�[RnGmX�"'S����$��*�ˣ�/2���mq��;�YjA�,�,-ǂ=�T붭�N]Xэ-�ܤNU�n*#��'2W*rN���8qP+�DM��yՍ���~^����{�����{��y������{�����������x�ǌ<xg4f�d���8�����^	�������	&K+u^id��i�ו��vgr��3n�w;L�v��0��Z���y�`Q�(�5�4���$l��%� ��@㤤�9mRX8�4�p��1I�XH�!�qF��#� �%�MQ�F&䬲�'82���-�uu�Ҧ+(��w�����b�|�>G���D�T#T�mO?�|$�Æ�؟��C���SR�6�er��ά�9M-��J���� L���i��a�B����0٤�#��/���f���#(���I�L��,��Z�%jHUc�V<c�>z�N6�rG�gd�i�Y�3xg4f�d���8�ǎ��x��� "����6�Sk`�1Y|�ϩ�&�(�"q��gI'�
��J�&Ȉ����I꯫�??~����Z��eV��l����~��qmE�.Vp�<��C�ㆄ~�ѿݭa�~�fd0��?>k�Μ	�s����t��3(��<h�<xg4f�d���>>:f�zYG�Mm�D���NS�y�[��g�����T��iN3RI������i�q��Z>��};�	Ha�Lm:�%�ao6�Ɉ�5\���&�m���0�~�ӳ�Ki�ΉaS��#�4#����Il����0ҫMSuYEܦq�-��0ۏ�q�^t�ƌь��qGx��}=ED��K�U��4h�)Md5��7��tHw�$��Y>�؂� �����\2cSԫos����6l�:�Ӕ��껖�0�.��ușk�Zѥ%=M<gU���F�	J; �0D�e��a�y	M	����o8f���kG��\��f��s�v�iC8e�i��xь��q�OG����>[����$M`�}�t[U�	=m�ܭVv,��diִxb^�Cr�����٦�e�K�c�]��l\)��)<�t^���sp�Rම�3��:X&`�uZ���ʭ9^�c� Y�)�� r;9"*��ڪ)XF���+ht��෇��|���u�a���8n%�)���S���N�B"nv"`����2	�NTDw�|H�LJ���� ��Q�<��t��=7*��:̑ʮ�l���>:x'�'��L1-j+L��s+-���9���v϶����5rT�u�a֜i��6�κ��:d���,�Ǎ- �BG\v}q�KܒV"nu4��[ᡂQ6"dJ]c��|�����#����d��\:'�<���pK����!a�P�����[��m��e�s�H��4�RA���8_߿�eh�+�U��p�y�#��W_����J}�b�I�Gx���~��z�,�$�Ӕ�?:�ϝu��1�4�#$�4��G��
��Yy�mӬ)�U�����j�Ms�˔�(�>��mS|�#��M��{�����K���	���,8�]��:ؤ����
�S3I��bȮcXX�Lx|>����#��n��T�2�o�E��|�t����(�L׫�Xq��z$�n�Zf�B֍�Q����y��uן<�ђ2N8�O4�w��II|�D�*��|��fd�h����=6hK��20���?�3��0��"ܸ6����d8r�z:6&wM��-GQ����T�EjF�l��0M�Jk��:j�^3��hl��;~�U��������jG��>�V�ॄ<I�x�af3xc<i�F2FI��W��u_~[�c|�[eMF���	&�;�[��V.u��6tԑ�J*�7*�0��Lt�N�;��a�kb��be���UƮ+�R�e�⒭;�I$��Vޭ+%�M5$��r�jJӑ��8��T[��_/��D��JZ�nxy^[x"" g�J槁ٞ��D�iO�l�
`�=-L'�}M��mw�]GϢ�-e�&��繆eΛ5�u�"xN�:C�>�M=j5��i�K93�H�"#�^a�v�4����m>y�3xc<i�F2FI�i�Ɨ��K޼�i�j����-�hz������bwȦη�b��V\4�ќ4����t��b}U�|��f�=����};5,��n����b~��u���[��v�8JG[vv��~�D�:���Ιi��r�O��y��.�|����E{}��?��Y�<��8g���(�X�$d�A$1�d�F3�1�+n�ˮ?<���δ����0��[��$d�9I���f��Q d`�bdc(c��B0c�!`��H�Q@���K22F!�c�4d�`���3Ş(�<a��8�1�0f���h��a�8gh�4��Y� ce���p��ac�1d�C>`��e2�ZT�
2�#=\]�d̬�_j��S��b��hBY���`����o\�M�w�uD-��4�63�(S�V��Y7���}�LX����(��������J	���`�b�<֋��K�[	�F=�O�n�A��똸��x�r+	Ɖ�u�լY�u�8c��،O���m��2�A�����ˬȽ���|_x�Ξ;�M��Rb}�f` ������Z�&�<�m�}���u1�[�(�Z��ӿ{�j�Dere�����|	�t�+����M�j����w����>s|��O?&W,n-��6G߽�{w�&�2�{�����#n\FmEҾ��3d=�!�X�u�����D�\�xI��⭓D{�?����;h��d�YYy�����n�{���m���{}�{����wws��{���~{����{�<a��x�ǆ34��u�iǞ|��Z�D���J���SPѮ�R�&�B�zx*j�G4[�WȐ�6R]1M>F��$��\<4lЛ���J%LZ5�3
Ե�)�j)Cޏa�a�&# �?N~१���a�:%�<����3M�)$�Ֆ��S茰���̸�������<2FI�q�ƗR{Ъ��D9���b��E��jy� _�<��K�����6��Y�ɜ�>u�.��+N��KmV�H�>u{��M	��B�{��iu�6p�ɢI�&
0y����3M�*v�4�}Q'!�����Z�~�6'��M	�7'�E,)�&������	�\_����0��3�0���Ǎ<2FIǖ//������G��
�]�^d��j���H98g�LŐx��Z����$����Z]4�µ�RU�H���΍������7t���:�a`\��ٴ�^��J�B>8+c�m�t] E�0�	,N���G��Qv���ٶD����en�<>>�a�=<'�E����&�Ây,EU�]�x�Ѕ�����o��3��N	�x}>������#ӥ�3���`��S�򬦄~��)�aO}�B~��$������F��L�Ð����K�D!�=g,/�"���s�'i��p��<1�y��:ì8�N<��y�ܤI)r,+!�Y'́��@�"��Lg{�]f��_UV"xrJw�ق'Ӿ��\L&�'�聦C�D���`9]}�i֑�F��Vm��tgO��~�0MçU��l��B�=��^�V�.�愵
���X�$�VY���s�y2	M��0��9i�X�6���-������W�u�^y��<���[y��u�XqƜy���kJ��*�D��}y��L��8�==1X�6���8�L7O��w'5���R�`ĝ<0О����q���2q��I5s]n�(������O`�R�j1_C�l�3��k��ޕ�y�W�yH������|�+;G��F�C��,��q�4��i��#$��g���N����V+�k��[�U��n��v�U��^����>>��&�ٌ�ۢ����n�����Z��Y\�#�����|=s��L������,�6�3L��%?yn	��(���y���ե�_i�4.�E|_�>��%��$��t蝃'{䛗�mޏ�<4l�g�ƞƞ<a�2N8��4���T�S�a�y��Mݬ�1�5��Q�x`*��ylv������w5T�$¦ⳅ�e���j9I3�4�QΛd�ܛ4����t{%�%�j�+Z���UU��kli:�-��)[Mji�l��t�4o��V�a�w��/ne](�p�*��
l��9r�)��'��SF+U����/cL��iu��)K=N�V�Ϥ�q�(|"t����ۻ�36�+m���k6���}��=�Ϣ!����*�ݪ�N0�θ뮾y�<�o:��qŜx������*�B�ڛ�.^��)������Y�k����6�J��#���IRr~O4�-}A�����C[��r���fC��xb�L��yC;�R���n����v�#Og�~�5S��KWG�6��NaC�_�o��Y��r����,���x��8�Ǜy�a�q�0j�T�*D�|�X��y�djBrA��Z�b��S~�p���nyY�j`}���O�����h�/�El�nMC��\������S���n��t���7ql�\���e�ӳ�r���SF}�qwmSo,��y��m��1Ð�W1Ku���ns�='�6�VF^y�|��O<㮼��\|�ͼ���8�ϙ�-��˒�-kX����U��z�'�����1D�����9�!�k�#;�|e[f�N��ِ]JSf)���!C�ߟ!>�.ؕ�9��kZM4��2�i��,�&�ֵn�"��=��Ơ!���~�"~���314�<2rD�ڱ"$�a𔺆���M����g&�a��O��F��a���4�>�������ª�v��>��$HD���I$�"0QF�>/;�>q>�ȹ?�,#�5���b�Q� �HlH������&�dsd��Qa4��� �dA*����"���R�S �D2D �A�P����$dA � �2 �D!$B)BRBUB)	D*�A�A �"`�	H%T%!��BR	HB���� �P��"�"��BR�BR	@�B�� ��!!b���!(�A)�!R���!)B��B!QP��BJBR	JB*��J� J�2 �� �dA� �dA ���"$"Ȉ#" ���#D��2"DdD��"ĂDdD�FDd��2$#"0DdD�ȈȅI(#" #A��`�@F #B#"$F$FD�ȉ�D" �"0H$F�"2"�#�D`��F�#A$�#"$F ��A`���0��0H"2"�#`�#�#A�dDF�Ă#""0D�"0DF	`�bDF	�Ȃ#D`���H"#�#�#`�"0B1#A��2""##""0DdD`��" #"2Ȉ���ȐD`"#"2�0A$ �dDFDH���H �dD`��FD���A"���DDdDF �dD���A"#H����1$""#D`�bA"0D`"ȉ�"A"Ȍ`�#�DD`��"$FDD`�A��D� �	�$D�� ��Pb2"0DF��`�#"0� #""0dF2##H��#"$� �"2Ă0D��FDdF����A�F0"0"2$FAdF��IDR��"R �T�""1$"DdFDH���H2"DdD�F�2#��2"#��"$F0ȉ���#" #"2	�Ȉ�F "A# ��d�F����#"A�"2#"2#"$FD�FDH��2"DdFA�H�!HHF	$A$�P) , ,H#+�A�H�H��ABF$��B" 1IB@,���bB" 0@�H�� `���ӌ"ƳcP�B!)	HD%�HQ  �2 1"	HZt�BR	P�%!YŌR�%!J@H�"	T�� ���BUB�b�A��B!)BQ!)J\R�BR��!	U�"e@� �	D! �20�
D �"��%!J!-�BRD"D�i*@�ADA	���*!)BT!	UCj���D!	P�A �A��0A!)�BR	HBJ�!��!k*�BUB�HEBT"	HD%!�H�0A"dA�$A� �H�T!	HE!)
���"���d�E!"�)
�J �D �AD2�H0BT"���"B!!R��JA��A(�B� �J�A)	U�TB!)B!*���T!����%*���!*�PA(�T%*��"�)B����"�)	D%!B*�	HEB�P���J�B���B��B�JB!�P�"� Ȃ1 �A"ADAD ��"	`� �D����!)���!)�D%!	H%T	HD*R	HJ�!*	HD%!P�UA!�%!JB�!*	A)B�!D% �B��	HBB�!�	HB	HT�!��ʺBJBUBUB��!*�QBR��EA)��* �A*��!	P�*UAJ�D%B��JB�!JB��%B*��T�JB!R��%!JAH�`� ȂDD%!%BUB��%T"�B��B��D%T!	P�%!JB��d%!�P�J�B��J!R��J!J�!)BR
�B!)��� �AdA��� ���%T"��B�R��"	b Ȃ �A"T����P��T%` ȄAD �"�����T*QBUB�P�B�P����A"DD! � �D �20K@��JB����"	PD%B!)��JB!)��!	HB�"����!�!(�J�B�P��BR	P�*T!	P�%!)�R	H���!*�	P�%���"���J�BP�*R��HD%!	HJB% �%BUA*	Hb�*A`� � 2! ���BT"���D%AJ�B!*��*!)BT"B!)�*��D%!J�!�HD%B�B!*�RJ�!)BT!	U�*��"B��BT!
�P�D%!JBEAȂDD ȃ�GR@	����5�lp��:�F���3���V�P #FBETQ!$R��J�&߶��a�2�v���|�pk���O�)xQ�r}�f������!~i��<Cp���6���m2��(Y�9t�j�|v]k�lk�4(��/_O���bP������k6��(�"m����^�O���T<D��J��QG��"1�7ҏ�K� ? �q���)|�O�l�Au�3���0��v�'�QF"?#�G�B�PoU���B&�}Ex?àb6#�Nt�Ow�%%'�1=e�@���8a�����7!}i��[��^�Є`H��_��������H*�Q|.�E)AKȪ(�� �-@ ��j��Z(���*�ؗ�x�mj�?-إ����?���L��=A�SA�vCPF ���$A�
��PD$�� �@Y P��Pbc��B`.O��@w�H�q�����4P.�f^w�����"���@"(��'�a�`6�5{Lx���o���@b@<�9� ���\��� �G�����Z~	�{D�|BE��B�@|��+r��5uN��9G�QGrR3_gB���5���u����� �͈����}*�����"�>��>�H� ��;�KYN%��5a��7+�FF�0HQz��](A@�ѭ�	2I�lI,�X:���"

�(@`X� �6Q�� ,1�s��)(b}iHP�3�1���6#h���b	�	/�����TQF�0>RN��ԀN<���QG�-�/G�AX����j����!��=Ø��B��	�;�yj	�zӋ@oP��z���H^T�C���=��]��K�Ev���D�
�y~�z�Eq��9�l�p|��0��7&��7��)����	� �A�"��!÷#yx!t��\PP��4��G��n�.H'OV�{tMQHˁ۝�X�0L5�pؼ���� �(��&�v��䤪N)�����6 �5�m�x�g l2rMh�$�B�p.�J��G�y ]6&��D���w�z����ʀN@���)�6���7�Pj���\|0��)�� ���iOJH�ʔd��]f����.�p�!�A�