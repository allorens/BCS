BZh91AY&SY��!ڶ߀`q���&� ����bI��        j=�j�m�I�٪�6f���&�Zj��l�M��e��mi��b��cT�X�M�UUcM3Tf��IV������M�-�`��V5�mh��}��>Ǯ[j�E�Z�UmFZѴTڳ[l�,JM�Pc3��im�`����h��V
-mJ��m4��-4�2���m�-�hU�`5UJ|��ٱ[s�ti���\s�1��1R�u�Ef�5��Ͳٍ����іclm����vԲѶ��cZ�m��0�IҫS-[dٵ�3M�����Z�kAR�    w�,�u�'����8�.������v:�j�m��Vn�컵���zz:�O^]�{�5�
N�eop)ҽ{�m��W{���]T��f�fmEka�X�ؗ�   s�E*J
���utjT)/�^���f��7��y�"�i��s�RJ=���#��5T�������ZSٕ^�����X�ן}��R��_}��ޟI*R�{�镖-�SR���L��iJ�o�  f�Ԫ����>�Х*P�����O��U)�G�z�zjJ��=��UJT�>��o�|��������}�B������ W����yW�}�3YP����}�*�H��O���%�z��MV�  �>}JU>�������AU(^��>}T�J�x{��T�_}O���ʥJT��}��7�RQ��m|��(R������RU*U]����Z���_>���T�P��k-M�6Ͷ�-Sm+�@  �w�"�F*_y�|��f*JJ��z��PQ�O��|��UJ����Ӿy��)T�����>UO��K�S�=U��IO:����J�Vy����h^�N�7����*���/�Zm�k6lm�mY��U�_   �>�%R�����TPJ��m�����R��y�}����k�W�}JUv���R�U�����ꀅ�L����_m���	��o���QT����>�T��｛SX�$ڥ�f��QXE|   �ϟB��H�{������d������"��}�O@��/u����R�ϵ���N��׽������ޭ����D�$��mjƴ�[-�|  7�T�$5��N<�z==�K�:z��:���r��A���n�E5Gs������;�t�ކ�:4+ǞpTebV���5�h����>   �_ ��zuB��{ղ�OA�wzѯZ�w��xPOz���n��Ѣۧ2�����p=Z����B�z�@��F��E+�Z���   =��
=VW@�kμ��
QF���B�f�6��޼q�̀oT�� �ޕ�z���n׏Z����ף�      � ʔ� �0 �`Oh�JU$�      "�����j�      O�IRP�&   i������J�      JI�R$�dG�i���� Q�$�_����?���d����}�r)K7�����͆w��w�;#�/~{���PW�u���� *� "�� �� ��C����_����j ���U�� ��Е?�*
��?��������ɘ?����`�O�2���<d���0������0���/�>0���/�>03�/���e�����������22�0���'�l������L��x�x�x�|`|a<`<a<a<d<g�OON0�2�22�0�0>2�0�`��'���'����2002��M�!��	����������0�02��x���a3��x��/����22>0�O|e���S�!���	�=0���!�!�/�C���C����C�_�'�'��0>2�0�3�'����d<e���C���_�<a<a<a<a<e����������'�'�'��S��N1�!��	�/�'l�����00�2�2_d<d|a|e<e<e<d|c��!�f<`<d<`<`;ox���/��02x��'��0���!�0x�x�x�x�|e<d<a<a<`�������x�x�x�x�L�2222OOO~2��2�0=0>2���'��3�)�	���|dRe�S�O���O<a�G�U<d��&P|e�S�  T|a�C�@�A�S� O<`A�S�AO<a�C�U�xȡ�(���0*xȣ�*/�C�AO<`@�/���2�x�	�(�����x���"'��0"x���(���/���`�C�U<a�C�OP��'��9�S�DO<`D��P_D|eO�*�ȉ�A<d��O<aD�C�U<e�̂2�x¡�"'���0�x�	���E<`�G�@O�	�*'���0 ���� �� �2�xʡ� ���2(x��̪2�x����0 x�� ���0�x��� ���2=0�xȩ� ����|e��_|e���>�x�f�C�_O|e��ǎ<e��_�<a��_<e���O�|a��<d<e��_|e��~3�/��02���/���200��x�x��q��C��C�C������C����2�������_|d<d3����_~���x��/��2���'�|e̾002��x����Y<e3��2>8|a���>0���������9?�}�|�������؅�cj��S�*�i22�ܬ���\�h8�&774�+PyK�q�ݡG�(cS�h�eF&G�B�C�Z�L���ͼ�m�rR�sh+��ϒ.h`�G�#W),��V�r��դTJI�����jӖLz�" \�4��z��vS�맹{Xd��`��.!��f	u����(0��YI�!L�4�[�i�R���V��r^ܬ��j9��Za��X2=�v.�I��s(8�b�mP4�M[Gm��bKZ��3��سa}	O�/��f��WV!ÖH�r+�����dT�yuAѠLLJڏjH$�%�������l��V�HꃂC�v��&�,�I��S�4-�[���zv=5r<l�Yr^�3 dm�Q��4�]]̬�x�CK�G��km*�`j3V�Z̭��"�E,ɢ27c��ς*�ڎRzΕz�KsH���,RIm<l��Y���2��pe�ƭ#�)Ōlu�-vE�9�E=m��l3[j���%cj���7I��bwy��n!Xekb�u)/)7�[>�ܚ�$����Z���V�q�$�{(V!���_��W[R�q�	A�ws1kuq*`�t��.���� ����O2�fm�\�N�Udr,{!�J˕�,��D�2ˉ,7��<i�(ZءmV�^�,X�3Nk�_2��5+]jded�Y��]PQ�M6f
Jf�or�[�Zr?���J�@�-g\XE�?�!�.44�V�
y�љz0ve4.���4<��	T�ˀ(�r��8RwC����B�
��fFkg
lV��L�8d�	R�Q��u]����Z�������r��g\q$.��l���n�)dU�-�;,\��fi4Z�TU�`:���Ő�WX��͑�S�T��� ki芥A�-�f��U���%�����R�Pbܩj�<�4n0]n�����T��7c�/)��!��R�0ᶴ�ֶh���ɡ����!ARZ�k�4���cp�M���ɿ![f�I�C��z��1�ރ`	3��	�{�(HٰT���i��Z��PvQf��Y�C[�����c=�d��SQ���J�Y���ܫ�n��r�{V��,c�Ñ��ܡj԰�T�H�h)(_ӷ����֌���Mۊ�F!���X �k:Sћ����:"��F)���KV��8^�ʳ[V�*U)+q-*{*��
Ӆ�o]\�
QLة�LI�Mky�EE��	�*;��E& �4%[x+LYb���f k,'��(���*Ap�Y�Alb�lu�r�kp�)��6��cf�[��d���(���uI��fAF����[I�w%<���Z��w1�
�{���[6�Z�r�'a-�DL���,GaɄ9N�8�*�:��Ъ�z
9,�#�P����TL{�Ӕ2����3A��o5.�a(% ��*���չ@h�*J�(YB������l�e�ۍ����j*�6񸑬�
�ySF�OhH�oBm���+0_�FҒ��ybJ�T�P!륺��cZ�������TB%+l��p�(�BV��"sS��<3h�,�ݹ-Ap=��aYF�%e8Se6p"Xr7$@�TNk(��[�OG�+ï��v��5�T%	+��k�̚nA�dF�=X�$�]�)�z5"-�Y�K5���3� �`^kW`&豢LVG�p���n]��DM*57jU�`RZ!�J�۹�v�w�5����n&uE�6�Yl�I��&���u��eL�8i�pa6^c-
p�r�ŉMe�J�մ���e:�,����ZkR7H;ʰtVڛu��� F�& �bnZu�@��1RTi�ٺ��{�og�}r zLVQt�vC-��B���f=��	J1U�5���(60�ŊI�t.���"�J���&��>�g��-�m�,ҭ���z��W%M�.ؘ�p��ݳ.!����HFds4�y�m&��pb���T�3mQT�w �vV�' 2۰�+�&�Z�(�f�b�ޗf��kE�j7b��3wi�"�F��[�M���z��6��Sh���t��zv�Cy�^�HAVv�.���mk�BdF�5#p�<qI�Dd��r�+�{D3@���mH��FI���'l�[�@B�e`9�$j�A!�2��M�m��zݢ��w
�5�n���汖�7�V���|1��Qz�%1�֕w��A1*Q2�b]hb��s�|Aj��>�����nX�l67�S��@���[��z�:F�RM��=*eƍ"�ܲ�Gz1�2����iɶ2t!N��i`�v^�0�PD7]E&��I��z~�B�E'�sym��mބ���f�h�����^�,L���V]��8�e��Y��a��mCV���Vӕ��/�D	s	+1L���I��˽iS�]D�u�L��݋�+�v��z����9/]�*�S�ɕ�pG�@f��^�V��
jF p����ጊ���*It�)��Րu�X��
̛��`` ���c�\S%�Ж �v@͵3DRx��4au��3�Q�!�`��I *7If�Ƭ� �70im5H��	d� Q���w+E㩊 Ը�Ъ�ʍ��c
�*k(f�$U���mQ�m˭�ѐ�HQݶ$xs@	T�-S^�ٹ	�r*٦��KA�ղ���+4K��6-�R�1k�4Y�t��j㰨j�2��ӈ���+ufDaF��A#��/�%����IBf ��a.���bU��ԓ����M�R���$?�7+1�$FSjz�ER�3i�3mY��TT�6�u���p���?�9Ae��L��V�cJ<fUe��[Y�ē�,��#Z��a㹇�-�C�a���O.��4�l��7��gl��06���9`m���z(B�6"�wn��v7C�3��Vip��)�~��`j����[�7P7X�����6`��~J>�D�cz�F�۷˒�L�E���R��%y�Z�����ݭL�� ��&��5�k[�O�F"m��f�S/F޽����V��EWib�[�'�T��D���%fm�-����B�f)碣�*]�&� �eF%��p0*+DS�wwP�c1�l�2�5Md��C$� �@K���Ŋ�TvTy����_��lAu72�ŵ�ے�0F�׊����v��6TEvS����q���&<-��ֹ�5�9�I�Y��aR8�1Y��ö/:�R݇2T:��yPm[�+v�I)�+3fHⷮ��9*T��cu�V�m  :�l-��zݵWRԵw�[J\�̴���\� y"�f�)@�����b�'ii
����G��1��{���v8��d���[`�I\�-3K�f�nBO�5�˩Fn� "ڰ�Rz1�QA�l��#�v�V�+�."��S����*o3F�j2��Xf V��A��2�YI��-�כvIj�e�ilʐ"�m�("$�Af��2𻣅9��%(����˅DJ�u��w&�.��^�rn����e\qYj��U�u�L�X�ذͼ�B7�ы
mr��n�k-���A�u��jD�]=��
ׂ���j�d�p��P�ʉ�=Ս�7�S���j2�\5)�K�����
xiEF�TamG*�R@fÊ�2h��%�e�lM� �.��֚:�FR��r�N��6��ua��Rj���yžI�J�#ɖvi���'I��)�zҤ�����HFmh-^���,W6�n��t�m�t��L�b�I.�魨.[�2���*���[�%+m�:UƂօ&�P�r�4�����hP6U�n�Q-��!���N��V��,���n�SehC*mmm�f -����(
�������XPƌ�y�S�F�V	RƼ��Ⱥ	��7$�L�O�Q�Ic�ёҚՙ��X?jG�]��I;�R+��u���j�m"��v�qݫ��6KKu�`D�hH�(D���n��\���۠��/RGi�V���q�PS���kwz�+X���Fb%2�+�iK`Ry��-��Ge[�3o ܕ�P�E�e�W�L�)��p��YN��EᖩdR��Iґ��$)���j��iH*�#���.�w�n]� �b�Z)(ޜ�4�7IP%��7j��"�˽2�}  d�(ϋ4sQi0�;���`ȍ�ہ̵�����iT.��J��u��aQ������Si
%�ׯ�𺆰�xRTA�j�DԎ�jl�+ׄ�$J�dp`̉��tʚ�������n�`w�V��3bT,Ma�c
z����gsE���j�n�Ӑ��Vb�ci��%d�x��׀;�A����Cլc%��M6+p�U���`�t�^xS�ɫy�-)=a�2k$1��p�q!$�+���1�[�E�Ӡ�zq����7W��]�ޥGN&S��uU�ͣn�8�3o!���͍�,5a��i�YM�vU������Hh7t�B��u v�]�fm�R�`*�nRp���f���
:��)��#V��+$�㺶\[M��� \x��4>rj�vq��e�`Q�$X~���4Gٌ� J�"j�q	���D9*V���]!۰�N1�i�%�j^ݍk.�1��3z]A"߅������Z�6s6�� �7�W�����K���Z-0�(!G�lha`m�-�-ǘ�@��vm�*c6��V�e=�i�F�;���6�l��
,ۤ�AHL`�j�V��f�ZA٫�0�����3r�d�F6\��^Ԁ]*<�@�e�P%ތ[B7o 5�m���b��-3NX�	���*эl����T-��IWYm�����hӱy���������@s6�5�g�|���+ƕG�(��1!y��j��r�V;Q�-��`c'4(�"�@�VH��Yv6ʖ�Ґ�S���ǎ�7!�bb�O�������vZ;Ia�VF��Gf�D��,zM �H��5�iV�s!t���
��N��
���X��K1�a0+
�)�Op�t�f�7Mb׌J����#%-��d�93P�x͓:i�N�WJa�[f�3�$�*^�R�vi��Ӡ�"&]��F�Yb�9��)����gv�Yv���JXmm�
2�V���q�F��*��	�{�Jf�%�E�y�ܒ�LZB��� ��v�J2R�T&ҭ��^"$8�D�9B5�iތتE��ۋm�Ub��z�o���eS+bڐY��%�N�U��J�1��!{�V���{na�P�%3�b2h$ӓ�٧Tʲ75ͦ���Z$V��[��oa��T�Hf��ձ'��%�T�ٷ�Bг��]�2�j[#,̶�����E{k5�'1�ˤ][������^����yZس ;���;gp���#2�E=	��ᬚ��"�V�i���	u��]�j�O+�+$�W:E�Z�wmʙ6�V�#��@�j�<$�Kh�n�9�j[�s��H
J#0�*9�Q�RkIr¼W�Zf���}m�w�Ph(p�TvV|�Zu�G5�ChV��re�t3u$�݋�#ݖ� 2�M�6�]�l%r��N��ب�PTR�Էst�"0�N�k��6#�d�vK�S-�n+�5v7� ������b�1Iu�n��b,44#�� �m��6`-;d)k+p0���x�
�Զ(ޔ�5,�EFk��� �nn����� ��.�L1]�o1�<{z�
� �Kj��Th�!�D�ݢ�%�2�[�����C�?n�c���K�A��D�+J�r�ԃ2*�[�qY�6����){[�v���B�f��j�v�N�r�-a�PU~emё� ��ҩ fKp��
WA"ď(���ai����%0���m��l,Ǫ���@ECNŎ{�ͦ�tԼ{,VM���686��}��\e!W�ҵl���z��QkE	F'f�R��]O�|��\��Z�T����Rd������7/(�TT6�	���H�
&�MXo�la�`a�LB�j��|�hۤ������2MpA.�l*��^�P[�1p6x�nS�O��> "5�*ۆ�kܰp�:�5��'֋˽�Y��D�>�VI��ڎĹ5��(�Ё��t�f�Ƽ��j�D�>�U���	�<�^wI�V��ke�V�=۬Á��\ɅP��f��հc�t�	��<nz��;�@P�a-Q0��:���g��P��#YxO]M#hW#��B�4��~v��Դ�Hd;�:YY�a���	RIע�y5HA��.z]�ћ�ɿ;!�JS;?K�e1Y�aR���gt3NV�CYi�6��]�?kG�kS5^52���G��Ƹp�"�S��goh���}qBB)�V�+;dq^"�Ewn�����W�C(���mGF���؇�e@�E���G�G���V��ǆ�op�;R&h� �@�$�v����Vjl�8Ipa,���2��1�x]����͚�Ur�{������MXg�w���JQ�'C��6�윫��4��%ۦ>�]�|�' :���c1�Z2_���]X��f��H�T�eڍ+,%̲Z޻�j�����B���/ig,��ާ�&�� ,
�ȲY�262�lCW@=�ةp�fi"Ee̲^k'N�)��_���u�7TѸAF��cAl���a/CB��f��lǸq�����ø�JI%�R"���Rk3mj&�'�&}gK��.z����Ksʱ09�=P���q���A�=�.=}f�Iv��oh4�%���h���VhC+�n_M�l�L�I\h��e����k$��y*V�b�oQ�U�zr"��V�0���W���S���J0���x��8=�:a�����=_����9��@���Gyx|W耘������Mfp�P�l<'e𺱂��In+<��Ԉ4�ɇ���t��46o{�Τ�N����[��}Tp�R��ɋ]���{u�&M�歲P�\�=�9�e��7��W��w=ھ�RAۢ�:d�ղq�Ir�N��\B �=�{	|��X�t�&��� $��ǔc|�Z�Q�Rl�y�[!�]Dt�%��Haf��+|�>B����1���$�,=�-�����<����!%�z:^޲�tnۨ-�X"��m���끜�J۷`�4�ƣn.t6׫U!� w!��T{��@�i7vٻ�(Y��r����8T�R[Z(���5��E#V9�μݮ�Z���{�HfE[�:��6h�m�_Y�r\�ז�d�x���4���(�Wf���;٫�BZ7�F[��3W��vSܒ��"O�-�8��fr�2[-�2�S�:�l;vQ��C�EX���9�h�it���'��,�z������)�]AVi���m^�	��
=@�Sqbw=]t1]����oP����8%oV��YF�;&Gݽ7�U"�\�j���r���zbꓲ>�'崷wϙ�	mv^E+r-�zV�/x��ŵϋ���6Vd�Y��K�YT:��ڏ2#r��v�PX���ꄺ7�u�<t��u���KǺ�n�v�d�7��n L�{�L=Ƿ�ː�ݳ-[�#��j�������Y6�20hU��Jԫ�}���l� m�Z�"t)B��u�}�yګ=ϑ�C4t��8+�-�h-��J<�TVZ�����M�C^���*��V%MT��(>ଛ.-�p��5�]J�:�P�;t��U:��<0<�i����"8S�ܩ�^9���f�r]st��9���6�F��]���wtgfb�-WQ�ǜ�4uleA��E�}"�(ρz��7��8N%����3s[YF�{7Q��M���wT5��"���V�5�8fL9������k�����XW9�����B=�7����|!�yذ�`���-��`s9���D�r�1%6AMW^8"�K7��]��:�w	����嶱��oC�,�(�����Y��/5-�:�ӓ�DxR��#m>'��v?��,F�K�`E(WG1űk�v9E����h�l/��:/Zr��*p 7*n�|ظ$���(�wN�@I�\q�7�u�����2�s���:�
�+Q���=�'GOE�klD����n�v�=^(3��ƇeaھkO ��f�۹��]:��d2s��e���)T讲� �Yx��\2����Cw�v2����Nkds���[�}�v͙mg0�$#Y�i�˭�']Ӊ-͸P��q��Y�Y{�-H��+r7��d	N�SǤu�D()۪L����Y���Z����#4'R�)��o]v#��*v�b;>�f�p�]>�fpj�㮛�_X�����!�=7�w$�c�:�p�LkN�>�0������tUX��Q.!P�5�Tl>��+-2܊�eY$!��ذY�z=�3��`��d钭�guv�R^������2�����x���K�����r}�u���/k��V��J���pTY�˩r��v2齦��lm�=c��(���7�����$,5(��p����w��)GE���]��S�P�D�i�e�
.��n5V�����V�uFr��1�>�d�zV�$i���� �(4���'{�(ap@E����ʙ�V�Ttw�!8u;�$�z��ä�}��F��-�J�t���^ͲI]Jv1�T9���J�I�
�B����޶�X��m��h��H�&m_��{C�AG��urv����_G����Y5[Q[;�i�a�G�qcu�g�j�y�s���k���̧iD/e+�u�fc�8��{;m��{g���3��<� ��t���TÅ��&Q�l��5VeY�����[�G[�
�D����N�-�ur���kU-�Z�InX-b�Ǡê�����S?b)�T���7廮�t9-�e�^-��t�p�*5����@٪�gƔ��&��W�>�Ni#�9C6�h���C�w�ivCٸ���}P��u�:�T�b_3��P4�U���]�a�;[,v�,�J��֦+mL#��O'V�X�0[Y��l���
J�>�!���+9N飩R�{p�`Q0e�k*G�BZ6o�����u:+��74���#36C�Z9R������R�khL!c�T]�MF�O��Q5�,f��ǌ�7���ݹ�eA*=5��i���N�h���wD��D*<՝�*��b$q:���N��x��.��M��k�w�����h�J�Z��0-Ã6m#��4�C��v�<�k�/�'��.��S�_��-4X W0̢{�I�zP�o(��?^?��p��CʻU"G���f�9a��vjCV�b�r�Ǭ%�.᜞'u�zԅT���I���09M7�����ݦu�9�[w[د��s]Ԅ�Hj�F��Éz+
�
�&��%rӮ���42:�Rn]ft���\��5lܧ>(u����>�1�s��HX˯�e�#�8��\e��PTL�9 m�D��t�Cѳ:���0#�r"�]����,�s��f��`T(��/7�Ew%.t5X��
��Z���g�8o�M[��q�5��
Rߍ�qn��G�h��{lR�Rw]���չ����L����Y�$[d7N,�n�P�ur�j���	�*�~����W�/�0{kz���<�J�5�ʁ�ŹY�oKr��
�j���9��]�t��)��wWNo4��M���E�l.�)a����M��r:�s��.�wa�. F��h۷�i��5���=���Q�P�����u���0�͝��si�ڻD�P��b��q}i��v1�J02�/��#���Ww	]+nWnҥ�!k3�����c�u>��S�{;]dGd�k�7�c��]���wnP^/���;MHۼ��P J9�֢�:!���T/8h_B\�bHrt�{�����ﲸ6�3}�l��}]�Gne��k�EH�B����)%"�<4a��H)����"Vw9̣CK��(L���N^E4�}ȼ����S������}��+��z��լ.1��/>`��\u�i����ʷ�3F���#�Ƣ�l:t1�i�u�o�5�,�\<�V�m�J�3Q�5"�-�� ��Q� �U鴦\g��݊%NK�Iݷ�Kz�qtF8ʏz6ʔ��:�jGaZ9����U�pF��d�u'�^�ZF���
��=�>\:��ѩ3v؉X1K�v֠�R�@Z����;�}�EV�;�m�B�F�(%m&��嫲��/u�\y������TU#Z#M�|��$*[����]<|w��mƐ�N�6r�-Ns;����b%r�L����\�7�n��1��UL�C�޾�N��=<�L�h+�$��ãNWV��;kn)&��QJƫ��I"�@R���f��1�\b�_@M%�f�\��Y�_�mR>��3�N� ���vE\����D�Ϋ�U�û�Wj�_]K�s��+�ZP�q�.�Еd��:R�r̬�]��ˍ)ł�zq�V`�od�@)边�w4�ұ������7�ޛJ�.'��P]LX=�u�"��{+/�l���X�6|ֻB'oR��zD[ײ� �S	�Y��tt�c�@#`$�#�!�Tɒ���Jv�[�%�£����)�4/x�{B��ݼ�����]�;n�{��I��0�)���jj�9�T����q<�Dݨ�L��C(i��oa��us�=}��D���y��x&��s�,�{^uwl�ʹ㒌�Y;j�%��g�:K9v)���t�Ă���G>$Z���kX�������q������u�vk�-�!�Cк,�wm��oX�룰�m��E�� ]�Z�vYv�fQ<d�d[���-v�k{�em�I
P�iV��Tu\��#�Y�P�ܧ�_s�����ޤ�m����)}��j�4�A�,$IO����d�=@����M��o�2�M��0!�]�Te��� ��o]��:�h�UzF���dK�M�9ҁ�s�T�e�+tZ�tީ�lٽ�jLW�Aa��n���V���ĺ5v�� U��c|�6KKev>{b�ov�֮hj�ܥ�А\�Ǔ�-�w]�)��Gl=�mh�,�91Z�. ��s��CI�����|��θ)��3q@��^�Ef��S���)�~���x[*^������4�V� �El��j����4Wj�쮼�p49a�W��f���{�i��b���B�K�d����R�]���H6M3-ʶ:G�S��D0��Y��m�3�ܡ�e��rN�)�`B��4�Is��S�Kgew>Z+!�qz�/d[�Wq¥p�7a���e�G�	�˔Ӭp���ʋOl4�%�D�+��~�!��yAis��a�����I�c��KĖ�<���J.Q�j�e�]>k{v�K�wQ�{,�0Pq\et��7�Ȑc쮮)�iHwU��P��p*j��R2`����X�k7�T���Z��Dݞլ�D���t-�G_*d��]ޱ���nXs���+6������
F����l뚞�Kؔl�j/���-��5��#��%<��������R��±^R�ۄ=L]ƲvP�k�ǡ�W8:��*��fw����	��΃j�נ��w{ ��Y�"2�UYM���j�O����-���t�N��yg,�aw.��|���`߂�~�jc)@�*� x��r����, �Zm҇�nd/�7kfc��ӯ��a$:�����G��>�C7*r�(Mx����0�������XG�jޮ��쩺y y�5�j.��ț�wyZ%�.�B�:wo^ru�I�Js3���hN�,[��e������Mqʓ�p�wWb|�,���M碦9G&�9�����8c�����b����]�>��u9�}[d!L��S��������4�,g��X�lIG%����̶�l�"������g/��~�-�wP<�r��]�s�7,	�u��3��x�xh���T���ɶT��N)nf㙎��!7�|���TGsm�&2_q�70���McK���"�z���-8w��vY�{,�۩c�xjP�QU�:�}3f�*��L�O��xZ�l:ӄ�A�o*�&V�Qζ.�XL!V��tߎ
�6dTLɮ4����=�h���T��He�C(���cvlu��]y}�@[�s�ig'�D�h׎^l��^�]�u���Ĳ�E�=���6W}׼޽�w0VD���݊�KƑ�M��2�e&诵 -=�u��&�`�h�>���N��\':�FBV^v�l}b*^���xq:"�s5�V�Lr�A��Bvi�8����o��8`�����@&��g9�4�S�=��r@)/Y��I<�:�I�M�6�sn.��x��Vu>Q�x1$�^�ב`��4*x{i��ɉ��=���S���.��[�sp���ΣٚEc<�dn�vK�|���B�I�vi]@q�]6�Qz����5}�Jv���,�R�ԥ�Όf�Z���ɰK�����;`��ήՎ������}\�oXj�Ϋ�4��(�h��c[�j���`�\� ʘL�`��{����]E�1�
�]��'�5>�8�k���=�����dX��*f��yPok��]-�Y&�����V$8�[z�%*>�7�g�4�vo=��j��No�Q���@)mE�7�������,8�o$C"�-;�oXw��oug�h�]�[-8�`�:{a�r�*�P�&�|����*Rdq9փێ���v�c;s���xM�B�	��hO�ƺ����K�C��$��<����g_F�+Z��Y�d"g>WF���>t�뵕�m�b�p	x�Ӊb٩m���t�F�F���"A��&���ƅ�e��{��VzS�L.K���;S�f�+=Libɪ��w}�L/��M��#k/ae��s���5|t%�]�ڷ�KE3��Gl�N\P�(�C
��W�o�'.��s��彎�&��gxM�3f�$>��Bj鯻���#����e(x|��v����+Z�����`���ة�Ǖ�}]mt����}/8��E6�d�璭W]����37���BZ�z[����k�tە�v���w"����ÇN}�f����r�V�"�����T�e�{캒��V���)v�Cj��0�Ŗݫٹձ�|�>�N����4�T�#I#X�鶈�$�u�3OSr䠍�����q�����ܲ!���`�5h]�����Ad���T��\��t�iD�2�m�0�L�>�,,H��A�
>g�@���7D��B{ViFVYC��� M#�*���%�LPb w[��̄���J��U��T�x)�	�,<�
�f�����F�1�E M&������4B9^<O����XdsK�Kc"j���9��Ӧ�iN��[IQIav(9����Id�@@�QU`���N�>�t�um;�t�x�'��D��v4UD�iк��E"I�����&��t�:*�APd�) B��A'��.%E$i#[VR�a��Ut���J�5i�l�V�t!�v*�
��0�	Q �h�uSz�tj�Y -5�����Ǣ~J�����݊m�I7�?t2�K�T��@|Š�r�ɤ) ډ���L
T>m�(�,Yժ&����ʿ�>�p
 P�@�A"~c��$UC\Z 4�ܮ��Ώ�o�����������t���~G����v)���EQQ����� �������|���N�*��t�@��n�1��b�E�j�{{��\xޤ{�.��Y{�krn�L�
���{jwΛ�����$˺Y\�������f���a�J���|f�3�G�*��!�h7���&K�N�׀iIZm�,mN{O]t]���W�o"�ƪ;!FL�L 测F!^)������!��QS*�x�I}T��"w7��k���=g-�&Ή����b4*���b&^��n�h/�sM������f޾jw�~I�".�-6���
c�Τzj�t�,�:j�G�:Ɖ�����4Ѯ]�1�24���Ջ�y�c�x��3�KYʰ��E��>]�]9�ktp�,�.Y}����Ƴ.4�.�$��Z�&��c�]���M�y����g�R��5��G��K��bX�ʉ��؉�Ĥ�VI]ʝjɵ3�	��Z�r�S�Nu%7u����]��v�u!N���J���:}j��~ ,�e�����#�^�����U���=2ھ�n�ʜ�/�-���s�MN�K�5Ձ<t��l�����J��qE:�C&���'��)�p�)�뺺�aZ�Y����Q��G�
.��!)��0r���*�#�#�9p}s^0�����-E�ʝ(cNPY}[3գ/w���|>����>o���������>�����������}}}}x������}}}}}}}}|}}}s�����}�w��}�w����?-L�`	;7�x�U4᰸<��zn9��I��YC���}��[}��	�u�ݾ��D��P�H�IX�e!9_-O�
F�nJ��fK�`W:���WS�2*����@�=&�u`�{�!
l�-�Mܬ�B��D*�^d��:����FPr˪�`}�0k�F�Ø�Jx��)2fP���>�sy��V�]pJgq�7� �A�;�6z]�U�3X�\N�):�6�()�5r���
 ڑ=�>2-��ݙOq���=�F���06�.ݦr��C!�D�yŎ���UX;	�t�9���Zy4d˔�9ą���/D��j�3��b;V�ǜ�.��)ӮB���Riɮh7���r�}h���I-[m�;�s�S��n�Ծ����s5��y��d�F�qs+w�JR�����|f�{.����^�5>�ˇ%�F�P�!:r���k��2���U�ذ��	��i˴F>���D�ෆK��NӫG)�R�<w�������	/��x�TӺ�'.���3�iw"V:U���s��ِꝅ�� ����Gol��ǝW}6�s��f�3y���#]�4�8�Ϻ;�;Q���`YC	a��u0��߿|��:�:�����{s�����������ϯ����������>����x������_______�����_____^�___~�����CK%r|�/�_��;hl�R%���](��i3�]:e��/7*X���jl�kJ/�_����h�=�A���~5z�G]&V#]6W�|9C�F&�����z���nFq�Ղ�P׆��ʻ断��{��{@�S~L�����#�hm�Д�hc��+A�w���x^��;�{[[2�G֙C��-t�׮S2�7�j� �͞����-�Y�����}��<G0r��{��ǜ�D%M��(Z�8nq��>�A�s g"Y6f&݇F�Z=�4v�]�%>T�0A[�U��6��>�u�ӵۚ�)xq���T��D]�νK�G�0<�����5g���嚋�WK�Wo��gE�x��g����J@��h�mV�vU��]1J��+zNĕ��*�����w6��Q'ݼwv��UL���DhŖ8��[Mc���{So�4q���|���Sp�`k��9.aP��I9[����t�>$��K��|)j�����]$J��%��돳n+^5m)�s��+��E[!��tsHXE�!�5�iZw�z�Rm*4�f;���(u<�_^� .v,�B�y�@K�'b���9��U�W+u���g.;�s��o.�֬�"wQ$%Mv�z�	��]w�y󻮵�77�^�3����}~������������������}}}___^<x���������������������������������r�u�xp�oN����{<���iO���{FR�Q������҆ΰY����ѱ �%Vf^ռ��H9a�7ie^���ʶ�V( �F��\Y3���ꬽ��3����J��w;rZrP�@4;����
%N���k5��|��X��J��-*U���,�{���j�8E�p�8����`4�$y��b][Vv��+�9��f-X�L�n>d���ʪv�c2����B�JԬ	Ni�UfQ.�vH��oB�D��W�Â�R飷N �1R��ݓO睊f�9��r�-*kK�T�/��&��եi\I�k���}_(I"LK��c^��cn�@^�:O�3���V��q��M��qq޼������%���Z��-���ӱ.�O��9���2�ӣt���*��^�λ/����(��l��\%�ڶek:���Ѽ�F��gz�����TQ��+)�=Vw'-ډ�$��s+T�FD��A��L�th\�d@>iqL]�CE�wn�i�-!��E}�ٱ�)�}:���A���#��6.]���/ ��# ��D�Q��Ya>uxx�#��B����<��1U�R�/8�#���<�ԭ��Tz�.�J�T�]so]٫�uh�s�>�u�<��O�==>����������������������>�����====>������___^�________���������Qˡx��|���͖29�:��4�ďw��1u5�]�}�l�i�W�V��6q�snL�(����޸ H��|�]܎�`=Nޑ��Yd��m�u�1PH��g&u�CW�r�㳗���|�Xyo^�Z����N�Y6��;��y��˕۰U�t@�Z��ke�\�1V#���4/Y<E^���d�1����dN�\�57J�5)�;9�,��3�0oq�c����/g&ZO��ᵦ��z3�߭J�-S�_:�d���bG�	iu�J�[�(�)��B�s^@�Ͳ��P��Q%�y�W&�|��٢�Ҵ5u*֬T�+۾Ǭ��e�y4<��SM��s����)��F>C������ǰ>�d����JHX��E��ֵ;���ЬVPZ�k�TJ]��;��t�$�͝)���*(m E��v�_N��Ql��j7��(�:k����N3�koEڅ���s���@t��[BT�76��KJ�$j�\�F�l��8�f��M�O+,#��Kzz�	E�8���W���)��Fo\m�r���ul��p]�4�m��r-��l`w�~T�O ��D+cʘ�wGa��O���Ү��b�C$&��6�첧$)�oQ�X�%Њ�)����6��1h���_�����>>�������>�������������ϯ��O^��������������������������____=�[Q��v���`���`m�A;��n�4�Lئݪ�#�,���yO�d� a�j��{x���1=�u+u� la����N��6��\�W`��A�+�Q��s���=��m�:��-x��O����&�*/��c���ݪ�3q�૓OX�(�I�(	}���͜;�;����l�ɶ��8­a*ں�S�D�sv�CSa 1���������{ +�������id`αo=��*L�ݬUΎgp�ɽ�U�ks��
�Ϳ���կ���4��������dwN��ǱWi��F��jx�9]��cO^�ɢ�R2*�xA�i����#7�Wud��i�=Y�1����5��J��$U:��	���o[p̹r�6F1�N�3�첞����O�荒-��
�4��BZR�;p�]�yCrȚ���KF�(5i�"�	��:6�P��u<��7k[��:�{��CջT�uI�l�4�G��N�(���}I�|�ͽ�T|���`VFc/\tT��5:�sĂ�T�:X=eD
�/fn�r#צกb�MqE퍏���q�C%#:β�k}x���yI��9p ���^���Ď��z��+1QyUY;��HŰ�q��cl��F�}��JcX]X4=�НT��٩yθ�=GM�}>_z������������������������׷���>��=<}zg�����������__________G���ר���u���yաӣL\�;s��v�
���ѽ�PX�Zʻ~��(LQr��ջ֡��#�w�Z.�MF���3�X�OR�1ڍ�]5	|�kA[{xIM
p�t��B��Di4%�O�V�*�5�KoTҔ��V��$w�{mUn��]�e�EN6>���Y��0R�j�u�#)0x�Ȍ���XC��-�hi�:�j�J�r�Äv�ׂ2l�JXVwE4��ќ�L{�.��VM�5�E�mv��T��;�K�k�,�mdR��L�uX.�ׇ*�Ǣ1Y����u�����hl��f��Ҩ-��gxf.x:[���#{d�3ҡZ�[F�+�&�=w��x���ic����U�r�C��
l���2��(Aδ	W��%�+k�l\�/�H!���[�^+��հ��5~��YX���S��s.Q�8�9�(3*Z�9�i��:yz�Zi���c��l��i.E͚K����+���{�n�X
�x�h���)��%����i;�&>�Rx��r�<+h����Aǎ��"E��f,��������������z�Kjſ8�h��vh��:�*�â��>U�����vD�]���v:���#���]���Տ�l���� ��|�6z��,
g����U�5��ǿo�.����oϽ���=l����������������������������}}}}x������}}}}}}}}}}}___________Y����-u�W�h}2�op]������uT�yBV�5yĞ���$�[��V 5��صC��f^��^4�4_?��T�d�� �1�Y[�L��@��)���:1�i��:����gc�,��h�ZFu�y��#7�M�&������y9a>�}�$&�*f�Z����r�P�A�E^hڏ����[,*�V��R��ES�]��ʉ�g�z�UN����a�l�I���E�*�HeKu��Bn��;F
`[x��仢�E���V�id[��3��7y�t�=�$��1�څu���;:��9�5׫X�V"�W�s�<hX8��Ď�ִ���ud����:��Z����ۢ�o&k��7��N�QG5ǐ��A��j����I�_J�X+_&�s4��n��Y�O�%�u������Eɋ3j*����9l���k�6��E��|�r^��� 3oe�P�Ꮳ��9�${3�t�H��oGH�M�&���*Ww] 6#������UJz3�w!�F-�y��hQ�p�[Hu�+�vН�\2o�{5�!�FU}R�' �qD�V�w��u�����#���]/hf1�`j���t;n�t�u�ᶍ����W4�+qFњ�
�g �Hw��ɣ/Z�����g��p��VN�n�������F6���R�7{,O����~_w�������������������}}}}z}}}}}zzzzz}__________G�������������׏������;�Ϟ��뮷�f�:ԡ�Fow]�˥�B�D机B��t�����ʙݲve�2{TҸ-��{Y���nO'�gX��$�`���Q��vL�&:��<��Uy�ѝC�i{"f��;�I��C�K��ʓ�}UJ���n� :�}�mn�l�G���IMS�nþ�ze@���W�b�vS�D��	zI�<�g@=WC ��
�Ki?��7���Kj�*�Ye��`��(v0�mcm����mѨMA�iv�坆s�c����UQ)m��w��8s�F�F˝ �h��qHu�d�z����0�oSU�_;�\WY�ϻh��f�.&s��5#�"��s��,'[��8<N���/+H��GVݎ
���m����Z�+�9�1 ��������%v���E��'Ya�V4��'Mr�뷟3�{7
��@$>g���{��{m�c���n��>���Y����Zր�YX�q�Msʖ2{�a�e1���Y�ɼ�MY���s���W��:Ӛ5�OU���\�9
��nV�"WǴ��`=�,Ü�c&'eE̳����ff�zu�$`��;&��{Z�=z;�L���sD�mI#E���Cokf�\���U�fn���n��刭�k�)F'W�$n�X��74��R�UN��:��]K�׃{o����wx��諸Cxl��ʌ}u#O@TT���ثL�N�z%�]��"J�2`*L����W�\�oP�������C���_W�]�=��gr����)vBdՍr�8C�0���r���dw�P�ݥ�\oGI�wyt�Twz��S�	�,�N���]N�@`ƶ�J�����:��F8�!�A���̫\�U׫P�`�AՑ�ԽT\�(F�y��r8d4�ݩ)t�J�R�r=��0v�n�)�Mp3���kt�;*��b����y�ٺsC}"U��{�\seLX�\�u/)owUm�Mfu.��4U�t���m1v�<�VUWgdB	C{����Ϸb-�O"�Q�%�ì�/��-�Nl�Ő��h��B@W%�42]Dн���fC,��e�싲�ԧ��Dt�Ǻ�]>yW�kڽ��u��q��Bu7�>pU�k'C�A�P�ɩ�����u���z���
�9'��w:��21I"F��u�ڞ�����:��-��2��6�'"�*�]g3���X1ϓ�ޒ��\ޒ���4�R�KW��b������\	s��}���2?�S��ꥴg�7 U����v�^v*BD�PVNP����!`��K��v����:�9�t�FrV)HR1�K"�,�|�]���_>�-U�N�k�s�K�,����9�)ɰr���s΢8����;�����Qm�ͯ���9im�2����*�ոl�o'���y6�!y��ʯ��������� |�Ч������������_���~������_�k�nu������Q�hW�1L�e? �^ �L���(�M"͚~�x~n>��7�r�TΕP;/N�5������7M�K��К0j�u������dk�Io",R�Hܜ�w�� ݀MN�����:Дgd��s%��9vtrV��}l*:�-h��%���[�5���elX���[�B�P����3c��"<��4ީ)�
W)��w3Ӯw�j�9�^�l���ɯ�4�0�X�j��nb�O,,�
�O&��Aah(�����1�ҧF�!�7]���w�N��)�A�h�0p���8U�Ie� 8�����w�ʷ�a�]�ӗ<]��v�)�-�u��R�%ε��l�(B�g�e�hmУ���q�v�Y�M�����Ӈj��\q*��hr��ze�:`���furPb��,+{�#"�d���j7V"�xQ���
��u�Uq�4�!R��:⾭p��Q��f�˕٧[Xx��&�nfsҴ9�>{��Ҽّ[5��>��;.��F"���l�
�Mp�D��Q(�w^]�-n�v�s������[]Q�'H��U/��Fɲ���2��G)�����M�]���RoX���9m�xM�[L�����r��7�Ͳ�M.��� �����򢝖a��m�`
�<	��Bd[�D$M�O]1c���$2Dx.,c��h�5WWN�l��h����n���]t���/w;#���}�ժ�98��q�����îu�*�cZ�*��:�D�Q�r�5�����x��׷��O��9����W*�Ϙr�ˈ�mh�I��sc�s�Er>[��QW�g5���Z5��C=?_�ooq�sʀ�妈�qhԙ�"���V{�[b�����c�qխ��՝V���Ooooa�wj(�c�-QD�|�x������Q1V��s�����|�\ƣ�j���h�m]f�:��<{|~���O���'�\�O��|�9%5u�ry���]���7{L��G�j����mn�._,E_�E�zs�����'f�дT�LsN�ry}�*�)���s��'�.�¹��t7DN�>]�gL���X.}�9c�ϝ[w�t�\9�X����~��w��=�K�;���p���:�n�pq�\�A�v؞[����5m�.X�D�F<D�sX*.��>p�δu�#U˫��E�9\��O���mق�x�s� �9ȍZ�3��γ�ƍ��8\ڃ�6��c[ƹ����\6Ѷ;�9�Ù���8�Ɖ�nQ�U�:�]lqC��6Ύ��ۜ���ȬA���{~�C��6cm�f"��d�w|�ɭ�����Z5���6���g�b�h��خ��ܴX�]G,�᭷#[�ʨ�ծ)b�n�sc���)q���
*����KQ��N�nZ+�\��u=s� +�X�d(6�󾺣�<�s|����Upv��r�s�u2ܵƮ����QC���ͥ�W�y��E�K���e�>����C(�t`\����ju%�|�nV�ެ�q��B*��-�B,R��'I K ]���\i��<j���\���}X�tO9~]�/wXUZ�s���:b7����i��{��W3�Dt��튫 ����h,���{�07�a+�1�J@>����T\�w�Kt3��{��y�����ϗq�&�Uw�oxQ��|_��w���Ǥ��J����W�}�A�y:���޴��j�Gn=<��3��w�����U��֧�9=Sj��b�	�E��ڏ�:�R꼛��D�}W�=�`��7ٯ���:���ŲcD��0ݼT����1R���Ӷ�U�8�#/0����,���{���'䶩�N�Zw ���j}���hLz���_���������Fw(�ǻ�C��.�hm�=��zM��˷�}U�`�~�j�e0�� Wc�Ӗt"[���wygs��ɹ]�j����N}�꒟?�:˪p��{�3|�!)�W�iZ;�X�[}P٥���v���b���Χ�M��S_|9�Fd���}ʎ��`�`�˭�إH[�@gSպ�uˡ6ڜ�Ɵ>����9�Z/��}
޴ԲR���]"s��K=9L�7�l�bZd�kά=D�6�h�v.��]�DĐm����4BW.��������N��	�:U��_�����U?E�~�.[�Ǘ��S��b}6�WY������t8�c����}b��^��Ɇ>��o}�rWǾ����e>O��:
��uF���)zq��@�+Ө�_m�\G=]�6��ց��u��������Ǭz�T{{G��oG�����l�������:_���ʟ%�b�u�z��x��{���i�Ysďo6�yU�g�ƍ��r$�5�]�U�/C��j{�7qF�ʶ'&3v�V"(�2P?��S��z*� �wѝv�|�����U�c���ϕv=���	>S���y�G�}�\�ɠ���o�M��j42_��_o�|��s;����)s�ݞ���Nx_�Q5�o5;－]�j��n����D����.�H�Èo�q����p��<t
�7Y3{��7J��\�'Sǻ����+���75k6�F�.X��-AN���/�)�:��*�ֵ1�r�s)]���>#M	:N�n���X$���@�U�K;Vڹ��>k�&ŷF�òh�4q��oZ�X��a�"9z�g���<.��|v�W�^�Fcec�o��{�}&� �'��c�s�%=����]b�m?��{���S��L�m�c�"���cª�^�}����c\��܉'���q廼����z�".��!��۹4�Em|<}\l$�wޕk�u#ga�}�i�){ �e���y�-��%�^3����v�\B�ǻ˺%Ł���Ͼ�xs��E�wj�@­�EG(�ZWݹ���pXC���G�T�~�oF7����w{}����*[���Ur�\�xӆ�wՙ�w{eq�7'-���J�>cn�|��}r#7�O{sf/ON���WT)e���&}b�	�ά�{�kP�:[�Uʵs�,"/��wZ�O����|U.y��<j�@M�juύ_�L#Ն�+;��P��I���[�z��zK;�>)��;�J�oS�཈��%����{'=ŷ<��h��%KWg-B��1^ͼ���7/C h���p�9V�ܭ��B�s�,(PYf�!#{�N�uu�u\>7Y������g�n6��,�g��	٩��گ��E9��+��z�=|pjaԊ\j�S�@N�o�GkFka�U�.�P��᧪�s��r�og��|'
9�[a��f�z�q�z���5T����F+��P���\nr��޹�f�͆�)�|o��59j}F�����x�j��~!��R{�|���ލE^/v���W<P�4Sz��{�q��@���Xz�˓m\�y��{�יZ|S��j�r���]���S��px���P/�Z�o%���q��^�Ӛ��Orᾓ{d�R{2�e�{��v�s<&��[�hgzmR�݇ҟuP��P>�+�_]�:�9�����^Gޙ��W�z��X=7�߽8�ٜ,�˻����4tv���1 Q~��w�ǵT�:���(M#4r�2��=�o���7|fƞܯ.9�h�����^���[��5Bn�I��;�^Y�I�6�����;m��Ϭ֘��nx�7��-o>��j>G+�݂GKo)�q�����a�v�07�q���XB:�j��(7���gI�b��N��c]7+,���Ɏ�=b�(��cL(B
foN�|FH&shk��liv����Ec��WYP�ge<�C��[Yߓ�[��C���0:�`��6I$Xi��A"ۣD���i�7N���G�~4�4X�
�������V�W&L�Q��`Ʌ���f��'������}�T&�*{(SW8ec]����Q���
�&�����=��]A�ϲ_�:�|s~�W�|�sធ߆c=�Vj�g��+�����/v��|�}ϣ�v���ewη��u	�2�.�{�m +���vO{��Ng���j���o�Y�*����0��i���e��텑q�*�o�{�I�v���}�U7��|Ӽ�����}�w�gH߾�kv;P�X��������Bm�N��_xPx����~]������ʸ,J�d=W�|:�Ͻ�@nC�^�ח���oO����`�M�;G ύ�~�^Τu��xwG��-�U�p|���1�W�9K���6m'��J��'�VGnW����Xޓ�`�� �fף��y�CT{�b�W��2�}<:sB�X����Ul�t"����@׏��Q�Q�Rڏ0��M�wv�k3�ѣ�Ă���Y��5���%�)u����r7��W��r�)�h��E��+AU��=����]����j�`7�MWeu\'rW>=��`�.�-�2s�{Z�����wF���9����ovl׬yw�ݸ1��N}����)�)_s��ꬋ��zxׇw�{#�~3���·�Z&�����v��:/�r�慎Mt̏Q��힍��xc��,��b��ٛ�c�k�Y��4>��{ߝ%��'���O�b���7���w&�{�
�=�v`��B�3xX7��������=���;�{�j���t̝^�t��� ��Q�k�N4&ϟ`�*����kg�U�	�|&�X_۽�$��&�靮�������)�}\�\#9�(bs���m��C�e�e�%K�/Fr��3 ^[�ﯲ����2�﯃��}�E۹�k�bݭ�}�A���:Z~Y��'�wU�O��)�����+`��SP�G�f�d1Դ��s�E-�-QΏ��_|�ί����~,k�n5
鈫OY��Nb
ej�18]��`����ߔ��%j.�dT���ް�ن�+��̐�.�{�+�BwmSu�s���r�o ̹d ��o��
�}��=�"��r���]�\�o78w-���&����V����wb>���)B}=�1_�EC�w�ϣ�Ϯ��KNz�z�x�^���JWS�݋ǹ/�]�	�`a��I�+j�Ӿ�y�.��~��~O�8��W_��h�����'��q�W����s!�7�n@ff������b�kk���7����gha�H}�7~�G��T�ȹ�B���������������q�J������O�KΣ���}��t�\7ͪ�t��ߣ�}�	<�oގ��\{=���X���%kt�{�V�:��=�\G���Փf�{	�����s���^��|�\�3ӰE��k�mN�9��d��I��<"����Ǡ�;�:�`�P �0�%@nW�⑚���jy�z���}�yi�~��fz��>O(*� �r럼��_�5\��֐�g ��Qk����d��"�6O��t�߻+��"ΪD�N�*_��u����Z��k-�o�9�`QW|���mVM'A���t�t��3!Cв���FveJL��-����_��U��4�n�Bk��=\�έmdo�CZA'נ*}׃g)6�s��K�N��zt���1�մ��m�{��:�1��W�7���R����ڊjS>�����ս��|�u�۷�PǬ��W|e��v�
�j������d��ǨWw���3��ju��y�����,���r�;n���\6��<�����o��X��u����uݓ��3�lvzOz����=,ש�{���{eOePǟTK�~.&�j���̓�O`�2��f�Sϳ��Ŵ�n�|���mA���S��G�1����4����^{����C�yk?Wr��y2�ZR���ݍ���ɾ�{��墠ߴ�.x���A�{����y�N����W�sWA .����7Mٺ��X�j���
6�)]�[ZEw�OUy����y�{�����T�fA'Xg��Ƨ{�Y�-^��Q�/s�'�R6�@���o{{2^}����b�Ŝ�/{e.5CuE���)��Li3�$�e��}�u;���uǺ���'<��b�-�.j��B�LCa;a�栩�[5!ӠR�� ���\��v_PA��Tt��8���H�k$usԂ��j��'Zu�gƤeB��c��.�6i��ɩT����-�,��8�wj��4Yn�����x���t'���ξ��w�ǉ6�^����ȇ3sӮ��9�V�Y��IV�9�˹�>������/V���Z�W�3�83�8y�s������霨��T'��>���"5�t��P}�~r"�K앏�� ���3�z��]��/�7���(>�N���i��9�L�[j���✝W�0���ZF��q��RL�쁯���4�JM����Q��49׽��/@�f�ҟ]=�p�k�z��G>�Ix�y�eYs5�_םz����}\~��vR�|��̠2��]�#�j�t�7|��ޓ��NS
�le�==�}��ߩ����u��mOh��﨨�rQ�0Ws�mX�|*�"�C�7+��Ϯ�f^�ؗ�T�%y�p���ay�%��.��)SZ
��ro49��=W��V?��Q+����>��^�~�w3�'��
��Si��/7���R�W���AH+�	V�j��@���U�1��;�T�]��]�>��������0�O+��<�k�V>�U2�ٽ��ů�����Y]�Åk���A�ɦ]�a�^�×�8�
V採*!�é*�x��o-���"oT��7Wi�B� }���t}n���O��%����{�N���L�fE��$O�+	��87v��[Tw���m��]G:���ɏ�jG9���{��������N�cjI�b������n��u~d��g��9�'k���y���	���v�N�5(Y��	�^j�a��N'�>:�s�Wc]q��C^NW��H�s�������;�59<>sw���� ��[�_\�#��h��OmxI��%�g�p�Q�7��W�$gă����>��Myߣ4H�z5���޻���j��Ǔ;����6����L�1���0ь�z=�)���G5��>ﴙ�f���CJ�nV�uc�����~��u��O{~��3s�כ3�'������Ѥ|�l�������1~�A�}�΁��~�`ΐ=>��}�T�
�{󲱖����f~N�ݔԠ���.(�Z�w�m짒�4�B�����07�p��3ȟ)���h���z�6j=X��Nm�,:v��������K4��)�ʾN:ہӬ����ƪ��u��nP��K�x�n�os�Fڍr{�&&s*�U�g�8����\����Qk{%�Oa���F�E���֒2sqp�\]֬iU-�e��l*��HɣK��Ô��R��i�N�8�y�Ax����R�T����됰T�4��X���P.�v)�$���w�u�K;�պ\{+���s^��s{[��PI\ �lwZx�+]�rq�kes	8-�}�u2]ٻg-�6P=V.�F���g�VS��P�[��Ms��oK�jԲ��&ڎu� �[�n��CL�o)'��m��Eq4nr�x�}6�8+�����/Z�I�b03]
L�gF���r33&���\��p`,���פ.�x�t�C�ff�HNyW"ͤ^r�]De�/Ky�'E���L��K�ʝ'e��/�w���A]�^?����0]G�z!F�<83�������y6�&v-u��r�cw��qO�F(�����u/�L�_v(�AXhZ��>�i�(�,t��WeE�:�_k�C����|q�޵�Re�t�w&ԇ9�85	ʥ�5� �Ӊ�޵�N���*�u@p$3��u���(�T�΅,�F��|4Wi�DMj���J���1�f�v��WK+SxȳPj� ��(�!��M����;���ݱ@w�|��9��s��O-Ҙ�/��s<�\��mG2+T����p��T{%�Z��c�����D.]ۘ�[fhj�cvi�C/�+(t�fd���rs���d���e�VF� �'LG׺֞k���WR��h��k�Ӎs�,�d�7'7
�ۍgւm;����"�:��|�pƤ)wrG��ä��Wim1e���tk��4�.|C乾�+�6��l�(����:V������sw:��q��r�P��j)�&��h�+m��S5y�R�uH��8�	���m�N�ѐ}��ٕ���F�æ���TyE4#�4J�V�j�vaa�ﭥrr�P���x�V1���ʰ�me�M!E�v:�}^c�fp�sy(�9�1��� ��\uII.�Z����m�)-��Yv��&Z�a����6�{Y	�䧝:�e�����W�����7K��O&����H��U��[�P��,�3�e���`N���^7�K����B�F6�uk��ʙ�o�k�X��y.�5��ך�mKz��������Z8���dgd���Fm�Ŧ0���bvp�*F����2���aG��i�,M�
�x��P�c|��X"sz�S{���>��������|7_-�GϿ�
<�غ�,η#1sli����Ȉ.mV�\����9=q8|����χ\�DS�N�O#�S?=��߯�l}�^luֳN3lD�r׃Ѩ��9���ǜ�3m��{ϓë��tحur����:��$��t�~?�oo6��w�U����<�}b�����mEUu�\1E�G{��53�\����>F*��{~�^��D۲�60h����1����-��ID�W���֊�J&��ۜyus���g����������{{;1�����673͝r�QTshn��S�������k��S�|��KQ�s��^箷N~=�^�ߕ�	�����TUUv8���6>�b"'��:ƈ�3uj��`֊�ʃ�N�����tF�d�߯ooe�:$���|�'�PM���y��UN�QM�%1SGEZ6?��Ƿ��h�\�*����w�ʪ��kj��Ǳ�3�y\�.O(�b�)�qX����)���������w:�J")��������3<�QKMQC[c�h���<"�uEQ�9�U����BRӶ
-��ÍiuD��j��U�F�R��4�M��=��[�����w���֝`���׉-	��G�6ԼP�L�y��)��J�P�����u���|�N�k2������ks���/R�'b�pυ��(ٱ��Z�f�?ؙ�����Έv�O��;�a+���w�ފ k�42�3�0Ģ٘7r��t�xm��-��ZF7�R�.��;y27���=�[~���.� ~^$�Ϻ�T����NF1��O��� v���v���%~�a�z��6U��t�+����h�=(�G%yi��*`W�}�.�rp��]���	D���7�@�z��r���]g�� J�a}M.�q嚾�DUc�n5J@{T���-��z.<~"�P.�����]q�nZ��[b'F9�#�[�tL ��z%�M��e��+(��2���d�����R�J��Y�ׯ��t���m%�rܐg�;=���\�@�o&+`K^�)�{�T���ٮ�@h�A�eԨ�e*��Μ�T���e��n�d �f5�$j������Ti�]t/9mcj����C�-x���/3�pL�_Edp�����<�|�c��T矘1�=� M�V8η��+�s��լ�=�����)�c�Q�~�3�Gx	���{��+�3�ْ<cv���R�\eM����RQ�
�6V��^S+���}��Y�^Z��H�6���M�`ޣV;S��w[��Y�6�J�αΧ]���[��ax������6���L�":�t�ַ�,]�:gK��(�Wd�Ͷ���sSP�p�֌��!�����¼=^�r��7�&�R[lr�����C�0��l�	�)�r��� �r��ǫx>��6�nb����Kw9�,����;t<ȏ���&�['�mP)k�����=���fr=� ~bӺ�s�0I!���`}���g�ݜ"�^�G���9��+Y��сX�-aU3��ٛή�=ϣ��,�?n����r�7��(�/R��j���Ňrg�@l��%ݍ����Z���a&��wi|R�
�����%���Ϡ��-pp���a�"K�#��Fk��Nj���%OF0ו����K������|HNS�ٚ��̑�b�Ϸ]�v��w����vn��D���Q6��T1BV~����k�Bh�_-��D��mvK�Fμi�O�ä��>W�����Kex�����D�馽��~��!�^Cٕ�˭�o]Qz�d�)��Чj��5�'�������ƽ� 8�7��>/�:<����L��
������@fT)g�xWb�f��ny�=P-T����]t,z�A�:�,�'����&�3���L����U�5ޘ�;����,��u�<E��YYy��:k�V�]m�o�)A���f���{���F�v2���������@J��ӧE�	dj�h�u��F[v���7�����AB�ow7�;Q�Z����V�)sJlQ����K�����=���M:,��@� �U$
	�Y��D#�́�#��RO�3}����"e�Ra���r���W�\�Z�������̉-��t�ˢ�ʊO���Jj��Գ��z�j��^���;�Q��DvcGvK���z(�?5�P�-'���\uso�儥y�r��{��\Ne����/�6�yA\q�k>���q�4�@��A�*����Y{k�<�^�RqH�W^׸�4�z��������7��}u��y�_��=�5R�Xc���2Cw=c�)���3#�B�7A~|�e0�jKqr��d�H�W4�l%K�W���m���-z��-�����=0���l�D�c��K��� �.(Y�N��Og-�0����*�֜EZ_&U,d:4��5���4�m{8���Z��$�p��t
�B��ʌ��1�gNmGs����������%�bT7�~���Ó�O�4���~ ��/}.hS�)�U%�=ڕ�Ĥ��Z��?�s�่r	tYgE;t����/,�v"�_j~Y�o���>���'�Ȏ�01�m���-�]�{���� ��
�ȇ������5�s5�h�a/��or�� x <{X��o#�Z�DIR~�b�`N.�ۭ�}�ޚPeiW�>�0;,'i�!�%#�7�h�ￏ_Ms����\8�ˌ������&���zļ8E^���<H��+����\"���R\ؔ�q� ��:`Q�T2M5�r��u�;��@N�+͓8�OlO+�LV��l��oztҖZ�L�Z�Ն�>�UD�q^Kr6
i����qь��Bҁ��#-�,>ނ�?
�D��|������L��(����T�VB~����?��;��a<&�jFs�nwL?T�����Q��D\JTj�u4j����g`(��-��{j��oR�y�Z���T�[X�!4Q��AWB��2l�}�
�Y������A��R��/$�{��|��X*��^j�X�7��R~��0���rw����F����B��.'�馷}O���ޘ��˒��Բ<
��I6�/7�֠֏s[%oW.`X�G���2[���2o8���mz�V0��2`H�5�r��_�"�{Ѥ}�{[Pэ��יg�!��p{T����K��n�T��Y'_�I���-�M�{���"Z}�El~�\�����p~//�V[P�	�Y2}zh.(u�`c=~�冀�00��GZ���5�̤s ��NK�Oٽ��i�=#�A��2~�=�-��6%�zӛ���1"����XQ�8H�uT˹
��^:ӕMb�3Wa��	��a��8���y�fG7�=e:�nL����C�-E=ķ����^=����_���2����uQ�9n��6��
�.qr�`u����vx<�t����\�%��A(��^m�\,%� �>�s�#�#7�Z@���X�Wb Bz~��y�0��E���`*�u\��UqM���'��k<�� uh�:�7���XX���<�0�����T�0ý�6�f�M#�SY�n�]ė��=��3L8�Z�_,�`l�6,��6��Ԧ~ K'�l.nʹN�󩔷u���)����cg+�>�X'n=�{7�Z�����m�z~m\\YץX��L׳�1��i�W��	
z����צCǉ�i���ar�x`Ҫ�^�^�;� ;A�������}��y���xY���	�+��&�}��ل{�3��jcƤ����F[�v�lp�+��f�&�πv�T%ff��r��}�b]�T}������֍O����D3�4���+s�^D����˼�W�O�&��J�#-�W�[S ��P/�]��k���3�5��)���1�W��̕e��ϵŋ�yˀ��~�boG?O��<9��]��ySg��Z�u2���뇵|�p�p[�D+z���W�A�:`/�K*@m�޹����,�Z8���Q��=��*�^���X�>]�7N��J2J�uzpX��&�Q�����ʲ�4�lx�%]�]ϵ���}���&Bj��a�KE\X���U�Zi�L����f��!PJpNsݗl��o+m8�}a�ޠ�u������i,��äT�}��'��������YP�数_txo��n=ØE|�s�}+g))�{�T�SV�ϟ�;&�3����l��K�ei�1��p~~>_)/�R74��vE� ��h~�K\������,�g�k���}o�;v���7�� dF�����W�(!����^��&>����3�Ѥ���ߏ�n�.�8�f!��ʛ�bo��#��u?�vy����^�!��L�9�?5u�@w���M��w�:/�)�ݹ��e���09�}��0��`��?�6~��F <9�w�UMIqRm��P�^EJ�����[���bp��t�7�,.w?/��<���pzWbU9ׂpn��t�J�� ���TXm�gA�,m�����4Nkg������@̬�P1T�Zu�egf������4���%����
o�N�`vx�IN741�Z��}�j�����]���(�YM�Ӷ��S�N���f�wj�te5U0h8������w;�N< i��`�q[���`�U[xX�l��%�|��)��o�0m5�"�{�����f�=�>�wt�{�ܛ������yn��\�����c,�i�d+���W����j�
�b]r[D
������x]Ҕ���`��k(
��'v�5P��6 �\@t7]B���}�R����:h��|:q���H��M�mM��4��{�1�K��C���Ţ�3'�(.�מ�н�r��8�[�ڎ RU*�	^�b-B�����T��(��4������X�����������aBΓJ�K���J���覻`�K�g0t�*����y�-d�6	�{�J� ��1N)���e�;X�`p'������ϫ�餀^�-3�p1�>OT���Z�C�꿪�WaR90.Eh���"��)#�Jix���W�z�0�F):�VP���^�{<��5\��O2 {9�1%�]4jk�4\�7�/�#���X��<���G3�Fs��\��ǖ܊�G&�f �]R����Jm��Dw���%������ABN�s�E}�m��ᕑ���d���!��J���	u�}v�Μ?�t��l���.�`�Z�f*U�N3�2��H!��i��/����3�F�&��@9�Z�>��@�\��S�^��F`��?j�^R����-1_��\p����"�\�8`��I �V]Z2}����t�n.^a'Zϭ��_|�>�����)x��]���ߚU���բ#K)lS2/X�Jp&�|d�;�##� �����aQ��h���������Pg�{�K�%�F���o���IaeG/.�X��ߣ�_p:�5�`%}�av�dd���~N?��kٍ��A�B�cmf;����D�xQV�)�Խ&�LYy9���j&�ۙ��ےق����	@d��\�7;S���L<�=Xx��[0��k\�������9B��|l[z�@eY�t�-Gs�����Yv�[��C�}�Wb�
�4#`D���,��X���N�ױ3 jsu�D^�oWtx�Ts�t��k,��um}l���垐�^���Д��+'#��u� ��0��'(����0,ǜZ����,��O^eHYS=�o;>?Oۯ
��M~��g$cޤ@6��`���VDV�J'�6B멻�0�VN����Z2���|6 Z}��	x�1��L����U�;�p"\��<D�r����m���B(��
v=���k���wj�������B<�i4���}{ >S�ծ�m���{�b}W�*�vGI���|��� D�w��Q���*i���jFs�n~�0"���i ��#�����s&��w�2���ͺ1�3���`{�Q��uf��2��WcfLֿ����l|8߭mi�ϥM��Ds0�ەm~�nSÁ#��������fڡ�S�z��
��ůaN6h�x��\�7���{�����%0�ձ��^�W���r��~>4�]�,j�@�>1��x�4�Ҫ���!G���Zy3{CY�\����%47�^B(��W�U&E�n�����=h+I� �ȭ|���Uk�}���Һ�`�oV�g]�#�ҽy�1�]R|75"U��4#�ջ�u�� ����w�}��n��=��޾�+�33����ξ��V<�>r�^xI3%��UL����Ҳ^���N�O������B�=���mipnJ;���	c��A���}0��(3I���ڮ��SM��rq���m��\M��Q��ª�'P��v]�x�����E� ���"8���"�_���8��5�����؜lJ��}��5�+#i���7�:)���/�&���Vf0md�px�U�O�n߃��N'�(�\R]a&+&��)�, 0��g�q9��Cv\�5�.u�3��qBĕ��?BxBK��	�7�d�v̷����͡sR����r���7�7ώm��zk�?�ְM�|��X���q|���}/-�qv^�j���Zz5�2]��s��(U�j�	�j��Glk ����@%��`(6�UEs�|��Q7¯F->�}�R�Z�J��T.#5U�n8L�55�nZ���އ�4"��SBº��g]�bvì����nF��mUW@�8�21�3Vn1B���p�e�9��	�*��3�]ټ+[�G��2m�vY���8Ȅ(����5�R���4�m�x�-��/6k�#a��H��Q���m����S0�j|���ƻ��I��ʔzr����V$�4�)����<��@�򫝽3`<ޛl�yJbX�$8�2&oV=��+E���p�r��̾޸�׽ ��v�f������qG����2LM2+վ����Q�:��<��O?#fBL��9�A��}��;PU}"���Bܝ������g�W=�0.����
xl�?1��@���X�����	+˵PQ`M��8"/k2wkCV���A��#V���24�S��^7�T�$
��.!�ؤ���H�#|��uM�U�&z�s�X����wK�B]���i�c�ɦ�K&Vʦ������|ك�cLǐ9�>K�^py��ǜL�뱌�b�����CLNT¶��̉�ܱq�N�`H����Z�/t��p�SM��/tf�×�����ZT}��P�!��N��<���TZrqu7��KÛ�[W��Y&���yKbj.��t�]�f��j<�����(�DwN� �(m���r4�7fƪ������z�i�b�ée�jހ���ܼ-vt5������~]�)��A�Bg:���[�f��
��9�쌇����e��đ�?>��'�S
9f�������:c(�h�B1���[rk���P��Ǟ]�j1�Hʂ�7�+�
�?|��|>B먭�Q6�ؓ�A�}yqsJ�=In�	l��N� ��{�*U"��v�6��I|P�6�E��s��r�묵�ck*d.�=���SwJJ��/#��R�L����;��ޭ���@�2�[a;����W��z �9�=�Ʒ'Mi�K�f\-�V�x1��G�eM��J�}ǀ3L��oeq�}ݳ!�2�|y �����Fʹ���;J�,pp�J�4�f�-:�G<�õ��u�ݻ��%=t��{C���g	�͛}Vu֦iÎ��t)��95
(+ة�P�� \�]5��b��r�)�Y!����O�YgϘ��0���7v!w��sۼ�Cc�{bu'�X�]Q�k����dx*=ǢB�%�9�ŗ���;���,_b�l^*K-W{܉�:�PZ�
��� Gy	��p��­��$�n�wCҠ��g��kMGC19��Z\�n"���X��c��H�:��b#X1�\}UƤ�X��� �U��u�O�R�Vøōk�dD�T�&�Y�|uHu�[�m+V*�	m�؜���&�����}",����S�u���Y;�J��\V+����h������u�f�L3�:�_H�P�YiV�غ:ǚY"�N���N.���h k8H�d��z��U����\�R�&����P�v�jjw�
0�jn\s�L��rɅ+(���PU���.=q�,	.�Lv;[�)�Xv�7N�mY�E\��@����!2����K�L��[Y�~����7�,i$�
6�z�eӷF��yr�lp+X���ֵd�Ήgү��Fo>q���vd7R5u�����:2�6��3��Nw^a�� i�����oT�β�ia]���]�z�C�ke_D7*qQ�x,Z���n5wD����Gpn:��n�Nu-���hv�'��̓��M��Aw;�%��_JB�=�͜��79���*��:�1b&���u1���N�:�*Bz$�*�"Gj�<�T�}MnW�}W����\�i�Pnn[t����mXd�Ob���`�{Z!������l������l����L��؀�J0Hh�MҰ�(va�\���/vv'ʭoF�}{;�J��c�م�D>�|�$+{1�2V2�%�U�|>�9>���.��^�}\�
����a�,s��Ήf^99�q�M^���)�ޢ��Ǆ��Q����m0*�#2�!����b������i:Q|ن˻9�����ɻ�F����0=�m��e�Õ.L��'/WQ4�f¯���Q�Rց/l�<�:tڎ��Gֻh�؈���a���-R�L<7���P��!V�|�:�'�G\ѧ���-T��u�g""!�m��vI�.�X�i���2f�I�4�+2���V@�� O�&�y�Vu�)���7�0����Hy�_oT�N��TE҉�|��4i�t	>!jI��b�7R;�h�aL�h��L"XT��h-^
,Z�J�0�*,ҁ��@
�T��u�ns�|��~���u_��st����գAHb4e��)�*(i5��9�17,ETEM��~���lGv5X���M�4�T�G{���5u�s��]u�]T���ʪ�'?�������l�:"���
#�b��+N�F'W�q��Z���A{$O��;.���oa�w�4Z3��9�r!��15�4�T�EQRs��*��D�ӟ�����w��Hw�D�E*���-5W,�nZ���TR�g������
.��`���
"�6\��5�+MRrqy�Ղ��n�<�EU���q�ED���î�UA7u�!F�:�;�իckS�>u��QP^�^]\�"����]؞���U<؃����Ƿ��qR\�$�
� �MD�UE�i�jh �in�I]W0�8���{{vb�Z���7��_ �ѵ��\�	��*��h�o��TV�h���I���s4��Pj�*�)��RF��n����+o�h�Q P��&��ό ��n�\��]P��3B�_Sd��VJ��q����|�h�3z�vC�S�s:���(!��t���#�s��E��Q���*H�?�W�&I��bi�e;�u�������H�J��/��Q��xJ�P��3�b��o�:z���=��\��0���X3��C��|c�kuN83l�4�*�ad1�������?H��lx$hcP��`΀�/D�s=�������R�j �v����)�H�z`B�[K��tn�G������5��Etj�(��DkqHp�h\���J��a�|��Ɋ�f�7q�z��:���om��>�9Ó�K5��k{Ѧ~Z�W)�	^�Ɉ���p}ф@��j&ߪ6��}��k�7��� "��w�	��M�Ҩ��{Ҋ���]8�7��P�����N�sQ��S�o4'������-���v��q$1���(1oX.!�}�m%_G�f6Z����^L�9§�,�˳�|P��;�se��b�/%x���m[м��ޘ����N�a,�+�7*L�N��#> �����%�PGT�}s�3��7��;ϑ¸��\z׹E�9˳�w�q�_/z&�����oMZ�e�"���%�����P�|���\,�,�Z[�8�*��H9��K���l�_���A�fv��	�{�J,�Oh#��2�ʞ̃�3{/Vԙ�L֥���Xn@a�s�WUw�#��tC������� J�����s���6�hv�������Ht��A6�4�Y�k�}gtc����}�9��~�	�a��&I�c�kw4�9�)��S�J�5[���E5�I6��o:4Z9,� +���T4��oi���	�~�A�Zg��8��^)�?`*}��P�f�b����vlk�L��Z�O)��Ӱ��Hl�C^Sȳ��&o6��m�&*S.�#4[������09�I��Dy��S�yGd�(�_ƤS�K�i�Z0��,�^�� Rd�8�0�P�^�m,�nڴ��u11Yu|bs�Hd�6��KV��#c��
�u�6;���j4�=���}�q��E�=�Qt2��]�3u(`��G��V�|P� � ���x�|����q����h�i�3>������&P��f>�r^�����l|D0��'�'�ub�.�r=�3/9�ƭ���.,�u�g����/B!��:� �F�Hy�^Q���E�j�>��˗�)@���#L�#�,;U�f�C�X�Lg?f�D�DiT��g�ਲ��ĥuUu���Z��y���� ڇ��չ����W2Cu��0ISl}�m�>���`Y����=����=Gؤ�*��SMD0��=�X�}�Ld�O�uҍ=�a`�Y���wkZ��U��>z;f�Dh��'RL��)4Ej�3�b�"�����yc��Y��*&�lL_ueg.��r3����:��~|��s����ϟ��٘���	��`9���?]��<����o͹}��ݐ�v��N���`�$ϩ�֯�p-"K���vHy�Gu�5�4��.�D@�h��NA]��]=�da�OG���D3��_� \U��}�N�P�N]~�������hқ��	���B0�u�W������܍��nWW�����u�y�_��Ye���%wB���<<���0�a��{�U�^!������{���o[��=Z���,�)�Y�JU�o�:�2踸�6�Ʃ�ne�R��`��7Ց28�^��^�:�!�ڤ�\�t��oT���J��?T��2�p���2��9x���H�C}����˶B��t99?S}��{�J���|fm?6{sn�u��vȉW�:b"xߖ�[P3%�RB����d�mg�1���	�DǕrsYvD��	�Ρhc��+����7����V��+��xC���D̛�2T��a��^�W�uctG#^u�Q�TJQ��c:���%g��sc��֌��`y�p>��	�����<���d��?x'[D�r�4_�[e��X����k�H�46���j&lE�{��o.WT����0�:V�Cսݱ���w��Շ����K��uH��b�/��xiw`I���\.1tw��y���߾y�o���a�&	��`y�y�����֡�XžM5w#I�5Ig�
�C�1�<Z�cF6��D�����
��e�.j7೯�0\F>�L�[��5pv��q���l}������:n�O/�d;k���O<<����7~쬂(��W���8T5���:�4�.��,��gב��q���I�^H��{����]�i#>(�p_`F�idV�7�w!r���#���D�Kj/C���/�U�HC�=K��Ͼx���J4�3Q�yO��d���*��������o�p�����'.k9ú�ɬ���"��λ�Hs�R�a�����bJߩ�+�?��|�J��crk����.�
X#zkۧ���sTq<��ЕL_T�+����)Kڵ����U"�$�0AGv�a0�5)����ͳΦگ!�1,�m%�m��n��tSLǐ9��]1C�[5=�������!��=?cK�x�����tRuι�?�E6%oNXLt���f��&��YZ��N���yvkG� ���rm�AR���>���\p~�K_<�Zrs����283L��7�6ۨ����/��QZ���u�߅5����b�\k�;���:���O���#��OK�O�d��^���u�隳�c�Ǭ!�h�n�+�1u%ۼT��V���p_TTy�;�J�]�q�(v5�+��T��
�:E)أF�>uξtg��l��̤�0���������>�4�I_D>3�4���&����ο�C��}"z]?^Ab����f�6 �1��,���7��i��3L �(�J�{�&�l��z�K�6>���Zx���8n��&[ -��um=���)�rK�	���]�H����a�Ցf\�O1n���}{S�1�V�����P��QB�\��^=z��4'(�e���hD�P�I#p݃ݲ��*���{�@�a�G ��K�t@{��y�2*��TXm��:p-ly�8��c�-�������㉘+n�^M�4�7$�o
�y����"˱JSȍ26}C�z�pu)�)l���)u�ZN�o����6n�C�-w�y�+�D,$M1K��ď��(�z��?�a�ʅ�zmq����-<A��g�
�:��^O�_�}5H��F[���a�;�1B��Z�6w��� 5ƣQ}��ǉz}��k F)(�W�0M��r�!_�:Ԥ{az^�_��#%{?&����t�=v�S�Vd}�_j_`�t�D{ҌZ�(DgG0�_N��T�覺v��Ż��-���r]|�(zW�X�m�� �(�]��/ڄ��ws�`1L)��O����͔�^|9p��L��9o$���p���
�ډ���I�$��z�1��G�Gt����>�������b��!�K���������`I�&@�e	�y����������\=E}��z��qmWp>�R��82���m�dKej�wy�:<�5Brű��#���{77<�o7�026
d�d9o��+�^y@��}�[Л�A�=኿(��+�T]P��;rٛ���{i���C�LCϻna���3�/�����I�~��g'��9+�k�E�� ͉q.��SvHw������g��y��'�cB���F�ʷ��4�Ś�N1b��Ƹ��ۙ�H�Z�?L�}�]�m�ǡa0����V��+HI��~��]�A�T�cdhƢ;Ӽ��b�@���|�Ѷ���$���S�f�m�3q���r�����wk�rP�$�DA�R�}W�=*��Ko��\!p7�E(�݀�{c��y1��Z�~�++�q��:����d�[IfzY�")MG�G�V_;����7�d�i����-�с8 �f�X�j���d�8�0x����������4+����"�!D�Ts�Cv�Ȉ}�a��/M
�Re�p����K�|I��j�qmt��A٨�Q�+�sc/.Nh��;=	�ƾ(��\j����K�����݃�K���6^>&�������1[G��0�r\�$dx�Y	d�	�NէÝ�a�"^���J�:H�5*�=���p�l�o�T�ƴ}Wf���T���f�7�Yhg��M��
2of͢��d��v��Δ��VP�bp;�͝u�߿<�ѽ��|���+ε����+�2,�3*L0!2,�3
� ��ԒNݓ��g�)O�V����֐3\���4��0u0��(�����V}��K��p�����i������pGצg60�S��u�C98�7�F�]��< �}1��,��@i��J0zr��Ebn�O�{ʠ��X���߾m�tg�P�����9�%�:zyWi}�l^��dw��m$�cS�ԍ)>;�^���Xi*jQ�``�� �E6��P�5G]ܩ���*��
�i�5jfǗ���&%�i�R��
�WkN��h)�-[����mf)�xtNk���L";鯾�J7ԜL_\�/CL������!q�5�ޤ��=��-n+B�L�72���k�v4�W�M@�+>tI�F��x�����s��u'���^y�o���Ǳ�#3�d�U��ճm�%fX��/�[�;��ُ�����w1�*U�s��CԬ7�<E�hs�a>�L���\�Z�WXQ�0��3Z.�����[���0��Ӄ��@��Ӷ��砠c��qJ����U)��i��qm���gMlD��V���$�z����p�y��ޓ�&Y���'G��]��i�x\�v5�N���0�l8F�w$r���pr[ku���+H��|th��hs��r��[���ӄ=bf�ܩ�ݔ83']����u�[+p��b��A ��Q�d�f�`�R�e�y�=�wƕ����Z����-�Y�wa�pO�1����_OB�5`�畚��r�2heut嵙�>w�E����a��
g��冾��<��8~�y���}�;:n�\R�}5��nr�O1����=���#܃�f�ZK�@([u��	���{��#G����p�}�"o�p�y}Ư[=�����xs��C�"N��(`>v@V~Y�bi�_�z�%�2%��V+_���H�Lն�Bk�a��O�ק��@.�;�Z>�=� �s��J���9�����=G��P�����<O�9m��UN������Q�i�z�G�]H�����ܻ�̵"�]�G���%��bDu���J��t�YE�Kڬf����	�3�ד���#�W.~��l�.f�
xg|��;y� 	������?�]v[5���$�swc�c�L
�u
f)�	Y%ؙ}�c���\�P�,��^e[�m�r��5��m�;Pނ��M;iⱨw����ϹٱO�#�50�ǖrZ8۪RvJ��o,�i�j)�U�wI�JCaBi'�P�Z�eA/q�Rd�L���^��O��03�+�)N�=�C��%�]p��x�,DQQ�?S�Â�=݌���-3��5�F�p�����M���/_B���P#~jb�����M��e3�k S8l���CL:E0���~�dY�I�I�� �� y��{k	S�c+nʦpҼ�[��>�5�y9�:8�[ɟU��9D��L�h����[^E��(/no��t-��3���
uNo!-�\D�m�+ʦ�m
��r���z��Ӱ�4���n��G���y���\���-��9�c�t&\��)?Z]B�w;0�f銚˸��+ǆuC>���D����f~wЌ-�:"+�b�:z�gs�����J#����b\)>�	9U����j5_m��^?
�/��DF�	K1��l�����Ӽy�~��\c<��~�
O�ZU���$�i�_�&;:�W�Ec��TMz]Lv��8�z���dNmNyt-��-Q}����6�TE��Wq�U�}2ҋ���9��V{f�G(����<�9/���;��>~���㤑>�}���U��g��=���~�^H�P�H�zA����0�Γ�sV��ڬ����6'�Z���YTZ�+eDi�cSZ��~������;�2y��+ua�B�\�Jy+�=�fF��#C){V}�@Ʒ�jNgQ�R��ٗIK˯KM!Z��~M:ʷI:����۫���EW[����S��ZW|�|G�`�۝�=nW7�C�M�;R�{�����!��� ��CW[��82�Z�Om;��������}�n�y�����f&@	�d �� &���|���~�G[��?���~�Ȓ�H�A�I5 ����J���q�g۪�1��M�G5R��2���/�/
ޢp{-�j��@܆�q&� O�mAK�b`��:Sś۪}6=�x,|L�ݱ����"����)P(�|ik�\�%{+��hK�p���E��B��:rgҝ��|}���jZ,T�/
��[�����YA�r��Ty�BeI��K�Q��55�)���)�>BL��@��%V�c@����ɠC^Sn�2�6�E]�p���|�ÆK^W-�L���o��$	~����J���C(y�L�ƞ54����B�[zm�n��&a��8o���)W0� V�6�d�n^>�Vr�>X��~缢�``<d�������׳]�EfV�8�6\��¢��:̧amLu4[z6��ۋ8�ϋ��Ƃ&�(�cߏѯ־no��3'�8T�am��^�{ʟ5_�i�HA���袝@��Z��W�ˤ�d��h�2���^�x�OZb�k��S���v6�Ѭ^�`�� <���]Rq�a�U��t�����y��A��N�p+z4	;�����aΕ�f�,��/^ui��W5��:���!U2>�Z/���q�d���W^��"�ܕBVI�KӢo����dĊa#�ͦ㚨,
x�9$���pw>�c��d���fƬv�*ԍ�(��%iǯykDwSkF����<�k6������Vg�,�3�E}Q�A���p����
 �ӦNW;t�k����
��WTw"�2.:��n���*��=��-t
b�gnK�}�}�#Q�y��EC�����+9�ޱZEY��g-�*<GA;VŨK˩|�|Q�y�u����YOr<8(sj���Jڊ��m�ᕩ��[Ȯ�5�yJ�^��cy1�m�%��f��]5)�K��X]�%�}��֨���|z�;Rb���¹�b�ڗ�l���	��mx�aK7�v�q�/�p"V��÷C��c�6+�´��7k�=�(�v���+��x�F	�*��:_A�wuЍ�� CK�[bLX��;n�.�5\��}�؃����3CR�;��r����
NVC�|��	�%:�v�`����]sVL�P�ډ���lN���T�fԃ�%��)�+#��f��MΨ]��n�CgU���T0��6��¸d�b-�[�E�j�'<TPs��ܢ�t�]�����N�*ZFTF��߇f1�(�!�A�*H���Dk0ӊӔ�B��IY/-��!��a@��y�iD���*�8v��� ^��a������٩��L'+2�|V���jBˢ�t7�I9\Ұ�q�t���N���1Wd4���R�,`
(���.c=��
T�
���g��0G�8ݽ�ѽ�dت:���[W3�cT%��`�wA�Ω�o*pފ���6�D:�t��$�wLY6���7�jՉ��	��*螃� 7��ё-[n-ab�T���\<��P�JJ�.���%��#����s�o��ם��,�+n��k���e��)��H�$�o��u��]A��VG4Z�)Y�)��h)�T��E�Gd$I�V��9�'/ ��n�Q����Z��(y����EB��e��2n�^��2vu������Nu&�yCX@�.�}��v�\yM)�1�I$|{��`�ђ�X�4�O/jf�s�@���(n�DL=���3�wEU����msr��\��pfvN1)�uh6���v�\�vp�fN�1wg%��/;�V�*j��w��H���o{��O�.�ʖf!ޱ|�o�n��ģ��S�Ukj�1�&=�i�h�}���)����b88�ˑ�T�<����C*���Y'�K��N�F9���L�0���K�f=�5�'Eݪf� 8�ө ����.G��c�r�
�|� (� ���|�U�gE4�Z��svl�0hu1�|�Q;h�劮k<z�^Ӻ��`�o�x���y�-4�SZsEG��j

��AUL�����|.���TQ�����Z��{i��k����Qr���՞=?_�׷��fc�j$���ti�$�ERA|��`���s\�h���Σs;m:�E9���~��w��9���.��:m�U|���ĕ6�EH[:�*��g?�����RS��>�&�r�#y/	".�D�W]pD�W��9"d������b�^F"������V�QU;gl�Lu�sr9ET�5�||~?��;$�����y#k3DSTN�T<�lm��1����\y7Q�	�������@O�_yT}ܞ��h�9#M[c�?#�Zߜ�M<�AS}Ë�&�%=�`�N�:ٶ(��'�u�MTj�;M�P���3����_�����F��7Sh��C�����<��C8�2�,g�A}3sN�û��%��7d�Ю��j�}-� f�y��T�<��
��Eff@	�Bd@�T&PI�T�����_7�~}�.]��y� �_�k���<��S0[��1R�m���m�T�p�Ln�k5K�k���1�=E����"�݈c�Q�ݬVU4��mO0����f�<�y���2�"s�e��k��9��޲�t�%}����%h0>�����dNgF�9��c��-�r���>��.mŠT��C�f@�d��Ɍ� ��z~S�)��ɺ��T:�ޕ�22�0�O�$���!�ڕ��i��8i�Mi����^������}��N��<���éCB�@��9�s�k��b�#�F���5���U)�f`f�`3��5�J4��e�d[�f#��8?>�0��"���rk��}�T�Ҫp.��`ߛ�ϥW�G$��������E�+ʸ����qι弫�F�{�T��׾��܂ZF�x���=�쳊���`˺<],iZPn-#���a���|��U��-��7 ��Tt���T��JH��kCR7/��ޚw ��a;0�S5�ɏ��4�І�u�B�K��/��_��]b6#��&;c6�ЃR��b��Ǫ:6]���͖��W*+`��w��˯�
�bӼ��t��vk��$�t3y'$k7o$r�s��z�d��OW�@96M��Y���y�>{�
�Ȭȉ0"L 3*$�)2�L ]u���_��t�a��D�A&Bm�*�6�/S�zd��j��a��w���^�L��qYU7X�Wi|�C��=����6醵�%�Z����Y�-nK�恐2��P/���W������R�H�lH�{�ǃS�
�4�S�������Ɏ=����{b�+�]c
	4fL�H��o| �S6���v�~�A�Z�q������key�0�0�<�L(SO�T�[����4�w-�Pz^yKr*m�^��j^ PxƊ*]���ۗ5���E�R�	63VOx������6�Z���ĖmG���!��cbK	O��9�Ԡ;A�rl�+/ F�y3��t�����wF�z���$�'":g�\�V�Aj��])����X��.~+����;7�Ѷ���g%�̞���-0GCȖ�]2�} �����A�2$b#gX&�b�=n�=�Er�7�^D-�K断=
�u�&Uݱ��%ᮏ���3��֙h��A�}]�Ǜ[���:+�<}ꐤ������#�S��C]��'��>��Q�}1>Fg�/b��.p\��b0gS��9�Hw��<�r��բG,q�3�R��7�]���i�9�:mV�2�]����9����AY��MQ�A�=c6wP��8�7�e������]�+7)tJS�a��uM�3xm�B}�V%t�0�(��CUYFù���lUj��K�Ÿp5n���
��`T�&QI�?A3
�)0��n]��{�.#�^?�mM���1�)֩�G`���H�a,��7E�*�[5[��N���;܄�5\����m�2i|��E��a���u�v�Y>�V�m�C�c�E���g�{j�:�-�\�%f>I����ʄ�ꚙ^r��
P�{b3..��N�s �Z���l���$˰,U3�ar�Mv�"� �Ę�gZ�":\r�X!\�8�j=S�]6�U�O���W�J$[��P��" WykE��C~1)�e(���{8}/,�] @���s�*a��P'T+|�1i�ɲ��*�l%�(��ŝ�׼L�d-�י��3��O6��@�8K��zc!�����ǣ���b}Kq�-zY�g�)��YjMN�3o|��W��I��-H�v��MƐғⷚ>�"�c	��^4�7w*��v��7�rj�k7F��3���r�u�P�����d�iF�ÝHja�SO��,�� ���f=��ʞ1޼ұ�k-��f��1�t�ʺ�an�4����uπ����,�Mx{n�9����t3u�=�oO&F��.e��)J\6�^N8>1��H�U�����F�]�ή�+�|.� � � ��u�<��~efMWrs�B����.�2G�GV�k;ݝ�>Xi�Z��\��W��`T�&P�BdP�D&A	�D���{�����o�������w$|�q��"�ȝ��p�y.��lH�u�DRH���&B[{�ʶ}�cDp����wfD1=�8�j��o���&�i�>��v;q0���lݫbsi$�\`��</��^�ϵ��K{wz4���+��?� *�*ʇv����ã�u�m�9hϾO�aL?�o��4��U�F⯼�������!26DiU9"���=|Af��|�&��c������@ـ�6ʝH�3�!����$��]�F
��掂)��U�Tm�ՄT}���+<!Z��N�����^a4]HǼ<,�O,
���c^;75�3���yN6��w�q�a��M���c�aif�(�+<��g=�b:�,�����o���a	����?_�+���(W.&���D��ސ`n��Q��5ku������RW��zT�kϟnC��/V�ڮ�kٗk�,a�r��&D�i�<OP5m��3���b���Iw�����\��0{�L��7��Sȧ���+z�C(|�25~�8�ˢM����t�ai�� �:C^[���g��z�贙�I����au���b�r�*.�Z6��h��Y����fq�iSL L�C�}����l��ۑu	h�π�d�ٸuڢ�ғYN�'��wv��%���+����U&Ef&	��Y`< o0��𫻾�J��݋Z~�ۓ���!�����֏�`����뢽t�d��C���l�~暥���C�(��뷸�wE����`x-�TUǠVyn�" ��������Y/� j��;!䌙W/6'�Sz�Z��Npȣ�1�̈�[�4$��^D��X�-^P�%����|wO�����m{.�.���;}P8=�3V(2�6c��yeϼ
��W�ʻs��պo�=~�!�*&�����$B�!}p�.	ip�����"���G��!�2�i��_�T�����бQ��[��J{�y�u�κAjŕ��C����S6��<���has�7�mW0�j{�z�%�.�h^Z堽����AԦ����a��E,����}�=��lF�F����u���%�ڤeƓ����e�),$b=�{.���1ˈ$¾^!ޯM�s�{��>�k���Ө���j��j��=CZxŴ�A��œ�·k�{����1ϼ�j+�[$st�D�1��B7k9��;���ذn�H9ba��d>y��cj�O2ar�6)��P�n��-�@�(?�ܡ�n��<iخԔm��W�0��T�W�'�q�,��ɹVZe�e�Omӂ~����g}^��`V�]<F�A�i5�gx>�����w�CY�}��giZ�8]�j�8�[x�m��,uME�UP��UI�Be@�@&I�BeD�QN�;�w���>�k�|?g>��0��"*�.��n�����LN9�Q1�tΐ ]�:��ꋯu��B�qk�2��[Sz=���E=�"��ޟC1K5Y���1�*"�S�gf�����C�	���H<;#�ꜹ��T�<!���LK���3�a/��3��u{����s�q�����r�Y��D@���[C����D�w�~f�[�dЪ�C�c�尫���d)b��XMn�-`q��{�&���Ԑ��*�t�1+��_��b�s>q�GL�b8�B1��te5�hu�7T�z����iN7��̱v�e5D�%��=Y�����s��K�m0��`W��j����a ��ݸUS"�˜M�ܫ�`���I7���F��%�J��t�y�C�ic��֠U���3�j8���{�s�8��ֳ=-[�{����)���!��8���C�Ol"#���c̀��;����n�A�����N.��jQ�� �ۯ��԰��{�N���+<�e?�R��I����c�ڪ��Ma30u;RK�Z��t��	�W�@�\�b���y����Qt�2�SZ嫾�{�G��
�,z��!2�eͳB ���	���^�hs�����/�����l���nV���rDF;^W\��$̛+����}{����;��պ��\�S���0(L( $�	2�L(����R掎fwa˛ߖR�@�\�;����2�8oU���WZ"���B�63�O;�)��*�uT�)�.�oۑ��r�ܰ�Sކ=��X�>����@�l,Mˉ��^}E����!���"0dI���_+�xWh�H��k�[��zZ�٬6�ܒ�U��g{{yTP� َlx��2Jh��ǜ�3��])���V�W�7`_��G�#�l��o��~���ܴ�#�͖Z����H��|dB��< sz����`\b�l��Ǘ�1+mR�b��s�=#k�3[�?>t
'������d�6�-��#���&�c�[ͧb1�'݂1��s��78-�ż��2N&ˋ�O��i/}
�ҕbfs�O�ls�u,׹�_��(!W��E��4^�ӗ���i�7;����0l��X��(;T,��<�uP3�a|���p�T$��ȒK�~���+��%�>�?��y�?Mk<�f��w��}�DG��ʹ��l��ؗ>�������Jqpj�Y�&~~�'�!�Or�'T��y1`(1,�J��Ŕ:}��YU��Ruf1������C�V�����ɩv���}�:�7q���LNP髜�[��fFFF<��|�Z���c��츨�����Vuu���z1��
ׯ6�Aw,:8OK����;���ם^���W;�޾��P?l" ��)2�@�ȡ2�L� tH|��^��|��~����~����O}p���c�����,�&G1�V��gV��	�9����c]�]�x;���b�� ��cԼ{��c�ծW���&����ۃX�S��G�2�»�nխr&�\�c�1��ϟ�*�yji�{]���������g�����U��椼�:���o���o@%�͹�"��ש)�
��B�t6��C	�|va��w���,�w���_<L�:xy3�&/e�����q�E�M���FxC�\��XւH��[��c�/]ɌȲb������m:��+��L�<k~�mOFK#����|��1Y*��X[�jD���H���3���4	�Dy�S
9v�����L�ogB��,η�|Sh�ǋr�ꪐ�U�c��zx�2�5��A� ��-��-@�B�Zk�B���r��`9ʱ��
6qgwd?mR��*�5Z鿋�ؓ[�J�:�6I&�S�H��z0�ߪ+���Yj�����{!#C�Nl��u*Fk�.v"u	|!bF[El]σG�
#:���?_wj���~pI�L�
�G�Z������ʴ(���[k���qƎZ�u��0�4�C#�>5�lq�4DO3x��X�Z��
P#b:.q���VE�yr�eɳ��Ts賖��S;�1�D��o���}�׿� ��L*
3 �����0�L��>}������_o�Z�xH}e7��@��@����n�.�8Ȱ`oLi���q�N'M����d���:et8{Q~�Y�p���񉞉!5㸨P_C�J���
�I�{��1���}ۖ��jw�2����o�;���9_�֚2�!��I��Lݡ&Ǽ�G��Fiq֫��mq�t3�hO�o���^ԇ�����4Б�ծ�����2��ډ�|��P%I��G�N��obg�ޢ��V�U��8�!I%1K��f���^�E{c�A������+��'�}���g���)l�r�c�=J&�}w�[�����9��u�9{��E�9�&D{� �B���B��f
�����6.~����~��j�zJK�bv*�Dȷ� fGO�*�KЫzU�0#��1B�탇5xŢ�BЦ�^�^����N ��ud�,�f��_fy?i�e��G��v1­�������9Yv�4�ک�^�O>w��i�R!`=�iq~݀��8�x�zsV+_^���G�T��ҳ�����Fۇԭ
�z߂ld|���1��4��{�u���5��n����S����M�vs��=q�0֝N�#�:WGX�Y\P�zB�[��f�b��A2����2����M U
�~c�E��"z�W��䶡�be�9[=��J��"-�ty�Νu8boyl�J���ݽ5�]^��}�un�����	�BaVdD�U�Tf	� �Wn�.��l�,>)Ny:;����l�դ2�$(�ʎz� 6��z_��v*b��SGF���Mϋ8�{O�=F'����"�La��y1a������(ŋC�gz��.�LPn�b8sNdDEB�u�yd�z�k$�n%�-8h݁G>�uD(դ��P�Ѹj�<~�mo\ٺb�s�P��TpO9lp���CV󐑚��@͌*��1��i"`�N.`=���꾣��ysF��>:���F�>�<9��lx��m@����f�d�y�\�����2_iAj�K|�����@q��$M=�4� ����<���t�4^�M�knV-Y}�`p�rA�r_+���Q�h�' zD|�^0�����ݡn�C���Q�ǅwa�PfY��p�3`�ͰKP��Ώ W��im���@��A���]�[�}L4>	�U4� ��k�j�V!�G	� UЬ{Ս���<=�ӽ���[^�Z��#��ۜ�u�k!�H��X�C�j���"�דW�E��b�}�L��{df��-�xt ��<=���T;����X������D�#K$N^��꾑��,,v��qy�(F��t
Bu�Awa��=[o=��x��c��9|��3���,��-��4�G���˖��Q���-"�`���S��]�vKU����� GK-ex�+=�^<]C԰c��lǲ]!�i� 9�[��zNiXj��m���]բ�XNҠ5�S�*Ԭ�=γj�ә����l�NٍR�ڲ�r(�/*�A�CRo6�u��a���U_&�5x��z�rP���4]=@R_\b��3�K}.�wUmY�wD�@�tFX�� WJ���A'h9vS�K |+P"�U��ʢ���zK2f�̅����i�,t�1�$�T�{�P
���;�7���0�y˗E�n������NA��֔\/�s])� �.�&,��Ѽ�3B��a���d ���w�A��l��Vt��X3��H��Rd�w�����GI�^dU���q��t,mr/7T����d�ƫ����sB�t		����r��ݫ߉G2�\�FJxk',�]Ή WV�䖐�B#Ki��:���Ӻhw^Ӛ����UԾ���2��l��qJu;���M}�U�����kX�0�Ml&��Ns)PX�b��7�����{����I9+k��*�	[��M�����ڤEv�PY�}�-AC1\qh}i!^V��U�L쥀dÏ��q�1J�T�௅�iu����i�� $#52I0�g�^��T
�S�դ������B���PK]��$�ͮm�]�J��-���u
ʴ����[bݵ/+n�#u�F@�f���wjk�7�ry������Ѩ�Ey��'Fյ7s��:���!�sf�N��*R8�<�WvN�n�܂����t@7K��C.c�mN��̮B�i|�m��mc*�Pm4�^("�[�7ö�v	��:�͚'P���≺��R@�������+���3���Uk�{1N�$9�3��v�j K����/x�ð���a�ٹ�y��+��8zI�
n�`o�T��B�\�X��1엳�bW�Ec��Ǳ]9�m�5�5��r���J]2k��w�+��u� :��Hy�PY�(E��M�
"\��f�.���SNs�h�|⏰����P���Z�ݡ����btC��}��9�Ɲ��Z�� �ݚ�#ۆ��ȽZ� e�jo�O�ug�>�{X��&&��@��*��Qgm�շ;8��ݪ\��_v��G�X��]/��u�v����X޸i�W'�1��}O�2��x�2d�5�6U�:�X�ڐW ���ŗ`�Q�I�%%���d�[�ᰴ�[�+u�y"��HY�V6Q���f�5\��rN�)�deH(c�=�t�Sr0�!>�%�K�g'�1�Z�l����N�3��an:���.��M�-ȧ��.�6s�ϖNF�,>�G��2��E���4]���@�7dV@F��.���1��5W��h���;��.�먩"����&�`!H�� ����GȚ)�mѢ�*h�˦"��]���yD�݂��1�vOv#�4lf�c� �+mw.�I���<{�`|�o����*�n�y�E��тi�.a,}g?_�oi�)��(�h�.UG}jJ�����>�.%7S�9b �[1�Fk��>3���oa]Gȋ��kml[EG9ǑG3���\�5np�Z���O����?��X�Eld�"bb)Ӯ��0\Ω����#O�?_�oo6یrֈ�73C��ѠձCQh�Qmj���=�=����u���-��y�r�A�	��y�q�Z���Hs�j�������᱀ų���m1��r4��
9�G,h��=����ݭT�Q�>XngE<�+�M��s�:��F������~�sGU�����%��m�E�sVےrw2�E�b6u�l�*b����ߟ7���5��盁�G<�qD�H}])��݂��7G�u9+F�u�������&��ԓTW5��#E���Pۚ�_w^��QZ77[���+�aVe@� &P	�Y�I�BaQ̨?q�5>�GŐ ���g�����b�}��_@-W��/�s�q#��2K�YbzܚN�G7�������!N>��C��\1"���0 �P=-�=k,�A�{�G�n,�䞮 �g!!�ԅ��k7S?mI֬Hյ�Nͷ_q���{�����*]��GM�.h���BsJ2kn=�U��3��D�b���E'Ƽ��z:��#�by�O��+3����Ȁb5���کŽ��6����6!(��Dkb�s��z*-��i�r�j��?3���;:�f�M�sv��Ú`�Dc.�*e��̉imuKU��(ܶ8�Z#'�3f�;���j��ڻ,��B�4��(�����P�!ɣ.2$���^�ew{��f7b�LA�U�E9S�y|��L�G��4z �����~/��Cj�)��N͙n�5Unǭ�T�զ��`��s����[�a�30�Z��L��{RRӷ�G$M�q���BB�/^��c�#wkwK3���]H?mR��Q�D�fh�y�Xga?[h��L�r,#�X}v�딥�~�N��E��L�,�*E8-M��;�M_wn?ǆ�q�ѡ��%*Fz�0פ�Yz7��`���U���f��r삇0��v쏯$�#:��u��*��*��r��[W֦��n�e��S�Ā���md�/z^0/~���޽��~�O� 3
3(3
�@,�,ȩ�_��}�������s���� ���b�0W����\�%ff��LؿP:3'c�Cw�כ_��K�G���*$�>C��j�2��R�Aώ�a�%[P��g�Q���T���Z�(]��R�w�Pxt<�Ę~{jDK�#�rFg����y�����C�S��D{��F�{�q�I���MU�у��k�J^� 5�oX���niz��oB�b��Y�d�QxnH��+��9�?c�>�R&���p����C[���K��(	�l�uof��i�I/�$wC.�9���؋t
������3#{��Q���3�e��s�Gѽ����]�r�p���o�j�1,�d3��[|�q٩p`���������w>"�o��A���Ld1[�>�|:�O�����Na��Y���=�	`V�Y�l7�r0]�>a*��t��nE�hqc�-*�'-wt�6�+~ѝX)���{�:�&<��N�"~�l�}k0��m�DE��$v���8�J���]{����wP�0l|:D'ؤBӛL<S�3b��������ǖ��ܶ�Tx��ED7�,M��f��A��]C�b�i۹��&r��cq�v�c��jۅ��M4*�N�����%,G	�*��N�{����W*�KJd��G-.9��Nz��X]f��-$z�U�ո3_<�\�)�pɜɚ{:U�5�Ŏ*�`���<�s � 3"3 ���/}�{������W�������[ߕ�a+�vD:w�D(�ڽ+�3�Uݪ�#��Z5���e���c�U,;���O��xgQ���O�`n�f� �,>7��R�����5û�c�GMx����:ۦRq�Զ�kX	&)���Q�H�e^�Mso�u�F�M��QOd���d91�Um~[G�a�S������~>��<%��M���c�Y�[��I��g���G����^����%���~5T�,K�kޘ�+��"oy���g<_�%��&,���g�3�`������{�����t!�ˉ��Z9���3v_�%]���bg�My�\=w��9�-�*[�)�3����'�Zw�;����L�k��^?u��6�#��a����Jly�S�?W���]F�~T���e�\4áW᜿�G�0����s��^��m�t+,N��PJ��i��#l"�~?C�Ļ����9�f���B�w[��$^��cX��\�2�탹Ch%7�-��;��Ok���a�c�t���'��~|D���)�Z�:�~�]~<*�w�\�`�ﲸ�1V�e����%^�Ux;����v�����4��E�:��ð�q��n��VsT�W&Zm]r# 9�]2����҅	�W fq�h8�m/z����zedRaaBdN�S0)00�}�}��w��|�u~����c�嚶1�N����p~�)�3�J]b��(���7= �F��Uc���d�����E�!�c�u��߾��_S��O`a�e��G�f����ԬHP�ı�\��X��<7�?Sp��i��C�U��=�@��"/&4�opo.C�7<d���Tu�e6�}+ÄLqf���Hb+����㚦�R�=�z�K٥��m��[��H˄+U�wk��q�\�lΫE0��_"��'\Xs	�+�#O��I��?B�/iT*��qga�h�S���T1
�jٷ�ņXA>��Y��f��WW�tND:�u3��������n1R\�Nn������@�R5o8Ɲ��s�N'ܦ�ފ<�PR/�|dB�[5�]�}���f������O.~n�v���{ ϝ����=O[.5�tl�L-��Z�B<���^9�b�5e	º��W�ˑ�����������ʥ����݀�:�*)���Ћ5�Id�������9����Ŝ$��v�������/���`�8�t,ۉj=-mj��r�op�v� i�G��3<{�f�rgj��[�|嫤(���|�7II|i��Q���!{]���
D#̷��\�}ϷS�פ��RxY��Py��(�Xmh:}��g[���T;!6)�Rg������00�0�0��3*�����;����^��^np��p�s�@/�jg����t���lx�Xҵ_$~j���y��~�u9e�ƞU�[�];
�=�k�6w���U����W�5�W{���q䂎�J"�G|-��+����O��4��*��fz��u�O9�EM2�ze�j�4q��h��/^��"�־��+<����s�u�q�P�����e?�c��8�}=�z�X�Y�e���٠��@�}�=�Q�o��0]�Mh�b �-)���<}��Y�7U	���i�g���^���}!���?M��ʒs�r"�sZJ�Nc�=Il2l/f����-OԳ~*v@�ˍ�k����!�Mu�8�g{�����nKu�4ز)��%�cmFq��US](�x��O���2�_d��Qg����:;��5�)ɞ/~1�Z�xnGtu,>�"����l�+$2;n��G����-S��f��(�TE��:��@����GhEx�\�;�-�bg͸��1���w>�=7���x���əM@3�op��5ok��K�0�	�7���`_�&�Ic�q���ۭ���օL���RM�t����3��"wS�>�`��rޖ�!�To�s ����-��o⽿,�%�˃ޔ����q�y*�C����H>������w��# �͐��Ɋl�R�F��2X�ո6Qh�"�A4K�L'p�.w]u��{˿�~y��߻��矱��)2ʳ
̣0����_~���Dކn���(4>�?y�	�%�^y�T����Κj�Ԭvlsb^ƟK��K�ܧ�sw������#�D l�c�>���UB�Z��S�z�G����J}�Y��Ԯz�S���<��s!Ǥ>P�����;��(�Eg�|fu}��L�9�)�2K�����o9��Hd�����I��s��B��P@�ѭ�ɡ�"|��5SS�9E. ���B�὎ͼ�^_�Y#i�s�Bl��,jSi��O���`�p�:zd+ݝ?k�;��길[���O�7���`]gJ23�~�ݔE��2�\���[�����yϫ}�$EY����w��I^]h
/�.Xl�~m�_�zX��(b�f�)ץ���3���mT��en���"/T����ӵ�Io=� �lJ@�ԤD���O��=Zo]��!������n"�Ԓʓ}��H���i��P9���zz$�
N`�AJ��A"'F���ޭ�[-êQ�C�w=��I��Ȧ��Sx�a)Ҍz�=�n�5��o4xX=7�a#��
�s7�æo��?�Y�:䋘��JV'�)5���6^�~�;ySR��*;Xҽ>o�ro�TuQ+3�E8�8��oo�j�bU�\�]F��� ��Xw��rcz>$�9�X��ح\�'[�����J�4wUܓj<��zߴC��2ʳ"�o�x��ږ!Ь7_�1��I���&����^.N��{^�V�Z��=	,6}T�Qt�Ӡ)��sc&������y\��,{ ]�ɴ3����t�����nE��q���˗ؤ��r�[��쌒�V�L,�v���R����,#R6�r���}�{�;�����OhRM�1��+���?�Hw�e���E����\���d��\�;�jP�ݘ1J�!6�l;�Oi����	�H��"�T\~tDC�R%F��ef������VՇu;�NLw���Jg/V�}u�g�G���Ҹ�
�J���O��U0�o�u&�]}{�?B���.PS���sې-�lٍ�%j�A�$M0U�VwX�\P��Ϸ�9ȳt�Ġ���ǒ�45���ذLm�?�ff��2�D��+Yݎ���ם^�ͼU8��K�]���ly���=�O�/�k�3�w�d�UIm�2	x��]j��x��eZ�P�\�œ\�� ��őaã��(/�R1^w�	�I���׿+b����%�m}}�hܣuAȻ�K�s��W��2[vO\�A���_�{��o���,It���
����k�]����-�)l�-���	V`�|�өd��*�&���|w+�����w���#��ckh#�=-�w}����/<�ﯼ?j��RdI�f�aI�fUz���}����|��=�@A?���ڏB������!�#Z�Ʃj���p��m��B��p�z�?�W_��������`�k���Kty�o�Է�3�d7��%T�O
}�GL��{�.� �Dw��[�6�������{�&�/��� WT6�7��^��?�"�\9�V[��x:�Ҧ�}.��:�چ�&<��)?X[�ᵅVk���i�L^K��v��D[aR��2;4���~���+����Ic�l���'�9�)?|Ǹ���z���c��l�l��UGaq-v�HI�eqe�;:�٨����	s]
E��S���,�{��x;�y�h��F�����ּg70ש���Մ�s���&t��'i"�W0ɬ��\��������W7I��5�PR�GC,��6�&� 
�M7�ŗ��ƞ���90%������J8������ds��3	��������(�y�ƕ�Gto�ؕ�MT��~��k_%�U�]���L��r<�Q��b���\!��"U�?;n�g� �Pj�O�+���+��
ŝj�b�'��?� �׮�9��߸�ѭ�)�5�Ws=_8�f|�Gj�U�2'_b�/�d�
�}8r���z���;�lÔ�1h�P%fpN^��Rh9R	��o�"�m��Ȭ�g�]ެ@��܅DO�hc*��Q�2�L�[/�V�?j��Q�e	�f�f�I�z�������������-��&�=�'�3�X�d���n��n%�*����c�u��뼰/�}w�o����y���|�&$��dzD|³�=x�dtQ�n�t�}z����kk��W\�k� ݣ��h��C����ϫ��	1�Xv�TG�����G�(�����s����s�n��W�^!�x������b���ki���{��F��.-���R4��7R���l����'�3.Ȯu�|��Su���($�X��_�/ܓ	�X
c�*��rD0�F�W[r����nz�@v�����B�	i#T۸y�7N�G�a�y�~>��͋�,׻��X��Y�س�*�@ֺ�%L����+Ì��E]
��mBۗ�kð�y˅t�b���ڡ)<���x��~"��g��F>�C��6ݽ_,Ĳ�	V7�UT^��n�-ɩ�;' �p��Bk���G>UH�:ԙ�^�`�`O\������qo��}8�S�b�!߷��6塩 M�0�~�bG���-���`z~�=j~�����k�v�=�׸hĜ��U��sN�;1����roeG�/�\f��֯'(l��Qގ���i����G�ת�_߰�����7����;n�JR��8@��E0g9`moQ�������I��/G���h�ױ::9���_�#0�)0�!2� @8 ��Z������J}o�i�>N�ĵ��k�k�%ŵ��*]���>7�������J^�l߭n�GV.��2y�2�����yO�S�a	J����#��`+���{\>�:���eZ19�Y���L�NF�]g9F�O'��9�Y����sh/>��xH<6eV�g9�A�����J�5����ԉm�]Tݎ(�Tsyy��`�&�1mk�*&6z�]�:�"�'�ɋ��D�?lf�\.,�`u�&�ϫc
훴P�c�nf<P���c5���$6��7�,���R!g|�����(����<'�F���da>�U^��k%B$ZD�Z^H��j���Le0��e��n���;�:��'����>���6ҩ�=8�Ӫ{L�u
Z�L\�8�Z�Daz����>�S'��'�m�	�L��si��;b����N���K�?Dc�b�Y^�nj����i��?��\���+1���Q������;V�Q����3$��HM?�N���<|�c.vQ����Y�L � �i����Z�vrN�;)��l��а]-!V�/��a��![��T�k8�ߦ�`5��W���hr6�&����1D���������77���f����(���Pݨ�t�Ve
���h�@�������ӗ�����:����\�L�Z��B�_%s���w��.kU�H�^N��ō���|w�9us���\Q۶<8Pӣ
�*��'�nVr�`e�|ɍbum�u���Yu�$�P�RDtg8�^�:7h���0�ɝc�ޮ�;%{<�^Me7�k%�[��޷�4;sd�CL��).k_m�C2�C����R.�b��7ŚH��wsn���J�:���xek�K����Ѿ�#��g���AY�0ܭܜ�*=t��E�kkuK�\H�Բ�r�a��wZ�i2����;�o�e��u�l2=e��[]�����p�t��M�K��+����<ο.W�b��1u���)I^���84�u8��`#B�=���ۨ��(��l�s6�u4�c;�@��]̽����hϋ �=�(�尋t9�1i��c8��TT�4H�y���׋�	,����z��%L�î��cw{5<~+�"<�o{]�Z��v.��]ZѼx��Ֆ�(��S.�WY�{')���5�v�Ƹ�}n����}J�u�A��:۬�d"�$o):pV����Pv��"AH�z��`�E�K�B�.�Jo3W8��ʔ�[����&�U�>�|�Ҏ+]Դ4�q��G���k��/bv���#�-����X�y
�-n!םn�$:֬r�`�=�xRכ��m���ro,��O�D�aI�'H��k�</yM=�L�aCRnٷ;2��:���`үnj��l�)��Ihj�tyń��c�ksUNG��^����_s�8�2����i��Z@�\����:UZ91�+��5�Ӂ�M�ǻR� �'oL=TS
��N��54��HX�3��&��3��{�{�/4����X� ��[�-(U�1R��c9n8p�}�Х}[z�bppup\�uS��c��}f=�(�w�[ٮ�� ˊ��t�nN�&�Ӈo�MҒ�5�{!��ܫyu��2,��1��,����]:��lR�T�$z�S`|��hκ߆�u�mҷX;r+���D.�ݘW�'W&D,��@0e������I��&�]��!v9pz��M1ׂ]k�C���[����`3!�kz�	�uYE�����l�
��.�1wE�9ҒzVN�� 8�5�Ai�e�  ���M�|�vT�gK����ԧ;*�+v�/}ena��iJ�0Rۥ��W=�He����q򓝕>� O�Գd��X��ps��\�gE`Ʊ�1��[mDA]�9:�ѰgT;Y'���|{{i�͛cF�O���5�;b��V���1�����ܫ��<��U�����{
��_.I�f����	N[�5Mb��r�b�778���oOooǰ����9�r4ru@W$�ɶ3%;#m�rq�����Ƿ����������6�.�ѷw�b�4j���5Tm�뜹�����ꞟ�׷��]����PQ�m��ËA��5�.G#�s��AN�Ɗ堮\��'�?_����|�(삍ܵ��.�79�;󮗪������+�Y0�y�8�u�Ϗ��ǵ��}�?ql�6��[V�.�F��]m�1͹\�r9���$�G'9�E��g������cc]ڍ��ۑ�V�Gp�㢢F�F<����֎���c�Ǝ�9���c����|�&���.u�����4S�LU͸kF�4�1�b�1����1\�֬���X��m�-���9�<p-<�5�3��)�yC0���RA�o!oq�R�J��b��{x��[){�w���鄘Y����`	������y�ß7��ߪ�ן��u�!�4�.>/Bj=T��n����/<T�2y��c��%����fꉘ�8׼l���Λq�R�)kŮ�??@��/TZ��w�]	�t��U��g�CAj�nn�s-�\��:�V��[]�X��YL��q˵9J'/cЖ�/�]:cp�~��CS8�9d���'����G��}��V�n|����R|f�JA�܋���y�*z�;�t
���G����Uӌ(1��^�P���m�SL5�Q��������������<�&p�� ���/��礿d_�]�g͑?H�c�~V�̬ԍ|����kn��ӕ�\�Gx�?W�.�[��h8@�xg�y�wK���T+�9���)�9o�;�Y@�ɴ��~v�mkܻ,Pـ��h�g1��/\si�j��A�c�Y�u����k��72t�"�Qb�rR����85#$�	P'��^+�!ή�I��y�E����ye��v�y�!�y�=[ާ��j�\� �[?� =���!�iP5��0���U�ϯ����nC��"�S���5��q��4��F0���	����B�7ak����li=E����8��-�w�����M'���{��Y���%��tΰHP�J��j�5sz�����t&������dfVb���e&���HIB�#�zO"9ԃ�n�)��H�F}�\�6c��%j�D-"k0��Z���5�UXR��V�3Ls|����R1����%򝽼g�m�.+�lK��eq�����.�s3o/�My���a�~j'�"�0)���D����D��s�mz��7��5;��A��7,�Mq;s��q:���M�+��J(�LQ5�7��w�LQ|�A|�Z,W�}xX���Ck�%M�uX��2�	��^&�`͏5��?��H�/fD���/X⚅�ӴB���T����'#I?w�Q��fc�oPFv�<��}hkJ����Cy�K�-|�G#Ӈ[�a��op�F�t�Z�Վ����j@��7#{�&���A��������]^%'��!;�Y�����k�\����p��[Wl&\�^S�ynP�T�8���0�ua��tiU�^'n��m�5�Q�W�\C�`OE3w"q��^*|�[B���rg���z�=�ͪ_�)������I	0��|b�"H���Lh9Y�'�������<���Ȯ��E���9�C��f,���4��=e�\��f��v�L/�P�ӅhD����)[�"Mk�xR���+���#CE��aB�:���Yͻ}4����uI���K"Y�=�9���:����$�aj����<wV�1�YI�w\�V�t}$8��hD���*�>l2I�S��C!3I0	2��^5���[�,��
B�H"OQ�[�-���]��u�C�K&Z�/��*<gu�d���R���-�n�Qx��8_Li�U�c��<5��ԁ\�@�C3�hq�S�i���]Ԙ��e�(�COH�0e��\��Fg��O��¹I���W�B�g����l�7�-��R���	ON��NlTx��hU{�ڬӋ�lbz*;�e�%��j<�g��Ʈ�f�-G��g�`��\0o�x�X^}�b ��ye1��7�QT0���CF'Cٙ��-�[oan<�{T��k��P�o�w��b��o{�m�B /�x��f�����3^l�����7�MU��0��J?I��2.�6z�0M�A�<R�`@x�T�E�Έ�*V�*�����ۙ7z���r]3Y�c45:qKh����K%��v����Z5P�9N���-�r���[��r!��v�F��&���Y'v遂�x�:�K����@I���E�,oqOum*��]����p��̋ʀ��E4�\��drtk���AH��K�$l�ߐʖˍ7J�_>�/��+���s;���Sx���S2Y�ԭ���/p�`h���%�^�i�2yC�.`��]����j�uS�{��7k[d��S���K�gZ��wfv��]OQ����wkYu�K����_>s���[�o|�w�9�>�����	��I�`��	�}�����>���|�V����H��֩pZf����R��tׄ��&Ԧy_x����>���U��b��}���I
P@��F�;��w�Կ�'�U[jv/%��+:��&��\������?��߳%C����`�X�E�SW��sG������$v/{��a��K�=�r]x�M���u��8N��ŏSW�){0=!�ǭM,�}��f\R-wv��c���^5�*�7��7���&�{�~4ִ,���w��ܯ/�H��r�����p��^��z s]�ѭ�+>��#�:��#���y��N�sd��#��.��`T������T1y���&��y�^����I�*#�u�čǠ�ni�F�"ɪ���7{:�������B����Cf��Q?	9]�=�b�;�W>���(cF!{=���yÀ��[�@LY����C���Ŗ||�"_�E�Gi�R�`ЗTM]��S\�9J|�0	oN4�ld?����u���� ���5��<�
���wiY3ܮi{����w���H殝F�w8#�f	���<Bʋ�e�%��Wۆʥ:%��1c���L�19�Hkgv�E��#�59�O4$��s�� ����keLu���ș��h��n�e`n�޼��w�L��334��sjI��
o�t��2���v܎���e�
Vd`F�H�e�фKU��O1�ژ�.�2�d|1pN"~��K�YV�#V��g��r��r��Ak�(���(��L��U9RT���5����x"�ܖÉ��͆s+ۧ$n��>�[lqi��)l�����ģ'�<��Uw��arJO$�}R�L�Z|���z��.�OʻY:9B��al�v��D�e�a��ݼ%6����+B���X�}k�͚d@�FЦ�FA�MTS�#���,S������1���2�IW��L�/�\Z���"#<�J���g��`����+���4/4��h�L�j�BRM���!�����鶊��6VP��!᧜2��ms�7!�����sf,�T�;SVr��v����W�d,�	���ؤ����Sx��tZB=M�/�!�ei0f�ٽn�.���62�]��kь/t�ޕ+^ʄ����j���#���������مu�d����y�|_�E����Nldj�k��S�A�%�>aR5����)N�7ΠÖ=�k`�n�9j��D�R��C�,RA��`�av�dKӇ��Y�-~����?S>�io�k%JT�V�'v�I������t���FV�7��Q◥ �u�ҝ�ݭ�ét�\٢S�'e�-���O�{��|�}�?����D�30A�L$�u����~��]Ͻzy���9{������:�)E�K��5�]��7�F���.rα�[yJ�����Z��7ͥ�}�������񖅤ڢ(�]P2a>��������@��;���[96���^;^T<�bYL�0;aw�|�J:{������pph�#��&���:!r�U
5}�k�	ǈ]GS�^iA�s^Ҥ]�����R=���1�}��_`'����`1�	��=O7I�v%-�&eE=2��PǤ�����t���%�1�Z���[<LS�j�`���NM$�pfku��y�]_)�=�|
��05�F0����?�b�A.� Fc���ȼn�q]zn�t�z�`�Z�ሚ�L�r��֩���y��Y/�?@�#b�AS�v��fgo�k�ea����oHFU��~�-�Of��X���x�9{���a��ݪ7c��\��¸n�ZY�/���f�D���:���ؾ9�>j1@^�?�S�M����<�#;������ P̄@bm�֤f���gMXΊIo9h_�T�:��2M��XNьE�m��DRW�/t3E%�f�|�#KN�~��.gi�sr}V�Q"Pa�b�&s*AK�2�
)�9ڪ]�\����>���vX��
I�v�6��I�޶��v����>*oouG�	̠^��(iÌ�w����#�+&�u��jt[KёD�E!�[A�ERk�Y�lL�0IL~l�?{���#��J"�D�4C7������Ϩ��ox�1��0�h��Y~�X�d�<����r���ô�J��\!ܹ� �q�.����42��&�Y��Y���C����T����܁D[6�ն��Μ��h���p�d/>=�|[�$��[�oXOP�uL����%^�C�{a�D��+��Q��m��W�+���Q����|�J^�he�z~�40�9עƗ$OKV�Mu���f螥��(���~*=���a�7���@�yi��e�c϶钧�eI��:�T��\�Ѷ��2XI5'|�_f*Sm�yQn��[�� k��)�"��4��I&��������7X7k�����3��߱�֘Iw��=����y?!��d�ը�W1�WL1�Wd�q��n�O3<7HG;՞���bT(��.(�:w�Os��*�T��ao�����R�b}߶q��z�S�*��XA/�ϱLC�S
�S�����G=GY��p���i���ox_�+��.�D�	�-f�P���2����}x��F>�q����0rGߴ`J�������l�'VR�Z�l��P{�CMYwU�-�+jm�"�6v��_5*s_Gy�3���"�9�pl*�?�&;�ߚ|.���U�R��=3�8�B�n�3����m�7N�OL�B뻸r�n�����n�y����	��f�`�<L��<Y��߃�g���f�,�`��4m5��Z�<���}�ȑHf��Wb�v*ljE��S#s!6ߺ�7S�_�7��c~7�l#T�J,�����:�!n?nZ��̡0�c�z�����;Fdry���Bj��0O�x(?u|)�?������%� �۝�2��toVnB��Ę/C�o4Kڸ��>�O�T�c�0�9Bk�&���6}!/B"��2bň݌��]�~�g�������I�*a ��ű���
�%�*�&��.���b��gu��4}���4՘Kǂ^>0lx�B��3|��k
�n�b�4Tܫ{S=r^�(������6�C�kϔ���)���9�.��;Q��7������[�H�8��f�QjLi��/1t�R��2[w8�2/alSaU6�Qy0(^:���3�1�B &Z��>z�jʺ�:�+g�BoL�1X�]0��Jn�*���M��3p��\[L���=�4��ׅsv�L�C\��A��(UfHSϵgE��ݙ�ZhZ�Q�J�G0��#�f���ƍn~%w4�\�-���jy��ě����Gr�u+M����Nu�).f��@Â��h1]�����]Uo�U�7\��t{Y+�Om=�Vn��68�@��SC^k|m�1l�)�OQ�y]G�9�0m����|*��`�Re����:���U�oE`���O���Fbٵɞ���oV�y �Z��b9������������/��0{�T�<a�]hl�xD||o �ٺ��7�G��#�L��>���V|j�̎V"�f�-Cg\!��O��b T�@E\�P(�+�њ�b�0��[\���=��k.�����7�s�>��3r,���#�4n>lQa^@P��0�֥1VW6'n��M�q~���"ɘ �٫�~bL��uU�I��n9�s�d���2�T}���ŝ���I��)�y�ͨ��亥G���>�cu�~�j ���ʠ��E��k7^��(&zz;f��ɮ'��E��3RC��-sS�O��}#o�m�ZFJn\Gk�K�z7e?<�v�K�>��P{�?<W��Gs~��k�v����^�6�Mb��7�,��b��2�9'6K�.��}攌D�Bb-@^bL|�����PE���>�U�jǳ˻�!ϵɹ�҂UL��8Ķj�v��y���	���Xj�]]�V1�S�׍� �+�M��la��#��`y-gu�Q��2�u^�'l��¢��R(�:Q���k�L�����m_(�	O��
��]vw@�[���%��6�����QSE��od��2� �s��a�n��3���P%�
����{��������}����a�&i$`���I�������:�����9�?g�8m�^Ɔ-B�K&�-�no`YdZ����s�F%�����i��#j��իK�J�qK &�����t&\��m9�l	l�Ua}����agk��������s����d^_�a,��^�t ��ra��W5'��;�P0\R����S%�&�
Ul1�*s2tӆ�h��L֒Zj�\���_G�u�c�Y�s焿�{��(���Q�ҟ2�����z.���嵙�O,����g��11�DF��P�0<��s!g1�~W��=�4ʽԹ��fB<�y<x���Lkey#�*n|�,�2TW�<%0:T�\sdTw�u=��ݰ�6��h��)��4i�*&�WF�O����㤑h@���$>w�O-m����*��,�ᰮ߹�+]-�ʋ�8\W4'����z9��5��k��;%�Wh����q(�q��iM!�<㖆	(�1�<��4+�
q���]#�����֢b�ˑ��[c��5���d����n������"e�{6d.2&ώA��%#w���b���e=x�,7|ǀ��_������`A��&/XK� )�C)WD�*���t^�ɋ0�mZk�`݂��6��ָ#\���[ˏ=i7��i���K��Ŷ�8�;L�̹K0��z\uxE��
��å9oNh:{C��5WHc"��K��hq�Ȉ��ˡV�i[��@�ܐ�ԊY�}/�ڎ���¼ݲ/�R��k�]FG<��
��ٌl�h*Ė�W��Pߢ��kӆ�|��1C���E5�u�����u�6b�EY�����)˓Cd�{�̖�J��aU4��2]!!v���ȓ���/�f�m�X�^����G��+��x�Mt�f����f�s�K��q~#_x�ӆ��	ǒҲ<y`�b��FmrG%`��e)&7���W��5ǅؼg�q{nn�@H-d��Q<+�K��9�����Ы�((z�U��!�oE�u{y�s}VCkW�-�5y�p���[�p�Rg�c)Z6𩢹<f����wb`�nbT.-hW���;9%�狨qa�#YJ1_(���X�J�v6qA�ڄ$&^t31=�� L����)u�m �*�-1Ei�-�Vॎ_w��ô�ۜ�ZﲥH���Ĺc㮉�O��-"�^[�+7�u�=��J�G:k��(.R����ruv���ԑ}t�Ծ��N_0+��|���$�u���ꚞ�KK%��t�T��R&Hά��wp�K!k9�멹3�ȹ\�`+��S(Eq�M��SghESm/�{�w�
��ۣ�c�@1ZR ���n�vGL�GN�[�&�p��4���$����+�,Y)�nd�►ޣ"�t�җ/����4-=��Im�B�h��f�Pe�8�43�	����/�1�Q3v��W.b��@Z��\շ�)*��Bp�!�Y�7]�>��ht�Tܽ�q���}Qu��bW�gͺ}�r��p�V�4��7���j��s��KQ�µH��`g;�[�v�F-�4�0-���:�%����mt��i�+��6,*�A�EH)�P^�̈́r<��xō>���P��D�LP�Z:z?-���0Zv�@&[�'Z�}�Ϥ����Y��8&sL2�nuSܧJ�*��:�c*����� �9B7�m�Q�Qe]Y����9�w&�	r��n����Ƭ՞ 4H��o#W��S������k��\#X��Z,����k:���vJi��L�3�=�q�Fݳh�7��ws���B�)�oxڄK�:MY[��u����~X�p�p���PQ0�N359@�f�q��竧w7Gǟ��t�uq�Mε(�f6ԧt����c����uKH���Y�g<A�y�`�h�4^�ze�Hr����u��V�� 1đ��L��7k��q�>�]��e1nͥ�GDv9���)��x�5��){Z:��Ť��,n[{����r�	ޝtKgs�v7\+\�l"$��6�:��ڥM�;����i����-�T�I�EHrq�T�!L �ѧM%M�>�͔�M��藛r<�T\�Ƣ�m�j�np�[,s���V��m�� ��t:lj��-4T���������IM����'9��Ŭ�5FƣQ��n�p�j��������v!ѯ#\�ڱ��M�N�5A�M���^۝c�ιm�85���%�������ܚ5��5Z�:
�1�1F-Uc`�S\�ˁU]:�h������{H���>󆨪�P�Vu[�������A{���tF�5���O.<|||{{�j�CZ`��kb��Z���}�Ϸ�Du�U��9���nm�ѝ�.X'����oa�=��}���b�r9�r5W9Ɠ�槕\��,s>ܹm�X:|||~=����~q��j����clh5TѪ1��E��N� �;c<~�_�om�u�f��&�|�O �PRh�Z����RPV ӌX4g�m��(6�Jl`�*�6�b��#�N�b-|���宺�l|6�߾�ŃqY��U�9iN�/�@�k3r=@�":K��N��A�*��Q]�%����=4��IE��<�Hh�X�W5�?�?L3�A3,3�0=tE��w������ל>�y9�����n�����*R)|P6�s����P�'�#�;�ٸ�AyQ�i��&�.��E��p!����iީ-A�Y\��P~F�Bb�U��Dy���^�_B2}Y�z��
������/�G�o�T�x�[�x�ސc���]#���Q{�T��t����A6*���w�J������[�6L㍸j�Mp�9Bh"[(_G�Q�hcJ����Y0����.$l���zoj3џ�?|�t[� ,&O�%��)ռ��#K���~U"n�jp+[e��jk9e���������סu���d�|
�_@X��-�z��O�����<�î�]d�^�V��e�חc6_G���DG���%��Ց'��g8�C��ER�n�dt��R���з�%�{m��<FDtR�� ��Ǡ/�(S�����g�"�������_�}P4�l���T�cqe5�����r�I�;qpMխ���=��㽾�}�J����ǭH���?M�C�N�D�WG+��9յ����ʧ�t�n/��J�ӣ�ͱ�8�R��r��|7"��@q֬V�z�~�M\/jǱQ�Փ����()2�lݫQQ��K����6�N�6aZ�I���L�l�t�1ݩ����+������憖-��s��;u�ϯ������2� ���|3��7�f�5R>,V��z�������Y�V�]^=�������'�����@L24�M{�������	�6�05�z��}|����dˊ�}8F��=�/g�2@�U"���w�2q����]�6F��ɪmM�e8wt^����
�K�j�b�|~Gs�*ҷ��ȏzf��B:Z&�*�B2A:Vi �+yGР��ӟo7�V�ǸZ��q�^P�j��N�^9"_u�UA³�� j �Bb�Y�|�"Vo��.��L���A��{��3��)(f�3�n�Jvff��9>�ީh�k�@�
�A�^ ��.0������>=��~���*�/�Ug���;���krL�Y!����(C��'G�9�nՈ���@��C�S�SH�a{��S�V|/"8���
ޏw\���Xڵ�G��͔�'MB�j��a�t7��5n�l
3���5�<�xWr��x܌�S�Ϳy:��A�jyO�ppg�"-�f�85�L约�2�绢�5�8�d&�F�)Lh.�`76W]������7�/��O�ܼ<�ӽ��>�lf3��l}�����s�Q�w(�C'��y6�.F��5��T븃�E̚"�J�MwB�_&!@��7t�����V��&�7��͟V�|���F�;�S�ʏ}Kj�3��Ι���l�ɫ;k��Ew-�����̌����}|�<���W7�y�~�����%�;��I�����(��&m��
[�3�<ۓؠ%� 	���%��8�7b���B���O�\�!�XW�Ae�
�d���6QWX¼T^L
���&��y�ʨbm'�Ǜ��T�TW�:�#8R�O�a�����;s�tÌ�m�8���͉��-�<���.ǝj�į�j�=�n��\��:��B���k@��:es�f{V�����}ϼ��P����ХJ�ykz.*sr��B(���y��,}��fcY�L�	��_;��!���;Ȩ�mQP�Y�_��u�>�j�.߇(�&uO�l\�����{���l߮e��X��)�����X"2�ծ9�p8���V��}н��e�@XG��͏���� %*�c}Q��
"���^�~גw�;��IOW��1>�ŭ���nHs��Zq�7'b�d�����U�ۃ��<�WM�1����܂v��z�����v�n��0�\�wMx�W��b.6��.�u�(��d'.l�Y���ك:4��/6C恉j�s��Xb����T�\���7v��-���g2*�Q�����gbA��g'p�44Aj<��<يI���#�O�R? Oƅk�v�ܱ�!�kyЈq���|�X�v�Q9�W1�Ǿ�@ˁ+���#��HӇ2���|/��Ɓ\�W��|�|(�m��ҷ�5_�q���持 "U��f���g�����UCo@!�㦞ھ�k��-��;�^3��Ђ��ɽp{n��&S�ڇ�|D��[�����$��&r���=q��}��H+���y\�����D�Ȫ��U�ӻ5/�3tJ�Ku�L^)eʝ��}�ǘ���J�JS�6_4}���k_��Q��^��ڲ��J�b�|@R����oN"��\>�T^��s[�dM0F�V{�\����rh'U�Y2�i+F��c"���O6�N�]_��_
U�Z[��V@)�t�f�i���Iy�VLl�T.&�І3����a���[��<�Z/9�nJ2�)U*�/�j9s>�ѹY9�9��$Nc���u��{Ϝ��7�&�C"�D枼�8��=}xy�]~�����C��"~\2���+7�*��3Zd+�䏬F����]$c�=x����4�;�Lcz�)R��pi�r�hR����l��J�W3i#�f��@���QV �)��Kx���m���juz뢴��k���IJ���\\ݡ��KZ��G��\��*��x&��"����Sw����H��Ecrc�[��7�Go/>�������nr���S m��ԷȢu _����a�^թj�Q4!��KTGurN
��e���N�gL���la�T����El��������=�ۼ�y�X>j�v�5�k)6��n�Z0�hA�e�@����W��";y�w���1��G�]�;`W[�jF�JU�ic�G<�y�qn���K�k�e|{�_�7X@t�=�T��ʷp���$���sd񎋘��[�<������ƟwP�3�������Mf!�Y�|���,�*d�]�Wd�n���ok 3;��)�>	SB �N�Sj�<l �[�,t��(�=S]��t��˞���^��M�y�6?rʷa��������i����	I���\�Me0m`�3)��fL/s�0B��Y�R�jʣ{�O*��ՠg�wUMeK��S`L��]\�(��>�J�e��D��^���b�QZ����vg,���{otX�Yv�ר}�Yi�v��ǳ+D���C���=ڐ�E��/���zC-O���wX�hg7�b�v���PE�v���st�N�(��u"��s�id�y1vo<֪���Ϲ�.vx2������=槈�����uC3��wHk�V������@�����=OM���yۢ��r(���SV��Ϫ�Ե�����Y��l��.j^��e�qg��=��sL������al�ЃW�#�u鄴�fK��sؽ`XzVc���u4@��5�ќT��<l����r|�G����~�{�[�m+���aJza���|�����*9;�m�t�8��J6�H�7�M�D���g���u"o)�<�˨	�b�����qݵ���/�z�6b�^��~����$���H�[��@��x#lVP
���\@`��7`)
=���U��u��96ۺ��a�4C��@��}�A�R ��F%�2�E�P�ՇL�r{���� �����i'qg5`31�����٬��;oH(f^��Ǚx1��;jͤ�[=Z�N���4KHz�s'�7��M�ѷt��͟��j��:�M6��Bq�g��x�ٜ�h�y�W�k���Ҷ%T�=����aUa��V%F��eV��4�W��4*��zm�Ɣ��|�TW,�n6u�h\��5�灩�!q�M�mL�if�0�58�3���|��=��0�z#w<�7�"0�UM����r{��T��e2�'����������h�jL���@L$f&���Se�=��-��KX�J�iy�=�\�K2��w)�N���-�eg�x	&�ed�&�jo�����Y�J�����ڹ�F�3��֤=�;�sK�
��E���.��A��E�%grf�1Xє"H��,yd���B̭����Y�An3�a���Ik�VVT�H���S����]�[��v8��R�dV	%��[**�&����iPz(ya�;|�������{
��d��4���1��3f�\����m��O�}A��jݧ�N����K���P�YY��>�x�zy�.��uGD^d���
��5�o	u�69�[�79C�+�7C5�t�|	��;�6��`o���$�����"�	���eO�\	Wo~��i�v�c������P�Ka�m�J䉤��v���}�۳�T��ۅW7��r2����WX2��zڈ�$t���*��Su{s�Gc���Q�.�[{zΞ�������{����zsu1w���t�w���g��Ĝ���ZR~\�ĭNސ�.c8�lI˯��٩d}ձx�j(�w/K.Π��\q�"9�����k�<�ӽ{g�S(sʹ��=ȯ R:�����bq	����n�x�7;�5���/�G[/�#ė�l5�8��f�VnbY�`�7>Fqw.ґ���Ɂ�cx������@ҷ�_b��qe�\T>�d^�����١#Caqv����w!+2����I�V��-'�����cn���N��H{�9Οn;�)���dGZ˖l�[dif�c�`�#y�IV��t`�iИ(W9m��_��O�<�\Y�9�6�ﴻlG��[���C$9�zw�y�M|w����v��(O��uۭ�soր�P.\_*�w�><eT�rJ�=j��Sja9n��A]�J�`��y��6��?N�����Է=xh���r�y3ύ�&�2��q�-*��*�Y\:���L������.��:Grf�Y�o�p�� 5o*������g�d����e���ww �3�Pu�#���ooBհ瀽֚&�s5p(RvN�SM9�2��t��"����W8�g�_+Lު�u�\�u��Z<-�<�D�J		�@�Є������6(���M�ۿQ��$�*��M�f��t���v>�T��iq�����udGwG�%���dk^lB�����Wg�!4�y0��U^[N3��q��S��^��w�t �	e�ָ��{N*�Js�n��E�љ�򮆺K���$nC�s>���Z@�C�'nD�'<]�We��	�h��^q�&�㌎�����?p���H$[�#Թ����m@=O/D#����;��ܟ�2�J̳�DK���q���ɭ�dZ�}n^C���1ݐe���7���Բ�=
�Z�7Wu����ҜS�
�}�ۚ�����4uy�؝¾�Gql{��U��➚v���q���cY��x��Җ4��	G��9}>��
\"�)��<Tq�bxOAM��[Z�[	���/ڭ�XC�Sﭨx�οbޞ��^���v�&`p*[��W;�F��v)���Q*j��`]��ҁ��
uv��w.��� ��q��N[V��O(t��7_U)�X�#����|�Ve�ŭ��w Z;:0w��Ң����{�3����kjNی����Q��F��)�n������������PiԍM��yO
0�+��޾ؾ���=�HXP��^���^u!�ܧ5S7)r����uJʭ��,�M<]��]=�]?DFגW^�^p�(�+d�w���l3J�Q��5.%������3�7�d�fe����dLv��L�QG��ۣ��m�N,\�{�k�Γf��o�������&����P-h�NZ�����j5�̱��%�ٸ�Z�Sߪ��lEg,�:Z6C��9~�+z�,����Re�]��}�kL��%l�x%�x��q�4��!���X�)�tY���	f]|�4��ǽfRz�~֐��P��6^.V\��gWF�6hȍ,�w��*WoP�P)(xzz�wg�bN��<LD�f��Hy�ڄ:��`�Y�!��d�;vў�c�޳������Fu �:Nf~A���.���(u+;�eLPm9���(�hVs��m�`�<yY�M���Xj
�;K�oz���m֭A��Ym��,b���/0J{�^�k���Ʋ�u�������{�_;�����R��=^�\�ʈ8�޶j�دol���U��V�t����,�+{~w!)ND��n��6hIs�GqR�N���:ҡ$���B�+��a"�fw*3�\��
sY��eugYw �wM��;"	�[�I5VwvP�8b���Q�HG�o�He��l��4���L����]����]{vZyez([έ�X�a�t���b7���=����r��O���S,�0$���3��s�4o��
��Z(�"޸��h���m\���HSm0N��ɸ
��̈Zw\V�#ݯP]JR�3e:��%i��nCW�+#޽;tEk=�!������h�yH���vCA�]�ht3Af��}pU�`�vp@d�(�e�]��4��z�/L�J��y&�%�\��[��I�V�=}�bt�9ܐ�C)����-�)�Y@N��+x�0��j��X��f�Pz��	�X�L��[�Nua�V!Y$]5�(�{}�>����(*�K�wȰ2E�;��]�F�O9�¹��;;�{z�@��@x���)TĽ]t�B���Z�n��e�ҷ����y4�7X�o��«OcU�o[�5��\��5��D��v�T����x�Cg}��V�N��5#ɒ\��7���nT
a�D�>L�N����l�Q�^�G_ڻ�1ڶ W�n��z��u���9z�&�'�U�KX(gvu-dn�N}�3ݰ\%�^2h���s�b�[����G��'�7ϧwi���(-�X[t�}Ս_{9�f֌��A�D�.I@�>t��VAӬ�hO��#�%%�Үbŏu�*�A�PHk+�<P4oX�\k�]�t���6�2�ދ<�ڹ��$�Sw�v�+c,���d�rqaeU�j�}ёɵ]�}�ۄm� ��,��ψ.��*�U���Ó�4����(b=���R�'C��6j�Ԫح�X��d������X�S:j��|���V���ET��V�ʺ<q
����RYT�����sGJ��Mva�W��oV*Z1��w"�d���q*WE�Fv�R����ZΡu��.醃��o���L�S^ڌ��<JGW�Ry���C�\��ԟA�݃��oS��g+k�U�r�ެΥ�.���QP���۔��*�T��TJ��+;$:WVv�5Cٔۥv'r��k�����C��vHE	6v��.k�Ňw�w�뢫y���Ugc�ᒜ�5!�6;����4�&�b�T�p.��]��9u�Yك�3O,n&��k�N�u:PųG=�����󻫝r����~�N�޵� ����4k��<m��i6Ɏ��I�����{�tZ�w���:�:6y�K�:#�j8�05��p�Ѱgg��������N���yD��j-&٢�Z�jq}���5�������:pq��~���p�ch�V��:��f��ۜEDmE�>�p4���ӣ���S���Ƿ����j6�.s�9�Y��V�I\��r0<�9����:�g�oooǶ�������#Vt:h��]m�h���5|ƈ�u�X�":w6t��s�����6��������kO�EɵV�V�F�s'�d�r�*&��Y�p8����{N��w$�E6�Dӳ��IJ��ʱ\1�9�����<�������c��M{r���8j��n��F��&���α�tE�ι��6M%���ዝ����r#�Z�����-8�6�4i�,O8a�7c�=^ ���$�
C�'�f����+��M\�g�����x���k�������0��&�T�@鷣l	ڻt���k���z��}����|x{�;_����7 >m�Zg���X�I/b*��d#3	;����o"O� I�:'��v�b}� }�~�n-�L�u��T)yL�'�^hM�����1Ks����U=�a��mo6�qώ�T�{~�I�����ѽs�xF����f/�1����ս��|�׿P�S��\ܞ��L�+���^aNp2���5ɇ��M�����t���$"�#�&@���k�2֯Suwdw�غ�{'�jdAJ.���o���ek����5�jt�3
��wT˼;$f�,z���&t'L��W�"���:�ƴ�s���f���1|5ȢWu�e��PՍ������o�v9U�U�+�]����t��K��,(n���k�^�x���n��]`�%W�gz����\�6�wXsOf��Ò	����ɾSK�ȧ�txq_��+ �FP��N�gPbԫ��f���S쵹���O�1�3�5�{Z�,P٣��;��Ƶ�˓f��V�=/}�X�����졽ZF.�Psp>ڗ�����ֱ�Q��'�r�:އq����B+B�Ϻ��c�<=2p�\
i���W��,��cm��WQT��N+�1�<^� Y�����~ꘃ��C[Ɩn/ժ�� Է��/���}�^��Lxz~��2����ɟJ!�.�ٞ���P/%0�����@��6ϱ�	[�79C�)L��S8����^^a���^ѽ9e*�6ZD��k6>o8��[L/KV3L�U�����Ѥ )����]P+�e�)�] ��>�����;�!��ɢӘ�gO�"geG�0M H:VU����O9�/�ť�������r;�Ԗ�뼟��~�> 9��	/��M�,�����=tu�N@��{5 �)�4��k�����ݩ_�P�G ّy�21lxs���Y�=��e��5�#����[���"�]��C��ψ�Ѭ<G���������f�晍ˊhYD�C��.��oQo1�W�ؤ<d�x�%�	������%�����pͲ�*�Fm:e�-���yg���(S �r鉖	o�Y]{l�z�Y/6������ѕ���(Y�oY�ji�{EA�=��'X�-����.^��u���Ӑ7����S�ӥZsz�T�<��u��ݩ���Y_QI0"�	���-ݤ?l�Pםk�ы�d��KҺ
�t������Y�:z��w(�^vW�UsK7 
��e
��8��*e>�n�:Z̽|���y��G7v�f�1�Kz��t�9J��hI`���ʹ¿K���9r(L�y��O�30��[�N�]�����-��^K&���8�s�`Ds�k7)R�QVx�h�n���5lSX�%_=���3�4�gz�?t�w��at�Ff��.�����//����\�!l���ʳ6ᮦ$�zN����Է���~+ *�ʎ��|0
��}i=F��ܲ��6oL��p׭���ܓ�|�j�z�� ���d���麎A�Y���Q���w�fv�v��%�ڨ��d\m����5r���M�(�'$v33�H;�MMFE�&; u���}~E�B]+����Լ[o2?�>�߿T��IH�Wrfڑ��MOK�y!��>d9�*z���jN���p�G#J�n�/��q��"��d���c1�w�=�N�%���𔤯��}�k�LJ	Ww�v���vQ���7#�8�7N;=��"�8�s���� ��rm�����K<f�ѯ��!3���ۥ�K`���c�#̃�6���J�KF�ҫI՚C'ֶ�����%�����ثϥl�����/�PM����+9�=���t�NE^���n���?mTq{n�VI�2�6��i�8���� 4�����/gU����O᷷�m���q���0�*�Km �\EC�)�ݕ���g[P��s�(D�D�G��͓�����*>c]�D�tǯS#.�]+k̝<7zC�������k�5:�S�5[4`���y٤
��#��껛I.,���?��nVإ����ĥ�[cH] R܏M���ٝ����>�g��`�UB�`q�!��+*:1�M�c�2q��M���os��Z'�oOu V�{iÈn�H��|�p6��F>���Ne�����mo/Gs��3�R&���S[��G1��!T:�i��K��A�o�w��~1pƮf��b&I$.��:�-�szl����k����H����D��u]��}�~Ż���S�^�<̓�;�Pj}�ݨ}�N衔�ZiӜ{Z�K������7zȃ_٫��Cu,�5����+��3��#;�>'%��Q��;���f�V�Vr���3��r����r������u8�.�N(�����s������h$�*�=3E�y7��|�0��Y�.��-Z�P(k# �����.�D�R�Q:���[�ާ��DVY��F�r^1jG6`���mfJ}�9l]��okjު0��ٴb�/vf��If���y�ὬW��񫏕f�!;imW脮�P�~�v��;��Zy��]�q2E����杨��b!��c�5cI�K�}6����N�`��\MEF�G����T差�\\�31YA�F�� ;�ͥ�P1B|����B��ƿP1o��x~��?E};0.���~����l��l����_��a��U\v�6+3dߵs������������uT]n�`_z���m�����'ͼ����d���m�{���J�f���S?��I�z�7����C.W� |&C��Ү���r5��&F�'Z�ј�������˟|�Δ�;47%�_f���^��ER���i}�c�1��6�or�-I�w`I���J$�$��s��m�{����Z�����Y���ͦ/1J���k`'L�g��<ȉ�هp��U��;Aw:W�s8dn���U{��62m�hJ���N��o��Z0����~V����S��q����mm{�7�C�?*��O�Rފ��r���vU�m����&�ҜWyE�������,�<��K���|m��A��f�C�=X���#���䊕�T�iMS�fn�!�`|���F̞��b�ߚ5g畫ן��,ud�Q<ݛ��c[�o6n��w!f�vު�G�{	,�Z�?[���p�[�!�|'����L%.�?S���^DvUt9=�-�_N׺2�}G��va�� 7��'���i��=~�в:�XgԖ.=��'zB.F�͗�^e�� �!�F�oq	�a-2�\T�jΛԮ�IM$r��KG�����跾M��-zu쮱(od���A�d�P�o����$���(��=�K;�n�E�>���Ц�ϳh*��Y9R6*34v�u�D�Q�t� [̾�}Ա��s!%�M���}��E*�;4�rr��O��WO1���|��(��G��`�4��ԍ�TBt$_�{�T���Ҝ�L9%"���Y��}��u�e�yg�4u�L㸃8��$�Y9w�
��z����gC��:kW��	8�fQ��Fn�N����^�}[���9���z�l2��g3���s�(��a0�w������s7m_i.�hv�oN����t'Cإ�0���~�!����y39���l"�,��w�@qCwO����/:W@�ͪH���n����AWY����{��?I-T�(�Ȭ ��C$1s�T�y[�������i��ۻk8e�s�ږ�V<��y��*�@�em U�P����������t����j��=<��A���O:��uy-����]Z�Qʐ��3�*4����ﺀ`��ẹͶB���5v�4W	W׋����5��> kx<�Y��إ]�|I�95��-�s|wjXp�=�o� :{,<��+)�+ȷop��Z�_����b3�m>ʴն�!���X3g]d���$)jv��x�55!����+y{�k�� ���7�N�.����C���a�:���B�gN;�"ɝ2wH%>!�Wr'+��b�p���W�5k�=�v�o�;�&�y[�9l��`mz;����lR>b;��P�]�{�C���y�DK!@9��5*=�{M��\�W�v�{�e:�'���jL��b�]a�"�`�H��*/o�+�-Wq�V~����''9_v�{϶L��y�}��~��[I;�9���Z�_:�h�ޚ�$]��7S�s�����e�ŸR��M<�1Fc�<��|���U�ɭ�۝��z�kukx�b��&Z}�;�`8�e�͊<�WW$�<C��#J���f�GK��`����R���l�4�`!H�ïg %�aF�s����8�I�-��>�}S��i��cH��ͶΟ={Av�5i��׮��>�� Dϭ(�.�</NN��Z�R�j�N����c���uw�;9��Я��'lj#0�v	�� n�w�-4��g�Hgr�h���a�ҥ&�XnVe�� �ټg�n�7���"Rc-�C�ǖr�#��P�,��]y�i��<f���$���#K���+�5c=�F�x�x�b��78�k�v��fu��jl�Wڞu��!vr7�/�Y�H:��<�\�;=0^׽�S�4x��نd0�Ǳ��%�@djW�`<�n��ꚷk���0�[g�ϝnwh����j�۾t�d5�y�x3ꤔds ����aw{��Ӧ�T���u�2���	�gԱ����>uY�FZ�j��^�1,Z��M,���5{/��6F�%%��k'Ԫ�����e��̗.�w?о��~y��z�삘���U�y��!�i�Gk��<�L���&V��5q~��[Y����8x�4���eG�TK_%�t�畴�)�P�89[�u�D]Op}���ٸ+Z[���d(�B3��>+y��;e]�nʹ�[�ٷ�����k�uz`;�h	�/7O�L�Ӧif'������Ӓ������[c��,�F!:Fn��m�`��7�a����Ǒ�4�6��,sf�r+o�����#y\ �07<�W����w��q	��й�Jy_a�[25��������Ll�'Wc�Be�i&)��m��<��C̺ w���zpbt�U�����`�
�뛓�v^�դs�݆ON�9�t0��%Oa��Q��4%9��N�R�C�\��K��|��d���W�5)�ʇ�WK�73�v�q�30��8�a�}��f���-���<��6���� 5]z}z`SbҜ��YZ��ݫ�U�����=*}VwOS�V;?H`�k���n� 1T�X��g��OC�T��tl:1'ox���4�4�@Ͷ��Cl3���T��×��c���Ud�l�W�nm}PЂ\6x�ǱS4��pg����Y�8��~<��l+�e����{3�9�":�М�`衼��j�΢* U%;�;{��b3�K{��6��魬�e��H��j��[��3Gei���ҍa�v1l�ڨ���;a5E��v��8U~��� au����F��d\{�o&j�^�3L���1N��ۧ�� 6t�z�+�m����z�g�������k6�t��V]Q��k�9g��\������������Lmff�s��A	E�(J�3��f�3�k���]g_��ov��D( �cCV
y�����Gk(Kl8En�
�n�Ӕ���s��	x.�ȱ*)��%���>\�p��Ҷ�����r�!Zl��*:��}�Ğ��«}�KD-�q4�����t1.�>�sg;��w����A��^^v��N�#��9�ZsS4U\����k@)p{N�A|�k��h#�K�������\��C�� v�g��j��}����IH�сa�Q�,�=\N�X��O �=[%�u�t@a�2kgF�|t����"مc�8����9֋S�)��HZ˱���i�rq����o�v���R��u7���Q�p����=]V�e�3�F��ej�M���o��/��;��\�����9�:k��-1Wj	l���psh���1SG�|ݛk��f�}L�h�N��N� Ul����TʺܓA�Z����cIɎ�Df�2�ssQT�[ e�u�B6�����O8�K#-j�90���i�͖��v_(?���.�\��ij���Է�1qsI�����{��^��h$�ьm�,�'I��[�u�#�7��^M�6�t2�1�|��2���7u]f=��W�V�_����j��:Mc����![w�53tͦZǉ� �]7���vT��2f)�Q�Vri���x�FԷ��n_M[�n��&:3G-�֛LD8݆�Zɋ�WR��S���)�{kbT�$���tإ��dAJ��#8U'�F�&��0�e�wv���͢E��5\�M햐��[��[@ຣ���RW�E��n�}�U�f�1�u��ɍۗ�z�u�WB�WJ�|����P��j u�6�A�20�	O^]	9Z5j!���ͼ�+Q��Ʌ��P��z����D�Z<��F��}�p]��SG����Ci��MGZzZ�t����XŬ&M�m$����*w�J덣��T�Lp�,���<4��"�N�`�ɂ�6�\�0��P���N�Or����Pэt�9���[D�ٖ�����ɲ �=�X�ع������ѡ6+v��]m�{���V��5�����N*�{�h�tܶ|�U��@쨝wF2���c���zHQ�ǹÐ�<�$(C8;����&��0b�e���ɰSsZ'p���w�k������M]�Ys(�|t���y����Ӵ'�������'1�ޮ�Q��̡���Em�7�P���X����1���4�wL��lH��`�e �Cv�|����U��>��	4�WY��Z��t;��u�]��T̜p�ˡԀZ��ަUA<Z� ZYev��s}Ηk��s�v0C"l�A�m�|��:#!��ː!��w�0.f�i�y�ea�È��gj����r�z\�)Dz3�)	0��F�W�Xb��*tS-V.���R�S~�C,�<�-�m��$�t	j�:��4S�*�J�
:���W�>mu�ˮ��uw|��q���C�m|ቛ�ꪣ��m�"�6����lYζ�k�h�G6��UY���?�����jc6�[Vݜ9����������b9r��sb�s��x����{j�ک�f�j�o˜�Rh֏�"��\9��DDA�rӢ���s;������;�F����\��g�Fv�H�wUAGw\�����Q����Sbہ����ۻ:���6�"�nU�4�#�m|���ܚ�kr�s�+l���n<����.��:�m���ncQx����w�r�E��\���ǎ&#��͌i5UsnL��UUDs�y���\�ߟ.tث_7.9���{{{��v�ڻ���uָ��]W,r��j��� ��\�DW���
�9������:�4�Bi֊*�s�Z�������|�wnZ("䛑�&������p�4��nsh��C��h��Lr�?����w������h8���{{���sr����\�5��X�l�Lu}�|�8�`�DE���r�ι���\�utsu�rNlu�3���>�.��*ۻm�Z�lu�����rqW ��Q�V�QPEh��c���b
��o��.��M���;Tמu����I��>��\ ��9���+�y��b�)� ��z����f��!�{�0U�u ���w`�C'tZ	2��-�UR��:�WX[磻�'��Ǳ#Z����e��p��
w���G
�j�qh��H�)z	r��ƇF\���6�#����w%��a��~��Z�<�fc{��L�ȍ��\������B.u6kh�q{�%�I̼�����Т�LB[@L�q�4µ,�}������--{�SV�da�2×��w�w�a������~��)�涣d���Ǘ�r���yƝ�\7�zR*�t�������+a�\.���',{r4���Y�I��՝����gbyz��:�c�L��t�"���m�"(%p�aߩ����{[���]F��:;�M��������]:`ba�G��Y%��:�/�N���5�}?vF���U��w2�e��G�S�gC�N���i>�����m��~_�t��Tw�����o�z�!���S_��Ȁ����bZ�"�slf�{QYN�����KC(�Il�;�Z�9���B��rt�T��˃��7{&:ٖ���[W]m���:��y�2,=���.\w���eZ��]���"��x0o:%9��3�j;iF,��W�5��菷���-<�\7t�)�վ�P�D��ĺ>�urm>�ޱ8���/7Az~��4ۼQ�p��ۣj���Z�u���/i񄦳E�|{MG�~�ܒJ��W��BƜ�u%���� W�q�L�^.]�W�xJ>��!���o'&��*��;�'���
�D�n�ڴk��yh�ݮ�G=dF��"��0��z�B�����O���Q�v�񳱮|	��*���EMZ[=|��Ҹ�r�s�=��j��S��r�26y��u��'�����<%YX�=co�$_RH�#�3��Υu�z=gң3�{=��+į""�pm��Hț�@�-��P�T��eQ�V���YD�m��:���iԢ��gٿf��vo 47�#>��h�>};�f1qgmFUn�;n*��x��N9��������)|li����˟i=K�nN�����ƶq�k��<�p��8p�N�J<�?շӸ\b�pI-�:��%}�����E�*�]���94����n<y#Z�1���֊�G0g=���,����i�5	�|!N-��ͥ�	\A6)����B�f9T�P|vs�#��/#�5՚NL��9Cbv�#kB�=ʴ�^���UQ�w��t8���!#���/{6�ta;�gC�-w�r7��Ĥ�ý�^�N�$�Yc>���������Di�ֳ��՞#��0Z��jxe��ȍ.�G&ΐ4Z���J���g��9�9DO����~�xz�����j9��l�$$�a�����
F3��L/L'��1�K���D��2�nq{X��'z=��s���l����M��Y9�_.�?M(�R�e��u��o#x�F��}��/#��q��4���Mg�<�YO�Y�$?k��bTV=��M�{��ݔ���~����7a,�)kU����sȫiS���Զ�oq��o��o�|�4]���L��K�ك-�-<G'�7Ue�;��,&�� ��]K[�U��<N'�Z0�>�ŋ��*�C6����s���.hU����^����=�r�O?�].�=h!Z�����M���hj��E���]�27�*;�;`V�kЎ����y�����J;v����o[O��IÔ74\�V�܁�B^�0vm���(L���=g��=,��������niuC����=�g�r�e{�z��5X1������/q=<�s�b�^����K���uQ>���ݽ`D�J��ŭ;x�Z:�C3=m_Wt*8�x� ލ��w�$>��i̓wʪ��T�䪷�W��;DUi�1Qبo�
�6ҳ)�o���xncݢTRs�;ٖ<�Z���@�5�:�����=�;Ӄ3	���O���s<���蟟���B�Nekf@��8ۍ��Xi���z���N���-z��p����dd�ߵHm���n&��NxFb��K��ܝga:��/M>�\���YV�0�e��y��	4lNd>���3瞚U57��,�� �2�W]��#Ij�8�7��|z�t6��z�sT�]9�4]��V��St����![�"�Y���Uu[����>:{Ȭ�\A�\�^�m��:7�]�����H��X�
�" !4��vu��P�U��y�N��3��7Ee�@���ݞ���HGڨ�]�� ����������-�+����1ȡ@�<�����Y��Ro��ja�]/�T�	�u�0���4V��#�Ǒf�j�YtVBE���3"� �<m��h����(��L�wtW���;�0��8���&�;��[Φe\�޾,��e�#̪����	X�X9S�ԕ�R�dWmDn�l=��k��a���i�[��|�GQxe�u�O�Wm����Q�z�LF:Z[SC�Ud�lzl���}�K��fn^�AM�(��/�����؃��vqtzC4���3Y��������<�VWl�%}Bs����0e���_y�����^����G<Y��#��rW.O�hs咫��{�!��]6T��K��ÙiJ#C���ʔ�f����=Z�����x?E���8�f��3�Xk))����z|�B��>�ڰ_k.y�﷽6�ފh�9�^�J�(��`U�2M�3fE�l9z��	��m�n�m��M!�KI*m=��[^�!i��y~��Yٙ��ӡ?J����ھY��}r�.��@�f��"����{�q�6*Z;��)[ӄ\�S ��Sx;Em�[gY���H���f"�g�=*SRh��\��
X��4���ݯx�_��S|+��3f-w�S��E[��%��ѧ�`Z�J��~��8=���i������<k�g�3�'�z��4�#�<��u�U�X�.�wz��SV{}c4�czz�=h�Rt��*��VM�ޟ����\Q���|W��I\}���;�Ҥ�f�8&�|F!�#b��-wy�YϚT��	��"_�d�Wl�qW�;�-H�F:qS $��2mB������<�]��d�藥Ws�/����8��[��6y�``�;�]�oM=m���ӓ>ͷx�ǅ݆5�&|�@��9а��b��k|��U�8g'����W��}ݺ{z���)c@�e�֚�r��-ކ��"��i1����|�ZIʼ)wW�U�[��̍���g����O�U#Qw�� ^!�p�9m���^V킲uG�����m�NS�@y�Q�Ty�F���>�
��}�"�N�.6]g�=�����|O5n�b�=<N��0.$�w}Ֆ�9I�f��]'�l���@Ǔ�PОY�|)�U��(bC�_��3;;����2p�#�!����wSO�vU�H��&��XN���I�t��K������Y���O�ꖹ��u{���ݥ�q�A�Է C���^EVGG�Z�y�7	��b�0ɉx�%�^�eQ-���Bwʸn����j}L���et�5B_�"��x/B���l˫:CΊ�mCIW@���"�Fg8`����jʿ�r�KQ�~貘Y^]�M���&�z�����˅ͳ`e�{�X`��bpjf"z���^b2v���#x3��F�R3@�Y�����I~�u����_�m����K$�{:Z�W\�@b^�tR1�siq����	�5�O`B��r<����Y�ݷ�{��1�ڰ"n8���Se�f�0����߳��'|74��.N�[��>�}B09�����&w�3����/��\S�헉�r�_mU��#��A�r�ަlh��>�����tq�����]YX��r�&���h��ך��57���,w�m��h����:��3�ޤ]����s5��t��zM�}�7)Fy��:��B��s4/(ej[�OF��Y����t�j�D(�ւ��>Ϗf�ӧ�)N���:���`(�Ξ��Gw���fd�R�w�+������j;�֍�^�fe��s���^�|y�U�^Ev8�����U���&�j�v�^��0��Zn+�z4�v$0��������>M�V�H�W>F�ݱ�lue`1;pr��b�;�Yb�q���
�"�ql]�_�L���WP8X��8�n��yl»w�gd�"��O����z%�
S�Px��%��sLR�1��/h�$ڨ)�ϻV��f9oVo�ϭT����(�鈺��|�����Q�?tZ�%�/������3�L��UM�;vIе^����x]�)�j�01	�#:<����7�B��ҭ;,�e�W��)�0�l��V�(��~��������B�L��wk��;���N�j���aS�}�r�,�������v�V�U�?��E�,����Oq4P>���+�_lϠ+;>l������j5�i�VU�덻BW���<�Q��%��J�!7[Yְ��1�֝��w8�Cb�PZ���e����s룸LS+�=l��l�ҙ��Ԁf�A٪�뙫;��*�ѕ�vWw)-S֗m����2z�m�Y-E]�v��=�����ձȠ8����8$�SL����^��M��;��m^}����m�k���`&��a������j�tN�ӗYy�ͽ]����5��I��m��6�jr���~�nm�ή�׷5��י{��c�:�3���6�-x���S)�l2�AZ���sy׼K�L�S��b��	�����GEo��=	N�\��������Us�b���֒���YM���FQ6��̠�Z�v,���GS����PUϝ)ea���^�K��\��;[���4p���n^�A+���l��Dr]b�qTug�S���}���ssxtOWrAj�NyM�UW��o��<��S@~$V�����^9�֛�gh:�⃽����:��j���&���==mf ���}�xOE�(�Sʣӡ2H��-`�B�l��ǹ�g�vfoe׸��,�j�G>=�m܂6 3si,��#�u�b^�]��k�*ohT|K�7��.��+�p�=��������}_-���T{\-ޱ�uY��V:�4�z)�,�?g^�V�lF���f."P^�^bn�٦�F�n�a��Q��t{=1�@)������>+u]�ÊB/,���1�L��7}�k�\��ޏ:%�R�3��Ι��_k%���6_�ܦY���o�,��0X�|s�dX�(�m�*<�ru��y<�����ܷ�껎�sk�l��=+��<�W�d0�i="1р��%�6gv_��r�(�d>t�Ϩ�5�G�cM@�4߬MzÙ�j2���3���}ݼ������ί-my��X�W�ܳ�X�<�e;�C���`IPm���:wl�;�N�h��A#���q���-(�g��ܳ�f��Y%[4r�@)��3-4�yB�40TV��:b���/U9ꭲ��^�/%p���c%�΍ꭌ5o�^_Բ^�� �>~��=��)��7���w�R��B�{s�b�{ښ���J;&�I�{����o�ݍ��7�t|��&�K����Ǻ�~�[������.].C�\�i�L��QbSifo$*��$V��9��wF\ƮQ�u��[e]�c���֎����Yc$���f1�Փ&p,GA�C�S�b\ɮ��62��qRf�L��+��r|�t_ӄ�Fe��)�F%)Ѿ|��N�������$|�͑Kz볚|e�ç�=u�AP��Ǽ�PT�u���x�R�)�J�a��Z�@�!qw\�����e&�
�=�c�8HUү��T�PB��CV�c\�д��p��\�4�ҕ���Wmk�|WQЕ끣IoR��ή�Yי{�J9�\�4�f��d2ų}��}�ey��a{������K��]��PiSnmu��^l�5oW>M!Y�Q���V�3��{�[�;��\�.�1A�,v���}�dVZ������:fBsGs��2�G�[r��
�G+/��c�eќdm�Lb���Z��s�WRݪ�4n]
�sIn��������t��c I=�*u��&�Z�l����R��fF�Yd����[�ڤ��1\�MPypfоd%��y�*�۷7�.Y�����X7X�6���� G7lt)�!�#27;�����&�� s����xv�[,K��,Y�y�.��zj�(�	�e�ܮ�PNAN�w��^�^�SK����]�,�A17�vy�N\�6rT���ː�ƝM�)y��tۑ)�y��Th+ȍ�Lm׆GVh�wB��)�UX9��T����[F� ���
�: �G�\���E"����Yc)$ �[�o����JZr���h�ٲ�=S�|���1�E�OB�M�\���4\�/}�o7Ե�.��%`[]��{�Q�i7E�[Gc3J���+����6=�.WXy�_�8Mr��tu���a��u��Z����t���n�"�n�{�!�݀u4_v5"d���Ժ�#�_v��R�4ށZew�B�m��'n9&��9E!J�n�"-�����}�'�oM�m��O�۲D�IȪjќ��ź/r���4�����Is~�f��ENZۻ�H���h[NK�$2�u�t�`�gY!��F�h����頜���ys�D�J���%7�}�� V��d;����
ur�w/;O9����ۥ��x#m>��a���@��L�\Cߥr�	O��yӥ�v��svr�2��h�c]�zs�rdb*�MZUx�t�Y�v��T��N��D4k���m�Y+��1$Uz:V.�ӛH ȳd��2��r��[}W�5ʉށ�aA��@n� r=�|<�N
�����n�-��-�A;{B���Q��§aZ����螮jt��SwP&SJ�r;������,+�*��1�\^f坖-�p>���7o�ɧ�N��cΗ�,�;`��1�{��^??>�����b���Ѡ ����n%p&�ֹ��h�<�I�3������~V��Qƚb���1�G'��R[��5|�8V���a�Mb#��9q�������hwx���*	�8u��'ݒ�ۄPQ͈#g�m��������r����x��{{N���8�h�b9h�--ZL|��u�F�)�\��˓F�*"z�9�\�l��Wv�z��:�m}��=�?_�]�(���#�S�ѭ��sum�9X�lT�u�㣫Aͭ�luͶ�7mLN��*y�m´�8������q��DQR����0]cE]cc�ss�.cQE7'P�͂��uclu�q������_1��k��*�(���mU�{�<�ኃ����G"�6ڈs������Gg�7��Y�Fۖ-<�F�����p�uͬ�9j���͛��LQZ:�b���rx������ՋDc��
�����v�;�91���u���T��[�]Z��#�ܵ�sq�j*����ͭ�k��A��s�61�ULQX�F**���k�nQ��Pm2Ch�o�;'+}S6�{�~{}��
��&����)c7}9����(KM���J�ϑ���0�<�Z�J���.+C�����4�J�������U�Y��d����
�Z{M[�Ɉ��zl�����[�â�����{��
����w-�^���O��2�'�g�u���oơ(��Κ��|dZ��ᭂ�,��y�<���YUՕJ�[\�6����|99�B�F�~��@��w�F�ޮr����ᘌ#{T
���{O�&��	��H�Pdߏv4���^�]��*�e(���]O�\�S�ۺ5�0�ʾ�cM���\�"r��f 1����0[�肍N=����ez.�rt�Y0�g��i-��;�C�'�"�Gz�� <m�G�<��'�M�UZW�l���,G�B����n�����%t��揵@q��Y�^�7�
OtOm������	�I)���w�3{	�4d���\Ok&iηa[�����CRu�����
G���~�JU߯�Y���F'�T���bi%�Mr�!ҭlb/΍F%E��F�L�2Ej������ʬ�.9�nW'E�(��3�Z�sIx�Y�}'�z�,kZmE�=u�'K�G#��A����8�ק;u��}9d�<��C�N�I���f{�-�/��|�`Z�z&�P3.گy�}��4d����\#�Pj��;����z���.�!؛V��k�e/T՜���
U1E߫\��eX+�u[�qB��D��Ą�|p��Oy�٣U<k2�1U>f����U��Z�^���l���Z�����S�0��؀�~��U�tZ�$Qujn��ј*����v}No'��Zr�Uu^s�ʆ�:R+c�Ne�J��!��K�.���{��� V�N�W\R�kK��������<xܜ�+}��|9��|�3)��g�
�3�Y�:�h3�i���M�h�nټk8�@��Hq�5���M,�����u-�-ޟk����jL�^�4���������mmI�����+'��a+��~���[j����p��s���:��Ro��b���� ���zA���b��'Y��]~��w����o�l��U^���c�Y��	g�*1Ԇ�Ifiv�n��4��<5��m��P�P=e��y/�RmL�6�]h��o(��K���#����RTl�^h��zR�]\���m�;쳃{�9sq�b+b�z�Q�9��K��.>�"d8̖�#��,fn_� ���3��*g��āGq�_�n���+�k���Uc�U*�M��j�Z�3��+o�S��V��fo*�[|�W%�T������[���r}��r�:�lD�qq�T�����Tv:�����n�yٞ�����	�׃�e����b� ��5��D�5��
��q�VZax�ˋ��ד�rA�}��"�!a���X��0�*���b.U��;��]v#�&�l��:[a�#�}�oSx
���#p�_����g4cǠ�1�S8�I`���M���F+f=,��-�^0U:��!�z�wN�X8�Ӗ} -��otx��U��F�ZUE��mY%z/��p�؝�����&ɞ������\���P����6�ds��X�(�mf���:�z�;�����b�*��Z��J�>���M�[0\Ld���͟�G����0��!���8�F5��me�S3ee����[)�E��%�c�z�R���g���t��Jsrp*�ڿ�}�ѹ��OT�3[�3;B�$�t���;&���Δ��1}�RZ�,@����4���i�\v�}I3cooC/{ӗ�0�$?H���S�M�Q@��ƕ>vf������Z�a��nC/fv�#z;lv+��.�֣��V���1K��L^q�XZ:�#R����32��{���j�~`��ͫ��[V��J�A/Xu����OZ�3{�M�#d��a/��@�3��3��-%�y��%_P<�m��o'��4�n��G�K�ץt����/�)>lT������{������ͽG���X`/�4�>
�M��^}[sR��ǝd�t؜��86�1�'J1��^]��.�g���x`�������~=�_;��\s2�޽Wp�1�L&�s�/�3<})����^�s��vPm���-��F#0�u�2���Nn�����������z���蝐}�l � y#f>�=�k�̒�|v��D����r�`,�V�U\������4��>4�d��^1�'S�V?cți�KJg�f���'_T =Pe��������Լ��A��1c�p(mμ��s�yF���g���6�6{�����������6g��R���z����ft)b�Ri���{u��ri8�����^��x���u����`���p�������J�hc��Q@���4zh�Ԧ|1�Y�v�{��Vģ���rG$1���S���k;�)�����2��n�r�<�U���Θ�J��m-��+)���un�>���L���Wej��.��L����桺%r*��"�deQS^��MK$��M���5�V��Y��㊶�W�V|�73��k��k ���(�<.��;ݐ��cd8��9˥�/�iK��X��]^]��Iݬ5��%Ck)]f��f�����)����\YY^�>F��+v�Y *��n��gӝ��sVǵ���ʅ��C>�e�(i��+�j�~[���V�ek���ALfq~�vݪ�wn|�$���C�5�EM�A�����L��q��me����a3W9�$�?(�+$�3��������'?|����;���ېXpr��w-Юrq�Č�%���#2����c�ҳJ��֩Q�/��c#b�*GI�4��/�-ُ��[N��k�N+����$���|��̽#�o�)���S���r�u�p�������:ʭ�{�y�qԶ��)�-ۭ%��d
��O�[ ��Z��FC�j��f��U���)��I�Kl$N�s��%,{س�*[���P�H��<p�Ϫ.�5�EQؑ%�I�&4!��=�C�r�����;S���|�_���b�GV=���ێt]���&VS��P���dm��s�ilm.���9�xt��	��Uﱛ�
��k�ɀ�����P�ɯ^Rd�~�)tM�^۫-Ň�0��2+���m6�}��iLMuW���w�qҖ���a��*wN��f�[�##�w��d��ړo�2��:~c����M�5t呒�;g�^�S�Q^�� ���b�X�ߣ@}V�l"�VV4I���[�Q�t���fu7p�_*���T^H*���F��}u�d�Fp��	/���F�F	]�>��ÏPTNt�~�t�8�M��_'��ߥ�; �z��{���	�nΊ�k�#�?y*��:x�pW,qz�iR�έ ':7�;Vnm�7�ӗ}�qMF�+u�hr�T���W ���3U����޲nT���,y�X�������]ݩr��Wq�$��Ƕ�������Zo���g��C�$� ��! �G�	�>*L��g4�o��4��̷@���W�B��uBz*?vO���/�Šb:5�F�k��y�l�D�Ȏ���:Vɳ�Pj�z*���එ�['c��ٲ���=��D�#RsW�y[An�N'\��;,��}��\y[�,A�lg���D?C�;t^8�w�:��)6��[$k�g�/����VoU�Yמ�y!�ч�V]�Uȹ�{e>Ӻ��F��;d5�U��=�r[x���i���Zh��h��y��J�+���hT ��B`;����sr�%�q�š����d��"�M�jM���7���֮�6�����؟p�*�8_%#��n's;���"��3�BBɟX��k+p�2��i��8��رN<e�U(q��Z����8ѐƃ@�k,|w$��b�;a�CGs��a��fng�A�%�@J��v�����̌�v7J/���ؚ���ަ�y�G���V޴���(��ss��s�?V �b!�Y���6�=�l��{�.��ω�����˷��[��ԡװ�tf���t�b��0�4�����\�/�^�A9ݨ9v�a{:&�\x[É}�OIƴ<�:�mN�����%� ?zf=ٿo�O_�R�w@Yz�q����HA-V1S4��F�V����t��ʫ�|��0�#�S��⨙�w�����my+��M'�t@�tŕ�y�ǈ>���Yp/hk�s�u��3!9�ڂ�R�ʫxg�t�g4�����32,�_��S��]2��mU�z;��#�O^�-�Q�Նſ&R�뭣��b�����u�r	�F3��s�U�����g�â�m�T������J�ZCtt��R��^й>�m���S.��(��{b��j��9۷�-��E^,C�KF���w�v�-Y��	+�y�.�Q2�:�n���*�s ��W��]u^�"���a��PYz�**��r�]��6�>�����}l\��ob��2z��/��Զ�·��wZt���s#k@�-	����{r�T���õR��y���oLe�Py~�e	�5����1�9
<�Y;-�ԺHt���:�>�3�T<�>6X���7�W�^��7K�Յ����<ܖ����[���ݏ�m0`�-�I�QoM��@b4�����[ڜ0#�P-��S�n:mu��^��WI67�K,�wu��V�ߦ���w\ڇ�O{�44�y�<�^������3rT�nع���集w� �����U��Rqu@q�zr;��3�w���8dj��5S���r�>�ӑ�t��MB����߯;8C�m4 ��1=~��(z��5��JT����\{�%��=Tgja����y>��x�����6�;"��`]}i��v� �mxS3��<�� G���]��$rC;�}%�i[�����蛫��g�Y��{��1��e5���R6Xo�r�fB9W��QuV��Gӥ�6h9w=&�i������3Y�g�V��:@����iM�mF�f�:k��w��+�)���p����I��>�ft�e����>�����U֒�Я��Ftu�Ҳh�4qV�W8Xі�@ >5�r4nfOb�أT�g�u�W��Tg�t$�w"r'�Y^�w] %��@�ָˊh�φ���^T߱�8RĕËV��d}[B2��u�S��[Oj�B��J�l��1֓z���PR���d�U����=kkX�ۭX�Aա��b���{���c�����˖P}�.C:��uͲy�J�<w#8�wWg��i�:��� =p�VG�;��y[��+]�cyx��f��q��b{'_�B*�_��)t��p�빧��]f�WѺH�&��N#8泑x{�����.W���1苼�Y�!�{�и���Q���-�TΥ�G�'���E�6�����N�x��HNX�fs���0�^6��q�U��Jn��ۚ3������>.��ՙttY�}������j2�Z�sk��7tWKDBԨ8v��r�"w��O,�]^}��	�3��+fȷ�����Ҭ�����]4�7�{"�]Cw��ߴ�V����?��/𝛙�ҽ�ǻ�[(_�@g�00����� ������_4��uv��E#�+w�]�Ojߘ���t6��8���Xs�8R���l��
�d��3�����u�n֢	��7��6X���4:��]���������{�H�@PW��������� ����*(���p� >OýЎa�&����` �� Q�  R�Q �C� � � �d"TzݏC��"`D �`��� �a �`@ �e@ �� � � � � ʀ@�D0� Ȁ�! �@0�  @2 �@0 ( JĄ� � !@� 4�+ @2�
 CHA!
�EL��ȀHP2���00�L�2 �0��M+�*�Ȥ4! 0�C)1+(@�H@����(0�Ĭl d!��&E�8�T]�r���;��P|�;���Q�ATaPPf����?Ug�~�3������~�����d�{�|��� ���L���;���__����j� ��A�_����EE�w�� *������聐?�?�/����?܇��W�����O��<Hw����g���q<��?�?�?��o��T $�D $B�
D!��
@) �&	�

P ��
!" R��A�Z )AQ�T�) �P � �T�IQUĈ0 �P �$�0� ��! �C*�#"����B�	)�A ��@0�,J��0�*H�� H$��B� B�"��K$ L�J��(C�	�!
" �"c�����������U @( @)D(��7�����������@�������
�����?��;��O���v��?�:?����
���C����?�}�_� *������?�TU~���; U��?�L������0`��o�|O���?�A�:�V�����o�(�
��>���w���3��__������� �@�8 U���ܢ *� ~������/����X>��������^��x}�_@_��A'ߧ�L����?���>���O�QEQ�������EE��������/���O��(+$�k*�5��F��0
 ��d��Iϗ�f�J
�R�6�٩�*TUJ�E��P� 
�)]�+�Ul5�$C�*DTQd���-��UE"���B@�vu�b���s�R�ՓF�ZKYUc,,X�Y,�
iv�.k�镡kUf�Y����f1�ф�V�*m��6����ivʊ�-�X6���-����gd-0�L6�m�V-�6���4�����l��
��Xə6��mR��aT��0�ml�X��+��ڛKE�l6�k4�[m�oX��U�ʛp  ����:�v���%R�ٞ�㞹ލT�/q�w�:���ޛB������wy�kmKݻ�[zc�<z�m�p���w��;���g��Wv)��+۞����W^�z�-mPJ٢�ں]���iҪ�_   ����aB�
��nć�u�i�(�$+O�z{�"B�����BD���E�o�2��=�]ӽ�vޝ�y����y��v��+j�Y]������j�;�^�Z�m�͝r�w	su��oOY�f��q���d�,�o�  ��}�m�Kl��޶�����{�������y]w�u��yj���ǕR�d���{ҕ��J�n<�{�v�B���w�^ixw%�z�u��{wS;w�y�7��Ul�7�ʦ��K���cV�W�  >����{v=�j���S׫ٮ�Kk��P����u[{�h�x� �����C���y�QZh�mk���G��{�Z���z��.m�����3n����ݕ�l�\�π  s�Ej���Z��^���N�Uu�=����j�����;n�d5[W-ڠ=�^���j)��]U��Aeu���N���%�m��5�m[�M���Y��Xͦ��   �&:����à����m[{�5g�k5U�q�Ӎz+TcЇ�^疸*�7W��Z��g��x���Pk�늡Z�{Ǯ�����Ӯ��H{��d�  o>րj��v���P]�v�U f낀K�ˀ  �s�� �� �k�  is�p  ݸ  �ٳcf�6�eU�v{p�־   �� �v�( ��`  wi�  ,]�  u :�  w'[�Æ� v�` ˛KX�ɦ���ս�uZ�   ��  ʰ  �` Ge��  �a�@ 3�  �uS  n8  9�  �7{W  2u�ֱ��eEvfl-Z`��  �|  ��  �����w �@pàB��p  up  y�  �:p �@���t /|���R�  E=�	)*D� �SR�Pa2 S�A)U4��5<@*H�@	2��T� �j~??���c��_��㋊��[�0c�[&�J�*�Z������xc*i���{�xx{ޮ�����m�����0�1����0co���&m�6?�������o�#�)���?q.ɼ�سbVJvv��x�^& q����7�Rۄ�:�!uk Dl�MjF��4:L��m]4�n�6��m"��)�R�](6n�*m�kh�	���ա�����YݦQ��+2���7c4�9L;�Q=�2^�gea5�
;�4ƕy|o�ؠ8�$&����l+:12�;
Ah�&�-�!N��zE���@Q{�B�Zƈmbae��w`�v�m�"�uk����q]ń��vCxUL��J]����]�٘e7>R�c��)4�bX�YkVGr���I.��e�W��r3L�t́�75�������:�K���,�]ń���I���j�6��� ZM�9�S���P_Pj���(�i��v��:�Y��w$&�1U�]�!b�eER,8,�t�,u�EQP���X�7Ѝ�uy�r*w�:�i5J
y����>�d��t����`E�nY{�����x�ˡ:ۓ�r���H��Y
`0Ʈ|,��/YŒ��Twi�zC��8wY5�M��FͽHa/�r�]cWW��4S��^��і��n��R�#�(,p��aXh��X��겋�>U�Y�(���I�Μ�I9W%S�m�z��6ŵ�����;{yz�K�qU�"a�q4])ydV�[pR���R��`�n�D��y�"��4c�b��N��C0n�.B*ֻ��Sw51"�����ZʬR��cF`�$�S�
�)k�[Z��:(nn��m�ӓ5��+/n�i񡔞���������l9K[YKmD�c����xp�ONE����5��b���ʊ5�+B��r�yMb4Y������,1b͘[�]��Œ��@ݘ�K{���`7�n^�i`��n��h����A�B��$�{��
]�'fU��E �$�һ'E�R�+t�6(1��������f+U�e디�90;u��%�tڣl�¯c���
˫��+q�����x/+"[o��K	Jh�hn��l�Y�'�!��oRRjF�6�u�ɻ������V�f�"��^-ִ��b�9�,�n7+Sv�.Q�w�w8�Bcm����V�2�3L���Y�!�����Cm�*�P��fh�!aU�u�60e��m<u�N����(lK�bv�òk�I�ú��D��9Q|l�:�Ŝ�v�Gp���Ÿ*�R1*ݬ�_)��#�I'�;����1�k$��P-�6�V]��u��*9*[��k;ݳ�W�H�,=�/ �O}��� R�nބ�V��ㅭQ^���4*�z+-I�*�ղP2��V��D,����I��[�̇�L�unL!��K�M:���Ht(�L�(�;wd:u��<9vW�̭��4aB�j�4ta`c�L�8��m�à;�ILոt;�Z�Z�(u��wR��͘`%u,a=P�KU��[��;&���;۽�
ݥ���SP����K�D�v�5��Uj��$��a�t/D&
�)�L�*��R��@�������[� �V�B�Uo��VsuF�0l�q�w�`h*�٢�oo)'ch��T�n�hmQ�}�m����Yl|D��x�.I��%�	Yh*��:�Q.�̗�2\uw�h�V�CX�*�%Rf��Jb�������B��j��M O$׵��)���-Z��W�q</(�6�ͭ�-'�y��@�
I���s�;WV�ی�V�	 [���0�j�vY���6�X�xb�(͔l��C[%��K+#^
BT�Kr"�4+jV1D湷u�$fS�i�}�-8�	�FZl�Gq�72=b�캔LmX�^+�o4,�x��p=��H���tNHĊ�B����H�S@�F�Ґ������退F(����n^�b�.;�6��Z�o5T�]!Khbn�*i-+�W(}o]�3W��N��n�jV�t��ݡ6�����X���U����]]�=X�h#�,��'�T�\��DՏDw��&��R�[����ZXF��	�Z��G��t�B�	��n��P͡0��[B-��j��D��2ط@@Ʊd+,�P��Z6�`3a	�ld 7��^�I��p%hGcbz2Wh^`��h"w�\oV�$����+��(��SƤ�+v�t(}�Y�*MI|��B��ڔ�s3G���i�ޔ�S�����6�(��)IIeͧ0#x �AYj�r�QI��j������OF��fUډ݃B^n�j��3B�D��2pG��x���Y5&bj�[���@�?,���*l���m���� �CM�Bm71-Y���X�RZ2���(�[qC`m,o#�2��L}�c:�K�Ӽ���E�%�9��A-p����i���|Աe-cL�J������p�r�x��Tת�YY7
2f��A+�f$��RRhn��|�wrуN��և��ڹ�i�����j�2�ug+6�e�+�2rP�h�D�ی��t��U��z�'H��"0(����R���q�Ia�EY����C'�TU�\�ض�k-����^��2��iU���kyt"/F%1���AlS��l���R�b�筴�P7��'Q�X41�1	۹iͲ�,on�(�hf�N��F��R�5f�r�{�[n%Q6�4ŭ��J��v����r޺�BY���[�����@�"kZ�o,��-3��Wt��$V�N�A1��@���xB���Y���-݀�,�̵��5������A��W7U���YY#m^|��C��f����4õ��0�:ƙq'�ܢEm�-�@
q���VQ�� N�Zb��zah9FL���5��´v�q�
���t����n4Ɯ��������ٚ��8ҹ���׷���cp��;J�ݺ��l��F5J�F��u�e=��' �1e:ٮ�a�F�d.Pe��l�F���� Mf2��Iͅj�#laG���ǭ��巊�XV�sX�	̵I�T�p��=�Uػh�ܙ�6��D&PWK�N9�1P,Zt��0�/1^q�k���6�)���0]á)�*3�:&F4�B�7Rcq� �=�u6�f=�a,���S��e����M��q�t��$b����4�L�h�T��:�$&c�E^f˳E�ʂ�dh�&�#,��H1TBk�ʍ<s�z�#�zw4i0�#pa�=tt��
WtEe�jf:����T&�&���c/$<��=��`�nJ����AU3Q�r�!t�ċ	�F�m� n�B�4�۴����)�-��4�L�Y��ʲ�锖
��lv��R5�ͭC/*EEK��ZU�*,g!Yz��٧�o4a�8�Xce �,�����Uw�a��r�Sdە��0ZY�V�˺�#����<Y�v��z��H ���C4��dVe�@SXyr�������m��GLmn%$\gfŊY�Z+/#b��%:X�)"�׶��D'�*^a��D)�X[p���Y{�rK�����VJ�Yj���R]$s%�Q뻬J^*�c�όRĔ��Y2��Ѐj��*^��yD���0����\SUJa;�o/^���!�*��HM�F���V��b�,�T�ún,\��$BB�{��OX�QlV�U�i�P)Csr��������q*�v8���	�2�<H*�hS����Ϝa,�#W/�v"�)�v`1�gV��V����k�B�ƞY�X�w&[�jY`.�é]1���6�⑼
��daI�F�6Y f�^兂���E�F^�)鴉z[��>Z&���Z�ĕ�9o4��R��f'c1�t)"r����X�fP)Ǧm�4&7��obs��2ݥqk��G4nU�ce�+4`f�JPjx�ՍʳN�M|�#)n��1+�X�~�"4��/���q+�zN�ɑw��3"7����{�P*��Y���E`.�m,T��k4"Ũ�l���w7�@Z�f�.��H��f��֣CX��M�++T�k�Z����v�hܠ�4�V�:F-U�&|��t�1�KM;"�"(eikz7!)u��Ţ
E곑+��nZ̊a�ۛ#����ٳ�9�C�In��g��}W��܀jB�f�a�ٴpm�r�V]нE@�KM\��Ͱ�1�Y�gK�� �N�Q�XѳO.7�[�C���f��D�GK �f];�f���i- �ܢf���#�I�N�1i�y�5�٩��� �X�vP��%��G�d8���t-�x��D�*�LF�P	��IN�e��ua.�����$�n�q�B=��f�U�פ�w�2�EBa7�p��a�
��Q�7f:F�$�zR��¤7.�ڢ��Y�^�7ȉw&ՕrV<:�J9uiꗑ�Z��J�䗔�o2͗^ba�Sx&q�@v��B��@�`R��gU#�/cw7s`��tNج;�U���e:_n,y����W�1Yp��-��L�nSR`�qQ"���]�����8�Z6��{�un�s��fd�R87bx�6�F$^ͥ�6�zN^��2��Bի�YI��-�PV�É���Bv�+tn}v)���v�J�xel��e�w�sSN݀4d��%����ĘIfAf���lf��X@Tw7++��K����-ap��9(�LYd�pZMYOt���е�6�%j�&,ןff�X*��fS�� ����U.,xHYe�r̤&���z�C�;$"	�5(��E W�#b��6��L�"o2�=j�u��31k����9Q���d��p�R�Ĳ���I���f��e�-Q�KB�[�a���;���Gu�y�
�Vr��0�R���Գ�ߛ��]b�Cq[U�i<Ą˥���,U�_n�����9V �Λ
"��Z]eXdBU��bUq5g����z�7�d�����:f-9bG{H��d��g&5��Ek]�nIE����A����uô)�]Gcb�7U8��]�yc��JS�6�[N���JD�����M7PK��sB_�[9���L�Z���Q�*�M����Gf�O���N�!�4�Jh�&=��1w�+��l	5�Z������n�z���(U겡i��Ȋ��	�ʳ��y��{p��$��ȶ�@�@�{���"��	��@�$�k��X�EZ��.���yG`
���*�8�B7�j�
؉��l��ޭ�H�zŉ
��n�e�j�V�N��j�	�F��ɛ@����oF!��*򌂎�T�;v�Q�w�QL��J�4ltR�fڍlaMe[��&��3�飖�hP��f��SQ*�Ct�T�ASج���f�6��aV:�m,={�p��Z¬YgQGh�չuf�ƴ3b�٢���+D�>�����Q$im��)���0,�ܫN@���"
�j�R���g5�ݱ��,�C;ia��ZȪ��e+2?�V9AF�\�Tb5�hH(l�)�Xv��t0�st�ě�F}x���z�%��� W�l�uy���Xt��D���٤rQT��IXj�ۡYz���m��W��×��-�}��3n��Ym�(��s)���^⻡Bh��G��Ke�mK@Py���@�ł� ����U�KK�9K���F�UV�Ѣ��)"�w��i]6���t��
�i;{����u.�# b��`��8��&�Fe�n��i��1��<W�)�V�k�	S
[Z������k���N�v�ݹ�T�<aʏJ4�^K�/�C�C�/�T�T ߚ5j���ź/wM{��7��j�v�ƍ\�b�<�2���o�&�ٽ��P�]�����K[ƶ��N��%-k��+	R�۠)�uJjФ�+^���e��K9lᕇ��k��e�v�V��� ��3^F� ���&�GZ.����5S-��բYY��ʲR�	�Ȏ5����5��e!j*ܲbĈ�1e@�XV�����o�z�׆mZL
gb�kn�v���ɍ퐷h�lӟJ�0�t��Ԗe)��.�@�e��Ҷ1]����os֙�(V�P�y8:�.� *�j0Q����ʃ#,��(��ݺq��f��qS�)�m�rR��w�a�ijP�3v̰k6����� ��ơ�'��ݧ	�����F�����/rl!���wt�D-���gX�+h]���͕�-T�������
�S��cIj�4�(�"qm�d� )Ԭ�@��Jʄ!3Mi���=��oh$&=!�Ԓ�a���܈/������e�$�#-��Sl�[(R�kc��$���\@�����!&��Zs-Z�a�ى�A�Yּ�VnY�.��RʈLߠ$�:iQ�Æ�<p;�)�K^6h�;;[glZ���Scph��� %Z.�Jއ���]��E;{p[�c����&,&�O�ۭ_e�vk@Qu�C�l���.�z��B�{��b�lP�Б�:8�6���Y�ٍ�3����:Q�uǫ��r�U]����+%�V��ׯm�� P* �D'�_���H����#�e�l�[l����ݚ`+r�l�h��)�i������fd�ۢ&U<�ܕ���r�d�V�ɱ9�2�׶P�֋!��	�
�SN�0S�Uɶ�x�XːR͕�Nl��
���Qc�\Bla��0���)4���xm���/[
�Ĵ�VuMK�Y���D�qR�5ot]d�b�.��Bۤ�&cC��^\vi�Gpj8,[Ù��R�>��6D�t��pdg�ןCR
�p����aJS�E�����K!��b #�n�ʽ6�f�ak �Q��C#Ǚ��WRdt!�	yJ��1�/����bU*w��M�*OG�y���f�*e��Z��g� n��� �]m���EW�S�2��U�/�iÞw΍2���w+_e:4"��X^�c�7�v+�^d��� �^�w}�5�y���w2�q47)��ϝ|�lL/���3=3.-��D/�F��,я�כ*4�Ӝ����d��R���痉�]e�X;˫���~1W7~����ʹKr5z�X��V
���фb�6��B�\�/�&�(��[ {EWtiM�/�q��S�]V=�Tm�]t�$vubN�gI���1������tM36�P�:7�Q�}m���e�� ��[T6>ݐL��M̋{	e;��Z���QzW��CO�]��F��9Xf_!4eL����T���mڢ��Wf[��1s�Im���w����F��R���D��}A�a�Yzv\�d\�c�H����qVi�ԑ2����\��'8����Râ�j��c�W����ᥣ���f��Du���=J�&�f=�g]��s����\��iXn��C�n��1/�9kM��|&��jV#u�����r����uv�e�S����݃�@�s��;i��u7�Un���u��V���o�nb��Yŋ���+�p�ܗfYlo+�yG���n֊ӟ#vc�@���:`8��:��]6QԷ�m�����"De����i��/I4JEk�9��U�����iK�8�B���&h���Oo"!��.j�|:${r��r�1w\ӻ@�Mu���B�a#o��c��3U�9V��E���a���k��s���p���ԶfTL����r�z�-`�����n�#s�C�;�u!�y�o�S���0[�́��+3c��ǩAKrf�1.�ن�Ux���m]ö���T1VK�����>N�L�+�WƸ`��W�M��c4�A���w���I=�V;�[Q�w��ˡ͉��gf�	���Aw�i��$��4{� ���.��KM���gD��.ybVLeԘp���r{eê92�յ�e�T2�9{O�%�R���Ժ1X<�a�-N��t���9�ց��y:��$�;�_n���f��t�u�ڛ�%s\Tf݉^s�1զ>�/��nYN��;���
�����6��]1쿚ᙢ,�p��vT���6QO�/�h��lWR��]4V1o+���oX�F���jX���rYΛ���_F�e�f�ucN�.��'�/OTF� �I�h�a������W���� �Ŋ�o��Uk����bn�i�qYec����(bg1Ә�#{ʒ��M� �`�*��i�� vm����>cn�_h�iEi�#��κ9�b���>\Q��]!�����7f�/�hW7��G�K�3�A�aO�W.�)�ˊ�A,�,ռ.����1D��u�Z��V�Yu� �)*d�7�����RK�ig�b�i����q��-�T��_�[fy\�жf�#�HT�aŁ�Y�SAu^�G��u�1S"�r�3s�}�^�jJΫDP*���q��c��y�d�����H�v�C���:�ګf�I��
f'[n3ZVV��Z)�(YxW�5}su�}�r�RLjt�t!���q�|��ܪa�(�"S��P�����T4�n��j9�d�8u7{��uĦE�*���Șvm�r.��M��������2f Iۣ��%�R"�����:�jHf��� O����nZ��g����� "����8�ߔ�{�Mb@�2l"�P��Eb&�C��*�͠F�x9����z7�X��֘�b���%N��]��j�޼���mό�N,�ڰ�W;vbǪ���Yw"�Z{%(���fV�(h���"��e�]�p�z���j5o�O6fm�*\ӓ�����Yt�X��3[��W����U/RD�����6���ଋ�R��N�2�rsh�%�TU�n۪*�
+f�3�&ŗ�2k����>\���nR�l@����,E�1%l��ep�����6$fI�t�J�;k���o��E٬!k8�6�f(�q��b㬮�49��/W*!�VQ�df���,9��ɴ
�7��L:�FH��tmpYұ�Љ{΋3M���L�ψ��c'0�w,��Ѯ2�)�3Qܷ��*[u,�B�Pb���6i4�S�ӑ�S�F�Fh�ş�!�8o%
��U�ƀ%�ںj�0��R��J����.w�U�aє�?�4���Y��m|�[�b40H�3��c�ו(c9]�\��-rl��-�X�=��m��H��L�6�%�%��
�V�:���Y.�
�)���e2m��`ŷpAH��n>j�g�G���f�n����3Gk�����(.0�w����_6��P��b;{�.c��kCqsm y�z�ngٵ,�|m�z���$�y����;���2�q8�ߘ}*�`���k#ۧ�eQ�˝�
�v�=��j��*����H&�5|�'jw�E�D�)Q�+��3a�[aA�|αÇg�WC5^���"��@����=��J�݌om:���
(��1�0�$��6f�Z�t:v��g�G�ǁ}����M
��I�E�B����@m�d"��R.fe��k�b3�S4X2�Tz�Rm�pŃ*�5 ��O��C�pNi�bݏ��7���Ȭ�0�ӈ��Ԑ�<K����ڱ��d�w;����P>�ק��t��o��0]�@���𽫃XѺ+�(��j�n�&7�<�M�ئ�X��2�.�'���ת�#`#�����Ly�$��@{;� �n
�Xb�tPX5:���rm783�4o����h�񮹼��K.i���9r�Ž�昩�h[+B�8�{@���л�t�������-�)�j���t�ڲuL��5J�PB��5�h����a��^a����N̾-ID��Aں�ٜm��F�������<:�AO���Ӻ�龏H��V�Q^��$o�=9Ag��n������q�a�f\b:�� z-��Њ\��!��ؔW�7��p�΃�1�ŭc�]�J�rd�����7d��,���7�U�4�"t��xH�P;����$Z�A��:��u�����8ޗ�V������pp�i\,�ơr�qR� �
D�;��S�ȸ��?����e��s��mZ(ٍ�v+�`51�|��&��-o�	r�t��D+@!�F�8�*K��U��t�\�m�ؕ����`�y-+���oY��GRy.=%�id����BT,�6w�!6��g+�Ǚ�bVK�)��Mk�S��5���M�[9m���Z�ŋ��M�bJ}l_�4���ٌ��C�%����ۃ/Rl�.��p�x%�){���l�Z�c6����a	Yl���nn2:���I�� ��zPstC�]��b��a����JU}�!��f�$M�\+q��ڕ���RΜvA6�N���)��F����O~$��Ē엃*��.�F�^�ֵkC���r�C���B��qu�=/��r� ���4���Ջ![4�5�:�9�+�uf9�5�۪�l>�-��Z��.:��"t�������B����g�SY�{V�U�J.g.�N{�`쨾�"��k��Pu�7�jXJɨ�����:w�
C�VɎ�UJ�GC������H`��֔�� Q���x6�-��;�쌇x�
���p7�0��5-pb����|o��ԋ�+�v�]p!��Ha]Yn���*�Z �d2�0��2��ł�#����j�2�1\B��ܜ�ɧZ�9.�$op��ҝ[g	�:�[d�n�\@i�鯖R7�<�1;���92��Fs��9*������fQ�2�� l�Z�G^����гá٥��*ǖ�8RG�b� ;кnt���\�ĲJ�Vm�6�l�o\�5lB��.�4'Y�?-8]��ᩔw��WoLC�\�w.8Cv���E�c�˺H��g��+����dPLc�h5�1�u���m-�8q1_q�clgJ��d�WX���֭ͽ�x�|JhM�>�+^���2���`��ݲhf��l��˃(���n��R AW��'���Vvu��,m"h:o�f��`0��a�k��2�v�r�Aj��j���"i�3`�y*���lj��	�`�Y��~��Q�����eԘ���d �;#�m��>8�����2��J�ܽ���D�)2�[(���,��x��(��1�9m=W �gZe]vB��%J���AJ�q�Lx��[Z� ��&n"�a��Щ�S4��ޓ*�[�b���(�ì����` N�|�.KԔ��QS�%�dQ��ܾͩ�ܭVm$yئeFi���]��[h�Z'[�FTS2�tjL�Qk���\��63q8=Z�+u��)��QJ-�0��N�{x��*��.����01'����kO��OjmP�r��:e:B<#S�t��:���e»�f�C񹶌l��^D�v�����T%�it�Ɩ�w׽W�I��.,K]tUh�*^TkLy$�HuѾE�<�:�"�[O\|:�F��:�
�;��MV%�h�d9˸�jz;��E�E3K��`K�������x,p�6��Q����͠�ōfT
�Y{�K�8�b�o n�P��"Y�m��Y��Õ���)ľA&���[8Pl�,t��1O��6\�++o�Z�ڃ0P���*JC��d�;o��-*��Իg.!��	�	���q�tdBen.�pdT��繅AUOQ����W�Rq#�s�j9u��0v����"K+���9y�^�ng�˧,��÷m�_Q���;V�S��U���u\Q��ĦY����3��b.
*��.�˙���c�E0��f�[A��[}�ڵ��1v�F�׬O�e� ���to*��e����"u���ъ8q�u�=��P
龗X�:Hχk>ܳ�:��&W��B���L5�Ū�&�S3���,���جCq �U�ĥ�]Ӳ�;|Q)��m�r�e�J�lՁ�]]�r�B��Ud���,����r�ۤ\�q���E>��w�sb��tC�V�Zіj_pmT`�ͽv��x��81*����"9�Ҷcrn�x�O'lGR�wZ/v���51��,�ByU��\�\�ze^����Ŭ�E��ii�5_['�vvt�*ۖ�72Mީ��ac�Hl;J5�T�[W��@U�ꩵ��j�ʼ{�$%�بյR*�-�Sl�
W,�*�G'��1�h������2r'VŢ�.7�"�e�Vx�yx���'۾;�=�L�c꾰��}��J��c��"t�h�g3��f���v�Y�!��$���O@k��fq˼�KxF�д�wH�a��NLPQ}�f�nUH�w1��oA��E��M��d6�0WYFwU[���j9&Vmap�˦���G�]75�RD6�WG�x]l�{O{�1���v��ST�z�A��!k�:4�J�ū2�է\�n��;ެU�v$m-�����y�k(H�+a��9�.�h�� ��'���CBI�����P�Y��U�2i�K��Tښ	Ήi�k����s��A �1³�p�5-"�Q���+8@��U�[���>Z4Kq��i�0�#.�uF���).u��R���v[
q#IW1��j`�����
�}�Jt&5�H"Ɯ��Ҕ�*֗��U&ASe,���u��9=��k��g��B�Ph�4��~4�ҺM�yʳ��٣F��ΥMu�r�x��'�:�>-At�x�)=Y|�x��o:�6�yM����ym:ѳ9`��[:���N:�b�,�Ԛ��%M�.��)�=�vN�L�c_i�k3D;ʵ1��R�m'1ȷ-��sr�(��{�`�p��S��{���>h<�c�|m��OS��X���
����R�L;$S�͞���4�G��]
�f�c	�X����U�wT��V2�^�IWt��j0c"	 �(�j���G-l�ԅ@�t*TN�ɩ�{��U[ѫ�0�wv��e�is�@J	<9Ee�ز�;Ť�$��ӯH�D]����j����F}�&ۛ�{����9/>������i����'�\���:��ҧ�] w�]�w����&��&��)�Q
��d�4nM�6�1�G�h]�}K�	��.czl݅N�4gN��E��D��h����Gb^j�\���N�[���6*�̜�qKC� 6H�����eM� �I�Xќ�+71}�
�YZ�.4�pt�D���
��D8�ʷ&�i/�=b���p+��
�U�,|h�m�G9�H��Y��z�8u�=w}�*ji�96�$v�aA՟H]�_Y<ʳ��6���}җ�F�w�1V�Z���;�Ff�伖
Bߜ�7^��[��zf
��f^	u6\�e]j�p͗�U���})�.�d��L�v�]�̾3SEn�o(��,�Ӻ�f�D�Yy��'BE��ݛ�%�`z���m��Ɂ*��qm�9o*�Ag�P��HvT�[�>Z� ��Z����.Z�fƮ���Y�L�t�t#K�Y��X��׻V�.�:�`���}�1��5I��=ki�\[.����̩܉؇d��X;�,w�Ƒ�Xݛ�Lux�TW���l��7WD��Y��5l��q"��hX�	�'vFo�w+�[���!YA���u�wt�;t̶K�t���Nol[s���n�jȥN2�$���ٕ�Rev\X��Ɏ�TF#|�q�N�:=z�|���K;%�d��|�w&P)b#�����wZ���>.�PM��^u�jok���H��#��פ[���d*��&���<m�6?ݱ��}����������������m�X�͢K��Y�¥�M#���R��(H郘��3֐Ê�nP5��8n��CNY�v�����v_q�oA��J��wv��λz���wܲ�2�`�2��[(<��|��Ѭ��6:0RO��B�w*��p�k:�S!���
��">v�糣�{JHe��8�ǩC�2qd�5S{j��7K�+AQY��[�M�-=2�Uܹ��
�Au[�t�����)^e�,ޮ�t%��8�L�3seu�i�T�Y��R��u�5Z�y$j�_2ڨ���z����,��U1�
����;NY�Y�l��Iӭъ�!������2�й�SR1-+I�7E��t��ޗ(vP�<�Ƅ���.�<�Ԅ���Ja2�3uc�I���p,i�����Xȹ��pW�)����e��MPclZ���*�|5*N�C����=�q��oM���.���{.˥UJ�7[A���A��a�.�t��l��sj�J��}eK/!�ţ�]|�m@�a��Q�,\4ŏ����<�+�*X2qE��}��lpI���+Y�8\���R��E>2��9�KY[mMJ�W]@�e��1ՑyS�t��ʂ�����DN�1Y(aB�_6�1V�']��P� p�a�/P�n�Z���	�8mN��
&��	� �]�z�h+�
�����]��:�-@�N�3N�8W^2Yn��w�����\U����j��J�'*��8�pc;�p�.C^h�&��@`���=f�\l�ϝ��Y��1��T��O�tUaV��
8뮗o6'0�rE��(RU3w�W�PN��1*Vr��M�`m���:�ef�2䈒��6�>���I\�4���HV���
�+w�`��YI/ڗh��RSR����U�n⻏�2󲙫p6s�j�Ŝ�P��Q��ܙe�t���Z��F9�4�8��곽�v�-�;я��9���v��`�Z:K�/�LLW8�!�n�i��D8�
:��o,��+y,A��I��>Cz����ܶ��޳k�_-x�r��nk��$��) ��ދ+�A��0���J�7���z�9�!�쵙k�V�.f�hew%�������c������K���/�s�פ�;�$ ���f'bdѰ6���b��0T�аڧQ��#�2��WZ{���63�0�9��s@�;Y�w�{67�-$M�l:w���N�j�*�Q<�A��jO�ŵ�+���u��77n0�O������2��c�JYٳ�^�E����u�+wM�)��*�-g,����]����1WWϳf|�{8�S���L,
jT���C�Z�%m�k���1�����h�\�+�=��V�S|�Ү��w��7]����M���繺si���n	V`�f�)Y�5*�ώ�"Cxu�Ë"�G�H��ֶ ��
ZBUr�ؔ���R7��֮:a�1�Շ��ӮA0l�Ԕ����{Ō,���q�=��Y�g�X���#��S2Umk�Fpb>z�Ph ��%>;��yk1��̍���\V���M���[!���p�@��e������5���9�'��^9Za��7�}KgKTr�%cׁJ��.@��6�j�U�η|RP;�	
����w��,^r7EL��͚
�PT�o��� N�P��c�k'�"a该�n.�3^�5�d�{6�Dm Y��~�f�����.@XwCSUv�;�sAb:zl�+8i�'���7{��P7v����F=bLʻ����M�vR+�II2�;║�8�G�qn�W;�rY�	�u����]���+�DS*6ďEgeU�!�]NDͫ9E��Xk�nf�6�lݪ��G�v�+�̣�݆$�����.Fn\{�Κ1ug)Xɴ:��WK�[$f:���ٶ�����2��a�O�����Q���z�wl�ަ�6���Tmq�|�n����r�4�ڳ���0�AQUg%��\����Ĩ�ܹ��AAnBM^�Ը��t��R/��|�X�wJ<�QA��ug4P�޸�p�n՜�+Y�E`ӗ�;���*�.�*�I�UtUHLs�hu3	���I��u�
�`Տ�X�v>�} ��IeGe�{��k1�ޜS����1D�3���GY;sۨ�5EޕoM�@��ÄV��)�!�۔�X#J��є�♑�v/GA繨`=L��:��f����s^'��uα"d�Zr�B�-���fvN����60�)JWs��=�t�Ҩ�w}�1��(��:��BՋέʱf����͆��]̩�v
d�Ꮁ����ݜ@�۰�h5�W�k�R���[�pb�9�n�ea���=]��9F/��p,Ԩ���!��E0���;�隆.��զ�eLM,V�-7F'ptWw_H*,�Vi4u��R���{rD^�EU�.��!ӛ0)ql1�Hn�����iO(��Was���ޔ o5&�e#ժ��r�{{�:7��2lrD��ڻ�q�]t�3�XG�����S
�Aː&ݾ3�D�:<Y3�V���a�j����������`�=[�]owd���)ڭ��T�����@��!��۠Z��,1�ǖ�0$�@�7��Ww�B�������Cr����($��hA���2�K��K���n�aN^�A-zH������W:�䚣`�gǦ���-!X�wUЗp�eX���f �Kx0
�K����V/��r���l�vo5�� �o����:FN�LʋX�x��:�`�x�j��MESL-Ѯ�cU+�ʖS{�ҳoE�5�xz^�`�s�l�p��w�hJq�{k:d�����3�hcE<��7�K1����qw�,�v̗�6\j�GbM.r�R���[ʆ�uҝoaOE���8������o���Q��¥��@��,
�jt�\���tw[kC9Pk�-\�z�R��I�b��O��c�h�A�"
&�D�w*�⪲�z���'GkF$`�~>���7u����Js�����:���/`2��{���]��� 9c��+�z���F�)1���u��]Ҭ�ʄf]!�E޼5�/,s��#c*�E��˖@;	��4Cb���X*�V3��6�+3�m���pnr��6w7ƶ�5K����7l[���	��C���b�gy��x���};W��@۶E�}���8����F�JL�:˹^WE��M,P�Q7X���j���l�ҥ��KݽG۾�O�1��S ����v��M����B���#��x\��n�\��z��������/��Yl��	�N��k8n"ydl�7��[.�V�
�Q�����g�2K�r⻺aV�ޥ�b���k����'�H�5�M�=4i������8P���Kb�Ѩ]�!sGwY|��Wۤ�6S���+֪���/y	!�Fm��[��ےd!\�rњo.ne��Ff�o9VE6_S�X�9��#m�CM�w˷kH�I�q- ^�`sƸ�LW�d�R�l���jx&C�Ҡ�n_I�IL;�-��nRAK�ZU�z�����]�z`G	�4�:�i�<�|��$Ҧ̐;
����n�ܧG�����4�|Xɤǵ�K�ٝ�H"��!�t2�f=�#�]WSji��-��MފĲ�`����q���nU;�%a�/L�ǖ-�]v��KY"�)��܏�m���M��IM#�i}�#��gGs��}��:�W+�,�Y�%��o.�.�t��.6Ղd���+B��p�F�G/�jn�������	�C��kUmN}`.�_\%��8^"�{}{�d�d�)f
.�D�&l��Xȭ�.-�Q�L*�
�=�3s����Mr�fv�L፬���*N�.qk9�v�0=Gn���W[�+F�A瓩c�6S�2�{6��'L�������s�����`jdv���A�����C�b'�u܌G�S+�)���u���P'��jF������(i�0���5��˝8_#[�9�AQ�@�7z�YH��"4���13��ȥY���~��s6����%���-�}�$���{�;d�RmӊWYV'"��=u�hD�cv�&v�2������bzR�m�WI֖Fʚ)Z�/+j1�)ٕ%�nmT��8!s@��$�x�3B� �빍�vwBn�n����X��
�n����؞pY�:ƻ5�A��I�����:�I�QhSkZ�b����r�L�|�_v�FV�s���:W"�;��(���)�����]9�u�i�
�QD='���Z�c&5�*���clcz�Wh��:ޞ8�\�Ѯ����K<���ھX���s��A��M��ֳ�v�>�,&Z�0cK�%���2v�t�2�;����:�y�0RnE�98���}�]�j�:˘r��m��3;���WOPQ�@�Ef�L;�}Z�f.������1ېqJ5s�(`D�6�l�p������|�OT�f��yu�� 4E�yͰwk�����ٽ.��q�Uԕ����
e.�'����sm���gv������6���)x��2�F���:Eڮ�S�����>+]�H�l���>1Vh}#�]j�� �=�vtU����l`g@��F$i��=ۆ&�%AE��Ŝ���c�e�}s�J�Bmd�-ڨ��Yn�p�[��{�[aF9�e�6�Kr�aֹ���򺷦9��������z���A�Ff��9��V�J(T�n���v �x�]�t�uh�vQ�f�p�u��ۙ�˕�dčV^�U]S-��;�8�*���j%q�f��@e6ӹ��vL���ʜ�RN��(��ZFͧ��l��"�$ �`��rK�6%^Ļh-����)p���({K���;u�/�\+�pɳ�=��zY�m����R���(�&i��Bf[t�;��Ya�iŋr���j�v�6�F���Nx�L�'vt3!�՛�,F��* kc�i$��m4bt�ƥ��&v\Z�*�i������w}K�:���w�&����s#�7��F���r�����T�g	%ۜ����w��ӕ�L�/��:���<mW��-�S?m�-�X���r�z�����:Ҧ���6����3:mDA����/���
C®l�	Ǖ44ũ9R�1��� �ϱ:�o%k�\6.,}rͰ����ƀ{j� �V��3,;�y���V�rm�+i�υ֪���t� .���\6��w�)`�.C�yFZI�6�S!x���r��)�μ)N.U2vi�v����Bi��$r�� ���fQ�X1�yf�ú%��Ss+�����'���g���p���d�d>�e�uтs�	g����lg�탄ې���Z�?�E=�)�N�7��t^m3�5w: �pf��-��FWU0��Ƿz��X�����[ڭQ�,��`e�8�x�2ԊP_h�1$"�_��R�+�Hd�:���$��i�h�[�9��wTW���6m�M�q��T�ub����b%�=%�-��Yas��r�=C6i�vص/y�×(-�(�h��/�-�_{ӭ��-����)[$_M��8#[�q�s�^���rh�˷M�����*�7zlMm��/䱩]42��cS^h���s'm!hS�V��$�l3��_<Z���x^�����Քn٭���ͤ(X�@&�c&.g-��Ù��fp��ԏ�_bH�QVL�:�j��Z�u>�t�����/m��~sv������_�@�1���:n������]6�[)��Y�Z�N.��|�R�����d
uA��U�!V 4.�GY{B.m�P���}�Y�η5j�'s5��%^���F�������C,��T�K�S�����\\2*�l߮�em����F�l4���0��wB�Z�	J����XWْ�|�-�Iq��$�맹`St����չ��t@@c*f�I���N��,	���� H�ݒ�Y��X�0]��$�����S����M��o��E�U�dObT��'��Gޯ)�cޅ
�J�w]f����|�eX�[[@����p�"�W#�+�E���u��V%�Y�}�)�v�caQ�K)�`���rsݽ�Cq�j�,����]K�M;v�ƹWSv����|{.�|��;�U�ᛝliL��F5��6��ot�Fl���='j��U�,*�r�!�
���N��!O�S����qX�k�t�tKg�v�mg5ũ�B�������^�``�4��q���j�c[x�Yje�,cӴ��[gI���r�"H�bZ�uÇ$I[������L�]����n���dWfLws�� !vY�᛺�&]�����Ѹ1�u�b'��&;�y��]�v�uꣶu�ɢ���l�a�t�8H���=�o�4�ژ֌�(5��c�naS�莨if�b�I޺X��k�3h�v�t�ܻS�HX�֧��p�5���]�&I�	}x]��r� �����M�-�M��EX6�۝!EA�`a��4QwƣV��bnSr�e�q$��:�KP'g`�
#-XE��R1�xzM��zU����S�[̓��������щ��\<���e�Vq9�T�9�o0��^Ff�BS�sVa�;�S&�kǧ��<6�i�0=�S���܋�WS�e,�(7\#l��w��z���K�ܺ1����JR�ٝ\Τ^�e�a�3��zZ��,N��K C}iJ��lNI<�e��vt���t͛�5��s��[[-�WbS��"3�sY8[}�l?]��|8��3�s�d�Zz�u:�Ѷ�)�j�U��jQ���u�7p�<�J�ڒ^�׽�HX��Z7��(��[�y�����;�#�lm���r �+�H�9�
c��$s ˈr=v;+Y% /�<ɠn<�8���>|�������/� 6 ������v�����5R���eݐ-մp-'�cw�����<��^��ˉ@�s+�rJ�ۛȺ��a�ٕ�&�9�2�	�ų7r�{�������c*�L9�S�LoU��6��қ��.��U1*Cv���j�؛���R�sͱ����i��t9P�����+�yR�$Ӧ��f����D]7��/Nq���:tf'��:p��a��hS<\ۼ���2Dق����cX3��b*}\Ӫ��������
�KĹ�:ٻ(P�ם��Y.M5ó����7��kL������iҨ�V��/�O�%��5r�t�]���ָ̡���(����ω��])��A��ת�K���z۫X�t_5��8�Ra�%��%��W��p�<+p��=�B��cq�4���.��+1��0E>Mj���٬oI��?�!mh���ceդ�}7�I�C����E�q�\���cR�x;+�6vm�h�no��r�-e��xۤsA�m仂�����(؍�����Шv��;oU!2�c�뚔z���]t�t�T�ϥ�0I�>��Hm�� ��D8��]��]�/������mN������Y�!��Z�9E\��5h'	���v����f��\v��� �l��"�]�u.$2�2<و�/��{S�0��V>A�¤���ȓv�6Ey�ƭ�*�2�MWD"�������]�p��F��a+���G7qܓCNU�Y�ww�f(��D'���z��pW]�'�ݮ�냞:�'RAur��V��2wB9�sTaHg/\
�(fI�n���=�5t�r�)��\��0�V�t�Z����r*��e�qQ'VUF��ū@ԊwNx�+-"�%S<ܒ��,�I�T=\��H��ui�9��fWKJ��J-9*�
�1�%�n�EJ���p�j�13C"�*��GP���Ҍ�2�̽/q/D�%������2�U�W<�$�T{���LȨ4��'Wt�+(#�-$��+��+MCD�f��TI��Y��"��;��":�HVl����M���{"���t�f���w2ÚU�w,$��ﻓ�`�pN��� �%��s'40�C�ٹ0�����֝��Ƶ-�s&n��#S56���Y�̬��o�]��d���_mU��@����x���+�{l�@�AnJ5ne�(��(֐�{9��i竦Y�w=�	���A(�̿����;bz-�;k�`�(�D����p�z]�T���3S)@gK�uP	�uX"�+ 4Y+7��X%<-�s��S��
Z��B9Y�`�q�{z��k�U;*�+WD௵�|/Q�Y�-X��D�]�Д�V�%l�>��"��f�����j��5�ry�Պ��Θ�����q'���Y� �����n�[&(?�g-2��Es$t[�^1���S�N���U}����z.j,�c-����.A��צ��L��o�hJ�6y�+:I��!�Ϸ\b�Ɲh����u,�q��Jx���2��<e��Ե���4��Q��1]�Vc���!/S��`|�;S�OSuox�H�����',p�ޓ�g,?�c��M�<벭.?8k�宠*\s-�	^�!��nhwF��ZXS)���ƊF��^���\=�)��[��sH35�I����v�o��K�Bg&F��s�cl
E����Q�)W�m����w�4ū/_���񍙢m��{������x���ē�L�:�����I�<��#ަݛ�yH��+6�-��0:�H�.���a2)�#�]\���"s�1�U,lt��N�)�ӂ4�㹼��#���A�-Os�R5D���Eև��,d�!��Y�x�/f�f�9�YF86(�4_9y��O��h�|ڿ���9�X&!�yq�k�{��3�V�֛B�\x%��O�����$a�ځ�R0�q�E�@�n@C\7=QW�
���v�w��=��2:E�y���F80�u"9�~ar�=�%���q317�B�5[c���z ���]�$g�T�$ ����z�W��Wh���&xk����%��|�յ��\�dM�&��D�����"y���^�D5j�,�_i�o^�+ï�X�sD��.a��s�bZ������za�6�w�J��Q���%������VLX���Y(\B2\�6�I�z��y*�Q���]±qm�J�X���|Ǫ �T�H�:���$�V><dn�q�t,����<SAn��qU}y��u��Oݺ g�!/��r�XY�S � ���:�4.� ��ܣnȽim)�"���ة�����Q��R��̓�#MsR��O ���wyݑ�()0:N�B�@:֍K�.n��-QU��{�����Tݘ�S/V���\{����#Tq�,u������ju�Q���frN���qNfG�^��Fr�i�Q�Ws�9����ںN}E<�;V){:E��M&o�2we�C2f��OMS���e͠+�Z�i�P�j쑬���މkJ���q�q�Ba���[��ﭑ�L0F�2�ʎ���e:�y��U���&G�*9�`�=��q�7MCx��}�x�#!"h�;2�Ո�g,�����V�Pф�/&{��ܫqܽ^�/�W!��<�>޹\�0�&�U�V�Y� 5s��x�v�Y�q$�}����c�ؾ�*�妱�4k�Xc�n^�5<�T��2hWf�ئ�ge�&���z\���^�e��3�9lo�'�n� v�cK�n˃�&�a��r��bY��"ÍWP����\A .��P�;)���#B�����(�+(�J�vN,��)9��	��f}�����R��W>�`�|b�5�71�n-�����q#��&�u�7ƈ�E�S� l;v��bL]_uq!�{8�̺]�znC0yk�BAe�͜=C�6y�d�6����HYS�uI��-�^���b�h_֊�EAɻl��u�q�HV�M��t�Jwx0�(ګn�"oZ��eCbظ�X� �U�V������]���U�zh��(:�#����c�ʖ���壆���]��+d�d�J,˺�{�����y�g>�g��N3 3������4�nt�+�>��؎��;�:�k�P�Y��Y��Ie�>�`>M�Z�]������]����`��4��:L1_6��f�F̶ �Z�fGM7T�5]T:˂l@��'�X��b�0i7��=���K+�;��X�z5u�2ݼC�gHq���Ӫ�K����]xe���������╗+��.�.[
a�*�^��G��;+.'5ȁ�ө�cs'����&���S��4�ոh8����oL��	�g0W�3��@c�Q�]�@�7I����Mb����$f��n� $��W��=�)��O��U�Z_��jC�� 
�b��2΍n놾�<+Wg�"���<J���Ƒ��F�mfB�P:�3��L�Iw��e�1�.��7�)��Y|z� ��_tO��a����'��uБ�\K������u�E�\�9��}�����iN��|����'���+dVJ�y��mg��	�L�yp�;JYH6=�8~�+e��òJlgZ�4��Y�y�ʤWt�]�o[��C����n�L�na0ʳi<hp�FA�]ϣ�+)|\�&�87r�&�=S�����s"�PEb���VClQx�1
��Ѽ�V�F������[b�$��u��hNPˑhc�c�:�N��Խ\&��S\G�B֐��O�P�mL��2r�#Ǘ
Z��9K.�}��$}�3C�;ج�xl�w�u
8lo*��.;%�֏�r�v�Ջ�4���\M9��aG���Ϟ���Beu�=r|{'��|��u�-t-q&�jd#^�0���z֜�&l}[=<�^֘<(K���6vU�����+rY�#���VX<�`	oT"��������'��-gq�6Nډ��7"�Yfl	�"w��.!>�g�nܑ�g;i1�Z�^	�pX�]�j�ȁv����B��['B���
����f�E�-!P�\�OWY�mH��uX"�Y2�YFX��_E�|��2�	�隋cP����O%�W�M�3/W����z�� u�k��=�=P�A���Z�����	�#>�Nۋ���m�z��� W>)�F�W��8�u w����A��w�Q�]�a1[�Ń �Pή��U��=1���,\���$��zK�j&�8���9#��ֻ̳��A�'��Ju���K>{�CK�Q�mBf�X�W���Xhk�r���*=o{��*HBtP���Z:Y	^��x�Jm*��c�Â)��»ЧioVa�v��GQ�^CBZ�c������!zv	R>�Lj�Df�@	�6�p��N\j���Y��ע��C}���lW?��C(p��4<)��+��g[0���4�R�hԛJ�
�%�==N��g�E(���[}���y���8j�]C��8Z(��;����9D� U�.�c�>u��k�	�{m�;}��KO���J��(��=��]׭c)uEJ��wU����+Kܘ��F4s8�Q J-j���cuዯ�ޘBsz־��޷v������t����4Wj{��j���	C��WGz�s�6O^���kz������C%X L��\#���B㹷�dq��w>r0�v�R1f�6'�R��x��5����|�7�%���k|�͓Z=%��u�Ѓ]�q���r�u��ї ��En3��P׉��eu�<i���M�a���(�ګϽy:CXxKkR�.�O��|�Ƚ,��`��:�S�"a�E�'��aa�z�Po+����ɔ� k�����uo����T1p\�.NJ������t�����!o������[�zZArQU�T��==٥�T��R����2�ћ�it���M��)R��T�{�#�B�*����/�A��w�l����sU��Vmӄ.�,�{�p�Z٠����Q����@��Ȯ �os�j� �9�o��9���:^9O%��qgt��9���f��t�K4G�8~�bGs�b�{P=0L{m�[
srƕM�L�Tc�No�N�1��v=/�� 񢋥��ב)iҗ1݌�4v�E© ��0w���6��j.rS=�<�T	uHl�j/����L�dq�.C�����do��UsĢZ�q"o��~�~��Y�W|��"�ϐ�vvP~J@�D0e֊��<�@.���5�ِ��CYGLYr��C.2��2Z������֕Y��7M7v�5+�f�MwXqΣտ:�C���
�����7JՂ#��蝞����زG�Ǜ��S/�kym>��6��=�`X�4�+���Q�h�H�4+bk��.ktg_�=j�`u�7�+��.�L�~�MS��7��S}e��f��\M*+s�K�1bOx��m�&D;�LO1�.����}��"�>�$w>7o��qWV�C���s����Y�AB�zK��K����ǙT����C�P���W)������鏻�e�2���g�$x�k�5�]���h��ps���;;���(CD��gzֻ;fY|�����Ç���0��\��­6�W��y���x�Z�@�X���9�,AEdl�X%L��2Ң�*����L��j�+��Ӯ��m�=�J)��(wGQ�'9�����5]DI����Xe���	MA<1Q'�%#��\^tmBDB�+�f�����D9���~�$���Տ��@��[��_Z��	�A
��	0y���|a�D�Һ��UuI,�>��E��$�����-�U�c�"�U) \&&�����~S�;}�{q��.-Lh�pzV�+79䇅�Nb��*��f#���5ji�iZ���mRJ/�WϽ:���ÿ" ���ύ�x�5 c��1��<�.�=��а]��`���F�>����;D�\�;�unEE��O;j-#��4Kj̤%�c�ͨ�ތ}��S���L�P�64@!'�X��3�鿳v�^m>7�4A�Ʉ�]�*]���S�p]gLR��;a�UK"�a�M�C�����0�\O���b��a��ٴU���.�tQ9��^��}�*���.�	�{9�S�˹��T]��I
#��*^�^p�y��o�z7���PwG�2^�WH�7PKn"z����)�W�t�5 n��M<��ޮ��zƾ�k��D��>���ߕ�\��Xt�52r�Q�%=������0�	\��y�dЂOX��^�t3t���`��{�ҡ0��V���`#�(���CNf�cgI2�;P>8EWNR�cU�o;w��*٨�'gD�J�/���m�r��2���{�99��/"�u��ʥ��n��L8|H�t��PB��j�o��� Vt�.��v��>ծeq47����k��'�H��t�|�2�Z�1>�]ӆ�C�淪_�f��hwe��M����)Ʒ���{���l�L�W|g��ܪ�@�o�2p�����h#;�� �sȡX\no\,�]6sO�n��(�<c:�}i�4¶NSh��V�U�_��q��u~���
5z��n�|���s�<�#��v6\�0�H�O��h	�]���n��\��tE�� c=�~.a���:��_Ơ���o'����ǐ۪1s�b��Dүx�9=v��AH��ۊ�LM���X(:��i6"TЊ�><?�H��l�>Y�t���;וAi�@F��['mD�a���7a��0�f��Yq�x���zRNf���\Thb��7��u" !��~B�^Q
��ɨҴ�"S�X��)l��e�!'��\�I�����4����mL�����F�-9Z�l$�*�|�<y�6�W^3­��@SO�(��1�|��j�&�Ng;�/��Y�v���� ��]/s�Pw��mbGO5Q��+9�zX��<#���)s�L�H�,k�O;���B�����3���q}�T��o�<�8ԀѹuLE�d	��d�ȹ�#E�(1�y_.�v���:Zҝރ��n�cs)�O�N�&���f�W�^����*t�uZ�l�Ä�j\�c���)�_�+�c��������ҁ���;�U�z���=�ڣ�Ȑ���*��Z�R�,��?p���P�XV]���p�T��Q��؁�5\:��$�-�}���2�ip���w`�墻�dY��_X���U�l� Z߶�1�@�Ƭ ����|�`��>6��B���]���'�X�pk1Z2���'�)xi�������%F�Jv�O�e*ꍳ6��������\0J��z6�X?�cAĸ���5G �C*+[�ݛQ������jn5�.��r�H�<��H���P��V�*��A:js�E��o��&�s̱�(;��o>y�p`y� ������X7R���}�|鰴�ʞ\���IHn*�uL� LQ�{j�H{=`�vǶ�<�u�Ě>����&��?��C�؏_\��&�����o�^�j��t�"�Y��ps� �s��(;(�y�G�(�	X��:�<�uM�N�no���z��Xj���=�d
^lX�����j�28�+�� u�eE�N�u; �x0>�w�p�
��2�T§��n�dmF�|�]{����I^6t�`FS�3%�C��T2NS�sh��ҦT{Y��^�J�>��o�K�k7AF��,aVlT޵�>�t������R�[v�=�X�^��*t�A51^��SgJ�+y+5{%X5{���
�%$_���&��.�MEB�ŻVm�;�a�46	��wv-�V�Ҳ_b��E�1�f�`�o�%�Edg�R)*�q�5ھAgX�RL)y���L9��/x�Ճo�i0�C�AdP�w��#oC�uf�V��P-[�S��C�.�W��+@������vTZ��˵�0��D�<:B��W�5�j�i@�Z�Y-w!����j����]Asz�Pԓؤ�nvb����U��f�7N뼫̭�R�A�%3l�8�Mj��[Zv=R�����G
ΛBN�Av�!��Xx���S�Pv�w�5��7�M���ŝYi��q�Г�`�@�j���=;�v���1�ve]Ů�w8�N�o�Q�啭>�\l���Ot�>�6�����Q��u���'�vQ�N���:��n����Ҕ�u�n�םH���R"Z��
��a�]���֮�aO2�����Y&<����Y����qT-��s[��f�r���tJ��(������L����}�wM�������m��[4P-+~y2R}WM�3��������tK�c���44[���s��3���0�b42�:�B\I��72l
@�l�d,�ˣ�(��f�O�
�����)X�v����F�!�w���&�&w�$��Y/Y+!����K�u���� %J���M�n����6�A�5�\T�{gnP�t��@�"1��b�5��*�1)��f<Q`&��b�r��I)���j;�v'�"[�����YԻ��W�d׊����W���α�I���@�W-軏�"�ҵ�+F��ꥨLׯ�{n�M��r&��7��۰Ή%ϗe�s��8�S{*�a���/���`����inr�ʭ�E��`�}	�a��4ЌE���p��^3$4j�Z*�F���F߫���N
���#���g2F]c.��Lv-u{.g��gb�����H�j!3�p�3[�(̾�{��]uWi���k(Y�mkX1�PhM�	e���>���F�Q�����U'�7�y��j�3^Nӈ��[�R�UB� �OϡAW.5ݖ�Mn`�2á�9A9�󧖝���L2GOu68G��Ut�9Z7D1Vm�)\˰�iaz�M�\�Z�f��� ��oz�'R�h�|��`�]lo/��k˗��uh�#�-�Q�sknY�v:�ho�к&�3�щ2�w!�����b;4�a'DL�����j��#�	�8�6�¸O���ƀ�CN:�ܠ��
�|rC��h��!����2]uR#�JL�U�������T�ܡ�R�W,Ӗ&�2���IJQh���+�!�z;�XsH��=ܻ�D�T��\�4,���Y��(�h]P�Ȩu-�Z��%�r�ݹFTh["�C"2��'�wY\�+!+��.����C#ԃ�t�B=fX��Kp�\�*4���1P/2�D���Tᢥ丅,��	9��Fje(��T�VI�.������XIT%WI���Ttr)���/'L$�;����BRS5̼T̍T$����!*3�r��/K(�g#+"�A�ģʱ,(�؝R��uܯSd��S�&bb(��y�+���T�QN�zjs	g���ANi)	`TQ��uu�=pMC3�,�!SG=#1&�.��<�ss��Ȯ�Z$娡����l��$0�i��Ey�;�x�NV�t���O�֔&N�k6�⇹�q-�QW.X�+`mFio]�Yʕu��@��t�7n=���5�toS}3	���#��i�C⏠�IB��D�_���q�s���S�z<ǔ	8>3��|w�<��=��{�ܨ|q'�={��a�c�7�}�]�4��A��xG��>�DB�=C���!�ڛ;b��4�$
 2${�_��	�ݯ'�>?8<�ô�?y��>������xI��@�P��~8�����<��Ǉ˂w���?�ˏ����Aq��ȳ�	A�=��Q����};�'}}ٙ<�t����E���
0w�����������<��BN~&���zM����Wϯ޼�7!8~�c��,�������봏��.ܛ��I�Įǣ�����Ϸg���n��K{�<���n>滽"(}$F��ӟ߼v����z�;~�<�q�?��~BpwϾ<������Î}���'�iӾ��������������]ɤӼ}��a~��n��^���}I��4�.�Z�k:�}�}B��>������S�����|����q��ޭ����:�:90��>���o�xL/�߼x���?����@Y�����I����׏.��r}C��)���z�7�~��#~�� D!�{Oǈ���C�z�o*�i����}M?��ۑC��]Hzq&���v�|��}\��>��o�|o.'��0��ｷ���w*o'�߼�p/�;=�j������4߹�%8��"\���nBO>;�r�F�~C�B1�$xH��E�,� 2<	㞸< ����!����7�s�;Ŕ�P�N.�Ϟ<?�$ߐ����o. ��HU�����3-O���?������������.�o_߽x�w�p.���i�n}8��s��&��Ǐ�<�}M������yL*�'�=���Гy=�����?�(b� ���� ƚ���u�I"~���7���P���"#�+���� ��>)����o)��۷y�?&�i'��y���v�z>������y��xM!>��'>���>��i�Ǐ��G�}�"|c�,}C胃VN$C㳓��.�̊-_,� >�#��G��"C��?���$��q��{w�9?����w�¨|q'�x>!�0�P���ߌJ��ӷ߷���&�����ǎ7�<!�5Ԟw�nM�	ߒ��|��~?�[쒗���[F��-q�L���O��vyXXjn��� QŰ!h�CU�3n���jy�B�l�g��=�]Y�FM�����'�h7P�W�-���
���� 4��͡��M�n��j�{6����i�Af����Z��IA[o'Rr�QA��:��!��������__����H}w+���nL/����|�ۏ�'�=~��(}C�r|M�9�/_|`�|C�G����zL.ޏ!��py>�/�@0�}"�G�) B������g���>&�	��`��P�6>&��yq#��]&G�0�H1 ������q��? q���ϺW�8�Y���}�`��dyY�^��N�J�� ��G�"$_����O	�!!挾]�';�xO'�y@����|v�~&��yެ~w�>��y�xC�a��]������r���8�o��nӼ���C�}v��}���ߩ����^�����ԏDh��D�߾������bC�i�~��o?��aw������ܛ��ra?��)����w���P�$��Տ��|w�;�o/��yL.>8�����yL/���;n7����r�#�Or;���h�0��ӏ�������ǿ��zM! aS��H�=����lT{���@�,wpN�}~�$���I��y�&�G������}A��\|IG���Ć����Y;�D��[�#�'�@��G���$�@��1��@�9v�߭������{��<&����y��SxBt��X���}��xq8��l��e7!�����=l �}�Dxݛ�ʙ��{�x��I�>�)����{w>���>8��O_x��S�aw�;���~�8/� {I7�}������Ӑ������}쮘��q�<�� *�=�}#���8Y�Q��9y��t���"$G�I��>��܁���<"�����}n��	�����[)��>�x?�q�=?�&����v��<&�w��}����F�F>� @��G�������,�C�fZ�k�����#P��A�����r;�(xL.='�w�܇&Ǟ���U�N������������V<&����<�<p��I��>O�x��������w���˧����{���L{e���=�z ��� ���S
ay���������y�yA���3�_�YG�>�P�`aAɅ<�����Os�>�s�Ă�w�<�G��&����^v����an�?T�O7t�e��r[-��&^�ţ�)�L˼�)9�Ά�%�5	�O�1fo��v��Fҹ3;�0�IMQ�Nnܕ=#�E�EQ_|]v��E&�.��V�y7^�E.���b�Y��{���F��Z/t��O�$� "=w�>�#�����C�iH}No6܋�i߾�!㭾;�Ǔ�pxM���{����!����������=��|����؏� ��D}"#'�g�k��Y�����C=M�"�@>�"$G��h��`�������{&��|�����һ�5������OW�^1'�>&�~E$]�3���<~��i	>;{y�x����D���G�X��AE^�>���(ڽ���..!�}L��=�G�}����	��+����_���_ɾ}�|!����	/��0~|�þ!�追�hxL*����ߌyNC���~�ǎ��r��5�?�$>&�h��|��׻9�s�łՊ�Y�}���",G����8�]����]�7�>�q�����|!�|����$������P?�\�q�?'��'���!�9��n=�Q�H��̀��#�������v����uː>b>#�"0F��w���m� ����x��}I7��G���v�ߐ�X����;���P��q>���������}����v�t�>w�}��y�m��W{���7���n�bz�'*���������!��Ϟ��nO�Ʌ?ｦ�M������+���>O�~�~N�>>\rԝ��xq��ߩ�Ƿ��oΕ�P������ׯ��o_-�ٟ<��㽝�V��Մ��!�O�'}w��}BO�oǏ��\
ohO���ߍ���8$>{���������۝;˵�7��x��p"q�����d>'�9�������Wӻ����@<�c�� ��P�"0U?���>��M�{������������P?$��i��ϯ�oI��!�}���I�\
o�G��˧k���^��t����OG�w�i$��>��@ G�F ����ז�o�������|q���ypH|C�rz<�����aw��Q����P�G{��U7�H'����<3��<����ސ>���pxN~;ro����xt�+�"�?C>�>�����#�ӏaVG����]�k}`���=F4E�|D������叮9_[�&���!��o�����y>}���7����~~���M��O��p
�{IǏ?��X� c�#ӕ"<(}"!�1검J:��T�F�ڃV���dZ�\HOHv3�q��w�@撮;J[�.��L�^B���8��R� �nڼË*f5�ٰZN�7��������v��p��x*��hTM������X�ս����}�1�5yܚ���+��k��7"����c�t�s�=��C�^��P���]�?oxM�	��������}Mϳ����]�3�>�q�&���|����\
nwϾ9~;~N~�$����B},���z���ǌ|�J�W���SI�Y�x����">� �� {y�}���0��L�S����S��������P�90�=���O�{C�뭹�������@���Й��!>�4#��T��Uf����<�|���.�\��3«hL���Ve��ņnEC�܂Ƒ{χ0��*n�a��:�U������07��_��9��A�<7A��q���V�Iq�À��-�vr��'��ï�;�-��Q.�XV@����.i��(1�l�N2�$4��\����W���9W	����3_i��+��Q��({�.��u\)�4a� u��Z"�b�!��;�{Ou
���]]"�qN�4� ���ƻc$	�z�Ϻ�$Ź��:�U��UjARƔF�8�@J�G�/<���ִ�����Ь�8��g׏m�0�o[��9���DJ	�ng�'7�V�Տ���W#�'ʰ-�
�����1��ʸ�dJz^�*�lQ���x˭����^}+����l��D�.��|E/qe�]yI�m�K�:	��m
�od%_i���p\�}����xƔjX�={�0�GX���V�.��WP�DWf�:�Ӧe��Ҏ�FV\t�)�هC��hd�rK�eV�c��'����8Λ�'f�ٜ����Q�-��{�pS=n��oI���D�z5.�n�sܫJ(��_,ʁ:_��Q��Ӱ�1�n��k���W��ӷ�k�KO��,�i�焻���y�%�}�1���"�w)��SA �����R;&4R5�3T�A�=��sG�G۲��\^(�5��+��X�،z^��&���}��»T���S�q���T����t��/bU�9��t���3v��dg�*@X�˟D3�� ��yl��Z(_6����ue^B�F&�ȴ��[|��˻���Z�Z�+�K?w�;C�6���Ϭ�Z=%�]P�ㄋ}{�|vQ/1�B���d�����ܑ����嚅��c���B��x@H�Url��G`Of�N:KJ��զ�/�0ٯ���y��S� HMPe���<>or�C�us[̺��zie`�wN|J�Qɚ���b�.q$��;����A�~\t	͘v�[xsm`��Fޝy\��]$:��b��n��Q�%������ܠ=r+�)�U��N�a�?_&�����r�(hi�qjG��/��4�F�i載KN����e��7P��U#�Q����X�W@��}t��ӓ�`9�1�f�8��=��a>Ǜ�4rS-OU��O+�t-�Fӌ`��=�{E�c�]����b�g.� �l^ȃ
�2����E�B�@�Q�%%y�	�z�܂󁪐�S��,��AS���S�)������� ��m�T���n����Wf�U�֢��NI��ǉ��*,y��֎ոy�B3�<�D�0E�k}Q�8d^cNJX�ϯ��rՇV{��m�X닻ɯ��Y�$�L{;�i2; *P9O&`w2h��V��d�%JRY�:F��"u���;�;��u��;겾��n���M~G�{]�e��{�F̓>5��J!�b�~Â\t�=y3�cY����O6��=�E��ݪ�_e=�d��_A5�V�;�/w4��U%

��E�ǥ�<`Ku��|R�J���ٴ���������.��#u��s��~[p�8:a�ȇ�'�����kz#I~�x��<Ƙ����Tc(gL���E��rHޅ��v�[)�D|k�v�9ɣ��*��1�U��^�S݂`N<�B��hP�����ـ��]�83���B휦7u�&��h(kN��uk���XQ��3�Ա�pw]�rĨ����?5.��Crr7�pU�W"۪���@�׬[��Q	�u��6�sv�tҍNF��8S�S�6
�q�2�1��9h��h��/�؞h��gkg.��z��-�oQ*�q�9�Ӎ*3��5;YN�����l��-��Az�6��آ��YJ�s)}�+�qE���D7��ry;s�x�Xb��a��l�ZJ�n&t6CSQ��N���ۻr@��k��.����p�eD�nX�g��6�*�cM�%l�yч����)*9���M;K)�����u�+�Oy�{���z�_$���ƪ��nB�/7�yI�p*���g;��4�kX��}����F.#�e;u�-����]U������i����:�Y�Y�l�b���S"�	~�-b��.��֪��*�NI���`�[2��9ُ.(0���w�mr4�����:Aم�@�,i���V
�7�1L�omz��y����~��Z����/�uf��D�oC�"�Y���B�݀
WoD~��Gu&7X�2�: 7��Y�L��/�R��o��@jڈ���z��+�>j�Xf�\:�$���Ư "t�"��H�se�qKL�M�0+Y5��걗:A1����&ήe�<��J�r�#x&�/�gvCƥ�{�F�ƕw�j<3�Z^d[dQ�v�;P!�
�P�0�TlP�hdM�}�r�mae-��T+;!��GCe�{�B}��ͣG^<c� jơKsv������I�p�z�q����y���DnN�������1]W��c��ܰ&Hz�@�d�9�.U+�ĩ��}���������.u7�m]}���yu
Srl%7_D�Y�Gj��@6���������o�W�+��K�f;>wLh��l����@.�+ �Hp
����FU��Z�=**�I����y�t
R8>�\c�"����3�ɤV}�@�u/��եL&�L�W"�U�~�w-��p�W,4c�R*���#㥳q��K��[]ϱs���ֻW'Oa�)�H��l��W����iqͩ�>,���ǧ�9����|$JF��-{ݘ�
��Ո��rɎbG�Aaۘ�H8Vz��%��H+O@�9�dJ���wU�p��nt�;�'w1�YY#�I؞�ħ���w�l��<U/����b�m���΂h�.BQ}q�,�ᾫd7 F�B�P�X<'zQ<r�?i����a��՚�#����'����q�U�&;�è�N|��	��;H	�zq]S����0��݉ǂS	gZ�(K���ƜS�I����ٵU��!��D;R;�,��
P9�*DF�4$*�!@��.�Fh�M-1i�o�^Xz��=z!��%^���R�|�*���|�<�E��yeq�s4&�5㫬�k���sw8���eoT1��&%bdr{�*�ǭE�\v�K�!��nF2>��{v�;Ay����c53�����I6�_s� G�s�����E�
"+_��s���z��Pe�r�Ka'�F1�7:���M���.6��̀P�/-K^�P���֙ �t�V�C��@OLR ]sr��ti�|�]�9n���O���F(�m��T��W-��W1�n��p�U�pk�
�x��ӣ�m�$���__E����8E\��[�g�ZV,�����iv�/O4���9u�t��6���.7 �2�;b��n�tz�@�zlχeB�;l���p�<������+�nU|y��ۙ^�K��M�Yxo�΋(c��b�w�T����Xk�s��U�\�f�'����K��w���ش�Hu���f��TGUK=��,���܋���v��SCH��|�`8%Ug����fT+s�*9����.�!��y�:��q��ԥm��F�q#�ya�?M��bDxe-��>�Z=%��Hf����Z���8�J.�D�����М���0T�lǻ����-2C�n�2Ύ���МrG_�Tk�*�2Z<b����cycb]]WܓMB=��MF�&E�ony��o)����Wй"G�<F�챋� gw�ˡ��30��I�{���N,Vmڝ����V[4$��C:�h�_vp�ܞQ,V�U�V���D��e�b@�.��9�ڌg?GO�&4�$�l����n�D[�#!�E��2�Q�g�a��-��k{qn��R�Ә#�r �������X��8�%܁��\[��B$�m�y����kA����~�W��i',���弪�+i@�!�2�z��r�R���<f�jE���8wb����{ ��"X�iV�)WK�uc��xb,T
�<�	�8��FN��;L��[�3u/t�/A2���ǦQF7IyJ|>ՔߥÙCg��Z�/]��?q)�z7l��3G8�Հ�=��qkY#�d?v�?hGL��i�Ku�U~_*qAk�5����V����==< �1���ꃅ�fF7 `�jF����p�u���oq��>Ĝ�;_ɢ6�R϶�=�`P�q��n��P�^�U���Me�i66�^^�c��^���c�2f5���_e�6+�R|z��d��
��1��}���
t�f�.ӹZ� Ib�hQ�\�*��\��Lz[�T�bJ:bF"��bT����&s*����+�\y�
ת5-���b�S�s2@���z-�m݅#�����gbj_p�X3E�'ϴgӆ�ر�˫�@g��L�pĤ+pݍǵ�
OxN��8@׭�cVoEܭ|���|�z*�sG:��'%��N����E�(s7p����z,���Ѩ+���ѐ���-��yX{`]�uX�� �c:N�v����4�Ccp�Jg��+��j���S�9n��U�n�7�[��	ҬNw�aA�4�'O�t5.ͥ�b�jһ%佗/]
(\R�,F��Ybb$2�i�X��Z˾4+�x�R�L	�)a�zuq���7u��U՛�Y׈�l�y��ƋYp���J�n�:�Cs�w[�8�F�F䬸ڹ.sTa\HN�y�t1���8u7	�g
��;0�'S��c@�H��
���NV�ְ(w`���{Olh9Yjnx\���|N���N�h �pתuv#e�/.��a��)��WLR�,��=u����؆Ŝ� ����Y"���ǰ�ׯ+-T��XICB�Z89���a�MX۹}�Φc��]a;0v��V���ey셉�ҁXO��[K]���5z�Y�k�*쵷Im��N��{�1�2�d����n����4�N����]t2�.�g2'X�ƷS@��8s���{-�̦�*��,�^f��t�t�X��;
����b�X�ԧw�VX��R6���������2�˗�vs��]MuxC�i��_I`�<���=p��a���r�[�	�$�C
;��*/;i@ȵ��.�Ȩ4WP�Q��W0��@F�Vͻ�\J��`ҳ #5�߲@e�d�������ۭ�6�U�{��wu�	�Q�㔖��2QU�c�U�Ι��b��h=�ĹL63�JNm�y�C#�`�\z��F��aԈ����`ѷDٻI���:�՞reF�����>mlo`r��_/�)Y&�q��,B�U������j��S=�\��n��CB�1j�����;I7E�$���벝c��i�W�����a��Vy�:�{� a)�&����D�^�4KoE�$�6�h�ھ����ΐ�ϝ^c�=�7��ܫ��f��1f�-�`KE�6��w�`���SM��_Jbjz�O���+.���V�^��\gL18>};vuj��`�X"f�����ݛ
܆��O��եV*�����w(ݳؙ7v�HX榻�E��6.��U�r�T}}/{;��@ �}�(l��� �3_��b�}�U6pY���j���k+HA�uݬWS�4A�yd�rT@u�����rG�o�\��Ҟ���)߬n�H^2�VM�6\z2��4n!E�/�7�v0��	w*2����'�E<}w8:)+hꙉd�/2���_;YV^�X:BN[x1�2b�$Z�6
Ow��LLٺ"�R�v��{ʈ���X.���h�WW��kyr`x�g�V�R�l�⫯ L���������l-1��՘�hQda)$���;UUYE���!$�LB9��s��U(�\t�n�����ݻ�H9�E�ʇt�͎M�P�RW2=����c����r	����!�'���(�8�&8n�wV�V�z%:;Wj��Ա�H��x��ud^�qB��r5����]�*�H��z�D.��½XWq�w<<��������B��Y�"*�J��1Nu���#4J)ML�R�D�˚��-(�ViVQ��̥�ܳ�R!-L�rwR,Tˬ��K���r�]��!9W��r*Y�B+
�*̭�%�Ҕ��:.�ŗ�Z`U���Ne{��	4�0RL(�6r�"D��"���-��"�"TV���;�A�=���Y����sN�J�I,E�j�����'-U �B�OP�E�E���(wGus�nRr�J�Vg��FY�C��;��-�f�J�U�+2�ͩ��de���FS�����7sBg�����|�AW&��v���2�������>�w�)
D���?�< �'���q��+������r���1�j�Da.�'��9��k'�\Z���5dnL�����
ō��a�è�Wz��Lm��
5�s�
2	�O<�Ѩ���w'�u�<J���?`uٷu\c�cw5�h�n�����( �'@$��Ϊ���n�ef�\�ew��,��� 3��ZN�;�rDs7��*�O*�2�S�熭~�f���=P��:XJ���E��Q;�!�n��sc��܌*�ǖEwl�U�͋<�.���+�c�!���khϒ�B �0�e����#��n�%F�m����6�;�|4L,;֢�'��.չ��LC�m��V��t
hq^��B�IX���1�os�)�Iv���A��JK�;c��U�ز��r*,���MD�#���t�Va�]gh�l��S���CRv[�F(@��� �f�7�&��GVDiL�z����5�/޴0�(^�̪�5��IE;���Y����1��s����2��v�:Ւ܎P-�����֪&��e�P��ۜU�;R����v;�Z6`�P+��e��2���{�]�v�?�􊾴��$�)��
��uCƉ��*̴���	�XM\�Gw0�U9G�	5
F�3�*ެ݋j��g5������W�w�x ����l�W!Q��gi�nq�C�˺ u�c���54��W� ���!��y� �\�=Ӱ�����ΠLzn=�/LR�Z��ZKP���������*���*������g(Gt����O�"�X�2�!3�q��Mm�z�.t�_w<#��|�̾*�5���a�����{h,���p�0B����a�����
ĺ50�mY�[5I(!8�ݶ��1���2������yu
Sq&� }[X���7Ln�����qΦ���l���ю�?tj�fӔ�v|��i^,��pF�9U�7�.��i�%����+ڈb='Z�#�����兇���nP��Ӷ2:r�-�N]�3�9�GVm��F��NT�!�����b�'��GK&�'��ߖ*���g�� �y40n�na;Dc�c�K���V���e�|�U�q�ſF\�@X{�Z�KK!�s��\����f�adb�w��ujC,r�J��i��Gi��/��o�`*�p�vD|�s�v5o�^���b)��;��8�Œ���Oa���Vbѐ�ԡq�1��֦�.Ar���Q��ڲ3
��"��d��aE蠤�<;�p�E���mY�v�I�k�j�T�t�ar�������� ��u�{��m��C�Wq�H<�P+h
���*̈�}!t�}2�V��z)P�-��<�׎N�2��X4D�f��o���.X��(X���*-_�!B���C߾&����=�j6v^Ru���.U5���[�.�#3[45u ��J�|�Q:q6���k@�{{��*�!O�?�ž)��'Sf�+��#�S1M8��m�hk�L\+Xf�)��A-�W���_J��.�5>B�?Rx��|S��'2:G��Y��JXWn��2_�q���,��O9V������a�1�]k�h�Tx��(0ɣ������ofOhc��|�xvъ;�^Z�>f���Y�n��=5���`+���vl�8UD�tq�GCw�+殸E�яG�j���V�B�ִ��9^ή�Of�q�5v�pc3S��D1�p����6�6�@B0PQ=�9v�_��=7����|݀��W��>T�{9V&s�ԧy�!#��1�QHP���a]�݉����y6���,����5��j�RBĄ:hq�m��ŊA�Ǹj,��vο1YY��6]�S(�}�{	��]ז���	�������:��x&��g��:�g��~���xə�[�UʁYX���ShǗs�{�D��o�Ǫ�V���|j�R�*zK��}�H�lv;����6�u{�-��7y�ݸ�2���C�z�
"Ȏ���d��@�CI3�W��J�+u�:KU��G݂�����9�J���+N� ���!�������֓��K�a�˶`l.؃������^�X��q
�$r��[ X�]����Ck��B�r�E�/�"R����^oۘh��I'H�i��xnd�/`w)�,��Dg���u�dW�Pe19wYʧ3`��QN��A>8oM�yӟ��ru�F���.q�mH_C/.4�����Fm�nڗ�<)�5\�1�O$}p���p+MGM
�S��s�Ӄ��u�[��VIͼ����V��r:=�J�dM�\�V9���<j����	��u�\*X�M���Í�������-���1���U��!L!��R�TSQZrR��r��U�(�"�p �̢8�����D�&=�-b����m*���VԷ�7ו��mۼ������)�O63]��t���G���Η��N`R�|9ߩ�p�^F�+i��O��"�&���+���>3��Y{��k$�#x/�x�U0U�-"�n
 r��.󌼾�_k�� �9���Z�f�H#�<�� �R�cY���Xu�6ޫf�l�1y�8��(��Pg��͙��h0����.l��d�v�їB2��Y�#�S�T@�Rt��'����|�}��mE3b0E�s��9����ֲ��\�ZFiq;84�e�aw�:؟^�C��cՏkJ�k�Yj��X�P�ܼ�)-S^n�u�RP����I���Q�B����tԷZ���[^���-��tY��#p�L.��9�,ú��TF��eGb��H�GѴ�E�q�%����4�B����QSk'|y,�8��N1��6̡���.0�Þ��æ�T�b��j�H��^y�m]�;��~G��O2��:���!��?a}�r:�����.5Y}"�t1���0QY� %5�K.p�J9>�Wϻk^�����w�ݘH�|~�I�q��#5H�w�OX����f}�X�
QR�xFfm�D�.�-\����FF�6�7�j5pt1-�`��eX�mWo|3�>����D��d�}	���l���c�J�a�yӇ��6y�8EV-K�j���AY�.ى�����.[Q/S`���I䳓�����z���P�WɑVgb�";��t�[i��j҂�]f=6�F��3���-���zM�[F�8$ީ�vؙA�*�dY}Dv��4�dƹ��g+�ִ�m����X��~{�����Tb�e����옎�Wpj�Ӓ���V%�|�b6�3Z��X,K3ˣ&�sW�������6Ԇ��LX��Գ\�S���o+G��Iđ��ĞteZV�V�wnH�޸�Gz��a�mP�
��A6 	��q�������l��Ń��*�j_$WE���=hQ	�X�Q��u�Ʒ|�rE��3
�u�e���"�UX*4T�W�u&tRv�����0��g���B���uf��D���x������gY�sͦ^L����,���I�m�@���dK��V�|����� ��;\� 娘ڊ�}q�^ڼ� ʧ��_��[DP̚�/�"�1	�<���[7��#w�0�qx27B k%a��s�n����[e��
0E$3���=-�)S����a���炄k�]T#/��:�1i�\m�w�jGm����p�����4x�,k�.3�oI���gF���g�Y���g�4���s��c�cE�����Dm�t��6�g�EԺ9�|I�i�p�;v!El���g�϶�a�ϵ-[!���,TL�~�t�tH&�^���57\�ʛ��TE`1���g�Xd_<Ja�(����ŧ�ʃ1��i��&��(;���ѻ��"Ω5I�Û�4�$�[���xx{��[��͠�z�I�lX��2{\��9����)�X���!�/�Ϸ�|�ʼ!9��2�c�{n5R�;Y#���������؂�]�<�����ƿ�.�S�K��7^5C�g'�9(f�JF�d���&�^���8̊zr'r|���%#�Aovs�_h��p8�K��;ݛ�'�trC|{�ygv}��t;7�+�b��_<ue��s&Μr��p�o���_Sp���tĉ� W�Y�wA�z�N0__f8,�����7�V@�o��p��%��i��X��#�p���Ԉ �;�+�8�GZī�oyֵ}�Z�!�Z��Q��|p��=�D*��l���D��"��	=FRj��yv�;0F4�a<"�x8[�o�u��k����g��1-��F�ɝ�/���]�ᠨM�n�% � NҖ��*|rBKeQ�,_;)�F��d�2Fi��O�(�L�e��) ��V�9.9�X�kl醀=g�W��P4��֙�4](�|B2�!�o-��@E�G��΂���;#S.���3��e�+�Ҽ����Xf��-��e\�
��n�3���������=q���?H,E�J�mᗻG����`��k�-�,��[}��&��� �-9ҥ]C�)�r�"7H����/2�w����\^oľڽ|z:o61#/� ��&�xt����1���S�ɧ3�gݶc1/��h3�=���D+��B�q�Ӣm1��UK�,�5޸�Hb�`��U��8Dٌ0duُn�vj��V�+꺈��=2e�=w�����K��U��c5:d��f��HGqa���@JqM�`����j\��#�&ł��oUø����E�|��Md���r�\u�Ƌõ`��020��Eu����z�P���`>1E�����Y�8��H�M���m����q�z㨑e
�3���H���f=ťƿ^KEϻ�zGP��5\ L���>��pݟq=I��s=��������i�I���k�H���	`;S�!�dv;ϵw��������b��b�9�F�<��"�:�8�J^9JdT7L�,�2��\�qȫzy8Ż����S'�b�o8�|����޴zf�>�����d:�wDPRzH�6�RAD�����&��f��O�;�T�r	Xk�W�Þ�`3|\��y@t��HO(l�+tf�o��	{��|���J]�j�p��veYׁ̆6�M�~r�C�x�m� �u�c�*����=#�C	E*Υ�2��@],ʝ�+V�J�mF+t�e�ٔ�yXH̥��dhGj�T;y9��~xx��c��s�Y:`�?.9q7HE}nH��R�j�U`�5$6 ���/k[P�L�fDj��kk�S�j����_��9�J�"�i��U�ǥ�4x�ic3*Ndc��j�2ة�.��h��5�@�����= ��(���U��{�_bߖ�ąr�7(�Nv��	��^kIm�=0����8Ⱦ�;3Θ�}.}2#�O��ӑc���u����3�x팋�R�i��Ӳ��!���$�|��͈L��
�r�L�s'4$��i��*P��4�i� n�^�p;)�[�h
�gA��{$������u�	���<S��Zs���jMU!׶C�l���X�3�nL똸�!��>�ֹu�\��$W/U�i曯#�5"��=g�"��u��p�g��y�j�����񖗴��"�Ył�tW��,�s��?j�+N8s�D�Td�vR��i�/8K�64�.�̙UÈ_Ԣ��nr�=.�i(Xx��ϝ�*����F5���@eG��hљ"�)�C��Un��� �A��f��T�1��j8=��J0}��¼�Q(t-�֝��L=%]�f��I!&�®1pC�憦m��1��̷ܶZ�� )�����ԣ�.��>b��^�|�:�W_v����J�3!��y��<=UG�������!8O���g�׍0�8_آ^��j���J<��N�Oz�`bvH�NV��̛�+�>X-����$h_l�Q	:H�k�#��q8-Ҥ4]��E�Ω���� 2���I��������}�Is�ȧآJJbN����p�'i��b�`�Ο=y�|�8�m��ݹ,l0��	Z�*52ik�BAy��������;&�sgX��&v�a������![����9�V��~�!�A��kW�n#�ԔwFD��<�ts�����Ҽg~*Gc���s� &�o¥�v+�P6�����id���z(���:�j��W�������T1��l@Ӣ�	,vcVZ��5�\:��η�
���p:}W�B�O���ʩ�[���D�<��t�"݄϶�ֲ�"*�=����\h~��=�"Lxe��{���q���W��:���Mއ�u�kks��lv��;��~ꪅJ@�i!F�pҧ�k����K��V�|��66�@��y���h��s����n��u�i2-d�J�zc�δm�$#U�*�v t���Y�7.�,;Oj�% �	��f�%b2UDV\Ւ�WA�Umk�[l�"#�(�7r�y��8����QL鎥��so����O�]oI����^�m��r���MYI�n�o��c��43�_8���]��Xc5A�ڻ��:�����Ɯttqi�is�A���o��&�{�.Y��4��cX�H��3&��=�L�6��T��Q�-p7��p�ZsZ�0��c
j��Ť��	4��Z$1]V�p\�V�p��+v�֬�viЋ͕�ipl����M��c�V�����B<�D�Y�T���
۹�_�U�L˫�$�O��N���AK���c���[�,*�X��ze{��V�[�p:m�/n�;�h�A�����ަv++l���4w:��!0���Ol�7]J�0���<��l�@�Q��U�-�nC즖[�}��	�cw+e*�G^Et�yk.ѓ����]����Ѣ�OTcy���������o���w}\;��hHm���ޠ�I���>�o�Rmq�Hrz��X,�AOgEI����ܭ��P�q7�b;`--մ$���n�bl���2�X��&��s�Vb�k�*�8Z�oQ��v��F�F��+&���X`ڼr��n��c���(�o�R��I�Z$���E��OP���+[���qV#��rX�r�j�Tw5��Ńk�WL��=��.$���C4Z��ܙ(9���%dO��VU�@6�U�t�R�̕�I��;n�T�EVɝg���_}��[�S�Ҳ�1�s��=]�����D�<�1z_��gi�u�n���2̅br]�E˝�ń:�s���K2�{C+7'k���ݷ�%7��;L�y��F�V�n��^��1I��M���>�ʻ鶳[��0i�ґ�v�s�۠z�q6��TK�y����L�]aLr�B��ٗk^i+�5�sN�P���]�.f��P���<֦�"q�W���*d6��#͙��uy�b��}2(`!%���+�Y��T\�gψ�J{�� \�A��/��eu�V���u�[�[eЎ�,j>R��>��h�Ӝ��Y���(k\
n��ެy̢��_Wto5�Z�K°.]�ٔ{2����o�ۼQ�8��s���/������ŚwcoO��H��Krw�j�v��Ȓp�ҭ/����]�r�!,��s�V�{&�p+�f� �B����׷�@GY�\���S���Yǰ�y:�g�gk��тA���<}�����L;�5����0Y�{9�O���d/����\6�!��>�[�V���b���3M�K�B��q���;�{���I��Dbj^;���U���.릺�\�qβ���+]�G'22�N%s�w!$�,����R�4.�^a��8y9b$�IRWwwP�L%,��@��+%�ͩa���5=ĦS�g)]�="�L$1"�T��%���s�7U���繊*	�w=#ғ%5	$Z���K�s�L,���.�Y�Ee*��ݔ囹�z]�3.���l��ܔ�KNG%iӉV�J�����N�[�܊��.t�Lء��\-���E:bD�����)�U26�df&��\�t�*��-(��]��ՙDz�ܚ�g5��0̓�j�]#��H�"R��wq�'<=Bu�NH��FR*fTXE��,�+���R��D��ODWeQ�fA�u]4)V�	f��w#��MY)'��)�*{����}����ϵ�eڧ0�rcs*N�S���y��Eq����P�R�r�*�Q^ǯ�Ï%WT��΅ޘk�Y.�k�����>̛���l.;�P?�j�.U���&����!�$VHi��qKL��"��e��"40�"G<=��������H@�l�e�k/�5�Q��¾�PV:J���5���[c����1��'���l��#�fD]g+L�>u7��#�Vus�-��[0�Ⓤ���S��C���vH|j�X�s�W�����ҙ�ʖ�U{|3�[DG,��A8h=	�d���f��������S�0��# �]���A��ݒ:���������"��ƫ`����֑�o��?ccNϳ�
a�@mʦ��υ���	��#_.���A�5c��ʈ�SC׋�r�2�WzŞ:G_�LsXj�y�B�H��l�|�U�c�ȧ�xާ��Vk�{^�4)ý�Ӥ�Z���t��#�4�E7,�W�%�f�T��A:�Ы���aY�����cP<;���#q��;+kzl��)L�3�O��W}2�QY�����Q+�Z�Ni.j�z�=�*��7�묧<7�p�U���1!@�o,T�Dʬ��^ë���@o��b_&�0o��5���c��2e�*��tFcMrk��0Y��dQ�T�N�*G�����V"��`�K�x�zS��Aq�a/]:LӾ�v�t�T���m�m��R�2В^nwL�M�K:��P���X���\�4�:2�|�Z��G��G�I���Vˋ��w�~C�q�Fk��y�@�
7�Mˮ��%yH��@���jݎJ��)�c�UĞ��Ieד�,�t�xMG�%��KM��=�'���CƢA�7T�2ܼ�OB]�����	(��	�P��!![�R�R���<D_;)�L-��4;��r��v(�=�j!"�K����o�b�^R�Yj�cҺ֑EJ����.3{�V^ff����*b���{l@Ϛ�5���1����{�r0��q�\�˦��N��Xܠ��l�0��i�"wQb�K���E�y]yi���wha� wy�=��4�<U5.�����[;TF�f�L���m�>H:����C^���kwM>�cs���`���dxB`��\����ia���>SqʬPa���2�֡KJ����*y�5"b��.���u�l'{�gV9G};��'�>}��k=G�Z��,�l�}��n{Jk�
5�u� ���0��t>�^^���`���ۺ@=�=���Zr���v��ɷ7)���f0��.�!��j\�um�J����5��`�T�t�1�&���%��
�8�Z%�ύ0��3���{�28��dp�MA^֭e,�2�e����U�v m;V)t�pw8�ՙ߃�����M���}ǽ�vjH��Ѹ�n1�O��s}0�a��c���^g�{Y�7I+u����m�}I��/�ێ�x�'�t�7,��	9��$��觴M�vT���H=�%���q�+[�g��[�o�2N��s��![�>PO�����;�4���s|��p�YaX;�m3��uܫ5�]��8U�~�z�cܹS��(=�p+z�AW=�V)����x�1UHm��d�eƤ�p7�nVu�����˟(ښ�ط�qc�~ɭD����T'�d�f�N�6��	h��f������&���Wl�'n�gn�V�1��Wmq.:1���S�B���u�q�k�7^������k$��m=��Jr���v�#��O�-�Cx1td��uǝVm_>�I��l�<��u��ط9Q�1���d�u��%m)���1�m�E�������Y=��F�Er���w�GPN���U���R� �c)ר!�.u�ϴ�`J5#�fA6���JSDn��-<�ԨF�PZ:u��T��2�MٝYvb�m�Y�y�i��}|1\ͮR��)�۸6�������8���ן˩v�婾�+$=u{�+��үvR��1S��k���Y�q��f���~#Ӆ��cVY[t�𳶱Im*���n�ې��B�쿛��zp�}e����P�t_}U���{ϼ2�l�����N�V�d�Z���F�����;Ջ�*��O���a�4�%r��G��c��qֳ-�oX|��ǩ�ri��P���ʓ��>��6<sc����J[�HY�G����b��*�W���<c;"����b71B���J�א�~�y7^��/r/]��"�o�5B���yave����@����U�-J�ko7�֘�nӛ5Ř�.u�Y4ĭ��i��y*��o�ݩ�q.Za�'��5l����&)S</�/��6��eM�/�P�jVGtNΗl_�7T#o7�,* �Q��"�X���;y��̇���`���9��sʙ����x2}�}iP$JђA�`B]�/�.��lvD��0�Jvymֿ��<Ec�+����0dK��xNq�/cQ#�V����X{â��!y�"�G�����wl'���]���{0��Ou���oT4��- ��Xq�M�r��y�^1�^����%�7��+�+8��]�]%�cP6��y�g���^>D)����W����x�����_^NV/1�'���ӎ;�җ���g����</�?6t�NM�m���Ҭ����b�z����zZ���K���Fߥ���f:�V�ܭ�T=EAڪ�.>y��_O"�stb%$3�+���*���V��=U�W�o�u|���ݍ<�g+T8Zg.ab�d�O:k��U}�M�g4ާ����s���w-����+Z�;U���z�3s]���.n�S�Qy�Y|��F���P����=�8f&�7��'�v糲A�YZ�<� ��į���k�Y�;0]+nx��Ǜ�g_n5"k��#am�Q��Cҗ
����������/5����]!�)�v��=o�Z����xa��[Ĳj�͍S;;h�Q.�-�������C��t*��M�(Ehh+h+�yY��E�v2�Ƙ�Ȩ�ۮ���6��(�7TV����_�O7��*UBP̓�,uѦ������g�����k���݃����;�-��W}a*6�����ΜVH���"+fj�X�o_��v��B�q����U�� �ڏ<q�'�puu*�f�ܣ����v�X�1��Z�z:ἅV�M)F)�k���f��F�u��ZQE�X3�2�r̰�c7�w���i3PU�TD7q1Eqxi�Y��]��`�<�e=�k-��lAr�u|r��Ӽ3ޕ�&M��f�K)ℤ뫦�V��[YO޸�磼�*�'�:�)����2V����m�����gp�z�R�:���e8T�qo�����[�k�zJ�� �,e,P�U���K��P�T�5�����}oQݵ*�N��k�4��<妾�y�?'==�����S=/W�[f�z�)(GE�U�ø����.���O����\+���7du�ǐ�u5}4��3S��;�vwj��#�܇BJ�dm��)�;�Yg�1F���Ñ�-�Jc�;)���egݦ��W<�-�1�y;m�3�	d��U@�n�1|Z�D콈���N�Mꐋ��O!	�ʨ�x�J�����N�s�'�XQ�-\Ԗ-�Q�f{菢#���e�x��|n�TD���,����͍���wО>�D��b�ՇR;�g1~���FҨ=cj%EkY��V.�R�7d�����[o:p�{��R�Y�v�7������:�9Y�����Tǹ�������(w�����cyJkV��Øq�Ҡĥ���PKw]�֥yY���v��-+�v��q��{��X!(�V�"r� ���=�����	;ߋ���dͥ/��a'w�Q���3�6N�P� �W
�8�sA��9�9�Bw�3��ۿ�9��q���u����ˇ\��If9wQj.}�!S)�[fO�\ҵ�W蓾3���=�iV�r ���1���4�+rX�1?t�����c%vMF'�
�`���Mc��6BX���.���=���u�uK<	{�U��V���n�#}�wXu5X��Sՙ�=Ȝ��ӛ��P\Ix�N��˂���w���𞗗y���n��B�)�s�B�-���X�|nҧ'n�U1�{	C+u�]�^���:���6$`'�]��zhH�RQ
ܙ��o���_Z��uUϵ�yEj!�j���v��!^����{���k�An����){��9z�Rڍz����]�]%�}�n��@V�T�2aӺF���x��߅ȏ���/'*1=:�":黎�Z��:�$��C.��ɐz�k:(/�\N���AWL	u�<�h��z)��d�u����c�(�igK�<{.s:��jCiz��kC"ś
���kI:��}�@e=p_iz��#q�܅k��w�Oxw#}ҁ6��;������P^F�t��5��\��ڍM���;{P��&��[oƷ�}*�͵$��o��$�⼴M���Y�G9-�o{uC��	U���9�z��Ukx�zD����Ρ��D�w%q���rh�ǚWe}o��L���u��5k�X���r�OL'P:;*K�����Wы�_l�M-qڬ�!���X�q��	��ƒ7�4Ô�;���t�[���0h浺���kB��E�w��R��.�ʰ����{�_U��{؟�F�S;��x��A�̙}]�z!�"�P?e�}Ir.�[V�g:��&ب;���.���u]�&�H�h�<�T� x =\z}Ӥe{���Ik��>i
�ں��=6�� Wc�q��=l[�̌q��7x�8�p�)�b�☇�B���?#U}�İ���w\��;g�<��jzG<�8su��*7�a`ܩCi�JK�������<[q����=͟�q\���ơ����TC�2��Z�Sʏ��8>��y�2�N�y��ｼ�x�ud�QU��i�x��p��&�� C�f/R*F'�m�yQy���X�'�T��:�n;��7 ����Ρ�j�p6�n?[Yp_���^[�����g�P~ަ�s�w}U�Ø�ؘ��nT�7�)��\vTWQoUἌQ��6f2��"k.�¹\�a�;����ꋲ��Ƿ�ޖ�T���p���A���S��)I��T�u�W%��w�߽�?Cr}�_2	�����q��<�>/4fsl�!;���3���H����mÊnWk��`�9�j�
��s�;�<r;O���A�U���b���v2W6K�z�b�w�+\�e�a�Z�fɖ5�w:Wf��j�4=Ι�j{e��n�p,�G4�?| ���ox�,{|�y��-{D(z�FR��k������چ�G(U��;�yܷJn�.F.�h��+S��ʢ��z�hN�4��>v�E��hW�}�++Pfw	�}�!�=9�9��"�g�?��u���6Ô\S`z�?��ʂ����Z��hYV�T(�!��T_5��9����\��x�Ul�ږ����d�M�e\a���Y���c���NFmkn���9Ϸ���C���q�2b)�4[�VjDjY�Mw��v
���o{qfˀ���ٖ���h�ným�*�݊E�dn�vgZ�Z�\.3�G[�V�Cw{^�-��lbf�
Q�\U��!Ra5=�������p@ןY_[k��,{p�IYɚ�z爼�����ӊ��F&r�k��%&;/��(��.��aW�
��������,r�����ɶ�ܨWFС6����Lb�k����*���,U�h�+���7 t-QIX�4�������v_J�%\u�G�I���B��y����u֖���V��m9ZV.��R�V��7A}�X���w���tWH��Y��̩���&*��DDV.4�qk{%+K7V.M���:Q��]�kj�N=q+����2��V�mF#C%m�dGr��C�5�{Xo���^X����I�Cnﮤ�Е�nc�q�B�Z��s�%�������)���QԖ�jթp���p�д�ڸѻ�0�v�m�U��*��`���Z'$J_85��Y%�4���CN�tw&�5h��f1��WIӂ�2��)��Yj���E�GuU�h �L�yUam��g^���.ꮋQ�8��Γ�T�і���$�Ԛ�r�
O���XG���jt�S������� �a�Wt$��j����M�@̃{ ��n���>n��u�5V%�L���ѥ�����,Ȝ��]Ѯ%���ӯZ�}vvE)���v��eCA�������Cv����z����Wn�v���[�eM��|�",�7���ެ� �(�]����u���&+�u�ej�k-�	�H��B�k��b�����%tH��p�l��=˘U���\ymA�H���r� �SӍWnc�F֞��\E�^8��R�ugt� T�.%�nB]4�L=�L=ʭ-D���w[�Ȍ�'����7Vf��m-�8a��صQ�� Ȗ�������I�M$�aƻ������Y�ejQ���nC�bĸ��f��~���_�j�n	�*^�ڿ ����s��ʰcK���[��W"-4_GdNpL��@�ӱT
鐬^��nt�j���D-��&jjևmK왲]��2�+��wZ���_���{�T�H���$���+	I�stU�RY�zNՄK�:�^Tz(����:�4s=������ZpVVT�=&��2Y��6N+�ڍdܩ�}��/)om����AV�n͏E��!�'!-U�9R�W�pw7���V	��Q䏬��x���ʷ��6���M��\��{V��V��!�2�fK�f*�[D+WY��S	��S��ct;P65�K2:�ơ�^%O�H��x�Wq�F��T��Ȳ�=���,�����P]�i7��ܬᲇl��hdc�(74vU'�իx�gsDG���vbcm�Yź�7�z�t��8T�C��sf�M���۠��<��K]��0��!l�՘����a�Ёb�$�=�{r+�/=���ځV�0�6V�+�NG]�Vnj�捭�fx��/�ҩq����VԴvp}�t�c�. 3�����v�c[V�]mg(�P��wl��D���9\��MeЫ;�%�f���l�K�dYQޱw|�P�-l#V�ic�s���.v��H ���m*^��*�n���a��n����ey.0�إ���p���dY����=�8lSy^r/�P޻�)�ẞ�;�2�D�1R���a����Zb��9��j�diUi��]�=�Gw\(�%hbg�#��%����^�D�f����'*,Աtw1'0�"B�1U*�QT55���ˢPU�����������(�rO)��ʈ��n�t�3�"�B��\D2�萺!8fxyz�E�H��ak5Y��]B��ӭP�\��S�I�N�9�蔑��Э%+ws���IItrp�M:��5-���/tw,u�es�0RT�VZX�V�f�T.�;��I����x���+Wu��J��D�V���NNK��K�r�b�2�(�dB�H�Y�sܰ�
[���l$��,.�(�ж��ŉK3OP��ܪ'�I�J���:��y��4�aR\*���!Z��TN����y9p� �EJ�!�W$ȢN�����"�� �U�lM<�In��:�p����/�W�Tέ�>k�s5^��2�v�9�1+��-4Ok:�������� N�m�;��/�N3������g�K�:�}�u�孈�z��ZX^N�;}��HX����	Sw���hm7�-X�|�C��_V(�1\�t�,a����Q��G^R���s��;մ知�����tS}��r�װ�c��GׂԎN�#����Ӌ����>��%(QR������ꓖ�.����s�����`{f�mKvqe�x��Diy���`��������c�Ƥ-v���;��W�hos�k�m�ߧ.��;�9�zf���)�f��6�[�S[��z�u���������*�S��Y%�e��W&���-��8[���g5�1��9�62������w6wa���7!�.��ҭ�*ZM���Ҕ��0v�5�YS�o���2�x��Z�Ǚ���`YA�z}<�˦W3���{�$^��?u��~!]��P��a\}LU�JP/e��ng(����B���17H���to�H;N�"wu��T0�]�r\n�;,��>%�;B�,���O,U1:{����i΍u<��͓�\$Ѯ�Q�l��嵼s5O��y'��3�J��!6z�z#e���eo�{�{�!�w[Z����WF1zr��za>�]ux��78�-n�
^Y��]�s�[�^W#Ѹ���,�p��0�b�J�xfXW?o>b��p�F���]���R��� n4l���n�ҖD{�*v��x��)ǫz��Y�f�-L섢���W;�Z�w�����m�q8��#��]�^�L�Oo47Z�T(w�M��)&�ps5�/�ﾃ�Sn�+~h��fr�:�Stn���������T�����F��J��Һ���M�h����-�f������_5�DbpnuN�Y���_j�t��)��f�ogv[�]�i#8�j�H���j��_���\t�}�u?�R���c��	U�w�R�Csޮ�r�t2o��0�c�U_lJ���QgF(ŝk�@Ͷ�b��\�j}��C��s�w��������]v;�:]�5�U��v�`_�}W�s{��|�kaG�V�͆fA�A�3�خ�PO�����p}vu�YC�7ģy�#���Q��]�o;OEA�mCCr
s2�VB��鏧8�\��V�^ݎ�ֈ��[�j�^'��6������]�O%D$��d�8B�6��G�y�=�{��^��_�ƚ��}κ�ʇ��㷴�Z܆�d�0_7b�c�)�u���WD}E靕I��z"�q�j�Ρ��}S��˻���aqyک�w�M��g'ܳ�[��Te3��_NĥO���թ�Ko>k�+��p�o���[�����
iᄣc�$���¢�Yx�b�iI����8�"?�Y�O�����<�/��>�0�����i�)����-���X�̲���׋n2'R]���Pk�y���*�v&)J=p�5P!\���V���#�_U�}�ٖ�gؽ'���t�z����_�_!��Ch5��+���*u�=�7ӯ�w�^Dsԧ6m���èO����Y
�����S*���kU����sҹ����^�E,3�<sz�w�*��Ӈ�T���蚪���`ۊѽ����\]K�4�̯��]�	��/�S�jŏ��ft�
��u14V�୺�wIl�&\�`��y���1H�����.��<���z���cr�;�Q��,!f��m�UBk;+��o�{�H�.T(�.ZgG���Wd�6�T%#id�̞lՙ6k���C�˘���M:�q��C���>���Q�͙j���g<��%���������P'�X�.�2!�1]�|��ܚ�;`WU�ޞqj�Or��o>ohz�и�>�+��X���#��W�N�Ʃ#�;��To<zn�}}4�TCX7o���%[�L���c�6��Tb�z�n�/��s��W.ڇ�6�`Z��[=���j%�^b5َ�D�̛T�c�q�E^sN��ې�v����Q����n�d��w�U���_��Ǟ�ֳ�<�,�w��U�<��4���ތ�܅�:�;Ϯ%�{m���ң��;ѱO�k|�;�v�i�͋;��rp2��ݰ�Sx����an(Sã�����^ў�An�zv�[<^�[�Z���{̼oxӍ����M�q�>��g�~s�Z#(��ěN�0gt�޿v��xol��O��O��o8+�1N��啂���h��{G3�HX�s|Fs��0�p8U��	��.�=�����@�*����tRYG7�M�}�1o�Uy����(ʁ����\���]6�D�j���
���%g+�\��*->���dg6�=�}S�/�
9l��# �v�N�jb[�)m	��O�{��~x^p�>t��X�*��j�5}���������S�9�@�[�[=��7�s6O\�#�hQ�9�q�~�i��$j���x{kޛ����򤒒��.Hwe���͸�,��+��d�0��,l��M�G=����S'xu>�����s�elm��f�����-�X��p��W�%m�O�b����%����v�f�uWz��(��.�Jξ��_C{��-��'�F�b7\O�-�%��66����o7n:��9���l����a+�c٩}�U��bzk�Q�*7�=憽��oA��і�6���Y^
��5Q�4�n��^�~��gV����U���5����3%K�[J@b����6ӠM���Ë���]S��-�z� l�6jeH���sG�2���v��ۆ���ݩ������a
�s���a��\�F�,��Gvn8�T��L�Й"��c8���Yd�.5kr$���*:ɻm�T��`� �f���-��]�'	OUp5�l�zy��h�-,��aʵݘ\!E@�`���3�4fs��i�͞����O���U��^�7َ�t�j&Ӧ����OݰK�CJ*���V\.a��7��^Cx[ؕCd�us��{���[��O���ce��j��W�<�p�nz���6�p꾹Q{}2ƽ�ز��ކ>q���f����4խJ޴V�f?����"�_t��T�7���Qx�B��$�-����*��;I�7��`��5 [@K{�a����S�0�T#VTOL'՟�x�R�5kvC���ز����{RU�;8����b~�(�yC]pad�W+^X}�l�N��R�ۡ�onn[��y=ٜ�ˤd�%ƾC�Z<����g�r)Mh�M�86�F�g��W0��ˇ��uBa�KT��e�٥��ZW:Ր&�w-��R3����~��*�������t�0�r�>=����G}����%���I���ՠ�bs�Wn�]%�43a��Y���Yx�yBx�qJj�!�C��Tf�݊�B��J�4(3���/6COe�ɉ7d�u�LY�V,k�9��B�{�uq���f6��K:�	{������F�͊!�ڐF*��Dv҂wab�>��):Ͱ�ٙ��+�̷B]q����=��0�4n�1�����P�U���  \t:=� �+�o �������+�y���,4~�s��	�K-}��}x����g|��z4�����=\���Sj��b�z�Ƒ�_v>�(<����@Ty��ک�7�C3|տq���q�8���'j�Jj^��Nm��J����T��M��}e�m��7��Chg})��;����笜J�A�qŪ���5N�ڛ~}溫��j�6#���Cγ� �5Sx���{����	�q�W�y�ק9�ޔ�"5�ݔ��*�EF���0��;\��k_��2-�� ��`?9��g���~�>����x�n�m��c1�Zq5ݕ��0����H�Ć�zF_��r:#�}5xlx}}�
a�'tpk>O1��9x��i���r�6�}ˠF�S�?p����R���'NG4�s�51|�H�����B�P�%3����Mә��x��ܻ����=�*=��O����@�4�,��]��<�`��{�Y�#wh�P��s\
�3���H��īk��4J��c��[bp��c6��\��VUԎ�m�t�zwB	��%^�;BL�K�v��lp���J�����P�t{`w�<<=�?-،�����Fm߾�ʗs�s��,c�{����<*�t��5 }����"�Θj��=��Y�\�0�>�p��\u7q�@�U����ͫ�i����j�:�����{pme�[O��5����˕i���7ձ��h,���q��m^f�CT
�,	��Y�Pi�孋�g8��]������hdk˺�{���!��@ڎr��s�����n ﲢ�^NV/�4��{'sj�bJ�W{M%;+�8��/:�����ܨ.;(⺈��璦�4���=��u�8������_�]8����wS��{bڱ����M��bӜ��g.���y
�e�T�kf�ZQ^Wۉ
Y�w����m|��n�	�}|�o��Z�B�4��ʝS��+����79�;����;ݍ�_3Q�z��	�c�*�y���Nz����{�A��O����]���j�{��('�͓��[)��r�O2A;��� �ooU\�����)lxp
�!H,i���6&I.��\)uq<�y�pc	O����hQ��@�C:��w���{������յZ�_'���_R3.AV�8e�����89t�ݵ��{��#����f6P�Y��[BB�o����2SnAy���ۓ�uj����c������-E�
�k�i����'��T��L=���tq���jm���\�������si^����-�w��W��в���-k*�4�oC�_µs@W8�ǃTyg��"�hV�t�|Ԣ�� �n��C�vzn/�}�Q	��Fve>�
�u
�8����z:��S���r�P��P��>�"S���<��2�'�a\�2�9�ul�88+ܸ���x:�\2?=⇾X�k��gE���ͬ���]�c=��\�ͼ����y�,��MW5���
b�����47��K��FS��/]񏥜�Ƿ@��p����n�Zpz��8� zXx�G^^ܟ�G]�i(��yA����ovV=Kk^��/����\TcCk���o�I���@yh^Ou��Z_q�`�ٛ�����o�}��/X���I�㕈-��M�4u��q�\x�dv��,��l�:�e��,31�f��aPb����.D���t��7O]5�+�L���ۖ�<���fR���燇�,��í����m��;��c���Wy�}P��_9�C}�_\����\g�3��7Z��c��@����髨�z�����}g����|^�1��8�\�TE�ƭ����?m��=�^uK�v���Gv�Y�I��ݨ;ڧPA��C�Ȇ���_ϩ���"ڮ��}
�V���Oo56kD���x����8��{��{��^��q��wΰ��Qx�y設t�>��	7��_1h|w6���=:)�����6�j-_+Sp�����վ:��d��{Mz�V7G�}8�����"��2�Z�n�ɫhJݽ���=�V 0ji��Bʉ.`�¢�<��ܱ)uCq�'QZ��n6����Ku\�pS�V@��F�S�0밻/��g�mS��Q�U��j�����5�q��݉�R�T5p�y�p2��ُ�أ*��E^a;K����9��I�����6֦X6k�6��ʧ�X�6�C���J��]�/�NMއ�n־7vڑx�so��7u'd�i+�[ֈ-��$ּͨE�E���g�j�on�T,�#[�ڛ�K��j��1�+/A��ޭ����YvWt׎�h<kv��.���K�(L��K�y�L�uu�k.�P��`�zGFF%�h��0 ����!�����ž�Q��49bBc��������6�3xm��I5�^su�
�ng�N�Gm�H�Yб7ْ����^f�l�p-ܕ��c��E��@��w�q�ۅ���-�ы�������ka�c�oR|�b��3�.��rwDv�[51����*T5U}��:�-gtk�V�*��3J��K$p���ƪ�1lX��zgU1��le���K�N�v������;�x<d'm��t�\�`�u�	���6N�vpk��_�����<�HQ8�U�R���5X���ɳ2cu������H{jp� �&ޢ�x�!�h�+����(��n`�rU��o��Q�I���+yF3�ci�yH�E����z��m�Vդ���( �6�rE	J=]����Ĳ�i��Ӧ�g��-rD��kD�R��of5,8�D2���NGf+�\v$�U��C�׎�z���>�ս�r��GX����ݻ��WU(�٠��҈nQ�|��#8����U����윴űܭ�er��q���|Y�Z�Ѳi�kP�O���!�-�ܕ.��7B���Ġ��k���Mۛz$��^!{��8�U�޹��]i��\Q�R��9NJ��b��J-�!�����j�,:�n�C�2�9��+�IYϚ�kc�T�m^�y[�t�gL�ge���^�v�����wظ<�pR� �@L���=��jv"<]i��Y�,[�]hV�m^����pc*�:|n
��f��]Y�X��A$;Z��XP3�a���U\�=�_��44�Vu�����̏�&[c�7cu��r���ۊHA��vhƞ�+
"_q��Y�M�׮�̽�#bZ��� ��� �"]X܏�5���〪�u�I�n�ċr|��a�k#u�A�et��ݜz�6ohS�<He�BE�|$�1��ż�Ӑ<�*d)�.�(��|��U�uQ6O��X��*�����F��+��|b�ZL�*�X�I�9�:Y]�a�u��7:�����o'Y��'�Ȼ�H�zr�iM�����EOs`(;�HL�6���4B�vĘ"���e���[�����]��p��-���;�f,yb�y/�9Aj�;ko"]�l�d��|�<�� -�wS	fՆ&-5��K����Q�q��f�����n-��e+`��sP>ݰΕiw+����(]�������.�,7z�_.��|w(�%\w)�$U�E4����Y]"V�[�W�Z��GtJ��f&Uu��*EYr�iI���Qk,��@�f`�r�Uw]P�u�
)�gµ̯0U*R�!up��:�"��]R�i�)f�����/\r�U!3IgMf�Tu$�*3%�p疹9�f�UQ��M��UDg+	9QeaAQ���u"��(���Y�h��zjp��뙗4Ғ�2�+R"2�p�"9ZӔV�VK5,R�Y��^��J��S5#B�B�B��i�
*�L�*���ԋ2�����r4����,��xZ	=<ܮF���	��ud�,�*��-AqE�*�q�\����052��"�n���E��U����qK U�:f���%S����t2���E*-H$�C�H������]��:
g_oN��1�<���7	���X1��\��PY��t�;*��\6��|5u�V�@%�}_UR�ǩ�{=$���s�o�!��n�M&"~�]�me[�:�r:W�z��t��[�y3]ٌ+�ޠ�9|��Uà�%�g����4ӭ4y��L�۫z�\F�;Zw�x�ד�AT.���OB�:�RU�� �tJ)��x�]�����TR���=�Z�&�S��\V46�Nuwh�ȭ<�@�w����F��}[l�G=|����_{��ؽ�j/y��k��6�c�-)�]��d�v�w�M�u�UF����(������ʾ�h!5P���ݰ��A����i��k��r�~�]�7*��z�H8\ǇS��<�'�yV�B�b{��5��}��f��v4-����ȱРM�{�nq�Ϋ/����[܇ɭ�nT�����v�pS���ɽY��������{~"v���;ȯN�W���2�zAKQ^�C]>�륬�#�W�;h�]�׷h� ������y���E��/H��F"+*��@p�O����Ǖ9|�e'�kp�њ ;ؒY0թ�nK��ę㪳�hz�4D#橗�
�q�u�n�4�"!�;;��W��WX�>�U�Y�����kypN��}�Rn~�L�|2|�� ?9���J��d�Ţ�s��a�(����������R 6ÄSn�@\���MCc�5�}�xLN_t�cϟq������,�oq��Ȥ7}�4�������y��8�[���Y�9�n�s�R����\�c!YG�������Ը T۪��.��ϵ���ّ�N���6�G�zt�����n�u�JY��Urj�t�|��gk��ɮV��y��n��U5Ct��$�+��fkb�=���(u �A}�V�ׁO���رΫ��*�3F^P�����:&��(�F�o*ss�]�?$�ˊ��y_^b��q`9�&���`n�o�gPͦ��/:e9Π�i�!+�_<��=뫷Vos����;�2l���c۠\v��M����ڇ�R݋|_Aq�Pq\�����WZ�Y9,��F�1�WgQƀ�YG
��H�Z���u)�!Y��ګ��	�m�C����ze>�Լe8��E�pz�x3@'k4�`C3��kH����j�We�\�8/�Ղ���"�liz��5ү�Zwx�DjN�oK�opR��u�7��MIM�w����۫�֍��wNTFtb�Pb:�F�ǣ�j���5�h���.��L��M�%��dNI�Z�b8q{O=��u.ߘ�ֺQw��6@�'����~4�����CJ�9[��d7z��n�Է?_R�����vɉ������z5]��qyd���ԅ��m�G�楛L���?V�DN7����ꓲ-��y�Y���kW�}�����6�_p�E�����0�H�H��]�U�2����ټ�8���*���k��#ۭ���T �3nc}Ǧ���yÒq�_����玧�W�od�M��m����ns���F�ĝH�х���\]���~]2�M����<����#��b��b���-j�Ә꣼#y��YS�]`]�as�����g���tj�/[���}ܳo���:��9f)�k�<�2����;,^r�蓩L��
�zc^}�V��1����B�%5b�X2���ܹ;W'8]Y�9�YyS��K�޷"�3���\V܍�L�ؤV2K9!�[�v�
�q{{��kF:����կx���p�����t�SNf�@���\}�琭�X� Wf��������3���Ef�	��s��__-��nm꡴�U}8}pUÅ1m1�%�	Wט����b��<鼳����^惉f�P�K���h��vI}�����d���]۪�r#/IvqOw��4g����]F�'�_T�V�S�[��F�,����\4�`c�2�k_�!�|qݽ]y9X���P~������*�5Lf����3
�'&}�2��[w�҂�B��u/m?R��WM����Q��%fcLGl���G.ʇ�6��[w�md�Q��ם.��,����)�l�qX�.�)�{��5�[p�R�	�j��k�2�Ku�˱�N��^S|��q��^�U���Z�]��'�]z�k/�h�����p��
k)֤��Z��p�m����_z��ȶIH�J��dr���:u�j�f�s��m^̱X�[̔���M,U|�S��ܧ�2g[��uyo��m�e��Y�	�X��x�8���,�
�Q3��*/y�}WU���=�qVd/����Rs�㻆��-N0�R���B��/?}� ,ϖ�g��9D>��C��}���l��cv��on�;*�ï���Q�YO�P��}{>�C���p�����t|��P��o:g�ܨ3L'�A����������;c'�T�Crʸ�0�凍���������S��Z�-h�,�����	Mb���K�Oх���l�r&��9�e�f짽ە7�e�G7���S�������5u���Ҝ��R��y��篱>Κ��[�������C�s�^Ŷ�
��օ���
�`j��+=�=��ڵ�c9�ד�����6���6��Gn�l���ܯ` ���>ۃo*�E��ՠ*�K��.]M��kn��gq�ߪ��1p)����j��v�X�w��}Y�	��l��lT=�r�:��l�\2a幯����u��B�����_�� q�Q�4cNyGܷH�.�v<���Q�=�f[���ΐ�$��
��#o����*㞛�Xo2	�"u<+u�1�q3I�!q�ua�<�P��I9��˳��G�Z�zF��=W>ld��_}��<`���/X��X������eß�}_^k���.��Q���x�7��}}5��M��n�)&�f��ة���&�y�S�#�U�1�iyQ��X�gD;�n�5�S��N�Q�~�.��u�"��mS�ٵJ���wڧkS{p�ې���{�ZȱanH��Z�Z��z��q��'Z��l룜ք���y�m�Q�����4�M&����z;*%E��a�Ȇ�}>_�4����vO���R*wܶA�$�״���\�m�'"���L�*Vೞ��J;����Ͷ���w5�n�����C�$�E�G�9k�u�f5ѵ�j�>�0�v6�2g���.��w��|��K��*�b~�(��w�S�[ܻ�3�Z���Ŭ'�e�ٗ9�I<r�jp��6'�Ҏ����ap�0\�ݰUpv�0����V��'�p�o0����u{,���m�a��إ��bw�)��5\����kZWfl����	�
#�(+3^�zFcW��H���6�����;o`d\�_RŽ�Eظ#�ojb8C�*bc��]u�d��C$ Wj;�:)z�uX��Kf�Ԑھ�v���e��,��Ui5Z(�ݡ�P�r>ͩ���g��:H�c\8�=�޸���<]��^����;�';����v�L�u1�j'��ҝEn��Pz�Nq�L,��4�ʼ�Qx��������f*j�o8:�]��]�@چ�����%�}�w�Q��{�SC����^j���k]2{7�x��Sv��q�t��Oh������X$m����T����am�Z��Ծ�/'1Ž�Qus�����6����5k2N�Yঝn�vΝc��PTW�qq�ƺ�[*�R-��$�/w���{z�6�(ie��=H�-�ͽ��3��}S�������ݡp�B'Y�.�>�zA����N��|�8d6]q�@{�[�?�Hz`��tsx\��Q�(����t{�>�>��¹�U;�����/���w�뤰�\�w�n޿�w�5�wŬ���n�ͽ���|(,��
�Gat[��߱�z�1:�{}�H�X�j�*��ُ���6���
�޵n���d�P�[�
��a�����jR)e��˺��ٻ�ls�°�(gX}.�"��������/hYL��c71:n��Q��h�o6'2�]�T!/S��m��!e��39�{���[m.ݷ�?�����t����G6��aH�ѽ�g��a�Ɗ]�E���˫z9���)��=�b�����M�OI=�/��,�le�W ��U3����0��ï��U5eOL����2����r���e�j�3�ެ��W9ݬ�V�S�a^�E�����y�V���<ˀ��讵mj�LƉ_)U0��V���Š�2Gl7qJY�ev�Y_[�)�sq�q���}�ܿ|:*�l^�w�@whGA���NT��.n`�a���7TUk��UK�l����x�����ATB�.�Pu�o`+_��h�C]N�T��'G�Xq+qx�6��=���]F���+���Oͪ��=��yʈ���F��Eh��]#��㺷��'+�OMF�~h�}�����G��2?������}{���J�~V����hz��ڎ)�Z+��C
G�o�(-���=<<��Wt'��n��帻�oh��LPH͛α��m�W}P!Bn��m���.n�=��P�����Bț��W�2X�T�ͅ�Ui���!N��63t��%Fu�J���|���\T��j�s��k����s�'m�r��m��qv���c���f��i�l�of�qǲ���x�g;�n�l|��v�V�q����vf�����nP87�][�-TY�z��-妟n;{JU��y���Jc{e��5���>[w��7%tR�#'��\x�yp�v6�zk����#Z��W��Ⱦ��¶��8uy.%(�|�.�V��-+�wu<���������q/�T�lHi��%�K�E�yb�ŝ2��U�[���0i7�yU���[�?K�i�E�a
m��]G��|��m��pߦcm��8���w���U��1������+���[QS��{3Sۤ��M\��%�Y���*��s.�*��Y�)d��Nr��i�o0;W=[=��ܼOv¹�ޠ�9}�{p���J~7YN�+6�'�b��� xa��AU���v�����P���������i<L����V>�3����"���~s&
�{��ĶVDi��֟�02qxAО�P�z�>���[qj��K_n;Pnm��޾��$���}Q��Wb�N�y_6�8�ʻ]�r�����:��A3U�#��g����у��'��o-��0�/f��m���i���;��p5tM]����Qwa�a����ʼ�x�щ�WnDk�"�ӫՓ�]���R�@#��P��9���g}.���B�.ߊĻ�N{�z��}���>Q��9����m��5��ޯ{�۽��B�pzZ��8a�v�=�Y����gTk���o�����ӱpm|�ۂ��E�����*����R�[��t������-�q!_%���}��]��G>�Y%8�؛��W~~g�p�W�7EFo���Dzq�������ې��vԴ\�Dog[*�>B�<�6"p�E�vFAy�B�{r���}�<t�*fj7,M�p�3�&�8���������� �d�<~rm�jqb�{%SQ[oi��;o��x�n�Y�i��a+�0�tu�0R�}�6���M��%m7�ڵi��g��s
�tY�17A0B�+T��1`������pdR��nZ;�c�Ƞ��W�����e3f�D�e�3�DH2gZ:��dH��a�T=��[�Z#$U��u�Ƚ�-�w@�AUm�ԓ��Z�r�,���I��ޝ�	YV޽�MCۣR�	s,�8���+r_�BX%���f\��U�1�w���Da����.n�nWq�J�&^�l]T�M��P�Q%a�YGQ�Oo@c]:V��8��cjr���O���5����L<�A�X]u_wo��6ҩ�m�
 I":4�Ft�gdܹ���e�bp��������ʕ[�z�3�ΒQH�Pf��#��,>�R�'�h��nf��I��wO�L�:��h�(1J]�a��\��{}6�N�+ܨԃ�P�a�׫b)&gVq e=>읏o#�Z'O�68(��R�L�0�Ffά����	���M�|�X}wkN}}�Q˚���o��C^��gI��£\�v�n���*2���J��c��m0hݲ�2�dݴ���
��%y�NO!P=TFK�y}��tX�%K3L��;T	v{ef�ymʒ���j5c���d;�����UcTݛ���z�w�}$�@W|v�kX��a��Hգ���0��^v�kiU��'q(&����[�+u-ȄK0�1GD;)�[�
= �
�����7�� ���\*�B:�u�by�$d
cF�v���Y|̫['>�L�@\�d��@���A�=�ҧ�[7������1��i�"�r��}�w�w+�3k.S|XO/��#`]�v;Kt��K�hŢm���c�;r>�f����!���Ͷ�6��'w��1�q>JNF+�-Y����D���O�.�\O:�&�eeJF���a��w�БQj�@�,����KR�Y��˹,�]81*&�e��j����s����]����%����Tة�Íx������BI����z#�]mG��m��{2��V����K���#��q���q��ފ�ش�8�g�5};\���k�B��}t9T6]1!~*m��0�ѝ��;�͡���QU�(��܂N+�x79c	�T��u�*�0�WGb���j�$�2�!��d�@�H�-�R��ُn�5��ev,�	\�Tw��g=0:É:(�{����qu���X�N����؇��;T�f0Sl^�݀R�8�urA��L8-f�G:���\�G\]�H�Ԭ+�@�u�(�zmљm����d�6�Վ��Z7�������9�K�y�e��O�+J��x�G���/^<.���W�J�SSA{��mmlD�Pc�K*�#4t@oz6���AM=�!�|��#��ΰ�{#(O�x(&��ֵ�W)��s=ނ����҇v�N��gs�ʓ�Le�bm�le�pAv�q8�@�ˮ�}��i6��8G
2F��@��k�)U��k5��׵UQr���W�i�d����VȦD��wIC$*�eT�r�qSS�/E�˔���+�q��J�4CF�'4TB�C�\x��)ʊ��DG:jV�R"TVa�KT�":tT*�7�wB�B��5ա�iRir4PU,D��Fͫ<�$��#-2�M��l�B5rC�Q:U�&[HLˤy�x��c�R��Z��#�(�T���Y�L0�
�s(t�¨������"$��^IlYa<X���V&H�Tmg8�
�Z�]2���E�l������D�N�ux�z;��S��u�(����M5Q5����^�.I���xO	R�����TX�IiQӋs�+��3,�%u�(�C����(i���E��7;�)���
ώ���;�����<��|$��) $@ 1�x�v���u�i96� 
�qX��zP*��R�CD7������eUE�Zņ�mT���a���uzc�x*�f�$[�����lx�iTc�k\�\��e|�Ԙ��Ի;�U�ɞm.<�{�nV��3zA�k��_c�V�e)G��K��f��?�d?t\�Ms.���PI�!����tG���9T��͸UaJ���+�Vcj��C}�&C��>�%nM���\�0��a�D�q����':�dbg.:�\LE*g��}�me}x��8��F���w�g���T���5���v����m�Z��$�̓O*/1TE�=�&�1�[�ՂT��7kj�ŭ���������C��������^1�c.�g*��ȯ�54���4�y�s`��{�e/Pr�\q�kCi�ۧWy���ܭq(��_�S�ݦ�T;����V-�z���Q���z_N���*�atg&���!%wWמ�y_��(�k8�]��WQ�ǖ�]׿r^l@f{]�ud��t+�;��$S����\�ם)�[˅����n>�>��@<״�L��x�e
i���T��i/yqU֔���w��]wx��b���[�2zr�Y��[���D���=-%��\�K
w%t�d����V�/�:�0��9\cX�>\/�{ҧT��W�;�3�y��#O<��Ug[�UmD4�pVJ�C"�D�e��U��v:�<��-�E�B���Y��v3Ŋg�w�&��}���-�i�v���dި]P�'���-�:����(3|�ܷ���@כs�%����-_}�oV�O�ۊ�Q����c�]]�}��<��rr~��¢�,����Qͥz�n1�Kt�h�2����row67R�@e�b58*LkՐ;��R���u@o4*Z�8����3��v��59�j�EЇ�Hz�fU��5}7���֣B��W}B�p�K��η����:�<�V�M)F���<��b%ne�O0��l��jI��P����ni����4[�V��lR������r�]o��ķ;���Y.�[p:���.�3M�{�\:
�Z��~��k��8Oq׹�b���4�(�2\�W,����w��a`げN��R�Ei�|�cu�y`���Q�J���F1mVF��2 ��!�F�����7[E�S%YJ��̱��:vh�X��_�4�vٹ��Vn�z���v:�-iŀ�؜�PU�����A=�()�-�-ng���������ڈ��Q�u�;��Sv�K�Ɔ�>�y��*o�~�;��I�g����{�mnϺ�@�AĦi����۶���@.�.��	�M|�\�^���@�k�Q��5Խ¶BT����q�|�a8�݉V�l�}�WK��%���&؞G 馲��յ�|�i�C���/:w�͉�|��;ݧ.��s�����d\�� ��Ǹ��^w^��?�Q�ɖ���T�x���^G�=��.iTf��g�B���j<5�-��INr]&a�D���UpSȁW�L������c#�?g��|{#ޯW�9�GNɵ�`m�w{FQScS��}�nj	��
�+��}P�y����XT7V!)�ܛ���+lC�oк�Нz��,�% p%��n�7-nF�4_��� k��@h���Ӱ{���o0�Hlw%��%|���͝ju)�=��+sՐt�-��6ۊA5�a��f�>]��ص����\�]�q@���h�1@�WL�/`��D <�J:)�7E�N��:w۸�7�0��H�����UWh�Q��]k��um�_�%�����_E��ȿz��^}�@l�)��23����\T��Gz�T�j����R�!<W��k��Wr���}9ģ��/=tFź�$�8�2�ba���n<�㼜��^v�X_g/��]����l�և�=T��}��2W� ~��qnk�@�#C'�0�(�����{�uo)MVѿ���ݑ����VK��׍�_�{��`4sS���{>�$f��{z>�hS���#�9P�'p���WI�������Er�L[US㛦���9��j6Mx^=T1�F��(�ϫ�v��7��6}���&j6���.=���M�I�v�8�yt�w�z9�q�Ƴ�eT{��8|�(�}>�����Ng'&�C��3�-�o��h�3�P+�؄���'S���n�U��gM��{I�3gi����tf�m����QxNF���j5s��^�O�O���~�߼�d;]3�?��W��mdNI��Îߪ�ed֔0���r�����l��O��=�ï�{-�}���
2c���%JTP0M�H~�!_u�;��U�{D�����=չX�7�&�Uڧ��~�r͋u�;��3.M�V�Y��͠6E��;��4��E�*n�]��|N�7]NҼ�$3��g!,���Rm�L!�V�j����xn�V���%w߄��=�$5�OƱ]1��=3��GS�|�~�y'~eTK�ꊿs뼽;��R�bPX�e��}BP���R7&�SsP������S6K��\<��D��*,V�+y���7��Y�˧�)lG��8\:�ld)�,�}�P����`LSwϓ�T!0V�mk��:���=����O�Ȣ�M��Zo�����Ы�ul��5��*�z�u�y�т�L�z�v�w��>S����ς�x��[~��gz&w�a�[�y��,dlĶF�]:Y
~Y��t�þz�=�o��h��V>���ς�jЛ��x���H������ �w���wj�"�xݍ>�o���~��1/����H�����8KGw K���#��W��H~S���_�*��ؓUٴ��R��ѽ�W�~�nĨ��ÿ_�����7���݂a�^�/��z+%ޑ`Jw=����i����徚��*b��7<NL�>�3a���!ߧd�F���p��4>y4&v܏k�h�Q�>�Q�޹��9�T����Qgļ�>�Mφ�Fmhqn;=���2E/U�G-,P=�����pK|�5�����lE�X��o����GI�S{�w�����b��'*���y�C�9����W<��Ժjо(cp�"�5��F��]��,͍��*w`�hV���,��]�p���y7��y����W�Z8���+��|ꏦ/����w��yen��zrO����|d�n(fX���{^�^R�����ZoT�f�i�<��W{ gz���mX��{l�w0{��=�.��ފ�����$3���C��2�3L��@�.����@^����*�����"k<$㻻ˣ��P���׽��;'0�Ȫ���+jzz�27�uH�����&⾲���7Nx.�n_��A_��Z<�J	��g��zn��Wp�2g}7��"�.++M�my�I�U4����%~�����ct����G��Ac�����늦����޵]5^���zg��O9>�ُ)��=�!����_���>������YE{ J>� -�r�R��`�����ՙ�f4���dޑex��}R����d#>gFo�Wq���C�׏�ƸMu���c<�T1�ԟ�Ch�
��T�'�(�¼^����ւ����}�{5�c��;��;��ޣ�&t�0����GQ�*����CspO@{uR���Xs�Z>͘iC��,E�ϸ���ҍ�1I��]�crݸ�,C��^`y~���n�<�/G�Ի%��A���B�/*�=XV, �s��z�5P�����b��;}����ߠ 6�۸��rF�d�k�r��j��ڶ�86��H��#z�N�ל�P�����+N�S�̃���)�A]J+bziAH%kp/p;�j��~�R6#ޯ���9_{7��G��{A-��L?���I7dw�=驼X��J��O�W[�q�<
�z� ��DS�rB�:-���j���=�}tе��O�o������>�w/x�z�U2�>���y@+�{,
�w^�������9Ll��3\2�י�[�[,��O#"�N���Y�z��s��'��e�T@w@Ty�zK��Y�ְo�W�Չ�F�H驇�9�},t��:����VK�\_��=7sC|��h���;*7=\�`&A�*ʒ��z��q��a�f׸�zx��`	J�~���~�8ޘ�ا޼���~B�uʿ�D�I	�����f��k�+���xg�|1�. ^�+ۯe���_��Aׁ���v��<R�:}�κ�{�+E�y�=��4�,^�V�+��̆��"��oz�ﯖz�j}.X�~�:�7��>��G�ȗj�r!{o�ȇ�Gi���=2���W0oݶ��q/gG��yL��_��/M��~�~�~=�c�=���w�[e�	l��ft���^�Z"Q�K��.��_�&�x;�.���=�aK����V5:�f���5�`�ڸ��{��nTT�wj+�n�b�2Ԋ��z���s���ÆCH�v���qree���J��e	=�l.
�_k���&��,=Gvr��uƥ�vC�q�D�׸��X�s�,\d���FL�����:y:�=�s��z�d9��g�����U�b=ʲ;�L/}ފ�o�6����D���^mT/_ǩ�c:_�Fo�_;�T>���/�|��}�ԏP�C��<2=8�g��7��[qP�SrZ���f)���Ѽ�{[맫ގ��n��f�%�^	ly_�W�����+`��(�AϢ[���!z��:�NEɍ캻TM��o�8��+��u�H�!�o�tU����W�w��� s9�R�Q�}9g��z��jZ�_��������o�c��x��Q^~���n�_�e���r��&�G=>Z'm�r�g=�B�:�g�S���9�_r���L���>�^�ȟN@W�\���-z=u�J�m��@�*�{"n�nO���)��:φ�	c7�Y,w��^7ʇ�>���;��2���W���H���p|��XU���?a��4��^_�`�Sc���xh�BX���
;ޡ������������E������{>������I��'��w�{e��k�_���nɠL
+�[��-���'���&.���jcGF�W \�*��s�[ѝ��Upk�X�*#L;���x��v�݃U5���a^�U������'��r�5eX�w�`�Ռ�tb���l�4�v5�����>9�2m��j
��;�$��웕J��$�8�}�2�ϩ��Y����wq�`��}���Zn'e���h}��~Sy�7��k��J��ܩ�;�xx���bs]���Ҿ�n�U��gM��Ӣ��(k�z=�xC��s�������Y�FO�i���7�|X_-y�e{}<�u�TG�TO���̣��v��s�h�>��u̱{5��	��\����{{i�C�>Ӯ�F�����7|t��\6(߶�a�|��[e��)�E�=�UƱ]1q�:��ςy�S�|�~�*��쐉x���A���'��{�����1�}�H,��)��&�Sq5
�T=�2��ɖ�w����	��s��~X�_�Om,>�L���:Z���{#ޠ)�@-�������΃�5�:�z��Z�^�wd��SC�����q�G����{�F�_��_���^i�7HS٬�/=��z�����o/��9��oy<��acξ����3�:����~�[�y9NO���~��c"k7WEos�B��>�ٞ����2�mFς��	�u�({�(�o�u]��j3j�˨���{�l�]R��y0&�E	X�-v(�:����ާ!�t�&:a)Z���3�k���ة���jAN]=�e閖G�N�DJ�}��� ��bF~D7����t��{RRnؓe��J������v�by�Ż1�*�����]�/A����Q�>d@��g�����"	h��	cԝ$|1ם���#ދ�������V�^�o��@����&�x����ñ~�v��i~=�&�ѵg�}w�[��V�C]V�:��tG��[�\�rj�d���f��;'m�S�M�50��z|o�����CS�7����=������{>��o�|Kˈ������D�zw#�=}�y.�k���P�l�i���ǫ�fC�2}0�|�zg��6o�Ė^��ȹ~¼F�;?b��U^�:T��s��:+N���`/�f{c�[�쁑�������V�{w��Eʙ�@v,�+��h�b"V�I�v���yy^��i�8��YV����' p�7$g�O�>�_�������|(\.�Z/��Wqϧ�0�Ȫ������z���5�T�����iݻۯl�V�)�>��Wx���¸N��p��Zd��3�M�EV+�w3���}i7���U����z�O'Frt��#�/�v�.;����]��S�{h�4������`�Όi�\��zPi?�vpd�.Ʃ���T�hv��Z�#5�q3yd��++e�u\*$�ׅpZ�f�7K鬫#]4��Zn@�].j��q�P�� �s�SN��l� ^#f���qk�����\Ҵ����^��bu�ݏ�S��	�ؽƷu����J�ĈN�5м�[J[�411�ù����"�+fM�f,܁r�p�5�i�Ū��[���dyo3��l�����CyW�8�,���[m>�ǫ',Kܜe�^�%#�#7�[ˁծ�I�,T6m��7�y}�I�T
P�W�� m����0@r�XY|p��,�B8�*�Q|��qq'T�
���w:WKu�����5ch�������\V�Q��sk�;�S�L���ܹ]�M�l�N��x���'�H�� �{m�"��X��1��k��5�U�;�έ��r��̥�-��]I�o�Ÿ��:m�j�����c�ב`����'H��%ȷhn�mc���8ay˾�х(�μ��"�
���6�������SB�[83��2I��QnVw��K��j���D㢘C��	��o��j�b�T�_p�yu�~�6+��������G��ޗw�|F����� �(ǚ5�Z0��*�ڌ�F���t�u���cd���R�3��6v��:驋�� �g0�lI�
��Y�ʬs�sU�Bټ3#Q����"ї��ںM��9��Lv=��_7߰� |�h�X�n:AbA�E"�Y�r�9����׀vv�h%�l�m����Lћ�� ټ�Z$���{O�L�6�e�񷃅�ЅĢ��"�)�̵@�o���}�V���نI+B+��69�jS21��b[s��sk.Fh]g>:^�^�Ki[	��)P��Ԫ]����_P��A�u�Q��ab�Y[�բ�緶]^LBtt*0X2�H�H}dA6�<�o�	���g�gGn�5!��#���! ���=�T���8(��ۇ �/�U�/l��\�Fv�`��M_^%6#��X\�e��x��7�&#M|�ӻ�/�\\�o�.f��V��X4��k���������;lscz�06t���F�*Q (-�I]��qoAݖ&p�u�y�&_=�z��9E�������Is�!#QKX��T�0�b�/D!B����=���Hj��ݪLE�����UP��é��7�ty�D\�}�OYy��*��^.��$q�������q��f� �:����>5�=6�c��#0#�#UY�㬊���ɧw�W9��G�ka�!��&JbY�Kr���Ό��ch��w���ps=�!gY�6J�"$fn�3��5-�lQl�/5�9V�~)IJr����6� �E,���q�{���I��U������ۿTwMp�[`g�_x��E:ݒ%ӣ	 ��Q�3�B�'*�$�Q�T2��4ʶZ��6��B�>�r���̈����"�f�D��̖��,�(�D��'u�%�g�x�Bt*�*��SRԬ$9r:f��t5����L��3���Qs���--U2LԢ�RNV�#����"%����(�ҊLD�Ґ�5��@�(��J��H��*��t��U��Ԣ�\S⎪�@�A�U^a)�J�׆{"���Q�UuF�������L8TAFT��Ht9�R�#�$xM��Z©R9h��4��].D]��̔�!\*L���W5l��
�J&r��D���-K�Q�(�)0�E��µ�K/�QQ�ݛe��Ӣl��Q2*���:*�G.S�%�jQ$�,"���
e�B�:΂qB�(�ζPUh�d�1PV�W"�$�"�S�UT]�D�$��AeI��NE7\h-ݵ�z����ʼ����'�W8�s7d���ڱ;�.!���ݸ�e����n�x���j1g�g��<�/&Rs�惸���q�_�G��w�ˍE���}����~0W-��a)'y~���L�U`>DU�G��=��p~F|Ό�B�������G�{~�[��:���.�u�VN���/E+!L��l�o
�{��¦�؅��~t��xꌏvϲ�_>�����V���+�2]g�C��PO@n�B�K|KGّ�TC�H�+�WDҖ��'ݽ�s��O��N{4���/#}`h��[����5��spH	��)�_��9��ݔ#'ȉ!�FГ�}9�qR��>���&��g�vO�޶ w�[�H�����L��D\U�:�l�~��r�)��:��F� �;�	Xj#�5�y]����>���W�e�_[���9��CG����
q�eZ��t�X��q~k�������p�:��ǽ·����=Q��H�B�7Bv�k��R�I�>�]㶣�d��=*�~��,:�����mQ�Ǽ�N��h�s��X��f�4�TpEXt6��ܲ���J�G�|�dOT{�+t�͟i����m0����=��d�Q����f�����.�O���+괶b@���JE�����\�,�j�����WR�O��C�[<�h�6k��������k+�3�@�t�l�/�s5�9�9�<�
�Ъ��ֆp��H���Ҿm��V��<-ѣ�;�ޅ8���,�OgB3��jP��҉�D.�f��kG�'��z�����{��ٵZn4���33���82�FQ�Y�⧼;��Y@z#�wŜ�<j=��BߴV��=�ǲ'�i���3'jg0dc������Ժ�̴evJ\��j}�����}j;]�Ko�V��	�ˍo�A�,;O<%��|5�	OH��[��Y�'Ƿ���2=��}��_�iY�k��p���:z=�^�5�m賚f�y:Թ�N����.�	��|.#&u�ɟ"�9�G�����ב��W��«q�S�&�+©B��
�	X�qnM�SqT���D
�/ҙyU���c'��4VW��/�X��T���ؐ��B�c����wޑ�Jm�C�1�QjW���j9�@ُG��4�E^�A��o���F�'û}@`�z�~
r�/AʂPf⌏W�-�laɊq=�wuo:���Ruz#��3ڌ���ԑ�O�q�v=�:*�~�%��2d@l��m)[�"+m�Z��gc�� ��~����x�����K����%�.��e�ne� ?{�.�>�mS�4x�藒��8��ߛ�3�J*5n�i)�I�Τ׭�5<�����r���T��n���t�舝�S��B�N�:�afv]hʇ�'U%8n=d)�u��)�{��ru�;s���}܊��<�*�:�;��v7�LU�n�S�^V8�A��H{Q�D��mE�H�86�i܀^���cޙuS�W�\�p��m!�Ջ�b����/A�F�$
����\������n�b�*�X���_��R������w,���uW`�5ϣ���:�� �n�m�U�{"r���n�y��8S���G�+.�j� �w����{���s�{��u!��{E��ob}^��i�ݨy��>�Dzd�m���^�Wy�}�L��<��w^UO���0x����ǲ�8o�IG.'��q;,c��������٘���c�L��i��L����G�3� .�^���q>Rl��{���S"�}}�b�yJ8�^o+�p�D�ᗓZ}��p��F�o�j���}�����#yb���:��Ff���9}�j��W���/O��#���8X�s��=T=��u6H�x��=��Y0z�fg������3�lC}|�dn	lܕ���C��t��γy3��GS���� h����^`n5:��^�.�y߽����:�CG��P���9"�S�P������S&.�����m�#.�su����E���� ȝ�c�ǲ�\�KOp��� ����D�� j�;��(��O)��s���av��m0*�Bʵ�Ou����R6uv��+/.ޘZh7ہ.���bu�ܪ���ʹ�����TQ�x�#��g���gL�|���_�vG��<-իb�Uz�����l��Vg[��{�-��A,��Go�z-W2�f����~W�G��Ϸ��9�|o�~�nK-Di�;y���x�K�>7��'5����$_�v�&�'���}�¨x��[~��w�/q�5~�p�nĘ��+�w��${$�荘��  �b�ТW�Å��̍�mR\�<�*e��T w����_Y������=�``%�wz"�^7#�'�ق�ۊ�LM>�i�%���X�r��\����'��Q�{-I�gD��+!�g��J���(E�{��$������������ǯ�{�>s�5W�ev�Ggr�^�>=�~�=�M�C�X���&�j���p1��D5g��-�[כ�[�L�E�ˣ|V�J�G�!�\ٿ��@y�l{��$��9�]W��ǤZ�u] ��mN�Sε��)l�vq��l�&Mic��wa�2}0���7�Uh��l���>�yј�,�>�{��ㇼN��{'���ͭ��;������z��Z��@��3�3�ނ%�=�s���]�����i�]�j�W�L8\��-�;e̓_g,2��s���2��]G�guZla�ش\yY=��x�P5("t>Ә}Ru˕;:T�`�p�X�i��-r<��ug�� �gXoN��=�T�X"�E��V��h{�+�,���Ͳ�=w�����3�k��Ō�8q�3˩�+v�;,�ȶsh��yz����#����t¾t��v��y���ueT<5[P���u��\��w�xٖ���^/����В�q�����A_�yhpȏ-���,�L���QCՊ�ԍdtU׽/3����=�s��>>�����J�]���q��w�ȔyC���f���R���\Zڝ��T֕�|@���L��\d���s��8�����~)�O�۫W���+k\j��V(+�{�t�[�W��>��;n����DUϑl�Ա�^��N"Uy��R�߷������8��55^S�Y�G_{{�EWUW�G�]= %2G�e���+��m0�z�P^�.����I��ɹ�yJ���3�'~���S�7#L����T�R��z��Z>̏����zbeA�W��L<Q��_��}=�3��H�z�bi�=�1�5�2<� ɔd��9�N�:%�o���޳7�g���	��?%q7/��9�\
���@�=�EE��$y��|T��ܥؔ�[�%��p�	�<�2*�����ܮd5j�,[3L��x7�x��ov6�_=/��u!�1�a������{�j�>�q^w��>[�B�2��έ�wa���dit(�S����鹈�vЖ���voLf=E;to��".��Uշº����Y́�d[�7�7|G����3�p�a��x�z���߈�N��.'�@?)b�칒�y�Vȩ�u��w@������{�t¿�Q
��#b7Ӿ=��J�C�N�71G��yIf�{r����n7G�߻��+�G*D�Q���/��~ekc�~��?c��Y��1
h�+���O�V����^>J�%O��X���J�O���DOT{o+tøͯq������ 
����Vbw̘�5j:iK΁��]U>#\�w��/�Eh���QGo�ڇ��=��6�NEN�	Z��u���y�Θ�_�^��G<�>�ꡱ�h���(��њN�.4^�L��*�������
�l�7���o�,��@ڈ�vB�[�վ��F��\W�(�o$����3Ӣv�>�_��7g��^-�?��M���ó�S���Br�ώ���~Ϩ����k�������:F���.�{�g��Ӥ����ze�G�XQ�:���>E����}ヾ~u�{��dR��VQ�ϻ�ֱ�)�%#�gʭ�nB��fG�*�"�S�T��ȁ��M�F�����ł��ι�W�ʷ"�,I6k�8q���o����.
<ۻ�]����j]�΋)U���oc|���Zz�]Y.�yK�hy	.�v!��Ʀ;p���n���wm;��v#]�*u�
:���T�t�R,�ʴ�7��+���k8�d;W��;��0�.)�)�=$ǰV߬zD�<��S�A��Oq��\��[q5�StDZ����Z��W���-�튿W8�B㽽P�ґ�q>������)L�Z�L�����ё�X�e��n�f[>�Yץ^>Ck���)���F��Wn�i�zB)��~�r=�Ij4���P;.xZ���X��=mj��#����s��D��l���o"s�J�F��q(��aw�����M��Ы������ g�H�q/�g�10��YN{�FJӹ�,er���U+��A���ϩ�O����g�R�s���@/ofA��M9 _ШKG�麇���bb���q�}ǲ 2���,M���G �����eF���<T�����=w Tyߍ�rj��dNT=���L<�����~}��]C;�ҏHC���1o�R�Ǽ�,����!ؒ7�IG��o��9�0�)�J{ڲ�z�q���^�}S&kj�Cy��	����*a#�{�wmQ�^BJ9s�i�U�ՠ�?\vx�u��إ�ϬW�*Я'kf�4�zM������Nk�@��>��̨��{l�Q�w{��I������t���t�gF�lQq��d�_<�<���ش������3G*.幌嘞�J�Μ��2�5��[	���m�s��+���dN�q��GYr�fN�h�Go���	t&�g�*s����L��3�\��&�@�M0�;E��3)�og�NY����J���ϭ<*�%�Ӭ�����6�s�}~�B����4��^�*�5{⡥"��~�-�F2	�'�YK��ʌ����3�:��H�(��n9ѧ^���2՜�m ��}s�}�hvym�a�	l�`jڇ�Q��'Y�ɟ��P~qE��3���~JU����u�z������!���=�*zM���j޸s�Rv��K��Yݶ�n�u�}2��Ȟ�\<����r7ҙK�^έ[
r�=��N��;������<����g���Qԥᐸ�9�\{>^�����Q�h�z}įO���,�{�_�������tw���x���_�R:���N<�-�D<W­�[f3�
�9��6"33�R��k9�=�΍�:�O�d�lĠ hW���N��><��V���Z�c��<t[�0��2~�9?����� q�e��{�o���B� ��0X{qH�����9�wr���ʺ̪b�{z���R��⇧���>�@��z�q�̂*�x��T�$�b�&&�V�j���73q�Q��\D���� �&
<.��ۂ��������O�4�M�sw5�0wG���A
W���kK�n �m��A�Yvgz�ڻy�Yg\����o�a�)<4��XTQ�eo,;�v����u���U��-�ts}cpx{�����au�~�X~��NDς�6��X��g�?��J8W�P,�\��^|Ǩ�qzk��;k�6n=�@y�]Vg��k�|Kۍ��ֻ�3�R�X���0��"nP�ͭ�w�k�4���_�G,ˇ����c<�N�ze�_-.9��=Ge�x����O����x�OW�;��:+M��;,���#���@��}?�R6?��Y�����v4�o_��+�=��'�ۉڇ���,\f�i�r���`UT{��R�|*�c���B.��n�>'�堽r����z+���FS0��V�<��Q�U�!���Qwי���|�Bk]��{;�ݰ�h+��C�G��B���g��g�b����X��zCw�
�w��3aP��ls��O���ˎ���GG�u����;W@��g�̞IyV��W��c����~�q�+��>^��Х���s���9���Z��m>��^�U����:�7�J�w�
F�T��e��<���|�g#jX�{ԇ�#�t�up�5����y�oM]���:�[�S?,��U�R�|a]6��4l�WpkNjR�V�W]�F�D����|Sv��Hn�⬼'�����gk�Fˊ��n�Xں�;��^���R�p[��݈��}��UV�˹"<��eh�:R���+C:�q)�>���ǲ�,�dF��f�l�șl�n0�9�,%�؅0�+��^��_�*[΍��n���G��>=��'޿dxdt�7��!��T�U!�*����g�e���}y�ޮ�'9b�Fw�v!B�_�#��m ^o��w _���ý2<� 9��2%4VJugՆ�ԻۙO��7~�>��Gv&y4�&�SY�9���ǧ �$(�uNH�*>FȚ�ǧGT�߭�fy��]9�c�'�-�&+�����8K�_r����+�>�g�s�y@+���ǽ"F�z���T�tu���AN��Uǲ')��I���Z�|{4�q���g�S��Ӌ,z+S��̾���.����W@T{g�]��"�麇��V�x|:N3���c��*�X�!8�<}��Wڪ;ͣ��z;]	�顾�,�+�	Xo���Ϧm~f��+�=���%��­����鵝x}\�� �����~�>!�+��v,s�8+��h�ܙ�v�j�=�9a���������O�{��������^ LB���q���(��+ݝt=���$��>�3L��u�DɅ7ۻ�w��h�\��x�tc��1]�e �Du�;�A�����gֺ*e<��sڌ_ ���U0��E��e��!���#/rb����ܭ27c�;W-�W�X*�Y�P�}.�:Wz�u���Sj�`�*�K�������;��dZ�\��Xe�����گkN���lp�(SE7]���/�C�:c.h�vO��Ԯ�L��6�O����hs����F�5�l�B�t��t�`��G�ꇌ����~b�_dg]iά%�͈�¦���!�����7B�A���Y�F`�0)���*|�A��~i���ɪ��Bv��ʹи��8,���3�OC����"kC�>S�vv��+���ص�^���ts|a7�N�C��l(�*3���U�A:]u��8噖����h���WA(qjXSF����|�u�
�'m�KtX�j��:
��/*���:�Z�(}�jZ`=�{�8W:�^�7Ȋ��U�݊���om����We/G������T[�MXW���^����6���Yyٴ�pl��޵@1o ������u��8�W���w� �o}�eJ�q�V� ~:�95���x�*�������gt2�r�E�Y�*�eV�#�}əPi�
75�Z��"�:5�Y}�w{�2�ya��acP�u�B�����D,�k�Ts-ת�K�):w�#l���R���P�xt`�X�cж�u�jN��lp̼��r�s&��ɏO�+FR\��*��6�J��s#r]���ٍ
r�L�*���֔�2���\X�)YDmSPzPw6��r�b��7o)um�e���n5�f×s.�ޔ��;:���F�(���fcF�J�}܁���BŸ�!׮n%�4�@3��J�=î�V���I���^��1t���=apu5�T9Z�$1��'r��5&J��٩��>VP���ϻ���q\��&*�͠�����D�*�n��4E�z�-�+�kJ�uǀ�X�Hj��3Wq�V)5�����nɜ�&(3�1w��߶	�q�p�$�s�H��WX|�(�Un���ȣ:b�Y�Ժ��ۄ����ףxsUn���N�%=��H�y%��ݢ������m-إogU�#����'m6y �o�g`{�RƑ�ofۗ®��f�nt	.�r��A��"�]�,�kEgc�xLN,�|wsV�K�6��$y(�ֻٙ	��V`���0��и� ι��(��@{6L�,��_Ȼo	j�v�v���y�5��w��.g��9=�Vh3�*h��>5��f�(����;��ufvī���(sݏ�.f��Y�9��ؚ�cR1�n�ڰ�s�����E�NDDUxI\�(�D��rdr+���� �S����J��L�f�G�I�Ld�&���r"�\/"�V���^IW��*�DQ�r������f��#��9(��[���;���Qs���(/R��l��"��
�+��"���.�"���2��si�N�V"$����.d*��QG"�#�����<��]u$�%�\�y7���=��䎷<�T����*H�K"���y8���*�J��W!D��p��ՑNĴ1s�(�D	�u4�g��)YrP��n�L��*�$�fE�:9�p�D�'�8H�4J�����T�Ȼ�ʂ�܄��]�#�"+���&kwhr*��*u<��.�j�Q��a,�X��K�N���qnjQ�m̭Kʣ�"+����rUCM��H��e�k9!B��faTMR���^��\�z!DX�t�=Jq�5*���q�$�ܥF��r��-��@j���3r�K۸��Ǽ{{�34��!V�:Th���:'*�W�Y�f���q;���_���sX��t�9�ضh�ʽp�2Z������@��v.�}⫽농��5ym�W���ȟt{��}]�|��"�Fi8l�C����L^�	���~����{�ǲ{���Th�wS>>��������� %�~�=����%��98\U0,���:��L��d5�}㠼W�WU��E������n�>���vyQ�lU"E2�~�`LT� U�S/#j�z�玜�����XBQ~��GO;џo�W����\Ԡ�6F��z��n �ۉ�p&��;;��v^ym����_a��ʣ��=�Ȭ~���|do����2%VYe��'�n_Hc�Q�7oo7�uvMV�8���'�{��+��u�H��#������w#ޙ��-}*���u^��(6����Kc�i�A����dg�T�s>�XZs"6_�E��&���{�~'8�o�zC/X��#"����L��u�@��3�10���3N{�FDJӸ�ԇ����c1��u0g��;�d���l�=ʷ��ϧg V�d�5� )��un2�LM5[GY����91�N���^��\Z�+Vp�����R/&�%�]��f��wcŃ�t��@�3�Z6k<��6� �}w�n�(B�gT��7N#b�+)Ik���J�[ڛ}gy���r�Z� bwBS�ﶳD٫
�>�]oy�h��[7�Z��\r����@�1�v�C�����h����yN��=�3�;�MW�순�{en�w���Gޝ�X^�c����:9�U�Duxh�^�^UO��΀��.�g�v$��1%>��g���b�3�f��z�{ez7T�>��&kj�Cy���T����0x߻ݙ�7g~�Q�ʿh��\�zg:��7�W��%/ъ�z���ٽ,{�n"K�|�Q�fs��=ީ�q�ݸ��",�u�r�<^�j���rIzn%D����5�^O�i��#}7X_Bא+����'��������%k�#ɟ-θ���g�[z+����ueSY5��ɝ�r����>K.3*{=Y��3�� ��j]�#�wz��m΅Q�e�y[e{�[*$��0�v1]1y3��w� 4}��4��t֥��WyuЎ����������|5C��6�}�D��H�$P�+�`{��fb��u?���V��g�3��L��r'�\<�z]�ӱ�!��}��)O�|�(��ޠ)�o���5$��w���۫��l��8oT����٠���Q揩�����K��W��{wO�*����{ � j齥�ĥA��#ݸ(�U���G�l�er���fDP���n�!0��d��MEwVtg�vG�`�xp��6�rWy�����\�yw�ia��.��/;*o �ō�t-,ՈT��C��{n� w%ż����U�<_���ʐ��R=R�o%�3�����V�ϟ������k�g�w�R�R��ݹ��>�}q��t�O��ĶDL�<J�Xp�^9�l�*�jК��T���E��v���A���䶼\���]� �r�B���DR&&)�{H�2i[P�/+��t�����c�c�����R�W���@y����T�:Cs�����L/y-t�.��q��}ݫz�Q��v@�Xk�LW��*���������*-߮Q&g�l<S<��G�]ׅ_�ַ�p��C�[��Q��}F��/MD%f���/ea��P���X��=���.���%���Of��wW��~��C�s������猭�4��c��,̇�ꏦ.#�⧎m2���\�Z-j��(�4�g�e+�?�§���잯�p�vN��k���F�*�ǃ�n%��q����}��I.�F��ON?uX��Ѕo���X�?c��?-�������}{�$���%7�͇s�Q�ж�H�����:=�+G�	�=�ueT<9;0�ǣx� �.�H��֯b����K5�ėB��-,���~��Z|w��`SY����Wk�S����͖����~|k/��\�{�dv��M;����x��D�jX]��)˙iiZ秳&F�;i
G�x)a����G=4}�@޸=T<79������W�y�p؅��c>�Ɠ��L��Rh�ֳ/���?A���?ho��ij��.f�e�������t��ˎ�k�IG��dmcSZY���̀{�OyZ��O�l U�x	�w��Nc	���2����ǋ�\s�>�1�>[[)q��!�`%�u�x���@S7��e��<���|�g6��_�������n��Tz8�.8��W1����%/�ë�Ǳ��v��E -�#�-�*,��y���Վ3ɽ�
<��U�(yo;c;��\sG�~���9�p�#L������H@�J���;��)ݦsv�*��o%�d��G*�ZF���$}�q��4T_�܋�����i��6H	��}��Z����f�����y��Ҹ�����+�Y~� {jlm��$l[�e���:��+��%�q��cj/���)�i��x�闦�x�z��U�p\珤�rK�ތ�x��Ǵ-���x��H�_:�h�DNSq��=ei���wǰ2��pӟML'�k4����ٵ�b�*��9f��^�N{(p/�\�;b
f������^��S"U\���3�=ٻAS�(���źO�B]�)�9�V6f���/����bJ���{����R)qo2Ko��q� ��[�͡�V�fڹ���cKW���s�c�~ֆk�o���%�)�]I�X֍S�8��g�N������n��U��#�un2�K���Z�A��=��Z�1y��~�#i�}�l{U\_�r5���i�D�A��'���D�G����0�3k�n�z�f�\n���R�b���>�U�	����cUS�7���{*�z+E�~��?~��{^C�wF~ٝt���Ư|�v}�3�ѥ�����q�+��#!��i�s�~~�Z<�O�z�G�jc��o#���r�����\emǰ�T��|�n>����X�|z��z�#q��/*k#=�v����<� !�Oh�qȜ�����gK�ɝ��된�#����}]o�"��}�s�����Z��|������Q�Kdٰ{b��1s�,^L�8O�j#�Pin�X2c���5���9֠=�tyw����+�mի��{l���D�$W����@��:��ǽ0�OUR{Tz�=�D��K�bFO{ף�9��!�j��>^�\<�H�M|O ��MC�����ug�=7O2��Gg��<�W�����uǲ�6r#}�=��0t{���F�֙�)���o��(��J���G��_��gU��k<��xE	[K�Ü-��Q�U��u�D��%KF�%���$�[ *XV���u�'�͙�Xy��]���R5F
b�Y#�f.'���X���y�\�Du�t3fUŢ,X�����dmD�Z�|��6��O�����~��S;�8&���"c�R���~�΍>	��ϱF{$�}�@^6`�v�U
��#� �����W_W�TNq(�f�G�N��KVb[g�BydT}~�R@�8�3f<�t��s�:2�i܀Xʎ^�=����=�g�^wr��,ُA���L�ty\_��H������mg�wE�����銌�}\��,SD�����p���If��]�&��)f|�lNT=���0����F��vnVw{���2}e���:��j��P�T��y����-]�����"�ܔr�}^�{�*s�w�$O1�~#U����f�&�k�o��gf���~�US�.#}L7{�Q����x�+��>�G;�6YR�p�~�Z=q;[7��t͆���k3� _��R�t�^T{�;3[�;�z�e�g�~��=��Z���姇��
�z�o�����Z���{���;y�J�����y-��j�7b���v��z+��O�a�2�ٜ,vL��5�;Ҥ��/߷����`��K�tK6+�_[�ot�#�"v��c}�7]��O�a��5��͗S�M�G��2�nrNYt��Y�V�䗁��#{�u��u�Ef�����R�챙�BdY��U冸����gQ��m��S#��m���CZ�+Y�/7OK��vv��[�gjDz�?BV�H��>�=�����7�<��1otSg"Na=3�~�t��齎����*�ݯ.�M�F̠�}�"6�zߎG�ב�exu�����Ac�f��a)��c�;�
�o����W��z2g�x�O<�y�״��S)o���j��=E�7�U�����5���]��+�m��nO�(�M�
��r�M˥�q��H�����{mOh��L�>�Jp��y�ݯx��^ꠏ�4��= -����My,y�϶XOp��I��`��H7Z1���U�"���!t�5n�p��+�X�����R&	�g �^9�l�/r؞���s��x�;�]e��j�߸OL�({ޔ\�»\Q~�n�2�̢c)�{H��U���>�^J̼k<��z OOԑ�>S^*��+ެ��dn|j�J�h�L���δg�'��o����z-�u�Jg�z���y����z�T�
����w�L���o�ި��齴
��+�P[�3����#������>�q�餬�6�SG��t�ȗU�ܳ2J�4���֩Su�e�5����ݦ:�|����wu^�"�!����lV�d9�R����A]N8J1t�*×��R�9/k���zʹ���O^)��qU8Xji�t^փ��s�,j�N�Pq|3��^�LG�YFX�>���ی������cL�F�=Q�3!��;�釽ӕ�=�k���ޙj��W�Ｈ٧�K/N}?�����,�(��Zn5��f���,c(���/7�-��r��u���վ�Ι�vՊ�{l��<���q>����Cˌ�qb�3f��CKQ>����=��e�ל���x����J��߃ϥ]��>�����{D�F�a�.�����Y�����%�z�Y�� o��G��v��N{g��H+���C�Dyh��vsL���@D��{��,�~�Ƨ�GF�;�xN�z0�f�e���>�i߻��_TųП����w�zS��Hʋ�>Q���Y{��w�
W����}�y2���L�zy�qu�9����ԟ��pyT`�ُv]�exW.��=x|���r��+#�@S7��L
<�Ϯ|�gd��������5ʮ��vy:��f�k����}��z����,�p\�H�*�z�e�E��O��5�}U���8���z-m�q	���+N�����~��U�P�L���'�=��o�B�d�5Ee`56��/���[��iܸ���n�9'dZs�;�I[�SL"��OIIU���;�t!��k#qX�;{��j�����A+�n����{���kP*���j�_�]w�oċ-;�g}���ޡ$�������M5�eA���r��P30������z�n�+Ty����~��{�H��a/=~���wdy͛\}c�s�f<��I77�k��V�
���<.����޸��__�G�x�޽ ;�=�@���*-�;��{��ԧg�0��${�}A�����"b�����%ᯣyx�{#ʫ����;�zｬ����k0�7���멒5L4z�n������i�Z�|{c�P߳�"6�{2'M�P1��=��w*S�>����;�+���U���<ja��n�d�t��:��s�O��݄�����VK��^Fy�;5�4�<�� �;>��]Q���0�"M�;F�]������(��}�����3�j�|E���O_��b�Ǟ��~BO�Uu�B�-�c")U�\�\]%�q�U������ YN������+��>�L����_2IvI�fC���@�8�b�ם<0%�=��-'�z�W���N�ry�w�j�/O�>��ݕ	 18�ܣ�О��''�C�gK�s��Bs��g?_�Y��v��j��C�QV*{c�wr����znb$���^L<��V�iR�~������)�ʞO3E��Q�.��x�ܷ�Z*b�mP�|j��\�{%[�������x^�sN��!+��c>n�Ïw�GW�n�q2�4��{��B��U�qdjH���g�j�G��{:Kg>�����1s�,\dγ���lz}�(u�}���JE{wO#��s�w=��ګW��|c��2��6���T� k�l&��[���w݇�3W�^�c>�~���\{ޟsU�
p;�����f�% ��]s�Nǽ}��]��L^uW��}YPѭ{��}^�͝�;����^�NQG��O�*6�؏wL�s�y��B�9O��l�Q���Z�2Z>�چ�CĮ*�׭#��2�7�:=j�z����?۳W�����H��x�\i�"3�J�W�ϑ���4�m+��Mg�篁�*�Lm����*�XN���]4꜐?(>�P`��t���=�x�9���}��%Te��>��龔�[��]jc �izg"}9\{�pj-�zH�-ț�{q��b~��h�zc�T6�]��}�ݧc7�5��|9�k����s�z���*���j���ʇ�B�"bO��+���UR宙��t��iz}W�ᢾJ�1qUO��΀���x����1%��+��P�L%U�9�Gz��)���݇��<�3��I���ye���kAͳH�Y���{~b�"݋��^wBP.�sw`��b�!}ß�9-h����X'�F�Q씎Q����wgf˺�ؙA
�|6)2cle��U7�K�Q��V�q�G(:
A��:o��T�0�q��:��d�5���w��1����l!8�Ϊ���]r�,(�tys�W���Q��i��Rf�|p+$SH����9rfp��������x6р�v���<Ԯʽxɠc2����5:-&gm#��|���N7���Sk73:r�C'kx����0е���Ň�)Mg�!Nf\9f�f����1՝����V��,;)��t�s�*��l�YGL|��0GY��X����� �6�����ۡ���$�>j+���{���#�r�ƙ�ȗ:R��c������H��RY[���m:��%�l:�i| 2m��@u�w��`��am�(3Aٍ� ������[	�˗M
��Џ�t��Z2r�+�L�@�b���I�$�*���;]�kރ��1FgxD���zWg�i�(ݡV�|5���5���Mbievo"l�3-dl@޽�����2� �8�#��Ln���`�|�Dl�;�݂�h��֧�����^`�E�1�1��4�;�+����2�T���y��o���X�{x9���=�����ns���r�u�/Q�Y�WjAb�n��[�n�P����\�uۈ���"\���*���q��sQ��Sܽ�7gEW0��L�f������w(�����r�r�6"�6��rP�>@V�ܻ�6��4�z��`J=�EZ�i��3;;{�������L ����
�I�zǠwUaav(��K(2n�429�/s���� �k{���Aڀx,�-���;Ol;lc��F���.��n���U1|�|3�=L5�*��kW`��gV���Ot���z���_�QoW��KjۦYK~L�8ڤB��HZh�V�-(E�Ǹ�S�-�O0�Sz�^�X���F�n���;R����<XVb��`���V�w�_Y�nT+9J5�g����Rܓ3�a�uB�s�!��D!�3��q�>}�Mu�-(h�ٷI1��^~��.vW&#��m9�^<�T���o�d}�ξU�n=Hn�]�S	/�S�;�[��;Dl+h,}-�m��ȸ�&B"j�Jn��Y�S�X����y!����#r��Ȱ�X�\��L#���M��B�D+O�,Yn�,�6X=&�Z�NH��%�k5[+���q�&m��о���r��$TK�o:i�'���v��&#�r�����ҥ�H���JHb���[�oּ)՜30e)W�uo
Y|*ɱ�0��'���!�̖:gT�����NJ��nd3m>�5Y�΀m��%p7���hQ��������I�0Z�Hi�|RmC>@�"�J-iwWP�*;����3��櫢�js�Qr�RU�䜐�7$��3�S��GR�CE��(�A����^V�Ց��C�����wJ��q��w�s�	�J#���UjAz�H8�I�ts����L�:a�J��t,�,����Ԝ73���^�;��^�Ne�^b@���*���e�U[�wtL*/s֢/=�wp�H�S��!;/-9;�(�!h��M]wR�N�I�9⇝2"rs��	�Q�:�*k���wk�;��DE�r���B�tT\���G���(��*���'Y�r�\�"]3"swqVbS���S����!�i��ܜ�{WQLBr,u:Rh�s�s��wӪp�(�wQ/;���nC��[��Q��E%Tz����wK�����p��T�i���⅝"���)x��u9zܽeN�r/#Z�����u��ɥIUS�o�W�=ן\f�VM�Ѯ�<l��֥��k���ʗ̥���F������ibn`ՎV̬�gd�f�T�"��/2��˻���o�������5T�������?�2��>#
����q=��Y��+,�ꇃ{}��!����,�L�ZnvX�b�+���,	Y~��Bs]��Y�J�v�w�k,��SD��+ҏ��n){(��9'�E�O�Pۉ�c0Εѓ�Zu������g$uo#{֓������SF����~]�va��)eSY5���&wǶ��y�{}����|�|^u!�����\�N���ý�7ݔx���rs	�~;�������ݼ'5Z�5��3�o&P^Ϻ�F֯[�ȏs�#��Xq�e��#�JohR�P=�Z���m��w�^�7�{�Rf0Ey\;�+��2e���.qu�9���^��Сիbg��k�f���=�Y��2ǰo���
@�N��M�
��'/#f�F�?<�ϗ���!��[�~��T����#Շ��x��C��e� 6B rت��t�7�Kgr6XU�_
=x�y�2���lw��6N{4ǡ(�&s}#M_��<����3혖����ۈ��x�;�r�s��h���j���ak"o�ˎ]� s��T_Y�Ɔ^��(�w8PF:�)��ltu�v3�{��|��2o�_�2��S�zSD��=tBT-�Q�GrdGj7֕wqJ����Yx[�u���xBB'iB���^	*�
�Ԝ3��@��!
=���c�w���<�bn|�x���E������m��x�����o�D�~Bo�˚3�KZ�J=���W���d�Bt��ȟ*��
�� ^��dV���\�Of��>kLW������h����;���v@�xk��x[��þv��f��T �4r����½�ƽݫbU9D�"j��a���!����:�Q�/M%f��5�7���"(!�]m1�=�����f�C��_��Qޟ�>�����͈ͭ�k�j6X�3ZX�r��pg�*�o��-�#���zc�v���o�w��.rϿ�¾���ǳ���6���>��tV��s���J��*/&�/!Wy)��ܯ��P;}^=7�ڱW���������t�û�ib�bN��q�:��R>�r���*�@�^��'�xr���B���V���]���8�<��uP3���x.v��g���}
�P�1�Y��������G<wޜ	�ye�c<�R��j,�*P���^]��+���g7E�Q���N�{�&x�3y���>�K�]�G�V�o�u�>м3pf?��h�u�����wnr8C�l)�ؕ�v���kB��#-�K��Vof�P��iȊͰ�y��|7A$%ɵ�3�r}Q��*�֊�a��L�32���Ɲ邴ZZŪ�:_7���U#�cHX��=O.����-T�brsC�%�QO�	j�@��T���\;ɔ�.#&|�9�9��z]��Ҽ���ޑ��r�z3�x�z|�Z7��Q���/=�3r��T��Ȍ��-��jX����<�l�i0���v�K�\��h�Q���*�>�����q�r�1ٮ)���d�t�d{��a���ʸݸ��Z��֧~�;ޏ;A�o�2=�Lo�Oi����e�#�>���z�Ķn	p��w�/B��?���؂�'%���o��h\�RG>�{i�7���[��W��>�7��Ӵ+�kos]�+_=�+��nL���xr ���	��n�S�~��x�`vG�����Q.�{��s���y߉����LV��g�����8K���c��+��^r�3���7:.�6.����I��P߲���u�"��U7,f稏U��"�5�xt.}z��\�T���W[Q�b����~v�&3��	�e��|=�-��K�qu>Ed�Cی���'ä�[lU��V�3~�[~�g�ux*�z��j��/�t'���� <�� %a>>Gzz�����s�3"�b�'�s�SH���@	d껙��V�����;�Wڅ�V)p�n�,w�𳹁[���<3ɶ�g^v���@&;�����64�:g/����pкp{ˆ臖��{�6�:S�t9+1qv��Z<�v[e[�r�=�گ�UP�Q}R��f\�%��f7�Ο���3[L1	_��!����nJ���P�hN
��f�����".m���w�ˇ��	r�5�Ӿ�P��F>��l���Q��-��]�3ʠ��箆w��<)�99��F�z�q(z����=�*��7;,fN�.�����OOO�m�s�&��]~UP<X>=�||�s�r=	�*�삾���y`�٬��C[���<�f?��Bsq�G����0��^���3�}�
t�;k�=�a�����vG��F���/�իe7�[��O�����;+�I�W��ԘͿe�UA�S��|����*!ի����x��D�=&����`O�=ʲ(�sJѣ��߲��x�2f9�����do�W���î!��d)��;#ޡ딹��L�ޯ]�4��o��`LEwPjW���h���?C>��o���:�h�����>�^&��Ӡs۞���^�@o��2���ٸ�#�ݠn2Z>܍�h�J�������"�����&��|'7ݞ]�y�b<��v��\?UzK�2f��L�Ҫϑ���26_��{�R�����}FGf����+�b�P�⦩�'�,��b����K�R�Ѿ!�Uٝ�E�y�-!��b�M|*R���t�0{te2�m�6�R2�����e��ls��,sS��i]EY���Jg&#�h-�ʽ3j[�ֆ�`�ڳPM�+����:gl{Vx٥iJ���q�ǧ<J8ߨq�m�s.Hq>f�yP�L��>��m��+�m�Ygjrzx��3�H����z�0Ͻ3�>�_��*-׉�P���a��+@lY�Ƹ!��)����ҽ�}�X��,g)�|5?U���|�{��`z=U (�@��U�y��S�U[����n����u)�0���Mi��U�xh��&�Nd����zມ�9�X(���d]킟/��Y8�{��E/Ӕ������ڇf׸�q|L�mC�n�������^߻f&֊}����>���8}�Q��a��vX���u�\n4���&1n{c�(��Xkx�+±�a"� {���YQ��m�>d��z}�^>�����<3���M���;R.�+}
�ܣ��>�Q+�����#yb����m�1~z+��gESQ�ZX>Z<Y�1q/p�&���Y+����j�7��G���$&�ߑ]n������)(�z�?x��ݓ�����U��JS�(�׵g���}n�^L�72�yR#kW�����^G�=�����ў��Aw�>����TXO&�)R:�oY���G�;V��[�����s'Gc�(*��t�G�j�q ɢ�{2]]��qhb�G9;���S��8-[w8a�1�#ڽkȺ�+/��Ȝ�|)�S��5y�RGFl�>��cY�,nl���-�͹2�ѐg��]Z� X̟D���pʣ�0�f�e�㒓܊��~ӟG�e�o�C3ޑ	��"U���[���n��R��oM#��.�� ���w�ԙzd4Ts��B>����b7N+Ƕ�c���3�R��Ɨ��ϸ�z�����e�2fʐ�UH�K����c��F���3^��{<�%��^�yg�cT��ǈ�4������r|/&%�fo誐x�>�ve�f̡�S�����gzt�(/}~V�ܺ�3�{i;�5�{2��L�/>d@������U�ݻ{۞�q1K'���[;��z�:H�d�U��=�����\��I���z�=��$ܺyOsV�E�oO��&&)�m����r�~U~9��=�̀�F������Q���K�� ��(����a�߳h�Q~��Z^�Q����	�Mz�̕���]�Y�~�JԌ`k>�wz��C>.]�W�D���ͭ�w�j6^�&����y�pw�}ѭ
�(�L�����ڪ��.!�7�Uh�@yF���%��>���ǲz�͜�tV�c��z3bb�+j3�ՙкWm�z�n>n%��Ԫl.��rn'
]5nw�c���5����<���a��~�^�Nxk^ �׶�c�vj����*�%9GF^��O6��YN}�(�g���y�� ��+�PW҆��E��o"��z��B�a��lxk�����S.oݵb���:b�=�E.9'ӳ�i�M�S\s�w6y�(zMi��]�0'�l�q��~D� �<�Сq��Eh��=���TĞ��n��_��ETn����㮳�����xm���
Kk|{��;��5�Mo�>Ÿ6��ʲ��Oh��}3�M���b��d��o���	��6����>�K�]P������������ؔ�C��vz�5�Q��]�̈́]So�p�2e9���R��sA�4w*r��y�7'α��>]>�H��8�SϨ��=�2Qf�T����DW�>E�5ddq����9���&^�F׬w��փ��lv8�w�q�W�V)��uƸ�f��d�HQ�9:�]�s�W����ȦR���U=|(/y�;�+�f�������<ni�ܾ�~�3�0u�M�=|�o�ْ0z{�aȂ|��fI�6hd:�6sޔ��X*ݫ��<�A�eR�����g�����ٔdg��{A-܁0�jJ�n%�����u��𑞧1銂�"�������1qպ{&�D9gt0b�ȳ:��
���f�.��꫔T�ڠ<��Xzk<,�}Y���Q���KÊ3��W+V=ZE��]9Ȼ7fVx3�Qn��aF��/�5X�1��Y�*�R��ewn�m���� ��,���W�����Ș>_Z�)�Ӑ�aD�5˽7�{��<5>�����{�����T�ɿ��O�`W��$[���gӔ��z����F��wǠ�^:�o�6{%�Z|�����j6�z�71q�:S�.r�;�y׉XjO���&��V�}��+S����+�z�R���	���@�F�Qʬ�-7g��t����M�d>@J�O���zۣ��#�2d��>��[N.�
�L<�z{��3_m0�W��ƪ��^��=�eP��碴Цo���G<�`m;݉|����2�����G��{��mV��/Ǧ��0-�`\/N���^W��������&{�O��}��[��>��x��h�D챗��
�Ԭޖ�n8��ݮ��Y��&c�����������?�K�;��o�\G�l�o$���98L��ɭ/	�Ltk���4}�e��宑^���`�/Ǵ�:����y,��C�D�rrp���s�,(10�V�;�oVz��ocW1��>ٕ�#�T������{+�nZ�܏���#�L��m�	���������7sc��J�Bj�nރE�4Gh�&��乹A�[��ԎZ��pb���{K�A:�P�Ý�vZ��Kf�Wp�5�{NA��c1d���a�\���m�r��v��U�=�F)�k\*�E�ҷ�������� ~�S���2ҭ�8׋_��!M��^T�������ɇ��=ޞ�Kס�冼Hw�j	���
��+��mCF����z[/}�ݾ�0tO�o�ك~7�0���F*�
�.�L�������n�7������%1��i���Q�=�=\�t�xaZ{P���~�'�Z� 6l�l�Ҫ\����4�����W�~��2�o�p�FbZ+\Iܤ��>��Q�zF�y�-̹ /�_�<����=��-/O����A�>̯V�@:1w�ly�2��|�zg'Ӏ+��̃���I@|uM�8��ِ�Շ�({�N���Z���j�Tu��`1k�Y,'����8���
�;�a��q�ﶥ N�'㟷��X���-lT5K�0;��풼4T%f�����x��=���?ݩ�dNLy��w�dz9�,��K��p{NnL>ͯq���&kj�|�e�d5U>#a�MT��x���1?j�h<}�Q�=tQ�hIG.}@-7;,g���\�t�i~=&���ﾏ�<1eߢ�U�ȤHA���3��M=���F�
��Ҝ��u1�Kc����2���M��U�#%�X�-7֛#>���9�l��!݋7��f���ݼ5H��Rq��1�*hb&a뢂�W�9�Z�=gBh�R�w;��ZG�d�����Ђ��+������u��.���ջ�>˘���Vtߜ�{I�0�w3�Y�6�Z}�(��gofu��|�D2��{쀲}���=�H�Z����m�1~z+��O�a�2ŵ�V�O2*_q��º�gG���)�3k�7��T�m�m�H���ǽs�{�W���V�pKf��c]ϳw���,�x�?�n�a{s�����i+���~.5O�w#�Lu«�4/N��=����� �V ��/w�R�(%&a��]뇀��[���uC�a���L���3^��<�ڳ��{�H��U��Ϝ�{ސ%�(�tXM�
���r��hοu��@�Vw�.�պ셈����f�A8�����:�ޜ���L�ٸ*@[uR=R�o�<κo�$ȿz]�'ůz�_
�o�َ�)�^�F���[�u���,i��4<�#�ԧ2ۼ�kW�j�⑿Dl��ڴ%K����J.}���Ր�����P� �z>��t��y ��fO;��uY��0�r���1����9H]1�gtQ9�鐟����c1���1���l�����m��l����`�6�����m���cm���1���͌����co���}���m�����1��P�1������l����`�6��6cm�a�coa�co�����)�̵�� ��o�),����������1��}�*��$�H�
UEPP�DT��P
H��RQ
�AB$D*D@�R��T��U*BUED�"%owJ�	BR�P%"��� �RQPT!%T�I!U*Sl*��U@T�*J�*�B["��ADEi����:Ĩ�����%*�	UF�QJ�)%QU(��)E$�P�IITIEQ�R
���AUA"��R�;�9�(P�  �U���X�5�@��5ZiZ��(�c(�E�4K���$���T���HR�H��P�PJ�  ��
������akQ�m@�(��(wB�E��)%:�Q@R�(���t�@����)EQGp1�E�J�㛊(���k��R*����"ARG   ꪥ�Y@��#f�`4Y&PFb�j���`����P
њjZ��@)Y��TUĕ"D�b���  0
P�Ҍ ��* �L�V��M�X*�-��֡��٩i�jb�CR+j1X��Mkْ��Mf�*)����"� ��  ;�jUYkX@Z��jU��	���4+kj��&UB��e��j�4MD�Tĭ4eRj�X�
`�4+m���h*���*R��T�   �D��D� �Ra-�5mJ��b�m�i�-���jZYViAfj���*��5���E[V�6ښ[V�m*i���XФ�*I)@E"�  fu*�j$,j�
��Ͱam�UM5��e�-��ֶ��ҩ�i���d��Zl���d�)����kTf�(b��)D�Q-��  3���V6P�I�ʚ��j�ak
F�h�6j��mT� ��d��M��ڀ��*��Z[V��� �T$ �%AI���p  r�Z���a�ڴ$�Z��Zl�ҭ64�T��mT�بhVV��5�UPj�ҍ �&1Щak,�QaUU$J��*�   ��*R��R�֩-FE��V��m[L�UMR����@ғ-�m���TԴ����2�[d� ��   � O@2�$�@ a h�S�0��%1�4L�40�� "�2)�OQ�MI�MG����5<ԄS�A*T��ڄ�4 d i��1�`&F F&&	�bi��I eR��1��S5��`#	��������+�_�9����;��e5wOV����p�
�"pƷ���DD_�%j".����� ު�"�O�"-������d�n��A����`�QDD\�$rB1]
""-�;z[t�Z�1�p��헨����ӕ	�i4p���zc��̖R������q���y�z�/�=��f���ލ���Zvc� ����󒖍e��� ���-��z���֊X���s�Y�)�Ђ�I�j�l��r���w^���� ;�([��9�ƬԚ�����[dn`�d�2�0��e0�b�4Z��h���������tq#X���a�q]�Sv[N��(�PX�è�)�KcyVj�兒�q�;g��e�K�֚
�^�`Yǳ]3�T���uV���/v!y���B��Ib�a*A�p�%i�n�W���u`e+F�L����, ��*��#G3t���p�	6��(�����I�ߎK�JJ�=�n	D�;����	u�l��i�ط�șۨ��y���Q��6�'r��fK�j1��^�y[5 j�<��wL�=ғ-�7b3�~���R���L
��f�^9%k[p�*���b��Ln͑ʳ�%uD=�ׂLyVMx 
 ��P/����Pd�/1bɱlR��,���i��hc*iGnn�1VX�r�-�z��x��`�6�[KfN��b�śs�hQ��Xz�p�Q:]$%���ʖ�u��������LR�*�:M�F���z�k^�4��-Lω��D2�Ҳ%MȉR�B4��X �ӛ�M��M���3iȅ r�B�݄.�=��:�t��nZش�|���4���E�u�`��+L����Z���n���)�X&2����2[��������Iؠr��JU6���4N���$Z�
	{�:�����1���"�K`sj:QG���d���f-�(�U�m�iՒ���c�ͱ��Wt��+V�P��re��n���|lf�E�-�Vn�(���)d��.��Y�h:meO�6���U(�9)�3k B���v�wf���a7�XEd�֘���Ȧ�E���A�͙����)����
�+�{���6<q�Kr��5P;��f�m��0�F% ��\0Tp�}3tn�YI�d؄n"�M|f(2έ���Som<`[�A��k�Yb4&��pR��f*�����R@&6���0 �A�����d�� �"��am�DYlg$�WwL+n����TU���Xي`Wr*Ӌ+c���E��2ݗR�U�/W�-9���KE��WtŊ�P뗄ee�����sӛi�F�n��*���H�)z��KSq3(��v���n�]-u�z+"9��r%O4niBY	��b�M\n2��6�8�[�ؚuS�H��:��2d����U����d­`��M#��r�ܷc;Z�"sa�wilp����+M,!�ӈ�3jݭ��0q�u�Oe�R�&�3h��JIZ�٪Z��L-��'.�Ȃ8�6��wz�E���6Ӈ]�,�խ���@70�Vȍ���A���B����1E��� bN�śf:{Q�:B�bw������4Ψ���4P*fjai��S`�b�n}�~E,Bن1��Pͩ�X�åi�0�����e��.��;��%`��N��h�!�Cbi|0��;2�ĳ���fȭ�/&&��-y6Z*h5��ca�ܼ
�^Q©G�PY��eN��#Ř�R^�u����WRN��Y�S%U���������B\E�����xؕiR����$c֘	��K� �h�x���Q�kq���8i���{E�:��4U�N�5xB���Y0����	UR�T��u�J��
�]�E��tĵ%զ�٬�	cź��Ȉ���֦�]�$�'p�#����pJ�F�wZ�k������+32�]j��yYD&0B��ǰ�tfV��	���R[���Y�[9��ں�^<���Yj|0
Ec
��iܻ^%444�uz�c�����R�5 \�Qp`U{��*�F�J�'h-�9�e�{�#�t� pI+�[˭	$����R�c#4^!i:J�&�B7zDkJ�X���$co5`UJ82"��B�n���݂RS�;���7*�J�m��U&������������Re����^) z0a5��
�����g����#fa�ܗ%����T,�e���u�3 ;Xp�8����SU�V"�փ�^��5�wtZ*f�Nn�J�u�`���J^,�t�qbŢ���@�j�#B����4�ו��6):a�ND� �qbhiA�9t����A
��r��7Pc8�Q��[��;C0��h�:fҺ{�W�RRV���Oc��Ш	��F	����u�M�*M�3�n��u�%�m�[tKH d�T"�5�T�db�����z��wr��kH�D�4�ڻ��ԛrAtov�ۅ�F@T"�ځ����I\��S��/��%:�[w���f�%2��9p)"{wqAx�X���n��p�ӶoP�����a�y�S&�i9���tS[m:	,�iV�.�h�&��`T5��sj�hR[/MK�&̣-�7#nՍ;�w2VGV�d�m�q��Y�,8ۄZV&���ɛ��1�P��̘�4��5��ڈt�1Pc7h]�N·LZ#��qM�#�i�wb�¬V;����ɣ6be��0�Sn�;N���+h����Rl�wwCe�3��N�r�5�[*BRK��u5�����V�F(q�W���f\Ѵ��/bw6�P5(�q����iպ����\k��Ex�m[`��3绕�H�U�tK�D���qTc�����Ą?�h�OC�4T�Ѽ5�5;��o%�Ҏԗ�kB��V�;���b�)+?Bt����)�;�j��G����K2�wU,��q�,�&��n&7u� ��͒���z�5hF�rꮯC�rXnX�aA��Ok���͡t�H��揕-Y��M�r�͵lG��Yc4�0%N*��Pb�n�(,�"c�4����1$�˼��husif�5��f���9yD�N2��Q�����j��Q�&=4.�>
���64�%�*vlӴ^n���1r�Xͧ�%��{�R土��k/^X����UM��[����A��D7/,(�=�H�L�sjKS��Qn�<;k*��)�����Z1 �OlBql��n�.Pk_�0o+Rbą sF��YYV�qaw�^*P]�6�4*2�IX1c!P��r�
��8��CX���aa.��V֛a��SHh��@4����`�*[�(:v�L�LI��lR�t^��j��5[F��J<̏B6�ǈ��-R=�m���8�O����[O��(����m�2��z�+�t��h%�X�IǦ�hM�Z�������*�;y`n������lcڱt�"�70�1�֖1�S�.�8	��Ko1j[�ťd����p#odV�L5*�v����7�c�Af���50��6u[(���YjR�Gp	�FNP��/S(D`�,�k�U�%��%��)ʱn?��e��1��<P0�m�@�
��j�[1JiX��3�^�{ǯVO�^ؗbچS���<`���u���˂�D�BX�g��+��&�j�3v:��S)ZN���m�e4V�eR��b��܍6*�Y�i�q�1���cD]�7^)ݬ{��3l�+SQl4�?w�,ܙ���W�2�� ����o��fR��J`Y��ϋ���=ώ�v�Ӓ��7X-�NS�����
W�#z,����P �8�"�F�бǛ��CIE�q��IQ{z"�P�*VU�˻b�O�u�I���]LR�
|*jx�X�Okf�f�,��Z�: -91,;�JZ��zA�%3W��%KKK�Y
<�	ǂd4��{1'x�+�!�˖蓮��!���+l� m��l
R��ve)�BNڬ�ҭ �n��(3��u�*�]Z.aUd�v�QFVP�%2����Z˥9e�����w���%�16��2�ɻ�,�B�U������F��;��)�hɽu�O�2A%�e������[��X��W����cI��P��F�a�Bm�q�i��T(�#7�͋�i9M֓�/wf5l�n�|��h]ݩV��U�j\�� .�^�$O�e�F7��)�WN�%��t��P��Xp`w{��7fjy�G�p��'�h����Rő�QeG.�٨\�T3C�	e���4���Ғ�Yod�3hLE�r٭�E�=�EX3v* J�m�(��S��j�+�x��r��S�6�p�+0B���Ϋ�F*�WTS�Ib݋�eA2�G-\��)���"���ɵ���{���(֔�nZy5Ҧ*-�Ki�V(�ܼ8c�s[���)�7%���k ���"L�+%��x!�N��toJ�$�w0�u�^�y)Q��&cȩ庑����+xj�\t�Z̵&�LT�H���	��n�Uo+X*�V��>x�htt[��(bT��T��s[�m*:����tr#�p����j��eӅ��eG.��Z ���;����dp�P^�-#R�`�ӻΩ�U��ȝ���4��	J͢]$�ԕn����*��Q�B&��c�f|��[��e��6�f^
Ɯz�:`�*J��݂��@1�7�m�l�3~���YN$x]z�ʉ�ܵ��P(�L�U�$�R�F�p;��>��"'-V�pJz��㺳�D.k9�[W��M���G��!��ӷR�+�R ?1��/T@��5��7{��%�8��Ҥ�W��a��;�X7NX���)*Љ8��jHۥ.���m��HS(���re��keց�:�͍f)�L�"�0^��
���Cr�xi���Y��>�,L֍�2�;��аM���:�q�􅕴��)붣���`����m&�T�2���,`7�i�n�X�s/�)@�B���A(E���	U�A8��E@��Y���/t,�-���Ab��,?��y�p��x����!`���Rġ��	`6�L�@T�1Q�z�4LJ�
���ONޜ�cCF �����ESv�@Y֨b��mް��X��(=F��E4n� ��ֶaҒ�e�v݇�K]�폜���j�d�#�M�V^3�L�F���Yز�XS�%����
�(�bR��5���hڦ�ŗ��v&��t�9vf/���(;�Ĥ6��������)�KY7.�qJ��]k-�r�1aT)XN=���x +x�a䎅fU��7X1:��5m�
0v�� t���)	�e襕���G�Q��k1�ԙX�]��С��/��2�C��Ú�l��h����4�z��.$a�b��li����¢.��m*e�x��e%�"R�l����y���,O�2�F��1K�	�LX)mU��SJ^F��f�e���X�^SX�j1���V�uVva:�-�b��j�Y2�ÖZ�r��L��,��T�G/JAz�hN^ʲV��P��`;j�Z��ͺ;�Nn�cYT6n�T�Ȭ�;>��g�4J2dO5�f�^0��B�x)��O\'B�5�&ۧw]���.���k�o^�p#���6�k�@.IVHt[�fc׳U[��SB���Iļ�]�wlQ"��	�tSυ�;
�sY�q�G{E��m��R]�r�TQ�J�
R��E�Hl;�R���z�l�m�ƾ�F�M�vpt�yBШ�\E�4|�FɆhԭSy)+E�(]0�P��p�NSY�Ai����R��m����X��#��n�Z��[j"�Km�o�)D���%)o�X�9X�Qµ4�ej9YqX˶�� �ƪbVŌ�-N����|��von�BZ�i���:;w��q�ƂI�߲�Ȝ�YE���i��-*�	��6�,�A���_Fu�ݗ���)_ۄV�"����J�N-Ԫd{)m<�ܕ�t�*�X�7u��2��ch莤�Tw���N�n�Y�+s�B����&q@J�ލEf�H@ +Q�j�<�r�J��zĹ{E�Fa%�Ʀ��2kɭ��Fc�M��L^����9$lb��e�����L'O")�;�.��Sek3F�fՖ�S��@���3%�E=��t������p���hn>�mʹ᫵�F)v�QkQA�m��N$����MT����!�[����cl�*Y� X��@N�]�u-�a���(�l��֌�y���ݗ��e��l�oh,ƱLWz��m�i��ٖ�㬷zr���8�,�i �mV�)�%ohd���p�����3"�5hґ���P��ʚ�k&hh)�\ݦHP&1�A}��i�����ff��J�����j�R�*Q�52n��t^�LĢۤ)h�vP��v�ދ�`e=T&���L6Pw�A	Z,B���q�\i�	v�Q�SD��(*KF\g0k�j�.���{iqm1m���g~���˵LX6�yY�Ymk�{0E�h(���ttbR��� ��y�K���fcX���{�`6���(^��b]�b�ZV�Ӄ �X��sK�[U�u���^.7�[ˆ
U5n�Y(,�X��'5�˧��aK
T�.!�b��峚���ߨ5����������_�T��7�Fa��?������$µ�%ګ5r��qh�*K�i����y�5��o��l��2oVM�<�5�Leʜ�;w�r�%�eIx'V]��+�5{�;H5XM��jʡ�F�d	v ���K���x��w�:�������� �;_D~�H�&��D���&�|/l�M9�㽑9J���r=�o_U�SN��(�� �]�:�k��h�Օ@%+���c���-
P��mJ9Om	�g����6j��l�Y�^Y����J)m��=�Yz��=`E�/`N_N������g��̊�\��&U�-a4��ꏺ��=9���w'6�T��fX�Պ����΂=��+�f��De�-�glJ�vw ��Su�6PF�mHiH�}@�Yr��q.7�u|���F�-����A��]���-W8����6�WXj��TG�)��sGv��꘻6��:%f��z���hk2�]�)ܔ��8J��M�&�@�HkV�;�QU�:�R2)�X��nJ�{�sSiw[�A���a���mn�AJWu�ǥ��nH0�B[ʲ$Q�i�'AHw&w]�%��lY���0��`II�X;�p�Q����-���F�l�gS��L���%>�Z.	O���&�'e;���J
�ő:�cUծ�_bewL�ɇ��%��o٘�c6�
��Ӈ��[|��7%�tO`h6���O�;5�����%Ӭų#/~�2�n��6���l`����F�y{<�q�0� �bk�@�ɜn�Z�W�8U��8�49� ���_J_�f^Q۾ˡ�W�S�7ݫH���.��M�ݾ]���s9u��ff ��K�p��|��;��\�p+t��&�gV�ӡ��F�&D���J�3J�����P�]m�4X�f��3���lu����g>�w�yz�l9 �|w�wY�%��J�­:�-h��3Yup̚� Vm1�XQ�%��3]���I�X����a�nP�<q�6��r�ܧj�ue�UlW{NGR�b4���+y��b<�����m�6��&���gf+<��Ɲ�*�m��r���d�i�u�գ]��ٖ�ܺt��P��4qV��B�6���¨<����na��w���l�k A+���n��-�ou�D&�PZj/Ur���	��=�݂��4\�}��gXs����"c��D���]K���n�4l�+oV�u����&�&�N�u�v�a,��J]��p�m�v�\�bˠS�Lt�o�$�[�h}No\Mͮ�Ǹ];���GT爦�)��q�]]�L�xC����T�#X���|�Ғ��#Q�I�[)|�Ơ�r�qA�kj���U�4��8�F� ��f�.�w7j��o2���ðf]R�;/�㿊�d��S��{q�AX�{��O����[�C�A�ŗo���a�[�/����#`�$���PX��=��T��t;�	Q�ީwX�JcF��j�O���㽶��-nk�/��V��BӖ;����4AZ���Y�6�N�8>�x�2�T�5�)�K^ߖ�#o<ô<�5a/H/w�f�q�,���Kt�޺͒�e��rꌵ,�K:�Ef�β1�c'�X�8��q�u�E��JQ�\Q�OOZ%uu�m�pg�m,����s�|�9
�g&���-$�δ.�#G����3��T����<X���0$/:c��=�u�-Mڹ��pA�J5�R��m
�%c5��IX�h\g)ak�X�����N
)o͡�Oe��p�XA�va�1��=�.�y��gt����=}�R]O)�.�b���F�ax��d���Cc�}M�ύ�l�[�bx̬V7f�,K�ǫ���H���v���q��{V(e.�Mq�θ��
�ːMQ���j:D���@)��i�Ų��P`��{Hc�മ��d�����}V㡅���&'+nL��ݖ�F�h�]�A*5����}Q^,�8��F��ξ�Kj��o��=��-VF0������z�V�ˋs<��dۨy���=�#���5��M�+z���[� םĩd�m�Z������R9�To���Tn�Ÿ��x������ �*�2�`�����u�oT8��.�8'_b7\��v˥�Cf�9eu���D������O{@�x�i5���rܤ���lm�N��j��SY������2��I�⚴>��軦�N�)�P5���`d�]�8Wcf�_c�ˎ����S=�E�R��4�6z�$4�Q��]ӗ��9F�,��Kn�æv��e>a���8x7�)��9s�Y�3J�Q`U�k0N���D��7�a���v�>�a�sDXҖ/�U�VU>��lU�m�Upm��yZ��Ja%޽�\�Z�u^E�����K6��Z-�]a�D��;E\�Ԯ�;�ʴ	�%��Tx�X;�o]ʻ�S�)jD���V���Os�1;SҸ�5��8v��u>��A0�!u�M��.Ľ]��ɖwz=J�Z�N�fV�3�6f���z�X77y�,T��}�T},�]�8�hj��D��E�V8��ZkP��R�3q=1Z٭Q���y냐/�m��V�Rƻ��X��ܘb}�,&Dξ_(�Fi�ӯ �S�Ę���r�w�x�W�Z�RGm�؄}8I2�4�q��iX�5ΡS����Μ�N� t򭕑�@�v#�j���U�	\���E�e����}��ɂ�hVVѰ��Z�\F�:�����n�:ӲJm��1w�#����I���]0o��뤜���U�Q�갇Iu{��m�K٦�BP{�7k+Mb�j־����ui��̓��8����e�R-�z�ծZeWY�X��t��Uv�x��u���(8��l�J�����vΡ�C/c�t��.;�����Pv*n<�ܣ}[�8�TmpAa�	L�<7;�ǯE}k����BT�;��91p�F2s����"���F�@�oX����`<�w�����(GI]
���!���6gT+B��<<���[�U����U�/hY���"�]�|��|�o|"�ٔ�ź'���-ӂ��%�[{u�"|%xf=�e�k	37�B�m�a��TS/Q���S)*ot��K4Eg'Q�J볜���Ί����p��ɭމ6k���vB���B0[��;��5vg#�"���m7�l�P^Kq֕[v�����Zh�;kiu��Q�)���@�Чs��Bt�yz���R�#��+Aъ���x"��ݩ500�p��S�l[ȹdɎhϥ$j!�6�MZu5��̡#�vR�5�Z�U��<�Q��9�g���i#��G �\��<*��{LȲfS�Mؖ�ī �2s�����+ڳ�Z�iٖ�7��"��.�}s�m:N��5��+`}J&�P��+o�q�Ԛ��[�{)9W��{O�t%Y3;a�9-c�EV>V4b�]�����\�¤�;�����ޛ�M�b�c��	�P���,���i������+A³���7�|���(>���k�X�M�OM���n���M쵽gc$�%���L�y(�n�x��׋^�0ԧ�mǝ�����÷K���wacxgr˰��eC;�̫$��؉@��WU�"����V/'���a.��e�u=��#�)�S���̡�q�`Н�s+6���!�9
����K�@�b;ч�u�Z��@�u�o�M=u���2ĝX��xY�_�Y��"	kKޢ�#�DG>3+.�Y�-*FZ��3��oY��v�S�Y'L�tc�P��ѱ�Q�wd�)��u�����Iq����ek\���e�l��w_M\�ٹ�v�;3�l� 5ov������^������$�D��R��ڊ��wNN�a�f=��f^VM���̻�HU�@W�s����R�N;L�6�ګ��x�KD���N�s��faz�n�w]���ߥ����)	�����I6�;Y�q��sT;q��P�2��D�J��u�%q�����.��ӌu��EW{1W
�:
��t�Ͳ�Tc(��"�w�ᓦ���]}v͠M ��-=t��wB�V���R�R6;��v�γM����
t����l�j����r�0Y]�N��4__ ��Z�&z�f��DϷ��-���x^,���̆
�V���e�ij��Y�A2<����f����@(�N�g9�E��t�u��2�P8O�]�&f�s�U�
��Ȕ�6J��oN
}݊g^r��'Ygq��(�����ʾS�܎�9��b��������{�n)t�xjaa�t��a���K�D�� �4+������7�u�p�SNʺEQ�aG�{\Op�K�졬p�X��O�Ѯ�+��m��" �*w���^- �l�Z(�u���mJR�
�{�b�@�@2��̮o��E1�Rۼ���k�zQ�O�\N]�uH��X;��&�>ݳ��P�hv\���cN �g9`2T8@d6�����28Tr�������G@t:�큸��n�w\\�)���M��4���L��N{Q��[d4�s�/+]ܾ�E���RV��|��p���ӕ���Z)ql�.X���+X���Wyr��}Y¶�g���3X����h8�&;s�����ègYYw�p6k��Y�ƒn�>U��GY��Ш}cl�]b�uK'Y�_B]؇���V/d\X�)���������xψ�K��f��YP��6��2Eӱ�S����vk��U�l��k8�e� �(�J��!m���,=}A�������gB�-�W@�VyX���|�-��-Y4�d��5wR��V��|���������Mu�Z/�)QRE�r�]HomD��j�Om��*^���e����R�`V*���;��P�)����n�E�sR+������a�������ZX��U�e��j��1Й��5��=uʷX�T�>ǆ�����֒����Y{��]�B��u�u&�|��pC�8^��7����������D��rt�����$j�����Z���hE�L��ϦR�-�79S 
���>⺂d���v;Q[���J�>�EH��Ɏ�� ��ތ��	Iq�N�
nc��$�C`-�WZ��ǵ�������O*�w�����\�h��C��P�X����|q���Ž�vk�g�5w3(g-�����+ܐ<��&��F��V�5uvƻ�f�5�ҫW�#qCW�n>�eG1��d�o�
���'2#H�p�^u_ε+;3{�ڻ�J�mB-M�L�R'�7�$��E��k�jƪ������27a��e�V���hfN,��6%�m�*,yt"hpW�LHŉBk��:ƾ� �s��^U�9>l6�=*�,i��U�����r�&���<��y=!�����ŀ����L���M��ד,Sѕ:��[�Vd��SNĞ���r,�9OK3��v��LB��m�j��V2n$*́:�L��E%|.evc#�������,vW���N݃)XW5�y�])pF�Z99�_��]�Vmژyh�|��\a|�y����/g)n����aO^�T�T�d4���)Y)挦x�Lj|�l-G���j��H����;i����s��*�8�B�x4���ծn�v�V�'�v��q��t�f��w�#T�2j&diK���0ME[�
n��r���tY9|�v�9i�ۻzSʜ���oIU��l:چ=����C�tXX]KY�Ҷq�V�/+q�J������|��T�����3��x��z:Py����tg��e\���p�ʸ��^gJ�]42���\��eK-4� �,�ޤq\ ���T1Z|��읕,+���\/5'���.�l����B��̕��aՓ3�\v�d�2���A�?��^\��|�eE)�v��]��x�ַ�'Ӕ�I]<�4���Y���gJ�KS�Z��]傢�k��=jK޳tNzŒ� ����4�r[�`bv�W8�$U����oz���*H�Zú;H���Bu�u��)K��`}�W����,tQ�X�^WqP4�"K�������v�V�E�9�`�W҆I�G�F��I9�Ce �yV_ RK�.�6��L�Ź{�3�Fv��(�޷h\�X�4]�6�sQ�`h|�1(A��a��L�O��hm��� �ٗ���n��hS�|��vPf_N_t(ZOs]!�F��S����!:]^;���)K�ҧ�X��2�m%�`Vi3z��M���m��#�r��kfک*�Kr��Ω:��kQ�����ic���Y]��S,۽��;u��N�\.c��)mn&ru龆��`��Mp�X�'+%��et��[���]�ĺ󴥮V��LYk�Ӆ����]�((P�%I�X�bQ"�J#�Z����(�:����n���v�a1�z�=����P����X	fo��u����enR�(6��:�`�Ր�]S���]-C:@�y3��9���Qk�v���a1�L���Z�f�.��Y��Kp�X^_2鞗�Z����Y�����z��l�"溽����}Jd��������{w5^Q��S�Q�������6�|��6���ֲ���'��A���k^��Q�o�5ɬ�mX�csm�b�q�����q���+�~��۰�SX�J৒�"�u�T��mKTETE�բ pK�I�PD^é~��Q;;5ږ�\�7�K�b��[�ԩn��;t��V:��l��P���F�Z'3x7+�F����L��g�+$�f	�TCng'l5�TG��	u�0������m��%������Cf.O�a;.�e4�7�pj������ʂ�"����Sx�5�Վ�z��Û[0he4��X��f�eǹ�a��:N,X��d�pҶU�	Y�+�VDh]B��Tv�j�G`;����Nx/7Q�3P-��em>���S(���'�d�Kb�n��ޥx�ͱ�V�]1W�Ʒ%�X�������̖z�����``b�U��7������Wm���O��!�]�o�����zDr�)���fԥVk-	���8Ov�F����2t�y������O�faÀI�'TJҦ��}C��ŋ!�n�=y5�-�n��T�aZ4GX@�{�3�۹im���c[6qQ���&V����>���bӬ�l_Lj�l&�Z)��Iee-���r��%�`���D�3GsWc�ydN��e��VaۈGu�u���Ne�	���56r6^]\W�s��t_;��m��U�gfh�ܽ��1����잫�Á���s{U+l� �)vE�uë$<*[f�o�w3�1U`��1�.$-���Bh�"�b��h� �[(��;A��YÀ/����(٢�P3r��Ma����m�Re`���R�A�ܝ&7�eS�����^q�'*����6�$u�7����;i�V��%v�}�x��Z!���q��M�]{�4�!:}.8Q6�N�$�wi��i����c�E�-[�''KZ{�g���ou"i��Q��;)gp]�p	ѹ�8.�t����ܡj�qѧ��[\MZ�*�:Za��z�QC{��ѿ_]4���Z���t�f�{�)m��\W5u��a���PW�g>bV6���Q�G��řpXn�K)̄�@͝Ym�I<��{F�����\ᇢ�G5�ҎC�c���_G�F�̗X��dAp|[A&�}�B�1�d��C�K
�:�/�&����ښ��)�7�t_C���fr�v�7X2�5 ��o%�=�[�j�ft�"U��$lk��(Ƙ�r�f>�;�����¬�n�鋻���3����PAAt{@X��y�S��;)��Y�U�v�����κ���`*��b�H�V�@Pd��;��ư���mSͱ]kn����V�'[9F��Ԍf>��U٣2���ժ"(q=�N�	��;ԧ8�F��W"�-!T�'^�����3�]�(�s�K���]�#������1���>ֹͧwV\��a=�//x0tcI-/L�H�{Ś�r�K�Trѻ���f�b����E�Gem1�mJ��0_(�u���� �W`'D��ɪ��P�R����Z�+5��2�6��b�ׇXi"h��"�lTvU�c��m���h\M��Yt2�X��1T�뎝0GcR2�2i�A%F���@B侂邔��e^J�Vեz�� eO�tNT_��-�SuĉG�N�wt�l�2��Տ4P����4l��eN�ю�"��p!�bO!X+[˚��#�-�{��ñ���[�a�U������s/+K�������图�1�37A(��4��cj��F��6�'a��WԊ3S�����]��C���wط�d2�<�M�N�w��,��R��V7 xri��5u�P����e1H��K.X���1�ٺ(�i[5:��ֺ[��RȠ�s4jm�I��4��Bް�˼�v�p/������yo:�S4�a/d�kۺ�v$�����Σ�0L���\���X{��պ�&��
�@� <G.��ż��0YֺՔ4cÆ��W˱�`�ΟV�ݺN���A��{B ��͢��Ѣh���m<&�^�Y�
��!C]��4hv���fsQ6��G�t�(m=�]Hj�[�b�O�ܲ[�խ�q�}�ڽ]��}\�W.�t�<��v(6��75���o;�����4��7Azw���wz��a	i�mA���f��Wٯ�f�� �reAIRy�Z^�DN1W{u�KAet����,7yD@�M��'Ds,��:�u��f�mm:�oNӐ�̲itGq����:u��Q��A[��u�s ���,u!-�ܴ�6��嫳����F�e��M�U/V���j�e��#��a퇊4E!�6Ƴ���	�1.���'�y[���"����w\2oR�%p�a3���M}�`�+-��d,�A+�w�]��P�K�������v��5�)��*��[Ɛ���&��.����X�;5���Ǚ4�WǬfs��(޾�eN6
��	
�5��Ë�� ��ıR��k4��ys��^�6�A@�˜��
\�p�b�i�`e�=V��͜rM���n��`��v����U�uԩ���ݙ�6��E Ƞ}$�,�;o��f�TI:=Xӭѫ�R��w#$�M�Y�n�r^�y�B��Sڿ����%9����*j���x�ecH����t�������h�p�;�¤�;���
�w*�Nw����ڮ=Eza���Ȋr���Vqݓe+��ŭ���LH�AZ;r��ʕ�-�@3.7y����ʒ(^�u�{9�e���&��@����m5���vLѿXR�g,���t�
PjW�o'f��cQ�u�3k_l3���Cv�t�^�����7DS�ԫ�r�'i2f�U֭u�V��g	� �E�B	{�kQ�or�cP!���ϳ�Nx/E�z��	-���NT1ʙZO+oJ|-��[\��QRĻK�9�49���tk�Ms�U7;��C�Yz�<��.�����3�3���:�ܠGM!�Y�㙷��T���eԗܝ��٠��v�"��cʔ慪7͖�F�DY[v�bmIV�����5|�wZɩy������p8��:� O6U�2�↝��,)YD�'�N��b��C\V-��b�L�ab�b�{�FV]0Ì���읚(!3�ĝk3�.�y`��4m�Sf��罴��Sp9��QYh� ��\�1�l�Z�!\:n��j�٭=�*�5�v�PUG����Ju�|�K��TK�ԠG'8�xh�!42n���#oOSR��D�w*�6�S��]��.��G�k+��b�s���\�_JȻ��Z�oc�"%�3d�ğj+��v� Y��g��%c&��e֒Un�&���������%ӔHAeъf�sf!5�Q���@h�#�_A����D��:���o`7�&unǕ��k�m�3ײ�{�u��IXM�t$��o=�}l�+�Ʀ۬p%��S)i]�Q�b��(�ha��*�l�A2(�-b�s�Zv����k�wLO���t����#کM�7�v�ϐ�Xee���L��)S4X�Oi퀏!�v��j-hqQ,��}:R�ɹQH���&Y�߷!A��:���`\����U��\�x�;�u���Q��$q��S�µLH���ѝݗ*�/B�ΚZ��٭��ıOh��ى���t��5Y�s-x�[�����}]����-{�jԧ\O.��t�k��������(v^ފV����Z]�;�|+�����nV�Qj���"��PѮͣ�`�[zU�xWWq���y�VЁulz�8�qk;
����6�|���&M�t�4��8t�*uw}�s�[ys��{F�I��n��CB�F����m���YY&VJ�q�����f�#0G��+©�5aF�ђ�V&��y�҆���]�D���O���U��a��Ć�W]��~�`;U�*B�㳠*Z��f�Vvw�!�v1�c��
��Ċ(���l��@�v�%{�m��!�#Y4U��GZ�q�4�N�/��&t�Vڷ}|M'�Z��>�ʶ;Ɣ���,�:��3�yA
��p�l���ՙ\���:V����d�f�`�wI5C��|ȗDĞ��4jN"��ƨ�W��Ĥ��cv3�84���vr[n;�m��k��5]J�eִR1��BзcB	��0�do�h:�wJ��G�p��L3�Q�p�v;����ه�_��L�V0E,���%	vo���;3�j
�k��GS/��rm�T�}ԣ[2֜�/ ��(:])Q�E��+!
��d�B*3jj1Wn�D���il�xz�e��Ǜ@O���tL����4d�Q�c���M��yJ�-���X�h��]���Ʈ��ç�iI9��mT�y���r E�LJМ�DtcF�{xk����-f�TW�At��)e��ȪR	�r��ݼ�U�Y[��CT�3ӥ7��w_R��eFgD���݃����A������iKi�N#jaY��]\�y��*�]���e�.�k�wel��/�g.]}|w%%M��bkv���z0�\c�2�����A�s<�.O]J޳GX�n�f��٫�� A*`�`U�Q���q_SNs�!��v���lΔ1�f5�X����&�0щ5���v829���s�x�oGuj6k-�ar}����I���bg:Q�c=�.��]r<ɤ{i]ofn�,���+�wЮx�u���u�6��	6�M��W ���3�pW݈��N�n+hU���������e5�v��-l��fâw�N�Y���H�>�ƨ����	�{{����*���� 2��*d�"=�j<2��
$��a�)f"�un�P�I��7;k0���T���>�����X�N��������B���,�A�5�~���ѣ�nÛ�t��r.�n����)Q����W�=euv��Ӣ`���'Sz����|��74e��A���(�\��WZ�n�
�0lU���筌}pn@��p�+��xr��G�� ��t��]A-��+��u�E��Cػ�gN�XGa���4��V7�b�'-��u����ib��p��{	��$�v�����5�����h�q�o��ՙ�u�҉�Ů�dB���2�1��rW#/w��
;R�[�$ue���A'���v�uul���)M� G%��AٮI�b���p����}�[�v�ߍvYZ��^�uY&��ѢN@݁
���-E'gbݕ��)w �ł1-k2n���ۘ�ح��,.��l���ƒʶ�;)�+g1�V����H����B����K��.��&�e
�#���@w��5P�o�и��N��K�[�������.�wg,<��0ǅ���9�n5}V>r�뺊:��CF�+��|pv�5.�y�mY�cΉ<g�v6RU�j�+�jefd7\���Dv�̗�[Dw*��b�s]jڵ�%f�jB�,�u�H�1ӫ̒�.��%r3sc}�O�E#%㏫op}6]�;+L�v�9�b�X�!�v�����˺��W&�3�w��ֱfa:�úoos�P�h�M�7�'�݄�����Se�M�4�H�ɻ�m��Z�-�}u�*bDoֻ�f��u��mV5�a\�uY�5���m7]Y+xP{��-e�>�ٝʮa��9��ң�7.��>�ةص|��وń5W2k9s�>:*eB���f�;qZ��h�4���4WQ��\5g���o+y�Ō����Wo
D��8�Y��62�I�9��<�lgGSz�We'�o��+��'8�sS�7���6&	��k��O����k����L�֛����G��+��Uy�͗�v �Yv�9�'[�K�u��Sp��W U�F-L]`Е[�#�1�D�(��5�"'ڱ�!�Ǚ��Q�jVM]��v\�Iq�ҾuvjZ��zܙLfih�!�� ��m�4�4��'NW�v���LW]��Rr!�P�̔@��VQ���ҷgC"D-��ƪaL�n���+�*��n��(N�8�w�e>�E���J)��o,l��w8���T~UxD���n��T ��>��f1�q�q�
ӞH^VN=O�G�Φ�]�N���-�x�����iWK��Y�Q�:']�8���r F��ќc�e�%	��հ& ����	������b�S����Py)�b|\���E`�#� 琮U�7h����t��$^-�$�:Yb��)�����!}������&5���zok��K�c+1���W�s
�������@m��kZ�5^Z��@Ѣ�Ή�������b���:\}��w�7G�P�$:Z<�j�B`���b��'3/��u���/�)��p�f��D�8r�ֱw3^R�2���U�����c����k"6h;��o}�iѶXL»+`.���:V2��KB$XѾZ����h���˥�ʭ�2h��)o^�׼�`k{!��ݑ0t	8`P̰�[�c����X͵��(TlWJ啹���$j�Z^G���D�RSw2^���!��Lb7R}pe�f��Øm������B�(�n�֩Ws6�]$��Y��+����5�,�}X�Dh�ԭ�沅���iK�[g�R���c�E֖E�e�\h��t3:Gu� .�fuF ��0�Ȩ�˒�;ϐ6+�``.������u��l�/����ɪ���3�`�����v�S՛۝���X�X�p��jzNδ�!E:�6�Zo�f:�PDX"#�
E#�|������y*���r�vNjK��fJcEA����%7)�TlW
M�����*�x��J#X�D�J�f�;^J���܍	c��y��R5К�u����ZE������F�tl�i!A�8mY�v�6m���Q�5C��ާB�E��8�{��#K\�8e�<U��*����D �5e+��s����r���	kE*"�>Ǐ�"�/[�R���ǽl�ч�7;!��|ٽ�2$*�����]:��0Hs�Wiҹ㝙����ݜ;B�
�Ղ��VZQ6+(G�ފ�C���W��y��^���P&��\V�\���5����򮡤�:���F	W�,u�x:�6�X��ˋ�fσ=��U\�Y�:J��)��]O6+��	o�ޛOT	Ag8^�D퉣�S@U��W��8�F���r-�4�5yY�\9<]��A�WI.�L=�[��J%-_!N��p�4*��ޜ�z�)�噽D\�V��hp��B�`�ԫ]�j�K����,�r�WlĴL���e�S��"���x�F���'��2�p���\�=��A/c�Mֻ��cWY ��a���t�Ω���s9JC�RQ�ݥ%�klp@���T��ӮwJG{lPŘ������.���}C��1��/4�.XxK5�������C�ܥQ塩��a�*j[���:� �.�J���X���t/t�Iq�����ݕ��/���'Ltq�3����l}aq�S]x�2��ֹ��]λf�#U�ϳZ��^���qgS�UUE���b��ц���LJ5X�m#m��L�T�+���ؘ�Ua���5�����I\b��5J�\e��#�X��iĘ̲��\��U���*37++Z�Պ�j����%E&��*��%�[�.UE]\0im��3%�6�����Q+[J
�U�*��� �b)�TL��TUƎ�u]b&7."���"�FL-QEb�n�EM!X�YE2�+Y�Ynd1��Am��k�SN+�k�V(�"��j��E�E�]0ȋPӑJ�UAD@X�q�M,[J�E%lQj�LEuA�1����kF
+mb�L@����%SE�QV*阘#�Dc*X����T]!�,"J�A]R���J�DUFe*$L�b��2�Pb�R�Ŷ�b�[q(��I\J�.[��0�QT�6���(��*UEeq@Ʈ��`�X��W�~�6@�v\��a�ݩ;�2���IV��D�r�'h��V�q�b�\ir9%��2��[�g�\/����I���T�
���=�w1B���R�q|�ӗ�I�Dw§Z;�R}�m)�q����P��NY��)��21�p�{(��j�r�;��#�����z�b�n:x��z��*t%Yr��0����U��e<��J�53�T{���B��<1۲��&�ٻ����D��ml0�F#D���_��O�L�]�=C�!HlF�
�_O<��d�>��w���!%`�Wy^3�ra�oAU�*B�e=�\=�kS�{�Ԭs��T����F��!�`5��A�vje:Qdu]^�]ո�V���b����OMy��|N7n(!��GE�Fs�c]ϹeNVV�ڥ�6�x�u��UZ1�W�[rЭz�ʅ���'�1;��ʙǵ�.rf�O��VЯf�*i�7�z�V�����*?�_���u������\i��)�뛳Ǻ��K�1x(���2;c\������n�'´#y�lMT6zX]�sC7�ns����Z�˘w�%[��q3� q�t�Sa��7�����8�b�����;`�M���a{�nU�a�Y�o��4�p\g�]{g^�j��tZ�˽�rz���'6���V����~Ϸ��}�����J0GY��]��SJwi�uq6���ݜ�.f{dnP�6*#[�ǁ��SO���}��d�[I�w[O��H��{W�Q�=�@����R�}ou��Y��Bj�1S��gX�"�m����#���	��pq��gս�6���-H4�*j��F'{b9		:�}0����Q&I��_k�Q����=J6<�C	[�����e%r�kМ�^�&Z#�ޜ�:.�uu,�3��9�dr.mV��1��n���l��R���0e\-�.].kw����3��s��B8d���	ds�S,DV��L$�����Cm���cXt
v+�Y2L�#�+Z,O	���7� �bO%q�A�k�CT��*dd;�٢�Y��i��[W��[{B�����6[ȑ��3�
�]�h��Zmiz��e�a˽��+gv�HR�"qp�9WBj�(i��1T�HS��͜O7k�M�������{=Ƴ(#�q�ޝ��C-�vCU�2`���&���8H��+�B~����C�A�Yu�g��n��	ƃy���j.�)�G����on���8����9r��#�3J��k�������$=W��aql�u���U�c�*��,zvc#ۙ���#m_��ϝ92~��^�Ȏ�Z}Թ���4���ͺw���q[��a��Sxn���J�93OdSBo;Wґ��Oe�cY���S݋R����\��j߼�xj�P�Aa�y������ow�T��C:�I�-Z�.w�+���uϻl6�)�[]#��"(ts���]ųҞ���d^e��t�G��J[M:s�ߥ��Z���U��C�S�qԖv��]�ON�-=C%[��M��s�v��7}�j�i������b���]Æ�h�WHq����byרL^	�:E�~�x]��V�7|�9/ݵw�Xϓ5<��@��>l$�3�4kö�Fn9/���f\�I�'��{*�����3�e`)&��i��շ+��غX�Kd��W�ܸ�YsJZ�:�K4�~}W]�J�w��<^��s���v��t��Fq<'7{l�c�S|�&�IFS!ȴ4��~��E����S��O�{U6�5*�n�X��(G�Lӿ!���r��� ��K�3����3�!&�X�8�gDw8��Hi����6fn�����s"I��̠��;Y��V)�*��r&�'XѸ5�������+$�z��F�`��4k�X�[�D�U�]7�����j��>�үSW8�̉��V]���E\�܊m�BO�;).[�z%��q�W�W=^oۑ�n�Y�/�д�3x�F䍵�.^d��u��Ud��ӝ�ins6)ǻ,unw�X���՚38��0U����3ˋ׎kn�m��/9h�h�Un���������P��u�xh���{m�Ruؙ�	c1��F&uؚ��!�]�2a�jc��[Or��Klw�.����S������'}�X'�}�wRZ���n����E�v�p���(�V��k`0��r1��9�p9���:`����[ɸ�Y��Fz��Rߧ���K��x�?��H�y�48H��d��K��Q󤯃��s7�3�o~2^�n�N����j���c��K���0��9z���TӞ�L�4�
p��=�Wn	��}�h�SNw/�mHe��A��%m�r���\�&2�=�~;U-w4���Lf��+�\�J�_�Z�47�(�<�=sQХ���|��^�fl�uJ6�d�z��VM��w�1�~�E�6*���uK���%�շ7doK�jEn,u�-eK�J��)�H�e��w�^l�N��5Ԅ���ۗ����n;�l���x��;uׅ
ڪ�*u(٦�#�=��:!�B��7�Ι��!���Q�@��)Ng�|��Oi��pe�J�xN+�����>t�R!]P�b7&��Do ���v�3�Cbt8�o��OJ�Ul��w����<-�u3Q��}�� �V�Q$!���oJ`d�~A�l�|�[I�7��#O�c�vurM��}`�w:�M ��Ng%!�%2g��*q2�s䫐R���i�6�����!�pe�c���(p�>���J����j���K&2���ټlp}ng����T>'�Vc�O؏:=b�3���)s��=�ŝ�侻����b�[}O;UO-y��ey�u�*���z���`�������<�bEM�/�y��u��ޫ�<���s�+ۋ�	S�XKs�Hܧ)��Lϯ������H'�����t'"֢����V�'��fμ�6i3�1"yQ�w���i��U.Y�3}�nyf���M�g���lϜ�́��B�#\�}�qC7H`�YLW�׽w:��:w�nB|��8܅�K�;���SB�Q�n����К������/ ���6P��i%��tq���.%Z�"�����&˔��a|'<=g��-�__zdޣT��~�in�$�R���o��B˘�H������N���ٴ�"!gT��l��E�&�t����x{��#�Pt��m�w���c.!�*�Y:X�iݍReA]��L�[�[ZM��ح`Ic���%��)#�g8��y�FV̮�&}��wo���v�{/�^w2���0�؋�j�K�mZ��{((_u��4���om�RC�߶e`�;�1�j.Ϻ���NqS*z*9J�zQ�km�gK�9�e[p[R���:o��T��NN�����/n��J����@�)�������d*�:IN�V+��ͬY���*ͺ���0맦s
�;xM&b�@����W^��0nW'I��Q��]u;�B�.�4rB�XY��B4R8e_Sk��^Ƙ��m�xʐ��C{�(Wix��9<4�˛���0�V���Y�ػN�JY^44���P�n��tح�#��Ȏ���]fv/�4�쫨���˛�����m�e�7�2�hM�rƦ�������μBx�I.Ԟ�}�1��+;��X-�Y�o���C���!��^U�'��<N����Ҙׯoͫ��ջ*���2m���滄��*谪4��y�~�㳲��������]*�@"W�?u<�"k��Nt�Į�� �X� &�Jښ�>6뫶�*����=[��v�䔜�ޱӜ|�3r�U�e��c]*
�P��I4��r;3d,a����&���X֡��f��1����{F56�4�Ny;7"�iܻ���W�Ef�(��e�#�����j;OV;t2R�8<��U�]��XFT�X��n\ҋt��ࡱ�JVh�C�s�/q<�����Jd%S��M�T���1̲���}hl���G�X+i��F;�=����Uhu.�T�#��QS*����L�Hi+4���vU�r�*ڈ�'���ӏ�����|���`�Jy�(G3)��޼2R$���oU��R�'*���T�L�`s>ǆDkU��Zwe2�fYh�sz����XΛ�%��X"�*-2xo0����n��ɝwt9�*	i�\�/�Z�%��ٵ��^����	�s���K��j�k^�ݮv�Yn�V{�x�i��z��>O�B�0��l�B��Y�q���0�[u�S��D��{ݥTq(<��2	�j�>z:�l7 m(oy8 (H1^���A�ՖQZ�V�8���*��3��|�7�.�>ps �)�}�������*��w"�u�(t�:2v��0oV���X��U�����R���'��a�0���=���X��$)R������E{-�C���U^X�--ۛ����\���z��]Ԫ�bX8���%i�*S��������5:�Hl�G?����yw�%����������OT��f�J�tc�m.�l7����ތ���=�{q13�t:Gp�;,F�B��Ο������<�IA��7�����]�=��:K��z��\d[��!�x���.��]桋Wv�Io&��Ç<�s�9$���+��s�k"�3_-�-�G�������5���WW[�t��	�[g=�3����6��a��&����SN��=zT��}�&�IT
�ת�2O����_)�讘�m��Y����a�ZS��5��N��L�8rҘ�v���d
��*'�rD�������Ɠ��)zJ��g-�,5:�w�����%]�r+�Ю��M��!�w94>h���"�k:#;
���h;��!��է_Y�\�7_^@��n٣�'���F"�*s�V]gy
Z}�ho�毉3��^�;~�P�V�'LԼ�� �qV9�xN��d�klQ� �a~���W��nN��k�E��h;�fp��C���'G"�9��ofjvx�j���>i��<"��E	f�������o��2w�i�뜼4C�Ʀ'��A��e�`5���:����rϙ�'w-ŪS�Bnr��{�����j�k�ý�mw^>[J�gL�~����@\�C6xW�ۯu����ǚ�eNF�l��{�kg��W1/H�;A�f���FSsP�մ*�y�N|;��U�4�x�j�B#��{�A]m�nC�S�n20R"��i��q&\�v��]�Jj�.*�*��z��d���4+(F͝x)�Rg��h��b}�}Ogf������G���$^�)�B�D��#�^Dp�Boh�`�R��(DT<^^_]�)��B�Ҿ�Z��)�K�ZՎ�`�#/�o&�'�/xM<�\W�u���P�E�3:��5�U�}y;��데���1�<�vJӥwe=�C6�A�н��XJ�l�F7;+k+�yo[Y���K9R�F��w|�	��PTMI��9<��J��a�f�0.��{�cѦ��]��껫�geAN������>��o:�ܵ����Ȣ�[�l;�����4�'���`-R�w:�RQ��J�L��C�+�ve�g�2_#���h�Җ�<h���h�z�樣ML5b�\#K]o+��f[��ytQ��)�6cxNBQ!�X��i�M�咺��`e��J�0�5Ύ���[�9����RΈiwW�J�B���Y �Iq�5��i�:}�`�%�mW!*�͚�.���7�]�V���Ԫ�ZƜ�6E���6�LN�CR�����E�S�.f���LvŋF�ap!r�5z�u
�ΦM�w�u�]|sz>�#V�1������8�Fo�g.�����K@de=�z�o:�U������n�S/��c�n��]�n�FV0c����j�p�f)5��Q�����㜨D1+;ڪi�9�2�Yk��Q	
�!���r]�pJ0�NQ�+(kN�x�g�1���;�;��X�B�N�\�����$8
��u��Bg4�)2m��sN*�"5DWVLB��E�����R�,�D+�Us�-�ѕ��lj�gi[}Vb�Ń`����.S��M�sM3x�K@-W7ܟǡ��N�``�8q\.������ѓ`�v��5aV��$e��#G��Ux���+8ګa՚_�U�d��m�\��j�L�����"����$�� =v��,:7\�RF�T� K̡�v0�K���[-�'1c�2͈#љ�P�`�s&�ۙQ9uFZk�h6,$i�
 �R��'58ҷ�i�sAVA�<q�#�T�Z��]k��f��S1��Ӥ[*�}i����	�WV���+6�c�>���;
���x�0�$XA�,���C�+C�zp���[z��g���;��h!�(k[gV�|����U�B��<��n
HU�9)��VWn���9�A�pk�}s�tH<4E@��5�n��e
|�S��j5c�(�1/��h'�!�����f5�E��u%��ŉ`�}��d���?��ww}�a*<��HO��JX0Lu�X�9v�
b2)�ׯt��ˏt�;�U�`�tu1P����P6�;����ז��:���	��On��e�MJ�T�qd}� �P�,�����}RE�H���F(z29j�
ǰ�;��O]�㽉K��Y!������I&k��i��/o�K��C��go�@]�w'��|/�\�4�1�*��E��[h[`�#-�[J��U�#AAT�F�
,4�J�ա�EbAV�Q�-h��UTt��eJ��m�(�+�Duq�DEU�,Z�աm�*�*��TX&�TTD*[\J�JLh�+�6���`�` e+*i���X�1Q�-�����3�UM%H��U��
#X�F*�:B�Ac����c!Z26�d��
�IP��̴Ī0�ڐ\B�f\E0���H�,X���q��Y\�DIZ��X������(:�A(�+LLAQY-��J�)Z�j��c1�-.���k��*���#I\��dAV
��f53T��LJ�\e�(�RŘ�+���&��)1
��X�jJ-k"��%�V��%nf��DM%d�VҪ���(��˘����{�'���T���ƅ^*���(�:體�>�f��P*�n٬���(ܘ"�a��ho`���U�e$`w��K���{�;�˰�S����Z�;��v��ֺA|�|˽B������V���볹،n����lȷC����0�E�mfS庖��I��ݫ�c����;��i�&nB���(|�dpݫ���m�(��ߟ�y1���x>Ϸ�4.T3�X��X� u����U�����\%Ʈkܒ$�/�c�D����'y�m$�y��F8�i�=abM*���P��g;�}hi�B�4\ώ�����[����-��$OfD�yOSԟ����ᢷ��2�pBغ�i��06P���={,l�F�J�;Lz5*͊M�L�!sC]nel`�TJ]!)��pksV�̯3A)�3¯�Pjɐ��=C�r�p�u�nh����9OMN��`�t��!���0�(vi��2�k]��5�'$c��.y������.T.�o.\v8�Ox|
�U�Lq��u�~:��m��ED�E%��Wz����;�g*��\����S�i��Sl��O�]��4Ʈ(��ft9B�F��N���f>�op���JW��p4vP���+�yk��U����[쩉��?.'�Èf�;Ԯ�[&��x�Z3Պ߻ �/��¶S�HZ}�M��"��\;W/��|��1�rc�֞lZX^ӝ�Y`=y�����C*f>��'���GǑ۫�[�]��SYR��3>T�صm�ro;=��?�r��FmO^�kd�n�=������ơ�)�V4s]-WʀS���m���N���޳u��v!�V�T���S&9�p��=^Ƥ^%or��j7!��W�z��,l�n�8�U�E��$Պ�(�;B;Oc���P��F��̨p]��ץ�������M�I��A[dw*��=�mc�� �9{�(ۇWR�Nh`s��7��;����+t�<�(�&�P�"�]Rռ��[���mz:��T1*ɿR�%�gɐ�%er���wOF,m��&].F�vby��sD�8]\m���*��YK���t-��̈́�������iTKm����ǡ�+�5��J����W�֪/b���Y��BE���#nJ}�l�δ�&FS6��Id��������F�#{(r�)�N=� ���v�F�:�֖�LR��7a;��g���&�3���oVӾ�F��1-�vR8�g��`i���`�D��Uw��¥_�D���؍9���Y��-�.z�����=|��g�;�-�6g��M��,�xB�T-âR箽�>��f��睦������Y���4���"5�D�&���*��u��9���:�$�ғ޷��Q�)���n����Y�7�:*=��;�����6��'���Ue�1
^�@e�k�H�UK�Y�:ޜ��̜$�p�zW9��J�W3%�Om��(���Ԫ����pu�y����v��HI�z���i^�֭�S}s�\SCo��ƫ�.�y�V�BqUʜ�P�]�_&����j�b�ƹ}F�w�9��O�if��`���4NfcA����g��n�L��%\wږ�]+7l2k\�.Wm�.���낫�*��O�,�1�r�؈���Ȁ��6v4W�Nx�(�sp�a|O�:`-[�}O�;���Mvo:Ǩ�����U��pb�A]=��xEo�=O��<�z�0������{+�y^ʿ3[A�}�ɴ:]-�\e�XxT�x��g�ڕ{I�K�A��٣�#��C��|W�q��\�>�bw���c'~����$��7���I��VM����C�3�zy�@XL��<f�;f�;7��htɈm�ـ
O&�U�|�7E��$t�@��>��Bd��淹���0�wi9s ��:��C!�r'M�f����=`u�d�$힧s�$���x� vu���:d�Y�9�8��*�н�u]��e��naW�~� ��>|d�$ї�;�E'��i�^a&��ܓ�Cl:�v�Xe�a=a��7��d��ރ�O�u���(�}�u;c��ϻ
������y� �����IX{��5d�a�������=d�j��O:m�������!�2`bx^2OT��wu]_/n��������Q(���,O��q'�1�Z��awG,�l;��E�o�';́�J�ɭPYY��O���,�&��Kï{[��͉��[���i�@��a���"GtÊ�8�]��h�9��L�<��C�����	�M_�,4�0��2�v�:5a�$���w�z��9�3��~���[ֺ����a�2z�$�`v�2qS�H��g��qX�o���l��L�>��@���9��'z}�>�d}_>�ʪp�������@�z`sV0��딚C�'���4��S�'l�I�^��"�i��d9Ւi�M�!Ğ�����v��>��>�#��+Kǃ�6���l7�m�^輙��|ҫ���ܒ�
ɶN\�����q<n��]�T����}�B�sr�@ϫ޽�x����,�]���[|+c�����ԩ�J��A����@U�r������m��:�[Z.7o�-ŝ���]�s}�{sx�&08m�q��>{2�vɞu�l��哌��/�i��,�~`$�N3�	��,7�$�7݇v���7�/�)���z��|#�t����O�0P�����3l��L�T'�i��P� y�d�VI�t�d�,��Rz��-7�	�'�o�u��!Ӌ���\3��>���l�#�k!���z��Y��{�=d�uϵ�$��=a�'l��x�2x��Y'�:�h���&�9l��t{������q�y�/v-|=D Ͻ��we{Ï�����i'�s�z����9��a������;�`i��c'�������u����==��0c>��qW<�o��޻��O��v�ɴ����N0�8�o$>`m��O!8�����|�Y��� �9�Y�$�<=�E��x���dz���᫨�_g/��;���7U�3�=�I>@ѝsRn�'�a�i{���t�;�ym57�5�6��'��z��1�z�0��+sx(m�0=�:"	�QU�w�]����Q$}�=d�P<@�&��Z�|����0�gS� t�`x��C�|��,&�珬Н�xM����5旚������xӺٯ���>��A2M����d�A`xɫd��=@��]{�B|����ēi�Y>d��m��>�,�x���q/�y�][�n�{���nu�ad
 �*���$�8�d��(�M���Y7l'�M�z�����4���'�u���2T{�0������Gզa��߾��u�'��s�p:f�'G�oP��i���I�&"ε���%C[��q&�ِ=��Yv��{d�M�=I����?����;��g�����9�w�AX��W�O���;�-X�Bm�Z�e�ZhE�1��5�m.Q96I'�9o�{wz��FM� �:���Z�I���z:�NEn������%��=�1I9F)��4 �2ӝe�֤�pZ�j�G+��U{W���(�O��C�z��tk��$�Vh=��6�h9̆�;T�S��q'���:������$�7���	ǣ/�G��=W����?�+]��������{���P�2 �����f�M/'�Vk>��,�k�2t����l��st�*v9a8ɣ����Oг+~��m�����:G�|��=d�&������y�6�h�0�N���)d�jn�,�O}�d����!�o�v��3~g��2������@X{ߛ�XLd���}Bq:2����'Z�� �^sRtͰ��l1���N��ORi�h�}�E'>�������g���^�W�t�6���8�x|����	d
�Y3{�ڄ5�2Vx�P�J�i���y6�<C��q!;d��T��D{��|A�Ʋ&~��7�}��yY��m}	P<O<�ީ&�����'̆Ӥ�L4�C�}�+�ۭ����o�'��'l���L��d���Y6�{�o՝+�a�S�<U/�*�� &�d�a>d�n�|�������xý��Ğ>�;߸z�����<d*����<;��Rt�وO$�Ҭ��j�ف�_��| }��H������N[�)=a�ڝC}`C��y���	������	���o����M2t�s�Y1��5���u}b�����{ ���{�� x"=L�r�$�'�o	�I�זM�n�<�	�x�Y�MM����S�<��������{O�����7�!d��sg��n���,�v�a`v�i
���V2��'���,'���v�>���M�=;����t�M��m��o�Ϗ����J��-4��]�l������Ι���ď����t�Ir����<�]ճ8#oN�U�-Y:��.�55�Vy��*ݴ��$xe��E��.è���A���@�̣�{H�����3qI|��m2z���Ϲ\��`��%\�����,{�5ﹹ�0�vs��z�~{��aXk~�BͲM�s(�|�-�I�'����l\�$���'��|�Rq'oXm�#�"'Gl�}��7W��_� �xi��m�8��'[̓�<I�q���OP�<��s�)=E	��i=d��@�o�M��xI|<��5�t����b_SX��(���(��>�Ǚ�� k8��� ��n�`i���s�'�:d�|����IXh�(�M�G{Ȥ�$Էh�wl��a���{�r�dW�����ۆ=�>g�z �>�3�x�і|�:f�Ϭ:f�'��wt2x��;7d1��0��&Ь�7�*,&�k�`�{l%������o:���7�~{����:٦N�;d�R|����̄�]{�Y�htyd;g�:gZ�N�m5��6ͲN��h:d��z�C�<d�.�� O���P�nr�����8R�#���;I�Ł尛�ԕ铚�m��&��$>d:�
��m��+$�>�'�T��!�i��!ĝ����/�W13;/����i)��� �3�L@9�!�B�G,!��Xi>a7�f@�%|d�j��c4u��C�N2c6��݀�$8���	RT���b�goտ[��(�}�i�:|����tɖ�Û�@�h��I8���aRi�$��靲t]d>d��ݓL���)�d�a�/>�/:�5ϻ��3g��d��v�]�J��s�E�����-��sx��La�o �
���iXN2}iP�!6�	�:I���'�>_7v{eeF�˗,������a8}N��'��ty@�&�8�_`C�ϼ��VI�u��8���;`v��L<���T��r,�`}�T;g�W߂��<�	�{�a��<v� t�K���6sU+4�æ���k:��g-@s�£�5�0>���~۳S��"��S�t�~loinK�"��W�:fż��oE��>��|`R�
�,lt㙑v�JK�w�� ��0Fx�һ�!]��*U5?��(�P>���z�I���ɴ�E�S��6��N����q4}���������C������r��!P�Ϲ~ǫ}�\�>�;�����}浱BTOl�4͡��l1���r|�z����m�]���ya��7i�XN�8�r�^$���>�2=���'w�5V
l㣿"�c�<�����7�x�<z>���x���P�'hq���ɓ[Œx�]s$�,'�yd�����I�06���$=Hm>�y��4�dg���W�����#O���ot��@�>d?�2N���QH����M�ćYa�d�Hz����x(C[�r�'��vO�>���}�F�gE�\�۽ެ�104�G�D% {��d|>���!�N�y��=g��g7�a6��`��I�u����I�ӌ���G��}��g�� ���,�UY�U[��u�~�߷�����M��x��w���;v�&���f����	���C�J�'�=֡=aP��|�qsX,�����dy��>�������![�hEUg�x���$� ^Xi�I��Փԝ<`x�|Ι�=�}����m��i��$�2b{�f;݊�O�o���0��b��	�7~C������i'}@�H�x��M}a6�זN0�&��v�Xe�d�3���~�v�:�}�l٤��I�,��A>�o!"��1�۳��=�*�)^Qd��L2���'��դ��:z��m����Cl4wI�;g���l'�8�f�:C���xxq�����ﲵ��1�r��s���g�
����Ę�:��q
ɭ��$��{Ȥ��%`z¦�:5I�ĝ/(O�r�gl��|ya8ɤ�{.��u�T�^���R��&�&~\!���u�wL�]���P-�ٴ�����6.	��5!?2�ztr�U�k�u�vM�����ݰ�_^��Ч8E��k�0�&W:����s+��;�ަ�5�Fi��I͌�%_��O����B�F����wgrh�P�S�nI��8�+�/�_�|o���!�m��;���:d�f�8����7Hq��Q�$���8`����f@�%|d�j�z��5���fvĉ�?3���ZH}Os.��.;��l�t�d�=M��{a�d�'.�8��,n�@�-n�q���o��#��OM�f@����|��4�ɶ�;���c�Ï��>���z�^Ӧ�q�I���SE�$Rq;=�C��6��2whN��jb��htn��XswƤ�d���������ζ&��{J�g~|$�>�d}��v�:Ն�N�h�xN���t�2q�IߖO4���$�&���s�$�:��`z�C���tä��7��w�9f�=��K����� �}�Ҍ=&�=¡�=Bq�2�t��<��2N�y޲N3�ORc&�d���I�^ z��>]>���k�<~�ssv-�ϥ�]��ڼȨ��� {��q�Iۤ9�d
�Rv�=��큇��x�Y;f�ިOL�h8�xð�&Ւa�xN2mN���l��ٮ����(g���,���>��!����g��'��|�X��4ó��=d�u9������z��M3�y�!�d�nA>���W�����z�c^��f�c]��]k����v��O>d�F���8Ώ��׉'�w�d6ô�����a��y'�'���2):CćYa�d�C�X2i')ޭۯ�����|��l����޲=��z��=�q��"<큝Rx����Ӱ����l�߽jz�	Ğ[���2s�ē�:�X,����X
�����H����:��sK�o���Ov��,*CĞ��谞�s��[$������Hu<���t�;�!����ϙ�'9h��Lf��� �|�6��ǟ^�L��fA��V�o���Չ|�v��tDB�҇� J�:l��QL��g�eI����Fa���	�~�ΈmT�3zq��y���Ek}�WX2�9�;[���P�2�q���7]��h�7W�}:+�������<<"������$����Bj��OY;E�S(@�&���I>d�7�}l&�ך�>a�q�؆�C�|�o,&[��a�g�=q��*�[﫡��º=��w���\'l6Ɍ�夜B�ÿ�Qd�CG7���Y[6��N퓫@�&�:�Z���9���$�w�'�:OX6>����ȋ���f!��}Rwʫ���:�XNy��N��s�rN!�&3����d�h�(�M����{l&���=I�Ru.` q�'�&π�}#�~ {���'eh��`�ϗuu���>I�m��5��'l�>CL�$��{��C�i���q'L��:���2T:�XN$í�{i&��@���>��y��z�����L�]i�U����Y�OR�앜Bq���2t��d�!Y�=��I:9�j2x�淐�O1tkxC�*M����l>r	��#���g��Q���$��^u����NMY>`mf��	�C���M0���d�q�$�
���d���2v�\�C�<d�aַ�8�P}z���^��k���W���j�?XM2p��t��s�����M��!�1�yBm���'!�����2q6񄬕;�xE�m:�s |}���]g��ͪ�(dw���T�ơ��z�Xh�|�XM�t}�T�}Bq;��;g���i%gs\�:f�N��ö2q�a;B�6�� $��ig�(����������U��ۺ�����
k�E_Z�-�˔��aY[˖@ݪu��>�V2��Ww/I��_<�y;�v����a����� L�xi2ۚ��X��D
��H8��"�g@�P`ȝ��1�����T�A�S�X�p�"���Wӂ�	KVa>:a)Z��#;����ZOM���@��w����M�|U*�-����;N`:a��o��5:=]���}����'c��Ǫf�<����T����7��/$߲g�ʱ�:U��0�ޠ�r���,-��gs,9���O 0Z7+u�Î��m=�x��l8� ���d:"��J����GFnk�=}J����׎n��@�ڳ[g�F' �j���B�9��8�i����܍����N�����~Gv�I.+�Ws��'�|��L���XϮ��-��;jSѼ�Վ�%�9���;��ub�4s���r��Z%:$ٸ��ٗJn��h
G%�(�>B8�R�����`�j�7�xW�����]��k��M��F��S���B�N9j��3�M�������l�)��"��Ù5�w��T���6�/v�j�Cm��}�볗�w;��9s�ԙ��nt2j�4�:�_nbB�#�뮥��<y"�	�j�W+-�o�v_N�ý8uX.�S���9@.u�RH��f�}�z'�uq;_-��X�+�*-سcM4�!)���~����ۋ�t�K8���z%�eEV��y�Z�
<ܢSº��/�Y�ʺ&��K�������ո2}T���}O��Q{s�V�N���%Ժ�˳j�V����q;7כ!n���6��ʶ����=��;�Lus��n����0#j��ܒ�槷8�e�)�7MO��}�5;{���.�EJUlЂ�JN�P1��JlU��64oV�(՚K�Y����։�h@,�@]4E&j"�7+�TΩd�.��WOdGUJ/Y�6���h��>�yL{B^7���X�hҝ�{yFPuv�s�a�-�]�́���2SK�L��YaMP��܏�k���:
��.�C��A�B�[ȭ �˔�/�}e�f�,�HT�U0�[Nɵ�������GM���5=�!�����Rhz7Y�I����\��x,�$mh[�h�:5��m��(�y#q��<�9�"0���lJ44��V�6'*��J5uۯpP;ʺr�r�I���O�P
��� (yQ}�;{�ookC�D'�0�G,iգ�(��VKo���д+77�k�.�IA�a}����.��s[�Ӵ�3뙙���1=C����}&%ؘ�a;������9�����[�a��|b's8Ol����E�}Էxt=/Z������Ι}zz���5O��[�s�ޔ�:n�d�ո��WGN�VI����<y��C���=\\��wfP8�}���~���k����σ�İT�;j���!�"ʋ*V*9KA�R�TVk(���(�ȸ�t�
�r���"*+"�����dUC�P�(�-��M0�UFc+YX�be��Q�P�]%CJ�&$��X�5Ӭ� ��et�TƸ�TkUD`�i3Ib���)R�KZ[e�R��ȱc��#-���ƍed�1r�)S)`�EQA��%l�0�&8�������B���][4��Q[Lf��J:em��-�b�AE�b0Q�iq����,ДJ��mƪ�ċ��Qf\2��չ��(�1�+U-U�Z���(*�*cQJ�̵��H���EX��Xjو���2�FҩmCYPX�At���%MZ�ڰĭ�����Y�K��"�E6�Q`���JU�UE"�A�b�TTF�%aU�X�,X�#�P��k�0� �ڭeQ-M&8�iiuK��+EX(��A
#8��?�gGFx�@����lͶ��y�Vv��ڙqm��pz�+K�e	y�u��,�&��Y��lJO��99�� <k���n+#���C34�݊����{�mw=��ά���Kt8��;�[#���UD�,~��7���Hҫz���ߟ%�����kD&����p(�o�.mܩ��I��H�k���v�9"���寻M��}��ČӗP�7�5�C��H��f���M6��+���H︜�}��5I�k��T��f�5O���n;YrKz�����Wz�-]ϐsm�x�u�9���$�h�͙)���"�^���ZB`���8�m�B�:���!�g��$��Q1�4.�[I�2�9Kg�kЫ+z�%7;�m��f��qf\Ѱ�+y�5���#v��u����c�PmV[�'��Š�d�A��s�֧&���gUz4��72���:E3����<8#[j�rq�C��6��9�F��ήFwJa:ͽ�WX��ȖIN��p�8�`�=�̎n
:��cǀ��z;�F�Vg)�Dt���`���;;��H����mM����im��Π8f[���}X[�̔�b?hn�=�B�bw5`3�i������ov��vþ��q|>ݐiR��W�f�ߣ�A]7�Q�;M��^�N�lo�)z�5�zY�m��ƭ���F�s��W�h�x��o�5#���,cD!>��S>��ך9_m�ᚌ܂��]���U�q�|��NVWKJ������@��ua<2�̛|L-����U�wM\�z�\�Κ��fu��N�͔(e�k��#������͜{02e�{�����j�%�y�����ɚo��(H��Ł�
�׹��ufuU�|��+ۜ��fMy%���Fͻ�>��C�ؙ�։�{&'T��z��u�W��wwk^E7R�K��S��O���Ǐ�svc�]u�讦����xNC��ǻ8jo��y��s~��5o�?B���{F߹����b9�Χ�bT��n7!_�4�h'^r8?x��.���ɀ�
�5"��W�������y+U��8�5*]vq�T�VhC2��Z�Ԙ"nk74d��Z������9�5�髪Փ�]q4�;�1
�ֆ��vȝf�n�csz�w-�2q!�c;�6��)O2f���W�Qk �CIw<y;�����l��&�WE��'wh����ENz�V��k�جK��y0�=�CY]*�i��Ҧ�O
�W+����`����sw}Q��t�ϵSڰ7�y����C�6S��z���Mr���?gtVO(������li�]BV����3&�f�".��ۯ���b{I֞�6(4�	LȄ%4+_�+�&�����qF"*�kY1ys6uq����x�A'���K�tW.�Kmg.�긦'	u��v4B���Ts�m��8�\&�K�0�:{�ۥZ���"Ho��yKk�S��{����+q��OOr�b)��{7{�U���Y�/����no%
�[c�U�������y[e�c��Z�ڳm-ۛh������S�iS���]J_����F�`}�L��ԩ�v�Z���y/G[V��c���Nj���H5Jn��Sd}ڌ*���hv3�q���*�eW>{���4�P����^��t�����N������=\��`�ȝ­k�+9����{Q! �G˟7�vvp��*�}��Mv�Ov-JÓKW*߽�yAgn͆�(>�ݧ~���!�l�[��>�RyBJ��d�Q�+޺I��׶ڽz�'��&�6m��wXT�M�Z����\z��>�Հ��8ݸiv�$:�rp
gU7�%k�I���OЦ�O �:E>=Y.��)t-�^Sɳ����s\��c�k6����-��C�p�^ب�"��\Vu=ĳ�j{12�0OL\�ױ����������xח�Ɖ)Y���O��+�����;j�V���^���7st���Ϳ%hi�!m��pZ;lɧ=ۼ���Ή�b]�R�SX�d�'P+ґ�)pu;�v�S����:�f�>�'k�U켪��@���͈N�Bg�1*�p�5�75�SJݦ�i�@�qf��+:E�����"9�@�b�O �3 ꌝ�j��^�B���f;w6mj���
L�m��-8lr��\�����f�����V
l��5;w2�)R��ֳ11ñ,)3-�к����Z`ly)R|�5�-کtwa���`�-h�z�=�+t���i���L��v�Ņ�y���i*�T"{qg��xz/q���%�F�h��pV;4��+��v���	��[�Sҩ�����Jr�a���fA�w# B���ձ��%�W\�~������:��8��1�=��i#�4��j˯(9��_Z��9ev�.�a����ުE �3P�q��ic�K�����V*y3�X�^l>�DWO-�ʺ�~(H��+�m��[��Yk^jԷ{��ץ_LUs�Vz��#�<��F192<i�X�U�hg$VU����z�[�y�h��Oc�����)�^tc�o�5�M1��lubFs]�W�F<��,�3�2��_C�wQx�}��-�t�ñ@��C�E&z���I[�����%�7�g���0�����da���k�
�vP����B⪥LwmJ��n��O.U���oS��9O��8y�4�z�w��(ob������MK��0>I�vLѹ�Q��G��Q̠TX쬐KN�Zջ�\l����w�X��1A�6%Q�5�[wͷ�OHS�]f���>ѷ����&@/o$]�n:U:�>��;n2���n�8Ru����9*�3�L�6L��fOr��{�������f�_|!SV*��j���S)�G06��� J��s�;��}���ه�[�?)����z���޵C���@�6ͧ�DWG�t�X���"{���[f�mW�S�ӊ�^U��]J[u��r՝/7��p���!�!���V���,-�s�b�%���V'��܇^�k=6+����BU{��v#�B��"Ô�7~ͩ�����v�hm��cڹ���Hh�3!��48N����*�ئ�:��9��s�����w�~ߕC�ǆ�"}��9@|L���8��y���kfk�^w�y����sժ�v:���j���^=�;j(85V&ۇ˷�R��5��ڣ�������� v��X�{;}X�*%\��h��ջ��n�?N��W�ҧ�k���Klf�yU��n㘡R�Q���4�)7M�"HeaQ�I��`�b�1&3��2,��r27Ey^�:�x���R(+�ӕ�}�ș�[�u{�`���63�ä�K'�G�Jf�%YJ�	 p�]ݠ��Ks6k�`�X��i��9Q���W��;�����հ���@�٧�D[����􍼜�W�l��Ȕ3E4;+=�jݷ�y�[���Ӌ�6�[א�Vf�YQ�b��s�Ca�7��h/	g���A,�w�3�ƻ��s��Qݷ�ڇ�p��>�G
�v�����h[�=�95U�����G�c�X����>N�fB�������դFcLhɌ寝�^X�,���z�W+��bY�5�nl$�M��D�A9"�n�5u�|_����J�4yHҨD�j��aU�Q�e�]�]�&ٝ{�1j_�L��~�4�-�@�C�z���g�8�M�ύt�Zg����F�����Ss��@�)�<���at]JڠZJTk���+W~�s�摻�v1��:����L�L��%SBӸ�r���5}��f6j&/u��Ub���'C�F��Lϡ	zsH�UVb_Z�7��]Fs���.U�`A��������M�]��Y�WN�A$�!�̿M�y�3H@0���=m��Ы�]��v���eoCE"�5]�$+u��-Ԯ��T�����7v�G�Ċ4T²�ݤ��/U��`���!��3VZ�2s9��W�{�=`�U��ʎ�ֶz��O��� {��56�)�l���F��~��=�ϓ
T;/��9�p\Z��s�q=����Y�K����3��yBU�:U�n��,W�(�u7��=����O�����c���q8՘��滊�k+�꛽�$^7ꝵv�ޢqΑ���,\^�̼UO�׉,k>��h*��f������=ɥE=aD(�ۍ�Ƴ�U]Z����eM<��m�L�m���k}+FPo|k?g=���Lmob�۪�P����FUs��[ɻj�ǟ�XF�s���\�ӥqO�f�]�l1Ll�I�Ď��ڰ��)�������4�{pg����3�:��(�ƤfP�6(F��"����ĩ�i��@�������J-�r�HR4IJ�<��:|!qT3m�%���n����UՏgm>9t��+��C�W��F/&�ye<��UC�[�j�:h�.�3�v�[�7;1%��fl���m�����k�|j�a�$���M�in�1�6��MI�رwu\�Q�����N�U�{�TҾ��<����oR�W�k��$$�h
}Q�������|9����9�z;���LF{�'*�S���{����$q2ڧ{x8�a�F� �v{�vV�]��a��sqX/��	��HC���1*%�+�Al44�x܉[�Y��Oe��7�c�TS�j�+�z83�Ћ�1ʓ��Pc��F���qli���W.V�2^nK�������r�He���91��Y�J2&J���<�6��W�弝��ALA[ɗc�F�#��M�|Ny�.����E\�ֱ8�����)�Ҋ\��Ջ�:[ާ�����c�Mfd߹�r��|�i��3�si̪s�ҩ��`O,Gi��L���Z��x�ͳ��v�{�̘�3����Y�V�P�B}x��H��[���>U���l?�Xg�]s�M'�Ob���|�ep$�ݢ��ϜWy怷CG+�7�{���
VF��Q;��[�α&��+�[ãtZ�OH�Ӄ��V-oh��.u������uG�+��s6�[�eeG��#�a���-�B3o���'fN��A����_ ���sE�Bl���S��²�6�zgԆ�M����^;]I��rtcWn��Ws�]�v����<�
��#������R]뎗u�-����T���I��K�H�s�9����V.�:�H�%m��\p�Йe\bg�}pKDv�Odڣ��|�8w	��/���bJ�9؍�*3�uC�3����~>����Ƴ����mT+�C3�~Y���n>�.��1w�=�a[Y^�h�Յ�r�^��d/h..b�ZU�t��vfߥFҽ{��ں9��Ӽ�Hoj������En��u��D��$	�+�nS�0��s�ۀ癔̻CK��s+h�u���΋�T�����[������3.��];I�S2�NЭu���%tO�b˸[��m�bmVm�Y��9�� ��F��z^<'Qں��������\:�����3B�ґ<r1b�u�q�n��h�C���n��{��{����o]��Y�aK.n_c4�r�s5a��})��h�c��9�����t䥡�@0s��wFr%�w�����KU`6��;pཀu��笄���E��F��5�bD�p�]�`�,��p3��j�/�f��g�&)M��q�cs�u���]yt�;e'�����V��J��wWncZqJ�+ ��/�-m=�
�Z\��������3�~d�ؒı�Ӭ�W���Nt�CJV{���d徂��-�� ۶%W��!��>�ys��]
�7v펻!�bji"��ԫ�]g���D�/����E*�S:�X��¬b��+��R/r�f����V��[��_&���(ZWMJ=}��V��in y��Y֔�f��:뱨�9����,�ucFr\��:�傥X�6�\�����eB��,�.�6��(�̻?C�\�QċT�p�Q;C�Hˮ�a�J�ʣ��iGVԾ1�dVB�f��<+$7�R�{GM�}r��)V���;V.*�6�rײ�D��na��.�y�/�WNo,���Z�+�������@a�(�8@9�r'���H�\B�pȊ�dV��X��ӌ�,���}����QӇ^��:b۶�L�Ҍ8'�&�ԸQ�׆��C�)�����Dj9b��]����o̪�����Bz�z���.����<����D�|�
���X��;���ʷ��,����Mp�$���R�".�i&���q��N�r�A����(/G���]@�[���S��(w���b����8��ds����3�֯�kQ��ޙ$�	�)�SoT8J2' `�IRըkw����74��BGR���u}�U�5a��'n��B 9yT�ᵗm��Z����w�QLuJ��Y2:�W1q�l�Nc'��&�+V�v��Jq�YP�8-�B�86欩��% 	��@XyV���p���.�ospjyB��YV�V�RucS�]'��⺬�������k<��;�=D`(�y�㗨@	�2���*a[�l��ْ��k̬g,��I�e)`�.��{�<퇵���#QvdX(�q�s�%��NV��vz�ٺѴhV��R'W��'�Mw�ee^����[W��!|�2�WP�&=]�Haz���'RvmR��촪,���n����1�a%mR���nX]��
$��3�����`��w�Ѹ��IM�ɏ��R9C��ǭ�:���n�d���|"��;��Y����nU����C���M�ӷ-t�3qN݋�)݀�����;ŹԻ/�l�'ğ"F,E�
�4X8­�E"�dR�U��QĕX���"6�Uc\q�1,�h���хA��	�,���V�r�[t����TE��b��aF�J�YJ�(�Tى�ŌV�Ub�B��B��R�\r*��(�SL
�U�X�����9�S2�X�E��t��Cm%t���T�1Tj����Ւ�	a"��
j��JV�l���������1�ЕXj�J�qI2iX�T$Xc"�����i0C(k&2�� �qF.���	J9t�"�b5�h�4�YD��[S,�FI[ZVV(WNlq����6�����c*��P��J��Ve�n�t�b�Y���Df�q��#�"�dDZX#���B�Q��D��XV-F�����UHcY���0�,��X(T�f'��qyE�s1���K;��W;�EJ��P���1����u�wa�����j�j+˸Q&����;T�w+I_������5:q98��U��t�z��1�����9��ǚ���1uyv�m9��5��E\�j��B���v9�	=4�fN�|�'���"f�Y�K���5���o*����L�8�b��إ�C&d<λ]�yr��Xk|��\؜�o����f�ba��̈��U��il���Fs�j���zV�c|�&i��+8+d�����O��Z�Z�f����z��^C��E�����v������^�'<�{/V����[�vo���h	�^s�ڎ�m�N���v>�ux]��%��\�Jz�q��W�*v0�c���¡���B�26R�CYk����#��S��2㑙�ܛ�u��Ȼ&�T�EM�\���on�[P̌�)�c������T#i��ٌ��ZV��<��<�����K��"�;���R�q����Cpv�1u�xD>5}0�&U�B��ϋ��]��<�!����O���}P��)���Z��}�F�t��˷�Љu2hASX3���M]yX*�`kCy�Cr�>���l	�U�p^���7�F]��7��T{0����䍛�+�d��=�=�z��	�o/��������W2��ٷ�b�FD-�E:�yV�!��`C���ʧzR�ak�GR��s)��d&eա�D.��%mU�#	Ȅ���k�mEm�����T�2#[a�i�.!KB�ئ��Ŕ_w��w>�4#z��P�Ub�d���S�M�!�uV#����YovS�53±���frzݺz
�Ʀ(vBڱ=��>h;�}]*�
����]�3�'|�K.���t�}�x�Ok�cF�Wغ:��ׇ��Nu?j�!#w4����s_E\���.[�f�"t�Cx�SY��_*}�h�I��Zݹ�4M��`r��+K��Z}a�h����Xp�u��ߓ����mh������8���ϕ��l�ڷA��®b�gM���{�rY�	r����E��N��(�d�R1a\��W<�W�~U�6�e<���y{w*+v�¤�e?kz2�f.�F���*T�.�*��hX�B����
�e��(�����&�a#���i.��,v���B�yW4s��Kν�K%JW1wZ�����C��K�K+/�	���0��KC����������)M�<ʔ��;j,MD���AN)䢶�aL1C$wH��=�ŃBc\U�<jԨ�uŸ�Y�x�����][;׽�JWs[�r�ftODP(z�UG�
�X>�ӊjz!�v:8�MtM����1o#}��Hkz�F9u�^(�b��pAf����M�qU0	�av��8���]J����f�tWP�R�ƩV�	܊��Nz�yf?C/���EK�9����]�.�Y��7U8F(�ÈE؎͘(ӌ��
�qv$��$o�PQ	��Ybw]��jo���gK4�>������x'�X�Tje�V��8xyC)���[0�unc�E<��J��JkL<a:�ݧ��O�#e�-	�|�F�}�K4�L`��
�{).����z�+�8�:��P z|J�]Mנ�&�뤴�b��4/m�Yr)F�Q�tҎ����u���0�X:N��Fy#8f�Fz�<4��q9�5���<j��˼�t۵夦�b��%nf}o6�'c_&z��ǨԠL���z볪��L'�ǝ�t��v�'�]�׋����3pLb��H�i��/�QB�8(��]��-wC��f ^��zj��57�`�s�s����+��=Y�#������=� +��g{)C��"bg�7�Fp�XMd"�eA���f�!�{3Ӵp���{�^k����~�\�Ήb4lat
+k����w���l�hD[�C{NϞ�D!��u��;7�8p�fui��,͖Xز�;�e�r�Y��w�W�p�h����]'��Z�7����	�;2�4R�b��ҋhm!/�W���~��z��8���	B�wQٰ�iV������v�3sP#r�0x��*"���p񧰭*��[j�(�6�Z=F��̢8��o��pˡ(��Qq�禰D"P�Ǌf�w�X����ݬ:����mH��yW+g�lM�JћwE�6	@Ї<pX����eA������̫ˋ#K�F��
���J/�5	��\C"
ٱ�8t�AО�p��\�q��c;/�'v�p�0bYE�#�LQ��;p��3HT��-��f�%j^$���B�����{=2���a!ZB�9~�,�q�ʚ���l8%.P`�xeU�9���ts�f��4�d��]K�\\��f`��F�i^���M.�7kN�>�y�OFI��THUR��`1��NEĶ�,����Ʈ;�X���ս�y�+wMvsGQ�na��:��G�i����)�-���8M����bn��o��ٳ����v�/�=��E�v�n�*�l��Pޠ�):`L����
x݉�Lߺ3a�7�[�U��ޢ]78��u�Ǽ�Uq͇�飀�r�2,
T�W��!�!�כXu:g��C
u<1�l�0��Ot�=#|�����Si�}�և�n��a���.a�xA��-&��7J���oW7��=F0)�����DD�y��u����1R�0fVd��!dg[˲�[p�S{�uFи�~8`ө��%��&��DLP��*zb�����Ph��<:z�8�g6r�^��Đ8,��s�T�����i��W���0F+j��	S�h�d��ó�<ÓO�bY�֋��b ���)"@�T2�Kq^͚(�E�X\���c�/7�1��7S]C��[[�XzOt ���6[6�2�^�.�K�0]�V�aW��b�{�ja�����Qƞ�a�kv+<��{Gzzk��i�bF�`�G\������痓��6_��q�]�G��i����ȵ��Y�+z��>Z���'���m�C���>�/.��̌�W%���e�ُ�s��3SQ�A3|	��M����v�����b�.٣9��MlˋdA�-��]G����fY�^�Vf�0� K=>v�>���-�n�,��Lᖻ����K�K�Ug-��� Y�,�۶�=�mH֐��_b�;��ݰl�ţ�)��{����K�����Q��ڄ驷D��hċ�^9.���k$����G�9wR�ي��5�C���X�.�gԼ���%���9������PpujU��$���a��Ĩq6�Y�����LCG�8_k3���yX����.�Z�NK�/)�ͮWg:��7��"ܻ�y���3�5.|D�8:� �zB�9�L9�1~���R6'��3�ob��2ph�/�ۋ�Iկ�����ё��1 c�
5�I"AGl����#���NH]�W5��73�{x�P�MκQ���ʊ�4d1ᘧ&a�B6#eH�}]���u�˃2�^RV����b��a-jd;�uVP�$u*f12�GD�������}�X�����(�;*���yh'{�)g�J܈�����{����ԗ�n�R!+(�>�%���|����e�4�ƈ���\�
l��5���/G7�[}Sl^�Э�Q%w`u�\Qz�.����[�*|t4}�,!��`|����zy@s�˷&��u)s�ݮt�J����78�v�!-���.�v�ih��٧����-�!�)�����Jڔ޷	�⮫��ۦ��g,�⺌�8R�Вͮ߇��<˾a��^{���9�ݮ��`(J:!\��d�p�o�=������Y*��욽�z��n�Z���`�/m(X��;��Ag>�R!oc�-
��&��[�����'�5��V>�N�dk�
�[����[К�����8�,5=�y�擪8�-y
�=�Ui�B؞4-K�l�M^N��eB-N��5�oU�z��&U>s/��'������fi����-�����^%ު��tz:s���+�)�x5k���͙Ѝ���\�`ߗ*���[j�)��Ƹ�E�\o�B5�qōR��4�=-��{ӛm�w���L�a���<�1B(�Tx@*�+E9��+`cӅ߇0LdE��&%�9!Ǜ<3c�'��oz�F�.���R1Z��x�x�I6"8�#�Fd
��x�=�͸�bt��*���w��"m3B�ʯel��y�~���v�-Ѷ�MOm��˳knw@�"K�(׎�2��=g	��x?����U)�$�h�}��U��"��H�����dɂ`"��S�}rH�gں?^���T]|����ek�HM�	����1ضox�J�%��K�,ј�:nS�.l����:�{�{���S�On�\�.Sd�9c;z���j\R&hi��ۅ!4-UJ�_{���-�ѧLA
��HN�P�Z��C�k�z��P��gN�5�:��.��.q�ii�y�*���Ҡ��q��њ�*!�)LdK�3���d�Qx!��gLw*E�N-Ɨ~�g�"�_Ҏc�ㄚ����(M:�]�i��u�>��Jb��vz�l�����Z�q��'b�O1;,hBu�g��"�(��$x_ڃx:��9)��l�{|�Ɋ���nd"�2�� ��v�RQf�04gU��0d8��)9Z^���k�*}<�*b&�,鼻�G2%����1�(��ubֺ؊)kA�K�i����v�E�{�7<gl4��{�U�Mf*�yR���,��e�w��>ͤ��̥S����D]�PJy3��她M
�Q��gWY14�q��(��E�`�e�;�DS'g��m���t���mJ��:9ݩ�<�v�Y�j�7鎨��>�L:�Dl��ͤaJ���>����]r{�F[s:F���:�7�b���H�'S�3�tR}J�`���t��=gUt�L���Z�r�<�m?6�kq�(L,A�xm�a�ͦ�WKɊ+x�9�u��H�_0z����i6�d7.���NdT�*-�}5�j���2��oy*�����p}W�_��3��gL!��w.�W���{�Uɦ�^^tq�u���ν�Y�[��3�`.o��.��OP��nn�&eY��!���N���@�۵�.��g��+�零WӚ��A�(f��"�P�]^ֿ�{������ȯl��~�t:��g��ሱ��[����g@;<�9��s5���/2i�]6�	.�mBl�^�C����8��w�K|�?	���u���G��#Ճj]�qK�Gkf_m�ͨ���F�E��5~�W�Nc��]�-|<��p�L�غN�fm�|��$!=Xj;{E��6��}ǉb�N����|>W?R�i�N�MT#�`�"+[��t=�E�X�d�E�"db��vR�zV`�f*�xK�g�`��-&�������N�1�t��?j�h`SN/ ��DE�1AYN�\E��T�����h�ϗ������-�,�>�[�,^V��e�Ӈ��M1l���5�N�!���� �;C��c=���[I{ �*�A�	��y�Y�sn6�JYa ���r����^����8�l��6��x8y��0�XO�����&��q�9���3�ӹ�g����[��'���ڝ��K�+8�Z��ܡX:�C�`�[�܀EbT�S�v�v�.4��M�����]B��|7ʭ�]E����{��^���컨�F�mn��n�;`�uƅ��
T2r�'�9x�����5���(���{��^�Ȝ�^��Ќ{Jݚ��_{�Xg�n����Q�TmE�GPT��RS�������WB�4�~Wx]�H�oϕa�kv5T���z����yn;�&尠�f7�q"�E�L�ң~�u]2'X�xp�H��+O�Q[��ٵvr4��&�)��w��I�9��R>LF�P�b؞5nIC%#2x�(�8��
U.�Y�|�n�T�N^�\�2��Ξa<P�%���o�������Ŕl
���D��{�8��Ě�)�5T��*uD�8�*�*�%lJ����ӛ����x1Y|�Ι@ޭ��²;�5�M.=U$�7,�#�L�ﴭ�|럗�B�,��)o�p-�p��&��Riݤiuڇ:�cSQiS9Q��Y�~�e��$dZH�Q�w���fOP8{'$��YN����ʇ�6�hSN�W{QI�)���A:����u{�`�H�/�W'��|����F�O��R��o>�nom��.k����r]����tM-�"J��to��2�z��ݕr��������6��U�]��t���"�:�2��9N��gP�H�X	˗Ѽd��)"�sgp�l-���\�����&�s�f����Vv�FtF�X0�H�v���&\t��G
�=�U�b��23�M���kC�� %=��a��-��;��m6��ƨcq�`P|(徏U_n�6LW|E`b�2���^u�x� ;G��(�t��4^Vg1�L�ڑ�����
�u�����w�IO����VS�x�6���_��j��Zr2(�\֧EXY!�b��a�T�;�[��@,n=���p�åu]"r2�V ��7@�5v�Y1�R"v�1:�hB��ib�;
�f�ᴭ���[����Ó�>5�k|��n߻MI-�x�7��Tn] �TC&��\��m;�>s��>r���jn�]�J���1��R
���:;��U�:�(�0��fs�s;K짶��Ζ�Z$;y9�Z�Y��Ĉ=�A8y����œ��,��ӻW����+M"��nR��=���WZJ��������G��PtL�7�1�8v<�f��^;����Z͹ձ@�Uư�$ov*��{ o �)�Z��Ss�0�B̭��E\y��Bs�k�C����7��J�d�jw;�Mk$�e�˨RHJBWV�ݏ���.=����U��ΏD�����d%����d+�!,�N��n-���4W�Y}V-�tj�i�u3���/JT��+�}O(���s��in�,��8ps����n�gY:���=��1ڇj�ۑ�HB������_E��l�@e���}��j}�()���	J��v��,���!�UNOH���:ٺ��Bm�5�^3��[�+��r{��p�7uޕB�`/V��l�)���.p�&f�˧r���њ;j�a��֞B^��.pZ{���1����r�ڹF���(fl�\���\�����BM5�tΠ6c-�[8���t{]�7��.� ;ǵ6�4Qy1듨��1��*�D��sp��VQJݻ��4�$(�X��ξ�omW4�
| �֝6yٛ�����J�Z�s��]��&����Ģ�WWm��M���1�o˻������f�vȞ5���4����o52l���`Y�|g7�'pЎ�����,��=��Q�$����+�B��X���ݼ���{��E���ά�f8�c�Dz�*�7*Q���h�$Yu�ֺ����ַ�ƍ�)�	v�c���v$�{�mMJ�]\g�����)�ox���ڷa�c��E*�ԭTu��`�'(������f�;;g27�hȹ�ݳڢ���g.�R�A �H�+R��\m�����T(�-�*��V8���ITbi�)YE���̠��[�%[B���J��DDX9���j�B,U �,���`��H�Vж�Dea��MI���Zܦ$U1�`�m�*eV+���V(��Qb!���V��QeeAJ�U��-H�Q@F6�DE�JR�R
6Ɣˌӧ31�V���*(���hYK[��L��[[�h��J��(�D�(�TX�`֨�ʊ���
�Db&dmmlh�����Z�AV���ժ��%J��Z���(�(V�QB�Dq3

ԥ�(Qm�LZ�JF�-����6�f3j�"ѥ�5IRf"��Ŗ�`-b��,��meU6�-aU�n����-J��X�PZ��iE
ыZʈ�(fP�l��m�F�-�f��ǎ^��A��.^����N�0,TL*��}�	��R�p�M���[��N�p�V��+�!�ͳ������-��z���#OL~�2鞸һ�8���؍��L���j^ċ��>R�\��S��
��lS�����薂)|�j,X�U�6UZq~��X����ȰoO*v��SY���Oh������m7�u����u򢾧�q��񺲇S���'{o�h�#1��?f�2H���1^j`ĵ��@���j����[���i���o��m��C���rJݕQGq�ёe?k ��B�G���r����yݡk<��7��YvUh#�c���Co��1+��rժ��@Z��b��}=Y�/uGn��]�DV���W��b��:S<��8��N�{ս���VCHǂ�wtn�@3�V>�K�Y0�78m`��F��6უ6Y&�F��N�|=k}+e���<�nP�z�w�ZQV�^�ۛ+����G����Fu>(����e�V9R����x��G89�<ϫ�NB�T��_���J0�
b���)���֥D#z�g�&�I�Eu`~�vd�;!��w�ڪ���a¹�śzui�G�hFm\����Ԕ����w����V�f̤1�W��e�L��sV���"�����s�oΏM�A+��xN��Jv_uf��Crx�椋��"�c�lC)N��=�ބ�g;v����yڏ�Oa��"�蹆�'LT Q�T+�!H�h�S��9۔��l��(Sn#J
-E{����d�{�j89u�^�k�:X<	Q����`Q��'��<t9�L���8®��T����!��d���\Ŏ�K"V�f?C4T�waz����o�Hә�
ʚ�c��۸:սmj88?�3Ɲ_l��|�
�^���#�<m3���Ԏ��]	~R��١Y���I@��+Al��+�>$h�kR�'�}ʾ���8�}[<D��'�����OI�>Fˢ��)�b� ��ʇ�s,�f�+睜����KKh죀�
�MK�b��4��t��g
�"Ϯ��=�����S�:�<F�L<P<O)��3�b�
G��Bi��8��2�ժ��~1sO�R���F���@̙��چ,t��Nz��	�{^�A�
�[c`��9�������`J�y(-�%��v�X����:E���hZ�,�����r�[*�Q�:�Ŏk2�<�mpDDҜ�����׌#��f��x�����r֚t�C����˷�z˩��Ե�wtLH�8�jL/Kz�DT�N�hرh��7�8yF ��x�-"lKs��ַDdܰ��W�.�_���Ed-i�D�& �ôT�ӛ�N��u��ʔNm2���::8��43w�q�4�SYS=R�k:��Mf�j4dj|;���L�)q�h��=�P�f�."��,���\��=���\Ud\���{<��G�wb�yZv�Y6d3�Q^(�)���8��!�����҈}�\uԢӪ��i_i֕�/䆞���*�s#kI���[��r,q�y��+��<�"˞T�y���ޥhͻ����R��f�����
���Ӂ��Tn`�4��D:S�!���Pv#�3Ne�L��#�C�.""]�����"4�OE�,�^�T���<T�T=Y~�����Ϩ!�;�[�D����T�P{�K�w�*�}Oh:���d���W������۬�6�y�m>��O2���3r)�jD2��[��zWVD\)�v\�W�튁w3�+���c}x�Z�Q�S�.�*��n$�;��L��H�d��c�JkM���z��9�hc�7�%xq��t�9�k1��Z���3��&��}.sTY��^�I���/:���P��!��{O�w���įY��R���狁��/�^K�9����w�b�m�I�yeQ\møs�je�N�j{bos̾ô�ڒ��BNNq��� �n&��V\���.�ۈ"\���3�Ve3f(*f&U�l�e 5���ث��/@3)��h̎�c�J��r�i���!9>�b��S��fp�T���FsYTLE5�<��:\h�!����F��덬�e��&X�[0D�1"�ܩ�V�H�#3������O�v�B�,.�A^Uq�����4P��,�jIp�l&�^���K"C���A�Y�yأ]�^5~�A^�����y9��_���U��W\�����`�+�Fu-..��`maT9�y�(�ԕnE5:c3)fk�P�r��Jd������gc�x�A��eŅw��
G8�o�a��.���'��pJZ��y\D\�
��1q�٣������u�X�xA6��}\�喣5�ɧvTiɼN*tN�5��%��72���c�(�^�'�[�GVR�`���eʱc8�K������-gqiX��un�k��e.L]O����<������ǘ������W�
	|J1Jm)ꄺ���QK6���þ��W��V�h�.*q�+#���A�}�W��qo�y��V�<�+�p�Α�j�w�wW
�{#(���j���쎵��x�a��o�<�ywۥ���YNus�����J"w����}��=����KYsQf�q/bz�Q�C��V�JQ`��R6�0�=������]�C���v�W}��u�gλ��PO�S�܊9�*c�������:�_m
U�N�	[�S�g&��U�n�s:6�8�s�.\��Uq��u۫2.f2]Q���scI����m藜�\MJ11l���������Z�sƯ��fN�T���4�0̀*1�ir'g"7��+:�h�V��B�pZt'�Xي��ʰ�Z����WB��֔��Ssn����w�����X#�)��ԴJ����X�JW������]��)e���J;1m�+^�j�h{M��n�%�.��!�S��,��ES�8τ�VQC����u�F&Ƭ�ۗZ�۲q����ҴO�#g�H>���q	��v�G�KNV�
�l��Y�r��o`���2P<^vӸ�~)��PM�g��g��B��ǣĸCazq�K/p9��no��VV��CH͙@���_�Ys�J��9��4�a���Lnv�֕$�.�z�\����b�ѩB3�\��ò��o	ow�۴�uaY|�:zrd|븽��73�Tk���<I��3z����td��;�Y[Voc��Zav+ioot!�cB�����	�֬�Y&��J�}�49 �4�-���������]V��n�}S��n�Ӓĉ�����)��8��V��p*�6\�d�q�ޝ��=����*˖	���-yz�����ґ�
�j����(ձ0�iFu�z��=��Oz,Ǟ�6��\��5��Q#~+JS�h)�����;�LU-�)`1ϟC���ֱ���Q��q��:}B�)��Ƹ�#�ڕ�����-}�Y��I�ur�oZ��R���(��Y�=[0�tO�@���Tx@�!H�k�qU<b�j����o��f�\�~�N!�6�3���"}oz�Ƌt�c�!���Pk6`�^>���țzgie�i%�aU`#R�,���5Hz��'����s�آ��\Y���ԡE�}�~��� �,�W������3�����K��iN�)_���>6��S�>��ڎ-|2���O��>
��i'ǂ��=�^�c���Q�Jp�ԥ�h����[�e,�/��`��ȀjT�
LHXЮ�f��1e�?-	�L|Y_�u��.p�F\�h���h\9H�K�"�`�X]�fٔ��I�K�h��z�I��^q�G�T�Z3D���M]E�4�>KP�Oգ�MW��Z���fb�㝏�][`��ZIt���w�{�v%IM���V�d�1NX�C�;��l����}nk���'�ѭ�Μ1i?,�4�$c<銱W�od+=��^J`�EN���=޿cŐRt�!Bn`�B,k����ќ3D��#�}�7���s�Ϟǩ�K'�Ou�c1娼�����mׄ�l�i�㛞���^L��b�����=��_m����ˮfH���U��f�We#�%�=�`�8C�8��ub�k���v�S؜�]�O�z"N�gݡov�p�3��zt׳i��(�l���g$����4�Q��1\���]1��-!mu=��΍m_��F��ڄ*���*�_?y�R�̈́\G16�b��OW7Ov.Ur;4C��Ec�Yp>u��+N����ؘ�6Elʾ�5�����癕���c\�EoK8�<�[��0����>u�m�eg�J�1�<"���nd^A��{6�[nM�OgW���Eb�q렋,O*e�nD��f��p�q�
���+w=��K�,D��D��R��Wڊ�E_Nj�PˈdB�����F��]p��G� &���|VUI2A�5H.��k͑��s�u��6��SR�dr�W�'x�ʺ�z���/5�o�Zc�T���k �ANr�Mun�	pɸJ���9��j;v������t���X����;WVxJU�D�^�� �-u�i���؏�H߂�(�<r,E��T��L|D������v¯[z�hr�t۝�F�����P�B��2�1zh��tyh�G\|:j��%��ǐL���$�N1��G��F��^�`��D�~��Z�����*8�p��װ���I{���~���	��~�J�qe����ftȥ(����(�|*z2v��Q̧���M�ɮ��`�D[;,�$Gt2(�n.f��S�3����3�
�Y�|���g��t4X�K	��������'�,�iVߝ"]V�s`�Fp��IbF񞊕j�9�
��#՚��P��5����'q�w���&X�PH�ĉ�p�	�g8�Y��^��=q�6�w#���!�|��]%Rˡ8�ryߍ�C�լ,>���y��'ש��ݽvElu�U�R�A���k�Fl3bcH���a~�VsJw��[ήl�1�ޞf�P,nO��S��{C��r���ݷb�/8V�Z�'�l�t�����%��PC�!&��|r\����h+�Y�T����o,{K��;e�3#c+������d��|i%� G^ʅ^���^I|�sOM��}�))��w<�ŷ�$��6���S�o�x&�{ctڵW5�}���kV^w,_�����?|���kn�H���H^3�(�eEv��#�q�ӽ#7'2+�����iޝM9�������\t�5����^R4�@�y)��5W|Q�us�8}���O�y�,*��3T��lEd)sGGtbxչ$u��a�s�t�3�����n��-�O��o�s�C"���oH��lp��(ۙF��g����v�#�V���ԣ�fqH,��q�t#֢wbTgL�E8�^t+�%lX1Ѝ)�(K�P�DM:i;8��sی*5���q����ʢVlѢ;�f9{�xƷ���p ��1q�&&�j�f�=�k��c-Ÿf\^�ˑ{c��EbT�Tg���"�b}��(ױ	$a�KCݕ���*ao���rɱ�w�9����y�b\�%D����j�28
t�Y8h��V�����*B(i��԰���DGF�c#ǅ��%p~)yT'~X�+҇��2G��$�=Yۘ�=�&���S���Ki�
��-Q�Վ��l쪴��7��#�,�OZ��%7i%�x���ÉV��+-d��CM��ͼ�Y�i���blR3��_v�xS�.�m־"-�5��#�
$����_��VmE�<�R��n�5�C�@k�.<�;�R�H�j�����qQ�xҔ��.ҵvN���k彶�[�#F�@�sM@���OR^㴧]%���ʊx�E�e�q��v���kjuv��6����Y��^Q,�)�9&�1�kM�j&+��=y:)��^�OB�N����c*�b��u�Y�����vӸ�`�K��@��o�_["��z<*�p��ǝZ�~LW������������!ھc�\����ٳ��`�]yG�ݻu}˟_g�v�D�����鯎��b�f�@ײ4�UP���N�z���Q|�D�3�n e�̥t}RS��������N���Jy�� 2��<Lظy�y&�G�~�k�{���LS��n�u׎�y|쑈�z�T�Z�q
��."�^�kA�r3��[���:��K�*�e�r�q�[���c�m���X��t��82�x�`4�m��8��J��辈��b�P��<]��E��]{0��!�huQBR,�cA�t��p�^w�6�C���e/>'���n/��Y�������/<�����n��O�����j2���6�+9Rzo��VD�$���۸��$�^q�k��mp,�β�n�UvN�6�fNF!��6�h����"2�@p�ö��m��7'PݳM1Ǹ
=�ռםy8J��D�Ε����u�eZk�����(����R�%8�ڗ�6�vi�[8޳��i!�����%�RTmd��CB�i�"�ٵ�a6�L�����v�) xv������N�u�L��.��O���*�Q�8٭�!�4�m`�T�Y�k�R��Ө�+�V�BJs]evEy�	ҙ��3^|P j$+th�����ϥu���Z)����!b������t岜]+gV���_*vV�&E��:c;\�>�B��7rV���d���L���@�r��ֻm0����j��+d����W�b8��������	�-_q����i��m���}-諎��V�$����"o�����U{�닖���;�m�>���J��W�.j��G��w�E=��/�B�U&�J�z!�W�T�iL��3�2��Tb	�q�}W&F鮬�هfYQk�3��k�B�'Y�jm9Em�+����[��u2�L�V� ���s��%��vA�����9���8�nP�X,9�Z�)w�����(�5��_�猏y��<׀����O��y�V=���Go`<�}t.E�'b�@�Y��Y�Vegj	hs;��c{Z��«�V���(�̗�O�eV)y۶
�e%�)�_@^��_)��SL��1:���v����f�����8:)�X����ҧ�9�����|M���Ggl�!3ʳ�CJ��a���嚹���u�14HBE�V�u�7��t]J`��n�-���_S�tc��g�,[��o5���w���N�j���|W�!�i ��T�6��_[�r��EwS;�)����٬
�D�jIf�7����Q�}i�J��@`劝�+���e^�Juo�Vp��Ҭ��hNK^�R�r�tn�<�&�=}���Ϥ��$�.7�VV���ĲW}X�\���X�bw݃O7��F��kYOq`9��6��m�����t�������vi����j�iot��Иv.�/)�v�%��v�$#�jӑ!��'	�[̦&;�5�� ��)��ȫ�>�ʺr�T�d�z���T�����c�X�T;Z��Xt����b�r_+�qJ�e�D9�u����;����"fk-�*��ke��q�Ʋ�:�3 u	nG-���y�/������b�q]	,���vvRu9���_o-�0�$U�J��F2�R��	@�J��{�4���d=�w�"pAimjě.���l�=����ۀm���qI>\q_E�3�a���b�lУd����,�n9��.�F��������1oko3۶��S�P8�9�r'V厲U�S��Ʋ^Nx��Sf��ԂZ$�ӥͼ�V�R��w�22�r�KT�\������{*P��q5��2�}��w��Z���0W-[��F��QY-[m��F�(Q�����nY+Y+
ъ1�Z��X6��F�R,�J�q)�(VDeJ�fcaQ][�ue��[K�Z��T���s*TR��V6�UkJ�f$�jZ�����Xֲ�Tɕ�`�4�b�m++���SD5�r鸢��TB�UJ��lG��W1˙kT)E��j��B�iV�e��m��us㋔�L�Am[U
ղ���*kU	jҖ6�X�%�m+��[mF)m*
[b2���J#r�m��s+�ժ�Z��X#�Q�ƪb��LJ�����P��]4�5�T�Ʌ���S����1n"��k+Jۅ�aE�Ub[m��+j6�ZQ�e1b\ɂF�Bڵ�c�(ְF2�VV��F#*X����`�X����L®Yb�X6�DLK��3**�(~���~�T	��]���i-�мG{rj!;^��w9�g*��;~y/{�7p�����9�VV��g\��.�W�=�xF8�I�wז��z�&�C�C5.���]W�{J�ծ�܊��s��m�N%Mht��|�)�f^�7�6#�G B"N�F��2�T�F��6�p6�m�� ث�<�q�=&�s��K�ЪZ���w�/~������f?-"���b����������P��3�`���<����� ץK1^N�XhGD2�t�н�J�Aڥ}��I5Y�}�(�tˆt��SX*Y�l8g ���������f*�KN*��α�,�(˛ٞ}�_&��
un:�6">��A���N�#<�p�S�ȟYP}h؜1j��裚��3kx��	[�/dÀ���F�O��U��xJ�l�����RQf�0���7��r	(���'�7 �+b�z҂�m���6���C��v:�R����W�\�]�w?b���&�-X�}����3���N��u�&;�,�`l�d�>tsjէ��������:���Ʈ��/cN�K/`FS�pp��ɉ�7Z%��"����P
6�+����v�s��G�0�\F?�b�IL��fS'�IavXfY�(��-�Iv]*���*E��Vo�����B�B��I��W9q�x�an9]������MZ��Y\v��zBZ�Z2�0� �v�=�_+]ֳ�����7�̜uѭ����>[(����E��z��dq�λ���Ú��@�'j�7鎨��-���ի+[�
�ΗZ��n��p�/�Ҿ8���[�,�����<&�zd�/����6{�A���h��1R��1J8��E�{|���쉡�_�Y&g[�9��½��C�	�j��~�� �8�2t��*�V�!ӞP��3�kJ��b�:M�ʩ�\�"-�EC8u#aДxC�9f��*b�u=pȯ_!':�`=�3���7Eߚ�+F_Hw!�M�HY�P%F���B�n�����5A\v�չ��*{=�'hg���ŗB:�]U��Z�nD21�C�Tt���q!OhMN���7���<�X�f���0�9`��x���Д�i�a۶b�!υ*8`=�ȴ�[�ڳ7gw���!�/�s�~�xcf�	#-؈���3bV`�f(
v�v�R�e.��j�,�a`�gK�ZM�k�Qs��Y������7��ü���c�C�@�(B�C�S��]�������>��
�b���Un.z��ƞҥ�y�؇��U���Ӕ�L�Ʈ��T��y�d���g�їҞ�:�[�Z��֚z�wga]�q��7��UҰ�yL�}�-ts'2-�qJ�JCmX��i��9
u����W,M��"�:�ˠ�Z%Z��	j��׋���)�͸s0u��(�!V���Wa���\O�s��ex�Ub���+��9���L��n�˵+i�WX.����u�����g��!y�Y�nm��IAԈ�On[N�5:�:�AGC�I.GmQ^i��kkv��1!��A@9��#ڡ�k�9\�=9e���糓Y:6�h�,d"�J/|���X��4���r⭪F5�&�޼��.4�����9�}��3G��]3�qC�e�w�ߔ�q��#�ݦƪ��߃��u�"�OKM�oՖ��_�`nm:���������-(�V�G"�:.l�]�v�˦/)�5��^lC��R�g�SR���=GFU�$ud�c
qn8����L
�/1��������\�U��S��2��:+]=�*��R���ў/���{1ǫ/E���n�ruG.�ItR-�܉㵩i/ګ�z*[A|Oa�O�pÁ�*e�é ��؝ԓ��Ί��b��
^�Y��`)���;�G��V���ϸ\m��.^���t�;Q1���H7�tw;�uΐ��<G��t��Z��=���Y�B���ͭ^�����xػ��H@�שM�`S�Ǫ�����';�����3<o�{�j�KG�'�||.�ޖ��\ΖN�f��2�Y��: ��Oa���5M�l��U��O��b!�aHgo�m�9�r�q�SN%U��N��}��{e�B]L����A2�֪"��ڂ��t��.Ñ�=,�Fʾ���ͽ�X��m Z�Q�"Գ�����R�E%�Qb�R�����\�:��b��Z�f��{f#��U(>�D@��/�u7�R�}t���w����g��j@Yq'/�%�q��|VC�P�v�P*B�d���ɎnH;aW��p#e�ݢ./g��ݼ��S�9n0��A+ �qD'���D�B*m;�ߢ	g���n��U��wJ~���X�nL�F�f� ldc�.� wu��:��88GM�隊A��4$�n�, Ӭ��ykq�зL鼻b���iL�]�p��/hS�'yeE�s�N�.qC	uq�R0�״�-b�=m�a��Z����U���C)�����6��3�^:ɺOWM~�5��u{ �ż��QZQ��~
�����oh�S{=���,��M��`��u�ן.U�%���~�ʎ���y��'˭{Y�]��a��h86M��k�u琠s���Y�O@&j�Lw+BiGaԻk7����T��Ț7�����/^��U��NU�?(yfx�=L:�'�R��[C�C�sۼ�ګSZTC Qt:닾��^�(���t6Fl�P!LX51�y��Rk���n܊����q��3F�qM�Z,��Ɇ�`�mu��۷(T��(����|�(���0YT�
z!ӎ,m:gV�D�y�j7�Uq��)5���JzG#C����GH(�P8�:t�^�eW��4��*z�oT����;���}�G�k�7jl��r۽�*�^/��6���b:"D���!'t#CjYwS����|;��U���)�{�1^���I�+�\H�T:!2!��1=@K�*�~Z$�k��z��d��X:�[׽z��VCӦ#U#�è�eC"�\� Uu���>�#e�-��ŋ�p���;3{w��!�<n�υT3�'���V:3��6I�	R�(	��^���+���s�b������5��~�����"�\�qya�u$B,j����ᘧA�^������˨�d��u�p�,���~�����%I���ffM"� �����k�SQ�TMz�.���1��u��"c]�#��N�Z�]���K�N#������H �u�i^�v�����N�Cn�\�٠<���]�#!MUr�{�^[oaӹ��(��j��G\f��b�Ӏ�d3�͝�@�q��T�������ۧTV�;�%����E�զ!Rr������H鱔靸`�Ő�@��;��h�s�\>����A���t�]�4�:͋g�	>�B���Ui�Q��N	���e���2�Wv>}pt��S����{ў}<{*Q{3�
�9E(�De7\m������.y55�Zܔz#zp��C_S=��dq�:��V��!�Y��!���}������a^���-<��6���\ �u����O��WI��s�w�����YZ��B���{����g���A�fNW��H�@�`ub�^�(��:�N�[8�lN8�;�����>�ӷ��a�9��������8��v�
�]����,b�	�Z�������q8`\�
9�	Sk*>��|�\X2�5j���*�S�u�v�NުZ�!�Tnl��}�򡐦(tˈ��}�WP��D\)fq��&'���B�u�x�kE%�'Vms��n�7�q����n�ay��#���Cc���ڵ´Qn�26o<h2^�v�{hkd45�u��ͽB���`)�֓���|x�	�I���X�*���+�,�P�;mX����9�A�Ѷ� �2ȫ�Bs��v_u��;�rW������S�uu��u��Ľ��2V���s�]�9�������0(J�ȃbh�\�_�}��U�nQ�s��l]���M8��Q�e��#E*F+�̐�j��^�(O{u����a�����|)�~�$��t2*;������4S�33��yT�$U���=\���A�����,'_�p�Z��J�O�Y��*$��}N���>�c��i�k��V�C���V-UK�?	Gi1]+�Y���w��ɧI2�Z���Ύ�e�*ݞ�Am�!�Bh-V��(݉��ј2V�j
���U,���S�x�t��WR�>�����]B�E"��ڢ&�9������N ����jNy@9���im�̧b�fpخo�,�����Jدf���eŅX]yu;��=��M��_lR�1}��L�:
5uk�wc��xﱟ3����*7�)���/6�.����ʰ�v�b�;�Yx�O-av����i��.N�[X��Z ��Jf(�R�⍎�w��-Nٰ�j1�#U{Z��J�<�2p����H�K�d%�1�yu���M+�޴�6��y]�0W-[�S�^gӧD#DX���ꉖ�>��u�oe�u����VF�p+m�W�����λ��8~��iᮉ[�P�7&m�?fK���:���.R1�jH�8'��s�S�t�+̓G���e��0Co]=�)y1u)-�|"��z{s��o����V�QE�O\=RK/zBa��ĨΙ�!ם
�hD-�:+�I���-ĉ����d/2fp�P�����s+9���m�;�G���%�wʹ���ꙮ���=y=�r��ۘ�0J�3ŉ�ʋ��W���um�C��m��o>�.���B&n���AH�Q�1B!vPF���UzYW�M89u��i�v�e1���s�qt��f�hJ��R Fk�2ϗ4,1_��ΰ�]j��*��A�ኽ��U�v�m_�fh��
���ש�	����EX\u�^Dk�¸�d~���S}����A��j Ԙ�n�"���4!	���=i��oe�zd��\��^~�i�l�N/DIb�I.GH`�D�H�4f�/܉+݁׸�xU�=�w��!�,��<�NN����)�7�m[��E�AC�p�j�k�U<�%��#+��% ���#	���&_t�]u���Ek@}�ý���`�ǯ�a�u-�
��i-֝�q�̊%k���Y�fCy�t�ɫ�������T=����Z򛟼+de[�jD7�K�J�wu��.�����T	�=nNaV���s ��膭��/oҽ���a�ײ���Pdf̠lۆ/�UEZ�z[�j�����,�`���{�gm�:le1B���:��v9»��6�*vP.ڻ��Lb��SE��W�7�`�>�n���.�,�T�N�����l�H�(�1%�Y��nŭ���s���cz�ط��uJ����>��G�+J:��Kޒ����w�מ������pSsi_�K��j>��*R�9��f.�Hޑ#��,�3����1\��Gu	{À�^�|���lr��]h��z�a��0P(�܄�^3:c�g��wthq�C�;��:�S���N8�rά�K�E=���������*�QS&��<M`#��t��&���耋����O^Ψg�'�Yq����qؙ���l)�l���QL��~�q���@�D���F�2�T�F���Ss��a�3ǋ`�u�:��Yz��z�VGrC�̈�޾Dj��x�?{�dh��s��F������j�Ћe���x]RӺλ��e��^�*��:0ʍ���ө�23\u�o&���@���eOw������i*�c:��G��>�2R<��|�}�K��R�O���-|psO�i�ŷ�'���p�F�90�)�'U�~p�`��� ץK%��']+�OI�������Ώ��w�w����FX��;�fw�Θ�OS_�R��d�P�L�4ȝ�0�G�I�bpǔ�Y�<��f�Y�֣��X�j�8`��G'Yы3�'���������be�C�oT65�z��9>k�O�x�D��>�l�MTO�X�)�']�r�j����Vnʈc�+�wu�C�x.B;����v��Κb,law1r$.�+le���g�G���[��m.}�	W�+Z=,:
� ���N��8w*P6mԴ���K{�)ޫW����4Ytj�Mt�9��%Ÿ���P[�D^|���U��!�J&u�{����o��}COٲ˅Udw>�y��\iz�v���v��^�J��{��L�o��"5�~,�J�<lj������v�V	���h����K�q�h6E��F���Y�*u>4%�L;��k��J��
���V����3\��9 �w��w�ֳ�h__n\Zrj��2�aM�r����ڣ3Q��
� �l��KoJ��9C��kvjz.�wJ��٘*�#��OjF������e`�
�h`�swu�	f�r���ܒ<)8��R*]���gN�n��6)5��bI�.��غ������ݙ�A���N�u���H������u��H���N���:�<�o!I��`��ͨ��">����y�ó0(r)�kF���-Ecz&3t#Clp���S��Fb���gR/�U�ԭ7�uϻ�Fc$�\��\B�����h���h,�f��5>[2ͪ�z�&�Y�P�ޫ����7��c0�앚-Ku�}B0�5vEs6�Z�u.r.wM�,�y<����TzPO��D����C��A!��;{���3z���<C�{�4worq���5��sz�ua%��[��D��'Wn�����j���+�����}��1� 
�܃��e�Hg`<Z;J7��d�ӝ.��<�0����̨���/l���բ2��]}iAH Zb2�7�}���(���u�vU�7�v�nA��+�k>4�
�#2��0X	�<��8�jvs�}��ӫ����')��`�0.Ӧ�@
L�s���m��IyYϪ�rZC�4a��YS�W�5�B�j����y`uf�< �ɼE��g��r�f�szK
U��3R�h�|4�*�Y�Em ��S��i�i��u��":�N���ҞOx2�X�`���(ΟfR	X�͡2nZF�,`�GH�$�8 U��CG�@�H������HF<��k4Y��n�7��&�h����m���P]1v�I9B��@�wB:�1��(߀a�K�=F�!�٩[5&�с
wdD�$����u!#V�vDނ��biD@h��!��4�͊T���R���{�n��䀸�7Z�Rh�X#��lI@�Z���	veƕ���0�Dn��˫xh��_ea
���#O"7A�Ę�KY+�R����[y.�D.Po �y7A `��� �A�R�V�3U`��̺ �]Fh������ò
�4b������J���mea{q��9JT����┲�<�;u�u�Z{.w\k�'GGL�V7�zK���9��k ��8�`!;��6m�+A���hٜ����7���o��*�rFW*ᥪ]��T���T.�_5��:Zɲ�v��>,^�I��Q���$��U,�WVr�.���1Z�e���̲ο��m�T��vQ�ǯb�%Å9՛I��;��A�_S�����PLWl�}wF\o���w!Z�-�a��Qч��e[3��A��u�-��+[�dӻX��=�\lB� Q$
>P��$mm�j[elU̗V��meK�r�n6�TE����)S�	U��P�-��Q�1T��DV��ь��ڔJ���3(8X�PUq���Bڵ�Z�������-V��+U��e(�T̰13p�Vj���RYp�"�3�.%�UX6�)��e�e��QƊ��`�!S0s,Q�E)m�8Z��ELK����������mUT��m2�j%iQm��jV��[V�*�c�R�Ѫ�*Q+QT�*V,��-�6Z2��DZ6����*ZQ�Z�h�,���*,(J1�URَ*�օ�ح[ch�jTF��lZ��iX�)R�*V�YR�F�Kj�h�ֵ��-�UF��iQ[U1�$�Z4F�E��:�����u�]�Qf�[�do[��.��}��
M�����t��8:ഫ�B�����2��'JԷ:���a��4_#oEM��;kq�Q�ׇ)oH��Wr�o�� D-��q��7��B��<T�h�OԫC�k_ԯ�8𞎇kʹ[6v58gU�0f(�w���wO���TK�����aP�z��)-u�HV��C����5Tا�0!���P�]��CR�q��Y�K�%��k��K�?���0��W%����8����{�<o5J��"J=��I1�X�*1����ˈ��
m
�J�n!P�������w}ַb��kY�Ӱ���]	��g�_s�]�9����Ȝ~��Z��=dl��L��ٻ��:�)vHá�����L��+ᒟ<�$���74p�'ZdX�H�g�.�Q��_d����F0���S��@T#�6Q-��o�`�2:M�9��Cq\��R�u����U�R��τ �薓h��n�.]y�0%9�i���B¸+��m��r$!�w�kg�	E�0��8#��
����J0g՗\o�&�=ȶ,�ѕe1�3^s[Lu�'pE�C��&��؋jc
%׸"+��A^�J���lA���gx�H^��f**݀y�\j�RĢ�Jd'���M�\�n�:���b�eb�o�k�B�c�t�EP�Օ��(�-䃌
��qwVs�y�R�d+��Rs�p�����>�ޕ�޻�œ�1�:�N�mie�e��)K�Co���TlD��Rh ��+�]I"r��R���u�y�$!�P��h͚,ܔ\Z�-t��y"��[[�MN��q�gy׸;�����m�E�c����\<+_���(�f�*-vf��8�A�V����VE�q��h��_����o�q��=5��4���l�GM�f+��p���L��y�Z������]�e�����E�����ݜ�69	���GGt[���<��uk�e�<�.������c�
��J~oV�T,���)F�P�؇l`��[�F�B��r���>qДF�����<��_B/�N�J�3��"B�cy��dD \od�{����/ܪ��sl��k���]gs�S��/�{�G�i����p�6�VH�}�����>N��ϕ
��pM�s[�)j�>�ZwƯhr��������n�ȑK�,���.Dp��x�C�L�`=��h�D�;����\&�|6���ʴ3���-��$g �vva'<aV�Q@�Ok�m�*>����o��k1ѾJ��!{β,�E�Hh�!I�!����5l��vvĬ�J��܀l��d(mEqB���Y�a�8AmwdE�j����I�y	���ՀΥ��o=�{���MD>���U_*� ʆcC�0˝K	k�(WF�Ǆ�pvUb�۷�W�9�Sғ�]E� �u6��a){.�3��T͔�;��"eOLP8Q�B�<�]8�5Y�\:�6I��s�*S�"�j ԘjB��ܛE�;<sc����{n������5E���4�ƈ��t���0c�M{�h^�A^��z���V�^���g�B�p�#��>Un�����}�t,!�u�[�б(w���Tׁ�y{(=�����9x�C՚1���,������۴�#��vҸ���|.Mw���~�M�o=�g|(ټ�	��$z����G���U�S��^*@�F��Tӷ�I��iW/%M��bġ�Sq��9��I�檯m;��Y�<�oV�4-	�BܰC�n*���ׯ�΢J�O3*ju�}�ٱ����j�wyϩD��]4Z/:�N��73v���M�7�s<4��j�F������^)G�ɇC�n��C	΄����S�u�շغ'�6��T��"��&��6x�R U�yR����n�������P㿘�B�}u�G���V=����8����^�(�`�
A��q��pxւutEo7Z�F^;�ת���l�5��U�S�����1ޞ���ϟt���R ����P�b��P��c�q~�(ٿn�E�J>��v�����:���3v��5mL�㘮�zq�$N&��EM9��*�!�^�gVxs�D�޼P3���{����fq��b�Q�,O, 2w����I�l��:�:�U�ՙ�^�]Z����Z��-c����4й���u�S0k_��1=B\�ȿDQ=�چ[Kq�u�;/�c��LL�n/��
�ؓt��H��TE�/~���^Z�O�D�Nͅ�i���֍aڊ��ʮ�X�e�P	Ɍ0�j�q�5�,Ru@4��J�TBTC!�.��:k�� �2�s���NY��L׆Aإ3��=L`�g��&��f3+�(�����T�U)#hs��������^O��O���X���}w=�7��';������$��"�#��DR�-����;�k�PsN-���T!c��T��z�۾����� ����K@l��֟�Ћ!Ő�'+Kɛ9]����t͍ɦ!=7�g�x�6����@n�U��)���}]HvfjW���K���M�����[Zpdh!vé�������[�.��D��Ɋ�l���u	�.9OOPMI��'}k_w;ۣO(����n��w;fnr�V(&N\��(��]r�ޮԩ�E�`�V-Ub[���"-���^���ߞ��
��S��r{75�+A������j�7��>�Mt�9��L��0-o�h�t�P�mgk��4z�bq���T��`bu�򧁬�E�oC.U��ei�{��64�o��D����b������~�VА׾Q�����������>&i�~����Uio�W����4���H��_riK�Ҟ�KS�2��J�	Bfh�J"�J8��E�۹�8�T�u:�k�-]�^aaL�����ff�{΄�%�6 �IzW
�s1g�� ^�eHK�C���=]B��w�
eL���,���s�"̢�Z�Ds����f͋�Y�;ݼ��X�wB.�I*ֻʌp@F�L����P�D)���<Rr����Vw�&��b���Ŋ�u���D��;5v�����l�=�F]J�莨�n���7�=���װ=}L'b�ip��in(�2��X�ͬ�ע�m�`���ǹ�m��,>ϔ���V�BwQ�ok�2צ�v}�3��R��]Mf���J�Wn��S�sqe�iU�ۙc�H6�]ќ�L
���I�ս-3�����ޙ�5�̙B����t��.�L���5@��K�x�&=�ᭋ�DVh=�!*�T#�1}�x���穠�����s��]�i��|1�&��dYnEƈ�n�ʂ���v�^��v�.խ���Vog�s���'I���]��ד�B5�{^V&���T���{q���PԜ��n{U	�aK��	u���b�Q���\ Ȭ��XA�Y��-��eo{�M1�d@��	�ʞ��۩蘅q
����x��ER\6:\+K^&.�9Y]s���&��XPK�-�"R�����jq����x��k�F7��t�{��=�׎�Vu��ˆe#��Vl�@��.9u�w��2��t�[Z�﷗�}�`Φ����w���mƿ4ϳ��*2�j(\2:�� Ep���(�UV^���THR*�ި�!)=�{wv<����U�bJ���8�lH�^r�S1��I�"y�tru�MZ���DQ���m�:
+b�x�j��82�}Ja��1u)-��h� W7G/��Pb���ګ[*"Ν�#������ᐈ��:�'�!ě&x�~tb�%n͛VJݝ)�P��{x�ԑ��/`���l`�eM~���S�P� ��n�*���;Lo��`�muBn�SS!%��}��B� �T�F�;�҄h����V��9o;�X�oSn����|���"��y���|��˧	*u�՛�6ջZ�Nϱ���q�}*���>�N\OF�!�Hp8�^T)���z�z����`*T�Vꑇ���Q�+ا����c�,]���ZV���Bו�seԩ>����
v�X�j/�Q�<�����^�K<����T�~ϻُ�dU��9^>wyU���u:Q��I�Hp���x���/�l����ꔽ�/�7�w�!ڻN��yN����W{QI�)�0��iȍ�A�ٌ�(��B2v�a�q}�R��uf굴�_�P芖��6U�@5/bE�R�`�X�fЋ�w3��J��^E�rF��~��{�{b14+�ᰀx�r�N�:�4�v�v�$���c�<�w�Y��ꎮ�7�DS�Q��4��D�+�$�!��r�d�ad䘠Dק�����77xr������h��ʭ�T���5���Cդ���X��p�|�������e�ODFՄ�T�ݗMGh;
o#q���UEf� pۆ:���>r�Լ֐FT
"�G`�/n��.�U�,t��{����G�!ë[%o�j}F1���Rq�,����kHނ)9�]�Z���x��Hɳxa�'A��g'!���Pսr����C�fs+�`�SM��hr��|7;o{z����X�v���>��	�X�ۜ�M���8@YϽ��C��dTƙ�tΛ�S(f�@���g']�=MwR݋U4V�j�R���[��^�wU�X*�{i�Złz�9Դg$_'s��wд쬡�׀�f/�\��W<YU��z�wT�ް�=�e`z�3|�u2l�ln��s���'8Nz#��e�P�"��u� 'i�~.{��N.c�����:�U%���ZY�ʖ�X�E��1`ИN-㾷*!qn;\�f��.î�Y�9�ه�o��MeX@�+�+[��Za������r,�TӚuJ�!i�c�w���ӛ�u�>s:f�w--f�^%�Ta������z��G� �N�tu����[���:R���٥�L���}�7x+OÖ&ӡsNz�yf~�hc����D�ҍ7U6�T꧴���#�:8?�3Ɲ��HOO5
�D&D2�q.x�A�Y6�u��8���Q�q�Ȧg
"�$�8b5R������]s	����_=V��7�/R�hb�z�8��y8�]��ЋR����n�0ŗ�	��LKu���յ|��+���;c������1�v�U�n�_�θ*|/�^H�1+�b�"�2�sK��Ep��(As��{2S��N�y��M5p�x���5���.3pr)E�3U�OJW��p��2��a:�ܾ���/ }�Uc�
3z�Ӊ�U���<)��O��O�:�
9';n ��ŭ��;��u��)�G���֖�(��z_�]�W�[��}����;E?C&6es9B͋�({��d��[�{a.�HuY���6s�Q�r吪�V�k��Z��s;�H�@�8>�e��ub�k��
��f��n�i�^�����5V���'��ܶ[�z�d�ǵ�Pt��U�< ��.��Ucs���x�ʩ�����Ʌ����q��o��dĊ]\ra������oK.-���}L�y�,�8��tU��҈�mNRN��;'N7�UC��1�X#i���T����g]J-��evF+���u|�Ϋ���Zm�n���CO�J$`��k�5�ˉ�xO,׶�,D�o>��!��M\�lM��Z2�K�xBP49�#��"B�Ы����n�z�5��W�-�.?#�OC;k��=�	vr�,��=�ӆ��ɕnes:��Q�����.(�a�����L�WL��l�;�>�O/:�v���}׫��\\�ڰ���Z����sO.�7c�왍9+���,HK|W˥����s�;���s��Pw����D=;Cf+��+f@�<z"�#p�ړы��5��ͫ��,�eUJ�v 3�cU6��Tc��7�."���{�MDejp���S�g�m��؏�9f��,���
��\i�JPd;���/�����^6qs��<�Z�Mt�7��+}]լ
0��vK���)���e>v=)k�0{ŋ��y��味a�
�m���Ҍ���F*�Z���Sѓ%tP�Du��ΒD`�d;˚m$��s}5Ѥ�͂;A�s�'�G�����ZM�k����409���d���v^>�cl�;����(;)�ً3�E�0��93n��d-��!R.�+`�<��@:s-;&�t�,E($@��	�ʞ����D�������x{ű$X�{*�5�L�؊��0ۊQY�E�8Yu;Y�E9]��Ov<ƽĂU�Ɇ�*����n�L��	{`�6�0[�6h�orQq~U���QZ�æ|�dH��Ƈ8B��]Gf����.�UF�b��z��������$hs��c�N�O�������'[5!i�wO�
8�a{G�m�z��陷)�Ժ!�1xm��
��_}	7�u-\M�}sq���ʲ�����N�*^@5oJ��s��fPv����b�����ͻ
�G,�>���(�#�F�n�.s��L�g1�3ͱ�M�K%�ɩt��=Gf��ֳl&p�p�-�%dy)-�A�E���8��T��u�&��̀�f�Zy�'76=��˹��y'wy5��$)o;TGtu�ā �$F����[�愀��(p�6C&C���Qřonԇx9�۰20e��.���k�e83s������`���Ԥ�X��BQ���|�5�+�����ɕ:AW��&>�8w$�	#;:��Y·�t�k�"Ni������j�o�,yV����6�aYA�fnsB]!�Rn�̀:Y�x+aG{�Z�O����L(K}�$�K_k���'�x�T)\|n*ݴ�o *��u���s�L7O{[.k�{5�c,��E)rd;���0-���o��,�}au[Nʱжym�ǎZ�;]���1՘*J�4h�/W�V����93�<��^�i��;k��Z�o"�[�m]
�UL��
\c*uY0i�Y��؝��ls|���B���6�c�V�lԧ	�z겆���e�	�����v����b4���/�l%�\%�HϞ+�V{uw�D#��(�N��[�-���$�R������A�R�O�u@J5uͥ4s*���S�,��ɵ�AJ��FmlvE�������/��z��e`����[ Z�'.��0N�
�m!�kAVP���u���.����HT��P��2�m�ާ
l�5�i�h��)��3A9�̸wZ5(eD�I#+LF�^V��
Iu�D������o���H��!*�xE��n�����勬����ɻ#�M�t�h��2�$��ҵ��t4,�5b��R��q�� 2ӍY����Dl�q-�A�x�g�Bt����h�	� �A���Mf��K�Uzp �4[(Ve��^1���(�d���O�Zt����˸eʹ�ʙm����0��R�/6�e���r]c�_i�=���:�uz.������f����_2��\����Sx�\�?=ʱ�d��c�����:��(A�H���e�v�V��:�\(�ϖE��!�u跴{M_�{�*K�U}˯7fQ�/��X���۸�������-cgH�Vi4ݩ��^����̐gBΤ�Oj�DUH�C8@⮎�"��S�Ĝ(fd�d0<4!/��mR2P�,�(�+�跋�ƤZ;u �La㥽���cUJꗅGn5ˉ�\=�+6\u;n�\c���u6����_m����q%`AA�kw�*�E-�m����*1�"��b�UR�Dh�aR��E*\J�3�Qm#j���jR��Z��B��T�l��D�TKQ,F�RVV
4��b�ZER���*T�jZYZ5�)mj,eUm�*�̸R�իmm�⠘ZB��`�������Z
5m�%�Z�Ұ��7,�-���[e�
�2��%�[im�Eem���PF#Z��(�F��e�-��
���m-l*QEѱDJт����)+��c[j6ҩiF���Ъ2(�*�W2���J��Z4Q2�["������bU�W3&3�ƴXŶZ�#jW2fJ�DE�mYn7,DX"�ԭ�(څ��X�T�����FR�h��q��imE*T��-�b����b,LJ(媡l(ѱFҨ��}wnϹ�{�g:U��ɉ��$6kz��u���%��Os�)��L:��C*S�#}P��f4;VdT�2k˯�]��21u�P�bȯ��q���'w��B��|+Y��
w���p�+��㾄t}Q�H�,����p�zX�u��.�y���b�Z��[X��ZC�+]U��>y��T��ο[�ݙ#��m%�w��\�8Et[�Cf���F���K2_�O�%��j߽[�e@��=���͖Qt�2��},B"]��6�=��4p;ٝ�hCv��u9o����6X�T�˗�l�(��*��Y{S'v%F{�z"�C=�M�*'�'�4���zV~�{��:�/)��ֈ*�.�v������;KG����h�G���=�72��m�ѭ�ސ�=���Q�yB�Hߧ��3��:,V{(��’���H�lR���Q��2.f$c�
4!$�(�%@�S^�����e�����q�suuA�7�q����;�Q��/��A�	]G	K���dx��$��M�����9�iu��钟:�]-\+�y�B{��$]*f12�@�C�3�i�N������.�F���F]ʻ��j�Q�;�N�R��T=B��[0\�c*�<�#rV;�,����"V�>�sJx�\����ytw��-҉tPs��54����wĻ��Hw+�$YؙcZa��/)fV�8_	D�n'-��X�o������v�$�l�؞^CHl��edM�˅���s�*S-T��q�.��ĵ�߃��!�mK�f��{}Z��%����E<s��A��oDIB�Is�)d�ы�AN��=��B�����������OK=��R��[����3��Á�T�-��X	D2��ٺ߻O�t&fP,6a���ɡ��qx&o"�����H��]78�&e���E��ԫ9�{B�%��o���ݛ�cC��9����病��J�n�$���`L�7R}YV����¨�[����69t�sWxԺfVj�{��n����^��a��{5�M%n�_�λ�Bxp�r�S����U��z�wT���s�ȫ�{��Mׯ�R8��1q�fޟVK�R���\EgH��O���@�Fn2`�'��oI�,ʔ9���\�aP�a��e�isԴ59�<<���bi⛮�Y㕡��˧�M����1�İ]��_���4�<�P
�)��ع�uE��rέ�E4A��guvlغS�P��Rܵ��E��"59�Nr�yt�z��-��	��nL�h��@Tշ8��x�����iB$�osQ�uuAn�-�3tZ��ݥ������'������gN��GGo�-O9�S��VHcu+ΊR�L�e�$p�}AQ�N�gQ��������{7Mm]�V�EB�(�xH�-*&S��V�q~g�>�p���0\swR�{�w+n/�v*VF��6��[�X�ؓb����nÈ~,�=�����0�	EQ�ǽފk9��ns�S�\Ьt5���u��:��wQb�� �,�鑒y*��E��V�\�9b�Ɛ��f�LdW����w �R�3U��`�*Y�gK���6��g'����,J�1AW
�]�B�Ӊq�V�O
�������y	��d��%&S�k�O4�m^_���%���
G���5�u��r5��~s�Zʠ��NM���j#�d��h�.NX�F�d��{X�4�������}P`�Y�9:_	�9]���Լ�1��.a^U��d1��qu���\-s�εbٟ{B"�m2�3ә�E�i^��J�����:�c*x͔X��,�]_j����N>�=�9��b���Kd�F���k�Z�j�ek��Su���oP�o��t�]�������c�<)T�о��\qr�;@`ݮ4':��^�*��|��0�VR��*R�X�vS|(I���8�U��ܡne�aQ����..�8�6�d��wZ�z%#��ot��쎑�>?Y8oWʔ�E�X�L���3^�)zo!.��`{H��tR�0`Ɍ��t��k�P�����TQ@��S�P�8oK8�<�\����&����9Ͳ(�v�|p>u��g��Q�D�wF#�������/�W����j��1e#ݽC�.yS7�3�{�ћk,�g$Ba�&x�2G\!E�|��q:p�����{���1�M���N��<��e���1@g�o΄�K�7�٘5�����A��C�F�1����?z�`��GT2W����b枏�
��y�w¦��
�t5�Q����@i�	�\%q�ɪ
�Il8'˔���_t����*;řs�12�����Cn������遳�Yp����棇�T�p��,t��\G�.��i�.���(]ƴȱ��L3$:��8�:b�g��1�S������m���fô�yx�e�~�����Ѓ�l"�O�s�5D��G����rg�'4����<p�j��u����!��ix2�x}�qc��©��cq�(Ꜧ��ڲ�J��{8�R��5u�);����Q�����QT������İꢲr]�6HɈ�鎲�2�GiМ�e�
�q��P�^�����>����'1�/E��Ą�3�b�3�a�j8Kµ��:��2eۜ�v�o���G���J��&a�J	��69S�DdL������!`q9���~���@����^�6���4P����/�I-v�)���d����1�=㐩|�s3t"�a}Z�AA�x�'��Y<��P�Xؒ�̈́\)�ߗS���/y`{�#�2*��%Ki]E�(���"�%\cZ�`�ǽyQ�Qe���@�0tf�*5����K�&�]���9VDɶ6Bq���z`���v\�|2}�bjv}t�ꭊj�;S������ך�����Q�C�����s�8��o]�Tn4�Y�&�<Y��5L���FFrM��ܺ
����6�O#S�qŔ]:Ō��)t��,�Dtu
ގ�ٱvu^̊����Ⱦ�a������0�D-"��T���.a�qH��K�3�QK4·Gdwa���da	�B��[8�No�^S���S���v��l,%�:�b��e
4tc\�bܗQ�����Bum���㤯r 2�j�d�ܴ������>K��K�W]�p��Q=)(���qx{�[�iP������`pS����1P`ͽ�9����ٔd���ܯ���a�l�Wܺ��K��{wU
bډf+Z��~�ph�f	�.��/��3��U>W�R� �9�4ےo���V�7	����iՙ�E�c�
8�0��b��� �j��Ѽ�����\�mEm�R�yu�w/*�ΧƦ�I���aV�?�@��԰�ƈp�f3�}}����Ė'�V�T�dEN�!��P�$J�`��*��w���jvN��9��ۺ�(��Q�(�=*�	E�T�,0�P8���1@5."m\nܒ�E�����$m�����L�͉p#+j�X6Y��$��E�=!��D�[����fؾ�o�����j������U�'�}������
�C��ƈ����_f0��|p��i�u�d�p�o�=���r�+-*�(�m$%����*}�jaFp����Y���x;vl�{�, ]y������ݲݗ��<���vh�@�$h5��3j�c�-����zl���CH�𫘡;:m�yQz"5���;C5$��C_j,�&���׏p�;\{�R��֮s�x$�h7ed��]���5��FT�ӟv)y��s�ˋn#׼J�bkA`�{��O1��ʴ���l����W�6��۳o�feBx�R_j��r���3Dk�s���uܙ�4��q�Ǫ�i`3˨h�d���r������
�y��X�=���z�<Z�w����`U��sihs����^%�z��]���-��)G�7�@�sWTwb�歩���>��n�U*��W��#�.z��QJ�F��p�2x[�/T����}�)Ħ���w5�p�S�{0��DH(;C��*��T�sC�UtB7�S�+�մ��|�]ޡ�y���-o^(p�L�R1Z����dB�$Ј�Duvn�57����]��m�Eub��Nʐ�/;$G��1t�n%婶`د||�,%���gDm��U� �I=��n;F���rZ�<'��<i�J�I�R�$]*
"���Bqk�wP6�j�9�sZ� UD9��9��`35�p��g*+ԧP����,PȀ&֥��_tr�_jtkj��ͳV{��<�x��:�'�]�>t�VV��[�YZ��J������8It�q.�Su�ZQ����Ӊ��W����[H�o�����K��mF�d���ʊp����}tf��e��R��*JJ^����orU�VW��̢���'mo�*%ã��O<��R|w�w�Tw�5��eB����9�H����������W�( o����P��fW��&ӏ�7�8�k�]�N���2o��Ք�m�D��\�:���rȤtz�L�,�U��5�?���/μ)�G��A�t�������O�W�+\�f�h��Qͬ(�b�H.$n�RYf�0��ʰ������f��������6�)�Rq�k[ʜ��Ƌ�u�n%�݌!��Egk����`O��x��Q�ҰZ|���+x��$y�׎�ي�����`��y��l�d�4\�ɡ�;]��ѧn�����׏3�.�M�˨E���
�U6��J�l��7��:�'^�; �d�+d+��	�i�Gf�,6��+!�i�bk F̆p	��%7�x����j�F�,e=Ŵ����Uy=�b_��/���S=j���~���1�H�$q	�&�2�i�Z���;S��9gI�a�]h���J��ŁoF8鰨J�F�Q�j���[�dafP����J+���!��\���dC#&0f��l:�!F�m<W�زwk'C2�6�Q�1G����v 2�:��D/�g��~5��	Z���0���&����z�t��#}3u�j5`g)���z ˺t6��B��:xs+��~�6��E�wg��-{���ॻ�-�~3öRA*���M�*�I��B����d9f�f�(�3=!\�ވG^��X�V/�3%:��F��.2��t�ma��DE��;�����&Q�J^j8|%a�2>x=��nئrF��^�ګ��W����o��
��szSZm2�s
_O~��٦�)EQ9�����(ht�3~�U��N0�PV�LR�0�y����2 �u�}�Yڛ{�˽��M�S�4���nD^���`6fp�P�Y�"Vf��"�p�|+m�̓�]�8��me���S��O-�0����2�WA"=���W�/W��Ș������Vm�Mve�	��s��e�����Xܚ(_�p�^��DM%OL��l�=el��C��竻���ƅ��
_d�W(��W1��.�.���w�� δ�e��Ý�n"��Ұh��p�^����� !_�e�l�Ez��uH@��E�maR-�ꖛt�b��9n�#�q|����k0���%{���R���'�֊� D���=j�ТެEo-߻į��XK��Y�YP�[Ā�.��̺�y�������Z�V��������3r���3��3'LR���]�xv]�\�w�{��*���;��+/��(�ڝ9S��h�"JG��&�����I�N81�}9a�ī��;�o����4:��8"�/�;9Tn4�J4OM_<�ւ��x�2�j�4'*����N��Ւь(�s�,��:Ō�	l��EAP��r�T���>08�\�:�Yb&�ʚ8.eZ�F(��(���U�͖Io���'v%A�.gF�ӣ���o(ɜ؆�����'�r�����8��q�<��aͬ�O<�tLfEu$��\�r��)e�nt1�Z=+J�s�5���ХG� 3�w��w��n�Js����dE�]�T��
׽y@-QL�F挊�1#x��$�%���t�M�W�V!�}�W5�K�u��1��+��������O���*�:�K	k��װ{$��;G��N�P����:U�㋱N��GC!�uV��6$_���g"�Bx�3�����_@=��L�!Ø�(͈ʋq8��Bb��
�`���ړ99Ů�{��:�3�����x�)��Ih��*)ۜe<�G���5����KTˮ��ē6(
uTv�X�[+��_o����H���UsyP�Y�Q���+^]S�p�M����]=��b`YΝ�{\�Ѽ-�N��S=kpZt��ݡ�	y�����\��Xp��*(MWee9���ar�,�����P����r��#��vSyS����DPw#5���:�ą@4����p��|tuN]�y��\�M2�H�þO�\V�����P�5�j�i�����y_��3.���5�k��xo; ��8�n�eU�1�gV���b��o=۔��<���]Y��yf�iC�ً�Vͺ��Y\���^���*E�;k�^,�)��Y2t+J�uH�a�z�!���np���2fbɐ�c�k~����nV]s��[�kF��H�;����������Z�n�f�����b���K;* -����i|�f���gq�:X��Nԧ`<v�r���a�*�+�����L6ѽT;7DySx��%��UN�j��q����_�±e�.W=S�A{�i�i�R�v<��
��C7Y�n�1�����U.淓5��A�tSc����Dsx}b ��b���k ���Y���meD���I�[����n��-w�M��T���
�ղ�..Zя 8��"Vw3�z�P�Of�a����X�/b���f��k!��(�꘯�2�8,
N�ýIJ��uK+:�]����y�����N�ݑ)؆l]��C����|# �u˴7��m.D�3�pۃ�������xq4;^'�ƾ/2_3�s����n��@�`4(M��VEjcA�l}�%��yS%�֝�Q.+�Iu	t�7�/���Ț����&ڼ��Ċ��+�u���uk���[A��JɡB+Ȉk���Z�Vzʬ&-ʆ����w�a�&�y���[�f�S��<��@1#q|rU!z�Zp�A�emL4��[�^�K,�S�t���t���ޕ��S@��j�2�Xx����n�H���y�֭���p�n��uu�*�Z�xA�W:S?��Ab��E�C*�8�l��eYo2�`�����	X>9�m��kaI�J#sn�����lPJ�0]�JĎ�����ג�G�ʴ���/[�	��sa��[�l��컧zSz^��U��+�����%�0��nO�L�ಋ���]&�y���YWEԨu݄N3d���y+s׍���v}��nuΕ[�V��#�V��L�����r^��g�`�;��:��珰vi�ַ&�D�P�sD�LN빏^V��R�n,;�l6��HD�� A�"� ��b�-B��������R�2����#m���DS�Ɩ��US)S��m��C-2�[cj����L"�j���F�j�AG�Lk\��s(���TEEDQB���\La��-�D��.Z��1��hQE���b�cEH�kU(�#�,E�Q*QQ��l*�
e1ŋ�4.\e2�+j
ƥp�3-�ET�[���\TAA�*6�EbDb�8��\����1*�[����DQ-�\QTb.Z�h���P�"8�L`�D\n2ێ��paQ�s(�ZbPƱ��ZVZ�kKn\�eQs3�dʈ������Uq��UV�����\q�`U�̖�2 �"
����P�1-q�#YE��7+h��**$mZ��)Z�RUF�LTX�!��(*[Q1��SJ��AZՈ(�i)'�	$��h�Q������
r�A�tqi�Q^�on���`<��Ӭ܏�3��Y�z����Մ;���|��X��媕��)ʤ/��>�3�a%$g`U��^/:Z���У�E������,Q&g{o���p�~����Fx>�1-e�3�����PX�d�n�*P�'�h��=�w1���K��/a�e�m;�6��~q���,ޕ�o�球�[�؞T������h��|,i�e�{U�p9��9�y媸����-蚘�ё�BQ}ٚ�d����9�Ui�n8�,͖I���#�uϞ-Edw���5"vE�dq��%��������g�#��6�0�h�]�e�_@��+�*�V�"�U���CX�]S�)���9�8�PK�I��q�u���N�:C���s�`sW��>�,�9f�2�U�ٌޢ���gm�;G6]#�F�L=s�*(�yU(R,RH�ձkw)2"zEҚ�o�y��nچ6��x�!<���ũ�bÒY�X:�R�5�*S��1�N9�k[ݬۋ�1N�g�z�ީgV{��&܊���'��`���Y�bxΓWi8;+�>Ǻ3�(qK u-�+��q>��n��Q�����O��WҞ�� 9[�B��ݸ{Z,OMʜTOZ�"������������?p��r����X��KѮ��I�v��"rk\*Ӌ
4��ޙ�'V?����*�l�iM��
�V�`<�w��k���}�ۦ�
�֍��85(�Lo\�1}���:��,ّ�?��a�><11��Ih�g���R�������u���P����6�k�;����C�k���X�je���Yӄ���wGvS�Vv��H��ݪk2%" ��}�f��Ю�eq0�?-b�a_�σt|0�g��ƻ���Ȣ�L�8~6I���4y���Ӊ��^N�O
uf�wW�d0.z{x9�F����SE��V�N��h����+&8:MV���d,�4��'��]����\+�n�oٳE�)�{S&�3�ۊ�=`��xn�oTv�eye���>I�Q�j����ɦ"���1C��Gc�����0�E�3��s��w5j���\�ؾ�U�Nb�:2��͖X�l�d��l�w�SB��^l�܉[hq[�r�ʇH�m{�;��J�v��B�*����v���<&r���ֺ�>*���4��Uq�M���G�ve8Ú!�Y�j�0`�(�)�M�K��ThN 0OcU��������iP�Jl��^@�e��M���Â�al.)aĦvM�C[ݻ��Ǧ��b1$g@:֛�����_���(�ts�7�a�5��f9[9E&s`�.��uߍWz��*�a�3~V(ms����gϩ|@gO��C�9���oz�ش*��'���<Teʖt)�Ȗ�#(��>���-[G��2:~2���ܘ�^�
����Aaq��u�Wz�����3ާU��FDH|6�!�����a���6\�t=���r����7��4v6C[^�.��Kf��3\rLjqe.#�e�:s�zJ�@��+h:<�Y2�/	��*j��U%�����E{P|sޛ���	�^>d<<7�8=�*���@i��vH:�W��3��ֱ��	+�r?O`�y�۫�fM��f�P<����L�r�h�d�hN�S��0stKf��t�`^�B:�Fqu�>3p�����1v��Z�{uP��l&����!�L`�K	�z��^�7R�
�s���_M(�b�;�ŉ���6g�J,��BYL�3t2Y8��s���]|)����b�nQ�\���b$-LP�ru�DdLAuu
�ؼ	�p����5)+�>a
nr��X��ݳ5��̹"�������f���ӸM+�D�?Z�xa]�q�v��E��d�Q������jg��}��m����ޗ{�b��V�M*�8;�rV%�q�ۜ�Qkt-���������c����v���ф�K��8؞/�<��������fH��"M
�7+&�l�b���K�b��k�q�'܉+�a���x�"?|�J({��x��-x{�=sۋ�hC@����������(ڷ�z�V��>�`ϓ޼���Y�s()ۨ�nkM�-uuj� _�mqq3E��5�XE����+|��S�7�l�>�k����=����v����8xGx�c���,��<�4�W�UQ�ӾhM�^*9�dʢ�{���l��7m,�~KGQz��^ V���f����G��t�B���p��إ�v@)�Yz�!�D�E	SG��g�5nQ�nTB��,�^�*�熺��X�b��-�[Po�z�mҾ���p�ˈD".��,���7@�ѓ��ߟY��/����;��o�������Y�R��X�O���wι���ХTM�Y9��M��)�1�5L�2��b}oR�G:=K��"���~����2�N: �@bM!� .��3�牌���d�Yd��w���[�g)r��A&��$�>�Õ�Ȭ�4�W��֣D������^���M��f`��O�('=�/%�[�t5*����paJ8�Fծi�����N��C��f�.۔�3y.T�P���E�e�s{���~p������=�%��]w�m��"������/��]%+ʁk�~�SY�BϨV�e�|�<
��W�J�ΰ���{ά��H�T��؊�O�Q�ï�9Pk6Ǫ�P�斂(��g�ƅ��L8@���LHz�`�F㜊���Ώv����}~�D���3Ԧ]%�+��@dҊ���(�`��%䴁��#/_V��A�6'�#��Ɍ�R���w����Go�~T���֘ϼw!���Zo���{Lu�Q���*}���!��ƌ�3A�A��Or���~���XꙔ�\�,��	����uW]z�uyL�>�Lz��bvy�6,A>��/�L���<uLt.9�[r��SS�Q��yHP��!��&w�[�)Tᱫ���l�r���qm�KřAl�QX����14�����~ A��f��W,��U�؍p��m��Tf򉙵[�{׎�i�BE��o片Sih�>���Ŀ�UA��G_��V�dT�Xg�5&u�� �� X�7-�mK+�+9����#�Ӿ�:�5��D�6Tۨ{NPl�`����x����/�+�J�dU�	��A���Koc�m�&�떵��N��Npέ�����kD�5�؜�󄮐�52o7�so�5�]�$�9u-��,�>F�.d�����1��w���t��O�q\k3]:��Q��'R��Fƹggt��S���mVk�1<t�9ZQ��Ɇ5��z��W*��|�\�ԯ����@��u�engE�F��qE�Rʱ�����k�\e�QH������gЧI;3��9�y�}��G���S���Hz�9�!�Ͻ尬�/����xpu�U��oa�7�5zl�Z��b6)|upt1��Cq-��L�N���#����t��]v�۲���\!�X*!�k"Y�3��EJ�"��%P5c���fk:p��s�R}�s?��4{?w���4���AF�����n�{����+�C��j��Qc3G�j��uWuʰ�N�\��0��#�c���6IBT��BhV�7�	����9��dHxZ쪕��[�i�ۮ��j�8bc�����^e*�z2<& ވNCt�%�n��������#U{�*�66$�C����JȊh�}0`�!����+w�}NVu��z'jZ3)�G�m+���F�
uh��{,�����u�����dL��S��5�xRb�N�J��mt�Eӓ���K���,N/"ᒉ�םZ�k;x��[�z"�ޤ��CmՉ�^���FV��myP�4.�w��VF�Y�k�GC�3п^����tP=��[��]��������k�]{�U��:�k���:�ҹ��R�Sǲ�,�7��3�J��1MΝ���ll2��e�	���S��Ꝩ�Iv��L��<la����5�+ӵA��� �FM:@镲�S��z�B�zN�N�{�{�K��~*�H�m�|q�3aء���b8H�S%�ĝ����K��~�5�����fU�ڈ��ͻtf��S6��8�eԕt*�Ef��S/t@w���f�.�g;N&x���8Ԯ4(립qǭΡ�<��s>*�(dD΁�:/)MŞ25��0���X
��5
x剖Y����:5��QB����3����n6[���ֹ��ՊP,�R�&�ƵWu<��.H<�2��=,W����m�=[^l��Fq��}�u��L�+��{��E��������OH�j��e^|<�MX<4��G��n�w=�4�xW^�}�d]��/�uQ�Po %*]6y��	��:h���M���k7_9,Y7�d�M>�����8eWW��W���@�6˒��v˿���_7Y��Wo��6��.k��֍�If���V��[�vF9q\z�(����\%F�N����6�ۚ8e9�#E*F+�x�^��`4����:2u�A���Ԟ���u�C��tΟFt2�p�uX��a��L�J�P�"��q&G5�ݹۇ ��5\K��]y>3�!_7 ������Aǳ�bf�w��;_3��vêRD"�h�!�2�*�5�"�Z�^�e��($jbE�R����C�.�)��ۃ�/�U�a�I�.#�Q`ڌ6�h�E�Ye�RK��t�v����ICVy����=��n�fs�0�xjJ �K0}r�R�I~.�1�>^?B�=�[x����L�_q��ʨ��:S�ˊ֨���	�^Tg�6��	�UӓF,����YK.�xR���e��]�v�t�ެ"��n�`M�=�M@=��:���u���v�4��[1`�Q�]��Y��\l8㦞:�M���F�3[��T,MrK+,nd194r�2�4-	�^��1R�����
<UX��.���+���Tz�g�t�Ū�g]���nO7}˶��w_`�[�����:��t��!��X������׌g��C�jۓZ���it.�v��qM�Uɋ�����j�`��gZ�:�QF��c������K6]���o�OH��|�^���W+��ťb�5W�t�\��������Ҟ|O_Ƙ�jC�T����
���Y����=N-!�R�j�p�*�v�gb�
D�$�E������:%�.�Q�8wvU�7g7�EЉ�m�W<�Q���2X�յ�^ϥ]e �ƀ�/2\=^�!x]�#�]ݭ��%��}�g��{U8�6���Um��.�肍bH�v�i�Z�d�23���nX��7Td�=!uԏT<���ouVT+N�ȗ,ƹ�q�֨�>�[��tc�v�xyƋ��m����J$����7(Or{)a��콱w6�Ԙ=�,��t�tR��"�Xо�m�P��}㠞�J�H�g�8;"�5��V�C+hfdä���x�)��豟._�7��2���݈R��(<��,y�m�:��(l��3Rb�H2��l&��ԧʗ���]�FD�%/;�����GB�~8d�^�%��d���1�"̾�1�e�9��/��'��(E��8�ݝ��y�ۜ��.{V/�`��g6Lڲr�)v��S%6������"u�~���tUv�i/80��QHk�.��ong&��P�iJF���^v�kU�wS>��G�p���'�.�q�IT�����f�N�Ol��o
}T4�ʪ@��0F��vӸ�|�Ӆ� a��D{(���X�kB��{���,�׋cc��>޷eo�i1]V�B��2�»����p.�e���v�\^̚��G�չN"x�{�M�bx��r�͆I�^N��IG=x��rb�P�Ǘ���U��/�V��y"C�N�-�t�0���<|:χ��j�8=�j�'�9��U\m�c��6����d��\�%k�V
!�T����R��j�(��������3�/w�y��V��c�f�*E�J,�9�ً��b]���R4��\Mؑ��x�ݼڹ�Т8�S�,k�V�'�޼Q�]q���5�,��Cی�rq^�^5�'v���C*��z|!V��;nu@x�������<u����!��}���H�8-.�2��Qi	�B�ȿdQ=�X��d6��8�|k*���*��"߮r�+xԺ˜�`0�Qȉg���l�<n�����8U�@��4*,�{�^��(3�z��}s�{P�YJ���=�+3{@"�����fX̢�jt1:��h|�u�}����N�u�x��e��m��۹nrG��Q��8�fpk�����Y�U7��Ȧf�$NNV����	��2�͊�˂Ύ,	��]R��
z�k++��i�(GK�K���ԝ��]]K7�K���#�`�!v��Q�J�ɨ�\�[�滲r��[#�*N�s����ٵ7Dwg/�#��]��#�=����V��L9]|��MD�,���,s*O��4��\H��8��\���
�ʎΎ��&81uJRV�j���E]I�h�@#lN�y��ܐmqz&8{��e�ݚl������|2)]�ܕ3�҂�Z�v�frsa�{���5F�q��u2>��c��L�
�*��TB�s����u�ǡ@�(�Jwy۴��wU�
rR����-,��Wj�q��Sz�d�)2S:��l�_5�o��N�/�v�r��n��.���P�;��*�A�2[���ҷ:���z���Z0%w��mu0�;�!�ΐ��f�nX�d����?Tx@��� KRjR)B��x��Y��&��i$�+8̖�#�z(ޅ�0�R�r�8cC3���\�`��d�� 5Y��ѻ���q�w�K�o��������g�m���]��d���j���1SÕ����f���M�Ψl1+�ԆM���j�}p�z���v1J�6F��F),�;zut���}�[��{W)i-��oi��o�\E���%�]+�gJ7�hD���bo%��;9s[Զ�0
ّV�;�s-s`�Y�F�N��X�7x{r�Rj��M���s�ձ;��R� q���q���Z��E���C�ђ+{����Ѻ5|Q6m���٭�+�.�%�w��o�ͧ�+u)ÏHvY�K��B\�7s���-B��шvͽ}��l�]���[nvQԳ�cu�fr�QS�]�P��[CS�AV���QQw�2fJ�A�sD7�im�	�����X�+�&��9��T��(.�ywj�Mv���:���Sy�tpPt][{��&w)��(�R�ZW!B�F$��m9z�fji��2sx-�=Q�7�}�gOe<�e�5�*�t�2��g�����wp2S�-��v�yT�ɦ���;|���Q�]h9ל5_���n]�(QMh��~��
�_��IN�Y?ݩ����˸��O�s&���g�`K��/���ޣ��/X�ھy�*o0U�*N�&P�h��C�Q ��N�N*C{�It��:�]4���~�:���IJu����l�v����ٶ�*��l湒��s�ccN'Rqieu���|c��y���Ԟ��r���:|�	%;��&���e���u0��ç�X��uy�}��Ϝ�g[�ԥDJ�E�LX������̬������,*ڣ�ĭˆR*���̕��im��+.2�5U��T�UƂ7.
�R��bD(�j-��J֨)Rッ1����Tb�%L��L�F����TTJʀ�VcU��WS,�1�ƨ*
$K �T�R�j��PZ2(9q�Qı�TB����*9�ƈ���5��fYp�[Lf���J��K�`�im�n\.aMj-C��"4�*�j�V̵VGZ�ek-����Luu�5��f��TA�-��V:�Kn��bX�"�QCL���q��iJ�L�1�Ʌ����1EWHi4�4�\���Y2�p1ӊ��J�E*�u��`�kT���m�Z��麵Y-����SH%�Z�ar�8�mX��0uh��:���:sVZ�j,���ңXi�s
�˚�fXڠ1m��)�F��[iZ6�̶B�(��
�[Lr�+TA�+%�j�`�Lt��fcn��f\Z#t�}�G��@"���&8�z�t��/�Z����k�@�촨��tVۭ[6�Y�駃��Ǔ�ǯ��gNZ��j��wv`#���7ϋq��R�E��PCX"骂 A���Е��)��ևS/���c�`��77s;��c�LO�i�3`�p�R���(M
����&z6hR���n�ctD�2��ݎo�7��/%Q�K����U��A(�����pV}�DR�Dx=A��+"/,��S{36�E�����ڠ��IC�D8��ᠡ���ќ3A� ��-?MO���n�!X=�s������k֝3�2�݌!�>R;X��N�"L
� 6�;}"��&"8�}�
�{���K/�X��w�������w���P�Ws|�ͩ�Ja�d�S{8�~�w�m�=�8���Ug���L����kh^]�g��:I���%]mI7�/�7���1������!���#1�}�
b�線�fVlGeֺ���e�w\_L�tM�G�Y�BE�IQ���5�����f����8ӓuS�05	�����(gK8�:�N�3aL�ț+Fm����bhN][E�՜�Ovv�s@Z�[����y�L��o19�����1o�T((e�VP�9�lh�|���5�����ە�az�~���m�k��Y֭oq\���9{*�9����Z��n����}�Q9h��u��R�v�����ʳ݋>BG�:�-�ɮx\�r�>X.�"�zTAdK�B�5�z����ބl)��!R܋3�m�v��Ce"8>^O��	H����}�~�q�z�����i�8���Ncwe�]�C
���dZ�Ю�
x�APΈ�Lϴ�\�Ka�R�u�w0FWQ�����V�wUbgn�+"�T�ȋ"@�~�^�#�v �3\\��Z�3�5kwZ��΄�8ElS�K�*�ł�1b>���>|���y��0#[}�W����v�N��OS7�˅��h|g�C�x�X>j�N���O ����tۆ��Z���S�9�
��y,&�UħkC��|eU��/yP��H'6F,���iP�����\�ZE�=��X�B��m�ւ���/x��M1���{s�ҳحU*[�[�/A�v�ZQ3�������I|�t'yN3-1�Ǉ�����u�Zj��y9���D��DMv�i�~Js&Z�0ݚ���sa�>��B�D��F4n�vԵ� z�/�՚��7S2fj3o�8l��F��N��n,+-h扫�>$g���ΧTX<uj�;�
;h�]ni�w2n�Έv�nS{��.O�����Z���b��72�hk�5n��=7q��]���]Y���9>|Om��J7���(�<Z����.�-�:m��ȬM�;c��2޼��*6��{p��DE[��m�ސ�"@5����e��]�j8t=��/�v�b�5\v��CM��n�����u����|�BءƮ"n1^#tP�:��OҎ�d�T���M�z������FǷiL1rb�Z8OQє�������9A��?�߯�"֟e�s���˙�˶������ʵ��t�	ÅKC5nQ�nTB�l�(�P�r�siX���o�C=|��^
�j��[��	p8��z���;<ṃw���ͬ]l�c��u�)˴AV1���{x����Ҵ��~_m
D��Ni�p8n�;����(ި�N&/��{"�K���ˎ<5ϯo��EbT�T`�Y�N�rAF|-	$mfxmj��7f:&C/�h_L��.��ꔳ��Ʒ��e�2:f-A����l�mM�p���k���c�NDP� �v`��Ӕ:�_:�N�u�7(saO-���'�a�2�t���ǐι�/cq3el��EؓrX� L��Z����㷗lWY���K�w�����[%�(lo^s����+����{���Oyt�H���b�zy�={*T��Ŧ�B�5�(q�Jl2%_s�IB�N���M�KV�(�%�hX�|��)W˖"ѱ�FUB8�~��^z;Q6�Y�m���[�y˻'`P,�(�ĵ�߄�ԦZZ0?�/�v� �jQ��k���@�
%�Ey�9&(5 ���Тb�Y�ד.s����;PQ��>����r�AGC�T�[��fOt'k$Y���YpEgk����R�}�Ԝ���}qQ���nL�F���и�X�eO�i�QZ�OU�?z`�G��׮bN��{����uí�"v��ԎM|0K~�N�uWr0)��x��[Њꃚc���g8!P|�.�E�X'���ÞZ��x� vs�>���Y'3�?s��qm�O|pt�>��[�_�x���̤m�Ⱒk����,��� ��t�����[�jP�oe�x'i��4�8Ɋp+�$a��1�(Z�-�l;kz�nL�I'W���_9F��Y�a9Eߝu�ˎ���s�*(�< �蓚��_Ea��P"[CZ��]��V���X!.=ƯRF�ٱ�w>�:x�X�ѓM*�0ceQW�P0��pԡ̭ޒԡ�t\ar���E��]JG���b�`���tb�9�em��C�l�,wqo;1���RW+ �+I��[�}�ݫtrMon��C�^�Y��8[�垽TO����Ιw�\�9���G�HyQe��3/��&˔t�^���GLzD*��Vո�R��X��T�u^��V�,գ���tT�v�|�Eu,5��Y�x�)�`�"����b>	F�i�i�9�<p��I�z��˝�$�WuY�~�"S"Y�ax�T��X>:U\<
�J5�O�:��RK�S�9U[�M��q~�F�EҖD^� ��f�����2+��X�-���q�j����Lpw4G��t2��g��$�s&1P�ϟ���@����* ��qM��y�7j��R��.��bu
8!:�a�8f)�dL,�,���5uE�i���+�P��X[4��^�P��\H�LD��s�Fpȍ�K�N�+�ͷ=��hBe�0_l�tdi}�9^졆��n�̉b(diW�/�}��)��y��k'u�����z33���lضgۡ���C¥��Y�S���,׆l����d����n��g3t����y�ԫlW���P�:����uf���G�'b�c�p�fb��,�5�V��Ό7խ�ﺁ&N�L{C|.���������v`܃�f��{��}Oak�c]�]X��+S����2`��%��W՜DW;�����]
��;����=���N�M��F>��𨊧�<���m-����i6������e�X�E�yݢ(s�g�J����0�]�!�f����"�5�z�`'Fꅈ��bk6�u��"��0t����ޖ]��]�U�i�6���sN�c s�Ўl�AYf�bıf��:B@L����͖q��神�q:V��7]�#�AW1�XQ���	�Tq����\�aq��:�qǭ�{P���(g-�E���8�C�Ë��{w+ƘQA�sAS+�!>�<z��,ЋQH٣�UO\;�mƔ��l�NRQ�e�==�؜��˿R�N�u������V���
x�EmC5�D'2��4]��<ΏR��Q�iM�L�>Q�D��H�p����,ܹ}��v�%�>��r�n'�L��؝�*����>%��aV>|>W?���i���j�+)-O��n..]Gv]2*��gO�1�Ȩ�n�uX��a������^0P]@3�u�t�����w��4s�΍����B�7m��ڛܣ1 �5�z�Z}��n�t��C�s��9s)AW(�^��f NP��ŗ;��j�������Q\�3si#� �� ��Ӊ�*���
:��YŴ���Q�~9���R����/ȳO� ���t�t ��^�-`N�\�Z'�=��%���i2�\e
�0k*E�ܷI�`הf�~`+��H9��+��r�k���"���A`��_8Y3������L����M�ջ��I�]�U�u�����PUl�M;؁a�̙M��<5�se���{)P�v�+���\��ɬ��d��v��S���woha�a��Ȧ��۱}�p�f�&v�]QV�Z�d�٩�f�8V��Y��ª�ҐΟ9��y=lo��X�v�n7��ns�%�2���̇��MP�@���q��:+����δ���w:�RK7k����қ�/W�xwQvr�jb�8����rH�HƖi@G��{IҺsu��ٹv�����U�6U&�2y�c�-��'����O.yq=1T)l�(�U^��ڼ�1l��~�AЇЋ��Y�q�KI�|�eD훡>X�8�f�vm�%�_�`9���mgh��녹W31gW&%�;W�gy�`��Ԕ��4���3|�w^5&�u��k������k��8y�-���N�icq���ہ��5P�͑>��8��p:������c��Ƃ�\v}�控�K�G�tI��ql�6[�ؼ �:�� �yf�v�G�MOA��!ϴ1F6c;�ݢ�u�ˢ�4n;�����>�hu�_L�p���~��y�����B��<�c2���fŜ��^@�C:r����ӤxS��|~�����Q��L*:��;|�6!�#���B��Ա��G	:h��k�iy�Ȭm����XI�¬���S.so:[Wu|�~JVċ��0��9�����G�#>4/�e�q2�u>{�M���6�l�u�j�A_{��;IxQv}�h��/��nq�K�̥\�n��c��f�t�qY`�:Is�*�K$�h�I��CZl4b'����f�;��ȾA����B�n��]r���NEP�g�,WI.{i�!8��M�f�p�YPA�ل�*t,��2����c�P�T�(�n��ʷ�b}���۶��.�����hX#�%`���wX�>�[62��^͐����駂R�B�Nf���Æ�V���g=��~6M�r�Y��¤}|-\�M�Bw��4��;R
����0Wt�w����
b 6�2<�i⥕S�u��Y�ۡ��b��N�anK)^��[�O@���y�s{Ո%��s�W�:�o%[|��l�r�b�〮�!�{�Ӭ6�t��Op4 U�k9#ҧ��ѳo����*�U�8�ֶ�]z��Oy!�6r+ʫl���Sj
c`Y�9�_�|~�z��s����t�H쨊�t��y����}�n������t���{<�;q"���B�]F��^j�q{��a�:%Nף��c�X�P��'��dzS�wA�c�X�ک�V��F�O͌��7�tX.w�Um�	�W�
�"S����j.��'�bP.����2���7Cy���v�:��^>1��5�IS��l�k��ɺ�"BH�d9����[NN.��=6%�[�gs�C�B�2�jY��`�)�,`B����x�-�^��g�u涞�V\���Ku�̌xf5��i�L�!3�±P�n��i�����ʫ�=��3D$(w)2��:f��m���b�`�G�N\M��C��rBE�I�\��,��,���2�����=��k9ͻ� �q��qm;�MV;���ʹ}�Ad�{���G-ƹ3{!�����U��3{\��t�f�.�ڳLN(��/r�07SI܆����=�d�;����w���NTQ�o�*�J0%WPW-�Cx8����8���.)K�R�`�5���\M��E\���n�.��Ɓ˺�h9�ʻ�Uq��Yqjsw��UK��-7��r}���\���3dT�I�j������s����ya-ۛ�9A�7��ng؛����uB� �����Mlhcmm^jf%��Է�mwnż��ꍛ~�j����n�\��UR8].���֨*�C�ߛK�=yFB޹��W�S�i+��F���p�L�_q�|��&��r�35KA�v�^Ɗ�͋+�Q��}�ӆ�A|�[���ߺX>٦=w�:Av�Ka�1
��빫��wPV�����p����p�M���������_��EO�J�UU��B@�$Ɵ���"���IqArn���>��Y|��Jk��~��ѣ��m\�$��� $?�$�\��3#��SΩpfh��e����U��R��IA}DF��c>ӻk�_D�74���i`�w�E�.������!}�,�(���+(j*�[ۯ�EE�&�q������x�UA~A`A���$�F_�.��7��_���O:�|������U��$�ޢ�"���~�}���ʣO�%x� ,�2[��@�T�SȚ����g��B��t���ш�4���0Zí��;Acƨ����"��"/��.
b��
cQ���I�iOO�K�qT� �\duQAsl�gyn����qvo����$=�����tB]���������?�ZE��Y3�ʊ�^�]R�h{SKqO�q�j.��]��K Kx>\��e��"��j����=zS4:���{[͇1[���0���1��gT��"�j�u!�#�(��V(�(���O�E�P��LJ�݁�.�BA2*>��D�c]""`}�F�l������(��D��	'�?��D��>3{��V��~v�
���Z�ui	2��V��P$=���".-�y�u�]ɼEE��N@}5����	�{��#V�0>&�p}c�(	ϖ���c�vAB6�W�.OvQ	�O`��ؔ��̼.�}䈠��������#�&IW���$zDPDY_:��X����O3����5�n�hh}Z��K�l-OgK�ZG�{ǟ\�
ۘ����=��q��uҺv�TEE���T1��ޑM'�œ���k��h�Ds�������J�ېl�!UE�X�`؃�<_O���PD^���vv��5�ep!
�N�yҕ,�D�|I�,��k{��ܑN$j���