BZh91AY&SY��K�N_�@q����� ����bE                  {�}�ڭbQ��l���T���SF,�R�	�0�֫kj�*�[UZ�kAe�m�Z�Um�@4�  (   �  ��vՠ)�f�[fm��I$66�M��IS"��M3����B�[U��kmZ�h�V�+l���4�����kY�Է� �r%�eW �]�b6�� p�jƭp =�yZ`U��P���U��D� 
ڶZ6��j�m��f�LY� @�z(Z��P � �`  !��^���:m�n��]uJ-��R
��;�]�n׻��o{�ڡ�]��4�mI���v�Pl�r����ʻ�{��G�^��T6�HaJI��|�H� �}Ҩ������T*Z}s�{wf�4��:{w^���y5J ^^�i*�j�u�z��hQ���xt=�
��A��׸=U^եM�OOJ���;��hP�ަB��mbLɛ�E$� x=	���﫱�:7m׫}�瘟iCE_r�s�OmW`P����N�� �eu�>��Z;g���]�����{�G���:;�R�����=��{������W���ڎ����{G$T*�����l[X���$� -�}������{�IP5}�{�{��m��lz�8=]�_B����� ������>�_[�t��U�w�  k���z�����z
�У�WY6�m��2�i�5F��JJ PP�_P )>��� �;{ڪ=(c}���T
��W۹�h�
���.Ƶm�>��H�u��u�Ь�w����UW�w�xt=j�M��25X�Z�S,j�>R��7o�AA�9��=k��G��4��  �� 4�=y� ��K��X���=w]�@�t�f�eM�ږ�iy�%H��`ws�h���x{��p���sS�� ,���p �=��\�m��g{�@ ��V�l�&�	�ly�)H_  ��W�����P ]�{� ��� ���=�η��.�\ ۻ� ޫ�4h�Cl֐0���Y�T2��JR���� tm.��;��z ��� ��=�x �8@ZX �X Zz�� =�� N^ڊZE�,�mj�l��R� {�h �=� {�ܼ
4�� �=� Ӯ�N��^ k�
 ^���=��C���	R   @ J��RA"*��JT�?T� ��  &Њ~�
R��&&`i�&#�� ��P      �))*�LF!�h��0!�CA&�D��ڧ�4�#!�z� �*=T��Q)�������A�A��=I��~��ߜ���D;D~����$0¶�5%��߹���=�ϯ������bH��	 XHH�HBH���s�Ԓ$��c�D����_����s���g�'��$I��z����4 I�S����D���r�$���������?�_ʹO9S�9c�9NT�T�NS�I�r���/*rǫ�ʜ����r�)ʜ�,���<T�9NT�X�S�9j��r�*r�)ʜ�)ʜ����UNS�9c�9c�9S�9d�y�ʜ�ʜ�ʜ����=Y9SŎX�r����ʜ���r�,z�ʜ�*r�*r��W�<T�T�T�9d�T�9c�OU�,���T�NS�9c�NZ��',r�)ʜ�z��'���ʞ9�r����ʜ��',r����c�9c�9S�9c�NX�NT�NY�*�,r�,��ʜ��',��ʜ��ʪ���',r���r�,r�*r�Uʞ,r��',r�,r�*r��T�X�NS�NX�X哖<s��U9S�9c�I��O�Iʞ���ʜ������UNX�X�X�9c�NUX�r����,r�,rʲr�,r�)��)�r�9|T�S�I�br��9yR���NS�9NX�9N��*r�9NS�9d���VI��NS�9c��9d���<T�X�NX�r�)�$�9NY9Uc�Iʜ�NS�9NX�9Ud�9NX�9c�9d���r��xr��r�*r�,r�,r�9�U9c��NX�9S��NS�9}X�O9S��9S��9^��<X�r�,r�)ʜ�/,�g��������,r��S��9c�9S��NX�y�*r����*r��x��ʞ�ʜ�ʜ�*r�*r�*U�T�S�9S�9c�9c�OVrǋ�����ʜ�ʝ9c��NX�NS�NS�9^,��r��r�*r�,r�,r�,�J�r���r��*r�*r��sבʞ,r�*r�*r����US�NT�T厊��ʜ�\�9S��T��NX�9j��r�,r�,r�,r�)����d��NX�NS�9S�9c�Vr��NX�X�T�T�Or�,z���*r�,r�*r�T���ʜ�*r�,r��ʜ��NT�=T�T�9S�9S��NT�NT�X�Y')�r��T�X�9S�9eX�W�<X�9c�9d���r�)ʫ9d���$�9NX�9S��,���z�NY'*r���%W,r��,r�*r���%Y�r��ʜ�NX�W,�S�9c��NS�9NX�J��)�$�9S�9c��\��r�,r�)ʜ�ʕyc��T�9S�9c�9c�9yR�r�,r�,r����,r�*z���)��*r��*r�Uc�NY'*r���r��rǫ�ʜ�ʜ�,�9�rǪr�,r�����Փ��d�NX�NT�Y9N^UX�NT�NT�NX�X�U����)�r�,r�,r�,�\��',r�,r�)ʜ��9Uc�9c�9c�9c�9S����*r�*r�9NT�NT��')�',r�,r�����*r��r�,������yS�=T�NT垫�<T�r���T�d�NX哖9S�9c��*�*r�ʜ��'*r�ʜ���S�OV9\�r�*r�*r�,���r�,r���ʜ��'*��9c�9NX�NS�rʧ,��NT�NX�NT厊����*r��9S��*�)�$�T�X�z�X�d�9S��NS�O�9OT�9NX�T�x�X�V9c�9c�9c����$�=S��r��,�$�9NS�:,��9NYʕS��S�Iʜ�NT�:,r�9d��9c��NW�')✱ʓ�9d�����,r��,r���$�9S��9OT�S�9NS��Y'*����$�r�)ʜ�9c�*��)�r��,NY',��NS��9c�I�$��S�I��9NY'*NY'*U�9c�I��,��'*rʩʜ�NYVNX�9c�哖���I��)�r��ʜ��,r�9NX�r�9S��<X�r�,���9c��r�=X�r���$�J��NY',r��NX�9c�VNS��r����z��$�NS�I�$�9b��I�#�')ʓ�',�NX�*9D�!��r�$�"9a�RG,���Y� �G(9R'�r��x�9dD�I$�rȎT�XG,��r�O�Y��r��r�Iʃ�ʄ��H��":�RG,C�$rȎRG)#�G*H���r�9RU��#��H�Dr�9Pr��G*#�I�z�$�G�"9dG)�9c�NY9c�NY=Y�'�'��'��r�,r�,r�*r�,r�,��*x�ʜ��',r�,r�,r�+Ŝ���r�,r�,����ʜ�NY',r�9d�����rʳ�哔哖9c��X�x�r�,z��$�I������UT�9NX�X�X�X�O�$�V9Rr�9Rr��*�d����,r�)���r��rǪr��)�r��,��NUX�9c�9NX�r�)�r���rǊr�)�r��)�'�9O9NS��9Rr�,��NY*����NX�9c�9NX��S��=S��S�9c�9^���c�9NX�S��=^S�9NS�9NS�9NX劼���*r��,r�,W��������	�@Q�&`�m����!�*UL�hB��Y���%BҚZ�^�uxUR6�i�{d��-�/$U�^E�2`8�+)L�qU(��!�Q�&^�*Ո�$�K>Y�d�R�w�"�O\XwEn�XP��j�)�km�FKk)�b��?(*�M�n-�R��^�]�r�LY�ZV,B���� �92��}���K7����闅̆=�ksW�T�nP�%Q�u�+6
ו�qX�P�Q\7J����{��e7Ko,��Ж�4F�-�]���y)P�VUچ%d3�^�ںY�X�2���
1H��xa�qI��'fa�Jh��o&��
�4��ze������VkT�3��{���mL�"�J��#|:���A<�C7Y�#P*YBm뙵���+˭H÷a�9x-Eb�6�fQu��E`�bպAU�g�y̵[��ޫ���n�w����l��lnڌѺnĥ�(�,�� �,틹I��ˬ!"1#���Y9hw#�^� 6�����s1:��oL�̞��ͩ��#��]6Ve�d[�&4��R�<ccVzh�Jn�kN�I���7Nؽ�zʣzr���c/,�V�Jp^�wvYpBnZ֥CC2�u)'yS&bK^]�W�Z�Z�!�5f��Ӥ� ��z���i�Pd�b�*��[u,P�^�U�n��Le��/A�q�V�E�Ԏ[r�c����◾å�Ɓ�mf�z�Մ��SV�R�ӎ���4�ɤ�lԙ���vl�� �0����RGP�kF=�ӱ��c6D�^��7Co3t�I�7x�R�!����`.�
�Vr`P�k���h�\ �Vt$��ަ�Gr�N�(n��J��S9�t쫆eԻ�\P������ӚӊUn4ZǶuu<�,=Ǫ��W�;��R[����Ǧn5S�{c\�8�Wx�ŚE��p�bl57V\��8-tN�2�1�X�eh���M�8V�(�ϭ˻��{p�C6=�����"�����&�OKm])A�Ǘ�8�\Օ��Ǣ�^���ǘ��e�r���������4���۔�mEt���7��G��2�z���Z��[̍W�w��sw�i��E�1�t�[kt��-n��7�u\j:HT��(����6�8��%����Ђ���1+�r�� s���u^�o�-̬�l�[
����S�%ᚎ^v62EFQ�i��8mRMk���Cr��ʒ�=��b\��2c+c�K�,� ɒjW�m5x(�-���n^Q*=VE]��1]j���R�+��4km3M!���4��J����TZ�j�������SeΧuL��+s4�&汣p��RyyAK�TB�u���ó.*���\y����p-v+h_�ۻŹ4]ڋk3���M0��֋��.�-�;��C�(<İ!y&��g-�SY������̨�V��i˨73r��ۺx�=
݇�uKHA䆶�i�b��,�B�	d�vo*e���
rkת孹*�U2�V�u���C!%r��,wY�� �k.?'i��kf����v�\N��[�ve7xL��7f����K��Y�.ct.��R���E��=T�0��YCVԻ2�5Y�&Q�Ս�i�x�K���[WJV�-�#e�>��$:m���=��Y�bNΩrc�0=���ڳv�n�,���{�Sf��yg^hJ\B��e���-iy�]��Cu���Bݔɑ�̔��.�,�ym�{v]w_o`ޤ@�ήibT��֎��z�̸4��"ayCl�����"[\�#I��[J2�{��ނ�K J��&%V$���˵6�^��[ke2�n�f������h�T��ffQ%8�j�J�<�{���հ�­�Rp��V]`�[5��.ç�ӍY\��z�@���'lƥ�]Ң6X��H�� µf�R�p���)hU���n��o)�D�v�l��Oe�����P�r"^�cԛ���9z�Ȫ��ne+�q�V����h&fShX��z� �5�f�����<�'B�]l8kj�̷�� �w3(Cu$�Ǧ�P� HQ6�㪴p,�݌��h�7w�I��R�GǕn�z��ef��`0;�d�a��	a�y�@�ͭ¬ˊL�nї�E��M�آ�͙
T/�kUb\�mh�'ٜ/�]n�V(��
��ȜY�272�e�ů\��=��Ǩ�3]�8����X��OFn�li�
q�t�зl�y�q(���f�re�X
9Z���R�C�zfݽy�dc ۫�����Ei֦C����m����kM!7oT�\c
v��k3t[��)��f��/Dn0u�*=թ�ƫ
�K�ն�Z���}3�Qt+)(F�.XP�"�U�ae�1n��2x�j5d'���1��ۙ�!v9m�C.�����Ў����(Q٫cjM��ж�������6ů��_�*5�j�7z��`�a��ܲ��xꂅb����j���xET*��X5���^J�N[D�t)����U��3x�� ҞK"б�b��[b��)6ɂ^�����j��*j�9��ˀ�U�-��R�Q32��#^^��v��z���j�/q�ef��2�HMv�Ӻ�\˧x�����"I�TC|{8�k�]���R'9����ԅ4� �Ԗ٫K[6�p�-5���K��w��x����i���Ǭ�n�Ҡ(��U�h�6dle]�2�B�"R�֮�e�x��	v2�����`�*I�`��լ��NFA��pQ���nm	HG�<����b�؎-�'�v���&�8A��T���b���[8M �)j��,�Ղ���4n�F���ݿdӷ5�(���+�"V�zF��[R�lT.]VG�Y[����N�{b�.�����wx�)�ifL7qA5�IZ�ح8��36��U��Jf�
����Fd���N���ե� ����Ď��6�H%��t3o����@B$Ķ�ɚ2�H.�9��!��z)r�����#�۠H9���-B��ŵ�r�⫨���&
{w�R/o���y0�*m&��j�t�������I.���qh6��Ef�C�"�j.��4��ŵnơ��B��Ne���q8�f���mM*�^������,�9&������.R�{aJ���M��U�^Z«[�h����%�+�"�ѱ��R�<�yf��ȫr!鰍ق��ǁn���	�R���V`(ө��ztb�.�^݈����ۻ�kd-��l,Yon��7t�b�oէ3\��1Cz0n��)5Yݜ��Q�}|�4V'����t��3��1d�-���Vw[�v^�N�D�X�]Z�;(ay!�͍͔2��Q����s];N�YJ�(�Vݺ�̄-��Z�BQ��i)�b7�mm�u��C2�"n��Z�x�fm�3�c���b��jX++s&a��\R<�v���JY��J�/I��8���T�'v��U�U4��zʼV�q�v3��)�V�Ls�l��Y��˴��[vvV*�U,�f^mW*��%���U�J��
&��ؚǐ����m��l��J�5.�M��,ܶ�6��5�72<8�q�L��j�=�S�3nA.K30^�E�l�yZ蜤�%��]y�����%��wN�N�m�S
ݕ���/AC¥��YYA�4.[݂�[Dn�ز��,с^�b��VP��(I�4��2CR��vv��PY��7�,<�س �Jհ<(�yPf�W�L
��6�[6wq_%ƶ��}�z�.���i��2�k�^��`��1��Ҭ�R�f+(��YP��X�j���,�m%/-���0ԴZd�r�$1oHŔZ�Dl�zԫ3��ǘ��b�������M�e�-n*��m^k�\�
�y��/e��f���嘡R�]��-�j���N�Q��8�z�Y	#z�K���;�6��T6�z�RÛ�u�.��̬Ź��B��U$WQUG��iVҋփ��UN5�7]�oV����9�p�R��4m��-��:k��X��������3w1o�Ym�j��z�բ���*�+�˼N�ͼɍ��h��ś�3j�
܂5�j�r*�zF��5bȖkUt"���GuB����3)��{�f�T�l�N�p��C��D5;�;�du��
Eo�0���jm`ɦ�謱x7w0\��
�F�k��EM��U�h��ݴ�n�E���R��z��Ī�YpRǭ�p���/.uj�A��)%u.���x�C��"�ILM��Ul��ݡ/�X�cCk l��ЭRĬ$2���ƚ�b4�˕~l�IW�`Y�3�7*-��y$���%�T�.��#"z�]�Z�͖��j�խ�J����Pu�o	�-\�3NiB��k�y�v�B�]�J�VB����2�v��{���S�#Y��h��#�x�6$a��z�w���Y�ǳ�74�����ZD5H;r��Ă���ĲJ5=Yu�2B�����e[Wz� �٧�� s��V�sc�%ۤ��㹙��?%�EYϹ�L�%iv������eyz��=o{Ik���B��"�d��ɗPʺǁ��/��(���n�2B4�%)�߫e���][ttSrD}�x����;�������v�yIު�ūO���-Zn������ڀ��h�9��͢2�#�Xb(w�MS���|��y��M7B�:u�η(�R@��'+4jl�%im���WF+�l��՝Lüe�
�ՅhIRU��+�{��l��e�ehN��ϐ!�Z��mx�-+��܊�E�3*��WM����;��Q��kR�Z]�����x찤���T�R�W��e�&ާ�j�ST��3���J����ʣt����0fXP�;���
»)�SDx�Bzd�����\�H��1h���u��j�V�Ja�ֽ	�د6演t��Z�kK�:F� ��-ӻ��K�i�`Yv��9eҫi6V^�w������hJw�h��(�&2��6s�/��3u�ƭ��
�IJǧ)GVH�'�M�*F�8�;��h-�ۭ�*�Ö�GZ��-�D�'�5Qtb��QrN����6�5�K�32cJ-�o{���R�檴�i>],I�(����6���Uj�MJ"�DV�\�r����Wk��(�]j�4�Wij�Yj�QU��x�*K(d�o�7�-l���I/�˥�R!9>�RJ/����e>}��ޔz蝩/X�}wvY9E����UKꄵ��U���u�9��`&�J!�f,��V
y�j��+1N�w޻v�� ����+����ս77��:R��T�(�B�j��-�V�D�Ց+]�%��om_(�]n$�Z�OR�\K���U�bԔQ&��5]�K��N���R�z�%��ݡ�4�]+�9rO���O��QsU�ĕ$���q&��fq��&�tN�Ě��-�(�MZR;�Z�iE����q\Q�;Dػ�J��K��@�F����sj�ilO$�[qJ��UiD��;����#u�]��N��ilD�h��4��qj�R%��R�͈�Mbg�h�;Y�9^(��5��u���27y���
F��T�u-�;(�h����T�Clڸ�%�I,R��إ�w"��Kj�h��|�#��NI���4k#�t�j�]�,�]K�0V�Ir�W��7NK�Qm�5��]�b�Q#��V���TĖ���I-[���Rj�]����R[���Z����,�%��Y�J����{�Z�[ZI$��E���%I� �OV��H�YjE"�Y�b��$��1V��Z���\�+��Q_-I���,��S]��s��bԫv�]���δ��ڱB�p��z������R<��ʺ�ʔ�f#IjX�,I��֮���SO�ź�$kbX��%��Y�j���:'��O�U�]�Ŗ12�Tֵ#j%)NI��l�U����WH��ʵf���U�R����2]�M��}�]0�hŜ��Y��q$Z�W���Q'I�:�,���hk"�ƋE�H�t�&��ZZ�%�ԚMX4EV���)U��4��\ڣ�A �:�Z4���ʹ˱�;yl�Nդ�溓�ڪ��K�E��l%�h)�J�mH�(�K��$�$�v(�I�3+���������m ^+o�6��>U�rܿ�e���x�E�$��u�,�/��ϑ��]�)]LľF-K�]SH��m$%)&�4Ԥ�KR�R1(�*-kQe��%�dW�i��
b�YJ5�`=I�:�U��Z�弣Q(B��"w�7�wW���k�<�N�K1o'|�*Yk"�����]WyN��\���/�;��J�2e]rKQJ��$��kie�I�7�+�+F'�l�i5ܤGUݵ�t��[ݪ��8v�R�d��)98�vrP&�r��V�4�ƓG�����Ѭ��κ��V��io'�A�,ԩ-T��e-IUf�y>�w�#�W?>�ҧwX�ܲ��ĝk�K������g1ι�L�i.Sz����v���H���j���ש:�fWUD�(�%˱,UI%��j���R�x�Z�bT�R��`�[�Jo'y���jJ�1#ٝl�Ҕ��Iq�����i�m&�,�Eȶ��g<�-0N%�j�,I�J�B�T�W)\z,]Jj�.���V%�ڨ�ê�tOݭ�|�V�;_)�Q.�rOQ��S%��y�J���1-U�b�ZZ�GVrlmL�T�M���I@wfmTI$�-W;VR�N���X	J�jU��sSԭ�Z�I v�JRC�$K���uv-}{V�֌���%'�]T�Z]�궴ե��ՍZS�$�_%���)�R���4Q˵�E�^�\�\R�����rNLRr�I��p:�KQlV��^�o�h7ib�Pț�9X�R��T��*R�%��5��U%J$�4�&6�f+K��YڼOR�9r�;��KS�v�KT���p��`�X1+�v^�v�5���i��T��ZQjD���Y����#���,D��-dF�K��YkR��	�<Y�-w�"V�TհoI�+	��ؗzI���,�_^�w�����d~=���&�~@�z�;��:�L~_���0���K�5a���=`���<�p����3A������osڵǙΐ�Ni�޾��T
�U'�l��VM֓��R�9\en��7�]�D�OrCWQ��Y3̲��٥�&a�0T�5���Qצ�k{�ŗ�e���3E{+��YBl�[h�gS�{[OFʈ�{	p�`�}�������8���0�����"��K'i츛e`�5\JZR�p�v�z��Ҹe�ۨ�VQ�$��Q�^�֊�p��`�`��rL���̫)"G^��헭	!�tywb�c%C˹���zQ���:q�Ե㿒�Vj�7k�F
ѱv�,��kw�CI�'`\���[���}V�C����
��qm;\����Uc����|
����k�@��9�z
�Y$�e����
,��wfL��y����	Ռ��y�}����=yS'n�Fs"��t/�6ŻW�����b�Q�[.�Ю�o��:�7�����#�r͜j��[*�U�4�\y1��e������%V������^8��iXʇ\���-T��/6��}�23�6!����FV�M>�<��r��ڳ�;�'!f���l��ie9t"����v�[��Ɵu�e��"P_N�y�J*ʳCB˻�.o�e�|��ȹ��n�,%+N������8X0ᶻ=�Y��+��7�F�i���6V�-36��d�*��I�o����d�7���+�*D��»�i��ovX���Z����pg[�8���+����*��f��z�<�R����)L��p[�̨.�r��y�o`��/=�$K1�4YՈ3serHwgN"T��Q��f�,��|���6ś}f�N���'���R��@Rg]&s	}:�آ�=�h��!Aau���qe���J��q��6���-`ӑ�z�:1�d�3�Y�,�#����Χ�'�Nu��C��4��8�^�8n���m�윪�8�V�ʽ �����!FS���{�Kw1d�r�i*�T��;�Gm��2b��vY��&�֧׶�59%K���2³��
��d뮐�P�Ř;\��־Br��,�{v�D�GMH���D��1Y�}�n��� P���u����ЪΚ�[��_JK+�\f���R�^CW��I]�1���4�|^:�����JXnd1oLP�Z� 6���+�]\\u�3����#��ia}R�R�W2��tz�Թ%)<�U3sJ�=1u�հ݅n��L��K;���g5�ũ���͇��KN��xk7sc�y6[:,�(�:ο�;�t���g�Q�5
T���J���Ƒ��EV"`�eN�G*OU4��u:��%�ƛ+"o,�~Sq�CA��""�9w4"�\�Y�Wq+�o\��P�7n�$�CDIVw��]�ױtE�SE=H�Ȧ��M9L�WB�j�K�6��"�ŔA� ���}�An9�/_���л�d����ee�vVT�q�yD��>�����{��V_����7G8n��T��E/�!y��SI�{q��9	�
����y8��܏����T����p�-ÕU�Y��ʗ�QՐ[�d�69˃*�VI�dY��t����vu���Q�}��������8�#���TF��ݹX/!W�r1��%k�w���޵��k&����|	�jr����$��[5|Lz� )v�@4oWz�ڳX�@ӎl��@^���1I�S�i`�i*/�y֑;����i���s\�f�e'���gW750nbI���3zs/N�/�*rӳWa��Ȝ�lآ��Gu���V<�Ԭ%z��崆C�q�C&(�c��Xj�a;:R�gJ��֫�N�C��6��<�s{{�t���櫧fuPz1��wR�VoXZ
������:�VY��S�Qj�wt˵$ĵ�oJt��U.GwZ��j�\��Zj= $��=�^usG��^M���#��'WĽ�ݗ�Ə`}3hA)]�4��ֳi�*�\�[�}� ���6�[�w�l�1�MԳΣ�bG�³5���zPLg=��.cVL���n���&�)D�G*��0�b����[����Z�1�ɭflք�隭@Z��L!uu֍$o1��V��:"
���퀝��;�|z��f��t��}�]�M�ڶ��oB�]�^�9��ݡ���i�/v�8�d8Ut��n�Qe�+����10��By�ֳ��8(��dڢwn�.İm��#i8�얯)�g�#�vT�I��A9�wx�Ҫ�^P���ۧQ�B�q�j����Yn��i�]�Ю��e��=���l�;��'���ϕ�k��>�	�Ku�\6s�4��4A��o]f�Dl�IW^�6#!&nd휫�T$�*�����[�R>!ns��G{X��;*��Nq�`�wy�[��T���:7SX�9Om�f�"��/똥���u���s.�i�R�z\�xy�˔묠BG%�yu��Nܽ�dz��[R�\��
�+V����,��ÛR�d֚�9}Ө��.%�{�n��+\{�����;jѦ�<}ݵ����x�D���³���w�����X�kD��ȆC�c�J]��V�|�4+��t�L�Cf��,D�,@�f���5�����+�hHw`#�ݘ����O$I��v�yɴ��@��9�L�����뒣,���u�E��;��J8�\�|�2Ō���2���V��Cb��9#�%F��N�I��;$W,�3�'��%���x�8����ه���,�&D�*wV��2���˶kN:�Y}t�Ҡ[�:������`��57��f��-�
om��YRrEKժ���=WE�`�8_:b����GT�����^�Pb�0�O:��6��ށ��mVd�[�N+�}��ǩ����(�nh���GM���.�D��;�"��Y�l�^���s~��D�k���C�¨�{g7&m��һ(ݹ&1�9$
2�m�ZI8%I�OgcsJ���k_S�;f.N�b��Ê�c7i`���W���>��u�6�����q�Kǳ�"1&�b��y���zQ�X=s	+P� 1L��o)��41v�<��2��8ǈm�F�y-�P\�
�WjH�d�b�X37�w+�@�˘:fҙ��;3���3boj]=t%�[)�������Ĺ!�4YC'-��/}K"�pH�z[�+��}�{)$F���S�nw[����l�������w�n�������A�#9�g�l����X�m��\�N���!��p�o\��Y{9^��0�vUᬥ���+/�"�U����&����{�^ߦ����6�C%*f�������x*V�[,���e��.��P�=4'p��f%O79���tpLإ�e�.Vq4g¢qc��t��Wa������b��sd��I%�CO��3�"�w��x�N�7�Ē��u]-���^9>��B��p��d�.C�c�����tY���2t�k2�����ٮ���l��d�j��ul:(��UV�Vgd��X�oOIJ��'	¯fb��^ f�[ܰ�T;�[������
�YkH����I�L�gVp����u*�tfʽh��xKlʊ*U��Y}B�x.�j�Y�=�	�7u��!���v��o�aL�a
��lz�b�q��:��G1F��]f>}H�}�6����b�cb���9���K��Q)�Yإ�d��*k[[v��FtZѾy�<���<���T,d�G/:����e
���1GE
&�y���.?{��{���0��nm��V;wC�Q6�@uGO���F�F]�&G.�E��R)y�1׭a��	����`l�p����>�+D��c5.vo3����D kxN�t��F��M��N�;��a�O_Gpue��I�$�8��e�Cs���鰾�ԹXr�4-�٨��ZQ�ۭ6Gb���#������C��*4z�.�I����ޔ���BEe��\e�?B�t
7�Q���aZ���O7�*����As�4"z��M󳦵rv�Dl+:S �\�^�h�k�R�p���K<���l��D�wk7鉼��_L���t�bV%K���Z��CY�9��c%�k6:��5�hS-�C�h' ��洭R����ꃵ9Ӱ�Xj�wm�L[[�Z��>�sX���0#.e���t˕��|��W;�b�݅��H�v���l�W6ވ�r��^��GaW�4�6`5,7�s�q�0�^f���`�:�k�XU:�.Ŧ�q[�;f�bAkN��=���͛d�$�u��$ܪ
����Xp�7�=榽҈uUct�2>�vd�ˍپ9	t[�3׆^���}��1��H�5EG}�=�9���V��##�Ox�W��Ok.m`��B��۶/�U�*ܢ�=�9!�9]̾oRD��֑�3uFAݭ�owU^�IX�GIb@;���z�7G&P�J�K���.RD�J������������̛�w]t����Bu�e:܈_Wu�!����\'
�Fպ1�Z�xL�b*�<p�	�FW`z�����>�ͻ��\O*��M����;�T�F��^
�����GP6��WxY�.p�S��k��k��ڔ�S�����Vм�	4
�}�KL�n��R�0;+Nb�� 5�FLp���/6+��z���jr��FQJ����F]i���R
�Ro�.	SB0g�c�'f��ܶ�!+�hmEb��S����yztot���zu]��E��GS
�}{͐��.��>��pc��;�z6]�xg��m�5
�i�"����M}�àU51V(����':Uv���1ZɳF�]d��J����lmd�B�A�u�ugC�hӲ���;)w�1�kU�8S�$N���t�d��ҥe��&aec��k�"8D]�/-�i����[�7V��fN�yB̼��0��˲�u�L�'s	WD���}�w���X��#�f�wv�x�$\��u9�mĦWv3���9�����ʩӵ�	\��n>6��7&ou��QvhWȘ�lS�MB����<N�ܠq���NI$�I#�NJ)9�U�=�K�}s�����|�)x����"��u6�d���l�Y �w�8�J�9���N���x{�r��U�q&P���s��vβ@�k.�ޚ�T����
�|��G��`�G�r~��,d�<jyn�Xcy7��wA$�7�L}I�ݾ�9̭����!����=�$ݥu�k[s�}d$��;�e�,�:&���{�>�!����]&7���٪�!=C!�3y��r��k'�)�=�6�{�0�d���$=`�Ņq��V@֬4��I��f�6��� �˦H�2�Łut��w�q�"�Ck��%� <o:q�J
B��� pC���.�	>a>�9�>�uN�d�����Ǟ���a	>g6ӛ�[�x�Q� �@}j��5�k�0����ў�ڦ������W��"����yz�˽w����`�͒���M�h��7ή߇�S6>]�X@���i�@���6޶�,`q��<I �d�!�!�V��|�>q�RCo�Sl��倫�1��<���� H_���h!?��������>�O�?��"HHO�?����?�O�O���~_�q����Q�џ�'#*�?NQ{�ӷ40I�lG���],�٘U2�5�e��'�'s��ѱ��5�c�xd�Ƈ�I.�]�V
z��
*�.Ś�ݎ��4��ڵ�*�28�ڨ�1��gp�k�90Y��`O�:l]�9��b܎�nk�7t{����b���Cqbun��̬�{�a*ۥ���vN��f�86:j��Q�7
��װ�0�|C�DWB�L�t3O�ê�uĵ�����mf[�Wq��:�^�.��#[3
U����M�SP�Q+�n��i�������ʊ��e�/QYa��3"�-��&�:cF��KCg8�0NDWY�1�rf��(KY^[T�^��>ՌgJ���"�.�<Cs�Z����jޣ#=݌U����]k��(]��Z(T��v�@�Lv�/��d'.��Z˪��}RWa��ZK��r8�!a�u��yQLcA�����i�W��<f��4;ߌ�L���画i�80�4j�q"��qI�\����{�k�-uK�E�u�dr�_vj�h3O,Tq��c��o|�˅���k2db�u|��\r8���*!J������߬�~33�ffg�33�ffg�33�ffg�339���L��Y���l�x���fg�Ffffff������������������Vffff~��333?�3333홞�33������������fVfffg�Ffffff������efffg�3=ffg333�Y�����������������fVg۞�fg�339���Nffg�>ٙ�333陙����ff}333��������{����{;}�}��ﲮחF/�T�:]f�jj�z'wudc�O5+�/u<�5]Y�HֹV��mWfKMg�r��B����a]-����H�Q{&�� �r��Zse٘�k+)i&��Ԇٱg�	�1X�͑X3u���7!Ӡ�ͤ28��n����Jքq;���8UL|���i�ftӧ�x�n:��㥧0V��R�z�1-���	��Syʱ�,ٍ0��=P���B�y������;F��fn��*]ypQ=���Mv�C嗐><"C��j�y�nZ2��<����1w�t��);�����m��,����0��(�!j];2֚�rN�rgQ��b�i�dQ
�e��Mf�SU�B�[8~n�wiy��Hܛ�^�[c��CO-	�LU�n�t�����wO�w"uِ`̧��
��pnu�ُ����t��s�ٝ�9��^`�8��y��1�"���ukw�B9�oksr��e��W.U���V�k&s�8�4���"�h7�cZ}�t��:�0��,}�����i�;�������g�9�������ffg�33�������Y������Y���L��ffz����ffz����fg�̬���eg�333��Y�����������h�����љ����������fg���Ϧfg33=fff}�3�fff~3�39���������̬��Ϧfg33=fff}�+33332�333홞�3�z��홞�333?�333334ffffg�+34ff~3<fffg�3=f�|�1���M��,���&�uz��:�N׶�w�\i(����ڴS�|%�L�a�2�[�d�7��Pف0��.��m�����0��_90^f]JDa��ls5[*)k;��®,[��\�q��2��u����p�4�3��j���v�%g�PU�xe��^7tF���Oa���7O�1sH�y��A�h-mh����l���4��w�:Y|*�Z�x��ʛ[2���х����8�-[xB:$�'!4`�*U��Wu*!����M]���9��f�W�M�G�,8��"��'t��Z����M_AJ]V,o�ٌPfq8�o �Z�4[�1ZΠ�oD�$�Z�h�}D��.�V��.���L�Z�D�r�Y�ҝ��EfF�q=gr�k˾�>���A��m��n>h�;�Rʻ�x�~)	���E+���\����EYG�JI�|4����t���Jz&�nt��=����t�fo,��ڜ5�2JZ�U'|L+����ޜ.�`PX�eRg[�g������}���~2�ffff~��3333������������������������ffs333陙����ff}333������������efz����fg�����fVfffg�Fffff~��333?�3333홞�33>����������������љ���L�fx�ff}339���333�3333?YY���z���333334ffffffVfffg�Ffffff������efe���w����+��۷�4��nQ�Ðd�j�o
qtΧ���:dIh��TX�O; ����^E�ۥ��y�e��vh�ҵ�^:t�g2vGY��-Ժ����ټ��l���9���H7#Mn�ȅ����hJ�r��<��3r��bGj��X;�G�h걼4$��n�m��Әzbʀ�rP��ɦ-�|/WTL	�*':���/��hݒ�g�wwN���Z���
��b��Kͳ]/�v��]8�A��ϛ�����5�e�r3ݴ5h���%�*ا-��w�n;:�Ț�K�W��󧇠Z���Q����S�I�B��p��X�K���*t��Yq���z�.��wi��Se]��ٙR^A��K���L��܃g\�gJC�wgc���e�"i.VS����Ae��]�n����BlX���r芯oX���t�.�ff����&US�n3�猖p�vyTGE�j���(�K_v­6�k�\�hu%K��� ��L��-^�-ȶ�u�O������?c������333334fz����feffff~�+3333��3333?YY������������������Y������Y���L��fff}339������Ϧeffff~�fffffh������Vfffg�3�fff}�3�ffs33>���333?33333��������������љ��ׯY���3333��333홙�333홞3333�Y��||}�>>o@2�9t��Aʳ,:��f�Diࢶ:'VY��M�Jր8�M�D�Uqj����'IX::V]D�'���q����^we�פ����M (�1h��4n�t�e>r��ⅿcEdҏU<�]��tޫ�Y���{��]S5��}s��99/r��13����e����z �_�n��+u+pS�Q����6���ܡ-U��n�«�&�ה�Ih(��Rm�ܓ�ި積]�W�F2<WD)̪K�a���=U�AH)<�o:M��L]a�5gefB�x� 3��kUv��vM����A�r�@V8\�˂��Nw��#B�ka�X�f��;O�xۼ7DR�bnCy-�ɢ������L�ײ�l���JG�hfU�J:�e�$V��
�g��x{hmA��.JZ�^gR�i�C&1�MbJP���y��d}Ыt����p�����\�z�$��eiwxDαڨ��2Gܕ3�&�ų�kk36�b�Б�i�Q��� �r�;:��ۡ)b��kR��p#��;9V̝M��v-�C� ��	k���@�xxSv+- ���@_K5�ͦy��a�5Q*�I'P��n�Ȱ7a�
��8���/DӐE�kÈ�$|4�"9[��.�g�Y�Ore�v(��V��e��=�k�5�Ch!8����j�!x��XYӨLF���x[j��+�Ÿ��0Q1�h�8�ꨓڴP�˫V���o3TF�m��o��Kzn��TW��ڑ�wa
��I���Z�/�a�e�"�L��8�����<����v/x��W��;g%�v�<��,KЍ��jS�vkVr�+;ETh%*5����1���r1��0�3�2����q�Du���ҠCE٭t�O�e7R�ߠI>o-v�Y��7 ����Y��R�88)�x��-Қ�󕷨�DB�L���B�UI�#�':�4�� xn��:�	7ބ��s[ԻH:���OۥW�r������սƳYNB�ͲΥ�O��b��}ev�{�þ0mvE�[1������CRk����Sܺ���)�Q��ڡ7Z^�����S�G8j��v2�6d^���0�
l�ʗt;s<�=x��CB�t5�xI�*,�Q���#,7z:u(Y��0xy�)�U��d]�n��9��v¥������̭�2ZF�P��l���y�u�6��2Z��\�'3�Z�#N�l>S7/<�"�v���uuyx&�Q�Yݪ�m��i,�Mb�u9�һ�P踷�����W]�Pia���L�;�Y���d�qv�]����]:�Z��v��O�w�\�25Fa�v��WѸ'&��nj�}����(-��۩t���V�1�{�������;y/rq�+�m���L�&��̇Ē���f�"�<�qu�J�N��v4�9��������
U��+"�8(Y
5�:vr��ː��"�m���.ͣ�F/F�	�����wzi��uY�S���щ���YRƴ��ɇ C֠5�M#��j��F����FS�|<bKjKx���e^�N��@��VaG�A}����+f�wW풰��7K�&"R�u�]0�(�Ώ&����"B*��&5�A)0�蠀v1����]6�����h�u�.���ʒ^`8������ݺw���x���|e ����4U��Ho���Y*����&�����2�+�l�z>���1(��s�>�i)�ǉ��5@�'e�Y&�u+.o`�1	:�7B]®T0�צ�I+�.����7W�gb�a�C<=9����q�~y��%�r՝(�K���cV����Z)E��Z�#q����aVM��ϭs�8��S�2U����i�(�4lm�����a>g��M{˳��sS�nQ���t�U9M��LaQ�*��{Qc�0�ɥ�t �C��5�=d�d:V��8�%����,�uӮ����Fj��j �
��c Jʛ��xr����*Ϸ n�eL�b�h�s�{�q�E�!�qu�ix��������bJ>ښ�c��4�͢��d����mA�ք���}�頣m2b��1�E�]K���e;��m�T�3�%������� �h��xS�T��kaC�1���컽Y��mO��֞۝�¦���^R�N$.�����yr!¨��"bG:�P�qmX�N�뗘�nnM+��ǁ�&�Ny풃i+[׊��^n	�4�.r�f�FZ�2�fvr�e4>��T־$��+�&lY;��z��}��
�-] q����0X���d�dg�Z՗����bR�;����_�l�+�-�"��@���Pb�p/�Φ�IY����+X�gL�f��!�o� �b�L�X
uvQ�n�^M�Ms^m�:�5��^��� �D�Iq��0ڽڸ�u
��8l,�N�Zх�7d���-:"���.U�:��s{N�Evq��T�9z0;+P�\q^p��2%���GT��������)�o�H���X�P/JT���NԬ�VZ	Q��Ŝ�<+o��s�zӄc<$�M���3*�d����TȢ���*>ݰ�˧bt���e��duLZ�k�����������X�2R�Zk`>С�wae��5�ޮ�ٮ=�qe)Z'b*h���%�M-�fӥh<8�a�*��e<�0�۰l�ن��&���ƹ�+*�F�\9�dEV:m�1����Rj3q�5Rh� xu��u��)�ā!"7Gs�F��ރ�ö��ݙ��ˆ�^5D��
f>���L�58��q�M�}t�h�w�I�IRۧ��*�C3�o_�4�tr��6��/�]ʎ7N�"���-��]��-Y�2��P7����B/�J�<�_H�'Vi���M�L����	�[��[/z�����7�����<�Fى�Š�����Gڶ��B4�ue�Aw[�fny�!�/����0�Xvv �'Z�lsc�"�d�J��u[ FvK*|�iP�l_;�WEI������˺�$Ũ;'�>v�p����.+	^I(;(])X�l�b�K�	����"�7�����{{]V�E���8e�=�������G��?���R��w��Q�q|Ɔ��1O���KѼ�&�����,�y�iu<�%����GQT�W��dN�|-�����w�z�%ڵ�\�'���PV�-�A�"�9�#��)j�Q��V=)Hlҝ]�uY��۪K�m����.�ab�3���u`U-a]��F�u�*T& u�Į����d�L4�uk���.0�P�u���.�;׊�r��܃~�Nb��r�鳑��ugٴ\���+A�g��t[yrॻ�%ޕ��%Yr)lw�܃:�,4oLM�kR�rq�j�5��F6��4�RĕK*�*�;�by�@���+qR9b�%5t��f��I��E�Qn��nKҨl�sH5r껶�SɏJe͵��]��rI��	uj媂T��[�}���K#�c����Zݵ�\d��P�y��r��uM]Bi�\�����$� r��_��O��������O�#���'�����_�Rp1��)J
-0�����$��`�0�?�T��� �d�(G!��0IH0�>%[���،�Zp�#��s��hAq@�@4A�Q� �l�B�&��#�iY�ՉE�	����jC"�$�a6`@��,��*'��a$YID�m���~,�P��#%�$h�RM��ٖ�ɳF(D%
!���f�2�G	L�h �!�d�	�$˩��Qq�-Ģ��Y&f[L4B-F�!4�f"I�TmOOn&
� *�^~m�Ri(܎"X���o�bz�B�BD��"҅�������H�0	%�	E�D6�$C�ad�Rd�`C=I@�BZ�9"A(�nF�K�@7����܈C��) ۀȉL������J#f���QiLH��d�cH�)"���Q"\q�� �"ЄƤr6Q0���!	
FJb8Q�[���1�~�ќG�>ϑ��K�^�O#�w���j�ՙ-'��[M�ݓz�X���]*�E�\��6���-��aL�G;K[��2�7jM�f<�v�Z����aw��� �l^\ʽ��:1!�u�7���@�f�]���̥#:xm�4CX�����u�$efm��z�]�!�\��{Ɲ�r�|�+�ې�ꏀ�ѷvm�XM�@u�Q�Q5ݧ/�Dnԇ\{/��ݢ)�ݖo���8��R�5�d���D*m߻�NT�6�7D�OR��L7�4��)�:����`<iR�of*^�#��������Z�In *Y�lwf�o��ݗ&�m��1�����`
�YG�بVu)�35���*حI;�;̭�D�&�69T��&�f's����E9�ܜ�9��c��v�U�PmT5�N� Ι�՝�k\�vO�;®�re7�	ˬ����d�L[Ѹ�$'Vt'"����z��t*;ܼ�Z���;-1v�ܷX:�4&�����	𝜎��G��G/Q`��w�˛�N'���	��L�̐�#A��y	P J1$T�' �@��1�B4�>P �l��q�Sq( F �%�K��d4!B��x���-Ľ�#��&�F\M��B!dĠ(BW�H�*QF�q	@�K�DBL�Љ6T��	*@�s�F��#p��b(Io1Z0�i���A�����f�]��JE9�!P'�$"q��N����kf�5���EfѭUT�!L���2"I$��!�"��0�G�8�C���1JH��Q��P�|��܍2IM��~��Qge�,1D7=��\�%B�q٢�)z�CF[(�.#)����E���YfG$��D�)ϣ�u8b�	a��J����Kn[W()jk2覵��S5�ZT,j)b$��ဒ����!�Ԍ&<\)� �L��"4Z�y5l��%�f4
��D�}.2�q0��3m��(� ����7^DJp2�1��,B�24� ��܆8�(�P%�\M�#r'Bˑ"��~Nx��%C�r"�%F�f�2r4�6�fH�F�'�8Z�C���R!�FYHBߌ"I(�*$(I)t��]�+0�9�kE[V��SD*����B�n�)�Bv����V�*۷3(747ZLM�bl�lT�H猍Fd��#A�%�'��*D"A� -Ԍ��2bP!+щ��S���D(F��MH���.2�c�`d��q/ B�$�h��5��[�͡pˎe�4�A L��	!lj�@�bH�Ll�#A��Q�i2�yDɁ�b�͎%N���E����i�B�%�Jm�q��B�0�,ƽ)x%�D>�I�i�b?��h�0�r8C%�Qi�J2Cr(�&`$&���Je���#P4!%�14!"#j(�a��eN{Ӛ�mZ�¬S""-�KV�p��+5�iD`�V�ZXQ{�=�y�����g�34ffffg�+339�s�����~��/�KOPD���b6���h���d�����վx�O=��~<s��~334fffffh���s��~��b�YU��6�l��ZM�r�:��KSێ&����й52Y�S���љ�����339�SSS��΍�[zՃ�]7-)J*�"w~�[T8Ѣ��<���:�~_y�����ӟo�����Ffffff����9�g���B����D�16����q@RB��3����@TL��5��dyLIh#�̢$Z���
�D��t�%Lc�	+�ӹWmH@U[d���q�j�
�b��Q
�UV@�f�XHb
E̍�9cl	1�)�J�S�	P�ZUF�HV(�f#�F���Z��,ư���J� ATYX,�� ��rÚ��B4�$o)X宲��	�])�!Z�Ʌ����Fն[�L��I
.R�N�V����*�d���MZ.$1r>kX0B[*	@_.g���r:��h�\�+Kn������WX��t֘�2��5b%����k$ö�w%i��g�a�_3�]��.E��k0�̺�V�%��ab*���J�h��T�.	`�әQ����5J��t�X�{h�ڈ(�ʚ�2�Kv�W-�J�-
�������D�V�R�L*A@�PHH)zKS�B�fF�ny�E��,�P�Y"y�!D�j���ȯF�DF�l�� ��d�R�2\ �$����૬e����t��Kx��ƌz��Щ�1v�cD��3�;R���%��N����/QBI!	l�ry�M�#1	��m����@Hp�༢�HF�&HU�n-d�bZ�ۆp�Q�T�:*&�#���a0@�	��-BRz(�E2Le2H���d��0D�d��I��0��d�B2�
6KF�JD�2	m�,�5 Y�&�F2�%[d�O��m�RQE�FZuk�]���kq���1�̺�n��{�!�KI�����n�\�֓ug�H�/^�IT�������T��*@�f]l4� �� ��z��}�fD�)$�ᴅtw����el���L����y]���7{�9�?g�Σ��[DY޳�Z��M���+��;j�x��kT�̐J ��[�4∬KR���u*���.^���[��eU�yz��
^>��� 7z��zf��G��_o�R;sW�����߈8��)t��mȤ�w޼͇j{���aC���t�}�Bdj��m��RN���F�@6I�q_����0��[�č�U�u6�+V�x�i��B��<�m&�z��U���9��F�6�	�g�N�
��ņE\�$���}
t�HˏT�.�/����:���-N�1Ad�o��hR�����71����idu:�阋�^&����ɟnWKϏ�ѽ{"��YM�"�s��r؄�Cɨ�[Epɹa�T�V	2��z�E�/���ͲB�33�f�I�@�w�Ƅ���G�@C#�5�u�˺g�ꅹWm{�@�b�e�N�r�1>�z������|=�THKo-V�+;��&�����¨|>
�ill�a����T�~�p����!�����B��q;��S��)bՙR�g�:ĸ�j@��7a�Q�����F�'2Dn��%5�0 jH��}��~�������^��c(p�y�[��8�#3�+V�kŖ���/��p|�/�����AEC:�����(�(-�U-v\�����O67�e��Tp,���s�����*�;�{/�{�Xs´yӈ�Ч5P�q
��;�jy���6��//v��mg���.�M�oO���[x-B�A��3�Jݼ�/�cL �����(>7�@���õ�����Q��H#�J�;$0k�(J�*RIN��ܺ��<S0,�al�U���i:gJ0���'_��i�>p�)#�k@�_���4Zh^��3�I�Ǽ�2_r�ы�3�i�gL���>�i�¶�J�H�KJ����x������ǯG���+�o��J�>�5m���i��	S�s:��K	Y8H���r31>����� �{�<|������.wp�(kH�"S!~i�C��M���.���R�a��<��o�]5���U��9���a���4	S�6��^I�v,�Y��L��c�6���~�!�R�CY�ws��Υ>���f���Zu"M7��\���L�_�Cgg�Q�E][$�O�ע�y����>��ǫa[t��܏�H�gʜ�,�����}����������>za���]��Yc�䦍�k�<��K���
��F������Mײ5�ϙ�Wnk-�vJ<��ɋ2f�#-��,g[O^�F�ǜL��%zR�84�װ����2� (O}���+�;}8]���QT���my�.b�U&�	X��� 7U/mS���s�ZEp��R>�_���^w)�^���dY��)&|2/�<�������s�`y6�V[؃��	D���2�K�Rضͼ5����$ڒ��t
�e�lP��9�d���� ��3J"	΋�o������?{�||||||G��1F�7t��f��[>ݪ�W���鸂*�8������S<����3f�e$d��T�ܨ�2�n�lۿ�M2�ïq�}_]��߻Th�Jw�,���x"�U؋�dvEy<�T�S>��t	�V%ecT+S�t�S��}��c^Ԣ�Q
�D��j�	�Kܚ�8���.�������hZ�N�ީ�Y�©�s��ߣ^�g��Ƈ|P�o���By$�v1h���U�Q³5Pg.�;�[:en�"�}!Cn �M�����#�w��/��3�I=�'��� �w^�y�u����̀Fћ�#u~��!a�hȅ	E)2��-����ݻ���=�~|��E9+�n�\��O:���.P���3z}������5��K8z�"�ye��=�l�<�����َ�k��Sk��/r9j����-�0�����u��y.ug]���,�siIg_ܹ�od3\7�)gC��;��Ȼ�z��9�.�;� q���Y���{�K��c����Y������}֚?����+��^�f����r�Rc�yw7��A�m�ŝ�Â�p	�A˘�b��咳����WÐ��Pɗ�D�w�Fl6�H/7� ��w�Q�g��2sf��|5`��� Y�y� �G5��[��zQi�Ĵ�S��Mb�^��/W���+���joǧ�V�b����=n��V�]�}�kM��8��8�iq[��,˟}3Vn�1�3b��
�r�}9+�%�����\��D���N$����t�>U�1x׮�:[d���aA�42[׷��17[{��DJ��E�բ����y�鿔�s~1$:�{�jZ�zIޙ��t��ig��l������"a��W�B����[�l�}��_���eo �wsX.�G���}ݺji�����%f��cj��Q��!����>��`�hV���6�� �_�2�ZЕ��;~�����gwy1��� �8��6g�1�1|>^V��}0���,�3Rnwkf�/ȡ/i�.�_4��7[����7M҂l�釖>D ͟^G�G�d :�Zt b���U�j��P�Õ���������Gb��v�xP7ŕs���w�w}�{͏'��1����'A�R}�"���ߩ<��d�p6T?����im���-a�Τ�p�`̕��H�`��)�7}�k׾�j�U��`�"Ej�-�+��m��H)>x?7g�ژ���6�+�����7��UZ������ǜ�ȧ��x��]��S�e*~�&yU�]��+0�FkD��Ck�hb�R`n���絳�\Ua��F�jTц/p�[{k��oo������%_�����˄�����}.ee��N��[�LLKD@8��z��U��tP���H��< �y:2�'sF�pn|���J�W)_?_�����d��ò'c5i�]z��{�1;TA�{��4~�I�ԙ���;�q]G�P��>�T)(Q�=Cz��7�+�Dz� �?}���*UA�.�P����a&D�w��ؑsuW���z��R뵗����N�׃�3/��Ͱ�]K�đ����
7cE�Ԗ?����Yl}���ڕ-�s(�[L�M6
�s���3;�Cͬ����}z�(�c���|@>>�x{�����n��RGyH�E�^��^�X��S��p����Sz���&`�=�P|=��z�*П��ަ��:��rqL�o=�m���yzsS�Xq�e�F���V�GA`��/QS�>+@)Afc=�o��ֺ�k�I�b�<,���;���ULM0E#9����C>��h����V����j��j&Y��:6�%�l�حX��Q���.���5mni�^���Tys��:3��cU��+{�+V"d9����)K7}X���uv���]y-����s_�h^E���o�Yd�Ď��^
��k L�x�{T�z-=2�Բ{IY���֙��&����Wvb�w=qY��N��x��\��T��wќk��P�ڪ�rdں5�Z(��1O{[OL���r 0���Nu�w��{4�UK�;pv�o�>�o;��ԥ�G�r��J����;��*��wQS"��@�DXb�c��5y��њ�ieK�nwK��g&';����x�������ꢭw"�h{�]t-�����w��䁍ݱ��L�a\�g8miZ��D6x%z���ϺX�A�����ܔ��o|���I���Nf�V�2�62Y����nҌ���U�6����n�v��-dH�5�N>�����8i���		S�KɖcUl���Q�JJ���L�8F��V��7-u�\�����~yW���í4�Z��l�	5���5T ��:��/vɾ��pϯ�W������C����>/�����+6���k�-g��d轝�l�o�` 3T�ċz���ꍅ��>���j[Y�� �m�#"FAF3V,ܔR���FV����F`�Љ��R���h�6��E=aҰԿ�1�QP��*�L�����HOI;&֯��#�]7�h�/SP3���>���W���8�w�;��G>Y�V�;ں�0�N��%%,��A2�kU1��W��|��������,���w����OC.w[���׶革�\�{;�iϠU�� �H��0�^�s���k{��o_9�1{lF:fڸ��!�9��*����K��[rbEe\̽�p6vѳ�^�</sUܾ��9�g
H�7&K�]P'��t���ݏ�~����7
��.�]�����{�	1�;ɻݐn�>�w�
�ff>v�ni'�c��A`5��[��J���ѩ;�"��t�W�YyF{����n�9�~\���	q� e*��Q�R#��W��q㚖}�9C���7�w�ٳqD[s&��m�J,��P�8���$߸ۀU
���>�V���aܓV�b�u�.ˍ�~:ޕ�^�	��R��P�nL�@0�jX�Yz҄��/�}�/ox���]�� Oj�d\aڳ9%���q{�/�PKO����'i��l�k�i�5,u���^�VᄫX6��nئi���R��G{��zi�+�N&a���t��N��@4�i�E�@�~��5ZlE_K���P}�\��mH�e�8�&3�S�z1ƈY�+s!�fM�z���44�R�(�_:t��5�S���v�AC��Mt)���
�(�EdSf�wa/U��4<�z���N{����A�1�A�~k���`�3�y�wI���*������D{�7A`��	�õ�y2�ew�����<����F�^w�#\W C��_fe�#Ue���ma��-�����{#*[a����o�-���l�57r���$ߓOB�I����b�U���uwXz�m��ufiA�pX�6qN�
�dl�$�t>'�1��O.��ٍ���N%�1��@170M�]�f�V�b
���rV[R�o}�r�f֤�W$�}�AjO�L��}~hN�m�ed�*[>;ƯӔ��=\���G� Wݪ�ӵG����G7�m_�нfA�L��I9u��݁no���o����AP�^y}��>������&������>(��l�E�o�����d�즱���8~܆��7B ? m�!r����4n]���ȩ��ڝ�#���W�!�:�n�@�N�L��T�V&�B����WTȰ]�1���q%�Sxq��f^Ń���:B�7��Y� fc\f�iE3^��wd���$'��w�(�+�"�W\�m��u�[�8�B]�W[�P����V"��c[;٢�@�F��۫sH0�3�x��OV�6K�fZ���Kh��M(N�v�8�\���+N͡�k͢�sVSђ�ۦ��*	:5�2��X05�ෑ��F�V�3=��(�����c
�h��H'����W�${[s����'F+�*��4�����MS�N�'F�r�QK��ښ���XM�w�f���.�&����٫w�zv������;����uf�^�����p�{���gml�j+x�� g3d���
��Rt�X�:8��q�����ݝ8}]a��Tf�i��W���@�[����5x���-C�^�tujâ��B�	�����)\l��m��yQ�H�F��Bn�ݹC��似 
����T,�M]d:�e��(wv@�ә8��U�/��`�_��,ه��
����lY�/B;�f��U�oRw��iNˇԑ7pcUTXKu��J͊,k!�
.ҽ.�����۷��ݭ����(�Q�HQ�@�d����O]ߐ��#	��.O������}O>'Cni�~��X�9�먢�[�6שּׁ�{!����w�r+k�ڊ��B�]j����V�lJУ0���uW��δJ��db,y�F$�(�P���m�A�o�@�Zs)��\�,g�@$��-�o3z�#]]���r�R]�D�Ƀ݅:�HHu[�m���kjЌf�ϸJ��v���i���ҷA��6�c��.^���sx�)����#��ۜY���� $[�V��(E�����D;��6��%��1X#�@浹������28�]�y2���O`f�a�:���{s9S�s�!�w��N���_+���'p����`e��!m����w�����p�z�yc�MI�P�-ax�F]"	�jw-@�J�j�Lg"�}���$/����o���c^wZ۞B.��]�3k�����賶v)1��$l��OU���b��v*�.��;H������k�w�j��䠒��C�J;K���u��N��'N��<���WD�ߊ̎���:��!O�m��	{ς�7k��T�_���|����F<�)�U���P��T�1Ou�mx�8�~W�[e���;����3>?Z333334ffz���|z�x�DEQ`��A�^��[cKī=�UX��_s#��{<���׏_O�g�~�+3333��33ׯ^�>+������ɼ(6�=J�h�e�R�z�H�U]#aTb�,e�1��[|��~z�W�s������fVfffg�Ffg�^�g������,�_<�Ue�`�j
E��"�c۷zm��WR�E]�)TVQl��),������v}>��O�>�����љ��ׯY������-�R�%���iiEEUX(���1ZPZ��
������0��ZcXj��*�֠�X���W��[�b�-�H�ƥ�����ḿWVW�EtԊv8�j}�ekU#[UUEb�J����*K�ˈ�FҨ��q�UDF5�
#mUF��`��,EAq�0ciU�)J�)fP�����(d��ȱ�Tc��c�`�(�T��T�J֫KQUݳ�,��	!P �',fpPsv��.j�v�ގb��g,d��֖벤e���|{tm����4��Tǻ�w�>�//)e�,�����C{������@�d߾���H��NW۸}��i��c-B=����^>�L�{���FI���v�ȶx�śC�S؎NoYKx Cx|X���N�'�5(�c�>|��o�#:<��Y����O{˘ӷ���s{����K������ 1-��CL8>B·g��G�\P��}���F�S�M$K������s���p���K�~�ߦj�Y]ϼi�z��kC�$�>��cߘ����6��r�ԇ3i���{{�za3�g�Cx\9/�L�
O���)�ָ�à_z�M7�;�r{����e�)TAAQE*DA0��l�^�`%�s�al1��b�,lߠ�WY���(��ϑ��O?�@O��pM����d����M~��~5����;�z��x�߯�r}�'�s*�}[��~&�W]�z�h6�3{���ok}��`>R��ϲ�Ny�%����˨1�
��M��^wP�ٖ���Y��x>d�j��y�<��og��}��{�'��9Q��N��ˈ�r�ӯ<�m��sg�XIꞂ7U�n�^���Q���ޛo	O>gS�m�Hh�:�9����2��I���y�ˌ_,�o�b��dQj���\q�L�r�{�L��n"��ay�`�"K���C>�}[���KR��r��� �SV(`��f��M����W:��;ӻs���λݺ��Z|w�/!����U�ǒ^<x����~m����>Y�y��@m+�|���jy��(�?/d 4�s'^�O������{��qw�O��I^��{�{m�x�a8\,�]7�G�=a�04	w��r{������+�k���~*N���b�T���DMQ�e�1/�`|W�����[~�=Zޜ�և�j��`�6=��*b�{�˼<<4,������$�e����O�xn�ķ��>��I�`$�dҞ���=8���ǻ��7�w�Sw���o�&`:n`=r�ǂ��A��4x��G�m��q��q4���n�����$~�=�����$a�����L� ��4+����㎳p���R�� �}Y�B�삔�^�@�|�O�!Q�3�x���/�XF%D�T�랪�a 3gf4l^m�̋�]�����X`|�'�U�l���!�;�{��5s�P��XA��	�+.����y���`)�&o��*�<�
{��>��������=�ꇸ�r���3voy�i��%�	�ލ|�\�
��\Bii�g����������A�\���}5��m ����_段�}�U<*֮��N4�0_��"�V����Y��;�����h���V��N���`x�t��}���5�g�g[ʳ�'=aF��	+*V��p�1W�o�	����ݳ��e�:�;�D������c,��e�V2�,����f�����Qez��]��*Ξ.wC:E�N�YmUt�����ׂ�Zw���6����ɫǝF�Thq����쿹��W��U�������4�}��_�1+k�=ny��Q�^	�bw_�6k��+��x�}�����n�Å8��zm�x�^�a���zw�Z�b՟��R�]�Sp[��W�\2���z��Ӧ�̝$p�.���"���Q|�`<1��Y#���5=���q�^=f���u���ƍ�����"٧/��1 ��ƆW�8�y��φ�Fp�0mp-�#�
��U�p`C�	�Y������g�	R�`&yqU�LLnx<�������͠#��	C0Q���z����Y���֬��q,.��*� Xk_����M``����6

]�Ě<}�ﾚG�Μ�%������˛U�ܸ <Y���0�>	��^���3�3�Q8\_?s���v���������Z��b�W_P]&kqY'��1�u�p޼�;�>�ȇf7P`����FM��9<�8�C	`�CH��x+f��=>�XN��1Ӓ8a�~��(>��O=���P�/�����w�?%�?j�6յBጽ�"t�{���o?�`:�~���	�U�Q��Q Y#����r��:Gߎ�(�j��ƿE?��$u!�r�"5۵&"V��k:=�4Y�+�i`2��1�wrM]����ƍǐ3+��������۳"I��L2`�z�6wv�X�R_�v�5��	h�� 鸲�Orj�.vZ������y���HI�3��$e��X��0��͸E!��ݼ:�����tx|`�d��X��;X�?Y!x9�w�g{,0Y�\�^����{�Ň�Y~��MB���o��L� ,�ю��z<xk���c�:�3�ºn:y��]�(xYU�|�T�ID���|;����Q��iz����^~��y����c��z���jr��u]L�i��Om� ��׷�ucB�r��@�S�\{�$���'�����t2���x�!���+Ȱ{7�՜+�<I21=ہ��Zfz�~H����v���?~ I�L޸"|3Kg+\�I,9�լ+F�p �񉬄�7Q�aKb��\g�{ws�Hy����
���t��oą��9V�+`�E�K��ia�� T�vh�[g�����y�QM����\7�9�a �z�9�\8�����oD��tC�W�4{�<�
�r�/H�9�~�?���5幽�H��K�t�k�f^��l*���.��]{Yǀ���=�Ɉ	�ˠ ��'h�@e�/�Ԕxl�����Rq,٥�ӵ��R��=����G��k�8�r���,5���/:p��0��~�>���ڇsj��S�Pw�fI�)��l�t��=A�ԙ_��_B~H��J���[d^ׁ2s���	)|�ǝu{^���oi�<���Ϣ�v�ve�$QK܉�\.��r�XG��5��pw�]k�[=ﮎO�fJK,��Ĥo?�{�;yk�C�I3�lf�=�_���^_ >�.�~�Ge	<!�<��E���ޖ`Nϯ�ٳ͹��j?�_�{���2���/'s�<y>���½�X;��a�[�d]�L�.�oC���X��=�ޔ� `mO��o;p;!���͛���흉|���Jo� ��s�C��|���/S�~�[��E�<۝�ý���0/�:<����ѕ�ޙ�~��Fgݞ���X��.�fJ�oC�VI���yvݼ��5i}�!8�\�]�k�u�����KƳ-�g�Z��ux��s'o����Ί���8�d����Ml���V3.�L?1hԤﱏe8�h����� ̀32u�X�T����z��Bn�-�h?�5a�@�{��	�? -� ��^�$�BcCGۻu���RJ�]���O�Q�^V:զ��{�|��ڡ�{���T{��C�%p=�3�LѴ�z�8���l��"Z���J$0�9 bzG�Wߦ�����~�����<��-����k�Aw��3ٲOpT�',>��I�����{��b�(؊��c�����J�)�ߍo牺ؖW$.q��Uf
��:Z��}_�e�ӐC��a2����t��ufC�D�V*��g{Gd�$�FŤҔ�
��f��@���4��I�Xh\ ������9jx�m�ۯki��3��e�R2�K,a�?kܦ����ɍ�y��1�`o����ۛ�ύx���8��f��\�^�D��El\8�Z�]E��W\��Ž��x���Ň��^����~� 8��Ev�T0�7��l�n"�oOG�K�SW�&i��]�+�L��^'���G�(��r9��[�1lhnmh�Z빥�T����</ᡸ�yy���|��<6y��8����]��I���^z���T�
�+3Wxz�ŧ��i�d����i�m59?S��<s��m=N=�r�}|UK9W������`*�ϯԯ��#'cS�
��	6[V�;�X�`ΟXBy����]����9���ޡ+Hd�I��Y���W�O����Gq��Ʉ=H}�lw+�^'3�+���{���^g�-����o�h�c�c����&Cʞ w�=ώ�M�f�*�Ǩ�n�<��o�^g�l.��H��!���,s�۴\���+��ff���klB��&捻Gy���'㞙�'ڙ���9n|Rv`�p��T5�;򶬁���<m ���z<���[,���z8m�,�1���հ��)�{�-��b`�v3VB6�޸wm�d�p��}:%��`�'�s9f��݆\����'��h�t\]o
��4��gr�ܥf�/�?y�w�_�o[ޛ�O��e%�2��6�_�����l{����>��^�;�jUG7G�g9��e��)��1"E����i��mJ���a�s�;7�TH�oaK2
�8�����Sh;�{8s����jVmE���?Nƿ�;����3����u�9��H8<!�z ��{��d��v��g"vv{bk/�	@x�`8'Z�W��=P%���{8�ޯΞSӽ��a��@����5%\�f`��á��@M4r�Q����M~��=����@u����="#o��va��ȹ�d��a`w����;�yd'�ew9k��t�%�Ҹ��gi7���氼�4��6�p�e�bp�Rs�}�+��h�{�P����� "�@��L-�_�|yP����40~����=�͸Ύ�o	�zgF-���M{��~�3���<��}/yX����4Z�"o�b#��'�p;�Ʋ<$�{�u5�b��޶���9흀�̈�ɽ���k�N���k��\�Cwt.}hd��'ͱ��l��n{S��N��z`#��~rxk˼ol�m���%x�I/@(�C��s���o�֍k���K��,�G�s;
܀�mņ�Ôz�P�=��'����椁#[�o��oF��{`9RU�%=��Q{w�y��2¹����/���7�0�V��2�]׸�(ᵺs�%r��z�26�:g��7����UM�c;R��ܽ��n��jW(kpT���i���ob�Y��`D-jwq�G�͆J5_����]|>�)cH�{�����{��>�R����<��1��G�0n ��<�K�t��^������8�;�fV����6 ��{e>5����� �c@��	އm˄��/��%�9;�J��2��n�[��w`��#x�x&%�y�P`^a3�O�~���*���/��ʱ NVeGc�W�5������M����@·;˹~�C��-x`?�kS����d#6&�%Y�GO��=3��`� 'P~�A���㼎y`���e��Y��޳�n:�U��~�[Q��x�����5��s�@^*5�����f]��юz�+�<lm�>Ei�{;e��r6{��ѺA�*hDEV�!�C��?��o��^�bߩ�	���hu������.��/w�������ݏ�>��ͮ��E߇�?/�~��*�BO(����O���/�t2h�#:$ʋ�U��gJ�=����۫(q�k|���S�~ (��$�}�����Fʠ������ܮՓ�y`�E��Ioι�~��������-k,!�?/ح�����j?�G�|v*�{W.y��/�gp��6�ƫ�{�v.�Y��٨	����滚�w���iTO�p�Y�'fM��p�Z�%�Ƭ)�7���r;gm���d;��܎�6�y�y��������e��X�Ȭ�X,U's��u��߂[����h֛Y�ď��~a��S���� ����0b�����ۿ=m�zB�y�+��7��+[5;jR��y0�f!���,�1���8���}��XE0IuG�҃N�
�f��3c���F��v�(�-�8�:9�k^O~mu��.|dNZy�w���c������u��M"G:���o������a��=4h�����-���C��'�ejp1����^:��%c�Mr�xV����w�����n��*JZ�}ma��>^�ǩ�s�N�
 s�.�=-�"��ʱV��($��=��r{�\USᕱl#���>����<�>�����ci4����\볠���@����{\�����J�s��gd���|wW�4��\�Q��Y����=�����C����G�F��g�0��=�J���&RSC�@���5�&j��Z'�J��xo<C̰�a��4>��5��K&�8}^�޼t�tW�w}��㠟�e���&t�{t�ckm<��G�4p���Ժ`H��~YT54���,#z<�5TF%�/s�r��mZG�@��R�4��t��7��Z�E�j�Lء���
�n��.�=T�uԜ��׼xMs3Y�S[�mִvw_'S(�H����F��J��KȺ���j�[���u�����̓	�&J�,�Y�	�ɓVH�`�'e�~{���=�ه>�M���n��Ö���`|�osd:�?�)�������m��Q�I���>��zo
n�>��^��\���AI ���+������;u�nk���3��C��\�&>�@w~�G܀�����T/c�f�'�%�7�!B|���L�1�2I�k��l�Z~U[��x�G��` b�$��*�)9�dc&�v2�S���t��3Ɵjx�*�7�)�x���|ab��&��?6��y���W������c����������9yg{���M[�}��Ҙo�Cg�kF��'�e�O�*9�����y����\��qs�|w�5I������Z���vzyݭǞ�-��]3z��LF�9Ƨ���P�MM���t̺8_6���y4���|v�p�t�ܚ��G��C�)����.��6z�7' �O[8x�'2�����ts5 �`'Ln�{�=�2 ��_Y�G���K� ����Ӎ����˨q�ՠI��
qM�l�F]]z�G�����a�d���׈��!��}������}�?r��d�6�������-�x��7:��9�w��pwbd�ra�����1��Y/�
��ݸ�K�ٺ�M9
�}2t�e�<o$
��x\{J�Q�}��-�.լ���&)lf����S�D;j핂����oX�10��۸9Y"�3k���,Y�&�]W� �I���Z�[�E�j��Ϋ���&�w���]f��u�{�#w��J�)�Ce�E�t��L޻K�%�}��j�Y�e+��Η�C���P��rb�ٵK50�e9%��c�y��xma��0o5G�����;e.�ǫ:	����{���ڏ�qn`9���,��q]Q�m��5&U�rP��Di�{��vH;:ff^Q��؝Q2d�W�~l�2J�ᦃѮ��)A4��
���6�&)�WN48A��r��p��j�\�˚��,�;o��Z�s㫢!1y��t%��8$�����wL�֦(8EO
wK�	#�32��uRzT;��2��t2�}�:#�T!�Ӣ�:���찛��[�]�bR̗+�K4CG�C����3�j�h ��
D��r��I�b�isb)��q���-��nꏮ�%�=�P!f�v���DP �*��
~+���A�9/Q9D�� h��5@�@����	�����6J����=E���x�jZ�kq������Q��O��N ����U،��v(Nw�5��j�^�����m!y��x0����'�莜��Ab����Ƕ�J�7��7ׇ��7r�]�1�I�f�7�ݣX+s�;T�B쎏Z';3:�-�����p; p�Hc�.�F�:3e��1[������{L�{�N�Sܻ�71��:�q�N���+���]�p�zH;M%�Vm�$��G�]�s����H���ة��W6�ê$,-����ƻe�^Wv&Y��� ;���M�mf]���)��flj�_[C2��s:L�oH��k^�K�[���;����b��u����؜w$��{��dj��'W]:��g������Ol�¹}��c�#��zLaNn��n�l[V�m��%�i�E�+���xо����2����Gu�t?��z�=�������	�X�_^�ǐ�|0�ޡ՗�4PI��J��-�;�;iJ}�V�S�gXO֭�.ty-^����c��gM��j�҄��N�s(��,Xɸ�sK�=�M0��[`���sˣ��5t�jﱮ���,ܝׇiZ�w4��;�H$�	,FF"��Y+*�<d��]8��努�*��$E�C3o_o���������_�����fL�2{>���,��*�{l1�et�m�cH	mdX����M�˭d�t��4�b��rd�r~>3>?_>>>>>>3�33׳&Ogӳ��@��ő@q�2�h*"��JŊT�TX�k�g�:�=s>ٟ���|||z��������h����׬��~��|�m����hu�cr�eB� ����J��
c,�&�_�����3<g���������||fzɓ'���ӵ�Xv��&j��ł�X*AX��5aSV� ��j�F,E�EU,�"�R1DPV((�`�QTg��d~�3X�V+Y>f2e�EQ+S�*D���ݤ�TX1QV˦ՋX,���,q�P1�PiBVZ�"�:`�`����P�T`*1\���E�`Ă��(
��Ec�ő�TV:j.2�#Xժ*�RDAd<a��0��ݕ�^�/����J/F�d5&I� R6b�q�b�#���IHBe �^� �m�ĉ#�e��*D&�0�(���$x��`��j2�Б�n���ɍ�<�J�w[�V$A5�y���%,x�푊��Փ�N����&�H��C�Kh�K^dD�H�&�*0�-d�j�-�
�4Y�3��Un��ʱ̭�D������P��&	�R�Ѩ��G������"!�$�M(d!��`�bQ���J4�ĉQʄ�DA aB�b5r	�bID؆(�RF$��E�[����07����3W�!?��%b�d��0`%�Ɂ��2X�{�%Q%�$�$Il-=�}7~�o)m1�[3�w�U��\R^C5��R��=����Ơ���̥�Ċ<�.���9{m�hFz�.�]{�X�?��g�$���<?�F�Rg����}*y�p����ؼ��������b�����5�s���-�\pM�p�y��ܶ���ƺ}j�}��G�2��ç,0Ջ�!��P���i.���UrZx	�Q�ڼCb~?Q���
�յ}�b�lCH���_���'�/���o��z3ooVb�=�ـ��}�}�S Z��X���o�Q0���M|���ش��,���F��ӝC���6^8p��2Ho��5��9�����{z�7~܇�s��H>D�g��?�_뿰�Eq��㽲qƜx���;k�#�q&j[�=1�^{k,#h/.���+��%FZ�J
�<���)�_���j�7�?8H/�2����7y�ҝlN[�¡�[;�=۴����0\,A����y/<��s[m^��o�b�\dn?�L �۔6.�z�������K9�),�@�2�xԥe?�|�>�7�0?}u��ƛ���Y�ߨ
 R�Ysb�����.�r{�O�\�aj���]@3��������Mw�(&ya��mz�TDꯖдT���H�2a�)�Yכ���4��"���wq����?������Xm�ūJ����gH��On�R�23ZP�}��a�Ift�-��ŗܴ��ں�*��á��̹n����c�z\�T	�O_���������m�D��x���#�O^+ـCA@�c2d	�d��0��(�Aa!���|��;���yo�e6}�	�I�
��Js�>3��������e~� ���M����7���f����{�/?����7�X��[`�������t�^�$�V��p=
�ƀ��L����8dV�&����'���?5�X߭��JA$�Jz[����Y�ot�xoS33D����'Ӱ^�
���c�g�$�Ł��N��U����ܳ�e]xv.�	�Ma"��*	V��kmmy�xp��kS����}���~�.ߟ�A�%�}���vU'�6��}� �:^����=��zh�r�-c�zwg{�� �/j@,���~�w����>~��*��Ѽ�>o��t4Q�@���7�{��^���w��Y	�q�u��kP�n)ރ ��5{T����-���80���%u}Jř���N8�yǜ��0�s�>b��Z0/��e�k8�{��ƅ�ڴ�9��p1�C�q�.Y�4�"��zz<9��f��<3��3�<�>�do��C4Ot���h���p����|W�@`U�6E�ܙ���M�0�0�����`y�e5bz�/�h����5��AV�yϗtwRp���A��,��������'8�%���3��.�=��y،��7�QDTXͶ*�m�1/�Tm5�] ���"�;.��	RR:d�+Q�wm�dP���t����Zx��� ����M�u��\=�����=${R-C׊��{d�׊��1���d�@1 ����,�$�
@�) {�|���xy"��Ri���y���:Xpna*G����������ߐ���sZ�~5LKwR��\�9o�����f�`Ӳ�MTS>�,?��;i�+�X�'�������h�K��o�=�a�7P	vj������r� |6�����-�O���q�<]����y47y?���Jݭ�y�>b�����z�l��f��G�{y��Jۛh�Y��?�&2�7�~ϥ{�Ip٠ͫ���?����0��<���� L�$�'��A�����¼�-�%]�'��-��nZ����]wpt�@y��-���i�3Q�'E��k�sA� ��K�|��i��mQO������6�j�<�����:=�͓��-%Ʃ��r
�Tv�D<���%>��:�'^��woJ��H�.؞�����OO��|p�l�>��e�`{oT�a�"���g:p��eO��^i=1�ⷀ�Q�ӌ�ޡ���=0������6��0��[3ݢ�Sג�k2]y.{l�\�=��c�=XXHW~V2砟:����@�����H<�d�s��m��~덎x�S.J���t�_��F��n��#�]F�B��\5Y�K�l��È��n.�+������0��l�Y�e������ב�"%Ű�s��qX�rCb}|NZ�+qs5׻����� x=�>�?� ��^�D<z�^ȓږ�'��؂L` ������u����'��߷C{���!�|�P��4n�~�`5\/A��{�ǃ3�z���*g�܍H`l���j����s�ֳ���=�v:r4@7~�I�K�������nb���߂>}h�9��<L</��s��W<�	��7���oG��y�����Ԕ�1!�*�iL�����ɴ0�zLSZ>v_���xC�j��� A2����s`�5�@�!0�������]������gɡ��b�L�.{��3����@�~�a[����2��mfEL�'���\��`/��@E�L���C��r�����H�;ʃ��0,EG�˰����!O>�����0�g�%�l�=�	q \���ʶ`ե�S�4��O9q)<ކ�ڢ�u�)ɳˀ��;�9~�a������[�
��1d�X�QV-:�����xk��O-SV��ͭ���~Y��k ��C��6�S� ]���?64��tޥ�����l��RX{8]?��
Y��~��<��hQ����
�z�=�\�-�s��n�J�s]A��R����)��ղ�2ʔ�WϪd˾3dw��˱�jt`���1j<��G}�܊c�̇ɬ�2�R�.s��˧_-V��j�N>���3Ax&J25�W(k�E񨵺m�����4�=F������'�/��$<z�^�����{$���z�ؒE��<>��_�gT���uU��ɏ��v)���e�܆��'�8�I"9`sЁt� �f�L�jDNu�sl� ��X�(�%��q?]e��jB��u�0�18��Q�8��_�0`�߫����g�ho�̶�����]��~ɗ�b��
��*�����ꦰ��c��-%�y62`;��\�vZ���<���;�|}����k�ɞG;b���m{��a���t"� �;�{0pK���W�w��d+����-^�^�/��	��F=�!���Y�A6�}��G�}�a ,���a!�&-]ᓌ#�=7qN���?
Ǉ�~��I��}o�- ���Uٱ/P��ٮ�=�zO���00�n��{�@a��~����ᚲy~�ci�k��M�^�BbE�:���,�>{�c������Y�|��s��}�.=��>,�:Q����_�U�|G�-��6�� K`�>%MU�ƚ<�5 =�����������מ���{�k�?����}y��o5v�7,��I�ow��kip'�-K2i���hCx������x*��C�\L �ϬL[g=��)�o�f�W����{���I��*����xp�����C���>0�o7s��¡��{�J��R��u��o7�b�.ŋ^�5������m2�F���Q�o]���e 4���Θ�iXk�4������Ѥ6�,���}���>�o�b�~k.��^���_@��XJ�!,��j��}�z�Ci��{��x��EN�k��>�o��Y��|�]�t�D��M�`�V�ݎ)'�ӻ���*��Y啇�]�����o�/��O,I?������^+װ�x�^�A��z��Ȃ� ,������}���>;O����[�J�xo�G
_^P
W��U�F7���a�k��{Uj�<�O�$�?�7 �P���vr�����?�j�<*�����?���~��Ԉ>!�n:��ɼ�y����a��۔���v��ȫ�vR���`y�ܼ� �gܾu0ǅv.�R���o̯��~��n��=@Ѕ=� �����������a�9�?���D�0�M�t��ey�s���Jn/��`O?����)s�T�Z�3<�����D������tPRr��"83
���	�q�^s^�7[��lxsHCX/uc��zw��1xw��ɱ���3CGdF��=��3<�p$y�áM91���+oG7�z�㖡��I@�=0�y�}{yx���t������|�>`��&���R`l�0>�wg�ۻ���'��/�����d�b�=����%��3�_Ϡ�$���?>�����9�ٙ����0��O��M��V��W-�<Y[�T����O����p��|�X~]��!?�s��e�#�Y��������_0!� ���lI����0�j�nq39��z��E�(BV�Ǚ���i�Uk���u8b���R�h��|�øq���ʬ�5�Ӹ���]Md]�no.S��76��xQ��������Q'�U�ԑ�G���{Ql�fL�0`EA`!X��xzz��=��Nj�Dx4��@���P_�}�i��/gT?b�$
�r�*A�+����u�<�xd�)�Q��P��q��w=iW0�l;��D\K`!߁{�[���goq���i!t@~j����a��. HT�T��/s����7{ExKv�ˠv&4:&��6iR+��oj������*��ߪR���!�ԍ������f���DFZ��Vg+�=&$�DL��p9��ߖ��O� V
�O�q�U#�r�o9R)���>vCq�3��1��!���v���D@x�8�m��3�kXd�S�3��^o6�>0㓅���e1�s�$����e6�i���[��{}�C��kt����p.J�����p*�iŻϧ������g�<;�_^S��ˍ�"4I9=����y7�&���#��S���	�кED�[0c�n����z(;�y�$?��7:�S*�U^t����ww^���D>?�v�O�W���Z�*�ΏP�>��]�N,�SG=�R�l�nW/9�����?�
pyۦ+��.�`eO��Q�{��AO�,���� �������)��֤��IR��7�C�1�Wd�ܻ5v�����3�*�f̑�oR�f1Ͻh�^M�y���i �4!��w3�����?Ny�Q�%���%Vs����=��L��	7�h��Τb��̴ƍ�5�������矏����$2X̘��,�3&H����{I$�Z�lB�"�TR�����}��{�&�v�R�Q
���\{��D�w���H��Q�B��R{��X���'�U;������\o{rw.Oo�{�^u�S�C���V�C�)���Lz�1NmO���fg.�L�qUT�P��vYt��dn��/��DP�zy���~ζ>Ě����l־}g(�41�be��p�\���xd��n��t�������r�2.�,��[¼���2��a�2�����"՛Qˀ�fז����5���_�XUxf��t_�����h�5M/���/��onou�ż�E�&k��b�n�}� *|��9��RU����-�x��L��	Vf�([�hx�hh>:���B�|^�s�2����o���,�p't@Oc�A���{�x����3�������6\�0��/a�ZԷ��^O�T���=S��`�93v#��#���-�k������0�v'��V�=��b�+�3�����/�jz�2Z-l�)#�%.ŀ-�l����@ފhdĿ��ɴ�^�я	w�ޱA�>��^�ܻ��+X;�Z/�<L<��R���VzPۛy��F�s�M�)Wf�}���&��3�ԔK��w͔V7�&qz��·+x��+��V�keK�st��8��.ܲ76�l�����1��7�9繯5���H��XI?K�d!�ױ=�=x�^���{${Qd)��X@Y@Rxx��o<}�B�ה_nF��E�@��VM�G��Id���P�38,$�P�^�]��M�
�jZu4x�����!���u��*?����zCqݝ�m�ir��G�q�����>��Aƚ�EZ�S{���uۙ�n��F��yqY�� S1�׻#ä�h�A� [�hŒX~��U(8��1����)%ԖO����������ǆDL�<�z3]����y<��??�����O��4�3B�3����6}��7��*k��r�	�(�����5^��C����8�����k�]Br)Ol�J�VX�b��n�X	]�ް9�BYz����gpN=O�5� >~.%��#,�*���S������k�廝74�� ���O�}��P���[Ol��jL��C�Q�1���F{�ΛO���vd&Uq��f�q����M���b�;ߣ�����s��%�$�~���ް�vor�1�bs���o6�d���s����t��^�׻ [�~]�Bc�b�ӭ�^&^"��#𰂈�|w�	^xV}<+�\C��/�c�������U�=�{��b��SzCo����;����<�>}� �4�+���Bԁ>n��ɞu��g��0���?Wyo�E�;*�����nN� �M����)�]�BJ��-^�jF�'�س1�1��G�� C��ɝ��\sGY	��Y�eR�*�|����d"S��oD]�t84�j��m����_[��������+�؉���z���{$Ol���z�$�ʁ=�ؒ7ݫ_�.����>/��!8@�{[[�ٌޫ5k�?d�����_����5�i�l{if�K�4� ��3z�x��~�^7�5Y��"%_�X-��@����~ť|!}������>Z	�J�ƌ�����sr'�p�e�i�!�̬���Q^C�����>�_^�;_Oh�a���u�M@�5U��@N���Z���Oehk���ׯL��gkv�ke�Y=����P���H�/0���-�~���������:�G'���G&��ɬ";�W>�ם������
ܽ��R��k����������L�딳��2�O#o�>F+��C�����tR#h��k�~��+��vϜ^��j���e4!1�xH�޹�0"��	�֝�2Qח�T���ŽL��x߂�S�������ܨ�}��	6H�����~� n4RwnG}*�b(�6I�׻�p�= }�[��c��wq6��a��u%^�,�5��x^O��O��84�|���Q+[8D��ΐ#[�-�կ-����Ҷ�����p��� 4Y���N�x���Y����*-��ˣ�М+Uj�,Rh-<i�]�SU��7E"e���H�dJ��+	��������َ��0L������r�﫻�56��S^ ��םmod�z�,Ԫ���T�v#�����=5��D\���6���6�JZN ��x�T�bn�Q�v�+e�[�*Vnj`LQQ�m���6�so��y��>#;��-#{�^�oW��U&jv�*c��%=��b���]2��#����;�8�qQ����fKf�մ��ά5��QKWh�^�T�z�X�d��`#���
x�_n>���5k���s8���nt�[�S��1�����9�V�r��v��t�nPGT�۴Zt.;�A­�b��)����r�Y����"D�q�5Z9�p�f	\S��\��;��R��R�Nw��2ӴgpE;���ne�c4��dZ�Ӛ"��t1H�̱J���!�7���b�Z�դ#q�W�H=j
�w�/�T
}�+��wD��&,R�T#���R2����Lߴ����f.ܮ�7��;{gm��u˅W)sq���ˤ"��}��XB�4�-�]Zˀ��œ��Gx_0sf�({5+�S�i�F�h��/jj^Hr@�E�)���SP��ʷ-��'�	.�Lڷ)!#	�6ҖZ'�A�Dx|���f�Үad}�Ј4PZ��×B�uD�򚨉��8*kd�n,�d �9k��������;ٕ���J������_�ԂV���|&�{|#��ġ�IsZ*Ѧ`8�]a�ճE�V6���zX�i,a�O���.��*2���7���acKETSo��
�;p��^��s�$���N,�4ft�yFoL�:�lm�]r9��[6��\�9��Sr
��	,9;Β���x��pծ�_�r5��؋k���0i��Yh9o��PU�
�\�	t��˶�Y�X��"%���j5(�����Y�.zp���͚���6�9sO.�5�x���sȼu�
�)�K�;^o*�m���Þ�x�V�<�B���c���˸����NOwt��%:�.;�[��!���:UqM���6��6���چ63b%�ڬc�\����Ø�vq5�y��A�5�5���i/�iI٥ggj���N�)�ڦ�;5�(E���FE�M�K���_nKsxͅw�\]d%����fIk�y��P;#�i}�㔓�a�✹��V���Μ[2�Ժ���@��އ�Ub��*�0��͒0Y�� �(�ɦJ�U!�VlB����_*�j�z϶g��홞33��������_���|vvb �Yh,DS�5��v��u�`,RM�b��")-�RZ�u��㞾�O����홞333>>?_����^�|~��QE�I,UX�<�TUAE��F-d+�,F�d�����~�_�����33�ffg�>><|||sׯ_o���dZ�_*V����*E�Z�Y�kQ�� k,X,'+�3�����ffz����fV|||}9������ڶOʞZ��灔�R(E}����T���AH��t��]�Y2�SPQb��a����(�)P��E���*
(*��fc��Z���Q�Q`��*��U�B�
H$F	[Q���m��R)Ag����1Q[cJ��$�U"�����FJ2VD`��(�*���Q�ְ�$�DPU�l�f���)!P����㈰P��E�E��C�V�0Ed��,��*�Օ"��Q�*E�� ����}��a%���ts��&�7W:��]��#��U���bxT�[]{<���8s~����:ń�%���d�l��W�dG�U��{a'���$7�����K��u�-2������ǓPlgd�������
���u����������a<�2z����4�F�Z����Դ��yl�S����o���O�9?�oF���[��b�
���qR{oVhqM������u�3���j4���ʦ<5�E���x����o8ܲˉ��՘O�I:k/,�Ǹ���X
�>��b��٢{����pʾs?u�ם?�+U9z�{uc���R�NR�?inV��l�O^���P���}�2��j���0xB9�Mp�]b�k�������߫����A�������1dS#D�]�1��������=���n���8g��{�E����O� S�A� wP�|)�*
~����O3�`����U�uȻ�W����~����E�ҙ�����|��w5v�0�w�&@��?D8~Ɖ�����}�>@
�g�߳xv���j#��4S^׳�,{?g�����鿼����������R*Y������|/��n�B'����[R3}��X�C6q���y�N�3��|����	��������MФw�z�1��swg#�C����z��=�z��,�n�E{���*��r����:=0�v��f���^ˣ�-�M>S
ؒN���P؅��Zu��M�}�y*J/Jo6o&���W�*%�'�x�Ǟ�-z�^�ؒPL�d� c ),�fB�'��7��1y�_��� �o�p�R&�cMc��[߮�]��H��0�{��D	�	k��������Y��w�. ��x3E=�^4[�p8�m��b%t���@�z�� ��P�"��Y���?��1���W4�E�{��^��B1��1�
���_��[S�@��m��=u�EN0�Yjk'�f��e֞/]�p�L�{��O���ypҒ�9��aC\��lSsz�E�U8q�vS���ç6�[{���e������S�#�N�|�?X{�
�.�c�'�7����s�O�	�-׼�;g�3�����)|�s#?�/�C�[�'�U��35�œ����ۼ��`���;�8J�Nޯ\s�~1���;���pF0>`�s������<]|�WL�Ks�v�0�u���\޺��_э�>����Ls^�PmY���[���;g��j�_0{��8���<U���P� 3��8GT���l|k���Q]v��f�	�x3�s�z��_7��%�[����n'�wBݯ���S���Hm���[$k�p����=��p�A�W
���a�*�
���w�����eo�O {=�K[Y�Fq�՚�t$��=����v�>��I�,˸.$>,^�v��Og��^����� ���Yr YfK0��^�z�׏I=�$�$[-������a/�c��5���9T�<�i�1�������L��њa�Q`}g0[�6Įf�Êfɗ�GУ�����6Lۻ�,����z���꧴/��Of�^�^�@3�-�����Ӎ�����u�C
q5���ɼ6B��K�]���=��g鮀3�|'�/�>.Ź��C�?+��R�iPݷ�V�T�������C�g0	>(8A�>3kn�H6�s������3������YY7�+��x�h`+}�+��/�	�.%�Ù��,bp->3�dS��z��$��v��=\��"���3y�$����l�A��{��!�<俿g���Б&=y�yN�y��osa⭫w�uj<���`�o��/����[e�-�j;$.O��P��l:����h��fI+/�X���%�����=��c�̀(Gz��'r��'6��?� w�G��vE�~@{1\5Y������kk��k
;�ϘX���cˤ`�!�\`��Ţ���9w��o0y#L��	����x��������guz��W��/A��Ű�_XY����|�S6�m<��M7D�]�>� ���:_+�Ǡ�g��A�����3��y�7��_�'��;���w��~T���q��J��v�ՃV��Gsv��v����q��s�-����fu��"� ����M�n�k�*�5��Ԏ�̫u%�j� �e-"V��le�n�<6�Cg����>:Q��=_G_�����$��Ǐ^=D��׏I%z���Ԓ���?>��7�������]ٟ�0����m��}�CЛ��d/677t�.G9w���w�k�;�-�}�+-e��[��T�v�k� �#�m�	�lVI`+�wwyhq�������zG\��Ne��Y|L�6��D��S���X=�)��K=��w���/�����\�vfh���q���ׇ�����5���ˮY����72���K�oIO�������mz��J�kɋ�֢s��=B�v��/�L�5� �dҗ��xk_��l&v�Ϟ`*g��[O��7d��	tw��_Q�̎�Ã���v�4�)=a���|����[ހYP�)&>
x�Bސ+Ft¤6��D�a:�D0x���D�3����"M��ϗ,o"P�����F^z*�ds���/J�����W��#3S.{��SCH.�z�������aNM�b\F� 6Y7�4E�3T����>����yo;`��B�)=Fy*�V���[�����A{C�Mk��~����V�\c��.a���fs��y�#��Sf\���^>:�NK4W�'>�� ����,��Ό9:��T�]�r��Ǘu��:���w��H���F9�a+�.Y����$BZl`J�R����-�����
>������[���n3yr���5���{�揄i�ǩ倶>9x�IS����Ff���������I+ׯ�W�^=H�^�z=�{Ȁ=��5����|6�eQL���qi�*�%|'�ޒnm��C�-L��z=���I����##cb`�Ln��eơ,d��u�ۧk��)�qw8�u���6ސ�p-�s�v�b[
��)�r�������`k�8q��-��8L�`K{����/F�=<0�y��{��&3��G�{[�=��z<ng�w��`6�34�v���q�B��0��[nQC�?9��9�gn�p�E�ȉ���!��pw�`}`X�Z��@J+̍��xS}l�*;�
J ,g��N����w{���v'����3�r�3����9�8�w����M� �?�	�o����ٺF.b�5���VY'��L���L9����7nja_ϏY�Yz}����!�M�=��ϲ�EfP����n9?�v��[��E���t�ݿ0����y�����A��f�ݮ�nQ�cZ3t0�����\N5�_s�^iZn��N=`��F=!���P��hCn�_��G��~@c���D����Æ&]�G�w/���!�5�?���w�
7RU��Z̫�%S��3�n�*��,F�2��o��P%�Qv�4�$�6;�����A�<i�Q)v銗Y��8g	�S�[˂�sY��z��W��ͧ/x��t��C��W\p�g������e���3&K.,�%��W�^=BOh-�lO�����7����=�#����TC��Ƞߝ��X�<���[��志��@3�B�˙Z��v�pp!,{*%���;w�!��k��o�W�q�r�G5|��lc���Pח�赸�o��Ƙ��w��p���-��t��^��{�M������<�%� �	k������Y��=��>�	^��L�F���ān;�w���Pqm��Ij������Y���݌<z����@�#­�4c���J��c1����pQM�[�;�)�oq�����\ρU�>��."}�gn��.�Ùz:=�*�g1�k�?>>Xuʍ�{-�vn'��r��'�t��^!{�u ޞ��֭q��/�#��kzq��]���~�,*S���r;���W^n%�=�'��3��O�}�-��C���1�ڛ��<�s
�:��K��x��}Ws��pߑc>�o�<7�cy�fp�ZY��*�XDxL����j��oF�ӽ�7����(糕���Q�c���#���<�h;!���8���jx�sZ���Φ�n��N�ơ��ő-B�X�V^���Ӓ��m���p�7{�m��ի�I�]��D���T�I�7Q����`}�v�(����ˇNuK��􈼄�.ި`���L	�\-S�Z5��̙��[+��Q�`�����W����$�x��ǲ$�^�{W�^=��'���>j���O(�4ab��1W����T��N-b�6���^AK6�����Nܝ����-�uO%'넑4���������c-q-��[�]]������-D���y��C��\����/��[������"���D���L3��}�p��ӄT�צ�1�+Z#k:V�ߜ�m��d靃m���q��9փ���Kx����P� �.5͍��ν�ZJ����!����Իs�G��s���zX�p��"�ky�7[W@{׈~����ƹepE�te#$������?0ϋ��~�B�/B�C	�꿖K�wdK>d�7�����-r��7t���61?����}�sl��zc:}6�ޒy��Ai��摲�*ߖ�3a��g�]=}�X�w���h��� gE���#e�n9kYt��P7�!qf|"�y�U�?�GӇ]|�CD���/)���xx0�!�<���������'�'�u ȧu�꺫�;�k�������G�u�w�s�df�,i �.���:<pD����`�햮6�y����9c�~�f\H��^�UBu1��~��g����bӽ��UMgm<�hX��GD�	�,Wyw���tT�0���kz�8&���l����(n�v��^P>?Pk=���^F;����	�M�S�%�~�³��=�է��x��^_2bE.�ݾ{������$�%�$�?�xC �G��<< W��7��wxV}����z1���r-�3�f9��L4]E�{�66]ͽ��v��r�ӕۮz�}~Uˀ�kk��=C����a�z}�B�:_Xt��y��WiӪՙ33T&w���-�(��Ȯ������Matc��y�d[�^~��/i�oK����v{I��Pl`��V�4�r�������l�O��g<�Ϲ�y�f��B�d�Sl���N�����5���	�wG1��O��n74��u�s�b�w��&	��58{�I%w��|���t����?o�<`V�5VGqX�Ε_��=��]-bg.9��7�����8	�w�G>7�z(����ޥ���X�W2�&��~N���&v*�9�{�Q���o�ځ����\3��bϾw��A��dfH&��&S\mJ�w���(�a؜g2�a �$��Þ_��}V��}΍���Q}���Xvٖ�ɛ�sOYY[���[7�ӯ�i{��ey?��h�Ǯ��5=��%�T��������Z>cYq����}��)�S[sG%����F�"k�z�]��=B�J�ݷN�T���܎�д�cV$k��U���E\��Z�3G��rp<v�;5�`�j�˱���{[:3&�:���:m�� 4������^�x��z����<x���d"$���t��~s]�+s�����5S��s������¥ܯ?1��"x���{�������P�߷5+E���BqB�>"%g?'�P�P��?|�\G~�A�`.�����5y���2�p-����P>c�������D">�8p~�I3� a��.�Q�"�)Uڣg�����0ǆe�Ρcf�\_�k��A~�ey�7ʇ�G�M���xJ���9��Uo-Y4Ńû;��1n�M J���7�{nm�T\<��?M��RBOZ�mNՋ�Z#k/iV�
5���o�~�zd"ʮ�6d���=�W�f�H{j��yY�o;7/��xێ�:�<Ӧ��n�Ic�q�^���J��f[х��-�:��|���Q�=V�����3�:gw��t�cGG��{ז����qa�M��5d��O ����;M$sh���vw�R8��S��5p8O����飔�\��8�j9��3;����δ�z{3j�P��1w}v`|µ�7�w����'�	8��1��L�� ����MVF����G�a���_��}]�|k����=��<rE ��UaQ �����o1mK�w��+6��|�ڲ��q�G:��+�t;�v��|�P%:�;F�7���d���{W�^=�z��OlOz<��{���Ž���&',�ʳ����-D��`�a���/ǴGߗ;�,�V���t��O��ds37Os���z����J�b�zb\0.����le�f��X�5]N��gw��߄;7t��i����X:ݑ���l�G�OA�v6m�u1o3�k�q�"�3+us�^ٚ=��=ʻ�=�_����Ց7�����)���B�[�\�����C����B,����|{r�r���uF2fੁ|��O7��0g�HN'��Owz3���mX�[��xc��Z��n�t�;��v��o����~��n����
�ZG��Ş̾/�W���a9M�q<���fxK6�����я��:��l����On�^Y��9̹˝nw���Yt{p�֐��3pQ@2U��Aךr sN�o��o<~���O�~WT��	���(���L�\C*n�XτW�v�0��klm��	.���8�3��8;g1�x5�xxx ۈ��ܴ��/�2����w5T:%+�-��ϲ%�m������v��g���:'c�5�}u�m!��r�Ŵh��9�,22�/+j7wW*]��99ʫ�B^=;7qU�2�[�§q��N��'8���awAD����i�/o]�Ί!�(��Nx����S�҅q�.�+�&�����������-M������UL�uz��"�Wat����uZ�J�RD�ձ��8C��H���%� �۱�fl{�K{"��ߧZ���T;�������7*\u�f��EJS:�C�T�wk0�{���s-i�W:�"��F`�Շp�2�đN��o���v��;Nf�x�x:���g.�0	]�7�2��R�����h���ok�3aO���+��ױ�/.e��+��C[\ڭ͕��5sB`��Q��he��l��F��=��v"�&�Wj�c��Ai��� �F����ᩒcS�M��fs%#�̠+gJ2m�*��"0u�{0�ж���v���ɬ܏/��r>��=�v�L��]h��%�����6�	��Q�]h
�LĄcn�@�`D����S�aէm*�T#uy�����"'�bՑ����c��	)3����]��Y(�[c�s���,2�%�����(�y�0�E	�})���ێ·1�q&���N�CE�Iǲ��1>	�)9�dT@�";A�_Tޓ��f�[(=
2h�խ�w�V
f�[ޢcFrj�0��4:�涱�2����jf���jF0ݖ�pV	��v�3�mu�%���Ġ���sD�������&���`��1R��]G+�����Cۺ���;uz�U��>����k#���Z����\��w5`Q,;���[C*u��}�I]v�q�v��i}��Y��5���KN��;^�[�N�ۜN�a���s�e��Mץ�(�'��q�&a�n��]R�
ݏ��v��)��Of0:�t�ц5o�ͅң� 8$Ҕ�)[����f6�:/�v�6&��I)-�k�S�	�Wz^�ˢz��I�T���Ǆ����]mk..�Z����n����j��:tF����UZBX�F�E�j�Z�Iuv�|a���k��S�N�0��í�VD��r�2q�F�o�*��A��Ώ������f�:.=���ͣC3m4s�1�q�1l �ʱ
��x�7� �K���Ÿ��4���]v9$JFL�;�ښ�� �z�D 
��c�(�����DD�ݛ�uSLJ�d��/�9���33陙�333홞3?����|}?$��նTT����m�R�e $q���{h*��+**ȧ�,�}9���|}33=fff}�3�g����|}?�Դ��O��=��Qx���H�E�--KfW��s>����ffg333陞3>>�Ns���'�~UUE��T�{KE��iET-%��S����{>g333���������s��S�q>JΰYQb�
�+c"�0F"�=���54����H�(�J�"�H,PQUQeb�]�)$�i,pIU4��*
�i�PD����� (�" �Ҫ�*�Eb�B���`�1 Z�dPģ"�MM[�Ub�X��j<B�v����
�+V(�4��
�%uj1b�La�4�B�Ab��RUb�Ƶb͵1��AV"bQE�y��kX�f�0h$ P�Y��^i���6�&�MZ�Tut��Z�TGZ��Qb��F�I�I|a�=	5�@�ߒ�g�I')��,8A�!<DF6�pl=��[b�)uv��ɸ�摰��|�$�Ȇs�2�7��o�Nq7j9G��j�){��&�b9z���V�̚�h��Dֆ��L�g�( i2��8��$�b	~q���E��R���%(�Di����DF|�� 	���4�ĚqƐq�0�+�&���)6�Q��1¼R�̓Ő�J@�E��-��D��.A�(	pI�M�%MM:�t�6�V�W0�L����aI"RP%eF�j(|� @B3� �I�<sǱ+ׯ��z����Ǿ��π��\���T'P��~�U������ި��=�xX꼺���������BC�]�}���a�dF8t\~�ʵ�Ũ�@}>@o,h|oՌh����{�y2ڜ��y��X^��ɮƨ|׮ӝ��D~�?]7�����@���p?c
EF4s��&�[6um���fwa�qo7���T��-�j�f���p�a�@Ɉ	�s��.�z���Y��Vˎ�����}m	O�e-�����[u��y�8��q-��*x��7j���q�e��Gz�1L9��E�OB������/]����(n�f��]��]�5�k),���{����nQ��H�ˆ%�G��I�_��*�[å>�3�T��zz3�#��*q�æ�d�'�2���v��,��hlz�c0�ήr���#y�v��[�`�)�h��!���qx�;Ǻ'Ǫ�������8!��R�x���m�i�P#F����������
���� ��{�c]߲�E+�W�|G̼����w\���7�rҳ�ټ�Xs�����/I�l���|�y_��F{'j����<ǯ�f������gC[�-E�wY}�Ș����S�O��+�w�V��/pW��vnR`�W�l�}�X��f����_Q�T�H��-��IrE'BwT�'N�\�Y9#�2%D�:E���".��yo�$�_���ԕ�׏d��<z��{x?����x{ye���O���T숛�"��0oBC�{�r�L��w��hP�T�Lou��J4��9կQ�0�v�yj�i��ެjn�<%����B�=�t*w3�ּ����8�7I��/߂�Ay�@Eǧ���;w'˜@���[���-1n��vx�蹪���}�ާ�x��s��*^�{��d/U�W���~�~�Ji]0���n���\)	���ǀ�U�\����w��R�d?	q^Ǆ�����24�(��u��]:W.��y�Y{��k[cV�J�>\;����A����ǌ������/;�C���X��=��X���h��i��.��x�,%;�pt�<'���	d^˵���pO�K�<��!^��:d�!�xoDPh ��"��[�M#^w�ǽA�;�n�4��m9�Non޿i=8 屐l�\8ր��%�(�E�hm�f��Дn�'�p�*�h�zg4w/�>0/�w���������k�3S�{
_�c�[	��y����O$��>��q=t�U�a��w������t��mƇ;���ˠnB��y���bI��w����R�E'k��d��H����xk��>w+�}�)����I|U�Mq��e��\�{�uH��΋][ó�5M����^,uo��\�ׇ��x�%z��ԕ�׏}��ǯ�X �y�aV�Eᙗw�w���;^yxp�<�:t����~���Ƣ���&�R�a�,Tn�u�u�fr��Γ�lzg���OA'^z/�{}���̂���/Ǎy7��ٸ�,.���m�H��΅��(.�G@�a}���Y��Ǝ�U��`շ�M3�=�*��;g��b��VN�f��ި�n��.��>4��vnm���l>�^��{�zUͿ �����.�ޗ���ԉK�����G��}K}��������������=�AiAܩ��O��;h��k�S`�^��o�'^7�C3��wvcB�Dc/4��SК�L��j���)�Ѭ$�� �5���6���,1�߼7���1e�\�W��c>��<�Z�;y�H���H/�m�=^��\�����Z���F<g�i���0���s\X@����v����@~X���e;�=�:�U�lѸ�wt�&i�����o�/4vGu�U�%��no}^�W���3�>[�?��t@��jv�׽�5�w���O�4u@��o� [�~oQ�!P�=��~{��ȝ�XU���7�F�J�r��u*�9i�a�B��l����5�(]�����N�>C_(�BB7�m楊�l�aA>@^��
L`�b��E�u����{9��+Ι0��G�t6�A�Y�e���`xm����i��퇙�Nr={}�3^%/���׏ez���+ׯ�z���$����_�h\��������)ϙ���;�����zEs�\��(9�.�#�w:!\�]i%E�0���`Q~ǆM6",%���cO<���w�%�5�*	��I�������;��VY�o��!�;���z,��p?=�֘x�x{���\�
m�,��^v�[�K�9m[>U 0L��6"}�}�0,���0N�aG��9��S��_z��pJy���#��i|���V�>�	_,;�>��=�Yq�s���*/�o�1�}G����N'�����;��~}�L5��{k�y���a��nx�n��9�8v��"��MW�]�k����;�7]Ԗ	��K\rz�����Ɗ����TX[Xc�P&���'4��tzdE��un�L�ǟ�5��a�,!���6]�LQ0.;B�ށѦ�3[�f7�p�q,Cϣ�j�4Kȇ���j��X�Sȕ)�ձ����I��Q�T�a�-ؠh({D���x�lg�5=�A��$Lņ���ߛ*�F�߾�~�&����9� ���J�c�a�[\��i�n;leu��ћERl+���97�n�2��W�R�'��Z 3>��L+��Wr�|�RQ�W��^�x��ڼ��Q]��[+��&�M���f�]�ff��痯����2YX�,�fL�d	�=-�̟O"7�۹d^bW.�o��㐠g�@��苷�m��;AjK���<�$rl	N{u&�߹(a��~�8W��x��3q�XYUa��/�
�� �XN���nrv�L�?�F KvO�D�{(�QcA�쎂���ޑ{Xy�f���$[Vг����X`��p��&�<�,I�>�=�~3P�o\��Bޭ�n�����W	���:�[���w��6�z-��g�DS�u@��	�H�<����=};�������g�e�$Ϗ�Z�M�#B�~_��Yl\S��\n)m�䰳3v1��@0�-�}v��Mx����>jy�0~��\�Gk6��U{+l�#>�d&oM�dN9�T99�̈B\3<�1����~�c1���bj��Q9�K�o	\:Qq6���p+�Z����C�.�b\>���[wsV���|�Zv9`����ئ̬k�]�f
��~�*�+�; �0_�$��9U�i�u�X8���SӼM�x�7�fo	�kˬ,��^���fz��{y�g�b|����a��,���s�X��~OaZ�z�{�#)��&����M3�/����q��K��f�%�� ��눼��w�ﮍ��<ޝ�ԭg0�TQc�SZ���J�)oy�o=M���o_	�vu)}Y]��]������i�OsL��w^�H�yv����I�i���?�sǱ^�x�J��ǲ�z��=�o��$��|X}.3�@���B����C.�Z��1�ߑ�~U��4��[R�=�����"�cp�rt_�	�3��X4��N�ZbY���u�5�oP7����󫛝��f=֒�)��G�
'��������)��a�Wଆ4/�o�s����0���75�\Cȩ5�x��`��{��Ѯ� )&Y��t�ޠW�
g��g�!�[�E�k����r��w�St<���1����q����>C��5�;�}l���o�g���u�νG�����:��x��!���~ﾞ�Z
��Ę�4����b�k�*w6��/36�!I�����RLp^Tuy�o����K~����� �CſVt��\����ܼ��%,�Tg �n}W/Eٟ�.Xp��I2l��=����p0ϔ���Q,qD���5�x���sՊ*�|�՜�+(�B�&?��W�]�����%��7Kھ�kz2>tݹ��~�<پ�궶�ܑ;���~��O���
!������+�ٻ�ͽ����z&��I��?��δ�*y���ll�A=NJ-�n͎��Qx1��(X5^��Sm���tWV�X��1/��Q��qD�7X�-PwN�فo0�x�Ő��%U�l7wx=����/0|����>~~C�����ݵ��WU�h�w���������SΧ�@gM�!�����ޔb˵���ȶ>h&��tf��A��V[3�s�w�L���x�$�=�ܷ6�<󁨆R9�f�F%�?1�L�����y��p�C���¼=2.Z7Z��M�k�����s;H	F멝�瘎���w~�o����?M<Q����2�	�����~�#�#`y |���_�ɭG���n�e�޼yӮ۟F����qx���� pp�쟋�cr�'�*!�j&�<����h���ǭ�{��v=�������
���^3i��^yx'�x��6i���縩�Ύ��=;�ښ_{�D \>�N�!���q_��P!�X$�J��<��.�E�O�ĺ8/���WWu|�r�j�5�.�x�y݆dĿ�� ��z�&�to9Ñ�;�4dA���x���yޟ�8��[�	>�X��K�����L��zE���س��^�Lڹ�\p���}���!��
;�R ��V���;q9C|e��~?c�+�%�G���f~=�k�w�"�%|�P�T���f�ss�w���P���^�J��ݧD@x��$"���qn<|��� G�W�><-}�%��
���稊Q(���S�2�NA[t_m�tX7����Ǻͦ�z{}���{<���?��<z�^�{+ׯ�^������P{��a��Ŀ��{6ʌ��#TJ�9
��ߟ�7j�O�_ܮ[_ar�d�5w��w���vv���;�����ڃ�Ej��N,Q����
'����w����D������w8~��e�XS�=���c�������Z���g��y�-EDkɩl��F1���������>���:��@�)��	�E4w"%��ڶ��U�yoc� ��5�q0�Z[CP�#���'��eڹ����tv���IŹ�������%��Ɓ�F4æك�?�&����Z�ݮF��zWT��W5ڜ)_�?�}!�ߌϑ �&�������ɧ���<�fY�:
Xs3��OM��p1<{�@`�X�*���!��;���ݮ�`shOǚ�l����<N^�8����c���ΰ�o�������<b[�?%��Z{�Һ�'��?t��'F)i�09��"-�218���:����^qyw�ᚽJ�����w|���_n��w�l���t+srM
B�kL���k��ȹ�;��݇6���;ܻ��> a�Q*��6��gJ�`�9f��r�)��f���;m.���!�S�wU��9G��q���/���^�x�^�x�{^<z��"%<�n�2RQ�/��+��UMbf�\���c�%��b����1Y[b��%�MZ�N��
���7�����i���zT�$j �A�񂬮;R$��\�	�=�-��$�b�ր�i	G��I�.4�������y�!��'��d�~	��[kj2~Ady#n�O��v��v%ߠ�v*�E���8P�Dg�bqL,c<�z8;�����yOl��h�J&�(/��R�m�'�X��y��~�/ؠ&垇lZ"��N�w�ٕ ��;��HzN/�,Ot�y�^����f���p�%����߃{��e�d�1���	$׬��mSY�ai��1��;��2�YK�-}���q5>����a���ͩ7˟t�|n�f-R]�(/�����ٻ=��"���Sry���[�=��L�@�=9S��F�9��t����Q�7����1	�|��)�b�!*��8=ͬ[@$E�zDF�Tzu�dc�}�#G������qT�Aq-�N�k�x?vͥ��g綷x-�s�{�h~3(hs�߯��!���:=)�7�f�9���x�qn��]N�΢�O�܁]δs�>�G�'��` ��'�`�� �7��f�E��*_���x�6�C-�ᔝVW7���or^f��}�0�|����bfʹ��m�Ϩb�ǃ G��#��{�a�,��.�r4\�7����FP��p���}R�H߶'��2��*K���6�����=W�^=J��ǲ�z��?�����"������~aZ�+`�m�d���J����נD;�{i��1%�J�/�z���Ϭ9M4�qc��p+�Y'�:�y���ы�zU���}�ln��~a����!���!��������?���U�ե���)��x�'�w�Fv��vI���>n��K��¼ޏs&6���-�K���}l����	4�d֬W݋+8O�l�K��8x��1�$.,u�~4��x��� ��֝9���r�K�7[׹޶����������N�_��|�k�U�d�땵�Y(���������������7�����Ӷ0u������y㦋��]�BdZ���ZO������Τ	�U����y�>G=S�����^�U嗏
c����E�Պ�����!����>73�S�̟R�4��;O��𭑤���kܷ?�������0��5��;��G4��5�t��9~0v�= C�:��X�4�M���@�����N� �z�?M�8���:��|*U��F��G�V��١v��Pľ�ݭ6��t�)�s���4ӮHb�N�yu	հv�/-H�����#T���FAɅ2�ul�Y{:mM��6WYus�V�����qƂ{�"��7ј7&i��c�Y���ҫnؼ�L�у��	w�z�`������ub�ɲ�
�ʗ֋L�ȡ���5����Y�C�'n��w��#MC�n��`�6f/@�Aҵ�{g�n ����Y��<��m5}�zhY���Qm�7q[ۼ�¶����*�Ԏ�b�u��W�PLKt�v��,c��Z��7Ε�Fi�}o�3A�KUtx-��t�;@���K9��-N�i��my%�����qL�{H²��]�GVvKh�2Z��uf��C]���t)^�9���#�����<�+���fG�Yͨ�Xk�:]��_E�h�K�j��N�8� F�*�%k�J�2�ip��=��Q�K.�ߙ�~ȳ8�W|��%�s#{�ػPC�8��'\�����.͒�#ϫK����R��~��V~��5	wU�l�>_c�9.��w[�>|i�����GwOY�ʒUB�8Q�q��(��(�h{��;<S�Ĝ��֡NcH�;�-m��V�[��OV2�0 )C�\-K�bp��R9��e�}���|��X��/�ì�״`ye���ߔ��}m5/p�[�],���Ԣl��Q
�T�F��ܺ8�,�kBTׯt�+���(]���Y0$q7A����mH�O�F���=~OO�,u���Ccz���]�Ӯ�X४{;gq�s���:�K�5�V�s
�ṷ*fq�WL��,R���F+��S���b��%���J�1ʔ��6�Jv���UϚDK;}��c�.�M�[2�xn�+���%lv��IE3:��O:n�抇�R٩QmAv*�K�b��{y��c2�m��w�^!%t¦�Q��n`�Zp:�+��tlM��:K��H��ݓ�����)g���u�gy��LZܖ��������u�>��V@,�/ZޔdM.4�"�Ao��NN���A�);d����l�ذ�ۑ�ξ�u�y��h-y�,!n�}kEuā�λ8���Н�zc��Am�z�T9o�䘗��_Z���T���!�ձ�:�(#ډ*������t�tq�|���o=���y[Z5�=�Ww����u�Q]-����G�\�M����Z)А�S��ݗs�	˄�,��Y�M�'�q��6��v����#Vyw�PɎ��Ԋ޺�f�sN.ӣg-XvksF��S:<�]R${-��2Q��5�zp����*,m��SY`�ĬQ�A�`��1�Y��l��<x��ϧ�?_���ffg�3<fs���|s��՟��=e��!Yovc�H�JŞW�l�y嗞<z���||fs339���L��Ϗ�9�Ͽϕ�)>��Q [[U��#-
�q�����,�c��������3�������ffz�s��Ϗ_��,�����N��RE��j�<�O��Ϸ�����333陙���Y�|}9����J�e���|�HW��Ѕ*�|���QZ���C2��6�
�)F
��E��1UZ�XVhM�("(�US�b�㈰F"M��*EUPS�(�J��F1�Z�O5b�Z���0�$R�A�Օ8Ց`�[7��WP�������UEg��DPQ\K�q���s:����J^j�eL��딗KL�e���8RY����C��5�� ����n��ﾞ��˙�����d�%�3&K0�z<���`�%�Ov���S�>��Bڀ`^Vߔt� ����}��O8����"�"�8�t�T�%�2Oa����~U���?|��q=W�Py&?�� ��H�l� �{�@�|��5�c7R95u���fn�g���N�2�IT)9�dc&�v2����s:qqކ`h\�X�֝��x��2:^}7����O����OwW5����i��zo��~�[l�C�����}}��ק�Th�ce�S�?g�"#�h��梼�ޞ���Pc"���0v��Yv���D�LO<�n��[���-�`��	>��z����_}"��Σ���an�m��[�D����P���r�՞�!^�5������}5W�{�d?�h^
��<�?7k���~e�[���}]�[Ϟ=�����Zk��s.��3��3&&"fDo��Q��\�,�a�^qyW��,./4��4�[Jm��w�ݛ����b24�SՔ����|��?�<���U��o8�!���N�N�]��g�U�
�0.�����7��2�	V������w�s�ą�yGˆ�@��Όܵ/fn���?gK5st�kJ�,m���u�7���<��R�mb�ӹ`��������>~~^a��?�7����{�m�7Ov����q�x��y�ߗ8�\,��
G��,����0(2����/��3�����X~K���]J|g;�-�����Bɛ�㤙�h�w>%�9�Qh�ff�Q꧗��õ-IP�"]��>�s��Z�o�B�S�
���q������\ry��c�#��e���5݋x��vp ������[봊k�vߴN�R��O�����?�n������m�ɸ�]���H�~�(��);�����:C�V�'O�{�s���� �i��
����ҽR���k�N��&{��.����y��9�;�eU4�ٻ�D��wt����!��j�
L��R�S�_ND�:z��w;�2�:$[�`�;z(	���ǻ,a=>Fzk�K�@�|���aś�>^uhff˞ԣ� e������U�w򟳳������:�Į[�vZ���3�Ug3'g����)L���?5*�e�1����V6f3��$/n�:��s�ψ���fZ
�ɮEO�����a�*�&Qc`Ŵ�����(֣	o|����'�Ie��Yec,�.�?^]���?���o\Q��]4��7��@��K0���UKQu]�|��\K��X�t2�]v��M��IW����5I��}>���l�?f}����|r<�ܟ��a퍸Ց7<�F�Xq-�9����y%�e~&��?M^T�������x�d�X��[:�;ka�}9w����:�HQ1,����zR�5��z�!���q��/y�j�,�h��{��xʹ�i�ݻ�#��y*���̿v�#��>�nΉ̆�&���q�[;�|��0��x��!¹�:�π�9�ӕ�G�	&Y��W��y���V�p����93��9�`��/��b��C�\A]����;�A���1?��ꋖ@���\<u*��6�y��D�0S{��uOy�g�-����<XL����^������7���"�X���pg�5;�=�l�L3�@`�y��l~��RD���XnS�C=��y�9|��ZP{F��Kм��;n-wzu5��ԌR�����w�/ky�I�¸����׸�8[���&m6��
�Ȧ���8��hN66m���泉�XWM�{3t��3���_]�S�ŕ���p��(�Dπ.�C����G��R];!�:��WU����2�=3;��{<��������yy�������o%}�=/��7���3�#��>-�����������)ţ��J���b����&���unj��K��\uÞ����º�[�Z�����m���o�8�����㗛��\X��TTS��g�;�O��H������":��k7��_l�zyOw*����V��p���Z�W+�v�-)�N5�gs6��{H����\����ِɜm8�*�ڝ��V_�2gv�����zx�$zY9�tu�Kao>�3���"D�1&��Sm���n�m���;�X@�"/Ž��Fv��KwB���a��TQ=��׍i�7�?���zyߚ�qv�6ri���ᡛi��)�r������J�7���'#�1��]��א\:�/�X�4�%�O����P7[��4י�ǃ�V���o��y	̑o�f��^�P��,kVݚ�<�MPQ��x}��]�Aؖ������'hz9Ѿ�Y�R�
�|�-�n[��P��c�ھkx����>�af9�г)YjH-h�|����V��N�?�d�Ie��Yf���.��}�����ޫwv�2�~�q���a$��d_g�����ɵرn*z-��f��#jlCC�k���|`1�j��oh�?�C��!�׹z�����?��q1/�M�#�-Q�w5	��3(�F�z:�����ITlD�T�bv`ԙ�.d�����z������fs���[���P�磱�tϞ��n�������|Ξw�o
������V�F���ѷN9�aP(A�����1g�k���$����@�q��<nLy4�G2u�Q~�g� xM*ۃ�A�+l������ ���p-�e�{�swpT�q�GP_@��z�T{���'�G�6�Ļ�Lz��ZW�23���b��x@TX6��˸�>��A�]�`��36��u��g�����^,�1�:��Bͦ��w�����>�(�E�vkF���+�u��B<D]��].�H<��]󠣤��o`��K�e�����?.�Єi*'�����e'�$����v�a�^��7qԼ�9�&����_uX�8޸k�[=�汷?O���YIe�,ɞC6^�iKw�ߪ+���Ty���d;8k�# :~[�F"z�DYzNI�o����nŉi�{��=�e�{K���a��e���w ��o,��T���Wh�� \��gg�u>��T�fǺ��+�`׵�|��7�ˌ�(���bU�;X�΢}o�ʥK�����{�����yӓ�������{��f��L�-�p2��t���7d�U_��}k�M�bVK��Ƃp;';b\tR���]9�s�]��z^A�S�^�?������j]���G�ݷ>���Z�fo���.���"j�j�b�VD's�,�z}^�W/7��)���MEC+$����ݔp�Ӟ���{+�}�l3X1)/O���.&VA�L���	��ӻڨFvw������J�O�m+��g�W绑oU�ѓ�U��@6a}ffڬ!�od�� 웚xM��8\ta�l�D�u_��i�az����<�*K�Ty+{��O��>� ?j��W]�k1oL6��,Ri�]K�����W�XOT��7P�M���e�ʸ ���{��h�xC��rk2:������,��%�c,�}�u�p���5'[_�=�2Ԗ�I]O�%Ŏ4V�f+�Hc"T�kXs�;�s�]\u2vb�0XyY�l��m��a����Y����T&�=�G���L�O����b x���C������w�]Ƙ���>EM?��=��H���*�ee`zmV��w*��U2�}�C.���9N����f�~�׌��o�Q�5��z�o3vI8oxn�׭x5S��Ѓ�>��܎�o9q�����X��b$<4LH�3[t�m6 ���
�p�?�c������@��v���`�wף��	�x(�@��έ��jZ�ZA�~�t8�w�m�1r��C�-�y�&	���WtƘ�饳�M[׹BD�8��wg{�a����m�(�;y��Jִ0��;.���=��wvݕ�>*`<v�r
ݍ��I�3Y���f��O� I�O3�}L:aV�_,N��b2b�S����\Y��ށHP3/��g2W�@����a��}�0��t�*杂Ϥ��[��ٌ���ԙ�4胷X*b�ӿ�B����i�K���|�ty��iZ�|�q������F�'�{=7�,�N��BC�E�2nK��\�F\R˸�����|� 0��#ͷ@��`��ǃ��7-����<�����������No�[ٕ-���A�s�^KW`��P����K��{�f�
ׄ�N�ĵ١��B��=�x �A�^�䬟|W��Wf5ܹ��e&�N�ݼ�km%��+���	����y�A~���g1�M����'7V��z�f���`E���6	�՗�'���Z{7���ٛ�0�Ⳝm[������K.8	���4��	�7���׉7k]L��:w9iݲ}v�ոA�W6��o���"���]�T�h�	a�a�;0c���ZFV}1�l�i���;�꯻2{��{ж�q����Xp�M�쑖�ar�t��a���ؒ��W���S̨�_z*��u˵�xQ���v�uqR/!+	���k��r�Z�Hg��m?n�u�ڞ;Z{��-�W2��[� ��k��֑��}�e��	MM�3�oJ��d�ԛ�P��4˪B�w}lD%���w([0d�*���s\<v�Ў"��F6��js�g=�������e�n.5�qg�����"B%�����{�����|���̔�YIe�ɒ��������I�%�#p��K��Z6А��o}�~G�C��v����[���n@1W�qc�9��~�	�?9�����w� ��}�����':b�����nU��L�Hc!���;�5�:�zv1�Ov��=t<�3��$��@ZmW=������7�1�,9��?q����m��u�5��Y����=:��B����6g��v&��ϞaҒ��#�}�LJ�-���+�@a�캊�;�������ntA�,�zoD�d���<[��C�9A����Sr�i��G��0�6s����Mέ+;Q��|	�
p����LE4y����0恄@=70ї
:Σ���F���5�Q��}�A��,�M3���'����9����s.�S���������tÝ��8e0அ� G��.�&����v⧙��٨�rERM������0w_�\��",�=w�U��_�x�p�O��� ���N��D^��by��:b�T�$�cd&U余��
q�b��j�@&�n����{�P��}����z<�������>~~^~�]^oӾ��A���=�}X?��[w#U�KS�K���NV�N�>�U�0k�	��@峜p�t�wT ��z6}ut�|���*��9�l=�L�%@��2��0������"A�k͒���|�64�8J�h�˅T2��Ͳ��ne�%�����)����+���Vy7�p?�������jv�u���f�5ڛ΅��B�q�6��v���*�u7YEnaE�eS�\�"��������x?ux�0��S�6�:n�fVa*�f��x�h���D�݁7�����͑���(��f��9wf_^̊co8�m��y�V��Q_{�� �`o����{���z����c��-=S<׍�S�fp��Z(L����\*=�����v��y4W��j
us���.5����,F���f�g'�9�}��V�O����׈�=0YmL��\\SU���R��:1!ɺ:y)�ab�w#��P_='�y��g���mꮜӫ0勷��In�m9Ž��`����ҥ�̚�*Y�z��L^�p� ��̷�pv�S���OQҍf0����v�ud��D�"����OQ�娖�X8����aG�S�:��wM嚚]q.[�4o{�y�͎�K[�7g��p�2P%��e�QN�����0�on� gv�ƛ[���zsky��++˅�f���U�`p}eԲ��:�n�A�I�7^����q_Q����&j'��w6{7+^ e�;�X���4���6�� ����o9�޾�;��AuŒzUպ�Ӓ�NW��Z�2]Ґ:���]K�-��v1��k�T���$���["e�D�u���e��tu+�3�I:����*ɥtA�鳸�����)[!:Z�Wx�4�LZzVgo5-��o ��v#�p����DZ��]��Bf*��g"�(g^O_=F�.�Q�Ů��`�o����ht���F�f#��@˭�F�\@|p�_G�Nu[H��źH\/W^�o$��AK���E��BһDB/�^#I�yD&�gi`��M_3�؃��`a���Sy(�2���jG����Q2��V͇X�d�b�*��?e��ɴ�B~�m+J�� T��*��2��PyN9�/2����5nL���b�9A�a��ƫ{w�ɺ��\Be��^���;������Pq3��j��R;�%�,R����۷�5���ծI8eY�N���W[-�=��9�l�[�K�vE�LJ�[y��62�SՕ%��j�{�}x�ǰ�;2\&�f��S���J�a*�rv���ܣ�7F�Jw��"����x������V'F7�����e䆵�6&b�6�x�r�kf7�pk:��s9yD�h�۪�-0m�Y�)p�p��؅ݰ�q�P+��-��0/�f%_*�I�#�ז1g�%*��mQ�({/�B�{v��"��3�M1�C	�;&�Q��+�fef�]HD��<۽f*ڊ��D��(�eb������z����`�r͂�Ŷ"�Vc|�u�齯PF�zZ��[��s�1
5��a4�;|��t����t�"P�o��kl�"p��T��$��,ح�2��3�U�N�+�)�3t^wVH󦧼�]��ؙ����*�ʞT8�V��1�V�{Ԝ�MoDw����ә���U�**�yQ
D�F���w|y��׼<qF
.��b�a�հƠ�חq�����϶~��ffg�33������75>�<�z�d��5ի��jʲ�%�wǏ^�>>>���33>���������ӟ����G��AI��X_�X�ʫ>ݙb��2�W%�d��}9>3=fff}339���9�}5>�y��+��UwJ���K��'���Ϗ������33>��������>9������'�Xǯ��کհf�AF/�<��F(�aR-�X����D�ۧ]��c���j�0�

"���E�-FE-)����V���&�b����!h�, Q�R
*""�DXi�7���v���(
�4�P�bȈV��M5FAA��`w�ɶM�H �����I��./D�.�)$&y�L�$JI h�c��j"�AA�$!��X��L�Q(y)���E*R"ϑ,�HA/H�jF$�,��k��g4���F��f�Qt&m�7,�&��us_���T=+x��)6.<�[fԬ��CK�(�m�"�D��P�<`IFDE�i4Z2H`A���pC�i�T@�
%��
��1⃐! !��m8\F9'�B�)�*�U扇�0ؑ��e!I�P>�'L=@��#K�4�X��$ӄ��	��0Sb2	Q(�L���b(g�f�9Q2��3H@�N���E�Nc��<���x�=�^�{^�x�W�^=O�ο+��_��֎?�)jF�'L��ov�l�*V�.=�Ȱ_	���4��2b4����3��(Uk�-������P��U8�T�0�׷��=��?�,ϲ'�Њ�o+O�6��T��"�.ӱ��k�%� {v�������</��"�<Tbs��{��X�����ѽn�b��
�FA��&�3K.6�gFt��[�n�Ë_+�F�D�#4#w��\ܶ=Q=�i<�S���n�,k\��M�o�Ri������7��y\�ٚ+<!q
�>���+U�Xه�s+{i,�t�ٞ��{��=�S��R��vYM&�D'�@������Ipu�0�@=gN_�Ԝ�-q���ϱ��}MǮ����M����(��{z�Lz}Ƽ��Pw��N��5��K���V��D�nS�ϸ�bN#	w�g�邟�g3i�{��߷TYw�����F4EhP�h�~�G��P�B1���8gerU����faU�}������?V�ͩF�;��4s[8����n1va��{�]��t�Rzl辵�����|p�����w0��� 2�����T~����Z����][;o�U䃓���dt5�V�[Α��œ�N���	��;,�d�f2d���0�����~��oO�����2v��S gb���J�y^ǌ�Ь��fjT���v`vaC�{}Π��!��0gY�B��l묗v���_.�|��g<���� j(Ͽ|}�y�ym�Fϩ7�� �cB��`��j�٢oN��T��#oˤ�{���0��p�2��`.�W�+j�H�|���r���ͦI�F��c�
����|�ZU�ܬ\a��F�S�9�Z�Vv�0���������8�����G#sy�sZ��I����*~�f~����+� �/Ls���}a/,�2$�m�0� k�#v���!�ĮQ�3`������M~4֣�]�𩧟Y�����^<��u�M0�;�6x!��Pof���i��9��f�½�m����dz�5���X<geu[�ge�&��OZ�O�}J�m]�]d/	�U���Њ��e�f��մJbVeY�sE��g�GЬ��x�w1���P�^vO�aޛv��.�@��|P�\��a����ʻ����`3&K0fL��Yfg�{�����6q�^ffDϜ~4�V���*R���2	�/F��@ɾW>��3��e�fLcK3���픖������|*x�s�%����
��W2\���hGU%P9��8���̟��*[f9�.�&̲b�܈���7v�s�_��-؎f�j��ƃ{yf﫳�Q�5Y�-��Zl��gl��1�M��l�H�˿~}��{�-�������c�NI�Q��t=Vk<T:���[�Gh���{�8	N�q�-1��G �*|�vDo���Nҩ�h�7Wٙ���Z�*x���WH�҂�@"�_�1�ni�x��[:��즫&����U��oy�!c�ҝ��/�1w�ެ&謻T�LJݗ����*C���ʁ��}V�����÷w4��`}pޗ���3�Է/8�܅�4�4��kqR`Z$����_�nYWiG[:y��;[��z��X�R��l��xG[�1P�9{���hT�o9f�+���@�[AkߞT�W����2�>�o�~�&T�Y�ڻ\vKv�kV��,���]�/�[�!R�L��𑯮o
����0fL��YIe�w���w���y�c��;���Ϩ׺��[�[f&�f��/F�xn�zX��n@/a�
��t ��`��E�1��Q�pt6��ŇTx-�>W���m)L�e�PW��=�fn��`�;�}�q���5���\H�Gg����Y ^��N���2v�\�y�T���u	�ܘ緍ɮĭ^3mz��V�`a|}Ҹ�^Rpi+�	[��K�h
��F�umbTt�t&<��B�z������G��q��g,�cs���G�w��=9�p��o:��'
�x�Ly�E�Uǫʼ<9J�a�z4F[X��¨)j���}|�{���h"�S�~�q�v|�=N0FOND�j�8_6i����d�����[�ǲ4��k�9������,��<���=��O�g@Ö?r#<��ܥ7��O����9�t�R�A�gd=���-��#�fv��ٹw���N��3r�Y��v���q||/q��$5z�V���&;ݾA޴8L�t�M�$p}$�b�8�I�z3��;���9����wɱ?MM�K,���K,��6|�4Q+�o/v�fV9��5a
�O\�H�����\�*J�޶�i�В͚LNSK����
׳���){�A��Mͪ��Zzq,��@˄����^Ү������9���v��������Zo۵P[J�2����pQr�@��s1�����8q �\��A�����_tS �FG���&�yߍueYZv�
������=L�ʯ�1}��+���~]�{���k0�s��x�h���t-��->�������]O7�=�Ӎ�����"���*��wO�f��aU���S����(��L�t_oCh�"�*h�a��\zy�AӲ4f�!@��T�O��゚�ݡ}�Y�h��#��}Q�P0�Ҭnѐv��������^���N]ٺ\(-�;��z}֪}����4��uj�ԒX¯x���y�2�M<�<y��:G�}�܃�8�P/Q�q��#� ���cE$��H~�&�����8{�nuo#z�X�9�NK�&��uP�������#�}�u������s��y����HD.)BH�k�c �2��V�P���}�h'ً5é�^��#����?�y��q����13�������{�M�ٴ��"�+���~(X��>S��X�wl�&��@!�}+W��I���Z�G�-��p�l���hv���,��#���E6��p��=˄k�ҿ*xY��|��er�,5�p,����t{Ξ'v������C�$�`��M�s���ݾ�w%>�.��73��v��l\��07Sq��R��5��o���0g��榨wi��q��z���K��~�w�v�%A���a��{��2ө�47*�/�ѭ[�^C>sp��ϕ	�*����=|)����8��Zmv���S]�����nCG��i�A���`�H�z�'�Gv�Ɖ7��7N����^1��;�hi�,�"���1OO��¦Z�/	KW�����|ق����V�g�1�f�y� ��Zbj;!��;��6�̙�SG��0��N쵁�G�]���R��zwvoE����7z���i�@�k�&�Y�Ư�5��\^X� 8� ��_]��<��;�l�Lq�A�F,�����<�8��������JY��P�Z�2�Yى|�)���/��/�!C�8��=Ǯ)�i��Xs�ёá��\ 2	���j*7�j�Q��ہ�%��#�Bȥ�v��wl�åO���X�c��¨r��PC�el�̻�X����N���Vϓ<rؙ4�}L|���&�q����*�����oV�v�"iݞ�)yO�{6�� M��F��Q�q:�x�E�
�!�m4s�VxD�o{o#zE�p�:���fd�݂�K�6󺃚�1��Yz�C�f��ҕ���:�w�%di�>�v,k�{�3{�3c�㵧�{����^�n�0ga�Q��1��R6{:��&2�^�ff���^@��Sm�X������J�u�D�����ȵ;[�8�n�ޛv�)��J�^��.���w��Z��34�;
vܰ:5�WX�*��"ۺ�t=��|iocLU�f�2%J�]�S��g9l�e�zĶ�r��c�np��66��{l����x��n��JS})����Jҳ��39� ӫ�5����K�D�\�b;:�>w�_����w��rYIe��YIe�>��;�mz��e\ށ�����̥�:��k�x!s.�\j�u�ԭ屉T�1�>kKz��v+|�==a@^�P�5���􈪪�2��]�\0�O�@ہ]u�1�;���|�	8��g�-[�=��чx��� �Fg�\B#���xk6ǲ��I&e�q>����޸O���s��������M���/�o�׏{)�p�y7��či�a�4{*��e�!�ޫ�����{w��,T�߷�j��EȒ���)��1���^N/n��zϟЈ�g�����q�Z�>UC�L\q�ZQ��.��������>���Ü2
}6D�\��=z�',%��J*�]������v���~��yf��Dh���P}�_n�\�d�q�����MG'�^� �7O����~��v�P
#��}\�vV�+�I�����-Y]\��J���ּ�h� �n��Dw�mR�C��ǖ씔��M	:ZB(�}X�'���C��agt��ޚ��;��Ѭ�H��vuA��~�!���<���������Z9���L:�ݱ>�FT[��`�vf�[�vh��sm��k'b��58l��E��r�j�B�r{�C��u�H�֋��l(	:�n������C@��ffj>��&1Uq�5�9�;WO&$?EV�Q+�^p�6c��x���[vP}�Ӝ��ϧrݍ>D�b��l303���ҹ�ǖs����ύn~/~~ƍP\5��5��f� �:�oZ�Ws{��n����������ç���[��u�*�Q�S9I�X���ؿgt	��F��V^ǥ��8����u]x� k{޺���䵻���f0�������2�H��c�9Md�Jp���q����}�R�$���/�A�XQ1�۲xRO0:�a�Z�`?���4�����WO��y�|���6s;L�VA��^8�g�ײ�з��x\�\��f.�ջ[�x��&��x�1��H�
���ӜA�)Y�Ζ����6\�!���2��z�%���w�v��s�N�t�"A�V����3�q���l�Ī�k�3^���������qT���]H��g`�;��,��K�|�ۯ5���/�̔�YIe�,�ڪ��Vn�0Κ雧�쑙�!�ߐ$�:n_�kS�}m�[�����S���w�U�ݛ���9���2��מ�\�4�ْ�6�SA⦧Š�?��"�wW��z�]YZ�:��c���^�WW'r������,���C�Lz��|��P�4���i xYO��skdC�4�<Z�Y볫ՉK������n7p*�r�h��1�=r!dQ��Ê�R��r	%-����9�qù��l�*�ON3�4�f���(���;;��Ι\K���Of�=�k{���-�fQ�Y�r�%I,h_:~䦹U�����t��d�?O_�|�<z�
�ި�5����,�G��X�2���T�v)�ټ��w0$��Εy�sNY.�Z��㏶��0���v�J�f�vcl�mBOW�u�^ðZ��������b�6s�+��� ܰ��[�y���Gln��5��v; Ǉ�����PngnD�潩���Й�w)D��n^s���7����w�ۋ���[Stv�+�}.��U��+��H��k^V��|�iZַe��UT=�:od]�e�}}�Yíthn�8��A���]p$R��6��k�f�Y��W�Q2E%��K�IJ������v�C#���\~C�����}��^�n`�yK9D�u��u�V��~��X0T���B���̴hnA�op� \B�Hr����\l9�Ĩkk�t�9d���|:��Zm����{���S��A'Z���EYJ�����Y�yw|�&��ԗ1�D�.%���I�V��Y����X��W��OF�{I�>6�ֱ�&a��x��t��J��QԴoQvq��1�4��CkB(և�ATֹkY�va9�)�57W�fQ�pH���N�@�i��%�[Z/�p�˃��X��zs1��C�ə�y�s���7/�$��i5�K�'Y��N*����hU��,�|O����l�c�#r�r�7B�u.-a�O]"|��(�t������S�HH������n��\�l�(tH�s`�ʿ�#<�|���2S�J�؁Ɍ
63
F��-���O(Q0��7`Sf����a�O��O�o��}Q�u���9d!���08���97�iT8DU��������XHfefmY�(�O�^�Mm[�q��fsh|�2�R�읚k�x���N�͊��Y+��U�ˋ�g��DmH����^PÊa��\�n.�k���.�˔r�`�R�{7#-��wp��܁]-����W��G�+X����(+[aWc�35^�Pb��zT�4������z�y��%[�Vlf�/m\�:��Ѭ�adʬ�����5��1ؾS4�UwK%L��ͭ]n�(�����#�r݅�X؞8X�u��j% K�����K����Q�b鋲�%�C�kX!���B&G#ԏU��R��m�>��n�*c!��{�,FlW&-���+���z��\j"S����ռh�g5��B�8%gH�ĩ7���>	^m�Tc�G����ݖ� �Su�Ɉ־��A�1R wXZX��8��5H��K�vp+vb�Yw��!R�aV�b�K�Lޒ0�"8�;�ɗ.����/\��r�{9��Lߟ�4�=J(q̲-B��
�eL�Y�#*�ɩ�������������Y��Κ��Mϥ���,���C-hc'���{��W�=�������x���϶fz���s���|x���`�<�b����jJ��*ʶy|��ǯ�����||x���϶fz���s����~~[m��,�؉��i`�a�i�M�23׬Ϸ����񙙙�l������9Ϗ����?|y?|���l�_U~�`|��UR��a��,�"2��U`�]�,`�4b�j�(�R
�Ae�!�EbAm�UkF1QI�����T�9�b��8
��q�S�Y�R"�
�$\J�Z3n��P*�AH�#Z�TkX�2���icOYʸz��΃�T#��@wv�R�M��8�N�"#s�ލ��:�O���~���ɒ�e��YIe�}��Kb/^!��jɵ��l�0vL"8b3��:�N���b2aM����m�K7i�\�fi$��J��
�<>�����a�D�̭���:��p��y�
���z��;���M\2��TtC5�nǬVO�L��Sb�KWl�1myQ�tD�˖`�6�����^���j�.��ÿWp}�S��ߦ�����x��������L�u�{z�1��CP<�ƪ��1���7�J�7���7�����n���y}~��O���� ��9C����*��b��1�����Cq�)�����:n�e�ߥ��S��̖_WDK���V^��7f%�fffbyu��Hz���&੔n�ƙD����F�|��2��I�RV�R�T�\��dzήM�씒�w ���_�EU��6�~!J�U�jۡ�#eK�v1��x�����*�s�.���)�g�<����z�e������s����yg2�FweLZ'����_Q�o�qj0��/A�W'�=�����]k*��}�:0��g����%�Y,���7�<׾�����e@�����6 �p�wPӦ[g�.ة�����6��h�d ��=t�^���oMg�ڪ�+�eѠ�bazs�.n߮��D��3�#5����ߗnȽm�5��Ƥ��x��}����ʙ.�9��:c|����AK>[?�7�=�|s��zY�I��Yt��w&�#GF�op�����4��%�<5� B�.�3�w��\}=�i�3"��v�� h����̪�5r�Q���v��||�C��������|��j� �]���21W��+���; W-��u���\��}"&�mVoa7~��-�ֻ=#��ի���a�n��#�:��Y۝xy>�L���!,��Y����wV˯>�"�.��T�2ޢ9�p���Ks�p,�7m��a�E�0���\�]'LѸ�nW`�M��T��R�����/�.�=�_l3 �'��]��x�ܘ2�����,���P�A-X�{�F6��u9ȯN�aY��@�Ô�glW�-IM�����uFvY,���),��>�}��g������?nX�w�M=g���@�KU��
:|�g.�-ÎY�2Ѧx����Ee=�^%�"g^&m��� 7y�@(>l�P%@��e��eS0V9G����b�].�Ý��I&���~�^�3o�}];j�]��}�JIƆ�j�*�Q+�W�����qz6.�`:�r����{�z�mۢ��՝Oñ�A�B�2!(������a[���^(Dxx�W:;ح�Sl<<ü8ΝP
Ϫ��E3z=i�{��x�SL8�Wv�O)J�l�D�{"����ƻ�oe��8�o;~Ɲ�*.fZ�deV���t+U���&��0rUf�ѳ�RF��sB�C10}:�Ur�Kuj�F�v�l��}X��&G:1m����+��Ȏؠ�a|]sw��������R▙���'�U��ؙ���qJy�د3���m�����ĉ���ڕ�1#�W�������2-ވκɕ���kM�a㟲�}.w1pW�>
k�5���X���vYMBp*������yr�&�U/�ai*ܹ�K=`Vi���5bd��+D�=�ˡ�u��g������RYe%�RY|�^ۣ����/�y�0]����2�9�ܧ~����p��9�͆�vh	\�W��jU+Ԭai�`��{Qk}��6vd�@�X�*[.�w	S�/"EK35�1���(��Ќ+����"%wz�zT�X%��nJ(���W�j�[�X��4;��}��,�����yfۺYz�N�;�m~lU��Lz���w�����x�Bx{�jU�Y��qg&dpy� ���r�l���^B,��S��+��zj3���v���j~/zЫ�=�QZsC�,�f�W�y�E8��wz���+�ub��`�L�����u�ct�6�Ta��{����x��_�g�����y��[Rs/o����z��K����3nq�nWp)a�Ɉ�S75Ik�J�l�s���}$�}߳7 �I#��+͔�cg���t����K���<L�|{uv�ou�p����.�MhMK�k�q�*�I����SR
v��gGZ�]������u�C�$ܫ4��AD�M���b�W��e_���/eg�3�g=��{���䤲�%�RYe�����d�r�͸�q�Oy.כ�g��{TX`�Ά�5L݇b`�j.����s|�2��k�M��|wkg�qn��uі���7�&���v�axn<��:�����8f{Ū�o�����ǫ���,�3��V���;�N�H�g9^�`�ЦmI��}Y�Qg#cb3{��%��8o����g��3�K}8�����<3!�][��Y�V�	d5���7r5"}!��0�!�}�q͞�Ù��x�g{2)@J(S������N�%>H�y����w���xxR6���v��)ƌ@��x��/L�b��i����h*��Ȇ��"�ʳVVa�H�g�5n��s:��u�蚕W<�(d��gR��a�r޹f�}պ�������@��]�,'�j*}���twk����im�����wM��}V�a�bl�x�:��Q��r�>��ڥz-���K�T�ݳ*�}�;Q*�q����<0�w��-w�6���f\�]$����`��r��u�<�X~�v�w��Vs(�q����2YIe��YIe�5���{��w�|3�y�$�_\�`���Y��9@~�^���]�Pz/�ƒ����u�q3���-���o3�uV8*����3��b�[�j����3�z��G�e�Evx�����bJ���P[��5�|��T�=���IRJ#�ur��"t�����IM�����eem������@�qN�y��}�!��5x4�o�U�s.�����x�.p�Z}���h�չM�柇;!�Ɏ�
���]���9����EY����&�Aop�{K�#07�\��>�!�;��Uy�|w�r���������[��ޟQ �	f֧�܏X�=�i�N2�c9������Q
<�ł�P�;��I�Jyo�\Tq�R3{k��#Ez����o�. ��h�r�@@{��Y���_Zgsv�G�+�(���B��/�$^�]CD\ѩcL��
|�h�V����z�<Yy5I�����(�0�"p�JH�ϼ�c^����XF�����ne�f:"qe���nr����MK�y̹u�cҧ̤�D1jb�hB�(�un~�NJK,���K,��������}[�oc�h�����1�mIdJ�J��|�]b繑<:�\s#Ցdгt=�k�N��a{�J\�6�wv����Ԃ��r�@�F�%� X&�Of���:��ox��d�v��F�Q�	sH�u&}Sh���.�����K1a�0���8:=����p�|틝�33[��l���2�����jq��$��j$���ݷ:{̓^G
v���*�]1�w͹���B��&�G��q{��}&�ҍT�22�6�Ua?�����"{v9h�����򓓊�E�W�V>:5��n[�*Y�O����~����QX��O�LY��__�3����{$�����ρ��g	Ywx���i�p.����X�~�vO�Ȥ�Y��,����f��Vf4L�rop����XL
]���	|R�=�6/E]��9�Z�Ţ�a+�4ߩPJ�9��o/��~��O��9��T_�����_1!�wt��w��u�%rU5F�M׻��^�K]nBM'W�l{�d@��wQ`)m������|	GH�4��au����Kn���eQ�ˏʣr��=��yL���e��&��;���Vog']�yc����yyy?���?���U^*+o�x�rY�9��΃��#������o��{��hE�kR7	pw:�F���b=+3hY��?w��� O���q�KcvM�>������/RZ�<�D�L�T�S����ϱvi?�ӽ���5ѳn��"w>r�,}~@W��30�����}�){�׾��[��Y��A�w8�_���2�+�Vx������s�f�$���}}�\��nմ=]Fg%��3{�K�yyhxPd(�xy0�`/�@LGK>ҨK�������ow���¯e#KF��w��x%Q��0$�p&.Y�/��t
P��7��[L�T��s] �,�}.4H�^b�z�K���V_�fM��̾�*�����g@z��Q��}M��w�����o{V�mcM��Յ+W�c��y�m�橎�lץ_z�(��B3LU����w���G�/g���ܕ��m��͚n&�GQ\٘��f��;���WVYM���!#/�-��馏[z����˙�v�N�*搙�k\6Μ��H�U����cgC�c���Y����+�;�z���˭_�vrP,���),�����sU���e�<C;����ϲ%�y�!U��;��W)�z�G<>@��1�D���Ś��=A,K��p�M�ZR�"�;{j&��d՞�[Ηtz��-�]<C�1U�����~�u1���^i7�^��
im����*Q�Rhm���N��^�N�]e^\.��w�U\����5�)@r+�2���٢��7j�)�23]���=��`��?$�����,t�c��v�s�5�O/ks/wqY���5����]�@�����iڴzE�
U���8�D�0�mc�F�wf��=��3������T����KF�@g�]�Y~�_'���#+j���q&o8C8J��r�e$tF%]�{��N:�n�ǒ2Z6���gzwaS��!Jg��8t��;�Uߞ�����۷r���ǂ�'x�}v��Z{��٨ZTe�cʕ������������`-�V����Id$p����U�ZYXƓ�`7y���2p���{����JK,���K,��{����ﱙ��F�����M�\^��o@���G���,s6��oQ2��S�Y
��S�a��-�R�v��>�ZC{c�JfhxY5ǖP2���T��E��	^���x�[	���vt��a���N�fם��3Cv�Б�%��-��#�j��{��v�n��������9`e���B�c��1y�l�M�Y�4�7�ܣ�3F���>'�����#�>��٠�}�k�'ϩ>O��!�^�����$w�����-��F�]�j��Bl��'D2�Y����Z!���zj����Hu���ܰ��ń	�Gc/kʏ/_P���#�j���6V�X���׳^D�x9�"{:�{�N����9�]Y�j�,;�sL�dsP�~�\��G�=��P������ʲ�Tf�������9.�%�G��Y�;��}�LS�&�[Y����7�7����/MMV���ލQک����S��!I �}���[�·��.e�k��$��j*,�ŧ��>��_E�)�:�]G[8���k[ϙ�\�`���Y���a��e5��t��]ۄ�H6m��]�h�I�����3uNwu�m�r�����ʮM�ʡqg&��Q^oa�Z��Rۭ��`�r\
�r�K1�UfUAʶ^�ibOw��H�;�jMi%gz������Z�s7�I��͵ԍ3����r<6�3���)�W*��:)�ܣ��GzQ��d��ʻ
��$u���{6�[o31�3B��2X��+�}�*5+Z�3�tCF�Gm䃖Ѭ�bx�M��3��IY��gV����gtM�=�S6[{I��Yc�42fc�[kJKޱ ��uVt��v�ee�b�n�ѴϞ��P�!���Czr���Ηe�O�;�:���7�������v��5X`=(�&����8V��l�]���ӯcV��M�X��K�pE�#Odʺ���<}B�^ܴ�#+6"���t:�R7m�R�HS0�:�6��|3�\l�7�Vr{!q#c���tU
&��Q�U�!o�ɷ1�8��K*��W��.6g�U>^lNL��l!��CU�3b�'�1a�E�3]51�����Lˬ!�n@ВESoJG�($��wV�^Z�����&5�_�if�v-��v#�1��8	w[��<��;{,naA�[{ݼ�2,��V�L�X7a��x���w��3,]��������I�u��9������F���~ޫդL��lP^ߓ�]kT�D1}tJ��(aۋ9<ZV늝��67����\����=�Kv��$40��7�Ur�̲��,XB��2�R��vt��8��9O�ڃ:�0Q�xe�%�o.#[�ĭi����}}�Egx���ہ��;W(���R�C&�5U:��2T��\"QX<,���l^ʜ���\:�F���Q,Ԅ�3��i�R�U� �:&zb��r�[��a)λ[��DhB�wݮ1���HČ���mp�CӦT���;�uP�ǉt�኶�_t+:_��!�.h`}Jnm�0�'��Ed\9�����UHs�v��Uvq1r�e��]צ��m1������_6�v&����=Rjp��z.R�v��&�e��E�d��\��Bm�������*�JHI��]K�1�!���R�JZ�ʱ�j��x�I 29�@�ȪDUDbu(��cP�O,�y��>>>>3��������񙙜�9������j�?,�G�&ZA�h|��M2Y�-y,~��^߿'�U�������~��333?�333��9��_�=��(5���(��e�j[-����Ǭ�Ϗ�Vfffg�3�ffs��>>+��[)TQU`��J�L���[��m_�x��������������g����9�g����?+��$��*�V��SwL�Ptն
�qf\E�*,��R�7�#Q�J[
�*bm2�TJ���QQ|Ja4%dF,uLC}s˷1@b���j����13�c1m�3YLU��>ʃ�)TM9��dP�X�Tkj+�L�����Y-��
BHp@�	�P"\i@[@�FÈ�g�A��H9�l4`�B)� �L�(�Q�Q�2 Rx�AĂ~�$��TD��BD��@�M2U����{�"ͥ%)P&ҳ3��ܡjYr���;�ȇh�I��r=d{¯����L�ey�Q,F���!��!�	�"`�M�iFC�L0R�b!"E��."�y�B�AB��i�Q��FH�B8Ӏ�B)�H�MD�B6ȅ��o�HZf13Ģ�m��l�Iby��e8H��2�� Č�1��2d$�B��I�24T"��$�qԨ)��	S �L���A�����YIe�K,�����m�G���o�tI�q���X�D�QB��u�4)�:m�c7�K��n�Za��w|p�
K�;]	�(��+��N��qd����p�=�?��O]u�eG>��&|�|`����O��.�η�@��4w���Nu7��Rܐ������q�a����]�|o:n:yJDF����w��Z�������Z�ous�Rٝ�)v��N(n��\
���7z�H�7sA��(\98�skI�k$��̻���y�>g��=H����d	Q��U�^ȸ>j��(j�"���\sV��^��^�~��7�:�o���2��|���L�V<J�ڱ����L�ʞ���;p���V�x��k�7'`����6oUf��n�z�����@� ځ�O��5��b~g��;W}/7�t��֏�aċ(C�;�w\��SI� !��(%m�z����Fn�h��5�Qzow�������2;�c��`\����׮�j:�;.��-��ې)�mh�s��c�00J&��g�I�Ss&��|>�7����f
��{dg<�����2f�����|\C�.S�Ywćѵ��UO�Ff�w�V�=�D��H*�^M����xf�K��g��$c#g��������Ζ������-`�P(GC�����w���  m�9��w#7s��ݙ�w�}���SV·s�,/��0�y�����7 ud�;\v,Ճ�e�bH[E�W�w����w߮OV���\u
/���||#5u�v~�g��z�"�Rä�P~H�M���>k�2߂��|�h�ƃ]��Y\��'Ŵ�Ooc�_Cw@Yϒvx��΅�o���O6fb)Z��C�:~�+�'������PH����
�i���S����0
��/~��n>��*۶k���/���w!�?��^�z�YM9�7��J�M�n�s:3W8�O�
��U��Go�H����P��71am���3��t����]Y;@n�t7s�9����ۥ5��W�#�/-�V-�|l�c�p��yA��g����_~�'c}��zN��,���N9{�@����M�dlT�r��w�������ܝ�'gR�S�ɍ蔾�� <A���I�~�V&p����V_�Ew8�;j�)���Y�YUq�'���>���uL�w���#1#=�w2�R������h�Q�7�1�����6�n�/b��ʢ�^oh�O� ���ƽ�W�_�㠃����~�̮,���D5���%YE������&,
�\o�A��oJJ��U4h5UW��l��Qá��s��MG�$�{�t�$4t�~TUe���Ř�x���t���W/wu�p>�:{��fY����G	v�/�[��gk4��cl����ܳK��X[�6�7�1bۍ�ۏ}[���A_�t?�^��ǔ�|��m7G��"��搥��&�l�;]Ф���e�G�eo�u�m�.��t�3��a땳y�.�]��c��O!�txϟ�>���_�ٸ���w���[�`�N�-�Fc��A����# ?q����Q�#g��2/��"�\On���r�-�wj���i����V�%�5q�ƃ�YK�x�<�h�Y���v�3+�:]ALW��#V[ϑgп��M6�^�|]��E�mИ\�j�YR���&0�D:��n��T��ɚ�ۗ;��)~��>#��<�o[9�F�[����Nk���ζC�-����C�8t�(:b鶣r�{s:{t��-�w���1��o	��i�,shWnf��UŮ�e1��m�e�*7��N�^�$36yw�_*U(�>`�pW�h\�7+B�F��2h�NyDϗ*����'͉�5�%ƗF�k�(��ue��u�5RKo��u��ݩm3"�R3���K���:I�u�5���ͮ؆�X� ��=t�|�';أ��l\gi���ʡ�9sѴu��!�4'�j#���R�E�\�W��6�XOhb���\7�ۘ�9�@ܬ����^�ʤ17x~�'��:6�k%e��p�����=���:�F��e^ݓ7�n@c{,꙽C�f�E�	���[ӻ�9���Nj%V�sSO���P�L���U����T��:Wkqb��R3�hh�*�W���9A�Q�:����/n�v�����F����P���洘а2z�о�f�c���	y��2��{��]���g��0%y��r����������y�}�|��7�}��U���d�e6�/��m�l�o�V�^ɵ��'�]j�(����=��Z�K��FՁ0��#�&������Z��Ϝ���A��PsY��[%�ۖ�%�5�_�7m,��l�s���R�U�A�=�����z+5�1���Ջ6=�w��:���Af������~�i`�dwuuD(ۧv��#t�.H��a�q�8ϖ�gY3��[G� Cz��Ij���<�f�Ĵ˳wfvq��B�\�>�u�y�;�������t�վ[�q��=W}�(�8pRU�)h�v�Df�*�dDF�������.�_}��R����Jl��J8�q�aܣ�P����[ϗtg���W)�7q4�q�\�Y�4�Ӯ"e�D_��9����玏2�a���Y8���}�ך�� ��A���Rݥxw�T����R1�,����wp���
��N�C�����;d&.$1�e�Z��s�U�O���*�0�߯z�"u]��m�#��NG���{��Ne�0W�Î@�@��CC!X>[˸���|�gڶ{��up�"v�n�4A�K��̦.=g\�5�$ڝ��/0�y����7��P����YJ֯pb�c ����6[>�;L��>��fX�;�+Z�L�7f�nl�*FU_{������q��3�ng����-P5�R���ZY���d�32��R��=�w^�Ҋ+}{JNz�E�j܍�5%7�����z���2*[מ]7�#s۞E�dZh-�A<�xNm_zb^�ly�ؚ��u�uz6-�s�=�ka�L�P[��9�Z��۹�>ݛƟ`Cu�*�9G�������X��V���Z~z���y	��>\�qΡ����ܽo%��^�du@8�I`ܯ�!gS��Y�Mm�Ξ7˄xx-����--���J�<�f/^"m�V@��蓰�մ�wg3��7�Ӑ��X�^��9�@7t��'@��5��數妪6�?o"}�9 ;�be�(������з��&d��ze]"&�0z�h&&�����G�
��/�)Y��h�R����H|�Մ{��A>Պ�ﳎq��{̱>}s�GQ��L��h�N�e�\.U��M}�je_7y��CyƁt	Y����ʉ�p�'�����>oy��x�*+�����?{�v���uy�����3��M�'n��u���&rvͣ�����j�0Y�o�-��w=/�ݩ�t-�]w{��I<�����7�8��{B/�4G�.:=y��bL�.�wFi��۟X`�@'w�T�m`��ϯ��#"QW�[*�"+�7n��O	��	�=6���cهE���6{?&S���x���v/L��n���b"3C���fKom�}|���&�:��+��"Ҙ���M{�̟o��AZ�7+6��:��U����!��R`ܚ��XpA�4T��Q#��:�Uژ��X������uՉ�'�ہQ;�7�؅��A��z�J#^���\_x�	�\�%�`���5�g�4���Y��$.VkC�l�����ՙ�n�E�Q���۫��U}p"�&f�VL;���_)���zy
ܬ�wװ�+�k�S��|��me�ѻX��P�h��nb���Ψ�wh~��>#���> �73~��xox���ÿ�$^����R�k�z�����;L��ԡ�r�7��*�����>��%f����J[h���m%eofذx���_`�nmA��D�vl��F��w�e--5ݙgVmO��Y�����@�8Dd:~%Mr�8gjkoJ֭~7��ٽ��>�ܯ>[k���~��=j2���C���7U�;s n���Ngzg�-�ݧ��r���hZ����0ݧԬ\;�p���/���*��7 �Thϔ������j���K����2����.���!\U�9gn��8����{���ݟmI�
B#��}O��focv��0 �)����{Y�ῒB�ϻ���&'�ڟ�d�=7�q�&�����|��F{9`0��^�/YLG,g��4�D�ys�9m��[�<qQ�Z���)�s����o��	,+V�@|,�����~?���zA��P��*R�,��B�7��;R�
��k�ޘ멛x����w���y�^/�bF$bF$�������goz�m#v��zP�{+���vn�gv��J"S��U�r<��Ŗ����9a��n������O�I�y�xD�"|jU���pw�
,�_�jM�*�V����7[�z���`��jE�ea��O G��ϴ���|�7"GV]pk�ی���1U��83W���7l���,w���>��sd��
v�I����ڼ�S�@ދ�~�V��b]TekY-��.GsU�a�Z7� Ҿ��P�&j�=X�|+Vu��5M�>ɱ!�I�����9uyުe4��ϥd���h�唳mKͰ59�-�gNmon���7.�*���`����~��r��-g�O7�[aHJ��D��d��8��� �_Vл�x�t�v�ɹ����h���f���ò6o���'�b��h�B�p��Sױ��y����9��O�2(�Iƴ����ޞ���})�>��M]���Op8���gn���Un�D�҆�'� �j^���$�~y7���<����ͺ����y��2aw��gd�V�Y�N\�Hptļ9F�L�S��>�������H�'|����w���� ���)S�2�N�m�q���������e�·�Y��$'ە��D�t��#S"e��1��m3�w	x�ޛ)���#!��<oy�!����P�j׮�n��&ػ��s{Vv��� F�7�F��3�:6��{~���z�8��Lm(ZH�OFb�Лč꿢<�א��;�T����`�B_�w�sǧ���}ƪ-���P"�eӜ<�x!����]z��Y�4C�x�a��k��׏tLߊQg���U��7���Ut�n��dJ��j�yH��%�U�oVz�Ւ�����q�� N��{��t���;�������V��*%�X3G��~1��+}��4���[CZ���%d��X���0߬��}oX���`���P��vCF��m�nj���E��N���s�.�V1eE�ގ|nӇE��:�XS޸��v�Jh��(��R�7���w��۴�C	u�YMs[�^��МB�����X{��f]�$Ԋ�`Lm�l�Gj�Iܕ�]�hI�2��-�_r��eh��b��	�!��f�:��6�r8��;��](P����0�dqZ���u��D�}Mfr�U�EJ���tP�	�pr�m�44V�wd��}�7+�!��K��T-��G�";Fk�/I�9�3rL�.��e�Q��yTy,�]|��A$6�;Gr�Pއ�]�����9�E�ˬ�`n��`q�Z�Cfp�b�S7�����g�]d�h�U�Z�9)[}hfڳ]_1��������q�0�%�]�.�'�`�����W*���1�8�R�f�K�RJ�":N��	6Vj;��e�'X
�j�ܞL��͡�!i��/f��M��驊%[˸JiE����Ͷ�4Y����`�J��l̨ޤ�6`~\��GT��e�2Z;G6r�';�Znm.�K�P$Hqxn$�Ff��HY@��a�6�<d�1]EfkA?����e�b�>4-$�L��C೴*�ګ,Y],:A)��ta�k�mb�/t�j��(�+2-1&��)+8��
w��o[ʝ��Y)���/�G_�7�����ݾU�ʦ��v.ڷ @�H��!�i�nNIe��Kdݕ3�"�V��.c���>`�d[mA1�1&�o]�(L���DA0�@3�c�qys.0e; *x)4�L`㻹�7ڛ�aH��X�`k��Z%5�d�A��_K'`��`Õ>��S����uĆ�:^s���U��w �ܤ9'��nj�{6���O#�!
я��A&��Y�:�ڎ�l�n�f�sRc�:�|��f��v2�/.�B�)�b�m������qS�{[�������j%�q���x��/�ي��Gx���j����.o��`ŷ��T]k�d��;�W%�<����'���A�B��WMAC]���F]Y���A��>o��/:(Ns� ��]�s������Ճ���uܣ�_+�%v�i�	Ă�l��V��CT
Zu�pq�o��+��R�a'C��7�=�N�]��JErX\
�5ЛQ��*�m8s^N8��J���Ɠ�&��L���t��{P�1�D��`Ù�45V��S-	�]Y4�1P,e�5793��������fx���s��������LQ����a_�n˫�c[�e��X�f�������zL�����effg9�s>G����n1���Yԩ�V&8��0�eJ+-�Q�5�ڛ��2d���љ���������555=��D�-�3����²�/�iCƉQJ'�UrYg>�o���h������Vffs��3�~G�ղ����וeUĭ�-�TR���ƹ�-A
)h��,EbJ�m[Z��@uw����*[ePi[HkZ��+YM�ait�3Kj�_r��!��
�4u�mt��p�-Kh%*�B�Q�
�RQ�3v��E�Q��USl6��^YFLm)R"i�E�(b��L`��jJ��P��1̚��*�eeeJ��K �� �֛/]hw��N�ݏ���*�Qk6� 򃈎1�q>5�5nk"��6�z�֒Xw��<�a��<||<�y����3��b�6ܹܼwO˳����v�q�]?H��»�S�K��L���&΁糽K���%Gs�m�WR[��,B���w0Q�M�N��Dj�����6y�N87`�1�$7t���gH$����Qw<��1L�ف>��r~��f�O^��Ij5Yq1v���:��a;�C��g]z�����`ќ-�ͱ��Pa�x�]q��ҽw���-Q�o%��$����u�36�3�E��x�gR���gz�9f���b4Xo��D�nl�7��k�Fy�
��#���NIٽ���b�3�1ؖ��0�`0��C稚��}�|gfvMތ븮ٰ�GEנȌdI�p����͑=�N�`k��;�q�q
�k��ߥ���#4^d5��=�U��z����j�-���sƲ��h�Iت�Ú�e��u�m���D���C.�	IM�Ǳ�؝�N�_kB!Uת;���ٶ��ȚA�	/r����D������[�[=���-��1�C�6vJIc{ն��
!
S�X"Z�EOW���y_V�:�I�����7w�Q��X���8k>�[�b���<r�.��W�Y�K�v.������|��o��%���׉��y�,��N)FDD3�u���4]��q�E=�Lݝ����9�o�@��Of��i�i��4�8-����oV�0z<@���l�ᚢ�U�t�)�)k�ݦ�u�]e�����p�ԭ�f��{,�'e$�y��5�J�Yzwۨ����xx��[_{��c���\?ch�T�q=�ٯ�vnr��=�x�յ�����0a��T�*�sS�1�� 0uY��v�3Y�jF�it�=�;=���n�T�%�j�Я�KPڭ�����Y�W��q��9>oKV�-)זa���rٙ���ϰ���V�Fn���0��*�&�{E�����2\��nQ���K4I �v���4�/UJnYUT�QEgȀ��N�m)��ڍ-�s2�g�@�ٗ�M:5gCS���.V�bvr��rl�$�.�7��{�S��|������qD=w]�N�+⷗H*E�|�J�:��h��NTv��N��L�6���'!��ʴ�����nV���*Jv��������N��G�wO�2T�G��ѵ�7���i�����7�:�����d��z�T��K0k�T����!�7;れ�v�z#�5�9���{BtP��H���d6�54'k�n�f;�V�N0�
@��K��C�0��֣;��q����#��Q�:���v��K�$�SzNp�p�Q���tУ�˒������&�1�w]�;v�&�z�ҫ|&�Ea��eD�����b�[������}�赛�*��W��6��u&���ǠK�����v���}IĦ�^���{�^'��A��&��z�-����ۇHĔ�V�$`k;3���0!W\�40�r����2�Ƕ0����m�n�[qo�������,����tyr��s�N�U{c��ܲ���T�\y..��GQ���:�E�Z{�Xe՚ŠɘL0��x�;�d(5���i�.���iR�~�&��?�!/0���)P��C"����5�+�mgS5�]ba<\Ž�Z����t/���O����y����'��7�Y&QK��n<O�㨸�R��>h�#=��J����ӱ�$�sɉ��%�$��M[O�� 9�y��S7��Q�mn��b,���>33o��mOI����=���[ϲ���x��r�P'Xw<��ZJ�F�Q�����ޖ٭��v��ݕ}^�L���NL��L���)�vE0��î��;�": {5�C s�>~^G�v&�-��V��Ó���_n��>z�r;���,	e7]�z��u�k`nT�f���	#6!��j&^���$�g��zYw
����ϛ�UbF��Ԧkn��{�=�f3:�tA�1R7w1�.�F0n�3��jWd�^��Vouz�-$j=}�7GA"Ϥ荍���77���{}�- 2y��m{�ޗ�ܻ=��B��m�t��O*V�1�=�d�ed�NW]mh7u�1���묾�Ȇ�I�sW���P�3�v�$r�����1u���i��ں2��D;�q���3v��>�b]�;z�kVn�������|%N/�G�Q�&�%b��U
��0{�y߽��w��陛>�`�U2�\�ס�t�&�����tf��Vբ�n���[�������w�E�O��&j��β+�UU�58�"�et��o@��Y63� 3�~0:�U��M�u�^^V�H���w8әo+�ߎ�Z��M3��U"'������/o3.�{��x�/��d� ���=��A�ۍ�~��(�dRB]SS�-�'+��&;$P��om�SHH�l�]�ܝ5��+���o>�\Ž^Q�N����ޯ���X�9��!����yVӖ�7��Y��qM�����bAn�D�z�{G�X�����R1�2�^�`� ;���g)�N;���p»�+�#�'�#z��]G:8�W�s9=�Z�ud*�f�P�6&����r�N?��^��~�n�A��8���Iw�Z��/,>2��ׂ4�V�,�Eq�j�C�8خ����.��/5�Q(�x"�0��f�:�Of��կO�~:<�S��m�,Ǔ��q�mG&Y�q3�x?�r ���y�y��k��jΰ���O>o�$�Z��5W�Mi�+�]3�SG'U��J�˧�
ł��&�OXfc@�x����CC���7}��]���a;����"ʐ��j��k��T�w�C���]=���fػ�ش�ܙa/������5ʯjZ|(���)�#1�15�.��o�?i�|����A�-P��+��wM��O�Ya.;�r{�3��r/��U��yL)}�cHUxr�=ԧ��hx��"m�Y�T���b&C��i8�<'�'9Hۢv�TK���P����^_<��۫���X��W�=}���;{�N�HYvbo�ulu�qƽy޼���7'�~��M �E�G��<����Z[��3&�� DeĲ�����y7��[�5��E	�*dYoj�vP��ΝR��Z�͐^��[&��
�[rTE2c��M]��J�H���^.��C�n����j����y3+�|4�Hx��ۂ�_l��_N�N���)[(�����F��6m'w�3ӆ+�|�QzQ��I�s�v ��I��~�o�������i֟�G ٕo�v�gqsM=�0���1�)�ήg�lk�|��<�e���[ӫ�AH�A�}V*�L������@}�Jh~7ʸc^<���vx�}�ⰽ즾o�eю�M<��$&���:C�Q9�n�����Y���-�:�����u�<��l��GJ�%�����u9���q��VK�g۝S��Ju���>��i�+γ`�ć�:����q�IbS!�;<@hx�P���l(��wH�3%Q�NN���C�v&�2���|��\`v�x?��P$�:�݁���nǯ�`���uU��N�O��#HE����������y�8D( ъ�7̂n(��wnv��'�z��������I��Ⱥ�u�����;UK3�D�FDKK�4D��=�F4�<=B6��n�I~�rj��BT��ݓڴ	��Ӟ������7�=Xw%�!���n��ʻ󯦞r��iQ�YZ���r�T���t��f��HƱ�(��	�NW���o2��y��tL�����j����Ǎ�V���W����'Y�-��n��I�*k'�!��mt�6�:m�t���7���� �`�I%	h��+vȀ,%������3�Fn��he�z틦�O����3��`;�tN4W�nz
��8˸le�"�D��IM6^�66�wT��gn
��.TmG|A$���P���sr}	��c�d=j�1���D�O�o�َ�����z����h�@r�z+H�5Mٛ����˽�M�Y�0��K�������~�
@��ff�O����I��iWuINrۯƗL��̒��aS2�*R�&���L�ϯ�߲y�n4�*<��.��)&���y�g��`�ˀO��4yO�k��%~��}��5 �6Hm
���ح�#^�@����p�����J!O�M[�wV���V
��v5-�eb7��^��9K��{"{��R�rDGC�����ɤGnt3�W��U�G
���v�N� �<�����g�|fwoe7\J�T�9�W�V��r�&�d�������&�R�̳Qnk ��1�R�V��9�5�Bj���ݭ�SǮ/��	AA��bE�_b^�@B�}����O��3��*�n1��kY��iՊћ��+8�X���%�QF��Mc�������<�o7��*u,�Ć1���wwq���ߩ��i�8~��M��o�Xc�b�Φ�3\�PO����޿���܏^���5��K?V��3���r˺̵�Y6�%�,[��Z07B�C��``�rÔ������.ק�^�M7K-�����ӽB0���B.U�|op�ܨ��:��i�0�$3�o����a�}���T�r�f�S0�������=Cz�r�L�-�P��L}w u��W�����1wT��\^��:����o\��-���~/@�V��_��C�q#۲��U�͒�Gp��Fj55�|v�u[���<	�:�/Դ�v������m]V��x���a�|`b���^���;���6��_�o�0�G]�YV���Z���q�4J�c>4�\�v������t]ۖl̑S�éU-�YX����<�$Y�YB���v-:�C��be]i�>���[D.�cѨ��vd��6wDi[n�ژ�Ȋ<s����s�7Sc��ڳ���.&o��M.Qv.�}>o�x7�y�xt⣨�x��8Ό������ג{�u����fⅱ�ٽXw7Vz�Fw�WDkO��ͺ��z���,46��R�No4���C��}�+�M�[���=�k�H���0�t�ۜO�s�����7=t��'��K�{w�F�VG��N��B܅���WLx>ʙn�ټ6�i��)�Ԩ<te׹n�T^鬑��7�oVw`�x�ܤk5z���3�)*��j���x��R�d �T�{i<���n�Չ�L�4����=��W�P��\����l����e�c�^��Ús0H$	�\�`���!�4ag]A撠�j��{���l8�8��Ê6�Ѐ��\�XZ�|�W�zs&�WSRG�؋������â���'E�S�ߞ��M��{ff���y����I?�l'� <�r$���{������$$'��O'���K'�}O�;ȵ	UeZ�Ib1H� �`2H!$�VUU�DU�jʤ�VJ��IUVłU�j�$K$Z������j�U$U�eZ�EYbʰ��ʨ�V��,H�Uj��UeZ�H�b�A"	�Db1cA��1�b1�Kń��IBX�eTI*،X�A"� ��@�VX�R%YV$�eT%Z���RTEH�-��T�`,d �X�H�X���H�# �X��! 1H�	"�0$��Bb	"H� 1#�"F준�a�@d�#F�@B$��I�D���F�!@B A��#D!F� ! �I�A�#F�@B� !!@B0��HA��"� s�&oa$� �BF� ! �a���$  A�A�A�D!@B!��	�B!�"BD !@B2B0��`A�"��$#$"HFBF� !B$�	 !B0��a��D!@B A� �B$"D ! �`A�F�B$"�!@B A�"�! �HA!B!��#FHD!B!H1����G�$�d�@�H��Y"�Y"ȂY"�A$��AV
`@�� f`� � d�2@$d H@����$��%@�H FB	��@�@�@�I3 &I2 �@�@�@��#��@D� [$� $ ���$R#E� A0 ���"@a$���!�H$#!��@�E   )�H
FB	H�A0�B(F- �	�H�*�!RYU"U��b�*իVZ�jĒT��BFHF#��?�x��C�������?�!"Kb@J�0�WB�?�����O��;����������o�����?����ɧ��'�������{�}���"H������?����h��C��*DI�O����EI>������i��G�$��$� �����>Y����I?䇁�Y���C��w�C���M��I"��*Y"X�R%�	 a ��A�`A�"B� �@`@`A��20 �`AD 0�H��@�@H	BD $��� ����b%��,�H���BA$!	@�2d@�0$@Y$F��RD�X���$E�$�������,$KR(B�@F�H2 �Aa���$�� ,  $��0�� 2$��HD2	 H A 0��$�� �d�`�����J��*D���D����,�������j�BB[$�B
  (HB�G��g���?��@�����h'������� �I&�������������]!���?��g����'�D�4�ړ�t�����'�D� I@���Rt���2������B$���D��=�%�� i%�x���Ry'����}Ɓ�4?���4$�Y�h��=I"H�O���O�ܓ�_���$I����������ÿ���a�����?��?�� �'�y����$?�y,��?��RH�����i�����?��a���?����@��y�{�	$�8�������������~��}�O�B I�	���z��W�?����w������b��L��<�@l�K� � ���fO� ćw|�A%
�R*�HD��B�)TU%A�2J
��J$��@�D��
&��""�	"*�DU�i���5M���cF�ن��C"U��*V��f�#TekZZ���mMb��%�!6����6Ե��Y[e��V�ٵ�#Vkڳ)�w�K٩��@M�����m�0�6�ZL��)-6�a+k*4�+6M�J��U�&�6���Xd�cF��ک�cm�-6����H��+i���ֱ��  �q�e�1[��s]�i�ւ�n�g[�uٝ.�[U���mv�Ѧ�e�5\m�C	���Y-G3v�5�l�n��M�ڕܢ�u�t�e��\�MeB�V�m�]�Y�׀   ���
[
\\(�C���B��z�kl�Xh�J��j)h�Nݪn�昪�ذ��R�uv��5dԬa-�i�T�Pu���]��Ц���,�6��i�m��Z�f���   .�(uF�k�Z�Lݛ�w:��gu�)�L�:��]j�-U�UQ;�]�Z ��u�Uu��Z�N�Z��H�Z�[+!�1�j���h��   ��{4���j�ф�W0aZ�@݆�Y�]�6 ��N�E �L�
�mS�\:��Ȧ�[3ʶ�)2����S3Y��f�*kU��   Z�J"����!��6�U�J����9wd`�Sv�dPT��N�%-w9sY�D�n�U��t:�*��kK����ucljYx  {�풀.vp� a`ZPJ�h 	�q� ��� �vu  �0��6v� 4�i�  ��iM���Xڍ��R�֚k� o  �=� t �v�  #�� 40  �.P  �v����� ���@ :� ���Y#j�Z��e��5��<  稯@h�7\  �1� ��  4n� �\PA�S�  )wSp  �\� ��� (�iZ�aY��J�&����  �x4 wW\*� GL  ��  v�� B���  �  r�S@ l;p (��;� (cE*%\�lĢ���i�,�<  ux4 5{�lPr` ��m�  �+  t�p 

�`  ;4 �`���h( O E=�3%JT ���a%%*h  <�b  ���R����S�'�U*��� I�"�ʪ� 4���� bA�b.k�r�*5���		��Ef�b���n��?���������r���m����cl�?�m�m��m�m��6��8��l~�������3�f�(�Ղ��Z0X��U[F��,3��d@�Gp����s�r�4i�Q��f% �
�d��5&�5�e�����"����i�.��P��k(*�����Ĝ��!ѫX��7��yv��2��Ţ��L�Sla� 7L�9�-c�xeB�H�Qݪ����TT��Ų����+Z�^͍Ta�����1f�cJ�d`M;:� �|�'n�eajU�*��C�ꤍɂ�RYv���5c*���D�W����7�Uh̵j�+z���.V5ĳXe(�	Le�oB��v�űWķ5a���>�T��YGM�n��U�r���k]^*D��[q� �y%]�P8�s���OP��y�6V���U��Bk7.�,T襚ƣrE���k��+�,�W���[�՚�B���P�ʕHkd��q�0BZݳd���v���H6�Ǻ�U����l9t�@�x�� � ��dvXem[1�o-�`�m$�����єd�r��7���ʶ�`��sM�B
�oh�,/m�t��B'V^�c)gd*�V�x.IzYz�@�W�T8(`�UkEHY��n,u�觖ma��V�1��+����$�����Ve��f�a��vX��S$(�T�b�0�w��(�������Ƥh��Y�m�X5�^�Ҳ�CcT�C�%譁��$��ʉ4l�^Y[d]�)5}�,�C-��	X�A�ƻ�Ei��2�H��e,ۓ0iz
�S�l�qHm�mK�^������8�Ѳ6�M�[j��Uz7 �;3H�dkm���#��h����DB��W����LR6�r=Z&�n(�W��H%]i�t͘z����:$s*��+�#�Ix�b�6-;����$B}%��YKj������
�61%E����O��r�����R��d��
yQ��sif� I�q�-��.�Y�����V����y�me�b��N��l;��N´c�W�&2�RE�����dw����L��f�([F�IH��gn��D8!��J��=܏����ح*2	w�P�F}�����n������ke���&����o/��ĶKT�wM����ŧv��mB���j(���d�R�j�٫���,�{)U��kB3Do^/,�ڼ!��)F��C��AKc�0+n�?���Bw펅�bE���7v��VƘ�hA�z�bR���ՇmK�E���ͥwWI�EZTf��e�Ld@�s)xZwx`쁞PqS�x�� �7G�\�61�R�/&�3�;������Ɗ�ǳD��9yX�X/L(wx
���ӎ��7V��q���u+�#IF��Azշ&?�&i@�����-�4ͻ%��K
)`t��t%1�7K0��iD�L�LT��k��hpbI�am�z)l�n�]ԉ���5���wO �1hܧw��X��z��ݛZU��w�T7d�������v� [G�%���^Q����±��ƭ��Ne��h[�sX�1e�x����јb;��)�1�L5�i�M������+9zt1s�v�U� ���m�v�)Off,z�!.�:���J�,D�섷l"���.-�S��܍�s �6�e3	�c�M�s`��IN�h/y�w&���u=(KBC%�q5z,M����.�2[�wj�VR��Y�N���E�( B�2n �S]�H�ͬ�N�l��s[8����M�Xcm�Ow(��զ�r�,Y��@�ۆ+�r��x���.���JI�g~��B7@��
v��%㡜~��t���>J��ViP�`�M���N� �v1���t2�;h���s*l	�.��CB�cd�����Q��1Q˳�$��F�\(݉z\�
ْ�ٖR��('R|�P%m�+�*��ıyFc�cS;�{&�Puy/nw5�E�p�+29���s&kDm^�ݫ����ͷ��e%و=�������Դ)��	�P�2Q����@�hW������2�v�I� ��.�����
���#kt7�Qǩ\�*:���#�rI���R���6�1Hb�SB�f�l�(u��S?"4j���Â`�`��)[ܗ7-�KW��m�޿�@�!�5��;�ɬ�Z�6kV"��(����-�b��u�b�T�m.�L�䄈5��Є�)��P,� Ej�n��F��:0�ݾ&��gV�����h�.�+� �T�,Wr�2h�uYY�KV#8<G^���`h�]�n�:y]f����%��&��Q9��L;�
��[��i�˩�Q�)鈉W@e�@�,���,OfL���IA��25bm�w@\�����$�Vܽ�=J�T5b�/mÑ�&�8-�̀�a;W��i��v2�+r^t��/iBV��6L��mڢ��x�04��U�67���Cl*K]&�����[r2)��H��!%��^�u>��TNT��*�3+	#۲��[���MI�Xݠ���kP���$����v�ۼ�*M�:Md�0E�7I6!�2���
�l��f�b�6�s&]I���&�(�Tކ�Ժ&�@nf��U���A	M���tK
���sKǻIV�Cr���O`	��ˁ�L�� i��`��DI,������gsDm�-���m�%<��!�:�VթI���Yg6�U��)Xn�j/��m�Z7#��+2�t}z#J�7i���ZN:��(��1�ow^�ܡH3�0ټ�Rjc�N�jׄ�e�w�f�qU��\:���
N�u�TJ^�Dk���*Z�kF�i2�D�*�kMԔ��ɷ-f���b �U�u�nX�U)��*ڙ,��u"����)j����*�=�SJ4��WJڲ���4�WS(�ѤCBh��]f�(�D�/h�+J�R�
nK�
��6=�V�4N6m$򅼿��,\g�N��5,ЎHZ͒�; f��ح�4�����j�ݦ�Qʎ���q���M���J�q+�mdw-!E�6�Ҩlô�7�,�����W%��8��x�a�j�c-0v2�;����v�ĎEp�1��n����nVV�m	g�*Q�M90�nt�ō�v�ű(�����dS$�Z0�������IY�D((*5��;H���Eh�oL_�&Ve����^�ä��2\�@�kZF�;/u���2J�J���u��eS��Pא�N��ݸbp8�ROXr�츐:�ųbQCn�!  u�sV���[N�㷰��C)e8	��˛w{��&�a�t�U�Ȗ(�	��e[H=�Y�yfi�x���Jmk�BU-4xm�-mF9"�)�2�4V�Ւ�%B⨵R��,�#@�W�m�F���ouLX2J*V���f"㔡���z7lc)��%͈�h+�c8��5�J�NZc�"Mk!b�*��5��Wj�Z,�gr�V��Uf��n��e�̊A-�*un��Jͬ�kZ��%b�LQ�mݻ�K�c'�tI��׮��C�Ѓ�j۰�;_�aN
̆ӭfb zD���oٳ�E�k���i������7i�x��&����e��;���إvն�*ֶӬ�I	9��x�/l��fi�r�0AOA\�]�S]�@m��7�qCt\�^�� `]��b��G�P5�wP�E��b8�M@�*��P��;P]�'0�&�L�3(���6��l�(�.�o ��!N!�)���HQ;`�v�h8e0��F�[LE�M����P��RR(!4
_)Z���쌩!���,F�� S[�U�y"T`�o
X�*��V�Y�W�zT������ɦj�ܘ[v�n���x@�liÍ�G.�Y���.C1��Tj&5����[3(�#�ڑm*��p ��Dr2�*&FU�vYu���V���V��EN���))�h�5�r���[1�a�k�s�@%F1��le%�R����Ć�l}y�bϋF�Vʹ�P1y���� �{l���
V)@�����7�FdÚm�5&3F�ܬ�M3Z�6�ª^R�\yAkۄ>�Y]bh�^,f�=t�*Ml���AٵDbua4E�vٗ�;����	��^���ԤՕl���mh�A�H��Q#�
&Qmb��P�]��V+p*5�X�-�"��ܵ�JYf���Y���?�Ȧl�f�&�i���ਮ���B��O]1У7b���t�3&6�r)O���Q��ȣ��V�^�гl��sq!�K��d�m=�q�+6�'��#�j���m�}r򒺕0ݶ]����j�ʬ�=tB��T�!��n�>͚�ec�A��{om|��tJ�6�U�(!�C�6�Q���A�����M�T#v�ن�bF�^�d-h{����41 ��d�y5�n]��T@�er�ěM���,#tV�Z½˷��y#�a�j��j`1m*�`� {	��FS� w��]E�K;I�a�7C.F.�+t�Ib�Z,눚N6r5Xem<�O7,�;T�V� ���g>Gp���ZՂZ�[S�nRYH�Ѳ:V8!E�z���	^��Д�wa{A�fc�n�r�!Ӆ�0�����{�a���©������V�6C:�=nY[�[ӏ6g��a�2궚)���Q���]�bTŉd�l� y�x��:����L`y.m��w�-�Z�8�P�'@U�+�n���Z�$��;	Z�%`Q;�2�$�·ɹ�I���m�&1�)E�Yj��� �F&�Y0�/{�P��0{ۡ�<&H-�9ˣ�b�Kq3�jh8��(�leWX����D`�c3[�`���;ҭ=�-����n�:���P�H��F��Y�.���lU�rїq{��R=�R!ʻ'j2�*.��AM��v��)<4�ɦ���y�TC���7�VmE6�!I���Z7D��M��<�R�[/5�R
���0�H0�*
�ň���Ȃ��ͫ�JɘPi��c���;W.��&�R��&2h���۹r�ݫ+,S�l�.��*}OJD�jY{��bڙ-�u���I`�b���Pi3k� �T��Y8��!�b�ui2]Cu��1<�F�%D��RW	z�/l-�CF�f=u�m ��]��N����Y�YR��[5m/��P�O�F�v�|����-�J��[N4^�.�aHz�� �y��0��d��\�Nd;{�,�v���V�h�귰z����\yn흔n�;�b��$��ʶ�l��఍K�d�7M�\�u����k1Ĳ�)V�6��f���ݩDS�۽�f����R�ςϲ+���B���f'����rS�6�:]�4݌f�N�Z��0���50ڸ���>ԩ 汦����1�/7,��qn�+F\�v�t&��k\O]�4�}xq(��U��-���4Kx^��t��EF�j���U2����ʷiK"���ΰ̳wz���V���9��"����	�+*�Ye��	��E���&�xU�R�r�X�%&=82�p6���+��볕0f�3T�R ���*Abh�K+42]�Ǳ!��$�l�v��^�hPb�1|�h)$QE�i�)`�V=SB��n4*
�]ފ(�D���k	F)aEX/2�Z�jcGLQ �@���"3v�/=��僵�K�$)r}����c���Җ�5X#hY
��[�f��f�Vg֮'��2����{�e�VXy�#�R�NV�ʖGL^g%�G>_;�VF��Mˎ�d:~�kB
1Xf�ZGd7�+�mІ�TU�RF�n��h��Z���F��6E���R�:��YKso5��>��գsae�Z,��X>!TB���Y�e�vt�K�ژZ���yI:E,X=Nk(�LY�ks1)sk x��Elߜrm�n�K�I�z�+�˴&ѡEȒu�����b�J��C��-����$Iot��wr�w*:y@2m�����^iYP�k�\�Ԟ+�(�]ݦ���'���ݡV�EP��4���̪@�B]h�v��m���&���\�pee3qY����7����yN6��M$-4g��ԍi���<�zM��T,�3$�k���f��B̭�v��+���ݸ������AX�2��n�U�l-�����v�3q���.����a��[��`��R��/uV�2�ٹ���i� ի0͵�"�;N�D��Uաj��淕%���GĽ���*��Y��-jlӣ��ܺb�[X���"�6�l"��P�	ܙ���R��qjM�NX8�?n����+)�c2��S&�Q����3#�ٌ૥j@���1�7�M,%m*#.
V���D����ћ�Z�~��˦��NJ�.�����YraYyø�2_n�ݔ�0&F�Ȁc�,y�+W� ��j�^��*/��.iܨr=R�i��d*�I���,�)$�ⰶ�J��p�lP82�݆܂�
�m`�N�'&Ј���m�r�L��^k�����sQ[m�:$�^ЗR6(EL�ֶ�����S �hnb��Eix��,Pt��]-p�E�{n����7N�¨�#��\UfQ����T�ڂ]�W���-![`cj�)n��@�U�� o�b�L%f��&��4#�[MKb6C�2���n񖈦�v�\���f�#�&��n�)�t���v�I��
�-M�j�Q�2�&Ƃd�"�Z��x0�k�a���X�F��^�s�Yn��k�����)�NF-$/eV�{+�Xa�4�Θ%��je�5xY�
��*r�9�W��+��ml�4Ҵ,��H����[?nb��i�ɸ����}(�Ƙ+SN%�rs�/��W�5�y9ؗ�ӛ�x�o!;OV�T�m!�&�,��Kw�[��_����x1�fopW��>�p�h�vd�dX�e3WJ�h�VB��ҕ
�8[�w�5<��H�?>�* J y��;��y�/���5�6���[%�dnI!�Qhu�nMH淢�gc|t��ph��,�!�}g�n7�F�����ut���)�"����{�����Keޫ<�}Α��Z��˩�xRZV�=/f@nP��Q!���λ4����B�
F�,T��!��\��;�a�u^<�r���!Z���@#v�NP=�V����j��$ש9�|,Ǜ=և�oz:ǖ�ְ�)��c9u��i-n�Hk5-6�-���[a�ݷ�\\R��[q:M�t9�<���o���2��9������.��^����'*/o����W�ǥҒ���/	�d�M��8r���IT��K�wC^�(�]�Ű�2���BDy��'��G�
���//4��]1���ޮ��W����I�i�9U��0QX�вf�L�7a�q��ڇ_JD7�!锦W_X���:GI�i�=�.*���[� ���Yޚ%�ג����tp���m�	t�AcU{s����{5<�;p�i�*܆V��&�MhѬGG+[�.�k��Z��l3�<q��c�q�[�BO�;��E���7����Oq>�A+�9vS�[��'Wb�#5-�H�q���D��s3�DvIO-nv�s,���f9�ʊ,�]}�����pf^�<��:lڨ��'�w�A�p=�0Kd�%��F���i�D��Z�xߴk�b���X%(i~��:�r�^է�#�"�[����HR�칖>/��&h�Y�X#%�D����o�*!���q3�V��E����c�I�P�9�B;�9��`r�� }�&͈�[�{��W�+U��z(�u�<)������qʺq��G��%���V�WI��G�2ٖ/^e�G�|�ѱ�|r^��=!�L֊{V��o�:7MT%�4�w{�N��;�2�8��>.���M�'��	;X1�udu���������������sǦ��௤�w4��'ż����Hؚ�p��ܻ|�wM�o3f�m��o{��z65�o\��5͢�j6�E��3L��5��oڃ�u�� -��B#�ojuN��ח�1;h��c6Yl�O�I�z�>�� ��Kx[�1>u��.��f>M%�륧������O�^�t{���E�N=�-^C5���KV�e4�&�n$"9� x�^�S#^�u�VY��U�ҳ�v�<�V�X$��Ƿ �#[՚P��q=M�l]�G�8��6����آ����Uw��Z;�߄�)��o����v:�`�6�iV���.��3 2�[mܐ�H*94�3�o	�;��7�5\k�;[��h�NŰB�F[�����+9{6������]gW+�z���GF����t�#ei|宮
��+Q�4֪M�i)�tC�r��>���]�E���Wq�M���Y����1��s�Q��҂���r���Ⱥ`y�s��k
���gQC���J'�J�X�%h�bV�Y��u6��N�H��
b�:@�3�niX��A4^�B)K����J�k�[8u�o5N�<�*]^�	�|�æ��?
钡8���e��+�4�ګ0H-�F�Mg�$IF#r��*�n�L�!�(��W��R���^}��P�Y�/�iUٝ�����Z��������]/@ݴ��.�:80Ǡ�L�I�����ϡ(�oV�\�w�\�!�Ȯy	�f�Es�Y�A��w22S�D���ʘ�f�W듛�ڣ��]֩6�֬\шM�j��Y/���WB޹!�F^��jaMc�v���<VB�u3�Y+��7l�Y�[���QJ�֟G�le�U�՚��n��U����ܝ��2}�[��5g���bg�!k.�W��g�u9��l��R�w/�%�����m���tR'�1�G��ވ:�����%v��R�.�e�����I{v�QLG��{U~$�U�>�������:T�h��cn�P�+�mu����t�p����kA�f�s��u��]rїan�*�U��s4�:�e��e���'�X|j�'}}��$3������K�ׄ}ohܲ�P.�R����pDXm]u�lef�if5L�N��J[������ݎh��[4���dJ-��P[ٯ=E� E��2����Wu��J���KkWMC�}��Ց�]����'v�u�y��"���ē���YZݬ�n��;V�)��"$�m8��j���VI����87@+������s��ojk��7�NN�3̷�jX�pې	3e8&�Q
���{��KmꝚ�	+8)�s��EP��b�'�c����P�U�\���W�7,E����ɁYWYu��[9�R9�i�b�s����M���A��nw���f�S�{�5G�(`D�w�����W��j�˙2l�7�l�}�6��̥��9�e�L��!�y�wP���XV�A�LK),�!	_^3Ij�-��\[��y��A�l�I�,Ծo��&��Ւ�Ű:�E��+]���4#��_hq7�6��"�����'o��cU�#H4 \�r��Xz� �����V�k�u�CFۚ�2��]��e �ڂ���x9�Vo�w\�}�n{ƚ�Wq�
��Y�;��b���r�U���!��M��{�c[sHH�����O�ˀ�
ˣB]Т����v�u�d��&zZ�d���}_��ޞޫF���>�f��1
`֧�S�����Ԑ�#�K���/��rl�K�Ȧܔ�.�����Mb�̰�d��RV^�� 9���}Ȓ{6���9��-��&Rװ�ka�a�noV p��n�3���B �S�'Z^����[|��m�0�'��f7�Is��^������:�)v��xͦ��!])�g�W���.��u7'&>���"�ԙX�)=�;��[�橝9m��Ac��u��VF��E�o�b�*J8�hL��b�xͦIbѨ;��̑�AK�}����d��
R!��%�J�
���F��K��X�������V�v�e�:�.�7���kfg	ݪ����鐛���,1Ӑ����z*�gu�[>"��W��5<k@|����FT�&P�Ȋ��Qa�]3Q��L��v�Γ돹i�<Hw�ҨX0�*�)w#Euq��g#�{2V\Ԯ�פR��uk`Ǩ.��j]!Zv2�ff�XV$:��Q�k���j}pa�ma��yØ\t�&%[�>��dW$v��ʹ��]V�����g3ȋ�{3,7
�z�_��#p�KPm,�+q�	m�:�O^�!��"�vX�q�r�c[�SI�ΣS�; �0��gL��F'o�}r�Ҵf�sC��x��V04uJ�Pت-��LT`%�����l;�g���%l;G����(��JEe� Z�S��B�Up���V�8Ƴ
���J�����u�i�[+~c��ֻ�Nr<�S�r��S�C&���ѫ�O���y-�zņ�#ܙ�]x�%
&ή\B���e�%S\7�@q�]=bÞ6�v�E��n̥Bh
QVZ��Y@��7��3n��ޠ�ٜ}�C�&ݳFe�x[�۩����ʷ�+P�����=������M�`��5u��D�U�96G9G�Jm�+a�T7x�9x�^��՟2�8s�:��95����F�sn[�"��F-JS��9G����O��
��ŵA��`Ճ����U����:we鷪ſ��#A�&��#>D��f��F��N����,��$�護�SU.M
]٬K��RH�R�Ϡ]��������k�[��S�]�nf��&mɓ��۲W)ZE*�n�X+[�0�bf��q+{��ʼXF�<���w^f�dQ�Z&;�}E��$Y��ܐ��n1Y����[��ee�*�Hur�L�Bõ��O�^���]ʢ����S�WvzR��Ks'�i�Ӹx��+x^$z��������t��[�%ɢ��]��]������G�$��vkVԳ{�b�Qu�ioV���M�rC�p�Z�@�XV�մ�6�n�5�c\��*�kg2�lJ.��E�\��4`ep�#,��$�؆@2��bM�+��ub5}͞��J�dk�9��x���ZMii�U�7YS��bd�χ;̬�jV���Ā�Ly�@�I]��;�	f�AH��ج�#w	�Y`N`.�����O @��Y��ڹ��T�Q�b��u�S3��~���[�x=����"����ᙁl�1c�y2r�]��J����!X���igvU�v�8oY�i��VKg�=�nd�Z)JC��sw¯f�fجM�<�B�Y���8��5�X�Ĳ�N�yW23���)k%o4�H�0]��tfgga3� {�hB��!�m4OI^r�����M�r��5	��6\0�t3����˕��n1 ��gE8��V�m��v��ޔ��+���5��"�*����P�[H�CV�k��,l�q�u��@�f/;c�xaضN����ڎڕ:ٹ�92��Uԟ�Z���m9�ծZ^Po��[#���b�ZiJ�оst]��8�)s7R34��r녳���꭫����@��1�[�+�V�n�J�(Z���B}�A̵�0!��ݴ�������b�����gެO �����bf�m�ab|��.۔�}G&���zR	BfDN\��������~5�I�V�\ܬ)�KCL���4T�|�[��ۚ�p�v���wzͣLŜ���+���f��wb�������5Tx�������r���Xt#{}Jk��� 7�wcA�o-q`n�H�
�>��{�7��z�Y����WfГu혟V��9�wj29k%�������"��W�$�p�
Am�_���n=�Kr3�wj�r8K{�+L�<�s��ϣ
��7�@�k�{dΫ��:Җ�E.G�]"QS���9r���Hr�e�9��f	Tbg��G��=�Hv��_S�~.�)�}N$\�y���&�$PX{��FԦ,��
�3{��;�}�z�d"U��!Kl*;qk?wqT6�2��,�{.�F�M'΃�ǚ�ܫ��c������^K�.Z��`��׼9l3�fkZ�W5;jm�L� �|�,q���J�Zz�ڬ\� $3+��α;*K�R4�P9�w�f�̡��p�e�1�8�-��Ǐ�Q�؜.�s>ݹ�7���fv�4�\9��t�k���u��ͮ�Y5ߧS��U̽�q;�uj�c�a\5���'1J�bڎ��K��z���P/�|k*F'nv3vs�
��@�(���W'���8��n̝�.���R����e�3F��_�0w7�ܾ���[���pA�ukG���:���r��pr��a�x�m�a�b��8��zrfm�Џ��V��Vu�t�P�7�J�8:+bs�Yt{-"��D\�6�3�j{>��^h����o���Y]�Aŗ�J����1n�t^�����`�Z����G6��H�kQqm���L���U`�@�X]��/)�C�ݚ�n��؞)k^+{[z.�H��1�T�ԫ��N��2�m�i�\��s��1��Y��3�f�+
U1Vև|�]L�9}G����9�K�N��t�$��Z��� a�;]]�>����[p n������I�aw�h�v2��s���.a��<�\�&�^�2�K�{M�]�����ɸ���ci_s鷖�������jj:lC���<��a�����0l\4w��!���x^��X.�k�u��ܡ�9���g��!����]�`��4� e��Q+���J�%"\O>u�Z������&+�o�����l ގv�
�c��u6��e]4��W$��/{��3��.�8'��IYS�u���2w�ӓOM
t�GwL��R`�gG'�2֥�Pyu3R�R�Q\qI�d]u���E]�X��eMz�D��u<f��BfD���I��8ٚ����v+����Px�z�l��U;�fݦgp�������@��u�׸S��4`���s&��s���K+�wp1�5��"�9�mKD̝�n�*��@��&��i�ޝ6��^5r�f�m�l��:����z���*���f���s�C����*1Lo�\����"�o���K|~�s[�|�ލ�Wb�Y�#��!���[��A�Q63�[�Չ�v(o�J��6�	�Q��9�@�hU*�v\������.U�7�a���^΢����f.�Dd86U�K��Cij���l܉wW0b�m��˵�	���ʙu*�ӗRw�cX�#���̹{КU�[o>�H�@���;/W�P�=2�+^�2<�ףu*�����ڕٯ�;�;��x�imZ��q�܅G�{r�hsX�v�p{��P�-�+Z��^�K��q�7,t^K,�(��t.r�FA�Ϣ��Y����h8ûI��G\{�x���XQ��:�an���v�[���V��M=����0���u¸n��	���n��%E���H�Z�Ɨ��f{=�8F�DfS;�}P��u�׽}��S{��˳�:V�;Z��=\lM|�&�E��8[��f�r�;���ٮ�X�as��pZ29W% MC��k�w7em[��!;<�|�!A�B�,[��Ӻ~Zz�"�k��h�X�#w3)��d
�&&����e��w�;C�'t�W�`sc�U���偽�lc.$1����(_ �@Ee]�l��rSw_�X
-8�TBx�V��K���������ݻ*�r�~Ѳvl���V	^��{�b�}G.���Cfu���V�_Q��|�������I�5�$;�w�:l9è��ѹ�e���x���h~�W��o=�u�m�Za��i��[�3e���_w�����6`��M�m����}G�}�s�}�o���[vv��@3���?����띦�2Yw�9Z�_�v��I������Iqk*�K�-��aK� E�󤥷C-MN�v�h��3(e\�K\;��e>�vV'mq
�ZW�0��H�(�Z�]˔5��P���z\���J���~6):f�3+x�����G���vӸG-�,�w\�v3���i�e���4i��ƏMT�Ó6��2�[�/IyS	x�G)�l溾�*l�s�Y]�S��oQQ�H�@wR�lL&�!�l4{D�[�C�n�����]�+b|���:y�s �N�� ���IWgB���x�Ay��o٧�w���y��2ٰ����\4�c��X�=�"������S��a|%���G�Kb�Q�u�M���k~d����dMȗg'A�xL1��9/Lf����HX)��r=�v�锎m���:�iI�yd^�HY�-{ӊq9cy4]��܀�u�
�A���c%:��U=�]� WQ�o:Ζ�ܻ��'ಠ]d�9j��(�u�ZR��w����ݬ��0[`�	��f]��� ��i��͡vxPPS�p:h�Ӻ����̷�D��v���(�Q��%��cHe�l�uQ�,�������j�E�y]�,������}�P4Q�n�	e�؇�	q�,s�5�j����-	�\�ɥT$�o�f�=�M:rVܼa�G3rάM,B���n��
}�^��#�wn�NƘ%�5�R�4�]�*��Oй�.mйi�f cx+af13�2!j0}b�0�ۀ�2��O��b���l^Kɦ,̋wn�B�pڃ�훕���d�@�xt��k��e��y�fG��%��Z��MD��+C�J��I�;su�VT|�Ǧ�]^R�[������(���>�G�"SU��ܖ&m�_��P.c��gb���`	vt%��պ�Db�YiT`��y��&��W�/�n�f�����vf�^4�`E>L��x�&ޣ�����ʳR��}$o����Ѵٽ�I[�8�j.�+
qȷ
YGpm�!{}7�n��[�+�vVNs[y(����u��9��p�_^��0��Q�vb�{X]�]�kv��f���a7����c�Y�:v�	خQU���b�~zގJ+^�X}.xb�C���wxA�3ׂl%�S�����5�vr��j�3�bH�M�+K6�����݉�v�I~�}�#�w�d�6����y��+Mݦ'b��cܫd6�#�ǯ h�}�(�Om�"v{�\�e��Śj�}��A'G[�ӑ,b�.Y]�A����j�q��U�ɱ+���mѭ����k�|��Xn�j _;��ZE�	(gt��V���ge�.K�#���$yo����E�e�����j\�{�����5� �Hp�
�N���k�μ�-�}��#48؂��]�N;Wg����>Z(i�4�݋�*�o�u*<�֙�YoI�nE�*li��?�?K���gj�g_QF�[�uN}w䶺��05�t���ӸZEE�dT��sGv�ݰ����]�j��"�vU���0e������8��+/���M��&_;�u&m�՛Q�ܗj��n|��n�/vc�L
{��r�� ����������B�,wt]��vx��I�ؚ�+�=��ʼ�"��.y���O�ׅ8��Nj����0��(�P�,����ı'[�]Q�yZ�]1D���*���(]�� ��{����0�nRk: N�-\�l��V��W�98����Kۻ�8���1���G��{�*����=�a�JVqh��7�,7���sk���MJ�#�Q�}�;�U�C.�� g��9\oYC-��%�{3�B��A`�r:gu��1V��ei��]|TS9�:5ֹA �gxxo/T��d���:�vaُ'_?�܇�3N��[Q �-T���vt0�A��I#5N!�Y��9��Qe;�"��W��qek��u'�kf.������J���6#��=���U�P�_Y��RdJ�(��A�%]��q�f 48�Qzz�E�lG�"���L�н�v����::�"K^�%�3�ޕ�E\�fob�rMb�h�&
�.��L�&#�x!/��-(k6������Ϣ��o��*���4��ު5�]zc̗�Pm]ʍ�
HCQ5z�@����읫)k,޺���8Ild���3S����8��|�,3$���Z���!���L�Q,���*byB�ڴ����]�@�I��{u�MdX�ڔ;����]ڱFm�h�;��D���1��U��x�=�v�پN�+xA�2���2�=��m.�ˤu�VX��,i�q̘��՝a��mc[��+�jZ/i��Pki�g��:ۓ{��P���m�q�G{#%�06->���.���g�.�5�Qb��i���fpo%#s�yC����r^��MK��C,s�/�sC�J�^�y*��AA��3���xn��f��v����gq��Lw�o_I��!-�E4:�WE��2P��7E��{��9�ni��!�+S���n���r����NKwu;�S,�ی��{�)�dUH��1�`鎱GX�C�� P���
]s�X��Ok��N"�r��\�띻���Ӧ�܆V��-ۣGô�y-�(�Չ2P�D@��_�H^������gC���%���;�Ǡ�̝�vϳ�t�3�Y������gN/�lX6]��9�p��:��3�;!��<�^�����O)lt�U͗v"]-�S	��ǖ�N|��483Q̓F��{�3w���-�;���-�]���6��Q�S��7�R+:9p��v6��OM`�^S#$2;�E{u�����#妤����h��q��׻l�[�A572�*=����8�:�J�Ktf���ힱΦR�wcJ��ʻ�+v��rlWV�������9Q��N:4�X� �"qXō�s���ͱf�.�±Ϋ�A;� 9.k�$�W|���A��W��Է�!��%;	P�U�.j[�dݓF�b���+��)�؈��r�[��]X/�IT�1}-4��9��4�'���7c���R���t�*N�s�u��a1T�p��r�௶��a.]�"¢�۾�;�	���h����GA�Lu�QܨR��8�/��R��M�Fvk��$�b��ܸ=�{���"\4_:���'��2����H�[s�=���2�F������=����P�)mڧ;C(uȮ�4�;��1j�h��C9��Q��V��Q�4���z����:h�v���2�tcެ{�Č���*��e^@ީ��3͝�)�ݷpo��
6i����׵u�o�i �Z�`�9 /�DG3��.���"ty}��u��9J�β�ڄ�
����A��e�q��ը.�{�)w�L�r�� X�NtWQ�"ܩ5�6�-��Gu�."�u������AN�]K��`��Q��W�*���m��u��ĩp�Q�B�(�h;B��)\ý�6_;B����M7�d����CZ��{,�U��f�Qa�.deЫ��*]���j���J_=|w�JZ�fom#RgZ�Z�ggP���`��-�d}C#�o��Fu�Mn�Z�ٶ�ըv���B��=(��ɻ�lU�RV�>�Q뫭P5�y�7��x�K2�{��(C;����6���&��҄J皴���<�`�1�U��Y�_���l��04 �ٸd��9�]ƛ�uQ���|1����׷�Rܷ�!��d��GcDU��؛b�L��v'�y�96͐¿����|F.��=tt�Eȸ]$hM�a�.�<���	Et�[�n�\#����nS�S���������/h�/h�R��KM�����pu�(�OoX:%t�}ĦwkfϷ
�����AUY�Q�����y������tl�T�u��U����t���K]1���Np�ƛ�&��xc��蹁Wyƭ
���"�۫�U�;m[�[�y���!�Qōd\;Pӽ��w��l˵Iz�tY�b��\6u>O<�b�/J0@Jw��e}��
�L�t���+{s t�vھ�uэy�u��|O<�ޙ}Ŵ��>|��d"%7iu �'���#�� ��6Ȋ�.�opہ\kJ��ӒܤJ<���)����C���u�
�3�X:�sV�m�R���Jcl��U���2Z��|a#Y��-��nQ�2�f��ae�5)�&JkX����� ��)�ܡ݋m-��m�Y�&�>����h��p+�oZl���<֪q��$��޴ҭ!oZJ�]YmSY�� v$@j�-�}�uO��6��t�Ô��̅�al�U`��E�t*�Jo�X���cvBx��؏SŰ`<�H3�/F��_=ۇ�Ԕ�lv��J�i��,�J��԰_�����Iy@��N`<����-�tK������G�F�ruՠ�c�U��<U�tg�'Y𶪹��8�y��iUop�L�C�����ݘ!�$G���5Yݣb��n�xח]�,�gqǜ�Y�/g��_Z�`��g8\�n��Wս@�c��������fK@β6�w�_F�G_n�hp���cI�0�ȿ����U���P&�{yN�)d��*�L@gP�:V�v�:�j��%�9�ݗ{^�58&Z�"�`���v�2kk�@�S�1��dӖ/��Dk�I�Y/�1GHj)�;��p�-�z�^֏��E��~G�b��ϔ�n��tü�����fn_W<{�-��v�=��N��5O��_Yw~�6�<4�Jx��A	y�) �x�s�Dܨ�dK��՚���w�Fq�ܒd�#ْ�� 0L��X���"-�ѹ��Y�4�͋��z��'^@2�mw��1����S�E٭����|��:#+�
�z��k)�UoS���Q%����2m���g>�#`�0��Q,���{���/0���%}�񈹁A`c�����	qWhT���o%\{�ר�����m���bĔ<�Ʈ��'�%cү�\�ۤ���*���6�
�\� ]+n��"���s⅙��@w�c�Ԧ�*}�.v����2�=弉O5�B^^yT+l�r�v�/DmZhudS*8vIX^�q��Z�7N5�$��(g<�V�Ǯ��*�C�*��&�d�R���n��Tv�ޅ a@�>cf�S�(��#54��}:�4����#׃%��b�'Z��Zf�ѣ�A�y�Mp��kf�;�3�p�q
��g'���#h�g`V{_%C�K��汖�$���=�F�1���R[�ṵ$8�����1l�j]^���W6��7�.Q��~*�8"�0��#�A4Y��:4o����Ѩ4�����`5c��pfj��Q@�JAә�A.�sɌ�bB,P)�Tw��meqRiwJ�s�f���յ��ξ�Տ���v�<>��>�%]�K�t�J=���SMn�t;�R���Vf�m�,5/&9qd�\X������t9b�hu�sz�����32[���vDW&��xc1�=�8[�r>9M�;�-�ڴ�X�wc�0k
�rE�ģ��DwVq���V�v\k��Q�'a�@�̞^���
%�W�������.Tv�7۰4�ke9R��ݷ�"��%�^1E��5����k-��vìu�'�BD� �X����x6�N��o$청��V��
�\��_Sڄ:-ाC\�u�ji���ζɸ���wJ��n�/��*^��9Je����s�<їBR�N��fMר�M��+�����M����~V���P�L��m��v�l�FÏ�E��utfh��׵8
Ȭu]6`���	 =3�A�&)y�㮭	�W!�7{�m��E,��t�u�SC� 1F�5 !�w����\�#��o�wk�<�������8��v��鷶��Z6�#V��YV� ��jS$���S�ەD�ʳ�Д͕,��|tb�Y�7ss0��[k�8)��:�9lT�f�1�M�a��[� ֱnY��/k�i�g=&��嵡�.м�ɻ������#��F��b3qh끷�s{W��<{�+�u��A+��	�,��	/��`��"��Ji]f���i!yXڶ6>�f�����X���wM�����t���FSc�E�x�7݃V�/ys�yd֪�S��1���h��s�,M7ރ{��z���nm��tĢF�Гj�E�T"t�c����fMLK�Ý�Z�ul��u\�V�c�ǅAYD	�aɔ�OX���e�ױ����9۩��y�'x3x�6�5s���tGS�٩5w^��. �.:�/)P�:�G�ګ�kٞ���{��起��7i(�!O�<��mX�DS���m����6ݽ�e������]��=�)�@z�$���C6I]ś�v[�ӱ��`�&^�n�_|n,�]-�,n�s�&�kS%:����H\c�,���;�*��A��Icn���yt��)�&�w9{��1x��I学�F$��;)�o]R�ؘ�9��`͔ٔ������F^�jql�W��f��Z�����u������4N������#��#��gn�4��o���A��@�6�L����oy��maE {þ���mܦ�rV-�Q����+ؒ{���/a��D��-hP����*��Nʖ��U�eݤ���
�!E�l�E>��b=����ić:t���Q͗��<:(��#z�Q���u�q3��Y�
tr�A�1��b���˸�Vt��2�ӑ�E�y�'��̩���������}�]����sՅ?],:��RT��w�z\e�Wx<���%q�{�#n�0�b)cI)�;��W;7f�IVt�'r�t�4*�8P�Sx��n�Q:������9Q�쀘��ښ���j��v�4��k@���w&I}�(�NR�טfq��5�;�����vzt���Vx�lzpb�\h�.�������Sn<m���CfE�|���0�s��\h�#�,=sCS��&�D���x�OW�ͫ�N��n�r�V�`_pY�K�9ר�ާ��uuʽy�w]�Hu��T���&�t�����C(mJ�盠b�U�ژC�G�L�ŭ�,��҂�ۍ�o���$�Աe�kq��*^�G4n75�ɂ�r��r=�L�m��E�l0F���o����x{��3F��&db�#3a���(�:��
�r37��n��{n���ފ�/<���i8����c(�ys%�����C>N�k��ȕt{,)�zM�������,�{��4Ge����|�U�ݶ�"צ��5΀N�!"󚃝��i|��U�ڳ3n]�ETe��LQg{�[C����2poZ���m3�W��S5��8C��!?��w1WcHZ���8S�oZ�.�g^�(M�8��q��Q�G}̛h�qƁ�ֱ��`Z=���z8�;�H�:���ۺO2�Sr���l����\��IT��V&Y*���O<!q��T�3�r�$U5ç.���7.qt����UD��4��AT���(�QFA�!$�`�,6��E�jf�Zi�-��4D�U�	����Z��W�\U%��2(�+
Pʌ��5.����ꓗܨeQū���ha�(U�*'���I���#\mŘ�Jl�����p���sZt��Pn�<V���戢F��t�A�.fqR�NkM֊Xi�*�	AiJb�3)eE�Q�BHt��/�r"�ER�I4��$�9+���)RaXe���ǙW
�(�!]RC�F���9I��DUK	�,��冢�S/L �'���9A�,�IZt��r�"��QUiB,��I�dGT�.G�U�$�Ѥ]2�u˙�DG8��p��VU�u6�b\� �3m���#�[5+��;�H��=���o���[����y3n#�}E~���\�<�6�Wk�+�]&�F�!�!���r�<~��zD��������ډÏ�L��}h��S"!|/O3��bl:) �y{��|��j��!���s��Z��Ld�j��g||�
����s��7{Y�Y�ּ�~��j]�S,�.fj����k8]
~?/�џ�E}��\��~a�C��u��m��Fzs�����֚��s=N�M���ΐ�^�L���|>��^U�"����yh*!���jMi88t_�3�ۅ6���Q���g����84A�j	�c�3>s����W����7r��V���I��x�Y�֫&+�z�&�*��[g�}��v`2w��}��W�!~�zՠ#>��^�.�/�r�k��^�g�xū�T����;~Y�g^E^^�܆�'���U=�Έ������O�54��u
/��K� �"�����>���ޅ秹�!�j��=�s���d���� +�UB��'f<C�@y:�#$���gG���rF��^��S_[)�1�!ϵ�����J�-3�w2�<���dU�*�xkD���(v�G)�ww@�nz�}�9-֠�7��9����rt��%B���V��S��k�#���6 5���Zv�����z�n��U��縗����~^�r��J�n�������Q��fd�x:�)[�B�\���r,3�cr8��;.���?jQ�C��'�k0{t��=��&a�=�m 3x�Z/��{�����;���=�5 
�[�|ϼi�BǸ�z�T;�y����Y��qX�$�V�߼$�e���lͣ��v�CΡ@`��U�����Y�[������J������Zʝ��F�/SO��矠�&vj;������G
�[�@|+�԰��U���	�ֺ�w�YY�݇����.�L����Ɂ"a`�O�Q/jf&�D�C7��6���.��<����0$�#�	��Ϛ�+&j����Urȿ��b* �9Q(�~ԲC�X���S�j�ޫ���������:�[ͣNj�ĺ�^���繜 1���td{q�g�'0�,ل��V��]n��k��E�kin�N����^��C�����zS���0���a��kk}z�n�"6����Z�Ac�8�x:ƫC��bn�o��{6�@���'�݌M��O�w��J��s�s8�<v����EV�������	X�hk1X�G�3��ȕۇ�{��^.��o.�u�罋\�gl�au]�� ��{֑Wi�k�p�:C�qL�e-`��;�;��o�B�<������Z��g�L���CS������.�1��֥e���Ǩ8�����h�ry#���oJ�=������(��g��6�>�����t����{K��>ov|+X�p�39I,�RY&f\j8����\ �|/.����l࿺�5+�X�^-�#&��M�n�|e%�Fv��=��C�x�_����U��x�.�¶�[��=u���r�35\�5\�]�[R����,R�1g��V+oʪ�w+�p�62�m\5�����n/�5��yJ]:�?j�� p�ɚ�1��&nw�=���?�\��rc�.�:��h8�k�z��f���l/��Y��μ�uX��ͭ�Z+�6�9nR�:��Q���vE[�Z�ҏ�>��7��oɎ��ה�� ?hT{
����p�>�e����6����y���A���ͺ����L�MCFZ7�f~X>�-a��r�B�Ugb��.|���,�D?�ɍ���1�
n>`\7Y2ٶ�uP&�t�+\�ڞ���.�^8���wn��3�)���α~}���"�S�Ǚ1w�G��n�2�?#��xT �i���s<�����}:�d�=䗗��֭zI���z�=��S��yL՟f`�.�CiV�<�f���7�!��:�ɵ�4}�y��Öv�{U�բ��7��;Ӏ:����uCЙ�����I��
�5�)�K55v<�ݹ��O��c�N�B�����A���w3.����Ƭh�^WY�O�n�J�d��۸C��#���Ê�½�V�@�	���b��c�m\E�U�G&U�y�/m�k�0���f�??��k揬@k�!�-�leҺ6��[�q��x0��)�&n�ӯ�R�/�-���7��S������뿯x�c8N��W�����G~���^��{�;D��S�|�mC��C������6K��3S�EX����	{tZ��{tyu,��^]���5@Eˊ��`s'�'��3�D��nm�</.��cD�,L��X�>��oojy�i<s�8�2㱈m����mg��D+�s��<~�����P{n��i��4�T]��M_��O#�i�YWu�����~�n�)%0Ϟ�+l��~t�����s�cyT��g�)��A���sr��$��O�_a�5r�P:Ixf��%��_��pj�Hv/��	�&g^ţ���-�7����?�p��p��,�3���>��dhs�I�G�ͪ��a�Js�ۥ�X�˿Z\�U���Q9�xè_Y1Z(��@�]�¶�a�=���kv]�w.��~�ν̐=��\��jyr�rƼ��ӊ(H�yôI����z��G��K��68�/:���X�������-�{;F"�Ӗz�-��O�h	��km����q��]{�������Hi�P�UC����Z~T�6,v���y�R����I����������d�C�9S��5������~�ݥ׹���P�hK_D��LB�[�O�sAH�`T6��N����������/|:E�\ܴ�2�����ta�(W8�����f��=t���9'�7Ҭ�M�;�����2ש��ɾfV���+�z%փX��܎�R���?��F.J�Y�G�y]W�c=�3�M:��j��hz�μK����R�N٫X�5�x{Ab���\�kz��,����o������09��
�y!.�����B~^�ώ�"���v-1]Yت�./^�[`�`l4*#*����*��p�K�f����ub	��Qu��nxK�<.� ����v��Q	���l}�g� �������'�xJ~���O�nY���
�;}5p{M2���c����h�Z,�W��g@S�?��҄\��l|���MV]U�ܥ	��t��l��zwQ�V+�*�П����K��g�g�u[�U��߱n�y+ۋ	+/ҏi��%��=4�w�pci���F��v�$���sx)ned��m�v=Mg;����B	]d�d��o(iqGcᚺ�Z���8�c2��[5-i��tS/�O�灪�Z��|G��Kh�@��v�J� ��<oLJ�*iW䕘��f����������?�Ou�2��`o�N.��O����WU���3��ʋ|�ºD�#9^eۂ��eN��0�l�^M����� �T*�F=qL�§���Y�9�r�ۯp��R�f�}8�SV��3q�!�\6�<��j��=��!�.=�[��hT��l��I=���Ձ7�w2��֏�md��1��H�6Ǵ}��ÿ�.��íP�75�j��ɛ7�T?V��:� �]�*�[Ƨ̱�+O�C�lI[41�U�Ʊ�g.�B����{~�ޛ�~�Yʎ���7��C���f�x��V�{<�Ɩ9y���#ݛ�:�k�;z*���䅮})x���T�ʫHig��l����Z���JOf5o���Zt�Y�����#}���K���7v���U2b�3E�2~�z`��|���]\+��ڨY�fSe��V�1ۓ��O��"�g�b�G �s��ϖ�|h
#����E�{��OK{�6�L�av��ƯNV���=(?s�s���)��Qm��sCIe{2T����yf&A��g^��6n���LO�����L�zqVP��/*�c���d�������ov��������+e�4���-�����n�j�K���<��Nj�Ŀ���g���2W�� 1���B}˷D~wQ�}���(ȶ�m׈���+�R��I�U�y*^��C����ߴ&Sȋ��3���KmO%��ɩ=	���5�j�ˡ���V�x<j�:���fOm�fVҋq̣yD=�qg'� ��@X�z��%�י��f��a��iEV=�l� /��|;+����1�:�3L�^�����<��^˘*Wyb6.��f˪�ޔ����>f��l�/:�Ŝ����ձ�8��m�s��[�&�W��s>�^��N���}x��J���o�7�',���-�vw2�Z�S�f�5�:���{��G�[txf��yxR�>~�筭62�=��7��w����X��|%S��V+]��)�Ҕ�i��5pנ:�>Mm�L!@+�*��kumވ2�p��iLփ�d���Hά��Ρ`��h����;�ֽ^H-��4/ma�C%M ���8���щC5]A�,�@��r��¼'ͭ�0�N}�!�-��>�T�gy����k��F�X���r�mu$Y���k�\�xEӸ{"�9M��+F��#ֳ�����tv�e(.�+{��M<_��m��,�#
C)K�zN��f�1#��+�0c��G$����Є�ռr�s��S�Q2�f��B���Ug��W�Q���҇��)|���~Џc��E�*���5�,�އw�����1���$��a�@~]r!'Y"�x�Ζj`{�`������F�<��v����4s������߽�:{W�!�o��I�X�t #&�"|���MR�"�tC��y�����^��w�2����!,�T�q�H����Z��c̘�5&.6��U��٥u�`�3gN~��noj>���THC �H_��z˔k�������q�0p�K;��ߧ�y�R�6��cqOM?u�~�#�eR���]��R�+�>g�y;|,0h)������ͬ�)6�2k̝[��&���20�&jb�{>���$�.Cң2C^_V���WJ���Z���;���ԕI�w��}����G���`W	��'}�u���w���6���:W��>c/\]���/�^=�Μq��Q���y�f���O۾�����>�(��6�ϼ���[��[�����O{u����Y7Cd�Ɲ��O�O�#�"��^��ܞ�n��;�:߁�"�1=<4d���U��9���4G�9��OxZ(I0A��X�<�s$�f���p�V����(b��[��xA��a�kP�r��˷J[ŧ-������}�nCx�u�7��/��%-�]���l�AɃē��f]�zf����J6���5ٜ�������,�U�\��S�b<LS�\���^^t��s��ӱga�8���g��L�;���'�\�^����_ye]�ogǆ�7��Tҽ2� +�ZC�e����$Z�+'��{y�8�پm�o�K�ۦ|�o�;�x�Z�OJ���U�8��T�^œ�O�tM�)����y�t@�TG7*�ڧ:�糇�+�)���]�+W���,�1(:�z�������s=�i�+�0�`����Z��s��CU�*u����;��nc�MJ!�{�Ei���!�-�v.R;[�4'[���U��z��d~����6�q�ZoS��*v��{z�>�.�\b��g���Ъ�}�՟��}��Z@m{�?W4s4#VD��uA=iR��.=F������8:'A¨Wl�GT/���p�cDϔ
����y��vP��	��^]ro��i��n���(��h���Y��.�^�/kE��}���׽⬈�
D��"�p? rf���a��Z��IC.�c�6�x�8�{��menJ�͏1^lw�nI�{vrP�qzj��tsڇX�45��oQ�/+mj>��Ao�h{W�&��Ϙ�����Cۜ'�?�^��6�g?JןLbE�E�qUb���+�Dt;�ˆ�vw+��*�Z��)c��l�i4K`i��{в�v�lCd�Z��N�F��+���Y�S�/~I��eF�f`��l\����:�*����F|v�_yf�+u�P}>��\#�S�(��DhX*����^�O鞧��5�~�1��ub��`<[:ϼ>�P�l���M�6�Z��|=5�~R�dܯ�p����*�+��#u�1���~�������y� }���G�g�&��?�-�:��;+��g��X<3V��yT��f'`p��һBR�K����|��S�W�ka��	̞O���
O�aY\@��c�+��W��+uTݖ�u��<P���À�K�̆��׮�<�X�nǾ�k���`Uu�}3���ץ@[��к9ʿM8{S>b�|�9LF��Y{6��י�I�J�%r�n +]��z�g�>��scE��#�4��Q��W���3��!�\Cj�͆}���ÒPm�"���3�"�mg)8�w�]����
��>����o>^�2]�<!
�Bua��#Db>gF���Y�k��A�n���x��1w��5)�=�=_g��
��Mz����B��e�|w{AVe|7�UI���������9\(�Ao����@b
��:��1]��������fQ��t�+f��K�+ro
�y������A�W7�
��7R�lC�'&��G8��m����T�)f�K��@������O���ogQ����mO_[����߷<o��L"�aMe�z"�(A�TV��b�ln�Sf�VM��np]��ȸ�.w��o	AZs�����Z�]�/RjL���E�;%�<��4���w�[���մw:H������Fح953N��1���*��>ҾÈܠ�n�7׮��'!C��YN[x�d�
����A幰��@)B�ۼ�}f�j�$]�REWC�N���e�~���s�H�'4A=���v�\N�V����S���(� =���	�9񽖰4�����j�Cc��lf�-����%�l۽1�Z��Q"��fҜ]%u�軆�U�pҶ�֋�<�k*@�U�X�%��1`�Y��	=��w��Q4S��)Ԕ�l��<5ڭ��8�Glr0�:v,ol4>ݮ�Q��1�����.���+�;���V�L���Q��wҢ���{h�ԭ��kA��k{yR��ـd��H7��Q���;��V�����M�qW"�u��+6a��sSh,iK4������Β
#���U���R��ƌ��9�Y0��W���f�J�mD���Y�ښ�w�$�gmO�r3.Ɋt&�(}}��X�9n���]tx��q%],�3�)y}}��L<�� �;r�t��z�9P�zQy�2�{�9�lW:��V�tSM_V>ۆ�c �qr�����i�|:�p.|3��|}�_��,��أQ��f7n���]��3�]���b�d;�����E�y�Jz��i��+��S�2C�o��\W_t�먐Y�S�V���ˏ,Y��yB�壱��k���&��%8mM�S?6������.��W|�[�J#��.�!�ھ�L*5 �ڰr�n�M���V.��m�꾩�����s�nc�GQ4����>p�-�7_T��C�^�u���5�RGb�gjP<�Mй2�E�݊�p�I=�;���+���J�+Q���χ t3��A�5�Z��K�ھr�����	��,�H�u]m�.��>��KfH2���ڰ����U̧�A�xuiճ
���sr���=�n�kN�e����L���Tg�UD�#���`������'�����Ј���-YZ��`�=�h��VL�<�kގ�T,%��8���:��D}���]tT,1F�,�މԽC7�)9��V�Ɉ�� X+��n����S@�C��6脣A9��`�[Z8�]=6_Qr|�.����7���6�U�h���5���;P�B�o8=��g�v���Lu�\~��h�z�p7Hˢ-�7��70pp7��?�f\(�ȩR��rME�K�yJ�+�YYQU�t�9UAr*(����L�6��@J�ft�E+��9��R���1�,��F�HI{I�\�J]B3dU&��^s��J҈�W"(�D+H�-l�¢��N�p%r����Q��*
�`J�D��Ӓ�\�(���2�9):�G*T��ep��AJ�H�g�Q��l�8D2
"�ƪ����E�i�F��.Y���V��"�I.��*9r��;"R%K9W(+�L���D\�Y�9L��4�%H�QF��\�^2�G9E
�\�	GG3N��&r��`D\��D��)�Բ�2�eëJ��B��K�ۏ*����,�+$��DEI��B&C�9�*���Us��\Ib+:��Dp�8<Q����J��Qe �PB��񗔪Zl҈�
�E�Tr��r��(+�TDsD�dW"�TQ�[pr{�p���/n�M���ݍvIۚF��0��
&�w����,X�7��D�٭%���ڱ��XRm�}݊T�}@|���K�P���8�U?{c����&��9[.�����p�I��G���@�C����=v�s�`�o�^G�o�n?�Nx�w���}{w�i>_�t3��9g�ƥ,}���FL9���0fS{���o�O�n';��{1ێ�_m�߼����]�s�b��|I�#��2o|���,�^:O>����y���ӼO�8���W=I]�4��\ ^�~�@��&�j�w�&#�D�w�p��8�{޹�v��-�o���hRw��)��S!$������N:O���;M���a�n;J�����z��+� ����0�������s��~�Ξ���xV���HX�;���|�bN&q���q	��ϼ��ޡ��q��[z�8�I����pݠ}I	��{�/��M;�.��5�Ӄ���ݸ��q�pqߞ]�}�y����T�g�?|'�1�1X#�7�z���.����N=C��}��t�]돻��;qۺN&��9�����۞�.����y�h���?��s�s�$���������|�J����ªޥ��
b����ڌz`�7��\|�9�qۉ�����G�o���N�z�~;z�T>����!?�>wÿ�����}���~��aw�����u��$��y��P=d�����<~�sV<�}������'��&y�4}�$����>�n�:q�ϑ�q�+�8���q�&c��t�~!���ĝ���!��v��N�����39����M���O�)�o}���R��T������h�+����WySA�һs�s�|��+�~�~�����a��p;�c���!��z��0��x�=������0����q7�$�7Ps�ޡ��!�@�'�?����O���3�ضgnw3/�ⴞ���LD)�1�n���{��iS_/\��ޱێ����>}��t��iߓ�{���}�J���:M��<M�����`����ݞ���O������|N�v��Ǯ�.���s��)B���-^ꙟ�����}=�s���� q'o���|�ۈ�u����	S�i?�8��ޡ|������'
v|��'i�۷���|��@}N�;x�T���M�*��T~���֯װ��ꊝ~�VlݍͥzeN�%1�%aV��WoRy���|c9z�n�_c��(X|��A��P��A;6ue���A���U��=��dFZ�79�,�+LL�7�����d�tgPL=�|�.�#۷��zȷ*s��^�h^=@�n����_����18���㯖ݿS���q�U��I�������΃��X:�<���8��O}���'n��8���'h���|y�?\~C����`�|\>�(}�}Һ����K�x��M�߆���'����󏩼���$��~��:���o���'m����m��X����w�o}O�'�y�������#\��o��owz��>��}@߸�o�Hv{�ב����?�ι�@�'����t~|v�ԓ�w&����vut�Hz��x��Gn:q;��X�w��#n��q�
���VNw���U��C�W�+ӟx_��P����{���S�0���~�}N�t����s��(��<w��L>[.����_ q$'}w��n;};�N�x��]���n��7�/ �<�0�^�x<�m4�GDF��S�	�;�s~I=v�㾸��t�ğ�ާ<����I���Oyc���N<~���[t�� |�8�ڭ�Ğ����~�y�����N?{c�<�ߞ��߇�ė���W<�?��t/�to�˯��_$�Đ�xn��>��o�[��&_P��y�=N����~=��]��:Iߓ��y���n'~GIӷy����$޾=;�-���W�����O���?����G��c��#�3��=1�1�MAX9����!��q0��>{n������:�I��&�	?��u�7�q8���}���q'�׼ݧ��n t�<b*c�?D	��xl�sL�/J�Ϟ��q&�����Ӊ��=�p�L.����q�s�bwgv�M�x�����x�a��v��t�L/g�8z��8�N!�޸n�P�����s��'�L�yt�j��/[�����a�h~~��Oz��;�{շ���v��'~C�s��n��}B��P;qӉ��w�'��;��XP<I����xv�Sx����6�;�1;��89��3S1���I�7U��/v������~���:L.��{�1|���A߾s��c���y����;���s�t���#�n��>!����I��:wg��ĝ���=sv��U�3�ǉ��~���C1�g6E|���5�Ǥ^���&}I<68�n��*�g"���ʍ1��좯ޘgv�uqP�J�͵�%��Qn������3\f�v��g}7:r<p�qv�n�/��Hy��C�[���:;3��o2�]�q��N:;��+�Ք�g5�	�v�K20�6jb�{>���j!�}��ݕ���<�>f�X�sQ�W��E8y޴�q��G�5h�Ӿ���
��خ���[~hc�޹���vJ���~YY/p�>ɺ��:��RuCP/��T(ǵ�� -��~ٞ�s��7{(�x�Vl,ץ���U�^�wt�D]��D�`������UV�}�9Ɔ-�>zӓ�\����΋�AS�-z����Vt&}\j�nJ�v.qO�牊<G���:P3��Z�yh�Sz�/a.�xm����@�=��
ߗ�������k�Ӌ�'�Ŵ�L��
���<6}|��t�W�h����d�g�N|=��p���+99nſ W��c!�����:�V�����m�K*�0�ᩫe0me@���T�|^_���W�S�4詚�S�f��*a����FwM�x
(2Ϥ^>|�y�\7��0߶��'VÍ&c"�жr��U��ǅ�0P��.�Ƥ�S1tb\H���DL7���r��m��kf2j!��-�(OF��`�Ga��w�V@{=���mhn����3�u���T���E4��ÆQ+��M�K�&RJ�U��i�b9F�^TKLf��d�N=����(���ͻ�_;��ݝw��#��1�n����^��"��:l�74��Ԙ��,�:�꙳�
W�E��5.;�@��(�� ]��`��
�_j�d>���Z@/v����X��̷��W�W��JS�i�3z4=�, h"(�
��KDp����K��1��W��I���2z��|=�tn�{���M��Z�G�ߔ|%Q�4�Z-Ϯ�L����sR�o�p=/ޒ�`$?�hr'Ps>~@��B%�:~���Ld����}:f׋�Z���?���aP��1�0�3j���S<B�31��6.{Y��U	�������_z��w-�{���ޭ���E��ǘ�A�kӿk�53Թ���ߝ!��P0*%��⚶�C
��E�1��������_n6>��@$:�>{u��R{_�����]׉����FF0-ms�>����ؘ�{������n�ُ���=v}��n�N5~�4$��yJ{�fr��)!�]�s��{�Oɭ�}\)������<yRW=������[���%�.kq<�^��f\j8č)��q��T�\c/.˯'��)��uy=}�]���!�� n>.��.i\��e{nhe��˂�ܫ�9K\�i�k����F���=���x��[w�cMּ��Ȫ{jY�}��#���zλR���w(;�ˢ��K�3�5ԫ|��N�l{�%�d5��u�˶JDf�zZn��%`R��d��u�+�B�8CtrU㩓F��*r��9s��fY�{f�>9� �۪�c'�NY�����+�O�4�
#�x��_���"�3q>b��ڸs,^��8rJ�⬞�Łn��M�G�+��8�e�D�1tLkC�Uf*LG�W�1"����h\�Ѓչ^Mβ�o7ӷ�g�F�ʿR}+��
� �q�io���>z����H��z�.�y���o��ozR�|~}�G�q7��043���Y^��X�̭7]y��{�����&b��Q9JlaHCb2|Cn��ӷ�7�2�^�@{��Hit{Z�k���U;�`ZL����/�,�?\B�h~�DiU��
�r&�b=2b�rB%��f��?n��77/����jk.8�c!!<6��� ,�y�����ݿzՁ� 
��8<���=峅vQ��1�/u�M!��,�a�ڻ�[�H[TDWק�$\N?BS��\sM\�n�s�:@��ތ�����p��|�ƥV�8J�<�{�.���u\�@i�+˩��U�]�J7X�0>ܮ��>�G�@��8��{K��
n���<�۹��F2b)j������q�S%�o@��gK�[�xJ��Z��t�wׇ�Y��#��g�Lt1ࡥ������;|{�@/S%F�7��Y\��d���޴k�ٮ��W�1�=��.�BEk��k�MUٮ��|<5\8yY�~��3/r�����_�Ǜ��q�00o��+�����Y�*��1|�E`��3�"41�0�N�y�=:V��G:��v�M���z#ь��˯Lbg���,g�Ϋ����[؛a ����P��aЈ�+�b%`c�&��)�7*��cuwQ{�薹=)�&�������{��\hg����ʧ���xm�txg��=�uK��U�R���5��={7}sX�Ͼ}�Ҽ���(T��!��+]_�R�wt�9W��F��#w�N���
Ȥ��G��i��
����p]4���%�q��fc�1�g�V`sT|e]<��VTÏ2���,>U�����U>�:���Q�"��J8��ip�	����<��]c����,ճ��ʹ��/F-"|x`O�c�JV��_  ���*=������)K�r�s��M���t_����0`
a�ZN�C�Fp�SD 6T5Z8���=��ٻK�@x{e��Z߯W��
QX�rb@����f��RnV4�����x�)�3Ցg�df��G�L�ɔ-�W/�@�k�Wf}{x_�!ڵI*�^^�vU:ձ�ܻ���I/��BTx�t�
Zj�*�7[�OS��к��?/��x�@}ڧׁWg����	�[�w�7ט2�`hд^j�o|�^����Ł�r���pS�g�_��%R�dEj{a�C&#΃�D�f%��z����qN�+��W��g����y��l���T{���w���{�w�l�8��j��)�p��f%�ޯ����?��s�ϗFG��Lh�P0���)�j>�)���u�͗-d����wꠥ`3��R��
\��_6jb�z-����N����+KvW�+�C�xqa^,�}��t�x����	@�Yu3�SqUNN�'�߯��l1�Ѯ=+�V#r��ؼ\� ���k���h��LU<�Pg0,�����]D���eƑdt�����|�������ȷ��LF����Ճ�ʵ��Y��U��q~��Z{�tb?G'6P���q�5b�'��s�>,O�&)�R��G�����ɍ��b��-4�M�h��˔�UV���,ܼ����OY��;~�����},]SJ���
�i��{��XM��=Lcq��\f�&e�����] >��B%7,nߥ>k�r�MA��m�G[-Rpi��#�)���ĕ���x�v�t�͵�T}��4]�Q"�r�S���w���RV�']���ڤ���v]Kץ8��Ҷ�v�tظ���h�?���ty�~G܆)��<��F�4g�`�VM���� �k���"̊Ѱ���?�w!,!sz(�����	^T�}����h��<4������*��g�o�w�̱��Av[+�x܋G.L^yW�uڈ�:��B���>���k�]h�s{i��0���ݒ�2�P�t�!1�DƬ5b嫭��:�l�M?:��q�&����
V��c�j�Z��U-2�H
�P�5�a����9W�V��M��]]��N��x*��-�<z;3��E@v�£E�te�F
����BQv>�yԶG�*ܙ�on��n��j����S|����Bc�+�~:�ߙ��G����{R�V�w�dQ���bS/}ٳ�p�}�������|�>϶���h/s��j�za�36څլ����ї�j}�8��rZ��3�gAumW<�h����3����|ع_{Y�yT'�}�-�(o���*���sF�8 �֛�!�</�e[����uS=O��}��*"�U�w��y��紻U�i]��� "(`��Oڇ&]8�r��˫��'w+�L��p29Q޴�ً�$T�5�=	��'l˥�l͡�\��}��u®\��]A�k��qۋ;�����9I�.f���2�S\v�k�jY�f��U��qh�G�wb�-ه�0Q�<G,��.VM�\<���>��o�{_��6�Mn�gʑ�}��i]�Ζ4W�L]{�����\kp��Vo�|�Y�����رfg/k�ㅠ��c2��+�[�.��[G�}خD�@�S�^��_�ee�*�˗�TB9�1T���w���Å�gX�'�B,#R�1��k�S�π��m!���?T;�w�h�o�.����<�0�u
��;x�d�r*�)��ÜҲ�nu�!�R L̇;5;�if�C�i=U{�:��=qDʘ��s�\L^usQ�Rn|�9�m\9�/C�%�F���<����[vvM��H��c�f܈�ЃR��i����7�m��"ܧ�9��׆Ԭ��X��m�ޡ��}H���� �]�E�EЩh]i��I��-�����e�M<t0+x�%�V��꺴���k Y�t���Z��g1��..1��I�K�c{%��gl�^��ۣ9qNߠ���SQ�h\x��P�0������4O��9ve	����1�IfX6��݉P���0���Ir�k�]ig�O�[�*!I�*�G����Y����7Ȳ<.'������ӂ��݅�Y�,��f�u}7t.)i��$��䂶z���a��P+������I����꡻z�[�����Я��V��K
�ժ�:|��/��L����$"Y1����S/ �T_��o�
oެ���9X]��!��/>��}�0A��5��2�*dF��m�ل���s{n��ޓ�#�+��B���|���8�Wau��^���4�j��o������9}]����7��5+�Wk8@CD*�FG��{>5�l.7�O�:֭�}e�Y���^I'D��]ӵ-���>�׉��/�i�#-;������{��_á"���zګ��p�m�o��]	��b��fl�K�i�Uǧ7-k��}�L�~���/�Vs=�*$f��I�3S{(���^����Yz���k�3"�R���&�@�s�/�Ꞛ�3}�0T���l]��͐�q^�Ϫ+����xϫձN+�H�z2<I�X���*aˉT�=ߦ*#�VP�S���}(x�w8J�ǔ^��* l��7|k�����xn_:��<Poy�U�w�Q�d�V��yמ*N}SA�E-<�wܝ��(T�%�ս����_����Q�����xm]�HlT`���������$��0�Jw�pV_�8n;Y��z+kD�k�M�pW]L�ૌ�&� ��=x�BC�y���!4�1ƂV�=�H��g.�	o<9ޙ���s���ܾ7a��`Ѝ��h� ���|$��u�M��d�,�z=m���ж��i���&�����`�[�H�*�\.����͏Y	+��Gvo�s\�#8�{�k#���<4m4����v>y�ͩ���X��E�H��Jk;��ho�:&>X*k�(�Y�ط{Ό�;��kE#���5�8����.T��RR�,�y�V�ֆ�B�:Xqɓ/������1�{���:�3�!z�FKV�3Y.��pl��� ��ӱw`�	>Wj�������I�uۛ����zZ �Aʹݎ29�u���"zk#Wqpa��Q�$�����W(��{���/4B|�T&Õt��ȯ�g{/%����{�f��@��&��Q�
��k�yV=�.O.���{DfZe�W����xtk���EůU4�Y�iI�M�]�>F�a�
�h1I����>�=�p��4��]����O��Ѿ-��Y�}=s:Epd�Yx���a"�aPuɹB�piH��������c��=3Z%��ׯ��ل�����g+ݟe��,Ǖl�*5���R�(Vf���AZPU��wӆ�v�T����Kf�yq*����2�ʋ������a_+8lY��vHE⌤��i�7��I�g���v.M#�d�r���]^w7z�c�jt;�U7��5ץ��j�I��+�.ҩs����U��[978o��;<��/��|�^H��_�㙞U�R����uy4kö���j<���׌�1�&��J77CeM{�1uҺ��o2��V��)>��v�$;
��bi@���^{�7'������o{#˸#�P�ʴ��;�7L��v���dvڝd��ú�2���C*�_hM��+6}��Z�!L;,O��3�1��-q�ff�����P��y�;r��A��7��G�d��@�t=�V霞Hr:m�k-�%�Z��o)�5�P���.>]ק���>��71).u�{���u%(���Wb�֤���5�Z�͡�nӇ�H5�!�b�.�֜ҕjb"�#:�g���օ�u��[���s/�-m1H��7�7�՘�����k���U���.�%���CQ^��vΟ5�=8֡{��vp��6�q��^�ڵ��x��H5+t�l�5)<�wb����j�G��I��p�"�莝3����@��J�9qF��u�+	���Kڦc��dռ��Kb�q�h�q��Ec�����'��2�ܽ|��n�-���<p[�r\ufл�-k���h��87R��)���E�ajjւ�޴﯅*��[�蕀��l��w�w��ή���|7��!:W9�A���R(�T>�9(S�Aʀ�*"��UEDQP��Iʪ��YU��f���r�&kC�T��e��QZ�A�2�*��eQU� *�L�0���tZ�E��+B3*�$r(����DjEUD�9S���.�$^�D8���P*�b�9U\�9PA��T$mL�Z�A]2*�dp��W�H���	ȑ���"+2�r4.����b�S�f\��AR�%Es�����G�;9�r�PJ�AvJZʥ�e2���gTj���I�HfEE�DE�TeEQws�J,�AQr(/W
Ta�[������dz�pE�UE�*R*���*"L(�\M�\*(��d�W(��5"�ND�t�hТfap�2��,�5dDj\�D8��VeS�+�U�<�M��*��[F�B@DQJ�R�
��T**"�eEr���U�̕��?�*�
u�c�
;Bd������ BzP)`��ˌ&�UR�������"룢�7���9oz�l"��a�"��; w�_W�UU^DY�wˣ���Z���w�
�mL��T�d%�=8։��������a��ΈꜼ�G~G�)�����m�v����^�k�ޝ�~�f����U��Ӣ�|y�����cy���󯟐�|꒸����ڪ,�����ee��S�4�QY�b̏�����eD�?\$�_��e��)�b#U��z�h2w�����^��|1���E�Q�<͗��ۗ�o#f(����>�����ڠޤ�n������\Xk�Lߥ^`���R��aB��F��9�!g��*<�ݹ�
��$= �u�;��N���pஅ��坮��1��i^��Aô��BN1���}�G!��Vz|r�+����@���]��潋�\#KX��+N')��{>���j嫈1��q칚�2t�������T������*��x�Ǒcn#����񟍍��c$��(?A]h���/��1a�2���e -�5�ʇ�J��u��Lyf�e-sg�O%<���b�Kq�0�~�NN޴���Ւ-Q�_0�� 7+���ѷ�L�g�v�f�����ou7�h���r�Ml�#v ]��F&����)i�O6��K�����ﾪ�����l���%��@{Ʊ&"���U>��Ԟ~/��񆲏7��z�Xf�����>�F?.O�3f�4l���;Q�-d��x�u[���[.�ڴD��;����'=��5{�B�ұ��C��T=�8�����l��T
�t�j��i�O��ꧏ�gޜ:�9���{k�z���|E�W|�2��	,��v�	4���{o�u�s���v��� +��ҹ������1���-�yѴ�^A��^�z��5�پ��]H�P���.=��='����^�V������a�{��k�P^���9?cKzY�P�"�O9���>�i�Y~u�fxm�{G}�6������o9C�$�C{�2߼�X|��`��d*������|�,��n�p��࿏��u��7v�}��|Rq3�Q�o"�;b��HU�5~�%�"�
��y%{�"���μ��+���m����5*�i1t��(���(�H�;ʷ�[Ɛȋ��s9V֣u����O�k��8�z��>��y��}Q݂����o����|�_�w.99Pc�ˠ��z��Z�;OkqD�B��{!W� ]����S�P�������9��m�g����<2�5��r��z>n��4�蕮NlKѵu�woE�[v�aU��\�R�	��YKҎ��crr#S�v����_�[j^��yf��� )}��]�Sy�:��cW������L�1�R�<�c�?'Ì\=�&N����x�
HJ�/3T��f��Ǒ~���<5,D&_��q+���ޮe�yXϼ͉�x7�=�����w�叶Wi�gcΌ���U;=G�n��3ڽ�M{��e���h#�o�w��o���vI_�Z���S߆��^5�8���2�=�6kؖ׆vmbŗ�W��}����j�<=�)g���^��N�Z?g��ыk�\�؄}�@ڊ��/�i�W�^�,[��mgW��Λ��I���w�{�j��=1i�؛�ӪjG��j˳��xg!{ �ݢDϢ�B��x�~#0lL�v��G|��=b�Fj��%�0�z�8� �	�Ã$5��j��f৅������f�B[�i�Y�
��u1�h�z�H���?��1��?>�sǱA�s�[��	P�7.J�-裝P^�3Q��S���@��1�39�m�Cg�G�}�Բ�����kKkߢw�S/bPp�\��7}��5�U��q�cʘ44��6������y��'M�Ӗ}k�Tʬ���>��.s��c�-�k��i�ޜ�O�Ʈ�ϕ/1��
��uk�Uf6Q��x?o��ו�ĤY�آ�˓,�I������m���D�MT��/wb�Kt*="&���Rh��1v�})m_����Wѡ�C�U���X�y���,�^��Ա�)ݜܾr���{꿭3�G��؜�Aǚ����6����;�����J��?������@�A�j�z��y�"��W����Ƨ7��b�1�'�uI�ſ{֫>�q=���c��U}����7�r2�%{#^����U���E�cg*�U=�����~?bKk9Z�;i�F����G���tY꘽���?����x��x�}�����1a6���,žX �XbR0�^u�"J4��~����B�D��;�#�:y�_�+��A�WB���6���V����o�f!<�jȹ|[�v�J��]:�y�ڸ8�O�>���M=Ej]�ē;H��S���w|�V��C�j���������wCǾm�/��ϫ����qFD~m���f�^e3�y���y��{�Y/neM:��{����͟��~��q�����׼c}KOq}�����륩�g�!���N�gަ
5��СnG����ֱ��S>�*˯[z���
r����>�q�6�~:�L��mS����*5zwm������ԻL"P��|�4���w���Շ�w�
�S*�Ppb�~�!���}��w�	��}����Q�yv�_Zŗ[w9��ڪPpb��B@�9���&Ө��O-,���	m�SunR}���-{~�ණ۽�����}9c��q����ົ�B�!=���c���Yګ����r����B�R�=	�]��X��[y�8[�:��^-`���~*�>^o`�5�z����a=�~�T�a�zؔ�2��nK�E�%?_��xg+M*f��q���/���b�!'0psN֊��)��a"W���tM.�ζ�r��;��k�����zen�si�܌�-�>��g�Ȯ�n����__�.&ߋ��Ph-ɡŎ$�cE��˛��E�VE�ٽ !S��z�LDK0u֢5-3��%F3��}�}_}T	���R~�\��bR�E�s_LTF�� r�`#���"צ��iv_��8	8����g�;�KҸT=�Ajب
��q�]Ԡ�Q�V��l�>qַ�R�󸑓��-���4����C��T=��Z��?b�����VYnt�ި�����Խb��+O�V����"��߸�Gu��u�����b��ߣ]�K���^�I�yZ��|״/MF�ǌ?b~�3*}N�'<71��b~���W�D���7����L�Èw��]�IǊ/�ST��UlRztM�溡�:^<�����!�*���%��A��}Y�N��W�����jj�+�8�J>)�N�?!=�w���ޱ�V�]Y+O�ꃚ�,x�Up"�B�&��z��/e|�p�Jej*6�+@G�Yr׌�^Y��z�������i!K�y����.�28���d�~(���jV���Vֱ����]CN�+2 D�d��vڒ�L�[���\_>��������C�x���*����*:!��f�أ�Y8�F��\k�<�`���	�G��RL�+P�KL�Ec� �T<%�Ωx�o3!j;ٳ������v�ޛ��V����pt/���J��U��6��&ڼ�S��y�߄9�v�{�Al�����|�ߏ���9+*��e��s���mdoj��C8��kك�R�A��i�l��2��B�!կ�����z�?Y����������Ω=}gRs\X�ט�M|�Ƞ튄HU��W2��ly��_]�X�槧�e"�^��Ӫ�.��nܠY��+n��n�	��֫p�,�jkCߪ���(�����95�c�=f�ڿ�+m�+go[�Kg�;�vϾ�i�yf�X�{~~�����z���=�EW��U#�zwv���@�{��4�߳��~Hg�<��W%J�5�����f���Ԧ=��(��c+�؞��*�'��֮��/8��V�h�)�C���u_����x9K����G�PIײ�p�7-���{���g�,���G�\��'\�)���g��;f���Y_�\�I�%�r��K�.��e�4��,�F��c��V�Aᶖ��>�e,�����#�Gi���?�V�9�ne�V�nL��̲t���#J17#��v�=Iخi�c5 ���ʾ�#���ǽa��cڎ��Hc����۷��޼����gި`�]E��϶�dp�F��po�S�꘺���m�\@T����b���W:���.�No��w�U׭�8��S~G�@_���5����	4����fՇ�6�۴Q������w=����V7��N:&��tb�B�y����swt����)[XR�(���Nx6��Cc����D�5�;k&��)����t����#g�&�یr�y2��XV�լ�1/ ͮ��W�hz�˹"jǶyƽU�Ӌ׻6�y�W��	��-}���l,�ޫ�-a�����-H�o��|���u}�ו|Vf�Ɨ�g��=�]1H��2�u�@l���z���u,��Uz_��j/ҏ��%Zr��A�퀳�����V���>���2��6m�AtZh�����I���p�/l�ؽ��3��&�����Պ� �VK��:�;��.���7nן�ݠ�ǲ�u�g&E#��w���D�M��+�v�|�7�>�j�t�=:*w�b�J8MgJZ�sCt[1��L� ���gN��L�����p`�»/��P������yֱ�h����}��}Wɐ������W���o���1����{rq��}�Q� ���.js}�Ϩ�Mi1���Q�ȿ=�Ah���7�@��A��������C���z�r��٧�O��x�
�T�6=�J��@eW�؛^��K%⣝�k�-}��<'����ر��'��xx9T�_��U{�	eĖ<�Os[|��~ƇJ^x�Ϗ��6v�s���V�QP5��{���_y��X7���O���U���<Yd_�3g�1�c�C͏(E���N�� *~�!w4��7w���w��0'K
ur�a�z�(�
o��(��4��{�[�z%縍�sۣ�H�U�ͤߎ���ʤmS�Ƚ��W�v�'��t��)���%� f�{�����,,��ʤT�%]	������������^�ϡ�����w#���>P����,����ꑺU�mXų	�zz�R��U2�U�Jվb��kͼ]Oun1���&��^�r��]V����ɔc�QV��Qz����G�&a�s�=zL���_����,�i��z�߄r��/2v���ڋ�,�&]��{��M�����is�H�%)XX��}U���n�H���a��R��U���<�|�!�S�J����9�<��{k�����1
4�z�xm\�����_/#]�w������1-��d�7^�K�=_'�Ub6�kKZ�__�V�`��~�4t/q��N�gT�/Cب����+n�2�M�+{�E_[k����P�4��x�����s�8�C�a�sP1_i!���DJ�b��g���p=����b�����T, �^�)8�R-|�}歊
���Ƽ��0M��/٪Ӭ��{||i�|_W���[��_zZ����j̞��:.nYg{�v��� ���nr����W���Ǖ��8��s�Lv%������R����wb��r�w��W�q'��k~]C����ܞ^XĽ���^G=�]x��/NW��>3j��'��7�z�I����5�}Fv�+��*��\���4��9�ˣxs��=�C,�s��Ĵ�����V�Um4�Q�v�/����h1:��k��=��z'lG�S�ä�5�E|ۼ�d>�YuaCF��U�i���umv��]�Z���U���v���4rxP�M���&ޫ�5�JX�wZ�3�S�9�/dn �HȬk��rZv�����:�R�Әn�2֧��ގ�)�W�h�x;��><��1>��W���v�Q^)��qA�챬W8k�]�r6���6�S;7u-�x{�2��=�t��KM�L�K����rt��Q���J�}�����Ko2mF��.�&��_: �ImG2��mw�!Nk��|�����=Q�e��wV�kN[�
���;�uЋ���v���p��9�D�wy����x�xmHo�=�����"���+iܗ; �.�^':����6��|�ȶ7�pZ�%�'���=gN��Ul�6�Y��: �;�q�7+�hX���B��ղ'V��̮�x�Y�(Ch�%e�
�GO*�X
УB��b�{����WG����Q�y��	�޻\���95<��s�á;0.2�ۯ�6	��x�V٧;�!�,��M����cRXʫ�(�u�n�|06�=�t·�8@2g!��A���!���j��b��i�uvbs䖕��v(�r��N���6pt�]�����c��j�&�E9� ��L�F՚�QB�Q'�x��#ӎm�
��/lk���!YXg��l-4d��r�f�C/���U�N:]6]�Qʏ6�q�A���Ԯہ�� m\�����:=.�.�t��D]	�w�}���3y4���!�ŀ���9���Ki:�����;�J�.j�י���)�}�i+`��ނ����t���{U������xS�zx����\,)ۦ
�$Ǯ���+�����wh�C}�}�l�d΃
:-��^�h����$̱���9zJԷ��&�/�e[�th3&���;�k���gS����[�6L�C�\����J��NrX7��$�ˍ�'�]�]��zBƫ�t�))Н�8�ੋp�y1Z۵��ٸ�v�n�j��of��w��\	w=<0c��,���-.���i�av��E�KX�5",�ע�w���&�st2s�Uq���Y��*��S��2wm�6��HZY�
����*�T5�����T�H&��iIc�F��[��	�p���{f�4�~#m��=�G}�M=ɭ����sq���L��3�+�(�;L6U]^�KK<�PW!�U�;J�EZ/��}`X��z�ćm��u�H;�Ŵt�������ꊂ5��n�6z}�ڸ٥���1���*S}�/�>��m��?u����͘8� ���I� 6{4�Wo̕x��;��E]Ŗ�9{6R�<9Dz��Ebw�B�5X!pΉ	�|:���~�eʡ�\��T+0�]$�(3#�Ȫ��j�D���]�T�9��L�D�u�Kąr�F��U��Q�f�*���й�+�Ӝ�0�r� �ҽ$��9Õ��Y&������ȅ�T\���Qfd�h�Y�W(�D�kH1i8�"<�E%$%EY%�aUEPE�e2�Ԋ
��I����D�\��jJU��+��8�r'�er�ftȕZ�墮<B���2e���B�3T*&ru���i�-�%LBN��r"���13�(��Q�r()Q�AjR���J����P�P�u�A^/9+ȕp*�"�i�:%EE��+��F`D�E�Z-!uiAx�D��O
�"��UF�Q�d�Q ��r�U�ZUP��r�b�$G(�9q�A�+�d$� �K')T��!Wn3��1R��R�N�:�Er*�PD*+"8��TL����DwA�s���ɬ��֎��a�Ǻ�Y��0��c��3���ӹ8��U+��a��D	��wx�a��oi��G��舏���nO��e�~UB��o�ڿ8��ߗ��<U�5�K|3�kM����􈇉x͛��3+����P�~��C�חU��u������s�9��� jL�Y"�&��:<��6�ה���I�a���/eB����jeG�l�VO�),T|_y���^��k��3ӎ��^t~��^A�[O/����[R\�n��<�!'���Aq�gi���<�N�'5}�q{�K>Ѣ�)3��py�EM��;Ԧ�hv��i�Y����W9��<���-�K���V�3�R�^�{�����*!�����VA�X*Z�11{+5N�3Gmd
)��+{Hn&��9����D�_k���xF�z9��{te�J��u>3��/�\ʤ�g�y��[�p���sgD��>BKq9t=�����Y�z��`S�w�/_D���u8�ߐ���ǯ�0���"�k;:�;�iS�Oq��5�z�zQ�3�>M��I�zf�yJ�=���]����5��TT~�I6(l&,�:���
�Y}�-)WF���n���͗�p�f�T���Չ(;�a)�_:�E���}:�y���P%�3g��諭��[���mno�|6�����޲ߍG���*�A��C���iR^���^����Zk-VWx��^�~��^ߤHr�?$3������)bWu���T>���%w�{���c�l>��q'���o˼����WXܛY��%�9d�/f��)��O?���x��x�~�&_{,�p�	Vy�b�;Y�� ��GK��\�"�o�b���y��z�f%�1���Cٯ��1��y�g��.��*�yƟ(�Pժ�
���ڶ��1�5z���v�Q�����>�Kk�<�6����u�������I|�䓵d��~�wb�t�{���.��\ˠU�_��ng��I���T{�m�Tc9$gR: ^��-Ya�\e��ڙu�1���`�������E;��8�]�����ڼ�-���}_'M�PY������\Z*K�~�z��n�����a��1GA���q��%�	֫��m��)-�w�TȮ��[W_c�ӭ*��R_yzL���@��@�H<�}�t�Dl�g���F��e%;���l`Νi�T�F�h;�#��LR�op�Qge]N_�������ֳ:��N9�����o�F�����.���!��Uǯ{h!:�6ߒZ���V�=̋�:��ʍ��m��.�������f�z���KoecB4��`[�S�M*��ߠ�5�z���:���/T�oZ�P{�m-��X�%nB���_m�;ʯ-�UU�xs��=wE��d������k��c��-������i�� c��o�������bcz �٨����Mx�t�1I8�qT=�Aj�?5r����d��欭�e;u朙Ǽgr|�z�U���!_E�c/��SSꯞ�\��x7�t����	�<���=�N��I�ʠ�ړ��W������≯r.yuٛzѯ�zq�˽��8����>�V���xy8�d)k�z��^;��~�_qFR���]�-�:�5u�;�~}[T'w���{P�b�����{F�'n�'���D�@o��oڳ�z_�w��rxb��\��ϕu{�:�6��Ґr�4������O��nfz��m�Z�m'ާ�UЈ��7.���j�Y{���؝2�iܬf�U���q�VJ��#���}�����_xZ����+��n{꯾���泃���R��g鮯��*�b[᝛X���yϗR"rF�w���÷i]�M;
��|�m|����Ӏ�U�s��z�3Z��n�W�����Z��k+���6��==�o�m���J�!�L�{cH��K����=����ސ����P��h��w�ݰ#���mu��f�{��
��Qn{ƷgnMϓ�F���mypL���;K"U�m5��̵��o���5_Y�1/>�b5{`�7ޅn���q�%��c�QU{�]-x|��"F�%�*��-`�kj/ҌG�e�s��ƨN�ȸ�fL�cy(�x=�P�ȯ��* "�@�}xT��@�ͭ�x�h�W;-��B���ys���d��y�!�-ۚ
��$=�TJ�����>[�˻��4�q�{w�Wo�;U�A����N1� }Og�~h�h�E� �.����\��jy�G�ݴ7"�g�m�r������[@r:3���ȇ+r룛ݼ�Q��T|�K�a�k6Ʒ��Vu6oR�ﻪ�<���)nZ��qw����w�:{��ΐh=M����ʺyѧq�e��7*N)�O�
yr��UW���R���>���u���K~Ƚ��!�j����*�z��{ض�-m]��=�\���)�Ӎ��m�Y���y�Ly�]>���+ں������rmD��W�_[�]��������DyE�^������|��g�5�g�ϼ�n���9����Q?W��mW��p�	Vw�j�����F�k2�X�n(p5��5o7��|׎���&}�
5�n��>��2v3%�:�cż�|�}���U�?g�ꧏ�n��_B6�MC�ڇ���>>�V�*��{_y@�I
��w����<���s��*�8��ݫ.m��,b��{D�W�Utm$�~�m<��i3�=��)Z�5��kuc�㎧�x�]a��}n��Joy�j��[���fN��ӂ�y����7G�����moǾ�D�|�,������wH�3�Qr�1˾mjh�h�U7�UQy����v[�.O�˻�a�z��A2c��<F��N>�^|��jL޾E5��>k�����
.Wb&��c��Tz���y�/�R���q�Z�GC3�c�
����1���W�=?dۺ�º�N�T\�U}��U���s�}O���<�~c*�)2����؉Y&� ���d~^����˛/=�TQ�Z�4��zj!��P�H��5�k��'=%eH�������b�
�k��K���Fk�Ji�؄=ӟB4��Z�u3X��퓷����p�RAtZh�^�_E�>M9:�y�!��nY�pظ�K׹�SZ��96�fwp�����vs��ƕc#_W�܏Fp�>�,���:����Vz3�q�C@/l�^K�|�{�Q����YS��<�Y�;%A����{���Q??+�lM��o��I�՜�	Ϭk~����ӟ�o�b���<��<^/~��&�Ɇ�/_�a�gG$�uN�z�?(V����>qO�^e{�n���~��ضJs=�zqp?1�	Vz�ߗT����D��v�5U�s�x��yߺ�U��:�v�.�B�̶Nc'T%�w4�r��
K�m3[�s��&�'c���ۛy5�Ւ4��(�Y�bKs2��~�{H^�PPuu/=�̡pU��Jw	�q��:��M�.+�z�@��p��X�:X�;WoD��8���$pY-�O6~��������v癓�d���s��-��/b�:�!���i1I4�kNМ߽6��k̇�<�5�����M��v�UB6�0�"�9��M�{[�~���������N�y0��m<�����S-��%Z��I��&�Cg.�/����V-ϱ���[/-��e�9aU��W̨?KϮ�w�H�jv�J��Kn*�����^ݟ5�/>��
�2}k�B�����<�rv�����
�Y_]yQy�+P�zk����Nø�}�G��h�����GI���HT�A{�?�ޛ�W��^{�w�y���[��u�R|�ާ�
��lTxh�~���~����g��eE���H��L���>��u�۞�%/�U�{�+��l���+|; �5o_��H�-�ל��9��$wi_�Ih+!P���UzZ�����q�CT?�Jc�xa{���/YRU�dL��;wWot�)�ލt)O�����H�v��n�Vx|�<�ZY��T�w��H��`�ޯJ��[��c�\��yd�J��$���;�h��%�O����Ι:�OaF����N��}&��M�b��� g(f�ꯪ���x'�w�꾍�%}�N��}Qx�
�Le�6r���S� k��79�;�3���v����|���yZ]�.���'���g�?/��sp��E���ߥ�Ol�����s<��!�YT��>�VО^>�yŤ��=[�N�+x5���"}�}Ȯ� K�y~2���
�ݿ:��?J7�W��[`�~��o��{tb��o&��eG�ö�ҵ��0Q�>;_k��>�19NR�Q��_���_����*=r�x��D&�vݩ��/C���ډ�o��]f��5�j��w��U��B�O|Zj]���ڙ[���*�T�\^�zҋ������V���:'o�nUw#����ϝ��Ԉ塬k_�}/���y�[w���p\?��5>~�#S'V�����
9U�H�"��y�9k�΋��u�O}�EZ�vR�7�����w3*�_�^at����Y�������όAQL*�h�OI�F��R*�׈���3+���C��@��(�7�Q����1��L#3��٭K���u�4�ʏS3��T	�[�l^�8z�����lQ��k�Gz�v&V�3)+����Xww���������n[�����WY�<C�!T5�W1����������(�1�м��{�]�y��Nm9���sP�Ȩؠ�L��b4��6���Y���k�1Ԣ���5d��y��ݹ����IfF_�(c�p[I+�}����[~����[����$��~���0ձ�!���31{¬bNG���ùGl�~!��g.�\��Y����~����w�c���R�@�۹VG{7��\^�����39Z]�K7����1\�-�q�y͗[�K�`��ʎ�w�r+#�t��=y��}Q���!9�����n?h�<�����}�qS�zwޖn���_q�N�Emw��W)L������u/ۇ�&5���y��w�k�u_�c~����%�y�Ka�{�8\�*v�T����,�8��'�}��?x��F=j�e�0XB����̂`����� ��.v8�Bϴ]���U��DJ����RbJ����F$��/����,Ե޳+����t��5=�J��{�����e�\��������YJ0?�m�NÌ�u˙�N�����\�	x���}���}�P�4�U�3�xM/D���RH$�v��ٵ����кӔr�+5�Z����μ��aιH�i{z|����ͤ�B�"�7_�ġ�NW�Z�(����g���:��Xs����O��ܛZ'����`��X�����}=k��Q�w9���ڪ,��"���Քv�62����vZ袱��ƽ�=��5�욇�2��)2Z�����Y��7����{==o��=~��\(�Z�?{֮ry�H��#]��8v���UI��pn5˰`_���W�Y���y*��-�Sq���H���ؕ)V�E�w)[g�6m_A����|�,�rj58��[kޯ��7Uf?j�Pߦ��v�|6�m� r]��ڵ�J��E㖆,��Y���)�s̤=Ju[߻ط�KU��@�q�K��"C��������g2�ն�6f���.R��/M�y���U�����\��F;�Hof�﷘Q[<�nkR�[�ʍ�<K�-t1.��5�[�3������]xS#E�b��S>��wX��j�خ�+6��tnc��mcI3�w���@̎�vf��ҍƾS뺘M�cV��:'�0
b��t�KU*�GR �ӆF.n���{3r�ǖ9�W��O-i\sa�\��\2��7c0�A����ЭSE��)R�wNUڹB��f��bfjã�vVn��!�m�T�����|7W��w����a1�gg6��]���J2���(�?Z坱�U�9@��ǌ�u����b0�{����&�7�}���-��G����%MƁǙj
��Y�&�5a�e��z�4Rԗn���T��Y0�XGB��]^�yۭ�.��L�����'Op���1��cyFI�fr4z��^n�F�&���'%2����z㖩�2��e ���7��۶I-;�eY�P��OK���k��e�����[��j�ٖ�Y�m��cx�o��DxEC������ÿ%��y��"��c��׮N����q�{^N���;|pnVp-�#C=wN�;lD�SX�z��F�n_
Q�nb�5��( pV�j�{.�ێPWvL��w�j�ӳS/�1h�¸�}͠�i�C(S��J��ggM���J�� ���k�ō��9Ww��m(�����ڲŒy�o�w�aR���q�&*6F����z��i�lK&�\pݶ�S_(q��^��uoj ���I�]]��S�"1�D�R�e�
�s�q��li��T�a�{m��n!W\��p�k�,/��Apބ��W�N�'�g2E�4��Oj���ʥ.��6�.�/c���X4�τ(b%S�r��x)*ܚ��%j�d7�(�@�U�齳=��q2��'K|�:�ʑ����>
��x����֡
O�LD@�7�e��T���9�����x%���sF��;��%)�tw��g�5<L���
�;"&�GL�H���k��:[:p���Ziv�x3�:X:�/�
�>t6���k�d�<����f|����Om���L4����mtj�ᣵ����̏E�S���}��j<8�'��A���'�"6�ܡy��غ�Ԉ��TYR y�t�-���t��Q__{"���y���m�'��7o��j\��ോ���
�1�]�o�qk���H�)�������ז�=���u2��Uk]���;�ݜ�L�
[\u��3�z����y=�6����{	��tC��QՎG5��A�;���\y�>�и��W���Nz��FF�@Q�P�p�f�-�/Dх΁G�$Kf�kPVRua���I��{o,f�dkB�Gm+i�ns���,�U�ӹ["��+`ޛZͤ�-!6��d<:�cw�x���NT4��+��Din�`�h�4@�PZЈ�bլ�UT]V\��*$˝JI:r�H�H"e�r�4BŊaA1,9t�QUJ!����D�0��"���'N]�Zr9L��U���Y�ZTH%��$C�r��µ6Ȋ*.sB��,�P��G�Bq���ʪ9DU3�J2JJR����Dd��.u�DD\�5YӔ��Ċ:�Y��
"*�$�P\�r���U�ª�*젦�J�!ːDQ\"4����D��(�Y%G(�I(�Pr��(�U	*\�#3��2�uYrCeQ�"�D�(�D\KY8�r���B��UW#"�*�I�QA$���**� ��Y�Qr�Ȩ�LD¸WՖQ*�.��2�B,��J*�r( ���dDF�U#-+������Q�H"�RI��H�D��B��0��p�Ԩ�U��d���? (��|�32�f[�-��m�i���N�{�F)].r��ib�5lv�k��Vs؊]r�}˱����Vg)�
=������U�Y���<���� �W��X�D6r��]���ˑ��1�ǯ�li:� ��
��Y�~���1㊴?Mn�w����x�]z��/S>�k}:_�/t�!����[��9�p��������N^5^��xͯ2�B���/:vSڨm_��YdW�>�|�gqb�����1u���D�Ƈo����F(Qt}�\�o<dY�U��Kk�9�f�gWD=V��O*9Lm��70���j��*Ke�w��;S*�U��_�^�ĽWP�?�5�W�)�o|����W���.O%޸���̦����`�Њq�޸=ܯqp�.qﶷ(�>inz�ʷ��N���r¨����Qw����' ehy�ŉU-�^tCYuIT�'�ݛj��|]!I����ݹ�c�E��ت[J|l$������z��Vg��W9���������j��Ǵ�L������j� Dq$��s,Ƙ�h�xu�ON��0�ݗ��^_J�V~�WB��A^�w0��O^J[N)�����n��L�V9sp8b���6��gw����U*�򁂧c0�	�ő����@G�ي�uیr�Y�b�jG��:��@��}�W��=����iRX:����R�����Ŭ��_�{�3�%Sw���[�{{�Ωǃ�a�b�"�蕸�l=kn�x���:�@���o)�4z�{�:�GҐ�����V�藹 �Yu;$\`��>�Ѹ��v�~j���v���RN1�B��}�\�� �����S�{��dܽ�>Y��~ť��m���ַ}[�1<��MΙ:�go8�jw�%������>��>���i{<"��s��Զ��Θ�y��b��2[����2-�꿱���w��~��o�5W5����:�v�/O;���i^��	e���f��:�.�y�S�P
�0E�h�����C��w�T����j<����V�w����A��*�f�.��-`��-x%{��_�y�1_Z��bM��õ2���;L-���gq�X������J{�����9щ7y���c����DSՈ��o��71Y.aӍ�x:b�[w�_S<6�)���AK��f�� qgQɗ�*K�6I��:'��w���|3��=��o7)����+��f38�f����X���Z��)�#4z{w����T�coU֏w�Fm}�����i �����޽��Uڙ^�X�FL:������cF�c�h��pzq�D�Sp���~[G�3A[y[rrDC����u�^��>[L�8^ծ[�`��[���n'ޏ��-+��o�Ƀ��О�\��s���;j�};k�U�_	�5��{�T�0;�1��W�'�՚��[��d��P]0�	����R��1���ڷK�[ܬ¯{��4�^z|ֵQ-d��B��Co"��("Ɖ���Tϯ�y��Q0|���oz�I�����p�!��V�����n���3��6�+.��k�5�̎uf������꿭�ǝ�� ����I�;��٧�l��k[����j��B�_w���(��^�'W־���y[�gW�����y��A���i���M����Ȗ���mR�!�X�˞���z�ץ�cE�t���v���QV�\�����)��x{�r s2B)��{9�0D5e�Gsh���Y�ǽ�c�n؏��J�AӰ��@o͔�5�¢�e�����3B@o&��p!��ú�Tw��؍��u8�TUm�����4mAS�k� v��_}_}@'^O���viCo���Y���]vN��<����zſ��K�p���Rw�j�{Rw�>������y�O�y��^�a����W	3p�0�6�k�+���Μ���yУ�y��{�������yqW���SQ�l'����Ϗ��6}EC���7�.1c�N�hv�5��'g�5C�S�D��ᙶ��C�Ƚ��W��G�ZHzi���ݴ�ƋB״饹�n��Xv���]P����`%������~����j�[]WOl�,��=���I�~=���8���	JԾ��-��'�nεO�J��f�ǽ���ʒ^ ?����g��E�Zs�|�w��-�T;)	�0{ئ *�_��u�{=�¥�^eJy�I����`e�u�=�����ي���U��y�I���sv�Kܫ�-��7�3�M��t��G��C޺��$��:�^<�������Ėhs�f�
Co�����.���t���Z8^�6��w�Ǥ��F{-.�껛��O\�9�?U���i-���s�����Up1y]�P��Ѡ�Q������o��u02Kͫͱ��#3a��U��Gr��zN�tR�Ɍ��E�>N�ҏ���ג�r��;ډ�Vd�K}��ov����3�;eqz��/��:�_�*�EU�x!�������:T��,���=^*7Ann:nt����+=�)���^>4�����K�j��o���^4Sp�BN'+Y�ٸ^��q�C@/l�mg/>��J^�o| ���K��ϵuA�o�����W3c��"u�0{nE���r����c탕�~/������u{����xF稼�����U�%���|}�gN�m�y��]���g����k[x��1�^Ķ��voرmgW�ꎗP����N�r^�H���jYsz��^�18�1mx⫝z��P�^��/k�l������LC7�j�#��n��:�"�mBo
�jeW�ڨ�W���%� {ޭ�e�.�t/ԫ7UԖ��6f��u����e�����ٜ��b�[hU�����/Jˬu:��H�Iضr�����=�V��N\���ͬ�c��l�}V뷦� ?C�qQx��+ǎ����WV^������T�Q�ȪZn{��" {�1���Mex�=m0�����\�w9ੵ2�0b���Η�yb�a,��%�;F<���ж^U��6[ߧ<E��z�č��˃�ҟ~~��)Z5��y���mdYW�FK>�\��{x?^w��Z�Z��o4'���1�^A���N���*/3ecI�����[;��uQ�կ���x|A�1_"F�%S��#L� Z��E��K�w���h�Kb��J�ߧ���y���A�튀�4�����z=�}W��H����.�J�N���<�N!��W��;�=��ձCL���9_Jˏ(��*m7�%zkRQ�uX\?xǝ�� �b�)'��{>�X�z1���us�|�m��u9��܋��k7���^8B�cͳ�������UM�?N�߽���t�w���8���V�w��c��OR�^�	��%�j�Y�302l��R��+��3�\�$L�;���n��ߘ�����^¥)�2W��4�;]������!����u
���wү������T�4���P���ɴ,�s���.�S�@�(�Յ��tE�䒦�=��u�C1S@�LFQ����#�n(���#�}Ȣ}��ΟS"м��c��#ߥ�2��ja3��lX�Y��=�=��˳�_?祿��$}�}o�V[�^�K�ϥ=w����3���q�\W�Zv?g���^��}{����Œ�����ċ4�%��z�C���Z�(��(�����yd?x��p��3�x]Fu����T���*����i!K�=���z���}���n[��^���ͽ9�1z���������F"�^��K������rf�cԏ�y9�'?_ Ͼ��ά��}{k����;rn'ތ�	O(M;�;̂�Z[�U9��j�uI�!��N�9S/�eU��S����$���k}�N�)5��'f>��}���{U��T:�j!5�[b4��kW�R����z\�s����~ܩ��u�v�5��ؠ�L�s�fO����BӝiP��oh��j��pʶf�)�⯥6�&�#���L� ��b��:�E�$����9��z�����5�¾><ܪ�B��G��"�l�pc��������:JTWζᄊ�a�.�&iQW'����铻XB�p�F�Y����f���8�C�[�41���L^ɋ�E�n�t�4c�*h�
��|��w�*z�ſ[�cR-�+=U�<؝�c֕l�8۶6���4>4[���������K��8��.�Ju{n�g��+�<�a��/}�}�{����۷K�[��+O���u�2bk�y��O��O�vxC�����{�"��t��w��/��y�'�Y�c�7��b��e������c/7��o�D�Ɇײ�p�>t�HvG|^��@}�9}��@������v�9���!⯞��d��ճ�N.�cQ�T\-�8��1cV�
���jj�<��(��R���Or�]��
�e1K�����*5Tx=���E��BM2������K����X[���쯞np�L��EFN+���W5W�uv��ׅ�s���I�s#�����vR>O|i�z��>bor��4�="��5)�aq�w.�=`�:?�J����?a�s�K�*G����H�4�W��+aJJ�����屎��;��xV	�>�bؓ�X)�n�\k#��:֫r�Ϫ���/G���#��l<����?'s�
�lʦTd�D�z���B����=����e��<����^����ѯ�Z�����hx�Ӵ:�|��m�t�OT޳cv���c�*G�M�A��O/"y5��C�&C�_5�@����?z�WQ����Nl�䶘��*�j���:���w�!��A^8�H�z���~(Tʾ��6�'~���5䫄-˧��+<�)?Iwr�U�{VR��/[��ie���l=���N�W�ʶѓ8Yh{A
o��һ��=�)�R_��;c�^�����R�de�컋�i����b:���7�����<��T��I� �X�
��Nk�n5�Z7�h�	���&��*��J=�Fn�J����x��Le�6r����?H>f�w�~!��7zoD-�ű΢���򵴽쥏���{��~??g�^��ޗJq3�ʭ#Nyzǌ��W�O_N�%��gheDv���4l�o.���W�g�~�0Yx�>�X}��u�+
�6���R�@�
���N,ï��F�i�5��w֦k�R�o �=~��~܃�\A-:��}xb{#]�.Y�F�)�J���}U�)�sc���Bp^���<�Ëk���m.���P>��9x�^����zU��(�cb�KޑΈt:D�y�ϱ-���%Y�躣������1[�7h�+O�R�u@��=����er�x��=�z�X������1P������f��/^�I���Wۭ;��@Y�	�*ݩ�P���W��"���\K��VF{^R�}���y���B��yp�ya�\e��ڙt��R��=���_���[�	n�ݜ&^�t���m�Ӊ�Y�2'*�J��^����+����cv*|�'V��븒׶�����֬��������ܻ�Z;�Dm����+ ͦ*'VW�u�P^=����2�^����=Z�d�8����Xʂ��FZ߼#L�k�[ڋ���\
������q8��u͹[���v�@E�em��/D�m��#-��"1ሌ|�P�F֍��2�v���2.;�T�S���� h��r�	���v�`Q[yd���OE��|��Y��ks�J�'�Y� �B���
���Ur-۔�6�˱�<bI��E�ǻ�y�{��kCe������=�j���m�>Dȷ�.fEP�4t�����滑ܩ)O���w���Vk0�����Z=�8���e|�Ynַ�2�A�2!o���8
��tv���ٜefkU�gMX�l��FE
��1�݋��_;�a�t�V �Dc�zxCp��X-�}u�&];�5-w0\j�'��Ul�rB��E�ٌ�Ծ��n(z7�z+�8is͡o����_L��97M�&�����hN��`䔙��t�})��Zs����h�9��|`}t[z�,���Қ�����=ו}�y�w{�yr!_HBTp�[|D-(;H���W�ȵZ�]�:jr.���R����eST�w�^ћ�b�+(��R�����3P�L�t��o3��)ݒ�E�p���b��U�`�F�)��k�͏}���G� ��to�ժ�vTGZDp�F傦�MN�@H�9v���Z�gsC^.d�M��Fv[��N�1φ�L����t�{�"����{���װ��� H��]�]CҌ�fK�'t:-��!�k�*Ʒp�u�(�������E���cwL�'5�O�y%H��綯�npv���+BR*����s�2�aj~\�4w�V�ɼ�;%[6� C6�X���u���ڎ>=C�\�4��k-SY_��"����4G����M�bi4��;a͈olƚ7�p�R��17��'s]��e���DF�g����[4�����N +z��j��|pT��kN��M]r����OO������,V0�y��D���v�KS���mC� 8�,R���zc*�\��C���,�[�bх+��P1$L�	Mv9���_Pm�,s}�{���x�`�������K�Gb����7��<?0��~U��� V�[hw!%�ަMnЏ�fG�Q޹�� �ԛ��)	�Ɖ��-�N�t�2��!��^Y����F�;w2��GF}�ηاl�Ʋ�U��<�*v�B�1�u�兓�u�ԍ��n,��������^2�����{fnF�ILgt;>��֎�������.��^��:V�����q��L��(՘mx�0'%�[R�ãAлwp�w�=�a��� �X9�4�f��e�'�.�Mg�
GV_L�#�K���uδ	Ih��w���ުr.����َj���}��*=0LV���^��G#�H
|V���o2�i3J��6ރ;���Mm�[�rЁ>��9aR�kG�N��ktTot-��钸nz�����H3���k�]�	4���=�e[KƝ��L���c��=�ѮZ��V�Y�ü�Ģj�����V���r�u�nn��#UY�>��[��Q�n��P�b�*�T$�,U�Lⴳ̎]D�*���aB�((�Fd֨k"��9uC3�Q���(�E�*�I!DDQDEQ�s����*�S���Ȏ�-��*DBa]8�F�W9��!�L��.Q�s��<\��"�*�yiDQΠ�W��҈�+�Y,#���D2�*�9"��m5�"��I�ʨ�I�+���*Őr3���9T�eL�QT�U�V���+P#P�r*�QZr�5���ejE�I �"�PUb���Y	E�Y��2�w)���0�2�K��"��R2��T���UD���(����r��L��E�
5�qa��tz4h�U`�W�I���q٣������I}$��y���r^����`�e���iZpآ����eg��6s1�j�bem�~�;�:�p�~��ŝC�(��pe�rB��A��P�n���~���nb�C�N��^�i}� *����x�r	Ct%�������?x��*���ݟ���(߭S��ux�+��d=��>����olE��k[U��.�X�`�ߤ�?4��՗�ur�6qkO�@1=J�i����{���C0�>������(����σ�hl(�cتq��~m�>~3|��T���M��3���&���-����5R��#�l��ySؖ�L��v�R��7��G�ٱ�~�7���c�5��|て*{�s�}LQ�.�T7��t//z1�L��T��_ś��3z�>�U ��X��Kʢ�dwY�-C~�KUf�9W�﨟1W��(ʕ�jr<�97+��z����J{�x�[q�;��z��x�祀��Zu�g���Ҙ�%K�Us^���=�=�ՈػN��R���e���%�����*լ�mp,�m&1��ڸ�I���J}y��8;o���R�_�hEa�����{}n��tDP���*��6����v~Y�.�XN���%bb�M�4oB�����w0>�n��M�#�*�J$��C�^��D�Åe��b�r��Sމӄu��̦x�3���(�/���]�.�)U�V"��^S�.��|<�����^���џ4�OI��Pk�S*���U@�~T�����w(��3��;��'�^r�]��"V᭞�/�θ;u��uTX�pfy�G�L��A��]��M{5�+��&%���J��[;7v�c̟p��p{�pl�\E�UBZ��o"B�C+�gqeF�[�jtʞ�ޣ4|q���粄�y��F���=3���9�w�� ގ7L�W��n���{�noi����MV̽&p��va�fw������zE7]3���k��x֜���H�/j��Ky>�����&�7#��&�{�k0\Px:��������V�#�)t��cs(wE�k	��Fdg>����C�*����C��A[=�VN\Qx����k�=dr�j����)z��=��ފ�1��u?]N�����/�@�~�%l~[<FxlϪ6i�R�`�7Hf��~��l�{���ꁉu�}�k�����ҧ��W9�ZF�G��Xgf)��^�~_x��Zj�#uU�c}˔�����y>4���=���fvn�D̦�2ZN��v4@����m� �Z��/��kξ����o���]�۱�%��nn���2��u��^=�7�������b9����ӎ�ϳ��3V�}�����?�Ɛ���HW�WL�:�Q���B/�v#�����\��9���Z3���_gn+Π/1�����B♙�et̪�u3�o����]\���/k"o��K{ö�u�޹X����S 1:>b�;���.��L\a=*�L�2�:�L����b��\z�,�U�k Xvw��^���[C��z��ês55�g���1u]I�X(5�~΁����6z�m�[{��8�&s��X���w;��|:�����,\G��!�q�3Z6������픿T [�K�����<�Y���+n+�.s����#_݊���u��N�_��� ;��O�ź��P_~Щ]��y���Q��|,�q#���l\R�ٿ����Cu�gT����Ǆn
"~�򦡗���O
��Ł���`?���o�^ߪe��ݕ�z]oϸ����f�~w��D�J��oRT�t�U7�l�(l|9Q��������_�L:���+�][!��Q��1����=�����\���5���ꯨ��UPh�*;L=�}b�x?�:L;آ���L~�m� �b�r�0d3�p�4��+'8�v�NxAGz���]���@���Ϸ�ǯ8��H��9�h��@�Gx���H{�oJJ�y6m�w��w-�Y�݄W�r���S���Ô�o	���@i�jTsv>:;��/���s����NY�pWx���}S;�b�f��	�u��. ���z5;o��#�}Y4*0�^�>*j����r��v�ή��$�������葫�ϳ�<��9�ڠ���9�ň��$���IB-PS�\{��J��j\�Oe����M���w����~���G�a�y���O��:[��Nr�W맏4�~XO��~���r��eWs���ҳ��c|�s�+�X���G8�Y���oF�>�s;�@�+n(��A�
�̟v�M�"u���
�Y��׾>�6�{j+zk<��]�k�J���֑������wqYU����y��U}��v�;K��tz/��A//+�6'����:=>��5�u�6|���C����T�=O������]<!�������X�����O��7�>���Q֡p���c��t$;f�.�4c'��H�$r'ݳ\����$��jD���۸6���w;��|:��N�/��w�O���.�n�u���/yL��2}D���.�S��g:hnCT8m��H�}���(L�-=y�[#=sU���2NVqc6���{��\4�&��|��z�������};Fbm�<M�Y��K9��mŷ�9t5�q���|'63T�l�I�-�w$�s5kO�JH�T�<��3ۈ��{��k� h��P�g�����:u��zj�٣���j��8��O+���� )z6.�K�U�,vĨNpZ}ڗ��{.*4\��x�o,7�_Ez�d��Ϙ��͑:{P���J���8=�O��!ܨ��k]*r�o)�ў�k'��c��d�}Fsb�����UD9��t9�F2�Z�4O��7;�J��<����;7�{�kkVz\g5\��/@a����L�6���긋���-t����I�11w�pv%>�{"�'�Wy��B�H�K*����Ǚ=��ǣ>��3\�\E�UByy{w��Ȼ��:�cPk����^�8��]��fuzzn��fx��L��.+�)ʉף��VϷk�s��{�no;W�Ow�S��v�����s�_e]9���X.#��,�:|%W�t��>�I{+7��]�k'��wVy��Q�Q���
��0d������8�0"p8�<W�ո�L��5�9+�g_�n;�y>�s� ��$��-z���3���a�fł}��Ѫ�e�5к+��\}�{��uoUΪ�51-{�`��?Z߿޽��;�������E����ƭe�jRC]
�Bd5�6&Ҙ?^{�r�D��n�PAډ���z+w]��]�VwaR�@E�+,OU�K���=�75�9ėd|4�����H/޵&y��dqDg�f��3�/M����%N�]._S�<�UT,�sw��u�ܭ,=^�Ӕ}�fO����������.�=���Nsʤ���q�����z+���⮖�|ѳ�b���k�3<�kDͼꂩSL��sܲ!��"��e�/E�^B����{|��� ^���Ҽ���\fS�%J߳��<�96�Y]ny���@+�Tf1ܚN�nf���s�VQ�qŀN}�]�z�x.(��� ����-��[0puP�����^��u\H���j���A�[��N�!ߝL�f㨹�Ѯ�\N��D]�o�YA䉻O�����wtOC����d1>�=}�����0W��cOJ���T;]UaxPq� ޺��	���W�˓����.[���tE����l��q��z��T㪢��83<�¦W�����Ǎ��Ԋ-�g�>�t���+�P����ٰ�l1�d������bn{��k��S�⯭t�(��;�j����^�2�R&}ǴUc��K���f�uh����C2�.�9 "�3��;�L��V���:|}w�_Q�&�7��Å������aH�m������v}'Jt�U�$���~�U֓����;��w�{Cw�ߣ��84v�5�wg�,�Z���q�r�g6y�[�5��}�޲��q�5k��ܰ�v��W����Q�}�M��&ߩ��W]�E�_�
���e��ƴ���M�dIB����r%�6�|������js�}Q9��Hb�r336��Bk`֏1�A�<�����<�-ب�{�!���$^b�������/Ϫdm��u9q�`��U��dpbp��U��E�=ֽ!q��H�w�-�Z�B���@���oEk�U�W��~���������_����@[�ᵳ�'l��g��4_����JO"==ZP��meC���	u�F���������_���̯,�N�8�uq̷�+���+�*n+ư\V�����s'ζD�������s>��rJ��N���̋��v�r�����C����5�٧qG	C"��処en:�:��7�*h?O��99��I}��/����s}��e{�L �ã�/�;��P>@ˉLla=*�1��Qk �!����f�
�m�X=u��x����Sq���}e��T�kF����b꺓9w�9ez1��wp,��B�x<�����n:<7�w;����9N���ǚ�!�s5���#��f�V����5�=��/v�1�Q/4���*���ʷ�<Dv+���w�;��G��	����c�s����n�Ħ��2ӨI���۱A��z&����Wl�,�l���ȡ�ٕ��9���.͇��HcX2�j���1-�"����:�_Y�$틠�΂L��˧�:���ڎWI��ym�׻�Bj��-s����e���89o������ǹ�}j��=����(\ T<R���n<ny����pV�z��/�����������>����F����o7�D���
�SC��hx��GK��L����h���d�������R��{oպ����A�w��:�(�f��=��9Q����K��&a�7�f+��}�M^FG���]r}��*Gz8VL�w��\C���UPh���W��5Nr9c��[�>3,�赳:�?zzG*�*5��P����w��L�r��<���U����gpd���V5A��ˆ�O�Ը�o�^�g��ӵ��N��Zc��E�g�F�ˮ�9�3���H�~�<�o�}�6���aV�x�Uw��xzz>�s��K��ʫ�7{./��,�1\ou��y2���K��xգ/�w��9�`��	*�V����L䌼�=5����Y"Ү�>��S����9\O�zkK�j>i�?����5IW�k��?f�Ckض⮽U��>\e9�?{��n:��q~�=,ƞ�>
3=�7�ڪ���я��,�uzU�o������Y���N⮲��O!q�Ĭ���=����닫�hX�9��;��3$e��U	��[ϧ����t���~��d������T��.@ds�{C'��m�#����-��Il=o���oA�>~U[!�oK�]��sː�t���b�mnppl|�C�r����J�'ͭ������gxM��)�}�t��S��u�6]��7��d��
�9﨟#�)r�� �ޭ�f�������]�b<��2���z��,��P�|{E1�Ȑ�5�w\�3ʀ���4}ӻOݍ=�.z��f��-���u��y�pm�q�Σ��:�������ʶ�k��U�g{U_w��L�cӔO` )]�W)��F泝47��o�u)5��Ԧ�?W�̽�V���5toK�:/�q�����Q������tJ���g��*ɝg�{`�,��\����ª}^Y^��N��]Fp�S������ �)m.��]���O���3�%�G�PU��z��ku����sv�E�u�ۊ��Hs��3��fUD�Pj	��ΰǖ��xί��I���y����90�2�B�(d� �+&j;���U�\T%�p�������6�{���ݔ��ɞ��S�~�\+4�u*������C'�s�TdW��C�g�� ��n���[O�-){u��L�9=v�6qW`�x�ʌ����$�E��[���Z�ȹ��9/��ؖ���i���
����S�~3§{}�<7¦��Ľ�{s��������$�ťr���H�FQxb�~y���&_A�܁ӿr�,��<����q�¡��{��QH���F�х�F'�o�nQ.���r��ön������eHv�*��Xg��Ų�����o�����Y#�Ȕ�S��k0\Px;}��&�*���>���X+j��*���}��������,�ь���N\]�ʰ��\��}�v�YY���<=/���s}s���[�c�b��y�������u]%{:�;wz�}��XA��ꠅ3��W�z���xOs�/M{Qw�Y=�z�y,���+�8wӚ�z�*㶽�g�>ͺѹ����
��R��q��{*��1jȋ�������{p+z����>
��������yT���5}�0]o�d%r��zϚZ�7��H>'��X�7�0���q2~�޸7J�g�Y��X���gtx��Qӧ��)��������� �ƣ�_���Q>B�)����R�:�|�r_�!�5;�J����G0��[�`/��;�x_q`���G��@�Q=)�Y*]�*��aE���O���]w���w�_Fuq��ʺtuӞQ:p�q�S2����j#F���E��rTY=�*a?\_�/H�k7�s���kx�F4F��fp��<}'���Pw꩕LN}�,��==�@V�"��8g���]xT��ҧ"��Fr"VKdٓzֲ��/�,��14 ��캾�����G�/�r�D@vy!f��Q���dg�S�VB��š���ٝ�AP���_m �2���0�;�J⻇d}Y������;ڻz�;O�X���{�yH:��_lrҳ��g)���l��_���݇S��|�̠��'WY9G�̔gg+���-��a�G"�L�*��ksm�]�!�����.��A�{8;o~��:�<\��?wm��hf9f�rP�90�K+�Ag_ Ñu�r��0���pR��0fB'[���v�dM�}]O�v��S]��O�̞�i}(ܙvٺ_�d�U�3}�VvvkĘp�Z�{ةf[��sz[���fޚS��+�k^�'��f��������u#�C�d$Iї#��f���$<-���س��(�^�w:p����	9�z1Q#9�f�ܙ����Lڷ��/�&+<d\����4�k����W���w�ouY�����#�i���,ڽp!�^.ԪR�ƯY�v�]ЇZ�,��-�C�RON|@o,q�$?*ڶ̽Z-u*7��	�[֩��>���z����׍��fuC���1p���H�/�N;��hs����&lH�;W> |[9-�pg^����3��ݚ��#^�M�v�BG�c�Ԑ��1�O�fy�b���u�5�^FR��R�]R��Yx ����+پ��ě����X��}y��.�֑5�ј��Q�ۙ���{�Z�Ѵt�9g�ݳ�����*�8t��Y	3*���������x���Ϩ�z��i�-�흜���h;W�G�폦wg#W�ΥG��q�Ɗ�.c >�Ժ��ky���64 �3.���s�Y�8���� ��[iYB9R%Eڮ�,l۫��YAs�܎\���h+IE�g�`��!�uC�2u\ET����]!s��$��M�;s:b��zu���p��K�w%oEәzw�G�(3}nw*�˺�Z<}:f�Խ��r�Zi5�����������P��1�(�ś�u�ݾ��9uҫfu\�+���R����zxg�4P���U��h�B[R�{��t'�^�O�K�<[�E�3�oD�,�G�9@x���Ӑ˚��{v�φ�T`Ws��E��Z�E��꽔�w��D'gx2e���B���k��j����)1�n�S��f�Q\۰��%Z=\�͵����s��Q^"�۩�\�y���_D!����:�ˈ�#5��Yw�eZ�D��F�-"�Έ��2��N.�}����v;	'Dn�>b��]vۥ2��|j��x\u���Z`�x�v0��O��^��f��.�ŕ�)���FƬ�aHB(�[P�@P�/\Zn�uۜ>���&�Вw]�[�sU:<B���t����a:��M�rBs�����}�����H��U(�ZȎU\��˲*.YйA�黴"��*
����9r9I"
����vQr
���EȈ����2����V��^$�˕EG"�.EÔS(���W��r��E*WdUȥm\8Z�\L �ȹPE�9\�8*Qs�Er"Up�e�(�B�EDE]��Nr��*��C�vTr�ZĪ�(�e�"d2*<�sĔ\����"�Ah���ATQp��(����eEp��Qr*�P�EvUUp��QsS�*N��Q*?u�����߉�����e��%�r�`�V.�����cN��������,t��]�^�}�v�1�r������b4��y����o�*�s���l��[�����;�{�%���`Π�}]w��ê���83<�r��nH��n[���pw�\O���&�$s�D�q��Av�c��p��:���	�0zøG�kG���������4�>]¦T�j�������1٤K�{��������9֫*d������VK�������3����=vȸTh������������eه�ާ7Mw���t�U����}�޹ю�Ύ�p59r���f��,܎GĚ����Px:�K���eT��q�qj}S���~��}ʫǷ�e���dgu��C�> �}��8?A[=�U���G_Y�:|-�7s�JV��C���Y!�Eトw��J�?]N�~�^��������iRH�����M�?��������Eq�2�0���sh��	u�F��z�*n;}��sכ�	ǭFr�x�VgY��@�p��M׍`���HX\�y�ȝ�u~�йy����VݿUew��n��}����x�}j3�Ɲ�\VU!qL����U�d���s �ˆW�ނ�\i2�e���,���x0��FQ�{zD�b�[09�T��p�s��k�O��6D��{���Qҧϔ�y�<��'6�랎� n�ƣ]�Mp�y���/h �z�1�VV.�CaX�#�-N�/����K�`ܾ4d��_PW����z��y5��S�� ���V��f��{w�����r�n>V�㷶̯w��d[Ɲ�z��AĦ.0����J��������ʂ���֗��C�J�_T�<=��㓭��ːd��5�g��#��Cɹ�D�Vf��1ر_y������x���}��;}����,o��!��i��j���̏8��k��z��GH�a�|v��w�+����v�g���;���ў'�#�Κ4��ҟ{Ջ#��:���Yq�&�ɘ��3��������."��͇ճ��n�@�ꃂ�cٙ���|_�+m`���[�{Y��}���K,ڀ�k�T���*���3��nu�t���»E�E�uY�����=����Uo��9�P߇*3P|^���l{$�ɸW�{
�����k�D���w�t�����b�f�;�}"�uW�bʪGr���Ph��rŨ�%�{����Z�mf6GwI�O*���J�(Z}S;�b�f��	��^�"ૡ�{� ��.�&��o�N�</�������&�
�QWP�z����\Wm��p��r�9P�3\�D����Ⱦ�R���T}�[�8)����Tf�T�.J�6H��_�2�m4:S͜敨���� �a4�sg���{���	KuoP#N�&��)�R��έ=��wS��>]�oTe�MB.ˏ�t�L`��Ԡ��9g H�5`M��o�������"����Z���;�� +� �'�p�>�5.^�ˋ��K&��7�ﻮ+E倘�	}*s���H�w�|�A��U�[�;Օ�/�g$f=;[Nnu�/䫷���ɉvF��^��W�?3��Gӷ���{��4����V�Q�8�VS�����i=�0}���$e�~W\lO�����`����������2s����N⮲��q<�1"W����z^娮Ƴ�$�=���xNAT�1�.�7#�ܻ�;�h)��$�r�S���Y��#;�)��Y[��X�p�E3)���_��'̾q����z��)gP���c��BC�gr�dQ����W��\��2H��>�<���)gTT�y�pm�q㾎�q��ՈGE���{�c}f�ڋ�oum���K .��h:�O�����T��R�ߩ��Z���K�l�V`��*4;o����1�[P�w(��3���Zy\����]�����w�'�����Q�7���f^�9�Ǻ7�N1�ɟ�r_Ϫ�13)��2��S���
^�}�����?*jovu*v6F�*򤎯9$���Ŗ;���jӸ�K�Q�iMq���[��!oz�R鍺�:u�08��\�n�1��(^�=���Q�D3�te�in�]��v��"�鬭���RR|ۻ�ᓰ�t���9�#��ꪥ����t���ڷ��X
!�����g6����UD9�Ds+	�Pт=�}�U9���~0b_���L*��z/�Ohz9�?p�������u\E�UBZ^�[�%\V�mz��85�+��I�9��/�=¢3H�P����}A����&=�X���x4l8�;o0���u-Ʒ7����ndɕ���W`�G�������ڣ5�S�[3��&p�/V�W�s�m8��r�jz��?P�S ��o�k0]���Nrk*�����nd�UƉ~qy�x��ت�>|jv��\]�r�$� ��wn;�YY����
'�����LzVFR�ܵƞ�{�y�.�����Q����M���83�T�v�j��X;}~�*/�:����)��������i����7�]Y���UӫMN?��p�6�F�DOy��5�L,ww��V��歞�O#`����X�	������ϻ�Ҧ�9����~S7dWF�Z��W���t3Y9q��
��4�bX^{|�&_�����SL����r� t��7<��E�3��X��*�-��:��wLt�-�o��y7�X9iS�Ё�E�%d�䶱j���pR�]�/}J.����+*�fm�4��L��Ί�e�Yؠ�ܷ.}��YۓF��s�qwV*�i�X�R�t����
��~�+�1��c�������TO��fe;�2�^u\����ɥ/���w�pj�Rʳ�����*�R����ܢ���X���8��:�0�~OJb�R�nG����{��{� ������3�Bg8b����WN�e��}:p��fe3�)���w�p���n�
�eB�5��Nڵ��/
��5=�{�����vg.+��wC�W�C��U�QW�/�N�Y�tyo��TV�OD��0n"G=>���J�DK�����:���rU$Th����z��Cٚ�m�L�r3��#�윐�^�%�gV�̮�(d������bs�!��lL؂s���-IR��"�dq�-y��SC����UŜc�3hK��&sWV��lV����@4�Go�]��^�F����������ٗ���|=k�gz��-�����V�s�T����w�t���tw�59r����^�o����@w��6"���O�����w�^�כ佋�htC��w��\{z�Y��26���.9P�wʰ�5�C��g��{���U����٭*���J<׻�>����������w-�E+��Y3��:�W[�w�R8��R�l��cw�;c ,g��l
��q9��q�vu�z�0M
�7_�A�܉�3��g��q�-���}}��g��P��vzvۊ�Z��&Xk���쟪WQL;�ƌ<�����Z�2zN��~���߫�=+��"�$�vrSp�o����d��M�?XZο~��lK�����T9�E��������p՛��S;~F)�>���Ed{vr9�{<�+H���P=\)!Sq^5����S�1�["k{]��O8�y��鄸���4��<KT��ϥ^s�R��=���q�qW�eR��,=3+cL�v�ޛ�KN�gb�������\�j{�9�)v�ٕ��S 0ȶ8Q�"�q:�e_J�����-��4κYY]�OͰ�=�K��ʟ;)J��h?w���Ω��h�q��<J��U�T�����<u��t��u�z,�jm�������w��Ռw�t�.<�	w�����q�1#�5^?n�{�g��d���93�b�;�W5��hƈ�������w�8!�6)���/zgws^׷�A���T�H�5�p7!1�<��Kkf_�ku� OG�w�I�^*�Xm�`�eA�\h�q�f'��Tʚ���j��o����g����}�k�{�2�V�[7'5��j��"���Y4�|��.���p�P`�z�2,�ă*� �]�yc0�u�f��l�D�e�&��/B�w-	��b��%�9Mm���"��w��o����b�1t��ٝ���"!^t�0֕��y��|�2�8}�d���h;8��ճ6{��6ꨳ|́�{	�'�2,='��1��R^���u^�	�Y��Έ�\E}�l��b�=#��L�w��[���UPh�*;L�S1�J.����듩q�%�G�lmgI�K*���Op->���1Y3Qʇ��:��
�ะ�}�����[��U�v�����VM\ax0ч�I�}z⸋��H��g�ʆ	��"w|rD!�cK��ksx��j�	������`ɺ�7�zr�#*�\ޞˋ��K&������Ξ��+u{k�m8���~�|�(]��%t���++4\S9#.#)�MDem9�E�H|x�f�Dɬ��׾��q~�"x��dN�/�3�n��������@�AmEa�A��ͥ�wx��j�-S����C���S̕�n
���﻽]�.7:�}xF�!��6w�uV`��Ӹ������S��i�ܜ�����%wѝS:�𜂩�c��t��u�w�X��G{(0��s�
|�^�/P�ʿT>�~~l��\��c���rK~�Q'Ο7�>��Nyg�֠�v
cyw�`������x�~�s|��^j�Khm�J�}\k%�w+C�{5,�3�,o�E�ӷѱ��	�B	��H��0R���ue�j�!�ow}-��!�dk�A�ZսpM�s��nl��WD.���[O��A؝3M�����鄗d��u�V�I����=�קo��2}GԦ��-3�R��닚��n���+��w;��)����Ƿ7(���K��Ε�t_�ŀ9��sA�2}��]�u���H��s���u/V��ʨ�����U1���R0_����ܢ����O���i�s60�D�z=g���Y�8�s�̛�����Wp��Bs�����\W]�6����̦o�e
j&�|_���敾�S�Ľ�y{;Ӵ+����p`����fv⺯��UD9�wC��2�����}^���sN.h�������`܆Ѹ�I��������C'8��5��o�긊�x��ium��l�gq��7���b�U�*L��X/�x��K�YTDVk�0:'ܘ���F����wb��n.*�^��pBg��\@�D����(��b,���C�y����v��ߐ�E��n{�k�U�=�sx�۽��e.�qX.;�*'��#���'��5;=胵�.��ۥϧƋ�9~\cs�+#z�G��������wT�7us�O������r��#�a&�����v���.��0fM.�tf���շ+���5��;��kY�<��虛0b[	�Tͣ�J!j{�!_]����/[8z���^X�����[)5n{׶p�wD}��k�%~ٵ�����6��s��{�$�WPj:��v��%f�y�0��}&cI^���Q�6�{�nR���+��=�.39��OI�οN�wz�}�����$hL�l���*��.&�=�w5'x�tP��� u��+�8{���V��ו�6}�n�o�[3�:a`�3�}gW=W��g�6�9M[8%S��r���/����ޭb&�
v�G�ٱ�~�#b�����W��|�oy{�]X��'��Y9q��'@�,o��׎�d��\��4�٧Y��'������ix:����D&�U��ŀ�Q�.#�u����Ļ�J��gU�� ��hA����q���c�c�Eu��=����w(�Gq`����]�z�x.��L&�'�1QB=DQY�BK)���j��_zY��j���ǲ����8C�:����vq�
r��q驇u�>�c��̽�^�4������J�k4�F4F��vg.���.O����R�$���Yu�>�o�5INe��&�����;���u�+���=�g�Ψ9��|��e���O�<���ض�Yc��3�~2�Gh3QζM�#�W�.�:�vn�ǡ�� �����&Rt�g:����A��]��;�+~�6�Ȳ�VP�bn��|�/.Y�sM-���e5y�;��͇""*?��Mtw���W2�>�:勫6���k ��v�' Z)�xbwE78��ʶ�����\�	Ç�҄�\;�s�ԇ0�io�N�5��cKzvp�z{��i�pUP�]&eN�9Q���V}g��6����:���n:���U�)�6=��u;䍙�sQ��������F��=�l��f��/ިx؛�)J�����`-����{��)yWH�n�gGz59|�.&��^�n7#� ޜ>�����S�4���C��`�ʺ�j��{]L�|fFou���*.�9Vg���瀉��rl��Du]<Ģ��%ued����LTe]C��{\{z+X�c��+���S��W�zf�PSF~
�l�㻹�5�7�n�\6�_���� �F2cݷm��K�x{��\5L�2�1|�IUx�����{ߌ����d��c�ws�ѷ������|����/L�9"v7��M�;�tVT��fK�T��Uq�=��^����\g=�!�~8�Dq��i�Q�PȊfg��WL�ػ���~����^�7������:�0z"��������<�;�ަ a�ldq�q��( �L<���W��-����T��:�L{�`�u��E�Nm���:���r v���0F�EC��׆N\�-X�٦�з�n�}�Q�u�ump�ڊ����Q�p��O"�\�WЯ�mn9Z�o��
':����۵S+7A��F����:�lkg.-0��v���Q��=+#Y���g���>ݒ���".��
FЦ˼��+Bi�M��)v%�Z�ld�2qݥ�󖁌D��;'�{�SIR���2RZ/�D���껏���Iƃ&�͓�d�Zhm�]��OY�_c9[�x$�o�vq��U�ʅ�1�o-����]�P�v%v���r�����C0 %�	;w�1^�ccP�{����.�b��e�����%҃宎�~~�Q�� O���O�e�ܴ"���M�tУ�Ԓ���l����=��[���<��=��e�Vr��Z��-��^���lo�c��\��+�������ll<;���8�?��'�&�'i���O����ڕ�PQfg�׾~��&�@U�8��.��z��NQ"��m�d��������7Q�����[��,Q�Fp�� ش��w�S���tX��tƦ���+l� ��]`8h���ճWYH�yЭ�ܱ�]V��,��a��x��;]}�ж����I�{W�76�mgU�<o���WVd��o�&�b";�g�`
�����ى)��K�{);t�8��ά#-���WWR÷���6w�����ֵE��7��`]�4��)A�b�:��t��=t#�_���7�ҏ�^��k��b��X�P], �w�}���Omr���=Į�I[�h�XBnvtz�5_R{�z�����yu���L��w֕ih:�n����q�[�7L��mu��m�����i�c�}�_8�^wQ��V�9���7������+�ab����q3w0/v:��c{o�� �[�͍(����'!N�R9�N��n�d;ƈ�HV�.��y6�q���5Ӡ/
�7Gu]�fV@1rվ���z�r�:(�y�6�E�Ut�i�ف�}�ò��,��\|L��v���ӛ��ut|nt�.��LO:��jV��x��z�4���n�3�Z�V�[�=JP<Qd\�j_µ�Mr���;j#�q�Q��eo+1��6F��vF��А)�	�ٷ}��Ѝ��j���s0+�^a�M�}[��K�����S��4c�`"{�:��v9�-��]�1bj ;A[�����e�����9cN�	^Ö��V�nWy�x�A�C�xv�)�H�;���(]+�E
)a[�vo��[��c6w8�����fp�$���8���������
u��s�F0f�.�=Oa7�)v8�EYPKrܼ�n��_;��K�Nܓ�/_�\s��5HXA���|-\�c��٤$)-Â�C��ں8)$s]�	�Òs�[�]Ӹ^�,���NU�f4�S�6d۾�2h_D)��EuK�y�[h�gi3�c�U�\�gNq�)�u/A�.����'����{۠P��r~�(�9���Uˑr��Pr"���T�\�E
��reT�
��PD��
��.uI�G�
��\!�YQDW
*���TE��Dʈ���TPp��(���2Γ"�W.E2�#�%ȣ�TTȎr��QȊ�����QS; ��*(�I%s���E�QTTTP�U�DUEr�Tp�"�X�8EDD\���r��B�Ar�ʫ�"�2F���J��N\�.E(���s�*<q��
��T�ʈ�����f��9�TE��TQ�"s�r�T�Uv\�$t�x����N�w+�(�rl#�M�ZGl3]c)��q������{D��+�+�o���</�WՍ�$�S������&nAW��j�J6R�����=��ݯ���[��Q��o�Q`���깯2�3p��ᾎ�q��Ռu@�</�G�x���2��S�~$~6���\��1tJ\jjS�W5�w;Z1�0wb�>�뎽Kj�EU�f�5/4�l/���t���Jf�=5<W�$���x���߶[�r�����3�1C����F��:.���|	��EޖXk Y��C��u�3��I6���Y����=���Q9�{�Wpy����ճ7�ނ�%��lc �'��_���.f0 ܺ���,ιt��+��N�CrnzG&+&k��_H�uW�bઠ��*P���"��C�,���SX����=��V)0�eQ�_B�O�g{�VL�"���zx�T�}����=a��W�7��ܣ� _��f�5s#���sW�������QW�+���D����S�7ꇼ�1T���su%^���/z��D���~�V��g8o�ONVU\����t��fw��	�����n��'�q@�*���;�����lv���p��謬�t�H��s�Y[N}�y������q�)L��֡��c+���V5�=�U�mZ܍m��WKȩ����kku~T�����HP=羊�n�u$W�:�pBGYԒ��җ�%NS۾����h4s�^�f���������+m"xP���lF�eۣ���I��{�1/yY����q,��9���G��a9�j�C+n*��U`���S��������ZV���|�+���'`�����v���һn�F�u�l����;����b:g="M�����lu�d�J�3+��;�l�r��O�����״�#��Y��'+}�,�1\}��Voބ*�s�D��<%����+�Q'�:|�7��{��NydZ����t&M;6�{����
��~T$;�^�q��>��SuG�>�,J�.kͻ����k���ٚ�y���V[�8�ë4Gz"w(𿻋 u�4�vF��Ȣ^�%J�]\�.)�w��Й���'}�K2ۓ}H{�z���R�����;�X��3�'4���3�%K�#tv
��wBfo�uj�{9��ٞG�{a��;3��NK��G����L�ޣ(P{Q&3^�\��J�]��"�ϩj�^��K��G�仧[��x9}�d���3�]W��Is�wC��D�ͯ�'��v��ps�\z�/�`�H�ǲL:��������}3��k_��s/-y�����er���j��)��f
&�v�=��֑��?���X�X�Tk�"yP�
�)d�Kή�WdN��%\݀��I����ѻ�Gj�/Y^�;�V�r��뙲��oJ��z����������=�LP�ZGP�����(��oL��7?LI��p��q,�3_t�_����%�ʢ#5�'�s��k�Y>�L^_��Vc����vP�}�dYUBZ��f|}���/�fկy���'khc{,~߿6kGcޏ
̌m=*�}�����|bTs��9��@5;=�;Y���ٿm9�ݾ6!gȞ�=SI,�j�Tܽã��,��:}�jv��9qwʰ�\Ϥo���z���Q2�gM�r�xj��C��}����=����Ϊ�+���������ΰ��=�A>�Ȯ��1L�󥙏x��k��T����q'ݵ�$c4w��z;��uoUή���Lu�w^�8]��;^WV�P�W�)��>��t��7�2~�ہ�u��������������6�<v��~���y�˞�ۦ=�5�5����7��,K��j�����z઩�����>���r-<�UƼx�mg�oP���e���X�C5b�u���'�&S��2�)�GMC	e����{����<g�<��k+������SѾ%����٨q5u�e����G�b�hzl�)�M�)�Fd�U6��4�s2�r�Gx#,-�� K�nPq5�e�7sX��>���eYt��-{�	E��㹃�p�5A���z��{��(�An�{��v�oF��fl��G�W�f�]��d�w��7�Yn�;g������N�u�d��=��DՑG±F{B��ޟ!�Y*v���[��#�v�ӌ�[��!��u3)����r<��j�'g��^������c�B�}vT���\�Fi|�����v;3�]V�����x�'uT�\�ڮt�\tЮ�UL�N�D������㵘#�������g\�'`H���c<�7�wȟn�%I�z6������<*eT���:�7#�W�.��gf�����{.��x���Ԏ��Vy0;\lH�ꃐY�"ʪ�I�S�����Uc�6��������;���
�O5Y�3��\�3�sQ���@�.F�� 'f^:p�o��%��de��A#��E���mnt2:;�Nm�*7ʺE_��L��0js���y��Yf�r>$��{�X�n/�7�}P��>	{�w�-���F��*���X.=��x����F}�r���a_��{w�>�y�����s��qNx���E�`���a�Ѡ��oEk�U�W��g�˿~��z���Gܐ���_vԀ�!����Q�7\p���O�n��P1.��Beotqr*��N�CY᫡v�{e�i�vF�=K�nk�+6��wYz��E���kmI�)%r��t���� bFᡏ-֫�,o����h�zL�k�~䇫øol�����ک�u*�7�l��{��
�z�q�h�4Ӷ���H������̛H��I���N�<U���*�wei����b�7^5���
��s*����}'���{B��Z�����'�Wgs>��qq���群<�p�{�#�;����B♙�1�\:��njnu\��{q�왓�=����Ҧ����o�չ���+��`�q�q�浇j)���A�f�����eD� �{L�2�-�����O���jy3���9 ?E�'z:����{ך֣{�g�+���`�)������̶�d����;}���9�TҬFy�y��ھRhtB�BB�4�kFӑ��	qv.S��qsY��hƈ�}�L�;��V-O��Wbº�WhGF��7�83)�3���+��LnǍ�1R�ٓ�^��}f����e���+ �θ:/��w�����3��fT�{S5��zOK�q|�>θ���3������:g4t?u9���x>���7��fl���l����61��e
�ʌ��\������&�E5�1^��=:q��&fS"�ul��+��;�VL�wz�@f�����M)������g#JW?�q��ʽ1h�Xv�渁��lt�*��n Q7Qt����|�7ujO�2e�7�V�p��o���uU��;)��q���OR�<z�w��
��9����|3��Pks�' |���n��ùt�]�Ġ�l��{*D��X���:L:�eQ�i|���/����T<'��:K����J��q��S�qWC� P���65���9�/ax�J�ͣNo���葨D�^��q����b��K�0L�>�*9���;��&��:}�Ur���\.p3 'yb�jz����f�d����F�:����~�������	*�n���6"��q��kwg��=l��])\��imU�O#Ւ-�����5<Q�q���w���}γI��5¡��u������g��GE��g���ٙ>�7�bB.}�~��v��.�J���/{f	q}�u�5������߇
�dO��W������8�B���+���F�:���ss�ܻ����	����۷�~j�X�|�r�Ut碉�1t̴n0Wx�$���f�����sȯi����-��ΙW��o+������I������J~8/�����W
�?J�^m���0�V�l���e�o=���>+����X�to�cc��\3Nf�4c'�D�J��jS��9Y\ѱ>�Y��$M��e͏S��![m.oq[�f�'�J��7�.���+�	!�G��F��*�T��=q!�	)��"v�.q'�&�2�Ļ��Ǥ�WDZ��no�2B���n���a�p�B�V�3kF���N�4d��oV�3ОW1��{�H��]Q�'r�fbS��P�tr�������e�0�2�χ��5r�/f�ʱ�v\��]Y5�ޮљМ�q����'!�Q�~ffS7�2�����mB"�ڮ^�����Ή���t��9=qպ,���=Y"���3��p9��$
��٬�����R�������Pj	�i�q#���&a����2s�~��7�)���e{j����T3��K��=��Wg����s�I��㥂�/�h�eQ_f��e�	 �GW��ʓ���g�K��Q�Q�C�g��# ��<� �����7v���������ͳ����ˇ�⽋Ƹ�}�ꞣm����1qX/��D�s��*9���� jv{���e��1v=}s�.g���/bǳS�����|3�oT�oήx��w����\]�*�Ms>�Q�;������Ӌܔ#�HtPL�xa��=�����ꮒ���7��]�ߵ��6�!že~x��d��}Nj�U��o��tO�L<��L���7���Vo_�W��'�|aߕzf�oĊ �&�K�p]��zV��M���X�����e|L4�{����
�7�6Tv!pMw��{ӂ�]����n�( ���و�Wgh�>1���Y�z�`�Nv
6v?^7|C�-�x��24I�f�ޣׯUw�NX,�)��F[QfȎQT����~\==�<ۭ��B}L*SDx���fy��Ly�����X����5�Nw��^d�d��%��N��~�7���D?�}Ʋr�b���̰�0���q3I�aZ��V~yޔ��e�vA�uϏ�7=�!��"�v]!\˸f��_�k�$�hg�Ļ���
�wY�ƍ�wKf���s�]�W>�zN��c�Eu��=������,\w v�C��:�2�|$xh���"�ڞ��^IW���O�u���\�{�c<����v���ާ<�N���L�N��TÂ��Y��Ս�o)����xeøz�w��K�d4F�tg��u[��"_v�gس{kܤ�Ѱ'��fw�Kꉯ�yq�r���*�/������;�M�z�*9���A��ʩo����� gI&y(3<�$���B�f�(��Cs��	X����Y�x�Uهx�f��Xc��0;��"G_T��P�*�K^��S*k�ʌ��z*�,��ȍ1q�?)=Z��NK�L�>u�?D0zg;���L�_\�����F�� 'g =�"2J�<a�]��~���6r���bK�:Q�t��i�;Ċ`��p�k:ӫ�r�'=o&,�B��ݔ�}�\�ƤU���\{����-)�4N�8�gY�1�jL�+����&�wO�.�a�j�8�}�:����ZFjg���M;7/��+ޡ��<.Ic)q���K��C���ߟ徾�0=�WH�����N_)ˉ�u�$1R9��S�Ï�l����Uvή�ef��,B��YWP��ު�q�S<E��L��>�G�%�RDtk4�0���[��3��C�	Ӳ�*�ˊ/ �`|0ч��E�z+X���J�y=��Wӝ���[�/��'��r����� /ӧg���N�q�2���L{���� )C�x��[��J#"��ո��������e}��O���;��:6�_qbS������c��z{�sBn�f;��ɮ��������}=��ˏ�^s�R~8�G��qƝ�_ՕH=�'u8����4SQ�:����9][3.�:�Lk;��ZAus�7>�����e{��0��7�w˗��]\��:{������"�:(8���x�d��������O���jn9:���#��Ghj.�����R �*������g�T�1�gU�G�l����s����&u�#��y���t�/f�����Y�:.=ʄ���4�j4m9#�%.>�r�Ҹ�������L8�D���4�w�q�%l'����[O"�t�lc��9��=ɣ8�k{�ŝg�M�4a ��@������<:KN�꧷I���>�󾽘�'�C�;	Zg:���VPe9|EW���hdp}�|p͹�M�T]Gv�"�ND<�x�Qի����ᝉ\����ܣ���2�Ǎ)���L��\�Lo�O1y��t{ގ�gև��UڼNs���=��냢�����<.<����4�����`*�ࣺ���R�y{�yfw�k�u2ب��ٴz���>~��ّ�� ����61��e�l���KQ��8^M"�������\.=�c�3+���ul����_1Y3_}���]_6��c�ٕ�}:g��Ӌ�^����&�_ҕA�'9c���Vt�t������
�T����ɗ�'�t��yt��r�4޴�p�;f��x�S�<wO��ՓW�ଫ�{đz⸉�t��j��ܳ��u6��������q9��H�������@+M�L���팪�sX��y�Tߨ����,�٫qm�d�y��w�ƶ��&U�������yƿ�W��k��9#=ݬv+�{���SŅod��*��z�E�%]�}��⏣8�v������i;����P�ۊ�����z�C���4�����5 �2�fO��M���&�*��Gw��,]^�}��#}֑���C	���iث�,��Isw�~Z$�;�^�b	U�2c����1���[�JL�����A�Lș=G�e"���3a�w�$]M�V�5�6q�{��oPT2��}� �ՉF�N����\�����;��;��l�IOs���֔�p���WQs����}J�}��S���f)e�+B`�v1��G�2�{��,U=*�j�e;�;r���%��G�I�=��#VE���mt��5$��� �
ۛ�sp�ya��3B7(�1N˳��zU|�	������Pk��Z�כ��[y|���0�PN�]<fpԣ��_D3�_\u�����*֍�[�ޕX�T��r:Bf�Ww�2���5)�V��V��kp5K۶R��Wkۛ�U�{IY��m�q��dF�mP\nmO6__�c��E��ή���i�:�\\fR��"1����D���r�=���Ē����O>3N���������a7��rB�:'R�f.��:��[�)��}�X�|24|�����Q��,շ�yݗx3����<ZdT�f���^C��޹�J)�oH�`�Z�D��g*�T�;E�û-�I
�H��3*�;��EGK��:�{�'�:l�ng��gS�z���n�e�7Bb�A$�|ha��u�fZ��+�H$R|���/�
��Av�*C}Ep]Y]K[���{h����V �e
ɋ�%qg �\$��0-�DṪWjM�������ﺂ��^K(�ei��� �iL�VzF^s|�N-���Dƪ���:�N�|��xt�=�w��m������7z����:�^)`\5�N{P�W����nK_�ǹm�*�5S��l�v������~Ҵ����N��f��'J6�ʍ���+����[!Z���,3�cdv��:M�)^�=�w\.l/o4e���Y������z��n������x�ꍊ��\+�wb��7bӀr�����u��G�eh��2Hff�VjJ�f�p#{K"���j�٢jX��jr�cAQR__@�S�N��+M\�ؒ���:���=g�.��n�݃K�ڷ���Z58�F�f�!�Zxt�B��9]
w֖),��v�W8^ΠQ��Vm�|�ێ�t,js�z��k���!Jۚ�o)sWr���g��X�N��{�u6��ቁ��6ڗ��M���`�!���)�O3W���V�pSDA��B�pK,mf����c�֑6�k�cf��*�(�y=a���Y����v�3hg��{d�}�t���Y-�W`�ի�w����B�`���K��M�A�`�AS;1=T�{�sT�t��n�J�Ns �.*(!}�e�(pe!Ǘ���r�~�<2@͡�v.����[X�ej��E�����7��8��L݁�<����������Ij�^p'�y^iX��4���p���h[ݛ�'���G���G�6Pw<w+��	�Vꁌ��
� DU�r�Zܩ��(��A�
9y��qPU��Yz�r�6RpJ��4�ĕEE�q�J�Ejr���QTEUʫ�yB*+�EE�*���r���2�kN�P�\�)�CG8YVHp��QTA:��9D��*�����r��ʊ4B��TҨ��r$w)G\�E��]���QC�
��8¹\�v��p��9�֨�E\�B����q��]*�9N!r�q�)�B��AIZ�C��"�9Ȅ����9���h�������*��q�k/4B�.i�&R1bNVF�r�J�'(�G*r��H9n'r��1�S
�t�J��R:�p�A��T���*��"��8�I%��>@��G� &[�X.d���ӽ����Q=냟�g���q�2W�ܹ�Q|����ӏDɢL���wAw�K�{[]�RONHA����ӌ�����VU`���q+�̨�;�l�r��w]9��n]�.�/|$�}�ou{Ǖ��젃��U��©�z(�#̴opW��Ly��e�/�3	�z;�|�$w���k�\j�h�:�f�>�ZS��tվ�_���C�}��A2�\W�I��t���;�U���\x��w��ՈGzw(�w �f����=9��]�tc�n�����W�]%��pua���\��T8o�����w(�~fbS��5&�O+�^�rA <޹���{�+�ƁJ�T��Y55�h����;3����ɷ�G���fe2}���;я0�s�䮖:z�c�4�/���q][��x98�F�u�ۊ�L�Րj�:�X����yȇ=�wCx�	�Uʠ��Ov���3+�\"{@c�2s�u7��)�X�fgl��/�[�9�y^�f຦E�T'���W*��*L�t�_�_
��%�,�"<frg��Q�s���bJuW:4����X��?Wi���%1�Q��<�Y��^�M~\/j<�I;�a;�3��u����x��j��,ܢi��,��3m8���
��^��%n����@�+m7�6��{��l����^�+�b����[V�R�K�چ�����Um����z������J����ʾ�ȹ��|��h����d��~�߽���~�tm��;�b�\G)ʉ�����Byz S�ރ��s�nh")���\���%V���}�ӓQ�u�z�`��
�:���Ƨo����*�Ms>�Q�nuԜ��y����f�����K�w�׭������s"{��3�=�U�W�3�ӷ�jO���s���c��{�^�p��:��G��>'w�r�o���@�6WVp�wUt��7�]XN��[�ž�/��{�C�ۭ�uP�W�)��>��qL�#��m�@�ޭb'ތ
kL^.}��{���tņ�]P��>·��Sy�n�v<J#�d�H,T���3,+�5<���X{��&�N�]�5�]:����<Y��Yޡ��H/�ŀ�5b��^O�� �A8���6�>q��E��3��N�~�?U�}�t����9dW[�c�{)OF��6#���f���.c���'ӷ��z�+=�}��."�r�z�R�\׸�3�=�Gh�j����=�ӄ;9�{w�s�]\����̚:G�{����P(>AKإW5�_��<9����Tw>�d��g�V���*;#�̺��,�욕_N�w���s@4�������"z����l�Um�v&�ҴպY��w)���9���&�KN��:�̻�[zE^�D.<6�\���H��x�x[�4De0���:��faYێ�����n��(�S3��ܤ�ڿ`�-�j�͍�}%�A�:�U2�^�LO�1)�Q�s�q�tE���6=�^}wB��S�fr6�-���`tj냧��d��(<�L����5��H���/���g=��i{ڷ���3i�Ѐ�wu�Ď��8��P�*�K^��L��ʌ���謨�@�k�Juq��ws-v�fu�]�s�.k3��F�Z��s���L�w{��.F��=�l�5���}@i|}��)�fz>>=�/ިx*1z���DW��]"�����59|�.&��^�Mr#_Z�Q?��+N���푾=���@������~4a���X/��g���23c��r��E��Z�9^)H�RU�g,� �}��?|F��{�U��^���_e]C��ފ���1�0ɑ��鳴�����+�;�ۏ߫�=>_����� *�����3�gb�����{��ȹ�~j�^�3����:���@�w^���\5g���Sv�/�ﻲ����P=P�$*O����H^����]F�2W��Z1-w3�-��4�z�o⫳���}=��ˏ�g<�AC���8�f�R���A��18�f"��۸0ln�B�V�C����tDZ����<�%��jr�`A"Ebm���<�%�O>��͖��ɿv�f�;L��{�S��Up�=�uwXw�vo���P�~i����VF������gQY!�՗B�<,�ں,Nw�Y��u9�q����gc����7J��]\�������fW��L ��T+��Ҳ=��RU��GB5������үL����������R����^[�����Wg�t?R������}�]�{�'��<S�����:�|�`��'�_,��/e\�3��ov�]�V!ޝ9'���H|��NE�ǆ.(���ԧ��.UףC�vS>�Y��'/�#��W;��G)ܣ����~L�������Bcye��N���c^��ݜ�pu{�f�����`�θ:/��w�|h�������ؠ�x�:�2z ���������-�ީ�b��l���o���/����A��7�s61�W�;6�V�z�Z��}҇����FKb��&a�25ul����LVL�wz�E�u��(���uuU�Gw���T1�}�ܫ�Z�4Nr9c�gI�_,�#4>���3�o���{��7Exymf?j��2�E��W��pU�az5;K;�'���j���VU�;�z���{�Y�듼����ƪ���ߟ�s�V&�{Ϫ�T�ͥ���gs7c�V��T�WNi���r�NGWW���3�������`�ikQ]Om	=Mz"��(�;������j�K�"����nM�mu����#�kL�9;�|�u^�V/aUv�#�#I�t�v�$u�,��f���i������r�P�3Q��H��������+M�3�7�i�����.;G`��&aeJ<���u�>�g�����K&���;�Ppls�_���@���	*�V��Eef��b.��A*��n�v����F�GWK�:\�#Ւ-*����S�gN�w{=�s��ws�@�u{���^�o��X��WEuz���+��3&=�]6��$"��7���D.�J��^����N���Zo"����_Q9��񮸫���tO!xJ�u2cx�	�*��=�t�/MVm]�0�W:��/1�n�Ω}���s��PazVN_�*��ь�e�x+���Q'Ο {�X�����=���u`��:�|{E1�����ziO��o������#�l�ʮ>]��6/"�ٯ|����=	�\YL��Dw;���B;�;�X���lә��X����8�w���Y��o�ozo:.�V�§9��5C��{�H�}���q�W�(w�ߓ�PX��e>d!�Vyw��U��L͌��'���E�r�985�h�ȟpq����uۓp����B'`���o��	�~Gz@ＴǨU����R�J̒��Q]h�䕍��������o�->����m���n;��E�H�ń4
WҮ�ݖosf�_�9�����z��r�h��*C���=�<�f��n��E]��}}K���	�K\���a\n���O��ꭣ8(n�MO��bT�C��WV�C��d��9
��95S1;3�U��*M�=�#&�]�2��j���Ď�n=�a�fWh�D��í��̎�E��moY����Y3�o�����"ડ-z8Uʿ���4q��~�|3@���h�Mn=>Җj�vDtw�XC�OD�y����,L�#���D�<�A��k�gv�9�v����8���Z�s�ٹs�j��o���lt�s����>1=�?Y#��<�A��p�o�⌮cloNg��Gz���;}��&�*���`���R���:}�jv��9qw�	4��ǀ< /C��m�� ��#����.(<�|++i͢{\fs��:���g_�N{����w��	[��>�S����=�A
�v�j��X!���O�T;@�7WVp��*��#�<�YҼ��'�uv����~;�n�o&�8*SW}C&��o�1���ܖz�zc�T�/��gvוW=��.�7��vVsۤ� ��Y9p4�M�B♖@�4��r~�n�4[��'ʀ ��|q���r�fD&~.���J��|�A�N^LX�ct��ǼO���缽�����nS�ܽ���H�����hĄ�2�ø�GM�c���v弛�z������&`ӝ7��'(�y�]^���K���˾��e��<7�����Yޜ��6���j<Y��Yޡ���w� ;f��_��g-6�Ї�Z=u��U�ラ��XD���us_y�rm�s������R���Qb�;� =wY{&�=K��y��ޅЏ��=
�qD��=d�w��}���{L���Ut��S���q㱾�v��ڶ���3+Ou3Q�]����]��벥�*����-�:.N�g����qO�����謫����X�(5꩕Q/j&'ˌ���{��~���z��'���՚�ß�Fqz�u�ۊ�m�Qb��w2�C�f���ɸ��*U�#o��&���;�14{^{��|��\���'�wTdN�{�pn�UP��*eL�&hC������[am�j��[��z3hJ��tf�WV�܎��&.2f����]�j��(����M�[=�J�185���e�8W�1��.R�DV��H�n�gG{�N\r�����r���S���nr�{���>$�����{P،0��U����x������o!}WM�d�%��ۺ��c+��� A 6�/%^�D<H^���Ĝj��v���;��E�[��=fm�(w}dP�qv��:��y�.��=Nbk� *P�\�l�{YL����{Rp4�eu	�z4d�}nuk:�1�*�Ƣ�җ~������g�?D��1�4�a�����~������X2������⏧�?�
�*�ƃ� ��oIn3ټ����Ѫ��^���v���W�w�с�o��l���o�`;����ˆǆ[��ѯ%��^�}:�5׼7�ᛝW;.#��~��#3��:�_qaYX^�ٝ���/���������w�S93l��Z�&�y��ϧ�\}*�^���~8�=�<���nY�v��c>�WEw����+�)�ʨ�S'Y��4������[����̠@]�WЛ��y�Π�:>���G�(!tJb�	�X��}�[���Ҙ^��J���m3���n���n���.@|��F�w﨟#�WRc�
8���+�m�wP��Y�г,��Y��q�]�\=���;�:rK�HwƜ�Η#"$c�D���.S:���9��oI�JV���K�t�Mu��@xs�W.;��Gzw(��2��S9�f���o}:�'��V<��y{;4W3r�\Wml������냢���w�'�Ǚ��j��>�����a�5��+��J�B�u5�Vr3�h�	��4T�r�e�>/X��h���� t�dP��qsxw���7��d�Ĝ����s�{}q�=w��f�ϓ-r�"vi���{[�7gxM��om�%J-���zwD��:���d! ���js����/�H�[~��ᝧgQu�p;8�wV���{��6]Pey�>u�q�>b��v$V��G2e
���>="�z_��a�ٕ�Tj���1^���b�g���>������R��/u����8������A��MʎFA9��G��Y�a�x�+4��_gm���U���ˬoL�r}3��C�j9Տ��]�z����p]?~x�^��*��a�
�^�������Ǭ����/�l�H�]u9r��f�9z���'��9;��������M{�n$��R9��%���iR�츸��K&���;���|�����P��"J�>�· ���ڽ�^�S�۽�W�EiR2�zj2���.�E�]�}Ƨ�>�8�v����3�'3{���;�����m+��4Z����V���y]3>�=(bTAT�8z;�]�d.�J�)�\6c<j)GfU���j3�_20d�v8�P���U�v��d�3�HF5�(t��W�Tz��^�u��r󺲂�~!D��#�S��Q>F�����M��=���&��YV4�ej�����O�V���~r Z�J�Sp͹�Ù����y�G���ǜ�4�܏�A��y�^~�d�k��S#�W��F/*�W������ c��/�1�e�}k�h;�ݾ���	�,�B��u����U��wף�f;�X�/$���'��i��tT��j���c��t$;�e��ҟ��������o�(g���ٿWd�Գ�r�;..j=Ϯ����Gs�����#�;�X���lә�X��.|��^t]˿B��X���C��s�F��ؤnj3�45�8c�R�����:7ı�fbS����QU�K϶j�ƕּ�5�
'z�{�V�z{EP�eJ���FdCt'8_ݎ���']G�"^�s-R��~շ�E���3<����C��j|_D�/E��9,����y���]t��m��X�����ׇߌ��L�C���7t?3��fT4`��=0n$w#~�0�3+�q���v8q�=[���fs�O;��I�t�L��e�U�H���\����t�]����T�����,�%=$��k�1�=��*2;��3�~���C�Y)���؝���t߻j�����㓕�^�7���F�����L�y���q�r�y�=��'��V�&w��ښ>�,�]���V`�o����Uӛ�5���R���ήx��q�����FUT����~�ٖ����`y��Z��k����]O2��D��i���A���)�rVq��q1qlf9��QY��&s6�&�zv�hu��QM��7Y
kܦ��3�k�<$���W ��FtcmJݹ����3�����y$"m���;�n�7DՊ6��,p�R#��E�@BąnQED��	e��'j����n�Q�If��l������<��Z�6�[��q��Z?��=�|�2��"H+�k��q��SVilڽ��>Pm�ژ��6vQ�r�\e
r[����e����k�TT�6����4�#������^��ժ�5���{�]�r���-�� �!K<�Ɲ���7q�7�����k�Za��WW3t&��.
�����%�,eP��4Ls���̨�z1��Ĭ�Z�S#N�N"j��(n]��Ũ���[��F�F�0�ݱ亽��3�,-���^>Ը_0`kS�4t��f�I����U�.�VV�}�{���IHY�V�c�@�Pu����\���{y֎�ј�ǍatLZ��xu'5����O	��p^*�5����=�{��9@E�u���Q���ă�8�W0Ʃv\\��F�콮iz�^̹\��]R�T�N\�w8lT�l�H�������
��sA2���!)]�=�[@k2M��q7�Og`{����m�7��������W�b�Pu�vxp�-�-,��p��P���#�ᆧK
��ՍbHb�q����<�����g,��j�Y�xpX׃��:pn.��Y@hWw+!ߙ^��G���Z�y˥Ȋ���{[��q��N�-d�Y�'Vr�ub�e��!�����D��ݭ��q6����:Bl©���me�̐)zv&S��t�v�C.�͐Vt��
e�x]F����m����1��K9�i�wt�����*]�Ov��f%�o����sޔ�R���wPӹ&uEg��{R/|�E/QrO<~��I��[�5:�|���j����u�79����{<��Ka�o���r�_Z��E��8�`��9{3�D��W��49�J�.I���������G��^=���եį�1�٣���o�}Y�a�jC�7�Wp�ii�H���H�B�Y���tz"�Yda镙�ev.n\��m�!ڭY���L� @r������Q�[�]o\�4�HcN=j[����&|E���B���w��⁆�w=��o�Ur�n.�&����{[�S*�/P^7���h��fgH�I�9��)���5���ֽ׽a���4��I�^�z����vcV#/��r�]Tt��q"0,�z�x�H�_�E����+�����	S��}��TAV���4��C��$�\��=���cI���o�O\|%K%Qأ�'{g��ݝ��飮N3O֨c�k,��'w0f*�4��2�o[t:�9��)�qZ�m�y��́=�����|&U�Y�`�9 ��� 8>��
�0���')ɚ&*�W
��r�j�p�T];�8"�^sH��)��+!��ġCǀܕVy���YV�aR�S��\��n��yǇB&W�8���Rk�2PҎ�\��gu���l���*2�0�E0�unp����<rΦҊ�"�A	��8�(��<�U���4*eӊ�9˖��J�N�x�D�uǛ��0��QJ�e����	,Aet�#�I�H�G-��"
'"J�0�K*2Y&��Hx��#�f�QUȬ� �F���5ǃ˫��N�Ǆ�Rd^6NB0���J-UI$�	��%fJ�j�*<Ԭ
$�陦�mP�FNr��M��N0�5�\(�C1s�5R�.\�ef��ҢH��Qέ��$|X)�:��yg\2�L�w<4��J�W��i��]ܝ'q��=��X���E��yӸ�o^M�
�+���1.����t����3���+��;��VV`��<�²���'�\%�3�=gUt��!�p��!��۞~ǵ�_|�ד�.� ��|̠Ɲ��z�E��`�$������ʹ�� 	{��7���C�F:�:�7�ү���gϳcӹ��-��σ�5l��?!���>�e��T:����]'��@�N���
�|=�t��U�ʌ�Hz� ף�d��4�M�a�=�#�{r.&=�A�?/g��аt���뉟=ꃑJ�gś����o�.��x��j<ǹ�D�I=�!���q%���b_������e߿�T��:�|�rw��r=Ny�;/�w(�j>B�L^�T�|�[���؞�<dw��=)�E���*��Ƕ!�2;G��WN�,;G���B���Eʫ�^^�kw��D��mǺ�eq��}�]���/�(>����Ԫ��/��^����޽�w���*�4g}�ٜ����~�'����(5��U/j&�yq�r�~=Ӗ:�.2]������[���D�/ã���q��o��nU9���¦UD���||�d��2�'I  0:P�;z�fis{.�m�U��8���lg@��6.%ml���3b��ꦊ��|<r�q�}���AE.4R�{�n��2ʫ83�rs����0o�;��ϧ�;Jڢ�fލ�HG13ßFUk(q��u���k�����wӝnZ%�fw�W7B^q�ٔ�>�/��6$u�A�tk�YUBZ�3*{uӺ���;۬�y�z����,��D��gQ��]Zr:gܘ�ɚ��z u\F��Bj���r,�mr�Y����l��3�p�va�{��_B�DTo�t��n�gGy�S��nW���U��
�֕l�D����$q`�-I1����0�g�3+���zO۬=��k�)vo���G������
鐻��q�ʰ�5�C��[=�Y9qE�.#�_e]C�)����[���G��:Y�����ጞ�����������V�����M�;����bM�2R�*�y��wٌVߵb��gw�y�ˁiu�o�7�ҧ��W9ݕ�n���b�9~���WD��rށ�|:���d��["w��HE��B��\}+��� ���};�M�D�Ex楪�\���+*����̵et̪�u2cY��SA�����i�^�����z�3�%����x��� G�_w��\Pq)��zU㩓��l���ҍgi�DY�r\o�m�S��q"��ss�v��K�1jhѤFz%q�9n������ۖ�`+]s��VL?�;�1���m׳�m"�M�����b]�Z��TF/5���V��9��-��P-W72�W�K�2]l<�����,���𸵷�E^驠�o'Fe�V�G'[A�;�� �S���3�D�����HA�u\���V��_�������P3��c:#��v�V1ѣ�X��Ho�4�j4m9#�%.;�y�D��eJ���Bz��s��V\\��˭hh�mA�uLC��pfS�S1/D�=�|�g����,���f�X��%!��s�.����}[8��Gg\����G�����[t$�Iٕ�+���o3u�Iޙs>�3��4���Ǫg���ٿ�[����\wul͞�z
���v�.qʹ��tc�-�r�(c�0�B�5FG��rFK�~�0�2������zC��ڪ$�#ܯ�t�[~��9�y����1pUP�}�ܫ�U�}c#���0�eQɣ�x���>̓�(�6�y�;���}²f��!�����e.��=t�ce-Â߿<ax3�У���WNz��ҿz�}Ψ����Cc�Fl.���G��+$���'���N���'�gS�(�M�Sw��WN�oq��&�O�OeǷ��W�f��u�h�~�����Tv���jF�ddegZ�����{W��n�k¯��]�9H\m(���yuN���7�پsM=M5:�ق�����4����v��%n�\;��F��I�_�^�Bm���#ތ��צ��tz�м�w��u\�V�upj�����^��j=�y��gN��͊��z���a�����9�.�BG����S��s���Џgh���'I�,W����f�xTq[qW�z���\e9��i�ϡ�HEϸlwz�B�O�<&z�b�«sۻ�վf_<����2sz�0_�i�U�U`�'��%W��d��*�)��s�C\��n�ܥ���`��bt�w��{AO��A��uY9|*�碉�1q�3-�\�g����Vw\,��:��MtN���]O��=t�Z��=���dHk�k��A�2}Gԧ/�B��Ǻ�sԫKP�;)b��z���:����A~<x�w;����#��Qb�� u�4�rr�"�D�ɮ^�Z�i����s������75Κ��~�R0_u��z'r��Ͻ}��b|h�Mr�����Ě�c�=��fpw�E�����wJ�j>�fCt'8_����e�Kg��/��x��Ռ�s�N�~r'TQ���\n=FP��=���|D�/EǬ仈���p��<P��\OL�	sD�t�b��s��b�3�]W�۪��9�3�Z� y郑;����a����.���.{��FּQ�)��	��:���e�:�bй)5�m6��Lѹg���.�[��<V!��W8{y�ؕ�m>��`���3����"v���e��֕^�.\��9�_s���S���[��3�fnD{ב�A��}���&R�sb�{;)�|.���M����c�J���Np�+&j;���u\E�T%�p��s�I��:X.�����탊��צ��֭fs#��=_<�"*3WXa��>�&=ȱ2ՖGB��<� ���Y�Վ��7�����P�ol�2�.ßtc�OJ�L�����L�&.+�)ʉ�~�GF_�/�9���㨵���� �������=����E�p>=�R��:���Ƨk��[�g���dd�I#��в��Q�} �3�qފ����>t��O`K��p��3ө�)[پ�SeV���W��s��ד�.� ��GA�;4l�A�/�?{����-aw=�D�a�M[�{o�덉�=՜=Ϋ�V�\�a���6�F�uP�WJj���M�3țu�geєײ��-�L���nB��7���z�����J��{t���Qk'/����)[�G�~��b�f,�gY��H��O+�w'�=�t��|Y��Y�7�E�>�C��, �-���{�d�z��X�U��tt#J�}��.�̮��*U�U�}��ɸy\�,��s��S�ݞˬ�g���KΔy[�P�1mu���c��4�a�7����=ep3��3i#��*�� ෦�@0�u��ۮ��W�PbC #�ղYV`���cN3ջ�!݄V�;�������o0�"�Q	�Z�N�זݧ�d
׾j��B[R�l��*I��r���� x�ͧZu�g����Lz,�/��qlc�����:�b���k=º�����DN�#�Φe3q�\�h�p/���]���*]�R���:D��c���珷-�=��B�0;��fp�����peq꩕R��jG�7���y�zO^\V�ܹ���utEz�DXYO�=�_ݝpv����f�U9���¦TK�g~�ܜ���kzq^�������P�X�gf�.�y�����bn>=�,��0��-1�8����펬��ރ]2��z��b�,�4�s���f�5uh����3_w{� C���i+����޴V�[��GB�Dw 	������p˳�3�Nmi�+|�U�}3��Vl�q�些�g3}�+�/�;g.&�W����r9\�(Mlc��ǘקk�~�`�"z_�]c�@�qy�a=3�:#�����r�|�3_s�N��QJ�r��������p�<wpR�I�UN=��ފ�=����G��S������B����2��kg�G0l���_]H6�+�ػ���V2#���q�2W��S�_e�~3�uF�R1쀈�< z힡�v�[�x�GSֵ�]҉;H��m����/�<n�����X��s2��K^K���M(_9�����jݽ�<{92rȼ�^�f1�/���n��sQ���|�5nJ��;P���?}����ۇ7�e�������pսW;*#��~�GvV���j�OQ�pq�Duݿf����
���@��ǦW�l�����M�O8������\��{⇳|x8���(�=��=�Y��=��uՕH&yo�]3*����w��T�~���o�R��ҽ��=w��w��s�z<�]JvP��G�_wdZAĦ0��fW�l`����[��f�� �m���P}eH"T�N*�8�|�_�]I�}`��M�]a�Y��8>�]�K|G�L�+<1w;���c��$�q�Hw�s56�����p�>�zMv,�{����{=��\�������v�4�w����]���N���2��S+�*F��^��oj�m	�w����xܶ.�ɯ�����J�@�y�E�[�7����c�6�2��B�����~�*gfV��|<^�Hr��g���]o�����ճ6��#/8�H����\*�4�J�΃��C��lǰ�B��ʌ��z�#%��I��x����CU�r:�>���1n�X[��Cp]�1�L-����U�΀��ZJk+��Z�1�gţ����4�j�t3B�Fkǹ�dn��z�L�X�k�	�uЁ�4-�⬥o�Y�g)��Rb����t��<i4NmD���|�d���0��g�����AY3]޾�e��1pUPh�+b'�A���G,z<
Γ��]�mL]ȥ�}Ο�x����/��m�L�z���E��nx��џǮ�Ll����{����v��#�4߷�����!0�uQ_^�S!��#Q�v��3ܽD��~�<� ��ME�+�U��#��{�j�AOEq��*r���Ύ�F{z��y��w�w\V�����>�Hf#Ić�
��/U,�1'9
�#���.��q�禲���Ϥ${8��Ƨ�>�8�v=:�g�D��ď�\o|��I��5¾�⮽U��>^S���D�pU9�x�C����P(���^Mv�]��*�;}y:��=>ߺ�0\q�qW�X.(8�B�8�X�e�)��X���r�<�=C6וS6$"�1��t��u�w�{AO_�a'U��©�e?��~���o�s��/��LF]b���`����ͷ��z �ӞR� ���Ǿ�td6���i��ŷ�� ��Pw5������E�>�y_��.k�6���<w���ë���Qc�0�(?{s�q_��r�Z�Cuqw:�Sd��=�Ӭ]���W�G䱻k ���-{��-�JPO&��Nt�8=E/¶pt-�e,��!��ķy,��o�{	�nJ���>6���(����gG}VsW)�AH��A+��u0z�YC�	k#܆*ݝ���o�3� }�'�J�tOJ~���1t��Fs�8�Q�[#u��!�(�S����Td.�׵{Ƈ-3��ơ�֞W3c�qD�z=g��*ɨ���Fct'8a����T�O�F����/,7�_}�w�W��ה�� w��hq�B�Z����g���l���zRl��l����������Q�!��Ϥts�3��|ê����3�&eTKU��=0n$w#��9�39@p��z�ҭY�q��U�\q/@a����VL�u{��.���*�K^�r�x�3�b��������ތW��5�}���J�ʢ"�7���OD�91�ϻ�xL�?W�&y{7�rܴ�`e�#ֳ5A��S�����]��=9Q�^���[Tg|����L�z����'+�}NT���קn��*�9no3l�o�5;+�v��C�v�s���}ư_��X7�W=�z��?���ĳ��}7�Gkk}�XI�g�
7�v�YY���0^²���'�r�{?5tG��'n����3���3�;�UNJΫ�ߣ�ד�����(�r�h��2��0d���#��`���g89�㐪\s��ȸq�+h�y�V�EJօ6�����/��;�m
���J&N��q�ȓ�3jlt�� �j�9_h�Y�}e���[�U�1��+������^��>�\�Xפr�f]W�K�#4=t����䴚��`�鲺�����uoUΨ����~�om~l��9ph�l��&?�o�Ǹ��z���2cݷ�Uk7;|�����J��H/�� ׸�NT��� ��v�?g��=�*z�k�3�^���L�y�\�T�>��sܱ��"��e�k�B�Qr�s���U�@�����?'��W�? ;��hp�Y��m�'~���w�R�B�愫�{��᧹�n��tJ�:.;� ;�jMF�w�4p��=d�x�N{�c7�w��̞��姳g=����#�;���sу�7�S2����kF���P(>������zf���c�|����K��z9�ôg"0;�����}V�����p%��P�%�D�H����횽]Y�}]WS��������G��tz�X}]���{�tW]Ț��E��pfy߅L�y���[sck|o{�$Qm��WI��rx���VNM���<��}�q�7{�pn�~�n���B����[���1 a�>g�Kdpu~D,�<'���d�u`*��lcm���lcm��6���m�1��m������co�m�m��m�m��m�m��m�m��m�m��6���m�1��6��A������co���6��6���m�1��P�lcm�m����cm����m�1����
�2��-Ә(0�� ���9�>�5�#��M�*�ԣ"�&�;�D���kWM�u�(EZ2��l�R�U.�4�::�:h)Z�QTUKY��f��tó4jZԓ)���K�mmj؋j`h�MiY�)5��ڔՙ�X����-�Y�_l�z�7wsn۱�݋7s��V��)6�MAR�mJ�i;�]fš��յ*ƭ�J}�Y�ۧZ��N�.����i��U&�Z���鶥�ڷYW"�YX�m[lЕ2am5.�]�6ۦ�-kIZٻ��E��V���Fٲ�o|   wO���1X Ujq�9��w]�t�x��J�mc �\���F�����WAhwn��9�Z���j�v]����jͭ��    nm 
׷f�5�&u��E(�(�����  QJ��}}�E �(��Q@ QC���(��(��HP(���x�
((����ѵ�̶m�l�ئF��-�i*��    ޽ӭ��b��ʕ45e��{�:�s]��[�wn���n9D�h4�������f����
t��OSY�
�-�:��[7�������iZm����-e-��;��mm�ٛ��   k��3N�^��5���hl�뼠
�t+h�i�5j{�P�mm�ہE�Z��ww3]���+�v�]��kg����ֶb���W5�]n����,�k�5\+n�:�|   �������a��)�GM��$���%S�z�C���ҋ/n�fh��ӡ@�ݝOX=ۻ:l�u:R�QkdԦ��������1�hV�ol���Z�ݔ�ͦ�)[5��  ���5�e�sn�>޹�MQkC%*o5ι�h(���ղ�ݗs��;c��ͽ�U�6��w4:ضF��v�mT���UإgT^��S6E�ڶk(��*_  }O�i�ԫ7w;(:E��<��v��(����U���V�^mv=4��{ܖz��GWj7.�+ݽ.��:��Ҵm;���^���޷���H�Ol�mov����#-�ٙ���� u�zZ�����b@��鮭+zàǋ�
zt��+v�X:��q�ދcUM�7Z)�N��puU�ݞ��R�Z�)�9�tm�kն��d�髛V&�X�IZ� =�^���V����iE=1�������:�X�6�t�����8z޲��{y�ᪧF����s4�݂맻çY
:���ǔ����:��RJ�͈,ʹ�I@׻u_  �U
�h�Ӄ�*��@u��uX��Nٍ[�����m�݅6��xztQ��� ��׃�����eIJ� )�IR��x�10���L�TH  )� ���@ �~��%U4�# �Q2�*��  �������e�2�_�3o�R~�cƋ���9�o�a�>ֹ�?�B��}�d$�	&I! ���d$�	'��$�Є��$I! ������>��~�s���&/�D2�2@6��y�fe��+̋"�u8�yX��T�h#>G�R�H�;���׊�7��f �̭e�R�H��/R5r�*�x���&��uZIJ���/(��X�e���i�â��#d�(�śV͠1W��T�ݧj�zl"�=�eP�ˢU�Ѡ�PjՑy��_�9��w��J]�ցtd�@^��<bP�7�@D�qs���[���9X�z���{Q޺�%��7��:Wc눭	=σd;ɪ�\fM:�z'�D]��E(4��6)�-fk�jP$��ʸՆ���[n���ۙW�%Ә��m�ܢ���3lFU�!�sE��V��O%��5ڑ-���q�ݼu-�x�ʉ����L��KИ����
��k����U�YvQ��ܡ��d��\�.A���@��;�ٰ�o��5.΃H��4�R�0���]����shn����[��6oc�����w�J�rȚ�UփfPq%W��5	��yc	7[4�/�%Z�#tr��,���M&��r���4+��WI�4^��r�ڰ��:Z!=J�:�� �N�$�I�WWZj"`� �]�DT�̽4t�ףv�Q#Aۻr�L{��ձ�1����*ҭ�U��}��%��l�����4�b���q�����{yx*X� 5�,Q1�ԭ4%���	!��y� (Jh�E��qY��`�%���"��Y{��뫞w$ьn-[�{�c�b��䱐��F[�AMï�Nnlq��@uR�E��l�3��ڴ�!�^,�dȡd�)���9�ڂR	b;�*]Fm0Cݸ�zebЪ%�GGe�'�-��H��ٺ�`:�
2)W1��)�Tktotڴ�3-����7�Z�}��g���$�*)M���S�R�V]X��\*��4�WL^�dE$Ջr����V(��)b�B9�uojz:v�hv2��c#�܉Ҍnɮ�8�n���Q�CY*�l �X�H`ar�5j�m$�����!29We�e��u�[+k5Է����U����OFP��f��W�o��T�
l2��&��Fp��w�K1��V4�F�aلhj����i$]�%{��)��ԡe҅j¶ٕ;e��R�2l��n�&�`4vŚI�@��t�j
յ��ْiJ�� N�Tb*��o1�,D��5��Hx�A@6n�9�4:��j���+tm����"p�+� "N�p�c�2���.y���t18r��-u��"�c��0� �F��nbUy��
]�W���Yp�3�S�6���Vf��n�eJ��3^'��`T�^ �*���4���9�eYSKq�v��(J��Ш;gb���q;�~�<'v�GbT!�f���;�����z��@�sode�
u�[�p�m��nM��qs*e�+�ݢ�(SSdڅ��s*IQo&�f-q�޲���	W�e\��r�!ٱe��dur�����3V�7t �P�b�De3��#�l
)���5SjE�����:��0�%��(�uP��3*��6sܹt��.dֶݰ�h��VtR��Pf	41,ԣ�H���5�'6�|��[�R��%Xmn����eP�E��dk�c�$%m�Qe<Khh(+@��M��T�k)c�$U&�؆��!I� %øn��e�I
̺F�*��7���2�Ba��![q9�5���� �l����B⻕����2�ͣ4�RSY��,f���ʁ��0�f�edc�`]���C�5dzU����%�F]i���J��N��۸���y6ͪ��{Hѵ\Ul�iЌM���N*�S"Y�{ B¶�V�b��ģW 
��+5�יQ]��p���!�&�q�(GR�^<2e֍��^ao��%�s�p#�ć�w�c7"K��N�y�6~�*8��Yz�֙�&U�Kx�b���eYjZ(�HX�w��UڳH�$�x�*�g'�GzkC�J �-��	��I�n�?�6�Y8��L�HIw�U��Y9��=!�17�e��q<�]ݸA50\�*=³q3Z�v��0S0�*��]�!�1�̔�^Yuf7\0�.�SɹYX��L:�:��J�ŀ�G��f��#ØP��`���͵���M-�S�{h��ѰIfèک@*���`[�Dd�v��ݷ��Q��Z��C��-:B�^,Wz:WM���t�߷03�w�riQ�O6JW��:r� xfچ�]mJm+����S/a��֜�T�����l雹��ne!d��Өdu6V+���u��N+��sxt�v��qY9��V�V�d:]����e������i��j���a4J?�9J"D�&����(�����p�`�a`K
*T����{P����vu;�o+b:l��[�p�*��Wm�h����F�;��)�fV�	��U�<��+o,0��;��I
8̂Uݷ�5'�=�ֻp0rf�.��6l��à��Ъ�������QzwT8
WxT[�l�Ċ�5	�W`�!̴��f�3V��!b���c��Ub�K�)<	::G��^��:{�V�(]h��G�r���&'E�o!��zpA�Ld�K��7���j�j;����p�Vv ��5��M�u���4S��q�zk��ɸu�x�N�i-)�e�hL�,M�֓�X-��yJ*Q�l������WJL�E�lI�kl�Juc�(���i�Pid/f0����P46n]B�L[��*8�]��&1�ķe�s3�[�Ch#�j�f��9Nm[7�,
6��3$.�:��/5m9���j*����Y`L %Mf���Ju�30��%Xİ��Wza4)&7��v�TX�SM���;�&-i�1K�i57nf\��X�R۳xh�8槫� N�u)�j]7�c��vk.����XՄ�fU��V�w�"94�'�O���UZ)1
Z IwP�٦if�W1<�H�J-b��^�bZ�˫��h��$H)Ƶ1�����i0-�S���RV��R�������=ʅ���a�a���A��A�o3|L�_�]Zj*y����34���1,�@�ͥ�@K�M� ڼԎ�P�ck�q뒵l;Gn�\V� �H�[vk
�,(V|�Yݭ�ڑ��ޭȠa�Z���ʖ]�\ʲm���0��`�z�����I� �m��m��� ��id��oUU�[Wa����K�5�y��1�k����vKRTS u2�i�R�xd��Jr�7L�MW��[�
gj�T	�T[YJ��p4hk�Va�V�[(�f��V�w.�,V0lnk[��ր�v&���s�x#ɒ����D�OD�2�v*�Į�Y��k�ib�;ڋ:��QF2Q��)�ِ<8lmE�7NV��)�V������AʸX5$�#�gf���{*�d�m�K�ml���[xv٠�7nã�R)ĕ(��G��9�7�Z�b��1^��A/��]��ӗ
�G!jH!гbb���J����B�0\�$9O��#]lK�Vj!��n�D��Z�eҦ��Ԏ��	*Q7�����Z3 ǿ7�+�=��V�/�Й�aN�C�Pm��"��pd���׃Mc:�nI-V�=P#,
t���
S&�͊��Z�-d��1H5,��Û��u,�-��6����[I�+ae�3@��Q��Kd�R�Uw�j���5*��iV��xຠ�eR�	����P�L�{��Fe[6�[�i8u(�7Fc��i��
(k����V����jm�o4�3!OT0���c3h�D^�v| 6%����[�F�DgkbN��Vn��G��0�F�`�ʈ"�q��ׄ���N�|�Zb����7�9��3s�yi9r*hV�7�[�2ĵWi�oq0�#����Q�W�c4,9tUfԺ�����֗RL�52!����}g�9�������j���ej���m��v�<�5S��\O �*C�^;���e�YMR�A�Tu)I]��t3�(Z�Xҽ�6��CQU2�f��O(-yBV#�)�/wj�5�`���;���}��mɖ�ʁ��aMK9��ח2I�䈖��Pb�RR�S L�[[���k�_\�6�����·�̤�NU�D��S~yLU���� &��*ȼy�5�x�PH�osX�f��`U�Zf*N���1łj�dbrM(�J�n�P�ob�Mc{�m�m�&:صSudw`��8�v�R�}�z����|��Y�s�[6	)�F��u�ڤD�O���ۧQ+:�,jTF�Pn�5,��L ��JJ���M鱅K�u-fQ@,� �TwcVm�dW�e�-��.B�3p�W��q���fkh��]+q���5��i��O�"d�:^�_+���W%�^
�c^+���/ �F���p�(V�P\�Na�%��Bmln����|�<���˂�bZh����U���n�)�&��6Q³&�,6�[��P�Xr��2Y�m���Y/3ₓF���ܫh��opLn���x���j���XOd��o2�\��5E�8n8��.�'yV%��Íf�.��Ba� �walj��:-ʊ[Vqܽn��{�
��s  ��kt!�[���a�k7I���sE�2KF��,ң��XH�@�e�2�A�Z� C�X��q��3\.��R���Ih83wz�r���Qv�t4����;���P�4E�m�&�n<�4c�BL.���e U-��Y0D�0�P�E�y��
�"n�mJ���
7tw[��3e�T��K�����hU�	0��8��T'%e�<�+�Uw��2�SZ�X� �ya5@]ٙ�W����Gr��ZӋX�a{dlC^�3b&�i����Sj�W���9R�`4�V�),6�%\4���n�k�g}�"����������zq�=�h�㘇�AL#&:�����6�	WY���Ĥ]����X��,$kCV�m�U�jd�eKy#F�:�$-��XL�kv^͛U��7P����E�u*TF��D�K炶j���%�"KY0c�z�����{j�=��Sb%�H`i�ad��6�!!����F����Фu�7n��;,��=#Z�Ay>�{,Q�=סSp��کi����z�dڀjwLV�����R�5����8]��\:�Z��I�����B�+"�Ͳ�6X�0V����԰V<u�Լ�Q=ͭ"n��D�о�L��뎅�E���g�by�1��Lj�͉��ػ�Qe�G�U;M�H�%1AZ�zk-kwz�w� ��c��N���!{n�-���`����w���`��$�k�YgMas�e�	K�M���c��3)�,n����&v��tSQe�pY
�Tn�e�%��9a�y��ChQ��0�[5̤vbF-w�`V���h�8�%��d�U{�wi:�U͔0��% �啔��*��5�u��>7*:"+�hP/ld�8�l��S�Ww��1��;J"�U�ѧ�/�Β��Y��	q�U�W�m�}�	�Ӂ��ĄHtl�N�N�K��;�ȵ���̕��݈]��D�*�Y���b��/i��٩2��iN��n�̤�,VYoj4�6���9�V����G���5�4R��[��P�ёE�TgV[-]�eMִ8Y�э�������vM����g¦�{k� ��˥�ә�Ņ��,ݠ���nʐ��jA��SV��f��g�.��lHZ{32	{"B�dIӊ�hb �A�X�i �`@��WODRؽ�3�{ Y��5B��m��v^ֺ��Ug�Ф��ۘ�Rּ��p]�_:��L^޳3*F��Z�sQ{b�6J�Eq^R�)��ci�)h�!�4�t�B�v��ͨu�ze%���sD��Q��MV�"���9WvC�N�u��]d5�du1�i=�^	ε��T�«Y�-��c�d�r"6a;%�����olm�YK)�c����̸�ۀ��OlkL�h��Y�L-|��y���4^�[��'�^�y�o�-j��[I�°���x����Ud3$�Ø�������ƊX��HYE҅u�,�"_b̚&�deݬx1ˁ�Ql���Y!Ջ����X)F�"ʎ��̹�8�Pt���a����b��-�g��Q쐝6l�b�j5����e�n�;�� #d����Z�2���H�YRF���i�ɮ��j����G!%��{"^I�&9�vܧ�Z��g2Y$j����E0�o�QF�0�vcӕ��[�YUd^��&��8�U�衱��84��e�e���f!�-�s�A�Alݕ�Pc�d�4��>śڊ:����0ϗjC\8����EZɔU�*�˛4%���k^R�/Gf�����ND>;�TX�,�]3��]�:,�Iu.ad�� �3ofj��%]�t��t7w��c8��D@��35�0mLpdݨ"$�(V
��H�kKw®���.�C-�IV�KV٭�Ldq�˹x��1欣SM��l�*�p�YBMڍ�WI�-��X�Vܔ�ܱXK��.�D��5kT��π܈ն�*0�QOs.�u��r<��QRZ��t#��5���Ut���������Mc����w$��"�0��)�i������`����eB�lp�dcQ)Y�i���:P��ʙ�O�~�(m�S�Q*��2}zi;��5=LϷe�RC#�̵v���b۹��
�[`6]J����2��E,61l5�o1�"RE�-%
9��{%d����Z�vҧ��Êi���(��W0/Vv�ˀS'wu�6��=���'�l�8�|�gӰ�X��vl��n^SI������x^m6�F/pn�t�L����N1���b��h�f�g�k)&��lb��8�0h��%��>˘��4�e��V�΃9�_w�E�X��w�ׯZΒ�?f��s�<��i]�8��-�*����V��r���իiD�:��PU��6�4��ˢ��KQշ���OHv�2����R�V������S�i]��@�J`]�>��]b>|s"kt|)��w����}S�@ᕜ5��������L�������E�=5Y��ZΚwDH�RI� ��_`��E�����z�I{>L>�{��%v���R�b�"��|ƾ�%����s��d(�;�S6��{���,agF����5$j�"�&,�%	����e�;�/_l{�������^F��S޿{K�P o;��L��-N�נl�og�*c���:=F�L��N�oG+�J���p�_q�J��?�h�ܾ�o�~͉r��u@����o���}�ƣٴ�+��ދIs|:��Ş��o�S�扙6'>>���כ��r�\$frR_�W< �����OM�C����=�2^]}���e\���8��5xZ���1aG����xg5e���.��tL9FjTa`Tz����/j޺3�IkE�'n��)��A��Y'��o��wQ��a�C�2�_jF���)"{b�ͫ
պU��
d�:%0� ��+6��L�>@��c/y����\�3��M�e����AV�J4�S������'Uc{Q�ٙ|�6k����H�V5�����2}��9�mҾв�(�2�9hu���G��{*u�[f��O���cJZV�ȣ8Y����W��2�+!�
m�{���2:�䢍h@u⠲B;r,F��D9�e�5ݒ���{#��Rw٘.�Ņk���&�FR�(��8�A��r=W�o�g	��+���H�}����4��^y��W����Pl�c�����������WL�[܂�t@��kd��ݎ���d���פĖ���zr�NVb���w��_^��!�R�4h��ж���&#�t7�3&�KO�w=��>*ͫ��1���T�����P�"�P�#YY�FMq�M��ui�g^i�(������l���w*�ݚ�����V�uu,��,^�����{�5y�7\��-|�}�7X���e\,1�H�>ۗt�m\����x�L�Fv/>��9����Sh��E˾Y��'�)�W���\eֺS�}�50\c��]a�X�)�È�c8�bk�Χ�I�a�E��H�V>�m'z�`�d�Ԏ�\�|�Gis}B�Ƴ�L�:{���%4�J�Ҵ�+����tK
[72 ��;�R�Y�P�³.3��T�	80ҶȺ�Pٙ���u��a<mభV|pNzo���َ��9ɢ�s��P��
o7	k`O%:���)u3��	���C� u;�GlM�4�K�����8��g[t��մ3��*]Oj���Ǎ�a�TK$.+.����\0��h8*��X��X�9[kV�[�3�����dI��(e�h ���)i���W�fr$��>�L�����m>ȕvl]��ِn�	�f�vT�:����}���}'E�Z��F�e�yoM=�{UQ�T�iYn� ��wT�Qά9)Zt���jv&�0e�дt���z�|�K��k}�fb�ށ��V7H�[C����t������"@�,�'&m�
=��O�
�b*�;��r���f��aU��S.ƹt��rt;����9u5��x�RN������2\絅u��V��CA
� \MA~��z��=�6�_�����1ە���.�#��w�y�\���`�9(�$�߯����ܰf��ƣ�ޓgC�o�XZ1��%y��d�[�.S�]]򽮨R�����7a��;%DbU8�:�cl��/ �r�-�,mkJ�"�`���nv�dp��"�5c�V�vqs��\��Uml�%q}���9��6b�1�=���'\�vz��q�-(�����[���!�� ��s&�3��z���Ѻ�,ғ��P�<�/~v��Z\k�DM�͆�v�ԁ�j���<��V	��KD��xP_���MF����)��Ԧ�'�D.5��N��R�qR�h��@FM\e2��˷�0�զ�h�;W��F,�u���"��BT����u�/C�9�uv;{�4��U�IɋX�~��(P��7o�E7��8�����jȌ��	�c�s�q��#�wn�-y[D�����b�/��~ۂ��,>�A�.���"3{��5\9gf���T�X�o��S�Af��xT׺��� 𝆊W��}�0]�(e�k�˭Y��P�i�X��r��;;�׻|�,��.Đe�%�Y0d����w���dж<�2�ps��U֫(�c7����
�IV���-Q��VC;N-��_eK�3������ϟl�{2�S4�A�ɱ���|^yNd ʶ�y(�,TvU|�Z�u���Ð7����oE���x�y���޷�F��]�c�tF5�/��e',
���9ML�ٺ!I)�]b�f��2��&�ɧm�������dv��:Ɏ����Q�}'�׽�V�y�Ww�}�QHgOwE4�������7�"*py|�'�5)ںvQ�xj�&d��LǴ�85S2�Q�s�@U��3���H¹��1ȶ#Jpq[��q�S�gX��+�4�&nVt���d�yk����b��C8���{�aq���"$'��RS�#8s���h�Y���cx��8u�g�H�x�Nf`�H2X�e��(��ɅL���7�N�)��^����Bz��Cݵ�������%�ha��	`�+*��ې�dY��:�R��Q�U��X�70�4��n�@��-���>�y�K�t�"ҡv�H%8HMQ��ޗp��W݁k�0\�N�{ճy�mU�Gި�[�<3}�A�ND;��a��C�*ǒė�-���R��Z��F9f����ab�Ŭ3V���-�wma�˵4�u��u;�3b��)c%�k�����,�YLE]�BѰ���yW� �Oǿ .�������/`0�b�Z�����ۇ�s*�
T�)���]*�T��W-��);�ܜ�f�ٓ�5뱖Ɣ�a��^r�'2t�ZU�Nf��߱Q���ʾ�K�@k䮛0a1r��Hpn`+g#����ɣC�q`��w���f�V9�#۳i���@��*�h��X���6�#��N�6e��z�ǋ%e����0,'0��Ίe���G+*��V��K/�3����@�˪Ssٕq�*���j�P<�f��"[ϧU�ΰ͹{A!�Є�j݂���Kb���t�m\(gat���I��rKkQ�	���C�*�Ov�t3�B�f���
{)�c���Q�Ƭ��Y~��s��Y�wnN#	y�h�-��S��&ٺ���eh��|�8����ۍĐ���4&9�f��V���+Kkl�{Om��/�v�����M"���V{B�"���m\�g�;o�Avb��H�0�2B���;���<��X:n{��zj:���'7]j�F��w,t�!�^t��dM��r��
�&�
׬�z�Ğ���@���LFa#�5�b�N�՝�8k|��3��^v��k�t�`g\8\w��`�5u/S}l�xɥrL��U���C�\4v�ff�]�F&��eE�xɿNX�RYQz���-P����oƟ=��t�\��g���͗�
���Tt1�؋��ؽB=ɺ�����
]�!5kvb�q��]�7��+zk"�	7��]�M��
(τ��"�z {N��R\ʭ�n�������3�����%�;r�9��}�.)�2��;7�o���w�rm~�Þ�~K� ��&���Ж��$L9�:��W���727/��-����ayL+��.��j��q�5�׈܊S���0�+���A��ܰ��i*�-����j���%�}m��=`�ݰ�Y�E�
4�\�ޱ�{���;y�_ Y���4YD�LE�6�ps��a#F����Y|8]����I�e��$��//[��և�p{h��5�#6*0��C|��i�$���>����G��X5�ǣb_m�C��������3�I�`���P�U%3ByhY�\�"��T�n���4����7!����ж���sʻ��}���p\}g�Ё�:�ml������o>Glۅ��~:�����]+�#Ũ�[8�We��l�i��YG���{BZ'n%��#Z-*ͭ�.���-�B89�*��-@b��v,1eFe�-d�����vebVb��>fb����6���Q[�����L𲨷ʶb��u�H6�S�����s�1&6W�����8˲,��rۈ-z|�n�4iގ\a��5ʻ�J�����J���x"��VO-�:��p��rqt������!T�^����Us�k�;����-������I�"5҅�8��&^{]�(7��YR��\F �7Ó�9��:�ե�sVrQ4ǎ�}�w^݃7�OEj��7_f̏K�]Fiq��"��)�LCs �Ԓ\(Q�F�|�ҵ�K�B�u��ol����>�j�.V��n�K���{���}��C���ß(�;�j^a̭���8��$c*]Kku��͑<��L��w��D#9yv�03j�����%7y r�ݷ'k���gDL죷g"�/R���k��N>fnuC�;����$��yZ�]��.��k�6Uՠ�� #�y�k��o� �������Vbgq��\:�gm��#�e)��۳J�&��&���]�'+��e��D�uU�t��w ��Ikٯf�i-��O S�:ܠu +4�D��Ac�b��F;,��f�v��Ύ+2�12�8fh����%X�S�ÂXq^�5rM���^[�-����۪��@2@�=t���ܴ�c���w�𪹋C��nD.c��գ���U�O5�O���+i�dC�E��U��mK7���]��z:YfC6Y�O:���J����1����0sܦSÂ�����Kz�q�G�;:Y᧠���v�K�����L��
���wI?w.jS�2���d��1�Ph�Nm��	���-�>O$Ek3�rq��3�z�s#1g.��Ļ��J+W�c\�����5�׫���H�"N����.��wz<�A)��*�;�4�qQ�;]|HE�(�j�˷��-�;*��vv���ԛ�MN���vj���3:�Gug��̻A���͔���$C؅�	����$�P����!�P^����J��d1w�=��#��~�&g�V��o0���Js2;l8����@"I�֨�Ǘf�eZ��Չwre)㞑����nYAգ��)^E���&���Ź���^S��ڶ�G���yn��8�u1���`�Q�o+�\�4l�S.&��6�FCI:g�QnV�Yz:	�����"yDm�l 3���0Y�K�u�c )���4$�fd�Ϧ��ﱥu�엓��2��6�������ld��èFp��0�O����� �yu��˯/Q�ٶ�h%��%(�}�������L;t�3� �e���W i�1���SHS�>ܼ�;�2�\��7r�O:n!6��]+��Cz�!bcu��n]6:7%*ȝ�vBo{2Z�vٵs�C����Y�2æf��u�j�ݶ��T�J}4E[vy�ۼKs[�b�&h�܏];���Ks½�T�������w�ȇ����	��a��9��l(���Y��eY�f��s����i��8��YKuQ�m��o�����:Y���^�<�-f�[;5���φ�/�JY�8I&�Y��Vv3K�`����'�y}�K��U�̓���n	��/l�k����C�+����,�g�t��jH'����ܒ64�e�6�|Y�±Dw$��8sͶd��Q�Q����H��x)��F^ҵJ�y�o>h�*n��o8�N��0|:���{��l�]�V�I)��n��iwt�/ɻF+��4�y��i� �kT��h�@��Q�QfgYxh��.+r�N�Wf��f<�k��?�\�g)��)�ɭ�a�S5²e����\J���zaJ���w�����y����ٸ^m7�ud9-V9b�f%k��%�3�|/#�����0ZH ��u��k��3q�x���DG��b��I�O�+L���{n0���
�^#�<�_
C�A�.��	d�5����D�,��m��=��f�t��ʹ�-�lm�=�Jܧ�;��"e����K998"��Ɠ�.��oK��;��1+�f��6�i|�֔�}ǲ����=�����ogp| �X�ᄋ����5h�:>V�X�P� �{�J5}�1�FL��۪������)�x���H���&C3z��Şέ�r�'ݡ�K�]r4�i\{��ut��Ң�gk�ƶ����A��)�kh�%��-��<uxlط��3�� j��Bp�x�PLk�x!<��w�TgK��pu�L�8�汎R��>���t���k��Z=/3zݦ�׷��s��39����{�=G�`��{��ϥ�ݼ�^l��:�ł�%���!�&���̊�=���5�9ܺ�+1-��M��۞��Ssk��Y���"h�M[׶�u�X�l���.�e�j2�\�YӪ�si���w��W����X}w�[��%Iw"mRZ�1uع<���b������		�BH@�~�{��wz��E���H�q�ͤ��m�-�I�D��fi���,M9�a���*T�zllP�D�D��u"eyӱb�n�7�ND1�2>�ą��[٢�7'K��`o{>�u99�x{'m�TU:9��>�����P��+����Y���~G
*�mg:Q<�)�W��K�����^Y�	{��92�N�6��sr�[T�ʘV<$<X��x-
Eݔ�G����%r��ܹ������,��P���Y��'@���ء\�:z��:HG����/Vݚ����Pa��<��:��0�o����9yQ=�Po�6;y�����>dn���TUE;�tkv���D�L�P,�� O���:���>�E,�[[��B�g��'}�0��]�/�X�^�<�g����4[�K�
��p|#?d[��X�y??��+:g�̫���ちu�{{e�������<����̓��'����H`�4�{I��O2��W����:.��}Z��%Ԉ�**_�!nR�r	at�\d#�i]���f��m��	��2!l�=� &m��s�`sbGZ�T�u��Rn�����_�Vw���0iҳQ������2M��ʦ[������f2h
���FU4z^s_p�E������i8)�l�r���^┷u�p�{��<7%e=ejsc���"OĽXA�fr��Q��p��9�YB�����壆򄃾i*K���)�Ӻk�kcU7��
�Ы��t��h��bԝ\��13a#xr]���#����k��tbCt�/�Q݊f��e)�MR�CG�,��־D��Y�e���m����1��B8^a�$��+�S D:b���p1C���ۇ\)ij&���;��ox��z��w�JcbӢ��|k���V�!�\5�m�E��'��b�)��Y΁\�8�5��|��z�i-x��n��#(+-i1��7�Qwwp՗mR���]�X��n�S�34/�RG����	\T�3��ӠJ���X�:飵�H�qXձi�*0>�ħ�����@@�4̳v��qi;Ģ��T�/t;�����ݳۘ��l�[�Uu���8��=}�CK�dR����e��^�]�U�MV|f$�>_�({�v}}YI�M��[ہd5��-Oj��Cw$%�|Py��:���G�9�=&Y�%��وeuP�g9���d5�����7K[�vw
��lV�M4��&!F�v���%�����&��C�FM�|��<<���ݐ�u��� Ք��z:�#�Q	�MH!�����}�/m���z��z��dO��!VU�u0�J�8��I�,H+iV!�oV�u농�]&��5|�-;㒝pB�j8o�kr�1�Z��IZ0�'��E�U��D���8�;y�ܰ��h[c��0,Z3O.U��o&A���[����,O�����$y��Z�.�U�� �#0��7�������y'�!K+j��촺ڴ�a5z�"ݼl�j�'1Qq˱5�9�WY�W��G�zGy���x�	&�'�7���J̵�C��,�N+���3]����rB�����cg��}�J����^F�!}-[��7���;�.!�-�\�uv���+��mϮ��,���t#���'��a�X����
�L��0��B�1^D���9CW6+vh�Gn�bL��=�Y����l~Ćf[@��D����˭�A"�G�P����<T*�,�����7��f�6ڐw�q��򽈾�{�Y�}������ %���X���)H�qZe]fJ�q�t`�ش
��(�O>�2���|���sN1f�&arewoh��ʛС��lK��<���gㆫ2f���(m�ۉ%M<dY�BG[�+��]� �+�[)�YV����!	� �˖qU���u2��y���+V�P��$O��x��k��H����_$��t�.#�)�z7�`�vf�Ҥ�v�B�0�v7E��]����yK��']ijY{2�sc�(�P�*q4f_`�N�y!�ic��g̗�V%rߘ��#���0�3ٹ�8�o�wcL��O��1sm.̝XEa[}h�h��GQ�Г:.U�4�5S���:�7@+75���c���:�]���ΎC0�cz���j�3}�HI�oF;7W�4��z2;�
��|p}*'6�[��8�Iжc#evv��i�n�7��x�+4����<���>���ǝ���tZ���<�r�2�Éfl���}�o%r4I~��h=&8�[<�R�+4	�'1�: �_q��F3Gu=�v.�eրV���'���H�\^38��Ԉ�Q�Y�J�g-˔lVK�j��LYL��b���vp��s��lS"��W��p�2�,���xx��N�.yِLI;�ɡ�f�yV4�@Œ��)'S��:��X��6�Z�Ս
� �ݝ�A�3\��� �i+�����B�2�͏��FL-���ӓ��e��s�DEգD����^:k{*p&*�ѽ��������
�5��(x�rd#��M��Z�ٮ;�[�ŭ�s(�.|0z\3{{�����}�5 7�K�Kp�T��V��p+`nr�8�+�31��2��h��nS�*%f�ε$++K6�������R�(p�o��Ҁ��#lØL�Y�6��e�ϸls������L��˃w�m�p��)�i�!tRƜ˵�W��w(7\� 3�1�� U.$+wǘ�ĳm|jRݹm�����3%����V�V�nm�6��|
�8����O�k�y)4��;��i�V)s�=�2	u���O�ͅm	Fv��(Y��A�m��tح����ݝd��h���e�a�<�vU�S1�uю�&[8_6����d΢�p<��{C.�M�[��+���-�Y38��&<G(���qQ+�������m��D�7N��絝�r�Z���S�\z������wL3��C����F��I������|�*X��|�⣽�����ݨ�,��x��ܙ�Wh��3"应̣���d?<:u(�;­̷G&N�Є��I���F���b�Q���v�!։TVqɼ҈����=�شRc�뒏>�Z����0�C1�b�nA���K��6*N�n�3�3F뭉������ +�ͯ;{�7���C=q҈�wePʵ�f�ș�k������Mټ�lД#weP�3�����lo.�ٴc��&�Q����ǎy���n|0���5�/s*��\@�72:ȌǪ�m��(W*ʚ���VS"j.n�quq����%7bڙ���0v9u&ղ�ω��b-e�g5�8VT{�s��CZ���4Eh�u�oN;��f�OJ�1nx���4y�y�����0D\{'To�h�M�V>��V�z*��va�WW�wxW"�� �8�n*pV�_n(�ѻ�y�v�{K�424]��n&K�n��s4�l(����em�6�J��dt�F�[����4�,ԣ�s��{�HuD��Qr*����ڽ�x�۳O%f���`br���G{8;��X�WPô��4�b�ӡkw(WHUv-B��#��.*JJ՗tcƴv����k�¾�%Wv�e�ׁf\���{N����~ �/oJ�yz$�������i:�B*s�05�4���K�!�	b��I��]Qg%ؽ�K�݈�vOgj�9bU��J��*�ϤIV�,r��c��*�н���du�WA�y.����d���S��0��A-f4���y�բ(d�u�.�;tm'����Y;3�j�ǡ�y��`ً|to��P:b⯜������ �k㰔�3���+Ud�T�B��X�f�n�)�ԝA�Jm��������7X��Xm����hֶ졠�c�.�4KWw�
�(:4�jGv���x)��V7��ն�)+���A�e^_�m�N�F$qY�.8���_��O��rn<�U��e��1F�aNO����/*3�qj\�\qh�kP�h�R���{fj9hv�!:gW�{��}�.o���e�5Q����͜�Qv���|3�+(��ڶ,eӹ�3�"��vJ�x��u-��J�k�E�|�HU�dkv-iM�5`���I��q���x.aS�ܠ4T�e��M��M��7hfI�g#ᓡ�u]Aދ�����kv��R��Sr�R����)�0|��,E}|��m����E�-W���Ӹ0g�,^]�v �ށ�V"P���e|���,Eo]`���Z��W ���îJ�/��>3&Tf���!��|����l;wi:�*ʑ9Me�5�Y�5ۢ���C�N�`�@�Lɬ��8G��z��+g�����u*�e�R�C(�Z�I�4��{'>��ӂ`�dѐ�P�D����E
�	A��g��8yޚ�9�$M;�q3Vu�'\Wð�=�Vr�Y��U٣�C�`�஖���dE%�.y�F͎�י\j��h�݃0�J�p����ݤ4;J.�CZ�sm���F|�k$T�MV�u��c�S7ԓ^ឳ��8L����ܽ���M-�Bx�|����������Op�o����Dh�J��,��3�ǵ���+��V�{��Z�9�1�z:�/�[���@���'�i\K��K*aԪfnATVVX�U��R#0��%�W��M�a���mL�mm��ifb�J��E��i��!�V�$�r�*��x�Yh��hQ�Ћ�+w3E�S�c��17
�M��a�w�Wf)P�oy�;�U�n�*����5��6d�%eL��k:ޝ�`�1&;b�g�+�\	;bX��s+q��;���V����m�s���O��r���}<�Q�M��y��:����F��\=֫�1i��j&o���8r�<_2�EqT4i�Ȍ��U��?�;�jRUh���;)ִq;M5�7jN��6����b��s''��:����ty�W���xJ�p9�Q�G.��r��ՓAJ��rCKh�;�[�c<�F�-�U!�H[��r���eN��V1釨�a�d�X�戱73�I5�"�"~d�?2�c�'��:Y����o�^�L��4)<L��V���V;���3o8�,ӞУ�Tuy�O`������}��3�nW����0�}|�����Fm�
��]�m�lV� Ul��h'��c%�穢�BX�awDȯG��~9U��S}�Z6q�i�栉,�N:�k�3��r�{j�X�M�'��K�/�a��ފ���Ԃ�������&�oXm��E%�1N`�)���l���h�:9�~���d ��ͦ�ZXB��Z�;h'�#SV]n�%�q3�<��#ׂ�c���ϻ3�����
o���N���38t4�m�t��+#;��C^<�B��n�ovҐ�P%���f[6���ӐZ+6��z�C&��q�2 CFb�B��VSxur?oi!�}{]��O�V�zi���,���M��Z�phf"9�ǻl'I�=6���v�i��T�#U�5�o:��D�Y,�ɖ���`�6�P2mg�Z1|;P�����|�VBl�Qۮ2�G�ի1�]�&Z/~y�B��� �{M�V3����Γ[ˤͦ���p�]�����;�څ�,4�hN
&]�+�rZn��J����Ʈ!y�r7���6��M���rY���|x�m���.F.�[9�(i��Vwֹ�YAb�n�*�;����tLA��7��\��s���N>�)=*]��]q��2л��c��ᗋ�T$e`8)X-Yu�}i��>����$4�/�AHqm��.6�;�.RId�{��S��d��q瓪.4\́��x�=�� �a��h�	f��,wfՆS]��b��v�+WI�87��JW��WV���-�7��-Dӄi�a��hD����4��T�ɏ��2����m,�֓(��]�kŮ�w�MP�4)���$T+�G��R�Bo�O��.m��9����!�fp^C�E\�,�X�3!t}���G�W��fc�Q;G�ov�|����B"ٜ��M�z[���dX�����.�r��hƚ��&��ٕdާ�(E�����c
��[pZk�ѭ��^��!� �EF�U��S�8zx>�Jo�Q��V��l�ɹ�7��BL��3Q��1�b2��t<��"�U����3�ۚ�i�IG5���V��[��5���V*���NF�{.X��E�Q�d�v��IQ��*h�������h�VQ�"�B�O�	j����e��H��	��D��w0ZMж�����.0��P�S�.����T�,�uZ���Da�)DK;�]`�٤��t]z;ݱM��϶�n���<}�Ӵs �5�B�hǔx���a�++��`UR1q{�S��� .�iq�Y5fl6��}��Su7�zhMg�_*{�w�-���F���0�2�
ᶋ�]P�0Sջ�X��I���ts���iS!vn�z�<�_ :�W�0 &���Ef�լ	(cв��4�-�,fլ�\c�	̯7C�#�E��`��[�cSvy���-��7;|�Nkj��IaNvwu� 奪�#:6)�m�JEi�Yy�su2������Ұ���O8��{p5�\}�c^��˻!��k�D�y��*��(={��6K*�8�m�C��+�Bz]���[�Z K]�gz����ݹϵ{��H';��ڡ�<�*�3�Z�t�{�`�?h|(N������g�L�[��{��{�^
�Qoq@~�N�Fƚ7�����-<���ē�.;�$����\�m��Uٝ.�.���Vh:��2�Ѵ�U�SPv�!���=�v��qז6��r\_9���f�8h��Y�-��k8�����6/{)��2st�c��WDP<tKYM�@/�Ӣs
�f<�kxm{�_�6�Wi�Yg���u�2�`��i�S�Q��{�|�Ջ�}4�a3}!�E�>����Z}��wr��3g�ض��g|�����`�P�2�a�I�v/S��wZ��~��e_bkcM�觢��]��G�����:����v��1⸘��jY�ǧ0�b%���{秸x1��������БE�?W�I��k�n��K��]��w����ɽ�g���C@��n�Cb��\f�Y�L}�Τ���r���q-�9�9'�o��OS��<��0g$\݂�C;>�B�j<��h��s�!X��{�#�#�P�B$���:ӌ97���r\f9{^QڞR���r�`g^�[�Ɓ-����6N��XT]�^�w*��hI�/�Xw���X�Z�[`�W�H�h�
�@�\7d�x�]=�8������X¯��>�ݷ�ۘro,��oi�IPj���y����B�~K.�|�����ޮ#~� {m�Y���o3�mv�m�J(�λ}���3s�(�\q}�ЂI(�$��@Q
��Z�?�DfQ`��[b�+"�1L*"
&"((6��� �[JF$kE���"�*��#YYX����ب�-�bĬ�DF1��5��s�8,�aYe��1B�ڃ�b�TJ�jV�X�R�*�em��ؔ���IV1b�*�h�T��e��LU�Ų�V�,D��"��R�("Fڨ���Jьb+AV0jU�����0F(�PDc�*)el�J��ie��DkU��,c`�-
*��[J+R�YZ�`�J���1���,UQ��`��h�%�1qeU*U��A�bTb��QEb"��(�����Z�ͅ�j�DdU�[elQ��QE�ŕ�D����X���m���U�`��6�*UPTe��S�[QQDb��1TU��j#*E���7���Fe�����M��|�.�+`0ZBQ�E�w�V���h�z�#�FQd
�#H^S�)
)�2���ς#��w��V�������9J��D�v�Ց>��$%�P�F��oh�1ӊj�ʔ�oue��ý�-W6%*�!P��&w�������u�R�����d��s�㓏1߀�{^2�y�1a���e�Yg�<�����(쒻N\��K���u����k"$b{@�)p���(wc"��e�N��1{�r� ƍ����	[>��B�{�b^B4�f���9u�u9|'0?6{F۩��o��r�r&�G_�7��<z�v嘰����V�~H��Z��CG'�%f�����W�/���#o9Mi�����fՙ<��&z�y+~K������|���ϧ@{�A!�#�7u�3��֬L*�/$VW
���r��msf�=Ϋ�m潋�Y���B�a���(��KL>�8�ر6#ӭ
���r�R���k�b��S��ѳ��*�ّ�ں�R�sƳ�u�S��Om�1U�:�tĔ�É'�n�T��2�
�錦�
{��)��v���_]�bu�]`�1ig_|r>ʅ`�q�u��~Ǧ��x 敏M���:Ml�	�� �;-q
�Y%���吣�{z�uy]��l=T����f��5|疪ɒ��s�'u��U�_bCoY�U�eE�a�[�[c�c���aC̚�$_@{��f�����~|����x�Ϳk�ݺ
)B:�YB\��eY�n����h-�U���q_����sY��=��c�k�脛�8���v.,�)W+`��(R�D7�����}�`bs��P�9��H6�tFM	��%� �2���-F�1��ⲵ����
�n7R�\�n��RnKb%lf����T�ȶ�$V��S/�nVM����O7h�^|/���oVc�����<��V��!,b@�&C�x��웕�u�B�w[��ȡ�����-��O%��7b��SojS���@��/�oҲ��/:c�R��*Q~r�g�G���/WU�����	�;a�`�려���u����A�l���z��۽H��>K��j�Za�f�K/\<��&b��p�s>��iz��Emt�Я+g��-�����m�D��Γs�Vz�ya�*H6���y��أ#.�e:S=��7gS�V�;J����[wbƵ��6�<��p��"`�j��U��5��6��X�ߚ9/of�Í�U�#6L�K���T�
O�^_��}YN��!��k"�2���{�zoZ�GSѥ5�ٝ���8�ڗ�y�tT��9~�מQ�_p�M���e>�/��-�a�m5}��:%`��^B�����ؙ�L���T�a�yJ:�Sל�e���S�����Uy@7}ahꠢ҈�s�����J�ͨ����fkj���R�}���:�|�S�����E(�luu�L�w�)N=�=�"Tvm�	�fm�jґ�P�؃�|�9��R�.j���>!{]�ߜyw?�}�m���U�}i��J}[��'�Ʊ˵�������[I����W����/�^_xFw����W;�cU��J�sb�ލ/���89�a޶9�U�Ȥ���=�ڇMz{�i���^���T�I���a�� M�o����o.Su�ֻ�XЛ�DU�XG0F����x#�0N`	+=��,�őb*�r��[���1�o�\,���>5��Jn�*���h'q��9���.G���&m-��]�sk$�h��k*���Wu��y��o�c�$
L�ڸ#��u�V5	��6S�{׭�y��8v��r�l`�������s<je�M��ca��Q���t���jI��T��U�Y��bFlW�Z�ed��V,�i��jy��C���ʣ��Z/�	�"�DN'�hPH�8�KN��Ï�q��=�os�% �S�s��j�U�Uzӈ�@�sb�X�ɍqGs�<���a���x,�ۇ8p�Р��ʹ�P�H^c�Z�h;ۏ����]��V��a��}}4�ɠ�ͯx�ܟ.���-o��g��Vw�4���g�5����vs4-��k5��'��+�j�:V7\��J����<"�3k�(���<� r������>��ݾy�_F�7�аH��<ɸ��ھ9*ቱ�
ɚ�G)ZS�����w�^���qf�������r�J�5����ڼ#�]�{޺x7���35"p��7�a�W��<:��=�K̔�-Im7��D��;��K�h��:]֗'�v( �3�ǣ3�K���0�$��yC.q�C�_o��=�^�BV�ʪ�+�P�ME>aW8��CD�f���z�����?�ϹaQ`�,�/Z����U�{��e�J�Ù[bnz���W�Ħ�0�D���+�j6;6�SAfs��z�st�(�_��U�Gp��v���'j�G>Y}����0���[�i���xc�$6���؁�!�i'��a�4��Y��N��J���sxc�$
H�-n�T.����0�,�"/��O�zU<�<�J���ܵ\ܥT!P��VI���ّB��,�L"��~����꫸��[W��{c�w���qL[o��ͫ���g&ۅԎP�]+Q�*Wlܬ�ł���y�͉�^�nLQּUxj�F���vC�J�eY,p��/�pJ���˿?��K&N�ɪτv�[��޷A�[����G%����v���Om���*�Oz��ru����{{vB����	ь��\%�R�L�R���qD�ʩ"��wu��ONPT�gW9��Ii�x_�z�r*���E���A�1qX�@2e$���VaL�P���;���8me�E�k1���W��\�Å�;���$/@�h�X��h�㽊	a�h^냗���l\ٹ�轘�о{U��]ke��H�.}��Yo1����מ��țJ���3j����H�Ë͋{$z���Ɔr�9����[O���ýc=��<���ոR�8��Xx7��؊:Ы��g)�+Kw�nԮQn"�s��iu�w۷�W�ݸף����L�$x_=姞���s7Q�'wi$+%�Gvgyͽ�
�PQJ2�a�[�[~�4��֧c��Qs��5Y���g���ϩ⮅�~�m����*ބ��e,��Q�*^�Be�,�s�]+v�}ttC��,�c:��	�@쐰����;����k�F·����z] Wm���5l�NlK޻l(�U<����K�%lNL��'ն�a�:iJ[pMqSZ�>��!^߽��:+_.W��f(}Z�jU�;����i�H��v�֍[+k#HF�/����������Ն)i�T2XY��)٧A�g�p�ژM�Y]x�����^�uq��� �o)���ۇJ������(hxy=�b��z%��Dy���sl�c��lz^钌Rѫl��Ց4��S+�a^[*k�N'�p�r�����;.����=�J:_��ld���x�e�<hL�ɱ+'�Y�l�=˾܋�&�d�U�]����~*����^m�uNʲ] xu�r�f�f���݀[3o��=�a���F�>\�H�u!]�a�$q:��+�<:�.n5�v�÷�-s]�
ۍ���y�B�ح@Ƕ��X��h佽�R�h���ۨ��ݧL���X�d�\*�Y]n��c��]�gV[҉����F�%�u�H��r�dK}n+�sbi!�A��ەr+)V�uE�oנ{"WӮ��ߠ�_���uy��m��tM,����˞�.���w|�r�`�/8��9�I�'���wrש�'ov«��4-TZQsb�Em �#�'gvu�SCqiy�}�U������;{���2��6:�b�t��y�H��ש�<~�9mAQdBz[�"{j�܆v�X!�WP}+J}v*�
!�3go���{]D�U�+�>�`?:4�Ń���k��;ޛ�*��l�65t&l��ܑ�� �+��;"5�T�|�䭼�,O�3\�ep�vu�[���g??An_n��Sg���(q��R�ih窏-��η�U�Ǳ1��Dh���,�Vqj��z�aGw[�[ss����i��JkqP��X�.�p�U��d���IX�6�^��e
	m��������݌jk5g-��y2v)\w-��i|��*~�5P�dM$xPp��5���:��`�5�:��`�~�mgf�y4���V���]��P�dRg����b�eE�QS\NC;�S��kQ���OV�nG-V�K{P�u7dȮg�2�$�v�qq��X+��k2ZviC�߷�>�-�o_^W�����w�R�L>P���Խٱ/&��{k"18ޤE����h]��5U�1w.�{���n�xu�j�p��W�U�N#7��SS`�M	�g2��of>�S�_3���i,8�
�N����kE�R3�ؗ.OVX�v�SWhD�"n~�Gx�����W��N����2�����m�Q��;�q�=4n�)ӍqY~W�w;ϸ�hc��ӡ�)�8M���d�8/*��Ť;� a\�K����酆�a�shf����G��S�P���.���*є�c��f���p�ך��J���{���ֲ�D)�8?+��Jn��F���u��k;m�tM�8���Ļ���Cl��]W�'�[F���~s�n������q��߹��}}��NqV����j̴�
���E�A�_&hg>P��h6��;{�yv���ne��y��6���/]�m�]jem͈�L��pϷ�u9�T=Ž���	�����=.��U�պ�Q��]a̭���z��仰ʷ٨]]� �u<���q�՜���z�uy�t��!�-�D,�գ���P)����ez���͞�t���Mf����ʗ�������������]j��d�n��n��#U׎��OGf���NlK޻o�vE$x��l܌yW�;s���W[y�uke#�[�@�{`B��-W7)UT4��n�a��Z(s��j�ax�|�!���WN�ǻKx���]����]�˺ыk��aC��~��v�����b�f��񭔣�����goS���A��Y��O3��,���b[�iwsA]2]،�c����4Ȃ㡒t;[r�q,����٤��?��~�"��,���hR7�S�q9w��ANÙ�Y�[�:�1����)�n#ѭ��R��+��˿X�(�[�1?b��[�#�G�xVK:�9}��V�V*�Ƕ��͈Cj�BGSҶҝȇ䁅ɊH�49 7u4�vxm�=W
�[1�^��:�⟾���߃�b;�;2�Z�8��e�4�=6���b�ÓM�\�y�l��8���5���Yl	w5��-m1��k>�H�Y�w o����Eմ�aj����.�ݍt�MD�c5͍����B��B�r�st56m���S��c��*���t.+;�觎��M�O��({�ߨߓ��~r�M��K7�Ay�l+/�Sck����t�9U�y�q�GO(�4�@�L�$fa,*�����^�s��.�ik{�������<��ov¬U��w��V؛��T_d1��v�B�]�Ш�=5�E�VВ�V�p�lj��S�!�l�q�sG'<2=wv�ڗV0h�N�p۶R�]���q�rO�|�;������yi��>A;}=v?h��'n�e��ƀ��hS=�;����#8�vp�����^X��u�!�A���Y��+�g�����[#���Yp�f���:Չ�U�Z���a}t�h�b�޵�ޥgi�)��.?<�q)R���5ك��K����3������th~��pY�6�]���2yY�y\����Q�>v(��E����'q�9%m�q���҉ݺ�J�
9)������j�Ϸ��J�G�V-�O*}yCn�!���8_���;��N2��t�b"�:)�7�2����9�@_�lLKOw���S��n�d��P$�u  �R�Z��-�̰LK�""qo5@&�u�4���?� �c�n���9D^3Z���!���FeX����g�[ؠ<���׬�����b��<�6�}�����HKM���}�Ϙ͸��Y�:��V�j^���I�1_I��ޏ>�#����R�r�թ�9��'ZU��	�e�TK�F�=Ee���A&��'s����+Yީ���u��\5�CvA�=#5kH1Ӿ��5��;$�蹹^���̒�>�k�H����qA��Z���*��M��
}�:�K?-q�<�(.[���(�X����ɡ��f��4M�WL��ᱵ� �7\��� �]�&��iyw���}was�&C1ʆ��Q�����Z��Hn��[�����x�k��J;|�SV���(z/v�Uיe��gbF>��w�q�|���+��}k�"k�vǁ��­%gZv�t�2eG+��Q�J-��x�f�&)V���%c2ݚigg����-j�xG���3l��P`vR�T,�����Rq�Sb��0`��>i��8��٪q��J�d]֜س���f2�e����#w���G�D���k�x�vݜ�t>��jF�;���eҰz��v�9�,e���-�qɫy0J�������Օk�q��J�r�i���8F���5����0���檳�}������C[3:
[�_r��2璭y�8{2P���.ݰH��A0�H`��g�y+����:�2�U̍f	���S��+���9�5�����:�ݫ�1aZ:�'�ҩfS���͛8������P|���޶���B�2�[v�jK�&{��*���V�F�9Q�'����|"i�Q�|��嵐X���op��_`�I֕�;jF��}�v�g:����^�1^�
R�Kh�۟v�8ңJ���k`6)@��+l�N�o����d2m�ױL9]�rbX��ĭgEё �I$�wy�]w��c��,�>ם���y�W��W��[͇"�F��=9��9Z���>�����C� R(��a�b�j
\a��TQDE���PE�EX0�-����R֕���)R��EE
2�*[,eZ�eF�b��,Ab�P�U0Ѵ�֪��X�*R�R��-�kib�X�`�[D��DV*�+m�U��X�m* ��kQAB�Q�EQţQ��jU�Z����Qm�V1��XU�����j*�YDb���-�PUT`�m+`�+inq�pجTm�J2��*QmDV(�b�ŌE-��T�+iQX�#ڈ"��j,X��aTV(�Q*Ҫ*�+QV��Ŷ4���K�X�+�V6�jTH��	hc�DTWiQFڪ�A����(�Z���`�Ѫ�%k[V[E��R����Ä0�T+�1X�KU��-�UTcZ*�������,(�ʵ�J��+-+aHT���5i\\`����[kma�P\mQQ��+UQU�֊���(,P�����1J(��D�Qf���R�ԕ+**�*����H�
"VKiPDKj*�R�Q��
10�V#�I���ԬZ*"��)YcK,-�Z��EB�l�EUF
��	�'ĀLrLW<{$wP����el�i�S:�s{��D�b�ڭb�W�R^��*��V�9^��Ź�?e7��R��,;���?Źyʞ.+5b6Ʊ�^n�2��K���7.�Z��~�3�%��=�};^^%5��S�lr�b����in{�v�8��<���j6G3띎b]�w��f��9�/z�rl��ݫyiw�KwԎ
JH~�GM ���d�"��׶!^�wYm �`݅9ݺ���HU�L,T�
�7De&x����m�5�1;�G�Ȼ����u���-L>N��-�t���Be�M���;+2bb��c��V�RY��]~�q�5���B��x)���uNʲ]xnd��E��B����/�r��붅�*Ǳ��ԅw����N��Xm�k6fy-���7���]vq�,���nw����b�c�mV)
3�%S����2M뜑���Ր.�쉣Q�^��~{E�f=b��3��p�_:ѡ
��栝5{zF<,��"�Tj�g]$�u��I�y��/mM��v�ݢ�����Z4�:-=��rp�t3Se<ř����6^Ui)���̚�����8���d#Bh�Ys+�0`w4na�ǅ��R���zޚk���ۍv	���{���V�Ĵ/u������+*�O��ｹr^����1���j���^�"}O&/vz!Ӆ�}��=+�j/-���.���Xc�[��oy�S�t�8*���mh���ek�.�]�
F�<!�X�z�#C9�-\S�{�ίOfNs�.0����&x�u���DxR��;�6:@����#V���9oZ���Sv�ۅ]دz��&WFP�/��@�4z�*��i�������������1�ή���c�V��(W��=5C�ܡ�ۿ/v$����8 �7���Φ���%s��]���I�i
��dص��f��&M�ϝW[���L<�Cʵ]\��݅��>���]� ,Z7bL�H���񾜵WR��m�8�mý�|�S%��t:�ݓ"���>�>��cLý�
��%��������1�����3oЛTð��f] $Ɋ�4b��jAO��v��Hn՘�xƅ�=w:L'iŢH(04�w¾2�	mz�:��v��:��j���f�+9��Xy6�{1;�*Q�����F�o�Z�}�m���r�̈́�&�3V���g�I]�3�y��0�!��@�Cl?�P�`l�q
�Ri��	�6���г�y��_|��G3�׹�N^[W���<J��z{��J������q�?9Mf�u��Ψ|�$�j�l+�&M^�6��3�Y&?��L�@��mτ>>��뭶��m�{����w�wF�!Xe����|�:�E���ud�9dY8�����<�ԛ&�l����2�	ԛՆ��|��ԇ��0���� =� ������X��|:���;�vc��6�������d������6���`�I�M��%ݒy�y�)4�`|�!XI�i���4̟Si�̏^G��4��� ��S��h���z��J�R+��u�������2#Ҧk�<��|{��I�O�X{��m���5�2L�|w��%�$�{��M?����?3i��Hi������s���P�J��R���$"=�P �q��$�a��ɖI�|~�'Ru���]��O2~$����I��������o$ㄓ)���E�ް>���jK��뎮�ޚ�
#��0�H�
���!����|��O�@�d�l'u��S��I�|~�'�=��jo�:��N?�o��@����k�`_�������s��k�5�c��x�p��N�(y>Hz��C�~f�l4��g�2u�I�O%N���a�9N�RN��~��{vG����I��&����9bEˢ�o��Ԭ_��d{���a�s��<�B~CG�bE3�f���Y'P��͆�RL��u'�Xaĝd�T�!�O0��u��:�������=ܫ�'{���`_>�����}$���&�{y��3S�k!<���!��Hl���$�5=�e�uɠ͆�,��aԜe`oVI�N�f�8��"���4��M��9��Nv]q������[tB�D��W9dfH��ĥq�_u�e�2�<��&qBMb�b�j���b'�����G�_�G�$���l�z����Ydd��؅��6Y�����y�j7�T�[u��6�>��I��\��r���IәK9����7՛�w��D����>Gޱ���z�h��,0���_��)��}�k!<�|wd�d�s!�:���.N��>����$㎝�1{��n�}�}��9߷��C��YKC̞d���8��>M��N�~�py'�L�}`q�̛�"����~�d�(L��<�d�Z�u�i�������y�<9͍��z��G��a�{�6�I:���;��ݡ�N$����X`y�So����?0�y	��}���4�S��Ad�C��Y���3ӟ�5�o���烾m���y��
���=��$���5��u�l�5�u6}a��{�Πy&��51`u��?}<��y��u4��h�p�|�>������{8��������tI�<{�̕*I��c�*N2�cO$�&��̈́��Hy�'Xo�I]���������!�SN�k�����??hǱ�u�����>]����$}� ��@��8������a�^��*T�ܾIY9�8��'�M�y3a:��Ψ|���C�+��ίY���ߵs�۝��_d�\�_ۯ���xa�d�>�Xw��C̛Ag��T�d����I���d�RO�,���߳�y����#j �>��\gO����j�O���ߋ�g����u��'̇�v�y3m:��*k|��O �>��!Xy&�P�i
�L����|�e��wy��d�9dY?}`w�O�3�>��~�+-Q��p�Ǯs����xi�G�@Gȁ��j��m>B|k�$���PY%M�d�T&��M��Ǫ{��I�M{�m$�y��a2�>�~������}�s�>�I��m�`i�Ι�C�&O��|��M0�~C,�At�i!���1I4�����N�Bwvi'�7�O�� q����4���ƽ�3'PRs����ˑ�!�߫��yg��ww�j$td�s��atW<'��ʍµ�=�B5eOAn��7����Fu�u�<���:WN����3�h3!6XT�N��y����rCI@�^��:<4��H����w���ދ��UWQ�Hb�z~�=� ��m|d�z��w)6�`}�bi����C�&SL�'PY?�m2u�t'u�,�e�i��O2y*��&.�����h�����=���Ͻ������a���k���I?0=ϰN8a2���H���`v��!�?3	�44��1��2u��VM��O2��t'u��=��C���g+����4�z���̄}�:|<���O۲{�'P6�o3�	4�������'�4{���|��w�I8�O�CH,�?�d�V;ӏ{�gz�^�;����ַϹ���2����P�I�=O?�N�峩<�����2k�Ğ`~a��~�a:�����H{�E<�Y?'OgY'P����<g9ɟw��oǹ���;���+��P�'R�>IԜd�zn�u��3>����a��1:���[�I��'�X,���{�b�\�8�2q�c��~�5x��9�������u�IR���i=��Y'Z��8�!�P�'=���d��v�I:Ɏ��?<a=���É����|	����ŝ��)�H��U��;���*
���d�[�8�l�
IԛO�q0�u����N:d>�:��Oڡ��C�a���I�z�9@g�=Gx�����J���ϼa��'�{RN��]�$�(Lϻ��+'䬞��:�l���u&�?Xq�'Y���<����$��L|89��7��.��_q��ɫ>��(�6��|���<�'��&��dI�>{Y��Bd��<²q+'�9�I�M暙��d�gVjHϪ���:}�y�쟻.k|��f�����)?<a�Y8�i�4�	�ܧ��>d�9�bC�~d�� ��I�}�d�RL���
�Ĭ�g8�̜dځ�g������O�v,��6��J�M~�D��z�b5I��^��P�x�����������Һc/����ؙ��pG��c�:��O*���̘�=�;4آ��1]�!;��c�M�����)�{
n{�q�k��IAS��GL��.&�A��	c����괮�{����I������d2j�`m��>���d6��b|��)�{�T<ɴ}�bC�?$�Ǿ��$�MK�fJ�|=�R<O�����zr3f���SZ�}&�:ɬ�١:��d՟;I<�����q��n�!��37d�I\o��$�
C���u�IX~;���#��Q��z����Cc���f�9۝��Ǥ�RN>�H���ذ�$��a	�ɖe�	�Xm��C�W����a�~�PY%L��̞>$x' a����D��'奻S�J���s{��5�&Y<o���L�}�o2Wi']^�E&��Z�ğ:M�i�L�M��'|j���>d��&��>�;��w��v~ߖ;��w��̛J�{��i�?%a�w?2~d���s�&>�����)����0>=�`m�����!�CI��m�$�
�6��:����k?�����{��:�z�w�L0�=N�)&�����N�d>���y���&��6����{\����sy'$�N�ȡ�u�����Cl?&Fi0�־��뗆����u���qޡ�� �~d��Y?%g�Bq'���:̤�C�}��O?�O~�@�O��w�Ğ`~I��~�I6�����q�	�����8Ϙ�ߵ��������n9���Ͽ:��!��g�44��`��d���8ì�JϷBq'��;��:Ö�d���8�䟞$ߵ��=�<��}�}|�\3�~�����<&O���bE��N&��I:��k44��q��Y<���N0�'R���d���߬��>��ԟ��`�'�|G��=NT�]?P��m���d�����ӿo!?2��u�I���P�'���pe$�ɬ��2�q�ŇY8���T:��N�CF�Y:�0���I:�5���ǯn_����W�y��De*�ơM����ާ^�LGu%�ПP��MY�m�U}�g�6`�{q%�n{7Q�5� �J�e 0&؎M���wl��+�1E{��������ۄL%���%,ڟ� �Y1���4�i҈��=�:���M��)��o�`'Y��'��:�����d�~�d�I��}C��I��b��8�!��:��=��WR��sKr�ڿ�]���}�e���x�q'��'����{��u�2o�!���ؒ��3�8�d��'m�8ɴ�`�N��|Ô���D��/?&o�歵&Kپ~�C�ԇ���$���8�������sg�:�0�?��<��M{��)'P�ߵ�*
'�ǒVN%d�9��}�#~�!tk�c�����i�	��I�zP�J�����6�CX�:���<��<��u�I�o>�O!���{삒q����G������ˋ��;u������2u+'��̛d۔ћ	��i�Xn�O!��I]�2n�`m3�|�Hm�>Bu���T0��kr����ya��4��5}6�R��O̓����'^���t�ﳂy�?9M�`m35C�i'P�Va_!2j�!�0�!��:�y0��#��������t���������=����P�&X���$+�d�5��Iԏ~ė�$�瘑d����y�6�M��y��3>��'R}�����!���O��ѩl�V]}G{/_ܯ{�۫{i�޲#ނ>��q���H��I�O�Xk��
�l�����$�d�u�.�����I�����$Ӵј��>��H���G�-'d������s�_���﹯CHi�$�㴓hq���
ISA�X�I�VC��i<��+{��'�Os�q�e���$���N��)6�`z�V��6���^���ώ�����/���!�<z���'iha'_�T�Hy��ɆI�4��ԝed;�4�̛v�ݠ~@�����x�~`h���N8I2��?�w�����I��᏶�[��d���s��I�n����x� �k�4�U�Hf��C%�2�z, )_Z�@��A�J�쫖j��=��mY����鴂�Q$[�C�F��%g\fH#�I��Hb�gW|out,�4�-yG��b<�Ь3T]lIݷ����UV7�ċ�`���Ch~f	2L�Y:����hy��_�a8ì3�u2�4σ�q<���[��y��������%��8��ֹ�`����WyI�����|þ�fH�}��'���bi!�?3	� ������'PP>5aĝd�T�v�<�"�Ȣ=�|/�2�����j�P�
����Z��?��5�3�"=�O��=�>H��߯Y�����a	�?���8ϒq���$�Oٰ�
I�?���+�Xq'Y:�4�u��?g����r��|c��7��p��I��0q���&�T$ӶN�$��f������L!4���C)?3��2�:���l4�>���Lx2<���
��Mw�Q���驼����އ�d�{�C�����v�y��{�q�	����8�o�M��)��}�k!<�}�}��a��,5�`�H�ȌG�φ�J����}'2�'��x*u�u�1a�Oj�}h~d�']!��@�&��'Y?g�<���&S]� q��4~��?!�}�k2T'�O!Y:�Ü��������Tα�go����y�m߀����O`�O0�3�&RN��,?2wVC���'i��X�:���6�a:Ɏ�����NL�@G�G�ﶀ'�� Z�}jpB�W�������}�:��	�{T��Rw��&Ҍ'�4�P�Y'S?X~d���Πy&��4b��H~�l��9��u4��z�|�{���ϰf�dwq5��i���]��������I>��J������IԜdۗY��@�i5���P�J��:��>a�b�䆐����o�N���1�o��!2�����a�:���y2}�}���a�{�d�RL��<��sv���y�����̈́��:���>�����w}�s�iÜ{~�t���#��o1�R��؞Bw@�יtk�BN>s�y��J���k�(,{ȴ�;���V�|q��;�]��p�b�g�ε�]fl�G��dR�W���u>��]�������^�C��Ŏ�^�S�����h�9�{�ZH�)���H��m�4����=�|�����|ŃYc5~��Y!����8�_��̞A`|w��C̛Ag��T�d�=�d��y���fJ�$���H�sV��	�DG���<π��1��f�GVVn�{�a4�Ӕ?0�u���C�f�7O �J��0y��,���+$�*{�!Rm�'���0�d��w�+�I�1"��V糏�i��������m��@�OΙ��04�>���'i��e	�i&��~��PY%L�2u*ݳI<�l�~�pB��>�o�\G�$��~���SV�����y�|�ǉ^0�O}��0>�1
��;f�Hu!����>Bq'ڰ�~C�N���$�C�<�$�������Ȃ�=�i����=H_)��}x���-޵�r��~��L�x��g�&P>~�I��	��l�M?���M2C�a��!Ԇ�?Sl���,�jɴ<���t'u��&Y&���ֶ����ߟw������Ƽ|��*��~d�'�Ԟ���&�m�=�����k$�)�����>d4�ل� �Ln��8���Փl:�̩����=��K��7R�r���#���"����Z�	���M��y������������M0:��f����E�,�>#����}�u,��x�j��	��7�^x2��V�I�'�q�>��N$��$�a��bu'�����I��'}d�l6�N���u!�q�C��hh��"�C�N&�`�|������]w�1�s��7u㬓�i=�1I?9>��N�`i'u����vC��a�����C�}y��Ρ��9s��$>Ƨ����q�����P��ms�K�5P��+�z��+x5_��Fh��:�2�^�i�Y	�NeX���tiT��!)���'et�c4<KY�dk�R�ܘ�>۵����ȞU�᳋�U��!9����yK�K�/�3�>�(Dcfa��n<n������7K�P��[B:Nm;��N��Z7��,����|�ܗ�;nĉ��FoG�B[b�ҋ����Vj��
5�b�r\].���:�
�KW+�tE.:w�R��qU��7�͵D>'f�_v��W4�'^����)��v:��$Rg�zevM�Yl��l���o/7��{�6���2���[-�C���|���7�d���u�liDz@�y�ｑ��{���G�
	���ڇT�%ͥ�g����wZ:0�n͉y>��W��ض"qΤ+��5��ɾ���C��u�w<����X��kc�6\]S~�R�Ob��v�fn��̧t�����}��(�g%m��K0�n��.U�O`򐱘�Y�\�Z�n�N����Ж)��c�I{��7���h�LYԋ���D��C����l�k\��ܣ���{���O=텍����r��	���RW�u�!��2J<f�Yb�]�Z��,�Y�R;}sg}��������c�e5�gmn��Q��/.:�S���O�f�#�u\X ~��{4�{�z�L�u�a��s
�h�)[�g%����c����F6���f��؍��r�5��n(:{�=�j�fxz�Gx����@Ҍjy�rm�(X�� �Yz��"�����p��j�^*�,�WV��EN.��.�ws��}�l�3�ǝ�r�i� �޹�[
�tܠ��$�z�1.�. �DZ����f�CH��e�E\�xq�ngv��C��]�s���1)��H��c�w+��#���Q�zX7R�燏r�[��y@��A�j2�����=��e닛�{�p�9�uMO��P�}0���g�m|O�����@�p������){O�S�X� ��8�ڵ��dr��X� ^ˊ���]����̆zڞ�������Y�msJ}嚧U�{��ܶZ'8CDј{4�����]p���퓂�M\G��9����X)x��7���r�C��]���<!�|ދ1w:�Z�Ֆ���� %6�Y9��b��a��#�&gt$v�{�ݮ�1�aD=��M�v�ռ�R�f�+��f/>}~�)�=2�m��=L��؍\����"3�v�|pU�L�Iy�Ţ���8j��:Eı�|����\p��%���u���[��y[�s_pqk���u��)�yd�lѼ�[ۣ ��[v�i�3����|��ղ�<�5�N7�'+A)#ߣ��(�}»���|�m�:�N�3L�D���xr�r����~�+��~�̯���� �t��'}���o:��G8.�����y��9r�����'����펢�L�uuB�9!Nn��%�8c����Wf�Tl �*ٖ�I�d�+)�9x����<�v�$ �w'���$��U���E�G����/����YV���l�����}�-���on�t���*a�e!���s�|�A���y��O��~�g�&q�B4�c���=W�����;��a
�O���t�q�S���E�{_�t�0i�ėa~�����������Q������t����'�0ݾ�Ge�J�l;�#�}i�:l���\�m��+�+9���Ba|(t8��4�u_N��Ř�	1C��y��f@@��YeK�h�h!�;�%{�q*��u�`�i��"Ժ�@nf�LY���X���O�ۃ	�ʖ�MJ��G��(o_��-��f��C�,kq[Ԍ�B��s<{9N����"�u/�y������H�V�C幋B�uL�JN�=S�wm�/����uwu��>��񠚽.<�P���K�U�Ӵ�v����fMژ5j:ev��� �$�	��AA�AH��l��DE��iP��KlR*Vō�ł3h*�%a*�SS�JʅJ�EeE�B�Q-��H�PcT�
")4�$�Q(,�%�����E"1Bڱ��"�- �������
X4Q��T3� ���((��H�EPR��,�F��D-�REU������j$R�Aci(�X�R���$��A�b�+��&0�b�D�-E�U��Q�QEJYPP�*��EUEEd�����C�����QE0�Q�X�X�"�H�Y�-@iE�U����AKKX�
�[E�UDAdb!iAS�F�*���H�6�+AA-�#Z�m
��&��E$X5dR#H����,E�$W��%�`�(��Q�YF)
�AAb�AV
�T,IY*	Z*
�DTE���Y%eAIX�m!E`�
�QdX�DUF*�1eÈ���[Z[j[TDEA�mZ؊l��++X(�b"�EX(��QPP\�B�����!PTb�`�b�V ֈ�V�"(
*�(1J��TUE+>#�����ݬ��ڗ�#�)X�cy���~r���
4�ɂ�Q�Ɏ�7X�vz�0C��S,--.e�R:�Cek�T�w�����"�b��W�[�bz�<I����)���N�F�8������Z���
`����pZ=+�-��V���oD�X9��N	��[�����[A_D��5�{������GBB*�r4>חx��fpƸW��SL�|~�vUsL-ʬ�Z��q�L���k����
Z;\�VL�=�9Ε4��p�)�u'�fג�c���\����<���M�ɳ ��Җ^���Z[�E��;=Ή��)�����\8J4kE���Z�^{d,��"^�^���[�f��P���f�>�"m:�3���ו շP�ߢ+bĈDu+#9���S�G��Z���*�^�����.���a��ɳ��#�-��ypZuD1
���CvVZ�m�<�L�r�+�h��y�D����%H�،5�͛��9���:R5\�r��*
,vԹ����5�3w�H�DX�T��
�v�N�#B���&��(׻�҂G��\��#�hd����t̑ň�&�r��>�/��~�J�+	:���j!P�2��>Z������qn�R��z���H��>���X��"Ҿ�/֯���	�-��g.��/��cݾ�W��Ly$2��5�"��ȴ���7��8��f7v`3�j&���z���}���\]�}�<��s����^V^!������1�)��Y/�l`)܃����%���g��K�ef̖u]�~�=�u'�\��F��Ý|�s��BDJ�l+!��j�鹘W����,i{�ȉڬ<i�٦���d=��9����wnP:P���]��o���~0�9�=6fj�/|��w�ZoIC���{=����(�������N^s$]�H�����ܥ_N�Ze��h���t.��E�Wz�
u��|-�pu	���`l��:���<�o���'1Y��{[���Q ����(lҰN�6)���b�B�yu	��������&��.�V6�a~mR��r����O]m�pkesN�TR���ı�x�j8R��m�>��g<�:PMWr�lk���P��3~�w's�3j3�f۩�&����^�o���h|)qh�1E{Lߔ3�,k�H�"�po-�
mܖ1D��Y�<���EL(.w�D�]F��GlL��G;�!Y�ҧ�h�9T��~�w ��D�s�3���� �<������]+�!u�������t�D���w�B	iD�p8����JZ4�[�U��V��4�l<U�z�����%���E�=�g'�+ɗp�Ze�F�V�f�M����3/�9�w�c�ϔ�����{Aub�1s�����	���ӱ��m��xc�����T����\<����gz����v���c�|éW�w�9 �JANq��~U-Gd�gnC5�vo����^]ĐV!��]{�'�V"�U���8`�c�`;�{CtG�ṫ��@t��Gg�kB�wx��Z�Ç��f�N*��Խ �@�~>�R>m!���J�|���{4=|&�oZ���}�����^=T���hn`��]Գp��!��F�R/�vQ�ܶ�d�oJ�<�n��dn)�b"}�H��-D8��j�9^�����(��)<����m��c9���ϯ,H�re"��7j͌S�3�"��$����~�0q�e��ӭ����s��t���p�(m��b�G�f��{Xl{<���=�@�,:ne�.��Ԇs�1b�9F�c��2���{^��|5x���u�W���A׳.�~+Ђ�x�w�<r9'��t1�Ǣ-)dgu�v07���X��=�ܺ���&V�*OUu	�n�]���s�:�$+:�P��[���уvʓ2�ײ���%��_$�G5�QUH��nU8٭x��Oi5�߁�ތ_T����:����HfEq��)v�Ew�N����k=�/t��2�а]p�mw+=R-�x�؅�|�<�f�s�6�ǛO�bG*�oe����۞yl�T�Y�7����TYqr��gdTZ��+l��m<:KW:I�\#�Ō�p�[Щ�f�,�Fx�v���4��La���=DQ{���4��66Ѷ�k�ee�\�k��c!B��D��#�!/zs������3yQm�ξ��n�=6#aJ��WG��ϗ���.r�r���}���~ڍ��Ҷ��tG��q(?� k�2�l6��r�.�y����Xu�'n�2�g���Ӆ�UƝ:���(ۣ$߭uA%��́!dU�����+����Y�����s�E'���{!��EJ����������3���
�`�/�Ń�*�!P1l=꺕�	я��M{a��9.Fu�j���B�c �A�X�b��� �����Ԗ����O�z���{装׮\l��e��3�`��qX:��~�wa�<���`=m�Rʛ��=K,�N�q���vxAv|��N�p+> :��z8q��*Ǟͧ�y�D�T�[�H��=����U����h���s�q�����ݔ�"Q��dv�&�p��S5`��md%r=�1��ᯮ���z[���ϥ�:uV�Ì����z U�l�.�B�p�Fv9�{׷���St���S�����{���Ĕ�x7����U����d�p��ɖl���;�f��P#m�ydoD꼍?y�Ǣo8�l�D0�AkhQ�֝���IΛ��Y�&�^��F�T!3���F5`�}���׮Ю�
�gK�׻LC��,X�\����^��%����TٞNf�(�+*֤�v2��#a��W<�]����g^=U���M���K(�#��.3��LZ���u�����Ց,T�>�4�ڝ,����������Pc�c+�/dv�c�7�i���Μ*���8�_J=&Ȣ�bUŀ�)(��+��&�Kq�D��
�D��0j�)ʅ����f�D����b����i�n/NyǺ���T�[�X��P�,��e�x����(t�{eV+���X�fqm�Z�<Գ�=5��W)�u�R�[+�
�1��e.zN(e���18\���-Og��x�܎Qz���s�uE�yL��0�B��ɦ�2q��}��{;t��au��R���%(ۇ�Y�^�3t�������byE�^TV�B�q��J]����F�
�͠v�z���ոt^SFApT�P�1�V�j��jP�Օ�·�5�I���Y��2�Dߪ:����1J���&&���+y��\Ń�u�v�[ɩ}�p�9�*�{I�uU���/:$X�.�E�`���GZ�Y1��1�#���{�sVfr�ރ$+0;�dЈg�g&kz���<�9NG\[x(-wP��nO���o���wh�<ߞ, �y�L%���\�y0Q�CAH�r��NY ��8/�{�g$h�ˈ�|����t��U3�2p��hYW���5�x�c��>���.Լ�)��̅&���+GL#�u�����XM
��ilg���L�^��g6#K�nH�`x��_4G�=�S�W0��7q���/`�j��9�E���:E�����Ռ�k�'�XRp���T���U��b̹kg�#�Θ:
�ga�!^�w��H{hK^�"'s�`�F�e�N)�Ҵ�{�m��;�ݹ`���'�Ĉ��n"�Ju�D`+cM��Į�g�������0s���:�ǈ2���11�X-X��G�������x�m�Y�U�ѫØ9d�τ���{"ǲ�����(�s\B^&���.��9|�=�8,N�p������=�K�(7����4M���v&ڋ�lh�`�u�:q�ňϕ�]�t�U0�Mv�T�E2�ǧe���L�T�d��#����<���l���O��t�\�(2]���	�YT���׻E�A%��*�����)�G�om�Z�N���D�5�ƫ5��{6�hd�n�X΍5Q�m�m�����xTn���Y~򞡆�T�;^S=��7��Ŏ:OL�SA
ڽ��������q�kMxu�����v��GC֞4}LڗKc �'ٶ�u�yLߜ۹;��Lڌf�<�p��˩n�%���'�f(�<��BQV���(g�^�<t��'[ylߔ�ǫt+�1�|�7k=#�s#���s%���B���S�Ͱ�]>SgW65��fzca�3^_K�k�i��47���8��T�1���|����[��Eף64)jx*�O-�k�U���hg%�Ì*�@�$
H�DX��nb|���yV�b��rw�5��D�5��hͧ��BFK�5uԍª'�Z���e6�N4�����S��$	�/�z���ֵl�5��tA�5�9��c�!�z���Y*�����U,���G8xd=C��3ǥU�h�Jv���6�ḏ�}�z��C��:h�G��}>��&ޘ�!^�O���^m6�DY]�Qۭ��d��g��:�0R�qq�د7�tekP�&�+�����p����`�ǪیQ�_^��Y�R���	DN�@�gX���t��=3C��{1�pMa�-9�dcŸ��m9�joN�t�y�˹/8��c�ˣB��)���sd;{�М�MY{��6��N�8��tNq�S(��ֆO�{�����ν�L��Q�$�E�џ^\�n�YGFnՕ��� n�� W�o���*�
���<Ր���x2��e����lQ�P9����b#�:5l�T�8:������b����o��sk�|V���,���cSǬ5����M�Ξ.lģ鴺�
��7o��\��X��׽��F�*��qQmS#p+�;��N�kX�{G�ۙý3��Bg��f����B���p�P,�q�b}�'ÕR66]=�g��g�`*��m�=����������ڵ����ޚ-L��`*|�I��)��q@����y5�gz3Ÿa�nW�nd+֡��)�:,��-lŗ�*��ĳ�rJ^�j ױHYQT�{6E���5.7[�(s�Օ������Č�U�4L��脣`�8�K�F�ʈ�r�̄W�Ҍ�N�eR�u:%�ru<�H+ԃ�`�Ӯ	��5�@"�[��脣6D��=0�˕�p��^����؛;z���>�y�ci�t�v�������	;Y ?����+��B�*ǈ]9V��Fq
�z$�^�������%a�5�����r8�i�1̆m9�}2w\8<}OQ��ᣩ�o������=_�3���tv@O2���Υ*������f�-	{sUŗ�O��z��H�֜[����8������}����m�cx�Ut}�GK9�"Q�]����C���}p�G���y���%S�u�9M�]{/��7������i���oNK��f���!\1��A�_�د�6�g=X�0���5�W���g�\o��Hb���<d�qs��<�hv��70FM�؝s�S����Fk��G+ps ���f�	Y�.8�X�DO�vxU��_,E:����֚���^VP�6��zJ�P��B}������h%dXteٖl�r�y9q~(���ސ�y]����uX�u}��"�����7�^�Xj��{{b�Xr�
�^H��+¦}2NG���<�Ň�0��%�.��P6dn:qrY��:t׃��&��ۓMIΞ󙃽�b��(C���t�y�m��@�F��d�q^�7E����n��v=^U���lƄ�]d��ӻs�}Βxz���S�gԦ�S��k#��/5;}��U��h�Ž�\}ڹOu�^y�w�X貈�oD�ũ�J&b��]-�7�[��n/h�	�q�Ѽ���1#C6���c2��k��^�ө�CI�"@��eP{R��m��A�OMh�A�'x�
Em܋��cɄV����>�ӥۨLR�᪽P��0\�Y���(�upk�
�'�3����= �غH,�*to3��e�I����P����/{���$�g�<wo�^b!C��g�?k;9�]�������K�^2��}�����'��U�UE�gkz�4X����/T�jY�p�6��9�(��$+��q�ع�5���������s������\Y�_m2�P����I�z��xh>'�����Ѩ[YA�S"D����֬�Fʸ�#zFr�^�3/����u�dk����m�(4Bא���ړb[�<�e���Ҳ��f#U�z!͜�[�ͻ�y6r�����
	��y�YL��OW]�yP����B��|�����`Z�\�y5g�{C�^�O��B��3t6ƌ����7χNzD�`.ˈ�|����<r�|��E�'D+/���G��|���
U1u4����O-�5�l9�	UD#b�B��il`�j:�YGr���f�ݜ-�M2J�����
����W�F^�j`湳E���g��M����Քφ�:�{�ϛ}�kyC4h�i�S舐1�#9��VC;���^}�tm��ߏI������e�0���܅,a¨Y�<�)����-4/�����Ofn��<�ӯ�ٽ��b�٩�9e����d&��6-u6&��L���}�wn��[�tz��,�7�U�5��mY�g_�ۮ�3.5��b�*�s�1^��G׷�+wɮ�q���8�J�V��/;U!�5��x)8�J�&���鍅�gϯG�mX5i{ �t1ig+�b�����{0mf��	��Ә��TPr8l���9�0RVc��|f�����U���$�q�f5�N�R���	���\�,�Ԟ�����~��b�[�O��O�=�^d��N=��7���p�u��=on��.<6�@�{�z�ިyv��5��W>��ݦ�m�ד�>6K�4����7�]���
8�'�,�y�u�0d�Q�$j�Bk�˹evV\\�hW1��B�f¸u7Yk�z	٥	�|d�N�.�����Y��fF�G9pÊ7oFƽQ�\v��mM4��t�=�m�S���Qo��]��N;Α@�w�%��M�|qu��8VY U��p��Fm�Y�RAV'��ܦ�?3E�!��]�K�_w}(V�5��Op೫羃���}|!.Kϝ���e-�r�,�Z0N���T;�"���0C��8��	:}�+�B6ϗ9c
�9ڌG�c4;�1Q�A�Ά
&�W1O0���yS%�1s�묷-l�Ho������z<����;u�d8V4rC�y&��{��{;u�[�)�x��a[���g��xDP2�����x 0��\�a��%�i�.8�� ټ!dԤc�Ŕ���!��������s���3��c�(�J��:/M�F�U��i�h�EA��7�({n�vϥ�Aۙ���t�s����C�K<XgƂ�1��z�^�{�7�e�A3m�y$�=]�.cn�8�V=����v�k�����ݐ�*�u�үs1D�vK
y�Ki����%���#򁙤�<�5��qlj����i7Ln��iI�맔�s�B�&L#ܾ��Q��N�z�`�>~G�۰��˛}�A	Z��8W�YeBY�|��Y}�р/�y�y�6XW[�s�yٚ��V�aݛ�ƷXK Ǫ���w�k^��&%Y�����M���+lιOgؓ�6�N!}��&hlK����+��V��9#l[츞�u��&���Vɲ�1.�P9˅�9��V��I���:��&n��{��܃7�ưe$��s�w��C����)^U�yI"\��:��o>y�}}�|���.e�uJ4?�ݫT�(q�}촇W!2-�pٍK����ME9,^TPN�8r�x^����BmS��nc�&�@�%cNZ�4�y#S���U�(79�1n`��dq6�����(�Q��R�.]�q�)�G�ݴHz��H�������}�nb���r�}#x����H𙳻z�~Ƶ�疸�����*�NZ�D*��mk
�J�0R1
��b�$PYYX�ڴP��R,Uo�AETA�-�-������Yl*"*�J�V,[V*ʅB��Ա�$QA��Q@m�i`a0�EQ^Z�D�ʪ[m��1����X�*V�VV��IQQkTV%j�p���VV��(رH���DV2""V�*,R��Kk+[#e�F�@F,YP�X�QEV�U��EAZ�6�[aUP+PF%j�k
�1T�KmU-*b�E��R���`1Qb�+(�T����-��#*VZe. �"��	R�TQTQ\6f�Pf*ʪ�X�"��(�1-��UDdb..Qa�QR([*�b�6ª�Z��(�DTdPb�V*�F ���,��D���i,Ac*���լ*"(�E��(�[
��X���*	Z # �-FڳF(��TsB��b�(VV`KU�hQ�(**([b(��`(��*��UT��(�EAE�J���b�QQQ�X"
*��*1b�%V�,sja�TEV,X"�E*O���k��x䢮��8AE��*��}���-N��h��gR"�J�]�ɻ��I�H2�\�tR#��Sl�[�{�����U��r|�L��?z��P�v��ۗA2�?Q��{|N�u�J�s,zl��#K2��k̎7��u�=*R�/!�� �N]S^����8�j�?$*:ŝ�����d6#�u�/'��}k#m���M�P����K89�B�����H�겁�3e�;�N��qCF�`sư�z��C��}K�u���O,iѳJ�+��r��N���z�x�H�M(zoS4�;aMԮ�{�y�ʨ�jU-�y�Q�c���OX�'�z�Ӣ�E��q�� %���߿z�\C�F��e"�y>�mK���X�fߛ�uë�yͻ��Ι���]��s�Q=�{N���^�2�ϹoeE�������QcX�:E�bp����c��=x�i�9�˙�V:��|;�'�1J���p*���R+6�U/��^p9\�kg�>���P{6��J��>�Ruq=B}���Mʋ���- �0�w��3\�w8V�Kȶv�Ӫj��W,��,r#)#]aԵ��.'��՘a��g*9ZMm	uyC̜�]ט�G]�ݸ*|��)vfV�g*�9{36�?'Ob͵<������|�aht��=���K�թ맸]^��k������f�>EP;��0��`��pQ`��}P����U�@�Ll��+['nѮ��]��U}�UWٻ��ҽ�N�����Y\ѭ�H�ʻ'D�0K�΃]�U�g��[���X}.GE�j~�fg̾,i>��k��*��w�ݒ͈Vj,��کg����V���r6�
ZӆUmc%GMc��3^�>���)D8������^��O��\�>�����7�vp��0��ܩgh]�c'uȱ�zfu��U
Q.#CS&���kּVn��g�z� ���vzI܋
����#sYL�c7j����D��Hԝ�Gk��<�W�V\Z��Y~ٕo�y�gu	�>�
ŉH��ճ��=��Ń�ӱ�E�'�^��t�����~{�7c�=`5���B��;�`��sH�qfu���Z�Z� ��I�|�+�t�)Uo��BڦF��9��N�X��Xh�gze�aC8A�і6Tu��:�p,\f�EϹĎUH߶]=�Qgqy��Wx[�Rv���l��xc}�}�u0Y��[�v -����g�f��"ߪ�({ņU�-�+ʖVh
Q��n�Y��8��GI��ټ�{���������;�5oOCXG0�C,*�W��]���~-������+���%�������z=�/o�j���ZCR�$B��-�{;�5JU��r�w�A(�0�:�b�uh��:hY���W���­�c�z������0������i��
�%\5w�#�H�����D�r�ZeIK8���2g�B�.�_1#U���)��=�lGK�FĹQ�r��(�Цw����޴�����&�a`��rN���in�e(��nza�+"���72���!������w�V?:g�Y�����f��(�!�Q�n�^���+n��zl�v���na�����il\9G;"Y�C�C5�+idVR��K�H߁v`��GD��JD���s���)Y���͸]�{Ӓ�gY�f�)
��=�]��̼.�dľ���O�W����E"|%�,k��;��i�͔:OP���+7�m��$�w�N��y�M(}K�J��m�O	Tz�Y����R���(]����S��ՙ�0%/].}u��%p���6g�5����	�XyⱖG���7�O+���+N�c�YL7;Lz�vU�a9;�6ۭ9Q/�P0V'D�a{����l5�l<�Rs���L߅n��]��FK��v-SؗI���3�/n�� �]���Qa��^JB�&~kj� ~�ӱ�"�~�W�0�m;�gV^X�;���y��С���)X]���\A�ӀJ,�1��Վ.��)еta���o0�S1s�R��1=w3���|��������U3���������Xej�\k�0k]�'y��ʬX�jЇdƃ�s�"˪=���[/7yޚ�=w,T3��H8C�|s���Aq�eovxH^��6�T,��̶A�Ɛ�Y�=��P��a:.8��މ�dR�pTid��G\��^�o�Ҝv����7Mu1/O\q��W��^M�ꮗ0O����K8�uZ��#(+=�������~�|�f�z��蠾6��ݎ���n��IF�+�DXSj/Kj9��:�S��q��!���N��
���R����GIok�{P��p5,��5����Z:e��H[�[�SnI�����t��������7,�綑f�e��NG(��O(��D�w,���D��׵�7Nq�c1��L��I�#&W��dX�]#�f�{�����%9��'�Xו ڒ�;f����R�e2�t��B��Y݋���2�hD#y0��}l��M��#�(�"6���<�u�.�vFJ�~��G��J��:����b�zb�E��t1k��6#,�w;1wꉨ��t�j)�>o%o�:Iݵ���?�����D�[��Q��VY�3���W���o1
�_KW��pSXu+�ӳ�;]u�*�%,���ձ!qŕ��O�K�3��.dlv捺Iʵ�7g<��nF%2<���4�� �;l,y�!C;���
rȨT(u���|)�>���V��P�w���)3�rC�k.�j�Z������y��6���S$#P����[=u-GVz������W)�;�}�Ѣ+�l^	?�T��@�F^���A�d�T����ɷR�ޘ�^��cb.�`Sqx7�����p�T��>������ld3��Aï�F^�+mj^SVg.��h3�������ngJ��oo�,U�U�{��_u�J�E���N����vꨱ�j6*��إ!^����nc�����g�[��{���3����8۔��Yլ��}ƹ걞�z��)`���1F�[�k����-����}�`�����c-T<���9�(��5�_7~�+bN��b	�'J�=S�r��bE�"u�4�Ă�W6���+X�J�:u�K�f�K���j��o�S=ή���q��OZ���<2��h�j:tW���N�Ѝ\tE�p���E��YP��>Ϳ7l����:�>ٹ�f߱|^m�8���G/>���}��3�!�Z�(�z�f��¾�⻗SS�|���0�v�Ż ��͔�bM0<��4��Y+ـŮz�Mo��;z,�৻i���R���b�:亘�O;F7��it��]NsR,Oӓh����}U�|���3KV�{�d|fcN�A&_�9�ȱ��[�g�3�,k�H�k��O^��٦�K�Ƿ�����_��\�K-F3,�Ҫ* u@�S�'EH��
º|���.�\^Uf�TE�C����ױ]�4�����=�D���P��h�g1.�ZD�oӻfx*��*u&���[݂�ԫ�NU��O�#]���"Yۅ���wbY�����
��ҷ9>�b%�ve�h�Se�\R� �>� ��3��mv�v�s2	I^9��c2b�==�n|ݞ8�zt�B6v��F���C,�z]�,����¶�4��ĩS)��s�o(�m{�pc���-x�w�X�y��:�PJ!��wR��^[�-��D��Cw�z�:�*+��"��|���2w\�q�3��$D�j����dBK:w�.��Z��8�^��p��廃h4J3~��<���U�'oÄ��pK倿���W���G�k���-s���V� y]�3�LlPםb[ʌ�:
6)ɛ��[:�8:��x��j�f���4Cތ��a�����W�K��ٗ��G�7+E�/S�Y=�}t=EG<+;:doWCc+.�4��څ �w%��d�e�W�XBwf�a�3c&����#��Ny���������뽈8zʪ���y���>!h� �f�O�̹�R��x�	�ҫ��V'�.�l�;y�{�7c�=a�X(���V��65x�|>�B��+�H�ΧG�mgsQ�j���WK��`�BڦF���^��7ܸ�fמ	�.v��XVF�z\��u�������~�E����\��O�ʩ�t�08E��yl�mU�<�c:�^5�3��v����6Ӣ�͇6��i=<���Wr-o���G?���3X�w�x��(���1���n�i��T�0�l:����=�VQ*�Z�41HY2T�����gT�r�6wj���#��b{zs���ë,ҙ
!c�R���Ժ�l	r�+�3E?����18�W�y^���Q�O�y��g�Ƽ���@�锣s�$-�����׌�Ɨ5�sxnVts��g���\>R�������nπ��0�d�A�En���A�oA�}�yh�S鐪�=���gltJ�Y*[�+��R!тF:�vޮ)�^��=T�r<JKED}�
�jx:�Qi����j��#8L���+�%�y4R���.�q��xYh6\en���W݄M�z�h�xƜ������{)��sN
dE������2��gt8%���G'?`�Щ)zD`���k���V���L˘o
�kC��Y��trn:uI��QL�ϩgB��m�Yg۽�:������������L�D�����z �Dʞ��0�c]E㊝U���*��fχI�]�V�s�*f�s8��}�A�}+`�n�>l��O�R�2��ю7T.����ϩu�7�Yz�~�o���u�O�~R+ �i�I����	�Xad��|P��aєss�L�]�F.���pj:;so���ˆ�4����Q��E�����(�Zv��T��9Du�V�pzA�u�|GAv��ge�S�۴ld�C [��gqK�Y���t4�>�2V�Ԛʽ�����4��<n���{���&I��஧Uj�Y��ZW'{���7�@o����lb��t�������	U�X�*Y���,�^��r���ءbq�h��|�qN�����^լO4V	�Ka�r��U�WAS��'���E��A�ܮ����m$�n�aD��5){�͖wl+�DZ�QzqǺ��*�����\x,���|��S�9�Ϸ�ۣЧ�x�������y5��)���F�s$-�**"SiAA�g�c*C�������k����.t
�m��586�NI�Qz$N��
�݁�o��.4N���zւ��S��\�RB�� �>����<ӗ�G=�ʛ{)v<o[8;�&6��\�DTWE���v���ԗE~���=W*&��Jo
��OS��3����5}�ͧ#�^�<��s�uE�k�f����Q�1�uګ-�Smqڒ���xB�
��싈]#5�4/z���Ɩ�y��7�z���'9_LՖ��5<_t�1o�hN�Y$p�Mp�F�֙<6�]#���͞�o�A�`,�#våc�r9޳���$5��bG=YqA��#��ߟ�T�1�E@rk	��'{Vx&�&'���z?a�k>��G�J��R�t��C��P�o."_3J"e�9Z*�܍�GE�9�hm�
�`�F>7��\Ǝ��`�a1����\��>HW���^��Z>�i���!�f�7��>���`�$W�+	;|=1@���2����sf�%A�OH����=e)�~�;���wc����g2���"$b"s��o�d3�m\5��wE�r�@�Y��[Uݵ�ʒ8�ɸ�&f�T3�z�;�N��61D�z&	����w��������ǽ�-�H�~^��q��&r�b�-S\.bc���KV9ג/�yJ�N_����&�V|Hħ��]�"@�[�1@<�z-֎�t��v�4���߷�II;�o _=��B���F5���ĳ������'kL�V��<#\ٕ������q�޻��C4H�Qqc�F�'*���
Kv����*�ǎV>/F]��z��47)E�����֢��R�N�`��.�k��^x��غm�\�ä�lA���Q���g��iA��j��6cy؛|v�e�m
#oӢ%�6ëX���ֶ���;(��P�����ڗ��<�{�y�M��,vF��=7I��&��>�u���1P�"��8���(QyH�I�3~
]-�b=x�#�w���陈{3AAX{�vY뾓o�:F�`30��L��2��x�p�,d%�{Lߔ3�,k�H���8̕*2W�˔�H�9�u���rX�K-F	�geL��du��B�y9�U�A�D��욼1x�a.Φ���6Xp��b}�1��4ܸ��.��,닙��KE@���r�V���>�;w��6��i�]��s��U����N�yϸۉ����O��AS�QM�g,u][���ۉ�{fYd-SF��Ժ@4J� ���q��qޮb��)�;{`�cܥ;>�o������K4tL#�y�Yc2�P�vK%Q�_>;�|�WXrP�ƶ_�����{~�����Sx�n�'S�lv�L=垏�1]J+;��[P�\�w�<#�k�kʅ�zI��oXG.���,�飽9t��"���ܻJC&�^���*c��W	)�⽱��A2�ѽ'0)#�m<�g*��!\�(d��/Z�:��M�Z
��ç�s_\��c���*�l�.�j�t���
�ۮ�>A�%�h�Z�u�!�eq����M��6T컦�#'�x�|�9Y��BrB�p3R80ڜ�b��Z�����/\]����k��-��M��Z9m�aӎ�ESrV�R�W�3��Nnqs�o5NsL)_���=�n��⋨t,�\��i@������I�U_
̕�d��7�*���DiwV�A���N�{�C���)gK5��.�t��0�(ʃD��`Ů]�|!�R�:��g6:��oQdڹ2�F��L��`�l��3 9�E�݈k����'p��L�����k��r!!ߒ���6�_h�0f�c]��,�/��\���v�TfV�L��8��n�
;'\7��z�Q���1E��KR:ٱK�>���������ߡ�����T�dF��P����L3�QPڮ.�g_q����d�-��v�ɵ��/p*�=b�w�V��5�N{`Ի��)V��Wc�Y�m���!��7�y���d
9�'-ʉ7���ջ-��d�BΆ��٬�:8@z���\�M�fh�S���:2�q(;+C�wx�
y�q�sd��}˶�b$w,�Kc�oWnf��b���L,J����Lm"��c�历̩�V2h�ӫ�>b7�5�N�3�E�즔���<�{$�"�s�m�eG����������t��X�xq��ګ�\u��V��2���.	�ˑy�\\}�b΂�{�F�F�p-ձ��][n�{�E2�c�Fr�7����-���x���ᶌ�'*ɤ
��r�aq:ܪ�v�YWC�˵g`�3\���t鍊�u���XV�E7o���T[u٘B��
ӥ�{��B!�ֺpR��)弓�R<�sF��]��.�<�Δi�����T�,��6!Y*'t�Ƭ�5$JE{f4*h�u]�te��T�S���ّ���T=�CK�p��o{G8�ܱ�r����1�ݛ�|�fi۲ou�)���e&Ͳ��\	���_=���(�k0��4f�c�S{�p5��XwrM7�Z�ɫs�����*�����/w��K���������5�Q~���6�9(��k��d���0��fr��&Q�3gu7�kl$6�)��n�䝶N,��W.^�Л��dd�>ۧ{sn
Q��9-r�,��gi�f �;8r�/j$�Gb�7$���Ok+{<�d��M�kv��M���M�[H�Er�wK�p%[-sâv�m͐�Yq��2��`�A��9N�-5���]��*�AH��Q�Q-���DDc�R
�V��Z0D��-�T-�QQ���X������X�T0��`�Eb"�2�DrѮqEA\bkE�R��"�TE�UUR"#�(�0Q`�1r�D��+ŌUEG4��lR҈�E�**
#H����QQ����`�J21�Źj�`��E����L%H�G4���PQAX��,V*�+5F*���D��e�X�)Q�,Re*�b��*(��UQPEQ�b\�S��*�.Z�U\���,V��H�,Ra�D1lQE�b*�QH�X�(�-Eb�R�J��*�.Z�ְ�DY�Ab,DDJ��Ƞ��QAEF(�AAG6����UTV*�E��c,
�"
���DPURڱLU"0UQE�U�&����riǤ��u�2�,TC�/
�`
�.�h���9���4�o] *��8���z1-�"��4�q]�^Fн���UZ0��}l��?
�gv�O�e�c%�Mr6fk\�h�H	L8�m�\B�?p�p�L��|c�L�X�[$�|5P:���9mp�&J�k3ʦ9�� F�]��n���*�>�����.��F+�0��2���_K�܊�e7j��1�7ZN�#{hOu_m��D��i$P]����6(w�����,A�/�
ŉT��[:.mn��8�������+�������{�7c�=~k
/���7'6Y0���%A�������;�X�m-���pc'���Q��8q�j��]a݌�{\l5�,V�p���3xƥZ+�/yX�8���:�r�H�]!�B�8�	�(�UH�˧���,���}��-y��_v�]�OQ��/��\�����6�)w$஖�qF��TY��#�����j����Gv����Z0-9���Ņ5Jc �ue`u4�`��Uz娃X�,��ظ93�˚OZ�+�N���	{Ӄ���ë,�
d(���Q�1(��י�*����t����~ⵣ�@`]K��[��X���3�K9�s+`����҅^���YY�tʼ���[c�i��h�\��+˞P0h��L�Q_vl�vF�+��'��kM��E�>]�p�Yx��&��a�Ѩ��┌ޮ�h�fG��xxW��k����/�:U�ҍ�|�`,]65�;���Qn�锣pH���M5�gX�4��l<P��/���%��O�6�����N�Fd2J3n�B�T_^����άk6;/Ywӣ���Xyl�U��[�Q������W�|��b�^�|5�A�ґQ�nS^]R�3��,;�%%��>�^�x:�'�gJ/:xK��f���!\15��h�*{WZ�%���}ծ��e>㱒X�$i.���E(�tX��/T�/)Z|�����e�"Z�]֭�Ǌ�q X+�d1.��²�!��!+"�2�Պ�E��Gd3����g�V�z�rQ{݊"��,}���t. ?����[��mF@x
�-єsr��08e�WK=@�==5U��7�[9q`��'a�7�l(��"��AkhQƴ퇀q�u�ڷ�J�r���F��J��J�&��&�B����b�F87���_��3с�Ӧ��3�;˩�r)�j�?OP~�1��y"3u!�����Q�d>/<�]������6��{ �'�̦t �PĆ�t6sl�U{^2�Wn�1�̀��doG�~�|s�rM���� B6I%�n��'�ښۼ���NXZ'jIN�w>@�7KP��_������7�y�u�>�q+���u�=�^�'t��������h��۬0��~�:"k�(�#a�V�L�:)M86�,����W��Ʋ�#�׵�*L9�;O;����1���.լmx肘�usO��pT�3��n	��[����$���H]]Jz���z�m�(��Fj�)Y��.�u�c��e���檳`�x��W�pL��R�Y��1��P4��9m���K�8Գ��@eE(�D"5����u���}�=er��Λ���|�"��/pm2��o����O(��D����\��z%���b��\5��{b�+����P��OC�U?_�k�f�O���	��6�L@��F���m�J�W�٠��<D$xv���*����G�g&t�����C��}p#w-.W��+1x���+��x(-wP��dq3���eҥ�*�XM�T8z�ip!&�J��n_�fwB��|5׼kK�� �;<ˈ�B��QT��o�ְ���S�V)�^��7�^�u@�1�.cn9�%��iA�!���\!����}��^�uI�/}YE���0���ʍ�,�m\�*)Π�`�LsRB'����x�_*U){�~4�c/�i��A!���4��/��4Gs�N?rm���r�(ʽ�UC��+�ɐ!د6,�D0�*�k��
�;̆W"����S{��u%{��ӗ��G�� u-)�i��\e^")T򰓫~E���:��D�26��4Y�
M�{ʝf"q�ǡ���x�Z;Et�R�oL�w�w�͌�ۛ��8�����~+!��j���FhFm�"8˪�N��ʋ�q�avzM�ډ"'k����Z����F����2��m�t9Wr0}ϊ�Uo�}C̱��'ݸ�+ʪ��
����Lpt��f�b��z`�������v���V}s�`5��4')E����o��b���W��8vn��겁gcYXD�yGfv��¥Anx�7Tr���5~���+bE]�a�9�2�u���]�8��źi�Ղ���0e oا����-C�gz]6ڧ����Wuc���;��!q�y�����vT)��44���p�2�(��Y���P�dc��ݳ�.u�6���z��|=\��2������4�k��Ab��ȿ����=��]���t:�5{�g����6l��bp�o-�Sn䰌2��e��2V̎�G;�"�{���u��c�n��*� �w���K��Q`��6��Wg�34J(��\���c�i��G'!\��j1��n�0��f'%�$�IVGک�d��T+��\I�K&%�ˍ��u�z.a�k��7u�eG���8������0r�.��3� �CU\��⺇|6뚛8W65��c��p7.!aK�z3��P��<E�Lw7&�(7	OB2lE+P�]]t(�S�����W
u�'<�
�CO�#]~u-Gd�g{V�m���6=�P�m�G��d�=T�������	�/;9@�.)t�h�Qd�\��^;D��n5S�挽Q�23"��,S�s�I,����*���%ݒ��ًMc5A�U�ښ�Y��pe�8F�ʵ�S��N���~T̡�Y⩗���諷#���*z��=#v]��XI��q���z��w����g��":�i��9��^�d��a�����51���#�Y6}�2̮a}.*��;��e�EI%BN���*os�Z���tLJ�D�Mec�jcb���a��أ`lPrga�����3��&;7a�Ʈ$�y<UtN��{�7a�ӽ�`�a��X��ޓָ3&���{]�y^��r�4Ϥ
ʤ���b���P�ul�V�25T�̍ok�����$l����Z�B���j���Ȑ�_aLX۬���y��*X��8�*����J��������m�&'^�mQXw�J��%FU��Z%�t嗗'wj���hP����4�Ʊ=�pA�ϲC�
)�~t�6���V�I�SӓVB���й���������,�fS��cܼL�m;�K窺��o����(�2�xl�{��ڊ���Osx[T2��[��7ݎ��>��ˋ�cG�u�� �p1ベ�Pi&#m��U@���*��]��bQތ�Ӷ�F��)�8�ue`u4�M�+G�Z�8�+�G��z�mV�n��ǟ�v8���v!/zs���ë,�S!D z!(��ģ���=�r����l;x
����(�?_�fG��)�0w�X�$�_��@"�n�e(ڗW�u��W6��K�"e�ʄlK��p�͖}՛H�-V�K�Qe�x�-٢a�+v�q��u]h�[ޔV�Q�\;�!P���b���,����W��M��zM�J�b����ኺǪ�� /�k:Lm�U��	u<s���u���U�*����4���؀�z�<��p��bT����p��S��-ߞ����V�j�����w멜�z2ҋ�m�~�{^篓|�i��]�6�#���C������f�!+"̸�uH����U�{	��+��Ω)l��q{ڨd2�r��S;�Oq�U��E�;6����)�ٯ=�\��pj�/t| :�v(v��Bi�B�ÝE���"v�����n1+t����.�r{�d�A8q��w�n�r�n�u!A����U�kj�;yw~�15��H������A�ʰ��mF@aW�FQͤ�0U[�vglA�:��[Xh��B7�u+bhl�`��vJ6^Dhj����-a���av��Tdou3�mKf���De^ݳc e�k|X��]�'y���{)���
�n���Uk�Nʅ��*��x�M5':x9�;�8*ʽ�`���j5̋�����3H�t�5�����'N*���������U���ƞ��iH�.2ࠧK$�Gt�ei�Q]��Ιۣ�s�'K�.��UPc�y���vn ��KTb�Y�t��&��'��%g�i�v�������U�UJ!���@��Fj�)�l��`+�DXSj/N�vUsN�ޫY�굲�yv#�od@(���+����j�O,�9�t�Գ��@f��Qhߙ&��nn�L��Q�H��H݉����Dv)e��,���r9E��;:'T�k��*�<��)3xn��K#�����g�Y��.�"�C��r�^�3t������P~��]���7/������16P�ШM*�����jA�����OM��̣ںY�r�_]v	�l*�ն��0l��5̭��7}�r,��Cn�[Re�1���ؐ�:(v��[�ȪF�+����P��R�`)�5p��_T��c��˱Ξ����>����kXsOd|�/^TV�B�Ic�wG�_��e~W����=-�Y�z��oSts+ZXRTUF�͖)H��x(-wP�i�uN���gj���67W������}��A����y�Y���~�T�j�`�9dT::�ˈ�B��Q*�#�2�y��������ɝ��Oo�$��*���k��A�iA��#�*��J�d`|�-�lk�x���e7���銤t���f��r����ȱ������dc�M�,�����l-�7j9bΦT��C-Nk�f�g�]I��}g2)~_qy��!\3�ˣnUk�8B�^���K�i"Ǿ^[�6)	�	cK�6Gf�
�r�z�;;�,D�bDh�Fe��4{!�#"�w>u��>�޷��s,zl��<,�׮�3���k/�ϵ�E��#�^�ճy��U��J�?9�.�+��a��	�Qe_N�}���>쥂�x�c��^�������7w���+�`��j�/�uG-�M/u�;�+bE�j�����؛r{kLq�����z�XV-G�mq��+2;�3w�(��J�c�t�����`��y��;3�NA�#<(I����{�y1&L�C��(N�Vwl�;WGQ���n��}o8>����� ��ܣ��|,=��l7=��${�r�NW&�J���$X"��J./�H�a�.�mS��yLH���Lv{���~�8�w����;'�:��lH�P�,�2�f��fԺ[�O�b��W}e%r0�L��)v��ޖ�q~h^o���a#�'����{�+���W��2b��o{W�ot(]��M�:bQ�5���f�۹,`Q,�3,�Ҫ*���B���4�(�c	���ȋY�R���V:��r�9��α��w �r�6��=�%��r�����a+��pu�9$ip��nL�G62�;*w�[�*�:/�=
�q��! �-���G{|.쉳,y��#n7#D)���%��Y��@�>|$���}� *I�sk�Yh�9	�z�U��V��z�v�c2�z��ƸӇ}͝��ho8�,Y�N������r{65�92O;5�![f6�n4�˙+�Z����*ē�/�K��J{(��H#Y����?I[���1bki�*�:��[)E'��-�.��뽰�d�5�L�ގi��ۙ�����c*����s1#�'7G��]�����?�?0�J��-���RŚ���ͫ7/�f�N\�>��
=�:p���/����*�0t/C���,�qH(�����e)�sV6=��]��C�َ_p����U �B��C
��5����=[��Z�[k�b? AtÌ�����y���~+",������6�p����*����k<��c�������SY�g�g�*��Y��6�}祜:�g>��A�BM�Q��JS��dd��(|6t�\�=��{�7c nx�V�Q{�)�'u��1�9AFO3Kj����OR�Y�N���о�s��ϙj���:�F�
��C͊q��ܼiot�n\1F/��O��cyO%c5+�t�鮠���/��u��g��㺠�Q~y�%Ҏ�4�����m���x�O>���m�3���=^ 8tw*���2��=���f���$�l	aGWlog6-Ɲ���4�)�9�ë)�K;²�T.Z�89j�� ]nۚ���z�����K��D�#��<1#U���2GP�{�m"�bT�I��/7���w\�X��(gJ#/%y:Q���2��/_��M
��B�Ǘ��8�k$��"�f�u����/.�<xl���sZ���u�32J/���tWV�M�O�o5v)�v�b�T-��R|U����n��wd���ȇ�Q��nҊ�y���A�p�0�0F�^��虱���q���r����Y�E���ڄ�hj�"0V*��ΰ�jKHyWC��5�dD�]c�,��H#��,����+&qs�>q�>z6�b�o�3*���4=����k��|��Y����iU%��NU�	�������p�ç�v+����;�"�s�G�a�5��M=u*�)�����Ӊ+�ƻ�_�8;ݨ��k��j�R�A`���"5�ݙC^~�N��_n���z\�5�T���Y��#/h��Yo3qc]S�'�mIˑ��n�� p{��̹�>�0<$���6�u�R7XxO��(�ֵ��}����F�Yrv-�� ����U��Y��]"e�J�ݞ�zj=�,#q;�������픲]D�@^��G&�t�gm�-DGA�\*ڈ��(���S+��Q�4Q��l�����ǖ/B�ۻ��O=�WI^�vPɔ%�7W��;z�F�z������W�#gF��P�^^�z>־��{!�6�<HO��(�4hsh�GR�������q��n	��P�� c)V�D�p�\��佽��jzC��Q�z��a�,���u��|}�ͳnQj~�A;�6Zfj����+R��r�s��\=�ۼ@�鹛�_n��.դJ�\4�^�[}݋������g.J�bN����#jg;����I��Qꂯ�30��Ź�w�^�{ƈ8�:�F����'��NZrV<Aۻv��<��NX��3n���}O2����5d��P����(�Tw[vɽs����[��)%��S�q�)�z���,�=b��q�h�����v+"6w�2����]���877��k�r��[;�1�J�E�#�$qjb,3*;z#�����Yѳ�+�&��.�\�m�*�\0�GH��A�H�1�C&0G\��3���5�����[ō)�+ ڴ0(*c��HZ�ĺ���7ۮ��{䖘3����ݺ�ϲ��^���nE�f�H4M�Ղי���Τ�tt���b��aB��\��N&�ȟ��Ӷ��meh|��U�F��^
�J�b%�j��;/���r|�Wdth���G���j�s��2I�7���u��B��ݏEb_�Ft�luB����}����s6�ˬ��]�5s9�����ĜR����܅kY��#�J]�O�?��1�a��q�4���c�!嗳w&�"ξjŁM����2�_|C�.��O-���w3F1(�ۊ����qsY*Q�r��Y f���O?s5g��T��⛊��};���Ž�������\;�����RC5���9�ᛚ���ra��q�>g��u}9vֵ��8f�u�49�;�3{��;��^c��A1X�E�TPQVUDV������@QPdc,X�P-�Ŋ��,Qb� ��*�(� "EX*�b (����E����DV�b��ED1B���EF[F1dQ���-*ADTQH(�Ȫ
�b��űV(�*�T`� �T�a��bDŒ�IUDX)0ʑX�`���(����b��e`�D�ȥJ�"��U�DTPU2Q"�PQp��E�(� �XKiF$X	hT"++QDH��"1V
Ŵ�8�UE�AdX�("�1KTb�AckJFڶ�+�`��J�F*Z�F+ik[eci(��Qb*5����kK�7!����l�\x��/�&���a��ኵ>�>K'w[�s�s���J{�tbV|eB74y��C���o��ն�Y����J+l@��/�����b����gv�f�m,�Zf����z'm�
{���U�Vp߇@@_>�:Lm�F
�s�W]E��g���W��,V�4�r������7n:��;�0R��,K�L��"�y�4�ߞ�R��aqx���dG��	��nd����e��O9�v�n �[��r��<�+*"�J��T�"�7ػ��b�mU:�i�ݘ���#^�.ͳ��W�	 � ewY+��k�s <	Y+��M����C��K���z��|,FkEԵpχaOP!e��	\l{	�"+>�L���ɀ�Y�k�����'�s �9�a��Y�,��۴o eB�1���>�T�/�v��]7qI�/�g#��z���K��4�ܚ����>�Df�|-�2OP�pWS�U8��R��Y�6R�+x�J��t��g+a����<6��&�`����X�W�^	�~#� N��^9!�7�#�w���~jhg%Oa)���<uǕ]`����We-�r��U�W@�0~�I�v���8��<��k'5X��Y�iZIķ8��fc�Q������g<�������{ס��<Z��ӏ������f&������!�}@�c;���zU�SzKj�uaL��}�%R����K*\�s���Q�}-�?{�*��;:�[��pO�t�ce<����Od`֩�E��^b"�ڋӀ8�Tw�+���Զ�+z&�7O���*�4-ˈ��YqyL�R4�ymq�B^��5,��5������gF�k���qH�x���H[]P���1C/;i�h_m2�P���dU�9r��g&mv�<�MW�WB�]�$
�Uf�}~Ȏ�����߅���p�ő��{:�
�"Zt���#T-yPzۨPI,���DWy4"���.��Ac]u�71��xd���a\�ɳ��#�-���m:��,U:GrD��r	V�5���'Eoff�U�E��f��qͱ��5UK�NY�nmG�t8��|��ǶZ�����z��;ɱ~��`��ږ��hׂtP�+t'�J�\1���p����cv/[�cy,������G�n_��w���xf�>�8fk�)1G�4���Z�9tnPb��ubͳ÷���vΞ.�5�5�>�^�������<'�s"���%U�**����6�g<S-�d��Ć��uӁ�]E��$J��[m�S6Yh���Mn��wc�Lq`әEPZ@4�{k�����0��[��㇚����3PS.�Ԃ}�ϟ^�]%��M�a)0��NFe+9ENk
ޜ�����h�K:��x=��bS�}¦0�}���Ϻ-�\P�=P�-�"v��<V�hy�,��4�K���ܽ�������wT����a;U�o��s,g���k���mz�> �S��ವ�1'Ъ�`��tߡ�g֔��\#�u���Y�MSF��}ѡ9J,}:_d��Z'M?,b�|�Q�8t�,�o,���YVP7��J�-9�m�`XƩ��jؑWy���Chg��{=�c��Il��A�;>�r,:����t��e�]C=E��^F�<�{�U��t�����Z�O
,s�;i=S^R�",M��q�P��f�}LڗKa�16��e��r_��*=�\�U�VT�M�������N6<1+n����d^BQ�QoH�VM���Ujֵ
�ҏ����kg��E��rX���o�Ixd�͎&��������~����V�����,��4���
���6s�+���>���ˈ@ߔ�g�H�v�edq2��2#�p.�L<o�%��g�nL��3`#B�����r�f�V�B}��'M=�ۡ]+�ñ
�Mr��j�o�^=I]�S�w\&��o�3h7�t���H粀>���=��ɝ��s[�l=���惫��W:�m���M�`�d�s��%z�!;�Fk姶�F�f�����ϫO�=�s�f���9��?�h��g�m:`࠽���Fo9��F�(��'N�ˈF�7#D9��kt�,�+T٫�#p����D���NE%)<����
��n�ecA�P�e��1�C\��K4tL#��p��\�Y�jf/c��;kE�u�4x�����ck�q�g�;�+�U�W�N������3���s)�tǏ��o��[s
470p�.�Y�*"�$Q�8b"��N�^�j��tm ]��z��c��nv�fXJDJT4�q����wM��u�g҆�2̮a}.R�۳}&����V��Ϸx?�*O��j��1@k�bF�"H��S�Ddv��a��أ`lP�rr�zz��-\��2�0����kf�Η\�5������n4�5�5�N��nX�_a�>��~�1��0�┟������W�x��K��9È�mS#x��N���WǛ��M�0���X��=��Ps8w�pVH����{�o*�B�hÕlu���66���Q�����ګ�7��ܞ����..Q�yDϫ��h\qH�ގz2�6��#��u�h�#s:O��� �2V��R���eJ�/��cUaVǝN�X8c����]�� L��.}����w�����n��9pu���]���ʕڵ�z��������kkx����{��)����l;-�M����Wn���  }e-6jz�G�҅Oc=�K;х�Ӫ�#�MR�Í�VVy��=���]1�sw�VK���S��h���:���{]��rE�B^��čVYf��
!�	F۸��'��m��?����v��_DP���U^V�n���M�\��`k̂���Yp.S��� Xgv7$H[s��Y�=}�ϧ՛Hإ�٬���*$I:�GM�:�JQ�M՚&��U�C+6��W�B��{!�9���v�fiLQ˳{-��n�J���[�:�r^
D:0N
N��-�­��x:��O�<=��f�[T�$R������(Zf��Hwg��a��)�J>����F����J%�OW�}o��V�˩�xD�Mw�!�K�����*�n`����~�wa�+*"(B��NVugY()�ʞ�z�b�㐱�#�)zݛ�,����D�)���U�L\��^��!о�¢�7�΋[ѝ9�U�éx9jჇ��X��/ހN6=������6���Y�+��M"�侻2��3�����=��]��Y,x]:Ѵ�����N�B�X3K�v��G�h�ޖw������j|؟�"k!d�k(�Ϗ�80�V��b7��M�w�çS��2����JQp߮�q@\xx�����|7�Ny�}Z�����Ӷ��K���"Y��x![g����^��Z��2�b3��<�_m�[xK��U�!��{)�u�y~�/V���ԇ�ɏ��8+�֪�1W,)�{|������e����	�y��X�����+𞵎Y~4�\F�v�ݢ�����ŝI,(a�7Z���Р�x�+����A�肻���R����:��&�Ӭb�z�)Tb�X�)�X�DO-���y#��O��6Yݵ�����^�\�GL�Gq������N����K�i��JP��T�{C��hF��~���p��¬7"�Ί�҅Pl)N�%������
o�N)�G_���b��+�]@b�^��e��{�����e�w	j����,�Y�~T�Q˖|A��l��'�߉�|�~��hV���W=;�]<].�D�<U��'�k��t[u
���؀Q+��P5�ʂ�';���U����M�0QO�zٰ�y���NG\Xoz���AQT��H�w+}�z�y�;�թ0m ���I:�Q=�Z��Ç��7gl���1<���F�`���nԋ6^K�M�U�IZr�Ht�裮*+]��df��N��S�H����Č�sW<��Jfit���ڦ�����,�Sd�q�Ӌ����.�/��k�k��M�dG�YY���.���j�g9dT:9�����iDm��8K��S���G)�U�k'b�E�H�90�Ex^0���B|D��p��
��Ѩ��7��X���垒x6Ѯ��u)GT�82��?	��"��a+\<���:��CE���].-FN�:|F{�z0pC5���6ԮkóV|φ�2xJ���>�����pOgE���ie�[/D��X/#��U�˺,�^��q��`�l�B9z�>'v嚷Kc���,�m<��IF����>�Y0s,ez)����U0��0޵�獵Ҷ�
�˗[:L�ݓ�gu�0���<iA��-��GYo����{�t�����X�b�1E��I�U�sps�vwLX�g(_U���pll�ә6ԇ�5Mt�y:{���6�
8�1��q�=5E�%�ۜ�lX�`�u���(��E�P��"ζ�� �J�#6�7�u0�K���[�'�jT��r�ڈ�%M)Tؑ �B�(���)�����f���ʞ�֕X�)S)Z�0`2��Z�\:�R�Wm�U�f�%��_6��.��h�Ɖ����F��\l�D+L�2͍���Vh�5�%�E#B�/h'.r�t�軤��D�G�����nb����BU��q�lg
K6��h�ƞ�
�>�>Ͱݳ�0;�f������3jD#�L��w���i��G��L^�Q�A��q��Qz���,k����jmܖ0(�Z��v�*����f�*��uGI��(�� �Yr���Vm�a]>Sg������V;�����.�ꀩ�NC/6���|�u^��z%�P:>[�"�Flj�����+��B���Oj �� l*�&��9�	���T�xc����sVa��鐮%���g(|�I�,�G&qL/d�坓�>�� ��Y�ck�q�]g>��8�-��`��`?K�����k{����/#x�p�=R��f��f��f}M�ƭ��d��k�S��IZ�טc�Fb�j��Ǯnv�����n�J�ه�8w��K7*"��H��=q��v�h(|a�i*�K�U����ֳ�.C��s3�f�	L8ȋLl7uX�J>��h�݂��h^��}��VT&�sц[��nMq�;ڨ���H��xc|���kα6ۍ�;WmN�3l��R��'����&6��L&����Nj�,q�3sN?{�)���H�sp��9��=j�G��bSpv-��Ӽ/;Kf��Kku�u�f[�1�@)���ĈX��AZ�pU������l���J@��ˉ`�Ş����1��v,Q�rgl��f�M;gK�9�8k���~{�7csǍ�E+Ƹ����n��V(��)���5x����;o�J~=N�h�>F�<|K�ӡ4h�Q��~8�?h��{�n��c[\m�Qb��Sng��
�	ꮠ�>2����@�ez�-z��KV4+.�S���{s�-�m�Wxm�w'�Ϩ������L��d���:]P�M
��o��H�=��{W�=���,�F�i�]iMR�Í�VVSL��:j�8��x��IL9�hrE��U[�
�A[�/��9�bF�4Y�2Be�l��jr�]<��͵�_�Eh��3���9~\*�-`�ԟ,�M�rN��أvYzfo)��<�$�+F
�Oi�*U���Y��d\9G�e�M䢩j�kb��'{���K�`C$�6��5}��+a�]e�
��~�<xM�+��o&#���
�S氤$��k�/=]M�wK�����KIIp���#�U����ܓ0 �x�]�����r��yk"/���� ��m�rV{#�C�a���X&[��n�	Lk��i��p�<�:�'k������\��kH珳?:�{4�M�H�p�m�ްs�om��ޛZrK�����g. `��u��ka��M�.���DZ�T�t��)�T�v�F�)
��{�zS��ђX�4���R�K��}J`�#��uՂ���0i���H�.{���*���u�{��<VTD3p�����p�t]ŝ�})���?7B��Avt?��"�.. Mи�^J`�y<�g_;{U9���J1v�W�&x�WQ�}^ap���,9pu-\0p�7����^���P�$>��J�Z9Z8�n��s?c�b��ӶPo�����L��۴p��C@���J2/^r�W5F�ou<�z*�"{\z3Ω�1��#9��3j�����KX|��w#HBQ�Wep�̴+�,�X�О��P��
"��L�F�kk��Ѧ��D&�xo�c��e�)����i�w�1�<�n��A�҉/�]r�k���Jp�0<uǰ+��aŞ#M��z��&�3��=��\�_�]�NJ�mCqe>���S��S�:l����%\�Q��YV:^����#�P��(��u4��xթq�Yq~�e�p�`T��ϯ>�̷�=H���9��6�A
t&��י��i�g�9s6�3ts�͖��{�u����+k�D��ЇkK��P���W]3�W�n�b���dz���W(��u³w0�����ê)!&`�ge����^���$6���gp��ۙ�ֱ�~_^u���n]H�� rś�R0�j���y}�ī:�ϸY��e6�f\�n�	ƛ0����*���H�Bj�Tl����0�[��\�V�/��/L_7Q����48Q���p�� ��=�ю�'�����Ґ}�hg�[�g}0���J��
\�f[��nI�w�#��:�Ƭ��ci��b�ڨ��[n���1�f��6ku("2�kL̧:���5�'O�`M��g{YBe#J�x������&gf0��=��Uyz������a�3�a(�aۆ�1v�SU�_N�ux�^�Nn��75pv^�jK6�0vj��&9�a6�{3wRS��@� ^<��N���]Q�Xݩ�k�T��}�AF�-=�/�������
��t&-9vD��{N��STu΍����l���Wu���qU�Ÿ����#�XF=�-2����X�BxNvg`�xMmj/�ެ�47iY��R��w�nA�b���
�`;WL�E�����ƆJN�2�)i��; 6[ܕ(�|��\[��C2
s�缁I��6��l�#\�;2��or\��R�>#x���)���W��o���o�z�y�B �o��rr�z������2�>OЇ�"�;�_���g�c���G���'��G�̌�o/z9���j6�wʶ�����&BAԥb�6���g7�gAt�Ҷ�"9L���v+�x'�N�t�8 |���|sGn-�t����6#���wG��Շ���N<TH�.C��x�Yu)��8֭����Rv{���Iᮻ#ً�"�Gu�^�̱�%<u+�.��O�W+@��_�}�yVu
�Ͷ|zVk�79d�wWֲ��>��Oyj��V��6^��G��e��c�Y �q�3��n��H�� ��s&�}�A��y���k/������7��cķU����L�^����%]��i��U5ת��>���k�lL�g�y���W�g��vJ����7����5��e\��1�;g�F����0����٩���fh�k���g�>���s}��K�
��}n`M��A��}�5��rT���{}[[8�w�7b�v�{��>yu�-��ʎ��D�<�W�~��P|�~LvvM��d�Z7v�D�j�y�i���z��xw/Rx�/"Ϻ�٪].I�9o�Ğ��nc�}�	�X0�X;n� (�����Ւ�S�*�"8[>Q����i9Z�v�[�o��-E��c�{!1��{��!�OcB��S�6Wu�z}z�s5�BK�w�e��v��}E��pp���-��T��b���u�8ŃmT+%UVE���E�ԪŊ�j"X"��(T�bE�"VVA`*1AE�
���X��Qej�" ��c���Q�
�U0���"�Ҋ���ň�`"�Eb�UAE���F
��*"�����"*��ň(�AU��`��bF(Ŋ��
�X(*�b�VacX�¥QAVDDE�E-�"ȱ�`�Q@PR(��-E+X��� ��VV(����I���Q���V# �ڈ(,X��b�$ATa
� �(,Qb*�0�\�;Ѳ�Z ����W4!����1t�;84w����khuE:�J�S�3C*�V�r�+�к�w�Tb6�q��z����n�n���'f�i|_�K�l�$+�Ϝn��WDW�K/vYe}��D���/*.3]>����	���:���)����'�* �V��5���v��B�̤4%�2U�������]���R��&ӭ]e�w��[!8�y�*�^]��[�!"���j�e�T�*����iP��b!��8&8��޶m��ɳ��u�v$.�\4Ӽ��e|ߟ&�l���G7܊x*̷ �5.#+6o���.��#U�8)�"�С��D@���Hٸ�޾���\O�=l7wt���i����S�ot���4��R�yyzި�S3��Gu#��qb�A�2�;��Z�wM�`w1�J�DR�r����#Z�Pb�j�*�t�J��ۗϖ�+x����Fr"��8C�C^�#b�5�٩�2xJ������q�u����R��d�e�kAg�ذ�:h>˺7�FA�C���#o����J�g�t�[q��Ʋc%F��.�x��H��H�m߉��~0�C�c*���q��L�zŨ^c�9�e���FS�_F;tO����CIk.z���b���rSn8���ѐu�AY��[�XSDu�a�	;[u;n��KM�dO�����V(L�o�O9����2����R0y���V���v޼��V�iW�Z;ʴ-����=|��%Tb�]�c�F��ڳ�2t�A�d�t�^ܤ���w����U���]0�Ĳ¿
���k�sg/oyҮb��8vn��_M��n�e�ɼ�j��1�k��a��f*&Ӣ�MfcJ�)�8(�]����6�+�"���HΔ\X�E�R���CF���β;zͽ����4��7甏v}y�Jv���k�<���q�qF��[��ا�;�6m�)�mɺ}�m
�E�U��O�l�p���N>tͨ�h��:��\c{��j��w�=.jUf7o�u�5Ž�Qgz�'��cX�=m�jmܖ�_B�v��3�L��mI���I�S���W;�U�AhWO����́�O����4���=���j,���>�����J��8��JK��@B���(���<��Ny��*DgG�|g�*�Wi>��k6���XU)Gd�gnC;��݋�>��W	��<���ig�G�w������L�ҵ︤�=�5�i�ێg��eoYg��4��o^�*�o�V���ʄ"�*5��_p�/�ȱ��V1V4��T��\Iv����	sU���d59�4�e� h2;���Y@���y/���r������,��T�6�Ky�{�c�z�-�"��T���eU���W1�	Cju�/gY��j*�w�.�n��N�uR�<�U��X�O��33S�X��J�OvU��3-l�QUL�`��A�^.�|���D��/,���p�ߙRv?m���#��ݷ{�;*��Vg*��RN�����Пt�,+�&޺��XY�,��WyY�W�	"q��/ޞ��OR�}N߆���8%��^s ���A�������:�=��ƲQ��=�t�[.�����X9�^rg��7BTq�-�YC6t��=��v��R0�V'~y�"V�b����P�fɥ֬Io���_���6b�f�J>�ʤ��b�;%�
��%lxӂl�rla؇��������y��6�(�V��)pt9w+����ei\||(���m�sĩͤrn�us��Ui�t�=�p�=��϶�����ܞ����7�9Hŏ,�w��s��*��o�{0 ��1��(��t*{�bYތ-Ɲ�tQ2�,�l:��z��x�y��=��tb�6�(����b��,�U[�������寧������VDy����
�k]Ӻ�9v��.ۏ��!���k�"��hy&�wg�k��טv.2_׀�h(Բ4���y+�<�·�uw����]��-L^k-�T`����>��og��oe��zL�Xr��gN����G�T$l�Mr��N?{��b-�z�� ~S=���i��S�ؗ*"��#/�(����,�9�A��,n�!�R�Nڲ��H�zxWPz�q˥J�z��Џ-xy��i�!b�Mi��Wٰ����ya�'��IF�&�}��B+���TЫ���2���=��	ʼ���vvn�ͣetXU��/)Sq��G��@U��i1�­��x:쳑!އ����}YK�{/_�c���['�3��Lu���¾�T?*��0-�-�\D���/�%u(�Z�k�qGN�ʍ�YӲ�9�U2�A�ؿ��וXI�c}�^�h�<�o��>�r������u|������g2A| ��wL�bmWxGZ�q���y�F��u_#�������м���Q{Ce|7�G7�^9�׼�9�K������E{�z�Q�����3f��de^ݣc e�V��sȌ3��n�+���=���xB����9j�+݁��$�l�f���,:����u������o������%�n��m�D��5��[��W��rI2zk&��{�,���ׁ�W0�t��$j���ib
�F���� �b�W0��l.s=�����$'s�͗g����`Ժ�xv�xut2�t+E{��X�9�yZx�RW�Z+��J�V� ��;�E���
"�{��B��A�x�X�K�M�W,����+�LN���ż�u�=�>"V, dqt9M����S��Oq��6���֙���[�Ce�x(U�c�+z'*p����P�B�DH���Odf�O��6Yݓ��h�Ml"!>�O6�YԸW�T�0_�~�vsN�/�9x��)e��2�(�r�����]|_<��q����/��<�k 3JmE���Q`9�����UtEb�^��,���"{w)wڞ���i.7�����k�5sig�g��B�p�4�\��5[�d�r�����R
v^ĥj��+�ܳB���}<D�:z���,kʀh[u
���*<*{Y�P����m#��ny<'8�hDi���	�]�l۹�g�qa���E�PTBB�]6��B�s�������� �v��̇gb0�]��G6�t#U�9�rȯ쬩P�[���:}�����v��!�w'�O��e�~X������h��a1����Zb���{��z��A�)5G9,a�{Z:J�7u4rQ&�:k��qX�J�wh!�Q����g������q�LX>���9�D��">�S������i��	���C��)��~�w�bD3�B}����z�@�λ��<�Ow��>�ʁ�HV��:{�a�׸�o����U�"�	E�Ȝ�)�Bv;y�k�%��g���ӛxC�C^�P�S�5�٫>g�c���Om�S�c�3�C���[������ld3�a����e��q�av�^�"'j���~���E�ϳ�x�s����ܣ�ѬH��ڷi[񄯇2�}��ޏ9����^RbtR�}N��wEs[��ѵ��T���ڳ�2tӃ~8S�"�nRF�n��Nm�*�����WB5x�A���a�4������ó���겁��-���Zs&�`Xz���:/�t+����+n�̚����:�'���6�+��P��ϨJ�\<f>|�υ�bL�G]����7��aK��9��3ݎ���_����kO�:�R��J�q�.�ł��)ޅ�A��7ug��X���=��ض3�X�f�vθur�yͻ�����˱S��sp^+r�?qV��ѹyGz��63�,bx��Nn�Sn䱊%������@g�n&�_��a8P���BJ�w�ff\�q���`Ɋ��eۚiaԭ�6���}ݫ
��K�~�����)u|��f�	�$����B*/w�t�����h<]������-��b�v O���FWV�4(�q9aa��P�:�x:��jY�l�wͣz�x���?;l�@ꁂ���B*k(*
��M����X�wwpM��sʦ𺵂�,��T�B�uǠC9��U��f��=q�2����KS�X)�,��=Z���N��ˍ�G$�a�:��E �_B��8��SVa��钊�2��u����'�3an�HU��R�?J�'��R����D��[�n;~S�\_�V;<�5��]�2n�����C�0G����Y�uD����p�쉘g��EB=�h�����u�f�ë��~I{O��s3C\�h�RҘq���A�E�K%\�C�zIi�=���-gd�*7z�ʈ��;�=��92熺x�p �d��(28VOsr�-�\���\ٳK�mg���d�﹅���v�xe^c�}|�3�F\�J.=������a��9�"��#���d~{V�aG�������n�eG��e:]s�p�kwf�U1&����jn!bc9���[9��<X$�}�b��9�`��Λ�G�+3:��^=H��l!~ j��*$:��hh{�D��
d,�3���k����J���:��.�)\��*@>�pE��kuj!���2�.�k��WwC�5���^SI�VH�ռ��W����{c����P\<�r!;�[����JA��9�x��bG�5Q��-1N�u̇#�q��W�C	���
j��n07����*���6�霬�5�"����e��!��[9*�ּY�1��۱#�R7���2�;�<�}�]��ܞ�>��͇9H�F]C�f��z��F��:K
�I4�<�_�9� V�U�Oz�����+��R�`�1F���a5�5��͍�m�S\{+(�W-D�,�(����"�!/zZ01[�Ǔ2�M�q�m��Η���J���()���:�g�T�B6%ʈ�r���EU�c����ʽ.u܁^?=k�ɚ}մ�~�$�Y�C,���J6�u�ߥ�ȸr�fm3�gi�;�8�4�������\i��Q��d�fݚ&��Ti�Ei�_
�����C��n�|LS�u]j����d#^U��.T�`���@@]<֒��Q�\,*Q�[���o7/��K���c��\�XοT�r���!�w�ئo�� s�4�.<�f�A������^S��,8d�x.\l��9�s~�gz�Wl�E��<�%��z��e���MF$oV��v������ۑ�[5���,~Dc�o�(<qt�tR�VI�Y�L��z�{�b�z|�]��M�Q�ٯSz7V�ۈ���bI�|�`&ٴ�n!9@j�"���}�Ҭ�S�����n�s���xLӋt2N��|�r���Բ�N�ip������w�O�S����ԆQ��/Y�Ńz7�Vx��d��+"à�^]7�b3\.���|8{
u�������.(��<�J�#'}�Ey�GZv��T��3fĲ/}{v����o	�ǲ�t�|�tV,���
�eg���h{��F:t��<`�[�rj�`r��vC���|��]����S������ZŊ2=s��<�]�����!u����u	�V!�]��v��S�įMN��b���Ӄjt�M�*�M�.v�0�N÷:uU�����h���+���dQi�W.R��S�Ȯ����)n"��#��[�)�֩��ֵW������5��f�c��^�=�j���XP�-C.S.��8Izs¯�X�X��I�N��%�bV�j��5�6����(��2Bؚ����(b�^�"�'CKܬ[˧��x�܎Qz���tN��k�j�G����yr��n�7�늸�x=g4tN�;�;r�hF CN�u]���s�(-��0'XHׯ_��]/��ٻ?k�k��$�\�	G�ek���%fu��~�u�`��Q��O�/�}���c�����P�c��JNu�����qM��&�P	Й������gpNa�x�/:|��z��}\D�<U���w071�P�,��31p������!��B�dЈg�g&kz���y����G\7�B�.�$8�Q������E.�ĥ����.��b�zb�G���y׸�s^�¬��5Z����Q�N\�\�E�S=��?O,���,��Q����g�����V>,	�q�/�ϸYJ��q�U�²hS�ilg����m�`w1�K�E/�+	$�^���zubi��ڵ��;L3w
� �T~P1�(�נ�6���ׇf�g�\�<7��w7h�Ț�+�����q{�|I� E���`��v-����e��#�uD������)r<�R��[�mwPW�(�li�bDm�q�q�2�W���~����!Ó��}ޔ�W�W��3�J���Վ~s$^�`w�����(�p!c��ȘI��Z3���/������:E8��f�ʾ�(͖���.�uG-�`/U_Z�Uۯ+W�;4�(n�.^�i�����IԢ(��v��}X�v+p m�,Wd�;*j����:᧬)�[C�3n��l�l��Ũ"J���	^3�F"2���L<=�A��(|��Μ�O�)}'�������i�h�C6_+�����ݓ���n��fRU���p��bΨ�E��0c��t�>�):Uq�\BW��M�������ni�X�M����W/�Sl��]���l����7>1K)WA�e�=���}F����$TP�Z�Xzn��*V}KUyN�z���+���W�9U�Kw	�.�E�z!	�a����d�`�p����
'`��6�;m7�M�Ӵʜ)�N��丽���K۵�uQ쥧黺ි__�!h4P*O���) �%�ɜ��c���OH��|/z]�
�r���wj�Ig
HV`��_]5��ר	m�%8d�P{t/��J��ݾdX�� ��[f]>Q^�C�U�����@�!"}@LV��3V����W'&����Ҏ<�V˧/��+Y�څ�zB����-l�ݐF�`[�:[�vv^UX��Й#����8T�b�-4G��� ���We ���t�!(Ke�&Ɖ��د2�6�K]�oc�G(�����]�>�AO]�݋�PB�5�d�1IvE���6s���>���5�}�ÿ�̋;/^)�݅���6N	��{���tFm��AWX���6S���@��1JI��\��	���B�t-}g�]9\��m�ڍ�e�)��K��.6�u^���kGqDݎ�K>��L���dp�Ԁz�cɺy�7�A3���;48���\����p��B�ޔe��ޭ쵅�x�s�r���"�Y�yV�_g1cU}���c�,��n`��q�-(r��m�u�-���-!z��cØ��V=s���{��4$��[Yע�s�+b`���8'k<����袲-������p�)�[�f�4�dѼ|��`�:5Xv�0`S;9�٘\�C�k���i�Qѧ��[���]�ШaƁc�����Õ�Sg-Ӥ��7GsMl�o�[�M��C<����O�m))޺���G�ۚev 4��K�E^���/)j$�Y��ƕ-�pbb�^ОC�va+"�7����!n����=h���͟Z��gH6�af�(1h��8�L,�邂���v5F\\���W��Ӱ#%��Bd��5�8�,�˥B̶���CrWPip��+�\!Fy�]�ɔ����kq��|��_%��e��Oa��";�eY�k����=���|]ne�h�+O$z��#�6��N9��rj��/��W"�� ���l�c�o���z$�H��ˣ��*�t��p�8eZ|�k��e�iR��>9O�+���U�2N�	�2�����rDz�-�}'0R���e�d���N�����+��j��ڮ���]k+i��O7�F_b�O%k&�f)˩=�J��a>$�I�N��,E��E+TQb�,Ae�Qb��R()T�#��HUb�*�1DE�l���`撠���UU��+�Ea�UE�T`"�*"1��*�(�(�(��X�"�,���b�,T�*��J�TF#Ub�#����Q��AŨ)UE"���*�"��2� �dUQDV(#�XDV
��Z�U ��V�A-�1L4Q����V��2*�sI���W��<��޳٠�-0U�0�j�����k����v�*p����"2�K�e�z����zi6�k]݁��Ծ����5Po�l6��;n��{b/Ӯ�9Ћ�6�{u�-�'dN�hj�޶�VE!u))y�S=��0i��Ŏ�OT�RB����������=5,ʼY{|����ci��T9Y�z�7l�W,��Rq�o�q�	�Dy=����ef��Db0�jF��oi�P�(��O"�����[7�6�Kt�@����y3��ޢ��e�2^�du��S�'��l%R�M�����5��56��2x�j�7z�����9Q�t�`�,�z�T;<E��)덈E���Z�
��i�+<��.:��hg%�Ì!V*�B��I���Mʋ��MY�/�J��LU(�^Kko�r��O�w��#%��l��������aE�EN��<��Y���/���,�rr�K��/dSS�S�����ʰjx�����g��Z�xC�2��m����j�g�2FyW5�~Z.���TӇ��3,k�h�%0�E�Pt�.�Y�z�'����3�Q���$??��4q9�{��ܭ�/H��+�	{������"SqK4S��;}X&�V���ݬm��w���M]p�:2u���WY�D'h��ۗl��Vv����G�;�]E�^�	�=L�mp���oM�h�F�Q��Eu���^�fd6���/y��s�.C���gZ�0h%0�"-����2Q�a�:���o{8u��xz�h���/����ʾX�`�[�?u�`!q�<B�y���>;�r箭�c�b�ʌ�:
6+�L��~�F�Tq�[ڲ���I��k��4�γ���f����˂���݌jx��x�I�ۦS���[�0��+���>~=JMv�nE��/��SrC��b#}U��حҢ8j����`ok���(�Od��霬�9#w��1q	�VX�Mmr��}����yU#{.��(����5Wxm�w'�>���׌��z�D�-n��ޘa�>�,�g�F8ds�+`*
��k��g�q�m]{[�]�ۦ�At�l.��G�.b�«+<�i��+(�p�A�\,�Uz��V"
ޑ~�%�LUB�<'k_VH7�Ys��X��A�P�C�.��^����~���+"�:���G�O��PXNn����H+�A�
}7�I��whp�@�L���!m]uB6%�ȱQ�"A[}C��d�q
�\nW6��w-Ϋ3�& ���v�����'ʍ^w��/�����-^_��]���̆{������ch��T�
�o+ڔ�.X�����3��N���Nb��Y�Ro��Ľ����� KR�4��'aة������hcP���Y��Wޓ ���l�u�0�J=�vh��$뀊�&��.�45d(Z���=y5�|�������s�D���:�id^R��;��@@�䴜m�D������DX���y`����q���Ξ���S<�*�;��=��S6;���9q�\q)0��v��G�o��(�e�.�\l��)�sc���*���u�l�ȇ{�?m➋;��-����^���:��O�X�Q1C��+���.�f��u�� *��&��^�Ȼ�]��a%�9CVU�����<P��n�����gz�B7�u
/bN�4���j�v�dP0Xw�d�e�F�PD���6֝���IΗ^h�de^ݣŮ'z=�����o�uʐ�i�����qӈ[���y�Ӧ�O4�6����;�a���龍�r�e�y��rͰ]�`did
q�d_�
"��L�E,�,��H��h��wU�7Bd�"��6%���4�߂�,�^��D�\����G���z_T�ۻx27��CË�T}�d�j��P��W%�ۣ��ގ`0$W3@�o�v�JK���6�=�����}np�+��t��!�u0��oDh�=g���m�kd��g��vM�IK�9ݤ��aM���ƀ�|Th�b��,���_f���y�)�Qc��#M�螸��)(��N]�:1Kq6Q�h+���U��]ǻ:�^����KvY��v��",)��{�9LHY�X��P�,����ե�Lq��*�j��2_��85	z��y��@f��Qh�B#x2BؿU����*[�f�{w�6��}Ӥ�6��Ư�����Q~���tN��k�f��O��Th����Y���9����\�����
㽮Y�{�����&Ӯ+#=�O(��*�m�(;j-u����WM\�\֝:VC�dS0@ՓB!͜�E�[�̀�y��u�87���Q��\J�B�I�|1i��,�O�3��U"Y� �Q�p^lؘG6�t#U�5~ѥ���T���d�>8C"Fns3��O����g��.p98���ra�sL[�\�����j��ru�Kl�t�GhJ�!�B���ZZ>�/����"��p�����m�Y*�v�j���\0h$e�j��9�E��&�1�z�]K+zv��:5��]3�E��J��z��zm;�lD&Q��F.�����L�E������F�[���P��Q�?�Y��pT��Q`��x��*��!y���5nt��4{9�B7}gnP˝�����{�ma-�t�t	�ꇘ餒�ζL�za3r�rn�ɻ�E�Ҽ�~�ȥ���~�F^�z��u�3������Z=����m_o&=����^��+rd�밬d�ܳ��k!d��g��<t���p:�^�+.J����>���WOv�#ҡE7 f�&s�Q�2c��Z���0v}�L��mvg��c;6w�R#Gg��~C�i�8˖{���v֢��R�N�`��.�:���[�����Q���B��M��3Q���篊�47 ?7ԗN����O,i���:l-��7�+�(��:Qq�v�J{J9�7S��݃�ʨ�b���mS�Z����0i��Ŏ�OTҕAbv����2Hу:���o�=g	���FR,ד�fԺ[5��m�l�w�͇6�N��Q5�̎�א�<��qYɜ\�lb�6�L��閌Q�d^BQB��7�����/X�=m�f�ņ���;kA��OK={�PF8�C2�ߩU:��Q���
���6s�+��W����V$��O�ҝ/���Hhf�E�]3�"Yۅ0�8�=�
z�re^��\�we�L��TdE
�,NK�]�CóH��<g�ɮ��C�	�K�}��3,�v���y:�.R[e�m��'�lC.ܴ:��F
,����p��9�[�^�@��1|;}�E7�z��.[)q�=�wcs��i�6��mޙ������N���(�gr�9֎�V)�U�%�!p�@�'ԑ��sF�gk�*!����ňs����W���q�]V��u+�6�Qf��6j�*F�J�KUqI(�{��W��i�ێ���,�Y�.˗���(�1p�*���%���e��;ޗvK%Q�82;"f�-��c�{&#w��s_��i��\NF���}��P8�Í�:k��K7*"n4����Ԩl8婝D�-�;���v��ñ���^�陭r"F���ϊ'}�Yv�`�����z�^pךǨzɳ�5�y󖫄N߇3v��1���ܔI��t��ʹ�>�S�fs���*�{q�F�6)ɜ8na�Q���;�:]��IǪ��Wkqv�G��M#k��6W�pu��	6��Vtw��\ىG�,Ρ�<��<:�;|��ʁ2���P�,�p��L�U6s!��)�Qb�=�:�N�.�Hfj���nz��휍����b}�'�R66]=�g��3��*��a�w'�*�B���*��^�{�m���陹�m=��ʂ[�[�,o�H�낔���V
f�&�!�Tt1��ͯ)�tK�����I�K�}7�	��=�~�����y�U~U��-:��ԍ^׽b��Q7��!��PDm�	��}��uB���v�{��<?r��Ͷ���)��+`*�S��bYހ�aͻ�^�8o9[��jಸ{��e����:�g�ՔJ���(
�FB*��`�٪���x<�s�Ի*��p5{ɔZ�
!~锣�SL�T�B6�Q�Qy(�s&y:f�{K��7��qY���rkx�ytߵ�;��y�E8d*�.㖩Wc�=g����h�M�X�R��X=��yۻ�+tϦ�i��[4�yE����vh���M� _����hN�@�O��,���<f8~�(�`�g{�C4�id^z�7a؞��/��p��s��6��a�;���F�#f#M�AP��٭�^���j��T1.C�b]�d�����T�^�~��$�O�v�0��z�R�IxXB�eˍ�^�;.o���*���j#�M��&��>�J�ΚZ}�_�v�P�	<!�]f�\)��v|��S�\b�*���K�b�[+�d�7 ��i%tA��U�L\��+"ã(��S8��9j�Uh,��mեh�r�6^��6<�˭��������ה�B���ȕ�gl�3w/�B�O:��a�2���'�W��cp8�/t�M��)ُ�r���5����[�8��/Ss��,�f�-�Xi"Nn��8e0�j�+>t�{�7���8n�v4-�vJ6^DkUK��l5�l0��O9�+7=4�λ���#�rp��s<X�Q�����`ِ78��[��F:tןO+ojMkTw���o%`�-�i�.{{R�5T��υ�o�+ն�qu�n�������R�҃�����v�"��},�
���8���^k�>O�q���gG=*�v�N0�N�i�����'(�j�����K�&�4V	�Ka���m]�{�M�R�E��D���I�v:�q���<N���9��[M�b��ܪn�C�=��q�w�SAnU`<mC��Rˀ����ʸi���V�u��<Ð����Bt�Գ�&�3�Sj-�Do9�Ŋ������[KdƊ��3qإ����t��t��]Wߟ`
�����+F��֝t�{��ox�J�Ax�2�FD.�����Lا��Js�\/k�/�^Ta�DՄ	����{8�x�`B�z�<���ˀ巓r"�o[6�<�9�r:�#}TU���D�tGf�垠�I�z��,WΈ��񓹊��'�l{]J����[fN�݉�J�Fv�Lo
&�����ޑ�2��Av�`N!���~ޣ���,:�ņ�Fvva���XuV�G���r��mq�ڗywԭDj�/����d�T���m����(�ߟ�K����6,p��#�򜆌ۓё'X�vL�+rHP��*m;��W�҈�r�V�3��'��hY__+G�@��j�=��Xo��,��5�m�GjUQ�D�|���5�:��\��2C����oz[v�`u�342�Sz�I{ڢ1���f��CmO5�٩�g�fϰc��֞�X�6p�s"�~_W�	#9���gb�WM>˺6���I�ą��/�����X���v�Õz�;��ݹgƑ:Ĉ��n"�Ju�J�̱��o���{]���;�c��.}ʪ�A^����nc���\D0wyX�Ƴ��-m�䲼�,�:IJyU�s�˸�5`��Ǩ�+��
~0X��sSC*�{�a��*`�P1병�8栵�4k��=�ߕ�"��ULҬg݈lS����U(Q��}A^��z���̬���S����X3ܼτ�t0�mS�Z���y�M��,vF��/��r�-���l�5�f�Ӯ�v]ݭ�|��X����GxT����6'G*�DS��bv��/r��꿭������V�����-ug"gQ�N�L	)�嫙���!�F�
b0vC���{�&�gns\����7~Gō�K��kEn�l���2<Rׂ��Qp�X�E��}L�R�lf�>Ͱ�u�y�S7�6�N���Ίus3�D�k�u1��%d������T��u�B��7�����,k��m:�1�u��f��jo�OD��`2������徵��w��WG���s����=޸�����O�{�A9sR��"YڹU��f�
z�pL���s���ј���涰��[݂�O+��T1� ��tE�����%�����ݍ�X�*P�h�'��+s���%�bG|V��W�T�ؕvV��)%zMF|���������u|w��3�k���f#�<pX�xA�4���zg�]�,�F`�Gd)��|.�q{l��e����������{O�g�935�s��H�`����e����;�{
���o��*f"�RH�P�k/���{\�^��O�.�)���>�����c~�²�N�OWeK,���#�M��P�Y�s�qW�~o4m.�� ��
�]����??{�.���s��v,񚽢��F�4eG[�£��Qӂ����`�B;�j���Q︙L'�= ��N�㫣X�bz7��cK�ᷭ&�������7��Ԟ����]�wD$��;˲��__!T���Y�7��)7j�'>\1X�]aؕ):r4B�L�f�Xysj�|�}1�@���כ�w���4;���(Щx�:�(��'����vT���qq��q9�ϻ���G��}ݟzTݹ&����R]ci�R	u�y�h۽����I15�Y^��;�u%�Ԏ�V�\�ċ�����0��a�79������]Z@�+x<G�v����Ku��nij��l�k� "�XhvX׸��6��#%Ӷ���nF��a�_�i-Ǜ�#����"�Q*��%*�۬%���u��������3���vT��=˂�p��S�ʠY߻O
<E����eH�w`OKD��V��C�W>�4M���&?��oD���/�o�}���|pE>��B����i=�~0��hc{��{���騋 : w[�]�sxgY}��j���S�U����|����K��T����ٵײ�TlF퍹4���� �@���}���,��4c����F�5}n��<�f\���$(*������{�f�|<�B�!{�:H.�+�oj8Y��_r@"��w&p�I�D\�p\�X���w�`��u���[z���g.XDݭ������4oug.;���<��xC��^�;��,�1إ眏�+�;�Ū����S�}���̉[q�V�M�:��~!�=WY�
�̦i/27+��5z�������2�D��� r��}��ʽt��g�%���/�����{�JW58�������U-Sn�N	{7��y������v����9�񗷮z�L��}w�n-j���#=D��ו��Xp���h�G)R�橌l^�9h+�T�51�g`�����f��@��i����%'��m[x�t{f[�7{�M<����C�����rʆ>X��_�3	P2�WFm�	k����[q=�3�a��9�V' x�F�q����T�9ʹ]�	�SqQUc80��Rw�f�����$r��bgs�RV�V7\�۸h����Z�L.��u^�Ÿ���rW`'m�'RVZcG0��"�N�:VK#66p5��CP�)!�g��ՕnomY9Vgd�.J���V�2�hm=��X��&s�M����崏5o>���++�^������#+e��ȣ��']�y۷��6�i�t�Na<���x(MWmVH� rlk$Vt�Ɣ�h�D��s��O8hX�w���K�7��� �T�>�+$��9r�N3��V�)�D�D��p�7�C_r}�ML��gby�o�7*9�PPP�%d���2(�����I�Z�*�0D���)0�X�UEF ��T���T`(��%*�UX�X,R�jQ+F�ҖZ�mU+-h*�[-�0�Ш�hV�eKl��ULb�P2 �ͪ�Ah±Z�QmR�eB���X[VR�V��J�
�[m��j�G8��Qm�QJ�U�A�H�E��TL�bQ�ʕ��[!Y*Zږ�ւ�V֔m���(Q�ڭ���Y�* �kQ,��μ�U����gWI-)^��c��}�`�~t�i�21�Lz��i��g�����ϥ�7.9}Oo�;I���Y����~����J3�M�����pm�����A�����V�����2�e����J�.�u)��,>�=^o)����	�=����X��ޛ1p3f�� V+nk]p��S�&��f�u�#Tp���WK��c��V�27���7���W�S��7�����0Z�پ�/X�IB�!W�ŉ�(�UH�˧���,��-�m�Wxa�Hy�!2���3�W&�N��6��b���d��⑌<�f�*�2������P��m^�vKX��n��Q�R0�:j�����h�Q��I��WY�g�?��W���ڄ��q�4;����t�؞ޜ	�:��2B�e(���=�9P�߯�^<+Yo�e���hܶ��n�n�F�>X0.���'{]��#�2d+���nL<���詧۝�);�[O77�����᷋��N��֫f�O(��d�g���4�Th�N��Rp���qh�JZ0T���!P�Ob��(�dK8k�C5�[K"�R�����h >~;�P���qi��r�xO{xe����$�4�g(����&{����k��i3�%Qe�:r�sMz����Xį�?	�^I&�����{�*2ۙ��)�:����o
KQ��^׸�&q�#�2���w�l[x����l3����;�%G�E)�3<E�|rE�A\tl�E��8��3\�+�0S��7�I4	�=��ͼZ�Z���ђk4����-���'eˍ��6\��޲�٧��44ىٗ��G�s���ྕ�c�������O�R�2��ю7 Vx]��^�;1&��A[��)�f+����xl��Y�Ze�i�����<mF@yℬ�te��S8j�B8�B�Yn�Ӓ���:�\5YVv���� y�T����Zv��':m��Y�Y3Ll������d[}v����]+��^��Z��<��3=����{&��ڐ��#��輵��i�*"n��۶p�p��������
"��L�F��㕵��oDv�(d�E�C���=��W�hi���H�y�~"r��R0vN�����RW��y�D"�Lx`�vyL�/�ڵ���D����)D��k��'qKq6Q�����L5��U�\���O�%-��KޑE��y�����q��
��ܪ�t:��M��+	��u�;�~�G̺�[}W��$x^��F$p�R9"ѫk��1������g5�͜p9����3�Қkj���W�ٗ�s~�C�KB]�q���,K�*�6sy��s�kp;���Ɛ}}2v:3A�ϼ}�m��w]73b��G"{�c����[tz�߃����ǆ�/zZ�u�5�^�u���
�$W"�cԟ��_�ȝVw9�Q�Q{��(_m3i���r�C��5ܳ�B�6-w+)���S\�6��Am�SW��싈]���s</���[J�.��n:�/+w�����^��s4U�aS(��B�@דB!͜��.�޶m��ɲ�V�/z���s�҇\0��U��w�Loφ_ԩxc���Ma6��ŵVx&|߲U��:�i��o_�9��W,�,�
~��@��i7�����N�V9���\�����ԻY}S��*h��4��R���F�Y4(>f��u-GV
�t�,V�.7��Ow,;���EN6���P�A#/`�Uh9�E����%����>�{x�X�p�;�'rtc)l�G_���8w*w����@��LY��=Ќ�r1�v��x�W���<�H�!~.MƳz�w¡��^�����T�S�]{��{��d�,�#<'x���b4�os�JȪl�F���
��*�Z���ɝ�VJ��?n,��龛��c~1ڭ�PM��"�;�nk�������i*�� ��<����&�����Y���~/=�o9�	v�Ӄ��\���*;��Xt;|�T1�弩cދ�c~���|j��
�����-`|E�;đX#vT�ҍ��v�[��]�7�n���q�:j�+ۏQbWe,�`��U#��겁�f�pOb�ܘ�U�R|� �Uސ�yꦺw�'�rycH���^9_R�����'��&+�w"f�	T��P�,�,��m"��K�f�6T���{�����x��di=�����M����kM�9��+��B=�C��
/)i>�l)t�3X�f�n���3�r�6����;�*0'�<�,��I�t���3튙#�eq�s�q�!(�[�f�3�,bx��꾌��y'�w�\�bF����aM����Q�2��*��du�*9��EH��	�G@�w0��B�I#��l��'sz���c��i9s�L�g4�P왁f�S�/�b����Ga���N�w��6q@��]���r��B���HV��"��Z��H�v�TC4-s�g��i����^���7�E���N���/;9@���J���q�
{��;U+�jØ�Z[�[�Vu�Q��5U�)�vڥe�@�4N�z�Z�>�=��Yoї~�n����^K�ÔOi�蛋;f=�
V��ĥsw4���vi}�y,9;/�����_;�?\����
�[.YEv�ޫ����J�k\&u�x����^�;��K%��:��ƥ���7�xۈ��S�I,�� ԣ[�*��e��wd�U�6\h����c"��}h�!d?UK;�9Q�h���t�935�}��P8�q�ۨ:Fإ4��J7|2�M���N�A�`z��QI�x��2��Gh]텑��c���5ȉ��A�]�^u��p$C�=�������,�둊�L>φ�2� ~r�p���7�7���~>�>]f�9�ś�{�`�:�H����jcb�gX��"��P9�NL��s�Q�N[d�|�ע�˅�S����*�`G�a��7Ɲ�x�I��z,U��;�~1p3fv�j��VL��1��c��&��j�6F(B�����a�:q-�dny]a݆�t����}	�o>檳i�Ǘ�X�8�����3��$WH`и�/�}�'ܪ�����c�Y��<�}�׷K+oq7��ٴ�����<W'��l9�F/�OO$�"�]ȫ7�v�s�t��г�ںU/T����2}uT�t)�Sp6YXM3���%\5tb��-r�/����nﺈL@��ދ�i��X<��hz�]����ʎ��y�mA�o%D�N:��u�Ճ+:ӵ:���+W"�䈂8n�'�-M��2>���N������ ����m�вH^���@@WS�5���<-6֘9ZI�Sr���5п{'�B��825_�Yf��
!~锣�ĳ�S�ؗ*#sj�F,W�a�(J��sz���mΕB�)��M�w��� ��B�L��D���m^T���.X���N�x׌�i�.��xz�e����N�Fg��Q�FI�/���;���Z�>&$]��æ9x�בʶd*Զ	�[��E���yV�ȹR�{j�͌���_.%k��M����6"���g&����cf��/zpL�.��R�}�d�E?������ծ��Ke:�h�cx����=�%�(@��2FS�����~9-�T�0�nru���,}+b�]�XV�D
�BVE�ˎ;VR"E�d#`�gsۛ��v���E]ۆ&�{�^ٸP,���!����O*����!\s�G7*��a_`�+:�{h'7�d]C(�9��(^�_��"^�	-Y��:bZ�Vk��u��B��;X�%n9�]c�:2T1�-�`��.!�-�4ߝ`���B�q>9hصS�V]�2ED��_�t����giL�wag���z'�/n�<mi<k�v��N�.f�.ݾb�V;��v�:���>�i����͒^�_;�F:O}�z^�<5��e�R<��3:������C&�Υ��nC=�����H��W�3�s���m8�i{��P�8R��	�6�ы*F���5�ZN��=���+uV���l���*����
���S�)����*A'?N:�w3\$1Uy[g���: �7�����9HŁ3`��PN�Jqz^�<r��C�hɺ�����>��06��,xfs����`����Ӯĥ
K�ƥ�}�J���gw�B���Ga�"�(�Uq��K͔�lMdk�mE���¥lR5
�e����8y�SO��Õ�����5oi��r9F�s��':-��Dn�"/�rb#�CzZ�Gp8^��j��F��=�.��n���O��R�w���Vn��%r;��R�I�4.�]@5ܪK+"DN�K�5�ע�ق��c�](�[.�׷����4XW!\[z(+ח ڂz#]:Gs�%���J�Ӈ
.�X��fd�՗�W�kowS��I�����r"��N�w\$����mh��	Z�<<�>�3�=@{�2s���h�˷���cZ8�tˌ3ǯ3T��ǂ��6p�fn�\9��x��&j�drK6_{�ԣ��|p[���E�Ymލ,�a�F����=҄he��n9q{�׶!{q�>o��묥4���i�#����KT���}M߃�5�{@��{x�(*9���ЅDР��팺���8&D���݈\v&�Z�[��7�`��8fk�)�h�B# �0q�(��B�dk赃n�p�k��1�����ćn�z��+���:���#�7���s�p�iT�FP���u��T[�#�1j�B9^���פ,X;�A!���},��[<�;�k-���K���q��nM���*����6%�\#����V�="}j�yi��iE�9�V�Wsٹ��z����w���ʾ�Or�b�B0�,�ٱT�P4P1v�oٍ]�L�׏
��<z��8ԆC���-d���� ��H��N�ߔ�{c��f{�DJJ:�g���ЯW8����K���W3��g[T�u,�pW�4�n(mі���}��bO�j_�L�#hG�È�P�$3�r�F�J�����6�vΑ���=\d��^�d}����<���!���;b��"�q�s��c!(�{C���l!�b�N�:�R��pG�Uh�����K�tQ�)��B�e��a���dx-%��X��dZ_���E��Eϓ�X��$7V۫~�3['�#r+#�	t�ު��0�a��]��)h��|k���2fL�r0�J�;��9��gi��]$ڽxp+�F'
��ٵ7PP����G�TU���M�瓄"�JO�U����݃,U�^4��;*ut�F�K�'�C�A9s	�%�%*\-Ŭ�K U~M���/���3r�ݝ#c�G�*2�posz��?>Y9�R-� �}�JQ�$H���C9OI��k}։6=�������^����L<�τ��D���3�����ql1:��\��N��2�FS��X����Y�q�� ԣ^�ue��Y���gu��-F�-j�U�oVK7G`�F���ɹy"�:�l������B�E�n���ƹq�.�FMr/R��D�*nW_�ߏ+��ʭKع��MKu!]���s�g��G$7uA�6�����qt_?r�#߾��.6��اB�~���Տ�1�yqرX5*�7r�a��i�2�[fuY�C޲_��諾�B���YO5��]�R�ؚ�C6�w�2�;u��Un`�&Q�qE��b��2��U!ڄ�Z9���Ҧߕ�5��^��.ËC�o�j��/�E�φC���ۜv)sgy����x;���(�S�L�sB��k�@�z ��q�s�W2�dd��T��v��t��Ք�^s�������p+͠�����X7�p��=ҏUD����͈�Яv&s�����۞�Z�n� �X�'{)=}y��B�T�aT�5S���F�s�u]�Ga*�\�ռ��_co�Sy��(�a�;Jg������4b����&LѷS�.��[��-���X�m�ϳ�7��R�/�	u�VǺ��M��&M�`���o������s��#�ް�����Cl�]	l�y�t��`�[�r�D7�>/�-u��Y��k�Oz�tC��-L��G̨i!
���V�a��!�\Tּ9�9��tj��N�iT��f��R�ܽ��vE���x�>��i�5�$by��\�"m����y�5��v[䐼��*CrN�g�C�����?��c��o�1�tbi��W<&�ޫ��\���1�KFP{8�Ύ�b���p̶��1���.nx�m9�2� HIQ���j�"+,��wgq��o���\+^���=�hG����2j�M��C6�Z�W�҇�u�>�)���@�2foQ�4u���;6O%a�n�ۛ���ݥ#ǜ)���Hy�������x%�.,�a���-���'�o�xI�.�|��u�.*I���BG/��e^~I��I�og$���mZ��kt;�@CV��0���:fb33h��;)�Y���+R�5�Gi=�eir��[.ܕ-F�:��D�SL���'o;���h)[������}S�uQ��35v�_����]=�[W$��q��Y�u{wX�͟Zm&�	o}M���'f�X�y��I-�TEOz�j�7��S�r�oL5}d>f
�D������sH�;ZU*�B�K��A���7:�VI�}��i�﷑,f_Flx���˔$}���&�^)�e=�vI�9���cntM��P����ϬQ�.�vU�	d�����gQA����W�Uc�[��s�OE�	��i<Ѣ��J�Pշ���Py7�j݉�n�6޷�رl���Ѻ��7�{��\u����L�$�ݴkML����߯ͅY�X�G�>��ɤ�u�6�dُ4@�=
�rfr�L����9g)�����Ff3��,�5�S��R��<ffC��Xc�W�X0dc��j�b1�71��j_�m.��+����;��G�A��J7�w�[���wV�;Ǽ��eܕ.�l7}�E�"��XW�oT5FA�ي�syc�Sz�L�gw���6}ekݘ�#�W��ȥ�]���r�{��Ln�1�l��}ۥ�fn�f�����Ŏ�};(��3�{�A��=V�6Q����ͦ�/o���%�<&Gp�������[��]����s���7n��ڷ�l�StW�rS��rxU|e�xFJкKĄ'V�ѕ��V9rH�X��ʕf��(�����u�;�jB�N�{Qʽ�s�I>b�s�!�rԋidq��y����6��#����}�܂��JԺ�&��b	���)|{*���M �#SB\d�D���y�jǹ��.��^b��G�n��;[��ct��3�c�_v�ר�=V=��^AՍ�]���DuO2(k{$K�؎-(�6,��4�_+�r�.�W[Bn�w���p{#g=R0����}ldt�f�c���E��.)���?.䩷�[5`-x:�y(������$q��DI;qy��ڋTo��1~]{�=��=�m��@9�u+ĶV��B��aWb������Iє� N���e���{Z�&o_mN@(�4Us36���|��Ne��tb<b3,*;�2�a�}��\WU��b��W��0�{��=�1rw���y�~�֟ח�PȯնQ��[R��B����KlB�R���hԍ�A`��hQ�QA%J�ؖѕR���BڢR�fm&e��)h��������Fբ²�(�+� �rዄ���R�Q-Acl��iTQ�X�V6ѕ��-��A����֤�m���X��c��D���-�Tam
�Z#h��X��B���[[[eX�[lYm-�
��,���J�E�(�X�+k`�V��²���-\\�aU�V�KJ�s��"��4Q҂("Ķ�(�TE��T��J\\"(�A8��Kea[��#����QB��PX�Z�ڠ�т�V.3��p��K����g9���(GjwׇOxy�b��Vr�X3&U�"
;k����Vl�ag9�v)t�FN��ܑ����ԭ.�4���++	��u�r�fR�_G}ǟ�V��"Pk�;s���r��E�c6�w{�JwN�Vw�î���y�55�˨!z��e�y�?�2�[FF s��X���=�j�;�n�c��Y3���!��Lउ��騛N��!`f9�{m3A,zl7�3��)VF�&MCK*T��v�_����y@�ȶ'm���5W����{3�$^V׹>��I���2���Mgm�ΉX���_�r�����S���횆D��{{y��`Z��S[��9��n�6֎�i�P�hh"T��E�F�*�;X��ԍ��y��c
�yR���WXIvA!m�/���}����z��'��s眺U��X��[���BZi�Oj���Q{i�J����S;�7*���}t=}�O{��z�m{��n�ke�i�!�Oqe�IJ��Wϥ���h�wm\�{����Ж�ڭ�d;��o�S��7=�^�l��֡��Ȧ�u�V�:��[E8{zU�6*���	�x��"���5�8/yڟ<=�<x���!i���ͯ�f�?Nt=�����Ոݮ8p?(kl�+��C뢹݌��z媼B�˧�Ĳ�Qm=��7�a޷�m��i#���`,�+�ֻ���ǡ4��5u47hۦ��-ݛ�S��*�;"E!�\��M2��:��UЭ�x���q����k7��΃S�U�%�
��	Y5���L��u�s{sH^��N�9+&_�
�x�j��eH�2�$��XTL���#�N^��Z��vk4F+�7 T۫g��DO�9ԅy"�Sg%��z]�͌�x��'�(eWOvl,��v�8�03���ވS4���u�8�7���Y���k�tX��r.��~�q]I��,�x�z��.��[v��-��-^�u�@%�&�U��c�q쳔����7�7�#�}+���ϻ9���4��5}A��MxZ��O���{��g��������1�{+��e�&<��]bV)�)3N�0G�zn�>c)�����{m����r����v
;��%Gҙw���ӯM��eGq���9����esTڴ���������O
}��7N�ݷ]a��z��J�Ի'`�J*�ɩ��ͼOo��������蠰o_p��t���M�w;Ӓ���O4(ZfE���-�|��O2�U�a��Pf�;A���*�v�B=5�aUy�b�~�L������69��6Y��'2M��n���@���z;�|ж�_���SlƧ�ݰo��i�o��|4n�Q_��o����z�uy�u࢏
�����s��} Z�t%�sq�b/����t���|��c:�;"|p�tv�;��t:iim)Cc�ʉ�\��Fk�ohg9��R�9�/z�6�[�'��4�R�E��{�.����b��-�*�1MeW��W#[��U͉J�B���7q��T�Զv8[Ԏ����̛��[1��_<w�B���L_�zk``�*)C괣U3��tL����9+&�:�l�������B�'��$t�#k"�#�׬a��A���d��¯dlGv�37 ��wE�8�۵���fP�"��5��
�i��-=��7�>y�X�
ā;��� �E�@S?AL�p��q�:}=��s'���� [3�f��g'��#���޵�&��\�dvC�U+�VK�t��؅�6�ט�ض"��[�}�m���X��KK�M���5fݞu�'�!VM<q�j��צ�zo��u�e� V5^jޛ�G'�of������7�Z�)s��Qq�+�|�����ԱB���1s{�ז[�ov����؝n���gTK��M�;%?8�۞��e!B�X����H��y��j~1nl�f�b>[s(�߫]��x7�����kC�3�9H�217���}'��j�~��鳱�כ�{B��j�E鮱u���}T�*W��M�Ō��HV��y�5���Uj�R��{Ա��m�+��y<�2f�c��ϟ�z�l�,[x�ͷ���Т�!>�ݾ&f�Z[z�5at����;|s�g+�JkT�Oz�����u�m�0��!v�A�����ܺ�e��wЩ����$~k��<Z��ߡ�vӡf��Bަ��=+�'�vt��9��/r���D�[O.�ϟbV��fJ0�x�t/j�pg9�nHhF�@D�|.�;Ќ�����wh��	>f��q+�n���ɪ��Ig��~�²)L��;UZj�UJ�޻l%�U��y,�oY��0qm���ѫ!��k����,�\T�ה�Ts�n6�UTtt0�Ys�y����hj���5DJgLB�BH�T�Ә�集�we@ٛ��{�#�����%=������Be�M�VO�:s��oz�܄く�DE�2o���-�^*���[AMR
��>t���vؗp����<��{�qV������{")�»��	��ӿ�ݞt2m�盏���{긲�-K3��]@��T����]y�8��]�bf3]ԞҔT��X����剨�]V�f9X���y,zn���C�2��8[x�uՕ�����uK~"�"ت��;k*I~��� �_X�����}qH<�bmޫ����}�^�y�ӳ»���c%�țK�r�F���
�ҫ8�]\ ��	W]�=�z��Ǻ��=Z�e�<b��|7��y�b��^�qŇ�o�]�wҜ��7.���V�=�[um�YؙzWt֑δn��*U���;��ٺ�ƭ�.3.���n�A�0��%7�VI9��u��,yϱU�����-U����2}P�8=ǿ_S���]	i�_���=�v�mU��J2�]=f��ĩ���$��b�KF��ﯔ��@t.�h;�mj�:���j[��*�W���w�3s��d�Ro Q�f5�%'o�>KX�]��;G,s�o<.R�"m��!�ꃹ3���M���T���</�R�TɌ1{7��:�
�K�iݍcf�!�xPp��Mr�u���warݧ���3<�ġ�o�^{��Tb�^�>��.�dH����r��BY���ΐ���EY��1�UR�U��^��b�	eB��䬙�r<jgn�;l��did���O<�Xq�H��t5�ѕ>�2���������Dr9&�\ ~�=�sv#�V1R�f��E��\�Y#��B�>����+b���2�bQ�9�f̔)��T9u�Y�Jn���}~�-.OL�z{�I�]]�˲�RQ/����-�/a���*}���&��!��㹷)��p��p�V]�5��_ڊ��^��\f��[��$]C7���������z.��ۈr��mν�]�@���ͅ�U�*�׭8��g6,�ݾuإ�����d�F�]zv׏�}�R5k�5#�%C����י�']����Myv=6Y>�Z]wX�^"��iǲװn�3\��f�1Oo�7*j���+��j����{[�$13Y��_�6���`9����-JW�+5�)�\�[O�����m>��VD�Ԣ���B�r�X(ZaE�E�lG�Si��R7��a��צ���V#B����3�Ʒ6cO9�wo]�m�T���V N�h�[����灴���/2����h��[��*�讌�����V�vR�|��$·�	O@���ݎTֽkP�W�_��cXί?OpCj���v�/-t}��ۙ;��CSIۻ�k9��T��7˖��^�dJn���B]lm1n.�c����2��*0�� �v]m�u'�ͷ��3<���5-Y���0e����í��L�@�N\Ҕ�OH��n�wA.�"+�^��J�6n&B3b��W/mow_L�cKaʽHX���eޑ�M���廠g_��]�ZҎD׌�eX�����1��o_���M��>WѦ�1R�9א奚7V�@�G���'[��x9j��Jn�C���� e{���٬/���S+�n^[7��s|�؇z!o9~U]3���{v軃g��J����<�N,�+��7Y��gg�e�{{���N�Y�Woz�u���)���v
�X�Վ_m��MΗ=tЈ+ކ��y�9}�!��o1}�a���nꚳn��
O^X�k62�8�����������ye�]�CX1���r�����{{4Ôнq����!?U������^����Ւy{���ie���k��aUN��	q�d؃Ǩ�5��L��K�m(��W7(U�/����z�{��m{�y*��F���G=;V7��T����v�|_��ꋼ2�����vze�W���]ϖ�P5�u/�.���Z2*��=9L��3�m�0�ؽu7띿(��r� <L�|+r���ݭ�0�Xu�z��at���L��u���VJe��e�{v�m���,��[�a� 2���%�Su��Z�E���������ڭY�hYʞd;!9[��{6w�w"�:�\ʞ�B����zy��QN�cy����Hʋ^lNה�e͍���˶0L�KZ������ yoX�u����AE(B����fʜ��ՍŸ�&b�ib�y~ħµO'�~lr��uxc��FEf����},�(?8�ۀ��,�G�݌NEf�Z�B{��x�P�u��)Ud�,ؚ~jȟV���i
򸩭yGk(G9��`��	uK9�V��^�4�ުb^�5c�7dM&x�.��}L��i���&s%aYo*ҭ�J�3��t�K{^�B@n�����7�Y"��b\�ѥ�pS�ĭU{�6���=R;��@$���++	��uӗ�6x�#=�y���ڼV�"���A��h䀝�
�<�N��Umɼ�z-L^CQ{KN�Ṵ�p�R,dt2��4�{��Yv9��y��>�b��Ki�Ɲ�%C~6֦��=�.���J3���\����^劺����qO\q�՘�ac�|@N�����S��x���=���اzR��'3t�4{FR�����XQw�e��k󜼍�IмʫL� `g69[à4qWajt��#1�7�e��gn�f��[��"nmu��4ǬX�L����2$l�w�*�n��}�f��v���k�pĀм�7b؝���M���n�i£'1�oR���ʫ-�w���mf�}����+��r�]o��6��?hֶg�����7K��������x�tb���E�|&裂=���wg�;\�s���#��	�����(��R�̨V��tUf��b�1�;�6 N�h�zӞZ��vX��m��L��g2�V���x�RaEte�u��2��7<W�e�R<u��*�bj3V'�1^�n��V_v��M�Т�!�-�D,����������:��ڪ�F���c��~2XP�7}�f���avו������xx{��BH@��!$ I?Ԅ��$�$�	'�!$ I?�	!I�$$�	'�H'�@ �	!I��$�	'���$�Ԅ��$�	!IHIM�$�	'�!$ I?�	!I�IO�BH@�bB���IM��$��b��L���(p��R� � ���fO� ē�%PRD����**RHRT�U*�R��TRJ��$ *�E(J�I!Q��
Q@��I
��R�G��MU�
��Ri$- �-f�6�m��Q) B@)PE#mP�j�T�jT�:�%v`�*J%B���2�B�{�$v���*@PU�6eY��D��(�6��Em�j��BF�ZU*H���(�(4	UUV�m�҈@��������p   ��i�6��Q�*�F�� �m�mU���Wl�5�2�{����i�K�b%��V�Y��a*�Й[[	�[4�l)�b*�����*U���   Ǌ�Fƣ%m�M�`ڂ�wb�kI�hXRښ�3����[mU�f���Zf��-��v�rِ�j����:�G�MոhhP����B��OZ���$i�B�cK�   Z�
 U��
����(P�Сq��E;Ӄ��t4(t �m�
�С��C9��(P�CЮ��3UKV2��ZجT�j�L��*J/n+�[mS�T�3��R�*�׀  6z�Qlh���*-�=�42�����i�T�FյmV��3@T�UV.��mY@֓)�%��j�&҃6�6v;`���덵��l�@-��lƨ�W� ��E��-m�S�1*0j5V��ڒ�(����m:s�U�¶ճl6ժ���Kk3FK+[S[Y�[��
iV�n�v�CU����v�Hlh3-��׀ ]z����lMR�j�T��R[55mSvu�kk4ҭ��4�զ�P�*ʖ�hд0 �f� (��΍ ��[Z�	����)(f�  6���0QT��QA��V��j��()C`�ѕVj�����@�.�N��P m�*���҂�^  � �X���e0 К@�B�0�P�7���:�(PZk`h(f Z.��Q�R�R�T������$
�  ������ ]n�i@څ�R�-�X�4[\���1@�mDf�UJ5��ТR%!V��%A   ^ښ��Ɠb!�M%��AjP[mFzq�e�
�˺��jVƖ�-��[ib�ʅ�%�wqN�2�eT%��V��kmJm��4RR� 4 E=�	)J�  ��
f��2 &LS��)Rj   �m��&@  �I6U)M40<RFc-����������X��NCF����m����1)lD��� }����oz?�	!I�! ��� $�	'�`IO���$HB!!�������O��c�aT��#��_ȱy2��,�J���T��bK77�S]�zJ�^�u����6j�����!�
�m*.�f�֙KPe��`��5)e����N�z������@�ǌ�sC�����դnO���	!w]��$(��3�L�4�B��7F��\2A0兏�Q�i�&ɮ�q��uvw�D�5�	u67�PҘ�+���E|�\�5��Kv����*�=�ؑ��y�G��VFj��V�h"5��n��*Z�{�V�Z�Uv�ͨ�0l��47*˺���@ض��A��M��o+b�)��ɨ@���fHStl��kJ����Ux\�Yd���Z��{Lg��)Z�q���FM�>�D�cPa��Z�XF��7�#�Yb�@��U��i�7*�p�;r��ۣS/	��Vb:��٢�K�֬@�J"�S2�h7�]�m�Q�թڐ˧$�f���ʫ� ��̍RӬ��mO��7]��5*��Fn��xF����ȶ��ñ�Cou�#X�,+�/�� P���A\�[�T7���eG;�X�ޱ0�9��3w�.jufM�9�jfua�f�w�����U����h*	��wQn���<	��jx��6t����D�ڬ"�fC)n��H����f��+�c=�X��;��f�d���a�,�pZ���v	'����++kYԘ�/lD/mE�L�����k��7qJ���9ja���l�#A��Y&e �SL؍m\˃#��N��t��٧c!��sn��cV���s®�V��+��t�	��$�J,ѭ5)m��5š��Vf�9w�&�s Z���L�	b��k5Z:^iҥc-��t �E2�Zf��#n,uB��z.]Y��B�{�$�5Z�v�M׹��2u[�ɼ�r�qy���kb�*4'�pTb��N���B�����&\�p᷒�4��6R��FS�B�ލJ�7,�SdD�R�a	�J&NJQM*�)t0dХ�5�l�iSl����aM�Y��%�G��$�\�ʤ£h�(�n�ڨm�����Y�{�R�֍�&�C��xe�����H����sM5B�қp�q�
V�CtM����U��Ս���d�.�#�k�Jl5r�]B��#&f%VpҨ6�/M��xq��,��U�6aK4S��mB]ȋ$�mE�\U0�L6rG��E��/k�*Uܚq�3\�E%� mU��0U�)_��)�x�\�ua����b�C�K��4���ňi5H*V2�9D�xV�XI�whQ��b�;�7%4ɨ(��+������"#��F�M��b�nm�,�6,�/ohS�����\�U{X�x�-����I�[�Rk�X6-��S�mݯ����d�;b��%K�^���+K�3DD�z�-�O^��M���U��������$+�V��պ5��b�1"�`,۲(�,Y�Z�p�����|�+eѧ%cv2������P�sϹ��ޫ��(n}R��+4��ܛY������y����cX4ĻEU���%�
�o�N&�ke�ږ���e�D���t���1���6�J��)�������Qz�3�P�(9k��nՠSl��JF1e�ܗ�mQ5��R6p\wǔ�$���1��SE�R�5�����Sa�,��x�j��m�cڬ��1�dÙi�5�a2�Z��ld��3j�l�b%����h*v��B�� �- �
�ܧW�-�ʛc;��I;�0ӃA,f��
��ԅ٬�9��h���N�۴���*�f-nX�r���~��aX�� (���y0i�`X�-�V�D�����[N�����ޢ����Z���R���]�{��7]kf�8)���q�B���4����sii׉Q
��-j�L�g
��7hh{K-�B��zl͊�v�/6ӂkyQ�V�R���6Qo!��3Y35*gD��Y+,f���j[f`�1�W�[k���֙p�$��6&ٔ�
w-5X��Z��3z2A݉l���fkC�N�l:A�%��,��)�pS��XT ��4����0h�E�w)���2�f�76b;��4�+�aԕ�zy��*ӽ�M�Y5��rO+-�v�j�kf
�Y��x��ͩ���o�gEf���o5Ղ�г�\$��U�l�צ�������	ـD%��*��uA��]Q�2���d�'2<��]�:ݙz��ݹ���sT
�^�)�;��â�����m�v1�D�f���Xn�l"4c �+p�b�ib�˖���n�����mڹ-4����E5;��cy� �jU;�w�$AةU�(]J�e����d��Vr�h���[�5!/��.�Z���#+u��\��8B�/wc�2��l[���Ŏ5$��e֍r�cf��v�n5)���u�n��$7*�+$�&��a�S��e�$�H�-���tݮ)r�$v�m��c�e�M/D۬����c7N���^e��&P�[Kh��˚0����9��lV�
��s.�̙���65�n���L�֬�(5էQ��
�Y�̍`�5w�#nk�z�����v�&���b�cg ����y����MyYF�;����qa²�c:��06�U�Vme�+&16����ɷ�D-K��;�RԠ4�����LA�&j9�e5Zp7����v�ƴ�W���vd�V6AFnLe���F�a)���j�c�~"ݺ���Ql&�\c1�G�v��R]�+^E�7��RF��Z"��;��fV��CaQ����oF��2ф����,R(�����j��CŦ�l�b���J�kn��2�=V���1(U��hR�W�P5�[����3��f+��coF�ۼiU�p����mPō�v�������pX�k"m7-��ѫy{a�[�>ݲ���,���L5F#N�
�զΚ�b,9��f]�ؖ���T#d�+ Bi�	V7p�v�m���^`&� ��+)YYtTX�r����*R�cmĐ�*,��Ei=���aJ�^Gf��ز��G�Ĩ�����3�```U�Y��.���'N�%�W���f�)&�P���)��4ꭶvf�4K���76G�r�Wr�:�.4��V��G�*�(V�v�3m]�ɵ�K1��B�n5���A��ofj��k����e�XÔюٛ�f0�.���Xi��ϝi��th��,��6��'cM�5�y����ľϵ�(��NZ��fnmF/��!�q�w�^�:�����������*`����dj���I�����ܧ���4�ӈ*��8����(T���Ҧ�Q�֊�I����)�gVE[Ish�<��.,lf�%��O v���Eu�5�ϥԉ�ۤ[Ő�1�KA�6u��x��C0�4������K��,3w�IY�v9�B�NH��v{�F�40���t�e��H����UmE�mĨ�ͼ��CT�R�j� v�&m�8��XWe�b�wOU�8��k"�buw��<������9T(La�50�͢o^a�R�P"��iٺ�2��j��GIU��ղZ;{5��ȥKU�4Gx��fى��55�Ҏ��n��	��XoH ��1х
�kB"-8����S���!0��i�ݥ���2�{�C��m-�DY��^jO5�0)o�F��6J��9�fW�fReM�롸�jǢG��e&)���*��)�L����v%�̕	{��J�e���.����n�ݏ!�]���Q�Fbs
���Cw�*ؔd�!�CoJ�V��v�*�afQZ��C���1���U�d��^����*�&�R��cy�Gq��n�2�a��Z�%y�� ��.,���.%�x���U2��h������	_!Fe��UC1н��4�hc[�Y��ًNR$0��H�B�tEZ�B5UxT��D[X��M�Tv�]�mCOe�q�k�/�� ݣqđm�1�^.L�˛���vo���7���̀�B� .]�����iA�SoL��Y�I7Ɓyg*���6v�n�,[�fd[QI�&�8Ǫ,S���Z�0^н!.�h"�^70}��K%`�b��Nէ�-��ܻ�Lv���MT����r�Mi+�~âڽnhZc�y$!]�f��&��FThK�nS!�p�j$J��V���5�����v4AY���M��Q���Ő�զȓ.3d-3�+���l.�tfl�b-��Dխ�4 �nb�0l0��4��H��!W&|oi�5�G\��l�ٔt�a�IN�䚚2ݼ�Aۘ.j:᫸/@,IX�4�b��
V���#����Ҥ���{��4h��'mf�`�6�7V�`8l��1H������Tڽ���utpn�9L\Zv�4%c"ZSӛSM�F���yk,�������X�5���ޛ�.<f\�`kH\��V@�̃)k!1��EKt2�6��±y4��K[�
���˸�7��Z�C>�uJ�:�I�n:�Ϋ_F� �O�0��WY�9�c��f�ua2�\�v�� ��-���l�	�jDm��)�%y{nr�֫),���� |��*�=��U�t��f�BE�@n̋l��(�Y�������+u�!��;�X�̃�.~�pj��=s�͑�����mG[��9p#Y��Xu�1�6q6�Z̥Y��ۧ�D���3,��RS.7�)t��an��k<Tj�o5<׍��${�e06n�Qk.�+of̈mȅ�CW6�Zap���"®�u���.�"f!�-�;�96v�DZRY{v�"]<P�W�KY�p�.��Ӭ��qY�d݌��V��r�4�i.�m�M��&ґS�6�qM�4	����!B��.+�h�FA8#���
i�fM��x6�e"�/�)b[�0�i���?����l!���k2*^f*F�����(-,RU�~+B��̀���&���X�q�ʺd��i�:Rt����$S��Mbs(��}�E��ܧVS��n��X^l�K��X��AI�CMk136����G�a��i�[��W7uG%�bL7uڲ�ygV�6]�[z�n���CE��3`
=zDI�cND�KCqVKJ;�wX�B�j5`������e��1�2Y��q���m��J��6��w��PyH��j��nG2�iG	�C{���X��h�Ӌ��Y#�s�Y����f^��U�EYw�.�"��n�	Q��,��N�քNU⧊�RC�k��d�P۽�)b;o�i[�kdч*6���y�h�ŗ�KT3>��fdAۖiS+N�X8�fm4*����)��j�&
���Z35��#r��+q�cLmܫ0�,�z�,��W���M�r7Ll�íM[�S^#��2��CvU���1f#�k�]G�}z�]���S�F�:�S	N�*�M˽o\�Z6�n�0�[�
�w�0b��[M�K�o0J���h�%e���KE�#q��ū��͵�Uuj��%U��b�z����aP��ۧ��U=���'F`�n�gh=�Z�㸣�ֽ�N�X8&��[-�{��
1�X��;���*�jM7�Bi�ܵ���5�2�'VL��[�GB�1�i��F6��.载�tygp-�B�Z�m̶��@/��LJ�wn��"Z(u#Ճ��PKDl�ȫcM��i'%��T4�-�ʭˬd���q]�C7V�l�u�@k+*�6���d��X޺��N�8�p��q�p^%�ݲ��YqX�gD5	t���i�{	z.,�$�Ֆe�.��X��f,E�X+Q
�.��w%��]���xt[��lm˴]�Ժ;\Q�IԦ:�@���G:�yB�dƃM�۵s�Ԗ��S�.jHඝ	v����3���5!����C��+p��csI����"�-�Y�//ne
$iM$⫃SX�����,�c8�^hp�6�Nq-.f)Wt%#ck�&=��×4	�P�z^X��wF��vCe�ac%J���XP�p=��؈����5%ܵ2AWIH̋)�bR�W��)!��I���Z�nd��͍p-Ʒ��Y�M
���j�'E8Cbw)��`��ǿm^ǎ��
���F��^�Q���n�}�a�.黦�T-���J�U�eH��خ�U�K��ڬ��r�IX���4a�����;��1ک�-�֩���݃y���C0�4���G��i��ցJn������aԭ��g:Li�dU�L�1�9�{2���/
��#�&�5I����	��B\��[�t��.�9�0I7r�C�L&�&m�l�R������7e�&����GD�x�m
�
t�
��GM�^^�i�b�)�b�1�fR��cpX��Hݺ*�ǀ��R��c�5jm��s4���g@
��M2�X������9z�f��S�ǚ�Z���'b�i��	h�-�vێ�7G�J��n�3o[�Jb�};��VtD����a�f��2�ɬ�9�bJ%YImh��X�R@�s*&��j��r෹��S(��o���`���t���k�x��*�/�h匓0����1xP��+֧&��;x�E�k���^�-�)��pYF(7,:1<�N,�p9�Y6Q̣$��KB@jdʠ�+#OGo-l�!Rc&Mj�R�[b\�j�f��Q\**��S�SQf��؛yj��%�V;N(LYI
��1�ɠ:�,iŚf�@wf-(�X\�P�n��$�� `�i���HB�Miy�]�t��&�R�9����l���ʧ���G����݅T=8	���ʱ���6�wov��o�=Ù����86�*�M�+�:�x"{�17�)���=�r@�,��d��x�տBɣ��fu�n��V������g�MK�B��Z�JcV�ݰH��Ώ��YJ��3��v�]�G6�G������w����ᓺ����nG���u��.�$��yI��+���uhgt*�-���!�j�NR�n�w�Grd(c�c�l�4;�	nCջ�L��A��|_��2�Y_���:bm]�9�3���{Z���4+]���"}�x��V ���}3��O�͏6��
�hL4��{�1-΍�r��=�ޗ�Z���Jc�*����
�Sy�ng��
�5�8w�K�k��#�t6��@�nm���ι5�Q+�#+;�s����U%)�O���X���f����|�[�EJҨ�Ǩׅ�h:�j+�Orn���<�}G�c���h�.��\�V�Q������O+{���\�HU�M�t=�ʈ�	]��Ǽ:���,�,o{0��o�D�C4->ު*�
7�������ѼD����o7�1�>}$��}fm��]�7��w�qE�6NV"/%�S���6@�*M�[Fq��v���ٲ�0FAΫmP�XѝR�1`�����lG�z \X��'�}���Zʝ\���ЇEf�5�{o	w���X��S���Z�C���Ŋ���ۆ�6�FNH"̳�{���㪩����fb�m�˗Y����|�b8�uѴM�׻����oXs�ItX�V�1�1�Oxs�� �b��e���ciKv�)1u!��xY�1���-�v�Vܡ�4�9�V�����f��,�j̬z���oK����և��2��j��Qi���eN=���Ü��j[]��y'�gn�d����H�I�R���̡���թ+L��f����<��V\*Aݛ\c��E��R��Ѵ���2��vM@��u�r�M�7��CG
��ӻ��V�<oB��8�H�=�l�[�-��ÜE<�nmۮz��;
���ٓKbjZ��_}�ڰ�ڮ�����W�y������E�_]�'fr3WJ����RV�v)5�p�x%#RM�1���+=+�R ��k��2>���9T�ٻeŕÂ�T��͂�gs�7w�޺��4�5�}P� �\u���Z�.���MҞ9ƅ1�ȑg�z��>ޘiԥ0nfZ�K��O�����7.�+r�䣾�y�UJzr��FM���H6��{1� ����9�\�Z�r��,�����ƨ��	��a}��ŦC�6�%N�Y��ju�Y/M�f�p���1F�W�YV�Z3j��W��OP�u���e�oڐ�A���̃WDN�C�MX����Vj◲���%�%��uvM�!���3����h��Y���A�}�9���N.Y�iJ�U�Z8�s�|_֩,1��n�ш2P���t�ozQ�N���ctվ��c��Ż���AV����7@�CV�*%j�d�M�@�N���:��7�l����*f�ֆ�3�z�>�%+5��H�,v�y�ԽRC7dկA���w\둈�G�w��I{�{��ۻ��A���s/�t8 �5�s8�sX���Q]^r	���O-��Yal��9�\k��d	�1"!t3T*�n����&�0j��6)��p3ۮ�7�$���q����o%��.�'gNn<�J��u��܅�v�Mȑ��}yTn��S;2�7|�2��zC����&�̖��+{I��n���$��	jg�^WFv#*���{^�+��BAp��ˮoph�e`]J��ۙF�w�9�~n��y�p����z{��EOv�+ڠr���NM<uǌ*,f�_�6��ȳC�9�87X�J�/뤯>��^cL���-�7����AE�k���Y[S�ڗ0Q���՝#�J�;�mtjv���,!�>��$��Ҩw���x���fUP�Bo|�l�s�u�w<D��^%X:�}�d�9�I&Q�Q2]SM�Ы�}�}�y������u�C9Ĭ��N�3�$e���Y{�Q=�+��,qD.�� ҥuq��	�;7���1��f�Q�se	;�ٌ�iʪ�eCiӡ� F43�i[�-�G�,:b���Z��%�a���:����%WK(C1�k���.u���o6�ӽf$3w0�"��q]�-����$9�FX�)ں0�38aWG��R�i�ɝ����Z~�5m�B��:kq�^�+�'��:����澾�[�T�-l:�W!�����1�Yk$��h��Q-�|�����t��{�VP��
���.�m{��˺jn!eXƜ�,�thJ�*a��կm�5^��	��ں��ؽ�𷳩�Cu�r��r6��yb���8�z�¦]-�W<��Jlۃ�OY��N�+r��J43���µ��-E��<-%�m�3�Ř�޺�x<i�eʞ��k麞�2�lx3�N7�g��X��NX�B�l6]����8S���peL\���2��W�N�뾤釭�kf�@ṹ�>W���[���ꦬ��(�#Ʈ��p�X�c�c'����]�j�{1�<��9����VZΫ2X#$����)�Ġ"�!G;�_>�[�}�=xB]�$�j'l�o���g82�;�xq��$����f������Z���IV��Sy��.���^�ݫ����[L�ԖS�J��[��|���Ξ�q�"��[������J���Lޚ�����jL�y]@�{��mN��I��*U�xƩ zVV�7��j#2�Ř%!ʐ��:����Zqc�Hʕ|��vͱ�n'go��]� tF����h��O���e�4h�0-�L�ɔ,����{,�����P���5,�̇�e�&Ռ�	��5��|�x�~ťU)i�nT�6�z�\�譥O��=f��@�]�˭VΚV����D�(J�v��M���eʆ���T�ف�R����}��In�`'�^�Yж������)�wt�f�<�e�i���K���ա�y,p<�3�ٰr���W�h�͂��-�خ}:K�l8]�=�&d�_�Tch:*�h�]x�8��N
���7�ی
��6�W��J��6MC��+���	�WԢ�]��8�݈]b��L'��闌���a͇��;K]��H��'`��fgQa!B��"� )����ɐ���)r�F�������U>
���Os���5�efJm,����j|���-T;�k�hvm�8����Ч#����nY���X�Dv�7ntq_Ȁ4�ʰ�[9�Y��ݡ��T��Z���V���h[���5(r�oB�ᵓ�NF�#Qo$t�^o=�W����PROl�t{�!!��D��[}�-+7T�7Ek�I��&'��E��O)��;n�����1�)�8�`�>M�H+��^���#z�ui�sN����5���B�JT��7YƜ㓳�]vk�V�7	�z3�l�o�[[�dgM�x���#j�KN��f���/����r���s1�n�-�:Inq�%+]�@�uGw��I�Wf�]�'�e�i��wuiw.>�9B<3��}�1>��y�y�u"����W:ڬ�����׻�q���ܕ)�}�;�4d�t(A����Wr&�2�q�pˁf{����ND;�&C4�av�b���v^ve2� Ł	$[:��v�Rzdv�Q�To�֡�nl��ؒ�i+�{W�M��.�@q�g��o�;��� )f
��Mq5ݸ{j%����\��3PեŪ�e��ө|iU��y[}����S�%Vc��"xڛ�f������}*�ZkWyQ^������R�uG���R�X�jj\u���h��3��$Y�:�u��P�ݎ8��;k��ȄkT��b�wk�t�ID�Ō<��^6n��]N�>{M6�h�z���f=���h�	M�4þ��i,Vn1��n����7�n�X�A�1��m�(�i	
ͧ�c�L ˴x�DviUu�j<�a�7/U���R{n�Q<ŝ�{l(����#��M�Ɋ)݊M�/�>�[�4���~˺�ɳ�i�-�S�p�<a�*�Y��H�:�������}C3y�f0'V�̀����/
r��[ôsݥ�ZXʑ.M<��(�vأ]�n-�>��v�tx(;q��L�<�Q�*Q��M��x�%K�{��.�LYŚ�R576��l�CxP���F�����
��J�!��*�^���ܸ�{�u�p:��+5��.���NV�9�]�_f�;!����-�ӒA�kX&}�(R�=cI�C&�����2�4��x�֮�I������*Ǽo�Z�L��������
��;j�\r$ɩ��Wݵ��g�a�/`f�
|5IoI�AL��}6L}{�xT�gUE�7�)����A�i�	�[��m��Q�k%ټ9;�m������W:�,��>�uM2���g)΢�*��gR:6�U�:��XrV���:��0�ɜ��8���ȆR���O��zEh�ڌ3��ݗ�:x�ƻ��)ݜ΃f�i;;8��uEͥ>�w�H��/����}y�,�#5t���z�6�3�M�Q���˖�stN�ڦ�H�ǚ,q�9�X�6^�O[S��m��:�/6��TN�b
���B*�kJɺ��.�������Uf��؛��.��R9W)�V��q�we�^M�uo�R\�7��z�l&pp���<�1�ztV�cy]�pj���WyhL=gvYu��<"T�s1�e�ws�C#֐�ݵ*mC4��K���������gE!��Ҕ����LV��)�40�9;n���/����J:��#�����T�
��V���X�A�9/��Z%k"M��6���P�K�l2��\�z*�voZ��s�-���OP&f�;8�Rq]��v�l}��s"�P�δ��9s���:�S�{*T����qJ�ڃ��ݻ�ˡ���0����� w��m\!�8r�_}�s�-����6ў�!c���Z�O����vJ����y��;��D�q_N�̢/^t��f3�j�ѱ��Itk���u�U�p�Ν�L7+&dS]��f��<Ov�_<�Kꋯ&=gLm�
%����[N�u8�盷7N�K��7i1���u_@N"�Û�G��U��U���D�Uŧ&m5��A돲kb�q�ո�s�2�8NQ��(�D&�i�A�9٤��7N�bk^�W//�NoH�ќ`��>3�h�u� ��e�b�>��XUs�˔�����u�kC���ߪ]�V��%FC�d~S��t+@�6x�>�b��Q�&=�.�Ѵ�n:��v�]T!��)���̫��o���	�Ns�C@��!A���k@B��J�@������vf
�o�Ҧڣ%-כn}�%V-��˃�j��ބg-�4//C���!ǣw�n�Ӆ��ͬ��R�=K:"ogӯ<�Diܴ�=vyP���N`����bv���۫��OMs=AY��R�f��}v�����|'j����u��հ4���5�4���W�n�[��[����/��)�k���3��ӊ����M��Fͽ��r�kaؤ�DI��I[P]Y��r5ԩR4t��b[���7%��ϕV��1j�M�g�ܡG0���a�Q3.>�X��slܷK	�����>w;^�׼Vt�!Ԑ�;r��)dVi��L��%$�������jH0�_rm���$���[ug���ce�| an�����y�T����o7�ݖ���D6
��	��Q	��䕶ʁZY[�w1����;ʴS άA�	��oh�\���u_��Ktxs�H�f"�2t��R�6zZ���U��y;����ɽ���v��ғ[Y/��żw�Cj%��J p��w-�}�xL�UsjK�;qf�����A��X\��v]t�k�K���qk�>̲��8�q��^wMΎs�/�a/�ȹvh��Ӵx��y��4����o6��Э=�N'
� �Y��и�U6�N`բ� �2�D��� �[����y]��E?��V����޺��+����%w�ѷp�S{{�h��{t���c���4a�+Ur��X��Ӷ���b���<����jV3k�*� ���K��u}G�]׻�|ޟ_��˼R8+�p���L32��G�sđ�X�]�ɼ��-���wt���9�=����o��M��E﫺Qꆚ4��x�m��!�Rn�2����&����:E�G�"�w ��"C*�q�2���G�li�[pAm�#/�՜�p�������eX�wh�\`A��T2A&�j��~�:e)1�7ȹҺխ�7I]X�CGqOH/��p�ټyZ<�G���ou��I'�6�9f�5��Dh+kHwsW[Yq�y�n�wnFvY��)�Y��M��q���-��e-Q�^[�6�U2>1P{�Cq��_=P	���T1�-��@��	�!�I�A�����Ύ��r�-�YS;!	�w�i+n'Ѩ^�oI���DK��&^S��NwX��]53m.�Ԯ�du��9C�q[ ,%u��.\��)��[qw8�4��a���AS��5|��:�D�뽬�NI�O��:ty�R=����p̎��9ؙV�$[��� ���hR8a�Sr�w�9�q���DL��}����=�j��Vn������d$����H���{��.��eZn�z��\Գ�
��sXywҺ��.���߾ט��߾�8�HH �$��v�o��*T�7f�.JÙY���pk8�a#�t�"]����J�0&��ڼU��,����L�BdUD���c�Bsi����zL�ի��nlB�UͿ�et�ᜢ p�jn|���9���J����]��)>0��&2�tykM�(��;�l��	�ctN�:�GOYX�<Xi�[7T_]6�8�V�>���=���.�G��ܾ��j���73�Ú弨�ZQ�)A/q�L�<��p�*7r tÑ�:�$�u�O�%�n;$�o�
X	Xk���2i�g�a�gFo͢�}�mXK4'���kt���-����+��\
�Cz�@���H���hn��^N�	2�Vs(*��G'>�����iWH^�!;.�6T��i6`���� �}�-z�5P	ϟO#�-��6\0�\���b�ZȽ����n�=8��q���mɩؠ,v��ڥf)T9�������V&�U����tc����p��$�iWjT[@����y�7*YR��}հ��B,���Kmu�UbZ�OnՆYc���E��ܓ�y��x�Եngb�2k��NYT��Z2n�P��Ghi�%�������3��s�:�óP�W��E5sZ�.R�YyGzc�pLO/�ݿ�!�zc���n�l������t�%Ǆ��z��m�1oK�P�&c9}V�a��]ZV$�S��k����=Me�"�����D�+	���:.-�ɻ:� �	aJz�	��MqR5,\�q���a�u����a�����C�7�>Ѱ�r9mga�B粬�ǒ���Z�Aes���2��Q�R�nx�]}!mR)�EP�����;��l���,�*�&�����|�7|��T�u��ˏ�®ԧ^���]02�x�q�u9��8�u�gP���|�jױ���ye*�6������5h�U��,s�]Z,A�W[j��=��+z���*��/����bd�BF�m��`|�����v̫�L7]BV�j���ҍ<7dp��e=����VB�C�Tzb2���VT�㶳�AZK5��� �$1�I_Q�;o7pp�3Ҵ��!��%cO�����K�a��uu��y���غ-�	fV�/���[�ʒ�mo�1ds0��L������F�m�weŐٷ�bR6sg��ʹ�O�Li=�"t.��U��@�ͬP�wD��Ln�gd��L��0�u�j�PY�s�`�[��eއ���K����v�����X�`�v�x����7Ԡ5fpF�䩛���Z��̮�&�x��G!�ڇzЃGwwn]*ĺV�
���p�x+�1�Vgd�m�lU:��}EjP}�����5��������  T�M�d�: &.�t�o
�w�>〮n%�S�2t9��'�Z�qƵ�9c6^ٺ�X{%Z*�rAn���b�����
ͨ&����n�i��M�O���*��/t��t�goWu����cӾɫ���ѱ��p���ke���a�8��PBMx���D��7Y:�/9c�n}�n�[u�6��j�^�}{]}M�c��h�l�	�,���ad�j��M��M{z�#����T9@�u�vʱyY����9��8A���Þ��ڕrY�O {�k�w*}�hZ�Ə^�ٝ�t ���fQ���݁�2�w���a�A�u��Mr����H�����������Ӿ���F�\A��vm�r�]r(ά"]�#��g�e0w����[mS����2R��������z2FCT���NN����wwLG@��V�kIE����*K��-�b�&i��bB[vl��]��w/m�D�j�_��G�>�u�0d�
e��$�U�C9�wTF�A$v���F�EkZ�Ƌ�}��ۍ��6�p2�D-�D��Xv�]q�`�i>�g�b��|���=a��:�X��,������D��yq����q4�����°�����n�h�aʴ�w6�ò��wV^�[ b`��3.�L+t����=K���6��2��*��t*gJ��UJ�����i��A�yf���NK�.��v��Y����/$e�qu=Յ���Jg9�Hc�(wl�B�sAO�CY��^YW��
AE��k�+������e�l�V]��n��aE���A�q�ѻ�RU�����*�W�sGpj�%ދHГ�[�	�\<��X��F�����vây����d���5}!޺���vf��6���vlŘ���e鷹)�����%A�����'D%�;����݂�7[0[��Ϩz���U���BCw4�-�V���ƁfV��#N��QS<���o��o������ZАs���-ڏ5��#2�"�YiR��|�k�K�'mK����+�`ʱ�LT��E�ʁ��{�['<nٶ�C��k%ϖF{%��ۺ0�(��	o&�@C���N�)U��0��J���rքʸ-S�����B/�_5ê9n�f��F �h�e�YV���	[]I��UHn!�]��ft����\ܺx�U8�A���pV�����ֽ.���x�tڄd ����v\bf����wa�7B����ngG��5�R�"����yt��oDw[��3���yY�X�w�9}�8V�*�`�	w�ܲ�u�%R*��_n U#�-���]��r�Ώq������s��i]�D@���/{��=P���X���#*L�(,�TY�f�J�W;w���ۥ�|Q��/K���wn������=I&��gC}Q�V���;ۦ95��P�t��9Y�����M�'_u�!(]f͕�xЪ����;��4���Ӆ;��l��6�ۥ���̫��m�a�4����}��*�>����K��u�R��ޭ�f��c)	te�yVχ���'W�~N�n!nS�;�=�1>zvٷ&�{H��}�J
ޙ{�"%�e�ܲPz�"P�QN쩝M��ԡeQTB���Sl�;�4��պf��41��uڦ�I\��Y-�R�(=����i ���wR��br	��P���)e}�i���sb�A��������j�"�d�,��Ϥ�(�XlG���y�H��G� ���n�a=lmI(jpx3�
:�s����=;���3�
������I�������N���F��* /:��ר��v�������|Z����+GB�����Bz{QL�}v�����@����?LRW��>t
C��k�Ԯ��׉;�8l�7���N���R{��K�Ӆh��ܨ"�A1���8��{��֓�\�E�7p�-���>7��v:��U�^Ą�OT$�E���&���}�\�2_
f��Z ����H�Zz�Ѵ��7BWGG��j�]Wl��@^j��z%���x�k�i �8<�r}s���='��q
׆�ݫl��b�4V[ p��7P1qk����bF.��+��t��A�H� �|��?���{��-{+��%��3�E�Q�2�`WM(�M7ؠn����U}t�]����d:�nf8<�gv�9�ѐ�޴cD�ম��㸊�-sU��v7TKBf�h6񑜐!`��״1��W4<!eĥ���7*�!X�ҾRՆ��V���L\��:�˷J<anc��&�Qja쒩�vsVNKfoCX��F�%�ӳ�̙�����9��2���[�Cv�.�����́�B� ψ��TA�t]k{r���C��d�m����!V����Z��^�Ú�ži�\�;A5�F]�i�ry����mm�)�Z+7X�K��5�XkD��G�}qvL|}#�e��Qʇk;��-�P���M����â����ѵ*���<;}�on?)<<��չ(l�v�Z���ݖ�(�,u�d���8{^]������ĵ��Sٴ��OI;k�+r�0w�IC�����N
eVi��oU�-,cy�+���NX��pY./�ҾU�u�}�8Y��m�ܗN�Z�����9��;�iȞ<��/�mt�a�M�{���]�-C�o}�Bt�gd�D=<�ݗ�]ګ=�%�+��<�*p���0��{A�uW5hwmj��T��@��W|����i�*9|v69������p�v&pq+N�JR��"�]da;��<b ���iw9�L�vMv�C�0j��Z,GE���U&g^�O�/6�M�|s���ب�޹�J�h���2��Њ\NǘN]�]N4yp�jEl���x=��-#N�j�Ļy�L��5/w<&�*hV%t���1��db���Ee#�0���Z&T���wO��ovAe��W���y�f���N����<�H��K͌�C�ہy��-�}w9�D1��M�
�L�=������1_��B-%�7������n��q���N���]oi���ؿ���%s%�k�Y��k.@�\hw-��JL���w��[̧�{U6�qۤnc4�t!��Y��>W�.y��d���8�d7	v��\�B�-ʕ&��D�S�1/ 脗ݤnx�!reۏO;w�/"�&�!m`���(,����rʓ���b�Am�Z��Ȑ�)D�6o)5���ner�36�ip;[c�&q��q+ʼ5�JƵt&<�:4Zd�їr��q�6Oܬ(�sI<��ظ2-�f��1m�r������ӵ�]�nM�F�TZ*M�ڟ5Wۀf��Ωu)�܃N���G}�]���f Dv�[G&��2R�9ztHl]i���Qx�E�����]a��3�Y�¡�{tKl*��N=��oǶdlj�+��l_	�}������8����G1��>.d-fI'��$���������J� ܣ�\���w�g������#ݯ� E*����û�����5�b�˓v�p^6����̶W"������V�W����v �4{c%۸�0�[�VYD��o��,��a��fSF!gh�ȼ�y�"w�*�2W[!j�pΧ�l�PU���%�1s� �IMY��h�V8��_P��ܶcp�GigPr%n�j�I��X�~�4a��Dj��xB�D�����֭����&�aw+z�0���NϤ޴8�A�E�#��wI�����x�a��ÝRl�	��f�Hü��	w���ܣ�n�-�Yhd5�$'r��Þ��稭�w)��d� �ڲ;���k5�$d��Lx�.7N���u��Z�+qؙҰ1��9��uQ�ͫ/�o��C+�Նl�3�X(F
�0U��Rǵ_�c��N�LV��:wk��J��r�.�YJX.�����a��(�<�4/��.��梦�Y�T^XNS�pl�	�fD�I �^v���B���롊��9֮�c��#!R����u���pn���-�E��*Q�Q�Sq�L�6�ǗNM��8��FJ������41Հ��k�a��:�}�V��mteq1r���ο�W���#��x�I��}[»oY��8r��M���ƾ/O�`�	ߍ�N����;l�!�E�5�(n�Ȩ�6ޙ:�N[�b��e�Jr�G�\C��U���*̣y�B]`.^>9�"<I��J�z���9gX�I����k.թ5���.��8�V�G)�%�X���E
��Ԑ���_<|��u&.��)�0�����I�nV푽&v�	�l:i8d�ܦ�Q��"����q��5(���r�T/sxJ0��}�Ϭ��^��0��Aa���$� �wv���t7�[���*�#�X�ï�2q�� ��^*q�Y])�8i𛉉`�:'u���]`�K�������0i��g�{�N�ޤȻ2��o�&�$��vJ��Ղ�-�cr�i~�/m6�y(��{"]�7�S&�Z�7®w�4"+�:��hx_:�x$��ӝvV.����3��U-蚍���܇E�3�䶦�~&�Np:Z	^�Rv&��� o͊sy��t[�7|��(dF��
�P=���ήT���5�EQ�[S1��w�v��L��9ک��Oxɤ\}�� ���Ζ�u��;�+}�$t��ء�[������AY�wɯuu�?%�1����Cc&�i�o3�X�Y�V�X��F֊�� �\:_$����:�*�N�/�+��m�=�����C��h����d�F���v5���23Ϲ��
حK[+/D닢5a�&Ԯ�vw��/�`J��[nQl؃)(�W�/l���ħ:�.ٖP��ַ�V��w5�bUӒ=����w��w>�Hwג6%^�@�MA��ɉ>F����w��^�}]�hp%�m`�uR%M���Zl\��(%b�G)��{�i�zؖ)@3�-_A:�^�.��<س r,��֓���Yt���2��]˚A�����*s���V7����|�ղ�"�#j����nc�x�l��l���'�55��0������Ih�H��TPxS�fй��y��J.�j�b�ɍ$Nib���Fl���p�_Q�����f�lM�YuˁtdD�ڋ(�D�دk�����:o�b
p���8hho�(����՗�pvZUЊ�t �|{��Oy�CK�F5�C:ޖ��-Wa|e�%X腏v��ךs���=Bw�cΧ�{�L�*��2�Yh�-��v�Z5���x9i����Beq�/ M���R�b,�[��,T�}Y��5�t�V]Z�,%��Y�f,��ۭS�>km{�<�#�u�S��_��� o5vaI�on��K�]2�d����;�[��PXKkc�u^�=0K�\����>�������v�:�N��}���a_Q�� h��2��
����$�Xe�e������Κ����޶���s�x(������?���$�M����a��y�����+_����t"�^Sg+,"לhEh��{F��F��՚�e�8��Ⱥ�^��͇k���)�ܾ��;8����3dg�nԽ6^)��WQ�ڑs5�鯲��ֶ��K1G��vҔJ�t�n�����k8��0�H�٧
����ub�܋�<��Z�ʱ�[�"��u���]ճ[̗nu�!�Wy�
�彆���z�cu�"�i�y�遬�͕ß\{�_[��Õ����o������\a�Y���Wv����QY��D�����5t�G����-���q&f�{�Ŗ3UWY��9�N[6)�[ oJ�o�s�Ѵk�O�s_�P��Xk��L�o����]๝�ّ���HN�~Ա�{�[��X/:o�O�&aOaT}C�[[��ĺ.o,���u����\�KM�/B�ֲ�R-����;��j̜�SI��e^�ޒ���N�����}g�@^��a��M��P�/�j������U�rs����^S�OU�,��i���isW2e��'6|:=�7*��p�f����$tcb��}��'-���br�	o9�)�D�q)}z�G2���}p��|��=����潮�������O�;l���fZ5|��)P1]n��jZ��z
�P�
W:=.x�NPx"W}y��v��~5*�wJ�ٺs�����ou�� Y$���RD��1Z�ҢQ["*�EH�PUb�-���#X��E���Q-F�I[P��FkD�m*�(� �VڣX��V���#
��Y�Q��
���DEdF(*�"�X�KeJ�EU���lm�*�"��b�(��
�PTQU��*�
²�b�Ŋ����"�T������",V1EEb(�jX��(�#-�1��(*��T��X�TAYPV"�#V ����������,*TbE�# �J�(�Y-,EDX�ADb(�TQ`��@Q1�5����H���bZQ�EEX���+F)iEb)QeEV�0DE���*�FEV�"�*���@�Ub*"��D�QX�����QEQQ��X��
�PX1m��0b#APTX�j���R�*�H���,Q@T`������UDb��D��Q���V"ł�bD(�(� ��F"���UT@DQb��j,�m����QX��~�Uv�UӰܝ�q'��|�~/���a-��ev��}xf=�˾�n�*
��g���t����g��vκ������6\��و(D:zg)�z@sc��go�u�}�cuV/���	��z�ޙ���j3M�[]1��I
`���� �
Xx�)b��9�����%\i(b$µ��MNE�~T�6�@��s'�A�!Q��茛���A]n��x\�y��h��$�(>�J�d.b��P�v���{T,d�1�R�F6g�L��S�c&��x�u����}��:��^�H|�o�u������ƀ^v�KhЌx���O���>�$���]\���x#�o��|��̗�O)AɊ���#�b NlFy����ո�[b�D�Yf.5w8����T:�lGF�����������������nz�����dC�g�{�C��'��X�	^TR_�AJ����b����T�7�[�9<|:bx��O�t�Ž<I�[��l�`-ic��8"�G��@�S���b���WO�/y^c��׏�Y��s�(s}Ns|gN�O]�ɕכ�i��t����A�,���(}�d��}��{.��(�3o���e�5�1���v{
e.(�:��OP�P�J������Z��c��>���[��`s��7.�y�����WQ�tMp�s�r��{��J�H��2��%�V,a�f([���uܷn��μYq�y$�sQzH+LZ�7�r�#��<��j�!�N����>��8=s
��v���b�i}��oJ	�7U|��Jk�wu���fz8FA�P�`(��Ԃc����خ�������Z��0̷{1Yׯ��eC�,��T(�1�GX���w��j�G��j�Xސ���yV�}]I�%J��]u��10�|GP��xY��3�\�U#/���[����9O���vm+._Qwg۽��J�u���!0��L��GM��"szl>vL��4����{U�)1�8M�K��ڻ7�6t�)�c�U���ԋR:^����茕�b(�no*aLUsЈ��nRŭ(�h䎆Ml.��������w5H�*��I��T-!X�xl�,�k91,�/��5�+w�h���ӪLl
\NC�Z��5��!9�����[���]3��nWb&�71$���fK^�~5@��B�c�s���D�ޚt7gD^:���|�^��]��ou.ZcJ%0��{Hb�R��k�O_=�O��P��1��i�v7u�ɞ�3��hUAtqR[�E��9j��X2@�zu�&HP�:�*����yK[�͸8����4��a΃3��&L��h&��ٲ�9�b�+����Gx�Ź���ErpY�k��N����IլR(�z�v��R��c��VM�2�ٸmn��}�Q[]�!�.;S~.�%�<�m�C�&����i�oԺ�ꈦ�΅e�F�oAד�^��b}<��ڀ`��+�4l5�bc�D�nj.]�PD8*D�t�vnE���ԻM���p�d��z�p{�0{��A��|�Y��֪ѕ�����.l˷z��Kl�|Nl��F@p�wK=\��gׁ�^}���{a���˞9s��{��Ė����2�H�>�렄8�*C�|�yqw�;�"�E<�������(;��\�.���5;J�����>��aE�0����N�
n�����׹3�3N9l|�J������AX��`6*�l3@��Y��وV6�Y;ӯK�LFv4�ҵ�B��a�����%5����`�&گM�phY�+M�3�hp9��aj�Y� l?f״�&���2V˂tӷ����z��g?�˶P+T'��k����Ve��Ջ�}�-`�U��\�-ҋr��T�3X�XN� q��aJ~�-�BrY9��*����ܴ��,�AzD�ZK�߹�7�o\>5�'e�O{�{i�����\(�{�G �R���On��M��I,����9�(P͕;��^-}���8Ԯ33�IܮDć4�Eo��]�(�N7Avo+��裶�Ŏ:�,1�e�����u�«�TS�l(4���,5}�mW��+��x���Ty�<�4�łYn��t�1vDs� aC�xx���]�-����Y��GP꼩���VR��Pi�=ğF^dPkO����>0�'O�xa[��q�
��U2\=��~܄���̢	>���k�>���+�֘/��s���Yg�Ā�u*9M��=�IE��uj�j����]��E��2��Rã 4��M)q!RyS�XB&+=9Z_8�vg-�y��{1��+3U��}���g��(<��<�P�89H�4z�L:W�Ҩ5��[�r�]-:�׏�(�-͍P�B�,���8�}�4�w9Wbd��*y\rc̓J�m������M�>�<��Z����l^;>����r�w�Fӯ7�4{���v�x�-�\��cgĳ�慙�$Ò�q�_\��m��cՒa7�U��UX+�z��
SQ+9�@I�z�2�{(���Ki�}�8��#�{�M��ݯy���F]Pu���J��t_����.��s�u8�௽����2��rQ�J�S�0V�%�V##7Y*;��O��w�]%��WGp�:7��!��!���^LUHê���Qî��q���tWn�Ē3l}���mv]f��)S��8���%�l����8��Ğ�d�� �<u������������]�+�7}|�y���:�B��H@ "��UA��c}5���+��Hd���=���L�X�\�*F�����:���j���b�R�Y�'a��=�UP؞��D��G�W9Ub���h�@��:�yCX��&Te@�PE��*R��g����ȷ7�\r)mm�b˛:µ~����~�b���yY��L�|@Mz`�L=���cu{W��v2)�72i�.�MsY��&]J昝�9{���/�}4����@ϩa�D{q�^��H ��ʅ�{"����hu!s�>��X/�>7�C��mPs�U|u�:NVj.������w%tn�#�1��Ϫ�vǽ+|Y���z����Z-A���v�s�ϒ�{�aXߋ���ֱp4��d	��;�ai���/I`��LhЌx��2x�D��a�T�\�;����c�&�2(ޗѲnLT�~�H�X�	�=��/5�I|��{v�r��b}s��p��,��t�V���m1-l�����O �7��������B����f��D7�[}1�K��eoT��Z;L��f.�Tʍw=֐ɷ֎F^v��;y�_:RA|H�RNu����y�J���f�wlXP>hxف6.�\tn��g+k�J��A1�lo0Tmh��k��n9m�r�{�V�+��)	>�<`I�5���9�vT�-��� Ǧ	�ۭRҢ�%��LG?uӰu�5��Rc�z��ڗS��B�"�����]W6�OA�O���R�_���b���wS��=r�3=Β�=���h:C�b�mS��Bm8fT�+'��ݑ���;KX|��>ު����ೆ��bN�bK`�sU�f�C����Aˈ��|�_+ޞ���f憟OC��a΍��D5!N225�Z����(획��H�Ai7rܾ~�r�����s!EA�dqA��R���Z�v��N9�#$+��v7�1���%[yS��q0GX�����Ҏ
oMyU��R���nt��S
�IK'�n�M�m*�↰˽�`9����%��E�")UtX4��5� �a槩�����e;��ZX}�,z�u�[��>�{`uN6���!�/�c��.|M���	�Ƥy{�����}�-{U���7W�K7�]�':���w0�:Ü|�Y�ֈD��*LƎ�}��W{�#��a����K4#��gst�2,�)L�F��\!��:�آհ+����tɮY�.f�A��s���ՙ��*f�G:[��;:�12�+diF�R,�]˰��fZ[Tw���y������ԙ���ҧ2�xmx*��d+�f��,f-y�<��N�J��f͢o����7��TV:�Y��zg����=���ۻ}7���Qy7=����EC��Pf��N,)�#�4m8�CL�\��`nΈ�;NޜK�]��I>��bC��iD����!�>����řW��Z�u��E��g1�߉��\���f��s��_o�0��y�K��(ۖ��UqP����*M�;��B-V����ž�ܫ"/z��b*�����j�05=��U|�&��X������l˯3�sms�:���bMnO7,�b�k6���!W��q�p�MT��S��<��3$�NW4�V#�9ȹ�$�=\��Rf�B>�	��܂�g�a�[��'��l̇�6��ngZF��sYf)3�6����]Ϯ
c���_�<K<��
��6\�+[�:h�|��6����f��/��m.ǔ���+ރ��0� ��� ���k�3�z�>紅�N�u���>�W:h��딶��z��%^�-
����� ү�O��v�/{�S�8Y3Z�I�ӏM��*���#�ɧ�׃����YI\&��r۴��C�7��Y3�,2�
���2V�}1lu���rԪ��(����^��9ثٱN����=���6وV�
$CL�Z_�f7�����v�Zcԏo��v�ܙ��S�q:	��zl���h]��.�,]6��C�xG�Ϲ�����Z t���n�,d���1ѕ�~�J$����
��"�^���Qܺ�v�Y��#�*��9͛R�F6�"�An������z�冺��=���sWd��v;�9�э�9�C$���z��`TS�]�GF�ɝ���Tߛ�bX|{��cr������ŶQ��G¼2��q,j��'�r�1x�!���~#�;��(��L���u��m{w�;��p_�~3���]�C[��ظ�a_��utu�Y�����VU8���7g{R�1�U��s#j�M����eU�������yu�ߜ罈/{�ܸ�iO�]��!Wૠ�U'!��:0�zXj���P���;εaѥ��&j�譱; ��t��u-Y�E1�
�����=�6���=EZ&{�?t�|&�N/�/�
W4+Mod��v-�VO<��ݎ����wqw>c�;�|�o6��=]LD�cp��w�E���V(��^�����2m�=up1֙ml5.>6���tqɹ>�f�[�����SV��3���E�]�e�#9��׬n=}�w4�Hx͓��4��Q�[�&���,EAI�ٰ�"�
l�kb�<���%�r#b<��<������o���[���cv#�b����<l��5�D�7��5�:h��d�}Q^EmI�ط`I�%��߽bg�#3r{��2�Z��SV/?{�&\��3�n��j��s/���
�fk԰�a���l�X�Ϋ}�[зz��&��+o���~�{ ��(���Xw��'g{�����dq�p̓�a9���>Fc�9kk����1�Z!d�C���EE�TN�6�T�Ԣ`�##>^���^L5I:c9��!�ܔnk`�T)���t���r�-J���Q3���A�����ۨ::BLk���c��ttn�����GحL��"��ʝճk-Vmmr��v����+��.	����`��@��=�Gaeչ������ދ��d���'8�Zz�}S���ϝ�g~�?X/
,^��~���>�NR|h𥇌�=���뉑5\���h�=c1�|&���PH��V�����v����49X�&i7t|Ep��⯾#�1Ұ��Bw���)��˻+���=�W.AZpELfF�ݒ�\]���{����k��Nv�d� j>;} ����$&���I�����i�U��y�cm�\��R��P�Ob¿mr�P$An���?R��Tt��u�7E�o�C���	��w>�s��+�[	I��NFCB�ێ���P��<}J�H>�ڑҢ��Z��TÄ�s����j�|�u�$��T�g�T����.!�X�3�1`�q�D��x���ϒ˸���n�:�.v��D^�:6���-��O� �؂�R���&R��a/ja@���LM���ѹ~�,重iy�+X����W����t�1n�-۵g"�l9�c&ß\Dך����5�����eA�m�\6.^���y�X��U�GG�D'�N���c��q@ԑ#�A�v����P�ȡv���Bt`+z�O{^�۔�Q� ��sg`�S�7592|�:�`.y�3��;8:��v�����V/�f}Q�"Zxx��PUg���9���I�\§�%���	�4�cjѿVn��lx�ԅ|Ց���pF*�;D-�!�*�cc<ݝ����7���j�`��|#�jB��;��Ѻ5i^�j�i�?F���7�U������]wrQ`��v�9r�x!���W�O�̛N�d�J������o�k9
���g�,꼎Į��d�No1�E,�F����٧shk�crgSZsy�˜��Q����-NJ�R�:�b�$��e2�df>�5��W�v
-h̚w��uG0p\�e;�E���򤔭�l���][����>ݭr:]-��ٰyݻ(���d�}׹1,��`	��cmQ�q+���tht�zH���Yԡ��r݉�ؙ)ᣣiX�����qI��Ύ �9�Z������ͦ�������9˶��s�ia����\��s�-�R�9�yov�@����޾V��)q�G��KO���Kg=���V��nt�{)�@�x-������>��������r����s�v�,ˮ@l���f�V���b&����z%�>��̼����8�M�ٮ����9cN�\�l��u��t�K�4Z��V�lRYAed�,�Q^h��8�AͲ:Ы[Ne�;�Q�{Ui8:��S�����Ri"�l��i�J�rk���w���{�C��b�7�P��燪��1�Q��tViC�Y��5��m@rB_gt���2����o*�<>|���XJ�s����g7#�c��*.w�qu��y�Ek��W�@-����¢��,��Z�Pqu��n��(AVO�k�b�t��U%�rL�Ԏ�}9���s�e�4��d��]�&�n�Vԙ�c��kc��o��zU�a	����#����vӗZV��nt�o�]��p#7-��wM�vΆ#}�:���1fG��ތ'�73%��k��R��g,�zL��4�hI+��6���х�T�����pr
��dt��b�[w|�ѹ�_���焙��P�����g��RJ�Z�ވO0�/)�J�v��XNܚ2�>[�L�Wt��1��\���Ӡ�2�Xk�u*��pF���7�z*��t莃9�v�p����un�s�Ŝ�V������<��a�t��Be�/T��OGLvы僷|��n1���+��ٷ��H���<&��B�ao;�{��r^�m�Ǥ�~��T���8!̓����;q�M��B��SUt�+q�]�=��Ӄ&�:=GEa���Yވ�K�/gʮ�-�VS�}����1����/6e�lM=��]u�7J�����|w���5S�c0�W�T홍�uڻޔ�����)�-���ևJ��S,!�����3��b<������o�9�D;1�c3kX,Xs1͙�������d����Ҳ��V(���f=�κ�����4{�Z� P�"Ou�\t����ꄌ������+7iI�a�:J	��kmV�蒼�v���v`�@��fi�SU�X�*�J�I�.���A[�y��r�puc��b�����Zt���ß5{F����e�-����mn�H�?A?/��Q��"�`�+l�EUA
*�b)YATF"*�Q�J��
��*+Q"����cDUQQPX**1F1H��AQ���QDdE��("�
$E�0TDQDFTQF�UR�"�"E�Z,VF,�Q�l��ҫR�DX �F1PH��(�Pa(�Qb�UDb1b����(�TUTA�UXʖQQ����kQEFڌ�b���"��eE��lb��QPQ(+EV(#AA��*DF#X��F$DE�QQPDEUEcQ�X"��KFՈ+�bZKQ�mTQb
��(�,1UA���E�1Q�lPT���(�Q�`����1`�b�X��EEEEDAE���ڪ���b(�Z�+��2(�X���EH���0DQEPAFTX�E��#�����c��0V�1b��A��!�|+f$M��ZʾXRu���ɇ����9��`������Yzwu?:��kbik���u:���H�'+�ٮ���cr�Q�E���!�"]�b�Ţ���P`��b�(2:
tf�=c��=����YwWU	�6u�J����_�W@�L�Lp>!P��XY��y�ς���\ߖlb@��9���%+x���II�w�����Ba�{��C�rcR��=<��F���Z���\ Ǜ3�8��t��\��h�O�ܤ뮎�Nf;u��T�jE��z�-���*#g�^l��u�n ���07�����/��Cj�ت�uJ�sQiQ�]��I^f2lo\���\ެN(F�=�٣>bZF�~]K�_	,�y��3�[U��(X�~h)ԛ��(�e��o��u�N�0�lŖ�e�|�
.�z��b���	��2����\�8Or��f�8!���D�.LERA�P�w Y�QQb�	��6b�o���w�|��vR�F@bKe��,w��	�	-p9�r���E��/P9EI<8��}��vX�{5�ʝ`[%�:�K�`u�~��sF�S��)x=#>(�U�Edw�_D�o���ϜxZA���ݕ�C��rf������qw����f�����6nq|�6c�����@hħ�}����>���x�N��pb��o�y�b����<�]�KjC�+\S�e���cS:���V>yY�j��"�ʧ����o3�{/�$� p�B|-3ܫ-�µ�ֳX� ���I|*`��<�=��.�<��K�*+��KP+�V���mT�Y��RxA�,�|��U�s��d�����S�3�6�=]c�1���1�;y��s�S�/Ӂ�A���~pWy�<�ܼഎi�T���s�*A�8W������>ٶ��^�t\`\��(-a���nҗ�{-�Ӎ9����x���P�3�t8�rreȨ��z+�Ml[u��pѪ�f��r�n��{�xb��ɿ;G���ⱼ��"��=J!�o0����mժ����sN����?$�� <�Ol^�l�6���uW�Mۅ���^zf:2���(��!W�@N<�O/��މ0T4�-�Z"rLC�}^=P����R�Q�����Ct��r�g�a���r���4��Y-�H�-��� ����q�+f�*l�*)�:��_���v��pB�M�C]�t}�6^;G���p�O/0(�+�<k�鼬 ���W�|M��Esy�����7�9(d�a	q���WV�$�L�D�U�cs�!yF�QU�:���>V�u#�燆�n��ű�λn�����
0�%���,�;�q�`��wS!�Y�E�6%�j��_�	�Y���6��koO��z�׼�&��Hǥ��J9�/���xѸ�a���N!��t]Z?��u꠼=��*����%J�.wv�$o��gT�;��}\�i���'`��EF�<�"2j�A��7��i<Ҽt�/:_����2����U7!�5 cLੲ�ă�@�>N��`U��E�F/R���s8gk8���9LMR��9P?(l��EW���D��Z�Z���yX��v	��nE�q5����e�gW���
8KscD�! ;ň�)3lF����38ݝ�"8�`��u�k��8�����]�;9w�Y��O��8����4__�xb��ξ��o�h��U4X�c$�}Q^z+jHf�ż'm��j�-��E�Ϳ����v�n��lh���q2�@PW���<vͫ�2�ݔ@/����f�a�À�TQl�����WKf1_3�ϺtB��@5Tc{��;��qQ��=���=�0���xv�7���˿�Κ�j���W��R�s�,@�QQj�<��m�X����"��=��e��������%5m:�Q�~�9�E�(�t:ř�z����FT��t�9ڠ8;�K9d7:�*�^+;--N��٦pRi�Vl�v�T�:�љJh�o�������q�Nz��9�W�����)
�gh]\���:�n�VN�l62�ڽM�p'}]��4�����X4�]'��aϷB�cY�;u�����;6{#b����Me�������A�F��g��p:0��E�d���k�b�29[�E���g`�����`*Ӆ���>/��C���-�3��\@��װG�����<�Dޜq��ټ�N��V��B�Fǵ���R���Rz&������}_>�NR|h)a��)�4��m�V�8/z>��۴��.p�q�ߧ;��h;�jT	�ә#�F!1�!��Xe���㙹��{�=��Q�)߾F��b�P�t)]���{T/�.x��(�ؠ�b8a�٬��ݦ�Ff6�bC�L^�|��Vy`�����ף�X�ܸ�Ub1�v���T��WY��7���?x(ɳ�,��m:�@ଞ?L�h��V�2}�x�̬J�š/\��7=;�ݥ�.}��>1:r�L^e�A����ӹ�1{�J:knu�,�5��y���
�~��d߹}D���ǎ��^�>��Y��N1f��4�+jވ��(";L�xYon��|���'0{ W}�M޻�o�B�Ӳ鼃h-���ٝ�Rw�pV������,~�6᫩-���|dK@��ǯ3\��n�����]��1�7��"}�v�}<q���ŀ�X0�v�0۞�~��|K���I�sWj������#f!P�`�E�����~T=�c^k���6M�g��5����{Rզ���Uf���1e�����v����ʴ��:K>����"��*�=c]NI�*��Ɩ�^Ȩ~,ɅӐ}f������Q��C�茍�}Cfh��bev�a�}�9Ö4ε�%F��6!|���Ցғ ^<�|ϖ���Uc��Jg:�o%V�%8���\��MnE&����ؿŝ��{u�T7>�(:����͠y�؁mN�E��F��mL�l{��mJ������#�"z�h,�h���syT��s�[�Ʀ�(j����������!�Ұ�]��r;$%:gCa��@�KMo��\4��o!�;����՟�)�?<��ߟd�}�.J^ػ<�`���X�A��*U����3F���޹ZN/4!,N�ʭW!ƾ��������uJ�sQiQ�Ne���������}ؾ�.�9k�irA�a~Y��``��#�}cY9Rj(M:�����N�ދ�m���>��T/�\#�P�s��6����d-�bR�ݺT%�{�t⡘Jώ4;v���x\�ۗ�P��ܹU�ѣNB�[C��sYnsY���2�V��]�Rp��ܳ.�vfaj��q�خ5��� h�h���{Mj���o�'����6be�4<����DŘ��ֳ�׬aΉY�wz�Q�2�c��"x�m�w�!G���,����g>���5BB��wz��4{�:>�v`��5�z��K�ޘKU<�%�<�l䅞���ϳ��ב�H�w�]Է$�[r�uDSt�"yP	z1s~j�0T��t��&+f���9�8��V;�U��>�����A������F���1��%��
>�[��4bV�a�ƽ@����G�-ƻ����b�����*7�({�Y�_և���n�=C�~~N����tT�w�e��'�zl�W;�~V�)��"��Z�i�>�t��B�
!�9_�&4a3������g&U���^ȥ�bs͘��|(Ԑl�R�xd�z�h
���DV2t:	�ܼ����7�yf���G��u�k��P�f��b���6�M0����2�#��Nq'���sv"�@�2�
�kf�_���]���ǩx�#y�����`ôԊR�n����ϻ��\�����C��k=�!�W}�j�Vu>�Ok8�.ȝ�Y�y�P�9�ẵ|Nǝ375Gw��v6�OVͫY�\�p*��Ȁ���<� t��v�P����������ɖ�3šP��|G�έ5�\A�U��S�{,��5|:7�4��Z����BA���7n �[.":.���(��unq9����5�2u���P#<������$Z>���86mH:���29�Qn\�ʗQ{|3�b���qwxӷ]8�u��W�P����9���V�"Tلe���w�>���Bs�2%�F�f���Kv�����q$K���ڋ�ڥ���>������gD���M�X��	��u�Qh,Z�X=9s�9�ʛč���1��B#eUh�* {*%7ד>�r�Y�<4�+�ǵЭQ���������֩�Ћ#1�}I^[ʷjФ�`4�.c��o>|�8|��@�e�	�_k�'��yQ� ��
��T�A�
�ױ�[�7��G=����qc`W^�dg��k�ʁ�|�'��J���=EZ'�P.�]�}v�_GG%Ed��-'c��(�sG�����^��
�%���j"@r7�Q�cl�V7n9�6�+V�[]q�܉�Fx$E{���I��^���}C��9A���篫I̎���%q�4nV������E�d��rQf9�Z��[亗9�G�y�N%�;���=���~=ڙ�K�4���W��q�
}�i�ˋ����x�p{oqGU�ͻ#V8P���!���r���Q��t�݃*������zz�gk<���G�.�y>�ɢ�+��DTS�[RC46-�;�J2.�#\Kj���3jD����x����;���=P��̴��))�W?�K����'j��*(�՛8�s�JO�q7��k�m�k���@#�M������Μ�J��|�Ҷ���/�h]�m݈��r���\���o�o��3��p����7��TZ�'ch�J�>*&fo���8�k�����:XB���1s�B�d�F��T9�)�/���v���ъjM���ws�O����dJom:��ƾ,m��'J?���/��%�6^}��#e!l���ۻ˜�7��F���sa��X��)�
\XdWV��E. W�^����ګ��|�r�[��j�׭,Wӯ4��8���LrT�i���7�/���z���r��@�~�r��Y6���ݖ.Y�0?U
v�x�v��;4��A܃j�	Ct�H��Pq
��P+�����۹���%���[��"�GPPp�Bs�#`�6z�ێ�ٽ���>|P�6=a�E4{v�o��K�l���]禄���U��V����x(Nw5��ľ��'�Ǡ���7.�p�\�kLJ�Y��],�"����l.�����l��ΔH[Pn9�[�^w[�^�s ��<f�;��ox1_v!I3E��yn�S����e�}I�ZG
�g\_�b�k��k�Ɉ��2�[�>��n\l�pB�tެ���[*��{�Mc���~k̞;�%�oћLV�VO��1�3�E�{^�Q�D�;�e���A
���p���P040������_��0_Z�lm;����9fb;7m�+\��F h`Ѕ:ا%37�>������-
7�5�q�h��B1�w�,����;��꽸/ʊ�ӐcǦ!vK �E���ETz��ڒ5�-d��wb�e�LM�A+�_�r߶�c�sh�@ۦ�,��+�8���MA���=���n��A��B�g�{���<��f����VeG��><����UYv��������S���9�K1w�G�ˡ��U���m����!-]s��>�FF)�;�B!Ԋ>(n�|Н�[uxsEa�Z�]Zࡷgb�_�����l��W��d{݆��\�Q����J��� ��
���λH?P��C�"<�T{Δ�`��S�ߕg+�����|����QH)��=�:�C��Ùa�Y+b~g�{���&!^�G�M (��5��I��I�M�A�0���y5t��w/��� c�=�>�?R���G�=l��R��_K7��љA�ܴr_8�{��d�/�ד��E9;����ܖQ��i�[��X�A��}���B���^px��Ig%����B������5�J,�����˹XtU4�{V��/��M�4wfZ6�7x������{����Rz����y����?���I�?e�����6ùM��!�)�O{��$��O�E>d���<��h�����H}l<��)�qRT��?}��FH�;1w�R�~��{���;!���m�?}�m��*O>��'�gRz��u��׈I�>O&s!�2��>M��ɷ�OS��;��J�ɬ��Nf ��a�y�0<!Ͻ?h_w��]���bw����{��{�>T*C��7�k+?!�����M�!��C<i�Xq�"�0�����S��6���ɯ������y��βy�����q�q�x�@L����N��|s߾���c<d��;�b��S�����H<��s ��?&0�V� �l7y���
�Cg��l:�C�ug�Y3���fӎ��C�I������}�@�4}�TͳE���,��<~Oڠb��>Cm��7��m�T1�������%Om_�
�O�T�IP�Y4�ɮR��<�։��AOʓ�:��F�������؏kZ�:�+3��{Ny߾zx�|�~L��9��ć-���C��?*J��{��d��16g0�:�d�[s�Y4Ì*w
��Om�eA@QM�y�si�
�HTfϽ��xLןol|*dዬW��kό����z���_�5���a? Q53�+6�ya��C���P��;�ֲ�Hg���4��+��
����z��a�E�C٥�$��>F���ߵ?�G�������^�������1E�{�ӷ��o��~d�}�>'�L+
�2s����1�������j�8�r�&��,�ć�y����Lf��$���'�~(��A ~�����<�~u���~��|�S�3�>C��3�%b�y��6�դ���}�b�=��L*w�|�a�a��S��&�V�G?d+4�g{�AAE����X�#_
�D�9�&��|�;����}�,�)
�����u���5�O�|�O�Qg��bx��<��T��z��w��ݿ[&�����G��'YS���P�O��O�5���&0�
�'9�^?���������� ]�>��@%7�Vk�//j����^��ԝ:��lO��iMU�J�H���k9�i�M���!�9X^ֹ��]��K�Y�ۻ�;ri�h�=���C)&����r:����X,$�/rl7d{�ҋX��'}}e�^C�z�m�R�lq�$w&�ƷV�V0�)j�5�۝�٬��Γ[�ಳ^�x&�N��f���*��k�VffJT��)5��g�;��ύrak��P��
�N(�4�:����v �G���TZ��N0j�Njps���F*f���pb�i��|����+�����WS��fh���31�U����4��4`�k�#k��xd��wpa��xs�Ҵ��=;^���7�f�����I��˘)s5-�n�R�F�P�V��̴��H֖�ei㒯Vbv�k$v�6��T��XgL�dy*_�S��B�.n�Z�)��}��m�1ۥ��M\ų\޾�l8�^��E��qJ�wu�1�p�Ob�٨w�Y��eZ���D��7-g��{��Ӯ�%S^�]�C��o;�BYA��I�YYow��ޞ�fe��l��>D�C��,C�\�T�Qk�@���Fw\,AZIj��ܖU�Ss��{���zw4�m����k��r�f>V��Eb1�È��A��|#����F������Q)��'Hp�muuZu�P���:7Fp�X�����gL�wN���&fqf�bw�	\��i��VQ��D��Y7�v��>;�j�W>�ǰ>�8ON2S�1�[�����63kQ��Ep�[s1V�S����o�<�k\T�iV���J����>���Ԯ٧���2RlΙ��c��	�t`�t��[��U�ۊ�:��T��=�W���k���t;	#�wX�8,�tq��6�^w��52k�ߒ|��Z�y���"���9�]��3r0�K��U�ن�p�Je�=�[w����ټu�-��sq�T�`�E�oqN|"�z[r�s�M�|�=mw�/H޺"�*�W�!���j����5Ǚ��8o����!�ӨG�.M�;-�c)n: �:�l����A��j�_-�
e�Z�����n>�U�.����+��jw_Yrk����(�V�٩�n�k���3�W(��7��K�VuqB��F����6�dW���Wv�P?j��͈��B��9$M_v�4��S���plmMکi�n�;u�oQ��&�x��h�bU�V/p>}�S�m:+΍oG�'��{�*�d-[^;Lp�ӫ{�ܝJ�,�ң�a��V�k��<�l���1J@oVnS�}eb�u�)�J��C����`��	���8s{�����9��v�P�`c��Kuo���f�R� xW���맷�,�of�b���6�7'`�gm�y�no5��EH�Ț��@AF���T[ZDh�%�Ub""Eb�� ���"*��Ub ���AAUEQ��������ȥ�UQ"1U*��QUj��+AE��b%B�F"��b�"�kJ�(*"��ZU��(��1AaZ�m��"��(*��(���VahX��X�TT��+R��R��[Jرb"�+��ŃTb"��U����YQ�UVҪ(��RV��,b4lQEQF1����DTIZ�j�cAEUR҃l�EAD����1��A�#UQ%K�QUQQUDUX*�X��PTjU+U"�� �UAUV"��EX�ZTQX�P���Q�,
����Pb�,Q��E��+Z�*��QT`���EV*1"-��1U+*���1F1X ��b�(*�"��-J��[j���T`���b
!YUQ(����
��_� ��$�H&l����*w����/���*��ϯ1�;�U���5�ƥ�1��4Լ���-zt��e�����-I.�xtj���{���vu�N&���!���[4�C�a6����ݢ�1�����z+'�j���w'�6���wV��1�2W�&��z���y�'� �g��N�Ê�I��7l�Ǧ=��G�}qB+.")}��U�~Kf�|�����N~ͳ�<OP��!��a,?0�Y�g}��C�Cw�MO1E=��)4��!�\��6ϙ=��f0�³L���|��d���xM*���\��?{��S��ׇu�s�߾�����������@��3��z�ϓR�Ag��q6��TR}ϰ4�0��CI�{������(��i!���C�l��;LE��T�VN��|�a���������_���ĸ�)�ݥS�����`�;�{�f<��O�i���&��(ŕ�֤xLx`Z|��:���,�N8�IQ�w��i>d����x�H?Ro��M���`}��}���e����:��ǟ����@�+?*J�%E��T�:y�M$��g�ɫgY1��y��'m!�����&�S��;����I�ӻɴ�'�;H{��>a__x��>�'^�8��* ��j���n}=���>QH)�N��'U� ��k�����j�����9CH
,a�f���1:�P�����,8�M��a������d���L@]�����?�����e�B���o��os�CH|�5�d;���8³��r?y�u�ûފ����̲)�<q����R����6����)�&���E�M�16Ì�?'=���_|�/���܏�]g��k�?a���ϲCl�VLC�����
����6��V��w-��Xq�M��I�v�+8����

/���)�
�H?fI����g��x�}r<�R=�rP�����&;+���O���1'�q/M�8���wOP��<�����{��iY�a��sh
,��4��I��B��̋-��&0�lי6���.�>q�L "@F;���i�X6{�a���g߽�I��a��P����9@��i��+�'��{�c>d�S;a�������+*<��!�XiP���@��k+���Ch
)5�#G�?F?�>������!}���G%n�p��H����3bte-�'b�LO��z�¯^˥ux�BKt�	�s�7�c��ȇ�Vlr��vS��y)�'b}@e�}rT��nV�w�O���ڤ��Yr�LV��J����6�hڋ�8 �!�ä��!F���ۻ�������~a���2x¤7hlϰ�'̘��j�����o��*�d�w�a�
ͦe�{�AgX=�&�UT�߰���i�w|�5�B���I��=��]�������SIZg�a�xÉ�~B��j�Ĭ<f!��Èm �ɹ�,�q�06�):�f�d���(��;�7���T+&�}�}��Xq����<�X���|�/��������=k�=AAE�;����
����pwd���!_3Xa����ܳ���R~q&��E �2h���� ���&�l;�C�ԎP4��Vlk�@�~�����w��'��Z����=���IRi
���!�n���v�&�m��X��P��5��~q:�Y�k'�6��?9�0�0���yNn�Y�%~��'���SN��hO8����.��VK�wWl����V�*G���Y�I�����:��P���>v���bi��O����YXT��4���O��&0��P���z����O�V~d��sD,xlxL{z#L��%[Z>=������j�q��&�UTC�bm��,�ܰ3�B�g>�Φ�����Vm���i
��$�3}�=Ci�'5�bͦ0�M�OwI�Ƕ��^���ꈯ���z�{T� ���N�}�@m'P�<��!���V���M!ĝ�X�|ɤ^&�o$�x�Rl���<�~e�����a���Ho/�� V~I�!��0SHH�4��=��?]��w�`~��ީ���+��^�6����bxn��Jϟs	�M�&����>Cܲq���LO��|�I:�l6�C������)�OOP/��蜀.�x�9��u�����õ�3�o����0�
���
y��Ϙl��6�O2�Ay��	<VT=�����,8�hbC��7ˌ������N:J�0��<��P�A�é����u���a�}?ek=���ל�*&��J���1�e�"��+��t�r$���g}��0�a�����u�s\�4�IUR{�1>@��l��H?R�������և䕚`P* Q���9��#!A���;�~9��i����+��h��:��+�m�GR�Yq�f�6B̸����yj��Xu����5i^d�<�q9}`�03euq�<��V�uq
���|�p�4�(�et`���k&$�����OOu�\����˛���� �ݒ�n����
~a�y��&!��w!�,�:�y�d>�'�Vk�9l�AaX~�w��:�g��}E��kP�|�ܵ��J��|��H�1�|Y���i��Y��ݯ���;�&�yI�1��{��3�/wH,�N8�fC�T��&��C���VM��5���5��fm!��bT����M$9�+4�"����k�6��zf}��P��"���g���ܾxd{Ǩ,��'��	��~d��@��=d��f�'�=f�}��V�zÌ�d=7�O�J�5�`HT<�U$���8�O/��2��v�^����@d|_� ~jVx�����6�|�����,�
���7���S�����?$��>�)?!Y�k\����
��{��x��Z����bm���_�����K��H=Q�r����wUB�.���Qv�X;�6�>LHr�++�!�}�	���a��&���C��X��1?OhꓨVy�zya���LџaS��bN�|w��
ߨXϷ�;ٿw,���G�� 	�}�a�?$�Z�YAgY*
��4�N Wg��x��,��{C��4°�)<��5H,�Og��i:�H)���~t�x�C~�e�i1�{N�_��{�_w�����ϯ=�Hyh�O7�N�J�X����)+N�*d��٦;�<a�& ۖ��l�%g�k$�z���4�$�<d�=�o��a�ߟd�'<�m�}�Ξ�|�{矽�����߽��=��:O��M�2v~��Q'ʚ�� �C�M���Ci[�]���1��Y����Gy抆!�vl;�E�aXo3!�Cԕ�:��t�ACԕ����_���!w�O�Z������y��z�P����4Ͳw��O�3�J�d����Ĩ8���4ξ$�<s&ޠ����{�T�Ͱ�bn����<~t"=p@0G�[;ӭ�1����k}�{d�Y�|æ�C�I���y�Rm �ߚ�i>�~Og�i��^Q@���i��Z��I�~d�)��`i���;��M��Y4˺{�0��h�q�����<�~��cR��Rz�V}��tgfA6M��o}j�Щ{�#��N�lD���e�l����-@u���g[��M���;�gB���T2��qI��Z�&.7���9�K.e�8��u��	�:2���uaw�a�{lb�m/o�*S����s�>y�g?s����(_i����pZ��QHjg�h�����*xj���6��w�����<�1�T�OOs$�*q������[gY��0<a�
�������?2W]�f��l�߿jj�ws���2	~��D#�s�&�q
��ϻ�w�!X|���͵��֩6]g̘���QC�Rbz�D�w�d�A�Hlι*!��N:egP��Q`q�Y�\�=�¯�x�Y��t�Z
o�6 0@���0���XVt9ܓ�����O���� (�P�<�m|@ğ��{E�z�T?�q���'�5��t1�d�����b�S�Mo�:� �C��׶��n}�MH�n0d����ﮪ��u��ߏ,��a�w{������u3�8�0����X��xw�x���b�yd��?5��I��I�M�A�0���c�>aP�N����=3(v�,|�����\{cޘ&@Q}`T��4�2��U�HVa̧}�甂�'��_~J�'��ȧ̞��x���h�����H}l<9��i�T��h߻����٤����5�s�q�(������'����̓l:¤�����$���u���׈I�>O3����a�l��6���sV��i�d��Me�)�y�~�G{�KP�a{��mwn�O�G��������H*C��s{�Ʋ���Xb,�+7����u@�{L�Ì1q�|݁�P�%z��H
(|�����1'���egY<�a
��o��w��/�/|��>���3�My���L�%La���UH)�sz*?8�yOw ��?&0�V� �l7/0�!QHl��m�Y�~N���yd��JśN>n���N�����{�<���\�4�Y1E�~�����b^��1��]QCf���aP��qݬ
βT߹�����S���M$�o,����)
��^�D�e ��I�ĝJ���K�'n���V��}V;!���
�{���#`|�)�i�5�C���!����!�m��%I��H�zʘ�3�T�B�c-��,�a�>�T��γ��
�xɆ�ͧ*M!SZ��^����J��t�����`#f_��Q�e�ѳ��N��f�Q���J�rׂ���FB��zrf�!�[N�7բ!*}���� ���,w�]�zV�fcPc�9�M�=�՗����^�d�Q=h�t�������;��֖p3�{7sy����B���i�2�{'���
�����&Ӛ�y�c+%xɼ��ل��Dџ`uY���̇wa�P<;�;��YY�3�}�E�Z��s�O�uI� Q��
�� ?�������G�ն�g����������~������M��i��$���g̞g2���f�;�a��Y*i���6��S�7y�I�x�C��j�}Af���{�\��d
��U��@_M�Fvw��ا�z�E���?3�x�=7`g�JŞyN��CV����}�b��a�;�>�=CL6��x}I��C��s�N�k�I6w��_X=��o���n��;�o�/}��������I�e�O��f���6�>�Gt�!̤<��j|��~J�1���<q��fq
�}�y�i�{a����4��T��=��Y:ʝA#�������z�8�������������}��/\��&0�
���:��C-�~�&�R���`�L@�?!��oEd�5�7����ߙ=N��L+>d���y��� |y�	�eH>�l{��q���PϾ�e�~W�7���r���ϓ������w�ٶq�����?w0���b,ӳ��m!塌6w����������)4��!�s��>d�7�zn�0�³l�3�ǄG�{� �?g���u�g���]��AN3��'Y�7=�~�+�:��w�<�Af�}����TRzs�'�?3�|������~�)��=�<;�4�?Y1'��� ���#"��(SM�wU~�����z�a����`a�9I�Z���~�H((�`k�a���e<>�!�7�!Xx=�9�OP��~�gqĚJ�aO�1�};�/&�)���v��;6r�/�x�\�aM���`vwy��<J�ʒ��Ɉ�zʜM����O����5l�&0�'뤜A��֛��4���f�w���
����M�?9�C��!��1��g�ƞ]q�&�7���~��?2W��r;��S�7�`�>VT�۹�d���P��VO�`x�Vo��mE��|�%gbu�����Ì1����?3�Y����2 %	��^��_���*����޼�{X~nU���遧�ܭw}�����:dݶ��!ۦ�<�g?�e�,o=U�)9�W@�zj1lNb�f+䝬�os�~wO��=�_������N��:K�BK�L��je�E�o��>]Q�iL��{���<�KMm����_�ĕ���wXCl�ɬ�d=32��+1�#��Ag?��%UH)��sY"� ��nj�9HW�l��6����)�&���E�M��q��� t�
4��W�}��-K|�ud��y�i��bC�|��!�{�&!�{��Xm�L퇇3&�u
����@�8¦�E'���Y���i�Ne�I�4_�}�K��1�n�����'s>��$X���I�>�N�P�|��q.�R
~d����`i� ��p<O{�I��09��Y�a�w��Jʚ��0Ri'P�n^dYm��1�<���@2<7��ت�]:��^�+�>�d�
)��I��a�S�N9��SL>a_�<Nk���|�^��܇�QH)��Ğ�*��v��,4�W�dn�Ʋ�;�6�"��C���]��Me�ꏯ9%Y�_�Y�O�x�:H6���<̝aR�7��4��d�OTP�%t�~�	P��&�|��>aY���d;��:��{��i*�A�0��d��Y���g��Uj1w}˫�{ߩ
��^`��Z��3�&!�
���񘆷�!���'�b�'c�k��B�|�bxZE§{fϬ6��Xi?}f�E #���<ŭ���@��bS�O+wq��C��Or�gN|�AAE�4~�Ci�
���\�ݓ�/i
�f�6��)=C�g�nɌ�'�o��R
c&��6�x�H:��ɴ�����#�G�~o}���/��gj�>��{ڿ|v(
)�����:���>���������e��41�c���v���E����iwC�
�e=�\0C'���fa��u��-s��"���VԐ��xN����Üo6�Z֭4�uf��u�d�a�)�|�f,FAɨ>j�̾C0s�$�ݻ�ǌo��o�����n�	q�����#zv�A�3��o������]�3{�/n�\QK�v�b�/�H�K9�Z�=��-½���u�x��y�{�]���ɬ�7��B�n�=�371٧9c�>0��;h��s�s��Lv��������<�=���4�-ta�}Q@�=0����D����n7:��wK��l�^�x2����T�p�{T�Ya{_��㇢��Kp�Z1<��|O�j�8T_�Py;Ob�ׇw��
�Ԓ�R�����yP�3y���=�����]Ea�U|G�T)w��u�j������Tv�6�k���XTc��uCbz۵C�8���_N�~�i��4�æ��sn�$�h2����&b���*��+��]��|X��������u�"��4r���;�������7��~��;~H���K�v>"c|�;�x��L���	�p���J�gY1j*��z#��E����K�65˱u���]�!+����~I�HU�gu\�9���Gہ�!>Z��T砡�q���˩��P�uJ��`l���g�%;�C�pkk����~�t���A�_B5q��'�^$u�o& R��N-��7w����n������1OC���l�LT��1
8w���b�E�"��Ǐ�m���;���R��Q����0,�0Xh��&�+�S��xﴽ�ӝ=}�Lis�7�L�ow%���\�˵zʉ+5iW�gN��Ll�1M�#���k���0��i�|�T����B'^��p���<8�Eu )/�m\����\����[�Nu������Z�˕>�[=�xa�%��x�NpAj+"*}�a�)��:7~~,��,�>󾅙��!*���L��8�Q~���S눖�L��835��B���n�<�����'�"�m��{E��Ӑc��1
�)�7�-Ċ�ur���g�Lt��bM	�׻���<��qиȫ�>���7�F�6鹋	�"v���U�`I�/i\�l��kgo��j^`��x!�<���(��ʏ�Z��g׏������]V��6^>ԫ*R���l�,����9m�-[����Rc ^<�|ϖW���{�5#�{)ZP��4.#XBr��cc��]���J�\�6do�F��<�1�|�צc�=�4�R0߹�f���͠]��G���8�W@���`��H�u��n���'o_�t�7�=]�%�:g�Ƕ5�(����.N$�,�{��m��PԳ�4��:���&��R�{|�X 5T�X�Y}h�B��y��5=;K�����m��^6��C��wd�蕙�F��b�<�j�%�z���q>YU.c�MsU��{�)�m��G�HWm�R��^}\�5M��\���.�)���ڥB�2ld�8�N����n�w3[�.�k&�����d��T��/0,�Xxo����\hL�������2�z���+�:����`T�^<[��M�
,Y�>�X��%��-�#�<ow��]���~��O��ߊ�c�w[C��F*��zF�9�=�s�
=J�8I�)3�ũVC�O1}|�47�,{�:qS��h=f'���缆�(	��2-���p&��M�~�ސ���&�;�l��~b�q�D��	��ϩZ��\�Y�z��EC[�Ŏ�U��3$t��@O0B�	�m3�6�(F���
��w��~5�]x�v��%j�0�B���T��epꈦ���Ur  ����Ѱ���nq�dI����wس{{�d�bx�Qx��4E���3��%�[�ܣ_����)(<ƽ�p�?n��tgq-j����(ԟs0K@�Oua�Z�R�.T��,�.����J/+FG���d�������.�/��_MA��b�h�+ρ���5�|{Tte�z��!#�8�d�Б�!>�wբQyߜ��l�{"�Q�n����]�iL<3K���U��P�0�ݧF	�u��4rl�'�z���m�vz�rb��`v��fm��S�\���S)�o6�.j��Dq{ۜ�闔dE���c�&��N0eU؂ݑ���˫Ok��w6��O�]`���u��NSa����}_ =���I��&ȸ�M�ehs����FG{{��꽚�G���g"�b�g0[Pj�)K��K�z�m���d��;3��ʮ�X�`5�f��L)Ԕ�k�R]St��������K�7����'��z
OL��-�m!j�2v�g�+e�3�ԇ!�VK��Q�GFFR���-`>�{�+��=tL�O���/y^*�3�9���<�A��$�۩\���kiE�r�*Z�������Ә�j|��i��/�L�>��{��?w,�YR��.g*l7@ĵ�tK���ڈZ)�0�!ET�F��K�b���H¨賔�_�{��@ݞR�v"n��FⅆϢ(c�z���c�0�V�3�.1�ё�LCUpl�тqK�utu�1�����������y���s���#���_z���yH�/M�y`?Y}.�/���U7!ߡр0=�Rd���w�Y^������	o��O򚬄LY��E�T��\7���dq�� ��K����,�j��f y��������Z.���;R��c�=\W�Dl84�>��`�u>� �rT�JNJǩ�Y*����:��!����<_43Zh�X�S�4��J�򛺖��gR���nvF,�;��\��M���e֍Y\�YX�AL��ו��;��o���3d�L�r^��gC�{y뜲�f��pʜQ"Z�r'�zK��O�d�[�-X+�4��3�35���Љ�	��Sb؎�F� [��=�昭0��%n�Ksm�͎��G��h�{�a���4�u��]�g&Y��Oo-��්VL-3]�hZ�<!������tC����x�����%|�pQ
�a�x�� ���Ke	�E}o8����[�
xl�ǧu}���X�"���#v4�.��T�s|"g�^�p����dy�q��s;07h��.N�+�aOl��Pko�|L�H4m�i���ۗ|��}�Ю�v\�^.�Yx�w�1��b�:'(Vd=��S�&\�����[/%���m-��X�r���c�v��ݷ�\;��5�WZ)��93YUv�u�3q^
�e�׽�oV%P�{/��6��M_b;�"ls�]Z��sY&�^�|�Y}b-���iY\�A'G�]8̘/���oͽ]6E�����`8���NnS{�k�\b,��(�cr�FIJ措�s;y��҆����I��а>��s�@�๖�AK��ܷӠ��fI�,ݓz�nv�N�V��:)k^�<�YbN)vC���ܼ�{�͔�v=�m���,�7&����YH���`,.�`xޘ�r,3y�A�.�� {��G�)�f��񜱃��c�;f���\A�y�fHA�V{�����&[�f��LkםS���v�KΗ�����DP���[f�"��wS�*I���Jcj[.�p�#M7�����j���.�=}n�3e�UR�F\ʲ:�B���t���}]�/��.�D.�3�Nv���M�~����6��3=t��d0F-H���9�J�L�t�	89�HЂո�:rm0����g��f��+0s����;��AU��tfK�@�{A��9c#a!(bi*�e+�zLw/I3vv?��K�y{��u�r���б�s&��\���8jm�1��pR�_,l�P�Rc�];�{�8�2�b��`�@�s���]��̰�h��7���,��Q��3�ޠ��<��3.SDWRu���ib{��Df1�)We�#Ob�ʦ�V���5�z�]���U,�k�R�N���Gt%�V&v������I��My���1��;�hյ�lOH�������]%��!e�0�-ഞ�b���@'v'J��Y�:{����i����f!��\���ra��|�JV�N��[�U�v#�˜ǖ]nc띞ފ>���]X_�x���䢖�%�8�-.��r�l6M�N�tuJ��;�ZIem�: �-���	�ՑYIQY�%��7ʽ�g�{ٯ�M_��Ǹ)FP�vV1S�A�Yf���U}�n9��@'�@�"�(���`)YQ# �X�Qc����6�V���*��Ub�Kh�b�#���Y�0Q��5��#*�m��E�"0QV(���"�"�EEDX1+X�U���*���(����*
�
���*�P�c��#V1QPV(*(��`�����b1Ab+�H�cmAX�`�T�c(�E�Q��EX��D��D�1UE1b��TF,TcTb��QQX�����U���
�Z����TV,Q ��UEF(*���EEX�Q1DUdF*���"��b1��c��F(��( �"���Db�1Q,0Db"�b����E�F*�"(�"��b�EQ�*��H�>C�Wl������k�\4��u�cv��Q�go�',CpRUip����]��aǍ+�3�7�M	��6w���� 
��v���X�8�G�e�����T�L>4�Wɚ��_���2��[��R��h;�|���󳚥v�cC�LECN�'��"��f�PǬ�ǭ�?��K�;��}fOIC��+MF���{�}Lu#"�P��fN��Td��5c$�芊z+jHf�źȴ�^=���Q/OL����v���Ƥo�L ��Vô�ً�d���s%��4E]��w���6�<>����.0�>��q�0��-�GoP�p}���;Wj�4w)���r�ZF�w.�/@�CY�g�x�j����U��ρ���"7��Ȣ��R4���{#��e�9���ҡ��z�c�b���#>s�,F@�E�lZ�s�S
X�$-����
;ا)�|�^�b�k���v%�j$�B����n<fz"\�����i���"�N3��]�fX��ح�~��gحL��ȷ6�E,R}�)p���TB��]x�v�����r� =��>��������JWO����L7,�&���=�����M:�����殰��0M��Ո���y�B��m�HT:���="�r�l#U�"�f[$�����U}����S�,��}k�#ܯ�m�2pޮ^�ԬO6�*ꉾF5e.��9��R�4�uN:;�b�Po\�p��ڔ'(��1+��<�螼˹��0b�A���F���e,<h�b�,ߗ�)��7�����>�J����E�����ţ����K�=2�� \��T砡�qϮ;>�)3��>a�W��T�ڸ�r��}ڗ,�VU{vj<�҉6x�J�Ln?���,�H|��~5����C�����t�jP}�L=����:ʘ�<�TB�9��é��ʅ+���F��h��M(,�\���c&*uXG`�R� ���=��/�<P8���b�u�y�ׇ���k�q������&�uL]��!��
����
}qM\L�C@�y)�R�xz{!���:3���Ez�E�:˃ch�WӐc�e;�E���q@Խ�+�q�u�n@wʛg�%�G�H�Rƚ��
�vύ�79x��`�~�4;��v���8HAy֞���ww��i��-)��6-Has�A����{ʍ���׏x��N$=�����wK��siG?>�261�IϽs
��v���i����[VGJLl8B.:%�֫�J�ӃH*�ۋ����B�����Nw\�{75|���fޏ�:��j�^?d���d���gn�����u�+�Z��go�ɠ�5yT���-}�%���&g<L�	4erɥ�:0U__Z��+7�_g:n�h)��q7's>��<<=��Ov���Q���#O�HS���n��v��WPgcv,2���*g+�����g[��q-)�d1�4�~�������<y_+��i7ޭ(��?�smq�kt�+R%F7�,3с����ɗ<�xe���JwV2�`[��!(��#�fڥ�2�y��H(�k(u]xL��/����z�Ca^ןI�]	��v3ت��g6�y���L�)w%5�0�(��l��Q7RA�nn
��k!��G�-p��R����K�T��^Xz�3��J|�y�?�1��:�~�1WϘ���0�,�u�zkc2�L�X����&L�'Z��5��6!yBĝ8�=�	��ѳZ�8�m���'»�GÓ�د:��Z�b���dP=��M��0�1e���X|
���2o�k5�qZܬa��1�J,�ܚt~{��E5!������h{�0��y�N�\l{��b��fwuP5���9H�Fr�D�9K^��k%�·�/y��y�R�M�F�U`rsO��{����,���`�����	��v��[�:���#�����V�)�fc�j��,�0kdy�Y��v�b��+��=�ӻN��3�z�덹��9ُ]��.�-�RQ�ef�ֱk8�*�1c���^h�W����|�}�̩畾��������M?�NW��WF`�r�L�ʆ[���p���n����3�V���1DW�z@�+�Ơ�����E,�do�U�."�BܘDd\�[{WvK	>�|68���-L�Xa��=��~�é��Ϳ<�.mR[�ʪ}�{���7J�z6r=���Ѡ�f=p�����%Z�(��uJ*wCk��j�)u�U��`�t�i>[Y�3�������Hr������(����L,d��]J�GU��l�x�E@߉H^$\�v����[i��q��a��N��9�o�Ckf�*��-�ڙ�Dh#n�g�Wv�M/r#��6��(�6гғ�+���H@�:�̦���B��1O9(��w�˕��ӯ�1���~�J$��U{�E.�=& ���P����jFjX�V�"䷼��.u���c��*d'J-�y�8׬$t�|6�P��:s-F�Ђ����k���]V�g{^�SZ�Ed���ic9�Xh_z[^��q~+��O\2��^G��%���g��8�(Ƒq}8,�d^������]���f ,�i=��Y��@R�ݮ<�`	�M�p�4�v���ǋt>�p*��rܨ�Z�:e��,|�̵Gk;r._tB��Z�B��*�+�sj����[��r�_Ͼ��{´��i��X2/�F�GB=\�\�K�F��p�w�7��ע-�\sMe�1r4�vo�-�O�����T��z;eA�8��WGZ���f�_��d`�j�M���}ґ�#��F�b:�y���|�4���1[�����O��}�L�=�^�<�yh���Hc��s�]Tm�i�⇟	�w�j�1_�=�+�z�������K�Rؑ}��)GDk�,G�CQ O �qv)�ⓛW�"�P}~'��8�~iuژ\���)ns��c$�Q� [ԄT.u,y@�hH��{���A<���#����^m#���L���F���T�|�߱
���.X��0��6�x����j�K�E�>u���b�3&f�����&���%F�WFE�djF=Y&s�r�d���2��� '��-YA*�O^;���N��t�D�.a���؛馮>(c���әU��n��r{W�,aX�J����ͥD�dї��S49�����}�6+���z�?��ρڷ��f���^��B91��gLw�;|@=��F���l#��yN�9���:��l���@�$��4�f��n��ws�����R,��Ť�}�v��ܙϡw&^R{�:�	8�n�jW�+O-�Wx�����dƙ����')A�*����C-�ޓ�u������}�  Qͣ���
o	��PY;	�ڞ^|TIb�i�b��7�X5�k��\ϗ܏W<��ź���N2�s޸���ɐ�a��:P؞��D���QqC���F=�=>}�:زj3V�\��>�B�d?^.6)�v׋#����.x:�K�E6aK��"�B}`�-Tf"�9�\�u�:��
�����]_��:	J�����L7N暊��Qݨٛ�{ՍwO��
��P{4�+��a�D{hCyz�4�ذ�h;�n���sswf�N8��;�ܢ>�u�J����|� ^zM�z
�u�6՟yh���}�x�yA|J�2,ۊ�1G=x�����(���*$`l��`t���7���0�Z�D�ɝ*�C~�G�wyج彻̺;�Ϫ��R�U�i�T�4z�TB�9�Vdf���v�ֽ�����v]�Rՙ;��8e��)_��L@	̓��]����@����b�u����(s�{�KP��Gr����V��dhق805���|']�m"�{��%Z����7EX@Jr]d
���Y��Y�c�{u�"�2��s�e4�J�D�J.?�Z�Sľ�e�c5{���� BVT2�zڗ[6�݇wbl��9���yD����\b�����椲U�6.������O��郑9�9��/��u���� �;a�^�B���WbO��yѻ�3��.��P]�E�5���c>U����#&v�c�~o|&5>����Q���G�ꛝ��a�-�kg`F����<>izI؀�y�ZP���>��u^T�-Has�A�m�>�*>K^<����j�I�L����櫷�*��8,�k���0�x:;��i�մ�S�47�'+!	l��S��v������UB�6GD3�CR�#!�X^p�����,5�
�|�˦m���i��]���������8(u�)���u�G���8�<W@�����}Bf�9�|��y�f��ΰY��uJ-NL�1�s[9�GAR}�+.���vHI��D9΢�Md�B\q���fZ�ˋ�"��
z,D�1-���Ca^�ށ�'ü��:���#�l���%�OΩ�ԋr:^���R**��	����rhH���y7U����qf�)���.W>�2�̫�
栋H�*s.''�%�F�W�g��ҠH��i��.�u]��AÊ&r�k�Y�(��ٝx��5����mr2�y�1�����뵯pD�U`�]CR���Ѡ�E�b5�:I>2�F��[t��p$Ƴ�@��yL�S�*;�5�˕�a��E��C~j;��r���v���J�_}U_WF��u�� ���tz��G��>�Uu!9���*%�Q. Wҳ/F���8��sn�<R���C��6��^�� ���w�CL�6z87gD_���|���W�u/&��d�f����dh�<��<Y�{<k�g:��Dt��S��8"�gb*y����TNFkU�k:6�q�	"�TrB�6M{��[��}oԺ�����J��:~�r.�g��u�'���<�LF���6E߅0z1[6��
h�C���P���A9�6����-T�k��F���"�2Aj(ԟ¦B��&�VmU�<E]I�(s����Xs#V*����kuWF���ԉsP�^����DG=��g>�ٷ�E�h���2�LE>���k���sT0@�ibC�x9_�.�o'C�{"�Q���d���l�Bp]_?2�c���C�m86�
84d��rvR(ȿob���j�o��։��
�]SN�=�&w*�}��u����M0�O�Bx��쥎��f��LE�;o=kΙƮ��u��6j84�;^ΡE;��:��$|�܋c�Rv��빧�5�ٵ��&�5�8��]x��i�,u��`*�2��%�ʜ�L��t��V�}�	Ĝ�!�"]�]Ge+5����K2�3%J�oKЈ�]ѓ:�~5�9�5*�n�@Y)/�y#g��U鲎m=Ei���n�:�����
��-GweQ�m5S]��+e�������D���^�J�@��D�^�19�^�<9���n2L�Y��q%��A���1�2�˗YR�����ba[& �p�ʕ:�����Q}C$��޽�Bw 1�@�d���tv�ɝ��&r�����K�>�!EZb<�����T��uV����d_d���lਉ����;=uƟ�X.�7��g�v�F�n�aF`�=�������|�S�E��@�\r¿/Wë��V��i����0A��3��3��c�rnwi���.��}��O��,�_�i�\a�[��|~���>kڰ���Su������;��u�Q�G1F <ٰ�	���N3��V���zH>W�	pT��uM�w/�>J�r��vb*��!��Fy��&��qr�l8�׊j-��F�s=�(�1��7�������~&j�	���l�,�y�^$�G�$Gs8�h'�1xٞ�w�{o}��%Lj���z8��l�5�?!�u��zp�7L���#�{h'Y��=crwv�gɺiwwe�yQ��D��9��U��f��5�wf�	�М=��B�#�R,́��ܵ��rolc��B
P�Έ7�����}��Q��u(χ=��c:ϫ$1���3
�i׋|cf��c$�}P�`܎��1\^�%cklU��H�8�����Ⱥl�٨����[�����]&n�*W<�MXi����Ph�w�}�,vuV��z�t]J�6����@"7�%s�=�=���WV�G0�Κ3`FF�׹
�����uM��r�,��x�B:�����aE3z�K�P�$kp@c
.:d+����)�(� ����ϋ�#_�vJ6���>|0�:O?k�ж>�ylu�D[�����S��lO6TO<B�C���F=��C�y3ݗ�,��T������^,�V�G[d[�=W�'�A�
\9��X�GL�2h�����;7�����E����?��]:���A)C���c��ӹ����˛���Ps�8�[4ba���S��ԏA�>4<r��.����SÓ{�#<��oG�׷�z/ry\�F%Ш~N����Pq
��D�茛�Ȼ�����(E���jOηp�;�����:7D+k^����ˣ��N3A��+��2�{��If�<�08���u8��Q[�G
�Q(麴�����>�*��«��ێv�]�C��m�ɓt-�3%𧌹 0$o���p���b�,��,��ŎE�����y�N��u�Cq=��4���w]�i�
5c���ĕK���:�I���\K?!���V�Q� �h�L��a�2��}�p=�E,�&3����m23sri�S��z-<S'm���"~\��pT��VTԷ�Yw)vs2u�0�U���履����U[��j��nݡR�d5�و��F*լv!5�VMU{!�
�n����v5����gbG�&�[c��K_܆Qa��W	H�}���3(�EtT3����b��)(�X�P���Q�%/�N��Ts�w�'Q�f�O,���ʏ����a̒N�	���͘:�B	Ț!���.:d���rb� -]�z=����G��ؚ���Gyۣ$;�x[��{�򤫣�8K%�xo/��9кx7J���!��Xn�F��T�wr�C����db�{�]����KYv�u�g�I�AFXH'YnQ5f��r����xU�����^��w]����Kb��⮧BD� ��v6Xű*2�Q|�s1a!���7&���87��4u9��}y���sԷ��N��B	rd~��uGRQ�9��.�:����MSՐ�|��ԍ)����3����:�ep�%rř�Ⱦ,bSa�U;WPܲ_Z��:o��z�rѻ��r�~��w�)�2������_e�_��aw�7��{�����#��r�g���ru<��`�
�:Ygq��i�T�,�~���$YL]�2�\���z�mF�6kȢ#���;�_}���V!��X�J#�����*�k8E�;xV�W-����Α�Y:���ft�5np�[�nڽ�
΋�i�r�P7J��B�We�/dRּ�g��qM���E� �Fi�p�����pI��&��9f�9q.뀾�XE^�|��ɸ�ۏ��������ޡ������N�x�� L�W7i*�q����u�(N��n��Չݚ�È����U;�
t�z����b0�g�VLa��a:�]m'gVܶ�7��\�]��wK:4���ٜ8g5�[����=����`R��3��s�v䂞�A�f�Y��(�Q�A�;#=��WLqĎ�uu�4��	O���*�t�~7b��NȠ��5Iֺ��k2fN#er�:��̎�U���L��#���y		Ռ=��._KZ��gW�|0��,�����V�X�Χ���;~�-�$]�ҭ��,jހfm���S��H��"1����hf�;����e���7O�m�W��C}�Pi�O%ʝ���'˱��˫�c,EX1U��E�(��ň""�UPATX�1TV")mEX�UDUF("�"��֌�TDAAU��+�A#0F+,X�QT`�-�(1UE�������PQAF1DcX��*�Ab��H�DU�[UQ�2*�Tb�m,U
��EX*���Ab�1ATQdT`��V-IUV[X�EQ�b��b�"E�((�Q��¬b�QQX��QX�QTR#QAEm�X���(���V1Q�QEEQR0��Eb*���H���E(�Q��*���ԡibEX�,F[Eb��� �TX���E�+�qQ���s+O[]i����بNj�@1�<u,ū0R��T/3���[zZ:D�zy&�0�>��S,�+�����a ��Tw�;y=�޶(|o��|��=���#Wh�cq�'��<����ʠ�+UW��{{��E\��]�zrz�,�a�v�,�q����P}����Q��5G6FK�"�Q��z���?-;Ѳ:7�1R������yX3�]�纼P1���C.�d:L��k�ܱ�6���>�z*���18=`�1��8��Chq�pn�m��j��okSԴ��	��#b"c ��>ȫ�r/��7�[����`�U��N����1�q��3�{Z����6����=�cPz<"�h��]>�߼}V�{��X	��/���N��Mu���qG����L�"GG�5s�A�m�>�G��׫7n�U)��+r9��Y��o�ī��fҷj�2�'�xW���i
Y+��n3�����,�p[��2ͨr}�B "�B�v607gb�_����ضŝ����,f\D��F;R��ݺ~2��)}�����p���bm}�Z~�����%�s�2��mY���<�-&5�Ɔ���,��#�ingMS0���k��o7CDY�tX�γ�=�ޗ���������2䑜���t�\z��e�O���W4��깾x���Ժ#�����j�V��.;c���X�u,t��w3&�����,W�\����e�Q��AF|E"6i�@K�fu��\ɮ��Iĕ����m5S*94J�5��53$��L��#�h�B���4��2�4�\�Տ�j��N���Ld�LS9���J�vf1��c�2�*Gx)�z�-���*#f�RE-��q�+��:���"�	v��>ɹ��7�����^�rg�J�sPE�n�`uN$�x*�����b�U	���A8q�dm�_Z�c듒������}��_���7�NLP�J'!��agf-�n�a���Eb�G��Ǿ��ɾ�r/FӀ}��!�44��g��X"ԋ�Тb"r�O,U��ɨO�5�C��9_K~,�¯��A���>k�!��u��y�	8�6ںX-�gw���%�K`���9�6��l�,���i���el�Kt��"��R��A�#41=�sn� �(~��.o���
����&��X����������Ai�y#��7\��(�=�˵WVG���q���qq��=�o�&�V��b�w��1���R���gN�ǨDO*�M��k
wV$���&2���R�N�RU�2�-o�;;;��'sGۻ�;˼��ݍ��d�Ѵ�t	m�s9�8�X9ּ�����ap{ۂ�=+�{>
���s���C�o#��;���A_ʯ�����x��~q�6�\��U!N w�~
�9�y���hh�)�3C�pe�l^��(^]=4�o�y�N�ſoa� a�>�
!�r�8]L�N�"�E��I�f2|�M���Ԋ7�OS����3�J�[�J���yAkU�2�c6����-<<gM/G`�v��E��j���k��b�U>bu&�z���W�	��Z��lװ:�I�rW.Q�ؕ]_W)~n���c��)��F΂m���G������v_�c��]�z<��{�r��=�q9�y��7T�Z������J$��U{�iu���q���R�E��$F�Yn�իR�y%KS} �tclb.d7*�����t����^��;��K�q����t�H�������zv��Ɏ�/<A��CUd�ŌL�M���jK�2���<m��nk�afgG���g/v�j�y���qcV9<�}Kux�3o?��]�T�č��d��b0�6/��}�����Q����[���~?C�\N	�/������_�_L�z\��������\�ǉ崐�ۡ����$��=�>�������BuJ!^�ݮ�h���.�(~n��.Vt��?�0�W��bU���yb�-Rg~#�iٹ�\�-�ɱ���tֲ}���`\�R].A>��^���2���ٴ�T-���\V)���߽�).�Z�o�iC~�um�OtD�xO�Yg��ӥ�k�X�_@.轩�H}G����n,|���A�b��j ƙ�S`�q"P���XE�ѥ3�;�垮h��r��Vi��������w2U���=H��,Ǻx�����sj�3V��)�z��tʮ���W=�����F@�0����Y��6xg�އ"h����Tl���S���[��}�,�K%0j�]�p_T��-������������j�Ol�8s�D_-��y�.�Dt1�)��H�*�#7م���v; �1��0���a�T�ĬY����w�LG����B�3��)(3�����?��;j�1���xiݖ�#��}nn�Vo#�qs����7��:��h4l�Ox?���!�\U��U����r����O����rR^O<�˴�H@!�TXUA��`m�X���6-�����X�o�6�=��x!�������iL���Q����/]�!Cu�����;�ډ>x
�"�e<#:x�(j̷`������Js��g�s,�K��Rw�`#���ĺ���V_�����+n�b�5�b��h��ݼviȚ�vY�MR���`��3j��t�)��rM�k�6lṱŬl젖t��R�J�eeEӥ�Bn��s��}�},NG��(�����e��{Ӗ�]����x#�{'��k������n\�\R�#�'�9/w�!��׎Wt�\����Wɝ�R�	�L��0��u��:	J��=������P�ײ�E�ܔ^JN��(�g�?���>�M')>4;
�{*�lk�b�cMCAug��9�1���)�ȱl*
�n�	[�2E����Ρ>^zM�����y���֔(P�n������p25H��Vx��Xؠm�4�B��/aHf��it�H�}g�/o
U1wY�R��Y�T�7.,K'4�*c��1
,s���/�����U*;�9��_�cVD���h(#&*[��`�%�9��Ȋ-[����N�F��i]�6|lu-���p^N,������Bb$pkɌ�	ƾ]�mv�H��~�?i{���"�]�E!%��L�&l׮O�����|f��?Va�}���Q����.���yO7�d�`,-,t�	�S>:��5c����,
��Jo�Yb�m�\���^�#�ng��H �d��Fn�,p�hC<�qK�oԣ�(���y���ө�м�[a٢�K����%B�Ƽ�N��N1)�����f�40_"{,�>
��亘��d']�#̘WjC����7��C��������!s�P���_��={�x&�U��1������!Ἒ�~|rd�"�-Has�A�\P����9��	;���,)E�.zN�u�{I��p��������ñ-���PB+��}UJr�~Xm������g�M����qT9#d(�|�jA�v63��خ���f.v�+0���+��dYP�,�S���)}��8z�����16��O�h\]�.��/a=G �}O��X��X���/7/�]��ʥ�>W�/x.�������r�:M��l�O�VO���nHj$tζ�E! ��@�|�+�MpCn?��,�wΤ%�i��o,���9�1��W �cB��4�}��&��N'|Є������v�� �f��Z��FNH�~1����c:Z[K��3+�S��V�K���������
��.F�����l���`'�T���*�9�GZ�<�5���b	ӊ���ě�C[�9��3w{��i�lŜ�e�u�!CS�vwd;�g�=vtE㡑#0���e�+G4��0���.�<��� ��1u�(,ܻJ��2��ӵ¸���uKF
X�/�4��0�̕:�+j�}�����>�6S�W3�S���aGv���Eޡ.79�fn��q��������[��j�^�Ø����Dq0qRj�vgv�C���� ��Ş J�<Y����g:�K2}�6O0B�꣼�'�5k9�ǹ���KU�����hu��.+����QRle;�}Q�{%�0پ��Ư�O �5��4)@�5S*Hi�K��Qx���VC���0�7���n,�nfZ֔���s��;�2����"��2j(ԗ¦	�nj��n�`(Vl�r�S+�����Gˎ��1B�7hx�n�=�sə��.}������
.�N�U�����bH����2��a�t��BaD29_�y��Ƚ�D��r*PL\�����Ӓ7��GY�7lCp;ʹ�(�4���을�2/�د`�決�����A��I*&�撯(X��m����@�U��a_�kbۨ��X���j|<��I[s�yY���3a��_;�}�ܙ��^#��a�-��e0.��*aΓ&���nߠܴ�WF[�{� l^O��*9�J�x&c�+k��^������9v���D��v'!ٺ����;V|�%�e5W>��n�Mm�F�x�U�
9�fZ�J��Hv�*{,��xV�JgG��e������=}ATG0�˞1`��1W��]t�n,2�s[���t�=��X��h�2[C{%��������/b�F�`�Fۃ�P����F���6�j��ш��ܨ.xL�Kɘ��:¶L@
G=�Ԧ9C�Oqx�T��Jc�%�=��g{]Ճ%ΧC���ɝ�N����bZ�q<0�m�{g�_ef<�n�Ag��z��g�Uz:�^�<��t�^27g��'�^�Z��ѐZN�4���J�\��]�����O��� ����%�ٷ/�r՗ẅ��ZR��]���^~����3��:�8�� 6�Ը���*��e�������5ܠӧgP|�>�J"����&�)�:0N�5�����q�w�j�,4i?��@��6 �ۙ�9w�Μآ��PW��_q�U�X�~��!��'<�qv)���^)g87��"�,ڥ�9t���zOP��a-��D� D��o"��&cfØ�	���FA�2��읥��^�XJ�����˿Ag>�8-����7b<g�����q8�V�U��Ӛ������-xl��X��Aь5��;s
����ݚ�p�0���a�W[�����j�9���]�5 ��]��^pu�|�kS�e���h��Fj�5=^�k:t ײ*�ڽ�j����U�c�J?=�P#2�fΈ1t\��5�ǎ��|L��V�N�}p��R�;�e�3E��ǳ/�=��E)3��gA�9�!]Y9���5,jNfjV9Ns�&ߎi��"W�.�D��n7�6'�z/!~�nb+M(��Aٴ�\�<�C��UO�wM�/8]�Uݪ�m['�@=�0y��v����n=z�\oKZ�R�wy������cz��QEE���v1�z�c�H�#O#>.�iU�b�V��4=�$j~�Nw�u~��pmTt��R�k"��;�a��:�����j%�
:a�s�twal�AtZ\���Y��PA�tP(#�`l�����2;�"�ۮ9�`�y<W}p����w5�{�߃��%_�ˈDʀ,�t|Q�FK���!)���ܸD��X̗����4u��fW`�k�\����G;�����}O���q��԰񔇱uH��-q-Z+E������"���E�ch+�E�P$A�t�H��P@�*5���T�C�q��y]������\fK#�􍅾�v㱳{T(~P�>�=�ǰ_B5q�Ѥ}�!�)mq}3������kwt ib�f�9=ˋ�N�4��ŃAǫҪ#�qa���y��i�g�xwT�nŌ��L�y��:��T�[��o�Ez=RB�2\�7������W�Ԗ�W�q�}��� ��b��k���U�@d�V���Ŭ�d�ԧ۾��=ӑ�x�|p�5��.���uŵvf��*dw���˥/{�7Lz��#�]��=���ɴ�V^�:6��옩n��G� �،EdEj��uʳ�[us^�}�Y���
�ϛb�sTj����l�&}�Ԅ�H�������^�-k�ł��5�|9��]���nd�&j2-��E�r1�P{�E�Z�����EO0_ez����w{^�D�t��P�⁩1�=U��;RY��k(\dU�>���wòs���ݭ�G:4C���-���PqEἚ�~|q)��:�k�b�W��[�j̛x_$����~F�@#'a�#6�CD�=:##c<����ğ6G[F.�\
7yC��s�9��ήW�=�K�ȹ�����db�s�l���!�X�l7���?XT�i���u�M�{|כ�冡J�7������� eA�s�(28�
�ᔞV��&_�P.��{���1)�p�e�	M�!`G�D�����
oMyP�K�;i��4�^���/�r���Z��y*�↶]��؇W&5)��k�|<��6:&^�epc `gg�9ys��Î�3\���S@#.��.;���X��.���v�:�������[W�y};]j��ۃ�d(8���`Ȏp�#pI�e@k�;���Ym�U���$̼PB0+x��=�l��μ�ujE��n7e�Q��vAfUmqc\��O$��y�u�
���7���hѝ��tm<�j+�oc9�Rx�M���r:��@Y���������"���q'���Nu�*�[M��W�4r�v��0Z�6-);����dK;$��ͽ���XG�ܺ�z��s��ǝ���`��8�v�ӧ/�]�V��!)@՛w��r�>ၥ�p�9���\���i7{wܔiY�(��1�в�t�nFPE�3�4E���'-���ˀ�Ρ��*>�qSKr:���7�D�tz)��4\���rY���uw���ҽ�#�KvmtR6�R�9`%���{n���h�������V��Lq׻M��<yFג�:Vy1XV\��W0�6�t��,��B�2�cy��Q�'<!��Q�R�7��+�wozQ���40h���s���k���w�(U��e��o/v[.\�}�m�s^)�
�����ީ#�)clT�H��r$�w*�Xr��PM	��9��G����iu*��+#���s軬�J��	�f�rh᫆��1��J���}��b�"�]Y�ӛ2�+(���	�٬���\���X�J�����ƍb��ŝ@چ)�48e��n���S$3���*����o[6*�-
q�������ۅtv��!���(�`S{;���j��§ZN���}S��u03�lnQb��lg�Њ0�0l#5[�˨=��n�N�z�/r-<�[ۃ�G{eSf���¶��Bǋd)���ur�0�K����Sk �WX c
����}f�5�/gm%Y�3j�� �7�*e���ZwҸ�گ^>�j�:�T���]�e��mgte��:;;���`r�ou�bҷ��\bzh�u����^,��/r\0^:Um��\�"�tvou`�Gjܑ��m�6\1b\ėT��'�r�d�j�{�\���ʘo����,��6�j�7.��t����N�=�r	�J퇦C��x�WgK绢4�eHn�$�R]B��9X��O8�F�7�gj�քח8�;@V�m�͹`_^����m�:�6�z2B�]�iT���tK�yΒ�'o^D:`m\�ՄQ��On,i� ��Mb9�A°����N�{�oh=l!|m��'CfaomwAY�t�ސ����iMv/y�g^,��Ї j�bo5&���ʼ��q�xPw2�I�y���j�����U�5�%74���^|�j\L��U���!������3�('�-�WFe�Iu�,h��S	,���V��q�vn�˳�B����8��۝�+��yT�;r5O*V��m��Y.�wY���O�����_<���k�AE`" �*�1�QTbE�#DUA�Ȩ�1�ڥX�X����EF
"*1AV�T@A�+YX,H�� ���1�[h�� ��+1#T(��
,cPX�V
�dEA�R �*�b�V(��EX���TX��cc�""��(�*"ȫQX�����U���QU�Ĉ�QQcTUDEU��TTH��V*�
+���AX�DUF*�b
,b3�PAb�aYb�
�+*A�kZ1���Q�M��qf8���Y��(V�����K�DK��4^�Z��E7���R,v��遨��X�f���.�/����a��vw��~h~��θG�ͥ틟���C�1��A����hK�܄�+�����r����=�0X����>��ڎL��P�j��n�c�q;>�h�+��2�G^��ů���P{&V�T��T뜹�_��|�\�UԎsQA�TM�o1�6݋�W�gu����W<�ϻ��%�bǣf'��j�=�+?1f!�dP=��O��aљy��B[�i�k���6&!���C!ߤ��EA�e��*�l�3$t���n�M']�݆��-�0P���l�-T���P6���4X�_9nr�-��	$>��0�x�l~����y}��LEP�@f1sa���RCL���� (�U�`Ed?�WFj\�����Խ��d�1X���ܳ���.@i��C�!hZ�"�d��5%�C@�@��K�U�X�N�P�ނNc��](*L�|�����t{�^L���>��30tvz�����K,Ŧ|2d�ןE�g�s�ǁ/Ӂ����~p����E���<eo.]ʠ�o>+��+��&;���4�c/��Ē�)"ks-�]�Ff֬�I�+u�54@����x״��;:}^�m� N��)5/8�%���Go�3��p����. �#��qx�YZ�J^f�Զ,f���tz���н�}'#8.jq�������+�u�k�5��6Ա+ޡ���p��Xxr��i�2�WDǺ��MF������Gr��s��#��x:�O�Cn��L+"v6�1
��Htq��%t;{R��y�7��맍|��>�ȡ�z�C��a�+�e�B�O�'�`~(���;2s^�Ks*6o'���ϓv�:���GM�u�����s�A��ԇ}'0�È�+ܡ�~�߲����6���m�Ê�(�.]eK���C�	�\��2�s]���f6 �-@׍	]4�*l�(��u�A���jv/9Sm�1/2&V�vxiG=�ض��A���!=_>�\C�xz���gD��kE67����D�d���(�-�k6�eK�F��3��?S��F.�S&���q�XW����s��̈�T���:�������s#j�K�tD�xO�Yg�Āڣœk�]*�ܷ�o��7�u�$��.�6��U�MRrsP �8*lN$H����,4i-
ǽD����fE0<&)td��mÝ�R�,��	�$yT:����'��$�l�!�\�ؿ�/<�Z͍���*ɮ{��S�!���Gm-���:��t�Q�� �x�Ns�����;�H��|7cc��J�u���ʡ1�;\����z�eo(,,3U�=�d���x����E�݀P��Y6��wDv��ל���]�jׯ��̃�;o�X0&xD��x�$�lۘ� m��3P��j��|���WP�b����k#H�����8�<�+v#���`Ҩ���o�^��Ǽu9�u\�%��5�#`��i�F��an�`�1�$�g�riIv٬��!y��2竦x�՗I��)(=���_4���7.O�Ozi�.>1c�l�@�rQ���{7�7TC�@i��˝�r��7��ٚ�!_d���6+���x��jUCr�B�u��_[tڴ��1�Z!_��!���1R�
d;���=R��Q&l\�#���;�Hj�7�������Jt�rS���A��7�
}�aK�d[��8s��jxYN�>�� -t��>ȸ�>Q5H+	��ǭ�z�����4���MSV���Da�#��\��$csa���y�R)��;ue׹O��yx��A��7�} P=]}���z.��W̄���[������7�Rk
�Ư�Y��pnV���6�ɼ��W�֗ݪP1�XJ��V��@��s��R��m�罗5l��1�� ���`s	��g�4V�ێU�;7H��Hl�O�]�0B�2��<Q��O��j�4�'3&�eٌ�Z�}S���>v&����<Rz&5|��;��>\��+�E,<gԇ�v�՛��`L���¶Z�Db��#��,-�̂�@�	�s'��J�*:A]tFM�,�=m97�X5{F2�i-�PFCka)�r6���Ԯ�str�p�rcҥD����7f�f1��ef���mxg?�՚�h����oƽT����qr��:ʘ�Aǔ�̵���Һ���5�q:-��i�ٯ_2(����6��2b���H�X�Bs�7��V<��J�u�v{	~u��æ�m�������f}[]BP��BD�k½Ν��,!�N�zćV����'~��G�Q)���ǎ$͚�Q���g��z~y��4m�(x9��~���\��?\�:�`ߚ,t�q@ԑ#�^h�,������Ev��4L�5�ܹg��܌������ܭ��!��s	�@[!���x��KK���!��� ��w���MĽ��FX�\aY���!/��eD>
�!�tFF�>��4^�lU�S:�g�#�4-���L��B�ۀ�1O^Vձ��A�����^n)h@�1\�q��&����B��6���*�UǲnfO������He���m������n�]��79Nu�c�r��P���芴Y��\�Yҗp@S��`Ð��g<�՘^�\{�v�� _/R�6
LdZ|�/��b
!CRU�����W����tyƳ������l�ˍ`�F�on�ʃ���#� �}�@���G����7��������1 wA���X�*��;r�,�h�Ut[�ʥ�>Q�,��>�'za��˓9���t���7L��:��ƥ�zw��".zl��H�ȴ��5��w,68T'�r��u�М�wc=���8ڑjG@��
��4��q8��.��u1'�W���Ycb������,��o�P�rg�J>�̮�O���?���].&Lפ��{���  ��ש��~�; �'!�G\����7	Ɋ�L휬b��j{�r��*۷{�N������ppzr�~6���!١�O�sw�Ñޘ�z欞O{ZͤpC�2$/K��7�1g���Ś�?�<UlD:�u��+,�IN�N.j4\�< ���e�^�L%��X\y$���&�>���-�S�/5ub�5yVU��Q�-O����)!D��x�{�f�bܡ/��n�f�[,��:2��BR5��c������X�w>�[+�����8������T-��*�tS�]��z\�*��T�l��e���ͮ]����ҺsO3�w���!���v�]O��E�s=��2�mW^X�4l5���D(�U�qYU�W�q��g�K0r�N��q������=�)3�5��;=D��@,���;��S��NED_��4�八F�9Y�^���
�|�����V
sP|�A���)�X^܎��t�/�L�����߆^͛c�.o�o�n�0�B�
!�W���ɍ��u�*p�[�3ɦ��I�Ludk1����m��=�4����喰�傫Z�zQ�w^Ұ�Wt �^'�]��z��3�ѝ�ժ|�6�@��Vn��G�6m�|��ͥ����t�^ӷJ�q�l��IM@{=3�B��"d����=e� |�K�y.�ާ��n�ި�w�#�1W��%j2V�ɘ��ڰ9R�x+ܧ�  �PqU�����Ns��D?V��-�R��#:j1���|���v���tH��sy`�{WY��ۨW�HH���k�
פG��ا,��s����Κ�x�ɋ<�٢�2N��|��UE3ӤzE޸�a��j����)Ǻέ����=�]���a�[�˫+e�������;�w-t%m�zWs�_K���{�98�Wj�H9.��֧U�\����Te��[Y�{A�3D��͝X��<�b���Y� ��'u���SJ�x�|k�2{>~�Y[��v[<��t�FF캲!�<E�ٻ҅^�os����]�M�FⅆϢ1�\Y�N.T�R��|}���x�:��[Ӛ�ԒW3����S��_�d`�i���tDϽ�>c����rj�|���4�"F#�={�|��^����	�+���
��;�F -3��ʧ T��Y�'+��;nv��\�闋�����,-3�����Kc6x�P�"`�c�<U7�o
�-m:�/a^��~n{���݌�`����z�7�Ks�&� 9ň�I�d�ݒ��r�R�W�R'AA���ZJǖ�D��#1Xؿc���F�\�`w�o�L�/c�\�a��9٭���y�f6h��c$��DTS�[RC46-��i�aP����5Ϳ��yJT�k�ĸ��>��wѣ��6���ً�d���s%��5O�g ��c}Q@�z7*�w���7qK�r�9���D'���oHB&��.yе��4f�#fk��i|�>r8��=�~�.`��hL��ѭq7Wz6+x/��,��81�!�t,�%��W.mF��oδ�NXW��U������������	^H�9V�ur��#�yV��gX�b�����;��7��'U�|D�(51XzV�ui�����ܜ����sL��~����2�C�7��T)��s[]*��
��9Q.�q��ݛW1Z�VE���+���A��:�)�C��J;'EK/��y�c�i�VC�����R8#�X/���3�#�ˏr7LOp[�K����R�]��v���	�C�*������	���v~Fz2�j����W�J�Xg��:;�6̻
z+�'���(��.��Y�RCR���r���{��whYq;�J�6�~Ukڈ�d�\����i�m-ٶ#���*̤��
�7W(,f���˸ȑ2��u1sX}ŉS��ϰe#�˿�@O6�X-<�G�o�O����ˏ@bH�}qe�u�oFʱ��U��a�(���/&���Emv�,Mn	CY��e��m��Q�2��(\��
���ʹxuS�G��@��v��З��o_K�Τ����v[̮xLYf������:��Q0Bw͸�u����Š�lq|��aL����R���D[�Aa�M�th-�4;	p��1�ӗmX&�Z^:�h(]K8�t������L_.���88c-v�	�/|�������&�B*�CY���&��aʣ����X�7|nz&�W�Z��T�Yٵɍj&p>U��[���y]U��i��t�&���\�m�sY�ci����������Ѷ�)�^|:Y17{���.ۗ�-�ۧN��r��4+5Q�G*y��٧��K�R�9�]z�`[�*X�]f�e".v�C���|�l��l��ԏ^tԚT���޸��^��8��WR"�h���Af�a�(3�t�3�Ѯ��I�jqc���_��ar�ֶ��@�,����툐�Y�����w6��h,/����x�iʷ��d�
z)���C�2��C��Vg���8�7;��Ջ�]'ޛ��6�S� c�W�/%ڞ���A��eZ�
����kXxk�"��E�����.�Y��ͥR�8$�ך�^�n4;���9����ݸ��1���m�TXB�^BU2����t�x����������&�<�oSY܁z1�#ʺ�g��1�^��~u~�.q^�+��'3&m.�b�ݺWH_�bH�xfu��$%L�ft���ھ���9�����G�^�t���\��ur� �t�˘9�f���2���ʀ��Q�lb����T�������[�M��'�%�oZ��������o$I��AW8���r)8��[��=�:bFLd��^G`��.�@���%��'`��I�C�z��[���<Qu����=�]�.�̦;h��	���0���Ĵ��"p���v�t�L�u�S�9��Y,=G)�2�����Ơ�`�PzaB�.�8��ջ٧[��X�{x����n��C)��؊�tC�5H��wg���\�����CV!PLt��/Enлx}t��
PdrǋdDFM�:w;��ɔ�qɦ��l^���.�YYU��.��1Fl�s�3º�F����kn��f�9;�z+���b��9SҶ�_�,=dS<GY��+t�[�r�F��vj���.2��uں�3�*:DX7����r�B���[���ճ͉�D�Pºlȗ[����<�St'S/P��,U맻�*���{��;�V���D�O��uZ�Y�bdt��[��W�I��9�m�bd$]��:m<$VչfR�r82U�R�soMɐ�,����F*c�}�w���&�d���>��5^f	�6j��Bʮ�n-�{��Tkru'����Ј�s(�OKo7���"sd�»��|�U�Yk��Y��wǄ�5XM�7VD;���G|5՜=F.놴�*3ˎķe��ʲZs����)���}��WWt{%�b��As���>�����dP�S:��լkuן|�$�;ՄS̬�$��Ս���T��t�7`�%Y�K�e���ʂ��і��{ie��`���`�,Ӏ�2Z�"��q�kݐGRa��N��3e�5��biA�h����M�Dt�]g\��9�R��A�%+p�"�a�6�"x�j�"�ږ8�*cy��)T��-�WY��p�Mm^���sk.�:kK	���4ں�xx0�A\�X���[�RN���3(���}R�QU�E&�زao�Wur=���2��*�>;�+�6��Ɩ�����q���9.�g]키�|`�.N�w؍�4V�[Y}r�];Ƞa����방�d��vn�a9O���j0�c!:xh�(l=B�Ǣ�hU2<7�ֺG��0fEn
=2��e 2�n��N�9�#�Y�';3pnRm/��V`���э���"���'֟��\��; ���;���i�lw��V�ޗse<���ӟ3��T�ڼ�Q^�t�!�b ����̀�ǰl������6s�lVgίc�&(�*⍆!��n���%ɣ+n*ݭ�͕Ԅb�"�ƬY=��?L'-c�r��}e�6ѐ򺃱�K�s����%���j�r'
{Y7Y�p�t�s�:/�r7\��Zђ݊�h�g��U��ܵZ�w�H�wH��QՌ�\A���4���0�N���o �Q^�n]�}.Q{+K�箹r�g.����v���v�C��7�eUF�8���V��6v��5!��y���P60���:����e�Z�K�u:%.T��θ�á=�Л2uʗY&�՜�9��v���U�/b����0��-u��j�ov!;��!�r���>{��53KR����2�d�c��a�3r��Z�O�9:P��3����7�C*�� ��1듲u�,��E�v�Y �*��o�!6挦fU�[��1h9h��P4З�yNw�ME�|Z3� ��V,7O.k����|�`L�=�fq�!ͭ�����r������#p0P-)��c�&2X���j9�,����z�a+|�����U���d�J����[C��͡k�"q ��mH� ��F�U&4�
������W�ܧ��TH}��\J
��Zʊ�X5
ƴDFKkAEUV҈�QDk*"���ȶ��`�T1QV�4�Q�*�lQ-�U`�6ڥ*��B�eQijDjU��m+-(�*[V-kk�Q��E��m�i`�%�[jҖՊ�(���IKX���F��miJ4e+E������[j���*�QE�#j��l�mii+H���J�lm+m��Q��R��h�6�cXR�ƕ��aX��֢+l�b�e������2�U�l"	J��R��k+am��U+Q�J�m-�-�DDmm��֕�j",X�4@��$�@&��07}أ|��Ι�7��N`A���D]��/~�����ytt[4���y���Ȥ�p3ws��G�$�Z���9�s�u��r�-�IE��5Ҟ�s����z�s���WZ���6U�oa��֥QC��؂��E�mX�;���J9�]Iu�Tғ=g"m�r��r�5�-`2����A7~Wj:F'�/�����'5X��ݮ����
��:�Up�*��nEn�����|��xњ0?X��%�j[��/�r2��\W��P�4#/�B��w:
�Ω��K�~-�;#&�FwF�֪����rM�d6�?:���oF4�z��R�:��um�ÓJ��y�zΪ�o����O$I@��t@�rq�D�̓�˸�V�[ӬFb82������{�u`���M'�qUҩ���jY|rJ�h���e��`r�`�ϸL�0�'��&�
3O�l��[�;�Rӱά="&�ܛ�nh*��l��p{�I�ث�ky��鼭��� �����W[nV��V,��B��cZx���im������qR�VbH5)�ۥfw��l`��Z�R�&z�GS���V'B����)�r7�(<��B�{�)T�-�Gl=ʊLWW���mgw.3{tt���-7�����[\7��5��dD���W�j��tFR���9���r��jmq�=�����N�O�����*�z6h:ݷ;�v���ms�u컂C�������y�].��&�W�^���ɜZ�~��ǯ͌�潺�=��:i9o��+٨"�G-{����B��7Wd+A�C{�;S���v�)�7:y��b�XD"�S�7k�[ބ@�� a��ɞDߚ*wg-��R���m3���#띯A3��m�q�!N��ل�G�H��=��Ɛ�W�^ �.*�b�R8����P\r�NqY�2dh� �z�)v���F0�[�=��OE6.�UvDWv��|��?mE�������o^����z�q���2�OE^T���҈fxPn⚉�	Pv��X�D�Ë������ؙ���[qC��j��W{/�6�+b_!wvnkP]v���(�ج��F��Э�,�g�\��S��'�X��y3�:��N��׷��������L���L�����������V�kbu�'j]ܺ����joCl�д���i<|O+b����k�-퓡��&���YX�Ҭp��ur�3 ������5`���s�\��"X��FA��H��H�1�`�G6�X������c���I�Mt^�*�zXU�9A�y�'T�o}�i`��v��Ѱ�e@�c�N�^=A
��F��X�8�����ՙm�x�T}��4n� )�9vIg�K�T��B��	��E��Њ���o��O,w/ju���^oNu��99�������@�Re:!&4����>T��s�R`R�t���Yz�O,`s�>����c)���2��<ӔZ0��B�o����������#Dz�~8U�#t�cCsPedr����f��5�p6�Y��V��܃��>X����ص�T炮�7YH����È<���r�Ξ[�2e�=�Z��\�w���
��ls�gu#띢��1o�,uUk���\a{K
Q��cR��.��{�j�#��L���]J�<����9�/ɛ)������[�#�2㰞�{v�ճ#��o���U.j�]�����G��jE���Sҕ�ȇ+`������.�/�y�-�w\A"��)��-�l�u����x�B�b��@�,������pW#2����z�f�7��,�m[���X��^W�]8T��f����B��'���N��g�k�������1����OEb��F�7<f��뻮Zف�9�2&l�VN7~]��Yq;�J�.�o��;��ղe�&�M�_������!M�����wJ�:�)'��뾖[��4��ݩSQM�����s����0cgwKʻ��O��=ו����bJ�άm���8(.p6܃V��7�zt��ꢧ˫ۆ���
���O ��'`��I�
���rd�\�Ӕ�f�a^��9�y,vY�ۢS>Bg��"!1e��4�1��~+4=O��q,�}�iE=XQ0-��%�ۤ8>�'�cQf�u��5��ҿi�䘡j�	��/�ۻ�*\V����<��W���U�A�xn�0�����>��y`���E��d�h�������۾�^�+S�!��s�����HK��[-.��;�C���*�j:���\��]�u�g3��`ݶ�k�oov�	�H��ŕyWo�t}��Sc����u;��'���3<��Tk�M5��Fן��m�nлyr��ƅ(:��Af��p����-ml�s[O5�ɮyp�;��3^���VQo�]!���к�æ5�u�<�[cHf�{n׳��PV/��9V+�\��d�{��^*嶑��t#���f��IE���k�9y�]8T8���;�`���N���ǧqr���\}���I��`xD�s&�����3�.^�Q��A�g��"�]@w�q��w��V�*A�Cc'�ʸ���m/�Tc�:U���<k���[���#���u.���R{p+^��w��Ҹz��~UhhF_>�Iڏ��WO5*Y�3�ݎ�y�Y�*	�V5��i6⽏�׵lތ>�EgVDt�/�c[xifUu��*�Y��M]�F�/ub�ؙ�`���pSѼ
|qj�#suI�h=�[��"Ţ>wOB�Au-�[[�ō��3�7��9dg,���TGL��x�&�s%l�I1�9d����,.�Jn��MVqD��U��ngG�ez�>��z}Z������A�H>��6,��绰��S���χ���o�Lv����/�xO6�C�;��c���N�v���=5/���ı�VnP��l+���G	����}�\^\�9W���K���ў�b�K�`�cx���ʼ�nh*�[��h�e���xs.��>"ľ�18"q�����3��=Y�.�l�>�C��L�U�N��;�Or�>�}����.�7�f�����)���[��p�sJ%��\�,�:Z��8�����^�|�g�i�ɦ�>8.hJͺƑ��j�����=s�q�k��y��5|���|⯽Ōگ'y:���]�p��Շ��}�ȴ¦p�eq����8��k	RZ��ml�d�`��m퇛�vUC������8#�m��A��z�� ^��US/�Bǥ,Я&D�y�b�W ��8о�F�B���Hi�x��n�!mm�O}�r��e�4V�aq� �Y؏5k�\�y��Қ:jWZN�4�������v�$4�v�'��ޮ�E���J�^f����6�u�^_<�#��@d���{ӟ���F!�{�+Ɨ)jUX��(��P\@���5Sp���N6��W{�5B)�v�J�����AP��u<J�G�UA�[#�:s{��ٜ]V����}|1��m�j:4b�N88Z/��ef�M�\�q�����W]��gw�Gh��m*����~P��Q������c5^��E���+��@w:8ݝҬp��ur��̃J�3���R�nsYWH��o	w0���)�˰v��oޮLN�¨��MQ�ݒ�w�ۺ��BTϟ^�ʲ��_\��,�F�v�3>�:��K9vOu�`c��Tp!x&k-ef[r�׽���}��\kYT��NH��c���C��o �&,����B*�CX���w:��%t�@0�C�do���d��ʹI��`�
Ge:I�֢���EP�Vx���3k���"����\�e�r���]�����;��c.m��\@hq�r���� QQ��,�#�dmJWʯ��f��ޢ&%�VtȎ��<�\�"�Tee�̸��k��Kc�F��a�a�0gev�0W=�H����x���s��{��Wz��Æ����L3�Q,�����<����<���Zm�\B���j�[�79��ә�>�j�06�2xÝKj��f��#l��<�+"T(�bx��ps2jZI%D��u�09����:�~��nv�ha�����V��F��a��ډ�X�Ǜ���[ޅ`�b��q�b����K��]�Ya�ۧ���;u���t�ŁOl���C��|�v+�'�����I*N���$19�J+��q}�����[�=��)��\UD'�l�\O��e���,��爢����}�j�>���֯�^K�=��Ꜽ��nƉO/�K}��~�"'�a��(�m��u{Ǥ|�5�"ct<����=�J2̞���΂���eUGj:^���*�9���ᷜ�/�V�����jsm�9$l�"��o΅�j"v.qPz�W���9���f$N��J�U���Fm�)*ƕ�����>�1r�Y��O%m���QQ�Q�@٭��J���9���Ѹ��Z�XyX�sNXUp]�n���F� ��[EPgZ�ö�׋�l��R���+8$PWP�C�0�#���b�կ�&D}@�H�ݎIr1�;U�-����E���8%^�q�5�DnT��������Ž�j�����@�Ԉ�mP�aN��O�NJ�'
3�u�q����ܬ/�.�d�:z��(��[(L���	��E���0o"��-���bln\f�j�^8���y@]������t���ޢ*�o�	�\�~�;zt"��j��i���x.�]7De!X[ք����"vb��y��FL�?,cf���W���My��ڻxE�q���ȹ��<��qo�hk}��G1y���Y���h��l���JYE���
U7�C�$��ȷm��]�PU���7��5qA�w�h�z���/��ڝYH�>����֥�+�b
�YV�%�7��J����������3p5e"����s$_0��h��(>#\F��M�~t��p�t�F�{��ݎA����쎧���_l�t���ku�:�]��]ѫCPR���o�R�5�e	Po��o�8��ٍ�Sn$Ã�r,oB9�E��;�A�4�eؾ�c� �����ۇ��� dśfqQp57P�tz�TX���Ix��m�4N;퍸W
���Ȟ芳�m,����4�pp��	�(���nƕګw؜vQ��PV��4W'�|iv|�d�`9衈r?P��U�!~=�k����<��B�B�/yds���1���K�)q�ȡ�t�ec�����ױX\��w<����{����_���-# �6��kڏ��b5٘���mqE���^�jj���Ε�Ԫ�Xl��F�Jó<��3�+w*c� v���F����v�soD:�ӱ"���o+.9k\���1�m�.@:��p���8%��dw0�+z������4�5m%��]&���Ϣkm`�ʶ�t�#)��P�òR��.�R�o����bhkC��O��{��hׁ*����u"�9���GK$u�v�[����4,����٢�|"m�٠�v�� 8j���h��y�ۛ|8I�m�/!�Ӷ2M|f��7� ]M�8� �YwA]G�I��A�8���^nw>��'\�׋"�r�e�	���d�<�hp@�T�\s�����$n�+][M�z*�N{܅�΁J᠜�1�3HL�Ʊ{i�sˮ�6G�AR���vGn��)�u��B�I�-Mݺq��D�iu���(Dn��=�Qޢ2�r��3�e9���|*+x���r��t��sy�=�zVC"�P��Yr}ֆ���Z�o���f�Rቃ.VNɫ���S/TMo���\!��n��q����9u�*�t�-�����4�ޘv�� 6nT"�ѱm�,)�?��gc�M��6�Ika�3t]ؤ�����徻�0�k��!w"6��&^�7w�Z*�m�Ǝ�V��=���8
锫9�{�۴���w�,����cpê��&�e�;n�nrf��Νob���2Z��������X�c"�+�/+�i���D���� 7��N�_3�M�D���rV�0�w7�T=t��Rsh3�֗��^�X��r末��9[�WuY�Ê_�I�u��(�W5��VZ�`��G�]���P�͜�J�i���s�$U��CM.���c�@���ea�\�O��{yZ��r�
�oJ��ƚ�[��]W��P���^��Oz�i[��]���{�&��Z��@��U��"��Ӑ������%�ZĬ���!���V�7ʝt	�l��MfVXy1˩�>�_R�%R+�˟Ṕ���r�N��١'�7�}2�֛��!ŻJ�v9jc�<�
�&��1��KM�w�����|pU�4W;J]�bٳ���G[�܉*V
/4-���U��
�3Ѹ!+o�OjY)��\�����p����Βh���n�{���Z�L��=�I$XI����$�M����|��k���T72�v�����z��u�n[�w��ں����Gj"��&�e���ꋋP1�r���Y/��Yںy�d�D�y$�5�许cA�e���\�yR���w{\�v�8���賮�m�^�#6�+̂P�);*Q�mjZy��k��)a�k��2m1��f��⢍X_t�͜zo��ጕ�w���/��K,�ù��|��yҦ�X�um[���f��ӫR�F�۸Ze��ح��8�P�P.�m�P��8�qe��e-uLH�Y��]ٷ�]��li%�����b��co;)!oc7���VC�wW�=����N���p˵�ˤow��P6�]��1\X��	ŕ \�̴�L���]��ݚU�DN��-U��*���A�	����}]��J7\u�6t4魰�������,ڶ�kR��r���w
��Wׯ�`z�.���"O=��]��s"=�n�+��9���\�S�A9OM�
��-��I)��D�K^u�FT�9%�N�nU��iٳP�}�jvľ��f�E�Z$cR��6ԕP��mJ�5Q��+D��
%�Ikh��T(��[IKeb���VQ�m��U�U�նV�mZ��-D��*Z��(ƥmiV�j�ij�Q�XTEkJ
im���*V�����ګ�QJYQb+�Q��QmPmV��[h��-�FХ��2�b��+km���J�ekZ���Ң�m�
,��J�EZ���J��P�F�Z6���F�-��Ʋ�bԋ
���A�kF��Z�4�R��T�Z4���j
�QV�Dm�QBѶ�%J��%E�ʨ-�
�-)K+m�Q+F�,��KQ�R�Qb�
�E`�6TUbV����kT�m֨�m���clX-B��)F*�eJ�듙9r��m>;uҶ����$w/�e2�XM�*�ãj{0oN3!���bf��/� �:�Z��M����,�s��/��Գ�����=��-9������ц4统����f�V$�/n��� Wq��@��f��������X�'`L����q�'r5�����G�R��hm���a"��y�yeM���OgW$�Q̔���;��8��	�F�J�b	���W|&&׷ޮ]u%^$��qaN,y�=��j)�\U�b��D�����T؊��I��OGaI,��u��5�����z	����B#6�踻���Q�b�+�Ӝ��v���Gc�-��ѱ}�i���๪]"�>[\5��(��j㍐�ydv�bw6�N��i�P����[
��\�ώ_�9�&78��n��V\�V���������m�[�O���~��9�kڠVZ���b�9���b�y��m��DIR`M��klA����Y�p-��c�ܕ۷J3K��RX��.wܣ�;pU rN���Q�ͨ��!�v[���f��œ����]����.d����y�Ӷ8����͡/!��;7w!4j����ř����C��\�=Mj��7_,%a&s�촟����H��d��s��~�g�8�Ѵb��^�dlŸ�K�P=�׵BZ�v"04�T���f��V[�t3N����dV�#���Us�J�O�GИ����B��Ng"�s��z�2�����<�z��M�m�[~O����/h)�I��������+��-�����^P��7M��*�cz��u:/7f�@X��or/,�u���c���݉ˢ�]!�cB�\�ا(ogM�Rf�)Y��VT���^�,�����*�u�^/h�bD�\e�7���	�#V5�*���l��ͅ�`�{Շ}�V�y�Z�$=��g	ta�sO=JTLr��K^.�����y�]6�*-�W��$]��-u{���ë��1.:�!6ՇK��d�ˢ��邆I�����0e����wp���R��g�ʺ�ة�^ʎh����q;�4�v���Qn��r��i�?p"֞��wz��+-�C{�uu�H���[��a����R%�u��Fa����̓w)��4����46���7�̄�`�JVwo6(w�u��M	�@�涟v���Ɛ�Z����+���{�gy��{y-��"�	�W2��΍vu�[v��j�Gke��^m�۪�䜒�kԷid�.F]�q^��K#Q�a���4�5���f����<�Gv�hX�*����k9$Z�(�ߝZ���s��U�x���u�{��<9$��3x�,��ucm<�izZ
�8���z�\op��ǵjޗًOXR���dpi��I��CjH�f��9��:�5z{-й�]4p����xL���	�j,NU���z��vH�N}�\�5�1�4�p�gdX�����buT-+k���ۣOkU��{`��U45�ݷ�������G�HW���S������;��j�b���N���F��)��z6i�e��B�a���3D��4���G[L�xv�<V��<=��Ͳt=S�`4ĸ*a/!��z�PQF��z�3�op�h᠝e^J�3 {�U������;M���7��U������$���	]]}m�e��pҞ#�4�O7雥[���]�#�������זg8f���z�̎]|�h��y�>]O,=94Z�l��?�dQ��2{�
Ҫ^Uv�v��n�֌9��PD#u��5q��c�9������p!����y�;_-���R�ej��VkD"��w���V��o�;�:d�Ǽ�ew��˫'�.gzE�窞��z�A��+ܝ�\�J{2RΆ�.!P�}+�OE�A7����<��zݖ���痷t�7<@���݇7��49o��]�J�{��gT�)؛g�S�1��S\��g5�_ucq����.ԋ^�hhP�^J#�*^��g��R�����bn�)���賎'�@�����V?I�g;�`�t��v�n��f�bj��[����`jm�u�Zy �P9n�u�v�%�%�iv� Ϫ�1͟`�G2;j9����^9�ݜk�E|���w;zƖ���h�P���EI��.�5��h�*� ۡ��Krǳ��{�?Hw<z��(�f�N�jx{>u;�����ح��SZ����r��o�p7�H7w��a��a�OܰN;Ow'��~-��d&�T���P�/m��rB�noi�k�W�*XU��<�r�[Y����I��qo(�F&r�^�Q3�j�%�℡�D�YW�m�3B�ouƵ���Yk�w*C�!ζ)�,�&�M��|k	�'����*y�t�pc���f�u���)�脘�-|"l>�2���Nq߽\f�@���9�!���n���>V�.�D<94ч�-�v�u��m����[Dx7�Z�V�m�����ͷדFPSD�\Y�����]ra��kX�
{����Ζ�z�t�G��w9��:��]r�0��rUu}Ɇ�8�إb��9꼘�h��V�z.���d��>dY���S�Y��X��c��{g�����)��e�r�#*�ZEm�2ޭK������"�%ŵ�Þ�V�Pl*R4t�Ɔ��Q��L���깙}ã��.�$$~d��:v�̂�a{���{-k�I`JRǀ?���]�h>�?�V���V�afy���S<��v����7�Y����� ��$�὏��qN;������8�
Լ�jgp��}N�R�Sn ���g_,u��&W�]��?q��u�@��۹|���yQ�&�=�i�U��=h����g҈=�l�W㍭��;3�����|�Y:�[�;N6�M�W�oڌ�$���-�;�Ys��A#y�0_>�U�Erֹf����!�j=kڠQ��{V-��M��59��sE���5��qF�j�%i��N�h��P���7���8��j�̂��O%�.ݎ�|��yD'`��A��dL�Z�W��m�S�A٫ޝ;�{6��«6�tJ�pr��b�j,M�SCX��'��\27*���{�QOV�L�=�����+��I�>�^	��X9�I�Zı�N�s�Xu���M��˖�%
[֖˥y�j�ߺ���ʉ]��Q�ɦ\W1A�釺b���0��1#i��v��9*��f�x1�q�95֟<4��ha���<c6i�F6�r����D�a�7��x*���Lj��c_m-��B�*�(��4��Ǆ�
oeuq�+�tOG"��^�Ø���� h�a�&����*����2�<!]Z�ac�8gWNd�eCy�4��k}�����ɾ95�b���*�b����Z��m���C|Gol��{�X��u�X�p7{=a�B�[u֜6+k�N��3���Ǐv�;R��O&͓`\�T���w���C��=ՙf�OB�1>X{�=p��Ƹ�E��jå��^���]���Q�E��
0���=���KOk)���8��Z�R(Y�=�����0�%�FђԨ��:lpFW>�E΁�ΰKn�p�C��6"Xg/m.US���d��2�.+�V�����ʏ�y-�	P��i�Qq��dbL���I�P(4��o΅�j"v�q�AMYS���Dk��+�T^;��g	���8�<�}K�
�8���)�Xs^V0��Ǫ�oh��ϰ:g��y�	�-<E' �����mN�]n(�H�Ƚf��W7�Y�����1t�����g�n�f��:m~M�V� ���-O��X*���<ăC�V���k)i����)0�-@���hņP^Uʺ�����Ń.�8���6`���Ɵ)�*��R�wʭ� �f������u+ܡs�h+��-��w�X!;9fw��+��'�m��1�t�?K�&����4*����C8<"n"V�}���ί��0O�cBqs^�U����M໺�D�+��0-ҵ���x���]��x0/{��ލ�-\>~�:c+ؑ����g��h�vҎ9���or}�V�X�]O,�&�W�PZ�:��`�3�$Oq���kT�~]���q:5���ś�]{%f�r������w�s��"�yi�l�Lv g(cO������c����}�ϒ���ߢ)�:��e���x���X��3<P:5�H�'���*�2�.D��`)ܝ�j(;�T9+�GP�_P(&FWhA�Ն�:�\�Vj��y�	�v�":v�·Uv��v�\�1Z$�ģ
��q���Vy��C�{3�����a7j�]x'C�3����M����c(�x�n��Ν�d�g!r�e5�	�3��[B�s5hܜ����mnZ�m��
�p�0�q�cL�'j���_�ooG8)>�J�3��p��Z�7N�ם��inﳔn&gCl�P
�sCB"_)�$��z�;�학ٹ�Y�w�݀whY؝��FAm�{�&T_�s5��mvuE�}��uGh�4�ڎcdn�W㮕[�l��H�tw,E�ٗs����Xn
�<���ղa�pe,r�&5�Q������1��vN�7ܳg�?ݒE7V9�ǔ.NĊ��H��[�G���n�����)�kD5��"Zq1���YW��m��b�Z}� A��:����0���;�PI�-E�hD�CYg-�]��yC��������ո�ϸ�d�[���tBLl�Q��SCdt�t2nr^��J�I��b��7u�vx]6�,g˩�xrh�o�('De���N��SUၦp�YTy�P��hVoQ���+��Q��L���.ц��/i�!fܸJ�f��[�4�R
�z�`ŵ-`��|�v��)��]c�5�O���wLmO��u�o�8o��Q�W�\t#�Oc����O��kϼ@c����s{�6,����	-�e=������g\�Z�=�ׇ;��.�3��2����مt��b���{�߅e#s��Zh:�vQ��8��M�%�f뱦�S8�p�8��V�*���=���(>鷫{�2+��٣��]�xn����Q��=��bC#���nu���K�l��Z���>��no�}���b�k e=9ő�q�v�J����
��U)Flĩ�7q.S����S���������F������y.��\��T�>ދ�A�9��˺}O�2�F�<Ex�F��`�g�v�dq���N���c���魈k7���������V����MUF��;�xַ�~�zӝ��o4%h�M�^�o�I�̂)(��ukڌ�;��CڱmMvQo\"{�e*�C�g�r����Kh�Vw#i8�AW8�wB��H	ig7zx�⻒	��,�O�1s��P���CNJ�'
��jyL��'8�,��t�R�2�:K�9N���u^lz��kE��p����M��3OHQ�&���}������&�xX��J����g\ �3�lgh�N���KG*�X색�9�\�Zj������¾����V_tc��W�����N���}��H��ǜ�����s��+b�Y�9\�3P�U^f{=��}fN��@�3=��Ǘ��f������H����s��{��f��<�^���ov�cԚs���cVɻx��R�J�ǚ��m�L�;C����W#�Mjד�P�@�C�cLV;!B��L�۝�jrˎMnN�IܩGcJ]�[��V��'��[����A�`s��xl9Y>2�%�Z*0m�*�Ä��3�/%��������ޝ%�{��Er��qm�@�b���v�RXݭ@a��9.���}�uе�M�a��6��;"��٢���9d&�6Ş�ٙ���X�[=�n�y�yo7ؼ��K�Hk5*d�pj
�_neMQl	Y�f�u�H�Û�,,���:%qNv1�ZS|��.p�����.uq���I3X7 ��$��k�&�Fzd�;�X�eLˑʬ�q�]QJh���P�����siѢf�&X�ѽ},���!�}aAt����`�Pz������$�Xnw�lCNN�vS@��`gێc�<�r�����[�Л���W��E��$��쩤�y�]�+{�A��YW��ܤehʝd�nA֛�<83u�u6A��]0ȡ�3�L��]j��E�Uwg;k[�et�����:�"wi��R�dy��Ou������k_\9=�p��G-���|ťܙ��)�(}��Z\D�]�
;Tr��u2Q�E_}���d�����]4��`�t����YE�-��������]l�R�j�Z@��o��� pߑu���C�Y�����;i�2�q1ܦt-���s3GQ�36�fuP���	}����_$�t�L�P=���0^�L�r�]��!M<���GVM(���+�����*�����<���l4��w`nퟛj�f���u�����,!�:�i1��w��=�jY�F��F*<ɒ�Q��0;5��ӹ���x�қ"c
��]�s�uNaLR�uv�|���{qK鱎��5[��]t�zVEp��Î�$,�B�nl731�F�#u;��g`k��u\�]�j��x�)��ʳ��nl��D���|i�m喹9l�Z���rX^�� +k;�"*�x[��dw*ge��Ĥ�����Y�Z��� ������kN��gV檾�O��#�G ��_J��'JA��W�����;���r��@aU�!�ڍ�{���K@�J�{%�2d�r���A���]wc�]�%]	.��d�M�r�3ePV;�B��$3tN�jz-Ek;���#b��2�M��*M��y�ߌׇ�O��E�b#j�J�Զ��ZZe���)PiAaZ*(,X6Y-�Z���X�-b5"!F5��,���+-��DE"ZUm�UJ�5R�m
ª-eKZ�F��Z���
���mT`[j�R��6ЩX���V�X-m����
�PD*T�[m�P�m+m�#i���R,X��Q�Yl�UV1T��Rʪ���mE������F,F"#iX""�ch����E�����TQT��X5�+��A��¡DV�DPYm�`�V)QA�P��#UE�V�AU��F�TYՕ��Z+��IiAZ�`��Q�����e([j6�h����DZ�*�YV����"�VV���$B!��!U���x�欵�`���ƻ�7)sw[�\k�������8'I�����̆�l�:h���`B��.�L�Au�.ѭogf7+�n���J��Z4K��y�D&,���4=ՊE�Rw�]���nywq4W�d)U�x]���t�n����$�f��X�a�?�)�Kӻz���[Ꮦe�������2P�-�7�U`�Y�e=�oYS�_9ɝ�ǳ\�c��t��;9e�ˤ0��}Q�L�f8����U��'��Y���h���Ya�2�����/U��Zu�_�l��v���ݡ1�*���.�,y������X-�:i�]��L��5��Wm���;XR�㊻�2GP.S�W�/<k���x^:{��_.D��.�GW�<k��ϓm9V��{$��b�}T�g.1#�����4�p{�]��	��xsW����N6©<U���4��ٝ�d��w#^��7�&��W"Q3=�T�͢b��$05�������j�Yl�؁Ww^A��<n�v�G��q��e�ˇKV+���C����(�����ZUX�M�y������B��AT�*����+TF};�[��ge|��oOmcU��;�6Ι��=V��E�t���j�_.�Bz�t�2|FS��ʼ�5%��*�j����]V��k���*�X����8�c]�g$��@�Ҋo�׵l��R�J볡%��<߷�֔T��ͽ�^�=�}��m<�iy����؎v�\�l�ck�W�%Y��,�s�0e,^�����	�-<ە1S�j*-i�T����Ӱ��6��(\����H��xL�0�e��#�bxNIv��+k���bhkd��Mmؓu�Z��De6vP��Zw6$��swUN�]<��ibkZ|�\�|"��f[�W�.�n��;����\
�[-��a�{[�-�M�ɭ\P|"|�l�u�o+v�dK��oTf����Zky����7�Xg�3���ޜ�!����¤�f�ND�ۭ��jq%��_���nx^ct3PE�\���X���x�a��-y�\ɼ[\,���x籘�T8�nɩ�DK��ub⻚�h+��;w����L�{�Nu�G���Ω"Z�&s{wT)ιA8����Ō�=�r����*̕�Cb'\�1WD��0.ઋâ���b�/oT�m[Zٚ�T�Yak�p8gQʱR�����浨�T��ι��e&[攪9��(Dc�c��ֻ�3H=��Sf:�zwg��Q�k���,)V��w'l4����G-�x�/�	�����41ic����Ifn0/�j8��n��#ӱ^hr.����Ք�G!Ʈ�׳z��	�u{�J��@g8Ӊܖٟu���ҕF��eL��Z��^zs�؜�r6V���n�whr�8�M�Rw��2�5f�h<ON�>�3��Cu�i�!j#1�7t�:�U���ћJ�mw!��^��|dI�s
�@�2��'��#R8��P��E���˳ou�Q���*����8��gq�r�[X0:O�4{�qԩŽK�P=�\�|�0��Ĵ�%f&��
��m�FSZ��ww9:VQ.|�וXo�F��4�LZ*�^*ٕ�L$rw���$���Z�_�qY�pGܳ�a3���+x�.5���8���0����\%N�<�⚺nܐF^�3�;��U�厃�i��M!,���w���P�]{�v�D�;��[��2�Ui��t3���z�si��ʕ�I��E���U��3�����[��3�qً'���4�/k�r�{c���tBLl��>7�[TvxyZ���x��/k:�d�zϮ����^���2S���=Z�P�WB���n�띍#�1�@Kͺ�ʢل�B�oQ���]A��e�Ы3��YIs^M�b�B���s݆�e+��Z�A�W�a3�E��v���	g#V5�L��Y����b����8C�9`Ob7:���]Z�p~���7�j�z�J��)��\�.�͍����g�0�!0�m�W�ol����w>J�P�9]�8�1.m[q�<�S�A����.��I��y�ݵ��F�,K�@��|�O�uw���|u���(�7��3�s�[&��(>��ϧ���/U����kܲ;0L��[�nU���C}���7N�nM'��\st;���Iγ��Xe�U)cں��kP�6<�����$2&i�u��>�+j�,�%n�ꕩ)]�m�Gy�����8`�].S;��RT���,�6U/�w_�2�.�w9$*�z'˹<�#�'u��l�OP����`���z�̜���Y�3e�.��H��Z�xw�9'֙�i(�ïZ��$��&��Եl_N�v�RJ��`f�Vv�O&ܑ�<�E'�����q��+|�j�����N�6?>P}����g���Y	�-X�8�C[ȩP'FJy{9�;�1a�V��^�1.����	� 5&	9�c��4KB�V��|�-#����'Jʼ��^.�����[U+�/��M�����١'U��X]<�M���ݵ&��k�l�V[�v���V�2\�C��1���Ⱦ涝��E���7<���w9tkh�R|[X�xK��x鶯��Q�;dT�sϯf���c�S���߫(hL�9�"v .we_u'�8����}��!\��rw�ޅ`����맥�`��Ed��Z�ZC;�+&�ǒ&��P.�|��U�����=u�F[m�6��S;P=}o*e�mMU}W@�1�Sf��;�D	j����W�2r����6'6��<'p�&���o�S#R�l�s�D�Φ�\{¸>[�{N�:�5�j�����}L���Ϗ�^ͮ<{��ħD����{�X�	6ɱ�j>�*���NՃ:x��x�]�wE��s֣\�0���j�i>�J;2Sz��������B�}@w�v���y�y5w�[�2w^jW3��r�~r�Z��CRt8#�\2��Z�U���c�����,9��*ב��mԵ?*#B���Uk;�K'g���G�R1:�gY�N���v��iT�m�?<��u��^-��ޙ(�9�}/P�v����U�t%[��g�H"��%��wf.���]�e�`_@y���#у)`t�mPͻ�:��%�=���C6�bn�%�[�d�%�DJ;�Aîk�
>���[<'���Q��X���A�������&�d�CY����U[�y9���y�(s�����ʞzw�5�58f�lG��M�u*!t�*ʧ(<�:�n�ͧ�@����4�S/��g}�w��zO\Qk�}YV�*�s]�ԂэO����	�euZd�{Փ��q�v�'�S˄�J��;X4n��S�]�do�*���U«fpq5v�^Yݎ]���~!ζ&�c��@>T��@��Ǖyv���{лl�uu�.׽f�R�P] ��!���%���[��8�ri��9�t�{�ϫ��ݿ]om��2�x,k���=��>�W��7s��g2�#ѵ����'w�b̭��R�����..)�,gx�z�;aĬ=5�[]�\�c�Z>�+�U�R7:Z�u��E [ꋽ�{.QMbUu}Ɇ�J{��;��^:�:ь�P|F �:.v�N�d��I�r�ͼ���bQ�:�B#��P�R��zx� ��t�`��QS�^+�)j԰��4��E�j9�_y�d�
z+̈́�t8"v�{^�æc9e����h,��[�������N8�}r[f]�/}Ƒ{AS��y��W?v�u����Rj�z����׹dq�ͥR.|2��g��wbZ�7����W����.`C�Ԯx0��1,65L�wt�D�v��sn�@ӝ��^��RU����w|Fm����_ҪB��r7��iS���P|�Z��w9�i�7���{��UͶ�#y;�wOY���;�y�������D6����^�K(�c��FW3L��Da���`�So�V`�Npsܢ�Y�d��2��d� ժ�C�pe,�NŮ��7L��y�ԧW5\��bX!��'�ζ�й:��������o3��>��^	Զpu �'�����L��;��WӺ?_A^����Y��o���K�*�iZ!5�BZ�A�A�����oy91�9Oݍ#��γ(]��茦��0G#��cd��3o�����|���o&������`s[[���]�7M퍤2����車���&���6�%F��ۊ�#hæ�n�NN [�.��1�^�A����vV�6�Ύ{�1��y5^��߼��l^�8���R7:Z�Ӷ'�0s�y���^W.{����2�
q��w��ފV/K`��ផ��'d]mL�����2�;-j��T��B86���ꑚ3����Mȹ�7*����	�,�y[D�G/#{��|*Se��z/kI�;�.�����	��[q�k��u�N��ݍ:�;��2��tf
|vE���xs$�R�Z욫���RS8�F�����*KT�Ŋ{g�7�N��v*<ƽ��k�Y��;��\��8x��@�\@�ʾ(�grLq����q�Ǣ_Mu�]<;c͊>c(0Ϻ��Q}�|�ի���;�joa¬O��7[��e=���'�a�<ދ+U���3P�Bn�zx�۽\�� ��\�U+�r��^�e��4��Z0�aED��u�h��Du��i+�\�I>�>�Uu(Bra�:qP{��-��f&2����yjnkT2)��lf��#�@cgvB�d���vtE���T8���*޽���)_�~�W�xƒX�s��^ΔY�ǧF��α�چ��:�����؊�Ȉ�OJ�wb����Tb�m�0�hޯ�Ҝ�*�R��K�>�J�5����J]�?(��k;u-�_{R��k�c �~H���W+��b��#��i�yW�n5��{��uk8�+��,̻ھO)��H1�oV��5u���9�ڨr�~����)��[.�i�-e�5]vþwV��La
*qŻ��9Z5̻�\'wL�$m������`��/5�G�iՌ▔���j��0\y����S���ZuY�ʹ\��ھ%��d���״$^��|�&�Va��)q �=� Y��k���G���}GBO�_���;�P�5<�D�4}1�񎚉}��'�%���t�"}�V�P6{ȹ�)�	��1��W����pH�tbPl�O�	����K��n�vQ����o9���o˶�ѕ ^��d� �S�����꽚�^��Yȋ��:�H��f����������@��0�d֘+�	���o�_ml�E_;�{Ϲ8�)��n����V�eML��8�=�t�G������\ϖ�>i��̦��9�sy��m+';��i�����Pz��g?��>ڰi�`�P*�Ks�6�]QՌ����.K�N��]�s�L�t���v���tMbC�� v|�贏(V�r��ʩ`��ڷ�^�]J�+��d�����93��9S~n��v�e�Q^Yb� dQ�'c'�5X�O�V�7�����z�h����]q~%`+�M��>��~��*j<�T.7N��������]�ZTx�'�&&n��(�z��&�VS}c2����+u�����wJ�L�id�:��̆�u5Њ��$,̦[[�����PA�ѸR���(�v��B������fp�sn�qV���wCW�K�1��+s�Bĵэ��.�}�0:�����J`�����X�D��v������b̺|�|%(2����xk�J�R�u��	�o�V�³�<7Z���җ�=�R�I�9�U��(9c�;���ƨѱ�S|@ʙ[����q`u���(��pٜz���fa�˯6�-�c�=�L��CB�NU�Y"J�h��ኖ����$�ve`�u������'��!��R��mR%���O�1��T�؆��/�y+�a]H��a4։�����+{W�N܍��m��w��WXP��5�Ώ>nM�.�D&n��;"�QSX�F��w�>*j3�֑�%�@�Ҕ�|zs�Ãw(J�z͎;�+�j�o�Yj��]G@S6�`u�,7+�X��9vu-����K��G�G(���r�vJ���gE2�Xֹ��j
T����.�V�W���/k���/���d����U�����Ə+$�#|m��Wf�s,E�gȧk^rVimQ	�5���u8B4n-'o�tE��M���d=�#��*kzC�ҋ���=�2T�vvf����$Urˣ�w�H�my�v�ʴU��X�}�>ܙy���q�0wR!�rm3`[�X6Me\�R|�ᘨ�n�LN��5ջ֬:�M.4v�����r��joO�l5/3z1f�h����Pp������J�e�?H�U諼�=�	��,=����9I�(���֜�69L �a�]�V�QP<�f{��i���VQ4K�(;����<���c���M��ͮ��۹RV���v��8�/���AAp�V�Q���`���̞$!|mӜ%�qi�N����RF॥f�z>cNN1ٵW��ϏG*�QVv���	�J+�	�_aW��S.��VW,����e��m�E���h�1T̝����.�"hs�̩N�w0׷�K�.����9��f�gYQ}����V�/__1Cn�ꐆB�Lw��V��tw>��[�����ă���l�N@]�����к+�(���*�mT[���g�V��t7p��
���ӱR�(�B�ա��#('�;sd�-`��7٭چ��.��$�=�s���}�Y睰ꔊ��a�L"s,�b�N�cBY�NfP�5ϧװ�Ӛ�'������\�gi�{�Ұ,��:6*�9{�������2�RSw�J9pO["�-$�ٷsw�k���.�5)�!�[1d|��'L��w@ₕM�����u�����=v	�,�%U�p1O6,�N����TU(��Kk9��-�e�١b�WP�Ɵ+�����JB��+D�-
���F��U�´P�m(��+Pb֠�l[J[bR�P�Z%`���ȫA�
�X��m�Db��h�P`�
$`��c�EX��-j"�"�EQam
�F(�T(�(�V1k`�*1-�B+R�cETF,�1EQ�T(�� �Q#RU���EbE#Z���U
,(���E���5
�A`�E�dX�b��X����(��B��Q������UH�"2" �� ��DDPUcU�[DH����* ��D`�[X�"0X���E����ePF�DPDD�-*���*���6�D����QE�Q���B��eUDdU[Qb�"
�*�"*����Z�R�#��Q��EUm+dQQD�E[m�AAc
�E(��Z�*2
��"�X�B�vs��R�������̗�%]K���.V%��Cr9}Ɲ�Y������T���|͜���[��#��E
��*���뀝S���!����c�T�]����Y랆E<�u����y�nn�j�>ɐz���9�"��b|Ǭ����i]/M�y`?Y}�	���/v�=�^��2j�В1rq��i�v����Cτ�T��Va�I����)���r��>�3ܖ�J*m[�V��(�}e��
�!��'<���������f�g���bdCcvy��4��fۅ��^^s'gLhrޮ��3k~�&��#܎/<���HǙ���������3$��q�ʗ��}De"�K�;�aG�u�����j��?�F���R����K�33:��"�m3�.��i�~��z��vioxԃ/恄��[�T�nr6/f���\ɐT�q��9v�.�˖XDc�W��[�c�<�FT����/oP�n��ӷȿX�<�ۊ-��w95�qx<�1>�������0�'�]!yJ!�ަ oP�w��]��T]:5�9���C�lu�=�x����R7�����@���fr>_d�i�4,�);Z�%�-ɇ�IK�f�OuB�|�@�{�>ޛy�q�x�Ԙ:jI��J{���;��D�;�[����.�w��w����Y�]*�)Ӝ�N�N�X3غ#Uu���*kx۬�y�lI����W�Y+E�3�l�m�of�0�,'��u��s��~�ͣ��5��u���P؞l��P�H렴n<D�AVL�Ң��mOg1P2�R�mʱ����jdst�u�"�'�M�R���0�iT��"bkc����G���~0�+;��s��x��c�7N����@�0$��ҭO�|����=�NP	�`����=���N߇�;n�;5�W�Sڂ�{������ܢ;K���������U󞂨c��g�[Ha��r�:2{b*�'lݼz�T��ѽ��=*x�~���Ȇ��b#j�|�<�D�ʋ��_-��z3<��y�Gn?���J\X�N��ژ�AǨJ��{���=54/�˫�Ij��ʜ��S�;�������d�<��V��'���X�w�_�Dpn�Qo��o�x�<�U��>*;�lT;V��do�b���	Ƃ�Cj�D�t)U��� �md#�j�X�b&���	�E�r1p{h�VNA����,��:kMW�ĩװ�m�r���ھӋ+lm\[��rM�ćv6R�v�0���\�ܛ�6:��U�U��ˇ\a�*�
�ɞ6V��f۾{ox�%�����+vNi�;�zo,���ή�Z���oY[���`��C�ٰ5���>��ݵ�P����q�U����1�����5\��M��/�At�Ŧv<U�|�r����j�u����&g����
�-H<�fڳ$Cs�l��p�*��z�F����j�9�.��26Hɚ�bH~����i�>/V��:�je�[��������U
H��D5!N2247gb���#Pg!ŝ��(��j4ˡ75�gt���K�#����(q`HAK>�"ի�!N9�*g�N������W��� &F���x���Л��OJ8)�5ʭ�4~�-�YHi����wW����syn�Jb4��>�Zq%��f_�\["���z,F
U���$l7��N�����r�[�1���R��|�.�ݥ2�*Cr:{�"��z�}8�H�M	��Uj�-�>�<J����,��.���w�挿F�V:�}��֌�����Qq�O�;e�Z�!!X�R�>��n*��)t�Yys��NT�'&(QQ-��g-��-v"7�>G�1����Y7[���ٯ��'�h��u���̫�8��w��m��w�Y��J�	�^,-u�ssm�<�0�2����o�y�Z1"Gc�A�ËLю�|���̋��b{=z_:p�ݾm$c�{h\���\Q�X�Z�(!�oH�>p�}oi�κvدM�z7'�}��,c�� �*LE
@�E�hWoo��WQלڬ�� � \�\T^u8��x��l�3=`G1Aub�gb*wFQ��a[yǽ���4|�>Ēv�Xl�/�ܾb[��[�.�d�yב/*v�r�g\>�r�\�Þd�=]0M��A�M"|
/yXY��0C��d�77�F��5h�靮3=�Sm��`�n�b+Upڊ5$¦	�7ȥ���U��."�=��k���nQ�/T��%��R�o�گǘ~L�^s�>/�"9�gS9��Ϳ<3ѽ;&��|��2��,M%���¡�f��a�3���.�gC�{"��q$6c'�J��qlj�yɻs���_d�4��D(�4��d� ���-w�3Ϫ�k����cg�8��:��������!W�`q�c���
Â��OW���X^����_;��dڇ3�{&&�sR�������r!6�}鲎m=)=0}\ϖ����0U楧 ͠�	��z��>��tmօ�s�zK�!��Y��v��07�\|sC�?_r�O�b��1���˅n���b����� �Y����@{���!�rY31�p����ъQjqXn4�IŚ�7[��v�G�n[r�w%S]��%l�1ѕ�~�J$��S�A���&W��Ng���9�켷r�)Ov�K���1�2�A�Qnq�;R��1�8��L@�*8d�f�K7�Ϫy��'���RՎ��d�מDtV�ɝ��ʛn��v��`^$,u���5�=�Ժ�v�=��m�I粪]+�kf8=DH=gE6'X]��*oؑ��a�艽�g5<=��[��������h�Ѽ0���>=���8��WGZ�������!B��uSv3ل���i���>�^DL�	�YGy�i`����*�/�	�^ե��tή,�;�vos�T_H�F #����?#�7�򚬌h�L��|���^��m���:gI��ܞ���k�!��Gy��&��qr�l8�׊w�sg�K�-�6�f����Vm�kw�T
~OtߴMB@S�X���1�~I�C���s8�h'�1zVUI��o$��Jz�c�>��y�}De"�K�;�aGFӯ7�6h�EΆ}PJ3t��Eo�w1V˻���C����¡=�f��Z��ԩ`͇���+��iL���=)E�j�2�]E�l.�;kE7���|3��b�U����Zv�ۗ�=Y�Nђu+�J�w��.��VP	k0q�L�&t��N�u��An۝ma`�mc��N������m���z6,an�gQ�dT �=ʶR�\ҽC.>��`\��1C��/B:��KC�����8	�An�7�iݖ�#��|���HT�r�V���Q���]Z�;�z^�g����(�j�t��ɯ(Go��C�w1}]:�0�R��Cx����EŎ�'ch�J��D�4E9�z>^ɴ���Q�1�5�-��OF�LG��ж>�ylB�h�����=�L���n�IP��e~(�zv�h=�v ��*V��Y��E��=�jWO���jdu�E��\r)b���)q�j�U���%sv�y�3֌���� ^�;B�ye{��T:\{�>�0[�sLG$NH�Jt��9.)�}���������|hKJ��];~�8��Nvk�ڲd���`EgobY�Hc��	@N���J!GP��I�Nz
�u�0\v}����y�d*����c�z����,�oj��d�1�R�Fy�C!i�Ӫs�c&�|�<��~/p>��yHQda�1w^�a����]�g-�o}��&�\ia��^G����hq5�j�bF�u��"�Sp'�|��:��w�o��2���M�]��U�)P<�pʹ���o]��{\ �}�eVq�`��<�%o<X����ٷtH�y,�;�g�_xx�7@��Lh�c�湓�}���>�ͬ���Ϭ��pz��&%dX��HS�U)���q�$q,G��9���"�V�A�>(_�Sk�ѫt�Ǻ��.�گGFྚY���%c�!181�'��T\�c&���$�R�xK��LӬwռ��&��u,�՚���`Ut�~��Ѵ[�9<GLB��v�)��v��;Q������4�ARa��S@�If����E]��ns}�a>ۦ�sn"��Fx1έ��n��ozd��xo2��҃�>Z��瘃4��=�opu]C�l�O^ךO1�Jێx�V�ӈ�wy�tFF�>��4^�lU�h��OON��D��<ue�\��5�؝���0�}�B(��X�l`n��vx>�E+1s�m�;���O�}+-��*���g��>ؠG\����-_�ڏ�S���O_��/���~�Zd���E�i��Q�{啞C��6��d����:���#��đ	x2�`���/~9U�9�\��Y{r���{�Z]�lZ��z�1���'-���6/��Sz�EƗ`��_0i�|��_7w��qwm�-s�s��=�,q�����	�LS��pg���o�k�g����	�?��`��zt�����bMq�f��ȡ�7�<8�<O3V�hO}ɍJa��BU]"�*Ȃ-���H�|6��N���̄'d�1�i�H��{����ϼ����Ϋ�ڑjG@�^��`��O��ɩ��T-W!�r���$���e�K*�;���Z�L�ʇsPm#t�S�;^
�h��
�3�fiP%F��<���*�����kn��	�wE�'!���X�NT؄��QQ-��q� l-�[΃ӗ�-�}Z������6_*Ȼ�\�^�� ���vhi�+�������D�*LE�״�(�wU:��YaT01@��� \��qP}xˎԫ�贌"�[�Q�K@��t���f�ן�y�²���-�K^5@ۖ���h�}���)V�K�Y/�t<�~}X�\���pWUV�ܗe��q@k��.S�4�=��U?	�B��^V"��]�C��dL7;ν4�.�*U���>�z�8\�'��q[ d5jK�S�x� wKCH�8������_����{�~p�6�\���~�U�
{���揢���/�t�S���:ڬ��AX/�/w#D[T�;Q}6QB�;�mq���gX�|s�`�i��Eʒ���-EW�7z38?�4靇�=nE1�v�U9��
�+l�c����I��11�*咩�ݩϣ�c�̦^��BO8�`
�h�V�����A�}&���WE)�W�{}�+�����{"���>l�O��=r��JMqs.����ܩ~�ɺ���J��)''a7��]���k��g&�k���ԩV!i$�׌:�N5��P��7*M0�iႽ�OV09�xf��٧MԞ/������ig{��ݍU��r��%5����(B"m���G��B�JOL�g�h|�QQIWP��f�p�sU�����U�x�[>$�o>ϊ�z��g?����j����-הŕ�Y(�Co������y%K
o�tclb.d7J-˗YR�1�5�u�`2b DJ�0%�m�c��헗:��G9R0��d�ׁ�󝥆�Κ�y�W�r�*/\g��[��.�Vu�rɞ`XՇ�=�yN\�K��'ܩ�Zɺ�J�Uyr��ޙ�i����s�f�w�?b��qjX����ظ�a_��i�������V�s�;aI���n�k6�����>�艟{�}�Q�^�$����� ,��p�E�>�;����~/N�JI�솫X��	���e�qE՗T�ՙ�fd��p0�,�V��Ot~���;{���9
�w�����b=ݒ�w�gK��{�a�xS��eMx�:av���X˫��p��9i���$�7)ףv�ݺ�Ã�$�+Ngfkhm)��l���� CLੲ�ĉA�,~u���)�a�19z6n+χ�6�QH���zǯ�o���A�|�W����X��e��|�ھY�zWj�$�4Ѿ]}iomץ���+*��0�Hw�P@I�ٿ9���`5Q��
�5T�G��]�I�C����\i��^��E{$�b��N�[�4Z"ЮHa�!�9Y�����'NP\׆F2/���i���SdlL{�zsc�l;�ő�;܍_-͇z.N�;7l���J�S��a��7����V�#i��] *q�;��U+f�����},绥�q8��__{D`�b�6Q��>������;���_g=	,�[�c�2X�H@t�F�TN�6�T�{8�B!�����1@��m����1괮�w�0�Bd�8���ި���uC�`k"ݧa���b�UCbz۵|�
,ETY\���4�J���9������#��`�گU�c����RC�
�Ac۟�9�$ I?���$�p	!I��$�	%�$ I?�B��$ I?���$��IO�$ I?���$�p$�	'�H@�r��$�$�	'�B���$ I?�B���$ I?�B���$ I?���$�	!I���e5��I��� ?�s2}p$s�=�uM@�-0HA � i��J"�)RU%J�%"��AAR�)*�H�ZHR�HU@��m�$�Q �P��%i�[&�[k-��l�Vɱ+�r*�֢̣)�$���6Ƙ��Zj
�ֲ�͕����3Q�@�d�ɖ2Shm��6�pr�z)��4`J+fUJRB(�i���ښ�kj�م�Q��+Y+V,il��R��I����V��elժVm�M�B
���l�*��   a|��U�t�k�z��f�D�^���:��ޝ�@j�wVqz��j�a4��a�swi[�en*������{:�mww�.<�M*����]�V�]�eD����z�]4A���vH�    �y����-�og���{f�Y�7{N��f�5�{�޽e��2�]ꈑ�:��^�)���l��9������ަ��w0�O]��J�[cs����ƹ�9�=��Ҫ��;�+j-��4���   ;�_nS��׷����47��\��c��[cVi�w^�l�dո9s4�[�/x��( QE��:���PQ�����}�����:4h�E>�(� (����m���o���%4i&�ʞ   �� >�>�QE�qѠ(��(�}z��EQH=�iV}(kZ83�kl�  ۗ�x�e�7n(oC7e
+��3�h��5=sJэ%-�53���  �>�Tܾm� ���%��4�j��
��2��=m�w�(z��3��״��U����-��5M��k��z�E�M���ڶ�+b��E4��  ����A�7zz��5��smֺ�w��zP��c�ٞ�r��fkH�h�P�G��)��j��v2]��)�vN��:]^�ٶ֌�Iݨ�m�[FC|  ����m��vٸwvh
��K��Q���w&m�q�qú���
�iѮ�{�ާ�ԥݻ�z��[m����IK��`뎤V��ٺ��w+v檞�U[���g����i� 3̟T6j���[���*)޶����p[n���JY�;�y�y�N۝m��w������˹ţ����{�ٕ�]��=���eE�뽭+lW�����FKMb�,�F-a��Z|  ۯ�>��j���]�*�m�=�A��Dҹ����:�뽛ݍ��mv��*�C�^�z٠�N����֪vi%�{[�]ƴ�֨�R)-�N�EG�j�Q�Z�	h5h���  =���{��αEMo<���j������zU[T�״aQ�;�Wod�Y��:v�46�wi����MKm�m��wj��ʻ��=mm$���� eIT� ��F�Oh�JRTa0���l����  E?�P����4��U@ R@�UJz@A�<S��#��������٭�����Y��Ot5�����޻��ܻ�DTA^���?���TA_D�W��TA_�"�
¢���?����+GY�?�_�}�����Hi�e��nb�Lr��yd7ol�A5�Z�LT��6i�*���v���:ۂ��٥)l��u���l}{SU�t� !��S�P�OH�M�N=�֒�;V�6��[�N�;Ŷ��GaS.���ְv�ß<P-Rˎ5v��Up�S++-e�/K1Ӂ�,�#a��&��h��D��:�hKsr:����af�=?m�Z�>L�~�Ya��U�B��z±�1�rܺ�[��sn�������j̠
��:����gٮ3�4 �8z6$�������i�����j��u.���;Rk!"bjl�����b:�}41�[ �0��i3@m䔃�CF�N+�Gʥ`��!�H@���Me�:H���i�ST�[΢-V%E$���h��-��kPv�ٻW4V�`���	����7,�Uȅav�J��Нf�!Y�+��M�����\�J�.��;[�������H�ݶ(�v�5
O�[�%[�Sn����O�͐���Gz��^�pQJ&C�Ad�'�Xտ���i �K����%:�:�9yCw��ڊ��8ӳn,HF��7��e�ecv��t�nZ�R�{J�J%j�n�K(ݍG4x5��CkZ��QLa��QXoo5)e��l�����1�(�M�B�u�=��È�Y�&�M��9t�R^����5O�M�eM�j�@e�Y^ڸ6�M�	���P+q������܋�y�!��ᙪ@DWH�O�J�z�o>{�+F�j�
�(�x�s\m免��t�v~jӆf76���v�JP�';5D�{nJ;���с3W����QK9ɗ5��GP��*\xӨ.��?:󳷡*t�2S�f�\ȯ)���윰�k��m��e!����)軫��P*�D�J�`lXtd͐��v�[O7tj���}(U��2�X��@�w�cUZ�SP��2�LCtS8V�{5���hM-��34+�vt�e�÷lV�&ᡏ��)0����N7��hn��B�)�m
Oߥ;*���M�A^8��ӌ\�u۫C^5�*�m*�8��u�6)��tZ�E��Ǚ�@�b[,ؾ�t���u��܂�u:�!)��Y��z���51��S���SA�W �s]hĎ��m�&�5�G�1VЌ�N�kź�)P��Qd+�1�c�6�
F�H[��階dbt�:{nݹf��vEz�dw&�P^<���Y��@A���L0������VE�$�{�����Yx6B ���tիό��[�F���vJ	f��	�m�S�M�y���+5t�(��ӛA(��w�k��]ul�fȗ��ʐ�J^��V����T#i�x�ܥ��z�b�Zh�cp�T+-H1+�d����+fc���&��t|�܁��7)����ܲ�k���t������M����j����݄m�m��jw��w=y��O R�h�{�Ch^mD3J+�)аi��\�+NV����wQM��v�F�K{��r7�"G$�#n��+!m�gv�V[*?��Q��[#�X��V��k���y�e�]�8�"-V�>�g u,>���m��	����.�8<��F�ְ�TX�d�x�_�"tZ���k�X)�����n��"�s ��wp��ZE���0��I��^�u�	:ȳQ·r4Jl�ݛ��wI�ި���8�!�YH"�1<�u�J�sB�8���T��V��[5�(8��l]�D'�Q��2�˔�Y�dj�������7xē	����4Ey��ъ=���RUϕ/C@�	7PC��k�7V5����)PR�i��[�m�Sc�j3�%v%��!�^��L��Z�Y3r�U�NGX���V)�MJ��'�uV'���d5Y&�n�P��Fާ���}�U�ò��t�*���1m,�2[��6���*h��Cv�۵4J��XJgJc+k4cH��־�Ph)��U�-��E�9Ct/�!�Y��ʆ�I�r腖Tv�Rݬ�8�#w�[��v'��P�/`Nl�h3yVP��N wXT����m1�J����L"ū�YL��&��Qc8b���ibB�mֳ[��"�m�x�ci;I��!�l��4l�sS0�]�4��z,MAs��޲#rЭq����!��(@2��H�*en	����
^�Q/�W�S',�T�(l���md�Y2V}1
e,�[$�M�Z��/S��-�3�K�������eh�t�%�\n�;YH�5eN��U�¦�)��#פ⛇C�//o.X50둊a��@�;D���*9�ܠ��k��Ma9�����Y�X��FMm�le"+h�PɎ;� �lGC���L���
 ��4�i2�4Mx���V:+i�Mo�Ь��rd�pSՉGW�k5����1���6]Ҙ�a��5�Q�V���륶��Ia��.E+�U�N-U���(�{��]'"8s"��
��WlnU�`�f͒�V�ă�,�V<:�&�hA��r��c��ۓ(|
),72����`*�t/[T�V�2:�om\j�+.��^Ղ�T��U/kW�AQ��Xz^�Ks�Ʒ��d���6t�FMn���G�7�K3m4K�B�m���k�x��	�
��7kic�t��4Xմ���;/ZV�I�«�B�h�E�w"�˒���SfcVwE��3�!p3��`%�X�,[��fh֡[i5*(����͉��m�����%��T��Ѻν��v�k�HO�W�-���̔�6��ֲӑPz�F�]Q��m�Mh'fL{�V�����\X�����}e]�s1Ĳ˕��5w��4�^:�7���3i�Yj�q����Ɗ�*ub)�Ĉ=�rk�!ڻ�u�Z�6�8������5�h��T��tmXE(Z7�-�ݑ�)7I��m�f�=O-G.867
oF��1h@i�-5�]��S�� 9�i�i՜�����*զ���E=��x�K��N:{��;X�cx���٩O$�h1�Ԧj�.�N���oIg
�˸a�nԆ�o
4�ƈ���Z@��cg!*MvMK���Ғ��-,e�����sI�X��j���f�N���݅@����.������;�[Ѭ`�aKj�݋��r��k�F&�
'1jh'i�̻`�au�����*++�v�]+�G�I� 	:�ˬsM뼦/u��Փh'�y�0�яc̋[u*;�Vܭ�u�[-�f��5�n1��͡bR��@d�6钸|u�&�K�LCD�(ݡ�����)T'+-�2
�J�v�Ŗ6��'Y����-]�ʦ����hD�)�;k��YgD,}u�� S"}�qds�5��e�e���: m��2ڰ�x!.` hVe�m�����SF,0Vn�ܒ��-�룗yHh�iM�+uO���廹��J�l�V	X�Z��A�{>�DL��/&)7�(����
3)G�*�]�IQ�V�߳B�J�\7�ʼ@���$c"�v���yF�3a�f����1'Y������[V�e��j\���#$�D��Uz.���¬�DPYZ�+�5gU͹�c��@B<y��ՊP�(&�P)ZU7b����n��Bi�a�R�C�+�,\�O�"&�����*����̴��+dCjjN�L�,�K��b�CrA[e�,] $;%�
�ژ-̺�ܙ�F�$�N+�j���zlZY�
6����"��jUظP,��L�7Z�y��`�u�H���i&.�6�L	��
���a�ϝ����ӯ&���hD�t#��o3Sl�ף3��(0Y��U�7C���r*8�M�_�ee)�V��@r��%�J�m����U�J��e��L&ʗ�q�QT�׭hH�O.�OrkU�K��Ų��d[�J��_�] ��Y5��P�Eƃ7�wL]��;��0�Jl���A�m
���[���'�IK	+M]���7V4��ɺ*�1��$�/[*��PX���
�3���$h[����n�p�JۦOʊ���*y��X����n�I3�.��шe
����M,�	aK����)�aP���h�b�����Sv�t���
����Cf^Lt(�$�n��uk�6�B�*�+6��2�t�fLs$�bZ�I�K~��v��Ցu�R3[N�!ZPK�)ۤ�P��Ti�i��
���%n�fI�G�-S�v�^7����N�O0vg[:/a��!���bf�1��+7S�hF����`ۋ#�� -��$i6S�˛XM�85j��{����-'`ti���g��b���nC�[hhd� l^cO�D-�Z�LB0hfTu�Z��:֪��SAe���le��4��VYA^kj^�R���iʽ�V�Ij�ˈf�;�v�oS)��M�ѶJ	�)�*2=��^Â��M�n�3*�+�6��*��H�KJ�$Hu�f� f�C�����+�u�+K����U�؛q��ŻC����䧺рfQne*�W3F��Qk]fF�k}���CyWfw6]1��ЏO�&(|��l��[8��T6U���f�Z��eҔ4��KiH-a�Y��i��2���:|����>B�K7�S��& ��^��;���z�F�ǗZ�o)�����Zo]��L�j�"ʆ�����."]��YGV$J' I�tڭ�@�n��Q0~�V�z����P�"�h�[�]-Ǡ�R�j�Y�- ,ekx� �l��T�и��CM�x�U,]��tB ��+M�kn�ٌ����eMP(M�+o����xƷ�o�u�VW�vd�iدo't�웩�'�F^��=����Ϋ��᭫9�V^F������`K��D����SG�]��9�Zt�Nn�@��E�d	r���jy+�Ye7���M�����I�0�D9�mh&�;[BH�F"%Qj8�Ri�~��4�u*  vS��Ë:Эf�əOtJą"�J6��-n-����i����k!e���H�)J1	{�]^�a��w[W�GC{�SL�OuR��ߥ����%e�E��; ��g0�Q2йO<���0�z&��A焘�7Z�Ap�Av�q�H�x�U�mͬkq=�4��¤H؂�M�:.zL�p��<r�5-n�f�)۳�B��'��`�
��A�������o2m,l1�/m����A�hh��J�ڊnV�{.쐊)��KT&m��9���6��M�z�=�h��f1�޻�n���1Yօ����QS�U���S��[+-�0"�-�deMqb��i�+,��Q
wyY���dUa��z���uz����QȮ	dUڲM���N�t-S�V�Z�P�!���������5� 4�D��A9O
��N�)�l�0�Ӗ	��He:?W��s7^��#������BQ�(�F�y&�2�+TyN\	���`����w��&ӡ�%f�T�B(᫤�DU���l;s@w�A�J��*{�iM�P��!�;Ǝ��H!{.�j:��y.ؔPYwN�x�k[8��%9%�J$	����#j�������uf�Z2Ȭ�2 ��M��k�#/i{{�Y���&^4���SF4�P,Z��DT�%�hڦ�іJW2�8֧��z�Rʃ
Mn�h�I��-)V6�SXq���oTGe�I�Q�Uj;$h�W0֦c̳y���D��j�8�7)��1�ڇt�w��.�7h�{o�	J}�n�k��a5�F��2�&���a�^Y� ő����B��%dL�����&�֥�l�h<����f��ki��$�j�)P��n����m�TwB�jP�P7���Y��3Z�A���Xu��A��+v��l��Ť6=���p�5[��J��v��e-)քB͵$$Z��4s&�W�U�+,�m6-ܕ46Yŵ�J���^�B���52�X�[)kY���7)���sM+63jģDh����I1��u�6�ҫ9e��^�iR9���MމY	
l�B�Yusd4��f��DY��
�p�����ѯN|�+V%�D���y���U�V�j�X����ɚ�e����ARUY�%^=�F+z��~7��k'B�CS
(��|_.��DH�z�bFnW"�et`��F�-J�6���(�4-H���h݋Q���U��el��	�e)E�E9r>aıageh���N��Ud�����A�sr�����-��/��tڣ�V4�{O��f�rHN'�j�I�m��x�S�
k�ʍ����ڀ)x6 K�1���ǂ��nҼ���(eZ�4�`lͤ�fn����zh���?J��js�;͗u�^-1(Ȑ���WH��xb,�7j
��f��^lzΌD�.����$����M�YYX�$P�G{D�j\7���Q	3h^c%e�9A&bxsE��q	c`M�'帴�C4K�k�d�(��tӭ8��<��i��n����*Ʀ��6��W45[�~!m��e�����,m$��WW�ⶦGm�Fռ��0�y-Җ�
ø��ŮL����ߌ�r��,�q1f7f߭�M�0��R*���MUÀe�V��Y�x+.�Y)Ǵ*[�l�-J����Y��%��4���&��>։�5�-l٢�2�w��T�ϤVr2 40��Ô���;Z�����ހ[*�`�2���aM�2�轣CTn�kEf�ފ�ǘ,-��W��'�؜�O:`�Mu�E�6�w�;�*8^���[��Lݳ��k��H����b�)\�ް�����t��-NF�;:/v�h7�n���7.�O5̖��2���}J
�u-�y)�,m��@KEntެ��𣏕�9��y�leu%�^M��p��1��L��Y$j�^���8��KHٶ�)���T}�r�PlBw�`�\ZpCj=�����6���,+ۥЃ;r�Xp&X��v�,������uck:��b��p�Ma{��(E�}����)�fn��imB�{������W3�'KIJgyWq���H(��|�����a�S����J:2m�be�v���R`��7���VQ���J�m�3cҬ�W��1��;�;�%@�d�s��'|~7�D�b�a��b�$=�8���|bS�;gx�0�q�Dn��2���!ڗ��"�m���5��Ӷ��(+��6��]b�;� ��r:j���eKM�;��WM�j�?�k�7\΃ᮣ=]�wL7�7`��|��n�y(m�=����$��lb��+���:!��;[��� \���B���(�1FD�U�Ƭ`"�1V�	�q*1e]�-�h��k���_�B����]]{97cU,q���M,��n>B�v���2���ڮ����w8�4J��	S��Uv���=����0�+�)K���"��\���Y��yu�r�e_s҂`�k��_�4�^o�5(��mcu��-��{�mۢ��ș�VY�\��DN��1t4��I QtVvV��ޔ���b4�(^ǳgeII�]�3;Q���/h��>"�*�ʅT�^C&�i\���Z�7ݏ�*��Kc!�Zc볦dY�47(�OڍՀt�.�)�0،�������u�R�7{�139L���I;ЌV����c+�����8I�%������r�%�h�Ə]� +@rg�]/|����_*<�.�)_oAxp��33�GT�g��&k#��t�E���\�wj�)w�m�N��=��$'g[x�<��t.�e^�C�`Kon�Q!7��G1sN����B��0��wl+n_^k|��
��Zg�^���QN���E}��c���ZX4na%��D�ݝ��>}�g
�ZCgG�%�ԝY[f�j���u�K�p9E\����G�{��h�?E�u_Z2�l�Wj��,{�JY[a�a�a.wf�nV��~���������ǅ���ڥ���mrw�j���9��WaQB������D�b��H�u�����e��[�v�vn��ê8X��6h��e��bܰ��9Cw�8�U�n����̋� h��GӅ=�eɐ9��-Qo!����x�����y��˰��b�f�;(W�3
�۸���V�wf�ޓ��O��v����C�"�t(`�޺�Xq�@�s�qn�j�΅�]F���̨��e<�������-}nI�h.у_�[������^H�V�;��:��b�RK��g->mC�B��Xn��UU�乩�	,�廻���J��>��{|��F��"�Hy��|DW�*�R��jaE7g
=��
�н}��Ak�Qs�>��m�rx��w�l�=�I�F�@�I-�}}O1��fq-�WN���5��qeem�!�Q[yD�hQ]{���bd��i�����+� ��ӥ���dD:x�y�2�wvc��*��V�\6�+�2��
������v2���jZm[�Ǩ�|*]w�hSw6�����VIs��ʤ{_�KUk(s-k�6�(��ms�Dy��]|���H��eT��L*�J�I�q�oUe�?���s�pK��*9O>3�����t�6h����8{���j���2�)7�B���D�ˉ5�x^�� ..����؜մ*舗G1�Ԃ&��9���6�"k�4�+�XtVVY{׎�T6�M�GZm�9{��s����Hi%|�=(�}v���ܵ-�宼��-�Oy^+\�e�5qRkc���#8l��.뻳�u��b���`S�v��I(�!�ae���՜[���V5��%��W?��z5R�h��x�D�꾙;6o<[SxY����i�_p�rW*�̨��Q����d;��3�.��ǫ1���r�[Ɉ=��\���ӛZ=��c�X��K%;�.�[|4#�x����w��]MMu��3���Uި�I҅"���e�n�7wW��򛪧s�G!U�a	�^E��}�wk�!{�]��`7���gn�������}|�%�Z�J]'�r7��fu.���?s!���e�]�wR��m�ҍ]�.�8y����J>!�i�r�!���mo�'LkҰ�Bc��mG���$2J�Ʉ�l����?M+��ڝ�i�B��r7�� +�n�S����7��F����ˈ��^�8�,�,����9�0��S��%�J�އ!T�͎�lo��&��_�������6��d,��.�n_dP��ZW�$�|F�VRdg.��Ȫ�V���@��^;�-\VAC^��H<.������ڃ7����e��^�����:'-�@�g�� |%����e�w��X�ǜ���<Ž�."���ܴ/�sk�9{L��"�!4i;+���oph���LH��ałQ�V:�t�紃�_r�ו}/�EV^k�R�Tp��������r�n�9ޞz�!�%0��J���DsY������r6й�wYuwѧm(u�ͷX:� ���w����Z+�O�1Lb}��%`uo��N�u��Y{�R����M��s���*�G�v�}{O������2�<��\s�u�g��v-ls̐�z���׊���':O�øI�=C��r{F�Ygf��X�J*~~��g@��5�`�vd=���d�؆��)F+l�'"�6��\��
��vS�0�T���h�Ԃ�OX@��5\�ͷ�cg����i�y����+NPK]Zu�AyJ�:ॸ���yH�4L��F�ki*��%D��8- z�:�,Õ���c�e�_&0Ӝr�/m��'��}�չ��rwH��Att-��ḍ�-���
ΒJt�%»,�p�^��N�t2��9s���+qJ�W�芦�AAJ�+�g���ܟZ�9��=#\
����^���i�s���
����eQ��HJX�-�4��ە�5�������RE�;�h�hs�T�x��'��7وA@K���w���uwVՄ(]u�Ď�b�u%]]>������so�8"�j�W�,@"Fa/q�-�*�6)���ΑϹ�N_�y6X� ��������*Z
��Ǝ�ҩ�%�:l�q�F]�!�ʾ��s9���Vþэv�r�=Z�����f�̓�<�7�+)S*'{hȭC%Z�&��%���ͽq�T����U"%�J�c����Ϭ;���ȱ��X��;�J�h7N��xI��=�+�7mx�X�V��f�8�8�ηw�n�d�;v[ãa�1d�q��{�l���.dc��r8m��e�j;@ab��4��h��l�q��t�LyI�5">�]-��FĨ�u���2Q��&�GPQ��jt��ډWGyy��WC�6޸K��ԅ^ҏN%�;y{���3�P{���L7��Z&�h ��O_K��υ�I�Z�ǘ�՜\T^G@Ԃm��ÐXJo*%F�=θ�'&otkN�TqY��޽|��x+�K��y�5�ࡧ���s�8ߘ��6i5�X �3�ժ��M���/��ĺPh��ю�X�c�fW-
ﷶ�h��j(,zC�4�$�L
�-1575\�yV�-ɰIS�5u��=����.��!��s��׋uwU�TN��Pv���Γ��)JAd��=��Wj,�Ν�� -s�1U� �o,�� w6�n"-�zy�oqr/)ƹ�׻]��=��R�� ����y�vr��d�Z�;v]�)�6c�߱"-;"�=�R��DR��H��)
���6�i�Fu�] ��K2ѝHg��ݚ�If�v�gt�rG���]Cagb�98t���Ӻ^ �e�U���آ��dG#��5�G��!þ�k�wtK��9_ G:�]f*x��4n�,�Z�ITZ�	�k@loc�j*�m���b��Ytׂ�	E t�yX�8�{�v��뼭�R��J��ܾ�������(��Lj�����Cwtj3J�/q�[8����e=6���շ�x���n�.�thb��U,����.��.�SZ�1�i�ǉ}0��U�IÔ3,쾺�A��7�����r
���TF�:�:.V��V�����i�VpU6��*ozf��6Mf}6��z��m���36][��{D��pENh#�,9gpo��{ -��Y��D�]l�P\>�v���M�M�B��k�]aWMK{^��(�/fv�*of�
�6�ƅ�������*�s0[I�kuI��/h��Mۭ�h��Vou���s�xcJ�\�X��╚��W�M9���γ���T��wWm��S�f����ڮ��9H����qd�o	��T�pO*�ח`�\Pw��̫M�ſn,pD�Y��&jpkyyVru]"�^`I��_7�9��SZ3��˄G�Ԃ�I8j��~E{%��P7*2�p'j�=�޻��_A��A�Wڰa5-~ꦇ�ټZ��"��B��2:�WN��,��qի�ݬҕ�֍,�A^������6m���L�i��7"֮ή`���j�lF��F3�K: �'���-݁�^�1�U�O��k�(���=�.�W΢R�Y�t��o
즩���hC��ʎV0;a-�����u�h�O+v��,r�`��up��;p_d��ӗ�66�m7�0���[u�:�36WU��W��FÜ�|���Wl��v�\��y�L�z;���{�wf9d��+�@��U��V:־ywk�F�F�ֲ����H�	ؠMm�=��`�Uͮ�<)3��N*[���e<�;��Q�*U��व���5�Nf"����Tj�eZ�'N¡Az��m�K�2�\	U,��m��&B�ޣ�@���t�;���+����V��b����׹ĩ����ꚢ����o�_K�M��.�,\����	����y�jͱ.��?i��<�s��5�׍�u�v��;s,u�Ц}�+�W{�5֗J��c��]K�+ѡ*Y�D�}L�E˂�����Rl�����BF�� -eIZh_Eՙ��7��I�9f�,2ɾBJx+�%��DN�nQ��c�r�W\�k��Nʧ]��x����ʡt1��͏?zf��J��C�����s�J7�F�i>o}v�}X��u�������ST��g��'�-]��u�7�"�ዮ�S^B�X��^]-�d�97̈́35����m^�i�p�op�N�ԭ�e���gSݢtE�P�Z��Ėe<�Ǐq�'e7 ��k��u��]㉍�BeK�ղj��pӇ�3*L�;�N�K�/��8��*��w�KC9gd��]�,mmA|aY���3�y�-�8�P��k5/6sD���}��N+�Gz�����!\9ge�L��r�e�[v�R΢�T�go�!���˫�w�z�U�����r�8�(�?pD�FJL�̒�ũh`�AY��T��n
O/�R��%e�[+�j9����ʺ���e��w;	k��q6#��.�K�V�������묳ݩ9-���}�g�`r::%H-t{WP�
`KT�P��+�e����$j�
� 3��:]�թ_	��Ӻ�>�V#�2��6�Q��QR}���뮶���:��҂���Ics�]��#x��"妬8�F�xc���L��w{�n���1�#����0��B�վ��'9n�G0�ʾI�H
Y0gpW�ge<��3J�U�^蔊3��K����N
����9�\��L�?6�cG��A��%�����u�9W��`��r�L+����t������i+�V0���������b0�[K=C�.�$��9:e\a.��퐢�ѹ��h�e���s\��~2�;�!��jn28��7�f���'��Lʄ�S���M.W�kx;�k��`Ņyk���e��@h�m�wmּ�����gn9ϵ�;���8��|r)V�u+�@��96 �}��2����HCM�b�l�ʶ��ݝ�z�]C�E�}�;Y@�C�'2��8i:�SN��f11�X�.��:��W���ۇ�/��^ջ�t�Ju6��Y�"����1Tih�d�MK�#\°��]�=K���9lV�4�Dϻ3i�*�
\�i��ʓ��Z�
��� �XCaV����T{|$�(jqV��K���۱b�����m����ｙD���0����4{b�Vj�Y�2����1��\Zmݢ�lv^���>�Gg���Ɏ�2��X��2�Ď]s��B��ˏ���FƖ|j��QF�Rf�1�Vp�]5��YZ��%���(�pgmu>5Əm�>#H�rr�u���H�V89Ƀx�:)&o\����l�}���Ps!�h���Ы��۾;ۤ<������,�xo�j�;ݕ���[p,6��8�S�jĬ��
�z��9��u%��_iZ�A;!{�}��ol�R�6�qsVRv�����s�f�eA��[s*wehw����u^ZאZ�����v��v�fE����'��X��j�ty{��;u����wn��UT&9�h}�x�͵[7Wv�1�=}��i2�6�h���g�л����8o��2Â�fA���S����H��%w�ȸ��(��.�3�N�5n$�����+:�.PVf�*�9/��{��"* ������g�k��5����7��r�����
Gy9<�D��wյiZk^NBJDa�m���s���!y(U�7)��f�wC9^���!O�b��]1S��C�#�ڠ*h ��̳����`��*`Y��m�_�o[���D{%&�U�)�Բ�i��۠iml�ŵ��۷����I���3kL��n\�m�w|��i35�����6�^6�VQi���&�59Vf��ՙH��	r�lǴ4oC�
G�A;��}G�ڦY9�X�Q���|:J,���Hr�v�T�ୌ��L�´M!�=׺�$���خ�`]�x���2D(�$����Ӗ*
��N�"4f� y)YtՈM�ą��R�.5cH��n�����nQ����b��+�S[svF�a姪F�rqR;p>�O��e�<T�Du7���׳�G��61v7E'M�1� -�@P�+�f�t.��Gm�«\���z/�"�ִ�m�o\r��\�e�ͦ���v}.ȃk�Y��e'B���+����aS��/���Ƈ� �w��� $WTrPi�w��ޞWV���'�t�.��Ku E�pқ�ݴ����HѮ��b}h�'��mPvq���Bەv�����������Ajh�ƈ�R���d
�2�$�����
�����J-�Җ	63�4����5�iU��=۝9� ���hH@�G"
����>\�ݢ�Lf_cbc9O_ت�'2�(N/�������ۻ�l�U6]i|�Yj��l|�
�������7�Ӧ�*��L@�`�$�G(�8��u��3��I��v��F�m�1�U�u7�nBv�BVEI�T]��5ǯ�G� ��]�V���9fW6�q�����i[�:Yږ���v��N87"˥�R#D��D�Q�f�ʏa�Ͳ��4p�8�o��,�V��,lm�i��ޒ�if���ME�˦:vw��������{ܬj��`(���D�ٱ�I�>Fe��N�]�!��6�Ҕbx���RZ�mn}/~�RJ!-^,�p�J�N-�t,>e^���f��L�:���A���!�Z�@\�H���4_�������q�Zk�4�Ts9�T�gC�k�O9�w0e��;�����"���/�*\]N�G�,�V�|&]��έ�'8f�&{iYt����-6�ٹF뵯��n��5�o��YKF|��է:Ӯ��V�p�ʆ��Ԕ1k6��Vuj,"��14SJ�����s��s�е�ON��l"�K,]ki����*Z��aar�:+=�z�+3p:[�Hx�h�2ګ�(��z��坪��k5�
�2E�ѻ9����-�G�㮹�--��}ݡ-���KЎ����{Zq-���.�b6J���R����/%����mi���7I��0�\_h���X7
p9���l�k(?���EU�ɹ��-�j��k�.�p��]�:��2Һ꒠�u�ڕ�J���;�^�mD�q�U�\���©����񧼹��J�y�RV+���Q���T��R`�U�CKG�5��@���|�އM[EY�{x"3]�0V��⍲�{���6XnWH%�ެv4Ac>��hBXG
tVn�qy���C�*u��*o���--pٺ�,$ot. :*�)��e#qc��e�368���3T�g��QA,
�\�4G�RFec̄d��.7�1��A4K٪5�:���K[ =.p��#/5v���P�K
�-4Խ�R�R3)���^�Sg>���E}ă C��敗}@u0���x:����d %�7)ս�9L�}R�b��쑭���f�x�.�1V�4��MԵXfq�w�r$�N�H④S)`���ϫ�l+�W_;�Х�Q���e������Tݛw�e���-U�:�f��0C�c��-��!�e�Vt�]Yע�M�TX�.b����ҽ��WbC 
RT�ym��C��a�� �tа]�/M�U�+Bw`w|/���J; �M�vX-.yV!�o��&�p��r]
}&�֘�	�#m�;��*��!�M=�-�-��ͱ(qm��Ћ�W��R����䫨1h4VXn=�Jbv�~��%V �\H�6")���!L����^�nܲ�$��Ҡ�x��Ɓ��J2p6X�%�*+Y�-[��(��>��p��N�˗��9Mb��<�R�y@���R���iڳ��a����L�J�4�1\��H��
׽���un�nJd-R�Od\�=�m�X//��S�1]�[��5ۺ���X��B�I�%��R55�m�3�JY��͐	��-�����a�;H:F�n��'�Xͮƶ�2�8^P<'m̹L!l�C�ӑ���2:N�-�(��΀i"���;�������O����[�)_d�V��;+^�޼{,F���0|�$��II[���Ò���r,^�Cu���M���p�T�:+�V��� �y�N-�rl���2U� �B\��.�N�J�����l�Rw�)fށ�]�N����-!�]}�u�[Jv�Te ��]ku���_[\�C���@�Yɩ�xg��]s���"���#���j�l�j��-#"��wI3�wr�{��[��֯%�)���9�g$ǘ��!#�n�<����-%�T����ԩ[w�m�w3v%�GZc4��8��+��z��2�鎊�j_���6�޼�(�"���yE���0���.�71�P[��L�2����$9�lLE��)'r�<7q���|H0஼O+�r��H���'(}�������d�tԨ������4`��6� �>�v@��mWȲ���58sі�mY|�k,n�ŵ��[���d�U��m܂5�;�s&��^�Ӣ�F�cs}jTᇠ#��LI�w3��7v���uN�v>��gq�o�� ���/�z��3�ӆ�U�b��=H�,�l�L^�����5*�D�-���n3�pږVc��b4ƍ�&����*G�V�w`0��u��#�����Fu��C��_|ѭ���k��(����xSd�V�y'E����0>���⛺�j�S��_�4�m	+G�$�]���b��CR�i�M�;��4�WAn�CWMu��ʰ�{rG��+ww)��y�*s0��[U*����&�6N1.KO���D�7�g=�ǋe�+�入6n���Dz�oN]�J�7P�|@=m��JV���l�e`/p�:�@�voTej���}0�)��0xR�e]��G/`��#��,�	G5c����Qԯ��E}Aչ�����򻎔�w	v�P�T�Q������ڊ��=��9��#�
���ۥ�ؘ�u��i���hoڶݡw[E�v�>���(�Ie�O.
}StJ�C��-D��]��K��6*�X�v���u�8�-�A��L�('%m?�/�]m���q6�7�*+�ouIf}mV���jܾ(��ör��OH��W&�/�Tr�|-���!�)�ּV�q�4��]AL4�X��c!�ePTw1c�#~qe�ԩ����Leݲ�c�M�D>k�N���r\�nK<:��,7p�u&�����=����V��*@���1����N-ᥦ\�6�$d|�
q����'H��45�e> �v��L8�V)[�p5��_Q*O��RSH���J@n��[�,��;���s�q�jΦ9;<�6�9���E��p��%N�����M[J��c�����2��G�w\���\��h�렎AeG]rWZwzn���ؚƙ�t��7|#��9fh�����:+�J�l��;��u)����S��υJ.��v%(����Q��a���[�ՙ���´��j�;P���S޾��d��Va��t�iS�㋸i���6�P.��������W��"I�o9b����-g�R����v�'�+S	���=�c���2v��*��2�����]��f�R�3B#g�w�U_h�� ��:��fẺ�U�ou�E��;��]�D�!�����kqn�D�pv����Z4�X�F�$+�V���#�9��]]B�ڋ�����ȨVVfr��J���e\�/�c�Mq���kyQɹ8`��VC��X�*�]����s)�kOY�t8�U�'XC�]9�;T\�&b��N��;.^h���4�D�Ҡ�T#B��;�f�ެft1�(bo:_�(,k�{�� uS���>	՗r�Ƹ�Wr�]��g�z��恈\up&��O�.Q�б��df^�N<���:��.���tE��|�hS�,�R}p[�[/vAZ��ŕ�vd6�e/J>K�)��֧����C]� �������@"�!l�E٘"/*���6�,�r�	_f��?��Ԙ�����WO-��0ЭT@�t�2����!m,�z���9���Wrbↅ�Z�9gu�յw�-<�f:� �˭�6(A׭"�����ɵtF�v.��hf�u��5p� �ə��1m+(,��b7A�l�ٴ���WE���.�����k��VK��s�}8�4JdB�4ămϥ��㛪s��(��2ɏ��M��n�@졝ݙ�-r�=5i���\h�%Ȁt( W�
�T^�ð��p���lr;�jI�_7ȮTgZ�;��ٖ{)f`7AF��c��RAf"v��]4@�@�&�����8�yNא�dT�t2��N����Wp���M��WϞ�]�g;��Y���G��{Sh�H��|� #1'��[�5�no��Jú\�G���b�GO7Z%`��r�6�|�	Ƨb�-�L�q�qu������Ӵ�4�Ձ$�8�":e��kRh^�bH�P&�s�e�'MEp��[�Yږ0�v��Lwǯ�U�7v�l<1�R't�@�[(9�)���ҕ5u���77N�j�3���N�	n�kc37����b�Afu3n�U�n�P`������}�2:����E!���;��������o�_��Q-|��l���,y��\�ºv�rX��2�k�Y�a;�ԯ�Z�n���r�Z�h���K�Sw�SO��
�������׌�-��&Ŕ���W{d@�v�� z��q�h�6��s:L�8A����بQ4[C���Ht��(��hD.�orP�ӻ��=���Pa˛.t�����fBT���'�����R�tR�Q���mjIF�o պ����LXsb{�w��(����l�Y�xz���8o�[�����J]��MUiD�Q��2Z6��q��:��1�gL�v6Gvdj�jJ=��ѡS)0�����(>�Z_\U� d�j�r��������U|���:7��x�խH,�6��ӷ�8�ۢ�e���'@N�2ҋV��`k��{}ve�0*j�AfV�ci�9Y��v���W�i�s�XµiN5�2|�;�d�}��'�4to17ۦ�c���iL���[��0�ZKv�����t/��O�w8����n���C�n$5[��&<7O���O�w0h)!�)���*u��!�H���Z���+MD�r�Cz�qOr鵭��PK}�yM �ۛ9�[�����+�z��o~��t[�K�}�sW#��M"�N��w��Ϝ�i�#6�Ok+;J��1�g(s�p����/�W/�W2��r5ԅr����|BC�Pkx���W�ʸ�5W�#
]��B%d��M�8�.�� +aT!�TG�^��E���k�ft|�*�:HeŚ ��BZ�����2�r�0-)�W`��:��X0n�pu����㜳�:���G�^M,�ǐՁ�M��;�Wu֤��s2��Fh��d1�6��ʋ� ��2�d�s��ʎ�k�,O�0ԊDҮ�n��%��9�D��7 I:^Fm<��'#���.�2 ��p�)R  �4ۻ�䨽�o�d�c2�f�y_w@�;�{�)��g|)�r�4��uv�RV���=��ݗ���M&�[�o/z��U$h2��Ivf`��j=��|��ͺ��������A���{u���a4���1٪��9=�N,�4mG�����.vpɩ������Ϻn��i�P��m��yc!lH2��`�dOE:�.];�$����@��k�K�Lz�c��q��x,wǎ���x���Z��G�J���2��h}��п��C�ǖFM]��ε�n��[�]ڢ<���#t��A��M*��zR���,����g5b��r�9u�#�Y�h�:�|����7�3�ufiۡ�<�%.a����b�a$lQ�CrU�������x�Tuw�j�r�E�v~�31u�H|��Z��}��s���p�ݸ,neJ��2���ۢ�3��p҂*���(7䴢�xv�ą,�ݭ�����rݪ�ߒVv�yq���;Ev�*OL�
��BT��ٝO���;�z��<k
�h51ˎ��:��{����2��m:�n�q[���,Y|ssk�������G��n/������Ι�����8u��2􎭾 P�:� (���.:]M��'!���/�e�K:��X�RV�xM��:ÝZ��~���U𦲠�f�s9%Q�%fWXC��ʊ��'kWi����T��p��
̱/@8�k��u�u�U�L`Xo�	�m�Yr^NآB��&.��ղE�����ay�cv��u�v�����j�?1���K��\nd���m�����%��N"�?�����h�Nj�V'�����W�_}񯥪tބ��{���*�6י�Y�H{}���K��r��w'�w)�W��`;t��ҳ;Q
q�a���]
��V��k)m7�I`�N+��)�j�f^���u����y�銻��f�)��ʊ��X`�Έ�L�R-piu�<(J<^�������3�m��Ix+�)/�oz�R\ʼU,-�3R��ª�b��j봺Y���MeƉ�Z}ggB�̮���U����"]��Gz�_w)�\D!�|�ڰZ���M*u�P����9S����[�`oy�A�=O�e�ي��A?P�%vN��/�/R�1q�N�]�]Q��Ӫ�_���Щ��F����(�Z��6��o3xJ"��j�gU��6	Zv�����17����	"$^T��.�m���V�bQ�0`F�S��o��7��w�m��VAy��kW6���q��]��Er5μ+tȍ�(d�����2�q��̪���-��x�N+b҅�{[Ngv�ј`�ldiTs�n�mj��'��D|����Z[�_�ͯ��J��q�Y)̊	N.Hf��c�׎��voD���MeGś�����j-�|pe7N��rXZ9��	���^�ڱ{(�������>���Ϻf�k�����mήE1�9�'��")/累C�rnf������ �o_Mh�;���u�^+�R"o��Ž�r������W������e��نfeT�Fe9�Y��~�uDUYdQf9fdD��QS��VSVF5���ј�f8�DD��QPUY9Y��Yaf�Y�$UY�X`ŌY�EfSLADfeTU�%�RUU��%�U9��T�$DEI�&��L�(,��02 ��*�����5��$�"��JJ��*0���,�"���*��(�JL�#�
0�,�
�,303(��q�,���j" �
��"�Z��*���ud�D��ULQ%4DT5EI�ri�3�(���"����30��(�K���H���,���p����i�*"5d�D�EDMAM9Lf��Y5EAUQfa:��!�(�5.U�PET1%5I1d�CPTf�QS1U%��U3SESMD�E�YQSQAT�QE��E��`EDD�aYeQHQA�I�¤���A%DEe�Y�@��+�fk�:0N�_l}���F�L��u8q��"�bh���k��f����S��x�RYCn�ذ��M)�H6�=_t� ��X�w�2����ӊ�\�q�&3�����+ �(f���a�7�b��������yT���7�_ع�bNsS�nW���F���R��{sަ��~�w"7h����`J>�W~0n0������|"���J6�+urI��[���:�8%�-ܱ8�u�D=�ng���<t�s��p�ޕy1Ōi�Q�M�K�ox�]��)�91+\3C�[66��^��x�a�t�+������1B�njY�3B�7�q���{�y�:ʫ;��� �ڠqIS�ծi�FǝD��8�=g�&���Yݗ��+�ٍ����������n s3�fe�߽TN�}���ͪ$�����g��W��~╹�iி|�
�͕�o�x.�&R�)Q���d�7�6󲇮��	�-K'nAϑuI��|4L��ʁ9/ c|�>�b��dc��)_խ������a��j�Xf�ɽ�m�Vic����8��]g=���s1 pq=���6A�c\�)���,�R��j���f=�{.��|h�b��1�K��B�/��P�/����ey1t~�o����n�]��?itS�����G��YT����s�����^����}���ѤJ2a��ަF���/���u7bD�K����;�f�S�6�تyw��>9`e?.667�b$,ꄪ�U�]��Yt����V���t;���Ug��򪆖Wp5g������i[�D��t��z/���jc:�H��չ���g
��m���YY'}V�j�Q���dc�iy���W5�g�A��,����]U*��"憺���}QsP�1W�y�����/\\�����u:���-�_�$���c�ue_�����[��5�B��\>w�~zah��W��'(��0i
�x��qu�o;��*��]�a�����{�C�P�6���/7�ʗ����tP���14U�ޮ�]J����O���^������F�r5�)7F�Q��;�$�Ll����4{eI��̷Wo�k�(5F8[�7�]<��׌���,zPe�)q�Phu�r��wr���;2�k}
(�{C�wo�#�`�1+���(�Ӫ�\p�\2(	��*CF�5n�߰]D������;�+�q�(&N�a�\�a�J_�$���i0�`�b��2���]�j�/��,,�
x(�����C��=-9�z��I�q�xs�')We�j����^U�ݒD1�u{����кv�l;��X�Ts�u��0�s�8TX3��0���k�*��:�]�bYM	�k1:Yu/:N:{���JL�-�L�ŝE����&�m{�;�nS=NAa��~�%/
�G�ι����<��J��Dɠy2E|Y�G���X�\�㘴�3�P��_�h)�Wv�)��`��0�JZfܱ<*S�C�x5���b�9�}���ej�H��ZE)x���¸�Ǩ��"���ĶʄP�i�rSȂ�y���=xcyٝX�i�Q���� !��JF�e���*߉����X�s=Q2NB�'MS��ɷf�#F}#^�sk�U�WU�;�$�;`i�/
t���v�$R�ӗͤ.�fnM'#6�	���J��Lmh�6Ah܇���\*��%،��`����Z=-��<TQ��8�%�C�Qs�i��I����M~5Jeҥ�"�0߫Șz����hvKޒtVL�ߙS�u�+D_���_�(��vs��F4�D���O���a��K��e�fik����O����/ �V\N�ĭg"%���|�2o�Wvt�1h��]/���9��W{�e��[�N}֮�6&Z�3�13�#X����_i�=9����wHu؝2)��fׯwL�	���[�5Z��������n�6)�2�1�h�J�s��'"=7}O=8��F)^�����B�"�6��ۂ����k�CԹ���[E�����*J���d^lZ��H�`�����e��6�;���8U*���|��}�F1J��f������H�񦫎j�j��0�td�J�.g�сZ._v�v��5#gyR�6])�i����)��)��Uy��w��g��+�M$�W���zC0�jR�~��7ԥ�0���s���.@�sA�9z`�>�*ͥ؉M�u����C�˾�SR�n��ѥ�vw��Q6��{w�5��pf[T�t8.�2(��C%��x�,�2�.>z/�&�����Eu�͎N�1������[v�7�C_e�=�Y��S�UD����P�D�ʄ Y�h�Ϻ����q�R�'v����F�MV�M%:�����'�Xk�riI��
�[4���އ.���+�Cج:�������)מ�*W��[S.p���ʗ�ŏ%>Z�=�ı�/�)ķإ8�xT��v��ˍǷX�n7ͩ����8��KX��Cr'���"���L-l��H3��Tb�<��û�&c�5��w�p��MUgZ�W����t��2� (nrd>�5�O*�E/td{l��rrv��bGe����1��o�U�㘕udMcoz�Q9�M�"s���5���or����r����`l���;�oP�F��I�n��؅�u��<�kV�4�����V^r��9�Áu�>��ocl󯯳�C�sģ��R~j���ɶ���cԯ]�ܵ�V7��Vb��DT!LLD�>vp��D���|�{0.U��3���X~["|tj8���r3���'��.{Ѭ�3qF�z�»+=��`՗������e�OTpZu���D��#&�k˽A�q�����U�_�U��L41ւ]��4ma��6�%�ݸ��s�MD>='KH�]��Q`���p5��Z'%V�%�v����.��2\�`s���6&t�;��j����yz_:�>"��?c�т�֯e�:��������Uc�����Q铪by�z�EC���.u脌w\0ޮ�O�����ٍ�BR?z`O�/�����q��n�R����f���@U)�����8U�x�d��2წt禈zH�=�N�]����V|p��XƑ�$�,�6��˻U�6Qe�)��[�Z���V<#,hk��>��|.}k8�sf���{��-�ބ�wK��0�67��D������X7�\��A_�Ϳ��j���wϠ�Z�n9�W��Oy;�(��ASܿ7C��U���g^�9
��W(��z9�݇�B�\m�3�P�#7N�Kx*�qw|��Ε�E<r�[��,Pr�kWa؍n�r@��v�v��x.�L	����-�r;�)_fr�&ls�͒��1s����g��᝖�_d=U�-_�Ϲ˸|�$s�FI��z��f�l9U�+@h�N��O�������ѵ���j����K��6�C��~��.�&RE��&N�n=/�Mg۔|=�nsoF����ë9��h�f3*������v&%����?J�[F�o��g��zv��4��<������"����ֵE�R�5@hnra8��Έ����ha8�W��
�h"�d^]����05k������N�	�o� (�^ ��vá�{������g�b���UP�ʛ�?&��'�=��y�� �g�nE&[���j�ã>Z��I�윆�I5�H(�D��Y��`�K�����!ۧ��);O2*�q����:�y�S���.i�V�9��x��1�*h��1Ȓ�sr��ث�uH��E��3T3^�|
�!r�:��zah��+��1�-Ԟi�*����N�svÌnv- Vz� �����vyRj��9�=�Z��=��΍��|`�BB﴾�b�6ҾʖЋ[啋"�7�XƆ��3{��u�JΥ:�,�3p2\�ށwBK���T�
���ݭu-�/V4��af�*�wVOw	Kk�:r��D��^p�֝�����*�{jS���]��d���������\ ��F=���|���m�*�L��C9Ȟ���I�iTvyV����ip!w%j��X8�e���m�@
��M��q��kTr[ˣ*j#���R��ݼN�����;*�j�O�����'�c���e)�
Ļ�q�Jc�c+:�ӵب�]0\���]ׂ�v��ّ��=Xf+����-/����)FI#���a���*���S�0h�m�{�d�EWK���Vb��ϖ�"Θ��凵�L�J��Dɿy2E�b�V�y�Ã�Ԋ�D	�%�9�d���тgS,cO!��R�͹bxT�臾S��e:�Fn�Sݕ���E�@IN`c��A�c�c�8�}h�X��[�`Cc�Y�F׆:���L)��dG��=}J멥'�t�sm�D��\䬼���H�j,���m�n*
����#�{�z��J�ɕ6����d����\��c'ǹ8����d�O��R����c�Wld�	��|l��VHh�'g��1{��2|�Kբ�+MH��7rQ��qZ[f�r�Iݻ���O^mN.��;�t餍5�P�����xE`8��QX7�m�a���*m�#�g��v14�u���Ʀu�.��n���e��Pv�gc�	�#��'u��4R��i��z�3|����C�-q���Nw�ʉd"��\̟>u��$o��6x����I�u>��߽��59��8�鍌;P��
��ű�B�y6���f��ʓ�-�3��z��n:�#[Ƴ����z��%ו	�g���b�Z�K�����d���F^b���ݐ�7���0E�H`v��}z��:��:��|�"}�dL��\���mwh�{�=�#/1�Y�ڄ.{�U�:�e��MC�5\sWZ_-&\�bu2��O7DfF��Vm��ёwda�̹]h��!���7-3���;\_>�VJ�N��.�q�t'YRҺiְs\�!�7A�󫛌e�o+��ɯ���9p�+
���%���U�W������z�{��a�X����Y�+���W�}�P�=�S�.�f�<��x�^��6*��޷ڹ�p!�{�vD¾�08䨠��u� rw�G��zT��[w�0�#,�./70�OE���$�|.��2�z�W�%�c�X���]}͸|XY�"���o�<��3�{2��������˵@4��(���y	&g�N�PP9��d���-�^��E։Fh�PX�����ҭ���t;a�jV0�����-��!��ޏ�Sۀ��_��U�j���)S˩{�Bl��T�����3b����7#�]���@��������EbJ���&#s�8b�����-����b7.�e9j����wV�vu�]a�:�F#b��UW���Mʌj��ׅU��0�s�<�h�X�0��Uu	�:�<���	5��⢼�����l��3�j�E^�iZ]��J*�w$�z�Ta�U��9�f�$dF����B���GD�3"`�WB_>xP�Ѻ���m+)��w��`�k�;������Y�p�0k�1a��C�#r�X�ޤ��J&�����2M�?D��=H����4oL6:�x�F�qG�v�2u�N�n�o�M��."^���U���D��B2`yw�˰3}��p>u��׽lz�sk\�K��ղKfj��Y6�wdt��'��������Z.V��s2�Z�q{����k*�ўl�\�"j\�Bn�o�S��tsAg�8.x���T��A����x�ٻ�{l��4)
�uQ�������;��'T��S����u��k��{���-�(�pxi/��luFg	��ڞ�-��sb�pS����� ���|o�C9�������b��s볰]jgm��<�Rb�\�g,�x�P��]N���ǻ��lt�͝��a��v�NdR��}��h��������M�����lW��D7��x�;���)#���}J^0c���ΊE�"1=�t���� �����4�����1��rDm�ᡇ=�+/瓽��V�y񋓓��׽���l��#x].S�D���Jؑ���j�`��X��v� �>��%�w$���\�mrda��5�n����zu�1,U� �yP:�T�ƭsUfn�;?M�͜�{��.�:y�4�R�:�n�s�|:�m������/G1#$�W������~K}�=yu� �b�������Pn�����P�&Z^��D6�B�U�ǭ��gȡ�t�`kL[�F%�N��ܢl��ͻ�U8��X �]�#����`%��݉�jR�IuY���|-�����>�n�o��G}D��b�,E���wY�<G�X�֨��
U�[��[�c@E��NLsO�=̝�6LB����.��Gm�Jb�Յ�V�Ϯ[ᒱ;\ocxoe�*�7C^^�͛ �^�W��>���ӗ�U��*��x�S�|���aAB���i[���o���W!�P�}�*�O�vJ�u���e�h�i��0	�)L��{��b���J�,嵬s�v�F�:��T�n����ɠhP4*��\E�r�g���c�z/�{����v�l�0\���n�X\�.��3\ڎ"��z\d�Q��bcr�a��s�+.n�*!���[3\�F��>�x�Sq�c{z�!����e��&��H\��YX�rU�uc��v /$��;��Nee�n�o��.��F۞K�e��Y)�5sP��X��#�3/����͝v�oE7Ԕ�AX2m���K����{��bZ��F+-p�_:��a�01��v`�}����$��q����_��cDȵX3,�[X�9�+;�A8C{��3�WK�K�ΐL��_t�qoF��)�*\t̼tt���xve��������kk�	��pn�d-v��Fc���)�9��n%�o��+�J�楘�{�YGi�7�V�*<݌��X�VN-p�6�6ի��"RPXk���C/���w0�|Ǖe��ZK1�6P5�[���/F���&j�|�:6/M�g1z�������b��Yh��[c#-��Z��h��b���L��X��xj�N�2�;�m��U�4H�Y��mеj�<���-r��.� o���5�Sξ8��1x�5);��/��.T��nv�I*N�.�*iܠr�7z1��Y�9��%X�e�E��[ݔ4�ޯ��'�a���S�E���x��چ� ��jQ9��)M�� %1����>8\ύ`0�j�v��Q�uʕ�9&������B��]��F�!����j���C���/Q�FT���f�v�sg�yJ0Q��-�E^�68,х�b�Ij�8Ծ�˾��^lY6�ŋ��q��t[8,�tQ���H�ܝ��M˩v�˹)�Of�\���ܜ2�2v�fEZ��JwR)\}��CS�X 鷉kOpe_	+�����9Dh��kf[�t���7���tg�S$>�뇩Ly�V���h#4���=Y$]��η��v��X���7�y<V6!	�S��;�o<�b���'�����^�<�*��a�o{ [o�1cH�7|ci�nd窖c�)��!�<�䅱|�xH��-�;�������.��Ҿ�����C�hYk��ʺ������8��Y6���r��gk^ᧆcRk��&��vS�����`1�V	�ʨ1ޓ�5��Pm�i����������<k��ζR���9<,�:M1��c�U���m����P���zÃ$���ǻH�neAP�s��r{j�^�|н�2!0�cu�8�GC' ��"]8{��s����o���Aʍ�ӳr�EzALL��N��c���{2����ڭcq�6ժ�w�U�x֍�J�1��5۹�+E-�>���#[���řĘ�M�;
�=�, ��L�v�qS:o9��f���
I�ª*�,��� �k�VEZ�(����(������(�� 3J���3h�l�b�s0����f`���d�*���&�&�j��u�AQLQA5S1IE�TAPUIUEU�3�L�3�rʒ�������
��(������%�(�B!� ����"��*�������Y�4TDD5MEf��M�DQ��̠� �*�����lq�(��������
*��kFU14�EUD5CQ��Ta�UTDD�TQESSQ�PIUTQUA�M��&	�
���*I�a�*�"X�f%)M5DTSEQQM5CE1E-QM%1Z� �(�����)*���TRF�*�b��a�ZD��a��9�9LLVH�S�EZ�)���p��*(�(b&)b	��(2\��3(���(��
�i�d�����+$2��Rj���Z���|���<��^w��6b;.��/��ԓ�S�p��d�F��G*��>{¶Vqb�ŗ��m�S{�Y�.�G��=-y�T���#3�j��V�f�{{'<�i&���(�H���cg|C�1Y�������O�-��Ҡ����K�n+�E�}T�cꋗ�s�7[���J��.$<�Hx8��ޖ��\�����p4b
�G���^�yY�o��lC�F�y^V���j�I���w4�+�g�S�r�>������p
oJ�����qI�Tn^�r��7��n���:q��(���*c����b�K:�����/_Z�D���>5hN근!B���w�^�z�7�k1�����-���]D����������y��W�n�k�[w�Ґ\�ܞ��N
8e����Jb��9�ptxaLJ�f�D֝W���ޠp&QkA�Zp��;,�6�X���p�pH;�%s�n-/��5�OJ$��.���Lo���멶�.�D��/�Bg9��E���"Θ�w�,=��Zf"TN੖�X�ۘ�\u���7���WU�S0�}i�cj�������W<��JZ�z�ڔ��j0zr�����E~:8�}�v"�7�c61�`ʑ��h7p>Jۭߧ-㕏o3Y-��X�4�/g@�c]u �s�׶L���ƌ�91��[m'V�
\.���y΋����X&��Y{�_Q���44*N\96&�f�ת�ok9����{��Hݰ���E"±���h;�3����<Ɓ��az!a��k��JG�)*�hJ�A�
���Ȋ�cbѮ��6�&�����0�<yff7ӡ���p�iT	r���璪�ʝ���5xج�(�\����3<WRl#Yܒ9�MS�����y�bkM�j����N�\�U�tA��MH�&�bO��#��qk������G��(
47�}P�_M���VI"��:
|��r�d�CV^�wɲ��+1o�u��ʄP�c����ű�8��wA�=Ef��Ə1�:d�}�B���>|�M6���z\Ɍ1�����1~����7/���;��7]{o{�6�U�i�I������&��Dޠ��|����c���;��`���; �����ΫZ�'�vf�}]�=�,du�t�Z����b�ՅK�o7`T2(����C�D�~L��P���5<�z*a�z�^yN@�)NL\�F6ݚ�!@ͭ�Ǿ�z�l�h�5�}����o��Pշ8��y˺�!qR���[�pb���[��XC�)�csΊ��i�cD��󹩃��4��zD����h"̼�h�7���pp��]�j�y^B�pۯ��I=Q��a��Y�_ovo#�h-��*B��a�Ta�B���z.{�`^+�<R]7Īj+r�R��m굕FB��l�Z`�\�MOqJ��Kl���s4��on�f�<=�q���{���*��U$,��FH��4�w�ܺ�+�6lrw��=/B���,^�~oc8�Krvw�cx�c��)r�zQK����P��yX�(+=�A�sn��E�7~��M>��rޗu�Fu*��,�HE�+�[f�����͜5�b��X�O�l�����E&y,�~��R5"\כ��2��'O���MʹƮ*�O=9�N���;rcs8��]U3�A��v�*����g���y�#�|��2�A���x�I��/��F�F�F}�w�5*�Yخ��ى#u��yB�@�qd-d��f2D���s�����^�S�)[���%Q�tV���-ϽP�ݙcL^�P�0k�1\taU�&��=�G��B�������]qv2!�0g���T�'eʄLd׵��sfH��U�{/������h>�t�x�\���X�;ƈ��G˦��s�Q��f2y�o0�Q*V�9�^�]�Ȟ;��}�u��7iJ Yl��9C�x����h��qq�\:#�m�����9�VsJ��VF�wWL8��E���ɸ��j�ZI��BL�B���x��Kُ��ꚡ5��N�;gsb�ҪĂ׍;�|1�z��;|�I�V��O%����^L���,l��Ƌ2T]t�ϨJc��K�7�LÞ�������@W,>�z]��H�������6��y|��Sɡ^�U^�\�A�ay�ם�]-��Vw�x[�8��'���nz��>INc���U��\"�w)B�پt���K�l�A}J^G�1�ܕ������o!����0>g��9��y���!�Q>H�=�OMME��74�dM�c�Y5ܛ�Z����L��lm�L^��/�=�%1�bGV��IY��gK�Wk���j�SxV�no��x��=����d/Ua�R�{���������/�j;��J��{ۡ��~�����LS2�>5�{l�9w	6I�2Lg �툛]qUt�d<3�����T��5YqBg9���}c$���I��q�To�yw�2��T~���~��n�5Y���^��:�%wRC�u�S���V~*���QH4K�����p���+c����n�f`甚5[�,�e����m���Mab�x\���\)јyAA~;5ym���׽�p�ۢh@�Ք��=~w����'ZSt*9; 7�wު�Mw��u������W��N�3,#C�X�%���LK�`@�u��vZ��Oɥ@Ԣm6q��ڙ�Y��g,�Xf- α��r�;ê�:����st�M�|�RL��	�]Ku�f�*g���^����匧�����̹��"�(u�$糶��Y��%a*�{��yspo�V�j"T܆�NN·.|�{P�{��]��jy����/̗��3��>
�L�4��KG	<��nA��`�a�xT�}�z�M�X�]T����W��ު�V5�9����	�Y`Oun���y�@���[�nv�v�N��H�DE�����I����o�5�5.w���M�0�l�ʿwՑz��'A�L�����F_��������2o���Z��qITn^�un�b>�w�9�<ͪ��>c�0��rI���CU��E�/�tEZ�g�:��9t�&�s���6��73���Kp�e1�IA�X�o��~���ڱ�\hp�҆+�0>�t3"��g1��WCCqy���>v��.���W3i�v�*ɗ�u�V����\����M1�mq9ϡܼ��Z�wt��:}n��贴���P�(��K�[^�K]��H����7s�����F+5)�5�/z��Y����n�o.��@Y�&*[e0pk!�yr�=0l�u��A�%1����|:����yJ{�wn��sf���;���R;7�N^�=X{�N�lE��W��(�F�0�<�py�&��8�wwq�Q�k"_��E	�|n0\�-^��q�Y��Z}���˸��J�O�)�8�v��#�9uA]"d���_*ȝ���aB���ӫ�YN��8�^ք}��͹;zw��S�z��O�X�FK�d���)x���¾R�D�edFw�΁�'/M�]Ar�k�T]�ƙ��[7��4n�\�1rd��4g�{c��x �J��SH��H�;��������-u@�5�e��U��(�S�a��
��lVT"�U���6��YTt($�m��6#9�F{Q�f�S��as��|`X���9VHh�'g�N��&S���o�4�5�W�mV6�lu���O�u(k�$��V&�I �B���ŋSQ�T���9�\��tql��;�v�\p+D_���)����u#,Y�Z�]fg�4+$�Ie��&>F��0��m,�u��'˹ՄD�\����J0�og;��������K�@��i�V�8��p�+�ݦ�I��v�u�1�٥[�\�Wbj{���T����zCV�Gw�	��c%�����w����L����	u۬�w�+�Qgf�u3�+��N�|��%k3wz�(��Y;��Oc�}���>�K�V�iUxn�[�ۼ'ڌ�WNd�LL�mB� V��޵���ȎA�%��U��؅/ۍtsI�������r���J[�,n���+��߳ڗQ�Y�F���P��P�r�w�����3�c]�<�I�O�����M�$H��%�ݞm�%W�5�X,bf�}����B��R�As�u����`[�����{��/T�@S.!�sD�6��f����+��-����.b�mA���a2�����{~��I ���� 7�C�UC���|��՘�X�w�>[2�wn*��ͬ�k?'�$e2�(�V��9tP�_�d��d�"j'�ec�X���!Gݍ��ge`?k@諗��Up��W�W�m;�&C��PB	�`7�*%
�ѳX�+a}6����X+e������&�=�.���1�2�.F�6[0���H��7*�q�����ԣ,J�zexwv<�<��nY`�3�&�,���gW�ܭ�; ��`�j"�Z����R��qǋw]�p�N�a*���0!h�)EgE�u#T���t\���e��7y���W�
�����:W&	dQ��k�sdM�$0�ދL�q����g�9'�M��G곓��!���I�GD�5Ě�r'(�Fu}���l�N�`e:�Ip�Rr�8���r	���L�b�&eU/}����794_du�����W۾̵Z%�DA%�i݌��VKV~�ڼ!��A@�_dԟ'a�Aw�HE�z�E)�e�	=u�F���T�+?-b'���1y�x��|c���}T<MV��]�cC�=�JP�d��H�-b�ɸ��j�U��n��PQ�F��M��|���̭N���q���F�����;N�_�βn����x�|zA�l��5�V�]�w��:v��W�)9�j�Jn�D��'#��-���"j\�Bn�^�[:��\�W�Y�^ R�]��K��zl���+X3SO�{y���W(d]�v���=6�槮�=�}��^E�fa��S�a�
D�a�N�.v��L)�fR>�숾wq�$`�m�����An���_Zv�iŃ���36�@
����<�Nzh���%qTfoî^��}�iȺn�]�*Rc��I�m!u[+�M��!�ʔ��{�T�Ҧ��4to�L��壁���ɗ7�W����յ	��h�O�z[�=j�g��⓵+]F]�tt�}�+:[:�Q_X�}�T� {N�n����7l�![yI�hgQ���o9&v�?���BY��N+n��OSҹN�t���(pĈ=�P�g$fֹ��:�m�t��j�$�vmچ��e*��^�9�X�Z�l�:� @Ţ�{��SS�:�ӫ�w&<����z���4k`o�k���s�k+�L�B�����<�$uz��l�=����b�8Iκi���J�C��n�nuo��1%-/:,:�Cb�~��.�&R��zznU*�u-�T�j�5><���V��$���V}ҽ����#�Z^Z�kv&%Q�~K����i=��f�W ˬ�@�D�� Q���
���Y��2=3Vң�e���HC���X��(9`tKo@���Y�-td{l���z��ծ���m�
gp�q[CwF=w�ҁT���wQ!j�V��N͋�*��T�*u��`�R��d��ж���Lޣ�eB��])@v�fu�'�![��i���5ZI�1���9;��,�N�5�k[�5R!�pC�2ϔH��w��C�kf�{�Yb{^b�+ب��J���{��)�T�6�}(�C���u���eI.^���uъ2m*�-�m0��ᩞܰ�A�32���ة>��3R�C5f�p�8�����ǆ��ic��Ov�wc���~�%�3t�L��s{F؇Ov���ݶ;�����{ʱn����w�m9�#ݢ�'�`Q&%h�u֡q���b~�}<U���c�Y�p-,�).n�Q�]�z[�v���F_�|\���>��ծM�AѮ�*Z{�`��"Y�).z�	̿c���>�L,Os�a���$�,c�蛋O���y�����ky�MdK:7v&��� v�p!��Gg��8���x	uLr�8�kz��K�~w��qV�Τ'c���lM�~˻Y5;���e n0�َ�ų�js�\a�1*��(���W �A:VoVpC=�t�l@̬��ЪwŪ�x����=��d�f���_�bRǣ���3�ڇú:uԵju��l]����� ��=��0J:�*g��Ou�O9+�O��n^���#p�������$Qfb,�"���jǑ9��+fP������>��F���o@Svk{��*�B.�j+ Ƒ����ڇ"�>tgJ�v,�B�ju�3���ۦm+���p8D�1,	)�AxWz�+���Rz�gKW6�DK^�����}P[���N*��Kԏ�8W�7�^L���hg�/�*��E�(���I*4ʴ���v5j����f��a��>�M�p��pڔ�4n�$sE��Y�o�_��Z;��C:��Έ�S6ޓ��oTv�x�vt-�^�w$�e�:���/L��Wn6ux��ֳj�cIC��X�<:\��P�NC�2�3`��=rj�2�7-�G�bo�+��sf�v0�X�'1�G�]���Zh�zi*V|^�h��U�����ƶj]v��rNd�G��)8iz����4����筄��oV*`e��A�O9��k�aߧW\����W.��Ȼ�o7��ܑ��(䱋�b4&�<w�fpB����ˡG����;[Հo�[�j��fw1�C�Z1h����萮)S��j<vy2�
��Ŝ!��G��C@�%e�R��^Z5I��6!�����+t��{Gz�|.�Q�Cr\��ٖ؃`��W0`2JL�r��a�N�ǷN�v=�0(�(epx����ī��'Wtήm<���8�]��$��z�a�z»�,�-����P�(�3�mL�0V��m#0եg�^]�"D�<��lU
�:�d*W�
'�*��%Z����9���
fmݣ��"�����+��q�X���YˡL�g{�Hʘ/�SՓ9̣�;[u���\�i�pq.)Z3�υll��
Ȥ2N߯*��9��l�ݹ�?��+��甞�9���FX��9:Q�ĩ]n�����e�,R��ԯ�e��kfu�A��/[ܬ��wQ|y\��ZI�@�,
)l�{�u����d�,Ӡv�f�Wd��:C�:Q�Z¸�ڻ��9kEb��&gsrܬ���%ۇl�G�)�̗Z����m�V�_��5&Z5e˩�7�C�����%�d��˝r��ϼ����Ar������si�Ivv⫂(u!gkW7^���G�������ܵкK���u�[�(8M;����7�dC{�Q�kQ�yU��N^T��,9��m�*W"���R]BU�4����r;�[�BU�+S]��F^���Hʅ@�ط���R��qm�{��z�f�WL[mB��e-�k���H)�L��q�4�7t+��ξ�V�w�"yuou#�^ki�{nʰr;,�}zv�r�Y�o�A���urߗ7���qK *�D^��)JW[q�",A��d���(rkjf���i��^�}�RC��:j�2�AKt�9���c���Nٶý���
��U��{IÊ��b�1f�_�P_�:n���2�c�}�vr�ZB�Q�u�������nM�)�+҄���,Yv"�#���k��&9۴mY@ť��<6����]lq(֋�q�^߸LѨ%��H�+7]]Y�ͳ���O�E�w#W��+*�+�~��D�SCQ~�*i������"�����c"!��)h��Z
""bi� �Փ3N�%mf�R�H-%%��D�E�Mf8E5Q4�QMLPRY�f`SMRQLIIED�5TA�E4F���d�Z̦)��-baP�UQD�fEe��3AKLT��RPSMQI9��$E�ILBPY$�Ed�M�j���
5�1�T�LMa�$QS5D�AUYcPTLL�SPQF�*����
���+X�UEEQIIQQALCKA����S5FfQDB�DEk((��*�����J� ����Jh�����$�d����i����i#VQD�E�T5Ee��UTTA��UEE3SDT�A����DR�T1k,��BX�
Z���Ƣ"*(�s2 �"J"*"�)�����3TQ6�$��)���jbj �*�
���&hb��J���*�"��i"j�g�<�ߵ��|����Ú���v��	�w[׹
LC����2��и�ʻ	n�(͉n�i�\Z��oI�oa��ﾪ������ۖ(U� )�	À?�s&T	s^z׬��T�2����5x�7�^�y�o2t�{�Z��)Ж�hOf�I�����8I]�������J����]5d#��w"�����3l}�S�@8hx�<���֑�Lb��'Ρ�:�'����V�H����1�d	����K�����V� ��]bǵƠ�b.K�� P&��GcÖ���z�Ń���;���#>�rЮ�E���X�;��+@�1�*�K�ͻyM1�K�]5d��EĹ�|��\�����S��7X�CU�=����U�gn8J<�61Q6�{�:O4&\1�B% ��fo�"\�M���mP�ˈ�#+X�³X�K����7/�D�ٳS�U*q33�˘��V�\���0�9A/�o���*1���=�{o���d�1J��P��z�B����2�7|Я7ԥ�KU�g��HJ��@���Gg�oe��P�I���Ux\�T�JuW���:���T���6�{��A�0���B"��<5���2Lc���
��5��q����u��.LZ��Z���E!&�!`���NW����TT$ς��E��I֥��p}���ڎ^tO�T��/��决�'�4��ȚjϽ�V+u��zu��Ū4ʼ�[_{��G�v�v��6N�`�3<��vL�����b�N��CN��w�"�=���gi;{�#O��z�J�)Ǘz����V=(�%��<����mg�
>���*Ep$��@W65B�,ʖ�����t��F�Jq�5��JOb`�+�l٬S?=y�Er]_d�'A�nc'L/��R�VY�1�2�.F�6Բl�	�Mʠ1�OVbÔ��6�'7)��1J�.�yT���w��q&�܉�EEy'?�ʾ��<���ne��T��HA2O\�W�O=0Z���XD̪�዁��"��&��x}�w{���B����ʬK�2;l��O��h�s��^�=5R�O=E,CD��5y���vp�Z�a��>�՜_a$9��ކ+'a�ј6��q��czaU+��,���ROt���oG���枑(�Ǒ�r��Ah�%�&T���.�e�mĵ�s �;��E�E�3.8�n<���;�|3���M�����s�Oy���
���/4R��'�H�Icw�Zݭ���p�^<�כ�:�e��Ob�zF��R>���>��m5�aߏ���iW;.'���z_Yi讣��f-���u���q��w���u�]���&������+\E=����_}��_V�2���� x}B�_\mB�\��z8�0�U3t��L�zw���+��ݘ:u���g�.���vD�.����`����`�sث�2.��i����4+�G֛��_z�D��ɡgWI����:�u�
o[b�O�D7TAyΠ���H��p����9EW4�M�h���P����Z��G	�����Jb�������nӭ�}�3��Y&H�e�%�A*IV���F��y�V=�A�)�4���k\���ak��I���Gi>k_{�\Ē���pA"���՜��d�Y�X�L��r�=��`�bT�����,��7ُo۪;���F���;?F+_��ev)�Cg���r�GT��%{�רj��}�h=$��4�;��Kk}�ݞ��]�vT���'�;r!1Yr6���{�h�Kfō��T��2�d�u�
�����εYN+�+� o�u��NK�j���'����â�FhUa�Kj��q�eMLج�������Z�`u���-S�-�X;[�p�iX2�Ru���^����Y��iӌ��	�m�Ȟ��gYr���8k��ף��p�z�T�����T}+K���$�,��;f�t�İ̭w��rڵKc6%��Ѿ���0p��e�c�[p�a�j4�4L�-tZ�DيT���:�jM:W;�6#���ꪯ������s��lI\�@�.vtD�X⮄�� j}R�E�x�XYS��;6ܾ65�LYd��~n�f�30
.doO\ؽb�	�*���ʜMx�0 �d�C�ʪV�>
�� S�Q�i�ӜJ�|�ζD�bu2ӺRv�$�>= ����-%��}ʟMT���Qf2\���-�B�h���X|K�O�.^q�`�q��m����O�J5wj���j���qz�y���u1�������+�\�/Vaܱw���`�/�z�����v���!9Gg:�S����|/��x�oJ�<�\8)���;b�T�#�(�S;�[�r�p�s��}rI�Xǻ�7�Ko!���=�
��m�» �7um1f�	��S�bF��P�B�9q�8�y�Q7y\v;5�]��
���}���t7.v�]s�A��R���z(�ώ���.��C�<���;`�l�$��ob�FB��፧�(	���<]Nvo�N^�=X{��:ٸ��W0�'ˏx�������U��&t��;�M.ͽ�C������n����ftaP*�BW� �M��?}Gɹ̓��ht*_Z�e��,���Ln��74�E��f<K���������"���w����������[��S�F��l��S42y����1x�7������*�V�yT�33�32cB뉽V�d�R����:�*	�о����DJ�����|��VQެ��L�-@&ML���G�VE��0��W�Ns�c��=\�u������i����^\a��$���)�!ৃQ_�4�������׈�X.�ZΤ��쌀C��ޭ�\Q�-�@u�C�+�T6�� h޹J������:M�l�!<�z��b�N^x�{�x�cg��;;���� בs'˪�|E�N5ZɿAF�5�TT��M�r�*�ժ^_�{�ƛ4��k�T���U~{��g"e>p��v�%���6��gW��6�ٳ���v�Ӕ�d$_�*T(F/|N�1��a��Fx	x6\J#}
��H�p��l[2(����G���>���$_e���+���v�''ؼ)Z�]|
��ű��Y�]U�����M�F�����p���f�>�rЮ�VxoUEiv�Bhz��9%W�m��{�"�URF%��7/���ɷ��:u,:Dݡ��z�����{�tL���ǿa���@ z�E�jŨ"��Ä�n�a���OlY�n������J�dF��(`�a�v;��0&�V��&\�`��>���n;z3K�������c����_^�2}(�I"z�q��ݐ�͝�j��Թ�rvq�v�%���z=��Co�\��+L��☙�#xp	Ъ�_�)P�>��w[����h톝s���.��i���=�:���/�J�-P�oS���:��`ұ��P��h]��ѢsՖ��s��IY5>A��kȡX`�^����lh7��9j��x�ū�W^��<�פ�<�GZ����X�g��Zb��jj{JWz[gg7�����;��G��\8l��\s۾�� �8�¨�#�}��� K�.��+��f���1��NM�k��*b�+@�.�}����d�D�&�Xŏ¢�f߻&Z�<�d�ۡy%XuU�
G���=C��ԎY����`�14��j
$Mp鄂�[���05w��aBy>�$��ZS�9u���>���I�?A٘���~�}jW���u���������Ԇ~�� �y��U��\��շ˹%��s�����Rvk�7�v�ށ�y �����K��'o�������1�K����R�����׹�zdtw`��W+��dҠ��y�C����$�>��P�G�~Ӹ�)�k�9>��uޔ�w�y���y=����:���7-#Rt����=3�V����Gi�p�(E����2뮭�a���˳��m�ש�|��<��4����:��ǩ�6��:�6�tܫ�,L���|�h��O�Brӝ��M͛$��xq��I9� )Sn^�:9�ѓ,��R�C:��Q�5�|!�Ԝo���ꯪ�_��7d]\��g��>�ox���3����}5!����$��|ִ'P�Gy�P})�����/'���ܞ����L{�}�#���v}���Q�x��vs�o{��~��6}-/�Rp9�u�u��o�h���C��Oo?i}�Q��oA�&N����ie>��)�_`�_:�ܞK��v{��NA���w��w��5�wߜ>��y��^�����R�=�������;��˯M��������}H�<���ɨԇ\�G�9:��voZC�_s�z��:��^g�]���s�u���o{�^{޸�&���9�Sr�k�7}+��a�~��~�@r_y������~�9�:G�N{�I�{)�s���:����?�2u������g��nE��ɪ�U#�>���S�W�#g޹�L��ZG����4���H�=}�!�x/�P�q�|�Z�9'ׁ�s�|��翺wҟIp��w���1�^�6�X���������Ͻ�FI���u?�z�wރ��ۄ�O%��~��pN�9'O�~�+I��;��:�?b�q�{�Z�9<�w������s+'N���iԪ�\G�}��ﺢ��ި>����7&K����ҾI��3�N�J�o�R�����hwna2����b=@~<�rn7#�{�����F��~�J��?z#���
}��b'�s\�OҞ�
N���o�&C����H�Z;�ZO���s�R��S�˽�u	��볣��}�5��~�g�}�gR=�p��q�Oc�q���^{�����9��ӹ>�Oe��g�����7v��b�|4���/j�G�P7᝱9s.�����rֻ�8�ܝ�ps�C�M�Ѭݹ�;��prS����w>�ۿyӹ^����?�y�)=�.@p�ZZ]ۻ|�@���~���Z'�������	�\����V�� �5��W�x�R�R��<�gF�v�F�4�w���b�+��>ݒ����80�lp�۽��m31�{��Əwa#��ɒ)�/R�d;;�o$�O�N����bd;y���Ӕ�a�R�WeǛ���W�_}�Vjտ�o���Z��O7���by�e?����NG�vy�w	���X~��C�0�ϲ�g��'$�]�֟ҽI���K�����j=3�	�>��m��lm����������-V�y��O3���z�z��NG���C�7I����׸�S���y.O�w����5���O��O����ͫ�Y�k���I��5������4�k�hz��y�<��n��~��ON��{&��O:�Jy�x��J};��a��S��9'����t}y��w�u����y�g�Zs�tjW�{?o���r9ޗ�y�C?`�$�n>5�)�'��sO/�=Iޱ>�A�g]�gs����>������*f(�?�x,�H����'9�䛗-C���-/﹭H����.��k���Z����&I��6kZS�O�����{5����>����`���~�V�fQk��pu�#���j{��x�Ò�{���^F�܇%�����B���]w��}��/�j5!�7��C$�n<ִ�;��]F����+�(��߷sv�뺯_��5��;�'˷��?A�jz�ܞa�y{���_w��o �%�[�B�y�t�F�u<��䚍_�LJ#�'����Gvwn~�}B����<քܧ��?j��}��5��\�/C�r�i�Gһ��d����X�!���ܟG{��#b���C�?�����[�b�}�1��p�4���jC�����~7���+ֹ��^��C�;�/����nZy��r�Ò����jp�r<��}B�<����s�N�?G�cЧѱÛ��>Bvo��;��~��}�}��Ի�f�}����O�^��}'�{�	��'p��?Oa�)�h5����]��l�n�s�.Z�F�g�l.�KZ���u�c�)�Ê5}ӽ�aG�7��@�e�U��EHK�t����f0T��J�+��.=)�{ػ���b��X��7�g��}�Ι[��s@�LAY��f�ޥ��w�ڕ��\�t8������ܐݖ��6.�(�#�����Dz!�Z�� ]��}�ǣ�G1I��=�/r����қ��=�O �S�=yސܙ.GF���|�q����G���zN���'�X�CK�=��e	.ɾ�#��n=1S��;�CטrNF�u~�䛍���Z�?A����Jw�?t���;��y�9&K�����;��ϵ��7>�Li�΂ q�g�Z?*g莟z�f=:ǩ!��<;�5�:<�H�/~c�7nGW�N�俹���'ǚ���;����)=�'�=�o@nL�xK�S�[6l¯���睅��{�}�y�ݹ����]��s�@y�u�'�=��~��^�Ǔ�����n|��y�~��N���/s�}:��Zj��<����7���G�cU[�4���>uп��y���-�kA�����
�7A��!܇$�[��S�������<��rO%�_�M7��}7x�ow�"��_yϽ�G��އ��#���������ihiy�{�Z��gzM���vsZ��{�YBy&��<����G |��F�s7�WC�����g�>B�}�� ᘧ�y/G����G���u����7�!��p�N�2ss�?G�w���G�;:�I웽��<��}1��̙"~ǜ��芫��阏\��?a�y:��x��r~�Srr_M��J�^Ü���^ޗ�y�C�~�����s0N�?G�y���G�ё��p��?��|��rS��ގ�)�P<�)�ϰx�� �O^��N�:�rr\�_��K�����/%��huyG7���!�~�w	�L)�N,�B]��?-���>�5'�z.|�9���Oe��'��e;z�H�O$��:�%w�ǐ�:��7-/-C���4�����Z��Η^`�B�����l�2���Ρ���1�:5̙c=B�p:]����}��:�t���4��kB֗/�]w-�1��Ѿ�a*�RzEk�ߚ��9�Xw�̴��1ӊC:������I�B7��.�\U�oa��j�"4k�$�F�,vq{z"=�qĹ������>�0d?���y	�{G���=��{�ڧ����Ogpy'���G�{'G�u=���!�y��<��v���>��G�)ӂ
���=w�_ڙE\���@q�=�=�du>�i}�V�:7���L�A�;y�!��ٜ�>����X���r}�=�w'$�5}+�?O���rb=���I�׼wy�c��������.d����0@n[�z�OC���}H�|y�/������)�j{���I��z��e�~����y._���p�s�u���9�����o���5�Q�/�8�P��#�3P��b���NI�<y��#�|��I�})���ޗ���;9�G���<9�'S�W�޷�~���!�]y�ݷ�o�����~��]�޸KK�sØ�ט~�+C��n_����5�7�z���{�Δܧ|�}'����z_g�5�y�+�G~k�����^�����]u���>���zN��9	��'����=��u!�:|���Z��7&�:���䛷.���'����S�#��{��O�S�1�3���U����"_�rd�9�r�>��A��_��bj^��|u�PK��x��j�a��p�a�7��ߘ�'��n�Чއ1O��˧�YU�_uӂ�k�/P{��5I��<�����%˖���}>փ��/����:�wҞ=c�%��O;�;��Z����z�G��s}����WA��gG�}��]��k����p~���>�Ԝ7��^���ry{ť��~�s��i�ϴ����b}.��>:�PI���FE����G����� ί���SP���{��;���GR���f�������y���yӹ^��}��?�|�>�hr9ߜ������C�zg4���w��I��RL��W��A�e�g��ن���u,����!䗐�W�s�Yk�%h�7��v;Ht���Y ��*c�|�N�u�X8�駽�"Z��1�Lʉ�gCe�r�*@�רӫK5���c<a��������F,�O,u,x35"�G��Y�)&���G0�
8U�Snf]������{� �aq�T�>V��B�b�7YM#��Kmi�JQ�{wϳ0��S��>�,���qʴ�'	����i�G���jT��v7q=�4�N����3~����oB��N���i��$ͬ�b�g3ܣ�k{-��(r�Ż�To�x������{ՌFs2ԣ�J]l���W]�z�n3��N噆�s8�7ُ�`Z��D�"^@����u��p��'i���V�r���R�c=ю��p'�2�pcJ�j��"�扃��e�����ỷ����箮��P�¯N���I�fXT`|��Fە�Q��� �f��;rdy��eY��f�m�4ZT+%E*v!�揌
�;U.uvHf�Tv�5:�VL�,��ʺ�!�+2�vT�Yb��ͮ�@�%�?��B���vv���*�!w��ԺE8e�F=G:F絼;6�G�����)�G���R�F�Ѡ���T�RH��~Lf������x��,�u���)հt���>A���M3�Ɲ�'�)<�[1ov�r\��]��� �y,�j��=�Kv�oP�\(�bի 7@q�9>��U�h'�7+~\;�$5�����d9Cd�@R�U�U�yY�N�l�Srl�a�me���,]j�֤k�����{�7}߂�``��;�p.䢖�_S�z���JJ{g��݇6ל�oV�t�h�|�l�z,9�,��؛{gv�o_y�����Mi:y�ٓ�q�Y� �K�"��- �o�m���j��镹ؕҵW��!fSn��ƭLz6D8�Z��;^k�m�G�b���9�ӧ�%�1w��%,$��z_7�7��e�|�{���!��ҥ��V�t��̮V�lU����V���i�ʲ]ԧ5x8�l�b�B�v}oH*�gM�֥��GǶ���J�m�$�]EJn��?���.7�:�%��\��Ҏt�J�Yw�^�t��0	��[c*��d��f/��u��6����{3OV�����_SW,)�����SN�_4�x�k�rʂSc�VlC�o��J�c��R�=L�t�����lU�z��(�x��\�ײ2�+�*�#�1�wkz:W���gF�^��&H�����~#<�"VV5�c�,��p*��N���a���Nr)>T��A�g-鏓yّcO�4��(��s��TK����u��.�"�����º�˱���:m�Υ�V{a��w!���n��V��
�����F��ih�DH�+Q���nE�ˑ�G�$&Z��p�L%���96�Y�n��P ��;��am<9\Е0jޥ��7OK�a�}C���z�r�AE{�d4ĕPD�E�S2TTD�DM%��11Tj�)� �h�� �"��
hJ��udHU�D҅�D�3D5SD�DECUS5UTQDE0CN�(* 56�2���
"*��j*������j"��)����"�2h�&��J�(���f��)(*�H�)�""3X��h�bcE4UT�RUSE5QQIULT�fE@PD��QM5BP�TCQ4LLP�T�D��U�ČCA3L�5Z���j�(��f(�������"�����h�
��&)$%��*����9U,�	3Q4UIEDRDRI0PARNfDQM14QSEDQEfMQfd�RUQT�H�T�$T�ED�TU%144APRT�PUFYQUDV�$��Y�LM�ʪ&��(��*i��)b(���*kXd�YM��EEAED�^g��h��r��mi������*��
삖su���5n]Y���TL�Γ}��an�O�v-\B��d���������;���N������,�0�?B*?Jy!�c��}���s�K��}���ԝ�|�{�+o�-.[��9�'p/9���������k���߽s�wϷ���Y�-���h=���SQBw;��}�-)���e�Hvf$�\����Srr^���J��s����/��:ZZ���s��{ߙ�/;�{��������\N�2^�Ç5�;��/1��z� �NG�����>�����;�>a�N�:<�ܜ�'�vf!�i}�jW���Ώ<���{�����[�ږ��\��c���c�������i:��7��ZНB}�sO#���������]�Ogp{����y=�a��N�:��C�Ԟ��g���LZ/;�
�口Ц=3�}��F}�����:����K욍Htsz!2N_��ZНB}2��N���'���^O���#�=�����]�ou�Sx��P�dX��o�?>��?��`��}��i~�'O��˯��J���:^@�y��5���;����?��!��ٜ�O�����ܹ{&,����c�3b�q}]=ˠ(��s�9�z�����Կ��ϰܴ>܇p�u���h�	����>��sx�I�ԇ�>��N���ZC��x��$u�8�P��$�	�D9��|�9�/$��c��ܴ�<���� �����x/o��%���旨I�9�4�p������S�=9��~��E-�ϔ�-?>��;Mt닢���2u��5��y+������?@y�'r��?O~�;��^a�����?o����ܛ�K�`�	�=��9ף�1����Ȋ��3�q�sg���d���8�K��:��xoZܯ�{֓��վ�?KոMIܴ����M@rM���ⴝc�~����!�ß{մ���G�#�L�$uVި��=�Y�,il7�]Y���9��8�x��� :c�];���X����H�;��k���ɝ���}.����;�7+Q�8@�] [N��g�\�k�[
��uy��:�^ڜ7w�=���v�z�:��U�=s�/��<���N��}'�z��=�rd���+ܛ�L擫��G��AԾF�5r�������'O�~������4]�?��Y~ܽ��ԑz������7�9'��/a��>��;�y�)�S���I�?C���ɐ���\��Gg��}nW���:��`>u��2}��A����s�<%m��3񛿣ѓ'�trG��0䛍�{�}���Oe>��Ú���;����)=�'�=�oKKC���:л����r9�9������{��_������u9ܞ��u!�'�8�7~����>���Oc�O�s俍�Ν��'g:���@��h��\���4���\�\9����:3w~�W6�obԫ��`��sZO}�i��i>��Ҟ=e	䛏����NO.����}��y����{/F����Rw���럧����7a���q��^|�>v{*����#�o������4������N�֓�9Jj)��~��0hgwG��S���y.O�w��C�G��I�_�
��7���I��=��#ܼ5κ_/�|3~t4��!޷��%���`4����r?H�'}u��Mǲ�w�<�s�<���w{>���}蓽���ȷUU�Z�R����!O����
C�hy���ԯ!�5���G�ޗ�y�C�_�=@d��ǚ֔�蹏/�=I�{<��O�]�o9�Ϡ������{��>U��g�>]���z�Bu�ɹr�?�9-/��֤r��Η^����-H|kz{��9�3�'���?@�>��%M��Vw��Y|�]+(����+�w��O$�u>J�~������y/#Rto�9i��t-�Ϲ���GS���_d�jC���H`��
�J�o�qJ�t��S�����t҈���7$��J�.<~t��;ǆq�n���I<�@z��Qd�|�D�(N
��#|�XVMtj��j�R��6c��o�f:��4&P�6�Հ�d<��D�Qܙ�X6#�.�{�f.�/g�WT�-/wDG���Iw�͵��G�}���Jw/�krw.O�`��p{��w'��j^^��}�!��x���5�u���b�<�:Ocg��>ûz��U�>�)b�
�O��Ϡ�jC��Jd����Z�O��P{���`�O%����ܴ�Gһ����w�=�u�9���x��s�逨_�
*aD�k;>�AQ`��y�s�����GS��}��ԇo?h����{޴���]�s��^���y'���e7-����G!��9>�#���^9��?L�����©8#'�1�=_��9���~�9��#�'|��N����}�}��Ի�9��~����O�^�z�I�^��y�'p��?Oz=�s�L�3�~��33>��ߝq�S��7P�<���1]��ɸ�;�/R������M���w��>��Nw�7&K�����|�q�5��y#�y�Ϣ���s���8Ƈl���Ou�P���'>�5��1����ܛ����!�?G�v��A���7>c���~O�_�*yF\�n.���o&�?�Tں��9�����TZHT^�M�wv�qs�,R���[I�7{��3����\���"�ߪ��Ս��Օ�����]���m��ņ���Ҝ�v�����m0���lﲇE����~��y�n�jvk���]�=]��˟�S{�ߛ��ɥ�Lk�1kj��ZA`� ��<�~$�V�� f|2��A����}˦�l��n�O�n��=G�i9G� 	�|�3�Sۘ��zj�P1���!|�f��(���3�^Z5#����Q��(�;6������]��l��F�c����
�Njjw�pb�N�]}FrqH{>_�U}�}�+oK��B�}�
��U�X�
�R�7R���>��ƼN,"Aq�{-�P�T��e{ڨd���=+��ĕ�mu���)_��qM����ց��9,�����j�5�/إ�q����5����5�w���<F/%�Ws٧k[�����ݺ�����1��Ё�Q#ݪ:�C�PN����Ԓ�V+���x]r�g7}.:����v
�5��"/JĪ��Q��8sB��sY��`�lM�N�H��mmR�e,}B��K}��u*�����Wc�+6� a[��Ou_ӽ��7J�9nS<��Y�U�V%��	��wBn QdC�z��oW�ӷ���yF��s�}#F�2f!Dk�/K���[���Ǚ�}X�E�����OSiC��rf����aA�t�ɢɪ��e��Q�*;�7���sJ��W���W��1�lU��q����U�сc �����	O�X�����EPL5����d�Ա��6������\�n��]l�k/*u<��I���]���<�X9����r�C*T�I�X08����<_:���P�ܑ:��B�7\�,-$��I} g��t2��}�z#�z��ߜ�..�U�?��Z��+mѵd�W�}|��B��/�M[���V�$��;�G�Zz�g�s-��:�V5���ު=����nEze��kyUVݐ2�mT<�[��Q��גaF�ŝ����#�����a�\�iAWySk\Kj�U�|_����%��%Qf8�}�.{��=ݨ���������c2uc�g�p��;���T�Kg%ֹ���y��j�ܘN^a��n ž�Ź�k��v�S�Cl[5����n�bK��DT �3�|+���O}��]�m9u�d�����
Qf�R����PM��@��ƬB�}pږ�%���W#K��M�7�y��	^�|����������ȼ�%@N�6�U�~�t.>j�*�JC��o�un�7_�9Q������� -\�s�]��2��������	yhj�+�#g��2�H^JK�=������]��٩X��8�漎�O��^�C6w���X:�W�SѸ:��ox�õ�Imp���G��Xj�G���7��r��4��ݡ�݉{�K\��<��ม�XN;���BgG���W�}�E��ͷ�^&�\�odpYZ�B+u���� ^�r��ڽ��2��[5R86�����(�WU��L=�C�u睻�MR����l]6a���
�tnE׸w������P"�ɍz��v�=�N�3��I�M�S`���Q�����q�UԬ�w`y|�ŭb��8'1�IG<Q��w�4��}M��r���:�0�UVn������Ur�/���f�i�LTZJ�-�~A�8�ֺge�d�ct^ͽ11�nbLa�[O��n�֒��M��Lv��=V��
$D���1�=9%S��x�ѐ�\C�������5<�Ք��L�u�q��
)�4�)̘��wy�ʧ`�boB��E-ۦ�a��Ǚ��+�7pfYwd�Xߝel3����Gj�^�ͯc�9G�ѥ�Kʼm��;O��\jdI<��P���Ĥ�G0�u;�tg�I��:'֦0pY��wl�������2�c��k'��Z]��g�Rs�����jh�B�ث�8�j���㫮��!rRp������󼔱��(qR6<W`=qj�%��q���{���]��7yP5#��#j�*��V�tS���i=���.�Mf��4k�d���ӊ:O�|th�ȣW���\L-�:�U�6�;�U:�Pfo��̒i^nk�#S��ls��ǀ��\��J�x��:p)�H���ݱP޽��LHo��-}^�z�N�y�h_z 'dM2���wjo���u��%�΍���y҇������`�p.�7;y�o��]rIR��/��� b쎯!�^��p]�V(��8,�����aUe������#�����Y����dSC�������[#��
��Yw��[tR~a�'Oz;y�3��4+�;r�<iWR��p���M�]�7�ۻ�Y��hFr�Y�{��#O/[U��Jd�����h֋�7,w��"�j���n���A���sJ��W�O��L�^>��?Ar���vۡ�9[5�;��͵c�֭wv��.�Y�n@�Ղ��i*.��.B��1�b�o!�������<ͳ�cO6dJZ��S�ܷ�=4����9s�����X��Vu%z��è�=A���P�w��ݾ�V�������Sk[�d�Q����i�L��
�:�o��c�e�]x��]�Qۻ�3O�̪�Tl�ѫn�w�>�����՛sVz�H���8VB���-��^���z���Y�b���0b���q��߽�N؛�tk=;.��S�k��&���Y���'���>M��!����Uwa��h��=����X<�n�tS�]�����'�KU�z`�E�X���EC'�?�J�F��O8��]Oo�_��޾���4ܚN"_i���Ǘ�Q�#��;ݬ:��23f�;�.s��'�_(�>�J��w�����)����\���q;F�[��Q}��F�\҄�T>� �r��mz\u�*y���[.�f�6nv�����%Aé���(1�`�}��#�ͨ��YT�޺A�Ꮘz=�+ ���;�Go��eb�\�H�t�*y1{ ���x�tV>��dNɌo�BZ�R!�;'wݽ7,[̜�X΍�n����P��5'2�y������.S�W��(�2�R��n�q�Ռ-��q=��H�Ng
���p�����B��je����0񎵰����'���E��X�o��Wg=�
d��a{��J� ��3XՓO\Ϻ\�e����of�}۔��*�+"C<3y&��Y���\��jV(|�^�����F��mW�)��wQ���ˌ��71��1�k�Sr�'�j"����.�FE��sJ��G:x�7J�[3����|ھ�w6bY�S�nd�֮'JۇF����E󪈴��H�]��W.�}��N����Bm���a�!3@��X��x���{-����H~�2��JE�2i�|�5�4C{]x�e�Z�Tʃ:�6u_qڄ]w�u���&�eU8�D%�:��jō��{&��s��v6�T��g�[���|3r�b���*/N�}��g�`���5}ϥt�l�p��,|��SI���:��[ꋌY�w��v�ʧh����x����E��M�ʅKi@��g_�sr��6�Y����O�V��oELƭ�/1�B�=�;�n�+��v~�����u�*����x���t~�{��YN�����l�)dk��[�8�л�t�Ws8���j��}�+������Z�M1����}_G�v���{�r�mw�q q����|hj��N��i˗\�UXNenge�w�K��	%�cz����0���J��[���,�z�V���+5�X� ���;�{��0����j�������mz���.h��D�S��{���E��|Ŋ�>�5r:���|l��\c��\��T�F�x����1�WK����P����4�CV!�(o��j^y��-���l���<�+'+آޮ�];�e��A���st,1�Y�(�qg�k����NwHVqx�>��P"����U�'@�����g9�:�v<͋��w���v�8�xsG�&#�i���ϯ���|��I)�wt��4�����i��Jg��W,�DR	+�Ė^��V��̸��:��9;�ǳ{�����wCT��ŝ�}��z/s�'ܩY����6]�� f���x��I1;1�m�7\vS������'/���H��ٽ{l�	<�h��O���P���k%��d��B	�a[x#�i.a�XC,Z�v8c�6]�/^lX���\�-5]+/�֒��	����0�}W��E�d]a��r�lir�����;5�S��)V-P`j�;T%	���)a��4"EovUhKqwl,�I[�'�\nn�(%Jh;�r���N��j�{�v�HZ̰�}4.����ʃ5�4�T�y���[���Wd��C:�_u�ujv#"v`2���b���� �Vw�֠�	6:�����)����M���uwH��P��v�l6\i+x<�jC(��k��Y����s��o~���
K�+�b��p�Yc��^c�����Κ��A�&��E���k�-�@��u��C��%�9��T��йV|%o�����������HGµ��
EY�.Yj]՚kf��LyP�d�9���3�#J��Zbc��rn`��#�,>���ǩ���X_XKA�w�[�WT̊��Z�����8Xx�b��5f��[`�2B޺ɥ��8�Y�tN�Nu?���خ�Ǳ�����2yc�.!�ޞ9�S�`�mM�uc�R]*>��2(�n�	~ʁ�k8R�Y溺���m��m=�3F�l�]��ε��@�F�ڣ�~og��H�2K�>c%�=�8��6TK��{�G�H� �\�o�G��ĵ��O��S�ڰn˙��zX��x\�����Ys��s��Թ�@}p�V�]�ʾ�ˍgn�\}8�9��xt�%ƖFT�Og�u���0+��(e�G|��m�0���[N�gwS�5✇o ݵ5�W������*u�睩��Yv�Bˤ�蓮6��%�����F�tw���<��e�sB����xZs��
[��n;���U���"�'Y�Q���R�:x�	�J�����Ջ\��Ʋ�
�aVD(Ŗ��B��e�>����W���=�N�����5gJr�W��`��rsr�7�'Z����4iq[�$����f�m�"�#�J�y)�ڷ]�k����^q]�һ�UD���|��W,���S���.���E-����u��Ɍf�ݰͧv�KW&�I����K��#��ō��|�+w��&=�Lݑ:;R��OY6�n��O�V���W9�gX�ܽ����'�Z�=�F>�mԿ��w�>�)KM_,nڳG������iu��A�ZE�ճ0�/ 
����ѻ��P#N��ף1��~h��p�(V!�x^�$�^�e��/m�v+�	"nƽB�h�]ū���ˈ�;|6#��+��n��A��D�P��yq�.�[�O1R����̏�My�՞	!�3$�A��"6��m���n^D�+&�r2�e1�N]��+t=�%�L)W%��f���8��)�.u���}�n[�p��9�Ǹ����d��$H?A.�*
""!�(� ��J&�"����������,��*"�`cPEEAjƨ����
)�
����X��3*(�(��	����$�(��ETլ��"�"�3"*j"��b���d������,�	(����%ԙRD��HT�%AQjɘ�")�r5�����33#�"������*i��c0��*���
��*)��!��"����j�35&�����j"H���`��&���ՅD�YEEQ�Ȩ�b��IAT��EUTTE2STQ11TĔZ������&�*���Y�SE�4�d�A��CE�CVfE�
&���Xe�cUQfd��1L6�ʊ"(bJ�h�aE4CT��Ȋ �&�����E�TUTU1�|���B+��;��U���Y��<��C�pl�ƫ3�g}�o]ͳ�,��O��d�#��n _Nא�^�Y!�E����������ʷ��V�1�9���M��Lv��q��k�:x��}᷹��69{73��\ \/��m�EW�^�O.3VRƍz����'�U+v�d�تۦYpd�6��C��F����{{N�y��])
�Wv�y|N�ԢEU��p�V¸��ߛ�X��Zrע)v��ǑL�|��W��wr�Ʈ{�9�H�,S^�p�De+b8�>4N,�V���n޵�{��ȓUur`���㵆е,+b�j��-���F!�z\u���s�ڳ�Y�̸Ǯ�H1��1���	Z��W.fnh8�<
V��L٧��>���k6��e{��g+T0|�H�'!�*�\|�R���v�@����g�a/cF����+����{ ��޹��T�`�V�ޮ�H�n�u��ߩ&<ĺ��S��:h\��^l�im��c�b��ɂ :�������,��Ι�)vs���ؗLd��M�f_l�pj
��.,gOs�Up��y����qǸ��.���'{��%���C7�p�l\�2k��Rd�y��o	�Hd�k���)W�n����ȏ�ގ��ASpFL���Պ������A���k��R��e7����j����CSCI�~o�0����D<廐�4+�c�-��)��0�����`�Y0J_8>լW$�y~��C��qҙS������0.�15�n���vn�y|��HW4���+�O�.(�'}�{�r�6��2��ȭ��Q�d�Fz�4�������5[j��z�r��{m۹U6i�K�JeS*�S^ѫn	��ު=�߽�ܗ�jڳ�:��&'�/�&�כ�Og%��%Qg���+�5m���]p�t��ѹ<�[��i@�Bs=/c�:�SڎX���H��6�}���y��*:�ou�}("(��Oذ����u��XR�X=`�3%�K7^a7 �e��6��1*�Ew;�F#ދ'�`=(v���l.����2e\��:hW.�F�_}�ygV����e��S{[��4-4�o�%n���'S�w&�)K$��Pt�s-Z�ԍ��Jvb�/�����2��vwk Mh]S�,�.�7��J�kg��XP�9�gT�
���W,!bvG�J�J��ѐn�w興���L���C�}�F��X������9�v�ƆVÖ�����˫맪�=ɀ���*���Y<�����xg�)�wV۽�|�:�^���,P��a��)����3��9���>:D���Y�/{Ne��r*�V��Q��C����0>�}�lM���I3U�m)��#���$��%y�����.�P�eiX�Ђ�-��3��&&�V�-�S��m�f"���bk0���S�1@���j�pX����|��n�Dr� �Zs��0
�vڍ�*�V�@�P{���.�P=|���Ғ@�~M���Q\)y��n�1���R��;8�{S���'�n8jM��>�Qi1��b�>�7g�TK�s%T7j����4�Je��o�Ѵ%�3�|�H����/���6}I���;��׮6y�2��5e���ǚ�A�z��ZX*̈�������eHÌW�ͼiǗL�_�lNZ��x7��&`E|�K4 t�d��&/�®�aA��r�[j�[�m8�#<�YTS�9p�(�%��N��2����ٻ3�yZV'�Y��A���/"t�j�}�4�J9.��-�G4����y�����l캋^J�Pbu�[�M�GG����m�{�H��^�N�#�bƏ3���K��䠸�κv��}{����	��^���b��]b������.�r��fc#����m n�'c���ĞFw^�4��:��ž�ž�{'vSqbp�^���&��j�N��9�������}1�|����4�� �7�B��ʓw��u���Nz�`\cX�2�l5U~�D?-����+�~���n3�/$e���I�2�B�v�'�XȨk -\��2�^A�SڹWYOwS�Yg��v��U��F�@�,N�,T=�W��w�	Rw���`�����˂�r���:��W��:�>V�{��p��j�bּ�D:�M ������:��b�oU{�����e�G�`�eQ=�-i�� �a|�����*��/]B*���.���\#� :�nF"�}p�_Z[,�}ן���`	/���%�e�	����̺�tevr�:_N���k���E��2ԕ�8_kVEӝ��4B�%w`������ح%[S"�c#�õ�z"9�Ԛ��{�C{���Uy�H�c��Y[f��(�Nߟ0+���cu��u�=��j{ټϚwQ9n�*�	���`�*�B��c����a���ii���!Ԣ?7�W�$�Ѝ7~�����;S%�r��E'Y�i�!�_^�i��Dŗ�9��iJ�]>�qs�)����d{:�H��r�.vm�l�\v�ȼ�2�n�;�'ӊ|k�p��W
{lb!>��ݶ�2��卜��s�ѫD�{�0U{٩��jō��p�S�[x�b7Gh��쪵��qa�Thբ)hlm(�X�KM�wϙ��w���q�]+��+����q�����{f-uE�-Ox��nKF�a�<e.��rf�-J�`��+�J؎14�����$C�a��3+;��������}N��������Q�F��mu��ѝa*���Eɾ�O\�� s��dj���L�a���V*w$I���R���W$+2�R�5>B�h���c�x�Cg�C�F�����q���VhqX�K��)#ү��]c>v��q��C;�J�F/vZ|}�� �⦍a���e5�k�1����u��ʈ��ޮ�o*���?@���f,y�v� ��I��dSXƩ�ՎV%�sx��ۦv��㧖�������S��N/:J^i�×˟]R�\,?'��)X��tM֦c*���'{�Y���Lhk#h����gpp�A��� ��P�mDK�Ͳ�[��5=���|D�tz.���w�m�{|:���l,{����EjƼ^V��,�
��b�b&��V�+��&L&9ot�{��[�t��*�
�ܿ0f{RU���1�ķ<P��z�צ�.�|��V�Q�$��mTC��r)�S闙]*o���Z�9KY4Y5\�,���j��Y/"/�E��G4��W�dY�֍�Z�M)�T.�p�L!�+F��tq_���(u�i$^�{=G(vZ��h�G���ת2zҙ]eA����ge�W��{Av��j�ۊ�Dh��h�橏z����gvC�.�<�Jf���Y��$C{�.ҥ��D;�o�Y�+�%y�u��B59���X��]�u
:�JE#2�Z;��y��v�����_yV�0x��zj��L2vd��T3L]OB�g��}]��{�U�d��x���o�=���o�X�r�%0���fW��1q�nV��%m��d����j�2L1s��6�}�v-��!�k��/+V�_:��gذ�s�4G�y쿔�������+ޛ�n��M��Y��7ԗ��(\�c�Q���ד�)�]A�g����uҶ�1�:)P��3�qº�mq��*b��(�0�NFr��U#' |�m�fM��@���޴6T��Է�q^Q�ud���� �p�QV�Q��������vEa�7�P�fm��`����_���K��h�1�������$k�u�yrpa��� /nGS��3jzE\QY9n��-��i�Մ	���r_<}.�㳼��zK&�YW8t��}̭���+8N�Qo^p�ߠ�����O(�����L��r�{*v'y�]Д����z�i� �t*�Vs!z8I3���!�[u'��W�}�oƂJ��e��Z{�U�������/�z�����Me�J�3	V��j��$)�lz�O�:�'��{|(#������Y���Zzw� bŬͪ�F�}����<B������A׮�8$�{��eؼ� ������m��w&��Sk�5^?�p�ڑ��_(1�8)������]j0���f��}ͧ�:s<�Z��Ҷ�ѵd�Fz%`��-���\#C4�LZ}�I�,�ͱ�a�!3@��Cw�u�{w��y��ӻb�[^z��
FǒY~�N�h0��-�����2�^������x� Z��<�-��#vTN�wڲ���L�u���bGB_,�ۼ\r��>X�[к*4k�1kl���ά}��pn�n�]��q�i�j��
�Ъ��d�<��/����sX����յ�Q9�؃^}^�"�����N���(q���WT��P5e��3}�i���w.zB�7�X����cr(䡐ձ<%� �7ף^,�*u��o�wמ�^�-\��h����-�y��~���<H[(�M��x��7� d��ՙ"h�[y֞����G��t�k�����z��^���G���,5[�Ǝ0�:jc�2��kʊIy���u�p'��-+�i�5CAYj�܎w����D%O�9Js$�W���Dn�cT0c��%k`�6�U��uK�3�Η�қl��孮��4�Y���@�'1b�������
��v������F�]�W9�������:�0��X���-��@�ϒT+�����S�<�5��+[_.��ʠ}/��tn;6sZ�ec�/nA&�����3Sn�n-�K�}Q��l�D��T����z��2�Nm[4��w^y�w!VhW�㑫9��T�n�{�{�u��q��<�F՗�N���.F��p}P�zw���Z�`���ˬiB,�O�#�靭�������I
}��W�A�F8�چ�ʠ��*J��a���|)�mB�Y�,pE�t8Ů����55����#+���*�dܑ:ywa� ��s\(b�8s�b������5f��������W@�y����o�R"y��:N���c�>ZI��9��h���4ךe3�*f��d��Pq�v�3L���d�j��3w޴fɐ��N�x�S���)�mћ��QG�Ǖ���JT񇧙)�Et���ȷ^�7u���׉�s#j�H��rS��ߗm������r�3��Ȓ����R�{��u�̝�o�Y㐋�
�V����q�Zi�{pb�8�����k:wq�O����\�M�6ϼެ�%�*垸b�I�v�>2�;x�z��yc�s�S�K+��EC'�0x-Ȥ�����P8�B�1P;
���K���Iľ�;׆����[�NA�8ڄ��g���-̀��;9p*X��`*����v��ͮ�:��V~>��_ܹa�����'M�|Q�W4��x,W���Z�6�.:��T�F�pүhy������ufv�|xt#66)��Z�	4���Xs���I3Y�kj�S�T)�t��ܣm�>t	�3\0񎴥bX�o4S�uw/+Y#y@<bv��b\�ݳ&Sn-������;}o��<廊�B�c���e�H�
'wkʭ�����M^��PΡ7MAt`1	%�E�p�:>k.,�:):�<O=�wQ�7<T��R�·-˫mX�����|c0h�+5�GjS3(;U���[`���w�e>\��U������L���@���h�0�0\۫	ֵ�9j�B�:�K0�3]Z��6�yf�<9N��%9&�j	�{�v5���}0�@g]�i��'��&ٚ8���̭upr]A�:�(��
E��;�1M���}�tp-Nh�+NV�8��[h#�Hva�᭳���`P�M:O�|�.��h�;�WL���DD����)����S��|5CS
Tr1p%SU�����ĳ$�\��������AjN�˒�v�-vU�<C��xU�����Ν�#p.���>�Tsr��s �i�;{�j�o[t�zs>Ԯ�k�uW���A%t��ޡ{�e�Dt�
2&����b{�M7��K-N�u�f�t������Y*-�{�ij��V�cv/y���Bn�itj���t�(Fv�9���:b-�kEo[�d[�s[Qr�>��n����Ifڬ������hX2QɂhגG2���-ǜ���wr]�ak곎M	�\����A O�cg�\��b�-�����A:�ʋU5{/�e!P����M�m+&�tk;H��ʍu����K�^A��+�=�����5��J۷���!b��Ժ�� ��	�Y�L��qk��Vl͛R��]��|o�rL��Ww.N�#�f�1U�Ff���:�lW�la`����7X_wd`�`��1 ���״q9%[��:��O]�=�D��?�"�.Rŀxo����}���K���ʜ6#y��.�]ki����t����7��۵�<��|Q�b�y�D{ a���`�}b�$�F&�M^a����Ё7�w1��0uW���-OK�\b���u#�(X�]�R���0�z�����]��n��Q=+�]sV�OUA+���@_e�.����}�p��(�v��:y&2���޵�e�ݡ.H���X�p���L���Uev�P7t����y�dԥҺ���Eu�7�+.�띨�j�TZ)�U��D���E\��P�\���j���eh�w*dr<<�2.K��Uk܇�aw6�7��6�U�n�Z�1�0gZNþ� U��X��[�(�6����ĢX���b��zAX���%v���x��7��iմDgv\i�v���:�\�CT)H�3�l�K����kJ�0���e�&� )c(V�`	umfe,$��&���6M�KvT�c����4����f��/��mQA��ov=u��S}}ي��r�)AeŚ�RYg�w,�͡�-�+�҂���P�
Ǎѡ2m ȗ���OXN\z��k7R��Wn����u�qǺ��3��vbE�ί�3h%��jasWU���ss��G�\�w��~�h���fXPSPKST�Fc`ѕCILM�dE�UEQQZ��h!�"���u�Q-%EZ�5�Z�����J��kVF��"j���a�fEKTZ��c#V�H��`�d�T�FfD�T15U34fS�PQ14IY�-UTIQFU0U4Qf�1UddDTEU�dES5IDIQ�VfL�cY8PD�T�U�1TMFf5��QT�8�a�U�ED�Vfda��YdU�LIL�XSM���U�E50SD�S�dE1VY!�8��%U&Y1TPMSLQY�PATVc��E3%D�A���W�����w֓[��5�u���ysO�4�5PJ0./{Pks���o�0���:��SQP��<��!�M��F��@������C��;�u�����F(��b�9%^F�kk��L�u��6-��C�w�{Y���\OX�Om�6��U�Pb�B��*G{���^�z-^{�{�F%ܚ���nR�����u�e���/Fӳw��Y�Êۺ��<�4�tk���ZS*��Cqx���+�m���1��yHq�܍H��M6���X����NJv��E����ѫj�i�l�ȝ��guf'ȃt"�{H�%�:��G;Vt縺w�K�~n�,Gn󴂋��
�Ws�t���>�~1kj.1xbuc�u�ʹ��%\j��O�����3�d{����I�͈���PN<��\b9�k��O"Po ��0��}z����W��*�8e���o��k�5�/��F'!Ft歋��n��]��tR��6���	c����7�O?�����U%җg�(����ZV��!��f�n�pJN���ws��\��¼4��B��.�r[��.����W��.j�]�g�E��m�ϔ�"k*iǔ���ԧY��﮶+ }�>(��Zqd�ܩ�W8�󹝅E���K��t�UX>���tOk�Z��y� gY�i{���1Uc,�8�f�2)QGK�4�ܭP�\rp_<�~��ڑ��3s/B�(	�jo0�H�y�s��b0�಴�jPT�G'�-�ќ�8f`�ƥU.����*9#��A�
��[�ӫ�[i����2`Y���v�bjs��Y�[�48}ۗ!q�5�_(>׮��I��*�J��n��j�I��s����:�
�[�,��)l��3��oy�~O�o��' c��P�r���O
^v�LBj�J�E-�6���� ��꾝d3;v_��U������w/��\l�y�2�Ptj����40�~�<dΛ)J�S��u�( ��1������峒�ג;.�R������}ӡ�c������g��|eD�w}�*4i����l37s��T@]n%Wɔ/���f���H����1��r����EK�牃/����G'��,#�6]�Ÿb�`�yW�[��7*�%�k��J�W��{�fI󙼮�>���a;�ko%G7Ev��ͼh�ުOnT�vG�
U�_���2>~���I�W��S�ʝ~��yJ�<�.u�T�zJ�[��,���V��
n�w#�^�����/�m|_m@��eCK���Sx��b,���4ܒ��Cl[R���R�b��m�YF�7WVғ'[�"rv�Z�I����*�����܊1%/;�?�ћ%X'��3]u�a��):N�p�s=�R4���t��1�v�&��^k 0�����^�5$^Xb'7{��`���\to/�"�4�5��p��X<�|Ł�[�-�� ӲN^���h������+˂�r���՞�+\c� ���[�48�2s��ʥ�٬��L�]֖	�V������ʈ�ުᩱ7Nq��d�{��xR�9[>��̏g�3=&jsvE��!Y�5�+�읇�*[϶K�S��C|鄝�4��7o9fr�М����Z���_-c��9���6����vM��ĭ{	�o"
���,p	ɧ8諈�}9�Jr�����¨�v�A���nǞ����U{o(���'\�N�g�������{��y�u�h<�G%v��
;ܵÖS�'wڵ�/�����u�Ϣ#w����� /�F���Z�{�U�7q��y���yڙ(u���e�Ƈ��v���{qx�����n���Qm*y\ ��������j�cys}ۙJ�S-��Z5��*/o�ZW:���ޱ����͍Xxα�����^K�1��N2]Z�Uʃ�T�hբi2{�.����ޱ٦T�7��6E���i��X��C�1s��.���Mb��f��}�t�Hƌ7��J�R��3HO���ds®���ؕ�*��u�f���:�^ևn:�`ԽI.r��b����a�s�)��n�3n�\1AJ��vvM����3��F�P��7�f�+�F���ד���Xt��7ୀTv���k�=Ĺ��Tɹ\��;�hj�5�/��W�H��g���Bx�2�N�鮥/�g%�mY�<Bx��ץ��@�n�V�����^�i���"|/�����i[K%�j�:���K���^�j�hZ��]׃c�����5L�wA�f�>���ߦ/yUm�:S�}�z�bk�<�&�e��dv�y4MIxF]8�gj.���W[�U������uQ���k7w�%��irU�Z}�wj���x�K$O��䅊��j����q�(�j}����Q�ٲn��mr�J�q�Q�҆y[�<�o��#�͇zM�g@r�gG43��˳��i��9pew��Amyc���t\7�)�H��C��4p)y_^$�	��.�1@�['^��߹��Ν�f/*�	��bQ�$^�a�8�\�d�k@�^�WS�A�}X��Eƭc�\�<�mN��j��7^.\�h���U�κeN�Ȗ^ڣj��Y/=|��HsJ����EElݒN>y�Pݪ=��k���J�v�T�ѫoΎ+�&Һ}i�W:���e[�TNݐ04�S|����z�'�)��ʃ�T֍[d_2Ü{�����Oh�Y+=A{w��r)��M��__�s����	��zM/�Sցwb'3�WH��Q:��s����GN��Ļ~mǧ=o8`��'F,�c���Z�V�o�]_�fR.֯eock�yúT�P�+,X���#R��ɞ'�M脯
'ǰT��C� �n��������Ք�d�ީ)`�����g��-�kcK�U�J��W\�A�{i�H�m��9.wL���_�U/7舓�7S�]W&��"��VY�[^�ŏ2uc�g�s��S��.��<��G�Jy�+<ji_\�U;ү�����ډM�"���F����Urt�ٰ�
�e''�m���,��+���H�Wl��6���&��JӔ���K�������2o�|�y���
�L-	s��)����T�� �.���p���&�*��'� ����h�{���-�3V�Գf�TS89Ԫ�7�9�hm��|����޴*�o9q���ݷ�ê�����+wQ���`�W7����ON�
zBLʦ��
��r��y
�u�p_\��j��o��g�}���@��w�7���po�h�d��#����]@ά���nɻˮE��v�Ĝ����4�cu��[��m£j�n;���Ml����<��r�d,m��>ZW����FV�們��mNwj�J|�s��%Kǩ��g-�>��)�G���'�g'�
�s����� �<_1�DqǦ�U�����<*�@L��Ի-n�ү���յ˭.U!T�8m1P�T�r������nd�֮"t���F՞΋N��f�I�gN���~������\�ě���܃�t	!1�p�^��2���ӵ�FB�Dv?|�"���X�{ɿ��;W�C̝�~�lvYq��9��,l�݃��d_+�g�q�N�ez4Z�&*�䁈�]Uט�iʭ���{*�k�W��F��xEvU�T^F��ǆ�.C��MM�</N�����C���`�H��4>����t/)�۴͠Z&W�	ˋ:O(���ϕ6�=�pġ)o��14��Yc�9c4��Tj�Y4k����o�3��X���2ՀtXXze��Ξ�?��k(�H��&��5k/�^� �`����$��2)����ҕOkֲ�<ޞ9J�'����m�:EWY�Q��F�a9����5�����=t�e�(Ywjt����������nA�<5{n����-^tU#O�-�w����`HQCn�-��y2�����U��W�rT���'�}*�.3�C(Z}6�KM��ΪY���@���fesk�*{kt�ɑ�����.Ѽ/ː���tz�A:Oj�[�����x���@���Y��qזU�Tb{[EMq/�3�t�Ŕ�f��]���¶|Cyq^��N5ZI�|zAF�D�}�7���$E��\�[;b8U�[�]UIK�K�Й.yCꋚ�έѐ��m�P#����#:(��1t�O�J�$������2]a����[��A��.v�7y/D,<�+HX��� ��ɼ��XT�d�'���}4;�j˺�W/_+��Y�\RF����O6��� <\���轝c).�S$��sa��kn�������S��P׻�\�o]q��q3]�+�d�jX����HȨ=��a%��+V���*�|��K.���g-��N��KU�������GqO�f^��+��s�u�:Q��_i�U����]�	�������:&��X���yO�GE���ħ�H��M�oኳ���>�Bd�[
}��pwg��Q�)P��Z���|�ٳ�D�NAD�~L�����X��i�~����=��1���:�.��<�B�-�[w��^�ϪU��ļ�S��/C�����S4�ݼ�l�zI��Z�y7�9ཌ.c�A��#��Ρ�|�0oU��9�����S;���u��%�,.�l�9t�寖�->-��qŔ5�Wꭠ��rz1�Y-.�5�&�����x4G$�r`3�g:�on�j�H��V�f��X.=B�Wfui����T6�� R�|�t�\�K�OB٧B�"
�ie��,��͊By0Y��_�*j7MQ��qs#�=���w�0U�=L�usJ�o\M��j&�Q�g����<+�N:�3࡮y���ѿ�_?Z�{ݰ����'jG��S����V��^�O���N���ǬU2,���ͱ��nt�z�u�O�@3ˎ��%�A��CN�`>7$���@��'n%����	�Zg�;9�Xt���}�m��,�^��*��z;7��FĔ1'7Z5��)o��}���tz�*�K��&�,�*gl�F����+Y������r���cC!�ܰ���\�޳Ydt���xjoP|���U�3�)L�<��Lk�	j���"����^���'s�c6��L���tH߸��Q������n�;Hx9��wˮ���{��yJ崻�2�+n�S�Gt���0q)u��T�_<&��u�/=	N��A��%�m7���g��683��g5�33����+�"'ΑV/���c۸�t�M�ʤ�m?�h�t�{%��+(�+C��v^���LV�c��T�6�l;s��������������'8F8vk�P�	���Y%�u����sR,�"��6S��͊o�K�aWM�\��T� *�S5��Ն9�6S�ěn�]�/ޱr�u��r�J�X�������� }B�Ve˶�tҺz�|��k���3�}1Y1ug���c����b7*���wlFC}
�x˛�%��O;��N�3�0fr�B�3H�9��
�b�݃���yg�C��{���'/���ǽ{�g{i�<�B)a�V+�B}���qfkA�Vz�t~�8������Y��+WU(�R���o:����<��H��DB�#A��W�7*�q���q_]/X���$-���(ᓦ��\�m(�j�M�D�"������@�c�5;~���p�zc�]G'/����&		��fj�<�F�01p2��΢w�:�7(x�*u�f�%C44�<�Y/٩����c��;�n�O �
�LrqQ聛�zo�R�����A<[<S%����0io�X0R������h-�l[�}B���:��GS+��Z��_L�2��-�u1	�[']B:Io�&[�w7���m���*�7��C�v�c�8b���v�g�ӂXKaZ��[��]@�[�H�p�-�B�I��$�ޏ�S���@���

-=|��X��/��ψ����D��mUG~�*f$C��g��5����*�������dkl��wX��F���QYX���jUԺ�ɮ��wC������g;~&�T��X��1�Vp���g��s�kݼs;�j	n�<��Л�5"�U�ɤ^wk���i�YK�g�\�;)�<���Q�o_3VD3�M�v��]�cs%�wI��e���YINɬ@�K���Gf#L� ���WǞ>���Տ��b�
Yu�A�{'ds�:sa�[����B��ΰc��OP87gRM������{�\|��}��T�X~�.XGK�;���k*[�WaݛdcsP������J�1͡���9���c8�����}ݽ��M���� z�S(����,�MLǪ]����5N<��<�,�����F��W�k4���������z�ќқZn	����nX[���*�ZkrnTU�mwd����CIŧr��wMR�W#{*<^������ߜ��z�i��L�{�U���)*�nE�u�1�~�5z]w��hc��L8�'W����"q�;f��MtR�h}lA2u3ڣ3��/,콂��l%(V_=�����eD+A\�J��C�>��),[�vݝ�v ���ύ�ea�1ޗ��QZJզ�Ew�YK0swz�
n�5�y�Y� -�uuoV���a� H}�cT�rr�k�k���8��#b#+[�+�Ϊ}h��\�z��Ѫ:š6��ٯ6�B\����͞���c@���T�Z2Y-*+`�*�^<���z�q�ةݲ��!�DR�xC�*�K\��Q���p;%sp���݇�ɞ2���w���y�"-(E�mmrg�F���k�{+�z�;�h���i��gAy�����<�P�S�O;/c�d@��Jsk�{�bN� FO�[(]�ܼͤz��f�]]���0����L^clH2X�q.�E��vUS�Q;�/����J���'/^H���r�I:��aw������,�"	�ζb��g+"��5��2�=f���rT�PPf�:w3���!�͇8��+;Ohj�p���J�JC^��/I�v��0��mֶu���J��y�\U�L��2��a7KJï5`GI�vL5)-j�;�0�;N��XSP[�;iw<�ߣÂ�q�uďR���1�30S����T{(Fu�A\�o\��ze��Η3�2���������&�̰p�"�*��� �'((�� �js ��332i"**�"j��"�
"�*i3���*#!ʩ�(�������*����$�&�""���������
	���r�b�*�`��*�,�B&*
r�h�I�b*����������&�&���(�����()�	���խf�Rj���jH����������##"5b�QQ���4QQUD5LP�EUE$��ʊ*�"������$�������F�2���@
�
� (EO!e��w��E+� ;3/y���ˇ)��{�n(�g]Qf�7Ƿ p-$�p����]ɉ:�}ܳ����3bO���8����C�@nU�Ĵp�j��f�(�Ǒ��o;�D-��zڣ]f�����ğn�h��n!L9�^jy&0��e�s~�yD����(��RF��=�Hcy�QW�5Y�$U�3=�9*��=��`j��c�}ȗB�v��̑ܚ�I.�H6K�,.sSv�KÙ-��/ț�ԅ��,��qTo���ĺ�ݵ�`�����W���j�M��j~�[��j�`(ʝ����^��z�5�xT�Ɍ�E�}2�/���I+B���/=,���g@�p�`��lc��e�H�Tʑhd�4}�SK��n�w��Yx�����=�.��^�<���XL�xfk:o`*l�ȨA��i%�c�/|�x�3&�WTT�n㎡�{� ��0�国2<��ga�:�`oP11r�=�=LN/t�4��;%�>�K�¼�+��vg�=�K3�e	�����W�f�w�J�#��0d���D���m�q��H4��b^+�����7����^ ������u{W%F���'23������r����n9ܵ�pE��
ιc��v�{UB��)�#Q�Y�S�5����F�f�W[X���+�ۼ+]�Y�Z���bݝ������!�O��s��o���9�-\]��Z�j�w���D:�<��=l#C��^.��'���uq�[Hn��]�F�9��:���{DȻ0$Ŏ�Eip5��LK�J^%���R��ч��w���$Ք�z en!k5�����fJ�1e*8DJPs�	��.��
����fڨ:�i���� P�ڲ�R��}E��Zp��%c|@������T��&�Ы�Y.і+��UX+D�&�#�/0<�AQ�T׸���V��",�8�{�Ij��5�џ�\ROod�5ZI|:AG�D�>ʍ���|�k:�6K���P��ˍl4�S�&K�zb�^��᳼�n��\0�MF��1W�-�F�s�1�'6��A�
$�� �V�|
m
�;p����=0�l�+��������ʑ�=�|[�͓n�+7�]m�&��v�F/��ׄ-f{�H�*6e��t�9�+�t�}����=��}�y��O����	^m��h�B����Մ'u1]Xw�� ���3&��#JtZ��5s�����KW��`I�긪�fe=3CHU�YC���NM[�ڈ���,z�S��4�bK���M�1�w����ۨ*���h������íH��P�+��n>���}d�G�F��@4-z<�s�����{���J��j�pV���D�D��_*bx���t��2:�={��������?3�js�^��0�r4�<V����==6s�������2z�Ǽ��-��b,/U�:ĥ�2I��L���ջ�i��7�v3�HÝ���h�<m`c���xW���z�����g>=�J��L����hs׋;�r�����y����+Â�to�J�s�c��#ŀ�E��EW=b�K���*�I������kx�>��H��/�m_)�Nv��"��+�}���0:�eG�X��~�y�ɂ������B��������,uϭ�pu��.���_@�1��'2wn�S��'fR0&$2�m*�M�nCS&�xV��a�5��w���򼷜������S���u�����'�h(_��h��v�ZK��us䘨g;,-�6�u^��jk<���Q#,�����T4�ꄚ��
���T��(��FN���\x�V	ٛ�L ��čL9E�HLc��V�D�W�d���WWn��T�V5�t��/X����	�lj\�cy3�z�wO+�LZ���p�z�Z�M>��&�]C��j7\��6T�����8��[(+���7J�x���n�=�����6��E��;��E�c�@�P����;�Ͷc@ѕy1<�yGR�6�~j������Mk�0�0����+U��1��Ffs�*�Y�C���+0ݰK	�W���|�Z�L�/!�ݬg�z��͜��f���|��>�PȘ�ܺ��QW���c�g���:�=�Wj�����H���V�X��~��?�!��o00qc`a�'��f�e�I]�fE�u��B�]7����9�
S���B6�٬C(V����@�����β��t����R��k�==9��@�<R\���/%�z�����K�d���c)a�qD�F���W~����
a^)-��}��!Τv����)����8x��&�a��qA����J��C�����4���:���������� �D�(LDŕ�AY���_y���sȻ>*M՚M���[��]���Svk���J�B�]a��M);�LF�����+a}��-�����M��]��/����x���&tھӰ5�lr�3�6�Rwg7lӊS&��-��F�Ks+�t&Y�9�VPhcZ����BǮh�%��9]��dH}g*8'-�&ڳ+R>�W�NBY��X��Gc۞��
�w:Z�EI;5l�jlZW;�6#5�s����se�'\#R%�dÝ���l�	dܫ�Ʈ*���J������U�W'�ּ˾�M;b�oUR�v%�lnDḨ�#:���[t����c(g{�����4��v�>wV_֬��kt�ؠ2�"��M��y�<Q'[Fl�Ȟ�`�r����K��jF振c�-�T8�7e��O �A]I�qS1|��H��m��j`��U�Y5ğW�u���58'˔�[��Xޅ(��hx��(��s�V2��>$-W�q���b�w<I�7Z4_܇�U��z2(<�
�1e�sq��F���3V����;��!�����{�ʣ�u���zd�~]c��~�j�ΡD��D#fh���T�&e!�4J�7�MK��&�'Y9��x2$!���WM�1�vwW�>��+^kD�فp9>^�@�T+;�i����ܜ���VJ�Z�ܒs˵�r�5@ha���>Fo)B��7Ҥ��w*R��'�_�e,J>KTwt,va��ī4��S��ݵf���9�s�������%2]�N��r���Լab6�5��.�����D��'C.��j���X�4S���)O7��w^)X5�m��Q%�w��METX�A�3b1��J9�v?;�Wܶ��0�#=S�Kx�� u�w�"�ج:��_͍���e�=;�fL�D���7��1Ow+�Z�(Y8b��j+�Q��1�I/+b���t*\��2u7	�(��9�bI�Y7�7��500���lıV�ĥ~�P4���҄ӯ��;-1�Zt�֢XD{xr����
Y�>0)Y�;���%d��F�~�'Y��Ul�=�<�ot��wV��3��:<�U��~��OPR�6ī3,�A�%q��{%�J�7�{��'���d�p�Nn��U�l扑v`I��\ �L{���a��4�d��5b0�]]�%���S�~��tԪ9�ħ���=�Ǩ���$�v�P$�:^v+�;�6�'�T�Wq�*����J�:�0?�����.����3���(muy؃ui�]+�,X��j���
�N�UP���1����w�1�1�p^��[9���!�rv�@�����Fgz�Q���T4��KG	/F�<W�-^W��vk�
�}5���B���i�gb�38�����wk�*qF�lK�Y��{L��zƤ����ξZ����ݷwΉښ�5�.5t1�bv.��x
c4�=v�x�Tby�W��F���8I�ryu���sx�7���,A��3��vC���X��q��
,xD�yP����T�	�瞘�o:�FCgx����
�����u_k�����j"8�-0(��@:�P�p(9Rf/#��6��ѳ��+HBd�>��F��&����O�ǯa���#X�	{�!�(V���s�2�ڇI�c�N�^�/oxۮo+H�#ZIq�W�	�6�ƅ(w�+֕)7�#&�Ћ��R3�5���ܧl�H��61Y_ӫ�Lj�p:���2�X����01jco������y��Q۲(�p�a\C1��[=���^K��s��_�Y��Z�W�j��߃V�VU����u�n�E�a���cl������������/����,QV�������9��d�R����tqp�&���2S��A(u�W' �d��r���|�t�ww��5�}�C�K8�F�T� g<���X�{�z�CbѪC2�Hpl�OZ�Վn:��ό���L�`�"����yX�h;��U���g@��-���4 D�x�׾���2r�m�r<�)�D���/�]x���E"聽����Q��M�͙�o��]���Ҭ*y��;U�?z�HCw�uD���n�Ŏ
�wF��K�u�<��j��Mj��/1r�{�wl�w�Ķ�3�u&��zZ���د�5� d�Ȳ� ��I�����!<�,����8x��t�&`��48[�g1�s8��z��钕@�Z��KG%WWU�;�&�p��+��*CZ�S���Zn*��@߭43���;h����y;��|`X|,���d��vz�¨�=����X{kz��@��qs<퍿�G��(�P�(I�ӣ�
��Y$�zd�3���V�P��\��E��}oL,�V��,c�
����ܡ�Tqz���d׻��s2����y��V��5���o���X�5�}�ϲ�L�~�~�~��襆�Qg5tzb�mWU�0�7/�/!�5���oPw�N�J��\U���5�,+������.�l��0����MJ��GJ�[q��L��1hK.�5Y�C=C"Ua2�ߜ.���X�*��̸L��H�J���-]7/��	�r���P��vk�il�~��x��[��ӔX�,+��Mz�H�>LW��R��*����ǊK�o�B�N�.��T���e�3�m��+���_`*{�t�AL].�zB�2K=�.���P��
�:lk-�9�5�:yy���e��+�!R똼���̊vSu�4+WZ֎�5mey>�ax�4�?Ozh�6؋�Ҝ�%󅮘n6�	w��֚����Wت4��a�=Οbhd�iS�jD%�|3ˈ�&�ωj豷�9�U+:ek&rd�A\'dy`�!�f��]q�c���*v��&��|�}{7w���:�~Bt��^��6���h��v�Ř+n��945V����
y���0zߋ��K� �|�|��\�M);�LL+�E���+���F-���t��0v���m�Q�g�ò�u�r�2%�CuP�P�N�5!"��]�Ʈ*��
�v����u�1�)��&��l۲J�bY+�5��U��9��k-�5;�:X�03R;I�ݿr�5R7�1��������U�mC��P��g�s�J��'2h��dC'D�[���*��Zl����xݜ!؍p	
`��Ls�s����J�H��w��]W>:��>C	�경cόxޞ<���)�C��Yf��y�n���\C{��r��A�j�
��BL����yw�=A�¦M���Rl����<*%ݹ\�=�S�[5:1C�*l�R�Z�ڳf^9�@�K��� U���v��hs�p��$`@�bd�v^IM�T���=`oN�wU+��f�<�}�[#�LZ�j����߶���ɐ�[����{AY�|��ͳiv�rF�V$'ٷ��&�c������\sj����bUi�izc2�����:��/�����T=\�ɈL��%J��&���7p�:�Ǹ��:�h�n�5������}ݥ6��y|��S��{y�������������s����Q]����|;xn�v���;�
66+��gr���w~0oB��R�"Y���dU��4X��Vor���$�a��� T��g=�4��Jn�Qᡋ�s���ɚ���7�ok7w�@;�ɕ�c&�����A1Ui%�c�T��8f+����u��/�m���97�٥�ӪE���p�`�:�bJ&.Q���0uE9��V�7AY었��k�U�v�wu��AQ�1LS~B5�{tn�]�K$��2U���f�l8U{|����[�g�ə�A���u�2L@
�˓�OPS^n��*e�d�[�rև3��zu�\�r{ 7�]���{���w^��1v�.�D�'��۱1,)F�5T��D���Q֋�9o��)��|����{��u|(-�]}��i-�m���t�xkL���m^?�Fjsr哣�y�@��»lʣΐ�X1<����)���iV۝F��M�E�F��0T�sjݙ��4�L(�]�X)|�^40�صp
�*�_
�����Q�D���t�Jj��-L������KDr��N���Ey�Nz�7�����J{�����v�����3�D���l#pVM���4p��+�᫰U�W1{��y�Lͥ|,lJ�����GqPC",�R�`�L@M�4�6�f__7K����Jr:h��ɺջ&-Q<}�YZTVH���:%�Z�[+9�$m��:�^��vT��Š%�S�ۆD���������Qc��<��\C�̥W&Ư���|uz�
oqJ}|U�v�g)��y��"`#C�2�݁�Ê� .r�Yl�NNoL�ٯ40�m����0�eYp�4�>�i�F���x��o�|/��}7*��&�:8X�o���%_�D��G�jw�/�ʍ�����؃�d� 0��.�W<�J����WE-��v��4Z�Ե���3G(�Օ��:Y5+��[E�]�A�6s)����yH�lu��1=���eY�I��o�)F�óx14����딦��t�,q�R�S�Ehs�]Ζy�l(������~�S�FJ=-�Eu^=��Nn�8�seIxl�n�b��f�R��=�]�'�~����m�&�4/m-�b���	���F=�Q�k8d�s����˩bǲ���۰Bל��w����[N�u��U�ݭ�j��A�F�H
"dc�L��S���hb�p�=F����u�)��9Ty��tEI��uē\��|�&���7z!pP�o@��;�Xf�taۀ�%�6��Zh�v��������v��(��!�+��{J��SQc��;9��SU7XYv�E�sKK�xF���k1�Ր�l���qw*n����Put�$�*au��ME�i^[�qJ��%�ML�������c�bg��|���gbL�v���ϸ��b�.��k�o���ʫ�+)wX�j�ۉ|O�e�d��hp�J�F�c��7Vͣ�^�|1�
�܃�ruy�7�]d���1cs���"%����fK�fʫ�o�N�����֢݅E$�G�VoÛ���F��P�����
����~@G���t�7�i�;ď�O%��iQ���\��yޫ�_[A�K�VS�Y)E��Vr��7������������=
Tܱ��J!lI�{�o�h�䅽���o�z�R�vѰ��Z*;�r�s����*���i2�%��Ԃ�7�\qt��f:����O{��d���t�+�*�ڨ�>Ѵ���I�p�ڗ��`N��l��WiHU��|:a޴��Cw��gn:�5�Ͼ���5UAD���$U5^�EQE3Q,KDE5RAU4E1��8�a�Q)K-USL4�Qf&E@E$EDEE%%̨��PL��B��"b�$�j���d9�$ATE%D�QEMU�j�)
JX������������"+3Zѩ���cX�DI���R�UY�4E6c�T�!�ʈ�J��2��(�Jb*��(�	�Q�EDk0�̪ �L�A�(�)�0� ���s1�1�02�aEPD��O+��<ʹЖ�=5of+�!� M@Xް:���ǡ�pאPݛQe�����"���G�n#0���JsB+�ћ}��gn�vBB�0v�P����^��#�,mkTt�������<-��It���0��dXhO��!UwFG��L|ꇫZ�>��[�N��7�QwlP�Y�I��ރ�c6�I
J�v��/�/X��UP����|G4���zR[޻b���*�9c:[%��gU�Q�
݇:e�	�*�ͭ*��|hM�Eh�F�G�I�7q�z2��@��$E����Uqԡ��tn���^9�E�TtM֩z�k���Y9�Y��l��[�]!t�}ڟ�G�C#�ZW(w�0�H��(v,<��y��7�7׹�nY�L����X.UiOK������k��W�_+��Y�^�6�ܽ4�9��7*�S`�䥇f2_� S�-l��:|�����/@Z�D�uq����M;NJT�_t�S��7x�v_c���!���$���{[�65^�[��.���&�\��}��Ι1R�**��ȥ�COEbV�����CH;�Rb����b���dư��hs���g�p�`ydE^V��A�R���r�.��� �c;#��}�f�#�W|F�W��m�lN�u��#��v$*�w\��r]�f&��'_g�B˲�3{f;��i�-T`G5��f�+E�z+�C�_nT�r�U=�p+ݾ�C[��/7w�Q�l�>��x?����a�����د�u�qi|�	��)�D�;E��_�n]��JV�I�ʣ"�D�_�@�j�`�^�Q��PM>��㧟kwldD�!��%]:*��o�VVL	5�D����|9VE��/v׉9ے�2��; x���{��������O-�O�Y摒��:�7P�,R�X.�Z���Ӭ��ty	�NK�trO-I�W7�f �?r5�@Ȃ�r��II��gI����'�,����8�����0��=V��I�#�����k��asZ��Ny*�&T�I�v�SW��T#=j��v'�����DU�-м�PgQ2��	*�e�5��Մ��h�v{�0��Ù{����ҫm;k��֑�X`=K �P�P�@M��+��j��S�K��w-�5�uJ�h#�<�T��E��\�0�B�X�-��,w�Äe�*����X��%*����2����ۭ��{�ۏ��W��ʄ�1L��F�g?`}�{Z�J��*YN���,�����y[箨�3v�z�3�"��9���j����Z�����BQB�8�Q�sz���3��+�9r��M�����9W��v�����Jr\O}��s�j�'��͢�n6z֚$��)ӫ3̽��W�*Vy�[���פ�iW����<OZ���c��ޮ���i�	����e%wt��E��3}R!��t��oRt���;��Vk��i���@� e�>+���6h��/�J�'�u����,EҘi���<� T!Jrb�J1�;	�I���ӳ�v�CգP�c��N�ol���C}J^0����d+.\�в��R�U��bW�� )�"�8�o��E�����ߴ���F�s6��7�|ЫQ�:s5�k0���0�}�������H�¾�4!�n]A]q�p9;�Ȅ^e���Z�ha�wݹ�P1�{�/W;�M^��>0J �~�O&�|2��.��؅uT6B)L>�}�7��U���5t+O��wƊ��Xk��V���<���̀k�l/��fo^m�E���!���l�C95���q������lя%�r��%A~�M��Ր����f��6{�Vrvb� C�$����q'r*�����.s�'��ʋK���zr_^%��]�t�BUIl�kC�:�	�Ĳ����_f�t/�k���J�EZ�)����
�Wdv:.͈n�{]sDֲ��4�$u.[�ޕ0�K�]]m�D�P������y��rGt������f#/��l�*����J=�M��S���m�6����O-1~�/M�5���ТY"�94_du��F�:���y/_1*�}-W�$���x�������՜��;j�]��Z�)
`�bo� !y�z��l�SW4�Ko,�3}�D�B��\O�,�8����Yc����`"c%�U�k���b%\�Թ��x��P�dd�J{�ڭ$�>�f���5�ރ.��*dK�z�5t:��e	8d`�p����N�_�ܧ�EQ�[��^�/>̗Y���"=-Ozr|�5õ��Y����5Q%7P�N>�5�1h�.mR�Sur��w���u��_eV6Q�����sv��{����DX3W�r���/�sث�2.��_ڣ�bNsS�&��=��=�|��:\P<9A~��خ��R��o�L	#am���i��t�J��g��j�u%œ���M��C�Ѓ�3q��94C�qD�"D�=55m+��M�g3�#E%�չ����U���[ʗ\����u{����#�k\���a���ɱH���ST�a�OnG��wӒp	y%֩{���PaJ��ɨ
����E[ðv,ӆ��y�>X�ct�/+{Yi�5�Έ9�w
���x?M�G��2�W�|E�A8�,�ٖyPhQ��>í�,������W�'��w��e���I�/���s}@�e��Q�����,��.lX�M�(��(���@��*u�z��Z߱��{�9K3[r��#�j�UϘG'���s�}J���t���I�FI��U�esڙ
�(˝ٹ��[3y�]�v�A�yCƒ����C�`r���7�])�֤櫼ik�ru������dL�	�C���b�����<���D/����4U�^;QWJd�8��w�ȎkR�T~=J�[G�����ʚ��+#�qgP��].�P3^�b@!��v
�U�����[x*G%gDM�X�ё�S1���k���1;<Ҳ�P�n�R�T���H���Gt�N͋�*uz���YO��(x�k�1�u���˽�ݴ}L��}�y���69�w��n�ZyY'|�i%�ҫ�AG�X�I��#4ھoft����Pҏ4�}���bi]����krVF��W��:�o1j���u���w�3E��^�K`�.á沗uY�t� �]j
�!r��DlWg��S�X�@�٠a�i,l�-�*�d�n��ت�ᢊ���볝���}�{��p��W8u��ZIly��g���d3f��1��-�q��m�H�صrό��]�2�hom�]+(\�|Ue�Z7���.�������Wl�ơ}�3x��\D�x�x"��碧�Ԯj�5���k�ްZ���qI���p<��΄�mU����ǯk���$�,c���LuW��'ޕ�
_C�@�#^<[��ޤ����P!7irý���61o��b]rKL0�w�+��f�������j�:l�1�F�,��ɩ}�*m���:�b:S
�9�ptq�Ħ(���W �d8\�Av���yCF��@��}"�k�����;+E��u7t��N��L�]��щ�r�x���s��@���#�`�b@	��V`��{�uxT���2S��'�V�6{����[n5����G�,�E�Y�kĜ��cS�a��R�иo{�65wQ��97�)�5��r�?j�R�A�#'���E�{��W�y���*7sݣ�ǳ&fzt�=���ޥ����%�)�A.�).T��)t�sm���e�J���XEjȫ�N�T�E]����@�E̘]P%�y����U��(�S��Gp��Ƈ���-[Jr#7��{E�tGz�̭.���Ċ�q�h��� ����������v�P�:�T���}���w5N�%��Y�v�tmD�%[\;�|��C���:��� �
�ӝa�J��ۙ6�ț�k�U���8���sz2&�|l٪rX�Fv�ėJ�<:a�0�\I�x�5��P�	*�l�_�h+E��ԪuYS�o�6L׸�WV뙻���W�������<oT�~v�ZFy<P��:��T$��l��(:<���S�73��Y;rH~o4`�ù>��lE[��4��YT��q�
��,cd�P�΃n�v.�$����3p�������!]®�l���p~��pF���u�:�a��{k^��{_T0ٛ6X��gn�O#D�c=�oP|��[�~�g^8K�	���
�R�{3&�Ps;[M"B% �ʪ���)���G::w��H�j����}WBJ�M��n"{�ى)��SQ���{s��������t�k�'�)>O��F�8N�SM�Ϯ�+1_}f��+c",1|jm��q|Шo�K�r��]W�{c�ȝ�ת�)�2����q�Ü�0V� W3�b�
W~�-�����T<ڂ�y5L#:�4�i���V��̷dʙ1��~�|�\�������ӳBw�/����,!�ָ�<!LIٵ��(�l��%��@a����Ṿ��+�������axo!��<2�(V�S6��{�Zuu�� A@$�[Ҷ�F.�1����V�i	�@Mto&�ٵo#7vy�r^��/9r�(t-�Ml/oo4��Sż�����!&
Qp��d�=L�MD�+"�g��}ˏ�޽�~��|�Gq]0)��p0ގ�|hةN!au��\�iI���\���1d��0�{j=���'A�n��1�㸘R�VY�1���F�mu�d��R8ɹVų/��#{����Zg��V�'7i����>q`�R�ה���(�5Ě܉�EEy��^Wg,�]�K�q��2·I'ê�ܑ�2oJ��-�*L��b�뱴^��X"�ɣ��� G�M��7w���Oz��!e��ȕ3����UŜ;[Ur�8���
#T`���0��|�YÅj��$���2�	#X���"~9(��^}^+,c��ޘX����M�N�w��[��f�ރ<k݋"��uڮ�]v�C4Պ*��L(11\kx8�zS%�yK��Ŋ38/ȞB�>�i�KᏝd��ݑ���t��0qd��ˉ���Z�ƹ�P9V�,Ɍq�v�X�[�T0�U3bn�nu����)�_�&t��U��n��z��ò+be�g�кa�c.��XX�j��
S�[z7�Cj4�f�E�k��7����u��2�����%��������l��/Wv���3��an��u@�2)�	D�F�\r�P��2�Mk�lq��Ӌn��u��&X�x����\pT��_�\O����=��uC"���4��Iwܕ ���G����K�#��^��8]W�;�P��ѱ\%(�r���7Ҥ��0n0���v)�j��G4����wӐ���G�b�:�$�G	�U�i����2�_wJ����B4{-�hΚf����ywI{��	RJ�|p�r����(1x�ĥ~f��p<�����"��sqe񄛳�����wy7.���l)ˌ:�ߖ�sSrv�M�%���1)_�:_��PA�eY��gx�Ȩ_8c�e���:�����S�ξ��7�t���& +�����82����Nz����a�V̭��}:�x,1�����&=L��걁y�8Gc�Y��/�5'����(}�+KX��9M��Ut�� y]�!Y���>'�^C
+S�6޾P��AE0���v9�������^���g�	N,���QǨLz�YX�k��s���!s��&�,�*�K� ���Ƌ�8V���sIrwWs�]�WS�wc	c1�2���<��-7V�)R��cռ7�Y���r����|�Vw[�4t<�U�9�]�i�]��<;2T��\���[�J���³_������Rd�w��_f���CӔ���X7���c���� ��57�gj�gWj�]ځQU�M��l�Ff��zx���U�yUC�*v�p���V�㙤i�l����� �Y���%�Pl�rX��ʇ\�X�^��i%��P���D�ҩ.o��l����aF4��W�
1��Uد]C�xMn�����1VA瘸������T��Béd��2�7@��"�R��� �yp4b
�G��j�Yુ�\�rv{��ů���F<w�)��j򴅐®��!W�t�94&c�"t^�����Q꼻'��VC�2�����ڟ���G=����$�,c�%TXw�-�E�,c�=�n��y׫j��G�:�4hL�⤱	#E�X>�,q�[�4ƹ%�P�Nf��%��Y7R�T�ݧ�)&�������1����R�����Ja��S���
�)�U�jNLd.��;�9�i>�xE]�O�P8vT�j�o�!���Ob�;'[7�Z_+�k�<�%�w|j���Ko�\ ~�*��BV�� "��.Xj�wË�����ڊ�x�F�#X�dS̷\���$R�D0�ǝ�v>5�cY:�i�zm^�Ђ΢�R"�;<�nBǌ���}���f�b������H�����ǅ%o�5�^�d����e"�bU�z����'��4{I�1�݆��.�\��=)[�P7G�g_<CY�Z�1Cv���N!{�	d�Z	�̺�sO���=7+�^�w��X+o?��f��,.[���w��}	P`@�'JM�74��S�#Gh��ĩ�Z����x4��&����4Q6���I��8'�0d�Kl��Z�s�����%e-�������K�5	�n����H�����N�ڑY�d�9�W���0ŵ�)+�(���"""��-�v�	�IYݤ�6e;��'oь�.�7`G��
�M����7��-�Ա�]����ء��<�E��M��"��U�e`�8�j�fc-���fÝ���d�u�n}Y�mr�]�M�q�*�d��Ȫs�&�-���1z�л��-ї�]K`�d��|m���쵱j���Z�!Ǉyڤ���{^ŏ��Nחy�p����@Xj�U+ʰ��u�EhJ�CoU,(hO3{9- I��N//�ʡN�K�w�-j�AL�����}ᕝێ����{���ʑÿ�-犡�B����=�2h��A�N��rdǊ��-xHN���.��9���OFj���-o�6�S r�NǛO�ͻ#)#KIzGD��:�1���^#����˖��q����ec�]��HRPR�%F�����9��z���.�Z��Px�]���_������mɕf�W{ ��b��򬦸jˡ.�=���Ꮣޣ�&�m)��gQ/@��V\�������>��GWJY�"4��vy���o;�;����GWsꂞ�#����˞� �v�wf\���><��Vy]��6Ӑ^$�+��p{z��gm�K��7�����q﷋7`Vfe`SW�j.�w���S/(.�y��Av�a���]�6�(b��E{|9�ar���ZJ��Ύ�En��t�)��᛻�K��ܫ�M]�����$y��PfNR����*�F̕ī6	h�Ƙ(�����q��rlݐ@}	��d��1�T\>�ً��)Q١%쇶��9&��|��X��#U�kJ7�N�$��J*鷜��S�K�wtkr�M��;V���¾��l�\�a�gJ�gxì�d�H�R�aocǒ=�w�w����8���z�1q�����x[��Y*�1[נ�e�c)渲�޳>3��Q,�PʡϪ��[����mB1J�����b����;���ҝ�v�;�������F��n�AL��?h�J��j46���c����-՘�q��p��Y��ΛT�V�޹��8�`�H�7�e�J��,���A�N�B��Ҥ�*ǹ���Q��n�u�_�/�����v�TESE>�=M�a�QTF��UFUPVY1���a4Tٖa�p��k0�ueD�U6a��M��LQQ�3����"�����#�0� ɜ���h�$�Z��X�+3����0Ƭ�̈,s$r�"0��#Q�METX�1e`UFXeA�Y�%Xj��'2�,�fk#,0Ȫ�Z��aM�d�FefaA�̃DD�FadYf`ņ8�YY�Hdd�Z2��ʥ��0�5��ʳ2����,,�'Ȧ �,,�,���2u���������a��9�SY�4fe�f9Z�D�s2�p,̪�3,©��h�N�,��"�$�P����s=� ��˵q���
�ayʟ�w�ƌ决��×�2�.6�|���v�\E�{|�u@q�n�Rףo�tǺ��=W�.�&�d���Y�E�dXh��������B��w��X�tX6�����V($���*���<�JH�f���"�
^=�`0����'9�����%N�h���Z���K *C��%�O"»�).T��)t��m�R�,t�R��M�[ĺ���ǩic2�
�E�i2WT	r������Y6Q��L3��ى2����N�+5x��z���:j��B=���D��p���\����>� �Yɞz �ڼ��NS����pIR�ҡTe��FM�x0х3.�P���4��'�-�_<�}�'[}��Wy�H��e�V�Գ�^ޗ0c�+�h��,cf�k�i�Kw�9��7�
YW-;���F4
������aǆ�y��]����j���g3.�7[�֘"��#�a���g���̼:9a���g�"oDR�T��2���YrH�ć*2�̸☙�#xW�H����
^'���CNv����Ӝ�\�V3f�_����V����j<�����ƻf��t3��6ow�J�!��`�/��b��I���;���� ��o��]�[�*�o~�x� �i��+>&]a�w�opX�r	N�Ǿ���o�<��u3�9�	I�l���-��x�k��Xم�td��*�) jy�.�ߥ�v��yN@�an�H�兩�IY50�Yf6��bB�$2�B�:��a�B��Rܣ�o7�>:�����v\�Iywlc*�p����0�7��K�TiM�k�T��ggx9���T��U�Hmjj� �YU��.#�b����ʙ1��~�|�\H�Cn�˨+�6yt�}�v$�������F4V
����Vݱ�Pjǥd��d�"j'��g��]�<|K������U(������ԏ"�a���Jq�5����)0�<��U5۹L($N��j�H^:�P=��d����R�V_Ƹ���0�ʣ,��<jBG+h&������8\���a����a�_�u]�I�:%�M�DḨ�#�lܭ�ݞ[f[/�><�6r�Ld�+.��b�N/Y�5����Y�$�z2�<��=T���V�V��I���hx�(w[Fo�T�A�Z,�<sj׆?��=5R�[�k[ʪ��;�˦������i��~�N�h�����>��I�k('x��R�얭p���AҥԢ�uon�b�r��7#N�ݮ��5�q�!�p��{�x9f�A`�ש}������-j3*���l>���G���B�Il���vV�E���+��tf����D�tl�>�$T1s��VNܳl6�+���Ղ_���M���v�q
*��l��2c&�ό�*D����d�y�Z�$�>�eLd��k˽H��ǵ$H��w��<��̘��)�"y�D�te��|�&������x�|zN��M�Xv��co��H�,<�ڰf�1���kE���+������&��N�z�ĭʵ��#4��ua\�-��>���-�s���|*P�6�g*��y�ȹl[��;�{��uO{i��6�3k�Orz�E8���Q��:�#�h�V���߫��S3�C+���8e��j��#w��}NT1=����(P��3q��9���|�������).�]��%���x̙�m�[%3~��,{�����A1�j���mk��5��BVj�3����oo�6Xc���pVq�V��O�%�̓X�M� �bb�{���ե9]v:��}����}`������-����]�����W��O��%.��IY$w��ao���M��;�O�C��}s�s ,�K	
/Ws�/�w�9������Y-�+kv���(Re^z�G�C�	�r�(�ܞ�F'�` ]���:�W��y�2	������D�W*B�$u9p�gU�L^8���W��Ԕpq��Gw�cbdQc�{ۉ�.$��v�r�����@�r�G�Հ<ɘw��� �+������O��Y�5���3�Y|ӓ3��]5~��Zc=Vq3��e�̨c��W�TU��v�B�e�x�ɍ<��X+���b��a����ʚ���#�Mg�~�~�+�X5"��Q�pz��k�2�=@�Z�܉���X��yJLW[Fo�T���+.�]�;VpPz��on	�t@������F���$*�uBV��O�ؽb�NyUL�YO����\(���N�M�8Y�i'>�������\s3:����畒\5ZI5�P���B�j{y��5�
��k��Z�)u�����c���cC"����I�n���*J~��Q� �zF{��
3��+�kK��y���u1����ƺ�/�CXf ��uV��֝��i@��MON8k�&�i��g!^V���®u������m����Wڸ*�[<:uv.S&��Fe�n���,	�p�>�$�,c���O�����������7��TR��^��'P͝#��8_��^ff����]���܃�� �qV�Y��2JZS���%�}�^�0���
A�f��%!,iW�F峴�R�&g.Í�yY�/��W�̂�K�ؤ�/8U��ys͵i[��AY��</k1���R�ǧI,L���s�bf�*O@�����,A�)�F��o�u�&5F8�ޱ��g������W�5C�冀c��C�ߕ0�.�FA�)�7+��8:�0�%�efY���}�uU�
%�8���|2(	��*h�W;0о�;+E�kWSp�K������Ws'*o-�V�͌�G?��q��
��l�}�Y���^�W�jgLk�!29+΂i��y��gp)���a�y�P�J��D�f��eh�`�9�:���q��ח�E���d���gk��Lw_X��?D�J!)#:&N�n�]/�¾R��nf���*��~&�}$��C�0��C�6kX��V["�4y�c@�����3�E�M���Qej0�g޿8�/2�,����k���2�m��M�nCGc�a�^^�哋���ɧ)��g��+0
����u��{��΢e1�Uv�%͠���/���)t��5�eҮ경�ꤖ���\K�Չ��}eێ�Q#�^(R|�X+#��ʺ ���*ex�̮7c6��#.���w�F2	Z�Z�v�v�o�K�K5��� .>y7u!����xk0J�CKL\�dur����#�'|�8�yW�7DuVӛP7U�U^g���[�X:H���s���H���Z�+:uӴ;/�0	<�B��_�Rvy�[b*öd��9�3}��õ
�8�5�Z�{gbQb}��PL�<C�U��(s�bNn�k�9=��ǆ�x �4����k;cY@�&2y�'��f�%x�fm͞3;2��,:Dݡ��pV�<O��y�{6�
.!�=��yI��L�Mҙ1y����G�H���R!��t���!����+��i���n[���P����1�2%�کsX�L�c.`pr�#W<�B.�ܴ��O�cQ�9��$����6�M�$)�Nr}���vk��!R�N�o��`�a�B���-VE#.��q���䨰r�aR�RQ�|K>��+���M�9.x%QY��vF��5Y���;�ۋ'.�c��/Ж��\���L�'
������/W�]Y���,]9�X�5�{��dd)~]�dB/y�i���C�hj+���TOaBj%��p��7(���	��gq�N������U���9�\7���**�gˬ5�Dғ�&!+�ƻ�;;�RF�r�S�P��f���<ȸ�f?.��-�|k��աVk�2m7�kz���1�ngYi����	n��RoED�{(�q1Z�ϳ����	QZ��*9��e+V��˃b����������.i��&H�Fz뷢
^���ލt�i�gca�>���������X9f����0����o��̪�kx�\y0W�Ί���]5H����nz1*��ٕMa�g�Wm�`��@��{�8NO9 ּ����ȧD�G���#���o�5;q-����L_���~����ZK"rjI�&Q1�.��B�9`h0Ii���^G:��"s�f�J�� �=96uV1��R������ө�)y�i�*R����A�*8R�%�;�$T1s��VN��0.F��4�m���(�*J&�K�Ld֣8��(ז<����j�ZI}�I�_p�t+O@�Q*�Lo'�K3hq��m�)�W6��/ȟcN����v}�A�y�bo}4H-ԢrO�0g�.%v�Q6���5��r����s������\�:HZ�/}��o]����+�6&x���T�g�X;��8��`�sث�2*}j��ۚ�Og�lm{{���c��s�����]x��%�ѱ\"�w((�U7ҧao��(優��{��jU�]x糯�(��
m�^�:�>�U�nt�	B���#^V/>��*y�O1�ma�ِ7����1s�O�[�n����w:h�d�c���U�7��=K��ˀ<o��ZE���r$/`�3�_c�	hΧ��eM<���N<ǔ\"�7�)x����f��~�� T �&�Vŧ�Ҙ��}ݜཛྷ����ufCFQ��ɩ�ReŴ�7#O&o��11�{�ҋG��=�)��UlJ��J(�>���0n��o�~����P�ǫ9e�;%�͚�ZlH(*"٘��Np�L�yZc}�W��yA+2�ӵ1o�/�<���~'`y��w�Se;�0��U��Ir��V��"���;�~�'Y����ͯ �8ѿd�^�& `eĘL:ftuiʴ�F��O[�5W'Q�e�f�*eh��t�`k�C���U8����t��퉘���s���u�wR�N;y1/�)z%b���V+[FHQ�eMNF��hb���0=�U�U%�J3Vң�������P��O�]b�yJK�#7�~`������gz��(�gw>��z�qyNv���)�NN�30s"�ș|���TJ���bͬ3d�\���[y�����K�<XsJ�19e:�O-�D��u�%���b ��uݝz�.����wN҂�H�1n�K��w�[�q�7C��"K{&^�J�V*>(�s�u�ȼ��$�[@zUp�3�ӡ�Oj �Fͧ]
�/�Չ��E��ʒ���mE&჉"��m0z;�`m6�!�3gb�H�Q��+��g��r2N�ʍ�!�p|�E��W�����<9_>��η��m��Aq`�t��0�o7*e��MFgΡW��؂��<�,�X�-�W�.e�\���+�b��\C�y7�]-�=u��F]x������[�
�T͸#3�h���n��T�
�q3��Hߕ����M<T�6q�S4��b�uLt��V1��ٗw����<�6��K ����C�@N��C^�Mr���1Ǳo��K�I?�F8�o6qY��ء���o9,��[�@�s���ʚ�b���E o���L_��9��@K���R�F���ֵ{��S��:��Y�F}�_i��V{��\/s�`��\a�Z.�u426>�n�]�o�u��@$5�u��I_|�a5�ƃ��P����\�-^��qs#�.e�<�*�<k���d�˄�n*�R�c%a �O��>
4�!�\,Jq@-CI����v�䬬���u��xu^�<I֦m��T�臔�j+�Ƒ�����U���^��_!�R�<`Q{j[=��yb�}�f�V��<b�U�W�����m]��i:Q��T"px�_Bn��j���a���r�j��CV���Q��,R�G�����2�pJ�2k���)��
�a��̃9�f��ߚw�9�a㹣�+1j���-tjJ���
~W>�'cǜ����-����OIU�@²�}MOIuή;zH��>���6�Y���;ɖ|{ޮJ���bs+�	s�}C.&��LY�7�Թ���v��k
�&�@V��X�
���9����D���U}�.e[��f���bL3��Z�V+�X�F�.VHH�'g�\*��]�ɿpx0х3.��q(�;���Ŧ��J�>�f���I�6s�
���T��5KaXw�.��.p�.`��E�Mn��d���5uJ�{D8��h�K��s�bLM֍{�n��ǆ�x9^K�0��;3c���"�[�&��rY�68������|�2m��Ε9;0�L#�^�V���皪'��jO3E瞩��:�8Mz�"X�2&6��w�����؅/ۍ�u�x��X�Yu�d�����T�z��G,f�W�Z�=�1��FK�LmC�}N���ꏋ�OM��{�5̜}\��ަ�A<�P�)ɋ�Ҍk�m��!�`�����2�7�����1(bb��I��S����r�c�g2�WZF-E�M����:ʎ5���fk3�F�L�����z�|	�duYV����p��Ɍ5�J�5�����%���F(���xu'�(��sC����^7{+����6�Yo�9@��O���\�r��ﴤ.�P3��tk�9�R�F ]���uܖ��>�у�r�Q#�)	Ie�Wz�9Ŏ��5���#Z:�i������@�GEKz�8���y�ǗI����u����q��Yrf�D}��x��7xR��{c�[@�vr1�Zf>ndސ���HdZ�U�M����w��E�kS^N��{�}Y�UU	��#�#����8-n+	&�K��K���F�����p�r�>���\rh���r���p�/��,�.=ؼs���i�o������|��gN�'x{��H�4��s�FEA'J��������v���P�Aq֜���F�խ�Gq������U��R�;��Ed�Y�u�ԑ���mA��\u�]7W����{Ms��kt�ȫ�5��eE})q�٬������%��v�C��t����"gbV2�㬁�})���1蝅��v�;��:E���<�[���Zqp����õ@I�<Gqow|蚆pof$��#�!g�L�V.9�uV�I��'S��)
s^4W,UۋtJM�p#.��b��퀻]0`�yD����;4�1fgG��c{���V�k|�(�KpٞV;��$OP:(卉_,�5הuG�h�'�-pT}����������h���7�;K����T��S���.�ʼY�(�w1L;��O�����"����X�����s�٩��t��R%������ê�G�8�*ӄ�E��iu�2���֔�GV�ם�Gl��h�JZ��;�V��Z&�f�m��;��Ls�ʕ�U��ch[K8fĺL���EY�l��;7]�����0e&!�YWJH�e�Zº/Oz\}R7yn�ۮܛ�
E��t�	ZX����Í嚺oE�Gw���Co���%[8�����3�I�coR��F�t�7�E��!s��ʵw������M���n!͎c7��;W6n<�.鸠��
��d���	��3&!�հ���O��1�3�P4*�ꔹ������o�1�&�f�ҩNRL�8��ӎ��%��k�.e��|��Ip��I��lB���U��j3Tee��~�s7�x�;��q��p�4�,��W�<[uѶ�^�o�gS[��n�	3{|�X%��T��,�J��}�gM��wy���]b��S�r����s�`Y�҈;m���;�d��ƪ������	"ѭl���:��Z�(bn�{��b5H�1�q�I��k$��ҬJ�N���p�z֫�m��y�C�ty-
�a�(���9.w��=�<��T����j�܏�Y����h�da٘fVT�䙙�QEY�����-f8�`Ff4�`ff�`fffdTƧ#YX�c�Y6FYQ�Ve�bRYeZ��Q�H�aXeae�f�aMj,3+2�+,3�p�#"�0rh230���̊���2+���	ʂ����NYcd�Mk2���,̢*3Ztk�Y�4��IF�+��*��f�9Y�TE-L��Y9�eX�fTLQ�9e�#VYY�����TE�UUFf4�"mY9���
H�a���1�0�������)��(�'"̳22���ȥ�V1��c�3(�30̣0�3
�	�
�0�*��ɪ�e�"̰�,�K2�"��3��*�5Z�h�k����(�*1̲ʌ�ըі99��V�ÄSZ���U�cS1Y��rY�T5�T�f�5XQ�FX�1�e9���6ff��f1�� �'U��)˼6��/Y��z�����䣔O�����j�m�{vvV���Y���x�C!��Z��'z�X&�-����э͖���>�pvB\�*�3Q��i����|�z���)gv��h7����rUU�d���\�<ڃM���h[�w�!�,+�D�+���q��
���v��w��(��p
������S�H��s˸����W�D/���
HmI-���j=��}Tq�A��A�F���sȻ
���GJq]qAl��u���Lu�5�M*�rlP)�l�Ʊv+/��d���b)^+/�\cL��B�ͧ;x����mdV�%�f�$r!r�q����ve_��"ǂ_]�I��(��$���v�Qk1jLɺ�(*����j7��0����
T�X2u���[2�5-{��G��,��;���6{s��g���Wo&�d��1(����T�Y����긳@�C�ܲ5�����*^��u��8"�ADT!L	��΍�9��D�5>�VNܳ:7FX9���ӈަ�A^fE�:�u�]*n1�Q��3hI���w�)���Kۨ�a�dc�)y^Z�vN�d7F�"������sYw���HF�����}u1%�j~Ix)����F��t�F��.��ꃰc/eGh���|qd8��/d<i��q�M�1`�%�(��d�+\����}>�ϭ��6_T�k�zo9G�O��-�ѩ���{�*]}�D������4=ST<���}r����6;���u�6�0�8�hR����BsЍ/w�fV�����^��2��c�������y��<��s��Y��R��i���m��;��8ˎ�u��
�pv�Dޗ΅r�,�Ǔ���{��\6�Ę��Y����Պ0����F��J;-�O�v��r$9F��9�D�)�A�)((�d��zT6ŭ��y=���͢�L���l�}J[�=�́���@
J8M�U�i�t�*�B��7·�5���궼����]�u��V��>8c,cH�p�Q{���1^y�Ɣ}���
��>�f��V�v��'%�Щ��v�7��P��9{{%��YU�@��5Ulh[pΙ����d�����X7�\�@ٛt�ӫ_�Y]�f}BW}u5P�C
��5������X+JR�VI��&J�U��}��ٵ��8Ѽ���FN ���{��Xۆ�/*%֞��UX�@YS,� ϒ�1@k�C���Ut�� y��Gz�]�V˃ݑS8��:s��N׎���j�pޓ��q�m�sE6`Y\����������h���(�(\��R�`�,�Q�_n�w Į�G�}��ݖ�X�+S�#����@��T���n���̮9�n/�p��ݷ'u�WS��U�ެI.��x��.��O�bbZ���\�e%�HÉ
8��51y��3i�겾�C�I�x;�Il�~�Oj�Tse�P���펼�=jR��h��J���3�A�ų�}�Sm�Z`�(��8�^bv|&���|�����U��Kb����*�+� ���x7�oY����q�7.��
|t�E�#�V��:,�\}��LV6Q9%#��3�C�7��{k[�G�_�<�Z堮@U��EV4zn��@�������x�8�鬝;.��(㕄aS��q
��~��(Ow2��|j���xP�Q�D�J�r�^�'aus����F��5�.z�;ɷ����yZBȋ�����'n>���#}FBX�����NGm��@Q�fe�wB�^�7�ufg��=���:��}�7��"�T:������>��\>�V���&2,r5�J���4Q���)^��+D��\I���U��\������J%�����k����FT�36�@��f:S�m���D���{"�{���J���_-`eZ�&d֝���M�@[nΠ���C�W�� �䐝�2z�]X�0s�<Mat#��n�����6i�a$���0��+���[��w3��B>t���AQ�د)���mG�В��-1ˌ�����YϏ.���j�ج��G`ʅ�(�;z�tj�;Tʳ�7R.{�{��X;�T��ׇ<L��=��J�t��0r��v��2I���hE6��U��D�\njZ�j�U��H���wqğ3U�d�#�r�Lo�,;��qx�D���(�/�&H��b0��Ɓ��g
4�{�ԝ�ŀ�M�����z�:�!`���C=�r�QU�7�<��i/ɓ��B(����-�핗ֻ���eXqP/�NM�EE���m����Ĕ� ��Yl�(�ުxꗸ�ٽt{q������������X���<7���c:�T�T&�XF���}�HO��<篭��euz1'%�^P�!�;�#��C�X5hs��&3��]P��_?�]뫅I7s/���p>@z��F�]������+I`�=\��^��h�9n:��oq���i1n����6'�~tPO� Wo��2���	�Q�^+ό����>K/*���6A���g[���p����z"���-����o�9����1'7Z5���S��8�)�L�t�=�H{W4���FQ�6�Z��6�_M��ˀ<�#��Q�.�	�S�N�F%��f�sE��w����ȳ����2�o���EW+�}a��WW2�s�Kbѷ��T�]iyۖJ���~��w2�	�g�Lw'W�دr�2��K1jZ�E;�9k ��{=w�+g���b���乹|��\��ݝ;�6z��e#̚Z��ەei�'��svE*ʮ�̵{Nd�LL׸F��$y7fj�2���%�|V�m����f��u�!"�{��=���_-k��X��/�=*�ڇ���vw�X��LOs۰"�v��/���a�f�5%�)h����Δcn��2(V�E��&jwl8#;u�f�T���6V���pp�S��*�3���� �S9)ˍ0VP�U{+�Z����0_��k8d�:ڒb�/���aD<ڃM����81�L�Q�p���_w����T��/��ry��n�MЪ<�W7��̄^=ZE1�.��CQ_�d��d��/6��	��'�;n]:H_"`���,PV{�����9Ցw��wƍԧkG ��/*0�Hӧ�y<|��s�}"`�j����O*�l�k�bp�q%K@ȗ6x7z�g'�yޝ˫�4�-���[L��g�N�������<���L:%1�u�>�]�Lx��v��n�Q�b]泜Cv(g^吜.��A�o(�054�(^id�>u������4PY��@!ì����0ؙ/����K�Yq���a�iwt���MJdi?3�˷|nq�=z*ӽ�l瓟X���i-������_]�Ǜ�>�\Ty<xI�Xt���s�&����
T�Y��5�<���W^��yC�jt@���yS�4����8G�'q'��\2<Q:�3|�r�����g?E����Z�mUM]��;b0:�/����+�?�Ad),	��΍�9�h�P�χS��4bd�.������T��+�g$d��xޏ&���!~S�(r}~��(w���v,�0�@��/ñ�Nl���Ť!´Q��Ɇ�g�����V���}�k��;N�_�βtq��F g�׶���ͪQg�ts�s�Mz�������'��n}�p5��Z;��C�!�a�����U�N�����N�u8�J�x�^-�|�.9�Ct�/���e�i�}���)]�%��	P�+������:�'���b.~0���f�fR;Etr-�
&����ހ̸닓��)�m7[d>*Z�t�36�h�yNf�c��J���)__v^6������)驨����L���:c�7e/���a�P']�� �^��6�n�j�}Y�+[2����K��IܥnP;��Jp0Z�L��Y%u<�ܢ+9U��X}��Ex�@��|f�YL:q�N���Q�R�#2.�u���</����}���R�{W�k�*"�J.Պ�}V	��G�M���W�/fV�������v�#9C{��Y}��b�hɛ�����!���;�=�:��Dm���ծj�axͿ;?F �d�Ҵ=�rDdȬ�2������E;�݌ʙw��%d�2L�z������ͯ4O�U�,1���K���1iG�&�[N���b��T7Q�E��d�H#���`mO-yة3;��uW%YV�oOM����ĩфx��%��Į%���R�Z�0�B�?����I}�!o<szt�N�:iۺ��c��,�Xf,�G�P)P�5�Ʉ�l���XUЗԻ��s�J�Xηy�h���>��Y���e����d���V��7���%^��%�6/X���S-�~�Ȏ��;^�x@o%�`�v�X��5��t�������w�F|Z�'Xɽ׸���kve�{��q*�My��@R��YN�����Vh�mt��W5-�5k.����k��U�g�X�����-��g�T�(��"�Ί.bxW�p2U3�:�#�v�3q>�o�pҭ~�y
DE�uY�އ�����o��m���lJ��\0�7qPY��ȩ�[�W/��/�Դ$y�ٖƷ{�-�I���-ۆ���x�\�}��1M��|j�ήj��)srb�����uN<�i�˯K�카U����ԩ1�˞�>w�p��ѳ�򴅑'�.�S����|&�;�@���h�����`��f�EL�:��@����)#~Tn^�u9R�1����Q�������.���ݞ�ҭ�f	m�/|�D��9	���I�#E�J]B����#���h]�ݽ�mY6��:���<�;!٭`�r�]SX�Tբ�85	҆���s�����Z|/ү�˖y�U�v`�+���q��8Y�,����U��pk���k�m�*g��`{����䮟��P��͈��W0�%/ђH�t4�f�|1Vv׃D���Y��Yݸj�̤r^x΁/e�b��Y��Z}����.���b%D�
&K�d�,�"⬋��Re��f�T�������1�
�C������O�|��QX1�d���޷�w��ǝ;��o&�'tR�F�)ќz}V��Ş4s핉m��֘��� �[�����eyH��:��rn������H���{��_#]e�b�\�߉���MU��J��qu@�0���,�њ{�bm��Ҫ�@��4�+`��ig��&w��M�D�5�^W�*��g:j]�&����"��J�-��H���V%p�	���t<��=:���{h��G��e�U�&sY��D�=��6+��e����}�㾖�Kz;�ߣȐ{Vb���[[f՚�{�u���F�5�EO\���X�(�\̠���$�� <�<����yf^�k��� {��ʌ!��F���T�Ia����z�T�<t�Y�lw�l9`�X�����|��>�=Cz�1�	56?�k�S.�-ȫٕ���sրk �����i�����B�&��~��1p�@�ur��`3�N��17Z5���SyڬPn�fofP
���L��L�l��'Q�d�3f�tL��iϹa�=&ݶ�*�=��h�s"��LEZ�v�z�̾��C��ơ�1�]˼9�3T�q]nU�H�Uu�Î��{�c`ޤ�{��Q���Oׁܼ���zT!1�w�羙ì��Cse�q������p�Ҽ�t�.5����+����\h�;�#8j�i��l���GٙyϘ��d#��3�¡>�/<®C9��
˗ �S9)ˍ0V��&�����ġ��qȄf�vhb���n��f�!�c&7�~�Ez
&D��1T�@�ܲ7�W?������QGG9��Э{����ո��h-,&j\�M����������G\w��)�ތo��2C�ūftYꟺ��e>�<�Դf<�H�_U�2Wb0�^nd��՚���]��[}״�<ys4 }��غq8�^���-'���+�4/��L;"��.�X!����-l�i�<��I��W�+>�c�ͧ([7�k%��z=�K�+`PV{.�>��>':�.�T>t��F�S�(�`=�������WF�	�/b`�+�l٬P��D���15*��Ap��Q�܏�o.���wPM��e�U6Ԣl�	dܫ��W<YN,.�r�������K�]��K#u.��Oo*�TW�bs�&���� ��6�0xaU��Q7ep�yn�E���
���dl7I��A�_@os�E����(x�+�:�3|T�Y��r@m��⣻��\�VY�ucas�MJ��k���)�A1_;8��ta����,�Bb�7�y6Sã����r�V^8cޘluP�d��\Q�ο]X�����_�;X�;�4u�$���dh�`j!Vw��Q���C�59�D��c�N�_��L۽�*���)�ђ��e�6�;��u������X���GD�a��!�z=�G�=�AW��W�h* �����ED��* ������ED����+�b* ��TA_�"�
�ED�W�ED��* ��Q���+��TA_�"�
�"* ��* ���PVI��T95@��M��@���y�d���[�
}�	(%TQG�ʡ-�B�J��k(���h�I T�5*A!���-b$mm��i%�o��Ŋ��CV�դ�Y�UJeTƵ,�m����
�-a�l�&��[J�bť�FJ�,�Se��V3եU�*�Z�-�KZ���g^�`;������0�����ۓ@M`�f2���(v���lʪl��� �z�ڨ՚�� -��Z(�]ݤP7p���Q��Z�ֲu��o ��&�ڀ	��v���:v��P�!C��Ӷ�Gĕ �*�Z�e.�Ҥ�Z��m�(< =��+�jRUl��^  =���    ޘ    ;  
  ���  /7��Zh�jT����R�[;6�k���[,  ���RؼˍEV�n�Wm.�ۻ��wuʹ�n�]et��W-Nڎ��J�l�9�]tNwjcb��ui���J�z�6kEPԚT�MM�(�fғ\�t���[��n����Z6�uN޺��6�ֶw4dsm�a� �x+Z�6��:���f�����!�f�U��ZjK�b��tSw7T4k
�t�f[meM��^  ��@Vi���� .��ՀvX
Yb���M�›e;a��.�u�SU�� o)U�,�p�s0�k'TɷwB��n�Nm@+j� �Q�M���mU� �=yw(jt��֝
� 6�M�ٴk 0U��Ԕ�"TT"`aR��   2   ���(�ꁓC@ ��� ����U*�` 	�� O�4JT�  � & ��E"b�4)�#SM5��� F@�I�T�=)�24Sz)�z�F�Ȟ��߷����ׅէ���Y���o��eY����/L���� @�0���ӨS���H?C�	) �$����@�����2I$� l�s�����������A��C�BX���HQ���!� �2T� !XN��U(��.�4��@U<�p����:��@��f�އ��'�i�V'�Á����H�??����sҙ�}o4h�L�i��eYQ���^(��迌u�{�ՋJ���6������"n�j{>ܛ,�6��Y[��6����R��#̲���GX*�W��v�4v�e�ít⼫������E;gT8�̱GNQ#~��,.[*�Ici�Dˉ�f5	yNM����x�ir��n^=�m@�[{{WZ�ld���w���JV�IK.���ݎ�%��5�tf�J�8*F6Vl�N�"w�&\�ҥŖr"Rp�����[Ŋ�sTܲ�IS)G�J)w�T8L2��5ia�U��u>�c�6��@)^J��Pg[h�D$\�,D����T�+$�# ���7*ԄnY8�\v0DL���SҢYId\x�%���[gZi�@�n��D��'�^�Bt��:���w0B1�(Z�^ط �5��,�۸��8��cw\�a�kl]ۼ�١I��ܦ�ړ0�!��r*ԵGX��"���ö����T��Z�3�J����9���M^`��OU%v@yI33)������rnm`lY�bĔI���M'���ח��%TIKZ��ݔ�d���bfi���Vs$�V�t�D�1��3&�2X/n�X����3J�/u�Λ"4S���,��:zt�*��DL����B��,���6J���Y�-���fT�b��;)�s���H�xKW*���,�m⧊�Xx�x�Yu`�׍��Z���y����rO��J�mjMr�`#2�/5Et
��%#2�b+r�l�I�yF��Y)� f����Z3r�3u �\�_g�RD�L�P�X,����\k��v��n櫂�D1fΓZ�e��ةA�`W�h
!b��ke��P�g	�2�QP�Ь�L@�Zw\l]i�T�惹����K\�X�w�XCW֕H���[��t� eJ�W/I�D���K�l�#�����J�,Ebܕ�P*^�f���]��0� �uc��Ҵ�""�̊�.n��Z�3��
��oN,�i�\@����P?n��K2Tـ�X�op���[RZ��3x���Z�w���7��m������0�h�c�,P����g6>9�,O2QG�[]^�<F<1�Zm��L�V�����.�Q�a���ѭ�e^ecה' x�	T�Dst�06*2�lb ��X�K�YZ�1�#j���skm��+NcF��xv�h�͖71>�l�72� �KՐ�
l��Դm�j^�v���R�|������	�H�r��c�Rn�ܭ�5��i�5��-Ɲ�X�M����ݧL�v�TD�m�1 6m˺y� GB��v�n�c+ӓ*R��XlV ��j$�BѣSu[9��Xy@DF޹Yzh��Ⱥܴ�D�{�b��Xh�x�B셌
�{I@�ұVe�yf�Ħ�e^�2CQ^���#Y��*�J�#$՛#;��v�Vi�-o�t7�C4�IO2-+_[�!d��v���J&��4nZӔ��~fTU���K�XV���B�S��U궎ᛃj�(���-�5�ܵ�j�'ie���{P���Yn�N���J���)�9�Yr�Ref$ƌ	�U��G%-̌a�q�"�sF�*������	fj9����包[�e$�+���kr�+�� Ѐ2=/e�$N��Qg�,��kfѴ�6.�j�l�9"�V�� �#V�DTܖ�h@sp���yd,����ŕ�>��//jYd��0,����\Qح&���nN�JFP5�B�Pd+4���r�����j�e^�z(2��{;���P� ����gN;4a��6��n��J����#�u�
w/wH�[��'z��wt�t e�4�V҆�MH�f�M�J㸐�f'b�ۥ�$��-Ck �[��3^�9!b�>�{6��+)�t�ݔ�E�eE���v��s�[!�sfCp��o�m��n��V@g"�*U옢5���:�7,�j��U��S���k�D�&��W��*��*Zu�6]�5��E��ꕙV�$w^�`���[+�Wg�)�*��9u��;�cԍ�6���WҤ�T��
���5�㡤���胕�ٺj��u�	��T����jTр�86Vژ�a:��Ϩ�Li�)3��h����`�XPU����-�ShIP cW���rT�E�x�L�%�&K6�Ɇ��ئuD���hr��)�us1�6��j�9W���b�+�YDaB�+�e���ncx���@ŕNP�Y52+ۻ̽Ј�o�#V<JV[%aѱ�h6��`����Xv��i@�;�*B4	J�T8�6���MFV����u�toh�n�W/�Rib���� %R�+�a
�n`�b5�Єݚ1�B�M�}�:ʟDNXZ��8�v����c8i����j��um�$.��q9X�D���rR��l���C+XHm!�L7{r�hU��X�
�ӌ^� ���f%&f%XP˽Y�T#��@n	�DK�ᛷʃ<.��]�Z���d�9Dk�[��ɻ5����ݰ� �[���D���C���F����V�ɘ�1-����K.����F��>(M帄{f��a�f7`^�k��PM�4"�S��1��{���lE�hڗ�a���0�F��q�4�ÁhS["�Ce�3V��t+%�b[`��a�[��Ah�h�--U��S5��Ok�V��2���*�Y��bs,$F�
e ѢH�@ɘ�9Hh��Gө�X;m͈j���S�ֳ��0�i��}��
v�i׍ݕaä�#,�
j�d��hґ��F+Fɣh�Ѫ8�,
��E�%��Ι�f5�ݨ/6QJ�CAT��hU��l
`[ƥ@a÷0ޢ����87i��J\�H�X�h�n���Kf�H`��4u`�&�,��b��HУ��a5�s&�Pd��˿�hB��<�V=�|���#1Mm���SB�P�kSh�Q��9v��&�!�ږ��2ݝ�쁬PT�$�r��wV��v����xP2[M�E4c��P�=��I�q�։W�u��SP�s%�tP�����z6ջ(�еT�� �q7D�d	˕�DJV��=8�S1������Se˺87	�ɵ�F����8�.�Y�[���輨�_6���/RtU����@;36L*�����̅%������Tb�f�N5��nm�N��z�8(�S&}��tB�G!͵3CS-�ƕ~�n�@��G lZߞ�ю\�4YÁAsA$
��ܬ�%���%a�{l���M�T����lʛm��v��#Z�CF�+aͨ*D����سIݸ�yvU%��8��{��L��zr5xoe�F�H&���	���ډ�n�W��� .��)֘�Rt�,�j�޲ۺ�4���[v(�W�ӎ�	�7�c�)���y&���Flو?��&�+U��qpN�{\�W]��_,%^��]�
�9k�X�9w��Q�"��A�RCXӱ5�̻�T�q���ZR�Ѹ¬tb�2�f��YK�'.��^IMf|�ZԮ����ܓ"�Q+8U��b����YEJ�+1ԡFµ������J��t�!�EYK�w�����4��z�P�m�R`���O,#�&���b��S剻�Y FPHar�$.�k3(2Pv^�kjj۸��P�k	�`J�{r��Y��z�RPjք.�ZX*�X &�a{d�R`�n�+*ʭ7Al*fj��X�sQ�6ALD��p�
0^��ټsU  �|��Gf<J�Q�2�����CY:����I����a�R���%I�ɣN4���oj������X�Lvdwi��"��*��@� ���F��2�P%�����M.]��x��ud�Ǥf���GcI���b���Ǧ&5R���>@��l��6Ѳ)�x]H�*�	@��� ���J�P����m��$���걀�`�P�[��\������n�;�M�k`�1�6��YX�JkfL�( �ZU@ �ł�d%[)K�V��Df���\�W��X�R��h;P�w�BL�.̺�&�����1��nQyX(�mE0�6�I�s������_W����~�����3�ovh�	����������'v��-4W�*u�W�_����E&��]��1�Ӑ�.�E�ޑJ��jN��9e��>��$�������54�+:J�nkup袋-�1iX���I�Gwr��(��]e���e!p9�S0:\͒FR�ʻW.y�f/�{��1t�����I������dMp#�P����a���n�y�xh*�F�Wa�L�p�Ҹ_m�x�zP<e���c7�	`����@�|�Or�r1����e�xFR��oqh8�O�7$��_>�1������;L�u�x��GWe��-���_`v�ԡ���k*�wt��W��v�C�ե��Dl�Geɢ��y%c6hw��s$��0�ZE�<�
�ڦ��nW���_YB:��H.-�w��o\����ɜ�f�b%N��ձ]��w��\�Y@��+��,�0��"��33����ř�l�5|q�譹�O�p�´:t��w.U�*ewl��1l������[�������d�A�S-�G��-�%n��N���f�9�����L��5YR�$��on�6h�w��ҕh0]�bv99��ޔ����u�OP(M��~�Z越�)נ���Ԭj��ỏ\�=}&V��fBM�V���+!oL�����f��Y����%Ϡt�G6-�Ky�xz�wm�q�G_K9d�F't6�v2�U�׽��R8���Z<�Fwlj���9�8�;���dT�c8��k�,�e��U�-9"�4._q�!�3f�}o���K{s%�v:�S� ��t���VB�^�C\y-t�{B�A[�Rw�8>&����IZ��JWS�m;pŋS��Kڂ֮]k��+��R�-�W��NHk}�rj��)��R�Z���Y{1���.`�&��\������kpV�>h��zNɏ����ʐ�(%�$��C�8N�n4V�/{�ta�`�]HfֵW�T��:��&|xӫ�LI���K/p}y>��q¬[8�v��\{k\z0�VIaFT�p� ��&_�hŢ��w�"D���ٶ���u�i������sX�H��)���]b+K
�K��D�[�Z�bw�T������.�u՜5 }�fZ��W��������#�v����$�)���޼�/����Y;0mE��qi��>�D��Mo�Z�^�M@��㢭M�$��L���,��M��%��W�u��]�B�!e��?u>8s0�J��%��h�ڻiE	uٔw(�7�����q�����S�P�{�|���um,鹑p3�g j��#�w:�F]a���8.Gz�L���%'Y۴��eVhp2Q��#��)Yyv$]x;h�H��uM��$k,�v�
�&}����v��U���126x�OD�)�v,B��N�k(�R�����e�F���>�v����؏���Xq�C�����������W�Y����%q�(��}:ve"��kC��]��n��&	�*�K2;�<�a�pX�Ǹ]X�n`�RuF,%�`���4CS\�ˤ*κ���"#b�o^^!cT2f�ѧ�﮴��NSf__�vk&4@A�ms�rȒ�w/�ڃ��NFx7��hXhb'�..��>ޏ�WC�Â��UI����;���wNK���d���N��r���wP�+#����V��W\�YXRP @o�t�Ƶ3Xl���<��� *1ɽ�t���wk,��)d���Wr���A����=u5����#�=�O���� �Dq��a������Y�]fdi8��8������^��Qa}���	Ts9F�P�dE���7d���[�ި�/p�:�.�.,V#�M*C#�%n�cy�T�� D�����f�U�B<%��U�豬Ԕeud�N
�aP��o!�6J�'XJђ�>Y�/��6��K"N��GA�F���9i�� M�䫉.��I��.�Ҩ&��8ň�AN��9���x�^�&�0ٵ�Ҝp$zB]����.��C��*p��W»`��H�E�̌�Mp�ϸeMڅ�]���݉���n����v*�v]�M�;Z�>���sv��P�.�
�:po�q�o.�d��!��v�	�x��Ǽ��[��9�����.2���$�帮>���XNC���s���9��re�ȒUl3S0k$�
����H�;xR�Y:I��5����va�nw%�s_�بZ��w�im�&��8���l��A�7��Ө���CL�a*3
9,�A��XLpo�dY��=��_�&q��헔ZH���I�\��6�&1��^�⯹
�����f�,�����*�rJk�Ԡ����6��0�P�����(\v �T��6v�T��V���������/��F�pܑ�2��D�+�*W!��K�}oW,<G`kW<B+��E�޾h�n�s�JD��\Mپ��}���V0�nd��2f2ˌK<�ќ�æ�$�FhԆ;3n��z���h1-2�o�m69�7O7|��(�`.9�Kw2�s-�ַ��]D�]n�(|���=�Zz�^�R\ʾ� eu,'.��^[V����b��b\}�]�]K�ܚ�{�s��CU
кD1��V��i^h���b1ՠp�`=�\{!�!kI�(���q��B�r	�2��&�p�8`���e�m���[�U���L{w�48Eٗ93"4�yI!S3orLY8��2Y�
S5�Y��ıIV���U�4���8K�dmvL�v���pK��C!6݆����º7��	/E��4j�8��
���1�}�e��(|cS��s��1��ì���+f�A}�G��d�ْmX�v�P�Ԙ�nBW-�zb},ݱu��os2�c����L��ώ�$��6�P���Z*Z�Ņw���J�d=\-�{l�9��0����Z��ZIx���uP�15��M.8�Eѹ��W�r'�^�WF�P��%ޔ��]cԦCS%Hze��Й4��IZ�\��T���8n��=�X7�s��g\��j�L���\Ć���7����p���l�Ɓ�*�(� _t3`y��B�T���u���(��NwW��ty��cʾ�É�n��:�Eٗ�!��cz4�x��y�0[�z'3s� ��bT�/F�0�.O��tyQx���D�vSP,�{\jjwov���"�Ւ����΍u�{pyR�e_`[Z&�tcp�]��3w����vC�/v4��N���4��9��WiZN�Gc�ᮣ�T��V�2ۢ�'1ȹ���g4��t&����éTOh�*��9��/���[�F�X��\�O,� �ʄv^fu�l�Ҳ�	�(��:�q�7b�-���`Y�U�\�+g-E���E��yz�4b�'l���{7x����Ưw��9�x_��o����H.�+`���V�Ky����v'P�e0v!��>J��gy�[��6AC7؀��E+��`3&�L�x5��oi1n�eYۨ�|���cI&5̣�,� yEW�씩��2�]\(�X�I`��gv��m��2���Ԫk4t��
�U�!y9L����4�t��Uˮ{p�v�C[��H�n�,yԴ��G1\H��F��ٝVj8�n��ZRNھ�[okl"%ҍ��
h���~��8(e���E
�0��	��)��o"/�g�N�;)B��O�990��.���h�fW[x���I
�:���M�D#���S��2�ű�A:Vȸ� ��ʲ�F�%_]�����!�#��o$�)$�������[rpPu�R��Vש2��I$�I$�F䒤�dr�Z_C�s��D}$�rI$�I$�I$�I�$�JI!P�!�)Ii���4�d]�Wԭ(��M�z[Cf,����L}��yQ�ؒ�0'�J�US��s#�����Y��&�1�GNv�vplM�bK�&�5�䜹1�%an�Y�#�l_16�*m�$�H㕋��}�V�Q���U�yyzJ.d��J ���2�{J
Av>A�v_(�d��s.��r�d��$RI$�I#��2�h�G�qr1[R��R�7s������rI"JN�)ZdqH�8�s����:H�H\1��8��iȤK��Lݏ������#�'$��$�G$�I$�I�H�rI$�T̝�+�"�V��}����k�kK�l0�0鷷3Mf�R�~���.�~_� I$�A:�}�D�	�~�'������`MI	$�?��+���C���'���tVp��{ڴ܆��U��BT�w�z�r���ŇK��u"k:��9��õ�`W�'ZR�p9��{x�i^��N�KR���S�x7s��-ٖ4��"8ظ{�_����VXK��fL�V�p*��S�U��Xrv��ݖ7&��0�(bR�Jq�x$�CUv.f�DLY��B�q�n�nc���=dS2�J��7ewf����lys���e&�[�
wj����6�L�Gr�4�\�m	�f��ɇn�"���1��v�0.w][�w܈J�K�H�h�Up�g�ƗU�%�5+�Vfd���t϶>q��ڄstV� cy\3�hd���Ld�a�j���U��iću&�l�P�à;T��le�˫ء��h(��;y��摍.��\#�Jv�ݷ$����fk�ʚbՓv��7���l�&�����+!���o�B��d��]�VF�,"�3�;�?m�<)��3�
\�̻��8K�Ǌ�^Ng�
ﳚE�
�$w�/��A4�+�����<��8bD>��#F^\�o-���#Ƕx4�����f�Pi��.G�t�ʱ��Mm�$�?K.��r`�ge�B	��������+*ݷ�v�G�ܜ��FωQ�\�:���*����S��+W���wx!�-[nh����\��k��Xi���|j=xF2p��j윉�],:&4>��k��97�k���=�3����
h��r�eG��2�>�+N�-�v�rO\�����WA7�J76��*,�����NFn�F�������jѬ��+��>�.�Y|�wJ�P�*t���oz��r��Jz�Y���U{P�D�e<�̩u6����́��"GI�dޕ��=�+�<l�(���`��b;��_1^�Ap7övU�C�\�FWO��b;y�,��So�4t1n��	[��h��;��7�T������}J��kz�X$���5�����G%�����	�(_,�Qi���\�bL�61
��=vK&�]�ǂ��&z���(�P�Y��b��X1ò'��v��8Zʹu$�x�2ݚH*��D;�7t��ĺT�-e��f��LQ8�K���� �ږ!�b��gu_����T�e'�өB������������"ΐ�f�����hn�u��Xض�]�|��Gj�dڗ�JtqJwH47c�֊x���m0)wU�b���U����_hqD�����W�[�Go�>��Ich��FTv�x)��HK���ӛ1ֆں�E�f��u����
]����c
�e������:��q:�YO��j�fV���nj���j��a(�@�W�(>��ݬ�E����˷��ԉ�3O�1��3�j
���A�KS�C��i]���{q�#�;j��=V�Řk��R,�*���.}l$��LY�8����^�3����b7��q�S��$yG.��c&J��V,b�\�-�an���HwK��P��j�7*^m�I42�K�9|s_Q�7`sAs7�3m��@1/@��Nylf�U����s��^�T���|p��������n�ś�z�I.0^�L�t!&N
�y�L�CyNG5���ݒ��}�
��ܤ�m��;V|y�g�am�z��J�K&I��c�h��.�\�0Y��J����ųDiQݒĨ:�β��s5�_�m�ꔉ�B8�V0@���7��"�S���k�J��c��6;��4qHy]��`����X8�8+�$B���.ǘ�<+�"��c0\��|�Ѷ��jΦ��Z���a^�/���0��`�ʎ�:\~�@���t*�v��2�0�jk�oQc�kw"������t%�E-s��ֳN�u�1&Uԡϰ�K���1������0�Öo_
@�<R,�n����>.�G�:u啜�d9GV�A�Ĵ8�r�6�]����EZ"���-��w)�ծ�}ا�M&��s�)p��5tܐ����8��LWV�L�v-�u�ٷHӃr�J@:f��]9�l1+A�F�Z����-�b�IuN���q¤��A�gRmI����l%�X��<	s�<��@���,����r";��_KlJ��	w[� ��}�N�	��t��H�Qщ�����|�[w�����{���V�̽�&� �(�EbkN�swn���E?�C�k��I:ZoS�Iګ���qd\���j��۽�@���f1��h.�|���$����t���M����{��A�5�M2QLԁ��?�)���ő`�F�_��6M�#�X���%i���	�4��{_\7O]���Y|D9g�w�Tf��C5�I$<��"��k� ��
��'�����	I�2�D7z�,�E�w�j�T�qq
W)S�5��%�f����'Vd:xU:׍��$��w��r�V�<�n�]!@�4�yF����ETh�m��n^"_m�L�����"p%N�! ��3�*�v���:��՚k!9�˵��r�g���.�0�[��s�i\`]رh��5�t8�Cu��(Ճ�&�B���HaT�.�Q5(���[/�E������A)d�\�oPr�9�j��@���Gv&�iguэ�����*���O�]#im�Y�T���K=Q�[��s��րY>]��wn��u]��dѩ]$.�"�RI}�F��nhձ
�"{i�V�-�_9�n�i���|���;�Y�C$�v��=��)j���.��["�*ڮ�6��-c�6ۺ�9��V�Ud֞����e���!S,�V̴��7c/O���*!9T��f�RRl+�DcO0pq.�sN˵�yti�үa=(�-]嚶�g4Xٺ�D1k�h4L����by˻��D��Q�N�x.S�|�o�����G\�]���Ɩl�z�3���E�(�#����缗k��]��ݜp������$+b�������"RN��U�m�
����m`}2#��`�����(fٷ��+�A��F�s�[Wf/�d%5��d�x̮,5��(�"��ӱ��q�쓒��h��̚�G�j�#�p��D���K��'4&q�:�aW��T�h��1<\���:�49V&l�}����4�����&�S+��ڷ&�E��:�I��E�5�|$����n��	+��ƻ��$�Tj���,T�X���"�q܉�]ٴIt�k�/����}.���L���i���洚�����r̽�|�n�VVFWt�%��+�X5� ���U�#�����Dnpv�q� ]��IM�y�'.82p	`9��R�t�ԷiWU�pʾ��4jJ��bX��bc{�G76X��	���6���u&��G�Y�N)�Vr�vM�Q�5��Q�G%�����F��n�Ρ��Hw �&3E�#M �X�squ0{#R���O�*$ݾr��ڸ�w�*�L�T��GnD�}}�r=[��>���v�d��\�v2�Yg��=82˓%��vs*�[�������Ң��+)����pqWw�W�^jqқ{��;�H��W*w�P]ɮS`��5���r����<�m�v����D]�_��^�̓G+Β���(
oU�u�ʍ�ƞ�N������EKMN�Sc�T�s��b�7"��B�R�f�	[�����k�Wd
��B���}�P�pQ(�U���Y�3%��i#an&HRՓ/!�3Bek���Q����=�!�->���wWA,���:���lA�
��*�,�2K��1�
3A�Y
�9��ύ��s3s�H��ֲP���r��(��x�C�'�u�r^EGe}յ���K�j�am��D�eI#�d|U�D�r\Hƶ�k����W�Y$�Jc������^�o;ZM`
2�j�����xU����Gd-��񑔫�t"`P�`���WW2�V��ҬJO4��.MÕ׬��Y��vL[ ����x������Yw�y����إ�N/���9�����&vU�S������1�N]�gk$�����n��|�	��7'5\�.�2�p-bݥ����O���N��Ղd�J�m<��ޭ��M�HZYG���Ģ��]LCtzV��^��R�e egX]�[�*���BVcR���Ҭ'k�vDޭ��lB��ƛx��q1�1|�W�:��λN��W?~ HE���� �~��J2)j_߇\6��0�R�[Z�1��u�U�}������}`�������wZhsӋ���*u���̉v-�f����j�xw;�x���F�;�A�,��U��c�y�k*_��V��F­�X��JX��F��_m�����<b���j�����-���.�+q�S;�uy���:�bJj��bɗsJ=���!�<vb��Y��x�JRkߘ��%�,mn��Z�(jg����.�+��#?��xjZ����KˡG8�'I?��}+���1�L�|kB�Y' ��wLvq� �k9�4Q���X�|��e1�K�b�8x��7pt�u�1�<%л��#H�7y�9&�65h
����:��p�C�dG��C��/mn��Hdr&�I��8"�P�PP�i���I�I$�	$�I$�I}33��EU�y�m�J<k"�$���%�T6����`0H.�R�	��PU"�E�5*T" MS0�mDY<jb=�Lq��*�T��5DdP*\N�*,�R�&j�Hb��++��SNe*e�%s/Y���L*���a��,�jkR���R�M����cAV0�fx�H����
Lj���X-�
���ô6��&��FDc:�@W,�+�C
�DG�UVE��]P��U{@�^Gmiו=r�#^P�s���{ހW���ׅ��	�l����oEe�BK� `�%��G���yØ}е ��Co0N�rG��P�b��v1���S1�6�L���[�f��魡w\�d�DcO4���-�|�Juc��*yeSRf�`,�:(�>+z0�bՉ����@� 3��Yef>a6�]����&�d[�{�k#z�{a�t�K��g �2���\v�u!�Y�`L����e�P���Xӯ�^�R\E-�w[�9��VlMlv�p��9״z�I����!z��b�����Lz�D��.�����`_^�����d�����^�vt�|�m��	]Ze�(�(�,��)�۫�Jo-`ʴ?�T����9ErIm�v���5���ņ�(��ѵsר���-ñ��0輊����!qD�_O�u�%%5"��Vo����*7*� ����x"��vOF� ���WuՁxg(p	�
�~FU��+����0)�d�ؗ6�؉if7�ٳ���k�7W(�P��P��D,V"r�Ե�lTl�*��k1�Y~�с��v��<�/Uv�n�;�=������^� �X9�N 
�"���OX�ؙ�^�O"�s[������-���Ca��RQU���V�/Gl�.`m�-+ڸ��XcnE��N��ժ]xdOLs�5��\Z�w���5��}Z���]r�|�l��{�x� K�9�t�W\}ڦW�+����oy���� �c^����t��R}�5�%��E F�{Y�urb��WǋZN�B��XUbW��m^�y���hgj<���q=p�9�nJ�*�ub����G=-�^'5�_M���Rn�y��Bo���J�W���e�CL�����3��܃O���*��vv򷶪����G��̍i��Gd�9Ҏ'���t�5��
�ΧԹ�\O��F8��u�< �䇕>�Ǿ#R���9�]i��5�A�`	��}y�+Hq,ˬ<��z�fs�IK���y�	bw_
b8n�{g�6ִ����1E��vv�*g'���pqP-߂
H�v3oD�k##Hj��]�u�i�gN`�pT*8 ���ֲ�l]��b�]=〆7q%&='��-;�V���5�q��]r&ӈ+N=�)�
/F,B��ۋ����E�M@#�iPYV��y��{�IĨ�Q�����n$����+!8ɍyh;��^��s��I�-�Ŕ�̖b{�=w�i,(���¢�F:dKcw����2��ä�dB̭��,IJ�>�`��3�Wf�Oho��4z���m�wX���i�x_�V�,�����9ujm�o
0|\�~߮���o��G���݁2mj����l��t�,�0�{���[��fI �ȴ�7�}�9+��T"�ŎS�V����%��|�����=�O]
��r/%���+��G��nT�bbٙeB��u����=ָ�NJ.9��J�
"�$�V�b�e�('\nl�x��慨���N�ň���ow�.�Wn6�&��V1�o@��Qo\h�����f>5��ȫ���z�?�>Wp`~;s��<��Z������n�;`oX�'6�Vk3����;l 3�.`g!37hiI�]�;���X�i�+��C";�w�
�+b����N������j�g��j��Ŵ����﹩!�K匋�g6n�}:�����T.�E�H:���S͎è4�'P�zE���-���v�T��!^(b��}ڡ��M!�0s&��T4�]�27�diۅ��܂�e�J��.�(�5�m�Z���^]��E��S}�Hz�7>]�U4��
���x!@Qn�;��uZ�:/b���t�V�F�*�:�:¾�sn6�%ʓ��QQ~$���Į�������f��rk4*��-7Ш�J	�o-�h&-�%~������UX5[X]x�m�Huf���&���=X�����^���`΁�xt+L������`s�`�kד&pͣ�l��Aa�*��0�S˰L�Z�;�j��=�J-`���Ħ�G��{�X�B���Kֻ
[�R����,f�l�rVnY��`�(#�W�V�o���_cL��'��ښ����l�q՗������h��n9�.|
h׏9��%p�{/<�7҅X���4��W��)Z��p��������X�V�}���-�q���@P�z/qe�+�l�w '��W����[���A��[W�+(���i{��R�i����/��Y�1+E[f�k
��h�RG;14����P{��QSe@��,Ɨb���+�M%�4�]hY�7B�@j������i���(� ��e4F�9�)�P�����CkI=�8h�t�y^�s�A��;i�K]ǣ��q��I���t���J�k�#���d�B;N���OW���2��j��2�-b�/6e^�);����w?.�a�؍����͢�u���W���E����eX^�EɅ�J��%���P�QBA��X1�וOgQ�Y�v��NFN��eR�K4=�j"����y$Yq�1�O{�K��1�̛E3ʝ��/�e��e��,��b���e�ù�x1��[�ܶ�b4:��.u��t�Zj�8ݨ|/��j�f�`m�Ms٪͈� ������0���q�JD:D����n$F^���Q��ա��b"!�!)me��޾B���5�$�[Q�)e�	�ӌv�x�q���9Z8>��fay[�#8�RN���
:�x:�'N0�0cVR�mȦ�)�z��@�Ǉo��gI�q������k1�F��C|��]��d�W�>�fc�z{��Z�K-8b�,\9��z���'VM��=�n������|���m"WlMMhB9��x�T����	���u+�	�7E�΁���'\�;�՚�eQ�q�<���] �S6�	�a�xKB\�&�'��R��)<5@f�\LB����W13�o2����v#k�&,]ŵ��p��u�Z�ʛu�J�tdI��ͼ��{�U�]��_[�[���B�^	��l�je�W[�����]�:�w1!�K �*@���r�g�^Tɟ3}kps��Ъ�3P$ŭ8���m:��Ҳ�c���:ł�t��լ�mQyq���ch�[ FS!�d�		.qs���"����������:IЋHplR��6��e�;�O\��D�V�VzY��P���tX�ӹC4�
��M�)�W�%��Mm�m�v��T��%����R4��&�:��V��Ld�n�,�L��Y��A�iD�!}zO=��]\��n��7׹�{|��wP��@�+�`y�kK{;�F��~o:���q+�}�g7�kP�{kV<�L*�Et@��;�Bb�rK�Xd�9�/���?]kK��wj<ºu��_")��xu�+������F])+1=���!a!�-m�/�X�2��>��j����&�jO�P��KtvLab�,O���g)KJ�F�������2�Yc��u�᩶�]�� ���	��ų��]O[u�k�u�c4mg)���.�6��@�|��ȴ�	�����x�̭x�D#�C��.��]Y;cyG���.�@��*���Ω�/T+m.�XD9�&5	\	�D���6k�K�������9�W����9/ia��+�+V�]|��v�52ݰO�mL���]b�Q�����������}IV$v�ɓ�wR���c3e��Y����J�]V�J�Ҁ�������cu�:�������8�)Y.�����*{y��=����2��� :i�o6�y��&r�*R�f�����`�N�^�Q8�od�km�̽޸`��Ҏ.2�Ao&�Ӯ��5Vp(w0Ks���]>R�^ �+���A���T�Y�}c�Q\^�ݕρq��ZC��Q��T��8H�aꋈ65���|Z\�ԃ�O��b���3 "�]18���x����au	��j�Y�f��]��P&��L�MIX�k���w�D��N�t{a����22��D�A^�/j�0�Y��H��˲�ݝ�RG�#x�T�Q"�b���H�ו� w���՛|�W|��g������c��=�W!Z�1uϯ*_gf8��x��D�y.�
�y̪�Ԥ��^`7�"y2B�X�蕚��H�G"Q6�m���-��Y�3NY9��#I$�E$�I$�I'z뢦=1�Q>�AdwB�c�P<q��QV,8ŅCl
����
��Őbl"�aP�YʡXKsz�CGVV�TJ}���&��Y5�@P^��4�Ht�uf�L:����N�4�HbEY'z��U*N�XL���T�#Xm�n�l��
c��4Ϸf ��X9n޳N�]٫a�X]Xm��M 
���M��x�t��T+z��fj���am7��L�,�m�d�t�hTAm,M�At�"�J��Y���QM�W7t��1J mϪ��ikKw����by8��T/(�tw]JJ �{�MÎ�ڴ8ss28�62w������j�rs٪�]Gk>jH��:�ҹ5�w�1�R�ʺ�5Y�z?3��/�>�V����"9%qnSH@��f|��ټ�����`���B�f/��T9�g1[���-�GP_��}M�9>��_��d*�ƖK|��}~H��
���;�^#Cّn$����~�������O���nQ>�-/��ɼ�t!��|.2����WT���9vSma�p��m=�&+y�p��=b���.g?F�c�����P��=T.�`�y��D�s2���w�v.m����gN!��5���	K-���g����.�Ǩ]\�>�%c2P'���Wg5\��tQ��D-�ؓcJ\���j/�����/`D-�s0-��_k�}���a�ӑ�e�ĭ#�ka7{s�q<V�b����ZM�h�ݽ�$�1���hڽ
��bi�H+Ys�7eGd���wc�h� ->l�.emd1�Be&�����|硷�BU٫�ʤ�������X��Mt��*S�Q�D��.��
�1/{�z^Dx�4���Yo��s=\�<�dĜ;�=4�!�PR��W�Jn۵ǃ-��u�u�c�Lg3gub*tGa0/O|�Wa��%í��upqA՗�ٹ�f�-e��Q+]�GH���uޒ�c���Q���co�*�L��oqX̭r9��䱜�'8����͡\�xX�vg��� ��V8%���7K��x��l���#���M��|�zy�hӌ� \���sEGjw���T�k���n��y=�6�FN�ї��+�D�2���ɍX��maH��M��zKR5�j1��ׂ��²	\���/����t�ld���k�v�<��{�c�a"�2����Ↄ��/*#Aȫ�J2l�j�Ƶ�H9m��\V�%tL�r���ThBAYo�.���ϮWTR(7�wKT����O%
v�br���W2�or���	W���[갈��[(�Y�Dc�ƍHwǩ���8
4�W@7��Z�gc�2�S�g=ڵ�I(��I8��T�X�Ϟ��L�L_��aS�E�%���^�y�+�j���k�V�@Pa)o5����\� �8��$^�`��Z����c����.�.�m@��E�y��dٳxsW2�F����xU#��B�뙭X��d�x$���c|P�=���gr��ȧ#�+R�$�{�ά�;}����w/�������,Rקj∿e+d^�40���@U\�VɿPn9��Dr����>+wQI�>��:��R�+��;�#j;�/��"Ԥ.*�p��.���z6ZF���ŵ$�'^&��jj�:�k�I]w�e�u2m��F��ip���A]^9wzU33�oL����rKr(����b7@�d��;���^*�m���,�NW�XP�Աl4-��
XGT��3\2��3��R^(7��N��Q��u��'5:�{lA;�d:.p��
�`a����Կ�G�W5���;��k=�t*7��Q�l�����+����U~�Nڜ��[���lu\ݸz���Ȋ��_L8YׂM��$5V���<p�����1��͕<WD��foN�7���y���YHA.��,RFE@��Y#�N�Ug-�b4�"�yP�=cR�<즷}S�}V=/��޸����QeO�C��,�M2�AQ���Gux#�/0���S�y���XX���M̅��56�:�JCgƕr�̎9;s7�&����<�oa��^�[��G��^ �/'\h�z3 "���FR}��[�W�P!��G5F	���Z�VP�d��&0�X^jI7�Z��mK����ɳ�r��#=yZZ�A*ҵnq�x�}<�Cǧ�KUaU�_�@t7s<�$�M��ڽ��w��n%IQ�Y�7��S
�4o��Ả�4݈&��Z�N��F��)lEm"mr�������c+-T[�<q�r�T3�Es1�f� P�,{ˣ��w�k$bvE�f�]��gM�C�qЪȤ.��_��X�(e�����bϒⷯ����[SsCJ�V���J�b@���'0�R���M*����ã��&8�c#_j7��.Z��UQ�
9�M:�ߑqk"�έ���}��pwwS�8�����2��*��K��=3��� s[�d)B��EYSL�gSM�f�n9�!������(����w6�>��pU#�w�/=b68%w1!���[]Y��hV�x�ځ�q� p�ʹ�7�ʭ<��;��͎a�}Zd2N����҂p�ZVC��x:�u尮0cV��yI��c�T�Sobz#�=x$�a�u�>�S�c���b��B��LyN�0ߺ�lx��QiыM�����)�.��ؒ�H��Tv�(�FdD����z���\�P�,l�$�2���?�"�Kܬ��+�r�YY���p�n9,�Aj�SA�^p������j2�5����c�r�4�Ĕ]j'|�]T�>�h<�P�oN8�ғ,E�A�T�([����"��}�����y���Բ�ЃD�ݏ9�	&�[�(dfTU���7��[y��̋x�s��ZK;u�":������<dl��ٚ�l�&8�f���,���qe�r9��͍��������__��m�+VzkhX�ŉ4�+2�Of��d��W��uO�-�K:>�'�.�zJ>Hi���K˦�����بb��c���c\�� �`�6����)��gtʒ���Ρ\�r��Cr��n�c9A��/a�f���ܑ�'go���ޝ�m���YT��ϰ�]�l/u������W��"g��\4�){K`�k�+���::�B��F���V7a��װ]�㹋y�N�87L1�]��'���u����5.��t2�j�Nt Q��ok�[G'��,�8���6,��x�q�bk�:ݞ��յ���7Vӻ����V=I\-�J/i� �m�)際�*��P!�V��r��Ҭ�b�Q-:�Կ{��H-��ܜӾ�댵�Z{�;�qb�/C�C�fj��Tu�[�%S�qc�$���x�(���M˩��%�t]ܜ7��4��jIkW+r �k$�x[/��+��g^=:x��ʘ�³�[�j������Qǡ�䟾�/x [���J�Z��gFEX�eR�	��[,P���m�1�ڧЊ��Ž���c�Y�#��>TM}g�9Y9/���P����E�x�Z����n��a���w�z:�Y�>Wͪ�K1��-���b�U��-��ΧUŬ��ԓ�Ow.��!GO�|�&��ߦ���L�䂘V�8��P�'����	G8X�0u�����ext�.� %�4!��\N�X%bZ� �J}�;��>*'>̓:r߃�ɭ4N���
�� ';�[P��%��>�Q���T�,���c�"��@��t5��n�qf�Z�+�k]B�vZ�Eԋi���sf�=G��S�!�V�W	�NA'$����2L��1&oapdӮ6���I.��JGn��ǋ35wS�]9�m�:���z�nf��a*anTTT�����]�J_NN���<"ҸޚU��Y�+*�[;V2n�;x�B�S�=����v*+��5�"v�!�^�#��/��/"N	%���T㷽|w"�E��ӗ[KP����\I��#��}���!{nE]��-T��؁�eB�gg	B���졷�Sl�3o��4�.�W$��Y?�fӔ���j��������GFь<yn��ܲ�������c���r���>�+p-��R��Xx��"�F]7�u�a
H��qwUgnAٹ�l�`���k+�U���'MC�Ԙ�����X�9�9����܁a��='�d�}!�p��~d����$�ŗ�ٮX�Q��L*g��V��m�To�ԕml	�΋�N�
��{�
�r�J� ��ݢe-�.�Xi����;soQ�sy�ۇ)Iz�{uWv��˴��i�$.s*��SbU�"�j�u��o��4\!J���r;r�+-��Wx'�������Y(wO��Y����;*�+�b�M}X�H�99-Օ�,��`�Pmcɚ�f=��G����ƭt��H�s�π�$�.B�X��ٸ�C'[uœ�0ܵ�܍p�2����oM|)ӂﻛܜ�LK� ��E|=v*�>.�f�#�l/P�A���/ܨ��\7�2��1�#F�ުVI��}��Owa�v��`�Kw@܏�l��2���$�I�&�GO�q9�1˃�U���2D�I$�E$�I$�$�!�Z<���U���0��+3�,؆��3J���a��C-�����x�bm�T�E�dP\J��je�̥D@Xi*�YuLq��Ţ���o&/VbcI�EY*�&Z6�T��1�eE4�L@�L�kWV�&�mX��Ee�m�I�,�i(�K��R��mZ�(]��YH�R��5ˣ	Kq�4�[��p�T�Yib*�h����IY\���L\�:��k%-+m�y�L�+SV��S�V��f1b��Eq�S��6�;b�B�.�¸�E
��LR�Į"�X�Kߣ�\������w4ӥjJ�k��G^���J��t�Ү�c�3bE/��z�� ��4u���ḫەk*����9��/{fGȯ�˄�#��c�j������[�S�y-+���%9��\�������izJTuE8J秏ы�!�R,�M�6q�b����I��}�W�2�x:��1N�g/�(�Qq����L�{�pc��h��m۠*��Cc��k=f�5���PT�V�bm-Q/4�{�b�X�d'�#k4e�Y�Ti�3V���-�K��0\s
��|�xW
o�KT�oX���ޏfK�*�KDG(��[~W���ny>��t�{׻��70y^β�'c� ����MHr�9���ښ��;]�#�im�K�jRN� �z�]Q��uo	/��D_w�gW��ey_hӚ̀2v�m��Zk�'S�u�E��p���q��Y�}ˑJ�"��q����ӗ,jE�u�A�J� 㙴�FEN��I��3j)1������y�"��v�|nvU{�u�%�nt>�i^(hk�ᾼ�:�MMoR����x*�k%�"�7P��܄La��.Oo ى��f+�SX˺5��u��Gv�Cx\V��Wݒ��h̽�Th=�S�f����US��3**�������X��@��J�ZY�q�CvK���6��α����|�.�.�'��]\�
�w`���]ɅJ:p����(�
N�G)�!�{�|w������6��쨔��y$������8��/�?���,�T~5�+¯�ɹ�����~����"�dYq���L��E�6���G;>����m�%=O`'~L!�W?I<6rƤ�����S��<����u8�F�� �݉���g8�sN�]p̦��#�+ڑ���YI�:�㼀�&�5���/4���%���?e�lDGQ9
a�T��"D,���ƤV�;��w�]	�kh�WY���p���E��NS)VAR����Wm�Q���q)���>N��{#;fň''�B��>�X����3sr�NB��c�9۔��&eIÏFr^��,���8$���I}����� ���/8VD�~k�\�
�p�հ5�^�t��&�B��r�� >�]C06CvȊw��هO��ⅰ����Ո�`nm����f��ܵ�.j3&�4�a�l�]5�����cF������і�*�͛=�'{����[�1�	���la��1�,�Qv�m�o0]�F�����θ)�~e����~NsK�^�M�K>5��űQD�ւKv��q�����8oU{Yٰ�i��ju8&�`x��~y4�zo��.���Au^[<�1Wv����*'MΧ*.�ڄ�i=9X���cQV�R�0�Ա��X���(�cT)t�9���eC�#�W�����#ه���v�JƯ�Ln��F�1����{�P4���\,;ѕ�w�q��S��x�>��G���圱�^㓧q��Jc��A6\^{��{����5j�*�c���䋛�`lΛ���>��or�t���q�ON1}��vd��Y��=~�k4Mh7�}9Ѫ�2U���u��� �)כ��Ju!r���WP���\9�)�c�Z��!P�rBF�g+5hh6�3�l�r:�:��0�e�)�y�w��C[��+��p�t;7�h.s�f�*:b)���n����\I�!	u�!u����>^ �2ˁ�&A�L���Ɉ;ZIfsn_X��n)t�
�I$�����V�u��n!~�w���`SD\8�Y�	%��9Kx,a�b���hw�&:�x��� 7J7
��8,q�.�6��/�a�\V߻vS��3i?vk�kKW��sq)�0�h�+ں\�`iQ�CN�@��G�קn.&(�[��پ��X�Hޮ`�-�r&(ע����=�q�v�]B���'��5�k3��t�}�D��w{!F��V+p�[%�/�|8��=��:���o�mY���K�_z���o�~0{�S��ɾ�&�$'�U�b�]E[����<&y|j���c�z�o<w�I��+s�`�+*�k��t�Cn<���`�\��b��|.T�F��JTt�!�Ԧ�:W4j��-=�:�Y[�������E��I}�G��E�v�.���l���d�Ԧ�]0��qk�/yR��T����fi��W�t�(����	�*�mIל�U2�Sa)#,�f�5>qoe�e��S+>�r����י�[���ޯ{y���+�q�?pЅS)@��h8ky�9�ԗ�>
� R��w�2��M��P���@��Y�� ���~��Cs7'���k���[����R��Yb�h\L����ړ��)\c�������x�|4!��7ִ:�O�D��I<�S�k�qwb�����׊��W*2g�hM���~J˖������Z������6jNc>��~�5[e��I����`׾qU�i� ���QQ|����ںWZ� �⤯�ӯ<��"v�~������J+�.�+7ko�_$D>��hqr7W@Eۣ3VI��������ѱ`����Z�"C$��U_Tz��S����}�p.:�eF*"��߮����=�'�1�iQ֓u�;�Ƀ�U3MWs���_k�ӷ\�� )}�C�{М�S3g>/�UE
��\lh�4e6�lZ*W�j�������]췡��Ê�3�pe��ڌF��NA�#)J��2z�u�+�eO�:�z�Ľ�j�
�6Oܫ�v�j��/y}I�E��73��9^�������%ų�"���S�Gr�I��wDֻ����Eh�W_��N������cVw�8Yj�&��a�+�1*cUX��|g+3#"/.��/-���wi�h��sGpŋ�4^��T����MG�T�l7a^\���^J������`ZFTU�@�i�cH�����б6Ȭ����G�����ײ*�J腓 �`��j��	H�y����Y�n)B�h��Xړ��k E۹�!Qk�Ǝ�(7=�*eq?]��K���G�w{��̍�3E�b�>ƀϳ���+��4�8,�{���?{R���Ŏ�������z�:�o6���3TYo\��ӭs�7��*k�/a�1V�y�9f�>�1���P�<��g��B~�*�̈��kQ�Y?Gc�(�����~��n���5����x�zpp�kT�w�t;Y�������{,�v{�z���8i�q��2�P��M͞�Uz��@o��~�>xr��1�WXĿ^]<�}@�K͛��N���j��
�/�5߶��ZW
�3��c
��Tc��B��KRf���ՠ��8�$�O����~�x+F�[�/%�!w�(�T�
#븴T@f���3яd#�3kU��[���q���<1���ث�±x��
�QV��%oq���x�=�����=M;[�]�n�(�$b��q�Ȋ+�K������n���D�x �<MV��ܸ4kk��5��Y觳|��
�
B�ר���*�\U�_.-�Y.���ȷ3�½Jc��³��,V�s��}ᢇ�R��x���h�������N�f+7Waf��1�fz���33f��=3�A��]�=��j�Ҏ
Zh��6�x{����@��}������^GG�L���t0&dFT\�ٽu�.h;:���T��Q��ת�uʫY�*��k����ڂ�������5ᢧz��J�ʽ�
�kE����W1���J�����hM�wz2�G����AMvKu��P;�,}�I�<7`�e���J� �훙��s�ʇp�z���9Fr}��=�w��߯Ws;�r�1
Y��^0.d��[�ˌ�	��>��|�$���ז�pQG��VQ1�8�7F�ڂ�K���4��e��q2�4T�ʷ ��nq7o:Nu�E��sT�3k8D�Ί��y*]a��*�NА�\��e��gq������u5^�*h�[@ws:蝜f �Ċ�`zmӆ�HڦV��^2�a�|���hY5e���
Q���h�ݹ���ψ��-�y+�'O:<ӌ����Zr�gf@����<��:���k*�R�+���J��jO�������z�Q�w�R4�SkSɿq���L����v�lf�yqdMe�Q]e�3h�����r���u�X�݄L�[����7�V]oٖBw�%gsӆ�*E+���V����o��=5`O�hj-�+���oz����+��b��O�M%O.��˻ט5�x�3̺J���$��Q�����2F!&ڜg;�R�t�v�k����Q�o�'�{O�<0[�ї�z�^����Wu䘮(nń��ɶ&s�D�����rԍ�$�'�3b��.�S7�����i���T����������q��r�����ۃ�o�+��������tn��V�v���8��
ޛ�4z
�p���olL�8����?�F�N�Wb�n�g5LmGJ���	�{7hYFU�;��H��Oa�ǩ�yF�QG�����b7��k&���\�K0���i=o��Q��Wy\�*����S�d,wc<�@�en�4Q�7��׹(˸h!����V
Χ���T	`�SGj��}���j���;9��p|�m��C�=2�����ᕕN���+�]l#�Lޫ�Dw\ԭɸ/�t��#r�rI#k�R7,���E�Y�`�E#�I$�I$�I�z�0�<�x�q
���R�R>f��[��5i�/�y*陘���X4���)11��l�m������Ҏ4uu�S-�p���AW.&T���ut��˔�������4��cf�qm��l�T*B�c.R���Xi�.e�ұ��T˔�+�֝fR�i��V��N"ѵ�!Y���&.X��-��D�8�Y�.�GV�%���.���*�-1X�S.a@X-��`ۈV@Q2�˻�I�2�@�i`��z�gT�tc�����E�����QL˻t��n4�,s.8�#�%b�]kA�\����,��,��s���ۯ����K�rdu}K����f7u%�8d���/�w��r9�HR����G�+s��Y���%ʖh�q~��}B���+m�E�%3yi��.�A��U���:.��+�hUÂ2`�ɱ�T0�%Qr%Ż��Zi�����q����K�Y�bod�X��r�\�8�JX�Eɞ�SB�������;Rzjl�Sw�3^�
&���&�){�q�d��9�d���Cu�\ECL��=�1HO�2�_K5U���;�q�U'^s"zmfh��lϰ�C#�cQb�2y��|��$��n��MZ�f�!Lt�Q�k��L�`�:�[�ɐ����>р{�\��=��@��Y�	r�<��	���.y�k8�-+�u��\SSf*_x�,UY��c��$�>&_�߂��������̜�G�,���yj�(TJ�s�zm+�1�flp[�NZ�|��
�rC`�ҟ�)"��!%�{ޏD{���]a��>��~������b��'�h�2L�:���j��k������xMF���Þ�V���(a[Lla�9;�W�h�����K��!P"px|����� ��_n�L�O��q�dd\>��&��P���A�4�����7��L���M�*����g��d�3N�v��l_-h���װ��6��H5�Y/�$��*1�S��j��)�����>��f��
����T~F���W��tj	�J��ca�S8#m�Mˍ7U}@}wT�`���T�W
!���²h��X�%�.l��z���E�OL��P�ɢ��H>ͨ0���ܟ���!U�X!�i�{�Eâ�)G�V�#C�^fS��܏�Ոz�o���T��u�YՏ7x�P��b�(ӣ�/!4_v���׳h�7&��oa�55��DQ���OGve�58�gh�I/���"=C=�o�uۥ�w��3p�i��B}a��Ļ���ў�b��/
|k�H��.3��?EG��Xmj��"�BW��vb�e�K�jL�*�aL@T��P�5!�جc��#�K̻5�.����K�EZ4 �/���dݞ�POD�
oɊC�! e���3]P�/�3j�9Ie�l8�)�g��ǝ��w�_3��%N����3���Ri�Vi>@�y��\�_�޻�������gܲb
E�0Ă�I�)��;C�,�H,�M8��)���4�X:������+�V0��CS�L`x�{��>���x��o���/Ҡ�Xj���O��v���%a��)�!�t۴�����@�AN��d�N3n0ߖ�_5��m��R���H,�]��W]u����}����x��bNeH,��ǗI��]ua�AH��RcXT�3v�a�R
AO:��q��A~aP�J�<=����C9�����;ߟ}�>!��ϙ5�jL<��,>j��
q��Xz�04�<B��Ry�<t��T;��Y6ʚ�{�i'�T7l�+4�YI�}�{�|w��2R˙*=e���"yj��[���U�M�j���D5�l��6�[}�8�*g�!�VVj��3�j�7+'"�E������wl���G�莽�����$��q�d�Nk)3�0%@�4<Ch����vu�1 ����4�S�5�r��1S�Au���j����w�]��~����'�Y�I�=a�8���T��j=�"�Y1�ISh���
Ι*t�R<N��Ӵ����bq���\Oy�u�������$���>��1 �a���m��P6{L@�*Au>�1>a�b
T*Ad�Y���F�I6�H)�
Ì*i�
��+��뮯�y˾��ܿI��I=�C�C;�z�Y��C�X03��&�2m��IY!���o��y��~� z���lR&���T��S}X|�3l���*O����H)��>@�T
�Y���V¤�N��v�R�tp�}>��u�o���y�$��Փ[��1&�C[GWkֻ�B�3�]&3����bAa�{t�X�5�ĊAa�
�i*z�����\�3������t�hVq��!R>>�	Ӵ����
��T���c�{�1 ��\��m��Rn�P>J��\H)Xz�N!�bAC�y˾o���k�:��s��Ad��.$�
����TהI�+�1 �T�i��$�
�UNά�� VVk��o�B�o�bC���p�پy��}�{뿾���P��LH)P��=v��+~\@QH)�,���C_RbAd�vbq���Y'���%M�@Ğ���x�
�h��;�|��o�OP*T��M�����J�_=q �y9L|`T����^Rt�!ĕ!�Iߔ1�Z��Rb ��d��0�s�Ξv}���b�v ��J�_��{q}��ʷʠ�E�B���t�w-�*�'k�P�cJ��9T�Y>̓5�I�KׁWf�i��z8dW���<��cM�ܟ���ꯌ뮷�{���bAa��Xz�
E"�û&!ĕ=gbM�Y�ϩ���\-8�n$kˉ���4�Rq�j� ��������0�^�����=������1Ҳk�1 ��<M�v�HT���Ì�Aa��v�'�To�1 ���:@ěB���H,<�
a�;�\���z��y�|������f@Sh��ghkt�I�t1!ݰ5�f�
Z���;N����N!Y7�����×�ԩ��1"�XZ��޷�������SH'o����L�H);gn3�<�4��H)�*J�NЩ�z݁���0㤂���_�ỉ��'Hb^=��ƹ����_�C�C��L`x�M}O� �Щ�2�gbu�P�Aa�|�T���AH��s�!�|��Ȥ�
�٤1 �wϭ�y|�7�|�gi=q �2�S�
�ۤ�����i�A`uˏ���08����Ĩz��������J�H,�ʐS�OI�����k��o�q ��*)�I�,;a���T6��}�AH��6��8�^�SL��t}I�-'L�
�q ��ӿ3����o＿Iۤ�!P�*�&2�:jI�PR)���S�
¾!��ef0�1 ��;q��zɤ�6�S�
��Ğ�S�M��fs~��������
A~��󴂃�a1��tʞ�_)6���AHn�G�`q�5�� �Ь��,Z�3������'�1 �����}��޺߾w���:x��AC�)�RW__�4��+7�2M$�
�I�05���|�^�<@�u<��:H,�:�2z�����I���k{�Y�_^�w��o�d�Ж((�WV�]�o��6�����V
`V�#�~�J��a=��k$T�R�\�x�}�;�v���kIZ�ޞ$(6�6O"��{�ct��~ �񟅧l�J�d��c'R��:I�����H,3�N�*N'[��t¤]��L1�hݓR(x������5��}���y��_}�9��6�C;�*};�bC����Ӥ���>jAHo��d�ĜB��P1E��c�@Ѻb
E �d�f��
͝Y�d�+1��5��߯����9}H)4��t�Y*
E���
�8�T*z��bA`x��\H(��{`T=�&%@��m��m �3����~�to��]u��g�t􂞡Xz°;jt�Y���N!R�����59I�H)ה1 ���SI�I�W��&$:��ěq&�AAH�L��}_9����ﾽ�=� �@��3N�
-"���c&��ۤ���������jw��IP�<aY>e@��1����
��1"�&|f�.c�"*cջ��Oݸ�����A�0��.$6����PR(]�b��3���U �;��&�$[��ɯ����q��!�
,����L��>λ￹�d������&�R(%d�8�^0���+<=�I����x�6�PXt��S�
�wHI�>N��H,�e~@�ߝ�֌ۯ<��|��?t��}`T��OP/�>����ɮYީ��}�8�
i
��,����7>�Ci;B�lJ�l*At��)i�����{���>~�z]��=�߃i�I�*��J�_�`c>I��%AH��;��AO;�N3N$��<d�1����Is�4�R��f�T+3�_;��s�y}�L�2��
��=OR)���4� T7-<B���I�*ACL>�� ��S��8�J�S��T�f��哌Ā�]o������X�ٹYB���$�a%���7����;��x{�]�&,A\'t{]���ڊ�B�����u���Jp�{0^<n;ݵ: *\M9gǎ��8FCu��Q��ܑ�'���ﰒR��|���Z�S�J�MH,0�'��8���wM$���gL=LAH����2tʜI�(��
��W[��4�Pה�<v�2T�{��>�]}���~󞇉8��.�H'�T��$;�Lt�ی�2�AH�07����^S�t��2íR
��t���)�]���������_Ӡ|�j���ELxLELxLE0�
���Z��u�1"�P��1;@�<{ݚgL���R8�N%@�)�;>��AOXh��$��q �_��}ֽ��9���6��$�Ă��}gɤ���������\`VM���l���5�xAH�4e�aS+���0�l�
f���3�}��o}}��q �����$��S�� �4�Ϭ:Ն�'��,
ԃ��ÍH)8�ی:��!����E �8׫d�T�:��w�����ϟd�'̩�x�$������6�R��\g̕�J�S��*O�8�R
{=�c��0߶��|dєR
q�����_}�='Hv�Y�&�H)t��ALN�t�A`z�\�g�6��*IX|¤���0+PXg�R)0��z�P�+<d����s��[{���[�y�� �ԝ�w� ��S:�bAN٬�FO��L?����6*X�3f�N3�>�����d����=|�H�}f�@
����^�5 ݾ�o9v}S�/�jZ>|X�@`�G��]a�,H:P���ů�L$be7���2.|
��F�ID�vX,�0�Q1s�3d���U®e�>��ec�~����uҾ|���9dq�p�'�#���#o�[�SLj�u�f�.�����_x�+dm�C�^id�@5a�]7�~8pp~��}����SU_��?<7Bj�cRo�����L�+o��~�5��TD��0�JN;Q/�Z�z�j�T���	��}Ơ�(�T�׹IȓsJ�1�6�2UH���\;��B�l�N�3Y>�ˁ�z���5ܩz[�O�Wq�w����U�TA�ó[�G�D/�'���]u�d�u.�U��,E5Q��ʅh@�,{�����hg�U��Mh�P��²���d���["a%��tsSݥ����^�d��C�L?��IU���\5����9�W}~��ڧ���2pXc�B��z��]yW�*ઉ���QR�S�!6{p���+���D:��!�+�Q�0Ӑb�����v��]�h5�%�	S6�!�J32nJޠ�M�[*ĺ��D��f"�_{������@m���S�uw_��XUg%����G�M=��W��_��p�Ÿ�0f:oU��uEEU�����J�~�V凥��OrX ��<�x�m�h��#��=��Nf-D�I�<�u~j����s�*���L��K7����+�:�������yة�p��ߺ�.N��� �F@�f���I�Ռ��io�A���eC��Y��hR��]�
ʆ�z���N�"�=�]�����L*8�C��Ѣ�/�C��֜���㝛6{���������^~����3�P���H��Ui��s�����p1��9S���=ƥ+GѲ��@��w��cF(]��j����a��f]�ӭ=�E�Zq�� ,!K2!V
��e�՝�=�.��]���P����/i�U2��%��sؤY�Cۓ�dF]M�:�&�+rn�{k�-)Fޥ&�� 	�(�=���x�f��Z+�|i�	yR�z`�Q�F��.zr��Vԛ�ti�9�W��a���=���ka�w/�</C�ӽ�ݜ;����zΏ]�0���4��Rg�\_iۓxuNw3<)��	;��X��%J����t&�
���)�x�@`�S�G�cq���C�����W��ꪭ������ę��#����S5D��ʗ^c�����r�*��}���.Ta�4�� ct�PF��M"�Eȕ;�j`�r�/¡X�57\97M)�@\e�ҥB��S���b��  �X�������9=�%Ύ��U1�$����]W��9�Ff<���[g'�̑#��
țk+.}qay�in�A�&{-�����R�Z�/qvaT���O<���I�IdW����kh]���9Mch]ZHv¢��7c�%S��&��I^��/����˖h�(*4��oG�+6��gs�KQ��Si�&�5]LXFk��o9o�`͔�n�<Um����/��q�1�\��25z��QȦ����j�ù(i��֫;Y�f�^KR�pX�MEleR4e�Z��a�8;9�uvܭل�G�خ�7�^R��ͥSy���*�����A���˺�^��sٲS�hK�}���qc�F<r��˧ח1�p��E��1+�]kF�xv�pE�}���u�%�mcއ
롶�F]�u�	����G�<9=^�ZWZC��_)�]H�9d}�,���=�Qx��:��a1,<���t���\v(��vf;(s��͘.916����-T�%rh��dT�N�F�ӧ9�me�6���
[����~M=5z��"S0J��`�|ĥ@B������774$�u����R��)m��5}�����Ӑ��s����)���Ol����R$f��[��VLδJ�y���K�j��7�s �t>Q��}AD��p"�v�B���S9�B�^�J�ڷm�]�UnD����TF�]P�븸�#|D/))���3̕K4�0�U�Î��ܻ�R�0���7;n�#|p�Q��Î^#��:;�4���:��38��<���=�*b]igH�lXI����q��Us�­L��U�,>CFF�ͭ�ZJit�9��o*-ZI[�l��0\�T
W�6e�E.�b�|L�?_	"��� ��K�ssid��S�cV�ї�n	:I$��"�9$j=N&�1QaI�N��G��8�rI#��$�I!�L��[B�
��Ƭ�P��R�iJ:Mj�6�q��\h�ˆD`T��mDV-�(�3&T��T�Q�Q�e��Yr��mn�q��w��J���E��Q�\��-�)�Ă&2�V:��!�f�(�KZ��֓E.93Mu�00LK��b�{��\��uq1�)�Q���r�VT5KmT4���س�Ӥ��s$��Aa��.�CJ�j�V1��j�aQLLB��m%�B���]�;Ը�q���,E�68�3��CY�[�H�f�R�	X-Ƙ�D���q�7�����04Ɍ�m�bRP8����{��y��>�ݜ�
�U՝�Xn1�X�w*�_X�Q܊e$,�I/؏z=����_�ja�����f�T��HT�������3���ܮ#c�0OLu�i�i�0`��x)
j/��t����~��?\<3Ơ�L�.���R�9OEz�
<���#~ 6��v��~UY��� �f��U]M_GiC&�/�37����?�
T�L�a�"u�9"c�J̸��L�Z%��-��0��^V���*%ad�k�~�B�v���������nJ�&_��٧>�^���Y;�*g�U¶w-���s:9�O�{�t�.{�˼���H��Y�	@�W,v��I��灮T>�
��O1	�T�Y�1��]j�O��f��|t�yV�e&�S���̕�Na�uμ"%���D�,�NE^y�@��X�3�k(E�!�`�e�zb�@�	,§'}�l��pÔ����ZXw6��F�H�N���@+�����K��-owI�7�Ȳ�!%߱�{ ���꟨vFz��g�+r�ͼX�|iʙ��Q�O�:|��c�=W��*ƨR ��i
�.�1�H��`�\����{�v~�����oW�
V`}��@�½��<�~��eh�O�ګGι-:��BՔ�;>#�m��[�Z.�If��3Z+�S�pԳSZ�����ˬ'���-Ҙ�5�&vX���ّ �c�7]1��i�����s�tdm�5P'yJ�Po�eDn��u\��8&��^�0/�Q ,5ਗ਼�/ܩ}P�iKS*2r�k�q�\�5��{̺\�ʔ����@��^����ԺŸC�tWm�Rm��hKu�]�K��j6��P�g,;VP��<���C����&CK;+{�����5�8��+�F��t� b�p�>dv��^*����:���ZQ⥬+q��[�˾��t9����V��#�W���z��[��}T�/�ʸ�Zkʯ�ƸR���@�L�'/�AƳ�8_����s�(Q�]Ժ�t|�R��^5�W�'A����ۼZ2f*|��u�S"{]��*F�TCu2�<�H�]L.i���\,����vph
B��<z��˕p�+�]�����5Lh���#[v�!���,Pn��9��	�݄��"r��W$
��X����i�f�R� 痠�&X)?{�$�pۻ��`�f�*�[��u&Eқ���T6:
E0���f�d�p���+��3M��C�O-��70�݁[������GK�k$q*2@�[-�Wi��n��J]3P/��H���^���о������Kh���;��<0����n���;��.���F����G8*D,��'k��s�6I����!�5��`dn�-MN�WV���ܣs6H���z=�ѣ�n�A5�tبɞ������/g�����v�m�x�j�Z>5�^u�CT�H���x!^������������6tz�:�x^V�yђkR��}.H����9W���<�A�^�v~Ю�3+��;WN�\����v�E�0ھ�َ��qj��֚��~2hY�t&�lQ�Aa<?(~�M��H��ʨ�4tkp���LKY5�8�4U	��VC�Vh�T�؃]C�Yʘt+����H]��w�u�T��UVn��R�Q+��1b.਼֡��2�h�b���Ƣ]��wJL�8>+��a �a}�e���� ��KǙ�[�wd;�>�꺾B� ��	{p�V�$�W5���қ��fq܀N�嫃���+�Ig\+�en�M�˂�Fi��q���g3�]��� ��K4�lJI�_}�vgh�f��Y����1τ��S)T(�FD�I��?��7n���4 ߁�}�Q��~M �����+�j�C].�*�S�{��N"bC���U]n�����������d��{"s��b��.�k��4�~�>�I+>`�K���+����z.��	�T?p"q��Aj,�i�ˣxNA�W���Wk�'�s���Ny�KqU��Hg��{^
B����$ay¯;��&`L\��>%\��9Q���k����n�!��y���4�&Yb�|fuҹgEnW��&>O|��~\_�y��^���'�٪#�_xX�5�ɭ���&�5���p�3`���.�*%a�F�G��ңj��滷~W`ԩ-;��*�g3"�ʚ5]v7�y#�Kp��)�kn$�q�:P�#��*��(�J��:'줱�vY�Xɪ=�ײ�p�fI?_}�P�H��w
#F��G��3�Ç�^?&pDX�ꃕ�U��6�g�n�[��YQ�I�g���/�w6b�����;2�S@�ӓ�Tň�?m9��v)mCU3h�_�i
�P.����JWݥ����l}����1Jp^�^ʮHk�.3�@;��2-�n������ ڦ��CÅMW\�h�� Q�5WUkY�w�����Q�uV*4�3b��h�aBu\�%m��+�0�~��{P�y�u��q��
�=�dS�X�j�/�Y����\X�@�(*G��*ɘ�Y�ʋ�y;��8H^ł��R,��[�����{-3<)7�V�����]e1�C�Y�ͳ@ɪ�O+�)����S�VNy�%Jojly����
Y
�y�5���V�!`'��3�mɘ`t�؏{;���X[�ׁ����[v��@�-����⾪�wy&���N��~,���/�/��N�B�@�疬w�� R�_x�!u"��+�<sܩT?Qp��=X�Y��d�>���c�̆^��*gd��5�^�
�� c|��{�xg+x�A�gB���j��by�38r9�����}vn� WO�6ƸR�����J������ۦA�
����`��VC�c�>��V*��up��m��o�
#�|��C�b|���=�U��)�%��o]���#/�+��UW�f1�y���.��J�øqB.c9��%�fbC�)��4~����,`�J%{σ�%�t�Z�-g�^�I�wq|�H�37��,4��V������ݰ+���m&��ن$l����+<����N����o��|Y9%u�M���y�-H�څ:]6Z1<�N�*�Vn��=Ep)}�����Ss*�O���>�kM��>5F��
^4i�*�P�͞��Ɔ��r�wS���f�[�k��A^G�lzu�yY��7�CHR��8�E\�*�����X�5Q
��'���Sp��ƺ����q?,h�3�8e�s���&��DYQ�����p�,>���8�t�O�/ƱU��l����7׉�y�ReφR��0�T�CT@�X<5쐗3��2}3��oM��i�<4l=���k�T0g����;�8?Q�MQ��4��^
�W^���ā�|�;�*jc��o$��ꠅf�
�5�F���Lj?A��0�эU[Wf����W}3>��,U;�wh;����0'��ͮj�Ѩ����'C��u��R����V���-����t�}KR@�}�;��1�*31�I����k�nܫkRCd��VI)���� �������L��Ӹ�t�
�tiƐ�y��ozd�U�l�k�򥼪�5av���J5}^S�&�P�8S/0�E�>��Y��U��@h�W��#�e�E��f��~��������$O�Z��h�F��ɟl:2�s��y�q,�C�jr[{>��>p�PƝC�~�<���K�ϲ6c�-�d綔��f,����R��E��}���e�����>e��?b��j������ב�����כ��U�����E��
<>�G� C��[w��To����Str6{��u�5%W��ƍf�5Wl��|y'=ܛ�X��S9���nLt�Xu�TÆ	��~y�sTk0�L�5{eƶ� =�u���+AJӀdzm��Y�b4���le7�R۸�WF�b��`����;��h"6�B%w�m�XD$��v�91����2����cr�P�Q�:��F:"��лsi��+�׫�D�L��ʨ畆 �������*׎i�~�o���yQ耤�L��TD�|���ܘ9I��u�Ǫ5^��8֫Hh~�@ }v�`��I���DV��hW��k�^�}yDp^<>U���	tՅ���XQ�Ƶ{ܔ�}�SB�
�	��{º��b��b���BǷ�����V�������dϋ��D�s1f���UQ�U&2�D}��~����Ֆ
j�uɊSB���yrC]½��:ie�w�Y�?p�[t�M}c�j����G��){	�5 |�����qJl��,�فU�cj��3Na�{���[T�0Κ�T�����W&�)@�,'�8�w�r�t*W%m(�t��1`C9-�8	��ٷyWH��ͭ�!�,d�EfZ0Ι�r���Am֐
VF�$i��t�V�%����g�-�W�.g�ݚ�^q�]���/q&�VD hͫ.WR���Ċ�V`��Lo!3�k|����P�\N����W�YKb�Y��W�	яZ�p(�����s�����4T=�if2D{������+��nжBԷ�r������pWD劺s��t�>�*�So��{S�vҤ�R�u���)um1��(�\';�2�c(3�^�&ћ�F�XH�u�6�ˤM٢�KN��8t���e\�!je���/������+R�U�S ��z�:Ύ�+��#e�G)�� M'�N��3t���a��a�*��`nGu�!B��������Ux)*��T�8j���y{v�T��9�����L�8l��4�:�ʫJP�U�[h�Gn���q��m��{��nI* N\� T9��&qȲ�7���k�񯷅N=��t:Ik0��H�oU3؆k�.WU�FdX����19ԷΜ�L@�1um�h> ���R��ֆ��X�����.,�,�[�D�g�˭�X����7���"��;��5X�l)v:2m�}*�sUW���Xk��wʷN��S�G�*5��yNKw^^夒�7�@��˩A v���q���I${�tN�\dDv�Ȯ���ubrPI,��!�0Wn������C��}�c-����2�V<�sT.X�V�m��e��4�R1��cC.%:��e��2� �/:��՞M��z�n� ��ݴ08�����#�H��'r�#���9J3
(��I$�I$�I.I/��8ԗ�9��Ɗe-E
�"�َ֖!�����C��Vi��"ȤQ�
� X/��Vm6���QYR��Ub��b�j�JуiPU DݤP�J�l���R)��b��1�Ŏ��(ɫf�7B�7��`���eUX��
��Fuzΰ����t�EDDQ��UDE4��ګ,�5in��Pca���["1�E6�ib84b�쩷��k���޼��뷳}(Ҥ���p�M��@�v��0������܄Hd���Wݙ��~�sbȭ��a�׌��/W�b ϡ�Y�68�r�f�B����X�Ś�'GΫ�� ���f`���6|=\~����+�T?E^T�[���[t&	qj��I���m	�sѴ&/��*L���>5ّ �d��_f5��h$�q���D��U���5�ʠ�~�ব���N�����#;o�ΌŊ"����v�y����F|a���ۜɊ{��������l�e��@zXUf����t�Z�
���[�S���M�)�8sKW/�T�Œ|z;���*9/j\�U�nz��U
��#��B�s�8�D�绞��ܥꤘ��z��&�Tr�[OP����C<��=���72�ux���Rǡ��m���y�BW�f%Ƨs}H(���Y2�<&��n�4��b���״&�F�\��%]��K�z=��%�
~uq["`��\\)���/J��z�*�xu!O,�פ��I� �O/+.k��5Ģz����ںˡ\�A,�[��qyI���UxT���:���,`�M�@l���&��<J��1*bU3w �T��X���@(hx���v�^����|>�t�9�C�5[G*�7�U��d���=���?A�O]9P*��������n�M�G��z��Y�)/+�u���*����ᷫdc�=u�n�- ��]@�2�����F�k�Y��4)g�{�
Υ����Ǚ����-�;�xS���Q��.�_xxV_������>��0}��`ChT�C��@
��o�`�b����6�mr�	�<�6��B(�]���cOb�iK��\#�՘�;'���i'nY��Ö�7��h��J裬d�-��7'�}��i��t���Cf�zlxA�i$=��A[~�}~��;k>��ǅA���O���-��2�>fEj���%>3a��ł�V�B	K�.7��C������S�6��M���D?{��)`�= +�d��Fh�V�G�l����\���y|]��E���6��43{Y�Z����'�(�޿�-}p�DmTl�FWT
����)���p)�)�.��MW������v��6��g[����S���w��Y(}}��ڢD�u��I��t�Q�>��Sx,԰��,�U���8��/�b�^o��8 v�q����o�������@��Պ��ELX�}�n��S�T������<���Ӌ����=�@�7G�a��Z�L��æ�.�N�g]��d����S��[&�A�TFH�[��}]}F����+H�VO"�碯��驩ͨ����5QP	��q}�?<�	��pw�{'����,h~?�c�ќi�t*�?E�J��{�z�%s��.	�����:2 ׏7��Xlh{j#WW���C���^l=�rj�����xM�G\q덜f�$H�b7���)��b|HL\ñ~L��D!��?j򩆵3o����H�T������˙��7B{�r���*rb�n�NA�ID2��6���7TϪb�:#�"��ޛ��v��[=�;�kÃF���\*2D�@>�~�kj�1��3�źk��^C��Ǉ8_���?�	tՅ�޵�q	I.fz��;�p�TT�EW��s�X|`�Zk�Y������2u��ҬC )(�1xt ���jn��X�6�7�]O>{��D�ջΩ�x�)�B��
q��^K�ԛ�V�{�ZL�ѽ�"��%e�BK�����O���U��0R��o�y*5�@RӢ�ͻi����U�����;7>��ɫ��X�&�sT5U$��O=Ժ��mP"�g����Bۦ��Ɗ6�@���^Әz�mI��XJ�f���H�f:��-�P.�`�&|/���VӬS<#�h��ؾ^0= `�����tN��3ڗ��xk�  ��K��4X�{1��Pm�.�&~C���ѱp�~��bA��X+�`�]W�8wd�J�hvf��FOO=�Kdu��%�ۥL|�~�ͳ@ɪ���&bo^�xJpT���c�L1F��l���`�ʼx>��;��|�F
�y���`��RD��b��{�e|��tM�4Q~W`.w��\��.auf�S�����6�'��P�Ďm˳�C"ݰH�}4�p3,+Bܺ�u|s3�oS���W��w���}��}0�.C��3Rr��U����1���m���Ƨ��{��猍`�f�w��Y������Vї1�!�l��t�Fzr6���zeLcW
�B�ՊsʡL[�h̛��g��b�5<�V���F�ޚ���3�b�7pj�\ˑ,T)s
rD�O�qp�����a��<k�ó�X}�wݦ�� Z��X��=j��M��f��N��{u�;�,��{*]�Rヸ��#]v�!���,�b�޻~����	�Rf%P�7q`��1�j:q���^�d�N���Z+u��7�X�uR�է�]T�W[�'���̚���PX��2���P�}���Q�1%���	�7cw_+Q(�i�YA8�C�FF�G��r͞�|��.�	�6�+Bk��!-�Ĉ�a��POUٵ9F��(���4	Ee��_G�ї۠6�FrT���L}o]p�}Q��~��'`�Ȏ��4<Bm�yąQp�8(X�>o�F+�,�G�5����ٕ��N{ֳ��K�,Vg�����߮�g��v؝��9��r9&S��ķPV�<2��l�~:9��Un��@O+y+��G�R�~�����\�����\�:2M%P��ܴ��e����F���p�֌���pL�^�ej�tY��Ww��l��,T}�7#*9И��{j�b�^H}'�����t���j��g��'�g����0Rf~UD1�&t�����ʶ���w�3��H�hRw�!�tkY��=��y���r�������J�*�*�i��`�X
�Qu�<]m�'�lk��hz3����^�X�qP̵	qɂ'����O�gE��OR���#c�B\����I^�"x݉7�#r~W�I�˓�?y�����9s�Q*�L�Q�lMO�oH R��[[���jD�VO�W�*���NUW���3ԥ�RL��Ν��6�F�����g��N�sw���>�Jd���w-��]�_X�s�4�g�\�������nK��ơO�M�2�UN�h5�ũ��n��*[Y�n&`�Aʅux/ϫ��ȕ�Z)R"m}�\��I�ϖK|(�ں��>�=���sK�2���f}��cGZ�]1n�l�����8�ħ�	to<bZDq���Z(ށ�G�Bƈ�ׇ�իf���##�!��I-[!���ק:rF�a�\�t;R2�I��[F|�\�'��x�`�X	�Q]P��o�_���u[2�ª=�u��jd>3X
�X����D*���ӛ8VR}c/��F�O/
��B����U��1�dY�\����Hm\�9��`�S!r�k[�:%N7�r�H��$��ҟ���?�n��?L���tOj�B�Y��U�2L�����6���vv`ȗǹB���i؀ ����y�x�
�)���}�pU��I� R�6��u����M`�JH���V	��2�u�Z�W���q/�����/�w�;��͵|BRs��~^Ϯŋ\6�]_@�Vҟwb���Ku3y�`���{���}u�a�d�+3�������26�2>�q�$�b���ie.hLͺL��e�-�������A���M�n�<[�"���b�DW�ۗ%*���6kU%Z͍NA�%2v���>�_�EC��6�`SP-ו���#���Mim;}0�fr��fDØh�NTV���KGϋCݻ"�`�&���F�v�����G\i|-�w�N��{-�<��]J���e<�ն���2�a�� );�Psz9W�(٬7�c��5$�U<R~���!�2��sܫխ }�0}'�8w_��W{�{8׾k�㔭����1.�G�S�9�Jد*4+]���X&��=�^U���݊a�C!�J���E�������j.Oz[��K~�F�Q�m@�0\� ^�O2�X�·���AAj�Q���A�ɶ�LWY$��UF� �Sig�4�;wޞ7^gG�?��Юcl׆�8��A�.DZX�\m�0"Y�qR"D��6�2��UJY��S��L2n9�۶�M�X�좍pR��;�;t��.�:A�׳ڗ��&��N@/�i�V�_���@hWˬ��ʕkob��9�zMuTC��d�S5Q��A���d�;�?��h3W�M����/n�̪t��F�9Zv�RĆ�P�Ś������P\	�!�����2�(����a6��	CKMٖ�Z�S"�e%�ۨ��T����ڵ�.R�J��BX9�� 4��rw<��>�s�QY6%u˻��	����6�D��&�Dbn.�Шw�E��o/k�v��ɵ:��	x3�һƯ�3���Yqiu�ȣ��t0t��\�� ��UAIT��3S��4����pk������$�T�X��������ղ��u)�e,̂����Z��-�N�����%�H_Ll<�V�����hQic��
_I�]���4��N>�V���o7zl�q┺7���fށ23+0�|9���"U�2�.�hP�sm	m\�I��.Te�t67��i$�f]��l%j��b�"�Sf��M4����۫�U�RU��dCxHD�q#.e�Z8Z�#C }j�d%t�2���
J�6���̺�6ͳ�r�*�Y�.a���w���J�¢�dq-��C�CP���1|�k�;G���S�J�sys�Iܳf�u[V"ށ��^_m��������Ԛ�@''���x��m�S����IL�%���V��˗LJ�06�-�����`�뷒����w��o�� ��3*^"���_Qq'3�f���Q���Ǚ�"�>�n'Ԋ2�:Wh��5J��#)��n��L8yU�ҭ�ʋ,PHZN��޵k���69mVur���IP-W��_��%��4ZBG�;��k5�����3]v���1�h�jQT����}���균��3Q�9[/X��un�d���fRn��͝j\jCjM��)$r&�1�$�1|�8��圛(ܻ�r9$�I$�I$�I�w��m�]]��`����$TVi��QQv�Z؆Z*,Uf�cTb*ƴukZ�Kq�,V1�@������%A�T��5J���kR�TQ�Zi�UL�b�Q*�(��UT��[DLeb��c���1QCEժ(�"ԥq��Lfd[\����,B�Q�]�շxb�̴U��V�,�X�ձ��Dj#Uf���B�޳z�TMZ���҈����Ab��b���U����m��(�UTTTF��1X.�U��2���	J�n���T�2��g�D�nt-egn����n�`�Bp�q�|�9M�I~D]�Â��V]~�>�C�e?m�wuY��a�t���7,��H��"d�����Lf9�b���*����4�㠖�K���wg�Cv���W�π\߇�. *p<h��?��U ��]Oeq���S�LW����s0vC�} "<5������==3��
��<>�(�T�_�C\���^��/a���V-�b���ڋ�5��׭�
ҁ�^
�dq�V2VP{+�X�������N�;:�
���P�� ��b]Z�1I`�Y7�{p�l�b��R��t*�O�R�t%ex
[���1Wj9}ӷ a�M>��� �Юp���Y}^��:��p�U���:~�xV�GD��ӫ5�3zfR�H�>+{ǡ��q8�k$��t�f�޼���dv��W*ۨD���s�7o,�[�@�{�TT�P؉������%�=�]Zn��]r�|��(������v(O�Sn��왹9Qy�
vk1�Vq�($'����_{��c�~�C�8K��>�G�� m������SI^���{��~��/�j@~�/�3�/.�!J���E�X`��Oee{��پ�Y��1�	�.U=쬂���
�
�5!�T3�,��>��Ί^����=<��C�#�6:pwH �ےw/�6-�a�W�~�~ۉ�������
>�B^nw{,`�^&*���<�[�s~h�3P����̽����p�!�� c|�Ub�j�r6��f���6��9�STLC��A
�/��X��Z�
�kEq*�.�B[�%Y�
�Tڡ9=-׉�����mvR�n�����EsM��ݜ��ot-�v>�X\�afI�*�CT�Z��)�ğl��{b��z�`�J(07c�32v�}[�T���{�����z(�bRO��u���X8~ľ���王ӂ��y}��y��R�d����R+�ׂi`��h�;M���:���X6Z��^�&���2����;Qq����Ԍ��&vVV��j/� 렸*5ұ4}&��]�1��K�
�OqZ�ѥ[{ӜCM�J�f�X���~v(i�7�nf.nb�h�[�`-U�-*�/����PpO����®��V����]� R���O���AN����ڐ��4�J�7%Qt�׵��m�3�/FЯ"��UʱW3GO�h��*�@-j��D�m���q��x��!\\2��j���w��@%�h���N�z,Vￃ!<k���A�8:�I�����Il���<�yC�W���:�a����WI��|��s����CRE�u���I�FS�:��]3���=����[�cfH�"�h�ӳ��g`PT�â�f������t��hxq������u��ҫ�
�T�.B�\�oʩ���*�{�wSgw�!��xP�
x_: ����<������V�{۩|G�z�̼\��k/����_%��F�s�]ɳ�ף}�gYtϡ�x~�$+: �^Ҿ�輩��8^$�����ZfW���]�+)��C|ˎ�^��r�!��['`..�8�ٹq]Ɵ��e�b?7b�B��s�J���Z��l�a\[�b��kgt���ڟ��E(`�lc kZ8���^D��)��1.��_�������ePk.�%	:iX��x��ΰ�ϦWxu�pRTq��
�y׵�X�8!HڇY�7��^�fb���7�a�Ot���W��I�5{���:2�G���ͩQ��A�W.�ёEm[�Fu�vԩ#�6��r�s3�sr̈́��DvŹ�#ROë�O�"�4U�c��Moo���2���̖n����Ц����"�;uL}V���7���3���Ջm�H�92��R�]�ڨx�*6 �G�Y��1�:�л��1nz"{���ݸ}H��J���
�� MgT{U��M���'�P��~�r��묺�=?X�s�*�@nl�j�;���}��_[S+�ɘ����dC�S�[��<�[o+u�Q�����&{��n.5�AV8�x{b�p�AT���Xx[��}��}�/�h�>��u�k�)LȺS"��vޑ��}S���K�m��E� B�����5��u���g1mq�YU&s�$8vf.^�Y�3�
���V���d3�y!Y��"n��@R�S�avʎ�sN�Ut��'���{�]���]���^���֕�uv+3��#/-�\���'G(�/ػ��c�9�[���[{%P�1���N����5�k�mm�5_p�5���p��`��v�����!�G��s�;ݕD��ɯn����n���rg�\d�igoJ�MʛT@��.��1��*["Zc����on��ȇ<ƀU+0����MI�0�\���]1�1s�����#3�eP*��,�1�-��|�־֛��)S0j����S�g�I��v�Y�f�+�J�u�%y!N��b�[�u;e�'���\ϴ�L4�����Q�Γ�TXv�`����j�	�u�W
��e�l(���o)k��sv%\͚&�����I����h�#����j�
��*����}�$D���^Lϟ�J��';�2�$V
ڼwu���I��z�Xk�2�G��b�������t��&1�b�iof��vޓ�%c�ajgmm��I;��o$�x�_����J�Й��xt%1��/�p������ܓ� �$<;���?*�5MS4_�h�����
pl��ϲ�]6%�Md��^��75&`�B��Iؕ���IZ��/�H�P�/M���uX�:/�>2�R:Gağ�/����׷��>F��]�nA�![*o ��F�k���Y���kC'�|~�C�U��
>�h�,��]e
˟@m!�KEb!�q��5�5���'����o=��E^U�V�V���"�Q����5I������l�<|=��v���Y��` ��q����p~�����s�i]{���Zly����{W
�Q� ���p���zk�r�vXí!
KRc�ؾrg7�n{zuvl[W0f{Fl�R��&���M���U{�Ҧ��{u�f���69"�	�+q�:K�<�,Q�'�}�I)�qB���J��~��Xr���2��I�좩˟�{��t�����xr,fQ�O��]b�f�-\K��&[��S6P:J4�˺�X�M�z��*��e
R��gG���Ý\
�5�i��S��S0�џ_����ߪ�&���E�Us�����d�>4��K���p��59�/7��B��l��n��}�p�%:�!m�8$�*7e�$��M�<cc��a�`���p�\�t�z��`�k�[ыQ*�k`)�Ml�*�L��p\(��wk�i7՚cy�.0V`[;�=����	ދ��{�^��!ޗ��=�o7ަ�A� 	��k���X��#\�����{����,6���\WWu�4
-ա��
Er���y�:
����3`$e�A��J8��W$��wcC)ά������|4:�\es��xm�8�-��=�N�^y�RK{+o��9�[(�p/7��w�)��_i%'J
�]N�S�L��.��0r�t{_�K<����ɩ}��R87�U�/Fi�E�TJ�r���XM�wNC�9��W�;q�^�N��]35�95vdԓ��8���+2&�2s�e���QOZ�A�n$��Q:�MI[$!�Z5�%���q�[e��
/˒C��󙪂d�����y�\�+�GQ�ڶ��檗2�y��o|s�!�ߚ+z��a�Ù��/� HV;��������,ͩ:"����Yi9p�Z��w�+�(�8��V�t�L�����QI}����[;�F�٥�Ȉ�
�
# ��[LirN�����1�G3�0�����Fs�o �^�pءf/`E��:�k64��O��j�n�tV�:�����W��x�F�v1���m��n8qs5�'*l��6��'�Q��wj/I�؎�eX�7^�"�[�*$s�L������8���U�+�5�q\��#�����ޞ�"� ������6ܒ���e���;�#�{��q9X��4	g$�zn��Gg����;�`�u�-��e(�G�wn��_�,�;�QP��w�nG�b��nW8 ���G!|hrM��, {��b��Ǚ�a�̕%�rm2�T�n�-�L�
�88��]2Ƹ�L���D,c�᧻A\�pgz�w�+*pWX�l��EsQu.�j�3��+�(�(�+�[/���ۂ�&B�0�{R݆ �wR�.{h%�p�pε�,L*5�U)���+z���R�!��;K���P�=W V��'DԶ�M�]��E���8��H����w>w|�3�����ņ��n�.�rccP���6�vrX����,t���nsF�c�x����^�6S��e�s()A����f�8sA�k��%k��S�F���ԅ�t��M�}g 8����R%��ބF����p\�v7���:j�84�P�fG��D1�jM�a���7X��"Xb-��ȶ�;�Ԭ�p-$���=�:��Ȑ�ƌ�ڏNY2��A ��_u+{��f�����S�x�$�����]���*X��P,z�e�X�n��)��ͬB"�{��m�F�et���dS+�c�mO�]u.�g5[��k��Cw1�`(�eCcs�5���� K�	N[\lZ׸ֱƴ���X���j` f�Mپ�z�.�5��mc����e��U/����4"8ʹ�[;dfv�fw\1Aϒ��L��
�*wwY��5G��1�E���]�ёU�W,ӇG6+7e֮���yh"�It���i�����Ԋv�Lf�f�a�����P)^wC��J��4n�g���=0� ����3�ሤG�L�k.I$�C�9$�G17ң��N�J�%\��ײ)$�I$E$�I$�I|A�O�6�&f&bgj*b%E^�����Q�E� ��*
*���FEQ*�+�t���ESm�FE����UDb)DA�b�(�T��Tb�(�"�Q�2V"�Q��ՙ�V

�H�"".�QF ��h��"��(��X�]�UAF"��-�ܙ��c:j,E�ʞP�"��q���%UUUAQ�6�9��
�Ub(���(��F�F��er�Q������`�X��S�11[h�TE�F�k
DW-\��R��ʕ��Z��U
�6ܻ�ʬD[e�UC-j�( �(*�p[ٍ��ͨ��E�ۨ_�y��$�E�DCq)~�^�-����΀]�R�nxa{cٕm�p}
4�W�k��z��nҍ�h�<�N���Vp���0[1f�Zr\�*$U�Y��z%N��ȼ��d�G�RM�#]��:�&��8L��vb�\o�;�w$�R�7�7�6:�sw�p(�[;���fF�{ ˾@��Y��8���!3j4��F�E+�篹5x��ם��S�����:x��f̻�Z~��;�VƓ�`�צ�^�c�30a��IsBʍs�V�7�+�bL����j�Z�,:c̵R8z\-�\r����J6v.��Xn�YrP��u7R���U��Ν[��	��[JwH
��n�Ô��vR@i�T�ٺ��+\�bj9?+���-����=8 ���z2��.4���=m����P!��7a�F	Q+�����@k���L�3}]�"��� ��s�����KZeY�e��z�0,VQE@5G���$i��7ou�z�ʵ�~��'A�.�뚰�L����3�Ψ=jI����r�Z�3�,Ȼ3���{Ԩ�)��"����R�&rk��wU��;'d%
_��H��k�k9C�R,��O%T[�<q�'=**+����;x��r�&`��SH<�{]x:��
IJC��OYU��C�ɋ\��hn�mC,�2��]�v,�}��i�$��һɪR��o]�f-�[&���	}d��}���ps�p Ee�BK�"=�v�5�|���+�u�D�X�6!a� ��;�;��i�|A�݌V�[��s<�t(ۇ��N+�ϴ����2���4M,,��Y��)��0����ރb��PZ& /9'�C����m��4�U䌸��ʲ�=z�=Y���l��ûN3B �p�R�6zE�l������7�k�Va��x ����O��w��=gF�k��'�2������&�`�5x$�Z�K4��%&[�O���Y��p�*u�������3�].++��MN��q�Vn "�f��ܖf�.���<uvЯi�_7e����\�������e=��Usq����ʎ>$�}_W�VH���$t�1����ksA��*����0"�mqn��4@�AJ0�$�|H��x�ߨfy�ֺx��|�����e�Qp�%CHƣh�$*L�e�d�+W�R�
2 ����
 ��|i
̛�p�k�80��*{�V�Z|���G}�T�i�{[��g.RG���*fH�B�ƈ��we����� �mPp\7��=�;o
�v{hE��.I�w���i�Q�xֲIupV߻M�G'�8h%�4���Ǔ�zq��
}��3h^`�]��XVz�%�e���ϲ�e-u�R�ଗ��]�/Z�٠��v]@WD�Jc���I1,�_'9�(J����*Uʛ��j)}��ݹ�m����p����f��[�\3uH3��LE����G*��-�D�Ol7/ V'�`�#����,^z7��I������"�j�M�W�$B5�m�N���lM����'2ߚv60����V&����j��x�ɺ���w䫵fE%e�ui@8Ӫ��r�s3I(�oM�\�i[X!T��sw�tsXn��u�tN������p��B$gBe"u�M���)������0�;�J���<��p�G��$��ptEX��7S��`�1(�U�Xظ�ۗe�NF�=��1��_gJ�L���H�${;a�q݌[�/n��Y�8�rK�9��9��C0q�x�����cM�ܟ�UXOo��]]�c��$qb��7�d��gp&�-��3�<#����5�#*f:�c�5�/br�)�f��z����4,<��pUC�F�{c�լ�>�b<rN�	��Z�}�pލW�Sp2��K�}2gC�)0W��̶��py�F1���3.UR`s]�˨���mE椚�殬��|����E�=�_�J)h<�u+V%�4!��\��
X.�Z��Ă���ēh�Y."�X���QP��n_�J�+�mj�O�'q b`	���Q�;7"��A\��"C��äީ����X9umZף��SP�>�*۫��^����7q҄�H�<�_z� !���l�����"�	������Fj2Zp���i2�\�f�?��ϖJ����š)�O�(T2Efn��p�]��!;[Va�Tj�1���}�-��w4���5��qQ��ƈ&/��;0��.	��F5F��h��u�]ك;��ꗜ��@�b����4�FN��=���*V����aŕb�������ک�ް�(a8;��!�.pV����Pc��W�4�cw��<9
i�x���Zh��#*Ct���S��C�f�S���8�U4V�k�!ڮ[��_��Bk.V�`��ۀ@o.=�@κ�5��[��4���Ggw []Q�sǰH�`ٳ��u`T�Dț���mQd1��Y����/�,�D���M+`�̏%O��}�Fi�E�]�A{xSJ�ҋ�p��壢��v��>kvnm�����X�Z�nC(փȼ�W�6�����2��J�iW�IF֢ZvyGn��(&bg��l��k�wF�T�D�1�T4Z�x�ẳ/��|��v�
YՄx�����P9�V/xΗM���a���M6CI+�a� q��}��i�t�jӘo�]�dx�K��7c7�^�"�ң�K���^����v��E���F�j��=BSV���W1�oV*�畒��h�{�m(/�!G��~}UU٨p-��������b�m��tX�}q��rqeZ������:��zy	6H���sgUN�ޭ���%�Y<�(+��gކ{�V����F���2@�sW�ݨ��A�N��p����f��Q�)�͙խ����x"H5뱌��m�]��^r|Po�VzI	�
�ˉ���9[�IOA ہ��ˠA:���z�ac�D:�O`��?~M�cq���k�#ɍ`6��վl5Qڳ"���q9�k9� }����V����N�G��t����A�Fl���x��M�U�iq�nL�F�8LĦ�Q���nR���0�Ӄ2���t�T6c�3c�/Ȉ�W^�zbJ?S�v؆v9Zr^0�Ҫ�x%�a`qC���59s���5,;ͮ�y��7l�/x:��2E���*��MV��ێsT5��T��FB�	(k��gxZ��u�O�G[�0ʽs=�%9�ҫ��O2;�s���*9�:�	r�>Xɏ������#@鼍|Ό�Q=����x��|��F�{�/�Y�5}$a�9��:�o2���Ӏs.�te:��l�9�[Uڹ�xy��'��6���,H�~ו���JR��Jv�m��M�""�*-n֧�GX��J���[A�ƍ�-��P�ei�+R�S5��`�p{I�B 9vR�n��n�2)�Sx�S�α>7\���)�Һ���8���B}���2�����Aǀ	��0M��k�֮��We��O�"�ņ�L{k[���N�%G�)��Ѣy�W-���326�Hݗ�o`���}�%!��PK}x�9&��-ɬI�lwe�@��벆�8n%Au�,c>��ʍ^���|��urVV�w^*��|M�n�(�9�5���p����˔)��;�\6Y�k���o9�ʻbIa�1hi��|�nޑ9��m��ۯ:��g^�V&�\,e_<��S�b�y��yҖ�+F���Vb���ʉ9Sy�)�w�ԏ���K�]�
.U��;�q��oq.��u��Aޜ�y�B%%s����^�b�s�d2I���vP�]��]���Χ/2�K�yf�n�b=,�������w��p���� �ٹ�Wu�G����b����V��D�d-7��O�Sr���\h�ϛ���u��7\�(#��*��Gq$�=Y� ǋ㳥��p�w���w�,iU ��b�a���f%/��;��@��d�Z���x֎��:�l�Y�g(�8:�\�%-�h�jZ�$q��E��(
��D����:�t�Ⱥ�T>^n�ݵ���j����8+E�E��7�G���b¹�)C�,�>��[���h��w�����|��rz1�u���.9��ZK��H�M�V�'-�S-��;	��׷p�����/6��u�P��n��nG�9rI$lǲ!���Q���u2�Ȝ�I$�99�s��9���9��(�-VĶVn�yh�kl<�0G.����bcb������a��^4c�K�m�
m��J�(��V�r��+TGL�(�)X�2,�]&�j����U�s,*S�EUEDE��[LʌEr�LՕA���kUEB�m�)DA��TDQ�n�[h�����F+���0c4�X��,\�b(����(�T������6"�Q���PQ����
+-��G�AQQƪ��Wkh��+�F���j��M�[�@K2:u%He�TT_s7��]�%��wbQ�Ĝ�����q%�0?���ף�� GN�h���,��X��ׂ�j݋�maE#ڏt7A.{Yl�Z�]�;@?YKx�u���mUหۈ�q���/��BJ��F:ẋ0#9Q��c+���h<_9=�y�
H9{��_��>�]�\���d΋�~j[���]k��Dʅ�RF�GL�����3���9{�u��^�{xh-��^ߦ���L�|`A$L�zA�8)�VB�lj�Ǡ�m���KΛ3�r^�pD
s: 3K��ꋷ�Z7(�J~���lD����{�E���(k���iљ��N�*%$,�I/ȏz�8���?6(Y�(Yס��k���Vp�%҇ڝ��!:vfE^"�h~��g3���ߤ����ydP�.
@�uq���}I�.7�B�s>at���45Dk�$���u�-%�N������}��A�}��U��ްfD��z@EƏ�Wy���U)��Ž��,�cr�x����u����KJ6�-�z������Hx:��vJ⩠uA���diY�з1yålq��8�L�ˏ���w�0��!%�N����8��7Rͩ
�C��iV�Z���f�V� �ס�f�Cn�F��\k��e%�2�ޙ���)�&
�x�jI�y-�xRr���I?_W�wII�����
nRӴ)�5���n�c���]1���U��5.��ީ���|K�\OS��#v"*��Ӯ�\�y׷9�|%_C�4��p(�[��3N�������<��q����Ü��#�ŗ�Ƹ����m���qA��J��xmZP�lV�O�MK5�t���P�i�s��+�c���>��N�նOtc7@�o�nN��rd���p�� �\2#)["�u�^Β��S���1��G=��W�NC�/.�n+�����{l�:p\v�[�b(\`�r�7-��}�t�^��ԗw�Փuӥ����Ӌ�)xU������Xʹ��5��Յ�q�e�G��䟕��x4 [��`Wu	!�U��'"��w��&e�N�V��B�q��c$@��qm��q!�k"�F�B�R�ǚv�b�w��$�:�����Z�q�$qL��^�}�FK�%xqx�MN����r��;�bcy���SVN���p	���qW5�Y���It��[�s��F�R�Q�fUX2.�9G5�sN�&,<.�%!%<z�!�DH5u��	&��s�Y�b�08����v��8.2oom՘ǻ�:�^߻��f������X�`�Lv�T�6Ty��әY��FED7w�"�;՚�օθ��p4�[7:�L���w٠���S�^����	F4�l�����V�t(�����z �Vk�L^��C-ffۆ����+{c���bxV��x�,��������M�^c.U�JQ�Y��/�Q��V��_k}�GM����"N����ZNy���4/��`j�;b��8�~V�����:�}�:"��c� iB8����Ջ}9q=����\Q�KUc&��$���W���^	��]<-3�\�b�U��������n�Va�k4]]h8�e�-�m�� uq��p��L4���ɝh��]6��v��^9̧�Ds�8�%���H���"�aM`�`�=��JT��7�L1v�HkFK{}���w-րj}�֘�͍I?_{ݙÁy�s�=�V�I��(��!�6"����v��F��é#L*5@ݡ^�
;�8r�E+��ҝnRy�f(A��Ac��tn�ju�"�Z�{*���V=�Ozxlsޖ*o�P�*�μ�6Bʷ��jk���d�D4�{�"��&W- �25Z�{�OێD�}�s�J�����Vx`�m3��F��s�a�L�'��mD�̎���	3���zj��FcL�xA��k8:�4�6m�^�j�}�hi,xv��E,�}90�ɻ��9�8��Q���I`�jF���a7O8�Ϛ�b�Ȃ�r|�9����J�K�K舊�N��V[9pZ9NL��V�*b�C�4�_G'�<;�%�-TV1YBދ����*�v�R�N�la�
l�Ib�h:B*��,��k5����U�M���fE �)T6��^r�Q�'�E�ۇ�S�n�ZRa޺V�Gls�����AQ(0�}�e��3/d394m����w})ʮ�7��ʱ{�tȘ��`B�#Kj�&�8X�%~Pud9Δ,!�ʳ�x{��>Y+>����*�[h����t���ţ�x@x/��]��a�e�9��0M!J�L�l��K��9(�y��A�N�..!X�ݳ%����:�ر�]��>�/�ǀqc/�Wh������� �Oڦ��O5i���l������{�&��J��tY�GA����ٺr	�G�7����[Rs�J��G"�l%�s�afn���z8
�Y���In+�*U3������o�e��x�=$���1�)�Mw�$q�{��z{���ݼ���q�v����b�eY�ҧu^��-�eoF)"�cë�yƠ��/*Og;㫃n�8&����F�΃�b�k:��ў��-y�u���L�آ�����Nߙ/����`��q&g<��|>e��CY:�m�D[��������øν0�݀��J ���"�"�_su�TV��zX�4-��Uٺ -����L�!J\��7����I��.���t��taT*	j�z�w�X ������w�:�Y�A��e�κ���Y�Q(��۷��w�5��{af��B]o�x1\ɗ� �s��Yi��r�_+a��7�oX�c�
@Yn+�LR���a��x�,�ʘ�tc�̷�� l6����VC,��:g�v���7��ug�V��,]�����'0�s�8RTG6 ��9������6�,���YG�E����A\�,]�ݫ{����&qu�qu�ٜȦ�'�;^4���G	�5��	�P�t�;Lvnƹ�[�%�x#�YZi�$�_�{�ݫ�|�=��*����+ڰ=U\
2zf8Ȉ)U�ks�n�xc1����t���]���p.��Z9�}Wq�Yq��%�u�]d&�n_��#�p��D������_�^�k��jTTB�M2��H�ٕv�{^�^"��<aW�,����P�9�2��B��M��M��w�3�ovTf� E�[0Ҹ�u��"�]�ב�C`�7V��w ӥ^�M�^qb�,�!���t������87��.�G�j�#�_~\B��](/{5fO�Mbܦ�z���(4U]��A_4H=�ra-�����TiZԡZ���uk�"����2�.ok����a]}&�D��4���5��5�ܮ]�����s��d��
]�[�f�ih��79�.��Gu�5��-Lx�]��N��Uq�q��bd��I��,V�\�'2�Pkm���y����͸i�6J�n�"mp�r˕�6F��;�pO�sI{'K;h�z��=�+�ARO�(�����-Yѷ׸!���Q��G�X�y�̣\��KB��sj�t�a����*�EPݚ���.�ww�R�e+G��a���ҫ���
(��meG��[�*3��K�VQ=��V!�PVm���w��dx�ޒHs6���+t���V�(*[w�C I>��h�
�sx9["�b�r���/X�j&��
�Ӣ�)Y�چ�gj4��Fm� U�:��2�����jFI,�;�<s�:����B��\ԣvO<��-
��f3Z��b�:�y�q�q�^o
�b�l�Z����"x�Ce��*����q^�Bf��
�Wl�`��cܤ]�t+������A��MS]R�
�F�8bPb���g�(#�-��+�F��d�ZV����r%5[}tȆP�að�|/1a)X���c�]c�r����{kCy��rU��J��3�u���'hIN�d�%�6��1�oZq�)�=�؈�"H�*c��/l��z0ɬl�S�&����m�e:i;��율H�77�L{kvN�����vQQ�L�:�ņ ����N�k�ɒ���oi�U�뻠W�K��S�ۮ�%�"���hh�H�G#nI$�َH��J�Rt���k\�6H�I$�I$�I$�	%�g�}3阘���EAeXEi̔uJ����0�
���X���)X�*V;��Z��i,G-Z���+��i��Tm*�S*²
�J�*���ȱ�Ɲ�Dq+�tٌ��[DVZUb,ī�m��+X�:h�1�V"�1Eګ�X1e`�bI^�V(*Ͳ֨��U����9aF�\C�A��(�%�۬.�ێv�T\B�j�V�;�GT�l�U`��EcuvST{�m\v���	�7��d�Yg�}p2�s�V��)E;j%�4p��}���i�^X(a!Q�+
���n{+�u=��3Py\v�eSw;N��k����m����^:d\p�n���҇^c���I�fP�zl�`5ebKv{��oǎ�R<H�U���h�ۥ�p�۲�5���E��6ժ+��oD�
�!�I��}��1� �IF(ht��-�j�P��ε{H,�U��I]�u�/L8�M��3��FX��ҖC.�@o3���X�T3Qäc�9yQ�.�S�[��p�=|��֧+���z�]�*
�
Mҹ�i�vQ�%��J��Z�d�Ʊ���T�bo|yF��<�OR�owu��Ƒ*9��'��iSg�M����ܫ�Ndb�E���������;|�I�@�1�p�8�U
��Z������  ��A��,�+�K��>�=L�c�-qh=��u�}mP;��#N��Ix�u��t슞=�5x��8OQ�����^�oM�
��v�}l�F�mj���'A%N�K�{Gr�9�sn�fS�����}�3 ;=�(���Q�S� �ץv ��i2]�Q�n0<���*���r�:u��s�Sν0)��%ӳ��+SКj�V����� �#���C�Ք_��Z��x�J�����I:4Ez���%���Y��G-N��Jr�����ؑ�,�f�����l�3#��E����D��=#��Mm���6v1��*��7���w]Ŵ�^p���w �]���s�)�8c�"U�#[v�N �����oo�3�y-e:����:.r
�$��	���]�$�M'.E�.��x�B�q�-H]�j+D�d�E4q����[�5�S�>�)2R����!�g^�ި�Y��O��[�1��#��Ef�`�\�qUb1������Zv#8�M����4mZ�5K^F�qՑv�d�e�V�%Gp���80�򽽃#��"�ub�w���o��o�6�҇���AA���M�5'^��x��z{�g��X����C�'�5Crk��r���5י���m��[a�nO�q:I}y�j��}à�ˀu�����g/��=��s��p�o,�d�@4r�n���J%���z>��j����\V�@g2�Ëe�7^�n0v8�"N�e 
(����H/=6���=5604�x;��J�V�VS�U��ZY�*Zvg�n���AQ�IS�@n�t#���q�����7"��m)7	+��zS��zO�������E閛AzT&Po.�����u�yd�9������9h���.tA 0<u`Ĺ�b�MЗ�I�.��eyn���'*E)��(��c�p�w����D@��y;x�ڔ�$��E/ȫ�����Ey�g��4iS�:���ùg1���d��ud9�"���j�:�o�XW�CueC�j�0��v0����u'`A:]�{؛w�ߘw�Z���.a��y�wV�pe����yϤj[ǁ{yj��ץrmΛw�2�N�]��3^<��^D�+Y�����#�aN�T̓�X4=�<��}�8���}^Գ%#��V�q��k5�{̲8��`��e��R9Ĥ�$�Q�2�7d-��o��^+���%m%%+(F��7�j{�EΦ~H�*µ�nfv�L+����AA�6^��$���]�*>ܵS�cN3:.6pwnC8���g�XoBێnHԐw%HǨbʿ^�}Z�Ӵy$�G\tj�5e$�N�u{��M�:��R
V�3p'M��uO���ڎ�D΅�і"�J]�ʹ�g7RM��Nwh}t���앀�r*Z����o��NO\7F�A�n悾F2Q$�fiK.����A�P�$�l뷈�1:�Ł&��a|2�B�"��ʛXA,�7/n���}��(1]�3�x �c�n�0�[8�#��]s��Wx�"Nv31�*�i���P���|��:~4��o�B-њ�齡y��w72�>+ 2	��%���ƽ�wb�Ь�ׂ-�6���)
��9�7���hXʗ���Soo[���+�J��ѼKv+�h�`�9|�̀z8r瀿銕�h�Gy�r�y������"m��gm�%GBYW���-�
��@���Y��w�N,E@�-��1��.S̣�T�у��}ϧ�Ө�V�������D�B)V1.-�Z�d4�Z�^*,9��לj�b�[@b_�����q��_RP+PX&�̬�i�J�{4qM�3#O�QyEE�n�HסA8�s��u��9�*�9���������m��T�FH��d.�AP�$ੵ�Tmʚ
��"tA��M�>�즩��3�a$�,�&'�q\��ܵ�3�5�f���A�kD�1��(R��*|��7$�O�a�I��7k���Ը�[�� ��AL�=<�ԛ�ͥ�*���{H�8�w�$q)P,b�h�VqZ�5�怹������AU=��dXW��5�^V�k�v��V��5Q��ve��M�9�z��i.\�S]�5,��f�;s�����4����{��5\*���s�6.������]�k7��o��X�.Y�UCg)p���q��[9��5����N�Y�%h����Xث�bN�sì�����
��0o� �1&T#��𗞿��/=��Mb�80�RNX.��l%p�4��pᵄl�W�F�
�#�#w�1 NaD�Y���_�3��^Qse@n�t#Ȇ�ooq���D�2�d��� ��p��񖧯/o���������V�h�Ѻ�iwj����5UQ��LÑy��[���!y����=�Ra���Gc@�l�l���Oڞ��NE�E��6(4c��u=�"���11�fQ�A���p-XUMA�fA�T!ސH��j�`g���Ȉ8.�8, ��M@��y����'��{��Tj{Ǡ{��P�o��t	+9���b�^��F��39{Vc��Z�F�ca=Qb6h��1OB�r���
^u��WP�K0��8�tਪ�_6�e�w�m�*�n�)� �w$�I'�K�8Sý�={�M�`���q���SN��v�����W�V���a"0�k;+�훡ٕ� ��g����a�)ĥ������ݱ��G^uX������+5�\V��a���z����/^Zw�� ر�y���N�^F��h楒���bF���wn����
m�]��UC�����)��{ݔ �P�Gz��CXC7�A���[|ң��[�W�й5�Ol3Y�"�_�=�zgrF�!S&B�6ۮ*��+�'�?���p��R�*������-?�`H?��`Rr$���#:�(a�Գ0�&yz5�OW���4-}�OS�@ğ�sbk7ٛ�X��tj	�
�G���)����f���ia��_�?ȟ�~� �@��D��>2�7�����?�?��~���}?�DL�6�B?af�<5��S��(w�d����JN�>[ܝ���8`}�P-K7�DU=�c�:dO����@)'rO�HI @�0I� ?���I,�w�v�� ����A�ʌ��)���L8�G�jy(Ď=�
����a����~���`����`v�����O������d@��1�/�������Xi�i��a%��)��`�&g!'��X����Y�a�e�i��k���$� d?����ڬ��(l?��\����0��7'��?�h��	$��Ht"���s���?PO���?C�O����d��1���Y�l?0��?I���̹_�1.<g�YwIŸ��de�a�"�!N��É03J���P�����.	�5�s�1�	)&�:�Ñ]�o"���O���x�'����;��Ò$���dc�����"��q�nM�O�������i~0 12~����	�Rp���SE�?Y��'�IC��'��'��ܓ���p :���X ��d���"�xO�/r,6Rl������6M.��u��(��M�{$�u,��	1��9;{4y2/x���$� r`I�����C��~�	$pG�����j�a>G�!��F9�	�8��=�sB`'.�ڹHc��A238���yBzЃ>��K��䗅��q`H?a�����~��I ����'�g�����I @�=�_�&��O����y�b����f�;�[-P/a�����ߣC$1���~"M��~��9�!�vsS9�����/�Xp1�#W[��
��xpp4�S@���R�qT����"a��55��I�H�
�m��Y�Q!�?��$����$��d�D�?Ttx��&��������h��p~�~��I���Ԥ�F���?~fΈ~0X�2��XC��?��;����"�(H#�� 