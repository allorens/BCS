BZh91AY&SY3�+� �<ߔRy����߰����  `a��BJTR���%� ��8�>�����SJ�0�� @'�<:����h��R{���Q�w%@(�� � �� � a�(7`@ 9 � �� �� 9 ;����� <��x �`���@�  P�  (�          ��ꪒ#h#&hтa�0#OM2�%����A�4� @��"��ɠ h  4���OHT�Cj�M  h   
� B2hM)�4FL�$�M=I����0�M�J��F��#b 2dd4�M:���c�X�OL�g�� ���a�D��s򩄒h$�wI$2&�ο�.+�I��H��t��'���7��j����k�Ng�tw��,�=���"hRtq	#E:Xь1�m��w� ���&�Iڔ�h�9�M�m��}�&,�ń�'*������z{���ᴚ���?��û��NW��������A҃�M��ٮ���m����#�GNB>��"s	����&��t��6%�2���'R=��G�9�݈�D���C�H�K'��x\V���J��7�c�-9���_��:��d�h%�:��q|_�������o�w�ӕ��6��:B:BA��CMg���7�{����dYNI�=3���ǲ���L��O�#�<Μf��eP�Jd#&� �$yU}���I�Ώbg�9�x�el��T:� ��$F�K�Dw�G#��<NzR'�O3��d<ĭP�O��$%D��&��#Q����l�B�lYҙ��X�w�JG�<�R9�(�ʏq�x�S���m{�'��drj��T1���M��:pj'��	�&����g
eoL��"lx<;֫���O�J�V��_+H��{�c�ˠ����I<{�D�I���)�N�]Kw),w��'sr��e"���8�{x}�{m��2Yq)����-����&d�����	�ZIdd]"9W6���]�<ӳGx;:9���WI����{-�Ky�����-�kd����m���}���ݜ�\;żo����{�c����Y�rS�ݶ�d��<_��˓��Y�a2C�2��2X��C���8Zaz����8�Գ�bu.��wǺ���F	tv�x7�߃~6�L�J7[��I��	�zX�B�͖Yl�nD�NȌ�L��/.V�X�Z�T�R�@d����QZ�jW���q�VԮ%%�"_�����g�K8�fޛ��)�[H�iw�^��w�=����M���*Yse57���o�Ek��d��\m�w��mq���,7�va��s$�IѨ�Ԥ۹H�#ك�+S"0�����y�+��Aަ�2Dw�Gq<�W9(��:{'���,�Y�gY=�5�]�3��6pj�Zc|�x�<o�7���6���zN�V��x�-ޝfI����<up�7�0'�i:M�dٴ!�j,�I�����l+W������ٽM����o�����7��fyi�wW-����B�0��}����T؛W_f��������7��m�z���Y�*���𓽈��JK��6�/�ѯ��3�V��2b��6aA�2�7����~V��n�j�#��J$f�}<s٣0���3ٗo@4vp�K:l×��TYU��/�j�:�;6QY��i�O�6R��_5��1�g�x���x�x�'����{�ݧ�^ܲM��{j鍄�Kj�n�u��"��5�n�z%n�4��D�IZ&�(p��;�����#�xY�9�Zs~L�YTj�x��#qH��k�Y�Ś(�4K=aҙ��2�m%0�CvY�FQ����^J��ΟU��(�|��)�h�lՎ�~1��X��y�$�]Q��kO�6�Z�Um +R{�Vt����UZ����&a����	�j�8v�bN]���xg����������}���u�W��.S܌�����6fFIG
<m���4���Ҙc��2g��׵�L��Y�͔Q��"���eڸ2C��t,���a�	�������]�J*�L�S�q�-'���Z�1��*�D���>V���f�y��޷z
D> j�sd5k{��/f���i�گ� ����[|����
u>L�K����W�T]�0�Žp�={�î�+Ì��/
x���7�KM�'!5u�m�B�M0|wwx��'�N�kЄC�%�����6o�?L�vb�ǹ�*=�a�I����QEI�Cv�Q7��a�d�f��!�t�Igd4�h��F^e�Z��%qZ��X\1�zK�"ŬZ�@�$�}�mי�ǜ��K�`*lV�z1cS|-�lAԲ��It�s�ܱ��O]����ߙ�5�R�K�3�����j��K��|�n�5=���
t�=��� rl7�@Yi���>�҅�Jr ������*:�lX$�kmeWW��>�2�:��V�EYh���\]D=�`�D"��/h�d*F<ۧ~�t�53VZ����ҙeU;a�}8�Ǆ]��<��\6)%Iݜ5v��NХ�,kmh�Ef��|����3����o�z�����Zi^�t�����u��Y�����y'���±g����p�V�];z��ݎ�s��j,�OU;8;ܽ�u׫C��������Ȯ�I��ӻ�㳩��k�E�wk����_��&��hN�U+Q�\n%��kN�kJ�=G�+V�8���T(%�f����k2Z��s�[�ʶe���j��\ˎ=(�4�CQ���u�hɅM=FڣЇ�5���8�xv*�QΉa$��(�5-�dG"� ����1��Gk'�M&Қ$���[�Ra.6&`�L<��Q��%g��M`��j;hR�B�Lَ�f�Ȅ�&�Pm+,GB�lN�h%?@�C����]�6G�+�UPVӪÄb6��\P�{M�EB�d[����Vkd�`�M Ԑ
e����H_�)����-�c�>4�X�I1'Tև) ������T��6���*$X��H���W�}:
�tY��koN\q�x)�w9H�ߪ�m��i׎ �D	˗5b��$��d����y�r���Ǔ�ޏf$�X�،Tb�8�}~^�O�����˕��UqU|��U(��[QUUR��@w�|�ԨT/������iU_,UUX�U+Uqb�������{�]=5z_q}��v�W�Ҫ�Ej�V�U򴪮���i���1Q��,-�J�lMlJ�w���Uګ�|�^��T�ڪ�V�W�a�MkR5&�Y�D0! )�BJD�(������U��]��X㻫Uv��Ux��$�!P�@�\�	�@��H��L�B�	DE+����t��[U^*�Zm�Ҫ�V�^���&&�)iĉ4Cm1�)pĮ�$
�1����*���U��n��UU�Ҫ����t��(NF�dH����� 6�^�UUTUW�ڭ��*���UWz�Ip.j�Q�U����ʱR�qLY-��K�5�\3�ؘؒ�ըZb�S�F8Ų:�+�����A!J���Ym�~�<�_�����g7���y0�&��>1e����`�!b:H�gKe���!Æ��	��&���Yӥ	�(H:V��\;4����!"a}r�*H�2�n[r�U�+L�q3P
�2��Q8'F���'S��43R��Vj�����u�/UHʦ;CTln2Q��@��%��V4�T�Pj�Ӻ���J�mB�en��*�R��M̱S1����*ƕ��̵���EmWD�n�*�i��Ȣ������� !b�+�βf����H8�#�)�Q����l��u���
��"bc��j*�-��U��NK4W,{�p���yu̸E*�٬2�B
�42R�Mu,�X'�v�̦�Ȥxע"��n-x�5 �Ӑ�UE�q6���U*�:B�%j��[����F�`�p�I5V7-+V�Zܨ,T}�X�<Lm+Z �}I�dyٕܒ�lu�9�e#��m�n�f�-r& o2RFkR)eVMYuV��[��]6J'5 �cDsQ�4Պʥ�j:��Uo6��W���؍��������	DF����	-����	%�����Q�����-����y�A�\8e��:�9���ƙ�/�6���>(NC�u�$̽b���Eޱ�+bG5ش]�-Aj*�����k*�$Mm@�x3��^XD�ջ!��W���#�������ջ��=����j��Q�mY�I�Ŧ8p�gyb�Řt��Ϝ2!�7>\�����Tyq�K�&#��w��0����CkѺ�r����oF,R���DAq�8"�Zo41�V��� ���a+���:qI�a�1�#���q4�)>_#EA#�(�4��$��~r<��_+_!�+�o��,�B5��w���ak~l|�ֺ���7�^:��Fl�>����]���r"�y���(�V���u��Jː�v��n�~�p��3�֪EgID�$�|R�Ŝ�ا��}jY.�k�0��0(�}��D	W��W-���:��V�ê�m���Tjɤѩ��t��!��>/BW�:֭8�,�NMS��Ϣ"����y�yEy]��G�3��u*P��|�!]�p����x�R��?w�����)5�ѧ��`Q�w�L�i�M�CEb�Jϑ����9U?A<��7�1R�q����ޢululZ��e��AAAV��3n&�bn�[xM�cm���n�,�w�Q�e�m�GM���HTwU#��������r���'�>L���%b��ks$��1��A�GN�XRD5�(��ڔ6������9Ƌ� /E摪���X&�Br�	���s�.�q�#I"�gHc4l�!1��������'G��iF#ѳ%�<O���I��x�G���l�?�c�4��5K���Ɠ�x��<x��H��04��A��G�����+������)2iب�_����>��%]8��&_���_$�Dkö4��J�m�f�#Ja�^]G��h�u2!~�ϐ���x a��~��$���H��)"�H����E$^��A ��YK`�ԭC]Y�n���Xr�e�fYd�ÉQ\ۺ�y�롓ۗ9l�qve40=C}Ґr�湙��#�y��L�ҷ��8À�TH��>8Q�'�����&b�,���DĻXa�m���of9��1ӕč�I��I���ŵe��t����b�0�H��@��T+M./@�L�҈0��AD�'��T'$ʰ�,��[75��mPb�E =J)�6���J��R���"�h��,�,��MZMe����M�g���q��9�'-1&��q5��2k5r��3������J��j,�BacFD+�Z�e�|AaE�!g��q@�CV���Ñf��V��;�[�o�����e��h�f�Mt���eq6i���߾�f*5b14��1�Z�s��G	R��
L0��((��m��J��9%�)/~{�&{t��O�*L�e�7l̘��u���JV�X�E:,�%�q���]&�ƒɅ��$�+G;qT�o1$�t��H�n�t�cȌR����O����~~hQ���.f"(B�����/3��X�[�fkU�X�)Kʓ��ъ>�]M	棖�4S0�,M�X@���EuJ&�
���m4jƃO|A�Qf}$-j�*�^�6�F�5���7V��.%�g>�{Az��ʦSɡQ��R�D
�����Y�ȱ�&��T�X鈾k��y?�,�� Q�� �b_a���Ϙ���ɫ6 {�e��F�Z�t�E�&�a�v�lh�h�t�&8��#jħF'G�ط��5!�aetJ\CV�l�!@x��j�6�j��,ٙ4���4Ò�5�8����QI�46),��
;�2%�
�w=�C�.*���CD& ��X�)��qR���wp�v�B�m��qC�b��)uJz���"�+'�BZуU��ȕWV�\�R
SG�0ӤQ��cbS?���%��}���`���4W�66���p������7�C���k����Dŋ���0o1�*4�8���I�:0�4@���Jb���1�/�ǡ��#�H��6|C�������4�e�sG:=>"�!�h��I�!�4a���4v=F������<|B���X�i:F���A��G#"Ǥâ�
��~��N���2�6 w+J3jG��.��2�t�r�b��8�+d�}Zq@���Bo��r���W��v�c�JN-�c����x�+����1���e�N\DGЪ��i�x�w\A�=�&�X6�����A��k�{X��Ț���jM�I���}�W���̬ȒK���\��$�(I%�C�IrP��\�<(P�0c�a��[��� ��)�ʊ���1��Q��A�^-7��{�;WU�Xq%AO�ܣ%+�Sz��+uBT�{�$nf��íi��"��s������%(:�"�a{(軠�kĵRE�z�����p�6c�*͜ӎM���z�~.!���v����ѣA\�a��F#����T�H�X�8J���V��ц!�����+�����#{��ij`q1X�8A�L3�$�Lq|��%� �U�ҵ�p����uZ!,M}�<PoY������B/Twp���@i��6>Z�VA�$��0��"�X�s��Z����z�<��a*��ߤ%}��1��2��T��Pi����-0�uqt��R���b �%�Y�$��N˂�H�7	a��CB[�~E�-Ғ�����>G�����4a���agWU"���H8p�K���R�C�C]]@�L:jY�l�d�	�m TT�i[�sOi7
'}��^����2��+�lq��}V�%mW��!
��(3McM��]0\F������<Ê��6��I�Ht8�le�5H��] �� ��d�t����U��Q�U�+1HE��B�uD�U�U柀��F"���Q^m��a���7@�-첸A�$�������bR�L�t��)B�-���P�}��1 q��F��P��w���ߓ��nL�aj�N(��ߏx�I,,��J���g�"���+[\d�5#)��������cjkKkˣ1XjagL	�V���i'Ĕ4>����gę<L0u6b��*��ƨ',�I���^Z��N��e����W�.�(�ϛtAӁ��nZ�.��A"b�����Q.�հ�z�>X�V$��I �Yck���[�قW�,O�q�d�$��E�yqv�)^���%t��ۓZ`d��K��y��n��(���0��t.��?�nG�H���C�g�:84 �=�x���~<|N�O��T=!�@�#��/M%�Y%�#K#FP�p=0�<0��'�>#�<i:F��a�u��ύ#�p� �4t:��~��zm���%��H��]V�j�7�8޾*���nM����k#�M��^e�ݬ�>�kP��YWy}��&o�n�eoN�7k��9��[���$p�$��$��$���$��$�<k33/�$�H,,�F�o�9312I2&�tb ��#�a)_���,=�.1�,�#�R��CTJ��nŪZ4j��FB�������0�'H$��)��ǥ���c�#ހ������dP`G���>�a lijC�qFz�=�VC
(U�8i$��Γ��9G2+���a�ށ쒅j0D���wv�:S3�duBk��R��ADj8���Td9f6���
��R��b���		]iy�����Y+�p>ҎA��32a˶�x���<�;���h�,��R��*F:��6��m�}Ο�!�M�v�\Pae�p�:t��""���G���x4�Ո���z4�>>F�	��.������a�R�bߗI�m��U#�Z�0� ��υ�p�(��f�0�%�/��
���B�H5�6�m�#�vd����G�����$�T�4e7M��F���0��'I����W��8-'dKwl�B�v�V�����$��*)գ��!R>^^Vt��=�Q���\�	)A?� ��Fv��)�pѸM���[~�J(�
г|m���]Sy�|#YL�n���'��oJ����/���4�-5D�%�����Qw�d|��jt_r��ү��J
�tM�(���]><|P�-�B"o�3�EMD����%52T_R�A��Cȵx�Y��GbbL���.�vO�:Z%2�""o�[��i�j�d���,��?���LS������@�6I3ܗ2^��S��w�+,�Aѩ���9N�Q失�b����:�%2|��H�J�t����R�I �����8��I�ҍ'G������4#F� ��<D?x�$��x�<:�I<0��F���᤭:x����?���h�x�_8=,�5X��TUX�A��}s�瑊�aU`�k]�NK���Y��>��S+U��~R�14h2J�1�F�XLj��r\d��4h�.���f�����V+1p}��շ%�C4�4����J��Yxh�A��%���ALQ�[H����%�	N���%1U����YeTekNi��ˬz���;���	cߨw���xD�I�I	�H�H�2I$�H�H� �X%���-��ג�5��%D�)����Y���E6�y�ʝ\���<�:�v�ݪ��-�62�k���!�,IjB�uU���ln�/��|Ҡڳyv��/���f�\'��'*��0%eC�_z���.SNE#rHAĵ����_\�=G�d����פCq8,.�,�<�:�~ll�Qj�����u`]����ö́./"+�Ը���A�J/���Q�<@��gO����0qb�&�(a,& �C�0Pe�cmb��V3�Z>1Y��2O�qb�8p�N�����_i�f!��s3w2��S#Q���cT�d�B���N�}s*�����q�0��u)�Eu��K�����A%*S��j#�k&0`j�s��ZpY㤟��#"|StX�]����\#�Y��M��9�ב���a�R�I�&N�%���!a����vS(�+��^fhB�ÿΥ��H�0u����k�#�iwm��C����]QwDe0l�^�tJ*F/#�	�¥yG{Ğ(]g�+�(��3���\\R6��n��a~m�b3ĔA��C|c��j�.3;4Q��O�:p�#�m#��ɢ~���6ϩ��%���.#ʏ���_��׏|I��gc�p�5#骙�n"���|���>S`:���֖(4��^�\��&�^�q���,��(%)�$k��P�_,2Q%�Xp����Œ�;��c$���nAJ��Nʚ3����
.��s���I:�j8q}��T�uypm���Q���
4�w��>>$�8�{bSb;wj�IvC4��JU��ڙ�;2T����������Iˬ�tkL�d-E��Fxvp�=1f])2�J�I��H�E��Z8R\����d���˕�i�N�w��X���tqY��)TQ�L���z�IK��E�q30b�)}h�ÒuQ>n�&�WA�0����rGI"�||?���~ �h�4�>#M:OM#F�h٤3H��$h���rX��Y:�x~(�����<>��Ğ:A��x~����4|<|O����B����]o��1��c�Λ�Ў-ف�5M�p�z-a�� �l�y��7Hۛav�Ƀ�O��s�������I$�I$�I$�I.J�K�333331`�,��������A*�f/�"<�0����/M\:���:�1�NQ�k��v̵��+��y��d)���	|Q'Z:Z���	'�,, ��Ȁ�'b'틵H���Ʒ�Z�x��J����H����)Y2���0YC��Q��(g���5��ER�[�Qb9q�U����,�:���뭶/X�fY���k��Um���'��m��,�D"L윱�1�p����:��t��і�R�3��}pʩ+ȓ�O�* ��'	(0/��3��0E,%ZS*�!�yx���t��T�R����0�o��g�����[#Tb)t�R��_N풼h�:|�_��V}��rb"f
������#���V�œe�D@�+z�!p�Äɰua�8��*\��Ŋ�1YF�'�iќ$�`x���O�D���|����(�����,0���R�1�����va��E�a���qb,8Q��Jl�=�X��p���;�gߜ�Luf,M�wlSwd�����E8���m�n�Kpj��!�髮�)E��#����������J1y���C��ϖiF�w����7b+��1�t��:|W� l����iܖ�p��:���̯�H�����_uBω>;����1���\8��j(���A|u�d����Q!8���(�\,e0,.۫�9"f�F�=qҶI^m��`�RQ�?"��ú�ޫq�:��v�Q~i���Y��G�UU���˳ iѝ,�Xu֞��a�i<Tu{���z&r���#:B�+P|��%�>8����k��0�!�}j�(���ϖ=yE��H��c>p���I��	��5�"ΚNMѳHf��ÓI(��P�,�L!iD>#��>��~8x��Hѝ���~�#GÇ�����IE�=���r���^��q����e�˻x�O�f[^s��U%��ۑ��S�*��&�V/�xn�����ty������i��1���á7���1���WF�^�!ex������|>�+����a!��*i�G�DǜzQµ�(�qJ�-�p��H���s{�$�I$�I$�I$�I$�I$RE$D@DXSr��>�wh/��Y��G�$�ӣϟ]�z�o �2�bYb�R�#^F�MV�-�Cy��fe*�Ȣ�5��r	�)�&Pz�vU^[�y[l@���f���2	��Wo(ں��� �i��U8�?>��k�}E�G�������D��GU�"P�+>GWV#ݟa��ψ�8�x�P�-pgĜ5q��PZՋx�x�{F��Q��Z�c1vTڤe�I�
W���"�1-��~h��1p�Ȉ>;���1�����c~z;�ϳ�31n�fE_S_Q�(����W:���RT�}A���eM�⾑�6�I&gQ~L��cF��*uI�#|�+��$�����>C�� ����E� �]�$�6���(�g�g��g�Xc�c����D�a��]�t�WҐxRoG/jS��(r�f;��"w�����^̒:�i�E�2�xW��~W�x|�q|���\D��](c\E)GOm���*5p��>)>$g
:R���CX�3��|�_xn��l����C"�;��������OLM{�Qn�\�$�gO�Qӡf�z��n2d� s<V��LR95j�L.�.�m���^<��*��9H�:���F���4��,�,��QJ!̸�r��S��' fk`�w9�F���⬔RF.�׾nD!�޷
�j�e���v�uW��D#�+uE��|A�ŋ<^�}ZרW��X�|��'��ۉ���z�)�K��'�om2[r�\�U����J�)��!w�G�kQ�ӧ�����s�uh�ղ�����r����ζ�+6���EĘY�H(�YA�A�^vK.
��1o�L���|��8Ru'�ZV�t�66|���ɯ�dF/1�+��k�|4�$�tDC�m�A�ΐ������HӇƕ����0rhF��C4�4�4�����#K#GC���t>���88��=��<t��4~<G����4#���Q�!h�er��T�k�>�W̆s&���[½;.�9�x6��3TW~��q"��T�ܗ٫���J�&^�יB���y2"�`#[��c�$�)"�I�I$�I$�I$�I(P� `0�)��s���K��ϫ\�/�P�b���-��up��!{���LF��OAg͓�w��#�1Yf�תn��6��3s(���B��I�����Nt�Ɔ��K�l����+WMY�T���3�K���aB���'Oa�,�D�He�n�
�8���/[:�.�
C{}���ъ�uyA��O��|0<|���V&��pd���a���$�H,�Y���N?3�8�<����d'�L>�C�Adv�JX4Q��̹���^C�uz/j�f���׍�e08RƝ�Q��%!- ��5��N.++��x31���*��w�R>V]���V/W,]m2@�w��D�)b���||gކy��Ń7���)e��/;SH�,> З�e��E.�|�F��,^ ������t��P�i�>99:EA�"$���]���DnHmnj�[�R\��l����53P]�GV.qY�ڼ�y�oȽ��Z)�a�Ȍm�1J�]G�;�7T�6ۊ&�C�Z��T��)ص��ȃ�ǈ4��(�7�@�gnN�D'KZ�X�R�C�+x������r��ܺ���յ�Ĭ���ajNv/b5><|x����4���ni���o#cz�#W�g�VZ]]5���p���i�pp�-ٙ՘���I]>9���Na�f��q��:�\�E�Ic\>D�Qf<���e�R��R|�|�E.#��g�7��>:,�9���rGđ�G���6�i�!���I'M��i�I��n�pd�f��#M"M"�""�pQ��Dh�4�#��`�?#���#���gM ���<=<F���=��[�$$���6�D��Ai���P��撯��lUT�"��;$�
"a*�u ��(*�^IԼ���~\�)Z�e�&šreT�_�S1�X�2�"�:+��C��)*�/8����EHF�ɶ��ݲ�%�dW�N���Ķ�+C���"%�@+�DJ�_��L�QT���j(�4H?��ϾʒK�I$�I$�I$�I$�I$�B�
0�Yꖰ�ȕ�e�)� ؅���{��'4,�׊�5O�GpeT�/(�Y�[����b�]b���K��e2�Ҡ�ƍf��`TP��'�)\�Ȝ�V5c�����ؚ��]��v纴1�$�8̭7�m:���b���rj�:p��H�u�Ĭ�/�JT�\+K�Cq��)��uI�� ������N:lv��h�X���#)RQ�ln%QΦ�J$��b>\Aֺ7|�&Bi�.�Z�t����)�2OQ������8RɁ�j��&x�=�T7��(�1}ῌ>=�Iū�{�Qxo�l~��I�ĢY�Ae���ńD��X���n�<&c�96�|�}.�l٫�T��a.�F{��:���B�܉�A+��IE�t�Y��O_�r�<��*�Lzf��ǀ�H�/&�n�9�])��U��d� .�p��&���S21�{�yF@ϔ�U���p���Ȏ�c~V��k���Ӈ� Ág����Kk玝�~����
):�j(�ˊ_uC�VO��)��_�&�g��'B�R����j)O�,�ä|e�q1��(�%�>�<mٯ�5D���#��TĶ,G|�-#�`�PΧf��I���N����H8t,��ϟ��O��QW�*�q;�t����d�G�X�D�}�Q�Å(m��mG�˞XUf
x��G��ڈ�L�Н69��]�O���Q(&�/ ��y��QwV����G�+W��k*��V�+�o�X�Q�̳Qꮋo����*G��Iiۏ�|Q'�:ϡ�����D
i+k����)�%�^���C�Px��h�P|�P�׆6�MN)\E�p��,c0�b��Ӥ�"`�,� �g�d�$�Βt�(�Ξ0ӆ�i�O�:t馚t��,� ���{ɻ��]�b�ZVu��f�3�vVE�����)�ұ�m��I� �I3�<�O&������uVM�3��t��$�I$����I$�I$�I$��L�	((�Z�rt�qA�G#V�6�i�氘���5���O�o�>C�;m��|a���%F�n�Q�K
5{ͭ��
N�`]���/���!je
�2a�Ī�QK勇�OdW������VY�Ĝ
9DD��Rv�@/v���L���#�c�O�'��r��DD�6�Qs����)jQyҺX�v;3v�ߙ��T*>~T��t��!a��R�G�ժu��DLx����1[0Ӧt(�F��\7,ɡ�P�����#.{-��J�G<�{�`�)F���m�C��7�Vb򿕯J*I�ե0���"�gf_gm�y34����SWT2(�P�፮�W���-Z�a����\�zq<�]y���Y^}�>"	 ���7$h� ��d<Gʎ}�s���^KN�i��p���9+��T���>��R9Px
CXAg�4(�{��ʙe���~�tU�pʦ�*`�;���2f*f_��j:iŤ�q���Q*��F#�6ƚ5U-�&#�D#U��o[mu��!�:����p^$�	4(���p�K>�VZ�R��䖈�ָ.��k,M�լ-GW�Ğ�ɱ�����I�Ӥ�*�x�oІa�=]���j
��*�R����q�b���S�j�>���ǜ��c���Co�=�U+_,Z�Guyb��I(�'�Jj>o��=-2N.�}�����Q�G�WNx�t5F���#�rg��sz���:No+����{����$���ԯaR�R�m��h�� ��W���k�䏱9���,���_j2�F�1�c-�3d��A��Hxԑ5�cT����M�3*k�2�X�)��-%�[�-�)Γ���`�JX��JX��)B�IK��Ē�B�
X)b)IK
X������K
XR�*R�*Rȡd��JJXR���K
T�E,���P�B�)R)`��������IJ��JY
X�X)B�%,�7�Ē�B�
TR��B�IJE*)P�)0JT���)`�E))IK!J�& ���IK�R�T��K)dS
L
P����,���)bR��0bL2�������lm66�����k�ic��$��)d��ڰTR�,)R�%��L)R�E,)R�R�"�
L6��1),��8&e(�ZU�*�U�Ifpf�2���,X��bP���3L�3�K,�1(�ZU%�L)1��,�QH�cD @� B%�)eK),����Qb���Q,QT��Q,R�"�e"�(��UR,QeT*�R�X�UYUE�E�T�d��m�Vӌ�L��,U�j(�H��KU,R,T��K%�v�`��V*�(��*VT����%Qb�*U�,�e"�,�K�Ŵ,�R��(�k��X�eX�X��*���KX�YE��*YE�eB�,�jE�-"�h�IQL�1m%�E%�IRRX���%%IIbRP���Iab��щ&!K	J��"�%,��Jf�ȱ����%*�JQJ�!��͘��)RR�,��,�XRR�QRqcx,�N�eÜ����m��s	0��!�:f?rv���@X�$U�mY:�ŇV#����=�N[�t���q�~��zz]߿<����������m�ţڔ���Vua��h`]�?�_�u��XW��i��_�uɦ]F��Zsj�a����^�ݤ������l�Mf������經�����
��;�oY�g����W/�G��On����HH��)�2ĂC󑂖U���)��������4�x2z����<�c�2GkI>�����S��3���k�ܳ���;��1����D�B�$����{��=�US�ͼ�Gܲ2�o��8R4I���i��B�e�Tg��G����b3:�Yo���}�m�4ӓ^q+'�O3�Ѿ;���2kV���*��S���n��؍&�7�s��"�ڱ~ZI$2F�H��H��1L���Fw�&D���4����C%TI,�"-I3dHŇ���my6�ݥE�32�3�s���F2bd����F��h2��[3O�zi�u�aв�e$��Q!iT���BZU!-,��&)!ȑe��}�CW�<��S��O&��Ok�Di1>�iϙ�n�c쳪v*��m�C�4��K�:5i?B>_��a�lxx�%:a,���z��+va�&�Cg�7�jJ����d<?l�orpuø��V8�����Osxx��9o�6<!�{�f%?{�����'��1�؞���u{��\�[��=� ���w��K!Iz'���|�}�SOs���w$�E~/��#1�ܝ�b"D�V^q ��O�qI̿�T���.s#ɓTs})�ؚI9p�ì���(����Rl�̉"M��'�N�*��*u&���c��J�����a�I"C	
h2|8	�&�F�	����)�\ژ����ш`y�M�l���Γ�&V3L��9��m4aJ����$~&���L��ˤŵ�^繣�u����zbA!�y|��)>�I)�;�RO{��m��5����:����A�u��f=Ȏ�þ<Za-yz�ܞ���O3�9��c��NȰ4��,v:�O�7Oڞ�t���X��|�igk���I��W�0�$����#�S�	A���=K�e��������:�X���?I�}G�<'�����ѷqQ[�U>��I����Z�2ʓEL��v'��z���ڧx�X��{�M���;��d�Н�����o���>�#t��6OB�׷go���9ĂB��z��I�m�f#��ϋUzڝ�I������59���NQ�'(�i爝Ե���l�95F�FTq�������y:D��s�<�BD�%�}S3�2<�ß����O��䜣�d���BD���5�%:�~x�g�}��$��F��>l���g����0&b��rĞ��rGg�������H�
v��