BZh91AY&SY�46?�/_�`q���#� ?���bP���  *���P �R�+�T���V�[J�4����V̪�V���l�m����	TPV�($ 5� %��R��Ͷ*�$4}�;m�l�V�T��#--�a4b�%��	�-a�-�+!���[b3�B�5���Ē�45RkV��fɪ�amE �Y`'��Q[�z���4KM�ͫMZ�F��i#[F�a��ƚcc!���A���6Z��Hd�d٫A,m�35����ƌJ�+e�ٓ@dD��u�ڒT�M�2x   �O��x���P!�v�Օ���.l��D���4n��Z�i#�ӵ�u��J*�N�����M�fصڵ�mN���V��  ,����er���s��x)JS��S����$�Au��F��n�A@���p
���(v��^��r==�[l$�Q��m�0�K68   s��{"R�Kh��A�(Y��T%�O]��hU�+���
���K/<�t
 O<���m���%
��^��@Oz��ʂ�{�i���el�XZ��V�*^   {A������<���+�'�}�/�L��zRT>�X��J^�����|+�����f(5�\��@
R�����A^�f��|�P^�6�*ё�Ō1A��   uܼ���ޫ�z
P��ÝԨ�z�ý�M�ӗ�z==;�Ad�u@iE�^�WZ�=ӵ��V���y�%�Pg�y����Ɲ��Q�[`%�V�T�f��  6o���{^���(+���ABT�u���ܫt U�uqʩm�K�{p�Js�r�*��׼zU;1@�^�U+�Q��%Y4�L�[m��ZSjj�   ݞ�`
�p��m���8T%	�W� ����x*���EMή 
jw��@�w����\� t[��cj�[QR��U�d<   �h�N����� kE�` 9X 47:ۀG]� ���2�:
v�\ ;�ٶ¥%Ph�Yij�i�'�  ;���wc� r\  ��pQ�s�p�;I�jXh 79� 
uݭ ��� tw]�h6�kd%f���H�&%�  ���ָ�f�  ��8 `���g@��uw (��  [�wU� N�P�� P  L�)T� `i�T���%Abha �2��IIT��  �� �O��%RP      )Hiꌑ�2M'����� ��2�M$&�%P` hi������������6��}�������m���{s�v��ߖ�9��r>B���yZ+�!C�����|��w�IJ���SԢR��{��H�^O3z���[�/�7�w#��/�ffmJ)WK-YۈJU��������l��c�Ż+�����$�сѓ�'DD�0d���'FN�:2t@��0蒌:2tIѓ�'D�:0�ã'D�tI��'D�:0��:0:2td���N�tB���'FN�td�`tIх�'FN�td����'D�`�d��ѓ��''FD�����t@聱'FN��:2t@�: `��FN�: td�Ât@聂N�:$:0НtIѓN��td��ѓ�FN�0`td����D�FD�	�!D���FD��tC��(��'D�:2taѓ�N�#�'FN�td��ѓ�D�:2td��Ht@���c'FN�:0Н:2t@�ɱ��'D��:&ĝ�: td�ΈN��FN�F�����ɂr`�L�rePt`ф�ф���ѐ�P�$4ʗL�i�e�C�%e#L�i��$� tI!�ta ���i��1#L�i�F���:$�:2@:!�	ђi��2�L��i� ta ��Iѐ�FN� td �D Q� �Zb�L��%Ze-�&�P� pd2���  tB@����$:0�Q�D :2 td�td t@��D :$��'D�tItI$�i�02��Pi��2��+�%ZeQ�i��2 l`ф�� :2:$ �C��!� $2���
��eKL�: �!'D@��Di��0F�P�i��d@:$"$���D�N�CL��i��1CL�i��*Zb��$�
4�F�$�
��U�J��-��eKL�i��1�#L!͉Zb�LJ�i��1�I�%i�i�\X�*�*�1U�i�a0V��*�bV�!�*��2#L��
�ʆ�����!��D�:2td蓢N���:$�чD�82td��:2Q'Gc��:2hd�����'D��pz2td�'FN�:2td���'D�:$N��:0��ѓ�'FN�:2tI�&D�td蓣�'D�:2td��bta�'FtIѓ�:0�����:4a�'F:$��ч�N�:2ta�'FN�:$��`�:$蓢N��td���'FN�(Ό: tIсѓ�'�D�D�:X:2t`tI����'FL��:2t@����x0蒌��';���O����S��EN�U8��Wa�9O���t�˱`�O�YTQ�v�s�iMԴ�&&�����EH2.�3r4;&�����$O�gu�{���u��G5_����5N�Cf�1[4�鐿�Dm��yQ��~L���ڟ��<1��gb	%�����a�eЕNb�bhq����[p!R���ٸ�a���6%�P��և��&M؃/F��Q\+ۏ��0��w5
e�0L+S$wY���;����U;��G�2�k�����ś���b�>8��`Y L���(��tH/��X����5nr{�x�B9�c�p�`���@�-��в���\�U�Q�"��)�?���L��XHɻ(�Z���Xj9a�&��p��p���	���%l��P�ĩK����	�v��}�"��1y�AzyPwl�����ȉ�BHr��ٳr��"
���vpćVѽ<��]�IJx����7gn�ųj<�;�GC���]D�
8;�=ݜ�R!%�c1��5���p�,hd;!�5*�Y�5��ĩ���Z�3@���Y���)�W��V5sx4,ZAxuU���6٭Q�Ym�uY?FNE�7s^��u��]�1exfDi9kV,g����2l�[���*=tv�HXz�e��l�;��n��؎�Lg,=�z��L< ���;	<xf7�g�K	-XvC�G0�o��XS������1 �]�.�=��_1�#ßﱪYV��ʪ�_m����PT�0���R��5K��Wg��{A����x�.��v�W{�Vm�M.l���q%0�X�/E�h��=������I|LE.	K(��_41�fF�6�O��yE0��r��դUu��v�gn`�iՌ��v���n�IM�ׁ�r��t�ϖƇ��[9�y�0�P��]���+���y���X7_m镠�-'��c�W��]��6�X��vHD�gp��᝚���/_=�orу��Йlr%&�oKr:��4�x|Σ�ں�r�S����ge^�j��whsZ��V�I<�K^���+�{�]���� �xuޜ���!�h�8�`q	})�(Mμ�׺�s�X�̻����l�F١��9��n�n�g6	\�(@ 5�eδjrK���#ӹც����;%0�maq��;�%�h�������:O�t�7 ���� �?��饮o�ނ�k3�n�8�y�y2�����[�d��n�MA�LAk�c0h���7���v���@�0��31L������4n�xu�vZ��ԥ���(aă��UGal��Ir(��r�ئ������'��6�[��;e� [�R�B�����8u�Fh=�p���tH.\��f���v�\S���B����>w��d�4tTc=�z�kįMu��S9{<y-i�P�-�6�������x�L��fYV��j�n���{:Y*E�:1����_|�1��y��N8�9d�Q�p��׿�
;iB�j�e�CF�Z��N�u���8ٕ�X�S�w!7uS�O����O!7KCwgs��6Q���(EOa�^S�6��X�oE�Q�Vۭ%�wPA+SѢ��8˱�Y�Y��|���ǁD�cR@k.�Y[v���ӷб6�7��6v�*�-+64F�����{��3ܢ%�H�CZ��ײ�8�n��R�ֻ��ف�Ҝ\�t��z��]�3u�wq�b����]��%Z��M�|>wp}ɤ{�c%R�r�i����7	�xq�֙��i�8.������c/�C�v	� k�暞�8�M.oW��Ǧ�Q�H
��[|�εNu�"��-���R���x�(�O��]�v�b�zRy�F���N�O>��UbI��tWG*FuXC�;)�����vC���z��ڻ����[�\L<�TX����M�v�����(��p�G|Oa����kKu�|�;j�$��-�ǖ�=gbɼ���Bޏ���0�ĭ�hb�f5�]%a���=���N{�Au� ��7b���.d��{��޹ܲ�N�M�!�F���j=pd�5KV�:�ڹ��ð�X�W��mZW��T����yv���v2��Z����{��۵�� �{�sGR��3����i:5+p(�ۛ*ºXك�(Y;pڵF(�3�6�NBJvsq�IWQ�������X^�ǒ�l�iS����u4�S'��4/A���-�[͚ՎU�L]��ŃD���&�#a@�:���o۫��dwkx��O^�p���u��qZ��9tk.&BXr��^�X�^7�]U<E5Q3 ��3�ʮpKv눾!i��Sؒz��ҫ3K
���t��v O
ZkH��9Xz�}�9��[ư�t�apCU��K����5������й��UݽьP����J�ݼ�G��3�i��(�'#��a�9�X��ʵ�ő�Ճc�T��n�6Da�Yo��zUn� wY>c��c9�m��W�ꞵ�VhUb��!�nS�,<�j���n���n�n�K"u	��x�7n�p����2�X�����S9"Mޖ�Nu�����7�7�i���r�ڵ�x,������Ww^�sd�ќԦ:��s%����6�z,��hqt(>.�i��;�[K5e�u���0,�/M���d>$(��N�q1w��d���xX)�!�1*�`ݭ�pp��zՔxf,�_=.���W9�.�����M
Wьކգ��T٤���M���ݤ`}�����UGk�BS�N?L�t'篤��4�O�Q��s�,a|�ܸ��to\��`먀�#��v<ѽd��)���12�^�WiP<�>�no�6*�;��D(]�3�%\���I'D��U�mt�/��y��^+[�7�{�Nz���;�4lDr� OU�.�����f����/g�	�:>&�oi����A��l�z>rf����Xb���ۑ�+���i�pN�O|��Z��db,�3WQ9K���{��i�*��p�L�
+X�ƫ}�2�l�\�5�ej�cJf��B�C,­,;4�V���=�z��j2��ZKUwt0=!藑�q�.�OoY�8��}�p������L�P�o ~�7�]R�B�@�)s5i2s���o��'Hawi�c�6����y�eK--ȍ�b�X�)�D4�n������x�O��t��!A+�kG(&]����y��e�~yb^,,�Ie�"�nk*k �'J}7F���JuFT�������L������Q��~�XK�;��Ö�.:dP �k�S��§݋vǖ�lx��Иb�8\81a˗�	���q�R1=Q�r���3A���;ejw��7/`�6������oE�/���a������ņZ�Jq�|���ڼERn�T�S$V<cv�֖��]��Dfk�m�w�Gu�6�˕��i1L���x�6twjOI4�,U�w�|�uf�0n�Bͬn�#�0j�r^����+2�5��!&�ڶXA�.���X�}re-��ú"B.Ғ���wn�f�Ǖ����Q�u��[���v.P�;�/�X�Ӫ7 ����\�>�(e\.�1zj-Q��͋r�skC�}��Rط�
��B��p:H����l��_h*����2)�U����v��R����ksMݵ�Vj4�:Z�wQ�J��R`�0H�߷B����&��:c�k�:O�Z�Z�sFY�{�(�<AL-/� �%��~'�2�Ż�͚\݄Y�!�㫛�{X�Z����Wu��ӫٶ�z���ΠbbK�U�nL����� �|::�Rtn���6��X����ӷ�X�-d����fc��-�AW���r�-��M������8���u8ko_K�V@��A�;a�{��n�b��q��on�FM�+�Ž�u�P����®�-뻯���5�=h4�U{���ز�O� ��`d�2j ��i/~��)�.��7Q�c��>��G��ï���3wC�9B-�wQ��Z\�\�,pA<���l�o1�;֪�M��}�r�N�aS�V�E���W��Lq�ٖ�I�
�wU�l��4�:s�5����n��j����n��w����D�ё�N�`B8g[��n�Sp*^���:�̼���� �J�<՜�a�Յ��{�*�&M.�� ���qaG�T"�ԇ.�ea��,�;*|����H]&Ҭv�6���X�b�[�X���-�zk���5�0sd��SH�E"�롕%������&.A-�Bs��'��C�i�Ϧq�B�O೗#Mx�Dx�9k٢\ۡ�����x����YP�(|(2����bu�F����
˕����/4q+��B`��OxWl|�-��z�i���	)���_�jm��dLd��U�FD�'I�����(��c�a��%��0�fs6@�Y�����q��C��XI����.9	MQ�fr\������6�0��Yzl�s�M�{���j�58�N퓶���6C�LSΜ��]}n#��KV/ p_�^�sw_�;R]�Dd'-��i�2��&�[Dya�)f-u���l�M��m�uk.�0�Ne�ʭ��t2�+I�frr��%Ȣ�z7����R��M�sk/'*3����1�v��s9vl�E��DS�"����2�:�}bR��8kV�U�K�S�;���ɔ����-�qf�� 901���#��.Ep�� 8���l�x������1������;8�v���L������7�v��[gV�s�L
�����܈���"V�&��UȩΘ��2.�M�r����ڑV��$���i��D�-��.��Q�EC�f.с�r�Vb���Oۙ�M��sLҺ�Q:��1��ۆ�#fn��b��j,a�h��P��Y�2�\�3ٗg��Ѕ͗s�Kȓ�$�Vb��:�7���������Y'C')�y�CX��\�ui&���ԧ�l�n��i��x��� �H��fn��
H1����ڳU�%�P��6�S!"�/tQ1�~�l�n��GR:�\��H:$8��%�[r��ws(yN5���-<��!vLQ>|�l`_�`?A0�r��k�0�ќ�4
>�;#�u�0�ͽ�`��6X��R2u|�,Һ[�[ܺ@v�q<�.?�"��뷮�!N�6e��5JٱN��
R�`�_;���;�E�	uF(r䋤lF��`r[6(�i˭֙[kF	4���Ҽ����ZyV���(.P�Lp����o��Iv�Fs�;�GqfU�&���N�,�)�!�dXwP+�����Bfu}���i�!�������;:�6��R_��O��o(4efE���PhU8f��Á<5v>�gdy�Sg�|:�a�������F�V��%L4�F�<jdb����h
�Z;�?�]"|���È���&���k��s���k���^��S9Q�?f���f�i���^�m8% h�-�Z6�jn��O@kWc���{��{��q҄�ѬL`aת�]j�/B0��LmWjш����(]��$Sbs	�`Ӳ��%��<�,ݬ,٬t֠[�v�ˎ����يٍ������v� �M��;+�(ƳQ�N1�Z�m3���)�Q���XnP6�b�Ȧ�$�gV7V��w����ʆ?��<�V�鄱���N���M9,��S2����-�5wT �`q����V�)c�k?mƃ��MmR]�E�G�s&�L����w%h���;���l�7P�G�N#�Pi%͍��X��S�ŝ��)��yyB`�tzt�ĤǮ��ɶ[���4� 6Vԝ�y �9a�����y}l�=zKt�z���5��V��R �-��BV�Y��c]��H5��m�s�=���8U$�0V)�«�&��C�aT��۝;�S��2��lc7���咖h{���"Mꏲ��#��9�Vn���m�eA�t��&���/r�Ŏ��&��'��I����ESB���Q%���h�4p���5���7�)�W�ΪJ(��	�5,X-��$���9�(��`t���7��u�u��e��n�ɽ:��UHƍ�hmm�L1�z�ha�8M�*u�[�l�B-�y�ِs��0�;�����&.�%6%Y���b�����N��2)Ӣ#ׂ�7$5��r#}ںW�\����4q�\�V�x�*v*��9�a��])��N��YZ����4�ᘃ�a��� �j�ڻ��Ԫ��uTb7�zi�<�t��^b��ۡ:^s����7�^c ���x�l����S��^<T��>�Ã`��>b>���}�,�ٸ�W��#wZ�sJ^�C:uś�0������
��.��0p��c|	L�.�Jz(�ԧ� �!�Q��Q��@#ýź���ŉ��[��V��ƨ��Eө`�N���A�${'G��5���ʱ�{��V��B�u���<�?�)v9k0�����F\\6C����{"77��!�3���w�E�۽�8q��h�N1����41�糖�0�^�����\1}Ç�EWF2L�hZiEk�(�OA����߮��
9�V�ThA�4o̈%��.��G ⸑%Z�g�Ǒ�':�ޕ�V��]��"I�$�i=����{��(�V���r�,b渺n�5�eä��]�MĒY�L�TWe����v�0��}��n{�_�~U�f/�Ugc�9��u�qS��V��_�v�%��x�~-�N9�<|��}��Ц:e�[wo�.�Yȧ׬�l_L��(��l.��A�-��t��a�Ⱦ�c���`7?����sVjS��)���}@uo�	d>��9f�{���a�F��v�=�;j�E�e�Ը�P@��Ҕn�!wV�����z�3�%�,*�W�����3y�q�Q��
zx��T�^2"\�}y���V |�	��O"���G<g]m_1�Ҝz
ܧ��_wV7����hF���(Y�n��g6!��Ê݉�*����g����=9��2�4qy���d�ڑ���/Op��G,[���'I��0��,MҦ9���	l�9Ye1��s�����n�e�������8�܍��XOoN't)�m���5U���U&�+��J}�z����$d�G33;M�� ���v+�k�����sǊx7���8hi���]�ѡ��mJy[MF�v�d�\��Ya�u�9����F���O��W�Bz�R�
8ǳ�>�=���������o?Dh��0c�jT��Tv��[]�6�����{��26��c)E�1��2�T�^�4����J��/G�^���8{kB�%"�K�jh.]�ٶ�,f�Zpf�|z�Z�=���}��l�a�!�ķ���hc��spl�ݣ���fwN\��ۢ7-.:�P@��n�ǔ@��v�Ohͺ��Q��z�Òe�<��6���<%��>�yI�^��KYj�E���r\w[�q�,��\����R1���]����Cf�:��z�Ɇ�VF��"r�^����/��/[�����H�b։�G�Q��s��<��}�(��p��5%���&��2]�e����q�
�}Þ~�"#���9�1�\/�� w��zd�+&ǁY�,K�
��jc35���F6o7��6�z]�5�9�E劮Ц����f	��K����b���fo� B���Y�s��(J�<����LA�P���g*S{R�j�Yl��ynI�:�'�W�rgl���tS�.I��o��{���wx����,:���{Q	���y���L ոU�a��k�T�/��|�{x�9�맽w�m�����*g���r�?z�ߎ���ˈ�6�7���`h"��;g1"��=rw/%���v����ܡ2��۷r,��q�j�����:' ��j�2�1�86��-CT�gv�#Y͑�4�T�Q�,�}���N��$,[�ŬCq��9�>��=��,^�B��%��V�0{fV��wSd�R�}ڎ'��ᚣ
_h��uxP�1\��ZR����-&�dٖ�κv���e��I����xK�MoL�p�v@�O�8���1�AO#��}��&�a�<�F�!� �m�9m;&�uq�����C"�	)�f��W���R.Q��6Oj�tѽ�EWE���$c�8key��8yG|H���R>F
Z���ۋ�����Q�SPmr:T}F�";�)�� l�l�U-��.d��٦����ڄ]|��󣮒[)z%�J�5=�d�mt���p��ǉx��'�c�j�:V�v,Q���>J�݅�z�+��y��I7��]���3`b��w��>oڟ�X��}�0�9݆�YEP����%�I?y���]��M����aI���]vd��MA6��wϱ��y��Q��{4���I��.uA��1z��nþ�w�ƹ/{���T��SǊ��aô���f�����{I]{�[2t��LR{G��;)�,��.�V�x��o��6�-�8.�WQ��@�׋�e��s��X7��'P_=���k9�i�~��w��#V'crxj���\&��N��z
�k�|1�U��x�� �u~V�`�1�}<\�O}�x井ԛ{��#_ݎ���5{u�J1�,�r��N9'A�=)�]�|��j�s����1���WC��vz���/`��);�G]3�;�j�b[�W���g@ͣ�tc�n�m�]���awcq�>gy�,���t���bw�|,��f=y�ͱ�UB�ƥn)bt7���/��8*�3��e?�8�)X�j��y5ą��5�auA������;&]L	��j�����t�����J�yr�~���Uu�,�, �ˠ�o_
�KX�I}[]�}A��Y���j���P�zƅ�ֹ(�F�Wnp�Jr���9��A���Y���>.{��J�l0���y7�s�١.�sa�׵?c���rN�Q��C�ĴN��xX{#�3_A����݇5Wq�t��5��Z�Ll��.��;ʚ�
>��K8���V�Dwl蹅5I4Pݕ�o]�uC�rH&ó�"��j�z;�'��9����� ���g���	̔,7Sq�����g��s�����1DW{�j�.�MK^��S
A\�������E*����S|=7&�,eĈ�OX��Wr!#��3��̇/K�$O�h�V�N���7�׶��G/y�̺��<o���Yq�𕦁Oey���7[��a}l�ç�;}w���;,��f�ȟ^��඼�f%6w��ţ��f�<��z�i�:-{ۥى$���
ϮFy�L�`��&�{�9;�r1vsGƴ�.O�V�;d��,g.�a2d��C�FN%��C���yC!�j�0�-����A�o��{x4d�<�����$-`�ط\�1�v�b�z��/�=�����~&ǚ�(������0pךBR�r�^���'�5���[5a=�Z�i��/c����S;/M"�c��S�'�6ڈ�{�Y��۞�>(7M+Sr;�faP3S�e�z��Mi��H]iޑ��=9i���2d��z#��m����
o�1�h���L�^�7u��ݳS�b�:��,�:�ի<K�V�nv��^OD�s�>��+��Ǻy���G�ѱ�/��8�q������K�6�7�������=�?��>�H�3�
�+ֺ,�3ϳ/~ὶ'،�؝�j-'}������n�u�hέ��C��ַú���}���]� >aof��`fW��ݙ4�"!@�o[e�N�&C�W�J�� ���D0((��{��S�^��Y��/XA��x<��M��n���I���y|#�{�������7Dښ%QG�YY��)�s*K�u�JsP��ܫ2�ºh3�R:��HZ<�Ì`<Fy�빵�j�'+Pڼb�)�\ot�l���f��]��Bŉ���s�);�`�xyy��F�o��=���;�S����}OM���Q�w@�]�N�qp{4o�p��y;���5nrU�ב��qm�	�mf�ré�>�܄׳?���{�z��q]y��5Tu�V��f#m��ͥϰN�q<P�v08M��<ܘ��-#Ӈ���E���U���a7����>�N�|������!=�Y�^|w~.������ǀ,Շ�z:7�~���x�WT�F��PP�����x��{#c=�t�� J�w20���G�nQ}Ȣ���Cfȕ�pn��=�9�nB����[�ɋ+�g.[Ϝޠ�wi�g9�'
-�b��C�Q\�6���	U�d{���]�F��}]���� ����⚬�A�7�S�~*&�����(owp�y��,��k{|B��U!LK�|+���/�w�<���Z�ѼԅG�g|�Ŝ������o,A�wim*-�5�V�n�C9r�3;�[�"�7tғ6�yk��r{Z��ɂ���w���������.k�\WZ�ڧ|�j�WpQE{>���D���׮u�+�vy]$+���{M��ɥ݆�eH��Uu�܏\5�˗���&���v����=���&���jG��
�8�I���>β\���=�3؛k�<��G{�;w7�Sˇ>@�_��n�&�ױ���K�B��9<��]�}�{�F6�;s�:�n=o�P�$Qj����:"�b�b���Ru�WP��ܰc��-�~�}ѼK�k���	�^��h�������\�3���XM½�}6if����V�bK�&q�h���dr�u^��][�i�,n␪e�y�n�b�_����l�
YydK���6[T�LAV�ַ'*�;�_'u;�}�/w���wA���2f��T᫥���n���f�k��E"/�����vL����ʡ^Y��yV��XV����cL�p�����Ga+�.�_`��03���-����|�Z]U��>��}��}믚Hx�{7lN��=ǡ����mC�#P���;��z:;�
�f��[�y��]��xݷퟯ�;�y��
���w��;e�:���1���ˎ�7�|��=��"u�<{G:��Iڨ������f<��F<𤙾���H3�|\ȷ�;+x�n�K�z�6��	��ꐆ�E�j�rl"�^�����]OfG&֕�ls8�ñު<��t��W�(�G��c��p˲e�؁�`���1h��{	��ө��;_f����1K"oN���^�Tv��;�;�b=�#w�I��5�1	�{��oG����G���;W�g�� ʰ�]>���"��X7^��xl�w��=y,�ԗ"ҷ_Z�Z]u]����,$9���g�nnqBW`��Z׳��xr4'Dl�sBJ�S�)���c�kӻ$b�}�x<�py������F.H;�5�"�Ջ�k�'���&grc[�!��9+'w�q�$��Vs�H:nTc\�v#���
�ni�'Z�	MJn�x�I(�m���Nޔ��F�+QvP0wCz���T���;y�p��,��4������m�7�gdj���c��ŭ&{}�<2Tڛ]����8�܃���,Wo8�!=��F4=���	g�<5_Np��N�{��-|6�a
����%�Ց�e��5N��c~�N��#���fJ��S�9���w(���_UA�c�S;i[�5�T�M��.����&=y~n7}u|�{��{������qn�ʌA؍���SbQɘ5��m;m���YWO ��m�=o��ʮ���/�ա�����Vr��R-�R[��2]��V�C׊Vr����i��ywv�����cu�褨���X`����O��-�|���U:��$����#�}�N����޵��}+6l��m�[��J�Y�HwS�w�q=WZ���2�NmѺS�5Z�đ�SIfZ�����v�D�w2Xq�~���~��=�������zć�V�Q�O0��/��*�X�i�]��4��'̣��7�p�	�%�?`��Ӎ�xR ���a���������~`߻G.���g��mPS����5��g�y�n_M�r�v�ùm�\�T�W*kg�l'}{,3%�b�n����^��{��KHO8jdd3;J�E�8m�]��؁�N���)Ẃ���\�ljաBv���(�!��"�<u�>p��2�왧�����˽|�ݶ �wAw�x:�G�:��a���H�u��̎ؕ��+��:��=��#���]Js����{�#&��q�9�)�u`�k�d��4P9O���<�1�w�Q��Mmv33�ݮ�#p��׻�)ؤg]����W2k�ʹ��Q5�Uֹb'��R��o��5߽0*��N��e�ýv�4�<����U�`��o�g�9�]QY�gq�Z$xL���	4'vʖ�3�D{{ �p�7_aӯWF2f&�ɸ��q�7���T5���hr��&�-h�wB+ㅧs�WCtU_Wq<�S�:�h>���q�̳9kKFE��c�m)9匪�V�c)��Xz�>�A�����2MӸx$4���md����ßA�]�w/��7�B�Жnc�72��*�����ozp����{�3i�*!(��!|﫮�鸦9as���u�6���9��/��W��ԧY�3lz ���_ty�
UMk�rf��(���"���k3xPG2���	���ѾB�$.K�úg@ǛYiZ���+�"���4x�R��11.��V�>/�o{[k;�s���MHz�2�����D�����	�~�#o2�µs��>Y�=8y*��b\^��'i~�}4v�T *,��HB�Od˥j��8p�{V0����鈻���a��K�WW�Ժ�G��|m�ű|M����M��)�f�wCx�|^޸����.�q�n��N����Qj�ɸ��&Z���h:f��Ȱ�v� d�hԇ�T�d3ĕ�0ֵQ��ۺ�����'��n�O�7��||6{ۊOM����QN]ˇp�X �����zF:�9�sm^ٻ|0J�ܝ%�!�IM�7%�ǖ�����\�2W^H���v9y�w�Z�jٗAGX-�ZY��!�RfI���S���i
1�rW ԅ$�ѹ2Lm�t��ݧ}}�t�J̓�V7M�껪]'{|=tN����&;|�R�l1ŬN����#���:9���:<�������Qp�^q����Ͷ�l<'��$����~#U�tn�H�	MNl˸����b7T�sI��֌��7�n�8��sC<�q˿oQyo��YI~���e��[WtI!�Ƣ�EF	3l�@�ĉ��	aͳ���ʬ�҈�F*��`�y,��v!�q%�b�N�vVQI�8��!���| V�L�V�Z��LzN�f���i��I����z��˚Ƙ�3Z��L�I��st�G	3_9�װ��hmn�G����*�T�.C��M�!�** ���!_��Ǫ��ʉCLH�g�@ے)B�����	t��`� ���N����������]�āq�B����C�d�Zh�M!&�@�D�} B�\�Ka�V�2�!&`i�$J,%�ZV�:f,����l?�}xb!� +L��S���_�I���
h��a��noOsFޕbs0���r�"����BP��w�����{�T�+o��|_��׷�u��ٙ�m����q����6ͻ���p}��٨d�K�=�ʠr����=�^��p���Pj8K�A�뵗��wp}TO�_��Ѣ+�k�
BM��2�؛X�U��v�sF�}�vb�G��7�UG�g:ux�)r�af��Q�$�(�H��^��_�cM�6���S�/�[��}9n�����6���*�F��E86�5t��yŔ�@�'Y��XC&����j勢,�qa�Ʊl�F��v�ń\Nq�F�в�{S^�غ�d�n�F+
��8W<m���fp=R���Xn>/�Wg{y����,r /5��$����<���<�����>��D,�;]q���9-D���b�g4V�X3������Z�lX׽�+��<�-�V�>��~;d�KV&"��T��L��M�.B�� �vS�<��]��f������$�r���l��JͻÙ!�!g��twʫ��,����w}�T�W��,3ؽ2i���b��ɹ�/���/�E0�)b�;�7���z�{ J�]�=���&�{�>�V�Cu�#�:��h]6L�:K�uV*s���D�3s�k�����=�×6��+��
k�4Ȝ�ڞ�Bv��:���y{�Hc������x�dvj�5���-UE��ܨ�{���2�B<X�apB ��AA ��� " � B " �AAAA�9.9�6�>�-�_Z0.�F�)�ϖ�(��f��:�db�@ꖦ�C|`ǹO�W�G��3%��u��6.氊�<��ﯲ�΋������o7�7;W;9�{/�+�ݓ�l]����	�6�[�B�!c��V���۶3/v�q���������Aw\��Խs���]3��w
���F�u��u�''i��{�^9���u��p�Kg�;#��e�Dу��Qd6�V�t�]ܳvyE�V���W�<fM?\�{�uB�f̪,شhk�lQP<)��VFm����|�nM}��g6/h���ypШ�u����Z�=+<���0u�B<r�ۚo�&��&�X+��>��<�$�]�[����[���.���;�n��{6�jn�����ؓ����N�;�9��$H�=*���a7�i><7��<%�T���T{h��Q�˖U/<��	j�v�E��{�d���M-�7�����%u^9�K��lsj��soE!��$'�|�o~Z%R�ICe"5du�|"˗,m��;~�q���2Jk��w4�|�&6#���_(���J6b�{o��^��-����:����3@'kw��zN.��T�:1�k�'i�k:e����~G7�y~L���Q�.:��|�c�a�6��l@�8@� � � � ��X � �,AA �AA� ��Ap�
���b�aoh|�ٞ�E�(���o��!���V��f����Je[�%�Xd��	ܹ��=�ȗIK;�*���:o2:kEV���K�o���`&��n	�����iAԧw�.��ָ�:������pyj@y+[9D4,9F��O��G54ϑT���ǍX���T�طB�ƻ
7N�{S��Y�|�����Q�yJGd���}�F��3�i5���w`�Z�����a`1�X�f�HtB�$�7��[:�R3{�]�+��2�*L)��}J��p�45pJF=4.�E8=�a^cFq�����V4�0��({b5s'���`PV=����gGSW�V�o#��d�d��y����!�HD�0(��V��3��;�4�sļ}��Z�H�Y=F��6��iu�/v��u���e��j�
��Z�
�	����֦ B���_�j'#]ur:��5��5ե���p.̼�V�Cj⌘[b��LBف��:F� �#G&�l��)�k��f�L=Z>]����,g�2�j/�8�{�巼qtCq�b�{��H8
�<�2���i=�?�R�Lɼ��M����#B�vЖ?l��D�<=}���o��^O���=�8w.��zJ��
�MY��(k&|4U,�i�'�o<Cqb�CC@�A� �0@DA ��,X" � �A� �Ah� �A �ˎQ1x
�?{{��$Y���S?=��˳ܦ�0`�^F�&�������_B7UC�6�����;�l���z���yr~�|��N�;kM��N�y�m�iq�˘{�^�=��m
���Kƾ���X�S�v�h`ȱ����Q�����}�]:3_��7W/K�uq�v���R��9
������'����DQ�N��8�a�U7��7�+��߇Ҫ�.Y�.T8.YQ��ʜ�NF���h��WV0�#�^$�o��+'��i7�k��갠����/F�vce�^�!k �Q�ĉTm��Y���)��B8+K�ht�]k����0j�vn��e��N�HR���x0�(՛�[�x��}�Ӵ����y'wI������ai����%�ϰOwM�%���'�j��w�]���E�z��ѽ9����!�Ҿ���܊l0�u~}����OW�F�uCf�냱�;���O���2F �g3$Ba����iÕQ�d$Bҽ��ϭ]�=�6+�C����/�f�����P���VF;o����������(ݍ#�}t�=:�>�NՐ���g��y�lk9��EB>Kc�ne��ܷL�"Fm�z�o\K�݄�ch�δG�mMe���W,n�+)nag=�*Z37�80�4pb,AA� �A ��� � ��Ab � �X� �8A �6!ٺt��Un�bu��x���RAu�%W��;�"�,��ٽl3�� �f��<&���r?=�Y����"�,����:��2�^���]��-V��g�k�d���E���-Veۓ1kY;��������oGCV46���O3��V�$��/�h�Ҳ]k&����s�,d{��N݊����m�{/p�aCn��01�p����Y�JĘ�6�N<���/Ni::7R��Ed��-��J^�Н��`�D�i߳ڇ��D�L�͕��<�/R7�U�nM;�?�s��CH?7��{ޞ�Mazf{���.w>�/������$�����g]ҷ!�w�5>���9�Y��(�P��Sn�qk�7���I�;��&����'+mA�Z����_d2e���B�´��6��ׁ)k,���q\��`� P��>�����9�}��>���^E}��Z���䞛�iWb�8�G��^��d��	IާՍlM���j��YYbp|���;|�_2�}�8�o���'{RZ�(���^y���.�����6��VB�[9�P�)� O0q��l_\�I<i����#E]a�ѐ`z-�ڪnkO��a�j
�p>�]�]�.�w� �˔(x�D�l���d����H��� a�� �A �,X� � �� � �� � � b
sU!h�QХTl�O���Vm�]��Xw�
<�<\�a�Oi�+u��ٰ�-a�W��N�u��{Gٙ�t�cA󡜟e�J"�RY�˖�\7��^7����kYX
t�	F�Y�)���p�n�a�����Ob�r�{��k�a"Ş�j��=��ݯ�G}������P��`UЅ���«7_�I;�Jy�����׽eak�g{d��]�Wv���Vp�V�5�}��}�����J���������5f� �6-����/;re�Aו��O��ݸ�G�*���<G0r1fŬ-rߜ�=Cb¨eV�hީٟ	�N��]�0-L3R��]y���-_����Ѹ��+!������i�=kJ�lvC-�0�4��b�x/)��*[,�N��lM]�` ���!�Թ�h�~��o����L{
�~��Җ���;C�3���΅�L�9�⦎�l.����u���z5͓�KӢr4���g	���8r˭��۷D����nF�l��(j_���R��ϙ}�&R�J��1e���:r�p�l�3�l��^jw�G�a���o�p���rRڮ]Tz_ݩ�Ѡ����m��fl���\y�~J��#�2O���D�����w��;�h��
7b�$�����w�5�޽$����$� �H����`צ�m�ߠ'%�� �<� ��1[�VԷ�5��+���Ѳm�q�?A�1m�ho���[zD5P�N���s�귬� a! � �A� �,A��AAAB � � �AA	��4&���ޛ�5����n��ס�k�_��]��6�^�p
��!�>��1^�::�c��x�k�J�"G}��%�՟�A���}9�U�{��@���tw"��*B�>�8�󷇼�k��j� 姅��e��=��[��!���3����9�8���o��r��t�����D��z�ъ�4�B��x�G���v���g]^c���bY,��db��-,9��b��2�6�+��a��$詁ǰ9W�ƊGVkʶGi�(C��H��"�w^H��aóW\�J^S���U��/:��JT�/����[j�U|a�r�ʴ5���jv�z^���9��껨u^��*�]�N�(�
�/�����c�]�_=J/��YtO�y�8���7�+� ��;�'�C�A��Dɗb��:�.�%a/��{t1ίL�-X�^1�7%dAnc�v���o�j�f��
��ЦP/�AI����,;�ݫ�;o�� ����E˛wz�S�5_h8��)��W��Can��g�M3][I�Fq�\�*|B�[�k}��:F�z:�}����݉�G6ݼ˷]�8�$;��`Yx+��'���	e �G�^��}k��`Qк�p���������8R�<ey8����}j���!q���=:<��C���׋��hCH��ܽ���0����S��𫧰:}^�X&f���{J�mP.�}	=��^o�M��澾U�,�q4��>{C��}��M��%�sw�7�-O"d��MV�x���A � � ��(AX�b� � � AAA � � �|Jؘ��F��ٙ���gp�WB�����N=�z�5��<x.�P�����8��l�����H�OϷ���i{-�t���<��Z�9�%I>�#�r�>�w�|�al���&F��{��#��t�����C�Oi] R�ܼ��=xmPB,��+0h����%8�4urÕWۻ@�9��|�YS-�{�ek
�K�9�*Ûj���Y:,�F� �e�����Ԕp�n�����N	����yb�;[d����g���ń+X��r��t;��-�bL$�zGsɗ�S�tM,�.�V8`�dKk���{6m��k�*Xfu�0VM����l5��d��M�Ց����v��B#�V�a�bՑ�;����P{z$n^8��墩7�K���%K�)T�b��`lU���?Ygy�-}uZ+�d��
����*]����a�� QY&���˫�8최�{r,P,gf���ɋ�V�݁w������f����:|�N�����{\5<�,{�wyE�[Z{�cJ��.^N|v��Nħ_\M�����</�M��Wr����\��j>5�����mΖ�RNk�Hr�?���uӕ[�% �k�R2ӻ��GO�����6�UL�,#޴rM�q�Z�j.���������!2ɓ"����>��^ieq�;&6D�}g���,U��^l��.��iˤ~��U!h*-���-t�aDWT�8$@-�0�B4h�Æ� � � A,X� � ��
AAA � � ��6�Ftq�+��Wv^_=��ة�#���7��x��,���_�,�G��^s��^��nh٨)�p��ۃaaM�ް��̩������v��q���*�-����ror���#37f���!V�Rsp�ѽxD6����t0�0S�${r��;;[m(a��n�{�sڟT��`�C6��0j�pu`�`��m�F����Q�R%p"T�Ml�F;��D���R��(/~C�k� WV�'�1�����y/aճ#[�ƙ;���'��&����Nԑ����g�ͭ����ff{py���s�+׸�Ug�{�ݾy�!� �J�w��;K/F1n��X�°�b���93M�W��]#O��ǎ&n�m:����E�mH�^ڬ�*�u�V^:;M1��S��wۛ�:�ٲ�}��|M�h��P9��{L�ܥgl6ìǑ���Fd��ݵ.v3��`7�I�tŵ����op��L�?Q���È�ݦ9�|��\?�T�m��Q�Oz{�^(b~��w�s�������C����0u�Ζ�bY���j&�&��a�S�F�7��٫�n$7����������;�$,U��$�|�k~��{V-�Ǫ�Zp��A%�㩵�EDZ��_`�S�T�0�H�jߍ�D����ɾ��$>'����h:S���}�r�}'���r��B;��!���Y=�_k�:��դ�^!R˼&T�����mw{�3�0�F�*=��\x6���S��ἂg���2\�Q�&j�cg�&m�
<����:���~}���z�-���F9
y��N)�Vq�FQd� =��������&����L[��s&oN�,6;r]��{<��ڶ���M� K�;}:e��_T]��šd�N�Mjb���|Յz%��0=]�s2��uU1�{8jY�b@��IC���gOp�2���.�Zyx�߸����W��T�z��<{��#ל*�H����^9��+����:�WtݐW��C��J������}i��ʙ���xt3����GD��tdDP��.���
|�(q�O}����p�|��6�ϟ�>T�g�h���'�W��I}��V��>ۤ阸�����R���UV��z6w��zm|g`}��4�G���S{�����u4�\���->}�D���_fY]0�������Z��wmE^`��V�Z��n�.�k��n�����>�'�0@���%2-³�9���_/{x�n�w�O�$�/Ԛ���%�r�I��s�g��ʇ9�s�)�W�F9��ǌ�'mZ�m̓Ӯ��ҷ��uw5t�)�Q�k��P�V (���㳷8L�yAB��WD;���[����O�l}��)W����>�g���'�}�/�8�a�����y���{���/!���x�!���35����_��y8N�3ø���=�j	7���0Z��ڭX�6JǮ�D
���U�BJM��qi�]Y{����L��m��o���tE�(�o�\���`�U��Χpև)�����^�SE�;
Y �ޅpx��.ܛB�xp��b�V�ޫ�0��m�Y����u��-���Y7-�Μs��T4� �`oS���L�_��.n�r�T{��t��O<I���`��=�Fۮ"�|����sA5R�U�X06�i�����2�;���+t^�Wt�/�����A��5��ML����x���su��TY�.�KeM]d̥+���3W����= ��g��9ኟ3}V\���*��/cH�~�Y��V�N����0�^�fq��Iڬ<�ء�u�^l­rr4U�c)���&���v�!�ޘ7�4���}�}�������d��&<����y�o\q��8.���ʛ}��M���{VOd��wnw�'|�g{�=�z#�#��(�s(.�q�L��5��_��MiU�mns�s�V�#�fg+M����xB(u�6"���Kj��k+�R	FK�*�je�ؚk���3���ƃ*ʹЉ,��2��U�&����E�&��"���s�#Ϟg$mM��TLiN�l��\��#t��dpI���n!c��Ak�j�j�6Q)U�caZt�e3�!Aд#�TIf��X�l��`%���[�'ȥ�W�¬Ӊ��.�KE�04P�A�����:�ܾ�;t�Թ4Ъ.FDEHI�4�m����\�F�Ë7����e��q������ZVڐ�(����̸YP�=8l��e��*��ԞR��ұTQ&��V'=�3EP�]�n.���ֈ�OON�8pPQNZbX��B�K�V1��ƨ�m�GOm�,WV�Y\Ft�Ӈ3�Q�D�b,��	�R�"��D6�e���V1�:t�Â����6��ust��F���AA����Ƌ�����Z:٣���#X�xd�;��b��J׎9Q2Z�V�!q�m�]�H�mM7�M[�+�]Z(u�+(���U�XC��q�V�-��C.b�,tzzt�����`�auI(�+*�7q�[Z@P3*T�$̵�K
�F�REj�am%u����"��+ ���&�hl��A[�G*$�y�i`{��6P����<8zzxxxx�T�&e|�թiWVLT����۔m�3[J�\\XQ>��|�c�4�ZLt�8��-Y�����-M5��ѥ��4;t�4�8p�EC.8�j�`���d��b(�(���帅V�0b�[1*.S�+X�eY����5ۊ�Ur�qf�֪";�u5�����.�P��}xWZ`*x&ӹ5��b{�J@F��;8���<�oI����^f8[��]�k{��{ڜ�j��|r5�[��;�e�+���J�줲Au�m���>?}�p4�޾M�'IvX�Y��s�\6nB5ȫ ׽��L��G�Z�����:�b��Y�z.�v�e����{�zM���s�Kt��[G��0���$f������-��;�~l#��c�<y�5/&�s���]e��)��7�
�7�����A��݃��I`c��"�$����i��4��Ϗ�/�A���ˁ�Ϫ���(;���a��ff���v��ٓxs'I��&AL�-��2i:�gιzM��&�n�]_��zW(��9�w�w�GN���j��d/=t~j��'�}p_u��.l��'y?e�����=�_I�{��s��N��@��}6Q�\��K�ߖ�ۣ��B�O��<�`jg���eΑ�9�6 ��tО����o���j�:�`�'��%x&�F�׳]��M�<['���*/���
����lU�aBE��g��������3r��N�g䢌�T�U�����u�Es��MI�B�����J����P��g���ܞ�%5ն+N?7�S}ҷ��	���,~�wI�f�')\���p޶�i����W��{�I�oy����f	���VL�����N�bU��f�M<���.���
��Gk��;�����}�=�<�K��
��DxB�Nϯ=�oW���j^q]3������p�|�`1������lZ�g�exsc��Y�w/~�Y;�/K���;�%is5�d��`�Ս[�w���#�������=,�'����,n�{��1ӗP0�.���Fxά�ۓ}-��&�N���OɔW��q�U4����;���A� Y�-�[O?��N�C���`�K����}S�sSNd
��q��X���s=������� �9V�1/�c�^D�3�$ξ�챉k�Hn��1���k���f4�M�|�n2�;g:f���2ac���I��|�a�DM����wC׮���ck��̭{ٺ�㞧����	:eu!����<��7:��Ň�*��Խc�^��oqЂz��ۣ}�Ǚs���\�d�s�C m�ک���a4�P|+%�P�@�:��]�{����t]��*}oܷ~�pFO�N�v�SI8���͉)�93�N�+S���=��/??����) �b�;ߕ�����;���le������>�t��:_g����.�z�6�Cn�����f���T��1+v�k�6/K����y��|�y�Qy4���j���ʐSEX���9�o��͗����ht�u����i�.�n7�ڞ���e��	/�0����ֺo��/=�3�΂g?yzn�U3����ž���|+&�V��Ģ<$��t��v.��;�9=�&�{z�5�M31ʋ��1��Dh�_ʶ�`L�� �^��@x��gs`k�pI�`�KrU�ٟ;�<������%�u���{���M�C�q�wk<�{�����t;�ܛ�{[�{=�^��e�z��+w��nF�|D���<$8�ۨ���纯|��A����"��a�]`۱�?��@�wS�^CԱ{��� �s�:\��9��>��xh�\"��x.#q���Ư��)_P'�	k
���w�B�o|��V�)mn(�;"_V�����|L��̯V��d��Ut��ԕH�K����mr���������~@.��gيSsv5�#
�������=:������3(<=LP}s�z5�l��T.�����sN{37��Hz� 7o�	�=&���zEؙ��������մ�� �{��Ԇ������:$�":�O�x�n�h�\�>�ہ�NZ�)�p�"E}x�l��|k��xzE\C�<��}S��ߐ�M��-gּ�Z���L폜e~��L��:����|ty �7����	<h�Yצ{f��Tg�a�\�#�^S�t6*��w�|�}�c�{щ|��~�|�s�%��ݮ^��1�g�<jY��d{XX<z �z������pu5��M/�N��wY�މ>��xUq=G����uc�((�<��_��8:��T���b��x�w��\Oa�+���~~��o���N�T�r���Y�~�q��M�$W'�0{��i{�|^-�Z���m����Po|�)z�:��8�zAî��~?�kd�^a��b�䗵AM���-�+���_�����7�`�VPj��-��-��ksw<i�U��з�@��]�R3���U�r���:������cG���t����y��n��{���f��n�:Yǿg�w*���%�m����<VEem1�{�_5�(Hd�����7&>dڛ�~��ͯ����|�����߻>9��3�ֽK�7��q7�¢�I&�0��-���K�w�b�]��w��^�}���#����=�������x�	"�D����p�X0ϓ�YP�vI�z�ɓ^����NU����ǒ@/otf�WYث���K���jn{�?p���L�����/)��ޛ����{v>UҪ-G�9xk�����s�F[9�>8*�e$��G7ͤ���<N�k]�ſ�Hw%�x����vV������>�������Nn��>T+{�,@�+�Ķl~�݁Wr�~�{��X�V��DA��">����!޳��4���5/��Q�sw;�zOm� �HrdT8e����pA�Xl^˷��s��(�C���~Gr�{x�ߌ4�;<�zw�Ycׂ��d��=�a"�"`ð�!m��$c���-�L3����;|	�yt�w�M�Ow����^:^ԇY�y�3ЧW���i���pN_J
�F�7��ݸ�p���3�����w��᳅��;������p�=t�-�^�-W�r��[�5��0$K�|��Qn��7�;�(ݟ��`x�N�����I�"v�r�^wC�h��E��}���D��h�zh�n��oI3��ƚ�j�F�y�B��n>��Y�އ`8ʺ�v �<�>�����1����Ǹ7���z`��T` Ģ��X�]�[�ë�	��r����1G�o3�߽�r]�
����:Q��8S3��w��k�QoR��6�4j���bZ]Vߠ� ���/�`���lC�ԧ��L�[��=®��כ�RV�@s_�<���l5�=�����М���7ϯyyFj��>#:�϶�XF�]�Eׯ���3�j�𮾪z�}�NN�ٜ䰫w�f��UP�A�@C��v��H{�޸=�xx=u��I�>������6����KSD��[��/H�f�7ȡ(��$�=b{�x���H��(k��ɱ�g}�o�;I�1��ۑ�2{ʢwS(3���R����`��ܱ�7; *��	c�k���XN����8g�t,`����P:��m�}�=X�e�r �n��R�j��4�E[8 �؋��s�����vk�5�雬|����U?q�_(�5B��^V��Y@1���v��k�/��&n�z�����C]	$�sg#�$��Ю����k�=�*®>�;�]�A�P�lv�����v�m� �0�T��U���Ց��὾���=�	$�h"�P�%��^7;�������0/z�枼�jՋ��y=�8��<(l�(yX0; �,8=}�χt�K���=_.�u�m����ݦ��oW���]Z<��q����[ǟ;{�s"ܴg����,lko:f�N7�<9[����Y��ma}�����a1�'E�5�N�oޛ���9g����{��q�C�W`/�F�G�sp��Hj߅�V��jzA�>�*r���}:�Z�L~>����g���g�6L���z�G�9����~w��0=�rζ��D��~v⩹��H�yn���Um����P>���Z*�ty��I��4-��$y0t�ȑgfޖ�B�X���|�����'�ӡ\]�F���Crܺ�	� �J5C��;���Nc�W�c�`��zF��KP�l��	NJ����T�|�˻Y3���iAk�u��l���o{&��v��n�	�'�9�g��U�n绮0[�d垽-[��x#[�(h�C��j�ރs��J��Ps�ko��<5k󓫸e{@�>�hmX���_���(�m�j3RN�n�^T�6���уǩ�ݵp\��P��J���;�8J}��ߙ�p�2ݖ�F�l�<l�=���lӚ��i��W1��|Z!�'��<3�ϖ,�#o�i&���zOu;�~��-��x���.%#�r�,b@agτ�z���ݎ'Cq�M�sx�n�y�8�^M��?8�V�v�\C`�痢���'#o�{~��ڽ��ؤ���ٱ�}yÖ�\ՠ�z��yo���w���6�{nf��]^���p���v��8&���58�-�����9hmtq��ݲ�o/����8wu$���}*4��)�o���x3���y���p�M�����CL���������L4�-[6`���Y��-H�z�s����7-3���A������nv��)6�5g�u�乫�پ��&J
�ƗWmV(y��}��U4;�K>U%����ass�㦎�5����N���}𖆉�g����v���*@=`��}k�������7��Z=�|e<u���K��w��������!>�c�c��5�I��H s��y�]*���{�{}1eb�?Qs^��7i�\3�m@$����!��9PD� ��7�u�Zv�]�`�;U,+����:Q����!��f�Wz{���˞�"Fg$������~�`oX�Et=�6k����+/�{��Ii�'. �$<����4D���d����?p�_],�Wl����C�X�ߒS�X3P�&Hzɪ���T\Q�b��F���U�=����6��{g%h���	�31��"]P����/�	���鶭��؃˾���7�=b�/8e$K�����/���� �ZvSZ���h*�k/
���ySܡqi�jCN�"�4y]>�{'SG�n�|τU@$��@@�5.��o�Mj�.�ңXD�55UZ���������[�>�3��Ed,��b=u��0��V�	UU�]U	N�k>[K&w3W/͠sk~A��>#�����=^n�Kq�f�枧��~�:�x�{��ݩ#3��Cs��ܸ=o��S��Ǚg���o�d�S;�z7�tCdi65�QaD�6zک�Fc��q�?�ܳ}�=v��?޴�2���/���>�ǁ�$֙<m���f���;ׁ��͕�3߲^�h�+�� _�z_OgE�/ϧy���{�y�C{(��*�g���Qg�T������G���g�~��(;�3��|߯G���<*/.���赣]��䕣�X���x5b��C��]�*}�R�`���I�w����������=�؎+��R��@���������fl�hw=�=�*x��m⎯v�J�[7���#�0M�Ϙ���y|��J,oj_�4�?MNN�9|�롍i:h�v@& ��v�tl18/�H�� ���8Pgq��?7��Kڴ�-�@矀(�g��ս�k�|v;=�������9UCrb�cJ��g+\��.����QV�ݫr�@]�	��G�F�W�Dg�hge����+�{��*d��9�x��9��~����Z;\3e�n�
���x���M��e�䬾Ԍ�N��Q��,h��'w��:d�s�`ө7 �t
�vm�S�h�h�T��yJa�q�w���k�e�(�!�k�����ij�ל�Qj�C:Ŧ͸�
���`�:ì��,a���� �;m�<��T��7J�f]S�����v�w��zn �s�u�{�<Z����qGv)�v��a6�C��$�0�[��7/�><P{{:m�Gtk�G7m�h^� �%b�Sh>w^������~�wQ�������:DD�f�����v�ҟ$�'�0��<F槾A#��3�1� E��H�A�9Ue�[��n�r*�Z��N*g���
csq���;0�M��6�2��ۑ'i�{U+ns�	<H�yT��t
wo>�2>v��b�N��Y��h�0U8*]���B'o�W�i�"��s�⥖]r���i�'4m%Z�M�-�A
�ݮ�t��ԃ��&my��%�=Q]�p��@��o��4�q��[5'���j
ʏ�f]��4�U�;��kQ��g��Ô�r��85̆�!�EcT�4����e����・;:�.�C���Yxɂ�R��|�J�9�-�X�5�e���|Zkh�	$���/YC;��Ah;CvP��Em�yI��A�I]}�H���󖐔��S�􉎗�T�u�+�i9��4��x�J|jҜTZ�7�F�`�koz\<�愕UZ}zB���xl����kbǙ�9�[�y�7i��k=�圌�����Œ�9Y����p7�$r�m拀�bL���o�.���۩�c[S��������}��2V
V��n��tL�F�.0X�gvST�JĹ����ܢWz�:�����HT�����59Ƒ�q�מ�V��ˣ��P^�ct�=�7/���\W�<.6{�c΋S�Og���/;w ���E��;�#�9E�˵/� �b
�Z������������*�:���v��&�X����^�ٗۥE�n���e�7�����tb����s�<=�w��!Ѽ,gS�ujà��4�m��iĹ�-5�6�l�{&��{V�~м���y��">~H�=�4nxN�\ݞKˉ� S�%�[=��-�ڳ�w1��k�R���_l�Ϭ2�����0����p��o����x�a,�%2��K�����ґ�6C{B�}p�U��hS��&>��>�׌���۾��VAш�|�v!p�$j�J�}ŝ��ǬiH�H껈=��e�՛\01Je�ǡ���EvVCC6���<�jL�{ۣ6Z�Ux�Gn��T����|��	x����F&�e�k�?u8?�`L�n�v���D1,b�6�c��4�V]�����W)Eѣ��=<��!�I�Fe�xR����)�*"��0z�*����F�G�͛<,E8��Z��垻�hҘ���e�KU�E<��"�9e4ݶ8xxxxl�5*�Q/�x���2j�QX��UFjݎe��,On��i�GON�8x5/J=�O�U�Q�3 �QTE�K�1��f�e,�Kilp�Ӧ���rj�&��V�iA�fb�KJ�R�AiK�X7�8itl��ѳ��Q�ri���Vbb\����U�[F����Jʞ�X��X�K�ep�ç��-QUx��Qj�2Pc32��P�b�&!\B��YG2�ٽM��g�͜��
̯.,T��b�-���q���2���"��E�e�d�*X(�,����P]j���E���[-����k,b**���G���|0�����疏 <�ab���=�&lE#�JK]>g"5��)�]��!ж�්֝�6˭�OD��@
����x�l����z���{N��wPn���۹�����W�^v��am���T?P�����ݧ�s!�R;��> Xgne�&v����i��vF6����4U���*�!H�a@��V�I�������ɾޛ�{){�-��B�Y���M�D�d9�����܋mIK7�p�k޵7N6�R���)�b�<P�zd^�].�yf2w2��6a��V������tg���__��ؾ���]��i�W�MKhg^���{
��I3�aG�1��_=p#!��(>��\��Hy�ղKc'��u���TC�5�Ҽ �qM���h��1,�&���e	Jjw��{���i~�<�@>sȜ�(��(�݆�X쪻3������0Wm p�����$��|��t	o.IRkk;'��#��t��xMق�۳[!��u <C��K1����˰�l8�(�1���)d��A1���n`*OLb��;{˵���h�8�"l
��uv�j�:���rt�z��^���R^x�O���o���xY�:���h��հ��7y�a�kL::z_�Ɩ�p���\o���O�~9`�)���-C��%����묭��'��:��W�_N<�˻�KM�y5�*��$<�X���"W�F�x������g�cRT���B,�T��]y�M�]�0����x`C3��Yb�Vl��pr�\6�FL�b������O���AB�D����dmm�Tg�û�Y#��$n��E�)���������T�u�OH���Ts�ʞ��#;w]{�[�p�s�{<Lx��s���cK��.�ഇ�v(:�q�M9f_zn]�=>۝�9�ԻG�DB 3y��{oh^���w ^5���O�߲���_�?��C�Nǘ6��wS��T�ݮ�8Χ�f�ᡝ� !�s�.��F��^�{!�aV��0��psI��5x�r���08�4�p`�8l�Ox������{C�v�9�LLub`c%� 6�e�A3E��}	����v���,7��\��������^m�hP�r48ݎ[�a�S�h�7�=�u���.�0�5h����J�����^�CIk�R�6�޴�>R��l�<������m_���}]{����#䔺Z����en�Y�s�8fnブ�pC/g�ϛ��S:~��;Ń$`���f7^�m�FK�.��UMn�#�NE[z��A>��0�{R 	e��z�5qMp�p�-�c����$��ޔ�!��3���nU���osW�!s�~�ɆP{�1iՍJ�5�Ly��5�z.E�q��$�^���r�X�,��Ծ~��yg8�z��_m��P8�t8w�=��"�EY���c�2�K��U���aJ���Lz��6a���|���U���7Y2�c�
�2���M��փFdw�����U
2nS�J��6n�]�{���;昴iq�����H#��ל�o{���+Ð���b}������1���7%ۄ��-�A�y'�1)դhZ�*�p.�rD'}�[V�j��7��C�\[GW��z��i�?�&H~�]�n�a�>=J�,`&+o"�ME�QQz�f����@��v%@����i,,����t��ˮ0<9N�ʼp�7��,�y65�&�]vngq��Fk����S�1�9�b摴Msӿ7�|��^(!�����^�R�S�|�c��,��xsJ����8[�XU,�疳P��R�n^GjJxw�>;�� ���4M8�;/�|����.
������[�/8�AQ�-Y�:�0ʢ��t�yJ��Kݾ�sۇ�{\0l��u�bt�b��q�{�!sr`鵽025�z`kd����'ǜin���A/�e/�4���&��-�T-�,��l���i\�*�0��fѮ[���fY�%���ԨO�Z�L3ztN���嵺�Q����8����W?�{�|fY�ㄈ�Xq��a���L��]���;r�E.<�Z�&�����M��mQz�f�����W���~�y�4?��S�S�g�fߑ�v��'����5SQ����N�or��'����?1}�՝�߿v��<��ž��'���kW���u�F�c�Βj�Q*]�j��V9�/*mF���.'�#bc�&2�3ǌ���8�)loX6�׬���a�vpo!��0$��y��kA�@�i�����T��"f|tE��&��\3`.!a\l5�zX��r��3Jc3��/�CW?��Yydc{1�\�s�+(	��\m:naP�E3�TѢ�:3aqZWGU�P�!��\L]�s̾7����F�!k��A���+|
�G\>�z�SѾ��I��U��՘�Z߿k��~��?���Ϟ�{��s�5�d&Z1�5pݽn}g�sM��K~ݾ���w�/^b�!o�2��`p1m!8���!=��{�������7ԉ�x�TǷ�������	*a��[ฌ3�ص'�,�_|�9B|$ �=� �������s������7�T�+W��&y��c(�I�s�2��i�&���>�������=�}I���y}��.%���eԆ�.�X4���/ޜ�.�X�R���)��k�n�4��@}��-�_���3����OU:�yNp�pΙ��Dct8�C�H��8�*�zP�w�%�it�tߡĻ��s��S�f²����'� ��ǘ?64�q����Ju^ʒ�`/g�`�� ��Q��Sj�w9��k5��s��4kƭ���|~���y���ͥ�!�|���S������������/�7&�y7����e�|.�a�ק�	�`�ͳ�$��-��<�@Z|���e�;�#-Ls ��,��k�W�������P�+�s�v*�r<ou0�0�{����Nzt�r9�p�9�G� Ϙ�x8u��"%���;E����o48�NO�tc��#64M>(�==�H�b��XV���ەOe�2g�
���'�����_�;j����ʓn����ܾ=u���b�t��a��?�U{��O���`��9�J���>�E��k����~�7��e�\���!�dvO�~�^=%�h&+��ύ����M/��	^K4�7���ׯ>�,�(��E�s�j���}ա��]լ�:��q2��\��i��V���宜OM�a�r5c:<�U�P�χ����ʀ���]{�4���L�W���׊�R2að�����	��F��Q{YO�6�š�æ��y��\ટO={r=m#RSN�e;�Wq�����;[U�Y��>Z�K,㞠��7�X�������JQc�/���N0J2D7��מ���Ȯ؉9ϙ��M����+J}I�	Fq����[ռ�|wA8���a�"A�V
���Ts�{��輤��N	C$���er�&���6=�e��i��<$���/|�K���n�٬�tƕ�}֗9�\�9T��q{�.�hЄ|��#�T���W�]noTǍ����cr���N��sw��t��*�&�[p��u:5���H�#^��L�[]l�O;�ΐ�p[B�4���u]*�X&���J� �tO���,�l3��!vJ�nxN����rv�^IRk�;��kz�BH(G"�p�����^�"E�z{��צma#����öL8�ki'.��� �"� ���6�2�,W��T�yz����n�*�������h�"<�9	�G�n�vIjOaj�i!70��LZ~Y���ӽsPs�L:V!��)��� -)��c�����CØ�����p����z���s��c<��{S��܍c���tpO�㧜H��aD����B�Q��ޡ ��D�
��|֡Sl�4r�l��Fv����3YN[@��T��Txg�T�קvm�l0g��AĄ�F���U�A�}�ڍ�\��K��Du�C��a�Ʋ��=�3:ĿX	�,L1��l�J�MP�$T
�+�pXV΄������yl�vO���A��i' �s4�v�1\Ÿ[���z�9�f��]9l0w��S��(�����==���1��݀��ۆ�W�3Eډ�b�B���O^ެ��2�+��T�����h\J��%�q��q�>���_�-���Ǵf_P�D�ʆx^�c`�t6���Шrz\}l��$�}k����ݑ��{ƍ���-��9�Mq�Z��\�t吶K���RT�����ay2�d���;��l����)���fp�Θ�Iu�|F%+�g��A9(��7c�Q�ًk�([����/��*$\K᠂����pc�x�N��fq^;.�nM�I�hٯ�~�-?P%���e���ջ?���WSv[�Z��p�'���Q��Y�3!�C��A�qW(5g�6m��l�瞝���0B�|��������1GD}����� �9mZa���tJ	^|�7^�ՅW�Z�_����@�O3�ћ�yTi��^[(�q�-Z"m��N�j���^�wZڹ�\����A����X�hR�*��\�_Si����י�����*#�Dkz<`Ⱥ�I�<�r��O�%73s�I��L(W�E��2�-ʗ�]"�s�/��I�l�A�c���B��>�(N�eE ��e=r����n���T��k���娺7/S�����!��l�E�r&��l����Q�L,l�(!��P���G?k�e�i��Hz��ng�W{ݝ3�^T�z&*â�K��4H�f�t�m�^��;�_��G���h�����.��|���"q-�«�%s�P�r�ͥ>,Qنø�������Vھ0B�2s/(�q����se�����P�~1'\]�����̤�u#\P/6���{p�-z�Q:7��~q�!Kϗv�gL�;�)��,�R�$��1][�o�����e{��g���ݙ�MKܻ߳�si(�#���,���N��Kz�%�=x,U+�[��=g����Wx����|�/>��y�����tcr��B�x��s� �����r�Y�^qt1t�;+����		���أD�$�P`�x@r�@`�Ŧ�5�u#[f�еf$뎰_�s�PK�Z��-z9c\����)^�<X8��ɡ�#�����9�L3&#rKj�jT��zX�L��l�I4��mhN٨.�nj��dd9j��w��t#m���fI�n�6�%�w��3�/;[�v���o�$����̻
��������bhY�5>XGY�*�5A�͐ﳖ�Z��mHw���C�B!ʠ���0��m�<S��@f|����l�B�K�'��c��<5c�m���G ��}�r���4�m:m1p�ۤCDF���B'��;$pt~��A{LV�F}if�۶�e�T��iR�A�*�%��\�����ۘטNV��}�r�}�E�����|��!�h��>��\�KsS��/��L�T5�tI�Nί�U�gwc�N�9�w��7VI���Ǉ�����>CGmx�8��f:.�Bx_!,�־u�^�8ּ�f�:���5IP�ػ}l���}w�A�4n�|�'NS$HY��8خw-���Ve>��s����EV6WL+3.�M"��[�JPxUg�;y^]����z�Q���:_�t/���X�=n�+_ir��T��s{-�7)D �y���T��C���'�e�����Pn��o���/�ܨ���n��ج��@$A��t�)��\�>o+�D$��L�D�(JSǭq���׵�
�9�a�]��8OsS�y˰�u���i�vR��ٴ�[jQu��^eAoT`t=���b�_�.~�Z����hg�n��$ʶ\3kLh�n����v�4+ʇ�⮗������Ƃ�0���}��w99�¢"�ѤZ��*�?�0t��#�ku	�N�`�y�i��.�Te��w:��M�8����߫{d��NO��o�~�üƙ�� �cx`zh���sLڌ�je��l���:���<�Y��h�?�k���.;��p��vB��W��~���u|lH�%ؾ���Eo��x�5t���-[%��|@>�zc���Hr^�;�}bM�����N�}ۊ}:��W٪������&�
��
ߋ?��A���� :"طPwc�tK�F=l�.��!�����������$�^=��~�&���!%���$@"x�v��-�^���9"/�"�;�ޥ���%��iid�l�ץ�ލ���7s��<U������[ي����ƅ^n۬\OF������lܻ��aMʹ�-�����t>󋮏4L�=��zױ�V:um1jGޜp�
�M��0Mt�a���ǥ�v���!:�h��հ�nUG��ۙAlG=3���@N��P�;���k�ͬ�pc��tS�w���#" �O;�=4��MJ����7�@'�xmhg�D���
>>K���ѹ1�_4ͷZ�2.�6f%N;bo4��A�dSd8�x]�K��yc'n�~���ǋ��J��B.�^��cX�;W�%yu��c��ɭ�J8R3�	{����"K�k�	ő�%��S�û)�(}ù=҅Huvd!Q����N	xd�'��J�6`oڴו��R��t����W�8右��3�>�"z�djv0��gd�*\�Γ�xN��H�^���i�͂�jJ��c-��4�v�x��Zn�r�<�����������-�{�]��^I��e'��I���"����t�.ʁ��*����R�_28��6�,:,��_���z�|����t�RԶ-�]���%�^�+n������A/CRi�K�?X��p�Z}K�����qv���M����}�<�Z�G'�����U�R$G��	�U����!�f�P��a���uEԳ����!��OH���V�c�Jr،y*�ƦX�p�ۮ��|_Q!��$޷}����۽���w�,M�a �^7����H���&{�o:�]�o�U�f�m�h��n=�9UY>��}�N�W�K�[i@; ���-����斵t�~v��s�ڨ�U��s��Y�V�������l�;��ӷqC���
6�fn	A�2&�z�䯪��> �_[������f��(ƥaꝣ��]t�s�u��H��5��/�;l�����GS�m�:���+�]�7j�{.�z��v4Ǥt�Q�pZ��]5��*��5ZM�qVl��zE��wwY�w(����q~�z=7,�����7�m.������	�'�}/��sO+�R�U��c|�;��T�2yL���s��P��Q�"���s�viN��\N���W�$Wg�33#��[���G}����Ӧ�Q��uJ!��*��Jт�ۼ�y�ܛ��H).}��?_#jsc]��]ӹ۪�"���omN�yБ��#&v9�qM[��Y�c9�94^	�v,���YHbp�Rdc�$��u���E��opᗮ����,�ߵ��s���ᲆ��I��vF����#&GO92\�[T����C�,u��7�?mAu*ڌe�K2w9g�1b����l]+(��u��A����k�8=���Cs����pbq��IYO�&����_2m2��6�T�.�tbm��6"yrp�ψG�A_EU��'M��p�]]�&6͈mw_K����R;�j�����H�/�T��X�Q�n:��5�ߝY����ݥP��5�;u���z�L�{s���˵�+���Wݯ�%��셌%n>�����zd�P��m��c=�ñ�sMwҨp�f=�=t��L��D�!����1�y3��p��y�]1��b4�Pgn4�Ϋu�ZT�p�iV����q��v��~���] kCstyu���3|9��2����Rm>+Q���$@��zn� :x)^軔�G�AL؋���mYz���{��nz<�ʏ���WQO�v�{u�m?3%��s��
�,O#yi�8���H�n,c�j���z^� [|��O3�rt����;��[�&sa>5P�n	3�l�\$�֭�K�nF��0e0�Y�7ӵ��t��g ��a��,h�hA�����\0s�\	FK�\&�s%�72�������K+6�VN��#$��\�UpB>)_v�4�ގ�aԘ�xM��dA�J�;}B�Ge�_=�fc���5�$+R��F�Ц�G,vbb�ݥ7xSf�]��U�>�b��ym��i��tgr�4C��9/w��zx觐�kוx&�c3��Y��q�_xǇތ�ٻ��yv]6�N�ˏo�3��]�/���~��^��u(��Y�8�j��c�IԳ��mG��n�'��)qO�4�L�]D�1��6HqH�MU(3#�AT.H�㌶��",UH�*�B���˷1����:h�j�U��kk}-[k�5�LZ�ۼ
"�m;�r�QAa����᳅e[cj�[A�eh�ZTf-Qkm��*[�4�m��q��vh��F�Dq1�4�\�B�d�_<�*�t��*�*6�]ҰETz��M8���Y���6pX�J�jV�o�|��J�v�cY�Ssk2�Z�������.�M�6r'-�1��U��`����
Ke�媪��SHb
�c�a��᳇�k[e�����Z��1�XƵZ���im�[bՋKX%�ֈ���*QX�xxxp��Y+F��1E����Xŭm
����ND��E���)tˍ�,{�4�������Ӈ���UE��J���e�{qSc�������V�eb��V,b*���TEWfΚ:lમ6���*��TJ�R�
���m�����ҴE"��Fѷm�f���++FaDTb���,Ki�Ub����1�X�*�J���4�UEQkn���2&m�����*���,��V��P� Qtļ|�>�Xz�."0���1�/^U�����<e.J�m��h�
�&F3�/~߿~��4�5���3�s���{�a��C�CM#��0a����#���?aM]P�A�(�vb�O�.��;�����`�E�k�㙆)�n�����E���$V_��n����*���|A���O���5�<�DS��A��tZN"���0�Š��鐱�z{^�rj���Ԩ�����������^)��{c~�v����s��Pg�f~�r�I_T߫7�_F�jC��	�~�R��~I�,11�H���\ŶS��셷��W���:��|��{��	�����V���aښڒ#��OհRL`��
Aa�?yg��&$�U3��f1U���/m#�������#�Pj�(�3׳f�V@�A�9RNǘ������'r�`����L$(�B��L܄li���a��(���]��!��r�Omr�n)8s�d�[��Mj�<�2�����e��N���-^��+���2ǰLRuc�J�UI�4Mʈݚ� 6��UR�w��.d:ȝ��}g�"1� u0���ݧnY)���L�ۘ��i�G
Ztk�w:.oI�|@/'�Rӌ$v;/����`�����5�� ���ntg~�k�y�������5�oNV>� �Nz^M�an8Z1���3L�S/h3�S�{����\�]�2i�n��q������v!7����WjJ2�;��"ٚ��� BdW+�:�n���ĥ�Ǻ��gRѼ�A�ӾF��iY:�_���ו�(��~�P� ��# "@C ��(*9b�ۓKZ��9�����2	�6^����w BF4�r�_���@���O0��	��.��ӛw��Dܼ�d�.�B��&n���0-��V�zfä�0��6??2����~�[�k���gg�΍���e~xՃ�)0��s�U���o�IcA�a+�d���(��f\��!�f®�S��!�;j��sCEHv��%��Q�d�q[�J���G2��u�$���k̵��Vl�ݪ�}uE�/��hEïK��#r9hk�e1�$@���"����8�B�)����g8mޘ�]�n6{;)C3�O+	zs ����>1��/W���$nh�Ú��TP�m'{%�%u��z33����f��ƥ���.Z�9�dK��"}���<���fZ���n�g����m�^��I����k�)0EྀL3z&e�A���
Ѧ/�]|5C��"������o柎�u�gt#L����7i�Fd_<P�Hr� ר���L��m�{`3p�1B����a�^�s�C�AN&3%'�{Ǧ��Ƒ�-@_Aʨj&���.�G���m�����!C ���ӱY��ٮ�=�������v��]��+Y��"MM��!#]ˀ��}�;��DA�?�7���?:B�C�F<�����E�V
*�ȍ��6JWjQ�_]l�`���zƷ��xC�~1���{y�y�z���?�?F ��$��'� =� �)����`�#a��tW���G0��8���/uQ�]s�-m�@X�0�eV��.�&k[[Z���i=F�ċ\\:�a71�T6)�M�?`��4(3��mCƗxO�Y��Tb\ӵ�u�<n��t��%��L�/]���3?c�PZ��QGÕ���`�'Q�=���*�K�Sͼ9-�����'��L�S�a0La%B�6s�������2d��m���-�͵�ӓy�\�����Ɓ���脝pc�o�Ҹg�'X��|E-w�R��ʵi����O�a�3u�wp>%��_'a`�E�a��ݕ�c�酎D]y'��"Yp[��`Ӗ̝<��L��_��?6�m~����]R�����t��B���(➗���X��猄��J�C��͔��'�c�1�!c��	*W��0B�����O䳪K��t��Uw�}ݭ���Gov��Ֆ�+�t;���4�^�>��k���ڹ�p��'��}�!���-��[��kI`��w=����{
�|n�;C���� ��ÿ0���)��Z�=��g��f?��Su��Wz�:��9n��@"�R ��9.{���\�l���0q|��B���K��ub�0 ��#�3���;J��<�iJ�9��G�N܇,i�@��bl�}��|G60~:�*��6^���P��ko����������������0�!B��DI"2 {�o�Z��ߞ~~)�[m��ɶ�
SGS�1��1�B�]31a�����A�ꮌxHn��;���e�^�޽��/�92yV}��ܞOş�_G�v�1^�tE��W��;��c3�K�z�j�<q�fe��C���q"'��w�K�:]��&�;w����H�D�&����4)�{��EY��G?��鬯8T�
^:��ʿM�+�t�n�Φh��,
���;*�4�f*�������~^�h*�\��_��P�%�ǲ����G������y�`e�y�w�ۼ�k���zxgm&l^�ڊ��6��X{�9��>���"���h�%=�EǤ�-s}uNޫ�V����aԄ�W��%6X&Pd��GZ|�gXV�f?�ޭྲྀ;�
gH�Q�o6���� ؇�$6�y=���\�΂pK�"�#4������\��!F.*ČUwN�E�'vn��%�b��Z���G��%�"������Jt��0U��
�S*	*Mmק|u��y��o�w�J����)d���Xc��j��Л���숁��hOuI��Rr�u�Z{�{hΐ�*�"��\cxB�G!r�r��u��kQ��[���u��E�)�+[����b�<����p�}^�����ݭ�����\"�i�k&�/6L�)��ҹ��/�y:��)�iۊp��t{���	Ǎ�vȭ�BY��=Y��4)i�'����2$�FC��7����ᄔ��a:7����{/#Dd�hy��a  �y�t�ׁ���|�{~��/*��L�o��s��g�cl�[Ս�A�K�ܚG#�<z�l��X�#�K;-wu90�����n�h�\u^�l�[�;��vʠb�J����(�sׂ|w&%ݠlc;C`t.�<��p϶���������@�}R�P�W鞫k��FM���g�UA��v�;�
�)�w����P¯;M�81�ЄЗ׮{��k��KA�,:�^5��=���_��ƹ���N��F?^�﹗�����x���$F4:g��9�H����/�O��h>��N		��
��ֵ������իiT&�}����H|&Sp|�S_!lˋd������6�-sW;n�Qs���;����'�{��	������[N�i���g�I�L[e9r�;w`�m��p֎��V��^�+zQv�J�`��z#-a���Z~�"X<���xF�No0�/�s��ݵ��C_:�UϨ��Ɵa���a-E\��(k�b�h�W˼4��y���b>���Q���͜��&!T�e ��޺����c���EOݹ��q�_�̑�Y�ƓQ>�����|�����z�ѿ|xvi�d7�
ᖲV�S^S�Oso�vA�J,Q�gM�-�t�0�K1�ɻ*��n������z��@���	�!�"�����o���~~}>��O��y�>c�
���ȫm.B|n ��@�E�}1��ٙ9��:._�i���{ݘ�a�{`38#�\؉N2�'��j}k	�v�Piǲb���
H^��hu6���}�D��W�9��+xרcҜO��>(�xwf�����	�w�Wa�be�S��[/KuP�
Rq\#�v=4.����1�0�*_C.�v��l�F-٥b�]i�����U�nQ���LU���.2	�8_�,+v,4��i�П��3��ץ����x=t�gY�P�C�p%��*��)Wy����̃�g�`��J�Iq\�6~ʢ��<D4_R�]�'�C���^CD�~ʨ
���L'��\��f�'�),h#�%<;�n�Eo+d�]ovv�`�:p匰r�" srz�5s�*E.P��V���,*�O1a6ΰ\6��i�l��F��'�=>����:X�`����
������5�1']��/ҹ���Н]�O.�F��=s���\�0^^���A߳�0q�<���^�!���ؗe7(���^f���k�͵L�➛�Sr�1G4#gSU�9r��,�Wh"<q�)f�@a��^��)��Z��������Q����@?��g��h�T[����H}T[x{=�;����ޑ�̻�;���WC�eR�\!���Pē��;Yg��E�����>~��H� "<<7���r�uY]sa�"P߆?Mk�0�;�b��A�_�9�dK��]�l�	�j����|��a��/�i�5�_��3�ᆧ�Ρ!�d5Q.�~����sW���y\�g���[�Ig���w	���<��7�ov��f8��!�T@D�4�tE�u~�xco��D�@�t�x�i���B58|�E�^��r1�fB!���Az\�+Ț�C@��t6SK���5sZ|�L�'�kO�5��Ίx�0,/�T��h���Ol�KY"�ʤ+{a[=�=����&�&�rN���N�`.7Dg�~���b;����+6{��`hG<�d�NԷ6����Ƨ%�r������2b��B�ܣ�.�zw^�=[�S[;Z-�'��^*`$(m�[�8��A���S�ff��׸2��LĄ%����Ғ�3��V�n����y��_�C�e
S3�0(�|�W��^C���Ѯ��!֧Çu
����>�x�TJ��#by�]D'���~�[�T^7+q�KY3d��Óץ�n���%vI�����R��c�f�6�m6��X���.C��L��E=j6�Wr!�uA�̚]r��t�'C�o]�l��A&oE+}�	�P�=I	Y/��B���(�'f������i�@�v��D�A˒�':ٝi��`�؎�\�Kp<���j{7!�ԫ��&�%Z*P1Ɛ��?D��"�AD#{��{����S��U?S�^o��'��M���Bt8M�fD�v�8��z_�f-p�eP��j��Y9*�{z��5+3�5Ƈ��v�����a�>�4����%���h\l�����.��#M���ې)U:.7�M�t;���3�1N7 8�#w��^p�_�LKb��.*�RP����tUnQ;*�Z���`OB���\V>��]��vC��@ACØ	�}�|��ެ�%b�����䇓P���k�W�L��%�dϧ��4��K1��Ϻ4���C���k�sy�v��/���^����e[�]OA�OӈAL㷂Q^��E�n���k*��(b�Ӗ��Q.���@!��1��ޫt��8u�ٶ������Dq��g���ͻy}�u�qE�c�o�Q��
c������ʢ�U���CL�Φh��Bi`�)�k1Bv��eHи�h+�_,�-3��aqg���X�/eT�<��9ml`�S~��Nn�ޛŬ�^�f��L���&�
9H4^�挋���X���,/���9��wg�jW�%r��F�'�,B"���q���L�W��s����m60K�E?1�j_������?=\�|�~�uX>���}Uն O��;�fěM�5@Pו��׷�����m�tV���)��ъ��\}�T��5�vZ�v��]�a���|~� "�"0"0�F#�<0���c�7���mz�Y���&�	دOqa;�&Pd�h�'�Fq�{��Z�Oʅ�IS����!��|$��.�E�xa�DA�{d!B1W5�A8%�~#4�ĥI�dGc�dS�V4�,9Z���:n�.oAt�H02B�N͐��Ɩb'�O=?D�I��Juk�S)Ż�V5�(�wқ����%��j���=���������6��N�|�vDB��0�|;��N��9�{����kh����z�	����XsQ1��>��DHh� ��9�XP� ���-*�����;�.'e���սQ����]x1i�c)�jM#���0�@~�A��;�>Ol�Ap��1h�qR�&�wl�0�.��f��-��e ��+e/a(%��A�,kc���)=v~?-z����G7�'�@C�~ʙy�t	nΞ�k��)�_�6�j�Ʀkӻ6��}�����G�l*�'��'��H�ȇoX�%�_7�E��Ʋײz}]~5\� �Z��;TҦ�����2C�uvR0g���|Bb��~mǆd��n����S��j,SF��S����7g����Uv�ȷJS�:1�CsS��$,փ�`����iK��&t��g�5g{��|��E1�ãA����x���X�O]��,n�
���JI���,87�4ּ;�l4��TnbpR�Ϯ����YE����2I��}!�@F�# $���0o{�x�vb�G�	�B3�QZ�)�ǖ-A�w���9��',���Ëd���i޹yn���y��ݔ#��#�3��y�z�������%�!8[�>�}�Y
[����T�7����Kn��e�����M�]��2��qt���ءmA��K�k�F�i��"�n.�|��[b{W>�cv���AƋ0���Pj(�3�͛e�������7��h��v��SB.���>c�� ���W}X"�}n�k�ց,���O3��xs]Wu+{p�.?~�v���0����P�r0�ky5��� �ɊN�(v����Eʶ�]�c!Ȫ@eQaMG�q�uEÚ�����k��ȸ";Ǐ��RK���)����7�-ӌ�X!`	U ��*�qv#�v=4,���H1�" �D9��.�����s����]�~���6U�7�_T��2�^b�7L�'�a.6:�s^���H܁#�v���\ζ�>���a8��0,k�q����m����m�u�`sN.iz'����� h| �Ɓ,�0�,��H��Y�_���;	Ya���n+��gy��ŠQ�j�k,�..�%]����ѱ��n�J�]J�y��׸�]x]NM�M-$��S:�w.�ol�:���@��ڪ�����Σ��wj�rc��[�N�9�^-=�{{⯁k�r�L����ի�i�u��/�wJ�'��o�v����~����}�}�������C������^��_L�ү�ft8�G�tgf�EdL��wiƪ�n;�h"Tv��9;z�����8#����tI�Ht�;Vu[
Tda(Wg���,,��%^��h��Ta���61��{�YZ���I��M�*�f�h4[p��2���dܨ�P�c�@�̇7�j�<!(��c�����1:��T��_Ƿv!�`f�r���'�k�~�ֻ:�ϧ�'�ۊȷ�P��@l�䦛P�5(>kC�a�^������ֵ�x3���f�;IJ����(�ۗ[J�C��z��5��D(��������j��A[Pt��ɪ��nDܮT����R_Y�8k�v��&b�Ow}`I�C��SVj7�zx0?vh�����w��uA5�zl�Ҿ�,�{��^�;����S�x�y�޺<~���B�'��#��1]����:T{b���'y��.w�4e�-(w[\l�+^n�
.�X�U4��+�D<JF��-��rh����N��|�7w6�\GNwl�n���kZN����D�c�q�2сbèJߦ�-pM�b���MU�!8��o�����S�<�=��"��o��ú�K�I�}]�9qγ3��h�{���՜����q{��0���=@�G��?�n�3Gvxd^wڞ����q��֤^��kc��έ�;3���V{KWm�������ѣ����7�eƃ��;'|3�8\$�JڣY蜬;w,fn��#3=�����<�W�[LS��]��ZP��n������;�Y{:�ݦ��A z5�;:>�usjic���Q������Vy�9%c���m���4�@��y\ӕCwG(\{�z�cGB��$(���{n�En�޵���Jì��X`�^;FP����u�ס��ϡK$�Z�ӱ�����f����3�Ť����i�n	Tc"W:����^�����4�O�q�&[��\a����A`��i��$l@�.�����p�Q�}̶�E�I�UI֜�K/���y�����t�Vr���A7GZ��s�����;�V�Po��zy4Ժ�pv�Rx�b�TH��ɱ��VҾ/���OiL}���n۾ПVyߊ-guQ�aW�@����f�}&E�A�x!�)�v��T'�,]������s���^|�=k׻z��m-��em��+^K�,I\6�jM��u+�u�Rc����_'�R��y���.�P����#y"��q擟 FB��[�(�Q6�����.���ԩTEQH�Rگe�l��¬��+<4p��g+eKmT�j��:Y�blea[l��0�2��l+q��*f��o.0ĕ*-j��+6������g/sK[+PXJ� �ZZZ����85������QQ�"�c<���4t�Ӈ��S�������T*#mX�:c=�����*,[Z�Ң�>��=8pC���B��h`��ж��*�V�T��-�`�ƌ
alQ��h���Â�Z4��j��)��2`����l��-YQdV�����@Ķ�m�3t\��E�R�ٳN
�T�X[J�bQ酂�e��
����)K*1H�\%�֒�<4xl�Ŋ�б�ZQm��Fږ��ŭB��[Y�L`T��V6��&Z
�4lٳ�pUF�ŨQ��ܲ��V��+Z�	[ĹJ��h��R�V[Q�0¥T�u���ҵl���f(T���V��"�c��R��&Z,*ډj"��5����������{�7���_�P�S_���i���Z��WJ+Ƴ�L`Bi�y4�pp��QfO5A�6�&)����G�����#	`A$F�DH������bV 0���=!��~��?t�I�L(�.ynnRy���cH�C�PmW�v�#*"U���;��*<���7H���Kκ�m�Y���.�TXU��e2̝�1���i5_���C)i�����B�^��[sO�(L��6m�I�:�S���չ�U�K���]��R]{69=����&��%Ә"���~������P�IfR�������}u6^w��7B���A_�?Mk�0�w��sh`Yz/a�ɑ.�8!0�e�w�h�x��W�{����{�67��wBzܤ�/^&��f����,tP�c��+�m�MS�w�ǭ�G�|�O�ۘz�RO�d�<����ѻL� ̋/;��
��3�&a�'["e��<)���g^���gm��:�خ3�:��ߐ��O�V"�Tw��~�L�/.\�gD��~�7������^l|��Jb��<�ǆ,7�'ssE��-��Ӓ��Mm~Ԥ-~�f�Y��i�,�|�����1W�D5� �p�[Ռ+&*�E3�Bli�	���q��Y.�s���^����)��ӄ�����}��.G!�yz���,<�A�;��P�S����SS͗����ԭ[��1d�@�w3���9	t^{������^�\˻v���	ƨfXSx��S�ݕ���1�m�o"A���c{��ջ�^����7��q�=��$���"0�D"��H�$0Bg��0o{�4�����M��ʛ?�f�M�8�L�F�'�G(]�Ӻ��Ob�$C� ^�0��u;q�A�LC���](U
��lƲ~BS�JuiImd�%+�v٘�V�*�/K���oɺ�����,b�f���������ОGc@BGa�	�e'X�%�u��)�y%I�8�C
i���η7{U�r��Z=!C6LB`����7v4]rbm�L�*�I���SXM��N\P.�**�/����r��Ƃ@�����'J�Z{�c�ӳ�(��'�*�r�}�m�w�G��]OL�`��+���Zq.������`e���~|��?/��y�<_ثI>�a>o��t��Gq�R���Ԫ���(#��8{܀� B5�{��:�@ܧ�6�y'��[��'k�ٶ�Ύ��H�sߊ��/j�Mܳm{��?H��t]f!<�>LdU@{Yg���윷
�f�y}6���@�bԾ{A3���S��bL`gb�Ӫ��r�mޱwq~5��5F����l�#�r}��I}Z�&+��c+ro�N!�3��FK��V�fBZ�t�$&vd5���������s���Y�ށ�9��s�u^������VP �&�*��Y�ky���X��갇k��'���[�_r^�Xrn�'^�w��t���ܪ��b�xo��3�?4����q8q�.<�:�X�Tc
���F2	$>���������כ�g����C�?��04vq.�P��0�yQ����;�7H����	����y��a
Wu�6��O����#��k�svרp��|1z�+d�q��HƉ۷A1eo4QȬӛ���{�KE]�of��E?��^Y�X�iiABi���<.�J2Rly�+���K��iҕ3e�2�6��&�Q�W��*�mO����,����>��d���;��B:=;S���;��Jl�eMhħ�(�0�z3��[�|H�D��a�s��Uo.�P�dÃC�:�l�*1W5�E���:F%���I�ad�d�u&���U�nUQ�+w嫢�L�PR��%�O9�',JBS��� nN�ן�S�����t.�+��ׅ���'���zg��Gd�P|v���%'�c
�旴�S��;"#�Y�!�^�N9{������?�����u�M�)P[\Ú��/A�<��PA�a͵1��Z�[�7n�L<�\4�Ěձ����Bn��~/��2�t�$��Kz�{`l0Q�`/q
�Q�J�_^M�J�z-2Z��󽹥�hwq��^��W�׷7^���Ev��be�l]��8�^�dl�A���k;s��ֳL�
�|t.-�UQ�\��#��e�u��v�m�窍D#s�+~64��=��U{Fo�v��}w:���V0�����	�H"HBw��=�
��\|!ᯞ���e~�����E���}�O�P�bC�q"��D}u�Ʉ���>�[���I��j`�ö>����Ȧj��I�X�d���\�8�ج�����Uʹϒ�J[�w��-(W��ń�C�y�mt^�.��#pд^��'�Yk縙����c�ϲ�U�of}s�}kmGC�,w2�'^(��g��_PY[��!徯'�R�l�.�K�wx]�l���sW���&��<(���X>~1��/40��	~���Kڸ�̣�j�kt^*A��L3���	�^�<����{8���㘮���>�8�Hlp���^a�_s#��FF��]�6�5{��i�ֿ��W캵��>�~�cW��ޘ%S��84K0��ܞ�|hnʹ��$U�A�P�h(�3״K{Z����-�L��#Y���r��3��a��P��f&1�5A	�� �EP)���rS��9nDF]�=��u���Օ����%p���ÞC*9���M?�ڹ�e�&RU���4nm\��O3�"#�	͟�_�\@-����2o���xs��ɾ��O�g�f��c�-����15��n0s~ٷ���O
<2������RW<��^rR)�6��[R̻��ΐ82l��޺3�T`��
I��>�9�7�.k޾kF�f���9|_�?FHA ���D DI$����ix��@����z�^Ʋju�����z�9q���%�
*EИI~0nDx{��[�p��o��~S�6M,m�N�S��Hеr�'~��a#�-�W�q�cL:A��U��Z�����2�ܻ`iX�@�Z��:�Ը���3����o$n@N��Q]X,�e�[d4�.<(d!��504'��52�����0].��g'�c7�P<`��\�f7c�sCγ�}��$�S>��^����?�z���]F�;I�P9+�Z�ܤ�iIA�F�.�$ʨm���{��������a���T����Xaδѡz^8�%Q`��:c��؋�Trm��o���t��B��	Ot���h&5����Oc�������﶑_�m4�l��0:��轏߼�' -�����r�xF6
PX^ȍlb;�8aC�y����.I]�3���f���D�9��f�^��a�GX%@�~�Ǵa�v�ƥ���/E�3�D�Ǹ��%�K+�j@�j�D������;7k�n�6χnR`K�}�0�uɈv���/rW�aW��q��c�<-�&*tv.�c��p��:�ո�@�G�d�>w��hM�5�:���eE��8AT'~��d���Ի�P�dLi��*����us��am�nH�o�2n�3cN�M#���M�
��O���ۥ��p�O�۾H��>��W�X�S*c*�0��	HBN��￮�����W�,<��49�'���������ú��c�'@�C׊��"b�f����UooQS��Y6��4�lP��m��ƅg�E��̔�����#s ���/���e���k�����U²{�[�B�Uy�\u:j�sC��h��)��I����X��]`NT��<:'t`Q�q�:�e�7��5��?+֮�+Q�ƍ�q�ʋ���QL|�8��9�F��5]D��fڲ�3���1�'8]1k2�ـ!2��B��70��S�=[�H��|A��]�� YX����}���Qw�1�$�K5���%��	�6�%:�%%�gI`;k;��o�s���g��7���'wCC�巃�� ���ƊEt��½�R��1,���eI*L:�+�/^Ҫ���_]l�^w1�[[��l�DH.=�r�1�J��1�+�,�`va80���ޅ�N�;#v�wv��73�f�2�Cu(4�z"k�Ɔ�j^Pͭ0D&������"I�P�Lv��v+��j��a��{2�ˬȾvOa(,`P]E�5�,����d/���==_��_{Wz\ѯ�#H����.���7dG_Z��kf���?���G�o�S�գ؛��:���U�!�\{s.�p�j}���˹̜��	��η�����I����6�3�G�+H��r�ԝr���N�g��FK<޷�ȣ������зk���	�0$���"B ��" 0��� ����8�D�)/C���
n������t	��R7]�9�I�p��y�>a����S�Z�סof����%��ҫ��:�F��&��˪`���n��y��t��9c�ުd��d�X�!k�;k�?��m�S.�Rc`2���&}8��9�h7t�l_6�(V�UQ�>��\��F}L��8>�L<��{���O�3d;od$��/�Q{jǟ��9�y<��e���l�ג~�ҕ��pXx�������_�Q���@@����+���݂��XE�^�X��W��=!��A&]�`���EC�dK< ���C�$�%�މ�餮M>T<�v�h����ds.�4�������O2���_�
��3�S���
f�RT�\X{p�vx֨���s��-�#JU�&8�Hٶ�ɬ���ޛ�ƚxX:E;���:�3YlN�Ӗ���l[-��\zU	ꡎɨ�`��)6�S��W����[�1�m�Ut��D�G�/�/�ͳ�2��b�H�	�ݲ��VY��N4��t��>�ҏҖ���>��Uٱf�r���>�06�݀���]�r|�~��o3��I?��is�ow��J�M2Fw��|�v��w����7����v���ե7V�����=�J*�A)o��Փ��a�{��֯����=��?HB~�	���J�eJ�%X«���qkƩ(���-l>��|j0"�9�SۼH02TIvl�0�.ƀFvI���:��9OV�ښ��nWJޛ[/Y�%�	�n:�L'5�4����a���	��d��v]�O!�ʣ�?\ν'�����u���p�euwy�DRr��-j�k�sP&0�y���u4c	�_����n��תz�����Y�ρz�b�mZ���8�\���A���Ri^Fi������iػ4���3��U����(r5ĈxnO��[�ݣd;�v�e��#YC�J;����Iq�΋!�ͥ�T=hf�0W�G�a�,�(s�L��C�?*���OH��4�#;�'-x�M����7���U,R�}�X@&�S�߿cċP��n`�q|�;k��.��>�4-_�Ia�Ʋץ�cDLkNR�mgu���jl�����P����6���Vύ~�-��%�>N��g�d�&�������Z�\f�İC�@:K�6�_�9j/cbL� |#����b�:�q���Qh3�m��C�y�^B�5�Ef��0�[��L�!yϭ�dJO��~^�����eI���^�q�1ׯ��ב��sތ��b��n+������d]������pM��œ`խy��T�ڽ�X�:�6���2��;�J<}q����gV��=��c�T]Lâ�[���[�����-�K�*y�=��|=�� �� Id$�F{�x]��h�\U`o:��&;�B�Q-��~ݟG�/�Gt"�TSF]�C�R|�x"e�1���$�"���B��2�k�-�=���W^�cbt��a,UG�m(� �&��������g��j��,�Sʒb��d�(�b�(Ip{�'"��j��X�'�
���x�Ai��κ�t��)��X�Xg��C��p�]��g6"S�����y򃦈u����E�i~��o��z��=�X%'����x����q�J���
e��/P�.1��-�
��L$�0�ٷ���ל̝Qk3�Rv�u!�'0�'�Ȕ��F���*�q�3�$�[GW�q�A�j��/ϡ���׌�{�:{�5��A�6�l�i2��`7H�.2	�<�,��a�_��~6k���I�u��j�C��"G:��C���2�>�n�%=_�Ͳ�ah�RP�Ƒ�,ո!��h�v�^�����e��<�m^a�n�/)���
6v�
�q�57<5Y�I�SQ��"F��������2�𿶙�4�H1��/�;��ѱ��=	y�UFě$닦L;�Y4!����JOަ8��pe�����$�2�H�xR)Yw�~��{g;j��|�4�Nۜ5	"��m�8�W�,�i�E�ʪ��_i�s�l�e�O\ڍ­����i��ܦd<��t��æ`'qY��cݝ�iI�oVS@��`�n\�m�k��.���D�R���b�����H�$��������}��/�E^=>����H#���Ɛ[�W�������@0����̮e{����1T*�h��Bi��e�W=����������V�9���$�j���b����]���.�o4ݳ9�~@L3Y�j�j�D+=/�Z��i�3ͧ�5�-@��^��K�;Nd���]Y�2Wٽ�@�<!0�<E[�hfE��j�۴X�ϗ���^��G���j�.M��Q^\��m���g�T��	�#ϡ�0��߷i�f=����)���N�6e��.�p��P��D[bE<2�����Yt���,��%�r(c��	��q�>��qYIt�	X�^܎L�;oi�橯�s��DX?|���^S������G��5y��z��������(tjypΏ�]
V
�����	���:��hBli�0Z���2\��x={���.�,��Է5?!)�ɐ�U�B�ܯ��ǒ}���3�c0
s���0v'�fu2=�ղ�*�ơ����G6�?!)���N��RX&�	*q���5���_g^%��_��8�Vj��j�A�gy{�^��Ը�k�/t�\�LM��|�콫a�}�4�[g�A�y�$k�޺;���N��H�mL��x�^��n��ɹ������jPx�8��9<�ͬ�m�*�m��(�8���"��>#�n
��R6�:Ⱥ���|��b�bz��8R�9^���V��(����T���xG{�F��}D_ :���.s�~��(���>]g�}7����~��Pr���9��O��䝛���t��=��d����,�ȷ��l\�P!���{��2�qf����1��6��E�����=�������:���۩:�l�j�A0��R��W��S�#2��UG��ɛu�<T�l+�ݶŤB��(T+N��ݗ���u�eRf��ͽĊ��v�ɨ�E^�Rv�.!ת��t�w��X3����ѣ���I�;�#�yg�e�l�����[$�ר���SBvm�-����m��41�v��-��P9�eX�Ҫ�|8d*a�.�Tsq_^���-���&��᪪Ey�Ɂ��y��n�j6��q��9�$�*�|���$�m���2v%��MޖkpڮZ�D=�to�܉�⁄b}������On�
��yT�h�2K�(��F~~��q�iS�4�r�p��3��j�FzJ�73\�}�1��w+c@�f�ӯ}g�d��aUt��~���R�:��T�ܳ��Kp ށ�V]�:v��9��v6�T���S���ӇL	vd�З7�ʼ��6.�SOUQ7�{)d�+7!��WVy������w��c�6�@�~�A����O2�0ǘ����k��[�Gu�Cw����z��{�9�Į@��5�|w|���/��\�kp�U�A�aYe�m�����S��M�:D���'4����
8��ڳ�{��U�o�y�TH��rUmJ/b���(%�����?}�9�-~^��G���y������osGy^�9�|�K�s�=�ua.x{����{�����&���	��e��|x��n��ҝm�Dp�ǭ�#Le�%ܧ�Q����Z>N�4>����MV�zd؞_������^sA�&�&:׽��'W1��0�|;V}m�)�k�ww���"�S�Y�y���0_"P����Oj�������V�o>(�r�$��\�v{^�B&k�6mf��dr7��a��L.���7}��@,���aK؀�7��K����OI�{��
a�������l�K,l�ķ�H&r��EZ�V骺x�ܡV��p�;}c�n��w�⛓=����X�^������}�^2����w��=z �]⳷��{��@(�`{O�2�Yĩ����}�j������Tv��ݨ�� �kryG�;ӧ�]g���cy�9wm�ܤ�&4.Vx�₣�F]�����jI+�-k\��VY��C�V�*#��I��F8��TQ�c�c��+xK,���������yx�W�g�N@�b��$sҜ�<P�\Q��࣑��ؾ2 �(���Z�R�"�UvԈ�+"��<<:h��p��ݳ--�*��:�d1�b�J(�
�"V*	l���B����<8\b��ID�e��R)Z�g�D}�եB�Zfc��1��9��ىr[IZ�V)_Z��٣�=8f6��B��o��[i`�[
��9J�h�ab�"3�`)���L��醏N��ajMt�Z�e��[�ZUV�˔FF�m�Ԩ+)}��E�TQ�*R�1�*9k=0�ѣӆd�Vҭ�
����8��ʊ���h�U,VUe`�eED���8pٳGLµX�j�J�ңPV�0Ĵh�ci|�1�l�EZ�D��2+����H��"�%�+X�E���F͝)(��Ed��r�Ę�[X�h�jV1�J"2��5����H�-B�.Ν:p���~s-w\�e�*Z����E��H�,���*�bm���)�ADA�6[ejTZ�"�Z^8��"ѕ�ɉƈ,����Ķ�������Z��G����\9���G���m��<ߜ&b�ړI�**ټgt��ɝ�^=�	�ɽv�O�HP�훉�8���%�t�ϰu���ɩ���)es�?to5����<�f�� �H@FI"$�"$� !!+�*��{~��k[n!�y8���Rb,�t��	�By�hvA�3��xb\��ybOEFr�
X5����n8�Z�>E���2:T5iyB����o�>����%P�#�(�`��<����.�.���噧�b��ިn�4������Ђ�li����d��U�c2�x�]�w*s�����ׯz��Y�O̓�$b�0�-iĻ葆$<H#��}���@��L�_w�q����i�߻��*�8�d�v�߉Te��w:�R;��@�^�>��-�����۾k��)w�r��8y�v=C�aBv����&��zW=����{W��w>n��`��lp�{}[�Uk� ��A�������vm���/���J����:�I�E��g�v�}"h�*؈�4#*֚V����@f~�t^�<��{�e�����d�J/ޣ���}%~�=�I������@���?n<��p�dƃ�gH����,46���ܽ�	�Ct2��4�)�y�}��sd� �
���&���o�b*�a�3U��BM��d>	{d����}���xT0q*�	�m�4��N2�E[WP�Q��\�n�9��/{��9��Cv�tU���'-���C�m�ռ�{�WH�����Nwe�%���qo�<=�����YZf$vp;0�b�/,��o6��fG����~	!�DdH#$�0��`�� <tՈ}�I+�׮��7s��(_J`h$�A
�%�<��o�C��ΖQ���*^}�����h}}��Tϯr�f=�r-�i�U�n�`Aͨ�����؍�}�o
�kvʝ70ƶ �D�rӨC���<��yq�T%V0J��W�ø�M�L�ɪњO~�^q����ؿY��(��Һ���9�=[ƪ�&8y�"
p6=����Nm�N(�<wT�ff��G��5)�G�Lv��53��D'e�X��~O�Nd|G��a��~��}ʺ��t�-���2��F�q^��|�A�%:��)�JS`��Ȧ�ȸu��i���hLpe�\����ZcW(��'8�e;ʏ\8@J�|1��n�J��0�%�؇w��d1��?�_�9_q"*~o�`�ʾ�0�SJ���>#'����0�rt���R	zҤuf�H=�m�ԣV��;ۑ;�4�T�<_YC���xe�[]4�}����"�}jF���%Λ�[tҜj��O�KO5"��>?3���Ѕ��>]�U
�(N��WN�7}���b2m��l^j���k�q{�V��+�T=N�.^wvg�t71OSM��89�w��
?S�~�$e��~�&ף!լ!��h��zLS����
-���w����Nizk{�{��ו�~zu����ͥ���r\����y�-ѭ��tkG.y�S���S��!HA�D�$�2@D#!	�>�NR2W���H)�ݙf�pF��x/R����*���M��R����Yb�m�����a����n�r�Z�]f���|�yU���:�G��A�y�����5�|�#��Q�_oE���K��um��4\s�J��6�'�,|����
ǖ��,8^������ϻ�\��l	�n�x�������&��A��e3=X&p�W��f�0]���/^�x;�r�0�s 6¬�P!̈�e5EGy:�L[e>߷g����C�I1QL�o#¡�c�bv��zo��i��<���i����"���$�������W^�cbt���1b�l���Y�1�f��g^���:�3�Ցa��_�J�y���(�TP4x2�������}b���6˖��W��8o� ��0S��au����^ʋ�4.3��0���q�1<�5���!evW\4Ql�ޛ5���C~/)��hR�*��뜺�쉇Uᑬ��"z<�Ƚ=�<�'�>���{��e�S���d$,���Ι'b𜠑�j	I�5t��	�m��{h���^?�f���^�>�-��tZE`o��t��g�!rO&'����������Bݻ���y�A�k�-�Ǿ���y��x�y�=�>�H���<��i\À�ڣ��:�㠋�hr��2���O>+�.����ϋۇ\�}���^�S�� �a"2 � � ��s��4Ｍ�hr�����Fܻr�=����l^�e��&]a�E'K��@�8]�M�Fn�f�Wv����1�#D:	��0��˰�6�T��c��"�Ect�1�����|l���!h��#��#�i\�6h�_~k��/�S����!���L*�rW<�G(fGaS7�1N��y��^��K���}킡����(��ш3�7;��߀��u@uoc���Qrλ:7�G޺D��1,*�O2��i7����O��A�:z�Zx����pgÁȺ�n{��X�M!��s�{f%k��_�s�� F����*s�;CJ�LR��T���wۿ�[�@{�釰2$:��pB�T3Β�X�R9'�{�4�5-�G�Yr�ͳ���!�s,J��Wb�t�!��m��g��ݖ��#�(�%�A��1�&!��7=]�C��٪����b���l��.A��˚�|�՟��۴H��E��WO��8t�;I74��{����n�����FDM���:3�
�{.3m_��#)a�]���\�����MD���k|���6)�DBP8*n�b��B4W#>���|2�h�Z�;�Kg�讅t��@��W/��}�zOW�M�%�-��K\Fl���DGh���v#)b�9]���jN�q�wTԞ�\��.>�g0|)��L�nc�p[�!?$D�# F "D�#$��&�������Ͽ;�[������yo��	��܄("h8g�.6�5t�ê�x�, Xt�=�I+ͮ&H��Ӫ�g�k���q�;�cد�U��Jʣ����sƆĳ��[�p�Wj���CZ���$9�^�A�]s�Y�;R���D��`&G֍
O`J+Gw�6u�umצ_x�1�N����d��i��˩	��mE~�d��u�I`��%B�R�5���F���v��ŉ�?!��>���g��Cp�����D��1,[v+o�U��Y���z��QiVU&�ؾqOw0�[[�
&����z/݅���e���(�=�������5��E�K-��|��>�l��B�MN��;���� ���78�^���>������0c�v�UU��,ŧ洠�]�0�s���y������jF��~^��/�
�5��Gu!f��<�(�VT��NH�%��i��I
�w:�ť��܀��[7���\d3���R����G��)�zb[:�h���`��`:V?'�z�*�A��m�m�ؖ�CwEM]����l^�i�R��־a1c��
�p��]E��fEfY��'��{�ȰPu�`�ѳ�s(Q���Ƅ�nh��-��j�a�(�V����c��v�%S�t��UjKD�	�}{�hKSkDMל����|�����{ݟ��#$D�D � �!!7ߞ���~��>�
� �a04>򁣫�'mN_M���I�����c�o9���,rY�z��n�L�L�?���;�	��<�ǴB/"u�P��y>f���3��)ύ�u�w����1�Yu��W�lZ��;xwA�e�B�e�#��VZ�cF≋���V�Z�`� �"�"�Ӵ��-���ב$<H_���
�������5��:�앹،hPծ���֝�0)�o�����WH2�2����'�sͼ4��>��6�F3�̆�=k\�N��G7�FFp�*��_q�jJ���A�SlQG(=fͧi�~y�/����9Ù������q�Þyq���%���h&��aLm���c_.g���W�m��Z��*2����$�p0}Ct`!�*60�հ�F*��A8���TРC��f�+'Gv��δӭ�>�V%*Mw���9Y_*6���>+țk��c�r���Hs��]�1�ƙ�v��q����%:���e^IRkk�w�Q�p�G�@0*���GRbs�m:�y�f#�f�,<'�V6�˸,��O(u0�y��S��Y��wXgfb�����Kт�F���2�������!.[��*��Y~��{�Os�X��IHA����~��͌��X�av��@��|�8"��d��n;�\Ov����(�
��I���C߿>3�k�N�5�.��8c���{�Q��Bb�7H�
��a�@���"#����gNo:���6тk�W�9ljcC)�$�v���,��zOȲ��9�F�=4øvҋ0~ۻӋv{A�c��ÜH�,u�z%���=�ߗ@�/WJS3(zJ;��\Ӎz�Ӄ�E���pg�b�L�|94�����x1�Cr��{� ��|�=ϥ����gػ.Rs9 }�de{M׹ۧ������>���e{b�ٰ���t���[���ܪ-87=|���d�~R^?:�7)��~���`�X_��޲��<Q���Y�yїT�]Us�Gp��c�m�������C�Z>��>V���a!�/C�;=T�S=.ﶪ\LB�s��Am�Wk��dkv�k����<�D�f-$�w�/�tz�>CZ�&O�OW�c��k�Gt(m���� ��h�r������Ϣ���Wt��@�4�2�9f�4�����YWK��n�X�o`3XHfC<>عa�M
n/����o��nO���>9�A6�}���K"4�?j����׌GEXA6��Dr��X�8�~�8?��o�����>���|�(�#�|���"�(UJ'7dN�R��v�}3:��s�����CR��˹���ۜa+x�����CM�V��y��_|���}�����Dd��D"$�Ȍ���{߷����~{ѕR�)�}��!�٦5�-�?rf��Ј�
d�P�iu`���U���{�(/]t�U�^���^݂ըȣ6��K�B���`����nXs�F�#^�n���s�8�٘�z�72��OA� ��0�P�hRS%����h�j�����M���0s�+:�z�g�]��"DJ�&+]��v:nm�"��%:��A���Rqo�l3Ϲ6л�Bs����}՝���h0�|���m���:D��T�p�%���.2�3�+r������̾���JF�g�x �UX�)���!�4��˱R�v�c߸ǩ�uV��9����+-�)S�,3.���_�C�+����aў}���P�Mݞ2$�;J\U��ݚ��ˎ֌����fז^̹���+��	��F�Ɉy�6�^�	��ztE'��N��ɰ��'%�s>��-NN닲�k���u�D֑^
��9R��a�B�*�Sf�!��LNr��[�A��{+�Z�I��zW0{ �%�?0Ӵ'Z�Z]0Em�����۟\L���9��8���`��)gQu��vo3����n�&��T�fS>SEb��{޹Z�D�Uٲf����D��٥�1�n��8h\zm��.,pWw2�/���QK#��l�����WM���+�-K�uۃ9Y<�躉��i��V�|���t�.����d�DB"A��F�燚�߿?:{}�ֵ8��B��q{��s��LP�J���J�b��+�P��!^^�ݾr������ǥ��<�R0N� ���������1O9�͓��Q`ND��L3v�� Z�����]�����7�4��5p,����5 �г�5>VEN�ް��J��u�b�t��+����d�x/�X�3���{��'�_�`�c�H>����&e�K��_�]r�<�b���^�͖���\�x��
��K{K�]�5B���?����p\���qd��0��Q�u|��YR��4�^�A�WA�>�4M����s�,ݑ�Yn�_���
k[OXB��=2�8��όON԰�"Y0�F�'��G(P=��)�sy��ά���{i�ئ�\K[�D_�*��~S� ?!,�&%:���M�d�,�v7��ދa�]��-�c��S1|h�,�i@G�[_x>P�	<�ƀD��^�锝qQX����mOOSӽGMR֚u�ƒT�S�_8�=��}ab�3\�&^���.�B�q��4M~�����f�8�i�*uxr
�
­�qo�mSb��*���Kk��K;�N�z�*�>9�-�4㧺��~��c
IB�l<"RǹW�Zފ�|/1U�o;�<���:Y�)��ܟ'<|=�C]���T)��7�ܛ��o��w��:u��y?H~	��FDIs�������o��k�~�dW?0��J.��)��z�Q�� �0m|w�@�0�>M���+�+�+͘c�ol�B�л�������_�E��I�I��'�;`>��tj5ې�1�3l9�]�}�;kLp�gg�+�S�;V�d�2�j5�P	P�z sIzp�Ƭ³�-�mծ��X����@p�N��ثӴ)�{���W���r���uN*���n5Lf9�����6X]8�̅!�\HCh��ً�����6���4:�Ƨޮ�����6�M��vW�^/�{^��
�*��(h��5��i�'��!n���{3��F��y����!r�� zq_�񿲳�U��N�-
���ōq)�ง�W��Jq��s�m0��u}��>�~�,��>������	�4� �o�b*�"Y�е�R�&㵶�k��,&�)d!��<5U�mnףٖi�(wO�UJ�{����T;��T����9���m$��.��n+Z��`�i��ޠ�LPw���:�=��|z䲙�� Ĩ�	�r���(xU)vt��*�v�7P��]�{ÏFE�/F�C�0v�Q~��t�����ײn�\>���c�)=�{�S�+�8q��rK���cK��u��Ʒ��B�|�̗����1�sg��h��������Og4��q��8ִ��7��tP�=���}YhE�;�_t�6����o)�Z]ŝ��Y�5��0ǻ��;�d����9�vt	�C��ynW�=�h)T���C*��%6��V���/��nڛB�64�6"l����Y[�ŧ��s~�����r��;3r9��0������;�2y������2�2�ӘK�&%OF�O�S;I��}�{��X�^��`�� ��K���h�D�S��]��Oeև���s��%u�w�u��+{^[hEp�#�5�9��D��=~��a�]��jzEn3F�mؓgU�#�*q�gq�Z�I��E���"��=d�3ڮ5�tZ����-�	���3ja�ײ��m�֑�]5�dVVY>�b3��M�|�{<=3F�^�4Uܮ^�n��]fm�d��A�KG[�@���h\�t�·�����3�h�,�Mg��`���\�{�N�zH�yd�TMC k=	�v�}���W�ëv'�=���Ƹ�j(�f���LOvFQ=�漺Ғg+�k��퇰�Ǿ����V�k�If�]s6�Oh��C��;�`=.�w;������(�6&��'��_Ǝ��?zXi�p��ً �ƕ��'|�K!�BF�_z��rG���6�P~���o }OmG�)nk!uox�dU{ۚ׊B�lӁh�x�0�*���v6�[8���<rﶰ�S�wp��v��@����w9�ȉ��v5��u�1Ƿ��{�:_D�.���OQ���t��G`��Ŏ3y��d�"���Ci3ktrԈ���5��&7|�G-��w���c���r�.��4þ�\9�|���J����y�;q����Zy9,f��ȅiu���^�C[
ve���S\��U���oK�<Y��jB��9#�I<��l4���+����;��z4g.wO3�T����1���#�c�:�x����]ugE���K\��'9�0�'�I�x�cNy��;$ћs��uW;dʏ^L�:e�;Ҳ�����u�e�G%UA\�}��������<=^0{qf�5���B��JM�/-'�p��Ϲ�t�'<o�Z~w�F��}�<���=�Y�,G1�~=٥�t����2�ލ�]Z�SnŞ��O��-�Ѹ�cv���.�=�H�r��)�AۆZVE�pw:�ךO<!���x��B�ysc�v�����7���jN��jXF��ܻ�� ��t�/llm�n��KM�-3�����SC�Wum�u+�=D=�Q��a���;���-�w�C,L�?���R	�`�XV+"ȰY_2������cD�Ū����
p���f�b0_YDSm�eeKl�6�+%kU-�*)Qb�������Â)(-�jPm���_)W,%fe���a�m닃@XQ+ӧO�9V6�[j�������(�-�b5�ȫH��l��8t��g��TA��>Xb1"�)l*��)+X�'�2�mi9�aNYF*�t�Ç��m�U
��E�d�QB"�[md��Uq��W-m�qĞ<8l�\��.1�)[��
��T�*U��۫Fc+*,�U$��X�xl�������]0Ҥ�
�-Aƞ�P\B�9�(hˌ�D�p�X���PQ=>>>4l�ԉl�R�bŪ��UH-ejyn6�U@T��l���+PYm�T�M�!���BV����+� c4���
ʕX��������urGg�[؎U��U�V
�}�Y��5�u_-���\c\L���|�-��#}Z
� e��{��mkO�O���$D ���<kk�R��S^�Y��l��ȧx���,9/1q�B�`M�E{S!5�2�&m�nU�31�*��w\)�\;Mk\��Ui����~-8�D�:���ܶGP�U�n�j�T��su\�]�{CAѮt@�X���i��R�T������=�ă<��]za0K�#M3��:�:Z�":z��曦C����vN�'�1)ե"�PIRkg끃�.s��qM{��:�ʴC�O�]LW9R��=��hl�r��OC�ny2��1	��7N��a*,RQ��>@`�͕��tz6!f]�ic?���cBa���/C�L4�nY'%�? �k!����ih���F�%����ְ���a�
5�r9��k��Kv��P@�y�Y��C�餓�>��}�ߕm��k����H|�HⲈ�cg�ܠk�ީ,hV��'AF�U��kS,�s�ڭ�庲^�5�iy@+���UA�5�D� ��?�yO����=�_�bؼu����*�)e�F�Z�5���z}Tfu�#�,?��ۯ$DA�W�_�=�+�9�����>��[C)�\;a�j+�Eؑ�k���&)��m��7�AGyF��3h�����{M��������żOmk77�+�K�9�������`�&fs*G$M��1ʬ��&�qc�F�{�;������Ns�;�����>2"D`��Ȍ���>��~~_��?�폲������N		�i�qhhy���V�l`��[7&��ڵKŇ���{ǲ�Y�F)��O�&��cd6���@]���1f�d��:"�q:��8���E���5k>+�vM!�ޔ�|��7����ٗ�<�]��HA��/�����cs�]��e��/tT��r׎�)�lk�pB-���E�j=7�6�j	���V�d;�B���U7	8�����`6��2�Ο=;Ǭ��<��%���W�n`1�S*�P����u���הi��O��΂sj���c=x�!�(eEîp͢�Z(Eq��S�3#73zL˲�ɟs�~�$:ǂa2�Z1B��W��_��0�S���e'����n��s�16wpZ�Y#��v�nHB{$����2/��Jt���)I�؍�atC�oCK��&��Pz�'w���-xη�C�F�A�Ĉ�C�ݗn nl�ҩ2��%~n�I�n�Y��l�X��Xr畵O���D�&E�2��i����?яy�,���Xz�)�j�͉w�t�3a�u���hŬ�ˠr���F{S��Z���w�V��¦۬�q��`��x~�r���d�|��F����2���}�w��k%O1�;q{b;D�}u��ft!��n�`|����NF��Nuu��iŽ�ߚ�]��?���j������"QE������f��q���. -oe����E�m.��q��������.wbK���U����J��O+Ew,ں=�ݒ�
^��/-B��HF:�Ƃ�P�E��q#dlƽ8q�M�"m���4�;\�CP{�R�j�w�=�l�Kek��Uk�}��
�����Θ*Ai�^+���I�y�F�������^pcZ�pH�Y�"��q� OJ�)�zhO�;Bu�{w�t�v��֏S��#�0B�4��� >k�;2�u���	�f�@�O�Z踌�0�Ы�l�+�58&U�MHf/�+��\<�k���'��k��?�v���,bK�3]�B�4t��t��m&k��:"�s�gO����"B����О-ŉ��J�i��8�*C�Ά�+��Y7��ѹ��@!��0�����:L�c���|���N��t䕹�^����$��*?~�x`̄�Լ_A/�r�$k�"�kΚ�K���
`X|@v��=������zp��I�U@��0��������dm]�T��{Sl.aΎ*ޜBa5��������2��dXS�g	c.�g+���l�0��%n"6r����K�癬��{h��
w\����#!��)_5{|��q��U;]ͭ��jv*wS�k<�P�*�y���w����u�)]9z�GX8�l��v��C�� �<�n�(������4y��\Jy�(�J�;R�G��%6H&BeV�
R"�H��־�^s�6Nը=��x�����|gh!E���1�@�!��O5?!)�Q3I�s0�m*�.�Os��H�����1P�eyOԭ(��'D>P�	?c?1;��~3�=�^uF�D���x��bY'��˒T�PZw�H�Ǚ6�|����@�>�.��}����k6�)�Kͻq���S�ʥ0,���M��;�7��r���]��|��`���P��nxE������SJi�m�s�R�v�8��u=�1i�X�d��#;��"�}����A`Ww����󳓻58e�L74�0֟C�{�6�[Wj�`��׭Dk���祐#��CI��L��&��sR.zT`|����h/j��9�~�ȫ�=V�w(Z�
�^��#���C#��k.�9NB��ҋ`�}��p�7�����[��g�����6�ij����Ƴ�k׏�{�&~�T'��	�h��J/~���.��E�LR�k6����T�s�w�e4��et�L1�*�+-�԰hNx֨�叧"�"w�o�������ul����l>Y;�q),���$���E��;:��=5�}��7Jx<�o���4�ѯ�-��#��[��&�ى�}���د� �g�\�J��_L�e���vN��������ew:��^�0���G�K����yn/5ՇX�f�`͝���T]	t�׷h6����wB!� M;I}����~��,�Z�*Z�L%�9��6�P�D?2OR�oF��z=�f�������`zK����u{G�D��Y[s'�Օ�4��Bޙ�斐��1|����[�m#RT�e�o��S�ԭ(�z�-i�";;5h�?d_=�3���Ë�G�:.����.-�6��y�)�Jq|5�T��⤫#�J����$� ��`y��-��D���̆�u���0(F=�O��A�Y�7�􎡟j���X��q��W�ĲOi��Ͼ�J����P��e|��i1�c�	ٮ���\��kle'�ݽΥ*�R�i �%sן��Oa�Jua)ʼ�����'ݑhL=�]��6�k�>�OG��d!����>�wd�����q>&�+P�!1V�"�	I��k&7��||S�z��gj�����C#G�"<�9m��۾ܑ,v(�Q���1i�`e#���$���,Io�ᷕɰal�{��1.oر�I�h���3^�.�����ns.�uv�a����/�o�^�l`ѓ�xq�cX��LO@�q{���x��C��{2��:��#bR�.UJ��5��f�)﷦j���8�7����W�ٚa5�H���~U�P'���ߥ.lvC��a+�?y�O5C����k���7X�T*�J皍����<=�5�g'o8�E���)��K㸀^/�X�1���_r�|{��j���0Z��kD�������{��gR��qD�|�TՆ7�Q���k�x���z}����ි'���,���u��b5]H�No2����/K�a��<k-~<�N��g,��M���T��Ar���˾�y�K	���/C����_3p��풜i�i�xqhh�E�(Ab�?�6�[�t��zѻ���|,=(���X��Fp���,B�:���^C[&UJ�euQ��lUЯc#.����qns�XW �T<M!��"�H5F�^ݏ]�H�ӄǚ%1(�@���UVA8z��za�����{�m���fq���B-�=Ų/yy~��m�isϓA83��7��W�4���=�t�\Xm(�i�v6��|��ʒ`X�����b���8~�:�OgER�0��R�%��wBO�xa�0"��>��f@�����a�����sp/O��:\�[�m��^��m�����W��;��&�)�����ڂ���<�Պ�O]o�m"��� �y� ;�ۛ%~[�ߘ-�����x/,^�`�}�-{э��} ًV����ʁ!g��}��^�7}O�y������,�A�=`����!t�I���W��AEE�zsw����������?���������*\�ج	�F�%>��[A�n��x[�Y�a]�����ڡ�{[z:6G�T�S��@�;4����D�x��\�PU
Rqx���8]�"vg2�^v>9�Ԣ�:��?�+/�����B5�~�qX\�1�ҩ2,�2H��Jݴ�m��t�q7�z_B��6+T+��|���[1��"'��ǵ�w�q��P��v�J\����=��\�9���f�݊nN�`��ϸ��Εʂ@�xwAP>�C,xd�M- ��U��ۋ��n�0�%s�U�)<���"�*�S�:q�Q5��g���_R����3�;��;M���~�F��vN�`�
��d���uk	�{mi�W��3��4�EBlm,h[���פ�\ڼ��qq��L����`bN8�OJ粠���J�a>;Bw�;T�<���M\���W�w�p�C��p�-"�y�fW"���	�ǩP6�ֽ�y��u���Ƶw[�LZ��Y�/���,��d3p.C�&�]����Ǝv_��>�&��@�_�������������}=�t���̈́֕��t���ks_�w�>�r]��iv@�TkLе6��?��8�=~�V�{fU���9�R=Vz��w��w:9��t�uU�[	�9l:��K.�an�G{*�_�� H �x0a�7���It�G&����3-z ��'D[qL�����4>r�VE�f���˞�+i���6�8�o۩��f�z'Z+ǽ��!�O@0�A/�8f'I��	�>b9��}}Hc�ӗ�qu1�u�zǦX��dw���E諐�M	g{��W�=�FC�C:�F����P{�(�4��َ�']U@��ʖ��j2�� ʅ���'=ٶA[�I��4��ȭ��޼������I� ,�,y韚�����6�=�D��	��b2%;D^��=:���3/�������PUi�J�/G���'�zk�	��7Z�d�Bh��d��/W_'�0oo���!����GƄ$���F�c�m�'�|��3��j`b�a���Q�ȴ1�$���{;��3g�Q���K$��)�$�0�ؾqA��0�����3\�#�p���s�-��SZ�P��o3�:��T�-��b��]0�U(��7E2���u `�f�{w���w�4��Yƃ�m]ڸ2f9m���R7
Vv�88�GN�1���$��a��8��h����զo��ݛV�Z했���OD�`�G��	]S>��~ʳ|��GYZ�'��ad�6��u��49�ڊZ�T���[OTzӽ��Q4i��w�M�`��>���㲒1�K0��}����L������<��9���o�7��Oш)U�V	(���@a���4_��K͍"4F��x/@߼6�sP�[B�UzՐ�̪��]�f��3�u��WQ�i��6�}�+����5�A/�u1�Q
ghE:���a]�W9Ʀ;�\����0���GmD�T�e{b�-�>C~{��<�Ɖ�Pe���=�1�:�b�T�����5����ޟ����x���`��)�V�v$�E��K�c�0yO�.�{y���o�K�^���I��^=-#y�E!ϐ�_T�P�i�'>����n����On��ڛ��P�D>s�j���۰�B;���h{��A��# ��k��鮛�]*��U�����ҵ���M0�Y'�zamF�k������*�2���Y��鈳�}��T^�����إ��*-`o��a_�ϓ��S��[��q�*f�Y�%̵�mNܕ3���sW�z����m���6_���N�Hc`j:��lx[�)������V�E��J�Ƚ��
����'�N��a�N��ǬxOt��P3��D��14���9S�3�HW����R�wO���)����Z��M�v�U����A���+hgN!�Bb��f��%��o0f������ǇR��۱(��j��}��CAR�ӗB1ۜ"fe�Iw܎rT��.#k1�28��%잾�h��#��E�؍gg^cOm=�0`g��J�rx3=\���a���I��h5l�Ү�P
;hV,+�?ZĜ�'xŴ�ZR�ݥΞhp���u�@C �.v�L���ґL�%I��nP�{�R����^�4�ww���c�D��^�μ<���Ζgp�2هa�7'�����$��Bb�7zE*J��5���0�^l���r�:��e��y�Ű��G��M����^�-��S���Ju�۵���K*66���w�	d��ms�L'ú���a!=05��1L����W�ݿA>�;x��s�j�ݺ=و.ǩ�9�= �	�{��R�I�V[A��6~!}��=�ꞵ��V�8�u�+h���m�G,��ޔgj��q��W���O!
��3��J$�r �(.#A�G��x�3�*{�c5�}��	��	|n�,��Ė^/_�]}=3��f:�!\�4�EO���cg-wl���2�	����_�'���ool$����K)7L/���sP/���V���W3�3����F����D�|�8s�o�sC����ןv�D�4�@�f,@@{�ʜ��G���;+��9y���_�eW�.ֽ�zl�SFg�6�B�tu֪��1��B�̓����1b���C�Kj��`S#���wT���U|/4�n�A ���[;�PE�Aʽ˅;ãE��*��{Ք�J;.�0�-�+�ea�ݎ�[zGs�1�x,�z;��b5�86CFA�u	���嶷n|TL-Ķ�����r�!���k:ˆ�xRnK�6�F�=��.7��;��9�Xq��ŭo�c�_f�O����P��p��K�`��<f�v�͡}�D7ڼrOHf�@P(�7�t\n�Ϫ�/���#�FŔ�+D��e���y��,�K&��qڧ����Er��6�[垾��^VP;��<�A�[S�6o#hdo�Ø�>��ƕn�K�k�*�솶-cG����w� �w�{��N'�N�kiU]p�r�8�nҠ��w����*��7u�gsՂ�˸����
��h?W��2�^܊�;i��Wvy�m�ɛh�RoBn���ĭ�����p�7΂�'(5L���R~�P�Iמ˹�F��$�n��������z�[�#��w-��:�bB�섮9<��-#�S~�G���a#�U���y&0VNHm�Q�魯�q�qc������[�5��Ƙ��f��e��&^ICg�5F7=�G�J�ڪ�G�{3%r���Kۻw���4Q�0�'��3帒���Voz�z��в11=䎶����H#�o��<��mU�_&�2�X�wM0����oOә~�/y�CW7�
x��5���Wuۦ�Y[U��śn��yj�;�Q��w-�ܭB��ӄ����Ƌ�y-����
�e>�LtsNeU�#{Vo+Gv�q���RY�^��芮���q���C/�N�JT�o@�X{���~��
��D��K���)�@��y�2��Z�*qM6�WK�f`�Q�!b|5p�y���=��v]��"RL�z��!��pco`�!���u�]�?>Og��r1��B�p3���_"��J�"޾���}q����Pg�O
��\�x����
ȴ�X=��z݌%�����֨�˒����u��8	�W����W,��\A�/k4���=���������9'��(H���Gǵ�@�Mˣ[|6��D�,��5{}i�^=UxߵRx���$�G�x��I8�stj��,=�\�����6���l$���ё@�j|�vf�+%�4�O��>t��NP��w�#ͯT�^�~���;|��m��ٽ���+��җv��{L�x^�V�T�If�l��*	j$��p.J�4������u��16���ݎ�&U;����]���x���N�^F ҫJ�UI��[�:f:,6�EӼ��VA�۹�=&v��B �R��}��Ry^7�zv�t�H�o#�Gd�V*�f����;��w�^���a�S���ʫ,T��	iȶ5��o53Z�7���ʠ�N���%��<LL�i@Z�%�Uk+%�E�"�Ԃ�3-!����ٳ��Q�QV�m�*-kP�I�vj�(�Y_P*��]+�hAa�a������Æ���L`, ����̰F��[iP��D`�ek�X�0��Ç�Iơ�K��d[Z�Ū���a>�4��P��&56EY�E��,����Ӈ#`)�*�ì��±AA��"c[A�T�Qkr��N�@�dY�OOO!�Pk`�;i��%H��3-L�q%IP����3�.�b�xԚ��`b��J��#������6xp�����V^P�,�����5ER��J�(��X-VACv��%X.��<8r�b�"�Ud���lm�"�-��&�9�+jAm���ATF6��J��ե4p�Ç �hW�2�J��娠�@� 1Am�$U���d�����Xň����5,����(�W-�ZB�#hV[W���@����_Y�(�F���[�or>�<�O�ݲ�N^�����	^���<�v�o��N�;�Mj�b�L�x��bo�uU�vj���:���i�<4�hP�mn��j���^���T
7��=��q\U=K;<=��q:���?�b1��A�0[�|���^���O�o�~@_gtŐyR��ry��,���Lp?~�z3<��ʹKOհ�"�1|�°���uW?Wx��k�gS�mn�Vu���i*�b�U�@�!��i�tgO�.�`���9�\�L6f�qyy��C��!+Y>�ka'���0Lm@�T
5����x\���5��sv_)mʹ}�'��hZ�n&�Όb�����X�i�2�dJR�&�ru�%�Y��披�j�|W���t1��o0.��)T?l8����� �//��N�%`�Y��QtDH-ަ��2�F/����#�:~��@�4>_|��K��{nb�F�H��T�D�<EuF:�Z�9���:������Q��@��I�L�3c���?<��c��]�mT�hG����:s�\j�^���{=Ⱥ��P�ZG#bh��~g��{h���C��δU��Ǖ�F�캛�[̥�{/�V��L*�rR)�b|�O!'���<��7��]�v���p�&J��XY�`7NY�h|~f1��cwpn��z()9L;��w���?u�L�ב"6�&2s����e�"�t�j���Z���ˍw}�@�C*P�����h��Ʉ��=�ˤ���T��w ��KK��M���%V.i�撞Sx�Y�:��7g�d��i�����(UT����U�e`N���[q�K�F���vN���,(Z��S`R�a>/m�<���c>1b�p/���Xs����9c!��W�t&ʘ�"����$�'�sߊ�^�Ĩ�*z(U2���r���S}��2�]����̇9k�����]W0-C�)�;G�t־t�kM��̩9}��ihlԺ�2.'��e����(4?�i���2�?Fxݲ�HZ����&�=gi����C/-�Ǡ�3zfD��c=���C������)�+��k�ʅL�w�����N���ϻ�`�I�i���TL���<�U㗳���(e|<c��]R~�G�W?w�����a���|�	zd�d)^A��=om]1ms���_���3��V�����2���iqqw5�b�����)|=�e�U!o����mtkO3@ך����������|7/��ǩ�����C�G<�1��P'jXOqv��L�y1��c�u�����G�7O��G���r�L4�3���L&�!���|Cu��{�W$^�q��t7�Cj����˾)W+ί��52�yW_!�i�]D�������֗_a���Q��g�z�#��l���k��~{���#���r�eG]���ń�a�.��]j�jP:�j�9g5���W�Z7�w�g���S��`� fެ��sK�1��*K�!%B�6sZ��<�����1���tL�[~g0î��[sU�o]2�T��%2���9��:O!�7RJ�
~��a给��p��j�����vA��|��D��]z^�d�i
Gd�y�E�L&t���PZhux��-O"���Qq:(r��0��zU�i�a��pnu
��m|�{>�w���I�x�I��{�.���=LE��
�)o�?�¸C���B��M8���'U���;Vл �i�Z�eZ�����h����7N�۠/ Aw	�����#�ؿ��Pg\�&%�y�ѱl�l+d��Voj�E��˛S�۶�&��}�}t ��pek�M��@�a�.���5��%��ރ����\]��Z�dVҦ���'��j}�gӯ^���uC�ʁG��N�AO����^ϟ}b^��W"�����Fr�c8��sq�����7�u������9��).��j6X��SϷ>�>�>N'�;7����ݠg������	^�"�&�]�}�졔�䋎��t���q]�ֳ^�-]B+���Q5�0��e�ݾ�E�3>Σ:M�"k�y[~�4�:�@];�A]�y�b��s���m݆�>q�=ۦ���w����[R�������U�ݙ8�Hv?���Z^�9�eͧ��\/�mnbmoT���s=}����_����(��'?5�'�:��k����q,�� qͰ��$��o+��^̳";���.U�C0ÜW7���D����u��p��/4S�cC>X�ib�qi���}<��ө*f�1���Q5���u��8x�C0�Ʊ�mF�=�Rv=��"���8A�D�oF��jL��Z)�3:Q����e����^C����eMV�ӽy#8Fc�V�F;38��\��K�ot�[Kv+�u�#	�$�A���U���� ���?$f�_�*AG0��\�Ξ}O��4��f��������F���\�4W0�ӭ8�e[��Y+�s!BJ�IJǶ>��+
~��^�}��Zn�r�����a)f�~�;r��rz&�SI9wLV��bOE(NJ���]\���יww������'XO�B��Lp�m�1��}�0�^ �S#�)x�!JOO�zs_0������z�dsN'/#gǦ�8m#�M�y��|����X3����T���N併�wJ��9ݓ�R��/4�	�=%�^O���%+(��!��ܔ_�k�KiuFx���Z8v!�uʷi.ls����ˮ�V?�ϟ��<�{2�,{�N�[ts�p#��]��+R�ד�g4m ���u?Q��s��M�R���ɬC} F�k��Ow��W��j(��H��}*�,�]��=3��W�jȮ��{ܘ�f��m�A]}v,wM��~��"�5��ߚo��???y��H���yy����k��|���=����z����"X���W��<=
d=�^�ˡ����6O�:���[[���[�_�G����j�a�>��n�rc1�3\�����ɃH`�C�T��[Зd�;��׻e'�1t�E[2��/�\O9͚�ʩ|�K8Y���`H?��p�<�,�	��sC��ݻA��
ė��3ů-��%Ouunf���6~�|����������ȗq-.9��0�ȯM*���t���8}Yö+Z��T��ʾ7�(B$�j*B(����Zz�<���l���	��h{�	���L^[�0��)��V{��j[qe!#��4Q���ɄC��Ǚ�xz�����h2�WM=�O}�����v��FEN����3EJ�e@:�M�D����ŝD�s��3}��c�'CD�
)��a�F���J8(��yV�M6�h�c��5�4�6i�M<zi�G"��(�t8N��m)�R��P�2����?h��[.̫5������:���b��Pu�b�j�](�sZVwQ�������_����vX�=~��TE�4��ۉ(����������V�Ag��!ݣIm[��Q�aT:D��91ӛ���|�صt��e.��j��L-H��GfD�p�7����:��/%1�y�0��S;��F����:�7JЗ�ml����Nc���`F�N��ȶ޸iYW��I�ݼt�J��+�Ըb�==�a�EH@�jt�N�18�/��nS�?P� ў�!����ª��â}F�K���u+��km�t�yJ[V[ݴ�C>Y�ޠ�/0]�1W�ģ�vX;�ހv��W*[� �u}����+<̶�������y�B��}(��� ^�*�r{V���Y�ku'�Q�j�n��2{
���}w#���9�2° +��ػR1�'0U>=���"^_/f�����Th`pa��v$LM�cBɞ�[�yc&��N�b9mGjʤd��& v
��nyڇ��>c���|BҚ�fcU��L�O�â��^�hm[�!縑�H�Ĵ���<#���K 1�ѷU19AX��ˋ�o�O�c;��.��r�͝vM�<v�<0�����R�{�1��PL�{W�^�c���E��ǌXy�-���7]n�n�:O�n��j�����܁��D'Z��ꍣ��v�UOm����%,��d�y{T�V�v'�`3樰��'^������3S�fe	���g�� �)v��8��\����=�3f��ӈ��P�@�}b
��r��,��Eo������j��=���J3H��x��g�^�Ne%�u#��E=m�:��R�ȏb
�md=FNc,�x͞�m-**��PMώ��4�E[?�7Y81����x�]���s��x~��;�^��/��; ��#J�V�J�>]��g���8�ݓ��w�ӽ�1r{����OGI�l�C|Kҥ!�%Ak�rn���8\��u `�~��g�y�˶J���{��	Ѵƶ��di�hi��ű�48e$��sZa��A�j��[ݸ��e�с�[1Ǥvv\`��ѽtuHH���b^'r9^���Cf�o+6I�xfh��5J�}`0Y�#�3Cd�]�j�(�Fu<�Ƶ��x��u��{�re��f����4��m���`à���Ϸ���׾���b��i��~}�~پ����f�z�+駋ًs X�<���%��K05����oZ��8���AmL�;�ᣝ��%�t�R��;2��kR�K{�W �Ԅ���L�#��8���4�ʳ�\�5t�z���k5�G���A�[�Vgw�;[�}�������"(�2_~��6>��Uo~|ڏqD�)؊9A>��#��1���h-���m���%T��De]ee�}χ%�7�A��s���̆�U0xl�gS�q��CG�V��so >`�+(�O�����Lt��̚�o!ښuA�;r��t����*��~�}�c� ��&���+��K/m�ޕ6no�����t�y��B�]���TUɯn8u�� ����=�
�L�n�����v<��==�?���F���Ǎ	���˙W���^��|�ʺ;�k�d��3��4��4��R.����F���0�R�]��rl*���S1�}�y�Y �'$�#��3(D�6, �Y��ڂanD�q��d2\�3Dx��/ke����I]�Fd�ۉ�n�)f>z���N��}�ɜ���fV)��ʑ��;Hm�$C�)���� �U��8l�K1�43LM�v�C��ml���W����{:$�6���{���.�g�-.��x�o�*��MZ���M�f�N^�sZ���^���{0r��Z�J��d7�Yb��،s�pǓ�d����>Q�6�����ڛ=� #��������,�@)��~����D��}��<��߿~2Q��k�\c�^��Q��`��kj~k�=�%.eƁ�ek�Ė��������������.���m��;iȈ�c�T��zwe�����Y��+��[��Gl��Ng�1�-x�7GT��h���� ���xػ��ٽ�sf}�x�оKb�]һ;�[[�f�`����mV���۬�f�׫�I��3{0W�58;��[�(ҀVH���.(W��� �ln�λv��}W�б���o)6�-8�C��z�~[C���gcò�3��3�.:[#S>���y��g͞a�:B� ,����ؗP/���ft�V�.��i�[$o��*mz�_u��{{�����z9"0'gU��,��tK+�V+�65�dd�n�4F8�"�)&����1����@/��	X��D�MF.�˷�g{zi!՜�"'ƙ'��ڡ�ndha`�LŔ��TD�ܵ[�q�g'�e����:�g���x���w�An����m٬9�K��;��=�5��F�A� F��� �R.��:��`�鏪[�^t�OZxY,���y��2�3�N�1N��/K����U�c{��Ȭ�6Zc� &��k�'�k���SwK*���8�HI\"�T�]s=ܨdfϚE[���� ��c!w1]�#"�IYB��4T�i8:ݶw3�y�̼̉1��ُ����:b�(?G�Z4#KqY)O�����z"L=	s��Z"�o7����#����x�g"2:L$:�X�[>`���#Y
�����
�)]?v�_O�����U�ΌN:�xUY�.��"�A
6��L4:�q���-�Y\o:gM�n�d�������k�3��NW9Vy�/n�f�=l��g��Hb:.���~�)2��jS�b�����	�B�_6۽GN�D�dx'���>�Q�
��jUAgtQ��.��|��\�\yD�91�}Y۞�fx��0Ga��}�&�*�I2s���"���^n����'|v�:)��2�'���S�`�A���#��|/M"�b;^���[g&�x�i=��V���IyHe����T��w;���3�E&^����Ys2u,�]y���	�s��v�3��螻����8�<cƩ�Fɵ{��z@ᣎ6�E�}a����i�C�fN�I�vOƽ+$�0݈v�_2�fR���2_��6f7|��νâ��w��/V9��:j!��6����I	���VV#��Ԇ�3EɫI�Y`��]d�^��{j�p�;�{q�z2\��h�'aʂ�S���g)���Z297q�n3��0�@�]�VgYۨ6�c8]��]O>q����cʲUB�>�ָo��B�`WN��r�L�:>�W��]O�>�M�
�Q#T�,>�#�N�ķ������s����t�[�+�a'�5���.��)3�$�����y3sC:��:L0�2��������\U@n��f�R���)���8��ıWZkk�5Ӹ*SM8đ��0;�����{h(�U
��hh,j�2�ӻ%��]<{ȱ������"ɵ+�����v@���pht�s�޵=�K��޹�w�4�ק	�	�$�I~��㊫�κuP"6��I���_S��2*[
T ̲��t��%����\��J�{|�3�JW� j}݋W�u햲U�=�SI�l�lJ��_��VȪ�s���H��*$�y�D@�9��=��= �|3����B�=8���g�k�N����1S��6�dy�:Ed�|�NJ=$M>�y����{Ҍ���M<X�-����k�r�݀�*��c���o/���;��(��L��͂_{U�NS��P���`(�߯{'���k�]����b멈�74Wۻ�t�Ӵ-F@�x�7W�:��ܫ�fziU���Ry�ܷ�'��`^�q{N�ue�ˆ����l�6���pf�7�B����!%�xh���������nw�{	����U��6[����Xw�;s�cL��N��6�Uns�I�x�����׹7wRd]�i���:p��U3T-vhAi�کA,+{�Us���nWZ����B7Nɼ;gr��V*>��Zqj9t���s��X]�կ%�	�t�g;mW�r�9޲i�ט����1�ŝY�g��ݓTt�Y��wN�=^k��G��<�:�|Gq�-��ƍ�?LS��Q�P�G�{-]��[�:^�W6�����ۼ�<D4��"��ܝ��^�)I佬�<<��n_�*�z�)}�����ш8�/�"M{�Q�;J��lm؞�R·�<����Y�lO�K=1��6E{޺��K���϶N�����G�[]��q����-N�u��Wi��R黷��^Q��`��y��-�G�>˙I��e�iS��S����쾩�w�[�HV��W�wL�g�\�.e8�����X�t���Y�zʬ�ќ;����n���3z�F�4N9�;غso�[}!�{ҥ+!U��|hQi|��UV���+S	��T�J+�q�(6���)hǌ�h�=8r(q�I���.Zq*�Ҹ�YYR
����Z4M2W-S�g�'�RibϚ��EV�rR�Ȣ�iQJ�Adwj�X(����1����������g�c����AT�"�
����k"�;lխ�ADQiJ����*�JʋYkm6xxp�ȡ�/*�֖�f (?Z�L�O���"QF��Ex�ܲ,�e��b��p�g�>9q"����(��z��h�j�L��S<��m�-j��k��WL*8�LƔI33"�;#�V0��ӇwE�"��-JZF��T���h�
]f0+r�EE\�dɦ.��*jQ*4h��R�gm�l)��N�8.ݦak*}���uI[n�jc��kW,"�j���S���[) �4�
X#!��M<8rx��]"Ҕ�ۈ��EĚa���T&:CY7�����Y]��Y�D@�`x�'mq5l�4`�ZԊST���CC.�b2(�P��0m*.\�2�uj�P�TQ
��ϗ�a�n�*V�ww&�j`͹p���wbW�x�����^^o�dn��سr~��_{d�y+�S�z���x> f���p��'z���l����83����=����z���SF#h�.��f��N��׊�Z=.�{c�Q��<'�g0��B��w��}��ػ��h�}E��*��$�c�1��F�s=�me=���l6w��킎x���E�'�6�U����O�%��Tk�������\ݽ,=�����6t�(H�MOVfFa��\zyQrm�튧�|嵕sK��˫zrd����w&�~hn\o�/���@�X*��.|���/RЏu�Q�:z�"�h��*��S�����t�X��}ʉ7�X�y��4�`�}���h�L��rv�Z���[8@����$l�kե��e>ffi�\^)\��h�P��S�܁�t?�Y_��vcʣ����&�����;@���lDx�R;��J��U�(�&��2�O��=�1v��2�\UL�=�)|�G{^w����i�4w����)d����a���+}W۷�/Hu��'�v�������Q�6n�,�n�/\W��6�.���'/_km&�`��G���� ��k�A:nU��w�vꟻ���:�B��/�%u|4t�-���u���_v9-�m�S,�
%�K;D�x�|5�4���=^2k���1$z5n�AӉͭ�7��Џ�<����������h;�F�9?�|�`���%�>���}�I6?�MxJ�9q��1\K?U���̪���>'t��,;p���3�	XO�ޘ�DK��*�V�&�	�U��DO>R�V������Ut2�Y4�|��{X�[���.gMO�gK����_+a��t-��xyNׇ�!�KP���n�t������ߞ�[^�;�!���ͯzo�309[��(wGO�E�i׾U	�/S\��'�,1��
�8���1V�����D���ǐ�W�^�Ǒ���.:��7��FC��p�t����n�'��鷘���<�)�o	�v�Z*��[+)O�)́����x58�	����[�6��n�m��)�)���,mN-\��=�.K�Z�����`�[T�hUT���q�E�i��F��-7�6���"ܸ��$��YWuc�e�Ǧ
�M	V�аTӑ�^�D��;Y��zs=�^
�x>�i�/��x�a��sO,�uv�����������pO�H�2���g��j��I�q�qc\1�5v҆�+k��{ƱZ�I*�g	��AeP�Ĩ�"��#���F�μ�iV�瘺�v�g�.��oj���CjQ2�$eT#2v횙��C�@���j�M��;L�Pb:C��(���0P���%A�<�U$Wk.�������v_z[f��x�>φ�
�:A�*M�F�$*զ��ѕW��YNg���L������]^'�cǶ���P��u�bxt{���DT�,"��4tmL�Wa;�.��յ44�_�lkX�p�u��0�8k��^���}-o�}�s�y�
W�ɲi����$��������mq~���m3���{���y/Є
�g���\����⸆���(�*�5Y#i�4�J����V�՘�|@����4�q��6�e�T:8�մ�:���v������b��0�.��ṅ��8�ۈW������s��zv��I���e����0�U�xK�LMk^O-�И�����[k{�lܳ:��5�o�7{����&�O�T���fn���;��	��Z��9�� ��}��@��/Y��I���a��{|�!P��t��-�*�v%����d,h�L�f{z���֫6c$�dutØC�摁`��|�������+gZj*j��l��n���:��5�N�=4���1/��)R�Iw��Ї����C���Wt]�D�Q��ڡ�n�E#lD��[>e�l�"ko4�d�xP5u@fH�܅�{�R+�5dJ�V髋N2�Y�v�SW��|�Bx^���n;�r/RW\G*Uq�hl<�;^[̹��u)am�fա��E=Zbm�L�6��Z:��WD��l'���Wme�f,�ƺ��W�x��t��L���!co�m�nȝ1l�w3b�z��ՙh6BT�R�/^|�#r�vfH���B���s�r�1c��1�ٛ���ҥ�,��!'I�s��_��J\Hn���Os��@�Pg��;e\�xW{4���n�j���	��{�ٯ,�\��MY�$f{9��1uҧ&��qb��]������=apwU�]{��k~�1����{�9ҍ�~����
�u��+�h$�wZ���;-fn�<if3�hV�y��f��^^�3{ʁ�;���Q֥W���ZaoԤ-��09�COs��1zx���؍��$��-�>����s���{�*Y�(�T�t��Om�f&;�2!n#E�y���n�ݽQ	H2Iι�ܺU���!`�B���m�nm�5�J�*����qf�5�$dA�]�m(ۑr%�.T?P�m�&w*O]gw�m	};�)	\v�St��b7��(p��]���/:k6�n5J�7D�m+]��WӇ��oX�s'�080�4l�Q��g���<����g��c�x��V�|Ux�$�x	���i�s�Bf]�-�3-n5md�g��t�
87�[�o{�Ca�K��O?����)5�]���j����ʅ���c���q�I����,���1�323	M,�\F�b������`�����L�p�c�Qo���AH95�1ӗP1"��g�IM�����~/�f0\�v�֜�]W���|�`s�F��y
�5�&rԃW��<a?��W��;�ϳ_ɜ?v
9��b⢧�9E#�۵�ɋ���G��T�|t>�`���MBQ���\pK�X��EH(Xnv�b �����{��r�C��"�Ձ�՟r����R.MC!9���t�X�s1~��9N��s�n��3��ݍ�Z2����Tәl�k"�C��ј����J�]�$@�m$$voAu�ڊ�$��n�i�	����4ݫ(�m�<���½��@��>@w2��gĒ�����t�l���'/7z�9��pjC�������:��0�J�R*�n�6,�Ce�@��p�}��I��u��'�tϙ�=�S�p��>�o��t8�=�kcE����^2m�泆�ȕ�A(��(�{����p� ~"
����]Ct�Gp��]�ԅ���j�t�����i��^3��7�}�f����}m�}0��P��w;�Ջ��=�K�YD�P
�3s�}�p���:�)�%�Z;�>�_a8�C�cʠvm��A�����N���zD{�6��>��f�ٟ���{`��9q@��y%D��b��޿H���{5` �zy=���B�˥�rxԹOG߅!�:���ׇ�֪X��f���Ɲr��{4�;Zo/o�����$�y��;j�Y�Y���o"�^M4y@��t�|���yF�4d�a����i%��Iؗg��
�r<�fDV�e�q�@�- �x��4E���E,m�����M�t<�8n���v�U��Ћ���*嗝�2#�
좷jc���Zkt�"�Z=�)O�)���{!}�e��Cq�lF:��:v�%��K�f��ˑ��"�,㑇a}H��^P��B�j�?=M6�Uf�w](��)��M%^(�Nm)��(e����C;-[5�l`���N�R@�TDv�ظ��Y^&�T-A�Դ�d݊�-��jq\%3�=;�w���[BB'V��Ð�%�O�J`2����g�2%�c��Un�;���Z�궸˪����b�mH��H�aX�Oy;4Zo���my�;C��G�UO��.t�Dp!�)�.�1�kS��ެ{�s�6�fMe}&�l�'Wu��>lǁ�� ��r�p��0��zy�|�/ם�Y��Rk�DU�E�+n1{K��-S��b_���T1�/���y+P����wU	;�V�EH�cֹ�4sdHkt���:�_&��G:K��w�����E��gz���j>\��4u�:k�f�*��R����Z�C;B��6n���˫}�L�E1�:ًeH�n�0��Q0�X�޴��#kI���X�tuTύ��rJ8%�+��1��Ǳ�/���Ub�`G5��1���G]P�J���J�V�Z6�em*4��;����ߟ�p��Uh4d8+����o@��յǺ���Np�r��(۬S|r���
B��|ڃ�B�P3#�f3�.�S�/3�eC�a��.�����ّ����:9�8R��pT�eJ��ɫ&���y�����p��Y��BB3�;���g��d2���u��m�����f&]�[K �����.z�;uW�.���Ϙꢗ�>���aۮ�*]V�ca�����'&j꽙qh���*ПDVJ���6�{�K�h����p�p����<yPe�=T�zf�P����,���*TuD��
�6��>����ύ�I���u�����9�eGf��^>�wp��~K�Ő���-�M��Y(8L�ۈ�^k7|��D�E��������E��D>�MG��Խ�0��կ"iP�����n��F���bض�#k1�� k7�����t�<`5�2ۨ��3��+�,Af�գB1p��F4�k�}����ɥ���'���^OM<zi�=�A����&#E�
~���ܶ��Q�R���*󥀫s&����:뽔!g����0�en�(�3-@���~'�"W<�K���[-T�2�^�\�P��.�i=`pq!rcB��8a~�+4��3�ԥo>�����+^�/si'���V���A"��:��vhJ�qtMJ���g�����n6{��-��� `[�[��WA�t�j�(�M���,ꨢ��L�����w1t�Z3� t��a(f�v�<v+�()�C��ȑ7uP˻4�^r��H��'��ݟ���y�ږ��r7�8Ղh��d��bI�������6���ֻQ�t���g��G�l1�������޷���&ڡ��9�×Y1�#��{w=�4(��d^bY�3{ˁ��ޯK���Tz�°P'�&N�H�mb�<���IQ�Q�ye��H���5ɒe;��d���$���"t�M,���xo�1*o1b=�D}�;���4�YM�P��p�	��~ ]���9[���o�(mp2��2dH&#�WN�s�m���j7r�+g��%v[P�Gx�Ԭ`3[�s�t{2�<�w�O-@!@��\.�q��%�]�ɵ����iחٴϡA[Җ�&��ff/@V�K��b����fWH�U��������N�}v�C�	5�1ӗIDX������S��uY�V��*�7HSJ�*(�f���9��)Նj�����5e)v3�jګ37T�{������9ܖ��*��b�%͋��a_�gY�*��h��Y�	�r� ߱	�]-�?�B4O%P�� m�ևP/ǰGKJ���5M��3x�V�
�4d�=lE���{�%la*d�$��Ju�m[�L,xn�����u��U>�P��О��Q}��_*E1��yĈ2��jz\s1�O��َ���_K&�RAۂ��-�ΓG�ߠ� 
�<`UGz��#k'�M��Ş���>^u�@�f�g���T�.�����A�jz����H���u��ݡ}I�Fa6YU���1}��F��h �nh{��hP,��[�<���,�'����ӻyH���d���}ꃝw�u&���?����?�szg��kR��}ɭ9��+ļ~f�aMސs�V����y{Ūo���xFwQy�i���A8�|,��F�M�H<v�&�^f!���G���56��ri�3�̯+���h����lj�q՚Y��I3\\(�n@�^�~��f-]�@(�.Ժ�:�7U�ig���õ�y�6�b�g/z��v��ɉB΍��U�2��&O_l�6<�������:�+����Yyb�1�������r����Fn͕b`��z��~��}�c�����6�$�aΕI4sr��Nѫ��2G����'�:^���Q���{�-�6bq���y�N��������t�Q�
b�WWEZ���\�+�I�yM�E�W\]e	gu�Y}�1As8n�3�����o�\�t�zGIt�W��Ơ��Z�
�ΰX�V^=-����}n�F-��Us)EE؏^ƴ�">t�yd��/:�(rM=}V����5hm�}��%)�@ʪ1�F��Xrڣi��pjN=a|�_Q���eT��l_hx%\�ƒ�L�K�}�k1W�VآN��z���٭��4�H���d��!�zl��fVۨm�K�U�H�+SՊ�0Rm�3&�:AVL����c�
�R��y�$�[sFq���k�f�����Quje���{#wv�:�[o���F��-�tﷱ{'k ��;�g�f�)x��֟:r%XL����0�f�!EJ;��,�Xdr4�S_Q����wU�w��yջ�vw ����[)�;�s�՞�هFl�PRb璋��Q� }�<i�ԼI�Nh�-�h=��Pxf�\6�ܫ:��7
�GX�����(ܜ��x7�q�������p�徾K���s�OS�:Ygx�vf��S��޽��[�b���ޮ���yI8zf1�)�g�C��s[6�K��k^G����-�[Z��Ki�nR�݄��tА.֋gfx�+p�^����!���1��ywf�!g���>v���;���֊��v�I:\��G�to4�e�z3�d��o���3�����W�p���U;�^����8-u6�UgC����o<u���f�	������^��
qs{��l��Ó��Σ}$}Q/�b�Z�A�^�qv��L���\0+�a�4Ĕt�b�r�x�$�6>��E=��v
��h@/,��̧9��Qo.U��Un��77���uU0)��*��E����t�[�S�Z�rG{mE7��P?^WCEn��a �-F�BT)���&�	D�NkO]0����b�H�@c�cn�9�q����WK�1ĉ����E���X��!U����]9�j��eWZ,5KI�iK5LeAE��F?��Ҽk�GT�PRj�F�)�cR�����E1�A-�Hi���O�f'�f@|p��6pDc�eF�.� ���y�"�%dUUb��*�ckE[[UU�hWc�btçN����">P��^0������Q���w�%�5h�",DQ��qkJ1T}i4�F�=8p�q�
RT��TϡL][�+U"n��m!�\�p�e�U�����ON�DD}j'���6�E*4���AQH���Xb��Q5�T�.�RwGN<<<��p�	�Ld�,b",4¢Ԭ��1Ķ�m�r���U*�)ᇧ��q�C���Z2�X&�A�e*�o3lP_"�e@ynR��iըσ16l��Â"Ȱyv˅�YEcm�E�RґAE��U����\�X-j*�N���r�0��Skmh�Z�����+j"�E+Ec��)v�I�����q?H��ν���#��}�ι�g*�3J�LJ�n�`Ih�l�j�u��t��Tl�ٽ0�����+��7�S31!VV���gi��A���]KQy����u�Ľ,�E�	��9�{�D���з��X]C��N�t���N	���n��،���[9b��\������ ��>��΅�y���c�F�,fv!��=�9ᱴ�w�Q5��ު��O��ddd��{�]7zt��� :�2�e�\,��ψgr"w�g�1f~��v��ȩW۽�H5����pLA-�r��-����:�t�dx\USV�Ǎ��|�F�+M̤3��A����p��²��.�c���4�K>MhPeo'�\`����Jv)�r�wB���,��$��9�ڮ�̸3��h���j�M���R���UҟlS���������F�s���u��w�=�ؽ3*z�]����AT�F�si\������qwl�ҋ�����K�=�ϣ/��\d�A!e�"�'mQ���!���:��\�l�_#�~;}���Q�l#LUVeN@�3����}��5b��Լ��c������w����$Z���
��ߣ��|�]�O/(&�1��{����}!w���>�2�<'����,�V�{f�9Xg���"�����fdq���1���j(B�\/V����m@� �J�E���W6)�#n��"���=?!h^�O�%��b��<@�ƞB*-�w�H����ǎ�����'1Q����t�@����A�uѮ8�-���kgL�\�N�<Hm�>'WQ8d6c��A�!kv���ĩ<�gXh��Sن��5UE��ڐ��Ƒ �.��l��*Gst0���3z�$OLN�UV����|�1LG-���d��5�(��r�|�.Y^
�k� VV��:`��@�9�%dF����W]z.�Д���4���HBrf���m�u�*����L�0��<F��>�J$C���+|:4�mX�թ���Ls�]��=s���ĄX�T6�Lo�|��H��A�N�ۨb��l��i��'��"ξ�$�c��q�xN�F�Y��}]c+�����ˠC�}�;V���r)�Pb���kg�9�qSN�*�l5���f�r��ǑI���h-�A+w���1���	@�FuBb"��gr~+��g;�7Kpl���\�p��y�:�2�K�~�W�R���nQ��>ɭG�#�>tb�����w%�`�'����q�K&����g��J޹Μ���#m#]�0�4�ܠ�kksc2�@���"s�-�@t[�.w�5pA��U񳠋F����f��n]�#�_d�BA\;T3ꇌ�8'�U���u
��D�\��K?�c�K����͞�ȩRP2���9ݻ��V���V�f�m�����i=Q�u�� ��0���V����p���P��ּ5Ԓ�Y�{bp��f�I�g�U�w���j3�
�$72�Q��h�x��{��]t4�2ܒ �\�R䞻��>��NdzE��h��*7��&�.v��`�
�j7`�|�%|�R\h6�Hj�!�����&�Uc�Ui���#G���"��R�v��*���a��ҷ�t��͓�A�_g���������!�����u���J��D��2ZXne-�7r�9������Ц_��-�=�f�v�Y��{�*ŕk_�#�6ͫ�B����༪&5C��wEW�x~G|3�aj��0{)k��%�G*�����W�Iw�	�+W,���
�~��l}�+�Ǧ�L�|�a3F��D_N������y{ޮ����5���W���[����a�l���@D#�����2sq�f�l9��l�;�	fo(�+vM���������P�jދ�p��8Uj��|�w�/�\��x�J3�_�� y�L,UPb}^R����l��Sь���AqY5�WjF�t������h�p���ô�����C=n`�o*f-�2�4L�A��0�w���Y�+4GyN6Ĕ/��l}m�*����}xT^m����h��r0F�iqʌ�i���;z�98\�Ӊ��B�"���W��z���3S;�&�Rܣ�� ����n|Eeh���� ^ҟ����;�\�b�	��8�.�[T'�^�mrzNi���]hg dR�
�WcO�iH�����gB��!�(�Ȋx�l�\�_Y�R��T#";PW]�*�lR�GUX���m#y�/����2o�y<
��<��j�����8����V���nv�4��T��u��)fR��6��S�0���[���y���`Mك�OkZ/��̅�>9��@y��_��]ٱ�{�!���|-����E���j�F>�or=����R�zĜWr��D�JDp���]4M(����V��/���8٠��/�e�א��]M�#Ύ�yXW)*�붰݃fM�Db��ݽ�w��%�q�HɄ�u��Ǻ\IkA������Nl?c��|i��d�-
T'pk�r�Ԑc��Y{ݞK -��N�o�0�+)V�N@�{M��n�u���ly��8n'ѫgs��h��}�+�X_�6���=݂醱��#�]�+���1�a����k`�mt��+5-�5��i�N�իd�`���wM��i��v�@ޱ!�.��.]�1o��~~�.��-����<��
�Mͪ��Z��b�L�6��-��e^i�i�|�4��F�nU�`�����N�z�;�b2�ԗd苫'�vcC��h&CH����ZA	C��n=�['q��$+�i�D�u��Q�F���kU�0�-��A�pC�P0�J_�����fpj��Z�x�%٪����z�U�'���L㻻y�C��#v��+��u�}��+���뗾�4͝%��4�p-��o�����G���Rw���g��og��w����GB�>���iЛd�n��T�+�e�v\���/n�ot|q�~+������/�����F�	(�}<���FFE?NC:�W0T��䚹�SY�D�i^�\5�7Jԩ�E])�@�g���5���'��k�"��oXd��	��Cr��IBEr�R+���i\��z�.�c]�sWa�jR���`�5>�B�P]J�z�ܶ�Q��:v�6��Wƽ;4�H5�7��1�9oK���^�<M%}L��ꨇs����=o�*��:d۹�nf��Ni�š�G�~�^��YO���7җ{}��\ʲ��J�J�?h���}���H7�/q$�0��7^TJ���jYjY��"�UV+�m� �]GA�@6��n�v���f--W���� T���_���xh��4�[-�Z�=����Jk�j��{������ֆ���h�B#�vzz�Ϻ�Ċ�R]�c�dN���AM�Uz�Z��Z6.�nfj�-��bWjtjӜ1���,�30ޙE�rm������ww̚gZ|�#�w����mM�\h�����5�B�i]J�&o.{����k��e"���C7x�u��=|.�;r��XY<{{q���W~D+�й��������(�`����>�5�::�rSKt��"� i�7w2�fB@NџMa��6lpހ�# Fȹ�A�]{u`���d�Uy�]˭����+���n�c��&Ƃx?�?�A�X3�(�!"����թ����i����oP/�H��%��2:��3�!��9�Bօ��2Z�����y��Ǝ��j�#г�n��zo��|t��Tm���fꪺ���V��8���,�S�%C3�/�=�����������tn�cR�0�1������l�F=�U�2�=��W22�-:�|A�Hp�3�*)����5u�Z��6U9�l0	S�I��E�����{3��ܚ�}b&�w+.8��=��i�TK顚|����2��E�E�+�5��>+ʛ�Lެ�-X��2�c��^OM<M3�=�|�z0� 3��Is�_:@ݝ�U������/	I�{��e�=�wc�����^=��5������P��T��߈�����q��<����T:��J>B��<�+�ev����%A*e�\ʖ;�%ԍc���D����<0��m�;p��g\Ժ��@{���u���샙�RF�J�*C�i��|ܷS�7t��vf��D�N��BzO3��m�=�ѻ	i	%-%���Wc�x���9��c��&�wNTC;��5�yHV!�B'�7l���P���4��m�cWa-%��2{u������Pܒ�p���Y/�t���zL�ؕ]�#:��t;�V�:齙7����|��7 0��~Zk� ���]]mS0�W٠�o\wMv�B��*V���a��A��\p=�U
�4���H�5��̮׫������[\{�\�>=C���G7��7U�Q�-��_��8�O��`��;^�	t��oO��0oa���1��h��P����&٩n��C��e�8*���:L�� �b��իZc��z�'��fo5��T���~��f�|Gto�m��{ؘ:�*��!�;?kO3�}j|�:����<�IWU��d�>��xw���G�V�Hq�;(�*��Ը���I��P�����8QRpJ�%�*�z��t/q�Ν�J��c��p�k�w{\����_F�������Y��Jfvb%��$�*D��H�9��?_v߯ޭ���$��`�gsZ��E�9�a�)�N�ԗ{w����[蛧]#6���Oɼ@��<h�ܛ}{JGE<�xLz�r}a]�>�[K">0�'%^r�s~k`���)^�(-Z�m��E�9��t)\O���(:f衐�{0��0�G�Lv��=���hA�-��SNa���*1,PW.��g�cb���t�x�-B�i��y�&��!+����!�������olk��v��@�ⅺDu�6��t��a�	Hc��jL_���;f߳'�8�q�oO*sf|�N���Q�"SS�u��u��S�~��>�ݕ|^':1�	��̛�����7J���;��1ga7��}�F��[ۛz9�7E�ko=��x��z�P��������a]�bCu�d�����������&XAw����b��ܺ8Y����=�F�O�3�u��5l�]�M�o�⧛�$6!ׇ>t�f��3UsC���:��G.
�5�u�a|z�0��HTr�!�%a	�H*�������r���u��\&p�4�1A2{��E,�օ�۱{�b����sf+.�{/���m��/nͨ�
�g��۳�<fg9�x���0*��1ϰ��{u-@�`Tҷ�L�U���xx��e�q��y��ʯh1�c�1���_z�{�l�ώW�����[�Q�w�۸��3�E^�AHn�w3�����fDq�[7�)7T�@��9�eO\f�6����toh�����؎�q��z ZEM�V˹}�{w���5���b�V�O"$�xO��:&�b��:�;�/��^'h����q�y��&�(��YU<��I��	�@���.l�	kAxu�R����2�Fؚj��D�T��z�\���$Q�#7E�I�D��1RK�;�e7Z'7.�Wc,�.���j!Y(<����V�%l�ۺ�{޳��û2\�SA�P��j�>{[!�B7�+�l��d���E���F���'���[X����:+m�y�A-1bok�G"�b��y|H�ⳉ�c4�Y2�3�%,�U�iM�w�Z+��[��a�>?{ϏD|����Dܣ���#F�J�l:���PeА�ݠ�v�Ƣ�G;6�T�;c汛"�f�s��;總<�3ހx��9r�x4������l�`�U�a�[��N~�ǌ��� �m�1$���7�
�6�o�^���ծ!W�d[�x7�~�E��.��w�^H�d����^��&)�o�~������j
�`�������,�ۍd�����ѽ�t���9����|B{%L{��_���\�u�-����k�Ҟ�=�} ���-���p�2=��C��G{Qƭl;V&tUw����>�|�:Q���2J̖Z"Rz�aΎ��ѽ��/*����׸�K<��)�K*l7�`��%�9a�.�tų�\b�����z�~����67�f��k���y��T�sUA7-SJ�i4~��8V�9�.�Wq��P����Y�ocs��H˲�M`�rlb�-�Öa��-�*Ml�8��h^G������v�\�OlL��D��f�&��m
�Tv���ɖ�Xx���e�/|��\5�
����6�=�a]"�GW#��vm�ަ�������zG����=A�{��;O�+�����w�/ g40J�t�|/������|����$nTꍡݪ�
�w>��-!Z)5]��m-������3��ݺ��C�^*x�Av��6=˱>vU3DLG;jj��O&r3GD��e���TR�V7j�l����KrgC���s4��T���dL59n���M���p�9�g��o���9�5�
T���*Em��e����4)ԛ�5ܺ�r��mm'|ﱾ��B��Uc��1t`}x�h�
�Ƀ�����)
�L4�8�6$��y�˦���e�l�cM��Y|_<;�l�z�%�6�YWK�����1�R�˫���ܡ�����_��K^���U�0l�p|�{��o��rA{dg��aX&�>�Y�nyF�5��J��	�̨��u�C����y��{��^G�GXK4Z�'��B�0����3�v���0^}�֎��� �W	�cթM��{��=�ʡ��~��=_�v9��lr�Ǿŀ����<�v�oYBl��x��Y�w���,�+�{h�}��bI�9���M�Z�hV�[�_x :n�h����Lw��ib�'��:7�����0B�tEM�����;�j^�|�5$􂷕f�Z�
�b�=T���y�yJ�E���Bh͝��Ey�&�OO:�祏nxbW{o�4=�y7�z^�����������#eK{�\pȗ�:0��d������՞�4��9���u �Q�݁e*�l�Pt�a�t�/{O;(I�=M3�I���;GS�%�v7M�]�����a�I��Nn�c/x��U�W*,��w+nqcar�9�����d��GL�0�v'�U;I�RF�-(�5��X�nJm[�"~$�����A�lDKh�X�&2��̵E�U��)��xx~9���(�X�b� V*��"�#'�E`�YX(�A���N�8p�b��
��Q�}���f"�D���m�V(����===8p��imyk"���D�Y�"�+iQQ֨��\~�d2PEA===6r(�X�b��X�-Q-�U+:eUDT`�Ub�5Jٖ����᳂�(UU��".�>��m�"�GT��q�e�F,b	N�:p������G3�KJ�m�Av¾�V{nڌX��c+*�5kE&�qON8q��.5E�WƂ�Z�nS
��&7��5r�G-XŶ�����k:t��ÑEyJ(�[�M&�J��֢���������S2�S�E؋M%XUt�*�iF�e�J�R�q(��l��9�Z�I��j��ŋ��r�?!� �e~mU{��؟�v5v?x]��ݵS!Ŧ� i�Nw��6��7���|EB���*�M�+0�4��B,�(����</{����Y�Q�&�M�|��oƕ$��~�t�F�!�=Ӥ9��mž'���W7ٴ^̲��?t�s�4�&I����Gy�_�g�n��}�a��V�`W��3�l��*W\����q�;i�,�8UUv�n�z��nG�F�gg��h�[\�%4�p�=AƖV�.��}7���	?E�����]��#WD�vt���%N(o0�G0���;���j���Ud�i��<�j�dF�6Y�C+���sw;�sF�^.{��wR��vP͐lo�������8a��e�<���`A���%ɶ��0ç�l�Pc�g9��
w�Y�"�,��f�-]�7Ge�I���Ğc㢌��S�=���E�2���z�[
!L�4I9�Ό��;���
B%�z��a�򔚻�mk��<�A�_���Q��_b��<��á���UUR�U;{j$��8��K��uhT�i�}W�C�m^���j���/v���n+U;��4/&ĎY�*�{T����{��S��m�pp�*��,Z�,[��]U�㈏� ���gzx������aD��F��g.��#�����k�����ڥ����"��z�ev�u��g�^�P�z"�h��WdM[�f��m�za�k��I�g"��E��7����� �,Af�U��SN���fgu\����,�iG
=$�,���'JNp���y��>'� ~��s�3L4i����ggͩ0F��T*]M��r�^C[⶛ׅ=��c��h�p����8N� �T�����%��������+�Vs����,��n����:����1�#�J8�A�J��� �M��k^yuuk���#̿��g�Ͻ2|�4�VX~�,.�v4quٗ��:���o����=������o�zL�ϝi�p�ئ�a�f6�� ��Y�[��u�T��Oͽ��3+��E��%n���Dh��`����|�1Jn�e�j��뼻%�U�g$q�v�T2��3��Նeyź=����=��&��ˢ�6j�ܛ�d�e�A��@�͇���nyC�����j^5��p�u�@��8͌�1\u��1�3����;{�f�e�[|��f�e�2I�jAg���'{�ݝ控v�5�Vg�ѣC���Fh{�^R�=8�'Z}��1��()\{��a�. ��WK�b\�g3
�����ɢ�m�W4�9�6�}�=7I��p-Õ<d_<��mq���d��$��v/D�;]�'��I'FM�+��[�;Q�,�xD[dV#[�c�2٨�g�w�ڡ�uwC����I�h���a�́}B�=%>���}d�1ooj{U^�އ5���{�m�.yz�g��$隅#��yWb���`ظ>��763�Y~���T��l��%���[��l���׳z��ěPA�f�lH؏V��e��+�Z2����x��hS�7?5�k�/�w��8|�t�e#�r�ՄO�HnAtI�k]؍$�mükU����S]R�f�®IPl3k���'v/�{�x��ї�*'i�j�p����І�3��goL�Kd�����{з�
���[�t��յYyH(_PgnS�+<#��o85��Jk�%�ܻ�6s�=����]ְ��n�F�=���y�n���x������֪�G���3�~�.\k�ϫ"n�~$�*~��N��u����"�����T�t��ٺɦ+v�h�����H#H�n�>Y��C��l6�p�Z��Uݴ���]�f�+K*�.�v�'�mlN�V�4)q~�s�ᵷ����_8�O��o���`l>~�NA]��j�F&�'wM��L"�U���X쥽���b(wG�j��uH�'Uz:j|66��B[��5
Z��5�;�n%����|)�N���C&��^ �C�F� e�}J��>�_����x*	����ʹ�ͅ�:m �ԅ�}�0����tl^GT.��kr'B��a�����_O��mr;�"CµU�o�yS���en"[sQ��7/��H$��n�&��>�{6� A�2�X�{ӣ�,�4����͓�����j]�Zȵ\������(p����xu<����o9��e&'X$Y{�N����@�'��Ut����ū�G�%�ض��粭������ZӚ�m��i�$5��F�����^�䧧@�Qr,�?>���	���vR�o�o�)�kOt��#�9F�}�y�t���@�o�\A���bv��p5$&��4��"��pv��.2��^T�۪�뺓����+�`���TN�"�v�ʂ���h�ƪƼ�ʮ���qEgZ�ך+�V�na�� ����B�N���ݥ�f����g��9׶4Z[���2�e9����N�Uy��|��Ά�2�E���Y;[9y��]��ٙ��fCMx7A$�\���u�������Bk�5\V����=����J}��=�%+�:�6	8���[1�/�z/�8��j�'U�i�xxHPF�5>C��/m<�T�\������|�3�1t�ws��_�F$-2�p�BBa��w;~�����T���xU�;
0�ekVr%��ù�n��Q��s��-���t\f#�gE�]��{�P|'n܅�M�S�u�z�~�e�~�X&�#|�f�(q�
��p�fV���>\������������W+;ו՘���ޠM,����mL����# �_��|=>l3�~�}�c6���-9����R�&bG&Iݛ�P�6;��g\�3��k�*�����(B��Ǡ�O3���S�j�VN�}��IRv޿t���E�+���OI��z"�|�S���?�.�u!���>���}����O<��6�Ob\[ah$H;^�zw:��ݯ�O��|*K���U�H��Y�*2u�&|3p��;����Ė�	����bL��m&۷Mm�L3�Q�����|�ѱ�"E�d��a"J"�������f�wy��7��֍�a
7������gm�$9���e�fε]��y��i��78ޱ�EĝT�`���_0T�Iz8�y�B���>sG�價��w�T�ga�B
�%L��(�O�TTK�YА��ܳ��^nPy���F���A��1p�`%��h�*�ד�G�5���(����7w��s�1�>��m�<8�<�T���A�n���c6�:_) Ptj���~�V�=�l�������G��v�G[�J���l����_��):�LHzMk�ݬ�E�w���W��w+�gL�]�Ww6��[��Hu��ݵ|��dڮ�~�����u_yr�$�4q���{rt�H���N.���-�����H�|��uO{������� ����SA�~�OE�=����&$d�ܹ��N��C��nۂ�=؂�9*�z|t�b�D��_�-�Vѣ�v�l�#>[ϳ���c�z� V�sк:������4�ʛ���sÕ�%DҮЬ$L���T6�ll��������Ѻb�+1VԳ������h\�I��ǳ=&�P�ܢ�@�1�]L f0#r�bKe�k�[�}���X��j��U�J�`�ܷ�wR��vF��n��W�����tOUT]�=�$&r ^�q�� a!6Wi�K�q�}��{o�p'��=9��_�hs/;Ɩb���8q�>x�5�
�ݮ�Z&�2b1,z,�&%��^�Rμ�4Et@�Ӫ�Ϻ�.4YgT^i�icp��B��U��y���{]ӤO��8�����c-� a6��Ȇ��7!�k�Sp�ԅnFbA��R����0i"���1����T��\�|FU}�_�z�d��(F�[�/Y�OT5������5��:*gh���ޡ^�0݁pOmǾS�f����p�P�N���kpҺ��0Mj�
TU[��V �JXai�z�J�3^󎠸���O���i��w�v+U],��?|>�oF�;݄�i^|�lL�O��w%�0�f�)+��%`��8zͼ�lSl��lN,�Z�lk��C�S�X�Gj	�e�e:5;F�Z�m��%�GM��M�on6i4���U�tr}r��XD�.��Ѝm�=�mP�˚����j�#p�y��v���gCRFg�(lD�&��w���xI鶺�w�z�j��&��2$�S���t�|���p��R���̫��mD�]n#��U�%o*EXҤ,ݞ��b��\ �ET�z���d�s|L��x
��*�Ǎ���"H\��~�ކ�z��5c��8�wPX�̓8\3>���WjڢQ����wd��QڠKOfR}�����\���#�l�*N�S*v6��ܗP*������g�R�^���{o�eS:8�y��n�q�01��nF�R�����{=P&��[>º.�fq���Բ��'P}��<����:����4Z�����Ξ�>���:Q�V��g���#�^�c�\fiiƳJ��ꩽ����]��m�ĳv��=}����'c-�qL��e�kI���|=]��Y�D��f��f��+���y�c��5��c(*�/�V;"�ONN�Ug�p>����c8�d�F����E~�s��C�G��#5f.�y�聽Ք폹a<��#ăOU����3�۪�W�V��E+�rZ��p��%B*�����<��,dW��'ܱ���3���6l�������S��u,�� �U-���m��jKC_ {�+����`Ք"��D\o$�_p}�Ô�,₸��C2�'0����c9���{����:���M.8�C����Q��$[[������B6�ի/P[Έh�ǎ���j�ʽĊOA#*�;U`j��^[�4��Z���#B��\�fmtʤ.؈X�|�Q��*�y$����]Xӛ/�N��;��< 6�����i�͈{)�����RC�څ*H�P'
 jB�)klHkל�2�c<�@�Hq�=�yW�Ö/�둙�i�WZ[G:��:���3��k=g��쇦�38X�Є��Ǜ���m��iN�v�k�^jcbO��:�+�p�u� ��35C^Ҋ�I��x8�$�q���a��Ҧ+�M{����ۀ���n�[����/{u���v�^�xd��Ɨ+�]�
Ķ�ml��nh�6;i������[�ǜ�0�� y2o�X�Y;���},P��;��x���!�Ǚ�+���K�̀��#-��.�:�1�l����]]K0��xő��]wI��4wJa\������#6�`Qi�����������Y56@�*�ռ,�Q���C$m��6��tVM�Gk4L�dV���Gq�*�-�[����ʿ����A��f��)N/��:ͺi����[BKtn��3��ti��c�e.�Lqm&:i+��u�Rh<��+�����+EZ5��3/�{�(^NWN���Xz�D���׵�ndh`�l=�5s#.��i��EFwb��˹��������C�ɑ��8�L��������O���m�ƤR���Q��7���� H�k��-���M�E ��IXJ�J&P� @�@ �	
 �HQ�(@ @  a �	�A    �� d   @ @   �! � 5`� @ @@ `@�$�     �H$ �  @ � 0  �$� �   @ H H  @ B @ � Y  �0 �A$   �0� �  @�H�H  @3 � H  	  �0 � (	 @ ��!"�@�@
@$� ��! �;CQq��%)u�T�0*�_=��?�����������s����|.��w�i��/y�����ǧ��>��J��{�����R)W{z�J�����qxK��������v_mH�_����K�K��5|/�8,��^�כ]�J��C!�YV � a$` I B0 �  �#  �  " 0H	 �`���( ��E��U3"�y�@bPY� FH (@`B �d@ 1�DB�d�� � "@	 @`�	 H0�2 �2 �$��	  �@ A�FH�YS�eVJ�eYR�x{lfǟ����rQ�
f��K<'r���f\�=W�}O<|��U�6�����yW���]�h��zT�U�w^���]�Ʋ�R�UH�^����E�����
QJ�X��~�k��>-���_��ˑ��8�˥�ฮ1E*������R)Ws��e��~��W��Þ�]�.�w�nmR)W��}u"�{�N��p����8<Vms2��~�ǚ���_;z�����2�W��{n���z.����ww�UH�]��k��ߕH�[g��]=\���]�1AY&SYb��c ��Y�pP��3'� b@��/|^��`�QD�URCYU) $�$	TIJ��J��B���$D�IM��T�@�R� �$D��J�ͫl��4kKmm1e�5k&ڬI�XU��,c%�h���Q�ڴ�m�kmY�+`�ZڋF�)U�Fci�����f��jͶ5�2�6`m����s���l�6�M���Z�f�ڛi���U�ZeUUX�Dm�Uڬmd�[l)�Y`�C#[cQi�*i�-3f�ԭ���%�ډ-��ڃ��  ������o�n���y�YN��^�uuK��s��]�U�w��a��z۸�c�^��U������5�\�zܶl�j����=�=�jww�Y���Ɨ�U�zn�wyٴ]ל��m���ȪSZ�-�[E�|  ���Ɔ����!�ﶸz>��
4�͸y:B�F����B��{M��}uu���;u[{�X�w[�;�n��:�Z�����ׇv]��/oz�]n�v���v��;^m��y�h1�͛aB�-Q���Q���  �{[�ޔ:��սVe��{��z�ݽ��W����^���
.�W0��y�n�֝k�<�{ٮ�շ�޼��f���s�o]��gV�of��zv{sw��wV�V{�lZ1�yi��0�j��km�|  ���[k\�Oz�{N��g���^^�;��kG{]���z�^�n���n�u�mݺ҅���u�
y�\�{4�=�{����[��7Vºݺ���m-e�K5답VYj��Z��  ןv�sۻ�^��^{�n�U׽��n��{���{���i�Z<�m�V�m,�^i{��nv�{��ܯp����xgU]�m��v���[w���u㙴���E�D��ڤ�k_ �{�c�ۛwn��oy��*��=��ǻ�[Sݦ��o3�;yov�Mm��6�c��={���׶�omYӵ���޻l��ݽ�{�����='��������emL�iBj�Z�Z�[-�� ���E�Q�#���t�=�{<��n���vq�k]�z{�6����h��nҀޗ�5�+ '��z� [�3����of��
�oMVe$��ڕ��#BC�  6��
t
}��� ���
 ;w�����n=��&�@@�^� z�w�������2�C��=47K� z
=U��2͢�SM[A��  w�  �u]�v t{�� ��s� (�V ��*ǽ� ����^� ��� ��������J=)N�UW��]im�e��٦I[6��  9��@g_N� (�� �ǩ�:
���  ���� �׻�R��ǽw�
�� �AU�u� '�O�L�R����4"�ф��H��4i��<�FR��z������R�   M�����@%"&ʪ� 4����������0�p����m�9�kc��[j�:=�+(�h�Ed��"��< ����{u����_�PUE?����U���"��"��*�{����~_���D!�fUE�+d��{3ieZ�@��`��JP�&�<t�����⼨�����&f1��
ktn �e#j2`������!�L*�hu�Mc����%!�;*n�;�
�CS5�ɮ��[�RU�a�X��eX)+�J�P)h�΅l^r+�	#{t�!n�<�+cK.���dL��ݳ{!�J��z��WQ��7���ز��Z߲���8��٤+�3MM�ăU7T�[�sٳ����І�ɴ���mfl7 �����(��Or�ԔS:��� ,�i��Sq�d� ��w0��	k�v@�2ay��1E-.̣��Ť���YZ�סez��jhS�0/*�ބ[v���D��5r�w\.hIe��t6���8arι)m�á��i�7�]c$h6��-�V���(��WR)���/����/U���I!�^7i8��	E�ԵX�F��2*N�����lUr��L��%Ht�Y2D���ᲄ�L��ҕ)4�ˢ��0��
�m�e�^8��A�XN��\�.���.�iv�4��A��JUث���h���4�j����c4���ʊ���-�D���a���u����\���х��e;H�h���$�ӗ��Y���w�i�pB�]�x2�� �)�����Ay@e��R�֩SJ�p�k2ɕ#�6ؘ������sw]�N�&lI$�n=�dֲ�,z�7-)���Sv���ԫk	��Ș�Ge�Fڻ����[)Sv�*�ji�3�S�+���wz�ڮDn�>˸�uh0>��	�1��
�r�!��ᱸΧ�0���[X7n�9�����,S �J�b��w4����H�2���-�)Y�֝s]Ѹ��m6��w�!KN^B]�إ�(m����6��=ITo&:��ZI.��4J��Aՙ0�P� �OUF��w�7[��B���ȭ�E��]��r�&�� x�m���غ��Ц��c5�!�����92��J�V\{�iؤ!�x˶r�Q���~D�B�9�]h�@GV���,�t�����4ֵqJ�d)�ր���v1�aף>��C\�/(���"��x!��m�{���
�`��,��p*Ѷ�=����[�A�v��Q�	��+=��-`��
��]�Ա�Cl�Bn�Yt>t1�L"h
��lCZ3�M�|l���f��E�ӥ����M��y�v[0��X��LVi�h�J�(U����2,NkR�tl�=59��; @�(ax[̓S%�ƪn�����Zh�N��$q*�,�S��D��-J"�x/0�[(�yX�: 0[	�sDR�*���ђP����{�Œ�@�n��
��R��(�Ph��[�(�䡗��D����zU�����I�w*A��y��lƩ��R�s�^��m����Z�ù��j�h�e���Sy��nQ�"��+Z��mۮ����ܳ�X�-z1+ܸ���ZFMկO�K�D"���
�o~Bv=ܹ�z ��B�A��勊���{��,�i�``9{785�1��EZf\z�U��}�Z��Q�4 �S��t��⩱Aigv��)Ik�V�����F�Дt˥���:�X��$���a��˅Z7�@z�B�jw�Z
�d��9�V��,Y�Ɏ���v0̣MZչb�T�L�vsSݭ��:�]f�"h�.EQ�B�yO.a(f��&�ͬ��3U�u�qJ��T��	���l����"����S, ��y�,-DY���P�\g����`%cV��x6��p���+#�D�ݲm*��h�x�HVlE8#��,��m�� ��H���`mcy�T��4����&C�$���
Oh ��H�.5F�(6��c�����-TR��������<@�&D\(�W�7��ĺf���lL��8�phń�O�,I̺�h�/�k/	r?�m+L��L��\$F��6w%)h*�,�x�l
0-).���n�4	�sP Z@���5��� �̖
�j�ncz	,,"D*Dѐٹ�+^���Z��$�4L'>���EHX:C���[�%*�`,vU�U���":����[�&�/k�Ss���
S4��Ȥ[���i�.#�l���*�KE]����]4�
j\�wR���z�k7l;&bb��X����Z�,�!za���@)��N�1j�JD[Ѹ~шV����G@���Qۼw�*l���IC�V\98�ʼ��Q/�*{[p�iAJ�#��v�9��[	�q���&p��o0�5��̥�е�iV�i+|ni�f��I��-9S�7dJ��ѷE�t�R���)���:�ۚ�ld�r2O%m���̅I�{;���Lt�]�;�g*��TY	"�i�I����<����]?�V-i!O2H���Lm�QH�	�ܹ4V�.�nL��`�3S�mZ�6�Iث۷e6wU@���Zs\����qS�W+4�{���@vͲ�[`aͫ�������Ñ�S18��ma�fm�:�8]���V'�k_^Z��w6�w����RR���d��i8�B�Vj��D��顿h@�5�/j�d��Ռ�6Sw��Z����!�9��T�6�����a0H�X$�@#&���x��+��9	f��4�c�5�u�$��
���ND��b��#f�d�Z��n���IR��P�]���`v)��tv劼�K�[���$�Y���A���{e�:�h-�2U]#m��)!w[�I0hY�4�r�i�ݣlPtnG�L֞e,Ʃ��^��(��WOP	OSr����M��v��IYsKn�3l^��G۩Jh���y:�3a�3�)�.��*v��i q���GZ��j�%���ѥ�9�4,� �r�A�v�H�
}.�(V �O�������<�ijۓ#2Jp	���k˫��M��9x�Ӆ�{�L=�ű���oHF��v�M�$13�X��n��Z`&J!�����W{��^G!��R����c�ÏtL��@k�w�Lٴ��R��:�$i�hjY�B������l�L:�SW���C�&V^�U��-ꤲJBF3l�-ĵf�̆Qw��̄(V�H"�K�X����`P�^�n����.%���~�ZXӧjRl�s{�ӭ8��z.�
�-�y4�z,�Zn��+*_͊Ǔ.DUd��-�S0%��-vI`:Gf)�2M&���oFhG%���\�F��5Q(K�v��]�-n]��u���gʤTe�?4%G�e�7[�:R�g ��Á�yEw�1�/��M�Já�VReX)쵕!�f�fAPV2��8H�i�&3�bY��E*b��h��`����[�(U��N��[�`i������E�\Ԗ��ç�����<(<oH7+�[QPך�L%�-b��U�k)���/Em��a1{��ݚ6h ٘�u䶾��l�*u��N��ݥ�R,4n���ْLA�4n�"��܊10,SF��L��5~F�K�lf�Y�F��bщ�.��:���F"ט��334mh�C	�X��ukP�xȎ�Y�֨-O	�V�����ܭn����Z˷��*�Ce�V��c#bͼ�����ҽ@]�QWI�ʹ�S+�W�1nЁ٘d��y{n�I�,n�f�ؒ�j��W���DtkEf��I�F(a�d���p�ǔ&m�а{����Zi��-l�7,��x`�,�Z��`��ݪjyn�hƾܬ 
h^�5`^m��V�	�X�J�J���Z:n�n��Ŷ�^G)8����ު�Mŧ`��o1Ȯ�F�h�:OP{�NΉvhdU�����
+�$itA���/kI��mCP'/@�i3��Y��w"�EH�C*�� E�̡�6��!�@Z	lQk���o�ו6-�*\u��i^��	��ܰh�קUe�-:X��Gu�k*�a-ͥF٦��	��k��.���*@34K�J���`����lt6��N���ݹ��팘gט�j��uq�U�YB��ư�lK�U��7TV��ȁ�in[M	:j�� �q:�n9r�xF�V���M�4o��\��J90�y���u�7u).!�0�ɘkJJ��u[�H�oO�d��X���;�T܋p��0�b�GR� V�S0Q
��,7Z�J3f�����2l#]J��wn�O�V���&3PЈܹ%� 4
Ih%�:D]Ҽ۵R�cD�&�z�כ)
��qO�dٖH5����R�[0�L����,N�A�*����J�:f�B� ��V֦kA���FS7���_�k�5iɗiX]����B�<٭%ݩS*��)	m�.��i���¤W,�Q���V];8����ƃt�Rn�WS2Tr��۔�����s(��@��l�����	K�@���Z&n�U+�n�=d�j�6ܭ�[ֆ�4ekƥ��/K���.�]��+p7���"�M�.�n���5�єB���ί6+H��	;���l����4H5�E#T-�J�k�E��y�] 2�(�V��]�⤲�ؖX��eX25&�hJ^:k_�T��*hV�)]�����oe��X� �N�yi�p�E7�!v3�K�![u,�&ݕZ̓��͗��ieÊ�7Y��٠r��鱶�3uH�u��L�e$k]�r��u*�,�SJh9j���;Z区�a˄��T�q�4����e�6^�)���R�Ԭ�ށ�HpM��.�l���Í�PY�bW��-ͭ�t#t������p[8��QS���� Z�
#E���n��LZ�#ĵ��췊�[�C
��ܦ%��z�Z�8](�X^e���,�&(��9�:ϤՑv�y��V.D���f�v�����k��|)�[��mPn��XI��Vrd�L�a=��i��M�a=�,�ZU�RV�oZT�B��5��vU�Q=�cFV85�x�+6�Q %@�^�j���em��� �Dt�V�n#F�ް�A���]@u�f8��U�B��� :d�6�8]��t�@%�*K�.�Q/a��ka�lX�Jj]����7)�QM�]�n�<������wp͡�R�6ͫ�p(�VhYK�� �����6��:z��܅���]�P�p��\���� M��/k�v6�8)�q���Ջ�k5?��M���Oq��E��S���6~)8�8�I�h}�,1��ڴ2��z"f��v#�I[̫��a*B�Vط�%ݩ@��-�Zx�0��<���5�na�f���1�J���#�IiK��Hr������ %G�su�2�^���e�4�c��J8��-�7��6��v��n4�n�rEiP���@V��j�lE���L�S�w�i��\��WJ̘EӒ���ziҥ�N<��A%%h���7l�#�I�B�	�t����ӱFl�8�mnc��Fj�t�P�xnFdѹq0�)�Mm� ��Ǩb.Hbz7��Ǹ��[�m��9��ަ�=�:�N��[�ՙ!�1�*��d����G�L��mt��0N�x�Yw�c��2�=�4�X�Œ��-�CE��%���C�jD@P�Z��n)`���f�6�Rbl�@y�~����=i�}s3/��$Ҽzj��ͱ�]�kp�2�:b�{(L�l޵I�X�c�!��u=40hz,�J���MB�l��[�;��*���E�ODE������I8L������r�A�5��E�Z���Z��&��+>ଛzӨ�-cz�C.��Rn턲��4��B��.�n�K7��vU���E�p�*�MZD�q�V	#�2֍�b���a`���Z��l�5�D��gNʭC˔�j�"�lB��tdnCQ$@3�L���$�-QMH��U�R�����S6��K���(�V�'��T��MѬ�Se'/
�BB�]��!������mE]�v�v��0�\S�%c@�����G(�ҫM�;��i�&[�����#	�yGT��;��Nn![�]bVe��y�R�QF�&1�S��f�գ�Q17yd� ���}�r-LԈn�A�D�{P�4੤iUCU
7[y�J�G.h֤��2(�˂ͅc0RƳ.lQ�V���`���B��]�y�wH�x�
��e�4��nw����)KyY�B�Xw�e6-�Bhkej�L�s.�e�/r�e�nI���O]�0��AL��L�T�m�]j�\��+m�&����"h�&�(̺�$qQ�-1� 5��ɷ[%��e$2��On�})S:-^�D8�۽Vfщ��V�Rf���UV�6�T@��e	
���͌�.f�A;�tr�ȒT1��ڂ�7ia�q6mVc���(R�!e�C-�d�ʫ�^����l�D�*��@Vpܷ�ջ��t���@���re�!ޡd��!�ٌ1Y�FӫIE��+D9jh�9�i=���|rŌ���V�~I��޻��fG2�R-5�����o^�M�ݧ��v�.��E���
�[��V�P��(�4b��m�uq����-ҫ���J��e;�ƥ�����f!������)�d�-�[3%n�`�
Z�$]2�㭗em<b�	�.�ֽ	,�u�@ C��miBU~#/Vb�曚�5����^�H�x4��4^���r`os���ړ��K��y���$(9b�c�cv��G�e�&j���w��M�{&J�YD�҂����.��Kv�ږ���*i.٭��F�`}�K'/34m�I�Y�i�A`�[O��m�Ł�����u�
T1 ��A{�/ (�qt��չkd�r,�j�]��ϸ"�v�Dq����RS�^s!�U���n6������J��N��4�pܳr�̙�g�:�y������@�;
:ƞ�%]�c+��Y�9��w�ԝ�V��h�m�ޖ�֎��!:�5�!D��Է��GE/�B�����ۥ|H63����Ъ[��R;r��Kz)b�N�E�"[�ﻆ��,�I�F�X���\�s���5�V��}�����􂰞7�[cVh��=��\ѝ���T�y$Zv�\1���Z�ǜ+�m��Ƅ��]�5k{��N͊���8�Ե۬�f�N�Bڌ�.��R��54n�Y�es�H��˷U�l�տ6���m�s�;s��3��ͫ�:Z��Yx+zrX���Xj�W�:M��G�s�>=s���h��YOI�c\�G���Z���_.o'W
���w
�c#b����pP��w|y��B�V��<ty���R�Q:��*�.�ΝC�}�����T�����Z��.��eη�'WZ��3"`(�؃�����t�t�59�%��t�u|�ZQ�34�O
�KA�Rv���VT�}�";�!�P��5�f�v
�z�I�x���魬͵L��8�z��R�R0�����I�X����ƙ��)��{Cz��ܺ�9���a�燪h���[2��a�=.��REɅ|m=-%Pma8j���3���t���:ٲr%_n��Wm�����yȼ�c��>��v#߉�Ⱥ�)#15�f�tѠ˻�Y�M��N�I���Zs�L�u�ؙ\/��Ã�S���*��7�Y�$d�z\�o#�{�e�R�s�#��<U�>�^��Z,��zW&x������m��<mG������)��9[3]H�'lG�5J@��r��DoP<f`�C^����쩖%6|��� ���b��NOie��"n��P�����-G�\J�S��K���#���p���gsrL�T�&��I��m=��U�=���g�ѝ&��ApL�8�kn�ŎfAl�p�Xk���K:1�����1j��L�{����򵆝fs�z{���xt��[�ߴS�#'�5�NZ<���*�/�=Ͱ�[����ZM�;d�̼�<��h�H�{c]@�+�7+�f�@I(.����Nv�M�nK�G�Y���q�#��Ok��K2d�m�v���E)9;nD��P'�m۝WY�Y�)^���ݾa�;��Gyn��f��4��E��.p���Ѻ�X/ё�s��g�wf�7�au��_&�[��*�}��y��;X ұ�VQ�y��ܙN;�0��r�{�{�(3"�$�lR���┴uچЂ���J��þϺ%�0�)��j�d�اE�x���;��[@���G�h�fi���"����&�.�Jj�������9������$q��0[��h�\������c5{�ofU�s%�t�}�����r��N�,ɂ��z����b�����ՠ��E�_7�Z�8��ᆯ��طX��\�h��nخZU<`�ϕ��ʷ�2�9�B'S���$�0\��m�[YGv��k��B�u)v�K+w!t.u�0\r��֟NO��pq��Th���:A4;X��f���Q,'�}v��n��S��Pa`]��O^�������"X�]y��\#ԗ]I$�L\�c��{����nӾ0B���s:[[v�+
 �+���}�x��Ea�j�/��g1G���G+/�+����Tѷ���Lc:bߥ����Ұ�)0 v�3;�<�E� ��y�Tظ�)l��E�ł�n�+o�H!������	�����}�`��8��eu�9�p5�^�Z��{��9���t9�t��Q�B�ǢWu�Wf� ��[��D�I��u�9�'�+�da<y��s�/�ҧK�pI	�����,ͺc`�P��t��p2����a${�n�=d�������ZB����7��F��RM�~OqW�¦�s]���\r�=�3l;�\t�!MdSi�Uڲ�,�+����8Q�G��o����#��e�r�{�a��_#�5Û�P���{�\��<�e�5�Y��S����Zz\��V���)���v9��E��}4�a�q�|Vf����K�0�T��V��D��ev::�6M����/p�:�[4w2��|w*���1�W@:K; �x�<N{)�J٭��*Ƥ${��^����GEVR��Iā ��;l~u�9��ER��P+��v芻��"�Ss'1&EL+���|7��ڇ��Y����dsM�]41�uڏ�̩�|��J�N�̴�$t�uR��5N*�:5��=�[yN�ŰS7����rlb��,��z�o��M���Ó'!��xSi�˷"�j�'xM�z.ZZs�V��t{OU�Lk���͎�%5y0_,=[㉦�V��)rWgU�ul�hI�ˍ���k���ZP4��w]�L.;ٶ���Eo>H�w�hT,vd������K�&�[J9���}A�]�e��m�+sn�72���뒈�DN�k���J�n�ۥoWe�FPV^R�*�:-��C�������Yw�KD\K�!�g�f��!c6���ǆ�Sm��J�^��iIa�����w� �V+4h�7jT
̬dG��^.���MvPd�{]V��m�w���{��2d��f�-û��Epˏr��q[؈0�fD�n�\i�n�ۂKn�a�N��8b�8m�Xv�P���������]�8�SHnJU������}������w0H�.<Նƃ�Kz��5��w7*�AMn�h>٧[���(Z3������KoF'��-J�Z������u
��%�!���v��{fR士fO��	��g�״�Jq3��7V%���umu�6��r<>h#/�����"��1c�̌4CF�̹o��$n�Yj��GQr�1�.�tm��	��N�9����<2TR�=�_2�v���|�ތ���	����v�7rb�i���0�/�Q���1ڛ�3P�ZxS����R��0�B�乩���cz`�-m7��Lv��<�MV���N<}��eG,�u��N�:��e(mrxrJ����Gn�X+���e�4P l/�AlrD5l�w,S.�Y1!k��6���|�����u`ڛ�h7m��r�ۥ��:�����~�؞.��1ի<���T�D�����&��kۙ\��ՓD��B�ܸ���F	�<	h�4�� g&2�h�Ank���Rܯ�;�f��Z:7���rXv:v$�敃�Y���a�iF��J<	����x�IVn�u0���y�sy��`�i6�d6sF>n�Ac�	ykU�Ӻ�'"\�>�R_|��ʾѥ�}L[�p0�B�,��6ġ�7keøo1�;)�iEu���X�,)��!�Xkx�Y�[����#�{��0JD��N0KE���վۢ�*�Bs6S����5g�zb6�s��+�z�Æ�0����`ͬY��2��y����T��k�aMƧh�����W�"����#�kw��Z��/l(�Y��ېVe�@���{Cf���(e���G	F��J�e�s�-��W^�J*�w9�I[5k�����J��\wv�n+��3�6�`���U-E�%> [��Ϸ~�ޕ��%�������	�i�%�?b֞N���475Ȅ�Ն�g
蚽�תS�N�-�r��l����b����iL�v8����K>�5��ϴ|����l<\6��(���f���n&���J�2����t�+j�M��:�N�3�H.���*���X�픘Y��vPoLZM��`)��S��k �ɄN#cL���ܕҗ�ۻ�06�?vK�k��on`�W�i���c����dѱtr�k6��c#sq#Ӻ�fF3��b���[\fӫ�D� ����i�4��L��p%Eǵ���u��S.�y���y�i�8*X�'�떘�3�w����.�����J¥��yop�Ӕ*�9�;� f�F��-5uӁ���L�m#����Sc�%��Nt�q��\��.Ͱ/��FM����Sn�ݕ���� ��_Ak��#w��܆���>��V��X#le�ԋE�:�M%jq��8:�Y���-�ٝVo� ��)�Dڦ�[U�Y��Da��zۥ�@�� /��ھ xnoH�4��'}�.�2nr���b�ˠB�RE}���YO^G�#V�P���;�@w�&���޾�!:�|^:���r�#y�ˆ��T"5�j���{��>�b]���	.H;f;�KƆ3�{Ֆo9���5��SYÓ��pml��؆^�e�(2d���T^K�쾩%m��#5�{�R���;�X'��A"��f���(�z��@�Eg	Aแ[jVs�Nۜ���s��y�`�iNz�/���#۳�eћ���Α����NV�@8B�X%�]����5�
��̻���޳ڈ��7iP�'�k�Z"	u_7��	kX��m�Ԗ�%4	�5g.֍���i٦8��X�죘$Q���Z�9w(<����40��t)'3ْ���jgM�B ƃ2��A�V�Yc�WnpRnvg;��l��PCF�ni5��t���F9a{����Ͱ��5;/$O.4W'g��J��B���	�)]Ne���	��s�#v�5΍�R9���w�YW��&;�A�h�e�\��Ͳ9ԛ)�-���X��}���;�x�*N������ɯ�� lT6��Eါ��+�[��|�śƑ$&���R̦7R�u�ݵm�ᙱ���M����c*��_(��b�QIK9�K��\f�Z={�Np��}�[Zȭ�_�g��Z��9"30Ŏ=���ٷf�Ė��΢
�k��q��v���J �vLHgG��
�.�cT����йqyX)�;r��ǩ�6�^i�]�Tݱ��i��aZef��`JU���w2m٠VW)ʣG%օ���/TK��*U��+*4�yes����<�oUvG��z�e�&l�9�R��P��������+�E],Cj޻郷�ʐ-��3ͱxh(��1�x�����k�:C���UYL�Az��"s�v裖P\���Z8Iӳ�7���U��D���.��Lt��e����!���6�@�'�c7r��5dw2�|�+]1��v�����NV����&kc��B�O�ō�����ul"����u�L<c^;�v�ݰt%�8,S�,�����/����Nh��]��7�2�]we,���>T�9�iSYet��ٵ�T�q���e\	Z��ðod�L�ʥ$��4���K�+1�P��p��d:]��C�|82V�ZZ6r�:�*�F�G�kNn��k�#��`�}M_&Z˙�b��7������sd�hv��»���Ҹ��f�T�E���P�_��5�+��"�5�wS{@�((�R����+M����׹t#�mҴѨv��;����S�Â�nm74t5���-%t��ʚ�_^#A��Qu�#��VCKH�X�Z2���dJ����܌蔪���].�I�DP� �h�fI�+ �y��~ʱv�vE���R`l;B�^h[t�E�G�+aR�p춓�w;%Ѯy���l�审�U�m���m����H�Z�/B��5u�+'k6�;$x�|��v�	����� ��f޺/�aNizŋ響`�GN��V>L���Nqﺍ����]Lukd�V� ��DV��2p�*����%ڽ�qQ���Lb*@H��Ez��5���ls�I����z�N�8���<,�4-��,zxZj�nm�v�|i�r��n��r�e�Y=���X���ZIƩ�Ηp�]�XLWrml��E�i�NM�!G9��Ѯ�[�_�X�b�p�o�s�zcs�-�L=-h�'Q��xd����$���J�0�ɂ���D��F�B��rGK��l�ܺ;Zr���H`uyO���2�|�v�e�9V޺L���|4�U�H;�������0W��x�/pI���pn�`yɳ+��QTF`��.�8��8SR�	^��6�j���G�w��ݸr�����˽�⮲�{z��ʎ9� �����7J�-�+r���1lp�;~^�G��t��u���zX�5��FG�೎��`����Ŗ�7�_^ۚغ1=��lu�`ZѨs���f�x:�Z�v��Ǧ����v�l����]r>�t�:��c�3�'���#�Vs궈lW�5��U��SR�f��9�pǝ@����5ݙ�!�%������5�h�,�b.f[O��-�OE��(Z�3�mjkX:O�7�C�WVk+�v����Z�2���t�79J5�o��A��+�� ��d;��b,�m*�Ϡ�d>�C��1X���x�=}$�/�]�/��܆�%C�;Y�V:�]���&a�m�X1���ߐ����gZ�}���O.�[����F>c%T���#�ms��Vɰ6�^vܬ�p�|;������r��R��sEפQ{����O}�5VN&t}�8�X{�o�z*���ŕ親������� R�uN�(5'wg3�f�5"1�@7O�Dvxd��S��]z���Օ�ow3�6^]�.��4�My�Z9+�n�U��KOK)*g���gy����:��zgG&�Z�Y��JǈX�+ffI�.�[��:�F�wvv �r�;��ڝM�{h��ړ����8�nr�-�WKԋH���X�*g	gVӒ��f�i�6�:T�3���]��tn�}����3��	h��f�\WaŻ�ХlR�bU��>�m7�$4��嚪�K����9��ߢ����}���� ��� "+�%��~�w�.��Ȱ�Z$c��'ݵ���ŦxI�2��J�U���b�s���9��}�V>�v�g*�y�I:��	��x�tG�o6�2�5�Y���]��WE����WX�*`�]�9��=���A��a�[3��%Ր�!�V�Ȟ�����7�:|��Nv���{Ht�E� �1�݊iTQw}v�M�/�0�j"d���TC:`��n�#h����V�822o��g.�E�
ҳ1S�=��`�X���p��2�#hk��>4�������ޣ�>��k&.{or���I�n��Bn�P���zȥ��7�n@�W�p.."��]s<N�9մก�b���`m���nl�a��7�8V̫��N��mt�1��gU��V�%�:��(k虛5eM�_u.6%����Вy%�c\+�(k�B�e5J���h\�3ب:�i�::�� ۤ; �F�ߎ��[�_`��e�S�
��W�[�xlŻf�fc�x�q��4X|�^�X;e�E�N��rY�KPM'G1Ƌ�}@W}F+2�+�{����v�yR巜*VX��pe�C��c&@�bǽ�����՜���L��V�s8��e;<,@�<Z�ܷ!��i��+;:��ڌ��U��j��^�:l�έ��oxBkCA���H=�P�F��Yݔ3oi�iu� m��l�W�-hgtǲj��GK[����j�b�P�#���QFl���	1#(s�\�6�_q���t�y�^��#���=3�� z!�k��j��:�N:�LR���w�ӯd�G{u�:��;E���S4��R��m�k.�9���6�f�g@�� ��0��&�s���7��2i�iO8&�������y�tP}4U�/��F�8'H(c�Ԑ��3ظ�Yk)��;�I�)���Ą��'g�/8��z�솠���m�ȷ(���[��Y�_�kL�"�;�I@�u�i�Y�A�rf��P�i�Pq΁c�0f5�V㾘2f�YVGjn�0�|k9�����ֳ{�RJ8%���{�+ ��X�c��J��F�H�z�X��R��>��.���Ur��P�Q<CA>�5�-�y�9�9���Z��#�(�F;��))3�ܝ�O�%,���Еj�k�<���"T`� ���f�w\:�푊Q͡E����1��<��]rZ�L]�	��w���*�7�(���+2wOOL̰Eftd��'k��Jb��.��Ƃ����}4Ė��ت�Y�L�E�
x��n�c��t��S�0�T���,�w3�<���lm%Y��D���_llOgu��G6����Kw��tm -�Ƿ�����a;7��v-�u/t���kb����!�p�I�\�����kgq������k�
1��l#|n�%�f��8�ڬ^r�IS�KN�V���F�=��K5���f�	]=�`�+�WԹC�p�7*��W�B���%u�q�æ���aoխ��F���ޅoK9x���ṅR��s!��rw�
�ڔ/�
�ǲ��U�]�+�*k#�9��pgi�~7��݂I���D��9�G�����]�+'j�w�Xy������������� �s50s���<�r��N����}�S�ۛ�x���)Gp��%vm�4�ɖ�ߝL��׻�n�r8����*��Ӄ7��4g#��*�S�ʯ��)��\L�����KmƸ¹LC�Z�X���j���]�sk�u+r�7q_[��j��}��ͭ{��oj�<Z��f d��'�Nkf=�׹�]�EK��Wvg
jX�iT�Q��{S�_T�r�N���h3܍*t%X�t��vf���7v�v�f��1^��F.���=�_-����ڇ� �ȥ�V]��\�Z�@��[I'\:T�fe��@$�VkP�� ���+{E*[���O!���m/6/�'�_a�����bu�a�чpѡn�6&WA{K|�� �x�}�Ն�y�S����!�өM�Y򡶤�s���E�jf��=�y6m8	4�GV `��V����z�
7)�Kc���k�6������5�=��ԍV2^�2ff���QkvA��uػ&����- ���x��#7���qT,�E���{a�R���������H�%�,K��[��;X�O��͢���"�b�^m+�r�빥�f٥�i���2):�i -;�\��b�]u�-��ޯ�Z_NT.���#�bt��!�Җ�MNO��\�΅�Uc7��E��]���A�	g>�:4ձ�]_�a췴�
�*Fd9�fЈ�|e�y%�͗&DBbC�I�\Gq	\Cm�M�RЇta�
ܣ�y�7��{�@!������k.��2��ԫk��6�w��4VU��i�R���<��Z� b�2w%���M�����֫w�)��oi�j
=6ܰ�6�;2�)�Cr�U�oA}h-�5�{�V����xٮb:���2��	�
|(�jnX�w1&��[RB�_K�>����Ţ��z]L�]���4�ٰi��?@���Eb���IɃ+��}o�c��>f�=R�6Q��:�\�[ˍ����s���(�����r�з-���3��s��R��-Zgv�͌�dm��y�٣"E�ܱڌn3�YӤ��c`��̲��Ij�v�:2,]F7Έo��7����n����Bpt����^���;(]�h݋��+D��=��A޼�ږ���x5[0��ut4#�I�;3�t�.�_Ml�39�ãS�ר�W�j�W��f죐�oD��,TZ�V�<
g^����bxYc�ks����&5Ya���E-#>z+���î�C�0;:6*��0.\ma,��m㺎�D)�z�v��r��ع����c>���)$��;��4EetJ'�@���u0Q�/UGO$zm;jvֽ�n��u#�۬3)ev��Fm`�6���R�y�XA>�if+�m!�"�9厼"��bj`�F��9��(��-w��W��[a�N���oZ�ۭ��ᵂ �w�ݰzZV�)�`m���eh+�&n;I[9E�N�C�A��nևecM���;#y|�:�5s�2Ia5j��*�*�\Ok�*s����c@�m]��# Fr�u�]�
��Ֆ�@�^��WE��΄��͸1<Y>.q��̓,��x�7���ڡ���Vhېv�s���\Ϊ�����ڊ�π�m5�l�,٣d*毉E�X��L-í'Mc�;�A֬����vT�k7iQ�cv�df�R�m�
0�	9jov�i*�PQ�e��`�s�si<
N����Y�ȷV1����c�8�pu��{�\�j%��JMi0��yY������0�����a�؞���
�SC�%Lׯ{l��|�3M_h.��2�sp�0�ϒ8J�5�wk��V\<Wpy� Ӭ�;������F��[ҜZ�s��bm>?v�Ȭfi��u�4S45_NV���[���5@�l�
�Iƫ��n������i�Q-f�7N��Y� �2qɳ�3(�ɋt8�X�Pc��D�q�*���̵z��BC��7�[�V�|05n��ʮι��r���v	ee�M�=z��uJ��12y�3���2Z���%Y]�@r��K0hD.��Y�u5�y�X�ՠa`�����(�g�eX����I!�h���h-��ݕN�Wv�fgPb�F6�qr��Sw/�KЫ0[�=rmD:���X��Ɩ2�14f��[�:��m�\Z��; �T���Ntg�*���Ѽph���ɠp&�La�я0;I.}i�Z�kq���]�e��=�l�j�Y�&�}��밨��d�0�.����S�P�G��^��,�B
�o�^��j�M-4 ��1�Q"_��a�ڙ:�Y�A>ݹ��`�w�ò�B��XB����x��5
8���t�G���d.�os�H��ۄ�՛�W#bN�砉�Lx-��ɚD���6eܗ�Еpk9�l�3\J�f
X������mB��=[�,�,m����Őu]�-Ź{1�F�[+ �$�9�/1�`RKx�DEc�z������^��.,��{�亜bʚ8���6��[T:��W���Ի;��tK��c���s�s��}s\�p��R�<����ϳC�a᫄e�7_l�w"�
�vt�|��%E"����|�T��v�I�归����h���j�%$����ů��_����e�B'	@�����+�o\l�>}�Рujx_![WN�YL�FѤ��Q�u�,6&�W�R2�e�� �S�BQV��KC�K�vg*�Ϊ�-1B=b+��om_q*XIu!�i��Β�Uw|�T�j]�Zc�qw���<]VX�6�E�w7!���r;kIg7�xL�V�ɦtj:j�M��Zvs����6A��f�$�30-4��zL�*���v���)�:���ZUխf��i��b����ANy�Ygbd����[�Ҳp鵏��E#@B��f�b�"��"�9���[��Y؊%Z�	ĭ���8�9�*mI�*M���F��Q�V�GA�D�1u���1���m�\�͎w��"���RT����&�:��RL�7E_
�Uo�`&X}�h��	��5���r��-���Lh4c�Z�t�73�wWFx��+�j�4�r�7��XkQᓶ��s�e�*f�-F{Ek��ϒ�\wg� ���꽒؄����oZܭ3t�a��l��Sp���v8TNC��3�q�Bb�}�'Vl��ےfa������-���Y�K]��+J� ���Xku�vO�2���z4�Δ�,������rP�s Y�0U��&#t��#�@�yٺ�
�ޱ�^2Ù\0M�=�%cϨ�F�P$X�d����b��-�Z��tͦP��o�'��f�,��[�(�DW:��[��r���VaN�tP�'V�tf$U+�eњv;R�d�*+�j�V�I�p��%qՍ��������&���T�>T�۝ܖٱ�d�jb��7,�g4�'p1�����M&!�l��})�Z7�8��ӛ6:}����n�\{�� I�@���]u0yVl}��%� +)	)O`�i�Z���mo6P�0[܅�wE"DB����v�p�q��Vm4�=CJ$� ����8.٣63��^����"[���ꫳVu��_BND�j5�B}ֶ!��`���e+Qc��T�Vi��L�qg-����C�Tv��é�4rԯ]���������蹥b�_�w5�l�܈�Us�|���E�7H��ٍ?��ͼ��C��t�x��3{v��G������B�ja����R�ï/�y�7���U�c/�f�?�[*۳�f����I�7sD�˔������U���=VWU�O��r�ª�-�I�TEѨ�o��t����wx	����9����SԱ]�)ԣf�zj�Y�����D�)SQ&�q	et�<�0XrgN�[d���e:�t���Ʈ�|r� L�DZ	Nܰ^^+h��}�qC_c�(.a`1Օ���Ӷ����j�lh��od����hǳ�fT�z��5؜ګ|$N�_e�Αm�D[$ƥn�G���l`KS�i���v'�4j�B,�Ӑi�#Y�CywoM�]�$����RMG:��y�'p<I�c�����Qn_)8��>�ïK�U����Ƿ�䮮����5���,oC�bLa*v��G��&U������y��^��B��A��<��:���f��é����Zww�V6V��F�e�y}���p�s��������k��&�����oVԿ�!}�ЊsӼ>�r�^�\5�»l��� �<&�J֬�[�T�0f:w-Qvu��R��H�Qp��*Z�5�M��F�*�ܙ�fL�"z�7x� ;�h��:)��ͩ���H]F����\������n�bY��^i0rE�*��O�7��E�=ʟT�u�Ļ�9D>�K��k�45�)��*kU�	�M���9N{s��T�"�@�ݷ!R�7���-ԑKb��4�
\�!�f�Q��3�(��e��۠s��]Ҳ����T��' �%��B���Y;c9���Ѭ'�[���$}��C���d�
�����͗�Z�1l�AN�ݗP�ć-�lÙnɺon�x��i�Ĭv.a�1����by�]w���R҆�d�X����)�5m���4]��.�&� "�������w�m��y˕�n�C���G�>�|���*4~�"�m��'Z%t�}�Ct�µҺT"�^���T�:d9/�k7���7!�����2���,�H�7k+C��{R��el�dሔ��n_�.r��6r�S:�P�\Gs<�Rl6^���wY��Hػ̨�l�Y �Y��/�r��Fq�h,���t�ڹY#�<�&��%� �a�F_kYSu_3�s8*4dMɆ���	.cZ����:��a��5[�}�K�\�4�c���d5��9u��&�Ѽ�AȣZzB�GjP��7]����MO$J�c�m�&�R����Ui]��U�:la�z�%�*r:G_a��f�c�>��ɩ�Q],E���ZufCAgq�H#Φ�|O`�ӆKW�)Ǫ�(.��&q��c]D��
��1p����rm���w�8��[]C!��
R��]v8jc��s2���!�e�e)����r��x`�A9(pZ9�N0�n�� ��k�&-ab&i����M]����X��_X5t����<2��i�]Ed�2s�1�`;�w$�VfPZ��i�4]��VP��wYv�R��̧rZr���h�w}��[����I�*��aR��mś���}���^�W�4�ၰM�lT����C��Wtث�r�H΋�1�+!������ɔqg� >���}�Q�gG���J;PF�}3�e�0���JW-[,�{o����	�oF��BCI�����mq��Vw���z�J�[�N�-����T&��|��3"��.�6�{iu[�֩C%8�:E���-�hC�t�:ʲ����b�A�4�><gla�rV�Y���Rpi[�V�U5{��ۮ��Wa?n̓u*�o��r�kF���hŰ��I�V��ف���s��Ov����+��`��Ժbʥ�E��nn�i�ido	�tq���B6WlF�ꛔ R-,�ssҝ�f��M�wX�VN)j�V9-ʽ�X.s�ܦ�P'a�n�#Jm�tD�{�
qpެ��8Y9�󭦳yPu�0�t9��hSQ����&� �g:���s�n~�y`S�Em�ڻ\�9ú�������t��ᕎ�WU�w�n��QR�1�_gU���f��N*�U��%��)��,GЛݦ,ci��4�L����CKu�V��.�݅�kY[}Bd2�e��v���}��ᬗAid.Wg��JE�e-*�N7��������
WC�Ԑ��'��`8�#@�g.�������U�)Ƌ4j�up�Z�J��~E�X��!uA-�cvn�Y4��ĬS��+�H��u-e�t2uZ��mPG
6I���.��i�w�<$�u&��Vt��)6�R)t�m�]�5L�w9��۸���ӊ����������������QUT�[j����N
 ��O
��
*$��!Ѫ�����H�ꦧ��X����4�A�lL�4SO#QQQ-Db�j�J�J������[S�QI�O#EL��2E1N�L���b��
Jl��M%UA�j�
֪���"b�������#��h���.c��O3�"���"�� �b�yW.ITEUTQL�xO1����1��j��gUMEUKMPMZ�S��DV��
#C�m\�&bb��:u��b9�1D�Irm���"���(��X������W--mh4��*jjj���*��ETM�EW,�i�QPGc���w�~�%řòp�w1ؚ�o,����t��I�/3u�f�(*2]Ԫ�x�+r��m�8W���6���d�;;�7�eW�3��FB�*G�ݛf�i�����s���8��>W*��OL���m���3��;n�ᖽ��}yS8	�>�4,7Ʒ��z:A�)^j�u���A��'��r�?Dɛ�s�Fߛʨ�ix��p60�q�"׺UK�5���}Z|��y/��i[\��N�5�����xE>br79�;�"���*88��k���Վ�xeqxm6�mㄹ�>`#�d�[�����/�˪���05]�m�8�Y[�u��6[��9wQ{}nvם�E�]�����Z���Y�6��P_;�XNy��s�`��ˇޙ�1�J����<�x�1��'���P��Ap�Ȝ�f
[&$[\����ՅLE��7{l��2�ўד���41�$��w�+�ΐ�A�n��^|d�\��{|���<g��%@��t��~ˆ�_��1�ӡt$tdp���dr'��b�*~�׹Fd�+�+�>�ؠ̳x��c�Ie���e[ۄ/�3l�|��( h�cV��[K��S��dˡ���B "�4A��)�Uj�֞�7Z��S�7�n�d���k��n�Xn�t��4(�S��GZ�%�ֱ��g5�vπ-����(���:�N��䮩�m]Ci&� uA�ܡi�΃�B��෨�Z'oS�K��	�\meر��M����|��\o�n�y������%��-����K�B����4��n��:hX��c[t\m'v���a�m껍Nc[�/���o����A㠴Г,����z�u�9�����13A�C��;&���cP��ۀ<55H(r�ǂ$g�M�y7�j�'��h���WdG��*!i��f�"�~e�o7g�;���μNn!K�ZQ�ouGKd��!/�~������7��S���;��u|;�5�9&�j�0��p%Ŝ�-�KMR��x��:�GG71�އ3Z�P�\u?���xA�Mm���r7���-;T���f�_��#�����U�c>d�4���(֗�Y�i��laX�����+=y��'�
�^��bp�S+�z^ذ3��B��d�U�Em\�3%���ܐ��zj%K�+�"쌱(n%������2܇�3���{*xe�4ؙ`��a[���y��{l�rJ�1sR���7x
f|{�ҩ�Is'l#
���h6Hb�`�L�[��W�S���=�S��y� ~<��:�g�eZ��!J�9�J���o�θ���V�-��e)T�R�l��QL۔�Q4�6��,���j����J�M�	���|��ބ�C�����+�����_Z�c��.�L��G�2n��ʡ>�w��BN�H^�DO��v.�K��+$m	s<kӨ-��T!�|����3BP;3޳ů]%���{p
u�@�"�z�b$Ңtz��ȟj���zݫ���N�z�������h﹮��~��g*�/��<]<Dep���+���Ѕ��'St���M�OT�˨��ˏvG-�`4!������)�@Q\/ו'QƠw�=[�}q"J��xH�ӑ[u�%�/�Rǅ�ש�I�6��A��BW$c,��7��.����BI���5x�� t�4N��~�>ؐ'y���g�t�;�wůl&��"�nU��$M%�0F%	�)���H�Ҝ�X_�'�f�����lW�
a�}��w�lV����{ޚ��b����Z=�Q4�㢝#�l_b7����i<�C7g�ڍ]E�,�|�Z:C`8d�%�+��U�Ď�)u�79X\�K��tz0fGui
���&�xhf�P��H���tQ���q�C������ż.��J��/b��ࠝ ��g[�fO9�g�}����pH�QL�i�
�̮��Z��s�����8"ۣ*Ɔ
�g��c$���5x��O��)O����12�A$�P�q�4pJҥ1ݣ�8��Uu��٢��gOU��NZv!�'i�YD��ڄ�J�SZ������>��b�-j��,p����ս���rS�ӈ&u�.�c�+cc5gl|��d��C����}>\��m.���g�	V]�	��~}�<S�s�� ��k4���J.%b~�BbC��E�M�`�G1�Jv��SJ�U�z��}Y����Qr��sot���XK�LCG]Lov{C�W�x�����W^��^���x��t�:���:[ N^�暞e��H�:�O�_Ni��5�f�.��y�E��f �a=��x�1������ʨ8��F\�W�1ˆ���.�+�j��n��rƺk�xf�Xm��]����'B�1ǯ�T��w��!���Z�D����=�'�2��e�]�X�o�;?Yy)a-���A�WI]�^�����!z�@�eE�ś�id��j;+���q���3�I= �H�Wqۭ��Oa��.ȭ��B��7�ѕqݽr6b��/$��y�E�n�΄'�r���(�B�@!t���v��;&s1�)c�̭�����]c�)����ͦ/�}���.�c�9KL�yr�&o!h���Ju�&�\�P�t�iŕ��w{�Q���M9��Q�:����d��6��ŵV:��:����6��[4�a�!�&���/���1��]��Ǫ�)��+��M �p�L�;t��\�\�A�;>J!���T��SojCʩ�V�e��6!��l�ͭ�N�"����!ph+Ne�9#�zQ��+�mR!���˹5>�G�����)�=cep�Gޤ��C��,��w�����������骏��Sm��!m�>G!�>��B�]s��8�vO�ϺY.�4�5�}�g7FD�$��=��{0*!Z��'�1ԁ�WgdW�b[]t��3�U��8!j���ws���m�SC�$8Jp+���������v6�:���5��_�dU��ꔶtbcn0rtf�cx��s��������^%tC��\m���³մeH}7=�kU��{�Ck�����5�����<"�18�`�TLux]q�/V+��;���=xa�oY���Vű�['ҎC&�^�DN/r�Z�o�Q�v��n)�p��1�3-pڙ}�h<�;/DB�Pp�c.&iW��J��@Lo��A֝�K���=�1*��%���Pmv����T�n����`��	j�;\��e�]c�*�`�IY�䡾'F�,����u�G=�x+}ޡ�g�YZ���~K�8!�����K&.��0ћU<���3��-�.�Wq�r�<w�v�h�Ah��f�x����Yb���._@�}b�\�˰#ζ�d>'�Q_@
���:j�P	z4�"��l�^r��ݳU���S`�y-k���j�K���q�\�;cC%E��$o��Es����:��}�>���.��G�9Ǫ��BS^�!=u){�����h�K�N4�=��P���F3�g���$���S}Ǝȉ.�
M;zZ%����eE��B�Ͳ���( h�% �g>��*�ƹ5��-�g�`�����L�ۯ������,v�����o��kθW@��,M��c�v�zǦ�K���X�PTo��w�t	�s��~r��ⰸ��s�M���X�`},߻\��I�lk�n�>�R��Q�A~ǖ��^�O�4*��9�o��]��2P07N�7�/پ���[���
�,��>�3�F	���Yq�cy������3����(Еn3%ʫ����i��4�-���]j��΁�ꎯ�b���dq���Q���T��*���=��So��Y(�71�C���$�`juE��p⡋�͚��������;����
C���Ŗ�_D�.���/0��X�5@���&w�.s�.�vd�|�yJ�s2���.Z�o+;9
��S����;��m.ʕs�d��'H_�<2��cR�V�ϫ9��|�6Mh��Zˈ�c��7x��2��T`nS����Wr�j��3�ںcy�i1�2d
i�9^n��ixU�DF��������{-g:�,L�%{,=��jg]�;�LLX���W��8ԫ��c�t��Ad,�na�|5�rRX��̢��.���\�^�DD�:7�o�#�S��-���9�GjK���n,BJ���B����?�Ua�K�N�#�{��6��/�ż;�c���v��Y�ک���@k�ءz�>��NŢf�=���̖��=/��T�[��u�oF+t�H�`��!�̽�
u�^/H��#�}z���b$�N��r�4�~�ڃ(߳A;��j�U\���k�/�A�B8�湞�Ku�9�#��<]S�AË$������w��@���2%'.(NT��Q
 ;8����4!�o�<⭟'��R�#�Y/m��E���
��<I�Ehi!������5Ѥ>���祍f�CwK}<�}It���M�J�n��_���=�~(p�{�	�u����}�3���:�9x����Vwg���ۍZ�����^a�Vl=�D���|&�lzk(<�Qn*�N�i��)P�e��Yǋ����|�\X��X]�������\f	ǎ���e@h�N�N9n��,�>jv�ǃ"�m����[������+H\�������d�v�����/�pJ$���1?���6
���?->ǧv3"�/Ia��	uʉ�֮��Y�mex�`��
$�=�%l�0�&tG�/}ꙚW��g��n�p{�4��|�ۓm�h�6�z�`��"�G(1`T�V�kt飗�Sҙ�g�r�T����v�k������[ [�BGbvQ&��sXgN����c��KI�_y��ӥ����r���2�n�B����\�S4ܰ	��ܷNz�=�/k�u-�v�Ae������x�q���|,z��>y����V���T5Ɨm��hQ�P���mL1��*U�&�P0w�9��S��1�V+��S4�V� �c7ʝlS�.�!��^�b:�`��ׁQ�)�����D_����[�����	(\~��"]�8^��Pv)�Y9$_��W�W��B�5ad��]�Ge2���R;y�{
�u?��2�!��Q��}Uv @��r�FLr�Ao�.�:�8m��q����а��s��zhf��0��RU�i6a��ݦ/��ν�� ����n�t��%b�2�!��69�#��u۶��rm.�%��~s�Qf��k�I�jCۢJg��h�RUn٤��o9�mf0�ݶ]����خ�u;��|6��ٽ��l4-� �q�����E+��X���4�S�Y�q��
a�w��"�L���k6�ϘN.ys����؛���ܬ5DD�w)䥄�he�z�2fP�}�����D�aqߔ��3*�>K��9j��g����\(�����|t�̪��k�̮�6J>1�b��QG�+�k��h��o�����c��P��y&; �eFPn��B'��Df��B�rz�Ȍ۫PK��a�xz�h�9�AW�gt�$nɁ�����W$���u�@y��Ż<��Z�ֆ[�;�ba�;L��gcy9l��7�񶐸���2��#�uhP���@"n`�A��W�D/����)�=p6XV�G�Ki�����E�z��dT��\gkB�l]���sl'�+�u�HwT-�%���=�)���;�J�1p����iS%�&�s�XH��:�f�f��m�",�#B'���e�D���*�Y�Fk�q���+2��ˑF׎b�S�2��@�`ap��d���NϠ��ř�M]��]�� k9��ӝrp�ֆ[��g�tM�0q�%���o���"3�P�p�<$a바���2�&t�w���B�p�:�R��x��=�pE$�%]d�  �+���圓��ێU�:�H��;A��MT���1�̊��Z�
�M�ɨ�mm��֒#�"���f��.[b�嫁�7�V g9�hг0�e�/�����녣�hV��N������9rY���^��t�^�uz� ����k��<M/i1��6��);��Ĭ�ֶ޳�oGX0\r�u�W'���)�w�5�U�U���;wi�48���yp���F�ʻ�ļ[+�R%��h�kD�]������0<'�k����1�_;���9u��F��|�qq������f��MJ[g� `�89X��L�"�d�0��dU�Z�]��`�-���Phc�S�s��5�p��:̕���ϣ#�1X8�1=���:������ޗ��dt\&b�Z�7Ы/B�d�	9�="c�=�z�BQ�V�����yx`#_"�	ԩ��jK/O�c-�B�m��lT 4[m��ݔg�^�ɦ�dN�@�9�je��;u��Ƌ	y��n��{��p��)��Ǆ��sV��z�f̠�P5�$:'}����F�}^�o�mf���ⱻU�3��?`��z1�)Xզ�������p�@ ��5�349w�n>�����B�f%�9K�;�Ӱdy�P�;]Vb�:e^g}� �*�jl�V`���G�aέ<��z♿_0���U���n#�lKu#�#�siF뷴�<�T�0v��j��1R��[7D�ZL�J��͆i�P��;6>�B4�% �{童>կj�7ݶ07J�Z��V��N뵶i�Hr�F��Y%��Z᝝ U]|{�Ã9=R��։�O<bTC�3F�\Ŕr��mq�|cj4BT�9|���j���֍Un'�k�����iJ��]��!�'B-�ӯWZ��a���	�q����/&8[8.d�h�
pw;�6�m�h�m�t��T*�+]�Y��_;W ���э�d���+%�����-S7f#e�[X��.:|�[��/!	;(r\:����76��d�=a�N�כ��-�ov �
���vkъ2��D��b\� U�����#*,ַx�\�11�3Aݥw��o@�fJ�$�ܜy���͠)v�Gy�Ԯ6����5��͊Aok2g �N��Jl�㓛i�f�Xl�P�#��y�e�(����h�ֱ�E�:-l��70��9�
����^�su�����ޛhp܍��%�f��9	��ȇV2�z�+��S�$�m)K6[��t�0�B�1ƑCL��ifC�f�rν��Z7\c`�YC쑅͝���l�IG{���^�Ae�ĎL�[���^'�Vcf�л���x�w��U���J�VK[u�^�Q��m�v1Α�9|y�Ķ�G�r������+9DJ�4�N;�}�u��E|�q�b���bX�:8p-n��*(�s+i�(U���d�N����*9)�)H���*M&��f�ʶ�Ѻ:�B�6����^5����W�`��-�Ŷ��ne=<�:������ЏvV66�*��;.x����ո%s����`��p��.Ui�[9ծ�s��3r9Df%�/ޏ�m����M?j����N��2ð�5��=����{�Y���'��PgW�-�Ǖ_�;#�Bz��s�� ����n]Ks*�� �:A�L�6l{�ۡ��9IM���L�2������0��ԹMyF�N+Uf F�3IY%�k��eA���ا5R��kx�/ف�K�C��|ycWnsu:����S�N����ev�
?`!Z%��nާ�a�]Z�W ���xf��Ӑ������R�T#2�.�Z�m�.�thm:<p���t�$I�t
�d,��L\����r��.6zS8sT)��c;�U[��̔C{L��ǜ-f<�zA4��*]�.e�����b��T�N�3�ƥ�s��B]�B�Wm�@��Dv��k*�ɧ�]Cp3�:P�3�/&W�m������*uL���N�[�빐�WG�������yÊ�YXE���}|��-nj��;������~��U_�(���SEE%�m�(媉9����$�cEQI5��Ti�MUUUP\Ʀ���+l����"nA�h�N�m�(��mSAA�El��b��UUA1I͈��6�3\��\O-Ur�r�r�T[ h�����yh(�������A�kI��c!Z1����"�B��s8j*f�����"��*nA�m1PD6����"����K�9�55PP�Ʀ��V�	E,���f�P���PPP�5͊��J-�%1:̻jLERDU$�qV�Q�����s4Ҕ�T�#UG+�b�M�9���sb�j1���c���xsj\A����%)�"4j���d�-5P�f������������&!��4�r�5&b�ܝWDsJ3�ގ�ub�v�M^Ǭp�mK��࠮9�sdݣ[ͽ�dwM8]ˑ�����+���V~
� h|*��ܜ�A�z�9�ӧ���uK��%t��������C�?�����_��^c�|��)���04{���8��x�}����=0}XY��߿{�����.��r����4?`����{�	���l�={��{a)�>�s�&����T���r����a4�u��;�a�9��r|��r4DX��	O�} ���Cռ�߅�~�:��j_x(`xE�>�mH�G�{�<�{�=������v�`ӥ��_�� ���=y���0�y��w�WRR_l�]��r{�?I�HR$"�l
�2�H���!�L�z��Wѣ��>��"�H�� ����x�A�%R~<�΃�y����:���9����=��ɤ����ox=��������^G!���	2������ �@裂��Ǐ�_z����rt��C���z�/��H]�pO۸A���e��~ܓ����O��	O�}?y�G�>_��%}?�륢����ߞ�z�-:yG�}�|���������я�"$B�]�"�R~QYKҗ��4��v<��K�<��T��@y�1�nO�tw���;���r������ ײ���}�i�]����_o���������?�MϾ�:�<@����T��*qZmU��N=��9=˼�k�w$�:��r!��9'#�}9����N��}�����üu{���s��i�.�~������|�N�v�}���(}�G���{�ZG��(����͵82��h�J�Y*޿F���G�h���71C�|D?��s��'��T�?���>Gpu����O�ry��p�� �<�y�g�;��{� ��h{�^a�G/��m�i4�;߽���}����;#1j�d\������G�#����<���:����u�}���{�����x�����I��>��yR���<��7��:�u>C����u?�P<"=��>�Q�P��[�77�����~��tD{� ���G�->�G���y�z^��使�����^{���=��J��w�op~����}������_��u%���K�|��A��y���^C�{��>����G>n{Я����y�:��Oo"�M�"J���	��˼h�A�jX�n���E����߳�i�׻�q��/:K4 aSC�Ɉ�^�{�Gr��bc�*=���rmw-�\�w͔$��,.b�ή����e���6��]֯���>������9xot��bpwk&uL�Ύ�a4�I�x묿����|���=\�{���J��8O��d?�:�:<������r�#�9�����!(?O�:�_d�$;<���CB���P x{T��ڧ}yq�~Q���<�C��<�� yO1�|��{��}!�_��~��:��u��/�g��MC����	A�c�1�W��<u������M�ƭt_�:���(9	G��w��^���A���<��4�O��?_��<�Gg1�=^K�9'ÿ��p�7��;�Ώ��]�ny��Ο���|�����y@����;��ħ�Y��|&�~܇���4��/y��>��J}����N^��{6
���=su	y������y���<����~�M��)�.���{�|���ݾXAu����h�_��#������=�������xw�k���{��9 ����N�a4�=������:���9:]��rk�d(J�<�s�.�����?��{ۆ���v���m�����G��"��";تp�������O �}�_�45�{/=� �O�w1���_���N��^�;����;<�QԼ��]��ܽG!��u:4��t?�_߻�w�����tP�r�n��V��c�ǀ��T~���a�w�{�:�`�y��~�9���y��s��$?��A���Ϙ}�����d��i4x����伇�n�8!�����}������X�xwV��~��xF�"=�:���z�â_gOR�d��/���}���'��?���}a4�Þ��w=G!+��8y'��N]A�>�������g�K��|��|�wξ���g;�8�*s�>��>�C�D��i�̼���o�u	O��<��9	w׽���~u���=����7ܚ �����:>BP��y���<{�O����L	��8v�>s���������~���.G��y�%	]{����R�`�����9'#�N��BS�?I�u���9	Ga�=���`�?|�u�{���������]���y�i띞�=9o��߮�yM�P�|����(_�Ԭ;?ys�@,��m��e���r��.�甈=�)����Vܺ��vʩ�pי�����9ak��5�C�D��}\�fP�e�7�5p�4���["�A˺�eX[���{0R_+q�Ճ��T��̈�[���i
O?��;�/�:�|�4�.�!�������J{�A�:��:�T�`���A�O��	��=�Gǘ���;�����~�s��%��"<2 0=pH�%�T����!7�gm��[���#� (g\��� @1�fS���/!�|����^��9���C��.o��O���K���#�^N��G!�̿'���C��?.A���x���t>n�f0���'�������rC���S�O�䜽������KEG��ty�KܿN�맹��^����{�S�̼�����<��%Q�>�����9�b����컿ܪ��>�e�=�v/��2m�����z����]I��uR>�}n�������������:������]��|���Е@u��u�0r|�sy��G�r?O����hJ~��{�{�DH��{F!���t���5W�5_H�!�$�'�e���ױ������䝻�?�� �Ǽu/^�!Og_�|����s�?�'�t{�����䔔�u߿�M�ry&��{�P���"!�M&OEW�/P�&�w���޿z�i��zu��?���v{�A�{���9'ϙ9Rh4?֚��sc��z��4�=�:���y'�����{�2���:>C�	xs�;���#��|G����{�;�]�^~���?�J>���?������<�y��>>�ϕ!C��\�w����|��.�����3��'#�r�{y���Z(�Ǳ�B^d�rz�/!��_\�������/�߮~���V�-}��v�%��@
�D@�oO�_�c��=��?�|���p�K�r�����������(}�X9w/#�d;7S��/��:�ް�%��Q0���� #�x�oS����Nj� ~�׭~`�������v&�c�9y�����s�'#��9��\:��~��}=��:�~��~�����4�������|���G'��m!_A��G�h�b�-�V���9�����:]�ݏ��rRS����9'�j����h}���;|�����	��|�ޟ�{��K��?`�����G�޸U'�4���=��K�?®��V*����USt0���q����X5H�����]��5�hä�4�e�@ۣ��z<�gԂ����ɱ��Z�'qP�Sh[��9]Z��<�y��(�A(�2�u���LT	�!�ѻ,R���+>���].��· sb���3�����M�AMCHҦ8gl]4�'U����N�._�e�����:����'f��u �u�~���:�������:~�~���o2���:�(~�~y�����	���\�/�r}�Il�~I�rN^]��������4��;�]�� Ѿ���!.���'��u/�|6z��)�̟��a�!+����]�����^y������pF�e�y�_'�t>�����K�r�(;�?�����w]w�Ԣ�#���ptH�b��H����������e�{};�4%?%�'�=���:�������;6y�O��N|p���%=�y������rO���O���G~��	y�C]{��߆�|��f�e�A.�4}��D1}�w�z^�g�yϼ��ӥ�mﻐ��/۞���u=ˣ�4�ܒ�����c��?Aٷ*B����wy=>���x�2�s���v˥[��<��	��]Ϋ�9�h�(p-����iS8Ɠ��NV^�ٺ��O9��Y��t�;���+�� ��|��=�v�紘��F�.ɺ]z�+ʚ����M?��BՎ�[?4xq7*��2�XpZr�ʴ��MFl]+��7�7��l������$�}�<:�N�k��po�%-�z��`z��a^k6{�O.��/V��0k��[�3MN�3����X�5��KD�b<����]^��^)�tȵ�î\�l��gR���\�}���a'�wŕ��H��rn�09�)�ԚP�/;�@7P�J�e���ʣo����^vmC��V��3l��o�!ڝǑ{�CJ�-�K�8l@Q{�ȣnX�������y��wTcu'�o�K+s��h8~6�vS������apGl%o�q.F��hμ�=�h������/�@q��G2;�����&��ɫ��N�v�*>�t;�au]^QXj��d�����E	�֭�h�^p:-�{C��J�b&��ni�NWM�p���P�qъ�ȃ�׫�jg���ϔ�Ӎ������p�l�郔�����ݛU�-�8X`�fρQz�&$�Uޕ�$v9�ط������O�ɻK~|����=�!aP�����+L�B�AֶM�#!��;�gP1p��VZ�B_PF9�x�rh�T?j�d��"㉟��E��˫��t���=�V���P�{��(1���V���Q��/H��!�!��]W��D�5`.o�u�r_:w�:��l�b�BR,�D������K�I�i��y>���r�J<ڈ��Cl\�P�����`7�C�[k"�7o�9(x
�*�0���4���H�m��9�$ȱ�y�4�r�n��:u�tT�+��*�κt�,"!��ڄ.���H���Ef.��EC��t��c9�iIֻܻ~}S�\CzljA$ze̷r㍋�jB/%�/n^�4R��T�ڙ��=�kfnHc�R|�Q����=>]*��FN���/���{�o,�73lI��_Bc������WvU��x�������*�����{�7�F�*��-��;y�]7,�	:����f��(px��+� n�tj���O�^� Vy�1D���OEۥ����YGz��BƵ1�q���Ԩ���̂:��_O��ä�x�/���ۧR-�N������@
�muL$K,G��jpF��+E���i�>'E�K���֓��ż��1in�dCrgt�6��hbLGW�e�#Z�^�:�^�yZ�t^�G#+$j�\e�fu��@��C�pY}'a?BY��x��^�63a�୙*�"����񞹹�/������\;�-�H�����y7 ��^��t�b���k�Q
v:q���s�v� s��.���j����؛Xj�i�a��O��'k�(@��ʻL����}ס�xX�R��*�xx5����Ffa�a6q�C`�n\���E��xf�"A�&#Y�����b�C���'��{VfA��F�]��sѤ�x�����)��#H�U�����Nݷ�97KB.�8����͉����q�Y�`5�pkͺ؊�sp�D�O�Q�Z3D�YF�M���,	:�Xek�i-)��F�ʳ	H�MbbjP^ʵ��ܙ[��'����X�mg|��R��R-HB��+W�7Fʜ@��k.=��l=櫾zV�#U-SO'*�Uә�xw2�|���j�yG��*�a_��2�b����G�Zn�u�����pi1y	m�7�Ɔ6�{������w�ͺ֪�a�/s�7�ƍ��@FM��rO�����޴����"_s��6�Ƿ39�˪��h�Y��ݶ��R��Q>��u�_c���(���!�+�z�?u���'.ߚpW�F��v�CB�ԭ�ȓ	'ܲ ��1Ԩ2-2r}��9����ٯm.��v��dG����;��(R�׎���S��2�V�m	�R�
������h�����ӒZ�#R.�9$�*!*C�j�kٕ��]������@滬�t�>��w����:ja]�w�!\S�:hJZ��c
���S̲r(Ǒ�m_���N��1�WMI
��ö�L�idX'�KF��t��x���� 1�.U�\�Cx�E���3R�y���-�<ۖa�`����X�p�$��qPE`2P1��T<��q㎼�n8ȉ��˫�������m�Ŋ��k�[�|��t�M�Y(�5k��5L�L��b���J���{[Z�d�r�T���a�~/�w��ht�����Y��L�'m'�(��C:r�}z֜�|�����g�:eۂӶ�g*�B_we7�u<�q̀�&$@�����K�ө^`u�q��?W�,��	���:�vh�C�$������W�B���Q� :�յ~��kFw	���Q
�P˩u�|^�;4$�H-˳z�21�1�]�Q|�W�z��9DFj�艛����q)Z��;�5Lb�r@p2��sQ�ny�E3�hH8�6F�_�)��+�V��i�
��"�V�P�w<ì���| k:# hZVj��.�"��'��B�[rdkn�۵g�Q{k9��iPŤx�L��D�'^�������GG׉m��-Qb��������7�n�=2��-pZ�ޞ���;^��u[dHG!�"Oi���|=>�臄�a�͢�s��W:G�����8�w�0*!{����90P�0��:]�0�3^�H��>����wc3);~�ڄ!�^��ԕ��Tӈ�����-L��A�a�3n�}Yd��>�^a摫Ӓsic����B��wxq9�~4��o.Ƈ��:��:	���k�Wx{N�`w��Y��ڗ��n�f�+��y�W��'�ɡƞ�c��s�Nv�.l�Ǖ+*�;wDO�[vF&�bڼ���R�� ��a�/�y�Ժ��V����J�+�#3-#��H�vz�[~�J�}tb귲�r��J;�lm˶/gRi9��	NWfoNF�l����(��p�^�`H�1
�ў�4�=I���f{fk�7|:
?�$\���-\:�r}(�2oY�O��M���<�_�;�ak'���؊��'��ݰ����2�5�eWT+�x:q;3湁�b����`�S��Us%��d�}��n%f��Kez�}�7�V���T�,�����0X�Z�n��x0@�;ټ��.��ݛ�:ɋg�Y�^Nvm���Olhd�����;�/�W���w閂9���Raip,d�y��Q�_��`�:�H�G'��o�9["I� ��|k��'��9�/�.�½�9�����5��&�+z}�RYz|0Cojd�=ͪ.wWM�힛�=Oa��8X�b:�؄!��"�^���fç>RcG�^t����T'!�c1P��Ql��o�9��m�~���b�Ph�{D�P�����z���� v9�ط/��ъ�`!$m��mlV�cvwI����Re�H�#���		k��RFC��w3�(@�%���$ՠba�s���Nx�A�q���ȊN݅4���q�_(�9�i5�ہҩ�bɘ&�}*`Q�g���x��j��[�ol��y��֩�t������AV$uYv�_*�=U�%u-]�9�!�r Qy��5{
K];U 붭b��I��-&/���^5R����]�5h�W�� H^�#���F�*�Lφ#Uٗ���čG�5T2i�Z�3L��@9.uNK��#�k�}�wByᰕ#��b}�گN��zĝ�~?w���-�(����u6.j�I0���:��cN'����Ȩr����\MZ�F�]��괋ƼɦX�w��v���ծ��>��3�c>�{eV9���g<&�f.���ťO}�E�;��BQ���U�d#^���c�t���84��~�P7f�U5|J����cq%�ZVo%�/,��c/9l���\:��A�r�����;�g֥(��9�P�3��}>T�%��r�Ȕa���8�I��lD!M���CdÁ]�[��5��U��D�,�������[�D7͹A(YRw�ַ��1�s8hK@w%���ɑ�s/s���6�/H��5��2�D�d�����iF��ӽԠ�-]���j�
'��	���F�l?1�ʾ�T�������/�U�-HG[���+�T#�����a��%��pt���G����0�<�>�h��~���c�{�flଘ��фV���՜��"��;Bh��Tu�Ǝ��J��4o�簚3㪚3�"��oN�gC����#��<!}2�����S����w@^��B[;�
N���I;٭ڽX
^������@�R��`�3[�S�F�V��K�W	��F�h>����f�io��ۇ�U�&��s��;����fp+�����Y� �n�݌%e,�lu�Z���ͬ��/��Q�6 �+%[aV�W����@L�)\�X9Ri��Q�̩Ruo&��T�Iõ��2�7�m!����;��uט+�J<w69�+�a���,�;m�������+q����O�R��M�g[���E٠~��Ҿ8�B��[��*���哈�ykFv��3�1M�N�0G �2�v�ix�)���O�/ۮ��<.�#�����L��:cGX���WK:���0L�a^WK#�A�-βWD��
�A��� �u�͊��!�
ûe�ޗ���'7Πp�n�'d�Yvu.F�JVE��T��~�M(�e�&�V�#�Dp���-::S_9S�ڻg���>�� �f���Zxf����yE^�Jr}IoI�}J͚ܾ��6��c9EJ+q��� �D�(���]:�ƶ�B�R,q���ۋ%m7e���b?-H�i�p�/���h�κ��e����$l���N��C/n�5eMy���K�����KhlۃN��x�QY0KO���3x���8�'h��Z�!������T&X��e��Y6��&L_!s.Rĩ��Y�V�{4�9i�Ө�w<3JLk^e9AZZ��b�1t/�2��z'�X��r^�$�`1�*k{��N���Y��v�
�^zgCx؊u��Iq�Ɂ˷��SE��F��Trl��l�:MNCV�f\\���u����f��{A�d�p��=��a0$hJocJ�Ӧ�-��8�M���U����]���mȀ�=�ur�a�{6����M�\e���ݺP�9��Jm��ﯮ����sb�L��(�\$z\��Ue�zU�%V6��Z\%��֫ �L9��doఱy�e�7""j�)g~������fG[_h�0&��O8��ary�j=#�-��Ru��_e
�����6Ik`�Vn��D� T覫͜c/��egBPR75`#�Y�F��SB�����աC��8�(+f3)��Ů�\}bn��X���Lj.�1vFH(�X �=:�L*�."2#�)��v'��[��R��+3*��Z�s�XN}�_1Y`Y2��lZFj1g#�7kwQ�k����͠F�gk ڝ*�s��,:�4�S�wx/m)��j�4���;��޻7gM��Z��겫�U1���`	�S"���@"�u6�;,�����w�(٘�!�	�i�طs-η�^T۝��u���+y]����nvB|v1���S��w   |" ��Դ�I�5KM-1?���"�Ӧ&�m3P�I:�TQ��rt��H��ܢ�m�ALE4�j��� �mS$Q�N��UUN�A\�**(������6t��)������"��b��g$E5�$ID��!�PD��REHSE:�4%D���J+I����i��"�����()�fhJ��QEF�ACl��q4ѭ4r��4�:ѣ4T�F΂��*�"��F�"��IESIEUh�ѡ(Һnn�EPr]��D�@�M S�*�Ť��%UKA�
4j� 4j��T&����:��))JJjZ��M�
�`�
����MKȧl:)"h� I�!�ԇ՛�:6�%꬛h:uhh��r!�mN2kw��:A�pb�Ux����΂�lAյ{ �+{��67�?�%Q�;�(Wl��O�5'zVЦV���W'�?JWI���P;���#����uP�-鐼�y��Y����-ߛ[�����>ʖ�K��E��ǆj��&#Y�ś�kO-��2��;�>q�|�j�D�9t6(�^�mla=����S�S�1�(�d�7�q�C�gx3�r{��A�.�н�{6���,4�f�k&��ݏa� %ɪ�b�8z}���^T�d�`�,E�X|=ᒙ��z��rh6��qM+d��qE��5V�������z��4x�j��]��W�������sZP��Q��bl�����=ѳ���cY�e�B|�YDΞ'_�����4�v��x��lp�Y�}÷,I=�$��sc��KV�b�"ٍJCi�>րX�T�9"-�s�5vvO@yq&麨��+�s�_:��M�Cfˊ̸|�T\Lr�M�1>�r�iU����(>�p<Fa��@��jivIr���k��eu8�Ϛ�!���l~���w0E���o���X�LYŷߝ
l��@ը��74K��5Zl�5$x����U������c:���:�]�*o5���^�Lrt|���h>qOz�3�[M>銜 ��O��n5�����X�oT	X!���4�#H`�]�L���sn�r��/��� ���[�Ͱ�$~�<�	��5�Kx�8H+_!�0�����R���|צs�i0z�������)\ո}C����h�.���}���̯3�L��� "2�ʳ�r1WTX橀��;����!]���װ�p�\+u��:a�^�s{P�[�DbgV�3��Ř��x�9ȱ���l�s����^�=�+�DX�?w����D�e�
�}��&���Xz��&���N�~��uh�%jyD<n�~;
�Z�\�j�J>za(�rsUȣwǧ���%u[>�UA��VI�fƵ�x�u�6Te��#s~����?j%�ƽ��TN�MwU��P)��٨zlO>���wMH8�>�N}�㖎�O�������H�:��>�D8�!_L���u�S:"ƅ�f�����,7��d��j���.���^�hX�긨�4�2:Q��	k١�Ja�X�a_ЧG�Ki�	9��䄻���}�v�e���z�3��:
����$;��"��h̞����w�1zKt�A��ׯ�Rl�8P�Y[>�G\K#
��<Pp��Ցm2��P��S��1�./�oo�N͌��΄X#0tN�,�٢vq]��pp^K�ܪ88�wHMb[�����Cں���B0�u~�9�F�7aB|�ffW� ���e��$�����} >�d����F����yUM<N0P�0��?�v����~����3|��X#��:�?nz����������আYv~����}�<e]`��Y=��X�z�~ ��VLh��o~oVj�nfWk�U��Ah�2��i9콼�ڴ`I�i�[��@�g��B-yϕOE짤��������<��)���k��.��y��L���=#o+H�!F��Щ}��GP�r}(�2n���D���4��ViJg���F�|Z��[���ۊq�(Ӗ�p��*�}�<.�N�k��5�E.��S�N��OK7=V�ߢ�}��������=6��*�
�N
�G�i��+3����3�f���Kc�U�ɉ����Ӂ���8�9^�vԫg� ��	���r=S0��Ez��뉿0��3�|g��T:�k���d�!��f.Z�7ʲ�/d�v״�-����s�	6�q
3�4K>��F�$N�O����<!ȵ�#_���;��c¬���li�e��im���� �J-��N��1L�e����$xz�ȋ�Cdӧ�ή�4�gS#*V��5�wO,�R�@��̷/��Jx�����98Q�哻N�_>B�|���`#�!&̾�z����W,xf����ѦV#�7�A����直���߮m���7��l.  `d��}��)s.Z�a�;��qJ��S*110ܟn����f8����]C�T�k`��F@r,$T�g�
��֍�����]B�������h����m��&�:M	2ϧ��+�`Gl��BZ�dԑ���(V�31�HƷF�;�S̠b�}���/�9�EE�>m�DN����v��a��{c%=�rX{՝�,I�98��7;���A���������q�Us|��|�f��/gV�J��N���Ye�/ٸ����I���M{y�z���嬔k���k�!����"��qqM���w^�9!��5Xy:6�S��6��������;��w};��J��>�Y-��)\	S��c�rk�}^=eY����B*�U�����`Sc���͵~�e��m\��~�{v���G��S����]�E���8C�S�vXHW��TZ��Z��p����j0����7�Ծ��_U��zнjct�ǳ��QZY7x
fA}>I�Uaг�(�ŕ�M,���]��S�>,S�6���,�:Z�v���(3�H��^�#ޮ�`���T��_jM��s���n-�]�.��_h&�)�y�V.�Qfn�au���_`U�Y0� �l���%��s'�:�}�}_?�Ɗtr$w�3�%��m�u�6O�.��P��:��KY�`׮�-B���*%���\L���Y�<x�_}���kb:�e�:�2��לm���C�5"�۝i�nU婪���F��D����A,)��U��F�����|��!R���z�l���Aw�}!S�>�j���tQ�<D���\Z�,i�[�ք�N=W��:񼋗�֜���O�6��>g�!	�$뢸�!�*�2��G�R�w}��Y�&u�v�YK*5���7r��z�����6ds�A߽�3����7�;^Y���x�21��5-o���S�����lkW/N6�0�x����П$yh q�Uk�Z#�_H�s�x>g+'����PXu��|���/w���id͵�ph6�bU �e���:����˚K7\��qu%9�`��tEIX|=b1s#6�얋m��V�w�R"��&9��g��o���)��^��RЍ���8Qbm�7��洡���n�L��k��s�-�E��]���l:L��p2�OQ�Wϥ�/a�4��~�~�o7������U��l�K�z�>�#���@Ɩ�uk������)��e��:�T��7���P禀ϸf��	)���{b�Xvp�r�&M��7�١�iF3��>��W�s����%�j:��bq;(��'pE�`�$ c�����x���\�OY�1z^�X܆qS��a�QQ��$�q�րCJ�6�91hn�,��	���������=R��Lj�+yn�ƼX�ULE��Ǌr���*a�
vx��x��uk޻��T��y<�)'��9s�k�R�Sg2z\w���d>�񱮤�ݞ�;�"��c�O{�4r��^�L?�ώ+����4%.�x�Ā�}!�9=~��6[_{�|��F<�Q�S֯r9�Փwt~*��$?��u例�B^�|��k����K��1�.ռx�
�G�VP�uގ��o0�nz�3]��T��[�������K9�<�Ϳwht�'b��Z�I\�z!և;�ms;r�a��(�"|;nWX�?w�+_	M-�T|w��(t�y-�$h��eP��7x�Z��C�n�������R<dq�OHxJ�s6FC�Wu��-�c�פ�p��,���<\�����f�֡���Lv��^���:�'�tp]k)2q�/2zf�q���"�jub��Hm�21�;C��ڑ�>�sw�k����X��FQФU���{2HoZX�&�J�ʝK�g�G�;�9�&�8vM�p����r�����v��TMh�[@�KP��E 
-�2��������%%�{��]k��×uQI}�\@�=��c���sϨ*)��\�q�m�`l�t���ڛژsi�y�W�S��pF$p����4-4�kF�S>�a<��5J�<�RaO����@$l�A[]S*+ܑ�#�0��#�T�O ��ѩ�P��2��@c���7�d>��QUruuQE�<�LO��7N��)��	�v���h��!*����`-�kg+NtS�t���gh�_$����_���S����#�#�h�+�?W�n�5���������H�yN/�M#^��#�|�q]�)��'�`jd�9R(�.9��fj�6{�?s#��x�3�{O}ܫ�b�	'U���%��b2Ἳ N����[�8�m�'�:�h�j��0��jk#'M�f�+�� ��|��=n�U�2�o�>�u��V��:E����5l�!j�F������7/_ ���=T�h8�f"gz���#�[:�9[���9n�,Un�D�C��`�smQ�"�d�Vf��ر{$#�N��pO-���k�w`�0�$��3]��J�]o\������ �I�A�1�]����A%�+V0��]ȅu3��RI����o��E70�pVv�/��hKl<S1����{��^GY�"JV�o�t��v�?x  �f�����r�LFU��������g�\���<��m�,x��+� �\PW��L��J��.�(�j�x�H�9M��b6�ֆ7ʲ��[u#.�	8^O�bH�z/45��u
��ٱ�1���5�g� 8맔9�I����k2����Ӿ<t�u�Ԁ�Q`�ȅdu	K���b�caB�����Ø�u֓�d���ԋ�g�z���&�8ٛ½ �,�( h�%06t�? ̞�g�����u��Oj|�����q�ػ���r8z��}r��8"x��6��,$�f�#L�ܼz�˝��BSY��jN�� �c�O�����nwI����BL���#�`Gh8H���1�5"��Vxn��n��
�ꆯ���C�]"b�f<-�qӠ���^��ӝ��gH����=�������>͟pgqu{ʼN�ۭ�,��B�@��ύ? ͪV){��fq Ul���;6�
��Q��ei������A�Y2m7@o��lV̿x1kw�c���ns(��5��ZQ ����bݪZ,�̭�un4���^ٸ�C�iP֢�W��!�������V_ڞX�;[Ұ��]!��t�mӗP���$�](E����٪5��9�!��Ij>�*+�0�<�܃��֠�W�}_}�|g�=}ߕ��[��B�(44�k��&;Gǩ8��e����v2C7��~w��;�vV�
��|��r�;����T=���B*�X�^��l���\<y�b���q�\Yѩ�L\l;r���9�"��FMu\0��1 l�Ϻ�!]���G��+ڶ�eM�hiR6)��h�s Y�/\�hk*3��g�.jTV�M�:̡h�f�M6��9m�m��r�d�I?^�d\D�l�#�f�mV�3�e�
�M|�Q�l���p�&�*�]:�n�b8K���Y5�S/s���6�Wsm�'���u�1��{��>�Wba��H��$�d�s	duJ^�Q�0M;������g*v��T����r7F�K}�;�: }���p�G��x�8�+�T�pik�)�~\��Y[y��K
��A��� ���w��H�3��P{c��>�D��\p��
� �+���(yׂ�8�Y�1ej�9:19�Т�i�� �����;^hl29Ӡ��G�j(p��%�C�c/
r�x��[��{m��"�؟�[�wc��zZL����E�f�j^]���YQ[�Ĭ�#�ٔ7��v���u�CX�c��񬚷�įoN׏��DJ�S�ַy��,�Q8c;(�g�v�tv�yhT+N�f�gZ���v��=Ljn�&#,�}}�#��	i�����Ә��i4�
�<���{r�7�v���h�� a��*`��*�O�M|�E}_$�#�3�>s��nw�;/];��z�x#y��vt�=�{Ux�c���7~)��ǒ�r[1����th�f�V��7�+�g����S�����R�t#f�|�
$C��/OY�iCt�E_M�1g[���D�!�o][ [�B��Eƞ'g�k�"�$.����21��p���z���Ȫ��\=�T�s1�h�N�9J�L����B�?`~�Z�;%<�r����&���,�vz.;�fˊޙp+��a�r��v�ЫL1���A��:�����e��@M��BR���=���q~�	���!���~�^�t��VW���>��k��a1� �NQ���Л��R��x� ek��\�%�H�:+b�,fuj��/��j���&+���*���o#f�\-�K�iy���=�	�;�c�5�M��D�.��B�^V��a�֬����KW�Z�� �]_^�E�_>���f���V*ܵ�ֳU����r:#�c�.ve-`�sD�G|�A�h(n��d�u�]}�v��0�\��8�q���TѐA��t(��:ʼ9��Ɓv \v�7+V������d5�I=����l�Qn��� �g�Ok�n0���kF�Cx���BtEh��ej���+��4WV<�R�ꀹ������բn�
�mM�a�W1�ñ�(�,X��KN��`��/�.���H=�c�{��{���xE��1I�z���PwMN���������ѭ齹����m��Z�����G��,��3��͊�5�U�N�Օ����B��R�s�3^ݕ�_3e}���]
�B�v���sVmq�D�)��b�ֆ�6�k�Ƭ���ŖN
E5��P-�<��+���A�n�f���A��{>��S�a)��U�)��vjL�BwD������	/Sy�;���V$�(%i��<n�74�qb���3O�+k#��9�j�/���>�H8��"	�6>�Գ`�]�P �5z'[���C��9��+��%=���c��q��óy�æ=��C�u�3��f�/r%1�xJ�v��H��>�ڼ��/+3Gü�W$�/U�n���jĻ�̻c�>������791%��]�Q7�kmG��
��m�[�.ݓ4΂_1���dۡ�
spn�+�������	B�񗣸���A@,�V�\ ��%���9�3_��DLT��aU��7��q��E�9f�=ݺ`�J��6N;0��9Kz`�0�\��{��Y�Q��kޛ�`���y���7q�W�`�y7�����M"��O7�GLuwm���h��b��!���մ��1,�C5��7lfM?N'S��9���3�ea�ږ�S'��b�E��8����ȯ�A�v1V��(�>P=�К�u'T\MQ���q xQ����杲�n�c�e�١��9�8���Y�T=;JC5�4v��'��]Ѩ�`�[��a8�\��eڂ8�����P���7	׮��P���kE�aG_*���U�0>�n��B�P���x&ݽlc�*�2&&ؚN@uӣח���"�WF�u�3��X�� tP�Xgk_Z �1�[X\�,��pQǘ���O^���tHλE������m��]�p��W!F��̾�w��I.�W�"]����s���-n��1Z�YgU�ġ����s:�f�y����g�T=�������Z�\"f%�d���F^驦��M����E��y��������L%+�T*U�b�M�#.�rfA2���+z�:55n��G����np�M�1Pf9��s���.�S�Ҧ6�����b7�-�=JPҾq�����h%V��pr��vr��=����>�8.k����#��AKy�hg-��`�6n~/��~���UUIG'Vؔ����"����U.�":m`����"-f#Zj�JJ"
��������w 姘�QB�ڊj�lLւ�El�Ć�T��4DD�&�E0��9�������(�
h��l�Ri��(f�j���*�4�IM;d��`�0S����IUM�AI[e��X�ւ6��)��T�!M:MTEP��KDA�����tDl��� �rNIDEU:��$�	M���cEDR�bt��,Z��'#M$MUPhIAs 6���%.'IMDFƪ��A������[r���#gM�AM�DKHRQ�4&�U�*�-=�q�Χ��Ve�M�����B'���-N�n�X�� �U���x(�C&/O�2��uvs�#�>�x�t��v�sp����z[=~��=���1a�p�b7AB�(g�2��zeK����CBj{��01�ݙl��oW�$[zy���˝����$v�iX�o��"��M���	��A�߁-I+L��7v!z7x�[����^xk��c��H��I=Q�/�ষ�Nt�ش��_S��,�hM!r�N>��.γ�v�m�l��n��_��^�Y���.�fU��$ ܑ�\1���jc����
�L��q�m�`m]
1�:W+J|�sg������m�<��<�"�m�Z@r�������ˮbg��a�����E������6^$.悼�Tʊ��Ș0�4��*|2��)�Tt�� <6��<kk	uʏK}N:,�QdDS'�g��r�)��	ꅶD�#���x��Wl��4)�'�C�Y���}ۗ���?$���r���"���"t�r����q4��V;S�y�k�{[
�S�R�5ܸ�Ϧ��qѾm8�.�m��>���q�Ls=[^(�Ǥ��a��L��Z��o��j������=��*tرn��SpӦ7�����f_!mkd.�әx�����v�gtx�8�c�U�down��,f�]M|2gU��%	琴{��&�I���=9^����VeŌ\~ {���q˱o{א ��,~��ka��=���LV+�wzL7�w�FU�<+��=���kRD,o<�O�w��Ř}�]K�L��O���'�u�[�=i��.� /���=Hx��e�<��OC�ڼ/�@au���f�z��릭����dfUwֱ��
yc3���%����\:�LU�\NX_r�=h	b�w�#�OE�)�[T���ƪ�l����ۈ�xF�*n�PZ�ߠ���\���瓱�Ii�E���	�R�.�wǹ�YG2���h���7^���\@�rE[\�ܧ.�Nvm��{�R����|����W��'C��I�b��S�J!�a� �䪡h�O�az�\&b�Z�5k�ư��d�R�`��`�犗��W`׎N4�=��SK��b����C	־���,�7V駙���S�ک�����"�<ܸb�L�.�B��%05h,w/���>~_)��v`�����M�I0?�1�G>jNg���P�t/h�����k����j��|ך~��t-U���cTH����������m/��
8�Gԍ�ˋ/�օ<�ޖP���C8�w�S�h+���yY������@5	aǙ%v�\������4��@wlʑ⽗X]-��Lt��j�2�n�oLê�+�����{���$��^�P>���ؾ���f��nwI���Zg̿�P�zE��XO��*k�k(����z�Zy~,uM@W�H�!u���}]sĊd\q2ۜ����U�"	�{�T�R�U�м��]�#�6\�{NNl���;���oHd���|� ЄX��+����C,GVu|�z�*iz}���y7BW3�hs1�s�|���u�B�vn�83���)�h��{�����ª�1d��fg/L���U�oo�3sՈi��X$��h�Y� ��F��;��T���}��i�9\�(״�*�"#W���\t���H���|��=��>� �x�76�Zڸ�jb�� ܽ�`g9�"��^z����n X�6~�U�+��3�}Ny������<��b:*;u���8�qL���B����x�}75*+K&�/VV�9�{��6���#��ʐ��$��� �Ԭ���P�!��������x3�L�ze��y̮�C5�8O�ϒ�2VHu.g�N��$�tC,��2���ᒾ�wN滪i�!fc$n�ۚ����ci_i
�v�8�+�&��]I엓dňfbͥ��S��goT�&�s�tC�g]�F�yفM]�����ҵP�lWt]��h���+�!k�ڢJ���	����6j6���5����Û}ο � ��5�f`���·DުG"��D��;0OT@a>d!�e]��l�V<i��Uc!�x�����F���x�<��f���x������<+�%�D���r{Y�˫Zu�뻞���4�	�siǩ�9��B���9N3�0:$�+�_�H�\|�{����k��U�g0���Ѥ��#1�q����xQ	�V��+��P�3~ف�]��_^!�鈟l�X��lH�{Bk�]��W/N`nz4�x���'�H�|R�E��4ۺ����:��B�#5�A�=����On�gs��ɸ�d����q���b(�շy��y̒��~�@�Ds;B=���1s4#6�5�}�w�d��ʔ���ۢOR�'�39#�q1>�@ᒵϣiƚ��u{�I�n98������=�e��83͌u��97���$C���wىوA�݄<Յ��;p����o��w�1\�m����F-�\V���u �b����v���o��i�f>꭭�n��ȓz�����HL�eI���𝮶ew˘|է��h�㕷O1.K1' �����\vۋ�k�/YםsV(õf�ƌ��3@���x����	�c��B�NZ�oVك�~�����.�2���'���_9��ו��o'�|�3�Nx�y��Rf1��9iu2lOLV�1Q	�9��]�
�d'qs{�=:�/�jŮ5��Aa�tB�)6��v~S�5 k�� �(w�+�#�F�p�<��=����6�1��gN]|�������$)�%|8�7=�~��p?��T����Ipg��/k�}b8�Y�3���M���4q��� �Z�������k�]J�V\�]�Ű����y�}�h���)ȍ�a�H�P��.�+_TM�˕��P���n�����yM���j�(��V<�ߖ����@,�0/Y�vCP�d���k-�Y>w��ֹn���H�c�w3\�w$(���p~��w$s�y���ݡ���ʭ��
��d���ח6��Za�7)�8%�!�·�T�X*y�)ǟ	�����۹$���m۫+K8�	��r8�46՛�s3)��6�_�Vu�]�D#&��l%�A[%ƽ��#�
�����y�TE�
΁t�s��q�[��>/(\;Ϗ@�Ĺ�
Y�],�V�{L�LwZ�p�w��	���q��}}�uj��1W�ս�'+�?{���8_-�p��*��>z��D6�,��@�bߙ�;���A^���!��#T��㋑�_W�{�6�3a�f�����3�aӱ�9�d~��`�u%�5�jC����_=G;�à!����+��u��w��r:��׷'z����As�"�Fk�C�I�\�����ۼ�
uZp�t�5�
ќ�b\4"���<n�ܝ硹�f����_l���u�li��iʡʩ���rq�vd���58�TSً��N�vE�g9�\�m�֑i¥�YmMA�}�c�j3m�OM��ry���T�B:��*��� �B{\:�/�s���s_/����Nzr�}:��ƽ:
ɹs��ǰ�B���bFs��
�蓯��M������^��\n��v�*����,^�b]Xy�.��V��ۉ��o,	|��׼f�����c�+���smm���8f+4�49�����Ur����Y�����z�����������
A[)�����V�v����`�d.�W4̊ѽ����;8+:2��48�ݺ�d�b�y�.LU���|�eX
R�#*�u�*���}��=��y�Wm�t|}�L���2�Q�X��o^�����(��N�7zۚ��6��}��?,$�?������:���p���=����e�(��y��M�p(%�hQ�tCKs��M��.]�!���|��U�R��s���pb��5�9�
:�٫�2#�"�5������\KW9S7�OL��_H�{���o[{�m�dK�i�~[�jw`�lNG��n��.u�X֪<���4��^�3�%���l��J��&VC�W^)���#(�(�cR�-H����o{Y��æXǲ�q
�u���Y��ol�bga9Ó�;�H�Z��ڟ^�Nk�ϑ�ދ5�^���b1$u��do���9�rb��W���~[w!u�wג:��.��wjriq��Q����P�a��u޶���Y��;]�t�w��L.��O����l��vnL��^]ee�<�]�� �q��E<\%i>�I��\�ז{�Y�r$����u���.sm[<���V�����P���-����Z��\MV��9ֆM��v'�u�n�FT���0������ygi�t��\��n�9sox���5ׯ�c�m����]��ƍӗ<<�?Xt�sǳ_�m�нஞ��Eo_o����i5;v1�]���WE/T�cu7>!��oש
��6=/�m���M5N�,�y�^�R�<�.}.6�Bl��|p}^��H��N�o-i�2ҽ��9n�󏳘K}�.L��}�(NH�����/Np���ir�&�~���l��,��U���y�r�(�}�`t��N�vD?[�Po�����C�vp߫%�+^	_}�m<�S�m����0)�t�l�$מ����RÅ'놚���[P����qB�x}�Zr��:^���.�B����}��O�{��m�_���l��NmL�B:ki�i\�J�jv��c�`C׵���ǀN{�I�=K��d�}�:����ǫ�u�GF�ɰSs7etyn��*6�!9{ ]�ĒmS�E�,�w��r�Q[B�=���p/1N�X��!�r �RO��M��Aac��૕���Zՠ��Y�OI�9Wٝۻw��FmV�M����O,�ۿ����җ�عS�lwm�t���r����>/	�uq��6)p˗���s6�bД�UrS�����|¶}� 6x���"2��h�ҫ���s���mE��N�����f3�윈i1P��w�&�&5��ɀ��W羣�!���˞9�fZ�ww�]��Mst6�k61х�q�G)��*�r�M:�T�X������*����j���]��ߏ��5�=�A�x�.?ld��,������.�-x�EMf�����S篛9mV���rE�+�Z���?{�Q���티���*�m\��D��z���k*5����]ŧQϥ�������Ox�2��3�֖�~��s�py��y,r�Oۻ�-H7f���H�q�c�C����s�݀[D9��X��`Sq$�JU�}�'�͍�>�m��@7�h'�k���D�Z�X��ھ
��~� ���)�+yvN,>>�@�*]\��Lj�i��
�bWˁ������s��y��e�9K-���/y��H�e��5-��e^X-K� v�#�`��7�K5��S^��h���"*�]�v�~���{��ۭ�x�O����,q��V���o^x�����ړ��W>�Gc3;)R�p�߯��y��w]N�9H�bO��(x]�;JDl�xխt�c
cI��|oo����P��֯l��Az�c�T�q�V6���m��Wx��^�ٲ�_�c��5�vECɑ��TC	fV��f�R�k
]L�x��o7�g%9f}�9{Gj����8��
�X<#�_��/�z��N��'{�����mķay�f@�Έ�B�7����E\��Փ��(�p��;��/�s�y��p�b���C7 ��f�ȜYO��f��Z8#Z'3���?�ݣh��Cn1�V��Y�kh�z����s|�l����'w*�ξ�[���'t�{�/a���������W{�X�f�j+��e7r6{#+3�{ֹ:Uf��l+�G�7ov,$��J�kEh{z�T��"��}Sx�m�hi�m�6������X���k
�����9���c���ٚ,=VA��V�,���ǒ���-�u��W<��u��+�:WhYɨ�Y���5�Q|�W�7qGr���:4��	CTm��G-靑�ȷ{�*4P�Aޗ�7d 1Z��	��Ue[m텕�[��uD�>�m!��uCl;귇�87B���٦�/](D��H�ɷ;2�yL韑���-Vr��4O.�[����JF�[(_�U+/{V=��J*�%�a�9�!/�=h��9KAsMA�+"�
/�kۤ��X�ɝ���/��mD6��{jV���;�p���b@u���2�&fҔ��@k'V�W�K�;v2��x���z�B>�޼�rs��1��<�;,!�\�r�@�T���p�-˙GVl�ͼG����FX���i�]a�i�a���l �fXS۪ۨsQHQ�JV��W���Iw��<�3eY�+a��T�䏲k؂���������@%�1׼V@m�,Z�^թ���r�y�]<�6ٷ����Onξw�cc��ғRI\U��p��n�����i`��1���4��Sjq��\�y��9��]B��N�k��-)0���ql���<�
���sp(�;���0������.YH8�8�g0�%��}z������ ��cѪ)�t���+`���
l��8h�
%�yǤ)�Ĥ�WDI��A2Ӌ��݁�ٹXs(�wJj�GH!�\vM��b,���	oF<�ΈԴ�$V���mV�d�=BH`lr�����}b��Ԅ�}�w�!�DF�g�R��1��4ii�������JnV&���G�$D�y�Xm�S���;-�=R��b��s(x)�� ���튥f*�wck��,LR��nR�
���\E�EB�n���¤!0"b�"�ʼ�W���l�L��Jr�,w���̇_R����kֶ�K��\�*'3���V.���$������*c[�x^f6A��%G�Jg�Y�s{Q(� .�c���p�}
��Iٸ���I��Z�n6/�m^��)�h=���� �'L��x��Am�Ҷ�Z�\�n��S�*��[�����5H��7�s2��
�����GΔ{�7i��q:�{�SO|pt��,O�2*]b:�����C�f%vHE�Ƨn�k	��}�HM�d�MY�<�=�bu�®��e��,��d�+Qd^����N���01�h�т��p��̌�[(��hIDp��}�cO�`f��&�H����q'�reQ���k�s}�N;���K�Y}�R�R��ݼ����W�I�u��(�v����'��3:������m��������uR�(��]�Z����>�9*'��.�9u��b����^d�w����V���
����%ri3��hk;$KHP����Er�KACCI��EƢ�u��� i)��i�%cm[DRO,�'I�-���hJi(b��i4kr�MR+$F��)�N�HQ��kKI��i�
n\��9�cE��J"4��)��i"(��T:

�14(���2DU��LTPh4�s��bh4�J���A���%RS2iu��\�hb�`�PV�:�1��h�
JH"��gBr�:��k�-UQ\��SM��+F�h�(bZ���5A�SR�Nڊj��@� �s�֨h�����&���#l���ĺ���NH�(�h��y�~���^� ��7^��yw�o[��u	� ����/wI[Kgwf�ȭ���Sa��>�7q�!֬G�Cvf:��������6%�[�;O(>c_��m���Lϯ��A֢� e��}#.��� ��W�<��i��e�5��J��ٮ�·����P����k�̨���>��ar�E��1;�u�q`'�!����y��}YJC�׈��J�\��2����I���;�a}1m�������Oso���E�ភ�9=�
�^�3��[�T��[k��F7������5.�eT�g���leӉ�z��*
~XO�|��2��{O^��K�6y}�z4��X��͛�w�����޽�T��c7�tEzG�1p���^��i���^T/�BJ���oG���[r�

w�����4@�=b���\����v�ڈX�������{��.FƑ��U��~��U͸���v��ǹώ��j�-7��q�g�W���;�B��i�J>0:����. ��%51]�.]t=�W���ggV��EU�ЗWۍa��ݗ�1$d��(_*���w�xfۢ��ê���&�ιu���d�$�TԊ�sÝq��ھ#8�xd���n� �`�����+�n�Z�MH4�:�W�UW�aQ�w��mNi��3�1qگ.ː/5ϯ�܎�f[{Ŷi	�#�X�R��ծ�l���r�l��Z���j��j��3[Gv(Y����q�;Nm9Y�_����;�tC��
S���7�`/�?A�<W��8�H,��Wַ)�2o+��dW0̶�g:X��8�"{$E��bl4�9�p+�I�O������1*�=^z���p�����-٤R�̽#WV��0��;���xH���O&\]�T�oܓȡ���j���;��I]=��U�U?�����e��M�T5�Ǿ���$����s�w>B�Njz����-�q�p��y�@���ƨ�Y6%u_��c{�a�k��W��齣�$f u��E�c���`S:�['�����?'���f��q�u�|��o${Ud�Qٜ��Y�NJ�J���5n`@#1��Y2���/:��e�Lt�e�/��G�[�P,�@vd&�,][֕g�ڑ�n��}h�� A@��I�b��ۗ�IR����٢���wcs�C-�/��@�E��q�1�v"����&���;���ejܐ�(gowT%�nW���m�k����*�.�9�n��7o!ކ�ρ�'�]�k}|�]�ѱ�;��W�����{�em_JXBN�!�����o��ͭf�6S� �3��򮱰��w l�O�k٭�zYy��ۍ}�)�V�޷џfڨ_�Gd{���y��K�~uС�������	�s�='{.�;ly��U��V�:ᝲ���a�֞L�����`0^������3�)*wY�Td�y�D�����oC�|�bU�ϵq�|�EG��Fg�I�oe7j��}��k�~���e����q sc���y]+�N�Ӎϝ�{�RBڕ~���D��Ѭ~Y�,O���G�\gͱ��!��:>�w����,��������%��y��*/+����8w�/d��Y>�n�#�X�~�wѬ�᪰�WI�n�+�[�Z����<�Om�3��p\AK&%I��e���4��;q��Nm�*���Լu����iU2�ڕj�M�t��5!)��EvcxS�{O.m����׹���x�M���5J�΄\"��7_p]�-F
f�>/j��X�p�#eh;�ں��]w��	�Ygk[���΍T6���S�n�b�`���U����$�N{�������N��`JJV�om7x��=uF�gE܃&l�5m���'+���v_����.+�{��&��rR8��Ǽ��!v^�z����cԤ�q�yh��OfU�s��os�<$_u�D"ۉ��7�i={Ʒ;h�3��5J�=�NQ�k:�/j"q�l@��O!��x�C|��<�����;[;q�1՝s{r��� pBl���N�9=dt���=9u�^���`rΔ�^o�b)1ۗ#z۠"c�{68O�A�˛s����7�{u���O��u�X'�^�y���;f�]}1����c�"���t�?^
��:��׵�bM�yෟ(}"�t�\6��r̎1�;oё@�)�5(к�T7#�I����pm�T�������&��vǭѲ�=D�2�fs��x*5҄3q[39�ykk���r��ݗ�����i������2�L��;����ӬmQ����z_i��Cf��e���5ڇ��]؍�"V����XXa�B���t�� �il��m�x��H�ED�7�tPg�d䜋&���}�}T[~ޮ�V��*��f���g����X��X�$�v�w�utAF�T���6��9;��x���S�YY����_Zh��U��%���5��҆����[�'na�Jwr\���T{ǲ�Η}w�d���;�>��$7s8���B+�����M�ok�������e4��i���+{j�;�86=��f�^f���v����}ݜ/��h����V�����S��fz��'ݩ�R}KHʝd�:���f˚��z��X��h݄_mz�[�u�qa>�oo(y���v.�zo�*f��tl�n�� ې��Y��C�n'_7��)��F��*�I����U*'�콣�'"1� �%���;#Z��[��P27U±
��3�W�ݍ>{^�{P�)XL =Dm�H����X
��v��S �\m�xE������Fb�T�*�$�kކR޼��~6xeQ�T��;����t*�]˪�L72�jt��u9%�q^ҵ�Z�r��O�^+2��h<�k���6«�{����Q]���SW�t6�p�yDGE�}���#�ޖ���J��3^S�}!�;�9�e5M�c�j��nö�U�+���fۼy���;|����ך�=ڇ�r�%

w�ݨD��v������V�������|��D2�TSw�or)��	�8���ܚ�S�-㺬�Phc��`��(�wD[^Z}Z�V�6Šf�O-jœ�~'�k�*w�����i�`�?d�.��R�.o5υ���ݬl�{+���K�)||�wA/2Դ���T���k�V&v���Zu{٬�(�&�rP8E�)6�c����u����.����A�Vy����N��$^���V3�V�3�SGúv}o��{3�<�،���q�Ch��~���G#�rwE�Ls����ܹ���cr2���y���dS����ɣN�j��o�r1�V��5��\A`G7 Eە]�����yk^�I�kx�����{)X5P��q�l͈V�� �eD��+L��u#}*�s��}�vuƳ�R�]Z��5�c�FH��.�T�-MX���ŝ���bkSA:��U�:���9���n��X��S6��.9�J�FD���
 ]�:J^�|"�������k��uy{2���]��_:Q[G|6Y�!?O!p�z�`�MpV��s�fG���_#���S�ߖ��z���,9��Ÿx=�g��ژ#�DQ��+�u���`S��A6�o��{G$K��=Jt�������[�V_t�Ǻ�+�X��UhR�[�����m|�ʪ�2`�1�=*򊣊K�Q�TR*;���%S*�V�X��p�7�xWͧ��j�Aiq~ {�*�^Za�/Q �.�ث�:�ⶃ�����'놃Yo��5�vn�O�L�u��jw%�*1����������l���Z{��ͽ�.������V[욗�TFS�znBs�G�͠G��Ϫy��8�7���PQ��2;*oZ}M]�ƛ{�.�l�i�c��Dc�[�8g{b�}���K���r��[����^�Ű��D�FcJ9P���Ľ�dd��c�ŧm#���P�x��R��y]�sn��4:D7�;��������k,>�n�Iv�6d!q>�by%ن0;]Np�섎�q$ ����o�'pnH�q򈬻��4U+^
ŷotٷrc�TCH�݇����p{��G����q�gCa�Ӌ�-[o}����_k�a�1�P�s�э�r+	�Ƿ��:ﱈt���.v�]�Nk�ϑ�\�ط��X�B*"�X��rHs<^i9�C���*�:[rK9��9�z����|�'�5i�ź�V�7j���/����̫>�iv�-���o��oyV�7&�ϵ�T����	8ֽ�mG��S�o|$���]�QY�M|��s��үmҕ�����^��k��	�my�����uG����W�\���y�O�*G6BVrH���m�@{%SrU�}{�{�j��7Y�F��UU���9��N4�:���8�v�
|-��[��ľ{I���l�!l>�S�}'�R>�閯L�^�1N/����P�����կ�'�qF���%�e�~8c%M�:�5�[P:�n'q[A)S>Ğa���,����V�h��Ed�ZɹwɌ�#(��[�V���:�����"�_�����T���^�lM>8+�t\ְ-����6�22^Ō`�[����e�%�ӜKS�Fevޫ�.Ys�v��A���[���H{����guu䕿��Pv�;m��U^F�{�A�n�Lr�d\)�4�g{'����ÔFff�Lf�^S=V�I��L7���ؽ�훐�� +*?���'W-YJە2�����\�M1�Gcܯ�u3x����}���]B��$�>�ι�VkK�7`87���k�5��/i[/C�|�Co�隰rg}�V�]���wk�e���`0V9��g��5�$sV����61�m��͗[���r��B׳A��/< ꡖzN�����~z��C�Xg�Z�q�윭C�_�db��9�c�$9Lҝ�W����p��C�p^�����b���Fo�9��3M���w8�����Y�Is��VE��B�t�g�N�M �q��;J^��N1�F:��Ф1��w�,����j?<�0�vS� �˧��p�zyB}Ծ���L��C�4`�-˔�2cu���[.��>���H�6��Ꭱ�J�ݒ�S"��u��m5���
��A�B}�3�ӵ�P=9��ҧQ��b}�rNʃ�������d�1r�.�8�6���8ٴ���@O3s�I�"�h�:���ȋ%��w諭��<:�?W�������R��-�г·�#^�����}��,A�u��c���M�w�1�E�V](9���Y��ac���F���vg(���e��q���%��\���s��<�/��t����<��χ�����`�l+��A�wp��{^O��O��\��7ל�m��D�ǏL�Q�{j�{��7*�?�YSM7�CV���yjm��AJ�6J�lz��e(�勴f�i�qP���%�9�w:���m�^��Y��0���j��gi<7�y0�f��5�7+*y�Q�;������7��\Y����}����f�荗��b�)`���j�-7��f���&Ǖ[�V�I�K"��PJ�����sH۞]�RN����zB3���ɇ؍�宜�*{�z�G��Dcf�{����^��X�2b͛>�H:�b��k^��P�)��G�]:wi5�s��BA)�L
HWJ�M-Y(d�cO�άtLfn������� ��
��zJwLЏ[��WV峗E�P�݄&�aȥǗ�YV���2���5��ڠN��ƍ��:�n1βX)fĦ�JK���uM�ky�ʝy��;r�o_ t�����S��4
!�'Qu�ϻ�X�!۽N�i�8�#���K ��$wb�����Q��K7,;��',����Y'
�PlkR"���g���}NK��)�ezo�Q
��8�U�a
=���7sj��[m���IM����4��.�GBw2�m���0�	��ޛ�����a���h�R��]�%l�ݾu�2[��/����R�`������
��JہU�F�	{�G1K������7+����RN+7+V(w	c�Hn@{Y޺����n��`���+7Yo%�k)�ߵ�D2U8��Z�dv��Y6�톘�XQ����3�;:f�C[��C�9��
	ӫ[&Jm�"�k�w�mt��VW,V�Y�M�G`��KZ	�����K�o�/�M�=�-?,x���ri�3on�'8�I�˸lp3vM�����sJ��]kb���:��%9��X�x��
�ht��w!zƎ]qѽ1BgW5٨�A2���t�T�$�%A[*`-��&�+M燇�-�����Y�`kӃ;���T��!��h�+j��f��Ď_nX��s.���1���P�.(���4�2��E����..�eK�Qi�G1<f��2��R��v����ʉvEol[���Q����F�jmHL�|.�����3x����y����6-�E.��J}���j��aU���2��"�4Ӎw=��8y��A���BP���h�o�����5��u���ݺ5Ε��w�[��w�ƭjwK�:��k��7G�i���ɇy�֘�%�;pK��V��%�Y�q����wY�謽if�Ԓ�QL��yr#�#UҺ�l;8c�f�g3	}F��1��o q���=!��N�ǌ��6���ټz�Ѝ�_,
�6(�<�%��%�
�6��v����`�V�SCծt���%�Z�*M�ūZ�3�j>/q�o��+l�"�t�y'h��LAHo�%�����FT��<'��w�#��.=��|˜3�̊���;hچ��;A�X���fs ���������<ͭHr�'�����:a��K��܄��M��K��N�W
#��v�MWL�&w;dΥ��J5���"+t��i.�/3X�V[1Ú�NΝ&���m�ŷ�ξ�Gn0��[��Z�h�a����6�,����b�����s���3�������*;�յR��S��(��fuD�� �M+y�\����5���<�^�
��y���ۧ rU
K*�T!ٗ�X�}��9�+6��y����{�9e|��P R��i�%�PU@:s!JrR�C��%%4:5�EWZ�p��)4��I�lm��%1	G1��,e+Bh4�:Z�;d�:9'!�V6di)�
)iZ����ȷ8��4�J�:4R��'$1U
S�tTMPh(��CBQ�LCJSCS%	��!C�)M#C[`)ӢabB�)J��hZ2P�GA�
Hb������4��))�Z]�
6�֗kU��B���̠�5t���c�MA��7�w�}��R+c��[���o��8�����4�1�Er�b�S��	c�������<�*7���gj!=�P�`��یw\O��C<-e���o)E��xt�0>������v��쑻7���&}\�2������1��2�n]����MOt:\�>gn�kǷ��}�6���/�f}Nb���i�4��(�m�>�<�����.R\7·=Jw��~@B}ԃ���Ea5�&��r-R{2��W$��ii����yrËpO\(ud^��;m1�N�,�ݏeŁ:������4������jb����p=MI=ꝴ�FU�S#]�q#�7�yAv�Po:}{G���Fvr�;��V���tfu8d5Ek��Oؤ����=<���}��\ϳ��E5v1�2?%�?KR������������=�^�n�Cu��<�7�(W�c��Sٍ#��6��Q*�꟭��?]H�5������_��_�?l�֜�Kߑ/��� 9��i��L�ff-�Q"�UE�p�2�y���3��� u�\�aUN6���v@�8�֓S���!����,�@��VNZo.�
e���qy�w�.���u��f�*���r��㤹}�ڧ�B0vi�/����5Ҿ�����qI��Y���Ψ�k����BLT@Kj���JzY{�z	��u�����9��v��n���^���/����2���O4�8���ܔ۳6�	;����������l�i����y]T�Ϸ�ٙ����ٔ���g���4z�KZ�^�Ű��)F�J9@A�9񷵋�2+��9�w���!s�7��q{�d��àc6�F�Թy�>B��0���g�avգq������׎�Ϥ�1�[cs�("�1V�����ΰ㵬	�0��^��Pr*���U'=/W�֬:+�:��
�pme�`_N�7�:�Ԍq���R\��nNv�7�"�	x�y۲^�Q[H]��2��q�{���t���ǽQ�������O�d۶}BY�hz��ls�ட8���u����V<��Ϸ��A��x��&&�`Yc�U�rNH�!��Z�O��T(wÉWz/�\��C��R�l�p['n��
��#�v��` OX�������5�ʼ�ܷ��蕣�+�f<S�i5�w�KœN��7�{���o{f�V0В��5����fr��uG"]&<���.��}�-������}*Q狉��B��gN��蟼�z���'wy���Qa��V���I�9ûp����[��i={�ᦖ�>���[�l,ɽ���-�[Pw�^���}��#�}^�g�s������!�=1��T�x�=f�D��`%AUD��셟*U*%L������o��Ү���|���2շ^��^�f���7`n�86V3{(�	�.�gp��*X��R{uݏ����l܄纄Lr�f��sG/L���]`����8���Gcܠ���x���k���g�]��X��lBj稾?{���������P�G��V���8�y㻎�nIGL=fWkS�Xx��wjV9+.}���H�}�Y�m�z)x�ҫ�kV�;ƴl�4q^ތΣ)�h�~��׍�(�T�ٽ�%���\��1A;pn}!$�s��^�X�;|�`kή]�U��.}�4.;���.8�|�9�cz[�s�`Z�ב�G˗���Zn�� {��Q���8��G��໵*�2N,�uc$XpNEk�wuھhn�b���nWE�Ȯ{��(�q��9�x�_A�6�:��c�z5EvH靺��ֺ"O9|i����s�n�˛�殹�/����������U	��]��\g�wYV-��|N�,�W.�0v��!�}��u�y�u��C����(��3����xKٲ���{¥�|�ȯ�:4:f���$��u֯tX���1o�~H���ʸ]Mϫ�)��Q�z���6��rϰ��� �~�/�\�^n?�-�;{G$K���9��[+8>�,tŷ�X#��z�-B��������2�)�{Z��P�ʰ�k��d�=v���%P2�+:�O&3�&U��f��p��7�h'�hr���G�NDb��CԎ�T�k4��-�:	?��:t�k[x�5i�yP�x�7�����l-�0�gj��)�&�ϫ·}��'^�wO���b�]��x�I2�r�p�Gn�����l�g�=�]�����pJ�h�� ��
4�[�x��t����"v"k�`\�k��g�w/m=�;�*��Sf;+6��gf�}&%�H\3v�T��w�;n�����;���=��sa[l��o
��EE�#�3�W-ҿG�c���K$�9[����|��Q�j��χc�-=ފ{{��#��{���]�����K��ڋ6���j�=A�,;��|�ާ��>v�6fV<�c����ũ���<���쩝6݊�Y�#Unz�����'���F���	�FX��e���3nE=g�O��Q��v��E!n�Qٺ˺ŚU]���ffk/S�5&}����!�L!����1Od��Ɲ�#�B��!��ƍc�Ĺ:�W���^-�pת��$U�{�ya*�SHHZ�}!;���ǻ��.m�/4_0���V�fI�� �=�Ri�B�Y��qZϟE��qw��Ogк�����κ�C����Z=z�Ӛ��U'&Z������?Z[T8��p!,�
Sյ���_�њ�[�uKB繀ms�ﶛ���ڥ�-�����{�z�zV_K]_�-u���=�zqض���;��'����,-wݜI�0LC/գ2v&Q�6D�U@��\U��o�H%���o3����|��
S�}˙ø�&ul�����&��y��^�ح�ySsf�௺����ζm����%r6#��v�gծ�����e����&�P]��Ο^�ɗ�z�C�e�@=�(ɞ�j䛱\��q����s�/)IXڏg����ׂ5s��ͣ�o�z[Oih���'�l) S�4�c�+NK+"!Z�c��ݿ�������]�9�]�����~b��E|����mR�����ͭe�̼�&G�eR3�פ�yJ��fຓՂ�i�ٞw`V��^���m%Qx�z�Ѫ�/8�C�W�3������V2/B����v�[��{lr}����Q��p����rTv�$�vt�x����ԯ`�Fu���>͋�;��^à͸�f��O�9y#�"����kf��"/��|cӚӬH��=�M&<�F-���0���N��3���ӑ�7��� ��K��^�0l���_5�4 +7]<"�K��b��u��c���w|v�� S��.�c�k���ל�-�ڂ�F�ֺ�
;F�y�C��6-��	kԵcϘ�c�E��V�ז��J�pT������w^JV���z�%ǎ��9ݻX��޻�[7�r������[i\"j}[�5O�#-�I)�d<��j�Ҹ�}�����}�;�Cs�t�m�pL]��/�2z])'���8�9g(�dvknz)��
���dc���^kɖaF�v�D��#���kٞg��X�gu��F��cޢ�`{���c�}��.AJ��K�N'���]��s�ys����~��2������N����>ɂ��掛at���!R�v��xm�D�'u�����3�9�^��ݕs��lm^���8��]�8��s�%�^Ŵ-j^t��7���<��dS��4��6���g�j�uW��N o��*g�%+ߛn��XhMBuS��G@�c��ޖ�l)���AJ�0/���);���fL�F/�ܳku�-�)R~�ו�>Ǖ5�k����y}YP��3��St���2or��ͩ�bL�1W/��/T���C��=�~g�.��AN��� @M���\�= ix��/Sv�������kc)�mp�9aVvT��y��V�������-=��y����:06��\\[5,G�Q"`}���jE�����ΖT��,��h�fP�����:goh��;w����ȝ�v�2�f�Q���p<�*���5�,{�ZV�����]������U,�B�Ln����Z�xc��\��~:�k�X�p5*Y��	9�μ��}KV���׍4�J�D�ek٫3���f���P]��fk��#��Y[�oӨ��JS�m����â���+xU�er"�i���5�����U��PT~�B�c��'�unZΞ���[cG+�ta�����ߔJ#��u���^1q������{��T���bʅ��ϭ8F���^?����p�w����o�p�ʓ*K����Ք3����^h�c^9����L�k�#�[��+�^K�r3�=ԓ�_2��F�O(O�������F��^ܗ~�B�L�g�vWo_�+u�=��oRu���\4<s.*��=^A]�Ǜ@>͛�9"\m�=Jl��Vp}����-�M�H�Vu�4"ܗ+���:��A��Z8�9����A\Hƫ�|{9��Ƈ��vq��OA�K����C8����T��[�w�[�QٳR��oV�U���7wXƍFfo'�]ba�Ť��륒O L�Y����0����YD�-�"�_K,�.�t1]ϲľ{I��kΟ^�ɜ��u�:Q{�F��A�E��ju���^.b1���]��'�hr���G�De��כ�6��F�~V|{�Y�G-�c]mmM}�����[��O-O��q�F=c|��V��b���_�������h9]�gǹ���m�^��N磘����I��&iOľ�VS>����B��N�����p^�ŝq����)�f�^�_K�i�~[00R�d[_,��!\��4ͨ�g�Z�U8�m&=c!��P]�_"셵��`��Q+����ַL�:q�WCs�\��z�>a�q�Hl��5�S�	z��T�
�+����k2ԋo'٬��KI��یw�O��C+oҨ�-�Y�1�Qp#����E}��j\�M\jw�U���{>��f�v� �sgv�,򥒦��|�E�7����9�9/A~�r�C����&)���(W�7.S۸/��Em��\[��S�OH���� n���d�7���:�dN�띰&���o�v�y�v��U�uN�����Pƺ����he	P<��:��!�࣋��á�=T�<��uQw�]�[����̵O����e�8�`�rc%�{B�*x���\�ﴘ��Н�.���tX�W�쵾�"kpӸ�c�T(�Cy���2m�H�_���u~\J�O\�۽g9{0k�
t%�3uԶD��2�7w�^�n�IKH[=ih�aɞ�dy�X�={��q4hk�g�͞q#_7�z�o�JP����+ǽ�ߓѸ<;�M��[:_���-�X�u)���|�]�>~hC�<2���.��)�Z��Έ��zQ�8������cwB�n�C��u��%	���w�ޞ���S|�Q!�`%A��T���+h:�R�PR~��S��)؃t�kb*���ܗzny缩T�s�8T��#��7���'�d���o�6'�T�x��3orۋ��7)�����D2wdX�sPF1!d�,�l�s-���U=�W�4 1�(y,�̵*L{{(�P:%��ǂŝ��b�ƹ�>9�sSK��o�	�r�cO�+���L�uWsZb�]/t3oۙzz�p�XihtF�yɼ)Ox.[9�y�^T���6��:�b�#�m�(̑_�
�$�뻋�{�叉��e����.Jޕg��űA�ݞ�5\��Os�?]af�)`ڂ6j�u�z�{�8� gi����v�4��Φ�wZ\f����;��2iʰ��j��|޶�N��ec/o�2���b��h�'��!�{���`Jw�����"���dLda�sj����R�X��r[���X�dW%���\&)��#�NZ�n��yz��T���0e�QU�5�Á~�,uV���$�E�-}7g̓+�]NbR��ն������� d̺k'��7p�:v&OP�˒��A�u��y�bU�g��B|��!��8Pۤz@!�o�:w��}��:���V$5�ㄡ����.�Yx��[�^d�l��
Z�V��t{��Rw���Z���B�W�v�}n��t�]Yp;��g׋+._Yy� ��z�Sg���S��)�;�d꼡}��`�fA+y'���ܾ�]c�t�E-��GLVjæZ��^�eX�]Xi�M� �Ң��G�+�6�ЭHL��8���]�٣�h׫�2�����dgU���z*���z��cb��lѰN2���/j������~��{[}���iK��g;-�ɢ#��;�p��l�����:�[N���39r[l����S��7�����n\��!0�v^<���;��b�;�(W�mN�0u�N%���nmv�"��S�;R4�m_N#C�\.�D3J!%�	lg�*�V
�����#�&0n��9Y�Ӱ�J�>H)dWt������w(���������΄2�1�8�j�BoQU��k��ÀHg�����ŇK����$��Y���8���6��pмMs�W�b����f��{;E���D����h�K�h��}}��iP-;��5�)t�֦es��p��s@�<�z8�k9�X]�����J
�
P��@�Ë"V�:Y�`
���%!�.���ѽƅ�u��MZ�.�4�^Mj_)�x���x�o3�X�(8g�,Eb��NL�sE��WVwU�J�$j����
ȺݑK_=u�R�ݬJN)�4���ywb`�S��2�lI��ݒt�w2��
�S�<m6���q��i[]k\����]�.R{�D�5���@��u������؆RT�8*t
������v=����}R���c�OYy7�-v�wD��qwt\�.	�7���ߩȸ)SU�90�:F���WU�Ҧv����+��S��v"����<3��ڼ|�Pv6��AY}:�w�əlb����XD5ՠ�k���ܷ�]�1̡K�B|k��eu�nVE�]��I�� �iԫ��I�ͫ�\�?�u�=C_���CC�h��i�m�HU�Jh�ӪGN�E$ZCE1&�

�4�J�Z�6MP�:hh�SN!t��ղ:b4ib��[Yӈ��i�հj�3P�]	QT�X�Z�h
�:!���#�M!�ĕF�E�KT��3Q�Aiō�t6��$s\0S��ٵ�k/#�	Ibh��[YМ�G-���HU5���������q k�[<�J<����$ӭ&�ZJ�ȚӢ����h�j�%��4�ɬ�iѢ�@�@����i��1��4(jؓT RRK^��b�+�%���a�=I�y����P��0j��$ot7.���ܪ�/S�����c0*鱃?v�&=j�g��:k��n���\)i1x҈g<)�r�]2�^�
z�TL\�F�o��$��	g�PQf������vl\��|��>�6�3a��mCqB��N��`�~��De {��j@��#;��{&C�p�1��`�z��>xun�a��V���w�e�-v��}��ׇ>��h�i;h��/59IZY�9�:#X��Zʁ�E�]�c���e����G*�����k���o�z��g�圦�uћ��ơoh{ʦ߭����}a���S���OiAf%�ZJ�iƵ�t7��#u�{�����',�ġ�Վ��뱶�vv�qu��
��˛��w�ګ�y������s}�c� t��sR�_o���o�J�p{�x/��|�Z|�������2������ս���u��@�v�p�aO��m�����j��$�Thv[+� U}u(�r>�S C���9�*�\�hW��.9�܌^�3�h� ��'��j�:�`��F��is��{�%�hM�Vv�Vܚ�f��N�Y췌����v�a�3�,V:�޾��ԝu��y�2{3��Ku��Qquq	o���3��+:����3�o�AS6L�oq���r��M-�f�y�{�վ[Q��w�>�k�u�YP�:���/��nOA�e��J{��,��gf%�\����}|Gd�{�M[u�٨��8�٧K�<o}�5�o��q[�N�=�^�%�o���l��'=�"c�;�J���W�iܵ�:����eO4�8�w�/H�f���"C�pGo�df�
θfq����,�?C�l����V?Xԩf�V��׏�z�ێ_3W"�+=5k��s7��őE�5�"��[� ��Ys����+�B�
�Uz$�U-��b7/�=r��4*����P)�ے��S���iن�*��{)��Ϋ~ǚ���Z�|��G+�taoF��Zx`-�0&�;��x��WmM�d���{y�P�a�lB~��~@�\S�l?1o�ʕ�(`�U<3��TP�v/�GI�=��t���^x�����qO�<6�:��qF�*`��z��Ү�����[��lν����Q�ݍ�U$E8#��m!g�H{\@w
�wS��d��f��;�Z�*
b�ϤR���b��y!Ķ7�T�����z��ֿ���v��8^оc_^9���3�0�S$����S��$e������U6���w�7��D�=���y���Z�Kd�M���V�9[��~�9j��z���S����&8�ǆ=�t>��^������s���m(C��Ŵ8ոk=�q�{�;����J줠g��Tk�{��y-<R��k�J��ݼ�=�@�0�A�`���QZ�� ��t�6)�5����ͅ>��=�r#,OU�0�Ϊ�ދ�V��0�o�NS.ժ���a�k���i��V�	�vży�m����Jf���E�_D);=���JXj
O�[X�z=�h�����r�o2�h�J�?k�W���ԝYO�/��;̿7W��!B����O�糚ج�~�܉�ar��
w��,c���|�Q�����9�]y�cAS��'����_�"�������eӈ�1w)��k�G؆Ho/	B�5�ˠ�՟���.��i�CLSu�gM�k'T�NY�Â9�ٕ��&�j؀�|�`�( U֧ �`��v��]7��0��d����.ɏr�a�=�XW��N��	uʉy|�:��3w��	.���9j�ё�brO����^��x&��U�M�Ff����ݬ�oa�f�:�	��y/���U�X�t��MNu���>X�M�d����L��Clc葏E�B70��3y��MgE�z�Z�S���{��87g6Ts���.H+z����X�ʖw��"�l��b�\V|��.�@N�B�ǻ��eͺ�ۻs�:�*�Y4����r�x���������Z��]�S���\���-Xm��wr�D��Uw1i<�޾��c'��9I���@=HC��J�2�m'l���I���k]��~á
o�˛��w��'*'��-��Khq�*Z��������S����dm��ˤ"�m���8�|ظ��\��[x��g>C]��Um����hv�¶n�q�G���S�m��}Z�z�a'�u�]avU�#%�=.�S�)��j�8�e�,�w�t/li�fAz��Y�����{Ӝ�3#9	��u	��[o�0b았�Ԟ�\�f#�"�:]vu���N�w7��6�X:��l��H�m���y\/;�B�d��x�«zV(������>fՁcw��F���������F7u�a�}�����GN&N�ի�r�VN�r�\���L�s�8��Э�~�X_!7�vfp���pV�~�[�����������a/�|T��I�B�6����ܞ�M�G<w�����ܿ7�훔猎1�o�`;�՞h�{M�ޕü�K����I�9�jZW�c�2g*%�4�P	^�U��b�������c��CބI�}+��K4z�KZ�^�l���~�5�)�g�c�L�ޜ�ޢ�?P��^�-�{]F�Y5q���n�p}�RR�p���u{���*���O �Q�;�~���vH��{Y��W��ˇ��Wm��y����qǸ��9�����O9=�,�M�_�����'T����'���՘n2���j�����7#}�ܯ'�{<{r��|�]��c����xNov���=�>����d��Px�9j��o��^M���L����r�t ��~o�a���t���:鶠tؽ��9�a�X��R���9�+BՙQɴc�Q��W�����>k�waIf�����]ї�y�X�q�2���֍�L��Q�ϥ�i��9�'���u��8�:e^�`���3�Լ'F�w)Tr�S]�=Ϣ���pU��y�㍳>6��s��QC�,y�~�p׶?{�O::�}GԪd�)`(�s�p�K���r+�^�����a��5��[��v�h�it��D�_�f��xM��ʗ@r�a�B�lr�������O�>�U��Ѹ4L����ޑ���N/i,3N��f|V�u�?L�Z��i�gu��k-E���_{�v��S'�c��J�޽��]hp^u����T���Q�����,�T��n���*}�3��@�]��v����ˊ�\�e�����$�D�b*�}X}գ��v�����(�J�n����ytY�n�U���i�#���K;qخ�:k8���Y�p@՛��_t:�
�ܐ�z��?q��Δ5z��*���C�޶�"|u}����L�X���g����]\p� �
�.	\���)a\=�CG���}��u-'bHc���ۜ(�m�D������2Y��9P�&
��2��
�����dW���� TVvV]MȂ$q����g���A�ZIl������,�٭���Ws��L�=�
ܾ��w2�PV0eUt��]�NC��{�����x�q����Bvj�z���8�׆q�6���6��k��T�,^�vcl��u�%m�=�ÎIZA���螢s�4�&��h��'�L��d4l�2�����*�v�qɎG'�2K�o�.ONjBQ�./=�����H��������5�s:/�3/�F��/k���������oS�����zx��a�8�0�Wro�{��wu���P���x�y`6�j�9����g���WYu��`}R��t����2���J���Xa=讣q�o���ƞ�>'�S-e�{�5��kBU��HO}��c��Vu=����I�F�1׹w���N�z=�>��^��:/��N.9ы85W���t�l�T8�eܫ.7x
��a���5�Np�b� �s�g�1q���E�C��cQH�O�{�0~�ž�Lf��mƆ� 5��k����^>�� �>#���{���T�3��tO��99����օ�)�}'n.x�2�e�ѝ�W�uR=��>��0c>��[۴�s�i�A��:�������T>:��j�4V����9.������*��HIY��;F�;鎇}B\�>��z����������DW;�^��b7�+�Yʨ�f�����G�e'ׂL�%T���Ź"�0�����$�s9ẠK�vU�ڈ��{i�ρ�m���m:-7T{{՚�Ƹ۹��t{���DL9�a�UC���FK�Y�g�Q�(L�.�0�S]�$�jî֗5��<A�|e� �<.*z���n���?:�V����G!��z;h���w��ߙ��Ǖ&�=�lz���_@�:xi%a�~"E����WPz����^v�gX���,q�>��w][���ٖ�B��]}q�D�ϙ5��I�W�#!��u	��⯭�ĳ>��#wmc]�]c�r���4��wQq�lM��� 5#���t����է������J5�މ��{����#���{�+�����z��m̒Z������0���{D���{G;���R���@��7����W�n;��<}�9������$R�s�s��S����R��^�����¥J�B�����1Sӫ�G>ک1����=Ǡg&j=��.�:Ǵ�gopʌ���$�Y�]L-��0yexe9�5y����]�c�'�r/Ϩtϥ�QT' �Yn��Zz�;�=���ʐt�V|=0�a��՘n��<�!+��ܼ�^Ǥ�����J�Ym��Pfo�V��;��X�Qu��� �?�f ��s�S�p����va�A�0\��@5ovSu �{J},f
���Ȁə����F�	�������p3�ĺ7�w�WZ��)eb�rtWҔ8]�+r:&��&�γ�S!�uK~��r��)O�W )�*�����`�Z�31l�}Ss0_@E*M���T�_�{�m���}���+�`���h�w>�덞�>h|�TҕAަѣ��m'|K=�.y7qř|x���w��ƥ>Ӿ=��N����������e<�!<&X늜�����O�2e��0��o����>����G����l5��.U�����s�/c�!��_�xz��,I<�}Z�2�f�?��Gh�c�;��K�[�����.թ=0�J�#��\��
:I�(?��WK��#q[u�_�~~�7��&����{�7$q���Mo����g��f�n;����u���R,��'��! ~����_����̞tH��6��߳�Vߦf�ODN��>��<�}�D=7��e�>���ĺr �5X��e���D������1Ҿ>�ʱ���|�&�:��>��s���O��ιq�l͹�Y��iW#/(��:��6�-���U�<���+��S���U!���[f8�k�GL�q����_�_>�ur-)��y��V�8~�l�������h]9�9�
x7����j�1�Vx��s�c��K�1m����f��2�/�q�x�5�!d&�k�k�fk]�3�.�fSg��������������׷K:]�S6!+�9��LԘ/��hK�=��]���j
��Q�pA���^4�2�WL���	.�:ҺØh� �yg�u�%�X���J�������Q5�vNؙ��;�/k��k�Y���n�p�|��9��GC����W�3���΁��ldD������T=5��ȟ�s�Oq�̨xW��˷1�o��L��)b�9�ޫ�q����O{��\oz�SĪ�|�����+�0�ex�+�'c�^�G���T���g���{o.��>�}@t���u�w�ݾ�p�dϯ�>����u/]�°��e���C�}�u!��i:}�����W��a�}��uPw����7m���½�/��װ�7ܲ��U�K�r#C�J�9�ɼ��*3����������ﻪ�o������.���|��G�_s�-�EB�?��?���O�X��Ma��[i�K�E����^������\���[�����++�i�϶����t�Y�R�|gj��9Z����pn�}ǰJ�=ZѝV��	L��)|�r/��Sԇs�ж�F8��N��+�|eT;�<��w{�H�K����Юs��њ��z{�v���ݷ��9�e�� �.��$�,���P���՚��v���>��"�H�+PZ�)#��ݺ��x��=��A���M�L���Ԛ4��1�]=V�7�� ��ϸv�"�KL�w���n	 �^c�"C���:J�6�m�� [ҋW�)K�Q}��]�ѓsi����W=N��Ǥ�u�����5��=:�"ܦ��U�)�Lb4X�x��0�]��^��0�	j�WR�Ԧ�GT��7�լ�e}\V�e�T"�JW�o7xx��٣c45���n�Ϋk��f�,�=�<��r^jn���7==H��]׬nG�Gn�*Z�������s���T�YR&	VuK���}y�#�ՇnT}b���;!�E*�U ��1���g5ml��]�ՠ��x��Yl�����Y���n���|bJłv���]y�!�sZ�l�`x�H�0h�f�ܲ]�+��C�M�����'c�oW���+.�d�*t�<�q	����c�����ZӾk)3Ӎ�u�$h-T��s;�E�k�4�ȃ1�U�ϻ>:�t�{Ե���tV��(M��# �׳-uF{���M� ����GA�������~ୃ�n�%�[t-���Fe%V�>uY|��"��LM��-Ԃ�q�R�Ȗ1�1�m4�@���,���9����.�R�9���,<�$��Ҹ�%`�V������WX�3��[�w��/��u4m4�n��K�RBm�s�)�
��w��5�&T�����`��9ʈ�*JLP6u�m&���z\=ٳ#\��l�c�αR���A��ӥҽ��FT�{}ft���2�'�N�]�OjA%D�Z�\$��Y}�h���( ���;���g�0A�aƨ�9�5V�ۂ�7��Fo��i�v`BfA�m)��K�ř�k%�\�I+b��Ϟ�y%,&�v
�-���g>��)�>}��d`2��2�a����#�k:����qC��3��÷�M�;5�aAǹ�+e%�G�oo	����z�/�ǵ5�Rq�MY�B��չ��{��vjN��I�}���ַ�v��ݗT�Ü�$u�l{,:a0�ӛ�U�R�M]�
���,uc,P�e M�N���]��b���쾌�g4U��R�ѹEز�έk�c�&�E��J��3�ƻNC�pYg1��&��I�=#ӫ�{����c��n�i�У3��3�mm���h�҉��r��u�E�u�Sҧ��	<[+�e�]r�x�a6�r�Om��Դ��h`�xn�aT�kg-nq%�z%��;4�� z����/j#���ñK�H7�2Cö]E��`�ȞP����Mf���X�⃜r��Nw71:��-�٘ڂ�,o%�6r�����=km�`�T��52��կ�Z=��Y��k.ɶ�o�Ap˻mN׌�ż-�*���&V}J�O��;�=r�ڋ��rʄV��j
��t�ko뺺`X�"���"MZ��-�hh-��*%�Tk�i�m)�F�ڣM1P��	Jֶ�Bb�I���(��ւ�S����ƃT�i4D�M��[͊(���#�G6�m�F��h�ꀫjm�I�!�����F�F"��5KM�����F՚"��������ŭmgU4r5s%�kh��cS��)��m�AkVɶՋ63�-�X6�0��.��T��6��jتt�5h�����ZQM4ţ3����(���Z�)���)�X��nZ����KEm�Zj�Vb�)JF�����I�Q%4�Ӷ4��lPST�E!MZ�PQ@Df�")(�ј�(��|� zS�3�W:��Mh���<�׵2�`;-m�Y%�E.U�����l��M�\{���������UP�y������@��	K�F���[,z/���v��^�}���8�>���*��:k8���or����U�Â޺"W��6pt���O�������C�oz�<������^}~��A���>�Jg����\�k��� t�{$\�O��������0�6�n�O8��y�56hd��f/]ti=zKj�p�W_\M�QfG�$W�};&���������W��ztD�����?a�w���eu�R��~�8=�8�{�9��W �h��Vzo�~�n���^�i%̡g�z^��1��Oi�ﻺ�=�\ ��3^�wLi��ό���T��)Gy��$�8��G�W}S�r��t���]��|������]�@oz�{=�P�S<.==3$������g��3atT���xu+ˇ���L{�{�]G�?U�>�ߋ!{!^�5�^�x�Wq��:{�'��9\�u=�·ZN�v��ʯ	�/G������	A]2�V�s}���`+���X빛88�{`�.�9�׫��K�=��+=��\;�1�#J����
�0(�i���ٿ���x����l���y��C*�v���#��7� �1�,��oe�śFa��)��铘D(#�m-��C-��wavхǜ�޽$�T���ǣX��Nخ�	�2��%9�[}tt�����/W��|4��5*P�ʏaA\��r?к�j>����ʹ�~�<Ne�f�|yT9����|J����ݴ��~[���;� �-vA}/�K��Ƨ��Q�m�r�v�|OFPIْ�G.Ϧm�-a��3�(n�$z�;��������|{s辸|W��\f�v���S�:."�I;�N�!���q��S�VИ'uL�L^�P�8�h47����(�x{��+��&g���^<ꁕn�U+��(J�|g[��@�XةT���t���άSޮ;GJy%��H����w�V�-Bma��yЦ�L8�x�3��Pe�"@�ښژ<��o�$_��^���&=�w��tgf�Q¯���7�w_\w�\�4ȁ��Á%��n	\W��5�y��dc���՛jꧢ�i����9\����Hi7��#o��&��r��ϏI-փ������#�}�J���t��o��*2�o���Ӛ{�}ӕ��wu��o�4�q>�E�C+s9J;�#�u����c���%q�����F�/�����Ȟ.:g8��5�3L����b�_�:~�aI�^��:�>�}u�Wݘ�Befw�p�y�'�W�yӺ�J�6/%�"n�{\NlJ���ؔ�)��)x�rx���az�e��p�E�MPA̱�6��԰�e�T�[|�Z*%�Ϫ��eU��<r��G~sP 
�5���-��1�J�᝴�q�N��g��f\�
���4.�V��ON���+�1q�Y��zw�Q#���O>�qZ�~>�-���4���mz�'ɬ��=��3)��J����CME�ϕ�v�T+�3���S<��n#��,ozd<N�釶'0º��7J^�Y	_�O��u�ݑ~P��C���G�F>��}�A�N�mX�W���d�� �T;�W#O�j�U}tM^8״�y��j���-_:��%t��R�u���e�94�^����'e(�$�n��k=l�v���R�F�gx�}�.ys��
��Q�9�W�;�Ʈu�����8;��.�s������6��3��&Xw=GԺ��2�W]�6���WWq�E5q��"�|�nk���qx�`>�	���Ş% x_����L�7Z�2���\����U��g�S��L��z�X��譤9q�#תY���ό��FU1$�r+n�Kv�;��}%��V��u�x�z:7by��m��Lv�)K,a%#0�S�F[*�j�l}������,Ke�%�b��.M�rTFo�sEV5�;=D蹼����p.���_V�W�H�<%���B�A����s�@�X�E<�Wp���Ŕ��c��[%��V��cN�ӎr�':�]��j�m3s�Y$.F���)�V�|v���mD��_a������b�p��z�.��5MD��C��ܮ��rr�-�� zZ_�h4U>W}]it�qZs�Nq��#/��f�̂��+�M�b=�%r�V�x�8x�D�?���qC��)h�=T��u�c�ӛ|�t��7�q:0V.�B��#x�S�dtzd�Q�$5$zJ�4.���<�VF6��:yY��^(w�*���d�/�h�+�d���"}�9
G�ڄ�|���M	/�MgK��kw#�5^��^�`L������]#�X���g���3q�S�\�JY;_!鿏z���f��x�ťߺ�`�=yZ�ߟ�z�f���ԕ������=�he���A�SĪ�鳓��<bv�z�U���^�Ұ�W�C}w�����7����v]G�g׳���;��;�bg}�ޮ�]����-]v��ѻ/��*�P�k�ǣ�E./7��߫�T��Ӌ��ړ��5y�f��,���΅P2pu�S�8.�W��L
��s�p�������y��eF�?�(#�d��D֓6���y���W�˘��%�����X@所�e�E����3u[��e{�否2<�n�W/��z�k�(`Ij|��ػBe�n�n��Ǫom��Z\��"0���u���ߤ��Pڱ;�����f�nX�c���EDv��F;/�8nd��'�b|g}R�^�L
�c��U�sֽ���,]��{#z�*q�z)�q~���3O�}����V����҃� ���~�⵨�֫�:kOF���ݕk*�G��Һȿ���N��p���C�s�Cb�Hۋ�$騉+�Uc+������z���K������^��Y����oOx��{��|��θ/:�A�%ӝ���'��WP��nJp��^uR����z�:<-۫z���oH�����w��c���R�O]a'6�k�4)~}�@n��GJ�nP�����������Cy����'
R=�Oj�&ѩ3�h�K�]��1�D���� 9��H�W)��)a[޴4t�i�)��G��Y=��֔���;��ݝq:n+��%�Y�D�N�����E���P��dP���{OH��lL�T�;����OR'��p2o��@���z&�s=2��Ѹ;$LD���1!/z��п5�o���͸�n5�Q���+��zW 7�׀u,i��ߌ���x��T�3�S쮘���\'f��<�#:&I���^�qMy��:X�ҥʩ�Ҹc��Z㴙aN:c�����<$ 8OTo_Pk��/+J����bY���,<s��SZՑ��KHU�m��ĳe��v�Y[w���y6�\eP���c]�Թ�9�u���w�'��9��ޮێ�ϝܛ��ɸ��7��������%����Bc�/��t8�c��a�t�Vd�;�W���ޘ�=讣qu��c#9�B�_j��c��G�V��Ī��9\�Oa��n��ݖ9�n]���뗢�ߴWnx�FX�F���Z7�����@���/���T��aD�_�fP����Wi��Xb� 8��h\��~�O�'�FZ�;*��G:���Mң{i��H�<O�;:yT;�Ua��< !F�l^��b��9։��H_{��+��I����]δ.yH,S�;G�C�/�=�z��xf�d�!WQ�z���S>=�6}3�gO��_܋��{��q��-�i�8+h���f�>]j�r'C�,�y+�0���)>B�mЗ7悌r�הYX|�_<�;}��n٠�8TΤ*<����r��{�t֒������U!;S��ۚ����u1����_w�*i\��F��J�w\X��}m�o��q��%�0����)(����Lئ��B����]��f�n�j�8S�����h�:Y��ڦn��F��]��t�-���`��������-X��ՂṬ�����=6hY��]x��x7�)V����d=/g3�;��IXƪ�&茍�5��K:��-b�e�KY���',��xBWX�N�^ ��G+)$|<w�v�W2��*��'�w_\w�'�|ȁ��Á0[�&�\W�	�`��-H>���^��h߳j+�r���W#�ӣ	^�6���bn�s_" j@^"ج�u��uMNxa�ty� ��醊�z�F[}m�A��=�#�+����."z��o�2K��s/"jd����U���<�\s'�I��UԽ824�+5ڮ���y��3�O1>31�D����;��Uל��G]˞�Lj�
�;Ɔ}]+\b�����#���s}fJ^t2(I��w���Q��
И�eY�t"s��؞�k/��a�̦5*�M�jÌLk���{�ܩ���9gPS7�wO v�]�[ީ�'�ځ酷s+���7
����o�/y��F(��>�?���ڿ�JxwL������U�;>�ڱ+�H��K'\?�]��
��UV}"�]�jj^Q_����l����U]��W�r����F_�������{��>����z9|�����	��4%.d�I��.w���ɖy��U�Vi����7�RB�뵃|+�"�����d�D��,���/��*g�3�%��]ATXv�ݾU�k��јﶄ�0�fY���m�;��L��r��ɲw�*·6�XV�b8+8���8�C�dǕ$B���rɯ7*'PmF�PR�V�n3�δqͬ�ngGF�8r�X�@����OQ�T��	`/P1N��qN�;������}��#�s�j���u�1q��:n�%+�,z��,I<���q�hs�ξ�NFs�����d7�>{F�ٵ�W�����js��>�LУ� ��2WK��q�N�p���X�<�z��������j������;n;����u���%�gI*��8��m�,��X]>7S�*.��}yw��On&�[�����;��!��U#.!����]9 j��i�9��9��!^�M��@�}�ZUc��v�u�]iDt�qZs��8U��r2���fW�K�~�{��v����-�=`��A�@��A���{KF��C}��1�so���>��Ѧ�����l��i��o�J�;�J$�Ԉ���2��%N3q��_BͲ2�I[�(0�E
��Xʸێ��Ӱ�6~ԳIw>t�)�;^��}B���NI}�k:\t�\{��4f�7<R����t,wr9��y��{��x
}�P�������kk=5�����C��9�NK-���}�m�3\�,����:m���݌�I2|�a�k��M]QpS�k7q_�-������Ai3��N�&�>��ݩe&�6�|�թ����c/a��-�;i�Õl�q��:�����CP�յ.�5´�X�'7s��Wn�n��]��ϝ\��<��sq�|��51��](29|OO��=;��,N}v`��^�N���+JG>J^���\6���HOD{��N��}b����Թܫ�潳����=�sîN��1�
봝>ݗ��7-\w�Mv���;�=�w߬���u���<��ן��?�0e�ڼ	8�Db�h�9�]?��Η��らt��6���kkׁ{o��*����t|��b����z���������̯�ȱ�W����.�����}�cfb��L�ǥWS>��>��`�u>/�]Hf�힊�u��^��=�
̀V�k丣�|���p��՞�y���sxoi�?F�"�:_t�}}\9OR5C��.[CeE��.���ߦ��f_��C�psY�ޱ]�gp�= ������ޮ��d�y��|��W:����j�^�>�l �w��2>�w?($�.#�#:G�)>��ڢ���U���;�>ޑ���'�(�Wk�FDw�@�G�~�w�m��H�@6�� j�3�HR��y�Cнt��*㫭�����2�s�>6������'��p����Am�������w���]۴�����y7;h��x�=���C���nəY�W�<��s��f�1)$eyL�8C���c��5:�rvsndv������xl���n����5��((�x�
���+&�{=[���5���r��8�Yϔ5Q�:bod�)��)a=�C{�9�t�E���>�ޒ��F�u���KI����q]}q7�e����+�h�Qz{/�vvл3ۆ*�)]	Xމ��<9�v��O8�8=�8��ng�j��H�eI��̘��pn�{h��>��ێ�z٨��t��:�5��D3X|�4��Ύ�㤟1�t_������ޮxz>=>�`���9F��:�*9>wr|��d�9DT1��Ή�x�M�mM���c_N�~���]>4T�8."�W
��zm+ˆ�Ua��ފ�##��]7ʬ��M�h�=P�<��qXg��K%P��V2�9=��>V�I��c���|X�;�S]�3ʮ,��X�k�Κm�మ�l�
'2��t'0�Ss����Z/D�U^�	ch|kn}r�z�{��z#���G:���uX�}������y'���<��f0���^V=�5Y��S+	�F`
�nȸ�����uF5=�pj�����v���\�	���6|�E��U�'F���0~KPu�7�c++�kH}�
�jLMf���69\���{����Y[k���	�e��3w��yp����nGr��܇�]�M-��C��e�Z�}����v~�P��w;�´ �Nb��ƶ�+32�|�INܚX�V�{
V3x�l^c;��s8��d��w��ǝ�<Z�������9oN#�{�es�[299�%�1���\��J,U�$Y�x.	�pd���w�޻+��!4Eva��mܽ���ݜ�5c��j;t�����t�8�b�̨�!�Z�����f���흐0��͙-P�)���i%ߖ:�);xz����w�+ި��[Y�H����6PV��������^����N�y�7�i�����̣rF���$%*~"Ҥ�\��̔%��i���V��h����
�5��Q��n�i�.Fz�\K~�%�pC{B})d�Q\����n�[�����7B&����	��`gw2��݈���i�������m`�Ԭ}��겇[]�`Ϭ��(����õ�q<�A��¥�o�t��btك�Uu�O_7y�S ]�sq�a��W��0��7��>�|�H�~�;b�k\#��;!��B&�N��<��N�v��S6�"�U��sCE�ږ'-��Sq�S��	nVڵ��G�V�LlV����Sx��]FR���1�n���|���h��Hjq#�;œI�P%�㷼B��3�H������mWn\8��
��f�n�Z�j����r�I�&��3������Fұ����bn���+��cS��@�>콳�b��qO9�Zb��Tx�v�!�<���:~���h}\�r!�v7��I�3]�Z�b�}�;#����lNv�œ�ۇ�Y8i���!u�ed��S�����W2�5Ϝt>�҄�	IV�^��X���^����Ţrϔ	���Ǡv�;��\�ꆭ�	��g��b�#����Q^�CG���C M�uz{�w���nS�]��g2�^��5 f����8�GE���n�XyԢ�AӗG`�����b�;l9}���V�{���A��yj��}W�;�>�C�)H���tvr�r��\ش���u��Ѩ���W�a%*c+Λ3e�L�p��\�V���W�E�=�����l���s����{�@鞂��grH]�4��܉�J�v\;խ����V7F��A�f�ft�sR/nÕ)ݨ�����f�/ ��N���VU��Y�/F[s��B�?W����u,���qg���}بZ�B����^�q��)�|�����BL�çV	F��b�V�ƃ���C������9��ܜxE�
yԢ�����1a��B�;Qr��9�r,'y /%�ޙ�}���[}��0F'u�t5i��%.oL�^_R�1(�F��_�Mh�U�33u�9��%QIAPUUM5T���DM-A��V�v�5����iuT�U� �")(��]:����"ZX�F�4j��)�ՌLAK�t�U<�-DACCAI��������5lkK�C�f���"())��������(mLi1:5��PhuA��i��PT���4�%DQEUQU4���"�m4��nCL��j��b��fJ)KN-�6Ɗ����&&*��ѝ�lQECK��Z����

h63�KTA4R�tD[����4鈦���cPDD���4��cV�[&*���"��h֊b"JF�
+N��cM���E1R[����A��7x�==�^c��`L��Mꀍ�j�
���2}\���VVY���'�0h�o�!��͘�sh�`h�t�������3�_��~�z3�g�;����|{r���^��T3oþ�qJ���Dګh�_�j��zO؎G¾D��%�t�Ka��܆�P��sAX�L��YX}��U����;�_�{2p*-f�5+fo��D)�F���q{$�,	�bJ�2+n�\���V*�{��D��l�e;28T�&��j�w��f�go��v��g�Y�gI*��AH�_�����[ǵ�����u�/;���#�_^GvW2��Tp��'�_\w���Pȁ��3��Iw����xdUX��V�V�2��7�5��U��y9��w#���o��F�u�nd���@H��kQtx\�X�!�W�tN:�`..�*�F��p�[dq����r����@���q���b�p��5�]庠v���)��GDK�B�����/��4j1�]'��%���z�*W2�^�Lv�������6��;;7f;�M�K��B�a��T��j���ܘE�J��p�x^��h`3�Ok����ƅ�����œ�Zkо�웄��_f?ū�+���[l�_vI��;!VTڠ�\��Z8-_\O]��C��*U
�ѕ醓�*�D �^N��k5�آx�歸�l��vKni �/�gf.�e�ch�ᡊXř����x�Q��G�)!B���)ꎬp�zs�y+`k���AB�f�;���y�]���ފ���?Z��o����y9Gx�wa�v��Oc8����pߓ��}��q�t�s��ݵb���z�%��<Zc��ԯ=3:�����oC认���XN}�{��*��Wi>���s��0_?�K>8�-+Oe¼�(j�%5���~�(��/��Ր�M���<l�# ���w��><L��;ܪ3r��O��&ɺĊ��]t{�3��>>ɞ��L�W=GԺ��d�_�]��t�`�}�����$��Ԝ��R��ᾬw����S���)\c��3����y�tz�q:������9�r�|��wك������Eu!ə�1�z���������PeSJEdO�`�US��{�bh~���������ވ�x=�=�;d����is�A�rY�t���8�ђp_U��#��p:�+�z"��.�����Ku�;�9<�}�D==�d{_]��K��!N�y���ۿF�S���H`F���q��V>�|�&���>���t�*�:�gsȬ��HMVg�GP���ȃ��p����F��$x��,]��#;�u��D���-���R�����(<}}��gMjmIn.�3W<_������R�Փ܄�� J��k�0t�8��q�\��G���G��@jf��y��Hc�<WL�<��+
��Ւ\��?�2
5�AUL�����Rѷ���|뭳�;g�����9��M�O�(�z�=��'n>���"�s%��RCW��"bJ�4.)���G�y�G���X����R��t��<ō:���3��|d`����Z;�������n�Y5X�$x�'�X������ޜ����޹>UR7��'����f��>���,��C�:��>�K��T��qp�H��#p��2���	�����|����ˍ�\���d䦽=�4�==���No�;!��k0�\�-�������]��>�:MǺ��v]:���zvo��^���/��Ԧs�X<j�p2p;��\2���t�7e��W�Mv��s�ů]�]���wt���?e�¿���99q3�����p]J���0+=���pc8z�&mx���
�}��Uy�uc7��Q��2�S�O��f�>ȱu�7R�J9⊟zO�S�Mylg���`/e GK���r��﫩��%��:n�����QC&ײ�Z���w��Kqu��ׅY����C��O���9���^��RT^��\��1E�Crp��7E4��߆P�Ky�X�eYH���f��Ҝn�^�P�Ý�<7���!(���X����������Q�ޢ�r�ܫ��h��hu'w��t���	�$��7���W��}�5C���"�:_t�G��Ô�!�\��?��H۹�N�Y�@����w޵}#��Χ���FВ��Н_,�uP�ޮ���<^{���DW:��-^��ʸe]m���J���	>�`r�w2����ER��s�ӼG�����"�"Pʓ���Nk�7�S}9M{K�6�UX�`sr������҅(��CpӪ'F��_EG]b]:/ݚz��_ݝq9q�l��,� j��I��}li~qqRjyz�bﮩб�F��c�9��r;�i7���z��q�,�" 5I��մLPWgvTd,����i�ѵ��}��pʎ}���������O{��d��wuh=��K'�q�wcx�پ�ǂ׮�Z�GM*��+�U��6u�1����}�H�< �P�`�1��}EJ�5�����z�G���^:�'���MJ�C9=5�����w&��W&���ޭ�P+�#����~����ƆYۙ=��,n|:|:�a�S��Y���W�>��Q�u�(�ߓ?�N�����MP�`��P8Z^{�un�Vھ�Ck^�A�a��7�0Guv�T���B��B�Z��\M�E�]�����8�F�;^ȞW> �6��[�ڥ̀����ԵWN�%�:QGh�ڪ�_JT�˫2Ҍ�ʅ^���B6㪊G �������3�zx�P=0������Âպ�w���.Z�p:�ss�=}G�.��\���O�:h�
�+�O��Ne�f��9��^��*��(r�w���'��QW�ڭ�+=��9��b9�.��hf��H_�~��<Ne��~;�xQ���{ӗ�6�ѽ�S�f�w�^�\ �n�ؕ��������;�h^�p���ذC�Apv��H��a���Ț�3�5]C���F�e��}�=�t�+���/���q��e�ȟzmOI��]�-JX'����b��s�g�A;ĥ�!Ci�&���8:�K=�2�WA0��k"­9�ޝK���}[��5��+�Y�� �,�*�����s��V)VM�m1� }�d�����G�'��٣���v��Σ�C��1�%�gI*��~"EA�mKo����ɷ^6$ա����pn}��GOw^s��V}ʎ}������@�<X5��x>���*�kX�޹/���]����U����=r��J�u�]T�W�E���ʤ�a�Y"v�ߧʇT�Ҧ[�[�ո����ZD[��Y֯8�Җ:���(�wC�T�����W3\����[]�����C�|\Ã��1�e�6��a$B�-�w-hM��[�2���7�g1I%:�)��t�M��9cۚz=����?���@X�����{�6�
�o���Ni�99X��נn��]�Ìݻ��o�z���Ib���7d��ԅ_�/N����ƍF6�����O�
��\F����9Ӯ|�U�k&������J���&d^�xО+Ʋ1Sӫ�G>�mW;}v��K�v��m���rc�b�2_�������&�E��=0�Y�׫�b�������=0�ٙJ��;�=��x4{�O��\y����������s ���:,�����&Y�f.�<�ȷ�������G�#�.wO�%lh��//����}��q���V���j«���d���򉛹�[��¼�<r��gxU-T;�W"$�㘥�ܥ\Ϊ�I]<7����Pv�;=����W ��왞�(��ܚ�t9@%�d���M���ƭ&"��#�MK��J��;�[¥%<��˝R�֪��TE�5����L���ˉ�=�^���BS����N#��SZ�@�Nl�Y�	T{�}J���U������s:v��,\�����n��e�{���b��`DN���:�2�K���HX�-�ɲ�-�����5�y���Fe{A����eu��ZѺ���G۵��>W��������������0ը�w�hD��Ü��	PC�PL;.���x4e�t`�[��4��	���X��qbS��G�W����Ǘu>+�]Hr��b��K7t���|j�bq3�s�ϵh����yLI�[�#�=�W��O{�ޱ�7��z3�{�v��;����u���,��Oe��Ϧ���I�m���3���"7��﫪�f���&��6>h��}�D=7تF[�=Ls��=�zv����M�� ���P�΃���z�4}�\M�WZG�g8�9�'
y��	@��z=��m�H��׌�t�(�(#J��7:��/Kz��:�l��~������3Q�6�W�5Z=�8Nx���\N���|d\C�,�$5��&J�4.���@S��g���p�z.F�މ��"�q�=���t�q/�j2w{�&ٞ���jٍ���T���:��2�ӕ+q)�z�k2pokw#��U#y��{ç���3q�)��,��C񬓡����m�w��cVw���U�doV�ٗ��v�|��ɸ����_�������.�����X�wٞ>�RhO}�����q]Y�����q)zo�yp��ޟ}���q���1�[��+�k��"�fOP�i��n���{��Y�W��uc:��[�^��a����3RlC:�mhCCd���Ǖ�,�]{���s���C��>^C��wW�����ᮐZ�H��`��ټ�J�����$Y�U�6f��
��n_tRq�>;��?}�g����P},+8�z�b�zN��ܮ���ʟ���Q�'����<�d���w�u����xS3e�������d�w>���W�s�b��)j	G��ۙ�6���t1�9O��_M��nj3lk��+�W+{�'2�PwP'�b��Xx�s�5��};K�gU�.ۂt�ζ��Ͻ��WS���u!�o�힌�KL����(;-ջų��B�3��^��B�^�ΧU��� ߴ�ч�ȼ�}ӹ�×���:�A���le:�<�5`����I��>f�˨�<��l���n��oWa�ݲx��}���v���b��{�Ć�e/i�y�'$��'g�8�t�@JM�q[TQ�j�U�w�}��/J��܂�d���[9{�ٮ(q�׷}���`�N��B�|7(z��}�ԅ���A���Ը?zO!��7w�����W�g\N\W]�(�qAU|d��od�)�n;�t!G�vv��5G/��ʹ49�L>����KI����u���,�Ј��	�c�D?VGTs�^x�F8�k�5g����]�?@i�~J�z�4������@�]F�^�� I�4��@��`GE�:��v�>�%E�ˮ��Ȳ{I��֭8�IGF����i�U��kO%�N�S�VF��޵y
'v1�����eMJC
WG�#0�~P���W���:a��"{�g&����{�蛇+�E�>�_*W?�n-ۨ�?ф���7E�MFe���3��I��{�5��}�C��2����LQ�sS��9�`�͹�e����u/�Q��/MƮێ��Uq�+���^��=�F�	����o�T2��d���>�6�t�u�R�࿩�p�̧�Ҽ�k�ܻ�"��B�B3�|�*�'�1�z)ɸ�O@;�^��{��i�UDL5c+��|3�>�OǯjVV�*c}���m·�O��}������������v���X�W�Vha�̢�9�xC��B��c�cPT�{(��R��Dc� ���w�Ϋ�A�G:���Mӝ�����z��9����U��c�7�u{�kG?x�#�iaə\J�ц����.%u>�3�{=�pkYZ�ٚ�z�2�FY�w��$�ZJ�j6�(�)t q"\Κ��8�,GH�rɡ�s9r�s;Ӥn�5g��r�n��*'�����.1O�踽�N���[�)}�P�s	���W��:�������]��t�e�ێ��>��C0Wo���.k�y�2����y�|t+����P ݜ���7�E�:���6��4RF�bѷ�5ˎ�]��ɇ"����o�s�$�W��͸�;Ք;x��z⯢4������1�3����7Tʻ{T'E[Y%iU7I!u�Q�=�=�z��r��XVe��� �D�?��Jk�	Oc����]���\�V���z�}�g�+��ᣐ�c϶���q��5�c��_3��D���^E��ߣ<�����ֿT���w��6[���y\��Tp���Bp�u��z�����v��|Y3�i�wGc)+�0::�l���F��{ʢ��\��>�G>�la.�Q�	��½�l�f��
���nz���=gg�<@栐j��n ��
a���p�[g�zsOq����v�F���a���Q?���;�w� ��y�IaI?�Q�"b_RqR������Q���:���?z���=�1�^էC�&��rY���\F��%�Y��^��C>�����T���KW��C�Dt����;�1|�Y�q�={��5}e<Y;"-��DZ}����;��F��9˛�힙���ݦ5���'�r.<��L�����]�[ީ�x��"��Bz��m�0�.'�s�_��d?��n뗥�����ܼ�N��������U�;=�46��{#�K�������֒$�2��5�:�ǛCt�v���prn_C��q��K�ǈ��" 1t�y]&�Aʹɮci�͵²��M`7����s �C��vL�8���T<�3���R��Eƴt�$Y:�c!��b|�ƈ��{u�{�7�rg�j..5�a�˧i�v�휮�;�3b폩�v�MnAu����nd�8�h�U��]7y�u9�-90�� Ѯ�jk!{b���������*�uX�m�oa�f���
j���,�q���]Zx+�a��۠���hh�e<YN��ҏ%���}\��ˏ�Q�PswL[�� �PZ.4��葀�x[��z�W�{U�-�cۻ�wNK�Fa��):�I��[�^i�)�mbA��̘�����=O	$��_F�M��YZ�(�ȣ�r;ӹ�;\�\� .���fyLQo���+o��[F��HF�P������'�1��!�Л�J�>�.����0�E;��{���1!������Hݼ��C�Pu�4�E;̮]^5�J7�z�n��>��i-ŮKd��b�)�tY�''�I:�i�髒����o4�0Sy�:��(5\ịsZ��]=���q�"`��9j�M���|EWR��vum7E!+�����wZ_V��s�P�&Պ͗��k;Z]Ҧ�S͗n숝 ��L�Nt-�=d`�0��t�ge�]��t��xSjAe.�n��i��������wV��r�,瘣���Q^�(� ��,\o����"J]Н�JE�.��,a7,Ga,�PӨ���H-e�36�8:�׷9�Y�M���; 57��kt�� ���/���ef��ַZ#�������^Q�A�-lb��}I���Ecu����h�εy�j�7�mD���\^	�f�L]
b�`�Ҷ�:�n��:Rњz�r�Ej�!M��u�9Ҋ�ra$'VQ
Z�%���W��h+p��F�5̆&:�7���(�Z�V�0S�4�0k�}�f�x&v����!X�oS�J;���SW3�s��JCř��Ĳ�Ă��Mqy9�r6	D=�B�Dn�bR%���S���%+��V�b��}��V��D+��`��@�}��2�a�^�/]n�=ӕ'��ʘo]�W_N�vg�37N.��a��Jij�b}�%���os��N�gB��yWWva2�����،ѻ�#ح)]h��TV��;pա�����������#�ݶi��.޺�(���	��S�B��;p���>R��S[�ގ������p@�s:��F��
�q�h��lf�,*�5���J]��8�2SK4P��Y]}Z01����_nO����Q�.�C=�y�T�-�󤫵>J\�������buO5u�6<����n��&���+��pǺ��A��j)j�fON���XO{��4�j=2�\mb����8%J����Mf�"R�Z	������B��j�
H���(u�+X���ib*"h���#Th���4�Q#�C�h/�!R�6Ō�M�	MD4�%DD4��Q�;jhj���؃M�Ek��TQIQG-sj����*�bJ�&�9�j��"f"��&�h
*ִ���PM�j%���(�H�J6�r\QDSTi�AUE5SAED��DS4Us8��gUR[���7-Q5QQ%D5IDDs��"����9�Ert1UT�5TQs�P�QE<�s�"�����sq����(�-��b�*���ADP��1A��1h��&(�J�Y�9�M1Q0�4TQE��U���H�a� �P��Ex�������^s˒��R!볷��=z����O��gHyz�W\��\9��7�,D������<Z���:�l�:��?�ǯ��h<���4l���|sյ�L��yup\�!u��\��E�ق���ͭ�)�4�e+F��6o�(����ngJ'�'���^��4��4^bJ��>1�6|�Y��k�sÝ�޸��b+�3��t�9L��3�_�=G�K��}�,���ђp9��wae_��vυt���(E:Lﾦ�3}�z�^/T鿬�)Y�=@Ζ."�yYYM_�\���쫟&<w���:���u1������C�3�ca�T�Y�N��a���IH���hV���
ڱ=��*gp�;����b��^DgD��v���lv�C��Q,�a�5������`qK��I���t���I]���~;�oh*�M��o��m��M�b��Ei�Yz/����\������GHT��_��
Gw��ES�q7]iC��+Hs��\���ޟS�Y���8龎�WU�s �_(#J$��h6⇽�n!�4���� ����ݴ}�[��:�93�M�wu���u��K5�Hj��%r���x����a�+�-���7f�U�vz��6k2QS��T�������o��g�Q�V[��-�c4E��=�<�x���;��N>O�]��l�U��d����f�
,N{���܍�5a���Ŗ���LԚ|!D㢑-A7�)�F�����G���n~c��D{�+�ǺyY����k�F@���PU�W��z��"����������Q0
p��n����+rj�^�r8[�w"���{����b���}�P����>|ʚ�p����?��z��R�����\f\=:�+��ήM�� ���=��G]��5���^y2�Nt��<OW��-#�.}�r��)�Ƕ�������}@t�����s��&�Փ�;��}b���g׳��Q��Fk��/�t��;���V�v����2;����iy̧Wy鎆�)qy�pU��y���6���#�'.&x~������R��9t�|�&7�*�n��]9ް:ֿG}=O��'7�[S���"��VY9�C��.E�o�uzv@�}�s)�R���T��]�4�X�6%s�p9���Eu!�}��1\Ν�ĥ.E�ݺ7�s;��-��c�I�.��+*��oP������0�Y��N?���/Eu��ze��+�Sf�����5u����gE�pԞF���qFy��p7��?|7���;d�y�ۇ�N2����'�M�Y��(�u�Ͳ�fN��ZVЫ��Kzf2��oEp�w�maX"�����e��ُ���J��2����F����ؘ���w�f��e��FK�ٚe��������+�� `�*kf�ET��SR�f���U���d�:	:Kb*�qS-�N̔s�j�U��}��|3j̴��|F�R�j�|}��6K;{���Dt׸���Yp ՆX�j nP�/]>90�����n:k^S~���Y*��ﻷ�����]�Q>��a��D( j�� t�H������ޮ��Q��[��@����!�}����Nm�܈�g\N�������,�" 5���[=��c�vs.��;�LtN:�7Eqy�9���x��;c��ԉ�G�ɸ���.'�މx#ۇWF�t��V��L�x�\l�?K��7E�ʿ�n��F�j�M�u {�k��������D����-f��k�]��oftS8T�����>��Kӫ���*�)��}l�}
pcq���&Jܐ1t�c(j��29yI��k�>WP�ES��W�e=6�zꏍ��1���
z�{�z;z�Lz1�WI��O@;�^��{��F�%P��Q���Oa�}�n�o�4}.�hޥ5̗�W�˼=	�/F>��>� �G��j�S�q����!�q�;������ƝT��_�wX���Yƛ�J�15Yĕ��'�'H�N��6�m�ED)a� �ݳؕ�j�xuڵr(G�pKZ띧�30f�2�c+�Vmf[q;�r�C�����9}W{��,YhN��t�+��⦯:�f�+u�q�;|8W���4��b� �r�
!�u�>�ur�x�i��?<��enZ���j+𢏞h�\���h��A����Q��9S=Ĭ���J�}�r���w:ж}��T�F=޾yt�Y�u�n��j�I��Pˉ��;P�����p9�F��p3�������IRA�u��*��u-�+��}X�3}�Ƒ���I��]O�-�BR�����K��4�� �=�/M�j�ϫ���y�Ig|[)�����m��,��v��$E��T���j�US��׀^{����l�{|��\v����C���m;q�㵙��YpΒUA�/i^�)W�*h��0�[6LG�R����(����{�W2��*�)	�q�}qށrx����0{�|���+��8*d�/��y\U�r�s���}�Hi7��#qrFiy���Ъ|���	���SQ� ����A��z{Ц)��Se����r���
B�X�����)7��n���q�s$�_*����"e�!WR��������Q�4�� G{���W�w�BvBC��M7A+�>�m暡��i��j���E�joWni��-�$b�� 1+͹�����ڂl�pf4"�cn�j�L�8#t!�;��Zݔ�%��V�b�'\�_Q#���Q3r��Y��C����dnh��ԥ����QɢC�o����L�}3�O{�f�
sl�����30���K��B�������N��Y��}Wf�m�IVX���۽R�U&69��'����z4��'Ћ'hza����Y�鼽|tys����5q�Lm�Wx�}w"�Ϩt�q�j�E
�{� ��w���dSq�Un���W=�O3t�0����J�`�W��'U���f�h)���ڰ�z�j��ب��<U�oз��H�O���l�T;�W#f��8}��ܵ|=ꫴ�.�����������G�s����I��p��1���V���\J8K��\�8�哒�6��L�{��W�=�(����+���5z9ޣ��g�||�X��z��࿪]S���&���cr��q~W7��p*����3��j�7�׬�+��C��QX�:X�j�I��F���G��m{�f�8ή.���z;��S҇k3�0�k�,ݝ$��vt�}U9���TMdy�}�WФ�Oq���<���C���Ή�9��;n;�������h�er�ݡY69�Z��.��^�� �]1���3��JtR�_D��b�'3��Ue�'�:G�nh��{>Y�&{=���־j��F�R_3��+�/�̊�P��6�1+�O.qt5p�r\�6>�����c7�[��r�B �҉��f�"��t7�Y��E��U���Y%��a@�ʣ���Wpx�S{q7-�a���}�m�ްnq�n�̝��h��M{�{���?d�|��H`Xn�W�
Goz�4}�\M�u�\�߼�_D��Z�t�9��Úz��vuH��u[3ndiAQ u��A���{�R���q���D�&�>�U�u�|�z:so�Ι�&���v��ȷ2Y��IX�"bJ�41+/��������F��L�s����Ю�#.W��<��}3�K���_w{�%��Tpf��퉼W[W��F:&�e�/�j�p���G|��_7\OzO��E����e���Q��czn���=��G��*V�a��S9W�p���
:�7�����0����g�v��g9］rGO��|;M�'��Nx�F\�<�	����C���gYrnNk�]��8}q����1�8
�Ѯ�D���XC�3y���_Op=�W����t�v_��Za�}h����X�]�ʚ�1���K���*����7�ٟ8�}�3�X=>j��,wO�~�eP���V��U@l������#��$��n�ER}9^�T(ꇸ�y��fP�X�׳n~�	N�P�Y+��z�k42��9�-�6ʇ6T���㎤�)��$1��#Ռ�V�n�������S��wr%j���u�B�1հ��U��A�� ��|�}���~���Z�8���f޺�"��V�Ne Pw���P�m�_U�U�-��4̞��5�R�lq+�{�ϫ��~��3O�}��+���{��U]�{�<�w��l�&��f3ƌ�B��n����u�y���r/��)�C��C������?R�	�af}Q��T}^���&>���]!�Q�Ft���1��~�oWa�l�/=m�$�ӥ�k��z������k��VZ��5�I�	8�t�BRm
�'��V)N\�@δ����õ��x�Zz3d�z}�'��{���}�^�ވ�f�p@����̫����ޅ���U����*�����oz�9�)8U�g\N\}]v�?��( j�2^�4��.�΋�j�};��K���OkWb>N:�޴4z:������ӸJ���u��p̖Iq�z������Qx���'������V���*����`���zQ<��M�wV��Y48f��nwzk7�l�3�d$n �1/k��z}[���l�m�j�M�wu {X��ܾ�Ê���KHݜ7�aLs��*3� �xmDo)��в�9����K����s��pA΢��݂0���cU����,9\d������w6���*�$����\A�4�0��buVŴ�Q ����/�i�4Zۼ�����L�R^������)�r�_D3XT�>�*ilW�I�kǕħ��5�O�hg'��v�s�1�z���eP�T��U�<����&M�u���e��ޙ5
a�5����R��y\*c��e@�R�]�-��啷������ˍ�'�zc��+�ߺz�������3�zx�C�X����C1���5P�n�S�(w��I�n��.�p�u�я�oKΚ|�+�O��D�"�>b��ͥ�h'5텝0V]��7�`9�[ V{��s=X�.�]/U�������p��nr�3={���9�	����d�>���(��=�a��vEĮ��'>��Ƥ:P:���v������/�3�=�?b�I���C.&_�;0��~�F�\g�l�@v3���CQ����� T�ѕ�Gk�ΔV�Z��+���m��n(g+Gb��D���>�;�ܣiȗ*����۫*�5�Sя�U�f��J;���_��q���ex�7�A���`E����>�=�$� �r1�뭞�w��U�����u1���<w��v'5�c��g!�$�1q�B3�0��΍#I�4J�!�
���_r��k���h��{��	-%��ڸ�D�↕n�v-U�7}c�j��h�SNI��vJu�D��;��K��{hB�C5�h3X�,;|5Ww2���wv�?)h�L��&��7qq�鮭�]g��IE�R^�D�"�99�iT�{M�D��o���s+"9Q¯��Bp�Gu��C�.y���w�JV��R��8z#�@l�WV���y����Wur��y]Ԇ�^�W��0f�[������ڮ��[w�o�*i)�$�su����=�S�&<�RDt��1^3��u�Y��f���V|�����d��*���� ��+�R���@�|I��z�����Bzs�dJ7'����}&�y���,���g"$5L���֪ �;�W�K��@����k_]W�M]�]�[��WT���+�1��+�������Ej��&}œ���i��.W�ȝ��g/�_J1�ko��{\fSp��=�}w"�<��L�t�o�ފ��H��ɩ�{Cޯz�P�I�#]�	�0
�������������}#���U�;9^��UD���s]:q��r~��L�q��A�_i�O	�`g'�7)_:��&k=�{���=�=�'����~�w��9ԃ��/aɤjƯ����G���V���W��&\����r�C�['��C����ٜ�R�[j�=�ao3r/r�n<i�
�+=t	��
x%͡Q��]r�9[��]f�O`5x9�z��)Ej"l�(� �9��L��-uh�K��g��Cc��0U��{��=��Q���r��f�ϧUI�Q��'PV�=k��D���Et�+���5z9ޣ��g|�N��=P&t+��8���X݃�W��W-��gˇ�z#fP3�5I���e{�j�7��z�^/T鿬�)Y�=~�=%GMH�TdZ]�Q��T��/�2֙���3�����(��z+�^sX�[^�do/{OO	��ONf{0m���I�D�3_u��g����b_����~�x3��>q�Gm�[��{cƷ��w#��~-U�`���GL�t�����!В�j� �v[ۉ-�x�.��ueD�e��5jG��ԭ�G��5�#����]|��jKCu���M����Mkl�W������6qÿt|M��{�Nq��#.����2* Ҳ"d��7Z����A�\��9�1{�+��ox�M���m!��]m���e���7�w\N�Uq��9�ʒCQ�G>;.z�O��㲪n3w�*hN���t�v�Yq��ǺyY�莙�%��F@��u����Q�z3pG��y�}x+��]������֧��9��P�̘�����CN#y	����������E������E��5 DW�"��E����� "+������ ��E~ ����"���@@DW�A_���� "+����
�2��+��H��������>�������� tX�  �    P     ���=R(J$����TUA*%�1 %D�  $�j�DJ
���JIJ�QT]!A@�����c�ĥ٨�"��"U	A5*�eR��Rm�T8 \����  ̀  M�  " ��$(��`���QJJ2t��J5��t��v�iDm�#0[5*����J�.j��:���m͈뻧:��v�l̻u�f��n����u�wn�IME�s�-72�e��mӤ��1���؛8��[t���i��컫���w5v����pqH�4���i���m�;��v�ӕ��u2���r]�Ⱥ鶣�n�jWu;6�K��jP�SZַT!%
��*�m��;�gv�����;���ݺ�Dv4�n�j5���ZT��U�v�\�UT��$�6�T�B�T�M@� ��$�UIeHD�J�� [� H��M���J$��U$$�03R��B6���		�� W3 ����{�!QE $  � �0�*T ɀbi��0 E=��)*��       P��f��T�   �S�F�)EA�F&��@d1A�4RDh4i��Q�4���OH$�@$�A	���0 @`�0�l4��ZFT�Z4��i^@GAS�q<$����Q,�0�A":D�	.F*~��8�	;{��/��:u?��������[w�#-���8$R���&r���P�E�M�$BN*H�!�TR-HYP�B$��n�9���%�D�*gɓ%�l}P��U�R�	$�*�I$�$�I*I$�J�I"���E$IrIbIjI%��K���{�����;�@�Hh q$���I � Hq�!�BM���@��8�!�I'I8���@�$�`IL$�BIĒN0$�$'q��	8��,�qN$ q�'	8��I8� � a$�@0$�@��@8���@��q���8�I�0�q	'$�B@��M*@Ҥ�JJ�4��$�C��C��8���$��!$�$8�q	!Ą @�	��0��	Đ'�iH�� �4"F4H㦍6�$���\�I$�T�I$���E$��I$���I%I$�I%�%�$�$I$�$�I*I$�J�I"���E$���$�IRI$���I$�I%�kRX�IrA$�IRI$�H$��Z�ĒI$�$�)$�J�I$���H�i$�I�\��?�����u�B��W ��11�FP��G%�MSiٜ�MI��2K
(��_�o��_�<��ج�5�S�7�=w��6�-�0,���QK���|޺+�Zx�����v����թb�`�sWj��ysp&0>�Ӏ����(��[��r��$Ü���;h�oV����D]��Jn��IH�����:�0{Oj}Ϣ���ONK�0'����L��BwY��:o^�M�[tV���s�ǁ���n��~ɔ�у�`_�X;��ު�fq��������:�N�;̓;-��GJZA��v�Yr�I�wM�1u����l�.��j�빢���Ǵ�����8��9n22��wb� h���5���a:7�_-�怴wqײ9;���o;LƋuF�b��P;�9`NKg3ئF�� Ӆ�ի�!��$ܮ���n�ظ�`���bP���7��d�Tr�]7Ļ��J�WL����×uXN�kY�.�j�1rǚc%>�:�״��X��2]���dNǯ3@�vQ�nN�|P�ޯ`��ƕ�ˌ�Kn\C�N8eoe;�Lp�;-�vk�tʶ�*�/Y��2����70�)��fs�Zǝs���Ed��KǼ�	����6h�G�.ֺK��[����N� wocz�}�A��Ҁ��Xi��^��'�<+8��n��:��u�&ֺ�]��%n2�94*��*���|�4�9=R3�fއf�V�ҍ������˒I+��T�d'7Y<��G�r�w�WY|���#�"ػ7��|MZ]�"P�6K7iνራ��Xr-���H�m���1ĩ\%z�9�7�*Z��#����w;��@q_8Ƽ��{p���4����t�pot�AMu��3u̸FÇ�PV��źnjY�I�td��2��M�_[�s�D��k��Å��`�\��r\�t8��w��Yٯ��tJ�"�t��gq�m��>�3�ܫ*��ƔgnỚ���4Kͯ���nw.?����c�HU�__�[0n!��P�K�BSD墦��n�hY��zZhmd��w�J��;f�یU"=�{�-.<��(��n:�o]-ó�3��:���4���َ�1w�m�%�]�?[�J��Q��N����]�8�a���I��7s��@�7I�s7B�����Լ�o:�tz�ou�h-��vby�A�s���Yǣ	�-.����ymmjb�m.���z�E��9<פ�鯵�dB�גC�ڪ�ѽ�7���y�8q*�j���{YD� ������)�WN�u�D�kc��OLy��u�Ɇ{80y��h)A>8�j��p�mjsRŋv��/n]�����|�q:�>��/������"�G��I��E�#�yV�,#�(�7x	�vo͌:)ΚhXI�·Av�V�b�o���U�R% Xg��ݲ�ܨ��Kd��=ʷ2�x��3�I�t�J������.֨��d�#��8�>2*�(ok��pS�>M��jQ����spi������Ҝ����]�b�xF����is�o(�4���d_I�$��{sY���L2eᆳm�+Fp�!c�����|���h�3q<375^�@@V�Z]��܈ۚ*�XYd���ա�C��	��:�b>/����V�̼O;f�a�Lި|^J׳�"�'��2n1�����"f�n��V�嵬��U�ބ�;�v`�kq�o5Ӗ5�.��3pv�6tD5B9�Sޢ�Q��J�zx�����m^��\͠N�͛$��9�I*'�Nq��0�b���d�S��Y;_M]7pwwW6p�S�ٺ���c���sǫ;*��C����*C��<���`l��v��C#׈�-�H|���������Ө�#�=.<'B�j9�����$��c^Y8] ��e�[?uG{g)L�Y����zp�^@�Տb�0N�`ܦ��!�F�*���=�)�)=�9I���C7�W3� k��FmWb#8cqop�j��׽ѸJE�-oR�6ϒK�ӓ ɛ��:ÿ�_�لm�fK�o@N���ཛྷ�|K3V`�,���W���єO�ܺ�uV	�U��L}ú���:A�7%�;ٵSM�K��j��۝7u�3p�ҁ�d��&���V�E���P���d�Ѧr�p�����]�>O���0���7���ǻF�N���"��`�	�t���&�=ы����փ���p�tx,�����>V� {�`ټ��ɩٹь�v�6.����]�Z�������Q�V��{���*�nwn����6����S<��y��@�M�V�m���8Av�v!
�>λ�b�A�Nh<�q�&���sY�t.�$n.Y�����F���.��Ƹ:`&�4�l�إ*j�}:�sT.%|Ht��saUZ�0�<xn��%���רh�@�7��G�;oa�9�v�]9��Ї�X@�͚i�{���Y�A��t�gA�#^Yy&j �����A�ةˎ������t�;��82�q�g^�ă(P͌qdz���
ŋ�[�]�;�8��/����)��� N��,���݇;��p����jޠn���a	L�˻�7oUK6i�Dq,Z�d����g����[M�c&t\�J���om��4ݯU�l�W�î�QS0.ɺSG���5���b�:2���]]ٹ�t����3��Y	�z�ې�d�ӭgoMe ��0m��c/Q;�Z����t�/�5��������oZz<��3xE7l��p��t�4��Z�T�N�r�ˉa��d������11�jNwʎ��,8X��3����T�Wr܀G�8��p���6R'�*;{�*��@Gf��љj�ȴ��d��߰ >Ń�щT�em������t#�1��3�e<l��A|��q�W}���:PFG�4!�n��aË�V|i!8Cyd��;�Y�>��*���Z�`n��Yp?��މ���ic_}xhUՂ���,�^.��E�9Я�"�8QE��hߞ7p��^?�~'|�>�4�4#��� �-�1��^��>����I�X&o��0�gUl{]g�[�U�f���:��j�4�a��ի�ׄ�TQR󶄯o�upZ�TdG11��`a�9�;�����9krA"ʹ �:%Vཚ���Nw{YP��_Sw�A]��E�n���v�InK��T��𐍹6-�&1�L���N#��g��Pv^�ˎ�ux��?��g������7�D�5G��m8�8�ˌ��$|�v�:-q�ޙ&���i�*Ţ�Ev3�F�����lڳȆ�N��1B�|g8���Fo-]p,�=�O�����Sz"w[��:d=����K�=���L�!��}��L�+��FUY�&�Y-N+�*v�ֵ@+h�%i�0�TW���|L����^W=���V{.�6�ܓ�S_y6��~��&х��MԺ����`K�S�Jkw)�{��י �۶R��[(rc�;Q�Yǖ�2���y}�;��k�7���������s�#���w�5�"p͙�Gj��2V	&����h�۹%�����ݾ{-����F0V�[lJ�3Rܥ,γ�]N�:g ����˩����̊cn!��>#�3H�-�~�{�y�]�	�2�s@�Y�Ʌ�f��&p�f�'��;gz��6S.\�N��1ګ%)��ȹz����[�z��7�G�<V�2=eP������������<q<��^�~�">?C|E'lOޛ�/T��f�Cvzj��扵Qf����[+�gfCI+�n��O�3B��� ���4.���{�>[x���L�ݾ��M�|���
\t���YGZO���}Y���%)(�}W���%&��eq%�Ϻ.��7ت��7��3O�����v���(�,BBZه�Y�KV�r��ؒ�+iٷ#K�cc:�]/��*��*�Hn:OZ��GV�F��V������Rĺ�2tA�^n)Y{F�יѮ��S�E��u�}˽��-��n麈�/2µb�#KnX�6�Bt�ӟr�D��k:k���6j��1>��r��E"{�G�\�s�F���M�FK�V���.Y��z�M��W�NkaW��wٞ;a� W`��[?B�'cI�L����>Z��~�<�]�yh	{�����I0I}��=����N�
�Ǟ �-t>A?<���u f���4)����i�֨]���Z�&��'�L#�|4�@��H�[i�'q���y��"TԻ�B�oK��tЯ�l�&����g��@����F���E�?t�Rj�����iC�ss'NA;�-���D2���g|�̠�L��;���樓v.�9x�I��q�=�q�d�������q�L��U�8󺍕\!)�����jec���V�c|�z�o�*,��E\��\����*O^�b�h鶱��݈�b�]XgB.��k�;X�hS7vQ0��g��]4(m[��Ε��н�9=e�ю����|Y�ҙ+�3�r�ӥN�^7�~���.>qO�Ǧ�th�
������R�}��!@�����DCеG�0�ڶg��n�o��#�z�n3�"h+��Ř0Z��Sʒ\���������X<����#��o�Ǉ�����`�QA�m����A:��B�y�#Y]s�Yu��E�rkZ���z�r�M�R�Ʈ�ɍ�i��Nt:�N0*c2]��Ik�oL�l���hN�eb�!����8��:O��J4*�0�+��
���?�z��-K̘}y١�=2`Y��͝�R^\77#�,�Ь2x�V�<t* vG}���5��2E��	Wy9"�ʵ�[#���9`���򭓵*K�!�↲=w���8`��:���!0b7}�7�Qth��`^�^L��v�o���ʢ蠘��|�=3˥�e!���	{��	�
��N{ �+ԯ:��
��.��]e��{�+E��V�W:nr~�M�'��9������v���uOLl�Y����`^�1q^H\9�����0Xu�أ�B�����}�I}<����y�pm;�Z0b�*L��eܕ�GZ2u޸)�gS��3u�-�	�r´̃Iw%��zxhۨ�u$�c-5V_�!�Vg�{��Y��hR��kl��Uw�[��{ۺ:����&��56���yY'f��ON���#]�Iͮ�h��.�XB������^�m4��?c��EW,�W++J�CN�r��Dr@�˕����뺊vpSbK;�=Rs9Y��1���.�$����Y;����;7�rA�Ǔ}�jP<�<�.��W	Q���캱��A���)�Ľ��ͳyOA�n{�W���4�Z�˫bf�4���ݽ�����ْXrgE��9���s��^�_�3+�f�y,S�NZh�A�K�q\��2Ʈ�r�ͧ
j���Z����j"�0�=�;	�Ƥ�v���vr�S�;��HjB��ؚ�2��G/N]0�g��8�^�<�Ʈ����7;j���?}Ի����[�v�{��S���2�����W8�����a�χ��n�����T��]r�-����н~[�;����Tg���˛Ɇ�x��q�� �h����09��OB��`AS��'�X�ڡ��:l�-.ۻ�ݨ	�!.7*$ʖgSP��ޣ)�lq:��n91�2��q�]�))c���ncn�ufgl�\��]%G(_-Q͓�gBIg<�����&�3���]�IM�sNI$r^QF���r��[BU��q�a�M��Ih��M;a-��n�Ņn:����*m�jI$�90NmIP��:fԎ\� ��I��9$4���#/u8䙳�����;\��2�{J�q�s��{�q��ڜ���I&��go(��6�E&�lJ��S)Hniԛ���jI'D�]�K*J;�zSsDG�IW�1:�K�`+��{�VRWOF�VT�t�aIDgq͒k#KnԱ�������[��G���͠�*���إ9�YFA��6vc�s���-^n4���*�#J����ݸ�Cs�0&��p��3oi����Hjr
�S����h�kkZ%N�͑{��T��.�/��M�g�V�{�ǌ�;��[��̷pc0��	)�*�-�]�jը�$�^\{5��$��6o�j�T�D�M�o5On[\:1ŇD�1��4��������I����)��_&�˶_%.	�����y�=(ͽ��ܗH�@�8�I��;����B���A��~�yy�J����8�q8w=�B����]1����X���
�*��'�m�ǀ�ם�|����s�]eB,����*��8q�G=Sm1���{ �k}�~�^����4��^����ޗ�˳�Z6���^�ମCO��i�;�k5�@v�Jx���)G7�<C����ӳ���{mnu��1��	�'�n�&����`��, M��Mi5%�$�9R@�	$�) �I*) �I=�������eǏ�B9[{�����UvTο��!D/���p�g��j{���1� ���{<Ks��m��Zn�[]Sfݍh�~�n���/��ھ=}BK�8�Zkw&p�k�gPIj��ut,���Go�q�{pU���`�\4u������f��� �2�n�P���>���l�n���<cc��!���s�w�r{x���-���r�b��m�����S�Ū�ޔKv�[�L�7|u��t�Y �XW��v�4n�� &p�p���l�h5Z>�gu�#����̐I$�Ir`I2I$2I�I!�L�I��S�Yy��D��`�ni��R�x�9�s�Q��Mks-Wq�\:6n��vzo+�%�k:�]ы��hD����;�+$�i�z�}�,A�z�5��jK�5FY�ʂ;j�1vtٛ�_D=ё��X��^��
�1�yNRD�S5���J���_��/2��F��rg�h�~+;��Uf53,!qZ|��a��tg�?�b哋��=����Y����^S�Jn:��Ό�̹�%���nKu�E��+n��r�Q��I���ŉJ��nwe�u��Nu]>�ƭ	���V��${� ��I$�$�$�d�t�I�I��2Nه*�W�%;{���Z���9\���|�n��߶�&-՞F9=���KB��,��q��ED�n0��Ŵ�8�⡵��`d=B��Z�#���.����wl3 �iNS7\:G"�֪ù��
5g��|�^ĩN��g���̟J\�FA�������Ab��G�}�Fn�#�XAȺЇ���TB:���-�����ba�z�#V&�Dݥ�
�(}D�I�pA(��e!c���'`��g��:�z�o%3�� ~ ��C�{--���v�y\�V��R}$.L�I�I:I2n�I$��2I$�I�I$>����g��x`KW��pZ�ڦ�?ht��f�w+���+�ӱ���5jVWnLĳ�)���:f�Ň��m$ܢ��c�V�5U��&�4�݆g��%7�Yۻ��L=ؔ�E-w,�ѢUWB���eY]�L`�%��u3l�|ˍ[� �=}��N���b�� Z�>Ub,�{����T������K��J��|�����<�?e��_�'�ܺcg]	��{7l��y��ڄܡ���>� AEd�1�p��=��E
�,��Y�D	�ս��pI$�$�$��tI$�)�I"�I$�G.uX��6!�o�qR���ų��w��9-�g�J`�W�x,rP����i������CZ�l�/#�{�i0��	]�Q�.��N����K�����NMuo%�V�Ԗ%>ɽ���Ǟ>��O�֭|mby�o��\��FCT��_/E����̪�b�x��;p�sz2#y��H�.f��)��0��<qʷL�J�t�	7�K�Ֆz5_��}���ǜ.�3tUv�q�.�.��o+�b˿���1��r>��a�%=i͹G�R�q	ɪ��{xo�b]t�f�wJ�^P�5�I%�$��2I32m�$�G.I$�9rI$�J�+v(<�s۵�Q�o��WrN<��wa�lp�뗐|�[�u��yu�#�A�wyjqN�E���}�'��t�f���+�k�v� �ށ������rpx�l��oȽ�Ux�ަ��%�����2)���v���|��!���y�h�����[�8�e�5�ȡ����س���s6Jr�n�N�4�ksO� LG5��cǎ��U�Yi'j>Q��,���d|��Z��g�_	����l�S�a�x�<��*���纞�pn�\�^����˗�z&W�y\�,܈08Zq����ɇ_j�8�QIʒI$�JI]ݨI$�IBI$�JI$�P�[�2�Z��
d�";f[�;]6���3z�9 [}����/p%�pW �@h��
�ϥfK��aH��e�����&��n�R�/7���"m�,����!:���Nt
���Z0f�9��u���J�/R����祽�&��݋<mC�I���~8z��	@_4�c��fw	��#�c[��5����wen�Q"hxIkOp��*�6���]Nv���Q���P�b̝9�b�x����S�f����W�°����
 �٘�>#/�X�rث��G`;�O<�;J�w���c� �.!&�����ܖs:[��� �i�z��G*I$�IRI��%�$�9.I$��rI$�J�c�]�K;�.�0�Z�Zq��
>52f�����+�׀[q���P��+wo}���= ��>��gt��W����LK�m#�v�n���y��
�ב�����7�Z5�r~�]��.B�,ՏlL�a����ڔ�j� ��}�H�Yo}��Z7�X�)j&.�E��n_���F�7Q1�����ly�n��l����S~ɍ���Rdu��0opPM�6��46��z�mfø�B`�����t�xձ�2���5��u1�Y.�A��kt�K�VR �vd*��d�R5Wc���A�Vm�a%|���㷕qA����Ћ��+�L�jA�γαN^��!�1�uf�;~�����Zun	�6?�qm;�`s�3G(r'��U�����i�5����\����lR��m�&�ܽ�,�}b��2��%v�'N�:�qj��^��4t��3�������DvAÚw���DgQ��	D_;���%��}��<*�H�Ŭ\-�,0v]Awh,��u+5��:o�on���Z핅ҋq@�⛄�:��o�����|�
9���G�wuM�:@]F��W��Qgr���;r!�tԷ]>��ѝ�J!��!O1�\`YX��[�Ds�/7�ֻ�޹�Qz6o�m��I��$db$���	�%t���O�����st�t�c���z�?�i�V�����Ϥ��ش�V��TL�$�i�y\�V�j���j�b�R�E�^#w�qx�a����(d�i.�����){�u,����55Cog̽�MY����ڐhn&0h�&���N��C�8�W2�#u�0���RR��މ��P�����2v^�x���<��zx. p{Q2hws:����{8Xp�5I��o�����ڜ�����)���G�E�9� �X��\B����R����# .r�� �>�|v��};�b�z%�EEY�ž��4��΁Z��0o7�r�HQ�JT ?��%�	�*��[)�1����90�E#��������I̛�$q��2IRH�m�$\ӎ]Ao����*_zg�q�o���$�F)QSSI)N���b���^֝2��R�ꢋ��ӆ�^5��cF�J�U()��j�AIF1��[�b,TXj�D�Um
�-����M �EEE4�����ֵ�lel�]2ZR�UCPv�X��4�*���"˪5w�kZb��i�ҵB�7wk��Ԩ�T5T�j�u�k:TU�J���T�J��
��؋�]���#bR�UY-�(�M�W��9����y1V�Gߎ��	]��Lƙ�l�s.�����1&ڍΪ�q
8|������5K�q^^�]Q�.G��eM=��LM�A�ݙ��{��c��U\Wa�!�>W�*�V��ƞ,����g�LB����aS"��rf��c���6�~:�.���3�y�iJM�5�9��n_,:8�����z���j&cE�H��&��w_�uE�LQ�6!^i�s��fd+-簔3}��Ugq����L'n��yˀ�v�G�c]9��s��X�"YV�p1�lо�@�ޤ��m��k&^9�o\ى��4�uά��q&�{��-�{YƵz.��K��*��z{�5=���ގ}=���2��XR+�Lu�vŝ���I�u��F�'pT��u��|ˠ����5�#��-d@�Y��ϑb��T�i�3��z]<%�n���Ѵ��¾Gog���U}С�
�2֨��
�U����UB:�]�!7fC���U�wH�U֡х���2��X7���˝����wU�)1G��dLa���99�K6;�xM*�t���
R�ʠ�?.�~8�{?*)JX�f,0�^tf���P>V������9f����uq��m:��XܛT�����v��k䩮�Z��gr�.Ìr/�������с�$oF�ؼ��	�n�l~�#%ȋ
�'����-s����7��޴r������OZ��e��i���*���v{E�l� ق�-��H//�I����;��Z�;��p�	��)���7��t^UC�}�!3H��q<�ԏ#�"�Q���q�u�������RD\V3��լ�CsNw��&����� ��sQq@˻e��'A���T���`�������
���bvB˸��ގ��O�b�tN��������ee�vf�_Vgb�Y���k��m\q�/��.�9٘���̢��u/��x/�r1Tkѹ�����X�G�b{�PAn�����J�Ƶ�?����c/���t:�z�g�ӑ�h�?^k_v�{Y��԰2����!�Yfe��L/{�R����i����]�l�*P�r)w�͑g��s��:Ĉ������qnm�{0hΦ�	�x���ۑ�������2��F_vm�XCL--�+�ab����^GJ{�q������=�(5�7���'J}�%�R0j���hޛ�&�':���`��1�@�Wq�ˡ6Ղ�~�7��|��Ɇ�H�<�9[|Rq��kά�4ˡ��{�|cm�N�,L���y�*K��i�Z���s[��&c�Kߍ-6�}�@&G
}�VY�`g1i����ԍ��\��Ŷ���"V�$�e�s�j�����	j"�sy��	����Ղ��Wԫ;-����9��G�1����'Ԭ�]�.Q�7[�=C�K�U�fG[�5�C���-�s�;�|,ҍՑ�/tk$p;;��G=�Xx�39��q��ۃ��Rz1�����X����gT�仩�6��2��&��`�#lHo�X�^-7zE��ո�5�i�̝aSUl�v�#��u���[%�����A�E^%ٙVi#���W	�n��I��}��y�d3�'�R|ݘ�Q�-^r��e����I�и\ֹ A��-x��t�K��ĤT��m�.�:����u�L��Qv;��I�[�����+�0���)VUA3��I�����{/&�o��Sӕwx��޲�|4�9욃O��)D�WF�ğh�j3\u:��z���8C��n��k��/@��\%�7'�R�~w�uxE�l�u��� �C޾���E��W'��m(�ڐ�ܜ�f��M�11R��S�+i��������k*�Zmd)�����C}�����|׫R�싙�ߏ&#w+�>%l�ky�ٽfi7�h31���B�{?m�U����58���r+�7���0�,r��{E<v얙�N��r>����/�H#�U�n^�qw�,��]o��i�]o�*�?��u0�f�G�y0���Gv.4�뎃��m�O���&�{{���,��ss�PAh�5^Z����uh'�@�|�{���O������Q�n�)Q��s-G,��qn���k�,�J���{q{zV���\6�)G�}s�/����&W�i���k��o�����y�ّ�C_�&���O�Vվ��QP�Q|r�KZSbʔ�Ot-~���Ψ�a&[�X`2�N�1��T� �.���4
|��ub@�1Pxؙ�[�LL�+��f�>:����F��{"���Tiaw�~�(Ŭ2-ݳ��߷�3�s*�B�yB%Vxvr^���7+��hX\��!:��;Ά�c�J�V��
 DN�l�D�m+&�����q��$N>�t�� �i�N�,uB�VL꧉�sgl��� ���m�$��iΉQR�iY�2�7�ѣI��֠h�|�hI��d~c��AΣ�Bo��04˻:�(���*�n�NC��i����<]J���:h�Y�fG]˽�3yܱ��{4������������U�1��b~�7��q�;]�z*jt�^a������Z�Ϸ=Z�S���{�����vI跲w���W%�4&�\Ky�C&R�]�T������JsD2�3�`���֗s��4h��׾���w
����c��c|n�b��M�î�>�2)p�Z'��8��*�^��"{�dߦ����O��x��ڍ=.�x_����[�����o�9��h�Ƴ�`FY�9�j�V�i��N$�Ar�ܝۧ��D�} D��y*�`#P����+o�]�U2o�����37��f]
���UxC��\�o
yɎM�/�E������{��:��'#y�y����Y�����G�~��#���NWt �;�X�c��57���8ʬ�o�ye�M�!f4�#�_�累�:�]Օ��0�=��*���+��D����Ӻ<s�w���\[�G�Α�zL�寖��3��m����4#*�wq���ݼ;�c�쩮����`'Lpaɵ-0N�Y�n�+�%��˼�q�2�*ǰ��=- wvycX#+O�AwL�N��Ǿ�kܬN깯v�y��(1�A�s�:��e�;t\x��8�#T�\Gs��8�x��gkv҈Ť�Q̝�q�c1�RH�m�$D���)�n;֩G,K;��|]]��X�b�R�X�j����gZ��µ�.R���SUMUU�x�Ҕ�B�T-	)�Q��*��Z΁R)U�LX���ֵ�D�RȢ**�SEt[KtP��ZΑT�`:h�R���%ֵ��Y
����*U4R
"kZ�u��V���(�)�[L��Jn����M�u��TT�j�����.���*�)h-*���,R�0��Q*�.�m
*���!Y�7�}��լ��3�f�/U{	M>��M�/���=_P�E%�ڒkS#���6j��RUl-�+.�>�j���W�ь;g����H=�5NTG��V��<in��=��g���oG;��^�p�.�-�O���ҽy�s�&y�K�w�pf��_Ӫ�m���wQw�
}�G��ۮ/c�T%�p;��7�����H&io��j��"Y�������w���׍{�Ѩ.���j��k$*х��=����K�-�d��VU����v���9����K��1t��V��&�ȸ�U�����I;:���}�&d��q����Y�<LŘ� ����RHM�ި�;����|r4-�ۿ<]*ޜ�=�
�gM1+��ɸږ \Zoz�u�
�n��gw���=9�43��b�>��n�E�<J)ck=}�Γ��U��{V��+33�$����-��t����j�]y$����f�ݳ�V��B��]׬�x��0�=�r3�|G0ߟ�n��;�\)֨�v��-w��j.��zt{TϤQEj��{=��2��o���S��q��o޼��>����7��_����}r��#��N^.�P!5�X�r���	M�UR��^I�hm�[��O�B'����w�=����G7q3���=��n=4�t�T��s^����Ae2�ҋ7��]�"���jV/Nx���O�=+j�<�T����W�a�5�ڡ�7~cJ�p@��8ǋ\���fMw��wUV�d.�a�Y��h������x��+ۦ=���b�W�5�P�C|�÷A�r��qL�<�X
�#�P◧8%/a�$��p�k�4=c�V���=��uq�z��P���{p�h`�}����a-��o��֭K9�B�t!U�I�aix"S��ZM�#}ݰ�X�{#�Y��~C�>E>�J(瓺�������x;�������]r>��\2�M���> �[t}/Z��8���N�
b�q�\�5����t:�@�I��
B`z�hLr��tABW�m�q��!�O���Z~��� a����Bm�0$�ʀ�� i ��l�@�L�Ǫ@���>d5� S��k~�3]���@�I�h���� d٪-�RM�C�4��M0l��[����c}��Ͻ��C�C�V�@�1�� ��L����a8�Y:ɞ�!]�-�q�I-!�6�a��*�ｌ��x���C�'Rc�)�&R�>I� ���>e����Y6�8ͰRB������ϸIi0�$��I
gĤ,�Y9I0î��P�,�H(K;P2�m�l�d��3ߏ�6;7;|v���ha��X���
á�Վ�n���M���h{=�J�[@�V`ÇWܢtA'
EvO�Gѳ u��Hf������0��L$!��m!�i:�ֱ�`�o���2ɔ�� |��)�$�!hq	���=@J/v2d�;A>d2�m'�o��<�=���<�ޣI��I8�d�I��-�,�Bi�����J��I�>`RC���_���_{_|N$�Of�aā�fЇ�% su&P�C�i$���$�'��}�l�}�5���Oz����̆qP�&�>a�u�8�+t�M!�yDm ([�f��k}���!�I���Kd�qtd�Hy�e m��d�$�� u�,8����|ֽx��Bu2d�!��Oz��]P:�(q�l����XI���&�8=��~�k���%�P<v��$��B�lI�!'�Cl�I�'��Y����o\s��5�}����f�L]@:�Pu�yz��2m����
I���"�)�[��V}��;��[ �$�������B�K�Hq�a�d�S$�L4�ZI�M%0������p?o����?��1����#�tJ�,V��U��
�����H.RY��(�e��ʫ2�y*7��{��~HC���� y��:�>��l!|�(u��8�u&�.�_(�i��J��w�m�I�H{U0���	����L8�g�$>Hy$�(���-��=����Ә�z��^�z��@W�'���6�u!�u��@���D�$��Q�y��ý�W��5�!�<�:������i���&�&3�8�=Be'
d7�$�$�$1^���sw��ŰC�[$�d�N2u$4�O�ߒ!�f�i��
Hd�2�����=�;��!�;ʐ0���!���|��N�0���IL���I6��Zq�Y�~�}���0���N!�j�m'�c�H�<�r����B�I-!Z�i �	�|������/���S;�C̒��ԁ�C��HC�h���j��8�|��I������p�_{��>O�L��%0) �g���M��	�y�BM0����a�K��g׌oܒi�L2d��	�4�ȜB%�Bl�Ci�T�P:�3Rd��B�柱�`���h~�r��f��*���79��'Փ�֎��[}�0]c��JR�4�&��ٙڌ�%M{��,�x�
N9?�>��c�;�-�q �%��$�RI2��O�O��)4��Il�Pq |�6�oe�sǹ��i���L$�RO�O3��I��!-�C��'EBO�,�l�o;�s�o��aiRB��m$�:�6��ϕ��h2x��C�$�d��y��^��w4{�u�v�� WZ2d��-�a��I
����nt�OT��W=k��QGo�
��"��d�Do]P*7զjDHg�Xs�����g3��eBߋ�3�͜�Eѓ��B6�%
��E>�LT�ۙ3�,<h
��5K��p&}eM����7Y��uz"������]����77��E��3(�����jvfpvxb�)����:Wg�����7W���L�n��a��m�Ϥˊ��IC��4��w���w�aj�j��%�[ѼlѲ���W==���X'Ӟ���j��n�]uT�B�V�;��s3��h�����ؼJy��gT�n��6���n�)�$���>���<'�ސuo��1dS[��jhWc�C��
�`�$l:e�8\Cw���D�\���V�Dϼ<kn�v���ELgs�e\��u��@k-�a��z]!i��ك�S��
�X<,(~\�P�=cP��2zx��Ѵ�]0cV��x��gzh�$)�A,��X}.����\�շ���D�ndLb�$zV4�+qKx0#�%t��	�X�����/��~�X���[��J��XI��Z���m�l�������Q���� o�A�	U�`mw�R��(,�v�!Ǵ	��ڥN��瘰^J�c�����,�`\�)�ܔ{T^}���%\���޻�+�u�qEq���n�Gs��a�\�q&f����`����<ܻ۠������i���If/wJk�i�������鮓{�����
q)'葙����=:�϶	ܵ����XV �o|J��L��k�MO�\���X�\��d��t���.{�eu�*L�;�8�����]I��_�J���(�G0�o�"�s�H��ֳ�S�w9LD!�f;�r��g[����\0����>=&�ƸxW�w=�zF��蕏*�+(WF��x�|�5q��ӂ�%�K���$�~�|��sx�X��5Nk�����$*RG�D�F����_C%�sC�qU��0K�cWI޺�i��7��u��z�9�ט�F:�/xˏ�w6��q糖u��}��鳽��'���������ĝ�/�ޑ��f��](Ůky�L���=3��v1Q+�,�o:�C)\�~�ɔ���>�en)�>==5D1��|�ʗ�7��ǽ0`�]�4ﴁVt�p� �ݞ���<h�˷�JS{g�p(5��#��Q��� �[�o4��8h��l�v�o_Q븜��#�U��\�~>��{u=	*�����t�h^v���VG�͞��/{�%��<�`�����X��cs&� ��$���b9�g�U�K�3���_��,9YVޣ}rPT�[O�;�Vb�
[t93]�y��y�D���H�<��|8�����؆`:�a���u
�'b�D��hm��!�]��-��_�ĵ���^��Ru2P�o�(H�Ҥ�\�'dN]6���=��ˣ,fa݂ �Y٘�;��������|���k�n��
}��E�a��Oz{Ƿ�=%�Tsf�snSj���ٳ �ӆI��J���zm�nS���\�� ��FT�٢q�v���5(�:Nʕ��I��֣�&��8ےH�R9tW��O�Ѯ��W�wY~�����{��StU ����
b"QUEU�_�QÊ��kC2���W���(jҘ��ZU"U%^���E5UJ��i��n�WP��ѵ�kYҭ&�U5E5��Q�8Qaa8�("��ٺs� ��,�A8I#�ĉ!")�ֵ�i�*���"�������Q�Zִ,UQX�R�*��)��dTF��P��u� �TUU2�J�wv�5MS*�A-�5�g@#�����b�����EQCÆ�m����8Z�Q�)�ST�lU~�����H�E�l����/Ö��A�򸤏_5d�JPzUkq\���q�t�\�p��~��u��6&��w�4�왗�;㍜Ӧ�ե�)z3||w�MՄy�t���hx����a�$�I6��9���Z���ș�А�?Uj�{+z],.�����ȁ��0���GT�{/P���L\�`J�*ꡣ{��8�kK�U��f3����$tQ ��M�����,���£�����Q8rn����Ey�h&{�i~��[��1{��v�6�N]�S	*V�+e�������)Yp�?[hԕ�Bkw�F�f;�(���W�������c��:�V�K�5�j,�NC�\�ۊ�22v��_ �*� ���.����~��Fk*�����M��sD�7i�N�F����2����}?K[�����Tb�z��}7TwIC阯zo� �U�L��S+�����H�G2���i9��&�qu\��L�u�5\��XN[.rj�VX
	�s�OZ�(LvTw����2��*�-g���@��c���]��Y�Nk���y�,�붌����zu���f�P�V-��+�0�H��9+g:oo�0�R��[s���Z�b��{��|_�����g��f����G�4�����<�k|K02����=�F���|�䱹��,�G++ ��t�I\���۟Ϛӳ����Q����8F���8�Y��]�Qq�y�PV�q貆i�u/��^���
�y��AW]v��n5��w�NE���Si�՛S���t��`�G=��n������~�2��L�:��fn�ߓ�����
��՛���	X��s��Oy�J�a��G3g���kUf�E�Gn��;�v��s��;��"(,
)�i���;�_�����;�,�Ѣí1dnk��]�	��d��Ǣ��i������Q�Q[�S���G��/���#�����Ef�Z���I%zm�Ӈr�� ���Y?U���]0�(�1\Yd4HR�i�iiv�EÙ���w�s|994�z��.x7aVufi�KnM�y)��T�Y�Ci����/����,��W��y���:�bw�ѳ>�4E�v��n��CNn��5:n����=r�������},8��$��3�\c�o����O����X�(,��d,�۷?�26�;,��[ �*� ��l�gq�0z�T*��3s�jy���]>���~��Q�Q��zV/��y�r����)�]�SS���u�f�����̪l�/_�M�iߌ�^��o�;�	����Q�훅f��N�C�|q�v�#~Q<�)۳L��aT-��#�>[���[}�/���2^ϳ�+,����|A9eV����nD�9�H�p#���Y��j���J�EA�nwE-s��N�|!������o��z��x�5����~d$RE�E�N{����[�kߣZ�����)�h�Aj���
��y�y���,�?[��g�߽�7��)�v4�]�8���l5�yn&U>�}
�t֐���Й��gق+�~�Ѭ�gG�������A�s��R�M�7�#��~j�;f�J��`U�ݹ�<�=���#�Q}v|R���<���Vpu��Y1C���Eu���kA��{��8"���|Y��2s޿M����3Y�#W-�����*������`ݍ����ܸL�yad�ȴ���h��IgMh��s���,"�R)@P�@��}�>��{������o�"ع0�"�\�b� ��;�#=Wf
.yI��?|���\៊�6/�&�U��!��U<�=�]�,�g9��L�Nː���)�;������+k�RH1ݟ�S�Գ��ﺕ熭���"Q'v(L�ۉ�q����V6,�F�#OM:ͦ��������Y�Pz�Ȅ:QZ��_hNt^�^���Ԩ�ʽݘe7���zT��[�4e�.���9�^�jy��@r[k�Hd=�.뙳޻O1��v��k������E$PH�E��HMw��Ҿ�Ͽ�F��#[��:3[g�p����{�w��t,��w.:nu����u��j����[�:kI�J�����V{����CR^����$f��oWv�\�RB�I�FDp�wy�R5v�v�]�N�X����Mp2קFXG��M���d��D�u_d�v�uv�ΰ�m�$�Z%��cke��k�̕m�ϸ����4g��x$^E�Z�h;�NeM�s�a�h��u�I͹3��ε��=�Bك< �����TD�m��Q������d"��d"�E$����O#������Q6v�#lB�ed!Q(ۮ�w6��e���D�5�=�u�m��R��t��R�!��w3+8�	j���WA�"be�}��s��a�/�k$�k�..�6��� ��`���������^j��ǅx�ڲ:Oq&r�=�׵�4llK��]X�m��{jȵ���GI���8x��{<�ɏ��0��4�PX�*��h��̙���yݑ��-��������h�I;g��m滹�䁍7/bm��p*=�;��������H�E�	@g菦~���m�=G�|ok�z�>]�W�ʱ�(�[`��{�5�&J��qո��%a�1G]#z'~ܢ�z�W/�V5��s_�0���O?[M,���IdΧt4��p�5�{Rxy�+�E��}Y9N+m�~��Y���P���I�%�=DOn9����}�O����L� �&7�1V�9yMU�eŇ���G���ۺyPG��[�g8��t
��=���9�~���ߐ�ǰ������z�U��k�W-v����+;ӷRor��S#5�6�v�üONrM#=�����'�z���R�U�/�,����#�-�QɞE�{�hhr�X���v��~i��\�f�Wb$g��;��f"�
۝��O+����k%ȍ��2�.sGK�JŬ���>-gY$[%i߳ض��p����;D:�̇���D%�6�y��Jx�W�VҬ�|e2�jV�d�	���y��=�i�Ǿ�!���b�6���-�� {Q$�;�x3:�se��L�SY~UnE���&vٞx��Tg �����@*��0���矷�	�=bퟳ��ݹ"�]�{���M͗]u�[��Q>�A=���L;��h~����wwi�j)a~��,3����q�R���	c9��zrҸi�LA�5%����1`���s�]�s�:�>F�����x�������9G��f�R��zC����3�٫K�R���\u?#�I��J��ü�����8�I�y���H[9Xț��ڥGoSy�pm��W�vf�4҃���A�ԱC4ǳS��F��+���@��6nţ;&q&��u,ԙ�L�R	��n��7$���G�H� �Jn��i���)��߿W��_�w���`ȫM���������R��]kX�R���	m��TP����\a�u�"�*,�U��+��-R��[mm�kZѪ�����j�R�Nq"p��0	' 8�ٹ�`�!8' B$�3$�l�i
�WB�(���EJiKcx��:Fy���4�
��kuH���q��Z��ݖ�u)�IIUKTR�4�U(ƨZF&��z�5�m��B��1��M��`� �)Db���
�U��]���������Q;��ܮԨ�Nv�m��fٮm�ab�����UW���@�$�H)$XH�I ��߽�����G�=��O<v�%w�΁�#�^vk�X#L�VJ��ѪL_Z�����@��2�G�8Be��,.�ԘVvm�8ƙ���AfxEF��<z��5��R�������ۘ��ۊ��Ά����5�#
��;KD_�5=M�}��S�����ȣ�Ȳ�`�C�������lKpm��A,)N**'��^_��_����׸+�7�=R<��Tc=�4��g�����l�{�Z��mJ@�m(3��J��kYjs����)$P �"���"���?}Da^��s��Nz��Q�3���z#yܻ|D ��&����Pfݽ/�/K�����0����>�@KĮ�.�];ЁR1����Z.�G&EX�u�������%m�74���3;>��;]�nH�='1�\`Nŭ��s�ꋠ��DUn�4��W��k��<&���lz�����(s����[���4�h>��)|��q���8��QހNF�d�o�\G�c�bL$�yj=�ƨS���s����8]mc���ߏ5��ud�(G8�FUfv�:���r	~�>����}3�,�d"����\�?O?ѧ�j�t{�^[��0#�\�M6�0�X�s��Y7�̄U�ֹAl��7۞�~������x�97����'��|�{�
$���N8o�dI��j�]qC��ӧJ~΋��h��Up9���=�����g�o�&������N�([��l�˝̅�y2��B캚�it�ccǫ"~;�lM�o'r�ӭ�c�G4cD뜸�7cz����6zc�{��Щ8D����E��!#�0Z�|���Xi�C���o�����@���a"�� ,�Xd��I9�{����r��~ƍv�_�@�W�#3O��6���']�ț��Ԇ��X��C�}ef����'��Z*+������VL��7і)�xwo���0�j9��+T"�J|>T�W� ������[G�ޟVm���8�9���8��%^��PIxС ���`MO�
�.���s�$�g6[��(|<?Z�_��S������:�N��ьgZ�%p��F����c���G��)����c?)�C(��p��0�c���8�Jxb$f���8�Q��oVJ�k �����w�ޫ<5��[�;���!�  )( ��d"� �}�{�a?n��M�Y�O]�m�{r���i����%Ub�mZb�Ѹ�P���w�����D�E>�U�ʩu.U�hS�/��*�o�l�f6��u�
7�l����F	���U�]9Lt��_�xB��+����˯1]�R�6
ںPWL������e9�}U��=����V~_�ƫ�u����u���"���c���>��Hf�Fg��/*"�mS�������)����j���sy�����*k��������˚M���]�oZ�s&�P�R�t0tu,�c���K>�@�,�j�'ָC�᧢��2�z�'4�o!S�e*��լ>��[��rz�Ef|�(�ܡ̖������!�
HE���!~��{��vi�翌Y���x�Kw������Q�I��K��NS�W���0/��Y���
9����`�D�{.0ē*���;ʠ���f�Ի���	�$m	�u+���بs��y��.�}w�>��x���0T�E
�1
?�p���8x��X��d�����N����\�{C�/���o�p�ߵ��`�����O���z���S.��)�cq��.+��}=B�Y�yW,B��
�%֡w��$R����u*�m;폛0u�/+t}׷YOs׼)@������{�~;q�Gܨm�L�}F_<�oFgh��8��e���zQ)"���R�к�Y<��iN:������[ڛ�F�Ls��1��yKö���sZ���󿤁��
@H(IH)^u\��}���s����ml��D�&~��02�bdC�Twv�*�E�<�R�.uTr�(+��B&,T\�m��Ǜ��+��i��_:�V�>�ح:L6�;o������ ��x~g�t����������ӗ/3 �hgТ@��JnzM��=q�.���ߦ�3��SK������Y0�GM��*VܴI9$"�F,��{����Uf�D��a���1��Z�o�7\p�>�7�7�}�;M8��oc�;.��o<ؔ�7y��|]m�;S�;T�|��(׽���f�ͼT:�R�6k�K��t�~HW��+�w+{D]gN�!W��fEz0�}WN���&���.�fۚ]jj�BP��׮c�w�b�{��G[���w��,�Y"��P��s��}7����]%�U�Q*��y��㚣O��u�sW6���[ݞ�M3�Ui9W���.��_s~�w�n&�=��Sw�`�:�m��fsVɣ~wƢf�B�3�q�
�����W^fz��A�2��@����[���f
�n;WJ�Ң����-�+�pX�x����'��5���Ƹ#���K�u��r�
-xo��Պ��)����BǸ�`8���7������rw��p�V���TF��V�t��Ǥ{V)��G*�W��x�[��G�GS�td'Fh��,9�t�U�Ʒ;�M�}��AP�=�q�.�K�С��L�S�����R@��#(#a@�U
��⫔����i��������H�E$Xa"�� J�^w�������y{j��^[�YM��x�+VR,X��ޕ;?����C�z�����;?~�n���w~�5����)�
��X��
����Y����-ۼ��ZQ>�s�+���(���% r0g�)R��'��K|"j{q�+��>�wJ�͹W�$lT�=���1�����5c�mJ������O$��c�DG޾�L�+�����5^>��;ƫ��32��\6y��;b�3�q�uڼc�纺��"D�5Ja۸�{�?l3u�A�^h��a�`�ٮN�!0U_��Y��+������P�Z�3~!��*$���U�k�[��mS��Ms�W5n��S���m2����-Bt�����s��O�Ad"�,���
(w�{�}�X�����c�c�Rm��/-�L�3��a�CS`�f4UM���-֛�Z7�,|֨P�<^w��+=j��w�oޥ�t|%��n�=���"��Ə߼G�_@��&~�N�*������Qf�`�Gm�'nT��:�y�"'�1�Zi�b�-��ћ������MK�K��`*�繟E�5�UTe�����gn��Ӗ��Kw���
>���S[��|��ΨZ�Mz�u��m4�ꑁ���љU�8��2$�z����M;wN��w��NR�̟����t+.�ju�;[|Ӵ�]���	 �7�i�Pf�t8S��$،���:,����V��f(3�./6�o�����]**�ܩb����K�|���T�򹪄�;dY���h���6�).�6��a/ "�������9��.����X�D�Y��%��
�>�r�Up�5>�m#:��OB���>NgW���4r�Y]+*�ro\�wveѩG�=�۟�U�*=�Jml�m\'W�jw���|����ރSy�՜kh���S��qk�y��Z���4o�9,��.̔e����a��.��ٕ�hml9��|�OZ�v�]`u{��՝זx�?mxó��Mj��%�*���F�fy役͑�/������)g��p��	���=�њ>����ȴ���ݙ���BrA��6V<��ȕ�6A�,���M�?[�G��'$����'ʎ��C�=�m�XHe[�Vnd̝>6���z��"yl�r�YY��[�e6�oӵ��W�R��M~6�7���'D�uA]!趓����4Լ��[�����mL_q6���v�>xx��N	�upF���rv��?3|�m��s}.��\�{y��U^��{�?m�U8m���^cFp�ئs׫��,�����;oM�P0jiw$ʊ�2�H&�J�+��9!nIQ�$S�q��s"@>��r&Rȴ�~#��X�
��UQKL��(��q�P��Ѭل��ԡST�R8�S&1��Z�.i)�i
1Xŗq��U�R`���Lb��s�T˫��.j��cXH����[_0�`g���Z�A���E4�4��[K�ֳ�kVV�L[�YiQ��
�E�l�h���
^gԻ�-�Қ�*��AŅ%�j��3���"�J0�Cz�&)�A��l�JB�˫Ín��@#�	��$�y�$�%�� _�@
%�?<d��>!�$��mkQb�%��Ĕᱱ�.>c�D} �'����_�|��7��Z�K�1N3u��[9�u�ќ�J޵�s���I ��B
3��������z�����ƭ�u:�󼞺�2�~wW�H�ٚv\�d�񮙘�y���v��1�N����-d�?3FX`����9�����w~绖�YM<z��>�y�ĦyR�_WO�ӡ{��:k'z�a\͜��`���Ms����7��)�%w1��m�u9��J�ЯdϕE�G�SR�g���ʭ��vy���f��g�_u{v��0�|���᠊(C4���^e@�/�0�^޻͖����N�5�'qZc�w��Qu�}ʍ�ܛ���yϯg��Q�דn��0r=k)J�]A��������_!�b{��r�.�lї6�������+����D�	Yǘ����gMl�D�ŭX�q���y���� ��(A`
@RE ���}���>s�۬T���O��o��n���_�
�nKH���U��\������4jeɔk�BlЙ�M`�z�y�4n�uR�������.�s��WD��
������u�ȹ�#�z��{���R��xeh#�J~n��	�Wf;Z>x+(�^x;8�ޒ�G;x�\�A��b]u�YwF�__Rś۩f�^��:dr3c�.L��>U�j*D��/��͕�����=���[��F�b�u<.f*~��0/�J�[�5lg�iΊ���m���[��j�Y�%��-$�	��_b�5�yƮ�3�1g���;W��<n&Aφ=���3[Vbz4���n�NK���T�KƲ^�Ze팀Y�;y�a�m�z�Ǯ�cLw\��n'?����H) ��) )�	�-���L��9;>ꊓ:!_N~�y*?7�i��q���?.1� �������j��9�4fw(��AN�����9�^�1鎖j6fD��\��1c��{yb��I��
��J�z߬8)|Fp�)���Ϡ�m��|����(�vn���&nD���՞�j��J�b�+w}�䯩OO�"��ed��B�+��|)1Ƒ�8]5��y�J��7�6�]m]4+ �[j�w3h�z�;&Y�����J���>���k]U�G�7�WK"
��B�ݩ�3Ӝ��o����U̇Q��r��]{���:QY��~�f��c\j��5~?��mF'_o�޲�[$���ͼ7Ȩ�6�e;:�Eqs�9K��/u��6o��z��y�o|��� ,�XAd��
I )}��_}�w�.�:g��>��=M4�8V[���HV����hUD�6�d9sf�d|j']��H��,�r��ĺ����1WW�W�^�Fɘ;�����x��v�������p� ����O�?e���w9����b�t���3�a?5eO�㝻�<����d�ί�J�M��\�X��=1;8���_	Q[�n�Գn�V||=}����Ϻ��A��q깏�о4/E��C�tۢW��*��>�Nnceϥ,��191WXF�yJ���H��ʧtXDF����S����P0��]�Vӭ:�p.����Y���4�vj끍�}�`Y�y* Y�X�j�g	r"M��:gfb4�v���o9�;ε���7������ �A@��� {��/}�k�n��Q������j��u<�Yo^��]s����y�����P����)xv�Cҿ��
e�F�oj?�;��kX�ʰ�xv#�(YN{߶2ׯ&)'}F�f���q�>�����8��\3���n���-3����i�4�N�K1GEI�K;w^��1�&���P���{���j��z�]��K�FJ4�ϼ�f�T&"f6n2���>���L���W4�g�����_м�Yu�}�S-`0;�(�ك �4~y�|F�ek�i�Fq'�W*�����^��	�o�W�m9n�T���G��i轊Ƚ�-㹔3y�Aᵾ�Y/���{��H�N����P��#��]=�]9�c]�9�� ��,�YH
XA`$��ｏ�2��\U~LF�=b0V�F���a�(Noh< ��*.c&�\����͚S�&��bOw��ڽʮ��3�ݖ!���4��흲�j����L�B򱹵�Ut;<��4�����UGIqS�����3 H��̽�6A'��?b���5��.Dg���9�jr:���9�җ&T��������.&x*�~���uQWBa��J���������� .,}�Ñ
:����/-��1������~�������
�� ^���fE(�j���/U8�k���[�1�*n��~�Cy��������rGӱ9z�����M���fX��B��:os���7��2 Z�.*<ݽҕ���9�Sj9�_O�$Aa��
B(s��o���UgT~�R�R��Y*&��u|�*����v`�ގ�5
bw�&p�zD�������n+*�[�Ko��ntU�LY˃0n���r&�U�\ͥ.c�0}�XW��^�>z+��~�ݠ	s�<�G���#��Dh����9@�I|�9	u��j�8+隘���[1�ӑ�~����<������!C��u�\B��6�o�W70YSf�2�w�g��Z�&c̌�̬c�j�0�߬ޠ7|_��g(##q����#��v�=�.Ŏ�?���s�i�KW�A\��Ww�R��)ި����t:�z��q��{aϮ�r�W[ZY��V�`�:��Z"��;^��w4�pf`�J<�:9�w�|]o��{��̄P�@B(`E!$9׿{ܵ/���,QS���Q	ъ#/��d�q��~vk�`i�UL�����
��4%ݫ�]�����o�����h�(�<
�㇋	�����ߴ��?Z/��*�z}1�rڷ7*~Q1�|�����빧���{���X�V��ںuc�.�faS��S�2��l*~�U)�Z���~^w�=Y���ߑ�|����� ����b��l�ݱ�J����p�&O�5�
�؛�nhT9T�w�1e��GJ�����t���߫ꉎ��t�����2a����M���m�Tf"gO/�f��a������ciۣɊ|#+w9������fHH�j�	���o�g(��	�˭���m�D�JNO���
P�X�,��g~��z�bTEX��J���`_�߭K�2 �]��g]ݽZ�.r���2�2\���j{��yٜ����� ��3w�FlLQӣ2�8~G�pʌ��?���Q�~���UaYM�u|)\�t�̴W�0��e*�ˢ7^�+,T�%�2���dÞ��~�������g$ʣjvcf��YE���J���#�#�%�zڎ�d�Jn0\[���8�O�T�]A�)R�4<�w��|%"��xN�Eow<͞���f�������v��!v<>��.��'/�>Um�����z�U����p�᯶���~��omz�]M� U�&������(z��TX���2�슦#*$�U"�`�����F����Z�.�z~�{�o~oy���;�o<�7�w����b��X�����{�����~^P������}1S7�R��]���s�R�� �4����˾6�.`OٛHj�D�
&-ҳb�F܃�觗�}�Tɟ�^5�����T��u��U�-����0R�q�ηj^�Oo�%�YYr�ށ'��p�y��c�etv���3�����ݙ�*͋�����H��D�wZ�&q4����8�gC�0��Ոp$�m�n�Yօ���s�VG��´TP�13��|�n�n ���
r�����w��"MvP���.J���^��;�;{WYG�5�_\f������ǽ�jYU�V�@=�O?�c�#�i��
��
5�E�������QҺvX�o�j�<o�8���ƃ�(z���y�]-]���}a�5u�9r�)��c�ג��d���۵WȽQ��rg��4O8�^�G�IӾ�!�8����쫛cwkbé�Y�{�����3�JqH�ᇇ���y7���s���� �˰ep��/5)�o:|e�ek;�Q����k�6v��>���<��>��{��p���M�E%T�w�6�R��_]%��g$k�!kܬ���f\6oD���Y[�.���[�g�TY���n[}�se#������NB0�]� �/>'�o�~��?�RD譩ڳ��Q�:<��;J�Cᎈ��+�U��J��ȵ�*k�{,�|��=Zl�-v���Z��#s�Y��F�Q��d�i����^���Eh��.���SC49��h�53j�Y�0sN��C���S	���&����sCپ^.��_xu5�2�-��W����Y0|r���:;��Y�7������C��ϥ�r�<����2(r�2�C����=ފE�������y�y�R���t�8�֎�0�Q�B��tfY��}��y��RӔ�o�2��r	��(��rIrH�H�>�9sE�\�2�C> �ض����~�U�ة)*��-�ie��iV�񊲓Y���*L��q�`�
�"ᦃh.iUB��ε�b���Tm�(�[�V�8�i!�%�n���A���E0X�ҥbTUukT�B�� p$�M��:�ɡ��8pV.�
�.�a��v�Su*4[UE�طB*ޱ�c:@pҖ䪲�R[cv�ݠ��-(jۖ�Ԥp�
l��A?B� �B#1��_b�UJ�1K�-�eAVT)��3vnC�,@�������p��i}��RX�P�uw@�zγ�4�-�Ք��UV1K��v�U�����E
��V�i��3UT�U�P�U,qv�>�R��y��O}�Î�蘃Zj���5��J�]�w��!�((��őd������r��?ȟ�(�s�n�wpU�1�\�WsD����2�9���2'�Z"��T\�󮋨�h�L�K�z�L���z��9�n��pf��/5-o�}���tGo��	g��(��@�0�-7f��Q�_�ٻ��z%�ur�����8^ey޽���㔯Ŋ0V.=F=[]�õ���u��s�ĩ~�8*�&-�ę�\o��É��K�)�o�]O�v��7fOQi�g��곫Ǻ�@��=�Q��F���A�a�_���H��*`���Q�j;���NpTzjrꮬ�E[?N��D-bX׽�f�I��d�"�ы/����Έڮ��h�0�ab�q�}�2��)�[L�]9��]k}�;��̋b������}���^/�^��Q�ܣ3�w��h��9�J����up�����~�&I�1W�&��Wf�����o����Q�G�	Ƅ��40��,���l��g���>����>B���*Z�ڪ"�~"r��N|�T5@TLÞ�0&gf.�Yu�*Z�<7���++0;W��˧��+�rС� �N�^���;uW���s}���pɜ~?H������yq��=;�;�>yc^O�>�u�:t�}�\�8����x-��~�fm֡W=��&��Zs�~V*�t��|��҇*���� T����S��UA�ܧ���[Dy����Bc^���XgrĹp�����_h���x�&�V+g��V��U��%����;�W�8�������Y"�PX�׵��ǵ�GqZW�i����!G{;�V~��h��F�����k�g��p�!�0:���Z���+/(��K����9y��Þn�FA��`��6�����11�oTw-�YdK�y�L_%��֟f^�eW�r.��*�~S�f{�'d:�qQL�˗06���*S���Xz�+u����>���8+�;��F�|)\��*k�W�������ۥu,���\�B�_��^���>ΧLP�쪗^C�Ջnhۢ&e�W~g�d������Mw�?�a?t���xR	\-\���BraM��3�wը�f���0`�5	��.�7Φ#�/�n�;���l�r8��T��;��sDX�s��f�BV�f�����k��{��(
H��b�;�{��o5�Q��^��J�Z~&G�[�8��J��b�X:�)0���b�����\��8}]O�~�cx��_rTyKF�U�#0P����_�*�-�b��נ�W�G�;k�2�ۧUG�`�y<u4YMě� wF�_�_���\؂���^����fD�����[���~���=�LR�2�~�SM[�����1���W�LA5_U��\�W�
�w_t���u���ñ��]M̪��k��W��Tǯ�_����ޯ^�t�4��7E��>t��iC?g|~�����P8 �?�ќ�6�#jH�����Z5R!u��:U�:w.���5w��S�Vq����:D��J+�7ш�O���֊���o���w�~H�)��@�������ݿ�b������hΊ��V��F�r�j�=�w��g*�����ݳbm�1�(M�LT�Eq��}�H�y7�b�qQ\_hc��Oۯ�#i�~��ƈ�7����e������_WG�Kǀ�3�fn{�B�3��}9*A��Vfg�~2l����K'�d�:> ��@����G~��d��קd�C/+¤�
V��l|�Ǝ\�0�f	�mt�����U���3�;7�;F�<+�@��*&ө�p�GJ����%�qf�`̧�Sʟ�S��S�z���b��>x��*�[���c;�矤tД�:�~̊���A��o�w]���m%�Kt�`�ׅ�dE)̺�q�^�5��������H��Ea����O�A�?:���w[t�ioSi��/��o��ۜ<�|��WR�x�+��/��K���.�v�~����, a�=Z���(�91��XQ�8��N�1���^�]�HP�b��u�	���_Ğ��s"f�f�N�+
]oUu�?TZߕo\�_߶^;�B����.��9g�f�TR�8_��m�g���"�x������;Nv�f�4��*�*~��P�?���P�@�Q5/DٵuM
�o�VX�v��{U�b���F�T����~���������W\�������@�g\g;�V�����@���չ�^ޣ���3b��[Ƙ���r��%X������;+]9�_kZ�y�s��~H����X�)&������~7k�+�*�����(�lL�g6���}���o\�+��Շ�%�p�W�&�?dGS�hʟ��E�`��j��[��v��e�`�:�4�p��G���q����yuZEV���R���c�ej�m�?[Ϡ���t��4DL���qB�Tu��ݼ��>P��~��j���A���#���ѿ�����&����=�1D�'p����	�ܩ�������.2�b�ۜڀ���n!�c���кqv1.>2������Ub{T�;,�5����$�j��s F���M��U1g�
��-vS�����:p���ۮo{_�,� 	p�]Y;ߗ6�yP��n	0#���k�j2[�j|u{^:�O�����U$�������������~x��|�!��3s�Z�5w���K�;��CM;�en^6���{������o]Y�;�3�NFq�(��륈?x;��v�_��G���.d|O,מ\φ@��:[�gr]��*�\��e��ǎ���^��q��Ǘ9�u�6��*�z�l���������>֠�q���5���A���q ��~ҾG�f �u�J����á3ƶTlȠ��Ն(ٷyf���a��{�6}t��x�!��E g�`���?Ou����ڿ�]�^�9K%�&
�r��w���Td�5dC�90hcG�4��޽t��t\Z�ұ���-�M�ü�y���7[����iCt�^�[s������US�2ןw��Ͳ��ou��u�ó�>L]�.�B�ޘ~�n�����FD���g*=ꋓ�;�;f�	c�γ}r����n�Y �P�J�]W!�v"ܝ����}���|~@� b

?,���N]�T��E��C7�q*zb7��Ӿ"+o끐�����w���v��ԭ��ap"b&��P��&�}xP�p�*fe�+��"\��T�pu�{KI�E�-p�qx.����+�����{&�x1��D)�O����9&Ol��L����������nP��^|^VZ�]}ƅn
�&e���Ӊ��Zn�M�
"sc��0)�ltZJx��&�D�I�����l%ˠ�u�c{�9����(,X�X��c������w_��JMHu	�u��4f.\���.�/�-��VR�S1YN_�誀��6iM��T��ډ@���X�S�e����J��/�<��:#[u��~���L>��������jjo�q�S9�q�M��Y��?Iw?	אs�Wbt���+�����V/(?��N���W�=0�	�w
�"�ݚ���*�m{�f��~~L����ii��L�W�퍃k}���j�L�uCQ��."cU��]U�x@q>���U��KwspߧGO�G�#$����;൮�sSQ1����=E��;�_�;�Fy;\$W윎��_L�"HڔB��72�b��2-�Q���]�O^���J��ȁ���o���%�Of�Ȱu�v��Cs�
Q8:]��[{�̬��Ńs��=�:RJ��&̵������+MZ%y�ε���L��wWM=kW�xv,�w:�@�Ь�U�3�V ;�)�@F,A�Y��#Mr+��V.x3^��؈Ԋ,v�<{H��
�Nٞ/Bw�og�hx��%��a~��ຓ��a�@�{�V��ª:�O�rl� �!Xc���n6_9�u��k_.(��WLC�k͑�M�4s4u��/�����4�9�)�B��.Ց���j=S'�e�m:�bE	�FN)�;2� N-L��`acǃ	��Hg���e�2��V�\��6�[p܎��˕3k�Grm�zs�A�қ����g2�7��O�� �x���2�<_gy+�a����9{WO?6�[¶�(:�i�p�ɋ��o4^.�QرyxO0�m;t����p�EF5��|�.���i���z0o2+b���M��	P/|}*�c���V�W�5*�ȗ.�Z��8�^9��Y��6J܉Ë�/�tԆ��y��tl,&��5���ݧ�[3�;A��X���T�#��͓�_�\s7L���\�H��)Ѹ�Z�KІ�W�)ӥ���m�e_Ի��b���R�B��n�	?6NE�1�e��CaG�1���g��2XZ���As4�a�EU40R��S(�V��k֛�ڕWMj�a0��QT�m�ً��R[6n�Չ��a��$Pc���e�Zε��WCwTf���፥��
��f洰�q �pf"~G��[H�,.���ZS4j�r�V�n�[jҭ)���[-��R��gZj4��(n6U�^*T���)QK�����4�0��i]����cԶ�*`Z���n9�_y�0��ӻ&�<��sOs&^9.����:֖��ۃz�u���`  (���}����6���-�N�tc�ɡ7�$NG��%�^�a�w#���2g�9"P��TĚ�HTe4 e����!�<��stzUr�؛j�)�]7��K	E�����8�dd]�5=�p�MʺW��վ����Ռ]��]�;9Q�]|�F����Oc:��d̗�J�ToU�{�_�w�O��}^���z�	�T�빫en��ꕺ_�Զ��~�������9.<3�qC� ʿnу��*�[�^V2z/��c��ˀI���'k&�*iW��}p"�o���BU���? < A�g�^i�0�)���8:��,t(���:�Q�����r��|������Í�r7e�[�)��\ƶs9�^v�������Eb����^��w�����Y-�t��%\X�T���X}��<ӝ�[p�������/k����w;��"�f�'d7"�6�O���&b'��r�+���JsH��3����F��kWP��Yc���5�V+f�u���tjz�۬ܺ��2e8i��x��B�Z�ex�\���^�vx*#��f��������j��*�ߝ��̪H+�к:�O�0o�༬4:�^`�i]tts>}tm�f�߁�p������c�����x�w|&qr]E@��y���4g}^���.j��i<O�^|�O;xԪ����^�ͳ}�����|��s�vL5�L� T�:�!I�&�E>�+A�-`�""��
"�^�h�Vc�_�G鏦~������E �9߾�}�g<i�<�Q7KY�ۦ�`���R��C�3z��Yk ��.��������]�uw�dk���1o�I�1Ü<�p��f��O��-ձ.�f��úS�PE��sҫw?{�ⲽ���~��U4|)��р��y�o�.��v��6r���D��=��ù����Cus3a�3@�4�ZCp;��}����
�^���0_=��a�r~9����2 �X!�3�Ԯ��x왃r�#�&����,n�07���3��om�\�]�n�ܯK�鈮�kEE
퉬�4P;/�:�6����51�ۋ��|2�ujnk���ӏso@�.=�v"�[9'Z	](iE�?���������,|z���6����9Ti�3�;YVm�;_lv\@��t�ݷ���ѓrg�9�,��܇㟚��~�2��s�^�ɩ3�՞�70~����6�Ȫ���Ճ$ڿ����p�8p��΀���O�EB��%�>
:��[��W�Z�5:*
�U
}�d�	r�=��䆉����ʺ�+�F����+���L��\�������]1�Z�P
)�u���
�C�8=�
v�E���������!V��ޒ�)������H�C�83h �떷"�����ϽmJǻ>P�V9���syd���m�]�3(S V^_$ɏo�W.wTL5j΍�J�}ۨ9�[j9���`��!~�����{ﱿ����j�����do��=kJ/�ޮ��>�sXfu}���Cܠ4f��1l�ؽ;���Q�nv��>(�e�X-e���q-H�tM�������I[�7y�f�`�C�.�N=�U+}�y��n�_hܝv%���˟�mWS���x���˱����ʿ6�\�瑛b^GV�T��R8nh�yC��k��@�3Q��lt���Od�՝��qSc��}��z���'o&r�y���4t:�k�nn�>�j���L�B�1�o[�;���O�X((�V)9���{=�c��/�P�N_$�f��z�
��/(d' ����w�<�&'�oD*�xp��5��_XI�VSu���M���r]����4�z=釻�@�]D��s����V;�s�Ր�#.4�&�[@�ñn'�+����Z��c���\V�[��fo�,��LC�$�7�h:{�]vdt�ˢ�'fi�6Y�%Oq�o��"��?~���p��1:�y*�1���ז��ĎX��Ԙ+~�Yz�8�>���gi��Dۊ�{ѱR�c;�{�O�P(�b��;��>t��B����ң�]���Z�G"�������G\d;��w��0;��v`���Y��US�l�W4�e��*��}W0����'Ǿ�=^I��+�=���U��������$
ꑃz7��}��«9����UQޓh��Q>���k!���<o:�������Q�vF��Cy�k�gU�ǽ�%f�8B�?>>{�V&�{�����b�����=����k�|A�n�<��9Y5˔�����6>���b,����Xˍ��Y�x�9�s\�y��~H�A@R X
@;������s�~�{��8w����m>��M�O�+�{����Q���E���5F79���Ǯ�Б�{Te`݉�G�Ùv�t������r�hE��:5�U��U,&�6�./�B#�&	@g`W�r�lG{�|�'��PGzآg����[e�����Q��?*��#;�AT���d�����9��î[�'��G+vt��P��(z�U�ʏ~���Bw��h\M���#I��� �<d�Q��u�\9g����
��u�@��>�,����k&V=��t��Y�u���"�
H(�,"�d���_�{�|���\�\��_� �2a�I�	]��i�n�G~�{�����(���؆!�T̫Ӯ�d;w��ܗf��7b^p'1�o����(��:�ϼ��{1�M[�Ӿ��@��%�&��;���10��ձW�+������7��y�8�ߢѽ$W�o\�_
��2����c.�_R��3�+�R9��~ܑ�����R�o_v���n����ў��Q�Q�A�=�>cz@VJi�DJ�+�s���;���PD�
�5���Ͻk�+�#����`�GV���.گu��.�~n��Q%�^.�kջ���!?w�u��B�Wy�ё�}0u.�1I�ZK� ~�׳Ë���bՄ](5�_���b��a��裂+1 �y���Įr�2fOv�>�[:�OE5ƀK-��D��a��dƻg���Y��`�w��sjq��5xL{#�"�VVz~�2��e%�~5��9��.8��8����74���1�G��ǝU:�S�	fʹԳ�M��u���U!dg�����f��c�!=���ح���M�yN�R~T�6�<���ux�V�v�hފ2^�ٻ�ѻ>B����L��]j�w5a�8�_L�h�Ǟ�m���֫� .f��vc:�y"��J�3���\5{S�ev�q�Ʒ��n�{}�%�Rw�.�Z ,���&F�gnl�2��a���9&pL����j�..�=�c(�r*�2`vu�]��b��@��S]�*p��V��\yN�\����;[z��Cl��k���g�"�b���������,7+�]w�wj'��L[_j�5,֣ڛ��RE�n�ӏj(ź��u:��[�T�u^��uWi�$����D���UIx��F���/wA���\ܞ��f�2�)4�'�@,՞�;���jw��:���v&��_�c���|��=`oK���D��kB�������;�+�K�*]�y�΄dD�;9�A���y�LE,�^��/�3���$Fyf wW
&�����׆�rNׯ�
�	�f�SUi+��Y-�6L��YĮ�Z��`5æ@��H���t����ޜ��4�G�##N8���r�q�w�Y譍�K�Uo��N�;�f*�1v����F�]E������J	|��ѿ@p�A"��`8q5b��b44�ʬcZα�n4�eݣM��j��WUiUwWQh�֭ 1�p=����#�LX��@�	2Qx�>gvn�H#���ݢR��TX�[j7VUX��Z֍UTVe���e�E���RU]\�p�R(aA|
ӻ���~���C	@*�U���]R�B�]�4PRD��f�8	Ȇ��0`�I8Ix"�������Ǥ� �Ck��X�,c �`i�WȰ�- �Ƙ��@�����'��Bk@ �	p"=�~�s�Ǿ�^������CnfK[g���9������ʌUǽ����~�/����~��_g��y��/}�T�f���[��V��B��ni����s�c,�y=�O?P/?��`O(�KN_��㛘�߳���ޜ:̏�dcUX�rc�Jh��(�وwR�~"0���w��|E��Eg
���^c����_Q��o�h���4��V6	R��;��*+�gݳx���m|`��ˡf���ƫŰ�~O;�"6�������ެ��n�`�\�V>�r�(#�h+r�0r�Y�:I�ˤʊ��	^�!6�n~�����;�[T"�Ti��4�� �L%X�+;�u���y���~����ܽ�=�*����<e�|b�
�!}Q@��VU�Z�x*j��+:��ݜ92EHrX���^W�{WmC��ͺ��F<��=8֮�u��U�;�kb�"�QDV6����vN@�q������=���븶bn����)!�^sAP�7K��5�&�i�����1aV�����;�g{����Q>[;���v�"U����K�xaL�P���7ի�����Pa�d��9�e(�:p��&���W"���h�L/v=p�U�|fj;�$jLs5�F5�q�Vf)|bjP>�H���WU�47��WǮ)����g����.7g���]����GB������d��'Xˮ[�}x���Ir>���(��8�~I{#��s[}~bZj����j�G�&a�9j&K|�7N6���6=Ѕr���/�x-Q�[!�f4Tp=ѩ3I8Ggw�\w0�=[m�V:��f�_vj���I�x�Q����NVB�n�n�z�|e_&b�
O]�P�Y].o'��$�$G?��(ѐG�=�[j���Wg(C%�vtښ.�>��!Q�ȸ�Kg��	�ĵ7��%Y��`?W`�?�n��a�b�v9�\n%Պgd�,��n���:N�d�ą[���L[����ځ��2ј&w.B�\7]G�t2�zcw�����Ljፗ�ps����8�c~��|U~�ʠ&�jcVΫë��9wY�'=�fLӂ���{��7b(�H)vR����^�*��h9d��j,p��Un^!i$�˅v�D�@C�]๸'� ��,f]��"s����{8�@[s�L��)t�'�q&�.Ź��}|+�#�(W�q-�{Ob�sǱb��o��0g��h�
�7���9��2,u�/��xE���v;A�'���n�z��{^�g8� YT�z�'������:(����[��w{��^��*���MV�<��\���ڲ� ~[��o�x�����雴�[�ӜW����u7��JΗ�]��RTǽ�5|���N��m���L����(V�R�7�ڡy�Y��T�i�\�ѿ�<�R�p��zm0Q�����U��?y�k�prk6��A8v890��Z7�R�!�[�3OƄ�L<��0���vl�|��ǎ����'u�� /�4&��`$Y,��	�/�F��U6�m��4���^漰��m{+5��R<�7���\�߸� ^��yU�7~�������Ԝ��5J������j�MW��]nq�ߺ�uM���3��m��h�n�d��A�䇌����G���iBtf#�'��Z�/����gS[�θ	��qM-s?r�
�l�&���W��,����G#z�Bٽ�z��;Ii3}u�Օ�A&`�Tj��z��m"��u6�K�?{�7��0��D����O��{w��d5j��)��da�N�4ɔ��U��H��ɼ1�9��^�m�`�� fl�ם_:1>㞊*��
�_]�����j�:���5�\�g"�w�G�9@�V�O[�P��d���N.^-��o
� "�Iq��|�`E��v[ޕ����Ī��?~�����#/h)���ɾN�*0��U��jE�Z�h,�zi#y������6*�=f���9�ni��Pj�s�WR��d�?"6���De���|si�yo�:���5�e�@C��� ��^M��e�D��H�H��:g�}$�舫��N���5~�U�S��{ޑ�,ٳ1�j�ȝ�����u:'�D�Y-��N
�蹉��F�o�p���]EaדCqE�(J�� �y!}i=ǒ]VSQ9żM����S��o��-q;����ط1>��Q^�[�1��w�x"Q��=���� �od��̘�9"���7�v*tig<oހ����/ʠA�Dw�Y�&mq՗����c��#d.��Z�Zu��������]�z��z����pل��N�G��� <����}��
����Y����j�v�|���3оO/1�?\f�����[�gmc����&uo���,�j�P:��*��@�i�U�KRe�P�!e��R�C�K���s�ݦ�����>�ws��zm�X�Ay{"7F��\kL��Y��UڨNC�)��V�x7H��Z/�p¼�)K�ݯͭ��Vp���8�+l�i:"T�Ӓa�Kz%L����u�Q�p˕�Z��{�'�ݘ�{^zy.���5[T �w�OB�Xq�7.�*ޙx�5?�UN���
�v�^��
}}<3����� FK��ё"S~�R3���^�{|��2�>ެGs�Fc����^��Ύ��s���T�*��/2U��Fq�"��y��F�����u�F�֪Z&�mŨ���Ed��Wyn.��tZ�ԑ��:um=��W+��+&z�M]s����<�~C)�\����>�e��GV <��G���0����]�.a�`�������_�أI�yp�������cf��u��\�ܕҩ���e�b�^���}�YEvN_I��N4�ld-���J=�fl�	 ���-�:��������SW��N5n�ƽ�_�&��Fa"��Ӳ<O�2�K&{kc��a�c4�f�J`�P�o���K�n�gd�]�w!0zM�/
jd��xgo�6ў�}8?_d#�ڤ&�r�(.�w�At��2:�$�
:n��{2�=*�ے����6�p�m�Þ��w$fb��=n>����^�Z���'~�J���Q�ޢ��V3[{|����@�]�;yE >U�o��l�"����;���������\�zQm%vů��x������g������:�})C���8[��};�����d���I��"rp�\�3$�s��!��T(-��m��\����S�,%���a���,Da$��Ha�AM�N�0f2F��k[E4��*Ţ�\`�`hZ������-�۬^��#4�m�x�J�%2����cM]���UwE����X�k:�j�Uv2��-�X�K��!8ZH K	~Mn��?	�*���An��*��j��ʖ�tڦ1�kX�)�wIh�YJ�/Ux�Uwp�b6�j����Q�cZ֍4U�[l�Q*�����UE%�e�mYEU"�^+ZΕ�P-&��J(�iӇ�U��T�Ҭ�^��E�Ym�jT�Ta�����EQ�������V���Wf.ˬ!J-ܦ+K�q�X�[F��3���I�J����ݷ7�Cl#ع��h����{�r�����r�s2I�ԯ�ǭJ'�����@�`)�'\S��N���sp'�/yf���/�ˍep�5=��~[Հ��4,�m��A�m>�N~B�;�Vj����ڵ�����t�LƳu�K��w�P�� 7K�7}�8���1��!����|��ǭ�Μ�3�N�th�u�.��`�5���A �Tv��k@8����`��U*r^a�6�E!u�p�4w��dڝ�����B��$��D�����n�Ć1�a�Z��3x��_�^�O�$��"�LVP���u���w�4?�*^�b��[/��&�H��첝���܅:��¸��J�hH���1�#��z��c�3ᱯ_�n�j�|���z����O�t���j@g��#7׋��B��{=.�h8�ǅ���r�����ˊdS�"8��R�6�׻���a:O�=��>�~3��]�ݜ�ݯ�A���U]_�|���HF�i=ɛpu�]�`��Ӽ} ��2R�&^q�=9�]�����mA���)��r�I��;Ԣϑ�O�Hz�n��B#���aW�����'�c�Rg���&5��l�vg7"eg=��qQ��H��񪑖(I.��]]<*M꽯�TH&y��h]�7b�{�mGyot��}V5�)���[�Ό�L�O��xW��
��B���col�}�ò2�uf(D��Й9	�e@�\W!�����u��v~�+��.D�{ղ�� ����q��V&����xml��Dga�fXq��mɑ���:���m��ʠ�s��?+/���LUn�0]u�]Y��f����SڧN(��s�Wc�*�kf�����;�.�{�Ϸ�a%�{����u�8Z�ԸN��ς�X�8q �w��=ۥ{��]��tP7��dq����s/v�mѨD��x w_!��Nw�a���K�C�@�\R8V�	|v�W~t9�w��C���k)�B�y�&}^^m����,�iͿl-=@�nLb����ِ}�(3������a���`C�zY��^��ͻ�o���Ԉ�J;\$EE��-ܬ�
�9&9��F��V!�]G��*�����O�jEE�6��֩��X{��?�_4*��o�y�_l��»ٛnE��)�YIk{3�Ml��<����U�N��uI�h;�����Ӫ(پ5Eӯ�v[�����V�z�b=��
�����ʮr�	� ��0��>&~�X��8z���3Us��+O�כ�5�s"+����u늱�a;	]s.=FD����Ƚ�'e���ɉz�X��I,�n	5�x+Sc)3�D�3-��̠�i��N)�8o"��(��qGnk��~�f@R�����ae��8@Z��؄ozv7*h����5�<�\M�����xaD^�/�U��7`�������3WJ�_��.V�~c���������L�m��'��CvȨ���W̛Ɩ�-���[�r�n��DY=��h��{4��|�:���5Z1�x{��xV��Z�}vx�t��wTꜸ���̒�-���>�������<K��ѽ�L�Eڢ���]<�]:��ai���'ʽWt��Y�R�����,���dǰc�M!k}Z:b�7$x�M<�3[�����X9F2��$'N0ɽ<�� �\J�g��d����Eb� ݝ7=�5�9E��^�}��0Da"o����/L{��ͮ�ߓ�#�Wp��?�E��:=��a��&vZX�� o��%잙�# uϯ=�P�Ε 7 tN�*���h��WW�/�?Z�Ax�g�/�ڰ�66�rG��}=+MZ� �������*�J�V�$"�$�2�=�a Q�>�������]� 7��2��৅�q�tFWs�]�n�7� �[Fv��	��L�:���9�z*�f��Tv���5ϛCw9��R����9�
�-?/
?������I{�O�fl<�]�ty9|�H��;Q������{˟��oy�s�g�^;�T��V/֤~xR�_TCT^���j��6f��W׷��=}�hXx��a�l�W���hg7j�X�E��s���+�h�p�
țbe՚����vSrH���:Jv��C,�]1��Y'9�na�*�|@�2�@��N���C��[�ӈ܅ 77�q1>���N�Q֒+h�ItN�F't֜2��R�@�f�Vw�ߺ���Ɲ��
�aܩ����.�q����˞뗥�|�(��S(�;:��f��<[0����;X�?G`ۮ�1�Ή�MG5�|9cx��7y�T�ޏZ��-U��*�i9�r]���ZV�MKw+��V�#�c�-���pN@�m�ǲ;r��1ky4�]l�=m��&*P؋P�Tw��l����3>K��fɹ>R�K.v�x@��{��.S��yu�~ڈb��?�_�3:���(xr���a���r-�"�u�����3A��:ѿV�x�d���ZEE�\V�����"OWPwt^I��|=Ҡw��ׅ_��c����jH��/��r'��w�Ee��6ٞ���u��Ii��|dsڏz!D�����aǬR��;�\��H��O)�GA��_?D�Q�y�J����n����m]ڑa�
���G���?;�l�l��r�>��[�&��nr�r�w��쪵����'�����br��a�*�UlWYwWYܡ0��͚%�L.L�p�
Gh�s����(�MKFU��(]�r_}�d�C`���Pf��V�0�K�{�'|3i��!9��ܖ�%�7W1�F��K�����#�*�9��z�4�C��lL��r��M�L�W�O�K���o���^I�?-:�W�
�O��v�c�f��)�����#�v��U�u���'�SW4֪��:ݹJR�;��L4�D沝p49٬s5ݵ�N}�\��6����W}��XdpR�>(y�*%�E[Qx��b^��9i:f^`�.Ƈ+�(�Kb���=��e}�&\�4��J/��T� ����O<�#�v��Ԏ�κt)7����NDK.yw�7�d�����:�0��c؝x'�����L��c�Z��c�VNr�<L��2�j�T܌9Q7�S�<�`��,�U��
�.���0���M������II$"JI��J��9�o�����OR����F4��s�$�	˺1x��E�c;Ζ0ίU�Z�8��*�tP[UAx�n�ZΜ�muU*�n�v�i�NqT./ִ&���U����Iwֵ��#-)��+Qn�t-#��x�����ִ�sD�b�"c(/*�DF�ִ9i�WB�QT�]Պ�#T�j�Tl����xֳ�c�+IW��]�
Z��.�
����gJ�+TR��B"1����AEWV�Ac)�Tp˺PYMDqUm�Ba�)�����Ȼuu2P@ V4ey����e*�9�e��8�_�SyQ�Y���<;�	�#m�҃1�bJ=3�tW��$[I����Q]��Ȏ�<-�XC9�	8₾����u�c�\�+�.�ڽ��O��tz�4��gTOy�r�bn%X�s�8΀gT�O�A7�_Fd�"��X���0������0+o�u������U;�x����vl�D�1������˽�r��m��ѧ(L�<�̎�7b�}�_�c��w��x+��>�N�L�ۡ�%�w���]���p¥N֚�v�|̣r�(b���'<a�w��l}d��o�2�z��Jp`�?�vE�e�#�ƕΙ�Ɓ#�L�0/G[UZ6��(G�7rL�� ��WK.ސDg�?g������S�f�i�
=ޕ�?X�Ϯ���r�EO�#�0���[�Id�����0Z܅���Ms���^���*�����T�*5�5�4!,zNr��GY��
u�m�D����Md�;-#���p�K���̭�y��7�*�^˧�i��.�'1t�����@Ӣ�̦��J��:�O;	V��N]�k�m\^��O�wh�]5c����fܳ�����J�F�|���|���q�F�w&a������[�v�Y��v��� �T t�٪X�M��eV4,Ra�a�k��:)�[-��𸒳#���q�9�;�����yW��Y[=Hߐ��%�s�@%��-M�C�C˞WA�2��p��U����=��YW� m�-كu:��g�A\9�-�s���ٮ��ud��.]ڍ%��p�:,q��
)P�"�Z����T^oL�t>"�|��YSP6�|��c����9֌t�EY��7���k"�.�i��x[�U�%ޡ�y�`	�[��(�8W�.�>\�!LQ��lY�gu�f��k�s�/g6�
��Uv;����#�-/�Ю��l
�{�����(8�8���4�/uj[��-�S�}�꣣�9_w���_���]�G�,�ѿ�LFj;�.ab�q���m��
��e�j�������N\ն�W�����	m�M���4!<��z�FFb���p7��V�ZbF��Ls��и��oES�ŋ�QH�Q#��
R3nG\I{m��թ�LwW����+���X��'�|"|�z�Lf�U��ظ��i{=v�u�N��n�� ����P�F��5�[�y���˹�3|���撚�f����M;�}�>LL��{vк�v�:d,9�;�A-�[��v!���v7�C�/������l)h��Zl��z �;��N�#�Q��5$�ZyN.^-�M�� ���D�K�o��]ǣI�U��Yԩ�L��{嘎�~V2񐾺���2�f۴�o\�t��M!��.1)����=i���.����d�cY�j�J�mq�T]�0�Aj����D������)�X�d�
����zFxϱ`�����
�z�6EB=��Ш�݁�ck_�]b�~s(E�s�u2�6I�HӉbV�^�	x(5��apۮ���3G@ڵ�_^K7�U�:,,˧s�g��f�VV)��Y�]a֔���4��O����O��)�� ��=������G���]�iS�;���7N�L��{pr���2ν21�>�h�
��ϫ�줵�ܛ�z煅xY�Σ_d�����O��U����4Ҹ"g^a�Vy�5�������ۯ�>�b���ow��q���|"����a�Y�;���;���`�c������|�vG���;�����c�|�!V7����Q��?�PW)�y�X�F��쾯v�m�T�)�z0�y1���oy����K�E�� 2��-	�U�[�8��p��3��v�k��x�Q�	P&hc�ͽ&�D[~�}F�����+/��r}��Z�8�\��aW�X�:�:��m������\4���؏��N_����3�э@��y=`vd�P���a�"��cJ^��`��oM��֝q�i�W�{�=j�T�g�}l�3�+��1�1�����6,�,�y=#x��4���q[3y1O1��;����|��e��s�ky%�y�F���E����5�/��j>-�4�qg,玴��p9$� 8�@���~����~�l�M�}�� od�1�l���zU��厡��8��zȊ��*6p-J+*,SF��Y`2�xgC�^�uR��Q�h���:�;؀����p�\WS|x�A�c��듑9��p�﬏�b�IB��$j\�>�7��s,6�1TUo`�d�٦y���
W${�O�/:v*���;&Y����Ѝ o�o�		��}��O�!7����w���Om�a�r��ĕ��������n��F4 G@�n��������3lc�q��C���sk�!Qު�{��ׅ�������>R.i�ǰ\�Z�^W�<����)p����;:������܏��z0yLb�!i�٤F��o��!X^V�E�m��H�g�g���U����-�m�^�d���e`]sǹ�e����vБPet]SJ?t4�f�A��Fڲ�P`��`��ˀ�@�#tQ���9B'��,��5�Z>r��dl��11-0]��v�f�������gFq@z�%��Ԑ,�(Ub���"E�- ���$�/RI$^Bԥ���(�+�,�k@�d�d�*����
  ����AP��� 1T	B�
E
�(�QB�*@`��% �� 0@B�*(QAE
�P�B��(�QB�
J"����\��^�`�d�t�m������-�D�&�RU�C�(���D��
Z�T���gD�l����;���=����-�	16;*R�ŉ�-9�pXт0��۫	��Gar�Y�ES�/�R�m��ТR�͍q�e���X���BO�{l�����_���4�!�T��"r|J��)P�K�h���&�C��$��C���m�>SsS�.�k�sx���g3��$�g�萄$�����ު�Yܨ�J:�OB�g��3v��1R4�%��+�k���Q�'m������L*�X����vpQ�����gm����2���z���%�)�~KMr��-�`ʗ���ja$& ��Ł0�n�% �u���h�,��~Y��Z�b�|��T�Y��S�b��� ���ZE��@�BE�$Z��Z�(�J(]�dx��kjt���&�c�#Z��{}]�MC$�>
��|�vC�������Ư'�nf�>������k�����k�)-$Bb���$��&�N�|��ԍ���}mvoL��q�o"瞴�{�g����n�9ʭ�'$��}�q�֏3�v�=S'���{�4t9�Bl�����(RU�>}iEgS����к���a��:�E�����8В!%��!I�����Ԕ��4���:���\��&�Jhc$nb�ɺ�B&I�8/J*����/-r�IG���)YH����b�������rt�$��b�cn
�EFk���d�~�%4�L2�I)A����rznp`���r��:j�D)c��g{�����t�˪B�إz;�~�$�l�<�9�K������>ËTqI֛�od}�í:�\��XW�vҋ���(�-��ks��C�o���^=��<�{��k�c�ZB��뜱e��\����܋ZY���ҍqS�!Ih����4�~�|ƇBp�n<~��z7N$�oG�{3֌�*TQ��K�;}��pR������y`Y�C<=�V�uJ�#4��#V����uUe��9���5%��:%Uo��7�!Iw:sGJ1Ȭ-M�w'&�07�9�1*�z�,�y�6�'�Rm�]E֍;,���Hm����QY�^Sa�:*%H���*t���oJ6k�#�OI��t�m{�wD����O[����4��g��L�q��`�z�����<��,�q*�zX�GdQ_�B{77��z�s���"�(HP�؀