BZh91AY&SYS,�r}_�py����߰����  `�~j   (  ^���� �Pҵ�� (�*�U  *R
  7�"WfJ\�Z��H�0��ҁT�� 	P P
>�� �_zۻ[�gUݙ��ݚ��O���>�z��϶�!'����B����Ã��v�K�����G���w@.ۻ��F;4M�J^@${���� ��)�`��Z�@՝:6Zڪ����_{�����g6��$pw
=��K��va���yoG=�C��>�ֻ��wwV���Q�ʹ�� <>z�����e��.�l�tѹҹ�������۞��G��{�;R������ַ�u��r�}t[��[-��_� >,� �l:�l��۵��vv��w}���ރ��-�w� <	�y����m�p��۞�e{��:��5n�����]��W�G���� ���k�o�-���[�g}��k�e��u;�������#���l��s�۱mm�;��ӄ棵�n��B��P
 $)@  @  
�@    ��F��U*�LM�@2A�0���jx@���0� ` &�%*M
���&� � &   i�P$�Ti� &   #@aH�J�444�#)����j����Ʃ�x�*���(�i0&F 0 � 24�O���L������T�]��O������ vn�߾�8��� C�A�������  ���T.�������?�������G�l?��������@in��T�O��QU@tDOD�P[H	�@5t (&�����Y�������G��9���ǉ������L�=t�gH�a�l�á9�8W��3p�'�ޒ{�zIgH�A:�/�Rd��k��8[�m��&�Vq;`���2�_��D��D-�A#�E�C�r}���C�u����Z�S$�6ɶMi"u8P���"x�{��_pI�<���䇏���M�����%a:$Y�=�%x~�I���7gXJ5�<�,w�pzY�N0�${#�)�:='��d�F��丑�H��%�'�vO�3d�4DM������Q:'�Z��"hy	���O[�V����\"t�D�xI:M�ZH�H����D���NpDvt������K({���H��'�i-����'Au�"s�'�p�|Nu�>Fx�h�$D�$D��I�E}���DGŔ?pK�&��"t{�P����NC�҇�%�'����<$N	��P�xIbsI�I��C�i�|��W�%
Y9�l�'�lFB?t��9��7�"xD���p���Л�W
�IU&�'����m�H�O
x��������dQ7R�K�%�<����"q8W%����NЏ�9�UT��pM�F��e��]w��::�~�<^�InY�D�U(��9���Gĉ�C�����[�#�B{By�xC�w����6;��V�4xR���
��m8�N��;�7���U�=J��bl�=�*DG�Qt�x�Du��tNG���F��Du:{��O��K�T�L¬�U3�ӧ8lv����/SfNGY�|����`Pp�h���x!䲯�RCC%���_95sܟDO}�����D�:��;Sb6H��"q��P?m��pA��6[4Y�.DG������"5����P���+C��#�TD�ȝ�TOmO��TD�K��D}'���C������@���u�:hFO&�&��%	�8tk���h~9D���">$D�Mn�">���}S��ڞ8WZ�'Z�f�܈��Q�S��>MA�TD}uG�H��SŕmO�$����Dyʈ�ʉ¼M]O�wU�D~�Ϫt��S�
�S��U,Л��*":jp�C'��TMAr�hNH�jx�����?P��\�A�J���4>�D�"'t�C��#��ؙȎ�'�A��ڟ<�w�$��
<T�(J���;��C��v�r}.}q4h��=�ZwQ5��np�z�D����k�d:'�FDNi���4�;��>��jT��j|�v�A<I!�`����C�O�����f�+�O�ϑ��'�Su(~���ѩ��N�H�elG|�㺉gm)=ԤJ<y�;�:x����42Q.s�O�O�}�}\�Q�`����@�\� �"�wȊ�-y��b�+23�g���C�=m֍�K�)M��U�#���{�(4V�4S/�p#�����h��hwDkL�F@L����\	f�a�=���4����g"�R=�ݦ�Y׈�h��p��
0�[ø��;��Dl1�E��g��Yhv�׈���0���wMp��E.t�1M��5�{g�{���l4K'��Y�=���0�8�<�#G�vZ�����3�6m@4�Q{ZG�G���=g�D��G��h�5^[�.��q����
�=��p�6γ�'#���i|N6�aYh��F�,��&͈�G��c�#���=Ķ�;�m�
:�P�qo.oA����nODu�(~��4q(O;&����6Bp��J�*P�<��nn����,��DK�*����wU���J#�ODN������lM��+d�BhJ{)�,�ג�ïJ����4:�Bq�"<�l����"Z�ᣯ�,u�_#�f˯�lj"<䯑�\ԤG��|�ڕ�4�R'�D]�ᴳz�=��gYҎ�ȉ�N�e�"mԤG�(y���5)N�"'dD]J�c�J���JK5z�bm�M���2����D��H��+��?O:쯟�U�4�5��Оw)4{_O��R�4�R'�"�W�rW��e"k��bm䤴����/t+��W�V7�tU����'�r�O���,�H��d��\8`�h�$w�JIwa[���tDta�lM�A�x�D��eX��Uӆ�g�#A�Ñ����l18��$/�J���PHE�.CMQR�#sbm��<"�Wn,��+��k��r��4:��uD~��,jX�yU�<�W=#}�M����I)�9���5,����G�r'��U]䮚:�>�G�N�j��;���:�?x�Nԃ�|���;���>��zt����/��/�	�%�9��w��%� �\RO�'ԓ�+��qF�wI)I.� :$�ҡ;��>ԟPб$�$�$���u���bW����:)�T����t�Mp�P��"��+�ج�L�I��q2��+�}�o|��m��4	�S�����S�}W�+'�u��B�#��8G8j@�S@�dRp�$�u<�'ˢN��_�I�Ro�'1���t���+��É�%r>5]%�����D�9���{�:<)�5�H���x��<(�~9�h�m/i6���Rw��N�f��}5*V+��l���/�_�O�T?��蟞�Q?����B�ȥ��� o�^�I�)�z�VR�إ�3�K0�M�� ��Ӥ	j��;��*��at���h�%�J>F+t��X�~e\֫
s
g0�1|tZ�G
,���F�L������ѣ�kZx�gS"�8Y�KT��'Ý�����	8D��G$�d��6]'�gJ�#�:�F_�@n����ݽ|wm�"�_>д�6j�BB�U��JlzMph���Nq����r��ɲ����ڙB�)G�PLZY�]��c:ka�@|����[�R^�)L�!7���!(fdFτ&���ݽz��g��i�nL��k�^��.��֌>�N᫊Dv#��f��1�몣gH��_H���B*Svp�X��t=��>����O/RtY���������:u�a9L#�u�7�)�!��8^�Χ�{��l����kˏM�5�2�i�vrU�8r�wT&ܣ.�x��i�[��n�F�^1l�q�yR��ׁQ�p�,܎�*�U�e�����t�}�U5�S������?�Q�g�0���"�g��u�[V����xª��ݛ�gWvW�3�����#Nb�G%8��)�Y 캕a.6YD�v|	��n��=m�)�P�(�%}YD��e>���Z�[��������s���{>i�������Ǿ͛�'�*B����)�́�(Λ�~��G����a� ��$)yݻ��6 @!H3bmnl����㷒�b��3g��aD�3(?C�Sn���
<Ig�3�C�4p�>3� ��N���{?�k������d
l�gT�i�Zo[��z�k���١�x�[dֿS��4gbO���xv���t��*��,�N��Q�/��[D]W����a��	=:%����>m��
��
�>l����ϮH�^��!�e����e���l�{�	��2>(�w���->�)_e�C.���t����
����	X�%��b��f��o��l��M��8@�L�F�v|�`c��<%���A�B�d�%k8��n/a�a��i5�ؕ�q�x��p��}<�Z�[e�	�`X��,��-��Շ��8|p�%�D�@"X@YI�"��Tl|�so�(p[����љFp��8EoI�1���v��N�~��g6{y` <�Û=���j?2���š��p��F�P'�ڶ��/���*>����:l��i\�F�Æ&3Fl� eu�d5�݅Fʾk�Ë��b�Ǌ?���׎���=̟Q�#��V����.��pR�F��I����;(l��M׉�vO�l��$Eu���;|t�Տ�TYp�I(x�e��}w�kn�JoU�t��$�xr<ڣ��C_�I�pe}4�1SO����؊e!�Ή��-���Ivf�d���w1��҉����
(����?S�Gǣ+y�l
�y�eY�����ǧ���Љ�#^BiFO�F��KSꅧ�{�7�e������ڏ֦v��N��oq���IÛ��s%���5���^fv�����EX{>��k��K(�_a�j�,&�j�gPܖ��*��Ǫ�,�Q��6^7�a귤�t�{��DI�a޾�wY�I͇:7��$�V�N�jUu8��D���Y�� U�l�)
�O^:{^�:2�����ѣnN�n���貰�F�������S�,`h;��/�0v3��o�r��|��>H�@<l^�t,�7G���4h��p�p��:x�o���wU3��f(p顔��g9���]�h���d:h���)���6��O]?I�:p=�&�<8����u��=�YZ����o3�͒l��M���j7�>tr��M�a�jM�9�좊/#<R�zI�4l��`l��a	�M����W[ܐ}y�3��=��l�08R� 	���hjE�l��8&h�F�ݽ��/D���+��Vp�4t����dȼsj�$ꊑ��̛xl�Ӓ�" �:l�Ç�^e��=�de�h�����r��gWD801/;68�J7�es����G�/�ju�g+�!�s(�^�&C���ӣD�|�t�:Y�S<I�k �L�y��[U(�g	8b	6Qd	_T����;��
T��wO��>��.�w�|���m*���:p����q�Ĕh�ҍ(ͮj�-��ʉK`�M�x]c����^�(���p�:��aYTWm;��}�
B��z�Ş=V����\�ģ�΅�M��Ǿ����:h�U�qZ�W+�K&a쀽Q��0�:��������9%#��$�r�ILd*]�0U��+��ޮ,�-�j�Uk���N+a�OV�V蟲V]�H-6��l$[!�>8nH�|Y,&�LÒ��:\�ڭ����ιn�e�w{�On���F�:�Crk��p�-å!E��6U�V��[�L?�^��D������֚�uV�h�7����0�M\r�ǸE6��U���\��Q�����ѣ�U?��O�L U�\Yj��I�����.x�q����l��"��u���a�9q�͕8����vY�F�R��ӥ���HM=:wum���_>4h��'iV|(�t��T�g|�F�=xI��@�P��ˬ�E��Ԧ�<a]��:�c���g�;�~{)��y�^m�sP����E^�d���Yͷ͉w�Z��`�?�����ɏ��O�Gߟ�����!��?:�[��O�I�$��J'�?3����s�͕f岯�"eAj�씌e��S!�s�6�w�c��u�>���]l+]�Ln:����e)�T��f�͊	(`b$��]���}�j��[cQ��XJRK�����@.��7��Š3�=�j��-�eon�	���e�`(\N&��-��V� �GpOX�MtVTY^D!�]*��� P]ӭ4�i9���,�/��'���l!	f5�4����$ڐ����|{Yt�Qz�}z�v3���e��2Z��[bm�Ne�6iN9�:ҭ� Д4-�AZ��"��_K2^�	/c�J������.5P�F-K3"{xŦ���LRd"��u]W���4�hwĥig�z��~=�Ѥ�����iu�k�]������z�"�
�B	�:�C�J�Q��&KUo>�wa�қ5N�j�w�#{����Y�o�8�o������qey�b��I���������=�."�"U�jU�Q��=�g��%�*[�L78�E������b۴�;��z�ס���Tb��y�]z�ؒft�s9$�9��q�G%Pn*w���ku�W�Lj\��D��"��=�H�_��|����7T*T1f�J���T�@�35�r�En�k!x݆H��R��Ŋ�`E:��꠻W�/c^�d�<=��iq�9;���w
�' �)y8%��.�b�p].����=�l[��!S�+�3��H�!�P�+I5��U	|e��x���}�3�TZ���n��MR����ש���<�r8����{��?ց���g�O�"

��������z*�/��{Ä,�2��O��O������ ��P��i$��/��?��������UmUmWj��[UҪ�b���UUV*��Uz����t����]*�ت�եWj��J�����UU|�UUX���UUTUb��yUz��U⮖�@H'�	! ��!���9� �5 XEE�@	�U�� 	���J��Ҫ�V�U�U[Uڴ��U�Uz��U��U_"���*��iU�ҺEUW�UW��UګjӭR����J��WJ��]*�t��Uv�ڪڮ�i�Đ	 �YDY	Y >�O�>���@��>�U�8���*��4��|�U^�*�UmUmWj�j�UҪ�b���UUQUmWjҪ�EUWΩU{�t��kJ��U�ڮ�V�v����Ux��Uz���եWa�����|}'���}!��(�D��V�y)VI����s��U򴪯U�Uz�UWȪ�ե_1z���եU�]��UmWJ�Ŋ��t��U�iU^����*���ݪ��t��եUW�UU�Ҫ�����UU��[��}��H}� |n\�K�R��WP ��#�����,��"�B��I�'b�PLB�"�,���~?�R��$'�q�����������������~z?3�A�q�	�<""x��,�"P��<'H�J4"%���6'�h�6hMA(J,D��"%�b"xO��,KblM�BQpCDC`�K ���ı8x؆�	��:t�""pDO	e"%�b'DO���f� � �x�&�ѡbhD�����4Y4E����T�ؤ��Q�[~t�|ۦ�ɋ��r�]�Kv�
�}���Lul�
:`Ӫ��e��PD�+����!��j�(��2f�a���3)����jVV�� � �:!��2���a��.ۮ�Wբ:d�+�X�mB%�k�k��#����i6�:���%�����.,H�\M]�6"ʤvb������2�j53v�c�.*�WRU4���[���!mU�VR�e�$&m�V�-�RL�3f�t|*z�����xO��Ro��7�![��G��C��>+c
��u���鋮ѕ�tI*��ˏ�UJ;�����~������o��@˓V�� ���b\��<:d�@�C��ؖF�Yl �:��ë�Ck�6�P����Xj��m��]�E�;"i�SU����(B���A{��ʹ؂1F�ZA�V��d���FЋa���Η,�.��_%>�P�GM��vM�Y�����t���,jIx�L�5,;04�h0!�>k�_�o��MeX��j��d6�cf��҃.�L�)�0�m���*�aBX7usMZ��ٟ�y'֭�	�R��DV��Fl��U��-Z͵�&mİ�G׍Vf%��b�cQf��([&
�#)]�IU�ZJ$آ>\	�˙������c�rO/�li�ŷk�د./$ĺa`���kn�V����mt/Jy.�U�,���T�lcKt]�
@��]�p2�]��YXcjM�{Ě�3[�����K#��&iuH&���Xh�Sf����;�j�RShZk���.��6ʹpMi� q1+����e�h�`��K�R�k�Cn k){�543�@���O��K,G���q����%k[�Kki��l�
��1�ar��&V�)]/�G��z�1��i�d�O�����lB\���Lpe���Һ�e�qH[s�c�ơ�X�i�b�i�09ac5��6�#�&�$��h`ͻ(=C��1.�jB����n�����Ŷ��l[��WdݨU��x�öśq����%�,g�æ;Y~�xg��ٴ��o[�������eĔ
����ٺ -�,6��[	��R��ZB�m���f�|�ޠ(]��طmfm-�M�im�:��H\�ݹ��4YH�t2�]k.d:R$��2֢�2��ZA����%�0��ƌ��X1d4�N!�4��J���z=b �^~�,��-=,�>=i=설2�[�WM,q,X�k��E�k�D��(h��3J��e�a�M��R4;Mb]^�v���n��L����j�
-�����f4��1��9��i{���ʤ���U浻�J hR6� )"��s�U��ح�*��t"�Vx��p�X�.��x�U<�r�a]���Oz[~.��6���9TL��B�-��������p��n���3������*���ڹ��������V���\����+3333Ȫ�wwj������|8x��.8��:㭺����i��S:��-[��	���"Bmm�t���%����S3�I�,Vh� Q
T]�2k\⃌4m�l�2����tкQTͽm��M�Ŗ��ڪұ�Բl�̚`0LCQ+���V0�bq��G@�]�u��̥�Ɣ��(v*Ѝ�3�jYpۖR��i�8�;q����V��#u���>g3O{�A�)vؕ+	����;R�J%LKs�]U�+6��T�b�c�RD��#j���� /\Vc�`$�����I��������]i�%F��YH�W 5�e���eL��� ibB���ÕK���#O*ں��1�P��6�CA�1�
�U�U�ؗ���Qk+���0�.~�������ѝ�Dh1|KO$:o:#1f���6U6a8���L�9�?�Y=RW��k�X���QL���-�ˉҎ;�ܚUG=�q�(H���qi�u<F�\��ƽ�n�����4��>~u�4�a��M�y��I�nI$v�M��3�(�84�;��x��D���Ϋ��o�Kf��8���jh,����I会�D���@r��a�����%�ߩʢ�!���M6�k궛W)�ԕy���tPwcw!!&@Ɖc����̼�κ��n�q�m��Z���/X	�I�H� �Hbo��km��7}���>�{���}C�
��� ^}h��IQ��0>�O<����<Z���yJ�L��h$�@�~�O�T�I���/��ZF)�g���:ҋ�!s�C0{5�MoDi0C�h��<�(�d��m�u�\u�\8�6��98KR0{� eƶ�5��{kX��-�B-���Nf�5�����Q�é�f�,�*��\rtˣ͹M��N�ǲ�<zjY���O59$W[��jec���۫#N��뎸�n�q�m��s:b�2�ŭ~8ջ+�v���U56%�IE�A�wC���"�����4 4y׺Z���P�W�Su��Gef:�����e�1T�\v�rg^BpX�UL9q����-�<F�B
�����ٺ���I����R��ɣK�h���s�<e�0FBIBZd�A�^䝔ix���4x�e�4c�k�䷇�D��eȚwԓnf��ԉ���pR)��®�ŭ��r�%�խ��m�m�q�m�8��,g�K���B�.2�� 1w�����{�b���U٠b��lě��Uk��4߫8��x^��U�f�_M"N��/#�{*{UnI�LhA#�;�E8�urJ�R�=n�<;�*�!'vG81D5Y��%=���8<m��u�q�m�8���Ih�(�&����@�����Z�^&1��������Kd�!kp��$J�l�6n�Z����\��c{l�WkUk��ܑBع�ZX�ba8F���B���OtӠ����!v�7вh7r�[N��]5[+������t��p�x��xM�����i�q���d�Jr�uqqs�1.�J���.��&ɔ�2�޵&s._u$6ă;�u2P4�׳�Z\��i�6ǝZMw��Y��#rD���f���H��^�ֶ+��Z����4Νm�]m�q֎8h4��R�dҋ	�:2�6l�*���U0�>|n��Nd�N��L�blVX۵B],e�(��czI$�&�������5�mZ]T�M3���c�
:�L�&>���+�Uu�� 3�vw�i�ݡ��
� ��f��}��LgX���U:��i�:�<Kcv�k3ms�� Zȑ�s�̫�f:y8`Z68�$��!��2�ǋX���8O�q�1�I�c	$��M.�H@�[�v6hH��P�g���"�T��o�)�QIJ��QP�@�j��iF
/�r��JR��6��8뎸�n�q�m��[��Cc�  ��5y{qT�R'�牃!rIBݯ�)�bJM��Op@}��-��"l�ː�,(L.O��\����fr��p�E\���em?v��/L�һ ��]y"SF,�Pq��,�6{.-s���zi�Lo�,�9r~�Y�>|�I�<O��
=��&	F&Q�
y:��N��_���|��G��|��>[��y<�N��id�<��yf+l�L&I°���a:a_`�ܞ[)�<�E�[��-�y,���50�<V��+*p�D��L2��5�0�XL&	FL(�(åQ±4�ej�e<��<�Ⱥ<�ͧ�E�'�Y)$�$G�"�ZJ�k��<���4��y+n�YydL���"�Ӗ�[˭���y�N<kx��p���°�h�2��
�xʐ�$�`�a꓆�CRaP��FZ=i�����DOIQ�m*��y0�0�a���yyg��(����=�|3���-�SW�HE���ۼ�c*l��KF6^�	d�zpfe��so�7�\tn�Zv��[��vJ��l�hn����U���G�Ŝ�5�Bu�����C�[�v<�U�47a{��u\x���kN�ZۓD��(�_�y�Ҏ<��l��5�kJm�<��Vt������g|(���]��YL.�u��  ��??3?<��������Ϗ�Y����"���{UϾ�+3y�����{��s���ffw3=�33/{��s���:t��<'�� �:l���*��Ҥ�ky*�����&y$�0l��#��xE�	��䅘i�l�yP��X?H�-���(s�<��>4Z.H���間@ ��p���$;v
�)��_U[�����s��M�k�,�RD�bȹa�%&�`b|ZX��L�7���i���H|C���2�{	F'���p:D�d�x]5���K���a����I(o�^"|�Yo�v��C��ul�n/���Qb@���tPD�AH�T��l�\e��>y�n6�N:|8p#C �#�Jä�$�J�P��4�qHe���Q1a���<�i�f���r5T^w#�J��d����@�!t�r�e1Jx�A����Re"9!�vӐ2d��pb�N�I�`��e-)4����C�!䁒Ζ{Mh���#)t��K���␎ `��7�4�2#iUh�;IUh�JM|�Yi�EŢD��8�r�)&,�HA*H�ŸH���h��㧎�><'��!�GM�(��F�M7`R� P^-[Ln�nH�E�4Z8"֣u�{r�ȹx��0��H�C"�v�׫m��Ɠ���D}o�D�mFїf6������f�X�Y�,��3i�ȩ�V�э-7���B���Z�
*�Xk6��hoK�\�rV&�
�Q݈3�??�����HQA�@*ŲH�qAA���h-X@�(n�H�Gڣ�œG�I6�"�Ҋ�Hu"�<��Ds$[�@TK r/ҥUUJ���2s��8;jq"S�aiL!�w�kFs&�Dqc��d0�R����	��*Hb�Ha��^$�i���E�r2^�/�(�!���f���X�qi�B�&Xd���@�5�{7�xźr����詟��4d�>���-��!!@8Ha�)M�b?$9)qA���1C\����᳦y�q�m�<��.��l�o�_���{�m��Ʊ7� ��2���RD6^�oV�C]����NKGi�Wć2B0���z��d��,���I8�7���@�*��h�h��!��S%�8�d�,��I�B`�B�CI
�q"�8��,LR��0Z�K�dZv�m�I�"���$i�(F�>�PҠ(o�|c�vA�I	%P|�7A���gFP>"l��.HQ�r��6d��H�"���w��Ja�L�R|B1��HHB�,4@�{*���6h��1�����ӌ6��^|㮺ۮq�mvs�}��A+cC�rhy�m��5��IGи�.��c�e�B&34����	�4�j&4D:B�7��Jb�*�a������2T,5�;I�	� ��E��M<P]�b�����6�Zj����k�nX�+VT�]�M��3&1��H����
4kv�t�p��FA�c-�DC�I�	�!��C8is���YNl�K0@��'�,�4�7F��.z�,��]�]��%�"�KSP̥����MA2'X�"�HH|��$��#�X�J�ٜi�u�_�ϟ�tp��@ѣ���A��y��8��7M�'���H�7s��m��i�_b1i
0?���-��'R�$X"C$�h��	���&��"C�J0�G+ᾜ@�2������h��>��(ŕ�X��ϓ��C�<�Ɋ2���!���$p�䁧n��<�:d��c��������a���fQ�h9l���%��g���E�e�h��9���BU��f���d"c���>aDB0X{�IJp��d��-�B!Δ� :��j!�X��4�i9Bf |� �xe��Eq��HH:�0��y��8뮶�yga����~L����d����56Ey��$y�dt�N��b�Q(j
6i�
�D���D�a�2�"�I$�	���Ӄ"�&��[$SwjX7n��j+��]�)
i�۠�(�Uٻ���͋w��)j�b(:a\
�5wA8L�D֏n^>tXtUD�\�)!��G���}���-��9#��I�TZ]K�$���+�#ILC�0��O�"�!�� f-��0CL(�������т'ܓ�I8rh���H}��1!�&8"�2A��	�]J�BU�"x���1p�.�I$;���*�����I9����x�$Y�op�27���Y�Gb�o���b۳-��M�$2b��$-�SnoI	�9�%E���b�>X��h��j�6�v����Q{�g��%�- '��������k˪�)�J��y�u�8뮶�h��CF �:�A/R��!Q!I��B�N��m��Xo�~3.��6�dYe�,����D�/RJqC(c���H�2�V�]�.����,0��-ń4\&̘6))����*�e���U^��*a��A!���IFq���!d�)��2�B/��H,X���S)���)�p_��|��E�1
�CM'U�fHX� �(�2�.�`�[�%"z��0��4���I%-%�]Ħ��J�2�cW�.�/O�$f�DH�*��RR�|��y�Ϝu�[uÎ<����m�c�M�<R�X̕ËZu��m��_ylljV�b|D#q2E>&pQD�tD��0�^똭h�d�n#�Jv2��jrI"<�W#iUt]vL���)�Q2C�m!�4�H�����-n�v$J(5��6tUCo!��U.��ї�=������.������2�ᴉ��0e���cL��l�t���%b�B�g�RD]^�RϾi� �B�?@�D�&���Ԅ-�2@���2*�-
a_cP��'H%nn��d(�Z[I0�KV*�}KSYd�Ͱӏ�<��u��p������Z��kkQ�k4-����6�m��H�bh7R}	��~����B͘L��@�J�Z˪-y�٢�$M7��s��YL�h� h"��K_c޼e:����#��C�	t�=��!R�:ٻ�T`�e#\�,`���ؕ�R��)��5���0�n�9KE�K2Qv`�(��9r���:l-��l�:Zg��T��CP�%,��j\i) �"��Q�4�l�� �E&M}$��t�i��.���ǓI^ef��|�<�|��,���'��V	�
�&��JمBa0�MV��a0�0�k>Y�|�O�)��|�}i'�����'^Y�i�ɩ<�$�̬��(��[�y#�y<�ד����q���V�KY<O'���yo�-�k|���O-�>|�y՚yl�����%�yo2��-��]+�t�.��Z���ȘI$�D�$G��%�i��y+ɴ�M��������2�O#���x�T°ᚘV	XN0�J(�C
�a�50�'+	�Raa�mf�[H�]<�#�$�Iyh�9ie�H�H�#(�y+Ʉy��,�2�#,�5���׾��˄�)���J��
8�i�(�cL]����d��͐Z�*�.i��0�l��j�b���P年G�G��Ī�(2�%��P���G��&0y[CR`����������=�&Q���Y�M��xúKo���
Hm���z03x������١��$�f�v���c�ʋw��O7�qƗ�{#�" �s��V�L)!J�г�k�Y�]u�JU�"J��6	y�	TI�T"��ʕz��^�[N�xNx���2��rami�k�X�p�V��] L���4����W@G�+�k2�����FH:�@NR�F�mGUQ<rw�֙��V����X�	����~g�~g�&fe�{�f8fk333:�339��y���U^,W3�w������ffqb�r��31��8x�y�u��p��Ͱ�t۳6A=u���:ę�j�ì�J;BQ��u�^3�\��Vf�s���Kh��K4�i�ʛ�(ږK����=F�r��yٵH䬶�١3��l����n��G&[��6f�ױkf�%���3]Z1,�U�;l��A�Η�Ҿڪ[��X��pݜ,�5ش�Mi�t�$ɬ!ll����m�.�A�d�9�e�2Ҙ�en����&���)-�̙-��+_De�����D5�5�.�Q�&�,�L�$RI��>�J�SR��4
;M�
KYԘ-eiy�����rU�]b��B�锈g-U�zq��.���Ċ��)�Պ�Ij�U�b��2���iU�_�K��x��o#i���N�Lgݕ^&���&�)�-��ĬʩnN��7$m���C�!)�Ф�(4�벷j7�m��!�?{�gӈ����q(�L��92a-�i&C�ܐ8@�E�f�ۻˮ�m7M�d��d��/jX�7�k#�4��3#>D�
�K^�����+����/˸^I�0x���+i��t차��KI�6��ŗ���
"|B�>>>q��u��p��Ͱ۞�f%�/ҰZOB$�	�>�m��hX����-:�i-m)kM$ϰQ��0ĳ��UG��L�;���ET�UTu�iт�HjĉII���Y2����iz�=��->l��L
�Ii�	i�i&J������k�ڵ��)L��f�,}�]UP���-�9�ݶ��Y���N$bM�m-�ݥ%(�T.��a��Q���Ym����:M�, n'pY�\Ja@Q�6e0Bѭ�o�%a1��ׇ�y$�S(M�q�[|��^q�]m�8��������(�J��� �1D6��6�m�����<[�"S�J��_��a2h�-.�ҩ�v}�M;x%�=L�jN��|�锤��F)i�|c̗m0�W�.�@�䇆����b1hև��H?b��<��dG��^���i9M9H�g[l��.\����tINIL����j���rVJKag��
�]7�d�즈�Rm#�*QTV�`�M����bgrYn1
#�-IW��e��iV�8���Ϝy�:�F�0|0A�~�4$��ND��UUUUT@<�e�rx�[�?)����!���F��0�RF�}�)�fA(�_��k.�:b�]��ŏ��pZQT�PF!��6t��~�	D�.�RS�E��,�m�ĵ��h��lz�O0�N�8O�)���L'��CP���%n�!U(�m�Ô�c�;>--a�|HBl�t�"D�fI!��ܬ"��.�*�������k�)�)�(�8�y��Xci)�nR�%�i��8�ϟ<�:�n�q�m�+��)��űV���� ��^C�%��ʑz��-���%I
VJ�-V��Ӽכm��B[�o���yQ�ټ�����gH��.zfZ������e��7�����;����뱵�31�>d�����5�=eݖz�%�i&�a�mS��e�Ѻ%0�F22e�L�ؖ�|�׋�lۦi#�RBB~��<�ǜ,J� ��H\O㭦W�jf�p�5���$DE^�D�Vh�� p�f��e-�g����$R��'ړFG/��[E`x��Y:��e�/H����}S��]�U�(���ϣ�*��FYuU%B����Y�Wu�gI�]�b�F�r��ch�Yv_<��q�μ�ͺ������i��Ci�uuec�I*�)���|D�dؓ���Hu0�Aă�a�0wm$�ޞ��&��S?I�0���S-��.b��f)a(��G�KL�L�\Q�<U�V3Oa#Eѣ�˽��q�������$���;��p�|�2l�ѓAc�u�a��/L�i5���-Ft�(�rHJ�ԙ>q1�ŝ<q��<��^y��p��K��_��V9I4FZI$�@�>�q��!����t����K�[7F̗���Ix��,�m(
���_b���]YñT,���Q��v� [��S�5��C�X��d�J,�Ao�XhF-$�0j!�y��-��p�䣀]84`�-!�t�����^���
 i��!*��(�����Q�V�a�rm�Z�ϱ�{�N��/�|ێ���<��qiw��H��q�����.�|p��  �Hw̏�ԑ!��hgl�b�X�i��a ۨ�|�i�NB���m�#01e��/Ma5�!��؞0`f�'z��FZ�,��C������D�g9JY��O.�"V)~]lS���Z�$j�!�]T�(��ܸ��8�.�2J��V��l��\�Y����^�S�>e��uכy�μ�ͼ����y���#���V�7�'C�"Bȫhr�£m"O��  !:�,�|�ŏk~ܦ�`�Pu��=�k����/rΓ��yP���)I%��+��e3�7�.��ɒ�`�cz�J�\�*���="RT�M�-)d�)�'�O��S�]��|��7�,�|CAoԘ�MT�s[>n�8r^$�~�|ޓ�/�g8���N�����%,v;%X-��˟�qmk��b38��n�d'�� ���Ŀ�
oOJ(����ԔN$>K�A# ����G��Z��Ke��,%e���q��,!��ǉ�s�ۥ�h�o<��ͺ��<�o8q���}W~��$�!
����)!Q���ĒI$�=�D����
xС@ȯ��o��!?�{4��\��$�H(ȶ�@�sYʾ��=Eą�C�K]���vִf�5)/VE����H�M F�������D$�X}�2�!��aN���F��O��t!�p*0�m/+�t� ���oi�|�G��>ygά�<��"aI&(L+��	�'�-I疻�y<��'����{ih�O"��y���L����yղ��u�$��|���>Y�K2�&S)�0�'�-�֗y'���^W�I��D�ʘVD�a0ᚘQ���
�$��%Q°�F(�����1'��y{H�.�.��'�Yg���I$�Dy�<�O'�|���q4��8�%mş#K,�e>FQ*(�0�L3S
�aⰘ50�TM�T0�2�хa:NV�T�1<����f�[H�]=Rzҥx�DG�#�y;%��G�aE���a+�-Xyg���V<�yM���~O�{2�2\��Th���3��Ԩɬ:��r�vAٛ�3;4^�L�"=�ط�L�R�E�V`w5Usa�Z��+�UV�S�t�
2��X�t�HZ�=Y�uzbF�F����:�˪W۲�$�c��3Z�v�)2�����3P�e�+|o�BB)?;������������~qb��.��3��ffg�o9wy����W�ҷ������ګjҷ�����x��Ǐ:x��:a���8h���UUUUT@潂�5tYD?%*?4FÉ�^�c#4�Z���UQ�)Q�%F���/k��eu��K5]m���q����_��i-$�u��ӽ^�.�e��%"ݬ�,�I,�Ĭn�A�5�����;Y�#����X�������e�J�쵒ץ�v��0�d�#�VW�/^]��u��6�ϝy�yÎ#m.���ֶul�gV4ؔL��M�6�m����U/�\�z�KN�4YA����o	�F�T�c�ŢE�%�}��B�U'�7K��ޞ�2Y�.�Z��RO��c�,!�s�ۗNt`�����7E>tᖩ���冀��ILv��,.@����nM��)2P|��,�z�J��\M�w��2w)��K|{�n�����iǞu�q�8�ŵ ��tA����&@3N(�<�qT|B�0�J^�?V��}څZ�,ZA���iB��E&�����$�I @����k��E�����J��*�mV���6��ޫ:mf��
��V�4E��<̑e�n��W+�++�������V����e-����He7�z���һ��㷌�6�=jb��kD���ّ&��VحUw��tޘ=O��G/i/��ܚ�0�9M/9IM{z�I������V�>��N��^����1Y>M��������m��s�@��r��X�ǚ�Bղ���h�̸�6��y�q�N��4�i�iR֥-"ٜ����� R`��'�&��}���{)�rJ�p��Z4��J�d>p�ÓYL��=N�M�_I;�I��[��D2n��L=�p��`"h����s�s���k����n#lm�4��F�22�`Q����Q^9f���?Q�$kD%%L&[�u��p�.��m��n<�<��<8�a�����{�j��L�Xt�UUUU1jUJ���x����	��e&�e�e#f4Ya��|��e��rI2�t��N`��F�07��$rE?0Un8���U��ė�����v����!I�����i4a�C���I�)��O���U�<�a��1k�Bkx�Q)�7S�H9#{�մ��1^�0�94ei�˟D������|�Y]ǝ|ۯ�8��<�Ν^B�ڋo=c�#1o~m��m	ޔl��	��74`��AٌQ�	I�� �z��K��m�}R�.��}�x l|--�e�N�S��|�s���d
x[2����FBf�-�1e�=S_W̖[!
��O��f�m0�:5�)vV�+m�0��=���:,JJ�l�XZ���2㬶ۯ�m�:��x�Hx��w�̻���\������9�B�,ĝ0�PN��z���_h��Hڲ��~>� 	v�DY7�Ha}V�N��J���#p��n��{)��S�T��\���VT9����2��+��wht�`����w)��>&���[�l�����!)*�Lq��if��m2�/t�颃α&8s?xo��c�vk9%�B�=�{<"h�lbi8����Zd,��Ř>�'ۓI����_��U���=t�Y��|�D��T��Q]��]�![p�__��RI�c$_���S�_�R1-kM���ζ���u�^u�y似�յ<��`�cS�"o;��UUUU2Ӥ�g
04�着��^�iNMk�c&���Q*BT��șHl�/�D�F&�����Ӯ]��Ż8đ++���5L�YX�����v1Q���� ����������홗�^��E��a5���k�P|���������%��0s;��|�8�N��o<�:�<�Νu,0�	i��bH���I$�@��cc����B���-Ԣ޿9�«�s=�3X۬R"��V��ƛ�����/���/~��]�.-�}��}kn��T*�8z�B�����2e���!iJLN�l�!��-1gϼ��I4L�"�0�s�kE��9��mpu4�*�R�B���8~:���ϟ�^u�p��+��-�m��<�)wUԈ��.�8<Z5�h�I��%���m��Ƅ��i�b1�<�q��Ɇ��ad&�=w3*س��"=O�kZz���\��2��%
T�a�{�4x�Hq�&�ɚb��nr�wk�E���3L��<#�SBh[�?3����ܻ>�%SŴ]-S��K�,�it�2��.�yuѵ��1L#u�m�e�n�Qt�kR���N-]eg�\M�ά��uo!��
Ha0�BaX%`��L'�-[�%��io'�Y��i0��C
+a6L&Ʉ�$�+Dyyn�O,y5'��<�)��a0�I�	3S
хa0�eOh�$��5�*}�a0�0��S�0�	XC+�8aE�Wl¸L9RYf̓�t��������Id'ȏ�.��I'��D�����]ż��[i��'�iŞF���e�����y#�u>_��|���<��zӋa�a0�50�,�&æjl�"aFRy՜mmI�FR��<G�^�#��<�<�:�J��=%�zL-�2���yO#̬�W�i�����>N�e�Uي�B]:�NI�^'A��R6�,)�$P�Wb��U�m�b�O24�Q������v�%��w6A��FfϦ=���BHϨA�e��P�&&58As]�3��#*��[�Ү���7g{wǖ�6+��U��:���S��B[�6�
��� ����J��S��>6Ɗ0Eo�W�m�����wq��}o�mݸ'U���b-L�)��J����}�bC��b�ug�m����z�M�P֛^��,Gb�X%!��hx����f�R��������*Ą]�I(�Sg���k�����-F����r��rK���a�ҳ�mZV�9wy����Vեn���331ګj�[���fff;UmWKw�������m��N6��:�o<�Eť��ֹ[_D�\��F���9djk��q��n(�;j�Ii���6��V���SF� 9�m���[�e����OB�:���BP�te�5-vqp��M�'�-�2�SZ^v��n��ĩF>u�b���]c���h�қa��6�\]sn�!�y���Cб��Em����ƴ�ff�R����Z�/mP���ji�3+hhö��LD�����g*���ji��%�ɱ.��w�������asu�M�lk���`���*oC(iwZS}}�  9/��	���Ӥ4�G)TC�*5x�kU���������N��so\4.ۼ��I;:��+U�5���å@ہzq�]N������КMHS"}��-�Y��������d�'ݼ\�'JJ8C]oRL$1AD6a�΍&y�]�'�h���WSl��������3\i8[D!t�����%S��X����>����W>rUZ�N��e^���.��J ��O75u�,MXBG�'ƞ;>r�8Y����6㯝y�qÎ#l��\��{k�#�1h�]���m�B�6�����]�n��j���ujY�����Ի4�d�w=��'b�<�͎R'ɱ�6�]��-�a�6�ȶ�RaqX���~��qAq_���䲶�vU:6���l�$B�z���	�z�t�հ�2�]��a�a�VX�R��fI��8��Y�����a4l��|ӭ��μ�8���WL���!��o|m��xн�ŬZ_��M'u%!�e��x͖d�@�-&2D��|�r�����%|�&���};ʔ���p��Nb�U�P&��#�����u&E�e���+է�#Fѿ6�v��}%�F�`���Sp�x�/b�)���e$�p�Č�O�@�p�~H��Yuw�i��u�^yǜp��+���І��cAm��xЦ5���1��Ʃ��:��۴��m�RU�ŷUsA=!�h�V�կ��������]�T)@�(��DP�?�G��x_�"�+N�-��|�m�E]�j���G�f\���!���g4�),�:���:�d�#��u�͸�μ�8��`��ߒ�6�UYaܴ�Ʊ��vUQ�"N'���vREIt.*��e	A�))b���֧|�m��w����W�}u��gVT��ov��y���K2��s(�u��^���1�+X�2�(]o��r;�D������F�C�pq3�2�L��>1$(v�!�����p#�#Ie�M's��S���(�S(�|Ӵ̞����^���p�	�ٶ����5[}ԒKS���S�w���H�"1��c�~�"�R��A�>��H�bU��`��	�I�4[��2	F_٣��]�*H�q�LƻY���02�>m�[|��^y�p���ŵHM?@k�N����m���^�a�]�0�Oy[����#�.�R-6�a�+�0{+�/	�N��]qs.�v�5NU��N��|qe�ŭ���kIb�O�l��t�,�0D�����}d���T������W]Wc�u�zj�W�>]�ь����/y�}X�o,�����S=��|�θ�n��מy�8�6��ZN�X��@�A�I��I%�ݩ�%#-���MۓܓId>>(�TQ���_����_:4&M�e�4�4|��߽��'�Ql��X�����v�`��q>h�|�|�Z`����GH��:��(�<RZY�%��3���6���� R��P��hgv����Әl9�!$��-4BP#�����B�2c������y�i��6��y�qÎ#m.�/{%Қ�؜̟  Ͻ�v�w$#�i��UWgMY��*�+x��L�r@s+y~�&���.☚[B�N�5G�n�`٨�'9�^�d#�����&���#gΈ��Ӹl����C$�D���$�)��ŉ>5�0�$���D0�l!i�Yn$��1��H�ju7��6��ϝy�N:�μ��F��A,1]+�9Wh���j�Ӆ�H�d����(�Lٹe�)�'H���
D"f���$�Iy�+_7��S�dc1����v�m��a/tVC%�gn�w�7� ̹�^��RG7�.Ul�-�n]䛈n�yn�ibf
�b�Ooܕ��Y���7��a�D���:��ݙ��;m��Y5f
>/%��w�G�p�#vQe�B|��H�I�ˣ��]]XDx,���ͦ�B�%�Q�:>2֍CE����|N/�����	3=c*��y��`�u�U�	�pR�c�TCV��x�.�+���q�μ�8��S\[Q4�����J�Ȃ^�sd�������Oo� ���ڳ��rD�c))���C.a"J6^����nH�`����	����0�9
-�Q�4X0G��M�Bt6ybI�TEQW��#O*�#=�
�& ش�ڤM�8Cd.��1�V�R�}�!��moRe+)�YtÏ�u�o>y�\'��<"Q��x��B��(N�f� ��b"tAO"lM	�6hMAH�����8P��X���"'Kı6&�2t�blJ,�2|!�O�A(O	ӆ��m�^Y�^]8ӏ<��<�o<tЂ$b"pD�b"'�8X�l�AC�A(�JblM��'�	����5������hYc�Jсm*�-�=�{���u�Y����ЊӞ���D���kw��^ߥ�Q>N
2����$!��egjNr��dpy3Y��4.�����Y��	)1�Zvw�`>cV�W����N�/(�γ�����M�nZo�7�����sj�[�˼��31�]��n�.�333Uڮ����3331�]��n�9y�vt�ÇN�0�	�	�ǎ�F�nI7�UUUUSD5�~˟� _~����Hc=��-�^�[���.����b�Y_�V����,� �Q��hP#�9���$���h{��ץ4�8��ƉJ�}��\j������G��r�nm��_9�)FFu,��;NrL���N�5F���_q�>i�O�|�<�N8�8�m.�#3��)$��Ū��Js7��m�����~�pı�z��G��Zq,1����!���~�|&�H�滋�����6B$$0XQM��IG��!
n|x7�\��y8u��Qf誮�a2��+��ͯ߮ ������ϒ���6�뼛!��վ��T��j�}�ݔE}O�mN.�=\a��>i��>u�i�Gm������z�bi�w*��T���������5P��@�#q�H�<Z)]���I$��״
��c����r�ӗ3/z�������ra�	��v���r�]��y�'pҎ�:��.�1�%�"f1W��e�ȶeh�f`|�7&�I�Ig$j��Ud�)�h�˾0C�2f���r���[�>|Ө�g*4��P�u�Eї^�Or7^f��5$�{?�k���D=�k���GIUO�Y
<����,�e�2���Z�m�8�h��9K������͢��nqw�aj�k���V�����'�^��/�#UZE��t��i.��6��|�ϝ|��:ˎ8�,�K��Z/k9�^�ҥb�:�m��
f��Ƽر 8��Č!["�&0>x�,�#�l�����K>2d���C�Դ����5N���+�L]��O�e�3\�.U�
&C�Pg�����_?��i�m��H�Z۵L�-l��}�w��!k��!�B�r�<[ΰ��q�μ���ʹ��f �Z4/�-=7��Q4ex�$�Iy-�����g�_�܋�/�4�m8���4�%}��n-1�N#�;k$O��%�������ƈC�g+_�(+!j�.�uk�;�X�C��(�2b�Wܒ�!a���2M:�x�d����F\���$dթ*ȋW�BG���1��>�^�J�̸ӯ�h���a�Y�ǈx���#$���x��|�m��o�U�Z�зȕ�Uj��ꘔHu�U�,�؍&��#���.�-I0֕R�T�ޱ����r~���e���CƊ!�L\��䐓4����VK!m�4��U2攰[B��\��ut�UG����.V٫�՘G��1Wmיu�qמu�e�Gm��öz�d2��)5A!*�K�-R���#�.-�<��\1���CT�ejI$��Gr��7
��1}�]�O�a�'nuǇ2������i�fĕ�iѲS��Ppm�a/x�iA�8N��d��E#�"�9E������\�U
x���!�?>v�i��$�SQ�ej�6��1W�Sh����B��)wA$&����yϤm��<pY�O@�4C�E�Ql�t�D*QE�Ԩ��Ӊӏ��F�l�9f��7_I��O�4��^u�4h#B,1���iڣjJ�P���wͶ�o1kv�Q
���s�gw*�%��(���,���$>�BS�'���D8���S�2�Z,��~3��֊�:�6���ԏx�4���{_�*Z0D�>��M[]hϹ��#�S���+Y�4�n���,JKk�{�2���XEG�5!W�ߴ�u�q��q��^y�q�qf�]%�6��i�kZ��o|m��xљ�_�(��So��!�Hg	��!4�}}MXl�2D)a�}�7-��Em�����ҌoKx��!~��q)�-$�mϜ[#�Z���~�q)1Жz�Y��G�SM$p�2V��HT)�x��pg�&�u�u�ϝy�\e�śiv;_m�b^��H&��ӉQ�)B�MI$�^@�� �� �~�V���:
2e�I7���'ѽ�(���b�If�I'�v��/��}�pk���>����D����!�$���8�m�#N��NnKZ�����Z�\p�=h����	eӶE�Z^�֚��m�Ϟi�|��<'D�<tN�8hD��M���:D�&�M�����,M	���	�""hDD��B�D�P���"pK�؛f���4pM(��!eO�A(O��Xm�_2��#�y��u�^x�x�!�lDN��"x�	bY��AAD��M���'��Řz�9;�}��_�$̿��AؑBFLu>Q�H����;N�u���
������):ޖ:��5�p�I)U�J�`�6�v/9s�g��U�bjˬ�f�E,�z�uK[���vQ����C��(#�[�L��l���@���W���=�����u����>�-�C�0芶�
m�ю� Mx�ƨe����L|�m��9:鎼SkN�=��&r�a��ڏr�#X���T!v�uob��B��A �@��X�0�)3��J�K�#�i{�k��*ke�gXm�0��Fi�������R�)�[������J��ϮV��SZ@�`�㉠�t��U�V���mL�k�n_9�:Uv����fffc�t�������Ǌ�U�ww������ҫ�������e��i��y�u�q�GS\[S>���P�F����Hʝi�*�p�êfK6���ͫ5�vܑ�95s���ʓR�l)P�6�ԛ.���v��M2�[sy�d��ش�՚j ؋��z�^��l��;F4��4+-�L9�kmk�����RsV�k#s^��ЍfCEcI�U������b��hE\�j.*X�iwCLY����u�5qF5-E�Cc�n��]�k�����vN̡P��f�-��a��e4�5"��\ʛ%]e%&� L��oI$��"�$~�@��ua����������F����aĮ����Z�4f�z�Ƌ[f�3V��ؐb����ۺ�Tdem�-��z��]޹�c:�Q�q� N ��4x�Ѷ���d.�6��	6m�?`�R�Ԕ�`�!c�G>��C�B�	�zl������C���T)0R�����+�����@ݶ������\�/!XlB��6�l�_���>x��/_��4]ܲ�`�'�u�|��u�qY���)�Y�L�I����b��MN��n���>0S��̐�G�t�0��-V�UW�1���`�bםw'�Т�o�s��Z
!�ѕ�:�n�[9RY�����rV-B�o;ٚ��)�R<]U������~�^���KvN>-����}��Z���V��[+��R�k�ï�|�o�8��m�Gm�ܴ[s�K�׍���h��srT��I���ӉcÉv��pf�,�nNJ^��"9������ #�ļ�E�6�IUTQ+�g>0Qd2�L�8E���g��ӭ��$>t�h��&��>��0��}ۛ��mV��������L��m6k���&AK���|`����:��8��:��8�,�K������W%�࣐AjjI$��@�����>�#|�����֭��Z�lӹf�X`��	�M����!�4�˷A�iM�4v�}��g���+߽�Phl��LƜN�B��q�N�dӣ��xZ�y���԰��>;[��i�v�G4��C�ד��k��ϝm�_8��:��8�,����Rd����a�MGw$�RS�U����I��.ͥm�Ĕ��u�f
�Q}6�m�Mn��{ݚ��v�*u3?�ޗ*��ʺ��]L��w������q������}دz�V2.$�t�Z�+x��﨎���uY�.�+�T�6�\o^]6^R�W�m/��%1��Q�ׯ$��Z�}��m%Y�|�VK�|-;KW��svjɒT*�'�<y�|XYf�4=0}��Y�����kƟ`),��c�b�˵	b���UT�%RԳ^�<��}��ao�}(!�HIt�FM��V�
�K�㏙q��u�^y��q�]MqmL�)� J�l1X�!S��I%���~����>;ZĀti�2�=L�H�h�|�z/i{�8�7�y�Y,�)� r_KHv��OHI!5���w߷R���)8k���`�����U5T���U��9��!�O��]t.�vj��0�&��%��/%�y)�݅�Q�ΰ�͝<&'M<C�8h��2��
���hM��|�@ �����V�TQt�9���I��ߋv��|&�E�k+Y$�BO���:��]욾)���Ai���!��A��8�ߑ{N�f���i>\0�:�LW�B�1ԛ��k�at(��}]���]�i,�s+�RU�;�1�҈�&���Y�_<���u�q��:��8�0Xa[�"A"�m7^x�I$�,�.}wk4��ST�wd0�[	��0����ª5r�&	6���ԑ$#io�ʬs����V[O�q�ـ�GNS������6Rc��*%Tte{n�����C�D�Ӵ�4b��[�����y����=v�q�Ϝm��:��[]�śXc3�?q�i��nj�h9�7]LƯi����S�[�a�Ǫ|>����m���3�I%���i�Ls[3����%q�Spk�][�����zovV:ʗ)�U������ݱU�uD���z�����h(���X�SIC"��=� ��4�i��\��ˮ�
\�-%���{&L1�$��׼�*�d�b�p��pUUJ�s%�O��S����i������V\���{������8�D<�� �B���!����ٶR�����E�%��g�4��i��y�y�[]�śiv�c�9בm�33�ME�6�n�(4��g�~66���0��8�O�
X2���R�D�r0��`�3P��Y�m/	�����K�$*VL-�UK;H�r��0�Գ�rI�ˉ~$��E���Q�i1i_J.�����1���{��_!�2����}�HC)��8Y��{�Ξ?��<'���xDD��:YB$ �8"tЂhDК,N���pM�ĳf�	�""hDD��B�DM��GO�ӥ�bX�f�ДxN�4h��!eO�A(O<Q�4t�6af��a��t�H&afa�<a�<p�ĳE � ��E	�DЖlN��4`���:��Oj��!K��!{�2�>
>�ST3Z�ً���\�\���QjM��癚�a����V�5�n���Sh�6�Y�&�%oc��ʇ	EϖU�3��I��Qe���r[?ROQ�3�
�$�PP)�}��Y/wsw?|�V���33333�*����fffff=ZU[��������z���wwnfY��i��y��qמu��q[rmE�  ��o�H�G��m&/�M�F�na�(�=I���fͦϽ'$'���m�iѶ�sZ��WUu�xQl�Rm
��4����J���c��V�O%4i3��>�3��&JL:	�ܕ%J�Vx��$�Y���=�C��<��m�:��[]�ŷ&�NXėL�6C�kMd�@bl��&%X�J�~m��x�ٵ�Q��N'L'��l2u�ɀƌ��N�YT��V�k��l�M���.��Fz�;�od��b�l�Wb�0���9�1�O9-�i4m�$&����]��F�M��ȫ������c�,OBh��o����Pܳ�0�O6��:���y�^y��q�qmɥ�Lu�.�F��1RO0PR�GU�)⊔�&4�]q��R�&,�gRI$����-��<wꪾ%JŨ�j�pѻAltֺ�����"�m���C� 1�Yρn��
�8�B��J]->�>�9�[RHe�|`���0�7�iÜ\K9�Ai�v�*2��fS��*��Y��S����r�qf�J�a`d�<���BJjZ���)�
X;qyi��B���jJv�]f��mw�4����ǈx���C�e2	
ޢ�y(�DL�U�|�m��{������,��W�f�<��Ɋ�S��l�7Aݞ��LX[���<Q��&O&h�-�}��$Z&+�(�������.�H�6�Y(&H�r��6��e�)9���詧f̶����j'�Sk�t�6ɵnn�}�vS��e��m�8��:��4�a6�U�<�4E2�$�Ix`|$��	�Ϥ���$�Ӄ�h��`3�+����@�f�s�h>�A��^&�->��`[����Ĥ�:�s�BN,{�_ չ%_�> gƮ5!UW��s����D�u|�>y��q��8�χh�F���c�Ɫ�E��RI*�JN�NC���������){��8�(��\SKx��W��Qs��=)��B�6[N��!����������C�=�y>6�Ӄ�խk�p�W�q���3N�+�gW����/SFO%O&;'���S��m�m�\uםmgGܚ^�G�o�6�Y�$�Ӑ�-�BTQ�os ��7uG�P�q�fԒI%�.u�O�U���2��� ��*FMl�1�5��pF�fv��)��e����V����x�E�L�۔rP�����9;D�<���5��ϚJF�1�t�x+����܀d��ɜ����94�2�n �Ū����m��=�#J�.oR88�bRP^HI=�wWX���K�;�$�gW�-�A *�mH���I&�I+ВD/��ph}^�n�/�<��>|㍾y�]q�h�u>�V�/�eEuM�r��n�-�T��L�HB)R���}��>bl9�#<��Ϥ�A�Y���8��۲֭S����;v~䵬�u\b�I�䆤��u�x���g���?xY��R��-^�v+m�R����X5{�d�I��˂�|7�a�{RBt�$����+�Kk��V��m�2����'8ۯ�u�mq[riv��/jIZ�CFje���Հ.�Ͷ�KÀ

Zj��n9�{�<3ߋ�������&�J>!�m���)��VC����`�هN���������sML�^J'��^����M�p�e2�=!�h=��r��3��x-��m[� ����o����57[u�!�Z�2�6�m��>Ѡ���Ж$���UUUT�D�0n�td��+�^���u/�<)��#�8�Sg�RN���s�0�#$��M��;	�Kl���c�Q*�R	�<�a�I�;n'��g��w�n���.k5���luW��2��t��	�<'��<tN�P��"lDN��'JD�&���btDD�blM��E|��2DD؈���"A6"'؞�t�blM�6P����>��!�DDJu�u��av�aיY㮣�<���p�H"&�DN��a�t��,�F �"%	�B&�Љӂ!���x�#��Tڶ3.�z>*�r�j�C���т5^r�\�z3��^#��9KD5������r���f��_V��*oQ�y�亷;�X/�{0�N��+�)_;�UD���`�hu�i�:M8�K�Tw�0�zE r��Ώ"�����Y�k�R�6��]�*8�٨%��+&^<Uf��,b�3��_i'�r��Gt�黶��z�H9�D�ňc�K���w*���=.�<���m�u���7�w�����	�r��rS҇�ۡ�AѪ�Y�2D	6 Z�t�6*���	�3��D�ʊ�edEt@�1�;��9��Yst2�S��I��^h�{�Ԫ�kg%~�������wwo�ffffc�*���ۙ��������wwnfffff>b���ݮe�8p�ӆy�uǛGG]�ߒ�z�;�^�v�eՖ8*䢃!����K+j�R�"XT�E��L�;�a���yB�fu��m������pź�k���l�ײi���}�V�l�I������u6%T%��l�Cb-m��aģM�V\Cb˺��-:#��-#-��d�.�ڐ�հk��5Ƽ�-��]5�\�s���VR�;JӶ0+d� �
�t��L�HM-��7!�5�)i5+%a��Ʃ�+��`�mHh�sV`�.��bƺ��Z�=m���M3bO=y܌[��S\���y��պ��Bhfd�m�u|�I$�3�,"h���Zұڒ�\��&]�b4X��cvo*P�wx�9;L�CYl��f�[�q����f^:p]��V�`�R�
�-'X��T%n���-Rg�HI2��`�V	ʓ�� Q�-�}�I�+~�t7�-���k�,^���_9Xwɽ$��x1w�q���k�8�=$���ÓA�	Y2j�����}��%˲�YD�}�bc޵tcZֵ��v�M�`v�T�~`ʕ!e	g���<tD�4|0�A01cWe)L��|�U�/��֒JYfi�L�.��G�
#�;�pP�~?�m��X ah���y�i�	�fS���>3��D�t�n&�Sಃ�5h��l��#?m7	+Z����͖���6�4@ƒ��j��$'�p�pN�B�=�~	F<'L�'�:�A01c{�e�^IB�8�TO@�ڭ��[mt*"�~ǘ/�<$)ϛ��v���$M��f�G������0\�YA�{����U�Q�/��0|;بX�X~Ӌ��0���$HzN��+�4�n�\}���$����(��<�����-�ߊ(��~�	��N0N��<a�F�h�ņ��I��a��Vd�Sl��u�aR���I7O��5����$J&6	��UUU*U$���0��'\�C�n}�if���80sAIa�'��A����Y��0��f6�srJ��Yi-mR3[|���bŢE����ۀ�n*K	��nN�R��{2r�]�y��m�\u�h�F�X�o��+J@��˻�iZ-7q׶�����=���h��0T@#)*K�$��޽���Un���(N�0�%obf_qJ�]�r��6(>��ח��qHy�An�5i.ߐf�'F�;q�=��]j��Q4�Fz���Ԣ��0W�P��~�5#t�����1W�c��\���,���OS�$���]�h��f`������H���<HΦ�d��&Set�����A�`�z��jC����(��b���:ۯ8��\u�ဍс��h\�RS�U�d� k=���Şx�),:�w�=���@��	~��UUĢ�x�.a����}ºCN��f�*a�����PG�߁I;ҢuR��G���U$*�0�	fh��G�p�v�5��|�/�<x�:`�0O�0�WP�������W��E����7o �`��<Z�;�/}�G5���&��c�Rm�\�̕XN%2Ĥ�l+2k�=K6��b���x��^-�R:�L�Ez`s^�ǝ�դ�ڪ(��d�u�����w�Wn��KSk�]Yq��*SX��d��i�����n���Ͷ뮼�o:㮸�h�4`b��Z��E�$�#kx�I��/�=�;f}��w�M�����!����K�Fq�����ڙ����h$�ΰѧF�I��Y����i�.���Ѷ����dɼB�%�P]Y5�U=8l6g�n�����J�H�����r�]ID��J��n@�{k��M�����,��8�n��8p���F�h�ŋDu=.��UڦV�%�TeI�hǑ勶�O ��oOhw�P��2j���!9� �O���[�-�j�3脭ͫ�m��;�n����V��;g/GCiXy�_J�oX�n���A�о��]�CW/v���5�"#
{���w�| �05;;��~��>z�4Px�l#�h��p /)w���)���ڞb֤�`��)�>s�=�5]J�\V\>��#��)��J���I'2��p񔰴�絮R�0}������n:�Ϝm�\u�x��k�����������{� �1uD��ךK|���Pb��mPI�=G���zxA�b��km,Ƶ��>�T�R8^�iV0�J9f�F2}�ZR�|�{���E^���h/-0��Or|DN��$>��J�T��V��V]ƓF	!���t�>N���
s��I����bx��xO	�<'�DO��"%� �$4""p�'�D�&�؛f�D�"%����"A6"'O	���%�blM�BQ��A�	%�DGRX�'؆�	�
��a�a�'��B�B"X���'���8CQ�����"ABh�"lM�tD����S�'��2���}^Q�� ��"T�k-�<i*UAK�(XA�~�-��-��4Uj� ��p���E�YEmU6�"��Z����6JiAm��t�x�M��̽�S��f�d�r�d���"�C]ͱ-�ز�j>��YX��{��J;�ͧj+I�3�vn��Zt�Rq]�5Gt�[k�M������
Zi=<��_�۬�OM����a^��_dU[���������1Un���33333U[���������V���\����m�m�\u�x��k��ԔI$�}������_տ� (g��s��_��hav`��^:�4@�}�(���%Q(2�~L��M[��I��A�I�ܙs���rL��4;�`?�;`��g&�r �E	L�CO4s��t4y�S�	t��>y��u�]q��8�6�Ov��w�k;���NױE8C���bҙi!yD��-.��)�K��m�Ш�C����e��!��an�Jtiѷ��.K�1�R�]�q��S��sf/���CpR4�ӈ�J���1sY�|�nӦ�@�y{g���e��!Õ+��^�^��z�]��e��m�\u�x��k�\�=�a��{kUW/��\����J=}=��J�t�nWR���K�� �L_
�+ﲾ��T��]�ɭT�$A�]�A?V��E��j݄�U��@�rv�U�P��=+*���Ь��TM#J;ffS���2�%��Ej��q�[�%���Gޕ�n�����t�H��e�n�&�XwRHI4��>����M��Τ�1Z�п���M�"n��v:�������N��m�M��Z�n��V.��If�Yaa�%���g�<ۭ�뎺�Oqmv���z��B[1�Ff.9qd���kx�C��;��Tzki��=�����	$�Uf�]Um������H����v|d��W$�����}S�Vm��F���4����+ډ�I�3w�N���M�x��,M��V�pd�zW6�t�}*Uw�	_'S'�ۮ6ێ��o�q�\i����[���I��m����� g=��uUEs�X��c2CN��.Gɟ���XC��|�o��Dɑ@�զ���HA8-���� �K������2KM��$'u����O���nJ2m������;����8�i5Z�՚m��4��y��u�]h��4���m�$2�(w�i�� ʚ[F{0�\_���*q5Fe��2@Q����?ʨRN�v�����h��O��S��|Rn�%T��L�i6���l�j���\H����)��m�aZ^�ee��k+��&�디��Zj�^���h�ZV醯%�u�q��6��o�x�h�K��_��lB�)B�Xmz�T�� ��.ׅ�	���!Wr�\ ���)�I��FZ�w������L|��V�nE���^ZAO�}��sD%�'H̩p��Z�k�Uf��URn��QX�{.rJ55.f�SX��
��I����M�J�}ǚ��,���HY�N[8��K:�3���*��.��h�-�*�$�������u�Sӭ��s��h��l�� �]�<����?���Q�V���f��`��Ĝ�W�<H?��E��m�ԒH���]�e�m�:ۯmiv����fI$��-�G����J��Zt闏S��%���}v�I	V��÷��׻�[uĭ)�ǮB`�ĥ-(���0d�Ӎ�<>�t�t��eU�0zHH���Q��{ߍ�G�����i�<���Mj�=nfƪ�B3�B��V�;\]w�i��y�m׎6������tk���ZԊD���Ŋ�q;�$����8����8jhѪ/�]&ӰϹ۫�>&^��f�;��W����Ol��5c�<�L[B��M}��I'��Oɏ&��6|����|�����RQ�� �`�}�z�'���")�}�v��O:�θۇ0p��a��(bXۦ���$�S4�v��0h6��-�����)��a��ߡ ���+ݡz�y���}����ќ�[L�H��yم�5�iz}gһ�*�V8�to��^:(�2[��¥;ìnM����H@��>a�'�&_����c�����	�~�$�I 0ET�?������_�8`���PI��ᅲ��(� ". 
!��S3���Ja���]A�P�V��)	P��H��HJ�-K����P���P��"R�R�*"�*������D�aB 1�H�!aR��	HJ�U*�"TDJ�D�R"TDJ�D�J��� ���!��DJ��J��Q)�Q�)�H���H���E%DD��J��Q*")*"%DBTDJ�HT����H���IH�J���Q""R)	HJBR�"��UBTDJ�D�DJ�DJ�D�B%")�!hZ!�D�!�X$!*�""R!�*�"��"%TJD�DJ���QH��DD����U�H�U�*�"UDD�DRTB%")�Q)�Q*�R%""R""%"��*�"R!���DJ����D�J��JD"����D�a�!�.d"���%"R!
�	Q)�Q*!
�Q��D�B%BTR"�H��	H�RR"%TDDJ��B%"��*�""TDJDBR))"%""R"%E%"TD%""R"%DE%DD�"%BTJ�P��Q)�"� (�aD�!B�XF����DJDD������Q"""UD��QH�Q��"R"%E"%D����*���"TD%E"%B"TJD�DJ�B�DD�DJ��Q*)*"%""R!�IH��Q*"%D^���Q��*�"��*"%DD*!
��"T"%DE%DBTDJ��H��!`FaF��`D�`FHaD�D�����R"R�H���TDRR"$DJDD��Q��j��P�����������JDD���JBT!���X��B0�"DD!R�*"%DD�B%"��)�)	HT�`����`��!�E�D�B"%TDJ�D�R*!��D�!d*B���B�(�*��R��EAT,�X*���T�%�R�%P�
�PEQ��UAT��v���T���U%P�)PJUBM���K�D��
�!U� "�,+ �0� ����QPJ�A*�)*�� � ��B�JR	JAA
AP@�*�EJ"��AAA*��ARQ� � � �T�U���� J���J@�� �� �H% �%@�PD�����B	H"��"��!)�T�J�A**	IUhZT!R��JBUB!)�!*��HD%!J�!)�J�B�P�ABUB!)	U�D%T"�	P���!	U
�J�D%!�P�P�D%T*!)�!	P�%!�JB����D%!J�D%!P��!	HD �BUC5j���BR	UBR���BRJB!*�*�JB!*�Z�/X`D�`@�`0� E�`E���!R��%T"���P�JB�HJ!�P�J�B��%T*!)P�J�J�JBR���B�T"����"�HT��BR	P�JB!)�J�!(����%B!)�	PJ� ���D*T"��"�J�JB���*R��"	H%B!)
�,�)�JBT"�"�JA����B�!	HB	D%!�B�!)	P�%!�BR
�
��A*�"���T�J�BT"�)�BR�JBQBRBR��T�D%B!*���X�*�J�A*	P�PJ@��!*	P�% �T�!	P�J�A*	P��T"	H%B!*R*	�*R	P�	P��%!R�J@��JA)
��)��D% ����HH����i 1 ��-V*R	HT�A)R����H���JA)R	HT�% ��%T����*	PF	`��	���T����J�Rb�z�A*	PHJ�)�R	PJA*JA*	H%@��J�R�*	HTBUB ��R	HRT�J�R	P%!R����%@��T"��P%!xZ�JA*	P�JA�$K���"@c � #R�"��P������J���%BT����	HJ��DJ�JB!`FH`F�HF�B D�F	D�JDTB)	Q*%""R"�C�W�1��G#�k�b��JP�(N��W��b �`�I ���a�_�O����k�o�������������&q���=�%���~��,�)C��./�����i��6������j������N�g�'�����
d?���w�T~ *�?�/����������z�!�j ��@�����?�@��C�D�G��?������Hh��J�-�	�C��~g��w��?A��΀~��TU�������	 e+�6����"~�� ��(`b�؟�6���\JJO�M�� -4~�k|to�	����	5?,~�\�!�l`���m<o%?��P����j.`��6ش
 *����` � !Q����B6��}]�U���l�V���s���� ��@�P$AqA�`(+ B�� (+ B�K��������>����O��{�l���a��v�Ar�"��l��#�����W��ʄ�I�Zu-'�W�5��/�~��?�����~_����Wt����h������'���!����?��W��9�?$��g����QT������Y�|W�?i��zl���F����8'�?z������Պ�������%`~�P����S����ɴ��i�ʔ˕��$!��<~�@@������m"�
�U`i%%����"cBqr�#���a���.q�x'��U@i2������O�?vךTU���2'���)�_����,_���������E��?��i�?���u?p�0~�����'�����R
~��#�w���G�~By0�**��G��~M��VW��z�*����9�����s�������~���Z�{Gi �*��ϟ�92(0.|?���?���������v��τ�������߬2�����~c��0����?C�����a��1�?���~����O�B��YT�zx���)�O��O�EA?��?����vAO�?��t:O��qDO��0��?��)t~�jl��G�w�e?����y�J�H��������ܑN$�6@@