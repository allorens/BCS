BZh91AY&SY T��݆߀@q����� ����bF/�           �J� ���j��R!B�A$��6Ҋ������!�f֊SZ�i-j��ER��F��%"
m��(
��()At�6a$���$l�F���m��4 �U%6Ԩ-`�JV�Q C6UTR!�� �� 6p���U� ]��� 3WlI	��$
�$T�6��U�����k!U�F�EeZ5����(�6h���B���p nD(H�  �R� 
A����4�Imj�U1{��U��Ǖ����s#V�kb��kh���TVc�{{�4i�j��׻(���MQ�[Tj&��(�{��z::�h�==�ꧼz��@
3����{����ofR�K{g��XQJ���0�R�r�q�l�p�*�\z��PR�*n��%UJleDHU�C_<�  �`{�{JR���g�=��[η��R�Mǯ=ꊕ^=�ot������H����T �U��J
/m���
Q^�w�@z�UAsPjk�e@����W����|*T/��N���O{��:t4Н���:^q{��G�����T�à�AJ�� �omS��P�@Y9�U��B���m�)�%U��HD{��TU)��}�= �j���.(U4�E�Б�N�U+F�wN���v�հ4)��T�J���:�R�wZEUN�J�XR��W�@�;��Р��s��� ���S��S�J �7#u�d�q��^��Z�`��5B�I{��c�U�V�u�h
;�n GgUE+Z
�)�"�>JP �;> �Y����S� ��� 쎜  ������ ;�Xhh��  �;�hr*�]��hű�l�_>JH | /4
>�:���P M;�P
;�����S����@h��  c�ph w\��V�4Ȅ�Q��II_|�� {��  �_pzG�1�A�0�� �� �A���� ;ʺ�G8�
1%%�((�ƃ"J�JR 
�� k�(Ε� �� u��� �y���b�ànK  ��Y� ;�àx     �J   j`�JS5#�b =@B'�Ĥ���F���4ɦF����%*���      jxD�j�"`C��	�LL&���R�hUF�4h M  !6���12�SSi��&& f5M��O�g�?lD���?l7�x����/.\t�F5�>�������{.ek��U AAV"���P~�肠��h?����g����h��O��@_�
�$�;@@c��a�%QE��������~�)�Lŋl`�ض��$e�m�l؅�`��6��F�-�lKb�؅�-�l[aŶ�m�lKb�ض�,`�ŶlR��m�[#؅�b� �lض�)��J`��!lB�%�`��-�[�	lRإ�m��[�l[b�-��#ض�-��c��m�[ؖ�0m�[ؖ�-�lb�ضĶ0-�S��m�l[`ű�l`��-�m�[��b�[ض�-�lض��%1�0m�[��b� �$cl[b��-�m�l�LbŶ!l[`Ŷ-�K`��-�l��-�[�L[b� �-�m�l�1��@S�%�`���m�b[ضŶlb��4�`�ؖ���m�l`�ؖ�1�%�m�l�6���m�lK`������b[ض���m�lJalJb��lb��6����Ķ�m�l`�-�l#�6Ķ�m�[ض���m���L[`��1���!lK`�ؖ���-�m�lb���m�lK`�`�)l`�ضĶ!l[`���Ķl`��6Ķ-�-�li��i�lb�ؖ��%�m�l[`FĶ-�m�lK`�ضĶlK`��4�b��6Ķ�-�lKb��6Ŷ��1�l[b��6��-�`��6Ŷ[`Sض�-�l[`�ؖ��%�cm%�K`�ض��-�m�l`�ؖ���b� �l[b���`��F-�m�l[`�-�l[`�-�b�-���m�lZalR���K`6�-�[�[�؍�b�-�[bF-�b�-�[�)l�m���bŶ!l-�F�Kb�-�[��HŶ�m�l`�ؖĶ%�m�Ŷ(�T)��lb�[�� �P�*�� ��E����[b+lm�lb�lm�lb �`%����F�"�؊�b�lb�l �(`�[؂�Bآ��
�E�%0�0E�
�E� �-�lQm��l���b�lm�-� -�-�Q�"��F��m�����A� 6�Vب�[`�lEm�-��,b [[b+lAm�-����@� ��E� F �F�*�[` [[b�lm��� -�1�%�E��U�
�� �
��V؈� �(�� � � �P-��lEKb
[ i���)�-��
�E�*6�@� ��@�(SKb�S[`�[[`�lAm�-�� 1�[�(��"�-�-�E���[`�`��-�lb�ض��1�-0m�lB�6Ŷ-�m�[�[ �l��m�l[b����0b[؅�b� ��`�0b���-�Kb� �l
clZb���b��[0b� �lB�6�-�cl`��6��-�m�lKa��-�lb[�6����%0m�l`Ŷ-�-�`� �)l[`��6Ķl[a�-�l[b��%�m�la�Ŷ%�m�l`�ؖĶ1��m�lb[ؖ�-�lc�ضĶ-�m�l`����m�lb[�6Ŷ�m�lH�D�*>s��u����5G�{VYV�!�eYAP62�+��֖V(�*
7&��	�-��X�љ�)�^d;4\���X�OKo|N�`M9.��j�3]�#1l/%ޭie�z�����SwrG�C���$aQ;�����IZ� �z�Q1��ѯ+��\�2�5�1����!�o�)��.,,�7(#X�����豫qD(�T8���@�6)ǱP��)бE��k�mLґ��Hf#��,���6]�*.�ڧs˿C��^����[F�خ�+T,�+�a�Ų����	�F�r۳b���.�Qn+4ȶn�3ko]�����n��߮��tS�/%Q�jPn\�/�,5�:�,�z��&&Ʒ� mL�e�[�Ժ4�j�[�˗n��te�w��/!��ٳz,yoWn�p͔��th�2�n��琀؇1h�@n��l�r
U/)Y����/f���.[���̤�(��*�:�.�S�	mR��n�h��m ҕ��)�t)�1�j�lYTã+`W/ٕ�hX���~֕i�5��ŗ�74rŗ�zu�����n6���P�
���BՋ�Qh��PHj�wn�/E �G�nIS)AN�fnET�\�ƶ���\���ң�rP��-�7���җkD.��ê�S�S��{INf�3��j���6ud��o��$�b�
+]hn�d���<�����tc���F��o@j�(%�˻�+�m�P��YN�a\�Q<�"-;ʵ.�Cucd�P5���i�m�Lf\�Csb�5�BL[N7�TU��@靬ѱm�ԁݩ�rS�(N�Ǌ���966\���v3j]^���q$p�A�P�YL�U�gj��U��ϣ����˲1�+	;%V����&fb�Wt6v%��0��U��)�g[���0�1ݗV���S4���#Xd�)z�F7���e�h�ni�7�Q:N�'aWYT�rSB��f�tҡ�JQj��Ĵ^Q�5�Ջ�̭
z���U(/6J:љf��A�CX�ٱР�^��^���RXT���T���*`j�t7qF�lGc%��F�Gh ��8(�]�V�YU�T��i�)-@帄*J#0�M�î��V��R��nC*�
v�J1��,&�9*�f=�zz�a�]ٺ�,Pb�����Z!jPj82�c��!�6YrR������#�]��6�n��[f�(-�j���ה5m��@f�ײj"V��z�2I6e�4�l�v�ZSu2�u+o_�Z��f�j��ҀH0��[��pV̐QWr�z͟��x�݉7�l��xn��)��)�N�:YwP���zp��� 1�ܬ�%ڔ���3�݅aӹ[0d�72�7lFj���k�1�����Z�Ù�.��!���N�݌C1�tN��7�)�c+�f�w�2�Gs
1!�P�]��3hI�����Tubt�5dⲡZ�#�3�#���el9��Kn�����;�Jd�jļ*�(�1��]V�͌(�ˁH�c*PՈܬ�HV1qՁ(h����B���&SУ1��5	���&c�(���6�a�����B�%<�,�7��=���5-�q�Q�{�����PՀ93+LۣB\̎Qx���m'�Vk����=�A `+Szw"5��������:ȝӻPR�q�"K�e��.�m
�[W2�BYx��a"���K;6���
ʏ7L�ۑ����-�xH�Z�f]m
G@�Z`���(�I�ta�Ú��R$L��� �l����zB����%�SN���Rsi
����NMG��l-�L�GzJv���i�.L�@@ǀTl��L(�9y۶w1&	�u&��"y��n��i�u�C�4u�*�TՀ]���̤��ɦ��c�	dJ7t�&S8l:�a�c�,8�T3&��Ȣ���V-pG�F�7��ݶu�=hɖ��ڗ�Ӭ�u�q^Ayaz����'76���R����v����%�z�C%9W"��f(3nk�bҞջǚܓn���hӀ��ߔ�(T)�4v(�f*7bTXު[�氲�n�x�5�]���he�BA/ݚ��q̫A���8�-{�G��l��=�*lSU�v�ңK+R��I�ʫ�����B�����Վ��U�� ��Ø���a��n�sLv��@E�
\��

�1˭�)f�vv��ʳ#4����)�VK��$=Xu�F䡅[aUX���V��YN��Sj�'�6���n��x��T��'��tb��%Yt�g���b�T�V�"&\�B�R�j���FCzӔsj,*..�����%��[��^��I��WG�Gc�E���fފ�[�����+�l�)�ʩ4V�z��T�R�wnХ�i�A+ZUu7sD����Dܻ&�YJ��d��M�ǚ|i�u��ܽ!(�%��Eb���0W�5]؋VP��G7v(�X���:�X��ج;�n�qU�:�[$�	���f�(�j�)��&��p�K۹%��v�J�{wWPP��RY�&t���j��F�
�GKٺ\2�n�\���ںz����>zi�;B��w	�`�32,zT�i�r�\z^j����QH��\���+���3wR�ڇ#�v�d1#�O�5cK�[P�7*��X�s&f+c*����#m��F�Bx,�Y���vn�P���'sW���a�R�˺��Nyd�Z����J�bC����ŗ��c W�H=z��d��ö�kobouF*��'2M�u����障�Z����q��-�.M�UX ���fd�MF�h���*
	�D=$�ڶ�+ƨG0k��J�D�)�t�&����-����vR�,�ݗc	�f�j��7���*���2+̲�|t�r��FAl�\��3x�T�R���\܊�N�i7Z�ôF��ncϞA�QϪ\,�T^�Ke^�r^�Y�٧��L�2Ũf�Y�m���4��)�`���mQU��;Z؎:����8u��^5u��hY{�潲]6����$��h��X�Xթ�ò�`l���N�6ڷ!��o7	�̈́IbU�Vdz�3�×'�ՍEhH\�y�F�Z�5x�4�X�(m KFjڭ�(2��o�e�r���S
b�B�E�	�B�E�KH�cM���	�;a��M��B�
����*RY�d�˫�����u1��Q1u�J�X���kx��V�a�%�#4f���[Z��e�Q�Yk��&���2�h=6�i�ֳ����ۅ֘q1P�,S�hh75�:�ݠ�����V;brkkklL���T*-�ɐ��&�"[*92����ˊ�8q�0i��	�Wv���Ơ��{�Oi��=�ܖZ+*M�a�.�,�4]#4�#��%3�m�AAGsA*��l�/v�^h�hR�d�q�'.���hB�`"L�*�\��*��(���%������WR�u#V$RJCj�R��p[]hoa�(�SrZUI9N�YD����X�����¦��ob%M�v�MJ��^5E�(k�DV5��D�V��eZb&�"fl;1J�w ک�`�V4�*�Az6-�����m*��Vi�5�Pm���(Ř^};��	���J����aʗl8r�yf"$z�-p+����t;���X�d2�;������z2�l�K��s-d��2��˩Wv����[��y���yG�6�~��퇺[ �Ô��C�s%ź�x`V/lHJ;x��v�	��MsU�yn��]�`TZH���ATq\$�b0�����n*p�SVf����woCf��0ig�D�
ӭ*�شޠ��[�7��&����8����e������������{CRU�55�m�Ԗ�B����=l��SWAm��vj#%��AW��˙�f���q#�o������u�L3��,�*�N7r�t^���ZV'�4q̂+kE*�Z��9�5�N�����Ԭ�Vh"ȴ��5��	-cRncnD�c��Z��T��uv(��k�^=,�0<�4�)2k,z�FI5�ݻu�{^�0&���J��KuF|�T��dt��z��*���H0��3V3[Ov�XJ-f�Ǖz�.ȷ�ӧcq\D]զ)��q�+m�k �B+�*��9�d�Ul�n�i��h��k�����i�qN������j;���۠��Ǎ:7}�B,�!�	n�wН����K}�fM�T�c�C/M�7��m�lR�kr�(�����2R��_����lI��c�CZ��kh�q#Oo�ʍ����)7+F{�U!�-��n�SA/]�.�
rDt���5t��B;q!w�-��7n+؜`��vü�EL�`�u1M��I�cwm�Q�̓^�W�8�hWcQ��W.+&7��0��^ްq�UV$��.��j�{JaӐ87r��*C��݈���q�^cm�0TOxLF���L�ۺܖp�
�+/L��a'Z���n
HV��1��J�)LdX��II#\r�[�{G7u�*��m��Z�#�L�)b]ڼN��H��"�9q��E�w,�wc���ŽlceaO-��-�Ж�P*���+�#U�nîy��
U�z�U�vS^U`�S��.�kiE*CS6�mVI���.ì:j����0��^i:Z�ovjZ$ʂ�ئ�"@qڒ\��cY�&F\������r�*�¢��z�d�r2]����l����5�7Xֵ%U{�m[u�j�u2�+Cp�^�F�Y˙6�%���ކ����8�q� 9��%���-�V
���.ؔ�q\��l)D�t.��j�C@�M���ܕz�(� �'e%
�4-�]����0B��v�A.mm�,[��ui	&��g��#�guSl�ܫta��I$�^��j���фL�$v���n^�Z)�v7j1�/Hh�����=j[�ޅu�v^�V�[]K������p�Y��x��f8B�W�*<,r���VT������X��T�x�HH�{S ��&OD��Y��Pذ�*�0�:n�ջ��@��Y�eз�Z��)cl$/Vc��s4�0�T40��gf�`��]fG[����DY0D4=	V��f��iH���$�f%� ��R�
r�,a0,/4QyY�&	�7}Oy��˳���+1gCy)��	�d��ec�/v-��5, �����z~׸.� �{��ʣ�-d?��#:3r�e��K�j1)��[�U%)ͨ���z�h-�w�m�fF����A0Œ������(@�d�"�(,��#lZl�5�i��i��Jm�3�J��m�S0�5��Y�eѡL�3`��U=)z*b۽0��KәW�*f݌�v�׀��ج�6!��AfI�V�uB�;:������(�(f+�kwD&�zI-��e��ֲ%wG3rޠ۵���Rm�2`Xs�L�boVe����1L�ȯ~�Pʫ	J�CV��������,��e�T�R�9�2�2=��(���8��r�Ԋ�m�����b]�S�:��fֲ/UXJ�c�Z�]�ޘ(��nH�������#WL��+:;b��p��j�D��ɑ��G-V���J��Ա$U�h��5!5X�$�Hٽٲ�^b9x��a��K
B�ՕO��6�`��3����b�jR�ӮVe`(�^9�*�$��Z��;��x�4�N����/m��XՖ6���G��&�2-;e5���3p�ܬ�sT�2��JYx�vne��z~�Z.o�Ƽ:u0�5XN�yLj�4k�i^ؗ�EEM�؏˙��u=��y6i��`����wGZ�ɤ��ÚԂ�2R�	bAq�'O˶Y�]�u�yئ3e���*f�W�=��)���l��qE���DKf�TҊrz���bV�%Ƀ�i�U=強R��\��[��Gʢ�N+�����A�U\/yD�McY�̪�,t���7R�0r$ӵV����Ѫ���r��ܵ�k"�y��q�[Ƀ֟+�m,M#I*�}J5�X7j%M>J�iD�ĺ����+�Ҿ;D�x�3Kd�$�oV'�k7QWf��z�Y�E�G4�-���c9���W�`�MDR�\�4�V
�D��������Q-��Ę,��K8Vy�F�K�P�G���Uj�@M-k1_+��X�+H�qF�J���O-�"Ի�r�cN�5�*O�vvp�d	�c=���I)�m-����w3zoN�8�K�q(�:��P�'�[�Ie��а���6	H�V�"	K^oG���ʥ�8�-k�4�Ԉ�ԥ����h��j�:J�X�LiDR�PȤ�,J�%)m*i����ZQu"�s\���V�Ցv�����Nk^��f�H��=�Y�q��q=�a&��.��![���T�涖4��z���^:���\�*i!��ܕ��A�iP;��e҈�$M.����S%-44��!��<�eYVE��y�l�,��l���MN�;#Ň�Fov�S����D��"�1ϻ8
��S�O�oܙo�6��={��,]v)��o%i�չ*�`B��āz�6�;�<hd`��k��5��T�V.h�`���1R�JR���̛<��kM{T򕬴���G��8�V��6����7�����Y,����R6��4�8��Z�Zp�o���J'M�ɽ7gx�S0��m�7�4��nGn适<F�P<�%I�Ėgg8�x���(�O�v�&3vN�E�h�)�tG�J4Ҧ�NҤ�IjX�zo$U�;e�Ŭ��Y$��I�eD�ZQ6�L�=eY�Q!�Q$�;f�wZ�:U�QL�6M���*����-�%��9b�-����n�ӘL+B�6q�H�!�)fq�Nc=-�.�l�$7C	(�)�4�V
�����=/Y�pa��q�0�꨸h��	�&�5�rX�jJ�9��3������(*}���c����b)SV�F�4:�r��ޱ�}���{������=?������
&��?L	�����=�-wP�H��WC3nt̻7���o���(*ٛԺ�jU��/��F����ZNN*�$�t��ΝK�N|�ə�n��V����<9�{Vk4��p�Y1ʍe[�2��j閻�����Vz�@�ل��@��N�qU���6��H.����TY��O��B�LmY���a�;]ͺ��Е��M���Eʲrڴ�^�陆#t���i_!¦]3�J�p�+���9t�K�4h�V���b�S�+^�B�yD��)���|�6�%�v�Yހ��G�VD���ݜqӴ몸Gè�4a�yr��Ǡ���l�f�c7�޻��+<&)u�緰�[ɍV��孷ҭ1v�8�ʙ���
٧9�w��9��S��'~�J��7�e[�=�(����o9��}#U��Z�̹�
��`���{����A]��O�Wm�rk�<�ܪ�6o)@<l�;�ZnID�+D�Ly�K�w�aV��ov��3kl�Ok7u13u�03P�T�&��0:x5�ǌu�"�n�lfu�T��r�brp�U�aN�k���
C�L�7�X����gc7a��l�S��^�&���-m��
[.�P�Ps	��d��î뻓d:��or�{��B�]L�,����w�r�̱�X�MႪSʷ� �	f����Zp���a��<Ii$�r4�P�ٌ)6�%o[5���ܭ����ROu�8��xK�2d!��]�����Xa��H�y�G����S�A�UA�s]�H0����ْ�u�%���g uR���l@�gH�t�u�jC�dz���n�n+[0��y�`��텩3[�����ݥ%�z�;��t��S@�=:�K����U��}�����k	���CN�D�	ʹ"$���sOICך[�xu�4�_`�l3��#�X�eM,��H�d������<n1�]!�����6�ƆP�.�t�����ªu�����a���5�j�!ъÖ��p_C{W��X�9[k.�_jh1`\�JҮ�*��%�Ӎܼ�%j�8V���4d��x:�-���;n�,�i�������x�5n^��:�k޻�y+���k���WK3v��:J$c�K��_"�n��s��sg#iZ5��t8�v;v�e�a���>�p�&,ɛ�AG���xD�j5c��J	CΎ��S�ڌSbfg��"���`��n���A�w��z���5#���7Ve��)�5YMӡx��2R�p崤���Qn��KA����YNJ��);W����!�9�\J]��ĳx)���=��-�����Y��'�گ�M:��Yf^o�z�5Z�)�sݦ�a�j���ޕ��[H�E��9Y��aP�$�%P����|���.|�,p�&Z��X�j��d���90.�H���q�#6.�����ޓ�Lu�gu]�\��wtINQ��n�ǽ9?OS'r�m��U�|Y��X��^��i�|3z�)j���ˠp��,f�Ř�^5øɩ8���dɴ�����졑IX^���h��^� ��t��$��j�1+������{L��,�<Wr�cr�b;bv!�u��C���j����Fo�v$���оy7+�֊P��$�P�s��h��qu���b�t��  ���e�ي��Ci�k���:�ԏp��v�`�\nw^��6�viw�S�n�<�-ecz��d�]U�/�&o\Jol������	u3�l�ޜم+�32��K���]�u^��Q��u֎Du��r�g!���A�o+
+<��I���r%����"�l}4���e�u����zOpoƶ�m�}ںk㗴�_W�|(N���{:żAǈ�� �Y�.#�<�:��c���tÑ���R�Dm�,j�޵�|�ʌm��c��4c�����n���]�@[����/�����0�^lES����L�����&���B�kniR�2� q�mdj��]裆:�4N�r��k��]5ӷä�K�a�����}�n���3���mJ�M��$�B���le�*��n��ŏA��-e5�T�����Tz-�+�t�e�Թ��J�K�J�H�;ҙ[+����0����h���Fd/cpvv-��z�Xj�x��^�s�v�媝�e�X��ǻ�*u�j���On��8@�X���n�V�L֍��v���+�ND��;&~Z|E(E84n�&���)2�H�-+�6n儫�iKQD�&�;zA�;f���]r���{��Ĉ�D���مoy���oTo {�YmN�ī�q�G^5�Wa��D�k1��fo^Z�xC�;����H��p�q�2���={�1n�3��`<���S�D��%�MNr7s��C�]F�[�I�5=�>������,UU�W��^�WO6 e��vK�웑�!u��۬��fEܺ�]d�M�.�
�������]��K�&f��8�mgI���.*��im�k��k)�68m6�x{�G��뙴��E�<f��f;�����+s���Y�+���M5�8�ι��㪈BV��L�}�܈j�t^8����8�E�Ύ�O����9+�(�t-��3!&J��^a.�X{�\�/�iɂ��[��/�*��ĭ����;%����1������/j �<kta��k&�9���	���a�6�Q��IV�[��yc��y.�z��j�X�\�u+��xQ�O���SZ7�������l�w�q��R9�i��87��y9�,ݱ�B�bΎ���D��O77Uݺ�P^��Ǹăo��9V���D���y��� �W�9rɡk��9H�c!��rx��ٱ��pN�]ڻ��ӫYѢ�j���a��W7��J�Vs��jR7�I8Qz�s5og4I��7��	U�M0�}u+k�U�I�G2]\ɵ̆�"��\cz7yW<�6#����Ҷ�7��f�}�!2��v��ӻ�bER:m�S�D�ܰ%���6{,51e*�.���P|���Kװc裧��X����na�WW5��*�;F�P-k�h�*�j�Z<eޖ+��:%O�m�n�o
*e�k*nѷX�i��A�Ⱦ��s��ˑ5���mm��^��|bK��㳛A��P��1��X�f�XΠ�����p��j5��M�b	ٻZ�ھ)j�X���S6�F�_����.[ �gU�ҸJ�0fm�G�67��"E��G8NY�}yCl�p[˗�<s�< y�T���O{z���5�cj��-
���2l�;M#�=�x�����ݞ<-��Lv���Q��X��!ۦ�s�Ne���ם��`˥x�$�J�gX��wm�9RQ��j�V76�Ә��s/�T����]��(5N}���o��tJ]�th��V�]�1�\b���FXYV�ي3ӓ�K�UI����##duT�e�����"`c�/��c������ʽ�YE�o*G�$��f5����mWz]�v�^Cs\�x�4áp[�'<.����mM�&����.���OJE�I��aER���{����n�N��K}8��p>�qs%�ru��T��b
��yt���0��-E�oGJ7���;=٫+X���.#z�P1�9Vm<����Y��Vʼ���ʆ$;�r,���0�.�m��C�Z�Ltq��E[��.���U��C�d����A]i%S�4�m��;�ӱ��t�p7��GcE�X*��_γ�v����n-=���=ttV�C���h7K	��A4�q�Ӈpo�㒧L˰�r�i�Ne�#�se�N�p�F��,�(��u�8�l��0�F�:�U#��%fΙ��5gh3q�կa���D;鮷�3��mB�#j�2!��3a��4}��V�:�)m���4��f&=�I���Ygk�Y�3|񧒦f��k����wc0��̑�N�Z�[s���;�I�5�ñZBt�v�^ٵE�-��tx'��C�k�I�v��ռ�COʃ���#*�&�I:�xH�;ܕdA��5�;fYM����q��Y��s��4����k�rcN-��7k��k�޼@��pQZ�0��Ʊ=��Ҥ]38lY)m�\,6�X�(�:��`���PF���on�e�`���&���M�ox��y�-���᪲0v0%���zQ����<,)ʬև�X;y������=ь��kn@�F��}U���|�:�U9E}�g�
��Y�x��{�bOSvy���bTs��^�L��`��:��7m0;w��t|/�d2�+qu��fPIgi�իZ3��b�E{�K��=��N�G��k(]{��X:ο���/�^�Pqe+F4W]b:f�pU\����!��fe�*�h[%��n̾�2����ܖ�����pT�3�U��\���P�2��C�0�����:)u+��a�����0}�fSïn��|Fu=�4�|�ͼ*�Tշ�S�G�so/l�=ů],qaF=ĸѻ��w]f�R����%G.c��j�F�EpृX]�-g�sq���U����D�f�{{�RK(J���u��ǯU�����bCE]��+�ܠ]@��#N:�>J�m�Y���e�������T����$.=Q^�B���$u:h\M��v��a�|tX<��W�,��]���H��w�b�����]��U.���^�>��ڈ�2]*��G�:�Շu�@����/l�٦��]9ۓ9�wT�2��Ca��N=�[����ly$���Gk�e�F���ӰG[7#.�3:K[�# �,|P5��z�������$������[A�(U�{UPkÔşf���q,>�CuKi��]Ӆ�n�
�Tru�����p�4�7^�ٱv����ݧ��.@^h����AI@������n��m��vK�¯
�'�^��*����������Op����K-���^`3�D������Z�\�#m�����\ǯض�w�7�:��fe���!�#�C����O	2ޥ@��z˾#2R�Wo(f>��c�]]M�/(An˽̜�L�l�hJق�I�`�4�1�W`���<�|ý8̙v�=��s�hx	wwqw��/��x���_A�%�JI/�0p�s�+:W]V`t�E�bVg@�
�=��۵7��k��!qb�Z�^=�xŎFwwD�s�儮�K[/���ê��I�;���Ű��u%N���s\I��xء�����5k9X�6	y���.q\�Q�Kv�t��gUM���_Ch*붖#|�p�,-�Q�y\�vQ�]�Q3&�Nӏ
a�f�L�%��,����̙���5��c�Xĕ�m3J���cj.M�\v6sopUs��~�p�|B���,ǋ-�c6���Y}�QJ��o}��	r�̗��5�jtz$fIZ]�i<��^�A_fӮ��{��j��Z�Ѩo��#�7�Wr�߅�>��o"S7	��Kl�jyVp��7\�-��((#K����<�=�w˛��ɼ���]S-�`�������k7��U/Px(ĺ��Z�ܹH0��Im7!�T�^gN���#YW���V��\��`p�����}c?(	�4���zC��ؗԅS�%�7s�Ǳm�X�T�u�锳�h)n�%]���n;�MKޚ��m�R�Ж'ث8���S`�ݲ(��:�ݛ+��V��11�^p ��^�,Α{����ێw��X�w]f8k���F���]���ӫ]bMS#1�6�/l_�}���ݞ�&#h��JT��dwoP��V�p�V˙k�x�1_xE�7���e9��w�����/��H����I�]�mp��o����Kӭ�X.��oe�]η*���t���£�zF%*f�-���s��h�|���{�@�r���ZNs}�}����ݍ��Z��������	��8�]&l�-�xq�z��q�z��S'Fz�����+���r,��y��WC���������B���yC�)70�eVP��)p;3T\.�wUr���T�ު�v)�ȯ�}��]��
k�{����"fJ�(vnoV��SQ�kt������{��+}�NCsٺ�t���5V�I	���]�=����z����@C��wD;�jn��HTC'�w��Z�
yC��������^����5���v�CʤM̜��O�� n9�/P���K��'{h���.�)�V�wpCP� \*����59��:�xDM�d��s(^D9""{�^��u��o-O=�S*�)s�߲�	��y5WP�U5e ީJ�"��mR�B��� �#�����t�(*��Bw�ۀ����� �#����������>���}���w_�����p��D~��*���-Z	vE���6���׈�.l�[�[/���i����y*֨�έ3�l���ڎ؛.>o�VW%��B�+��XN5�E�M�_$\Q+�Z�utwq;�+O�B��ԝy�I�oq�)v�Wj̪�ݷ���Jd��IYyH�O=�y���_X��1J q�pYt�e2�)]�!��م�,ޡ��A^�٤P0��9��w.��l���U��=�Ev���wxs�1>���q�%��ꌙ��H�}+	�m��m����d�#x��g;'_-�UM���o�mH�P�-�;2����Yw�w7ʖ��]�)�7�˹5�+`��Ir���d�&�\͵�M���0��
�Y��-r�ʍ��3*��T��ս�0ԧ�l��������VRr#1����n�۠�r��e���|�ۓ$�F���t��I+�=��QQ�+\o^NEeŠ��.�X���alxtme�����z��<&�/8)˒R��I �]	�;fˠj/��(K:���(��m>�?W�G:ūI��3{1�v��T�1�̗aӠ�	pMy�L����03l�%�Nnþ(y	+�D�V���7]�S�=c�n<|z�\q�q�q�x㎜t�8��q�q�x��8�8��8�8�q��q�qǎ8�n8�8��q�q�q�8ێ8�8�\c�8��qӎ88�8�8��8�8��q�n8�M4�8�8�=q�8�8㏎8ӎ8�8��;v�ӧn8�8�=q�8�8㏎8ӎ8㎜q�v�8ێ8�<q�q�q���o�����j�}��o��ɝ�����7��b�ծ��]�;��s�heu+�����V�H\����9����z�_kI�OkXW����fY�2�y%�C4�+S��Ind�We�7���<Z-�OkL�15��r�[ts;�4�E���ˁ1E�虽҄���ѳN_zE؅c��nƖi��3Em�ΎѸ����f꜅˧Š��w�WL∗�Us՛�	u�{�C�N�)r:��s�싣�ǻN�%9�yպ�%'�C��gl� 9,��UF�"va8��#r�}����iP�ͫ�W*�#�ַ�DT�͌Ӻ\�:+�W��nWSG_C ����M
�mN�x��.���vȼ�(z�qu��#��y��������5�L�+&e�}�2�G\f������De�q�gMC�bo^\�pv3��7w��ek�X�dK���g"�[�{ҟ:�f�������j��<0N�V�������GfpI��)Y�*/%���U�ڗr���i+�^тelZk\�Lxʆ'���mK�.gfvg�&��$�t[���uu|8�W�n���h�Q�Bڭ�M�V�f�����wܘo����.��wx�̾��H{��Q����y��<��8��q�q�qǬq�q�|qƜq�qێ8�q��q�x�ノ�q�q�q�q�z�q�q�q��q�q�q�q�q�i�q�|q�m�q�88�8���q�q��q�q�q�q���8�8���8�8��nݻv��i�q�|q�8�8�=pq�q�|qƜq�qǎ8�n8�8��f��wy��2���VKǽ}�W6�͜��53��MP阶��vD�L����k׌�T���WW>��R]���&��˺���S%��7��t�� "�t!�G���M+��[S�q�C/���p6�I ��5�=��͚#ww����h�C��ʻ���=�1!\����]�v��]Wu^��JWB���Um�U2IB�KS+:�X'{`���%']u'��R���}�m=��&\�Nk�p�n��)�edkF��~�ͥU�k��4Rc�&�չEm��c�:5q�Vٔ&�o�y��Mio6n�Vz�!���7�w��թ�R��:ꍾÍ�Kz]+.���wp��u�.7���J*6�2�m�.�#��/^-t�sv�O(nn�Mӊ2�VA|ų2�����G��M�k(�铡巖��5�﷠�߅:T��G�j�B�o�g��I�yOh�V*X[��A�j�Or�V
����7����,e37	��0�1v�sG ��b�������R�+)��3R�\�rn<:Z�)s����n����Ѻ�j�z��9�`�v�vɾ��s�d=M���)��w>.�L�$���Y�a�a����/��\�puo^�
�q���V�6(g7��|z�����8�8��q�n8�q�qǮ8�8�=q�8�8��qӎ8ӎ8�8��8ێ8�<q�qƜq�v�4�8�>8�8��q�n8�8��q�q�q��i�i�q�q�qƚzۍ8�8�q�N8�:q�qێ8㎜q�v�ӧ�i�q���:q�q�n8㎜qƜq�q��q�q�pq�q�q�V�=��ܒegA۵�nZ;һ]���䬖5`u���1��m�"ӛS�G����ΗA!�M41�c����$ Q}or��t=�P�Niw$�EM�v�Vw�s�)ݽy��L�'*P�8wt9�R��z��ch_o�e 9bV�U�.�u�5�k��qS�9G�*7�k2q�)%�ū
Ub:{G'*�
�73��b�׫�^o[/�-���NԨM
��_!.}��N`�O���Z����Uݱck,�Gvte:�����ݚp�D�XgI�2"��N��yi�@H��g&N(?��UN;9��y�.ކ�D���C���`��z����fos�\�fUc��s0�k�*'F�y&t�G��"z�n�U�J�Ȳ>�J�G|�73�2ͼ�m�9��]�؍�������G5p��&��:���U�BΨ��t] ե�k�c�x�ȏ%%��u�pC�ӗ�2��-��
�RA[�̮�*�q��H�$U;�]����U�JԾ�G\���#F�-ϩ�ђ��Ml�@�*a��&�����8A.`�˪����9�w	N%�0)�ٚPccγ,z9;���6��@�ک�<�A���j�{����W-Ƀ����lv�B�s���5xw�B�m�z�Y��glK��m�=�6�w}A�@�̩Ѷy�7>�Ö�O�1d����ر���2�I5�1|�A�剬-�'�٣�����X��H�J��j���F�17*�7�_wL��P>f�� 9��Qt��E"I|ҧ�I<�!��p����e2(_H�e��gl�YON
n+�	�ܱd9�qeZ�뎎��c�"����V[iJ� �/��X酌t��ǫYư,\2,�˻%Q9�9�����}R.�U�#�����x{�ۜK�Fe�KT^�c�d���u��=����̫�fo4��R֑@��WfM���L�p1��I�Z�(t��n]�p�]��x�gfve]c�⪪�&V��rۚ�,�ޜ�L�k0+4R�T�̧����v���}b�b�FI@a��t�� ';o��8�l�3o��k��2�^���KSX.�NNΪD���h��\�Hsi���$T��V�Wi��	�.ww{2�A�6P=����k[��IUt�P��'�mI-��y�.k�SR����;p-��n� �UQ_dDV��{�r}�| Re�mnW\�[#�]f��0<(Q�4:o�v��{��| �a��7����}`BH,�D|�����u�nK{�\S̖��U���{���&E��ܙ��+�pl�|۴_S}Z�8]�&��S���9�/��!�&U���v�2�ko��&qN�ua���r��B�=?�����j�����;����rZ�*�zxM<WeQ)X{�ۆ�
��|�Hl����H��w9�|*��R��8�`oBŰ���O&1潿�d�|$Y�_<���\�s��P�Q
	�������"��,"�MM���:���^s�$6�oLT�)��)���M�g4eq��"5�3��{)^��U�-;�������]쀻Vn!����2�dc�Rͮ��b�}J��˴Y���z�GM���Y�t��'B��C�f��q�8]��CѺ`N�je��e��(�u�͙�u�xډ.��ཛ�dM1�+��O�V�`���į���:_3��uL���}T�a�}�[����ݕ�|����V"�=��:�k�"�쓵X���@ʌ���A�[:�F���|�3����e��M}�4�/HB��7KK̫iM�\�/^���]J�G��٫���Ǉ�ƅ�= �m��)��T���31��#���/�OgX�UV�W�R�N�g�ܰ��.��0|[1a�z��\�m�)e��n�s��������s�y�k�5��r�J�2j]��Uk�3p�8M��q�S�`D�V��f���@�u|����K�P;�ڬ�X���e;�F�E�����f�5	�v�yRj�H��Ӯ�Ʒ����5���|�K��2��d�Ԝ���r�U��Bʸ4��Uכ:�lV䣹�,!4TN}e�6B�}u�+�E�5�S��mX���
��n�;&rm�;��*��H�K~��1�*���'�اw���j���˯V��\���{�^����j�_G+�c76�(;g��#�����T�y��̏*���ަf��@pm-�����î*i��
���ޖfiG����\e�S�~�YJoN_�o��]�*�<�=�3:���t:�Lޛ��H���1�������tvQ�,��x&�`��DS�KV��-�X5��,sՀ�ب8�6B�o.�m���l�P�c��z�Ė�#��{՝���6d5v�u�� ��L�ںt����h�4�9tw{ܘ��3i�YdI1�� ����ڼ% �܉2h�h֎���	ё[.��c(�N$�����v<<ԛo�v��J��eD�Z弤]�y�쇄3,ரI�7��*���b�e�`��[�6Ҫ�/��1P�r�>���S�;"|��6�n�]��|z����`��S���z�Y�5)�2�]S�7�e��fҧ۾�� ���3H�Lmv�k�@�(Ǵx s5r������b����ڬP�z��w�if�h
7p�
�Xv���P�ť�Z�YBd>�nd>��N�������JUh}�Z�p�Ӻ���(�;��mI�ga�P�C�VwR�ŭ�B�������V
�<9��5;��n���0��.�cv�nޤ�^�kV��˿Z|m�3M�t�4۷��꺪���8c��m�nZ��([��f��yu�w�������-0��_�d��:pM���c ��uB0��Wb���<*#�3<���d�A��и1����s�Q��u{�uI�����Fȭ��v�b6�wgMգ��Fn���ӈ����[��z��c�0����gyd����ۄ���$Мl%譄�e^�Xo�2��(^�Õ�n����[�)�fť���O��'��fo6��FT�+(���W`ܫ��T2���vm%K���.S�OmT7֑|.��IZ��lwF��i��:�yU�EVQ�ז�����ۅ��$Y˦Zø53���E�"7���w�׊��%�����t�BM���nc16.�n�b���m�7�L�[��X{;;��VG�u�#�F����T��r��{�5�|��uA��-yoa]g�ك��}���U��nY���BԪa&3�ɋk)v�k�h��^�ُN>T�*� d�ZT$pJ� �Fp5��Ww�dp�ϰ{S�F��zèi<�D�l�u��S{�_7bCYO������j��#A��/��KwH�Y�AE��5ed��&86!�c˛z�U�uں��:�&�t��m䎂T�ʴ[g)�fͺJq�o����3�/�h���.^�9�>S�rv��贺Z�I��	 �'��T��t�:d18�l�����^�c��a7[���!;��]��:f�{{k�Ѻ����z�4�v�M�O�#���G�Z�����$�j�}}�:��m8��9��Q�m���L�)�E+�34nR�Ů�vk!<�C���F��٨���x]�Gѽ�
��\ȣ�ʡ���{���)�ԝtt;�����_g��j+�a^�� ʁV�8a�[���+_�T,ۗ���J����W��*Gi<��q�V�K��p��X;A}}��aخۆ�
ć�[��U���'[�'m����VԡF�Zr�U5���a���ʳW��Q_ �jF6Ґ�͠ޞ�՚�$̹Y�R�������4b�h�wy���.K�/7G/��gE~o���j�Uu��	S�J�-u���ג^����<OxŘ�4͙F�UO�}��H�R�z�I-@�Vʊ����S�i�y$l���Rʮ1)�6첍5K�Ȼ����X�ں��zHB�g����n�+|3	��=�UP�@�����x�ޱ����%�x&\���W_d�y�8�1�B��Ѿ��tQ�ͪ9)K�s��"�!����tM\u�:�.b9�җc4�W%�:uYQ�J~&�u*��.�.�S�b�>�,l6��N1r��L[B��u��Ё��+1�"��g6�Vр�r`����inS�8����==[�ǘ��8k��\#I<|v����#5�+P���K�n�2C�2�ޜښr"t��"�$�)>Y�y�5(M]��e�e�4���1*��Ö]��l��sl�+�J i��	J�1��=��RݬZ���χe�Y�T�뮭�]ꕫ`ʒ�`��C$F-4���h��\I�	�^��j��j_}������lӨ�ei(l�{Ѻ^jJA�z�U�e;�=͆Y�uB�#�l ��u|��++2��qX�&����}N�ڦ����Շ��^�W���=�) ����ܢ7F�]6\g���Qsi��ř4�ss�]���~��������������~����~���	�Z�RZk�#E�
�Q�dH�a��aA#m��E�6�Bbf�Q0������.q��KH�Al��`�"�F�F��4)�\�	�Gl��d��\H#a,0�m�JI���0"?�|�Pu)�IH	��E0� ��9+��E��
�b@TQ�E�
���TD��26�Jp�Q�ی0�0�S�F�$��e4!&�q����h����N3MD���iH�<\e�X�B�IIH��L�$%�P��l�c_�D2�i��%
@��b��i�Eh��2��-��k6���ެ]�ggR��l�n�r�Vڑ��Z��ō~��v�"�r=Ǚ�����_X���	?�MS��(�rowW ��S�w���Ԥ�)��V���<sy�냞V�s7�4N8:����kE��ok�fa�!J���G+Ug 仙S� �"R����7�SGxp���,;2�;ِ_f�}7h��u����3��m������Y�f^�i����6ҽI�<����S��9_3��Y�wmm��w��P��(�9�ܓ��t7Z7��>ub�<��ņ����lH/�ؾP٣��>y/;l7C��w�cW��(@�nqQt�(�U��ѹ#b�s�.�Ecgc9����/IW��}G��d|�����	W+x�:gc��'
�������V�:,����Ʀ���g���I��/9)c|3&-Ɛyvu�3g3���XNv:r�wuږ���ά��0U�1o}1Iw&�{nW^S��&�t�}d0���/�(d�ds��y<=|�w��^x��gv���%��L[�|&޶�ul��Һr�&N��VQ<�U�6kݮ�f���m%�|�Gk��r��9��mwf��g��V�K-���S��ޠ�m�f�l���6bJ"A����!��p�
Q$T��5f �BG"F B%Ơ,�ơ��� HA�R��ʍ�Ca�X��b8x�H�"#��r4�
"F�D��0��$�x�E��R�,��
)��i4yH�l�|�5����q���M������!��i��I��䈒�t��,�ȑP8�Q�h��.�""��J08�!�b �00xB���a!F5'-F(����!#(�ypl���ab,��
)��(Ȅ2DK�Tb�D�#���P5D"KnF��L��!2 ,8XL6K��E��N��ʌ �P��A�M��	1p6A\j��
*91�bH�e�a2�p���D��1�%���EJq1���Pb2$	�J!�ȊITm��g���W#4��a�[�p�Dh�a8�r$c\Q�dn4��4�7DCi)q2$4�%�Ӊ��.8Ra�b26L�H��"�0¸���)	o�F��S+[��U�c#���@��w^W��G9w$�$.�*PH>>=||v<|q�q��z�ӎ�v�۷pg(��Y ����.;��E��Gr��B��QC��Lv���o��8�8���N;i۷n�&���GT��ʼ�������£"Lq�x�8�8�^�t�m�v�rB�*D$w	"U㗵oϞ�'mY��E�GEX�wtE��aK��w���6����3K���҇�5����ɭ�Qi ���-���&�Vﯯ��eu�m���u�����[Z���N䫟���WH�E�2ȶ���d݈�w㎝�t�f�B-�B��/���ۑ ��9�]����v�b����]�s�.ںͻ"t�rm�m�:���q-��î-��^����;���wV�۷l5�M��<��՜�D����a��K!�*D�*�&���8.t���w��[��N�gNu}���~���P�wѴ���c��O����e�d�|^���iYM��ݵ�kX�K�;:���Ԑ�$u��+�/:�\�u��[�<�+4���?}��D��m�Xe0�l�I.H�j0�`�#$��!�M�

6rL0� �����o譹�ܻ�\�G|��S7N��v�<N�ۍ�O6�XY(�v:�ӭ��2�^V�um�hn�0E�b	$RI�$�(��eG$a��F2c)�a�Ih@�d��0�a&"��`��F�A��1Xn�p�T,�xbq�Q��E6�-�(�F�L"��0#�M�3����ʕ~o4�z���w��w"�tĹP�N�qh eQ��wl`e�������@b��S\��O��]1�:��7���_x��o�r�s;�b{�����v�)�:�oG��YN�f������=��x5��6	'��{-�>p���t fS��Q>���nzC��B���ܬ
��o
����P��L�����8��PX�=����UUUo�{w���1�q�/ ~��zO':�C�s��A��7�GL���7�Cǹ�xFn�W`a�c��a��W�����\NӶ�wn/���gbF���~��}�d�j0�B+�<���{n��#9�`���Q���y��{��3�$�M�t�[T��-#������3� �����]���=��o_}�ﻧ|=��@���3�.܂�{Vw��֎�3��\�������x��WW��m]NLu�o�0��]Kv	�H�q�S�m�*��`R]��8����Sߤ���,�i���:#ᦈf�\>�WՓ�u>���d�#��;����n�Ň�����X��
f��������\�s7�����Q���]u0v�v��PP;�q���qB��`���6o�Gp"��c���k=9����͛A�|@�j��7���ǰ�4=����>�s��tw� �wZ�7�ǳ{O`sZ��^		�u��'�m��3wǚɭ�"'g�=~���E>ut��MZhK�����x�zӪk{�/{�F�nz�<Z��&^�24[��c�MіC�=�Ki����9�s5�e��8��� �ꡇ���>|E��i���l�\���wi�z��HUo��[Ů(.����h����h��W�'�ݣs=�U���>��~�/��<ȅ$	0z����hۡ��+eg,����dS��[\q�2I&u��ӷndk:j�X��lU�H��.�}�[ݯ�C���$�z�A�L�wdw_jʯ{;%�:��z�M��xX.tQӯ@��Ů��Wa��d��ܚFW�E����OdL^��qKIp���Y]|�U���L{�z�5ru}��K��۱M(���VV(?��}�F���\�r�����Z}�5'�n.����{]��p������M�5������p��^�z�dy�7�=yzc�N�����=��d�ά�x;�d��pӃ�#c�����F7l�OY0N���ef�;�'ݞ��k���n�L@s��0�g��[ӻ�O����fqou��X��U~���^y��T{�t?��;�c.�L|.xzc5O�;��z�4[��/��l/eu��9�<���G���׺�u�Z�/��LKj�8��ÞwK��ݟ ����=�v����U��K���K�o�R�:�Cӄ���F@�?�T��\�y�W�mx%0��a>�}Xۊ���I�3N�GTĉ��َ-��7xc�7o�S���c[�f��?�n9�e���բ+�W,�v/������v��w}̩c(X����ם.߼��λ��Fl%��k����#�V^�>b�-C^�N���9T��˓�>��l]Ħ�\����LY�z�Y�u��p�z#�aR^��r���ӝ�VU�"���sڵ�NO����>2�m�R������X��J8��\�ɁLc1yw�s0�k*��羞s��=�������<xzT��I���Y�w��>�/�]I����{���� u�N�1�+]����wuֳ��c�Dz ��=�ٯ�<e�l�˧%�����y���H�8�s��h���{��zj~�������w|��{�=�1�.��|���'�" ��ۧ3#۟uT����b]h���r
���	ޗ�"������"
^����9m��@9�yޮ��f$�U�᥹��ޝ�	��[]y���w��~�w���nu��f�zI2^܌:k��{�w��Y l����wV�Xx;�tulmK��3ᱽ;�v��U:rs[���}o��8Al&c�m�o�,	�85��,�����o�k������
����.���h������ ��KkۻVM۬�ݤ˕ڡ��g��c��)
9���`k��t��!����=�X<�*�b�^���z���㤤��`Ţʽ��⸐�n���eBʓ�v������z��������r���飼ToZ���������Q'�%�p��X�d�e����ȀM�*�{F����,���?g�m�0@�9�=�;`���l҆˛9� �3�79�v���[;yEh��z4���b���;�|d�T+w7�����{WXs/ꕳ��+�z�S�U+��^I��}��}Y}�0��4���26|'�O����E�����w�+Вw�'���a����{�^������Ϧ�wY^]J���g�͹0xf4a:+|HއsU��h��׳�}D���ک-1��7f���s��P�$lu�P���p�l��qޣ{�f�VͰ�"����ި�$��}A	�u�Y����^�v{�zt;~����7���ڣ$4���|vN�:+e��������aj��n���ws<g�3����C���M�y�s�J���J�黖�u�W_i��J#gqu�-��Qֲ�[�T�ڭ�y{�W����bg�\1���(k���g�4�H��P�H�8�I�'K[�a���g�'3i����괮��਎vRN㱩R�e��{ebbū9���WU��3���¨xvMV��}�.\��=f�����۾'�I�}�`��@~�˶~��ںq�8�۟J���ty����Y����ސoH$�y�s�^�L�x'�Bm,~��wU�ԩ�U���z�t0��#�����>�'k�{�����K�Id[��w��{����6�!p�oC���q�jzFAd���?����m�y�����n_;�L��:�����P��:�#]q^�����ռ9xg�ܒz�d�Ci<k�*������I�Wl]�����Y$��34S��m�E��ǫ{M�(VRV˞$�H*gc����y��ؽ/=����:�Y��;�{��E��4%�mE�o��o:��ѓz����>#��5Q4!�wӜgv����O>��y�Q�Qi�re-�bxI<�w����X'|��f��txW��o��;�}D��e�/���r��y���R.��Źv��P �Z�ujgr�{kW���n��t���Վ�K�ƻф�WPmls\��ӭ��{dxd��%�U2�]+;D�/T�u\�/B��ĖK��^=��o>{��{|=�Y{5����9Ry�,�Lk+�<����qs��zW�T��_z���~���U������ƝO�5j�S��w�����fI�ͻ�u7G��� ��[��������.�cot���F��m=��IoA�}�C���^{>B�^a�$x]/]6籕fs{c�Gπ�������ݮ9c��փ�?I�y���X+)���}�nv�՜H��1���d��f�u��t��ϵ�g-�4��a��7�pg������������"4̳G#�ɃX�~�TTD����ܻ�>�@�V�@ �@Gh��*��dY����z����=�"�s;*��s�}��1g����u�r�k�����jټ�/)���N�g�=$��;few\���o/	_^�s���ț��ǯ���t�`U��3q��8s����y�ЀK�^�Q�\v_�@��{N�yFz��ק�SV��uUC>YcGI+{���h��^в�/?6�wNx���t~N��E�qŻ���\v��C����Q����wZm>�׬�~Y(<ܸg\�}�V�&�댾���|�0o���~?��V�K�w��0�Ñ^�{��@
^�/�����j$}y���u��������5@`K������'~��̏�'=�ﾠW��S+>�o����`��_0:��0^:���e��R�9OW�^�-��q�;�����9�`�w�L�&����y�eA�3ź�v�uOS��4#Y�I�&d��u���g�o�I�9�yt�X<=�q,{=�V��]Y��Ǫ�����uU�t��-����o\U��n�y'��i/��N��)����G�������t9�MxϜ�Uz2^���3{����E�����O�^��s�wQ���3 ����ֻ���Zs���{݆�{�]�c߼�]�9rz`�O�&=�#&t������p��t�t��?L������Lг�=�������7� �i�+�}|��WU���^��D��-܇eu,�¶bo�& n����Y����e,�ڻ��N������|IIH$҈%� �:��s��m�3{s�Ξ�tb�ٍ,�7L��]3\�k-!�w����ۗq�2}&e�8r��c<�ɶ�y�ѽ����NMs�N�Ƈ����Jޫ�Y1{td�&l̈���ӱ�%Γ� �x�g��k��l��KٸRgȟj��T[w���)�;��}�L���4d�n3�]�>��^���3�n�\ _�n�M�BFx��Q��u��{N���T����m�+��N1�i�=���sxz��K�>�fi�g����1���ݳ�o=gv�1Ð�����s�]fI�`]gf`�wvD���x�����0g�ځƅd�;sc����m�2x����9�`��cy��|���U��5����g��7�����;� �rl;z�_ds�8�/�ɨ�]�Gn�5F&(�?���x�# ��u���KF��M�w)>�Y��U|�6x�M���xq�p��'��.�ڗ���}[�����K�w���N2�4N�E=�0�k�ZE�h3Y�ȣ�k����T��ϼ�S^�<!�[]H%H�Yݣݭ����������tӻlq�չw��_F�1}�k�������Г�΃�G0��d�[s��]Z��;η}7ٵN�Ŵs�}���\f�+燰Wb����_�������}ʫYɹٱ�+GO)��~����a��]_�^�C��x�w�2,����/�Hw�׽`E��s��6Neh�8�8	}�vfh�V������{���d^x~C�륃��/�p�jnX����=p{vl�CL�7��2svGW�p��T7��M�bI\vFoǾ�0�͂��4�9��xo�7��{��y������,�續c���K��qaW�tu;��z��ǜ��N�g$m��4�>��߫=ڢ�Ҥn7���%���g�0��"���͑�N׸ϻ�hq{���Ͼ]�������k"{�F�E�:��r����m�<�N�܋�Fơ����+>�Z�̥�2��U��6_g�H9��Y=�Gz��VrP�,�?����!��G��V�_�{Օ^��C��?���۔� }�mW��3W�gB�2c�3�jL����~e�%�2h��������x�����z����V�	���7Ԙ�t��e�T'Ϻ*�E���x\Y*�3� �V���m�r�����qP�a��6j���N.���2��v�ռ��6�ٔ��c.{S�"�����*u���ZT�Y�*�Ӟ��H�X�^;����׊A.`�Q���e����[��n�Nu�6�V����I^2��7�fu�\�-�Uٵ\��˖�c���M$^�1��Z+�O2^�(ꘜ�y)fņ�U��^:X����A��bUA�Ռe��m��vd�$�֙���G�#����m�gG�r�H[sq"��
d6d��q�s	:�EYS�I.�I�Ww�te�"m�h�<�t��Xgh)��j�����(�f�Wt5�'
*���Ռ���Yb�X��;Aw
�r����RV�wE���S�J�$��ξ���ym��)�1n�zݮ=9�y�����V5InV�;S��g!��4H��³�m�hVN.t�Sd�q|y�\Sz��XK3��K��kb��M�'���a����ٕ�nm͜�>�RI/o���d�
��$�wt��T�n���0��F�QR�U�������<a�b��e��b#��ȟ�v0�/l�-
'�݄�S{WS�����`�f�h�Ƕ ����qZ5We�HK���-��:��]0S$��IB���Vx�Xi�|3��#��u�w�\�+hج�t��vDns������]��p"��C�X��y�w��7Z���E�h�B=�C�H�w[�9M0�VU�X}γZ�(�T�O����DfrY�:���C�cO]��Y4�2-�ǭ�6����jyqI��U/�4�V����)��^�LD7L��E��<��͘R���W�{������N���n�f�\HfdC�Xn�:w_B��C��������5i���(qz��(�����{�,ɬ�)�˸@ܛ\)J�ŉWrFG���;wGu�a9��n9΍1PW9Zֆj)5n�� �[�e�lR��PS,f����yM������7�=N+.Xǈӗ�n�r����^��H.=�#��M
wu�Kf��׋��K�1^l��ܜkWP|2��֊�1{Á�7T������0ʓ1Ĺ�62���AɆ�N��㢴�����:�"V��x{j���y�Ok#��Υ={�-��yis�����ش*�!�m���*�S�u֋�[�d�TYeE�wz�y>�s�U�f#�q]��t�ͽK�]����sw9�q7����Ze)qʮ�s8r��s�\�wU�WjAc��ԡ�x3�L�Y��#]��l��m�ܑW�iQ��a�vY%m����߾��~><|c�����z��������o;����]	'G_�vW��rI#��V�TdjQ	O�����_�����������㏯�6��{;�'�c���9/���Un�.-MW������"�"�MP�CO��z���N>�����������׏xޙIHE�F@rvtwEG���wS��"�;�����:8H".6ru�ui���H��ΐ�O�m^uyrwEG}ۮ.*������:(�ŗ�X	\wRQ��TTu{�:��*s��*/�*(��m�gsv���gEE�p_��ۮ�������;��/;�Kï�����@����(눎�p�w�	q$t�� Z$~�Y�7~�{}S�<�;��������|:j��r�g����7v��@[���<w�0�exh1�h)�����ߕ�;�ZH `��|�Cs����V��3g҉�`�=.�����p&��|��=�y��� ��s�T:d^��7��X�����͒���y���|�~O$��｝	W�>n[��&4����f���+yg�`�ZZ�?�x@{�N����
l)H��d@*q�E�&^��2��fV�<��{��y!мoN�+�b%��]���lrO;#�\}DJk��]�jkJ�縯{�s�����Ѕ��)F0����M<[�vg(ޑa��@<���b*M=d�y�!$I# IB~�;��<��c�2����q�b��Q�e��Q��}6�:W��+J�y?%�s╶�>�~�(��e0`�m���MBǐG0�s�u�H�U���`1�Gd�܋�T@��
���F�.���w�����ǂ���`g�����)?x�&-���V���s{.o/3^���(�͊�3���������Kx{m�췺��w2'�Q���)}Iw�i�������2Hɒ-��rh���� ׁJ�@�z��[x!Q�b��@�I�L��xc�9�N_�W||B)L��BƩ��޺����۾�ҵ�9n�K��8sY9�>]�%�?y^f6�q7h3��UU6󺃼�{������3sH.r@u��j,8OU��8捤��=֮c���Px�G�f�~nv軙Ի���Y���kz�����[m�����0oW�9��H{�\��_��_���1�i>���Ȝ�1��>+�a�����{�����>��4�i}�\��{:���!���'����e�B��t4.�@|f����ε<{z��pr��I�I$����௏_�������;��������/�c`�wQ��T�Z�7�&�����^��-��>��̟0Z��`!'��i�qh_��c��+�����.i��I[��k�=�7|�А����S�+us2T2Cc�_��\gtI~.�X��N.`�%�Ò�m��:��zjg(��¡��7 ��Ʒ�;-iͿ���Y�@.�;��!.�-Fcf^ ��>.Ȍ��~T>@KO�+ %t>}��`Y�-�x��]@�i�lRl�����Q4�%1jՒIy˜S:~x�񞈅��,j�Q����%��z,f�k#6y .�V#6����5����qj�"�XHֶF�c�\<Ý^��C@���B�#�,���r3���憂����H���K�p�9��Bde�N?g���)K�C�r�zە��~�/�c��}X�vG�])�5Ŏc<*��f��4Jb͎S7��{s�3<�����~���z������*h�n�oICU��B��Ϳ�Ǔ��wΉ����[C��j�ۻ��W�|����|������x׏�4Ƙҵ �$'�u��y;��9ʛ���7�����k�ݭ�(�/8r�ñ1��a�to�ժo���V�4�89�8��,����>ا�~���4u�t�^l� �D�V�
�
U���d8��yS�r�w��W7s��m (�V�/����񁌙K�bMz1��ݝ;�Re�� ����5Ԫ@��F��@{�N+�-͡Ac�D�t��s�2>�����������G��|@��%g��9%��5N�QL��n���+y�mx�ָ��y�%�э!�&A��%�v��Y�,*|�%�Sr�u���v�<���=��l�yj9r��PcK�CxHO���@}|���CM'ha��p�+�����9����Q]p�R��l����I�E�ΎeE]�$�֟sӸ1�|��Tk��˳(� !��`���*���>�㋷�x��p,����s�x�E��1h82��=��s�OX^ �ܮ<́:k�"�\��`ZF�T:��Z�\E�,f,˔X�X���3�r %ݙ�[+��M�!�_�p�0X��Wm����d���@��%�q����.����bkKΔ<3_���nǠ�zAp��qL��ѯ.����Ҟ�_���h��U��&��^I�{򣀱�Az�VV{Զ�]>L�uϰ+1�h�{��pݑ
cv�w�E//[�y�\v)�:�����΀ٮne�b̸!+��9�ۛ�;_�lV�H��N���8euj�X��ce�9j���;�������?�>5��H��!$��# ��;�MƳ�^Y�}��#�|991�6�z`ϰ0,�Q3�ΰJ���O!�����t{$z�7��kwG�s>W�P�՘���㖔nG�7��dM�j鋇�yb��O�s��v���S�j#��x�9N��q��<�|�=�!�<E̎l��$��=f�0u2񯵯Z��j�Q��qxϪ*_�)�4@�����o�H�90�dody�y	Mv;��V�
N<�p�skpS��xi6_���1KR�Q���e�������#��4��kO��h[͑z��GNX�-(xlע��])��X����b6w��Y^R��Y�y{�k�G�r�
K���Q)�cy�o�����2<��d���Y�QL���V�Xz�����
�|��#��t�ѯw���zu8��PkG�)��N�����H��ɽ�oLy��r����,�d�wR�GL���4@>�,j`&S�m�,��f�
Oa����-8֔+���)�)���U�6�CmCl��>���ξ������xQZ�n<�մ��Uz#X7�+N�2�[�j�X�C��nu�Z�q"�|�p�?'꛶+ۃT�6��-�a���>ɳ'�2EYz<�3�A���|���Uϔ�/�l��k�s^y>+�U��Oi�jv1+�T�:��Z}���@g��s9�Tf��y����>�c@F��Y ��Е�Y)L��y��+��j��qmSU����|3O��8A�-i��$��2{�5y��J��#h%�Y;n�j2�S�xυ�_i��z�VŰ��စ�`.f����Rd'-J��җ[��|��2��i^�G�Lc�S�ǡ� �h=���V�S4yi%L������J`�`�]�1^����k�Wae�s��^��Q �Z�=�\��,c���X��`����@��T�����'��Ɣ�ݱ����M�vg�\!Sz�Cc.�}�V��CNl�8���X�R��t�}_m�g����k��߸�P�.}p���M|}���<����]�Q�9����O��y�W]�a���Q���ZO�5o�v=�3y���1/�pЊŇ������3�\|)H
,w��;!�C���^���l�]�KN�x�:�F�n[��`g��ey�V�X_�ȋ�L����ng�w�B��=�^�G�nkxvx�
��  ɖ<&��HΑ��.�I��� /��,8E���P��Q�x�N��f��+��ό��!��@gD�/a#+��bQ�
O��Ă�'��i}��G��J���յ;�_�hS�d��@�ۢ�j�$�jEն�}Ƿ���3Na�5���25�l���,�Ycq3�d��6�m��u����5tД�C�\�j81�^N#y�u�/j�Ƙھ�3��;�U���^�&�畫�^Ϫ� �ƘЭ@��ҥ@i�4)QF@F@T$�a�{Q�j�K�se�ߦ ���e��d�����	H�T�������0�z�I&w.;�u��������yy�i���A��b�r	q$��N��h�%\�ȷ��=���}��X����p*ϒd��k"����	�B.�vx&��	��R�f�AzO���R�1i�b7��2�R&�u/x��s@}���W4���!�.���mz%��;�������և톱�� ��h�� ED�_������ԃ���{��Bcxl�u�>�MƄτ뮲Q�h�Bʗ�_�h�B;I��ғ�Y����j���USᕱn�1�1��Co<�Q�����֤�3s�t���r��Q���0j��@}��>E��M�9����z�z��.��\��k�̶�R��g��i���|�.���03nq��O����h�M�%��m�һe��1s����[�� ��x��"e1a�E�|��
ߣ��&��Y�}���q�bӶŹ���TL�\�S���/��qpz�;�|v_�͜&>2�-�D�N��z`-9���u�!�Gj��n(w �.X�ݚ2�-pv(�-�8�n_L�u��:�Ӻ�L�p�&�C]䬓M���I�>���.�wp"8���VQ����4'���iYݪe��.��ٝr�Yf,�X�iW)n�0s�&��:��]�v��ު��o�B,i�*1�4�D��P<������#ie����M���T77k2b-*�x�t���'yeN9/;����D���N�"����z�|U�]JF	N�Q��̓�f��@�|�ߕox�	�0M��ϠS��d�}��%��4ѻ\�Pa\���֕�)���)�9���A�#>y�Ξ}�N�lǅXt�D55�ܡ�[�_[�p�5��
2<�sma0׮A~`o�͚��z1��@��*��f�i�']<����|���y/��v�H��� �1g����t�Վk�&ѡJ��g�W��˿�g9��������5����;��{kg�������0�Ϳ�
t|����L/f"u��#^	B���V�V.��9+�x^��=ߥ���m
�Ξ1�O�y����� ��2��ݙ�d�/3��{yeM!C�^y�c˚�b�,{�Jj ��ȻU����5K������s�c�O�vU��֫���Ex}�*�OeE0���4��W�+��Q �$@�,��>��N{/O-���u����`�3W\(�&��<���tPb�L4������W�#_�9��Q��
�fe���mi�Dn熂��;>>�..�%Qo
gO2�
�XIp-��pN�V��S�{޻M-�Z����Lu��%�ǻ��g*�؈�-�˻Yf]���T>������dz݈��t^�ۧ��#F�]3ڮc��bN��ҨZ�{��3\q�X�As�Jo�����kr�q�%ؙ���h����\�@=U^�UW��>�D�1�J��M1�E*((��[U�E/�����"�'�3��069����E� R����ǥs�eA/maTs�XO-+N9Ȭ޵�T̅��Ͼ#9A��0xk�]�4O�r��-;�W�[�׻�f�1;2��jW$+ܢ��ʇ;I���,������t�0?���Z�����	��幷nd�Oj�+�Q���	��}0����xD�;P�/��������О����٪F��%�%�--e+��3"���#K�F<i�=0���N�S�vO�D0����k��&�YW�����_�F�OR��m~��G��k�P܄ȟ\�8�=^k|�-��j��m��<gdJ��GB�Xfk���ZP���ϐWnjd �1w�Ag9`����B�� ��k��N�GZ�g��|����m�0����}\�tS�b��珌�U�5W=8��%1��o	L�d&ZӕdEKk�l����x	�K�OnW��|��p!���m  cS�`.b2��4z�ɱ��l�����nVK�������M��\II`��^q���j׶t�On�$?��d_ �1����,�S���"/D��ǻd�������α��v[��=�n	��;���ڻ�ţghI�^�9ci��UDyQAq�l ���9��=|����/c��2j�����/���5���ʴ���H"*�;���Vv-N����E>�cEDYd�)�4�1�4%E�TB@Ey��F�)�������O�Dkx���)�TS*)�d�_8����'�5��S�k��ܮ��YL��I^�K(}o3.��.��酎U(��� S*z�P A� 0�#ϰƙk�|��<�Ջw����x�� �����ǂm��e&�0��g��q�N2V=�Fn���NAY$���>����	e��((9�!x�r��~^�#�s�k���m������F�R����Us�Khy��7��i��+{K;D�DP����kg>T�:�|����<���-��� C+;\�o���V��|�<|K�Z��=���'��+]��y���5�� 8�s���h�h�5�+���`�[�|��/(46��Ŷ��}:x�~�M .P�TW L��1�P��/����Mj�j�V�i�������lp��D�^�u`�8�@�,e��n7Pp���臨�S	R'�'�Vp�G����p���9.$*�y���|�����;*���}��qh}�@e琟E��"�)C�]��G"�N�v� q�U�S�� ?���k��Uj������ί��,%�A��"�1���3%����lp��mzh^-&p���#�:�<�{�x�g:�*Р�w﯋p�ˉn���l���qg;�{V!X
�3������[�C��
�]�ʭ�ܠ��
���(;��*�NwY�\�9�Ἤ��oy�Ӧ4"��ЁQQ#CH*-��ܼ��ϙ��+ʡ�V�U@KL��
�� 3Y��B�:�r`z}&(K�@ҍxg3nv7'�O�b6^��W��w��)��T���=���W:��Ns� �����a{���^vGņS��W=�lzKsx�
�8��Ik�d�5�)�������oV�^�n���B
Dȱ�����.:)M�����cxU:S쐢=�6?q�މc�a# S+�
����ό��o��V�)f��$'AV��9^߽�7I��ЯG�1]�+q�7��ݓ�Iؼ7�r	H�I)MM�GG��$-�ה�9^`Ty_/ ]���tH��/��	�t����=-�Y�I����/�E-��}mA�V�D���z�K����^ލǧ����y��>|3��`�A�-���	��e.��xJ�-�W/8L��3���x����WϚh�7X[��Α9ఱ�`���TL��rk �����馺(��3o�/�J�b.�O�n�Y��� ]6Q���ڮ�n-z�؋<��6'��B��'����6��0%�B��VwIN+�:y=Z��@T��n��ƽ&B,�
�+��+_*��~�Rm,U	��[��'F[:�oz��9}�(�*�;����a��܄]��u.����ۺw�9,*�K'$Sy��h-����,7���e\W@F��C�DT.��b�&��9˳i�u�]I�_�s�=�Q� ����zu��]�����,�x�Rx���mt8��m��l��T�{y~'����O��a]�o�hpJ����Ӡ�n.6�%[��.Wi�;0�I�*/��=e�R	���\8�ͧ���˷o��,&��|d��Tv������RدٝZ�;�Ir�\L���B��4*66%�]�aOnȧ��wE�L�X���̐�8i����Һl�`�ʂ��W[ݵ']��z��ю�k��'V��?��f��k����S�ϪAPҺp���B]��̾͞zhj�/�:��ק;m��{7/J뗹V�fո�9�[�=��i�v.�R�����䝽W9�`4��w8��p��i5���0��t�b�(k����Z%X����@6�n��5軬��ܵ
3$����IӗA[�A�C��pqS�M�7��,�}B�&%E�
��	dF
e��Z������v���B3ê!���M�b���3�\�p��GU��\�<�&�%�^�u�����N�z�n�|��v�`���A3WtV鵂r�q�� 2܋q;���ŗ��4Y�l�X\�dR����x��̎���JY��x����y<�r��Gj=���T�"��L��]}1t������L�JJ�)];j���}pw>_���Rpj9r����kk��f�������b�[�W�;��|:�7fJ��A�Ǽo� ��<�vO�?�ٌ'���O�
�����n���H\/PrQ�+�峐I��l9p�a�\v�]��a��	Wڡ�ݖ��[�*P�c�Ρs83WZ�O�� ݑ���o�|��w���]L�6���앚ݣi_`�&Ę:	Y��a��Y�w�����X^�����G��u�5�6���e�ej���.��={c wz)ԛSh���<͗M[ɧڤY��'�n]�q�#�x\����]^J���-�gz���6ˉ�V+YS3a������̳����E�uKHT)��1K�{�
SBM޹�G�0v�m���%ݨ���ܚ.mǸ*��*IqhV<�V̧
�/���X�4-N�:�輽�W���%f�I+��-F!�̙s`��QRs��LU��˰E��5��/vK�ҥh�x�Vjn�c��ˏTg3nЮ������͖���>6T�4&V�%�J�Ř{��v*[�� 'Dy��λ�}:�iM�N��b���X�m*��b}�J��A�Y��Etn�����w���O�i��o-U�[u�#�WGp���w��3z���EGW�o���%Dqq��Y!q{Z��/�S:P'��	<x�Ǐ�Z}q�����z�����ǎ�����d�A��?��w�]������,��;EHH��^<}|||zӎ8�>��׮�_^<x�֠H��P�ԒF�t��+ltqq9pH����T$YB�}}}}v��델�8��=t�������@T�[Q�O�jt_��we�p�a���^��s�Q�w~�^K��=gO�s����m��qٽ��b���>K�դ~�c����@/�_־_ky��׻�ZRY�����;�2����rA@�'�Ҿ{^G9rq�9�jp,�:C�S�+��}_������;ฎ�{^D6����\q�g�_}j�<�vͺ.8��?{^V�Y��ډ��]���kl��QC
L���&]H�L�<�QmJH��Ta2�I�h*H��"��s�tQ���i,�ٺn,=�su�Y�t:���I�;�z`�Nbq%8m��-`��Z��G�mgow����H��h�j@�,%�:h�4L(�
q�6���0� bE�BʳPU(
I�Ij@�r2�	�E#��FfJH�%T���`�
�n�IA�l�! �	�H���G88o��P)��������a��Չ����z�ٶ��۬�YӜ�]i*�(����Փ!���A^ ?�H�ا�x���}Bz|��9������9�`0ǣ)�[b�ӧ{�ܵۉ��;�{��s0d��v�sy�:d�?z�S�U0��f3{ғ���i�,N�+�9��[�+O�):���׀&���2c��\D���o�Zx�,��k~�^����;&��-�q='-F�3��J���̴��W>�N���A��oH8��ߑ��؍�	���!��
�<�n��N�/�/����#)sص�ˤ0|��ߕ�@?��}1 ��!<ղ/u���ƼN2�lFR�U��M��� ���k�b�%pC/$d5�S&�0���Ķ�}>� �~��6��+�/ks���ݯX(�jām��S]�^���>�z$�?���c�H���:E&i��QYYUM�4R���|��A����:��T��i�c�41��rƗH���\���kN��L��Y|�Z{/�ۮ��32�˯������])�=#�_����R�:"�6 ��	���"S��Ҹ���u�Al"��x	� �����#���F�[A�Ӎ����c��BN:�Ale��	��|}�?�v�}��{z�te��˛����=�i�-���h2��j�\���M������m�k��b����dY෸JЌQӕ�t^��
��/L[��"8$��;����oog3�A���A��GE�h��!� +���Ux�z���(�M !M
 TdA �D[ў^�>���3z�np���~�=N����|��v�xa#2y�����m��00��ˍ^�B��v�vu��E����#\Ky1��s�����X������x�Gz�A�$ްZ1З�H�"v�eC;\Qw�p��r�b��0���������?F]��F/���y��& s&�j�}J�z�<�OJ��,��Uj�XO��k-ۤ�aZֵ��e�E�A�t��9�����1���8+h���5��?����f��9�;&{��NsX���V�U��Vk�5���>f�1遅�@"O��O�ߖ�bˑ�3���nS�2�U����ᏂmC�Vǁi�3�ٶP��'�0�"�3�[�;1N��6a����T��G��-=X»�S�w`��t<O��?�cA}ǖ�u��f�sk7^����O�LTk ����{��ι� ���>�vg1:L�u�s��힩�R��`�3^�~B>�|��Z�V����L�܄ҍ��"���>��po�=1�u�{�l�,��٪ۋo9��� X���8C�Z�̗0�[��´o�-�����l���0<�~�{{z��w��-J0�H4�Ăo������Q�oQ/*[����36q�I�8"��2�c8[�h�43�T�9��-�<�u\�y��3�$�}
��҂T�44
� AI!���>{��"r]/�yB���>`^�pGw(���PQ}�爳Y�ɠ���7g�P~�]5�ڻs���:�� �魮c��!f������A�H	P������Z�[�L[J��gns�iG��bbc�:5]�(���q�(��űok�:{��Ce�|���]=�q�6yk ��5�\�L�	�EW�ߣg�T1NZ~Vi&��˴%�ϏTt���OM�؅˜[ ��]R�^��.[��K��:/��T�+ĩ7�>��w0_Xu*���sn��_K֣���/Dci~����T����ʥX�
e^[��`nY�|��iͅ��be�3���N5�ƫR6x{���'��FN�z���UvR���1��8ŧ�',kY\�zD�`��V��g���WC�!o�7����t�L�zV����9����a�ؔ�Њ�/	]�M7`�e��%ݭ�[%�7����Ӽo{dD����`�\��Y��*�gZ*�kWAI��B�	.��t`J,���WT���l6v|5���ϛ'�)ݧgQ�y�h���<��0pV4�Oy1���)CN�]oq��cO �DU��^�9�IL� s�XqK��X�����"n��kw������}ܰ��ML=�����r�i�\�#�,�<��l�5�g:aw��Ԫ�D}~*� #CH	M"%E$Pl皞�s��h���n��B=�ѥ�x������>ʀM�;�81�Vw���^���:Uj���v:��'Z��C��͠|���=շ���9�2�7k�p::k�a��r���R�u��-�
�אt�4>k�&l���5����;pΎ.��q`$�,��k�s�e��θ�+�^���5�1�a��z@�����*�__g.�`��,35摹�Ş�q�c�Shh\��HK����)i�(;|v\����j���{�|z���]�v�������Y���ƹ�<�J	l�E�)��+�g����:��M�Vp�*�c�{��I~��Yj�(��YO�g�-ݙ;�0<��)���A���!�}�Fu�ј�-���`������w3��{ݠ�Q�ρ�d�S���#�PΉd] K(]"W�n>757z'6��Qu�6��PkOf�Y.���<k��/����)ֻLy�~�.��	e�%I��e�M�L�E�WfI�1S[�5�<ř���� h>��X)��q=ԩ'���+q�Iz�6(¡��vl����RB$-����z}7!��C��좽E�(a�����5���$��0��GZ�hX�s;%�{�қ[ܯww�IYI��'KgA���Aѷ%q���m�7�V�_.��݇�f����Ac�4����҂4�DR@���%Ww�짴?p�R	�>��Q���8�7<5ꪴ4�ֳ�T��'~��LW�1�������~|?���̗*��ڛq���2��0osq��tTYt���e��n�zi��8~ƿH�|hNG8�vZ�	�aL���*s�?��J��W�$����Kג�Os��q����=�l�!dsu �㞊~�y˳��S7�q�����t�D�q�l�s]�INtrz*��j�e{b�q�A�XB�i�mm��.��W�ޯ���T#��ڿA^��a\:�������\}��Y\�Lk��ղ�ߥ�S��=�d��t��UK���2j��<�̟(���'A~�a^���>s�Ʈ�nJ�Fu�o+ijb�b���e1��(���)z�،|}����}�Rۜ�]��%a�mY�x�,���h��D1��W1YS�\����-���0S�P�֜�6�w�@��z�n�{����|��ЊgS�Pi��H/�i����_�f|��pȵ���Glnh��t�����zdTSEtpw�Hjb�%��Ƅy�6��qL���N�۟[�~�-���vv�4Uћ]�}W�8ܽ���yw�����`��ܯ&�T����4�d�l&�q��*?/\fm�۝�|�	'�ێ��,�|Ļ����V#�����x�fC���ss�����j���r�e4O� �7�����@
hi
�����_n��yEh�>A�|��T\�6Ѫx�5��Ar/ K�9,���>1a V�7R� ����� �Ε0��g���|}㚼z|r����v��_���R�$j-Y9�S���v!O��t7�C��#8�ssi�PR���C��/���弴4:~=3��s�u}�����A�^q�2\��^u%8���7��oG�=�'HǅJ�Hg����u��׫,A��f�OW*�w~�Rbd�^n��.h�.�>��ӽ�����eS��u�y���i��֫3�aN��eJf�I/��t5�d���=5�A�6ߢa퀼Un��i�FA�����x����%6S�wc�̉��e&]�y���OiAc@.Tȃɤ�]'0S�g�U��o�>�o<�I�h����d���/%�	3~n�.*ʞ`�t�*�+��8������aU׎n�{:|������$>2�k
��c5�ڑ]]�b�7����{�wg����&m\���ڰ��/�۝j��#X!h|%s�L.�@�>�SH��݉po�a�����%Vs̺���n��<s�m6���iN����ɩ�Oʻ�Ҷ����p���Ɍ�1�P3��(Ѓ5v}��L�H����a�������y".a3Ur�؇E.�n�|��}�5���%s��O�ҋM���"TA$P$ ]o9w��d5t@f������T	��49�ǲ�|���,%ĕr��8�N�g3�L2�87pڔ��6�Ǔ&k�[�G�X7���/��t��j�B����Z戉�Zq
ڼ�t!�\���߳}N�3"��`Q�@A�#0җ�Z����N�h�K�#7�*3b�!�x�<>b�+�v��QU�4-e݁^�FnW���Ǆ�t�S��"�eF�v�ve��C!�%���a���/���sWbi�iw�z���z�k��c2�_������C�Mͩ�j]5����{�9qWm�K����xH�������a��lWT��vf�6�/h�F����A2�F�'��#J�7^�=c�O�=��`1m)Ķ�	����%읍x��/-���t�He�5�P�l�%ե^��5�*��Qְ����^���zC�fX7��1U�E�2�xB`s@��D���S(����=�e@$�0����=��x��J�gw�;����Ca7Tİ�v!��HS�_��a�W����6�vH�Z+:���A�yu}Ϳe���Sq#��/77�״���T!ZW}�b����^�c/in��R��,���k�-�,�g��H*����,�,��A��=��,9����A��#x*��Z���v�ݬ���K���.��[[���e=5u��[ݗ]'���? hiT���P=����L<��g�n�>�u�}yw�B���Am�0m�9r����4�n-?6�;��b��j��]�J��c@x��oq���d/�а�9u��Z}��ֻl�vr�Zu���U�o3QR�3jqե)�صC��8��^�|ΰ������D����]�����jz��׊�k�кv�
�>T��T�W^���EWE����`��;}"Hx/U5}4�W�kEF�]i��;6��]ʶM����`*}:�?6��H�����in�v�C��|�e�+�w��aC�:kǺ�#��@��~�wA��sJ��k���"���x�,b�i���Ч'{`_0�PR���P��|���C�S�xld�d���`�'y�z\�qhq�;$ÑC��>L�Z76n��O�T)r[t�z�W�����~Q�jz�����)�ٸ��C�����k��`�q��^������S4YT,?�:<��n�������LFk֭f�y:���%ħdt�|C�*u�j��6-=Ǟ�t�w�`qmâ�;:U
��X��e)�m�{�����{c���gS���cA��ڏB
i���3e����B�r�/�������8r�"��T��}�l6�I�绻����72����VZ)N�)a+b��[f�*up�F�~��
hh�$hh����g��{����C�(+�ˈ����,�������X�;� ΣZ�P�1�7� ��q��z�=��5Z�O^H�0�ј��O�ݚ;���QpW197�ѽ����R����-p8��'�}5>t�-�W)P�1���a��k�X���B�~z�B���R�>"\��O��Bb^�~�.�)��f�;�3��ؘ���j[z3$H"�����"["��
�|��)���4�ꂷ��뼉WZ�a�����f<��¶�>���^9쾇���ض'��f86ȸ^��d	*��!>��sZ,���\���Pe#�ix�#V�L�ȃ^��3�u6<�����9�"�f���y��e�DK���,	y71�^J;��㸀^��񡅀�V�b�<����o}��d[�G��l;_tF!�L�7{�'��OJ��j�f�;�a���uy٦�.�X���A�`~O0�З����y�כ�Yc�}Nc[�[�r����}��e.H5�A�ЁC���u�z�l���`q�Z�R~�`��ٮ����o��/�r�\疆�s�Δ�X���&/�g^�|��l��YD�ސI�^4����1��t�^�[|͟����va���Z��NAI�m�}3F��g��p#��Ę�e��j&[wV%�߲�v���K���y�_J������ ���-44�A���<�L�+���u~6Z_#�� ^���xg�̋a����c���EuG����]�:�����}>=��H�.&O`w�����iP�A��oL?��Vyz��4{��uR.� �nR�=�ew�o�2��M�4��%�آ��x7�$;d�;-������m�R��	q�sx ��^Ǫ���w�`4U�N(nG-A,^������ދd\S9x��3%�#,ZO��M����)���oL*.깶�i���/`��,��b��M�w�ō\z�\�g�k����Y�����9A@fpB�s�yV�V|`���]xǖo����d�ڵP�SC�2���#J��[
j�q�uE��F4g�!)�FC�|�T&�m�ؽoW.�lle�ոa�� fj\�F��B�Q�l�=6�{b�8ށ4�"�2N2�P��z���y�l͟�_?C;37�5��G�,����t?��˚�З��A����f@�cB+��";=�G�cRA��4�
��ژ���1L���sy�4���F��v`���3�{��+S4F=�4�>��dƜ��j�e��xKZ/*E�D!)�C(�V�>f$�z�$��vn�����X���G2�o^X�AO�9Yg��Bř)��Cě��b��y}w�v:J�:3tE��*��ZF�B������2��<[�9W׷jp�.��d��;��`��eBmӹO/��U��sT�.����c�&�����jNX�	�oA��74ଗV�w6�g$Sy������8�pi��O]��5���3����vN_M�r6������Z\ʹ�mm��EQm�x��ʥ}�a�+�7jse��H���|3_4���(��{:�m+�j��%��6��oj����ңʗ́w��\�d���������m��-ʆZ��{Q��Ͳ��YO��톱�L�q���f]moY�|ʍQ7e̓ne��+D��˫�A,����Ԫ�m�$�c1
�91�Y�3yf�&k��r�idv��K�� e*g�w�#X�ֵ�@4��\޲.UKN��)x���Ji���s��p`����X��vܧ�1�����2}u�X��/�ƣ׏3��_ ��6+�J�ݘa-^�C�k���m!�6�:(�x�e�Sh�J�Y=�E���J�V�d���j��f�ʜs��%D5q�vУY�׎e�=�s�-��Sw�jv�̗����.Q*��a�u"�q�T2�"s�S2��6;�S�����q�/5�oϡzw��LnPK��hx{�Ĩl'
֩��#)nGX�s���{ŋy׻��U��W)t5�9������k�Q/
aeߗ�;5�����]Xa��F���E
�f]�y���=�*Cj�p̡+���wW��b��TP�9-u�Q<��_!����X���	�/_.���9�����Z챬ɯ���ƥ8"�&qΡu��Yr@ee6��ȅZ�����7Et�Q�/\�mV[�l�p�=���ur��ۦ�Y�'zfe.�p��u��BNԺ'rl��;9��W<��Nɧj�m�D����R���#�mVq�k)lCv����\*�+���ê����S5��D dO���]À�\���eTGz��]�ؼ*{Q�؅W����<�D���������SĘT�ׯwq���[�n��o+���m5of�4�m,i .(������k�ox��\�L���:v+5��l�s��O2Ό�0�����o{�V,@�:�y�������C�f]oA��G��/y��#͔���y:ו��W��m��i>����;Y�t�ʰ�O�fq����܃{ym��&��|h�rn��tM���T$�)a�qM�)]�]q�}���`��*�d��K1�e��X%��YB7KP�5��nn�j�U22[n�>�x���ێ8㏮8��O��<m���n�\�Gr�<�IKڲ����+)*i��Ǐ����qǯ�8�o��<j�u��*7�G?{8�6�U��g_�"�m����㧏�8�qǯ�8�o��<l.���P�(��������m�U�Mn��ͯ{p��\��=���Խ�������w���ya_W��6��X�t����tn"�33�s+?~��m�	ag��+�D&�x
���@.A��_�y�9���ӧ�$��Z����|Uy�wyqGwMW�J"��*)DK����P��V�o�-|�Yך��������u�������4��^G^q�z݁!�r�,����8D��Rz�U��Z�{C7E����Z�f�g<���w��<���N饵�י�9?��>����)��i��F@U����{�_+�ʽ�I/Q��/���i����	������<��p��P��-��u�0�B�8[v,U��3N�p��=�0�`���|�W�
!����Y+\ZV��!i�ʚ�N^:L�^+2���X!Om��.��=���N��>^?X�g����w�e���)��c�[n��S���-#=�0֫;�B	_zc�P4O����+7Ӳi�Mп{s�ne��|��27{@�n�{��49��ϕ��	�0|�|��Dы�yiG��e��{`��	�mO7>�k�Vڴ����;z�tDל���^��eguƇ Mͥbﻴa<Cxl=Ρ�>0y{l[��u�8�|>x�2	t� ���CW����ݱ�y#���7x�9;��(�¼-�W0y��8��t>�y3-C@5K��֜�1�uE���} �K<�n������Nk|&���ܰ����\��I�I��D��q}@Jkm3���)w�6�A���zx1i��;:͜a.:kqB���,�G�B�yY����o���Sz�u����������j�޿��&x�ƀW���}n�ޔ;�B�����pϧ8�������S<T'E'�G�<�j����R*��:�Mi�;`έ`Yг��$��c:��=�{½,Z��e�*�\̲��%oU*�
��SCJA#CJ�PA;��X�/vp�j�� ����ue��w���p�
>+>!�*��������[���E�
|�U{����DIn/	�Q�(EP�ػ|׶t�*���v�B�{���zM���dbM��ᬂzN�Ƶ��Mt�)�\�tK��)�JS}����CC����ej�<Т]��1�;hn���>�/��]0�U(��x��8<�G��M��v!H\f9j�mxޚ AG��B���M���$��.'݆z]=Щu�z�U�L�����/�.�Q���Z����|�^=1�x`i��@G�a��Flhv6�u������#��H��s���e�w= 24��x܀�Ӭ:�t0eoۈ��*�_c�7]3�>٣ԋU!3>fc>*��_��^��\x@K�t6�1�O�C�D4�^�T��Lfe�n�qЇmt�̭�S*��>���>�z㾞j={B��gc�M@��=�8*���wݨ3$��=���ʹ�v׸Q�d䯗Y|�sy�0G���6��Tph�����:�?;��i��nŜp��R5c{�vg@�|���a"����Ё�G��+��A���T�=}Tl�3���ih��gIק�Aj{qM�]��,@"�qF�`�T��Ӻ*{&�s�x{�����|�e���_��hi ����x;���G
�i�6�D]P̝�޾���}�Y�_H����i��3��I���� ���`|�t�B��/��?~WAw��jF9|c�U��o��F$ǌ�!��@/����0��D��@����Ij�MI�^���O�-;��a���zu�f{u�s�Ls97�A�����NN��,��)�����?@���e:�|��{'��iu���V:���]#;!T
�`��G(=����ezl��������3��h�bm� �B2=3�lЦ��׵	��MB�JzH�0<�o��o�Yt��,�W3�r5šb%����k +|k|�⽝ K���ebQ�HGd&@��J�e����ۿ�Xa�r�V�=C��T��� ���7���2.��]_5@ĞZ��]9��8h�)��E��=�o]���o;�t�3�v����)�a=�S<Ւd;���������%הF�W�"�%\���F�������g��M��jz�Mp�k9����@�kv:c/���y��iK��=4D�-��x.��b�s�8P{i;����y�rM��ڶɖq�&:��#�=4�?h�7Æ�H����܃^��]��m�=dľ@��a�X�����C����ՎY}�z�3��
ػ�c`WF���k�+$�d'پ��2��+�҇_��Zhh�O �����iF��+{˅{ }/����9�hUvJ/5�)zJ;��|wüxc� �;7����#e%�j�:���{���^`�/"�U2']C�m���k���Յs��FGP�
xb�K�t�n������Éf���!���3���xnm�{"�ts����G����	rzj>��o��Y��Y�
WK�����Ɓ|Ё�*:h��uQ��v
�x@�2Iq�)�C�y�w����-<��4���ƹ��2�z��Fq���o���0�����Ko&{\��e�a��w8�=�+�����0�ZA�vX`��7�զ��k~�Q�2�Ҳ���dy[�f5�؝�y���3�m���@�T+6	r���i������E��_Hfi�Z��1�V]=���IF�Ɍ�b���z<�J��V�z82d�`�V��~�(��M��-{�w>�^�G�1a{R7ja�H�ʮ>Z�/�_����09�3$«�Q�s��=<��r��xu�~!t,9��9���|e�7}C�����`ȿ<�m+=��y���P��F��l'Dt�ϑ��g�(+��j�6x/q���=+=�]�F�s���-߭.�X�l'�#6��V�o��K�pb��irpX�𫛷�:���ԭ#xj��/����k�#n��[ψ��!��i��)���+g���}�OM8���ȱ�aT(ܚ;����t�C�S=� ��yg��˘I�aD	�U^��ʵ�c�{�]��}�b^�����F��
Jqw8�F�s<��5���:N&�2�kZ7���#s��iG26�n�C�Y+�):D����^u��yo
݁F�a�^��Y�/D�>L�!���H �`첌���RS��E2�H7@'��#h��<���zUVR]���ܟ}�+Pm��
��(^�<|p�-�`F��a(�/-^9r��包G�0x2��.kt�f�`���w�f�X��k�-��&S0id�Rdt�O`�E�͏����������E���k��ᚩ'���
�-!����YH��Ǩ����8��!7:.�QN'es�J	{kU���`�_�0�f?���4���t�o{c95.��0;<;�)`2�S�5��8�������Py=�8������mg�AB��'S�T\ �3���xO �w����y��;^��}�_��C=���,htg/o�p��Rj�Ǟ�&����3W\ݶ-.�|�tҽ݃�.J�GO�ĕG���q�(
)�sCHu���ӆ�9٨�d�����#�ԟh�Y��ط���,���y��?J��I�
yn`��� ��&���+�=���/{[}��5�W�=��x�׏���7�y��x
��J0inyT?�0:m6��D��Y���HWu
w�w/�C��=0�ҵ��G^�n|dk2^�T��/���;@!��}ϕ��k������.�9�nAl}R�f,֔)y{���Ӆ�!n_�{��T忩i��ڃr�����{�+�5tD�PQ�޷��%Rt���/t<�k ��PY��^��!۩K�j[�1���VQ�	��ȕ���O����T���P3䓈MW�Bg�Z X���i��{i���Ol���)�3������HT]���A�T@徣@��i���|�Z�ėIA`��*�����׶t�Ņ�Pu�h\erk�ZdQ��Ɨ��>�{j1���`BV�<S(��7D�OcTS*IRaVvؼ)e�tJ^�}�O72z�n?�jy�7�1��1�^�
��Kϳ����S��O+��sD���@���US�7#�AP;�wϞz�[!���u	��dY�&�Qq�Xc��d5c�1ss��A(��%� �L?2aK�Ć�ZD�Μ��0�(�Xт��R1��O�Y�w��Y��C6,ֆ�"����Yn�Ȗ��܁h��YX27@�XQC��~��B�D��fMr��f򸢐k[�_W\:/�r[�U��oY3�ķ�
��7��1�����r��.����Jhh�zϓ���^b_R���~]/�
�}*�z�<
�e�a���ӑ��v�]��ˬ}e<��&}<��KZzy�Hކ�>���2��f]!qtQ�zސ�wT&D����a[�W=��%�^»�uo��X��a�{��-��FY�������p�m�B��L;6[Ȭ�M���C��j}�S�ס�/���,&�F�l�,�Y9l�Ov����������D$�����̣ј.4�dߑ���g�Ko3��ֽD*z�j�xZ�0��=Mm��e�:���m�����I��B��'�.��}�$6vN0v���MBb[�E��7SΫ���,d�П�D\�Q����A�, hk�I�Kս�h��Y}m+���K�z�B=%��r��6�,�4S�^<�ň����f�F
�&j@��:�%}t�9S��)����^���~FcX�3�XJ������l�K�V>z"�C���Z���B��p�($�xQ��xlY���	P>r�)��J��D��ZK��������[������'9]<c��gc�w0���lf�ut[�c���}�(�E�#4ˆ�#5��S�,b�+Qw���&fP�s{��y�r)�kE$��޽���������
��k��=�Hx,�K jܾANyw:t,���e���g:U��!vYRE�S��Yn�I��]p�;����[:^��?������д��Q]��>|��w�3Π��c�W��:yGӐ�I�\��\\:au�4MAǟ:�ľP�W*5I���(�F).P�M�)ML�p;�.P��L;;1�mp�����.x*�bـ��gzgz{���1��L��Ab����	W0�z0�>G�6-�y�t���0u���.��[���!�ȥ����&-? �sr��6��;�?L[x4k;�݅�^> ����n4�P���\H�ϵP�����	P�;�=�W݃��W<������w}�l���RK���VQ�;|�k�T�b�A���+M�ғ�:_ܢ�,���Q��)�\5p�p��O��fɲM��[���2i�C=�XCר�f���z�DX{/�+�ųJ�u�1�X����iʚ�f:gS�^�<X�Ⱦ`l�� �����	/��>k�2|�;�_�:$�~^��Z�۝��u�5�pKlK�Z<�<o��-!!C��д���:~��^����>f�ou)B������U>jފO\a�Zx�!��t:՜����^"��َs#�ϝ�~�ެ���̼��F�V;˲�Q�.�Ez0*����d�r˸LoN�*�u�W�0�����CL?������`��B�Q�4^��ݺ�f{�|���8�x�pǛV��pu���"o�)T1�[+�4�^�(��s�qs��<�����xWXYU��[�<����&8�zkO���u�#6 E���L6���O6���'�3��,����r�~����ȹg�]�|���V��B��pbԖJ����΢Y��=��ka��2}J�P��^@ON�b̉��<�|�� ����婮�.��~�B7��ڹ�tz-`9yv�3Ҏ�s}0�6>B�Xs�#OTx���f�@Tu�����1P7Mq����V�C2����ehȕ
u�� �N7K�=��1�-�
��5����%��)�h�[ˠ�Ami�����]XHׂ�j��q�#gN�[?VΞ>������Y�g��d�۞�BC)��A��nߤ�n!�d�s���=�r�>���w�xa;[y�sR�,���̂l�u�L�mD)�8�U�6ʞO|b�o��V����A6u���׊j��=]:���s���f:wϗ�x�� �:u�\�H�"{�S	��<���)<®��j���U'��v����3v�)!Y��2�Hg��;�f�-��9�>����2�A�cQ`%U���Fp�e����7į\M��w1+�ܾ��E�h3B�Yg��i��Z:,�B�Wr��g[���w[�F����N�d����yJ���E}�ȖS��Uݍ�}�%��9��~�����
ih@��y��s�O�6V_�-�;��WZ�<_9��0i>6�`����S��l�J�P�t�QA-6c�A�zy8�8�~{*	{e.�\o\�\�gf�B��J���yIt-�]x���c��j�2�u���>�,H���z'x���Mc�y���4G��v�}�N:-���S�.�V�A�X3���vd_mٮڢމ/����q^:"X�:�����,����y	g/-	{��?���'�6ENϾ�}�C�]��̑���C9��'~�%uU�l�طG��tws��]�fu:L��J����v�`��H	=��=5{h�����O)�֋��}"]��'���f���h9B)W�E�ۖ���yזx���I�,G{2��	q�N�ڸp��c2������m]����@�2u��Ű�y�;�L�-��Lg0��)�^W>�!4�'�J�|�u	-w�BeBѡI�Wd?r�X-KTqYG^\�^;��'�l�˻E,d�Kr"!�=��'����ZRX&�EP���Nc�{�Mp��q��G&6����T;[@�2�������S"�6�#��e������E0LѸvvL��I�,$�V������k�D�.�oy�k��1m;����R\+�&�+g"D���9i��$�͕b^�W�6�M^�BnqiKݫ[yŪ��:�,��"�9����]�+�W�_��\j����}�vh�6b��I�. �t�Sa>Z�K"�[�����q��̝�^���-Bp޹��_ʃE8k��#1It��s�2�XB�no1�+m4U]����/m�'D��^ct�/������X��Ton��d46Ȅ!ՌU���s�oV����f�rC��8�.��v�F���9'GZ�n���/�
�\y7\IJU��+��p~9��P�z7=*�Q�f��,�����X�7��j-�v�1'�j��_֠�Qm��:�&²7��l���}6)v���Lʸ�l�+�����u��,z3[x���(. Fo*bR�6�l��}$�����1M�G��Fs"�����n���MFgen�bmA6�6���:n܇�����L�Y�ݍ�KnT�y��!�"՛c��xנi�%�x�t��;���]]�s�ekYZ�<��#���I��:��M��u�c�^�&�"�yF������4^���Gn�9�g#�����ya�S�)k�aH�K,�fU#�$�[��w7�"�y},J�����ٖ�,ڶ��&R�����.�;`��v^�ƛ�ж�j8#��k诜Tq/�N�%�q�7���c�T���ԑ�(�
[!f͏�	����ܧ��U��� �"=�rY��o(������t1[13򽬵���6�|�	��Sz6[j����㬅�Բ��;�n������s8��p�Wۋ��AJt���c��[����]���w��{y���Lּْg��w�)sm�+Pl��C��g@gw�4C�gV���ݝ�l��0�tk�=���v�[B�m�����N㣂�:����B���]f]Ixŉ�bc��0g����X�vp�b�,O�W��Ԅ���k����gv잽�In��s}1ٷU��Ը0b��Žo�]�0nAқ�}γS�̇���M�ս��%ܕ�����Z�c(��b-�%�w�B����V�*��id5�T��%qk�幵wYbtމݧ�q˾ւ!Mb©�u޳.7�}jV�,ϱ�|�����*�V9:�4y��\�������s�ʇ��X�9-}�V2��=��T8�����:�����tS���o$��dSiQJY붹�R��� tW	e�Su%l�2C'!'fn�
�*.�q�ArK��%�Z*��t��㎞>=q�N8�_�8�o��<h�-����/'
�+�y^V�
�uI%��}}}m��8�q���i�Ǐ6_6\�RJ�]=�W������G|�e6���"�4������q���^���O�<x��!q��Q�T��u����sk��{n��һ32�-;�b(��:�:�);��w�_>m�VYGM���^��;�;;��}��]�}_~o�w�b��;�'+˾�%m�,ü��眝�e������A�e��n�2��������<����!l���8~�o.�m�������ӓ��Z{o,��+�,��-��5��<��m�����(f*,����$KfDp8T2�p�|�D�i��*C-!+2�-�H�b�)�!�u���lm�ci,	�.0�Xpn�}���rlV�R�솱�#�r�+���8*o�w_f��riU�8i��	kLF$2��m�D�� �$d�q�Y�0[M�؈�J)�D�AdU
�	��Q��n�H(Hj#|�B��'J3 \���i����M�M� �<8��\C����}��D�y\��XY��l�[g��Z�.��NĻ���Db�I+����'�N�n�߾���P�I�����ވ�ӊV1����zO|��)�<Ϝ�
�O����V&y�,�Y
���'�q8��,1�C]![���9�	����D��	�Y�s��f�/��n[�;k~f`��;�B
=�<r�9z�����ya���Sӹ����ȸ\w}J��Q���9�9[�XC u���|�^=1�x}���R9��_^窦� ;��Jc��]"��F^���SIP�T=��4���8�|��6	����ڮ���+�b����c���;yJ��oA/t�k$J����l4*~Y�Boe^Ѻ彁����@���9�;o��8�;��C��wS�,߀|}[��Q�q{i(�$7�=Z8T�&�%	i�K��a�ax/|��=�T|k˵l>W���~�����t���J.@�k��VQ;�;�0��"��>��xM1d6�;G�8�O�:�B�������}����e�=�&�Դvo'3�;$as�&�dq�h/����0�c"Y���.9��O�����|�U���_�\��Y�a��ٕuN\e�������]c-�;=�����ypt<w���T�}�4A�����"b���\ò�Y*笧/)j�{k�w��oH�.9�yۤ���6�^;!��C�;L&򱪣:�p��ɧ���)�BQ�<��=�{�7�!>]>�]�P�ҘH�� �g����|�xi���sKb�D@�'�7��_�5���9]���[�>4vj���2*-�d�����oL���`�}ܙ�����}g�7��>�-���;��+� �׮|����`�5z�Jz�D����LrS����g-�5Ξ�E[�{�f�.�����^����hB�$����;����&�
ٹki�s�T�P����-L����y�Y"S�q��a�<8O�; x6vo_Y��7��i�P����_�o@>�rL��B7$Od\:��8�`[O�)���S �Z����|ʭ<�/r��y�������F]��X�oH�^J��5^��xض��u׭���E�N��acb���[�:{�͸��\���Pe#��9�sͶfi���С�6��ոr��JryC|h����O��-���U�\�re.�z7]��/K���T���_~o)w�L�>� ���D87�.��z/=Q�M�<ՀwJN)gO'����p�SƲ���5{m7��������/bK^�u(-oyn�������*�D�;��[R�Ék��RG�M���z��ms����s�v�:�paV��ɑ�θ�o��V
=K��+yhc��ڗ�eh�E�!Z����g~��8�yǮ�\t�mp��ˏ��:��I� ��9�9��/R��̳"���G,�����mCv�}�����b��.wh4vd0 t/O��]��5]�l���M<A��ӈB�'�c�0�qh(��-�[z�TU�?P-�W*�����w�Y�e���5�������j�����;��9��P��e�0��;�N��@��xUλ�:��-10�1M��r<�Vl��QPi�'ƥ�_Z��f���Sz�DH���;�)�nC2��d!���S�2��=J
L X�K:k�VJ�k��ً6rg��5f���&��:ŕ�U%c�U��(�Q�bo'(ֶ����>�`E͚�H�.�1�-�
��z;\<Û��P.E���a�@Ol��(�[Ud���б�/p���<3��^~�u�۰YZ2�����Ǯ.|W�9���� c�<h�o'1~f�a��\������o��Z�t� T7��y�DA`;��"S�		{9>��f7���ϧ�Yu��H��.���R���kjm��HgbAoj�ܝk+�,�9t`�j	EVM
E`�����]H��Q�0�G�I��,���]B]Xז�����t93�}Б��l�l��H�7�q�ϒ}a�6f]-q�r�n��~.!��8��$t��㹬����o���R�[�hl��7`)��@,���E'�Jٙ�,���=���iU���y{�/`/�p5�#cF(>A�A[4�gj�W�:d]ct�L\�Es�K���Wsp�vld!ɢ��ký4"� c&!���1>��5+[\B/-�]��D2���ۻ7���;@']#�.U����;�i|!x�CNj�|��|����썺�d�/3�r�q��%��ΞeVְ���f�i���(|��C�"��as�r�f�:�~���BZP�Q焜hzW<��K�)r�mF6��۹��[���xws��ZO�L��b�7>��x?[ϡٕ�&���JF�=5�Ky�^��Ksp[K�g-S���tT�\���3�Ö<A�6&����3n<���1%��c�|`fV���M�5��ڍ�|ޠ��TgO>+�P����^}?��Kح��*x��E�y_|W>�����L�o6�{L4�m�����@fp��2�Yq".z��zj-��@
���>��,GM���;����J����&��c`jGq u�3}W��]����H���y�ł��4�+n�9��܌#��b������D�#S(x{<��b��(v�_E�Ys�cPB�eD%@�e��T����������t	����z|4r	�������ݾ=1��(e�R��􊣕����Q��Mnd]"�}�3�{�ŏ�l|(g�\0[�_��mLP�a���HNzD�d�y�K����b�.�55\�I��~ax�d[^��S^� ���$�c�>���"cׇԨ��(?�I��Y��U�y��aX�����\��hd���	Mw�2+FD��+�� z3��z��Q/����JiroQ�3�l���1 �������'����XJK�!B�7:3B�?��� �K_���1(~��{��<n!����z?Z�s�	�񜻆Oi��{ĮT�%�E� ��(=��z��!H��D>�2�B�%�
ݕ���/0q�U/L;� q���AC�_�@�iQ^ ��?���1~�x�N'���Zއ�"z7!ا��Z~kJ��z9�8����Z=�:ln���v����pn�n>��'�����vyr�-�i��..�Te�,�e5�����4��3�.q��H�uyb��4� [��ʼ�yc�4����xl�1��wd���+LaP��S�
�F<4kj�)�~���$���$r-�Ԩ\�1�ѱE�1՝=S��N�R�o�}��C.��>��5�,���ev��� <*���v �&j���KQJq�{VM���"�!���:����0����Ɗ�F����6����mt�>�<�a��t�|678�a���`�C��^1�{j
�G�~�3��&x�w�^a\�	���+�b�96{y[ *�D���(��`����(��ߔ'ʩ�5`��r4h�'��',!י��K��D��}�;��sz:r�GGo�5�:FE�D�����S�s;�G�&gc/��R:%7���,���
Z�2͞���W5(�z1��,��5�_���lX)���5�;�S�z����Y�<D����o�$�_�S��E�?4����܎|��+%�й��t�qr��c��M-CT+�=$2*1����C6q<q���h�J2�rz���蚑I���� ��,�>ĩq�5����?�)��zPd�k���[Uc��˧����
~;�KX!y##���<�طf ����� y +|f�����-�8����դ�)b]�4Q��uF��W=���Sۺ�
DK�qu0�G� h'#���;V�[y�m^�O���s��1%�P%�$�5���>싇Q���3� �!�oS0K�u1ݑ=ˍL�]Gg��w]"5��:��S��_s[+p�hF��>�YG������^=��j�+pҽ�2�&\�#-vH�1�z���\]w��V��i�&ձզ�+�˷P�6ko�5xp��~.!�{�����^!��߄�a���ԩ'�b�sȤ��j-�a�C�y���]�Os:h�����G/5�-�w��A���<�[��!	�U������i�P�l�aQ>��1������'k��B
�/H|��_���g�U5_%��y\�{�����ˤ���$�r��β�@��}��H2���(�Ϻǧ^���� ��B1cɦ��=�a�g�m榽�X�R��cɚ��T����&�w§P����]�i��ǂ���*�Q�/|���ȳ"�UO��!kd?��4�w���L×�c����
�i�'����Ӵ){D4 x/ǌ������1�{8�Bm�]fSC�T˃�4vİC�@8L�h/�ZK�^���CDvS:�jq[�p�Yov��Ay�6�c2�&F�����/�f�?)ޤ|X�A
�\��+����=J:j[�+%dmz�<�S�CG��D���=5�8�˺ꦗ͒^�TQ醩���� �US6��V��|V�\u�=䐜*t�.��p��DPV�}�|�䜧E����Vu����M�3������SSQ�vD������^"�LӇ{jMV4�Y�Wa�{�@��㾢m&��H�<��z�_|�lTˍ�lS��rMѳ�������>��Jr��"{nH(1W�"8�&^�RwىKW\�fq�[���|}��<���|h���w�͝���y6Ƈ@��ZbT,|�ఽ��TE;c�Gz(>wV:0f�)���P�z�Kzm���.:k�%s��\�V��Z���j��'����I�O�,p�C�N`ל؄hR�U�(5�Ʈ��y��t��s*X��9;"�/5nQ�9<�n�TscK����tD�V�
�!IN-�-�,2-�sT;nm��Ɋ��xZ�*o$�N&3�n"��7�eRb9��@d��ڋ��W�q:r�ՑN������+�H����g;�y�Ƽ{5�>���]O6��'�0��E�a�i[��:.ې��0��9�a�!���p��=҃�h	�2�M�`Gwe&�C�j����ĵV/Y�
�+��BM�������(��.�hb!x�lx�z^K���E�����S-3b���i�ҵN'J�����T�u����������ځ���\Fz�-ε�j��Jɛ�4�T8�+��)P�.8�-~*	{k���{.a�Gu.Rd���*v;"�/�iZ�Vh4�E|m�0i��u�}ut�l,V�C�B4&�I|���yw5��C�����ԏ�����?=�ֳR�¾�|�M�`��us�V.��Ί-�T��:�;+j^���#v��P�/�;u����Q���ń�����^�5��R[?{~���vپ�B�-�>�5�{�,H���vU�ը��;���J���k����;���,'��q*��z+_8���49�c�;V�r�0G�ٓ�2��۾�x����WɝZ�?yh��!��ψ��\�0�q�5��}Wak��������s�YZ�(���0;򶧕�QQl������uf�G��Z��a�=�9��{��6��IP84�2�'[H׊xn��� c��F	<4��NѢ�Y�62$5YVxʆ8�xNq�O�܂(i��O�6ܵ��}hg���N.���j6��^�خ�Qu.!Mo�[HҤcWd�e�$秵���0"�*��z���g1���14�Zvls;	�	������^����i��P�g���+���v�	q�Vl�z�q���P�� )������=��>�zsb��gτO5oD����	�c�4��dSf�iB��0ީC=�)��z/��o��[P�E��MZ���O�L�sw&�cܓ`�m=ѦX��ymI*W�#c9�eD'�s��`\�&�6P ;W����s������������O��;�������;n�Hy
�:�V��׵��]�v�9�J8bh�v��ݷ������ua���,��a�����|Z���;xP��zb�)��|\7zW+�b���G��Eλqk,n�[֥.�ٵ�3m!P2�_]f[=p���#������]�)�3ˋ��r��M�~*�X9�W���35��r�;�/��iC�C0~���-US�ξszm	elrD��E�a�����Y%�yt�~jN%�\>��89�!�Q�8 E_R�ˎ8+��C�~�
[YB�>��OB��ÚGa�`���񈰶9�R���9�����[�0_6�c.����/�5�~#_An����� ��e���������*	{���)X�����<vVo����^jȼ@���<�~UƎ/&�V����l|�z�ymK����ʺ��|x=ؽt�v9��jD�z�f>|O�Z�?ZFb�ɓ���&�,y�����Xq�c^�̆}�r����p���9Ѹ5���Ē��f���S��m�2��S,+�������+q��������g�K���`ʏ4��\Y���=�� 	��ݱ��x�}�WV�`�X!��xi>Ȩ̟=�*�	����"���q"��8^�^q�e��N��9v�q�L���\[�Zus�y��0�B�dȨ�
��vHw n��1��Q�;��Ĳ&]�Rt�'`��1� �q.�݁��;��}xW)z�qi��yh�V��:B��ɰ]D����=�^m��Ţ`o���;b�Ů��{\kP�;�~K��A�����̧/���^�Oc�걑^nz;&L�+����N(y��c��j���R��9kk+���f����u/�ג��8>�,�Vv��T1���O�bݔ���^^!��ոanS�(=�[I��\5��I:�ِm���tdו
غ:�bn��na�R��7*�7�pg~�H�{՚+,,��R�w��;2*�95�T���ݡ�sNҝ`�RE�a�t��wh�n��&�����P8��(�nZ����L�*�[Kh^�ܻ�<k�5�^	K3y�y�5���_9�T2��-Pe��@�ޘ(I�{U,�p�Y���+�ٰ:�1�
��Ѡ�@�24��}c��ɖ�i��(�{������=���J�Kn
Ԥ���0�4�h{վ�y�4��~��%�,��w��N�U��{ڊת�}"�{J�U�eFj����L&-��F��=����=��P��T�6,B�
T�Y+��?K ��Dg7;'v��}Q��y�R\jk[tvm��gE۪�X�Z�y�F����6�Y*�ͦ��m�±3�����h�ցW��g=ʇử�9E��M<�j��%���4{%K;���6����ɠ���b��b��e��|�d E�] Fbw�.��Qto�jd`:X���v��e2�##X[���X�ch ���yݚͬ��nm�&]���<����̎u/�8p���Iu�[*�wu�޼kY�`�nY{��,U�ջ�%��#�x;gp�[�=b�7sa���:�ɬ���R���ݺ��UD۪�/Sj]����Qu�g7�2���ꥊWUݽ=n.�{���Ӥx�f<S��}T����b��ja����ps�Y����{���T�2�u��꘼��f��U6���m�}�b��ؒ��UuPָ���B�w�5IfT�kv�(f��.��Q���9��6��
�t��68�/|�ܮ�:�Sz�\�Gb�c�7o.�`�%fPtnJ�:W<��%N��79��y6a�ww0.Ξ�e�׮���.�k�Q�S۩��Q�+j��[�� �צ�M���ga#xu�w5,Զ���#*螮�̸��QZ�����t��3����8��=�j���΃������v!
`�:Jݫ�g�F��'{�D�*�z*�	�ez��ڒ�A\��q����p���W]�&�]�7�C����j-�	[a���duG��m�<.w��#"�E�*ƐÓ�N:�y��M,���*�C���G8Ӕ�[V&V8f~_#��}��I$I�2f���ѹZ��N]�g|_=��o>�z�����q�=z��>�x���	$��\�K�$a!EW�c��{vt����[�|�>������8��z���}z���c�<�G@0I ��D.ۢL!}=�i�����4��m����e�V���׭<|q�q�=z���>�x��3UEB��T�˹�k����y5��nm���2kA���m3ۏ<�������ڐ#8����7έ�d�uo��|��Rm���/9m�%�s�L��Y6����,��&�!��Ӿ���^�^�IuE��%%�	q�h#��)��;f����9����{�^���v�m$�so�3�":m5���|~>�����y�3^�¡'6������v�f���ڐr�:m��ޛ�B��!OlR��9��O�îx�XN�d9����r:��v�D��y]8L�t�(�y���H����'sʭn�[�}],W�7�y���&����rgف���Mȧ{-�^3E�2=2�a�r<�Q���6+v�E�c�-c�lfoF�K�t�����j�-���$o��\�$J!$=�d \c%c�AW�d� ���N���Fi�#"e0�K;�p�t�=�Ǥ	����L+#���-�k���_����A��R�s�ե"�RJ��]|]r	}v׵r�1fwU���5��)�2u����ڂ�5ӧ�˃�$wR�\��)sȥA*��Fl<U;��.U9�r/L�<��0C#��!	��m��H�����2/C	�NV��Ҵ����{e5ټgY��3��*o	��p��]���],/��gتk�(n*��x��\��N�S�M��\�vI=���5�����Ƕv�6�<�!�?�
&˯t�u���-e��2�>c)k��u�9�0eK =+�^�\�/�޻�fU�0�_��(x-��/�Q�l�,_Ud��qB�m��� 	Ng��hߙ>�`w�� �M3����#��
��\��t���:�}ugRyWn�J����%�2�����޲�;���q�Ʀ���-N3�<�z�-Xk�1��\;����M��Q$b_xi"Nj{�bޏ>��]V�H��6��Yn������B��D�E��Xۻ�j�$W�L�6�hw�sÇ�p���5V�,��k��}S�:�]����y�6"��)��i��q��:��r�^���xg�m}���|����iе���<B��	����bN�P�oD���Ÿ��f8"�Ν�I��VYܻ�FV�횝�$m��k��D�� υ����U����G��u�"��$�S�A�L������^T��;���Ef�i����`�Ώ��xd%nϾN��tX�?�C��9��V>��l�Y�塍���Ӟ��(����ϯ�,���N9�c��H�<�zpz�w�u[TԴ7�s5Vwb�T�-����������=X�F;\<�yθf��b$��S�R7��o4ٽ���j�+�T�Y655�����󠱠-m
W*��5�c�鋇�Ol���J%��@���X���o �Ҩdw���)�ݟ#���%:���
qZ#g+Cljk�Kh���}�2��JSz���~.��2�Q�����7aJc��<%`sȪ�5���?&��̫h�����"�T��ީH� �}(�rۮ��3��|X܏�,�|=�{�!�٣X�5+�]⊣Ls=Ma3<�N�O9��6��2D��m�/�6�]�����rnNu���҄Fq��Ej<�T�r4U��h\��9s�#�W[��v�ن����D0 ��Us3���<���:I�Ç�p��*�������i��ش(�o ��#ӳ��
���Sši�U
�X��jnS�����A�ͻd��qh��㙩��>�Z� q>"��m!?\�6�B��dO��iAK����n%�{�������]?%�o���I��	o��!�>9M��n��w��
`��Y��ָҏ�MKy���d�]������G�9ի�`Z�}�o�v��
�>2�x�|���Y֯�x�X0�3��p[��H�F'���L��<��G0���r���vN6��ݎ(���z��_"�K�#�AP�CM^��<óe� T�8,�q*~c�Z���{��=��S�9��������@���������ѡ�w�~�0�Sȷf��%���[�?!�b����_��3ȁ�xf����ŕ� �c���ݡ=�� T[#���A��X��٫]O(g^*B����3�q2�'Y\��&v��	C��$烿��v���b6�:�}��Tz%ݙ]�2O�v���-�P��\
�|��U�v�;#���ʰ��3�*]o}�"/=>�sE�j��3͚u��x���s�3��%�;�=>���>�xC�IE^��<�y�d��v�VK�%y��m��8s�,v1�*u��a����ǻ/����N�n�gU2OK�Z�m|���9n��"��z
����Zi�n����ǁ���3"33L�r�wݢ�4�L����j*�`}�t��N�]5`��5�O�~�^���_|����:i��D
e��3�~u�{dr=ý��H��8�79�A�����<O�p!|�QO-��ބ�z���fҮP޷�x`&��,h�;+�Cq�泥�9^}1_�i����5��<L�9��&��3tܷ�İ5�@Oj��#'1���>z���Hqe�{�և��������w�e	�>#�l����E�TS*�J�xP�|���'� "!0�v��yb�e]����b)	@�s����*�]s<�Y�4��s�݃;�y�SS繻����L\m�~��
����Ss�B�Ԓ�@�=�i~/I��%�yt�~j8��;`>�9�8P\��~<�`0{li�p�� <'4&9���2+ITe�dk)�$ިn����y��bo��u�0�wo%Q&�L[�6�������PgVͫ�8��+��
�^��!�GN��^&T���&�P�� �.Ek��: �^4qx��{��� �B�t}Cfslh��R!Ca��<�Lc��>�z ��-CˮAi�y�6��ȇ���.��Dޗ��V~��CD+�@�Sş]ުOr?,կP���:wyԲؑV���R"Q�^r�@��6�5�w�R��<���G�B43�T �&8h�9��]`���t˻�βJ�r�+U���#^oY�Ս����@�W�@T��������l�}��..�	j���\g�4��[����Κa�Ғ��?`���Aڻ��$ٷ|��M��Ը�A���֧�5��y^x����������C��lK>۹�*OH�<�V�W��%�@�i�=�/B^��d{.�Ef�aʠ�7��ŗ���B���D�jzw,��T�-��KX!@l{@:�Lz�=4aJ�/�<�<T�׋��K�М���7f���<�,�������6�{J1�}$1�B����|�����9p��3j�w��.||0��DO�\�׌t
^U�|��z���n��8�Ä\l}�u�L!aH��]�N�����Z�^}��q^�d�
3L�ҧť��lk_��5�܌���xx@���['�C+��/��m[��2�&%�?D�V�L� �Rkk�"@�oEê���eF͛���K9�(��័�QJe���2�Q�����F�r� CR�J��1��3`��Ue�荝�̼����G�G-Ѿ��p!<��K��o����Je#����j���_{l#��}�2�8����q��V���d��W��ʱL��''f�8ARmʺ�h�|ǀ���½۞��4�6��'
]��ȮBwo�(z�t��9K�k/��e}���g^���7�w;{�6�Ō[�{�v^�=�����w����Z1���|�3s-{z%��
��\�zB�>���=�曭!<�i�O�[y�y�<��Z������Wu������^;�	;�X�|�C��Ο�������7̭�
3��,��R��o�C��݊�"
H��y�;E�F+�6�R�fZ�eJZQ�'M����������ɟ�1���A#�=�DBΑ�5����{�n�t�E��>��^���'ɵ#$nJOn��vD�T}�ޜX�����! 6nb���Ԧ��z�A�7��kCX.)�:߬:|�WI��A5��-�r\�!�w3��&�e�Qܯ9�{ġ���d0�>x.������o��\˺ڿ4��/b�N��wi��p�Q�6�^�Q���P�-?P��A��H+���"��E�n=3Q@7"\�<�f�j�1.	~́Y*��55戺�V2�Οu��{��D%�,"�����\O�U(V f��ScWl �\�1�OV3׾{� ��G�%s��W/�Y�;�����NWfwlE!�J@�A �w7w�W�k���E����ڻ`��f�s}�g�6���NܻV~��9�v�r&���i�7�+�;4�̞��s�p�z�B�y��vtl�w)7N�S2����r�����c0p�|��^p�/��#t�̠����av�Ң�Y�a^R(�u`�f���,[/�_ƈ(�*li�����gO�S��
���_��dcoT\:����ݡy5�H��F�1��]r?j����[��z�~�`��έ#AT))����g��;����s%Q�e�[:x�V|}�/�|�<:�p��[�!�䭰�o(�sS>wu��-��bߣxz�-���8m-�E�k��ρ8�SFKQ��&���h��{���g���dS-u��i[��\Ձ q4��,���U��vڴ�\COI#"3Q�8"Ъ\k�Q�<��q˔�',H\�O�ÿ��|y���L����X+]-��՞���t�}_xI��ݓ�Œ��W��h���kO���0k��N;��Fi]���c����L�`c0%s�_���u���*�"e�9�|.o��6�zi������m�����c!�|$H9'��H��_*y�i�P�z';��ss:�I���&eA���wO�y�����NE�u@�fp�v����
rEkn2~򖉷�����}��1mˎ����|}��T����ww�,&�l��gP�5��M�ɋ�o�:
WW3�-�B�P�;��C�w�~��7�z�8L�]󼱵��:��]�{�1��Ms��M$�q��V(����?~�
�y��m����	`�[���P����z$0�
�A���5I�i~B<���ȿ�E�%��̜�|khf��`k����,�w@�#:G'�`�7��^�x	�����<ל��fA8���Җ"�]��0��$�{��+�QBҿ��]>S��1�/�>j�]׍�Ƨ&Wꖣ��'���*���s��q".��\F�	j�m[��\�9�ƼMzh|����iO�ͭ���Ր9����tS�CX���4��gޡ�ř�S]�3��bR&�J]-���q!N�s�<<�������(�>�����1��5'�l"9�t'� ��C��CGV���3qT�3+/��LTjT.�9�@b����i8��<���C�����⁌����Oei�^[�<\�cޚb�҇��z�E,v�A]��\�}� hd�a�|݊�6�͍�{�����HV�?s�y@	���:�,Rީnpc��S�mxw�P���]3�o�\�24r�}�	��f�D��EĎ�=/C�q��������|b|�TLs:q,���ڈ������x��b.Cw\t��szYI��؄`��\��)t�"-��]��"�Ռsg���*��.�{^�����]X�z���j��v�:���Rҕ�-�΄�u�UH�W	�7%���Dt�y����v��W2�{�xxW���3�����q"��L.w�������i��G�a����f*�� �5�ׂOC����5E
�5�2�5oiʞ�����Vã��ط��~l3�ɕ�W3}=��{f��쩣�M��N��e�}P��*�cb�l��A�9���:�$�H��93��x�\�Pեm���Ms��x�b}�T�
J��94����y��Gg5�V�!?��Ĉ�d!ҿ���_��Y��.���\j��=FQ}�1�m�q�����)����H)�9ഏw������׭U���D�{�#Y!�=�V��Cz(ϣ�8;�Y�8>j��1p���iM�\�.w#mj�7��!�!ܺ/>��z7�绮��%�*�Fi�w���=0�1*m�u�h�:��xi/,�b5����qi�?��;�N���@vA��<q*�SO�뼶��g�(a����c�+�+��'��G�q_,!e�+��.=)�|���]�$Ghؚ���7�H'���"�MV�S�H�51��z��x/V��:
͈�1 �a-yh��������
Fw����j��q�`���:�{s)��Va#��J�#:��yK&UE��McU�ʣ�o)�����"�+��?;�՟���nbp�& ���)�M܏���7	�{��bˆ�n43U�	g{�{B<���r�u�ty����=���&1�w(SdW�5�>���gE1.Tx˲2�
�XRu���t�N�DH�PN�U�Vl����u��r�jZ9���+�|�|��w���گ@��׆P�e{v�Nt��l�8'��7�bk^d�[GC�gDn�W����W�	�fy+�s�05�ω����53c(�9S����f��<��2�F��4%l
�F��ʒyưo��+._;��eS������n�8Do;��A��*E�_=��6����DJ*i.�����.|��f����7�bW��D����c�36��0�ܪ�(ϕ���XVl�g�C��f�#{c�Q�8*.�z�Ԙ��u�n�j�7�ޮ7֞��"�o���]�W������y�������#���)o�^����6{HO�S~���k��յǺ%0�e�c�	�꺽R����룝p[��<H �����kފ��M硤uΪ�ӽ���u1u�+m2^R\3_�Q25�%�z����O��7G��]N���qs�w�}ODo����"�uG�*�}V*(���$G���HCX���{ɤ�L1��u�=3��s��7O�/9o=��eu.O7���{��V�����$U��Y��Y����l�⭓&v��dv{Q��Eݸ�CwQ^�ze�e���Nf�R��6:��ѵ�2��{jP�9��G�]|Z�ٚ�>Jv���k���F��q;�㎒LG��k��^����͜m���ʎ�O�� 󔥪���,�y;��J	\�X���vf�4�`��bn-�fN��͠���Nm᝸�盾˻�1�W�i�������Hѹ)�K�-mp��͡pk�� �+O@.Yrl��ƯRK��*Sk,/<3!f}yԪ欸�y�e�w���3�q���qc��q
6+k�`����Nh�+��^�os-���+58�-��4���T[��L�8���E�q��5]�$e^{[�M_;s���Ib��qڏw[NAF�cl�ܣ�S�N�N����m��T�й����`6ܲ��}|��n�� ldӽ�8rYH��{��^م�Z���՗��]br�}�%v�)�F�N��]��7%'J����a�K;Z����{Vor��&��5R���2��	�b�r�~5!�fw]:WZ�ږ�C|.�v�Gt��S9�7P����t$quvr�C��6j.RKl1��f��oHj񞕰㱐7i���6��`�n���]�af�v��C�ͼ���_D2rݠG���%�������2L�7��B3��U�ۮ�R��%X�<7Ѕ�����N�!j�����<'�+Z��{���'����Nut��{[�`�͖������v;p�{�� �R-�I��O��R��m�_v7��������ﱫS���Z���Ho��$�V�����97145�&qca85�]0u�ȝ�\�!�¶��Y݊ܧ4�Ѻ"J��9�ER�o�ڢL����]-������3}���0
��$8�'�u�N�n�4�JXm�h���v�;�g�X����9�]�J��}��0�LB��yv�s��DD��7�G>�N�{
�<ܳ���cu��|���VV.�íf��)��x���^pm��t#�5��fXY%6�랴�E�)i}��`�n����:��Y|&��6���U��:�miեom�]m6�{�Wp m�WL�;N$&�tGk-�;���6�m��2��]�����;�;9O�+�/B
�7cV�E��xJ�+�6V���c���8�3U�#�x�fV?����?���Xu�mo�ye�o�u�p��q�^���X*4HIl��[x�O��8�<qǯ^���nݷz���˩����FIۑ�������x�y�m�|��{sn���8��班<|q�q���z�>�v��zd���;jkP?��{�9������$������|�X���8㏎=z��}x�۷�쌟u��N��[�����>j�V��U��s���D�u���ك��''�i-�8��Y��6�t>R�GG���'{ޯJO�]���>7��@�'9p'֝|c��
9}��=���I���G������}޼�����D%�[nI:��[d�¿��A��}�;��V�5�rN���8�ƀ��Bw�GL�YvqE��rJ%�W��'s��Z�8_-d����,Ήm����I���%�ݲm�Y��՟���E[m8��s�e����(�8N��Z�pc{����_ đĔ���P.Ȅ1���H[� �1�����P9'�&D�xA$�P��钷��t�qC9xi�uv�+W0�Wui��V�Q���jSX盓��{]B�RuDy�����+Q��
M�bp�D.�1�����@� 
@�l����O f1a�PhC�Q# $�� L2J$���! ĒMĜ���Cf3)�P�Lm��[��<EBT���4\�UJԹrM�#��,`�����H&A ���8�6���Μ��٫8b)����L���X�K;���t^Ϯ��!���������Yꚽ5���_H��N��޳���}}�`�ց�mP�247��03!-���D��KL]V��}��k��^r@�	*^�W+U>�}O�J�i��G4ftFF�2�7]IF%sCJ���k�j$�=�yz�\���x�Έ��7���:7K��]�Q�S��o�Ķ2�g���R)`�>�*ɕ������ezݖ�#��_1��vːu�ƥ�w焣�zU�k��|���,琇q��j��pN�.��\�|�C'9n��� �s(�a�.}���J��w1��s�Z�C%�j����i$n[sע���f���h<���Km�>zd3�v�Ϊnwf`Ι�4xߛ�H[~��u��!����s0��ືjc"�1���ֺ�v���*�v��nK����N3�Ǜm5�A��̝�$��I�V�B�0�o7j}����P�{qb�j�·gn=C���ץ�A�s�	,|�	C���θ��n��7v�\X��ٸs���(���.��]��Jp��Ώ��-vn:�]/o�)�0h��ߍ��{���r�\��):���^	H��:��{�rY��O���7��s���XT�z��}���y��6�l����Du�0���4���=ԭUs}�j�ߠ������sz]jM%8��=ߝw��KҖ�F_�=��>C�ק����.������LJ}�4͕rr���v�́�l�̍c�p�`Y�xܟvH*��y��E�x������l�6�C�lω~�1��q�F�:�w��yV�[��E�i5FRu��"���+�j�ς$�KA�P6=W�� cѨ3'.�3}��I��p�;�~�"&���$�?\K߻��.p}J/�����QJ�{�tr��ĉQ��{�N�be�{�vd�ϣ�0�Y�E~l�C�q�T��M:���΅S3��:BĦ�npUC8��)߶)�@0)c;�{quTľ�[ md/^�Q�"�u.��U	Q�?Rr�ng-R�r�.�z���Cy꺸S�K{I�����Z�w�{���b�;�C��m�kw���>��[��Zg�2��ʫ�N�Z��v�QW>�?�x?��ڣU�y�l���*ٝ0�+l1�vq-�(��rD�����cQ)� H_;9y���|�;�%��y�dq=��ESP m��� �g:�#�KmUN�dJe����}�\�H;˺ �r�)2I8���]_�`�pl@3:�jp���uӽ۞�O��	QIn�%��c��f�mv1m��ms�}�ы��N�~D=����K��u"���+W$L�/�b�R�����#;�c�ٓ���KԘ0|��l;�1ݳ���w��1]��f]��㛅��z{&��{ƭ d�>�`-��a��̟�#�ʛ���ڻ����5�:ݝ=�c�W�<�j+i����[>�7��#�]p2�-K�1����/�t�tk�s�;|T��li�7�Ǝg!�ayC-�ؼ��i��ɽ�wp�Ӧ=��m�j��87_y�P��Cw;�"mi[��b�^���>�˽���R�L<+5�)ŋq�\���g�i��bK8���T2ƮU���$�;Z�9sN<D���۸eݬ����3�l�^��GWѴ3v�s���d����!Sa�����Z��߱�t��8�:��Hj���gl�r�^��u��¾�� #98�k�\�]W���{�<��O��~1�4ƈ�d �$��y�7���s7acw�_H����$�n�'?��9��zǹI����8��wx�l��oc&�dmzYԌ�X0���R: �����rAY-մ:��p���y�2��8�<���o��-\��8>���� ��Y?z���ߔ�CKZ�����Y��9�/��P'��^��ՠ/f�*�U6S^��ͬ-"!�!Q���Z�̑�1V�F����Q�P��2vnF�B�_5���6��s4�'E\����h�]��H� ۬�y\�I$�~�ì�����k���;�O���j2�z��3��_t{�T�������l���}ܶ��-�{�+� Kf<m�A\9_��za@�`�s�K�w�<�"�����v��s�vʮ�s��1�н-�Ϧb�����J�}�tj��(�%ܻ�%��V�0`�.w��?��v�c5�|�;�,���j(>������.(��n���z(������x2�m�
>ߨ��h�,+ิ����
��m���<7��5�������i������7M���VR`F�=\�Z�sض^Y�Wy\�K��Ɔ4ƒ4ƕ�ߕ�~�b�f�����=�:孨v�v5�]u;^�C
��T��.%B;%]���Wc��;���JB����Th
��g�Ŝ7���D�j�/lQ5sf���)�v�Fw;;��ډ�tr�b�k�uQ��Vl��Y4��+-�r�7$�i���fj����1�"Ho|�s1��${|ڋp��xU�,���z�T�p)Ϣ��溠��T0g]�t���cv��F��=��w`��rgZ$��td3�т���R�H׼�S	��ζ��:��YO<�x��Č��h�,�@t[�����Q�=�$^���Bj��5]��n�q�� g�/c	�\ UҝV��S��W�ڄf�mg��=�h���mW	Ϭ�`v��:k��z����
ysYa��1��x&���E��٭�:�B@�h�!��R3y>���0ёK���&(^�ׁ�ч��eD�ڝ"��=7�x9B���Vy�R��0w����N;L^�����{т���v.��Q��(���n�7g'�g|��[yD��*�fڻa�LBj�8�v2�0�^*Ts}�A����!㴫D1H������/j�,{ՈfN��]����WJ��6��p��NS��N�㝭�^V�{Sz?�����i�!cB"H=;�O���{���>�U��F�����F9]s(���%�;����62`�8;�d�t䊱�~�N��l���̌�� :���r�Pٳ�&2�u>fe�q�V�R��my*
y��w��P�X2�qmz���1��>��ݶ4Cy��c/������������ԅ�q����9T���ԧ�q*��.&�W�*�ot�5C�r���T׷t�[f�;_��1&9Ǻ�L��?�#�v7��4�tq��V��u�q�z�$V��c�_v&��i��U����`�xf��R���;���yW������N�_n��a�$i��n�f�3���'˭�3�@1�L8E܆����}G��1ø��T���s��2��P@�,��b�O]mڽ��:�ƛe(��#b�s-�wzQ$q-��ח���[T1*�T��ݷ��^6���Ϡ����GLt����ð�ˢ�0�ـt=���j>yڰ+�cB�
L:�Um�{o�>�Yd��,8V v;jWG,����_nڸd]�j�W���t��9�|���7Nu�������~;h
i��ij2��wߙ��+Y�^���>�bj~�v�}�#o|{�������q{��;�Bi���q]r��C8���"}1�U^��6���� ݀T!�J]͚���Φ���u[���4� kK��	��!ZSl/��lŉ�����Q�{)��G��:{2ji�j�gֶ�C���"4]�j��sW
�v�FЏ���x�B*���F�(��8�֑���n��Oqh��t�T{�l7AX��������^l�����Yxz��g_��kf88:����pi�����&o2��=<5�C��`|����`ǯd\i6y1A���7�ö��V�lŝ��KT�J�����n���{�c��=�3�E�@C)/�8��۸���%LSW]�&��U<bj��#7���r��GZ�4��m�8] �6.3��秷���.�h�W����]7�7����i���K �>�EJOK�^ߓ��j���XRv���7�w_#о2��k�݅�o�ܮ�>�$�4��h ��@�G�{ gl�<3ie��)jZ��$�d<�ҟ�fuרT�
�ec�망E��)Z�	P��t�m�����zx �o7�Ә۱�Y���	�Q:jUP379Kw�G1i�.��G ݡ�k�o�<!�^���v�:�|�yV׸�خ��������i�;2yVj���c�^7�Q˜u��_[���s{�m�ݴ;D�`��o�A�LD𨌛���� ��8���^�>ց�`k��Gv�G�vp���]��(^J|�p:�)+��.a�hB�� ���w����g5����E�ZTU���~�4.��p��*�w�Hv�A�5Zx���-��a���f8vh�	 �J�G%�6��+-@��{���ӝ`��F�ƙ�V����/�^[aj�Ԝ�=r<ٓ�s"��Z�du'��i��]�F-}(߱	�Gnt"AF%B���V�Tfcmd=��P��KF��5"
��K 1G��-�I%!�ll��{��1��K��_~DI�V�*��W���y �иWh�ubS)v���^<��o ���A=+A�[l��J8w,}i�G��b�d8�cy\y��k���ּI�����qK�v��JsW}�6�{�<<<<>ϳk��G�T'{��u��tֳ��ݚ�ګ8��l���s��m]��셲�����Xcm�����賘}}��)+n\y�KA���`׸^�I�\Ef%@�lǍ�A[��n�9yZlm�3NV����������]ATR�[Yϝ�������HDoH�M쇶+�:��~����\AÓ;s��^�a���[/�3]5�`y�~�m�u�>[y��Ի��f�mS��)�MW���{�4w���͖����T�~f�x	�*���<-$3!ϙ�}tak��ڷ� ;���r�M�K�%]^[l����ϯ����&��(����GGl���;I��ɱ���Ժ��:�oG�_�$2��?�gU����to�Tc��&�ݚ���$ؾ}�8�lR�9�����C���׫FxU>y�U	�̱�� 5S��r��^@<U$F��唳���y�	5*����I��|�"����qY;L_b�˴���:�x���I��3s-g[BVtw�^�FK�]o1����E��(�R�T���{��9��k�5�t���u���8N��$�;�n��2��1B�#��WoB�e���tY���C�K���y��a��(��QW@mr��M�Ȼa�� �P��hO���M]����d�M*�lS�M����]N�2'��h���eB��"Ϯ=�o�Gv�0ib$ɢ{%��o��/[b��}�Kz����<n�2ň�w�
�#u���Y&�/R�'Mű��z
�-m�=�5��oZ1OL�����*�����u|�6�42�p�(*��!q|��x·�[��fD�)]��ff�tx��D[�Լ<�OeTM�'��Fw_��J�<�����j�23�_�B�Ǔ�^�`�R��ޮ�����bH��$RK�&���N{�ϖg=�`#��Ub����������%mLn�3���h�T�t���;,�#���'V����q�ݔ��I����B �=}zk�/!gr�U��s��:ڶ,��-����nyD#P�K����ٕ��N,�-��{�Xu!ӈx�[���Ӽw�̾Z�o������{n�|*4�8!�,�=4�t�v�Gv��!$�Tѩ����n1������쩺>Qܓ��[Y��oe��Џ���fIRc�%�#��W|@aCx�Ks����١���e��cdf&w6��ĩ�X�%N
�n�rS�X(e!���:�(���L��7��C[���Mொx����f�6�Z�%]�Π��6tf�:s���t΍��4Z�z n����#I�S�[����l�&�$�V���.���&�Zа8/gqۄ��.C']�؎�1�f�ˎV�59�Ұ�1�Y]�ܥa_��s�8���8v&t��9���l��əo �s��d��g2��kE��Ձ�]��Ip��qo)r�e��z�y��<�����p��s�X���ܧZGdש�^^n ���mK���i�Zu&]���i�x+�T+8(b�*�� ;p����m��:t�G��c����0Ut����к1Re�K$�9�,��W���S�B���w
۬�cm�eUg�������hX��LZ}f���}ݹYi9]{��87��خ���i|���~T�[V���b�gȫFEwΐI`oTs��A��ʐ�}[CJ)���>TNS�q���;�	��F7�턓j=n.�{a2�x��1�Y&�$�fuU�2��d���&fe
+�����H��
�Ud�v��d
X�g��.V�>�� ��Tv�,4����9=��If�"S3:fIB�X�s	]ms�Y5��4�LݵB���9����oK��l,T
��F�c�G���:����%�LN����v��R�F�U�x:�!�8������޽P���K�Q��{��o-��kNP���m��c����ӄꘇ��Ei.����vI��tb<hP�ú�x��}�]�#5$CH�:
,K�]Ue�[Nv6�"����a�[Xv0{/Fd1���;n�t�g�����A�QP���:��}ZA��1X4�ѹ���k-f�s���D��{����`=�^,��]�l��0P�7+��56�o
jb��ܕ����7��R�ͺ��Ua���w��2鶌!"�ʻ�g��.ڴZM���.��]�+���[Y]��n�=.���V�@h_���ī���P���G�KR>4��4��xFR��`�\.��7����Vv<�oP�L���́��A�]5WeӜz�YG�6{hMݷ�]�9�{���]�SD�iI|�ɱ�%:-��^P��8�/�#���7��4�[�t�{O�F*�����R����չ�k�yA.�/�2�[4rշ�3�J�Pt���6Mq�
���b�r%ۙ��h*X�
k�U�΋4sl��8��36;N��'~;>mmdPBI$����oX�����q�ǯ^����v��	���@�
d��D�,��v���A˽���e�۷�^w�}��~���;�q�q�ǯ^����vֵ$B.N$���ݒ�c#�(c�P�J�
�UH�=}}}t����q�|q�ׯ���nݶh��HT"ie$@!u���߷���J\�󿚼"�K}�rƶ��.[Y�n�B���I�w�k�����y@�;;��q�6�|�v<���V�����͔�ʲ��q�ɖ#�����nӄ�%�!�����(��ye��y����ϫJ;��Rw[np���੶@vvE�h���w=��~/�+�,���cE�y_�k�C�[`Yי6�:(K�+�������Y����O�I2b�.�g�t����a�̒�_0�=��ΛM_��~ד��ܔ��/;�]�N �������~Æ\����15��l�W@^`�9��a�*��/ ��	G���Ϡ�=Q�w���1������o{0�L�687��������+O`ጄ�sVr�7�c�&߆��,�M�^r�K��=:m��O��P@-�3�\�Rܲ�U�<:}��EZ���a��$�KAu��p��Ը��8���w���jx]�l=%"&���������ikc{�6J�V����\�fR�b��.�(m�I�����t	���s�x��1A�%�KN�d��k�e�?H�g"�PF��+J��N6��mg٫��c��7�UiJ���U�չ��c�edV:2fZ��GL�����A OC\�C:
�<���_nϨu���x
��3��,z|k���Xu#�t�:���Ot{�G9]�L�J��|.];��i{1��<:���ի�1L�N��j:�s���_Q�]��e��e�]��Ee�k=U��s�_[цE����9ܥ���ī1�M25�FǼs)�8�dl�.��7]�!�So-����ӯ�ae�^g]s�;2�y��o7�[�aי<y3 ;{�lAo�O�&�#v�+*���<�7=����sq��{��^��HL�7z��Al���hY�M�ޥ���O-:�%Y_�4�?���&o�N���|���Z��)�l �S�n�j*3��j��l๹��&$��6��-~�v*������Ј�jV�m���b�>���vusǺF]�pf���
&b�T�e�s셳�b���
��ˇ�c�W��ck7�m%Ut+�9#_V�=��=T5ﺨ�ȴ%�H����~���G��>!٘�:�9���\z��ћͷ=۞�s��bF��t�Ӷ6z�w@c�B�p]xVW�P���<G%�')��+4}�O�4|����{��X�9�y�.P�k�O7 Y��3,��w�Z��;���$�bD�	��Y'^_�E���E�@7GV�x�լ~Zz*��]��:����q]ǧA]�y/��w���eg�
��rM���eDj��X���É�,���eIU o�R�c���έxZ�W}*����ϔS-:8u�i��A��j���;��*���������eN���gֶ3������N��,����������������L!��I�[^J�fe�}9st�6Z�а��6�_TCl:�~�n�?�Ĥ^>��Au(2	�v+5�q.f�a�x�27_Wu3F����j�D,~7劮��oVt�EU�	;w�b_��n�>���/1��#g�Ԇ��)�E�l�����eJ֗ö�>����f��}��H�UqU�uә��t���D橽�4wJ��,V�a�@�w�v�m�1��F��yu�e��c�ƾ��.�P�6�[s�{��3f6yn:V�JW#�Z��3õ���^~��&�	����\�J�~�O��y/�Bn�������ČPK�v>l�{,�kk��by�UՈ�����|�K�u�S���Uܒ�ޞ����������I�T��o�:V/ڤ8J�n�FT�i��V�^��F7�D�4��DU���Yb�i۹�֡�ס�Zj�������x6�8�9xVW��|{Ai�Uڻ�MY��N��\���RG�I,E�ӎ�{���aR��I+��I���α;f��'�73���$�N|�*�����"��˝�]�����TL�(����fSR���y��ڗC4�Q��Ju��NtM�t;�ܻ��m������{�2���xq�㵇;>hX�B�T2�ۣ"��L�;���Ջ��%�_c��n���Z��YĐ0Wl�g��: `�g+���b;�`�LEq '��y�j)?�fϭ~��)��gϸ`/7��SSL�X�ڝ�U|N
����qW�5OX�hnp2�����%"si/V���f�I�k<	��{C�_kV�5���8��ʨ�d�Q�dg����x�ƍ��=ޱmsV��������z~ �pW!G��R5cf�Y����ϕ�!���m�1���"7R��4�=�xBz<��d)�����N��ʨ���T���r�Q=����O��r���d	�+�%p��0Z�>����`l%o��a���yRSx����~�'ꌸQ�������~�VJ�`���V&O�N��.tC��������g8�y�
C�X�1)f�U��z�Ir�� s�Ծ��ys�^^nS���Ef��gA�ywO)x��p����[t;�V�ө�Y�f�S5Cd�s�>o7�y�zY��&��y�|�'WXv�2��@.�y�A��a��m�;��pυ����<X2��/��.���w���B�U���K6m*�'#;U��WGsr���(�l�#�����l���w�e��L�T\i��"�a�����rVxl7�-����mo�%%d|�-Ν��7Q�h>�8l���;&ہ~���<f����-���^`�9�]w�b`�2jnUA�}{{����/r'��NV�������4���>�8w���_C�A�n���Z����>Q*��%�>��gğA�G��Psa�'�(q��7
��iќ7Hw�OU�pc���6gv"H�q-8)���I��u��I����n?���o_�_���*mr���瑷���"�ٗ{T32��LO޴|�wȁ���(oW�K�h�f�c=�����d7������e���ج�`�r�{1XN�dV�Ú1e�n�CN����yP��O�'�֫�K羢(�]�0Q�7�&}��L��ö����0u�=�ܧ5ʻ��b��ʱsרv���k��4�����p�>��C��+e�xs����M���i��ת�W�Y��p���L�-z�N]]�N��gu�U��EU�)�V�r*i����Cy�l{'l!,���&��k��u��jj�q2��G�Ǜ3�P'����>�϶�D�y�[�.8����7�KVHӼ#{)D�r��ך�IM�y��.�OJ�gE�i��瘓N:�`����ln�%|��
�ypٵ~wY��9���'�����d�N�}[���E���V���c�Ȏ8�3�����u�1�B��(�zh�Ӟ�-h��H��X%����v)i��=�9�χv��n��h���J�}�k����ږx2��Ug���1�x�(�Brfnqz�w�sh��[�����ᔼ�;�P~i�D;'_P��[c��=������(�4v��g�z�R4ӽ�;/l��m�Y!mE�c?}�F���)SO��0b�/�7�,M�wו�L �ݵ��#��O5Pve]}�'x����C	�^�$�:��Nfe���}T�׹��4�DU�R;�\�K�b�ӻ,�S�ft���z�*����y��Ȃ�����ߞv8��m��r��[�h�J8&�ŉ�*u��;�f,[/h8�j����*>0�ӵ������tv�u[���g1��Wu��O!T��^�$_�PD��\��� X���[<�[�U1ʽ���":�t�a�:�,yu��B���I���w"��,c9�ѝ�ǅ3ːO)Fȝ<�YD�����0Є��~�Q1-3�".��MnmQ�l`�����\���<��'����ڛS���>x"ᬍ�R�b*�UX6Ϟ���U�!Q��($�#�u�Zr���n]1�דZv|č�![�����_�ΒJ0�к�Y�Z7�&�{p������~��'��LK�'4�ج�^9,�49੷�ͥ.d�<��v3xϣj�d3�t
�]��
�����t���)��_qy�w��;�!|��|WLN�ƀ�g����E���A��r�p��Q٬_De��&�{hT��<��Ú��	
�[�+R"��ղ�A`9����{�nAW��Zu�.�mz�]�y4�ф ��e�<E*�N���}6�!͈t�Mf����sq<�#{][�U�)�c+^EV�(��w�
˪������.)�1W[�cO�P���K�hZk�v75�V��nL��� 6]�JIWth�t>t���F�gmL�D���U��k�������-��~4n����qp��k�a����a{���Uܒ�ޓ)U��#�Rqdmvч����3s��aԈIy�t�J�L�i�ڳG9�W�'7K[6�v�Z�����k<·́0�R�X�v���L;s�m�NP�j��ӧq�il��ff��*C����g����4�pN��A)]��T�z�ݣ*����r���#�A|OὯ�̒w������6���p�D`�>ZSN�Qqj-��Z�S�E�һ�ל�x@�nM��~�2�-��5�j�ܧ�'@$�Mv�U����I��*^�vy�2�<�ws�	��j���m2`��|JY��ꧨEǗP�Ԫ�,�5�K7c퉧J%��V��/��W�bvW>��0������%o<fB�f��f�_q{ ����9n�̾\;�T{�t����������o����̲�0n�S�ӎwb&��3AG5Vr]��B҅[�ŉ|޻u����.6]���k���{g��=`�a�O;���_������w���U�13�������^n�&��rv��݋܌�=f������UG��藩�p��Pmұ\*��+c�룳�5G���^uWBJi�l>��o]ّ!��Jڥ��\�11|_"w]
Gg�Hs��=ݭ��j/���\�����}!��N����;{V��;/G��s�aà�R+�� m�*O��n�>��}���%B���1���q�xql{	@D.�=E���5]������{��I-�ٹ���XOv�M��m�w%�����Nz���s���"�q�k�6��3Nt��K���z���o@a��룱Q>�4+/n��m�h�<;OE_<������ԯʺ����G1LÍ�,�m��=J������}!�f��z1��o`�7��d�h1��3�Aj�m]��/	�ͯʞ���S�u�� )�Q�=�s8 _��Lj�j��7�8�M����v
\��Wa"̗9,�����mv�UǏGn�!-\n�9W�뮢��B��z���FS3����T���;Ձ`��"�#ܷ��ٝ{�������y��o0�VK՞<8��WP�P�D�ޓ<X�6;��s��5m�m�Yד�K!�����GZ�ڌJ��^�=y� �!����q��ݧR�n��[���	>���4K��ԕ�������|���#)?ة��i:�{���,=�!&��~���<���n���e���y֠�
Uٟ��yf="�}0zЭ�a&�1��}n����~&zjl��H��I�UB9'n榜�/c���o{�]K�y=�1e`Ȼ����p��%�S�xv�PP{��nCgx�Za]�O�>����]�2f�w;�!����ǥ�!G�w�L'��p��q�Q#�'�RdJn��_#4�R�-Q�t�L6��H�1Yq���{��X�|���"����Ěu�����W�6ǚ�� �����r����*�+�����G�2��V]32�<�:�;�w%��U>��7��7z&�[M��Ŏ���f�CN�秢�*'��7�b�;����ՔU\˛���
v��^��]֮��)��
�����<l� ���X���
��NXb���v��wc�mCv�CӉe�'�:
��oG`��;ebU^��g;&ª�Z��G�3�v��u��ǡWܤλ�ҭH��a��u�O7�so�Ô��/�"�W���1�N,6��d���
�H��)5g���ӳ[��P��;*:|s�����0�v�$��4&wR��Ԧ��]'���5�Fou���*eb�r4�v�[��܀��c�.��Q�ȶ��K��-�2�Xi����w,��F���yx���b�T9��&�$��wI��#��ʤ��ܥ��t]���\��Nv=.�Ӓ����x�w8�3,0�:f�-7���	�E(�����ǭdVQEnX LM��{��k���l����w�	�q�h�.�m�NNm�oEW`ȋ\)�\�3�Z��21˽7f-0��X�yc�/;�ԼV��M�{O�D��U1�����v�O�c�7�c'eއ�(����3��T�Z�L���>r�p�S�`T�ה�*͟8���ZP�ۺүM힋�TDZ��ko�o\����֢����:��Z<��:5t����*�Q���֙�Wm�B�(L�:[#F�\�wbnX�UB	Lm�;+/3��N����P��F�QB�v@w&5@�P�d��Y���46,��Ҧ��;�e9��P�̷F����
.̩�cz��e� Q����%oC��/px�4ַ�ck�Dj��&wޗ����o.֢2N	��lI�s���჌㦡T/�˹PI�{5y��ԕLL��5d�i�JM�Y�ig���\���~Ϙx��WA^��)��ެx�$����b�1@��s¦V_g:�USDa����L�t���ғ\�;�T�3����Y��]j������,���QݭieȡW�D�3f�S
:�\��-O9��u�,��v�D��*����eJ����o7ٱJe����ЗA[�۪��+:�ɷ�����m��lsӳKoÜ0f�D�ژn�N�W]UJ\��<��Z�A�u�Y�-)�f����1����F�JW����f��e�Y\�4��S���f��E��FE��;r�K��vkS@��@�i`�J��93c�N��ר#�����):I�^�&k�+jD#�5�7|;��k�G3^j�A�'�ł�y������f�#�o�76u�Z� �w'V-���� ��Ŕj�h�z�S� �ɜ�����t"SΘ��' ��<-��q��\q־]7N���#�u�O��ۥ�/n�W;��xls��1H���Q�=�Y	�����R	�(y�I��vjvYŝ�h�	 ��	��I��z��������q��z���ݻv�L�r��dqͻ �n�6N��dpvi�'~.�����੩�׏����q�q�ׯ__Y�{�}����8q�@HWŐI���Qb0�aH�����>8�8�^�z���nݻv�2���Jp��D^՟��DxۿJĊ� ��?l��܄��.H���$�+;���B����:��Ӡ�8B�9��vE�q!�Q)p/k(�"�3��+����K���"�����I)|ݝ��ݺ8�+��yV�B\u$�~��;���ݠGr���yF���[n裸����]�gYqg�|Y�n;�Ό�ݥY&e�$Kk��X�vYD\Q�w7�w^w�����_�ib�h!�!@�Q@�4D	��#-��&G8�P��|�$�A�B�����;��ՙ�.��7������t
z��}8�8�7lr��{�i�/Uݍ�]��&-�võ�1(K2@�JN��e�#h"	��$mD�8(��B�L6�E�D��D�YH���T�.٠�l�!2AE�NHJ%>D�F!H��&2
$d�"1����"�}�p�xxxy���c����ðK�*�R�ݹ�N�����-�Y��;��}�5׍���.n����\��#0/�w����cp�w(�w������+^�\�q���j�TJ0��M�2ո�z�oj��,�1�B���~Rb0ȅ�S�����(��jسU�+po�fq{��ٯJ�۝</����8˰��kad�����I٦�X��1l�	�k�g��6�L����'}��\�U�86����G7^Q{�Rq�vJ�������/=
R3=b}� h=`�u\W����X�c]s���n�Ռ��,漣yz@���8bT��}��K�A������Aع��]��ϝ[������G�^��+(��?NK=� ��ވ-/m�NF�7չM���|�OT�������&��j:ٴ��L��F��%ߛ��VF�,4*f�=ܫ�5~|D)H��M(2OZ�̲�`����-�S��SN�ܤ�]#�ṹ�o���:���T�}gf++%�@Y���^rCq��KRd[MK����7KWJ,�y-�u�s�^�2�grۢe�s;&���Q�NKF4���o+OA8WfN����ه����o7����o�Nt��c� �
� �X��n��z�t�@�*,_�U:{�F�έ5ws��M[<�N[�.�Vh����H�-݈F�CK�D9��#���]IM�}t�FߌH9�9
&���ڕ)�`4��r'6{���i�1�����#O.=gCfg�w���h\�����-Zݕ�p$����Y�i)�9R�`2՚�ۧ��ù�<�>��0Q����s�lr����_l��؞(��]һ�Z���/�������P���;�O�9����Ly����5L��o�}�+�3�*G��B�Ǽ���坳hU6�Ho[����Q�;k�n��Wq��e�Z2������j �d�h��po1�^X&���ȭ�5RU<B���ͽ:��1�\��:|v�31���y�=ze��zr��_�����b����/%�z[��&�Y����R�nھ9^�2w��6�y�	��8���=�n>�د��|G�~Vzya�x�s�9��sWS�PS#rwۤ�g���=4ƸN���ip�!`LN��sB�^�.��`F1���|3=�x�{�UU{RP�=��R7����9�<�zߤh��Y�4���R�\�۶���܀xΟ<��i��<���O���2��mP1nH�fN�3E��(��z+{A�9X{��n.���'hnp3�	K��إ���B=�&B���w7��~�|�~�zю(2N�S��M��U�Gf<nRs�(LгŢ�.仵���Fo��Ad���g������tL��U�4�8��f�fl36Ys˽G���|�ճ�jt�WY�{1�BU=f�03l�Ļ�s�T*C�+�q�R7-��dH��0�-�X����3������Q�@��!5�nW/7$���%	;~j>�y��J�b���޼�nm���F���;Q�־ r�>��������R�}�Rم(�3Q�ÆQ�K�V�<뺀1���W�+Ǧ��	OF�c�����}��3��Q���5\��mm��W|vd��`s/1Jv; �wW7���k���y@�[|�qgR��۝�#��!�˻��<���[K�H�N-��{_#�7��[7���{e�)b����$H���r�nhW�~[�1��bn.�s�Y׫�y��o{�6�	�=��4�f��k�m�68`q�odAo&�'"�X�{�|n]�a����Kv��)BN5*�*�wQ�,�e���F ��`{�=�j���|�^�yḍwp���ϯ�}{�>:��(�����f��#~:ܨxok��1�g�Ztd�.,m8�����*�jޠǧ4��������d�c%��Ħb'z6�]��a��Q�1f�i��mɭ�<[<l���v�[�Fl�o)r�KƖa�agT�*���e�6�� "O�g��u���fue�M�&k`�2;(���b����O��kW~�7�+�o'�~�4"�V�u�s_{՚�3�7�_���gj��̎�x��f�%�|�.�]�S]�>FƜf��$v��e��A�$�ן����g�A0%�E���f1��l�SF�%�@�ҵZ�5^�%��ٓSN�زɼ�������#����6*���0��(:�if��s���??On�����͸P��gy��~�M��1aq�
W���1$qI��r[UHL��dl���z3'+�r��or&�,j�8�p��X΃���Ӄv��k���ݗ�������>�q�$�c�!��.�]���l_JĻ�0=c��d�#���T��d�u_?���1� �o,��GM��R�eJ��*>��8���g�/A.���w ����q� /;�'{"G9Kؤf��g=G���1�{��l���k�S�K��#A��n�o��ԯ�����Cbӳ]�60����<Nm�� ��,}[\�t2�;}ݽc�a�01�#��F�g�׸�괉����3����,��7�֗.��L�=���j�Z2q#��(ī�N��.�l����ܳW-�k#�;wr�[�򑪤D+�c��M��
&���f�V���ХZ�WH��0ÂT�0l��M��Y#�����3�Ƕ�l�w�,T��i�ޤZH�nǸ��
X72	7R�tZ�g7D�K��X��urw���kd����_zCP�gwG�#�xY6"қ��g�]#��Z�^Va�O>�k�+����F�ܾbm��Վp;�Bm��!�b_Q��1Wn9N�G� H�����>���yW��U��r�Iᅡɭ�	K.�؀l�Q����=%ܳZ+^� ��DO6n^�7����{����34���A��WH��#H��$��큐΃���a,O̻�a���uQ��)7��^oWO+#O6z����~�d���*݇�M���v�𚜙�gx�-{�P���.�-�o��8�z�m�Y�S�U����.�3�u���bB����̋0ȫq��t �Ԡ�=ktݹ�'�oG#�S��E���a0����U��p��#z�FY��0Y=�n�Fvq�ɓ�r5[��g��9��#�:(�t*�S+�FGE��}؀�����REU �}r�Ƙ�@(~
��`Xa��SY��%R�xP �XeT�'�^L�yu�-���Agi]��a
{Q��b��r�0'v2�)�4�ܱ�C-qєvz{[�;M)���]SԜ�I}�{�#8R���#�dm��[\R�d�s�Z�|v&b:BRZ�����,j���6�k�|��B��r|��Y|Gf0��q����_�Ԥ��@�Pw�K7n�|��>���_]�}�=���u�����n��&�S��g�T:񞭰�h���` ��Y�S\�_v�u�������ޮ�.��O���������������rb~sa�y���I^oLrshh<^��G����*�̖C|�F�Y�x�kU>ͩ�};��(nʆ���*��V�ܝ<���K���>Ƕ��8.n�rͻH=�;��X��qΞ�����	��;�.��ǌ�1�σH{N�Ԝ.z�����V_�� �}(��x����&��`×E�k��n;ŷ�tTο��r��\�==�tLOyݡ:C��R�&���u�>�&R"4�@�����B��M��Gd�i�^�oAVլL�`s]��W55I��(���!����[���\�>Uy��@�;�,���.�=T�E���J�ֳ]hp�SS�g{0k�3 �(��x�A;,�+���R.8OSH�6�i�sUe�dC�w���^s�\��'�q"���@Pmc2�&�(|헬�g���|���̱w+%��|Q�[���8ޓY����Ya�����J� �Wxc�7x��F3jb}%�g-Jʓ[ꃶ�a�i�[��m3��N��:Ԭ��U�\�7���)�Čc��{����sޞx���u��ZG���H�x�]F��sP�Uې���|��k�Iʘ�ff�(����H׉]m���^��Vې��%ɳE�L��;���d���ַ#υ���r�(��t��[R4[���B��<"�{�����{P!\ypU�M�v��F�D�򚙗����0w�w��u��w�-��}���C�ި���?Z�虸�M���������g�JYܤ�ݓ`l��a$fǘk��m�.�g��u�2���툆w[�OW����Ǖ{lr�j�l��ti��X�d:ޝA�d��W5�xe���I@Ļ��E���<:�hgv�8;���\<�%T߄�T��M��|G5�����(S��l���c��t���8�]�T	��&����ԃ�'�f<��/^9��t�s\�C�]T�WK�v�;����^��;�Ι��}������4�WV�x��ӌ�GeV�8lE���-b�(i�+����1�x 7��=+K��c�ۗIt��*\38mЌރ�uh˗[]4C˙v��;�ݙwn ��y�_vm�����b����u%*�v��]jp�x�^��шm�س��e2c�_���G`�hu|؁�L��zI�_8���{|m�<�R?~��ɯ{�4�	ؚ�tS�z�w ��BPnIw�Σ�_����ڞ�aX[�GiW��p7`z�=yfng��YЩ�Wi��7Z�ٯwZ#2�I�Ӄl�M�RZ����સ����Rz��X4�HOm���3�5Uqh��xgw$���7 ?
�"�G�τusϒ�Ʒ�\�t��6��B���{d��٪n��!bJ�5���p�W���Y��*#6٢B�ͻ[gz�i9���vT��s���.QU�uT5�����݃�:bR&�ȡЖnv֟1m�n���N�َ]�z��]�d�^�:vID����oX��u����0�:^ɋ���X�}ޡ5V��y�����D;������o�A���}��ÌGvS��x��� �\�%�Cc��+1�H�WA
T�[DJ���Z񁓴K��M�W�m�v:W�+u�J�0.��Νr'ͯ�Օ����N;+FU>tW
�b*�n˦�ҝ�}۶����w_%W^e�tN�y��o7� (��˳�����]���K��{�O���)&���L�)���r.�U���ӄ�B����O�	0�o��Q��>��|W@o۶�̓o2�V��F�b���D����A�:��c�wF<�#-̅;�#�4Kn�ŚZ=��ƛ���]��^�g#�m�"ά�	t���O(�f�~~���Fk���<X��6ؓ��#!�h+����4(�8��K��b�*�	�|��B�+"F�h��=���<�7�OG���ZA��<���(��G�%"Ű!O���,�e�oeNF.UCLN\K�f�45��2�0+G�.i�\�RMX��* �
�� c 1����=�xsH�ӹՉ^fM�?H��/+���E[���߻�v����d�������Ɏ�΍~�>;w#U��
�x��Ԉ��O�8
2d8ך��)TY���XB'�wn53-���q�陪��x�r�"]+"�U�&L�N��#����ʡ��<,T�Ý\of�-�y|�M<X9��]����bb�<���z�H�D܎�W-�s@R�ze��J�Wt�WHa�G�%���V���[xo�wY���z	��hNI�؜��	i���Y��Z��]l̐n�I��]Y��P���8#3�y�Z���ZC�F��w9��(]�9����F�«�#�&y��3�sH4j�����TVj48��UwtdBu<���V�NN��/�V�U�z�ش8߯B�,��7,۷OWJ�g�\�|�=9;�b�mt�y�Hǹǘ7�ҵkq���PJ����es"v*9N��	W/.]vvm�m̀���u�^���{b9�����׀�қu�Y�/�)$��F�;��g	G:U�[�@��n���Yg-�@���}xc��޵�z5�1^�k�����s���i��%Voγ ��Y�Ԑ��^,���ez�nMDA"�;�[:b i����Ř-��uhդ�k%�Fu�W���K�wƮ�\t��4��U��EP����@q�4R�/-�֪Nu�Q�e����؃(e���(��gN�9yv�u֫m��iB{�yp�WWGq�+XqԘ�Lw`d݈�u]n��=/���V�M�aTkWb��f��W
�3�af�\4GES":j���GLM��eΛ�c`�t;�ˮ�g�HP$'�D�<����o�U���^^�mi����᛼��AwNK��o�$��b�=z�ͳr�<��k%�}G�����췝�w��.�|Z/=��i�ЫzQ���h�ܹ{�TIV7�-��dN�e�/�N\�z�9�T�w�5_�M;Pi�9�^fk��y`$D���͒�}2�ˣ�C� e�m��)�#��ĸ�M ��O�WE!��Ni8��+!g4�(c#�������f�\q�|�b��^s�����<��:�;��š��T����E���.��c���ATS�G������Mgnt��~U/rܚag�=�E���ټ��۩$�w^b�jMk�Y��W@�"stE�kss[�hQ�4��n�|`VY��T�L%���wTo:��]_u<��Y��U��+YyZ�u���9ʔLP�q�΍j� ���R��u׬W^�0;��Vʍ�4IFu�mQ圦�p�l��hU�cQ�3G+ ��JJdh��m������l�af�oY��ڜ՝W���֠�{�e��ݵ3��4�}V�[]I�&��p��e�)���	چ�F��O�A��}k^u�7�s�$��Q��:��Tͽ�[k�H-�U���i�`�vb� ����
����'S[�[�ޫ��YI!B&�y=�������fF@�I1ӷ�]���8�ׯ^�X�۷m���*2IQ���Tw'��8�8@�dY������c��q�q�ׯ__X�۷nۈ
���GG%�_]�(ȕ$�d$�F���o�Ǐ�\q�q�ׯ__]��۷[F��_�ݱ�o���j��^�G�A�q�q�u��;�΢��8��mtqw�bt<��rS4w9'q�WYV}]�]�G�d�_v������g'QtG]Q����Ż�y�u�Du~�dI����9��̸���:�[�wqEO7gE�qp�����9((�J;�:;����γ9�ugvSj��.��ܒ	 ������l]E*!%D2�t]�Q�v���:.~l�TR�H��HJ��{�>�p�Ū��nP���z�V>us�N�ԉ�ʮ%�:�kyN:5�s�J��TW-m�\]=~ꮽ�TͲe��37�n�P���TF���t�Ckz�BUa�r��k.�c�3�܊>:��0;�%a�qփ��]@��ٿM0�LG��VO�,�t� +�Uw�+�AS([�/��g�.A`�ǽ�8`,��?��|��׼�<���X�H��u��F�L�mlWЖ��n33�������#������@�0]�<j#;ʼ&')�@��Ħ^�Y��=�[<�}�@�P6�'�L��f���`Q����˘���D�Pj����޾u��qm��Ɯ�VG�5��0�p>F��z��ًj�1��c
n�ݾ��P e��n�\X޹.:N�!��K��%�t��楧�����3�l0�V_�V�Z�<��h#��4r�,�D��7	����j��j����;�;z��Yʞme\lz������2"�|n3M�NheW=N<�N��|��l�7�c�	}b�]zߏ��m�K�N�yKO_B���驦0�/��=$;�W9�ˇt�\�5F��:����aǃn���=�F��FҾ<ȣ:�����T �<�ξ�u��[��7����z��o0� �����sMV .-̗�=��(�v��'.���5��.�;_3��ǧ��{���N����Q��G_��z	5Tu�/<z�����{+�u��to�vZR6�����V�T	�`$ײ.iΖ�Z�Zf���E��gac*q��A�M)�t�zh�.�B
�4��s�O4�:�&gb/&/s�B�]�!���e�z��}�U$S3���j��:���,��z�(Dτ��i�=�^C{k�eF���̄S��ag�����a;�L�.˻����f]_ƟۍU�M�[a���}^�i�.�u�]"�Wt�'�i�����&'X�e74hm����يO_{(3�` W��[�d�w�h�|�����B���ݞ��	���&W>�@K���s���w.�;�{L�MM�ꪾy��ɞ{�;j��yR�Q)n�7��ϖ�FlQ�;���k�7.��ȓw�ͧ���&��6v�Cj���+���ղ�cx`ۙ$����!���`љ/ꃱq����Ip��Qj�]�Xg��]������۪wς!,ve���H��N���eh��X�1Ի����G�F���=���xxx@�='�ꞩl%�1��w��y�D���"��qbXW����W���^��g8+���aS�������v-ׂm歶^�g]�ӡ/!��Q�
�O7��-��e1r7���Xq�ֲgq1������m�����a��\��T)�R��_D�9�69>�H��LX�k4�y����D�2-[�4�/��
�E�>�n6�Z��pf�<ory�/�w��es`8*5��E� ���)5ަ�ٲ槦p6g�L'�9��ot{�xO�9Ʃ�	�3�n9������$�V7���y۔��>
�l��h���/,ܱ�n~M�Z*���r-P�h��+��u���m�@nЪ�w���2��$��8Vss'^;y���e��wf����|�7,�܇΅j�[a9Еq���>m�R�wus�__
��ޭ5ws��&��?�70�un��3W}������7���n̊2;��,�{��a�gWA�A{��#*�Vrз-�n_n
��r���%�$=s����=ƻ~ŉ�/�GU}��3*E�\OY*�)�,�b���#�k��r���ʾ��c4����L�T]�c���7�;@���y�o0� \X�'��dw}�:I'���3�g��pg�"m�'�TD�D̓=��|4Εe 
��In���^^Q=� ��ٖ=�����;�!�ú��zwn�ʭ�)����&Wwy.�������sv���d[�g�Yw{p{Bc�;��F��1��t�#:M�Pe���lkxw��J	�c�7�M���";ҹ��+�U��7�WMyb���6�d��9����6j�w��t6=��s��t�}Y:��?N�.��5덎�ʌ�=���RTz�o�� d�^y��G_���Vk�SȁW�!����L�Ŋ��&7��x��z@����u�y�CI��2�}�a�q�-�)C�#Pۯ�w�#��"�ؓ7L]T'��Uw�2�u=v܃`�����z��^�eVx���C�2�H݊�O7��G�u>��|���,	9z�ҫ���y=t�*�����k*��d�ά\*��j�5�_>��9��F<��A�_�(8ͧ֋�U��玕L��]f�>�-�f�2���&��7�
wj��]���t�
���8���i=��^
�Q7����c�H߳����{�s	$������MUe����7���FҠ����^�(}�̮�6��3r��h%U*�m^��� ����r�Cztvi���H.��EE�=J�
�{x�򋴷GM^�ێ!!�Hʨ[3�w i��4΁t��G�y8^�,�+w6:fX\Dh��D5x�y�L�$RH��ۍ�u#y�}q�@�˅��[=��D>ia�_`�em(ּ�'����5��s�q7<��f�L�=�rZ�F}�(l�A��������G�k�me����M�fE�ќw�R0O�H�Du�tn�6�D�E�V-�8�c��[�5v�H�՟�SE�m������r{~��T��w�g^��
¨����	��@�ffTc}�9�/$���M�~0$<����'�x�fk��+P���yEf1b64��6�v���\\�Ut�r[0���4[���i��OUu�d6+u«�:5��v�2Z8˅Fh����w-��
Njf��k�}n�50Suľ�~<+������n��7xe�O$��1�H�y|���=�{~{�}����q�3~�;{r�c|�����q���vo��G�u��TN���em�\NH'�1����mhv�C
�3�]�gwwgq�@#�y�m�F@�n:���w���x�g~%��n�i��w���0�a E�<#/4��T�_r����s?T=3X}�����~K�1�����L�e��M?�EC��v�|c���M;�X������,q�p�yf}���:�	
��U^���3et�W�LPcD�v�vi#��n�t��d��3H;q�s��Nz�4�f��sW��
��I7]��pG>q2�8�� ��רt��[�v�u��E��U���N�0������D8��|��{�J$�s��w��P[m�u]�s� ��)��s�}��N�Z�� `��Y��i��̂��i*�J��0CL]�d�~t��p`~N��;L��m���T9n$F�d��W��1_wd<�x�3
�̗G���`趸�h��@z�wy�ЭM�˛�ۜ���H�/��m��%B�s��Z��H,���.�/�g�Z��|i-�/{ߪ��P����w�x�4��)��"D�):,���o:wC�0ky+Ӡd���8;�G�'Q�^�U�Ȅ�vI	GF\�u��B�rA���q۱�b�m=�D�~�~=ݵ}ڀn]+x=]�Ɗ��[p�tvn���A��m���l���K����*K�|w�HP�q�u73�/_k��5M���5����}"�nJ���o���,�@��l�"�,�N�٭�k;.w�E�DC�԰�~q��s��z�.=ԯ�S���P��N�a��т:�tѺ=�૙�XqN:�Oj���]A�Vw�q���QT��Z%<-�ojB�5�Ak��/�@*=B��G���
�DM����ͧ��ۭ��G`����C^0�#��=������{͡PR�eI�ݟ���f�٥w\�HC��s{�}憐���h~�k�!90l��-ٓϔ�W��ݕ��]���@k׳T.�3�����Z���q��y���#߮e����z��uw���tݎ���7zo=�X�_\[ oѳ�:�l��{�@9Gn�m\���F�,�3�L�ǉ}��jj����z��vj�.�ö��u�c�R+N������rbKv�30�L���YNμ�o7��� ���|NMW�P�/�<�o��G	�i�oY�r�X�ΜT�%�GQ��&������E���5]�*Y
R8]�j�0�/Q��[�u��5��u@
�j��.P�|�Gg:]�/�+���E�ǽs��T�?�VJ�W[(��?�^ә	��zBѼ	���M�պ�7O���'I� .; �S�K��G�Z��A��;�������ΟS{
¬��t��w��X�Ӡ�Z��lE�wϧ�X
�!j�u=�6ۓ�u-V�r����Osv��
�Q,c,κ�/!ys�8�=�n��]�A�ɴV����v���M�������
�[���P����JA]��,�ʐb`\��wsQѼl�{^#0��ǆ}�<� �J��N��g�g�����ag�\�}.�M�8�;�^B�2���{օ%|R�p��0��Zs7:\��3�xOz];ev-���cϘѕ<���ן=HH!R�'��(���"z1�e����2�V��![�n7"�O�=��o��Ի�L�|��M�ӎ�(�7��A��u��_U?Q���㣊]����Ha	������@91�#5����ϓ�jB�ek팱תp��*~�v�;c=��r;���]�u���N��0�\.�ﺳ�Ӧ4��n6�H�F�ů�A��݂L��[��7Mtp,���%���;��	�����*z���U<�xzG"#�u�$��ǅ�B���)�'x��e�4!X`*�~x��&r׈T �SV����ɕJ��r'��P��#i�}#o��$+�z��}�V�RV����/a��R��ך8���<��@�U�MI��R(g��:� ڡ6�E9�z��*�^�K�x��FS���y��]i��y}V
�b=YOV'k�=|����IJ�w����R�R����}��z�ϲ�Wc�҂�
oc�����{�{0�N#"��a#m���qLO-���=A��gc�5ۅ�v�.Ӯ��3�ax����UYrs��TՖ��6�̀�N6C�yF9c=oTN�Ǚ`��y�	�V�w��8�S���Ҷ*��[}�;�J�
�w�̽;��]��R��$Hx����	��y����y��`��|r�Q㇘�Z�n��u	��N�V��-���<�<��U;F��p����Ǔ�@H+���[�E��� �+�gժgmlZs33gAy~�}��ˍ��ϫw�չ�9����3^͎�%P�J�0��2��ݺר�<_nq�7�f�� �{'i��k�;���E�l�Ovҟ"��{M����#f0�;�w�t�3����:ۣ�ޕVZU�TZ�D^�sk�I1w�xn�L���R9֕�G<-�rI�8`sHs9t-i����-��n��S��ث����������^���l[�i�9���;ή�f|�k����-���-�t3�����摠��2�i!�����oZ_;����~�-����ǩ�+�{�H4\5���<3�:�G'��m<��M;	�ƀ ��&��m�;H��ۭ�]�ϣ�?���[_֩�T U��UD����U �D @��ae�A��vr��207BFA�,��"�F
1 d`���d(�`)����`��,B B�a*�FF
�����`A�,�b#�$ddb�"db��$B��A��$B �F(a�D"��$B(db!b��$B
 E(D ���B
 D"!��B*�D"�`���BTD)�D"	��B �D"!�$Q�$B(D 	��B �(D"!��B(F �D 	�$B ��D"!��B
ED ��$B"�D"!��B
�D"�b!��B"�D 	��B*�D ���9��)�!�"@�@!�"P�E� "�D# ��QLlB(Q�" � B �A� �R!J B �A� �� B* A�"��B*�]�!` 
�A�"��B �A � ���B�U(Q"��B �A (A� d(�A( (��wb�
�A��$���$B��b!��B*@��D 	��B �a�FFF*�b	�$bA��B �v�pb)��d�FA��B 1*D"A��B*��(ЋF
��(����	A�b����l�F��n�<�G'��D	UH�F1͠9���V�����q���?tW����a��0�R�g������J������G۞���( ���������PEvu�*��� ����0�@b�O�/����C�?c�(���:<?pOȇ�o
H��<���?��0�;�+��?�?0���?�~!H
*�T"�BD"A $D �D ���P�1@�)�P"," �0P�P"$U�@��@��B1P�B,����.�t먺���EEQ�F@UA	A�Q �U�i@�%Q�uRU�W��IWU
 " H� ��"	 F�X�@�$ H�B"�� �("!"E�(E��X�@ �"@�E 	�R"B � DAD ��$E��T���$�$�E@H�n��!(?��l�S�UQ@P E$��p�������~��>W� �?_�V�����=�������tO��H~ o�P������aPW�L��O��/�N�W�"�
���ȃ��w�:h��""��������*�
���A;�����W�i��|"l�۠�4�@Y�?y�P���h� ����O��v~�}~a���4�� �?�����J��?p~��C���� ���<��l$O�u����	A��4����u�>'z<�� v��1���)C�����^/���W��"�ä��,4���-����??f���!�'��PVI��jԬAݖ` ��������<J*T$%�!*�*PP�(��%EH�*��)"��!T*���QQ**�($�*$�(�mJ��Fڨ�BB�	TR�*(���!+� I)EJ�E*AH��D��UT ���B��ʁT�Bk%JP��*B"����(A�J�AT *�TURI%IJ������%J�RR�PIR�jT�*�R�*"���}`�"���   c�Z�l��6ؕ�i���n�Auۭ�E�,i6�έ���R��;���\k:uJ뮩���WWn�Th�ٹ����Ym���-�9V�U��������P�J��>  l>��B�
4/[��CСF�P����"�B���\���چ�R�m)N��mC&���m�5�U��7m�۴ӛf�gZ٩�]�ĭV�n��]J�,�.��N �RDAJV��  y�%�R��tW;������{�N�-Z(���n�vܗm��R��D�[7[.��F�s��Ҷɨ��V�T\�ʺ��v�%[��R�B����$QO�  ��ow����b룕]r۶���)��&��Z�T�����\+V�m�6UiU٪�:��h���d�5V�u���IH��c�ĩ$��E�  f�|S���nΤ�p;h�5��4��:���:����r������Q��V�k�Ҋ굖9�۬uEc�����EHJ����   =�6�4F�{a��lH�ݺ���F�v��b��e�ȥWQѐZ�WQV�Ү���N�m�SU5���@�Q@�8$P�J��d
�
��   {䤥B���
��T��-ҐPQgSq*��hV��*�IT�R���s��J�k�B�uwD�*q��*�������QJ��@TJ�x   Y�U(��q�@��!*����T]��@��MԸuJR	q��)B�B�@J�F�A
\�ܢ��UࢂP�REIւ�JC�   ��T� C�N䄠��{K���c����R��U�$P�3h� ��N�s�t��,��:�P0��Q*m�Ύ�:�FtTR�!J*"U)
o�  7�6�B{�s�R���B����P��]�nQ �E�.:)IJ[�7A)E�7ԢMʳ�E"����U^ E? �%J�A� �{FRUA� U?��h�TyA��� ���R�   S�i=J���di�M�R"l���  ���=����X(���Ե,�6֪��+Em��_K:+A&ݕK�k�������߿�w����lco�� �����������lcg�l|�=��{~0E��kyWl+ګ�Z�`��,��BL��۹񧦝�F��z$m��j���Ӓ���[�
�;X����1���p�F�l�w��s$`�,�A�,�Xx3�Sؒh�(�Hd�f��~6��2�c�DS]K��w��0�$2�� U�&�X�%[)<�A�eM��6�Ji7f}ѭ�/1&r�cyX��CY1ûdV���
�Z`l��kB���4&Фq��ˠ�tdۭX���H�h�9xZ2*CZ�)�����һѡ;%��M��q��ډ���,��P&�nͭ��6�&<��ݖ�݇V�D��+�0Z�v�2��Ȭ�P(c�P�4C^������C��wD����.��6T8e�-F�j�!�H��1�W���ш�0���oY8�%��v�)!��:Y+cIc�76|`s"W���h�MMͻ�$������4X5{r�#^|��ƬZ��81Zf�QǗ�%���T���O)â�U����Z��Mî�^ʽ��U��C4�0E��t�oL"K���*`l� ���2�e�[J�����Z���r�ܔ&^�g�� `�N,tX�9��V/��U��+��G+
Ř������+jV�Ҡ����h̡-��T�n����m�f�#��	�f��f�Qޓ��W�!��nZ��n�m<��S8D֡��$#!��Fp2��xh�d}g+v��=���pn�A4�]8^ʘŲ���	�a��J5F,q���R��S�K�x��C`8 t1�&m�պG�߭ޘ��V��=�R�SMf�$��xZT0!GtVbb�Gt�T��Y�%�z�;�L��e]dx���?R���p�R�`.�֒[��f�7W��X���V�l�2�]3��*�8 ���(aj��ɵ�TA��ˬ��&�wfk��fF��aրI��\��0�/v�gajI��v��.�A�2=/m<�!8����0fV^COc����%�Cv�YF�m�J}��(���ъE9��N�Z5[�bST�j����!����<WJ�`Rٮ=����*�,�ŵBj����{��q+������;���lPV� 4D�Nn7�F�,���v��v�@�S�XqF�jGE&�{�16����[2I�V�&� ���;NȒ�H��RM}���V�փ.�"�ו"Q�-�v��d![�Y��v��ԨƋ�$ fL���/ oH�+0��O)i	�?F�����R��x	)mXub�o5R�8��
9 M7����wX�q��a���&��N������6�3�R&���aU�a�/n�ĚT�2+p+�KR��&�N�b�j�,4-�-�g*&����C���fE�Z%�Vʎ�әH-������S!2�l���kA3 h��r)i���8uP׮�G Cr���J���GMϤ�@:�0�ѽX�v��BO���6�v�
ݴ�2^��
ԉV�RJ��e,�AH�rcV]3��UeZ�,�Ă��ZJ�b9*-6M�X46�/U��{j���Q��f�:��w.�B�B�Mm�t%�E�W��(�AnP��'6�#m�z��K#b���2Ri��ļ��hych��i��pv2+t�+�G^���Rݫ�X&	������e��X�twl_+6�˂��E�1J#�֍���ݕkf�F��
@0d��	���y/
��@*ȭ:�w�aA�a��2zNl�r�Z�Z�)�2IV����ܽ$�V�Sef�5�m`�-F��բh���k�ң7O0V�:��Nh��x�	��x)�ۿ�,;��e�⧂��ڽ�){b���3j���֥�`ևX�3i�LQ�n�JYX@)��$˶�v�,ֽ�C�i¯hU����Tv�ٵ�~ʬ���Ӵ��e{f��Xƃ����a��e�U�n��H}-8*�<&UgP#:�1� ��YkB4������⎫ѴKǸi4ӫ�t�[��zq����ni���W[w'�(�&�M����5Y�wB��^!0��1-�ZZ����`-;iuݵ��M�,i��	�Ћ[e*y�[̿���`Zք�K]��H	�kIٺ��8sPOŖB���GU�`�֑��ET��$��Vm��W3�������d*�Q4d�׮cvn����F�H�'��^I�En�m�T��1��cFY��#�M]���f�4ӼcAe�R-��2�D.Jsmn-�o�s-�.�x�0�x�[,�Ig5=KXwY�o��J��N�NXf����X�>y/ �/*\n�iE�w�G��U "2ŋ�e���n�k�5���ZYb��3tK��8imɪ����4��![,fD�EE{�ʔ�JE԰�כFܹ���H�����n��DS6¸9
�|&la��o)иil��D�bdoEj1�cXt b���إF��^eȣ()R&��B�v$�hLfe4ǖPբ��&���J"*��1�8��1V0�L�Dԑ��9Gt�R�c��������KѴ-B�;�܅)[e�ʀ�v)E��.�MU�f��w*LS���QM{����.����^'9,�Ƕ��P�)V�^#�RaQ�%��D�M��7H�V��y�.H�ׇ&�WE�T2�^m�Z5�ۚ�7xq �kXw��كR�5�b�m8��kj�vf�9C"���9�`��)�e�p�%��=�ۆl+\,M/-��LIU�/p����Tj3����Z�:���ɢ�0��!GQ�V�r�9�e�B嚑=��X�m���Ͳ�ҳl���G4nm�j�͘н�*6��ބ(�kaJUv$s�;�@�-��ʕ�Hʌk0č�hi��?!�����x��nѽ�+�2�BE�Y�0�xL��5WqBȦ���i�u����ǎ;�X2��-��n�Vf�[M��Rv�dq�y�/ja9zbZj+�����#�i���] �wV���.Gk
Y�v��l���X�a&3wU a���
foµ��[�΅j2v�H�P�sJ��V4�Y#T�[�bGDm-��c�����]��Q��̨۫h��\@bx��{,a���SO�#����V@M=[I�϶�V����v�]˴4Z:jJ�#�Q����#�0��&C(:6�	��$�����Fڬ���6�]�»+xY�W\�Pv�X��	�r^��lH����VFa�m-��-�I�[�h�Ƣi��Z�6C�o-c�,FN
:�}(�H�&������ȬĆ��s/w�ԭFn��4�HGA��jᴅ5v1d�Hc��$�q#��K7�)fH����D���[F^���A��P0�޻��D���r�H����{��޹t�����F�&)� \6C8�F 4�%��Ŏ�b��y�L�P�%ME�%�LT
'Xf�V\��]��z0�8ŧ�%ZPPUt��͙B�AB�QT��x���5�2S��MhIB*�M%��3@��G�ڂ���h�����F]�r�"S���>Y��+C�u)�iR�wY�3Z�50�B�)�w�SEȶ�g�"�h��S4�f�V'׶X&�	Lub� ��ܭS�o���ŵ/V�A�nG�kc37l��"5(PQf�lS'*q6F+��x]�	5O���Slj�VAM`�:�f`͹�S5�J��
DE�u�kt���a�OUQU�gA�_[�Zu=�-AL�u�ӌ�fD�'M��nJaXܱ0�:S��˺�H�Б�P0����˹��-R���:�^M���a3��â�n�+XЮ�;�%*��I+N�vb��*L� m7�+ֶ=̧s5�;@,�Խ�s&=Y.\��"&���-�G����&M�ŇiU��F�q"�r#�
Y&e�Q�V�r�S�6ˤ��`⻔4`IT2��FR6b�r/�}���ݺK@��ԙ�Ux�|���Pj�l�ą]��������P�&5{x˄��j��Ɏ��,V;���	�j;8"�m���H�I�cu\"��q�+��P�����#��.1�Pe,�D�ݟ]^���ۥ�c�O�d`b��PF�-f���6�=�p;�Ь�T�fB��(L:U^^܁���i�b�Li]�y5�+)K
�F�4��K���T��yi�fŋT��d�����q"� �¡��Ղr��(^�7��)t/[ob��-�[�'�AJ��x�fچ(�y6�K1{��ڙ�+���n��Mҡy$ܽQQ��9���� u'�[����q]��tsAgV9Q6� �r赇L��EE���U���#vxlaL8�Z��xM2Z�A �d�{-�<{L\Q��^ާ��(r��o%���Jԁ4��bJ���R)Wl��Y0aڽ����&'�1�O��-�F3��Ƃ*mݱB,��Qi�j�X\z�e+G�˖�v�2&e%[q���M�ż�jn�k2�ilU�F����/�k��2R���{v���+'V<����gZ�KB�.2�"
Ũ7PT���
��ʺ��2Q��E,�~]hXs,���i̘�۳�(=t҅h�q:����c4�����&��H������I]lWVf̣,)J�;��Mg�
�i�>6h�V#o��&,vvk ���ڭ��M�u�B!{-�p�v��w�+�Vc/i�ҳSaP˷*O��)�*��65	���hЌi��2*�f�"|FQ�*�ֵ�(����b�_n�2���5FJ2K��%m,��Qa�ق�w5ԡA�*$�c`F�!���V<�M[y�̺u�L&�W��AVQ�l"��X�t�C�G��9�<9u+p4�swN���;�5�k!�ح���{4�UK�`KQ�&�r��Z&��ע�fF�A'7Y��[�o#a�
�\TT��m�*Ō���Չ[S[�Sq�H�Y`�jRɘ�+krU�sU;"�4�wX�(�I�JQM�]���)�q�",���Nm��h�6d��#���nn�(ӄSeP��,�Z�d�麕n�Ԟ�T����+ʠ��;jj�X�*��L� cYo%�ɩ��zT� ��Qb�нb��^��MS�ʷ��Xx+VW�=Ө&��fJ��w6��I��!�!���b�r�lnX�b���BS.�Q��Q����4�K(�S\$}gN�-��T�b��V3f�!Y[t�#�ѥ��
c3KV�ÈH��{H��K�Ъ;��w{V�:U�=�]�I07"ytР1m1���4B�.�
���9 ͼlǹ{p$��ˤ*���')n�޾P���0���G 6f�
�A����1�E��*ҹS1��&�R��V�41̤2�\�5�5RfF�S1�It`a]e��=ݩ2�M��8���!�f���[�23���ȇ\c� �i��/H%��+�Z;TJ���:���De44�'1S2�VJ��ɼ�2��a:���]�+4�@e�!n�v]B�^ V��ݻ�y��Wj�vtĥ$>p��p���˛�ou��uAc;�9F�c�)v��*�5"�᭰u�4�J�4if�B�%� *���,Ӧӧ3Y��nh(:&�̵`�Z
/�����0nn�ӄM�T�,hu�M�eD��:�Sf;���0 (��Q���j�)WwC#mLԕ0��{�'"���F��KX��yGe��6�,���O7c6��V�j L�F��D���OM+�(;��hb�ˬ��5�俑�tѺ9u��b�pm�NK�u��Uz�����hm4�Ӆ3k7v,�u�j�a�UqF�:��fa8��S�^%��Y���E��%kə����r8Ћ-�n��$մ`ZY�n%J�����8�c�@�e͐�m��U�FS��Y{繙Ճs!nR�Q$kıY";���c�b�i��T��Y��fR[7�R�PN�N��h�q
��r�V�����ce!LV�6���	���V���^^Y(
rX��[Ly��-J,��.�n;�J�H�
����C̋5���Y.��&h,O$�NU�n-N�Yl�,Y5�7v�A����*�N�:��F\L�(VLC^��p^f��a6�&�"�H&VT��M���2���A�e�*֊���הhKx�˼����(��.d�s�aL.��.m�4�.n��-�h��K�q+q��Sf�ah8mJ+pmPN'j�dn�]ͻ�j�Y�[����oA8h��� J��'i�D�I�{��^ݪ�RBu�-	K,�!c�0V�wA�mR��%�g-��n�ě�7�!W��	��x�e�Q+tɰ�B�0T4����Y���=TS.��/��R�Z01m:�XޓB!��Sb�+�2�t�
C[�����VD]���ޘ�$2�	�
4&B[�H+[X�z���J�4hZ���o0�On���1����N�/q�^�����P�e�v١�,Yj2,T�oRGw��(J�R�Ȳ�^�Gj�Ɓ�f�g0�ƶ��E��Wv��1�q ���td�-�3-�n�(��������`|�p�lKu��*ۺ�����y�Z7r�B�:�ӹy�0��{0K�Ѝ��NɊ֋����@�w �wY�=Up��R��W�l���� �0����\YL�]�w�O���ܡG6@G�f�ԋ�9M2+;Qt��MfV��@�nXҭ�k�kN%�Q)D+P69q�r���hm,עjvݽ�2�2�#�Gn�4)`B�Kh�8�ހ�;���o^�R��21غyy�������H��j[3D�ne�j��A�^��r\��9KV��녜7�@��!i��,���>,4ĄǪeJB�M�
��M�����Yt�iVӘ�2�yX�uvm�z�����v��
̼1�Źf�@�@k&�݋tK)i�mӡ���"�A)���I��Ǆ!�KVM�-\�`(��Z2�̛����]:�&_w^�Ұ��'ؤ�y&>�9}�aO�Ek���5�c�拑�1�i6���_<��a��W��s�יO,o,6c+e��՞��s�ͮ����9i�+���(�ǫM�ed�����Ft��.���O�Z9��-�>d���HMw�3r5Ԩʽ�0%�;A����V;HѶ��!�{�}��p}g�u��+�/��xqQ�{-շ��R�6f�<���ި�,f��b�x�[�:�!\�u:�cú"��uv���%Ns狴Fil\j�v�=����'h�2٣x��bJ�`�K����5������ά�4Vj{��7���7h�M�T�F��{yx�21%t��)�t>;ĤD��O�0�Pp˩UY�a��A{ ��������Ɣ��yG�Gt��M�R��Xޅ^gfwg$������JN�,5�ΛɆ�<�ۍ���Z���;�A���5f�2Ԣ(�L����J�
��) ;^�=´e�nGQj5|3b9ΆT[E�"�c�/3g�o]�����gkb�"���}Z����`=q;�Ui7!J�R-d��e������޸U⧢U@����f��]��y��0E�qv	Q�	�Ŏ�X9��uՁ�e��^k�ۏ*l;��W��Pc�>�Ne�s��i��4��<�����a������1^1�Fע͝I�B�>Mr��(�V��q�xb����=��u�� k\�ѳafH��B��*<����ܘ%q���<J�a�8��V�xR�g8��Hi}E���|%��exs�YԻn0��N@1s�җ�L�2��*pk�e�;�a}�1IAS	�ؑ�rָoR��]�Y������Y�;��U�8���OP�)V_Z\��[*s��wټ���7�m��AW��̨zD$ע��Ȥ@h�Ǣ�_�Q�76��|�5���%���KU�;�pZ�+��R�S-#չ�8y�:���>���0��~"����ut�0*S%��@]^aa�óvCޏp�\�m��M�c(��y�W}W&����N�R��:�sG�2�4�6%?��:Ip��JN����ʵ=��6�d�xp�7n�$�ouc�Z����|rխ2�-��^g��}����4��A\�R%@��Y`���X����s/�&�ظ��!��`�B�ܛn��-õ�z������ޱu��W�>��*�ϪK�r�'}vL�QI��*���6���֦y�����
Y๏EY�����>Z��Ԯ�B6D)
v\z)���f��.�oX(�8�u=\��e=�޳���]���������:˧m��Ӹ��w]��<�!����-�/E��C�D���\9�^!�oo&�4Wo#I7��h9/K쭖�b�:��X�F��щ*r;��}Ɯ5zE���x�n�ȻdX(RN����0�����Q� 0�n��N֌Sz����E�x�F�Z{B��8�:�\T���ktͷt��;2u���r#���c���v��;[�A�(��]�b���,�	ց�+W7�ⵙ\6��s7�]Y��, ���5���,�Y��f�/?����Jd�Od�������,�nRޗ˨(J�@o}>�m�1M��n<Bb��P�ts)C�J���I�[�fc�2�]��R92�'���N������ ��R�Sn�n#�7���9i������j^���t���J�RJ�n���<]�&��|�������ynw��F�,���~u<:����1YD�*�s'>�k�5� �S"���X�5�u ޠ!�Cu�p�
�q�R�ԏ\:A,B�>�qʝ@���,���/�(������jy����c�Kz�Mx�N
�7�v� ��{��Gq��κ����RX�
q�@9ƞE��6�L�M$U*��L[Z�P����1�li.ei��P�[l#nn᷹���U��J7���T@��T��c�k�E�lm���BS[���cigiO�b�XVh��/o5-|�ܬ]2��H���]#{a�Im-A_v�1o&w0V�:�S�^7Wv�����Q�0R�6(��idt���,15t�+13.�����uUͦu(�MI��Y"�2��ov�,N�JE�v��9/����ٍ���L��K�9�+�F�n��R���9l���ٟt�j��$[�]���6_�\(��$��<�u�jq���	G8�`�{*gPAYP�ކ9����p���5�nT�k5��]՝�d�é����c�ٯ]�j`)���Z�v��W��/s��p�bk�,�z]�zZ�%�Z;q����Q��T�$f��ڵJ����������	�%�MQ�d�(p�a*��]w�`�0�k�����%h7�z����}V�0��˛Z.*S��syP���
ö�@�#�	��1�w��U����qa���-5
���%�^73@�����L/ںu�>6[��7MdG_\pY��#�s�S�Ǹ�ZӲ�C5,�L���Lμ�T�E���h�x��H�Q�jr���1��m�j��wIs��4�2���O�0������v+���k7z���V�����y­��qco�*�i��j�E�M(�t:aR�B�"�8��ep��:-c~�p��ܰ��խf�T�����q|��Dd�]�����B�:Ҥ�;���]���
����k <��z�O���V��U�f���
sOαfԎ#E>�ީY����^�+?I��"FӮ�m�*-��QM�QT@��A�vQJ�{*�����smn}��}��f��� c��t��HLǆ��ݭ�)��Sf;���WyP���|����髬v�I�ҭ}� ��>�}�VS׻[]h]S6��	"jT��O�9���#�X�Ϋ��'p"ub�R�TڳG��\�i��ô%
��<�\�j��n�U�:nl��i07H�˩�����X0�Vu[2�ê���j��h׬]���u����\j���U�=J)GV����+�>tN��]�%]lF���ѧ^Mn�=WuY�����m�P:rh'cs9�+��K+;V�}!��VuN����ǜ�U��;.�w�ZC�
�lLHμ�e+����L��u�}DIT&S�C�i�;KWf��|�wn���|�Ւ�p゛:��uw�͈�mQgfmm�`�_�,b����Bn�D�
tW'�$��A��g)�pU�*!
xGƹ:$Q6oM�u�gX���!��4I�Ű��Z��p(f4�Q�åQ��n�}��ә��◽�]>��Ӻ�;��<�`�D� #��ioc���9l}ς18����e���DL�i^�<�<vu�uv��UZ���jS�m�bw2����1ѩ´
\��^�OI�<i�����S]}v�ٝ�t�c粤p�urދ	���hS=c�f_R}���w}�X7� W�j�.�n�<lwaEsH����Xޗ�u	�O�򐁶�h�,[yx�b��T4�mr�imo,�˲�c���k�7����a.]7���R wT#��*��iM���Qg�m�XQ6:�����1��w
ݾ�Y�D-����p�u���F���؃�(�μ傚��=��VXv��[P��k>���{|�Ty���*�y�Ӽ�֮��R����u!�5�=����Je��n1�F|]�8�Fc_$��ӵl�p,\��N��Zut�V�ʊ�Kag/a<�:�52�ݓdv�W�3��P��,���6%O�:����r�ef�׽�������C�{��j�Z}�D\�׾3�w`��+j�2��(�o*�#��7C�]��&\`���d��	O��u§<��d��Y-Vj��i�S��8)�+��´���B�{�gr�d*ch]dx��,NQѻ	�H]wꓘ��T��Vʻv���q3�VP_=���4w'�u$�	7=�t�r�ʜ��wV�	�)`g���:�5P�k@�9�(��w���Sv":�]��e�¥1�&+�=����w�rh^qȺ�y=�]j�˱G�T�*�D=o`�h]1#u���_��Ó4#�Z�u[�oM\u��t������W(,��J@�Z�d8ڔ^曗7:���%���vt;LFT���H.�1n\��l�.������sC0�VM�~)��\*�!��'ɖeG�������\p���ބ���g$��sb�F�čL�c��R���C��e��X�XuS��wkv�73��ͦY�C�m�E�A��6e�{CQ�FYQ�*�g���B�f��H�%�,�u�Yڊ�T\����w#���4�<f�;��Xɔ����9ƛ��#ݳ�E}ה�^;�E��ά��.5��6z��o02�y�_9]�)��`�c%���Ks]�U�j�9�O�(�;����9�%���P�ըn@V r�c}��)��f���Kx��pu��+�뷹 �g�b�oA֣���ֵz�{ָ�}�B�hq\�\7Ί(���;��Z�K{ݘ,�"1�r`1�9V;w�ꁷtq�����.���}��Dt�z�Y�:����ٿ�u��"��u�����l�g�bZfq+9�������@޺k���j��� �n�_s���5|9��c�<�֬�	I�[q9�n����A��Ӏ�!23r)�l�'KC�m�11�p�gSEjw
��P���;v��)B�>�9�r���1�q���UÊ {�[�+�v�t!��#��ݐ�BeU���Q��:��B�۔��x�D*���������V���W\ߕ����� �����AZ-�\ܣ�r�,1��Vv������4L��������"4��P���,��[��3,4��6�����Vq��5�v+��L˔��s��n�5�O�u>Khm��r���歁B���V�I�2p������-�"��ʆ�Xtӻ�0��:�p�Z#��P�W#ε��ɨ͔�:.�[����,%������:7.B^"��3KK�Q<vu@����mtv�)�ղ�ͮ�Oi�ھN^c<�P�Q�Vv��iWC����"�\�Vr m�NC)���a6s���9u��&}B��.�#����kv�(�wa��f��
U��d�z\���e}v��D5��v��T}�s���W��JJ��v�.Ľ�1��̰SÄ��RZł"m7d�)$ɻ�(�e ���uةm��hk��n�pv��b^�r]��W�׵'&h��9�ԝ��7'��Q#����-
lxC�z�<�"��d��v͕,�E�SFiU��31.1�%r+l��*Sʹ�B�
��sv��j��OfKc��ĝX�`_Gk�A��Wult�Ô�#㚟ikj���'Q� e�̝����>���+���\Z�_l����W�ܖ:ԭ[8��7�Kʘ��B]#���Yuz��Wnl�.��r��F-]F9��ս.��m��y���mx��J�\nbڍ���wyrU��"�P�;kw��b��B���e9Ö��n'�2���ѻ���5we�v
@E�T6���|��G
sX����5|8���*Wn�֥�� vWX�bL�|5l[�o�V��ZNl�D�4F�Y���Νֶ�{���TNs��t�9�#s��An+o�����9
E\���8BKbu۫�� �`ޕ|�f�n��[��Ğz�!F�i��W��iV\Rl���;l�;󕖀���8�UTl@C�$$t�D|�)Hd��@��X4#n[�F�]cE�������b!�W��Rγ�^���p���Kk/1Z����:����Ռqʍf���IՕ����R�X؂̸9��7����'�)���W��5��V^҆�S����͇�.��ΰX۔�[�*⭊����+d�ٛ���=�W�a�y1�F�.���O�&��f�-�7N������;��UC�
iJ��Z����K���
��
���oNK�	��lޖ����x�	ݦ6����]^%%WӐ�Jt�|���.j9HR��{p[E,:��(>���ﰵ���sq
�PЄV��V���|tڵ���u9��^�t�GB#�@or�&�u|�wuE�s3ym^�㎺�q���Mbr���w*/�N�V;��`�m���<�\�}8�E>���JwW~�yyn
�;W�@5�Z���o�h�^\qOI�%�^U��!h��o���BE�1�5lu�{�E��źD�������k���S6dN�?�V��#�v�v(�2P���V����[u�fH��j�:����-0�癳`W��f�kIU5�z�Z��o>��#�-�Y�7q�t2ZJ��xyj���f���}�q����|.�{�Zs�k�=V[k��
��P:�߮�V��q+�͠��-�dUrV#��g�yy����RkK���ޗ|�{��]	�5k���#D����v�d���]�4�%-���LPIJ�[����x4[�E�W����i��&�{�dـ��Kd��;�n���/�s�FҾ��$2�᮳z�ǜɷR�T�8$���M��g�n]'�>�J�8�]�/U��J��.�EZ��۽����X��#&�o���1[�v��T��R.ꝥ�&���,r�ص�, K{s���������:�㋼�In�|_���Nu����69�P����*[ڽ1��w5-WA�"`��3��Hy\�z١�%��N�\Ĉrs�M5��9;5.ޮ��-��&�ur����V�n�á�+�Qھ�k ����u��W^)�\�N
�� ʁ���W�$��vz���w	B�r��.tfq��s��\���*��13�ob���)�;�c���w	�ۋ���T[�*��u�J�Z��-_V�g{i��tP��ws�)D��d��� �3�;�.�V�������` ��cc�y��׮����Q^z���t�9� ��S]��k���D�)�m����(�S/&n�a�n�w-���vv�7��.P���3f�Wۘ���kO�|�<<h2�:�ͫ�pF �Z`�����/���6�H�C���R�`77����X�[�ʣ�R�	o�&��wq��@$�e��Q.��~Ǩ�|�؅�P���4��m�6�t��r����m3pRޕ�c�JV.�6�
jF�e��7y�!U��jȫ/6m:w�)<��/ZX���ɔ �
w���Q�iI�U�g��8Gӑ���Gai�-MjTR�yGv:0��\�/�^GYQ������Ӟ1z �c��3T3$�Z;kzl.ӈ�h�|Ͳ��	?b͗��w��%��Z*������`���e7X����ؚ�A\0��S��6���ʏ�N���q�gb��x�Ek3���:�N1����0aA�%�A����ԳKc���ő�#��{�$��uu���>�
-�G�r��}��;T뢏F�/����8&�$cc:e��}էq�T���f�^��4���7��a0�6�T4�8��Q� �e��׃u�vZe�ç]��u�����*!x �,]3��C�g	YF�U�����^ \;[,ێ��EIkʑ!cJ�ݲ2)P�(C3���a�в�:�:quK��rY-`u�h�N�T9ܭ۷ʣ�RUV��i]4��E�s*�VR�����C���H[��qv()�.v4F���ԟ.:�8](�.�t�(VbwW3h@(m�e�Q˖[3��ި�Y��J���u���X˭��;�I4.v?�čY��U���D,�sij���ʂ�6���C�~+ �^�z�mvV�x.0��u�I��:M��jH*Y)i�7o��t�cw}���FNG��`�6K���/�k���g<�]A#\�јA��\�&v�7k(@J&�^��`X�B�=����>\�p����F����N�l7��x	�VV���Ҹ0'����r�C�0YJ�Ac B��#�����X��ʶ�M���������N�^δp���HV�@|r���U������{�2�_S/�c��ٖ76��H�\��.���N���'U�w�T���k�>�Xf�˗�����t_s�8�
��Ѿ����@�ml�x�-����{���BR쬖�̘zRf��;���1�d�Gr����h����&��g����������۳�0RT��I�T�7��Z�C�	/';u�t*��"�P�+�PYX��V���G�oP!b��2�ɗ9�rJ��[g�^ͮè!]L�wl�Μ����o����%�N����L$��C�e�R�Ju�8_H8�:�;7%:��g�h8��x�£��p�U������:�ޱk��Ĥ���x���f�z;O:V��.Wn���38`S�j4��3�G��f�d����"�r�Oy�z�����ed	f����S��/�EwZ�]�[Xz�=&�3��p�Ϙ:1�n=$��c%��΀VG��CO�=����{XX�7
��M���t}#�`gk�WWWAU���
|�=�҂8�U���*��҆\N�t��Imh�;ꁇǯU�v6�ge�T|�0 :E���.p���ǔ!�ʎ3Ƹ�Xr���F,BP��.9m *��𥼕�DQ��[���y��+ܔ�'��lŋm>aw_�qj�+�k+;+4����h�Q��FR��hq�f:K;���P������v����ڝȮ*��|u�;����YO�+d����μ���pi���)�"u˖�m�8��L�}Jz*h���Lc[��<3S��Ƹ+�a�|��0Q�L�R��IYx6�vS��R��Y]K���%�V%�-;k5���;d��p�9 ��^6����Ͷ��쿛"���n�^Ȇ�B�]AX5'L�(g��&N��b�+m>�2s}ys���˃���Ғ�=�[N�T5����VD(f�)�.d��`| �`bP���w_Hl�*����U݊cL^4#�cȍ�W��V�n�zf�h��e��ʷ7����@��T�Ioww;C�e[Ive�Qy��G5�����c��k(�v�I��H=c��2�m+k0�ÍЮJ�!G{����sr]�m�Q�����5�����r�;2���S@��P��t�d�{��.��nޛ�pdg��&��וH���%7E���J��`M}j���gi���+����v���"Lm:,c�Wθ�,��L�}�Z�IZy�7�D���^b��XI�<�}�[�m�S�f��Ih%�G��oc��ki��?tTb���//n����K=���LT6�<���[t���1M����K�e���l�6�Z1�Iq�� �7Gc�frA�U��	}�����B	���,^N�[5i΀�X��W��b�&j��I�9@yM���qd�Q$��Z[��m�s�D�9��8�,�㜏v�]���8Ga�7M���_	"C������/��9anYU��G�UR�P�X+��j#0f��^��,�kzL�Z��u��(�1�	�U.A�����X+��$n��p�� ��{��*,���2t|��ւ�&I�eǋ�:��cM.���5A��z�Zl4�4�-9oV#��h�l���u�+�Ŵ�罴�)��������2	� ݲ�v�Tr����pFu�n���Y�WL�f��6i] 1ժ(�� �]]>���@��J��u�t[;�.�ʎۖ�20���-�Z�F8�o-���Y�~#6�Z2��q�j��*)*m�����0fI�lj�Η2�X�\�2*�W���;���XGM�ڜ�q��(2)b���UP�j8�@�nSrڼ]��J-��{���Zz�jQ�ϠX�sv�s�I4�ݽ��B�]���Y���_m����x2�9��d�-�:Mm��n�ھ�52�M����مv͑-���IY��\��`�~Ͷ�Y�`�/2��F��j�b;��QV�b��b�Z�&��\y3�L�k�7ed�:l<����nhL��E�l{hi0MS�f�lw��K#r,I,�w�v�&h�&	�v��;r�Ƹ˓�Ƌ4�¢��f_e;���R�mv��1�kp1�@��'Q��59V��[i`u7�&��� w��<��v��#I�Ry�xa��Bvj�a�	d�Rͬ:nv����"���쾙�y[���AYs��"5�����%]�^�ː�������M3F�;��󃳧���ԟmEX[���2�[W-�c�΅��P�d=��M�rHa!�'E����G�r�$�K�����z��B	�̗�ۭ�%G[^��N3O�u�׏�����-��v�|�K��(0oJ���1�}u o�MG���G!��xnX��e�,;�&9���n��N�m����)1��1�m��R�i��u���ب���+7c#�5W�Z;ObUq�T��UٵvΣR�v��^m#J�b�������=��#5n�w@Ezh�S�?��5��6c���3�|����>сZS-q'a�j����X<�gg,*o[��}�����E���̫�d��9]ˆ_Sb�glX2y�9��9��uD(\:�������q��cѣ1�\U��݁x,"ͽ�oQ�/���F�ӽ˃�%qRmY�X�.�*�Ӕm�
K�y�7����O�m�)�B
��j��V��@��T�W�h�̵@f��31��zXs�Z�������7�P8B��3D����K�k��"<s2^u�1�A����b�i�켧�+]u��5􃢡fm�H#���t�\�g(���m�<�4���9֩���%�M���*�[�ŖVvkךX;��L�'�S�r��뮄l������Id`�Sh@�0��'1C�|�r�k@��]�J�r �"I�W��T����Q<Fk�
�%�ب�╚`���. ��W���z�y�sPP!����)ԫ���S2&2�H�a'ˇ�L=z�{آ�nG���|吳"82�1Ku�Y����E�*^�%u՟K���ŰS�c����v�5��#�w����nΗ��0؎�G�������@ޫ�w·N4[�4fei��bN��.�Y)���u�)�ul�V�m]�q;w�N7��Xyb�U}���Q����F:1`�,���Ԁv�P��ypb����Cn��f�l��p�0�U�2 �줴�Hs���B�4�	ф�2�pU�=�
��wqY�g�0m}-�ݚ�At34�CB�r�C�h<��.sn�[�V�����>,���϶ȘxPG��`=ZN]Ǚ��	���Ү��9 u��bT��,��4Vh�zt:�͠r;�,�ti�n�Ƕ!�Ϧf����∕pf�����Fݧb6�:*A�^���F0+]�f�ÛHz�<B�22������ëz(Pա�*�}���\�p�w�%�1�F�,Й�6"�����61t�ٲ��'-i�i��V��;�c*�uIO�vTU����8����M�cΰ!�#��h`1�����֎<�����1k��Ma(E�6�����y�]:�z�4+w:ȗw���WX�+�RD��bv��dc�����kr�A�W���������+.X��pR1�e)���u��Gpu�gZ"ˮ	���TI�6��ycpb�w����=&b���s9(�d8�Mo.�Z�\�&[�����P-�/�h�RY���[��n�FZ۩���,�<�5YP!���k0l����
�&���$�<3��K���'��:�����j=Ě\;L-�YN�[)�M�3W��:^G1j��I�-����Z|���.�|.�6����M°���w�G��`oT��8�(W���uy�fr�Q�K�fU�������Z)���%�9�u҆X��A����@�� jb�5Յ:z1ˎ�=23��kjl�Ƌ#\"���s/��;��P����-�F���m��Y`�ro���"MX|y�ێ����ӝM����܄�dU�Z�Tt�f �7��հ���a����}��٧�gv�]���S5����;z����%_a�rB(�����U���f0���!f�lV��QJ)��ι[l�
Y}�ᝓ:q�a�7i:=�g;�/57��+(	ooE>��NxSF�y+:7�:*�e0C9���ˁYYz���gĆ���WV�l΂9�c�퓎��]�̣���-8�O�j|�Q0�:-�}���a�3;�f�Μ��;�ʚC1؏�����^m5ƺ������7(�"wL�89G���+K��x�9A�����#k ީKV��V����Q� �WĖ�^��V2�%��$�5C0��#�7�EIX��a�b-K4q�v�b�$r�ito�Nk�g(C�d��94�W�aM=�5k䢽�<�1����\����v4*��x�ysǢ�tL�/6*Y��c��&;�Om�3���T���N�SI�����%��IT� PK.++iWWP�t�'RtH���LWV�|Y����[m�)ki̩w�"����<��ͫCW5�o$��`�BPC6JM��Ai���5�.2�t���^XDlZv�V ��Y�h�i���Ж��,�2��ݒ}��w;�;g^v�`Z���*�n.������AR^l�c'ΰѮN�KOz���X�29�Y�Ś�|w��3*����x7���0��٫�o|�+Õ{�)��\t��jmٓk��^��]�����lp�ٓ��+Zw}r�6�Wj��]�DA�♝X�a;�˭0������mJ����]�$�5݁Hyr2�u��,"sn�d+��o�yw]�d�D�Nw�l�'U9�� �v^-30�J9��|Y�S0�:ژ0!-����5�j�
d�Մ�$T��fS���VsW7n�8�%;��Hg[��.��3i��\�K�\6!��h��:y�mr��욶�B��܊�p��ofu�!b1mJ��3Isw�n5�����/P�
���[�7�����j���,LU����"-p �)E�>gH��y�;s���k��m!�����T���w�59�s�uŹ})T����u���IE&� ��K������~�n��"A�����1�vnPw�:4��˭����cш��\��'P���59���=�uIŤSR�k_Z�Fe�9�&��p���(y��1)n\=�#˓)�`U�؆�#h�$�Y�95YV/M�̉���Aȡ�vȸ��v��.�Si,8w���؀Ci�ևm$%>�Gk�� {��H8�V!F��9gtv��AtX;K�[�8X�q�4�9zhffs�	�끕ө��ΊȈY+6`=H
���AR�X^sFк}�g
�6����Q��et�º�B��9q�AVЕ�+b��S�>}ݏ���q�T3��i���-i��aj�@N���O܎����CkDaPb�;@;��ʼ��Ӓ�ޫ�X ��Nk��Ի7Gq�hƞ廆u6P�VC+)`TB�ȕ^<��%�o.��s��g�H�XԻ�S�h]��=��O/�]�4����_Xέ��9�Q�Y-�$!�;�&Ő���n��`��I��������:#ޣ]C�(��B����JN�N��Pn*�v�� Q���v8��x��t�ƇI��N��:������ ��e^v6�c�v�se���k5�m���M':�7f�m;msCG{�\��}oA�����3���[7�������2+J��M#]Kζ��
$���۴)l�ȷ��l��+ d�fh��DDk\0����7CA�Վ��h��+7�x�@���� �ϕ�K��S�nw's[W��R��@"���W�'ՙ.*����x���K�ͫ!���܍s}��i���iSO)���5fZ�u�@���|>��}�!o7�c|v�ae�Y��2������yƝ%A�-{��=y�ػ�M���>�h�E���ou[��vs��b7n�ps��9��\�dGh�ٷ	���iZ��y�S�}N�^RJ��P�5KȌ�0O�X�eA���qO�$?��y��뫖�J����=��Oll�ͩ�j��y�n�vDa�����쮪�
ǜ��gf2y�)d������Jf��և`��\Ngm�+v�u5l�r(�ھ�\�\6�lйQ���dfY;W�]�Ղ�
��n
:���-��_-!�u݊*h岷��Z\����fR���Ȣ���by)݀ؽWY�k�vi�P]�XZx���7��MBsV�n��:��� T���l�'/�?q��z;o�9T#}���v` �#%�V�5qH�����2�A��_�|��왫����~�e<KhSW6Y�P����/#�e�-E]��w��3�o�ٽ�P�_U�%���Ŋ��:�d�K���7x�K	���{�n'�+s�*nF�;�Hڻ��gk\���S�qvU�g�jaG�n�4-�<Fton�8����]Y)���s�wf� J�梲��.�\Vk]�)�H[l1���Ζ��'�%���.we+7E\����
�X�޵�](6,��\���*�2�g+W*�l��2��^��jӝ���(6���9VuDwu�W��d��f�G���I �ؐH�u�#�Q(�QY�.dG��#9��!9U�*�UD
��E\9�I2e�J�*�;(�GaEED��"�
�A����aEAª,������PU�r5*#�W
e�S�&�"��\�\�4��l�\Hң��8\.Q]�T\�#��Tr���HT.aG2 �
��À�*���Z%D�r��DU�*���N�W(./"Q�Ǚv�\�e�QAr9LԈ8��r畇"��СR���I�M8�I9��
�s�EE.�XQv�Dr""�*�Tq�U�HH* �*��hp��UTr�q�dȪ�FI�;"�����(��PC��
���DU�mΏ�o��&s��\�Z啛��7�գS��ݤ2m��l����:u��d��GWm��2�}�-���)3����2u�Ι���/�F��z�f��C�[7L�O�u��::�ĆÃ�2����q<�z��w�d�N"���2��:<DO׈y�@��/�Jz�
������PWg`[�ۜ�={9.t���p×HuN��ʳ�
��l\��1iHk´#���.p\���F.����T�
����Wf��qU���Jai���_؝1+w�@�ϫ<�5l׆�j�'��g�������я�G]�WE^�]UX>��u���:�կ���8n���إ�d�����_��37�g�Ӊُ��>}��A_��Bםg�U^����,��%6V�[
^���W1s��'/�W���K�|���l� &#uV�5�LB�=��,ξl�{8�D ���?���qi'K��g�!��P4M�c|�嶜/yc��ǂ·=x��U�~��w���2���ϙ�_3����{]tio�8<<��~��5<����Q�h���j�㚤2�r<~C�ڸb��2���܈!U�!�A�VR�W�T���!��q���Gz���avNd����M��zM���]��}i���P�2‮ٯ�V�f�v&���R� �t/�GY��/n�U�:u*���j`Vm��c{�v���Eq�zpv$���]��
��Oc�M�;��ͦ%��k�+׫s�uuX�z�U�:�~��b�k��>jO�ã����1=S,�"��Ɯ�������"�n������ #k{��<)T�<J]�>��x�˪���2����ʠ�/���1a��i~�����q/G��tL`j���}��
��ՠ�γ	���oUN��a+!����.�j�dP �����D�(���*��9��_xM�#�&`[����J1�4Vnd����燞O�/��xK��*���,������{N3��﬚zn �M\��53�>��u+\�L�M��!�������8<�]�)��\���g��޵mJC5�aN����ރv�B߮u�רjN��,s�&�n\��t=�F4|�fW3����|��I���^��gk��*#ai�5���ݦ ᚽ����0T��;��יUd^����b��é^L���=P����#]����x<���2������4 �4��uoE���gw���d�Q8~�����v�$C+�E��jG�I�&�Ȉ�ֶ0N$6 i���5~g堭������钔�瞛�	�:j����$�~��o�0/SG���=Bn�᩶E]�{M4�݊%�[�t�&i��-��͕���&��mq껖�gN��H7X�]9!ʋ<mfٖ�ʰ��HtU�_u�u��Y��L�r�}�D��s���y�%p�l�g=^��t~�=�~^z�Q��x��+��u���1��i��6d>�w��+���nKk
�7D��d?!킙���W�v΋������ѥ�TN4#wc�U�~LN
LC��6�P�(]�岲���p�3M'(D�q[$�3�85�՗ϔ�������WJ���uS��"�Ѕ�叶��3>,}M�����P茏|�2Z��nҰܫt���d��QX��ү�KF��b�
,4��J>�1�᧓_y]J�:SM�p�m�\lnL鏼��c�r.�_Xt�ޔ�.�Z8��6��c7iЕ�9B�7`(��7n`������'U.m BG��P+��L�A��׽_J ������k�5FXS��������`Ͻ�D6S��H��h��wtj焺���z��q4�UĔ՞��z���idèom��f4C�D�&�]�~,E��$�ڴ��4��s��\��ص���V��٧V{��R�塣�vYȇ3���Bt0�P�S��O���hm�,���ٽ�ML�T�)*D�ø��@��ʖF���Q^+ 2�X���͙���~T�{�wR��g�ǝ���I�q_Q��g���Z"�|��/~��^�»w�n��H�D:֓Hfvj��o;r4+����Wt��up�;��{�Y��,Y�f�����;��=?���/Yr�p�{�������
f��`#?`̼F2��ӻ�L����5s���g*C��C��;F@��"���r��TiC|���c
�Sj���b�p	�b�^��b���]/�0*����Z���E+�z��K^��Ӽ׍��#��RL�;� ��st!�e������1"�H�!�F�Ø��? �`�����_3�l�������:��@�,yn��\b�3P�k���8O��?v#,��ȆKe$���l�G_�ח&;��e��=�­.��Ϛ��;����yXZ`�+t]�u=o%��7��)"����=LS^A��n<U��:��E9l�s��B��f{��i���L2����b�g�P����(�~�^� +�ZCFϰ�x1h�c1���Y;"7�}Z�Kx_z	/�TX7�ǆ�t�({MsewM/�t"?)��������B�[hT�w�y�@/��7>u�����rR S�t	�t}0H�:S&�Toۅ=�����D�9�$=��te'�#�=��W �����sQ����[���w+���7bSzc�,T��ss�3�*V+p�f���rM��A��m���!=�O�\x9섎^��{�|4�K�:J�+ވ���$B�˦!��>ɅT��|�5���Pxn5�0���Ek�_����V��F�t�]� ��.��ݚ��ly\]��{L�W�ƝպF�4��ݐ�!��%Υ�\��:�����tr��b��iN��{&��_���?*��j�.��m��Nm�Sۭ��� ���#J*59�}��>
:py�a�g���A�9�%>%0偯��3��=����o�`Y�� ������Y�I�:v:.׌�f�-?��p�W���뻜d>�4��-���NH:�%j�������:<D^��8���P.j6�V�4�=���+Q�ѓt�ڰ\X�s����n�F=n�NG����(��yȉ<��+B���`��+ݹX�Br�<��*zX:4�C�5���̥�18�2�ꘔ|�s%�Leb�ۑ1�ybo��^�hʗ~Sl���������=�C!UV�'Zϙ�}��^5�B��ֱ�PE�!�f�׾D�ܠ7|Ux!W��Ӊُ�����/��h#e�pK��;����2�pU�0�^�����PٵK-�}�)����r�U�N����H@�*锱����N�^E`�w�^��X���¬���ݍ���:���ض�|��w]�JbV�[w�4�����Mİ�ȸ/��x:Ƽ����V��ψ����p��N��9[իR�{���*!̌��|���Ӕ��� �F ��Z��!/6���ec�*O��E��L`�C{cWT6�$�rs
m|������/
�ظ~Q�W8bV�e����J
�� �!y�Pم-SS��{g(£���3�$=�W!��غ_n�`����D���g3~T���!�������.�2�zp.3��A�<�X�v��t�y]�h�`���S1��S���X�pם�Z'����SuC�����L�O.4u�Ү��)���5`|�ڝ�(D޺�q)m�h�:=��n�p��'N����l��C��rn��;*�ڨD����
�cPa{Ѿ�MR���"����w1�{y�7�bƊBcIp�׀��bȫ�"B� Zj	2Sz���әa}ྛ��j^��f �w/?(r�YS'�%��׃Z1`JwlK��*����/�����{N3uۙ�ۍ�35v%<NEX��H��-��_%)�&�t�f�}���-U�;8nX���6��������K^);�
�{Y��ha���&���.�5-)I�s�b'�W�&[��'C!IW������
��ehs@�F׃�M���&��l04��1���vtv�fq9\я��|�w۱(k)�	�Dr����ާۛ�BY��:��H��N��U�S���ԑ��~�P���4/>�|�4|�w�<�3�ܺ�NF�1�х�E9�b��3�g���gy C��ޔ�A�
�;oP�qȻ��Ө�r,�� �wSM|8X6���yq�	�q�ew?o��溛-?^^�N_9r�,�W@��z����XN`5�E���Ua��'gʸ ko�=b�&���!�𙽖�:ww��[�֮n5q^֚"�%�p�&}⁖�ϒß3U�<�.*��Utҿgo-w�-I��,�1�u���_!�)��ZwTc�Z%��AZY��w�oν�y�Ϝ�&���Ffb�u��a�6���Q��eѸN[*Z��T�i���n+d��'5K;M=Fr�[����~
��-z>�4����鏟��,04�[P��ב�|o�E+nn �X�]��@��T ��3�& �	&əѯ,�r���=�������%.�vΩ��h��� o�Y��{�1�) 2�ڜ�^���5�;�K��/	E4�$�Y�x]��^�z��So"J۷g��n�5j�Nث�|itQGj���\��*���[�(��k+��G�U���bΘM��#�۴��F7�b���:f��;j���V5�^l�� �e.�v�YWuЕǰT��N�b]ϏW��cx���{��8Ͻ���G��N�ͯ)� 8U`ʅa�}�U�\�cK�>Y�m�-ʵ��¦�Y8)Se�b)ϫ�{ވj�b��O��>$��E[�����H������SԽ�lMo�P>F���u����&4C��u	�'X��uPEl�Y�ϖn���V�T4�D���ʬ Ǝ�V=�{���4i��:}� =�(xf�Q�)Q-T ��C[a��9:����3�(.�Bq�踗/B�5��$��l�S-� ~� S}w�-�|9��]Rw�wTT=޸Q�"�l�,�וٌ�d�����7Ɋ��њ 8U;�,Y���<�0�;
���*��R�nI6��Q�h�tv��3V*ó�4� ���਽�X�v�B�R�L��p��!��S��<.z�FZ� ��NN93�j9r��W�3���m�4b��5�J�1�����_:�{�B6+�8�7Z0=f��׍��k��Q?�՘���f�P�G��˭fJv�^���w���?b���xe��"e+�֎��,�\�c{J���V�ș�����/�}W��{ֺ>05�v�xY		+..\���WӋ�@���Mӗ�����
�/��vP�Emw-M����P���,����v���e�}0�N�4�l5z�]�<��fF�Ls쮢un]���!�K��=*
�����+�OɈ�R�ɠ��U�Ӭ��gW��CV3�{���a(T+I�߽t�Y�+G��
��4��>@WY#F�Y�K��h"^�&�}e��� ��c�x��7��Q�t���� �d�7�P������(Ο=ޭRL�]Z�%,�B1��t��7>u����ܕj@����������)��쭲v;�Hq�,ݗ���Ē���S-/I�n���ӵ�+��F�t�kx��h@H��Ucm����o�F��
���^�wV� Ӝg۲��%�[U�b��E6�1�!��]Ehİơ5k��sC")�1�
Pw���'-Yf �O�w�
T�V]{\L��a<h�E7SJ�$���4�92�Nd��u��Go�����}qûb>�[��׬{�'��S"����������3�ӥ���xZv�^z>���i��}^�J%Ր��σ&Xv�ʇ@"&���>�,����Zl�g����m�ǯTRI_�Qd��(7Oz��'e�3����#�b��v���s�*��הY��5��x��&ݓ�Z^���H��[~S�b�p�cx�g��T�U�b7wIOXG��n�agH	�b�M����8�c��9s|b�/�T0���uW�U�4��d��s�Q�}�.� ��^�t��&��w�3�< �u�l^y���+B1p��_q�г���ܧ�q���h<��ӏ��U�5}�Y�~K��R���*�q����z��?52��rL�H�-X�j�~-VM��2��n�_6�};����gW��^0�����2gڔ��ѹZ{�vp���Ӊٟ>^;(	�W�����Q.��論�N��ԏMY����s����Q��\/ܽt�E�'��n��O��X� � Y�k7r����ho
Q&}�v�W�E���ϝ��1�Qi'KG�����ѯA�u�s�e��j�ui+�8�oB}UF��@W�hM:��)j��B�^�]��΂N�K �j��P�q��
n�z���^������K�|�d2���D6��3���(�RA*c�ey������S'�+}�9��J�1ꙍFժ�BE�k��>jO�x�}O��6�n�Z�M�v=Swf�KS��7��*� G�S�xR�o�"����3�F_��I_}��*�_P4���,��X�����n��H�M�-
���nq33aq��"\pI��t:)��Vb�ɴe̻��)��J�Gm�Y���8𷳅�\G>�:�� r��?��c�\�t�y8 ��s�e��-ܧ��X�:}�Bۏ�Z�܃�l˶� �y�i�V�Шe^V��rn�{�i�j��֒�<Z���%	�Է2�� ^�ّ�xS��U�Apm}�=f9{K�ظ3'>Uջʸ=�{�gWBMƚN�aK]�wu@�:�(� �,]_e\[|2�U*w>|��.� �9�a�h�p��fʌb�v��ާW�WR�&E���R���w�sdc���_ҵ�m	f��V�;6�Kٕ2�J�O/���si��#���Ʒ�F Q�"%uk
#u"�Ɇn�wu��:gM��ٍX�|� ��.�r����Ćm����w&`�A(ec��;L\��w��	����&��D�P��l�7˱�q�t�2�E��Y��IN oh�n�Y��z��Uԫ��J�@ﳋ/-R�!��ԫ2�+��q�xl�g_oה��m�k��ʴ��X�`4�D��5�*5��n̋QiڲT�z&�7�|��̹��6�b��]��M��^ٮ�b�.�;��7�[�	�s���n��⭜�K�!�[7�B@��qJދ:p�5�����2�ݓlVp�,�	\��n���jj^ѻ��byn��c��6�3(���n��8��3zwD��&�s�^`z���'[0��)�f�ˉ�D�YԏD���ޫ7GX�+Evʹ���U�A�Kie_[�c���=d_ZMc��{i�:0ue���4N�F���nֱ9��*�h�!�ӺP��=�=����R.�e����mvY��q��MF��f�e�g��������(k���&�R���f�=U��i7�ϲU�4e#��*b«fJ��+@��eHc�}�sQ�Z��o
]�2l�j}�8)u�ֱM��i���dI��Q
Ic�A���(�q��Z�m^D���w <=uԖ*�@Vv�n��)�ئ�e���	 PpQ,1ѭrӼ�v�e"�U�O
zA��A�v gP��W��[j� 鈪�x����L�Rra�,([W�_��|z�޺�T�Z�,���>oG�vn=bv�ې��R'�q��3@��s���=i��Gm=MMԍ���Qf�}����CP5����H]�z*O��&▍�mwfn��g�7#�v�ޠ`F��Vne�{���N3��HF_,�b$�ש�ך��b3�� d�gz�=����3��6Py�k;�[V�cq3�
��m�9V﯀J�5L�Т�|�z޶��g�՜{\G�N�]�����s�1K�E�-],��r�l����;�}�^Į�:�>�n�V����_ooA��	��\>H�ڣ���v�\c2�����4�e�j�+����=��M�
����r�I}�V�۹�9�gA7��Q3(��j���>�����N��O����8A*���2��
�P��W�9r��TEr:w�**N'(��3�r"��T�T�TF��+�(�*��W(*��
���\(.$��*��*��Eª�����)��i30�$*
(.*U$Ī*DU���QL�"��G*�q����)9@D"�PȪ" ���".Dr*��I	DUr(�ʃ��^D#�*˄QND�샔2"�TAI$TS��#�U�
�e�.PTES
���s�2�S�(�����U�9�#�L���yFDDU*�UQDr�'��r�\����\#�r�@a��G*쪦�\�Ayi\.�(�_�/�O����ϟ���B|�P{I9����vi�h��sh��;���.<+Jɏ�\�"��؝�m��ĸG$|�lGxo��}%630i���?��0�����|�n��&N�<�:E	<C��<����޾!� I;:d��n�$����T��{ό&#�۽���K�iē����0|�������̿f�q�Q���'��C������Tޞ�M���v�s�}��N��V��>>������ι��i�$�*ɼ��V��s���?&�8��'x��q>��6	�@ }�> ��Ʌ9����YY���4g)�"4G�0�r��C�}���z����z��{��?�w��)�Sv����������!���n��o^���ێһy�8���:W㯤��P@�� d����1|6�^{^�O��C㸇hv�}�`�!��;�����®?��~�;M���<�^F�'����Ӊğϯ��pݠ$����s+��&��Hv�����u��>�@��Q�s�vKMv��;toN���o�����w�i��wo�m�w���8���η���]㏾y�G��q0�>��[(��q;�{�6��eӸ�'�`������n�3��  �xא;�}|]�]:W� *���h��I�����Qһ봁���#�o���N���t�v�8�|?�q7�O�n�޻�F'x�|���{z�O���C��zۺ�x�o���@�0>�B�.ƽ��������W	���8;x��}O�;N�|N!��xn�'q?���t�Uߜw\~������:L���n!��;��}C��@�'z�v}��n7�I��6����G�!v���9�ޘ���:W�����o�פ}��N��Wn~�|�}��;W��=���S�����~��ۿ!Ӹ��?}���C��r?�'i�]��|C��P�q�oP�q����b�����v�J��)aSw4����!�ם�n���~s�iS_o]�'_}�������{�1�����q�������n�|<��o�t�7�����Ӿ�����:w�v�]��;�S��Q����z2E�W�Տ���йB좇�}��s�eӿ���{Ѹ�$����:ݻ���@��y��
����|9��8�~��y���i۳��;O�ݼw�k�>p���o��N�m0>� Ǡ�XTY�xj�G���޽�Y�[��5m��� �=�o�l䌺
����-�-�U�t
?g���P�����6�{6 �-Q2���xj�W���Bd��|�R��`b��j�<����n�/S�U�} �M��X�G&	|��Ǯ�e��
s����O5�F��끸G����BG�z�&�q�U��I�����M����i��w�u�S����z�����y��z���x�{��aC�y�2�q�8;��u�e�=v�!��x=��;��t�y���=��~���w��c�ɗH�;�q����﮹������;��:v߾�so>X���ɻw���ݑ���lpF��z�����
���;N&���|C��!!�~��Ѹ���w�t�����E������I��7O�	�}]!��_�]���Ώ��v�;K�ל�o];�sq�폦�(�Lz۷���Wt��ס�����7����N�o�w�x�|L.�A�:qӼN&�P(
(~O�.����:�/v�$��]�y������a�����F�]�fNpG�E,��2\z���i��[��<v�x�=��ô	'�����1��B~'�=�;Ny�ӻ��}�t�� |<�:v�i�'��.�C���v�h݅o�x���D!X��`w񹼋�~�߄} n��O��pߓ���ލ��㷼�>A&_�ny�]��������n�:I����y��F$�N����n<�1?��n'x�zt�:v��^��ޤ���<MǶT�Hď���#莣">�}N!�5������;>����q0��?y���z����޹�o�I�BO�=�}��N>'��s�}IĔ7����  �.@T�&> ����|�a� C���n�H5�""D|Q@=��v��?�����Ӵ�շ�~���;��m��;׉����A�Q��&����S���q0���z�qާ��������n�v�p��߆0�\��
Đ����B>�A��������V�q��n�����v���L=��G�j�Ӿuc��=v��ݧ��
�?]������Sz����:��|�1;�y�[r���:M_>��|��B	�e5���+���^�\��}V����s�����g�y����y�}~;�ӎ'�
��&x��<�����8������8����	2���>���;��~w������צ��{�d�oݒ嚕oa@}��.�Kۍ�n���	����:������{SE+�A(3/�mjʶd��K�f�D-+�p�|�@ݍ�9�i����̳Nµh�$���+;��%��:���8�����ɋD��b���7������$��a���[w��
o�=�ރ���y��{�wn�x������=��۴�����v�������N'��o��ޡ��O�G���aw�û}wn���q����1�p���փ�rިj��yH�a(`u��G�z  ���R_	���ۈ<���$��`�o��n��S]_�������n�������:w����K��]���0q7�������c�*�O
�UT���o�w����x�p{��x��8��N'���(}>w�G��ߺ�7N����^\��N��ۉ�{��v�U?���9���z�b�>;q]��{� c�L|�oNY'`Žm�.�����nsݼ@�'�h�N������t�v�9�1='�ܭ�?��>���[|��?�L*����߽�����yͽ~;����w�7ē���|=���#�"D}rڧ�r�v��gG�V9����i���8�kg�e�O�X�ԝ��ts�;qğ�Ǯ�wN��o�'o~��}��v�'��??��_�i����������C�xn�}�8D��>������
\�v�x-���~���!�=:�P��L)��9�����~N8�Į$$ߙ�a�7���?��@�'|��N:O_��q�x�!&��o���BC�k��}�}���|��}i�y��v/�hA{/D���=ğ÷�v�}����ym�>����p)�w����|��;������|gw��n�-�~q��;��.�
�(�
=O�q0�c���x����R}�G�>�?}4���0w3X���S�̪�U���L� �/5}�q8S}����q]�����x��������n�<I��z��v�7������ۤ�:v�oω�~����T��E}@_?~�,�2��I���=>2n�A�ǡ�:�ǎ�?8�}1:��F� ��g�N��!��$G��pz{I�n�_}N���	P��)��Z/6��S{��my��n��kx�Uc.����wkt�4�Y�۲-��.���ˮ.#}��/v����Q}1��q�[���N����F�N�tVj�&;��7�"�Si�G��(^q�P;]A�wSb�a����D���j��[�}�p�H��jr�/^����:�M�饠�˺�u�2�W� ҂������O���+B��6xzA���ϩL1�
G|~Z� ���VY�F"`Ʊ7[+Pw6�,��)��}^�S�9Z��ejD{�@hTN"�dO�Fյ1�-����U�EQ8lh������S����"��鏨��&��;f��A9i�A��^C h�l�l�pr���V=GPU'jo����á�+����!��.0��uJ�~zj�Ý�a��*�c�؝�WU��zoY�=cz�Dn��9]@983Лb�y�JJ�+B���y<���ke���k>�梴|�,�gt�*_y܍�.18�g�e�Ӏ�Q	�`�*0å�4�Ӳ#5wM�\׳�
à����c/�g�s���&+�!�����N���'㽳���[�b���1�u9��z�nʳ;��p��^���*�/a@N�\F�O UX+��p��/���sM��ߜ������D 9���qV��ഷ�l��w֎�j1G�ε,*h� $�Z���bs��s���/r;q}G �p�3�X+�=��Ps�����f^��=��m�-�]Zn�L`)}�fp����|+DȲ�#d�j�	N�*�E���^��H=�80�ѷ���O�(]��k�/Nv�*Td�h+�`�M���r��J�������^�Ľ�#�I�9�U�����u�>I]bP�W<�������W�}�N=�uĸqq0.O}�=q��
� �Ӹl�^��\�h��l��:	:�,�z�����W��`��EL�F�gЌJ3Q�����!��?!�m\1p�q��V�4qЬ\�^�W���x�A�"�A���z�cYT����R,`����"�8uFN��P,��y~���{!��2;�����@�:+@_\ _Z�k>��^
[_l#l��^�)ᨡ��;���T֒�q:be�͘����b��!�ˉзB# �h��F�̘[v�������)��xa-��=�y!� - ��[F��+O�`-�>�)��)qW�?�3P�&�u���:�`�F,	���7*�̊����2�Oѯn\[7���Š���[�e�A�eޙ���S��&M�n�ן3^�6~�%���e����;3����0t�z�o8W��,[g�K��饜ƸQ�]�'E�����{=V�4=p����m�l&�$��#���X��a�W�S�<-�i�8f�덏'@�K�����)�R�X��:�30g� ��8���oه�]ַv���xu��P:����N\�|���=�ǔ��z�*��e*@��nu�[�xK�
u֧�Y���(��.�����z~��v;�94�++<e�J����C;o�!#������&oVp� ��`��ޔ�ϻّٽ��Y�n��5��j����|<�q�w.4�� �3^̻�t�\'OT�2 ��{λ��o���uEW��9�械��N�}Xʑ�U�kTݯLޫ�P �-��uP�����r�h���V�y9B����;k��Hhǵ=Mӕת_a9z\Vd�.(�o�Fj	D	���FD�b�.�g��C���b�N����Sv�ʺ�ܱ���g��(1=A.]��9E}�ڌ*�W�(]N[+!ڿ���g=��7�d"S��������������NLWOL|��j}U�}������m��E(*���l,+�UX�f�*��Ih�__^%.^�^���z<6�v�NdCQM��f����p|W�6�W�n5�}C��TUe{�Ǹ�4�V��H�X~7~�������[�b�M���'@y~�#(�(MBuR��D ���!.��`�L�#W�٘n��a3_F-���Is8!"�M��{���
,�D��Oj�:����f��Һ{+k��v7ug����#K���C�t�q�V�<�{��1PS���
����;������ήB+��o�ԛ�.����a���N̑�j����RC�[>�%��r������wL�p�}c5�=�O�����|>����f0�@�|j��X�鯰��Z��)�Ɔ.�D����yߋ�IU��[�{͋�����H��8�^?�p�5c�s��ht�RB�ff����|ݡ�r}��~�g=�!]��ӯ}�Őu�FrDV�q�.�V"��,W	^�}�>��^�9����|D��h���#&\': v�����U��F~����4>�����c�aoe�~��:�^Ix�W��m+���_�΃5e�
}6�Њ�R"��&�7�-�����jY�;K����i�}�͏z�6"D����^�IXT$�b�S��x)<�����+�^��{Ԕ�>�uZ��:�^�;/qf!� y�Ե��R�G������K`_��xa��J�*�����ںӒY���|����iFlG�=�a������y��Mꚁ榐XiT;�zwf1���v�5��+��+t�P+	��b�.C��C۵�� ��[��Ye;� ǳ��k���kN?��g�#4�&�u�,���ݥQZ�F��� We�4k�G���3oL�O�Lѳ�:o�R�Z72�LVW��fA�
ɩ���lͷq�ˮ%s]��6��;���.P���������m+
*$��^��E]��<�����u�
P�wo!���S�����v-N���"�k��5�T�HrV�"�*v��������o��T��Y���2�0��|��� �x�㤝e}F���?�]�g_�1-���;��z�E3l�}g]m|���/���k%_��{5������G��y4t����:�7s_����>��Y@�l�����L��R0��_=�#i�q�:�V8$CS
����\y��{�{�hdYd�=�hB�/M����[��²V�xW�D�*�����\�u{��1�`����>� V�@��B�L1�
Pw��Q��c���ۇ�N������a^�e�hJ&���O���t�9��t�;���~'�t�a��p�݈p�*��rdz}R����Vʻ%���S%�r�� E��1�tњQ>�>;Ռ�3^�8�8�	�ϓ��ōȫ1���ĕ]�:"����f����	�uJ�����Ǉt�B�z�7Y��3�g�JH�Uh�Af�^�^��I��;�#*� +�����C&m�4:E\��@1Fr�ߏ��A$֍�_x�-��p�;��.\�4�d_�B�/fv&�\L0EY[^�����[�J�����WGJ�mH�J�me���ͯ!^��*X��q��yS����Cu�o�i@�Zu'C,շkp����������ՏkнŸuۖ����X�!DF����p������9(���G���*uC�2K���ِ�¡1����@�3����}�}UUMhu�^B����	��Ư����dܫ\�~ۮ�6�}+��|pU�̤Rxl���We�I��lB��C>�U�v+��U���N̪|�vx��A��K݆�Z�4�>��r�=�S����O�V{�>7��
�Gk�������)�7�F�u;�:�� q���k��'�<�+�/=3}��퍌贓��=��ϯf��׏�^Y~�F���B�e���]C����6b�c�
�r�v-+D�Ci�ѕ~��WW���!�
f.��xk�2��kY��~9�������X��k�.'"}�]���v�w�\�&}]��8Z�Ǣ*f5��j���b�X�t����>�R�P0:�wd�7q�߳���?%Ǩ��h+��-��`�S|�!"R�����`�=5I�^�s+Xdz���u�M�;��
�?W��i��H�`::��
�%f����d�'��)M
5�mli��#��ġ��yOJy�AM�Y#
����@	�mS�N{�C�8I8,^v���e�Z38h^NWڭu�����"�v5q�ǡ^�Պ2��؎�τM��(r�]��7\Ot��,��:k�7]EclP#%*���O��U�Ce�WY��^b*pF�W�	��D�<�)�E��[��O�X�S�E�������|> �%����CWE0~��V�y#d����x0E�uL�U�f.��m����$�d�A�TU?�b�EK�Ѧu��J�}�jafNi2svb敀:����z���j�ה{����SR1�W�^�.[g��aʵ�_ٲ�g�f�"(}ퟰ�7gD��e{6/��1��]R_	�����(��k�aU������jV�1	�k��T�`'իp$�t�u2]ؿ{�N����<��Oe���g�l$+�V�z��V-����vq>�O��[/���[�ᠣ��N����4 鿱����.�f��2*���-��a�c���;*�7j_m��O�L �c�AL�07�{9�~��֍�����r�pa2�A~�[�`��ѡ��ߕ��|�e}�-Q}���T�yAvc<�B�n��Ɵq��-}G�@�"6h�,D��H��a��ªF��E2���_ޟ\R^����a�$9�F(��dT���D�OQ]�]�pRZ�F׷��-�L}?Hc��u>U�p`c�>Y'V<X�OM7��>�P٧��^����9�xc����S�|K�DuxǛ��N�jР|���w;�����kH���ܸ-�j��(�G�Pw�D$1 ����>�wZ'#5����:NH鳊�jӝn�<���oU�[5�r�q�K�^�$��IU�T4��m�YI��F"G�V�>x�s�N��lίqU�Z%=B�^�{�6��έ+��C��-/T�s�9Ef���WrL���k����u8���s2�%�.�
R;�����2ɸ��D�]\�X��Ӭ&�a`W�',Q����8�����*i=��`�5Lۀ��1�Uŝ�o�ąҥK8��;�V��g�Սd�.Q'�̺x�dr��\M�Mƪ��#�݆V�3�wv�q̢��|GK�:�|�,�VT�79����J�vsVťu-�oiSq ��Y��E�!۰]�O��\YF%��5U����u����C	n��FҔ3�MC������!�Ԣ�VU��_h�y�:���9�9y�d�Z썣�)U�lآ�)%Wi�f
wq�F���f��q�Fd��(vr�������V�^Q��kkѻ���#E��f����}.�⬭K
�d�bO 4{JYR5';i�]c@M��[L�03b�ƛ�K��6k���Ԏ\v]�oP�嗺������������ĹwN�2YWkǼ&{����/n�]�ڙMm�.5}����;Vq���fsK��Δ>�T<R��r#8s?Y_Ic����u�x�wa�V1^ۮ�SP�b�)5Ց��핗%Ķ�l�u���峵�V4�V`���\�ju�{csL�}���ܸv[�\p�Bp/g;C�kH�����or�Yss�.����*��f�VD� Ţ�z䚃�F��8vf�t�ݭo����C__g%�;��/�S��Z��TK+=Y��B��w�������mu����^ޮR���*�i66������N�@�����c �S��|ueg(�g�w<nu� �����l�ݪ�V�_�v��j��g�]�u�x��;�:e@�ܮY��]�o^cZ��<��sZP���%ŝg��!5��@˝�5������i��Yu�u����gGn�v#{@iNsG�57tHg����J��w�����7S�1j�ccy;��<Ժ��J����t�]h�j�	�F2�Y�v:U�QbII���e�1��m:4T.E��+�Jr���ށCU�P�F[m�����nSWB�-��(F�{��v\�0� A�ͧ�oV�	-�J��z�زm�Kw_]�c��Wr�*Ś[��P�S�dV3�y�X�R�K�^��^ZǧM�@�u�뵉�L�YW��/I���.vj[ݳM�o��wI��kR՜X�gs���VY0�-�W1vU��v �R�����fŹ�v�@iL�$�C�zº������_q�6�'rR �W��m�LL.���߾��|���QW���VvDÑI4(�W.�H�r
9L�\(��'9W,����(�EG
�.]�TAEG9��B/r!D�(��\���DIӸ�	Pr�J ���9�9ǘ^:ETEL�*�DG*r E��ʢQG�Q�8�yhP�p��Ȃ�"	R�UDd�A���<e�*�PEQQs%�UW.Dr�$E*$��.�Qp�TG.ª "��EG"�,FnZNaj��93����(����\��]+r�MQPF��T�Ih��b��K0�Ur�M�rr��ʊ��&AgA�����������g�A�^1^���e��i:��l�.Ǝ�&�8��xv�G�s	+�|�	d>��nܙ/&�,��~��� 2�ͻ�:��Vg�o��O�!��y�X�xO�U��KF�믯�Kwu�Q[)kR�v¬ѬKF�G7�1��N�C��l}��z J@�.R+c|�Vg���X�*�j
�ɱkˉ:�4lB����N��6�0FQtP��/,�� p��e��=G_:�^�����t=Ca�]��nϥ��>&H�>��R=����%���ښf[������I���Ǯ�`�����X|L*�5m�q�ƈb˜D�&��F�z�zq��r�J�����UA�$-�p�B���lӫ=��u���Z1I'e�/�8���V�V�T�"ob+8*u��|Ő����En��]��J\�e��.���\�7~���K��mH�L���?`���,�����PYg漮̪g�{2t[ÖA{~���ބ+�P{w�
�]�c����K���+�J` 6�jF٢�z�L�Q����ݤ6Qtn���|5"��!���:�uLN����>�D���v����}��DUJ�,���&��'`��Y�������Z��27ٹ%^6I%��D9*�E��E�m�]�j���7snU�#n[H=��sBT����d���P,������<v����H���*r�aũ�[ž��x�;�ս�nr�`�\C��t=̑,�$���}�����wfϕ��g ��4��,�́KZũW�#�N�îe��9����I��@%�ˇ���F��W�Ö��?u��>|��L<�V˭fGҝ�S�Bn��e��<��S~��53���(T�>a���rvU�=��JӺ��߶�IFߘ
Q'�:!�9H�s���df�MeV�x|�Q��$��ԤF��5�ͽݹ�wj.�С�>�n�b�0�^:a����U��`6
5�:I�c����/c.�w>U`{%9ƣ��:=��2M����b1)�8�f1���m!����1Dz}\������^�y8��='��H�� x|ǆ�_Q�[9��&��Cp��L0���"6�۲2�Z*�˛��t�b~�Gۦz�v����@b�A�k:"�B��u���n�1�ߥ��Cs0-���	�d�I��(�qN�"�ό� V��;�L.5�(p�;��N�B��j�&T�l��\T%�
G�3J. �MBn��sn┙t}�$%D��-��I����δ���yaywE\�V���Kp��ӹ�a�)�L�'M���-���r��ծ�B��Ի�c6�������;��&�p],N���.m�)�5�o%ب�<<��^���]�h��ݐq�i \Lbû����u{MS}�N+x��g���������-�S9Y"��9��M֒������9c�*�ɿ��/M����e��㎂�S�3��̏�����g�Q��Yhd$���Q�����C�tx��/P�9B�g~�����o!1#���ei���vP�'r�R�,V�����#(h�o6/�ic��{�&u�ȇy������k�t��#[��`��i���̯AEw�g�~��\�U��Ւ{{��&�'�j��pp~��uaC7�V�p�-X�_5~?5�ɻ�@Mc܄1UV��q���')�����c�^�o	��y�4�AY�{*�"2���	�8r)KTa@@.1�x��x$�N��M\��!�O^@ȗQ�w>n��>�Z/�m�b��} +e��Mv�����{�z�@+�> R����Z��9b5K�=�k���Ʋ�m$����6���m��=�ʉp�D�^�����I�F��k5�,m���#9�N�=��k��g��X*e�p9(�Eד:��`$�RZ�^�!����9\iqN���)�j��]wC]kq���5WMŪ�!��;� �ٳ�v�Z��6}#�EG�:�e*3q�X����S-V���O��^|�&�Y�H���X��Ȳ�ܳ�Cl�>T��;gGO�w+��W�&�Io��@�sz��3Ӻ,�!\�Wj1o>}�2�)w.���3k��۶���T��.��D7�Q.����U}�+M�/Я)��>��D项&H%�:���3ͫU���"����#��b�tԨ�	�NR(�s��W���VD�z���Z�k�
�-��`�F{]���>e��h����z����{����	��/΢|beOɹ��^���ۻ���9�3�Չ<�gk2��w�g�e��
I�C�k1�ǆM����Ӆ8=4itH�'���Y�e��f�4ue���$U��U�%n��^^hŁ)ݰJ�s1~���w�p#E�qf�����Nz����i��3����_,�Ba��&Nn�C��J`IY�W��+�h��]gy�'�Un�}���j�ٱ��Vw�^��:p�3�fmR"�������n�o�z�N�A���/��d��@z`�5���PUc�<8*��1~(e�a����K��i~�JOwJ����8M�U�����;���� N:��ٮ��{K�,[A���͞n�R�U�}і�!��t�Е=s��hAӏ'�|����s�φW���ָ�z%e󘙬`ۊ5���Z%�C��ՙ&�1�.9Ա"Z��������F��Y6�N��X�˕�L!��j�գœ]3w���e$Ky�oY�y� ���r5�vw.� ���P�����]^wF��2# ��a��J������g��%� �8{#���l�_���z��]�WUT0,�Ǟ�y>�5�я'(�G$�ģD�U<.g�h{ٞ8ۑ3;x\u�X�4�ex�@�1�oL����f3����:��4�����#9~�͏UKGM��PK�KکqD��ªF��FӖʫ���z�\�fw\Ç~~��M/yp�����
���Dm{y>(Wn?�`� �eV8����-��<�[�����5p�!M{�����I<�+ ��<.�U���o�f/���/o^�ǳ����z�t����%����}p�45	۸y}S�U�yYA|{��>������sqsn���e �;��	6������3J��`���4�T��@	��X��bŷ��_0T=B���]�o�g��N�8�pBG!ϫmԏlE:���L=�:��=.�M�'CU'= :"�J�c2zpx�^ն�Ϝ�h�,��OQ��v%H����b���s�ꐠ=��R�/R#�8�^1�l���xܙ���
�Q���>���Yg��[���]��䕦D���k��]�cOR޴p���Q9pWzv�E'^����W*�Ԏ����0�ܭ�.j}�/�g�L�<5f�g��]�ڠd�MT]ȓ���udd���\)R=�;��|��W�U_}~�iT}�Տ3,����#��f�ⓡ�
k)�D���ت���\�\-f;��r0�Y	o�.�v��J����j� w�|�~~��s�F���҃#��H��M�;;���n��X)?V>��*�y�S��x�G��X�y1N�����Iڈ�Җ����= ��V7�M�б6i��F�^Y5�35@�.1�1;������2���,LV\���x󸗋 :k����jǣ���}ĳL�KZre��'a᯷R����)������8�s��իǾ�����g-/t1}�(͉��=�ְ}���®��=y��{Ў)�M׵�p��w�PU�zf���V�B���Ep����B��!�l���k��o�Jc���������YB2)�edS�g�#4�Bk�Zr,��~Zf ��S/L��m��N�����[^�����8d�>�b���a��t��u�¦��T`�_#���>��񮬨���ۜ�gxlՠzS:5��rP��J���z���߶��u���M�KE:.�uʹف��,�]����h�K9�����e�W�J��z�9x=����z%�.�7c��B�֤*��1�{�+Q{�B���/���`%bA
���:�]f��9���mv�� ��ق�������]tw��I4��˲��+E��?������ފ��u�h =��'�O���1��:S>�K�s(nJa��!�m��,�9����^�K:���:"��uL�9��!"��
1��N4��69�fU�s��Z|�0yH�^���K%>��sg���j����U���U}r�s��yH,Ǟt���[q�݄4�QE�1ۯ��9�qW
���Ԉ�A��ȿ��4��i��i�2W�㊛��y�-����
~N�1a럫��i.`y�",	�鏪
�roN��~~<�W�=�c�=�CJ��F0d�T!�tǡ%WF��`�nX-#<\a�1���P/3tBuB�-����z�a��l�y�h,R�S���:|�����E�{t��aO�QZA���u�&���ʀ�
�ţe_s��V�ۜ�`��i���̯AEw�g��鍥+5�r�8q5W�e3Tŉ���!����]N3�D��r�%X��p�욝�Px�d'���@����l���|':�b�0����v�^��<.�Ņ����u18�MX�&ez�-����^Eؽ��.z:=8�G-*	w9C��l��L�F�����Tl����ג�Pմ��U�V�a�7��wJ��q
[�aT��)��}��R�1 ��@*�s�7}�����w9`\X�L+%'ļ�:����>��mg�ͷc*���ʚy ��g��}�7z�y��EY�%z��� �["9Ϩ;�i+����>�v';@nOR D�� 'uV�5���]h��׷�u�6�-$����׼�����A'�2��M|!��p�7�6#9N��
%�c��^�(y��AD�n�r2���\�ٯS8	<�,P������N"K�Q�bv�s�r~>!���O���Z~�kv{�d��~���*�x�<g�Ȃ �ՠ�}ܪSJ��WN&R,`91S#>ק҄��9��}y��NO�ã��'P�8�̳�Ug@��� wڞ'�������K{����x$8���q�:=��n�?;��*~���\Es
�s�m���Vcu��έCڀ�lX��כpC��1�V�F'�ۯn��U�dHB�� -6�$VЛ�"'%�|�!�Y��/k�n�g��?!7�5TÒڟ�|x0E�1`'T���gc޵:TV�r��������������|w��״�8:�w�|�-	�d�&�n���}����~�u�5��9���(�ݵ��]�b� +R�;-ӂ�G.�������b�NU{x55�4/�)��2qF��Ǧ�J0<�� ��Mn��1��(����-�op}U,:߼�;��2[&�]�_v�ʉ�{1DK\9����<��6��Oﾪ����YN�[���_@;��eQ��?�`�|�m���;}k��볻�3W������y�5��s�Ս�����>��=��LF��vQ�+�����Ԭ</�U�5(짬���}^�[�6���dh{� ­��]f�L���Qb�`�<~�VƷ+�W<�Ӑ��z:���A���캍
8���s\Ѓ��<���Gm)�$T3���u��@�����Z��ʔ��b����)�qpS������%�wS��y]zj�(���z�;���@>E�ȗk�Q�TL{^��)��.�ޣT�k�j�����:�+r�Mx*`�T���n�¢~�E��j����5�88�ۦ�C���E�f�����#�����˹`�n�&1*��Ӊ�
����/Si���2}�r��G��=�`Q�uu�̸�F�l8��S�6�H���4��?ꇚr�jݨ~8�}y ����(3{>��E��7�E=i���1����}�{����iCu9��I���h�����p륔��4ne��lBc��p�)�v�S:���$P�-_NO#�32�Uһn�b�j�f��H�۬:�S�7-Iw�܆\���T�����T}����>l������^)n�6���׌ߥ�5	�k=S�Fֵ�?Lm�Ð�������j���7��	����Y�>��8p^PS1��C�~V�gO�*FW�-�#V�^w�{�kL/��@6��sF�_����S�؇g����{���t8�yH;�����+�_��*�r^�0���y�7�\KV�}��6��|9�k;�
B���y33�w�r*�\cy��'\Cn<�7��u�}�\�;�I�ݺk�����]-��n���m|�U�Ѳ�l�~͖�E��l���!�����A$��fyҞ��ʪS؎������?�����g_'��y `��z㑗S:�Ne���&�*'X��.���lΨ	⋱�Pz��;����$Ľ�D���y�dx�U�ۅ[����w�v�B�����ܼ&H]��jJ��m���sa��gZ5n�!}S�eHK�<9�r�^'gKs,R�d�map����|��R�)�f���aY����R�Ә��\���u>1$��[vhvۖ�;����>�9�X�bĠ�����s��<���Ÿ�]9;۾X�].�s��=������ju�vu�ͳ:�N8���S��{Й�7KJ�kZ+T�����;N_�V!O;�rOJ�ɼ놖�4䉹��[u������J	0H�-��G��ذ)U��d����\8��}��]J���S�eL�@n����f��Q1���B{��,�6��o����#s>,�R�[��=X|e%j0�v��RV;�M|����L=���G���X���j��9������.�L7/$k��Wd(�t����]��R�v���>��:��z����(?vL�G���51_C�˶�e�<~���9s�fM1)Mm���;]Ţ�Dx=�A��ҥ�p�_I�Le�]'=\����q#���҉�GV��7��fVJ�n`c"PB��1{Qu:�k�]�צ���.��<�b����[{Y�	�iB���Ug�e�����W��(u�i��f�ڝz��7���	�CYc��o�8c
�ē&��_vR�!v�Q�X���ԶoK�������)�,oB)_lM�����;qrf�u�ʷ�Q\��F)�m���r��5��t��Iyhe$����q�';��z�B��W�]0�Km��GWN�\�(�Z��ht�f�S��%�'�|;&�{�,�]�XC%(jT
�?_Wc�����õ54M�6����6�T��cf��y�P���a}Z�k3���ԣaެ��Sxx̭)K�yJ<��+�Sgv����.��荍;����Cq"�_%%e��.v��D��L>���,��Jf�c��n��3�Nز�ʶ�O����jV���)Z+�%�x��؋;9Lו�I��̙tT䥅a-8ث��'0c٨���LgR�<H���.�ohY��x�d�EДF�zG�/�P�X���;��Ż�w�:�v�g$�\����nN�)�;�ʱ
�Z�Յ�wi<N�8�V	�)c��D����f�R2.yc,�y
�;�};��q@�um
��GX�٘�U�1�WD�v�M�k�Ӭ�T����G+ڀS�t��zu�j�哿nWV4|�5ѻ�;%�s����YC� �eV["!l�i���9��}��p¢I?�A��^�ƇZ1���W�M��V%�*r��"���[Y�
�4�他	���C���]��V��3��[N�d�B$DC�=��:DKGrK���V�.��VOV�Qd��l-�k�}/01И�8z�Ho!�'��&��̨w5�;�Ꮸ�H�00mm����<W/ ڠ�밴����>ϔ[�ĻΌV�d�_!+ymqU��ݘ{R���Z���EͲ�ZV� 2�U�a�m�*Vr������>�*���rr�D9B(��r�0�Tp�����m2���UQw��1*�йT,Ȉԋ�2"�Ue���p�EPTDE�ąA�"�ɥ]!	0�w+�:��-b��"lM�8󋥈b]%2��U��Sq��k#�G/�"�uZ�Ib����4.��j(�9�"�NjDU�¨:�QTF���(�99s��Q*W(�As����]<䠢�9Xd�Y Jӑ���*����s��s��r�
(�&ҥ���I#RL��ZV#��y�*"���j�Z��M5�P��&\���at�#��8vE\��pt�ʊ%ĮE�j��#B���W����;�����]w��َA3�\P_&\��Q���=�.�ۙ��f�2�s���Lz_q���rP�g^�[�_n�}_}��}m�%�o����������w��^�鹬�_��^Z�Wh�/����}���k-�UU'�x��=NTSm\Kר��!4��w/����=��7ڳ��ԉ�T�%Q���мˌm�Ĵ�jsU���}�ic���m��c���o6�����6��x����rX�f����hƆ���>� ��(��<�G���그3�w����D��D�N��K|RܸK���͐	��xZ�"&&%����k6�+*�ڄz�׳���[I#���T2ϰ΁�t2=����W��}.���!��n|+�bk��>����`�~,:U�٫¦�F��n�z��So�P��|���#���C��WoT�3k}ǈ��(�@{je��f�~���oC���a�#6��+J��m��S+Yr�5F�V�k�j��~ɩ��㼈�<V�����mǝ���}�-���!��J���\N*Y�)����^�NJY�J�'O\6�iv�>|���0e$�7�Sb�n��qv��\�(eFh�Wn��K���]t�����2�mp��op^��m��QG3RA���/��Y\�b�\ktC[�/�-�A��ڈA�mY[�������W�=Gv)���V���/�,͚Y�뭼N���z�unڅ���ڒ�U�J(�l�{h����7�S�H���Ƙ�zW�\o�N�=P�/�0���a~�%��ʴ�k��r���dn���!�q�q#��͝��x.z�<��r�Tc̜�o����lLVϺ�
G/B��2�o�ꀌ�����l�p���<�<��k'n"��7q���}�ѝ�J�vՌ��8���������Z��6���=��Y:���`����kAZ�x��ξ���Tj�����7Nm6���2�X��R괅+�]��s���L�q��N8$�������w��S�{�ۓ/��������5����G�,�#i1�)hd{�!��`�Ǐ,]�;��e�+�ލ�Ր�j���z3k�z19o~��ڇ��Q5V�P�����9|����̻��5�n.C�f`N�6S�
�E�H*4bz���j�[��bU�]a����Hα5�
''B@�k��2�j*�V⧜-�4p���Kc�M�;L��#��hZz;�I&҅V�K�u|�D�L����uO-V'�<>������^���{5飯v�{���^3�T�2Z���M�����2����Ũ���c��q^ne}���CwXCT��O9|�yY�\:U������=�5/ٗ;��Z巡�v�Ǚ�Ng�=k��}��	�~�ؚ��.����ƾ>�'K�i�}j�ǝwkN���ÛW�Bק�mL��Eb5�Į>��m��C�G;�6�%3y�[�ۮ�m�[�uQ�>����!ޚ��G������t�v�_���IrZ����Z�5���[��z�8f�-�>�N}Z�a4�V��Ϧե�R����ی׼���=�Oa��EkiOg��񪙜����������[�x�Fy��9���KvY�i�&fi��_M�T����7���=G��~���N�s�1 Lɬuz����}<�g�NU����WT�C��k�)���̛�a���y��U���۝�����o�g
�%-��K7�Jh}�K�J�W}����wWI��ι�K4U�Tr�j�PŷhvF^bn��fU�h���ڬ�:�+kP�.4�j>���G��E��]����3�&����\͖������_W�(���>BB��ݚ��ʧ��(揵�J���K�¡l���+}8��B�o@R��'6[ik�y����5��`j�}'v�&^�ǭ$��t��ݸ�����Jwp���/T6��Nj����Z��:���j�u�v�uz-������`�e��~{z_G�ˮ,���m����U�Y�T�Vd�iה(r'a�	ȟ�f��K^�v}RݸF��!��_<g*"[�/�n���:{�/�ڇ}�z�H߾_{Dz�Of��A=�+7S>�3f����Ѭ+�M���76x��.c�j銹雜����9��ჴ�=��IB���	�H\?��5K5�iXƏg���i�{�i�b@���Mn{�H�Ϩ�ƷSZ��q�p���qp�2��JxG4����E���p�Һz����{&#<�$�v-8F��w�y��k�u�}��C�H�[��h�}Wvμ3
̛�Ո�{6��ܱ�7��W]�h�wʁ�NDK@�ək:��efsF�	BeV�
�S#00.�K�����3RyXV��.f�t���^<$-;�#+P�+������_:��� A����0�uB.o}_W��L��ݝ���a��k�|����s�yuO>9+����=�\��~��K�܉r�Y2|��������e}���:��&y��S���nM]FתN��N?r��cҡ�~���N'�?E�Ss��3d���uG����N�wdv�ǰBK�������X���;l���S��8�W�>�������,���-�Y��z4������yIKܲ�roÎ}a�����VFU�!g��[N�0qǥz���ŭ�}M�q/^�)�M\��h%h��A���b���[=��nW��Vے��ûQ�����co�Z~��9��zʶ]Mc��-N����;������P�;pO�y\���'��z����Y�F��|f�bl�P�zţ{�}{%�"�&71|���t#�&���Uw<ܕ�X�m���\�L-d����62�SV�K�Rc�T�f�T�������Q�yIA�le��,E����'��]s�m!��o�����'������]I�I\Ic�k^z��>0+�U�� ��[x:c����Q'�K��>=Pӱg�uv��i1�ۢ��{���ٳ��ó���eM��⮬}M���Y���_}��%�hEǬ)����b{��.YEHUU>��۞y�g?,�zR��M{8�G���K�*�I�p����yӕ������r�+��qQ������.e�O�&���)-r��Nq�h�Jv�T�OY����Hվ,�\4�� ��O�=�Q)��,�;^��M}kX5��g U�j��5�`n�v�M
sf:��l�Lʕ�kf�,��u���%X�(�&EV���=��uܠ�Y�o}P�Y�5	�Is��%���j�ʤt���\s�AQy�s7!���W坿���	�Mߜ�/df*��ꕃ	Z2�si�N��4!���ڙX/䞿2���r�1�N\7��4�uU�xwD��z�#��^�^�K���}���{������9%o!�i=:7"�S˿jSl璑35l�vt�[����[�m�~�z��%�]i���Q���ie��:��K;%i�Tsj*����M��0�����̳i�(����X�j� k�2�����2r��"�s�]K�nڦ.��n%�,Z�c�5\z��m̹ɼ���v�=a��������������^�����V�)�x�b/0⻟��a�_���ڌ*'��S����� *_���=ݶJ��ا8sҶ]�u�~��$�����;5w���ҕG�id[y^�\���v=�J=�4����=eR��A��${�k��vϸ���#���c�V1��o�x��ћQoFW��w=��/�e�w��IG�|�w+��;��r*�s.�a����p��ZR��'XϚ�L�^�[�˵�Ρ&b�	ȑ�9��1{�SJ��y�|��T9�>�(���K=&e������	�i��q��J�e����j�:������K<z۔��@���[+���NW��=w6{P=Sy�Kܚ�Y?g�T�ԼЖe��<��i7V4��w�?z�*��5����Ҟ�5Y�Y���W�b}�o�蜨j��Ny)�m�4ہ��\�y�D������s�a�,j�ub�J����HGv�h{}	�]�nc�y��tb���wS޿(.���������>�p�I�&�X{zf�u �*ý}C��X�\J���۫�e�we,�� Edx�C�B��^��ӓ�R	�@�hP{ۣZ3�oO>H+��	����ՙ�g4f�jW��yU�w8�٣N���}���XM?U��ϡ��J��x}Rm8S��W�ڧ�&9YK�ϑ��V����~�W���X��^kK4���zI^�;���Fc�����6�A�z�:�`����OE_�%*���(�uj�﫼�f�9���U�^��:C�)Ǯ�b>CSY\�ݏl�)V����f��ڽ�!�7&��a�EY��Vz)�AvA���0Ѣ�ؒ^*h�C���nomֿ_�)�M\���6~/f�Rwa�+-E�'/v-��k���ח}�;t�u��o//Si��櫁�*�Z��9sR1��ZN�ߵ�>h��K�7R�r�Ob��/S�9P�7c�T�)��NT��_�̉������"6�&��S�m���^���^i�o�6���ݢcsD�&��}<�1}Ֆ����o�����_wl�\��P7K�q:h�:��:C/�S�ޣ�8�I�ަ�}u���3w�%��d�J������7*�<�v��zS�y�W�x�ܩ��	�t��I��t�g:�W.��f���t|�	����K��u��	S�"���lW#x����1o][�ȯ~����!rر�E)��6��������P��%P�j.�\�Sp�t�D��U��Q5�&ᕂʛZ1�gL\'NQR�ij z� �9���'S>O�P:}<�NJ����iY�]���now0�q�h�Jqq0ճ_ihz��<���u���?qQ��ViH�G<�)�λ�r�"ӄ[q�~Fr��2&#]����*�\��$�M�����-=��.�/_�}O�#��������d��ri�3�5���� �w]��tO{�>C��J{>��򸃲�i8�dؽ�ՕRaÑu~7�����/��3n}1TM�T�]H�K���:/l��y�3�@�����]�󊟢^Ӎ���?�S�	VuzF���3j�)��+�<��+���>��^�6�9a��Y%7�����dQ�u�{G�,��C�*���9�W/^�z���V���j�v��n;�� X��j�����Tp�|�j%�q��{�r�d�}Gs�>}����|]�b۫b���{��#�--��K]u�veam�5J��*w]�V��{E��ǁC,$�b9g����uw���N�V���-����̩�c1����꯾̛��� ��w���K�U���0�w�<�ߋՎ���c;�l���q,��������������/R��ؓˏ8k׎������Cva�G��jg��O[#�]���^�T=����}�]��	ɍ�$���e�=����~���t��e��T�c��&���^���S��㦯u��]e�Ԑ�X�o|)�>�t�D,�~[0!��"��{��松�7���cؚW��g�m��9
e�}Bڵ�#���rO����O��~Ȏ��k~�ҫ��6�;��y�B7��#�1g=CX*�7J\Q�E���+�5�MF,�����mk[q�5r�6,<���oi�
2�8�Tی���J��=���ۑ-�^ͥ��ƪOl��U�NU�&Lg��N	uC�wlCCv|�z) �E��]�k�mu�uW���-d���5L	�&kM�����i�=�Y|�]�5���i�Vz]B���k+0>HwkY$wh��k��3]��X6�wR���ᘎ��ީY���g.�k�3:�M�g@���PZΠ	n�0��s���A���*u5���f	uǙ|������{�_u6��$�y��Ga�)�U���o�D�b�{	�̲�w$R4{9��"���N�>���k\�9�M��7	ڦtܝ�����՞w�E�	�ï9��+�=L�
b��p8�j�p��S*h��֖��#����i�/(�j�ݬF�A�����ᕭ)���ȱWE�F���R�h\�v�[W������>��eXT����v�����)q�nn.f�cǛ�$)��-f�H�5n���Z'�&����W��蘾ڗYZ�9��ק� �Sޡ�����Xn���G��7Jw���ݐ(�:���P=���Ia`�F��.+ƅs7.��(��
8�wb.D]��p^Sg47�c=�v���Ĳ�L�x���ӎT�;�++*���� =�P��;�����Q�U�α8�e:F	�PyF<���XF�n��WZd�uۚ:pR���Kۨ)���@
�s��f�O��m�=Ϭp�-���%�;��.�l�O^\:��Iw5Au=����Xz�t�_Ko3���O(���v���,{:�3H�u��6�wl�u�T�n��/e�*�%�cc��;�������4VU�Kz3EZ):N�e9͘)
�\�Z�%t�Q�������c76S�Z��?��w�X��
%��\J]��="6�go��wVC��+������gQT7:y*7ǅ����탦pQ42��-�ޣ�屧3v9/��&�6��eJˉ� ��X[']];�����.Yn����e�c�t;v��e��l���X���Vq�Ʀ�ϰ�@��$��nY�1컆��=e���`�H���\�%��a���=�A�TJ��Pu*ƍ���v�I��oo�+�m:��t�%Ӝ5�ipl���D�؎A2l�q*ۚS��,8��)�%�� ^�j�7���"�.�LgE}�]��̓9==ܪ�L����ɠ��$�܍�-����N�s�u�b���1.[�=��:k�K��@\�Go6�s�M�$u� �Ÿ��;���)ttvi�S���>ɓ������o୦էԨ-f<�����`��;-�
\v�JҠ'��e� %u�ӻ=|,K��t�J��t�|��Ƹ�R��r�~U�i��wtU1�9gɻ(U���aJ��I���P���y㌑�yԚ�����v���Z2�W3�9u�t��=�O��D�%�r�4時�$�5�T�{�J����չ��-��k[&�Q�t�d.�J]�p����u3�i�X*;�'s9{\� e�����Ѻ���Sk�G���l)@�O-%�Vg;��^p��\ �h�h�>�M) CӮXRTs�Y�U�[��JpI˕+-3D�!P���$&R�%*X�ʕV�Qx��"�"&��Ҵ�fbd��*�G.'"`e\�E˙�Y�r�n%P��eJ��*�8H��(^r8��B��E���ғ0�J�A��x��x܎'3D�B���1ǃ�I��e�qP�̌�hL��a!�d�ev'�9yJ��T�R�e�#����Y�J��D� ��ig8VK��+K�U�ԒЌ��s�G��!�$	d��I��<�����9�Q��V�L��.\L-%5ΜN�8�p}W�_�>�d�ד,q�6�}ǫq��ܝ�zlDt���v�C6�Ȼ�F쵇�s�	�ޜ	ؚ9��3�K�oz߲�^�T� }�*^{���JR�ٳ�W�S�������y,/�dߜ��=��l!3B��˞ ��U)X|㩙��w���������#^����a�^��ډ��z�܇=/���JCqFn-��Ŕ��!�����cY:��M�,*U�.�"S@�ug���+�;R��F8٤:�N�������p��[�~�ze�^��VT�k�.�@�/f򯤽�Q���
3��S��ݺ*\��(Q3��_��^�l]��L{y������+�-T�0�V�T�¬Ǯˌp�P�~Fی����A�Y�!>fk���m4������ɨ:�\5�nCћQoG��v�?@gאƊQXm:;1_]y�^-���1�|My3PRݴm��xϪ>uJi9.į��M��7`�5	��~���'�ߜ����U���y��o!	�~�2�Ҵ��j #t�����-v�kC*R�v����E�Q0��AZ���x8T��&M�����2� ��E������S��msU�p}����D��)��]���o[�=9�ښ�K�!�.�9k�:fa:�Ο���-RC}�bhs�d�DzB���+�x���\�oC�߽�k�~�-��Q�w��D���f�u�U�Q�-���~+�Kۜœ�emoC�Z���i�<��!<mz���]Wn��	�衸�����A���}9���I���t��5�,Nhޗ��7T��Zp�|ہ�f�<�"c����R�@�Sm�fè)r{`����ߞ{u���M�V�<}����*-�>L��M����!�*J���D�9�e�fꤻ�}+*�{��fs��w���xB��oS�83&��5o���#.�u�~>�u�1TD��}:��ؠ���p�u��O��zMBq�MU�~�e�7}���䱚��4	Ϭ9��EC�F(��
�:u�I@��H#NA��z���x�k��W�d5���r��or%B٫0F}��I�F�[���eUV������6�μF��5��+@�����w���"��~����آ��l�孑ѝd{��hZ�(��Kܐ,E�b��m�*�
Uo6R�ۅ%���vV�]]��N�I[|��I��H,@��jl������Yf�V�_wB��b��n=�:�L��1	�����Yj�L�/2��>X1bY�|%��y�6e��J�嫏�߃yq��O�	^�c=��r�D͚Z�������9�^c���K�j���u���^�~�4�Bt�]��w�MPs�(>�2�}���0��4��:�:�����6���Ӳ���lT����5Y~��˭�y�}� �Df|�nFz��� ��I�-�Ƌ9
/�G�o��`M���f���6B��5��Ҽ��mX���7Kźi�;55�i����^�l�	����5
e�F���9�����J�Iyb�fVw�ͩ�Ϳx��-��I0�q�FBqq-[P_�smY/�6>D߽=@n��$&e��'5�ITէ�n<�7�y�Bu�+�X���_���|k�s/]����|�����l���o��!/t�/:��=�wa�Z��Y���@��1w�J�n�ʮ<�u{J�� 1���i�t���Z��1h��wWG��{�a��ɹ�%ը`2vE�)S�`xS�N��]�(f9�+�_��6F'���2�.W�(q�˗�O�8��wv�G�Z
S`xQʶxt�u`Z.t ��Ƥ��Uh�*�_r��'���*ϊ�E��E�7:v��s�˸]2�����l�N��P*�X�9�Chd�YZ�O�,� ��vd��>����?E��c����x��XqL�G+�NN�����u�}[���;��:z��w���L��ߗ�d͹&�����6��/��F��o�/�J�P��%�F����ީz����k'_���+2p*�|�.�'����q��ûQ��nn�1���N���k^C�6������Q���0}��q%*��**m'o���bvzkk�X���σZ7]�>ݯ������U�yW���;��C��eX�L0yW%{����
skƵ�m�2�%�P��N���V[��n�����揍Ύ�Մ���Ҹf��߰k�}R隂�*��O��6��xf��"��\gP��o��׾+SI|��ش<��W�m�%�}�w�����^6�0հ��RL�l��.xƢ�{��C�j�dt[�ظ��a4U�ثU�E �tUy���ht�ng��]׻A�Mq�h@1���jU��q�{���uf�&Ge=U�OO`x� �q��a����0f�Ǖ�����,�:�=��۹?]AVۚ��N��n������q�~�n�9ᅫrT��=�&�~�Ǆ���1�~��ͪ\�����ۛG��a�,�.���::��d�a{~�>B�xN-ܯ�m��֪Ȗ�/f�X�����,>�W?5��fnB9m7���W��Ty��y���ym|3yy+/�6�Ī@ϰ~��Z�>\��1i�O���<{č]VJ�(�����^��Y�Od�(8�k��Zߩz�~539Y��O���*�W��+���U��wT�j-����
I�g��ŵ��6��E���g�����U�'{�,
V��^,�=^�m�W1)�~��ո�;&�uz/ThueI���gwEn^�_��f.��Ҝ;,����m.�}O@�{P9Α�����P�u���X��%n��H�'=)4��%��S�P�~����`�x���&v�T��ڽ�qoLy��5�HZ����S�6���<}
�߮'�:�Q�#Ε�{�/EI�t�p�/γ�rqV�or%uW��z q����%b�Es��u�v�5���dvfW�N�3� ��A�>���pGQ�l��K8��N�\-�թ�]��-+�]:�h���]e��G�<�����/6�o�q���*�h
`�������v#������$H���Y�9<��Ʒ!�ͷ���t��=���U!�گ��cT��:������k�jpڸ��B^�F�����R���s���EӇzV�JKџy�c4L<{#�ϭ4��7����~�r���?������P�j��^�ԏ=C���a����eܡ�b��j�(+j�;eE��h��f�4;f�S��r4��鿊󚗹5����ǽO"m^
���;�T�E����6��z��pU��k=��g�-�cZvPԊ�hm��ݩ�����(]⚴���ծr��:bVi�7^�oN�e�����ެ���?,�<~{/q8e}�Zs�y�mқ�^�ž%���Y���*�o?U����r����H��39����~�	Z/`���9f����Z)L^ݭ�x��bޠ�t]�^�lY�VP�f^�Sd��ߜgʯ��QvR:us�o}�|j�۾L*@e��' �ce�N��:k���s��s]oT�m]	����Gw^5�Qs����c3*8�]ޮ�;�owv�\�a�;(�>��Se�]^���V#S�l�9V�maſd���u�<k�'�KF��8�GH~���ݥ{���8�w0٠M[������]R+ڷ��1]�ߧ��u��m�D��\'�X�N�EXݨ*�*�/l�x������X�6B��>±����"��&�ۭ~�S{I��u�l����>m��N�Zy�P�r�ěڙ�j�[���C�o//6�lB��p=ez�z��|ǣږ8�#X8>��T��N�UG>;�����^�(�{�M=w�\�{(�\L�}+��j�4Ow���o��w*�9��B�������_�����Ѯ����g+�T�Br_}9Ц*��-����F7ۂ�V�)K���n��@k�XSI�#o[cͳ�{���}>f�zf�s�\�S�X��U�y��t/�5�j�z��r&+�<�r^O�#������&�crxd��U⢙_�$�,ݹP��-�����lC�"�K�ɸӌL(��3n^�n���v+T<�P�����f��X�{FE�7ve�N$5��`�6�<.R/)�(�ǌ�d৷�ι%t3��ZV��ޱ�%|��!+.�]wR�%NY��I,z�c����^y��s�AT�=/ޕ��7K�Kji$Æ��#q)�ĵl�11�����Yő�Ek�*�9�ˉO'�k�p���N��q�p���<�V�gb���9�4+�8�{��{hͬ�c�}��V���o�N�4�@U+t��V��	��4ӟ'g�����U�M�o��֩�q�l�½��|���iܘr�&����:�W���v�eAퟆb��ʝ���8�=O#oמd�%8hC��ۙ�?&��l=ܨ�y�������U��-:G|�{����>c�b=�U��F���{�K��������������&���N{�{���^���Kڌ*&7�9M�q/^�{G<1w��Q�2��n����\ħ����|��������U�[��z�sd��c|$���{����b�~�G��]�����z��SQ�<=f�֪6�X���0E�F�a�XR�����[#�wFT��M?�9%��QK/o����XO�}v���x�f.�N,V\0TC�e-�v�8t���'97Q��%��$j�]a;D���5��"k���Zb�o��\��&���*|��wt9U��,�o��N�D�m������Ϸk�ts>�e�"�&71I���iuiL���o��ˬ�u<�xֽ�lar����}�G�(vR�o���IV�<�UJCz/���;����z��n��-	��}H[�Ѳ��ݖ�Af�o�DLS�8d�������Tji\2�;��B�~�i�?{�&)g�(_�>�i�]J��g����^����U%�i���n<�Vײ[7l�Z�Ide��s+B����H�R�e��֝_Z���w%�Oj@M��N�� �ƒ�����X)��Oo�������w2�c��X"���%���l<D�O��W^�UnhfϐE%��0<��b�y�dkUp�)Ý�p�=�le�ڴ�Ng��S������XK�ZZ=,]�k��˿Wj~���g+[K�a�����?g�O�o��bf�D��{L$��;o��5֕h��k���6LJ=�&���νg��{{,��!��}���Y�^�;�x*Y7��<��x���z]t��\)ӽ�x�E��fu�K.sȟs�ʱz��2�s��HGKi�p���r�X�'F󮻸�� "��O,>yȞ7�>�^��v��7��"�pzz�����NZ��=ͶԌp�%Ee[kr\�+<n��}�.v��q��0��լ��/Sn]�t�T�Q;Km�-��oʢ1���|V��C���|<v�44y�VO����qE��ezRK�"Z~�S���+k@�>���;����Ag��5; ���1��.N�޹p�c�����n�zʯ�h
O�s(����M�~�Y�`����W�d����k^��?�)1�.�.^Fk1.�O���\(t����Ϡ�=�?��Y?W�5-�F���`�xϼ�r]�5"/3�Bm	�����9 ����wϟ���1���=�_�*a�~�K�]]Gr_5��ښ�S%V�[B<B{5+ِ����<�ǂ�������eದ�ƿ0� <q��c��*�e�4q�;~���i���;Ay�ؕ��N���0��Y.-{	��������KB���<�^��Zanf^<����_q�Rc�)��_U��;D��X6�-�
鯛:BKE���c5���V��������w�9-ݥN�Ր���‡xJb��0��T�˫�&�lp�#�0vi6��˱�����T[��5l '��,*%���	<+��S���\�gsx��b�8lqv�h���Rv�cnU�g��q:���G\5y��[utxF�wMD����}gMnkd����kK�7���sq>��ݾ饽?x�T�1i�tkC��[H݃����E���0;J���A��n0������7��x�e#��{W��|�B�1�1'~�H.7�;��:�(�wonУz�����c�"\-K�:[�i�9��)������f^^��#�W�4@0V;�c��8��[T׀��rm()��޽�m;@��z]�g��'J|�$˧{���65E���2����&��_E�G?��I:Ke����XXUb�z�/���&��E48�ĻR{�>Y[8L�u&����Osw4W�Pw:���q�w&�@V�&�s>��C�t\%ܾwV'��)M��vE,�ʆ**孬4�b���
����lǯlI5s�2���4��>,]��g0':m��uҬ+�;00�|Q���6����E�:4�؇��i*��
;t&y�Crm�T����^-�CV9u�ji�3�S=���t���G(\Hr�gY�oZ��+b4���.ү5as���r�6u��O�k������i����Y��Ұ���zP]��'5ϲ.)q�q����i�X�̄��ť@�r'�b��lD���ۺ�6Cs��u��^ڹu�i�7]5�\Ohs���1�5��-h��v��@LWp4��{ȓ҃�v�%���C)1�Q�;��>��`���H�,�i��k�dݙL3|ngG�|a)�n9��ˤѹ�nT���Qr�	�4-��V��0|�cΫo,iE��K\6��ZT:�aV+4����a��Yz�@@�k�$o�2�{Ӯe�Tχ][xZ.�<G{D4;F���-ueuj�Pf
c3�P���t�^v�͗%�ekY9$J�n��2폺v��<�7Y{��i��/s7AN��]oX\�`=�9W���t".o��Pgmm:�ۆ�)��4�+g����_;�+���l����5im�
��DS�#���|��y9��y��|{;Zlر/�-�Y�"z��i�,cN���$��AV�fq�����;S`�wsks��2LS{���/0��t�FN�\�P;�ʝd=���[ ��;�	���Όj�5��9�;�+�p��B���l�t_U�|&�x��X9f��	i���
ېL탺D�8T*�9Va�(r���&���_�������nG�*�J�%M-���M���""��*
aEhu���I#�iWn2�	�C��G\��r79q��Q���PxR��w���qDN)Js�����(�"q��E�hgi��$P$Ut31L�*T#"����A�^D���Vg
���]�p���$s������RM:��M2�I\��ċ�I	�ia\���"�d�I�e� /(�4�e��BP5��J̮&fA-l�1$���Ҩ��Ĝ�ArR+U-!9vP�t��-H�\������Ur�˜J!B�2�fj�R�J*���e]4���		r279�93*��"�����EfD�����UL�DVe�����˒�.Y$��a$Q�B��D�
��3�r�ʓ*�c����B ��D(��UQHT%�\0J�[��J� (��%�L,Jx�w/�^Ց�	LdL�|�Y�]�v����LR�Y�I�̷B�:]�tՕl������ٳtu����+����+H�Kjk��7w�O�qq0ճ_M�߭��w��v��LAr)�ά%#��Y���4�OfJ�ޮ�{��*��Vg�;�A�f�ם*ץ���.����^�䶳�̾H��3Ю�xg�����r��r���p�9�;�'U�}g�Fc���`�N�q-�^	=~0u����u7��s���#�gu��γw�>���nBz�]B/O^W*��ƟOhԠ��e��y��)�����X�w0���Y��W�p�^�K/�rD�&�V��~.7�TiM�ϥ�z��Ʋv�n�r��7�O��~EA̴�'#}Q�������[�m�s�ڦ��5��+@ڻ��L���O]���r	����%��e-�n��7��cz��
sUy[������'iU{$8�nY3��U}%"7_����z�~�Y�6�̀�NF�]E<[�0�љ�cn��q�(���߽���ζ�ފ��
�?/H�Ȥ�	��f�v��9�z�'��}g�V �k{���2��gWv[2,������vX�ձ��S\�ej�kRI�۝��ѤĒ����)��,�<\K2u���q)�gS�7�N���C�_j��%U'W���)n��O�
��̟4FhHd�<�lf��r�]#�N��^H!��!������KDy�e���w��{������_r�j����}隂�*����z5���nf:��Z�o�HmO���b���֔2�;gL\'NT)�:ёn.	Yt�[���5.߲j"ud�~�7J�����L;��g�K�R�˚W�}��U5�n//S1"�P�L���[��y��w�N��y�ԛ�W
/*���U'�]�m�D�z�?c9���]~ɝw��,T�hT^�ey�֫R�d������ǵ=Dn�]̪��Ip�Y������jk}��5��v�B�RN��Mǝ��Y���S��@̣�#18��h�7+8j
��%���~�ٝQpS�l����G�뵓���<���Ƅ�^O�s�X{:�Y��ջn�%(AhS�+�}�C��rҹ4��82�}gi��Y��]u�gB�d��}��ݾ-�ZSu��y�� b�V��1�u������e�ҝXmp���Sn�%�\EF�f�P��բ�V�׶�G��=s�˘l&������}Q<�<BWC�>����OQ���Y��9���'�ߚx��|�c�-����b��"���*�d��¢w�2��/^���sY�_pX	�Cn�k�;k�{�k�@�>�@�);h	�x��_H_��V����R��|'����}Y���y��gKds�Q�5C���{�#��]/h�Z��fqì�^�Q[aVcN����j�Ü���!�]��9��t=ܭR�ħB�E��iR���$N�Y�'�=��zZ�Gޏ)ՙB6����@!����������u���8�L?{q���Ҷo���{�P�S�s_!fH��f-8�{��bo����#�d�N���Tji\2�;��B��荋$+��e�U��	�;G����i~���5��d�~��*��5��cwf)řq��	�5�Xᛍt�AV�h�Jy|�?���~\�?.W˖��</����gm���՘��,o��9 ~E��חnd}�Ρ��i�+43@�j��{��d����B�N�Ʈ����\�W�����A�M��,��/�ּ����!*���粻B����쏋��Ƨb���V�ޮ�E>S����=k���G%��
n1�B3�q�1�yt��<�ݺ]~V��բ=R�۱�F�sf���W�����j-���ϗ�E$�E���{�,�k�Ã&�i����mo����j��#ާǇ�<{	�M���
�����ikEbjA��p��=ȭ/R��@8ۮ�O���&��c��Y�G�"^��\�o���fC�Z�C�n.�K���(w�����������n�r3WB~��Y;t��Y'>���{ ��>�*�꧘y�sge����kc��!��&jy����]�2�>��Y�8tb�a^��n |ח-���ʪ�x��2������jsi{rUց��P�E�3��ZE�ݛ���e�3m_�r�17��y�Yx�z�m?#m���K@_IJջI�V-H�C�f�����PRy5�n=��eBt�z[�N��``��݆����#�,���R�9�ft�5,̑��f��JSi�X�j�;��'Ӹp�.���;b��݄��gN�\��k�zC҅�Û��u-#aF�����p���P�I�����H�����㹺���1^Dy_>�W%�"�bK���̑�TV'��c��/��������p,��͚)n�#o|߰y�f|�bצ�xl�4�VMF�*�ۓ��D<{4#ճ���;VLK��Ú3�zzWk
�x5{�{ί�ᐦJ��>�Of�{2�&�&���J��[Jh�Q���sI�����EV�,�Z�c�[7l��I�j�30=����|���2ԯ�3`��ha���������ݹ�c�d��7~��\U���2�M<jOn�p�w�A��-z<4�����·�+�`����c<�痙��,�է������}����6�f��7�r��9ϺD���j��bֺź��:V��T�zi���I�:�%z��6���#S�6~9Uip!*�닫�)г�&�f���7�7��sg@W���k�)��ڼ�3݇2Q���yY���7�s�bА���m���y,�k:�p� �@NV.�%��-u�9�$A�/��u�h��������A�.��e�"#(n�`�j_=�ŕqj��i���g`a��7��w�Lt[AQ���_\WI|�������x�t���}U0q���.'ڵŔ�ܗy��[۟(��6�|}�4�6�}\J�S�uu6�ěU��}�����[���ۇZ�����L���f��!��x���{�L�V�R�n���n6��$�]�܇T"���=�MM�e���X1ꯤ�F��B�#u�4�nj��tn\?���6�~9_5M���UB�P�PJ&>*�:�u�	����Jy��RۘgU@z5�^q��d�d�˥�'�t�'��k�
7�$�ƏH�=D)�W4��f��a�qĺf���d-��G� �~{�i���.�丟f�=�ڵ������9����˜����e�=��c�2h�-{�j^��bs��T%�4�a�q�~F��C���k co�ݶ&ЯS���rm��摬�,ߗ%<u�b�+4aQs��"_��i�妣#�:��F��]�onq:�2Gm�&��ܭ�e��G�.�й&'���C�)����3.T�t�����!
���ƴ=����`WC�X+��b�N��t�Ƀr�ġ��۳E���C#E��NGS}
���]}.�FC[Ư;o�����n��^��
<��U��Uҭ��澴{s�^M�G7����Z�t�n�&�s7!��Fܣ�N}Q��S�7,�mZ\���V��
��2�	��^�wF�ڜCN�Iǝ�9go��0�ܻ]2����1�QFH6}�x;+\�g����ZN�ʌpn���Ψ�)�\7/ګ�-�䱟y�kh�R��7�D��X��c�����%��F8�Z4�8PSOr3�3�yȻ�jz^Y�=Z$����vb/�9�}�s�宩uv���ug�o�vs廸�R�n�|[�E����Q��'֧r�ke��2����sBMC�{�b@ՙ��𶱀u��6�ۖ���[V��q�C����v��ӧ�/&Sw�K>������9�;����5��+�s0����}�`��F\�V�^bJ�\���W�->���yf�軏��SћQm�.R�e��B�jD훝�l1�`��Zq]u1�	Wz]sfj��p��;�ւ�^��K;�Y~���72��dm�e��`�2�(w�E�$'&b��r���̓R�yK/EC����v���r9S��r�>^x}|^Xx~�]ٮ4�o;�zԱDM��Vu�yotmr
��t�^���ط���b��[�
xϪS�5��f�=��ۋd�i�°)���>����2cWl�^��M$�����F?����x^�/��PǊ�\�'�j�=�B��<�˲����O?��ʭ��R\5�,9N�=R�0'�y���L'lL��=7T{-?�zӾ�V�x;��p�7˻�K\�ƷSoX-�Š��j�V)�@�����+��l��2g��|�L�}�4�7Um��fځ��Qqu�|<�
٨��Xk3�9s��ᑔ��̩X2��է�9�ew�yxx9�~�%����h��C}^��5��a����B�)�k��_a��39_w�����Ƭ�+)�h��e�t�E�ۆ�'��肮Fj���uK�5�Q����{}Q�<��8f?����%�{���si{�C��2	�ډs�C�}�4��L[����V�������wn;��hYB��ey�)����V.]��4��=v���)�[-m؝[-N�wj�\����4���PO�pom�Ӧ���ὢ�ac��h�aZ�0�;{7\�&c����i�sh�S�97p���C�M�8I�7��������[۟(�B�O����yB���JVuz�(⸍�z�✦ߗ�-?#{�^ܕu�l�}v`a���+��~밵z���x�������c������v=e^�~���ͧ��^H�1�}z(-dn�J��\5�m״^���u��Ɔ�V].w�3����XX}Q�k��������d�^l��-ی5��M��ԉ�.�=��F%q��Z��͓�>ܘ�`����[9198�U_��n�3G�2Vh�[{﴿B��;<]rG�j�d�Mv]�MT|uw�|̰`��h���t/��2��5�oC�hT'L�|���/H$�}��J��2J���c<���ڔ�5�#��!���s��s��^�5ǩ������$s��W,SO=���\7��w��j{.�����d��N�6�~ٌd�ˤѥO�9Zz�fK�����I�PP�IC��:=:pf��k'�CS�]c��H>��m�o��0H�w-)F�>�Ts!�]�;s:��s@��.�9;^�v�#���ܝ��r�����|�c�y��Z2v�X��O� M
�w���z��Ss���^m_���\{e���r�7`TY-"�|��D�^+se�3}�����	k�>��E�6}=�c|O�|��A����y���@�*Sz�')6u���ytf��'=�~q[�4_�r��7��Eˍ�L����J�u��_m��SMV���޸�9�#�+��;����������c�e�B�	�	�)mq��x�u5�K��{�Nc.i�����:���N�wk�A���0���H�Y�R��X����S;���˱�
>S-�[��<]���p��uw��Hr�5�������+�o޻:<V�9�G��d�FGa����S)��	����0�wU��'��=�ֱ�1R1=��)a��.��aS��tʞ7�K�1�)� �v*e�eDԥ}ǣU:�U���b<���;Ϩ��㼪G���r��Il���:70.Kf��/Nۢ���gmw�]�y�k+8O	ݮ���������>��@.U�w�D�p��&@����i�ϫ������`+C�}�,�ݳ0U�B��:�ܼ�fu\�������!�E�[k��]}9��]��7�X��F�Ew N�E\z������t�J ��Y���lϛc���>���Z�������mh��*��{�)cb$�|��%=o25]�ݫ[2�����RlN�Ԅ.�:�ܣ�ׇ{pZ�v��A�����έ�p��묽��l=R��ы�')[pT�.�C��V�J�V�
�V�:�7v��3]\(�Ԃ6�n���HW��f��Mk��ɝuv���3eYB�+l�l��ڡ3�c���s-ᓂ���5Z�;�d�
u6nT��l��g"v�-譻�r�.�ؗe����o��ܮ��)$��A�3{��bM�ԛ�na9 �r���\��I�Ah�De�}��Sz�/qG]��e�γ��,
2jW�(~��t9��X�wu!�c�hۢ3�f�Vk��X�����Z1F&s� =֕�)�+W �t4�-4�.�!7�t�zMu��V�e����V[x�SbCt�+W��o��i��5.$�_^�^+�}�R��7�V����w�c9�&�,�ݗ�����!\:�p�To-���1�V��GqC��v�eN�Tm�o:�F��s�D�h+����yS�����:���8��-�<4w�Nk��,o���Ҳ0�w�)N�1��S_)A�	�kvnf�hg)��ѧN��g.�p��.�T��(N���WLF$�A��r�m���V]��iQu��
��N�D����g5:��#Xź���vo@�/i\un��|�v��=���@s`��e��\]5�a["T�˨�@n���.�z�j>�gr��j���fuMX�|�V��F,��-	az
�t^8�6��\x��h�1�����)RH�Ƕ)�#��{4n�K{�3� �F�-�Y��J$6��s��-�\R���2�.O/�%�v��wZ�|-�Z}J���\c77T]m��!¤�M�O�n�
j�o���X��M���y.]����u�hZ�`�W��ϏL�D�	��1�)���r�2���:��'<����,蒦��}+��{�)�ܕt3�;ھ��պ��&�jk��xg���t6z���fm�,pݜnk����ѫ�M�Ǔ���W0�����V�{w�!B^�\���_-v5V�o-�NgN���®.d �bV�]]��`L����z��u�p,��v�FRT���hm����G��r����ζp�n��[�
�eoeJ���]k��>�*[Z� �l����`���r�?ĕr�
���辮�.=��Agd��-amU���/mQ��ʰ;��s���y��α�ku�ӈ� ����
݂^�*nt�ޚ�5&n�7��T���y���u�Pn5e��EL��Kv:�+Wr�k ��5��4��#�Z{y�.�cx�Pzb`���o���7y�� �h��s{��p�> 22uw;]�(w7��kEQ���P��H�Ȯ���s�C�&	���Y�RgQ
��,���r����(���&r22��,@�D;���Q�&��Y�
�!DW4J���2�je�RuTR��24�YDZaie�1U4!T"�ʳ���6hj����U��%�"�QR�S
%��b�I�ZRG$�$��R�)�'�Yr�D\.I#T\���3D�YӰ��YZ"I�b RML

iͥ��HEVdf'ERDҔ��(���8R�Vhj�jVE"&�P�Mj�2�6V�Y)��,���E�.\�0�*���Qk2�欃��Zd�$���9�d�ֆJ���9\�
+�`nRqQ$�A;B�l(���
,���X�*BaQfT�#�Ua���p�4�<yŚ�+��TW:T��Hp��Q�!��L�9sU��kM�A�DU'1 ��FT�RaKJr!˲��d�-:fF�����f�%�>Uy�k�*5��U�bs�'���.�2r�82�5�3��{-�Zu����*k���
t!ˍ���+�'9��]
iR��9�Q�
=��&�~�S5�kGd���=����f�5��&��0��H��&7:���^�C�ڜ�ᅱ�
~���>��lbې�W�����g�}�>d��Q�����jݸ5�<6�Nn�N�B���x�0�T	�����9T�:��\�-�wB�\O`��7�t�]�¿_v����%�8�����6���k�n�@N�l��w�U�CYO9�G�uR8�Pe����\Н�����xoZOp23���K�ʰl=7Ӂ��ɳH�=g�Y�}��ޞ����y*��m,�&��|3���r��4=Զ&��Hm���7|���A�����ep��>����j��t����k�%g��+C,J�zc������x+�Nq�8�H>�_�?�̣%<!�# ��GB�}��*v������������aL�pK��s�k��U�a{��7Vb�g��S�r_'b���>W�N������!��P��񿫤^��^v�
�v@�uϥx.^�f��.t��^ɇ��'B��G}ݎ�
>'2���r7�rXil�nPiGFPgTBǫ;�M�/w��Q�.�	%:�u2I����
�g%��{���[����뤑�ܺTRNa��w��z��\����(IqI��:ף'.������]f�iVT�!����6�`Ì�����TC:������NקA���������EP�>O�͌���]|Y^�-���Y(��IhѕP��3��3�PPu*9>�-�k�ʔAW`h�u���NW:��h<9%��%lL���P��ncW�8�,�N+3��`��:=���Py�����;g�>���y\=Ϻk�{>8%��p@N���}���ͺ^���e�D���"�S+�r:��[�<1�u�y�Tgu����#}�<PiC�K&W������w��RBn�2�� +��<�^�����]t_t�'9�	��^�R{.}�ޣ}�6��N�,����B$:�Q%���0�F-�\'��ΞXO?7�z���qxtp`��(�xvuhm�W�uU�7�2KD� ���qE�j�Cx��
�*D�z��s��k]���%�:�,�:����_>��hN�t��Od�75
vӅAN�h����M�н+Y<��0����:�ݪF�9\L�����f�z��x�sc���nx+8:5!�(�W�ٶ����͎��,��x����Ϊ�<���4=Ӣ��!�1f	��'��ƨ�$�n�2?~uU�Oܞ�f6dc��2�rkg̈�������\���bS�z�tZ�׻:���L_��;��!�o��XW��:�h+8�r��т�Kk�r��ԣ�#��V����ν�h:�w;rup�9��ܙ��V6�<�iQ�y�&ep���qԧYq@-�Kg#�*�0�Uv�y��~�2�;n+H�Y��dJ�[p�v{f*����z`�����Kˬ�[.���D����Ķ�n�t��!��3t�.�����o�=�wbq_>���ɻ����y#Z�L�o�؈��r�Ǔ��U�f�񲔃��H螮����B��AG�ר���zKM��;P�+����������럯5N�<=0i��˩39�*_Tg�n1{�z��%l�
�L�p�@� �V3�K����q���&�Jz<g�W��B��O#﷧��]�:�ϑ�{+ƙȵ$�{n� ,�q�w�ФK�3�êU!2y9ط4ߟg��c3�#����v�9�:�Fb짹��H�u�,��C	>�@zH�.[2J���A�}~�?W2�����γӕq˪������9����[S����uc`Oź��3`����-�C:71G��Sn��n��������G�x�G�:�ث}U=, 9��#L��D����#l�{z��g�x�~��$XA���9Y�?N#�� �w9˲��F�c!��e�]�]�%̃Ug^�2Xō\���]��ƢWD�P�E��n�a�ı7�S������=�5��[�V��2��)���E��ˤ�u�#]B�m���'ڳ�Lk+����s�)�º�k���}g��s�7��q'��ͺ���©-H l>�+:9�H5����F.ܬ��Y�Zj:�M_Q�<��8�%���_>��E�/+�ڙ!���w�C(���˼��8OM���W:ʠ�N�Lmn�R"���5�<"��Pa_P�7�1dOT�:.��l��Ss�O;��~!	�t��.�eW�v�W�c�]м}A��>�t/���]~ӛJ���ԗcW�ø4!�Q��#��[#h.M��=~��Ä)׫c�^%�sx��A�t7���2sYR=w�L�uX���3��z�A-��h�����5�GY,���FwNYڮ�_��Ts"�W�9�Wi/���{�\%g�۹��'(�]Z��K��Tq`��m�q~��ѫ>K��cht_%�.�����u4������weG�#k�k��tc{S�s���]3y�{5�_��߱�-���6��$5>�������}}�O]F{_^��~�G�2�n(Zϕ� ���N=M���:2�t𸩖��9����~.�
��z�VDwWqYt�-�sv$k�`�#�.LE�{C�gT�-Eh�[��Ш<�bb�%�ߔ��e���N�vV,6y��N��mm({��C�e9�W=[J.">����n)1on�jx+��Z�rWS�\�7X7���*J޼]�u>�q��c�ة���P#�;��}F�Έ>�Q.��u�\ÿј�羺G,�J�0Ѩ�*��R>��	�<�=�av��>\k<�ȿu������eA�06���-9^�ʖXD��E��{���r3��H�wy�Jh��bT�k�����xoI��Z1�k������r[� ���:[>k8�F麑���r��Vs�=Y��o�]i������:��r==4��R��_h1�W�1�󜎛�n.O���5@��}���zk�[ZD���dt���tͲk��M�]U�b�R:x�20��pD�����h�	w�@S�;�4'��̀x,[R�j�1�t�ǉ�K_q��[w�Tϰ�׶o���/��V�_�1�_D�/�r4��A��<�1������z�ؼ�~�{�ʽ��rv��&�~b���P:��(y;uܿ��j�CYO9�B��I�Pۮ����E��n@��}|��fhz�z=p�^38!F�`��l�����wַ�{���V+�P�㋪����ˏb]v�y��n3����}t6�Pɛ�TADa�<�{ފ~�=���B��%�@^M�ք=#�⬩D�[��kL��Gk����m��y2��TC������"���]p����k�i�j�W[�Ғ�w	͖W4H96�޶�p<�I"oH}˷������%��v�Rr��>��a�/sB��"�]��+k7�v��{1��̚-��6�f�7�?U��	�]dn�qq��+#�^
�Ӝk�?��݊��
�c���c���� ��������:x�������cRy%��9�\uz9Z����V[Α�w�N]�V�:N�|fW�|�Y5�qN@�z�����\�s��E�b0⦚�щ"�]��=��~�G"����xAه��HΘ��iGFS:�4y��՜��"|�E���2On������8ju�B�?]�r�(Ԗ�*a�<��E�L��tymą��Nt���ڌ����#OU��IE�{�;��9���փ���]Ô	*�g@��1�[�;���v�=��nD�������*�{����u��4�s�|g�y@��,�8 'y�Q���N�5�)�@��hNbI��׎�*�[�<3�����ܤ����>��a�e�+t2�JZg�6�����@����;+����/u���팎��ᾎ�ZO����]Mdf��d�g:&�C�wQ�ϡ�	@]2.K��a��[����l�>��밢�n��+yg��J����N�v�S���e������66��3%03�L�ur�)=24t���+��[[Z�}2�q��m��MvB;�a���T�m�ۤ����J�6t�5�y�8�K���<��ܛݙY�Λq/�r��6�>��-��K�3����Z�VvE\:���%�cny#�Zr7���;x=��~���Fr�E��t{��HχW 7�!��*e�7.��b�S'���f�D��
A]�Y��g����_]�|,�(=�C3*��b��ɸ��{���"��X:\�����Ѱ\���^�dUu��>��[[
��+����XG��]&�Ӡ��>����a�[�~����cq���3��Np�Hܯ��Jy���d�r:��x��]���N{��ʾ����կތݾ�9P⯡���z�
�	��3Al�ayu�[.��"���L�� �!ݕuǠs|F�fz_���l���������^Ch9�Ƶn��뎖pv��<:�1-��M�����q�����3�v�dP}�����زj���=3��k�Nbq�w��Ό����x;���f��3�7M�ޠ����9�E��$�XD]�m7#oT�k��|��ȯ��gK��,3�F=S����=�'�y��ۜei5Z������5t��Z\m�v�I|�J�V]m9%t���ʼ]�TXL���a��=����v�pA_t�L�z�h��d���qd���WMޮg�w�JJ�ٵ����D��m,��ٜ�J���Y�(WG}�&#��vWV�[�-n�o&W<=G����U� o��|���O'9nh9�>��u1�uv��vזkX�%C�v/a���~0�<�e�I�|��"�KfIAv�Ǟ/�o��>���V�Ɓ���@��U=���9\Q���V��k��;���� '_��%��;+��0�j���w��dyt\�����1�C��G}��CI�t��US��T��2 �5�#L��@�zz�)�ж�go#~����m�B�&Nk3�����g�{�����긊y{��Ԕ�.!T�� 4�ٮ4���uo���o��R}�t�qi�{�j����<�㇧�Og��P���/+��������:Bݍ]@�������^���k��!�6��Ŷ�̛����&23�gTuC�n�Ӿ��>���@�K)ɬ���{<��2�9�k�^��ΪQ�鍙�2���y�b�M��`3+�"W}�����{H��"�m��arl�:�_���?W�cp{SG�z�^�3r~����37�V��>�k���_(%�>��@�����5�:�e�F�|�Y�^WJ��]�#1C�5	Q܍��\���t�Q��Z�y��g'�*77V�v��U�K:a��T��a���#	̼
�F�C*\����`�\7�E�0�ei�S��
��^`G��8�'|��Q(��R�3��D.,-`˻���*|�,�EvI��u��I=%��^�W	Y۹�p���>�]Z'N��=�.\iӗK�$W�eC�=ٺ�T7��1~%�g�O��(w��Y�#�w���wi�@{g����Sf��|L�*��/t��3=c8L�w*���]!)���G�����6w���۟>�f�������E^-�J��ሼ��~!<j�pʀgO��F��e_��+�w TB�=|+>���+�#����=�N���􊾐���#�����*��r5U1u2��<�yty{��{R(��#�+ڼ�d=�}�@-�����\���2���Itf6�yT;���n�P\E�]�-Nm��H�^�z��.�1ĝT��I�;��C��S#;��>9%�9 '5tn`K�����L�sY�6e���3�#�E�Bwk0�����t�r��L9�Ze�%�DF�˥���D/V6���Ȟ:z�P>�<+ ��ŵ���/��>��/M�7K����)`Ì	]�S4��=�H��s�_)�qNw��p[�nC����c:yY�3�O��+�xӵu#��<?+
c�ȵ�KX�sc�P���	��v�m�95�6�n�+9�w<��~�پA��5;�e[t6�,3�J�	_�W,t1�>��m͙�)f�tU0�ʵ�M��	�߅=cT��q76���
�WF*s��2G:��������?��~���Ҝ��|�������[���ϻ�����T��ܪQ%*������28=z\O�;ľ�Ҁ��Q`>��
9���FI�4n�S��>Gx�_45�:+�wO*�����N��M�����H׻�F�wWDY�i���t#:h���Fنj5��6VB�s���\oEރ]tU�β��ˇ���9��P':�������L�v#
>��^2�d+��\��8b팛�G��:�f��(?U�ӆy�cw��9�����Qߧ8�V�:y"|��S���e�������ˎaO�qAt�>�Kk;r�T�@Ϣ_^���:�
>q���eR�p�g���{����\}��ɽ:�|�Y5�t�W�`L/;@�<���zaw�l{�×ÌZ�nO�������E��aQD�XF��f���rXh-���iGF:��`�8�6���_o�M���\��ÞWZ��6?]�r�(Ԗ�U��"n~KbX�:�ey���\�y3�t�QX����}C�NEs���h8�r^Ô	*�t8�����ߦ�t�y�;�ZV���^2ٺx%ˁ�6c�4��F��oi������Ry��Μ�q���k-�b�ͭ�o%�4�xew��S�����.�SH�`n5K5VU��]D���k�߱�+�ks18Obn������m&�]��[�7�1��}{��*�����Qwe3j�4]@74.�_lݠ��y�81�M������N
��{P��*N�n�5��k����\S��u+Sw�+^��k@�X�Ml����Y�x�qӡ�W�xU�L��[���WHt���P�z��T�`^���8�W���z��<X�+X+�,wm>I�A�h��G�#���;p'Xtv����:��!��&�]�WC�P�%VΑ��5z�:�t��1�^�_2����%����(ۨ�^pBd�����5%��������Xue�5�]���u���gV��v��"�������g=��>�㈞u��:#�Ī�����[��~	��e�:R���,�9Z�1T#MBdOuNd����8�%��6f��Yh\����՝|΁���8Î$�	Y��R*t��d �noJ��;��,��~�mM܂�c;-��d��D'l���JDR�,U��tn��N֍�}��۠[TL鼻7�J���U���9�a��#�ce.�5�|�6�Iӝ&��1Z�FЛ�2�6N��qN��dJڻ���}H�}��׭�`���I6�����r�(��pPFr�b���Ӏ�ˉc�7˳��GpZY/E��/J{	�bVP���!��S���s]�F�ros�j�L���h���w	�^ꔡ��
�SJm5F�c�uդ�'fĕ1�'o��J�j��)�v�,�+kHUdJ'Z��%��ӆ��;�E�)�m�A�:�S� 	�ӑ (�7w*k�΂�h�(Ԯ�������p�Fc}F��%^-�BK	�D��[Ğ�[|eî�u��2���aL 鞠���j>p#ٱ5It�ٷ��ۑs���P��ݷ}qj��ڲn�*r�V���:��b^b�Nt������<�r>���9�E��7snl|�{���ݱ�%UD��K������p�9�|2��s��j�\]�@�8��I*����Vx��F�n�vw���2����;a˫V&����%+����y��j��H�<���ە�^��:̪$Z��k��6�t��'�U�w9K��fp����͌����ӌs��:W���C�}:��t �J9����IM��:l�ȕ[��u��@�m�}�Rgp�R�d��3.-u�'���wZ&T]v���`�d](�
�S��;{�lM�ƃ�z�0��rmq�;2��t�DV��K�z����g��(����tG��g)��.���W�*��#��kU_8���T����ť�Ö�^��ݧ���M���=�_nN[ 8�~�����(�KK�Z�K�QsRV�R��~drdEx��a�CP�,����"j�.Qr*9S��VRp�G
��+2��\V��T&DA�J�(ȲЈ�
�(�2�.FaS�*���g�-qҊ�vQTj�Ȫ���G�
�����+�!H�9EQ�r9T�*4QNp�\�s�QY�YTI��,:Uˆ�D*�\C�"
d�@�H�q�"+ȑUQ��PI�DH��UQGr��#��V�.Eʬ���3R�T�%�+�D�ʢNң�AEtR�Es�UQ�ND��*�����Y!l""e]Y�gV�.ʢ��Ru��&"9�* �9G
�����Y�6E�UTQQ\.D�UEm�s��\ɢt*��E��p�*.p�"���J�Ү:�󧟓W���r����{�'
m��{�v	�8fu��:k0�wʞG�Ȩ��+V����R0��|^˘7�
z��X�dA���uȠ�q�3�X{��9�8�9���������ǰl��q!�3�M�C�.з]�y�P�|�Da@�<�bIO�a�
-�7�����d�r��u�,�4h3~�d'Y1��My׌.*t�( .�2���@W)��X��Os�3���2���.p�\��R|���]XO}��&���
���͢ 5_	@]2.K��a��[��^>��je���,)��D9��{8σ&������s3�>�d���4���d=9[�M�qٮ�9h��e�_F����Q��r��q�ԁ��W 7���)�_r�:f'���fǡ��Bk���m�.W���<�F�gYN���n�R5�W&���{����x��X:\ګ��R�|�θ���@s������t*�9�Py^���3�����]&��\��FtF!+]�r�xNߦ�v�&�M��qE�̨i�Ҟe���t�#��e�3Ur������Ԇ�[�Z�]Nd`�)o���BY��/_L��%�6���4˂魈������،�������9�^�~�R�� ;������
��i�
��Bxs=��C���߳U)��@X>籂F�Ğu�6�1w�Ϟ)�`͉����o�����_p�F�&�`Nq[pv�݈����*L����vZ䕗!�Y�V����N���&r�6}ރ�˳g�ң�%��N)��(~�ɻ��+���䙠�'�����\����S6݌��ǔGC���ϥ��>��h\�H/s�QYn�%�ș�5gjI���$Y��S����Y���@Zn<\^.��I��2�;/�3ܻq�s����$���qtr�������!Ȟ��&X���Z���	ρ�9����=G>}=�`��_�S�=�:���Za��͌gD��ѫ=�A`�#�J�=U<��2�g�:���C>���&�����1iP��B�s^�>��S��eX:�� ql��P\��
�_�{���S^�������kEK`z��N�����Δ}}q�}S��:��l	�� 4�3�a���2zxY�3���+ڰL�V8����>]���Ȳk�)�]U[
����@���P�z�Nԯ<�Bh���4���	�Ŧ��>��t�i�<}8�u�=Y�o�URX��T���;q>���;����yEpö�*���|=�3X��;����Ȟ#�2_3X|����xa�+d�b0N������Tg*f-��
����{K��q,�t}�->]᧹.��ԓjT�v��h��w�Fq)պ�zi��]9
�b��,���:b4�Wa\�Ӷ�q7�bMuq�o���j�ZH/��ְ�/���-@�;�Vv�dN�K�gV�����lɇ��Z�S�|TO�Mβ�w�ck��wF}FK��y��C�́�np��mۈ�v�)����8n��[�Y&��n�կvL�����^�:KU��DV(\^xRU^����z��鸉}����|��FNF�>�=>�ϑ�z�X�ꤌ&.��y�4�!���}U�绨q����e��ٗB�oP'� ��o��T;���Le̉�n �Y�MqD���Ҿ~����-�wg����]��8���h��q,�=���ΠEC�]�E�]��ZL�;��tD�}�;�I��@Nj�>����_����ӥ��{�S�Y�2��(ݲ����&t;��>]#�ߋW�������8�]��Ƹ%ܔ�ʘ���+:��G=��J[xd�����e��/�*;(3�"���t'^����:v���[�S��É��:��Mb1q����IUc��*������O�Ԇ�`
�׶����),�J�U�ù��}���u��qשs,�̢K�3O*�te��1�L�D�x��ja9yʯ� Ǹ�p�	tņ�w:+�8�r���b�$Y�ӷ�[��a���9�zVT8 �����ŗZ�\-��m�ҵ�!`�����vU�X#&TAMkc�O Yo��E��sM�p��V/U+D@�f�.�a��E���,��|�]�wX�V�t{=�%M�ov����!����nKߜ����/F��xC��Q^�gܑgɀs��)~7FY�4�*'b[��9����Tw�� �V����O���d���!��=�㆟tL��7���J���b����l��ͶϾ��7�q;+0R6eݺ��g�Xk���#��ڒ��MMNw���1m�w�j�1���G��=\1��	��Q��-XK︠�/����W#C&Ln0*��#_#��S��O2�6#x��b�C]];=vJ6�w˶���<�|��O�.G<��Xd��@� v���w�U��3\�=�y�E_G����z2utoPo���4�Fz#z=p+�u�2��l=6}8��[)>��'gzڋHU�e��=�sJ񯽗��������g]1;����˨d��r�
!��G7�Yj}���;y�13+�/�sq��C��%����]�3̋�q��'=߫Ы?F�1�r���ɏWR+���OF?����*r���������aL�_^�S�/Ujͽↈ�5�94��Ԇ	P�Z����ȗV*��j�n@������Ѭ9ovo\� A��y;������o'��0�]���I�,�B2c�{��K�)^*E|T��.7u$�M�D�;�&���j|C���u�έ�JB��쓶jI]�O�|7����Y���d�����W��^2�����^v�\��ˊx�WsV��G	�۳�.^�g�ֲ)��X}g	J���Fv����H�S��8ًH�tw�{Ok;OX������j�xrq]hpX�փ�A(�D�jKF�2��_*ʲrr��s��B����E�ٿL�W��b�zJ=���S�θn|�փ�9%��P$�w�'�]�݊~�Sq��Oz#��$��`)�}���Pv���u�}1��P���O�l�Zī�~j�3���Bh� g��:��@�m�I)����*�[�<2�[G��O�WA��-��Xb�<t��o�M��,eL�᠀�fl�Ger�����3��v���ݍUO#8�+�dz�;�{���}7u�\U˚,�ȈP�4I\�����$nC���o�z���Iv����
S]1Q�^�WG�����q��t����
���NA'p��řmr7Uz�Ux��<��be�b��cw+���GO =��k �}���K�阵2yJ"��v���o�8�X˝� �X隁Ԫ�+�o��՜1��V��q����J�&	YI
�Y�yD��>����@�G֋�pe��w1��u>%�Ğ��Wy����Zۨ4����� �aݩHdL�<z��1�&�p�x�t�,���km ���{�2�ۓ���|��
M��,y��t7�wj�����L�٥(t/�3]��j�s�+�E�;���F�O|OF�5��.(.k�3�-�z����XG���׺tA�.ȭ[��z2��B��b����	��\��CN6�
y��%��r9�U�=��d\�B̞�q]"�T�K������+�]f��t�}}0Ku�2;�l�����-��[u��\A�.�@�wr��t}[�s���rW.�_J���/�8���:P��r�n�dw�/��y&V�A^Y��s�Q���o���'}�ȵN��K��{�|5}�m�:h�jrv/�g�=L��ggc��}Uͮ-��������<#l�{��Y�r�Cee>�����/�s�QC��1z���uq>�ｊ=�;�@yę��::�e���r��*�]@��r�Q���V}\�;[�I��Y7B���Q�+:��9�G-IT�'��ĕ(L�N\[�5�{��q������M��yͥ57�p{ku�o�J|G��7�ӄ�@΁ �H��KfIAv�Ǟ%��틗?1�u'K�ǒ��<Ҵ�dYZ2fu�c����2�t��bư>2	,]��C����":����rJZ���f��ՆRՈ�%u�_��s4����[��|«yo����4EsλQ��4n�{��N��q�]��p���T�Gx`fWJ���ܡ|�ud7ڿ;�]��ӌv"�W��Y�7��w�[Sƴ��������PvW��k��H�Dx�S�<�.3�d�j�q7�b��>O�&��#��v�\C��d�@f�ɽ������Z|S�9��g|U`�zj1i�v�[g:g4�GNׁ����.'�8���K�>���r�G��3G�R �mp�������������=Ǒ<Y����5�Z#ʐ����ȏxU��Tӟ:%�97�!���b��xи���U:�w�cwq$F�r2n�o'ު�{
��f�a���S︠�t��n�t�ʑ�@D߈S��ǂ��U;�^�8�'޾Rl:���}~݂��'���C&hwODM�w�f�zD;�Q����[#irl�GY�s���{�瞊쩽TW!#]1��SG<���Ϋvs��CW{Ԣ�b$���h��@����_}�>��~�T[秂8�e�q��W][d�utg�'=�]��o4�y��Y}�{}���V_6s�.󤙞Tc�Ѽʯ��J>����L�/�N���� �q>2>�p���^;[�s�RُR�d�w��=\��%1�tţ[k(n��5�뾂�er}�tb&�j޾��#[�8�K���*lC�}s駸A)s������I][IK��Kq^|�bo��!-}�,k5A���̬O��b�Zx-��b�8�-�m.��4Ԓȡ�g`{��f��r7=m��{Yӷ�%b�J�()�\P[1�4��bghB�8����9����5n�E�Ѡ��U\3kQ��~�G"���c+�gK3��S�ʿMW.���ɱ쎾�Q$�!\��+�P�P���?]qϢ�TA��AR�}S)��	��N�Y��Z���;�Y}��Ⱦ��Oq�{���lv��z�yr���Q%ј���~���r#�Ӓ�Ƕfva�l=<�*&�R��̞s��D=7�R=�UÐ��.���78*�ȇ^�������B9�7Fx�5�0��n�8�s��ﻤ���u���]V��,�;�o$b��+�G<�TUˡ>=Ҫd����҅g��5��<�}m�Μ�l��tGֳ�:�]��0V����6��2
�#I#��u����7���}rƥl11�E`ݐ��fh�lv�c�{38��%�qC����
��\�dɍʉP/ny��A��)�������z�v3��;��wB�s�'�O��E��F\w]%�{t��v�g�
p��ѓWs?	�������,W�c4S��(�v�l��خ;/m7�6�Hn�AWN�u��xw6�Ę9n��5�FQ"��YA���
�Ћ{Y8%j
�!W�6���+r�j�1s7�n�����=L���k��v�su
?%w�]]��ڮ��]�7�E.�ж]����ho �u�{�ތ��Y3*����W3���Ϊ	�5i]��	j��>������i~5켸y��������T�>��CnPɛˡ�����ȹժL�dx�z2��..�^]N�|Xg8���g���೏��'N�R�mGZ�]P�F͍��F�*��0\����\m>E����Nv"~^����%����xU>$��d��:.�}gt͗}�Xȯ�7u�;�I��3�'ȱu�^2��X�8�mx���[xT��rs�]�O>�WViϟm!�yT��8JWa�3�6�%�/EWS�G��b�x����1�ODK�(غg�B����r����udpNr��|�t\�J5%��d�復�����R��b��ѝFq���.>%���^��vG��NEs��)�9%��-{�}y	�w7(�2{X��}�I���F:�$���ҙ<�f��v�#���Ɨ���WtD³�>p7���а-��]�s�Yp ]�g@��)@���=S)��s��[�<1�u�s�� ���`q��+6�V���UpqY�NC46+��1�E�`f���4�b��e�bà��/F�j�naΰ�%����}fV��`D���|3�c�۩&f�Y綨i�h�+�lo*x��r�ț�2L��]��X��>�{�0�ը�Y~��ȯD/J��|��{�.��=��S�����0d
;+��@,j�V���-�w��e�Y~�ϓפ�u>�g�Y���,���ٮ��K�,� 5�@�L��/Ǜ�ȍ�������U������|�=(��p"{��@����*�UuM�$�l��|�8nfϛ��/ٸ���U>h�6�T�|j<��m��+���:����O���Y�0{�������}��͎-HF��ϡr��Ѧu�����#C�9�ɡ��"��R��3$K��ԉH�2�A�Ј��s�����ç�U�Jk������qβ����gUa{�t������Ko��P&��]�t=k�a�q�A*��5�jy��%����U��)��x�i�{��L܄r�s�k�������:^>��%�2;Kdm��il�-UǶF^D�=y�����q w�ݷ�>uN����߯�G^K؜Wϼ�C�Kvdw�/�-�35���MUi�Os���i��Y7A�����1r�0vz\�sZs�B�νEe���6��WI� LX���Bܩ��Z���7	�=J1+�uM�z���0�֏&lQwR��Щ�2���H��2fɂ+���wN�	�A+��N��bE*�ə�I�vs�b�n����%6�����o7e�����U���0m���йZ)k�����PyK�/�����3�B+�n�z�{���f�_N��]�Hd���J���A�kF����j�|���p�Rb���F���DXC;3�8ҳ�K�� �^���p ��wp��!��F횃0^^���.:�s����0a�lOj�p݇d����l�ݳVI�ti�@4n�9qsN����|U�2����� W��9u�f]u�϶�S����so	��!bP��omiܡ�2�iE��z��(��oGv��rC��S,Y�Zb��׮n�W`�֦��4v���9S��{"X�y���K<���(Z��%�C�
���s(0�F�(tY�A]��6�k]&�u ��<�v���(���{J�1˨�%f._Aos �.��N�εx�WQ�z���dN��j���"+Gt�O�i����Nw)-V%̓3r��Z�%��T�f�w���*.��qT��ړ�	+iŉ�h�:;ͽ�F��vv�ط��"9U�x��r�m��qP0T�����ޫiea�}�,s.�nʐ8�]u�v�Ŏ6�H6"��j��)4��5ټ��z��:+�	5-�VVΗYYϳ��mp��(5�	Y�y!����Ƶ�T�1��:�*o�S�������('4�˘Z%[��v(�sFF	��V^B�gh�;���Nd&�ފ�a���j�N��8���Mmvp"Ʊ�)H�� V�+��]!���W�H���Cp��"�qf4|��r�u#!:�;:�blީ�ՙtm�0ݬ�Y��#�,޶�	��t�%Q̫Y����؆/AZ�Α执eL�ۙ�Wd�J�o:�3g�Y_J$R�H7,�EM(�5�A�d&��)�a{�զ�P9Z'��IݫmN�I�v���wԬ�ǩ �ܔ������nD��s�X��^���U�����'^����Ŋ��z{�4<�Ɋ/���:O@�j9�������۱�nm>l�u��54�-LR���i�է �n�7}��Mf�3
�5�ﾕiWq��Ry�02_X6_pT^I3���a�䮷���!&��s_��`�:��؄��Z��p#ݔXqTݘ�G�w�i���U7�'1���R�9��]_c�&:N^ym�nIw�����,f 9Y|H�u݇���^ӣ�ou��X{s3����������t�n,��+)o3[8��6pٕg><Է`Xj��!�M{����j�K�\�o�Nջ8M�����'�<LuӠ��;�\Ig4��&���ˬg/D껍��#�ͧ{#�����j4�ݫ�ru����e�_hO�q���������}��h �P� �Q�I�TQE\��B�(�J*�|e��q�J�TE�U�p�He�9Q�4YUWj��Ȫae\#��PU2ɥp�G)�'9Ӵ�X�G"�QȎTDJ%v�]�AE����G1
Njp��r����e��Gev�Er�9QEfȹf\����UJ�x�K�Uh��D�QAE�$��4���G	2�0�,�ŧ)PQp���P$���*�¨�+��Ar$��jȊ�.f"t+�U&vAQD�EgB.Qr"���P�D��
�D�"dE�Q���(L�k �E\�0�����9Q�4�V��L��RNsNr9QRItʂ��Q��pU��AB��Y4����\��"�UQr�˔˜��A3�����Z�����(��L�TDQÙ%&s��fQ	!R�""8r��QEU�Eq2Ւt�r�(
 �
	�1o<y]Ľ����65C����Ad�6�km��� ��Z`�Nv�2�����@j�p�zq���c뚙HIݗ���\�����=�x�Q.�I��)j�<�~��]kR�ݪ¯�$�\v2�g/�Tpu�]D�P&tt��!��͚�q�!��jt�;Ǹ�]��{�=�q yл΅�k��=��\rԐU|g@�y.*U!qU<�幠�����F9�9�T;�M��؋�{q]�r��Q�Nk�c�nT�l�K�3�H)Ϣ�P]��X� ��3���<��;@ϼ�����g5�q�"�W�dho_\v|7�<n�1�&t�F�G��;��P�/����֛����!�9��wϩ'��#6:�ث}U=7� r����kF�����b��@��L�g�a鯱i�w	��x���\GNׁ����.z����s��YGޫ#����U�T�����@�](T��o��5��;�5}F���<r ����Λ�o��^Ez(��)�H�YJM��H�cj�}�|TO�Mβ�clܪD9�q��_p�"�dȡ}xpK���Ni�v$xu��o�I���vP�&�B�w8��g�T�a����S�.��I��R�8�{�\�X��λ������	�83[*r|�)�����Y�B��sb��I���m��VF��ɒ�{�q�؟2��=|9]yz�`w�;!��6��
f�	��펎���td�8x��ci�}4�<�Y0V��*�v���s��!̨���N���>��_z����t"[#k�ɳJ����ӌu�5�EW[�,�>�Kp��C�^uXs�����˽졙�*$��������3�;�¬�]��d?��g�����Ė�>�utg_%�9���{�4^_KS7=�$1r���k}�;��\s�3_F�8W�������l��1z^�A��Z_Uy�d/u*�x�s��O��h���gT	�
OI��S��|b<]��]k���cY��vn?;���a�Uۧ���Pw��W�S�t��E�%+�,e:X���o�!��#��3=�~�����*h�� ��ǭ
ϟWqY�Hr�5�ž~��AV���k�*���H�=�5����%ש���o��yt8,�?�^�;D�g����u��qשS:o�8I����y���@���s��9]�=�u2�e��O�����9<�r;h����Fo�w]���r\�y6�9��M���7����`o�|:W��(�9��rݤs�3�V��p���\�io�B�ZPJ �̬߭E&33�\�C[�U��z2�iń�PD@�]�b�V�
�����Y�g쭜.�r���ץv�!�[7� �y �g���z�{K���G�ΗΦVko{�x�O����NGՆT�l���sS����%|5!uD�L���ބ����7T'J�퉐6`7P(}(T�ק�����c:sm����]2�r��8�p��ܺ�v�ݳ"��mT���$�W)�t�x�k�!��ڡ��ňۛ~��,)v�s�g�A��%��ƣ T�uCT�F�d��D���F��r�n���:�y��b�u��U��TÌ�I�m��ǀ�1Q`.���/��#$��"=n�MU�G�٩��skU�~<�-SCYy�]7uR>ޘ�����"�{L�w��C�zfsx�q��N���'AS�����u��Ag��β�����GϤ��:�܇�Cvc�0߰J�^�M�.XM�	���
5���z|:�����)�K4�q@?U��R���ۼq��3��X��}�Eտ	���~}>�W�0\���q�O�qAd�%ӝ����
_f���*M��������ɜ�M��G}=�xw��w������Vlw-'vʯ���>�xc��R�y�M>�u���2�`���;�~\:��sϧ\WViϟm!�yT����fa�f�1�]��iT<b��ѹ#*���=��`��� y�Y�L��
Q)��&��o[��	x��[��ܙKyu,��
�����F�?Z��{�AxFv�ew�g݅;�+���Wp��1�k�jv��GH������甃}�x��,_����z����d��ub_���s��c�,3�!c՝җOGf�����u�B�|�t}r�(���nl�ד���w���F�Q����	���
���/IG�=��r+�p�u�A��hWO��u^��l1.���J�pI�&n"~؇R�ݑAO,�ᾕ�Sݮg��vϟLi���\��vZ�s����p�N��l��7����'|71u2�N<u�W-�1)�+<��^��r}-��K�g��������#|#���h1�� l�����5�Y���; }��yK���]w����gNm��wR�o�����*��m���dtl��%vN�GϲlC좬y���E|팎��Odq�M�uhY��g�|��ѯz������ee��h�5��A�^F��-SC���
Cw+���� ��up{!��*e�=��x
������(k녮����Nf:��6vlT��B�����n���ݪG�s���wu�7�@˗��dQ���
2�]s��<E}�X�x-8*N��t��Uǥ���5��۷N��w����L:8��ƌ��ۇ`���T��IZS���r�º`�+�sUq`��(g�5Y�Bl0�K�~i�B��)�rA�L��S�p�K��Y���j���Y}�t�C��E��n`���c�*��wZ�
��S�PfY����C\�ӂ�u(w�E�lx�{8�<ϡ����r:����}\���l$0�u���܆{��gr!��i�}�]a�����Us9��/2�`}��|�k	��w���5U;�r�������t����d��G�Rv��{�.�&�wզ0g�O	ixТ�;�@/5qjz����}��в9��7'}�ԍ�8"jznkv�/p%]vIЉ�=gj��ȓ�;M�p7�H	t��7NyoPw{=�����)�1�
�eu�{^�El�_	��g���NC8��U@��+�=E%��OKgZ�U��t8��h乍·5�m9^4�}jH(��b�U!qU<��[���wбy6�Wu�Î�[��7ݨs�6S��!Ҝ40�'�����=;��}6�[[�p��D���+f*��Wu�g9�w;h����a���`�T�D@�Fc�(�ک{r�o�����s�#�N�A̡W�Bk���d{�.�oy��>S���o%=1<�4�5�\�f�7ʲ_ʾ�(�Brs��q\�N����d�������n^K�7Ɂ�o�QQS��"8SG�+O��|P2�m��K��E5pd�p3t��|{��w ����M�]l��*nfd]�8_WY��K����1�-f��sh��Bo�z	d�*q|z���Q�j�}m�����Nׁ��ױ�9X=��Ǆw+�cV:�L�����jKSd��Ή����� �8��=�5|/�y���'����U�Ur�J�G���D�q��uc1p^WI�S$5p6�TK��B��+����!�h%�B��}�U�(�Q�~tG>�����z+��0�\�J�`Nي����	g�Ս�oo�̎j��%��U�ODgu������_�������m�����Є3�FNP���Q.���5���ǖ�9g�Կ22��}7���Mk�累��5y�a���#ڻ.E�J���'��u�"q��jD�����;�VW
�/	�q�q�e���ND7<��]�����k=ݷ����O[E�W���p�@��L�\��^I���bbˁ7���)�K��Jl�/<�t��������t�tc{GN䪈Z�ѯ������X<_zP���o6�|xZ5��JɃ��dG	�Ӎw�;�ע+9e֜����C*�1Q=<�Ӑʧ��8(�����=�a��߳�z�7�>~��y��#2��,��e��"��O��5ϊ��Rƅ�}�F�A�㚮U�"�cfy��6�ݸ�c�җnO�u�5�)M�]��=�����	p�������а�J�;\�
,�����5���v��Q�]b߃���1=�]��u!�װ���El�k�#l�f�E�G���W����:e�3�Gw�ۡ���{�Dv��>�L?(�;K���,��2������y�.��&'���A�5���Ǔ~į��#���$/���=}ޮ���G.6zf�;7�W��%v�D;�4�t��R9gJ㖻�[�7�ns����⽔1�+=0�ݑ�rg:E�R��NpK7E��!��x�@+Ƴz�<��هW�����z����"��n0��ָ��N�!.��3��E��@j���
�����ս3��5�\�n��S�}��yQ��闤��1o{�*�+���1�_D�E��Qz0���{����+������H�%��\6����od3q�W��.s��(yu����Kͱ��	����8:$�9WQ�>��c~m���x9]��i�fT;��"�9����]�GX�Ѽ�>�Np��p�s�\�5�<�C������y�X|�@�.>Ζ���z����*�rvsbUK`����H����4��j�ߦkĳ]K�&**��[b�m�x9a�Y���8��Pӄ��w���]~�:Q�^��U�M'��
�о�o���.)�՛�S�2�n�#���|�#�X:����P��/u��ԫ�+�r�L��`�G�-��2���@)�K4�(�Ch^J�"��6
Ց/̝�g��=ܖD���'�Mq\}���O��\ $���O�[;��i��p��N�]�j�p�J���"���>Ҹ�1�Xȧ�Ҋ�KpGS�vr(�L����o�ǲ�9�Q��D����"�S]�2]w����҂���XTQ8 j$?fC&�_r����-����(�S�9zc����N�tׯ��<��Ѝ�޴.?]u���U�~�/���W2L�	�3#���4���4�z1�L{��(�>���q\���婱�%ʻ7�(t++�t79%\)@���,5P�*e����qd�5yu��}�#�R6L��/�\`2�,�롗����\��m�����k�y����\U)�[+B�g��ϕ�"�m�=��л�mr��3�wU3GeO ��1� \��i��Ng���S2��Q�D��zЋ+���s���N�����}wQ5�h�p���4g�CX�6k�u�El�,�y]=�cn"�,�Um�:*���Go=G+�=w�����h6C�O}�k}&�3���N�.�>t�C��g"x��YM�6�����9�R�u���.4�f!�!J���-��i���Q�i}}W�}ϑ�Gr��;���b�s��y'�|Bu
����=����L���.4��|��
����4N�U;���'�n�fWsDY���dp�ɇŭ3=����H��7���*\�yv@o�MO���T�����2+&M����;ţA�e}�v���nW'�ë�����|{=hɺ�~|j<�E���`�S�nx(�c$��xV�_�}�yp��e���o.<D~�e�*�0��opY'x����P���!�qC��PӍ��.+�}ŵ[�f*D,�����\��������<�5o���������4 �U����&-��+f���>�y�Ӏ�z��[�᪩ރ��.��7��#���{�gm�߶%h��M�b_�7�'e��
�x�*f�|��m��F{�=7�8K��}ޭ>綇}�u8��u�"0�x��y&���^������Z�bPchȲ�z��Q��9�(��Goޣ���"��]���ħ(�4�D�
�:�L�C6laUULs�;qA��?wb��S(����U�p�
ki�t�6&����h�V��^]5��歳�H����X��Vln�][�U��؍Y��\���6i!�J)t2�;�qnM���׬j���7����E�@�!ֵ��>��S�L�$�b�U�ũ�ke��n#'zO�f��;�t�!ΆJ�+��L��$Pf6"ĕ(L��)ݍ
챑w�7�ټ�������ͮ�G�ێ[��7C�hu�l�hC�8h6I�������ޏk�\�����na詜���Cb[����<��mU��	�}}q�7�!Wl�����sWV��уf'��MD"�4�Ȍf�y	�mb��>}1�{��#�]vġе�D<~��*������R�z��̀4�<j ��ҙ��Mbڇp�[g>����Nׁ��o(̱_�����5g?C<���m��9���	P��'�5��_Ŧ��&��ї9�����9��L?sd���������@�I��!�V;Ƈ��ᚌ����_8ܾ�sȮF�}]#yw]ы�Ϭ�Ǡ{���>��
��P�P}F6%��t�n���˼�냻�F�6c&3��1���ȿ��3�x.��/���@��fJ�0�.�őӷ1���Ӕ�����M�x�6�߭l8O���zξ�Ҹ{�F�Ϸ�E�w�b�|*�R�C��'���^�J����/���Cy�:AΫ"�x4�x�i�%��[E<���[B�d���Ŗr$:��7`�S�M�d��rh\�����%�I0kxUpbp��ԍKg�*��\����8]u�3�{ˮ�a���d5�AD
��ZwAÒ��M�ك跦�⒖��-�LMg���W�N+z�ф	�WoS�����n��+��\f�E��,��,APf^�O\���n��	�{�e�^���K����9iX�֖�.OQ0����u����a�i�rZ�8�e� �u;G���\�`TAFH.��xx^̕�������e���������l���	��'�Ŕ~�"i���͝�a�k�����U�TN9ol�N�d�)� ����(r���qi����n�ϱv��A��ڮ�!���ZJ`|2�N;�n��TnI�ْ�`��T�v�6�5�	�[%�xej�#*�qKPD��vt�z=���VDmuM�����hs,i�F�Pԗ��[��ܻ}@�x�v_rq�`N9�E(��S�j���L�oR���F ����=$o��;yK�$W���u��VZA8v*N���:��@�kC���ٵ)���4}��"�怩<�y.��N]��S�&s�"S�[�Lƫl��Uzn
������z�IW���e�؍mT2+��9AB/��V6�:t��/Ab��jSb|*:�u%D��� ��F;����,�C�Ŏ�&/�k(D�Я�� >�p���5���ڱ� QY.-���,.�}����-���q/�K�{-��Hj����6���Tj�S���@��]b_lω�M%��w�øhgp�Ol�9_[t�6��F�f�M{1:�P�r��|���a�&�sKT��tüт�3me��D+�d�.�$�����ѕ�g=HS���qWm؋Tt�x��ѴNᇶ}%�=�#����2۠��6��}f��c�	�Q����h�����bL�|�¥]f��k_h��}�X�%.σn�Ȥ��ܻҎ�/��:z^��";�|��z j��fuf�+N)��;moN.9A�`�;�;i�ʄ��l'����k�KN�W��/+r�T띺0)�7}�v�ħ�8��I"��װ��"�3m��kz��L�iI�I�;QvXoK�ΐ�x*�%���֮�ypvme�u�)w��M�lvැnSlj��frf�uWu��N�4�B�o-ڋ��Z�P� l{53F[��<���O�m,���b�6�Q�Ϯ+v�u�5x�\��湔��鮸��Ѧ)�dک]�9��ǖ-�D���u�I����n�����)�kȥ��7��Sm�3+
��Fi�5��.�^޵X�Ԭ������iLy��&����je�q��0��=��[����ь����f�H�[��N��ȅ��;N<X�?m��#�}��%��^18^��cvc�Y��y�/+� � D|	��B�8E�:*�Z�.� ��16�Ad�Ȧ]��W
��U�hgC�P�J'"*��t�����D��E@U�S"�U�*#�vTh��j 슂�����*UZVHZ�dEfU'"*��I��REr��D!	���X�j��B�r����֑̂5�Q�(�;*�*�U���".;3e\����+" 8QV�ʈ�t����QDN�!���L� �T���#�G(.*����aQ�ʢ
�EUEHi�U�H�]P)�����¢(��Ͳ��˧���� ��ft�!PPQa�R�u�L�Vau���fHTˁW
L��uMePr�9Q�Q�e2���PE�2�U%��)+��e	�*�E����(�*�j��>s����������\!!Sغ)�>���s�������5kG�L����o!��:��l�9t�b�v��e���u�q�%�$�� �;�@/.��h��+�{/m�UU�q���G������H�+$�����ͱӰ�{7��d&�e�;�K�>���9��:"j��o�T�d^�����;�{�����ٌ�:�{�t�tg=��r>����N�u=G����>pS����W��K
�7]��\`g��}�{����>�_g,�҈@HFu���������k��ƹ���[�b�8)���F�z�Bǽ]��ϫ�L�#���tt����*�@�r���B��%�ͅ��I6�����a���Oq�G�����lv�u�A�ʖWi�wӔ�E~Q%lq��&d[0���2O�~y0g�⸎s����{� �u�:�������
�8��6}%��@��N�!L	�ґ��:W]��ݡm�qZLk�mu�ܛ����)�9���#����ϧ�pB.�@���D�^9�:C-�BUd����ߛ���'�H�oM�hwu	���1:��_a��"�uʊf���=�����f���}(m�!�P��ە+�v��8��l
�\-���W��E���$[�ڇ��GqQь�����ؕ��z7�a[�V�h�ԩh��eu�	�F-]�\tf��;���wo�KY�t
G���a4M��6����˹�������zs�P�}r����<��}3�Ot�@�>θ��S]F��A�t}����D�6�zU(*�4x#mʯ��ry�03/�����������n0
}��e��F�P��2zd�Ể��N�㴁w.oY�ƽ��cutq��g��/��ɾ�b&*���ϡ%d��p:�s+�������bl�GY�k�u�W�o���>��GS����s�`̿��	����s��]C&nڢ
4rXW���;�N|�Y,��6�^��+0>$�����f쩛���&�u��U�Vw�Qߧ8�g���?�������qal�Z��^����.��\b;�?�}�k�>�Y���W�;+7I�wM�w�>E�7�4���=br���}⢷;�>��W��E���d�u�ҽ�uxj9�i�s��9��%z�]ʳ�2����>z�L�E���C�2����pTx��'K�k��Ü�!����=ybgO���
9Z3����:Id�G�G\Q�F�	��o��)zJ=���J����, ��!C��R�(Z�q7��tfݎ��ڼv�=T�YX�SVFu��͂�J���U*);`Q�]s�I��Y�vE3���ֶM/�oHy7r��ѵ������#5�Q��_:̮u	�64\�MY6�<RQo_VZ3�q��
̝sF�Č;l��1NV������%lL�9T;���).Y��}+J{˼]Ǩ�����"�b� gXxi�=��Σ������D���J71R��;�ћB`�u㭝Հ�]w�T����h���q�����vʞ6���:�و%novzn6�^6)����pu��Jcz��rڴ2�Z�;�Tw��t�S��}�4x�2 s��[�/�)i��Oc�ר
�[<��0�{l�7���9[Ǹ'{���늇������Ѿӕ
���ﰢ]� �� �,F�;e�a��Ŧ��&���wR�W���ǬM��wSu�1=�EW(����Bu{&Ed�����!;k�I�>E����#o�ܪGs��n�P}�=�0����/��2S�ϸ׀��EG:�ҧ ��V6pT	��\N���:�����H�>Ձu����jx>�T��w�hwO7ڦ<��Q���	��9aˍ���pF���^زtMzV������F�6X�{.�!�������3gM�;��⴮̪����0�.��!�{os2���4d�7^{~�R[0�m�	������FW����ǟ�˞]u�]+�����O\C��Ȭ?
���z�zo��E�Jq+�S�F,��*N�.�mB�3���+��J�aF4y�^�R��*���y�4�Κn �Y��Ҏ71Ϋ��Ŋ����:\6�:~���b[Wvz�v�Tr�y�^	^�y�nŏ܁��^���$��x��2;��Ay&f3��kb�*᮪��K��}�w�B�^�V]\��R�G֚=﷕ɸ�L��6�]uW�����p����"_��yj��^;.N�CG:+��۝ی\{�z�y%L��N��3�b��r�	����9dլp���կT6�}����}�=�<�(u����Ӭ�>�VI�@(��R��6�n꯮�m8Q~w�=��Y�����u1�uv��v�8�5r��%����R7��vi���zτ���EL��<y�B�%���by�ϻh��ޤ'��_\tnL�n�.�W�����y]-�2,D�mD#ӜiL�f�W�BhN�{#�>]��}@y�uH�o-o��F�{�������T��ȀMD��~-�
/��N-چ����Ϻg4�f/޸�t��s�X��E)�ó�b�j�3Z���C���gຐ�/O���Ŧ�弊���-�uc�EX��5K��W�=��$Q��$�]����_RB�n�S�-�}Zn���:��")�M�*�>��֟��y �(��T��Ө���sx�͈4�g6�\Hغ�Rz������]��\��AbB8j���;��a�e���QO�vsϊ���9Y��(�2Y�%w�)�g.���Hj��U
vo��[8ʬ��vxOrB��ӁW4{�ܦ.��ʤF��<w���҃�a��t�S1������-I����y�\&���G.�ePs��6�tn�J3�o(ٚ����A3B�4!gz��!�ދ}>���Ǯ�'R�fw�;�:�Z���G�{vX����cWMi~��gU�;8�hj������2oѼ�M�!7$��>��E�:}=����%��ߪ�c�bK���Q�/[���%��1J��}�z���Mᜢ.;x�6��Vf3��l���C{�qȼ�r8�7ׇgjI���Or�>�H;�ھ4�|��gv�ӹ3�#�ꜣ�t�r��X)Ƌ!����PR�];X�d��v����L���[�]����0��a��|Ne�c+�gK�x�`�-��I���ߟ��>�{O|���*;)���=��B`WWqs҇k3�a������*'��wi]Mӟ.Ȟ���gkE�L�g�	�B
�y���_{��l� �yשa;3���Ǐ<�؛�DMf-a����$ඃׯ&���K��{9�5���JǸ��h"q�n�g3e���3'0A�s-u[��ڞ*0
WIRY�:�xZ��S��������%M�u�Rn��W���u�{yn�r�b�:*>��qLB�n���g�$����Q�e�T��Cʨ�į���s����{ʨU͂$�g���q��C9ׯCϠl䞷 ��%Pk��٤g���Bk�ݬe�y����.Իg�,��έ>�Ϥ���u����l�8'��8!Hp���*����-�F�~ɺ�v�WxL�WxgKw�c:}u�Xk�}Bn�]U�b��GM`1�Hv�Tg�f�s�x�k�4����к#܎O��8���tϙ=�A��^�d�#���W�Itm>o�^���Rpѝ��o�)�j���u�C�����:x�f� }}p{rz�B:��^�ޜ�
�{Q�I�4���M��45��lxn�k�n.�4;�����[�66�A�bg�]6/��:�5�:!GY�j:n}�#��4β�y^���U���rz�����s��#�|��� ����r.f��OD�2�ˍ��å:�f�9��z�lgU!��]W��FdQIp��zWa�,���.�Y߮�w��5�~ ����
�z|������W��y5�N��&T&���2�X�A�w)|����p49�pW^�^!1����L�PJ�E�q]�YaX'2��l���F�bd��U|�U�]���ͥ/�$makf���^�ޒ��Վ]2(a��p�79po>ib��
���{�>"̗�Ҁ����C!U?d����#zk��G+L�����gúl��#�h��8�m���[��{�hul׍Ӗ
��<��/�\� =�_Guxj9�i�?]"�m��T�\�O�����uq�Xj ��9�g����^.���.�_WsԆ:��wS{����c�VWP�羺�8I�3hmg��GDf�g�(3�!}�N�o{(��~��*mK��9��ODWm!�9HlC�^���	*�n"Dv!��̑_%�4����)���NҊ��ண�xgLq�_��w;��g8�8%������J���7d�\6����}辐���=xU������mD�������v@�SƆ������B>�m���9�%�HK�Ȁxn.�6"[V�7ԃ�ܲ���K6:�h.�'��X|�D/ ����o��HL�PK�}�a���l'������=�3�����Z׈�#�Loo��k�v�tW|�}:$���d�,F��-�7��e�6�r������K��]�6� b�7y�4�[�fbW����n��)����8���	V�����U읛�u�Sn5��d�����!+%�p^��ӽ�9}1ٱs?Y�][:VP݅�&=%�K�qE����-N���1�e���L7n/!xB��������2�8�D!��`�K�阵2Z���DK��Ry����o��;��U@��Ś�U�(�Q�N�2o��@od3^�z�\�J��sт�G���.=��No���E�xz�4=�<Nl�)8��3uUQ��1�S��zw�m(u|��!�qr6�i��)4#�'s���=���l�pe�����F���vx=鎙�t֙��
�g6u���u~aȫ��%,~��y��Q�&쎟Oa��\@5�П��c�b[W�Cu˧#zht���mxc��Ŕ���1���c�S�3��VM߾2;� [Ch/*񐸕����þuT���u�yL�m�=�Vf<����#,����������;�Uɸ�	�x�f���rL�:#��:#̺ ��Uv�)/�V��R��=�GOT$VE>���>�c��(�VN�S,e@���yL\E9KȿY9�����2����g��-�N�G�z{�Ob�e<4��+��d�8��z0AñՉ��;��ϛq��.��T�s���<���Gh�c���w;�܇5�a�ܩe�Ir��_����v�#@�3sa���ت�ŷV^�}�����1=M����@����Ԇ7W$���
k����g�,u���+�Y60����¦��դj�{]�����l{��b���o+��Θt��'w>}���5���W����=�@���������
���O3��Y��R�����G|�=~[���n.�����"��G��u3��{�&�[X�9��wϨ#�u�� ��^�l�p�l��*��'U.m�sQF�-�����0��-ۇ�/��<�bQ8�D��"���C�/��m847��.�*�;32v�'rl�6B�B�����yr#Ӥ/��q�K���4k(�_o;�9�L�'�㌗�l�8йu]&�L���ڱR�xб����Y+�[��"�"����b���Uߛ}g�t�@��f���E�9���
f9`��kޗV����k��w��ӏs��z<�Χ�ڥ��3�z!�i����j�z��
ǛG2�铜"�nP�~"���y��Z�p��lj�.�5gU�;/�T9$�퉙��Ps�]�]�=SC�qA�n-�����GY,�g8����$��S~���Qt�<�gliQ�\x�uR��s�������Yta����^J��q>-�����߀˱w?~�,�ԫ�.]Z䫖l����܉K˝v��,^O)��ӛ�ȫO��	݇���U���D5XNRcq���z��@��9�_5r��)i}/�V���i�ֵ�[�.��fƦf59���zp8�)q��N"rn���ygag���������ܯOt�����>�57�K.�xeJ�(�M��1N����_�AEO	������o�N�������>�F.#��t�E�% X�V�I�V���ʂ�+�[��4>�*9\�3�8�49x:�<��g
��w�WR��y|��G��RńW�ϢD	�`:��I�3�,eL�7�t��ǪB
���x���up�W[������o4�9�j%Eeu��J7�J6�j���e��s�3�*�q*�>�9O�ni�&��C�y�Bg�T�����϶#(}�/_�9%� Nw�:����єw��uК�./���VyV���O6{:_��$��9�L9�Zv�t�'�h1�T���](Wp@��b��gS�_���L��,�;�t�>��/�rɮ}Bv��K>P@j�H��-{o�a�^����r�������@{.�6�>����g�GL��}�q�/�늿�J�C���gm�oK����ɝ��蘀~^�:7����L9�3v� ���n�����������6�����6������l�1��m���cm�����lco��lco����6��1��m�����m��cc����cm���1��61���cc����cm��61������6��cc����cm�661��ݍ�cm���e5��F�� ?�s2}p$u�=�%(��R�UUP	R�P�TB��@A)�DD�UET��%P"��JR��D��	$TG�}I%P�*���J�JKZ�H�
��%��T�])BQP�D٤�b�R�EِJ��R(��$�D*���+��DB*�*��B�H ���$J(
PP�����" �HI)Q �!$��P�"�)��k(�QH�2�   8"�a�B�ښV*����k3@�Uj�T��a�� *`d�`�AD�QUASU��v�6��)H���II'm<   X�(��a����/]�T7�N�� �GF����Q�ttQ���th����\E�@h��  ��� GG@ ]CQEf�⠒QABR�P���N  7 
^�]j�(P՘��mR���Ѵ�m�)�5VؐL�P��Y$��iB�b�5�3�(PQU�F�(T�  {�N�u��E���ݧJY�@j�Ww�ۻ�r֡`�wn�CYCZ����҆���ժ�m�
�,S;X�]��@ U*R�J�Q�IHk<  X�omn���mʘӧ]��]�*�֫k,�V��ݍ.�����X֕�� �ƚH&��t�]���jl�U�"����UACH�x  'tY�h�Y�`B���E��iѪ�m��vUE�e t�tک�cM���5f�N��F�Z:����� �a�@���%[bR��T�*�@U�  Yq�N�wYLN�P�٘��4��un�\-�X7l�%LP��:�V:iM�.E��۩]Em5�ݍiY��,ҩF�UkR2�$UP�j�R�U�  �yӻw[�t&��n���GW!�)L�hm��R�5`)M��h	v벌��j�(թR�]8u3J����Kf��VjEP��T
+�  j�
�Y�8�V�
i���h:�­�pt�n��V4������(Z�	�ڥ�Muк+��t��.5�vv�i3u���kr��(��U�H��O   ��Яv�,eB�֪�V���PSX-��mѦ�ӹ�Ŕ4*��R�m�ttpm�v���7Z��x)�4��J� 4hb)�IIJ�  *y14���  "��	J��� ���Tڀ� i$����  �K+��`x 	1�ଠ�b�r��\0tV*�~��Ͽ}�Ϸﯟ�B����	!I���HH�	!I��B���$�� ��E����{�5�<P��Z b_�V4����,VDq�x.n�m�F�����b� ��b��k5[9a7OD�����^&�b����-%��&�x�Sl�Ԋt���SR����o�Ac��Z{���E��=GN�C7��$דj9V�ʈ^KP�V`�����l�������"e��c!�i&ƓYhM� A,���P�����]�KM�����i�yH��!W��50e�֐(��U�E�y�`�Yw4A��g,�f��E!�fk�Zإ�[$jMV��*엨��+��m���`�S���ۦ�)�k=7���P�۹��x(k��F���`0�ʼ(�T�4�]Ո���Jr��2eAQݗyx½�oc�X��J��ը��z���2�6}�3P��+Gn����e�A����/�� �M��a��Eȕ�܎�O4�q�U�a�u�ǭKm0���R	t�ث�*�ͱ�-nB��,��X��m}e:�Ѕ'N�" ˿���	3K뒎 Z��܊Zݍ/�ۭ*,��妩��I9�J;��H�5���\;4ӳX���/$&�JICX	��ݫ��i Ê��bI��:���&k@ފ̡u���Gh;hrB�reY�z�7yDH��Z8]�:�`���:�6db��Hf��Pc�W�M&VCX`���k!��C�a�&�[Y5�=�pY���nF�[Y�5+6���wqyzCtq}��J�x���n��ٛ��rkk�2�ʱml��,[B3$?if�DHF-6�'r��)�{��V�HG�a�L^��*G���x�mj�ǢX��Ze�y��%E����O�6I)�"�a���Q�Z�M7co����iF�ŷ��i�/Xtr����H��oZ�cMJ�P)̡�S,�eЕ�ޓ]9�$Hb�^ro�rށ-�u ^�fBZ=X�S!em�@
ҧ��\�xi��"��`����^	�Ĝ֒���� ��H^��.�eX���1���^�+ehh�Vd�J�0�t��:�T�b�х\-��1���#�����n�C(��܃Y��X������m�{R��V���A$V��Ylbv�PO>m+t�4�Hq&�k���kKF��x2�J��'ь����պ"�P��5el��
E����_�*�Љ�U�sI�C�+6��E��tY+&�-,l�h��MN�Q��j0Z��(^V[ŵ�����wH=vX��sUi]-@9g(:#s\�ۙe�M�.�B;5��b��WStJ��ne�SoE��eՙ� �C�IJQ!��|��cŴ�`!������I�3 ��E���\f�ƛ��8�H)���,�bJ�0MPh׮����I��q(fY̫ƕԝ�D\khe�m]f������1C(X���̧�FU�� ��h䬉˭]��nݦL+I����c����ZbI�KpG���̼����!�A�V���V$L4]�2�ɸ�=�C�d���юS���Cx�Z��<*st��Jwm�c,������nQ�"Hj��+�B��B���M��ޤo�s@�
��b�ݦ�V�e�y�.�7z��&|���&�R�ncd�ۤ�aN�ײ��"�[��ĕ۩FdQյ�*��ln��E.�5��v��
�(*F&[ӚD�����u����)�(�7ݠ(����B���75me�-�򮣬(��qJ�q��N���Y{-���q�6ȃa���*х�Y�����R�Ak��7�JW�nu�P�s)����
qeY�KKY�>7A�:b�R�6�wQ��Z�m�K!ծ�z�
!�Ƀn"ْ��Mh,j�F�;VȦ�A��r�0��(�Ңj�f��� ^;�"��+5kת�ea�Vjƨ��)`�kiQ��/Q���B��ɛ������\���X�9��w���=�;Z�b���DK]1�Y��iV, k���Mm��oNn�놳R���!�~c�sR���^٬�`X�ts�R�Z#a���l$��K��j:IP�`����X/2�KV	F��2��ɛ6�=�3�2�4�X�%I[A��TʗJ7�( )�nS8��ik6(����!�j�|�b���Yэtp��[I�P>�G���������8�
H���Ӕ�8�A��O^n���X@_[�{�=8ij����e� 1.#���T2��͊�l�cUĢt5�.R��f!�ӭȪ�5���ͨ�V�i��f^�M�[�}��u'�m�7�n�VeE�O t�
f8�o>��V�Q�c^�Rà[�L$WLј�A�7/
�^+t*N��FkX4���0�(��z�Yz,�f��ha�6h����MP�o*�b`��an$f��V�x5il]5o��#��]ܦ+U7���`�u�j����\wY�I�V%y+o��G��f�b���1�1�e/��l�V��A�q���ש�6n���!�Xš����]�ݥ���nU�PZ����Z ؀+l��[�b�X�ÇT�,��%Ri�6��˫{�%xU�����7�3#W�B���#B���Է*x.M�!��Ź��+ZTV�������U��Z7Ն~�����VmI����b���T�6�T�j��eՠ�2v�f�Y��7f���!X��gSI].�Ȩtv�3u0l�cd-�+)�x��zӖ.���*!�c� �׍�ŷ���P�)᭔�4��[���j�{tV�l!3q�{��\�ҨH:�j��[iɇ�P*�R���˖��)z2��ˉ���,�FQ�@�)�Y��)j�If���J�k ��}oo�X�U92�*R"��ٴN�u�#kv&C�-^�vrd�����Y�X*jt��n����.�a�wU�B�MV�C�X@���5�AQ;���B�ƥ�[�F(�>�Q�q����t)���DD^2P[28�źlPj{fΝ;i�*\�@���?EJ��x`l�HʲP�twb໢Ȧ\nM�*�\�)=vټ!���=4H��@/�E*�j��'����*�y����Ee"UBL�o1]��w-�7ݺԜA�� PfҐ'�5-�wQ��$�҃���
����WrÄ��*�dyh7W�u����x����u޴YM�F��݉�ݘ�)N��f���`��ɢ����CJ.ʻ�W.��F��c+5�9&����H�Z�f��&2V�r�Q[��*X�i�h�w!&h�J��3m��v����t��!����u8���ۼ��i5fL��B�Zpf�˭���xun�n-i��u*QA*Վ��pڥz4<�x��I5zv^7�����G�E��wI:��Ou����ؖfՄ"�{;&�O�d�����Ӏ�	L���	� X��2�	�'m+f�ֆR��e\������5�)M���Qթ��% %h���M�V�-�/�׉7m؎��Uu*�N��?0�_s	�����;"�p�jp
G6�Ok\�dXÉY�3����N�D�D,�â�|�lطK�4�\�[��ڏZVT�K`,)�'s�y7v])��i�b�8��O���V-��`=7wP!��[�
�4.JaWr�p�Z����ʖ��&պ�m��{�R�%�w^�W�Z�,�������ձ//&���Q����驇��e��Z���5��v��?l�N�LZ*�ǣ崵Tn9q�,Fj[�h��HU�y�Wd�I�֗�5e�HҼFV66w��$�)d8,�g ����&��.�eԡA;�ZKm��u�ã%X[um����9 ,x�����`4�kId��rKY�ho4��ʘ��1R�72� ��n�H,=�2���,ı�ml%5t�����)Q�C�$��N�R�c2� ���[�( ���}��`�i�I���l^��2�lm���+{1[�(n�۱I���;KRgV���X�U+�y� I�f;�匡Y�v�ö��`�����*�ꩇX-�B�"B���yx�6�RJ����`ɲ]�r򁍣QPطY/r5���b�U�+F�y���ԥ2ކCF��R�;ʻ��x(��n
a�f���c�Ŗ��67.�^�wx���!��RRgV�Om�dG��h�)%��l �4ۈ��f&�2f�k�XB���{:���nA6#*�:�#/ �k]X�C�[J^��PL��\�(���%� ��kZ)��{r�!UiJ&��Z�k�q$/mS�.˦i���j=�բ� ��%��X�n�M�y��� �aЯM	��-Ƭ�t�
`VR�i ۫���6��䲷1�@�Ҽ��Pk*تǹK�U�*���J�2�ુ;�躴2�,�u/K�"=U��y%'�Ju�)Z��yk0�Kӻ���+LB�D������F� �zhAGV+m��5���
�bI�[�p<gք�S���4��,E�H��.S���� n�vV��Yz�aɃ�z�6+p��
�ݒ��0+R�e+�Q^�z�e�t�iX�ţ*3Y\��P�%�Q��3+��8[3q�i�f�ѭnj���3
�S4N--�	z6�˴�Ƌ��j2� .�֪����]�d�n�*�n�2^+���S��09&�̖+V]
��}�v�S�w��m�{����b@�R'YU�X�֚�VdT~�,��T������n[@[�v-�JGL��0��˽�N�Z�z�����)��Ra��n$�[d
mn.�7�:�$�L!�]�[��S�����X4j�Ƕ6��H��kx��]ZCT�
�R��N��V%�AVe�(-�I�v���"S�o#���E�=i��n@�V���,ҷ��,<����3S�@�y]�zU����mrK{X�m�Y����q�4�ə�j��F�:��X�1=�l��������e#t�j-8�F�%[�v�b�؅f��+������6v�V��z+S�jV(��j���-����)�3 �7��U�j^��� ,��
[h6�i8M�Y`�,m#.ħ �FG��2��`��Q�VҌ5u�jJ)%BCyv���ra�*�H�P�#��jRkE�����;d�4S��Y"Z[r�9�]�hֲ)��9���m�A�6.��ڭ�0ƊqI�*8i[���w�$��0^Ҙ"̭*�GP�F�F�`DՔP�<�=g���\��o]�-�;�)�%K1;�#�SrcP�!n+bI�l$i!����-h��H�i����ʁT_m<T·P�X��;�\osop8%��5E��O�C���l&�������e;V�&�*͂��SiV�F���j�YD��������Jޑ���n���6˰�d�ssEr�`l���+Zs80��ŗ���P�^�Æ㽉�U�H�Õ������S�$D�٫
C�N�sj^]�Y,Prl�KjL�N�XW�Jq㔖'�R�t2�h��J�$n�̭3U�L��1��QD��@��B�7���X�]֢0`5 f�W%�[LV`�� z�#�`d[Q�X�o��{x�U�kie���Km5�b߁�[&�����唱PL�.�(�,*x5Fi�x�E�ј�ք������k
/2ka��0�!��e���rS�`ތJ��G�h倪]��������u��3)���8��V�̷F$��Û*�:0,<>QڋHT4	˫�t��x�$��,�W�kUv�2��ݻ0�:�M����{b��j�]�#,�����Ը��4欻�u1�B�WK�Ud(㧹�������W���u6n��ᙛ��U�"���Fݜ���B8�Z���΄U�4�[B�U��0&;w�q����F��R�3�'ej��'.�-�(�5fƼ���9p*F��%��M[���Hf�&�k"{J�`dXb��V 5�;Y�ar�(���x�ܶ쪻v��vݻ*5k(ИB"�C���7��V8��"[�L�¤�;ڍ�R�ô��H�h���R�$����ˊa���b9�ӤS��v��e�`������7�iGJ���BĬy�ZҺ66�GL��n�7�f� 鑘F��+�ɿ�wX&9��j�.�����)
NTPP����ܔ4��aAc��0�F�%�y��=4t'{Z�k$*+�66�k(詻p�%-�kS�n�Xߥao��#ڗ{��:b%����Ӥ`�VJ�i���,g�j�F]I�6(.����L9�:e�4�IkW��,�:fV0�PU��j��Om�f	�䭡�t�-bmF�P%6��,�+q��em){�\xR,��Mk�����]2��#�a����FQ����A��9��f�]0&&X��i&L:1�$[BfcK>�,*-��c;�F"F@�l�2�̂V�)
-*_K�����2�f9P�+N���Q�*�;@+5"�慘�������X��s0�٭���$�u5"0� U��ѻ[��@v��w�x,�,�%0L����Z�Aݥyq�CԞԣ�n�
�uZ�B ���;t�M�G�D9Ԇ�r;�h�)���AL�Haz5|���ˢ��	0;P�,0&p7/���������/q.��}ԡ@S�^m�
�L�i$�fݚ�Q����L2Z5����Ji�E�J�L�
:�	��a��.�b \J���R�z���
��Z�fƝ�\ڵ�#�R�W�v/%��P�+edt�e��j�[���b�A�#�Lb��
�z�ئP�G�)7]��'q8sCB�^ڟ*J��6p!���/��F�D�z����Iܞ�
�#f�"�+ĥ�����fllEV��a6$r�,�}��t��N,+23����"�{ӹ;�`ĬN�߹J�;GGu�����>��2e��+��ٗ�t��G�e����I��^��2ubĶ�7��g��+��i�F�+�� 蓢�=;��h�|��vN�MgMޥ%��xc}�.qrS�A���K����$Dˮs8��M�8�]䷛Hd�}�@�\lE�k:m���~|a�����.�{ɲm��#��K�8�ǖ2�ݧ�%��]y��T��p���g�i�_Y��Ep��S�9e���c��t���[�I4e\Y�V��t�Y��Ȓ�'k�(#�����º:�촗4��7AN�a��qհ��ۖ\�K[5Ws�F��vf:a�f�ȅ2����G-��f��f��`nu
�C�H!���a˷L�O��f�j7e�@��5MY��=�6^�qͩ7(�̾R�$d[|�P��\�����gem�1���޳7�V�.�u���O�O��=z�s���ÙFhU"W-
)7ۜ�����-�v�[zs��7o*ƍf�%��$`#rc0�7b�Y\�v뎏BP{�s��f:-R�홝}KzF�u21=��1�����؏t�
9`i�EC�-eXٜ+�-�!���O;#��<�ǉ6�L�غ>E;{��j]���xdO.�K'Vf����(2�6)��4kNg]�k;�Y�x�d��T�����봮��+'Kԥ�1Ǭq�"�F�1q|T�ݦ M��f����K�:�s݄��́̕ˉ{�;�.�A.s�È��Z���tn˾Y�#y$���#@�\����R|�kF:��V�o+��[�V��[M�tO��^7W���'�o�R��������R���Ngp�;4ͽ�ƭrP�Ȳ��d)�pu�VN�#��7:�I�\�PǪlާ�r�:�]�I[��&�Ig��b
8+|l�9�����r�8���Ź�8&;����'C�8RC��YUu�Y�@A��и[�<���;:�p��_Xͺ�u�w%aDy�g�9̾Q��jQ�Kw���O�rU���xis�b��z,+ݫ��ٮ����l��j1q������m���b�;6F�����5�[�A��;p�p���g��!:�<h�̭����b6D��|Bj-�i�wA�s�n�s`:nb��Z�H�J;���E���<�5�p�0���hk�랍H�u��up`G�P��:��rҡ�V��rQ�u��m�f�Z��x�]d��ս5��Le^:�K_;�ʊ&�g8����Yw��>�6]�h�W�T�;s:�c+NJw�f�5t�X5�B`�F����{�+��N=��%ݤ��<{�'סӖ�
�c��7������ ��f���!Pd�Ԧ����}I4vdޙ���4,wl�4�t���-���˖���YBp��W|]n��s;/F�^@�����Q1>yii�����)K��z�|�^K�R�m���pR�Tt\��A-7HvooL���<.����ݻ���k9���Ԙ���J�u�C�3����2s�b$���M����U�SɜPT���c�ԣi.v�������T�_y��Dl�\���=5�f^c��&�y_7�Ү�G��ʒ��iw�# ��*�X鎘ÈjmU�x�-Y��X����x���D��H�z�wոp��S��m/o�� �*ہ���� ��4՚LP��Sž��t�P�Ԯ�9G!��n��]��4䕒��QU�s����7��C*��(�Э�ѶE@�QlWv��]�^����\�>���IC�4;�
%�z�q�h�Au*��} �V�Xn��Զ�$���W�,�A-^h̖�cwM���O�9�����M@7\��Y��+�LwU��\�H6�Vs���J���c:�V���m��������\�S���ۭ��|�콫m5(V<v��o�j3}F�	`�^���a�iܼ���ES�lA���X��Qb��ܱ2�U
W���k[�d�4Y��Q����s�a4�I��>`d�A��J�̺�b�E����h��V���#p^��L��t-2�Uu۵���aA��PV�9�F�
&C`ʏ��1a�]�/q��wZ=�
�\�:�g#@�4MKx�÷�i"ArЌ�l����k�F�m�;�9λ	��`hHA���eq�'(���3b���
���,�k��9�,�v��Ԛ��KX,G=3�[L��X|����]$�7H�*Qn_VMg��qq[)��MMto6e���f�QySyڷ�ը,h�9@�Ь�[y���d��N����n���XX�vKo#kZ���׷ײ�w��G�����-^��a�n��AG�<��;˳yO�(r-K�]��vb�Jѫ�Y���|���*�۬vؒ
�W��jዘ���j����9jx������ʀ��Q�{ݒT��CT��ƎSd'��͂Eo����h�*2޴W�y[��Yu�`%�1�iѽ���<iV�Ku�R�9���hw�Z���me�09Y0+���b5���n'ٲ�5���[h��Y��i��k:
F'̪���U����8����}Ԓ�n��[�K�60F-x��K'��)��.������t�A�����'A�*);ZpEpr�Feay����!�7Oh0MFc���:gtJ|)ԭ��Au��R:�R�/���ɍS�Z�%��!�{(TSE���9Q�˰V��S�E�f(ŧr�iw�`n�L�ܳݠ�-��r�>�P����F��!yW4�'��&|��v���:��8S����x�fA.�ukX�܍нr��b�q:�&�2�m<*���S����l�VGN�'+4�W�)���+4�b�;��%&���:κ�6�{B�,��9%y��ˣ>Mꫵt�Γ�b����$��¹���!�I�ß1٭��3V���5�� ����ZmlC���V��׻��˼д�v*�s���dO+Mh�J�;\�K���*�
�n�@t2U�'�:����t����{oO[ܢP�����Pg�% o�>O�Q}Z�����)	�k��	����zal���Qɸ`/(]�J�76R<��w]a���A,����3�$�]}�TVK2^��&T]���5�tt]؄"&l���Vc�$ܕ�޽� �Z�a����s���c�`����oZX����s��Ɵ�2�p��[v��8�m-��������-���F��]���t��V)Osv����Y%tɳ��\W�5���[	:4;����#�(Tu����O.�웃��TZ���(gk�z%L�fKE��58%�����I�P��-��.�� �۽��S��=q�ʼ�:�9��e��
Mi�DkGNo1�9���#b��|�{i>Gp��S�o7��A���<i���e=ssV�p���y;áѩ������p.�/"o���e�뮩���_K��X,T�k���������wy�B��Ag}ȁ�z\OVP5���vH�2��)�b��&,��uv1m��tsau�(��n�@Gk,-�tʊs�鵁gf�o�o%!}�1�����@��]v�+x��S|gR',��>��]-��570����J=(�v�:�D_��%NU��]�(B��m"��ި��f���֛��%oS5����X�.ޅ��!YE�l��Cz6�Ȳu\��|h��t#v$��G�>�#ݼ��D�l�?��9�jї�ž�B�jV����1�۠�ז�
3����6оc��i7���u�{���@�cxRB��@�n������^uuC�Xy6ʻ�*WL�+_e%b���ZHA!����v��7v�g23�t��@�vs���#ܕh����|Z�.G�L뻨�Fmb�3��Ç7*eN�5֝>�S�D��9@�R�9]�O@�ru�Hu�J����x.`����ۄ���9i-h*z���|,�`Z���h��+��y�cZ���5{G���®�O5-V�	3��ϡ]�%.Qj�wj��XS`96!��볯okI�euϵ KQ�qDi��B��2���:;��E�<F9�pY�� �R������a�Z�c�q���������� G0e�1gA��X�����(v[O�c�߫w���֧�cl�k�����M�x,`qr��w1cXC�;��yb��63��X&��ۆw����(=<怬5�Z�����D����T�]Z܇Y��2��TY���ɂ�9t[� 	�p�����T�3R��u��lZ�g��-E-��k�+C[Ҥ�ʵbjn\�kw\~)H��z��|p҈�s�Ʃ���+:�S��n�)�r��h<�gE*ӊv����f\�{65{�.������}W����w���b�
N��u���K�	O�-ȵ"A��Dѣ��e�"V�d��Ѭ�
�����eŶu�Ϻ���0o[�e�:��/.�i70qWe�w/}n42����^��m0�����������h�ɝK�S5o8zC��G�e�R�"����v�ef�B�l�4f��k']�l.��RSٻF;O�������Gr�����ul`k��A����Zմ/�+ �7�H���CV���a��7M��t'h�	HR+�5�/�i#6��Y{x[.MFt���ʺ���:���J�Rm2'$C۹E����1�m�})|�5ծ�^V������ٴ��&���RYp-�]]Bu]�.K��l����p��hF��Ofh�!��yk�W`wF��$5ӸV;"�s���O$ÙVf����wy�o"ʇ�-gq�/�{cy@b��D��@���pbTaׇ�1b�gb�a<��JNl�9�^����1�*Y�P�p���`I���W{Í�Wn�2���ymJ��Z�	�g+ז��<W<��]�VI��K�� �}ݵo�g��-"&�?7�I�=��1'˅���p0�2@:9.��V�����[٣S��U�OE�H[�U6��O�*
������;����j��՗�JJ7RT��e�`n5�V���o�9�攼bN�݉v�K'���^5���U�K&
�N��;�:|K�{2�,+1�)�����+��I]��]O�)2��)n�z�aũ���Im�X���ˣo�\�{/���y���Q��iZ�1��TL�z����L�^��3_�����SA�KPc嗋N�+������NfK�i�6�ּ�hWT��(��PU� =f�}\nN�"͋��flV@��e�2����)S
�-f.���uF�e�꣦�s�ج7�:G���� ����r��/���5F��XrAG{S�G�mF"�)��B��v�/� Y�a��]h��hP�k�������cU�1Xzl\٫��t�-ݼly�2��<:F���_vު����ű��\���#���՝��7�q:�(�ԥu"d��S�Uj��Հ&�Wtƫ6��Vn�K!�R�F���i��2�r���S�ȷ/b$��/5WƖy��-{؎�SV3�\��h����U']�ʬM-
�z�M��n-[q�B[�q#ƕw�ƌ�H�p�����j����9M~S�a6uz�������*l�8�m�{G ;h��q��R��v�f�T�F�j��2m�����?w;�Kb����d��B�)����/�'����ѭ짏>��i���%��MqJ��s����t��h���b����˲�M:���·_H���=B���jj�#��zCx�gr�h�W\ي��+�,���x�}`H����Qu]!W}ζ������ͧF�7�9����޾b- {+�u5�;АZ�������<6C�/syJRe��hiN��k�w�4%e�zC�LݞK:����L��<�]b@��F�R�t�hh& \�#4����搻�	&kB�x�s����PB=%>���g5��ܜfĞ`q9�|����\U��B3����4jx7Eul����i���:��]�1�i���vGghɩ�7՝���HҢ$�z��X:���`6q�6����WB�.l��;���lq�������hϳ*U�b���`a�$�E�*�6���w���W�"g4�h43 j���Q�x��	Q�z�vŦ�Xs�l��{]M��r�),��-n�]p�����+�gv�q�v7�q�5{4�8����du7��ÛkC�ܤ�k,��s��!���ݷR�[�ކ^����b�bȗC��BMJf��[OVڥ����b�����I��l��6��Kײ��i�Ԥʋr���CUNޙB�:��eY)�!�[�۽�9���K�i�0 �Z���Ag'R���ƅ����Z�7H��9լ�+z�vX�#h������7q9.�=�uD͝*��s�;��8,$oCVx�9��֏�s�C?>�p�ӈf��aq��y�q�q��L�-����
�jA`���eǽ1Է���ѧ2���o4���-
���1s|���F��n�.w���'�PF�eP�R�8#C��5�h�wvl���I�%��5�í�I̗���
5��*����:�oN}L_-����7�D�{{��,�
�d&��]M���g-h�t6��&Y�����r���_Z�B]�M�����1�b���|o��5r}Μ����\��%ԥB�[��o�0񧀮��#m�+s����� ��G��H�Ý��X��>=}��+�j�l<^J=g�����7�NQh*��\)����ˑ��63,r�,�1R��)ڮ�&����o���`��-e`�:�4����8���7�Z��|��[w�k>ln=le���! �����$�g�9���f�r���p:�՛݂���c=�10Э�!Ȫ���BYV��}�e+z�0���R{��� Q���fq�;9W͡�E�]��GE5��u����=+D����˼6�[f�A�jE��;LV�mF뢌ҤH56�N��c����Hܭ����X�U�He�0j��׬W�r�6���S7]v[�Ӭ�gh^؎u	���R����+8���	��<���DF*�^��l)��aL�f�#k��0��
�]!��6�<����+&}�ק	N��C��6��63{�Jb���A�g�m�ɣ�k���Nn+�[#����+�#�>Jk�3�8]Իe�	Rb�����l�³0ș94�t@_l[��x���������	)�Q^֝��
j=�֕u�%�ZE^����0����0���o��k�"κ}G��P��$���l��g&S)^��s+D��C̾�t}xN8�ަ�T�����j�[*���뤞VU�9L��Us��5�PENiL���-�Q�S�)��Y��	pʓ� ��}Z�n �q�}/$9��e���� ƙ��쮰:�ຐ��m��b˽�iS�i�ׅ%R�R̡�4mm������A1J�?L�ju�9�V�yl5�k9_>ӆev��ӆXĳ$g�V_u����Ӵ%3�v��PlַB�����-+/���
�/g*�����١T}�*y���Ӷ�G!aGL��ٙ��wyoC���T25��0���j��α�_�ʼV��������w��o7z�_ϑ����}J�Iõely/��oP��q�\K�WK�%���K�
�Cu�|j�QӲ�n\�j�L��%����pެ�[@ս,u�_aH7���m��̺ާX@)Z>���#��E����ݍu��ޗ����+�}4k�
�YI��b��g�M���S��۫{���[u��9�v�}�@K��	wG!���LQ�n��n�9���Q�W|ѫ��2B[�RP�$�oVZ1g(��W�����o9S�ZjV��L7�ܕ�!�\u|ƚi+��v��o䲳U	��u#�-QOr�s�{]}��I3�嵟m+���:�̰���1�����-^�J%�v�ZH��:�0*˫JA��gkv�V;{wNҨ�7��ރPƒ!8�p�&�����O��(y�"fR(�Pz��ulu�˸h�l@�哅V�`����ʷ��� ��X��H���k)�3�w�ou4��ڛI5����/��f�`�]����ZhA8�����F#T%�..��1j����&���/z��Zb !N�+�#�i���痶^�Sr��Ɋ�nM�]>���M��<�9��c�R֙zL)�Rp��#�&�Y	�]]�_[�ϡ}�j�<�������*L��x��3\u��sLJ]r2ĺ�����{�02�@��^k��J���+WM隱h9�.����/2��,-�*i��7⠐+�_e3{����\��ֽ�cU�yf��l����c,�CzU�T�����В��գ^NM3�0b�vJx��9�:a���C�9ր�563F�&�`�F�G�_f,���8@�zR7����f�Yΰbu���Y�D�C��0k��zh8u�;ҷ1��,�
}]ԥ,Y�������m�		oi}˹:�Tt���+��t���D�X0.��E�v��e���?-�M7�9�.���xk�ЇB��ZH!(��ሊS�go``�,k㶣��[�3���&�VJ�%U�+M(��Q��Twm_ �e�[)����,�Z�9�\y�+-U��K�\�f�����5q��lJ	֚Uݻ�r��%�^������.A�i|�]�tG��VHէ���Z�V�D������F�)Bک�(`��=} {j�fc�ŵ�&��[���\uVR����w�nU�i�]�%:7�c���Tk��*���vjٱ+T5���qF�ͱ�gB	-���	_nj�/��^-��V��d鷅���6�3�Q���Uɕ*j
���I��2�,�����eCN��z�a�w}��z:�-�+��l7i��E�ͺ�Kgyf�\.�����hU��U�R�o7��fnii%{��lc�Ʋ�.]�Kd���`4�V��Ļ��KYUjA]�o9p�{]J��l� �ef������:۷�Y(7X
��s�i}�f衼���RQ�1�����
R�!�x��@�.k�sv����-mv_K��J�����+�}}�kL�Κ|�p�Ee𾲨��8��E��e�V@@�o�v�%bY<ns]!���1����ڎ�[I���2\Z)ձX�Ώ�cc���ġ� W	h����$[L��]G�8�ځ�K��ZX�Y#���_]�F�Os�=�)��R벙�}1��YE�NU�GN@���y��	$p�����,�'Y��X���U�T����+�Wd�I �j���w\�(�ҰU��	XZ�_;�
�OB!�U�֌��B�=��\��m3 2���v���H�VU<g-F����6e�`��۫(Ы�eSY9�3J�Gy�!v=�΍��	ع�!��q��Ӧ�w?����k?G�P�+��3�ܾ"��c�o��7#�m�5����^���eF���H���7�Dj��=���[;l]mt�u�\������[*|���	�v���/���-%m�rΜ��Au=V��N����؈s�9�`5CHxi�b�؜��^cgy9���N�x0A9���ͧ����)oZ�D��w��������)��[�I��Zw7E��3��gZ�e-y`�Y`qQKn�a�bKn��YX���fT�x�uL���t��h�z�ǣe7�"�h�7qu{�nZ�)GF=5!}�(X�eL��t�P�ֶý�C�3P�H�]MY�]�%�+�m@�7S�cܕ��X�A�������m>�iB5yIIO��H�s{u=#�XZ�1�� `�����ڼ�63_av+�:�1cQJ_}Z�dEMR�]h7�H]gsƔ�ujd�c���˪tȊ�W5M!��6hf�4/_n���l�:��G(���QB;��������ٓl��	DM����;]/M����H����k�w.�:^�,4�"�����ab�x�+/Zx+#��t�r��V^H\�j�"�8rڶ2���Ŋn�B�7Z��a�_�!I�	O��XM�Q[�3��7�6��DA�ⶹ�<B&�%�N��赕��fr���Or�sGSw�@��&��U���M��*�nqŁ�31Pڗ/e4��-�%v��61s�2�tZP2�Q�(���i�b]��p(j3Ym�u��r�= ذ%����b�;1�^�-��f��q�X�`�E��n��31�$�������ٍ�PF`\��n�XV���uu "��Uժ�N�X�=؎tȸ@r�F�g1"ì��/M�tbwQ#�ۆ�rOz����e�Y�k� ��pl��kZko��=�t/'$�T����)�=�o��le���t�^��i��+Ց�7w��J�DNر����G;8�D��VJ�#��W��ȋ�Ft�K/��o�sv����*,�7���hS�Z���4wH�81?�&Fe�eb�%]<� 3Y��u2���APLJ�Z�i@��.v1t�$��`�k/wWmm\�<�2��(��Sa�VR�h�+M�:V����p����x�*}@(����B�V�(hױ�<��,$�u<�	Z�!Hh+7	�g��Eti�.53NT��c��Vٮ�+|1,�]�f>�:�N��X�����>�Ĺb h1�S�XBX�l�N��h�*u�т86�r�0i�G�y���TZ��wV=�M�v'u����
�6˥b�urb'ع|�t�]j��no]�J4�Ǜ�����0�^��s���1.�4(�u�B}S��l���{-�5��qf��5��0,_u���R�޶&d�|��l`�����)Q��bF�s7�؟%-]��U-ď��k��}�Ꮊ����YY:��5�K�q݌3D\Ne��D��e,}��R�7gA�kQ�Q1zh+�멲�sݪIf�OQ�M����t���0��펎�%��R�U�`ɬnu�n1�	�����c�f�/�k�-L��t]0V�����B���m��՛C���>mAx�ZS,���5�SL�B�l��	0��͗ʻJ�Ҟ�^�վ�r��Vb)178��I����4-]��Vh��M��:j���n��{B�#�
�����u��1���]+,LwB��s��ZR�	/s$��S�+
�Q*lkJ�".[fÃ��cˏ"Wn+7n�e�L=�����%�����"�;6��'&���G�׉m<�%��)�K���a�Q!�2,;�\f��a���Mm��2�m�d�Z�R�i�&�`6�e^�:<�cf�����;��oq�:V|����u]uh�[[3��h��kVzL�{���1���nB�r�����d�N�����:��E¾M!γM 4����u|{\�7��c1H3Ct_:�����Q��f�5:�`ĜZ
y1Z�9�@~���v�n��9��<+V�u¶j�S^��ʄs�S�&ڜ�	�#�i��Kuڨc��
�0�iv��گvΫ}�c��cE�V���THm���kF�i�w�n��'��bEN�Ͷb��d��81�$sq�T)�[��|4H�|J��Z���2�N�۾��VW~���յ�m&Hoz�TY6-#�\b>xZIH��aw#}�� >B�I�gz��Ӡ�&�J�!RF����d�4�͈��a̴8jeԺ���Z.��sy^Zx���!�R�|�Q��"�/��;�#'���D���
�+�,,Kkh�z����ʚ�Vr�s�9̓mn�$+*����+I}�b�}��.�vW��y�BU��[|��P��k��;ԭ�X�Wi����тT�5J%w��舻َ�ʁ�]Sy�v>�Rg+�h����z�:P��K��%��qFj�)�E5�]���o,w �Y�J��2��������n��z
T2���r�+���m�I|���V#><v�q�m��9�=+�iFu�V�Q�,�%�30<���i��Ģ)<B7ݔ��d��E�BVZKu\)��G�%YÄ9m�YA���j�5��dk�����+������"�c��J��a{>C{LIfB�`�N�I{��e�m=�8_n�ԦI��"n��-�.��A6x\ީ���Jt0i��|ZP�!�T�|Xt��m*��h1��o��"�{J�D�Xzơ�$��8�wL���B�B/�e*���
݃9�8����] �4zoZW�+���)��.1��܅Ҿ��v��-W%����#��
�8\������ٝ}�R�+�0\�ج�C����,�٬*�Ir:�sU]j���-؃�������]>���ʺlX�Ϯ��b�b`^��ԯe+/r�_Cz�et"q�5zr��|�i{q��!�r�t�KgrM�]�m��t*���u���n��1��iU8*��f�ٴ]��*u}%ꆵ=����ƯXȤ�����+k����f�wa���e�!���tYˈܥ�(�mr�c�g�Fz�Gκ胷�� Ѵ[Y�!&Tβ�a�r��'�v5tsC��iwujM&
�F%`A�۽�e���wu�;՗�(EK�Wp�����O��vw ��
�xfe�l6�bNy]V�;��f�7�Ɛ�z�sX���P��]X`��K�y��[}����ތ��d3.a9�:�G.Q˕�[ˡ5��8VU��[ �]:v��u��T]�V��Yū�+�h���wD����lWS=a��t�������˽bs7�ͳMԭ}�9�+����Z���(;Ole��Q��4�v�*,4���j�P��=g0]`�3lQ�:�+�|��R��[).q,��qKe�ًp��N�3[h.��j��:��`�W�N7l-�ͣj��0��J��j�)*�*Q���,�c *;�L�Ϋ��V��&p�xD][�%*T�wNT�I*�1G0Rj��@G):�D}��4Ix$*:��V,l��S��,<��]�V����r��-�,�aO1oeVfW-��C�Q�Q��J�H���;:U�q��4��S�u����%Ac+i &�;�-�a�N�w�Vr���������5��
��tho*�Com)�!��N��iX�w5�4Ү+fc�Y��,�a��Kv���i��L�����2�/��GUlX�3&�V��5�ܛoA�Zc���K�T�}\�N<�2*
�g�u�+6��vۡ�Sx������2մ���|P��&�t�7s��TX�t�SJ��%����m՗Z8�d-o	��O�;�BV��w*��&0K����(�+�g;z��r�s�@^ث}z[��B��VⱫ+4(����vXj:���h�	I�c�vZ��{A޴��)�(q�]Խ�Iv�U��X�>f:����/z�.'	�V�=B����8P�
�z�)b��#��r�[�
�D����e�J��)^�G��+T����A��s(�w��$vݎ"
�'Q ְ���q)h�����j���Rb1���u٬��u�ὴr�]Ha�|�TN��fkT�
��}k�-:q'�5�c��=T�%����Q�!�#�tdmT�N��ӓl�7�k�=
�<�ɵ�s������T���f���\�K)���XU�غ��t0�uY�$yx�uf9�;�}�f���f��-���.�U���QZg|���p팡C�_hXV�S�a:�ݕ݌&C���Q���t˙M��n�ZU]L����b���)t�q���[�(89�c�8a�]t��:�n#ma�[���*��wq��n��s�����#�--Icw#aO�חǹeb��:30`LKKu�H���e#�3��
[s��&�Ix2q�8d���1��t% Z�fݔ01�6|#�i�Ə�?w#�RŎ.u���]�y�mP�+ ����I�T�g��s&��(9�ż�|Ww(ɽ�8Ԝy��;���wlV�귣U�i'��ѐ�fI�Y��ڀ�ŋ�T�v��]e�uN�u$���Pޮ
��|�N���|����FuKv�S�%�s"��K�d��W+3=z�g5�<�p�y���s\�r$8�ȵbf-W�,b�8��w�W]�����H*Ǩ.|���d�}w\n���olK�C��/rm̥���;v�+��� ��{��x�˨�S�r�o��.�I{׋6%�����t�S(쮷4�(��(�����C��U�^��sf��oS�n�,�X��W{��6}��I�H0�I�W]b�[Z�������,d�*�gs��M9J��\���8�ʾ�f�S�Z�H�&e_Iéfo^�l�g�ҕ1�dY�om�����i.j��̽}A�8]��l���]�]m�P�Zzv�p����7�ֿk��ڮ�,%\����(Q���#l�,E�U�+	D�
��+iF��b�-����H�������Vڲ
"QF�Y+U��iKj��)*�k%F�T��`�2������()l
0�ѣKmIYaZ�C�U�U�(�*[@DjV�Q���ikQ�J*���Ab[
5�6�-jTrʂ�VVTl�����kPfe�5+Q���VZ�(V-`��(Ԭ.a\J���"�((�&&e�aU"����2و�e�
Q������J���q���h�E*)X���X(*����h�J26�U�fQ-���C�*�`T�QFժ�`(�̨8¡F�`ٗ9jTdY
����8%�,j����V�J�$PZ&8��1(��V��Ej�KAEĬr�&cj)H��U����Z��,%B�mJ���m���"��Q8��(�V�*,�Է0����*1k\��1��TX��bbV�ck	�?y��u�y���1�4���ʷ�R	&�l�S;���#F� Q+�� ��-�k�n0cN��[��=�-0�=��q�����E��<y9��ov�?q��\k�h�O��D�TY��M-������2���}�^�7��yS1{>��VSSʥ�5�< ֱ�w�0�x�����L/��-�[�W�<;Ԙ�����'c6�>�^��ɪ^(,z�z����q���e�8<e����<%����B��:UR��#�J����{:�+��|��k��T7�P�J�G�RY�o�x�U�+;ݭۚ���	w���rey#�ֲ���mT��Q�|�^ߢy޷B�$�M4yw��5�f���^U{�}����Ϳ�l����ڜ�Ms|��3�;�N����ݒ��oOj?.�Y��'Q<}��?9�����{�\�
�v���m-A�֝�U������k�7�s�s����uW��̳7�=���ϑ]�*��-:7�����
��˕Ӳ>~��Mz�}�U�A��ŠB-gC�:�+�+$����p��9�y��0�j�M
ќ���qﯞ:7�ͧP��%�{(ܤ��
E�p��Yj�d�[��m\|�Ǧ<P�Q�*�����o��jf�A�=:�ޭ�̶��OC؎���Ri.q��3�D����=�?nu}�_g6?	qΌ����}�i���}��^j�S��=�$��2�nXn�_"���A������emj�OLosn{R�U�s��]��buX��y���7+�t��X\C����jk��&����z�SS{��S�yT�j�����n�R�=�y��7u.�MNĩ��z������gӤ�fH�fjU��M��,n�X�GC�(X�f�\����3�O��{Q����u�/?i˭#F5˩[7���[��{��{u�;\=u[�v*���>�&]{����]�`�8vm�ץ�?�J���!Vp���y:]���s����U�r8ʡ⏢ܽ�������<nTa���+������]�E�!<�ut����{�z.���l�Oԛ�NP�7*�=
����k���un���&v� ��(Yk8b��h�D�����S�wx+#�ې]��U����Y2��G!�i�nV�Vε���_U��$gq�;LN�����/�/u6pЛ��}Ь�6n ��t]b�w0�� ��V:}m��R��93��eK�������a�Y폘[҅�8��o�iU��׫r��Mn�v�vE2�hC�&U�^-��+�D�W��by?y��@��K5��#z��FrM<��+o�����E{�qNڡ�cq��~�z>�uw��5�}}�w{�I/{�zǝ�G+�����]�߱N���f�]Y��wOk�W����#�nK�]v�(���hT�����RN��E�p����-�3x���UEΔ�̍�����7���rl)�u�Ź*��ܻ��u\��x��=���NsMݕ;Ǖ	������	Ō�v�ޗ���9n���8{Oe=��������k̆iמq�(0`QzS��ۋ�O�����k��;�[�>�3z�TRb�]Ya����2�q>=��MF���E�
����Զ{�y�N��<����e8��?6�hݺ�*����'��3�^ܗՖ��75{����E{ZM1m�2Sco(}æ�s�{��@��WJ���zT�4{wI;~K�sŖЧ���9Ce���G��3h��gD�iN�(a�����,PI��]�)��e�:���t휻wf�V�ه�>ݗ�Ӟ5}���Uoo wK��|y��C��Q��G:��j�:}��d77�jy��]z��g���]����wR��}�fkS�0��&���TͺNS�NM\�8DU]]����.���}���r�^/r�ƕW���Hw����g�LR�>�'�y��X�<�6BH�7��x/z��1�svx{�ӪI�@�T ��l��s��u�KM����7��S���R����V{�ԖumF��z� �f��rn�HL޼�-�{z��'���>ou|�����oҊ�������u&�Enz�C�-];�k�,���/{�k˽���������f�6�^{�q�յ��Ro_�f$�Mm�W�|�=��q杖�f��߸���Y�Ry� �ܚ)�{`��tP���R�\n�gF�:`~�>s�g���$n�x�q��/E�@��8�.ÁB9[������T�L�;&��[��*NZ$Cr��'t������𺆸{�^& �^�F�Z��b�� �2��mf���7ZX�i�`#�M��)�����9eƦZOz����9���T�����`\
���yޣ������Rp^saS�mΜ�4L��	r"�kJ�D���>�`���Lmz�ؾ'Z�|���c��OC�y�wK�+n�*إ��3��sc%_8�/s�+ëö*�\�u�3�}Ź�N��׼�ޗ��/:�>���j����q۝���+'\��sEOf��ER��Pcګ��m;���ۛ>��Ny��]y��I�T����t�Ӽ1+{�����t�r����J���ݎoj3ݲ�v�o��]��/ܑ� �������`ؿ|�߲<>�����d���{��NMť��Yʴ/?ly8$������s��{-[���<"U�0/�C%�}���.u��3��ǂ�W�����u��:�P�P�:�G�Y��w�~W<	jukݰ�W'�kr�Y�JLz2����x�gVm���Ʃ_�ymw���s\��ҟ�m�-l1H��F���W����6B��Π`�Zt���q�h-aw����U���k%��.��6�����E�|�e�4���4��65z{!Yeo֯�u�5�PĖk����m���ԏmV�4��7�����{�Q��.�ĥ{��}��K���;3��S�ir6Vz�̵ԉ���ׯ���^��5����1��b=�=���^�6��l��L��]��W��>Ξ��\� ���K������Q��r����Jn���w�ˣ�O��������=�(j!c�<-J7�Ҭ���/��e�ީ�e�R��΍O�w����zRٻ�����x��N�V��^�3�O�+:������9����?͎H��0�T4o����U��E����^��s�y+���:�y6�G9�l��d�_8�UB��U�`Z؀��w�)�VB�ޙ�C����ofu8��=�Q�����|X�X�ٚ}%Ot��J�+R�y���w�Nw�$�ʩ����P�ʵ�ȦV�wJ�q�ƈ{b4��o���8)8{T�cΫ�g���i'��%R5yv�F)U"��Ck��%�i.��|�gb�7Y��D�`���0<]�߳O��ʃki����N���wN��a���C���Ii�dڀ�[>㽓�,M��9G:"�;iq�W�e�V��A4]�o�=����H��9�י�冻k�B�z���0=�d�_ۯvz��Gj�	7빕j^�U;yם���7E�&檗�Df����j�]b�Y�[����]naW���s��e�|��1�t�iS��1Lg������_L>ot>�.ZO�����J�r���(]Sq��@�*�z����x�gV��/'^RV���:v���.<�_�S;�v�҆�8¯�ǣ#��3H��������z�u�~��K�R�*'D��v���u5sλ}V���
{���Z�߆]�����ߜM1���d�X�y^o�P�E{�k���l-��]�ʧ{���Ǘ�F��m��n��1V{R������g�����]�O�}�3��^�>��?H�y�7OIw>�>ПW�\o�׆�qU�u���$�M����\���J~���f��h�gW}J�����ɴ�*���C��^)[�k�	�HL��+���8e���^��X�!:9A�:�D]!Ok�b�`Yt`��r���c,���0��������}|�ݜ�M�y�T��ݍ͠��z�ڦ�nN�23�%�;���[�l�å��^^!nU�z�]�곣�=�M��4yC^�N�O]0�p�yqV�+������v���t�=<��J��oo�=��ߒ]߰z�=({�{R�(�6�J��W�G�B�el���v�t�����X�sAs��c��Ʈ��=�&�d�5�c�����K����g���a�;pz�U���s��E=�����qu�L�}/)�<k���/z��V@�ς ��1ܓ��W��f���yy�{R���T�8F�v���'��<»������=K{���pn�d�f�/����rj3�p����Ƣ~�_�w���yy��C�-U�x��K�����HT����B����	�~Ί�~䔏�F�Ǉ�|z���Q����Ig��T�U�ǽ���K�&���Ǿ��,k�~n�UF^mO �խ��~����g��Yյ��|Kl�10���L��Ϫ�(�<�k/,ze�/h�c���T:uG�ex�V��O��^a:��j��S[���{�����ZNQ��11�*:�8�jc4��.��6��\7d��-�7hA��8�p0�=���(7�u�ʚ�,�ΎD_e���������i��u�خr^����ҏ�?E����lh>�b�WwF|ӳ�R�����?u�y�[���K��B���5��y���ǋ\ܾ�������f>�s�Ǿ�'n[��S�+��e�=]�Bq�͋���r���*�y�sa����q���z=n���,�[9t�v�l����#��D�2���ÿ́��rx���nv�=Y�,��^��2��'"��2�mxM`k�\�UE��k���Q��z�W�==ü�;���)˪?y���=Puz�lF��.�FvOջ������n�ܭ|��;Qn�g�i};ũ��������=Y���+�j��w5�psc����'?w���*�rT�M�^�8=�+v�-�H�ջ�d��w���qk��7�9�IU�ڏ�ݲ�5=
��]��j��N�k�ׯk�� �w-�~�M�w|n���M�B�v�I���'�dK��1��k}�������J�MfE|�2�VYQ֥ ��
������m��u�u��YX]i.��k���Y�ΔZ�7�ыz[�Vɹ����`�l�U����Pz�u��N�m�H/i���7V�mlN���r�x�>��k��{-U�����%^����߰�O4Xk
��s+��P���mOV��=^E�kb��ˋ��n�J������.�W�np�kٽͧ���J^���ғ��Ǯn+U]<}3�6���U[�WT���=7���b�V�����ޔ.�aT��s�/%.Af�*W^c�������v���oWz>_S��*�S�s�v����adɻ����A��x���i������-��R��'.�[��zJ__��<�cq��;���{ͅMߧzo�x޽����sJ�\FxZtj�:Y����6�X{rmM앶��߽����o�UO�⣖�Q;U�7�Y͋��n������Mo���Y�����M���1�F[UD�Ur�W�!���o�P
�sX���X�9�R��\�֯��<-���g�\�Du7�fl[]g MFO[��p�a��3���,E���t���@��Le�\��I�*���/
Յo3�J�w��PI�G~���\�H�. J���FGP-�^,�dk�_n���@3x�8JRVA+���HG[�S������ �}�\/̼�M�oL�]�ɺ�sZ+��gm^�[�
�tey%�oM��Wq8Η��Ţ���Q#��㧾y�.�\�E<r�x��B��m�q��ۛ���樌O��Μ���0=h�u�ҍ`�Y�2��L�Y��ӝ�KY֮�RNg���H��w��D:��0ej�$����!f�c0֢���c�x��a.Ȃ1����0\�}8fr��w+�s�/:�W'x�+*1͕�:�H�wE%Ի�K�Rh�����S/���R^]��{E٥�� ��]��坭�u5ڣ��Vݧ6�<x�RX ���}�|��5pXU7�����M��gY(s㛺aJCÜ�L4�u]t�y]��u�"�m�Y�Q����T�1gp�alVXGN���6�[��7+���ťB橝F�t�)��w���q�^[�C���]�력3�wq�Ӊ���c4Yg-aI�ia��{F��WS�6�	�F���.�nm�慢����.'�m�*w:`��i�����4⤛[Gt�g��ʺ	�Ro!ڍ�5�IiuУM3WKn�8����aSj�=�[(_FQ���tP�����6k�p��y���Ao�G���q]�n�p=�g`�Kw����Ƶ�ދM]����Js�O���fiv�d��@]��"ҫk;����ћ�l�2��n�p(�eM<T����F�U�v1)լ�C6�)g1{JRٗn�^X�S�={��5[�_;��͏Z�[�{wQݫ,X�$���R΄�� ��xluG�� ����T*���#Vs;J�Jn_��RN��S�G;o �s�����
�6.�Ϟ���	C��Ic�c���@�Ѳ�.�'���8S^@�ٕo\͑���\:�eI�������/������8V���N�{Yiu�N+hN�Y-ڭ�s��m�	udyKr]�;87�>��aTa�q-M�!�A��9G�9��c� �m����4bquj������H�Ř�R뫙ћ�r�z�3
�����d*sޜA��t;u�;����:�����v��� ro'}b���|3���`n�=��<����P˙�p98�l6��c�$���9��ƹ�ܖ�r�ʈ�:`�D�
��l��"Sfb��*�ǵ��SD\�A���.��k
pf+L���^��L�� 췇��x�h�`��mV�'�1s����|r�왓�Γ\I%Y�W+��b�@P"�(�)
�cFD�m��c��$UD��[b��,`�X����fP�YT�(����+
�f6��`+R�"*�R�EmYPm���r�(��V"���1�"��6�D`��iR��kV����*�eEJ���**�ʂ�J��7b9i1��J�����b�V���(��*��Z6���%E
�Zc*
���ܡ��VKksa�F*[�+��11P��kUER�E*��4Qƥ�Dr�E\j12�IZ��[V�[�Ũ(�
��m+�f&*�TD�,*Q�Z����Us. �"�Eb"� �Pm�U�H(b-��0D�"�UV)*W.eF(�!DU0�Q�����fR�*�(()DG(fX �X�TH�DH��"TF1![�c�((�P��U"��P��Ub�e�F#�X)��Q�2�YQ1��-�P��~�����uz�'+2��ց�uĸ/OG�U�3Q}K����A�2���iEue�0]�N=Ǻ����J�o?�ꪮ��p�[��L{7���n9�����;s��B��QT����Q���s;����[�x��OC��֚���S�)�<�j4��m��S����`(]J�5��u�vg���Rs�rL������/�z27���8gWz�B��-s~�϶_ekKX�(�����MfLH��խ3\����\U?9�/��e�Z�{y���[�v�ү]:���ר/fJ���NMR�g��7{-gL��뱳:�Tg�Z���y�٪���@��H�J@����ϙ�"���=�.�{�Z�ǚ�SI�ܾs1�{��s�m�J@�*�z��j�x�
��.��E�؜��"����|s���S+�q}�4*ޔ.��$O�1�7>����'�4��<�:�*�'�7����_�'Ҽ��1���"��gbl��L����|K���GZ�i�Z�9S�۞��A�czKy���桷D�(�܂��Vè���4�+]2Sٕԡ)��n��r�Bd�g��@��:�uGhj|�N��9꾩8^ˁ��ґ����w�v��0Bx.̹)V>QoQڑ��y?}UT�9��ޮ��I��6r�iy<͔V�+[�ϵgQ^꘧*�����ѭq �	^�%gͭ��%%n�y��R�7��+��zן�]�w���'�{5��s�q���~�l^3���r�d��Qy{7Ӯ�<[R������|\�'�)��97K�����u=��;ޏs�n�[��UV�])�:<ߞ�t�l��9�f���g޹w��if=R>�{2�]!�(zp�W/�|/�}�w�������b�\��)z��F��;&�W�1�t;b�\�u�gb��}�S�=��4�s�瓒;mݮ����K��SQ��8]���E����f�Ԝ�Ǚ]���ܽ�1����|������D�^Ss{��t^���X�m�y��e]��~��g5�u6M�;����EՕ��^TT�zƊ��<�}�\�X���E[�x�k��"�Y�w�y�TW�Y�w�2I��7����x�~u�P~��P��(�k<���vz��X�i(��@�ҝT�`�H��5��%)�x1�K��s�Zo�|1��r�36`G$����j�ާ�1
�]�6������������zyz�b���=�uM<7ނmS읟3n�9Oi95Q�����КZ�f���E�ȴ{�eQ��}�ؼ�fD��`]{�*�N���_J�����=˩+J��w�e�k�l�T��۾<R�m7�nu_i�<���9�����'<mG�2�֯�N��e��κ����}i��ǟ{���i#�aOT�mv���[���^G���z�����mJ+>�}��%_��;��%;��� �O7Աt��?u�w��o7��򙚞>*ɒ���D���lP�\�S�.�H;��1����z8��);r߼2�n�A)�jvneonp�r���+�;DN�U앜����(9=�M����}KP����SZ��,��h�f׿��(}��(�y� ��u�u�����i8�ĩ��!Y8�G9�]�N����k8��^>Ĝ����'4�V�����x�i??2o�&�M��̓q!�a�VO�XjZC�|���.2O��y���&�É6����2u���s����V���h��L��L�	�I�]b�c������/a�o,�>�'*tw�!�k�y���V�?l>O8��g&'�����,C�1�m�k<mQ����Y ���Yy��瓔�����_K浒�ub�׬$�������I=��s|�9�>�Y��@���p��	�O������ń�m����Dē�yϼԘ�l���P��A`�6�̝Oa��m��(m4�6�Ϳw����7ϯ<��o;Y>��v{�2m�o�zwyl��w�6��'uO�|��ɳ��N'����&0�C�y�1	�t��h,4�ğ2m>5��N������߻�������8Ì�=�ƲOSA�9��y��N$��Nk |��N��I�M�{�rN���a��l�O�w��:��~�Rb
�}�b���0y�7��������{�%I�T��@�M�q(�m��{�5�u4ya�J��}��@�O]��sY�~�:��P?C}�8�2m�������>�{�D/����|���l�~�ﾂ���������J�l���N�|ɷN0�@�=?P��&�h�RW�C��	S�>9�?$�I��32q��=� �߷�J�9���~���C���|�̞o_�x�:��3�I�RM}x��o����N2|��O��8��k�XN0��RW��!��%J���Iy*��mlr�����B��}c��
�4�8���y��q��w��I������'X~��ړ̓���&�X)8ɴ��S�`u>򇏩?$�O?o߿@�J���_�����ղ2�/�UAZ>������$��k�a�IS\�d����N$���?2w�0�	�M�����I���E'������V��V��=���w3�q��}J���!R��'�6��,SL�A|��I�C����IS_��Y8�	���N$���� |��'���[I1������i�hO�k������_Eg�||BU��	�m��m	�z�d����'�i��/��	?!�<��u<d����0�'�?v�u��i>;́�&�;~=��~?�����xA1�J��:�(z�n����)����H�Y��z�bF���A�j�K�{\\��1s��)��l���̹X�Յ�z}q�E�k
<ń��]���ڶj1aj�g�So�����{�P�}�r9ά��ǄW�}US�1���#;��&�����m�	��Ȥ��&�ܳ��Ԭ����.��'Y<�d��u�׸i8��o'�I����ã���|��g���$��nɣ���R}�M�I�>�2|����}�O�~�|�Ozʄ�1��Y�I��7� �L5�Y8����M��N����`N
������Y������ߞ�yc?�o�U��O�O�i�&��'g{�:�猚퓨��ٮ{�OX(m��L?!�YɦN'�Ld�!��T8��3_`A�߅�P�?z��Ok#��m��̯�'�eN��HVO�h�0봓�?�:���'�9�=v���rN��O��I�:�P������,��N'���}���
�W�Ag
�|����}_'�I��8ɴ��8������}���9��~a4���'Rm�	��i=v����c$�l�|Ԙ��gP��Aa���u���_���_����4�ĩXO�8�5a��$��P�&�̇��6���9����a�~ϝ��d�s�:��i=I����N'��ߺ�2M������r~�3�W�^��B�
��Y��VM���hI�N2�&�u=<��i��<�2u��y7�d�O]��5�>@�;��ēL�Mw	�u�����߃�T����P�����u����N=��I�;��& �=ݜB�m+%@�O�m��a8�����mI8�|���!�هI�=9�!�	�|}���9�������i�)��B�b��w]}�>�a��P�CL�N���d�CÝ�RbVi��iY=�|ɽSN2|��������i+�!}{���w��E�?ot���_���W�}_�]x}P}'�i��>@�l*��>�rC�|���a:��̓��^0��?�<2��O�;�xj�q�l��|��Ͽ?��ۧ^@_�<��T�:�GI�}�;��^�%{%�PG�"���赵یvP'��W���`�k	8�*��嫤�C����Z�q\���z�Y"��_*�8�_�ZW�Yr�ٻ��t��W�/Ц�:���rʒ�͵�wu�ڄ�=|y����n&�yM�J��?9'�~a���M0����d�+�a�I��nM$�
Cý�T8��9�AI�'�����IԜ�d�����|�1�U^[1�7럻^����s�>��|�;�hf���ԓ�y��u��<=�:�*V=�Ad��s�:��)��T8��Vy�*ORh�jx�i����#��{�}����Z��d�I'�}�)8�@�Xq����S��N2�z�d�'~��=f�:���:�|�a��xu�T��a�N%d<;����D}W9�?z�l�'kR����"�:~���I1���=Ԙ��i<7dR~}`h�8������a��򞦙:��?{d�2q�^��a���۪���wTԩ��*�����r_r��g��M%d:{��d��'�9�6ɶO���$�O!�}�>t�i6Ȥ��&��e�d��Mya�a5�=f�q
���_��AT/��ݗz���k������&�|�s�=g�'�?s�q+!��p�'Y6���9�>d�'���~�'�~�|�I������2x�e�d��E�ꂨ
��ࠡ�N��㋹���x�`$�
��Cl�JΆ���I�.��i�����'XO�{�@�N?$��'X$��k����(q+&�����W��}��Y�{ �E�^����L�k�l'�Vt�PRL5x�8����I�d�Vy�p'u�N��:���ì�}a?Ozd$��Oӝ�:��_p�)��}P}�[����~û�+��sZ��m+&�q�2��2|�e1$�g�T:��mזd�V�Rm�Y8���d�d�9�'~�N��/0�M�I;�`u'��ϵ�w~y��N��k��[�2���Ld�'}��I�:�yhm�&�Xh�������e1��N'�T:�$�|�2m+_�q�l�}C�>�
�����;I4�󧟿}�w��O����4{k�Ds�����A�ڵκ�N\�0�����|�M����c�3
	I��ɒ�MV'}�R`�.~Ot��er���C=aC>�l>}LΧlո�ܴ=B�#��c5���lrاa���U�	;���q������}�Ui�mY�ӂ�~;{^ݽ��<�������s�I�xs�5& �4nΡRm&�`m�:�I��MyCl�	�T:ɷć����m�}��n������������ٚ�0>a����I;�2N�Y?$���i����CN��߼Ԙ��ѻ8�d�VMe�>d�y0�|�}�V����A��~ѫF�/߷e{��N��z���l�i??!̰=`~a�ߞ2~a�a�rN���I��w��2xw_�
I�<�}Ԙ���ԕ�hG�UP}Z>��=6V�_������ީ���I<d�w��$��(m%}d4}�M�:��h{�a�'Y'?v�N������u�$�?�uY;�`,'Z��*�����TA����.{���O��dĬ��OY6��I�&�>M�>��C��8��!5�q���7���M���i��)v�C�=Ag���_~��|��qT}��K���f?զI�'}��&2���"ɷ�����=t��m���?�N!���&�~�x�VT8{��a�ý��N �;�������{�����7����v2m*��H,=d����x�:��3����I��M� |a��~}Oڲ`~MP��'�I��c'X{��	�+L����FZ|���kםn���T}*w��z�������'>J��w�B����y�2M2{���3�$�ĊO�Ka��~}LCI8�{�=M2u�{߹sg1����뮞{߻o[�������~�OP����è,'����:������'�d�+�;�|��'���d�����D��I��E'��Ka�G߅3��j94q~�绿�_��TWߺ�M2q���P�N���	?!�No����s�:������:���Mr���>�}��O����&�$�P����sV~�C���Oڿ+�9b(�[�]��[siPho����a��u[�N�YP�1`4��s%h�� �4��:-博��pp��|r-��/���ƭu��\��_d}۵n�r� ��tw��nn�e����J�̢������/�ʪ��ﾸ�����~��&�8��(u$�*h�ì8�h�xd�'���q��S�^�&�q��7��I��ݝd���Ì�d��O|�I��|�׏�k[�F�y�w����]ﰛ`v��z�'�=C��!�i��xe�a6�Mya��_P�'PP=?Xm'8�<��	�ayN������\=�����W�~�1�Ty����������4����4ɤ�;d׶N0>I��5��DĜH,6��l?!Y�Ĝg�\d�!�O5a�n���N��5��i8�ĩ�l�d���Ϝ�����u��7���m��2Ov���6���߲�u'��;�'N3�;�Rc�<-��Y>Aa���P�'�\d�!��VM2M�aěe`g�������}����w���y���Cl�d��~ݐ�C�����	�Os�����qa8�d��ߴLI>g���jLa�C�N�Y6��Hm�:��Y&�q�����ﻭwS��y��������s�t>O'�Xq�������':����@��y�p��L�|��<d������N'��w~��q���&�N!Y6����s��w�}矍����������4���I��G�8�I��ya�'=����I��Y�P��oz�h퓩�O�i7��	�x�����N�����q�v@g���F�����P_~�ǅ}Rm�&���������3G�:�I���+�!���8�ԟ;a�5�>a7�9ru���~�rN'��Af�Q~�.�����U}��
�חT�}�9��&%I:�IRm��YI�O�6��5a8��k�Z�m��(u%}d5��8�T�n�$�I�_����B{����|����M��k:m�L=@���
��>Ag���:�̞��2N����RbT�G׉+&�X'>d��P�`m5����'~Cԕ�&��4z�Tܧ�	���E����(v��c��Ϯs��Rs��FL��+���@;&��U������N��;��hQ�����}۶��;�����k]j���f��Տ�S�0�H������7[����XQUX��mg@�^�&�����و�v��Q��P���L��}_}U����~��sy��3_ݲJ���S�M���r�d��;܅C�� �ü�'�����2N���ړ̓���,��`je'6���~5Bq���������w�yr��y���߹��I��I�v��M�����IYP�t�$���0�'X{��'|ʇyHT��>�ߴx�i����I������E'��k�s����w[��u˟��|��6�Ր�!��zβxé?n��4��������<>�Ad�4~�d�T'�{��N$���}�2|���}��L@�i����˽<���7��{�{�1�	���"������	�q�!��BzyOY�N��O���4���{�����N����~��u��P�~�O�:��Ԛ�|y��v��7t�����^�~����z��5�����T���L&���Ȥ����,�$�+<C�8��˴4��O'�'�u��/��m'�7���$�ǝ�~�̳uφL�Q?�2�7�W�\>�>��w]A��d�Ԟ�܁�'�>��$�����'�$�'��2��4���2�2OYSG�8��3_`u��,�OԛIĝeG��e�Xw������\�ꯘ��}_�*�P}S����q������N���&�d��=w�{�OX(m��L?!�YɦN'�Ld�!��T8��3[?s��9��v�������u�ֺ2m+Ԟ��'̩�{���4w�u�I��̝I���ߜ�Ğ�d�s�'XN��;�RbN�<�>ed���VP�N&����r����k�w��s���<�J�4����i�z��6ɴ��6������}���4s�~a4���'Rm�	���@�O]�~;�ud�NwY&$�C�{��g-�=�߻��c����d���d�<�La>I��VM2M�C��2Zd�'P�s쐬�a����i&�<�u'��z���;��O;uߜ��۬ٯ�5�i�,י���+�ջ�E�T�#��aQ�wg68)Rndţ+l���yY��Z5��p�-���ouN����˒��Lf<���;��<H���Z�����������)��hB�I[���ވ��ެqt�{ �7�)*��wb�E��,�}U�}_}O�������C&���~h����l��h,4Z|���m'^Xm4�q�C�N��7�d�O]�̤=@���߿[W�!�ҧ�}����R��};��u�x�6�O}���O<���u��	�(M��VO��l�|�l���q���,6ԓ�ז$�������¾�b�v�?�;��n~��n� ��	�O�Y<I�wI�i��vs��2x���qw��Ĭ&�N���Jɨe�>dީ�'>OO�����������/=�z`��&�l�عv����}�I��X~a�I�ݸi��>@���*d��Nw$:�̞���u'�3��ĩ&��aY>|*�*��A��>��4og���0�����Zx�	�&��l��I�<�aĕ�'�<���$�Xh����N~�ɤ�AHw�2z��v�R~Iý���Iԟ�����(����ޝ3iS��%��Ok�����Lv�ܲz�ğ���P�@�<f�RN!��`~gY<C���IR�����$��̝I����B��O���~�_Q���=�����/I��xV]����N���I��'_�,�O���Xu����S�d=�=N�x��6���d�CgXO��<>�Ad�4~�~��;Բ�9/�iǊO߷����_�n�(X� �V}|O�Voj�uo؏�^�ɓ S�p�~�K+ҽ��ǻ�;�E�'���ݪ�}��Y���.�'�x�����'6���9k���Owr���X��Sݡ��~��{~&�O�4�
8p_Q������p#Bw
�r���A��WM�2�v��+a1Ԩf��=�W]�.С�C�XԴe0ө�tڱ`�Y�[`Y�8q7x�XŊr��W��#L>�b�<읦�	)ų��4�ie�+��1���.��M �Q��J/����_e.��bN��߃��/����6*�K�|�.d���Ƚז�w�8[�R�Y��h�A��7���br����ZF�#ϻ	�y�{`#�$���Ȯ��]�WWo�y�Y�n��N6�K��E'|ݲ-�����Id��1��-�Y���c�\��0\��:�x�i�O%�_lZ���cSXz+�8�]�)���hwg,Ά�2��͇9��[�噭j��
J5�_������+m���ԫ�6Ȏ�Lֵ^�۸�K�0@	��Ŧ�x���f����@��$2�Ui͖v�n6���]�&��K)��*�%���.����O���=;�x�����'r�v3ofL�k�xq�K&
��Km���l���1�dU�qZ�u�S��״;z�r�aS�r0��y�e��D�}B�0��gi��ی;4��+��)�jt��Ju�,�ŏg%��9�c�1�;�I��W��*�١��W�I��Ǩm�>���aY3l�d5�i��i;���T�㬧)��f�RC�ʘ>���|�7z��LY6u[à���Zi�,V��3�Ϸ��W4
K˭���v��S���*0���ogM�7:2"�Q���M��6Dy�4y^��ĩ���kI�6��1�zRN��u]X�l`��P��y���]v�b�����r28vb�[c-r5��N�@�Ѿ�V����[�u�/]ho,z��za�+��;�P�[%��\�3r-嗰�D` ���G)�.=q]N�������3�8�r��lfP'-�-��/�|f�B&7���m)tw�r˧�/�
�����Xo�t�b�˭0����' 0ww*����
�&5٘36���S]>��3V�*=�	ˤ�i'/P�|��� )Q�Qהz��V�Q�m�)Β��W��wT	�L���v�+�̽�(���ݻ�e̥W��]95,��U}mh�K�X�߅3�R��2�v��Ցm����"Ķ�Q�(�]��=�������Ȳ��8�0SU�Mtڝ�ju�1�.ݾr�P�������z|)h�c.����4N��W$Ņw��j�ojI����/��Z����;�׳���HMs0wX!���+7u��	o��a���T�Dt�����'իŝ}��w׶�ۮQ��\zU�$;�)Ce[A
����x<TsM��<�)�SG)i[���>���|���;y+�Q�(��j��z�ťtW����\��kv�B\ʋW+m�&�l����vt��j4]3n�p��p������7��7���&�m
>)��h�����ZU��ԩ��A�(̷)Z�e�kk`� F�T��V��R�*�2����
S��Yb��Z�0ee`QD[lm�"�1ȌdP��R��Uej8��+"V�L�,��X�@c�5�Ģ��ł����1A�娥��qQDH"�J*��q2�����,���J(��C)j9L")r�R�mRe�-.2�)��G-
c��r��.P�er�Z��lV12ʍk�*[EUEE��R�1%�QQX�[�
�DbE�Ve�B��#F���1�j".Yr���m�m�����(�P��,�"����-�a��\�@�\h�[dk*�@��Z��3Qr�S2�$m�aE6؂�e�0b�)/��H���>+B�fM��Vu �����7}�ulCy-�z���{���sh��Þ�Hu�I��:�)�]�e�*�ƥɡ�.Y:�g�_}�W��X��o�<[_ǔ�Y�U���n�v9{�Rn�U�y6/3���y�c�	w:{�n�tݹFx]'F�y���?8��'��)�����ٶ�5My���Q�C�l����*'b��u�|/����=�y6e9�G=�4�;�=��u��`���FW�P�h�k�Ⱦ�c�xwsh;��T�����	z�y{�8)�u=F���:�s\_���[��۵�J�j��3s���p��r��S��E&(���j5u�p���_�����t�o���k���l~_C'���|����)^TȕT���J��[!��V|��Q���z�@s�^˪�9p��vM�To�nnS�ueE<�^Ta��תJ�lo�I�6_3C?b�9�S}i�]~��}pέ�W:|���W��e%��[�\����(~�kmek7'���ڢ}�u�S�3����Ӹ��X�{R�_�5ޡ��SZ(�xf�E��i��m�����+�ʝ�L�tFq6�ẕh�*�~!N;][��k ���+x⣄�}��uqal���D2�y;WD���@��a[��t��Pq>�༒v�ٝW���UW�UUtg����?{�����⛯]T��3��ʇ(t(���Dy3=z�{������Z�	��/$t����z����y�]E�_�F�z#�����Ws�Qt/�M��}�}{J������*�Ƕ{������?�QT��PV����Oc��i������Y��_����Oc
�y��~�K��m��z��.��.���J��N..�8:���;^��{��=V���&�����ޥ��g/cK��(z�3���^�^��ªz�����kUo�f��-ͩ�ҵ��O=��m�[�hp�#�`l���83���i�2Jz�N'�ƥ۲��������+Fׄ޻|��&yբ����1�+���v�&�o�h�;o~nsʜMGw��wݳ���j뗻=-��J��y߃k�c���{���y��Jw�_MF����{b���n����D�Mo���ꛛ����ӷic�]�wcv���sX�x��Ov<,z���p���A�7��})w���U�]�淬B�X".�I7Sf�����2��&d���5r 5=�3�z�՘�n����?W�W�}_�� (�u��7���T�K��ʸ��󽊤����Eו3���fL��>��<s��Y�N{�j�A�=�{uJt�y�����{�M�[�͗��S�M���gUoY
���{55إ�u%ގ�?���u�g���]�,̞77*1{K�&���e3�/�c���[����_z��� �;^�������{���R'J@��c�&)�L�ɝ]�E�y�����!@��G�S��l�'��3wx���]7*���z������0'���7����%�����+ބuD}�z��c�)1�Λ�?aɲ�o�}�e�+r��Y��V}|�����g�Sέ�{���]�ٙ�^	1���gޮ�;$M?}[T��f�>��7ݛ3��z�}��m{Mmw���x���w�6�^�k�}Jn�~�����}q�t��c�=J�~�wD�MK�9cѝM�խ5�(�Jm���2j���S�}.=����%Y9w$���qA�qۤ������o�v�u��­\�g�Eם�b�ٷ�Z�:cX�bp����� ���o :�����oNE6�#��T��卑JA���iN�07�+�t��_}�W�Q�=֣��3y�<��qJ��G5��I�^g�����v_��$�lvk�����[S�'�}�����t���T����*3��p�+35g��I��;���r�Ⱦ�q|gΏ�C�n9���N��')��{���M���[�:����O"��k�����?�|�+�������roz!��:�{|y}SQ�c��캜�gm�w(��,&�vK������K��%�*��/)��OT����p���f��֗��Z`�0}��L����O��*f/etk�>y3)�s����9���c`g{{%E�މj��R�=y�Þ���y{\�����D��jZX���R\�o}��"���-��]N���t�!�J@����}&)ɏ@7 n�WO9!X�|G�z�Y��.j^k2%^����7mH�7m<͓.�LT�H�Z��ͯ8�:i���5�#o���7�u|���kj6��.��!a;��q�R�;[&�����l�	��+;���ٓhF%f�y���.�� ��eN�Ӿ�k^��'66wӫBZL�ks:���4-O���_}U&��/g�q�'s?w �)��P�_b���Q�޹�6��֮�
�ow��3&_�1��.��/zͧ�-��>N׺U��dv��\���Cc����-f�z�zFOc��9&��iy<͔V�W���<�爫��ut���ڟ_�*=cq�<�o���suV晞��dW\y�8i��!�W��z@���s��:?H�yғ2R�1<���"R��<��>.+*�\͎~q|\�'��ҹEY��������&��ܗ��ՍT8w����ew��gG��<�$�P� ���j�d�\��v�h�p�}��q�����j����X�z�:W���5��|7�x�s��V�J^{k��p=��{\�VT��Ϯ?h��d��$�@���n6'-���{�rN觹��)1E���MF���E�0�׏ok�Gf�°+GYY��"��!��un�G	�	˾�^�i��x=ћ���}J�J�s+��	q~z+�d�)�]ǳ��i�G�`&�T��6�6��ʴ�0e�J�_酜��lM����c%m�\�,��s�����e�]�t8��?U}��}���C�߱mwR�Y[ܗ�ާ{��Ow�H��
��sƴ���OrNz� o/�BN�����>�k)���w��77)Ⱥ���!��{�e
�o�Qunp�G�y��w|��9�P�ۯy��d�f�,x��h���Sq���imz^c����#����{-?��TwΡ��]v)��:��"+9?w�H�$z���R�}ҽ"��p�ή����e�����������[#-5����t*�(^8�}&=Q�M[~��>�N�n�N�P��{��$�C-ꇺ8���}���~K=[Q��=K~]��<��y��\�cu�^��!Yľw����>���E�����G]~Ʃ�^ϼ�
����'�޺緌��7�x�����j�y#<-Ik�Ҭ�}~��Y��ߞ�I ��z�k|��q�7w�>[;K���+�G�|/�N�씲w_>� �+k�fPLT���(��'�Q������B��_^:��][�QX��c���.���o850�*p�"�@���%Xʌ��^��TE8%���W�ϕl�+w2V������*T�E ծD:����G��[M�6v�m��q�;.d�W��}Rg��=�w)����U��y�|�ތ�!�.Agi;��p ���]ޣ#�gG�/<wx���nt��{��6"3�CF�5�u�G�^mܚ�]��eOɸ��\�ʧ��S��M�y��*��U=G���Gǟ�b�;rWn��>5�'pN\�'tS��T[���S�YՕ����O��:���4�ڃ��]-pwKg�7���b����E׿M�R�����������57Ư�{��ۥ���[�o{�{��J��KwM����ls��^ϷZ��jyW��s�t<f����<:�A�30;�p|����͊
YY��_fZ��=�1�{��NMR�L���v��ٹӹ�v��z����4ێ"��O0׽ ��
��:U {J�1�1FS~��%��������Z��î}}�O{�V���y��T��dc�7�CU��aq*�mV]����diy:P�%�]�W�$�J�+Q�ݹ�rW0o�[c�6`?�U����%�Q.Aݺ>�z`��kΕwv/���.�q���I����,&.�^�떩-d����cb�+y�y�s;QT7ٝ�u��o-��n�?���諸"׺BE�~�]��>�e[7�Wz�v��Ja}&=�n��ŏԻޙ�7��٘�ɦ5r6����O{+V{���k���]t��W�[>�������3_����'*��g��34ћ�W���:�^�x�Rg��x��Nwc���������5Ǿ�7w*=չ�{���O��U�{�@�w6tkoI�J�w�*��.h���9�����>��[0��5��{yr�x���G��Yф�%�:e����H��0��~���+��M�0���n�UD�a�Q|.���|�;�y6���{+�j�t��鑋����n��v{Q��V;b��j��ؾ�c�����9��,�wfWN����6#�z%U;ǦٯW1�a�F���j����vEW8&9M�^y��y��e=��֭ɗ�5*���5|����qp{WOs+�;��z
9��1C(R���/Q�<�-���;ЍuX��wp�	yc'f�(���N"$W*x�m�ܮ�<�S�D��������Sdnq�cc����7��]��3(&�ϢWH�8J`�rlz���zΫ;��׶���8�������:y���{�I~C�E^���1{:5׏"UFe7�8�i�V��D�zN�|�ݞ�/�֕Sq�]�T77>p^�rj�^TL���EǙDY��]���`,{��}V/5�jU�0/��}�U {J�����3� )�U*����;����E�:�W�W�_��"_{��s�7���u�a]��r�o't	�\˻$>���Z~�g�/�_x��[�}�PU��L�#8��]X��U�oJ��ʖ��<�I��dR���HO�{Jr����w���]~�W#�
*q�����eg�fP���ꩾLwmU�ÇC���m��KOj���S[�w���n�㽹�9�ؚ�Ī֓�ᢥu_�s9��̯y��<��k.�ӣEi3�x$8�e[�0��wM��Aq�//����p��ע ��<�k)���}T p�*KѪC�X&����pz-�+E^Vqʸ�2��u�H�;���5S�rm�5;�5ǼO���4b�{��f���;�����-qƶ)`�;s�Q�S���S[sF�5�l̎�Xx������2�AڲK��_|f�Q4n��i�Ԃ�fo��m�;Eg@/�r%4Bc{H=m9�Ŏ1et�4Xڛ܉��F���҄�tXۥ�lk���]v��W����꯶k�&�����{��MA����l�^��Z�u��8*�l�^w�N�!�N.�hv���<�N�^ߨ7��ǔ��=VUK@��}@��"���W|K��#=t�:죾�6>�Ժ�7+^©�x�F��8-�ϧ{,p��P�ݎ�{�R��/�0�x0�܄���MO�_�<s��2���?���d˂�eL��9�J�r���<LB����e1u�\�#����	�C§Ԙ���~��p=�ߚ�K�=����.aȽJ���)%5G1{<.󺬣�ʇ��Dq'�����޺���z��7��y@�
Pw��Q�v�7+��*IG=y��V���R�yJ�*��iV�|Ig�[T��XX�WV�K�_�m��J��{*��3�.n��W���W�F �W|�U鴶ˤ{N4�xg�1�K6)���:�o5]��{-s�ef��c)��ޓ��^ d�joX�Z��{oԋ�V��t9`)d��zb�]�G��݊��ޔ���9��P�XӕQ��v1^���Ϳ��^q�|������]$�l��k�]��([u�!�T�l�X*oZ�p-�N����Gk�C{��!yRl4��iu_mNwAާ]�m����nCQ�j�r˾�L�SE�b]u���CI�r���+)��5ejYՐV���L*���1*�.ݐ�#OO3�:�I4��VVy;���sv�=V�E$����%a�*c+k1�v1o;C��x�*w5��Z��I#F�R��dU{L�v���5� �X�M�u�u�p�J Mbջ����:,d�Ϋ�9z�(*Te�vr��4%���@�^v�YE��^��y��<�wh����A@��Uѻ��C��XL�]mMD^䥹�e�;���p���q��w<9A���l��_c���@�Y�����V��t����"-�$:�Į��ɩ.�O�X�����#��c`����̷8��5�uA��j��^IH�Rl�.�tK�lu�S�u�-Q�+���A�㑀��Wm��3����݅��|/ꓪT�ͮ���N^F8��3l�
��78em-�P�"�[�gj�6�9E��e*��bt�y��N��^��4򡫲�|��cn��B�:�>�|�:L���Taj��i��Nc�X���l-��hweZ�㡑�4»�'B]5�5�;2���tn�о�Vc��\���ʧY�A�.1���x�;d��N��;Z1�v�2�ݤ�7U��:���N(-��0ӭ���s�y��sz&�K:(��'t��p�tC݇���)�+���mc9����**��w5үD[ꝷ윻�E�u4�Ϋc�@2As�^r�l�� ^;��Jϰ�*����O�4��#6����df#R[�u��a���!�^#ox����n�)�����ʉ�
�an`C5cZh0\�,������2���ι�S�4����} �^\�l.*"uu�G����ak�ު����.F
�5�d�G�w
1�>$�P�je;��F�u�њm2��(�2^�h]��xR�bv�L���+��o2W cC䚾�;���j��b�W[&׷���M��v�D!`���K�Kr:�ا���IG皶�H+x�U���*c�fm����dWp#kr�ˑ[L���A��hF�`��w��%���7:�
����Ձr�*ꂶ�L��c���݉��#B�Y�G�ѝ;��$��A!"e��0������ڠ�r-�R�¡��n��@˷J㝪�]Zk��5}�U��]�.�-vn��GKnɅ��6�*�F����@��&�>�Ot챺g˲[ټ���n���9{�Azi��WY����+�x��N�O��h��fL��z���=z#��̵��i��9��Vu�xa��88�����b.%���wt��f\�T�{Pl������\�
�P����C��Ƒ7"�	 �u,n�n5q->I2�@3c��ĉo�%���b�
�Q�l�r�\�nfDr��ࢆ%L�̬+�c�
������-��V[�UrԖ�[b��a�ULeq�W.eR%F�d�m�Xۍ��b��X���F5Sr��)�)[lZ����fS-��`9@����TKb�1̪���R��EZѕpn*s*��+.PR���e�Z�KK*EkTm���-T�dR֗,m��2ԭB�U�J��2�kL�Qd�UEb"֔h�J6F-J��R�\�0J�iKh��+��1
��)q�b)�Prţ�U��ҍ��A��bV\h#V�QU��\Q��D��P��&U���\m�aSUQ1�5�"�f[�n5�&7(�j� )h�S�nV�u��d��iQW�u��gX��:��9�;a�M�1c,R�3FCAlV��Fg}k"�ɒ�1o&�0m|��o3zos��S�\��"D�/V$���2�S��J��*�}�1��o��>�F��ݖ2:l���d����"�[X��ƪqG������>���"W����+�����Ng���[�xnG�} �kY�}�Fl�ȡ�<)+��H7�3o��y� ֽ����6�8<#]i�M�:f������W����0v�7գ*^�0�8�3ʴ�]B�yz��z�qI�jq:��Q��l��B�J���ˬ��OK�Ƞ}�7� �,[Nٛ������RX��Jc���N�+��I�k/L)�P��c�[���[v�z����c.x�2���"�{/��no�\�Hڶ;�!V�-�X���3��x����|<�NLT�n�~{�|F��J �2��k�)��}@�>9�]cH<���Kۂ�GS��K*b�w�: hݜ[����ǎ�V��Z�%�dWOve�PA��(�T�П��Q����
U���/ƫ�8+�\�@�y�n/N����
V�L8��_MThU��_��=�Y�7�9�={Tf6����V":�*�\�^� 9��{I�V+`�\�m���|��܄f�&@;-Һ�W2��A�WZ�d��*��s:mٓX�x��{	�QM͠+;��ݖ���h��Tҝe7[�ޡ������W�e�%qCy�(���Û��l�����8_u���ogY�T�2���Y㾽��4O+�<��3O,J�^�l}�!�ҫ��|��o�c�d���ӯ��)>>�ZY���e��w��1]�}e�����6��C����Μ��M+�򧎗k�^Q%7pQU&c��Ie��,��LWS�+��K����̎q�|H���\WY���m�1�۽ b�3�Y3���(0�e�B���g���iY���\U��^����|@����@��~ Q�U폭T�����ǲǪ���s�YY�Q��y1x?�~�Q�⬇M��aǎ�,����g�ޅ�F�[�0�L�H:�c�jy�j��a�+-vY�7�T�Z��z]	�Y����]9��f�����UmL>��zs�A[�Qh�7�{��[z\t�3�|0�3�=��_�Ot�kx��Mˮ���aƾp��3 ��z'��k�L���~���Q�����P7��N%J=��y�<�0���߄�M.� U��`��0�g�OO�cY��gE��2�,��s;U�G�[*��:���R�sZM��Py�����Q�f���u�3��˽���c�aPV�V���*�"W���P;2�څ�`W�	����3�ʜ�P�Թ5{֍@��jPI�,���g2l�b�`�yw8�q�s�a��Z��!����諭����oI�4~ʽ�8��m(�yw!y�?{d4�"��N�qn����7�,�*tyԺ�|�V��O(�jD�z��x7�W-��lVc�C�|��\2�rv���i�[�	��{G�]4UT�+��.�?�p��a��U���xE��M-y�u��z��MոV���Z��s�!�E<W���~ @�o�s� ���Q���.�@��\��w��3��6'�*����k�<���]-���~�0g�=J��	#�<Oh��p#�N��ҽzN
v~�s T��|v�n��^�O�B�h�r�;X��*��("^��=�D��9Ny,����L��K��!���V\;x3u�J����I�ʒȭ��{�Z-���3�1`7��6����[��&���׼����lN����si�7cg� ���d�+eE����������dyI唲�n^���a�Ƿ۾�ϵ�o	g�|Y��8����hx�sk�ָx����<#>��r�DW�������x����I����&�%�����a9�j5!�6���ڙ�*��q�s��Xwm��[�I����ґ��Z�W��>�Ή�Ga]��.0���^�'u٘�J�S�jjʵ�̾6��0W�)����8���c�j3yҙ*e�kV�����N�����6�n����G�-���^��C�y�ɛ���F�����ۈ,���]��
��^�̷�ݥ�L�%��Ruf�w]AeN'���������3�xw��:�x:Ld�n��R�>�KÁ�-ނ��߽z _��ʾk)���o�U~���/�U���o�9s}BaJ�b�v8V�P����KBV�d��m��=__=T�A��&��W�ŵ�i�Oz/S��,�W�J��]k�U�!��׆����!��9�_)B	G?_�41e��#b�y���Z�#}��Z490�p���Q��D�� p� �e��U�m?�9e��h5���{���2�o�l�D{�!���<5�+;Q�#�Y8'n�Q�x"���l���J��r��Z��~9�q��~�U=���ID����%T�WB�h�D)�P���}AB�d��K�x�T%�}��t�qL�ZaM�h���>�Yf�s�)[ˆ����p�rz��3�W^[T7�O���q�uj��֓a����~k��(8��9Y����}���GnVhiKU'1��k���]v*�c^]�]䧉�e����x�:�HĹ��+p��敪��(]��|l1a��/iS��3����]d�s�q�Ӕ�W�ΰĮ�_��������}R�3zt㺁����:Lκu�G��&�\��ꪪ��o�;����k;C�Uł��U�6�4��]R��%*��2�hi��戆zR���I�����;�,2W��@Εo���]���E��=�����L@��j�z����x|�A���r�+g�r�^y!��CjAoIϺ 5K��T����;�C�&���`�\�<����S>+�����U���Ey̔0L,iϣ�4*���g���ԫSD���u�w�sw����:'���Y|3n��>�(?������^��@�"�п7��W[ї�h�Eu��Ǭ�F�YTyX���:��>�^��Z�&Ti
�Uy����`�Y^/Km���Hnal{�2@~�P;4��hC<xRTX��JB�:�t3�n�S}On[v�s��н~;�=5��G֡�����U=�f�}VuT]�t�U�AM^�� �����3w�L��+jq��\U�7���"���S}b�ű�홵f�{{�µ@�����w��iR�G��u���� �\��]N��'c����x�)V��w�����egC�`�fc�
��5�>[��5ܹ������+�Ps���2�Fb�T�5�G( �֩|JK:���'����3"r�|з�ms��;4ݺ-W�å���qPѱɍ4�]�ⵋ��3�Pew1E�Q_Z�x��7���꯾��}�#y/�Nx&I8�Wb�������{e�T�����rK�뭯26��+��ekj{wS~9ݗ�du*�2h17�i�w]��[Nm�Z#���Y1w;��*w����Rs�?O�Y̯m�MM̺
��'�*.�<��badͬ�૭���T��8Do��*��;w�彜��ƏL�4;���Ô'��SU}�*��=�WV�a�z٘���{�,��#���Dsq�b���â�7�s��^���
�N��X<����9eeƁ����G�c�cq<eN��O�!�b���ZYR���yޔBWa�O
��G6&��d��{�ڹH��ٹO+צ^n�D������3�,�Ւ"4!1\ڌW��^�/�|Tl��g,�Lz�xl7�+bbՁ�m�0eWtD��R��EN�q(�+�f�\�Էss�4őb9�.��\l>���<~wj���C�l�#j��~�<n�(:۞��=XI=6yZ�0+��|���*����ư�3�m���eu�iL��d;�j�iH�W�R5쵮�;���f�x`��&6L�{�6�G��z�����&Wh@�#�kub9�	\J6���/VE��Fu�����]I���2�I^5�z�?���X�p�IҙY�(nRa��H$n�ߓ]Wq燑{3f%�;"X���8N�����S:�M}�����������r�����<3�<#�.��Gz6V�:�E��yJrоRU/:�p�Hgq���J��Ν~]1'���M�Iyp�W����Pp�9U5�+|�Ѻ}Q��Jb��|u߾+�Y�x^y�ig&d���.����)��*���=G�z}P��}� �r�߳�d��%��M���;�J=g�E˿�.�	r����ن	ƧPq=>��-�d���y�tу�渺�%�
^�[B�;�\�!�ߔH<���f�{d5��V��
�G�b�'��_{�o�6�9\ٍ6-��Y?@���>`�8s]e5�𔼺�>\*6R�5߅���g��"��.x�2����ӓ���]�~�[�N̺�WP�%醍s��ȱ�ʡO���ާ�yo����|�ײ��I�ϔ�x�O.�N� �M�@.v@1��銀Ch�ӳ9�Q��ʶ���.�c[�:ڃ^ԵCt�s��<���`3*��Eʺe<{o�(kZ�߉xe�O�-Ⱥ�']E�8f���ze?B�h�,���*�a�J�y�,�Ѕ��F��Gh�c*t�ٮ�w]�&�vep��;��u���^�OP}��ś`���e�R����]�ܮ��mj����=�N�v�ڼ!�RY)������QF�5�/�Z�Մ�.�:޳e�ְ��O�c�̝���;�J�]J������iG��s�:�?}��%��d�襉p�X�΢��b�8��n&S9~-:��5����n��ܿy��u�zE���"k�p�k�ryh����L+<,A�]]��_^�ިNuק�9�sZ�Y`�2`�}��Rye,��zjz�����l{n୥�I��gcxA[���ӻ����AU�J/���2������u^��V3���Y]c�j�cޘ]w����؜���i��jUsJ����e_���%���S|��߮���隐Y��x.Wؽ�-��K�i�⁻d��L𕚔��x�J���ϯ�e{��d�;�t�>\;�~��eVj���s���>�'TV2K��@_�W�E� m+\�j�PqM>��	�Cs�=�dZ{	��z6��Lp��g��Aq:��$g�w!95AF�7]@z���4�N~�/_VO�_M���*�����I��At+Q�H��F�CD����˻�jǗ>���/7�}��ׄ5<�DE��=8\�~��Xp�"</�*'�0o�<��N�m{��D��4e����GM�S=щ��B����.8�S},����jPfK��N�?g���7]o�uPZX�Oj6w]K��d���S\�s��4uн�S��-׃�̭���rH�f�\U:���W�U}W�����u�����5Lbo���@�{�!�S.�����;�c�>T�Fy�@{EzY��=��\�V���o���~�;e6�$,3Ϻs�)�l�㞺:~�L���7��y?ZW���[ωu>Q[��H49���a=].M|kg�W]���i������Y.a��� �������36�g�^�O*�ܺ&4���Ҿ'�Uibo_���=~˭���T���v�䇧�t�������Q��&�Z��*���)(9W�4��^44��<��}޷=�E�����V��^�Lf� g�U�#>0A��بD]OWU����I�z��3(���=�Rx��mY��R^4O����PtH-�=,B��S�0״����1����"���[Z��x{Y��iV�U���Ε^s%s�Ч{�	�}~���x�����J��B�V�=C��X�𘗇��ϸ[��斺f�ԃ��0?s�a+�Y���(�s���W�Q[���EJ5Y����ʹ��^�ϖ�	��+����w���OT�Ȟc�}���y�ȝ�&kK۟�c�>4ԣ�U%����\yx5���h�}\ksO}��[+���W ��1��W�4]�ʚ�^C��sdbP��]�V�oU�!�c���A��I]��H�Ə:�]-���,���i����}yV�5J������v��}�}G'O{������lRS����}�!�[5r(g�
H�^7IHs��C~�ۄ�#�N�\�ޙ��~�i���s�]?u��}j;n{+�}=�f�}gQ��q��N�@�V{��^\I�P���9z��jq��xM�~<�"���M��3�ű�Wz���O%z<��q<�A�.UוM�����89�3�/�vN�ʹ������E��Sc�xp�DC�wʥv+���P���{e�Oϱ���r���d��۩�90����Զ:'��u�ۙp�vC��,t9��bc�j�*�iͽ��E=�ԦW�ٗ+��7=��|���G���0p���Y�t=œ�Qw��,DY1��¼[OǷW)�j�&=Ϗ��˒�7:߾���\�G�L�S���=F�ۣB���Yz{*������[3�u9�M��c�v��f��f��\FS��E�������Y�U������K/��s_�p��\g��c��}����~�)�@lmuT��TY� �(���gcz�+�9�ۭ�oI�1E.���+�\�\Nk5̀��:���kO	$�'|��WCuͬq�o�yn]�K`ѧ���k��cN�7|��g4K�WL��]6�ejuh��*��rX��'���N���l}�D���C��Y9�9+(�v�`�|ȃGi��e���������n��V=�T��r�5\���y���p��s=��Y����rZ�n�YW�v��̏�~�\P��w�Oeh�h�(U����(����k&��휹�޵i��!�V�ekܗwx�$�X�jtWlc(��w��yy���X����I{��jf�l��nK�э���]�mru���b�%�\���,��n�ނ���T��J����Z"�.�������]΢i��ك�(�#Et�Z��������yoM�BU٩C�fE/����e7�&+�AWryE�f���j���U�Wv�5��Z�LN�|:�f�[/Q�w8����|�s�\:Q��ꎮ�C��L �P��|+u�i0�ي�.��d.;�s "��v�o��X�2����⺰�J/r*<�6��]g)���3�m��L�PM��ه���x���T�̱مt��*sa-bWINn�L�ם��[,�����1\�ə�����b�뵭ĳT;ד�k7��]N�G��y�uIZbb[]Y��w-Z��X���ss
u������{��v�E��U֐�چ�A��K��m�����T{9��F���)�"HB�L�4�6�^9L��*Ld�"e�)��!�])��6����K�{WN�\Íq嗸7�Y�e䜦 N�EUު��(�����V�e��ِ��jw����e�8"�H��!���Y1��`��U���
|��F�QEv�s�t1�r���#2]��+L�����m��ұK��L�4`��|v� 9Q3�P��%��2��k�4�0���	�x��Tu��S����i�A�oP�j�1��{�\' y���*�3��d��]��gh�;[�`�Q�Vg)]�g7�Wu����:�NK�핻4C�
w)Vd��e��b����GX�)cj��T��k��Č�[çv�z,�.�C7�ՑV����� ݗJ4�Z�SC�=|���Wk{��۰�����)ëN���޳ř�i���GN07s�kj�����DY�t�����X�$��P΋4s�u��B�9lP�տN]Z1��^�����v/JgU���Y[i���su�j�4y<�voIJ�/N%�e�A=��<��t(������ǰ�oS�wt.������K����o�f�N)�=Q��_\wMt]j�k�&����[�ܧ]�r�a�v��Y�b�vU}Yg��dޛ�N������z�x�s�:9olGY9��T�l�qb��Y˴���*䋻Bbvt�87����[I�u:QAP��Qάk� <GR�� �K��7I�fkHz�iT2��1IY(���.e�U+
9ZV��**ֈ��Z,�X�ihĹjf�Ad�TbT���1q�q�7�72��-�-�0pQ-r�TbZ�*U �E*V����Z�KKmDE��W--�5*"[H�*�J��(���h��"����V���F#1*��LAEULme�T��T��`(T
 ��̑QFV-QD*��Z�1��X���jT���"2�dU[Z2��-*ԡX�b(,�eQ�Q[Z5�ZR)*Ue���Ŋ���f3J���4�Vh�+�P��b-
T��kiKmE�+�h��k�����%�]�*�"�ST��a]Ü���3l�W�3q�T!xK͹:1]}xMզ͘w��)	��磌�������������0r�nSϽze�}�2�*��(�3���Q�{E����u�,h:㞝�f5�յg�@�3��a��\<��c�#WtD�r��ȩ��^�
c��]���uxB�w�`�|����M��x:<��p?+^���'�J8,x�VǓ�����Kf� R�1=�WK�2��Ҕ��E���u���X�|X�Gq��o��ke`������Z���w��[#�6Օ��,����
����ʠ��,#:���4��6�^Engc�ۭ5��J�%�0W��K˃ʾO��8^����Qh�>�>\2��V�0`^4I�=3�ﴤ��U��U���uԠ���Í|�V�d��81�M1�����)���}�]��ܰK%�=1]��� =��`�&�q�������sn���o\C�n���0l:&(��CCl4�X�F��OL����6����<�
���L\ϧL��8i���X��1����XK*:F���y`�:��˲�ܷ�PK�����
�x���b�hz��@�m����3+*.������=}�M��s����k�(�܇�{܍l[jv�G7�ہ�_��$���iUқdu:G�\�t��C�f:vA��j�-�����gN�|NDc����zYy�yC�z������H��{�";:]w�h���f^����'i�K����N̺1]C�Q/LϮ���[E;tys������=�Kj{R��I�ϔ�x���3�$��v@���R��W�+�ư[����1u���s�(5�z<�n�N|��<��}����P]n��c�,�
��ޜ,��I����\���O\�-;kᡍ�~�k�)��C���hHck����c���~�0J^�����b�%}߬��0�%�04a��*�Z$��C�gݨ��]��ݍ����ʄ݁����E�=y0���׼�B����'����m.�6�o�w�37p����2FI��wM��^����_�˅��~;e״P�Hk[���o<A�i�V�#���v���B�8���7���u�Ś˜���2���1�B��1�'�qqC~KE�k�ۺ�|uYT����|̡��d��|��ۃ�������U�".��s�WYo
z���a3����Clணj���7S��d���.�к{ˮ��.c�+��X����ָ���u�Z
����YP��_'���͡��Y���\�ѫ�ł������K��G��3d-�]���(+:m�SwI�*1'}x��:v��sbY�`X��kwnt����Wiꏐ�Ua�뤗ӌ"e�������G�k޻Pc޷m�b��9c!��s���"}k���>[�)�����o:W8�M�{�����zn���m�ɂ8S�E����]A|�.�w���HiyF�����=B��(�ݕ�̞�{*��5��f�X8WYk�7[.��ɹ�(;7aف[^�&V��휈�yV�2���N{�Ǫ��h</��o<�f��랞ĬW3J��m2}�S��Os�2�]o��lt�V8u>�f���q7W�'Ϙ�����É�닼x���P�0OsHw�9A^ȕr9�8�ٞ^j口9͂Y�w��x����v�g*�WK��Tkg�Uu��?�r[?��M�M[�<��F7����]�j��^����T��8�������z�j�����eD����F	�K�NM�IZ�1����x��^R��ϕ�Z��v������z�g����ҼO8vj�C�_h�ʗ���v�S�oH���B�e����=uܱ�XI-�C=�+����0hʃ����Aqyy�5�Kr׷<cˬ"X�Obc��KZ��1\�}(�-��T�K���P���Z�F%'Ϡ��TWV�+U��2/b*��,�3�(+|y��f�W+���cvT嵽�W&c�w0=����;0��_W�A����^o���\%��fl�W�62 ���D�x���P��Z+��\���xE�@;r�螗�F,Ǟ��uU�i9[Ε^s%r<#E�v�t�5����ڏ���7���ｈA�5�!�7=|��Y�A=[z����E/��*�}�1�3T���#>��(n�0��ӊ��KߍT��<�z}��u1>"U��=���r�������������>�S�c�/������٫�C+�xRE�񿒐��A����s��i�Ui{�gN��J�&|�1�nfGt�k'[��qo��f��,*��V�ʀ��Wޚ�z���I5���VЩ^Mu�!ʽE��8������{�@�Ԧ��E�cw|A˺r�'s}��t�E�k�N!7��g)��u��fh?f���<�u�wxx���ݕ/�-���JF�����.�]
��+�/��1*�x��j�B�o�oSz�nu�W�]�c�g��l��l�d:@�КM�Ɛd�#^��iͽ��2�ӗ��׵��-��w 9c9Ðz@R�,�[�g�����B�+[/<(ۑ6V�wH�t4���|\��K��v)��Έ3�Ķ�vy*;��i*�5)��s�1�_d�`⫊�����sĩ��{���V���})t5�H4�؄��Xi�T���}�Ϥ��7m�[�_�ql��5�4�]*ne�Uœ�w��][e�b��t��=��Á����7��]�M�o*��>=Y&g陸Âz�E�B��ZK���;.��w�Vf�/��ܲ�G�� ~~�����]��<C�FW��A�� Ɖ�t=f����s�����M�=e��l*���c'N�t\,e7~��sL��ڕR���*��_�����3��"Gp�8h�Ď�u�V��:Q%�r�w-�Wr:r�<�?z�Z��3���˨�	����Z'��mY�֠*���<=�d��X�3�"J�)Ql��)d�߳���sܕ�~�,,0Ӱ1���<�=���顓�E�P�l�:�D���Z�O{ֆ�����W��;�g�Uʭ���C4�~2�f>�2q��ڂ�{���m*�2��Ծ^\&��w��^9I��p�<�T�=;i�e��s�����dg����ͥΰ�U�t>�er����<>�~.�kPV���l/��e�K��7\�Q���m_{i�)�絘�3����wL2������(7��n���F�aR���N�p�B�p�/�3M��]i���Xn�.�[if}���ť@�>�.b�;��X�����J��*��Ss�ism'�Wj�w��hs�j} �w��}���\�i�.L�и'��+�=;�嚍D8��Unf@:[��#��W����ޠ��c��˖%Wj,�6�$�z|�q�V����*ƦK�M\)_��=<�òyֵw����pk>�!�*zX�X46�Ht9���{���Er6��_�Q'�s2����Ǐ5��M��c��U����ҩ�f��a=A�fUY�)[E�@�z�{�f<��e�+��|e��SQ�W;瓟�zvf�����ˡK��u�^���Z���s����J�7<�:2���f\n�Z���Nx�R�O�\3>w��(n�V�֯��(/dA���Ug��{�W[Pkߥ���ӎ\����1ݥ�Ѵ�e��\ݿR\�V14�$]S�x����P�6�M}�ͫw�߱v��^����*ae{ɞ}-�x-(�Oj��שA����]f/-�\5�b�:���9�E����3�p���|Wb� ����>vEm��=�S��Y0:����b�P��zI����ѫ�Y\���8��19����Ǹ:�������j�<�c9���o��ʔe{B�Tu�<�G��Qn�,���5*��c� mw`�1�W5R恅�nƈ;�b*��ٝƄQ�
 �r\�'WC��u;Qn��z�#�gu-C�>}y��U&�{GH�&=����D�`# *���;#�O,����js����/z����{my�g�{b�~��Q�PZ<~���m>R�q�:I��~��V3��r��\�.zV��Y���ܜ��/|N	�mq��ԩ��E�/*�9L�
��&NM�c�n7�mi]�i���n'��WX"\���W!x���0�_O/S�3���N��W3��2�����u{Ш�������Ʒ�߇0��0<��	���z��,��~V�t�{��X��L�{]�󭃹M>8^�d��_��&	���;$Z>�^z������K���xm)�j!%�)V�\'nnT�w&�z�e\�~��w>O޶k*��+��l�/���ví��}��K�o�%W��>e�騉>�U�.v1��滏�a���#����Ȑk�i�~���8)�Ez�iTˋ�U�lM����s�"5�y�lv};�c�c���c�)��;�c{/x���!|�F�Dz�5qw�W]�^���q�T�<C*���{��<�K;:�uTY7o�2� |q�*��|$��^u�
*��7C1۷�����;�Zx(������tE�2��o",gA����6��� z蕯z�w]��%�	�XU�wer��6˅7|���w)NkzQY����?UUOq����O�hd�v+����Uw3�E�����l�����{M_�Ao�F��z�7�d\��]k�ͷ��e<��^U��7.�r��]/-�~�P��l��o-�Q���_{-X�뚼���R��������*���1�d׵��U[�]��;��ؽ�:��.|�|J|�
�Iv��|�Ͳ��[�2�j���1��eu_x�ꇬ�g���h����%�-�3��������AT�ޓ�WD����O{7�u�O7$��GA��{���ţ�i>+���Iz����Ε8�o�%��=5v{CJ;��ۻ�n��zC�}���^)�ô ��Ֆ¬Ԡ���FP||+k{մ��?_�W��rwr��bZ��P@:իuO����ѤU/��&w�N�dx萀N�{1k6������m��g�!^�E5�\��j�_qϡ��W"�W��,W�����]�a��d���,:��L�Z��V�`��T��z5^�K���S}Z2{��>���?G�$7����F
��J��R��GW4��o��r��o���{٦vM��h��"�V�*�����PQ��y�rE�,���q���jV��N֥]5����4B�MΜ&Y�҇�c���u�9݃`���f�p�Y�vމ��ԣN�%J�[ҳ���Zj߻|7v
��UԡF�4�g�끜��1�8������j\�=�o���z�3�u����+g���p�Z+�ԫGu2�=�T�>..g�N��t�{r��ڜ͞���w��	W�)���x�s�x_��}��fv\+)d�V�ܭ�Q]�&6u�֭q�2��؂���*�>��l�vC�1���b,i�5�
7�$i�p�j���2�m^uڦ9cܥ)��w�;T h���E9�]}œ�<�[V[&l"����&}M����]+�Ǳ��/��8+�����y<52�I�B���%}e��uo�����=�ڭ�A��\N��p�����;Z;��G�FW�<Pl�@1�x�C����v���/D�����8͂G��w]�W�[%�*���c)��4໚zAhuCP{�驨�]�2�y�����<%m�D*WaVXدc�\�]-a���J$��^_�'P�Y����Ո���9�#D��Z�\;���g���*T8l6�eI��^,f��&J�W����Wm�OS��8���Ä�6��1���hǇU�]8��ކ&K�J�ӈo>�3�[иZ�;Ct�KE#�j���U�WQ}Z"fј�O��T� �����i��d����k$��WAv�Y̮�[�yi���<�	\=:I�{.D�,�;�|Mi�C�[^�����`/����������/<��p*ס��k
�'!��w�8.�ŉ��v��ϼ@+�@)1=����tוy�r����cG�\�0��{Z�}�O��iv�����e{mՋW��=
q��*�>�����_��Mv�cU�H��^�~�sǑg���r�*�.�W�%(eP�C)|��<��<>�~3�lW��-��Ϋ��ؚ�9�x3��|�m��I�g���%]]R�A}������LC�=9�z���/<�c�e��ϯ�8�]��d�\r�Z=���U��evم���u�����l-f�����NƳ�!�.]w�x��ʫ�A�x=�)/q �W�H9�nR��nw{fkki��#�?N�,����u�*�z�Q�TĳPi0���'���ò�g$_�;d��x�a�rߎQ�b�����e<����R颪w����ЭWP�̛��0�z�9�,����O�.��/�DXϯ�x�S��ײ��I�ϔ�Yw^��NV ��U,�Ӽ7t"!{�����f?}���rU�µևc���Ǌ ��(3���nX��v���<�ǔ1c5<v���%,r���fn@���Y���)���I3[Y/qo^��nW=n��-(�Z��Ͷ�S�}y]�n���v9>�Uti��L¶��*[s1�T5- ܼp.����9�*4�TǕ58��5�0}R����3V�c�n`��S]ӸU���u_6V�]񖊊*��Z�����Fɼ���"��lL��𷸆;�T��T�ܽ2Wp���,<b wb�sٚ-���n���d-�g��4Y�^�7dV��$+�M,e���ֈu��`�s&����ױ X ��K5��uXj���z��8J��F��3n�7������o�iuj����dX|+��T{>Zy�}h�� ��t5��^\�u+p^Yo䱇��e��u���?s���l;�lPugU�oYC$�Vr���;��x�0ut��P^��l�IYܦ��N�a�[C2�լ���Πx��xy#]j�������
�[J�vK3��V~�h��ڎ���׽�bX��!m����*�����r�A���٢"��`�]I��ne�6	Pҫ�Ԥ�����SW3F����W�C9�o����u3ڳ�	"'n�5i��9�7���r��t�9�`\�Gڮ�-�����ӻњ8���v%�`�\m�u��v-��n��Ʊ�����,���zr[y�i�Ÿ���L��Ӝ�U����t(�ŃP���ݒ���(K�/����7�����y��B���N���Oƒn]��PbtkZA�V��e�WɆ��K�l+�����d�uu4��/Z�]��o;�i���졘���پE�#{�r���5�@�Ku�~EHjq�8�81�z���R�VaEK� ��:���ö��9qĬ�BZ���T���Z������听�(gl{���Sn�"�]���9���d�]=O�1���yq��*�k�2+�sd�a�͘�&x�ˍ>�;�$]���Ӆ%��ʺ�6��ɈS�t���h��%��[du�aTͬ���v�ë��_A���3"q�Ak�-=�*$%C����:�==1��'���M�E�p��tyNv��wP�����,�=Z_b寫pJ�ڗI�)WRj���Bv�B������/2mdZ��B�5�\�$����m����h̩��H�
=PnK��\�QU�]d�t ȓ��j��6K��� ��X�\"��0���qղ�=��b�K��xu��̰��b>
_gP!�����N:d�S�]2ʰ� qv7l�&S��#�f���(��L����a��Mw�/�d��N4�M ��\����Xov[���Xï23M�����ǫ���c`�OX̹��G���
��u%�bcخ��K��CwD�o+x=̖�6/��x����N)Y��%Qim�Q[kwJ���ؖs���kkU�1)r�#Fe.T-m`�T�j6��TKJ���lR��eF�m����V6��Q���E�����4s0ʴ��KZĵ��c,cj��h�k-m�е+Z�ʖ��K�J�-�j�Z*�եm��Z���A��e�JQ�ڥh�n+lK#Z��+Q���(P��r¢�8V���ˀ+��ť��լZ�(�V��%���U�Dj)VZV֍��ZYkJV��R��Qq1\(�e�1�V��Dpk�hV�l�ڊXܸ�)j��X6�UiD�EKZR����*�V���(�UF�b�QckQ[kQ[F��R��(��lF��R�Z�cJ��j�J���+D@   :)��¦�ia���b��t����k}�E�����Ӌ��ѿ����*��|�i*�<����1�����9*��U�6vx��Uu�j�Ü=�9n����׿K\4?T7Y�)˘y\���R]��\ᗷ~�ī�Rc!�H��Y�U��U
cr�꣐<�w�߱v���-��N�W{��sz���(�f��>�~���]o�fR��I��B:����ߒ���hXk�]�v���ٖ��2��X�]�RY��<UI�ʞ�|��2��_Zk�޿��X��X�֒��<wu��Ͻ�;" �b2����I��{����W�4�T��Oo��y��ٌݽ�7�T�ꘪxʳl�}Z�0�k�^q� �N�h����ʱ��^W�W�ہ8
{�7�-��S�<�Ǽ�k!�ۺcj�uYT��б(`�/��9-�0>��T}<��t��9���^���	f���yr��"^L��ɍ����
�uJ�oT��U��pS���$39��mL�x�Jo\���._�V��>جd1r�g /��"Z��.��er���TI�F�[��4�֫ePqM>8^�d��y=�T01K�,�e�;Ts���H�<�t�ī8�_L�_)��[G�K5l~�=!jѳR�%i!{���BxT��3�ee`�!P�l�����ẃ�+r�J�!J��gh9\�VX��[�6�l�sA�(JW�vT�4&��9����>��,B!wZͤ��|׊��u�V������f��Nrm��3�n��7q?z٬���T+��]zл׻�Á�۶���=Iĝ�W��7�;��Z �N{�Ǫ�ϥ�Dw�t)���N���,r�(��
�}I�]�mq+�؛9���Dkx�S������ex�frN:'����ڍ�$��@��Q�\��i���s�l�;C���{�!+;]���6;��}�ᯤэ]��]�J�2�Ҙ�خ���,�`�v��,U�M
~Y�3��`=�Ǽ����xyy��6|}:��Վ����T^�M�+����W/�YIAʽt���P��(��ιϻ���|'�,=���y@�P�CR���pR�yJ�S>VMk��w�'���ez��)�/�&�xxz�U�b���Cϝ�����L���[�0���
��
��/2�dͮ���5;_O^i�,�>f,J<���
[[�(�j���Pt�ޓ�t@o�jݗ�}�ܽ���İ1�#zri����+g��]WŶ#ft5��haZ��w~j�a�!�E���[|��Ơ��"�M2�Rv��,�����d~�mߵY/����<�^�C}��u;6�1**�\C�v�5��Z鼵��#u����do}���3,���k�t ��[��N���� ��9f�}ϲ����uҍc�Q;FNyo"��;gWqcX˃�6E�ٷ���5��oj����n.�7��ň���|�����"��={��V��)�>x� �j׋ܸ��ѧ�TQ���en&m�Ex�����zu�rWF��Nݏ2"���B��j0k*k������@�=�6ʡ.�j�]!�%��_��Y*Y���9T�#����\	jbe��=��=5��G׵��}s�^X�ESެG��J�;ӽ����*��]B�����[�^�"��=E�^^����dPwMf������=������ ��%���Uh�KԫY��W�y�q�ªu��3�v%3��{^Ƈ�݃����e\�Pa�<E:O�Wb�}v���Ϟ�gr�NnE&;χp�ߪ�����_]DUvT��d2C���>�,EX�>��"�o�T�RI꘺T��ޛ	�_vy������K&.�{� h�$Sٹ�A}\Y=A|]�y�ձo7ۙ��a��B9;��6b�%θ+�}/���	����38/T�xpOQ���4+�<N'�O�Fξ�S����4�(]�򬫒���՛�]C[���>�2J�N�5H�p�����G�5Sj)~�r�±zv����Z�]\.K��{rn4��q�Qov��WH���|α=mN�����ظdm��'����[)�oc]�s�_�,���-���:Ξ�{����T��:*3zGS��ͻ�^��5����5�<��.����*��1e%O��7��gJ������Х8��AhuH�||(޿<qӉ�X�1ޫrA������G�y�:��k�R�=���@��=t���F��})�5m��l���	��'ܭ�>��P/����p�%���b0/]s���#��n�{�]ę���ކL���H����uR��[�v����~������QU뉷�ا�><'m� h�7z`y� �&'������Xi��cl��-(U�����E�V�r�V�cԋ��h�W��W���ǡC�<��2o�n�΍��\'�`�7��2e�{�HYo/iO���s�.��
T���(U����us00�zf����yWu���k�o}�����z'�z\t�3�Ixa.��S�N��35�[��{��49����l�2��{Ȿ64p�|�}gc�ݨ�r�+����J~`*z� p��S����o�4��i��?�ɽEY����x���X=���[�6��=�;�)�b+8��,�s��ʟn��y��������}�N�Jk��i<������n���U���(�U�[N��Ŭ}`5�����i�%�ǹsq�ή�Y.�T�/V��M���cc�����/�#�W���`q=>�p�5�P��.� q;������B�^����(��㹝�0/�SC���^��Ժ���}�~�J���@'�x��)?g�ޔ
^�9��~Į�s�m_[��[�l��ۜ�y9�G�]4T�+�;2�U��i]��i�Un��c`P��+�c/*��^_Y�j��|�(5�K\>��B䷅J���%Y7�
��[��|��N��m�8J�x�v@1��5t����r�9�[Pk�k���n�N��K��s��r��S��p��o�<�� ���4%�����~�yeF�CC���(���:\��k{P^�^�	_Ge�qT�E�PeK�z6�墓��k�Ŏ^� \��8s`ɽ����\�����$����I��,��
���OfT�>VL��U\�ѝK�{��8��{�q&�§�)�)g�{܈+y�# )��;#ʪE����8�x�
��Ԛ]���+1�W������f�d9���������G�h���s������G.��z5����k5��h �,�N�����(�JV �ްm\b|m�=��Ӡkh�4W���n�jTp5N�F��isg�����2�R�7��St��{��D#y ��ln�Eb4gbź����7}��YǴ����@e��\�u�ç#9me�6�=��o�u��ksR�2��Qu�ʽ3(x/8�*��y�p��ݑ�y�C�U��Ù�F_�#j��	����/PY�][�M�f�M��������v;ԍ?u�d��A�S�����:i�&a��v��+�h��!�+zql^jF�ɝ����cr�YO��4�@�z}Y"��& �N������yX*:=[s�_��o�cW��;B{-�#<��rj��s����ۯ}��k�T5�?g��<.����<���:����ZOZ{���'y\��夿��p�]��u��:�����tY�(�/�h�J!)��ө�̶�O����+��"���(�<���W��7�;�{�C�e���3e�<��r��f8�ԺfZwާ���F��,��F�pc��닼r�����0W�k�wЄ�ޛ��w]��yz�Vdy��q�)���/�9��,U�MQ���w�n��U�u�������c/W�Zѐ�|�M�/CHJ�^�"�*ny]�,�I��Z�t�%��D��/s��۠pA��<W�ͣQG��%֏�]�6��'�K{�@lb9|�V�gl�}(�Tuzp���V顨,�us�����*Z�&�\��&�v���&7������I�z��L���s{8�')9W�H��u(G���׽f�澽�<Π��K
&�����w�R�Г.
�U�c.ɭ�b��=��59Ow�l��A��z�K{N׽�������o��0A��$*
���U��M{[QI��>�g��W�]e��8�����*�`�7^Q*��!��
��[�k���띹�r9�<���P�8��{HȈ���.Y��^
�z+[��ά�;=�u�`�w���)�RQ�C�~�D�'h�&�8O�N�@����R�a}��O�U���~�rpī�Ml?-���5��׋u����<��� ��V��C�k^�Ea�����gۉ�0e��/�uxw��]	�%V����xL�4�{<�`�T�1�P�tg�5r(ez���%�w�@�\C^�4���;xf�FW�N+%��g�ې�Z��nfz5OMg�Q��VK���S}Z;ƻ-�o.�#�ȩH�(m&3��Ft�=����UmN0.�wޜ��Jy����-jve�u�[�{��x.*��}*��
_[��_QbVe�{�0�9��Ytϟ+*��oƲv==�P�����v���(u:ӗ����n��{U\2��l���5̖���^����E���c<��jT���_G��V�۩�Ō��ݐ��`ڝN�1�w�K���;<���a��vV`�;�Pd�S��1�1��{shy�ϓ��N�(:���2��m�[��Y�����xT�U�����}Y�؆38T�7[*ne��]��P,t&�q���n���
���~��x���M
���^��)ƶW��׾;����u�NjWC�œ�w��>ro��z��S�,�7ɗؕ&�d�+��~=�.>���p�I��zy<9T:�n���༌������v[��3�ʺ���0*γ�Wt_oy����������w��eƊ^�z5ϫs����*S�xVf�YIS����gJ��CM�A�������s�vdї���C�W��j噂|l�+ah��5)��d����L�:$�7�=��Z �\�:�y�R�f{2Pʎ�=YU"#B�1\N���z����#�R�&-XTםJ�u��E�����3˒~:&�"N�WFK���gI���Ҿ�܌J�6�M@^y}/�]B���q�&���X�#�S�P����*ޘ� ����z��5�^�+�C��6$���Z �[�#7�U�i�A���Iwˈ��)��D���xS�x����3E~ ]���\.rR�c�EX/�s�U,�M��%Q˩}+��*)�U���.殐N�p���8���;@!�x�� �%�Km��믰���Cط�k��N)���!P`�:��X�L�}���Z��l`�9��V����»��Y�֦���V~��9�R��/�>U�>��R��}B|*�}N��u^��E���
�곬���,&�oo+�dۥ�z��6Y�6�c��=l��WWK���=T��΅���q9�~����Gw|!�OO���5�&A�O�\��J3>J��Z=)���z� ��Ѭ�\�1���|��3z��S���ꄇD�U���U������o�W{���ڽo�.�y�O��C~������u�*�z��o��	�>�oٚٝs���2˕f�%�f���D,Rߞ����59燡��'yX�mc	p�S��6ǚ�r��.��/>���"�_\��w�Z����2)�W���s���U;/69s���W����
���9� �7���
��O:��j�ځ��ٲ���	��5㳒��{vVC+v�^~�0g�z�P��/��%Uۺ�6뭟^W*��<��Q��X�-}��d��2n)/��n߅*ڗc<q�詛�\��n���l�87�m˥�t6e�� ��Ǹvفk��i�*����f7��b$&Ά�^W-B�^���J,P��t��yR��{��z"-��H�u;�ɨy���n��	ͼ�fz��5�^e+�����S�T^�K�Ut�;��¯n��\��:�Q��r^��8?UZ��	U�%|:B���T�Em�'�*y�+&���/��Dزl����u�r�b��^,RϪ��+y�U# H FH�Rye,�#c��o�l�$��h�ͫ�&3v���f�c>fmu����(���3�p=%��-�C�ا��������"�q��m��ը^&O�]'<i�n�K8�R�S�+��Xx��pT���G���bz���r?��K�B����:Ƕ�4��R�<4S�)�ɫ�_�>��ݮ����VO��d��5q�z�p�>�b8<���ve۝�T��	��E>�<~;��	[l0���|�S�qM>8^�d��z�=����/�>F>Kq0'8�u���ZB'm�<̄�[��<ɷ^�W5���'�[5��[�%�g7�<.���gUY��*��8,v�_y�g"#�U�.v1�.k�U�@��P�P��Y�Ժ@A}W���,M��T�n�6�Ζ{�w�Bd׃���rr;�r�%���rv�E��ܾ;�we����z��U���qN+�ዱ����x��3����Y�0��q"b�,�f���\�����Y��IBQ}IX�X��s�e��VQ�� �}��3x�b�PR;�+Wu�z���ž����ī\u�\�nB7E�Ca�@��3d����з���4]ʲ�gy��q>K��(n����q���e�,-��ɜz�@�7�u� r�)������!�܇U��|֕U�k�v��c���4� ���;f2N^,��nѐ]��R�Z��� S�MH�Q��H������%ڮ��ó` -�v�N����|4f��R��^�ٹ;E�y�+�+&�#��:A�sC�H��6��c��n��]��zd���ktWd��.�n��`{��n$1KiiF����F^Lk�%5��WN���ǂQ�ǫ��]��VR�Tn��n�{:�>W�h��.2�ܸ�U�x^^V�o^�C���]xz}wlE�})�f��K��[�[4evq�k�L�,p}��(#�S���*�/nS���[�|���U�I�Y�Y��w�p����5�M����䃩"'u��� ��c�?W2�F)�����x���u�7��\��u%],
��j��Z���lq�Hk�8�	�̮�	���G\�׃p�������և^hJ�t��t�ot��@�r�-�U��#���1Kp�8���=��Y��v�H����0�.fCS�'y-�V;�/6��;K��pS��":3hԭ��S�F�}sz;e�7�er���4S5���i��6蓉�уU�ם�_״�m�k&9�-}�i�e`����v�[yk!��a v�����l]��P�r�d8�㔭�{C���n�x��2�&��h��� X$�)�}t����hmhqϳv�o�����:�M<K�'t���Q�k��ޫ
�L�o��&�j�*��&�����Lw\#���#�.ڋ)�X*}�:�:���ٖ���+���Uvev{��.�H���Ë;Q�o��Ӏ�d��1R�&oz�:{4K����F��2�=��=�k��%�8FW\3���:�5��x�����W���H��uS������y&1ӻ���ם�Yqn��J��V����D[^���S���6m�]2�絬^ٟ��u����s�x�����ˏ+JΕ����IR�����Xoj5��S@�h��l�}.�EK��k�R�97,���u�Zٺ4S�1ۤ�T��]���x��ԗ�U�0]�bܓV#��J��(�[w���tH��/�)3I�Lے���g��83�飶��X��zJ�Hp3�}��^�Μw��n��J����t3��Ś,�.�;�j�u}�ұk+���MǷfr_<yc9��9D����ٗ��N�;d#B�4�&%�-V��4�F�kYJ�m�J�Q+�Q�K(�6�F�V��Z�,�\�V%Fe�[`ZЫm-Z���4�hѱj�Z5-��նR��m+*+F�ZR�֪�m������D[-cR�YKjZ4)iR���XѲ�Qm�mJ�-�,+jZ��D)DV�[e�KbҌVҊZ�Z�ZƫDQKk[�-ҩm��	h[Z-�X���j!Vԥ��[Ym��mTj+m��T��mE(�-���ڔ�����TDT�ĕYm�[[h��mjTFVZ�mZ���Pm�օ`���̵0@UbZ�JV0kQjJ!R��F*��k*2�Q���TU֒�5+k[J1F�����������R�[j%���������i��-Y�6�]Co��9�2'1@bU�U����۾��i{}�3�t������%P�/�j�k��I�K��z�к!�ʱ0G�:�Ez�\ʥ��k�U�lM�N� _Os�7��|W'm��x�N�v�4WV��ps�V8s�(�Y��F�5��4�Ŷh$+
li;-+�Y�����k�,�#�PW�%\�9�1��]	d��ɡ�]��Dt4�ȼ�Y���]ڄ��mʨ���}/�}Y.a�S.aȽJ�|���NY�r�4�u:���C=�似�t٨��<��� �1/�b�[��^d�.�=C*e�J^R��ϕ�W���5����%v��D�Op���������}�dFP�x�J=���o��J][���9=�'w�+���
�:[e��qʦ�x?�c�6)��e�x���6��¡f�9[�L��̷�,`c��@Ǆ�H�^��m�8lŌ���|=f�v*�s�W� �\4;Z�澧�x�eu�N�cDxmN�b%����C��WN.��xPڃ���T��#g�;����R��U�8�.�ߡ�}P�о���Z�r(U/����Su�TiQ�����@�F0�{'f.ʉ�H�Ӯ2�*k�)Y��\�ˊMӎ�A:���R��=�[��/{Y����T�x: a��p�����ce����y�VI:���Q3�����s�/V�s� M=���<�	,Dv�J�����͔�iv������~�^�ϖ�	ج�55�Ms�
e��ѷ�a��=�&{��$�F�0�3v�ϳ�	C>�ۄ������:�F����p><�ɀ�{�6!t%M�udM��d�>:A����:y��}l3������ ��g�44�W����)��m��b�'��\���\y��c�2��p�V��!89�w�C;w�<�a;�SݙI�m��Їut>�p��ӓ��N�(:���3�v+��a[������X�o"�̿nԃ�yv*y�!����Ӆ�b��w��Ϧ�[8]��|U]'r��U�8{ٻ;ǓŽ�Ү�ң����f��{��d���|t@ќH��M̺�'��o6<��;�Տ�w�,u�-aW[Oǵ��d�gÇ�$��[F�Q�b�|��FWu��QHͣB�4-$��<��x[3{>RWf���g�w�\E�4O>�:�f2��;z1m�`sW�0O*�Y�U���RT��Ack"8^'r��W�G$�ڦ7H�>̦�ވЬK�Y�%*gq�t�`�T����GQ���#s:ѽ�5t.������o��Ӊ5�wP#3��>^i"�t�	ujXh��Lۻ��s��;�Uݼ���d����,�}G�=ј핢phb���T�*�O��c#���/'U��2QS��gnɬz���Վ�Qf`����+�����)L��s%t���o���O����A�zG}�ʉ3=lQ_t�t2K,�c�z5�9[V}u�
�P������\�����rgoL^wç^��+�"J�)QR*t�%�:O���T�f!�L��uݦ�.P��k�j��}��ɾ���{����0{��P�:<"��;�
ړ�}]/��MyV�@}���)���u�T�WK���D���^��=a�e�c�b�����b_{��n�t߯�2cGh����f*��8�Z�zvr��%R�1W
����'¯�ԭh���<>Qz�ֳ�=Rw_I[$�+��f�PV�E�tǷ���qX7�z�Ϫ�%VJ��]t�`�a�ý�SͩH�0���w6rݯ�I�K�Qq=01��L�싮X�]��r����tyy�n]�kb~�=�ķ��:;�ǶaUṗB���{�y��~��c��hm������ۻ������&^!�9�&��H-C++� u*�m����T5{9�sU����|�xOTF�-+������N��U����KV���9L�l��s.�_."
�f���'����܁�/��<�l�:�t[��k-�
�,�Z�N��;�JW3,.]G�5J'sG��^@�`A}49���(-Z�ќ5ݨ`���@wmsW��K��c����Yw���;d� ^��"�r<��o��+���s�O'?h�˦�"=n���y��sz�\�x�v�+�P1]@�5Ͼ�Ȱx�;N�^�\>_T�����鳥Տf=z��pn4ӓL�e�	>�`^�,��}B�9t+�y\f4 �����^t=1wJ�wy���K�}�<�S���J
n,�oA�1	�`�|��yd^d���4��w�:t�^�z��_9�ڼi_-�� �]�(���	ށ��e)����j�wgy�|bx��"�gon�I�f�B���Y�#�OfT�3�d�61�}~гz-��4۝�5����c��IAW�+Ō��"�ވ���h�} � U����2�2��vw}�8\��hӘ�V�6q����e�.�M�XLU8ʳl�V����@���xF���OV�t�қ�+E�=M��5�~�a��,�`u���O��k��GQ�V��Gݓ3k��1�1v�/^꥔<�l����%t�*�^F�/�p�g����C��荮�vZ�9��::R�GVv�T���x5o�^R�e�u������=���A�|���W3h��d�!M>W��3u�I�0.�i�"�S��9�f'w�o^�Am��ntX*�58p.�Mi��ɳ��tx��M5 i&�sS�n�N"sr��.���D++��n��IW�À���� {._�V�`{N+d��a�fe�/�8��r���{��X���3��>�)��/J��o'���b��t/2I�޿7���R.UŠ�˔-u�H�;������s����R���ϱW�zۭ��E��I����>�t�-���k�[g����IJ;d���	���DU<�D\�`�k�@���﷟�C�n�^�������Z@��
~��\�˺�[\J�&�v.T��оPE��_����o^�ݳ���:v+�`:�,��B�?P�+�=�K<��Y;ur�<���u��t�`|X��霠�g�ev�4�'(�|��>�!��oՄ!BY;��>w7��l���>˒�	�{M_ʢ�_��%�5c*e�9Qz�<��ˠ��=|��U�#�ߖ6�䒶��j%�*��t���_V�&��������jY�2�/)T�袜m�Ny&�qx�}5������~����U�U�2#(A�ͦ@ʐ[��x+��������"]����Y�EU���f��C�m�[���z�q/�a6+l�[^o��	{����l���vehF�A��d1w��X�U�P3хޔU'݃�Yd� �ԩQ��b�� ��c���.�gl)�qYl�+�2^Q�������	�ĦL;˨�D1�Vح,�^JȆ���޿^�/}g���T�i3��(�3�)zs��i.}����
����&Uw03ń</�H�^�6,�z�x�u�����z*��9�/�^m���ֻkI�ں3�d��P�Xӕ�N�b�5�1�ë�`�m�e��c$2E�����6�i�����T��J��sWd_�1��:���زvIvi��'v$���k��f�� �@�6�#>�萌Z�&Ti
�W��ʚ�>*��
p�(�"_W�d���^��iBm�+��p��׶�'>Z��V�`�wOƟ�Q��gޖު�a����v�ɷ�4��yA����ʃ~�t(�^�(e{��r�1�8�7_6K��zW�d��w�L{�oǥdPwyM���Oapp�c��Cl���(�#8�o���+���U't���.]�ߨ���}8_�쪝�1�<T��(A���ۙu8fH��	^�'�.���n��[�|rm�_�$;���g��s�Utԭ�.�t�:U��=���G���r���>������&.V����k%v��x��֫�)�m_7/��*b��*.V�J��8=���z5�W]4g>�;3�'mn��@�<�1qo���'pQV�3zmMj�s5[r^�R��զ(r�2����A4��7�dn��sc	�f�=2�TT�eZ�%�׾:���E9�]~O3����Ż �U	Te�f��l���W�g����bg���\�}�e�-��G<�Go}�\Q�i&Ba�3^���慳@��hhO����=�8�5��Ю��PT��YFx��Go�
Eq�bѹU��0�^��xfi�S⾯h��,�_wE�µ�6/YW-��[ogpy�j��k<.ޙU �:���-$ �;҈_+����{H�ʽ��n�����h���xn�ܗ.ӷ��}�IQ�dI�ߤ��VS�LW9w�o�`Vq����R�@�:.S&d�K�l5U�Ȟ�ٛ N&�����|�V��{!�V8 C+!��y7s��~�癥�l�����*�~V�eqpX��7���@)1=�t��w�1x�}�rz)������Խ��Ņ�^�xY�R/�h���կ��}�K[zn	���9M�w]�V�����æ�V�М�^u��\)U=o�J~>�kGI���n�[C�b�ӕw{��cΆ7����LCoV� ��e��[�����f��ܣW*")����݈��U���_��c�j���ޣGo˭/R���jAtL����]����ܻ�L��#-Z锶��ج��qvP}�5�%Mn6vډ�:�Jv\���9v7�;З�tJ��^��������^��S��3��^K��T��P$#��ݶ�vy��Oq���V��V�d��P��Ud�>ܫ~��}ee��~��~���_l��x�h�����_��< �Xp{f�S(8��Vʶ���-�:G�؊���^뵩�X�
�m�ג�||�r�߄ʤ�>��������=�~��YR�s���W�����z�O�!�m�q�=�o�!(�OPTN�dU�Xʹo�(�b�>z���̽�\}9;^t�/��@�P�r�V�Y�ז����EB����JT���\�__\�ϝ���Z���S�1
�S�h�G��׵��j�4%n5<re�\����db��F��*����
�(�x��y?{�9����;V�Cu�\1]=�`Ϣ�(2E��ēµ� ����w�sO���w}&���Ǯn�w�SB�hϜ��ӗSL���K�WK#�N���-v;O�����S�|�/RZ<�5��3�%���P��d�Em��=�Q�.��{��gd�ˆ�Cp����5���3q�q�3�7z�Y�E�$
摬Ww+����i�^Y��s�I���ۯ��),>��b�-f��V��n�W&�n�p����(/>e=H�p�g#�z�@�z����X�}0��\�u��E��:&�~&�pWR+Ō"*��+���d�[ O��nnG(��Ǧz��/��KMi��q�򮥶]/.�߅�U1T�*ͳ�Z�0�k�9@M[S�]��Y���b���� n0�K���� ��}��O6���교�m�1�㨺�b�|��x�����Y�W���_W�L��ln��Â�|w��Ú�⒒ᄹ��(�^F��ڻ��{�gy���D��+KԪ���ʫ�^fK���k�'���&8�d==K�TJ��W��oS��[dg�D /����_5��SO�@�zn{�F��B��W�W�X�<��.φ�LϬ���˔/���#<�Br��)Qs����6��*滷�^�OY������5�R~yv���j����f%(p_c�J�;�l�DsʴAkĝ�ᛱ����޻%�D𾠾'�0s>�Q*����&��=��m��q���E��/��_��5�)�p6n+�(NYd X�����k��烔�l�2���Wx��JkSF����~�l�߅�bt1�Żt�k�ԫ����S����~�$�vWh��}e�݃�o�^�ƃ#tv���jg0��c�x�'t3�`>��O3��j����G����k	p�A�c�M�R��Y��1�d��;�@���u�Y�S2��6�N�t%������y�/�P�w��N������.����o����i	��;�]+��P��_i��W�fK����!�.Z9ϛ��T��l^�VהХz]Dz�T˂�m�;�7s}���R�o��0e�5*���X�2�ڵ0�C���}��S� �ͻ����]�R��������ү��9Bz}���G���s���|�]��G�/�y벯3�2���P�YBP�����/c�8jgX�Z�5���G�UY�=	o:q�#�d�^vgWte��������E72P��;�xF�S��TF���v��~hxԖE�w�7"�g�y^��޾O�U�W�U��|L�/��0xxzf���V/�dޜm�;�1�i���;|UL\m�r�tHF|�xL�!^���Sb�>����~&����{;�Xm��ڹ=C��0Vq���P��܇)m�2����u�ڪ��S��Vn��S���]���.f��q�*��^HZ�ql��#����N��)[��q�P�'�pS�Qp�)݁m
-��nmА�-�,gS�x��ݛ{.���U3%����l�3�a�r�'��]
��=�_w�Y���)eb�2� �wK�e+��;+�����D��y�����Hi�S����ᗯY��k�p;A3�&m*�Ոa�p�s�����zeZ%����q�Zt��/F���+�6m�J�����5�YQ,��U͍�>sF���Iq�o=��]�1*�閳�޾���KVI�	�.\�seEDK���C x���F<5zH�h���r�n޸�^���E��!����Χۇ\���VZ����qx�R��GZ�Kwf�gm��d�/]jq-Z�h��˷үY�(����j%� sg!�U\�_�ՅlQuJׯ3.V� [s&"X�L5���lw��ݗ�XB��U
�23�ɼ�	SK3��ź��9���}o��hdv"X՗���x^-;;�ǻ�KZ�D�=t�LoAռ�;�W�^���_�y��jt
��}8��&ի9�S7a`�c���c���f���\�!�Vֲ�t�Dk��C������:�z0gTLW^C��<K�H�{k'w�1E��W�_j"��>[&��]�u}ch��:���-$?��y3��ܚfh�91��k� ֮�����)�0�L)B=��勩}��;-�!w,B�͔����N>�7�W>Ed�Ko�������]5y�5|m�h�qqW���`j���n ������Kh�=�ڱ��;�Z��-��ɕ��d���Y������X����S+l@�>���%DmD�8�|w,v�o%C��ڮĬ�@��w���%�E�gw;����^�.�9�'RW�E�pr�'k�:oxc����u��,鸉F�>��(]�g�0����XmܜL 7/��;lͽ��)uѓ�^��#�UK��U\�J��m�ā�/��\6uqa�M^�v(��-5��6���0���&�I���,�FY�m�ҙN�:0))U�Cz:��:̃WVoCw�d�	p�B���Ǡ��]�]��´.�)�M���·257�\0��Q�D>�~Gn�BU!H�JD�V!�N�Ʃ�R*G�ûZ�+)U���lt��B�Yw�Μ��鼆�n��<LT��y���ՆoO��Ik�������_��{���z�b��7:ՁW���ub��uD\�31�G��=*T�3p<h1�fn�P���YR�g��|r�n�Δ8�v�5׃��	yhs����[�eA�.kA(��;WX���2��U���;JΩp��9�}k2g$�����;i���,��������ɳ�8�2ɾ��uՈ�	ٙ;o���h��R�o���n���ꈳ�����Cݠ����KB�G2W%X�<�#��6����w�>+wRak����2-Tƃ�h@�+o��ljUkYEB��-b���JԪ�kYe�[Kim�T�UE*~�`��Ֆ�312�[QEUm�U-lQ�1J��E�+��PQ�Z�Ŷʪ��YZ�R������*[Q++"��Ԋ����[m�U[lU
����T� ҬDV�жŕ�J�ʑED�iB�E��a�⠍A�6��E&[���iKQ��eH��k2�Pm�m���-���m�ő�X�X�
�����VҰ����"�0Q2�T\m�*KJV��(*ZR���TeEi[X�kZ2*���ȶ�U+U+1�EAT�mQֶ��TPY��[D��ʭ�b��[���b�E��a�R���F���ڔB6��b�TY\��(�rʬ�1�R��R�"��b�Zʩ�(
ܬb�P�h����3
��V�,�mTT��PP��^^^pC�hl쮺mm*��=t���ľ[����f��|�k"��zxt����6eümveEK-�x��o�hq��9��c�3�Q��e�=7����|����;��L�y!ʫ�Ğh׶VX�����}�U}������z^��A��7�)F-�ʻ�}*�U��Q����D�>���S�)-��~x�W�2���
�9�Qq1�M�n}Nc���=g���:���_��%��%p�=<5N%�����c�~�h4�m��zg\j+ݯ��1uT#(�!���!�K���;t�	���UNlzU%[:<�֮��ܫ�mӟt~�ƃ��}�j�0]f�ɲ�ދmī��.jjT�r����ҕ.uC��������2_3�YJI���=�h{�՗�m^LE��-�S��a��X��Ab��3��`v�������sH+��z�kOy����Ir< �WypnUGp�@���#������7[���.��~� ��F[�_fZ��Y�ӕ
S���VT��UE�P3���b�
�,lW����,�'����7�g��'�l����fQ%Sw*�'C>��=X�C�xNV���)�����ޫ"H՚�탖+�t^�6f�}[���m/gl�V�?��g>��M��2Sՠ}�z�0�>��Â��r<��Eb�k8u�p
�i��J�|��'o�]��Y���z��ԗb\���OU�`�73��y�K�����{ë��%�]��P=�yɒī7��7b$���TUH�А��w�ϊ�=��e �^��r��x���"�x^����<�p�V���q?C�:�� ��5 ���|���{7;,�eI�)�؍O�yyM�1d�2b�~-���D}�U�cj|�����q�YRu�nq��b�/ͭ�ª��p�<�|_��Z��h˯�T�Z�t����373�����n�ݬCe��>�PW�T�Ѻ|�.�m'�f]����WK���s��͙�koI�P����t;W�1��ߋ� x���e���+��>'�x�W]�!7}��n�g^??Ec}<��N�a�9�ہ}�S�i�l�cY��U����&��N_=�J����H���{�h#����Tr�����C_?N�d59�g�\ް�{���Q���Εg���eF�_к'|fY��R��r�^��fS�COۜ��!E��dщ�k�b*_��p�9�z�>b����h���j<32��~^��X�5q��:��}՛Ȟ�{u�]�*�+
�v�ޗL��-I"ˊc�$=���p�x�$W�#������N����.B�P��M��JJW�u\G44�=.��
�e_[3
)�u�{�Lr����YGo�k�kQ��r+��nHd�(b�]L��C)�S�=���� S|P
�� *�5�U���C���k%v�&>~^�����$4�u˘y{��E�Pd>&��Y�W�lWYC���L}/ݯ]=�T�J�Hq�������צS�)V�r���M9�A�/����ڽ/�e�boK�v���4���Ih�X��[;x3v�5�����ȭ���	[y'<AٞZ�3�۱��N�o��O��}�=e�-).��p� �7|�9Y��(� k����Y|--}q�;�c�0����et˼59տ�IAႳ� �񧞷c3���-5E�nc>Q��O�ֵV/�??x��v��^,�	�Ò��D���xm�Ӟ51*�Ǘ�ˎ���v�5r�T��`�p�Z�]��y��zݻ~ź\���S-<'2����uz�z�IۻZ��]�	��������T�fW����5q߱��'����3s����=��L�<E�f}r�+"����U�� ���yW�e7.x��@�z}�.�<���g�/w�ꘀ�NG�)ԅ�u��w�(&p]ט�&gT#�ds�ᣳ�Y�A=;�R(؊��Ay�Yt��4�\Aھz�N�J����l�g-Z�/7vu8�MR��;Q�(j�KB ��,a���6ӹ�c��]!F������yyٻ��{�݌�{��c�����_�J��5�d&m�R���)�=u���ө��y����f㘮����Y®X�<(�A�LI�Ы:�+����MDK�e��n_����y����jbN5ߣ�O%� �z���MQ"���V�_-$m�L9W���3�c��K��s^jª��x�|�;*w����U*r�!�h���3�
���o��������+�g���~���q�5�ز���8���wCi�,�K�k����^i9���c^���A�eV��K��̨�L
�Ob�g���h�]�[\�n
WO]󳠎�7�x����Y����/uʚ�l?���j��n��poW��#�3����t赾>t�ݼ(�����dҪ�/�V�Y�Pr�X88hYY|���Pxm�C`�z��`�����_�����A�
���e���|�7�����*�|�ZL�gj�Z�Y���Z�D��͆���9U���/g��᩟u����[-!��z����GÆ�-�֚ur��6���>��%�+��ݨd�*�Q[�Y�L�-�C�QЧ�8g{ϲ��8$��f���GE�T�6ʽ�r��,�;c;x��z�T��4�k���/��$�r��k@������.��R�m�R���Ϸ��7K�c�uv�=\uU� ��)QT��B�,xƈ���]v���L�79wb~PHLd�Ѧo��w]]/D��m�2�S��[Ү��ĺ������vXKEm��;W�C���=�2��j��T�����76�9�B2��	�B��j0k&͌R���^L�ȧz6�]�3_S	�%V{�ī��_
��q����*��s���s0z!���B�$�~[N7�Wڶj{Z��r]v��џOqY���A��
u~��Ͻ��Nz���K}jԒ6rݡc��xh��U''��Eu�e��uw��p�U����@R�����3�Qh�pf�����9|��zS��Us�A���:��������������c�M!V�����{�����C>g*p�)�Un9�l�qˁL�3�#9�{y�p�!T�|���NltJ�tyo�p���f�9�E9��������_�v�ݲR�+c�ELԮ��x�����yulE�e�0����B:��~5����3���8J�l������x�w��ro�wW���auU�7�n�~2���F�(]�D+����x�r�[�z��qŹ�6*�B����?=�J��kn�vW_u7x�����}Ճr�d���]���L�J2�cS;e��wyA�t	8���L[����4R^��L9�~�Q}5Q�W�t�;�}u|"�.ν
�����Q���T�M�~��1������qǗO���P��)o��Z616�p����P/Z>���@X���{+u��\�O��5�+#����Jq����u��*w∦+Q��Xد��.�j��=��8��x�t��.�V��$�`���t2K,�eS�
��pg�����Ի�z�ۥ7{6k�k|H��b�"����ϫ�����Uk���:
��4�����W�U`���7;�q-Q�Y�l�W 0�5��Z�:.�q?0X�o�r�
���^��
�{�Sy�W7�B�W��K��	z�b�ݥ�>v�9������k��4� l�i��X�ɿg�m6��'����a�5�w�J^u�*�V��k#��O���3�3Gԥ��rژ|=�p��y�+���m�]��Pi�cƳ=lʖ�\��L�G�~㮺�L�J��%�L�p��6_x�X�������l�gt�C��ͨeBTw[Ie�� �e�8��o�к"U�7�n�����d��#Jn�=��̝����e�Υ�bY��v�R7�Z�L=���p7�eG|q~�����צ
�lnS���I	� �8oq�\�*ʻ�3+O]Z\����5ik��+��(��)<;�i�����3����ly�9��� 8tw+���q��A�4��e[τ�G���Ik��6�i>����CG�@D<ۇK��ˌ��|��j��z�����r�hS�PȢ��<�Ժ���42�;4� z��Ҭގʥq3�ǡb���C^GNU�r�0��n�6��B^�l��V;*veХA�� xz*U�#�*����x�uS]s��y���[�j�������<C>���O.��*U7� �� _�F��7<���S�����{��8r�'�py�k��/�˘yz���A�C�j류n� ��D>g�]��Բ n��h��0����T< �-�EMh�r���M9Qz�u�[���H����ye�D�$h���I�\1�,l>8�ϳlC]��Rt2K"��M�]����U�8]��=���O��=e��ђ�&*�Eac��� �ED����ގS��Xv@�� s$g�O,����~5���u����x��P�����P6$ ��ݺ�=��2�wY+̻�����ޯ?
�;�O��qnpj�U����csX�9������W.|�W]F�S�E��ub���p`]���"�7��]V�����9��q���>�y
Ğ��f[)A��P��W*J-wt��l�c�E��/{���&;"�/*���ʴ�d�ކ�4�L;��ɍ�Q�E;v�S�|�[��崼2���8�3r�����B�zU����P�Q�x�s���{/7u���7t�ϲ[5'C<tS�U~T��f��K���rv=��6eK�`kh��M�=�O��d��X�1r�g*����"U� ����y���]�8}PӅ�/l{�Y{�ա{��^�ҖpŖ�z�(]R8�ʸ���-u�k��L�b�s��>��/�$M���I�Z��n;��s]��̏���B��W��P����.�6�!��G�L�z�4����3��c����z��K�"Tx_PTO
`
c*�U����7Dyz�n�j����m��_^�fVWvR`μ�:c�S�*�28���������A��s6����N���65�X�t�_Os�2g/�8��s��J���P;�wv9���ӝ(^�L�U��WK�����*��u�`�=�W���^���(	��\�CaT��Z4n�]1u��+�<wU��0��ڏ7����62W8�Z�v���)'S�mi�MZ�9�e|%j�C��V^�t�.����mta���3�q�.�.Mk�;1{�J�W9U��"���p��!�����(�w�E��i����@pΥ]7�.��,�I��&�ڽ'�ibo_���f(:�C(n�,�(j�=�-��鳴=q`��t�}�执Y�i.�-e%/�ס������h��~f�O^5��k5����0f�b� ��q!Pqd*��9Gp����;^�ݪĠ��kr\��no�&��T(:
Ao��W�xNH�^��m�+�RgT;�n��s�|w���S>+���U�ʀ^�J�nd�Q<v��4*��b�4���yD=(W�V��+y��1i�Mρ�=.ѯ/r�{�FP||+kzR�X�d�r'��F�ؘ�O�Z�m�l��.ר^ZA
�Ϗ+��S����!KW������F�W��쉙�=]���2@|�?=�6�C���a���+6���}Km��^�Y�}Wh�n�|ۋ��c�X����z5^���$�V����O��4�.�
t)_�t:S�߲�,zy{o�K{����*�A�ڂ��U�$������R�hS��"XϢ*�P�O�����5�ZV�]R�ȭ�֊m5N>�$����W��/qT���ݮ��q]S;��c��r����V�H|� �K�
y�l�-e��>���[�+yq�O_l���j��?2V��d��p�s���L�IZ빬�X]v�\�z�-����c���D1�paq1�4_ٮ&w<TG����{�Ba[�k�{�e���+�4�y�^�_¼6��:Uw�b<��x}�Sp�����Mz�q�d�.����[�0�#�ÙϪ����J�tyo�_�WLۧ�{y]���
=�H�cI��^7�o���u��t�'h<&�][e�0�=�[Oǵ��OT���dcv�.��*/s���0z�ן�ѡJ����9*�-e�`Yס���m�A�r��u�����Ҷ։���:<#+�<�7*/`eY���$A�*�#��5��ʅO}��������a�5�eT�V|��4໚y�huCPzZU�w�T����Y|
��c�Ցgo�[Y�s^����Wg��y�y����:��S�
��pOs����s}�ۚ�H��1L*���U&K����M�2K�\�EH��_Ili/x`����]��n��Vx�2�bUq�l�V�0��*�U������84xE�0*�n�JNm�L�c��=����A�_SD�э^JB��Y��5/&�F�Y��-���Ūϑs����.�X�Oz�<�1�W��:�K�\�xѬ���v�so5��&������9�*.��Z�=m�z�y�e+QHZË7���\鯙�tXMQ�8��{7��;���j$��ɧDl�pݸ�A��;)�hU�Ok���=�tq*ϝ͸9&����q�Q.�����<*���Y�f˱�Uf�YU�\J+�V�G7�ew	���WP�a�]��B-�ҟ)�S�vZ���0��ER�`�m��t�.f��+Q��z�K�ƪ�]Z/��PtA:"���}���t�B�[�T�z��ӫ;_rh����0��~&��{w�qIY�*�Fգ�&��ͻ�yB�up�RVJx�����t�Wtt��[ɚGT�<�Z&9�i'k�t�w4��qwf7Q����Y�Y]W���gP~v��XWx�n��ez�Z��=�U��"��X��Z�mX޴e�;p�;a�|R�:k�F���#�}a�I���]����8��F����;��2��L��Nh9FE*�ƞ +(�J����ɯ���M���e+�/���;��*N�Ҷ��V���oS�]��hS�mv�K��;�Y:���t�P1L�����v�&���sSwi�ޥ��
減��`��d�7i�]��Ŗ�#�:t�Z�[��t*<;��V��V��@������4"8A})�{q�3��;��0iSM�f�J@�cyԼ�v�1lK2	�EEǤ�S�k�r��Y���L�%�.��y)<%�ֻ�tv��Eu3@��b�.v�Z� ��%<�W[��㹯�s�w%�󕌨��u���D�`?�-�Z��C6�n��G��(�y�ƾo�E��[��sW�V�7"a�Y�nun� �{���遄���d;��vAh�|t�]�a"���#;�����1N�&F0�Υ�ŀZ��*"]0u���o㸿C}��6Z;+��YO���u.�����2>#6u�i�{p�g���[��7|un�UՉ=b��t�	E{N�x��0�u�L��=�ԃgHd���śԯ���\��7��z39��us~Ί��-)�9,W1I��r��	�ox-�Gx���y�������iʻ��qi�^t�<����j�ܰ�dD��XA��gd���4s��2�J�t^$ْ�7�;x�[{Qf�֥�=}��k�j�1��8���u�:z�j�6�s(0���U���te��*��,�îb��V쭋!��8��Z\nŞ;�W2���<CL�=�G4�
�^�Y�/u�R��؊)^����j���{3�%��X��:�8Z:�KΡD��F���W&�[6�Oq����WsbG�G8,�$G؅m2���MN��]5=�n�}���^p6��&��=�F���m�m� �d�[F++
� Q��Q�aTQ�b�����LKmd�
[*TD�-�֥���J�TU*H�Zب��%��V�	m��QDH��
�J$�YA�+
��R�Vʭ
�kR�-*eC�
ʪ��ث!Z���(�mF,U*,YY$�T����UDb�d�AAeJ�Y
�J��"�B�PD���VJ�
�*V�Q��-�DA���Ak@YY*E� �PE��b�+
��(Q-�(
��e��J��TZ�ڠ����e�b�
°E�TH��VT�D���%�H��U�� R�R��d-��TZ��T*E
�DJ�*��V�ڕ%���(*�(�P����PZ�E`UEPV�-`[eB���j���*TQe@�����Y��)V�R�)++m
�c,+%����DD*�PU*E�~��_�v���A�*�jrRB��c�x��$��p.�Flr�u<Q�D��ᒙ�[�����Ρ{�K�����{�:q�&`�w_�;�]��_�5�帆��7�xث�W*#�2�1���@\u�-�^��壃a�5�#�&�׼u��ˏ�����ff�՞�`�u�R���]�qN=w��&�)�ԗ����a��
y�+����;Nr�����}�o�l�e]�N7���K8a3�u)t�`���2���1��=>� yT���g�VF���:6|σ��v	�G nٕf�  ������5)ˈO��:�x�8�]I�7��ՙ/0u�E��YM�9����e-Q��W��|�{Ү�2.�8����X�%���l%d2~��������*�z;�XϮ[�ج��)������q���׈��Z����CM�S��t��
ʡ¶���j�f�� ��K��@��\����äk���9�2)�.�oD�r�^��XĀ>�{u=1κB���KxڌG~U��8���2���5��FIu�q˘yLP!/*�c	�(�V���HV��3���ܬ���Xנ�ud�W͍��R?���nu-d����ה3�0&k��*�[���O:&z��^Jl]u7�q9wa��Z�� ���
i˼�����tP���)�g�MCܩ��21��w9\���4n�v	������ӯ��ve�O�-Ⱥ�Z2pT��X���|�Һ�ź�+��ʝ�0�W��Ye�Ƣ�np�\��H�Wy��-��X������2�+������2z�U�8�+���o�$Eu��J�Wh��}�z�^Z2}Ip�L�xSF���A��S����y���kXB�D!��$�
�;#���r��ڳ^����Z��ym�XCO�)Wgw����^�>���x��oF��֥�q�eC��9"�nnR�N�pl7&vR��ao�c����}�5��o]�	^6%w���%�&NT�><,X�o�ב�Xu�K�5п'q���@ݹWt�Y-����ᢝu�S	�̯{�p2r;�t�=\=�{�s�X�|���z����P��T� ��l����U�����~�*�������x�3|k�*W<\��L��n����L�ѫ���|�h�}<Ŵ9�����:����)�8�1�c2�?5W��%P��^�s]���7q?z١��(�T���]CT��x�Q�j�OͲ�CX]���b����� �aVR�D��	�W-�9���E�&v�}G�r���̉T׀(�Yս\��q�e��.J�� ^Ϋ!]nYμ}�¯gA�x����f̰�b���]����ڡ����؟��<��fw>k��x?�o"9H�D\�c�N5ߣ�O%� �z���M)��W�6���$c=�j��mq+�؛Ꝅ@�����K��c�w���}�Rr� ��L:\�g=q��+���!����4�r�n���]�	��	S9}�;Ҷ�{�N�٫�Zk:�w}S����H4���zN�:��Xl���߹^�K�=Y.a�9��sO>W3[�]��e��W]*Mˠ��&n��4�+�|�&�����\�T8�/ܝ�����������.�gD���t���������4<d�t7+_]�e�\��9ӯ�-Z#�z�p��3i�ʐ[�{bHTN�B�[Gp�=�,���K�������qk��;�g������ED�nHld(:
���t�5K���0^3.,K�f#'v�>�(>Ȏ����t�4�݊�_{�**��(e����n�e�;^�̃~�^�n'��d��&�-����Z���ߩe���PO}�����Rޔ��OT��x��P��ܦ���%a+�E��X��}:"�+�M�<�X gc*���lkY���1W��Tx=�g�ј�yw��@���-�X/��bx�k4wjO�'��w!�;xT��4n��j�t��v��ky؜�z�>���u2��]�n[+��i�es��6f+��ɦP���N�S�V=+#�0���x�Z�_�{�n���M�u����ܭ���Sv.��/���|7f�E��1XR�����x}㡅�����l�#ěE��ŝ��s�cd�U=��Q���H�WCfw]5�u�5��c
�L���Y����^\I�P��l3����ڂ��Vs����(yM���=�w��{|���~N��ML�C�
�\�����<s�aPs���c*h��q�a���⠩�y^y�c����Ԓ��$V��v��xl.������� p�9S���fK[�������)҉�l�l��\9E��,t9e��Ɛyw]��vO,U\>�.�V���K�E���Z(����S���䮆�'hi���p�y���֮}gjAt���Ykϓg�%0nu�,�
����e���"�Xn�vK�mc �2���_����5V�o���l1��S��{�M߾S��<3ù��tTf�������2�����X߰s_���#��"ȏԪ�Dn�-�7����Ic+`+��M
�^��<�9�E���w�]�^Ң}�p��W�s<"��gƕv�J�N��K��U��$�Eek�ܝ����jZ�ov�P�+1�,�UJ �J����u5��&�����^@zh�&�s��_(tV�e������.Z��0�S�Х8���j;H8�	wJ�
U����~�ӂ�2��q]�;~�nS���י�n̢J����n��%�z�� q�l���嗛��g4�,JbD��+�A���<&�nx=>���:�]�:z��ً{:{M�1)�<~Q�"�! �̃	m몗�[�u{a�,�\��*�p*ס�{�����I����l���R����K�1=���ײ����abWQ�,�X�>E�
X=�9�ٙ[~�H{js�o`J�b�j�<"n]{�ã]t�걕�z��e���{i��vLx��ϓ|��b�kI��������_)���,��pW�5�t������`�q�>3z����/sJH�WpBUd���uԠ����r���__<�<z'� �?�dmʒ�:޾�{�ݽ z-����Q�}wธX;�.� Xx6U=�}fq��SO���sk���G��©!�}C<pd����:NًS)�.Xr�$/;����}A��n$��Y)�: ��xzT��5-�.�+1�+�#u:�[�Y�A=hU��^S[�NCNU�S��2��ے6�6u�����$�=��#.3z�,�g_A�s���u[I��p+O��WGc��8�eZս*�Q�k�[��&	�:썣T�M���|'QQ����u�kr�YQ�7<�hk<�7�"�t��3�U/.&�>&����EI�����υ9^h�=���s����.Br�j�ǎVT���p[�����옖�b\��Rځ��G�}=�!�2)�/�gI�P
�� "����C��K �y��VR��<.�:ߎ��pޏ���)s)�%�\��ys�rmY�ln�^6u�Ͳ�W|)�T)���SU��mP��޿S^�OХZ1˘z�k���q��R�':jN�����窷�b�j~�pK�E'Ip�E������g�P�}|�j�]�K@��I��r-��7��h&�i˞̩�|��2�����v�!xXт"��ޙW�N�R��]���b�� � U��'�T�+q
�P�%}�δ�=f����V-��oL^u�te��ph*���B� ϡ����ٹ�Ht���NǺ�R�u�j��֤��Ƿ�7�_9k!�ۺ�||��ۯC�P��/��M�c���4h[/��z��;����wJqٛ���D��`����d
�E��o~j�lS�r2Wf��+�j=5�+h���-�r-����ғ��*����G�0�{�p7voVzo
���*\�r�C��8�lBm�k�b�fӻ�`Y��˛����a�v�n�/5�z�tl?Z����\�ԥ����3��2��[p06��}rF�F�>|�k�v�ǽ~��ZkI���v�����FW�D����d�9;M �fw ꉛ��x��oq3+M8^�}�.��є0h��Y�3>��Yn���^w!=�w�x\�*�������ٷ^��5���<�Y�~�,��̟>�\j|t*��U���U?fu\���ho9�昜�sڋ ��!�p�>.v1��滏��~z����wr�%;:�R>��霹�U�%^��į;�o�a*�}�eT�\�N�d�e�O��<ʯ^�+-e�X$�� ap�=@��(V���ֺ���s��3N��0*��eL�½�*rS��X9w�W$��Fk�*�g�w@���`�s��]R�t���U�l=�v]���b��t�b[ַ�����g�l$U�^˘q��Rw���r�d�����Wa��^�റ7����Vf/sp7��A{�zP�Cs�u�2�\�^R��nY5�Nܾe%*��,X�hWu+��(��%�C�gY�&T_,g��z�v�R��Z��%a��J�zil���ֹw�{l���ܵѷ�ib����_v�2b�D�8��7����p�qQ��\�*n�N64�a�t��؊��@]���`�]g��]bk��ޝVAZ{n^�S�����}���x�ֈܪ����f�:= ��e ��I
�>w�-b�ć�-�{y��3=/���i`�+q�3�m�I{ݔJ��62�A�_H-���^ d�j��x�ۏ9��HnY�=/��fnzi�in�D���Ң�R�	��1�j�E˛��̋ݞ)���Ɯɛ�D�!ϝ�;Bͽ��[6,O��O�{e]�c&������:vs��y�! �0���8��??=�4���P�w��c4�3���KW���9Cy�!o�dq���г¶o.��܋t�T���}��c�X�F�7��VS~�4��(�.�ֻ35'@��=�4�x�[���${�H�鬯��^���N�p��kċ��P�]OY�p��U���yʥ����.��y��ס����<z*�q���-��~��š�ǻ�^�e�ŭ��{�lȻ�5��S�&�B)e�>w:�[��/�v9�@3���p爗��SVal�����v���Wb��\�;o
�fY%��Խ3�5��R]��x�4e2���\A�ف��E4�,��s�b$�ټ���]ƨK�4�����;���.�Z�Ҳm��}op
�V��l��,��^�+C泩�&R�}���ě���s�p���$7�[;��>��Y����Ze>k.>���7�>yԺf_e��U{|UvT�����ca$��c�]�a�]����f�xg�*�M�gi�i�[�R��{�3��U72�*������p󨹟JKE@Kw1�2�֏f�yN�MոW�ir��5/��C27V�~�E?X��3��05�Xm44'�����ï)��$��L�ı6[ӕR����kG0b>�+��R/``� U���Wz�z�觓ʛ��ޑ�Z�%[
��[
��ҫ�.=N�!��R�}T�:������C�ol���_d�A�޻/�"�W#,��^R,r�f�<��^g۳(�����B���%�z���!�%	��c��(����_�+h�O�P!�!�Mh�%��~,n�D�Z��	�\�U�z�;{�ҹG�+*�T��`c}�N��!�Z��-r�\U���z��~;UL���^t,*�x�.�}�.��`�̀��_%3��b��l�g��cO���XQ�r�_cf����ڸ��r��_B�ȉS|�t����t�걛7�)��/�
�o�}b�ڞ�9H��t���:���������وDNF��T1n���M�1��#��fQ�2��7β��y�C��O>co�T�N�%ٛ�+
�kHSʕs�zR�j�u�S�1�p�Ŏ�Sh]zi�k��{kruoJ[-�f	/b��/RDt�ٚ��u����u�˫����|=�p�T�PV��W�t�s���`�w��۲O�S�m����x�Ixa.z�'���=���b�UR{czV��Ʉe2���̾�	�sY���v��ʤ�8r�W���V����9��g�K��:�������s<�֠��ޕ,"X46�f��u^�5�����ˌ������,�'�����ݍ���֑ҫۯ��@��u�M7���T��jD�=@��<�g���~8�7V!�g��������G�=��̽�T�s�� |f���S�.�*��u'��^��_S��m ^ɮ�MĨSr��:2���ʧq@�5���	S"�9�\3��n �<0:��W73[�oIB�U��oCWZʬ�u3�x�;�pޏ�F��|��<�(a�R�(����UɜDkR~���A�	�`�d��5��mM��^�N��9Z?-�\㇉y���q^�D�|��`�j���+h��#I>8)j\1�,k��3��������|4lJ��ذ.��p�3�|��R���QY#5����YI���W�WX�I�L�Le���n�zsA���4�]�K{�e�.�m�ڔ�A��S����S99R���FԤ^_�A|�����D��޶�]�ݤ�*t[]2uZa-W�\{d�0vm�Ǔsw�<.�"�,mU�;��C��Ր�XXe����U��8�N<v9�e�aɪ��b���I%���7��PZ���.��f+�܅�g��d��2/[+3Dsvi�pd��hZ��=�(F�a�';� ɳ�V���C]���57�;˹�V�Z�Z$h��
���flց��.yf��W"�]i4����e��­y0�B��M���9�}N��y]��O%��A�GH�3'iI�z2��hGŸ]���:�r�J�0�#�/Cޓ����JWV�hQ����i������H�����Sl��T���*Knon�0Wl[Yϰ�uE��}�.�yG0�2J�x]_P�(�;�.����5˲r�`�[��<�Y�1햻{u��ͼ3�a�Ԧ�I�շr�!e���U�=qV�������Ŭ�g����	9΋�7�M
�T�O.��,L����7;kv��e$	|1kp���Fd���*=�[rwu���ff�-@n�c	�51k܆^�!��	�wt��em-�.���q�ց8��v��}-p�Ry��?igU���O�hl��%_N{]t���D�9z:&&xu�h9Ք�ì��/zp�]�2�W�+%�L<���94��
�f��j��H�s�L�N���%(c��v¦I�˻=ʻ+�nuޑ��ȹ�T�,��;��]�w^B���H��BD6���ӛZ���zh�k2�*�����!�����.���3�^�J��Wk����g���	�b�co�]KP�ukr��vΕܳ��`4Zd�Ձ�2[�{�!c:�s��r�B��
]El�W�rp�:NT�<��(��rb܅O�䩯&�t�z_G�!àk�7��Uj��D=�|)���)���Zƶ�ж����V���-�Q��Z]��3S과R�[�j�OZ�k!�4kiH�å��cL���p^�:�ec�nd�Lk�	6�^7���!���:�u�������s	U�GYiJv^Ԗ����N��N��J	����F���gշ�_̀�}үr�ܫ�[���@ḑ�r���mԓq�!����l�X��j��R6�	8#��P���j�Ǐ���K��
�v�R����7ML`�]�ڲ܋:Ź�����3b��!���Cy3u��fR��/������U�ɳE�|�V��M�:����4� x��8�ZS؏�/�6�X�;�s�/:8���Q����E�:뚨�)���i
�3��T�'I���|�
�tY\��ow���.�M��nޚ�-�,i<�
��N�%iu'��ӓ��"�[�z��Tu����8��MpuɄ)k;ˬvSp�/��}�k��K#��*M�7@|P P�j
�Q*�ԨU����k*E�ªIZ�ʋ"ȣh�X��d����+��*�(��YY+�)EJR�X��l%m���k-�j#*DI+
֠֊,X��iDPPX6¬IX�VE����@�Q�EUZZ
(��Dm����Q*ԭ`����TaQB����
b��UU��V(�QjQQ��Ŗ��TVĶ[j���-[iQ��A%aE����*�Z�()Y-lD�Z�
�*��P���*KlX5VԊH�"*���H��V�J2*���V%ed��Jֲ���jQ���(�-��X�XV�*KKX*�R���)j�
�YlX�Z-J�b����h��,�UD�,R�"
���(ҕ�TKAaQIUQeEP�*���
��*��LI�"��\k�E"�Ī����Z�mc�̤�EkkTB�VV��T���F �QAebw��.������>=&�0���u�D�&Ձ�M�����egAw.sh��=z�ix���$�W6(�6��+�V�l�R��5��t������rW��6�>�����c���.�Wq{>����.L{L�n�
�2�dU � U��RyeF2�Nuo�\�=�z�����[��ry5�%n]g�7���c����#B�+̳[s�-�Q�gh+�
�oAY��螞��if�Lg��u�ګa��(x/8�3r���W��@�M �
l�6f2���"}���	��h�=�e��R�<4S��I�ؕzm���x�۾��_N������q�o��Lv~b�!�D��{"�}��#>��������ߞD4��]n��x�M��v��.S�z6�d�)ٟ#l�|��/躂}r&G}�_U�]ǽ:[�f�q2��
r��rm��s]�Lo�~��YG�ׂ�-U���g�J���r�c�:����;bbw�J�U���c�.kW����J������՛�>H���ԗۤ� ��M*�qq+����aO>HuIu��Ӆ��S��8S���bW��_7fe���ɀt�t��D�1�K�� %��.kU�L�[���{A
�v��٫��@�W#&�e�-ޥ^4�� �e�[��v��F+�#�>�yS�hc���k�'��n��>RƦ��oGG�uε��<D�xpF�p����Uqw�W]�f��=����f.�.�o��1�������u��foiLd�WA9e���)Q�OA��Y�OR�٫+���_�*������/;���oS�ꩋ��1���6�L�v��_9d2U���뫃�E@r��%csz.Rj!M���}��ڻ�j��\��y��t5,��pR����S��M.��&o�A�zs�L�^��&�k��%	��z�����L��:�j��;�
���S��R`�$��}qo{�[R����x;��J������%wd��T(:
�����B&r^�ez{�����{㞬��e����L=��h �VP�Д&4�%��rhJ�M��n��#��m�|:�X��!�1&xmL�{oQ�3�ע�oJT~y������K��I����o�j�?(r�Ϟ��j��ꋽU���j�
Iz�S�	ڼ]��Jx�k~�ɯ4~��n��E5����d�g>�}�FUl�ȡ��+��t�n��}���$�X\��	s5��>K�[w�#h_�=���8]�Vm'9��e\e\���l������]$��¸��W��<�C�O]G\[M*��9�]Y�s�`Y���xoW'3#����T�٘%A&I��̝�(�݉sċ���m��S-���H�驮�q�K�{�T�QA����kܟ_5[�ݐN�
K�#*�P��Ɲ��\��b*��=G���u�@��ǂ=*+z���'��KQьw�J���*��W*�Ƴ	Xy�r�� �\T\\¯KϔiR���^>�n7��2r�šF,�`�GNO��~2�Z=*�B�U��P�����l���bΰ��z���{Q���kV����cEc�\�WUd:U@���]�H<���4�.�z�N4Z�ןW9c{���r�@u��R�ا;���:ȮSs.����
��.���َQk�07�����德y�^�z�Ƕ%�d�g�$XT�xg�=tk��F�^�ZK�{�H�\Я�غfEқ�*x��N���Nu����֎�na��\VS�2�� �L W�o���GMe��|�ލ���6�ً)*|UW��c��}]�p��w���Х8��hud��pJ�V��6��iv��v�V���6�Q�j>���yH�ʫٹO=p��n̢Jn৕
N�K瞨3*�LגfD��e. ٨��aN�U�e"y�:f
�3z�g
N򋋅��M���W�RwrJ�I��m[��[9���u�g}�j'�;V�8o+�|������|�׸�i�ƟKpwNY��L����z���}�$�s�y��듹v�+Ԟ���Ƽ%r����@���5��L�|���6d��4��^��8'���e�yT���,���O���03H�x��}t��\����K����jT��i߯�k�>k�^j *Eo��vt��{��)��҆S��*��=��Mk���}�Z��}����Z�|zj��{��涛��Ϫy�����z���l<�͜�K6
\yWGZ)�^��^����=�S�����y�+|�ѬZ�a��^�U73�3Ϝ�ǁC9KE�{�L�xa/ꞥJ��������G�zh����w{�v��{��XwRA�T������Y�IX~'Ń�d@]R���`�=��ȼ������s����iA���k�cY����5E�8��꾴}f�L�DYq�%�����d��7�����i�^�#�S��T�59�eM7���O(�jD��h��d�4o�fI�FR}�nx��'�|%�d���OQ|���y9�F�eN��S�.� �u�FK({����5u2�n��`ՠƀz�\c��}Iu���:��x��g6Rs9�S���;ؽ�'{=��Z�</P��-���
⮦�Kq��	;vq�$�¢!��|����ӕ�3�a�IE��L�(˄d�����:�iY���y*����է�E˫��r����;�<c�S����O������[���N�koMN}�A�]���w��Q���Ug��9M8�(5��FT�W��������T5{sN_L��pŷ~���W�1�Y�U��W܂뮢Ӊ�0p�j��~�˥ok��j�I���iW�d�v��x�;R�*�r��(2��Y*�YJ�|*�cE��p<7Z䖛o�ΞpE��L���=kI�ʩ,��
���*�*z��`t�.���^�6w����"��v�os�~g9zY~�2�d � ����<��w��:�������R��l��C~]�9ϩ&<f]d9^>Fem���[�F�ǀd8���*�nnR��d�vj�"���j$��Z�if�Lex�Y]���(xy�d�e��װTC�i��ٳЅ�ǃ�������0�x��<f���7��஭�[G���&�剞W2_�0l3��V��W�z��� g��7�1��4+�z��9.��z�@ ܶ:�)X���˘��05R�5�W�P�0n�^� ���B�; �KC/+U.T�.#��_j��E�s���Q �^o�n���]ֶV���Tk.�^U�o+)�b��c��gJ��ū��\n��Y[5*g]���Qq��ೳV��czi*���1]��\����}�1��7H�>�K��P��:Q�+ד���~n�Z���@��m����S��6��9����5nR~��S�U�B���x���t��ݚ�̼CԜ��
��%W��}7�E\ ��c����GpL��D�B������{O��!���
��6���k�U^w�T�"Sϱ	s.�b�:r��u�Q���(}�;�	y�/�� �F�,p+�Mq��_]�f���`U=�9�*jW��[s�9"��Z�+�}[�SNҘʝ��*r�!}@���]*����5�ֺ퇽oN:�� 8���鼼�����/LP*���*�T��8�ҩ��.�r�d������˄U�:���	�Ѡ�I6n�����W���b��ӳ�9��J�^R��nY5�N�r�5��x[��g\kӧ�`�U�Ɂa��{��l�w��gG���ڨ�8E���]�U�uI{��Sq"���7���/��E%�<�{���T(:�Fƈ�{�Poa�e�l�Ċ$��L�7F�E�_ p�����V�SR+y�}r���]*&T�ԫ7�z'7QԖ�,���f=����{*����Ej����81Kڷ<�_e��wTYPZ��caS�r��wt�vS}xgn��4���Y�׈�@sIe�ϻD9����fjc�޲���E��3s����4�v*$��Ε����'w���ܔߴ�(i�d#�m���5c�C9��o���ł3�2�S��[R�a�s9&e�5=\�=�4�z�g�{�}�۽~P��iYxj��G�J��:�b~>�2�����2�;�g��l��nǙ����;�u���~���g�tg�5r)�طi�	���)��֮�Īo�v����p��Z��Ćo�*zjk��n��\�ފ�����4G^����痩�ܒG�/wKH�2�R�w(w�؇*�1����E^R54�.�[�ƒ�`��Y�Бm�	[���>��5»�WWCY��<�8��|�(���u��^��z�{v��ېA�s�A���ܻ�C�w�Y"����
�U�� �h쩚�~��ʅK�	{HW�y����n�9�p��Y����ėJ|��IV�Yl�>�<���׳f�~J��ޤ��w� jr=�5��:�=��<:�iQ"���ꖼ�hWG:�\��)��l����9����.h�T#���9lSp�o>��C�������P�]��bf3ɦ��7�I�>ɷc۩��!V�Ǌ�gV��������r�K�!G�|i&�z��gQ]*7��5Ȩԩɉ�v�`�rD���޷�ws����p���g*���\�^�/�u�,![=Բ��O�������U���j25ן<�O����}�(_-�$>6[!xp��ڷ�Y\=�׻Q��������>��|���S�z�FV���������U�j���t����7ٓ��S�j��{�v�7^��1Lg�\��ͯ����"r�n�n�%c�F�o�p{�/�Ґ=�ǮLW�M�ܲ�<X��2�g�kػzb�o�^�ޔ1�6Lz3�ǯ�4�×�Ej�c�������X���ej��c�+��ORߗ{�|�6��&���ķ�~v2v�c�Q�z��1�-����}���_���fU7_O9�n�^�Jg��b�Q��>~q��{J�<�7�U^�K<�W�h�ND��E! ��7Q���Y�L϶�:�'�cu��x�����TgZ�NkǇ��C��%0<�㒖*2�-�h4�[�JWf^|�}K�t���L,�\m������q��ӆvǏ�GÍv�ٗYQ�V�EN�XƵ%7���<�E���9�mw^=���zѝ֩�eP�^�'w����=T���1z�N����Z�p�/�[a�̥�^�&�xk�vq{D��}4N��ف�y4Ot�<����/ϋ��b~v�=�_9n��b�t�S��������Mé�4�����WB8߼gI (�uw#[ֺ؜�ž���E=��E&,��j�^.R��ݓ��������	f��_{���Z�Щ쭗ٯ�~�ܢ�k~�Q[p�3��Ks[=��\�f�הӞ5���mVs>�_l��M���QjL6��(�2Zq�~���%x�܎.�������ע�Z���n.�\�f8�Iϱr����5T�}�ۥ {J����1�".�ˢ�׮���%c���(?{v=��Y���s�{���p���ڌz��5���_`u�cw��QM��Z:^����ke�[F+�u����Yn���ʜ���3P����"ۙ]A��|k7�H��1݁����k���OC�a^����䲯�nli
�I�c̛����j�QM������W֛&�ޭ�	����%����{V�d���F�X�&=�xy`���:�WO$MD+������#��VB�9U�o���^_W�b�xԿh���)ik|�ޮ�#^;�m�`.O3e�_/<�!��g��U~ǳ-����3ʠ����;�cR~�z���g%��Q����ߋ����K��� �6��nvjd惝�\Y�S�����Rv�yS�+��i|1��e�g��'�^��jUyN�nng�y��ל���5+9ۗj��@��Jzn�;��v�9�KN���������Lsʚ'�s{��덨�l��.���wٖ�Pxm]�D�Ur�Q|/~�z���T���'�٨Bv���ϖz�L�|V��=j��}��*v�C�wy/I�_M$g�{���NI�מ���]3+��
U��
}�k���w�:BH@����$�ā$ I?���$ I2��$�P$�	'�!$ I?�H@��B���$�	'� IO���$�䄐�$�	!I`IO���$�$�	'�!$ I?�	!I�HIO�BH@��	!I�	!I���e5���i@��!�?���}����q�CǤHJJ$P�J���ET�P*�HT�B��	���"Q62B�R$T�J�	m��P$)FZQ�{Έ{5IIT��R��"��T��)IT�����H�{JN� ;�:4��ۍ
t(��� PM��b�n�UZ 2J�-�� m��c]i��AM2�#`Q��t�h�#�:tN�;5P�2B�%Q(� �    &�    d    -e�v��i��T Y�
�ۺB�(�� 2��յ�M�B[5��5�@�4��ie�X�
T"W  �siBR��!3�I Hc-�iT*UBTU� 3��F��A���J�A3P�60#m�٠�J�� �1�0R�*�I
ER�bF�5+l�E
�����P���lY(��k(V�[V�M`�jB�P�\ 6�fL*�P����*J�m�� mMTfU)@m�p��D%�$B	AQ-��cV��j��hUST2y��(R�)�J��Ѡɣ&&�#bh�`�{FRU%       EJz��&�3H��h4m@�4 z��~%IM     I��jc�2b���$h hƧ�?SPI��Х(@��M2h�`�8�ut�*ua����ʰ�T1��v�ZZ�B���D��TZ����c� *���4B(*
f*��TX�+������(.�9Ad�pEE�@��EQs��@�Ed8"*��~X�W�{����n�AEE�Z�k�_-�.�*wC��1�Q	/��?�'�ޢ�Kh��W��啁'�:��Ԋ��a;�F�j�L�ꬱb�Z�J6,ix1�B��vJ�{$/!�,Y_i�)��k>b誋o3 �I$e"2ŢC8���ׅB�Ua�$�%�����Qf�6]Sۢ3RX�P9�ܣ��]�2K��l��G6C6��EJ��j�(��i��;���BBYz٫�ykdB�.7cog7=w����nܭ��m2ja�a���A�m�x�ȅ���$��4k�4���`ڹH;a{�~���an$�"ksPt����S
�ː`�yt���vcmբ^i��z�yOn mK���Qi�f�n����p���+ܼ���Q��CCjPH����qK���ˊɏ`�Xg4�u���M��Aͳh��.e�*պ`*H��R��h���U9��B�Mncl�{���1	YP�z�`�3sv�f8�ɴ���U�Ty��C7��,��k�0�P��wd�iMXI�ZpޫDe�t���L��5���oZZ����,Y�ĆLi��M
2^�b���W��(�@�ʺf�)Jm�if&�3�c!P���2�� �M�����9cL�gm&�Z��X�YA���e�)��&I�77��K)ܤ�P��T4I2e�3a:)]�6R�R��5��!�*5���n�#�J�~e�cU;U**ŭ�ϵ���j�J�6a7WF�b��yq��n�Q��.�)�Y
ܪ��7`��"b��h����{Yc�"%#Bޣ�Ε���ڿ��LWi��?�3n�!Z�b;���q��7 %�N������U]�k�i��A��&]Ǧ��X5p�J���i3��lPL
�X�Me"v�'���b9�J����q��)
R9t#�m��,�Y�$rA�]i�&�1?�����{m��/s�Ef-e;l66e�-�e�
޼�/q��[.P��S����)��Y��)��zA�b��h'��Լ�w&-���8%Pt���M�2���ޱ�]��Jr�ʧ�)�j��`��B5�F�@;r"2�l�@��l��w���E���<fa�Y7qb�qU㖰Sw0\TԚ��x.14�yYI.ڃnT"�J�d���%4�fؚY�X&�:e��NU\9l�f�����`�WX��[��T4�]7pHuH*��a�HZ�;2��{a����7�����T�*j�%A��W�n�#���d��ˆ݄�G[p�mS�yB�U����5�!��Ѽ �����r����� o���	�ǎ�H �fRIP:�EC�[�f�e&�FCx���Kn�Q�aR���t��bw1�0R�'/eE�(�h�0���SE�+��8t�$K��Zp��ȁ�+Z��q1V鸝L�܆���Asw$qVլMm����憖Zm���D#!h)���`cj�d����m�� ǅ5�M�����r�H^@d�`�i�#`�1�J� �Ţ�7X��:#l��h��e��)4wuHl*�@�Ԡ����@��5��� 6�^)�u`̤E7���*�`�, �b����ˈ^SUci-�ܓ �`ۡ���/Z�ڍZ�[bJ�u5��C�2��HY��Й����nK.fSCZ�xAj��{���Ƒ��75lŴ5�w���5��B�jK�%P�����$��Ը*;�sv��Ͱq-�򒣲Lw��*|q1��fTp�.�l���#j������bz�=,(���ؽ�re���,V�%�v�a�E%"g&YJ�}*J��#w2mЗ1f�iZ�(U�#�mE7Wf��Z�š���؜���N��YS;��V���J�3e��mee�z�	�P�U��la��dxaܼ7X�i�J�&ޖo.ꆜBe�u���%$��Y#��0�17��:�8�Х]��e*��G1���B7�T����@"��c[�[M��cn�|-Ypn�O�4��n�z�f�Z�Vn`PG��F�����KQm��C.�e���²�Y`
D��-�9y�W,a�����l�R��1�)Ր��2n�l֡ё�ݢ���)m�^��s,�'�o*�&�ig�g|$������P�U��V��eJ��� 0Y�m}r�P�҂��6�'�o�2��6ʢܖW��jƑ�B��Ұ&���1[���Bd��nd�y,=�݊);��U��6�n--��Q�,�k$*i���fP7P��)U��NY� $��Y���0���6�Jەd�gZ�ɖNV�U��X�r�SR�`�eϕ�,�U�"��x�ZȦ��,i�36ܢ+hP)���7JqY+T{k뽑�ҭSmʃl��a�z��� ҆�FH�{,���fۢކ/t,	L��2���`��ab+�/.&@��A��x��&M�xJ�rvLǐ,j}��ac���ˬ�H��J����*A��SZ��� "[�]�;vn�9�FT���u�F��{Y�h�n�K�yrB���b�7,R�U-��#A�t�M
Q2,B�طjl�l�2@�1����n7W!'5�#Z��A]<�Y���3A�����f�Q����k�b�e�ͦ�Vm���vM��h�֮��o�#(]J���f2�z]8�%�˩�*�$�Gd��t%J�e���R��KjE�t�°���v&8�+��q!�Z�ݜc2;=�%��Zݘ�Ěг2����R0�t5A��ʕ��swR�u�$�j5�n�Ӈ/r-5o&f����dXǶN|9)Ԧt�N��Z�5%$��Rn�-�2���}uv��cѕآk)AW�$'%����6m)K�I�ݢ�z]e���d	�ݹ��	$|�j�aϯE�C�`�2�&3f�wONEd��N5��{r�0��$��1'�*n�*��MKFo��U�Z�܏urBr�^�z��Qѭ�\N���x�ѿE�GG�7r�I(-!$����ǚ��Ɖ��&�Ԕ!���r���eP�*n�y��4�Yٗ��j��n�̠���v�U��AJB,'��Z.3��Y0��`�(޼w%Zd֛�(gлsL��%�T� P�N�t��f�bm��;c�*�N]w��hp*�$ŕ*�^����Y.�#�H�.-H�#ne�(�X�Un�cq�u����ө��&؁��E���m�GT���*xۦA$`�5�X;b��F��IVgy��7nfɐ�t�
�i���f�}L��DL���d5%�ч#؝@]��y-�ɂ�N��i�"�\�7�6�D�ǘ��Z�\�r\)�on*���j�Sۛ$��9���dW��k�����G\���٫.,6�dU��[L/��<2�^ڞ���{ΰ�)��H0�9�� ć�pc��4P�����ݭ��k'.��n�~����۬V۵Ͷ�_&��=��������kj�8LR�ON�7g;�r��[�R�\�<���ݞw�L����rM�`�����bm�U�_
�^=����z',}T�S�F�Z�e*7�+{z�w|���l\�x��E�0o`��[�����8�ji�W{u��_V���Xz�4��p�w%t#�j�Wo�L̾��:�n6]+�c��(f���T߻��[�lU���h ���&�t1b��O�	�í�:�@EM�Mv�9�^[ˠ��7����i��q�UY�;�K	���j���3:��|徼U��-�B3+��ʳ]˺�E8�vz��}:�% p)�W�$��%����.�_�f��"U6�s)c��ot�	�Сݕ�olc]�L�B��%�"�vgu���%F���ӽ�ƽ��w��!�z����]E Q�\>+ ��˖�n������ǙH��I;af���<�H�r�n�Ҋ�}�O�=�]^9�q-�h����{�LrǦ@�i]�U�F���#\�%i�-�C϶�����j��-ouC*Rt΅؍J��mKUt��g��O{��qw[啯l�)۔q�n�D�d2�6�*�1Ki73V�ʻ!D�cQp�G
�g��\Co�n�1�᳃��f���gW)ko�᪜�7Ddb藈ma�	�δ�����n��fe��炉o���Ѡa
0��Y�\�A:K/AM��Kj=��Hw��?y�����E�+��
�z�0�]�nY�E`B�����ZZX�|p��׍�w�8�ǆ��؛iM�S ��n�o��&��-�w[�{A�`�29���+VZ�\�DgPH�2bR���ح�p��W�]�e���Z��hG��+6ٙ�	�A�ʛn�R���2�*.�˺�oA͎�����k�6���58D7&db3!��ď|*q5��w�XU�6�v�iqIr�9��˾X���'����;1�,ѷ�X�="��d@D�������֮^�=}�J�::�͍��̹�Q���Bb1��nN[�ADv=ͰJyK�]>Ь���.��*8��;��Sy"������eY�ά�]�8����n�v,y��MJ�R�@��f��4�O
4��D�s^��rҝ�B�t��%ƦU�MGt���㽛q��p��Vf4jJy���xl����띹G��]�a�������6^>���9<� <˔x��voj��<3�]O����E�W+���&����TE�3E��{�#Zڮ���\���r�W٣�,���'�C��ە}r�bj�ͥb�GՑ�bQJ�uA�D�y�7LW�y��^!}�+k5U%�[#J7���om�5��Yس+"�0��u�GY���v�]+�)��nD�`Z�:�\����j.N˼ڥ��}�΢9��u�����{
S��p�i����]=��E8�]����~������]���k���&�p��e6�A���YY՜��}���sLY�����X�	ueK��%쬁Ŝ��o� m�yH�s�﫥�iބ:�-�f1��k��
�s��C���Y��ك��"[ϓw�Ig�]�d�2K��kY�����y潦�h-�	B_Y��� {c��l�C��!w�����.���WYZ����GFY١`�vWD.Toz���sY�8	`� ���k��봁��{k���+/���4�+v���=:)��@�Y)o]!�H|k�6ff̹�O;o���2�Y�.M��%$�dy�ob�$R��;l̬M��[�p�L��	�
�	�<4Y0f�6��ܫz��nvjSgjO��S��/���W�S��;��؟i��0A\+B��V�!V�����S�U5��ע[#"t#]{�w���ۼX�I]����|78��)�-յ�0�����[�5����"=S=��ȩ|�;��&�����at�ޢ���nYf��t����u�*��hN�PFZŤ����TO���^�7�O˲�1��t��\=��ri鷁s�ڰ�R��ΠK�1����a��>�,u�sH��)��nAVurOLk�s;z��sT���]ij��Vs7��;�&e ګ��l�3^I֊}߷�nB0�P�Utɝ�%�j�6u͹��,�RF��[qa�� k����O�uG�j��p6ku��䑦8��W�G�I�FnS�@��eY�o�BF_m��K:���%�ͤ"�Z�pPᡓ[lYw��v<���z�\]b�v���$|ee�s�l]�Dë��	�Z�$��=:��+d�G�w��ɩ�es��7�C�Yxq���Qs�^#�`Vn�}Ͱw��U��i�7�8��ۦ@�}�V,�������'�q���҇ɖ[*��J�ȱ.��vr�1�9,������ŝ;��u4oFЕ����xh	����}�~t� �U�9N�/4�`Xx�S�N���;�d���'u �n�^WY��I��ʍ� ��z��ח�aB����R�������% 	��ݛm:���S:çՑ�w���qәd�4�pV�6uy��}+5�=h�.��W�[cNe�ԛk*s6�
mv]Y1=��çY�b@�ބ�*���EV�xզ�6gC4u���{m�t�{S1�m��42�qY��򛽧º��{��89�W�� ���Fgf�#�6���W)�\ٽx��.�6Mc�L�{�DŖ_nS��e驶�p�YZ�Y:pr�>̕
��]�XH�֕��k9n��ѹ�m��2k�!<��tޫ��M�b>�M��b#;=u�Q���b�;��)�����;�xh_�u�y5iؙ�"�ѝ�Q��ίQ�#�_o.�Ljm^'
���lȲ����90�uĝ[yf`���ΙozC7��x�[W�0��zȆ��j���6d��whG3��tq��w�g	tX��%��-�w9�+&'���{������r�f�:�]6[�OM;]�m�(�v��$}/Z{��H����E\�v��zw�vo+�:��Yle(�Ҹ����Qt�@��޼DK�{$;�  i��w�W�G��+o6��`��gskz��OHs�+�eB%��F�$XZ+�9��K���0K������/��yS�I{���K���Z:����#7�L�פ����>㕳������ߺv�Y�L�zf���m�A���Ŕ�<�V��Gmk��rm£m�m��m��m��m��m��M��m6�m�S~���|:ڳ&�}X�n:���m]��/l�OTv��#C��q=�nm��H���+�f):�MOvs��j����Z�)�˃��(���*�!� )V�u���I��j-����"<3�^TtcKOf[�'�7�=�e��^��Z$�i�Wi�زsLYk�P.�/z�H�£������ճrf�i����c}9n��he5�۪��ETT^m^��E@VUYPԶ� ���2�v_�q��������v�ֽ��ۋΩṱ����}�	6VαV*��n�ݠ�ΕwŬ�ܶ��4�*��j�;x^��<M�$�#�`�Lʺֲvm��::�B}�1,�U�c!}���;�zD�̼<0kw��r�R�V4+@Q"i�wi�8w>y����X6��A�t�Ė|����]p���h����T�rH�}��nͰ�66a�Q;ݡ�;�]`�|:�"b�&7J���~�x
,�A��:�o�C|�!�E�;�,�eg���	^I��N�]#���J�,T7(��D$m�c�U�X��\�\P�%}��ud���*�ۙ-��c���#��L�H�T����2�I�.����m��B����j̼6-o8��ƌRv���k�Fv=���C�ݼ�V���r�ou9�tJ�m�����+lіz�U������J���M�f]�V�5j�(� z,�̠�%d�q���۫�UG>��j�"�0^�
�;��%n���8@G���*A���|)u��ܥ#yP.�$xEU�U�g���F�d��#nA�c��Tޕ��<���1]"nƃ���[6uT�ty���8�ː��/6�`<�Ұ��[�Τ8���.�V��|Y1oC����<pop�x���qo�u3qI�A�I\ޏ��B=v��M�e^Gf��x���1ڴ�2�yf��#��v���lɩ�#v�� �
��$�S��mA�97�j��3����ᯜ�
��ܬD�0\1���vFZ&��%̆	cNbqIJŜ�����Y�8��>*TJ޶�]���W�w<���8���(��>�&-��w[�8j�wK�������K��v�W��Eӟ`wQhX�G�U�W*<�2�V�D��`:� �*�iRU�C6R���u�N�n�Om�Fa�rԏlK:��IC}����m���qc��#�W���X���.i뜫J��C��]��ڝ{,af�����33�,�0�-flD1%�<7�ú�d�)�n���3l�W����U�X�b�����l,<!�sj�T!�VUfcmD(#�*`Ʋ��\7�{Wҝϻ���anW!�D�
X��l�k@ٹ��h��6��\k�6��a=��WP��������/�0t��܎If�u���5�fCs,�M.0�.�^�\g�7!��aX_M
���s,IJ��:�43�s�@�{}���G뎶�>Q�A�ø�o5��u�U�Y8ٗ�&�)�1ژΣ�r���t3��Iեݝ�,���sˤ�w�S̓���Z�R8)<��I�.��	����hf��z���m9Sr�l�i�ٹ{�a��#NaQ�Ot�͋so�Hm�E]W�j��=N���@Sw��v��̌8ܽ؃j�r2���7Y��M�ɋ�J/�Y�����Kg	�Z9��M!��V�76�4��:�fS-���d�e�"��[��5P�i��w�ػݛ��LA��ظ̖��]֑rp����͓��!�����|"�{6���Bp4�Cl\�l�e��Xa��CM�M=2 5èKἔ�M����O(���
���z�.����`-�Ǉ��$�0�_qm�z�3�'��@p,�Ի�`%�nK|喫��=ܻ��oL�e�5'V�wt�e��\qϱ4�֝�U,%�^�m�ƹ�}P���U2�vWn�����Gf�g	l��2�i����&�-t3(�M�.�Y��F��x�om'G�c�P$�ھ�T�G{�)���B��2I�}Þ$Nд�AJ��Ȥ��ݧ^֜d�k��9��ZHZ/�b�W�i�ܥ�����W7��8�p9��[.;��:�<��F�Nݺ���+	wG�8?��ĬLw9�����-c������A��}RS5(������4�)���:���Gא���6�(��X$��X7NX�Ճ;����gz=��y�z���\��ɂ�pޤ�L�zQʴ�*n3��Jw�ѽR>�{R}v��ޙW+Fms��8�sT���D�{g���e@�lna�js�+��ܔ�X��Kǧ�f��Ů�C�z���f�Z��lÜh����z���D�I
�@���#1�˾����sZ��`���Ss�� ��vf��T�n�u��˻���x�r5¬7!��.n���vq6���#�TjAOY��45�oD�Q\�8�Іno]�ڕΧwCï������0vqY:�'�Vꙅ W�н?8d�ۚ$�',c�BCm�]�'�g��E��9��
U����>�VuGh��;���Et!��N��gr�Љ�XW"�֧ӯ�&g��um�hW5��3u�-i��y��U
I^=���o�լ�u2���[��Z%ݺ�'�G[|��,��}���ڬ4�7 �σ�����Ɩ��|��7� ��b=��T��.��o�x���F�7�u�/�v��b�f!E������k�5]w0]��۳Mv`��)u�G�2����w\[�Z���¡�\�-o'u-A���2����g�,��Uu���G6$���ya	]��m�&$M��9OF���M�փww�2���q��*�\��k�������HNS�ݗ���`j�٫@�cwn�S�pR�8�P�
��Gx��er�8g�gwȹ�݌�JY��W�$gv��R�9a\�5��\Iʴ��֐V�X�wml�('�ϱ$i�d�����E��1��hS;>,]�{�kt.o��[���s���Xb�r�I��[��L��]5V�ܱp�Ѯ�ƬJ��!}�Ғ��+`y�2̝4�4�c5vv�H��;��v�X;s6mw[�}A��FE"o�G��¸�7�U�@������ogfp�E��c3uɜ�T�]^��a'Z�u|�Z6KF�䁘���)"�ߠb��F<ƥ`�s坦-��!��>�����w�WM���������Z�;.-����c����f�V�w�C��n�wvi97/Do��i�gX��։���a�`Ӌ Ӗ��J��Ían��s�J�(
��=���+\��\�fr�e��oG$Ƣ�嫔tEs�0�^�6lu�k�]��i�J�2��ȳI�Q��Bj��Zf�z��x2�ϓ.�G���-�Toi)�1�.�b�1 B��I�n�ise��ٍd�}�*�n�k::�2�Q4f�����ԁY�4id�0�8]Z�Vb�&h�����&�H��mb���AۮRv���#�{��x���tIٺ�خ���阙�+i�<���S]v�Gq)���zK}Shp٭+��%kE#�7rG֨ھL�es]ιm6;:u.2��@��Jڜ���,zgPCU�ڎ�u�j�]��q��>��FK���Ԅ�}�k	_}B��u8���r��
2��ӹ��Z2;�>�r���i�v ����,��d��]�_?������~���b{Q�&��}v�A�3�r� �;�\��;��r+u)�����U�z��,���ُ��)�!�:�y8����V���,P\&����t�Y��Ob�B��R�=$�C�/�3*/����8X[]+x��v�v�eb �]T�:q��`V�-D/�C@�C9��\������̸՛8�ԫ��|q�>�Ed��(����<�N�뭹�8��6����'+�R0��,��3�\����o`�˦�F���%fǳ����ԟ>�\o�՟T�k��[�K5\!8z/&hdk�_+��u��n��G���80�9�vp�~��Y��%�z����,O����s�3�3z��9�V]x�Q�'���G[��V��ʰW�iR��X�(�m��1��U�lUQ�h�(�P�����;�������e��,�e�FK�̥�Fm�2�*[V(���Q�YR�6�*��6���"1E,�h�.5EZYE
���DTF�hQ�%LAk��
��"��FТ*V�PbS.#����IHbZ�V�-�J�J2�a���}�n}���w^󫞡�qH$�w�7[���*Ԃ�����7�9�����0��|��la����#��*������H��uD����֝������:���v}�W��<��s'�&#��/A ]�B��/�O"�����,����|�"����!�,����^�ms����đ���W�iˋ�lo��,EG6v��syȭ�=N��_�N�=�5�N��n��c}�����m���?e!�Hd�dSㇳ-���w7����J��{1�5�s�#������R�tvMB�w꺠����K^_>Zl�5��sw��P�!؆Ƽ!y<U�Y���?��0��f'�0�!�ۏ=��}��\r���ݭPS��rj�uqs���ɽJ%:M�k� ���F]ڢ��r�;D���}������x�>�l�E�ҧ��jgM���]۹}��Y�i��_nO�|�:Q��O��#P6�:�m�{$�6G�ZE.�
Vn���/V�������oN�}��E�S3�״�=z���N�����}���1z�����AJt@�}}r�],ɝ��ۃ���^=ħzQ�����1�x�j�-�dx�_c��a_��]�U���E�Xt�Uo#N��㇈�_j
F������_�p�_xRx�k�bB�]�Y��:ͻ�O�Vs���7����__�g$Er��?60�:;l3����_����W-!�i�h����(�F<��A���?^E�^���Ηݸ�u��!����]��+:W`�k�k���b��W*��7ww��Qg,n�G��8뺽5Vx�:~�C�E��	�<t�d���03��w�����|t��.�i�1�LzK�y8�9<{jﱳg����d����Xа�D�-���&:������Bm;#��C<µ�������=d�GN�9xk'{}�P�t���h �L0���������P>kշ�@o��0Ѣ������s���b�1U��
:��0a��Q���l3~Xa�Z��Vp��h2w���]�{����V�w�Ha!�'�L<ˋ��UT���_�O�޿!�}�
"zї@﷯�i��yW���(+����g�"�����(=[f.VO]�j��r�8�'B��J�ʧ�,7��L��E�i��d�t��w�q����=�2�{7�I�Μ��f�s�	��>��}�ƫ���y��~\F���MC�~AxN��yw��4C<~Ԇ�HY��4G����ee�t˽	���#�Ҹ���Ǘ�AoN��)C��7�}<�毖��!k����=�9���!�򪮯r7�xdli��<��ZwP�h��+���ׂ�qsR3;+}==S�?K�uz'�z�������4Ӧ���ӽ{�������l�-2�KA�.��^_c��G�W��Ӧk�b�='o�V��?����j�5�s��,^y�=h}���f�kH��4<���i:��m����xD!h<ZGZP0����O�n�yU[�x��~���s�:�&�e�����?BG&g'�U"�q|��e	[�Cr��"B�n�r�9����Fv1��N����	��?f��#T�Ϛe�_h�K��_����!�S���dig���N���k�:�~�W��<��=�.�>���\FFW��fϽؽ��޻_"	��DQ~΂Z��|�>����0�Zn���2u����L6E� ���7��~�W���^���̟��^�����KAd_�vD?MC�"��j��Kԙ���4�r������j�PF�@���yY�bR����~��d{�a��P�����<��C�A�$����g���c�#L<|~�CH^o��cR�8g�U����\�'H:@p�">[��,��p��ҫ�t�l�)?l���ۚ-R��pߣ�*���8�
Σe��q�PV^�ÚqT�8��}��@��W.�0H�KQ)�u*�W�g�U-(ܦ8�!@�b��n%���� Ny>v�D4~e�ץϼ�t����V+��������~ZF����di�����S�og_�{
<}�}�!�qZ����i~ӑ}5<�շ�f{q��}�{ޔ^ 0�*k�ð+!ݏ?{Ov#�-"��ǌ?e�����GO���$�J��H����"��X��ϐ�Ly����UlA����*�~CO�����8��'
�*x�>��A�]yq�W�At�������) <tж'��K���j�1}�����+5���;TC#�,�X���yf�q[Fw��/C��G\�0�3�]�
�Ol��
��w ��#x�=�${���T-�%J�:�f�{ܪ�MR��S��r��?O[��ӧq3]�l_3�E���f�o�kA�}'�#�e�5�{��B8���|�z�߶�(���y�����+��\����2=1��4C����?j�O-7���g��G�w��2W��|�;��:��"~&��Zk��dNﷳ����S�Y��Ǵ�/����ܦ|�L-��)�ٹt~�^<e&p�)i������
У��NB�}�%�s���!��t���b��2\���\��#�B�k�#f� uy�[�aҺ��<��B���+"9K���'���y��B�.7W������U�p�n�^�mǕb̿<^gX0��Q��B�q�s�J؝H�_y�ff�yrY�n�T�.�����րă�7�z�OO}%���@���C�¬�~~[�jbe�BHi���u/Y׫2��L��O�-�~\~�G�a�� ��	ޞDӇ>�:
7�E�v���m[�n��0�>�[nvl�f3��0������yq��#چ�CNK�;:P����r(�F|��kXG�_��S�9����Kݗ���y2�}���?P���f}����d���[۷Č�9�n��5��~f�dq�BO0�zϧv��s/�o�a�FҩP?|X^�H��U�=�-�'�ێkK�<��s�����g�fo�iۄ���=z^/��Fz�]j���6%����&�'n��>�f�So#�p[�u4U▫�Y�zp��WU�O����)aC
�<�L��SڝX;��V��e]��?��=�
L�6��<t���l�x����!_/���9�����t����g��q*��C�& ȇ��9�:C,�U���b��̀q�<S�,����p��p��p�O��(�<���-!V���(��Q;����g����uo�"y0��|��?wY6�:�����{�b?JW�H�Ǉ�C,y��1���7����4BK�x���!�˶���Y]�Ҳo�o�����4DHi�¨x��23��u�ѱ������5�&�8�<��j8x4�R�������+Š����I`���&R�	T���a�v�q�Ĝ��Π���k�-�Ö�X�GUAFd4��p���*H����O����!�l��g1}dW��m������8'��V�`�p���.-#ǎ`�!�sb��;r��D��x�~�����y!z��y�u��߭�e�����d-@U�b;~a�o�AX�^f;���o�xC�gH�L�8E�H�4��_\��[Ƙ�*,������0�,{sX^\yJ�~�]�#��%���ZF� +_#y}���u72��4�ɐ����,�+9�+jZ�������߻ooȎ#Ϳ���n��5�d#
��1����=�Y3��Y� ��#���z�!�p��T��_f}���]_�IG�����:���tm�D�.�q|P�c����.��v/sC��1�K��vj�:�:9;3n�;/���4�P��챽lm+{�ѓdG�:6	���Ơ�rqs�<�����1�em�dV�R|.��$W��j=���Y|-�څl��L����/I�`����6�ݏ^��q��Q�P�i��b�$Xj�]��|W��Gc��U|��zf��
VM��&F��� ��?��&�[Z]Wvp"�4�v�iZ)}ա7!ts5&�6��lic�y�\6ޜ��\ik�Tt��Q��:��1�iTEb��&M�[*3u�4�뗎�a�r���c,qݜ�Ɲ���<�feM\�ͺ<fN7[f���"�)���@ԉ]֝Cb��h�v�uo���w���@�@�?{��������$j0��[]���SU�[)����옢�mc��h#��/[5����p�x�p�{6�q����]���s�ZB6����I^0l�����Gs]�G���v��!�2�!v�y��k��%�z2E��s��inDwDך��U�E(EO#�4�L3�U��J�d#q���z`Ȭ�xs��\a�|r�W�rv�ElKG��]=v�b�l���IT�)B�.Gy!��pf����D�
���X0�ҏj��gN�I��ݻ(��_a��r������˦���U��jF��l�2n⻳���v5�W7�z]�vl���z�C�|����������j�=t.��E�3()R��1T�*"T��*�T��%-�b���([�Z�襈��T�QX���DR#hX��R�c��3VV"�����t�Qf�b��4V�F�����T۬�V.�QB*�,[�U�J�EXQ����r��TEq�(��*ԣ�\B�m2��!TKJ���D�1UF"�f�`��v�8ƈc����AV��"���1�6���i�*�����ǻ�k|4l��*u1$u���0�ʀf�.�.���HQ����/����6�]� S�#Ma��Lyb�oY�	���cY�����\pkm�=��=O��o8����%���(|�|����u�Uz�X������O��7�������{C�=�ݍ"� B��3��{*��^ڂ8a�����u>k%��!�ͤ���̺�z@��}9?!__!�l�za�*���Б 3|��A�������H�5zųF�<�{��Po!G�6Yys��XT\C
���}�u�y�H�i�,��ۨ@a�8�M�����2����;β{��Ӝ������c6W���׶�`��e� {�ݜ�J�a��gw<��sI�Y*.��-�g=\���U�ڞ���E^�;ϩ��rkS�ľ����W����?+Zp�L�&R���8��@Vo�ssҮ��/
Ao�~)6&����/���Owa<�����(Y��hj�o�V��F	����z��o�?���6|��������`��F�=:X��]lg���B!��g��E�]�y]��N�n/��oo��=�o����^��Zq�gN�zU�e�|v =��Z����G�e/�K�ȶ.Y<�U��h�+|��i�d}�/���t���)��#���<`�2s����Z�y|������[ҫL}�zh�ߔ����Y��wf�s��6yNrox�.��\�����Z����b���o�ߠ���"�{���۴��Ld�8�&k�Pko oI�'�\�/:YNT���w��,{������� ���߽U������֭�fa/���;�kF���k�����ge�9�۞����f�$8���9��!��営{6�� ���<w�W�1��8~��҈�e^�[ϊCO��/_�5邓?���i��F�����h��h�_F����������蹥�����G��� #�^b��õ�-��/}��v��#�v�W�x��0��e�[�������F
w��ꙷ��N�N��}������g�����?<�7V�v����ť�Ŧ���{o�pԫc__F#D�����[T���m)@�\�r({�Ѣ��h:��������_u�)�zX��ж�*A�����x������ۥ�W��W�(Q���(�]~T�۾��C%\����}���0���x����Q�t�~����꼏W����?_�]]��^�U���{�+����zB�)n���⻃Ob�?Q���VE�����U�w{7+�,�G�xԶ!�0���,8~dB+��WJd_>���ָѲ=HQȾ�lS��C�W�\^!k�#l-y~���a�p6Ǐ�Y����4�$�q�P]�wb��t�q|i>A�,s�� ����{�罸��>#|5��2�=H��q���ڕ�(Y��0�o��p�0��b5���$=�貤�6AzE�X �ZQ*g�#�������V!�&o���y��P&��+�6A�3�(������U}�Vy�O���Ӻ�
��k���1��/_��
�}��G�1L�z��L��laZW�^O�,�YC���z,��
��<��>^8��p�@+C
�s�׽[��Gb��	d1�/���������L�b�e��j�]�?n&E�T_����'�0y�{U�T�����,���>(������b������ӫ�-���w�]��<��"$�����r{��3������c�}�Ύ�U� :P۽^��B�2v�'����x񇏹}O�xY@k%��u>Q�E9y������#�!�ߘ�@w-?��W�jV�oB��h���w:�#z?g�|���kh>�S����������Z:�z)׃N듛���Ë6�T����V�E�#�HH{��}s�]?����n�uL;�_y�8��/�^Wv�l�8y�dq�a mY����s�;
����6d��P����"��|{N�����+����=��#Y\�wnJ><a'O�;k+K�7W��Hc�]񦻻ٱ��򥧌�˴M>?i���Uu���yo�~�ܝ���?py���{�9��w}¾�D�F�x�\��0=��y��y�r�v�x�^�5����U������Of:���#i?:hO}�>�/T�ą���x���t�}���g����"��0���n�#
 ��.�v�rw*����Ǯ[l�j�.��s7,p����	�FT�v�[�/f�狷�b�:ws�R��WN��ޝ��?C��{ՙZ~(~�Xn����T|x��g���l4�!E��AY���S���x�yڶ��Dq�R9�����<FI����+����Edf�#*��n��0�P0���HQA����5�����ʮ���܄���2��v��ol��_߭��1Bsݩ��2�-8Qk���ư��(Z��Ǚx�s��ldC���q���^\~�ZQh`�˾�w��^F�>?�0�1��8~Ʊ$���f�x�>���/�������i�����w�腖_{�W�0�?{���`�(��������-9��P恃1z%fx����2a�Έ2P݇YJS����돆��#�͹,����d��Q�8��v)�W�}_UWv�9���{gN��;�U;M�=�/�m�^1������2;�:E�1�a!b�,��m.�o��[�Hw�lJC��_sp���<OPkW��0r-�k�K(���;�i���Ay0�Z|t�v���ӗ�Y������Q�9���+��=x𱋈��W3�:�D_��B����B�>�GG{}�I|��U���}ዎ���	G`�|���؆�۞�]Uy�����CK?wy�<{1�@���ܨ�lQ�QL��u�����z��.�
��vF ��U�b�f���^h'ό��)
8~ڶ)��E�1�����Ȏ��m��Y���YQ�n�e��q�ԃkA=f�U�f|�."�ꚫ��2+�.�dU&��Y�:�ٔ\F�vm.�5�9��	���S�����fc�8������憐��&������7��>. ���@��X�Zvy�^��w������|0�ak�x��:�&�a������}����G��]�t�7y�F�gA�����>ݯ_w] �x�RC�J�a��SP��+;*�u�c��?=6Q#�di^XG������ו�����#Hm����n��&l�daGCyb��s�����?2"L�1}��z�h���}w�V�$M�F�ͫ�Xˮ�(щ>#O03�ܟ�R��4/�y�r����1����,���;�O���e��>ٽ瞸&�����F��ݩ��J��\<���
߽^��ǆ���*\m�x�	5[�gu�U�ݚ2�B��ɗ�e�_k�����U}㍧�[�_�K?,N�����՞CM�O���Eg�S*x�t8�P�h���+���a�u.��,; ֲOw�9��QV��`q~0�����,w�R�/�*#����㮧x��R�A��O��}o�m�5싵a��g�s>!Kś CP*:B��/�,�A]�W��ѧ�LZBC���gﻕ�s�k���Q�,�!D0���8Go��q��|$�z�ٝ�^_<�����������d�wf3�J��+
�2T����=f��H��f0<jC\� ��&3�J�Xt�& (�}��ε�׿u�^;a�1 �0+"ŗt�$�(T������*x�^u`c0�v���+&��0+G�_5�[���\��u��o�ߡ�Aa�e ����φJ��v�{a�_Sx¤d�R1�E��T�)��H,��<d�1�'��מ���]��=ޕ�0��1DEã��Z�^)�b�*l�/M{݂�6��wW9�b^�^R��d��wĶ��0^�]n���*	�����Z�^���D�6��_Yff�х��+xȗ��!����<�0�N�x:�E��Q��ckj+7�g���[��w^���1��i��(�9-��DBٗ����h���ǣ C*`A��Z��2�k�֧I$Y����][T�k�&+���&��?T���\��^�h�md���c# �+6jV<��;uQ�/e�^Tރ��jf�[:��D/�U�����Q�	�+G[��'0�������ojS�qs瀍:����¨)w�qA�+x��L�H�N�Ӣ�]�ےn��qi0U��mƮ�W��N�����ܨ��"+����f ً�b�mI&n��I�����!]���xE��]e-�؍�2��Ccz�D�$_4w��3�z�ι�V�ܼ��_Xϐ��}7m�Lc�����t)Ƒv�u�+�w2��CvV ��mQ����b����٪�e���8l��4��ʚ
%'ff��k�K�u�X �wg�u�Za-�Րν7���X53���{ί�q���P������j�p�e�P�"��S_sF��q����>�L�+�]�o]*��V�ɑ��P��@��0�c��f0��vS�溏K�#��y�����5)^uD'+/~s���=ED�W�0Q1���3,OmE"�\j
�Ҋ�V��EЗVW13*1AM�Mh�D���o+��C-Qe�kb	�
"��
 ��6�T]4b:�� �S-�F,���J2,Pıt�w�d6�EF
 �EUUQT�*(����&5J�Q����]�U1�"��M4b(����Z$EU�U�K6�4��0��W)UUCL�4D��Z��Q��AV�"��ATJ���hٽ�����������`�wd�\�R�b��9�~������/�����*�xöbT
��N�*Aa����
�_�L�Y��@���Y��'���
�e����g���y�_}}4���_~�g�6�P��&0��a�������5��A@QC��<@�lIY�JɌ�6³�Mu� ��y��)6˾����{�~Cl���}LH,>g��AH,�Ɉ
);�M0񘁾S"��P�$4'hbAI�Qa�;dѫ���L*?w�s��|��w�0�
��+��|yf (�05���9i�
�X9a�R
|�0<j��p�'��8�*AI�q1��V�.����s����6��T���LE�l��o��i �m��d�;C���
AN T�����d��1=@���z`V|�R�5�N`��}ם����� Q �����+>Փ
M{CX5;g�1 �`V0�m�$=g��I~j$��O:���.�޺�ߏ@�d�=��V|���!m:IQH)�L`x��$f��H)�읦�Y�J���bO���N����9u�u���¤�C
B���;a�bAa�|8�Xx¦���J�t�R�a ��)�n�R^w�y��η���}���P~�
t�� ��>La�
��*%`x}qE�����RbAH,�%a�m��R��
�o�y�y�mw��{�|N�+�l1>@�%a��{�Ă����H��}CBA@�T�-�W��
NШ
);f�c����\�Q��>��4�Ƥk�G_kT�n�	G%��J�	��\r��U�TO\�c���#��GF��I�/e�����{?_}���{��H,+
���q��
��I�E�(m%N o)��T���g��1 �~%ORTR���0<k7�&$n�5�����y�� �J���R������bAd�Y�a�
��Rx�H)�iXx§�׶H,4���$a����
��Ǯ�������였���bv�R�AH,+e �ᒰ8ԝ%E �dּͤ����cT;�4��b����y�v�xz������'H��=���钰�e�$N2�5i�N�+4�Sh�0�:a]�h��H)�,��ALv{dАRu��y�k^o�w�����q\H)��v�@QC9I��=a����H,8��0�*AM�bA@QCI*q�x��R���_p����{����:H)=��'�*(J�@���R
?3��AH��v�~jALa�18�R
��a��Ri
��}��������<��Xc
�{�i �����Aa�t��_���!�
/^Y4�@�>C̤%a�<�Ay-��8�3��AO�z�p���]}�ӷԂ�P1+XT�
��P�%@Qd�^d�|�J���=d��t��T����0S�
�@��*x�Y�{��yַ�o��I��W�AH(J��QH)�
$�C�ç�P�A`f�$�
���:�bvϘc�a����c0���:��;�g_}����|IR=>��P�%N���H,�%H,:a]�l��Y��<IQIP��
�}� �~��>M�:IP;J��O�s�o�j�x��]y�u}��#��`��ŀ�A3���Wt��λrZ�Jt-��>E�wv��:��	9�o��%H)�����AH)��c��5;�Ğ!Y4~Y��T��lLa��z,1 ��g��AH.��1;@��:���{�^}�^�'Ǵ1��s,���X��V$�5����&��=JÈo�IISH �tʛE%d�*Ag̖Boϻ���_o�� x��ô�hI<`S�IěgI!��$�ΐ�����s�:����:�߾���
�R
i�a�� �ά1�l*�P�%H;�*IS��)�3�1 ��&3�J�]0*x�P�_3��+��k��=&�*OY� ��&$�@�*�&$��1 �7�d�aSh'�V������� ����{����s��醒=N�bA|a��$��*v�R����V���
�X�Ă�S���
IP<JÉ�����^���p�s���\~��P8�e �(m�<E%a�
�Y����x¤C���@��H)�&��H,+
�v$5����z��}���v�Y>��J�Fr�AHwi������T�!Y:eH)�<a�� ��a��l*IR
ACI+׽_.v��Z��{��=>�I���r���%`k��<@��`bT
�L<q �|���z���
�Q@R
VhN٤�ɇ��޹�]����"Ň�*AI�+=ݓwa��@���L*Au�a���<dĂ���c��2z�C��S�
�s(u�iϵ������wͧ�<B�5n?f�S����6�4�oӲ��ذU��ыNS��yTt&�S\R
%M�D�O������=�����$O��qE!����q ��*IX?� �kZ�I
������	VP�g���>����%>���ey�,�0��#��l���t��y{_�����~��8gظ�_W�"Z
�F���佬��˼��`/�z?O!���i��E��G4�����64�9�z��o�Gw�Լ�P�>��Ft]Ə�)�^=&3�g;��sۧ��m�t�6G���g(~��\�!��q~_S�F����7��7�E����B�H�������}|�ދ�nK�F{E\E��}����?�G�X����Di�CRFVG���lq�<j�T�46������5:ptu�Ka'$�2��Mk�1E�|��ui��6{�3�9�����/K�	P�/{�]�?�����29�]~��?^�z�n��+�K,S����ǁ����}#���GM�H�#�o�ei�7W�o��o��}��9���:hRe�D����>�M���gw����)�a�A�>Z~$SCNCǠ�3�����G��_^"a��b��1Ն��Ҝr�;�~�@L�;��6���i�a�O�b5�t,܅��!��Q"��"�$
�őڍ-��ύl�/��g���b����B�;9��nl��D	g�1�i����ő�����Ҥ2���~�P��c���צ�a���E����k܇D��4�;�����S��;ᚶwMІ�A7�2���ܒgc�,bI�:���~�����W�.�I3�������bi����ȣ�h�g����ϥ���?)���^s�u�ϸ��cH�A�2�
)��b�-��o�\�#di�d=X}��W�����l�4�'�S�)����=j��C�]��;w��A�]���<W���"�y���\c���CǏ���o�s4`��� Pyг�H���~a�c�fO?UVf�,����=/�F��Z���0��U��f��`"Μw���F�0�2<_.y���ۋ�8s�ꟾ��rm_�G�C�Ԗʞ�h���c��P�y�b����F�+�ԯu�q�*�%UWR{Z4j��Њ�R�ʒ�(��5-�H�q��aۀ��.�����U��y�9�?>|>�I�����L1�7K�|�c�Xx���^�/۳���/����э2��O����B��Y�ʮ;W��]:~�l���Ƽ����)_���k��b^�+�u�(�ٔ��F�/��q�vz}�=�I3���_>�>�,�����	GN`_��6]߷&���=�!\�����?tx����(]�yu�����JCǏ�<t�C"�+?1��u{1z���ƈ�"��Ť1HQȾ�B�>?)�=�1����!a�����͆>ʂ�;Z%���5lG�������e��:�B��C���2�zSg�v6����赃o�u��j �e.�ر�Hd�&\� m�w0��eT��&����u���������iO�u�
U~�_U��S��>F�!�@���:��onX��$Y}\�Z~����0�ӐԹ~_#������C�J�cǹit�lm?w�{޲<�!�|�a������4�+#��2n̫��{�+@t_q��4��Ӏ�!����ON�V��HeD*��G�G�dx��#�Ƶċ�����{xz|�3W���Ȗ�$�>#!B��}��x�jz�Z\�&/��X���A4�f��g臭9< VG�}Gqx�=��y�l4s���e��QC�_�^<*J(7�E/T.���h�Y�$p��hh�޽�8)�wT��/����x�:_9�$uύ۝y�m,o4#��Ó�&K{������jJx����6��:�}�^=�}z=�xu�|^s��f����Y�C�!�m���y
k�k�����`��oL"���l�D4¢�<��G�he��g�_�s"υ�HLCN�՟�?x�������#b,*0��CH!����a~_k�~(b�%�X4�!�@)�0yx�H��:��Ei�7W����5�|S��r�����^<vץt��@mz(�ո��>�\t������'�OĈpS����f,�1���&"�0�^H��毝�W^˽ž f %����6�0-,;U �'j�n�9-cr��)>�kx�;t��XL�Q�_�Y��fY�㣠:�=�|��M
����ε�Y�z�v��! ך�}����������w��y������v��x;�4c��<ZAE�>?v}��"��ŧ��Mmʝo�M���$(�y0��t����C��n�Z�n�|��_B�(����!G�bM��d^�]71����\~��Q���3�c�z|忌��dQ痝�^^��#|��s�"4�l��(�9U^m9����#H�,#'=:Q��`Ak�Ka��Uw�q����.,R�e�o���8|G	���ל����L�*�5�~�"���O?}�%��c��d���*�4:e��4e:p��1�y�/��s]i��^a���*;��װ�&�.��e�if:�����.�r3�>���W�-�y��-wd�皅`�f&-��B�ATҜb�~�x���կA�m��s��B�^��3�:��� ��5+_�b�˶�'l&ݑ�ջ0w��qKᶻ���Te����4RR�p�jݼ��w���Öc6�h�vM��H�3�.ރ�[Qg7Ϲ՝���Ud��u]k����	��Q\]N�K����YܻRi�zڻU�yHq�9���6��J�4-�h�$D�����y����M�u#o[���CVEI�6�҂����o�8-̓���r)l�:'߸�gcyۣ�^ԙkq/V��>=��P��,Ɯ�w�����ʳ�W�;�z����JX����x,�/���
��uJ��e��1�Q��[�)Ͼ�*��M�I�V���&�m�ݭ���*J��D_[q�9w#[,V_S�Ee'say�zۻ��R[!$_T'y��m���F���{�e�"=�j�b�ݧ_��z�.��fɜ�}��p/s�s8��{ܙ��Χ/���:r�S's��V���a5��>�*������-��B��	;�ڕ�����D���d��2�X8
	�Rf�4 ׳����*v,���O����Іv�a�%a��}��pl�.�p��n噔3ryg�8���q�}.�Iݐ�vs��\긄�9���ԝ�U��_���j��nv�1����5��FcV#KE�`�`�)t�d*4�IX�UGWyL[b�ժ�"���fR����imE �,\kv���]������%U����q����U�\�s(i̪�.�Qwh��Q�U�EU�"*8�-��h���Uc]��b"*����X�i\���`��B��owH���v�E���\�QL�٤˧�ZWXU`��GZ�"��J��DO����M��3�7]��UY��UY��9Ti֋зJ�5y~� y�o}w���LI�:���;�՞:ݍ3g�ե��V"+B^��{�����5ic��lхF?���y��}Y�]o˗��_x���r�3Q"��C8=���o.�^��(�y�<EE�9{�B0��MA��Jk}Ya�^!��%����ڗ��V�h}yXt'Њi)�}ޞ�X��i�?-X��ڷ������ݧ�^ѳr���jꕋ6Ϸ<p���y��@�[���r6�ỻ�'����x�w1���������|�l��+�_��~�;��&o�T����غ�Fi��b���r�]�i2��� ��P�5ɬ�!^]Z��X�IS���5!\����r���sv�y�������$�t,����r-���g������ ����}�-v��+L��-N��3Ϯ�<8�A.�/w�7�����>��X�4\�1�d��� lJ�֍���浖V2��#O3�����)�i+��2�������9Ց]�]ϋ ��!p����&��5J�U��9��^P��,ɄxDk��[� ���.&C�Z���؛/��� ں�'O���p��&��9y�۹�)�S�movNS'X�cWp����9���~V�����9;{�3��}U��p��˚��N]�en������]Ė�._4��̦O2�X�_Y�W�Y��,�=��%��v�J���{�Ou`w�Sk�LͅJ� �[�o\�dj���;�I�T�2Z@���6��7"��q�a��t�p��so|��uo��چqޮ����=e�]�ea�4l�磔�[���s��ǤVͼ��(!:�VVR�Ƶu�~�sN��/=Y{�ƕ�ǩ��R�k��t���G�G�ݱ]-���u�|,&��N������ �=P�h�������C$��ZCᙍd��&>_{]����Y�B�ǂ�_���HR&�yOn�J�V}N��|�}(e+��g�c��燵;�&���Q)y�Ә^�?A�&|���lf�Q>�}���"�>��eḽ�+(0B��}�T}�}�=ݫ&�(Ᏼ��]�}�R�����d��.G}��~s���'s��'t�ۅ��G@n�Ό�5���L��AYװU����}��}~xM�b^�o�Q��٥�7n��i�e���x�l)�ˏ;���fY�y�d�W��>o���U�}_dŤ�����ɣmb2i����K׾�\d�;ai�6m�:��7s���Z��<A93W�3��/Ȏ�3�9���z�@,΋�c��Й��^��1��)8r�vk��=��+6�gz��o�*���>�s5z6���{�����5��vF�y��jϕ�!�Zr��O��2��+���E����W0�}"��eZ5rf�w���^�v9Ջfv�[��uN8n��<#�T�>8��>.��� �L|tdӼ�m䗁��k4�HKs����s���}_W�:K���%��w'�h�׭�C��D(��V�'8"X��F%��9��Gy]qI�,�;�,>��q�.흯��Ʒ�L�p��esԲ��k��,=hӝz:�|��ƴ[� �&=i�x��2�e&�2�]נx{�C�]�5zb�w��hO2�ŝf����`iJ������8��̓�iP����4���Nb�l��̆_�!K��e�W.��k��Ue2�r�T@����2���h�p.�<Ρf�&�T�w�"s�(Vv��C��U_W�X�4�߲�a���	�ZkTl�avFe^�pr��{�վ%���p�G�QŸEX���ŝV���w�~RQ��b�B�0����'N,�μ=�����v[�ُ*Xvhh����֎a�E̖�׽z�{����Y�#^唤��v��$�9��WdN�zn.`�P�Y��%�L�������c�n�=�^��-���lg��s�&B�nx�R�v[�.�}�/L�Ջō�t��FTڄe~��՛��@�➤�3|��+��Ɏ�e*	�W�{��{���w�}UU��֟e��G�}��[G���.O�9^��n�r��IV_��oN�RJu+[6��z$L`n]9��ݦ�r����42�y���9��9��c=8]���ϭ�
p��Fyu����aQ��������5�	4q����w���z�^1
lj��K���Y��m���!#�"���:�
V���:�,�'9�W��}�.I�&�7;i(�P^5�+��pd���z�B6s]��	� ���C}������*��ݣ�N���6C������͑�9�?K��u߻ �����̯w���	�;�(zw��tE#�Au�6t-����+���}6�WXP�;i�yr�h���_���~�~K�W�d��� ����)�m���l�c{�z�U���㷚��9`^˅tuf?t��>�G���x����a���G�y�-�¹�����vz6��]Pq�!\M�o�w��GV\��k)v�� jk��Q�={ا�<���j�-���!vy��"�=�T�����ߍ`�<��8�70������(�fڜ4���5�U�� >����5��_�f�=f_��ܣPyH@�"7����w94}������U�M6Vu�I|��nT�)w&��1��mY�`N�F�E���%
�/F���<vk�?i^úg*Gm�enl9u��u��sq&��ob��໦��M���z�'\����`��k�O�������uw���Ϗ,�N�?g��O<s�+��C���{ϱ�XtϪ%�`ŻŷZ��p[���,��$Ci��3v� L�s�r�������m�Z�K�NIÞ
M����p�o\nZFV6x^�9W��㻨h��4���$� a�=7p�����$R�3`]�2]��=��嶓���fuM��&��7�n�ap�����38���b���D�yGI+;&�KN䐹�Y�5_T��n1w�ڣ��9X��p����ۣ��S�\[���r�����A�ݓ��v��Q7�֮�'�hѠ¬]��&guῙ�ۉV��֏LY�C{7rE�1G�GOr����|ۜn�Ҕ�����z�l�Y�Q�YY.qk�\�X�71@��?PWy������ǐ����[�"����y)q΋]>�J�<�R�.gb�'{�dpv�آhr�����(`0�]����v�֡��c'��d}�&�}A�zл��y�,��Z������Z�Gp��)eL���PɄl�+�]�4�«�oy*y�g�7�X��o~�G^�F�GRU,ob�󫂅:��OvƎ"~;�[�3EmՊ���J�[���TS�d��u�!���2QLz$Ï*o0VH;�c����êt��䬑��2!j�׽K�)�μxcq�}�s+GI�7����Ф���O%I=�|	�/���̓�|sx��$�.g^C\rrV�Wں�U�s�!]{�7C�������a�y�Q �_D(�I$�����l�l��b:��%TXŊ���oZ1UB��Y���fE2��nUw�޲Mj�Z$DDQ[X���m2��*�,ESMb�A���faDk6�4U7J�A���.AKD�Ks)�]Z#R�Ъ�DSkf\�UX�]`f�TQb�5���-���m�k\B��(Ա�ʘʊ�����7�GR�k3v���Q�*�.���m�jff��E���U4�[��Щ[5��ETjT1iU�3(+(�eK�3!Mډ�
�iE��c�6�����J�U�jQ�5n�{�]u�y�U�]���z�r���M��ni��s�M�i�ﾪ�}�����RY�G1�,�{w -���Ν�(�s|��K�Gj�i��9�s6�Ʈ4�130�r<u�mb�7�PkW}��B���Ӽ���m�ny�i�j�+��5^��&_֏x�CP��FlB4�{T����s��ݦxN؈T�
Ʊ\�R�ءY����a.��3L1��ὺ>�����S�/X�Z^�ݝ�9�~�J�d[H\�_�Ys��o���	Uy�ሿr�ZK,��4Cҥ1\�
���#�7tˮ�;�"�������tr�%���U}{��_��g�o���P_bY�)Ն{��b: q�p�^U�{�,-I`�(��z�Sz�{�;2w^!v��VC�6�x�l^�.��<it:=ȝ$>g2��J��A�^a��9%B���F�~���X=0ySJ�9-��Er��}�/�,����f'=��k+8���^�Ev��5�NW�A����������Zھ
���Wcv�̀r�X�����I���\�e>Av��ȷ�A(��+p��]�ǀB2��iNe���$K=}�����M8��`CK��xS �5�]c_�y�g��2b;�^ڈ|�٦{|����s,)�v�bmT���&jh�ku�X��>�wU�����l�2M������'�-�Wuj,�\��줢��E��4(�[��ywP�iA���N��w=�kyJx��ux��m���q,^:�Ѩ�r��y/�"���~�!��r���T�o����^���;Y=��<<㠣�T� o;��JVO������,�N���Ų��=$ё�i��s5g�j���/��l)y0W���}�}�ķ���>������pËq��u2t<�/4��1{��_y�����Z�|�fpts��x�&��v�v�͌�=�� 4�V4�z�_�x����3���/!x�<k����^���l�;Q��s99xV�Ƈy�U���w&sNo��[��6|�ѳ�M�G�/:�7x�1�䲕��(E��=�:��=]9H��n�\'�}^����t"�W���:�����op7H7械�ؖp*�_m:�`bR�/�3� "�t]
�B���qٛvx������~����*j����vi�~�p�Zz������;�7����I��~W�5J�<��]}�B$X�{�y!jx^Oy�r}[B{��G�-����T�A�=�D3�؍/r�{{nznE��<d$�uh&ҏ�C���{ث����]II��};������f��u쨴��\G�N�[JD~�*z����N���cF�M��E��l>�rqU��_8�,ߧ=~��=����e�2j�8S�S����e�54��kw&l���l�=W����"E�qś���MU�H���9�fp�k���S�š���9�
z%ֵ�}�w��X\XA�f�q�]G������?�S^����ݺy�=�n5Ψ�M�p�p�wbӻ��~�7�+�H�^��9�������뤆��)� M������{�����ѵ�)��K���ζ�O��u�b��Т�t�������>�J8�j�(���_!z�A^)W� ZqYd>S��*~0{tp�+>�e�VF��ՙ\6��wBV�ߍc�YP���K��&E�W��ՙ}S�b2��
W��ϱ�H{�u���V~�M������r�u`%����Mb'�ɴ���s��/���һ��ƹ��?4��q��_�^J�l/0�G:��k��h�ߠ�٧�/�^�zk���8�u�ܽQk78��T�fE��ge�Xp�c�2��QMe�s���Y{x'^8+L��j��z�\��;���ІN;��C�n-�H�)��Imz�vAs���Vu��)��J0rۇs�z���<��H�Y"�^!v;�/r33���e,!�m��g?���W���	�0O����ګu�39ccy�;�$���b�0ˮB���;M��[�-�vf��n�ܶ�k8D#=,����ݚ�U��^�!yi�}mw��.\M\z��4i���V���^-�w#�mZ�wf8D5g��A=1��1��u|��dRJvj�)˦��8�h�y��G�b��K�x��h�AǎFp��	3��ѹ�ٰQ���UU+��toչRw�,�U{��=��b��Eѡ�'n�ۙ�ҝٔS���2�����[I؜��s.F��u�����/j�'Fl�DI|�%���[�����V��}dVu�G�}0�zg?C.w��;XE >}������9u!��Z���=��Ճu7�I}��j�s�	���R���"��+P՞^ғ�8���.�ں{��U���g��{��ἥ�~���VV�=�g]pS����_/B#�<�緟I�U;Ջ�����'d�'�ۤ�g��۟F-�W`� ʏ�=Ic��s���=j;*���W=�;ۄfʥ��X�G��dOj�?L��]=|�;�e#�Df��S����]�Q�
�gl��]s�4���F�=V���2���*�CU����iJ�����)Bd���֬#õY��)�;>�/�a�^����P�Ֆzt���$J;(�`�t�%�sK!g��\"kQ�G�{�n7��&nxg*��"��F��{!3K��7�_|c�Z�^�l�,�OnV��Eb]�>��S�i�@���*�j�W^��t�h��F��2Q��M���������9?��S�[�m���>�i�)`�֥n����q��
�qx��̇2_A*<ko��`GZg|һϻ�0:5x�et\U���q>�z����:�Z�o�
�ѡ����ċ;gMr�ib�^�9^�,�8W.H�ǆ-p�tR�0k�7/6v^���NM�\�5J(d�%�{y�Jֺ�W��i;�5֋CÛ�5���Vv�ȝF�x�C��ʆ%E��WOz��fs}f7۶v&��w	�F���]7M�͉����=�P������=r`7�8��n�i�d���/�[:^t!�S���L���5�T��}�F��@�*ѲNF��?��ꡂ�_.&�K��j��v'P�6Ce�*��������\/�4o1QI�j���t�H���9Q+{Yi꼗�����뢹��O��j]�fm��:�Ω:	�W:��CK'?ø�y<4PU�j������b��Q�GWIǨ����&�<����wEr:F��f�`̖�)G���or�a��Ef
�	�*f�9�n�Q=%J@�-���Ywv��]���j�"jG��\fep��t����6�I3��Z*r��6�b�z���5�IgjZ�qNo��U�q̝��]Ռ[E�=�{����8��[��O
�ٚ��h�S6*ee:(�����zk6����V��w����J�uO^���u�z�a��۩X����f��r�v�Q�.o*�yv�S��َ7��6�fM��z��U���I��CYm���4t��J�B��"�e���i��Dm)1m�\L�5mQ:ji.��e&e�[7��W�i���:\�uK[2�T���VkZŘ��U�SIL�M�d��k���.�4E.���Z�ZV�P�iuk5m-f�fe���hT�n�Dq�J�����L�Y��
#Q�3,�aR�Qj�S)L�0¹��8���-�iYk�T-c��jŬ�Z%@̙�AD.�pCE��K��1��[���(��-6�:j���ZԴ��V��KQTZ��b�r�0R�\�0�"��c��(bQ�b�����%��=?�%u��7��p����(̅_8�}�
��⯳�R|Ícy���n�pS��&�W�x�����6��&��X��to����~��(vƷu��0+�������j��T�D(��������c���{{aN(U�oxĻ����jq!���S̕M7��}�0�(�U#��kJ�4Cu}���je��8�]���ӝ����A�J~��{���77�x���Z>�o�ׅ缞X��[�
������[g�xfY��Y�-�(�KL��)�nk���U�`j8j��6̫+7�����|=���~%`glE�_�_�涉��g�g{��"�+��'e\�L��%_�^�^%S��+d�[�E�ޔ��bh>� h���B7<�Tx�xȖ�Xv.م�!7���m{��F�y킪Ƚ묹t�;*F��݇d��R~���p������<2ݞ��D��MgٻhS�paܼ�{�|�[��U��f�v
~f�v�f&U�x�m
��ѲϹQ��ߊu��G��IȲY��1f��S8٢�Uϳڮd�'G�p޾���y\ɾ�ڡv�݃ /�^A�O6���g��&-�ߦ7Q�Nx�&�`�xz��t��>d[XCU
���ovw�y�[c���v1z�'��z�U�Y��8�~���{ˇ6��Ly��=�Yb(f��n^
m+�(|��jϪ��7.�o�d�����7�*Z�)���1�\�"Q�d����䞞�Vd�~���%�L����u�ڛ�s �J�NK���mκ�������w��xOO��:�MηV�g�fuc;X%a$��Ӫ��=�ͺ���t:���G��ɚ�T��,5�Y��'�A�ʚw�ﻱ4�ly~��['hW~Y�_��]�'�g�����z�35�J
��%��ra�&�nѸ�Y|���A�K���;�o�O^R��fY�N� �J!�S$��ŋ���v��،�:���U�f�7�@SV�7�Oj���z_��6�Du�z�*X�.(����dr���յ��ue�gkpXܮ��-�PZ���B��9栱wX�^��Np"�.�ѯ+b:𾶸�;H��3+Y��j������ڱ.�D,��S����L+n��=/�ǖ��+�i׸�����}��,���X*��G��bӁ�(��˳3x��8�L�{�X����z��t���ݡ^�\����~Az�+��w�.��^�kޙb���M3C`�{P��qG2�����_��I�&�7�ޅ<��WQ滳�Lh�T�'�k�#Y�u���:��n��ɫ����ݰM3���#ո���!�q�	x-�w_N�Om6=$�c��;�C��:o�։�{����6�:��m�i��jBs]�_m�Lv�烷�����h]�Y�˧J�H�8�q!<��w��׭>C��4{�"���v3/�)��=";����D@8y����\q���:_Wp�S�/C1\5@�ew�F��"�ۏ��U��efz,�����6���ْ2pn�4"��n��ڠS�V�4A­u�+bH�=��.V_�'&R�p�k�;Db�m�7 �zgj?�u�<�gy�C�3J�獪!�=x�N̕o�έ���B_�������o)�¯ܮ�n�����&r*1eں���k,=�IVi�R%ه;��=��J9��w+o�nB���
��_����~�-9讻|���1��E�Y�+}>Ϝ/7#����5�L�5]�������ӱSɌQ���g܏���ja� :�D~�I|�~�]�ƢK��s�ǝ�<��
Y�4��z}I}���r��PD\�G]�Y��V����?o���Wa�je���e�;�g9�Q�~ˢ�<D�3[������fń+E�}��U-.�W��o�7���+-fm*e0�u�pod]��b%]�7��@@Z�����ܕ������=s�VU�7������V~u��+�fӟжnۖ�="�n�=���s�+v��7��̉9e�5�b�C/�:�V��ðe�3;;+\���~;��y��N�?�{�r��˭�}|+�{�v��硙���R��)��]�h>�]�Z�:Kzna6�hnя�{M�*c}M�d�0�ׯ�*��{���]q镳��;F{:߽{e�ԓL��U���;�����~/f�gc��ed5�b� %�♚3a�c��Y(S�D(k�^*Lv]�ggN���/��l���x��:x����x��4����4�~0�4������u�EZ��~̻�m��q%Z�F��wz�����-ޖN:|l�v�iC*P���yi�v��C]Z��9\�|�aX��cS��.��s4������`�ӵ���Y�Ӯzd�K� ��l#W�K{��b���ن{�b2x�=��E���`��V���
AX�2�M+{��r+�S'CR�2\�9��#�	������ޞ��Քq�p�2��\���q��K���:iY�%.��W�$W:��\Ғ��to/��R-���=�k�Wמ��۾�4���ތh�a~Ye�wosxQ�uVa��7��;LG61���Np�W�&�qהּٝ'_��vH�,�"uZk)����kr��+�ά�~7������J�ӏ_S��Y�zGO�2�ĵ��3�7�\���N^5��G�2V�i��ˈ�NCͽ�T�o��x����y�>�Q�owީ����'��?z��!dS�Ku]�,�7/j��Gܙp�t�:�=�e����n��{�y�&q�ӌ.��%�ۭc������ƅ�]��Ϸ&XL��9wp6"���;�6/ ��*��]-3�y�3q��kZp�F��.�B� B��|f�#�D'>a}��v,8�.���;V�������R��Հ���L��fi27����33�wѽ+��s^wd�0 C��ƫهb�;�u�$OM��.�j�ѶEt64��]\Ɠ����4\R�)o�^��W4.�}w���0��s�5��L�]�3�����7ZT�a��*�8(�ͫ����MZ���t�|�W9Aʪ���cJf%�]I��N���j��g1�SҞT�@me�
#���f'9����:��n��uk{���k�����d	�r�G�e�d���Js���wa�]ݓ�	\&Y�'s�z]J�Ⴓ9�����]O>V��[ݗS{�m�;N�D�3\�q�wX�oZ���s��Ư�d�V��Oq�t�]�	��r�Uӣg�B�s��\���`1;)}���}[�UӎuM;�����Ҏ�R�~�i8�8�}:xּ>N�n��6�n������f5ች���qF��K��Ư+����*�<�iC)crG�P�G�7�T����uƊ�Y|��FΫ�Q'����[Ю�[����s�u]�u.���0��$�5ζ�MAy5ut�;�cj��Lj`ђ���Z)D)�T�+A����X勘�.X\m�\�X�fUTKnP�6&�rfYm�aufe&8�Z�)iU)i2���%���nKnfn�tԩDY��U�1ʸ�T-3�i�ڵQ��1k[�䶘��ƅ�*Ze�L�ډQ�m�K��%k�D�ĭ�2��r�*.X��eef+piL�3iS4fU���-�c��Y\�F�D]�SV�R��R��1��*�)�F����ƶ�)L+�Z��f.aL0�-�m�0pm�0Un5qi�b6��of�AQG�e�;G�"��2���˕цK޾�ٿ�}��ӌw��Dެ�V�J�����g��TŞ��坢�尝�=[���jJG������]��f��j[d����ݜ$��gVr�����g�vt������ӄ-L�c�wx����ͽ^�os̳�pG�R���c��_\^�>"��~�Woh��x��z7tZ��0��z�z���ﲢ��<O�{��wOG>���X�e>9�:���x[lj�东&m���ں���jj���=��.�\�^z�����8
*�9��n���ރ���	���tua��}�K��S>��٣$g��#���Mx���	L���~��6V�� �y�$�k�G�rZl2���/������!D$uZ*�D���{����+�5����
�b�Ý^��j��{LU��]�˕��_	O����U�f�vp��f���qo#�6��N������p�w�b6��)���ܨ���u�3���u�)������uFhTU��s�w�	
����μ={�.�{�t��أ&��5���y�F�cf�Ԧ����.�aw	�{�NUS.w�z,Vs�܋��F�d�=6q?q�X��ښ�! ���In�2�a��g�E?|!���lz�QNa����fQ�z��h��u[	��˝Q��WJ������=%%�a+��L�������W�֞;��f<����\<]yX�k��l�X��w� ��"LI�4��֡�j���7�>�.�5��5�t���u��*4-�hט�`�0��'����(
�;����Y�V��ܨ��A�"~��lmA�ܲ�#PrY�J�����	|.vwZ����ꮛ�����Z�'>��՟,�"���1�yn>{k���)=	�C�7���u�|��/�Wv��9s�~b̾w�AQo]G�jKy��s�2�����Ӵ�W�D��iҝ���;#�t��y����5�
s1����tj���˫�\���|u�T;�d�5��*�"VU�)k&��!�Q�j�QJ竌귆����ag�-�:�ču��.�Vr��-S�"����*�N-;�{R�H�D���Fk���Δ�[8\�;5J���Z���@Eޣ��i%=��W�V�"�����^���T����OZ�܌ta��7u��vz�ܮ���s�O��cP���Av#I:�����Hڀ���u���{��awNd�����Eg4�3V�ڝm�����!_h�}�n<�TǱ��~�Z�p�[7��{�8�jI{��7p^�	�M:@*�sӡ��.��Cg�/!q4�xQF���hFOf���q��~�b�=�^x�;u>���*������ʴ��sx<��*f�r��h��c�1B��4����lb��.J�Ct�lo<��W��K�x���?;�:X�^w�X���W�����ҭ�X�#����,��ٓR�(+�eG��K�{Y�u�S���y��zM�u9��$ޏ�^���k��{/nX$];}��\�;�c\iWqzb�����5��/�tw�>���vV�^8�.p)��k8���V��k*۾[Ϣ�B�ٖ�w�+�d�.]�Z ��e{����2�v����d=n���.W\�S���@>o;��l�bΤ3�X�6c�N�Yٲu��d=�����i�g���� �4L�^��W�}��.O�{۩=�����\������~��w܊Q}4���
��߬��#������X��jsV���ȯ=4�{lx�WY5p��$�'q�՚ �a�ֻc�^f�+�\���2��^Nޟ��c<1��6�0s�Pl�A�<�IەOG���򶅇�o��}�O.+Р{�iԞL!s�<K��7�S_���wnh5�iڵ�{)���[˜�h��n�o,䔋���*;�f�
T��nG:gq
]� gi/�h٫�v�%�v�������S���n�_����J��n�#&��$�ͼ��\G�X�+N��Ƥ�sm	����}dX�t��T�bƘ���d������{設�Ԍ�{���[�d��#�	�G��C���x|G�����U������:��]�V�9/%W�eEa�6�ټb-�#Oy���;�����\��͂z��h�����U�������a���fJ>����k�rv�n�뗸Md�_3W
]������+N�)uV91Dq`������-�6tղ�/J�d��9����O���?,�,�������~�7Ǯ�n�
����Ѣ$O4���ZSr��5�q�t$�YSַ�"��,�/����+��F�
��ai����	����Gܯ�k\��1ٿf�U�X��7�s%Z��=�a�>u��^Z��=����o�Q�)�!�X�{�綱k^!�J{źk&�s�Cf挩�z5lد<����r�rŬ��m��z��6�̖��W�,��79��W�Yʹ�ecEU���Z1��;G\����6�@7y�uu�vu&�L����{�71������yr>�ؠ�nl>��իp��72��E�������⩾�\���^�n}{����"Jj�jn#�������zM-�F�Ȼ�ު���$@Y��T��*)���߿/GY��u�+�1O_��ﳷ�z�w�נN6ǔ�cP�u� ]�.g��v����v�}&U�|~��j�5��m!��bv�Q%Y��=EW���U_������o$��.5}5�,Z��V�t�36��ҽ�L �v��pv,�ǂ�s���Egl�ص\��u�D���T�t[�t/S��ж^�K@���!y�&j�oo$?:�_:淎 oz��3�p���TB���L�mK��z1�o�K�&�@J��f��4�9�������<5š�qk�,�#k'f�ζ �]�� ���o��Ko[Kv���i��j8��x�l�{��8f�nS2�qnNi�ɉ�[�#H����/d�M�ɵ�u:ɀ���)���o2kxM\C���=�j[�G^�殆e_�˦syS���]A�c;L�W`[�;6��'ͩ����VY��\�T2���W�=Xn��IZ�Z�aȯ^kӎjS���ύ�Ҩ���SXus�|]��ѝ�T�[�w.�7g�gw c��v�g��V��,Ż�X3�+�>P[vD��B�㳹�&�Y7(R���zx���ݒ�U�q������OiU��9��q���4:��؉�j󮮉���i1N�Aot�[��jyT��0t�oN�S������ v��|��ߌr��R\z��ݩ'%|�J��ݙ#�+��V���Hkq�]��BT�h�,7z�B�2�f���e�o6d��t��1�C[Pob3�peT�F:�6�]���oPk���:'a<�W�Wu�D��3����^���{��΂rG} �񩫫�y9'�y�.��0�G�LD�nfjV�oB�ڻ�m�q\���R�(���
܉����*�lk1(+KP����k��KJe�+D��&Vĭ̱r��T���*w�b���tD)s��h�4�KT�
S��ҭkV��ҥr�*��9R�Ke�ѷ331�Եn�r5���B�*X�j�Xf.e�V�m���eJ��Qj&���yqi�y~`���6��V�0��NWH��V����Jo���a�ܘG�KUX,�u�Ub��N� B���r��LO6���ͬ�p�[���pj�-k���暾���m#�nk7/��������Nw5�H����a�N�L�&9-��j�Rg�T�S��RT�k�����q.�O���;�wG���[�/G�N�N<�= ��L�zi#9�Xgǁ� �y02����ͣiK�YT�w�����K&M|��um����	��)��(��h����([<:�:��N=���ss#ݚK�Ց�*��'���Ԡ�/9�Op����*�Y�y�鎷K���>����u��g�Ig��굺����f�ה�د��S����������C�z�e��)ʸy��n/w1�vm�}�f�����¬���F�����u�//.#�e���{Ky9���	�&5b�^P]�	���o�~-HM����yG0���xN�9"2�M���K��Z�18�e�����z�>��^�� �_�o�o��i:�ڵ�{1Lj�ُ�k���+;��TY����[������%�HP�����Z�¾�"���a���I�v���	��;�.�	�e�@*��;��9{��ɷ��.\]i��{Q�=ӳ�%��������DnFli�7�����������q��d|��\6SKǦ�<�mbX�U���<�]�%qKݦ�n58{j7tZ�K}zw�V1�+��QO-j������S���]����
io������7����p�d�H_^r|t�ٶ�RA!�k���8�� �����S��؅`o]a�gx$ĸj's�zI�KՒ��W7�fT�a�޵n�y�d2�#l�ݪ�ϺLFo_7A�EF'c���K~�ܣ��z�^���FD�ft�ʋZ�w�x��� �f�t���Z�+����v:��h�Ň������׏Yu�qN��!���k7_n�����η�n�4"��[&�3�h����|7��&��O��~n\w�C\��K3s�np��m���0��b�iʴ9uԻGj5ּ"�m��/Ҟ
��gV	�龮;~]�e�NPg��C2� ��Xtp�/�ݯ^�h�#W��W�Í<�RŹ���N�	�)�1�ס�r�e�O�vڳ��#~�e:�����e=J�#�J�źH*kg��𾨖c��^9�i�M�ݔ��� ������[mp+M�Y���U��8S�.�zv7そ��+J��JH���{��ǚ��&�9ˈ�-�張J�7/���<-�f�[��	�=��!N��n����κ�+a�Z���4�^�2�g����Z�4���AFd~Ҕ����z��3.�ؽ�'��4T�͊�����ڻ0unϙe	���	�{�]�؅~N��>��g���������[Y�o7�����0O�c��f�����)�]a!b�y#��F�g�K�N^@�<C,E�X�x*�{�'�?-��ggլ��@�a|(Mq��3�z�]]$DX]��ݫ7�P}��ߦy"ZE{��E$ɥ�Oey�5��i)���s�-l��Εg¤w��Q�E���4�>���s�n#�5t�ZP�sy4�#��jY,�e��Do]d��r�F
����)��<�6r�O��v�4�:!�)m#:
���]6�:F�S�;h��h-�{g��Z7��M;.-J����Q�x�מ�f����Ҕ%�I&"�eu�՘}������ם2��ť���}x}�X�o���ZM�f�V��]�<��|�a�7�`���{���K/�<u���YR]��^|n�_˗�\�zo<�4�ɓ!�Y�G޷qW
��,�Kj����^��A���T�H�������M^��M�\;=�u嘰&ngV,i�?�h���=����&*���';�u��}�f崟�o�ܷu�����t���r̹	1��%�L�7���C���f����כ�۠�mA�a��73\�gwz����*ׄK}���>~S����]_�0+������N������Uvѳ/E��3�,=(n�Q�ѥ햭z��:��p�P{�WA�Yȯ(ںZ����:���l3딋���Z·>Oѯz�C��~��nK���ԅ�y���۾lR7��s��ӳ�&�q��=��!�e�ӹ��l��9o��`WqA�ee�E��i��R��
�T���5m��h�ξ+JY|i9�۳״��Xw�����&\��;w�J*=^���=�>�L	yG�)޼��s���w�>&��]q��3��f�}�P���Y{�(�yw"J^�{��S7~��Xqo�]�eM�g-J{y�.�'0�OYޥ��C�5C��Ӣ�Dh�|/*=^�g����5��#Il�_]�k�sE�\�!�0�/F�󮰲�4��&�r��->��>ږNj����<��y��x3vj�ˆ:�;�Y+V��x��������]�x8�M�ֻ/�=6rﶓ����v��:��f�ݔy��P��s�h+�Z�<29�]�lD?}�@�ޱC3����Lh!upX�$9&e(�|/�vu���9�k�!:��vB�b8�����3<�I<��M�^:f�3NϼV�kgY)|�����ٗZ����`�xu�����a��>�o�Č�UͿyk�k1F�腂���e��Yߢ�iնSݹ�}��`�vo���@�kBx	���P�(j����;���1H�a�{ �l+�UIX��ۿ�H��^�UrA���E�б�Q�Tol�ڇ~��$��yu�=��E���}Ull<��JRǭ��6b(�SUǝ u[����f^��qo[�vr��4�,��)��w��t��̓�:�#�JN2L�U��	n�����ӕ_e���#����;�e$[��}�dݜ6��46Tץ�������j�5;��.s)�,�'m+�����1�	���^�(���$!�����1v�����Һ�i�ֱ�\�t��$*�@tf���PF�b��Xޱ���P�/4�ᏧE}��i�E�a�u�br��B�*����k9|�.�'R�U�aU{�8�5x�_h/u,iaB;�Dt�$��N�]s]�)�3g�i<��	��[�˼¦wH����Lm�з] ��;�m3/W��A4d��f�:;�#�8��u�:��P��з�mčN)F��:P�v�ضrX���@L�{P��g`��
�P�r�VPm rr��W��T�!��>�\~}����:�Ajt8qݕ�b)��@�\;9�Ÿ�]�hy�ӘN�wm�ɀ�i��q��}��KI�yw_kyB�TW~�j�Ck���p�<�<�=ɚL�w#&a����Z��3�o*M��ѡ��c=��uŪ�U3wV�9Q�\�>L_rZf�>�5wRo�+Ltg���v,�f���3Y$�B��{4�0CCq�����Ӽ�i�������܆Cl�Us{8u�wq6gn-�'T%9����6cq̬#+Z*ڕ-n�^J`T�(e�l��cm-�6��Ve��V�%��*���b�,�Զ�)�2�ˉJ�Z���X�4Z--�HsV&j�-�U2�Z������E�,AQe0���%kG3��5Drf�Kq�)Z�TӎJ���4̵���Ǝ	s)��G3�[Jմ�3(9c)�6�i*V���Y\զU�����Mژ�3ʘ�e̪��b+ٌ ��^V��8�70a�4Y�60��u(76	���M���{�J�	5L�r���Kf�V��Y�'���[�MQ��no�\���2��KE�|�z%X���F��<�t�Z��Xs2�#M�q\�B��RƮ����V,��׷1�g/'J�Kb.)��Z����z"�ځ���'�ݿ�V���c��H��չ�ʆ�+D���\�|j�>w���Ҁ���K醲_+��4�+�c�xe�{�_�>#�}v�������}]���r��FP�f;wͷ�� ���;ݼ:�z�rZ���'�k_M[�囜�3�x�p\�@(�Y�����8߳u35ߵ(eQ�]`�:���U����Z�hG��u��`	~�d���v����*�J�cWO�ǣe��i�,,t��`p���)+�������:<eF^w��G=��}��f���U�{>t�i�K}��]���k�
.�Gi.~2%⫫��U����o�(�(o%;^[����*Z��{�G:���f�X9����9�� ���L(����_>�+�ۭ���w6�'��rV,5�r�v������M�������"]M��]��@�;�/\�ыR����Ҁ�:n��V:����k&j.��*�9�g<��t��z�<��3�y�z5�"6Ta=ܤ{}��E[�ge�+5;�m�Kft�tWiʾo�^�{�9���5nq���X@^��疗�_ؼ�;��<���6����0	야7��ì�
����)-]7V&j�͐��#t�Y�i��<��g9�����״�Xϼ���ʼ�^	�������q�,�]���G�!�^AyBb%��s-e�켧^��f�7Ă�I{��9�#��`��]���˔�wn�lg<Ǘ��{e8�(PkJz����o�➶�?,��[�)ՙc�6��z�82��d~촷���s�H��1ᯝ�ҕ�?jyot��]�Y�[ۿu[�yE�^���� ]��GdÞ*���3ⓨl�Ren�c ��	�X�BCρ�F�gc����%�n�4&F��J��F�Gjor]S��.��T��h��������g���p�����.�JOv��N7�XDM�x����P��-e/+��l6>]J�I{}Ֆ1�i�!���K�fN�lE%.�-�l�ҹ�ʝ�K�<$7u�QY�:��bx�*��4��+�r��3������%��e�t�О�^<tBKv�·%G�yd�x���soƒ�DI�+��	��bׯ�[B�8�h���Iec�)W0j��X����co|�v��ù�Kڒ&�J*�|6
�-#�5�=�HH])+5Vo��o=�Z�B#2��g��o5b�Vw��22�\�+x�^��ջ+��%vI��ʙ]�~~�>䫯&];�8�	�zO��Y�A$c�H�)�궍[l�;�d���ٻy3'M�Y��ړ{�{�k���g��ܚlS�cj��H�q��XwG0�o���J�=;EFO�Gכ9͎�Z����8N�ma��{����,F��te�~�n�_"��m&Q��+�C!�z V_@:]�
���Y��$�8z�8}[z����Uuק|{��X8(s�fI�5Sym�
�A�ѫ6��v#v��u��a�������꿆t[�RW��Z8S�Y�^�y޵�q7F^�,؞�Z����J����t��av-��ǳ���/)P�u�-���0��T�pL,.x����z���.N�*Q�ў�:�XV�N��9���h�Z��%�E/.#g�'��]�W�����w/��QCL7��\���-����]��u��^O��b�_G9ޓ	L�w��V������v7�ͅ�M%�΢'+��=�6��-��~��ѳ�kǪ'�^Q���쫜�f�{�|��sw8Ƌ=���F�%Bj��j��qG�m����A/1�q�mn����*������q�OU#����z�o]ܜ]`���1��.�v�X̥h�7��Xӓ�Jz8J�v?r W�N�:B���������'�T�u�Q'r��l�`�����Ip�����}�g��X��a�Ř�N�=ʄ��q��H�����D�Qջ�Dg��Gk(Z������Y��-,���t���^�Y��јߨ&�vT�W�7U��rap�9DWA�aC�K2�7�ns/5>�I��@�/���h�/�!��6���LQ[g8^�ު���S�(&���܂����γ&�'ت�X�s���O���l��I�D_+j�i�S�v�p�(��]����L�ǘ�m���Ӣ��]�������W��q)�b��x����WM���+מ�ppuZ�z������/���qv{���)�;B�ώ�\��6lC���e�)iiC4t�����MN��0�`�JQ^q���F�����^�6yd�mP��p�!4�x'O�K5��)�AJ�ʥ�={`��mxY�r��#~ 	�M�����u��$/�w�����L�f��O7�~y���=W�c��1;�7(F_;\��x=�Җ'�9��驙��	�T�w��Z4Z�+��{���JY禗���~"Gw^dm�f�^s5Wr�lc��1㗯Ym��O��)�V6#�"4ެ�97}��&/߇�����K��NqL�v�g |�Huޞ��/g$Kq��[p�da�N�0�ł=��Wuqq��yI�is x�{r�U�LX��{���i��j�9�'#�f�j�"�@����k���0
Ν�f���C;��|��L��~��U�a�&͈*���r�q�k=k��b��J��-�{��	�Xt�3�uEY��l.�.�48�cU��[�V���\�v]��O�W&<�yA&�	F�r�h`x�F���tS��b�ftQ\�.��K8ܒ�|Ec���9���x�<�Z3.W/qf�����qX�����j;�ʑ���S���f)M�X:y�3G ]bW62:̵����N�)�l��*��U+u��p�/�qރ!�Y��~�����O��6'Zb�xs��',<kf���&�u&���b̘�=���I��"�N��k�L`��L.�moaӺ @�����-�RD�M�L��Θ���t�ٽ����
[�Ne�uɇyw1�*��D��YJ�;L!��τ����S�{}Af���	��t�H��{ʶJ�;6��ph����}n��긃6�K't:�1�;�va79)��n�p��T����ȸZ�h�7��p��b�\�Q���«{)��H3;�ࣜ>t����Fx+b�A�w�{ݴ^���7����ƅ�f/��X �w	��r��{���#J�[�Y�{�NL��4�S�D�]=<[~6��ճl�r�[��ɪh����Mɳ%K[v��V_Z<��d��D�
�Ypu-�6F�v��B}3�z΅�6炃Lc�dwׅ���Nzwe��_:$nU�v�wú�:�ٖs�n&O��[���q<�����8�ò�{��T����!|I �Z|����hln\��T���,T�*V��e�V�(��p��]2�m6ю�ĭ
,ECT�TaTT�����8Z.YL��ShڹC�����Q�ƈ���VҬ�)[*[jc�TL����"V�V��+U����M��(��i����b�E-�hYV�X���QX�����U��=���<v�̵�hk�-������m���\Q� Z~�l7�r I��y�@Y�����s낍aĻ��1d��s�j���s�&%�,-����Jay�/�E����^����uڠr>$r���֚#�q��=ok3�(��eg�2���/
�] mW�{�'&�+}Zwl9ki�'�xT���e�~�,c���0�pE���u�&�ƃ��st���Y���x�mg6�A�1M�m���S�s�.v�=��w�Ē֪��U!W����r�=�\b��-�N�ʾ�IQ<����
X�V���-�⪳*���;�L)��M��5(��xF��ݞh��<۰��ơ�8�(���rx�/O׫N-�f�`M����8Ǩ�M����:)�^�"kY�[\���Y�>����I�t�.�β���񓛊X�j�������4g��x�%�2�^f"$aB���9�vk�t�cM�&�7^�\�(�o������������)_g�oH�+w{���^��l������R����9km�ҫ����Z�n�n��*WJ;f�x�����&r�n��^ MQ��fzz�n�ZR���>y���َ;��v�I�˃�N�t�Z�f-#�>��n�F�/��݄!t�V�}��-�w�_sOs��1��9����"�N�D�jJ{���=^�r���v��+���+�̽c��KwX۲�����*�<U1����{����-L<�dG?rx����m״�3'�Q���؊��G��˧�1i2s�ydvƯ�>]�{��Æ2��m���CXsʘ��*��1<��
�_%�|�gg^"�NL=�4�i�O{.��v�f�ltY����Ng{��<�;1��{�ӳ=�ޕBZ'�q-�C��@7|�n�W6�r�����z3��
���]^�ҽ��'�=,�9ը}��׌�^��ϡԫ#��L���z��u���%ry�bKL]kҬǻ"�[3O�̓
�{�Gp�z�W�^���!!�C{1��ю+�Z�&z�s׋�5Sۛ`�b��H8��roS���GY�^�����gt����J�t��b'��a�W�-rFSR��y���K)����u�ʝB\E�,Ɉ�A�$��e��Mi<�11�eM;N-J�s��J;k+�PY;��6�u�x�"F�ɼQ��nu�>4�/����Sn}$�6���1E�����T�`N� �/�X�����+i��y�u2=��2�Ť>[���G��r||��6�9lÉs�i����ggW��w�*^��[CWC/1�\8b��r��'������U�h8��o�&�|��Muѻ�HTs��rL_����ϊ�=�>�ϖ-�)K���7�ܰN#j���y��`��W5��k=[5I�m���\����6r��\����Wچ74ȤF��:y��:K=E[12���A=̃^Z�{LTp?F����^�C7�gۦ��%Rx����2=r[}]k�+�M``�^y�Z���8�g��-�w8#^���LzvL:�u�Z^�]�q+���w[�6v���Ƿ��h���5t�n�	K�m�Z���1��<��
�����D@���|r������`�E:����hǤ����u��pߌY���k�uxy4��^Ld��n��z@au߄�O2���9Z�,|�L�2�ҫruz����Ƴ����:B��B�N�=�[��zW1�h�E=��*)F|���+���η�w;���T⼠���ۃv���^��t�'F����9?^Dk�W��k�Cz&�r���2�����o�iB��$.��n����H�:Zq��w4B���
�(�-�n}�P�亃cT,��Y����L��9���^�%\��b�-�xWc���.;㕺6C��Gb�=f����������,�w}��!O��x��:���m�nq3}@&b׉����Ú�A�k8����z��r��]���ơ�ՎA��Wr�Y�:\Gr���|���
Y[�W���^�y_���a����xGf3�,�y}����	h(�s�	�D?:��B���˅�AK�,�6�
��ukL����ǅWOٕ� �-8B8��� 3h�/�{.^{�>�� <�wO�r�
�
�a�CN��5�V�]�(���JȂcӀلi����(ߕ�O{�d�RE#��|���aO���-Y��N�%C��V��]�k�ϩئ�� Z�{`��yq�n|�t�׷ךw�y��az����J�a~F�x�Ry��o{7����D&��Z�&g��W���������]t�Y��aD��$���l�p���]+�ɺ<e�%��qs����)r���u|�h(�wn��r�o��J}�ΐ+6j�.�/y���������W�굫����E;��^yj�o>f%�=>4T������Vsʁ��s�J�p����R�ە.�-�B�x�ܵH7��A���t^���p�����DB��YD4��a�ye�:ꊿTڛ����|��Ň�fǐ�� ]s^_G)�^�m��GEw���6�|>�6��9�Ymh�mx㠥���S������+����)aP�4�0�æ^�Ϟ�<�㇁��Zy��a�7���=7I�Z�M�'y�`�gAn�����������Kv�Wcώ��2y��pEqdY���u����P�;C���Ia W<�QC�!�T�Wb���<n�|9���^1y�̈́��������kJ_eʆZ,���7��t���/[�zo��(���a�Zv}�#D��ş'���]S=���0�B<��C���/��=4��j_ޛ7ޢ��KAr�SB����geY�]�����������@K��y{���Y�b���n��$agXB�����F:Ba��ހ����^rG�Z���CH�1���8~��g����I��b��9E��j�Q�d��V�Ӝ)�Y��>wF�/�K[��[����P-�ZUO��Կ_�1{������Y��³ec�[�Ϛ���#�}�Y��(�~ؾ�B�*���z�tv��C���	$�I,��QQm(������x�: ���~��A����C0����f���Fٜ�8�T��"�h�QEF�2���&����Q�]+�`���Nh���ᄤ�d���־:c�r�O`[-z�Xu��?�!̓����l�}�ï>Z�i��+�Z鬢�DQQ}�w�u���}(1C��*/�"芊���D�Ȕ�:����N������-�|�[����v�a֡F��T\�@�[���we�@,î��f��9�u���+@󅂫�جws����2L�fe��y]��ȤTY�H�gjہ�g��(�� ��Ț�I��E����!V�,�d��f���k;PQQv8�PDʹGfoz�m�A�ſt)������_�;>(Q��{�N�6p�
*/[��s�1���p�h�j�M���4"�p��qz^	�	����{�/#�>�0��v ���'���o��k�9��OD�v+@6"���' 䂊����Aa�/��PR��4<�ـy��e҄v�C��m�EQqq7ZI�@Y� n���ِ��,bޖ�D �:B�a������P��1b�qƎ����I瑁|3���~��(���.fͷ jL�QQh��~� �f g�tޝ2��o-2N�)��G��l���=��q�����C�9�;�)�^X���P
*/I�Û�FO_�EE޾F~!2"8�$t6�q��9�Zh
���<4`F,6��Ô�=�k��>�4���=�R�M��%7������2-��!m���3�,���p�R j��{=��h=�plR
����/������ �vz��EEֹC��(�A�}!{��̃|�O]aq�BA}��h ��-�����"�(Hv�Y� 