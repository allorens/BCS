BZh91AY&SYz3֯_�`qc���"� ����bA��    }�(})X#L�kMV��C6���V�!B�jVjX5*�-�cN�$��Q�����ֲ���Z�4"D(��&յo�s-��V̙UV��I��h���E�f5l�L�c[2JF���e�L��TV�C�1�f�b�J�`�f26�Q�mk[lX����(���լ4[h}��mUKmJ)�I6 �ٛM��!I�&�(�Ɠm�E(�V�Xcm��SVUK&�R�a"([h�2j���y����V����  ���>�ڲ ��k7�q��TvN�\�T�mP2��sQ�c�N�SS��T�Z�\umؕRvs`����.ҫ��jTPZ�#m����j��  >��TJW����67n�8�+S�[i���֎�SZw^�y��m�	��qꐫ�Jn�{�om�a/K�VtB�.��;�)J�Y�{�������)RmFcZ$mZ�fπ  ��׶�@;���(R�nz-Ž�i�m���;ڐ(*���yH����ohiR�{�e�[eZV�p�:���J��_w��2%W�O��h����=fi,��5Zl��J����   x��+�*���y�{WmIV��Ok={�^�-�<��u�C��>��za^�K������jUUqӺ�J�4���)�=�7ޏ��T}�T-���J����Ǎ��f�if2"�j�ղ�   ;���UIZ5��m�{jMbUS�U��}��wV�7xxyJ�+l��}���g���+����ʥ����\t��*�}{}���(	Os��v�V��W��y�{�k(On��굩���fŶ��*+U�_   ]�}��U)]���7]8EF랥��핳��{�J%QM���7����+��w�m5���r�P��/v�;{y�Һ�n���u�ʫ��O8�{eR��z*'��
������m�kU{�  �{��������y����ۭ�3ɺ�{e*7OU����-����{ҋf=�v���=��Tغ�<{ڲ�K�3��^�[{uֻ�m� :[��(z��kbb�6�lJ���&��_   syA�[w���·�A�w�7(���{8z���4��^�5����E��n)OV�z�\�Eܽy�{u�c!OU��ڍ�V�b�kU�  o{��M{��@���{A�מ�x� �{O=E��p�觢��Zp= �z���TWr��z��՜��X�2��f�Sm%m�
�T��  ;<o�������ok;�ު��`W��^����^�ˣ�,�6/A�Р0;�R��`u\�M� 
>   �   ��RU$  d@ E=��)IQ�1 0	�i�L�E=��E @  � EO�A%T�  0  	��T��OUT�=M      !%$��4�S�e���Dm'��������J2A�UG߈�_�u�c*�>���ή������ۆq���ӝ��� ��>L�l@}*�����
�����?c� _�y�	�����y�O�w�OJ ���T�ʀ�����_���������zS�0�ͅ�����0�/�0�L/�2?�ǦS�#����d}�?/� ����_o�W�+����a}���_��+�0>�_l�����(�L(���|�,(�����{`S��*	�P�ʠ{d=2�Tl"�Q��P��|2 �l"�U�(��@�� {`P=���@l����@� � �Ȁ{a@=2��l�������PC�"!�@�ʠ{d>l�TC�(���E=�"�l
�UC�"���d}��>�2(>�EOl*���()��ʢ{d@>���
{`@y�A��*�e=����@D��
{d=�"����
{d ~X@l��
'�E�
��T�Ȫ{`A=���Ol�L��P��<ʞ�S�
�ad}�!�9�=2��_L������}��W� {`� ���_l��ϦS�+����a}����� {a}����'�� {a}���_������e}���=�|?~�����=�������������*@ߢ�[��Ӗ�*f��o���Vw�b�dl���9��qlH�{�z��K97r��Ze��B�&ٗ$z�y���hn��x�Z�d�nm^HM��4<*�mDie�wZ	 �-S˫��(lˍ�^M�A�I2�e=��٧�+d�
0f�z6)�bܵ,�q�V�Yt��7�wn�y���"��t�P(]@c�i)3���W�]�� �P�o^P�[��#Z��K�f���̶hH5[:d?�5���ة�p�[vhd�:�b��:^]�v��n��sˌb�qe�13�I��η*|�݉��h�5nr�ϵ1MTV5���V\�l �ۨ hZO׃f5[�%�]�.��b9�k+["�(�j#4�F������B2��R�4����X7��Z�h��ǅ�5]���;�X�2ݵ��Vf�����*;4h=B�e8su�W�C��SL�n��`C :1=�aހ�B���;R���
�KuI{ܙc%1J+:��vj��&�,�&8�؆�a���VVFHgmY��z���Ct
��"��;Pt�%����LG�6dvr���!�m0tb��z��iaT�Q��v��@(|�W4Jn��0�ûTt����]�˗�V'�R��{X�ZV�Uo���S��5n�vO+{sRu0-dU�Ǳ��^ؐ����7�PR�X�]Ӥ�2�Ŕa�ssP�Z�gv�p�,�߃vŶ~[I����h���4fjS(�ڪ�Zr�ͬ'+����-�y�tH:�v��"5դ3��`RMV��:����}y�nͷ��ග����Oc�p[������@��kh ,mlFփ�լ�f�2��TB��5�%2l�,4w0�"���{@�F%`��D&�ux+QX�Q� h�
���fÌehȥ��W��1G2n�V�T�Z(ܛN�e�*�a���T��Gxw&%PTŐP�j��;���Dٔ�wL�%@�=ǓPe+B���sH���u0$�죧�".�wV��t^>�ۚ�p^9�;/	ʵli�&�mٌ짹���L� oeA3Fe3�)@L���uT۠[���(b��i;
�h���df�ر��Jb�tQ�,�`Ge�)�:��6��obT̸Ti�g0T���M����&5fXg`�^d.��o3d��X�B)��ߡ��3
-�KZA�O�8pX^UK��M�ڷ6��F7�eƴ��6��b5tk.ȃM+��b��K�ڷr�YUݗ1j%�r�iv�՞8�%���ӱ��r���Yv�P7qV�6���"y@#C+N�P�Y��{pX�7q]���U��t�J�`5y%��5���v�LӅugc���[�*3R#\����v��<AJ��Pvv��'�nS�b��+^�w5f�d����M�j�5]�i�6c��N�Թ@&�P�ks�J�O%l�*?Q�߭�Z+o%@66�Ĩ�, �ݎ,dcb����hr��wQ!6f[�oc�c`*~��E ۆ�K.G��V�Ʋ��J42Agu�f�K*k%+ݬ��upTJnVF�'ٖ�[����>ӎ�iE�^ԘFl��@Q�&�zk���3S2�X��-ܶ�Д,�s~t1�ي-YL:df�Ջ����&���nj���k'��A���:����4	�V�
��Z���q�zRա����	E�@�x�S�^��X�Ma�����E�[0���ՔD�bj���m��N��yi��iU�22�.:/�CQǋ0�Ά(%A�[�9@ef3H����T���Qvo6YNQ�]���Se_�Qq�@КP#�n����nT����+/f�Ww���0�{v2����obE0��U�R�9Ne�1�'u��E�/&6(���6E[P2^L+8r�&����΅�
�v|���+E�%�s�����#,5��-�4�p��n]M�R��%�dE6�(Yt�e e>���@��*׹�I�MՍߒh�Y���<�d1�+l���������R�&9u��xZ�f3LG0hƐ���ge)�%t�n̹/kC �C]��-�Qt�⑚��X��OJRt.ʰ����^<e�.�;���	۳��#1f�5j�Q��5�;D��M���[��&�7�,PCv���j�EH��/���,�J�&���0CN��r����� =qY�Z�R^MY���S)V����66�:bk�����QJ�B�O�GQe�uk+�&p�C�5���T��@$Eٺ:�v))�Q$$%�Y�n����D�j�hF#�t�ME]&!4��8w.�.Tu��ڒbYIT��8n�h�kG0��ijVX�T�\KƛT�eG���%-�22!�g °�U�]sIw�R֔�B��R�{s�Ee�s�=��MӔm钘�f��i�F�*����z��ôR:���)ɪ\9���#Xm�
�A��0L�k1��^c���fړlX�� AԶ�Q��R��u��f�m����N��ml�� Di�%�ٮ�a]�ŉG� �K�k��FɨhS�onPaV��ʛ�Xu8��{X2��s1B�̀�����K.TL��sB$W�N&���(�"1~��¶��^�ܟ*!V��#ivV=�(Zua�t����[���0��U�%�ÙL�T����3raj�|���p��V�s�(iL�4�	�^,�s�2�mf}�2�:���e: �Z0�^ҺY;��Sz�1�p����,����0@i���5�P���em:m��Ir�̷J�Dw3�S*��ZS�X����;������ØY�{� Z����6lÈ^�6�L�T�����<�D;��?" ʽL�Y��wE�jQ	m��2����֠�C �n�ȎV�gS��e�x��9c۰3��Ƅ�ǡ�}6J��S�B�d�6�ٸ����b�0�kuK!Mn�0[��X����䒬�,;d�6��Se����yO�n��|ή��k���x�I�߹��q��Ub�̖�J`��	��VF������	��PV���:NMY����r���7�8$u�2p�)�	�UC�X���I8�����
q�̖ͭ�oa��I}+��ϐ5��쟊jK8�Pi�Ѭ˚�-	D��P�glPA3J�'&җ[��0V�F���*�-ѳ���פn�
H�ӏ�C��i`c2�0b�����00E@u���z�;B�zW���l>Ӎ=�����Z�Y��4Y�3˝��XKas=vfv����5�t́�:dP���,� ���:�VS��Y%"P�J�޴�Pp��4�ڇ[ ��l�2}
č'Wi֜W���㖖�φ�E��\�4�1�2�[�,��]��k�Zr5́V���D�7���O�[JQu�s3i$�o�@˥Xڡ5ا�jڱ�\���[P�a������C����l/%X���@#&b#jֽ�Y�֕y&�)�C&*�WΆI��kP�����YJ�˭5��6���)��a~U��f'�"�������P���N��Y%�כ/p;�Q�,�Ȫ2�Ԉ�m��:��r���f�p��Z̼r̤� E�Y�����q�I�7N�
2�[Z�Ac�P��4����=�$ȫR���,Yѡ�S$��(�K��R��e��+dě��������ڠ��.�n��n�cw����CgT�M����{5P�մ�����ec���*ZcR�-�F��E�RBܕ�3�Bm�{���%�:í�1GBΌ����&bS1{� 5)PȨb�Z��K���6�a��^�o*�d 6��3�\q��_\���I�WX4]�u��vjڈK�p��G ���i�í�4�Mn�����A�,-3PiP��f	F�f�ue�t�V*���e�9��X6+���-+ʎ�����9�p�tӴ��;�!Yt)Ae�c1ŵ�;AH"��*(��P��u��{�a9,�d��+n�+3&!�����!_m�	u�Kb�;c�C�H�2eI�fj ���9tA��jmS�ֻ7+���VQ�ee�;��.ʛ01�U�� ��1��9��Vmv�C�wF�(�7�V�cp�"��*dH)e�ոf1.�tMY�Y�M;�4�qV�@�qY�U���!��u��i(N��y�_��1�̨/��h�{��mR�2�`��V��YC0�Ve����2rd6�(b�f�B�n3���/�Sp�Ŗڦ7j��TVL T�&�f�T�'�s��1�í �g���ZB�dn-!b�f�F�j��XÊ}�d;�c��2�1*��cʘ/K���["��%5A��#��Ҁ0]hh2+Ӥ�z/$iKG��+Za�Ă-�Ѽ�e�-�՚)����o\1ay�՘0�.2����x4T��zh6��{�Z����&�;�{�/1:�Ѧ֛JXQ ��������1��ʵ��L1�S6����0�H^��.ĬܩHTvT�Z2����@Bp� 鸵������%�DIS�����qu��z�<�4�?��2�D�s7
v�dL#� ݃6�f~:�+F��r�]�ȋC�N*WE��C�<i̳toJ7����e�Ǝ ��nR��42J�h�0�M��o�؍�]ON�2'P%�%�mm��
��.^�@c#�Sn��rܳ&��DB֓J�ՙ�[nf�7�O�Nӥ�;&<9Vڇv��t��;N�m�*6�jKji$�S Wb�RbVTe$�Bu�j]���^Ve�NISi�3g���G3ܩ�mg:[\o�b��ᠬ��mݵB��	�5�T����W��.��%����rl
Fb������
1�zX,���D�������:�ͧ�3�������n������Iwuv�Eٕ{3(�AQ5r�4�m��B-�]�����T�6v��*�[į��I��v8|�y}cR�>��5'��[�ʙ\����6 ���S.�����k;	�̔E��͵h34��єr�_d˖�V�)����z6H�)�r�F�L���w#��Hpk�D�OT���rD��;���v�B6l�n�wz�ƅ�1�^S*�d��mk\�&��5���SR�]H�H��$����M`T/�hc�2�4�m0p'�y��v�*]�N�Z�o]�[0Ѓ���2����Hq��m�l�j�ϛ�nLt�
e%�����#�1X<�>��wC���@��9@F+1�j��޴�ܟH
��c��e�)˖��V��Lc(��X��@�u[J nf�q�e�]l*�E��YWlDn�e��Lf �h+��[�݅Wu�Ȏ$i����Q��=ܻ:u%�D�f��/0�#�
��6���ok۷##*ava�i��F��0A�ɀ�X�Z)]������]L�״�2�&+�Y��8�yu�vS��$ٳ2e���*�[�����^@!E+e
,����5���9-�CS�`�b$�$8��)9�F�O+P�g�[XFj�j
�@n0IrHKB����sP�����ս�+n/�R��W�Ș��uZ��Ţ�E��'T (/����c���N8J�B��C�q�Jm����-44�mc�J��@jV�v�H�T�ž{ׇ%7) �
���	zm�J�Jd��{A;B���A��]85�0+4�1p˔72����R��L�Å=?%����W�5��r�{�u��Z��#��Y���ņ�9)�kF��Z"���k��m� �.:d��23��.�,ݚhА�֠5�����t(���m��>��u]t��ܷ5���rY V쿔5�HEI�Z����Ch8m��ꬡ-�`�z�ki�s	��!�y
tr`�CQ�9m�eLln�OnP�vd�$��3(�k�+	�� 3#O&Q�ӥ"�Pa�,���A��ѧ���O��U;�ܜN�n��L$��F�Պ5�6��qڣ��rƹX@,�0�Q��ǘ����h�0T�J{���p�7r3X4nȾq�k�!���!�)�l�q��x��X�sP��$�hǟ�����[J�%����@$h�ܙM����A^��d��n�&KS�0�,b.>���%{p�"������V�i�iq�M��F��m���f8�
�P��/	���k[R�
@�@S#e^��������]�X�^���fb�5�Ir
Gh}�h���!26��v
��mm�Z�3q�j�ׅ�4��.L�'
��V��n+x�q��v$�;�(2R�l6d�%�I�2􍺀e�\�ו�ŭ�.�Pɦ����R���@��i&*OE���R�;)m�Y՘r3fl����]CV�Q�W��0Xh݂�-��H���MMBl衲�Ҵ�r���n�t1%P=Tm�g�4X��ZG#�d>f݃m�mV:�9+f�Y{r�L�C0��V�BfA�Q�.�P���b^Ri!��e��gX�in,
�1N��miX��y�F��^mЋi9�����$軋�n��MY���F�f[��:1.��%����[��%f��A�����VY%oS����4en������Q奌�Wf��X��.&@�5MYF��nRڄ�&ޘh��4��D�,�r�R�cw �˂��0eF��S������S	�,Dm�U+D�q6��/h�yj�bt��z�02en��'-A�1�Ab�K���P�p�CI�	�xtIQ�4�5(��v�{����up���ԫx=�B ��*�ќ
�!�sw`�3I�ax^i���D��q� O��(�
�)���".o�t��������(a!�P��O�b/��(E�mU�g{�_��5Mn`0ba��*�h��uc�W�qV�`�U�y� ��0��D�����x��l]Y��9��}��������:�d��/OY�p;�\�@�t�W?�̏���^�oo��_�XZ��_�Ï�O��gy�K𳜿�\��MB��9k��<�Q@b�y{"w�j�t�޶*�]�h��]zz����sy�v0���\��c�dV�
�=6�d�q;�}��4�WyX�wfM�EJ-_M��\�'"��ڼ-3��.6��m�*��R�+�V�ٛ2�䆁�F����)��<5�Z�S������jb�@v��[�̼�j��{衬E1��[+�u�s�ܮ�X�]���yKqk�}��WH:�8��V���*�?܆N��f%�6�C0$-�VP4f�^^&YVz���׍���cQ��ڿ�6����8�]��Ó�W5js�1+�QZ�u�ˇm�5X�ˀ�J�a㴶�X�^���OJ��w#�u-m��c�k:�K���Yh��$�9,}�_m-.h��qm �	 ��g�O�s��l�azGe��[��|�	�a�rv �a�J���x��GpX��{t�����:�5{8�:k�x_g+�3I���f�Х��Y9A�4�Ih�	R9Zp�}NhCB0�ncJh��pR��5�����ċޔ�����N���ۙ5:��<�gwD��r�7�b��m������3O$;� m�-�m��tYgA���#:����R����;X��.i��`泲`��\�������{�n�@��2bv=�[�-@U��x�%���se�e\���YWz�:9��P�>9in�v��s�:��������4=���NW<�؞���=s�
���V0�3�VH�3i���`�9c�;ݜ�e�S���<���zF�V���76������[\�v�I1��/Uu�	A�m:�wY��A�5�F�s��;���sn)oo�ge^�͚E�iB�$�|�s��uњ0d]H�a�Q�9]f��+�(k��J�d��7P<�#᭡Ì�C�WpXR�Ij�G:�j�N7{�f�9�����%�(���h;�8uC�F֍�,s{o
su=�im-���\�8�$�<'&���n��j5/"��U/��We�+��$���Hb��M��t�\�A������
$�3f�c)����H�:�0R���s�%���c��,ؕ�k�0v�D�3��q�2�Ƥ���F�q�Q���]��g1Zj�%�������Q�0�8Z�*L5:�ލB�-�-<����}�5׮��OJ3F���8Ћ,�Y*�-�i5S=Bw*�����a�&vs�}1��W��lNHB8pg��8�If���g
�	u;��)+3-v9ɣ��"Ū{u������P�0GwUȡ�.,#�J��*��c�]q� ıR�-�6�ԕi�i�M��ܣ`�e�m�[J����J Blg�W�g.�-r]M�Yy�i��I�k�Q�VQul�����S��������ЏutX:k�� 
j�H2m�L[]�*ԓL{u�B�4'u"�{���Zu�Qd �q��w()8<[6nD��Myگ(N�BX3!�Lc�#����-�����p���U�rxv�%yv5)b��1h;�DFe�b��{�85T�2wI�VMZ�]e3�������� �[��'�c{?!�OY��w���B%��Q���te��X�W��r�s9���B9	n���ۂ�%
!i�1:.�#�ݥ����#WPe��N�f�z��+6�����#tu���>�����"�	Ȉl��mٓ0]1an��-%�l�&�JW_WU���6c	%NWWW�3������Nգσiw��WJ_*���(�0���řҡ	�6�,�ò�V!,��Rl��w^���;5>V�-X�0 ��q��}���rc]�
.��E��9%��X�׃E��}r�q���y��=$
1ߎ��9��q���+76��M+ǶIA�{���
E6n���/V޶��`���Yuc��;f���u�2�*�B�d��\��n�D���)����b{[�y#F��ąmӍ�3���v��+�F�wfA7[77'�Y��FDM����
m2\�m��S�y5����ns��F�ͭ�ρ�T��1���cK%L�HM/b�+*n^/��k��7�@�zkj�gh"��=�:L������M��U�K'R��渊xr�b�+��|g�4�%�7L!G9�ڒ�䅽�C&�{��s��7Anj8,�b�@ͭ�sK=L�h7-�sM�^�1�W�ܗ���г��O]��F�9�zp��y�.��"u��܎�	���,u#���	.�}�BWeg���B晎�KΊ��V-���ג��Wz_�	�J���¨���t�T����ѷ��z��m�weRV)���Mh�q�\6-�Ju�c��4�b���jv���U	{|�V����G*v�����v�ff�FT����bno�r^)P�B�iB%Ԗ�RB�c&j��yۼ���q�i����ؾ-f�<@_n�p=w�\�١��?N��dٸ��CMh��2t��z�=[���93i�ג����V]�{���
�Z:�Hy���y�Y�+t+M�v�iL�&fG���Vi�������VX�Z��3m���jW[�"��ʂ��@t������f�\��$�5l�7�9��ξʟ^�D��imI��̛!��hĻIɀ!3��e��j�jG�.:�蹺�f�7�׽��p�4��K�@![y�r�$�%r�0�������I�q�eqD�(n �3`��3bw8wI�k�����{Z4��Z]�zY�!���+�+���1�'ˬj�����4m�ڬL�-��닧�N�rȪV�}�<��^�����L/g+*m�+����z��D�:��TUye$�
�V �50��os�������/cٷ]Y�nP{V����}�fۛ{|����.N�z"�F.�S+���{�P�X5^���v=���d��LH9��R^��]ȃX��k5=��2mj&'W�m,�)<�`�9�=IwD,�bX�n���'��wHorr��I�n�J˛MV���V���9L�� Kc`N��9=�+7�ۛ��q6�7PY4��ߔ+p�[{O��zw��]1w��(+����\o;1���2�7��ӦT ��Iښ���U�@-��(�nս(U���o]8G��u�]��U�2�.I�/��68Z��Z	�[l�5����ϐu�<Ҥ�x�c�]�`*"���;i�@4G;�)<{��z�l��L�Y����n��p4Vt6������:�Ʋ��Hb����O�@��;e�^�z�(�Flqȕ�07դ��ɥ�\��3�:r���_e�ƫHGv�\سlBJ0ŗr[�]v�i�v�>�ٲ��\筨��|\Ȅ����c�xŞ\t���S�P����tS��*-|�u��i�P��@Ƭgv��=9o^���2��.�΋�s�n�����䕌�.V��f�:��6�9�
�Y+@��9g �1�v��/�
�p��i�f9�f��_������~�p�IE1];��	.��S$��:��ªʹ�%�v�Nk��.J�z36��]u��.���;�]���8X/p;F&Q�<T�Ֆ0 ka͋[����1�WfwE���Ȗj�s�V[��,�ז ����5�2'�/q��� �q:�%�=���#КZRl|*�V>��R���9�]���:
��*e)�����]�޹���t�F̬��k�^��h�l��S^`�z�n3��xu_R��ƀM�nƢ`u�<aؖ;����2].��,�ؚZFf5���#I�ʭըc|��zu����s�ٖf[�+���i�9��s�j �w���N�-i��;J`ogAYS�(�
��L-:�N�ʇ,X�e/�y���}ʂ��r4��X�[��(Q<�}��#y�Ӭ�"��w�/���9��]J�m�̙Q,�Z^��#���w���Kh0LSN�N��`+��+t^"z� ��@�#-E��-n������X�;���R���ݶ�ѝu��G��ʰ:7]��u���v�4ܝ�%�S11���=N���2�D2�V��:N��ê
��z�̜�xY�[�_3\�+�I�k���
�w�/��7`��,� ��OP.E ��ݗt&Ɉ.J5��/y�r� .%VŔ���ƴ��r�rփf�]�͚�R0D��ܔ3y��4h�Yk�k�L*e�=x���e{:�4�A�5�Gו�%p��w���a��*�1��=h�ݰ�Wp���@��r^LG�aR�Dۭ���/ٗ=v��þ�:�bC���RD`E�@�	u���X$+e���/�n"ݑ��1�k��;+���R�#���y�2)\�;9�g�����*Wgsq�8�욑_n��Zcɵ�KI�� �Hwʔ��/�[���7%�g Զ�7�bM��n�b��b)d���L��NsaE:c�{4m1�c�����1����n����Ԧ�z�;�w% ��Jv/��)�=�҄��I�P.���n2L�Wb�C/�d(��B1�p���[���.طR�H�8Si��uۗ�S����Sm��zCO8\!�2�w�I%��_�A�H{�V!�u��>��Q��0����[� -v#W`�� s��d��v����Ǣ���]�u��7,��Q�Y��y��x�J��|��g�V��{֬a���,u��*�.�bK�G<S�`
��e���E�P͚-�=�F��XA7�t���P�Tں_ZR|QiTg�V�M�g�=�RZ�PIz<TV�s�(eX�.RTk3r�����gp
���vw&�t�:����E����eo��Ɏ��)���!�Y�sr����:@�!�dV��zK��U�z���6��Z]YK2�C y7��.���vf	ˬ��������[ ڲ��;�L�WS� �K���څ����I}ReuK��J7r�,�*,�@`�ʓj�a�7��c�c�7�!�f�=���w�J�@�í	��z��ν��Ų�ȻP�n��@�v^��+	���J����8!B\+D�'����O+{�������Vp�y����F�2��{�*d������e���8]JP��^��>,'ll���Ӳ���7���}���~��
&V^�<!
]���(m�-o<����	ʚ��GJv�eF�D[�s��U��u��hR�^�UԼ��eZU�^]n�������۸����A�91��z���=oS�V���l�Un�U���b�Hh�uhJə\,
�	��,�N��x�a���"�k��/S��ւkm^W<�7C]�*J̥E�Y���VpJ��|�R�;!]��eFk���n��h�[Z۟��wVsΚ�ؗ4ʎ���Ϭ�T&c=E�JSYΥN����EX�Pph�O��f�ȷ@K�U2Cz#�K��ٷ�26*WJ��
I��s 9Y�y3V�3#.��5��H�ñ�W� 
�D��
e�ެ��E̹N��l/���up��4�$��eJC1�0��+�����"�2��R�q�!cKS�!�*�LI�e� �p��w�PT� s�����0# R�>4J�hZ9!��]b�����r��q�}.��:�L��c���w
�pǘ�e�a�'�#��Z����u�L87m>�R�	ludE\��n�R�ڻd��T4.�ĝ�}�1��iK��j�벲`��3L�����v�q�뱬u �Rhs.��2T2�Aed:G'q�O�k�r���@`;x��W��!��2me�]��![�:f�u��k��xWIsZ��n����)iu�jW-(:6�5'a�d���[N![l�q����-nԓ{B|��g�N��:\��t�gD�"6�wk)�b���,$em��i��j��JȒ��U�.�;�	��v^T�o��$�֩9���F:[݂k���Y$�s�X�G�u��F]��+H��>����R�v�Z�SYy�fIG�J�Pb�%gR�;����.�{�v�n&��d�h�ڨ��Q��!��Q��&!�l�0�Q�n�mͤN�fS���/�7lE��mT��.���`�%a��2��G8�}���qӜb�kIUaq=Snl��!�e̛�N���'	�DX�T�<�X7e���*� K�t ��5;�U��Hkc$++�l����ak��c�ө+�X�Fc;;o���`a_kSlxd���:�ߑ����"��uoE�'a	#p�&� ����'b��g�Y�3]e<��wC2�ż�e�����{\��{�=�ʆmt�$\O�[�i���z�R�&u�f�IEgJ1���6O�6�c]ܧMK� �.�i8�޺�K[�X�ژ�ŧpӶ*�q�n��T�
��뵢Y쫵թ�u� �f�AKt��v��f��Op�
�gR�I4�4�S�;��R�<�'n��˭St"orԽb��~4'ƞZmh}O8(^n!�7�D!��vٺ1R����2-��r-��c�Ê��S��G�@�n=�H�K�9��pY�j�(��ѽ
m����f�Hr�R�w��Y�4�}��i��� ��m��&9�a���f�rR͊��Z�ãz`�1d��`@儣J[Ŕ.+Ӵ�>a^˸Mܑᖅ	�V���1�(�e�y���=yI�J�m�xgus�W5vV��Ku��S@��o��������2�䛘�_ZN�K�+�2����E��oM�u;&)�u�b��߄m��Z��O�x�8�}L����8;��e[�g��3�ׅ͒F�9���H�RI$�I$�I$�H.��J���]Q��ꗷ�~d~cC�C���|�=A�z���R��y�O#���$��~�t�7��̏�P��?'���DE������ࢪ |�?�~_�~?��~���*������q�������|���>y����|?^v����  ���]��H�HGV%9Tep��fK�:�w�{��c�psL����rb�
c�+*�m#�.��:��̫FR4�4=�� ��v5�x]�̓��w�i����fp��.ju��6n������UdΓh�@M����T���+H����]L���iK�>]r���5�P��w8�Y�X�v�P>����A���;i��
�L�����V�<4q��NqǬ�Yx/VD�>��Dt�I#(��p-cv�$̈́�{1�����_c��;h��5��N�K�����-�\iQ�y]R��]���[��\�@^����W3��s��`J��*I��n�+7��P�2率#仭�9N1T��ν�ԭ�ޕ�6���!�,K���f�*5Z�0�v�wKCd�	W7N�V�N��FN�<��bڻ�<6�R�����|�r�Z&�J�HU�)�����+#��-Eˮ=߅���4�7|a�p�|vD,�����gM�ՄOek�l	��'����s�˓: N�ϥ��pW�wX�z+Y��3_d`��R��Yb��pt�]/�*�5���2�ܩ)�:p�Y+Ɂu�wO	lM�2��.F�-k��u�X�s�\M� L&q�Y6������f�\	�]���X�H�ɢ�����u�wm,L����L�t�u�ƣ���a��	����� �Ip;�lұޣ�ݖp.�#h��$�r*�hV��������[� ���5Ρ�H�d�f��K�����D1��E��'EI�^��8�S��.�t:w�������yRPL[��X��x��1�h�F�;�2��w\���N�|��nX�F8�J��]��k�9w(�4KRĵ�L#/�M�{N��딜��`�����1q�Ou��g�^2�
�0��4:�8 ��ZA�^��Z8y�K�Bѡ����@�|�o)���n�\��r�Wm�sK�(�.]����-DƜ��]Kn�hOo�t(Yl��1�%�V��4A[bȬ�]�$�^�֪
�372���L%S�9��a�������E�T
TEt�]bXp�9��b���TU�EW��e2A��5cgpu��u�X��aL
㋔�Z����g�a<O�	]��k*�*̾{�3���Q8>Q�u8D:=ʋ)�.̮�l��R֪�b������I���Qn��ⷅ*|�fnk��h� ����O��b���ǅbv+d�fK9��%1��4�hVmԃձdy�����������K�����u�b�l�~��D;'ҙt��}zu+��O>�D$cz\ܬ+j5�(��*�8������K�]Y�"����+ł|y+b������YBU�\RC9͕eXV@ϔ�-��B���|�h��׆T1a�Y�� l6�%V���*���Nɢ�������_izֶs�b�l���!����%^$��L<��eݼt��F*�-���{\#��m
ti�����ѹJ���S�;`�SWV�ڷ����f���{[�w<im���X�V1�"܃���ͳW�M�kut}�o')�vf������(��?X�����5b,wE��je-"m��N*WryHq��R��|۩#�Nf�j���/���̊�L��{
�u�k�{��Ҩ+:��u[�d|h>��4t�����f�qfQ�i�,a����]6�c;�&f����*J�N���y��E�{ї6	RQ�D�E��Pݗy�Y!짤�N������ͳ2���Q�l��GH�
�wܯ�@:DuO����m�:-��P�i���$��ua��3�ًr^L�b��;)���)�ԩ3QS{��]4N�3�?:��_k�tjb�S�,P���o��L7&�\ T�uh@�����ܭ�!Pa�J���®�Գu)Nk��U{W���GS;D:��1��`'�p��JXusl!bj5��lE�ά���7yv)uAO%ds7�`�W.��O,�*��X�ݝmC�|��u��aV~�WV��Ƶr�펁��Cv�ٍ��=���k/�WA��7�ӥx��m��s-Z��ގ��X�3���O�x�s#�]�ԅ��^qU]&���-H��j�7�J��3�E�g� 5��\J����i7[o$�j]�b�L����x����������눃CD��N:L��n�5w�9�d%��#�Z��g��MieǖG�����}X�㍀@�Aˮ�T-��Z�������\��v�ؽ�n�T�t��%�RX3)s��$7�X��m��]��,MP�m�\����9�.(]yh�w�>� �䫖��w y����U1:�q��NJ@�%��k��4�T9���2(�� �]�H-'�A�f��	�,
jz��r�rT5n��IǪQ�]��f��J��u�m� ��}��Y��f���qͱm�wn`��T+>b���n�>�6_-'Z��h�4D�CSN՞��`քu�r�%J�nӽ4r�u��)�1�PGkN�d�~6�c�0����ĺ4sp,�u�WN�f�G��&�h3&�mI�Y�b�V]�w;b��+�w\�.�,�7�?k9 G&i`������Jj�&:�-aQ�!쮶s1��ej�4v��w���5��%I�RN-sy} �8mV��4g��l"�#J�ܯ�i��pd��9]�����x0���C�ԔJ�SV����E%�ǽ����,�W9X��ԫX��{w`H"�P��Vn����-S��t��+ֈ5ǩ�bLC[m��0�{z�4�r���CVb�k��#m.r�X;9P�]��ė#�����H}[i�уq^N�T�6,�7k��BJa��{���,�MmǕ�e�»jƜ��9�p�Cv�L�š��1ćԄ�6��^����]a+�r�ӌ�)P��9,N�qG+�=��oVm�iѣ7B��.w���Id�,tTQL��q��ܭu(I���C�M���b��������S ��/Eι9�Ȯ5��#��*����:t߻�@�&�<�{FFWBC�F��\�o[��xSw\�յ�.N�^e;3�'Wu����fb#�e��KrrMGQ$�͙����D�(T.J���ERw;-u��87X���6/�r��y�Tӫ���F0��o� ]�Fk��Ǖ6��[�(\Z��'�Y� wnkJ���%I�,P�|_V �Ǫ /F��۹�$mކ��s�$<�{g˗%��{FVڴ��z�X�-�^���x�w`�t[���LV��n�Qr1�AԸ�,hÓ�͉j�Q�N�gM�&:2q��ىo�b�q��-��Y}��p��3ת�J�W3�1|�ʮ��+�����/
�Ks�t�Y�I�4zv��+�}�ݢ6���ݘ�Cʐ7XgB��Ʒ�z�6:�Hڢ�F�,�5��3yM�E�0�{%T$���s3~�Z!5��WH���Y�8v%Z�6v���%�v��O��Ҩ�=���<����:�a��MeӠ*K�׈�)hvn��K�J���<�;/�x��ˡ�0��QM�����Gv�u��˙����k�u�M�+d���
�WVm���>��7�R�Tj��\7)����jC�����[�;�?��@��bT�g.�]N�a!�e��΋W����bV�,Y��1٬ʘf#I���l��ѕ}w��ERA��1hg1YJ��(�ǝ߆IB�`���m����ڻ�P���s�;���y�ת���I�3Y�1��ݎ{�NU+�-8k�̂�G9]8���3���Y-Z�"k��ge0�Є.��p�ݶ_*0��][�n13cu��vf�gVVF�5��¾�>�{�J�A�Me٨Ӥ&.:*��	��|͖,�RƮA�Ur��V�fVM;%t���t�ꙦP���&d뱐��W`��
R^+(����PĳM5�M��-V��+0��9{�+`C�VkdK�M���b�e�^���-���u��*��⑬�=wZ/�*�X��;��ΧXT��(Lt��� �bM����H�8����PZnU��Hvm+=T:����vV�p�Π�e�ݭ�cZ��V;��Ŝ��ْ�36F��e����yYB�3�x�����O�
y��˔꧱u���G���R��0��i0.���-�R�*��h��u�"�N�F�EP���_bw�n��-�S�_p0�=h�u�N$L%�����V��E�jy�JO6�=%;�2VU�S��<+O\�wh�8u�ꏧ\�/.WL:���/zGg)ܖ��fq-
 3�z��xĮwۙ �	̊��5s�賴YGj���ݪ��	1�wa�f�����''<��jw����U���ۗ1L�֍t��B�{�2J֋���&|�cM�67����(A����tW[Ys~����󶮘t����a�%哒V+�R�E=�)�WZ�F�X;X�����M�P���C�k�!u�6� [4f,���Tu;����'�'���d���&�Xx��XE)�u��o�k"�F�� ط����%�yp�U��Vb����`�4*1`�����}O��QT*�ѣ�����͈f�#Z��G��x���M�.��?�_jR�+�
���,���+4wj	F/C�u`����{yP9H�*��Ü�*�*X��0(�J��i�M���uq� r���X��G�o�2���i��0<��2L8�h}Ϲ�Ԭ�B�B�ۆ³u�e"�o%b�CP��G��n�-�yױ%�k�T�(=���ߒ��v��1z��e�F*u!�yXyv(.7t ��W]�L�N[7:��kN�A���G��A	>$�	[{�}{��wQ�;xsJ6�p�SE��"N�W���֦��EA/�pA��䬻�XY��}|5�m۲�2�rNj���x�R�.j\���#�SF1�Q��k���7(�(&U���w�����٘��:RN7�Z�u�2��mh6�pU`���T	���V�K!���Uˠ�Zհ��u�]\�tj�\ޱ�w�t˭ٵ/d�`�yU ;��w)<hl�����^N5�u�+�iz�z�*NOk �w-���3�	��(��x4 5jT��׬m��T嗜��v�2�J���줄��DJ�g��7�+%�rMS��wf`4D͊ܥ��a;9��@�|m.�����.@�T�v*����Y���ȳw3bTe��ڸ�,�ՙ�.�t�W56�xQdv1������F	�O��x�;�l֭� �bO4�`j+
���8q���p��b��kv^�hMQ���6{�9IU�'p<{�* ��g^�R�=�ۺ���u���)�)4��/������9��O�!�:���v?h�RY��T%�X��������cP�1�M��n�F��uk��e�m�4�a�oU	A��\�˲:1f�j����lrf�YG���=�m|�˭�5`*�.�����`�M"v2+{�e�����N�FA-	�a0$�+0�C1��5�VM�Nu%����6̱H��r��z����|v^_p���襻KW�,��v��a���{ӪÔ�X��O���t��R�}X�컧�nhӪ�A �٩�%'%�l{�����ڷ3lK�n�Z\���%��僙��9-+im���0���Vp���"�Ko�էk������z�+X$�[�ƶ9�_�RɃ�c�D�!�n�'mh��ׂ�°�T8/
�[(�Π[�Eͽ��
�٘��3��I��Z��	݆�$����9��K�
�
�4�����Q���Gz��j*���Ŵ�c����O�ӻ�S�<���՚�u�<�%��Wh�[[ǯ����9q(!h��L�޳��#]��:��8�b���\�m�_��9^����n�����ׂuP�*��%���jb��OH���X&��wq�j_\}B�$U��؏\�,�B��")d�ߖ�����ۊm�Ǹ达��.��)WZ�2w,i(�V���\�
�*Z"��<�>�ٗϝ�I��X!���{���ȝl�y����zb�*�a���"�V��`�(�G9J\��Nl�wt�j�5��jɘ;�N��k1�ǫԓ�����b@���/-�$m�b��;�J=���Z �7A� ��ޛ�.�G8\=�&#��Fp����&�*Q�zJ��PK����0S���7qc��ė:�`�ml��ñ/^�w1Ӏ������[�e�.���@N���Cx-�i�CbZޅ��wB����;�/��9�ei�Hr����ߊ��Y����� n���$V��H, �w�Sos�-�2J�n�,t��FӁ�4��qJ���-�;7!���"�U�R07n%Q���wW�z��P��j�A����˾)��/7�1�J4�֝B����n����$�*)f�1L�r��Z"�sn�Q�:��b<6�i�!N��Kv����_g}Od}�����N�|E*��X�d�u�\�NS�cyV��e�2t��)
�kz�"���WNbM�����<�%el&�gm+��% z��Ιo���I�,���i��lު�1k�fɥ��r�+�a\��I��,��e������i�!9pxѣ�� �t��Q̸H��)�f��V�X=���K�κ�]�-r�\Գe�"���L�^��$K._=�b|8s|���]�Xf�9ڌn�:S��X��v��D=yGOh��H�ԮX�qT]���%Ӱ�UD��"a���`��V\����3bQ8�m�.U��e��\��m��IÄ�z�R%�tx٫������ϋ��q���oe��:�۫���D��ث�T�x8�nh�[��C�Q8�T(o+o�-���r�]�,^�#v +�t�l;Q�?ܱ=ss}V��O`�v+��hbVD��H�����T _փ���_��~����/����?������}?��?O���������~v�>{]ۊ-�P 
�]&�A�HS� ���Ӣ�I~tO�J��Ii�	�-�A/�%$�U (�e�}do�#A}�W�d�`�׽��ɾ����%Ճ�ݑ�F��4��$�V����Q]�m�z8�o���Xv5�Zd�%,��/��7ϕɏ�'����-o�ڄ��c���f���������w��\ѩ��n8U+���q_uk@f�>�`�����wu�
m��_a)u�	�JWٵԵ9G@�|*>��QT��/c�s�H��1�AT�9�Q�6w#�w6h�$U���Q+�e=�N�ƫCN7��0����-���Q<�y��Own�� ��C���R�e�B0��Yo&�U�-�J6�v�i�B5L뷐r�3da��/�ӡHf����r٨�C��P���7
x���B�X��K�R�ue��k��ޜ�[� Kk�J����2ིwc
�tr��u�i���6� u�n�nv��u`�uT����-���ϛ�m�T�u�������i��q]!-�X�ERi��h2�j`�_�K�T��rS@:�W��So�gp�/dY[q�Kˑ�2��Р�D�[�U:�1,R��h�\���QwG���T�׵�^�	q*�9�$��=�1�9	X�/�]n�K\������G�f�:	�Q�du�	�F(l�7/�͵
,�����psڇ�MQշ�5�����J�J� S(��6i�i� E���J�M�Ql����%&�,�i�%�QD��	��b�� tJ
M�	"�"��J�%�1���8�茗bۺ�n��c���d0���E��PD��HQh��w^]��'�b+��N�T[�#Z��]��[[uưIE[tn/�Df6�vź��٪��ݫ�۱��N ӈm�Ѵh�5��`�b��]]َۜ��v�1���1&:�3Phz:������mkn��k��ة�-V���k����1vն��Dth�g��6��h�)(g�;����u���QU��Ӌ�wQ��h�1�y�Ev7�X⊤��ѵ�n��UQX�:�w]�4c�j7mj�']Ƶ�#����-u��ƪb��v�.�]����Qv5Uu�Z���;f4��"�d�m�4�jѨ����Cg��mEIDU�E���h�S:�vj����$��bb�S�j�q�u���#cA���kN�*(����cB�_��?VV���K����n@C%_���mz�]g �cS;t"\+��2��CW�W?��S��0~�)��Nv�Z~_�:�J�eP �S��@��@�J!0U�8�s�Q�WP��X�h#�I#v�$�A-�g��+z;=�u٪�m���T*���vx��۹��Jqz�$:���W������+=-{�������s�`|�'�k@��LG��V�?C]�1���Qg˦�r�3�4���{;�1N�S���[cժ��ߺ�׏��{�t��L�!��)�����V��)~���Z��oO����d��gS\�;"�8��5�����ګ����Z�Vm�#-9��E	iz{^V�st����UcH��y���Vl���Ɵ��S��E��ֹǞ���g��|��=�z}���ʱ�{_;�+�q@�N�C�T_���U�A��!V������lL�4� v38k�r�ӂ.]�I4�b�v���>�<��u);�����q�9nx�K`�3;%��c���%�qC��חP>�K�W��D�a*�kw���Џ�~v��;��Ţ*wH���`&���4�V�Ň�Ӭ��z��.v���)���&�u�;��<�ܒ�-c�ʓz��Z�Fisv� 2�mr9��j�#H�CֻV��e���wb���l;�lr�,ږ���v�-Z�8���02�βʺ��Ջ��'�/_[�S��[�mze}� ��[��;1��F�+Ox�svЅ3A������
�M����x��wuޞ���� ��1r�[����|��V��A������z�[w3Z�����������!�m�~V�	0o�Ƌs˝v����0�{�M�Ӿ�ڙ��v**ttg���3z������g�?zm�O�z���g^��v����v���aA�QZ�E9�x�Sz��2��p��K�'��}��	|Տr��Ho�ЋѮ�t���u=^���5�E�kX�-�[�t�{}�'�r��o�>�c�n�F�^�/�Րw�i/O��^��c��}�{<��b����{��~�T�^��SD��wT��z{r:Ɵq���ǯ}Ǝ��v�E���YX͚��+ˁ�	���'��AT�Y�"���\΅?OE�Z���b�j�ۙ6M���ք���$�^�@�˫:2$;�Dcuہ��*Q���I��e[����(m�_>�@LE;NVw"��)̃qr�NO��'L�NܵxI�a���8ƝH��!��,|yX�MU�vN�Vr��]���(l�h�{����M��$гz�_d����.�W�����I����ןJ�ŝO�g�'�������?\K.N����wF����^�2�5WMߜ�)��N�����x7�˿9����1�o�5��W���]�AP��4<��}��2�e�/����vu���WE�p��G� ��T�⽾��w��}+���]��m��0�{�������{o���ӽތx����P�}>c���R�.y� 0C����5���2��Z�59k��ѣL�h<�S�|e�&c�.מ�L4����{���\b�)������;]=�	�&�ۡNOW�t���7�(j�_�P:���������OR��n����|PL�SF���f�m��k=c)�Fw�Q���3�Uf?"���~~}����dj2�0_Z�;k7mڎh�C������K��\�I	0�w=3��*�o��y;����;T���x�SA�&��U��dLeh�-Y�@����ے�lp����"��rM��wk�a�n�������6������یσ�8�kF�Da!�\�{���7�%o�`�j/�ӓ6m��X솻��Y��o�������	��v/����郸��,���a���d�*�M�.��4�j#��x�<�}CWxͪbL����z?rs|�g���b�זl:s�J�lN}c�H��L�~������������Ct��d��5@�Ƙ��0����Y�ޢ����<��fX�By�M���ӯ��|=�C���۶���_G~�ɲ�oX�ݑ�ܹ�h�d�`/o���2���ʺub���w��ٻ���vătv��~~ز)�{��a��6D>>���.��_�����=�y�7�Z��q9�����o�km���`���%��j��u���Ʒ�+�O���#s�yw�a����W�;���K�3�xE;����G�(��@q+~���}��y����O�Q��. T2fE�{S��u�6�5�ʗ��R�2�b���ByѭohP�N�!����Ba�ԘQ�LΒ��=Q��	�췰�S�k���N<8�M凣���߃LC�w,��[�����t���*߬�m���<�W#N��.+��*߮�.��h]$��=�A����Ti���a�#ZoZ�Z���V77.*�5YL�EI봎_��G�I�e_��	����?lÝ=��+}E�<��$�tN�0ڵ�_JZ�J��Z��cʴ�yP8j�;��Pp��¤�/s=�N�9�Ov*�z�W��_g�ٯM��,L��.߅��u���c� �d\�s�G�W�8̛�����榦wˬi����N����M)^�����oϲ�g��;E���g�v�&N����eA�Z��#����l�]���]�`��/J��U���>�_���˸����M�N?|�:�W�b�=��=��v|�)���[*>�ǹ'+]��_�#{�����n��#�����N�Ӟѝ����-z�ŵퟗg[Y�x�ϙ���UnN+]oM��� v�
r1�V�ҥ���{���y�����$S�#�il����nC�1��Js�h�&��Ji͉��C5lZ��fd4�c�-P���^�ƛ�j.X�N��\������M����;}����WAf�}V��ʋ�mU���U�<��^o'��h��̭�����~��X��/S�ş�x��矷�O>k��Gw���){;+�	Sv_
���DW�'�V�1E��!'��O�zeP5���Ԇ�딛a�W}k�����~v~��|K��'�ߧ�W�55����Ug��|�a��ز�;���S��oݟQ��+�ƙk7�/ѭ�
���E�-�l��YFa�̡1���ʿv��tU���ׯ����#��>�a���`�{�0�4���/���{�칵f���<���B�yO��.Nw������x��~��>�����i��˜���S���b��ޔ�ygl��v�y��sܾ*sq��o白a����<��D�~ٔ=]�m����^b�C�"��K�>I�W��ue��,ť�W��M*��w��h����k+�j�ѪĜ�R�� g<�LR��R�b����f>��C�B��u}v��'�J#�<��]��ml�M�Ԧ�s-�hu5G(�ٯ`������٘��Ư#�2���]7�k�K�E�qc~����㱦ߠ��Ɉ����u/`TQj�Z�^�7��~]� �<���i��5s�q��� n���j�d���j�n�|��R�{�3�k��W{����L
�_���9[�j��ߒ�v����o3m-]�����I��NX&�t�k������B忺�����bʛ����s��hF�!���=�OW�����z=�`����޼�ª�]�tA�CGz漫��Sh��ܟ���2�	ʦbհ:vn��c�w3���z/
-UqAm�>p�ϳۮ@��FS��Ji��Հe9%�������U�Gx Ŕ({Uo:K=ѽ��y��f�N�~��E��'eW�e{�ܯLy���wՖ�����{��V�3=+�fd��rjn�3��z_lu�'���g��A���j�����5�ϒ�j�֪G&Aڠ��I��@��L��N�p��g�'^]�Q@\�絙�a�7�y�t����Uj>����TQ�v/��F�b��'`�D��#q#�]�Y|2e`�fZ@�VA-_6$])���\x�����;O�Zj2'"9.p'$�]mCaiW� �U����~���ן�m%����˓��q��reA�"�i����>�M�3�#���-�P�R���RyWWCU�o�=����+>�������w�[ܨP���}P1{�o�\}o|�h�"+3z�'�b;;�<6[1�}����;L�Sq�������Q??{7�T��Hr��g5{����{W�5LeI)z^˷���
���97�o��-l�41n�1_l����^�.����Qx4�٧{e���'��]�ʏ��`\�לE�c}Uxo2�Y�D�l���-��I�Ϯ�*{�;K�{���қ&F�;�C����̥K|�d�=���~��S3�,�^�h>������y�#��U���FW���|ۤ�y�	:vb����}����2���b�M�/x�w��T=����ז����q`���~۠(c����͐��+�٦4`�r�v�2b��c���,�x�o��`�B?{:-��b��V(3��SW�ǅP�ٷ�LP���fd);�ǜ�K}8'��)����L%�sA��71�K��v����(5�9�X��s.!gVk���5�fVrou��D� H��*<�7�sD� ��=r�]�@^g����<��;���3����n!=\�=�~�y��o��������})P���&<0U������$�G���6OV@��ߜ%��s"����Iֶ������hì;�^�g�5��I���92p>�m�O?E��s�P������z:1�w�]-���@bXa�elԞ�l�=%�����:�g�i�2x9$�&^:F<��0�0y�� �B�30������J�ΰ��>8zz��w=�������UA�<Ũ�U���|s��1���E����Q;e��E�ǐ;x��#$i#��Ndl6 5�x d{uS S.1=�����/�^.H㚫9z����2����m�l��>m>��^>��,*�=Ac��p����[\�x���c��w����.6F��UMg���c��y��=���ȑ5��nMoW��K��lO	j����F�Z��%�,ިJڷn��2����.�Il�[���
����qc� �e�o�w>������Y�:�rjZ�N����5R,ݤ�=���;�d��eZ}4΍5u:�ט[P�I���/�<���We��Q�ͩ�j��Z�n윰8�٣$�{6��򽦶W<]�)�� r�U_uQ��'�{�
;�S��^]�v����y���=��wه8�'�G��O�����ʹ��O���j�^��拾r�^Y�=��Sv޵~r����do������I�tj���xfM8���ʚ�w���\�N��5����t�Pû>$����.m�}L \��q���,�E��Vx3��S+�/�c��~�x7P�zƐՐX4�����_^>y�/E2=��W��sh��Z�1U���g���h�E������5~�GK˞��U�K�N����_��TCOv���V]L~������CX3���ǲH�g'K[t��!nY��}鵔����v�FL���v>��d��S�-c�����k��B?�_>39��@����_�{=~�_�����{��{�|j�o�s�/�<M)&���R�s�w�`'B��N�j����U�޾����]������)Q�Kq£�wW�	��3chT�d�Qb�^���UIρ��V��oCt�R�u�]Ѡ���gj��e������ى2��D9P�@�2�Fuw
�dN�������tlv'�*��י�1c<VfuJ�^h��q�p�9�2��۵����*�p��]��(��ڂ9.� ��먆�wo]�`��s���&+Y��@�a��Yc!���lT�[�wf�'UC#��XyЬG5�Sj�]�x�;�y��ȫ��"�먓ቻ��±�ЎgLSPW.�D+r��O��h��w3�ײ�������a�e��ӹ@fWC������'�Tv_YP�H%�/���V.F�o4�����;Y[זJ�\��7u��L�e�i����׌ſutpDau��E���ˣ0rs���*�P*�E�u$������$9kM�*��<��p�U[��v��0Ʀ��L��73q,/q��ʺ�!��2�aK���v
��˥�蚓�=���$K�Tb���i�H�rֵ�}�q�Y#8����.�c\�B�3&Ǫjj˔b�p��2_��5��R*'�i���W@��*�me_��uʼf�"l$l����[+�u��k��1������kR�m٬�G�k|��y���]��HM����塃.�s�^�������Y��a�Z���p�l��«���d���ѡ�d+SMg��HT�����T��p��V3Af��_�g���YUԨl=��{z:��2�p�Pi�Z�*qޑ\�DG��!�oo7�Ղ���U�c�=�g
u&7c�ѩ��Z��b�ꏌÏ��{8>lAY���كciq���L(+��n��V'�s���uv��`�|P]t�{��$#3D:0W	d����:�6���ڠ�C��C	�Y��}���n�R��@ɛ��\���Y��{�����XX�1��_&7ptS�:�H+6Uڮ=�
ݫ�te,0ncҥn�p�J�w0u�����k��7��5Z�R���q 5�p��	�]!
��cm�������ͺ1�G�
�s�컒Kt�:��\�v�ܜ�Tee�K�}�����ª�`����l�+ҰD�ܝ�P7�gq�@0^3���������1��ȍ�_L��+w	˲:�Ň�Izh]�K�0E�o_l����WmGV�FtB��>�-�P����6�-�\�Q�M��hW��.[=�rq����YA)��)s�p�^]\�V"�3c�����d�*��\���&Q�t�AM�of:s�kF
9, ӝ�ie��8� �@�絔�V�Ĵ�W�|/ ����
��|;��j� 0W{�����faK�އ=y�2�� &��Z3sX+F�w&ۀ�^�C@��:fi�n����)3J����F���ե�:���h  �l衊(�c;wh��U[F3�㋬PV��ݺꣷv`�jӢ����1��Tv�؊�g^y�]<�]�x,��w���c�G�8�;F1����yxlxo8����cX�j�"ض ��w��n;:�g����:���d���;b��w̕�w����v-��ۼ�	��j1A��=l]z/#θ�-��y%^^EUES�7'�<��xkĊm�y�y�{�v�qᎱ�,wq�nq���*��4Q�����5y��:x�������>y�U���ɢ�5�����L�ѭ����O��(���ۮ ��Ϟk��<7`�6�"�k��QT�cڈ��E�j(/<�X���-h�n�ѭD�嘼���1ASy>Oϗgt�y�S����1k=��]�T�U:�4G���j:��(���
H������|�ͨ�=F��%�6�v�E@EӢ��5��t�X�I#���Ƣ�ۦ*��^�����k˶���(B��5~�%�I�����%����)�}\�����b��5��I���n ��o�ц<�S90|�s#���.f<�Ⱦ(�-;�d`Ц���`�'bΥ�[��u̗)V�^]��N{{Q{�o�-���B�|_�-������v���/ ��D�T�p�f���� +~�:����آ��w�ޥD��)j��?(_da��}�E�UKV�O�;E(6׹K0� ޱѓ�[����X�;��rK	��KyRZ~�u���3��|j<|sm���^��_-A�^=�dv�y���cG�t��W\��8��D��J!��5I_�1J�k"Hw�#�NL}D�|~�E��^]�����9{�{�?8`�[�h��̜�<�/\a��A(�r}r2���;[{_X��Z�HJ|�9ݼ3������{����樤��Sm}�9���Ӛ�s��\zv*PG`P�`��ʹ�pS��������ҍ��z�k�Qqa̪k�J-98���z�[bn.\w�����bB����^�^1��*,���~\�����23�� Oݜ��_��T2�E'�JGs��w��97*H�/p�o# �x�
��!��e��Db�P�P��xͨ,��@�/y��(�^��x��r�pZ��v��8uaK7�hG*���=頉�~�~��G'�?j7���aά`��Yڅ���j��v];�ゝ��X����b���od��.�9�+�V�ÏT{͘'6�=MSѹ��Ū�}��Jh�G�2�]��=U�v����;|IAR��wY<�~'h���/È��Q���*Z�]H�ߣ���6��cd}],��u�9�p��#�����/��ĥx��`  �D��o*���s���ֱ]Lu,s��7y>:j�Z&Sxa[<НfǪt��j �>3�U�UT�ͳ,_���$1�x/��}j˔/���.�?ft�SC}�(��PM��/5b>�'�x�rƃ�ܿ�>�5V���E�d�_�29f���:��%��iM����@<�h�<W��6VS��|�9�y�!�+���I}j<�5��\��gβI��y��{��/��Y��~��_��.�l�����Cb,�/��^���T�yR_-�����?W<��}�έ^%O<e�y!3^�㳩��'���&G��)�(��Ϻ>:��J�"�	��UU��N�;�:���O�����ޙ�_nt�
�`���"O�k�IK��P@�w�8G�l�|��s�7enw-��vbU����o"���V�H��:��Y�/�\��Sl%��S�3b���ǴOu��{��=�nսtv����9/d�܍K����æ�iѪ{1��>J��)Y�������8�MU�ŲE�����</a�]�l�I�kҭ�s�)��6�q����\���X�uG�mj��{��-;�<;����`ہ�}��g������E��k*u��`Ol�ll.�sը��xr���*�q{��R����&sVh�q��E�G�s1g��gJm�H�,˲u��3��lx�_,>\��"�LDQ��B����(m=����װ��F�C�v&e� ��p�f��(�-|c]V�ݫ��xz���7g@��^[��I�r���������͖���?Be��{��R�t�#�Q\�[�e=�<g^]^U�LS�uR�ǫ���8�	NF�ʠ ,= ��gi쾋��3v�0P��r�y��+�ɗ�N�^,���P�ϭ^/�
�M`7�{�\JV����>�=3�u���Tֽ1���̿�oM
 qT�g�p>����w!��琯��˰Z�/�lx��ܬ�����Y����,�C4�軶�2��GN�oq+hg%&.)dp������x�=x��w��5�T<D�90 ��_@Z�w�);����\Id�R�j�9�XF�O.�tD^��x��tm1��j�1��DA���	�)�	�DH���E�"E�e����xnL}����^g��r�s�ڒ���9ϮTcm�M��;����N�4l��׺ʧ��jLN��stA�t���ݼ�W{����g�*�>�(����dW(
������#<v�q������Z��i:�R�s���T�lX�O=���5���;3��t@�g��'#|U�!�ǝS4���tIZ�B#��"!FQ؇���W���v�5��� �̎�?wCir�D0w��c�(�Ú��"4~ ���<ޠG�D)W��f�\��5�1��5���ݙ2r� ,a�x�A��i����<��au+f�"*#�mk��l4k�D����VV'K%553G�y�;��x[���]�+TcN�2�W>+*f������Fυ7�
/���b��~�����W��O��t�ֲT�>���Ќ� ivj���K�S�\~���
�yQ
~��kT!f)J��_Jm��G���qC��/�\E�#٢љ���r�e��Kv�e��.�n�wXE7��'Q�%�>�\��0|������l�ު��$h=F���1)�	T��ª֤۫��ɜ�Ơ\[ ��Cմk⯮�i���N��_�����lmjC�q�.8Ғ�è�������/��Wu��z|�5�f{CwQ�he�[��,��k�dMy�B�og�	�\Urt�K�>u#���<ݵ�(��*�r8o��w)���nU�3�ܛ!��Z|+�ݒ��Kl$FS�ы�a2ADZ������ӿ\�c�N�?h~�kkx]��帾�Pyt��7aSo;8�!K�X�B�4¶����4���4�7�y�R��]9$d���x�;zm�tv��B�q��u"��V��T<H�8��dW��o����t�pr^8��;�S'ou׍��[�/��Tn֯Mūr{<:3w;pǠ�d8q���#�@��*���T`�w�e��FX�wy��7T�E�{<�4L|�1]���W��Τ��>f�&���|�N�f1l����ސ���(��,��=G�R�f�0�������Z{.F�q��Yށ��S�{]yG�?w��u�ܐ�|�+��
-�
����w�H�=�� j�O*'_{M&2���ށF��J��轆v�l��-u����ܟ���?�}�1��C<�	9>���G{%���V�#�6�>�=5��&Dm�.�ϥa���-$��ߔ}���׃'�1�����B9�r��%����|�Y޿J�Q�䭒$��Lgt���.:���,�\��G�t.&�׮'�����u�I�������ݧ�i�[)C�I�C�yVw�0�b�GJ��B18��� �[y�f�[g%��s���L W�D�{΂5z�K&�+*�l��w[��Psq��+�Uk��B_�BL�|J�PVm���2[��X�(���q�P������{��Ќ0�-�����%��F�'y:b�Õ�-�2�m�.h�R�.Q�Lo�<sjc7�s���_g����n�쎦WR*�A�=��,�F%�{��<�ܙ�Ǝ���x{�H7W�)�ݣ�|�&����o��|�����)�T]�%��6�е��O��)�j���W���Kc�w@�`�ݎx�\�������ӓ�u���ka�5�Y�ٛ�2������\
��,!�����}Q���Ψgi�J�_��EE�QI�J��f���}���#e�|Ci�[�@ܛ�a�=����=>X%x3��,���(��1�l��T��2*wG���K}��P��3_w����IG��#����Jܨ�]�"yje�㭊�-	����(�ա,��=/^.SJ{H�e�Ϡ�),��IKA-q	��5�y���M^�fcl)F�y�ۋ��"�ĪL6�{_��k��{�p��G_�>�N�t���a��l)7Y���nJ���\,QX�^GOX�'�7�cc����/5`�P��+��4��Tܽ���0I'A�H����BB�/W�g���y�rqx�w��i��t�P׺N��/T�A��_�<�&9SR��@:�/@F#b�P���p�~���{�:��?g}�/���d��m��0fo1lbkZȝ2���.e��C%�ѵ����<-[��Kz+��^���(��bU����Wv�Hr��>Y.�fҽ\57�  �}:���1����QT�n-���kiM��*hjkp.�����T���~���	��gO/�� �Iĉ� �_���I�_�8�,�T9 7�Z���Q�߄��~}�t����N[��`{#F-Lm�ɴ�j��M����?;�T��6������,~����Ǐ��]i]�޽;���s��|Íl끫t�C�X�(5C��6hFA��5��RR�҃Җ/`���ِ��������H�j~g�_TE�/������p�N)�y�
����_cɈP�O{��U��Ž��wj�3Am|������)U�dƞߣ�Y��&^�c�k�c����9\��b1g��n�ӎ������C��u~���gJ�(Y�6�k�U,Y���J���̸u*�F��iu�׾����ke�]鄇̑0T�=K�˲��2�q����"���ۚٖ�2�[��<�2�e����~w뱷>�Ɋ��
#�L�P|rܙ9�n���,>һd�Z��P��XY�LS۪��`�n��b����2�8ƂU��0��}�DoF�3�ڦ2OX�^}ӊ(]�2aě�Z���[Ƌ$��);K=���wg��n��Or�R�#@�Ꮓ
��h�Qԇ:��WAwC���𱏄�����wQ��&�x��u-����`.Ss�%�a���q�)���v���z�L�Q�Ej�6��t�<W�H=��VK�7iG�����ϋ,j`L|'vH�M�/��QɒM���s-�*���mٷ���G������Z!���Q�ٜpaP�ŕ�P���8��S����=���}	���wZ�q�O�DeƊgL��cy�LƧ2��=}]e�~'
��Sѐ�)���L�k&�����iE�ڪbǞ������z`<x�8�M�Ė}�N���M�躨6w:���Q��"��� ی6�w�������0}_tw���@�N�yWҋZE��ldZ3^�riR��E��1֚��!�����I�fuR���hu^�h��_�<ܝ㭜��\�ֵ�v��GP�32}�y��ӆ�0X�4*�<��5�0�?������f�I�gF�Ƿ��"D+~�Bj/��ufԴ4��cEA�i����:[D�H��1�������H�0�h�\���H�8ү}4}��ᱝ�,Ÿ�-bʑV�!����I�_����"�÷!E������|�O��@n%^��\��=��
�RN�񃯞���֍��|�y�Z�sG�����;�c�B�k|�,�?TB/�*���~�En���E:�u�ݥ�d/b��틃A,<`�������Yíj�,����S�(��hq��n8��6fɛJ����p�Z���3u���>�M�D��ݦ��mU���g:�W�lC`pYz슴m^d�5`5N��N�/��t�k/���� ��9m^*铊�&2�.^9�����p%T��`�Hֱ��8�BQ}*�\W��7.�6N��2���V~�)�������
c�>W��M25�K=�sGi�A�K�^ ���eg������������z�����G�\{r1��!wzQp�T�t����9�?7O����]�zG_]����g���N��9�[A�<�DF��J����D��۪彄��*�=��_Q/�,�Z�US3}|��FS���G��Y<��bA^�������gz�S-��KSh:�KV-m�V�Y��,����C��.��ld(-!k\�m���4�B�㼠�&r�\��[y�;���:��2q�p��-�zI~^�,r���s��kP��.ƌ0i�9����`=7B�J�e��t��=̱���4��櫗G@���/��gی��!��&k�ƥ��P���LA;����י���C��s|3}؜��+�����緝�X>���(�N�����^�;�u��gź��<����v�PNA��e���Th�f�#;lCH��L�e���'���W��mgLM����F'q��(�+�՗藎ӝB.��*)����i���a2κuG�+��ӝt��Ԯ�U���ĭr�>\�W a`��.�[#���46ՑnLW�mZ�@�s���yXz!c9V�[���b�������n΍!���}�k�x�t2P�C?,�bmO?|S:.�.��̈�[��B�5*:��g��'@˷$�2Y���SYʒ�P�W��dE�/^Q�`L�Y�F�j���f�]����8>B�s�d�kג���Vȭ������	��atw�W)c�>�� ���)]z%��FǅYL:As�S^Ń���Y��̜��V��ֹ�Pd}h�)]�[�=����U`o�C��z/�?nj���[Z՝�����&)&� ��m<`I���v!�ð��u�fCF=sS����G�7��f>_s�J�	&]������s�ʢ�<�NN�/�G;>9Q�qO��kh�2��+'%��c�a�}� ��=;'�.9�=��r�݉Ib��t�5�ڎs���Y͸i��A�,[T��)e�i��!d��=2��^��Y���J6�wOU�MtP�^�gn�#�+�p[�~N��;aj�x=�=rK
�0�Odz
�Y��O�;&_:̚�R{[��.w�j3��^��4������YR���I#��4~`�z}޿W������~�w�����<|}��%z�ͣ�cⶲ�od���w
��3��0[�;NJNC�8���jv(�G��� ��K��K
�}Y�r����ibu$�R	��+������Sa;9w�k
1B �V�/�gJZ�˜�Ў.0��R��ɍ"�R�P��P����Z©3�r���aϷ�؅zd�j�g)۴ �~"���W\�a2�2*�@�$Σ!5�5������9K��t�Q�w7]=��'�U�1�|q'\��r�ed#��+�6�lu\j��y�W]�l���R�c��[U�t��i1��ѷx�]�ٲQ��2�k#�)���sf�^�����n��ˑ|�B{��L����"��]�;w*����[����αhm���Ӎ��[�J՛��R�)���o[@�������m̶�wNT3F.ŗ$��x�\eG��)gY�iIYy�%�N��`{���ɼ�rv��k���"ށx�Y�Rse�)��ac���*�^L�Wc�@��M�:�����8�Z�s���w�u��
�"Ƞ�*c��ZzVw.�H��9�l&��)�WN�V��ʑ���q#}C��$�#��4Fsr-t��M�f��Xާ��t��R�FQ�}���utЋ2����NY����{K�P^�����ʨ�]\;ܻ4�:����ѓ�h���l���7�[�Ɔm�t,P�wo��+������v^QVG7�}6�m�Lk!��q}�4v�W���Ma��%C{w}�j����#'�\���\���3ʭ[���%+��kf�K��2Ĭ�H�2�-.��t�AO�$R_<l��|U�
�M���x�j�Ʈ��x�Pwb㈜�)J��פ�b��&��w����d�c���9K�9F/;yG�'�i�=�r��!a|6a�*���ey�.�4��ts��{v(;p��U	�Ōv/�k��KyLPV�ʺ'�γ�c�2"Nl�_XN�;�N����x7#�Fء�ˠFR�i��+�Ŏ�,�mj�'�V<�%CJ�\��MZa+�}�P�UΆ�ݒ�x���wX���P��l�x�^�{���[�ɫ�[��5y�BohPU�m��Q���)��-�S%קb;�ۍ:���7	���웯�<il��r�	�|�݁��\�Rt��F���[�X�ѭ��&�msx���y�4l-���]� Ҡ2���dMfeؙ�*�.YO�<JV�X��I��Õ˃����*��e9b`u���˒^��n�E%3�a%V0��n��wP�IJޚe����os��v��E^W��y*�%�T��P���`7Y�C�j�S"��\m�W9���|0H��\)3�u�͔`��å�ruZ�]!Y�㬹�o2�ٕ�][Gx��W���
Ru��GE5mn�K�%�%�e�=����)��+HNt�%��n���+h`����f@�X�^ڲ�;ذ�p�o}������{����QTUD�TTG��UZF�1:7���8�ᆨ�S��yuI]8�ֵAUQWF#Bi��EEDEU%xE�%UThՠ�PU�����Zh�%to6�<ڊbb<��Q��k��Dx�h�DQӪ����E4���(�<؈���J�DE:Ѷ)H�Ѩ�*tb���E5u��"�:x���G�j�݂�ގ�"c͙����P��S���u�
h�vtb��Ǯ�/[�P�]�]f*��N�&�Z�*�D��[�����(h�$t�E!4URD1�5E5F�Mz���� ��ELMQTZuS5]d��"N�h)��EI%%%RQT��4URiv�F�>3��AS^F��)x�+mPU��j
���Z������(�c���������:wH��4 B��@y_A�PI���}P]�.j�ԕwd�b��u9h��e9&7Ņ}(-'A�R��rx+��1�J��$)���(�L�(�D���61ݱ����"�~(��o��?:t�l�l�n�P}��2��|<hY*S!l�E�([1��sue}��(����C����nXK#�����Z��a�Ǥ��ƇYs:�jFk�y~�Л�w`�^��?|)�s��Li|Zj �8�S�|���z<fS�4G���������t�S�
�0a�M~��W%�
~���)/��ߥQ�uG�8�l_*�Bgξ�'�gm}�v�:�v�Ω��ܺZk*������L��g����W)K}AE|kV#��8Dt\Y֫���4{�#=���$C�>��^���8d��F�R����tG�TH��yfE�ws���q�������ӎ)���kͺb���A�=$dX�9:��R�6��X��u6��f3��%�3�YX�@���2�C�"�(��g9z��`�T7�]�܉��XEo!ץ>�F_��>�L�G�,9�����S�.ÇIm���)�>�ކ}���5��w�iuj��C޹��������kly��`wm"&�}F,����@J�(H��cm֟�����o{��3�n�5I�ƏK�^�O�.kVE��[�6��ɣd�!X��͟/7ub�<����Eӝ�w$\����:�S�\�6`z
<��/���<v
�ś�hM�������Ļ\Y.���T�IAn:�j�:F��=���{ʼ$�=]�u��>\m��V�(m��keV-HQ��̑ G��z\��^͐C5�F]��\�&�fC0��{邝[(�\��O�|�ݍ�L`��.���3�&_+�"X��㳕*"��T	�-�g<��ة0�jS��29��h��
�L(�y�+������.D��g��la���Zល�T�ܟZ��(��R�a�,�����*�/�\Fu�K=qo����S�!l��O�X���eN1��tvq�vJ�����G�B��_D`�|E�3Oɧsb8M9������ �D��Q�����j)��%�=�����p?*��%C��rW����GKE O����h�
������]�q�k�~2Cl&����?�!f�`�Ns�����V�Y��Fb,���8�wF5���Fy�^�Ԗ/"!��ͥݛ]����t*�R+d�TZ�[�w���������XwY��^z&3O��M@��G�UɃ��/��z�V(|����_�\�37P��2}�cj�#2*��{A��Ԍ
�`��m�>��|hz��v���_�]`Q��7x��s!�n�;�g7���{�X�~��#��/4�������s�S���$�t^w,�N����@s�#��o��J\��uH1���`g3:eѺc����8�U}qT)ok��hu��svN��X`G5�R�bf\�����}�W���W��=s>{r���,&�Bj,�\�a�؃gfϏ�Xi������x�V�ڈ��nW�y�+H&��?L#�J$��S�z�})5S����2t߂g<=B3H�ܜۅ32]�y�R�G�:x%W�����e���|e��r��F�Q�^U�W�'��|_|��d���vp���ץ��������L����x��=��"�$���䨳���V�K�v�!��k�՝��v��ߘ��� Z��,(�&7`��<�<�m��]c
�Ê��ϚѠ��{�~D3��:d�����`[-|m�a�Qʑ{bS��Jn�+�߲?T���tu��ݔ�Gc��q[�v����	IC�G�}< �P�	������H�����0����9�ev�A��U��܈W0����l3�B�s^q0�������q,g�T7��1B8���78^'�kא��v�;�׽�{�o�
���(�F�BAO���Ri|7�65���xX�����{3Jn��՘Ҽ[Y{���*9�lg�(-+M�;C�	ޟ����A�
X�������N��m�u�=���[-j�t��i�I�����:��U;�&`�:��AۡyPS�{����r^(���M�]���Ԋ�aZT�RJvje:ձ����jn�z�d̥���� �k�[��̮��fSM��#m��w�� �L����ʴ�M
4ϟ�<�cZ<���.��v���?F}�ug�2:y
<�*п�"k�D%����m:�yj	ż��^S��5��-=�&'݌�>hf��a�����
�a�\n��>���O	\C�2(&1>3c�����EӨ��24(�Ob�ť��g������-�u�iD��z�"}��e���'}�����v�(:.�9W�N��_O�|1Pbk��:�AVM�yW)KL��rAW�5�MFe���>�ʩ%EＭ�9����5U�a�s��?@�Qhk�!K��k���B�:�,�EZ�W�P���C4^��ї;}�8K
B*�w�j�'�����w(�{�$T��T,�!yȸ�}ӷjGV���j]�ę������R:��է90Y����ߛ۳�N��
y��ea3Yv���u�f�=�����F�j�@񁕅�=c�{^�1I�:��F)�@��{��/��k�]{�bc�nMBy��� ��z)+5-K�ײ82�vy���(��9�G����tTz�І�
řײ�_��p��Ȭ=�=��o��� ���x�,M���@�]2)`b�	u��\[��D��S~�&��)p��
L�^��CF��3���k��%$	��u&>�M�+�]�p��v��ryZ5cQ��q,��x�o����qu���qt
�\�
���<Xڽ�:�����F=8�5����/�k=��UB�1�����8�Κ��n�>^
U�$<��nr/b}�c�o>!Ր���@���huʺ�s�������+��PY������R��>�5æ9�Yh��ڃ@>�~O .>�b��Q����s�����mK�s͚����c$ͅ��ő��B�s�oH�ъ�ʄҟ�2Yn9�@X�N�^��wm��n�E&�*�����L���@K�~/t��#��S[�U&al�BzfϢ���sP;���z�R���bT����}]��*b#	����e��;V=7�OO~��qڌ�n�]AF���4��j��y�����S/��4c�\��'�H���/�}~��b���htx;վ��.�V6==��(�ť�#�U�(z�/)ΊJ=Bj-V��Ɋ9,�Nn1�)����`8��O;{�GR͸0	qKhr�Ԩs�p:�3�X_���OK9�I���W����^���y�U6������ʹ7���BD��&V�+%��W�7	�ݳ�N%��=��|_�.���8���zgK�|m�+��O�����X8����I���[�~}�t���O��l��9l�M�k��^���B�>�"�n	(�B@sm{{EǗ�,G���`�
�3�^�5����ݗ#m������z����H��M�ǆ�qM[p>��UW�C(z	B�����6��ۼ7VT&`�NZ�1Xixs�l5K�D�>9�*�H�ys�o71L'J��~�t ��E'ҮD�	v�3E�m���3P�[!�&u�>�G������.,���������Mz���;���Iu���	������Mf����ax�ڵ����iƩt���,Ѷ�X�7�i��b�e�����ױ��(�I�S���ؽz�(m�{[+�$��$k!�Z���G�4���j�;q�U!!��)ҷ���f|�)e˟���J�v6���Exs�e=��E���}p+�u�ΌvcS���z�<��aw��I�jS$�.�����!�K�/��l���ɱB��[���{)���e��yh�<���N p�F\�<ÁFK%���ᘽg�/ׇ}�{u����Yc��$0�姡-\v�mz���ӝ�@w�8q��Q>QYTp�e��P%6e��ȇ�_����Lr�"z~P4A\A0Q���jsb��tt����+\)�>�`�.ջ�i�k�ޝy�RN�]Zi�0i�qU�Ƣ�;F�ǒ�u!�Z���=r*�.v�!��%h���B^2ݪ��`g"�~O�w\8�����6b;ʒv��(�'�"uV�ھGܦ+�!�}3�����']�[����)h������Sާ\��2�z� /m�������x{��� xx«=��e�!��G4]*�mj��\���B�HB��dd��9ؠ����͜��|�fO4�憵�U�Xs��(��8�6�^K�<�4=9P�@�(��Kxg�^�*<�	��ڿj1�~�LJ6��'�
ˑ�խC��~,�μ?����T��-��Y�̐1�FՀj��Srr�{�l��PMd���uQ�M+�4����$s���4hw�-�M7���Y�w��吕�b �='!��y�|p*��E��<ݐ1z|<�{��s����ȝ���i���:ݮ�X��M��]"$�Gr~y�4"���+�8�DI��ݝ3ה&/\	����N���c<t;0ƹg�wS�Q��2*�{��H�Ia���fW9�P�QV��J��>+.�;��l�l���d
��bT2}+f�u�mk{h���&!Q��/W��E�^ĭq�1i�S$���ٗY�`�+6(�XH>�e�s%�� �l�n�)��*�)�q���:_�/��m�զ}�ϰ}O����元�퐺9��>P�#��g�
���E�8��̶Z�mV̕/�U�٘��9(S��o��T��6`Y�|q`�/����/��Ub$*�G��k��o�-�O��E� h����O{�}��9"�͎&�ogcˡ!�[�}�#L�I�e0l�V���d������j8L�9دF��V�������<�=��;��:��M2��Y���Y��(���z��϶�~��s!�&�`ڒ���~cS=nƢV1���f�5����=¶��V9kL!�U6U�x���o����&<������/";���&S�S�m�z����N�QtJ��8��P�BIF�� ���](�L��T��sW]ם�#�@��X�}
.mٳ�_q��w#�C�q籐���zn� N��A��!Iq�]묲�����m:�U�k'�k�
,�{ׇ���8���sx7����4h�窀�P׼du1�\U^��8�(��P�\�����C1x%�g�X�CA�OnY�����^m(�Y��ة�׷0�#I��dP��� ��c�9��C���`��F'z(�фZ=6a�"��nS�/�fp{Sɀ�,D�s(ì�*fL���P����͆p�i�q�v�S�[5���Q���"���]6�=7@Bz�}$��
�PT7,��Qg�br��Z����Sd*G��w�C.]��L��\��cN����\���X�@��`\��\�����{X��w�n|�xN�[��y/ī�`�6_��]��k�>Ϙ�qM{Ӱqwm.�V��b��ɖ�f��9�/B���/*���)2'ew/���T��]��q=}n�q)HR�^�6�!;)ڽS��GK��%2�>��eͯ��e�E�}ׯv��1�{=}����<HU��䚰hU/�u�X+ݜ����O
�ͯ@��l��)�H[>-q�ߌG0����;����߻�یKr(�L��P�{:,зY�;�9��i��!A�Ͻ��JZf��<Wkt����3����U�v�A�q��s���}ڨ[m�;v�)�PX��]�]��f��t3aۮ�0>C}���9Gkvx�G'��o˥��Y��]�U�����v����i�Q�[Fi�6wd�
�cՔ��D��.��-��>��vy��v��&�^n���;fr�U����Oݣ�/ +yCn}t �����!��J�<\O��q�=����LglF���}�)FE�N5w\��G��s����l	����H� '�=x��D���\�s�O�SΕԉ/>�R)�su	���FK-c�b),��I~�Nŗ�%M壎��DT�¯���K���ü%l3���JزU��ܝf��V�5�eVIxS�7�����eF��㥬+��u9L���r�.;V='��#����q�41�b8��É���g���i��(h���CSuV���g}�0���b��xɽ�n��^�n�n��4�o�r�`B��C��3u�i�s5�8�!t�Kى#���ȑ'2���e��;�
�lU�kg��"6���oZ�Ze���2��������������xx\X�P襭1���*k���y�	�
�H��>5!<^��{{y��^9���TyVZ�QQ�Iv�~�\Ǭ�N��g�m3E��0^���M���;O�b���1[ �&����~�9-���2i��������{�M��w,�*0�K=��VzD
~��q��T��m*8��Ϳø�߲����V�?4�6gvy�<d���>u(�褞��8;;؛�W�{#C�ҟ�QʁN}/ʾ�X��Cw�R��}�mx�o�N�O� ��f�+Bk����ܐ��+?0����P^��&~��3�"2��&�4�}*{)LR'���L��C��9Ho���s�"�gd�)��#���Y��&L���2��E|0V���H�Y��Z.]n�E�]x�.snEmX\]��a^Ƕ]Mލ6Ӎ^�)�M�fS���)��n��(싼ϓ&� �b�	9���q[B��U��嵲��}HQ9�#�V'��"��������qWҬ5IB�fuj�e(��@	:��)��§ܬ��N�ͨ�����?�����z�~�_���������z8�nx&1H[cr[��%!̝5,��[j�ܱN���m�����b�*��)f������&���w0���:�νF��N��"hT�,��ܪv;�\��F��5֬1m�KƁƨ�+������X��\r:�ś��T��B\�I�Hw:SzGA�w���ЫdѬ
��n���`�ӅE�:�`�uK��F��k:A���zVF�e� ��e�i�
d�䕣[�F�u]]�;d׀k�]�;�1l���sFJ���'y8�;A��@�jF�LO�u�]�|3�H̛w���.� ' �74sԲ�w�GF{P�����소ɒ�=��j��M�(�ڰ(]��V��|�}3 ���Yv�l<��.�h�V7�eD� u��-�+me138��oibV6yH�i|u��!�����-���E��!W�˝�Y})ł�NU�VV�t��4�(��kB�B>��Y�I���`,�x�Vtж�%$���:�g6e�y�������4�����T�xK5>H���f(�L�&�cy�e��`��ۙ{���j'�n������/d�h��]XaHwd��LY^s��ic�6�*IhʹY�dh7�Ӵ�̺x��N0�u KMf���R�#�� w6�ڽ��2P�ȑ������ϛ
gd�|��D�[��K)7"\�X�7hm�r��݉�'6��h޾��m� ��Yr�p�D��[nr=�r-�F�4���E��2Xy�s\xc�$n``7ï-��2�kE�<� A׺�+��䭉�	��u��B��u��^�*��1�wnel��V�B��rd��!���v��=�f�IY�J�ǩֳ��_g�vs�k� �B�������fE�ʾ$9���t��b�Ӆ�<d��na��.JB�su��4��z�]����������h���J�V]]���^i�L���N�t���ӗgTk@&��ݺ&�J֚�
ܤ�(�c-	rY0]
xO	r�;�J����+,��R� ݬ����壧&� �8�t�"��	�!v3��ݚz�^�7��"�r�xj���>N��]ev��`DRj����S��\o^bv4�������T�8�3�:�e,�;����C!�x��N s[ð��ܸkO�<w���|%_3��!5�r�m!��]Yu��D���(�TF��ia(v^�0������9��K�f@��փ7X6�^*�7LDZ�gPY��0�]���<FDXW�ޢ����W�-f/qD���W�^[X�%Yv`S��-hmppla/8�b�kHY��w�逅kmWM��aɜ	B�m���OV�|�����uA1&R��R��X���;��ܫf/;.�BEw}'0���5L{}������V�a�V0>�6'���0�bU��(P�?���횢�Mh��"��ii&��$� ��-I�330@i4UAF�����% ���f*j*�E������k��Q�i���V$���*��A�TAP�TlQ�� ���T%ց�ێ��E�!E4�1DUEɢ�l�Ew��EMLu�ZJ&��8��5E�I�E-$M&��0f
(�&�F�AO�T��*����E�0EW����"��f6����QF�kN�*i���z�����"J"�ABEMS]�Sv4D�]�@QE-TQAIGK��JB�.�������'w/UWX����&����u����(h*�%����Dw`�Mo8ꪙ�������(
**��45h�AUUM�TE���IA嶣=��!m��Q-S]�<آk̚�
�_������>}}yJ���i�gw�:����{0i$k��
���~�e�*4ؗ��ɉQd���I^�O��c���Y)ތSm���xx{�=�jf����mi������%�v����6�Y�LS��L�^�:��*o�X�4�nym��7tk(0�^��R�x%G��-�<�v5"�ݐhӋ���9�Mc�3�U���]d%���*}D{Q��Xࠣ$���Oš��L�+s~���q�Y�R�(b�.�1��G��L[�~��S��涍�.� ���D�Z�V�k^��,nvj,�v�Os(�<&r#�ڝ��-675���AUSkWƂ��`8϶$���(����F���Q�T{x�AKn ����4k���9�/��5�{�sLjO��O�R����h�=�؇���"����)�bj^*�Z�,/7i�� �?YxY���M���C��V����D��4�b��wKY���dc�H�q�B@���W��32\*��>V�m�BF�}�a�#A�߶�}���tA~ɲ�W��-^��; �x�s�J��b�vnh��3��ZS���f�hp{�<8\s�m����� ~�DH����2��0Z��?��������=����\��e��X3nCS�=z�Q��M���o��\�}0]3���ɼ�v�C������	�jH1�����jJk6\�W|ٳ��Sz+1J��ֵ���� �kyLd�kA�-��������>ʕ���e�մ���������f���{�IY!wr�[�+�����@�_�H�z�}�B��O���C�N睈�t�������ٻ��ʔ.
[~-]m�P���[4ˬ-�oiUt+1mD<�|w\��灨ۆ,FT=b#���It%�]�2F��6��������8y*�E��m�-]c�� ,��9� ^������1}D�_���FF���t!�~�t�1����4���g�<U[w���S��#�_V��H�Q�T�Ò���S�?C�����3Ր��^Cϻ�"��Ң�]U��K���M�[.�߱������f\�|j����ZlZ5���LD5�����ȓ���]��+��!��M�lD,�P���$M��PK��:�ܫ\a\�ˑQ���|��Tq�D3��37�z�C2�Y%��lM�}v�eD��^ZUK,q�c�Q�أ�-+Z��h�'zB���˺B���j��oUzV���N�9*O�4o����x�)�|�O��֮-��h��*C�w-�؍ee�e�LI5p��NQ�Wة����::i>�3��z��k�f��a�s�g��ܵ���A�Y4�,]�B��K�F���c ��$p�sW�{��]�ڝ��ú(H�c�A���~�^��OO��Ӫ��:�u���Z�s�av�K�?�}��ﯽPpzb� �>`Ml\oj[�}�W5��u����܍U�.'oz_:�[ =���  3x3}�`5�����y©$cD�2����D3lx7Aa"pǄ�_F;�A���Ǭ���a�sI��ʾ�)MM���	]�"�g�-�#b�AA8<�`�����k}���Յ6�b�f����ۧ����U���lmF�`�T�pg���\Y:(c���������1-�[�Un���aYƽ��f�~�vL[�H�$�]�	��5�R��@�a�x�|?��9�9�7�!��?ts&��ŭ�_+pZ���|N��Z��LC�p��Cu����˕K��픝:26�f�l{,<��"`�Z����j7��Nw�yZnd�YʈSh����SvpN�;�P]�}�!+6:�c��v��Mf�/�m�����5��P�{i;9Q�=��0�\|���_Xx4�����O�25�.��x�=_���}���ޥo�~�{�k�z/���c��i�����ǲ�D��3�Ǡ��q�ݿ�5�=N.��G.�����v^WQks�QR�vBT	z�Ŵ:ī�hk��F82�>W��}o�c�� �dg�L"����)u�7h@.��q���sx�غ�4t�@�R�܋½�df*�L�Nyb�#Lc,�7�4|G�F�2�JNK���8�ܒ���sFI2�\�Vof+v�9���W�t���5����{Ӑ�G����~����ŧ�]�q*��nQu��{�����(�~�PV��<5��m��QWWt�V��T���k���<�	8;=>��fZo����|ű�X��=5�N|++*]�uۄ��`��4�/y��e*�";M�J��mkgp�l�^�ޟE���ާ��,��Q��=�G������ �鍱�bxK7]����{��M�~b��Y�_��~r�'�W͚ٙ���^4��$NG�o$g��ƥ<F�=�>�^�n�ݥϸFb	;�볨Nw�G����P��(|U*�ʈKU�~�k�;��c9��D�vj��}_n���9Ķ�3�H��`��f��,�T9J[�
�>�A�j������ӱ�B�����ľ�|�#[��(P�'U}�F>wH���m'��\�����K�|kЌZk:E�C峟E�,��$z�u�¾^���bS_�pi��]��@�=���<a�q�(� 0v|O����ɞ��c>���7/Vr`�_|���"L�CmR5�geK�����h�ڱI���	E��ZեDێ3d\�]�]ήs; ���C�k��S5K��*�݋f�Q]�4�\R�0��>/>�]��M�Bd�U��L�uE 9��{gE���T9�y��U�[w��J��=���]y���>>�?UiA���(<`��<��t�^�G���a�Z��])ry�$�_�L�u��^j�r�X��ɭ\�k4�e�ٚ�:��r�|򖷃ܡ{cγP����"@��_P1m���iƯK��1�c�yiL���:p��Jvn�8Ő��E�(����ˎyt����l�k:����S�wI��XF����юIˡ/��ݑ��h��J^�a'VE2�tv�>2�]�mʛɌ�v�r�YKޝ#(ӛ�v��<9��� �+-��r�R��yHS��dW�RϚ��Y~�v7r��]��n��R�b=a)^��R��W�B�+1�ݺ����'�Q�U�;�vp�lN8�������o�M��Nz���	&�.��,K߳�`�.��\�*'R�g%�]�a�aj�y97��qH�Az��e��<��p�o��1D|WIky�f591]��}��z|!�Cj���{%RoP�#��A�#�漪����cyx�{��@Z�/T��K�
0�S���|w6b���3Z��Y~��h�}����(�Ʒ�5�����jK���X���R��A&�~�n
9�>���p*8�D�^�A�QAn�Κ����.C8e>�4��m!�A�P0W	��u��2س�fzܵG�/6r9r �u\b�	� Ç�ݛ���#�S���cJ�䍑�L��j��
����`(�JJ�σ���߯�����|�7��x�G�������۶�^@���wz>wL��=z��?R*�C�:���]ĕ���lr"gӞB�|�}���yNU�^iy4�66�T]w��^�m��ݝX)Y��W�����+:2�ҫTb����|�8�د��v@�v��r*(�[Kݒ4�l�^�k��3�k�H'�GBF�O��^k
���/}�g����S5�%�_�6	ߝ�Ʃ��8�M��Uؼ|Ս9�*贠ȥe~1fB���AO�u��ꦐgg�6�\׋W��ֵ�T�~���[�;O��]
�{Q
~��kF.�NL,�7e�N�]�iYz��F�$ �鵴��3)��UL���M�-�u�B�N^���s�N�y,;>����T@Y���cZEsC�O�\�nCG�AW�Ο��D�Ȱ�K=ԧ�E}\�]#��#%kR�c��9�@���h�g*�;���򐧻����˄z�f�5���H�վ��A�W?5�Lsux�X�n\AR@�����"��:����>�XաQ�jJ�6L���4x՘�T�+f11�ȸ��*�mB��K.����m�������&;��s���۶nA����w�vd��?��l�`V���P�����wUd��%+Y夀�]����o
� 3�޽̶}M4�xFu�� �7�<�>��	 ��V��F>���(@7���lH��R�N��u��F떦B:k���8H>C�%G�=�|�g�j���FZ�\��?Y�V��V�7Vt�Z��ĪK�6w�q籐��C�r��ހN��	�z+L�O���{U��ȾU*Z�R���t�E[_���~��KFPY^v�&�[��G��Mnl��dl�}�z�^�!� ��#�IpکG�yWة��;z��c݂g�l�g�l6�7m
��(;���f�I��u9 ��}"an$(�����Q�����E�Ύl�i4~6�o�f�x�ov��>X��"��Ft�P�������3Y�'o��4SR���gm���a.^�Pg9�<��
�7P�}�R�)A�o�k��c�$Ģ�)�����U�OZ���w��]��`n�b�僴��F�2�]&��%��P'U�O6A{F4�LM���)����	e��%��O���J���<%�9U�F��a>[��5���dK��׾��Ɉ^�+L����,T��FMH5�蕯��2b-D�m��������؝�yl��e�l�CY!�W8VI�Y�[���s��>m�%�Ԡ��}y���6���zuվ�~g�\�}�C���s�2��y^��c���JTy�jҭ_<�eڇ^�9���x��C����:!����T�
Q
Q(���l��X�=�k΋����7tK���.�e��N��6xeb��;�b��z���I���}�<6.�@�v�4�o/��v}��)9�#徊J�0���q̑��u�(Q"VOK�~=�����6����Qi���
��[bn.\���3�SO�2}�W�mb���UGol^�fYʡ����7e�*(:�(�Ĩ���*��t�h�pdB��,*��툨c�Z����Y��A֐ڊv�o�&�s��3�F2[$�c����:Kf��J���u�fU0,�N�����Jj��,��\�����4��L�Z�=9��2�"e��LN'���ޏ@��,ŉ#�"4N8��=�R��/~��y�vq��u)�_�k9}�f����H�P���<ڶ_����4�u�WkA��Of �\
��>���
jGOz�e����5(e�˕ۢ����R\Z����fy�{	��$�~ ��'x����{�&��B���i���J��ߡn���R�d������3����ȗx8���l=��M{4��?f-�گ����a��.���y�W���w]�;�Q�p��������A3�z�0&�R"oTV1m�����F�JǶue��:�"l�C���E6�{5^��OlE�؝����k9;�ee ���[i\�b�3f|��y�}|y}ߒ)�ʍ�B�����Pu'R�V��S^�3[���#��u߬��J��$�3�r�DY��r���t'-�es&��ù,.L+��C�&,����3��;�S8���k�!� ����罝�Dp�ׯv�Z���Ǜ6�J�z�����(�̑��3/���=6������|J;���WSS��S��҃Җ'����TE��e�Q֦�(�n-�Y�l�>�����`�P���;i��yz�~����1��4������+��|Y1����;k�;,����L�N�b�D�ưL&\��)?_���Sx�nS��wdt��o��-:Y��W�0�ws�������R�-�&E����މt���W�["i����r��z��zaKa�<J��k�w[ޣ�0"�W*�S��C�`3_r�^Ù��k(�\�c�}���]��.éZ��/�.��S0�x��Da�	���ܴb��w�!E�Y����^�|��zu�q�w0�\f�#Q�4�{>�(G@�2�+U(�=R�������<����*�a�.?�x���9�6醚`��\�2,M�a0(�[������p��'�6f8���\ظ�W�9�b�$�R#9u���.�k2��];#דIe�yخ�9�'{*U	&�wծ�@�`\m�'���,���k�q;�嫨EXl�� Vi����y��7���y��S=��x.2Y,�|)�ϐ����Ҭ��Aȝ<1�m��?v� ��ڄ�M�Ji�;7��е�2�S��.l��`�e�o��3K��~��Lfzn�YZ+�T'�r�}B���'�7��N���>��t��֡�1��f�|�^�^����?�%�7��݁&�#pȐ &lй��U���_��k��1�o�y�dԖ�&��Z��^d������i�b�/zDL��U(�i,(��P�u��Do�e�ag�`c5ڀ����m�8^z���=-m�K(8��4��9�3�"n
~����
o�Jw/�W%� �݆�S��>�R�Ҁ�$+��4�6ST:ajt"$윏�7ҋ����]գHyYm��ͮ��w	�������i����<�n��C�粁W���%����:o�="�Qx�ß��a�Ld�պꍜ�!��L�#��<�X�k�"�=�P��%�	J͙���ϝ�C[������%S�"�*�M~�S�D�b��˪�O�mK{'�Y�w��xoW�����z�~�_��������x�=�3kJ�˿I^KE��D�x3�e�DH(sgW'B���L6�iݯ����}V2`x[}FV�1N�delݪZ�5��a8Vc���,Q����=RE{��0�ڭ'���,9%�H�ʷӎut�f�ӎ�ҵ|�����zi.9sfK:�j�K�֌"�L���{�8Ոd d�ͬja��׼��� #�m��%#�GI5�-	}+���M��T�XE�*����5{����k+�L�l��`�������&�֧������cxH�wP�H��)��l<���{�a[�^���-aiz칊�`ר���� ����i�t�C���69��W��L6�%�66�U�8f@Y|�hRQjp��(Q4��G��[�IZ�dw���l��8d�*i˽k��%\��B(�i�q
Yj�m4�b�y�puN�r���k.�\3���񁸵N;����|*�t=K�Xę09�K�X*K2Ԉ-U%,���t$�-�\��9M�ƏV�xjm^�����"������%i2Yޘ�1|�Q���ya�v����me^
���j�W�;�R�9:�%n~�n�,�4�Pʘ,������L�jV���R��<�>���PR������h���ԭ�Z�኱�r����9�z��1f<6�b4���M�nP�boz�뜯�R�ޡ�Ŋ���)M�Y-I��/�v�7�)��(�����t'�4+�=l��W�\
�30��z[�s�'\V�'�I���WGG��]����*SJ�������7Q��R!���{r����e;Wj
�h�7r��56�p�W͓�j��R�'e[���v0*-,25��:�\c�.�pΚ�@򄤘�wфcA��ښ�gAQi�R���V2\U��36���)+�3k+x陽J��������F�k,�y�M��ݔ�h�E��zU|���Y���$�w��p)����K����{ [��J�9�t5�r�cM��=����+�����ٽQ`F�uJ&�KQ����L's�Z�6sv�B��]K1�.Ɍ��
/o��l����8�^*U���Ў�j�n�­���4�^�Ol��*9oj���$�V�b����Rt�ɕ-ۺF�C��\)u��0����5�!�Σ]R.��G���0���"�[5:�T*otO�0V�j���=�O@�]6��:�^$��)ף��N�݂���#̬��#���Uܮ���[|�\@�ݩm��F]@�6 {(�j��&�y���$�I�2�b��:ƙ�C-��k��Mc;�0d�[������rkɂޕpݘ�2��T,W6Y�02�WM/2�l�kr�M����#:�&v�����;]X|���u�a��fJFt��(L.j�X����'����!����l�d��5/bZ:V��;�|�Uʵk0�V5Ng�AZƥ����}E7a�1�[�L�t����UaN����۷�AC^�Ӫ���4�@|xb�"
�hhi�(

*�M==�S�.'RER[��-��b��%ZtSEb�7`��ԞEy:[Ո�*o2�vm��y��4]����)
j(��͠��&�榊|�Q5Ah�-�݄�tU4����X�ЕCH�5Q=�I�M�u���֗������AII]b���TRѭ1.�4:4��QA]�:�h")���zJ:+1E��왒�t�4y.�&�(�-5TSAE3!��AERS�^Z��%w�5��gZ5M�KAQkEA�UMQ�S�P<Hqt&���.�OY��EPQIO�4�Ĵ���M�Z���!4=j��PS��h
)�64N�Z4i:n�Mv��Зh��*&��kA���^}Q�]ƌAe������v>�7�,:���16^4�e0��K�Y�7(]�33�ͼ�E�u�#[�&tB�;q��a5xnfԽ�+3B��r�*H �I ������͸ݟ��$&�<�~�o%T*L =�Ӌ���Xw���.�>P�4M��=�$����W�E΄f،��̓;5rb�v�8��Fd@�Kj4���\����e���s�=��:~W�P��dx�L's��*�-�Żxਧ���U��~�b��i�V!JTW�#��3Ր����/�V�f_)άG/<�)�<�û�������.��E	�Gޘ�kLs��A���Vi���	�KRuCz�#�皤�o��Gr�q�r����!Cs��f����ZQ;��1�\������m���ԪYc��Tsr��<e�G|�;Ӛ�[Ք1v��m�qa��?��P�<�j_�G�Gw��=�J�-Aeyڤ��h����eS<��'=[�D�F_�.F̄`xzо��x�3��scA�\���?݀��kquϩ{]���w��6���\�C����fL-88#��N�q�&�P��<����t9�ͬ0�[r� �v����n.�Dg;�F��L�zs�O��#�@+�Q�J�a�i�/�>���ܯȟ?$`�yk�O���y^f��u�ɞ�[y�R}6���%<:���|4*�0Q��ᕴt~�ŧ�Y����$P�,KpI�r�v��� �3�`s�,u���>�1,�L9V�j�6��}l�;���[���;����|o�^�  �ࠗ�]	��vtІ�4Ox���0y�4M�5�ӟ%7���Y��t�2�s�{�ʹ�3��[fX��{�c2���n�h(���,�25ِ���5\�-z��q^�>��n�k�?@�|uςj�W�&�#cTW���j(�L�L	Po]�"���Ns�`�(vh�y���C��%���Y�G�zE׌�iɀS>�܃\���Ѓ&�j%�l�5.�'�؀�~�b(�n�>V�k=o����P�Cܰ�����dK�"�ʾh�[@ߺbN=�]��@.&���[��n��W���1�E�<�n�8�6�E����+7���;Cvx;�	�ٍ^��j��?lH��@���0���!~�Jײ�ӓ�u���kW���z;����h�{����U]ק��<u����ÆLΨ(��׉��<�j~���`Z��Y#�\�[ux6�9�w�������Z�-ʎ�)��E�>3����:��nQu��{��1��Q��wI���o�rh�=����I0W��!{�i�2�x�z����u"K�(�;�z.SJ{H��L<q6e��+3���2���S�<��4��ǽ^��k|���SW��ɛnS��wrwq�<�{�Vtf-�y:��:�U��o�-\QK�EY�6�t���љ\vd�5Zy��c��x2��0�89Ʃ�m9͝Sn�Y���]!�+�F����(z�����;��y�������D$KHP��i����o�����N�|�̝�6�����|��t^��_=GB�V�v��Q�)Pb$nK�m��z)f����_gut��&� �5�R�g��*kj�	��Iܧ��{�����h��t��	841����uU\�T`hO@`� w��|�/���' t�@���cz�0���iΩ������Mx���f��(L��.�i�6�[�������K��g�$�b��e�.I��v���w���w��~"l�g����X_}��;�$�<�-��Dz߬���0u�E/-�TQ������aR�M�$8���<rY�>&ћ#L�v�n<]�t�~�墛ɴ���H�:�Y�t'$���qMb�ecuMk^9��M��o�nvmߡoT�͗�[�ܼ��q�� 
��Pk�#�}_�*��&3,Tu<��0Sile6�x��v��{�z��I�e�^��o�e
��SPœ�	���rAx2�}az%,���\���5��ro�	_��-Ȟ6_�L��qMV�����f�i�R#~݌.hl��3���M�Z�1���Z1���+!+�wg�/��u�L�T�y\��+&(�S���.�X�z{vӊ�|�Q�¡��ϭI֞��f���]<����YWY�&��RU�v�9Q������ȫ,�NÔ6%�Μs�x�֫���Sn+H	�I.�hU_ʻ����7����
�/�ԌӬ}d[�u��E��@�U�g�2[�L��Tyo�k�VH����
8G����>=�j�=K�fʀ�|xn���;�i�r�^Ù���qE����~����?A3mF]vG��o���lB�gҰ@Xa�_)��)�)���y8i0�jS���r��K�;�b1��8���/��\a,[j�#P��}0�*�<������@ޅ��Ų'j���dZ�p�Y����@�a8��Zk�QD�&CF4���*�K�'&wB�.옫���}H�V.�#Jm��*�am_���ʇ��*� � ��k�����^j����b`L��yc�;�����cq(�9~g�UTp�{�N��A���C���!��+to?Cѽ��2$B������w�iL�8�3��`�}x3���z���˖�{s�Ӂ���	�S #��e��U��u�RTU���p�����];�f���{����N�7K2�U�O�%.��+SK�s�"D��!_Md���u��p�����
��-����S����'>K`3,�(Ŧ�]��Lp�UgA�����WG���$���#m{���x�2�׬;�8�w��Qi�knQ䰆���F	�q��{wi԰m^����Y�NlL��v��}}^�������R "V��
�(��wcJ���3u���lD߀lH��Q��9�W�0�:�������@�ME���-���S�3S9�g��SX��P�PC*E�NP�X�Q>�B��"iC/�>����_�:�E�>Y3s�1��YB�?�pt��������~.�&G����X�Y�^H���R�#�%����2��
"�b�k}�o'�K�ŔD`V�%�s^,z�P%K�;4ˬ���,Y�cx@6j_��Xm�|u���e�	�Lz�y�:��_HkV��J��Kv����x�􆇾:�અ�Ce�5~�����N���}r�T�e��^s�!Lv;p�"����ԫ�����5�f#�/lU<�c��m��u�L��T��A+5r����P�Ⱥ.K��ƌ:ω�OdT۠��Urp�T����iz�P󗋍ˁ�*@]��(��D��m컖6~3ϥ��4�>�n��<�A���#�#x����	u��Gs�VW-�yrJ�&�\����N�:�k��s�n3RĨ�$DC:��;��Ƙ�S,Xc�EF�����k\�k.&��m]H��[���u�FGi&�`C��͢�%u&e���zLx�Asܭ���]i1É ��J���V3rν�7�G>��Cbj�v�dC8�c����y$y�֢�N��a��p#v���2�u�ʈ���2[�Ϗ����~ ~�M!00����ކd}_D���8��|�<����:V�M�����G����0��mܪ"n����Z��\"����rQ��8y�U�w��j���<w��]�4;�����ɗ�GB��.�Ro��E�{��澑ީ0�k��/v���G��
���;c�x}�"�D�T���w���\ds{#�$hh��i#�@�5$o�A5�O�ό���߲<'��V�dYŶӆ�
��<��7��;6ķ=�{��x���c<��
�7P�Ojr��ǖq�Q`݊��2��R\d'`�К�c����/2�Z��v� �A���^�F��P^�Mo��ـ�*�r-��ゾ��}ES��*��_q�/�r�;�<澾����N�󹣞d�K��Fvf)-�y��x�z	��� ~�`f!%�T�595#�=��Nr`�o�lu�t�޼$5R�ƥ�*�x��V꜇�dq��ܟ\����M��1�����a;�.Z�7)o4�޺�}/%�:�]���"�W�s��ۜ;
�acc�BJ́��4-��l[��Ui�Tr���fs4i��"|�ꗇ)����ur)6f��mU�[ǜ�:;yz*fĕH�UCO:�O���ڹWY:R;�F�U[�Kj����jri�G�u�����ub�ؠ�p3��N'xn��8��;���j\�1խ!��\�^��S�_�/0�f�0oy�x7�4�����Ńw�*u���%���Tu��qu�SL5����=��g�a����7W'�����5����E��d.�q��t�F�����EE�QI�q*�Œ;��E�&�U�`���c��;S��ޜX�r] �J26�J=��N��/��q�?GC�;7��w��ؚ�*�+�:�105 ��2�G���T�ޱ�B�W��I��d���M)ʭ�1�+�(a��!�0�=� KӚ��"R����Q�p�������q�w�Yc�K}�q=��y�;��sH��⤴�,��]{�\}�Y_gut��$j��@�gƾ�a��E���r�C.�â�í�J��0��Z]B��Zht�US�@�v�$䂷�;2<����wY�Z��{ʦ鶖����r}ŽJ�599�;<^2��q�a�h��&�C���[�0,���{��t�|��a\zT$/:�n�6ۛ�����c����
�Mq]�}�Ǫ��[[�^���JY�	��y�o�E:�Վ��ݵ��!+uw��3k��$U�Ó���^�DNud�vVR j�^��I�"�Z�M5ql� �c�xf�\���a�oO[�s��t��fqv!J��[���`ơ)��v�:p��GTCoO����Y@��[�e���7)��������GJ�I�#���;'E��G��^�>~�~�~7�}��?����B�`7�7�{��O:Q�k�R���t�f��}{��B�<��U���� �6��%�J��[.��Q���{��^p�����$�}�q%/f҃Җ9��\y��Uf�d�S��y�KlM�fuu��*������+Ώ�[R�o�yB���F�Ǔ��E�r~+־�=P�Xij���ddOc�w���F��I�͝�2�^8���Ȭ�:�B�>�DM�#��Z��9��}3W���V4cC�f�S�[}&�X&R}������ѽUo2��.̇S�j��r������M!F~Y�$F�X�	^�d���Og9r���e�˽S��\1,��{�\���ǘ; ���ǏJϔF�_*W����;+�AW��d_>��R�*�ocU]�}
�>7����q~ߔq�n}�S�0a-3��ϦQ��T3���M��y�#X��sTN]p�K���ڸB��	
�V��q2Y,0}E�j����k�D�&~=z��j�թs�6ˁޠsz�i��x�?K�kozŠ�J�al�y��2�3��ysd�={L0g3�]}����ߥ�{{ł�J�f%[��#�7JC���37��A�{��LB�X2�S�֯jbzy�S(wᝥ˿�O/�y�]r5Zo�o�їK�k���[�%����Ib; �"��W2�4���e�S�����v�[ј.�5��ۏ�}��<��ox0�ĀO��ǜ��E�x�={(��
����O��ڊk��{��cs�I���jy�,*�lj���D�Vr�<s���9��{��m@6�/t�?��칣���uƗ���_�����ᨪ�<wWۣϾi{�]ܷ�]\.a�����A)��T���"�3���R����ܕ{A�K�;j5��^����NcE?���e�W�뒓��,���clR�."v
}�L�A�:&zn���#PyUg����d��;R���v��<��ʊk�ajt:f�����6�c��w�\F=U檊��+c��<ݪ2j��*��~2'5ͤ~�b�W܈���y�ܩXҝ��aG���8�%��v���*Ϯf���d]�s�!4RiU"m�V4���)��h��J�֏n���D�8X��6~�*���~�ʿ�}*��T�~�-�e�ַ�sE�Nn�P�<�?<�H���.,$m���f)�*6Q�����>"�t�/[8�67r�{{6����}F)�A��_7���1MP������/�^g��#�g����剚�N`��b�G�,.���Շ9�`��-$J��P���	4on��m"4p��Y�5���o$^d��w*ݽ
����i�K�vO�O�'ݡQ�wW�lY��45c;��˾[l�e9jh�N�4�[�a]m:�o��GX.�=#뽩��F�v&6f��� � ����l��s)M�.��|!M',/ڕ�buL�O�aۧ�3�P;����1�/�V�E��D�6�w
OX����C�IqNiWb�[�o(6��T!�?@����7F��Ռ���z_e��}؎���1u��ja�݄���W'��	u��ܫ\a���'������b�ՠ�r�L@��Wҡ� DG������Ijm:�K�7TQQ��c(-��ݸ�UvdN�0r�o��h�`����O�)��T%O&jT�+w��}��Z������\m՟�*�H˜�{����n�M ����A�䆚]�
~;ʾ�,�z,{O0x�,��ܫO4���'x�]b���<m�=!�$���������\ρ/���H��4�~9�R�^ �=��U�ꭞ�
���]��_�H����{�mO7<a�SԈΟ��x Qk"!��?n1M}*YK�Ϣ�a�~�n�v��ӷp�O ���m8zn��0��X)C��)�ڌ���oT2�RZ%�\z9�ד0��v�I�ð��M������=��W�����{��^���}�л���7yzV�
��9zc�WG �7��w��E8���
�e�N�2�y�]j�Ο:����Vq鵃\�uY�f�Nr�`ە$�R���I5{�a�H�}ډ�tz35=�7
�V(��Y�_2�\9��J�3�t���C+�I:&X�A֞K E[�b�8��JGu��K���Au����r��k��!��N�6rH�P��褱R�w�c7��^f���볭�sz�k��8ճ�����Y��Q�U���\\�����,2U����;��.�'82�����Mvu�[M�n�s���݄Y�I=@E��I��;w�`|�o�T֋nH�Cul馎�̉�n-�N���P-��!ov��.[�9;t�3��p�;W��G+M�ӹ|J�$ �7"� ���$�7s���b�*�+�5JC�'����+k�˾�s�;����
���0S�sB���B1��(�ݬj]����e�Yf�P�Y
�F)��`z�o��ڒ�&�#ڒ�r���#Uv/��ى��m2Bb�58l�Ck�>68�a�M�IdF��L���fº��NYbVI��;f�u�ے��|�(T��7j�A�.��`�XZ��C�erԪ�(�n��Y�N̔�KC5��a��e��M�f�pI-ӂ�v���V�=G3՜eGr'��mVG��ڴ��.kR�I|%�B)�9�@<�W];k�43�w��]ż�s)��I�Ι+i�:^�k]��1]�	!NM�x�d�1���
�fu�4
�O'o��l��
j�/����wipQv:<����͋q�d�v��K6kR�
�h�<�hf[�ݛS1Yz���v���X�E���:վ�pP����I�����ǯW�3hJ�2��x�2��FE����5]ŷ݆����=��j��($��i��<AP�uśR�f;�������k����3\F�TG�l�ʝ���G�]\J�l+w'=���37WH�>�rЈn�;r�CJيd̮΀&�O�����Q܋'U�r
+9������c�2(�K9�s 5є����x+e�ׯ��b��yp`�E����$��_I𭼠m���=�x��#$��$1K:�w�ɱ�0��o\������S�&^f�u	�@���er).�F�-����(A������B7�	G�V��R�҇�U��[�eI����e" ��ڹ8d'V� ���Ig��7�n��އ\��\
�5 9U
Y��5��]�>��)�j�q�g�$��6�:��L�lYnS��F�U�d��P]�P�����v�o�(i�]��OM�Y1ځ�#��ٔ%��QOhL�}�6��
���b��3�X����7���c������٘�eC��y�-� �nGvybU�Z���zS� �O�$�>,Eh>#���F�����a��z:(��j�.�����j�U��n���ZѪJ��k���L}Z�|���ĕ@Uy!���B�S��MPt�z��AD5J�C��۫��)�ݑ�u���$�@���EPU]cT:iu��h��ݩ� �����ճ�g;���� �[4Rkj:��Mt�b�:�#t]�kV���`��U�AZ�5$�50](ևl'Z��QE4ucvuQ ]����a7g#�v�lQh�ԄGqw�T�b(j����
B���[.=]�j6v�(4�4�|�vH�TAic�*�n�C�L�MtRhz:�4芓Z:��"(�ݞ���I]Q�6������^*Jt�	M7a�T��ѧTݴ�1SѤ�Z
?������ﾶ^�V
+ ��^Y�a5;�qAq�\�_I�	L�B�]+ym¦'&/~��}n����$�a
�&O_�ǫ�,����?��@oA�c(#[c���Vi�uй�>�J����d�@)�^gs5�y�����&�P�x�ͬ�	����\�v�	\��0{�0ҷ)��to�?Q40?2�]F[F��d>I!��}t� �o+��l��Pk�)�H	Y�>�B#�#t�2�t
S��n�<���@�C���b���E'7�E6QJ�F~���a�:�?�`KYkd>���`7�'3�N{HT��^�gWk�!a�IOa(���.�}^�V�Z�����W~��c�5ܑ,��M�u�ܫ��=�1�~�-?P�Ɂ���n�I����
R	r�m���y�iD�X=��*X�|�c1��%Gr�)��E�,��öm�+��P��e�1�њg��j�fuo����c�þ�#�HF����ܦT�ޱR'T�9k���X�[\�,3�V�M�e�N���{R��p9�G��RY[�;"#A���"a�yP�<���J�G�C�=@�yL{+}�s-�cY��ml�Az�Y��by��>3�x;k��� ��Dq^E���uW��+�X���ܘ��w?t��Hr0��S��*T��.�@�W��^�^x���Z��=z���k��,_20;���
87�nX�4�X(<�v^�xh{,s��C���nF�Q���c�I��٫S�E�Y\�5���DUt����u���oxo3xr�ݯ�BBn��i�^�zgM�Fu8�o�0�Ο�m:���Vyh� �'&^�������BZϫ=�ϛ$	�������)�V9�99�8��;��<�j�q^1B`�X{�H�D����dS����� �FW�D���C$�>��{_g�"����*�{�v���;w��.��=DDFa��y۬`W.Kȋ1��R��ES�����Elw�+(�噎!7Wx�kަ��O��B#R��Å�<&�Q��Ϯ�S���O��\l)�!_�]}9)=K�8��w �PtC�FG��wZ�=ܶr���J���#Tۻϑ�w�2�s��T	��7�����zl�����N��wTf�H`�о��V����(V�"N�y1
GT"��aɮ8o�uD�Gªjrf��dXq��ĥU�ܫ&4�~��g����cS]or��J�\_v˰��0��v��Vi�,������c�����O���pZ�b�#:��_L$�a)�&����Mn�+��z6ˍii�@���{lw�N��=K�˲<l�a��>�R�ۙ��5~���EX:��EY ��T7lkn?�Aea�y|�|�ǥK|�x�'�\D�X&��ic���ߧ���q%qo^��$���FVT��O*:�Tz�+2e�u�"��y�t��7w��Q��Y��Ӳ���"v>uy'֗Wo����y��D�Ty�Ӣ+���^v�q������o�Z�}�'o���a�CU԰h����o|[���׍_��&/b9���"#a~��{��k���E�S�9O�]��2w:�)s����㚔��'��%/�!�JB��V�
#T�g�	��y<n.&�a�41�_�(��7�U9����pї㖫�`�.h�b��}b�� )]���w�^���Z��u��������mό��B���4����j;�e�������N��`��0���20��5"�sݍQtX�⬂`*�������TS)��-�N+��z�>�h��֛�!R����� �O��/9
N�!���}]\���^��-4���4�6�+W������֘�Y���N5{T�����@o��_~G�^T�מ(���UߵΙ���1��|�.�]��*o�9���9Z�#y�ˌf�URj��PQ,��=���J�."r
{雉�s�h_E�ǳ�C�9�����dY�)ؾ;��<D�$���)�?C�:r�u^����>�R%(˓�����	��ȌV{F��6&}���0v��|�V�:Ԃn�_T��'�6�n��7�:]���s{�����tώ��.-1�Ǡ��� *��j����c�.]o�ڭ�Uأ=�~�Kk��@tB��K��~���|�x����!±<	uh� 8]Fۤ�Rx���҃�#��3���ws�p�D57RN�p,���}Z�E�}�Y��t_�S�^�	�jf��R���"er8��O�5�Q&kW�L�bFl��	ڤ��Vl��btUрSH����Um��b�Ad�-��/��|�-L��e{���;�q���V���8�F�}���r<M����Ė�G!�������ww�8M�۫�U1.R3m��S�'�E�@�y���M�92�h��Ufv�3@�x�a���-1ڶ2��uQ/nbS��Jn�*���us�c!�h�@�hI��Y!L�lZ���*B����f����H��4�5��5���z���\n\AR�ޛ���P7U��s��\�u}�BcoMR���dK��U��&(G<��P|�br;�q����G=�w�	��u�04O��˅A���r��*e�F��o���tl:����q�q�g��-Wݙ��ux)��G�8��!H�yWҧ�5*N���Gs�k��A�ښ�D"P{�E����i���`�z�Q�G�x�L.�4'��,�SZG���S����ZΉ�
>���*���i�|���<=cn8#�T��R�9�����-Q�X@����ûj�x;�z���_W�tl��`!�3��>X�6�鷇Qk �V0��<���eM��㓠�a�(�`1�nA^K�q��d��ӫѰ�*��ݶ;��/~��'�<LO����1>�5-�+�F�4��C��DnyV�>°����^3Vt9���g-/���0;C#Z���ζ��M��V´�y�*���Te��e�$��n	7_uE���5���c3aѝ�!���iۯ���D��Ӈ����M��+g��hQ�99Щk�~%`��}�X=��p��ݻc}�&8y����0ײc
��9��c׮�c��XM����=�G{�	�+`QV��MG�����*k�/��x�.ڦ�f��EX=wI�2�L=��W���"^Ũ�&�6�H`_{���ͺDR�IomA��%�F�$lk�Q���MYη{��Z�����U��֛�s��ȴ蔬��5�D��uq���L���m8c���'v�7#��6�LRr_E'61H����Sqia�aT��6P�Llj��lf��3��h;R�����V��3�z8��?b�/�*V��(�����-U��&��ɓM7�K��]�w�ػLu�Z�ig�"D>3��A��\NΨ(�su�k��&����K���{^3��"�eIj�ڲ�-q�7o,]7��s��^�9�p�I�c�y�S]�ňȴG3�{Z$�Ho]�O�s��]z8�����*�7�>ZX}L��{%!�D�u p��K����J��S���X�g�^l�oR֯��ݡ�yRհ�:��/R��0/��_�������#��}M�N�% %x�gs:)�s�ި~NFI�.����N�����p��9��9cЇ$�ⴌ2���Gr�w�
�<�/�[k:��ߙ����c�9*��~w��m�6��Ii׿$d��1��"��>�ԑ���c�㈘pyA�O�E^y��� �iw븓1x9���u��]�D�a�4���=kg�LW5 v���_��U�1,g���������^m����40��X�^}}\lQ1��rF�5ygH��UZ���/�A/���y�e3&U�]Ƥ���wc�Y����s��;_F����;7�}P�l�.��.�~��,�v]A����R�H�W��� oA�g�֫�������Ϸ6�N�@>$ߩ�˺;�ۦ`�!x�h_t�	{,�g��MJ��*�TEzk�J��T��ঙ럇*D��l72�l��/���ҿ{5;�a8����j~��E:�I��㎇�yfEМ��q�7rXZ����p��|����U/W���=x�A�# �k�I`~���2�ʅ���`Y?m
��69��̷���D�I��R:9�>�]�w���ɫ��d�@��뫗����uc�lw�/��԰`bG}q�Kx-��w��I���+M��_:�lO�����i�!z����;Ks�z*+٠�ǈIcD�ÖՅ�"_�P�����)�xw�t����-��o71L'ˌ�{΄C�Y�|�D�u�Q�y1
@ꅩ��F���e�M*������)��@Q�MW����O.P͝�ކ_+��=����f�k[݌��ɭ3�s�~�ގY�a������3F0I�Ke�+��&�X12��Q�ǻ9�5���֬jݡ�P�O�r5���nu_ڭ!&@W>�+v�;�i�R��:t-��l����ӑzy�sc�eǟ��o
F�m�}9�ˎZ���4�x�ܬ�V�7_�C1�Tƾlg��Aװ���LZ>	Բ��'Ǽ;A5���Er��F���g����-.��s?z*�j�Q\�vH��Te��\���h�LxWU_�@pxx�������� S3�8 z�)�Y�b����
�b~�G�}��߸�0�moT�^)�q�A`��M4=�'��6r��=�cHB�/�D3'P��1�́B)����-�VH�)踡j9�@��c��.h�N&�5��xE92_8��� ��@:�w�);���Ɯ�,控\O�� ��+��z����;�9�3��޼u��ō#�p\��o8�f.�����yy��uf����:U��ZW�QU��A���m�c���X*���F����e/]=��k9Y`�%毼-�em� ʒ֎��r�h3^�@�y�t�`�"�c+yl7���k*+�l53E�R��O{�a�⭿嵬������k��K�;kã"'���*�ZD��O�e����㪙��Lv1U�#u�C
L��Y��U&�7,�tK>���l6
0�s�C�/��Q9�����N�6�B/2`�ݏ4���hq0��E4'�t��"m��b�Yc+Y���K���|DL�Qk"����ݵ5�r�J�"�"�k�H)���ׇY��͜�����zU�D�
$�Vj�_FC�q�3G��d�ѝ�,Ÿ9�y�
ĦhM���s���d��w*J��+6d'�^�L�JS��k�Sm^%KI��<�L���7���:��mw��6P9��X����Sw�/LB�X���b��2!{��^Rh�[@�,/$S$S�tM�v��\�S)��UL���ۖT��� U��<��\��&/�w���t8\�y.ԶΞ����Cr(Ч��0�9`L�m�
�n�Rq�ę�|j.-�CD[5H���P���n�m�h��<��;0���Qq@�*���f��g��t����nB�����
.)����ff�$��aOwWn.wa�'���I�4a�>�0/$=�۳�2� �Η����������Z�Q��fK��U�{7��MN���eq�:����X��j���ӵ�*t]z��Vʎ��m.�6����zm��v~5F����=�"!:j��ms@dK)8�[��%�D�*������	��U#G���m��O�p�I���j�%G""ޘ���ܧ~��ɹ�����2�Tᔘ�s5,{r�9wC����l�WH�;�(.;ʥN�k�Rtȍޫ&��ay.���e�ӥ�v�Q|J=ʺ�H}ጏJ�8y�ZyQ�W�^1���lN�]B�c�N��������F�x}ý����}Y�Oa�=iJ6�6�^"���;E	�M�wf�����bEF���lu!i�������.��q�D���,3�����Ԙ dڮ�]�6���_J�����x����NW����w�n,�7�D��c�x�+|۾�Vr~�kS�,8��|���I�NF1̏snfUCW��v�J�3R�>}T�s])�d�/]�
sm�
�\��KB����0���?tu
�:�������R�iSR�^���Y�j3��P9�����-DO*J��@1K��]d
7 L_Ǽ��{��0����:�)Ϭ����{"i��׍s[�����Ǡйl]�d�~�}�|������q��BdFQ�6Uͳ�Kv����G'
��d!��"��/.��Hn"ek�sܻ6����9i�,��˫l]v�(��l;��CP��>V%�;�[�H��_�.�ɛ�?�7�n/�gG�fڂ�hm�������9
�h萕��}r1
F�8�����Jq�H��<f�du��b����~O�Rr����ި��y���)8\��tLL�ܫ��or?{�+��쓵Y(4������)X�5)��o�Ek���Xln�g��~H���n+�=r72�ٱ�]����"=��q��ۻ�,�\���9���iO���ݴ�ےm���F	���"��t��o�n�����#�|%C�R���?m�g��u'^t%���=���nv�(�:O�Ǯ_�ǯ�09%id'�=_J��R�?��xW=A]�8gT;3)�\�L���%}O�*j{�FM:�s>�N!6��ԑ�㈘�w���q��;6�YW��=um#���S�<�q�v	T�m��h/B�Ϟ�x��j��|g�ut��&0s%Zؕ2jq�[����_m�W��ΊǢ�Ɓ�1��XK�fy���3:���[Uc�Z�V2�����A��H�����8�>��g�v���rGqx�w�8�a��F{}ޟO������<�|}>>>�>[F��7��5̌�y�v
�R����ojg~v���
o%G��P0-ͷ��*���C6��O��5y�,7>���ڎS�n�F�B/s�6�L���+��_��7{إD���Gq�u��[�����S
}kO5\��d��`0�S�Ƣ�G$�Q���u����)k6�(	JH��Ƿ�kH�$3�k|*#W�[c�\�w �@�dvSԧB����-Gq�N�Gj�����D��o�� �o����c]�n+@7; 	
���Nc����Y(^n�3�5���!�5�n��Z����S ���B+�^< ZSܽ��\[#��5�����sY$�<h�LQ�s��ί�,g�󃎁����֩��)˴�v'5���|�Ow�~�:s�����L�i�p��y�[B���[�t�=�%�w1�A-xs�L:ت��q�����p���5��W3y��f�K6�ܚ)p��.^�4,=8�}8''f�e�(n�*<�����Z'�>9̛7�
��]�j�W	w��͆\��tEIW�h#�2ļaj�h�E|�+8�mF�%k��3�A:흒��CDX��d�X**�٫�C��P9��*�K��J�Ӊ�bQ��.K�}OsI<tx\1-O.�J���pwpV�c�+�Y	��9��5��Mӕ���,��$�]�H�B�᪋������[�(4�7�wEX+��w�5�#àJ���C�=�S��&��l�qn��r��X╨���r�<j�sw3�%�н��Ews��V�R_m��Y%��S]]i�[��b�k��\�,f��A�5���̝d�������N�R�t���iPudʀ��g7*�d�B��[�ҝ��-�=�����ә���Cgz�I�Q��^5T9�a�.�2�$�v�7YL�!{�\7�^��M�K�h�'.ΧH��f��s\.h�4���ò��p�� �<Nb�4#�u�uhk��Y���n��W�3Uw7��D��[��u�&��s�r.Mb�+��c�ub�X2�r��sF�w�VFg�Q�����R��w�4v��Vs�1#.�Ǹ��
�4p�OygT�CGuc�z��36���5{�w�89R9�9V���;G
�C
@u&��ѝ�vm��rK��q�gj@��BS��q�6J�S�iu��(g%Xʍ�ϳU_��eA}OHᗰ̧~�x����-�)�/5�h*��b%�C���&Ph���Ƈ-������ҙ���+�駡T';%�sv�e�Ǵʿ�����B4��e�����G%٦������_̛y�;�hX�QTb����	Gf���&*/�	u�[����^!5���g�Ӽ�.��À���<E����K[&���D�K��}rDI8gQ��p�!i�9�l�E�����[2.�an�/�B)��"H�VG�f��2\�ѫ*5C���7�d�n���轥�l�ȀB�w��]5sA)���$H��E��IQ4�`��E&�v:�N�!ZJq1�=���O<�!���ӣ֗T�COF)��)�E�:률�E��Ռ��ѡ�
��1%TI���F�l&�I��K]:@�n���h8�4��i����݃CLMt�R�h�]����R4�4��)��P:H��4>��5֬b�u�4����.����F���l�Q�n�]d�MRPI�h&��N�t4�����G]4WX�����M&����AI�"��#'T�7ZB�ր����&�*	��)i:1!�tM�CmSMh��qֶ�)�]�4xZ����-7a讝�ttJ[�iu]%t�K��M'DEih^���i9��[�m�L�t�5�?׻�z�ՏT@�"�Tܜu7�fD׷v�c�0%�z�(Wk6�(�Μ�*�b2�u��&��ә�6��8��)�Uq�6Ԡ��[�m:H�T��#��Q^�}~��H� X��n�5��t?�s��~5��*K�	����m3kݟA#X�k�!&����[9�ug:H"�K�f��u�j"��,�����tsΓ���N�V;�u�>矒�ϴV�l�n�G|�Jˉ����dy�"�s���|u�S�H����Vg@�}�5|�zo�v�0�4��u�-,B���@�y�m$����{@���غ�z1,�gw�R�>��@�*6�o�m�{L-z��C֝�/�����KYY3d����SMb��Ɯ���+m}!tJU�^kn��O"�So���=�QI�������
NuA��ɭ�i�o�{ix���~����_J�(M�n���[� ��>��L�����:�t��M�eg�̿����z����q��{��-�aR��%�e�2A���P=ԭ,��/���~޽�o�hT1vw%��8���t�F�m�3�1@s��U�QQe��{V����Í��4/zw����4�y�:
󬰳0���:�Z���8��;Cv\�D�l\)#��ٽu��*��R��V����IB�fF����gKZu)pw���kR��tǼH���뼓z�kFV���0��J,�
l��ߐ�3�2VnS4����9A����(ٮ��ܜ垮6��M�-W���&���w2����{([�r���eu�7ʰ�[oXk�j����������O@c�<�by^�4e�����
0Y_TH�y;0t? ��Au�t���L
���C='� ���ds]N�e?5��7�t_q�w�*�8ս0\ڎ�a),!�~G��!�=�]N=|��-�XH9�6$!� �<y�C�s^��R#��{��C;�I��Ȝ£{޵��c�������m�W�`�*� ��(Q�@CS!����}]J��N������8%����%Ɨ����NL���'�)Mu�#|]"4�G�E{DayiO�+ ;�/x����m�`�R�kR�����0���>*�576���Ǵ���^�+�a>���[x��}p��rj�9X�u�Ƀ;��.W�$7Y�$6��r�hO]0��u��tB��77wb��ǈF��Y��f��>5ufԴ4��<��ƞ�[(7X5"r��$�w���듕Y���c5���a�H�@��V7����U���§����8o�!��r�s;mo�Òjzu���H-��]���iC�)�������ߔ�W��S=��
�ɯ��U��t��sg�C�\A	�^�{��d�hJ�m�a�	��p=,
U������8ׅ��I�a,�>6�)�@&�2��U������[�WOx%���&F���;�b��v����K��PōI��Ț��d�$�k�8=$�~^�X��6>�
�n�;X�� ���0�|y���RY�R�faw����xH���}ֻkQʺ��D�w�6��S$�<�m��M��7�����(%�7ןT"��	�i7xtFT�p�W�f�0� ������%:aiT�����A�&b����s�nF�3�UV��to.us �p�e���	�tć��QqF)Wb���z�󗋋��������{�Ɩ,��s�|��P+��%�D!���M��*���"�\�����3XBZgqL�EF���+<X�<���~+ڟ��^#>ٙ�=yuGk�ѡ��ъ�A���|%�i4����;.;Ǡ���!AiM�;_z>�O��wHA���*y3R��K7������Ӊ�n[�����E��;J&�Z��K��a�s�aw�!��Nެݞ�'ݺԴl�f�1�\���9��E��ϻ�Y1"6��q�hr���\��J<��1$�pk�3��`���(HQ��*�),K�.����o���ג~#�P"���x�O�X&W��*��t�`
���:E�g�tr&�!�#�
�]��$u�뭷B緵;�.�GZ~~�[O����z���\��C.im=���}�v��5�8f�,�y�`��0����n��i�bTys�=p)�ַ��[�O�1�C�]�/�>����"@@ڳ�n9�	q�E	�f�]�1�v��f88-��< �]��~��w��:�y7Q���: #%a�������,e���^7�Ȍ��]���ymMD�-��-G�<rH��ڐ�P��ȸPЎW�YZ0��i���T����Vs�i�o3У����;��O��n{&6:U K^+�`��)pdߎ#�G�U*bw=/��z�;��*����!t΍@23vh���dg�q%���;m�i�.�T�-�H�e*Ç�D�Z��[��u�%���6�M���:$��k��)9��B�mEٟ|�r>o+���~E���(�>��X�|��%f��(�.;=<A��wމt�g�ŵ�����*չ�W*!�1�~��E�/�y9)v��8�">�L}ȵ�*8���x�"���Y��v���d��dd��6��P�U��?*x��X�t ϺaK��t��~����(�L_6��oy�M�:�l�ީd5\��(�#��@���wx�>�ƕ�0\��P3+���$��b�U�ۘ���\�x�ҍ+^y�DR�z���A�߫�^�!��yYC/�ܼZh��K�0�����ݹ���]jV��>�_]�
��c��e>]�����0���q��r�V���j�_�{�������'f*5��/ԺcP�;_�7��0w��:�hxTS�I��l��6?�9"�
8d˜�M)���r�����,lD��������=�'b��QU�mЗ�~/t��1�h]�U&kg�е�O����sw�gm~�Fb-47AǦ�����C�Y�҆"֟��SJsӦ�_�:�ny(41�t�
�����:�G1��u�v\%ջևvl���ݥ��jc�����������Q���MV.󚕎�sn3s�\6ȴ��5+T��eqd�ЪQ�Q	j�0Ht�P}N��=�^Wm���4�"2)s�M����\�P׌�z �f��T&��hj�)K|P�G=4K�"bb�5�֕W:n�U(����沇���t���a	p�j�1L��"���']q B�S�U)!�ߐ��'���9�3܁��SU8+׆jZ�{1��6�2%�TS��҃#�/e�};�A���K�{��^��S"�#(���B��ʛaC�-{~�+��w���<���XE�҃>�\�l��_�pW�:��6/��3�d��`�y��n�GD���	�>'���ۥG��eO/ �y�J�P�u�M�Ck%]ǱV�������D��p�~�e2��ۡ0��5Ήc�;�(2����P �N��� s�J8�Z���{V��m��Д��+l�U�پ���v����ku�C�k��<���_Eກ#EWW��t��j�C/���~��v��x=7�M��C���,_�G��~���x�<_{���u��ީ|���(V:YyCoܲ�^����C��¥��	r�d'1^�m����]��U۝V�/�s�G��������zJ��v�Wf~>� �A	�yҲ	��|��vM��҃��y�3bC��S	&�7�5)��tO7RR����D�9?~Ϥ�<t���_��-�8M��y����a�.(��,�1<����Sߨ��ه�����4���\(vu�ql����*b��0����������C��������.@�k��MI��ޝ�LG($>�R�� �@� � �N7�Bֽ�\��_���Z��eѹ{r���;�"y��t\%ѥ[�����^� � �P$F�蠨�&��f�i�:�18�hLJ��ulὩ�{�_8�{j|F��^�&��)��\��t��>�?=y�ʬ����d%i�ԙ��30�;Nz��XG��繝h�܃Һ��~*��0��f��JO:$�^ݏ�}�fg�<JͶTmz���E����0K)�.�2��t^uY�9a-]�Mh�5��������Z�Psixzs՛�ʽPflf�a����Ѳ���,�yx��B,���	����rK��J�}�j���ٌ��K�����p�ʋD\���Ό�Q�b�b��5g�v�>K�6g���`���#�ޛ`ܢZ�n�h��ӳ$U�C䮎����z"[d6Aa"�SQg"�>7f��K`{�,[����E�NN�B����^m�[X� ����"��FB�X�+�����m��F���} ќD&�FV��X�4��phB�Yt&�u�O~܅���6,:=�E.2T�Mx��r�z�-աx�7���.�Gw���K^�sE�ٳ�h�v1�D+8��+�Jif�%s~���(�X��g�������u�$�%�2��s%��|�l�<��)���(^Bu�?}x=�	�wUe��e�]��=Y�Vt1��L�{�%�.��m�fm��,�P�q�*��̬U�m��9���89n�	���} �\X1J�vO-a�8�N8�Q��#.�1�e�/.B�p+h���" �΀c��ۻ4}^��;	�C����gAY*�/����=�%����z�U٥YA=C�%G1���*d��:���A������m�!��F��a��{	��i��lu�;�T��w�i��_�^�9��j����Z�>ŷ�,-��f�[�]u0vx�i&��s���n'"��ځ��]��q�cr>]z�S����{���F�fܕy���X�������̥��[=�Z�t#��+��^5t�̌�量� ��(�b�6�,��ʀ�eV�G���˼c/��e�dl�v��?:�c+Z��*�Q��}���_d����N��G�����։G�!9o��6��ׇ���ԁ/1A8��z��5�tt�|�g݌�,��񩯻����KN�7RF��]����v���ǈ�V�
�эV�M��^�
��FQ3ĺ��W�y������8��(��{�{ADxtB=���p��d��T[3Y��=�[�a�6�c��sS~;ݬ���_w��X�רgΊ�/���~_=Oq��a�Ԃ$��f(C�R�	n��g6l��@�l�4�|:[�/�P��jo�K�V��R&���jk���ޕ@_��A$6J���e�n|���7j����io�旞e�-����eM)�'�.k�����P*�����*�sر(�u�}3enӧ��p�游��l��S���Zh?A���Gl�z���
̬-Rmt��s���`�+���3d_�s��1�3ܺ�K�n��i��k��z�	K����f�}y�4��!}��r�K��RV0��m�Y}/��Z'1�yL�FSn��friO�龏���*�~�Y�6��oΞ6��f7A��pr�{l{�~{�p�g@��;*�M>����n����Wy��6;4����zQҥ��9zp �X���|��,��G$��Pg�S\�!l�	�汩sT�fD�
ϖ$���%ޱu����t ��Tjhuty�˲���7
�(�l��&��\f��NAvï=Gxr����o�A�h�l�����?q��8ӭ��՛L���ж���3퍛�v9щ2�I;�,?+B[.�|�Ϟ�z��Z�o����i�HE�;��= >��t"��2��ǧ�km!��!�Q�j��&-vW�H~�ibL��.Ӱ���<�,��gl$��3�pU;	���6g;̠d3��qyF���6p��]>bo5��n�3'�w���%�7w��[�� �-u'�s=�|�N�}�Sb��c�V�����������[��ݯ�t�E���r��V�zL��Z,���ܝ�/��T�i��k�܊F��\���l\W9Z�*�M�Gf�Ӻ,�S� �W�g�r��\�Dnz����Kɛ�8wƽ��h�����4C��*ۛ[��#�i�3z �t�7	c7�։r�KC7��x�SE�Q;i���ov��}�/	�ru��ix��32_u�!��B�xLڥՍM��c6k͈%K�3��f�Gv���r}j�^)���r#$�r�[22ΔC]sl�:H��Y�9�<C��ך�\�OTTN�K79�)H+�NV�p�׾��aލM\Q�-jW�[�m"��WK��HdU�v�W�R�Ff2'�%����~���7#��^�ƍm�^�=��'А�C�~~�V?`����q��,�ޔ;u�>��ICg!Uvr���K[�)�}-��A���yA6Lg;��{���Ǽ�7��[��t�7� �����g�zW5S�s�|���T��}��i�o�&W�[�cvC����dȓ�ԡ4�T����UBg>۱7�~�wQݨ�g7����@���v��P�خ�V�Ꝉ-��g��z����	=���U�R��,���?�����=^�O����������o`J����Q�w@�$+6�l��0���W�:P@��0��Sh��I��Qy�q�\/�� ����'4dt��
��/�s�ge:��T��sg%C`uo�+���"n�6�Q��,s�W�[p#]����q��)�iQ��l3��{�
U�l��l�V]���#��aߴ����4uϒ�]-��8���:�^��6�<��яe
�%K ��.��nU⛸�(ź�'^^�����1h�ك��K-��/�K&JYvkaSP��I�l���sWloz��F�WH5��4��U�� e��ϴ�>�}LlxD���n\����RC��u`�2�W!b%tV�rN�s�/{6	V�:Cq�Ox��}y0��<�P������Cs���mC��V����b���7��.��DK�9��Y#���c�G�1:��ӏ:cy�K7]	5�m�n�P�X4��M��ct��1�䥣K�[&��v���&W,�����	�@n]5@`I�)Cz�O#�re�$�T�1����C.��
lw�LzB���1����{}���_^�r����I����i�^��z&H�J��EcF��UŪ�W��:�Ӡ�TJ�i\Y����rl���W#�(�5� �++/F��CN�3J�+a�u�S�\.��4��a.
*�d*X�ݧB��<.��㣢@޹N� �D+Pl^Q�:�gS��O1�հ����%/�H�CG��4��ĳ�9Kc��ʑ�v�/�Ot�YWH��s��	zn�1a�0v_�ksf��a]�;:�2��Khln ({f�K�7v�It�sm�� ���JɿdݧY4����d0�X74
j��bf'�X�K�)f�C܈^0��پ������M�!���<x�Xc��z��
�f���(�n�b�fZ���X���(�{T��Ej��^Ձ\D�)�%Y3��wQp�[LS9T�3s�i�� �>�x35�	�y.�{��|b���gpə�QX����͙�"�u���|�qB�����7���K[�p��-���N��	�kol`��w�u΃��!�����&�w˄1�so �ෘ!�����1�GS��3���nq�B��C���:&��us{�&'�Y�e��h��n��;�C�vk����gX���]`Y��Bz-������5��"q�kz�c(i�GV�.H��^8�82�V8mr��麺F*jWSnl(� ��=�5|��=�$���w��3��w!���-)w����s��5�/v���&���tX��=��e�ד&��t���x�d6�\�X�ݕn���r��`SS�S�@.�X.0����+�����EKӘU�d�%V��!)�.)/+w��J��W� 	8�d[�V��1vͲ�**�/%=���I���2����o�t���O)f`-ne��bm�ٚ��.�G�gQ�����e��]t�Y��K��zU6GK��v�}αC3J�OM`�K�w<���h{R��-�hC7T���� �0L-wm�ӫwb�տrd��ر`��'3���=���!�*���b��h4�lP��E6�s4j��tQvѶb�Z�KZLl���@U��U�t���"��u���j�u3��V ��t�b5�u�h*��Z����Q�t��\Z���:t�(44pF��&٧TD�th;]�;]�'U�S��M&����Ȯ�m�lcRk�=��uZ�N�b��4]wU%���m:h
v�j�"��o^nj��t�h��{��Wb�Gl�0�QӣF��ݕ�`(*����ѡ::�i���GAQ�QAI��
+�����4th�	��w��gAU�������=V٠��5�h:�ݧ�ՌmcLƍ%�kj1��UѠ�5LԚcnݻF��c���:	�ۻMk�����k�mKѢ���B*(���W�~�	�b�\���1�t�g��m��)�ͭ ���U��ꁁJ�f��j����j�r�q�녴oWD;?m^������hl_5�3����0����7����󾣞�PsI�9T��ߤڒsv���k4LQ�V�{�Lŕ[� ׏�Íp�XbWo��d��<xl���Ŋ֫N8�V�2NK�VNSH����&�=�-��hd^�o$K���[��4��d뉴�)�ؾ�:ݞk-t�R�4H�l3ølE� �4���蹾ѐ	��@�nbs��hح�}��_.�-�,k�nk�Uݭ2	�,�S;�`��
�y!FA�r#Q~���1q�SY�ĔB�v�w5��M�gB�:F�4��f�+�lS猆*��f��m\ٯj�8�SL?f�Ԇ|:�>OV�q��S�Y��kG�r�[L����f��q��R�S]V��M9M67h�f�(��Ex'�J	P�'h��U�V,w��[ 5ٹ���Y~�ώ~�}ރ�~'�2W��Gݞ����)A¼��A��B�,���u���6s:��3ȍ�4Y�æ������%�R�}EF�|L�.�a�ܩ��7�@���yNhdi·�
% ��Y�I�Nr��e  &���̙^gh��;��0)��:4��Zn	Öj��1��Sh��᧕2:�{��g��c'X5ڱt��J��4R�o������y�[dG�M{q�y������J���4R���SGr��'C�}l����u3E���^|M��!l�(�.�WC�<�N(���b��bA�#��ɾ���4g[��L� ��pc�9�&W�����}ߟb�)*�R8�ŝ���&�9{�{o臽S�2R�qXꑏ"ի��ތ��6{���\0���4�_�6��?gC��w	F��d�5;q���'�ҙ����qŶ�ܛORL��kc'���l����L��T�;���P���������V��k,ݍ^�ͦ3Ӽl=]��A\m�MF�L��<��fԼ�tA�6,��[-݇�Qn;b����=�9~�7����r�r�����B�0p�0�}�#��jh���Ί��!�o���l%Ԛ|b�H�lR�G���Bt�l�ٞq뉮t*;�����m��AMC�E�]�gs��4�U��n��N��?_��M��7u͝훒m�=�zTk/FZ̺IoIS�d���U-���ccc��x�����&�	�'n��e������vN��!Y�M#:�ڱ��x�촖tuJC�Q����J���r����j��e� s~��u�$����F�f�i��c>tV!~�_||�}c�ǐL�%�%�f2ot�er	�!x
����l��T�~��˞���p��s*����]	;O
��W�P*�J�J�+�-۱��SdO	sm�c1���F��W~~���e�r0�Gl������h�����	z̽�e�����=͞�z��,�i����f�8�Zh?$h�%�^�'5������KO���ίo�?���}wk)�!�k�!l���oSЀQ������ٗ�s�Cx�en�ڨ�o ҉=}>g� C��Ama��6$[4÷a�9m�>����}�#��b��6���}P[����H`j�=�����kީ�b4����*o���\�T�q��[rF�:^,��{�s�ǽ��+zZ��[ Dq1a�MV�+mo9�[�u�g�ykmd�Si�\"�3"��gm��wS���VqڳJVk����C$�b�/b�G+C)��:i�nK�\O{�q�WG���}նvo|�����V�(5��,G�@�R�*�e�]��jܫ��o{��Q�����K����Z9�ʃ���Z�3+{oy���/_�C�vE��3�=��W>��n�tN�}yn�B2�rqLj:���������]����b3�Y�8{T8(A~���Rj�GY���#'�l�ڶ`ўy�6�8d�#o��RuL˘�~vӦ7H�DaQk���� �Ô��W
�Ci�<h���"r�c���G����wߨ���*��r��9�&����,F�%��5ǶӺ�}0�)
�g�X��cFd�E���U@]�#7&$_r9p���j�l������5��eo���ߙ>��1P�U��󇕣�Yi-��-�Rq��_���!�ڍ�w3��Q�j�ٽ��6hĊ�pk����EG��8�v������)�n�����²��XOuYz�� 9l�^22�p4�d�
l�"������f{�UvV������c�s�zJD���WW�9^D��c�3]�xz7�}a�9Xs>��D���WU�M�khV!��(��"�,�#X���hV�L"�k��'���<��Q�Iou�eu�V�����C'  �yٌ�"u�8�d]���g`��	�r���V�4��s&)]/R���U����K|ٚ�ӓ;�� ~�sG)���<|!���ܑ�0���N��޵W� ��7����7�2�p�V^�lew�F�(.:˴�J��U������(�@XU���O�+]��x}݈��&�=6I�X#v>	q���֞d=:�j�YD�{�u���.���tg3��qm�\��f	��zb4$���JQ����������4�{"���Ya"���ϳ[���!�ڏL�m�QO�P���
K�[������Z� ���9duq��\7������`ݿI�K�R��_��]�߻x���ĶH�&y�?H��d8��&�0��,�nj��#'�%ϢׯjBۑb�n-�~:�`���
�X�d(��Z�����Փm���Cg<��ק!eut��T��pW���u;�3��{{2T&E[�v�g��Wt�	Sf���]�s䟼M}�뷒"M��j�����9��ƋIb-��d/�C��l��J*���l���X���yr-�ж��N�Y��o�K(���Nr�V����렐�u7��I��^���]wY<����Ɓ���7��$���2�+)���xZ����tjq� 2��n;�|*��)�UT�_<��Q�/�ve�r5-��ɡ���g�j7�:��}}��XZ�%aʷB���r��,�g�u׉@�(9\mmyT1`��Uȟ�|�D��=<�o	~�C�\S���n���@{��}	ex%),��5���|��+MwS�r�E����7q��oCJ��h���Ժ�t��*]�
�Ł�w�z �=�����qʥ3��0�<�׻�7����g&7|���͌v�����Kj	,����vܻ٘u�p�c^I�Z�]��d����ǩȒG����,���o�ض�,3�}�y�Y�Rڎ�����1'{fGfoM}m�<���-fMγ�!h@����ˍ�zB�}��tMuZS��3�oz�qW �?H"����������<α��D}L�����F�^�V��JAP8�}����>�s���i/� ��
86*1]CG��]0Qч�O}�5Z�`^�V�<��]Z��E���VS���#�	��W����Q��DF��*�IϷ32㽷j�FI$��u�^2���OF\B�4=T�j�����tA*�@�l�7r���7/$F��l���_�k�{�1�F���WM���=6�^����;qٍ%�Â���_��sײ�Yw�=~�9�2���z9@H^���z��YԌ�-�t�9^��/�f��dT��{�"*����ۭ�bϛ�;s��';�/���W>��2�n\�=My/��;��!����! �2t��
�hF�Oc2��
���kX��iȃ�x��<U�ٔ(ِ3L���m��8�r^|���7�1�5*5Uw�Ixȓϱ����;-p�Į�aK
�*���Z��W9Ed�\�nO��'"4p:<��LvZ��O2v�<�f���U@��2w��]���w�N���s�g(Di��� :��ej�ʶZi��SG���,���%�Z���h�oU|�p�]g^q;��r�h��Wq�v�e�N�>!l
���W��A�� ��V�.�5��_[�֕Վ��nRt��<.�7�oW6.֡�jV�j�c�O�e;��
S��1�H�)��W���`k��y�Q����d��������棝Su([7�hL(c������/�&�]���!�G�B㹟v�z#Sbf�5s�j���9$�������#hĀ��C>C��T�O�g�݄ڛ�7�tZ%�U�5���	r�-�V���Cdړ���'o3���K|��1��3��j~\[��a1&�$���w�B��6ɼ��{�u�Y�����P�Ȉ(О��5������V�o�F:��y�O�Qk��L��G����`v��b�}�ײTtq�֬q���MA�GD�+�s쩝��ߤw����l�t��m��^;ޭ������|w~��FԴ�~F�&�4<,�CmGї��8WD��^�R���֚�������[�:\���X��o�ڙAٓ�?�����&/K�C��z�Oʊ���1E{y7O�AO!b
��]�l�Ȭ��mǊ9�9>τ��b���Nu�]�∱XK�"2O)���k&;NC��W�b���в�h���+�3�3��W��I��ȴ�.���6�H{-+;��v��t}]B���]>3ܩ�t׃��S��y
���L��'�`+:L]g#f�T�۬S�j$�Ԭ�ĺ[YC�^�=�r��U-�N>Es�-��st�n��ܐe`r7a��ӻ�W���׬����W��H��SX�6߈N0���l���l�IR��������t��d�@�J�!���S�P�T⼲��i����3q���;f��𩩰s���M�m<�g+�j[��L����is��^|�ous��%���)U򧫫c2�݃y�.m���kM⨶38ý�cދn�7$x1���Wwg������'2-����{�1m�x�3��=
���z@��va��&V��ؽ�u=�c����X�PՖ^�=�Ԡ�5����dE���0:-D���=+��ʴ�Pppro,�YJ�cy� �x�w�=�����~���"����m������7Gń��-��f���i�-���O�D9�z�3����k�K�[��z�R�z2F��44�����}�I�Ĵ��5u]ZN,��t�E�0�vl�2����n*:���E����P{2`��:7�P�*��B�2h�,��k�~�o���`�*Ph#��R�k�ФqJ��NT�6�ܳeGۊ������kkp�e�PJ��?6��}[7�v�헾T��d5�7���r�Gl�A��!�Kin������5@04��=�"Z�L�۱��z�_8�����+����[6�eŮ���e�ő/ pQ8^������Ÿ�]c ���B����:��.��5��o�oG�q�6!��?{�|T�s�����x8�<�ԉ���2� qk�T� �2�l9�L�5�=��E"�.�>6t��{9�
��ģ����u\��&�!]�s��,�W���fw�(�,�3�q�#�Wr-A�4��j�q��Y��'�w��I9�Y@�޿I���#�Y�h�����}�$�U���ҿdd{��ɮ�En?�V{w�sk�n&{�}��6��B+k1�^=�p�<��R�h����9��M�!f��\\�5ǩ��+�g�SC�YZ�ns�w$g�]����>�W����y{���>>>j�a]W\�Be�zn`+⺲�n���krP�e�f�$�nq�d[`����f�N�k@�.bU�s��5�_<���Z\�+l�ͪ[����,�|�43�� W]�cH1ʷ��kU$�e�w|H�18+v��N�tr��7)5-�Y�x��P��N_X�b�KU�'o"�[3�T{�\�����CN����1����f���7����y�m��ѵq)۠�>�̣z�wi��GC9��'�ɍ�m��*K�pb.�C��wfvڸ88'��
�<�mz�ZO����̳8.�u�X�z�4�Ш�K��eۛ,Nj�^h�f�;]v�$�b�6`V?���.<�[c��u�uqeh�i>��Rvj^�.=��e�q*I��%*��PD�)�TU���k1��&q5����"-U�uhƸ;��*𙕝(N�͕���֍E��*�(3.[�n.�[L��;`�6�o3�3�Ѻ۝����إ`;j;�t.�KtS<��Y�0��(I	��愻�,� ���L��5�jmY��u8��M�Y�V���H��q)G,^IA�7pDr�*�8^cA��o���X�Ԯ�9y�VN� V7��~��R�q%�1��̜�"�L*��;�+Q�J��`;�T��>k:qoYw5���6��L^�.vt]�J;$z��f����3i٬QP�6]����=��H}C�(�Ȏ���%v���o� ��:������p;�z0��tٻ�f��e�Wu�2qɱk�lUޞ|�(��y�pB�uN���r�$Q7��Je�܁�G*]n�nՍ#,`��~�/]�b���8.7Rwvҳ(��K�[�7)�-�ջQ6B��{w	��M�6z�4ee��VV�"�=�޷������T��u��"�mp
�S�t�Ed3]ҏUð��邢���=��(�ا*�I�+^F����o�$����Yj,M�-��:��oVJ�m�N�rF�/��>#/��H�N>��;Bs�������3�;!%E`cXlq8�vV�,�K=]��s�XR9tՑnŌ��{-��-B�ב3�ɅԌ�"0�7+QDm� r�n�0�H�&b�2ؠ�^����
����J������e����i�iK�M������j<�[
�Z7�����I��Y(��4ID����v@�Ga {w�mWs��J�\����vjLT��6��RY��qV_Q�p��mf�iuD�͆�gS�5��w"_FZ��*ora䔻��u�f���ܩ�ݨ�����4]YR[kOi|��#y2�7JB��!�P��E�y,wWS��	�����'�x�Ů	K����쉰��͐�p�] )C�H���Ύ뇣w��2�h� �0�n�s�gi.YJM�m�`�%C2��Ev�6�J�̘<��|	���H /�(�F� k�o<��"�4;�ֻ�h5F��I���Hh(6��4�s��F��6�u�Pv7kj�4��uգq%wX��1�Mu���ӭ7`蠮�/OWn�J�wq��Llh60b�퉦��V+:hz�N�qh���b"��\[lci��`��b���F؈⠱���㱶)�֊
]��v튍h���mp]ڠ�렪9�%ݮ[ը�;���hv���뢃�Ύ'ͩN���"��n�kv�ֱm�����홚z:;�q���y��6�BZw��݃�J
(�Wv���cm]�wwEq&-P�]��n�����u:���w��m4��.�I�h��cn��'n����ۊ"�N�gZ*�jtmDi)z1�������զ͎�v������{����m����������춳w�(���B���6cS���ʆ>θp����@�>���7-V�N��Ҡn1�i��ۢzY���-T�t�UĻ�K.�`6I Y�l�%4�)4�P�R����ˈ�,B� ����s2�_��V{�AK:�"�[�d3٘u���w
�|�:_�1t��Ij.�
�,��?fO�����6�X]���H�@�[�ѧu}W����v�D�����Zk�fM��sehK<�_�;�
ʎ�Y��*��Ϣ}'U�Ƕns{=��d�z�@V^�=���=(y��^y꾝mF�Ҭ�o��?g��� ��G_�?[~R�����{ш�~�ҿڌ�g"�YS�DT$5X~����;���@Xd$���<$�;����懕N�%�҂���x��N�gHp}�3�WLr*������ݍ@�v�`7���4��ι�3ۇ4�͟�1��^T��r� ��󗑀�Ny�M����}��p|7�5��fn�P�M ��'�[22��G��Ƙi�|`u^gVL�m�MR�E�x��]�S�������=�V��ϟ�`j�Sv����>RoO����Z^s�>��坩�^y}��_�̯L���(�E@��%SS����`��xNA�r�&V/I��IĝwE���tݰ�S��-1^��L�F�x�i�ƫ�gtܭ��d��iPů�:�w��c��y{z�*��<_��zUu/�SFnF��>�U��j����s+�`�<'6+qg?1q=�r97p��2��n���MZ޷�WE��9"��n�wzɲg=�G���VeP0��2�H:e����U{�����A���b��f�EB���^g=�I�^9Y4imY� �Ԁِ�5Ȃ�=Qn�t]D�=miu+��ٞ�t�9{�a�J�e����Uՙ�
����\]�A���j�^΍x`Szר�����5��O�L\m�H��]��u�q��H�16mwު�6�L:N��6�U^�&$���<C��ȹL��^!�I�y�Q�3�cZ1�Ľ��+������+Ճ����r5�Z!��_�83g�|fn���U�-km�w����;h�1]b;��J�㺯�r؛[\�2v��s������v��[!��������#Q�`e�w���D��n{�-�#�=ᐪ$���^r��nb/խ;��1�@�j������e3y��]��ܖ�v䮼 q� ��hj�p]-��/���4���B$ �ՍP��Imk�]^�K��YX��zN�|��u�"NR�U�D��t)�07'e�PԬ�xo{����Tz�oi�h��煖>l�R��n)Q靆O߇�������d������ϸZ�6���:�I�I���zh��R�:��xh�ӯ�*DM�P�� ]��7x�P)!�f�x���Dvm�MՊ��ޖ��Z�q<h�^{*bk���da���%�/fK����gg~�p�ו[4�1�m��A�W�2�j�s�vU�LM�;�X�#�d驼4�F,w�m#�h~����g�g;��YOM�W����P���
����op����><| ���Oi����
,�Yz�?A���JD�K���t��U�5m'���h�*cr�;|o���wf���M����=3��)��Qy�,�J��	]ϴ��&���@�G�b�}�Z~����il�oyޤP�.���ە��b�E����t��~-ᴠ���ʰg7]�:�7	X����#{\4G.����k��JtN���4����e�]w2�m�2:�e�ݝȴ�`��F�f�}�ԓ)�M���6���+�8��Y�!V�z���1~�i�������wS>�\w`�w�zL��r�!���;-ǁ{�G�/��Sl��(�|��j^~�v��r8����GPYi+���g��݉���`{ۯ/��M��;���f�.qM�W�k��Iެw���W�8���=�#� ��4�܂}�C�8!��N�G6D��~��c��J`+S랍������Ov5͑`o��s����)����3g����*
�a�� ّr��5l_Ga�\�s���K^ƪs��)�u�J;��Hl��]��-�+�f�Ȍ�1b�v�Xm���,᭶cL���������,ԛ�W��O����$��6j�:;Td�6t���6�g���<���3|�\ML����e#e�σ�G�Ly�k9�Rհ:�����m:�e�G7�r8��T^j���l'>��o|5��{s&sR_О݅@)��y�wB�XZ�^�ʚ/�1w8v�<%��V�0�����`�k@:)�$p���[�����;6`�:�GH��.ܣ4ʈt���>�+C�ӱn�����@[w����e>�euy`�����i�X ��Od��R�:/�껝�V��,D�L{�b����q���yC��?S�e'X
�dV�4[)�a����ζ~�z"|���i����;Y)~�w�]�+��'cǟ�V��[��"6R&���bF0��P9-�_�F[R��JއIK2��J1�#����������$w]�󛐾W����כ��IkP���h����ͻ�\ѕ~	wH)gW�2�d;��`�A5��8�Ԇ��[{��HӮ��q\�2�4ݙ�_��nC,6%R{�яۢ�{��l���HDb0�{fdm��eB�%ܲçV�i�6蘾}�#����x���u�硎X}�>;�@w%���5�U��A�3լ��u��+��?�$U���Ρ��dZ=�(��s%6���VI����wx��B�(W�#0�̖�fT��é�k����B1QѸ����Ή��dOҷO�Ϡ��譳��U҇��t�r׏����#��7f���K�]�T���tn��3�|��m_�kI�X��O�������V��c\"�t|PZ��.�3��:�U�ɤ��ttx�Z���3*P��n�Z��WbI>�}^7���<Wpt}��g
��&U��ֆc9=r׳.vl�\(L�{L��YC���� JAzu;�|�8F׿.&������� "3�[�?q�����}�,�⭚4�@ቹ�g��U��{�'(�6�v������=s>�V�n�����Qӊ�U0�����kOp_�Ug�H���b��j�A��K��9�K�I]�R�z+n����۫�[�KD��g\/m�51����j<z�|��{�:�rS�����j���<.�Hk��3�B�V�K2��ʶZ�j�4
����nf�`U,��c/-'(��xK,$w��+$Q���2$ڟ6cos/	�'B&�:���B'�e�����$l1��`%���~�;�/�+VT�:�h���]3�'+M6���>�;��k���@U����mp�9o{��^��ec�J�W�[ڀr/��-*V_�l�}�հwm�:R7�\���Σa]���vS�
Gr���ڜ>�AbR��<1���Sl�!w$vw��aw���'���2��Tw���ȁR��S�t����p�7\�k��{λ��(�+;{;R0gwi�d�vZ�v�sǄ��Ī�t����-�b&��\^��u`��1�������H�`v�����4'����"��#KPz�*��^��WH�Iֶ����>��k�.����HM?��,����L�_o�woi�}u�ue��*gx���o��x�8�(�a�\zw}agwl<��NY�Xg�t��y ��N���4d���7x�7��6�������W2Ǚ�lB�e��u��/e�br����.:,s��
f��:�w�k���^���|�eU�;�8�Cg܅���5h�m���f���8>P"����m�E=WU��`�1XK�Χ���<#�D_&�\�"���)��͈�G�����ћ~k��i��a��w�黔�.���v7�d���D���M�U^Ŏ�\�ӂ~�×1�z&���o�|I���_j��B��u���z�_�vF[���f�d�o�pGJ�t�����mm\�";�H�k;O�S�]!����{0֦���h�$�; ����=l�#�"ˮ��������N��}���٘�J3��g!�"X���nh�W���6:�#�1o�o���Ҧ�]�U���f��B���k2	��EÞ�^͎>��W�ib��Gt#�)�sE*��+�A�[�{8̞l���7USS�������$�D8���y#La*FN���F�殴6�	�w�->t���oU�#ja��r��t��|�ح���M"�D	�Cm�3_UCno^̇�۲{`֜�l;�?%��O$F���ky��,�X�r�l��ۗ���'�*x��ɀ/(��ģ� ���^}Ӎ�۹�[�ډ�nv�Uۼo։[*�̂�mXHǃ�Gg�:���!_����%�q�y[VDEl�����^�8��/t�_t��,�@��hz��-5WC-��MTg��V¹8��IP�z��G�bu�A������#�Kg;qw8[7�_ޏ�ߤ@Vl_g��?a�/�����D?�_^���bg�],Z�ۼ[=am�	���9���]â�ԧ���B�Kg��]��EjRm����MPy0^Y��O�ۇ�f5��Z��ߔ�؋��_m�=�2.�F-�����C�׎����(ue�6�_r]�v�S���l��Y[r����hZZ��]M���*�֦C���|2Ck5j~�K�â,��}�������6޻؊� ɚm6���,@�I�V�za���]�H�T�ٳ�j6!�o䶦w �L\`���8�� =L�� 6x���a�W�Kv���j���:���깳ZbsPO�b���a{ *��'�~�]��9�쯦jK3OI�T�S�@jV�lwB��)�(6����v����Z*���־m�xw��&HwUl�V�o��g���9@)����6�`�������y$�Z�Mx=x�Fi�G%�pq=k���ۡR�q� �gIӻ�Y}j��w�%Q�W��ٯeLz>d�w��>�'QZ[Q�Cgf2�Ɂ�˧�_�i�iP'w��r_�n�����[��E6�#v�~ofp�h��Q��W�;ϖt�*��{0��u��^�y���!��o�Trȓp뺊��#.cU��F��sW#�ږ�z�����*5 \��A�Kqs}Ik�ٮ�i�IF֦t����fZ�O���&�q՚��B��mm>�\�� �����5�u�d���R�ʷي�5��+���hm'Dl7d��as�bO�_�/��	����:���朷����6#�Ѕ5+{�n���լĵaB��ߒƲg`loM0n��4�Mc�ԭ�䅘�U�[<�"�Z�}#��lbk�
0=f�[�os�+1IY�iʫ��-9���f�-�� ��s��X]�#p���L�E
r��g�c���˶�+��מ�#�j9ְ��A�N�1ٗѲ��z�:�\�#� v�m��{hF�T��:�l6)x���jT���1t��&E{�y[ta�\hsk�~?rXq�(��4��U�#,�\n�[����1-���x��i��ޠd�������|�r§�_�RC$��1yyb��nE��O윦zdR�s|�a����tǪ/�8�ھA'��Dn֬y{i�z�c�/��cU�D�\���z�ڊm�s���&W(k{�x�<�~�_����y{|�|�?{�|�-��P�+mڜ��X[Sy|Q�K�n[�G;bkQU� �ۦ5�2 �U�V.�\�"edT���q��C5��R��^Fη�%�8e9`������K�Hd�u����l�dvsN���֝��«���"��m��OC��sc�b�ЂXmr��N;�U�\�pJ��Ql%��en��wJ
�������6�u�l���.���WB��*k�5q�J��qg�eJ- ���t�ul�Y{W�BjY�)�;�4�7�Y'K��D��h͕�;+t�KR98o&�]ݝ�s)ԔΏ�����]t}.��{�ӻ����YbE�A7S���`��j�_��cG���6֦�	^��.C:�����]E�0c��m.L�BI}m�N��駰���(�69M�hAJ��Į�)������t:�Ezb�K�8��z�;z�5j�l��ue�A�𗗦�{�v�6�e��4�+��ʁ_c������_;ʺ�x����t�����I��(|�� n[���
�L1c�ꔓ��~�9ǜmWeu=��O����+��\���K������E=T�+��\j�,5W+L��G�7JfP����چ��^�R���7�e!�����S2f]��TW=]�Α*�ʎ�ݧ7fo`'��W5��i̮���0�
,�Q��߰>������w�����+��K�g(5�E�u�ĺ��o�^.�DZ�6�A؝��v��3P`l�+w*Ŭs�X�A�`+z�����Vj�)�Yݙ��]sV�iW�[,���u��F�2���"+^jO�rǲ�G8GV�ձ�(-Ģ���*���Ir�Rd�(b@V.nwWU̮��i��YKU���[tFpCɊ��C����m��,��b�}&'�*���^�����i�ۉ����"��vippe�KT�!��29Y��B#�W�΃l"wiV6�F����L8�d�;�wS�[[�+]��:�����:s�j��6#�d�:c_AP1�b�w��͔��Qu�,�)�lT`��rh[��޼�����֚���v �Mb�hy
s��l:f�n�{�[���^���r�u
H��� 
�WF�	�,j�quԻ�N��"�k���n��]l�/x٫.�u����-�C/�ذ��M���jtu�I�lnN��Y������]�.�
o���ټ�}yp���}��`�ӖE.w���M�w[#+pݨ2]���@j��}F+.��j9�Ku�D����iEC��gd�z�2{:7*�ˏ�v=����rٻ�w����+c��ut8���+�7R$ŋ��5o�f� eX"q���[��V+˺���W϶��\�n�%�qCgء���

��C;	�	P�ɭr*�X��n���v��L��&�
�gf�@mXFŝ��q �!)�rX��.%֎���z���>��)�ŵUD����<�G�q���۶�mmE���b&*��d�N��h������؈t�d�h5I;t�ti�$ݓE�u&g��F�����۠����F�k@Eh���ĸ���g��0Z0I�`��qn1�uӋ�ӫ�q>A���DE���X1=4��d�"��衶7c��������6�ٶn��b����6�TI弰�5�"J
+[k����qD�����lD��t��;�;cQE[N��b�ƪ����:�WN挐j{�����F(��6Ʃ5�Q�Z�ՠ��L�m��+u��v����[V��g�3SDA=U7v��T]�Lm��j�u�ڜESv�L��_������������j���)�����.�ȥ�nJ'y[͜�l�=�@of�O�м�+O�c��CX�{'i�j��y�l�a�R����*���$�����vR���V�V�A��l�4����ۈ�~�g���Oc�0�\]N�d��_�[�㕓F������y�i1�����?�+�p��4[�0{��!��7s�3@�m�r�l7�����q۶�O�Q���i��ݰ�P�L��Fd��k��\�(�}���;�W�5wV��_~���z��:.��="3ˍdt���Lp�(��
Sf�t��ׄ�'n3�-��h�QlQ���͑zDG��{o7��j2��Ӻ{�4��r�W?M-ۢo��[o{{�6����DN�ɖ����s���X��� l������,����~�w�Ìp��a���xعԤ�kL���5h����rN����\�>�ydp�t�WN�T`��W2c�|Ԟ#�@*=B���`wn���<l@�Ex�sw4�o�	�W��%�|�4�ݣ��F������N��j�� �]0�*�5�):����HU�JV]m�m��7A�N�1!�2`}]p�4�tď`1��-ݝeN��Zu�_KxV�7ք�eG{��¹�[����o�A}Ҙu+~�����s*�}��ϪNS�����0�{x�IH#�C�zu��U�lIrcHǱ ١����3憳쩉������,6~�X%���6��������S�V��A��!����Lt��9�q��3R�/��Hq����U=XmU-�x�Kl���ڎe�ْ�}'�o���չʿK���d�T-Jӕx��|�[��t��f�&���o/��nt�ѓ|6֜}&�:6JZ�����V�Vܴb/��4�O\T�xʨ3��f����,����|�,�O���&�3�2��e��N�Y�*h�nF��,�ĸ�Dp]j������YW�z�Ӄُ�;A�����K�zM�޷0�9=%t�Lkޡ��]Ty�����5:c�'���1;x��
%���M��%xD1���ν6vzj��]U�I/����#�昣�Z�g��]&؜x$ �ڋ�4���&�ث����Ow�G��[Y�ӛ�+:+�4":��T�fZ��Ê���=L`�N>o`+���Ӷc��}��N�i@�[�:���wd�Π�	����
׊��Cd�N��ٝ��$����ټ�,��%(W��8$akSl�Fl>�D�Q��+s4f����۾:�)���{>����wWrŷ���;x�ř������9��B��t�ߕ�b������1��u�a�N�q�{S@��[P�x^��r����*5��tw����=��fDfl_@�[��y�3�x�C+�(��v��L��X��<��2����dy��?���~�s�-L��@i~���^��������3<�9�� U���Y&
i�=D>��Z޸���TMd]��bF+�!��Z�T�ǩ��f��eN�x��Vv�M�.�{�!�ۭ����F
�ρ(�U�������"Vn�Ș�j43�t�(���n5!�z��\a�ݲ���(�����8�fh��p+`S��R��h�W��%���~Wq�Y�mE,4c�)nx�%�A��l�v�������?�{�p<�v_J�U�d���rQl/\����j���bI�̙�CB�M����O!~��y�`�.D�������P���"g�¥�(�@�*۩��k�B��Ӌ������Z�I�՝Q-�r���%�Jd���Z�3��@�R�ׯ�)l�����>���*�˔~�I��9��#3��Ŭil���L�;�=��n��;U�iwX*�٥Y=�q>�u,��5�!�u��ݢ�&�SMM���R���B�&�:�A��V]��uB.GN�=�,��p`���1�J�d�|>�q��,��f�w�W)e�h?fqW�y��t��q���TX[�ͷb�D��ݳ6�GYP� �r���ud��f:Ƴ3c�[��ڤ>�e�x���h�ᱛ�c����c&��5��V7����jZ�nu�}�l�d_�y�Uq�nn�6uEQj�'���{���#�+� �l��6��_�-�.�F}a��"��6p��{e���9�6�m%���ę���l�A�!w��W?Z��4^G?�{�`Ϥu�6�#\�Q�<~V�Y^仠!Ԩ~mv�y��Kj?Jm�:'����ϰ�W�e�s�����k��_,�ɏ�OY@�G!���7:���]&��f`^�w?�j�A���q���)x��Ma��|< t��$N���c�p���({����t��(��T�mMz����Y�OO�2cx���y�7d�}Q�X�S���ET�w22{���MwS�f&�׮�1b���)����kY��1o�_��ꄵ�s����XV(M]5s�*$�S�V]���Y���_p���IS�D��V�J��jde��1���!r��"P� ����h����:����9�YU�̤����Y�3dj�bc�mhɺƩ�<�D1�VSiG�^��G7������,�;��pe8���/�G*�{�Uݮ���e"ݛ���u���6݀\��o]udq1�[$���ïw��VM�?1��$��{�1�����]и�R�;poa8���E��A�lù>�����6��)��B�>���J�v��dHw���ۇy��4S�w��&���Z�#q��ò͟B�Q�=��-<zK���b��YS_�X+ӵ���u@K�׆�dDvT�]�i#�*���<�v�>�mX9[}�u�vyI5U��2�3�Ᵹ�]3�d��R�k0e�q/!�'#{WZWtRXó����0�N q���
�.q��*+;QQނ���7��Q������**g�;��o:�Kv���H:��������W	Xէ�z2Pڝ&�f 1WK�=�/���Yϲ�v}�ߤw��q��s;�f����N̲��r��f��U0�>phϩ.��=Ln�e�={^�F|^C�a�fJ�q���l���4�ohL�8�I�B����tfb4;� �%�B�X[7lR>lA�����Î�1;j�>�/0�ȉ�U�]�y����_Yn*��(�U���>�bЁ����S>�k0����U]Y�;�v�OۘOg��:F@<�׵[4#M���s����j�5��d'B���mf�,�U'a��[�9��S�O�ꛬ�����P��[ �׎*���R��1Haa��^�Z�+���#�Ͼ��W�JT��J��9��L�v�%���M۾��Tohj^9�[P�l����Zi���G/ĤM�����]RHt�֍�/`�G���s�[����}r�Xp�4��e�`C�:c.a(c��3Y%��/���W�����������n���q�1���r�O��%l�#-�Tu�X�i��f�4	�}�O#2�?�Dr��f�o5��v:�yԛ*�H�r�+��ٶ�ɮDD���~����}V�T���d�+f�p73�P䌱�߶���?�c������x�EF@-�]4M�A��yf���-6�u�`�-ً��n�=������roU��(R��n���i�8vp��yF��-�UxO��:k�,H/�淵�"�;����ܐ]֩�8g�e��u�f��e7]�XGML�A�z�t^�7e'��ߴ��-�=6Ր�_N�R��d�N���4�s���啝��S|�i���NTD�q}�`���ˢW�ڡ�����J� mt�r�b�O�mn�&!>��f�m�sb��cT�4�03$?H��N�?�w�3Y��7�c���n�Gs��"���u�5��A=���Cn�_7`E�B��U�w���7�G�f&o����I.O�����ܩ��g��=��%Ml���yk���<�r|�J#�b��Y�NDbGh�دi\�W�=��� �gnn(#B��s���⾣��hS`CE�_r���r^����Dik��4��X��9T���iR?�9��wP]y�ͧ:�oLoo�r/T�e�����`��`m7*r_�k;6�7�n��+.�j�"�1E!�=�\b�h��e;-��Dh�v�u��[s17?E�&|!�`=��BS5�.����
W9CU��N3o[y�����#vZ��l��T�)VĴ�ʹ%5�z��SJ�����SxZE��s����ĠP�T|z�B��ڊxh����&���َ"�w3��{��g'�ڠ��ϯT�o>j�Ko��w�sv���W�uw�MQG�w���/�R�)V��G��c�M�{�)�alH��wj#jλ
D��:��#��\A�6��$�k�yԷu�=d�wZ"���f��nzD1�)vS]���S�|�̳_�l>dqW��F�����n��Y}��Ӯ�6��~R"�Llnb�����*|�u��tɰ��ȉ]ѝ+;O��g�����������V&vF�w%k�m�WfMj���vL�7�#8���8W)pwu�7 ­:�u�!r�`,w�YŊ,�� ���f�����&c��Wcٷ�WkDJ]�¦:qR�M�J���7 �;̛[܆�VY9�X
ܽ�>m96� �CE���&�����&2���rP�czxg�.��Mm�f��Co4y�2#��̤a�����U3��|F�(gAGp�}GX�gd{��3��an˺c
��k4���?ӂ3��7;e��ް^�H��^;�C���g0���=��m]n�N�4E�	#C��6������Q>n
����&��5'�ş�/�Sfwg���V�Q�1�B���h�ɍ�B\,�
�{}���O�ܜ����'�z���FA�S�G�n�T��J:}��'�1|b���Ю���V����c�l?�`�b��5C�6Щ9J������v%��=:�`ə˲	����/ Q
�Z�V���&@�i@�_H7q��A�3|���엘xeZ|C�&�r�Q�hYU�]�{�oL�`a��}�{aq�z�׮.E�omlӭ}n~�5��]��%�qC<ld�zM,�Y�����GC�Yin���r�m�Y�^������|*T%?��x-�����W�ӣ��mW4y�#Q��x�n�yӰ�ֹ���p@ʋC��%ZH����Ů�i'-�ma3x,�͜����)������L�-W ���	5۸���ݢ��7��rE��m�u�r4vǫ����<�O��F�;�e4�\���g+v�T��g���4��v3�y�ق4۫ؾ��m򞅽��ݶ���\v��F?i�ه�x[����I�ݠ�p��C����r::�UO-���jJ���u\�t�t������-�;��?�fτ-�r���5�7�V�;�i~+��wGkP:��#;����o=�3}5+q��N֌�/}�Fi�b�AS��e��)g>����ߧ��5���\E���u�3�Y|��a��M$���&��z�|}͛螶l畁��4�\��/{�u����ѣ0���}p�]c��w={����ݎ���o��x��~۝upk���kϮ�^+����T0c�we��u�k���0���U�_kk=E�I���,@�Ca�-�|��W��������?�Ͻ�C�� 
��T_��/���%@?�
��;��q�<�v�B�`eY�f&�V`aYVaeY�	�fB<`X�� C  C  C" C C C  C�އ�<@@�\0���  a� �=� u� ;r� 0�|aʪ�" C C( C(�C( C" C�C" C �@ʀ��� � Ȉ���(ʠ� 0�06�U�
� ��2 2��� ʪ�ª�( C C
�   �0��"��*� � "�+2���L2���*̫02�ʳ*�@� �ʳ*� L�2�ʳ
������>/�~��4�� �*��������E��� � 7�������ѿ��h���?����c������������?��T _����������g�( 
����? ~�����#�D?�@ U������k�Ā߀O���?��?�O�������b�q߽�U@VDT� 		�@  
 �P� "V% 	� d@	!Uf ��  � !� $� " �� %� !	�I\� B �  @���$ H�����������?�

�ТR�����;�����~aA��� �?q���g��ߘ  ���0~�����#���O�o��g������:x~�� *���C�'����>`W�P D?F��A�?(�����=� ��O�������������������}������ *ߚ�����_�@ U��������?P�����>_����@�BO��/���� *����̠ *�`����>��
O������n�����@{O�����#�@ U�_������L��px�������}/��I��_܈�����׀������������2�?�1AY&SYP���_�rY��=�ݐ?���aȾ����(P� �P*�� ( PE@ 	 AE �
		(Pf�HTAJ%IE)T�*PB�J��UD*	J!	
�QRJ
��IP��PJ��*)"T�$IU!%B�IIB��Q)U*�T��R��@�B��R%�)�� ��UQ[fLP+`�UUTLm5mUV��H�cj���cSmV�laZTb&�k+
6@�I)E�iQ"$� �(� 4(�n:P��P��X��N(��a��U[H1E	*�Ƭlm�����Z����MUF�SUT��JU*I3 �!p ��)J,��¥���k*�M4#m!)%h5�X� ��P[
���h4Qp g �F�"�[I�*[H���--3 26ƕ�Zj���(i�T5h�RIU("P�
��  C���Ơ%5M	5L!U�!��[�a*(�hD���-a�-I
�P�R%p  7)C(*jBR��Z�CA�Ji���kl	K$*� b3m�RT�$�D��p  3��Um0���B�J�`6*(�J	IM
����
h�1� �$��$�%T��  s� 0AZ�, Um� U�(��J��  @ `�
�` 2�PU*��\  3�� �ɀ�� jm � �� h�� Հ(��h LF� �H�Ca����� � ��` �� 4�X4(��` hm  l� � f  � �    ���R�        �x`�)I@h�h� 2220��`sLL�4a0LM0	�C`F)� ����M4� #CF�1 �&S�dF��m#&�Q���jm��J���P       p8��3H�:�[q�W6Ȃ�7Ɩ�k9bIH�i4��M�1ez;EPUKN���c�"
��� dF�"��t�(��S�@"
�Abu������?:�!�Ü �T�`1��TSd#D�*��@��TR���vZ�X��q��݊(
���7�4�(SXa��L>��(�$�De�4�'���ml�kk��ҍq�xHl928��v
[X�{��xkH�.���Ǩ�l�\��tGE��Y X�L�Yd���a7Kj�� �Å�ˡ4\�c%����:7���8���X����y��������_A�\@�+�KX�£ډse��B���Z�JT��Xv�`Z�1<��uU��EC�nPF����O)�1�[jXT�,��[h���ҹ�a̺;��f;�Ʃ-'��t�3�Whmn��
D��f��Trl�����W���-L�����/fYZ��CB�z&4�F��QncR�hæ��fU�lx�8�<뉳k����J�]�̳�mc��u��X��R�«H[�Q��P��sq�!���d�kE�ʺ)�uyd-�ȺyS2Hۤ2#�1DU`ћ��������HhI��N](���-�BCZkZ���(�	m�9�H�Y���ʲZ1��J���E#-��v.����\��X�iY���B�\^]�+�JR����ȈI4���Qiִ���-�$��n
�Z��J��7�c�v�E. �2��k��hyOh[Z����8+[4^���YF�3^X��
ə@A+Ubܰ��bì̠��QըR����G,�:*����������n�f�RX��2˦�šEw����Ԭ��I]mZV���g6�E�,��]�/5�j�`��CX�U�Oh�_-(�n���tC���Xٰ��*a�N�:�T܊�⽁��u��ʷ���t�Q��w�3���Ք���v��nL2�h���mf��-�Z;b�Ҧ�T�X�܎�ѣ1���-G!�cqڧsTǓw*6�ȅc�[7%`T�>�"���q�4,v1���ڿ���R+ejF5��Y��r�@�s4��z�F�7gC�D�_^P6�URCX_fvZÁ�26Kd`[!U���.�����Z]bܶ*9*<��2"*��.��I��l�Q��[2�mc�R�A�h�|/Y���n?�5��Rkm!׷Gie�w��x��B�m�m\��˦�׏fnjhV��O�[�)7ww��S��S0�o2J�֋�����K2�+�6���q���al�4�����x��Ʈ�����{J����gkVJ��e&��[�^֙aH0]��VF���CB;I���yt��Qڃ[���G�s.���vo]�����
�N啤V�$��q�wKn�5)�S��2�n��Z/$���k�����\���0\��!����v�V����I�SC.˻��n�Y�H�����Ҏj�a,�
'���b�HJ�L��D%/M� i� l����Y�n:�X���{��/e�`�ɳ�E=	�b����aV�E����5��ɖ-1�F�Ol^���f-%�6	������B�0:ۀ��ek`q!�ӵd�o2�c��dS/i2Hŗ�)Tu���P\�\��+�-e�{����fWXW��h�l�<N�Qj��73F'Cq8>w7[���@��J�yR���Ta�c[�d�t�f�S\�b�W���5oMm�]ڈ�/7M�Hm�Vy�.�B��i2(�S$r�`��Y�4+�X(\��������!#B����Am*������Tj퉈壍�HX����u$�i\��w�сCuy[���V5�
]jIԋC.;D:Ġy�lz1!���7]�F�t��x3�hۭ���5Z��v����[l�]�\�/R'�<4n2ࠬ=J�_vbn��1AP'����u�Z29�2�^B��6��2 �F]�-�-/��.Mۣ��1��L�x�㫨��lIJl�R��X��j-�-���2�MF�9��`��vY,�V��Ѓ�Q�C[�e���6��vj�9ZrC��#{�C�o�m�V�O��/�V٢�eJ$�&�1NG�W�����H��#X�W�"��r���b;��`��*$�0ٍ/dա曭̭�N��� �;�YD�X���`��˻�|�Go&��:�����(}6 ��7�n�^�SB�E��I���^^c5#�����gx���ϱ��cKy��ԱcDs�e���F:E��j=�2�f*�K6nR,n�+�[w�x����@kui��ZL�N�cU)�-C�T�R��!b��J���ʔ�e�A�d����i˽���I"�[wN�4kwo>Z%]7���m��ǣ�����,Uچm��k	��_=�"�Y7K�Vټ��{�'��$�Z=M���N[�[Yb�p�t�Z-`ћbQh����	w�<x.�P��7�t+W��mJܑ@�<�R ]����+טu����re9������40����9/
C�%i��jd��f&㢜0Z���vFLz]��h��dF��9�w^����&۬�%����_a��5��k���e=M�[��uɷy7mL�H_f��-^�%%�v��4��
R�KVMY�7�D�.b�QX��l2������`"֙�.�L��Ab��ݚJ�ܷ��u���k.�x&<��Tn��M�0Q��
��EhLCD#2�]nB�����s;��lu�+�N�Ƿ.�E$�-f*t��i�	QKژ()A��`l��uD�S�f����i�a��T��$4�y�Qb^T���I�4#�Q�s3q|�mn��.FDg4ndbf;A��YH�;�~r�G�)�yKm��Z��;l�xmm@��ҳ-ի�nhڼű���B���5xvc&��7F�阑�4J�ZjÖmݶ��5m[�W&��+�Z"�����[�(mZWq٧��݈mV��n�0�B��Y��^�R���mj���@oR6X|��1k�t��>�k�z�c:�o]`�]4Xh�;��K�γ�5^�J���HޤA�]�-�P�k,�ubRu��nf��t�W���Z=��y��vޭY�Z�<�A�������N�Y&���LՓ䞓W�\������4j6(ɳvBl�Rb�1�^�*ٶ��4�+ik.��r�ǪJ։�[�݊8�ҙaY,n n|C.��i�}�F��m���k��w[�bg�\bd�7H�N��˘N��*�<�t�YJ�X.9GwE���N�Cf�ڡ�Vli�N��x���si��cT5���Z^�]���j*)��d�7��j��De�	�%dͳim�kI��F!����w�Ax��M��V��*{--�j�N�d��nk�3�+>ܺ�a{�-t�#5��P�k۳�(�x.â5��F�b�#L�*�Z�2���[wE#��:�˦�B�`��J�;�2��{B�T^�n�oUX�Ed0SP�v��Ʒ
{��Z��r��:6bu��ۦ�IXLG^�����kH�9t�
TV#X{�+��))s�v����2s�jR�7R*t�*���h�(kx��[�Y%E ;�B�G �������I���V��ÛV���kY�m�/5�t�b���\�؊Q��0�'X�WYOML6��-3Z�",�5cnl��d�H�f�jꥠ���W�Q���8oN�3w�M�<�������T���l@�-�eZā#\������v���2�������n��.�]������7�R��)� ZwXô�&�[�!��f��4����3}�� ��S)b�H�);����j�-E�7d;$I�X9���*��+ƅ�kXV��6�E�I*7��:7wCL���v)��Y�fB�[u���V;�8YVT���i^�5		ռ;Nź�{���nk���n!.�n'�ل��,b�:�T���+2P<�w47[�n�ҩ�˭_7����B�Y���I��n>�a�i�fZ����>�^_ȸ@Ǝ�N�.<<�.���eӠB�2��9�����I�򡫶�x��:(�� ��?�
\�5�yvt�)VX�N��4G�-�6�d�GC 9uuI�p��m�fS� U�i3�)*�F�̬yR�j���X#�`1.�9�2-I�zSt�kV*�V��Քa��PۨY�yi�r͚�uf-�� �5 �`�Dl�FՌ %2�؆t��P��3bAK/7/�m�a<OJ32h���U7J�KI�D��a�nЗ�6�d�[�v�eQN��z�Xb�}��&|t�E�ʺ��^�4�T��X��� �n��oB�t��2Re��2J��[�mB�cT�-�ͱ*z^U�j㥘�:v�#��˼��!�)"��]�"�(T@%i��9.���! iͫj�A���F	}K>�Kkۧ��!���|�٫Y� ��d J���/��v�!l��SZ]C�r�+uj�l�2�УVV���r�죗��
��^kiFĩ`���ݛ3N"VS�G��/DP�D�(�ÛzU����ugC0�ѕ���m35Ц*dˤ��wF�;�6�79�c�|z��Ř(��+h��Q -��c�; �)X��=�����z�o����L�<]��$Z�Ǘ2��F3JmЅ�
щ��W��a��͐jz�bɶ��xwN��K(�����&����N���ي�Q��{YG�4� �4��s`e��m�ʆ�BB�֌���:��
�#Ȯ���m^I��*�Є������Zo)}c]��Y����8%�$̙G(ڤn�G�7�/wd�WR9k����&�[/f��Y��I����B���f��ݻє�5�z^�tA���^;���/�Rz�᧸r唕/+w1+c	��Z�wf�ZT5-[1U�LN�v�~B�P������=��<�5c��4��:�_#�7\mPګ5��m<K�K9��{.�:oH��&�ˇ^d%�;"yB-�!�a�U�u�6��jٶ�LڻC�xx����	�zi-�-������'P���F�X��pͤ+H�Y�K%����4�ƼٺG- .��K+z��������TZ�r�Lb<�;9Vd�(jƤ۩�K*����bi]�Y�0#u.U�ӫ2權��L�c��q��z�I�� ������h;Y9��WX�U��̝��Y�t�4�I��]�Mݠ�ݛyWK���H�if�Հ�`��Küo�%X�cKk+ws\���K6��xn�[�l���%OH�9Wb��):T�˪���	3kl`������f�����t��h}s#�Bj��C^r���sSQ�f�V�n��B�]��;����v���,Ir�6�b:*�m�Qz��bUn��kL}��*;����o4�;�k��S ��⛼�u ���eB��z\��2��ʶ�-����x	�WVl�̼r��W�{�M6%���J�6�%:!c~7�kM��,ӊ��-�ܚ�U�� K٘�&V���c2�fZ
��=�Ö́�K�^�h����0��f�.��=�c��0\��N������̚hP�bC�]iѺӆ6�9[*�s	�8��ҭ��'6_Z�T���s{��a��~��u��e��qmA�m�]��.S��|Z�7p�ս0ݫ]����(X�U��A�/=Eg!��:%�JY�+1�������Epӏ��m�R�ꕐ����ՠX�(�N�O6^�*%M;n�I�����zl�fu[��gܻ^ �+t�?tb��Ъ%fY����7��k}��
��em ��&N�{HQ�rR�mQ�C'e��jY!�؅o�B�j�:w�et7t;rm�K��j��*�G`�߶��VөoMp����G�'Γ�沢w�!2�+���z��@(�/���.	��J�adG���r�|���HW��Q�{�o*��nt���2��Ѯ��Ǩ�f���d��oR@'����b�gV������0�O'�2H��9�X7WW��!��ݷ5.V��ҵ��;�z�Z��̡�d��.3q_=+�,�5�6;�e:1bwSIju��b��l�(��Ͷ�U'�<��s�� y<�㮇^%e\�w6�-+ͭ��6�DR'>��z�F�����������T��t��G��ʶ�f�L�3/e�/;�� q�ʹ�s|k1b8��Ԃz�&m�\Լ7�L
�`�dݰ䭬4su�˱�n*�AV 8��,';��Jp��.�t�q.�oVlǄ�uե�S����#3�tĻ��U;�3��"l�Jv-�S�uǯ2	���C��1ڭ�z�-fRR�Yy3�gY��x�O��#�d���{�$FՎ��Z!-��:�J8�7�c�C+.��5�E+к�[�+�c��9R�u���Wfe�x8�ܗn��bo�AJ���ډ�����4��Y�kr�go@t4� &[�L��eN�Фh�e�e%�.6n�z#��V�Ox5���xo^���;D�ﶬ�z�L�]F�WQK^@z����f��f�x3r
��b�]�9�6��I��'d�J����3y�3$]zF�5�����wסݦ8 @K`�t&Z⸻�u��!Z{N�bs��[(��tj%3na�5;v��.8�w�Y��f�{\e5�3��F�^����u!,6��1�0���]X�z���v�� �̬��-�7�1��5g8k`���[M��3 �uM���h�Y�Z*��l�Ɲ��r�|��-����i=��^з��5�-�k�>f��ܟU����G��Վצ���+Z���S�)ʓ0hy��ڲ��h)(��:��/2�C��y�8�}s��W�RN e�����W��PZ�(��L�e�ݚ
�B���ƚ�CoHF���;��G+��!f�}ׅu��rG����I�=toY�p}�5��h-ٽY��w���H��4�*��o'6�Zw� dϜ�4�Qv��}͝9�2�9Yj#Vw&l%��|�B����ݜI��Y9��W ��.���L�X�̫ܾE��
�n>��'p훊Z'zA�)�4�����%%;98��*�L�d��mM9�=���?-Η;y�s��������nT[|e����^��:WF�����ٙ��8��{��qX�L���X^�֑��UpW�FV��Á��Y��k�L
j��WO�Xn7����d�q��]aޥ𡰙��8;��8uI�۬�Ήf���;I=��aZ�[�� m�j�`�8����[7����N�A�B�h���D9��H��-�[;&�.Ҵ�`˔M�h}	������}�m���샙\L|�йMt��xe�w��P6٫S�37���,�Z����۲��<� y��<ʘ�}���6J����9��0nu���L۴�����B�ehLo3��K�,��5��wo &Vo`ӆQ�:J9v���Ӹ�J"0y@ �ZWr;Զ��QE�1)PC�<*hgs5�W�zZvT��������hKi�U�l����3�O㝚j����gŝ��'h�jf��մ\b�'ÊYy3/��!mr��̋��͢01B�M��4X�"v�x\�>�K�}T;������� �D����<����U��.���bѷ΍�ǃx�i�c�TR��ˆ�2�i�2����t=H�|(�)-iѮǎE�`��� ���0X��P�Q�P<WNv6rFB��@�䫯�����ٽ�K�L}Hĥa7e�㧢ک*m��j�gU�G��]!yM1�9�áfv�����vݠ�%['MI@��+7-��v���Y��V����`�*N�'V�{��j���;����8Pe1�B�)iל+��!�5$��J�{j�09�5�wN�W.��<:�t�x�(��]��}O��|�cG��2���Y���������g�t��WXR�ĴR�QB+����r����F�j��\��]a�6�4i��[Qʳǻ��2�譒^��3�
�������W�H��Yvfh�t5�.0U^E��jV����+0����cp�B�bp�[�]�ھG�8�5�������̠jP�SmB�ܦn�$��*6�w��F�DJyI�~�8+�`�Z���Fͨ��Yj��y����5ux^�ܧ��:�.Tp(x�g�P3X�Ҡ��e(+�;��6!٩e���[P�����c��n^E;X�!J���oE��B,TJ��%��"�܊��I*gbX��S��m^ ���W��ɵ��:E��y�b]b�[v�%A�SVvĦ#��=�ɒ�Q&C�4m� Y���夰gL�-�ᗦ���t%�\�:�:�����V�3"Y�n�n���tӺ�;z��]#A\=5ل9[���%�iwE�d������.�N�%u̓��2&�GVk��:ξ�xU]�H�{L�ظhwv4���1�뜷`��M#�+�WX	=m��I��:[���{�mH��%�fue+$��4��D����[�µ�Ih��V��\�Ў��=�T:�έ� &/m�:�+H�
6)�}��Ҷb�Yg���u
';`ƴ�H
��oP����.�ÑEĊΡJ��Ӹ�L��^�h��s��(�H�s�����w�JK�����n��0�:��"_
p�4�R�E���V��5���m�h�4�Ώs8�k$x۱4ц_V�ZP��%ZG�+����3��*QIq�"t��W�5H�Ӯ�q���E���Ƅ6�Z��gf�ާ������t����A��a�mE�+C�����P�y�A������Ƴ-e:��Q����{6�U��U�fS ne�ڶmf�y��cg��H�,��=�Y��\D���P`�1���'k2��͓lV��_wFv��i��iU����>�~-(�q��&�Q ��ʥ�#"�x�\�a�e����D1�}h�,8�VX�.&0w���h�0H�)Lݘϋg+T�:������	C��D�@�;YcK�LqE~�xk�۲s#ʱ�YG����Ƙ��{[*0��4���^J��ʕ.VX�O]�� {Le�����4�[z.�mN�Y��VA�ୡ�v˝���
�@d�J_X�T ��)0qї٢�nRopn�h�ڃ���؛��e:15�=������N�^�h��#L����Ӏ�i����ӽgU��;&�2H�2��en�v*�{r�@V7��v���
���]t[�W��	�.WT��XxS�C]��oB
oQҨ���)��.����pOޣv��ڵ-�8,�i=X愲�
�z2^u���_k���z+�����ؘP�x�y+hQ\��\E���u
	i�`|�����N�sV����^�|B��-v����v�փp��ɢFj�}��F���7k0�ĺ���]��2�۸J}}������W@X����Թ��>�]�h�t�q�f�4`�V���dݵ �LpnQ雺y�۹�����j���M��ĸ�8��ٻr*l�i]j���5�]�N�X��LF?v;�WH�K��$�u�B�7;pA�[͊J�a�]�����K]�u��G~�<Ec��A�|���O2;T(�[!�R�H��P�����;1RFX�S�2r����uu@�<:��E�v�t�t+}�@�^�ڍ<wK�e���Z&�ه��(���%��ktO�.�%R>=�!�.�u���NQySz�S���ҍK��X痪�b�\n� ��:1�Vl��v�r9����k���qe���S�#�����7mI����2��]0Ub���űI\k�Wu�����V�oh�wH��<y��]t���jF�'�Č�|�V�>�.ẖX@�\'��C�ݎ^h��o�h,*�>�[ۋ�im+g����kBU�/3!�Y�
�H�
���X�xs�*va�Vh奡��*Ѥ�{�]M�SU3�hgY{�m{�~�N�X�^j�ì�[kWp�&�^Vs�X{Lw]F��/xp6U-��8�A�Gb�,�t;
�ރ�ݶE@��,
�|�1}��]m]�t��Z��'�ݦŧ����L�QԨ��\�0���=W�&�>�8��{���=L��7v�ز�3u���d`�s�Z�ɷt:-1�〝���%'<|$�C�18��WS����>6;:woP�3	�c)� �J]�Z����Y��N�wv$r�ӫ��Uw1.G�����iM{'Bi�klne�)B�eB�8�F*�A��m��]���j�.9a��]AEd�򾛊i�*̀�қC�������r���^^���n��v�ɩ����������)D�Nr�Pù�2`�*�]ۻ9v	鎝j�>��ժ������Z�q�"w�+=%��Y�3�l}����2r�=܏{��36[��fT<N�����U��O�;n����� fU��8�B�E��']��Ӷ��dr�(�c��`e�1+4�����]eX�R�X�+z�k-Ǉ�D���Gm����Zk�֕3�[�TԨ��4�'cQ�d��ӓca��n���K�-Đ[��(�5�5�N�ȀgDݙ�-q��]l�{B��Y{@L��0��:�d�45��ʫ��I���l��eZݧ@���tm�KI��pڿ�8��Ć��]�J=��������ѕ�U�U�b/E'T��~�yʗJ�E �5�=���^S������7�	y�R�_f��7�R�`�g
]ȝ�j=������֒��!�b�������N��dw�9�,M��m�x�.�C����+���L���R�/gR���fU�U�����6���������I���:���z�zy/�W[�wn�\/aV����YK����0�-����$���E�,����V�U�׭�:�������TÍ1an�sa�|�1r�����ªW.�dr+��e]���N��U�Y7d2�Gz�t�n���j�� *u��w=���Q�0�Y�fd��T�eB���=qմq�nd����?����5����c�Mli�*�Fă;S+"����*"Rbw��T�<q3�ӧ:Ҕ��a*�u�3v����Ǻ,�7�����a�R�iՓjTT0)|�rD
N�Bu�9��ۀHim'��}�s"<k�6�M�z�7t��#��K6w�b��})I��u�����Ἵ��Ӆ�
�fr��!�+u��>��7��Yc ��v�l����w�-�n�7�r���v��w���@F3l��Ll�O�K嶹b��>�8�VLU�Pi���%�2��1[���{e�sbD�����E�e�Nij.8�N��ыGD�����~ �tmQ�l�T���}�VU1Y�Pb{�B�ui���M|�
ԫ�U�oNu��L���\���=*[X'
лEvk�d����V?��r'�n�4X���\�oF,���)��Q�;ue�rcFN�@=5)Xr��n��}u�Nm����2,�]*C:8��m�zk��X�݋Z����K=}V�b��d$�f�7t�e��e!�K5�:N�6�?M9�(�j��}���z���қ3��x��^���y]��Z+7�%��g��h�2�u����(�=1�j3]�4�5���m3Q&ҫ�u�tTǝ����m�q�:����T ����u�͌��/nS7g�-�b�X��b�K*q�ڑH�mf_�qZ��ɘ��N��[��! ��q��AVf�:0�7��K�����e��a�eJ[A�9�ۖB��1��Fn�j����� R��v�!��|���ݖ�69�����p�p;�i�6*V�.�`��w��^�i.��밐l��x�>K�� -43��;�&^V�67��n2��u
��aJ$�:����gV�b��]p���:%��L�+J4_ o7h�7��Y�j)���˘4���&g@CV���w��9҉�Ո��d�2�nH��ϯ3S���B�Y���7�8l)B}Ü ��=H�λ�Z��+t����GnS�Vї4�L����N�6�7��am��:_G�]�8dA����ۣ���޺o	�6�#�ݑ��waT��xGͮ�"s�#?My��e���k�P��^Y��w�JN�]m��aEg�iP���&j�J���V��u3.�-�����-֖�7)�}')T��It��m���D���Y0�/B5��>�FԠ�Qg4�m��6�ʌo�>8Į��V=���ڶ�P�nIU ��Oo8eP?:��a��X�V�Muk�;��G��o��Z�u�0�;�A,Q59-��D��Z�НN�穾����G�e�gdE�k��Ą�T�r���Ī@j�j�Z�ג�������+��bt����Fy�zS1��ھ�e�V��zλ����a�u�U���]8wZ���ǥ�1�x>�m��Π�"�C�gxp�ȋ���1��B3�/��:��<�q.�=U���VhS��[	�����dg�����/k��Ӹ�r뤱���^���z!�/5�
�6�Μݚ�)n��F\���ݼ��4q���'i4f�&�ֹ^_r��-�c����03�4gS��^j��T�^� �vt�8�KM�{�P�3N�*���ќ�F��.�͸�Q�R
� dsV$��EeŦ�����ooy�� �xTB�'ѪrN�����k%���F>B�BG��hmũ���ω�֛�v����f��W��u�[D ��Ƴ���K��\�,K�;K�s���v�c�a�<Zk3�7e<���,f���nP�"�!EY��%��Ӯ�m�\�/2,Pj��;�yQ�	z��w�ef�mgZ�؉�mƟɄj���c���v��)����B�*D�ɱ����P�u�Y���+"�C�c�p�堩u�'V�B�(hU��TT��f3���gJF(:Y��՝<>)_��b����J!۩AFu��o{���8k�a*��
�,	(Uv-�[��Խ���L ���_k���t;�s&:�:���e��-�Ѭsv&����hZs\���)B��'�[Sq��)vɷ����s�ʖ]I�+�֋Ҳ���Y���;K�A��T�g)fv���+��H�4���Ii�Q��gv�ۖy+�ZA�;h�	�g��������ȍV��F�U�'ݐ�c�WF��|�t����v���\��P���O-�;l�md�|M]���gT�����$��V�Q�׊^�v.4�����q�|.��;��y�ak�*f���
��7f�*Y�"�IQ��c�T���x��=AXWe$�bXooc[�4i�v�"��F�����z���O�A�`IKjR	lI�cm��R���j�4��:�(��].�aa�J�ⷥe�w��J�"oi�&n�ܚ�
�����.��w����H1X���@�sz�(`���Ƕ&5s8�`�pN��*���ʶi��N��(4TT����4�NVg��洽�fiǐ�fi�wCp��\���'`V�[8�CP��13e��-�j��6��iH�(�n_@�@�ꕝ@������LAϏ9G�Y��ʾ�2�����x�c0�Zx�}#����5+�JYi$M��$�S�]q5o�hq��١�nJ-��Z{��"�W���Q����&�b�]YX3)|��CWb �`��0�^�T�۫�pf��K��U�RJʗj;�-�V�U�.����M8�ˉ����]*Ù\3�5�J�`��'7�+dm{J�f]#Q��C��{�)ܴ-�{Xw�Rۋ@�(��������+�Yӵ�5s��vN�2Z�u.awl�Z7 �V�}��9��Y�C��%�ta|U����WG)*!nu���Y�^�H�C*���:(]튁gtᡌ4�e@��SI|i�ɱ��<��V&��W3.�ZB��%t��*�r#�f�ځC��jS5f���D���e��ƊH�*�ҾTj֐�������)�=����)O�!iN��Bk��>iцq�ն���ݠs2�yn�T���v�6���:���o&@Z�s�/��t�R�/����*������C�$�)r��_��긎 9iW����`Īfn��Q���E����M��R�c�-��.�݀�� �׆�Y{�]F�`%�	��i�}���z{'")��T=��ݵ��4Z��K�ԣ��Y<�3\n�q�R�|kp駮�q������[�5�$1�[�)\� �pX���Z�����Ɔ艸��֮�#
�����.ƽ�����IW$4.�V���=ќC|��өЮ#s�Z�"Sb����yX��E����
�w�a�vݎy a�q�Fã]O�;ʑh�A���$�l������B�L;&���*�{R��9�Uӛ`Ĺ�on��\G*l�p�p��ucEbTy�^�����ֹ���"�b�z�H�!������wJv�� �K�SՔ��w����mv�B��-��.5M��׳3-�0 :��q�v�/k��O7����gW^Q�uŉu�(
Ql.�6���ئѵ�]�o���6����j�)���녳�fN��Mv����QD�֭_6	BcIC�9�����%�vs��YXFР�0X��Nm�*c���ɣ�{Q�1��;4V�#r��֔�R/E�*�Tmoz���.����v���e0�O�Z7X�v��u��۶�5���[� 8w��':˳�����n�|M`�u92hF<kw�����4U�}1�]�Ʀf�$=�@�s���u����"�qѐuL��7�{>z�K��%�����#�Վ( �ixu0nm���^� Ǻ2�mwa�3�H:S,۸km���ȫ-�a-U�3ڴH!���EL-T�P��f	�9A��]��7�x�M*�2m��hV���#���k��QzhV���X4�s9S �j�υ�6�T-r��Pm�|�Gs��M&sY+r˭p;���2iy��u�u��v�7:�W\�EW j3(��m�rJ�$
�q���HZ5�7B^��&�H�ID�U�2�lx��[Z�y���=Rِ[ 8+"��HF9"���e�e���z��y�i����[�&����'�b�g��:���>Nk�a���&��(�ْ��R�x'(���)<.�t8�g:� �ZuҺgSOn]^M�6��qR]Z�Wngf7��hV/�2��a:��qW�om��%;�ty���b�ep�[�����9ta�gumI��^�Y��w�D��Dب�=�Fc3�Bki�!���)�v��)�������Ն��6[�^��pl�}�*)6_PQ䔝�S�kHo#���-"�����)ST��F���b�<wc�{^�{G�9dn��g<�ME&�s~�t����ڈK�ݴ��5!F.�Z/U�bu������sd�����D��|�V�YM�ҕ+�g	WH7������w�3:�e�ާj86e�L)���Q���#'w�j���3F�6�Jc�sJ�ФZ�����siN� ����Q=i]��57��
��y��w�)�KT��G��N^cU�վ[ԏF\6�mU�&��(vu���GL"�9�f�W���Z2��u�y�y�͢Y�|wz	����!*c�uZQ���pڇTĪwt�=W��F�eq]�w-7C�����u�H�q�35���ןb�"kZ��� ����a��m�Vb��S��0�/������ ��%�H�tb�w)MF�w>6
dc5��ȑSs���WlS]s�@�~���M�r��s�u�A�6b�a�6����o���Q�A�9x�Z���MՎ�(��t��J�1��V��s��
X.����k����n��A�oW�^�5��]0w*Mԥd����:9K0���ӆ��\z�q���\}y��L��%Q.�t^c���n!b�j�+����j'�go�i���e����[�M���U6]^�1���57Y�+�Uq���A�����lV�w,�C�K�ͥ�S � ��cܨVE�I�*�Cg�ciۮ%�Ŗ#�}o�'��2�ٖ�FҦtT�t𥉉�`PW U:��W���g�m���J���������/L� .cD���ܧP�0ν�ݮ�t�q-݋@s�r���S��jr�f�F���/���t�zI�K]H�ι�ދۅ�e�;.K�(�N�Oh@_Z<7��=���'��>��uB�	��Zƥc�^���L"�A�hL�5�9� ��m�U��l+�h<4���ီ��$�u��6#BL�d�Ǥ(z%q�B�W��ެY�*t�Y�l�R����7��z�M�xu
G6��:��ʷ��]e�Z8�\� F����y����*ݥt��^�B���m����5�P}\0����U�o�Z�|���Wܗl�W��U��U��"�����|����G�?%R�{��Vg�=��G2���a�W�`��(}�Ի��řʳ�:��`	P칒��A,r��YOӱ�j�à�y��)��$n�Շqp&�&+�J7vx��0}׳��W��\�8y�������7.�8Pg�[��R�Ø��9�ff�<is*��|d��]�)Qc:/"O��������hFGPc��L�����t��P�1���K;X���y^��8'NU�r��}g6��c�n����D�n���36��Ǣ=sk��O���j��am�-�#!����ז�����wv�;��j�\�@%.˵K��D�Ǩ1�t�	9��֩_\�xp�V��K��x��t]���.u��2�u襤�zVѬ+9�A��q��%L4�(4�t֎��r�U�L��uwfq)��v\KAG6�����55���;�6�B�6Z���M����;]/�
]�O�૏p��ʲ�V���l�Mŝ֯Z���nJ��ݥ� �:���L#d(��f�3#�+�I��on������(�&��"���H��%��d�"���Ú]��U��Uˑ%IՔ��2��N:E��;���D�D�ET<^<� �S�NFts���
<�Gr�9E'����.��w3n�x���rr�\�,��s#ۮE$y�Y$�h��nE�ꥠU4���JdȊ���j�U	k�w#���Yjݓ�E�ܧps���;�HE��,s
���1ur�rvd��/"�R9N�N�Tw*�Y��Z���y\���h��N{�S�ᣆ�N(W����w�D�#��u�hE\�:k�!�A��=�3]�1��p��{O'8�Wp�C�.�NE�N$��F^���}�����x���O��כ^�'��k�</���2��%�;N�K��At��/����8��&�I�������F��5�rb��a��5���U�C�Q5¸fRM�������δ��4�Ȁ��A�uX����5�+K"�qL����Z��Tr�.��Ꚁ���CYa�c�Z>_*�G����;\0�4�z�m�N���׍�G��C{�����+���@0�銃���8ڭ�3N�M�|UV��}�AN߀U��xJ䪸3�0�f��\����h��$Ћͮ���ٌ۪0�<*����W�����\��\�}��$U���t����3j&F��?0��+\��eP��U�+��`���g����%�
��_�b8n%��(Ώ:��L��p��Ɗ���<�E�L�9C!�^♂}_f��;zO8LÁ�� �zWJ��ɚ�8_����8�a��h�gج��O)�T�T��Q�U��@<v$�J�w��mϸF��+-��T�ߠ��ثCn�h^����W�K:��(
�rمc�.ҩRdS�"Ytm�L�W���3B4ye��pb�/n����|�g[�:��]
����]���	!�ܕ[��(�x1�9g���j��R�ik,�<L���Of�R�a�����h������f���{)ϊ ct��b~������1����c�
��!U�1�T\�mE�`�R�t�3��Y$0��qE�����Է���+�@oX�p �����D�T��Oq������*0�3q@w��mT�Eg${���\��IREt�rj��T�7d�}(��kY���Ϝ^L!G%qRr\��ڸ�`����S�l�k��.�e�����Z��2�
�_t�0����K�(�&� �W���Woy�ڸ�䛺�)�N������]4J�EBrMꯔI�/�BtRV�������[�ܲ��8��0��8��?0oe�,�D"JdE�QG�C�J����]��a"���n�:�2��p���1���`��.��o�Tl7(n�����umM�aM��]�n
�촼>Qv���k	�7,�]m��� ����{eW0�����Vf����!�����z���hb.���6Tįp٤�-���F*��8bS�G�+�M<��e>�0���CYD��p�o%l��]�����#^��i���}��W���w�w�j�O�5�ga���0pt��q;*�&u��*qLP���s�@C��N������(Tһ�ʧ6�υAW��`��B��'sY��k�#E
'��ɝbA}9x|����GF�k1��[C�k�f���{7�������Z���0�iU�y�hxk��v�:�[�s�G=#Ѩ;�5��sB��"L�1�~`�k�9��/��u�U`�W�x|3����h)T��T ��(�?�h/-��j�K��z�'˻���d���5Pl8�j�Ἠ!X $DrA�K�Z,ip]���⏽���ي�]l_�0F��K=��4���9�PW�I巉gr�'~���1B89J�2vzcJ�Jf#�˃V��qH�w6��x�����B��쏚�� NR�$��0�'-f��ˬ�֚ۥ�[9��.����;�p'�p7/Y���Yw:{��el���p��V�w%ZӮ�J��xm�h[[i��&.b1Lk��pu�.o��7S�qv�Q��­���W��j�5U��r�i�'�!���y'��܉��7Zlͭ�M�&8�4e�CY��T+}f�]geOa��u䊉�(�b0Kꨚܤ<�֌u!�Az.r���K�����l�I�I{���vv��+��<UCTo[�0�50[�n�\�ܮ�����Y֔������i�
�U¸�x��ΐC��d��a�d��a����(�N摊��c���}+��4p���W��d�۳�Oz�hl�6�؜	����w�σ���g�Ui
ns����|�u���Q7E��}���q}�\c�\l��#�M����֊�9�J����F�?z�Z�O|I9Hv�W��)��tUM���g�g�f��xX�/��D�מ�[�p�}���w+�j{��y�=�b�r���W������:���*y���4-oT�m�5+�ٜ07b�z�Num�5�3s�$��^�_8V=������s�i�9+6��nMZ������`�q�^�2l�{Ǩ�hb�tR�[��#ǀ���6Sh: #��Sˮ5����(mA�
uV��@�%�B�7NJG�	�.@#1��1��W����0����q��׸�{��\p�T�.&��:(�kE������"V8��������UonDW�X��X�h�{
GT��.J� ?��8@�k�n:~5�$���.�^���5A���v�2gs���������>�p���iNI�eib�Ł����i��~�^C���5��c *����F*��.S2��)v�J�&Fm����L�3f~|`#	��G*�VTTi�(N������=��r\�Ƣ��_c��Rsm�1�LA]%U��B.9	�;���׹M�怘�N%Th����AaYvxW�����\�U˭�D>k8y
�3O�/C�L;[|��b̦�'�cSJmK��t�����v�ۻ���*B�E���ѭ��5��i̼+r���v#�L���a�2�%ab���8d0*�	y�*�����oU�ĸ5b^��~�"�u9�ph���^�LS�����O�t
�U7�S��N�����:2�XóuL��V�ɚ�/�xf��3��[ǝ��;M�F�~�Z:0v���q���rS|�:�H|�5��:�w�*���9���i��W
�A�o�O� ��pW�%�r�v�~�f����Dt����}s0��h��Ñ�)��Uu�ab�Uͥ��e�r�� �w=�8�4��� ���kE1¥^[�Ã��S��!��t]t��gn�chp�N���2Ds�1�Y�ݺ�
;�a�+˅@;�Y<��8�$Pp.��NQ�P ��OGy�Oq�? �&��bm�ۃ�.ǾǴ���ݽ�yׄ>$B%I(!P`Óx��yÅR�Q6z�s3��]
KY?OݓWĶT�T����ـZD�!F�%�P�#�xݡy��;�-��>_Hn���י�����s,6��5X�N_P�hqъjH���d[u>j�Ig��g�)E;Yϱzc8�x5�����#�of���gs�-�wt�9��M���\�l��s�w>�WP�U���s;�L<g>�+�E�ck3K�7�ֱgvGk����.P�4"�y�M��<�@����V�@Mywg`���7��#�`�.	��tݘw�Mj�j'�40���D"5�iF�v�w<���{D<�>�D��7�u���U���qJǠ	�,���b��@�1�0�]<p�l8���q"u�!\F�%d�B�+n:��:�U`[P�o�u_�Z`}$\��Z�)aZ~��/�!�Ռd�|�OW5�_w!� R�xZQ3�s�@�g�k�����M>���ͫ0T|j'���� y^ri��1Å��a67j� ���}�X:f�\e���l��^x�*G�=F��tf��w��MAZ-�WҼ�4:�\ �5{�Gd�k�ՙ�{<�ς�5��"U�/���p�U�=Ʒ5U���r:�v���������mt3.�U�S-�TP3�趐iH�s���ue>�X�	���Q��z�+�݀sUv����!�2���r�۫4�u�8Vf@��^E�.lE:L]n�j�k�0ګ��]%5x��x��o`��>�}Rx��oL������L����V�(��E�]%�
�O�jw�!����uF��T� �ߌ$Y,E�x��1�RY�[��)�7�0�v��ch�K+��BwM�)����c�u����G|�#n��WO�(�F(Ciԇ�g�)d�C1�7FT��@��{֑֣�/0���S��k�� �ʉ	�3 �ic�&5�q��s��H`TsC�r��w]ڹ��,B`8R��0�>�2���G!��:A���1��=<�e\�o3α:��5A,�
Vp[�X�2�����a��p�殻s�¼���ޭ��J?BΪ:�nR�����Q�0���6���u��P����Y���hD8��q��@���_/�.PW�V�[˸WVnj1m���w�5��7�5���UF��4)��s��A��d�zW�mK�F/ZW��B74��y�w9�cY�	��,��[�1�E�g/e�`�J�i�vȍ�k��u�����Y�r�Q@2���[���oa�q�=o��{�nK�n����7�WUU����hV��L1���ók��{��4��P�ܧB�{4.�b���{�ΈM����E-��:���
K�L~�!�N��w����l��u�_�a����i���fR��|W6�<v�1op`�Lo,�!"��΁�n(�	���7���VwPL�����H�1�]D�f�7�<!�t�luPF�+�6��H�5r�T��ٻ��^��Ub�c!����1ou ������K���+��fT`]�+��j9k���[�:� $x~}sW?h�����QvhEi|s+=D��/G�ve
�����Ӿ��'���@<C��rX���^�T�S��<����3� �Dh�;�����b��F�bX̫�������U�pJ�a ;~O,NH����>v��a��O&a�#ӈl��+D�b�����iy���v=�����P޺т�v��J�ꆮ{#
+��5^����j�zuv���9J��H��\��ʤ��3󕫭�0�p�O-���6�J���\���9��v����qŁBw���a���L���E]���~�����1���U���E�D��A�I�s5�e�ЌΎUW��0�,�r��
�4@64����Qj�SSͼYu��e�4C��`�e 'i�0��XJ(Tom��m��TʹKyu�#9��,v�0N=(����"���v�l��W���%��|Bmh���1Y�~BS0V�,g(h���U��>U(<���&N���6�����E��"8nRZ,���K�L��u���V�;�u�yH*{=���Z��.��h�+:��,���A�T���w	���^�{�OWi��X>h�i��<6��u�WX]�����e���
�M��c�>�ټ;P�4��Mu�?�`�c7�a���y5���+���a&$��-sR��Y��ݦ>0��+��tFnW�{)ϊ g������J �1���_E���SVn��C��VJ�[�Y]:�h�Ҟܼ�]e��2�+ Ț��n.�}nQ����=-�[��]��QV�2=�R��:��M��M�Q�ǴF61�+����ה�57�q���x�r}]�(Es�i�:�Gv��u�`됨s1^�`ʙn�#�|��ӎ�F�ˊ�V������y��qk���<�Y;P�@�;�#F�$�"�妑�&�Ԃ�C����/��8��1���R���tIՒ�x4M]���V���ue�X/0���2�1�6����k=���,8K�r	�m��ݱj*w]�#͔�8d$�<n
4wNV���@RI�����g7[y]f\�C)G��j��� ���p��d��7Ay.p���E�&/�wu�'���� ��!�7/X s��5I�ӝ�|�Tg_mը�9xh���Kڂ�QO�U�ږ��S�<��k��0�qv]'��ו�>��z��VH�뻈��T�e܁[�kt�7> g]=	������"�^��z&���Vc� Zf�$�������+3KE,��h��g�������XA�R#H���=�B���˚�'S`H;{�9�--(���X{@	���ق96L����cq�2Z��C�qə�<8)�ι-�%��:�(q�vY��L�x�X�3��N��7jRv&�����r�񹔇RY�ڱ�xKoM-n�!�T��m���N�a6����z�:,=���Aܩ�f�����YՉeWm�c�kDa-:�ut3��Ю�#�fU���}����{��g���u�Bm�:x��`D�Ǚ�����x�'gZ���y�d��Ih����Z��˦aW3{��uH0��.]�;��Y��:���%9�#*�ܚ;�R��A�����Y�O�*,̷��ӿ�Q�+U�6[G��-�+E��n�8
��[��L�kiv��g�gX�(�pS��U���Ge�G_��]"'>YPP�I#�ƀ�M�9�{�X%��m�2Y�:�]Iv�b��.��]h[&dA,�� �E1�:��q�ÿ��B|5����Vҕn����sئS�Um?�KT���W)��Qج�����֗���� �TU�&��R��o~FR�H�׎q�4���%k������W��*U�b���U�Yyr��k���SI��I2-iJ�R^�0�Ȋ��<-ww/'Lt�OR3��ȹ븙����ETH�N\'7u��ʢ��3i�F���-���s�)2N�̮����{�TC��s�)7D"��/;���,��\O.�
4�H�D'<++�w��<=sٚ�Yw4]���(�)�U�JT��=G͕��[($�'WVz�q��{0���,��g�y$N�dn�7\'C�NUE��Q���C�d%�r��:�I�J�6G�tȧG=�=TBOQۮw\��#$ �iNbD~2Ib_CM��^�����e����N��J�)@J�����Бgdt(i.vn��0W��+�.��ӏ)���>6]�0�x+dM���M��9�pH|O��y�(L/��n����ѹP��M��pxL?,{C��yWzM |I;�~M����D%���;����S�G�"4D! ��z~�!;۵��]��w�߼��������;J���7�����`�Âw���~O(RM!;��}цD} 1�Y��@WcВ^�_}~���|���]������}O	�!'>�|��Ʌߝ�|�~�HSr�7�1��Bw�����'��ݗnL?�㭕p.#��x��A�*�}K��uk�W��C�">�"G�s��������S
��'�������~NC���?>�~Oӧ|~����]�:WI�ӿ���4}���E����O�.�8'�z��ׯ��Nӷଧ�o���\oHx~8��>�v�����|��<�}q��x�m�ܘ_��|;��ŷ?������I��������90����}���o�?�|�����U$?�_�zO����@��O�SO�����?�_i����������!�5��o'��0���ےv�7ϟx<+�M�/Gό�=������=~����N�rag�w�$�)!�������N��
�������C��� ���nC�S�zBN|!�S��/����o�B.���BY�"DA�ǳ����sFS���<�I>��z��˼�I���޼���w�~C�F'�ǟ�xC돏&��Ǐ|yL.���ϧ��®�����	7����9O�=>>$�:az)}C�i��<���<#���c�W}M&�v�^O����i�$�{�����N>8�v��z���P�Nߓ��`�>�����ǟq���>��^?}c�Dx�!��<���Պo�{����ܮM�����pHz�|��P$���xw�9���ɅP��O�\P�_y����9]�4��������=;w���9���O>/��!G�A���[n*��V(��'V���P��OQ@3�)ve>L�^P��;z�e7�Ю*��������b�y5y�c)��#�-�3�*�<����0V-X��{������]i�T�F�[��b��h��]��8c�c��バ��������0�Ǹ���'i]�շ&���xL,���?�����'���!�܇�������r�������Aw��nF">����*3{�g_z>�#�8D��=��͏���<��}�z��6��hyޠ9�v�c���=&>;ߋcۡ�驍}��]�l{f����<����L/ߖ�rohH)���{O	��o(Rv��ώ��ɹ0������q��90���_���H��@]��w��ۓ㷧�~�{���}�>ֽ�uZ�����4}�+ʌF>�",�m��xL.��ANv�I�t�Dޟ���)�����G����	$<����n��;y��&�^?q��#�����[*��ϔ��} ���~>��xC�i���z=���0��5���<&���g��6��x�!�=Ps�_��	'|v�v��:�Ʌ=�����?!����r�����������~�{��~��]�zw'���P��ߝ�I�v��-���?�w������y?�x����]�?�~�yIM�<��'�탙�i�O���P�����ʟ81�mfw��A��bp*�����~���C��!����xL.�����)�!8<��@��ohI�����ߓ�~�����;~�㷇}|&�����>&���?&r8m������^���Dh���0}�P?x�ǄP{v��'�o9vS{B~��}������>��|�	��{���o?��܇��7 (�����~�@"#��C�����f��#�"I?�'}w�9��Ʌ�����HI������U��돩�~M?����Ǆ�?�o�O��?;x�|ps�iߜ|>~���q�����ﯾ����;㴓��~9L)����ԓ�ag~�#x@����ׄ�]�N��0�����xC�<!�<��s�Ă�v����$�P�|��;xL.W�X�Uz�@�w{�����ܾ�U��a��T5ڟ-C�����Ǎ6��&N��������iZw��q�Ae���kx��wv=��D��uH��yO�@�舁��wRǟ���@" ���q8����x�ĘP>����=�çii�1+��$�п���.	����='��]��=X��M�	���ܮޒM�|��Ϟ�����?O^�|�s} X�,DH���E�d
��1�UUZ=\��մFeҶG�6��u�|aW�u\�e��Zbl��l���E�K&g�rՋCp
��C��Rx�tS����
Á�1
"�i�mTMF͏�\8�t�J�$�w �-��hi�Oᗨ�*��@�<)V�1PHV��}��{��~��	6k�ahtM1m*��ɞ7V~�i
o֮�eWw-��T�R���Te-��TCV	dn��.����:�kC&�����N`�KSoo|��{�@���tp�s%w@����Ufy!�#Tj�x#VE޾M-F��A'�ي�e��Dw��t�h@�e�Y w �����z�V�\)U3��p��vj�
��PڨW�3tGU7�3�cA�۪۾�Hþ�ǧ��v��F4���F߸���෉uv%
C ���<7���x�Z
�$��NT���'��;�i�]�]���$������'a?!�eejj���W�^]ѷ�����~��2$�F)��Y�ȫ����g����Ee�z�)&���B�\�L����A
'�Ŏ	����9��O��b�s�N/�9�c܂*̊�Xw$U�h�K-ӯ�%�C����ל�]�f��!R� ��9�R�Ȁ��d�L -��sڬ^�3��[
�]4ŉpaΪ�\�f�M|�2&Y�TE@jv6�o���3?y�w�{8'�1�f�O��U���L,t���t�c��i���5�N/nU��g��M�!�Q:-ѩ
�f|x����xNJ�q{� u�>�G�s���pW_����x:��C���<+�t+�2�/)��7Ϸg_8�Nf9����'�����a��/�N*�<ح ?EU=�f�ub<��Lѐ8O!Y�/���dGʤ�v(Ύ����O�Ӭ{�I㞩�r�m*�����}i׫] ')�����J�WX(0VQ��s�������Ћ��my.��0�-6����8*�;V�k���ʙ�-D�))�XQ�k[��W�P�<�w��r�����Ε���W�Oq�.�5�Y'F����I�羃��������~����j�`"�h��xi�5Z0+5/u�� g���G����uq$R�X��K��&�~_b�����/�Y�w�����d�y��su�'8!�:&D��1�UA� cY�:"YB3r~��H���q#k'{����DS��y3b~؁�q�'�I
F���ׇC[�Q���i�wm���J��PCC�CQ�o��XDGq�2<.	�/�]�����(��oMB��o��Qo(�PPD�C�5�F�S�N|�,r^���7���%3M���d�S$Wܝ���W�� ��U��;t���B��P��?N�7���*wS��s=%��Pî4'���{��qBj
�	������-��:&/Xu���7���C�Ӵ��D��6g��,�;�yfѬ̥�к�U6 j���\:�^��T�nN�7��a���� t�J�GMwbĹ+ݭ<0ۤ��z3�3��D�e-K�j`U���(YȢ�}�D|;䕴E}?��@F�ϾSva^L1?b�O�Z���+Ǘ�ʹ3po�k>��u\��k__V�պ�2����y�Fp�v�2�4�(� �f'�1�a��P����4��~2���{%n8�f1��؝ǝ�U*/�b/N27�B��h��U�:,�����0ǂ~G)�i��!i�T�`f��%m�t/��uc%+K���UN�n_c�x��eX�8�=�_TU��į���^$�x|���vyEu.׳t�ʾu����(�B��Ih	��PVMM�:�Ӕ�d��]��3�i�����\�EA�r��	�j���� 3|`���$����$�t����Kjm~"�dԞ4�J@@�� \p!:���\�)�`�h��	��S�m��41�W�7�+�|JL��L�-4�AY�VZ
\X&��W��;�ע��`��LT�n��!}�ŰhT�wr����9��o�(�2_
��n�t�n2AVl�nNxn@>8j�r�  vף���3�����lU`�QhN��E���U`�)�<�S*LsqPY�Z¹B�Q!�1[[Q,�����5��@�cJ�M'1�8iQ�������F�� �/��~[o�^��wtDk¸,�zs¡�����K�^^�F��Qξ�����&6�6���,!vP�/�Q���͸y˔Z
� �
���Z�ptK , Q�p]^۱P���_�,����*�N�>j��Q�u�.�WY���n�|���5&4r���^�1mO�sgt��6V���'DE�˨w�� p�13���(�.齺��qk��,S�U�
󋃳,�yJ��*�U�����wD��َj�+nm<n��@%�#��W��4�Ƽ2�~���b�����F-f���x����YRp��:<M1n�*�,!�U4����)D׳�'I��F+�H|{@�(�S7�����*�f0����G�+"�k�b��Xkq�g�>�X������P���ʂe�Y�7���*6kFZ��V�Ó���*/io�s�Ů<�d:��3���}�}}����9]?mb��n��	pZ6��M_�}J��l֎���O=����B����Y���X|��n�̻�y@�eWd�H�����8��q��Y�,QyV:�uh�o�բ�w9����q8v��?[]ל����&�U7Er���0X������
�7��~ݜ�_]�ip�E����{R����}�*�N?���8��U���-"���Ď���G"��؀tL5�����������Y��2��B��A���w�T5_[̂*̈�Gp�$�Me�~5�C� �V��`��QɄ!���Q�4���:S�	��N� ���� j�e{��b���0ԗ�x\q��a�f����̯���d�(�3���u6IшS\�[�)�e|���{�kgC�Q��T*��8��NXsv��z�Ҽ%p�����,,u��gn�M��q�����_	m�gd�2��WJ��xl�%�:�1��C�-_N�)򵕵�E��0wX���(^�{p��-{i��K��jvp{��%Y�J�W��j�2�?}���Dc��V�8��8z0�XlX�a�,���6�CLA�t�C���Е�+{ZR�Z]KPؘ�cj:����Pd<+αh
�?��4V��g���M����z�;�b��})/�pֿ$+@�uθ_f���hR��>Q�[�R�_-�pܤ�����2��g�t���JY}��_)�U*�p�Z��}���a�FD��w�J�<#g���]f���)�t��G�T�^�
xh����Ѵ.�G�wT���tK�v���arP�' G4�cF�J��츰h�ռkJuEf_c�S�na���7 b���1�	�u!�"���h���IS��fsJp��yo!���~����N]3��^��M"��Þ\p4�x���E��gB�Hb��o�X`Dv�ZPT|�,���Y�=P��2���u}7en�)�4A��7v��]���Y��7�I�-k+Il�-����=��E�w�n�m�|�^Rf�o(S�U�X�Պ���^% �^eضlKo��<�D�n�VYn�!��~������oQl���?`��eB&�np��p�[�"*OqC�A��Y�P�K7��dC��`�vn	|i9���2F� k���ـv�R�qO.���~����%��� �����K��3�baWK�}��GT�#o"��o���H���|M?�	�\�Z��X�<�u��S�:��d���Q��������s�Pv��XUg0�'���C^W��O���cPo$�S�r�y�,a'�� s$D��g��f�o���8��f�|yo�Gp\�rIw: ��,���`q�@��L"�"t_�T\)A�~�yC���q�7���f���8>�}1+��v����K\�1�÷W6���65��w<�8�Yg��A��P���?$���#~Զ����?1Z=G�&aQ�8Q6�ã��xP��н�Z#}���}�4O�n�_]�陶����[�晊us��͢�܏^�P����Dv ��s�d#�����#�<m��t(ob���׎D�܂$�]�]�ch��Ōmp�V�yɝE��-r��Bī�t�@��4u�����MZj'����mÓ��`���1q��z�N��+ZUj��^I�64H'.�5�`��qzrWRYtdvf�./���6��e'���#����.����T�D��@AC�Ô�
C�y���w��HV��(�� ���K2�:�İj�8���E{��,3�of:�9e@7�����6�̠&3b)�=O�q��ji�֭�;W�ؤ�¹����N��{x� b�VWP}��G�h��VL{%R�q��nrS}�y���bU* *� 3�Xf7r�O��:�cye�7\gY,��;��<h��k�يt�u�0n����z�Z]5��Ӭ�VFL��Ҝ*gA;7�_s4��$b�&�fU�W���7��r����*5�Ogd��O�e�;,R٭���U�Q�oV��r��vwy+�%�vFvoCʔE�^;�����Xtd{Ɋ�)*�v5�;#��B����%�m��ѩ�X�z��!��+=J7B��e�}���#i�]�����Ф���OL�(�`6��ݲ?�iX�Xr�9ծv��������5�M��I�b�j�n4���lrU�}ԑ�G�6�P�ҩ��2���x��],��5@R�.Q���t��V�ܤ������e����Έ3�LB,{��G)[�p�V�\�IU�{�v"b��u5��ݚv�Z�0���/.�&aj���L��g��Cv��ub�ƌ6tnhr��l�H�c�W�R+>���A�9x��%oC�{b�.�2}r��T������v�QQ��r��9��"�\ �n'yW�Yά�Z��gj���p�s�P*i68SyY�W�K�urT	I�p�ذAf^ñ���R�#ER�{�C���'%�q8)+���r��3����]9�^1n�� ��R���g;e�xx�`�z�)ͬ��,�΄�"n;�b�����=���@.��^�w�]����Gg spnj�ψ-=8oA���$:�Zwq��R��HT��.���!܄ΌY��?N���"�"zyW���EZ�AIQ�H�ܭ �i�Gr@��#w]����(�uh|tpIi�9�-��w*>.�Vϊs��2��s5�9��x�**�G��N�C��\�䎄fΘ\)2R���L���4���9G��T�G%�
��9r���@Т���Er�"��Hq(̣E�+OR&^l�:T���F�r	wwP��Y�]Y��J��`�HJՕG""�]�**�Nd'gТ�AG:�*�G9ʹʹ\���,XI� �l��"֕]Li��&l�?z?����wz����q^hnK�����E�(� ��on�BTїc3����H�4�?��}D��{-��X?@�ٌ�knG�pk��bZ����*�hd�w�VC�2�{V1�̘A�+L[<*��X�D��c���N�*(�*n!�fv7���:>!��ak���cs!+��C�!D%5� ����rLJ�/Z淰�}(m}sMY��u�s�<!
y����T'sv�#ױ|��'��׭�:'� �b�,s���u�s��ƬV�K5n�Av��ro�Zu;��ƈA�����S����L[w"�>����N�����"�}�tyU�ҧ� 4n>N�{*+���Xa�@ջ�ZN
:�y(*���f�7_D�^��VR������~<+�W3toݽz�Q:����!*��P( ~�@���@��K2���8/�qk�4����Lh�f5���B�d�B!Y������._G����8?c���+���w�'-�U����K�w���-����%�7�n@��CN��U�)�}�nd��8���uù<�Q�af=!ρ�ϳuֻؖ�=�e7C�1�w;��[3�������꯾���^g���Q	��o1J��$`�����F� O��}�T���%�B�q�g�{�-H��b�1S���������4�.TkR�:E��B�Q�ۼ�|W��ת����SQ��/j��^�)s�lQ�"������m��ɍѲ:�TO+="�YY�;}.�����`D�p��y�Hr|)���J��lN��E��ҷ�2(H^���r\ޅJǿb^�̜�M;a�7��~/��V��տ��b�~AL�����*�4:�gH���x�v���Y�m�{��MCX�O���w�/z"�����F��wh���Z�_^��)jB4�ո:�T��Tu�n��4k���ƭ|��?Jh���uǣ����5ki|J�}y��g��ӷ~�;�t�����9-�>&�>�}/�(t|ǯ���XΣC������kQ���(���Y�=������X�c�ٔ����V�7�ӞS��%>������;$�weq���lT��;=6�S_{�]b������f�.�ɹ����>u�P�LRb'��׿4���ep����(�Z4^��m�LR�X�U�aV�kǟ�0�<NP��ףP�9��7�=���K��s�nmIՌ��������2f�K�Ϫ�*�g0m��|c�;�Ť���"Ֆ�uk�صY���5J��A�U�X�ƗO{�ýM�L}���������d�������~dvqA�ϹߧA�t���U?V-��;U��R�gyc��;6j�[ �	��'P~ӝ�=9��R�Rn�1D]ܳ{:�.,��:I��]���3���K+x�0��j�h�N�k'EB�[��lvҵfsQ�K)�˸oNd���Sk+�1��0�Cs�E�Ie�]�݄<�׼�+"� �*i�ݻ�x���6��fQ޶���^��_*�k��s��br&1w�;��=D}��ީ��:9�v{��gV�ϵ{�5�7=�Ԟ}�Y�\��V���D��':2m	C*���u�����%�y�*[��5y�7����ڼY-�wlul�I��a�T�)�tD�kWv��sݼn`+����S*�jI�V,˪^}x��Mf%SN+��fuA�-�ڈ��E��9ˉ�ޙ]c����DW��o��5=�s�ᩊ��w���7n��Vv��p���F���ܞp��U��O}�Ի1uJn^�=��3��{6����~��D�!�����a���5X�r�;i������xR�|.j�d���nm����5��P��ʚ!��2\�Y�JV�"����y
ˡI"��U�k)-����B|��`r�']#JuJt5���)JKU��7+s��������/z�dV+c9է�"sN�ʝ�J����pݾ+��F�,	s����G�}�Y{��R���j0�쮍���ϖ�T;~�}�vr�iS��J�}@�&w����N�N]�h1�f���{QS�=h�^��S�d߆�������*�{K�ܛf���L)7Rg�Ǫ�Y��g�a����Exw��;�L�����ǎ�zr/�U��^�>q[�ar���o�d������
D7&6iKmA##D��������Ӊ���m=psAק{�R��T��}���{����kk:�#�Gk�||O}�8��9S�+jZ�q����R�P!LM6LS����(n�� �鍳���M;�J�!+�Ds�l���[ط�Ĉ�jb>��JXw�
�_��Ӡ4�����-�	�U�h��V�`�'(~~�%j�1�تzV�%\��+�d�V{m{�.Io���ۢNXwQsY F��$s-Gt��ݥ�i)����#��}��G���x9{���?Fvîx)}{�?{{%�w
����Aj�{[B�vmMo)�:\7Qm1�:�3L�;&.�`>�hV��]Oa��q����pS�9��*��R�����<qg�i����)���'����{����Kz��A�A쎝_�9.DM2�k�Y5o+��Q�1��r�)��$J����rrL�����ʑ�	Ui�0����+(.�{s��'���<�V�?c�ְ����uQ߇M�SsK=_gF:����1s�\�eU��NUk^��js�9�(Z�}g�\ѯ�y��g`�hk~{�������9��!]���J���]az�!��O�ˌ��Ě���/^��K}pϥcN�����nCA�|+�5I��NgFrA@��䕯���b$���B���Zx��
n��ib�;Xvq�W����y�YqU�] W�0\����9��nw��89�ym�Ҏ�m��q�y���U�����������_���i�_�H�.)��u����n��v�>�r��s�K�n�����~�����s�0����c�Y�%��Rw����}0[��f��Q�w�9Kf�Ǥօ2����D�Ĺ�[ߜ��R��}���y��v�u�&�oIQ�!�mF-ovE�Ccy>[��/���p��)��sW*�ic�K��8��t�]��:�N�i���-����qM�p��Tf97Z��W�f9�:��!TRU|�k�k�6��n.�VA��}_E�g-���O�c�V�`�<�%m��7毓F߶�<Q~�>}�xa�K��-Iʞk+�*&g/tR�8�`�y�8��~�]�~�m���1�GVi�nJ���q�u�J��7�L�q�4Mݘ4��2�[����a�i�]�����{���w�y���ͮ��f��eqѴlG��T���G%>؞f\Y��z����&+�.��(��}U�}U���y�{t����Eƣ�LoZ���+|UV�7��˘'ֽ+^��.#(�ųiq߫�h}���z�����j������<���Zw�.�7�;D&6x?	P+ D�`�BF)��v�\i���N��߻:=��S���zb͝=�!�-謁�h�[�1ЭSk�낽�:�)Ѽ���S�&O PM����dS�Ϭ��ZT~�ȃ�E�=C��M����8{���t��͛+k2�����Sa�7ȸ,J�Ke<Y��NVCv���Gu3'�}�u���bi�S�>�Xz�|�rj]	�'��7�4f�p#Ll}c����vOBc>��j�����3������fRP��W髽!�]J���m�Pf���%�:�Ҳ/�
 *m_�WF��V�l�1ˮ7ͨ�����K��Q�C7��x���FGfsMCaJ4���������jw#���]Я#Mџ�'�7���\�tΖ�8U��7�U1�{���lm�j
��1.����s�����2���׳��kkʞ�����U�NwNt�w�m���e��:蔩�&���Z���߹
�hْc��j�]bٴy֪y\�
�ʏ���Z�ҋ�OI��G�����D�����G�tϊ33O���V��ˎ�狹��r=�z4�w����oC�f��`P�/�D6��<���{������9�]�j߃)g8愔�B�oV��,=_\��L�>\S];����oЃ���y���m�g�j��
	�q����(�/g�ڽm6�'����$�c�X���&o�>S�-w��<+=��+k�v��i;�Iงv�au�+,�*d���IQ8Hͼ���i[EFd��=�u��7Ʊ�����[�?�}��G�^\�M�4��)���t�W8@�����[��*Df�䀖�E�G_.|,�[�MnV�gfW˵T,?7J�Aft)+i��j��F��p9J&R;:����AJ[��uV��7ӤM�n�9Ѯ+(Oܥ�]"9�+�ʨՍ�șl�޽Y�rwsT�_	֣��+���c`�T4���Ê7�q
�M�-X��*�.u��[��������Q�&Q�����/��oW���qκT�ꉍ����̻�l�m8ov]e�oc6���=�P��F�WWQ=¤�l�M��W�U��y5o2~�FV-����u1λ��Q/n�����sT���^Щ�Y�nr�:�Pc�uW�_�A{�$J)}gb�Ѳ��{Ȏ��ޏ�/kb;��t¤��HF\��t�� *�bp:�f'�*1ǖ��[�(�JP�΅>��Y ���F�duY�:�j%&rgp{L�&�D�7��ժ��9����2s�MЍ�o{A+j���մ�+3�]�WW��r�ou¸Qv�c,�3y�ű��.��n��t��ɝB�C�HۊԂ�F���űc�7�:Q|�!��;I��+`.���,Vv��qoT]ء���<���^���
Ä6�#8��W�'}�+ 5�(K���.�nv_�[E.4�+���cl�$�rúT�O��w�梧J�&�r
-�S�\�o2�o-��Ƕ��*���ú�����ڋi�\Mfl�����HPA��
$��(�dX��@�!�9�f�5��7�cݷʮaNN��n�D���9yI�O��{v�S8.ņ��h�NGB�7��* �wS��K�@ó)uL�u�\��r�i˰��m�V�2�� ҽ�
�ݴ4)3��]��uj)�sC3�k`�c�ēFW����X�%)� q#LЋL��n[7Ck�����L�'�R��K쾽��4������ɀ�}�d� ��s��>Em�36=��5/�`f�p�?:��]4�"��ݗ@=�*#娇���o<p@X MC+������j��^�*f[�����w�A�R�K����ɭ\��y�!��-��D��b��eS��cgw;��1��r��ѡ�\�����W�#ˬ�ץ���ڤ��w�2`쏾�HQu�"�X��i⥙�83j��H��� ~t�-�Y��S1�����(�x�V��眨�wь�ue�	����Ý��ߖ�����n$�F8���<o�L���h�f�5��޾�m��V�/���۠N٧\3�V�=��;��We9�w8�iE������QZ5Y�/a"�v9B�mJ��X/����,-��ij�����P�N����U�����Ka�B�!�̌lpV�;m��2��Y��}��d�kf��J|on`�wed�����Zw�S_ ����DÕQ\��-B�"*),B3+�eE˕]�NG���r��,�LJT"�Ԉ�0�TY%E�FH�9R�\Q��dp��*�R"8���$YD�r5:@�%��Z��DY)�҈��5B��A@Q(�(��AT��e+�#�2�����$�Ԫ�r��r=�z�Zr�6�g�G
9s�TUAZ$ȪȤ��"*��Q* �(9A9TU�ꗺNl�nj�ZHDt���$�Ej�EG"!�"�͹�r��(�I-�+�=�r�"( ���\�:I\*&y��r*�?P��y{la`�����˼,
��zDw3�G�IOf6��7a��N1;�S���nI��>��ꪫ�|ch����f/3�|��ȪO��n�-�7)��ڹ��]�x�,م�~YC+�-S�"�͡�j���̶�?c�$zI�;C�S��~��d��y����y�l�����m�{�`�>�h��y�t-;ys}įN�ݔs�Y�C]g�W\�(,���G�ѻ}����m���t\9���25W�{���5�5\��{}{���˯�y�>�v�
y1Cr F�����W�\ZY.)v��줆)�T+5�]K��ИjQ��nU]/o���X4�>ȕ�6���Bw�N51��uf���K����ph^����R������w)�����.;S�LA�d�s!ЩB�1[[�OYϨ��������r��GyZ��zӺ�����jen����8�����1�%j�'qS�L����⻻2s�ow�� �U��d�'}��A3�njnDDG�|&�n�(��� ��4�W�5�D8攘ލ�U��9w<J�
5"m]m&n��zy�+�nI��9OK��������iK�ѫ~�`o�<K��>S�c�X��B�+t�~O��\C�A�φs��������o��]��\�8�F�	޵ђ�������'�nzXE����)kY�TP%E���朗z���k�����;hL����}�z3g��`bo�%�-��mDJ1Z�YT3�,���6�i,&v��m��x�U�������y=��zh���_9�Օ����oOR��.˦��)�Zhv_�21�� �����2�h����{u��i�ӼBk�׻)���^�2v��V�E�k��w3�x��5�sN㯦��kI�sU�?���M�ϔ~�����  �U�E�U|k���`s��������j�H���p�1�$M�Uer�_�����kSu���c̽o:1d�M���O�;���Y�=P�@I�����AP������6����b8_`�4E�A#q��L�vOö~&+\����i���[���[���{��3�G]��������ИR���u����Ǫ�;]n"�˳�b�ї���+XN�3����ɦ��z�i�C�ޥN��/�{"{*7�ٸ�f��UM�lr�l�ϫ˳kܶ��mR�:حU�M@!�o:��pq�|e$T�fv��~�c'�q�J��ք�Rƴ3ʀ�&�DG=�܉w�{��ã���]�+��O�~�0�U�I'ۑ:���ʚ��f�S��v��.�P��FOr�%h�y^!���5jR��nL{���	6ʦ�O`�e����g�?j}��[9.���̥X�	��zl����s��F8Ut�߾�����o���w�'�94��yo�UQZ�����r��Nm=�S�ɗ7!%��7�#4W�Xd��=�8�����o��\|�Kz���=;y{�D+ʟMS�pa�p��Z}�/z��!��[�������&�N��mN�-ј�� ��u�ΰ��?Y[�k>�M�-��7���.��ƥ��a^_�Z@����dGZ��d��v�nLV�����R��������jb����P!�K�4��eh
�Y�u���8?����M�-w�L��?¥�3��u)�g* j._t*����rB����7b�|�(s����jd�vf��$��O �����p�G|�=�:�:xX��=��ɛ��8�g���KA{�]�tJ�kjV�4^6�;�Ǘ�É�iwy����	�:��pGm�9N�6�D-6.�εň��M���x�1��E�m�F�Q�����8�%�i��"�ԇ"��Ѻ���}_W�qu������bF*Pk�������6ٮU��2��篔MSs�yQ|�1i�W�5
��i�����H'�s3}�hEư?�k�k�b���u���Q+-'{�1����^�1���i��Jy@	1��#r���^{+b�x�%�;����:�w�,keۀ�`�ӆ�s��:�Ʒ�Z��,���6~C,��� 9�j��fI\��I��Nv�g�)���H-mJ�Z��o�ݣ�#�r�Էu�0|(��6�ZN����]Щ����j�z�/g�Һ��[�Y�&G%�8�$���O��\X׵�YY�tKjb�+����q	�v�����O65��f�Lu��.2u��a�(��N��Ɵl�rK�P�)׷��L�{�kz�p�����0��ʖ�rw�ogWc�0����YZ��I��v��������k�[�{˻�9h�R�g�T��5KZ���'��nC���[�xU>مo�.D>�i��c[�*w����8���=���ơ;cӪ�w�zp��I�2'�y���*��UY�a7ݲq󟔸��<:�4pOa۬��my������Ott�:�y�=du���Z%��z����`�ZڽP�{6��m�k��I��֋���}�mK�}�������xx�~�K�R�P<g5�!�~��ܱV����7Ӕ�
�P�x�d��-��S�\�X�j"U��rنP���rj������|��3�*��<"P�FKR��9�Z��[���X�����t��x`�����sg'��}4�r/���ouՊ|��5�z�w]:s.w�R������|h_>x�
����A�n���ԨL�ZH^�Z��@\N8���Z{	=�t��p���}��U0�Zл�o}޲��n�-v	��X����2N7����=�G�+��<r��h��{9zpɿv�:?$��]h��i�]����T�&1g���}�k�^��d�4%u{u�w��yM�>����>noN�HۨPH��F�cr���FV:y\�M�}�v2�!H���{��O��n���#��Pi��=�|߹�|��p2�9S�<�ދ�O>o
o�/�v�e�H�kĻ0���S��9�.h���^n'��B�w�~�����jm�vOqퟩ�0]:�b�ӝA�w���#r���dvtW���>ObM>�"�5�u�Щ��ɞ��_t�n�Zc�AW��z$@|��W����-N,�zhW?'�瞩z�]O�aott�ҋ��\hϲ��U�h\���G^��fYJ�4+�:��c���&�=�f*����ރ+zN�y0�Mɇ-�_����-DӇ����3Gz�1�U���?f�o`�b�$8[ڹΧ�8��rZ�#ң��B���=Br I#�}ެ�p�T⎧��^V��V����+�t��{��t5�S�p��x���J0�X�u���GI�Ny�SŬ�_i�yQ:���,u�La���V�t�16++�-����g���]g��ǎ�\�h�'�;���{1٪��S��&���r��^����7��9F׋=gƚ�	�FG6�T�#ޅJŻ��Vk�E=.�p��Vi����'������n,oo3x�5��k&�'��FØ'>��k�|��Y>fq%��d��b��h�n���;��|��Ի39uN"��H���{��s�1�J�sj"���<V����4�l˦4��:4��_HYS��M��X%�u��Y*�gdT�Ĺ7\fˢ��J��~��꯯w��{ �U�N�_.��
R;:њݯ'UG=!s����|j����Ȧ��]�#�;!�V{�tl�j�Ҝ�57Э�
plLG'P�	�_��`�Gd���9t�uO�[�_ٮ��󯔸���{�IH�>����������ٞ�1	��|EF0��=�S���<��̠����:��򭓝Oy_X*w�f>a5�WKwa���L[9O�F#�-�7ި��~��^�l��1[����n�\�{�3����C�w�C�{������2ߑڝ@�D��K��Ռ{���]��#�	�.a�Z��g��au�M|��a�+�}elYI'��ޯ��M�4V�s��&#n�uֹ]��>4���7}R�<5��Cφkͺ�����N�E��6�t[OE����ږ[av����)'Sz4�H���Ě{B��L�UUU|�I�~��k� R9�i?H�$:�6��;�G��b�{��eV��;������^���EY����/=�Iz��*wҠ�A�ي*ZٽBg���owfS\_���x|<'U�n�5n��o�zj�
��SLԮ˭ԃ���Ky��m�Z��n��Mg�s�RBM�iN`�p]�ޟ��Q�r��ȸjQ��i��cu��l��N�N����@�?E50�&�A1�ɪ��b��L�Xgj��i�����?l*���s۞����Q\�#��׏y�N�z�J� ���U|���2$�`e���(�8�z`*��C;lM˻���3���&��w��ù��K���z��st鎍��4hj���|�[w�Ư0��u>��9c��&�Ώ���uv>��uoI�'4'���3Sv�u�������[(���һ�$�t	eb�+{��ֆ��4w{9��uY[�6�����G$|r��-[�5&��EN�W|j�(!̙6�\y0P��HT5��ѵ9�E��R�����w`6�����5�Y�h��υnj]8>��SZ����m�C�q]1����S�Q�ޚzD��;��i�ʚ��۾i���Y�u��b��v\�@� �/��!�3�YJ�=�[���z-	��x����m/�T�O+84ds��%�"�m�]g��0;+c�YH�}�yeh��&j넭0���6����{�E�@('[J����7,!�i���P�2�j<��6���4������>�+����B��F�һO1�X�����'�R����1=�D�����n�v�@ǧ��v�kv���3d`+p�x�w]�|[��t�/��� ���=�j=��L���MH�qW��p�6Ф��$�|v��yB���r�f<A9���u�%���r8�]�r�N���ش�BT5je�}�n��Q��=��3jZ����;5g<�L�@js	���]�:���-�-Ú��2�n}��%2(�̫FTO���]��إ;R�#�5�]D�7��+z��{Z]��R�O��9�6ˏ���Y�2a�F�ýΛ:����W}��9�^] �&tb�V�RĐb�l��8s4p~Rm��%�[���Ew���ʁ��]/wh�u����oM�jeּy>��+Ԑǎ�W�%G���u�7��0Ӄ�� 3nJ*���t�:�=.gnܖ������2��V���J�1DD,�z�4X������+lu�)�}�ι�j!#�H"��ٔ×��^�n�����TN�Vټ��J*�ȶGl>���(.�M�G��ջ�*v�]�/�jAJ���
�C%�n�y��g5e�Ď�&�[�����:W�d�͞������� e�����B��&ʝ�rkNh�^�v	�+�A��k7�Pڻ�h�N�r*�bY�Q]���G�$v�=F;������t�n�:�K��v��=�Y1�w#��]��]����`�(��**���6(�"T�Q*A���^�!wwE���Gq�DʮW*�껞�+�
�e��f!,�W�U�DD\+�teW;"��fe\��TEQUWN��E��
�t�72��*�\#�\&rg"9E��B��r���((���p�b2�L�vA��DD��N2&QWf�EA�H��\�c�Qۺ�A�Z4��Y!�UE(�r��M��(���BqJ"(��qʹQD���E*�����q����r�r��<��
*�����@�ep�X�ENn:�p�W�qtB�*)�EPD�HC�2�("dS�Qp���yԗD�2.E��\���B��*<\�EU.\T.Q�Y���t�c�[�L�)䱊���	�f�;F!W��-GXy3Q�XΏ�o�P��8��	���i	���}U{�e{��t(�e>�dߪ�R�3NJ`o�_v@���OJY�Z~�}_qQ0���Vj�]`��vX��#��"�tһ�Ah����)��ҵ@�O����a�,NzB:���{��롪 �C�yT���%��.��3��7������Օ"�&�vЙTLrǯjR��<g�vFPcn��l�|6���j}�YF�/'[�ą���c^l��u�߮��S�g\���'�R����q�\,V���j���9m3γ,Q�i�u��g�zMj�w9���F��K=Ɉ|�q��#z�6x�b)e�o4��,�O&��f"�fD<n�C�t��0BFF�#6N�\��d}�#�|#�j���ݫ��ba%zt���3�z���Jv�c6�`S�U�ߢUw�c'_]K��(J�9�3���s+.g
��b'x�6f<�ݮÕ��#��D^;���ѿ��;�Ć��Gk��h̯?u��8o϶k�@i79Ś��x�]"�=}
f56؅]��RW��J���j:���LG.��`\���VݡJ�3xm�h����TB�s
S�s!6&5���x�B�&�N���--3����~�*�\LlI�ˑ�N�Ab�7;�'u2����ux�;�G%����g�:�>8G2��A"����OYt)o��εSv�״���!zh�ottt��=�B�u�����`]��|�=��M[�6�R6;��qC�ӵ��ʎ��w���g;���� AH�R��g��|�[dR���3�1G�|�p�&�K�b1��]��=e��e��*�]#���W�-��mo��HZ���n	k�@�3��8�bn�Q� Dj��U�4�R/��cWc�iWX^�-�L�S�҉!u��&�5�菾��u��I�fwꑛ���^*=�(�U���`J֮����֯{ɹS+�P+k���/�����M��y�����ɹ�'c��V�uե������63]]�G�]�z���1��S2:I�د��ɭ9ٟn�J)�ݮ��o�\�ʓt��%!)�O���V�vv�F:1K�{SL�����
��:ԣ_r���&���ɛ<�{{�0j���Of���G'M��_om�|_l��o�e>sR5��b7�M�
c\�|:��qN��4�_hmM�AQ1X֪u��,����Ǻ��M�s�8��r�Z��k[O�&�������О0�t�Ȯ�1���b�w��^�jM\���d��Ψ�e��1V	��Z}�6�*ׄ��f��*V��qת�+\��u�s��b��`��m*n���(�p�t��9�cH�:�&�iG�������"��=A���]}�b�dE�&*����1�H����1'},.nV�G���r��!�;�R��>k m���z���'����z�g�Uf��!�룭���wc�q�gܟ���ʁu�&W�}O�Pp��M�׸��ڒܿp�>B!���A���;C�2��ޜ����a/�ޙ����5~wr��>��� �ϓcK[3v��n'&h[뼨Z;*!Aك�ʃѓ�1EL5��kmC�e�J�!��m�]���4:�;�lk�{�[]��aQ��&t[������eD9�,����;�L��0���Rz�We[�n������D7��u�zl�*����K����FK�c�к���Z�G1�e�%W�H߭��U)*��|k>��_q]&q���C�cWDa�K��V���">ط8�e�6�e��y�,��c����N����ȉ�Cy*����2�i��5g��Bڡ������c�}'����wWO��}m��B=�r!8v��q՞n~잨��R\n�<k�sO�X;�]&#;]dF�'Q��Ncn�dPnz�>�N����{o**�N𵷢\���g���X�J��d�=1���I��C~N�ST��u�U�U��^��|��R�;4���uT(W��U*u�s�,A�~[��)������p���'G��])A�Z}+�O}���ڋ�M^��J�z����{C��t=�eKV;]o�(�zn���4SF�[[���}�6mvw�=9��K���c��x&ǚ.���6�),��2�7`�*�Z����v��Z���T�!V��B��Fg2�2��"77u�T�f�Ji%t�]�0/D�S�Kj %�*�w�k�{s�G��7c7�2#�-o�� ��.ƾKG}R�����Z�{��v��8�h��U}Y�w�a����ZI6mp�VO������ͮ]��T� OJ��c��м<x�۝7�,�d:���c�h���*�a��Y�LV��1�HR�]^�{�x��3CYQ����,=�$�s����b�fL;n�+�μy6��+��	��;�L.����3�)�7ײ���{���'ѽ��c>�(�S�n��q��;���Y��7��xA�>�N?��M|�N9��LD�進v�9u��;{V�p�U�MĴ��n9�1�!��i���O�V+��6z4S�}��Uo{4��EƷ�����մ�QaSw�	�$��0�}��u����ͳ�� �#�)�2�y.����R�9W�v�D��Ijoon�VL�V
G�J�z�k�Li��n֪�芖让��m�Zwm�R_7n�'3��jh��(F�>r��pp���pGX��UUn�R�����D7��p��'�K�[�C�Ub6���JIM�����CűS������_[���=�e���A�0=��T�͜v�^hcV��·���[��:���b��T�Ծ�?v泭Ujq�-b��:������t�m��e+ױ�ڶT{
���ÈU�^�<k@E{G��Zk�����V�8�~�>�,�'��jH8 �[��=H��a�?aw���>��V�3}��s�8j�v�΍����ޕ���BR6:I#v&�ɭ�S�v��)'����2�ʘ�ힸ�BR���vr�9
C�%X���p�A}1	�ڎA�S�!���|���uÆt��6d���S��5lJ��ذ�Un�5}�%x7ý[)��+��*$R>�h����Զ�jr�:MSY6��ۻ+5K�{�*8ٕ�aR"��1ف�<z���{��K�=+�5-U�z\<�}U�P�թ'�N�tϠs��E��	���tx�L\�è��c_��J�^��H ���Y��GK�n����7sQ����Eey���Ηf��Z�c�a�s�f*���=-���h�1�kn
+��	�0�mP�ߩlU�.�訢�Ư����Cn.��ʽs^�����r����k6bo��ZaY��C1��ԫP1�n��M<����wCy���:�Z�vv�.V-���!3SKlu����; �0�z*�G��%�(Τ2���&��zX����8��;�c������B1�j`���o���i����]��ct�9zn�7�u���y]��>|Y��pFo�f���>��d<�ʵ�a=�.c�wN�4i�_=�9�Y�he�t� ����h�F�-��V�Pź��[0ۍۚ���&��ɮh�Ys��o&�ˁ;'.�[�d��n���UUUowkm�yw'��j��[ۅ��ȕ�_Nl�C;�w`�V˵�9�v�M*�C���`lk��{�A�'��R�����u#�Xdb�{� �`��t��m���>�(Ş�������'�b��[�b�C?K�-O�|�g;PV$�\D�b4��#}mmW9�'~���=k���NZ.�R�5�\2xCߟnȇ�'m���?6�h�X3)Uf���eM�y;�Kb.7����ATi�u���*̗o@J�݊��nu'b�[z6 ��=���8۩��GX�k�JZ��b�_	;,�ͭ����yՏp�������^L���F6[�!B0��J�8���ʪ��. wN�3x�Y@�N���u4�����bq1�s�����o64%E܇���#�v�����j�AO�L7����x�Q\�˕���;��΋z��@�UU^:<�!���߲ '�O��DJ���j��N=�]?c���g�.�esTw��4��<��[ʿ�`��s�vU�Ռ�o�[�6��m�A���mEə�:�Y`������*z����N�:�_cv��g/N(ae9+�� w�2�ɔV�Է���-���]]M��vZ�7��J��O������#�-����N���v�v���2������J�s*/R�W��lk���*��M�X�@H������2��c�0/�U���l��O�8��8����[���i�K��F3to:Po�Vք���[�H��z3 ��)��d�[���܅��T)'Q̬͡P%���`]������g�KH���a�4��!��*��/�8⫭U�e�l8Wd��+�mYxzBJ�q���:��m����� s75����n��'[��E��P�^�;�c�d��V����3hM�lr֓Q15�40��txcv�TY��ƺs�U�
�[S��v�k��724�`����Z�������m�r�ް�`��t� W*ހn��Y��vb�[p�� �B	f����B�a�-��0�Ky+�"@�3��)����^S��i����M���K4a�V�C�7:�wYK]�èg<b�=\*�0�sGTo��B��j >�����'d+ި�ۼ�,�k:�@�w+�H��������
��������B�߹j�������-⨝C]z�KW`��I�B���O/-�>���D(z񭼨%����f8���z'Źy��r��4E˄=�g��}�*괡RY�����ԉ ;!C/R�xa۬l}�pB��.;�\STvR�����b�&63�F����K�{;ko��٧_ٗwm�̡)�ö��ʝ�:e�N��Ϫn�Rc�[O(/��|�t�:F�B��6���.l��)<*(�Mp[�����6)K(szwD��}c���
	��P��[H�E��WP��ݡ����F�Lfs䬵X��;J��,d����q^<�t;/Yt��F�
�"�c��˝���;:Z�Nӝ�6��/':��g6���#[{��,]h���ݔu=�Kh�8�Au�p`�s�I���wR��▫F�jh�9k�۪� N���RNu̳щ���Z3jP*�J��CF�U!���\�C��hG|��!�ܝ�t�$�2*�д��`dll���v�;���K{�yQ���}Ff.2���U�9d������y΢��lV�VΏ�m� ǡ�5�o.�Α�PWJ%�D5�^\���.靠�z�⋚�·N�q�@%]�<�˼F�.���"�F+R:Guyڻ��MtoPxztv�9���k�2��4��.#fBo�2]���W�@���0��H�u��d�//E�ۜ�ל融Y�h�;Փ�A����v#{h��݄oQ7�i���z�\v�F(N���|�{������˜�w]I���AE�u���S���"g-]H���g�P�&�p�u�bt�QTʈ����:�M֑��Ҫ��摢G�D��T�5�r�X�R�D]2��YAs2��E�T�Il45�ʻ��/S��{
5��B�'<�����N�=i�OV�B"�ܸ�	�S�^��r�1���YUQTZf�*Vm94(�s�NIE9�x��J�D2�M$ܜ�iTPQq��+L�!E�]:UgsȢ���YEȣ7w<A$�wp�6UU��%U®�CՕU���H���Vv�M�#�C�r�룅�K�;��
.EAEPT�W�۩D��N�W,�r��*#�"�� ��J���˫Cʷ'�q�͜��a˺;�I��^8���z�d�j��{���6:}a�I<�a\"�d6�P��B��<����1:����U}_p��'�� ������G'M��b9v���J�V�f�ϭ)���]�7�k<�<�a��i�~}ҙ/^]i �F_�4��j �s�Z�Vᠣnم�Z���|�9��CV��^9�X�����_1����_�?n� $wƚ��zog!=z],�i֚��G��_S%'S�ez�Q ���T;q�w�{�Z�{tJƘ�2x�4�`�0W�R~Ff�5m���P���O¶<˽3����k��3{��Q�gm��I̋��haj�n^W4�K�K�C������A[��V�1!��]�����Xwf����g��'�x������x7�uo��?���w쮥�
`�^k+���%�]ɷ��e�pJ�Z���nbv@�/,bޣ���Xcz�-�q�<װgW%���jvq�Vr��݈i���WlC�0�q���?}UU��zܽ/?~T�W�(Q�u����3k�߽�l�u�G��+��~��+͝�纞�����;���}�ȏd�2���PK׫T-g�Ij�����2�%?���W����E�r�s���7�j®e���	5��-��U��o+lzo���`�U��}��[�Ljq��4�EPkp�E�78��R����	��c�S��_4���S���{���l8z�JDu�bU�k�ΐq�\tN��Xe��Ð�8�zC���7�"Tû�OI�q~D�ډ%=K{�-?\v��������*��~�3�g+������2���VR�5r�F�b}9K�Q��X{�<��v+���d�se��ڛ��YgZ�k��]L��8%�o6�M.7�V^Gh�6����.�����J�r�!rΙח��I6]����w%^nJ���Ry{�����҉GB];����Vg�Ƥ�W���<e7+�ղ~�G���Z�G����2�M�|�@a�}���o#�.����ʥ&�[^~U�`M�Ķ�WsU���aP���N�:0��_���'���5�<��QǏ��������Ւ�����;���?g�>�'�i�{���j��%�q	X��/d�u�c�y
��ek��G��3j���x��]^ޙԶ�Ӧ��4�է�.��8V��������iǙQz��Y�%3c��ƺ2+6�ZAj׍W���f�^��r$����u�,�^�]��/���o��]<5C�k��̑mT�¡�S#Z�kWZƍo8��H���[u�V��8>5�{8a�Vl�C�Js���3�m��pL�S>�{qDMf��z��mנ=���i����G�I���J�F�`�+G�Sp=kxK(��8J��#kWJ�\�Ƨ�O&(��fT�i)��5�1��ߗR�*[���� ��YTg����]kQzƼ�����]��$���'xZ� KN7�^
�����z�^��O��0�ΫciK���/xE��>��{��+9���e��bQ��{����[ez�n�L���ݰ���S�:�~uY�v^ʋ��&f{-��uW#R;Uэ_3�SS\�_M��p��Q�~�����5`1z���`�"��躵�7�{�Jx��u:��e����w�H���CY6��E�l��(�kN ��\_K�xL���;�p�^�m�`��.�6��A����.$6�S+��oG�����LЄsntޜ���;Z�N��W~���97���;�[�`r��y���!�w1��R��c#���An�u�,�Y9[��K�|���S�5Z��=�6ڥ���b��){\�Y��$S\���n�X����V��]
u�չ%uTS~�v�0�$)W���9?9fyh#fT��U�W{fy�*o���go{k��3��s'�y�����T��W@�����������%D��1O�����}1��MHt8i��!�}xѝyZ�{<���/y��1<�u7�S�[N=�E�uD`��l�S�׷�i-m����s=n9���t4�=�v����L<c���=�5�k6������m)��s�X2��ͯ|kr�dj�v��,bٌ��8��zMŪv!��fL�����iz޴6�9��~�OXu�O�޵�����V�}����Ϭ�T�z꧐��맽�Qf��ͥv�N����e����sm�l�\o;Tء��5�
']��{%��6��9P�A<�8U�Ң��;���oU���+�{}Dp�^��o,�ozr��*L64U�o�rx�H.�z�o����ʲ���V!/��g��+�[��Rw�W��hu��r��A���m��ۑ"��G��o���ϐL�	<iG%(�;�y�~�6vm\=�=��a܊��+{��	�}�p)dX�m�JO(VQ�|�-�21���`���-s�g�>�}F���zm�OO�ȮEfڤ�,̢k�D�\��o)HM��	t��̟���v���m�B��������ŋ���yk&�By����:ԣ\�����b+9���3(R��ʪ��Sف��&rq��t�N1�J�ѕS�-ٕ5�!�R5tTA�I���sY�|����T&%�j3��heC��;�d�����1�N�;��A��ʒ�bQ$�J;d�ϧ@���[]\0�L�s���,�1T�(gn'�{s��	8Z����#��lۢkMc�#�m���D��{/N�Έ�o-W���z�Zϯ�ٶ��j��9�g��+�֠�K��5�x�5R��o-���;��������m5z��7=��-J�x�Z_��|��p�n���/��*H�n{�qe_�>���d�K��X�R�Q�6|�{F������߰��2u	��>>�+���D&'��/.��v=:��l/Ub��`�:�����ɕ��׃�2�y��/���v�`�5�t��-L�:����8��ncz���/F_��߹d��6��M�v+%f�1l�:a}"�~���qQ5�)��>]p��V׎��u|����E�}�3�e��a֖������:�u�M�T������e��ξG�5�}��OVi�Щ� �+ii��a�%8�Dq����oֆu)��f��Վs;g~�\�Y���/T�y.����v���t1ovK:��0��r�R��\�<H�=P��z�� �V�o(���V��]2��I<��l���ƤÄ��`��|�r�
bi��֪����)m<|�<������U{Ȭ��{�\�|�V9)��x���J/ax�zQ����Yjz���2�)3�u�[�!�p���5�c�s[WVu��P��T'����?�Y �2&�i��˜,���w?9~�<��J�
�cx���M҅�����jKշ�y����t���p���O���2s7�,�맜��)�*^c�~뺵v�6�l�Q�B�%"wv׍�	��aG�%y#�{�G]oG[J
h�t*��W�C֎����ڶ�_���۞Si�7��E���= �:wd������g*n�T)�L��nӘ{��tJ��Yƹ�÷�����U�TU4����KU���R��%$�6-t�Ee�7���Z:+�;[�����ٿd��~氮�/a�;�o2`��(���g��%]V�7V�v��P7Qb��J{�3k��؞����������
�X�����Ѡ/��D7��A��s�P����U�M&J�˫���3;�v@��N$ؗ�b+q��̽K'�p�=�:���u+�6:�Gt���$�o��훾�<�s���!��<�vw�C?K�M�.�w��ćѸM���W��浖��O�&�-��Hg.��3�%��-�ih���T�sݴk�-���J���g�;8�}"��^�곸Sf�Խj~�s<�q-�;�Qwh�Vf3�2�p�������b����2u.�굧�x3���m���� o<�Ů��A-H�yxՅĵS�{irA��ks�X��V>��%��k���r���[�,���]��0�CtpW+��9Ma��+�{��[���7˻xI�m��/ĭ����|3i�f�����.ָz2\Vpܵw���ڦ*E��w�U�q`6�%���X�65�Wn��`J���/d���"3z{�-��y�%ޝ��Ts�@��w��� �,c�C����ʟ��.1ZYe\T�\��[M��f��#�4�,�|�m#3h0����{CL����r�;7�fTG;C��ט|�9� �K+D-�6�Vz�}�+�8�/zc	�җ��S�Ί��Mտ)i�|}khV+����L�mWa~\�Q��*ǯ{T/<S�C��b�1���`�*��"`�kr���T�ü�� Fv��x<%H��=�̴���f�r�/~ї�i�H�����اu�K����q0c���$��^t�:R8!�A��)[�hi�f�M��x2im@�?�����N=͘�-\u�mq�I�M/�iε����N�\��s2�*��[A���7����S���)�s'S9iһ�L�䌩��V%���Չ�F�Έ�S��Np4�m�ރB���J9��bf�J1�����-�6Κ��ޣ�:S&�#X 9����9w�5H�����,M)SJ�\�x�U%ef��R��s�q�N���4*�J�s5�|��H�0wb��qSrwI�	C3Qv�5�q�{>�`y��ݛ�>��u��W�S�Cp�ɮ��D#l1g(MJ�!��V�)웍bv�pLF���+)�j�o7�m��,�I���#9`+��ut	m�=���v�X����HVon�ک����f����{�<��4"��җ)pË�ݜ�2�f͔(U���H������ھ���]GM������m%�Ы��3�#ZӶ��t3�iFr����cC;/V����Zu�Vq;a��v/P��:m���3i^��	ua�[��3(�CV���[��^�I��	��H����w�HH��=��/S�u�7�=�7K,��۾�D���֊��u�k6��os����,��:��� �	;���(ś��q����R�)��n^�3Q�T���G�%R�/t�Ew\]1�ܹpyN�U��A4:��'�d�mqM:��6�[�yVs��������:���
]��� ��y���s�n]���zRF��)ع5;y�9��6�b��f`R���jlܲ볪�Kmɉ|�A��\���Tuԕ������ӊ�%ZV�q`-l�K�2��D�0������� GmR��d�cRפ}Β� vVZ*��]�IݛW{�!m�N� �Mn�E���'���UÚeL�E�������Q[c2a�d"0>6NI����Q��ukh��wT˳y��Յ��]�*Sߏ"��/adwe�h��)���b<��Y��>�V�$;Sw��2Nv�>�D�#��wMX��!�"D(�'L��,=R�<��;k9`��k�nQ�^YՒQ�.���6P۷Q�@Y�S#vu�a�{}��Y0��w��]��;��j�3��Р(
�:��5�V��;j�!*N!s��UU���U�
L�*�pH�"'P:���
��H�S�DF���9�H����S�
%nW��%d�K

HU"�a�N�^�p��"�w*����9�s�\��$n��Qk�\���i((���$˧b�V�Dx�ܜt��EA0���3�-���)<��]�=w4��Jȶ�N�dY�wa�:�����;����Vv*ҹp���Ag
�T�r��fESrNz;�&����n�ӎQN�	$� �Bt���Fw!9�QBBT'I�rn��h�Y�A����;��������&̋Q"��twG8�v��8'��<==��������ѕ7^o1x��#z^2CQ���#�qBOb�U�C1��8�+��Ҽ�ʅڪ��7L����Iw���K~��ޠר<�_��x�k����N�/�iu�����xQk�)��FL����}	���jlI}���v�6�-��۲9�l�?4��o�Z� �GL�ɥu}%7�����g"b5\KLGm��_f��Y���G@��n`�ߨ���Z�*��dʶ�UnPGj��K��������Sõq ���z�S���7�k��;����_z%.ct�hLb���iQЮ-!�jz� ���p�\�+w��`x��*�)��
>}�[�W�/_j����!�������<跻g��1�1��	fzH#bef�8ҕ^%W�ʚr�e�.��H@.�W��{� o/b���/6�@��kS�E<�NM ]��h%�^���jW8ٻX��^6��kxV���Y���.�,���ٖ��z���i�cĢm��U����c�{�oJv-�|Õ�.Gd�s������Y���M�dw�Y++O��x���������^��N�.�V=½�+5b�pd�l~�ƼS������BhH��5g[�'��S3��Q���u������;�'������H6'�������͸�ñ��2׶�f��[0;OeJً��u�x��"�!þ��u�������)��9�sv-�e�Q����j�	��4s�{��\E^��f6�m��ݲ�8Z��ڠ�RC��:���o���>�뭤���48-pq���د���m�������B���{���V\D�+�&��O^@�SA�q
����"������Tŵ�v_ t��
�Z29�?���y���5����-�~4`�QJ�-Y�Y"oCq)v��&�Gd��f)W����N+-նg�q<�SC��>L�+��;��ҷ��H������eg0q��|b��/-��P����"�s�kFr�y��<�Ū�}Vj����z8�)r���J��U{�e<�)l�N�md~
&�o�-��E��}]/^9Ɩݿ��Zw��j��a�-�#Z��6xn�lx���=�J�{��7�A���ߠ54�Q[���3�{=�5��qʛ������,X�=���>�o6���z���3��Tae^���ޘ��
ὛޛD6�+!��L����:[�(J�����bU�#������o?q	��
gm�M�q��#�`dl�F)��U}��Ej�n�\+��|�[O��N�r=땔#�%(�js�Ul���G�l���-G���N��.�m��`ONƌ��JY���^^����l7����9ـe_lt���W:��c�rΐ�wt3%C��BS6k��?U�ʺm�U��Zi���q-��!\=�gm��O��JQ�]?r�7:���UNf755��6��&��잠���S�oD�"]�=�.*�v�}3.l��>7F[OlQ�aW��z\Jʶ[ǭ�iU]��}���eٞ�g9�}�5��⺳gm��.-�9�u�ğ�r7�ګǋȷS9A�5]�4�--B�Ϋ{�����ܜ�8E���{��Yzc���:���������J�:+Y����gu|6��ǚ��{�Ag*��2�'[�):�Ycc�5����`��v9�^�i�g�TG;h:��^|�t/7+0����O�
ޙ\���a��Eo��ћ���a�`Չ�ɪ��N�F�%��,j��+8�h��������Z���ޢ���E�;�~�·�Y�]�[�Y����a����,���C����B�Aq,pv�rNf��.mC
��XǱ{ӆҺy�y8�Tj��8�'J�8�[φlT��O�z'�m~7ݜ�)�c��3r4:E=Sy��
�YF����]�^3WI>�H(�������'>imBT�j:T�G)0I�4rcy���ƫ��߻ǐ>'���[r��W�\���"(�B&U��܉�Y#�`<Unn�
O����v'Ȗ�n`d�ն�oIz܈jX��T��Y���y����=.bm�&j�����DN��;���Ӫ��&g�2f�r��V�jb�j*Ci���]f��fa�aB��ټ�L�R�ƥ��H��Fe��t�
�U�X���[��X��&��a�'a��&_^ͫ��ҳ��[pۀj�0�W.էE��(X4u�|��mqӶ�����'�CM�hɗv��SpQ̩�M��]ZU-KZ�%����<b��5�����M]��/����n��C/7�� ���P��W_�,�wWm��`��!9ŷ�u�(�pg�/׵FR�y\��%��+x�w�nv����×�9�=��>R��V-���:�:���(#���im��s8�{F������@�<�n?Jf��W������M��<��{dk�5��pWMo]D7�0$�xx�KŹ���M�dw�+O���m�g�7�	���q������T�[Ǿl\Ri�r�ʙ&�*n��͔�f+��u��92o}���9�����~�c�r��$���#��'yH���Y�k�����B�dم�k�ݢ5cZ���\���Wz��\*�bt�f���ۮ�����n��Ҿ��'� 
���eb�,p$��+9˻V1t����Y��٬�e\��NƢ*�u��ޫY�6��W14�o�55�8����\"�b�K�6^�Ԥ\CR�}�#_Q棷"�bm�O��N�΃
���q�Ӈ��M�M�����1�1�����'.a71�=A�.:��LFv@��I�9�P��K6�q��UgeL��p<���Z������b���1IC��z7���m0��j�_�z����L��r4J�m>�w§�{#���[���;�[�7���2��׮	�O�i�hB����1��g�W�.��r�xjN[����v��6vի=~g�jk��4Է�c�[��\�.�=�}Y1��"��#�3�ϞOMp�����<2N�����������7�Q����ʴ�Gt��Ҽj��艵qe��BL�kf�{P�����ܓL5����T{׽F����ewv٩"���JT���uK�*R�냀[��g�{�
淶�&N2��w&�Y܁�K7�@���6�?Ut�����,�3:=�*�-�)]�`�*�˧�֗���^u�чej���t�{L�U:�N5�^X����̨�~�g[.��Y��ī��o#�^���4�8�}���{�����|�GP#z26����>�1�T�î�-\�pьy���i�-����d)lz9��]�Oyyh��P�C��Ɏ��xTx�I��χ�\�p�\���h��Z��s��N���ԫ�l���Z0Bz(?Ty�1�ω�����q��Aĝ�gNu/(b��H��j	�ސ"�&��RǺW��M
^��3qO)�7���o%��E���o¡#���W�kՒi���<*	���ԙ�z��-�Z���j;��t@o�@k�P5�_��zfׅ}��2���Ǯ�eX{^���D�;I��x�xX�7�[��t,�!������{9Ň��_ֲ�^�k
�������m�/j��WFc˒��-��ŋS�zi�{A%k�J��rbnk9mX���D�G�+�x�0<S����Ls$^�59(;��CW��깄�c������eN���F�D
�!���ުC��CbT���^�����NW�N�z��w�����,H߳�3�zX��M3�6��3ko��<bo5����af�&ƫ��=Q�Zb�w��"����y����{.�⊮�v���[�����v 9���~
g�	io��[$E�9a�{}ƪC^�ի�e������s�C��6���ӱ%�4f���Oݥ1r[����ϸ~��yb��J�c�Z��rY�r�:�n�b��W��m�����]��͗���\�����Jty׫áNQe�<z@^�3�( �<��h�1�Ձf�vE�.�n9�1^���",Ͻn�������뀫������:>&/=$����B��u���&[1^����j�JӜ�VO��f�J֟�#c終�p�L��Vb��V���d�ՠ6���U�;v��$ôE�T��{��2�CuQq���]���.r�BhMU|�$Iv��룣�U�x�he�'�^OVU���b�����ԫ�{,��`O^�q���^�vuϛ �a�/<�=�l��WW�L�H�0�j1+j+���g�b���������J�1T=�ٳH��4g��P�� #��2�c�)�I~��r<ǗE߻�=��<=��a�m��)�]� ���B�	���I�}��<�OwFs�l���oR��L�a��L�D�L0|��_ò���h��1���Z������D���]p�/Ŝ�q�����^���w K9��PK�j�Ʒi�{c_�v	��S9q9Qus�<3�p�7�,�,1R��\<).<�5~���բEy�EGP��G�?�f����s��Ʃ}u}�q�\�=��H�`zc���b�5�l�;�gf��f}s9���;k޸u�_���1^^���]���
����X�p ��X�j"e�����9��`W�F�6���T���>�t�ワ�2�	�4;�]d�$��x��sh�<�4��&������=lwdO�NV�ڣ����^�C)�n�U���N�E�0�5�`M�!GF��{�T�mB��iJ�PX,q+��aT��%���W,T���x�):jQ�љV�j��ڀ�Zb&&�VY�!.ة]�u�j��t��JV��y��Y�(W+��	��L};M�Fѻ���'&5>k��p�'�37�V��V-�r�'����>r�p;��A������B�]y�1v�P[6���ϫ��t&nǨ��Huarչ1� ��x�7�AH��f�btml�Ӽ���n�a9Ҍ�L���G�y�F�c�;}�Xͷ�-���a%���@	5����s4U�d4	Ve]�2�Ƕ�Pc��q96�$Zx�A��u�%��Ή�wJ�sʝ�(��]�^���cq�Vm��M�o�vV�{�)��cJVV���]N�=���x�oQ���Zt���p6�<��.{o7MYݰ�.�"� ��|U�K>u�U��x�-꺐2T0]��%�4��+��D��5��51oWL�E��OI�AC*,��5:Y�k��ŝC�\uk� �A�kq�1Q��B"3�V�5��3G�ZV�a�P�uu�[�ǽVW��f�ބ1wJ�)�H�J5)��:�k	�2�Rɕ�5\+��zo��<���7@�:wΎ�4���t�C;��t�W�i��ցrv�z]a��9n��]�O']Bu1�;�-H���W.�2�B�b� �N��I�!P*[�Y��v�}��X]a)XfA��.� ��:n��ݏ6��х��s{u�.F?��,|R������b��zzr���j��:WJ2�y��0#jeӣ/�gs�uL��Ɋz�]����՘��+5��s\�[vm@n�S7M|u*}��v�L�$��ΐ����Q ��������XN��:I4V��p���Z� �)���:��*�^�_!g.�74�(�c�Y#A��*�9nVAV�ﳯ�`̻�EK*t[J@I��$nD[+��Eܫ���F��n6��J��Ά�9�x3+m��$.5�.���U|.������)�#&qF*b;7Gg6�	ϒ���Fi�:�Rs���'_�������Nt�9��S�Ny�8��(�w&U�織���.��nE��*iC�r�b��(rHr(H��̒iz�M�*ΐ���
NAdS���se�T,��
�ևL;L�t��9�@�-&�#��F,�!-O9s�仮]-3�u��"�Ȓ%
"��s˻�2�J�"L��,�S)����S�vr���T�"��̩+���r�㹎p�A";H���A&"��U�4�<���wT�M�]�������:��:#tЍ��k�HwAuȻ�����ɕw<���3���#�����q9w! s��)����E���̬&����Nq�%H��,�$�3���ϟ>���=�?��l�C��6�����`�R�W����jWN���72�-cW�K:��tV�r����û2�����㔏�[�-�,���.!t�v܁<Gp�(�����yk�|Dע*�	��b�G��Ƽ5�kE)����ܻL��'�l9�^�$���^�F�s�Y�tf��޺����|�EǓ�Ft�Nc_+0i�[��z��]];�=����a*U"&z���}�G0�y�{�R�^����Gҏ�c�ol�
�]^t���G ��bW��%q��)~�*g�P��r��>>�u@�ȏ��<��d
�@(p#�@���0���ݧޝ�k�<ϸ�'�i��Rڤn ��p�����>$W�cC���o΃��{�hf�p� z"NّI��/�J�C��Q�^��*$Ç�݃7����z����Ʀ2�+��&�NMm1��M)H�EC��c1ޘ^��3�����̯��}�q�az�Va������S�f�ڏ	��W�;�(���6C�-�M=��o�+ĻDԕd��+p�&kX�5Ag�t���5a9��g!Q�F�Β��k��|�����;'^IOe���-XM�μ%k�TZt��9�#�"ܧ��#�w��ݲ��tc�,Ts�'��9P��.���q���y���~�kOS�� v��\
�'����k)�Di���7��Ks�q�U������K���zc'��c�3_q��^�QX��OY<pl������B�M��*yZY�����s�������b3�0���y��Y�=iu�5gA�?E�?����KKH(|8{O���ֻ�C۞�����9ޅ^�#]�ZZ63Ѿ��x���y�_��](f�D}�l�����}xy찏L1�
�"	 �t����+Ǚ�1�s�*,y!�Ź{�
��G\�o=(>��q�����d)�!@	H�;$i���V{��'ϊ�ޘ�5�1�wN�g�r������\�@�0xv�pB(�^���]�P�c+�t1V|�CݨW��x�I��w�[�r`�{3���M˟{�S��+�-����{L�e�ˡ�w�K��8<j��չ*��p�NJ��:��@$�8��>���Z��ȹ3��7�+�Vjw��p��9�u�T����0��4�ͬ��fC.�z��ȡY�͎�U����1ꄫ�f-��πkd�:����.�W��yO���@������^RǺW���4�O���+q�w�F�]>�S�W���
��¢�"$����Mz�M|�N���#R����=z���z�O�5@;S!����+�ǆ�1��̨w�mx(�~��˿P�����|������R
d�P�e:���Ls$^��;	#q����f'ּ���u�͛q88u;��M��j��� .�ޯ����������Q�vҭx0��_�+�[΂��i�=�b{��}>�rqL�<�b��T%�"��7�y�xi����g�x��� a�W�<g<r�9�~�$��;�n�4�X:7�'�N�T17�������jDl/ W�M���n����BKc��,+�=u�w|4g�����RX� .+}qVw�M隷��y7K.�#�|*V޹[&�[��v|V�գ���>[}ȶ�[c��6�d�����ga��@Cy,r@Ŭ���۱�4�<�k��_V��j'o��q��9V�>��۽���(B�<<����ź�q7�3����3���C� Xn?M�ϩy��@��}��~4�0��US;�#�νLz�n��o]��Lü��mZ�#�\��<\�ڈ���;�1����Q�[��G�b����7�j�$�p`� B�6	�`#�Y��VV%����s� �S�+lϺ��N�����P�3p�G�^s�{,q;f��>������={�����Q�3㒁���l��ND���\h�^4������s=Z�͉��>�����H�>�Z<;��q�^ T?eQ�� T)��B{1�ސ���������T����|V Ʋ|yz@^*L8U tq��ѹY�V�/Խ��y�-�Ez��z�}�Z^�'�k�Q���-�S0�vT��3y]R�}�?zx���9_��=Z,`��\�K��
:]@���zv���9|:��i�r�n|3��F���ڭ���m����'<���M.a��0�
;��j����N̳z�����A��s��c�r�.ޤ��<[ykr��ș�!�ӥf�`�lGB�7�;]���o��I��Bbx��\NT]\�<3�p�c<���1���K4�>�^+<@������c#�NY�����Tjnb���R��{~��m��}���Ph�9��W�V;5��O�P��qEYU	|�K����V����v���F�f.�T[;�mL ����Ƥ�V@\0�[�B��o�B��J�a(����8#w=HW��
����ۋK(��,�����=YΥ���G��7�*k�g���{��ܫoEj;Gc��G��Փ��=�f��z�T8); s���R xx:<2��^օ<٢�W�󺝗��䤌N��6&: �L%P�Ds���1���Q�9�z�}ٱ���|N��:�߯�#c��G�� ;�g�W��Ey�{lՅv��y��Ќf���C;>����zӸ�w��"�˒6����v�Il`���LPΣ�g\�c˙�<zo���f�9��m�8��s]�	u�:_uEAK��pÃ��嫶��nn䋱�K�RZmq%}���9��p�\ԡHB�:�Õ���E[�����'Uv#�ܳ<����u�ÐO���ǩmR6v_����_yTM9�#t�>����Vw���>�R�\9 ��2����T&t��T/H^��T�z�p�Btf�;�6�ϔ"��4�baƍL=��n�q���kNMm1�4K�ꍭ�lW��9�u�^Mg��G�j��s OxO��U�a�ϴ�s�k��kB�����ͯ`�J#�@S��P���L_9#*�v�v���L;ɛ<w�	�Q�U�^���~�=>�@	��E}��EGLfӢ9\���7S,o��;,gG�e ����z�,9��}��`@_�~���*Q~/�L/sΕ�kV�#0�Ҭ��ϕ��S��1L��Dd֕y3���r�2.�T	��PB������%[�4����ɜ����X;�C���U��2�-
�dXa�a���͊������}��'{��?^�����+%��a����[�g����w��As��'C��>��S`/�'-��(0���J�f����qs��Ky����a���m�J���:p-��@��|�Fͭ�g5]�X����ჷ
mX�q;�F�[�j8��Du4�H��mj�G��_����h�t���Ȓ��3m%@W�y��i�}dM=�����N�&O���+�Oq�S�ݑ��G�^�
�Tw�!��'@F��!�X�4�����h�z�Nx��L{�Y�1��������'E��F��ezK�g4Hn$��K*�� a��FL�%���J�م���c�O��V���;�8�sg�������z�ǣ��h��z� eΆ �5��z�x��0�>���>N�o����]�f}�+�>�^$
��k�1+k(��iހb�ı�����u�;m�������"�����?	������ja�����d��Wn�猟Q�3���z�C�1=�<i�z�MP`+�8;���#�y�+��h�����%3���i3�ʎ��-*��1��ϻi�d�ϔ�a�u�R�f�uc�y������J�"��'���l�	����:���O|��W��FV���ࢣ�G(��"��l�/�o>��
n�8�[Cv����J�k�4�yuYg�r��[R���ًqӻ��H�cjv�j���qI��3��.��̬�YŰ\�����"��a`����u�Iv礛���Cn'j.�һ'´�#==��w `_mk;1��iT�+�����}q���!���=��v�u<��g�w�#+e 7:������-�=�"�
leCt�߻,�����f��3�7�9r=[�q�o�����`�����Q��eL9��81���$OI3�a�[ꄰ��T�t���~q>6|�a�B:�|�;�u�5��J:܁*��ޙ�/p��/E��y�}�/H��S�5fF�~0�L+�L���9|o�^��S�Y�w��'�6�kڠx�2o��LAs�+�����
��]�.5u1od���?zJ��"gǇPq�R3ġ�	&�"��e*xX�˛S)z��=_���f��S��d/���4[�j�ѣ;�~/e�%q��(5=~����t��J;�9=�e��;���nAn�@�� /WCb���ua߱��]e5�j�\��\�8��ݧ!������r�<�y��T&�t�F� ee�,����g���ɍ�[t��ų�M�'!��Ȯ�ٸ��ǧ,p8�mN��gD���d���Ln��>�i<�Mx ����ߨ��vG��C;*v$#a��W;�3ћ[&��ic����L:��4� /�S�+�*8�n=y8}Q�r����9�3���^�cƦ2���m�gKfw�/ƾU0�'��|j���zzj�úr��p����y蝯���N�8?i�=�����ǂ.`L�����b�PyN��Mi�>�{-��S�2}��5�����`Fͭ�>�W���^=�`S���`�Y,%bw�x|L:88�@s�9��O�������=w��_b�qƼ|���τ[�8ݒx��2�������c��x�;՞��y�aC�x����G��b7�x�����p ��gk�g/��ŗbA^�`M�p��qe�ԃ�r10�y��6�n5�{��/=j�W�s�������ý3�$�"��(�n=>����i���ϒ�9<���?i�u�����ԩ�@��8�Jn��Z�m��j�c�x�Ҭ�u����Vx2�06�؁N�Ny�ڳ>�r�zqw�=+�A��N"�
�KW#S9wc���ˌ���.AQɕ���LN�V��HT�1�Q*�A��3$@��w(uFe1	G��5=b7{6�y̦�G��� _�޿dxdt����4%�R"O:��|Y��F�f�b�w��A�G��1O�����=�<+����.=�� #�H	�"�N�:ٹN��Zߘ�8͈^:�j�K������*ǃ�*"~�T��a������;f���Y���1��}r�nxm�g0����d�K�rnz�V��g�qxi���}]�B��#�1�h���� ĝ�"�)~=�����ó�10����!؜*n���j[>B��	g���Lv����+�I�8=5�Ǒ�X.�j�.b��.�^��0����* ��8�4L'P�0ü���<�G"-�Ku��ď}���e�ǧ[�q�,W9#*:[:va����L���k^�x�R�z}���=7���1q�����N��YLZ#M��,o��G�O��鿆�K*������Y�|qP=��.��u���nXb6�eЛ�X�h�b<%�4��f�}�kӎ���i���,u_q��l�,�������qE���K�u��M
��&���	�7W�Fw^欴X��J�)ťd�:�.W�c��0ɒ��ӡ�������6$ibmd�窷Z5�����'��-�{�h���\�FNc È,Uњ�B3�+����u5	�j�1�h���tf�w��0�++i�ϗ	t�o��>�l�z�N>�{u(�5�e��u��V<a��zz	+k �\tv�M2T�*e���j��� ����U������:�Vpj�+���G� נ`4���4�����u_�>��+�tu��s��h��L�(�=�8dv�"���ܻh�Iޭ�`ԡ5wvQY�	�{��Xv��D�&�_�-ӷ�7��4ޕzWtV�݃F�޻�Cc��J�s�Q�W�3nQ
�p�k3{k�-�ae9�c�i�H��=��|TP3d�+"�H�;2uD�^Ū���a�����q�K�8Ɂ�͹eW�p	а�ԛإ�6�^;����V�t�(��_t1���d ��t����u�Ty�p+FU�Ӓئ�d��&������
�jξ%k�B�_9���{�Ly¹����
�Q_Yޱw8�*L��E��M��'+�u��%��{Ll��kɜJӑ�RIĽ�R�ʀ���:�*�������U�hh�A�kNT���̾���`T�mJ]�Y/s�X�
4�M<,h��tO4����Ȃ����PɁY�Jl �@%�u�>F[X�	�h�1J
tf�o[���A����A�
F�v�� ~�Z�MNo`
��i��iW��_[䶸�����b� >;�t���kl@b�fP��i���ג�,�k�nW0텒t�"�z���(��|��Y��U�:���噦��`�M�BfH����qi��;�F*;@k�7j�}�ׇ]�ɒ�-f��N@Pb�b:��ܙ68��^��v&=��}׵��qEF��:�߲��+�f��)'��S%�O�	4ME�RD����8q3�u)�Uc��n�����]̝	:T�z�w3���*T�p��i���r�N�T�aNN:,����TR�MN���S��Xȯ1�Qs��[�U��I-��̤!�ʳ'V8WL�R�MB�K�Ď��x���p��M*����Q���s3DDē�(m1D�R+&\�������g�&t��9{��-'&]��S�ҵ"���6n���9ܬ����9�ڇ-0wF�$95ڐ�9ܵ��q/6ܓ �KԣR�0�Bֹ9�Ú��C�܍MBV��y��Z��E7Q���<����ǟ�n���e�<�'MPk���F;�ήR=�.g2 �c9ՕܣR�<&L*�דk�n��r��h��^�w.�F@�g)|�3Z�3���cq]N����9�>[]��v�#��$��qL:���댙�Lk#�p�_:
�g�	\o�H�g�G��_����ϣ���O��:��.p������N�ѓ<�̋0�ߧ�m{�y���eŦ{����"*�RX]#�:�7�*���,�53�E�
 t�����^BǾ�O
��r�*L۫��S��v9d�}sP��%@_���B.����Q>:}�ƚ�U�*�7����4{�����^@!��'�Eթ�`�ȳO�����{P+g�Xaq�
wպo���9���~�Q�\�J���~�ñt��jT��Ϡ����D�����e2�v�\N���'��''š��^=^��7��D�|��!{ eΆ.	�7�������^B����zc����s}Ľ:����u�@�Z5���J��7�>�&-b��ڥ=]��0c�ϟ��P����WM����YVGg}�s�����6���i�ۯ�j=�:m��ܯ8��%onnr&#�F�8��nV��F�bMEN)cO!v6�Ĺ��i��*1V,���mj|Fod�I����q��A9�>~���
���50���^��҇{��ٕ�cڻ�tj�X��Bb~�%���)�YY@Tq�6xm|D�i�y5x��^���^��L�T{ƺ2|i��,wp� d�̐�^�u_�DM�:�y��G��to�֏\d�lޟQ�5��
d�C3n`k����>��՚�I�|8i*Ϣ\�۝����iW>�Y�������M38l\B��~x{�>gں�k�yt��r$�>�C0Θȷ;�q�@�}R1�gw�P3O����HqC�񰼥���5*�-��NO���k�ZY���dϏO��ռ��OI^^��Pv���S�a�D�8�A�`1'#�e����;��X�EY�6Lk:#}�[�.��T�)Ts�,�r�YT1��$5O����G�	��b��MN��Y��-�]�&�gp�R�ߪ�~�~d	iUt��C�(�ׁ�_�����؄���q�SEw]b��ۤ���0(9;tK����o<��FI��[�]���?hX]d5c�!(�/#g��F�79�k55��7�;y]o��<}��Y�Q7�,���;�U"~*P1�����2�L����WZ$�{�SO�+��|(�Ө~�Ҥ�qF��I���\�xcf��T��X��ѽ�s%=�}7d�_����n�A���2���W�g�B=���%��1���W�����;�=�	��T) ^;3#�fo�g{�i�=��1�-����"��3�8~�ߤ��chz���n�=S��G��h�}��Ӓq�i����B�0�F�F�P�hß��$j���+��+�Qo	Xpp�Y6���j6X�3��l*�h��~���KiX��Y�s�#W��E~)��v�i��;������\�ki�1��ӷ靬��s�i�'G���VK����l��T<���3L���z�H��Ψ�<ײ��=� u�>YLH��ū�n$�>��vk묨X�����tfԌ���{���=7�Q�lÕ�OM�:����g�:�J��̵w�o�9i�ԣU�u�4��uR�:�ץF���E`��Upԧco�mh��ە����@Ε��_g0V����Ƶ�g�R����3z�
ݖq���e��MI?߅\������zKsݣ��Z�<��0~���(�gd��òo����t \�o@��_��KƟ��2�����~Ɣ�e�4o�������޸���g��x�N�wL	�����,�y���z����Ǖ��"���}�_ML=�7E�I@�(��	/��w(u�ޅ=����4#޵L^o�̭���^�����VJh�	L�����tDK����M�ţz.�O���=�����__�܋�ޯ� #�H	�?o�����/W����#B+۵��Ǐ�A�O#��s�m�9#u!A�Z�^�}��K�C�t�H�s�X>g0�+F{��Q߉~.M¯P	>��{��qN�^�Ndo��d�9���6�@1v̊��_�d�T*���0C��|�䀤� ��7����N�{c��;[V�)�<�}g����4"��{�a6�=�c�W�Ϝ�΂�4�թ,tݑ���6��4PqX=�����咧

�elM�׍e�w�P�7˪w�q$z7𮞓��\��d��|�A���[�a��8,zrX��Xj���LV�?Fz�������9��`����q�����{��#+:]���=�o;���4OW�Idk���P��,o9#)KGN�;>�r=�I��X�3�㽝U��zzPc���L����c�\���7��_zi?*�o��2Ͼ�(e�mǯ�F��3�zX��@L#L��#��O��5Ӟ+����^�U���Y!a"�o����&w��3Q�E�*�1�Z�6��>c_z�٪����͓�!�s�_���������ig���t���g����t���>�ǚ�Ǯ����O*Djș�C�ӱT���1C�Kϼ�����/Ѵ�B��S����橊���&�I�p��BQ�q^xʿW��q+|�G�Y�i���r��j��k������1NQe�!�R=�.�uա�(S�Yu�.����+�t#n���;>�;7.`KJ;ڝ��2��w�٣:���C��ߩm�L�\YM��h��ʲ���`4�0'��]*�VN��e�st��o����xv����
$LB���ɅƬ��;�}2����,u?g�&')�<�~�t��N��Ro���тès"I�u�(hXS=���+��+��O^6�*A�/k}��M���F,�-̩1��F����@K:�v���׽\=���اyV��R�5S���K��G����׉�����@A�[YG��n��9S"�����O��8;�Y��p�|}��� W��@G��Ʀ������b�����s;��g�*��
A�d���q��0,��@�<6q��:�^T�.�!6}����������ʇ��R�)���q:�Q�,6��q�qح��N����,'�n*�����<L07�Q�6��D��.��c���'�����:NٕK�FT�/�zZ�X�o���&�*�uC���A��w;�z]w�szk客k=��Du	�$+/���:c-��� cA���N���}����x\�F��k����L���,�幑�� d�ԟ�2��H���8��I`��X��v�`k�N�_C�ǈD*��Va'}8��܄�z���qEB��SEʤЊ@��keo�c: �"����������Y� ��ws�����K�)��g�e���}�}�uR"�O����;�u��h���#beE{O<�E�D嫮~}�/v���l�L�3�;c:����{q-�t�69�y�q�r�/^��o��/�x���A��p��1�󮜠�E3�qt�8h�\���U�W���dǂ����	�9L�(
�����\��O��r�ff�����W8��&ϡ;w"<r�%�0[5�nH�'�X��烼�ޝ�\z�+���[NŹ�⇡�*^�n��~�n�����%�0�v ���z��� [ӝ�:;Ǹ����6\���� �3ېE[�P8�:H���h$���;y�C�Rʊ��`����^
#���π��*ߨ���j��\q��:��{�_�} �c�e���G�|.#�¤yޣF���ïW����~1�(w�.��m��o���s�ڿ[ژ�\L{P~'ƚy��SӶP�!�ݳ�x1l�/C5t:��_�m)�[]��ٹ�1�&���h�y���������X|Lu��@F���X�K��cLΆ=��)�鎑o���噍�U����D׺�~�#�����?td�?a�s���`]t�}�ww�׵���.�S����4&�e��LO�L;���/6kI�g�>߮�u�F{��Gu��Ϋ�G���Ki�
�
������Tmtt*N�������T}���}��	�4˵8:����;5��$���{Vi�w%!�g��ts����+����5*��t��Ⲧ-�z��EP�=�G����|�r=��і=uL�T=�&Y�'Q�27��ǵ{�Kk5��3==����덾�C��X�\Hѿ�� ��!�Z88�:�O�MeӐ���9ٯܫ�0�*�>��K�Q��n�0�J�_�;��T)<;���n�f������w�b8#N��ղF{޿dz�*��@����	]T�Ϫ���#�����l~w�),���L���]����Y���ڶ�)��)N~}�W������E��\��^!���뫉_��0sonLY��-qJ���q�2��̄�<ϲ���9\�ڕl�*XGFL{�wJ>��q����#�������p0}���ժ������p�\ ��0�}��g'�.�A��;�q��#MQeL	����˙�w:�=�O��0�H"T�P���%a�zc�fQ��\��s��ͿV��l]��,�Ja�F���FFǔ����P��%S��Wޥ��ԏt�,{�{(3�c~Gȉ0�":�J���{NH�����׺�3ǹ����D�":c!�<̇�e@�M���N�U�a�*b_��Oz���w9�|��f�j<'�ׅ�)�Ȩ� 9n�EB�/���
Z;���K��S�~��6���l�T^Ua��vz:�Uz��� ��g>NH��È���E�w7<�nc�5�U+ZEn�x����uVx[�`/��/�L=�җYmZV?Y�^��͟R�.��*���#l������N�c�\�j4ȼS ��T��� �*wф�`�EOm�x�c��Ѐ�2�Ѩ��-f��A�WvON�6>��E���U����2M��J1��&�V����s�3���N�CS{�cs.q��������f�W�r�D�u�e��c����Fzf���p�d�`��T9��0�g�g��E��T�Y���yU==�G�]~3\�Y�[B�Q8w�}�R\=��tA��N�s��6Q0���*#T�W�V�JPj]��)��9�#I�7��,����3;�9Ċ��=|�E��5��T+�S�k%S�
��^������#r��V�,��k���|O��Q&D�~�����Y�:�tߊ����N��ӯ\���s����>�2 0�L�'��CB��W�P�=^��f��������?�&��Ӝ}�����.Lgȁ��.t1d훸��m�/�;W�ool��UzF���=�&��@^�T�u�@�E�D�������w��n�׬w������n|O��(��鶧�W��p?	�ϴᩅ���(�R���o����>��]t��H1�'���p��1ee������,�j����`���f��'j�n�K;��6�\|��KB��#�XO<����u<}����Օ�J9$�څV�D�J���!�)ae�r^c����ov��x�F�Ŕ��h�>Q�e����z�s��yR mw2��I���U����#�N��wc��[��=0m�u����T[FSO.;i���9HV^��vN����;����n�N-%�:�K��8lO������il�saa�����T�R�V���$�Y�kS�Oc�a�*������s\챯>����o��=Ň��Ĳx麜�owo�w��#�VhUAL��U�lJ�WZ���SR��u��m�nMW�oy�����;)Y5�Ю6��)$�/"�Z~J]դP��z�D
��i�C-(�qm�AdTCX���+U�{F���q�s*wO!��\�h^��Z�p�U㓚8�P�4M�	�ܽP���d��<2e˗�˧J�8J�{o����`�od%%Xqs�1�H,���5�Ny,����wbm��Dvr0ej�\�����x�����5��9of�\ {h�bIx1]ܖ��rH��|����$�M(Q�4��F�yX_j�HL���mh�)LU���Qq�:tƴ�l<������R�fL�*�hGPdq�q�ƞFR&C�7RD$�Ż١��zm��9xZ�9���HW�4]�������8 �^;m�V$��������7��ReMIw�Dox!�`�4�c�V9�Q����q�\{�%����[��Ý��2`��D�q
oseCZ{N��̬�@u[f�\S��v�\�Q�{vؘ�7���Ӄ-,��t>�]$���{A�J9�;�M�U`&�㼂.iel}WD!v��pql��u+�@fu.���A�����|vܑ��vr�	WCW�u`����]7�:1>ҁ۔D۝8�_P��Ga�����8,�p��Ņ�6)Uմ��F �8�P�g�G���
�.+T@+E���Xa��'k���K��6�:4��5-Q� �~g�������E��9���M>�`�������쬻���(�|_v]�H�}�ʷ�n���2iˊ�����B�("��B,S\�����S��z,�v�L*�ޤu�9f��nRDǍ�� ���J��sm]��28AL�_\
*�	k5*J"��#��8��%+�(FEhj����'"�r�RI�XEX��y����tЖDD$�Źv^�
����D�CD�dZ��P��ds�v�]åNy9��S*�dS"C�.�%WD�M;�U�X��!�I
�ܚ�u�^B�m�]TV�VgN�jm�
DK��9�*�J��+�9)�����d���F�\���q ��"�ݹ9�%6$���V4L�h[\��jEEu0U	ΑUwY����J	�!$�(ŤӧNЂ�Vz,-@��B�R| EQ��c׏%J�z�W �Qκ�FvaQ���]aФ۔�M]�Ü�p�}ܝ-��br^��p$vзj:�i������~=U,r�>?S/S���?�u��f�����^��H�9���rPw��ON<J����\z�q��=�6��o�cO��`L{�hp��Yъv����U��V��#}7Łv�䋮�~�z��8�0��b﮾�u	�$+/���:b����Ӱ��������;�H�|��	�>��Q�^���t ��QU	�{8˄�c�(���茙l�a���Y�c��(;�yp����џ4%q�'�yB|��^�|��G�c���m¸��ɘ��1�҆x�=���a�*�.�}�z���|y�s��<�~�@-�o�����i�����QM����G$J�[�|�6	[�{'ߝ��̳���= r�"�*P1��.xm\���UH[�>���;
�y	Q�F�H\=��ާP�<r�%�0[ Cx�D��,Ys���u#��3kj�+�$��d+��4��5㼊�>^�a��� X�1_�5)����u�j���>��=����WS�*;��HR�՚b�v��+��Ƒˢ���@��d쫵1:Da��a��_��~\o¶|���J��G��wy�P�������w=��ww;ޭ�'4�AC���A��6\�N�Y��"܉��+��F��>��z|�y'=1��w��'�"0�/(�> '�@J����~�u9\����ѳ �����4�����R5�z���;k��#۽��"O����|M��(������1ׄ��fkK�U���GG�z�w��Ǿ�'K�U聓��h��c�s��?��n;?�qK�/V�@�g�r<0��dx�54&��b/���/�\�C���-�"H񸛟y�j�;��P�q��%M2}�,
��k%����bw�x}�s�ndz��-�z6���B��]f���~���@Nt�/�������hf���\{s�o�����L���C�W��S�>�V�V�Εi�=+���;O�����[tp�;��^����N�SIح�e�;B��9.s9!�7=u��fq>���]�9�o	�WVztV2�i��ݶ���ek��TR�=|4�.����g)P`)eA���2&�2MR6igV���=�ږp ��@��S~��ü�f*�u���z�[��n����Sa�x};��e�d	D��`Q�FE�*�a��q½�V-��r��^Bٱ��N������
��bQ*��;�0BD	n�}��@�;��㧙C}��v��\�6y����ᇄǪƉA)�ʜ��UBn��y��񬨯��*�au]n�.'��|4y<�<)ҩ��������$��Q��<$�	��# 5(a+�E�L��ݨw/��n<t��<��>�6�w�9䠼@��2C<�=?t�~�8���9�5�ǩmR!�1�<�i�3�*����T�\?m�[�*�DIcs�'lȯ'^�o��.Vnޮ��q�rLy�@��|=_3�-��>�$�܇�\[�16��8<�$�n��\��G���M�)���G�s��ʀ9�C#��PL'q����5s^|{�Ʉ7���=���[���Q��WU���3��v�׶ q��mם9wMޫm��~��^��EDd���-J����K�)��+^���l��ʺгz'��u�sVl�t�(�-~s(~O��O����bc����,�r\�Tv���J�h����І�Xp���ﳦ=W�Xo�>���@�^��L�0�䁜=3�s|��M?R��m�p���L���ӳ�[p�'�p0/ӱ����@L#L����E7�����'�[��;�+m8%R0>�CۓZ^���C8�;=��Hxu��R�uˁ'Q��q����w:n0�:�F�튨ss�,a:���rN��G�u�.����ޙgÂ����e«�wބV����G�uJo���Y�o�z��ϢWg���}�����SV�b��9iR�]��D)��;!ȒUg8oG�������N&�D��_Y��1�i����7�����{B�߿O���������^�&�ŝ�#\�<�I�'��W�x���\j�)�[��Wx��i.r}�ﯖLzǯ/���伀@l��`��̀<4.�%3W�P��|�<r�=��Fu¹��AQ)%���Y�^K7moSB5̱p�[o1�L
>���]M-�R��epz�;d���`�k�H�Z�K.������Jҍqo �=��N�:�.��[x�h6�ݭ\&Enpr=�>7��|}�86-�91p�F������\�`�Yq[��Ӻ����Ĕg�G����;.b��|M'>_�����5�A0�������P�~�|�N������1\Q,(�M"<B��>�� i��������9͕�pY�7.~~��Y%�i�wS*	���O����)��"���������W�^�����m��z�k¾�K�f�����wL"O��0�?��*&�/qgV��9�@̦$Z1�M�<�8���,x�������o�ޜ\L/-͏/q z��5�.a���>'�ܹ�;Qu�ϴ���
Ӭ����ãmzmޝz���3����f�]D��Ϟ��:ۿS|-�xhe����I���|ԁ���͔ ��a�l����^zO�GA*����wn{Ꮅ�(^������:��U�".���{�p�����h�OM ��O��04��]e���"�)ԣ[��40�*��+��*����t�Г	����Y����Ն�CV����#j6�_=�򓋴��Z���hhb����~0��H.�w�]��B�FG޷���4#Fc���q�<����?g��cQ�[�1y~|co��Io{�z'ޜ����	Tg@�L�E*�1S�l���媠dq����mߓToӇQ�r�q�׫þS�Y�@l�ǤWR$�@TG�<��;e^M[��~b�瑏l����_��.O����&�R$��cgN\b����܄����?VVL���=�=Q~��*<雅�D@��>��,��uyeo�W��,�Jy9���Oq��Ȍs�y^ߕ��:G���J��Y��r1^�  ��A�/j)�x�g�a��>�i<�Mx ��%�>̽�3��oV����{��@�s0�2����I�x|��	�]�4j��R��N��K�[a�S��<N�l� ����������*4������9���T��t(���^vc�.��B�T;�,���|�E��;Lz�6�X��?�;��g�ɮ��7w�3r����I�/.��j� u��ϛ�Ϧi���v)��̫.���F�/��˔6���f���;lɲWf�:�STh���#�����)U<�F��Ntf�i�>�h>�C���e�"{�[��/�\NT<���-{ْ���o����8ppǲ��(��Paye1"�e1p�N���
�����^������*=�z�F�}}_d�&8�.�N��W�t{�g p���{��E���,�̡����<���3��r+�c+]D��*_zD��y�}8k�:�Ң��޾��{R� ��_�T�U7��KKƝD����n�ߊ��������O��)��T����IYedF��;��S�"(�Cϰr�ףq�K-��%�<�^�ӍK�n����(*J; w�*�=�/��;qF�}Z�O�8r=������ќ[:����_�<1N
� %%:�Gt�Ufo�Y�U"�ų�>�Ʌ�u�P��z�1��������N�9~��u6v���N�F���5�2����f>ݘ}��>���b��fe@��
1�XAb���`���N���J���ˑw�|-恠(j^[GL=��T\�[f����f�N.������Fp���]��D3��f��	ѐhj�+��r��bxC<8�_Wg#N8+ܢ=n��
X@@�Z�����aY�zc�x���t�Ú��R}}8���@]�e�[�����wHNّ^R�x���Âm�My�Q�:��a����?|=�}�>&*�5��V�X�gС��g���g�.O��:j6�z��,Wܨz�<G�'4&�j ��b��3.M��s垅>���1��z{��3[P�O���d2ndGGˮ��T�.(EUs����d/}�����{�w�6r0���� �^��L��,��:dp�HS���I�e���u>��;(e�m��L����M�cyH�{_����S�HX̸��%�Fmo���X)�#t�C�2�Q�Z^����!������dױr�V�g��VV���Gy��q�GMDY�u����Un{ŋ>6��-��;9��g�Ϝ�Ie
���S*kj�}m
�]%��iե��m��'w*[*T���ous�G)tR��Onrq[�a��h|��{�v~�����c�3�^"
�c/:qA�v�3��v`��5�^lb3��1�D�5*<ܦ�.O6hv��qdVuf�(^�=s�b�F��\��
�R�i\s��H;�H1jp;�}�"�G�����U��R}P<0�����p���
��՘�5��®U�u�w6a[�#�y��-��W�6�q� ܁�"A{�G�x�0���S�t��z@�>��ǹ�.l�w�Wu�q�� ��Ñ �PЯ%3N��NG��3��֫�L�>��NRⴞ)����D;uNLZ-��\�ad�S=��>.���������S�����e�ط^$;��=��N�����������qzvWt�X����7���U>޺�3�?
�{~�zvn��{�St}jaꟻb)�I�G�}],`RwzO�|� /\)�%O���s�����H=(m|gۓ�6�+K�f�*�u�0�>/�Ɏ{W��ֆ/@Õ3�{)�����;	���us�ӡ�����D��x��;P���]�T@i�j�b�j��A.F��Fî��Hm��=������{X�&�M�w����{�ۼP��[�.J �����b��kF�u��n���t�#�W|��3���B2+��y^��a�K�τն�OY,�Ó�ա_�>�����#/��{�<;�ѧ@�L�6�v���u�M��U�~g�Y��:��ͯE��)\I�~�1�Ζ���@�_�R2�P�:luO��n;���'�$�MO�}���%��U�Dc�b�&w��r�ڑ^�_�|���Ε3
u���;��e#���-M ׀Y��m�
�r��kU����S���}��:��=cG���-<��c�%�w�b�~�P&*w��5�����(�z�m���<�q�(,=�~ӔQ���8��j�P1���~d��Y=�\�n{����Z�tǵux=&�ǽn�׌���&�R;�%�=j��%��=�P��%���YX:�U?1zQr0��:������#�j�>����Y�wG�q�|f�� ���r�t���L�p�*��l�bc��'xy�p�bb""""<ReT�I���{�R\�@UM�e��"�2�5%�'LI��Ӣ��K\�pfB�P �%��ޥ�(��ʠ �aTM-�!�yt��ֈ�,������
�t�1FF�ݍ���g�6���3}f�[�H��a�eƩ��{�Hay�����a�%b�fe�-�\2EU>���s�J�u��� 0�S�� ���pF!%hv?�W�p������O[~�S���s,���u������ ���b vXi�b4�[B�s%�h�v��#$��j@��֡3�K���9�x�9�1�yQ�月��ܢ(
�m�쀶t�Sb
�
" u�"�}�P� �.LV"!Ll2P�k8B�)��c �Y5�:�PSF�xx曛o7���� j�_t��C_�`���r��2�o3�<���#���qdTT�k.r�pz&��O�u�G҅��������k K�>���Ǒ~�׬��n[�^ǣ��M�_˳��p6��@UN��c�Ǩb���Ɏ-�hD�$���C�GUTR�Q�EU=���}��LJ��3�y��	�X|��}PUK�ΊDD���B>F#�`"�AbF���}2)�i���)�0��Q�O ���)��W��UTTɠv�;��ޜTD?E�z�|�6����	�}ڏ۰�y�3�~�(	ϷxiYc�uAB7�ճ��!<��C�mJ|w�`�~�A@UN����Mѹ#ܓ$����R;�@UI_[�Xš����������:Gp45fi{&7�'��� ��H�Z���yxl�-~@dC����{��9f�k��dPS����e�p��Mg���H:2u�oLHt�7���
�!��`m� AT��`ڃ�<��3�ÇDUN#��M�p������eq!aNtyR�.��D�|I�f������w$S�	���