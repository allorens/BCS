BZh91AY&SYpc�r_�py����߰����  aS��    � 
             �                    �)�	R(�(UP@��>�l �� 	((�
P�J����k�7vW�^�Z�Y�C�n���b�f������S�  @|��SYHowE]e9��;Ժ�m�eR��ݚm�:��vn�vȎuuT��T����eە!NF�� P t V�糪���{MVŵ�E����ha���+FZUEEl�ÍT���  0�>p㯮��s\�]
�=h���b�V`ǗNR��R�6J%)P d ��
O�ܥ
/iR(-�
o��D���`�S��m����N�ld�һh �=<����j��Xq�[�#m���'g��Җ���	,����P � �ͩR�������vD:V�T���:�EAM4[P�k�^���  �|�u�iR��q�wr���j֡R��ݬEX�b� H 'PS}�@��1"��W`c����6ڭk������z�l�Jl i�Ov[�(q�f�ձ��-��[iLr��V�a�,�C/v:�                        @  � P���~�T��      S�%J����`2h�"{J��@ 4   4   	S�)�R4�a M4��&��
���	4�0���	���zFF�<�P��R��I��d    ��Ϯ��q*�����}��s�}渚͇�Ӳۚ~�ӱ�����3}1��}��|_WFٛ�x����~���ϯ���WoS���wK���©@�F�6f�ۨ�Lu��q�U_-�;�fl?��Vg�F�ŷYUUUQ���V;|s7�~d�O��O���pʙE���Q���y��r�ֵ��Z���mke�]M�kq�&mm-��Sm�kn�V�ֶ���ֵ��O��k���Zܩ��kZ��Z�=YkZ�z��k���w-)�ֶV�e����J͵kJ�[+�j\in-ki�Kl.0�)Ki*��Kmm;��u������i�ŭl:����V�֖"��ַ�R�֕��Z�Z�n-l�۵��Vź�����Eź�ַo-l�-kiեV�ֶ�R�+ZV����Zmn��:۬;fN�Vեis�J��R�ZZ��l��۫-kS�����q�Z�i�qKak0��k[�-;Zֵ�n�jel�V�����Ŷ�RY�ZԵ���ַZr��R�kZִ�n���mŭku�.&miZ���6�V�m�58Zֶ�2����8Zָ�۫[����ַ�;iZv����m�i[�jeka��56�����+ekc�m�����q����ֵ������qLE����qN-j[Zֵ�kZַ-kakUM�kZܹ�T��kZֶ��ne+ekc�kakM����2������ĭki�ŭk[mZֶ�[6��ĭ|Jֵ�եkZӆ�+Zֵ�Ű����kn-k[������+mk[L���Kbַ4�V��Ҧֶ56˫J�\qn-kgSm-kmx�m�kR�ꖵ�1<Zֲ�<Z�ˎZ���ֵ���V�-kZ��72��m9kRה��Z��ݷT�V��km�ŭkZ׹�-e2�Zֵ���)Zֶ�2������U�kZݷT�ؙ��k[v▶ŭkikr�)Kik[v��ekM��ֵ������mk[K�Zֶ36���Ê��Zֵ�+Z֜M���-ź�:��k[�ڛqM���f{:gs����4�a�#�
�
=O<8|�Ͱ�f%�⺵�p�OV��u�V��mkZ��̭k[���k[��Zֵ�t�𲵖�&������ֶ�6����Z��+�ږ���ͭl��s�XZ־OV�*[������+ml-y�Z��kR�ekZי��k[��Z�ZV�ݵ��aV��m�-ՙYz�Z��k�ak,�K�-j���ZV���l���ֶ�Z�ml-k_&�ۍ^�KZ��̭եlZֵ��qkek_gv�i��x������_&7����K��W��W��K��.F�3n�kv�aI\.-j[��kan7s��������j[�ng78Qe�r�-l/S�]��-�T�'�
E���4�|(�X�ф�H��m���n0�M��/�ki��Zש��w;R����6��6�)�D���I[�����e.٢�����-l-��m�ݺ�a]�ө��[�n�kWRى[	Zӹ��q��+�Ji{�R�\ͺ�W��R�[�������Z�4������e����6�\�ӎ/3����Yeq�֫��Z�ɵ��M�l�sl-j��KJ�6Z�_f�aq��^�ֶ���u6���ږ�jmkmz�U-kn%�����ש����-m.fֶ�s�-�ͭl/�ݭ�뭲ː���يZ��&ԷWS��i��ֵ��-kai���ek[��Z��Ÿ��n�l����3ZakZ�v֥�kg3kZ��w1+Z�떥���ͭkZ�����+fֵ��w2����mkZ�U�խn۪Z��s6��n��^y���<�mL馢�U��Zֶ][k�V�+��ֵ�g�ZˍM�kiqkZַx�-��y�Zֶ�ekZ�ɵ���*mlZ־Ͷ�ֽM�kSM����������M�+qkq��R���6��k��֫-{�Z�qs6��k���k^fֵ���Zֵ�ml-k���km}�a��K��ֶ�.�:��j^�ֵ���k�ZֶY_R���M�n���6����W=Rֵ���T��f�Zص�����V��Zֵ�ٵ-��j��ֵ��̺��j���Zܩ���kO&ֶb��ֽNV����Zֵ��#�.9��rmn3sTZ�6��ɲܹ���*���sj[���V�&���m���M��ݩ�j[��ۋew6�T�#kmmfr�V��:Z��ť����en��ͭkk����bֵ.�jim�s|�3K��Wq|��m��Zֵ�q��������ki�ŭkk3m���13��kZ����aq3kZֵ�3+Z�Zө��m0�%3;cS�ͭ�ˍ���m�����F�{�Lx�' Lh�]b�a�e�ZYj2�*��ղŴ�Ɩ�[�7kiܭ]�i�Ʀ��ڝ[�����M�������m������+Z�6��%��SZ�9eu4�R��ɥ�zm�u���[�s�S�;�݋u������e�2��-�6M���j�[Ku���a���k[�f�.���3.���E�sKRһ����R�k[k��V�1s+[�g3,��͸���M0��6�ש��}�p��ֵ�mkf.eq+^&���_f��Kf����3m-m�-�V�M������[�7����֮Ͳ��cjV���6��_&��ŭk��kS72���+Zי�,���p�fmk[�q���3Kq��b�[+fg=R�a����+Z��۫Jֶܹ�Z�[v����6�����ͭl�Ŵ��l����V�+Zu6����keխj���Zҷjm�-k�qe���k[L�s.�,�kr-���l�k[���kf�Yki��k��k[J��kqn�֕0��ֵ��[�ZԶ��l�1=qkZ�vҵ�+[<Rֵ�Ĭ����[i6��Z��V����ikZ�n-n-���M�k[m��f�[K]�T��Z����Z�]NZ���6��2��Ͱ������Z�Ë[L.;6��6��n-Ŷ�ٵ�kh����-kZݵ�ŭMZֶ]Z�N0����k[--�Z�[+i|J�[��kmk�m����mm2庳�0�V��iZֶWJQn�je�V���ml%յ�5kc���������[�/�/M4`�mjZ�r�[K�-�U����r�Z�u�L�T��b�ŭn�n�+v:�V�:�nejf��ڭ�4���ne��gM4�ڶ��Fm�Ka�����F��6�\����V�k��n-�[��v�1�X�FXM-�i��ܭŸ��s6��܇#in���O]mk�V������9kR�Kqk^��Jˋmj����ml�Ml��m��g��6��m}��猯�8�.3[eirҴ���qI��[Xelel%m�ήi,)VZ���Z�qqKZ���mml2�ͲaN�f\.&g+,�M�j��h�.Ɩ���ͭ�u1+-lbe���ֶWs��u�nx����J־Ͷ���Zչ����ʖ���+mm��jm��e*Z׉�V��L[�-���b-|�am5S��k_&���q�)y�Z�q|�u�b�Y{�ZٹҖ���KfWٵ-m��j���۫u����ܙ�V�+fV��̱s+Z�Z�n�m��M�kgk[�:J�Yknֶ���V��mnmkeƖղ����s--l�i��kZ��Z�Z�����%k[��Z���-ŭl���֦.ekZ�[k��[K-�Zֶ�=R�Z�:�ֵ�ړ3kuk^����Z�6�+[Kr�V�Kuz�Zֶ�mkZ��[Z�Ŵ��q�ֵ��[�K+�cs3]���X����+�2���Կ��_��|Y}_WO���o��J��+����n{g�<�ݖ�"Z��U��m�&�`{�uhi��m��	��&cd�!��a"�Ht�e#���^�cd�NiP�xt޷ծ<=��A��V�	:S�S�n����d��j0oP�V��H�s�>��S/_��U�ݸ{��2��eZʝ�/~6_���o��|���6�ޔ�҂K1����eĄ�IX�Z����jz�hf�Ĺ���t�J�%L�t�[���(��k�)������fy���y���2(U�	FHL��gc�氵�"�t�-.wf��sI�������;�J>Ho��f��/~;��^�<��f�C]���TEcn�_-�|@�&)�=�'s�sf�\V�p慀������Y�t���:X�f����I������1Y�ȭ�YD
oݙi$��1Ս�=&��¶�� 1[܃CF�X�O#g
�6�y�i
Y�c��tME��ҍ9��nI!6�-��*<oJ{[Z�=4�B�������ZQ�[����m���wfu�?9^�6VA��*��&$�,��gNdңe�f֖x�?�a<�0�d2Fi!]��q��VC�D-��V�VKr��"�;g&��gKZ���w˷6�I�Bo�	^k'ǘ+A�ic<;i�*Ǐ7�3/K7���C��+
%��g�]��OHo�m~��'n��z "b�pd��~���t����Δp��&��a4R$���z��Jݲ��>�"쵎㵷[Sӭ�>�i�lkgoJ;k�Ae)��)a��w5��%��GN�u����4õ秱J@ɏq��9�0�J��׾�z_�6{�ܮ4{�1�7��ˉ]R�^ ���5��u�H}0�ѳǋ�צ�cfa]0��1�Љ��/=0��OIP���t��ǢucG�+Y/5�NY�:�N���c�-˕�̐���A�̆S��xZ�[�g&	��2y�����l���!�r�oc7�J$��X�&��zuy�ǧ�:ݎiV��]x@e��\�]�C�B(���߽ste��&�k��5���7���l���^e�ӑ�[�N_�H�9&��i����"yi����G%�9�ҡ������%Ʊ��TJ����ng�E�4��fY$�I���@�,��.�a��[<W��;J3��a,��0�OO ej��k|p��O%������V�h����p�Y0�����<����[�:�]�vi���փ�r���@F��	�_�!��Ǜ�٧�ZY\d���V���jx�I�p�zx�%���45��.��,���:Ő�:|B��'��;Lp�e㇦��<��I.鐋Lx�~ ?\z�^2J���!�z'au�E�Sʎ)�gfN�ò��Y������UB^����N�8f6O<G������&t�]��u�}t�ø�~ C��4��M�|	�H�:e��fL(x������ϼ{���7��I�����V����!�q�-o|rk�����E���75Ή����9���R&�C2u��2�Dv���{��.�XL�j;��9P���9����?6r� "I���$��O��yú�|D$UN�R��:��\��� �����^90�,T� aEk����r�C�8|p�gXt��y�M i��<�l�Q>z�$
f�H�0�=��&�	��x@ێt�u4YG������Hg��	�(���gOe'���z2�2v�<�i��&<�q�ҷ�i�yzބ�s:���8|���M>��������a�;9�8Ie�,���M9?n�h����Ӹ/B]Aa�C�,$����0dE��E`{3r����Ҟ����{�ߨ�I����ՙ�2wOK=���ަ�W���
�/|љ�<)��]�z��x��Z�{t�b�,��4�V)����f�M>�Xr�r�}3v�b1����0���z�/&t�v831�#2��y2�F�v�iO��3����z���'�\5���*+�)�NB:�G��=n"��t�Ev���W���@�Q��uᥞq��n.	��ˇ5��tnl��X�����ONLVåΜ;���<t���G�M�/Ι�*4�'��EUk��w��G,�{�y7�	����p�a�F� ��_�x�V�Q���˯��ܴ��&Lhy<ۗL8�,�ݔ���V��aF�������r��O���W��%5u�ҡDpԷ�K:zw*k�l��X��#sG��T!�suuz)N0�|�j~�ʯu�-�1st��&d
��G=�a�>�zS����5C�M8�w�����~4�w����z�m2>��r�t��[;��}�p��ѥ�9�&���(�j���X����fr��h~����c���
%��4q1��os���z�u���zvt�[���>�F:]o��v}�Q7�Ǎ=��SBb�Z�#�5�������%�}�\���v��I�c^S7	��[ss)<�'�--H�rѺFB���$q�7\74�7i���(مx��������u�TDqc���h]T���Q�蕇��
U�p��f婶I��&����d���k���A��a��>":K���H|���B^:z�w��q�����X홏0�J��Ψq�C_Ow����Fz#t�8���OJ��G�OI?�7׸Q8s
��k�r���E1��x�����<�+c�����C��Ο�'=FŇp/��pɤ�)�S^���R4�V�<�{6떿b��{z����-�&�l�LVj#P�rS�ݴ��G����3f�d�r����pw�ܾy��vh�g��z�m0�zt�����4��I�t��9��x�h��B�}��":�IÆ��>�Ow�LW��b�Y��׼�	�1�<}0�Ius͗�ǳ��`^���j/���y�9�Wz�t&a��_���I�/<���L�"��:��=��Ozٺ����[4��zb,��M�3)�l�{��f��Z��vhI�S��u�{^F֐�{5��u�DDt�u{<2$h��N�>�L'w���#�bıˬ���X��x�p���9	�����q����_{������U����_	��[7���O2:!J�k~U�O�v�!5kei��!�:��.��כ�f>�!∜&({:@�wmY=���g�
b���e�E N�q�ٓ��<øM��;��v��r_vf6'�%�i�*u�Ǌ�@��8S;����Y�����;�ξ�!�y�0�$�c}��ֻ���{�Ϗ���7_gK�J3�a�o:DF���	����{״��L�l�K:Y�����}��si̝������i�����s	}:���"G�̍X��x�g-�vwrâ�p�Ů�e�}ُ�y�8���C����?�5t����@�A�f.��0��k��o.��<,�{Ҥ)��Ḽ���ɐ�GO6A��$3Վ�=z��ۣ�MoIh��S�DÝ9�s�0��C/w��B���RJ��>v6�e�.wn<Ff6��T�t�r� rkx��wFbe��)��dg����k�t�fbұ�g���I�J]�y��}����J�㈳�<[�I��1!6£�x���d��lP�e�c�yh�뇥/4<�B�Α�ݯD{{����11W�go[ݮx������M���3����*�����|}ޑ���Xw}:w�'�V�d�rתz nI��tvB{�w�����=�}6Lɴ\[X�״���U���A�C�{�x��=�����MKm�aG�������7�7�Mp�W��� �uG�WL�x�Y����[&�O؎exn�����ˤ�=]}�a�tjXMF��28z�Gf��H�ql��~��<T�P=�ޘ*���A#�srV�z|I�g����e9��go�����z�r���ٵ�&��<�T�ް�_�^�������x��}�O�>�?�����d���>���q������������A)?�?�?Í{O���-��Ysm�7j_Og���uu��s�U�6�t��q�\Q�}�vuՒZ�)4�B�X�������珻�t�S�A�؞��^��m��;vp��s��Z��/����ֲXnhg���Ü��gv��an��8�Һ���v�kR�V\$GNe���`�I(�t��ە{��;�7?|o�M��J4�U�����c��ǽ`ڔ�S9��!�+��<�ݼ���
�q���o?^M�ox�k���(�S��ܒs[��<G�k~��oIș�M��y���`Z,���m��B�V�4u+s8�W���K�̦]i6Q����3�f��f�+o!�MX���c?,^p7E���js̖��R�#1��r����u��q���^6޳z<>o�!�K�e��=�5��E��K['{���f�bh�mD��^��m�댗�u�s̜�N/Y!k���uZ���&�i\\Bi�IGUe٭ua䜛*����Ι�\��+�t���6����Ws�{X��Lqf��t�UCpʊs�-��q�ƻOG:x=z-囜K�g����5�Z{G{W�t�uh��^�><�����M�E�a.ك`���ˑ�-�ٓS$�Y^����Y����$��ɵ�Ns��-`�ԕ�����L��<�ǋɛ	5ƫ
»%)E�2�����,�w%�$��Ӝ~�vȓ��m!+#�1�	��ԑ@��>C������)"Il�HJ��D����]h�J�il2N⽝I����Oh�&3�j�]K�?���Vz�՜�9�.��]I]7�ڙk.��i[Ć$#^Uk	��:�|N��[�k���ݕ'{т)R�t`�D��Rl�
I��m��{�7]]V�&�)6%#��ڗ��ʝbQ9���kN(��.{�n52>���i���D.s�}X�I����$8�ݹwo��i�{��i
����#%�$��c �--X�M)a,��W��d�.-�Z�t�Ms̸��t2֓<�qqy4�a9ώ��^��\�^$cM&�hyk�F��^���ށS�м�9ŜͪW�$��C]`6s��]mEj:p�FA��e�9Jۗ�dP��m�F�^p�x�_3;)�M�>%�4���#��:s�ԔS�ּu� �{8�mFha���:���9<)�o`$��m�]+�K�v��Ki;�L���'^+���Ik�Ԯ�YI��9���#�9��8g� �z�z�^s�8鶡P�ӓ漯;�䓳�qb-��+��^s�
z�B�qys�?!��G�y�?D�H�NT�4���!��P�#��!dq�����E?pR0� �Ų(=��|���co��k躩�{��fm���v������_���V���y~��-������o������+V�յ7�n,�ƖجZ�9m��o��:�q����f��ת�U]y���}�{����������x���8vǀ�6�C��� ðhR��P ���{���0v�  �@/��]W��]u�h6Vه&�f�՛6������GV�(�BR��%150L̓Y]�.�ww���q@-�F�g@�@; c�< ��t@�x��^����@�4��pv�K���.LT�H0�LAɄ&܆�F��ն�S�{w��� ��  ��4��a������`c;:� p�� X�Zִ�: ð<�]����ww��!3L��L�&Y�;��V�c�ڝ��kME�qۜ�k�m̅m�շ-��8덮���B����J%J��ɨ)E+R�V��
���-���R���V|~?O��o�l̈́֨���������6ޟ�����4���~����Z�um���a����������-k[+Z�q�8�m�����kZ��֦����L-kYkm��l-kZֶ㮭m�k[n��-kikZִ�k[e��ź���km%�J�-iZַV�ֶ��kikZ�Jֵ��-k[�ikZ�Z����M-�����)e���l4�-km�������[�R�a����kZ��,���l)kZ����-�]u�V▵-l�kZ�miZ�������[��պ�*p�IYl%g���V����Z���VZ��ֵ-n�+Z�Zҷ�|����{�= ��K*C�4#���f\"\�"�ck)�Wi�fÆ��B��;�S��I�s�v�Y��`��A��v�٪-�r�r��W6����Kg��}�}���Μ���!h�g]�w[��x��D�8�Y�)8M]ɮ�G���ԃ{���v+m�t�"X�R�-!�$��ϙc���҆h��\��׭���M���F՜��綇��teCS��kg��C��g�͔��<����C]x��y9R�-s�xc;�~_�����+���l}���g���L�����\��Y�����ۥE�˵�gTĬ�c
זKSf¤q�{u�I��U�,r.$ܜ��sc1��Gd���Ǝ�^�<t�p�p8��`���ҏ]�+aHkul)�2�m4��
�gG�����y�ՠ5��bi{8&�ۭ�
M��3�/���7]%�nՂ�n/F�j|B%�qZ�ucOhG�(Z���tsb\�D�6Mm�Z)YZCeW�b���8�㦢b:�v�� 닣��V��u�����{9-���;��ے���cF-���ۊXHD�i)ޘ[$��:�����6���~��cZ���v�2��v��';5��]l:U��)n����]#f��j�V�e��s��(�:B6�������OV�EY�
�O/�6��h�Ӵq�4�>2�F����/qsZ=��y�<=Api|r�IX�k��l��"v�N�MC��l{0�٭=���<��ѱ�ͮ8s��i��f��8��Q{盔J��[�5�e([�T,�t:�E#�p�nvӓ�Zn]Zm���P\�]fv���n���N�n6��y�8��pWi��Fnb���VRYJ��&�x(�͏	�W��sۑ��a�tK�mv6�,�g�O�nv�r��0w`��I��n���D�Yu��Q�*���Z�EgXn�:VZ;==���0S�S�wb�=�ݓ�������*Rn ݘ�E�R&�۰|�ӏc�,��].�a��Et�,u13��F��mz<���j3��LU�J��.��Cs2jv��e�pk�6�ٹܛ:���u���/d�]&ǩ8��6e�qם�G3��ؼtj�%��+��C,vݻGj��:3��t����ZE�f��>6�8����8o"v��%�8����8K�m��S]���kF�W.������h���◲�ɮ!1� ��\�|v��������a�6�O*Mk��!��ۇ���Ts����u�Q�/o���\�T=���a���@�q���8E�oIm����˷N�%�B;���w�����sz�5� ����u$34���窪��RI�:�w}�sz�5�"8��8�̭�\mn�����Z�Zַډi�d>����olܗL.�&n��YE+��,�:}��nN���L�aUqF��U��}Le�e�7;\���vl�l�@`�1�d1ƌ�i���H"��򘖬�����6�(�&`�6��e�]����S�Zڞ��8���*��d[��S����1e��YiSv��4�7c\��mÇ�l�v�����9،I��&�R#��F9�cX,G�i�pwC�^��{.l�x܊���v{i.b�}M�!,
$�`�������x�#z¿K����N�x�F������1�~;k��hVo.G�)Y�b-I�m۬K}�J�ډ��G����T�јҔ�%3O4�c)�GꘄL�b��(('�{�a/����4:@�/���jˊ8����rßc�Х��~�K�"��52�`���H�����)`�F�����ISi�"p��4�(��R������z�=��Od��rޟ��er����!��@ۗ��^��[2�y��q�m�^J�um�n�k[�mD���u�µ��EK�<�U9��������2���qm`�6�g�iI�[����Η�Nے��ZU��g�����߲�^��:}��y��"�}:Sm/w�-�[M9=�7:����$���"�y�{�{�|�>q:!�Ԓ|#�44��@ P��G�0Q�N)�׷�iy��Rf���[�Ų£�i��iո��ZV�mkukZ�[j%�Xe��nH�2��&Ԫ��x�nJ�L�ڳ�9ڪ;����اQ3/)�h�c��2�@ ?�9�|�|�x�|�ȯuْ֙�6���a�&X������"چ��^H�������rF;M�l�`q���px<��V�Ͼ�Ђ�6!��l�����Cy���D� �C/,��Uh�:w���W|�	��T����yS5��h�ew3Qǣ1��<�0��[�8ۮ�+uն����oO���c����:����T�c���I�.0�?����:<�{���{�y��	_bxڢ�2����%$O�p}h%���a$A�t|�VH� xPtRf6z�e�jYq�I,�b99��/���RL���t��`�A�s9�0:< ��﹄�[l���^R��l�I�����F\�OTGV��x��\�g,c>:�a*rx�������ZqO՗�o>[����mkukZ�[j%�Xe����ɥ()�ց���p�%��!��E�c]���`�m��4�i��&Y���i���K���p��fJj�
�X���m$K�� J�rnźbK��{g'bh�Fwlh�ڵ�-}�۹rȩ8��Qq�٫�¥����������Ί�|�{(�8R8�%ry��|��Q)��y����T���aG�~���{5x�D.Fk���LZz�%�0QP�D�V��������1��yI�xE�IObNTq��+u��fU�a2���!)�\vޜ��kMeJa�y3�RoX�R�i;.�q�c(��a0�;*�/8�"�L7[��2�J*%���C�!���,R��	%�ntƌ^�υ�ݺ�x'��<�<)9��3���l�j��8��)Ɠq��K��8۫Yn��ַV��Ŷ��1L`�}���PP��Nqs0��733'"b7�Ɲ�t�r4�/)�M�f�nmm�q���w�;3�fLo�r��M�o���!χ�xG
]����>|6F��^����������?��q�ç�n�elCKK�6m���/�<�<�G��Q�'FA�4�>c'qO��(�^���J�S�6�a����&g]^1�R�'i[6�]y��Z֗][k[�ukqm���a�N�Z�̩^EQ;�P����c�s����1�UMb�a�G�)���E�B98�%��6��a��r9*q3t�����
��Kq�³�G$��>�<}ҷh;m�Vk�@����>6 �.�d�ѯ:=�`<Z��3H��}����#+�3XĚ�;2�%����To����g��.�8S�G&x(�'9O!y���'b��G�)�zg,�,L��14��Ï-o8��Z��mkun�n-��,2��ﶚ�nffILng�'js��sU��2�/V�{���"����un%�2��7��b�Uw֬��r��[�o�te��j�),$��,T���������'&8f>���k��&��-�����sI����L�F����,Ĭ���2���BW��V��U�uZP��O7=���,3�=�UO���z��C�U��,���]d�4��EG{檪q�a5��e5�0���	vg�N�ڋULV؉��Z")�[:��m�iuն���]m֔K,��'�L��籎��bA�ܑ;�y��Eo�G����l��N@�`<g�g}˜yQ���|o�|7�����9��@���]��������4/EL���٧u!�c�1$�&|p�e�q��!ΰ��B��-�4����lVD�ǆ[��B�v�S����id��nixd۷C�1��4v0xƁ�ތ�1C��sI���1��s�!��Ej*5��9�D��aU��L	��Xn��,�<*=:<���q��S�a9�Oy���bx�i,���Q^S�8ħLSͱ.q�Z���y��� L�#�R��i��
�D���-,��/�<op�qٚ��s�m�ϥ�%�K){:������{������}.����30mL��1�a�)Ժʳ>S^&ZL����yʄ�1m��8�y�.��ַV뭺҉e�d���IS32�j��)��Z�x���`�7SV��餢 e�\8O�σ鸇���a=)��7��_I��2�'�B���>i�˱P��;ĞG���r��3�M�ON<9�5ė����1┵7b"	&��E����GA���[n�q�X]�KR�1|�<=�y�:C�t�0`|�lo4�3��.F��I�Zp�CiL��1^�"��y�}���S4�)�e֕����V�8��Sj�1���1���K��j��1��ǘ��םcO�|��Ly�y�u=OYWWT���8�<�<�<�<�-^R��<�<��<�<�)�<O���~1��y�|���J|�^U�V�U��ZqV��YZ���>W�y�R��=S1���y�u�:�O���>r�T�O1)�e�<�y^����y8O�{�u9��y^y^O�y�<���2�eQ�����y�[���1���y�<�ҴҼڶ¼��K
�XyR�&^��M<ǒ�p¼y^y^'));KɔǓ��:N^)��ʉy�<�<��-+ɗ����|�yN&�W�)�p�����/1����[Ϙ��y�[�<�<�>|��<�<�O�Ǟc�V��<�W����y<q�#��V�O�O�s3��:�O�+�Ǔm0�9R�38y\y^m^K����+�W��2ڼ�)^O�W�W�2�����|�_:��Tϔ����&�=}�Fq�F�т;��O憤!҃Ho#�1����}k^uw�\Y8�AD�� �7���/&�!^��IH�{6�/���qf�0A~iJk��i��u��T^��\6Ӕm��<ȸ�HF�̹�˨s���|x�I�K�i�m>x���W,B� Q�j�����xzcXK�[gHK��G�Jq�ј����/��O>��?{ߍ٭k��^�k^�fq�{I�rIw��wꪤ�{�w$�fs�.�W~�Ԓ\���Is$��;� y��yku�\[�<����[�u��y��)��i��9��UJ�Q#h����㺝�oZԸG�ʏ�De1�T����Dn�iUJ����u��tXyӚnɝ2��Nx�U����Ͷs
�d��腛���ܹsV�Y�g-�=���J�e�o:y�&$���H��)7��X�M�-�n���	��n�~cH���sg=�vN��7KiӤ-a ���>J��>�v�-Θe�s����۴�G�0����eP�O�3�����$��������3��v�qlw�xtZQ��F�jM����,&�|��g�[o;ی�\�Gd�nk7�^]7��;��ѸXKr�翎�4��x<N�D�N?���w��I����5���wU�7{7��l>j)%�"�RfMʦĢr��IO��1�aTӎAH�$f"`�=���t����SyX�x҈���!Q% ��yo�8�-n�խn:ۏ:���M4�L�^׆��Ü�'����m�[ٚi>1�������/N��[˙������q�m͙��{Í�g�=�ֱ�7sqs�!��O��$b��6ko5�C���D)�d.H��a8 ��w���6��EH��5���qH(��!F����C���G|�w��1ʁ���?%T�3��%]�� �FLe<�2$��a��6��L��n%
K�a-��l��zs�u��T��P�S�*!Iq(���d����ͯ~3������C����Ny���X��}���ؑ����x�ӏ	��vv��ΰ�F�N#	��/��^=��\$e1&$T��v=�"���X@����N��y[r#��,:�\�i�t�I���0&%�m��-�uo�yj[ͼ�q��i�`��a���U�V��.8u,u"He�	�#k��J��3II_���8F��k`�y�G�Y&n�2_'%��"��Ĝ��xG�s.�V=M�S�6�!᥵�Z�f���7]w
�]�0����;JF�$^�(�{MRV|~Wp�'cr.�0��hA��^�󢾎�ޣ���0����%f��ZF���P9wk�a�8���|]��z[���)8�|ƚ��&$�	��xG��{#��[{i�L& ������I�LH�'�b���x�͓υ�ߗ9��7��y��𞹸����<����]\�/F�l�#U�(��#�,�&��8������;ZtP���y$S�m�lR%-���*"'���*���Cd��i�3����$[T��fq���ZQKl�C�k�{�u��:zwu�d�җ�U�t52�MD���#>��������|a9�C�ۧ]�L�6���f��7�E�̶��]��DbG���������'��6NKRQ��r���l[�Jfw���A��~+��|e���~x(I����s�S��-8��n`[�3�&TH����5<����%����7UU[ˉF夊�e��F��2��V�:��<�-��yלu�Zy)��i��<�u�ᷜQPx� z"�?y];����<�.�4��a�U�D*Y$f&"1(�v汍���7��[<b!��%�R:H��Q��pw��>.N�����M�7Ƙ�E3�T�IEmQ%�����'x᷄{���5Ӎ���<�{��E(��F������%m�#䘉Gx��刃m�#��o�4�w,�t�p�gnn�\K�Q��\S��O��L��x"'= @?p��-���2��/$��Ëè�=�X[$E�p��Ș�U$R����8 >���	lR=�}Z[��UG��F�
&"5#@KL�EW�2�d�*FX�j$µ����a#qkq�s&#	n$�b9\Nk��)��]L,�!����ȝ�9��շ��.\��='�����-���1K)b`����8��y�o8�μ㭺���4�2t���<��~B?W�'>����-�^�j2>J��_99��|�bO�8�#IwW]�*��5TQ#I<����"�M��Y�ؘFe(r%D�F�R�#9����Te!�>;�n�����D9ޯ�:<�892��N��C�c�����O=;���ڭ��^\|ko:�9#q1��DC�FY���E+s��O�c.�a�VҫRU�Ų^�J����X$.,A4P�x��)��-&�S�1���J��%�(��C�6F!�;KL)��ڹ�LҪS��YTE�3Ų�"7*�&)Q%�:�8�#l�n�e~��c:00��)c�۪�F �0�K���5���:έ����f�ʮ�N�ݖ�)0��TC(��J�;O�j⫭�đkfw��=h��ͷ�eH��TOX��J�i��G��G���Ϟy����|��R�q�y�[|�1D�,�]��"��N�)J�74�.�<�.�;NX�pO�������v̛]�G��zC�4���e�l�i=!��s�ⱊ�gC1L�
�3D��~9�,��J�5�"%�U;�=��)$埼��o��9�'> <��jwt���N:[�dt[4�!| >��/�_�mƿ
Y�`#R���nu���4�h�~�����YL��c��nFf!�JV�i���h����79�vvX��Ǥ��c�nOt����<�a�a �yO_�)� �x��&#��+��Ф�1�F����	�iFq3p�.0���ËSr�&$���}��T#q��w?*�LDm1"��[LF�/qP�1䴉�)faIFT4q/$�yռ����<�-�yo8�n��Q��:8{;I}�Ԩɲ��uϳ1@�bb?�#]��Q�v,&<��h��D�O�X�R1 ^����c;o���X����W�[L����<c��&a��4�5���Ǽ�T;�����7؛QיD����K!˫� &�Z\+�蕓�A�K	�l���n�.?10#K{뽗Ye)���I�	�U^��춓>&��vt���xu����]:ǄD=���\��u�(�b<�Ƹ�:��'}N]����O>������}����;�ۚN�&���eժ#�J�L)0'�IF`��79�	ï������8�ZN|����a�I0��Lý'=�9�s���8��?;���%���6�bb�����R�a0u1�%��K'y���9Aq��F<��&��R��L3�oɮ�}t��ZQQi�FGX�H�����/-)�LP�y~�Z���0��a8�f�Y���?h8+���y�^"th< ���	m)ʠ������LL���M��)LG��7���c=��5}�u��"0E���n4�����o<���<��u�Zy��Ji�Zh�3�V8���{JTY���N�㽻m�7�*�RgS4��Jil71�d�o�^nst;,�dr�q�H�m��y��g8�.7	��G��a�(����#q&�{�52���S:�tz��1�=��,y��-;;��[���-��ˍ�[��[J�3���T�fQJ.�(Q#�}�o�sN�����m�����<� �'�~��i�F�Y3�N�����4����y�8D�e�(�LDe0ļ�:9N�j#��Bb1U^&z����s��=ݳ�o$�u�sG	����n�{�w�}񹵧�+�<��%(��_'��0��9�CI�Z]a�D�LB���Ii�m���q��y��y�ӭ���%*i��t�|?W����K�G�Cӣ�Qd���]���&!��UW�m0���D�jjT�7�2�(���=0ur�a'��g�e�0�:���fGb]m�}Xz'!C�8�
!�����;<-����u��X�ӳӭ���wښ��c�m+��nہ�AT�#�8O��a�q`��b�!W�dF��$��N��h|zq�[=D���^k����;������3��f�L>�o�d}1%���t��DH�(�ZI���t��Γ�Im��t���xc�����ԡ��D�Ľ�>�m�Z!��Zni�޸=��u��=���M��׿�����!���91K,ki�>K2�K.�f)�`���!o�mź����yky��yo2�n��	R�a�h�ػ�KJ�ɧ:�L������ŝ��g�:ܹt<{�Y�M�"��g�#�Ȩa%9٨�Zb5+��e��j��:���Lh��=�s��N@@�ޒ?[��\7�J�7Ydڻ�����_M�3;�iZb%%�f�3(�ô�0�;��_F����D�J��
��瓛N��(�I��`���L�%������wÛnz)͢k;'��Y��X�1\�'�D�'Ϣ�%�����S�bTLBW���V��
c3:`��$i'ľ�)kɦ�]�D=��.kۘ�{��û����|���2�d4���I��{���|x���v��)��)*&�aIfbI}�x�E&�2�?��~Z��?'ɶ���\y^Z�ӌe��O�i�<�'��c�V�V�y^m�<��W]W\V�q�'�+l���+���������i�y�y>N�W�W���e�<�6�SΩו��Ҽ�R����kW[W�+βǞV^W�SΫ���y>eOL��L�⼵Z|���x�9S1O*^T����4򼗓�����u�y�q:���y>q^O�Ǟc������m1�������|�<�<�<�y�O��զ��ͱO+��a8O�y��|�����r�'	�?)_>W˺�Rx^�Ou��u�Ҟꗕו��.�-+��|Ï3��6�[�%6�&�y�'�4ǞW�['a�u]z��o����4��W�y�<���u9yO'<Ǔ���y;q�O�����^Z���p�qZO�U%��Ky�)^N���i�y>N�y�%O*�V�O)/+�+<Ɠ�����cǕ���y��>c�O|+��huDs#���q~5�>8e��D?��c�,�ZE%��=є���aڢ������1MCr5%� ;�`8�l�ˊ�)�ͮ-�[�T��rT��.���INlޝ�����K̍@��u`L�3�hU�/�2 ��Da����V!��$[1��[Q�I�%*�
Hen�R��c[Bhz�#\�����`|H �F���
�d.��d!ff̑	7fO��1����n�iE&��ju!/B�vXp^ξ��>oz7҉^���zu���e��×�X����I�y&�0��D���c�r��5k�XVţ\K)-p̆�X���1 �Oȩ��B6�e�ܖ�j�cB2�/mp���L�:4L=p�ņ5�6a9r���0�3�f� �����O��29	�X���
�3+̘[�ə���L��	Fmh������淢���J4�1�ՖE��Y
��<�(ӂ�a��5�)����PF#őѫ(�@����a�Bi�#���F\�;A��Gq��m�������j�d�t���*��G��n��V�N�8)ru؂�]1�ՓW[�CN٣�zƒ���[�13I+p���Z���᠄���]���7���=v�Ԟ�AsWF�L֦�ZF)��rĆ��j
�;d�^�n%Qv�7�E���LD)(��T��1����[}�ﾻr岻33�5��(ծۯ�.l\�R�U���:H�Z��������k�;��I�Iwz��RIrN�fjK��ܒnI<�jK��ߪ�R�R�Z��yku���:����ij$!ҝ)ӡ���ɟ�sǛ3i	sZ-��꥔�J9֫[,�k@�iDv��;��ے\$���nI���o�Ilؼ�ٌ�pv�\���;����V�E�a�t5�!�k�)�q���B�ѻ�X�K��2Fj]�j%m�^QE*�bL���:S;�����A����"�ی�,k��\غ볕�])vsx�XN���Gsڻl�D_W'X؊���k�=y�]����<ú�۝Δʐ�ܶ�6����U �I9�3�#&n���pz����T�PH$�L^��IJq�Me�m7۳��6rHS������Ԧ6`���E�a}��X�cb�-��z�=��GA�����R�tw�w�pu*v�-$V�&!�<�\j���j�:֋hSwq��<��k=��$��y������髶��'�M-*�wS5%$����YMVYTG�\�n�^}���b�J�[*�e2�i�b��:��L"_��c1/-EuP��l%�6�jY$za�&�/��xB�OO����q���y���淾���Y�Y;�黬�8�;B��߼��u5���i
g(;E��&OM�}>�4D2bv�,&w�	��U�h��IM�h�����Hx���O�/�M��qז�^[�<�yKm�O��N����Sߞc�EE���5�q�w���ʖ��M��D�7�1ٙuƌ&�Da.�뮰���-J�11	Z�I�q��Z�Z��&��	Ly,�Y}��D�����m�t��xO\�nxBG�������?M{����V�1H�R��A�|{��KEDS�x���}�����٩%1r��)ȉa&N��i��9L���FBa���.�$\y�\�e0�z���S��{��H���s?m�i'�EC���Ɗ�!�}���1���ƚq�Yi���[�|��yk[���<�������TC�:S�C�|	&A�kǒ}o�)��%�k��q�U5�;IB�ÌT�W�Ua(�cqqۢ�&cͪ#�t���OS5)�s����(P>������jTǲ�1��1g����ی����~�Ȥ��*D�Ek�����x�C��L�����a8�o&o��G����MJ�-��rUV'>a�ũ�#�<�1UX��e�N��߮iSQOi��zq3oGq�/0��e�L�1�zQ�~�ݙ�3�b$�?f{�]K��LFR�>mn8���V�ǞZ�J�[N��)���Mp�\���>
(��O~񜗞�G�>��\I(�+oi8z6���M�+ͰPNxN��_��hK6(�����6d��|���L��HˎUM�x�n��~fJ �O��tH>b�XK��J5TK�E4��I(�Qwr������d�wIl0@#���>7�����z��GA	D�'fg��>_S��l�T0�,;1�UNeU��Mb��Q(�9��ۉ�񄺝���?;���T㯛u�|����8��[�[ki��:C:�ƶ]i�$VR֕j|t��N���@�E�[<P��|�c����ܽ)M����͟/[�$'jyx�Ĉ�4]x]���=��vz����WVL�i�)�(m�25�R/z	�@#��.�R��nlAT+��2v����ϔ8x �Q]�OUm����1'�1м�Lk�x�qB-)�=�e��Z��t<�C���R	�����qno�8�e���O4�w�;����[�̴����v8�D�g�j�aM)1�c��q�9�Q�D�%IK�g��b�f㋩���S�b����B=ܚLWy�w�����#��xQy��G��eUX���G\K)%��)ޡ��Q�'�'��zz �����q����5�G5ظl��]�f�ni'N��ӱ+>�g35Y�Ѧ&4�0J9�!=�[�1k�Lӓ=��FYy�|�θ��Z�um���Ÿ��a*QӤ:t�|7���"��QA�/���ݝ4�D�sg�3)�q1�Vs	$@4t0��i?�΄����2�4����LWiD�R�+i�ډE�V��m��M�s���SLaU3��FqD�<�m�c�"�y�'?����'���ܹ�f��U���K5�L_��v�h];��/x�Y��4��unfp9�5٩��dc�k���&Q�@#���;����3���י%�����U5Z��gpϦ'zf�S�y�u��V����x��l%Ji�4�IuͪgzL�I%�g,2�m.*�z��Գ���%��r�H��'��ƣr�
%���L�!�S����	Gѩ}�����cJe��J;\�0��1��FMSV&�F��U�j�X<_ε.>wI��IG`.5��̘i�JN=�G����/���O��s1�im�Xq$����a�&�o0S&Nc��d��Oy�r�kOvz�RH��v�L����fbe2F%��i�y�qžZ�um�o-�qm6��SM:{_ן��B�EJ'W���E&I%��f�S����UJ⫟;�@N{�D>L^"	�y��,��5�CB��Zع����z���il�M;VOK�|�x�!���T|ʒ�Q�B�Lb#�Q�UJ��3�y�w�2_����!
Jt�7�`�^���ev�O��� s��D�T_�L�8�Zӌ1���V*���;i)%�L ʞ�ң��P�Q�&~n[�L��UǼ��1�$�z�a�}�Rr�m�<��y���[�u�-���
R�iM4ο?�M.Ո�omt��:v�M���򐅅�"�j�$4,����9�I�٫�gs
.�;gc�:�UE�k��݃xK��J�ƷX�e��֭�cG[7{k�R�PA9�Q�blAϋr����a�A�>��p���A�MZ(dn�]}G &T�Z^�-����u.�޼�.㸞(N��UP6ÈA -2`z>\r+�5��D޳U\2J>�ⳏi�&]�ե;��=_f���v;��e�j�f!�#����k)�q	p�Y�W�$�1��qzB���Q�A�����V�諹�*5�&��SSU�yd�yޭq��%�2z���ӈz'�BԼ�)�a�ǳi�'E&L��p�?����8r�����r��ktud$q\��G�Xk;�c1):���Q*�y���N|�Ug9��&�UX�a|�F�g�|��ۋuż������[���i�(�!E�֒�F4��A#�����W�De�q�V]f�������LMb|�v�b��d�_;�3�u��ʪUL7�R�}3��*S^�E��^1�K�[�'>%�t@�3�`��',Ɵ;�n*�R��&	e�6W��[m��K���o�H�ER�A4�g�/��7�D �+^=,Ļ.}=��V1��e��%,��y�����@O�:?~�w�����ل���/1mG
��]u�-j�դ���:�ϕ���p��>V_+�<Ǔ��>y\elyJ���c�<ǞU�]K�+��ż�4���<�<�8�'��|y^m�<�Ҽ�'������O<�S�S����|�ft�����Zy�qKv�J�ʧ�c�4�<�<�6�W�伜��������u6�&)>O\S��i>L�ɔ����)^O����1>W�����>f�����ʧ��c�S�+�VYVS��c�+�+�+��|�<�0�y[mZi^mT�'	�O*S���yJ�|�ZeY|������ZII���*R��y:O��*:O��+�V^Wft�'�T�N2�O�o9��y>R�¼�,y>O�q�'Ϋ��[��o���X���<�4�y^[�q�y>O�e�%���y=y�:�����������]f���t�0�K���y�y8yOL��<�.�*��cɦo7��<�Kμǖ�y^y^O�q�&^W��|��l�и���ם�hŬBqJ����u��kE.{�=���0ks�cPk} ��v�:���z�w�!>DVU�ZsW)�T1��v}��烥~N
��<�Y�7R	���B/���H9��{]��[cb|C�4=�o_�)�����45}���A�d4����}4��+E-YC�E9ѻ` �J�ry�ˉV�e7~O5�^�u皗��{C<���wԒjI<���$���$���.���^m�u�\y��V���x���L)Ji�4өJ�8�e2�%��0���s�D��Xd�]������ӛZV��
%��Ɨ���Lg0��F�>���A4��;�	�ѡA/������Z�kda�H�6�l������F�㧣����J��7t���0tgA�(8�	�?�7��%���>`�DD����Y����V�XW��4����/��< S������?h��$��G>���u)JYb"z����F�r�d����2�!����{� A�h��>JO>qן:�κ��Z�Z�[�y��[m0�)���N������"jש0iޞ�(""y�r��ޱ�bk���ދj&8��m)K�p��?�<(��'�{fܒq�[f��k��sqc[<��̾q�+��-E�s2�v7��)z^R���}���cq陊JR�#9[LKy��q)JR��7���Z��#/�JR�-s)�a��v���MM��Ķ���Q�<ⱨ��c�3�hDO�N��=�'2�S�ц%._�`�Υ�y�M�u��:��-kuk[��o%m-��R��JQGx��>�U,���X("��k$���NAS	5`bYAP���ZC&R�X�Y�{tْ��u�wH�B"�8^
2#�y�ԃ�i�N��s�g]��s��:��Ĵ�mWFLm�4��%��k,��PDD����~I���Ƿ���5�'�؜Ӓ�z#q@޳����|�$CG)t����o�N`ۓh�"�C
�LŖ�o��\E _Rq��'͔��a?����9竊xzxr���\%=1uM�ϸ�R�`��K�m���,r���DNw�[)>ac|���)H�DO�����'�^��y����W�������Oy����w�落���""�z���G&+4���L\Tv:��j1E:�r�����O��i�撮P�u�냯m��������'x������cy�qEbV\S��m��u�_:��<��Z��[�[Km��4Қi�T�uSv��f뿕(����=��W��&�f8�z`��2A.��j���cgHuR��7����������>��5��8��I<>}�Zfrʚ��$�f|����'�5i��*)6��S�3�n+-y�	>��^>��ִ�d���F�74�jVk9�mn��4�L�䩵4Iإ6�517�m���JRI1mq;������┒I�{Q���i��iN<۩M��V�:��V�<��uk[��o%m-��R��Ji�V���&jV��(���ϝ�)�����=�}������| ������t�����~�|�@A����	���U�I~O<_Bs� ��=����zB����T�;ss�lٓk!5���$�|���0h�F������O}����=�O�	�xc�=1���8��
z&;ƔB3È��Ų�tB����H!�f����툧��}�Ԫ8�im&��ڈ0e^N�e����u��<���-խn�ky+im4C�Ht��������EB"P ���A�糨�:( tQ�|+)�D{�9r3�ǙST����Z�b��>�k�v"�9"��I��W-�xTk5��v���:�|�i&>QO��<��$�ȵ�_���_�,>y�J�2���)8 w��~��?�X�C�(��Ǉ���(" ��1�8����}�#)��T��N���c�R��،*/1y�ZRRf���|���S�3�ѕ8��Sډ�5n;3���N>m��>u��<��Z��ֳ�im2��SM:�����Z�lm��^�׶:&�_;����i���U����^u�Eच�x���m�u�����^8a���J[K���˱ӱ*��fN3%��XK/�EA�~�����'��L�U�
�/p�i�t��_[�jͫ�\խ�bYyy�.w������1�,$�2A�Vr�u����)��ɘ����4�em3�V�靸���2��+SG���s����?�p���ߤ��B���rkQm0��n�*�:���q$��<ʡ�x��u3�܍6ҢR��u1�}E�<)M�"��0r��ʩ%i7�sZUT�<QQAW�����D/7���Q4#f��L;JU3"�ٟ��ӑ�����=��������`C���	m��s3�L���v���u��Z�:��<�έkukY崶�aJP��(�����!��Mu)���&%�Ze2JN�P��Q�����8�T�Ye��9ʝ))I�u�����Ϗ؅"5'/�jD4 @�J0��rfff�e�	9���6��^*������ڙ��E���)%,�%��(:���ڣ�@,@�He�)D�Y���ԗ�G������:ʒm1�ѓ߽T�V1�'q�>R��<��m���==j7u�$���8���{3��o4ӎ�[���-張�����-�XR��Ji�P��Z	|PD)�
B�ߍç��t�"�<#��s8@G�9�O�H�yGY3��у�@@<���$��4�ⶦ�I��>�Xm-51K�":�})kqL�Z�V��#M$ۖ�M��-f�����G��0�̰��vf��sK�\�=ǦX�a��jl�St�sSIe*JM�~����x~�pQ���Y��rbr�L�ߓ3�jڍ��׽3,�0�$��<u�ӭK���ͼ��[����Z�y���-n�k<�Ki�B:C�O�����HəS'U
'^{�QAy~��'�O�����.����9RL)��+�\a�2��nQ��1�!%�[G�I[6��d?2|Fy��V�:��𧧓|+f<ѶY����Q���J~j+V�Ŕy������!�D�����>E�"������=1�������>�
��R���&:�h�I���ϟU��ODD2{W�Hby���7
����Φ�����Q����%�I2��w:[�.2����o>im��^mkZ�J�J���<��<��6��%kZ�ۋ[��뭶ۋ[ekZ��ֵ�+[kZ�Z�Zֵ������ֵ���u����Zֶ�����������������J�J�-����m���ն���kZִ�k[	a�-n-jZֵ�kRֶ�e�VZ֥(��ZV���jZ�Im�o<�K4���<�,�kml�n��֗����kqn<뮺ˮ-מa��)孅�n��-kSZ�[�uź�ZqKS��Z���Z������T��ZT�+,���YakZ��KZԶV����x=5�S�j J/�\Y�� �Q�e=մdO���~����f�Ɍ&�f[޵'vZCjfSR|�7�=�f���mO�I�Yo)����S�	F�d�!�9G��;i��i�cf��Ֆ�M��T�<��1�%���.:KH��e�L�e,<ƺS��6������=.$\��I�3t5t���I4Ң5F �&���3i')wM@�w+qR;Wd9��J$d����Wڎ�D�Bё��i�ʩG�(T-�S�HA`N쓑$�oj�D�#�C�[�aB����#, �4�۽iߖfI�Y�����8��5��=���6�����n�+�Ƹԥ�h|�z�J�Eq��r�	�L��>B�L�-�0�}sF*�h�]��ڇ\LDT�8�z5
����ТH �(�Q76�nQ��2+]43Ǚe��9{��t�������p4�b4��Û������~�X����s���u��
���{w��@�̘pW�!�ϗE��5�nh*�ۭ���0�,�؜�8fr�M�4)*�$�n�݋;6����	G�gv�⤝��u���{S�.���nm�R��2��uz�V=ڲ��Xgg���\���H��:�]�m�A���.���<�2�wwu9$�I#c2���ԫ�\�YYR�����-�Z�Z�y��,(�:t�N����e$t��\�iK̾�/mW��ŊS�����^�Z�����.�-�>�������b���G6Vi	w%k{[n�ր���[�i:��3��֞l�<
�P��[-�1����+�:�7G��Ռ�D+�2m��g���Ɯ�S��}��JnܭZ�۳�:���6W"�)vm�
{-t�n��b�r$�0�2����n(�@�OX�t�g�IB�;w�L�<�w>+u�d��V�#���M�h;s�����nWG���4]I��R�2[K|	�A�n{{f�Ep��ޖ�6��bjNXWRT"�X��oV"�Q���k5����a��f�xP鏂��p#�JA��2 �<�	q��Ǯgq��\JRv#Lr�m�#�9x�J��S?R�V��5,$�Q�'~y�鎓�!�M��o�aI\��5�g��	���S/\Μ\K\Me4�a�q�}Ti�^m3�L�߾��9J_h����(�bu�bKl��Rc|�	�q����x��2w�t��;�V͌�f�V�Ĵ�Ҟ��s�;8Q�L�"fc���p�,��R�|�1��g�c�eQ�%��m�o-ż�^y���[�Z�y���
R�i�>?}�����:9����Ƚƚ��U\x��^��kfRNә֦��1u��ϓ�Ғ|���0ƍ0�os�Ҧ��.G�n���a�2�RK���ҙe3:[/F��0����z2��F�Z�_C�i&��f'�a�nj�.�H���?�z[|;�-Dʓ.A��A�O�����>RN��Y�~�U{)�ft⸝�ʒKԨ|�јe&b�����b��˫Lqh�c��|ۋyku疷�y庵��[L��)���N�i̮\�:�L���D�M0�,�l;�oK��?� ���|��J�����}Y'?s��|��+���s��""!��ܥ?�~s=$�kl�Ab#���*�8���yZa&��I���'�\[���JM������m�T^���L!�	��o�~��y���|��F�T���|��ߓo|0'�'*L}�s����O�<�=���\��K%�V�c��'�g*�֔�䙏�&ٍ�/�r��O<ێ:��y��yn�ky��,)Ji�4ӯyt�Ó*��[g.�-X�9��I��98t�C�-��	"�����\J\f�b2��EG�T%��F!�#�>���]���8���+�u�3��vjw��%=!y�C����zn�}��јg��/&3S����$�¡�e7/����t޽u�����aj�̴�Q�k��]�<�&;�S��� ��~Bz�:`���a���>���=멪mw����.4�έn�����<�V���Ki��4ҚQѽ�~Ť�p����q�T�м��h�!��2cQ;[����_����ssT�dn^sE^g�9�/p�!ey����g;�WX��3��|� �ɥ��!Xq���c�y�0����iT�������|��i�ʺ��^Y�3��jLKI^[��Q�b�b�C7oA�J���l'f�]Y�����C8B��S��v>A�t<��Jp���r�b��ᜣ��~�'������lC>���m�e'Ȓj'S*e�ӟSN�&���^���a8�4nXJ��Nƣ�/�d�y�ԧ���##E��<O��;�x4�AO>����[�?'������ȍ$Μy�io	I?�}>fRi-�p�m.����&��OJB|Q
�C����H��US]��Vձ!�=�T$�H{������)Sm�ۯ-�V��-o<��:���[L��)���N�]T���k�e2JJKa�#�aI�q����!�#v�o�1,=�i&�&g��1�^�;ݹ31X��UZ8�]���x�Sq�n���)I��0�:L�9o�A9�OL~)����n"!N�BNN}�A���cdX�4�"���u�K,v�р���x.��PC!r�>���_Ƚ)���� ��/yғ���ϧ�RJBp����T>���y�]uן:�^yky�yխo<��e�)M4��uSӳ�hfH��2�%&#܌<�|��\m��U�4i1M�ٟFMĥ'Lz3R˭�����ۑ*�RR|Hz<!�=�A���h��l�b�4 ��sm����>����tM�R��X@�V::>�=�>��T��^j4��S{�i��URod���"�'�}_�=�C�D<?�	?�r}�6�T��0�C����χ�<>�1�>�oq��/t�2wp�wn���|r��'r�t�|6��>yխ疷�y�Z���-�XR��Ji�ZC2gS��T�(��<O}ό#,�~'|
C��b��SzS������o�u
J�Qn��p4��)��'���euam����'�H�1��q�6=_W��V_�<>G>��|�'2��3�0H���)%�<Ѣ�����q�+,��kS8�g�O<�:��tǟ����ΞrB�%:�������$����D��V��>u�yky��ֵ��Ki��4t�N�9�a���MF�&��N�Nd�X�qB������NȲFH�Q��D��:��3�y2F�`��Wv����/e��jE9R'�B�׳td�Ӛ�}�s룅��μ�/�6p��p�$Me�"f�4v$n]ESC9]>~PD6ܝ���'Y���Ա�nf�cc�ᵉ���(�`�t�����r�� mE��T@�܅�z��#� ��t�i&���i������#߈��eL�a���j1W�Y;���M\�S8�>TS�:m�bz�coLm���!1�Q=��}��%��a�\���\|��w����q���j0x�i�!l������!���}:N}�:i*I+S���b��c�)l��ˬ>`�!����ᡂ|��<Aڤ�R�W6�����s�ܯ{�ś�q�=�h~���;H ��C�LQ羼��V�4o??���"p^��"e5S0L���3�_>i�ϝuo�yky��ֵ��Ki��4��>=xg��E"Nr<�x+�t�$��<B�g;j�gneZ�Μ����!J�\��[Vݭ�u�e�Ǖ(�=�ޫ�xt��!�I���+���Ie�ĥ'*<ì�agpþ��my���" ���1~(�x=�, ���>r��?����t����j�4�ke��$���f��S1�)"�qW���/4ũ���Ǉ{q�a�%��3�4��='�|9iie�$Ï��u�vj���������ʽ�I}Xss�ӽ��6�'��1X�L���{�Yc�N�&����>Z_-��ke+[�Z�����ն��y/)�y��q�q�S�Z�������kZԶֵ�����kZ�Z��V�ַۮ�պ�-kZ�[jJ�Z�Yk[�-m-n8��Ɩ�VYe�+mk[l�k[E�+Zֵ�n���Ka�-kZ�mk[Z����M2��ZԥYkJ���K[)-��o<��:y��̶�Z��+[����JֶV��Ŷ��.���yOy岵�k[-kSZ�Z�un��ZmKSf�Z���Z����[�[�[����Z��V�V������l���c��N|ǡ���������Gg�WJ17Qy�e���K���^:��I�$���k�����D4�ǈ*G|��O(��_k�uLV��9p�+	�XCo��w�c�������p��G�>"����	9�E�E�E �Y��Az��|z��W��^u�s;׶��\̙Y�o�ɒ63!�]���;c3#�����$�I#c3"}{����q�]uם[�<����ykZ�y���
R�iM4��s��d�o�W��z��{����%\i1)IԪ�Ty����h�*R�I�L���v���Q��9K*I�	���!��9����|x�^�ӢA�x��xea8����*A,;h����V�0�4>o?^i$^=c� ��1���:���ޟlws�[�R�s��Q�N2���K�L��,&.2Ҝˎŝ���L�8���M;2�N�R�3���fZ����I�)1��{�B��N��K|��Ϟyky��ֵ��Ki��4Қi�A����ELC3��x��o\��xw�ۇ9��r~5�AXxN�ޯO��y}?��S����Ԍ��Q%�	�D��D�"��'9��'�TGX{D��t�*Iםe����L�U5Q�Kk�3�R�zJ}l���Lf>��1�b��y��$�BT�{鮥ښL2��<=��$ ��~ ��ҘJ���*���\G#�2k��zSZPCޟ���I)�μ��˭�w���ƛ�u�qo=���<���<��o<��@�!EQGC���\I<	4���|���U���o�����,���W�k1ozo�xܖ3��.�\���m��+V��V�dq��A�4�Mû��{?v+"���H'&��ݣ�_�L6t�&o�ǛlJ��/���{�TA���e��H�^�(�L��+�c�|o�Ƈf�.�%�%�..�����UX�w�+ty�]a��JaJJ%�n�55�ˉa�0�*�am�ۘ����W�e5��m�K�ƌ$��%?qaӧ)9	�:�SB��=��-��e��1�jg��)(�"X<���:w�4y�A�s�9I>,�����}����RLfg4Ҙd�O����R�6�v�-��fm!Nu�XdU"���\C���̒�<�Q��I1ֺ��I�g��V0�ݸ��u�V���y疷�u�Z���-�XR��Ji�b+�4����5��d���j0���#Z���C���,�M���"�j��x�|J�QB�O�|��yU!9JO|Ֆ���|��R�WS=y�6�{�V1��	$�|��O�>��V���|���ڒ��c9�F\�13���a��Q'Y'R6�ˮ�CV�)5-�ݲݝ�<��a��R)�S�yL"	�H!��zxnt�??�ef'��%'[L�e����L��D�am0�R��L�-��G�4ꢢ�i��y�y疷�u�Z���x`�A
(��:#|�H4[o��?�)��
%�Ĭr�&����%���)o4�)�-�)$@A �����˨��a��	����2����D��O*�������e�'��-IK�,3"�$$q1O`�0��`Qr�dL�x�|ַ3jy�Jg���cq�bX�*4�c�&��C1�^4�|��H��)+_DϚiQv���m������[�ƚ%�y��ba>�i,�'"
)��8a�S8�_F���N6�לq��[�Z�yמy���L�JSM4�N#�uSSFfey�/�E�I��
&˒zN=��#��gW�s��ճ*"1IR����J�i�K,�ˌ�}����O���Q�ra!.5Ks6l��2�"������t����"Qy�L����<:$4W3-��ÉRQ�i1���O0�%��>H�	�&k�N�0��&��%&W<-�Ue�����[-%O_�kg:���x �u䉇��D��&)�����m��R��D0�S7�榧DǟFa�ϝqn8��u��y�yo<��eJR�P����DDi�rCL��2��\O�����Sk<�+��O����%���[!+g��B���~����z|�6-kGn�_&u�X�h�U:8S�c�Oh&�&	6�5�{�袂!�zx�����Sr}��owQ�]dZ����)��=�����d��%Ώ%��y��2��ut�\���H�k��0�;�^�i��UiJ�RR�!LS�N�{,����"!�>byUYT}r�>m�JIJ����q��赭�i�R�1F�s�_��R����WdL}y'��A���%��mGm��e��R�#��i�&��6��gx���)��i�0R	������V�I2\bQl.xH�h�X �������`�	}�0�x<�����=?��?.��9��u��8����[�:��<��ym�ʔ�4�L4��I��_ޑ0
�;>�("���[`�L71��L��;����i�]�a�b�L���k�4�$�κ����8�b��c�s�=���e�6�<#Id�L}[MF��ک�L�̰��q��"�I�*���L��� oߪhM��TB`p$�Eċib\9�iyd��<=9ӻq�!�*4��F"c���k�)�<�[�e������@��P�;N��4�����53��2�F�g�N����[4��u��yky�^y�[�-��!C�N��>�;-<PD?��􌺝?�x��?�=>FG��8Q4�u�'M�ԩ,%*������8�N%6��W�����i�u3��ḘI�Ӳ6sh�M$�[���8x���r1��ۥ-������Z�x���!� )�IO�����j�8攥G��	LD5(��kL{��1��)�%��R��>��iI,G��uX�'��B��[��̸�lC=N���.���8����[�:��<��ym�ʔ�4�L5T�&;U9���3Ng�o�EN@�����Y���_V{û��Q��O����wIכ3չoy�rV�՞��\�"%�#�G u
~<���x�qH�^-��*�Ma�xE���5�/�)a�G��zsڟϐ�19ӧ���%Ľ�+�U5����L\i|��$��Ǆ�<H��8?x܌�u�a.;a�
bYKIr)����}zz<L�+p��~�Eo�K��ȉ�ej��[[�S����-n-ka+Z�ak[kZ�[IZ֥�kmiq��y�]a��<�V�ֵ�����l-n�+[kZֵ�n-jek[�um�juku���k[kZ�-iZ�[J[K[�-+[�-����ZԵ�fֵ��ҵ���kZ�YkZ����kZ��ֵ�l6��m��YkuJR�-iZ�e�����Im�k[.p��S�0�e�yմ�Ye���kikZ�i�]u�ZuǞy/y疵���e�������]Z�[�6���l-IYkKK[+[+[�[�[����Z��V�V����������o��qQL�)��X�8o1&�Q�[K����NnD\yw���J���L�Y�
{u��l�nݻ՜�"�]����%{�N�T�;�hIc->v�3 �ۃ��N�m;5J]sE>9b�Y��sÅۅYY�,�m&�&�f�Yغ�L>�iI�nL`Aki�,CH�&'UP�0�Rā� ���d�$S�]&D��I
t�ws��;݂y[	��
xp��`xq�*r2��hN(O��b@�8Y�d5"�P���$p��iH��=�I6���6��p�)P��1Ό"*�œ5�\?[2��p\��y�����CFa��t�Wc�Q��?n��}����}�֝��v�u�̚����
�ێ��P�Q�x���x�/�R۝c]F���[h��c� #�2=��Z�8��'`�A�>����
68�V��Q�XG32�K.0�a�e{֞�y.x���82�B�,�*��"K61��U,���ɮ��Ws(�LJ�qen�e�.z^/�mz�R���ؐ�ȃ���W�u�,�f!:�j���_�`ߍh�l����d<]����[�9+���l�$�Y�FOU�X�߫�3��猦�t�m�Uo.�<���N�BVskO9ߎ�`�3=�s{ܒd���*s{ܒd���*s{ܾ�T�\����Wyn<���<��-��L�HC�N���O�!÷k#�ś���@\����qdۜ�p��T(�o%r�i��(�.�s��� �ݳ�eu�Q�t��m���7�;�]��t͠�l�:���܁��8�.H����i�r���u�g�sj;rkp�n�'_|c��)�Fg\�B%!mKH�5k/+��3���F��ԅ�'��n� �8{\=�Ή"� �K�7V\��,�!׌ɡYIW`�FTJ��b&U�mR�q6�8��f�E���V�H�cY�QAu�{v�N�v�;�|�$��ϺM��w�6<ѓ�!3���u/Y��CRIt��ąO��4�{=Uɝ��֒�Q�!�ct�)��~\|�[�E�э��L��>R�£	|��3�����a%))v_9C��rU���7SXv=�&���YJz�I�)~�ӌc�o=o3]e��򛌲��LҒ���X�R���`� ���0�����_�KΛ��%��?��J]�����S���zKg5sf�:N����MRR��-{��&��ʥR�r�n�뭺��8����[�:��<��ym�ʔ�4�L4�zQ陉�;rn�s�n+gu�n�k�J$�'����Ďd�xa����ؒ�fOݨ캔�DRꚗ��'u4�MJEǘ\m�T�R�R��,�2�R��D���??��d��F}���|>p�O����S��a��r���Ky/��X"�Z����^�j��0�t۱��/�p��,q�X��j:fJ\��Y����'n���>uih�b!Mjg:�jSI�:�q���9u��|�8�����μ��<��(�B�(b�����d���$L����uȿ�S\���Z}�L2��G�3��iu3�ZqEDƒ�����8��G�Gϙ��!
����K��L凚z2����]n��e��I{&�k�w��Btݿ��Ǟ1r�S.��_R���3���Z�%�2�RZSo�3�M�v���S����U������' �~<	����%����o���b�0'%�<��8����[�:��<��ym�ʔ�4�L4��7��T�fd�X�v�������)�8Z�Sh�XqQ,F=u���b�5���	��v�$�	������kl�O�yI����uo�s�_s;E-R�L��6m��z>�Ͻ37�6����4�N=����u-�mٙ�UO/i�0���~[�o��z�l.;����&Y�bf��K���ی�N%��S�5S5�&�8�U�c)�JX�1�Rf�U1��|�ǟ:�\qo�㯖�μ��<��-��R���i�����gs9�s�1��e��;��]_!#m��۶�R����چ������#�?��|��2aŕR�bZ�m���szv>�#�xw��#�J����)�g6Z��ד��==?�������y��u�=%.��H@�<�����Ѣշ�Ȝ.�4�B������ܨ�[��x�o��>��A-aX����1�e6�[lu�0�)-�E�R�A���	&OãF(�y���#n�y��4�G�ۙb��f:�Wi�v�Yww��O#�a�7�Ϳ�iu1�_F��v��a8jY}ĥ/�{���'ΙK֙eۏ|�rJ�|��Ry��54�]k�4h�*Wr������ٯf77i����S��>nf܎�y-0��-��bݔ�תf�Zv(����8��mn���u�[�:��i�)Ji��;� 5����	�PD���7���+z�Җ�\�U9ɪɸzS&�q���iMRۍ�±3L�)�fv�ZAlşLFa�����ǞkS:B1D�t�������ޝ>���vG������LĦ[J�%mJS���ck8��+�K���;igg[�a�R�>(�#��%�����<�w�m��%��UD���\v.㌔��}��bp˿L�]��zS��Kl�3(f4y�->yn8��[��o:��-�ym�ʔ�4�L4��v��f`S�����Շ��a��ߏ�=���T�F&~YK�
�|����Lp�DW*�gd�USZ���i>���E�}��Qs��	�N�A�	ie3�q8�1֧���6�ѷ6�I,����ә��j8�NG��(�)�[��`o<��)0�����>���Y<$��^4�iji��e��&���,^L�a����Mff<m�ӎ���in�����<��q��*R�a��t�;�Ouk'#SkHsNJ%���<>g>Q�?n�Kk��ܿ>]�J1+�[�7IOw�Uq��������`�_|-���k�<b���ɚ|��]f>���G�|�4�e���S�)e)�&fv��6ն�r�0bƦ��n<�ye;�zO�	�U虎K1jvu�g���J��}����N'8�L��^S$��d�=�nj���y�ͺ�-�����<��yǖ�L�Ji����=�����j(�0��A廸^�:�&�X�Mde���Lm��DT�+ �	 ����	is%�K[*2�A֊=c��r����[����;�~��1�4�oIo��{����sS£)/��@�tG>��{�msD�Q�)9�4&�k�˙���&�^��e"�Fwb�a�K�4Y��5��a�����!������8T�O�n�N�ë��S��Lb�H��	� ���ߚh �1��n��Ow�����q�{�J̦��g1��<�2�]�j-��?=2���7�';|Um���$�}�1�����D�!��Z�)�k�X�MFU��U�vi�s�B�?.���&�<���WyQ�0ө���wS$�,�M���q��4�]Z�:��-�u��Ҕ�:S�t�}F����/�I<|3��80!���M�� ��G�\q8�6�N�U�L�O�f>Ls���U��)&ڗ�S0�G]{���L�}K4ޑ��TL��ng��T��$�'[���=XVIƚM�C, ڒG7�nq��b�{�,�j�'�n������}}=)���y����5����|������9eS�*73����q�'m�\��Lb��L���a�s��ʖ��Xx���֥����ֵֶ�����KZַ6�kq�-o<��<Ç�y���ֵ�����m-kZֵ�եkmkukZַT��Jֵ�������l0����ŭ��-Ɲe+,�֕�k[k[[KZ�[.-k[��iZ�R�Jֵ�kZֵ�kem4�L��YZ�R�YkqKa�-kY����Z��\4�kJ��ͼi�yo4󌬳K-kZ�Z�ï:뮺Ӯ���<��ykZ�ZVZֶZ�[�����i�-M�ajJ�ZZZ�Z�Z�J�Z�a��Z���[kZ�Z�ZԵ��VX��MgW5��Y���]��h�Tb�Ca@u<�dqm�J�x�Q2��EWR�"�(
o�\�1d���*�N!A�p� Ws}����a���$�G��!���}ȼ�V�h��@Z������lo��,���L)T�	6���1��i��?�7u!��}�K��u]�5:a32T���rD�I!ffJ���$�@fd�{���U*T�W++�8��-�V�y���8��aHC�:'N�y�PK�/����Bǘ�Q����ct�Kf1L5�u����I����� ��L����e�c�Lqǌ����V9b���;z����K�ov�����GT?�6Y\|F�O�x���8��/���Qə�Kv�����|�_;��q�9-��k9j7�TKp�q�����ᨧS˭nʰ>}>u}4�gQ�<����8��[��n<��-�q���
SL4��Og�3�p,��H��xr�|UA)�xn�<���vftڢ10擑��b�i��]���?9(����B^���k,�m�̓iϧB�����ΐɊ[����멚�΢��a����)�B)�MD*`���^��c9�t��gN����y����/o�w����0�ı�q����G�/�L+�Ua��z�ʦm�E,�����z*f6��|���[�<�Kuխ��<��y�[L0�4�Ii���Mc
a�1~�����[aeu�>vS6��}��}=.r8���ۑߵ|}�_w���m���<c|y��ݻr�ۗIZ ���B�"+!7ߊ�%��|�G�@��?�������m��{C�t��:ף�&�3:QZ�S@�\M�(��{2�҄`ٜ`���SX��gh��a�� ?���k���=M;$TÊe�7�¥2yn4�kyn��ËiD�"�r�[+���{<��>��1�]y��U�$�J~�%�D��$�1��nx���v�����%��b8�.��j%�c��]J]�{y����OgYUK,89�Q�n�aA{����Ɔ���-"�LUהPF?w7�%߹��'"S�G�0���{��KK�nF��m�����ukq�yo<�-�R�a��ӱ�k�T/��2T�C<�*̄�睊+uz&X�������]6�m��wزڒrZ�=/:$�҄:}�D�E��A�R?�K��?��}A���F�+S��eķ�L�bgL&=<")�-�g�t���(��p9���@��G�W�	��m8`��ͣn��76���In�����ƴ7H�N^@�ҡ�y����=y9��$���|'���c��&(ߣ,��)KDd�_�{�h�-�Ϟ|㏖��ukq�yo<�ӧӥ)t�D��QWN�U��#/�)�KM�e���;�Wʊ�G�Bz��w1��y����?�������A?tN_@c��'�"Dy�k�;M--�f�O�>w)5-�`�Q����XK�I�D�\��:y���]sH�)�w���x
���,K$��c���Ӌ�i��%��\Z��J]��z��;�u?T�O
ed��,&>�L�ͩm�kuלq�[��n<��-�q���HC�:'N�����ϙU�m0�b*'ѳF�aKj0�����>�H��ż.l-���1OOf���)��|�&7��Ox��6�)�&ff��)1+�ӈTDF;n�[�f�M��W&��~ôe�KeQ�[2���ǳ���#ܙw�<�/8��X��<饺a���0e�%��m��8n9��R;ډbT£��y��e�Z�qż��ukqo<��y��[L0�4�Ii�^�����5ed���;x�&I�&�$�+D�lX��&�B�'a�k�ӧzJ%��n�g!�ZK{u��A�˘Gey�n,D����*��$����3�^�E�m��Q�O=|�uEV��YڨcV���(�vL!��9��b������o�N(�Q�;υ�� '��S�^�I�p����?�8�i��b��4�ܙ��/���s�#D��'����Z� �8�u�f.4f5M;����)㭔����O��>r�c�#�ϐ#�1����Xq>+鹏���RZ�'J]1p�hF&b�l�w��gU2�z���kLt�sm�nF~�6ۗ�]b��iky�|��[�8㎭�����ַ���2��a�)ҝ�y�Y�~�)�*��O=_���Ź]�bb;������b���F�yk���a�U-��F���R�MS)iN:�F\�ɦ��bt�V!�\J�8�U}�iS�V�Z�����ɔ����	!#8�/��'�E�5��'�,�T�A*<vJ��Q	SYut�Y-e_�R���lg�>��?2��r����>�N�c�	;^SZ2�._':��s�[}Q���2���8��[��n-kyo<�--�R�a���h��`�};�f�33$��i[n%�T�#-F15)�p�^&wd�e>Sʌ���<��8��%����_���'��?s�9��!��ο�]�$�I#���!��Y��ͻ3��'�����fz�
n�n;l��ϜKe2���Z�汚iP�)�1q���>n���2�,C{�3S���=2a��R�B���1�KƿJ�	�������̺��b��yǞqǖ��ukqk[�y���a�)�KGM� ��)�yPL�{>������i�]0��1�۞��Î���*��:	!F���K[k.��a ��/c4(��������\ZYK�>���̦��V1e�T���3--����8�)ؗ���5:�.��U�0���̠`�DE��}ˤ� ��d�!�� QB��!�"�RU���Yo�p�Q��"0e��|�c��������Ѓ/o6��]qK|��ŭK-n���kmk[�i.�jZֵ�q��mn%kZֵ����Ǟm��y��kZV�ֵ�n�kZ֥��]Z�Z�����m�kqkRֵ-�������-n��JJ�,��kZ��ֵ���l-m�k[-�ku�akZ��ֵ���k[,���akJ��T��[�J��
Zֶ�[k[e��J֕��K2��o<��:�ǌ�y�m�ka�뮺뎼��<�y�kp�ֵ�����[�ZV�ZqKS��Z��֖��V�V��Z���VZ���[kZ�Z��ҵ����w�2�T�-���ɦ�W���x�έ��7����G��u�2���;mfM�n�z��q�3;o:�y����If���<̮9+j�&��/��1�bRj�9��Fk�m�H�)�g|��`]�o;�gJ�.[�ٱ��FTA��i*�8F�E���G�(��X%����*�d�i���x���g7a;:�<��'���u�:J�j�>�F>*������!W�1CӬeҋ��As3/��1q$�Ӛ3'DF�0�$qAK=0�s�����/�iyǻ
��b�;�y!a�1@�_7������n^L��(�d����A*.U)s\7qG |�{\>�fV���-�D㑙�^����g΄��35Ң�0��,LB�U3�N�WK�9��CfTU{.�C0,�6�N7���yK��%��[UTBҵ�P'J�p��"�ٲ�aĝ�F��`� �E�b���
B��r���edc��M4��\���&[����U��ݤ�+,�T��Բl݇�x)�Ϯў{2PY��4Ս�ك�a�_�s�$�T+�mY���,�[ndk�����>�.;5�^�ASO7�������ء��m�,t<�[f�vu����8�6������7>�ͤl�v�y����\h�����ӵ��.n�۬�qY׶3{rtn�^��U��ā^���D��e'�v|3�}����{�}:��rI% q��u{��J �����zֽy��m�y��[�Z�[�<���)M0�Zi����R����X71��v��v�\�N&6��=�z�sº��'hk&k�(�\��A��j�c���*�����w^tJq���B�Z�r�W8k��Î�"��'8l�Cn�m�7;�6�C��َ�sv7;�yau��l���v�ZmÝ���v��m�5�5D��=)���땣y�8T�cm�--�㝪��.v7g�w�\q����p^=��YJ�=L��熎̖������2붷�g�[�v-�d3$�FX3M-��	᳡,�}ۤ�e�!��?V�N${�Q|Y������Te!V�Me�x�"�Z�n�e\���,�X-�n�&�X�i�V��<�$$<>�H�K�K��3��4RXJ�_7��i�H�R�wI�o��xkx�����"%u3��J\\\al�Q�'�¢�1R&j>_��*�6�Z�0�b�����o�Uc��)˝���}���|_G��y9�D:y�招�L������t��q�X��J8�P�C��S�֝=�Q����Y���'FS�L�ʧ��37�j�Ie���K�Z�mn<�uխŭn��C�ӥ)t�D�O��UNΫ�|�o:t����PMΑ�?�^��O��I�Mĝ���ͥ���ٵS�#S�>���Ê���節L*=v4۱Y�T���y�J_�ZX�� "	���g/
~�9�K�{�C�����t�8���5��U�]lH
qx�}���͙�>K���8����HʾNy�zS����,���!		N�Ü���}?
���=>��'���6�-�������[�Z�[�SIK*e�R���D\�հz�U��^z���x�G���n4��մi���ˎFi��\��'D��r��柯�$��&�<���G1K��b�Y7,���`��y)�s���X�;��c�{��B�(��jbT�6�&��	�k����OD���9���Q��c�����m�Σ�':u���iܭ��))%�����4�`m��UK�4a��_7�p����k-z��Ħ~uĒ�����7u��e�:��y�͸�an�����ռ��i)eL��V�9�&�4�<��犨!�O�����l����Ԅ!y�=���S�L�(��wi��]f�g�c{7"�t���j=[��5mݏ��۶�#j�Y��|��'Y��Wj^�1�'�����s��SX��̾a��z.���G\�aj`��ջ38�F����N����\S��rb#hFf�Ӑ�JFX����p�
(�m��F����ͻ��k��K�'-C�5l���mo6�<��ukqk[�y��Rʙa���^�fu�f�5"v.�w�q��~R���늮�u�i�mv<p<�Z�t60�K�l@F�h�������s��)�^�����d�۶�FY��q�_�|�[Ur�]W6�[�Q�c�UA��'V��IM�%�b̵��d��\�����-(����$��ǋ��E|����;��.�d�\6�G������&�N�XO�9�#k*�zp����>y�(��`�!�Т:Q)$(����-��>`����I��Y\e�vgm���/'4�H��Dy�R�%lCK��xT�ͦc���Zj�\RT�?s���x�ؾ�.��Ϋ�V4��U�����
��̝`geI��a�TG��L����.u1؄>���)9�C����ߴ��Fl�Ht�i��:�.���y�����ַV�~?艈b�O�D�zH�xyՙ�Q�L;*2��e��F����1E�!�xw�|4`ѿ��gʥR�kɚ�D�^�nYi�<��ѥRC�)��w��-���Yo�'��=棱�)*��gM0a{R�q]y�s�]�iI��~�s�ʸ�1��;��~[-*4��Y���'�R!�8t���g�w�}`�t�:��=s:4�n�uĶɖ<�Q�73T�1�3�ӕ3pˍ<�O8���yl-�V�ֵ���yM%,��0����F��Z�x�Ȭ���[X�)�������Uo[�;n��É녻��"RK�����L6���3�ęf0��.<����N4��!�����ϟك��m����w6���<6��e�����%`�>i�2�%o&|ÑJi��f�ى�Fׅ1�z^�m0�۩0�2���W��31R��p�S.$���aӍ:�h�i�c�]�Ⳇe��>p��7f/�>m�ה�|��q�^an��ֵ�ռ��i)eL��]:��ǜ���8r'��� �z��~��C�'F	��FI�� [�0�Xi��Q���٬%S8L�m�g]f�VR0XxO�}L����V����p�#+$�i�L�>����l�2�o���D��8�ft�,sqת}��9G�Kjq1q���Yi����!��3.�u%8�cJd��^Q��f���ӈ�1S��I�j<�kN�XT6�J�a�ZUEu=Nfq.M�o�q�m�yKuն��n��i�YR #�����<��+'+��A!f{n=����s�?e�����1�f6Eʑ�+T\#rjS�Ҳ�<U���)X�b�Q6��Uk<(m<����u���A^�$��_<�g��	|�)���Ս۪Z1�>�R����a���)zY]Xc+S:s�mZ�¸����m�X�u���o�㌵y��i3	0�)���F����I+�|����N�kN�2�j)��UzcM��!P���N�UMF*�&g�L�N%o�u5�Q�������1�c��>���ah��F�#/�I�lF�M�lӼ�ܑᗫ��`�k\�;W���]4I@�AP\b�7�(up!���]|�>�Mv1e�[ζۏ-Kuն��n��i�YS%0�>|N��UPO�D�>s�cq5_�y�O
_�5�'ݴ�σ�a�5�2KsO*3������6�K�>��S�L�m7$��Oe�0�jf�*�8�Q����1�׬�������8�y񊟡�I,�J��r$]V��]�^��*�������le��.$�X���\�Tu����y����	=�ל�'��ǝx(r{�Ng�Ĝ�$��x|�,0�7�����L�$�p��.t|<<=�ܣ������<in:��n-����ql-ke��n�����l�kqĸ�m�ĭn�kZ���Z�[�6��<��<�l�kZ�Zֵ�l-�]Z�Zֶ�uiZ��ַV�-kR�[K[�[�:���K%+,�֕�k[kZ��ֵ���n�--k[	a�-kZ�Zֵ���ke���L-iZ���RV��JYk[�2���Z�q�m+ZV�,�ֵ�o<물x��%疵�ե�u�]u�^u���2��Z��kJֶV��[�qkZ�i�Z�8�ԕ�ZV��Z�[k-k[�[IYk[KZV����kue���k���u�9<��y*p�8W���a��J�S��(��z��Wg^�*�E_!B}~*n�������_l�����=C���*g<F�t�t����}�8NsH��=�hw�4��|�S�'��ꏐ��S�Bk��YdvZ�)g����P����T�7���x��$�p�����ME#b�`�1U�3�nM�r�[��H�33$�{��J���o��rI%@��7����u*Tq�mǞR�um�k[�[�4�Lb��|=�U��N����yϼ�q2�檕�D�)�E1d�n0^w~����j����s���x'�)��4�����D����p��'P<��칚H���nU1Q��:�Z�:�-@�i����جb�a�uӏ��L�\�3d�:���g�0�fo��Yg�=s��(��֏1������~�WЇ=i�peɍ��-����n-j[����kZ���(��a�R�w>���̪��w0{�Z���xxsӼ��{�����c�K�rC$P�1���;A��o�����?gmc��@4o4���â�'�)h�m��䲺ܪjZ�i5�b^�:re�Sq}0�&P�4s���Q�O����!�e��
:�o�8S��a<�Z C����2ܐ��p4rFIjg�8۵���3�rMgܦ�[�k9M��#�Cn<��[h�C��U�ۑ��G�Ky��Z�mŭKuն��kZ�y��,0�]�1��>2Z)d9Ԫ�:���/zbc�^��]�b�Zuz�'v�2}B8{�y�^m��y�����%R�E�%\�1��0���&ӧ�K�2T�^̴we�kr3[�93�cs�U��ĢS�n�Zi����<vU���A$�@,l�y	�ȇ�1E:A�Qi�ʵ��b*�@�d�^����{�u��;ζc���A�R�C�A�����"DjAM"�L `{`�E����<�(|-���q��`_�%*o���m��W�om����q8����M=eԴ�7Ʀc�����TN_4��<�OU��u�����Hb3<��WTҔ�fZ�DĖ�>���HNy���W⑖XMb���H��H"�f��[��@�J��b�&m�)�w����r����h�Zc��2��׼�T���c���קu��-�q�Է][kZֵ���(��)L'���y�.J�~��2_�*�8��eqv���yqǣ��kH�q>���{�3�l-��-)G Ԣf&vɰ�`�g/��&-�$�p�D�L�)Ȓ�	i�or�j2���m[m�Q�@�Έ9~��5У����b�iDPA�"=�e_��2���"̻��>ө��E)�����4�nf!ݳ)c1�n>�U:z6R]ӎ��V��6�)n��ֵ�k[�4�Ze�K��3)�a'��-$���CDS�'0g�b�J>	��ڞq�>�����>s	�9i���MG
a�O�fj<�d�����Ë��Rۣ컞T_�V�OZ����N����v>8f�Q@�G�.A�`�C�:�F�+K,��KH�ʫ��ۋq�J�SxOT�e�[�)�FS�>�D���X̵	[m%���m�Nf4���ǜu����bw9��N1S6�8�0������:���n<��mkZֵ��J%�Xa���W4��G�&�x�D�{�W�C�	���I=���]O_)D�m�!��xsI�0�����|��lő�.x�1o��B������>I:%⋄р���ki�YF�,>e�G�jǱ�c���蔼>�1s�������9�g%%��q:��1�/�tˑ�	K0�뼙�P�!���S�^c�N*5-������-���^|�)�>"'56�n<�[k����Ӌy��yj[����խky��KL������([�*8��]����3"o:��L Ө2�6'k%�):�5��UQ^@�M��������@��(�z��*���<�����cV���I��@��}L>��'��Z��s[仸&��^��F�s���]�Q���Τ!�B ���
Rg���CV��7ď�.����	o��'8V�d�2���9���'q�}T��\i��.S����i�3��ͫq8�[
Qou�[[�ʛi�yL�T��1�\s��� ��A��B�����~}7�&�0��%��L�Ҙb}�F���y�n��ڢ_K��%|��ws>o��>�8�Y�O��vŖKD��ijbᬷOvd��{����a��),o�5NF�}�UT^=U��a�����i�V�o:���V���ֵ��j%�Xa����z��3"^r�+⪂�������ӧO�n�ə��Q��!��,:��.�������J�Ә��%�,��Џr�0!9�����XfH����f��KJ5R�Q���䧌q�p�޾��	&�YVG�����K3�k��ba�6�yx<���2%�r�X����,��[L�Ԫ-��T�����؜c����v}0�Beq��h��Y����|�o:���V���ֵ��j$�S	����|RNEUUV"�"
���đ���*+ە\��*��T\��J&�R�UR��x�::�m%����Hy�`��/k�K�;V9��gͪ;q�Y}���gЈ���#��r�5Q��S	0�55\\m���QI>ˢǑ��,JK�4��B��,S#)&
P�#)}��8a�D�����o=�%�wuU�[/��'m�fg�D$��h��N�3��(��饮2D)��o	s�*��OuT�&q,c����֚*%��2�uی���L�53��n#8iQ��m�)�^i�q�μ����Z�Zַ�Ǆ�S	�")̐⪝������������ط��|9ٙiשݵ�&1�T��l�w��~9{o��aP�Wt���=V i3d2�K�7F�=τ�%�\��sE⦻q�#O�N��%�M��%<�7��X�c9q󯦓��^�e��9�̦d�uqv��g�,^����!�_�s��BQ{��%�2�m�
��n�W^�r?_�G�?��&Q)����J��[6fÎ?�~������h��|�t���f�ݬ��'v���n��v��uٛ��Y��C�w3:h�&�E�DD[D"�m4YD�m�\ۄ�e��B""&���Ȉ�mdH�"-	�5����h����4["kml��hM���kmdME��-�"km"&�h�&�h���m�E�4X��"Ȉ���",��E��MD����E����E�M��DD�DD�"[h�""�[D�m�-�D�b&��dYm��dM���"�B-�h�DD�mDE���,����&�4M-��mE��"",�l[D���4Ym����Ȉ�",�h����,����h���&��E�DD[DDE���&�""�$DY[h�D�m�����mDE�[[h��h���"&�"-�E��������"-��DMDDDE�"-��[D��DD��D��DE�""Ȉ���냫3�"$X���Ȉ��km""�!D���-��""�&��h�-��H�"�,����[h���ӧ,�H�H�D��"Y"[K$�f�iid�Y"D��D��I%��E��M-���D��KIf�m&�,�!-�I�ufp�HK$H�L�K,�"Y$��M,�Y�D�D�Y&�-��D��K$�I%��Kh��KH��h���Imf�id�%��֒[IK%���H��,H�Ki4�f�[H�KibD�#����[H�$�%�im"�4�ĚY&�Kib[Y��-��bD��Ki5�Ą�M-�$K,�$%��[Ki4�M,Y��-�%��D��	m"BY&�K%��H��"KI,��YE���jYY$�$��Y�iĚZ-&�-��K$��Ki4�kmi4���-$���4��--$�$��ZI%���-f�$$KI������d�%���$�If��d�KI��d֖KH�,-ZD�ZBZ[id�ii			i,�K$��$K%��5�%�H�H�I��K�4�D��Imf�ĚY$�d�m"�d�%��Y"Y"Z��M$�D��I-��,�-��-��I���H��$����$Ki%�%��%�8�8KH��ZId�5��m,�-�K$H�[I���[I���M,�M-�$I��Y"X�f�[I���4��,H�M-"D�,�-�I��H�,�H��$K,�"ZD�%��m!f��"D�M,�Kh�K$��	4�D��h�K$I���Ų6����͹�c[#5�6��ml������fB��:qn�JX���l��3[,��6��6�[b��[b�f�4,C!�2!�ж!:Z���CYA�	
l[BAhYAd$�Z5�$-�kBBBА���dBА[CZ��-		�hMBh[BB&�!Bi�ZhMi�p�H�i�֚#[M&��il�ܔDe��Y4�h�i���F�Z4�ɤ�Mh�M&�hMi�5���khȚɭ�Y4�Zi��h�h�i�k#I��&�[M4e�M5�Bk&��Mm4��2&��Mm4M4�MY4і�D�M4�MI��������Mm4Md�M4��Dd��i���Mm4M[M�����9��Mm4�[MY5��ё4��i��i5��5�Dd��h��D�Mh֚#,�&��&�ki�ki�ki��КY4�[M4�Mb2Y4�[MBki���i�&�M5��ki�4Mm4і&���ɡ5��4Mbh��Кi�k&��i5�Md�M	���k&��5�б��Ibi��i��ki�5��Mɦ�ki�5��Md�M	�FM5��5�M4ɭ��ki�m4M6�i�ki�Md�5�ɦ�k&��hM[M�	����&���L��4M�&��M4�i�kM4�[FM5��M4�M&�ki�M�M4[DE�""�$�"ȑm",��"�v���h���D�E�MM�,��Ȅ[BE���mDE�"�4L���-�"E�&--$Z",���H�H�"-,�$Z"-�B�kbѨ�D�-���"���BE�"�DZ���Eۛ�!hH�-��h��Z,��!"�BE�-�hDY$B��D��$Z"شDDYE�h�mdY�E�""ȋmdH��-,��։"дH�"ز$-$Z$Mݹ����!D"E�b,��E�dZ!��E�mmE�"�m[k"h�MDE�DD[[h�""�&��""�"�[DE�H��-�Ȉ��DY�4H�&�h�m"����DME���:�p�&�h�����km4YD�dDH���նsDD""E�#���"�m4H�,DE�DYرE�DX���-�kmmD�b&�h�YD����4[""h��h��[D�b&�""h�����""""Ȉ��dE��!D�m�4[D[i�m�4Y"-��mE�MDE�a�=���z����kn��sg��{[�8�tf�4�1��m��;�>-ϫ/�����z�������ܿ��$Fؓ�G�j�����w�Ǐ��_�g�������-t��;O���ݸ������?�;�}\�?�n�ɺ��{���w���O��b?����_�j��D!~���|����������ׇ����`�#�?NCfl?�܋H���;>���o���}�{嗃��g˭�|��n���|G���/�I��|����|��lͅ����o�~YQ��u��c���s3��a�_��W���m:�~�o���9����?��6���������s?v}��x�����n��w�R����ϣ���V�Ú6l�s���m�A���3n�833�cmƍ��o��f��(͋L�go.�?f�g5���S9�7_��?_g��s����ϩ�����m�! BLه�6m�FٶP���BA�BF��Vy�����ᷭ�<|�������7���lϩ�;9�����q��?o�ߡ��}���q�l͇Y�n\���߳����m��-�����ޑ��W�����;����f�m�?v���n�s;7�e������A�~|�������_������7�������~������y{?�~O��h|��a�l;���l͇�����������~����MA����)�_��>v�J!M��d~�m�}�n}�J_֜�c�o�t{Ͷٰ����x}��gs~���D�)/�B���p�m��y�����u�m�v�L�m��ޛl͇6;����/���O��ٯǾ<}�fl>�����~��7ѳ�>��1��_�����|��{����n�-�l�����_�~��s>���7��k���ɳ�q?77���o�o���|�fl>|��}_�n������6f�Ѿ�����_�?���6��^}O�����L��o[��_m���z�i���?W�������Uۛ��5�7��s�G��e�����W��^�c��ݘ~��Ȍ�4FQ���6؈B L?�?��m����s����׾f���q����龍�ߧ��z޳�g�Ym���<�vn�7b���������?�>�m�?񭟻��:}�zM�i����g�������s;m�~��~~m���ǋ˙�>���w����~T���1�F�=�Y��������)���0