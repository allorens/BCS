BZh91AY&SYZE���;_�@q���#� ����b?��     7��ke)�-5
+jHj4h,�"����V��5�ֶ�ձVb�4�eP���
��UD"kj��bm����c�����2�㪊�imT�,�Y��jͶ��jm����k"��m����2�h������-�
�km�%V�f�[m�0m�R�F�AC��o{Y��EU��f���l���Ti�P�ѫi�m���х��k%5fѳm�V֭-f���l�Ȫ�mQ�mIIRmL�dm[k%6�Z���^���Z�  �����5w.�T�n�@4�5�.�Tv�붶��l�t��R��A˳vb�l��Mm:�.t��u��:��#���6ک���ڛAZ�i< ���h��g4�u�-�\@ �up� ���l� �v�h�3�@ �8CCwK�  �{� ���T�ԱY�ՙ��n   so  �m�{�ЯE����z [�o@@t���= �׼  ����zL��  7�ۍ�4 �<4  ���MF��ٶm����%k[p  f<�  =�o/@
����z�l���y��p=:���C� �{� t � R�]�h �5  {y[m��diV��jj��Kf�  ��  =�� �� �;��@����`��  �w : t�  �nֺ�t�]�P {s�-�Ih�[�Y�"�  N�t u.�  ;���T]�ۇA�n�� �;S�G@ݵ�  �������� 	ӝ��a:l��D�k$�%l�JR� ��   ٠�@��8��۲�4v�W �W85 ��h����(��`5Ѡ�v����k6VV���@���mx {@ ov�  m�p ܺ�tkB譠 �k�  [�8  ������@ 'F
 ��*D�%l�eiF��[�� �� -��  �X h,�8�@(� Gn��ѠS�w��-���� @=a�z�4�Ͷ�j�[�Z��ex ۱��c�\  ��� °�F�4 �j�NwN ��\ wa� ��.� �    
 
j`�J�bh` 	�` CB)�)J*���  �dhb)�1	J��      "��Д�H      %4�b����jiF�H�@4�A�A	JQ(�Sjd�I��F� �����r�JS�l��0��R���Y�֬�Z�|�~�^~x�z�g����=}��
��@U�DT�
���$PW�O �����?3��������ڧ�A@X?�UU��<"�
��O�0v��Ȁ�����~�/H��?�f���(yaс?F�,	�*�:{p�d�@�{a�G��}1�"��=�/l���W�;g�+�
��l+�
��=�l�l�L���{`�S�D�;eN�S����/���{`�G���=��a���|2�l�"��a�;eN�S��;a��v�=�'l)�
vȝ��l��"v���2v���;e�C�P�;`�S������=�'��;aN���==��W� �<��l� v���l!� v����;e2�l	�v��l	�v�=��l	��&dN�G�T�{aN��A�=��ʇl�vȇ� ;dC�ӄ8�vʽ��lv��E��
v½���x`N�C��xȊq��")� ��
���(�v� �{`T{`T{a {eP{a{e{d~0�=�
�����N�D�DN�@N�U� N�N�N�N�QN�N�N�N��"�� )� )�
)�(�� ��
��� �`|��>X{d���� �Q�EG�QG��G�G�AO� l�� �;dN��P�;aN�G�����(v��a�C��;e���;e~2vʝ�'�T�;e�C�A�;`N��l�l��@�;`�C�P�;d��7�z���v�iM��86�>���(����2έ��5���lɸ�T�m=�[zh�{0�m{3.���a����R�(�KwT^;�&6�ͽ{X.J9x�T�Y�.�Fr�)�b������e�с
V��W1-�o�%u�)o�·�����r�,&E��k�-1@�3^�5��d�4��y����M�u�
���$������r��C0��f��J��h�R=�q���ʵh�9$������D�v�]nh�F��4^5�X�?������r+�P��fkI��#s�-؂hr���z��6&i����!��'b h�O(�	�@G%��S&���H��Q)4F�R�Ue'��# ;�J9uc���7�Ɍbք.��4�w�J�]�Sd�z��ֱ6 V�M��ճO��:��e%C;v��^��=����5��V��I�WD��i�f��B�W`�J�{��WZX�H�E��F�D&D�3���^C���.�^�feH*��
޽����	bcJ�2�,TX.n�C
��	�'_�[�s������&�v���)��;O;�-f��{��%����\x�*��l^����FD����ɢ5���DˇW��Y�M�7(��P�ze��{O"غNR4�xB5d7��mۨe���7�y���X(jÔ�;
�r�C���d(2��mѩnVR�VM�T��r��{��&��i�9V�&���gB9m�Ay@-�3���"�=4h��M-�f�q�N:��3n�V]�#vԤ���ȸ��!�L	�Ǵ���vU��}#�Y��c��;`A�
�T�&��Ks �3��2\�7��1�mbș�(�"�26���Ko��XZ˰�-�K���I�]7A�KI/mU�A(��gi�(r���l��;u�S:��t����m
�7k4��� ^��0Xmڑ�Bv��b%aa���F�����֘<�`cھf��1��jir<�x�t�-�ǝ��t�<��}�5�\i2�%���-�8W����B��X%�в^"�+��"1@8]�]|4�����+�kF%V

�ZF��0!��^"���i���'��"e[7#Ke�v�@W����EǱQ��C�Q�Bᣲ5 )�*ml��,'�N��w+x�ڱ��#��]r<z���y,�)\TCyme�F*���c �t��{�j�a�l�u��X��}ʅ4	��S�Y�Y[N���XKJ����7w0�Uck3���޺8���i��An�Y�#�Kn�Yu�56�sưX��#j�̚�]�/5��$�Y��y�cJ��Zmͬ?dykL�z�RZ��Fh	G#��#d�v�e�eRt�]���̬b�gmn��ݷ)s����mif��w�mh��m�Z���)m�T�!8ۭ��f�a�6�L�)=
�!�f��n��֦2E����j��n����
9+V�C7fv��gu�@7{G��ۉ[����x(L,m��[.YP����[	
��T�Mm���(sw����� �ʌ+��w�J���s&17���8�OCQ�qҲ����L�1dIƶ��!����x�s�4�պv�δ9��8j��6�[��+!rE;X���۽�aiyy���U�n��a+tt��#i���["2�@#j�W��Y��^^R���V�VJ�H�(EMX9��F��%$�n���
4�@)��kx3@��K^f!��i�,MS��N�q=�[���UĞ)��&Qy�b&���]I1ܬ2�te�Q�Or���t���m�R��j�V��t�������x�	$F��wo(�27Il�{��W�F� ��l
۸e�Ef��VZҨ�oX�[�]�� �݃��n�#C[����u^V1�^�%L�Nc���4�©
0EbO��V�EGr^��p2��$51���&?���7el՛��i�:�Y�i�i���Įb�EiZ��Y�5I��-�dU��2�� )�EC,�%N��滮��u^�����[N�!b1۽;����9E%�UՇx쳱�)
h-����,Z;�[��vf�nY[�����n��@lVJI^� ��7�j&f���jRtۼE�r�&��Jl�W� ���F'��m$���/i^��PSo��w5ڭ�j��@fm:Xe\���6�k�1+"��vq6P�{�;8)�jc*�S�%�*(/-9F�L�q���5�#�/,Ȭ�p�ǚ����2:*�c�(���A!��c�
�Ww��tȕ��h�U�ɍ�9�P'n��)ڣ��9Gt�X2놣t�Z���0�[�J[��S�-
'J��_7���4��\e㡘���-ѱL�l����d�r��n�v�0�ۉǘ�J�w'��HmV��pP6q� ��oS63D�ʭ���A�����t���gh��n�2ha�Y&
S4�o�ʺ���\�#�dl�vӁ��-65���E�eg5y���ݲ�)���#��;��L0B���Y�(Lq�տ��4�u�^�h�9��:��:6鋗���c�H1�D���ї+V�57v�t��7������.�]e��5Qe"0�v �2VB����E�r�i���X&� ۹Hc[��)n棊��ҙ�C4�螣AQ9�m^o�P��wPk���%}���OX�깗�6�$7N̽U� ��x-(�o1�m�2�S�	�V(c�x2�ˌ��rݝ��;)�RN���څ�/bԵ�,���n�}	��#����hnT� ��Gy�b8�d�L�E���Ձ��[���� X�bP��[b�7�Ld�'r���`��m
2�e8��b�����i��Y�X呡���·�ep���qug'Mh�B	��}mJ̭��d����%`Whf^T
�M��p�=��[���@��@=���WX�8B#:aeܺ!U�,�Vj� �o,�Yhe*6�,��%�)[R�l T2�2��m�RNe)�M��Tm�ŷ��W�%Lp�t���e�� � 7l��,4\IZ�o�l6"VU�����^*�E 4V���A�I��}	:�cn37��f��]U�W��;R�*�Hic�%!Tp%�s
�Ɩ�=���[��lj�� hp�������{&݌D�zLw��ؔz��0Gob3rS�S�5$y�a�2�h)Z�؛tssH���e�|Ѷ���g,6��v|2�"�`t{B��JONʙ��Vӎ�id=A�r��Mt)ն��:ހզ[�H�TTUxUmY!`�q]E�񽣥�bX���I����e�1pnٚ�wcV����߲M����mڕu�ѳ&<�b5/F��G$'�Qa�Z�``�����[�0���ԡ��q�+I� �5�e����Om�'�Ӵު��o<��֊�=�V��72M��H��r���91St[eR���,f\y�.9�{��M�*cX4�gu��x��d���0m��	x�K粰M;����`��y���a���C,m/�.��1l��={4;�+Zj�c�Hfި�M뭔cU]]�cz.[c�r���S��q����[z5Dd�/Rӆ��f��h�hWYD���wt���U�Ϟ�y��;��ө���h��H�����dݥ���� ג�V�޽v�p�[	f�]༖�"R
<�o�e��N\p�MKذ<�.�ӻ3]be�M+�]��2�܄G��K,�w�BZ%c��,�Ә)�[h����q��iP�tԪStAv�t�K���x�A7]`ycL�0U�����;9��c�m��:�I*97j Э�C���c�C��n�# ݤ�W5��ŕr�9���ce[B�kd��M3�q����RR�o1^��اuz���tMU�Q X��R#AG�R��i01*�E���w������WV������a:n���=O���@
ʓs\ޣ(U� ��"ΰ�	x�l�M�QP`� �S��n��H]Z)-���]5�����bÅ�paw92�O �`�J���9J�:�m�0Ř�[Y�l5o��z�iM��a��]�Yp;���˔���:�-�7S.	Y[OV8�^n�x�b�5i�6r�V���z�����a�U�ڃ�Y�Rz��tجͧ[u�3�1��4����m��.�v�š&�j�~�=���Y��cb��mY���JmI�wk+S���ƊȨ�E���(�2ڏ^D�_AQ�`XN�{q���T n�B��wI^-�
��D51	x�$����1���zƚ`���˫׋6W7cFݖ�ʗ��!�a��m;m�ݩj�-�Z�ݠ��0���n|�2��2��D
�n���e���ő����zR'2��L:õ#Y�=y��y/^��۬q,�nՊƳ
���7pa7B[� �O�BIO[&<�,��.�m<��fpJ˒$u�Q4EI&Dv��ѐ���]���[�#�'�Z��
�0\��lG16�B�[m��V슁݂�1�x8՜�S&�aa&T�wF;���;�2�c��GR�XM"�e;���%�e`��
G3D�\�61=PH�nYot�A�R����	��š%]:��X�m�.,�si�B�����Y+b�5YAE�$�M��c�kZ�cZ�*^s:��ɵf��լW����8Y�V��U�G.�\Y�**7�lC�d`B�MƷ���.��]�5�|Յk#BHwk]&��8śe$&[�vn�vib�U�9(Q����9HAZ���,5�3�y$��{��X7�����åoh��n0�����r��q�Ґ��i\�cT�ST!�mi��d�TJ��aH޳�!�ҽ�ZY5-ͻ�V��i�.���R����i�EYvM<��9`��ø��w��5ni��V!���c��Ib��Dmf&�7Ykki�u�[.����@ܣ2�M]e��52S'w�f�3c���z��t���꼷s]J�yl'k���mS�Tt��-RZ�2�˷5��K�UӨk2�nYS-8ӳ��[�c�d��k%��6F 86���9��*Ȣ�P�Y��������sU@l@�M"\�A�,y�ͤ7�K�d:g�=zolz\ѱ�d��Z!���9���B��Ū�k�hVI1fn�<DwGm�"�c���b)��F�Ƭ�5�x\��w1���(�,�=�{#��g��p����z��[�]�qY���Y��1�]���%���]`�%@���*1m����5�	���z�񢦭��������6���+��ڎ�5X��n�T����n�Z8�Q�h1�'��^�j���.�L)�*�6��4�6�V�8�� �;gh��t�^�ˡ�A�Z
KL�)`mV�UE����[��[)�+�����@X�{��v�*S(^$ ��$���z���Ea}k
K��Ջ�r�,��h+Z����K�P@J
+WF��^|�ƫ�n��Y+b����a�l���PUͧ�L�t/Bm���ZT ї1Pǔe#�3�uW����Û��֞�2R�P�V�7R�o>�0��~r�d���⩩F�66%NI#(�d��I���
��3>!�e[k�u�� ���Uܔpֱp�i�GY-�]�
�MT�̴��--�B^�Ĳ�GA�.�i�@E�@e��z����u��t.�n��غ�`
&�ˠTA���k0�l�coh�B�j�&��P�CǷt��/v�Z�����36��c����r��Ckl��(n�6�B��.��=ӫ(J׬�P��Iq�rnՙ��Xi��.l�D���sT��@�D#'#���h\�"G,���S-�J��� ۆ�i��`�8�;{Mf�-������Y�N�)�Y�#��N��cBص+)Ʈn��$z>܋��b�|�lP���s6�5�lJ��4m����qջ�ԪVu���bʹ1�nR�r�ի�b"��:5QtK����7��O�������R2�� �*8T�aK!m�aI2�-��:)����N�R���S�o*��@�+VۺR��91��A�xi5N�ܹ`�QV����/k���+q��
��:&,��c��'/*Ba�)|�O~�Un�U�m5Y�Mem:N��:��[�xZ��)Uӣ�Hټ��'bO]�ED�6�;��q��2fS����ںv�@�ʴ��kP)a@��C+4m]�^�%�,�����\�\�\����r�h����
,���b��%R��MC�z�9P���N�; )K�>ݴ��W)h�OA����$��
v�m�w[��s6�:�a=jֽ7&�Pf:׷���W�n��ҳ���D��"s*�]Y������7H�C�|saN�w�=ML�n�^j�^�GvmSUj��ގ�'1m����5ޡV�"��/& 1,���U��G֊l�i��49pܴ�7chТ9�pdI0^iK��t7;�ʶ
ۢ����12+t�XrIV�-G�Q�20-�4jy��	�Z�bf��kb��5B
Ӷid��c�϶J�v�X�V���4b�0�q��l�>t�Ѯ�a��aXZ-���V/9;��z�w��>�g�z��)�c�3n�Z���X�T���R&J�h�깗l�0�Һ�@{��ķ���y��e.������{���V�&�Z�JqT*r�hc�6Lt�Q�ᑉP�#� 0��Ӏ+�e�r;Д^PR�񳮇1�yd��I�+z�:�;��${���`�\�{������VGFݣܲ&H�Ɲ��&�W\�F*,�9Q��ٗb�bq��F��q=Uh��xV;-�n�m�פK�N����H�VQ��]�;�X��e�\��v�Кy�@�P�b�&:)�V0�s����W*o4�5j���PV(t�����t4XǕ�)8��t�aD�^��"�S$�yK(aRȺ�{L�t���?�Տ���o����O�/}���n~k�_����ݎ7R�Vn�[n_=����ֹ8�_Ayr2�PuݳX�:X㷕n��r4���iݾV���*_d�֤:oos���l���N>�ڜ��ƓN*3�C+��3*��S:T�5�#,�܎ֳ���F���l^4QI�w5�ui�e��p�B̗�哕�]r�(2�n���6��j��t�݀�y=��Z9�t�|z�mU��άi��;�� �R���=[w����Ӣ��1��pϵk�����TN�*�ևMR��y�񺾫��K�C):�06L�kή��3i)�C\ظ��5f��'�*]�g��M�s�̾�E��Mcܗ+P,�XUt�@��l�Vh�nA$wD�]�[�k�.�{��3�����O��N��Z�{�\�E��wXk��,/C����)���l�\[clkv'e��`cָY���p�XGoX*����+F^�N��q|�
������KU�`�K�\��f�t��t��\�2�3Ji��i�O�v��.�U�,�6�Yo��ܸ��L\�V��'i�|���YK�AVA5_u�hmM2���HS]7�l���.%]���'t�k��`ӨkL�Spm).��:v�c��bKc#2I�E�(�m ��ʺ0�d8(ڰ�1Tzvwc��1�v��m�o%$o,Y
�@�qݎWt�K����9գ#T��}�K�H�&3b�mGu��e9>�f�;���5��f���t؋�ЅN��%�g�� k����	S�V I'J��Z����zv�=p;�9+n�v��3a�TTy�;ȑ�
���ֲ�Q�F#S�[�
Q����hoU ���X�'�̮Y7C��7�2�B��"k�n�%E��i^��k�X4�8�u�L�f���մ֚�1��X[O�j��ʳ���-�S HdPVQ.]n�4�=���8U��Hh�'H��}���2��1.�:��yNP��Э5���ӈ���º����v��6����-|[y*��z*یV}}q�1��ޙ��dr�\�{-����w�3-��O;)����"�)v��D���-��R�p��K�M��&L�w+�,7���.��)n&�Q(�"c�Ř�*!;V���2�7��W�y}*����8���G��R	���{��:�!8Z�J�7et�$�����s��"��{�g9�-qo~�epJ��h��㽲b���9��6�:8��9xc�[R��\��m�8�X|�J��7���	��`u�W^:���U�iv�R��pg-��-M�rZrY�F���k��Eb�ߚ�55����ص���[F��reޅ����Vn��me=�늍v�Z
��dQ�2PYl]��e��IZ�>�����������5�h�VOe�+�w��Ric�U�^.��2�)�;حgf8ki�#� Tj�ü��|`e]�j�b�x�b��6)�p)���O$������v
�ܩ���'x
��j��<U�����ut��VMc��p��R;��R+�ͬ�����6� ��m��c�EvGH늆����)ٺiJ'4�Y��2�7�X�K۫���(N7�H
G'��qL�bR���Pщ��������.�t���y��^e=����jStu���{��[IN@7L�fJ����]d��;�g���t�Lfk�p���b��>4�^M�z9*K�U�zS�^<��]���ۏ����x8��I�_C��AK}�ĵ�N��9Wc�]�4�:W���f�m�˭)f\p0VeB�"/����"�Ư��ĭ�I�Tܺe_\Qdh.܏���u�l�l�Q�Z/�Ε��d�ڬ%J K|�ٌf'A�f���O�O�&(�L�)�V��V�1���ؘ���/�!AuA�\jL�	�(Ը�H	�����җT��wT�9�(��L[ ��iP���w
�ٝ�%�6��1t߹��oӹ��K�9��>C�\�Y�30�s�t�4B��[6�bǴ����1dޠ��&��ƺ�6��v(�5y�.xWfη���u���	C��5d+
���6oA;몺��M9Q�V/��\�aWyY2	1p�k0��i_d9G�2�WٰT�l[��fI�WQ�$TC,�bzjm[+h^��zWQ�t&[������y� �NժN�"�0y�#�b�(n̐a��\,�L_WZ��|$I3v�n��G����o��v�gK�K.��R�Yk�X+%�%����7���'Z?0�E^7V��=:�-��r8������דf����L�O&]륩��%���5� SbMr쁐��S��x%#�̺ٹ�_`/;�"I���@v�M��:T��:4j���5�IMtv�V�C3hvh��޳JR��)G��!j�yL�:i�5P`Õ�˨�3)�.y<�GϽ�J>ǯh��I|��C��բ�0K\�rW&��x3i�����l����	�I��xW�u
�}w����������r]�Vsq�71'|;3k��e�meҔ�D�մ��Yb�%��-�5��-t啦ku���niV,R�V]'u��v���ٌ���uǒ�=��K+�Ve�&t���N��x����؍iv�fG����f%�%�����k_fo�Q�:�Ed�x�b�F���8Q;����.Kk�$gjߡ��2,kQ۬-X�K�+9�o�VP�үl�4�T��3���#R�Y��Uw 7N�ق�ȓ�3;!�iJC��F6YAe�d*�כ�6�E9�jO	��nk�z�>n��"JȆ�,ɝ���X׳hV$�㮃��G�:�)
;�Iǭ)�.�7bu\(�����ᛏ����]9�6ʑ[��y�^W3�l!�w�(3s�HG�����u��Dc�V%�{�Pi��_.�R�9��&���N3Zw�s��ts�-%�j��u��7շd#[�g��G^��$aMZ��M�B�7ՠt�/rE@��t��2wP�7R��FC�wyK���t��@�A�6�h�U��3��P �����Ah��*J��j[ru4N�L���z��F��3����b�xm�n� v�5Nf�v'K�ٌ҆���]s� �<ɺu�x̼V;���+��)3h
�e�����tm�	E�lt9w�ܮ���y�Rb[�"�١�����VtIgWL����@	T�������E*��Av��X�A4�w��t�j�P_5ۙ�g��ge�j!���^�e��k��#J�b֯j���zl�ئt������|Z2��[>Y2�n�ULM'8oi�5�h*eX/�k�x��Ɵf�u�f�%B�����B�k���]���Z&�}'E�F��6�n=��5Wu/�6N��MX1���z�����5�e���'r��U�cqd���]1�Oc��9�3b�%Ms���l�$��l���!d5�)LjHt�=�J��t4����9UY��+8�j�ܭĶB�v���4��c�}�)��]њ��������bjG�,��m�`맮gT��a��Ub��O��
j�N�����U�e,�~V^��L�p��`�M9�S�f!�����<ڷ�`2���Iȃ��� �Sql�7����U��4�h���*#����ٺ��0�M��w�9Ĳ�uܳqͮ*=�5�z[���h�4�}��̤^5���Rn�\�E�*9�2�I�y��r�hD�y)΂�B1K�u����o&Z��-��ve	��xw�}��x�c��u��Z�eG��؄X-�+{/��q�Vܗr Zh��==y�'�fo��rKY�'`M�]��5j}�����G}��}�ͽB�,�hځS�6���:�r�v��}��S{1����H�'�LvT-l���8�U��<F�����$�^�����Q�]�2'����;'5��R��n	C�K樺�5��v��v�Wbol�����t�Yk:��p��tj�
�b�rn���`�y}�љ���k��]�']R����y�w��ѭ�i=[�#����Qʳ[K/p�# '2�9�@�Y����M�׽�n��a���ʷ�Q�����X�nlV�u��g���o�B�4��l�{mL�Х�9׻�ٖf��Z4�K�m��R��Y�y̢��b���M�t��hY*P�!��	���Kk�[rY����rj��,`��L�S7��!��q��ss�r�
�͍�	M&k�{���{:�&������HY3�U��nAB���u�$C�V��]�~��x��.���������������N�`X��x�dNu��HXm��wQ��mY9���:�H�j4x���l⚧2����a=����T���Ha�3c�~��-��ENk���H^}j�#�o7��P��a	D�oEڣ��a���E�B��q������Z>4���'bFi�af��Q`�.��iS�����ٵ�RE׸ݮz�ެƊ�gdW���ksV:*U������k�J3Z�t%����d���䇓���/���� �/��9�	�(��$j��Jk]u��ܙ�陛���R�[c�c��������g..m[Eu	j�q]��X�4ɆP�}F��J�Z���&u����\�@3ڷ/Gvu�����qrG�����}��DoV�lp�Y�321�#u�&V(�:2k
�3��V#�C��6,�[�?�oIҳ�������D4�ۉ���Xjun�y��^����R<i�;�����vst���]ֹǡ��a�qg#ɥz�A���ۍW;T�ّX�ʄu���`�y�!��7��.j����p_ٰ���R	P����&)\�e.s5s�8DP7�S�Y�@��{�#�*u�u�� �[N�w�ς���U��˕�R���6'����l��1he��d*nJ �>g�a�x2����0Y̺��&+;�]e==�"�����n.˧��i��Yo���*mPMLw�Ӵ�9��SQu>f�UaQ��]�W���]x�n�W��jr�H�k��VFM��ξ���O�ҎAm<��se�;�^Ʋ��/�%�<Uv[\)NDݚL�Z6���w=��r�rK�nٮy&룫�#K���I1� ڝ�2Zp��!mMj�z�V�B7ym(�x7!Y��IѺѨ�A/����MKl���B����2𶆳��s+w$V��B�	ɘ;i���+�tE��\�iS�M�
�vp��U��,��@"	�e��ͩi��Ŧ.wk�3�5�ۇ��c�7$ʅ�f��L�n�4�7��R<���O�wJ��%��\
�ɸUn#Yc�ߵ���fg;�B����\޲TU���%�&�3#Yu�A\�kJgG:+N���X���*�t -�@M6��c�H"V��syX+v�(��Ͷ��%�m��{p]_czt�T�1�VIp�j�E�YH޽q��jC#��٢31j�%̣]S�n�^�U�`m��i��Å�47ڬK��]�0<J�u�|���:5��ƒ!\����o0�#@e�^%.Q�{ ;�y����4,�(
yv�M.}�F�)Tśғ�CZ'2b��F�ތv(�{������u[u܆'� "�-=�dI̮����qX���"V6�C���{u*H<J��s�I{�IC�}	��L�V��O�`���Ţ� ;��N!�W�!C3n>ʶ�>��7HCv��e���i�%���P!�� �<�m򥦆e���O��]`���ix����:B
vuh{K�w�#��E֌�Cc���4���[Or\��$fQ˰"�3�s"b�ׅPsfa�/7]%զ�N�Dڮ�&7j��C+�(nb�)#�yK�%�ˁ��D���@�s,j��-�x>�t^u�X07����z�aKí�!ɶ�C���ӣ��]K+(mAn�R+x�ΚQT���/��3�r���2�8��=����wq@Ѱ�Пn�Z�k����F�:�}*8F���ӧV'cz�s���]}1�=�֕����9��3�Y"A�vwI��(
[�0��T�rO;WENֳ�@�3�n�R��@����-�2��6��A]��y�a��VF��1�P��n�U��\J+(ɘ]�'Z�Y|�;��5��w������H�ɢ�9�*N���-��r9B�9���ڝX�i����"��LE�[6D�n��|���X.v�����q˨$-m�f�L_+N��T()�v+C�ה�T�@uk:c�P0ێ*k�Y��L}G~\2�dom�3�U].��pW����X>�͏���T	t��2�] �%C|m"������6��͙����֮͋�7+@��	���Z�1V����/C{ʏy;��@v����tN����t�5��FN,�KOR��Rr�׶k�6�ZeefQs�W9�:-/@W1���t�֒��w�yj5u`�����g�R�:3��m�:w*3o/Or�c�22L+f��{^료��]l�	\,��q��^ʓ�GqSt1Q�-31�׽�l�L��(Y��ЩmWv�w�ۓ��X�ξ�>�=ەՍN���>�S�L9l��9��$����� ˌֵ"�騺��B��%l�"��4�$�IR�N����*]!)�AB�����[��MR����)�/+2]*��ˣjȇj�Q��肶Ȁ���*�6�?*�v���&����T툌 �iR%X�;*ˡ(��i*hF�eM4)�d�A�(�Ii� �!Vp;$�����E��1$���H�i��%Wd�@4��m��:����J�B5a��-0��V#�	�l�lQ���5�K�	�*�x5��!]��橡H1`���h�ЭLU�A��FJ(?��8�U�u>�t�Nh�N��j��_""����?��xP��/�����?�HB\����˻-u�k���@�M0|+���H$(`�'39v�����c�E����gR���]ٱ�-$w�����F]@!���nv�#r�U�Z�^���ۘ]N�@T079I�b[�3l�6��v/��)I/��<Y��ޝ44q�T� �_ڔ�<�}|�ۧP�I��`�yŐN��d⥱Wd��u��)p��J��ۭ�RI��;�Nh�9��7�����g9a$��c�oH��u�xK؜6/�{)av�{���W�<��A��z�;T4s�\�q�vb7ƺ373eeo2�����#L�]f֓Sr��*hv�o$��-�0`:l�[X�fk���q����=���Gʯ�n2dPms(�q�i��=Ȳ���'�k�^'�0��Sxm<!N��� ���G)ew	|@��YO{*M)�wC��Wh�00PyY4�0�xG]�/5CwF9��.�Ь��U�s�k�y���%����RVc��KԸ�UQ�B�u��������îD��ٹ�A<y��4P��68a$�Ѝ�`k��/v��������&�֋�$ښ7��%p7�uc�j4i�$<�����m�ʳgx�06r2S��="ԣ�ڕ�j�L��A���p�x�
�uD�s�jҁ��(�(<t��3�=}.)��w����z�4O#�Z���3���:��U�G�v��Cnf�P�X)��>��G�����W#��ʅXfN�3� ��A-���R�pZ�/b�)��u'(o���7�r3���RX�]�5h���t�Q��:�ݱH�]���P�퐅K���r}|]�$
h�ݧ:�ZWv��ۧw�J�\sv���{Z��Z*�ǗR�`r[
�IG+��:�*��I�;��ACt�]�����>4�E�\�U�7	޾�`�}OuF�+!7w"����&�����Z���7WJ��>��$b���P�͵�W�ХPiV]K�D��ث��b��$7�%�S�XU	�]���n��ʍ1&a�p�rۛ���2��4�!�N���^��\('�=�'ѮOED����כc9�[��v�{X�)��[=˭3�9��9Ե��J� λ-�	���:��` m)L��w7q=w%]:�%.�n�vY��V���Υef�"��#��U�IK/@ TkqM����7׊���&�X�*Sl�goV�	��,tFU�HW�ꥻ���^0]���h�[Z��En�K��C����[tm��cz�x:5�R��&���ҵ@�+�f� ���쇖�&*#�l��E�
�a���*��ܢZ:8oh�{�Ju�������S�j��E���'U,�\%�!����bi�E�J
�� �
Q楚ӱX����L]��D�fMɱ2@W���u��8��t�?լ|wAs-�f����f=~��3τ�,ⵚ1���mǂ`��2������(�����RF�Eݷ����C�5&wҖRaf=�P��ǫe�|�9v̬3pJ�pP)��� �`^��v�\�q�j�վ�L9@t(���b&Dm������9��{}����M�D�gz���.�U�s�Gq�3�3�C��o%V)���-���:'^ � s�I>;
�&���IƱU��X��U�Z�D2U^�=����ǹ���㜺9Hl�KY�j.�9u<������h�0k Hy^�:�[���kU#��]�Yk�B֘P5�<w��b۵CWwI�0�&4�n��8��4;�$@	}6�w������؉
�l���d�v6叝Ӿ%�����\Z�V��Ҽ�����a�a��!�[��+�u����U��yJ\9�5�i��R�GfT���'�o�Ő
ϳ�R_jU}�r�=��;ne5srt��t�X�io�LJȹ�+��%�ƅ��ܾ�;MgV��%�C#�]��Z�/�t8;��v�h�O+��|:�WV��B��8Dږ�������Ӌ�c��8�/0cAۡ�ݗ�u>�� ��f��ui��e[��2�(&)z ��ƺ%�碆8�[����(l��}�i5�v���HV;���%U��-�7�;�]��s&�j�vv����T��[x�(�r�Y�GH��W%![�S�w�Z��u��`�)D(Sǝ+h���Պ�ĸR�N����'4k�:*8����^n���c�`Zr��ep�F��0����X�xχ��.&\��f�K��*�AlJ0�h���m��Up������"�	�9l��n�l�F�6��P/i�X+��,�軱�n!Zn6��+Q�]���j���v�͝f�ԕ2ި������:�B�`*e��<,L���(����[�� �,�#���Uݔ�:�bE��&;g&v��<0�Ŧ�'p��-��$>��r�Qy�v�*PtV<�6��wC�L,��	�Nrl�k�Cb����1i�Q qf��-T�fv[�͕
���U%eTe�`��Ô�e�Ul ܝ)�e�s3y��U�{D�#�G�s���ӎS�r��/�T�;ڪ�OmZ+��ni��+�-��g1�Ϲ�-Ӌ��]ISe�wFe�5y8�˕��GdMiaܝ�<V�$y��m�(U��Z�aSW:�:�d�<��[t3^<�����q��j�o�f��y��:ݷ�!,-��^�uv�^��Fb��V�W:"`L�}V���:͎vR���tg���R�ya��ʧU�R���e)��M�h��]�� B�,]�<�l���ʽ�#+kh��w�V7������b;o��J��j@���Ë�4�J	UX���_h�[CB����aL�42��c�.����f��پ�tXZ����/��	���Ӣ*;�/������^a���Q��)vyڰYhk]��M�ZC�Dp�Z׆+�AP��WlB�oP;�,7��ZԮ;�Q���ZX!�2#��ה� `E�VQ����71�7&���ԓ`�������0L�4��[�eK�[@gm��7��h�\���;�������o�iKn��oGR��2�;�>���:�����ӕ��y�đ�#�� G��\���\����(�޾�g1��w+b[�ٺ3�ŧs��fVݶ톯�a$L�6���C�sm�]���t��D$�͵�@��Ta��)��ej�ZB�M�K�Y2�y�]mT����T��*\��������e��l[�U�	�GA��sQtx�f:�s�t�V�JR�.�����F�5� ������&+���f,^s�G��ֲ������ǝy����񙃫��{D�y�5�"�v؄͸)����j�r���Y���Z���:�@Z�e�N�r���Vm��虌��>ڵɻC%���[0˾�;q`���)9��n\j���w[�ۼ~N���C�����P�45��3j�Q��#��e��9��}}&�[���@3a��ϗY��q��
*��ci�u!#z��f��M��j���:+]�Һ������%Q�7��W�-kXA8sQ�9t`��:;������Č	c6"ý\/��n�7w��$:�4�K{��������=���j��gY��[8`S��pđ��J�c��QңO+D�cg���pTnY)ޜ��7h ��ɔ'�"�%YJ�b��r��19�����Tu{x�to���:�O�� 7s+�1�m&B�K���Kn�^�����g���mj&xm��q�`x '�'��b�;�ꁊ5r�`���s��^�T��z@�, �	12�ZF����hAv�-�������2;=��G _W.Uu�(��mM?Qzz�����z�sM�&��5͗n��C\�*�t{-������f���]��p.�/S��X��˵|m.<Nd�NU���,{;5]XU�N��;�ST����}C��b�5�K���z�k��Am����dz����oj�Srx��� ��R��i�U�Ѿ��umLwx��[F��1w6���o`���f}.n�e�]��ᡜEsJ�W6�f��=��b	7-K5���v�F��/d��t��E�q][A_#���A{�շV�-����f��f��R5;)ʜ-�\�*ԥ�F��ߗ<_�r�:�^%��W	%��^:P����l���]*�8�b��=Z3\
�F=�d*�3���;���bڴ�9b��RT��������	�BW�t��%s��=��h��Y�@�A:�E�Ӭ�J��i���)���	v�Z.]$�k8����D��{X��F%Z�t[s:�(��M�J2�놋T�筃X�����%�/.�i=��o]��kTCo�,�`/�k�Éup�0nX�hŽ��+h�٫�X�ur0�V֦���d0J�m1e��]s�]v���¢Fmq��e��b�4�N��9����������pV5hY�����ؠ��:�d���ko`��*��髡jT�T�ӽK*T	,���ޥ�3���B�͛d� �QZ;f1LGr�̽R�ʙ)wV��Sf���&= ��⫎�Z�[��*�5�xw��7q5��R�0u���R�`���'/������[v3��I7,�E�E��F˭ڱ�NfN�J�gd��MF_k�������X�ej��1�7��R5/hQx_:�S���D<雷\;�v ����)t�\�&���+S[�k���nR�w{W���55� ;ǝ�v�1��R��v�h�T5<X{�����X�(m]m<�0��."�u]�lQuG%%�ۓk��.�mp�Q�MYwfu!Vr����Ε���K8��ڦi���RV�W7�zr��
/��5���h4��2��ꫦ\6�vd��0�%�Y�N^<����w��r�3�l�C�ę��-��;��}��J���)U�[ov�r��eG��j��W���<��1���5���|\3J��*�VwVS��ŽI�h�:J t�ܸ��#:�P�����t+r-yحGL��[F��|������l�n�Deg8*d���W4�
1�kLP(�s(���y�o(`Ǹ7U�qA���k��\���8�8����s�YcOi献�pj�,D�1�񎒳e�����j��4:�ZBf�5�O�f�Yne�ZΊ�ݥ{K)ˣ�ve*B����0.
�����a��B8ň��T���i2�L�Wz�\�\7/igK��ɧ�{�O�Ý�.�w9��P������S� �V��	�M
3����*���)Z[oN��B��E��
9�XΦ��9#���Jwi�r��Ƀ+:U�!�ѩCGLr``:�i���ش����љu��B�n>E�x9���u���[�F�mWYT�+�
�X*���_MUj�N?��e���U�U{�KK�F}c�zr��i;/�ih��$b�uw�0��;���	v�`��j٦7��5#�լe��Y`��9
\�V7�ۿPY\�J���ʶ�,7����Pa����s$����4pWC���5ͫ�m�Ԋ��sl�V����F��=�}h�M�:ֵ�OJ���D;�F镃^���.
��v���V�vn���yx+���R;�9�y�y�:��"�����Wd�|�R��b�B�B�$V�m�wڞҽ�9��b|eva�n�R�*�G����)F��/���w|�I�
�����f�ɍbŻ���]�uZO��Βt������
�����5lt����j!+D��>�h���Yb��	M�������jR\o�:�&��c\٪��V9���G\��6���9�v:�0h��pG�gd�b�v�-�KM�h^'���&t:,kykT�1m�W�n*���U��f��k-wR��J��p��%î2�X=d�y�M����⹄�S���%D*�c۪mS�M�/�+�ꔥ�n���r���P{��q�[F�?=!��̊tٽ��n骺��a�l�:��6�t�ݳ'���|\b:�q[,��̋�oP�5�,3yi�j���ҧ�i�)��@�m��}��Ԥ�c��q�>�G��Ǧ�s_!�£�}vy8(#�����V�Γ�ӎ}����}Cm�ѰK�N�D��{B�5�&:]�VVk��{�2�A�C9<Uh�t��Щ��*�(�Pc�s�d��c�B����Y�1Vn:��x&�ʕ1n�wt���93S}RԤ��xo%*ؖ�U����H.�>���
+�#�
G4�)e��͛����ؗ��R�c<7�a�z�M�à
�U�(���<�[	���1�/Me�N��ݩ+E�I��ս"��ã�/o���я]�#��I�@�I�}�R���JSF�:�	�7V�A�+at�����s��X�sMvKΒ�n�y�eo��R��1:Ս��҈ݰ��%�N;	�nӥ��셾W}Zjc��zГ��g[tm�*R	�^2�zCY.���L{jX�Le����ma��n�v7�s��wΔ�s)�:��H1���Z��߲Z?v�f�DBvVޗA)a_a�p���u[��e��y_Д�/�YQ#�'��-ҫ�ر�T۳���՛K1X��I:�M�KG�'�W��G��P���j�8�ጎ��/�#R��WR�R�Ŕ5-u�7��	�� U��o�bn��*Nu��u�V�xq]b�x\͓���(��V�L�m�1�Ri�s�U;So2��lc*�u��N��S볒�i��x�Fb�%B�q��K�}��՜-���Z�78S�Am��=�%�Hҕ%�s���C\�$�T��l��sf�J�M������m"�-�i:�4�R�P
����D�����br���O��/����q7R�*���oii�L֨ 7f�Ϣ��ugqb�9���=��ɕG"��Ch�F���凃ڮ�{Z�"վ�� $��#�˿�N<�4���?��?���W�k?���======?�����������}|=��&�k�vSVh���?2��^;���[G�j~����Dyr��4������"̤7�����S*��R��y�q���NV�{{x!}3*ڥL��Y��S�U�mKX֜;�Hu6aJ�4{��\b��Y�$�6Ka���'X�Gd�w.Z�G7��V�N�C;x�Sc�s�]��:,"6�Cz�C:��3u��%�_E�N7�t���Z	PW4�\�Q�|2�me�<�;c%�����hk�h�nf��٩m��.t��>ŕ`����"��4�d��5�����v�T��MJ���uh8��f�8��QlY5�ifjӝf�l��U��� Vf�Xf,T��c�J������Űp�q�3r��₎�Ď��Y��\�R�L���N���wm�NZ<��idĺ卩u��iT�]����81i���9{H����ƶ���6�`Q-s��Ο���]�vQ�|Eh�k�/L܃�]ҫ8���tD�����n���Xj�����,ȡ��n0�v�f�JK/;������p��5���)Z����������]n���ƹ��F��Q\h\rh[��]��vo�3�B^���c���H��VDώ�ź��͡��9ef����sE �5
�t�$��G�WqC�)�	�~q�&��;���/z�� ���b��Bu�T�{GTQ���B�pذad2�a�9�6��n�X~����7��IQE���#��V
,	{��׏\�o���׸K嚨*���+�h���$)q�UUI�nC��l�CAHR77.��LTST��DZ4���<#�rxmʹnjM:�T��93����4Z�q���C��ƚ(����V�k�"�h*����&*d���C��5F��ri	�h�X�!y�r�0TD$E4�M��E͚����(�E�Rs�w0sj�*��-�EE�����*��F**�h����
��W��M[A��4L<�檹�QE�\Ʃ���5@D�r�5TF�Z�DE��DF�2�TEMQ�uTTRM�M�"�-fi�����q�3�0Tl&�j�Y���
���`�j�9����G�>5yK�����=V#��ͬ�@>I,�djso��	`Euvf��n���5�C����x[�����Mn�l�Ļ%c��fՌ�����>a7��G�B���*oN��REz����5�N4�
h.U�N0�st�Xj.�@���C��w&�K���v�M�9U5���b�o(ɢ7��y��6��Dm����x�^'���'Z�`�~�����ʸ�+��j�oE�$��#A������$��M2#�3�i��Ǌ{�
�=U�f�z�Ьq������nMns�dz�b.�!����_N�{3[�ᦧ��ɐTL��
���}G(:���0��].���w�#<��;]GhQ.;�ǼyVX�[�/�ZhW�-��[Ou�]��x�~Fn�Y��Zd͊�(���U�x��^����?p����F)~u{y�p��w�a7��v�}Zo��у{N������;i!�2���.�y�#O�:j��1��`8�{l��e��7�Nؼ�,�ĝ����,z���Kr�%
����=Q�)�35l%7SB����2I*��D��=6)|���� uq�nDqc���@l�&� �J�_ҳ2nhE�}�]�,��.����}�+�<ǎvی#�4�+b�A�+�͵Q��F�V�ݼ1<�a��^��~�WN�������U����G4 o]����p���~~�`�r	���v�v��������W�Y���q�%�#͹*y�ן9%mIR��yt�^p�^z����_I�V�g��V-��Zd���عr5Q����o9��u��]�C@g�'3_e�5���a���l��[/w9^��>ˊ�����| ѣ�����/�*��TἎ2Ϙw#o_��쎖�S���� A�hFDk���z���7��q�̔7"��>w��%���v���������"����N�_y:���ͳ��nN=��Y�Y�O=�����[~͸�����%����U,�0^n�n:fv��7e?v�/���k����uG&��-���U�Ֆ��W���,D�U����'~�Ч�ޛ������g����}>m�T���KoS�6�����jS��x{���C3R������:c���I��`-�Ye�Aft�ԩm8�t���c(`[,	w85S2��-b��rA2(����z+<��I�V�CR��{�6MS��n2�܋�#��|��ܗ��
���l�:�b�sh�"*��c�p^h6�4t�������xu���u<Ǹpct��1����֛l���ö r����w�^}�za>ϳ��#��}������ ���DAo�.�bR�1uv�W��z��MٵS!�ޙ�Z��7�Z��c����8�/=;�ʧ�[�r�"����c����5���jw���{�{.:^VoI��ީ[W�s���x��u[�F��[�Z�����iC� ���K	]X\*W����J��%xMڒ��1�u���S ������S�~�J%����/^�����yQ6M��\Ϝ��tל!�l�w��G�N���@|i�'�]n��QU]��y���}��+U����입7�����{�l�Xr��R��KNv�de�F��l�xcvվ���1/e������Q�Rei���N������U�:�����毚�����G��r����)6�l���õj0l>%G$V�gZ�.Rɵb�c����]<~o��5ى�V����.h*����Dw�"�=p��v����g���hzz��m�R��Yj���w�ެ^�h^�B�C	���B����_�{�7�=�����EQ3�׫��J]���?7��-�{��h�8�m�c��Wt�g���{dZ��~5N��'rk�-��=ⷥ��Cn�{���b"���O3����:�����U3��ο:ʞ��]#ޓFq�B�?GG��Dxe��f��N�ƞI����ͱ=�Y�}���s�\�n4p��6���������G�-��yl����73���k���"m7�m�S��^J�Jok3�^͑{+�|#�u�d�$��G��;ޓ�^W�7.�K�
��+�b׾��
'5y�mk^p���vUq="���P�����I�U�}���B؛^gs�R��m��pѠ`�.�i�o����>m�j�T���_�l
#���gުU��+��\I��/zw���N^)U�ʟ*����H�%6�t���u�߱�����Fbyo����}ɡ�C�嘺�1�+�<��Ξ�T���^l.�/�U��Su~}�f�
:�n����*T�F����R�m�}�W*`Ω�י@�sv�⿨^�Y\���p�p]M�tH�mNY�����C�MY�{ꃾ�+j{����Dfɒ�ˊ������ٞS#�4V��okY�^Yc�T�F`��r���-���Q���������`�y�g9�UHi�~�����t�r^��d����H�����{_�7CvA��ϫ�w#�e�kP�ν�H�!�l�]���W����R\�� ���c���~kΫ��
�e��w��h�[��������x�|,����y����x�4 �U��UB�b�!�#��r|O�MI��=�U�Ͻ\�	{�8K���i`���Mt�{e�B�W�^�@�v��Iڤ����|�&�I��}v	5�_��׺�'���9OS���4+���x�]���o�y#�T��=�)�c��][�q��y�K`�r1����O{����oH�`��9\>����C<�����t탠p0+G�8��l&.qN��e��Ba�KG�t!o�H8X�7�橴�utHu:M�6pwm>#�Ԗ�я�=[�n9�q�K�
.h�D�SA㛚ʢ��t��7���e����u��Z	G��*�6�}�^�t^��g����{�{|�{�Zʫ�qo2���dR܁�>����<K�q�]䖚}��)ʒ��OL��~ίs{���u!�߼�z݅�H�5�kn��Z=WN���X�{�{;�`�����=��~�i���q�6�(�L=8Sݵ���R���N`��mU^������Ng+}�^��x�r!��4jM���K�*�φ#:�מ�T�����'��u�Jz�*ߤ�w�2����깕O,W�*3�g�b6��Ѹ�:��?ws�}�Ƀǌ4A-�+?Tϒ6ܔ��YNKʊ�]!�����g������H�o.Z��VP�=��זr�c�2�y�ot�XQ�f��:��>��Z����ޕ��p}��J�Tdf��l�.*s�]�l��ǳ���o=��J��d�6�i��1*�׼�6��g��4ܯ�=^����3<��Ֆ ��R�Ԋٙ�|��Vj�g]sT �iT[,��=��g*nKv��v���з���۶�H:o����i�CV� ���,��'�*u�
�/�ޝ1άz���Ca��L;H
�ܨGFn9��r�I�e�[��9�}ϲ�Y'eނ�3�Y%���o�n|J<A�~�s�Y����*Ϙ��o��)N���F��[x�2v�|z�E�U�۽�6&��� 1�ܞ-�G�c��q�xx	�I��=������{]].�J�G�8ż�g{��j�Բ��[8��_{��Cl�����_Hm�s���c�-d��3;#���;���^Ȏ/d�a|�|�d�?������u��.+�c�0&��[�#kɍ����������u��u[�j�E.:�ݝN��5LpU����� m�a9l�f�n��OxGOw�퓛��<��D���U{�v{fer��K]ܦ%9�)zmVsw|<;������=U3�|\���7]G�����a&\�r�d���,�>�k���E�N�9q8��mN�t��}0w���qRg�G���m���?C�Tۇb�u�6Gy��T�/2�];�uwS�
ڜڵ���^����'�Anl6c5�Xbb5��휵�8��|ge���&��_E��
�v�7����T��S}f��m&��7�h�{�r������u;sV>�ߩQx2v%?u7O#,l�+iˎK5QWG;k۽9�4S�*��*���á+������[_e$e	��w�6h����,N�z폇Uȧ�,���X�=q5;���I#��s�z$�j���S�U�=�wɯ-�j����5�`'w3���)��݊F'?'iz�3��IS��������z����ڑ�N÷�S	�u�#�gW�����W��l�=��髈�U�?�_�؎�pj��=���Ɏ#-�X�;!��\�z��������`H���������fW��-��n�]c��o���!�x��7��r�K��ݝ���������
<(z��U�]Z�ؼ�q_l}��*�}���4]{�E�Ԟ����v�W���S y��c�}�1s�!�(�+�m�'��J؂I���Ө-��̭�j	�Syy]l�['������yF1�qy�J��]��Qx��zdPù��H~
gTŵ����k�Dw�5��k���z���a���-�w��g��6LQ�����H� �Q�d����� �}^��T�������C<.�#g⺮��yˣ��}^�*Y٤q�TF�Q��r�o�;�� @�#i�z׹��lD 6C�;�&��w�Lq���9�����T�vP�mu��ȹ���'������=�����vֵ�^���z��/��k�!���֪2��v��=]�m�,��}as'k��t��*L�7ݴrӗ^S�7(����J���b�U,�T
�,6�߮����C�d�;�ޅζZ��^��{Է�J�:�Vy�	\�ޫ�d��rD��ߺ�7�T�Y�+���Gk	����WWӧ��{Թt�y��Ol|jk�"zd}���sǜ����*�0T"����K��W9QqR0��|A�F���ۚ޸�L�Dln�Ĉ�����Wt��V<�|wё���븙�M�����|�����D^@N
c3�L�l=��^(���cY�/����>��{�����t���J���Wd�MO_�T&P�^���yǝ��Ϩ�0�uO�<J[��y[���dl[�F��ڷ3�]��̻˥��Nr�����-6V�ƹA��\�5���sw�sq3SO�g:��s�`p�m���W<͆kH̀�L�C��泫L�����ֻ�DJ�6r�{�D�:f�c1��O�@��b�+=m?R�I�wB9��{��W���Y�뮨ݓC�ݫ�T�X3�z7`�p%{� �;���;�ƭo��=���%�"�LeU�<r�U3�����&�sq�0�4;����u���I���멫RJ�<G_W�g>���u+d��0���	|�9�����q裺c�kvM����>7��y�]��ȯUz�^���͘��[=F���v��TLh��-�b�����ϡov��[oΝ��������^�G�ן�G��i��?d̐Ld�=�:}���+G6���#��FK�%�&z�6�H+��I���+��rA0pO^�n�n�E���<}���������������~>�oooo������$Evu��/1A�����Lbj���p�������\�Ϙ�,AYZ��N��a�@'JU�1��4)�����9�r���Z��n�K~��::�6p������L`h�j���e[�vXİ�����CaPA:�����1�V�Mf���U����vG2���D,��D�u�[߽[W���>�!�h"ݗ^�]���T�6z�lɜ��TђSr����gF������b��|Z!�=��&��Sw��g��׬��F����쮫���m͠ɻ�=iA���j=J|�-���M�s�|��z]K����b�������M6��A5�0��N�%�eER��8��{�p���� x$gR�"tP�L;��"������3e��m<L�
�a�q��U��1u)�\�2#*Ąr�w�k��m���qY����ѭ�aLfp�U�F�y��Z�!��I�:WqU����;ݣ�����J�7�����R�Q�h�82�����˴$}��ٸ�6
�Le��te��	�v�x���)��w-��+a��cE��u�n�oh@B��j�ϑw]������J�#-	q�y�Yqqψ��'7{zR���6�8�.���{}88�b�qw-���ޘ�O`W��esw�ܲ�R���D#�3%>wL��7L�oa�B��vb����s���Q�m�ۋ�� `��Lv���ˢ�v�����Kr'�k�, N��^	�n�Bd�	uy'K36(	�6�ƚ��ED����}ҕ��_hJ�����S��yk��yi�� Mշ/�5u���J|�wY]��Z52"�����o���%�������x�Z���엊=�X�D
H�r�]'�s0�S�D��F�{��ʼzM��ؓ�+��1R��;�uAV�aI��$�'"P��9K]C��Mfo;%l��D*�p��q/et�'|�nm�ph��ЁvkwwzB�g�Y��c�S����w-�v3���+	}WLb��GE� ���@@ LN4��݌��N����vL�kz���Q�2�L��t
�[�7�gHV�D۾u#g�j�o�*�j���� 2�<�������ʥس�5^��:^���f�v̫x&$ʶ��dV7wZޑ��FQ��N��)����+c�|oa�#Ř"�6��L �����O6���%c���3j�仔VHr�[a���r�U���$�!�B�s{0R�Wo`�jv*�����t��������ޢFQ�u�}��c����j�fx�:N��ccC7D,�������H^��]k`��������`{�mݪޡ��s�wk�J�0Ppꗫ�5���[��-�-'�̀��]�;̋��'ӳVm[��O�H!���X�/��ȏ.��Ƥ�մ��To�Rˠ�b�L[��s83v���VpnM��b���%�]�����DNs�\��F��F���x�*(���}�PL�U��*�*�ܷ �
H�1TM13�y�1HQDQ%U<ڮX#��MT�SEI�1ĳQLE͖�*H(��cs8'��ULE��*��4TEMUA��Q1AM%�ؚ��&� ��TNώo���9CMEMq�Mf�ëm�9c>#�!ѱ�L؝E�&��qDE5Tė3����9���)��(*�����9ƀ�P�@I5F��>$$@D%Dr6tcf��ŞZ�p�4�d�D�ڦ�֠�6��،[d��;V��W#bs��4�8�j�i-®UFث��Ta�D�C��Ō[:(���1s�&��ѱ��J&�b����h�Xֵ��Ʊ�cb�M�m1��N�TDb��\�pE4Ӧ���EQ���x=��{�����u7H������̭C6j� L�V���(�N��zu�F�1$Z�H�Ҥ����&QŶ�uU���yx�e�A�Ú�	��tp�gv����$>�c��H�i�@/���6"����,���5�h3�7N9��+˚������GGuG���p�4_A`y+��{��p��ɴ�J�e����X�v��K-����|Z&���r����׷&m�ڒ�moY�A�Z�`�ۜ}so$�=X[(le�ӵ�r���/m4�P���Ŧ.=<*Uc�N�y�����sv��������\=�mE�U�Aa��ch=�Bޭ�[�y�<���0D�� ��d�}����ƛ�re.�l"{u[ �	�r�d��22�%'�Bz
 ǩ�J����^ `�����{�?e��-�g�N ���֐�� �<E����E2��&�}��kz�\:�OGjW�A�F�X0�>��2FY��e vK�3�&N�I��Rr�@��msj&0�����	;3�U�fn�ze�)�&,�BmxLpm����uL4��&�z$�3w�S�ypk����	�3 Z�o��ũ�t�]h��������
�(֐!��˞�U��u���x>�7����m��!����޼�?$�Xƴi�9�H���c��[YGew\Hݔż�}.d
]%x����G�sD��t+ �Ө���*�P�����R�g������ޔí{b��H����1j��J>ͻ̷�S�IY����&��Nj�~nz����,�O��@�x�]g�l�0p;�ٓ���άR)���[�r��7i�(���e�1������O���V���d�U��P]GE*���]"8��ׇ�nDZS;Ow���>�}�����z����è�k-{����5�E����H�|��x_G���iS'�W3��	 ]4C�,z����ڀ��@�$��s4¸���1\�_��b��1�!��q�y��[�j��"5��F���9ރ��G2�����u�L�v�q�b����M�>	�-6�;5���Jp����C���i���(ON6ۜ�Ǟ�~`[�]���"e���
���=X��_(k�>�������oC�"���*o�,�P~�b?��V�^��#�nNؾ��Ѻ��m��%��RFq��͜eY���K�X02FI����M�v����j��WK�͝.�t��b���A>��OCV��
ej�k=����r�3:
��ថ���{�L었��Z��aE��1)�|zu�?�=�A������ex�
W�T�SPV�{�#�|�oߝr���f�ڱ�dtxu��X��X��}g�k�Ky+��S͌y�Kr�}�<��շ��a��eYἾ��>W�P�qumM[��3D���d��Z�ƞ�_��6��7�f�|:b�B�Y���z��k��\9ֺ�`5��C�8�H$whg�a����6�Cn;;ΐ�ޏtd�]	�\���|�^�<��� &I˼'=�W�TS�of�l�]J��{����;�jXO=4j��栃�;$t>Y��a���m�4�R���LS��!��m��G�P��u�ݑT�k�͑�A�/@;�0����i�'�`���q�v��N�nO�n��n�h�W��쪷�1Ly���-/#h��=~g皁A@��F�B�P�7T��x|,u��I�DMv[|�^Kة0��+�����o�IcH�C	N�"�nC��p��!����i��-�a{WkFZ��5�]N�c���,ى:��qM�,*�O2�S�4'��C��<k��}��F����nb�*lL�D	�OH���4-XQ+\u��\�⠷�[]��9��<�j�Ԉ�wJ&�O�0�ja�h�3:
y�H|.jv]�v�`��8��I�ֽ�i��c[[2�c�{�B7OA��f���6�˯s�gRdK���D)󉉍��fI�����E�6!n�+8���w��O�_�V�"��u��L� �c]~����^]� `L�/0�Tm�_��y�W&ϲ������K��Pळ%���������A�v'��ї<Jg<;��K�=RpL՗�.u/��p�;��m�:�2	yC^��1W'2㵲�uq>�xXk\k��!����]On]�S^$��\�H:Ɓ�mKǇ��	��f��n�������Ɓ!�,��O�v��3[*�xcC`3>e���%G9(��4�k����/X�ݏ��dr@_A��B9�M�n��b���go7�,�m�7Z�['�X-\�}sZ�TcR�ʖ����Z�0��Z���Q�Cz@���&݋<n�Jwv]�pl�noEG�<>/� �4�	�j�9�qN2V'j[���Md�LPxRp#g^	�hDE1�����u�K��?W�ON͉L�E��\���@L��W�i�y�nB�f+��S7���6o��⧘�!B�F�c־��y5[㼆ɒz&<O=� �򰮐j˵�U��h~�v�}f ���Γ��<S*H�aO�|ᮢ澰$f��B`��Yz�ӂ\��S��:8���o4�]�a��o����7E2���4�Q�NZ��^ p��p2�+e8����:�}ɚYxE-�09���B��P�{�t�ȴ��䠱]
��q.�[̰v��y�\�wWN�[d���.���Y�}c�zh��Sm���v��*��z�t{�U����7��u5;<�C��'�A�Z��L�����������;K�R}7�
cu}�
�\��3Z�(��i���w�������[ׄ�-` WY��]��Њ�9o.{kv�V��B�HӣB��K,(jݬ�G0Q��AyuH]
,8�t䯿�,�/�ys�G54��l�`�~��:�ꝚmW�E���*��y����;��5p����|��5~�@�&�n06�AD}�hP���EW�]����k��S:�_ϱ�zg���D{�To�§Ҡz1����P;��k�,3��`38�`>�E�Cξ�&{٨13j�c�h��{�ϖ^��l�3#���1�I^$Ey����|���z%�<�������se�|�a,������B&�kߥFk��h1ݜ`�y�$�I,i�}������8|'�� ^_�>I>����6g����h1�>�� ���{9�C�wp�o�lgIauie�/�Ԗ�v�n����O7�z�����
�})kKHABi���6*���Crfڵ%L�޿�7�ۘj��qo���Uik�0��A�6p�4����w}���/��|�dzx`�X	��P��uCޞ-�y�u��wS��TڵJYa�O�ј�-��з�xA@���F[0�`����?c[�`�j7��)
8�js'�2O�#4�ĥI�߭�����=�������G����,|�_��K�d����VR|�%QV�le'�KqU� .:םM�#�fbѯo:`7!*+ڼ�����檛��T̓�d箖-�kuFv�FX�P\�3]Ic/�{�ۚ1����� �y�7b-�@�\c�>��^̓��R�W�)ٷ�`��H"{$���Jt�<b%:�j�L��I���-���,X�������)��ߤŽ}Q��p�f�����L�{%�)�$oQ��E')���(�[\Ø��p��hb�z��*�8ׂ�];S���L�!��Bm�Lpm����TCpl�s�}/䊶G�c�}����d����Sԇs�� �f�I���l�Q�/ �p��C.}W4�c�W5������_S������"^FG6Ò�Ͼ�(�pdTK�@��vk�w��ݙ>�'�W:o4��OP��V�i�[͏܁l@ʬk��'-~��^�O�W|zD�d��]b�������E�V�i�cn��uFA�M�R�	�|s@�Bը�è�e�d���zw�v7�r�Ϫ���
Y���Bh���LKZ8b:y[B���ɱ<k�|�v�3u���i��xW�v��j�[��eйهh�/��i�P���a흨��10�́;#Y+��A��ޠLQv�ŀ�G]�s6*#7C-�]�ֱ�/e�^m�;�8q�E�4�Ԥ�$�7[��;����4�������ա���K�3�|�+�j��Z~�L+�b7�W6{�u����r���v_��twz1+;�<X�[+ou�;8�U�N4M�$��OkVer�Y�َI��b�si��N������r��*��gw.c;hV'l�5�+1<R�j٧x�]ݬ�CϞ�4;��;�7����7�z�skS{�޻|�mEv�r5�=��xU�)�4��R�J�P~�L�c��盾��^��w��Ի�u��&0�qAd ɫ�,�#ϣ6q�z�|1�<��;����'������sOy�Y�1�8�^�!3��y��i��X�'���H�3Ã�O�">�TVFz��V�M���)���v�2�b'\ezbS��b�2as�� �^�LRu~�k�*�5��vu�Q2aJ��4�l\��	܊�0�ό����,�@L$�;���� M;Й'��Nm#B����Z��9�b�������*.5FN0�nE�.�od�#	��2ڇn��醑�J�&�U�*mtٗ�Z�`����-���:�#Ɓ�l��R�w^�w8ѡƘ~	���#�Gd	d�2�T��5E
wf�3����7v�d1T�z�aU���s��-K������ߙ��8{h<y��C����́�]�0�r�p��`b�|WJ�+;I�*�.xn�r���),h#�'��ݚ�><�|mot�QK���9��q��YFX�B S"�'�������:���U/ɀ��Uj�`��8��n�z�&Z���z��ɐ���3������}\l?FZYë����V&�Ѫ�ɪ��\w�J.��0�/U'��ó�L흂Y�H�i�;̸-;V��j�l0jݛ{�i�{؛V�vYM̊^+�}�R�E��{�<`�"�S�L=�����'���{� 3xx7���(��+jC��=3z�[&�
*��ͽ�E.
%k�u��+��%锾���@�x�E��]����[�w��$8�#�Ά�4�}o&4'e�mv�a�^:�i�k]��˖q\tj�S�9[�ʹ;����U-�5w@����̙�x�`>�L(<F����fI��K77��![��qU����u;��\�w��0_��7�+�x/��  `L����������nY7��ND_c��m|��L��C��HzJ�!�F]��d^)�lg�`Kz�����W���(�y<y� '\8ۃ���^=��ƶc�o���
�W#^^z<�ƶ���t����d�FJz�խ�@���u_�]e�J�O��ҩcMmCLy0Z�0�*�Е���8��ި�|Ӿ�='b'q�'{�ϥ�¦*� S=z@�?4���	���(�K�j[�����	q2oa��qjM�
�d�M��`<_�~��*�Q?I�M�{�,�6���!�	����S�x�5-��ry�.��Π�Ʋ��%�j�U�F�c�������C�f� ���	��z�N�k;,�Q����[�N�.���{��W���Fh55��-�ŉW7@ ���PI¹�b���:�&�.��rTl�������U�Pk�>�YN�+u���Cre$�@4JB���Q�}�P�Wa�7ٌL9R^v��o��B845Ik�� ����ߝ�~��~>�V�JI�_>|����}r�刡�ʽ ���ax�I�x�T4�¼��+�w0����A�lo[֭��%�]�!�L�ΒD_k�,����X��&�e~ǒ��.r���-3�`Ӗ��\k�MVY����J��ΰR�-ŧ�D&��}�hQ;*OT�j�+_1���RX�Fv�ޥ�o�WDd�n`�8�ͯ}�m���{�#�a��`鹧т5����u`���zNл%P^�Gs�J�*$)�"ݘSlv����9]!���t@�sӇ�p���:=7�����j��˼�V�2扮�ł�����w[Ϲ
��J	{���9��f��E�|�W�W���H�/0��M �˷k��\���̞��1@ʮea<u>����&g����h���@0�:! �\;֑mUT8�h�R�_5�]���w8���9$��ǦC�$FO���lZ�X�c����(�����{��������T���H�3m���;��<M27k;I�$=D$q��i�֯ojb"%ޜ��$�n��M�nB�Y�p���c��{d���^=���#w3E_I`[ԕ�AyǗ��/�E�R.��:��y�f/Ӣ#����7�Z��4�s�rga�T��]�8�VL3w\�aZ�WֳJ�+jj��4�l�+뭩���"�f���2�q�'�&gEi�����R΀��Q�OT��<'�.M��èL��o>|��ׯ5{�{�z��[�]s��E
U	λ�x��q�?���׆���kC=X��҂��No�R=<���5%L�޵�}�a�<�U��F�=��؇)���P|ش�1���N�[W�:.��8\��	?�VQQ0��L�d�{{�[�y��C��n9yiBy���Pd���%�Fcз�ྲྀ;�
N��G5m�����Dv���B,:��Ta�j�Bp�:F%���I�Й:���>=5���$�d*��*�3�7v8e�k�]��`��ݍ!	�y���>)�W�E2��&��۞`4��Ec���m�Uy��/lbR�8���l�	K6�ϧ�R���&HޣI>I���>_�a���3�ɑ��l��ފ��Y��v��ןc��{aA#�C�ۘ�l�ry����*��rt�����KDl����3v]I$�"J�T���ϩ�f�F(j"�kH�s���e�c��
nok���?�^�~Bʋ����Q��Ï�-�c��>;�/�@lc � !�:@`��0쟋�]	S	7C��S��KO!���X�*���JNXF<��?�m�T$u�P?z�
T�����>�~�Ƿ�����������������}>�>j�y�Tu¦�s/eNH�%L�uxm��TGg#���u(�x��%�Iks��YH�����/���[xn<�L������s�m�s
�*U�hõ2�QO�Cz����{3)^	9����-	f���#��v+T�q�W>�����m��K�9��՜�
���U��c��q�H��L,G;
��^Vr���0�7�l֬[��wܞ���b)[�'�L��`g��I���;�}B<�X��A�p2�w!ֲ��a���2���_n�:x]�ߥ���G���^j��a�oz�"|l>��nA�v9�n>7��
�/.]�V��������W-}DFef�p4"��⺗����u#�)���m&�u�"��kB�;MeX:��&*�J�$01�!Ֆ�Q�ƚ˳#�}����U�8��x�iV㦍u�4N�K��ZB(67��$�D�=��l��w�B �q�dSR��\���$+p��HF�X�mbq~?&P[�c��j,~�e�M]ݱiz�*kL9���g�����X�wJ�T�����hK{&2D���ȭ>�x9�i���O;� �K@�x��B��pB  ̅�xhC���>"��m�s5��ᙑVt��|���2+�4m:�+�����V�z��u�fJޅe��H�s��&���AB���O�2��GO�(�<��<��&=��=젊�d��y#S�ܡ�-W��e��V����.��&�;r�ɴ�9F�e��4VX��� B�n:CtF����y�=�֩�/4�Ӳ�BZ}���;@��*�cC^��Ш���L2)�X�9�A�هo�{
�#��S��:����y�����a���1���ZRWm��IY�2�k4�GKY8ǡ��4�u.�C,�h������x�)s13���,ϴP�����@�oE��G �!�_\7M���)9m^�vm`���[��h���Jc$ǖ,�;���t<�[Z1HyS�	�߄�SDtN�!$1�/5��d-*���R���Ǜ�������if���R���E"����$@8� ���!��{R�ij],�n�ڸ̂Oe75La}Z�e_%y�����,�H�t��L�	�(1[ٴSb��)y�&�bX]�2-K�ڈ�e��ד(�ogb�m�6z;�!m�N�b� �-@`h���X��s;��v�wϸ��rľ��G��'.c�����ܳ��75�QT�L�&�a��*�ш��2�ɺdS����x�g�4�8����Bn��/�
7�b���CHs���o�l���ȍ�z�n�`���[D��G/��2�Chav҆Z��	z͆�ҬO
S����ƻ�#�Ґ��4G���&�2�]Q]�5�5�WHۅr+WRǛ�kL���� ����I���pT]D��J�y ���仹�u��@L2��6��>����i��mST���B@Y�U]�0���x��:�8q�6H�"f
�"��Ƃ�8[b�8q��j��UEMǘ�QUp,5����s�rH8c$HV5�E�6�G9�AM��Q1[j(��[g�.Zth�
)�b�bj�Br(���tLgi��j�<�5DG6
��9�r����`��)削b�l�k�A����c�`��b���3�j ����T�EUSQ\�MD�UT�5S�U5�1M5�p�
)*��(�媚����*(�-�Qr�F�h��!��s������I͆�*�*X��DE5P�AMEA[b&��*�nf�ss��lA�Znd5Q5E4�bf�bj��)�MQMS1L�QL�M$IT�%1���.l�C3X��Y����`�"��f�*�X��*k�����y��<w����뿞<�����d�FI*�{��Z��ЦR�C�Z�r�P�V�gd��:v;I��[��]f��/dB�g��U>���<��]�w��װ����C�{��	P���H��D�Y��>���u�Q\�Q}������W��k������E^u���� C�x�ɦ6�����c��s@�$�1,4- �{�W0�Wէ�d_j��U��X%�-MA�����>�����ìs��5����'s�E L�Eټg��W��gai���có�;c$���k|��8�k�K� ��m��p2j
urg0�\�#�Q��
sU�6���{��/�vV����˴��iϬ�x�dS�x'�lu���1�p)[���̪4��Ѱw�,�j�^���+Z��	G��2W1]�Fl�*�@�t���^�`cz��>Z�X ����CvK�@E:��0�wD�U�{T �Z�A=yd	eI�z1���Pʋ�-��L����/jQm"�f@��gDIq��צu�VL.z~�k�& ����Ja,��C��\v�~�V�ۋ�?KQ�T|>��;�Nod�fsk�&I��G���Xc*]�A���u���G���)\s��D�
�:`h4:q��i�:A�Ð�v�ۃntCO�x��aj�D�R�>!(\H��Ur����n߾�L��F��/7\ה f�%��_�����(��t��wյֹ��}�f+5e9�g�tI\{ϥ����S�*����vg>t��u&[�(_��;�u�w�Mj�䖺���}������H�T�A�i)'Ǿ�|�u����ѝrq���m��I�� �l�6S���!�!�N�� �p*��fz�'��9��!MKؕ>K\]:z�L�"��搴��=���������gs����x���q8�0]Kκ�J�+;I�P9+�Z�BO<��(��S�W{M`!W���J�K�Ü��}~v��m�$�'��՚�lĝqv8�,(] s)�u�]֝Mk��|���Wi����������-"�Ƨ�sN���yD���9����'���#���	�����u��ֻ�6�S�d5���s ;-��X�d���lķ�T�1{���^Q�x�> �Ř�t;N�0��z��Ɂ���h�Jo	16�c*Y�Ӹe+`�0 z~�(��2�ɘ��
8�� �_��c�~��W���*����Y#�_�Λ�X^&=��F�t	�b����R�}`�mβ��a�h:��4X� �O#.��,�D��y�{`3vCgZ���8-6V��T�>��o�?oa@٦��NHxm�諐�r5��t� �8�~ჄD����Y6�{��"�ϝ�K Dr����t\��%v.�]Ūe��o�O%k᪕kʓc�s4b-��������ܡ��^�40��T\S�|�̲�d��l�1n��7v��Hc?%pqh��NF-h^���~�
 V��V��T�[��V�� b���!0���=�I|Q�] CSjP:aV�D�/�]�`߅��_~��}=����X)TV���S<!64��-"G;N)�c��MT�5?)����y����ܼ�e��hka���c���u',���
P ��)\�I}�W�ppuψe�;���ч{
���o;aݪ�:[h�Is`�M�d�(�qӘ��}�9�[㼆ԝ ����*e(l�3�����N��nֈ��z�q��zGt�N���Y'\�,�$i0mz�绘OW�����/l���E@9�X�Q�&nB 
`u�e��"M�0�;"���J.���L�i�n ��-�Zg;M�������qH7:p�X0���:n�1�[��У~iC�8����Z~kJ��X�⪢݊M�1��f��L=2���^��*�M�1�5��f����u���8Ϲ�.�2��o�ͭ\��hk:�w���@�\�m/NqÊB5�:|��8u��;4ڮd�2o\l��*5��mn����e�]y(%�^��4�d`o{9Рk��U�]�@��o¾p!�?��+,�Ⱥl�q6�kzƼ���͐�s�J��.������K�[��7L{.�I�9���
疨_ؠ�ᩀ�Wίl�\�㏏C��I��״��N7g%���U)�aԍB3�oq g
3P����vN�x*tD��ѹ�2��.a�m0f�xx{�2*("D ���tu���}�[�}kϗ�gl�#
S O��S�3�נL�5x�f4Xgc&3�0Vf�s@xH,� �g+�!����w��7d3l�J.[���	P�zA�ū�b� ���4�S��5W��;۬���׈~a������/s���`�c#v�����C�$G�L�vi�'k�v�^j��&�r�O�w�r�%� BKO��-"�'��p��!��;�i�(_I`TNˋ�>��V��A���B�*u�<�M��y�A�`�K����ϖ,��v����q���Γ"���j5xf�޹LڗJhZ�`����@e�i���o�K��-�â�"���Z��d�wF�3�f/Iv�Z�^�I������,�A�W���yF-�׻~�o����  �b�S`�յ�u5�ON1xDxj{`�����Ђq@�=���er�&�~���s�:}U<%ؤ�m�+3��xa.�`d��N͕�=� �vc�C�Jt�D�Z�K"�KS�L��b�m���OWI�R��b��������	K6צ82�`��L8ޛ4�Ɉ��^���p�}�ѱ�9�l��l����Z�Di�	��lv�<�WJ���]��ANRrj?l%�r��.��W�KX���gQP'ʠ^%VW�ȣ��@�L�����cs�!ˆ�3�<�y��7���ۺ��F�㓯V��Č�6�`�0%Oa���]��M"��D
������E����Q�����X̌���R��0�����>G�e�[W�@A�9���`}�{h���:�������+qp+�~�/T�K��-?,e �XE<�Xf��|@~�v8�����v�������%�Ѯ�̉���z8��T�dε vQp&�H�P��w='�q����61��!�:C�vګ�m܃0jksow��&יq��?��ɛ�c�ɭk�e-c�o6?G���2j����B�6M�a�~%�쥱~5���"�*`��������n}��Bը�Ë>���OO�������=�Z;�(�K��(�#��'cT�2���L�a���k�}�;M�i'ә�8��<c��M�R�V#�z�]"����Yx��#A�g�Y��D��7;#Y+���w:�trxR髜��[���XK���d��kIP]ă�,�4S���%�q���D·W����s��9�l$��z����V���>^��4W%ڂSl�W�v�o�i�y���%��#�F0�f�w�A��<;�u�<�m�Z�^&�Ө�ZՆ
*� ɨ%r�P�*�{ӭ��l��g�s�k1xdW�P�cۻ��!�y�Ĳ�zŬ�3k��s 1�8g@w$%Y�љz���va�I����r2{�&jـi�p��R��{"�r�5�/sKNd�}~�hfJ��F�5C�r5�nv�[�.d: �Cс�m���<|�x�z��~ �� bi`<<=������Ⱦԯb��/��1�E@�NE[W�A	�� ��@�I�} �c�v'���mY*�FE�wQ��S��u�+�p���p�����L��C� ��&):��ХE"��|�;7����/O>�Z���-�^��1�$Ao'0�w0���;p����<�	�z�����&�k3�w�[�lq����u6%QN.�H�hUӍ�DcL:A���S�v��fj�L��x�'A~�~�P�b�I�y<�[t�O^Ҝ�\��|������"����-��֑e�1	�z��3��%=_�L�"�<�4�/#h��=yߙ����q�h�rm���{ޝ�^@áA�=K�9��hQ�v�
�����nRy����v����ٸ@�{�[�2r�.���[d�.���1n�)a!���OEs� �в^8�*y��y���azX����@�W�Y6��yL榧���C�)[��t��m���M뎿'�\��Y�պ�1-p��CZ�q��{������{�=���3:���춽��+���w���g� oƑc�c��_1S/�z�ud޳ᙎ�b��1Qp�÷nf�(�z����R���N�e˼�#�u�K���s%Wt�5�M��(��6��3]��ps}l�mۮD���ڣx�J�Sܠ���QH DfR�)<��y��xx��<�]��h�u5�eC��j[��@���g2dK�p03X4��틑�a�55i����!^k�L�O�zY�ܒ���v�n� ��i��ƺ���yw�	S͉��~ה����*L�^�%���u�y�L(A��K=�L�=����	I@A���i��n�âm�<�N�O�;����n�3.�*o��4�c��S�0�7V�Y����w�Ar��ЖyY�� �teC<�[���s�݆��4彲ީ�u`�x#XXd�_��h���1��*�M�~�R��A��0��'�(�h��ʮ�{�#w��9�
�Z=��V
��/��k��#K�`b�d�NԷ7n���[�ٹ���u>mM�ڤ&4�ׅ'�(�=���o4���1m 'C�L��;�	=�3��zp��^�,��%_��{��u���M^�7�c26w^��վ;�alM�n�~mh��;�?^(����О|q����k�	�\�^%�:\�L�#I�Px`��~���C9���_����͓�=K��#��J��0�;"���E�7E2���7g�x��̆��p�QUh]�+TG���Z�KEAm5u}Ǉ+CdD��$����
���jZR���^�8&`T}���P���0�]l7�m��l�V�-�qLSmt��5���b�z��ܛGz.*��@d����e7y�t��½=�MӢ��\�7u��n����
UB��&T �!PbDM�����JƩYO-�mx������D�LdT)_�҇@⮗��i���g�'j��Ni��Թ���������=���kLp�n��.��0,N��n7o�?4��m�k5��S�ܕ2�(��l+����4���B5�O�tz:��ؖ�F�d�ر
f�����l~�,[��v�A/r��9��fk�^�a�5��C�w��l��(B��~�M�L���]�6�̪Lm<u>���׉��w%��1a�y�(�E�<9��뜚�(f�t�@C��3D<������d3od"��=$9!���1^�tE�e0�5��v��.���r>��w�h}a!�xQi�ӱ��g���vq��
����{�-7t>2Ot쐝��YT����N��7��/l����g�#�ZB�	��I�z/^�wP摻����c����u���Թ���䮆�)��+�~9��!CBQ��~����]-Zϒ��T^���q�ض�7�y|i���ml�ʽjq�jH��f�'��V��"���h�������XΪ�Vw��=Ͳ<4X�kxέ,f������C@I�a?����Y�]Z� ��{%dyS�N�/
����;~\���[S�������2��;��gv������>�Nǵ�6�a�.�Wkj�|/E��|�A���*Y�fn��ʘ�Jӯ}������l
,J��")2��
�"1(J�]�ru[��3l�F���9]�tBk�(2jXf��.�aG��u����o��y�YD�D[]e_��ᐄ�" j�`�{Q���N(�=�f�\�I��Gc�i�Ewb�d�^�-�����y	�X1)ٲ�#ݍ ��y۞������B�)�Cu�#�27.��@nd#2u�>Eê�󍐥��)f�7Od�#�L8��4��MYn�9����W*�%�<�����-wN��y�|�-�y#��"m	����Qv�ﭝ �3qfm��K���n�P�_Xˠ�Z~X%�@�g�-qy��i��^�äGS�X(-"�qZsz�TbjηkDQ������e}�����E�jF������>;�/ힽ�ga�tM�<l^[FޮʓL�^�js s	�]�,tɬk�zRr��FM���`5R͚��ͱm�Yeձ{rug^m�p��=0�X}O"���.���dRAD�E�Yk�'���j+��Zfĉ[�Ll�9�F���T!�g���xBD>���t�C��~���	�zi�y��=ԴTM3�?���Ʉ��)z�I��1ҷ����e�cJ¥��Qy������Q7]=M�0i%B����n��TO��_�G�������]�8�\<������;ʵ>�{��[9�9pѮ�rT�b΍���޷����7���{��^:��� � � �h�Q&U�ZJ���(@~y�x�y��>�x:�}�^K~s��-E�;��x���0(-"e�c����wHn~�Z����&��n�X��wP�9Mk�2�ZG.��z/��{dK�CF��i0���3�����~���7JbkW%7�d����{���f��K�%6�5F]���֞��6}��)�=���*�^T��*���]�aKW���&�Ӌv+Z�u� ���*�BFq���8ʲ�����Ò�m�x�N��r��5C�:@���|Ǧ3r�9mZ����0�	�,�,��k<5�q���M��e问����͡8��\d<s���u�P���A�e�`����v�6��4�3�}��jy��ޡܥQaLz��:����g�[��Y��v��.�&�Ss#7P�6NZ�w��m���T�n�Q���W�����8�Aȶ�X�8k��X���t���7
�e�u4g0f�����C�_;Po�/�D�"��<�OEq�lGM�f�xa��!''*�.��TT�c�K�یV!�`.�@�=�jZeIOVL�"��搴���[�|�O��G�������{��������������������}>�x�׎}�&Ll�J�#�eMZ���v\}}�4y�ӵ\���E�UL���Yy�yI,J�t��Ej�$�b�+_N�g�o@zOs}������֪	9ӷtbǥt��V�Z���K/0kM1Cr�[CmIϞ��F1�iԠ��[X���9��1M@w����k�1}p��6�.����-��v��'L���B�D��9�qB�4$�G>,�n[]�q�-Cg�u�2�q⚴��֐�ֆ�_�Q}���i�Ǹ���{C�� pi<��WdU�x+;��U+��9e�Y��.�*Y�oxއ�{FH��;�����HH%;k��\أ��C�m�3[h�G���d���:�`���
�ث�o%��}��в)7�`L�G��V1MC���j(J�ޜy����ƾa��w�!�����yV*
z�y��d��f5�.-Ɂ>���dz�Z��wj"�	il�91���s�b�������Q��$��x��,;\v:E���ҳ�v��� mVP��e\k�u���������ê�r���/Vu�Sj^S���V��w:�]���S�VޙO�.�[�)@zʂp^^S�kl���C[2��aj�<&.@Y�89 �R�H��^���a�[�m͐m��j� �_o�Ƶ�G����;xU��q��Tv+Ɠ6����9�1�n³�0{���1���ɫ�rں�Gt����eP�A�jT�5��[��i�F�9�ev\�~�y;��-��݂6cw�t�"#�γn���H���� e}�����3+c�2�J&�b�zpnt�:�e�2�+u`���l����&��=���3��%o	6�!]�ĒD6E+6��Af��i0�_,���u�;Q�z�Ʊ['��ʴ�u�J�ү�54�0����i��2N�������]�.J�t:+��b�+U^Q'Sҹ�u�,�/ٖ��7�;u�xѷ�]��A3wCWx��"�]���U��b�帚u���1���#�1��+(}�7X�ҷ\L=�UȹV-zgY�E뗥���]��<��r��[Vrћ6��iolU�k�έ	|\���W��AUݩܗf�N���C�����ޠ�Ә�*�F)�<r���C�T6�x%I�t��e�vɰ�3d��}Qu��;�$/�꾣畊Ώ������7A ��2����Q^��fz����p�&oJ˃�N��c�,V�nM}͛x+�|����s3m �&���
f�bޫ(v�Y��������-�r�r�e=-��ha*j�q'�muڍ�P��4��Sgpr$'Y�� b�	ۃ{g˷ϵ�)dq�ڀ��jt��mJ�Jhm����m�f�.@t�=\�bF�S���؎3�פ]w�A}þ��N,ź�y��Q4OF�ɷ5G�i
�t8o��UUT�ULV�PPUE�h��d��"*��&������*R���
H!"�&�l1�����2�4��EU-Qإ)	����� ��((���IAQ�b��|�fJ�i��&"&�mT�AE$F�)TґD�D�EDU5m�&��J(�9h����d��������I�fX��(h(*�
b�&��)����*���,�T�QPPL�1��P�SJRU%DITEE,DEQQUm��j��������`�)������)�(��������Z
X��� �!���( �������PDD�5T�PPQUMCJQ�MSAD@�4�44��|�U��m�#��l5^dp��˲e�s�ܖ���Q�F��T"�ܜԻ�\����	�-qKU��V^��{�<�Ͼ����eT(�
)A�d�T�R�E�	�(�|��矞:��`p������>\��_�L�=��J%s�Y�I缔�4��0�o�qOUK���v32����"@�T�"��(�q4������V��f�bN��⨰�Z��R}'y�ٝD �%�VN�Z,9���-{p���p�'�8g�c��-�Be@OH���"�(��:6m�'6�mt��Η܅T��A/m~U�Nؘ��s�w����39����e��dT�5�A�s�s+���V���PI�'��FR�ǜY}�3�끀��M~n�\��g$1��0_B�f�����R���t3w�E�x���D�1ׯJJ 5ܵ���`[:yחy�,[�����aÓ'҅!�/�D<���ۜn9�L�3"�x�zO��zJ�öl��k�he�'y�YFn����N��R*��N$Fd��騼{kݍl� ���/���T1��ХsU@��ѧk�ϙyEۦ�z�\��a�
��sE�
��{{�>�)��ܮB�V���e�!��Y�Q��ظ6!��V�*��zޜa71P�)��}�`�È�lQ��=A2"/)űy�����y�а8sq���jU�N��Ddʛ4�88��܂��N�׋��u�!J�ݩpc�9��
J4&�N�P�M��ZŔ��g.B�I�T��׍o	)�c�A@�����Й]��4���8��Z������u$~x|��� )H��J4#J�0*���B({��}����׮{�<x:��c~(N�X�!2��Хp�I��if�7
�/���i��/���*fp*��p��Y>!��5������x���RX&�EP������xO���}�;#e߽0�,t7��!��݇��'�u��@���3��s�2H�a�>�����WE�V����[�/l�%�c $t3d�!0\�.Cwc@��1�y�E�F�C�YW��=`���ވ�������T(k]O�A�6�8z�:ٱ��	��n��hQ����S����˼Y�5�Sz�dq�������ҡ��'�h��GX��*�Դr��mz���յc�V]�0��[�ܝ㬎�5F����u'��w=,��%���܀� B5�O�tz:��K���!���Rm��,^9hv��Z�X2�XR=+�ʂ^����\*�� 9��G�*W]�7�6�^���^�j���z��%ЇktΝ����c`ʤ���S��N�fy��K1/A��ձ��l=M����mj�`<X��})�k�~���#�Q~�Ǥ�$87��x����AM5�Z��fZnHmu�BT�%dSW�ö����2n-z��bRf����6������]QR䌒j�X�n�Y�bC�+I�v�&(�3L�~�	�S"���.�:���I��MEN�B�Ք��K�6����"_Xń��� C���+
����F����ߍ�h��ϴW�AJ �@�V��
�iZQ� "�4GQ0�͋f�
�����tK�pr�Caqb%M��ؽt��7fM�v>=��1��3h§vx,�`'e�}��lEC�Ȗt�5!�Y��'��{9�C�ݢ���'3�goKu�hZ�0�*�!\�����O��o#^Y��#�ZB
Lde9�q�%�tP�47L��v�^������l�Z�`�@H�O���3�J��2�
6�"����μ�=��:=(T�c���W���Jl�L�ɨ,3I�Q�a^=�@[ռ�9O������W"�wAo@R+��"zXH$=ˤ!B3k��� ���?$f�\�I������-9X���n��z�:��UfT�d��'�Jk�ϰ:"NI���>�N�	�^��(9^����Ų�
l'gZ���Yȸs��X3C5����;T�]���0�.�3�g�TA���wzp�F�҈��ct�T���㚼LYz|�>�a�̃��"m	���i�2�M�ʩmk��ۦ�ױ)��x�&�z�}8��R	u��wf�H=�=�6�F��_�y��#�<�U��9%LI	�#Pr��of�'xC6�V�]�A&:"��ot
��r%�.�sI.��5 8/7>ֱ�@<�@b��"L��8���û�Ǌ��M�t&�r�R<c(ŵy�z�%���lm48jW�򙄣]��|��������1 RP ���% ��R�Ǿ�f�q\��>�6���Kwݦ����/4-H��)�
���>;����61��e���vS��tm]bk~�F/0{瘯C�J�=B�ՀjE10fڳ�����o6Ϡ�K6!���Ә�ʄ��~ݸ���a�;��C~�d�ٵ�~����"�(�Ë>���OO�Ǣ�E�뢀�(�x^5���}T>ߟV�.�U��떾�F�=ki��G�����
�,����TľV���LI�n�J+����-D��#��h�gh��&9ف���M��r��I�s�J�{3m��r]{��C��v�ŷ�q'DYz�x7��+�AV�\>��ׯȸ����9Jw( ����~��GC���v��7]���^Jm�nF���?sͼ���fn1S�ݦ�j��
\"�5��k����؜kN�q��BYJ�A�#8�C6q��i��Zn�'���"Y�׋Ӿ�����E�C�0�3r�	ȫmNB�͸�1XuM�E��a����f�ь����\d9�23��`�.6�ėi���Os��Ә����ǫn��x�����`��l��I�,Sc����X��j��6���-��\V�ɡQ�*��r���W��^��h�Ԡ2n
���7|�.��=�,��\���Q��2��	���@��e^#�Բ�Y�eeno\��C��9w�^�z��ǟ=�Ǐ?4u׿��j܀R̊% �#J� �����u9T������У~�I�2�lQp��3Ĉ-�Pe���	N�#r]�SN�B�F&y
S����Zw���s�:��)��4-\�)ſE��ȶ�@t�z$��t����1�r:�7.��#��.� �p�4���&X^b�sȤ�
�@ߣ�x���OqW~W�D�/Ӌ���G����;H��&	�ݐ%�v���RSՂf�X�4��e��u�O;ŘQ��0�K*7"YԼ�A��C������A�7�W��
6�aTJ疳P�����ML���qW,���\uA���̽��>p��X:n������W:�WB����/��������;r�R���Fw,n���rQC��;ZhP?~���
:8:U��@���4-f������ D�sŬ�ع�˥�C�J�I�zb�9���֯s�w���4x��g���͖�5)<c��iwx��T�mk�R�HO�Z�8ô�R����_�|�s�&���~�lgc�����9��gx/kƥ�S��Y�R����R���I�v��-����>=�~o�;nQ~�=B�x�{կ��K�q곣�������i�՛Q���1v��hU
V���:"4I���pw5F��Ȯ��aI�+��/l��V��t�ۥ��y�G�
��<ϑ�Yʞ�q��|"��<y��z�>n�G�u�|�s� �AbP�H�����w������s����o����y����F2<;��@̋!�= ��8A���j�|�/+Kw�������{AKe<S�v8fC@���`��I��Qx����֟fA!��/�ꖦ�At?0y[��^�M���w�|�|?r�g�P3*�*P�����O�7xO�4 Z�EGp��KA�ؕ�;�:ȭu�c@Z����6-�C�9#b�z%�&Ƒ�`�È�i)��3^cΓ�,��8z7,l�5Rɨ9BSe�d&T-�ģ�.���k�U�_���r;���O[�J"�b!�	��O�W��q�g��~BS/�ZRX&�EP�ػ|��	�H4��&*�Ԝ�6��	w^!�{ؠ��` _�����=�):��,����2�$i0�T.�u�3!�Ǎ�����uje�uDc�ϭB�lwL>K��=�"UvQ��Ȣ�3�V�k{��B�@ܞ���T��^GnуNY�6����B��GM�&n��B���*9;�0C�*�]�.��w��+�@�Z~d��[Y�\<vǃ찏t0t��#�kuzvh��8�);:#�e����lz���g��W�6I��[�T_5������Er���9�$H�+���3�e�{��V`��b$A�����xX<�{��Pǌ;5�@�6��goº;"��
���F�U��bU3e*/��8u��;ٝX����X9�����|�s���?g�4�BR�#BP�1+@P�=_>�|��������opM����ñmg�1W/@Z��S`+���@�^�<� !ý��ڨ�om}���ŏpo�y��k��Ml�J�aH��{T��/�W���%�kݾ�a�1�k��ةoWY0�Pu�/D;'-1������Wz�`�T��~���>�z&g���R��k��ʎ�C�Tv(Tb1��B
y�<��{��:~�n�f��_�1�I^�D�Θ�#RC��d�ݯ��߾����+r��2Wߩ���}��\O�T�{���K �&�7�\��;�����&a��u�ڴ��U��B����O�؊��xg�!������<sս���(�uب�܄���4P�%����B���0��"���xiז{�}.�:g���Rz��Y�-d����[nUT�y��6�4�L�`�ʭN7�jH�w�,oN���V��Ȭ�C��c%�S4gN��q�m�����׮��+�Ռ
�ة��Jn��A�R�4��(ΰ�ј����Kdz�xͭ���2��pP2F��	� ��s0���LK$���d�q��(�\���7ïI(��u�7ݙ������{�z����JfN}�l�k7�'%��z'��t�9�	9�<�ԗ_QʝZ(>���	9Ȭ�Ӭ����mghǇ^7�0wv���GI���d/!�(��i[^�7dÙ�{B1�%R�xn���x�x� ��B�b)��E��#ј���{gOMn� ��Q%ٲ0]m ��y��%:O-{�i�܈����7�s�H�5�Q����'d�k�>�����ki���a�2��v
Z�9��h�	�cw.����t��d�&�imp9����#ϳ�l  �y�t�J�gT�w�]��!s+�T�ޒԝ����rt�{�Z~XH%��ˢX������)��:���GwgfO�C(z���q|���uv�T�\�I慩���w��p��^L�(k�ϔ���t���[�m���$*��]ً��=B�՚�Lhɬk�����2[��j���U�E�lG�{�%0�Ξ�xH'���U$�`��  �^a��Х�uCs�i�K��L:�x�Z�B��n۷iStE������������ uv��C��� 1`И�����t�C��~��kh0ܥP�"%�V���[vGZ�pP������sP/����3�Έ�v�
H���`L����ׅ�4�1Tq�/0�=����z�'��hC��5%ڸ˱i�q>�Sǂ���钿Q�7�_k���I��ђ}��8Y�'[����:�W:����kj��]�f`�}��(ɀH�W��x�_5q%�Ե���s+��vN.�2���s`amN�u{�*���'k��e�c�v&C6	A�.����Gs�@�ist��Yi�ؼn�>�����R��%�B���s��m�{�}���(�]�%6�5�˴�o�i�m��:�-��^iNf$A�n�;���20G0�����5��y��a����2j�W(5��?�>��P�����U�l^����W]b�������P����l��V��PB}k ��5�:�ܶvY����� O����ϝ��W˰��Q��qwb$���Ӫu�lk�N���~`h��|�6���͜t4�QI�#"Q�0���8�/P�.1��-��,ֽu0��B��CTV�Eo4aٍ�F[u;P[��59��=�)�FE(S��>Ű]�l.�o@>趣e����'3��c�w�f?�~R�({�tduU���j�,�x	���"�׊�@�t�z�[��}����3=E���U��l��b1�L��	��v�wc�=�%=X&m�u�`s-/h�̩Ɏ�����Tj];�>��mC��0�7sץ�?t�w<Z�
����7)<�m�ɧ�Eмܽ랲[W�چ�xwf��|yp���-�耛�О��Vj�Y/U�ǫ��1��:y����j�{"�I릳t�98��ݴ�oJ�]�ل1�����A:�[�W�f�!��	�B�z:ڂ��]cl���Ϭ�$�E�Z�v�%"���f�ƅ2��;w-����]�zP�/5����VV�����v�T�r�H������3x�o33uW:�.�'��L	��������(�0�UZhP>���4����Ƅ�m;xx*�<ٙ����읾v�s���~��`�%�Ts	;bu���Dt�����܎yi�ID�d�c����h��!��T�j���sP:�i�k^�v�&a����\�s�ȓ�o�� 4VF��Y¦r��c��uyR̋��f�;�XW��E�ęf:��;a�Į�ԋ��|�Ow��xu!,��]�@�9��!�>0�s��t�̋!��C�	@A�n%d�x�n��*n�U�.���lCz�F�������hA�2�aq1�)=�j/�u�fB!�4�!�r�x�V��4���tU��@�^in��L\:�tS<`��,:N$E��{��j���Eٍꋥ���"�(�r+��D����ءT-]
V�p��8�}su�Є&��b`�+Z7L�T[L�E��*���vB�y����nf�!5���A2�2%?	]�,�$!�e��|��;�M��|y?B?Kp��k�O��0	��{�VG!I��x��Ғ�5{Њ�vl�:?y{���}9��==�=>^����Ƿ��=�>�I��ʈ꽳<������7#9(�[����j���a�ó	9��-\�cm��K�ߢCB�t���6a����A"G��V���j*�J��s5ڗ`�g�}�f��Q�)�p�w}�SA��r�'e��Vi���������*(332$����h��JԺX�nmf������+{JԸi65:�d�շ�vh���o��ogZ+�ܵ��/K��Ɩ\�C:��}����C��\�hdq��Y..f�J^��`ԅX�rG��C�
��f҈)JGV�P4�5It���-�έKD��7N�n�U�>�W�p��LӔ{�| �PL:wI�ѹM�BY�yK��I�U�])�ON;��I�{�]:��^I� SB%{R��M�_�㐷ԗHs2�دvte��[�����oZ�+K�4�˫imvSR��4�σ�9�e� ]ͤ�i�C�m�D��Y��6;:D��75�<lEn�
�3��׀l���5��cVrb`��[����[
�C5ᥴ��Bl��	r���cg��8�n�-V+�"Goq/��ٗ],f��3����έJ���Q[y|��gF�j�fE&��h���*#�e,��])�äVg��Kk�v�\iJL��]j�����s�����WN��B��M0X,Y�v�Fp5�kt�溓kR�g\b�a��|��/	5t��S����0�1"д�ɰf��z�$~�]��պ̓>Cew*��hӐ�j�^�t h�UgQ:I���м.�P&�����y���B�N�+e�M�t�[5ͭ�1�r���� ������Vu<�<� ��t���AO�[��S��Nwg|^b�ݴ���Z��q����.��q�U�r�@�\k�/���~=�)#���+��ͣoW�h-Gi�a˖��V*�;u�G�����8պ�e���l�Ӥ�	r�v2��칩*�wkZ��L�$�2��+���[M*Yd�wȾ�s��]��sZ�\d��Z��)�Up@�w�����Iɫ(�Ǻ�-s&K�}�y�]�m;���&^�k�:S�N�-���̃Og6�m�#�2���2+�Cޝ�s�~�X�G-�5��i<g�7jY�d�ld�3Qx>a��ǰ�@l���K�Ѐz�v0z��|��<va*�3���'rv��0�5�Aau����ىN���{V��]�,�.�e �Z��4�u ���B�[/��!-0��ڕc�y[����Y��ʧQk�9�a�l:�])صq.��Ł�d�ۧ�_g�ː-S�G�l4pZM�=R�u�Ag=ѝ��ڙ�=z�{`6pΤ���v��}�6V�D8�ѝ�ܘw���h*U�5Br�I��	�f��y�-���к�7���o����s6��q�]U�ԁ>��c�|�4XLɻj� ,���k6���Uf3�6��u��O�aJ˓nl�I0��X,\+���)����mPm�͚HBY6��ܭo\9xG܅QM%RDR��QI��R��`pCI@U#K�QAQR��D�BU1R5E1RQA4D�i�TQ0�BUEAMċHDR5ATRRTI@UAT��4�R��R�SF�IH�D4�DL�BL��DQ5D��L� R���A�t1��Dbh�
���Jj���ih(
���)�������������J��ibiJ(M.����B�����!����������bV*Z͚��P��je
��D--1TDAQ�M��!QBR6ƒ��ρ������.{����:�������"�Pu����q�n��ۺ�1���S��V�\�v_��*[g����j%�'٠
\i"�ȼy����n��'
ʊ<<K�c�߃� �^ ���ƀGa�gt�N���Y'X<TyӥoHdv��X5=[�绘OZ��$fɈ,=.Ct���J�p�0��%�	�ƠC쳩W���ֳ���E2:f�z�5��7<8{h����:n�	��a�F����{��g���t>y�B4��,�T#��PXחJ�栜K�k������6�����\��u�ǩ��V�Y�kêm�jV�2L��aM{O��HWC��,��oϞ��pG��a�[tLmN�~��9�[S�×�����o�U&�W�*��#ҹ���ڸ�7P͹�l�,`3�p�o&��ͪ��HL����;'M1����=�f�Z�J|���[��c�����ڜ&��/����P���ݮ���D"�!���:~��!�{!�c�]��ʉ�f�� �d����᳁k�E{�=76��}�.����𸘕6^�;��h1�]���=ʯ;���:�ise� Z���=.���[�]�����B-A��l���}��zd�F��lS�s�
�=K���+��N����{tn���Im��X`k�{ڱM:�"�ǩT��ݍb̖�Xn�A\h�f��(�=�+�
��<�#fe�p���cB�8�ƥ[��6���{�'z�h��|��dl�Ȏ|	�wc2�M���<xr�uȉ_ʯ���a��ՃN�c%�^���q��>��L�W�X��B�).���m?4S�^����?v��S�8e'�Y�� �_����ס�3m�)fÑA����	�����8�i�s�5�8}��Jz�xa�/��<�\zz���	_�b�=�Jl�=�5��4���Xi��2�&���l��4�ޭ�=|w�
!��D�����[ ��b�i�� ���_��hf12e����R^��sr���k���ơ�l����� ��Q%ٲS=�� ���ϊ-�5U��òGF^�i���~^]"�W�4��os��f��u�=��ki���hLpe������Y�1�wC�Ƿ
Ntp�Uԓ�yNR�t�4���5]�����ٻ�ӣPJ�kb�/�H��,*c����MI��i9	�^�ŧ����B�����i���䥥�ue��d�?kL-S����'�K��sM�ګ���/޵#YC�	Gs�O�㰝f��53�5�L=޾�o�;*��1L� �d0u�"�~5=B���R)�5�vzRr،y�8�_'���SF��j�ܫ���F9!��%j�{QVo��,r�w�S�� �{l���Wu�A��}��c#pD��l��,\�5�H{�z�|�n���q���q]Ywym�]��ٓn��*���:ܛ�Q�������Z�Zr��yP���7�f]g=��emu�}�R͗�(H�
�G�/�{Ţ4�����hZ��u�;1�����F��s�j�^*�k�ت���Xt�v������D&-�����W�a��t�-��Z�vV����ʗ8V��0�Ţ��l%�������D���<����be�X��Qnk���T�d{�79��I�.��]�H`��:"���o�ȗuG��������uc����y	e���DL~�ON6ۜ�t�e�f�=$�PJm�nF�[�Z}~X�K�%��{x����[� .E;�d!��[�5s����ъ(0���Pl;��b����2/xi��L��ج�l��sӼ
H�	<�1�L܂lNE[jr�(�}-T�ⓩ���>�~���l@����rϜ��~5�^5���!V��L��F6�Y��1Saغ�tA���t޵�$�*�
e��:���\c=
`z�f�L��[e�6�+��"hb�P�p�Y����Y'�b%9HȤ@�E8��cŴ��N7��=��J�s �������!�����Z��y�FI�`'L*i��s���.�B9o�v��6�Wh�Lˌ��Y|��+c�iG�';�Y��nP]���5n��J��'V�Sr�SMڝ�+�7�m��0��{J�A����PW;��jT�A���cl7��z�q0�2��v�ӹ�#��&E�&)y���N<������b0�* �l�Gza�<�0<�#D:�A�`"�<���TuCOeIOVL�"�ն���R&��ߢҞ���n&��5�Aܳ��p��0Z��0g%̼���B���¨�yd��w��_w-c5�'w�_<�
�ʂ;P�Sû4�|yp��!o3f�p���WM������c��YÁ����g3dw.���I�Z��R�u�j����n=��gᣁ�����_m��jq����b��b��SR�B�xX�'�\�T�֪9���֮{�=���34�	��!�����7N5P��J�n��Ú�u*��ֿv��j[���#Kߋ�g˘{87 2�^IB�4p�)�`<`���͹��f)Վ�f��ܢ1%��~%�����	���߳�_N9�T�^@��l�����:#�B|aq�8��K0�Ȳ�@�C˱ڈ5Q����el6p;��It�H�l��n}.��bgZq"3%'�ME��^�kP�8�Z
�?�(R%�Tk?eEiWp����#ߣ�>�S�~�4�˕�n���
�̞�%=R�wc�Ǘ%�lfv�a��ي�0��oj[g��i3�n-�|�9{����b�Dib��LK#�i'I;e��j��U�Dr[�]�Ԛ^�oa#F��	$O��R�ݸ�3�K���p<6#���C�xϛn6�5��tS<XXd�\]���}�j��p�Z�M-�l�=mf:a��3�Ak�z2�*U"V�*;ޏ���.b���=�M�T�-������[e��V�C��S�N�7u�Է5�%6Y2*
O��Ӻ��V��6;�w�6TGh�������=��{�W���ĳ�u�I`��B���/8�]�O�����P��Jc�ޢ��WW���l��Խ���<<�d!�0��S�\GV<b�Ԗ�0���� �k�G�f�t�s����i�vQ��������6N��uv*��ڪS+�-�:a�~��>w�>�@�h(f��GM�0u���/�6�Ħ�x;��T�*P�⮗��i��r��t�~j	Ļǻ`>��@`鵪���:��6ϕVkxn�)����h@SR��־�`X��|J�/i��IWC��,��%���܆�8�'9�xЅL�&��n��*a���p�9�٦�}TZ�%�p�B�Gb	����9��3lyǥ���~��#�v��Xƶ+N���Ȣ�YO×��J�Cѓ�q�P�VG�S�:� ����=��9vsЀ5��ϡ���ބ��9)�g�V[�ef�D�N)���*8��[wsic��-<֋���t���_YwƄ���UA�o8��#�o�z�0g6�By�mtώ����l�ʤ���S��q�N�*|�M�w�v�{Ӱvdu�,�ܖdy���M�zb\3H�`<�ȇ�|/~��O۰��>�y����������Ϝ}6� nW����l[�;��tK�XP��\O�J�/����$�I��
�S}�m�[�(T�;O$9!��Ӵ���}fOP�^Ȗx�ZZP�-�h��������1kat&���p�i��*f��SJ�|�/R]��l�r�Oz�Ϲ�BfƜ]Py��^Tw�52�q�1���uR=)�rfڵ%L�b�� ���	�r9A�ٳ���K�ވF/�duk���5"���[@y��q��S��ج�
�JmJ82c�i?vc�;��V�-�X�uѦ�Ƕ�x/���(��؈��[ �����Ђqӽ�z7�����=wk������n�@�4��)Rk�����l���qxIvl�	��v4(
�g����(	��[���/�z�Q)�|Q�Z�^kg��&���j|��\�����m8�^nq��t�w��|�[ }4��}V,�E)�40i4��Y�1ɢ��fM��re,Ŗ�(�|�ט��He�%v��s��[ʴ�\��5���¹l�D$���x�GR��1�V���ݝ��m[���p�/Dwu�<яk���7�CF��7�Ub#{��ӛ���0�zL���I���V�0��La0���g��F0�
�Aʻ�W6���/��}�y �#�(	�w �KuL4�����Z~XH%�yH��3L7_F�l��2UA�[�gF�0��<����`���_��sM�ګ����BԍeIGs��]�	ٙ�R�˜G-�C���wh��<F�S�����О�\����sfMk]����pw�6�]�*ȅ��k�7ܳ�P1��큗���
��Q��#O�=�n}��B�&6ʪz���ޛ��;�0(s�e�a.�WY���a�#�C�H���h���x"�^��}} �4�ej�D����'����Q�I����0�8����o���-@��#��?3���V��V��3[���E�dLR|�N1g`�2W��3���4"�Mj��.ŧ�`��:"���x*� 5�m�L6�n�tc����!�s�\L��m�{�}2�3E�K�RN+������L��/�Q�n'��FJ��oP�Di�{\}���e��Ƚ���Wn�6℃���A�w�zck��Rk7d��!-3 �6C�{
}a��cpV��g�n=�Z��p���t�Z��/s��Y n��ղ�>���XUй�q ���%�R���� �ಕ#��� ��f��@`�����9�)c��ܘ�`X�\�a7J���}��y&�	�d>r�C��V�3�l�,qL������`���1��܂nr*��]�Q���R��y�l�l傟[�΂�ʒ5��c��^��8fA8�ř��i�1���qc\+�͸z��X��B��A� ���M�[FD�RXK%�8�����D��v郶��ۏ+��ǄͰ�]��K�/��5 �	�r�	�I���&JqO�l;�-�3	0��V���]�4�o FF3�Aòr��x>�DO����Q�!1V<�Z{�P2��-�
Z�[�m	�1YYd�]Z�t�m��7�pA���'�^d����f{*$��&m�tU�K&a��&�%��暙��Yq���;�?<��������z���A���4ҘN�nff��9�����M<�J�s�6�Ƒچ�٣r\>6�`�D@M��y�Vv�˳+�ܕSr󓙍}��;����q�!�Qak��I�7�
��teWh�C�4w�Gc�ǿLF7e���R�ۈY�4�=#�j�j�J�a?J粠����9���֯s�w��/�=)�7@!c�1�������z,U���i\e���G���s��p}[c�}~E&�JA�x޻�m��4�u�z�*=�F�����g<�R�J�q�Wg��K3��W�Өc�y؃�Ё���˃O{��6��.A�k�ڤ�.�N�u�8��8P�͓�`LI�m�f� ��IF���,�����uH����˨�v9�%�����Vz�;��$,��=^�Y��y&�_y�ñ�c�wR��UH�}��, ��~Ɇb�n�6��E�/�A2��<��_�������G]��T���Adh�/0�P����a�e�&��#���ű\Kv�Zy(AF]���e���\3o�ƪB0�}�I��5��"�
�_���d�����إ�ބC�U� �r�F��q�髦.s�=�k��Jp�x[Xވz9|�6^zsUPZ��T���c�t�WB���p�7�M�T9���<mj�;W��gV&��p��{=�cZc��'i��ن�����`�	� �Ф��Gh]��בMI��4.�,�����Je�}gm	�8���^!�v)��%1�1)ե$��g�Rm�2����$�Ɖ�B��V~��:�hg���ں-E�����;�k��	:<9�o�P���+��r��9-�ƛ9�'��1�Q�(i|k(ȯ�ѣ*�� �;�¿�:�!��4�Q��A��Pɹ��T,���Q�m��3�4�NSܱDƴ���L�P�օnngpܽ��5Ŭc,d*�\}�Op����,bD&ȯ#*�V2J�ge7�c���[����޷w\�J�RЙ��v��
A�Y��rkҹ-�#��N�y��W'��E�J�X������NZ��mvM!����wZ��}UC��l"��r�J��P��t�Ǥ����t(ys�´�(?���e0��܏���3<�d��-������56���h]���еΦ���s�qͥ�����.��ʛ���m�PpC�
A�G�8s�cb[WL��H)U�)��eA/r���v��gn⧕��w�Ǯ��K�nW��GH`�G@x��ݛ]5�2����l�)LJx��H�gp�v�)�(�ݵ-Oړ��q�-AnK1��Ɏ�;@�`>�E�y���{����ݐͳ8A�����}m�Ͷ���)脄�����-C�C���w��x8��Se���R��9�^3�7�w}��~nT�������&����q!�z��xgA�C]7Tod���]Q�O>V��s�zǥ��9�n��<�Ae�J6� ����љo��*�C��~��*��#c6������`��;;oS1���֐&ڴ�L�~;(2��6��Pw o��_��Ӟߏ����������~=�3����g֗���魺�Vkv�mu��Y�/��7	*#�kfX5)Q�Q�ZG�:;�l2���[G	RU��uf��v��TE��V[��W �1u�V]v�-_4B�]�O�����Tf�@C��J�l�����m`R^��8��3��ℳhM����foB�[�9!�ws���kR�b\�v�s���Q�[5��&7FV�^�D	1'�.T�`P;�3��	:�� �@�y"�v���T��lC���Vok
�n�ٙ.N'G���a�B�wI�V`�z�*�;�zƦs1��x1C!��2v ��})b�U���9ϊ���*l�يk7�X%�×n2��պ\�K��6fZV�u5���i������x4;�+��a}L7]�#9�[�!��Ev�vE�T�r� ��5�m!��f�Q�Bn󈳽p���S)-��;qs�\�N��u�+屻AV��ř)<f�^])���=n��٬�+�`㺗�5#Y�t�Ø�*g�_Y����c2�4�R��ǩ�^)���U�&S�ZPo�ĵ����J4��f�l��e���2F�;�m+vY��:S����#�7z�`��"�>q�ˎ�5/�̦�z��r]r�E�:rn��][�������-�x��Y^َ����sbb�NۿgS�n ���2�dPh��b��j��}R�����*u3��ʴ���/1�S���_�Ֆ��כ����U��W��^�)t�F:����x��j�0������75j�RPꑹl���T2���g�WE\�����3���Y�G:/4���YK�����4�Ԧ�{�"����:�v��xjg3�H����>��3�x�5BLF�mc��]:�Z�TW���c얲��aV��}��� C6nv=k��Իj�As�*b�^&�Z:7���b��j�!nX�������G)�sDͲ���&���$��hnqq�ͩ]�Rg�dV/�s��Ev�Чj�{k^U��Yw/z3:�)c�f��4�M�7���&�y��7�l���%�ɫ��6�(�o�`�Y��A'���Wi�bR��$)%c��P5�T$�!Ydy��$�ԛ�*&5���5]��,Lq���J�#8�XB��=�t9�Z�u�U���a�P���1T}G�^�R�]�T�e4N0+/nƊŴ^pʲ���/���k�C\��ϧW;wp�,�02ISfֶ�Dr�$�R;�{�sy�F�8)+�F��u�L�0*��N�=�5΋1��ٹ[!�o�˲ʮ`G*T��{N���k5�J���˨Ώ�*ګ������zx�TuE�!n����;e�ky�bT�7�^�3 m㨌�2�2�Y콐TM^���[�Z�u9�������1qd�6vip�#;���u7����;�V ��q��y�*���7&���1X�א�/P%�LTKHDISMQAMLJ�QIMCJP�dj�)H�FH���	������(j���(�hi��
���������\�4'*���5�b���U"ҍ4�AABSIIJ�%IE4	@P*QJ�3���h&�)F��)JhB��
J�J�"��bF��������5Q-S-�ZӤ�v2핡tM�և�2	h�4��(
�A��Z �JA�@��Ц�A+�_�����VE��T+ʊpM�fA���,�M���e`]�ڞ"LN��Z�v50VWp��;Ӄ\�x}�9���sW����u��9B���7�D�ϫ�J�`��Ez}�D�� �U�lS��?��~,�����$����0�{�V�o����0=K�w��[ �����-��[>Vu�kf��k
�sh�Z1�{.%��t�+��5�Gc�W=����x��Q%ٲ�(�w��w^;sT6�!A{6Qzs�'��N�.�L�2����y���ȸu]x������!�r$�wst^D`9Lhe'%��0�7��O��Rr��E��9�y%:���~�N9񮋲�;��N��`���z�&�rsry�=�S���j}bӕ���]qxz��a�:�F�<V?㭕J�/U�~�l7���q1�,��u\�u����(�P�#YC��?Zv�`Й�C��ޛ��u�[��xwl{�<0#o�a x�^�Z}��S��@�WqX��f^h۾r}�4���u<��|ja�,l[�6��`��G0�C�yXC�E��/Ի�>�^�������p��7u J1)���잟WX5\�_�?�C�u�0g���L[<��{�R;�.ٯV�E[�����.H�j�%݅�충o籕���\"���
����㸀٘�8������5ev�(ஐT�~X���Jmds8�	8gE��w�0g�;lw5n�G{��s1h
�2T�&��A3"Old�����z6��	��QjB�v�:��c��a�'�{:<��I��Fi�- ��@�Z�/a�G<3�Ӱ��p��k�#��E�0T��-��Lu�[������	�/N�eش��q eϳ^���:j�������ai���;�K��Kf|���E��<K��}tj��t{��j����%ڂSl�dH��K��˨��빗l��vE�>�S�fȧx���>0��Ƚ�\���kZG�BA�hC/LtL�9��UZ��pld
���Q�g͋e� [:~iw�H�	<��=7y��$I�[�2'0g,F�g��ʙx� _Z�(A=,�,�$kY��|j2��͌�̂qv��˽����i�M�N)�d/g�5FA���!�9/)��hR�T�SP�q�uEê��3�-�W$9�.�6�v8N�YY��
v܇b0_Jnf�L���{#B�ʢ�]�N0o86�jU�-�ב�o1U�\Ų��Jw|��C�Z}�p�n�;pl��nԩ0x	��sȤ�pWp�M����tT�N��2o^���n=�`"1���S �y�d	e]���vT��>q�[iRձ,*��t��yV���x�Q��_��Z��|w&��+S "�â�e�uwS�nZZ4�:���2Ϛ��ۿ�5 ��QP�=z �qu��tѣ�WC��R�9�M��9�6�Th���O=��/_#�+ ��M`����=S�	 �6�`���nܵ���e4�����zk��������-y�7sץ�?W����3o��8@�Tv�C��n��9RS�P�r�̈́��Gf&wvnr|��X:n�D�\�8G���Zti�_S�-�f�QF%k���Qak��Mx��)�9�L4Ui�@���xs[=�H"����-5�]S��"Ŝc�Z�XHM��E.Q+\u��\�9/LUG0�v��W��aߣ5����i�an�nm���p3!Ca4�t����Û��@�~��;�B�^�C�g}i�������\�ϗm��BK�-�3�.�����ƀ�����^�~��^!�.���|�w93e�1�ۢ-�����9�����dUh�/0�Tm�28;��M�3��d�k[zi��k��!pz@A�F]���eC�m����	�"��H��I�ԥ/<𩦫��fU��ay>\�L�ƴ�2	|��r�F���N�:b��<����A���N+EB#sC,���.�~W�Ʒ�=��VZ�u-�@bR��Z��*:��oN0�F�/�|���ť_�����Sa0�P�=�.�F�fS�(լ��;�>?��U��}	�ȱd�fS����	yX�mx%����`wϊ�JU��R�{2���S�<	�{GF�.A�l3� N���[q��6#ܬ��U���y(����U�h��Hi��2��t;�_C?�G1m��!�s��K�j[�����LȬ4)=�;B�s���=B��1(�6f�u�ȼxj��3��֜I|�0�n��أ��MɌJu�1ܝ 6퀔l��	?�ӿ����q�C���y���C�[9t��xL_������o'��.�5�l�m����k��I�<9�W�4�P���qA���k@.�n��"\������:�O6n�k>a�|�Bixb�"�Rt���R���LioZ��|4�UQ�a~��g �۷��9u�����,P��|�P�`�(qG���O�iAb.��IĻǻ`>�ՠ�[�*�^�j��:���0|b�O��&Q�%֚��8-`��gUW�Eʎ�S~WC��,�~�mR�[��eg!�
<K������8u�?T��j�}n,�2������`�%�]�}�T{*L��m�]�ֹ���l[��0�<p�G�v�M>��m��1L�T��7u�*Xj�����UOH%>�z	L��f:b�;ᚇ�h�]�5��`~����o��]+U{Z���~�B�����k����͉ώ�W3C�F��( 1�o��߰^'n���.��<����2Y�,i���G4��I���[�v9�� �v܏2��9��B�Z�k�V��N�Z[��GZp[u�"f���-��YdNU��$TP�}N���S2�|��=�c��H�r�LW��b���GD������Ƴ���lN�]���Va[�z3]&�ݬ`�y���H�i�K跿0���~�
٦z;��ۅ��'^5O�o&{˚�{��i�Ǟ9����ӻ������4��C�h�(+.~&lšm��|*9�y��j���,��T��!4�����FS�S��ɛjԕ3i�A��8�1�}S�K�5�R�`d+�k{��)������o:E;�ama�}��OP�X�+ڊ����M�\��&j���X)���s��3\�(ζy��n�4��zkw�!�2pD�����j�ծ^!�bz��VիF[8On�d�N(r�d��3L�JT��#��|�ό��%���?������X<9ʓ^����
B��! �c�5{�%�|
"K��|���U�l�q;�p�������Ep���h�rf�^�2Ͱ�2��v�8�{z�$��S�6�k�sQ1����1m$�i�Xp���ye�)�0�`��:�hLpm܎iNqD1��ڞ�ŧ+H��� +�<���L��d��!�X��_c4i��B��%��ѐo\ͦJ�i��T�W�"���u�Q1�[&`�ر�� }�G{Y)6�φ�3Uwk��J_wq@Kd'W�e�y�R��1�����Yv/ACGK#/� ��Ŕ�A�#u1�J3P�Wòi��0��[!��i�0��˞��i��Us^E�8�EO,g�[�zzٯu�w���u�Q�����t��v���� !�:C�y�d�hOP�uf�S�N�O&N9u���c|;�K�ڤ�-�������f�طvm��p���@�!�ȇmt_of���LЧ�*��::��)��omVJa~��y��s=����ҏ˝Y�P{G�[[3�G�E��-�:���=p�.b����xJ����T��N	��
��P&+�j/��x�� Q�<>�jW!�32�:C!�1�/�r��]��m����t4��t_�������>���+��l�N��kf�w<��2]z�m�W�F� �斘�:��m�<;��7u�f�&p�a��Av�|e��WUsө��CXdV˴�|kO��l�w�\E!��["�髟WXݭf|`Aƻؗ���J31���-��b�����A���=��U�-�<�ӼNI�C�=0����OL��%΋�܊�=��됲���jFO�xa��2Б�g�c��eE����f�>q�{fr"~���j�yܣu��u()��Xᢳ&���p���#1�j�.4�87ӊ���-��ԺH�t*E����kK��P�9 ��N,�ptڎ�T��Hof:��oei�W\���0T��<�M���GcU_CZ��8/���AMk��{������U�Cǉi���n�����A��Jv�ӬY��}�� �ɊN��J�RaL���T\:x��9SR�ϙ7Gn:f�z��-u�#�������i��p�_Inj0\JgOf"S�#B�ʢ�\n��썍�"s��|#�)�yA̫R�R�h�8ޏHQ� C�L9��ۃ`���)�x��Wqq�q�AC8�Ӱw�-
�@���(ǡ���S�!�!�O���|�%�a�n���M�T6��Fu^Ρ{*��j�d]c��Z^��vng��8{�<��s��A�{��~Q�Q��νa���n��琻^�I�,���7)<���`�û5zF似�|m�0t�_(̂v����#Ze��X��X�`ĝqv�Yax�q��WZ�Sݾ�58{\0jq��2k��u�n�l6&m��:c�zG6��4-XQ+\u�?J�T��_�hlN��L��V�3R��˩���Y��Ն�[���<���:a��sBv]���Ú�ԨO�Z���Nlc�J��[r^z6�j&;g�[^ bz�=�u ȗx�`<h��=3���jY�~��,�'r���,��C�x�(��C)!Κ�j}��w�r3��%WM��h
��[����e��a�k��9L��;5�Ǐ1&����%���<����fohnKE�èU���N޾�?���H3��o���ĥ���ř�b��Sx�(���q�ۯ��0>!�%�'?�!��6[��˱���:��ևt���ݡ>0}��E_c������^�n���%������l8"�W�&��l� �\e6^N���Vo!�p�F.��^k���ͺ���m�^�W!F|�.6�5{�.W�)��Qa�
_L�y�������``�������<��J�9R���FB׼0�*�b��%K\={y�%o��rx��n~�OX�G?y0v��	�����s&���'5��#bև5y��M�L�ʖ�3��w
w�i���í���u̡h��ƚxk��Ё�iN$�P�		��ا�������i���������w�k�ܰ��-�`Z�%B�6s���xOB��Hqm	�����|#<�l^��阤TMf�n�~�^@N'I9��,���ʒ4�S�_8k���N�N���I~��k�@�x��;���7�64���{y�J��0��QtÔ�.�tSz����-���57f�*��3��k��w��K/E-�&1��B�����Q�]/e�?7 �ƗI�栜K����es�\�N�>�5�
�p�2Ʒ�/�Օ�����뚐�ٲ>]�D��LpPE�
�AfH3kR��-qn�gt���O��͠d� �
��袰)��&��H���+X�ڜ��+GgG-�w�:�u�
��D��&Ø�^E�}[Sl�])c�{yI��[��_?0�_��Z���4'f��56���h]���զ�w:�WC��K6!�32{N�^��s.y��X���f�q ������֯A�WM�e�Qkd�N0��zW?L�h1�x��	U�D5���q�]��h�PQ�΅U�ʊ�K�Z#O��"7��8??��T/~�琹���M�eUp�ә�+��+~���עfy��f%�3������D"�:�]��3G�P(C���,ۆ󘾋�������HY$�ArC��LW��b��!��D��Xlv�	wt��Uə�p��
��X��1��`�c;�����$@"x�v��-�#W�n\ͼ�tF�u��Wϊ�i�sM��� ���5�C��'������;�i�/��=䮂����[i�4u�1�n6Z���"�XJ|zh��@c�<xX�ii(M1������Crfڽ�*f�;(5�`�ie��&�$�Q-y�c V���8^���t�w����"����J�`��j+�]ȃ�B�~uK)�3�
[P�(1jXbi<��<z3�-��վ;��e��as	~a�5O��*=��]�_�d��S��0ɻ�����;O�{c�<��)�U��v�Ѣ6A�xʽ����#4x9���9LXr����IBUk.�46�ɐ;��.�����0�(l��:�4�Y��u�\ʎ�9�Υo%�0�>}l�:��vU���SRCnR�4���A8�>$��b�+�.%�pN0�՘J��yV���RJ�c]]��O^(�f�|`z��'���S��D�V�E2�$i5��d�S�\:}a\c�!�3����&X3a��ͭ1jY��c��gd�q;�i'�I���Q�-�a�i�2���˧�5K����U.��y�CE�������Bc�l����uL5�mO�b�����N������]ʧi�'�`����l�Q��Wũ��y�c�?=H/ƳO0������F�x^JAn���al�����%ݠ�3��6�?sȇb�k��+�L�(��<�"ݳ�W[����fϞЅ)9k��y�s� �K6VŻ�l�a�8!����օ��i��J��;ճ16�K���k�P�j%0��/�^���u��c�g�������� +�l�Y�p{�9�a��u�-��6'�Nç�ᦃ���df�W�r��������ñ��G�(���f�'(��������"&9���X���w&$�o�˱n���{��>og������{���o���<}~�W��:z���48�B�tG2�ƙ,�n�}�ƺ3��n	�HpȔ����.�2[��o�x3��/�o.Ƃ��r(�ݠv�\�:��Q�S��G �������4�k$M�D��a���i��z��j׮�i"��s��F��:y4�oAJ��y7q�n�.j]-�APt�z�k�av�Z��ۣ)jtR�g1Z����J�H-uv,��>k���g1�){q ��7u��'�C��s� �q햚���n�z#� [���u�f�s]v��O ��gpU�N�[]�īG�6����v60ʈ]���\O�1���c'Tr�E��k0s��\���ʣ�@;.�L�`�'<9k���^����\�����d^cvӼS��3+� ��R�|�X�V��7o�\�\9�s6��B&�b٦ˡ�M�1T�3�ܾ���:eWP�C��Ǵ���jg*�WM��wo.�5�vW&�o�P�]7��T�Y��ڦ�G�>U�������QCr�CDm۳����:��9$���|���q�U�X��&��� �,�X.�w����|�l��T�Nw���>�)ۛ �긔5ϩj�:nr�Z���L!fʟ5N\���y�a�B���Ҭa(�o�u�g/9L`ǋՄg�T��Ws���횔��g�-�#9�����
��V�k���tZK�_af�|�UN�U��q�m�VCmi��T ��	)�y�ſT������.7�C�)��d��k�%b,Sh���A{lr�K	^�Tx^�#e��5��
}��w�s��G����e`�#��*won�@��N�xM��^4���.�K{�8(�,� ���i5s{�Il87��
�1�n�b��]��r��L�%����n�� �kYi\�ٽO�h���G���	��Ntm����� S��j�B��f��z��g^�X˄��k)2���$r;/���r�ᳲ���j�V*t��\ t��(g���mn�*̊	�HWi}�;a���TU�+�\��i���u`�F�Jչ���fŗ[�|�U����-Λ���jM]|+.�v����C9ZѦr�-�ss�L4�ѵ¢Zh�k��*s�RL��
�:2W�B��n-eD-���νK�b�ͧń�ù��2`t(�3I��K�����[p��m��H�J�FQ��ۼ�bչ�B[E})u��+mj����L!w Z7Ai���뛺J�ɏ�wƻq�d2��6��Ν�S������wU�0����;��L$�㓅2���)��C���$���G��H f��8a�^�Q��ڻ�v���1�r�v�[!/����!�44�������$ԣǤ���
�k�q��'��쩬x�2v�!�^��3�<��V�:�Ǧ�5v2@�4�u�q�;� ��%���Ʒ�*GJ�i�ܭb,lJӕl���Xܛm�R�uwK,�Bf}��@Qd��&) �Km�醐L0��x�<Ǝ>���4��H�()
���SH֊)4�
b��h�(��
��V� (�.���J"�)]@i)4B*�
����a)v��)Z�Ӥ��62�4�!CB5BQ�4�TP�4���4�#XӣF"�M-F��4��@PHh4�MI�H�SH��i@ZtF�H�.�
z�PR%�ӣCCB��4.�Q�t��t�:H��ɶ@҅����s�7�E��[�>�[׺�L��ع*H��������n�'%�3I�r���Jk�� ��Ccp��4�mpv�Fܱ��h������]W����Ur�0+�\k�SFN{>�ǐ��h���ubzq���t�2̳C�FY�i��v���b:�3�z��IE��Q�i�֞�<���l�w�_|�awX+����˾>�|�<��q���W2�l�<31~!�XI�PjQ�g͋e����K�X02pBOq�ѽR`;,�Y'l��7X�^�!3��ȫj��!>�A9�YRF�����Ƭ��sn���
�be۪�8؅G����2��|�4<'k���-B2;s���A1IՌF�+�I�2�l����g����Y�v*��1��"y:�k�0���K�	�����2N]�9�K�v���I�ӨFgK��*.5�-�[�ADַ���iq0�2ۇn��0�;�Rd�L_Q��ӏ�z.ۗ6��C�y<�/ǌ���@w�xa;�-(!�B|�xs׻ K)�`��L���۫N���i�j�q~�Mc�]6Ⱥ�09�-/#h��=;�?;�����0�7s����Euv:��w>��2$�z�����-�nRy���Gfjxwf������kz<��%A���`Ww:��,�t�('ۋ�t ��M"�M郲��ڛY�W6w��~9�f,�1uvJs���yVj
�FyO��9�����Č�����<dDޔ���m��YtY������+���ݭ৷���I�
��S���i���C5�[De��md����|"2/^��.�WB��<�3�U��y�ں���}�_TP�T��n��\�X�-�{x�����T��CL	�	��C�е~Q+\u��+��/��q�:m��%J���8��ܻ�����V��z������e��Xsp:�a?Mk�e��&pQɦ[�-�i}�N�\f���^�3� ȗ~��t�#l�fI��Y��{�l�vr���_Sl��#��	�c�D̻HD[�@���,������x���
jvL���^�C�*����d[w��i�G�vp�X��C�Pi��O��TD��%��`3?��h^���9(͵�M���ws㷙��p��W=�E��Xݍk�3�����Q�b8��[�>2鋇I��KG1�f����8D��,~����BA[��~���ʖ���HZ��0�+U"RS���͔9��/�Ը�=jX|}ꛗ�� h��F	��!�#��F2\�H�C��Jl�!2�ս�����6��S]ޡ��w$V�f:�o4���1m!8��@L��W�i�b�`�ز�!8w��R��Ȥy
�+RԺx0�ޅnWv��(��R{_�����w�ݍP>F���@��q�b��H���)O�>Uw]�;�_nQ8k���h�j�bF����sM�d^��%A�O�=j� d��wD���.���]��T��t������m.lwʿ�g*r���k���o�j~�T�	�%"�F�c־��z��!��d���!ꐄ<MqM���LŶBY�z�xg���@�d�`�eA#I�>���L��h�Ơ]�J	�S۪�������W:���c@����<�EL/�J.��)�yoT7P0i�3�wkp_:��=Bk�J�f���R�h�f-0D&�	��#�Уg�C��qWKг���K���?#���iV����R�B����puk]B��\�#���֘B5���z�:�S�1���ZJ�/V����s�i7�U$�v���ց�Adi�=8xr�F��a��k�N�6��U�W�*��eK�t'��w�Ϲ��PKܼ�����B��r��Իā���2�����nwqd��n�<�U̓?K��}:�	��;p�K�gc���x��rl�Ҩ>i�tv[ơf�f���O;��ݐ͹�$�#=%�Ĉh��H:"صu�v3�.�9���~s�/�)^_Ox�Z�z$ͧ�{��A4��ci��$=!��ONŰS�`7���yu�o&����mq3�?��u��ca�O���B�ɕ�����qTpm:�҆Y������f����Gf9�=c~ ����\3��#�����W�;�${gWB�2����{����ԝJZj����h�RyLJ�m���yH�!b��&�cw�]�P��ĳ�M,�W�6K�$�9�g=�C�wp�4P����J� �M#70s'��F����C�g��sQE�[60X.��G�6�\]n%�JY��=)ص��
���j�<�˃b�8�X�rFl�zǫx]]���XtO��#�h	U�5e��ij����&�{Uݭ�E�r�q͈R�&���'�Fu�ј�oV�^����0<0��]1#kY����oS�M���/F�nr�^'�X�2Z���|j�Ξi��E��U�s|���;Mݎ[]��`�S�Ɛ���O=x?D�I��"S�t�eA#_�����YP~.��ԦO�g��p�6�PP<�:���m��gò]���&HޣI9w��&�e_�&=J9����sTT�$-�4��v�ϸ�l D�}"��^���;��E��i!7K�h��f��!b�wn��~�`qs��5f�HXt��<� X`�Z@�#�H����q1���C�}�u�~Q�^���R܂2SŨ�'�r��5
3N�#b���j�b�quH�G�~��+7��C����Џ7m<%]��vW`�M���5�J��}��gԭ�]F�+~�[;[3�5ES+�x��g�`~Ȅ�ol�*1�-ʲ>�t���n*��vX����fɛ�VFt�Xr�g���LAd����ٕC��V�����kx**�7�8�����,|���sF��x�7�m��ʀ2��L��t�y�s��l�l[�4v�>��2N94c�.ָ5K&`�u��ˢ��-��H��D�E�Yk߉�uy���H���B�3�٠��E�u�n��I�2!�8��t�ɕ>	�r�]��Q�I��Xq/ �/<�Ьi�P���gr3�7���!oa�F<3�������T��_u�w
�1%�����"�8lI��Eܐw�;c/%�'tE��S9͑.���h.9���I��\N3�=��|�ن��ب��SL�f�6��f�5O��ڊ��O#.ű�>{�m�N�f�`0&|�[��E�Kȵ+*�X���5yZ��O^���hi��=GA!�_AX��.�ՑC��| H��d��ySJίCzh�yw��I�`S��=c�
B�(wd�U��I�� ���ʼ��g��&�*��F^3ùxg��{Ow��H��g3"&7�4�� a�dώ�ۜ��9.�o��Ҩ����	n����q;�F��+�Z��0[K���y�����u����sP~�Ƚ�2�����3��tʼ��Rj�n[�>SJ��W?W��xղ-��P�3�c.�bI�!��e"\Y�p��o@7�<�Z���-�-2-ݣ�+.�XY�LIvU�+e���[�L��6�V���.;9M�K��w�I;��(5P�](r�ݜ
���m	;3|_zo�<����g�lQ>,6��{j-��N7�5�x�AĈrO��r�Z�Y�r�G�d�E�o��ޥ.V6$�c��B�ܮ4(>�s�]<0����~�0�X���W��g[�0�j^ĪNT��	�d]`�O����zk��6����G�p���L�u�}[��CIu/��b�H��	�@9+�Z�f�'I��\nHO��y�pә�� �UUf�'�����D@L���Eњ�NA�|8�,*�O2�V�L'���hhЩ��<����;`ÇB\0b��	�tdd{MVJ��J�
�^ۯ��("�5��?K]���-��p���zs�W���y�
�ft69��y��ry�n:�7���؇曭�xA�u\o?l��%�b	T�5x������t��**���H������Ķ�ead5��ϔ�3:ۄ�b�\�.��1��Lȓ�-�tg/��046�i#qm7<���l�4��f��^���]�R�5���*����.��PU;�d0tE�3����x7��%�x�'�XmaI��v��9oSVK`�'��vWlɵe~���JN�N���%f&m�p�(�]�AYV7S��NAʶN��8�Q�Sh�U���oa�mǏe�V�����v����^N���WggOM���3o��y�O�y2}�
�p�.$C\x�zl���[��xj��I�+��r��c��jE�=���>T�L��;X���u�~�h�h���Iň��O2�;7*Zڴ�^�����Pgg:��B�Т������Ŵ��^��Yא�msL8�v�S���԰�4�Mwc�w��Vn�.����O�߱l=�']J;B���{i���Ol��KHN%�b<	��D�!6���xL&�>ޮ�l�1��g��!�#�	�O%BUA��F�)�0���TFIH���~���_bx�<n#��t���A���M�A����iCe�2�a�*�����;^�tms�F�@i���t�� n�nݽ�z�=�]���u�Rb����,��;�(�}6�7����0Ѭv4G8m����\l�uC�� �m�0Xy�l�*��]�;V�Q���gQ�k�n���#N��i������z<�oH��U�G��m=d%9�2�j���rf�y��{1]Um��D;�KT�ٮ�d�jYR�v^��X�8|����t�2ױ.A��Wx���~��+B���E���w1.��NkN����kU�<��\��5��{����H*ak��;�G�E�8�z��AB���O�*l�����.��58�y)���G?��1�ê��v"!�wB��H�i�{�k�ds����m� ��@���9�sU�Z�L��30a#r��f�ka��=DAm��M���s�Y�p�sl���:2m^ө����ט���C%>����a*pv�x6k�؍n��>� �"A�`i�w�ɞ�Nz�����������3���Ю����=�wD<����.�yj�?��zV��Ƀ�������}��9�Q�*����nE�Vor���f��֍��� �#I��#�#6ԁt��=}�=���h:�9Ȑ�!�b�"Ηm�� GB��(���OZ�{2ni��dE:M5�/OX�U�Q�D�����u��2�v@��a)�IU�����U�{��&a�Ix���Wo�g2���UA,��"�!��Q�x&�*����z4���o�w4��S�koR�����XZ��6�;k�а3سԆ�e/�=�w���v�E����i�i7ֻ�ݭ4�&�+x�S�IC��j��F����܏V�JDf=���ɩ�ee�ӄ��b��,�Ɲ��_lT��X>�%h�r�R4��wghf�D��WUi�� Uʮ�߽C^�62C\�M~��xҒ�u�y���c^��까$�ET���6d6c�۠�Ð�}66���OѮԆ5�D�A�$v��w�5+U.Vɽ�9�{%O���r[F��][V����їV�d�2l��e��WI(��w.Ǡ]��#g?Ryu�C��od}��r�+3y,��ZzU0r�;6��n2��"2�" &�o�ҏ�_�0F������K�U��y\�H�4��
�/�hq�nvP͘s�_����ȝ��\;��q�0�7�&",&�k.�ó��;~��Z�����#�El�r���=���O���3,|�[�.�u�Iw�Y�)S�	~�ֽ�gY¹�����P��;"�a�Fz����y�&ٴk�/�a�c�m��n��Kx��8�7��G��G�e��2=��� !D�Qǝ����-�ɢ�n�hc������En0�\��P@��;m��|,ȹ't�:-b���?:X�U[���:WF�V��u
�M,�7IWn��'�����k1�q� r������3�SWV%��I�ؕƮi���.6[����û<[�������2/��}� �*�%�=YJF�u>�~�Q�Y,z�He4����/Wʵ��U3z�FEO��|A�(��j	i=cV>꾜8OMy��38��tTC�re�d`��D�Z5�[�WD�&�M	-Xj�F�k=
ym~���]r����U�j���v!!|+V�m)1�F����;tυ�6N;��P|��N�ݙ-$.���3r����a�Z�����"$~���I+�W���s>�t�K}����n��SdB24�D�;�`����
8^�H�.%�)��� �����F��U�Gi�m��3��a�u�G���U���I.� �:�.4��_E���S���-�0������U49�9��Z�P�1�霣�5�N�^OF�R��&�1Cv	s�j��J����ڶ|'���x�G�����{���g�����_������i֑4-��
�!�/��ڋ7^��!�c�@{a�ͯ�H��tH�ĺb),⵶�@�p�w��� �yB��
�{t�j�`���^�gb����A�xS��ϸYo3+aBQŬ����9�Ss��h�U�;���V�\�3}�����-vT鬍�~��c��F��=[��=tu\�����8�֓�ȯUs���DZ+�Q����&u�_�=��*QM�U�19�دi�fU�d�أ��un̓d��7;�݌��T��o8��}.�.gl�x��X��nh�{Z���6����� �&��k�=m�;�5ҕ�2��v�3����c{����Z�:V��`Ի`�`��6q���2�V�������$Z���г۝G�6.�7u#G��Zu������F�u:������Mju9nӝ*��r�e�7���kh��`���a���5��T2�x�ԣ��;&��q$�V�{V-��9��K�m�[�pbi�7f,��	�Q�˶�=F:/��FS�k��|�D8�j�x5u�=P�Y	�ƛ��zc��T��?I��b�b�L�Ԁw��둈q^��\Olv�k�Z���/��Ĩ��ra��_:	Uێ�9�h�%�]c�����-��=�l�m��5��c��)]�IeL���7+����iZc��b+N�(��8q�r2�/{/���s	w �m�l�#��-䭷�nڴ��Z�i��\e�ٺ��ƭk�D�sP�r�[I��>�5�yQ�U>�au!�B�*�����������u��lT}AR`Ք���ݻ	�����}&<��ߒ�:�n�/��t��U�T؍�!Cԕ��b5�s�e
&��E}b�M���㫣c�p�ʮ��V� Æ�Y��)GT,tz�l��Mǖ9=�p�]x-���p�.�,=�?��T�*�і���|(R��uNw�1���k#@��}-Zn��V�.&��5/���YnR�m�c��YNW�z:�]��,�K��-� ��}�H�9K( �ʉ��W��a�$�۬�u>���re��)S�h�3���TŐ�X�����M6{V�����i����o/��.E��^��1gQ�y�cWcm��y,K2ɭ�4HYb����!a��{���.�X8�I�2]d��Z��T8+����7o6'v�Wv⮬��u�����J����i����=[X^u����˘��µ�"o{x�r�'Ϣ�w\�`��~���B���M��h�bծn�mT2�t���<y�+U�=�H��i���e��6ڦ�u�ݒ�ב��a�(T*��Gx'�vb�OMU�uv��a��F��e�wV�ض�Z��R:Fm��B�����v�s�b���[��5Kq��ĦJ�覑Ǫ��ʌ}t�c�M�����f�-(p�"rN�sK�0��e<�Ո'��u�ػ��jYP|��l@7�U���\W.9l�EV:q1N=�����N:<��G]`���M�4!�l�41�S��-!���u�)i�)�4N�	�i����8��4�Q4��4b�5�
�l-4��)CT���4-% �@�ҭ&�
WB�Pr"�:�B��
-�#� �$I�4�C[e��MPT�4�F������(
l��J��" �
(t�"��$+K�4�iZ])��端\���z�z����c���J�J�>�r��RY�ʥ+�����f��0�6T����6�t�7��qS��.�h5ܶ���}_|���������iG����St{}�vΆ���w�d��p����A����q�;v����#�6Gb�h1�G>y�����}��N_��K�Z,^�LՎ#��q�$a.�	1��M9�t3���U:Ee��m�-�"O�'��ķF�e����i8D��h8+@h~�u�509���cv7SP�ˁ�/!����n���z�ܧ�y5m�<��au��"�b����81B	G��MUS���d\��+laA(��S��t�Uq�ˋ޺j�J柶��PF<���Gڝ��-��y�����H�>m	�0�k��F�Uo�M���2�d�q�=���v��7��T/IA�sȞJ�$�����P&��u�E��yfi�]�=��x�1F��k�wJJ�^�A<U>�K]:�7���s�/kֽ�B�u�)S���6ʬ��kJ�=|��]{]r�>��*�x�<���V�C�/W*�=��\~�	����˴��Qݩo��W&C�Qr���U��WA���6�����5Q�1v�I �5�U��WY�C�w�-I�PC)����u�ٌ�S�˫�A���Yx��X�H��uf�wO��}���j���70Y6ǘS�A��#V��I�q< mloI�VۭO<NN�R69�7U�30�p�ܼ���ف�� 0���d?��7�{W�]�jLDlr��;o��ps��bc�q�'vM��i��3�7��N��Ρ��TTd(.*���l~���mRIux�j(*q�"�S��8�.�z��מ[��яك%(��#�R�al����G�� �I�:Cn�)�#���y�F�i�19X軀���1��۽�� _�Gp~�$��F��j,�ہ^+.R�ሇg�J��Y��n���$�Xٖꍰ��i��=B���x�d3�rf!0�OՒwݯwD=6�ey�kzq�GWsvRԕ�Z*�O�)̌�{ B	��©����z�6n�y��叱�y�y��;[���u5����z�[~4A�'�4��jU�6��x3㕭����-�D��:�N�a��j��L���qw�� �i��������^+4Ɓ��f��]f@�^�\�]-��Bڌb_V���jY�LH�|��پ�n����@�I����$���oZ��P6Y�.�=i�&���s�u��lg*��u*;�T\d�$,���pk�ظ���g��^��D��ֳ�ឃ�P�� j�/kgͨ^&R�����������}z6M�=���x�?�X2��*D�ۍ�=غCjF�<D�Aig�`��1V��y�z�����=>ˇ:�@B����
F�r���4�J�k��b�q����,gd���l�f<m���r�pݷ7�B��߷��k�����>��MxK����-pck���X�Yb7�v��a�3\��q��܇�dg]�5&��3"��ȮIEx%�+���-��M�
2���+�yu&�=�<k�E�C�R�[�(ҏ*���ëj�2�y��]���|@"PnO�	)=��V�+���m=�@�ן���ŷL�C{�v=  P�4��3�׎�g$E��J�*uf�k=猪�Q�}�.맶��
�wswp�L�1���#}�K��v�*�w+��ؗu)������bVSsFS�oI˙G�P�i�[k:���@ ��z��	h{�;#�i!Ts|»̂0e�;��W��]U�Y��5�0��ص��y��=�ٕ��2����8������}�9J6-��Ý�-�����nRIc�OKv�af�8B���E:�����O��F��yF��x�)y�e���x�*�{0f���KM,p4�y����� �gj&��fd)�_dHO��Y*�[�Q��;���������}���kUBɛ]�F�q�#����*U$q�~���L�͈߯�ՙ�2)C�U�Ke�������L�$Z�h����	�Q������^Ge����/8^�x������tUD�O�=PEȄ�{�| V��i�������*�kX;�͜�-'���x�e,�庞̉�pBn�%jg���/��^>����+���$���%|��q>��ڳ���~�R?_�H���o����H��^~AJ��/��Nn�S�0h����a�щ�-�=C!��t��I+��`:�m<�y�R�LI�u:��a�:���ys�N�e���;�i*�o7,�r��(�;bb������譳��l�X2�TXY�M�wH�F��y��yS�c��r��J�zW�p��:�����[��u8�� �$��h����.�=�c�Ī�.��I��.���u�Nf�Ľ��:�ۇ`��|���K{#d�h����\������7�hf���_$o`l�|����'��;]1���M$���K�s\��K�e����q���u�J��ޝ����MH�a
��Y\V�����ۓ�����rM�z^�u�g{��P�������s[72hu�!f�2����0fm�*�$`&#�WO��ߍ�/����+w�aɕ�8'a�P���`w3-���H�H�q,tIj���e��\�/�"3�u�>�I�pP����Dm]u��a��zw��5�{QJM�� ���G��1�+b�6�� �=ܚf:r�ؑZ�>v�A�,{v���F�<{��CUk3o8r��+���Χ�^G�����t�zk���~��n/?z�~^�k��{�#�-�:iXc�L�v+�u ѢAnX�DY���뎵KG��v��M�]X�&v(5�Q6ÈI���)�'��0���X��+�6�}`��v3N���~�=�G����HS�E��Pŉ\��x��s�TN�u�p��7��)*�F�9a�u�s5l�p�oS�
j�M��^�]<�k3氽v�'ٝÑf@F$��ISmU�i�	�H�M誻�bv���
׹�Ds�B�!|dwJJ���(:OA����se�P��m��wM��;�h�)nzx(l���l�V9R*ۤ������r���wT�TRۼ�ɷ�#"@Y>oF����k������<�de�����Z�(�q~�f;[o�/������|��f������L��g�|;�4��G�'vM��i���A��A��
�/"��7]yͳÓl�ݶ�g��K�QN	����>�O��d8�_�3e�V
�������'��6���х�χ(�;^&:@;p��{��.]��I���h=w�/�`�5!!cҷ��K6j���YUk��t/	��5��ꁣK�>�&���S� f`5k� ��M��@�`&m�O��sk#3]�Z�o$Mv�I��Ƿ���Ls[lq��$�:sq�,�]v��x��O�o�^h�[������*ؤ��Gf���>t-��u{"1�N�m��x�aѝî{�s>M�E�P��a|=7�#�C�h5F�a�Z��J�� vYy<H �ON�x����;;��c�JF�9�j��W@~IP���}�r�z��;�G��7L�^��B���	�9�yJGE:���,��R%�ET��`��[����������8�g��T8��jm�:��q@ކ��=q��RvӛY�Z�|-���2�hE�jA^�PR�$�����/Pxm�˻���9#*��z�o�1��
ߴ_����[P*�2�F��m���-�7�.���v�M+}�U���r*}����#�t��R49������B���9�s�{:["aû�+ė��P:�̍/ �6K��4��j��y�G����
�Gec��q�UtK�4g�q��	�>��0�l�cPZ�4�g����ޮi�{j�7�߃�
G��F`<5���ǵ;N1z�]}׉	kPg2q�Y}	SOS˭��.���.G�z�;[����F�WЕ	&���B�
�̶�P�')��-7��
�e��4f;]X�(��n9�5!�m�����rU�sj�o6������|����ǽ[*{����pr���6�20GtN�f����l餩�{-Pk7^�%仗c�!�mo�j���f��:����{�Nq�g���$�l�Ҩ�0r�JSKt����,��tkD�����wZ�k��l;�
K���	�Ol��J�`��x?ϪzN�)�c��Z��Ħ�{�T�
r�����	�:���òq�L��m$ܾ��ϝ2�l�\���b�������2���If�a5>gs�qP�3�m���x70��#v4f��Q%��>�c��`�^"r5�(�Z7V���7٘����I���robߤly�%�?4o.��9�4�ɞ��)@{�׉��̲H� �T�\0VR8�\�F'����o�������C8�}��0�MzfѨȩҖW��3�*S�}BzWZ�rB'�@�U���&7Hz�<?d��9�a�v���;�������z�$�-�|~䝾�c�²����y��JZ��P����\�{.��c�l8��,�֬ه)AsM̈́��P�h:�:��wa�Lv��l����z�\He�0v-�Ί�|�]f������� �,A�;��V�ę�=���Po�<�7��x�����L��ߧjO*;w�-M�i�=^PE�$ ��*�J��5���^.�D�e�{�<�@%�\���n[��fD�IxY�j:q��:��̮� ��" ��ݎ&�ΒW�*B\d6V�j�23*�v�Ty�0e-�Z��a���kV���ړ@v�u�U�Ҹ�@.���'��i���ᓱ*�t�dX�A��.s�:��bS�](�T�t��Ȇ���53M�so�:��m�7�=0`�V��*�ѓ��Cyri`��+U���V�s���ur�����Kl�a��ګݦ<)4@�o�,WU��sdwl��'�Q
��=M�7�4s9���q�p��m�ا~��\�s�4��Tԍ�9CLd��6}�p׍�0Cp-ޯ$��j���ͨ�v��AFmf��c�'�X3��÷��0�i�X���\�<(�J���pz��	*B��گYK�[G$R�u{CQRl�'%�۬q�CoV�x�(�늬k!��ڊ�v�%Jޔ���ZFd�����Jj�z�h�x�df��7���;��%�7@�՘36�ƈ�F\���] i�,YC�|O7�b`,��Ô�F�cr�:���o�t�h��G"D�-'��<$V�=v*$M��K����Ï��&�]�������}�X`��Vsf~�=8��'Ig��q��/ms�봎���J�ɩ��.)���S����x�ۉ<0�εZ� f��K��ז�%��e�
p(#��([\F�Y(��eڤ��Ƚ��U�GA����)�K�.���K��g@� �.my������'�cV0!�'݇�� �#D�U�IU�ne	�Fރ3�M'D{զ��f�H��9����L#��o���IX/	��I��-n^�u�3�=s���.�"�������󔶄�P:�GY|�䷕"����·�K���rI�3U9�z{��2m�0� �n$ճ�Γ@�}���ޏW��<��^^�w�����}��7����zj�.8v���r��%署��hL�����:������r�zI�ofֈ��:���	 ��=ʾ@@��9kĭs�'�G[�I�Х1� ��,+.q벴}�v���	�f �e�|�(qō�]@��]�[|/�7��\rB��V[�.�#�1�N�-g+_�z8��}���D]v�o)��趆v�Ŧ$�w��D��õ�@�{ن�LVM��w:��8����͢Ӿp=��`N�){Yj]N�΁������86�\�=��5�[���ϧ�]c�i%v<8+���_kT�����;�E5j��Q���{�q�m(���.aFc����o�ck��v�[V�6-�nVX�ݳ閔\�f�^L����{R���
<:blq�*q˨]�7:$��Pck~�+M{���/���~�o\ViX�ȝm�nXb4��HȞN�j��c�H�հ[���"�rA��Y�C���b���Jz�:��0�:�kL�:�#*��m��Y�틉�Ԭq�'>p�^_��V�T8�H4���˗��}x`C�}�<���}ZG(]3��zT��ø ��+;��<�'Kp�N�j&d8��P��}��r��a:�}N�U��%���p(�:���ߴ����o�]i�%���ӭ�ŷ�+W=��pB�J�W9�gc5�z%>u�6��D�эN�ڼ�t�n�Zd��j��O�LW�¥uK�j�&Y��k�ǹ������ix���7-����.�?"��p|[B�]ϓ�-ZE���Ԯ��Բ��f��ja��_9^�=�;(U����M�ǌ�V���*Xͩ��o�Q�F�&I�3�8��"��oo��4��.+�W���Qs�C@���+*3�P�=�����}���>�#��goz�7.���T��r��pR�Rj5-��)W۲�N���e;u|�f��X�="�k��ݶ���{Vw6�k���sv(*z�<y����@B�p�W��Z�k%%G��z{Q�eK0K�����-l��3�Nc�a�-�ˣ��-	q�s�W��f��܀�c0����#���h�ݛ�Rg��,6"�*�0h�Ӿ)%�T�f��x5.[��tL�@%�7V袉a��<\�s�Ѽ�;6�+�R�9����P�F�f�u���7N��3ǚ�N�:�O�}�p�KA-OA�B���j��\�7Xv��@ސ)���[`*��e4��Draw7
��G�h��o7!�M6��,n(�c1+{�'H١���:��6�H�Pq��Em+|(�Z5�ǉT��s���@*�.���޼}S�Ÿh���ٸց���X����u���x�h��55�72�T��K��&A�)a�eovv�s2�7ӥ|%��r�	r����M��{S��ڴӓB��8���^�Y�n�1E.���:�y�_ֻLK�_G�L� ʭ���ɷ5Z���[���c0QR�d:�Q�Udb�Q� ���*0�Qj�4�
����~KBr�-�ԋ�X�u���"�R����(t����@iV��l#�B�(�B���(�i�ih*�)�JJ�i(�N@�B�tS�tiJB&����R�%-4I@P��4�q4L�K���дh'�4��E%rt4R�PR�ѧT�4�B��AMbCd�cHPi�K�M:��(()
(*�j����R��MR텥hZ����A�P4�ƪ(-��TU-�Jn~p����s|����y��޾���.7�໣�yNoGd��[՘,�ASRa�N��n���'���.nռ��-����Ip�V ��dQ���fj]"���xN30ͫ��kyYQ�iq~[rõ�W@`����P/^��܊[�[=x.t7�J�Զ�F��X^|Nl����n2�O���!\a���,U-5���
�d�����zz:��ux�j(*tȼ���}\�E4���ɹ��6T=����*1*�Snnt�Ϲ��o)}�d��?*���0�!��t�*Nsթ�F2	S홌e��[d�z�����'#3��Z3V#l��]B�|�Pg��G�	�	3����0J��6e���+�P��1���ݫ���p Kgn�+@���u�p��B��G^Q��YYa�\��������{��	�Z=WJv)��%��D ����a�S[�(����ʹ1��Fg&T������:���)J�H�^���-��r�Y=�Y�SՋ9���B�
������=���q�5��t��$�*=�^>B_E̘������z�٘����l��Ͱ��w{���4��m�|�Q�� ����拷EV�C�K՗�,�a-E�{�)�SyAd���X�q=[�d9E�wfm��lRb����d�՜ÉAJ^��<��vd�P�9M�^��\�;�wq�Z#����s'gu�B6o�uJ�_:��Tw�5��ځD�\���7Yj[��/觡E���������,�B�L�T�q�v.�ڑh'�Ƚ�1����߹�zww��H��ꎺu#K���?M�0�f0BN�*�F��~�trx��<h6�H㫨fCf<m�A�9峉�e�;0G!�"Nl��6�S]�݃Z0�Yϝ���}]�|�&�'s�Ϩ�̟s���cg����Q��Z��:or]˱�`���=`�~WX�G��[p�.��*�k6#gU :MV��ftit��я�1#/U���et8�T����Z`��$��NH�Tk�
��h���8�욮����{��+�Fch6�|���؎�[�tn��oM]Un7n����G.�^_�eW�
�f��n:|z�GPc��F�껽��Lv R���z��(�c��mmuM�-��<��(�������W<��9i�W��u��q�s�{͛#X� �B�	��:1��*ƶ5���bv¶>�%栞�_n�{N��c
���a'>��7aU��VP{���g�����:�y��z��o,�='y��h��
��c���N�e�3fKFe�M�"Y�~�&�T�A�ǉ	~��ܲ�{�ܜ9녷h���b+����,���B�^]�픇W G�T�y.V�o����^3li�8D��Y�n��,���(%U=S6z�dT�K(_b��rK��Pmbp٪�Ǳl�W��i���3��qb~jѡ�Ua0z$c�TQꎦ����6�Y�zA��PyQۼ駉�p��PE�$��3���-d����df-�#`�"�s�-������eg�2�f~�ns�\�.�nux��
:ۄm��H�$��oJ�K����j�;���v���l��E�	C���p��R�݅���ER3�m����/���M��_v��c\��1�	q�,dd.�1��Ļ�~:�R�O��x���n��4n5�]>Y�4{`:p0�Vk݋*'-��m�:�`�'��Y7����[��a�lu��,���ю�����͛�µ�ۓ���s �I�+\���y�C˹ ��9$��/�re�����Ůe�b��W8����
[�z��{Z#87��v����{��\�+q����>��>�ڍ����r9�r�K+W�r��{��%/$I�U�l�+��`�l��������T���(��(�G�k�upllC�G�='Ru] �_�hu�G{���ʤR�Pɑ���ɂ,����gl�GR4��{Lb��]��:���!;)����`�"���L�	l�I�e���!��x��A��`��;V�Tك՜6����c�/�<*5x�p��e�{��O�"C�s�M�r�F�pnNֆ�-ݳ�lGP��ɴ�1���ڹ�����q��S��Z��X�mˊ�}ؚ%�2��X8�m��5�o#a�w ����Bf8�>�����@��'���Ȯ��7�[kPS�JԄ���@>Z��s;,�S�G7f\�<��oscbf؍FD{��uܒ�U���6K��|�p_�����������K=��3W'i�jVG>ʕ�r��3������ٸ؉��rK�Z�}jif�c����J�޼b��7H�aP���x��bQRZ��O��+��lu����1��8�U������d|�.��v�v�ZW���:N�kPA]n�iz�4��dRt��7�oy����ا��g�i#-�) �#@�J��I]����TC�3����2�0���h�c\Hd�7�>�G�0�����7a�\�y�~�b��y �%��my��[S�@l�u�����cxs(�b�Z�]#{\wTu��m�0�A�pS�'Vϯ:�D'�b* �K��2�f��n�z�� �:�$���B3����]�-�9���^���5�
���tGMߒ�yu%�8R|0N�k��Ɣ7�lO�A聴t��L9'v}%WL�����@�]@�jߺd\�)>�v;$Z��԰Ẓ7ĈyX�5�'ۜ}mFϹ���;^���t�?|��S�C�{힊o� ���ZHF��c,����݈�x�H
Y�oFjh�Һ+t�D�[���6��!݁
�z6=�_�E�7�-�??ڴ�r�].�t�Kd�ᕀ2rk�.Q�����x����%B���~��<U�*��W��&g|���){v����mG�fһ�8S�3{�v,t�!|�n&��E�8�XM٫ymЧ�Շ]ؕ@]=yj��yHR�ݚ&�f�gSl�t5-�,t�X�u���C8A��WH��aa�l噸3�V1�y�Xw�1�����h%hr-�t��w��C�
��/W>.�e�8�x�S�||�r��S��Y�)	h&�H�^?��?[ҴZ�vQ&)��ΡX�$.����½5����W�@�5��؜O<�.!dBu��y�7"P��3A��E0iWPx@ŪC�&#ͨL.��RŠ��qד_�}�[~��ݧ�z��o�[�9��n7�b鱅lFTEE	�}'p����9�x;\U* ����@�Zn�>i����Z�g&3������L����)+�\i�	�:��L\4ۯ ]�Awݫ7Jx��ͳ�o,N��`�t��<�T�4�Xo�>��Q��*�ů� �X�ݛ��xӾXI�]Fوe�D�'�&;��{�rב\���]���c����G["a�;�S/1���``�E�ԡ�m��/y�������G�,ʷcd��������M�T��D�ӂF�v�k�̪�˷Za!�	Kr�XA`9(p�W�H�H3N%���i��0%���X���a�����RiyG��\��7�'e�}�@#L��� �W}`T�B�i%֫LU��6Er���/��b���u��9Lg��f���
3���4��\�(�r�5���zܷ}�}ș^'�R���#h6��o���~�_Ym
<���ܭ�!a�ñ�����4���;�c�힐��G4�g.ڸk(T��z�{(���)g���J�^GނR��7�$��'�����d]�1�꺳�{+�vfnL�����z_j��r4�̲A�BDg��G,����b\6��沌��WO��͠��-@{�k�5u^��D��|A*P1�o�m�^�q�Brpwmu�>5G:�m�	C�OT͞�ȿ^��6���Y���m]�Q�_�E�*t�m����ߍ�,�A\X�߄Z�xL����2؛��B{6����C����u�{�s:%�M3�y9>>�,�P�ײn ����Cl6zNӃ6����VU����v���M�P5�)���`q�O ��z���Y�����>6��X�R�B ���c�
ݸ��Y�'u�<���-�=3֞h����)N�.��}�G��&W<�i5���е����;�5�{��:�s	�[�G�ݨo�#e�)�c�Z�hܷSٜ�m�F-�N��0��	��p���n�F�:I]�J�Xe���D�4���R�4co�w��7[	�J��h�t�D�f{��{�J����R@�U@�jN�Z�u�qxULuC�s��<ޘ#���!���{��X�U@tQ��^�Y��Y������ǌ���|���e�`�V�z6J��"
8���1��r�<m�ݱ��,ow(�[��`t�q����a���E��[�&�ʦ���nx�T��)YAv��8�R�����u7@�������Ve���9\�_��q�\Q�9m���H�	�s|�H���5~�b9�^�<(:W�<��Gg93��ˆ`��\hq�'ăr	�Q#�y�)���y�o�A-�V�w���s�F�g�+٭�'�u�v�����e�y`��һ_�zgYEr��q!���~q�Uv0o;�vn�R��[}�.,��~�FS�ZE��2\�ܭ���@j�Ԡ�*jj}����*��U�w+Z�jվP�5dc��N�d�b���3D�Y
��<��ޚ�k��1m@�"U]#�c�C7��;k��DsyhX���Q�y~�|�1B�=%1� ���ݰqK�hR��^v�����OK�k��i��DH�ɦ���S��=�t��b��0��m����5@�ɮ�v˞>Ί��-�uJ�[Mז��.���R<��U��9=1͹S�Gl���]B��Q�ڂ�K���P{%m��Ӓ�V)�4%�![��W1a�nz�ӪH�غ[�Rz�O%P����
�M}=]��n�Sd4��$�����u�|s�RE�!4��á���Z�$�E͟��>�K]9�gT:+k��@�e<y�f�>��d�3���c����I��x��&|�vGu���o�B�>��z���\���SX��03����7�Uq����3������Cۘ�O:�..�`++�sȾ��G���4q<�wd��,7���r�M�v�9m%���Ā5g,]�ڲ6�1��[:�7����O#ء��6��J�5�C@�\��ʶ�+hY W��=.��λ�''�%oĕD���
�M� nq�f⾉�׮xr��YxYX�~t�^b�jc�Ղ���P�Y�[����o��{���]2����o��F��QAWL��6��/:�߫6+	����u�bA(g��m��@�����~ֵ_�v�&{V�:n�ř��g��n���f��Hv"�f�c,�o��G���R��8�I����T�P̔�gô_H���gw@��y�Y��KCɌO�Ѹg]l���7�*z�����Ōi��ob���!��B;����g٦�r�����k�^�X��|�ߨG��V��-t���rX�T�������yo��yQ����NUnD(X7"�$7� �J�Gsm	�����M�z���Z�P�zY�+����&aZU���!f��(L�\λ/���-ß2�G����f\K���*�B:�A� j�ֶ=�}@��ۗ���J������'l�OOW��fA۹�n�U��1P��n�/{~�>ޟ�}�=======?�Ƿ�˟/����툀Ҫu��5�6fx�ꇋ�}˨�c)�����ʇ���=ک��Oo`Zأ��S�{7ywD���b�G��f:���͝O��oAFv7����;/s��[ �o$撕>�l^-�2!��}lA����)��Εfln�Ѫ�`���F�*�����}��Wf]�@�v�^!Nōf���o����b1YO<o�<w薗����[$VC&g[������ĝn�P��m��R2����t�#n���vm�|jc:P�L��ɫ(��Ɗb�Wn�B��-�Mt(W���_�x��=��so>�0�U�2�h�d��� �����s��F�r�"���b���Uu �V��/��5�$��ȫչ����T
���KUe>�H�K�U��5kY���6����� Ls�Ð��ks䎅O��c1��bW��k�b�z ���&�y�斺��a�5c�͛0;�
b��L�Ԡ����grͷ���n�Ѻ�TO1��ʐ\QC����y���۔�Z*ݺ+)l��嚶x�SF*UH�n�]�7�c6����cu����u��ܣ2�6R��F��|ܒ��85,E���vP�Z:�u~����x��$�-��*�������}Z�k,^L�t����8��K�⾞��+E�) ���eDr#�y�<��H�}����擽k����":��kZ���k]�:�t慷��t5#��M�fp�.�(*6�ʃ�F&ЎX�Y4���m���[������Gn�k��1�ڶ�k%�u,������.�޲�U�Y��du�#��9�{���{D�f:xL�
kAg���S]��mU�XcBU���Lq�k70�|+vTcj�v�����#��d&��urD%d�īk��e[yxmF�Vv�<\Y"��ñq���\ÈR�+(�9���:q�*$�oa�Р1�x�!8Si�H�n�g'Q�lк��[7]!�Z��ys�*��jEU�"���u�l��߮���&a.8� �(3���9u�����[�D �w�����P�B�Z.���V�sC��ѓ�ڲT=�d����������P�K�|�I�w��.�pU�L��]&����SΔóR��53@�gW�-5���]{S��ǝ���;�9���K��lR�w󧦎�44���Vv!\�Du��r���[u�9�WnZ��B�f�o(��Jg�@�ժ�A�_��;H��cR����|he�r�%�k^��G
K�<�����u�@{!������OQ�\��cb�ݹ�*�pm(h�=*-�p���Z�Vw�'���xk �G�WG�t�˳�P,v�k��[�{�,֦��1j��w�
]d�s���p��\0³�9I-��+v�p*BM�dY�g��G�ÔP4���+������YRι���6�E��2��"�qH�âA�^�pP-%R����i&�)�bF������������6�R�l�RR��M	�SґLEP��QCE4SJ�I�t�P]eւ��F��CC��4�f"�8s�j!��m�5m��Eh��:(
6ԑ���ִ1c�S����S͐����I��Dˢ���rxTN��f��hj$�
JJZ�6�shj�*�����
�4Z��������A��*��J��PT�kTӤu��i�)4�hJ9&!^?dZ��
�ۛ�i�p��_+�j��m�ɛ�P+�ns��ԩ����˾Q��Rnd��/��yM����Bvg{s��%���wo��OҸ�����]^���\b�UK� 5�_�C㈼dWax�R�uƃl�:��'Ԑ�� �C��:��~.n���GxG�6Ў6�m<m���ZW � ��:���y���r�n�c�6��C��Dl������5�^y#	.�5v�7�U�^N��xvf��!{����ͤj�0Ώ9� FΪ�4K��җfݽ��s��Mo�a�7�3���R��C6XVy�͏!�ސ�
Td��*2:fh���RN�v��ݨ�s��W/�������|�� �?b=C1��Y9�&��ub��k7�<kL��2;	��x��&:A�=!�����B�W����\O�~�ğ��{ÕOk���Z����r̃��w���Ic�M���R�N�XV,Q���(�2R��ي���L�գ`n�̲A�D���<�{|�L�����\qg�$�V���+yM��3�8�����ת��v;Ua���WG����o+~_����"�1%�Ф��~�FӴ�>p�9�+3.���{�2	�r�Q��O���F+Y�v��k{1�Im�/0Yt�C<@��'5��"]ѥ.r���W�ztX�(��8"j�2=h���m9���P�ȓoե�q�8"���3���J<�S�&l��N	x�p�����͞�#	4T�	c�u�Fp����D��e����U��r3CnU'�)�
�d�5�W��OM<zi���)��P��]u9�8�+ǁf0��+{F���h$T����jw-Չ�!�h��[=��O�g$�Ȅm����
Qs����T���n��M�]�V�캸���u#��!�.�#b�+��xrUx��1|Coa;��gSg8���h���S��q�ƽ�]!��	�G�+d9τou��:uZ����t��N�=�}��}��E�LGI���R0p7 0�'�1�Uu%"*��jٻk����p��O+]�
��
�K�`���6���OsA%��%�S�S���cWLS��,��Jmv:�yP��J�,%y��Um/�����^�׹�k6.����c�kkǁJS
s(_]�Bѩ˨�Xf���d������Y�ړP�݆4���CX�ȥ�;���<��v2�[N�#ωG���o�rgu����"�@]��NM��Ǹ�7�ᝮ����B����=ԯʺ ;Cz[��|���8t�y�5�L>H����^C�a��/�H�5C�r���Ç����e���n*�v�p�@����9@x�� ���KI�$H$�1SSP�oT�mΐ����=vz�t��
㫡�<-ylLѨ��{�]�sm/��z���n��x���aZ3�z��;l�@�x!f<�����3��y�#�k6����a�����滸�#�M ^Z�tSǵ��wPA l4���Fw/7faN�ep	���\T��KlAM+S���x\ә�i�C�]��D�l��w����q^�N2�?��*�ޏv����U�ʯB9>;wy[=i=dݜ�=�	gH�?q�ɹH�j��غ[�R�	�O%����d5DT�o��Վ��^|��6��5@VQ��R:Y�m�'���O��W�4�44�`{3ٲ��M���I~��jb=ї嵾5�e�ۓ�+#�s������tY�27�Z�#�J�v�y�]x��V�ܱ�f�ɝVÔ����̢�V��$�6���ݏG<�FJ�-b�*Mx8��<rۚ_�{f������Ȼn��zv|�A�
V��u�l�L�:�Rj{��g�\�rx�*E[t������|��aN���7�Y4�JP��᱅��R�2��Yz���[�Q�(8`�`\�auP��0�Q���7���;@���ޭ�]ڲtQ��,/$������m�t�Ai��B�qm����bD�0���l�腝f�<�QD�)������\�I�7].4�'��#��qa�؍m���R�g�eEV�nU;��Y*�(���<����߽��k&Շu�ϣ��FlȌn�������ɡ��K��#�����Jz���ǵtߧS>�!݁xVu4L3;Ʌ���.-�3נ����ĉ��O7X���9�A���l!gk���h�Na<�"��ZT!^R���� ���&��$�M�7�vi���v�g�ׇʹs�}KT��u6��3�����Ra{�|�LCgg\\�u�9��F��h�k��d7&Q���d��=dI4���>!��)�ci�0���⫄�F����=3�n�Ҟ[��]31��%m����p�WE&�qJ	o5�Bx�o��Qu/�.��[GS����x̆��&t��{����޴�%��F�����3��]����{1hU1�iń���Փ�q����	A5o�}���y����$���t�����
�P��xF�L-j��]��OU�F���y�RC���z��)L��ﺝ`l��]91~Eduis�V[�7S^'쨌��-��*����5���%�P~��uz\@"�0��`�vj�"�wW� ��`m2��災)+�:�#g��uuf@l����L�͑�}��ל�#E���n��T׉��^�lyg>hؾ��l��:n:�vOk]T�[o�|4-�CzDl����f�kϫ�Pq�K�B�W'�VoM�_g+t5�>[\x!���*㧺�M0r��̝���y�^�-�;��'�w`�P��M�o�F����wm��ukk3fNJ���{fm�/%��L���	C9*ڹ�˾��@ϐ�V��@a)�C�l�*NK3�%�4�� ��ŶKӺݖQ���e3�I�Y��M�I݀��v�K��'�ё�ܐ&ִc��n��[��WӁ&�WN.�z�������dZ^��.��U�7t���.���mq�3�;(d�P���}s�W�,R�qL㟒1l��D_e��Q���n�D���\X�c���W�~FQ}Юw�"�~i�V�g�`���?Q�r��9d�G��A��E���iN(fV'ٽ��̅=�uCl;
7�FDy�ٴsfYx��K�s�q��7v�]����C�dhn�fC�i�p�������#�Hc�^�H��T��5��0Zk�� VQ�V�}��`���S�z_���)�SC�#&����6p�����"�h�T���ׁ싉s;��+��,C�DfMӋ�r�B��x���P"�J�����׉�#@�I�A�T�OM<M6�j/�˹rr���S����#f
�DV���R7���x%����T�Lo32���"&���p���(�n9!nB�n��ow{v7ΑW�*���t�.�ݠ��m�6�>P�ͮ���O��Mk����(���M����� �e��filnI ʽnu7F�##/���)���:ϒ53i��j���H˩�g��{%��U �&1iV��O�b�OF>���"j�2P�{0����w���â(]-�3{��=�⸵�G�=C�q��WH�#v�+�/�Jum�㑆~�������s�<�):_d����?���Pf�D�κ�Y��.����ѧ���ݍݩEER��%� �:�7=��d>��p���bf%��)�	�>٣=�����]�(*�W����[3J��ك�tE�{�ʶ����{'Ѩ��+����f��j���n�����o�V�����g5C������xH�Oӕ�2{�eTU��L,����h��R��Y��=���0<�Ւ��2��\d�t۩�dW �\Dwl����=22�l�2:�Ƌ0�V#���!ZNr"�[��S�d9�s�_�Oޭ��ǎ�և���!e�)aa|.rŜ�m�/6�gb��Cо;(���^R�tS��P�<x4��n�y��]f0�~b{:V���9U�]\ݩ��%�m�f+G{��'a�����i���,Z���ͼǴ{DL�ϑ��p5��}YW�e�n�c��锇l�E ޥW[ڐ�7ہVd�-����e^�}��M���sט�ӥ1�J1��:u{�GJ����H�*{��|��k��kϛs���-���/�2ї�R��}��p����K�dG�HW]�%�B9s�w�Y�k���y��l�ȓ�u5l��ɹtF�'͠� �Xz�3��cսXd��j��[�A��v���<{`Q BQ�#o�v����Kp�z���ƱK7�nM����w�ejt�}���ڞp5vFL.�[89�9C崟_�O����QH�2n�W١�8A�<el����=X!�.�Fo[W�&�j��J8�A��#���	�?j3����Y�L9M�zn35��Xw� b�BϤFɪ��Gs�յR�'��j��i� U��{��\@v���ί_(����m�L��j�:eH��'�� �j:Gd�Sc�D���=��F̋�����/�+�e�"�ۛ}(����U�g���T�D���t�c嘵 "��]r<�pZ��WŖ�O_l�<#��;Ż�1]Յ�`{$����ö17qӾ]�}]}՗��kV�G�`�m�M�_]	*m���.i��U���F.{]����{PJ�^c<��N�D���|5��[? C(��L���	GH;b:Cln}�B0��a�j�y���s�}���Z�����o���p�����!��]���$�v3ߵ��m�7�H��iR�V�O'�y��b��d6��9LC�'��7�L���c.�^���c��wD<�v�4��<�U�����w7l�1}4]ݻl�ln��z-�6\��� ����xx�����Hu�tiU5�Z�n:�(�C��]���1ez��G4��X��XFC��TM����u�v^RW�꾻�8H�4_�E�z2x�*�1��9�PAO��+!��/�߁����?�N�+Lt7�0y��FUn�u"����9q�w/1�/:vP�uH^�p�ҏ3�$��+H�����S��N�*'��h���8a<���]#s�7��|�6�O���&���g�Ӧ�'�y�Pq���������$C? ӵ9ua�&��*�/_q��Q�H��y�W	C|�Wp8�v+[��IKGDQ��z2�#xmuN��<i<�����Y�M�B.�l�������(_b <�,s"���]b\�&��T�6��oL<�t��d�0op�p�m<�J��x�\�2ޑ���%�VUר��3P�v�H��-�Aly�ޘ����W_�T�\�7WPۏ�S3���n�����(R*Wc�vmt����ȍ�]J[�
�[Oh��]���|;�/�yx�n�2�ʨd�i�z͏�pQSY���뚷��b�7<t����<�w����U��ch6���%�}m٧Z�,#&�vo\��.�e-��ش�=��c�YL�R��v̎�Ǒ���fNf3��ǆ5��~��%#�:�2_Df����=f=�Ɂ�Y�Ej��/7�#��c�(����*����2�sǽ1oB�ͽ�g�X��P<u�b�U�u>�7���bq�E�no3;�;�QQ:&_ZlKڨ�Ge�k����h�:nL�86�x,Û6Lh���.��K6d&B@K�� �"���/�/�H���p��#�N�x����L�+0,����0,ʳ"�+!
�0,�3̣2,ȳ
�!̋0,�3(�+2��3"�2,�3"�0,ʳ"̣2,��,��̋2�ʳ(̀L2��2,��� L2,���L�0�ȳ̣2,ȳ̣2�L�2���"�2���*̋2�32�ȳ*�00,�3"̋0�10,ȳ̫2�³
̫0,Ⱦ���>S� (� L�0,��*̋2�Ȱ�0,����@��C(�U�

��
���(ȈȠ ʠȀʪ� �s9냅@!� !�( a�U� �UV @UXy.  �@ �UVUX` a a eUa�U�UV�� ` eUa�U�D�  aE�``Xy�dY�fU�FdY�	�f�O 	�f�V`Y�	�f�`Xt�Y�fU�VeY�f�V`Y��G����z��� i@D� &O����ߗ׿��A�\�s?GKGՎ���Bg[1���u��|2�����@_��/�?�xUO� 
���!���@�O⟾_�O����hP( ����;���G]��Ȟ������7�����b��~�"���
"4��Ġ!���*J�
K A�A
 @H�� �*�2�� J*Ȅ � �*�)  Bʪ�� ��� 
�, # A*�0���* #��a�����?$�آ(�@�� �
�#��`s�����O�_����{�h������N�<���
D�QՈ$ *�ȇ�O������O� ��
 *��~D=�>A��pET���<�dW� 3�?�0�����`��������|{| ��PVX��a�fo�$ $��dn����p����<|�? ��>�O����8{� *��c�?���
��<y�􇐤�U���? ,��p9�g@��i��I��y |�������T��x������k���v��PW�>�>� *��9{d}�������1AY&SY�e���ـpP��3'� bB~|�䀡$U�ik)
�B
�)T�)�Tm�R���@$�ђQhj����*R������IUUAiX�T������B���Me���]��m���Sj�-[*����^ͪ�P�j����I�U�{��ke��aa-�6ڔ(lm�%6��Q���f���F@���Md`�e���Z�jͭm���)C3m�6نZ�fi�+��3[fH�j��6L�3V�4D�2[Y�M�������F�X�6Q��iv�I����  ,���ګ�;v�p�4v�k�Fz�:kn�^�w8v][m�=o^�wN���^�۲����P�ov��l׻t���/�z���jv˲{��h#zolڷ������U[���[U��m�S6d֝w3�  �s�СB�
�l[�>��L��cKar������r:6���lkKcl��z�䮗Z+V��W]�OMS��9Δ=7a�x��v�J�������v���v�x��+��ܯz�ʭM�U�ضmL�F��m�   �u��F���m��Y�ڽ4�mׇ��;ݚ��Ւ��u��{�Ou�].�{R�W��wJ�vݽκ�v�b��ޛm��w[g�r7m1髮�n��m�9N�n��6�;�mm���MTت)�T�[�  �zj�^�U���ε2�:kv�0{wmUov�y���Sf�7���{������;۩ͷ�����ۛ��@u�
3���顧�V���mm��bfj�   ]�Ѣ�t黶�8���v�V*�t�Xu�e];.n5B�i��;�E��Q��]9p�\��*���Uf�-XڭUf����  ���C���x������ s]u�@�[�*�+mܻ]T6�ZgDg8ŭ۝ ��56���k��X����j�V���J�ͯ� ��֨�|�{�Ui��t�WGUөܺ�7s���7������v���@�v�  {ޏt@��p  6�EZ���ɒЪԫ6��>  #�  ��C��^�  �� ��j� =�y΀� 9�  5�q��  ��z:  �
�Voe6*ڌ�eR����;���  0� =}�j�t�ݠ;�  jc�� v���A�is�  � �` )����x  孍�Te�m�m�ԭm��  �{�  �2��К� OsÀ���� ���  ������h4��  {��^� �)���R4#MhE=�LR�� �a "��IJ� 24 E?i)U?T   i��R�4�@ 	=R�&eU  ������~���M7T5��]{
�����58��ң�L��N��ix�iܼ���! @���������m��m�mm������V����m�[o�[m�[e������������_��;�K"N�b	�;[r�mX���Sl��Šv�++�oSx�Em��� uZiT3���\(e����8v�n��5�cQ7���T��1n�z�mf<��c��oBa��Æ�ю���]j{�k�SZ/.E{�ڍm��{��kV[�)*h��7�&]�EH�kP�Ph�X�|�M�t�!M�I�V7]9?0f��ew�P*��-.��y�����n�-�eZ���{j� 䙧U�&]EF�;�+O��`Uͫ�佂�LȤ��CGF	cN�x�<�x�H�����X�S�u3,<�k�]޸s��-j���|.�ŒŶ�֌Hn)
S_Z�Yg,ӭ:�yZE��-t*�p	j��jΑd֞]3W�\
�4]gpCK2�D�m�h�j�t�%5����8w�fU�r1V�[���dİ�Oh�(�������t4�)�L՝�obm[�����Փv� �^D�W��Q��w�h�-��jfP�7K��0�$ti��j{k$���/��G�w �(��߄�.�!(^n���nVm��J��ҏo�E���a��Pf诖b�r*�MK�)�Ũq{�5� hi��Ĺue�r�`�i�b3֍$Ȫ�'ѻ̠��H��#�p�m[I�*�T�n.��'j���B���!&���1؄��Xu����0�2]��H�V�Hi�621�vv��;
��X��p���fܙv�i�к��Jܠ\֕6u�˻T�Ė �Υ��muvV��ZT�ma۸p=�'n��S�*0*��W&�ݹ����p�	O�B�e��͏8X�v���YZh�i%R'tr�:�tiג�1kuc6^�1yl�tS�x�VU��N�'ol2����DT���"@�hNf�-ֹ1+��ٽ�d8/o�v���-�#0D`��a����ڣ�O3�^�w%\i���/X��m`J�Ԧ��M��W�
��з@eMM
�Q�pccE�ةb�-��6��.��n�i,�Vs,A��L�-�Em-��N�`�4���!�8�ZZq�CKi�����$J�bWu���t�CO�A��$�e����٣@�n���	Z09d����*^H>�ֽ́�d<:Ue �9!�J��p<
4���SATvS�:>���CX�I�m�!�q�(��1�KM�U�.�8ӍU�N��#b�j�@�v��*�C�nCy�6l�ñ6RHi��Z /C;C\����(�b�I�X�t	ڛ���Cڲ٩�,]� TQ"[4>�6��zֽݨ�E��7r���	Sr���yY�[���37-*��̈́	fD)fc�Z�yl���J��GLX�'�^�����ؚ����#����r�nIZ�4����i�8��4��+F���J�૗2�lv�U�5�`7�	�AV+#�'f�ث�E�ZĦڊt��^���.nGZn��
K
V�j���"�,-��J]�{qXf�]�MKQ�bܰ��?f�sM�p���B�F=����bͭA,�ՑF�T����Y��x��
���wr��Ŵ�ør�aB�u�&�͙�� ���Ei!YD�����y �w	k�B�b�+x���sF^��A�b� h;�'k7*V!˕���|7��Zę�\*Ⱥ�iԘj5�Y��'.�1������fE`���Kt֢kR��(dv�(]��+��`�Vɚhb�T��u�T;�r��5Lʶ� ��Z����{yY�˨.��b�f9l��d:�YJ��C,]9f���1hf��\h̦��n;Œ��*���lP�ć]*J���M��m+��)Q�Ŋ���u��P��D+�xU$��am�m�De��AՍ��X�]��5��`ǩ�Ӯ�$n�8�SM-�`Ȟ��z����7h��NV2*�lPB�	�[�;gwҌ��Iy�,�W��,����X��+P�1�R�CG�3�+(�z�^�3+P[�Z�=�&�$6�V���b��S��V�n:Zɓo)Hm^�V�̠A� �9�u�3.#դ�a<�t�ЗfYޛdc���O���*�E&��[�B���Pu�+E[�"��f�sJY-e/�I$)�Nҁ7/q*{���*�h����Ez�g�hݲ�PoEj��a���sv� ǙJ�3U�hG�]�*�$0�u*�����ܭ��PZ�6� ���J�H�J6�	i�l���'Ijʏ�fֱ)=�e��n��ۭzt��`�,�U�^���XhkVGF�[�N��4�����*��u�Ɖ	in�Ur6���䛕�KJ	��#����Fn@[QC�k�u�=rӛ��PQ�;db�T������	��0��u����n
�r�"ސ�"
�
R��R0:/p�k0K8�Yp�ZU�I�pA��ٸ�xN���[y­��ۺ�kL����b�h�,��j�h��֭�jn�e�B��6i�V��*�6|qӢ�i�K6�wR�`�Z��.γR�!�Vh�GJ�MGv�k�-'F�Hm�T;{�3!�/s�v��f��p8"�sU+v�4��Gz
j�N�.��,�f
�P24V�iMV��E	�-��tL� km���$����+c��ڌ�J����U��������k*���g.^�j�*I�V]&'F��*���μʐ�����5��AD�[g1�7�yFF���8F�T54
wpM�ze���9cJ����R��6զ��ԭ���K�BR���r ��Av!�j��as�b(5b�r���ژ�Q$p-&b��`� �U�-R�L��4��/��R��fd65�4g�sfe\f�RH��m��J[�OKB�Z!�Y(*v+b[�bwkU����%�m�R{`���Ul��N6M��Nݥ���T�t��QQ�4�45�X���CLT��2$�EԻ�h����4]�uV��e�$3h*KL�c0�hn�N����8��I)͢�-��9V�ǌ嵖�cs��XjLU�������M�m�ሌ�{��]G4m�ȵr��؎0qQ+�+�Z,�cofdU{�Ұ�6���ȡ
�f�;N���)�Ũ��T��&�M�^��[�K[�4R�b�����֝d����j\�k2�-ҘUӨv���ii��4^��V)�PN��iYI�84T�N�/o[�����[�s5rn�I���*_;{�3.���wN���YR�W��{D�E�m�֢wqdM,�@�4┳qnfi��M�(����zX��/�㵉��B1d���w�� ݹQ�Bf�
�o"�X�l��
�wW-dH�[�Vsp�G-#���e#{F���c���Gi
��@�7x`;k[�Vn�O\��'wvPڕn�<���F�dP��.�K�T�@U�%�L��ҡ�����9h�.�H~�#�L'3!��6����n ���s�uØP	kM��5���)(�������dm�h�B�8�Ռ�r	�֋r`����b{���j��A�(�i���O�VkOu�b$�5�mB�٦�]��V��v@�GU2 코fڧV�m�p�T@y4Y9��OF���]-��t��}��ҫ*�miv�b:P���VȭϰȎ��,fͼ�	��ܭ����d�e�����030x3XX�]���vhda!�mk��Z$��\f�)f2Û�^����ٻn���N�/),��B��M�x�l��Q�lܽ��BY;�JSi1[�V�QM`;r�����U`�q]�v ��z2����#V0��Lwz	��"��VSݐ�iӼ%l)X <�U�X�a��s׏�4�*"�x#�h:����\@��,;���:ġ�:L|(۽n������*��M�xr���H�u(2��,h����2�29*�f�E��:�v�?A���%n�(N�$�(�������Sp6�ٷ�]��ٴ�r�%[��RŦ�3�hV^��ˌ��n��z/-Qݠ4��-m�F�:NhW��dl�8���	�n�l.g,V�w��@ d;Y �nRY
ulla��8R[�~�9�ҡz��S���(�PXu�̖%:	'{5
 ɖPx�b٣i��HN��uVE��a0�v"))ui����T
��@�9a�u���I-��������-�w�QŚ �R��EI6V�D�A��Ȍ���f�w.�87XY��t�:���
�b�[�}�k�.X���*zv�x��X��Mɨe`��O]ݐ��A[OB)]��Pt.U�`�F9H'��kw�$ѭ��[Ɂ20 J�p	G.k�
���my��`�7�!+ �B�]��6Q��g�ڭ�j�
uu�puh�)D���Ad4*L�dClVMCZU�"�v���� ��RCn��&��2c3n7u���ՙ(�f�P�������Iy�!�ӎ��N�D��k��&&V��<W��(كQ���˥��Ż�IK*,���J��(H���O^�R����i���1B����z����@�n��3�cIR�
��2�59.�����<ͅՋ�FW.�M� /eV��`�vd�z֊�б̟h��.�Y�1$^^��Nd�oC
^'pU�&v-
!�U�x�d�)���V���ۼ'0���V�fb�l4l[�8i☤˘۹�W�vYpS����B���9;SE�l=��t�r�����l�栦(�#a�5����4��I��(�-���YU����d�M�汔-R�V-�)A^�c��hb�Ne�f�b<��s�hz/m��3!a
�Σ�w"���-@l��q����.�2���<jyc0&�֜��^�Q�eJ�Ȣ&R��E�Wj�$��2�h�%��j�,�����ٍ8�h�����qPv���DC@�KD�1����`�YWH�Vf��K��H�7��α!�U�x���Z�3W��J��v��`D��j���D/1T�ct63FJ�l��ā��լe���j*�0��c'q��.5Ho\j�t6��%���2��vshX�^Q��JS>^$�bQ��i��źH�83=u0ե���LeGN�����f��b.��kY�OS�-ئc��E-�LK`�m$���n�v�ʻV0(����Xċ�F`�APe�j�%)�ٺ�ϊ�2^��i�ߓɲ�i��PR5
��ȨbB�n���z�8�����;�*Z� =yve�V.=��62�اCC�KEa˰w��k[e�ٶC�q(�9��k�*醡.ҢU���7ᡄ�����-&��S��EXu���i7A��2V�Ee�!����c6����]�n𕶯 ����*���[E���X�5�>vT�w9�ͬ����2��ƥ&��ɇU-��h�1F�Pj�6�j���q���(Z30���ݕb��%�Ҏ��EK��f�/+5���$�[�2����[�&�.EE��Ky԰�̊╗Vh"-)Y�����)�n��čMuˎ�k^!fEW��Jͫ��A���0Łe<�L���EU�A���
��^Y�w��X���m3�Xٷ�����#rާLGͥnL�E�V�v��X��5�gX��w�i&U�mF
&m6��oEj&�Tt�@���fkV�yI��~*�]�N�V�e�2��nc�ѱ�&[еT:�;�LM�������@w1�b0 FVQb�e�J�9�;�/�[����I���~�Xw2�(�TL��zH�nj�ͨu��{�Ȗ�O�5�Qn�鸤2��j��ը��q+�������x)i���p9)�+V�5�����2Eef�Z�ţ�Q��H�̙p,���vu� �z���pRG&�����@�La�),�{�w�eǒ��KX8�J9��V��*����%��2�dՙ��Z��fܲ#�w�h���Ű�u�%x�q-{dD��WoRF�P��Oj�[���[y7�n�8����8�,c�pO��[�n]b�5�"q�)�M+o7$�YF̻�*k��t����P��m3m�j�gpb���"WE���N&��<��֞�b��*�&朕�i9F���z�-��.��k5f���Z*h�7���l�j��R	*!�gsJ�+X�v�^U�+]Z-�)����ыAW�adӗr$�]֧ŵjo2��L[�[�6�m
Эm�/K�,�:У�CDԻ�Ň`WZQ��K��Y��m�%�T�5����æ�Tچl�7���S�Q�j�Qyy��L� n�%9mbhM���ƈ֩�CjbN�qc��<	�X��ڙI;3^�K,�p��҈R-Gl�xF�퉧f@Ӡ�6��Z{c7�������zI��:���
����/2�X!
`MnS�oV�Lw��CH'�0:�E�T�K��T�x��͈҉�nR���*��w���^�D�di��Z	���Qe+I�HJ��˨�(01����7-�V�۫��2R3�:�[��M�(�ս1����d,�2�͛-�Tt'f�f��*!�T�lܛb�{X�54j�W.�ǹ�a�F��d/��j T�(���FZՊ�x��pT����(�n�A���Cx��s2�$�����eiTu�Zj�+�ն�7a"ތĤ�^ 'ȡ�iGm<��AO@jɷ�mVC@�"�Cb����+��jݑ�j�Jӡ�"�� ��5����3�F�tʔѹ��r� DdR�f�6� �s&�a#%��rse���/t��}DEK@�Ȩ�E�I
��Am�����Zd���H��׺�(姵��Sf�t���ޣ�n�9���%T�&j�=5��	�*s����J�+�0������|�:�vhU��ds����[WJ�:�Ъ�U�ӈud��+�е�q��z��ru�a�KՎ��T7��C��&>�͝y�S��Q�M��K/��������8�6��h�R�WW�}:��c2�4�Z�
0�}e���ǝ�,n;��Qj,5:>���i��<��՝u�\peb�xًvFh�%��:#�U)�]����Z�[���m��$z� �aL�W�vt���L4�3I��z��f.���,| �^�i<p�;z���i������gU�������a�X�tZx�{+)��\�n$�i/����F�"�����]��J��C�Ӕ�u�E���n�e�fQ�%���Ԝ̭�ҠpmY�5��[���#%g10svrGyKY]{��-i����F��c�T4�UiK�����]8
��krl���2'u���0�H�P�ѓOg|�����F���.�oa$;�I`�N���KA))���4��m&҂%�[�:�YtA*]N����#hL����o[���E�t���3��T�Jř`(��V��l(Ng������wӷ��Z��{kY��O�'U����!Y5�X���2�ĻUrs��Y�{z~�s-�}�;���t���v�p,J�����f�܍Ҡ�-.X��|Q���\h8*��N����u�^�t����5��\��:2ѷ] �]ʺi�]3��n�T��ث�L��rj��3e�o39k�Լ����>JV;OzJ�8�<���Ӗn��x�̜=�n�=��O=B=}��t=󕂆]dIc�y��e�� ��5Jwz�[�R�Ʀ>��v9Mֈp�9�t���U���Y����b��u7��)irXɾ,�ü�p-�&��zy)b����=�]�45Q�FF�[\����]��ք�ͤ�����\��;�ח���k\�WS8.�7ev��n\Cث�r��(qu/�hCX�0���{��&�q�n����|d}��ҭJ�=�$�qn\�"c��(u�E�~2�uG*���5vW\��[J��v&���o��n����.H�t0 ۳6�l�ժ���\�|a^����i�v��q�j�'QJhu��-����W�*�GMd���냆�u=M6I����\%]N�����=��[y@�;�٭��l�M�GJט�h�М� ���H7�|z=~8������G&�R}t��9}���E����ן��୘|T��,���9��vэ��=�b����o�j��T{�YZ�&6i5r^Y����
w�^5b�i��]�Wyɸ�Y�&���$�Y�\��&ܤ�!�����d&�>O%g��ng3O)���T�[!�#����Q����[T�_Jx��(��αS��w�p$�����v�C��nd�a��u#\���Y_ss!�oR���%X�jHh
S�5�����Ֆ�]�WN�Α�W������%34v���7I�znu�Ϲ9��۫�e��]������m�s��d�c�o�5�c���Hu^|`)ݸ��f�ae�d|�J���'>l�U����؝�7RMO<}���;+�C��[::�Ec��h6����j�Yz���;�v{9�L(��f� �e��{%�c���x�T�ϯ.�B>yc��Ӗ��F�a��>ƈu�2{q.���"M���e���V�q���]��Ft��}̃f˨e��]���>�$}�+��Q��ߕ�c%���7�%�vX��F�ug��h;b�{'q�9v��7g)�ٙ�y�s��m�!�-TW:tXz͔Bz��핌��fAAxF�Չ
���`1�Q.��ͱ��tN:���)�^���B��Z����R�h��?Ge>�H�*�c�s5b*d��g
A�|��&C�n��z�2��`[�񍏮����K�;�H�V޲�p�.�u�Ň��MY�ݤV�(�S�d�h:�i*D;����F�ĺ�0��x{���V�_E%�vd��/�^gLJ����b4Ɯw�a2Ռ �q�Ih]����k�5Wu��A�a�s�n_}����TBV2S�۔�Vԕ�6]b$lFb�4ۉ��F��K�:��j � ���JZ$�����Eq:ί�� ���k�yjw˅3%иk��"��}���T��:g4Җ��e���k*�Ii�K���^M��=��U��B��+����"���b�:6�����N-<��o
�
�ϝ�e=��u�tYnd���óx�.�R�|��=s�A����y	����k�m��{���m'H�@�S]*tFr���3\N�LL�,��[��75��[G4�S��2m]���j���%`@H����U�CC�v�į���DK�4|Բ�Ӯ�À#��}7c���g8�R�rC���Z]b!�����#�Ve���1t����F[���-��j4���3V�u�u)�E��éTW�uΚb=׸!8��xn�Uw:�Kj�;i�[w�<Y�)䛔�5Ñ��(0ft��J��,�y�q�gsN]`��E�a�&љ��ݬ�|uu,�?���X�z����WT�����nvI]Kw�6Ob��鄻�ƍ*]�	Sp�'NҨ)I�e���\�Y��[|��v�3���b��U*�"���E�u{���X��\�u	��h:G��sӴ��;d<nY7�뷮�=��0B2M+nKA`���C�\c1�n��*T:�r�3��L%=�vIY;%��"�׺�FGk�]�3E��ܱ5M���w7],��ƈ�qfc��N`�ʾ�:]Dr�d��#���ͭx�8���P��qH츰#�`��\���z��= �Q�/�+��M�"���޹�Ex�J������F����f�;�b�{�j�]M{��%�������I�A�|���{�)e�(k���u��i:®qF�$I��.�`���ʸf� �d�7}͒��]���f��D���J;4�"'a�&/�+�bq��C�^��ki�8��Y�\�ޜڐh.�Ն�^��N�]��Ҏ륦��S*C�W|`-��m8�qlt�4n[�S�_c�9I��n t�����D���~b��Z���26��AY���}���fǷ����滰��E�M���a
��$ۚ9���[N
a�n�P�ޱrh32�E9�ރ!��Nl��X��㳤��F�fͱq.��һ3xΡ|�L�l��8������tx��q�뤸i��􉱀���^�0�_Y�K
�/�9��j�>z�Sc����9\��.�r�x>�M�q���m�\x	�9U�B��<|8�a�ܡS]s��4���;��Le���95X�%�Ը0�t]��_n�4�A���d�������Ԏ093��B�r����Opo^���{cQ�*�<*�Aȫ{�,�8����"�OdD;�$Ѵ���z�7b�C8՚ba�AE)����LHf[1vI�o8V&�){��v�h���v�[���F^�'K�wA�x��ա�h�K���Z�l�l�)v�E�ڮ�:Od+r�v��$Ub=<;9� �����Y%U��{o�NJ}���iR��mY$�9"k�y`�)�ޤ0��N�vI�4v��vt+Kq��Ԭ�}��FRf�H}��㠇��׫��Ӵ���U�%��xܯ�f���BY��v��,g�H�Tr�r�ƋX�F눦�ٲ���U�5*��KKy*�+E�D�*Wn6v��/w�Ȱ2@8��e��r�vh�FgŌ�i֞F�Z�lc����rܩ�C!�}�s`�1wj y���1�;�y�C���{1v̫@n�6�R���7ut���BR���Z��̽r�^wYIX��l�T5)�;�`��Rp}�/���x���PK�.jqɵ>�FR��&-dh�eLFh긖�\�J"[����,�u)��z1q�pu3�:��񙺊S��m����$ut5znW[%��|�Y�/ytʽ/�Z���Z��j"v3z��7T˱d�6&%J�oEnn^���	�^���{vf���o�e�w��� ��nM����I�R�Wy�鏉������!tzP̳�����.�\�G$̳��A�>ި;�bٸ�w�Fu��)m;Y��T��V�h���u��i���8RV�_>�/�H�=�]lm�\wQ*f`�t�靨�`�����ǜ����r�븫�Bݮ(f_O�%$��ʸ z�����2	�5ݙJ�%�swX�7�p�wxy��C9L<����-&��2��D�+T�lR�3N)o6ݧ++y��O~[E0��biR���1�<�k.�_�̃���jڵ��\T��fo
���W��tޮtӼ��X�Z�|5��VJ����<�yp�ι�t�����N����\��3!B�'�i���l3y9�W�8p�¹x�%�[XwD�v;��nWw!WjW�X��4�a��D�9;����;��b�C7z�GК����.:*c%>�]�'Q��-���z�ㅬ����z���v	���Fm�+:n>ʰ�D���9��}����X�z�ྶ;Ve�����F�f2RɍWQ�F���3Gq�5��CSW���j��&W8ck���k�c-�<��J�#+9ܦ�+�\��6��\Yo]�Y@�h!3񡱻���J��°��*t���Ҡ	n�f�X�,�A7���t��
��^�ٱ�1�\2����|5�ۍsK5:7��姎�;����^�fP]rJ�-�E��}$�t������'+��˷�7����-V��mE����K�(og�ҝ�dZ�v��OU�5�.�6nȲ�g9O5.&���(�d��ocu��c�*WX1Wc܋��æ��V�u)ܳ������?��h�4�wjcm��|���E����]�yLt��p�p��a�T�l��T�`��&fXv�r��2��	'={�l��tyn((q.��S�M��P�!]i������@Ռ=��K<��b"�.�V��ӥ�HN&�z�,��b��ݫ�)���"nX�6i�W��M��;�X�p�����Ρڕ�7�n�6�&�C��bѺ.PcZ��Z�TYk��Y݉n���D�uea�G�n����K�N��v�',5O�і�l�P�{�)��� �'�q�-ܫ�rR��ޠtq�f
�� ���ϋ��3��{�!��ۻ�H]^�P��v�&v�՚t�˟t]3�����$�Q-i6r��w����W���m9�̑�(��r�*%���fV� ��F��.�a�&蛼�hS�_h�F�ÜLu�,����u�:Ԭ�/Z��D� �ݹ
\v�'�%���
�՛����,[H���Yƃ�J	ː��`���(��kZ{3]�w@,���Pk���`���:�4�46^�1T����>�f,{\={�ev�5`d�E����/�J���� �b8��c_��ym�1`���/q}ы1�}�e;�<�8���NO��1�09F��)n=X��\B��>��k�a�;r�G5WZ�Z�5��iʾ��u_�"��k��y��&¹�%�����Zy.��~�MS����%L�t���zi��ܨ��|�!b!��,w��y!Ӳ��.&�ݶ��yB3e�e���R���]�q�`�I+�t�)"�1|Zd�6;'V��Y�f�f�ХX�5'�P�no�����c�F���%9t��Y2c��z�.����(�I�b��D��WX��n_N��wP'L
��K�u��H5t�w���v�,�f3{z��ȕ��W	������6�m�m�v�U���*G4Yr��k.m&;�Ȗ�ӎ3�dn�S.m���(Mh q��k�wE[�������\��^ɡ�d����S�k�WM�bt��-K�n��/(�F&��:���|h5إ���n�* ���AY�C��1����V��;,��E�qG;G0�n�JZb�ͩ����UX�ݩ �8���2ko�ń�f�"wks��nLi��H�S�[�Z�彌�u���f�r�Z|f`F�U$�M������YxzuK-dB^L�A[x$�*��*=�F�](�y��'a�ݧccY�iٖB��x[�GSdu␩���m9w(P�;�2�Q��RQY����Ck80�엘zv	v+���\Jc�">����"���֛D�=q�����|���v{��%���k���I����y\���s���F,a�ҦhL��jM�m�B��բF�ØƋ
��<�����Bfag�Y3H�.��.O{yL���eeI�	��٭�Ui�t�W�z9���Aϑ#���DvVR`c�(k鴬�]�IF)go\(�E� ,L��1��ʙ��K�酷�Gv��)��6�4h%��g7�����9�GK��-@���bS�C��;O�9�NU"V�^�5��Õ������w��/q�o�����+9��"+m��V�)QAE;J�]���m`zEm>7�����nV�H�q�C(��h	�e��|�N�WCE�;�N�h��\x�5��a�T��U�������wK�/u��B�:��C]�)Ms�bg&�%�S�v۰pEٖm�&��
���.:��V���ł�qN��͋b���1CFr�2�G�I�.�͑����R�Ř3kc�AT$��v�+_C2�Y���B�#\&��D~+�n�=K^I:����ȜY���$nZ��r��:�q�9�]�X����'���T��Tm[����gx���_B�akf��S3�;:����s�ge���vm�7S���Hwc�Z�
��&���y
���\�U���ʺK��N.P/�7�_sT�&zL�2�<�2:$���E\�
�z���M�)��BD(�G�rG���D@�����6}��]��'[GN2�nm�n� �E���(�|8(���y	��f�Ttv���.�涜
+��9"���֋�U��뼵��y׷[Ԧ7Z�b,䥐Q�B�[G�T�ժw�� X&�Yt���n���k�
�)Qc�cҎ�_;�X�7�qް�H����YoIk{@�#���ҹ@�U�F�G^�r.���s����q�Y7M��S�8l]G�(л��2%I)d��r�d*�d��|�T���U�R�亓�s�X�p�ᴒ&a�Y��u�ɔ)b�Z� 9�}�����FO��kެ�#&�q�&uf�o����mtwu�-���#C��]5V%�ik�#u��ia�\�&u��WaPy��,��ȁ��� nb��7��#c����u�`*H�R�]s5ˀʕ��U�L�.�v;�c�e�D-�}�(�T�	�Hew4�i��6X�}&��m�h=X��f"�B�k&p.d�y�w8�X�b
^p�mI��� >�#,n���r1m:x�8,U�h�ï�6kP�x�N�B`��W���w��ۄ�e.�u����9)�^hn� 7Lu��%��k"i��R��c�u
G���з6�n%�V��Z�Tb��{R<8Gf��v{+��u���ǹ���Z8,J��� [c�A��ϲ���
�Bq�#��C�!w1�R����A���F"j���u�Z��1wC&�'�81����N���`\Υ���x(	˨���4(w;�H�f�
����֭n>��/�X��&��8�TH�c4^NT���	�b݀2ޠ�wS�!�鞤~,:�w�Ga��7Cc4��R_uh��trf�
۴X&졏n��,u7}Y��Ρ��u���E��#[��:k�	"݈�|������)�-jv�-f��bK�`����I%�
�R�$`��A&M|����i����������̺�
v�����yie^\����h+����O��=ȫH�{s��x�Q�[�m�S��|�>8ek�ڡ�DT��OE�vو�X�D�@V]��M��;+_u(�
ʌn�6��fogR	0�vdq�r����	^�.N�0%pw�[ެ�Ob30
`*�׹A����9H1��}�9lᆑ|( �r�k��P6bu:^��-��v�*��YJ��;�6��#���7�8�(}%b'U+��x�䋻��**өէn�L^SĨT�j�:���ݾ2@�<�Z���X�:��^�`{�J��r�
�����d��$n9�s�e���m[�2�1�ё�.�*�>=��r�[���W���
:M�W��a�$P%���J�(��� #�RnR��ne*�e<�w��g՛g��Z.���>ǫjD�b|�P���]I�:
�[}D���y�Y���0�����ԃ'8�KG���R�]�����w�5RXPu�ˋ���"˘�E�fvn�U*���J���,\�:BS�Ho,�DBn�\񮽽щ#��M��V<���B��Le�6L�/0���ջbƑ+��x&���Qo
@Cg�r|K��1��H�!��9��(��˾�� e��b���Z�E�R
���(K��qT(kS��2�㌍����=t!��N�Εae��]7�d=�J�b���J���tee�6J���H�"�\�"�{]-�T�C5�q�S����v�
��F՗�������m�	�50r=���h��eL4�)�d�M�����ܺ�}X��[����"Df˴D5`=�O��ܱ���t���m��bnv�S�mܣCn�h
aVU��G|0��^�O]c��>�}6/�{Ce��WD�ȣx�1Y(3�̳�6�
W2����M
�6�����P�3�=JбZ�ޮĻ���كB�ܦ��x���X���S�=�;b���^�w3u�Ұ� ��A���,�	΄o.j�ngV}��ʓ�}}Q,��YtC�/:��
�f�����Wr��pwr��f�0�)�S�83��t�VX�GO��7.�T�}Ruc�M���yq��k��\=�C\�ε����Յ��F>��'n��p�-!��}���}��XS�v�%�YWq�h�n��H�N�y�lK[Ld��|�(��Y";YF�,�����x��mG24*.Y}�d�W�,��Ԩ�j����6���fTD
��)zoy�L��YЕvY�����71>�����8QśV�qާ��N�r���C#��D��ٛI|��e^ќt�sd�4���%���N�FaXX�{��r�E!�1�b������Ħ�����[C˶�^
�)1`�z�g
��慝}��,��o �'+��k���ɥ'Z]�:�0�]ʃ��r�}�lh��WN��&&^�I��>.fq$�,�[c����@�������[8���sw�+U��e7�F�9��x�7��驳�"���S���1t%4�ãu>]��st�'Yf�w,�&㙲pF����ъ�����QL�w+P�;f�T�J 8Q��_�c�)���8������� %���Vn���j�c��0�`Pqoyż�y�}+F ��%X ���lx-Ov1�HU�z"@U}���}V�՚�t���L]��	�|-حc�Y7gR���М�����T^>�ۓ��@32������Y��d�]�LeW:�$.u����W���%Ŋf���2�u�ܸK�8��
-&�o�Vfb�mkd*�\{&QU�6�̣��7��`���m'g��MR�+i�Q�SnH&p��w�6��QbF�iH��B��w;e���+������'� 6��T�S�Fh�zĆ�E)!Y���묳�2���Cֲ�Lԍ>�ƒ<_}����m5c�Yֺ8�v�"`|��KN�X��n��,n��d3M�wk�1
j�[��f�R��2���e���,��!ֺ���A��%�r��&ݖSV�w�AB�Ē����;��ڭ�e���		�����F7X��]n�ƭ� 8�����ܷ�Cu�����93�p=�H)K$������u���	�e����J��˭�j'k�{peӹ3�b�=7��5�����D�f�ĵʾ�AfS�К��b
��N��Bճ�
Y����jKC\�j��5��oEK3����A��*?��m���=WC�{�[;u���k�9KX�f�<0��VJ�a��|�G��+�L�u�n����z��1�����P\�nIoi�ep�l��Wk<Iv��f��ɥ����׼���AuYv��,�1���Q�(� ��\�|�&*<:�;��h0��5�y+��V���X�0Ʃ��^�
k'a�Hw>�S����	�.u�w�9�!};��{R���kiaZƦkN����L���,��40,�H�.�={i�yC�W������^����VJ��Tv*� ��Z��N������6���'u�{�ml��yX�{���#�
n����
9m+Yj�45,�"�7��u��gp�X�O�����ڂ1�nP�I�*���W[-�֑�i�o�U���-#SV^T�(���q�NйJ�	�e�w�kw�o����mK�3x���wVX���LV�@P:%L���'8)2o\U�LT�jt�G�G��5v�@A}��X��E�f٩����ʧ;y���c%u�-��eSE��ׯ$Urku۰�u�]e�9X�(t�N�U�t�[-��մ��d�}J�n'sYE�������é<|񁳍��|��}ײ��J�4$��Jp��V[5ғ7w�e��WG���mU�yZ��An�;�f"���(N9m���C��;!��.���8��Zk7I'T,��\���v.�V�%�AOnS5�{%��BDqH��Zͽ0wU� �D�޽Iޏ�'pd&�̣W����#��֛U;-0GL�H�SY�L'�_ r�Эcy�8j�p�D��y��]���41X#
�f�%'Kf��m���Rys���Wg5Y��hch�iH��&UYj�t�[8;@
�� �;�6U�vq�Ȕ��I����s6�.���1Z����Vd�1��s^+��X+f��Ѫ�d���ڐ�t�Wq!U���a�3�c+�z� �y��RQ2F����̨ 6�*����do`[�����[��&��]kc��ҚE'�F�*�
7����<r��m�Gtn���fd�I���p`�k��9���y�w��}[�����5l��K4pڲ��hb���t6e�Y�R:Q�y����"1�_ct`za��Ȯm�0��r�T�J����X�$pYܭ�Y(7��kUٵ3��{���i"`��[��n��ki�0WU�wŚ Z*bF�r��&l�)ڡD�n���l[���WJ�ixy�b�E7��>݀�v(#d�n9�U�fgS��U���m�=`��Sr�sM�~��p�ż�
(� ������Y�횅d�G0�E��e7�)QV���
Dh���.����S����K-*B�fۣ�%�lU��]�v�uʧVDa҇)��)'�3w�hX޽Vo�[\%�ću�er�.OiX�7�Rm��:���1Yѕ�AQ&
��im� "��!m^��evI[7X�q.�a���l�M���p��`!�JT�)�9-�u���ԖA��u��6o�8x7��n��@�N�(d������f��jzz]]QK9�ԕ��eP��F�Z{�oo=�놛#��Pt�,���mvU�9M7e�`Z��M/#�\��ƌC���,[���p(�*�x�g���Ϯ�>ԍ'����uu8��ݝCe<U���S��G�3�e��{�t���Z�6Kv�|��nleۭns���ޚE�Y0<٥�m�,����>�}J�B�i�y$ep���g%�Z��V�KX��������Jۧa�Ж�m0���1��8��)�f��z�;T�j�J��yv0��ATqҖM��gE�n�qs�6@X�"KjP6��:8�Z�&7i��Y�V�b��� qѵ*���-ڬ]8ăg0dz�qj�;-��5�N����`��ۺ�O���4�fp� �-R���evR`f�t �N����Cۊԫ�K!W�ok�䱼����dY|�<;C��F���O�8Ӄ�!�,)�n+�Y�v���n�{Hi*����by�&�S�,HE����o���7X��%��*wթ����`�LђS�V¹�U<:{Sy�F�1t��4�pn�b[yˉ�Q|R����3�1ɐ��(Z
��M�����N�h
���]�� �n�����7 [��EZ��b�ZN��Y�~0F4!ݲ�n�����!����i�7.���Tu6hŦ�+fc�� ����`�4ƽ�V���Z���Z��	>�Y�]#K��;���fp%I��uϭꐸ����V������]K��:�qq儹��	j�� /�vf%F�Qۗ�L��L��Վ�_,ՙkq�fg����-Yѿ�n�7���RL7�8��)Ѽ�8"����-�ǘ�l�qO0=��+4R:��t&GD��4d\�\�:��U�:cmG��e�ݥ����a��V�GR�5�x���M��ˍ�)�Ç����)�Ѧ�P��J���\�i�V�Yx���U�e"��W�Rc���0s�2��ag3υf����QE:��&^\Ue���e��	�JH����;�Q|�K��e��ñ�7�[J�R���4V/�kj�U���ʔ���+e<`qݠ�Y7��>�5�Z�3�E`���g�꿊 =�hI�o;�U��t��me��3-b�F��{H��p�)-�y�K	��Q��@S�ö؂]\&��5�gY��B���|Ԭ�z�^��kWD�ͮO�t��:ٽ�ƨ��]��C�Q��
�T/�n9�&�M ��/2�E�k�Tή���a�'\�\x�;@[H\��:ՙ��4�m�6ҥ��Y��$6`��R��H���*)��7���Û)46�\u��8�Zt5�r|��p`���1�+�^g�wr����9[f���+dzr�W$5ǗL\B��n�r������,"�c=�\N���``�b����z"���v�-��E��;��&�V�8��dR�w�*�>�kj����Ur�9C/�^QP��)�A2+f�r-؀Rɽ
d�e��:��0�N�Z��mXGwdfɖ�+���Ή��ɒ�D��ܘ��v�B͛k�m��=f]���JwY���|Y63�2餷��-u�*5��G��j��ݮ��)ٌi;[��!�s����*���N��:���Jͺ;��V�!���Ż)e��X�����pن���9�W�+�vh��-�{�:�R�Q�a�t_g$��u2��f��e�.�W6�m1G,rz+h�/�"��7X檺�F���d>�Z}�^G��_cD;�mi�%Wn`Ӧ���C#V�Xv�`c7��B��ag;�Z��g ��Wz�oJy̞{z�!���H�q�y������t��Y���ܔR���r��/9uIr�]���氎(7�"�:�	wg#�]P�=4;yR�F$]<�r�6>(�˘w< �j����;�o4i`�\�: T0i|_n�����Q/":��Y�d����*�����b�h���\Ɨ[�Z�`s�����$T��آ�kaL�7�v���ʦRa�5f�������0j�t2��DkJR�,�*h9��������\ڳ�#:��򊛡iWa�r=u1&�m�@W
�.-I�c��N�K1\��wE!�k�5J1�WoM�i;��t�x�@��2:Q�p�ۮ��D@'ҹҚ��XkqI����D�"6\E,^��)klVjᳲj�8���i��-�%��.��F��wc���;�YD[��H�H�Bg{Y߹QCa��Y�Q���v��0-4���=���Ȅ�O7���e���Y�Q�t_3[;��L�q�E�晸�r�kV>kUh�e-8	
�wO6��u+]�XT��v}�)�����VJ�=���Fj룼y�
BJ��8�m�Q&V^B���ܙ�!�WRxD(o��\��P����QKT;�n�84�d�
��@���Wn@��DlN[В/;u
E5v��U��Y���"�y���B��X][�U�VYծC`�R[T8@���Y�	l>OVq{br��#���v.#�3f�Nq!5dͨn+u���}-m-��	*�\�)tҝ��]�_�T�OYՈ�t�s]��gX�X��)7UN2}f��n$�W��wxm����4�&31TUʤFf	���e� �_.�:U!��e��՛�,M�on��-NХPko[��ƭX"wS��W�NeJ�m��|�=� ���W|'+�q��4�uڊb��d�����̠:Z��������>l$��!�˻����rcԟu�&��
r���f.8Y��$�=�y�2V��E��לVhgI�YZa*��RlҏY�1��t��nL�2 ��;BP�E�4��K��ѮOfK��d@���(�ф���sJؘ�w��!Z��qΤ�:�l#�-!۽�mʸ-�+)m��W��]NH;rރ�uW�\³N��Y'7�Ba銤�b�$���]U[
XeD��u�K�s��HuݪBňԚ�4b�lh�A����Ӯb����C-	 !%��$1���M��"�ђ��e�(���ѻ���N�H���e�
�"&L�!���MH9pˉ4k��f*���s$��`ӻ�q�Z�W+�fwu��(�wt�.wn��I�̈��B,P(��6�d,�H��t� ���cs���snR�3)�sd��Dk����&()�Is\��E0�A$�J#$!��� ݈fI%*s����Et�N�L)�c3OͿ�??��߽Q+��|zG�1R��B����5��qS�)[�r�y�X��T|/-�ۛ:8��3{�ڛ��>*up;�̳u��eNa�<� M�T+a�������5R���j�t9j�����p�9~(YRgoJ�̥�=���]Y�(�Luc膎�l��R�Y�

��6�[Z�˫T8jie&:R6�[]�7~���3�iZ�GncB��^U�q[ϸ����0�
��߅hū�i��v�C���L<1�4�vjw\mFi�b���G�T�W���� 8��})�� ��G	�R��]p���;�#"\�=��XO���9�/���멌��ro��@��CȱQW5���_�a�|�3#����n��v�� ~�Z�s`�J�}3�T��B���ߗR�YԜQa+#f��0;��l|��/��Z��V�VN�y:K��ݍ�?�ݶ�˵	:]#<Y\�#^�鮠B����*?iJ��֐�U3�*�O�|���o���P�g����H+��JJ��Gc���,�*h��|!B<�G�"��k�D�����Cj�\ ��P<d���x��x��Z���U���7qa��״�u:>#��*���kB��D����EY]�]����l!Y���YWMm�P�a�6���]�����ک�v���艅t�'�Ԍ�����//`J<������[��q�u���&k��o�g%z�Ҍ��s�չ2gOͺ�g):���	k���ac��sB�%��v�!�y�Yl��n��emP#L-$Q�|�u�����ڿ�;�Cs�븜n������f�[͊#����N4�ȁ��jP`P�ǡ��w��\��T4/�~s���L/����y��K��;�P�z�h
�Ĉc��ȍ$\D��F�#ןr���h�e��T99��rj�N�=/ϊ7�p��xX��S���P7<-��P�z���?�����$���̩�T31.2s>q	���2nl	����:k�-8��<,s�����.�W����r�u�����MF�˅���F3\�ɧ��N�w�o�����]��9Q�u.V�0&�by9��6�Vm�d!l�G�&67e��E�7��t�{��W?C���;V��L�q�g7oem�������D�����j[T��g���@
��u\#,�3��s1sɌ��k	�?[�+�L�l=R0���w^ZN��U0����ժ��]�fR#�;���r�>`9������K�x�>עXC����mgC��9�̕�᱗�^_i�C^F::��V�pRR��~'&��U��+��
����tU�)k!սM.���?d�b�0��KdŶ��R�Yf�h�R�L���Y̋��,*�»��q<.8x׻���k��ȱtω�����4�G��UU{����_y�Τ���82�*d�"1�xI�y���]Q�*b�#n��I N�3�I/��M�`m'��Ũ�t���	0���\it�U��岲)��o��}�0�ȃ���2x/nT��hO�wTJB����g)���ʖn��_jv����t�3�����ͳ�
�e	<�M�U.T�Փݶ��M���|K*�#Pvaq�����󄋉r�k)��F< 6hY����/5L�R�i�*z�5�`��(h2�fҤ�r�x�g�ثg��]��|�ޣ�M�Y��T���_���ꘚ�2T�10�ГU�V�1��1�߲�
�%%��kΪ��ȹ�����9��o���/�+W����k��@X�)��(��+�Ry���v1+(q1n�tn��[��K�8��H����*�e?��e-� �މo���9�x��!�l�1q�+M��ԇnxT��I;2S1�*���vd��(�[r����ƭ�/������u�L�\���)�,�5n�Fk�>]H�����B}k�Ҡ�I<�B�jXЦ<� �2Ԛ�4<�nTض�S��L�2�I$��t��ͷhl�r��ʈ�M���ay�O,9�����x	�)�ʺBS��|�nC��Wήh�V7��k:k�za��w�	:��2��5N�Qd>�[0��\�}�jk>�XO��R]�~>9g>qp�L��4V+^��lF'!���Y0+�\�W.}��A�F�Y~�]c�g�
炡�k�|��L��q�)��T�w['
|�9;X��?N��`l{���F����r��j����Lz�?�X��-O��Y��l_1V�+�k@�Q�p�W!��e��Eo��_E<v��B���5�g[4�[`F.aS�۲K꛶d<<^1�sfX
��1�S,R��:#1Bw����t�b;�U��P\Po�u�':O�Q�$��N�+"4���9�
P�4���:�� �q��D�	yuQz��Zg+,P=G�U��Ґ�,}��v#�n�k�]���Nc�ʼj�3�!uԯ�5<��,��Q'd'A�C]�����>U��H]��BUB1�r�&��]����M1�����FF�����Lu�:G�T9W��$��i�h�����z^��{��b/!��r+��2��ո+�ɐ��În�[)����+�B�%o�45r�R;//;�f�+�[�#sd��Ƌ7�����>1���fw:^RF�m:�}���b��D��w[M�};(Q�>P�E�����<9�.a�ҙ3�;��摚�2�@C3��A�_
�_��/fn��������6c���zS��a7�#��cT&�۪fED)��*��S�y'nc�s�>R9q�G~�ǛgSږ��/��\��Cj�9 �D�s�b�P������`� .{�E�C1�i�k$�$�Rf���ԃ�֮C�?Wܕ2^3,r2Ҋ}!Ut�U:�H�Nt�D𺐈x�+�)��P���'�evm�Q�屐ګ��c�����.`L%��XG @{V.>����AQ��y�ʉ�Uoqv��b�D�nB��s\(T͈�	��:܀����敪��1��R�,��}�g�)B��r���[��8-4	ɚ'J[7M�̯!^��^?B��!�Q�EiD�TA�F���HdcUx���}Hk��G��K(���@Wۍd1���1�g�xG^�W���S�-l懦?��n'�����J]@w{�B�|;O
*@cc &�ZfF+N����J��5q�>=�pV"���qX|=Xb�ѱS1�9�s>�lndf��5M�����&2րuS��U�7(����ɂw��N�ɫ���=Z��
�G���:�;Cts	�!�o�F�(F�lٔ/��̧�*'�dY�f��)6���\�'w�Ѝ^'�M�iv���X���f�%.3���tB9��K8������Ln�i�ɯ<��fc�Hf�g��7��m�2��^$�t��es��5�tWP<o���P7*��op,���-eb-��Yx�1q-S��̂� ���������8����P6�o�u(q���a�Bk���k\��4�+���Juh2V/FO�el\��J�����}.B�3�XR��lͳ��|jg�K]�w�r4���>��\+��ծ���� �1f�΂�Ɓz��$<��#:"�:���������q7��)\�Сlܻ6���W�.�?zUq$ai4�Nq������Ū��ɫC �H��4t�<z�2'"bF��N ݫ���c�|��;$LJ�tg�GoU|�֍F$ �5ۭO������EL\��i�� :`����"�\Oʁ�!��=���x����H��=:�y��V��${����mTH��<ɓ6�p�G�OF�#��qAN����z�:��TkegN��k���L�h�8��S�T���J��Uod�M���D�n�O�V��6���D��Lރ�kNR��=y����ݯ� ��B�A�:���4c�;�>-�NQؘ�ǯ*��!"���wׄ'�k&\B(�8�F' Z����2j7�x��l^Mj��Y	;�c#\���vJ�F�x��1Wn���ӵ!�{y˭s�R��&41��W*�b�e{401|��Fjt����Վ�Xys-H{Ej�Mp���R�'1�gaɇ�`p��@
�q�1h�:��Ct�*`��7�h,�W��I��`��f���H?E�wA�����t�VT�L��! &�+#v^uy&�]`UN�MNО��_��ٸMW���_�Ӓbo�;=Y���Ŵ����3�^����'�3s0c9k7��5�2Y�j��d��л��H�V��EkI��R�����}�+@k�{���[�1W<Ax�|�4�`�+
e���}�^���c~ق�阦��-�ώ��������2��1@֧l}z���`#����f��m�I�M�#��̢Pqk�Y)�.Y�V�b��RP��ab�\����h�F�z�̅�V.�6r�:S\M����&�Ƃ�)5 @��:�|���5����;�0yˍ)a�/ee�<y�ǠM�tP��8^vWlZ�dѶ��8�aJM�κ��J�@�>W���NN�3��{��=A���T6-J�<�1Y�ڜ6�[�լ�Y����32�M���o�8$\x�K3�L��Ǔ ���w,�/�:�%^�w���*y�&��S� �`c���66W��+hcM:=Ϣ�`M�c�XI�3�ok��.pCg"�`)��:؃?)�W�s�*��%Ӽo3����s�p�V��hj�3]��8��3q�������Fǒ�KF?��G��m4����Z���8��j,ʬT��$TҴ��wK�q�ԇp�I��I٣p��k��2+�fI��v��V�x7V��y7R��9�ڰ������w����T�������S5� �sH�[�z�}Nt �>����\�L�5�h-���0�WJ�#���p2�X��T�"�ufɽO��
�+�����ҙ�
9t�N¹ྡ�k�şp�)�+o�3�U�O^��*�-L���?-8�`������,1A�8Eczhŝ�)cz̯��j+vL>�%T��놤�e��ƣ�ڿ���VcD?`��K=ޚhgOgX=�=�ě�^r�q���(�D:)Z��Z]xS����w�����H�C� xYC\+ܙ�ʬ�J/�A�îAJyʻy�AVuԨ岨le<Ʒ��	���F�m��}}�?AZ����
e��m�K��*����$�,�շp�uJo[��V�N�@�����L������ѐv��մ����Mb�xT�NȲ��ү��Z
�'^�T�����â�P���A��Յ����U�o�]Wy{�e?8=��{��X}d�rz����5�ii���Q��UiN7F��{��v���ȍq0�9\C�q��3�x�Pj�LIi�W��q5::(�Xy%�p�CdM��[q���=j'�,o����]���g0��t�µ?�=+���,�� �h�r�
v�A8#��	)mH�0áӒ�_e�4�&��c��0�i�nH�x�E��+� E)DC/2*���q͙�E�������s�P�F3�.��)�f0�ґ�3"�um�3"��G�4�e�콹e��{&��D�WtОsg#,;/��ϩ�ŵe�Z%C��3�f�y�9SAv�$��TK�2�0��&a���"�v�w#���}և��=�w/�"�:�wg=���W�2�h���:"�>'X(v�>�Mt{�)�w�j]m)�>�,������$x�RWe�?Jӄ�9�I�ރ�4jR���Xm�P�6��R�Y��S�'tQ���8w6�S�>g�Dqg�_�e�tsqHE�Ђ����m6�S��q���e,�Q{7�p��GI<騃2��|�f��gz�2��LWfu� �U����;��WN��`9��"��:Џ7l����ޱ��Į�c�%r}�u��t�p7[Ӊ����`V���~�l��8��N����})i𕍥�A)��ޮX��@4zL�5y|����(�z��EO�Ћ(���`�B\6���{KgI�9ߐ�Dg�,�#�@�(���@n5pÙUC�:�cuc{=��M#=�i?|7����y�������B�<;O
<���5�\��(*�_�l���J�[�Ծ�*�;�N�x��Џ��YMn0h��Hhg���Գ�<j�P	p�m���;Tpٜ5��I�g{�b����^pxL���6��TSԕ�k9HOf&�mj��/�b��B��\�I���ONDi�����T>��~�鳕RA�Ғ�oIC��y�4��u�}z}=���Di�f�/�	�Q��-���h�6���M"��t�IMT�)co�emn�Õ�o���lͳ-���l��p��H�s��^Ke|���,7�42��U�uo��p7,�x���Q���;<���3�*1:������w���']ď���=V��?8OD=��u���dŲ��Ŗ�ө-����9һ ̱��\A���^�ǙPn]X��㣯)��7(�HH%�v#�S�[@��( :�N�!=}�wWP�]bx*��,K�0�k��M��j9zS�y��m�Dn���b�V鈀��|�U9#��mp*�X�J�J ]%��{�1.p�LKF=7f�J�؅�4Y��s�>��Q������}����s-+X�P���+�,�fW�ʖ�Ʊ9z.A��ұ��vS	�om��T0:���ۆ�D+�`nnk�Գ�}��(�4����O#N���)�8��l�n�q�9��e�ؚU�4�wL����w��#�X#�Q�ʥw]W��@�]�"�Qt�9�����0n�R;mpwŎ�VJ�횈�nQ�:����ך�Q��o����(Tg5.���X�JN8����y��>��P�Hԣ�ʂ	N�����r�(e'�n�+o���K��C�Pή U�Ĺ,c"��h*�eomk�4�*붖&ʩ-�q޵y�В��r	[��lZ��r���z�rwĬ$ D�L��	X�i�g��7-l�Dmo6�Mk�������Pl�Ӵ�+�8{���2Ps��Y�_�d���j��@�{J��F����)�]�#8�-/�v���rx5.0حݕ��s����p^���IGS#������R�8�_,ٝXu�]���sO�N4{AWX4.䥚�o���5}a��R�C����7�Ǳ�gbɹ��T�z�zts�X)�V�7E�d��f�������nE�ٝc���"⃶��=��t3���N��$���CW�f3(t��&GTN����3�4M#!��$=}cR�O!���"��L[L���22Wk8
�M�dhFþ#h 7��E�.։r�+��[Gt�Hpw�H�.�&��t�����T�Cm˹��ҷ��"B!��)j����9���{M���v����NW��V1=�JD9�g#w��xy��足�!�2�Ƃ��g)�pU�cU�膙������&���39��W\��̩�32��(o9-�����ȸ�&��KP�Seň�ĩ5r����\J��l��IX9̆�P�pFS3�v���S�aT&w��̱>�J��Ֆ�#OhB�Be����&a�4>�f�Nh|��ƊMN̬U���rg4�����\$�&/������[�N�|x�b��3I��cc-c�K�&�J�ʺ�x%*,� 9��Y$fG���lE:�
T�y�H�ky�����j�bw̽f�]�cx��k6b�Ӡ�@Jk/ �R�v�����Vt��J�9!pA��|�m�W$8+$C�Z��PS��vz˫��*��1��m�6�ǧbޖ ��w���u�J���n�2�f�ɨ@,���Z~�ܺ0w�L23�)'0�&r������񞺮n[�K��)�d���� �wW4N�vwWs�d�4$����tL\ܹĨ�5r�b)L�܆�ݹ�,�(h��� �`A�`�2h��0c&%&ff\ݢ��DQ(fd�h�D��,�L�Q�1J0a��4!$bB���: �l�2��#lHa�(���J�b�I,b���"BF�!�JH�BQ3��@�uvB@&I�ݘb�0�6�1�	�	(��I�pdi2d�L�7c$(�'9�4�C&$A�I�b2�����Q!!��&)�L�D4 �A� ��Ț
r聓w[��)&@��A@0ER��-��`��`�s|��Y�
�d�t�D�inٽ��آz��n>r���f\J������ӅHg ��lc�fK���N�c����h�5�y�)���������Er������v�����}ק�o�G��_�{o�oj�_�����6�o��W���_W���F�*�.^��Ͼ�c�}�,�ĿE�z��zU#@�9_��o��~��-��~��y����^���wo�������������}׃Qo�:�{�u��םk��z���׵�okſ=�y^���׋�_����`�� >����g�����V��t��?u⽭=�}��߫��6���W��m�v��������nm߽�˾yW-��\ޯ�^��u�+���ݽ*���F���m�|_W��y��^��^���"�F��و��/ ����n�,{�!H��7�_��^��x��7�7�������Š�����U�oJ�{�瞿��U��鷏���6����r�}�����so���m��o����x���.~>�DD!��\��1Fӯ{V>���U����ۖ�}�}�v��������߭��[�����͹�-��w���[�����ϟ}_�~>+ţ���׭����x�����z�����~_>�_��ߋƯ�7����F>�";��(
g��OV��I}��^z��^�w�W�w^��i�~]ס�͹W�����o���6������^߭�^
�߿�k��ϭ�?}{�w��s}mߟ�}�����������������lyLE�>�>�a)��L�l-�7c=��w�}��n�ֹ��_��׵�o��_���k��W����-�׫�����Z|���ץ������w�W���w�����y���nm߿ﾽ5��BsU���>b"G�#.Q{/�ǹw�T�;�ch����`w�I�1��1y��~���^ƣ{�ݽ���^��η�o��W�_��ţ|W�x����|W����u��K��{޽y^�u����"�[D�#��^�7N�����\sP��1��#�D{�\��?o���?<������~�_�>z�{U��_�ߞk����nk����_���x6��o��ſ�ߝ��v�M�o����~�K��>߬ǄX�,1#�X{����3��Z.��K���1�@�4��5 <Q��}���x����o�<ޛ���Ͻo�������~��������[��W���soW�~�K񷧍�mߗ���O�ID2#H�@@DNs\z�~m����TE�t]~U�x�9>�������sۂ��OC���OU1��lv� �XcM�ե�n���k�R�=�ňى�jv�o��"� 5-TM�3O}��	�m���6����"LKSD�(
KvK�d/��N60�yHc��<��=�"(�t�)[��u���\��}�ׯ]�����}���޻�����}�����?_|�M��yڻ�sr�׋�o����7�����������o�;�~�Ư_���W,x��� Exp�&������n����%�O�~�͹�W56-��ߪ��r���|m��ߛo�z��Mn_��m�U���<�|[�o���֊�m�^��_ͷ��5�����x�GD����DH�_{�ڹo�r�o�o?��+����v���湧u��m��+�矾U����x�ߝ�^��w�޾���o�ܫ�﷯�z��s�s~Wߞo���7������<��(�Pj`z!�����`�D�.��\�-�x�|�����|�x׏��o��EDW��޼�KO���"a�<DQ��d��c~Q��\∀Li�T��#H"�=~��5�?Nv�;DϾ� h��>�D�~�!���7�_�߾^��W?�x���}�k�ܮ���k���szowί^�o�_˛�wu�<c�w_[r�^^u��W����X��F����5��m���[Y}xͤ���G��"��"9����h��ϟ}[��_�o�������>����}��������_�>������������~u�[��u�zm�ϝo�x�顐,�!�1����L�ʫ�՟�EU]��>�ADz�4#�!��7~����j����W�����x�Z7�^���zߍ���Ư���=-��[�}���[�^>���<׵_���������b�
����3Ƶ1C���}^쟹�Z��""��(��1f!:ă��1�/8@z�0�1��6����x�������s}[���\׶��Z=��<�5�~5�ڼW�Ͼ[Ң$#�yD� �D=�x�����T�Wz��ҵ}&(�̘�C#� �kQ�����hߪ�ݼ��~+ŧ�_=_ͽ��m�����/k�o׍����ך-�Hሬ�H�	�|w��=H@F<�}����P��U�n��<�)��?+��m������瞛�ۖ�{�k��W��ۼ������W�x�����^���4��~�Ţ���ս?���_���5��W,}_����/�_W7�n�������#��>��e$�^��a=x�ފt\YC쇐=w[+@:V���[�˙vy\��{��0Qiر��<��AX
�ܫ¬�s���C�UM�m�31��R���V��ܖ�]�պS9Sݬ�*�)I+��k���vpA�j�2����]�q9�.:������w5����U�so�=u���}��o�ܫ��Ǻ����ѽ��{������5�^��^-�x�W��}�~u�o�}o�~��{Z7������[�m�{���F��#����R���&�ӝY���#�G���LG��Fm�k���ż_�ߞ^և���y�~��o�{Zy߫����/��m�{���^��77�^�޽-�]�m�o{�5x���x�~u�Zc�#�>��~�.�.�]�[{MGw翻����|^5}�������U��~��Cb+����W��{o��~�om��o[x���F�|����ޯ�{Z�}��������˺{���w�DG�H�}�G٪����7���z�m�Rןޟ޾��o��ƾ����5�ow��f"�v�|鏌E%�H�4!���$�q�.	��B$�3S"7�������yW������o��כ�rѿW�����p�b"D}��ls\��%b��|�7���_�x���W,~����kү���׻w^z���ž����^�z���o{�ߛ⽮m��η�����ߍ�W���Ͼ��h�۞���4_W��5�>�~���}�"!�*���O�nϤn�͝��2���}D}V
��,Uh�������zo�����x5��^���O�o���痧�oj�.o�}zk��6��~y�\�?�o~���_�~+��c���|G�a�F��~�hL�k��/g�-�+��#����D"��}��Ƣ�[���z�{W�޵��5��^7��������x���h6"/��^->v�o�^��||[���sܨ�@W��M�Q�z|*��ä��{�|��x��>������^-������_[x7�_��^�r�������6�����~|����E�{�W�m�^tZ��1	(���$P� f8�$���b��}���yD�]��ν�g��չ2�-�������Ͼ�=���_�z���|^֍�|޽}��_��W��7�|��n5��?�~���ήX�^�ﾶ�U�s�����o��~u�6�;��_ݢ�G�!(�=�����wZ�K&V������-�z����ѣr���祿���p�_<�����W���������7�޾}���_W�O��ߊ�o�|W�����C_�s_>��zZy��#�b�X���B|n(����=ѓAX6l/PW){}�)�����r���\ۼ�X� *�E]�_դa�@�rf�5;�nT���B�"�Ӝ�싶�U���Wl_dN��es���ut�S0�ʾ�&��3�M˷�l�g���*Y�cG`�bȷDP��*Lr����}�5�x�m�}�����h|�{��W*�^���|m��7�����y���m���_������w���y����j-����޿���ֹ�>��o�Ƽo���p�C0㗞���b���ٿ�_ן������lO����+���o��񿞖����ݽ/KF����z���������n������m�ο�x7������j�._[~_�~z�oM�o��|��E >�#���)���z�6Re|,�f�C!��|�I�1	(�?
�-�ۻ�_:����m½k����<��U���z�\��^w_V�^��������k�_���{��^���?Z�����1G�l�8Whxmz0�w�߷��������W����}��o����oʷ�#�" ��ȏ��b,������^��+󺾿4hܯW�oK}^/�W�wx5��W�ߝ����1�I�,�b����魪Vm~�rG�o��}���`��D��ꏢ��W7����~+��������{~��W��Ͼ�ms\��6��v�+š�������/ſ�~W�W�;������/8�� b4�!�Dqj ��N'h�̲}U��쮚h��>�>��X���;ֿ+���[���񿗋������}k����~}W�����z��+�������z���_~��B���(� �vVb�{7�)MŶ\�iGx?�%�TH��r^�u +q��3�T���:�cuc{S�7p��9ʫ��<1�)�{��Tr��
a	��UsXn�P`�r�fCV��0�,Yv���I���6�}�o���]l֡c��O��£��������]�!l����ν��NB����T��m��T�^pxL�����hc<IAV����
��#�d�\g�@��j���AL��ڹj���ܻa�� ���͢C�u̬R�[�D
�������]vL����ӡ�8��e��NWMr�J�t�Y�B��g(Ţ��Y%d�
K����0���q���LV��ct��֎o$�Ud�*���4\C}w8�zr4��ˈ�pً�Z�Z��V͂;� ]Y����jy�N��$�_�����1�V�P�U�6�i%o�D�����Cj�\!d�*����	щMd�s��N��8P��U��G녵X�E7_�-�/��Gy��vz�生R���/��%{P5}t�	��P@���EA��t)����_ �e;��������ʃ�\�.wL~B=D�N�κ��M;�cPо��:C�{��]
������,�����L1;�n��n�j�>�8u�k�6��2�V���J�U��;�Xi�Q��C�I��^^ h�����u�w�1}�Xn�I��ĵ���~�;�x�/}[����+�����m��V��2nt8s#xƀ3�͝3�Z��K��r��Q��ˆ����'��B�_j��I:�1���p�T	��(�0IX���,�������Z}����Z�/�:�^Á�ڀ��K�}~���5��lS�S�Y٨��]-��R0>븊y�3���*�j�����JiX��+�@�؝�5�I� e�:f�L�(Z�|�;�i��IX�l�������t憍H�ck�MfG���}p=a�����κB�vƘ�ͥ-n<�*eujש�����Br�t7/�P���嗂��ץ�YԽ�N9��!�,u�j�^�� ��u-�O+U�^����S�0�������oC�C�Q�Jg��\��{��; w��3�i�,D\_4z�����u�L$M�B3�m%\!��"�i�]�U��z�m'��7I:��q۷Ǭ�s��\,��S/��w�e��u&�nN
D��x��4>	v�#ff�^�������_�n����:�^�L��eaL�ySw�ًӣy����o�=h��#.��P�0W�1O��q�ʘ/{�������lE�UmN��ԓ�����J��W�1��L�*BE��6��qM�	�,t�Lvy�9�T;7�+�N�p��=e�
�0��Z�����[�iRC9o����-Yg��ܥ\���%��,���v�!7Y�@c�|�'P�8��x|Os��P��Y8c��NS�:�6�`��j1�9H���6q�Vi��/�6(���n�]ƺS��p������{D�*@�_<��3d%�w�b�^�JnǢ�m��FE9tf��Y
:� � ѕ�i<�մ�'S6����'Mv�{ɶ�qU�۸�5��Wݜ��l��B-�EVNn���*f;,nGҭ������R[����ｅ���\��@�S���݁�ٸ���Ts�tS1���m�����$`̪�W���{��H��s40��gV��(�	��1�V��Cg�Ɏ\��i�F���Ro5���|䩮�a��%�Lc���N�GX-g?i��\5�]���N�֋��(�a�q�u^��̒�Y2۝ ���ծ�A��d�@Ʌ�wO����7�t��;��s�1�"���ȑu�u���76uHE�t���U���dԲ<u*Nr�w#j}<��{g�z6�j3 �q��8'P�ۖ���c>%�7�5_.:�`欽�Z�-����@s%�Q�Ps/���E�j��e�k�l݂�z��T_�ןʦ�,���6����[��EY����1���-u���2�E9���&z�*C��P�4�1�S,��6{"��n�b�e^�L��m�{g��;���Fe�Ƥ�iiq;'V�4���K���P��]��Uϝ-�ER���χ����q������Z��H��		���ש�v�*�,��mi�k��̓4���l�(4���/��ײ��{�e?�jIizm���0�ĸ�uBZ�jp��Β�3v�KW�t���s��#ԯ�	3��wck���`.��S�=۔�!�z�1��=2p�7FG�Y���;Ǝ��,h�ξ�+�}UU����^�� �q0�^:m�w��d��'�GITW�hz�w�r���V�WV$�l�+��9vZ%���:i���F���	'��ʒ���0
S!�]g��<���lp�l����"�Wq2�q�*a�Ӎ���ˇ4��|�A��fX��G-rݭ���R�!.��Ce��b1�j1up��S��ZR+�3Xw���h�JN���ޕ�QմP�jGK�k�Ƣ3�b��^�9xz�?e}ϭ�0���Ƣ�u�E\���
�RI�P��/�GI¹��U=aL4���ɛ+�V�RZ�b�uN'^��N����EM��!=�Kϙ�����ސ�q�R�Q�^�"a�M���nBu*A�[ΝZǌ���1bk-��WG  �@aQ�4v~,����m�.|��k�'Jlۇ�dd�ǪvVٯ��QN�P=��`V���"m��Kp�7n�Z�@�*;���+���}��h����
��/�ve{E{�Y�К���s��Os�\���Ȧ[7[WʞN���o��"��h����(�8�e�c���Ve�"���we��;1T%p�{[������!��"�rP뤬��F�!&b�u:}�u�7YV6�p"V�p�:�M�,Q����-i���}G��;����;]L_�t��
�(�P'�'3�Ѹ�Ce�1=��˼��a����z7S5N�����N���h\*�2����u�������߯��dQ���[���W���	����n�o�䁞Z��kq�G��£�����0;�{�MTK�<�;2k�|�h�V皞طLG\K�<!��T�he�Z�N���Q\�������|��]lm��d�bwp����#O�,�w��j�܈��d�`�{�_*8sݱ�n(pE���Uq�m�S,��0Y����ԭ�Ƥ��ƈC:�\ ����u�u�kԍ}��Kr�p��:ER��,��<��{�/�X�E7_-�--v�߹�ҩ�Un��b���y�p��&G���s'�Nd��\��D�����o���Kj�k�M�U�5�%�M��j�*�S��]�\��+T�5�	w����S�3n*�۔9�wk��Pؾ��jr�9����Hm�[�D��������<��i��Q�?wu{W��W1qK_g��e�ˣ�r��̜T�q=��nk�'k2��X���U�tҥ�"M��AMI) zxs�F�]e��k6t®bO@��Իܺ�e�e�%�3t';캲f�Ŷ��Y�9E��U��]ݭ�q���c��/��PX�ݺ��}�G�]��^8Y��������h�e�%P��n��� h�(UJL�J& ��E�H�	��I�.X�>Y�Y?SLj;Gx�:��͵R+�S̙U�$�x�ɘ�%%�r�Z��R����e��\�R�;.�QE���~�Ƕ��дꫨZ��F3�s�&�J�;B�ff*�Я��i�6�l��l�?�]0-�	�:Lf|��G���h��� V1iO�^;�F�ץ�U�J�8�
����Z�V���u���D�Q�������r���c��<2�U���L����u�`�q�����wgd��`%�^�L�*�Q@�MY�0�7�B3�nU�-��ӒbC'�����3����'.䧖R�ݣ�{��r����v�\�)�{˲�8�.�=u#Z��hg�ݿ�����ҚI�Q8<�X6����֨I�N~]��L��ea�n[+"����ɟ��_g�g^��u\3�FN"���*�xW�Q���q�S�L}Ѯ!�";kc3�ۇv`-���|�i��J�A��]��{p� �����Z�AJAM��2�bcL��NK�c[Y��|�=/�wԅZ�Ȧ�h���/�,�The�yB�
˱q��@y� Z�u�b���*��L��n�"�CsFcb����w7�\��c�D�ͻt5�l��tOo��Y��<t��J�4X�w#[�f�ӛ6q��`��֥A3��K�^��(s�@�=磮�q\���#P�a��K[�^����R���w4N.rC����s´��J]�3�}e[��+�R�ɕl�ռr��4�B��:�ՄoR�V�e�k�γ��_'����VS�܉|�5�+w��/3ciP5v.�b����X��p�:S��Tv�1�r��AW����)��rʜZ=�k�lY
��#[w*}N�f�<�����b�ذb+N�Sk��fܒl;S[<�d��{���tmNǔ�.j�(c�+ת�<J�1�۴nf�=��*G_E�XR�N�D�0��7l�5t�nVcgi��օ�sJhSu�f}��|z�I-���̚�j�����+a����7coJ�D9)��W4�6����o1i���N��.�8*V�1��M7`ꜩΠ��"ڝ��:��*
�D^Հ���[Q�T��U
\�yV
�-*���c��a°A}R����a%0�Ur��uL���4��xfA9t0=��ue k[����W�;.�����v+u+t�X�-��ʖ�jA!���:�p'hJδ�f�[D�:A*�c��B����wf)\�d�٣&�˺Z9+_M��|j�GZ0���]���yLb㚀B����Ss� �
9�}�zt7���YIQ�TX6��p�(Ju�;���GwD7��O��]�D˥E��#�1��+6��Lt3Ё�c�Pq;���wu`ka����t	��h�����ѩc	ݞ6E`�
}Ѭ�y��s��E:�\��it�zE�ݔ�\�U�ǚ�����t�*=r95���^(Q�}m$�Վ����i,���Ӹ3�.�(yr�ܝ�q����l,�`�xB��Yp�F��{�3�)C$���vk�R�±��4���7��2p;�T+�#��0��������UĎ)룪ݫV�yJ�7s!w	�ssq9��K�{S�ϰd�\*M���ckM���h�S��U���5ג��q2�W�Ԛ��WQ�u���X��Kݷ1�����A��Y2u�܍�q��@X�7� ��
�LT+O��;����݂Wo4�k�v�Я{�%eJ�]�-@ը^��)��GZPX�k�0�y��L�νy[R�#���&`�:�䚃�_[�e1�P�0:���T�Q�Sa�����3d��4=W��ͽ�8���;�$䵃F�mҾ&���B���\b3��$F�5��2N:�R�
�8�G�md�6�*�`�)F>SGfLΕ�.�����?����(ID�D�E�D]�HC2�$�ۙB�d�$�LHDC��PJhF���ȒR$�	3�%2	"d"f$�6@s�	30�J4�D��0���PbR0T�\��M) �dL�,FiJ(�M2J��II
���"5&&h�$lP`f��A%�RR�B�L���S2�:r��@�	("��1��pSK���!B��$��Y&db,J1D̑$�3�4���!'u�u�Ȣ9����I�Ċ(�&��9��R&S$X�s��Y�p�$&��QAI�(�2�ےd���ȂaI &	�A�;���Ck3h\�x��-��q����:I�B��%%5)'�b�2u�A�'$�{V���GAv����6�\;������ﾯ��M�-:1 i��m��i����x�=Ċ;1�n���)��"�f���n����Y486��1��;�X�pҥP�kT��&4vm*Hg-�g2���r�][�c��0�!�4�&�;����w���<�~o�u�N� q����;Y9t�y�ݮ)�7V�x����ƣ�����|\���9��Su�t9�aL���'2Ҥ��%s������koˡ J1a>�f�{�����W>�F�9�Ź�d�
��Սu'�Y��-l�m#�hE!�-�\����1}Ҵ�s!��<*LW$���IŻ�
�;�Z�FOE\D�FB-�LN���t�ӥ��Y��o+UpӼ��m�8I�YY<���S�x���Dt�e�N�S��wRF�'�.�;��9��}1Y��NjҾ�۝;v�:�B�j����:�d:�*�r�2jY<�/ITs�B������[�3��x�=\�p��2�Ӵ�'��ڶ0������UL���%s]DE�p����qܞ`��^힖��-H�����8��z
F��T�w+5ծ�ñt��I�E�K�6ø��Z�{��r��L`�a�AiuᓬQk0��Y��W%&��_G�u1�]bή;�f��I����I!�%��81���.�o=��$���U��G�C�����t\��s�n+*��<�G�٘��/�\5&S,�F5�m_�qη��u`�Nի���X�Q�����KF:	}^g�_1�R�:����̰q�6{�0�!�u�`�5��QJ�ͺg�DSj��}���v�!,���Z��=����ei����S1g��|js�1%+$ʱ��#��Ys�:�q������*�����6�J�^Ι�r+��	6gke�Ѯ#Z=�N�oTu��.�P4�)ũ-��D
T���,��-���[�Wh罗q>7�Qz~��<9If6� ��F>dm�s�L����ڍ�snI�jV���6cDP����mX�9����c��0�i��ڇ��eÚF`��+yQ銠���d^�i�ZA�3ԣ!&��Qe2�b1�k�]\8�M�pM�H�y*�N��`A���y��u(�(�F�Py#�����D*Fz&-�u����� �?eG>��HUh��u=k;R�zd�V�\F�.�z`={!����	��S?���U������UC1=`w��W�࠿4v�ߍN�T�
c`n�,�7J��F��ͬ�I�ttcT���n�1�x�Sa\�1�uҜ������/���{&y�Y*I���`^[�.�vR.u�<� ����6+�s�}&&���M��M<ڿ�r�G�uµ�ﾈ����9��g�R4~������L��`cB���"/�'hM��+��Y��������h"�0U8n��O-�mUѸ��W��K���_ǩA��g�*6� +7�f	���y������M��k�l4m^]k��rV��`r7A�}��xe�f���i��e����5DV�|Z���b�M�Ϝ}	�*�Jf���p�a���̭j�%Y.�w�RT�j�k���뇪�4z�(�#i���]}L;�Tq���<T��Z��c>uN��cH)����t�xm�uc{�F/s+E� ]�A�BD>(I�˿[�.�����h���m�{���Xd7|��q�����é�p���dR�J�5	Y+��^�T�3�{J��5�*V\ᚡ�Yl�h�S��o��)c�T�hc<IӴ���ޤ�-,oJ�����}J��#Y��lg����������pً���7:���{�/qś�W��8�U�9�u��0���jF��ڕ�-�]�fQ�ӷ$����+��z�U_v����v�m1�p�X�`&f�M�APUo��V�T;W�)np|"��+Z���]��,v�JDN�l���S+�����@���[���2�p��2&UĚ���u�\Vu7X���b苇dחg`��%AE�[�2���G�}���Тu�8�������(	����iH��f�q�|jg����71	�i32��>DnX�H�8��-j�I̴�Q�m�d+y���]=�՜����^�6�>*)�bș��Uӣ��q7��7Y�Q���C����S�3S�����q�%����ts���O��j�O�	-�~'��=�d�Q��+h��zK�~'ڑ[���q)5�gp��_z���5iT95	��^L��ªRf�����հ��м�3m%�ԥ-� �As�ݜ�0��7Ҹ�r}[j�E}jy�%� k_T5*c'���r���-RK��j�!y�p�闞P��<i��ӵ�&
����}&坍�W��һ�eU��z-Ap�¨*�e���&0*��Â��V���h``j�K������i�:��������~����n�3�*��n��z��\��{A�Q�r��^�V��RÍ{� 4�G8��7\�_��i׳�FUԋ��q;�Uv��?�d^oj�����t!c	�bC��"L^u�i�u��c~�s|�֩���7��x��U���ϝ, ��.~�-�m/e��Y�߶L�M��9'h�I.�f�P�H��"]�}��Y�[�=@#*9�I����^��&�pK�\L�r�C�s�zwf)6�}�D}��M&����_t!�XJȒK��/r� �u�a��k�>�]�睂���/S�S�
s-OF��ٜ�pe�e�Uq�똄��̸
��Y5�)Lzj���AOW�5/�Q��F�9[�<�l�4tz��&����A-���諩H�����4�`�*�Cr�U;f�1N	Jt=U��r'z)w����cDr�"���>���G<r�c\n�*`�ڝ��m��EF:�)$H1�8,�W=�C���d�,b�HOI`�įB�lznP�b�@�N���(|�oA8q	%�	ܴa}�F��3*V�}�T��&�&& �趨fr齺�}χ-ɘ�5�:�O�$�Q�*��uÉ��0S�Bj�SQ� �=��]?C�L5�aMY���l�`�cbn��k��:H�lCe|�+��w�3B`Q��R��Sx��8�d��D��
�;��]��x��a5����Nc�19�d����*(mVX�6�=J>�=��4���Z�5��R;��Ҵ�ju!�9�Rcg[��-������8|ū>ͧLW����:���F�Q����Y�j.$�j*�V��B/��8���}��G�;�*��7i�9�n����#@G�&r�ovr�c{���`�&)W�U�׆�Ȫݕt��fl)����At�;�r�ވ��������-����F�����yU�V�YD�x��/������������ل7��ݐ�ss����9����p!L�X�S���u ��2��l��O�yf%�*JA��Q��q�rD��Y�H`c+%��9�1�'C�L�ά/�Tè�N��8��<f.&�){z��g�����T�rdc �tC��l�Ҧ!�-Oˏ}������\���uK3[c���^�jm�:P?�~TY:9���[�T���N9���*�Jkއ烱[���G�W[\��=��?M��t�9q3�&~���8�=ԸЫ§��Ғ簺5w'.�/Z��<Y#ێ�#S�D,�V��f�j
v��K|D��[����C�����\�ޅ�d��j��Ӗ�dS�a���e� F�� ���IHG2��m^�K4�R>�������BA�����x���w��MN��rxk4g���z���E�?�������=�.�Y��/O��xr��k�]��z�����n�R�OxA�Eb�2*�ig�n��Y8NS�۩�g[=@�	���,�CK>=��Ş+<���\�I�u�
��{����{��͞���V�]\��rm5�9;5ҡ9$� Y�C.��+M*�]16��foL��+)�.��׵[6J݂mZѦ�}��״�6�ѹ2 �_� ��*���v�2ގ����0�iL���܌�֧DṕǞZKpmґ+��Eѡ]/e������q��]\;%;l�A7�#�nƄT-�^!�=�ͮ�NQ5��r���|PrG������Q
�����9׆����>��ڶ�'�k�d}z�[�"ӱ����9 �D��:�&>R�'�RwD�s��h��/�k��tYXa}�L������o�w!���~�J�/"���ǉczB!�Z��L�]�
��T��G���{�I�v!�쮽/Mu����mMQ_a`)�`iyՈt~���VA��*#}��o�M���oƫV�11�#�J��a�f��,w��`y������w���쭂oz"�ݴ��kp_^����[��Bt�����n��S0���ӊ�VS��r�0��.E�^��&^�f����Q�F����C�����PP������{�d1�U��Z�u\/�Fn�2�Ol`�� ����O�и(���@�W}�2���x&U�k�g2��u5�=�ӫfh��\�3�\��(�rI.
�{^���ţ���1e�+B)R�.]yk�* l�z�+���\�,�A�3�0��WQՕ3�jV�@�9�U$tH�b�(֞Ū���pǺnm�m���T�ҪXK����_}U�UWN���m�P@䫸�Uʾ��6w>�_$��]��������ՊGvf+SA��ޫ��\:���P	g����F�)ܦ���T���ϖ?���g� �SR�j�׼f�š��~߰�鯣L(Į�dGON��V��6b�cr'+GU�jr��ԓp*��&��԰�9�:���9(-V��U=<Ԗ_���L���SS*Kf�7�xN�7�i��QTW,�>���rt��s>���+�a�=)/L9FJ�q�'
䓗�\'#J��c�0�s����$e kƻI���[�9h���SԠx����[׫yOh'��_+����eNwIﱻ��ĳ��� %Bt�<�쫥[����i8J�	��\��������0�H��f,jS��d���a�d�Tn�b�"�[����Ԋ-Ň2h�����z�/A���C������ �qL�3B=$JJ{ٛ}���{^�/zW�Q��*�L���詆���+Or}[j�E}jy�&�t5����n\��MH݃q[��'WY�뤘M�Ǫ)soUa�p���f5�tWX٢"��b9�wv��GZ���Vv��W��ٸ�g����.i����J�����k
���PW)����%��}�"ǳ7�9�5�	��=%&���Ns.S������� Z�J��Q&~S���B(;70>ugD}g���!���ROn�ZgG���mdjL��_�K�����ٿ�w��@�f��x��^3�6�����֙sSLkz{��H"ņ�.�~�7¹���~Nժ�L����n��^���J��RY��$��jjpx'��8�@
�u Y�e��a�Oa�����(���u|2���l�RŽY�e���O�ZRY�Z'	=Y��?=ʐB]sXd��ދ]���d�y*5��3H����Fv��R�G��4z6e�VK,��)�������/�f�`o��rܾ��9��{��E���w��J����ȟEQ��Vw���4�`�`2�͵y����5fy�|���z�p�ʌ��Z�d,^�h�����W�%�Ϧc\W@�6��7�����i=c�*C3��GSUxͳ�A�0���,���s4��ŗ�F��}�]A7�=.]�+� ����Oj�Ҽ\p�-z��kT��ƃ�h8��Y`z��X�OQj�4h�جs:�m�&����D�!��:%#H����˻�|vϰ��v/s�F�޻ݼ�]Yq.�����N��[�}���F%�,�7U�du�u�E�Z;.�����EҦ��fs���,�X.tN8��[��������s�c�IV�"}���s�Oj%�w,���Ob��3� <agI}��
�[��~;����&��x�[�e]����5��}Q��G �����Vp��vbTU�Lu�:��j��z�`H@�,{�
j.�F��.��	�u=-Ѹ��8Cn',u�s�uv��y��K)7������!�U�z���ʼt/��WR.�{�hy�ȋ�"�y����*EɆ��4o��#]�UG��!�8	L}��B�t4�c��	�j��/0�s֞ͽ[����Fp���/���&B��nX�58>���H:Y=�2au�'t���7. ���.��T�+ξ�(�wk�2�X�uLE�t��:�t���0��������B�C�J��q~�0��C^TY��S�v�Δ��*a@!�4�|��ڮ���{�P"w�A����^J����8����^�'�Y�,KN���㚕R��u�����>%
�;X4߼{��$��M�uN����װاf�9�p��\1���/3���=}Z��Z]xQ��_�u�1է��r½;I	;�w6�����^yG�\lȴ�����L>���A�Vʧeao�Z��k��F���v)%7;xc�b2Lop�J��O��Gか�F��ORqīeK��(bK�l=մ���V��lV���8+�\�x�t����|Q����/
o{R�ϫk��2��2�Q�#���Ħ�[ľv�6m������Ԗ�^��[����d��k�Ԛ�1�߶�9�t4a|*Q6o������G��ז	�.�.�Q���q{5 �p�s�=�K��(t�ծ��!ab5bW ����fq�Y�j�މ��^��E�-l���H�F޽�k��C������+�.TIBnR���͹]W���1>=Љ�_�k\�G\lH���ζ�&��3Zͺ�>���.�_|ڳ�vŋ7��iLrH���Kt9>�S&��CQ�|S��*n����m�vy�9�q�m5�{m	O���e�[��s���=���/�g7-�m�%��16�:��sn���ǌ��+(1���1��^�_/���J"�/�V�{1mӔl�'�[��n4�vuE}}N�vl����!��A��jBe
v�F���z��<њ�-K��u�i����¹Ea>䝖�Ɲ��2��xA�؅R�Z�E�v��pjl�m�p.M��]���K�)���5w�0���q�2�,q��m%-�X��8���(!R�AW�l�jԢ2!��̲4��Vi�hR-]�]Z�8g>O0��V�;6�AƠR�K�*K�ރ-Ztŧ�T�+���ko+���y9q��u��`k�(��	ܙD��V���=6��r���?��qJ!^�q[ge�H�*>{)j��|�KD�ە(��(�����]�
��W+�,��;���y�>�y3F7�T�J���P�s�i|&��[:����مdj�m\X�v]���ݳl��!��2�!k���jʾ��T����)�Y{��ZQ��l����Ɵ����۹Wٞ�� �w,
�F������c*f�z��0�pEoM��'ҹ�'ݢ$a/�k�����IN��U{���	�$F�WU��u�s�m<L��
F+G�\�=�Xs���`=���^.�$Ouٙ�ɜ�T���ԁ��b�M2o��q5�[���.����nnD%�]^�D��wʲ�Ǜw��fk��x�J1���ꊧk[(.�"��u��;�Vp�v�V����yrG(m҈S����h��%m���5Ťق;ĭ�uʘ�WaQ:}v����
����S��I�:#s�E���*v�Ϛ�qG����wd�ɐ��r���WQj��nSY�PӀvZ4P�6@�ȎRW͸4η�[)+ l7� � wE�=�.��o,e=V�٭��Wg}%:;Kq0hޥ����0D��M7�Y��ţ�'v*��l�,��H�0f�@J1{N��6h2z����p�0��u7�Y�(��4���Aqp8�������?{����4�JX%+���0�"�23cF��H��2B.]�e&#FL�IBX002��aI
LQ(��,�$�f$I�,�"C3h�d��2�Bl)F������@�Q��44Q�2# ,�Q�@E)H� �,�L�(%��dd���I �4#2H��(�I1$LH������4��$*4�24i�����B�4H�D�A�l �DH��2h�,�)DI��hҙ	K�@Ċ�b!�&��(��&$��,�
L�JE1*,A$"A������y�����;��Ja���'�u�xH��ܮ�%�}706��vg[�a�rYlӫ|[�u�XGu�ю�qk����}��|V��$�;������S�7m;�cE��ExT���t��Kk�8�a�Dަ��"��uݝ�Ě5�\"��*�:B/���N�5�g8�.ʔn,�����1�^���g�I�/�~[�h��N�Ggȷz25��q��[i��M�n+f��ci� ��L�S�;���_k{ݪ䭬��6���|^�˸�n���Aj�����@Xm쑝3�F?���_�����_gs�ޤ�S�I�|XKa��*�Ս㔚���c���L1�W{.�@&\m�վ�`�Kݼ�W�������\H"�Q���!.��t6S(B|{W�N�1b�J��"e�c�ʥ]h�f0Cn`�êfE|�J/����Q�g�aNUᒇ/xg�ѻ���w�ha'�m��c ��� R'�?�}˝'�+���%S��O�tyԇ�1{�U�Y��������#IN����Ň�?TG%L���\O�'PDLqD�!i��:�u��^ZI��U�0�R��"+f�ͨb:#S�c"Uto  �`ap�hC��dOi�!!suTÊ$�����{]щ:�$/T�];�֎�󠸥�4�y��gr�ۺǻ��d��
U��y��R�3Wn�Y}O`j����b�e���Kz��ޱt&�!scw��w���7�h{��q����UU�}����.�S%��Q��/:9Q97j���]��5�7�$e�ު���'��}*=�Lړ'GN��i�'p	�3�3�a���|pyF�|i��J���\2�5!�b�iГҫ��=M�3�.C��Y*.G�H�JE�HzBxyx��P	� K�w�i��9�@�v3�2ө�g"�s1�;�0�;^�и(���@���Pf��C*�蹄�
M�ke�kY&g/��َm;L��V��-�6WV��!=���kq��#񶌾�Z8�u���l���"�ʥ 5�d}�{����m��T�^pxCk��m�2��,��ۂd��ф�>G<Y^:F�G������O�,��w����cn�[5�M.�iBxR�.�p�,)+K	��#hKz�L-Cu2�*zW�ӗ��U[�wRxV>|㚊� F�mm�M"�P<r: ���O2�᫸�u��x�?y�Q��;�/;8�*M�v��r4���>�aQ%j���	��!���
�v�V^����w��]�����ɏ��t�7��(��l7�
�ءN���'r�{���݌�8�q�Ve;���\���~6F=�g��@k7qf&��i�c�5mn�}d��*���sW|,f%��]f1
��
Ţ���η�o6��FB魥���><��� �a2#��!�%5Xw���']��u|%��!��D��:LM�$V��,�������QS����j�#rj��-�&.����h�q51ٛ\w�sb֮Y�ۦS�#�˒&{����ު��Ѩ˄����p/#��4_��]�4j���=���(�2�Y5Wm�}��z���O�h4�F�g���Ʋ���]�k�R7�?wW�2��{����IZ���qAN���ڭ���菬�q�P�Jf'�~|�嶬kN2�MfqOȚ�����
��¨*�eZ��B������q�*˥�YQR�Y���-t|��+^��h���{q˝agϫ��;�b��N� J���w
���aZ��r�9ݯ}���ȸ.1[ n)�9gQ��X���m��>}�r�y H9�@{�X )�K��PT �	O�nc'�<@`
Q�T�*@�\��k�5�ڱ�<�~.������,L�Q	mV;�N�c��X�`v���v�\�)͔���-��vG�S��nd��uWDDf������.c�d3F���Vu�z������:'��vҬO��T�<�?<8!��{bh�����aq������Π����R��n���J۷����S��<�3�n�a��\��S�
ܲ��}Z3It�p���=])~������������M�xuZ8.�"M"`�	h릗����#O9��C�5(��T[����VH b�[�1gD�Te!V��d,OR*��l�!
�g��빔H\Ϋbc���1��'�M��_�Ӵ>�p�ϋ�M\>��H2F$��&��H�Y#�wC�V<s�z���v5FuS��!uH���j����QT�h�C��%���i�3r{d��X���`:&��O�-=��-�p����N�q7�`�s(JU�op��n�Z�Ӗ�1z��!� ���=Ʈ��@��t��}�'I.pCe������b]�GR ���Sb%q�S�@�!3�����k9u�Hzs��Tܾ}:�ʧ���'�^��ʱPz���>Ϩy�������ҫ�O]x�^U�kdKLӵ�1Q=oC�EB�2zF�<*LSi٣'1��Ȩ�v@��������D���Y��C�#2�۱��T���6��_k���U	��j�-o�@�^&:���w��߮j����1)��K��B�h��@�޾u1��������caiઇ��U�i�m�r�kHe^�lC�`�T���ol�� �ԼU�@��[�J�&�w��ck,
�gr�eZhv�.S�����T���&�Z�����rF�s�����>���ˤ�J��T�?zT�3Ǆ=��4\��/�uLE�t�ϝE����L8�Y�s�M�A���]���X���·�n����%N��s;�}������J�f7찼��U���Ĺw�ғ��e�m~8"�x0���+�e���9�U/�z]{9��>'9��SN?pR0]�ߗ�50j��ױ�ח����e�W�;'��ZN��䲥9�E�/'z��!���(�v��2���{�8����:]P�
��\-�3���b;E<I�oD�q�Ʈ\VUȣ�l��]|E�t�[r����pk ろtg8*�*�������o�`$�,�z%�7��γE:�����w�5��c�����M�N�����r����(0�!��n���K�8��k1�[5ȭ�e�K2��T���Ԗ+S��
��������j�tnZ��6}��y�9ߤ�$)�"��5�Lv�CXs=m�&W����.��k���zuN���R������\�"�J"�^d*]��Z{ǅJ�YΎ	��A��n�I�E��n���:�fhZ�m�Ϣa�܄' 4�6�����_W#x�lVQ�X����t�D�Kk�|+m��[��}�t�-���+���﫜�Si}�l*qΤWZb�U�[�5�s�3��7G{^L�q_�"  MO]��o
E����J�g.HQ��^o�U�/����B�����rmzҭ[Ҧ��y�2b�NU����g�Ki.��Z%Xu�"�&㌩; T��J����1�y^M����rJZ:K�+�Wt��kW!�}3��T�y�3��ύ��P�1 R�z�{xy���=�I|���v�oZ���<�K��S�cUto !Pܰ4�j�Z��������_-v��4�-��H]����1ǘ��R��n��sı�:��2�tE�yU]��="O���]��y3�����b��xyh��N�)8s�VJd������m�`��pҎ]�c����i1�ϭ�5�,f�zޭ9�-ڥ}EbQ��䃎�^�v���&�}/W77��{*�dr�U���\�kM��\�2��nz���V'�T�齹]�i�Tgaڊc���'U<78��>~kك�7�㵋���!�1�^�nE��y�?'@���ַfPi���2��O���4!Ѭ�GL��x��F�n��}��rKݛ�$�j'O<Q����>��q��v�J���{����e5�]��F�a|�5��� �F�d�u�d�u�pɌ)M���\�Ў�?/O�B�}��zi?�����cu�B��I�}\�����6�X�-�F8k.1��H���B����)������d�?ʢJ^4Ή�Y&�Ryy��^�|�$r�I#/\&;m����Q#���IP`w3�嵍l\ڬò9F56�q����_Ů��Q�3��{R��}�0a����
K�2ztم-s����-�p�܄�EE�2��(�=�U7� ���CV�Z��H���ȳs����*�1q���J�|�6�Boa�<�wvaZ��K@fY�
�@�RyvVjx��v�&�;�7@�_k͗k��ǲ�+���ʱ%=".�����qj�[jg%����"{o��f.R�9����������6+�`;U=�qk��[ܒ���E�P1�͆Ҏ�`d�8��u���/��5ٽc� Z��f*�y�`��s��6�j3�����,%��!P��t���XCܱ�-|q1V�3�GL�5蛸�1�9\,U��P����!8�s͑n��gS���Z1�3��b��gPk{~po��[cTD��ji\�5�Ӯ��7��uH�e0iFB�q�ٿ}�G�EV�t:h�f��n�r��s�ֵ�5�����Uf��{(2������������q�wC%���Q1�ӸS/Q�o��u�z��*�ţ~RJ|k��zx7~�����G>����;o=�g��.;a�n�'4d���&M��t^-��
6�	��Sï��w��=_m(j��U���7�8��vv��^Ә_l�x3-��g�#9�D�79UDI}����N��8<�fE(�zH��'C�2p8���6������m����|Wϑ��4���\�v*���E5��k�O��}��n#\5��ji�j���IPd��d��Y��J�oawm�A��ޚ-<j��qz��ʅ)T
	Mt�`�'�+W�r~�
]�Y�gW؟��u�v�S��<g$9�U��Vk�Y�_��]!R���|�ub��P�[y񩚙9&[t���3�/��U��8�;��{oq�U۟[(w5�5�?R��2mb(^{x�[r���'j��h���-�n�3̃z�Y���W,J4�]n۩�H̜����.��"���n�n�r�b2�kW�4� �����mfQ��DG��3��H2'"gB��t��AK�S��۹��|r����Oʸ����E�ˎz�b�u0�9j���7����Y;ƻ�ݗ��O`�p�)��߹&&�Mƻ��']�lR��Frx ޱ��Ҫ���S���潭Uj�u5����cW+]�:�^UD�5yBĵ��R�;(�]OfTO=}��k���s�׉�=ol�CyF� K8>��7g��=['@�q�/���1��o��y��}�\��2�\5��W@���Nt���Jv�A�/�f�*f�3��Q79P'�:�|�E9�F�y��3�*{p��	��k{*�ds��Zc��z� K�;�ⱈ��mY�F9��T6�齹]��.�;�1�PU���"o��M�W�Ӟ�Qݵ�nd5���-��e��\K������.���ۿ7��sn���F����N�͏+�����k��<���4����H����Gk%w��z�9X�C]��M^�tȻ�ݥvo�
#��4Ξ��.���Js�s��7R�z�`��u#�e�y������؋wR���0i*�;�[�M�4�No6������^���n���߾�	n-��޴��p�_��mBi����L���M,������g����O]#�.����.Zk�ˆ�[�L�'s5v�/v��*)u̡/�:�C���t�P`$�DIZ��)���pq%��m��ޥ
���������3�]�vA`%��jk2r�Ǩ�v��g��N��l���שc9��M��,�"�h�wa)2��Z�bN+�;��>X���桾C7ì{)W.*:�z�.���d�]�]�9,�SS|��;�֋�ꚎI�pˌwdL'D,����&A��ś����I��|6�
�˜oj��[Z�;��M���g®�d��^=���tX�Th^}޹�Z�?[P�?c��l�:�����#n�U�2��2���_Bm���/��go���#����c�>��b������h�<���Y���G�fx]*-���h�Ӣ��6��B�����*�ю�8�W��c�|{HU��(>,
�jX�����]k�d�XX��wWI�X6�(t�ò�.��e:-SN�ȷj7��� n݇��%cK��4iq�2�֮J��w��3!C7{W|���F�4	��X�i���\�k*'ȝ�>���������|Bϊ������fetf�,t�[���)���9�	�i����jXnT�X��C{@\��)e��y��8cӦ�#<����f�ٔ������p i�N[r͍���
�8�fP��t͑�XM��F'd֤S� �ѣ���m�D�O�Q8�*�R�X�W1)M��fm�@���>��<���.%�}�6WT��c"t5&Wa|9]B�V��d��p�E�v��T��Âf+�&��!�-m鈮��+Q3�&�e��H��K-YtNԬP�+X���.�o�<:��b�`Rvq�[�-����4S�(�$��C������m���zc쭓�@l������P���A��L�zx����]��t�ԧr�;��p���P ���T4�*,�	4:��b���A��&�BT=� vN�o9�`�|���4㲤��e�5�l��&H`�J�f�����w���^�X���uz7a�R����s/�1هA�i�:Q��qش:����z2c6{m���¶���z�;=m���4�2ކNR��+����$tұ��v��#��Q�u&u�;qg-N�9�β8uj��&@
�ҕΣM��:I���hlm�:�n�O8W@�Uev�`��� �Q�qP f������v2!���/�dJ��4�U+�#EmG�4ն�A���Iu����j������C�	���iWl�2JU.��\���MU�wi�-�q)Z�������}��#��,�}��+��P��w\f����Gj^��&���ik�7����)�;��C+�Ñڸ�m+�����"A������4>��Ѳ��5�؜�6Q@ȳ�u]��򅦀TᬇWBw�	�VJY9�ؗ�0�z:݁��c�0��_6+:�IR`�;�j|/sm���#:^=+�AW�[,3�x��{]EC۱���㋌3+1�B�Н*�@�m���+N�LR4��ˬ"�2Pd+n��5:��u8�"���;��}�s�c�Y)�V[սM�S����KP��������퇢U��$Ыu�R�5�&I#��+:�2�Y����+[�R����I�]c�w���k"1\WLS#/6m�Őͦ����v���V���X��5��ũ9��
���P��	sYF�kYc3JX8\h
}��.�Ji�۳��Y��8u�v�j����dZ�Z���f�t�4�Y$�Oe�uF򶯜F��P�:%�o�p���Z�P���e�ȳk���of�1)`�o�l��;@�qQ� P �@|���@�M�A&I��I4�	��Ji� �&,S�&��� $�!IE��Pb(�CɒP��M*d�J���CKA�i0"�aB#Fa$�B&	&Q��I��`#E"fQ� FI( hHH2!�P��2���&HAQ6I�d��1L#dL�I4��4�"42aBY�0�
d���J��4Fؤ�%�,L���
#PI��Ř%�$H),�a��!,A� 
L ���AQXa��$�A�I�l(|�gR6��ά�/R`^�P6%�j�h�.���Wi��J��S^����}ݪ�wWm��i�U�j�(N���~��>���;���*�D9����k��秊���G{*��8���֤�������	BxNL���6�r�;S)�^-noϷ�.�W!�s�i�7��o3V��������z`Q�|�*Sa̝��#H�'̅�o[wG��.ed�I�3(-P/���F҄�L�q���7��|_=������9}�����7eTV���jA�Q_l�+~Z�_ѥ��p�	�-�����ޛ�)�r+ܬ�}�Q�{b)�5�Cӈ���g�.�k*q;im,x��S\���=k�|��%P(t�|�J�������ɖr����(������p�5ٮ+޶}�՗ʧ�`�V��<��oOB�tک굼�k2 <�O��i\z�!=�_[c*�?"�z\��[h�����U���f����6�1�4�o��m
���c�[odٯ��YН�#���&M�*��%�A��Vݩ|�M�|odP��Y5i+{$���-S���WO/2�'���Ｗ�=��;�5����z_EXg:�K4���ƶk�3Ϳ�X�35�NrL�N�&v����ӷ�b"�k\T�m�Kg${�#6y�w&��'ѥ_�4Yz槗m^�zѽ�.sP���\�4���`V�cI@q;Cb�uCS��!� �Q�Jܚ��q�j5=y��.s��	��.n\7���k����vD���Sه�����yZZǭn'}�-�W�Ӯ�N�x��'���dk�b�sVn"+�'��n)�%��y���V�c�^�-q�g����}�*�U��A��"�#�5�19��{8e�_>5�t����;춝��^���W�6�^��v��y�8����X*r�O>љP]��_M�T@��\aQ1|�W�-6ŧo��G�'y��z�(0��}������X;�.z�iCW�¨�ز��2O`�V8I�[ ��q��ٷ:��dRd�u�6�+P�f��D���On�NĚ9���D[����DKO� �����]��>�3�O{�׹:�5A,�!O,�q�Pވ�v�b��;�&{f
�Vf���	E��=�/�LӖO�n�COV�W���tܺyXk2fK+9��ö��'��H��#wX�f��(�j��=f�]��7;V�՜��"_1�'��+���천���놭c���i薴P��.�\W8ޖ����2��|"���ToHi��]�\g[�z�)�*7��/_j�P3,������|֋�o5���1>5[�O�����O6{�GD�X�S�Q�%�AKE\�"ί�q����$hR){��U+�Mo!v6�)�(�%*���O���]��@����3H�C�\8��Kc�2�ޚm�vͰ�,���1Ԏ�Πu��f�#kB�j��jqJE�U6�kS.��I��q��,��tD� ���٣�MmJЏ7�Qķ{=BI�sV��j�SKa'SQi�4ہ��YU���Ŧ����QH;ږ-�N�[p�Y5�������e�T�z'ޯ�چ�ز�1���yщF��)����Bc&�C3��F�`��'y���_%�	OQdN����q�%갍�^����(�ܾ�X�u-8g�i�c��rq���i�br���t��F����(:2��708+$���w"��R�V*��a��0Z��y�ռ`���ͳլU+���36�ńƦa��}+@��͹�ָw�-��Л*d���Bt:���k�H�w�eq�F��	��£�64����3ѝ������C"%��mo[[ٺ;�����9a1���S��q�
���3�q\ចQ��Q�6.7�+�nٵς�����5�v�Y�H�<�	f���ruԥ_�]+�ب�e�6�\g��r���4x��������O�Ӏ_�'i�qIR�-��8k.1��M=2�FE�zJSך�:RH�J$c|����!.ߺ躉KMAI��Cݳ�̆*]�u
�&V���B����P���I���+���J|f�*``� �my�j,�������ͨx�S�g�B������TMfF]iI�A���Ɯ4�n.#�V�X�`���Y�D)�����������Jk2k&��z\K�[�u��TG>j�|�h+"aJ3�Ϣ8�.�ވ��Y�W<.f@�c=����g^Ҋ�sM1;�hemwzH��k`����f��đ}�rdSn�Wv=R���R���.s��\�}ݏ�oc7�f�ͩ�A����|������Nwx�u��/xL<��B�.�+uqK�쌶�Ƿ����޴[}3��0�q��,��A��I�{y|�[��B��A@܍�V�\Nsڼյ����3I�Ǚ����sJ��7�X{�[�J]���s͚����v��T�|;�\�ޛ���������S�����~^��V|�,>�����b�Ek=�F�j���6I󚙙���UG����\PGz�48%6�}�N�`1f��Un�5s;��o�N&#-s�2�-F~����O~�G9d�$���b�6�\|�I�}�4*����mVT}~�E��iRl\:on%v�]9�.��q��~�R����޷�ը<���4��alWؓ{�So��޻eT���%j��7��z�l���5Q�_9�>�_Q����+�5���oN>g�A��&�\��V��?rB��>D$�����gLe꿎u*tܘ5��]3D�$��y\}ݭ��-���n5&׵Q���~zί^{��GY��ˣۧΒ5ɲ�`��u�_��7��⿌$3� kBAg.	,��u�i5:��ιh�+�6���*y�.N�%���m�K�϶���8*FE�:al���M�.kn�ޅ��`�����f�e�"�k����&gi)��>5[�K�������_

{�����h�J��?zȶ��}�>w�gTb}�[Jý[�le9f�8���$���ޢ��IHq˵�j����jus�V�#��_�;��A�[��q��dϗ�^�H�@�u#(���*�j'�m\o'_kG).r{NpP9C��Z�t���:E�ĩD㖪獳�"��/�Jq_d��}�y��v2�E�NcMT��6�]�9Z�U8EB�X��ҙ�y�ת���y�rh"�*�&��]ZI��؜2�A��qѧ�k?\T����������V%я6�[�K*y����ѹX���y�[]�ݚAٝ`
G�^��*N8��;��Ψ�{R^�Qі�D�G�o����j�3�2b�V�F�1�XPc+����":`��Yf��p���V�)ٲ�ۡ�#Ӷ3�PN$��sn���~��W ��C�V��R�1���T�L9oI;{�@�+���h�	�D=������`�vs�z�z�E\m�Y%^�knc�PkqI�uHn�{�}��ª�8�b�j�1�TM��]-62��w�-�B6[�Ӯ0Y���Lע{\�Y�g�9a=�=�d�F��7������B��{��:�M�����H��Gml�X��)�<�Q(����]��'U89w�}J�Kb��cmꖟ_��c��TE 6b
�%]�9{�wz��q/�i�q���u)Q���޸k/-���-h���|���,�����Z����'��dR��zt���ƻ\^��]��ɗ8q�a���Р�6$cs�*�W�y�ςάO�����;�X�-��B��퍎P(��6r�r�w�w�������|}�D!�c��Z����ޤ-Mc�;|��	��t�t�᠔�j'�n�Y;�g�TSI�[�A�ή\m��S|f�p�2�Ҏ�·]&+���m�5�#�Z�t]��)0]*WR�k�Q�*g-�jC]iL��s�r�h�g)�gw^lU�$��CK:�<{�ў>cǛ�;�F���PK�I�y\r�2ǉ:���H^|U�ԏp����4���Ǵ�ذvk�xc�c\se"���&s�w�<�K}�qܶ�S-���I��Mƻ#\�~�-^V��5��/8�RϨ�l?}~3�]�N'�q���UZ��u5�#M�Me`�	j�Z*�-�V	٩!�"�jgTK�<��Gs�ɷ����'���hT�Hu7���ͮ�g��^ݯW;7�iڞ5m�^���s�kY�l�͢OC�
�f<��M���v�>t:���(�GxfTq�Y���@���Q��Kv����أ�����ȗ����moT4�?O[w�U�����%/�ӽ�tu��&&�,:�a�$ظt�ܮݴ�o>~�[f��@v�^f���j0b���sju�W]+�ثp�_ͷ������K�j7%3�y�b�d�Q�4�)�����'��'i�qIR��ۇ�j;3n¡�+2�n�s�!uԥL�:���?ʢJ]q�Eԥ��O�뾧��<���vn	�3����K����.��:g����C�2Zr�m)���+p�d��f���\ՙ7�@��nY=�p�]l[���.úG-���&]�U��4T�!��Χ	��u�3����O5h����+��$ַHjJ��_�z��>w�E�(w|� �0b���嵜� �^L��U�uN������8t�98ͨx�2�B!O��wL�d��z��٤�m�%Vgv��8�1�u�SJýI���&��9e �����|��rf�/1-x���m�����u��W>j��C6��"T���qQY�J媔�� �p*��'�I��[��E�7�<�2��cvOj޽���Z��&e<�v+Ԏ�j�}a����w~�=:}���H��e-�ʀ9	���w0�q�����<��vD��_T�ʜZ�7���5�ܛ��t(TM�.�����Q�����Fb؛x'q�q�P��o�>H����M�F�&�y�8���z��bk�)�驊S�m�y}7�\J����2�Le�v�Sc){z_��Ϳ�6cg+_R���0��s��q�Y�e�֩�*�f��ǒ��D	ܷ���VnU������22���f
=8v�wu�p�*Ů׽`�܎�u��'eβuk�O�H�r�
�!�/&��ĩqw]�)'p�z5AR��9)�eu��ps�C�� ��ސ���fK��}V��v��W��(�<T��Y�����,�e�9	"a�W�N��eUᐇ�v��C�*�ǿ-�!C�-��I���&a���I��"k��h���]����aͬ{Ke	�Ű��=U|c76z�����6}]�>����oz�P�@n|T�D����@�H�y/�O8
�8�F�KTk�{p�5�B΋|��%Q�LwϤ��v+�]->���^�<���6׾�{�=�6}�	c]�k���T9J�PK�7"�����)�Ϗ{�^\n�ӓ��>�}�[J�;չ	ld�9WS�h�}X�N���1}�6-��\��_b㜚J|�Ck"oR�{��"r&t.Y�(3� �_�sQ˶��Q� 
+������x7�Y7/���7���(�C`'�:��&���8�qʑ�y�x4�%&å��,�[D�;Y�(q5:�(�����B��/9��Tμۮ���!Kus��F��¶ು9-oU�v�28;�kC�+]|X!���p�u/C�V�<L�*�lV�*��^��&ꈪ������g:�]L�L�F]�����[�)��bv"�i=v��]SD��ꋳ@o>�Q��B%�A�2�S{*l
�^�� �4 N�g���<as�n�HPv\��ɠ�h*�gX���i	]��9b=�P�
'7���6X�{�i6mDqꚆ�g����/T�i�#�VJǦ\OA���;ם��/�r�A�WMѡ}(Eu+��mݽ�I�6-�#lހ�����/�e�2�U<ѝ�Z�(WwH:��<����e��Ռ�HS���:O�
Y׌��Kv�sJ
���T#1-��!{J��������ݲ�k+�V���X⎈7#)����̥z7c����9F�W.�k^3��>��ܘ���?_ܠ�f��v�+`Y�.6U�^��/��D��G>��Es9̸wc@h�y`�����d� լG�֪���ɭ�C&ۘ���ځd��c`t���]<���n�.j��̨��݁�ж�*�*S��X7t`��&�$,�I(d�/�\�D��uh�o�(v(�զȰ�Ջ��xn,��0X
�2�l1В.�Z�t0�,����;�p���\��7���GȪ��H.�E��\�s��i@�S�:R���x֋]J��7s�w9�����N���Z�����|Vڽ�|�h�	*N�	�݂�;���}he���ŭf[��n2��-�a�W	�]:nU�Vk��ed���O���ҝƮ�s%�n�F9�ڜ�TR�.��	魈�Pd�qs�as:k����Aq�qon^��#Z؋��/,���c8S�:^��\W� G�����������ד*)�=�WX�V>V�dP�D�h�:�]է2[.�����I�KF�r�Z]`��1#�.���.<�3�S}۔�;�3��vBa.��wuػ%�����kq�g��u�Q��	��n��Ӌ62��-��0��U���N�:�[��NQ�e��f�16�e�~�;�iV�Z��Xm#�A��\�س�Ou��_gd�6%6n	f�3u�k�^j���
tg��
箍!8jw1^#Ș#9����X5����Y@8 *�b��[q��Ά����Z�]�pHrT�N3sz��y]��)B-�^M��=�b����PFﺵ]N��ϳ�I*-j�}��L���ʛټ��;
]46�aFU�s��,��mn��P��1H ����D�M�Vc=]E��@�Y[�Ն�Z�fw$�����2ډ�V�ڍ����������(Q{�.��wH�nR���+l���*�MODK�A�zje�0�NȲvY![y��5���A���.(!j����J�"�*ԝ�ת%��◻ȤL�W������6�M�^�0�*2o7��m)��w�FBR"M����d��b�[@4FI!2cd,�X�$H�%@C	�`(F��2�)5��dL�""PQ0��1�Ĕ͈�@bH̒L�0�&B�p��2��9�DB��,���a+�� ������6C`K�di�����6,32	��Tr�@�܃F,�H#@��QD�TblƌT;��l!X�mw��EL�d��I�D�A�S�X
H�P�[�1�LH���v�%�Ė4rwFf�\�7���޽��ߞ�N��,Z�E8(�x�0��
�u"eF��,��&���7�̇�=\u��%�GҀXZC�H���]���%v�%�EtfW�Z�!�SQk�-���Nk�9����71P"��*��<}*���K�ӫ�5mj�V���N��(;Q	�k�Y�E�uۀ��yX�K�R:Q��z�'�*yhۍ��r��s��\k���㹛qN�N�����}��!�'����շ���3�Le����s���ke�ơ(Z�N��{5r�t��݇�PF���:�>U791�T_.1*�:�v&u�>m�3ہĭ[�gtgY���쯊��w�\�m(jK���	�v�&�ɣ�¾m7�����۶�h�E 6C�XSk����bO-������_bt�Kb�-�X�z��·��tRv��%,C�A��敺��Y.ډ;��벪R�Z�ۍp�c��	��i���X�NS.];����ˢbY�#�Li,�WEԷ��O.ƻ#\gi�1����a�ǾK^�O�n��g*�|�U}��;Sb/&C`!-�c��^���ã���!�t^�-Y��h�>�a4�$���6�@w�e�)�yXe^����nY���Ѩ!��Zl\偻d���t�֫��� /�\�E����j\�9K�5��������\T�P�k2Ψ�O�Ao�7ն"2kU�Bj�&�_�޹Fa��&U��Ef�~��h��홋	^�n[�NI��{�ýo>�sBob�t��!u	J�h	��AbV�e�UkIB՘g���ʱ����S|�pDq����ʉ03�K�{g��ݸ�/jjoV�s΍L����䘞��k����"K{��2_M��x��3��uCn~+�/����3V�ڪ�����N�m��� �C�y38듅K��7�D�&}k��m���;}I�5��*��@w)�^Ӱ�Vu*&Sx7�*@��IQ��&}o-O���/C_`�m��(�̨fEUd���TʴO`�s��C��ͧH�GxfTr=��nr��NJ��ѯ�ɜ���!�����)��ȗ�������Yvr���*��|��������+�s+��W�������a~Ö��6���N�V^ ��e��!3`/5::U���H���e4��B��AÆVMn�R)E�I4cCC��6��C�u8������**��T��rJ�V��GKy2v&�hY�]8g'6���P���B:�9�*{�GH��Y�Q{�N�=�(��I�n���Wn����:�дOg���3(-gn~6����T%����ب�e��\K��Ê��s}��,S= ���W���yݓ�ʔ�w�[��5�#�L'�w(@�[�}�u��V�{�����E��Q�:�K�:貖���E	�W�|�%EMs��[�u��[(t�wϦ
�b5$�j6쩷�T.XNN�8������ۉ�k�o\�(�?w���家�J�M<�).��[��[�s��]�҇Z������Y�D'2q�}�<Z|od��@v���s���|r�9�P���A\�f��v�^5p��_bMGjL	UK�
*��l=s�k��;��֋����&�S��#��V4�=�I��?'DLsm�v��Nsڼյ�㝱{t�go/)�+&-˦ghj�2��Ux��X�ʽ��-�^&c��Oձ��ڬ���m���7��h��֒*DF0!�N\H����k�1��5���������˛x�>êh��S�h��g�B�֥O�\�	�}G�Sc8��+�����C9o�v%X����%r��sr�Qơ7�,�����O\ʫ]���~��go��\�%�mk\�q1]�r�Mki�^'�<�;q	�s�Y�t[��k	p9�uJw/i��9݅wq��rS�S/m��>�Տ6�Uf�5̺��U=��	oyګR�pa��u�Qі��Sa}/W_��f�4��6�8�����;^�����no�79Q%C�
6�&mRl\KoU�:ULn�V��(�v����;>�U�:��Ol�K��-_х��͝.�j�ݨo���V�:Iq|����Gm���ɞ_9�#��_Q��L�8�������,rs_̵��Q���i��C��@l�>P�}���i�)W�=�Y\v�INS��<������m[�i*:c�|ܹ�뭨���֚�[Y>޻�U��%�!�������uD[c)�HC(\d��u���{���D��4zg]4��*$9�v;�J�0�	�}՛s&.�Ht��{�U��&�J�c۩��rR�Wư��s*�M��;7(�-T$�ڤ�S�c��Ù�fz�������2�]�����s��ל5*�X9�u��b�[�>�*Lr�qk���.�ߢ�Oк��X�m�҇Z����GJ����Y0y�gr���<Q@s��jF��f�W=��o��������Ԩ�zrL~jM�T��ފm�T:fQg�J�����kMRsϻ�ݾ�t����'<s �2L��M|�����c��&�1�l�m��1Ԟ�WD�S�������g9"�̪i����j����mƻ��+]�r�}f!���8fgݫ��ڞ��[����mg%4�(��SL5'���z�7�(m'�Z��K��
)
��h���!���ԑ�Rt3:��̩�ou:ܬw�_\-p�;�B�gw:J��L#�]% ��LѮ������ؒ�e�(��i�B�z6��4	[�d���bD^9��վى�\��U_�߰�m����	\-G��]ۅƧ
@�A��!��u������CM\dr��< ���56�Rߜĳ��/��⚊ڽ1�W���`�\�C�uk�����[h���rW�ץ�rϟ��k��7v����c5�ᮚ�DW0���o�i��3ػI���9�%}�3CW�iF��{,�gfk���{�:�<O4����7S�ГȰ�jV�NU�r�b��or���G����k(?_��y�Oj��87g\W^��¥�bt�6:�5���'�̂���¶�cv�񃎫8���ٓǺK���ˈ�jOf�!ee
�+UV=q�/�9�/�sT�&4�+��%�4Zy4����p�-�ܵ��q50#��Z2�JP��~��2�	<���;КV�3{|#�
�E��pƺʨ`�WV�����5,W�{B!�)�y�8���&��,�sBoi�(qҕ@ѣ��p�w��Tֽ�n��^ir�V�'oM���7���mpD�SԎ�lWA��N�'�/���p4�k
�ռ�S.������c��6su����Ș
�t���(Ԑ�0;fT������*���<�Ww�ޮ n�^�P�o�r4���d�xJ���A9°�}[(d�Ʋ�L��9,��cS�ͼŰ�e:�R��U�wu�m�ƍ�������9;;?�k��r�X�z�����̀��a�D;�:mn^��{pb�Z��GR10���=����ZVmX�SԲR�E�L��g����}T�o,ŷ�*��߫^|�K��������]|Sc,d�8iB/$�5�_m��/iNv��Bs�Cx��&��Κ|Y���s[�z���#]��w�H�t]��~ʿ�<�TML��*^�~�Ҙ�܃�+�8�\��2��K���mC�ܪ9�]��\�Cs��fsm7��[�ٷ\.�.'���G$طM���ۄ�����I��)7UG$��ξ=s�;?y�b�!C�%���yۮV���Q������4dm�ު��@�q_T�
�*W[� g!��+S+$˷	��ͧ���P��9 B��U�O(��Ǐh�7�:�+)��K�=�}���F8[Qo��T�@���|�~*�Z�[��j'5Wwg(չ3;N�w��Ơ����n|�f��r��R��EV����*8+�k!�f�>���X�s�c�~�cK�[Q� y��)�ֻ�6�<����<L:k +��Kl7LdTV �=���nY��[W�	�sݫ�#yd��Z��*�7X���TK�ygrQ�h\9arT-�&�ʀ>X�Εv�X��7r��k_��RI�V�8�Z(f��[�g.�)��sy�63\��6e �ew)n4����� ��ή{���i��M�o�P͠�뮵4�ٗ��8�����0��Z���-sS˶��:֌���fFd���mb��Q�r�6v1ø� �?�Y[��/ݦ����t�Œ�V���5���L�\\6�]�:����+�����5#jrbʩ2//���m�z�����9:��18f����ByU��7�tVdp�2�z�#�g'�k9K*y���u��{�^�N9��w��2e^��j����vq�넒Dԑ��9��[g(��|��B����f�gN���	]�٫Yu5�W͟{E�2��ƭcGޗ��\��9-_��^�����G�=�2�=<�����o���7*�=��bߖ��?!��a� ��Ʉ5��o��,�E;���SR�Sj��CA�4s����rpX���δaOj�M��ð�l^ͻ�2^e _�h����r�5yn�r��Mu�e�2�v�q����
��DQۜ��d6��c9�V��^eo^w4u�I�n�|'k�I���v��ɞ��zZ}��;l�}H����z-�k��/�q.[��pk��?��VỸM�-<�-)w҄�͊�M��\��z�K��9�TUDOu�������eB|�JQ#���[���5���w*6�p~��3WZT��ޚ����ƻ\^������*��V5��.i��Pم�9(��T�Ψ���}����ukdd9=/i=�8йqG��v�=��u�����c��|���t'E�k�m
���C�P�F����kVv�=n]��:�OV\ϧ��y���p�
��1�l��U�.���[��p���{=�9Δ���������ی}�Y:��5ݲ�^j�{B8���F+���PD��i��[�i'=�#_&��ByEKR��%Yb�~��^�_Z���h���3�V�A�uj�5�
�gtNغE��r��2{MYJ�Z `�en�"uCE�]Y��5m�I��q�H���W�IǢ-�v�+A�=�-�J=�G�%��㈵�-��"8O]�X�q�屡�b�����7�ԫ���vTD�=���r��9}k\>1bsfU(� ���I�=�w ��l��}i��}i#oH�ќ�2�s,E���Z<ً����z۵�܏w�o���OР�N��U�j���j�/yP��:����99cb�?�J�!���u����ꌡ��>߄9V�,uO`b�/�$�2�E�7	^Q�1Q�7p齹[�p����L=��jr�K{�Z2{g����N�}��Tbt�0�*-CX�z�[ڃX��[�ɯ{W��KL�-p�D�Ij�W��M7v���p���fw��[�{��R]JT�9��'�]Pq���uޚ���\t"���/h��oNkp�I��Q����*�P(����~�O��ә�}5/=�i� ����`t���a����^3{Q�B���!���UV8��%�%�'vZ��nHu�Z9>h1g^Ր�$�����9�q����kYo!��b7zQ꽂X�]c�
ѧE��!-�=��V�d��V�PNwc�+@�E{\n�Y�;�J�1��>�v�o�b�#J�49&Kh5��Ͳ���l�D�и_M��Р�,Z��Xsm<��,�N�uNl��U3��0��WcC6.ν��,�9 5���e�P<1��\���^"PfkS��/+��ז�`:�;�\RU�B��h9Z�h�����	Envgq�9)9k�
x\=�3ok���+*��-,]�Id�q��6iArtWrr��������Vw��c�WZ(g$�&Y0pQ��������ȞKvQ�8�ya]5h.F�8>� �du���4��A#�	;iؼzg-4���T� a��+�Y�y�P���:���q��9�l[H��b�7�ªi��Fw���F�p]��N�ۊe��f@t��jW�4f+(*�]IkȠv%���؞��KG�d,�z�
\0S-����.�.��N�����'�5�d��e�7�[����Os�8�(���>�kz�y�T�ɪ��x��nr;�\/6ƞ�l�V�7�O��d��pq9XI��kH�v[.�nJ�{k�9wy0K�KZY�	GN�����9� <��!D�w0����T�%>�a��À�j�Jj	v����D
֭�.�Z�aN��z�����e1�a֨�ſt�p�}��1^��|.�bp�C��4�Qә�߻���	��y9�S�SxKe<#py90�0Vs8��ɀYzC8;��ӆr��
T7]Y%�`P��C�km��%CŶ�L�G�8Z:��W�(�'�Jl���Jmִ�p ����F�*o/o�vէ ����ac��Yh����.8�]��u@�t��X��yP|(n�M�1��G�%=|zAY�n��i���vv��[�T,��h�R^��]5Ve`[CZ��+bȻ^#��8���|�W����Q�;~+e�o�kz3T�V#�a�[���)|l�޹�ً�kEw�+C
<X�'G��r��n��+5St�T�u�NZ��ʙ����Xz�<����al�Y,gu�B1b3nX���=li��$-�r\�Έ�y�i��gYvo[�,�;�c�2���
%��1I�,��\��b(�&�[Ngh��14
{�t�f<n��ժ<a�*2�֤�gxӍXG�Ż:���B�U�9,�����bn,B�qu�Ŋ�8~B�n]L�3�;����馠�l�c�l�q���4�Y9�Ԯ����ȋ�뵃-1��yfh�9dN�M�Ax�Νj��޽�Her���Օ��5���y��ks�W�̮C�ɦ3����p�(H��v���s�����[Z��9���4Qw#P/��9H� ���=hueݚff��ޭ�W)��\�R�S�o��F�U���Y"� e0 I��b( ��I2I�Y��]r$��1E���n��Bi2m�6d��س,Dc�q��F-ȫ����ܣE�s�$�ݪ�FLQ˚�U�j��F�69�4���6$��;�9tBZ1�Q��N].l�-nnE�lQ�h���6˔h��
.��r]ݣ��i"�$�#E�E��F��wfƹ�uh�*����T�AIG#�6������6�t�nWw�QƊ�vk�b���V{��~��j�� *��3l��ŧ���I^\�yΆ�Q2r\&�+5��՞j���r���R��ػ�ncB�&8��2ĵ�/��ֹ�_���M�M�q�:R�[y��D��Ρ��5��m���No-������}ϝ|�����y���sT�Y����j�M{Ҋ^肽�Ӆ��Uӿgm�.���b�q��錯���+{z�5
k�0��y�5k>����\A~�|���/����]fꖾ�T�)dco*�]�??[��$(��7�*�/ÏS�w��
sm>]q��/$�CYUb�3����Fbٷ021�V�4��AM�N��r��S/m��dk����iS�n~\|�w�Lͬ��<�7f����KB��D�>w
e62^��o5���e��ש��DJͦ\jzL�	3Df:���*^|����ۉ]��WN�k�BM�k�̀[vUEhݢ�`��<��R�Vܗ(��_bzp{EnQG׼�G{]������ԛ�F��l�]KJ��Vw`�z�;e���}ڥ۵qV$����	=UmШ���8.��\4�V�us����^�V��#���b��ʘT��Q s�΅�:��Oka�)-�+�$��JQ�͇:"��g�o���O��3ʁ��GK|F%Hb1&r�����9�O]�G[��L�8Nˌki4����@��� T>����	=�jS�Pv�i"S�2�O8�>M���j�eGʒ�wϧ�7�t��mK�����U�%��X�%>4[��+}��g<f�JB4o�i�z�+�;/>��
�jͨɦ
�o��)��t7�*cvc`�5ݖ�^�R��`
�K֬|Y����0����a�u�{i�owD�L�mdL,c>b�X~߭
��ٵ�5���^���8dL�17�z����g'EM�,A6\?*�u��ce����k4�3��NS�Ľ]�����NX��Si�ڌO�~�tD���[��w�y`��'�ݴW���`<��<Ͼ饹�O���}�i��;����3µ���j�#X�^�(��Z�jm��@2�!e͊��n7�C��3EkM��䷲�감����m���}\��od���j���x��.\�2�|2wl��P�ؕʝi(�����}G8�Z\�;��-�e.σ��;�"�W9f���.�{jNI���Jlޘ�ES��>�qZ?%<�<��{q8���{���1[Wp�|i�'���L����	�Mά�k��L�-�\d�]�ü�N�ښ�q�c$)�H�U��X���~c��Tb��bo*���;BV`=��o'�Y0��j���yk�+ݶ1s�`?^����ՙ4Se�m7�M�����;��9���<�-�F�q�ͧ+��.��� ��Z�_�[�p��Bm��>�F�O-�.�������،Џ�����.ړ�fJȞ�5��z�4�u����O��IȎ?k]�Ҹq˽�V���Gp��gw5/�-�����k���S�}��{�+��!�=��ٹ�[�t�BZ#y�ೱ>��j�B���?^'�V�L+�M��ʈr8���+�ў�Gz{8\Mm�<�����x>m^��3ӌF���^� ����4Ш���}�z�j>ݪm�N�('~:uN8�_,�Te((4-}v��'�Mj9��Q�B��������>�2;A��ӳ9x.��{C�����+xӡ�[ŔV�0p��l�1���2�,ͬ����r���^������=M�;�=n�fФ��D:fQ��သ��q�ϙ��~�;�5�(b���P���x�T"�G!���$̒.9V�.N,ʬ�5&�en�ڍM�}SP�0[q����]EV����9{�u�&I���^�mZ9A���(��4��NMA�R�@��Q;����'p	NY��E-��R�*'����u����/�Z��/.�#���BH03����'���ys�ip^��v�x$���%��c�OW0-vz��r��Қ��-���/�暿L��p�jÜ}2�tlH������m����Ŧ�K����͛�s�ʂ��8�O3f���{����Qz}�1��p��0�+�I��7�nf�����Va��P>N���	੘�g�9�.�P�'J��ص_|�}q/�e����/7��"H��AXЏ�#�����nV�� �SThY���J���Jg�n��ׯWG�����\��3�ɧi�g2�i�m�ˋ�;���b��@	-�UeKjH}���
���]� p��o[�ݘ�@�\��4��r����8Luy�x����e	*�5X$5��rC��T�^�}e�:����Z��r�SM�[f���C���F�ʾ����/�%�8��3$Iz��u�OQdT�8h5��վ�[�Lwϧ⠄�������S=kjV�C͚r�4S����q�P�(�!O}�0X��%S���9�w;s����Z�>嘎ub��)��%�
���Y@+���\y1�MLX}ކ��|<�5==�����>j�|�h+�>	�������/��%Tlq��+�m��k��W�ru�_7�5������d���|��Y��dLBtD�!��+j�+s�紧��{��^g���(����O-�K�Qơ7��+]��t�[C/�"^aůYƖoLf2wZ��;fr��:�NO(�D5�Q����P�In�2;o����/m��D��D��m:����2|^��Z�p��]������\q��]�P���� m(),�(��L�6/S�R��r��`��]w������Y�%L���m+;4��%�\�yc)�T2��8����:�ުP�����܌.��7y��'p�^�N9�r7��ͧH�s�k3}�B��kJ���v�*8�,ʛ���:�g(��|��ld�]Cu��:}2�5��C������k���j����ms;�M�AP�����*M���{X��S�x6z�a���Q��s�8κ~3ց�t���[��zTY��cj\Cv�K)Z��\�2vX���V���?3@���#��]��V�P�UMLt:"�u�l栺�B�x��o��^�A������zs����b\���~��^�]TJtj#R{o�[q�n�8��6���|��yI+}3��3��[��j��̭��i���-�w-�-�%mj�\gT<g*�7V����ݞq�.@����֊�b��u�Ҹ�ky��j(�2�M�4�P�z�N�\C!Lw�O�A<�jus�F.9ɤ*�Rl6�&���Y��LaEv��ޚu��'`e��B��i�]if�h��`�J�b�e��g��I���c��A��h�$\!n��;�5KUq�������FE*�tnY�]�fl�H�6Vs�v�,����f�2RAa��vk�צK��S�6��ۆoECob�t���}A���O.ھ��l%�����E��e��j|�n1�W��nD����'6]�ԓ{�����)�T���륰�T��`�6�]��k�'Pف}��n��6�=�����h��>�o�%5�LتOWbpʇ��ByZ���fW��_3���#�5.I��~���IZpoԝq=��Lz��G����1�G9O���\���x�Vzz�����N��=�ʜ7�>'t���a�VW��s��� �����31�86�⑄�f��;2G�M�43M���U�m�tUvG��,KN�K�`< K^��A��¶�9%2�]'�^��Ӎ��ϭ�9'���3~�xA�>�G�<ױ�!�sq?n�9�ʉ��@�}�A�����N_���Q�q^W���Ш�7�E2I툙C�=��1fj���w��͝q=��g�1n�	���U��}^��<}�>����ϫ��ݟ�5�G����V~Et(��Q~e)v�y�q�F��H<PΥ 5��:�����Z?w!�(�`r�ͷ~l���P���z�u1�	]h5�lvӋ8��m�%��<�mR�u��D�i����9Յg�;�>�ܓ"TC�Ջ))԰���{�g�L�<.�ԼreK7�7V&���8gz=Ln}��?:�n�~���Er���ľDx鎊'�I~2��"E|vRS�y�A����GD���dy�y���Jj&�^z�ƤELk�u��t��.K5���Fa���q7��^/v :�F�_�ě�=��͓�V�s��&o��\w��p�o=�#o�LMD9��sG�Dķ\qh�$�j-�����P7�h�y�o��gӜ}����m���_��f�̒ѳRٳ�FAC)ۜ��<=���QUWx�W�����K��#1���Fߧȟ��x�C�\�$R,���\�dR13}{^��7dz3a̓Ǹ��c����T����R=q�o�d����|F�I�$r��1@����n���>�2O��}P2au���*%���}���1��1�߮�^?Ps=)vبsj������=4zG�	�Dy��2�O�U&X��
�[���/���~/����6�C��/�|u8�>�<Ԅk����O���\+ʑ������w#��ڲ[�J�߾7��*�O�c߇c �G-;�4FO=���p��Ur�i{֭���z���ZF+�-[��6�j�Q��_i<�����Qb���p�9��F�(�59�&����v7�2��ü�9T��P��oo��ִɡ:y��<A�t3�씌���H#�3�g��}hdz���:��5=�瑡��r�rǁ���6�^>���5��{���r��|j^��F��bj���������<��y�r�[ư�&t/�+m�f)
��_k�>���/	�����:,ר59����ׁNW�޺��dSW��>�$���h�P�iP����O�,�+�e�x�]L��t|=4�>�.1ǩ�����*'I�oA�kKq,��ފ���0����>$�U{�uEs�iwڥ˺؎^>�轌n��۫�
e��̬�cۇ=�P�#޶=�>��
��F�E�U�b�C����yw�)��] �з��5�KA6S�-Wa�?I��HJ�*#o�TÁD��R ����u�}/��gW��������5���ٓ>���X�r)�\M��֑����a�F��o�F��2��
E*�Ξ�[7"��{�]��.�U�� ҝ0�3�Σq�R"_���������7����~k=��1�`�ڔ��̲<x�Ls���<�Д�x�f|={�r:ו�1�yY����2_��Y�}���z0���t�,�Փ��ˆ��n4����H�xG%��-���s�/s�U���*�νY�a5��+H���S��;#w��[2h���#N��$iɌ�!����9�㣳��KNQ�2�T{�9mx2�ZC���:n�} �Q��Њ*_�W#�&c��Oa����7Y-t�}	S�:�����~�����³���d���<��4
���A�,��C�=s��NV���Ͼ޸|}�Y�>��)�����
.2q���g�@9�z�d�b��eH(�����g���n���R�)5*n;��$߷M�h�;����v�k��7���ܱ����K�����]�Y�}�S�ܣVWMo��DS�6�W��9�>��w�u5�1�~�^/{�pU�׼o�ٜ#/�~9K����3��/�O���}3��6tz���:�|NlF�`V�G�:���;^�eg��Xޘ�;�Q�jx�^S������?V����>Ng��ʁ?�b����pi�Z%�i�x�T�0^�q0�#0e�e^~�-��1>\o��C��?u!q�jx��|J@ó�z��z���t|&D-׭��7��}����,'<G3�NӖK�w�+�.ʑ��\�O�+ƌ��Q�"}e�.�w暟v��e��M�������|G������Ϝ�i���(�_)`��,�F.�x�~�W߳+)4�)q�F�kP�O^4���P�d̩�$�[q_s�PW7F cb�2\=��鹽������=�
J�
�gך"���f��YK��flLQU�"�yc ���iG��Hʽ�dB�(�G�&�9������D67�6~�WIh`�.Z?	d]f�`E��޹4ob�yi�k4ggk��l�m)Q���H�_U��t�4.XAwL���B��G9����ÞSW*L��ؓggiW�K��x���/�h\�+�=Քh��x�Jѩf�iC�K�8��ڜfD"L�{Q�ɶ����.t�U��;�����TW/��/�oP�����u΋�1�"�B��$�媵�*�>G��z#��$�F�+�ѻ��,t���Cq\l&Ċ�-s#�a�qΫ��E���V�B����YYk�j�b�Ķ��egd���V� s��Y�����z����Lʛ��]za��nJ�J�PN�s�����]z�N��4�f@W����7������d��=Mu���al(cCz�G)%xpV!ؘ���4Ld6y����(��5�D�*��av�T�*�y	>6���Bi�N��j��k9�vh���0%3q�tq���ܳj�)Gt��)J6��H+y�z����KqWrҶ���|+�j�Jۡ�P�֪��x�i;c����n�:u�9iB^�1M ��|�w28&B�t��}�H��i�fn�ցuq��^�I��[F����05��k��sA;}\�ђU�-�	�7�-l�>Gx-���9�����	�*<���&Rux�����f�GxQ<���s�.k�'h��q�7u8�w���Y�۴\uʅ�l+y��m�+��(�}[�}ӓV�>g�B;W��A>�ء3bBk�g,��l��G��:�]ɮ��̕��c/r��<�&2䤲fE�4�I�R��=w�v�V:�_تလIn+��Z2�y�Ƈ��IL������H��V�����+WB���|�:;��S��+zv;�v�e3o��"�ެvv}w�#Aݤ�:Y�<�`^$Ь�Rە�ϑ����~]oh�t����xԤ�"E�t��h񝏍�����p�Q���J���N��f�T���OT�hC�+1�pR�hvn��F�ću�»�6#י��Ls�v��]l@��������ͣ^Ei�y���5b�:[Q>4������K�^�fpҎf��mt���>\�_��@g�=JR*�_P颕�Z+
2�W����݃�����[�qƶ�
|+���������Ϯ�s�G��]&O��,F�h9f�A�2���$�X���݆���M��Z���8�����(�]p�He�ˮzٝ/e���S�z�D2t>�+�k�9�2hzp���ƈT��zr'�RWCG����+����X�u	)�u���
�o�ޭҢ�;�����jwwunV�sn\�*�ۛ�\9k��\���r�R�nm�h���Y��s;�ƃN��wF��7M�`*�76�&����k��r��h�c����j�:�lk�\�n���\��[���&ۛ��6���������"�E@mr��C��bэʊ�����;���5��:nnm�c�r4E���q7-r��sC��9λ��9�]�srw]����TV.��f�cq��#n&ܹt�rMp��%+�v���cn�t��79����������������Ό�9N��Og_����̙u[�P�B͎ۛ
�yH���Cr���V#�#�wN&�չb�B��Lv���-�E��;��2���Yu,�7V&�������o�3��p��.��Q�G�F�p��fO�S�Νɏ�ç�͎����|r��Bn}�CF7���x�<����us4�?E�{���\:�Q�;�.Op@^
e���8��
�5��C"}�ldg[7y��S��d�_��R�Cr@��>�����s�̖i��<LLJ�u�������z�H���~��@3s[u5��|�ȹ����^'��87�����_�&�ϦT:zH�}^�qJZ=v�3�L'�&��}��=cЬ���j:����������}��N�ɔY<6��*p7JlA�t���;��UR���.Z;gx�>��~�{Ϊ��r�L�{���q�̞0�O��-�α*��Q]�9�N\T�:."��~�oS�|�.D7�c5�+�}������:���'�t?bW��t�Ϯ���q�}P2a+Z�O��N����c��w��!z��25�����Q��Td�U��^��T=bk���Xus6r4�wn��	�0�'�D��qF�`
�s��^��'��hN��D�T0)��77��5^م�"�(2f��@lv�#��+�;$�ݰ��%g��m���.ڱ��'۷��"��6[�T۠��ິ�����2楤ݑQ}]����&9G�ը�6��4�����t8�ԫ��KRb�=�g�7I��43O}�ԅ�eH��K'v��<5ʡ�L�ة��U۲�h@8.�;3{��S����ȿT�����5t��ۮ>��B�T䞻�����
;�nK���r�b�ݾ������l�tϠ;���6��uz��=>��{m
Μ����'�F@mKub�\�/�fj�	D�o�iH���ayk��j8���x�/��<�+��ݐg8�n=)�-pp����H
�>�3g�~��2��#�%J��Y�,�7V&���8w���?u{w���~w�+}ږ�+p�)��u6�	K��j��|K+u#+e%9wP}>��|�X=><�{0��=Cls���
���އ�U���:�p.K5���Fa���zW�݀�5U~����{=�Φ����r�>��=��\8��=�#o�LK$�ϑ 74}$L�\���9Ts��%+�����5����O��Nq���v�~�����f��-�Rټp��K1'|���s�z%:b���L�퀧�7�F�o��~�p�>D��s����#���:�;+�GH��+�L^T�Xج}�k�r���x	=��7Z�Z��y��R� ���+F-v�Y���U���O{lp&l�8NmcU�@i�����6t��6.�-�����)W��7�H:���.0�a���7kyV��XY`D0Ú���jU�3�Z����)�/�*y��g�q��T�������Tc�o�d�?O�w�V%�p#w��W�{;�HW �c�9fI�E�&Avc>�koFV��ޖ7]U�~��u8��i6����D��6g�����ࡱ�ʐj:|J����;�׫t�/��%~%�+\�l�t�]���Rͼ�����{�CƖ}���ɡ��e�v���F�����<����=yM\tb�A9��t�ޟx�m���U^�sΣ���wP{^_�s�s�o�/l�S�/6}{��D�_y��:�l������wؼ�=�ex�r����:�����7��ɝ�*}^>u;��z9�d̯_�gFT	�����N���̰�w�n���s�]{ǲ���[0Wl�����o�G�z<lǽ�f�R�����S>F��ty}V�O�z��G�#H�
�A>���tw.�2q�W���q��2���'���U1u2�ꩉ[�X��5��>J�^�/:���g1�Lא��Kgs}@>�~�=����F�d�Fa����T;��i��6/�}샴�7e~L�����2���/?߬��m�D�qQ� ����-�bɚx)#aP�!�gT4G�Y�U�l�p ����ٯ����Թ��p�ͱ���5X�ԭ�}x/�h]t4��hY�vkf�9i�&�'q��.˛	8/��G
�Yܻ��ڎWV.�Sg�W����~�i�9>s����|n>�*#o�Tðl�_B���I`S��W���vno���J��@���+\��T}O��O�IӞ+��H������fY ���v8�N��o��ǅ��O���j�>�cX8�>����1�}�m��L�o޸=�����}���{0sp�z��&G��N�u0���MM��x����������V|G_��w�Ӿ���ֵo6�q9��_��`W��TM#.OX���=�*_W���o�*c��w#�r�gރ�6�0�9V��Y7�~��>���σ��f}Tʑ���)��P��}�v���]�n#�Cf�y�����O'"��,����{ή��?Po޿���X��eH(��� �|o㳁{z��}yx��V�z���,2�E��%/�meB��v�Dk��7��<�^��
'=��Ku�������X���H�O\VRqJ�Ǹ���=����<��)�޻�����*s@��s���=�ܗ
��*2��ӳ��(Áɹ8:*�;���[�Yꟳ��Ez��WA����3�ڊ3;=+*�A�Y}�����H���)D"����Sn�
����䜷mx��o%�x�ZK�p��l%s���U��4����}-K�7�7��f<�8i	���/GS�\�Hj����º��C0n��&�t�:��Di�ŧz�2����n���?+���+��sB���T2��ן�z�xt/�:�#M01:^2t�z�V�ռ<�G`����wM�J�����յ<nωJ��<5z��W����tlQ�pSPN��T�=�Ěz#�>vE�zW�����<�ԇ�/�r�R�qr�<jJ�L>��^��{=�U�{iu����#�;|o_�����
����{�םxv}9\�d��,{gf8�z�}]�Z�J�z�5Q�S>S஦|z��q�߸��������+���e��6j�s�R�_�Z�Ũ×> ��GAʌ�&����l�����"��Bn'޴4g�ﭣ�ޑ�]WS�r�ѵ�y��=r�kΫL8�Q�P@J��cž�/�Ҽ�w�gB���A�����T�`Q�R�]�R�A5���Ә�{�,UO��&�H�A�� �W���t�}��kls�tk�m�սՙS���	9.E{ܯ� �ԉ�G��d�C�������d�e@!�4���z����6xf{���f.�,ז��{�����sj�E?z�>χ���XC�reO�f{���ݵ�ضK��"\z��)L���n�����Xi.�=��,4��R�b�����Y�P��`;D*o|��|0TWH#+6�i��)��X�ޏ%��������`I`W3*aj����]5[׮﷌M�e5˹��l�����;`y 'X�]�eVz�JP�VW3�s���?mG�{����d�ސ7�:�_q�̓�b�p\��S�շ�GW�����`�k�踭�_���>7�;ˇ�߮ь��I����OT��T�C��Nz�z/�i�3���3���*�L5���tJs��wS�۽��sU������B�*d��͜��V%\o�E�W3gC'3���@��ⲽ��:�w"5[ /E�)�sK��ʶC�6W�z=T����ϗ�^���Cֵ���vx�2�����yN����;���㱉=�3��%z<i *1��
JnL���ۮ<�и�9'�������~`�����z*�s9v��q}^��*��ܸg#�}����N_��b�q�>U��B��$�e�Q�!G�S�h_�yਫ਼�'�����e����B\���Vq�x��P�z_��y�y�{�����L���B��x�����7jH<
E��T�s�R��7V&�����w������˕.߶7�	�<m��[�3lñrQ�|ITe�?�"��Jr#������"����[�glUל����Lp<b���7"�o��^,z�Ⱥ���
�jw�J��h���|�iP�n�4�F(�n������.�v�J��y.s��fa���J�ٛ���ӝS-�|g܁4���Y��j�q�T�3KK�mS��LD��<u�K/���7pr�"���Y-���VzP8z:�b�H�@À�$i^+@u�Ut���ׄ�]O��0��M|����K���|��N�'��Q~�bi̗5����H����GMzjcÝ��a���@� zR/v��u�1��~��A��x�zv���_q��s$�}�L��ӷt�zyqݐ���H)J�J���
_���^��_Ͼ��x�C������E]�yR�܄�P�IS�30�t�����	�+M�*|o��G��Wtb�߬ɖ:9\o�o.��#�^@�د��̓_"��0��O��kkֺ���c�9��`8������ݎ�(�8�{�PS7�����,w�d��Ī0���W�z�L����ʏ'>�Ƃo3�m�v�����c>��8��<ig��O����\+ʑ�Y9� �^6wj?u��V*|�ur�9��2J�p�\�5y~��O���5=�瑡��r�rǇ/���Tr�Ou�Fג]�۷AW�O��ٺ�Lڠ��Z\o�C�V��-�̬���,����웍p��$�;���	v��!h���LS6+�UY��1�+fO"���{u_e:F/&��i7՞՛hY�$>k�itk�T3�A49h�XJv��
0���j�xK��Yf��6�K��wuӂ	��"����Dv2�i�k��'[SN���A��J�Ӥ�x���3���)�X	iw�o�����׼z����烑����T�p��:�b���M�gĵpe��x�$��!����=�/���資��zVH1����z�++ԇ�7���+���a���U1u2�ꩉX�� t߲,���r�&��������;���\C���&��.J5�,���8|��A{a�IN��m�{+n��h罗q>7�?u���ߴ�y���� ��yQ�X}�6J� )ͬq.����򹕵��}\i�>Q��j9�{�=s�ZG>>��\_�þ�T�fQ�E[�]��}U;��T�F�����A��U1>u����0s�.����1�}�m��΁�}9���e��߻{����7�fB$���2$�2)�za�ꑛ�5l0v��*H@I�ޜ�K�)
/�M�/�=Q�*:�@�=�f���ϥ�z��K]6���r��]�rC��y�B�2\��UG����<g�o�;���A�RɌ=����/G�Rp~XU��~����n���y�~��W%I!��̳fX���	W���w��U"&�e���V�J��S~��{n�X�k�����&НWՈB�F���*��3��Xa�6�.c{h�.8���X��3cZW4y�C��\r
y���ơ�$_�Mߣ޸|o���2=�WF�������q}��h�gޖV���x�)����y�=��U��~��KM��qh�%/����,O�h�k��7ۨ����,\q{3���ݼ>�Ǽ��G�j\�������ۊ�?�U>�@�L�દ�*��f��3��K����+q�+�c�`��[���7g��z|+�A���3�ꁳ���:��NgK��G�C�~���%fǽ�]��:d�f���X�ϼ�����Ӱ�'v��<��X�3�K�=�M09E�?4�&�T������k� d���i�>�׼{)��!��Y3Ǿ�ωJ��<5z��z��f�K��S���w�}9~ףƨC�>vE��Ss��������r�.���r�<jJ�-yÿ3S6mno�{4��\}�;⨨��kwp�z}�o�x���\{�g�|5D�pW�6J�*K�2��6��+�����Oz&|��Tt��>��Y���u�>�)>/�o�3מW��/DEh�~��������F��,	�
W���l�����"��Bn}�CFC{�h׼����S�W�z����-��Z)1@����<�e೩�p��k����%LJl������+^���YmN��+}ԕK�=�lL�?l��]�\�	��{����4�e�X�I8]������f�2��*�N:�B��Y�Չם�������)�(鰠�ח�q;�|.K5
	Q�x��E���;�΅q�ւ�T�n+�SN��_F瘲&o�<}����ޮ�n3޸:}>���d���މ�bbW���t�}Ͻۇ1�����X�f�P63�5��4[~v�z�>��ɿ��\��q4�}2��x�e[��矞����!t����h��%p�o��G[j�F��H`�x��6��&iK'��[>�����x.��t�!�'���N�:*n[;gx�/����{����d�{ޠ;�����3��w"�狺�>�f���%�l{jV�����oS�q����0��+�&�/��9���^ʞ�&_�^������a�7|J�0������t\Ru��t���w��� ����7p�8�9�=��'/|�ī�^���q���qaz�7>�%��?G�E���y�s�#�/� �?>�3�^�fwޥ�������AF�T��,��a���P�ٝ� ����{iz8���>��^��O����M�ȧQ��u�y� �NI�>%������y�'jf��;��3n��f^A>Ά��=�ɋ��1-�O"�˔z�QeU�WV`B8�sѭu�7]�f0�ʵ��L�Ξi�f7M�.a��E�ƒpfؑ����� 4+]� ����l�R�9�t���+n\u�Yr�L38s�~nP7W����v��qRzŪ*��l-�(��V�g�j!Dr��P��Zy���_�^8rTy{$9�aG� }K�N��J�Y�f�Mt�ݍ՛�cY'b����ۜ��٘�N�K5ۓgdt�,΁;�wL�u��mj��"���>���;��E�su����j�stS��0�mt���p!LN�d�Y5�ZADgh�za8�+�������ܒm[N��ս�v)���7v�yZp�y���_�)��8��{��v̮�8��E�E����*�ʵ�~���wM�4Έ7q�.�5}�=뗼R���]*�7ͺVa�!\T�r՗�E&�O�۲�
��t��HB���IH��6����D�yh�]Qӵ˄ѯ^Dm�Ҝ`cWƎb�j��E*��I�Yͦ�Ҙ��i8;ENY�w8��k��Ƿg#�����2�PQą��U����Y�gup�[�����v�}�K��81l�DS����	:mס��S��W������,Soq`�3���-�k������)�03�]�O�ij��ŉ���fh��,�׶LT��񽣤��^g�i>��)E2ybʺMD��qu��]���+����9�Kk��ۏ:JL)e�%�{�\ӐAԓ�q5�c}�cO���Jݖ5����Z���ŀ��#Z��(8f+�W�y+oNw_�h�j�o�����&��� �V����w.:B�ՙ��,�%�ur���(��e-�Wn��Z,X�u��S�
qOȞV^ia��be��6&�c�T�wxn�ǎ�}�
�F����ƈz�!�+�z`�ޚ�����_�5���_
r��HA��V� �Ļ��b�P���ɍ;�1�����B9����{Zj%�_�ø�"�Y�R���Y�.L:
X-��2�b1��J�7Z�Ω�ͽ��R���qu)��`��5q�|�RH&��٪ҵO�w'7fmrA �:��)yL��_h�YV�̩Xx���S�5�ܴK���iRɍ��]{B6{Q���ح|�GN#.Y�5��ݭ����,���r�b"�)δ�V�����ԏ���x��;�4`�l��d{C^b��R���ʛ�2s'�eB��Y�nDH��y]�bw2�6?Y�#� T�@\��=�2�Vf���n����K��N�T��R�v�o��`^�����8J[W�u&n��L.WZ��=��᩹�9�V]�a�����㽖kfE�Z@��X���L��L�1�C��O��M�Lͺ���w�Rb�He�}`օ�I8l=��!�j��&����^�2����7�5��f	eB " E`�@���Dےk���n�w"�r�ʹi�n#8���t��W7.bۻ��Q"7s����\5�H�(�6���p��5�ۚ�˛��5���s��]�n��]ݸksFM�r�I��]�;�Q���vc��Μ��sd��ݺbJSr�˖����lk��sQb��s�nk�$��'"+���9s�.�1"�ۤY��9���X����9wX��Q�rѹs1Q���ͮ��])��r��ʹs�5���9�wRɋ���㺹lc�3�]ڋ\��.��r�˕wv؃9u]��\���]F�g ��<�C�j��]8���M���!�F�k07�v���@b�%������ol"�Pp��q��NE3�����Ƶ�~����GL�����6��uz��<��+��m�� ��j���s�UG=Rtz-I'��x&xz�g�b��t%���X|=>}�����x���S�(���=z��"w���g��#Q��g�����~�|�R�x�,ʖn��q����B���<ݽ^��\}��g�brx��w�k�p��n��[0��+u#0����uLN�Uю�=�YR�ޒr|ďD��џ?my��ޡ�\g���:�b�H�Tf	-��{W�eP,�m5�ς[�}\mxz�Y��~WO����#��\8��z��L�;�K��@˧�*%��s5n�O�v�Ǖl��M��ll�^�1���1���m�>�����h6���/�~2oX������;[Z��e�{��N�qI�B��4xv�/����m�+�~�"|s�9�}��-�_����~�eD� =@z:i*G���ǝ����X�q��T����������yE��u��ux#$���l�p�2=>�$�Ȳz0���1R�މ�>�y����[P��½e~�%B�n���0�U��t��v�K��W��E����K��)��n���e.�3w���'6l����S�ٹ����4��i�hU*𡖵ub/S�3�[��a�Қ�Ɉ�pAW̆�Fb��h�u��P�<s�:�5�/waB���`��~wt.3ޠ�n=����4X��eH5�O�U2a���պo�hGFP��u\���g�$I�n��7~;k+áz����P����ɡ��[_nx5a�~2�r�J��*l���쮛��R��/	���>�m߆C��p��5=���F�U��-rǁ��GJ�5nϯN}eK�+�%t���'�6�%�ȣy2�Wؼ�=��������+=�q�%�&o�Lπ���8q��z��<s&P��GN�_�0�m~g@^C�)�x���	���1�J{��D��z�{��O����qݎ�����A���X��S>F��^}��aϣ�.�����y��2}��p��{������!�񍏗eJ7e�z���KJF�Y�!����͊��Ѵ�D�����<��޽���;����1�Z��ڃMj�\�҇��L���:i׵�t�F��;��+^]���{�q7>w�9�'�{#}@>7�TF�:��d�O�L�>�>�0 ��}�-����>����ucQ�~Wq�ZDxߊҟ�i�o�F7恸P��ڞ�;fE�nPS�����22��ïx,�\��:E���c�6�uqIv�]2�N���j<������K��ٕ�2�
�������gl�vu,�9E�wI:��4�ԧ�<�7��N�j�fwR".��>%�05K7�8�nP<�Eж�G�����|��>��DL�\��~,n�3��kT�ϥ��1���ټ�F�Z�|��kv�Vr�ȟOӨ;��Lȯ��eI�㤎�+�h\Rt�y����T��c���L^t��f�o�a'Eϰp��zώzg/>��:u�r{`L�������Fp��~�������D�6e߳q�'�{���B�y]�Mω����Q�?UH<Y:���eB���s'�[���UR��jϢ�>��ިzW?m�d{ή��?Po�z�Cɡ޹�x���f�4�+�Gj^{ܕҞ:|ģ����Z� ~՟���L��5'�n��m����;X�~��l�z�V~�8���̼�t	G�����Q��u�Pգ��exl�|N����}��=�C��q��?E/��&�N�6�<�-�jkeDנ׾���n<o�p�㓛3��4�{�NQ�f�~'sU0+s�#�zv੅]�p�9�P����*w�y��og��1{�S��d��O�b�&��t��09�4^#��s��dפ}�z�2=O��}R��E:C���T���`��	�+�7�kܴM�nS/>�t�����Ρ����)?����(V~t����-�����x;�	�R��T�/.�xt؟l�%�5ʵ8z^�\�c�S4���Y��s�J��T�u�}lܕz�x${H�ٝL�J�E5*���f�mk���=[��Qݵߖ�^���T!`n���)����{�z��F�ۙ�\�O�}��7�[��U'�����2�:����Y����y���;�<^=�Ǽ�>����r�.��y�n�Ky@���7��J�L�$%Q�%���]K7�7V&㛿qϣ�O����m�'��|�v�=ޗ��W�ߠ����`��B�UX��-���zP�>������:�~��򅼽
䓞�)���������f��,҂Td-��g�y���΄��>�쯬zgse���NKb�{��w���;��u��ꉨfK5�"px��^��.&k4쥙�r���ϻ��|=Q���$h����(�x�C����_�&���e\!�m�ӯ�7*�Y]��4�js�{�^�F�S=y���7�y����W�7ޤ�z� �C�~uNL�TNr����?j�vs(�I��̦G��T���l�/K�~�d{��2�L�y��P��o��r0t��l"�O�8eL�a�e�l)=���}~�/N����o�h�߻3s�:��D\�xv�ՋbN��,�xvW[�}S��
�ֶ�Kg�M��x3�`�-���Tr\�zV������]�W]��3�=��pŧ�x�\�20àU'��roT춠��GB�[�0��2�"U��#�����g��(3*=���eٯ)>�ޞ�=~���6xx�C&�Z�i��I���ǹ
��}���;���)��0{�~��3���/K�*�*�}z,�^��B�%vP߬v�??�X��/�̻���u�K�w���ny߆C���3��R�y�V7����̩�'3L�õn7�NU�/-���z7�J���l��i�*17dZ�M��u�[s���̳��MO�d��ަ�*�'`����~���_ڏ_�R�F����<O�5}^&�9~>��ǼVEy\ox����UO���	ܗx��OO@���C�}$���|��L�L_�n������8��������b�L�ѡ������I��o���|��G��7~���|�R�x�̩f[�L�B��x�`�����Ƒ3�'
P�}��?:�j3~0�G!P,	�n���}������pqz�+��q��ў{^eoz��q���t����" yW�a�Y]�b;1h�ߛ�j�U��'������F�k򸛈�yb��W������g�Dm��%�\�T;����*c�v�gaY�\$S	�U��Xy7��M�b�J��V����J��"����_���r�w]x����R����VM77鵵,>]��wf���Ɔ!'RF�q��ST�7˄�cywh���"ߣ5�$�}i��M�����wl������,҇�h�9�^��'��2}�I-Wc���v��n5�Q�	��8}9��;��߽|�h�_	�q���n��OTz�Ͼ�u�5)��A��
ȥM�/���#Q���F��|��~ŸOG��5<����ȗ\K�u�3(���= �^�X*%�xМr��}�����q����\w�}{�(�.}�c��;2m�}��F�Q�qOPɇ��a�����N������۪7k"��}��qW�=�=���2<�wB��9��z|���4X��T�Q��U�}bwL(�<����ENc��_�Pu����+����R�8_m��d/Uy�ޡ�K#�}x��ߖ�0�����x�;xଃ�������<g�O�a���72��9��~7����ϴ��槝L�{��5E���e{Ѽ���+�RW�O�ng�k�C����pJ�(��2�V/;�92�|K�+�̩��Z��O�b����+�5�Y��\�i�KE��t����?�%[_��t<�#fX
�K�x�/=���솹v|t}���qݟ:�b�;*tݖO���2����ϑ��A�����[֪��ˆ�"t��`��޺:�J���!��̳�e[��v���Ɲ������qL	n����;.N�cGP��{7���(��y��/��x��4<6��R�-�i ^t�w��]��%����f䤫dWbuw����xжܺ��5�Vf�a��e&���4}����`��G������*}({����e��=_��FU1v�|!ג�����ʬ��a�Dz�}qO�bx�ף#}�w#}@>��c�r&炱rQ�E�V����UD�\�4�\���l �cg�/���'����>u�=�'�{#}@>9�$g:�q�J��	W�N�kg�2ω7� �}Pμ���ϵՍG"����O�i>��\_�é�N*y�Ƕ�[�
� �Ez֙�2
4��UD��-�������3��R�)~��^���S/��6�U�&���=3�M�޸=q��K*L7����+�h\Rt�{a�������]��0��H�{�hxyQ�G�q��z�`S�Q4��=qf��=������f�م��n����W�no��!��;��{���n�O�����@~��s�,��C��:���ev��rܪ��z[��t�;y��㟶�2=�WF����ǽ~��ڱ}��=�}r����7��훪��(&F�V鿫g�|����7��>O�h���@zM�n�tJh287{���v
������p�S�f�6.�n�Vh^W(�NL�y�!�	N�ѦL���>�bG,�YU}8�.�_��{^�~�׎ښ����tO�K��nq�#��ϡ�����U�p�k�R�7���S�v���V�j0��gr�;��-�$�u�F��?���3���|r|��r|3~�T��=����wϝM{�N:J�F�s)�>�S$T{4矮૏߯xߍ�8n��ۙ��CgC�����*�N���"禯�ޅ \�=����V{�c{ʵ˹�)N�0�>�>E���kN�G���M����GW��`����x��x�P���z��=.P�/�<jڞ7|JVf8�ڄ�˪K�Μ����R�񿩺�#�P�x[�/�����q^�<NW
�vT�{�W������]T7��ຟ"O1�|g�
A�;s���wp��s}#��o�=�9^u��T�Q��-��~P���X~�l��J���50�[��eԳt�X����s�O��;�*��o*&����EL������\>�p(R��A��R�f�Ke�}u�9^�!&�=s|Ɍz�wtgz,��XA�t��;�4��z�����w���B�Td-��pzW��Ɂ��F]��ѧ�W����D�;c"������&�=냧��`�T" 7Qx�Ϣ/W���N�V�r=GB�����]�`�Zw����`�����!�z�s�^z�`u��>��n񊑐�!rJ|J$�ҝ����P�J��`��Tl�q|A�?��� sلg���t��G�� �E�.A�Ӽm\��.�������Jf������}��g���F��k$h��?;c�H�dx�M����/��d�eV�R��Y����������D��Te����q�3Q���~� }�=^ o��� �zG�Ńv�o�tZ�ܓ(L��l��
�3��S���7+�l��R��s�\y���x�9�3%�Z�w��4v&�&=T+�}s&��zh��Ӂ��+N�����{����yp����׺;��W�]�m(�>�1�7��K�;�׶o����>%PɆ�և'�pm'\O8�u�#k���{]���Ѿ~�І}�^Y��P^��yU�[��A������홅��a�)u<�NF�b�ͮ�z����J�uS /�q��ϝW�����x��걼r�G���ܾ53�%Z�x/�wy,�ܣQU�
�N�z�o�ʭ72�J��^ TF&�U)�9�:�]8ۮ>��C�DU.T�n/�e~ٲ�E��������n����*\��'c��v\�gsX�u��[�T���	�^�����gNI�qjI=S(z	��|�/��t%οMuT��A�:�X���ش�i�Qt���*p����a���%_a���f����k�F��tgy+X�}ke<U���mW�IcF�j��R��'(x�b2#���/D�6ev�K��3�V:]�-�번�U���E:�������N����@TU�;Ws�ݝ�R�A�Ә}��Y�q��3�k�{�q��X<�T�2����3hz�m���e�}��c�Gz=LnG��=p��=���b�P��*�2��R$s�gQ��u{�܆���]r�L���"�|�z3�k̭��*�ԁ�n�C�rY�D%�"�jÚ|k'7;}�\��q�9�|v|��b��o�~W}�h\�����q7�Q~�bq�١�2>�뷊W�N\���B r"�'θ-n��F�q����m����>��Nւ��y;����o(r:����6�ә%�$�g`��2�HU�J�<;`)~7�F�o��~�]^ꝥ��L�
�����q>Ͼ��d���3��`��4V:\o#�>&c���IH��>�����C���H�?+�1??Y�p�>�އ1��t�̓P�'� d���1R�ޅ�oE��K��ۧ�R/ٶ��UaC~��c�3~���y���{*A���*�d��fd���+��hU�����۪���OMҕ��a+���Y^�U�rz��,��x'���V-^T�ߢ���.�B�v�tu�A�(^Zt�if����2pR���]Έ�k�C�o*���kD̀K5��?�Ѩ�%*uF�έ�u��j��*IތUۄ��Q�sy����V��:P�"4n�������R�/�K�QD�K�{,����W)њ������k86r� ����c��;c�F��%G���FvR���[� J*C���
4&�� a��,ɯT�Y�a�b�|z��d�J��̽�`�ҋ��TC�Q�L|����2��W���-�M9�Y�M$s����
�W�m��aw��^��2g7������X�wgU�mG�D5}�.p96V���i�6w7�^uB+��r5�Ź�o6jM5%��**������J�g%LT��vRX;92��e՘��)�ڗ�����&�r�t�������]��p++2i3pwMB*��`�&�1�խ��f���Ƞ�ntČ�2Rik!;�;�ٓL��|V^�v�p��a]X;/)p
#�O_E�Zȝ���3qu���d��ͫrÆ��:���DZ�ʂ�7� F�)T͒b��["dW>b��G��v�3L��cx����BIݚ��I�u�_U�x����%�&>��[�V�VPC�ﭧ\�8��nsO�h9M��G�*� ���Wd�:���}�wp�5����	��'w)wuv�l_i�A���9��#��R�n���(0Wv@R�uƔǠ	�_nQj'u�C��Nnn�}ՍS셎_]�w%8�W�L� jʶ�B�x��\=6u=dL�*p,����ҦU�ה�TW�Ájw)�'�V%�Q]ܡ�{�fP��Y���L,g�XX�����}o��e�X�ts���bw]���<�B����4uc��nyy�s�!�1�����O�V.�'�X�>���Ա���:Z���im���� ji�1t��������,�p9R�bYP�
�7��'�3)�6t)V��q���>��E
�n��JCc,n+���bx5P����n���*F��S)jǕ��[ډ��M�n�T�0����B5���sH��k���A���:0�W�<���2�a��G3_$
u=
�W�E'	���#V��9TL;��m��:��^�8+��]�w���v�NK�^���୮{wL^���%�.Qd���].p�݅8������s�r���[/�u��pF��}jg۳[#UZ��re�ų�M�V�h�
�[�5�����hz��ŉև��ƫ�A��-`�Րs��K�y1.J��9�ii2,Y�&<+��wK\�JQ��lٍYb��}��H�k{iH���kW1\q��^�d՘��2��Rw�uYY]@��B�16��N^�wf,|����tI-��VԝR��h��i�c�jd=\u����*v�9�.�� #��cm4��7|�� `d�ÑS�rW6�}�Nb���uZ�+�gqd78Z�ەC��2H**J+S�p!�-v[B��&�I�
��k�.fb�Z���59u�ńNr+�0]�A�F.q(�v�&
���;�T�s��sbэ�`�&F";���st�ƍ]݌E��ɂ4$���t���1�j� ��F,�F�]�v�r�%)�\ţQ�G9��ʌ�#9Ҙ�Fb��FK���X$����E�$���B
*�����B���d��m�Rde	\۲�E)�`f(Ѡ��2��PQ�sbD�	 ��1�W^�55�ߜ��%�샻��S#Z���'�r�nP����6����$Vyp{�"JwVn���
�_-[�����u�N0�>�W�lg��ݨ묯#qS>�t�~7����ϴ���>�u��'�)<|��⣺���޹�9������s��eW%x�z#f\
�^WȇSO���mt��9uZ���<d�f��?;�X�|�ƛɝ�'N�L��O�>���:S�2�U��7�'���Éð2}����,�]{ǳ覮;�j1Y�S��|��� �/��7�����ډ�y�t}Z��~S4����"�ǩ�������!��3�b�eJ7e�z�3��}����񴽷���´���g|n)]A��%�!1�V���;�o���Ǵ����rQ���ث����|I��@�ިW]4�{��'���;��2|�s����*#}��W0"���=��}�:ވ����'��x���z�"��\I��"��<W�a��K�7��@0�su#=��s �P��UO���n�/ō`�8�xu���v�T�y�3�Y.�Ǿ>�Z��L�p�����Nd�Q
��D���E'Kǭ|�z�Z�fG�\{n���s&^Q�9f�4&3����B1ަ��[�JV���BzX~��_�W��,oZ���^��uwp|ju����)��7��ol�j���fskVp�":m��Ы-j*A����oUځ;�cW!+�*��+�r�ԧ��Pw��C�{�����=3���@�F���:���2�	W~��Հ1�-k�ߧ�b�VV�Q�Ez[鼄��w�H�^�p�����u�]�(�y�hK�~yUSGSXٵ4�D��l�V�g�7��~�����]��Ͻ^O�ؘ�u�D�1��;�o=V--y��a��m�u�U��!�y��6<��(���v�Dk��/ٮ���W�}}�Jh��M{��b�����O�Daal@���'�6�>'�wK�m�x�v�Vz�n׽x��v��(�>�0҉�W��]�W�����g
99�>�᳡��:��Nu���@�f+�y��j�;��@z�d1��~�>�g���U��+�b�72�J�̓0��b��J��b���>������&}��o4׀��;^2?W�q���dS�;�C�R�jx��)a��t���jf�}�lS|�0>���~���5F3���8�W���)��W��W��NW��1^wbD7�n��	�9>����I�̂�=�F|���.�z��<�>�i��H�{�o�=�5������P��і�9�	(ٳB<�eg�M὎$�#�1�f���c;|�����#_T��$ڀX�w�a 4Z�'h�IZ����#�.��!�z!��St���u�^n̩KyL�nW�N�Z�s�3M���Mk}�ڧ�8�)����C� �>E�OlL�$yT;��[���R��7V&㛿q̳�P���u���{вI�Ӝ}�%��|2��A��J�-�2]o�<�yY�SN��Wz��z	���|���h�zF�y�\�U3��f�P@J��~�o��/W�<�8�:d��q�U��u��x΅k�����0={Ho�����z���z�X%��D��+7�U�*��Lr[g�Lz&�*7��}�Q��Z���ޤO��O?z���뉞�SW6��G{svy�̲���F3g���]E��������m���m�ԁ�@�x��躘����M_�4�r��"�yq0:){��,���5�����/�����;�:�K������wrH/t�>����G�GT���<5�NqR��}^�z�<<K�/U:>���;&�����z+�n#�.���������O��nl�_Z��Hǋ���ס���'���u��ڬ�呑����yU�W��b��N�,�ۃ�ߵ���E�c�o?�B�~���٢�#�Rj�潸�BB��5�J���:���N��o0���0Zn�K$����;l�<ĸ)S������x%�n�3h�&ХHb[Jiz�����n4��+����,y]�f���#QSӤs�6�v�>�~�tѺ�V���������z�����S^���e��T��e�5*��.;�A��%�cl�uG�+*��EL�ĭ���-T���:�]9����ת�;E��~���p�z����$��D��3�5�W^�G��etϠ=�М�p��r��{�6Q���g*�)6�f_�l�o�i>����j�� =�2A<��1�n����~�.�]5	!>��JKd�A���Zr#ޟx��u��?b�Y��P�h��	�,��q���x���UY��^g�{��R�����V&���p��G��Ͻ�Y�~w�k�Q(���%T`xI��7�}��ҥ�� #ݳ���}��#�|�z2#�k̭�PҮ3ԁ�p��;�rY4�gRy�׃|7'���z�Z�M�zS/w��5�~W}�h\�����y�Q�9 r�.�3z6���j�Ov|���q�p6:Z>݆j5�h�r~�˃��>�۬����v<�����9>�}���/�M�,�Z;��8��/ԅ\E*h��
_���F�j2/����	��;��}���Dޅy)C��f�ā�3�K�ܱ�
Yk��)Ӡh,2�{�&p�w4�\Tn6F��<��ơ��WZv�NE�Ԯ�< �Xq�g3c���P̈́h�L�i�v�SR�.�e��9Pȧ�st�N����[/=���m�Τ-g�G��=�|s�9�}�h�d��Y鯌�/X��Y���o�Zm�H1��h�՞��=�|��C�����߬ɷ���@u>�$�,��0�`O����=;����ǻw�R���v%�zo6P�UV�7���ϼ|�;�A�{*A��T�Ǳ�8���-�*�I�^�^�1�S�ei�wW��v�߂�ϸ�ޡ�K=ׂx�{�VS0�}&�3��{��WK��
t���ȌɏtVW���e�:u��;m߆C��q>s�m���ũ�>�-��;r�נ�̽�s�r������2}:�eW�J�(�F̸������o��`����K��hT�q�}���X��9b��7��-ߑӷIxc��Pr?�Ѵ_��J�6�C��SJ�����2k�����K��.=u�Ȋj�>u��u��؋,�+2�P3Ņ�Ӽȵ�uv�z֕�]���^��y��a����z�������z�F1�G�9�|��/\����|�E���WA���Z�� F#C��j���Fo�|�������&�q�]��������T/T!�,����㚍�Twz���jaf�X���v��1@�veZ��U�8�(t?^�e^*�i\�\��+�k���q]��1�[�[F:|���#�v�3��J�Bm�A>�Gaa,��T�^���A�"�x1�<���h����%T�`�Q뮚l����O�׽�s�~Ӟr|�}@>=5�_��=Dz��z}
�̦E{�\=p�� ������u�nKe�k��}��&�޴��;�S���=���ۅr����=~�\���4�ә�PB*��Anx/ō�gQ�j��Wv��<{�yϖr|ŗ���w���zgt�~����W��s%��U0ݎ�&$�)��P��e�s:�|�.Y�{�e{�Pw�W#��x0���ώzg/ z�`T:uH˓�f��̓K���^y;i��%�S���tg
{7Еxz�;��x\{����>���Q�l?]�7�^9{F��Om��;ɺ�I;�Bf�eE}��L����޸|y�+��ST}�?Pn=��}���yqˮ�b�B/���,��|�Ī�gg��V鸊�||��/��m��O�\}E�nV���-��H�6O�먝~ˡ�}�9t�QXZ6t;�++�n�>'�Gt����d��]q1s�Gvzr��T������;�pW�՜{�fp�����>�l�w9GFͬQ��m����v��H|5��Y^����1�T��e9M�Sa�7NI��+�J�X�\��	K5�7�7w�]o�M�>�܏6we�O8�ӧ��i�����(�
����"��OPj��:���Nk��kN��$u��P91X<��D������_��ަ�ǂ��?g���s+ޚ���0�s*t����3"l����'�ם������}Ji�TZ%����߯�箽���:C����H^���c�/"��H>�����NF��f[%���a���C�UH�Es��2!Xn�x�7=^�t��1�T9jb�2��]���#��T�v�%�a��HOdu	O�Y+�|�_uP�a�{N���i�5P�f��lʟkH7����ً�?��LX��l�|�Lt��Cʡ�L�>�˩f�)��'�b'��]�����S�G�r|_�t�{<��3l��E@�~�,	��x��:[,O3鲻9�"�e��c]"2{�g�W�!7�hho=O��Hҳި9ުfQ,�( %_b�dghpVw�{��=u~|����9�gB���A�:a����k��%C�}AZ��ø��,O	W�B��o��}>3 �c��u��#�1�}�d�	��}�D�"<g&߽\^l���j����H	U}�s.�Č��W��-��p�{��g6��m�ԁ�d~��u]���jN��Ӫ�F�ݚ՝�Ț�Z�Σ�.]o�fwKʝa�ֵED���o���W�2@�77Q��[��\�\扴�������:�����2!���t��g�*e��z���u%�u\�+��^���_V�B;3��)Hm����wbߠ:�ʓ9�O
�2�l��Q/�E\VR��9�_�~�)MT"�/IS4�N2Eϲ���zy�&߽@w�̍��/��'���]���ӡo��._!<�ۗz���9Y�s�*��
uu����1���>��N�?^ٸ��3�㏉Q��ZU߻ܽ9��Q�9�-RqJs��:d�t���w��"��##_�/K���Ղ����ѥ���T<3�;o0�ϴ�˙��P�*~�{[rj����
��;��U��g}�^/!z�o�u!�˯,��c�p�y������;�f=��UrgN���+"4� TbnȸU)�9�5t���Z^��A��q��;��{H~�S�z��P͈�xh�T+��H�\�g:g���x����Qc~��yp�)Y ��w��*|�3z=��}�9'E2I��.��=�SK�*�����.��i��ۖ����<h�G{������<^������:�j�9ơ�(�$�2���X���͐��c�OeU����eO��O�bo�~���1��,����3~0�\�P�%?u$���pb��ѵ;(��0��r��Ez��]�ʏ�J^+Rm�//I>$Q�mi�Z�r���L�:�]��[��jP��:�FC���QǏŦu�6��Bd\��&�j�-oOI=%�D�Y�/2v�VЈsp���g�-�RFs"����X������A����GO��F}��V��iW�@�N���d��ҳT�@̲<x�:���pzW�݀�5��q7>��0�+���W'3�n�д�n�������W ���:�Nd���r<H�n������1��h�r~��s�$c�p$d�R�r�R��g�g'�{޾�7�,�Z:j[#��HUҦ��_���NgIQ��:V%(�%�{�{�ѿz|�����x�g�ր̲FB,��A���X*\��
��j%�.��׫.Ww����6���s�H����_ͿY�p�>��σ����2N"�ꁓ�V��9����,���c]V�W��z[w�"���ަ;�U��UNB�l���4X��T��^^�t���*b��=�����W����~��atR��t��|��Å�v�߂�ϸ��k�Չ�Txa�v\�2�y�8��N��0��E�ω��dn�>��#u2��9���vۿ�U^�N�䥱3����"j��`�����������9�=X��WK����x	��*
^���[|EP���&=�S�ُ��}���<�����!\�b��n�F�)u��b�L��[�Y���iF􄤾�hb���Ư�o� ��=�* lme����.��s���W5+c��9��V�7T�	�_U�3�.��÷C��t��y�I�c���ъ��֓�&�U�֯�]��P����z��L����VG��9/V���y3�פ�ۙc(L�R}'A��X@�7�z;z�	ʶ-O�2�w���o����T��U5qݐ�|�jɞ=|J@�{�}7���{���ݝQMa�$�>v�x������>�1ǥ�_C�{�dW�u��*�� _��z�C3(f����l�{�f7ƌ������7�PU�%�!g��z27�>gr#}@>��c�}�隁�潹��R��tO� z'O��D�Q�p�Þ2�Q
������u��O��O�>s��������������50<����#nS��U) yMD�7> t�^Dk���*��߹
��~���7f}�|}8�q�zF�����m�i��25
ETO���n�/ō�4gEu߲.�˰��7���^t�ȗ�l�g[g}3�K���g�B$��L7c��4��������8z�ѩ�����4=�I��f|=o���^W��|}�g�=3���=Q�*>t�&��:����c:��=��>=ۄ�2�0w'h���k��*�_kW!����������;χ����~��V����V�����j���km�km��j���-�խ��m�խ��V�j���-�խ����j����m�km���ڵ����ڵ��m��m��mZ�~V�j�����j���-�խ��-�խ��m�խ��[m�[o�m�խ���mZ��b��L��fb��̓� � ���fO� ď��{|��l
h�-�i� lA��UUhV��PV���h)� ֨�"� ����6[@ �4=�]�k((AIH��>�EJ�P�j���UH�fRUJ��mu��Rv�ED(I֤Z`Q
�4*��U"EH U�����UJH$TR���U$�H�إ�(E
�%))$( "�V����Um�I�RUJ*(�9�);iR�D���P(J_  �o;�]��:i �wP���P�1�R��:άu��k���S�l�Y�l��gF���U�vAJ���֎�%t4R�[b�� ��  ,xz��k\�ۻ��
�2��@v��=EP�뎊 QEQ�}=•�(��3/p�E (���s�(��(��K�[�(��(��Gp��(��(�uHO�	R��e�(�f�;g�  D=Qh��ajڨ֭ۻ��5;	��j�W�� ҹrJ�`j��Z���p�EJ�uҊl��B����4�   l��k�ͨ�S
����iѸ2��v�"P�Mu�m�J�۶��k4v*�-�h�m�r����خ2�څ)P^�"M� I �  g��[�(�ۚZ�����T��=�8�M(m�n�u�m�Ŋkj4 ��]�v�Tn˪cCN�]��gtn�h0b�S]w`,D��@v7��'�J�o�  �A�뫫v���j����Mt�����mu�5m[TXt 髗��vκj��7.΋�͠�av�9l(P6kUj��h�5�b���wn�MeJT��   6�yݴu�vwE�t��۱�V��uj�C
 �M�7݀��q�mֻ�����Ӻ�M�u �5C��2�,��v5��
�UT����@�J��<   �� {��9��4R�jӭ�7cLҰm����nР��� ��I�8��M;r��Mڴ�[f���ӷv����+]9Ԣ��lER�n���D�x  Ļ���كWek�XKee����8��v��۵���4黇5F�t�N�9��-v���e�:�[q֨���ZН�B�Z�*�l�!J$���  ؼ��(iۣ�
P�[�������L�ûi͎�g]��\i�V�:�:mv�SA�݃��lnC;�� ��]wn�s�So D�*QP�L��O�* �UO���1R����&�#O��T� 5M��"��M 0�RSUDP�x�N��׵��n�����n۩��w��9OVO��[/�3"�~ ��|�}�� >��������D��* ��AQdE7�{�����;������5�k �W�4H�&�_Ə+�8%�Ьc#k<J���a|�y��T�%�7���Şr������h&�X.`�����z�*�K����e5!L>O
w�|�������ᝬ�6�V�+��Ɔ������Ԭ�e�d���Hϖ t���9�l�s0n�F��lH���uuc�^�kjۗI�\)�4+<F����!eԮ��Zo3HyWw�DCV������j�r�_�2ŬjԀ��VKف��j�,T�ퟕ̰� h��y�x���v�id�]���u�)j7�`V���+\��mi�x��Z��{�u+��N���]���x��H��u�V�����U�a|��
�A��*�b1�ȓ���h�Z���/KE��x~v/wbX(ໆ�9Zh�#y#zh՝�M��X5�M��Sqk[�!�[i�b�2 7�����t�l��e���Pa�WƮi��$3�-b���Ɇ�e$P�0�2`vsA��[)�|��]cn��K5�R8�]�n�s#����pU`���y����Tjn�d?dy�j�V�s.��8-��Ì���j���[�"[Y,h�f�c���B�)�H���6��'XZv��T@H:ڒZ�`��<·N��P
�Ʌ.%.�kb����;@��L��m�n�I�2���%ٳQQ����؞M�XǏ�%�U~��1�Ef�1y7H��S_�{q�;�+�U�Z��i[P�YP�d�I����3��ҬV����I��ѷ���t�^dU*-�^��b�Q����үw4�-�Z�l^�tU�pӍb�9*�z�Z6'�髳�E�{R���sҪ9Fcj����L߮�_;.X���R�A/FXv���;J�H�t(�Ր:�ZXչe꼨7�Y�GI8�>zpi"fe�2�m:F*
�n�(	W&�LVÉ��0V�(��p̎72�Bh���u+C�k&m�xCs@f�t��p'ff/0`�x��Z��ueH5V�H[E�d�Z7*�WE�mɳ�7H�qn�.�y�j��,�}���]�h�������}XX6��{��h�7Y��	�1���n�F��؎�E8#֕��I��k*�;eȚ�S�^h���͛a��/[Di+1�l֜�B�7h��sr�;t@!���/M��j����ҕ��<���e����I�Z�NM-<P�P:����ڻ�Z����k	=*�����uY��(���mkՏ�wxn��v�H��%j<�-������RU�X�+p����)L#�lEi3G�vE�)R�J��(��W�ޗ��2:(@����f�^,F�����T3!.�ֆ��\�z㤉q6�\t����!b�(���qm�E��v���W��F����"*�C�خA�֗oV�N��i��p��`�GZ�"V�њj�B�\�Z��i�=��-S��P3G2�;�I�0a8s)\ ի0�2�,�Z
��x�5ЈF���.�ͪ��.����%ʷ��w�6Zx�o+b�� Ҍ��:ۼ���������ېT:1 ߌ�X�Q餪C.�B�V�4�Z0ճ���v��TK�ddہ}�k	^�o^j+4��Q�n;ú�4jHVxDZW|��A���;�C��X�D�4�n9+[�;�V�b�:EBn��Vh�M��z���Kvi8÷�cq����j�0�Y �ةϦ-��.��f�n������*a�U4�VU���![�Ɔ<�	���`�K$D��+'.���{U ͝ 
�Q�)ٹ�ܛwx��Ԕ�t����PLl5ik�iޱ���yn�d�n�2��J�n����ԉ0+�BU��W���65�*]�f�e]X��`��hӘ/r��F2�F�ڼHY�����UԼƒ�wl���`c^Ѱ��^�H�S�6��gY�peP��d�J�j��L	u����1�F��.\)(Mݼ��sjmF :-����v�J�̶�,�tn�Y���HFI7wn*9K2@��a`:j:XK[��D1��{)�V�����d�ar�Y���N��������:R������{J�����[�*�����f%{h�T�- ��v�0�
�+�r���eӬ�۰u�IaN�m�aR��e�3-���8eb�]��`���G��Qπf�p��%�:�YW!��Q�h
�2���1�Z�L��0K��"�r�u�dWHnZ����.�S�X�������Ci%����H*Pm�'#Z Z�[��2�h< f�n�`�b��Tr�9���r�)e����ǲ+�
�v�*�1if;ۑ�[�]�L�z`��T�{�&/�\T��s�x���g;���Ï���mS����腶��#t��yR��q�V��7�$�E	�9�w�����v�(n,�@����S,��Dg2ɼ�z�Øʐ\����j���dT�X&Tl����l%.���ׅ����)e�he�'aS�"3I��(^Q��Z4�)Z�����`���R�m\.&\+T�*�3,����ί�3����{�b�{���J���.ʩ)��&�E����{�1u����-NƽP�
�ܳ�u��v3*�[��(���U��k
�RÂ�u-�3֙�{��M�R��#5��*�]	�;K+D�c��4�.��*�&����S�n�m�	�fS��G	(�qLekK)KeM,��JB+v�3z��N��[e!wN�1���αU��k�#�d+o�iM뢳��ʰIC[&��.��\��MxP6xG���\-_U�v�Q���师'\��֑����4��om��z���6kH��f�w6y�������Qym����(�fٳee�KU�A�f���$y��+��n��ҵ*��A�j�����H���t݇o[�W�c��Рj��YB8`"�O2���=ن�8��ٹ���%h�XPbF��o09���	lAb��R|�"�	�ȥ�ܧ��b���,��{�6%�k�/lr��% �ƈNb�S�m�?7>���<�xJ���$�4+�&c�ؗMGYD��u�n�6+;���i��Z_i�[IQ�ycМ�lM��X�8lY.<��Œ��c*�c�!L1`ו��ڶe�u(HnZo5�Xn��C%�^��[6��i@�
 �%��9/f�,XÀ`��<�:��tB;kC�|y�4���VVXd�U�@���Ϋ9t�ˌ̽ts�ൠ9O������۾�7�uI�l�yY������*[`ԽH	��ݧu�#�0ٲ�=gq����P��^JXY	H�������l�uwh�Xj�CҀ	�ѣF��駣0حZ���FcS9N��r�N�#��$.���H�0<���]���S%�ƴ��D���w%�n�W`i�J+�m��#6,�+�X����O�M=�,����E����2V0�AC/a�ꄠ�/)��,~�'!��H)Gxn�W�u�l�t��+4a�X�t��t�U
��F3�V2)
�qz�$�y�I0��F�d��q���A��p�_C���8��46�[�rļ��U������u��נ����/�RQV"
�v7 l6�
«6���V���v����F"�F
���*<Ͼ4W�pU�dI�Ae��n)�k5���*nQ�v.��!��=JyB%�/ �+�<�XM*+F.�� ��F^�>�a�$:+`��@	�`W&�-��oC�ѫ���2�YZi��nɚr7$٢�ա�.�p�ʕ�\0�8 Zw[h�F��Ǡ����?R��u����έ	����&�t����jM8�}�V\4 9��zܺ�,h�5X&=ʸ�h��1��Om�Y9���ׂ�,ّ[xt�x��R�/��Ry#��awB��j�b�S5�X#2z�F���9蛻��F�|��������u�v�ln �=�!x�[��i�֥��U����Ƿ�������cīSAC�a��Uc/��̥c��ߚ�C�xO�J����,|~�X��W�a�UK�GjX9d,��1��d�#+s�R�[��])�[�	E��?3�J��Qg�aD���@�*Q���ŗ������֪���ܖ��{φwe���:��3r�Цd�uS��*�
;��%̃fh�6ō�51[t�VSM�7M��Ӹ�F�U��
�L�2H��P�Ĵ�Ļ��-.֒����͗1f^���{��6�nЩ����v��f���3kYCyR�X��lI���We��%n`/��Q�����:��Ҩ�	Մ��6��'�V�q�2�M�m�c�A^��5a�0嘎�WЦ���ͨ0#�3��/w:=��=T2�YB��^,>�ER�5���n�$*�ԱO�K&���;͙Ck���N7���LcPgUfVeͱ�r�-q@������6��v2ޜ�Dв�������w�1Zi�f�sm��wjlō %��Pv����\�f7���y��å�k<�Fh�f���
��K��Lk��c�'-.��u%CR� ���Ne^İU�T�۷�SG�/0���I�*3��Yu��l)&cj�e曭܅�k(�*]�,��e�+(�յ���<i�7�k����R��dQv��A��sNM� ��?nm�P3��(�X(ۣ��;4`n��dg�}|֜�WZh=z�H�X��i��
��ݎj�]�^��E��*���l�(��|�7�Z�m&<$\r^�$��
� f�Jɮ#��6f���n�[��G-�;�
}�}�̱ȄFP�v�A��g �R� �Va�i�z�1\1"cK.޼�Ub����rm堮�C"Cq�A�t�k�v� *�H]�9�m��-#��F�^�AI�8y�*�]{@�����w7ۺ�,^�k� 0]�l&,��Tہ�L�ͅ�*�^V�~��Dg.�7�S�K�p�.��İ�	��Lգe��]��1Kٚ�q莳��t�S$f1�#Tn�j&e,ߝ,W2d��@s4[�b*b	[^�,Ӗ�@���G$�56�k�n%@a+� �`�t�z��p�J��kf�
�dسI�"���Eܑ�kr�����z��O�� O~��,����.m����T�[܆7(k���,�����]J��2s碆�ĥ�e6 u�آ�������܍� ����"�4�˫�Od
0��h/�p���[)+��wjb�oN����.�
�L_-u�Em�z���w�-�7W	�����u��XVR�(1��ǃN��q�"��g^����5}L��VG��
k0��ڂ�]晒�����T����>���6���ׅ�+$�+w..�&�Y[H�����:����V+n��:$+n� ��5����JhH
�����hJe6�n��x�Y�98/uj�M�̂�in�<Vat>�[J��ezkR��+ 1"��*�f��Z�%fSC^�`
7�/lAޙ����+5j��,�G���{F��[CJE�k�ua����T	���R����3Hݺot@Q%V��츱:x�h�̷�
��Bi�y{��n�`¶��Hj-��[�mf�f� r
Ŏ"&�#@TVĲ�Q�T�ұaS�bm0xPx�νB��0��V���'v��G���A2n�Z�1�u$2�(��Q���%�P�8n�L���s��FwWw�1h��EI�Y'd[aIOl������u��w��Ӧ��#���d��˻<s�Ȫ̥G3Y�dP���-U��Sچ�3��6Λ�u�L�I.��|�Z��40�ڛH\&ak/6�l�V�:*U��5��bF�̳�K<;&PV)A��$�ER�u��߂�[[,�cE��ӵWF|u�ǚ2��X˩�H7 h�P�˱)�l;�󼎱�:tm�FX�MP�B��F�� \N5��QY�2��צ�Е����',�V�4u�l��2IQ��R�]̕����tͼ77V����Fd����V�ۀ�HB�h���5F����7VG���tlR���8͝�e��h-�đ�"ݕ��MGU
l,�AC�ݣ�ku�G�&�6��Sb*����sj]k�	������Ϟ*�H�%���+��	��n1e��CG��^:	+�Zo��D2�IX�u�F�ͦw:��+����F�+J�����Ț�"��C;���m�Ҥ�cZ�\/Pz�l��`N+�R���f��:EK/^��z�x���*�ʯ�^��#i����j|��ßG4B�;n ��(��ՙ��C��k7wD�򉰕Yf;�Ko��fXvv݁x4��#�t�D& N�;kkvҼ2ݼ����W��J%���̙� ��H��� �VU=F�T����6��RS�pc�!�SՖ�1M�V�Fm����h��n�v�`Su3t�!��<����l�)Y�q��5lcz69W���� 9E�&-��ȴ{L�mS��d����n���h��]�w���K��q�{@�'�Wڭ���u������1�5F��)�j�nك4����(��ỬW�c�W��V!Z�m3�]��N��H���әx����f���$��;�kw|��c;\�
�|I�$�v�Zw���o�ýݍZb͊%�·�鵅v`��t�v�m�%d�,,U���^�j�(��.�&��7q����1���[OU�F��R�9��<U[�Yo6���=��H	I�B�ͼ�͚lI:q���ߜ���<A�bjA����C�^^Yv��p�i�ѭ� H�����0�� �y.�1xV'�[wV�c�.�)DS���&�J��iڢmŐe�ז��������@DV۰��<֯��D����RT�j� 8D�6]����͢�0�9�6����%���c�G"Ssf-{{G'*������أ�D�A7��H����M��eh!^M��k��ju"�]��\,V��iͶ(g�!V��a`�҄��_����Ar�����9vƍç�]Y���?��Rٮ]�]�G9�04��/.sJJ���,M�1$䧏)��se+���� |b=Y5�D��Q�Y��?n�n�핻{GY�(�<�T���;ޫ3i�RF3.|oƶ���(��� 6���=���@V���TW!oEfٵ�n���G�v�r��q�Z`�-�V�9��������c_>[�s����9�Ǩvm�#�g����$4�7���,}t��1��ܘ��* Ūw[ۑv�zH�D͈S?1z��7��x����m�l��R9H��gW��T.�r�ƈ���L��]��8�9�_OX Tk9Ex��hoE��� 6⤷���+$E�cKx2�&������t���[�������w���9V�Hn��
wX�Ǘ��/�Υ��J�B�pD�Hq����j$k#�WCQ�������6���y�Y��.@�G} �ͳ���d�J�2*[��׊F�谒�+u��Axz�Yt^5+�VѨ��՝*�ƃ��;��4��蝜Qŵܪ>��v����c�U�4M����eL�������'dS�s��N�Vև�f�U����C��7�$I��H�X�C*��q����&*\������%da�.���l����>�N���4����i�8�<�5�6^+�eJ�Dӎ�S�]c�Xs����D�Y;�����!�D����:���Y/e��B?�N�L]���4`�f���499�[v
��=Y��9J;�V^���]Hyvu:]�i�`T
��9Mi����x�+}Xw�r*�ٽ*�>g1XD�u;�şY�ʽ�7��m�2�7b�fޓ@KP6�fj�++p�J��U8��.�XyYٰ*b ����)-��ȓ!�@n�8r>z�-�*���'*�&�9Y�K%���NX}�
�$Zlmn���6����r���H�m��Qt��:�h�֢����Q�S/(-�אUt���a,�d�	��U��e���G�]�/�<�C�0�V�ьr)�5�Q7���*[�,ս�YFY�X����?�j��2I�`�"�ʸ��E�Fn#�-R3/g}1m�e�ި+87�V�%���ɶ� ��c79�jVVM��𥮻�n�]uz*n���"�U�R��f�}p�ږ6���4��́ࣤ�������ۭ�(��Sc[x��MpR� �A�g7�{���;*g�'I73]G���}g�9Z�U��� �@��O[ '��S�s�d�v9��F�<�1K$3Q-������Uw�iA��Q�qC�Vk���$������!�Ԇ���p�v��eDB�����+;w��N�+~|]H:��r�]��L�m���څS���[7�WwD����;m-�D=�&֎	u�r4u��{A��mj�{�v�94&��w�cY��+��uu�[.����B�JvV�Y���7��6�-m���N��@�����=�0n��wϪ�2��&g�F��m>4X�V�LJ� �UĂ���V����ʮ���;����|�C|�<Y�~����u�����G7�[�|�@[(A��!6ͮ���*���:Yi��[[ܙ���a�K5�c��GѮ���tz��N�M��g)U�3��o����d�#ނ���˄�쮭�g\�7JM;n�ߦ
�C�j���|���o

��;6���ZM�F�v��zƪe*<9��u��j�.�X����輻�6��v+7�̴H���郳9D��X��	[��H�;��u�o�)=Z�؏oe���=���#bm�"ަ�3��L��0�4:^��؂��"��m8lf�R��@�S��Ʃ�7��Y)�s�0�8��5^�w����4{Y����A�,W������8���Ƣ]͒��+|���,��{xZ5����I��F�S˭��b�J��cx�Ŋ`\�K:��Ϸ��l]O��K�+Jjr��{dK��y4H.������Z^��} ��}��iͺ���$s-vjۭ�EKLo*U�^P0vv��84t���g�$=u�-��ac`YL��5@���AB�ܓ�u�9ݹl��7�Y�i��Wz^���6����K嶛s�:�=��L�n�;k[�W�xx䦵n���\��,9XCn�o'�Cy�iϱ1*"�Ʀ��pXur�V�ͭ(���,.x����n�P}\�����2Q�|��7�xv�GI�����%��U|��q�[Ձ9�����'���ĸ
�_շˁ�&P���]��7տX%���-k9���E�o��ͦ>�uD���YDn1S\��q\�_f"e=ϔcz����fm��{S�,��t��K<��)���@av�U��!�TV(]��.��of&�	��W9u��t���a�9�0�J��52���o݊J�`z햯��Uf;�	v�F-�0�۩F���(R}ƳH��ǴmfA&�����/;.���n��^>ܒ�[�YL�n��g �F�z�JK�GS�.���\�kBLL^��b�iô����]Q����HӲ��Y{kl��Kt1z�ڷ]�e��X�tcG6��qn>h��ӡ;��]���,�U!�'bC!�����m[g�m���8�,�vU��qԗ�k'v�N�ͺU[�B�]�����b0{(�Ց�C�	jƽ�ۭ�k,(ˈC�ʡ�I�I�7N�z�Y�*�!\�z��kguga�6��K�����*��S/aMS3аK.ZE�3��Y%���&��=r���M[��[���`-�̹�*Т��yy�q�y� Ք�h�P�e��t�r�y��ҾZh�P�-&��P�[t.��-�7|��l��qqץE-saea�\Ϻ��}{�m^����'؂5o�<MZ^��s�0��LO7t�f�wC\�<���]]�o4�6��l=��[]z��rA6��'(fL4��T=1������GU���'�[n���f^�[�>�S&}����_[O�K�%�b�$뫹$͡E����e���C�B���Vr��7	ǢTt5v��@4�^Vumn %nS:�%�{�\��	+���OPBvtY���B��jԝ�J�
�h�U�0����l��f�l\�9��
��7�.���)n�r�J�@�SZ�W�7�A0h�ˇRl�nA5i�E�3�_\�L�=.��Դ�ⶅ����a�/��ƜĕF�;/Ug�h���h�m. �蹼v��꾥��|�������b8�9�F9[��0�[Ahʊej����+Ν�^��CcZu/`Wd��V��W.L�����{�(����*CJf_!wfۗ�R{S��7�v+�6�޽�0�m����{��׻$7t��8!q�nc�n���b����[��MȧT4�i���}{w.8+����7�qh�����_n�u��H0�헄Ĕ��Mg]���H��/�����A�(�o/13�v�o�HYz�Nc\Bڹ.��][��B��GD��c;�!�t�.��x�Y�3%$�fs��E�^�ʆ��Wli6b�l�c�Yn��rE(WK˱/�sF�-)��>+-S�[�TJV�{lu���@���[��6��I���Fѡud�r=p���巆�t�V��wa���]��[��fY� ����gjT�Yթ;����vˊ��=�l��ua�[�if��8�R��,�C��Hd�啒:�������æ�F���أ�	m�6nӂ���X	|����˃�HzR�ʈJ���#_T)��
܆�l��miH�H�d�26rY��!6��Ǜx�]^]b�����2L�'q�+�B����$�@C���v%�d�/����(�/7�6庺� �����tu
����b^Apֲ3�[�$�`fŷ5��1��O��&_�ym*|{��3{]�c���E8�R�՗�k>m��vW<�{&8�7w���;��Y�ݗ1�c@�uH���{�1��:z{���k(v�^���;���Ⴍ��ƺj�x��I��!_)" R<sT��Ӻ�U��D7����Sc�`^C��)mgU�Nܙi�7YB�}�ђ[�gV 7c#t��ܫ6s'X�LV�WQ6�]%��ʱt��Yw�]>��Dg=�!��YD�3��4ε�(t����16�����s��
���4�ޭX�i��2� %�.���N����⧝\H���5r�(L��`ĳ��h�ٜ;1�fZ�ͭ�^Њa�\iR���F";�p��(lx���5�.�OPZ<^r�����Z VGs��g2$��]FZbb�ʆ_e֍��`�q:갷�k��z��mu2����t�H@���,�m������Nh-��U�'�8��z˽9�K��kg!��Js���Q�$P��^Z�V&�Z����q��V�@���C;n˾�ɗ���j&l�f�$��������۳��4�-bc�Őa�����ۺ�W-��n.�x�l�*R� �-�:�H�J��R楃o�q;��;�/*X$ej��+p]����U�����v��0��}֓D�ǽJpJn��wIcT�ų�'^u�e\�9,㇙��Ӛ�x�!x�����������6%+��K�Pع�swܯ|��+�N�������z$�-"���6l@=�t���W�r�1�I�w)�]�F.2�4"0��,FM�ԨkjŪɕ�."5]���=`u�<�gN����hm�7hm4Wwױe'��w[�Q۟��$y����PkM����Jp���N��=k5�JIX�e�s�jB���tB{�ĻH�ɱj�;HM�D��Ź+�p��r�Λ�=*�X��륇X�΢[2��WF��pg�]i;�&CTU�ٹ�5�"�4���l���%���	�p�]����z��y����q�'ub�9zz����[�F�Lr������e9��<�f�;N��MKM�{yx:A[F�nh\�r�4P����\�%;C��2�:;;�n��JVstji;���`t �Z���r�w�^��4�;;�F�\z��*]�>,\�B c��_N�Z�V鑃e�fWlĹ�M�j���.u����5hܺr��KY�Nn�޻cV��By��[��H��k4��)����O�ʈ����i�5*Vc&e�ʻf��
��2�J[n�ӯJ��n���/Gt眦���G���}Yx��F��7I"��	�:����L����P۵C���:٪�Uz���KY���V�P��Żx n��mh����2�k�+Q�s0�5�kȢT����±"����]\uY�@N�����j�-o�k�})h���5���8����"gX�p��Õ����P;�{�ģs�q�`��S3�S��ujB뻕��a�̜m����A�Ɩ�$)�}��vʰj��YG4��k���S���>�s4��(��i�̺E98F�]e�Z��۽���&Ƀ[�9XT�0����>���QA�
�n���0�5��Wr�J���ō
���1�gj\�=��)�ݘ"�+�+(ޗ�.M�o�YL�)	ضVhY��R}>���jǽ�A]���8˷�ֵ�N�ӝP���|Y"�V"��ٜ{��fF�����U�JC�u�I]��v���	:�~�(,�1�[m�1���՞�F��Rui�&҃a��փJ&�O�;.b趖�)gMi[፨	�[���}	^k<���lBX�S;t�\��+�����7`��ʻT]Ϲͨ�5�w'x��A�qU�vn^�1���j�ud7���P`|��عW;��*�v��5���R�u����벺�.<��٪�o��]i&Y�R�
�چT���P+d8)>�SW���L�S�) I|t\6����]a�����>(f�Uv%���iu��$��o0:�	}Ѱ����3��K�,<Hۃ5�ٖ�̙�F��֏JݰA&�ʙVOe.���)�%n�\�:��S��T)J��]z��K�X:��K�P��W��p�%�2"�OL��7
��ݓC��M���dW�aSU}]7���Y�!����9|gV���
Cc�f�n��p�K����f\]��ۅ��׮C��@�p�Wpm���ޢ����e�{��@�/�M��{�R4�,��Avr�B믹\�Ml'w���r<NQ��׊�4A\6�lv�P�t�k�[@S;p�:�	:�(1���'6�83F��s,�G��x�gR��(ew+i�6��Yj�Q�cZ�Zz6U�����v�}�tuˍ�v;��r�s�9ي>u��O3m�����p3Y)]�+��]�R��%�d�P<3��xt�@��h��Yː��o#�VbCl�`&[Ur]��[���U��X��Tѻo�OR�ܯi�<}�J�x��Xl]>��Esj�o������Y�FUX����:��k+�_�Sn���.��p񖱮��Aĳ��\����/6����t�h+2�wVbٹ�Xe�f-4�X���s�"YՊ\ftnQ�%]�^K�%,��p�X�5;y�q��@C��u��\�U�,shr>ug)V.��%��bn3+n�E����K���M�!i�uΗe�6-�쇇lO�Z�L�QWYp���\�0zwA��f��[r�Nq���zE�gؕ�G.�k�[�Y�7Ju��ig]nԼ胐�*To�O9}Q_V��Z�c�q�d��`�L��;�﻿{�������}�~}���
)������{&W�[�~V�T7����7���Yt8���0��bGk�#/�h�Y{�a�xB
���pkŽ��Ѡ�3�H*��@am`�}7BVS;ڛ�v:5�wu�3Ul"�=���m�}\owyH��1��u�5d�5��8�ޔ�������ȵ��Ws���ϊ�H��u	�s8.�M���C�q�C:�k%���<1���JT�a��J���0�J
���ŭ���]
 X�tf������Çy�,XC0�8L8f���V� {��)�,˱*9���U�"o�T�E��.�Ǉ>�-K?�6J�u!�i�Ί�B!j�c����ș������oq�ɭI��H+�t6��j��pW�x��۝��e5#���o� ��n��8�;3�5%��N2뾩P����W��6��m�um�.�4��[�5��7�qWV�Er�˘3ll�-�æ��u�v�q:(J<��*\��yTq��`)�s	<d:�Npe�Ź���!��7e�f�l�g���6��n)T�=�]廜N�{�o�R]�;��Q�b�������ˉVdk��兡>`|ė�6��K�]�͹NG�9�;��#h�*J΢�5�;i8V$[x���6T	��uw�7�Nމ�S7)'��p_�w�r�fn"DN�L�*p?'wTz�.��vͳ4p����W�:�T�A�ږL�mn���%Q�[Bj�y�Ruް]�[ã��î�v_n;�`�cU�ѹ���L|���m���Ҧ�E�R�3!cE�]P�uԸW;ו�B4'M��>�p�6q��ʜF��ۡ��v�Ogb��cU�iS2�r ��k;�͍&�ԅTgk@�L쬋:�F�F��7��o+�6khT�A�MF-��q���5���!Y��R"��"8��;|^R�/&"S�� 7�b�ތ�1M�2�k6�`��fL�|��r�uʦ�/kC�g\Uv<�낾��1�ML�0��>�M�c��HK��u"�oHp�M����\�(�HU-����]�ȃJP��*3*�K�c�'NLò4)`n��C�[��)�ɗ�,�5 �gn]��)���:f�opZR�A�U���`ǵ�eq2e�koh��V[CD��A��8*Nx���%_�*�D��=�P�w��kܥ��s�[ Zu�����Z��S�g����][����uuq�Zd�{fʣ6��ٕ�"�^n��J��)ݱ- -��{�������`��`�x�j]��#�e	��!�k��,|{�h��e���|OS/�(�i,e�h��b�����m����n�����W]VM�B�5��Q׮�W�w�0R7���F�Z�
\x��h��m=qJ�m�gq�B�y�Gn��'�lm7]�rK�7�\��c���vi���m��Wy��[t��u�&���I���ߧ�+~r^id�h�{�,��2�m�h.q<L����D[���xO|v-!֨,nc�Jgnm��M(��[�u(�ó� �DsWwT�u�2�v�+A��A�,ʇo�Ƕ�]�������T8U�*��� 2�_ �2��8e�~P��&<�XT��m�D,��雡p������Rp]](�v���u��40LX=����wa�y��`����,÷o�R���)�Y��mV��yzn�ü�͈�5����WR�	RU���f�vX�%Ǜ�I��9A,���X��t���Q�\6�F��`ظf"�����Y���=��;!7�F��������M^4,�gv%�n�a���|!F��c3kX&e>�
XN\i���J�����ZI��"�U�q�3�k%�ܰ21��[e���+���S�^��bX� u�G.n=k�#1�Qv��7]�ģȉN���Y�f�p��U�8�G{�Q0�l�ݶ�9=��s� �r�N3t�2�Ǒ��e�!�]"i��5�剾�����8�r�8�M
Tq/���Q(��#Wi�2�\Qe�|;;zb&jI��e;�Q�R��`Z{7�9y8t�)��V��m��;|��۲i�^G�,��+�����8�{L1�ۛ�ی���F�-�|�T�3A" ���7�D�+/��EZ�܏H�T��YC֪@���a�`F�,Pd@�Dv��h	J�=�B������wk��>/wV�	W")��4�br�"�����)7
���[a-�k�u�\���T�-h��t�Χ;̊����*e��,����	Z˖�ƚ��]��k3�ͣf9�J{
�x��V��q�gh�(�����ļ��S�u �5v�<
ך�Ī�b�АYc*�d]�o<P��J��RϤ\��Ѝ9V	�Ǖ�Q}[�ڶ���`�Zl6�9�iU�܈J����	��T1����G
24�9h�WnZ�/8H�/3yP] #��W���f�/��ns���J�A�;tQ�#s]t�k��U��*p���r�nfڝB2�T����WM��	�V�@e�Q٘6Q�:8��Tr����$��>ۚh����P�V�]�;�4r�,Ma�j+b�<��eX���Nb����������b�y�Ľ!SR\������V>=[U�8����jԫ�c�$�<�G͹e�n�K�|{N`"���̓d�W��9��G�y�0m��c��'`�96�v8��9,+�F�u��Z^҇�GXs��<�J��;1�u�`tt�f�Z�	قH8�`9uy��y,#3�3�P)���m���k��zy�]���X��؆�w]G��7%���Ά�_�@���."��Cr.��*��7��,q�����Y�DV����3�l�`�݁�����m�	ưfx�^��n�� �$n�)��
B�5��\˷�e+j]�J�.��J��e {*/���xB%/�1���f��V˛�ܨޑw.5΄��6N�{Z�
VM�f3qG������`t̵�r��1a*�-4�y�9:�V�<�ʻ�!x�ۺ+�й�y��~g`�Z�9-�0�	��*gf��I���*�����q�$wv���@n�K�� �Bb�}RV��e�s5��н�3u�Z�Cv@o>�z��rc̟4{⌻���\Ĳ���V\O�kq�Ov���C'W��L������v�R��D�Z��aj��w@wM��ld��92�M�� F�0m����K%�;�CU2ܺ�Kw/<8��Θ�o���'���ZHwѳy�(t��Xո�,dN��3s�fəө��o��3BShJ��C�j7h��}sL��MJ݀��`�Z��92s��:v_v�>��(`W�R[6�wdƤ}s8�U��&�
��v�)yX��	ux_�|s+xK���EX���WŞ�8i�ܻ\'>�� 6'Ww��rvԫҀ�.�����0!�� &���̈́_
�F+\1�[[�r�lƼ�I�pãz��%��+�ځ�ґ�Ɵ��a
����a�I�U�A�i:�b�M����S9Jo\�Q�j��95Z�@�	��
á��;�� ���ũ7m��wm]�j��@��e+"�UbRĚ�HӻY
*�Z�7H�̛�K��G���@5�����9xs��QC
'�<���@����̣t-+�Z7��V(�x1Yr%/�S9�����p6Y���nP��4��>��L�<6�Jhw�Z��&�nö.�����TV���.+���/�QK���뢑��j.g:4d$@5�΄h�VPN2g%��[F�\�-m��Ƿe�|Y��Վڗ�S�)\�ڏdƬt�#`�Uޥ{��gXQY|�uH����s��F�r��O]�{Mby]�0���y�7+�L�,&��%�![Vl�]��N��A6����X�t�-�d� �ͨ�T���.��jO"�)*	�vJ�E`�Ӳ��|��o,-a�.���dNؾx�t�8��@%�[*n��U �H�e`�np@H��@h��:�m^��s	xi �ηL�Pەla��j���ߕ	ݸ�s�W�l�� �D�4�>�l�]��ѠY���tŸ���R'Z&sAH[���1�.gd�����P�+����5��d�9���X���둮�
B�m��s���p����n�np�)�,�*_)u��W"�pf�^�meq}o����,��ު���+rJ�z3g+;��k��]{I��4��mwu�YV:XN�},mWW]d�7�8U��i]��T�[]X��K�cqB���D�_v���Gj�況O ����-�, ���lRฬ���}R��o��g{4}
�we +�2Rss�"��B�E�����>ph'\���݂������Wy}�l�f�#v^�0��v*Y��<.�O�=5w�옪�%��>'%�v��P�=��!c�8;Ud[�{�ʸd=�R��9�,��(�J�S��uֵϷ��/"� m� ���YVFm�v#�r�ju��X�_l4h8��z���x�CѦ�H;ʒ�[�5�7stʚ"X��ܫ�`g�=Z��[w)��]��o-f�N�@�D^�|�[`�)Ts���d,���EҭM#c����aF<�/��P��l�iN�V�OR�Ei�q�S�q���Gvfw8���l^���õ6��)䦱$��Mkt��YH��̱C���)ʶ�R�غa΅�H�>�)���/�h}�-�u⹣6�`9��ķK�/ �*�P���B���K��:�f����,���:��(F\H[;�ӫ7�n�$��u����*a˒���[]�D���E�����[v�{���:Z�v����E����k���mh�҆d;�O^&��X��x�޺ϑ��^��ON`������u��t�xl��t� S���Ş����Nqg�[vڔ�F���t��,�hʍ�t��+)�6��l�+� ��t�
�;1� Dm�õ�X��с�u��wRlf$���]���5��PX�*Ʒ(]��3����(Hz��	ʷ_e����Ǿ۩0�1s��8�U�p�\��c1��/-J��}��:��Wai�AZ�PJrk��H����6Mu���n��M��Q=Z-e�-���9�ޣ�X4� ;.���qǮ�LK����G��Ƕb�ל%�w��	۴1���ӑ�G4��`�X
]�Op�ˍ�w�a!]q44wR P���P�XOV�z�����$����Wux�,��}z�bN(J��0����t���\�e�;3��V�%�����%�K6��Ւ�7wNb���,[C�틭�ɔ��wFc��g^ۡ>��v�AzdM�.�]x%��xR&��ә|�WOiN^ 4����Koh�h��X���}�G�VY5�E�A��b��=(�;�F �e%�;H�ѓ�TK��h��u8 W�6`[����L몏��� ���.����jH)�r&f���v��a��ixck_NBձ11ε2�3n��t쳹qd0Srm�P�EegY�w�J:(�$kf��]���;aD:��e˷���36�a��2r��_(Җ�ːd�@+1��i�Z7��2Sg;��/�^�X��A�Nݮ�ς���2J݆��.��w��qmeY7������ɈL��|��d]�N�th�Y�!ٕ�Vub��Ψ ޠ9��G
�g�����*�Ug@|qC�GUe�u��ͱ��e��M�����=ڪҧ�yj�m���(i������PI�]�+�s>}
i����:H�X�h6z�j�\72f�Cn���
Ɠ�V�}���_bw�ݞ&k��UڶV0�r��[},�Mo��f3�J�.��+m[�o��k#�e�g��t���Q˲��Tu��&��b���k!��c�ۻ!��T�i]M/R�<�0|�}7�G�V�Ӻ�-T�*[�̼��f�Wm����fkT���8Z_>���J�b�7�˱�1_T�.����)ڍ���8Z��t:�o����0|	v4�l� "4�������Vڄ�aގ�W�>+�ҕ�J�
�!���ؾ�b�D���h��EL�ϞR�ܷa�����A�� �o�nY�{�R=�I*��и�D��L�sX8��,я������1�X��:�Iی�k�R��Ъ�3[��#%-4+�>ʰ�9� ��8����U2�Y�Ե�����ڃ%t1��D�J�q.c[�;���Z��p��Ѷԣz�Cz;b�jg�v�����X�1s��=��=w;D��Ky@K��S�2��m�P���'�{�p�$[ò�%N��ѥ���ݼ�7y�S;���B$V<؂���v��7}�"݅�Caa�F�F�oe���d
U�B��5�S�!�̅�x<����wL��؞͞��%Vf�vLa��X�������;d��$v�l�@:HK�AR��Ϋ�ܝ*�b=֊��V�D	)���7X�*%���}�ws�`q����6؇[��B�z=�jG������<�I��;�ٔ�zԛP"hu��e���l�ڧR]��tu�Y���B%I���ڎe�*�؞ݶhe�.���1+�m��m���)��0�khMXi�n�O�C�/�Z.﬌�LJuk��Hl�vg^���d')T�Y��d<���J��A��qV�\�(�ڡ[�+�1�5���҄�8���`d7\))HgW4������ۃ+a�"v(��3��K��Q�()A�h��Y�V�w�2C�9Nm=�_*�w+�-c�]�7�Ϻ�Hh�1��8*�p,�`���I].x�l�X��\�,}�|�8y�ј&��l'��W7v�9u!�iYUmPmZ�.�D�m�fJ߱��g�򦀆U\�f���d;T�ٶ׼p��U�9��&Ӈ�u�� ������ͥ:�ą�S7�C���+�(�`�!y�۩.��家��n�k<�f�a�xeFq��\H3y���c0@1��Ҳ�N�瘹B��d�*RWC/��y�`;K���մq�`kU��L�A� f�:~�#4��ڝ&+J�0�u.T���t5{�v��ٴw,'C�n�A��ql�H� u�h����tiCMu;��&��[�1�˵Y�/�vp�8�H��C_Z�A��5�VK���P�O�{ራd�@ܽA꾨*�|���ڼ�T�ͨ��	f&+�\��Ú;�h�Z�Ѵ�y#͐tt[x��ͣGM���r\��6�.A��v��b!��w
�pRy�>��:����Q?��Իn���q�Z�f�in��u%v!�nmu�7�X�K�uh�Z��+at�]^�L%B��7j�X��������#Ug��{�WIz���oTA�B����fV����G�<�_76`;u��U�����.��e��=Q�ܓ�˵����wƋ����.(�[rn�RoP��j�N�F&�e��%{���(l�" �۲7+�m���Kӱ9�:�p�[ͩC�|�/Gi�q���B��;��K��Y���s7� ���D�ݹ�� ��{�7)��r�����e(�!�qU8q
]�7;s��57�f����\7���+���8!�=f,�nv��ｪ>��,�)���!�ʳ�p�q��«#2#3,,̪�,+2�(�"")3,��,���2h20���333,��	���`��(�
r2�"a���3*�,��0�����2
L���+12rp*0̘̳%���*c,,��*�&*J�f2rj���h��(*s���3
`����32���ʫ*��*���l�lư�	�&h��(��0���"�
l�(21h�̗&���32H�22����r�������"��	��"�� ��32�b�
bL���2)�%ʖ���(���C&����30���L��p�����Ȣ&$�)ɠ�0�%�"((ɬ���b�}�k����j?{���[�>n��ċy�fc���0R���q%*�k��f�;(��&�E:t���v��^ru��ց��/�I�����p��cV�{��}k��'Dî��^��ޒ ������oM�m%�\# '�7MB<5,.���<�*��G`�d�A��������V�r8��Kt�v�����Ǘ:V���°���ZE��s"�2ꊾ��5z�;�I�]�TS���4��x�5�Y���S�!' M�]ƅ�E@��V�"@	;7���j�oyi[��'w�,!aՑy�k#\/�;�	.Y���D/������=�� �M�癚�^\��X6�X�@�t��~2�i��B�36퇱}[e�\�.X����W��A�^MWQ�3�&�l`y1�L�����k��K��o���8kY��3�����+i�Ȋ���:�q��1�]�����T�F�&�#�L���.b�ո����_���X&��p3Kd�V��T/a������G�y���=FǦ'�5B�:N���,�]#v�&�F��\��7�Ѓ�T������`��ux������8�"du#���ǂc�pu�X���8w>�,+��_-�R��Hg>g���
H�@�yDWkE1�X܌X`Z��X0�f��ɧ8�|+�K�	Rj��ӱ�ww��}�;���4v��V���5���B�M��S�(ZnǫGe�엾��v� ��Q1�(2j�e���C���%�(����t�Y5�o2�j��0�֮��sbxQ�(��<$���xK�{�+H�<ϧ�ɭX�\]�;�Tl���n�x1����P�W�И�2t��!E�3~�(;S!S%�f̓�S~����Sy^���Z����<�7��r9g
�C Cs&i�\
�҂�v�d֬�Ɠ=���o�,�y(F��xZ/����ݟ �����Sj�댤0���32�6<g��1�K�/
0P��K��F.!�Q���쀥��e��K�!�U恗�6��Q5˳@� ��K�Kg��U�o	l����4��nm�XR��j�v�Z���K�,l70��]PaX$]P�[	3�g�
�����<d�������F���'���c�]g��n�GBt��uLZ�8]�'��|�֪�(����8�}���V��Iq��A�n�@����s��5uLt&gڀ�4��|2�/��8����ށ+��Ku"#8���(� ����~��7��9}�ˈV-��ᥩa�1��W���"��I ��k��a�]f�ku:���Y2�5
�7�t_d.}x�}�w|&�Х,�j�XD�&'Ѣ=#PV�b��gG/�d�V�d`��u&�2]����8�ڶ@�a��`�T��J�w�����yg�KQ^��x�}�k����o�-u�����Xϼnf�=V���=�ŉ��1��a�5:;�;Κu</;��j�U&�u��"�Z&�_�q���unaαT�_�\N��U;82 &V�2�"�q�����I"����6*�}�a1Ғ�}>K�	sԩ}�*�����)W�94Z����O��,�|����5T�fD�ގ�4Q:%���w�	�X� v��M���$�ب�`�Rx�O���i�hTj1(�؉�@�}�uKS)���X��3ݸ�OZ�8ڥċ\&�{$:�O�
���x�=�n�^�V�������"�t.2�̻Ck�_RF���qR��p��Ӟs��c�#�)ej41cW���*5��+���-�
e洈�V�L!�	L��.��
�=8�i�L�`��o]�u^�?Y���$��N�l7Z��v�q������(2@��p�	���
�#�^{ΝƬsW���*yN�H<�����с�_;V�Ź���>��1P�E,�-�˩�jo��ۙk���Xg�i"�&U�m��q���0�}0���tf��	�Q$�'�"�����5}6�'
�l�w��"�ܺVb��-����V�����9G� �瞯Mc6�e�b�D��.9�D���hB������~;��W��┎�̼@���]Q���q	ȣ�i�>7"XtI7䅆��ML��P�a���gv^�.k9-���j����tI��
��P E���a�uP�䒆����}��^#�^q�2��c�ԯ@�N�T�C��䃉����	Ġ2��C�9y��Ai�&h�Ƀ�K�1n=+a��E��]D��0�-#<~��W���"�5d\ei7}s���u�u���)�={N�͞V�V�Xn�>�1��P�DV�YQ���� �v���]7����Z�L�-�R�(h�^㡊�Y�UJ�|�\{�nD�{-����ïǡ��1nO.�8��'��8q.ۦ;�ŭ��`�a�R�&p;7�S�ժN��ۘ3�P����joV��b��;(;���d@N���ax��_:ȣ>,V�\_��>L:
Ϲ�n1rŪ�X�H/�@�V%"E�h��{,G)}p���xkBu�w,u������h)�3�%uy6�4O�T��c{f�۱ Q����L��r�zp8��R	x���p��\����M�n�Mn�ˬJ�nU�T��R!�jC�ჩn>#Ns�ʙVJې��_.������8{.n�1cES%���%cp�.ܰ���r�E$��,��U("�D�-���C^�Q���{
��7T�<��UB5�c]��en�p�\�H�u�s�R�7�����Xw�J%�;�MR��lU|�[�3���O��#�WJ��k-�{TT�;� ː�79��>�ގ}����
9����*y��^�b�W�æ�(� Rx���>���'�#�[���9���@{���Δ1���''�Iˍ;}�^��
>֜c��/ڶ����/5�9�@&ZŠ$��&����C�w�S��Z�B�U[�:nڰ�EBp�+ɽ��s�Q��Z�Ȼ\�i�X=
�ɩj{/mg���s����'J)ۦ�':I���kgv�Q:������~���'`V��z���� $���Zѧ�Ł�8*�U�s�+Ԏ�K��gY����\��v��ˬ�s.��t�L|�Yf�²�ov���j�=���6!����&|�$���4ԅh�(.�3*}ݟn�}kgo��bDb��3�B�q�M�Ab���n<�E�lMy�ԃt�k�`(Tn.�����Ew:�u��s�V�Jqn�ڇ�X�58ʌM
��ZR�DP`=�VC��5��������9l����?�+P�}N{�3�ǽ�v���������>)dbOx�&"���K�����u:�)�����[�O^����n��癮�K1`/�J�9:;�S���Tv����w7��˺͛Մ"�S���2Hd�oI՝{#u%Q:�Tt��*!hl<��OM�s�fbK.S���{��p���y��/l
�%n�o��t|�R��(��e��oZ�x��)w����o��#)>��D�N�r9��Y������uoB����q<�|�[�s~w��5<�6Do^�<�w��W�\�%�;".u�JNk�8�����3�[�)v4T�p5�\��ݠ����zz^�	�!���[>�aW�b���u��oɺإa�k�K2"�1��N�vh���;�6~�w^�Q���k�#n��KS#��<�^�m����7Ѕb��<�zGk�;L�h)�(���	��Mpݚi��v���(�2�h-P��]�H��&پ�����&sX\����,�6�B
���w�C|��]�����������[U�m�@ɼ�[��]��/5'���Ejp��M�c�u���!����B���t=���Cf2��[K�]��3N�h��p�ۭ����c���w�aþ��X�omL��ʜ��P�	�MEBv�_��ϲ��GX�^ؼ}��Ef�m���|ǔ�v��[�- ��\�z�gܧ���OK���~)r��I�j�m[�������+��ޯ]9��o+z�\�I�\bhW���ݩ�re���)9>x=�7����ތ^J?L}�
{���nuݟRVA��72�^��k�܊y��\_	C°LR�������L�J#���xJ��l��;hrY~M=Y��}�P�T[��QУ%	U��ZΥ�hw
���s|�k5��T���07G�b�7�DcMz����XR:�o�];}�	F�>cz��B��t���!lR��1kuu{��^[辱�8�cM�Hz�b���r�tPZ�.�z+^I1ۮ�X����̛%c����3\ &)+e�k�����^Jj6�.��vf��.%OR��B��=�=R+�p;o�hʹ�I�����o�.�z��m�ׯ��0�^w������'�u�\�{	�yq�C(�"��H�	u9LWJ��yh���)}S���u���
=��϶�eM�|���W\5"+���<��';|D,]�+������*徵�l-�7Ds����i:ڸv�@C��Ӟ����+׳޺n���.�c�fG���M]Wڸ��N'b�7��wU u����h۵W@�z';_$�;^�)~Χ�=B����&Շ*+��ȨN1I]@,�;�N��Q����.Q~���<��%�}���MBp�s�[ŵ����b���f.�����C�q#���G�#�����gLk�	���U�)V^��hp;C�2�lE������W�evϾ�/B��;�}�!꺔�.*�Z��n�;8���|��wM$��\i�b�'�{��/����/���KE�������Z���Հؤ���K��1��j̔S�sDdb2z�ޮU���r�C0	ޤ2Q�M9��'�d+����'�eh��1��L��o Վ��'#�pV��~�D�O'�0��M�w��vC{]���]�7փ[p���<����P;�)*R��!&�[o�)f�9�Uu�͞����û7�oax̺گUB�����k/ɦ�"�ec�J2/>򞾷��ݎ��Bk����;C�'^R���ny��R�O$ﺷ4�Y�y�}��RKF�9T�PN�����ZB���އ1I밷��{tg�����O �P�;��UM��oն���:��WJAm���=�_���\��s�Kuf,�YYN�w���#s�Do5:�Ns�i�Y�Nގ��؀S�|c+�c�ҷʥ�UM�UB���1��\#��x����J�M�ع�D��5��i9��rN�!ۭ��n��)T ��l���75;��yj;׽;2巜E��z�M5a�ۄ�l_�=�w�M9�oO��}�����HD��7J�� �V�󖳇�1��V\"le�Yօ�*RL!x�k]�&��8�?��N� �2)�Ř�����ޭ4!���y׬L��`��Vc�����,fm�UkK���c؃�h>hi�]n��	^��
#�{&
F)6���#C-��K����K�Ng۶�9P�+��3�/o{\2 �^�\�ߝ>�!�WmLMn	);ޟk�~��6�#�/I4��^��r����X����Z�\���冽9�J�Aw9\�N㒌����j�h9+��V)�����b��`�����+ҕ{�����Q�ҽ��ǌ��}����<|胊_ъI��x��;�^z����}��|��=�N��B�m�ܥ�J��D�чq�V-��M����#9��Ux�	�sbTWf�.u0��.ko��[y0&���=����;%�b/N]Zϴ'�k����Z�B��oƘ0�ԓ|�s����wӦEW:����n��	}u�P�1KCb��qu����o�Ft^�B߷���O�c�Q�T00(��T���?x��� P�p��A��dI�ݞY˭�F����dKڄnE�po{*ـ|�X���իg]�U���s����(��lt!��t���&��|-q�j�iP���wZ%�ے�'|2�	L�1����8�֗n�GX�VI�A�/A�+9��
f޾{|�G��/>��������V�Z6��
.7�S׽��l�D
��+q;�9�����2������Ïi��<6��n�zn1��ie3�W1vi�zA?0�����XT}玲��G&K9�Z��v�ϒ�=f��O+�C��0�!�7�8eJʌ0�[�o��C��v��IFk&Y��׮�d�V���bI�@�0���CwǪ�N�%�Z�oF�n�An���"�v��Y��c;��/�_Md����.���y$i\'ۥ�%��+��6�ڡΧ��]n�u�:�]���������!_7������37���NΦu�Ӻj7�%�O+Uٶ���j��K�2ُ�w1��R��t܅r�=�u^E+Q�C��x�a���@u�p�c�e���ֈ������h���F�t	p�|0�	�[������TQ�YM#��B�m��ͺ�ɛc��H��y���I�|���,�y� %2�f
[[>hU����dk�UϱEOu�w�W�u�N���Ob+^	�A�p��>�oY��8Sk

��:�ڴ�E����J���f��X�͙��Һo�]hóD�<���v��e�,G��R���D��4�>h�wNnh�~���殺��A��O	�d'.Z�,G��ǋ*�ڗո7H6Kn�B�'�1�Ҕ�w:�������w��Il����VJ�+�j�\��D�QY��q��Wӱ^�敞��-��&����U��2���.���n�ocq�v��VF�ܷp�-JƋ�z�I��oto�T��Z���(^L8�%*Ŋ�g���Zr�:[R��tJݒ�ݪJ!K6$l�ÅfR��ba�V��A�DlwU�"
<h�Я���zq����Ti�5j��쾍i�˧�,v&��йr���Y�n]/��Ҵ�n�wMw���qHs�[e�ָG��;fRz�+�$wC��cj�� �5� T��j.p�an}�L9.�r�l*<���t�iv��o%�[z���eiv��6���vdg5ɯ:��	�Qx�ց��s�^�i�inI;��;2+o+E��%p�_l[VM֓�¥���h{C�`+d:4��^�ȹ���uE���"����Q;yŃ�q����
�Ri�7�Cj��f(S3���ە8�\���tq�Vʴ3���*p�jZ�5f��N9=�ҫ�/��R��*�_:d��l��{��u'��U�A���j��0�]�t>�כ�p���㮡�%(YT:�ێ���(���m��J���؝e�L��+���/�R�w��^䔢H������\��+ou9��F�U
��$U&A�E6FU��6!�LQNI�14��Y�D�UEFfCYUINTaEd���fP�1�d��EED�ae�TDCPUd�M1AEfQTUUEe�ML�Q9�Q�a5��Y`PMM�TT�a�QEEDMACD�TEUAQDCIa9TDfQ�5e�L�Q�1�YdIfa4A5LMVX5���MT1QLMU$L�TVFAUAIAUVbd��TSUMTTQ��QK1QFb�Y@EESYc4U)2�!DUT%0P15MUQ@SUEa�QPS1CPMET�aY�����bEALT�@U4D�5E�Q���TU31$D���FI�PДf-3SDDTE4�aCfd5M%@P�C�*�y�H�Wv�ŝl]a��g
�dl��L��ۗ�.���@�xf�li3du$�����OX��m�Ϲ�G c-�p5�~P��G~�}�m�V�-�t6T��
&��j�S��l�fy��9��?')��Q����-�MUrj��Du��U�w-5w��e�\�v-Dd0�Jx>��{h��Įv&����[��X$,>�����"��J%ZY�A� ����f6�K���o*�Y�zŽ����fy��4�׮�Cko�?���w�x���TT�9~ޠ:�u�d�^=�����^��a7���`�:�sR�m�Z�")���[@aQE�bN��(�����r�|�,��q��R��b�{aܕW��8�@몙�݆��r{J���}�	��JMEy;Z.9��eK���j��鞞�`~��f9�n�/+�-K
��ȷ=[��u���LZhRv�\s�5���!2�q�B�����`=��8t�aSs�.D���htx��_fZ������Q-S)k����C�ˡ�{h05{&�U�<2ߢG\�+͇�˾�}�w����!γ�2y��ZY"������M�ŷg4�,�P4�ٴ���We�q��6��q�����悶E���)��]�4���k��s��t(�ٖ�)w�8���č�}淪#�r��:��1MLu�QQ1����s�����^�Mv:iGq5�t�S��WI�6^�����k���|J�A%�dRؿR��Փ��V�˄��6�M�
Ò��pq�����'�-���{�p�X9���s|�5yφu*J�����-mea�f1����m+Gm���,��w`k-hSI�kz�h}N�����"xU�i����f�I!�9��yW������q<|:%f�T����K]0�5����ۋ�q�1� �x(����>��^�疎,�^���Yn:��rm��X�^Mˇz�����Bo.�	϶�*�X�\�w��G�[�Hy݈��ہʶ�7ˇ���¤۵-��罱Ǌ|�>�D��Hqy.;y;sM[2�89	�n��U:�K}��ԳA
Gvb���鸜��k��\{i�b��WJ�x�����=N�����&ފ�m�?��sh���i�L�YXZ�'sNŻ{�T�u����TXofKl@�t��Qfޡk&A÷
YJLNdeH����k&\�s���F�Rm\*)8Y�d�T��c�[�JM��Q'iv���'S�!�׀o�{Tg������p��v��"V�C��wX��I��)M�:�������{���S�b�ڕ����o�!��J��Tc��9Kh��1bs�� ���C���;�^#=����J5z�SG�Tx�/�xkx7����}fe��s���<��`7�sy9�����$��w�)uw�B߼��R�&�Y��K��CR��	.nr��#z��;5��:�NV��4�bʃA�Wuar�I]7�E����ge��R�A1Q��/��&����LOvz��v�į�hH���Ҩ�u�q�i����Rz�59xu�ٝ������<�]_}�]P�l��E�ր�.z�� ��̍fK���3޿x�����̈́�MT��OPn߲�*��!���P��CZ�_�J�٤�
Z���@p�i[y�m�#���d��/Fe!�7+f�G`�+c�^��&�s;T4�Ֆ��b���r�a@k��:+�2��l�w�M�a���nX�͕�&O\}^�[6�;�>�=Ք�<��wGF���n�=�/���-�;n���R��H���<��5I��&�o!�[�8�gi�z®�SY[��:s����y�)T"��N�ǒ�������q]kU�5=�����5�.M3-pr��u�~t��U�Z�7j�f�	��.ȧ�0ŗ�J�ܽkB��A�vՇ*M��Y����i(��ݎ:�Ұ�u��==�.?br]�}�W��.�����A�J~���=�gB޸���f._<W5�.�܏��{�K�)��A�{����hJ%���~�ܝ��r�W}{���x����z�����]�~�D`�G�G��e�_Oұ�_Wr�������G�����}� �����G��仂��|�w��r�愡�_ǝy�^K�X�u+�����d�����v�>���D����8���K�=����nz��>�ït��Լ������w��R>A���r]�@��z�p�9���_e���{���^�=��y��ؾ���$��3��3��w�G��z������xC�����R�h��i}���
����A����:��{<ގK���������[�K�߼�����?p�k��/C[�1�834Q�qHT�Pcm�C�1S��r��.�ќzld�a�˻��ح��Ɵ)�V���0�)Ԧ��3��`F�^�F��]���!W�rIpwۢuj��ҡ���il{��x����R`M=�߀T�h��k瑱[%=�:2�I�W_m��_�N��yt�_#��=���u�w+�d�:��<����5.����/�n^FN��w ����:��{7��K��~���
��n�����c��}=����"���W˭u��z��{�����sѬ��/#�X�G�2?u��)]{ՠ伂���49���t��@�I��a;�����{��/>K>���yG�T��H�oF�|����i~���k�.I��0<���n��5.�����G_�7#�~>�A�y!���\�^sz�|���s�{�����#����K�o_B�O�ޞI��~��X�w��δ���3�.C�'n`y9.�񘇰r]�FJ������t_�{���ι��_q2;���{�A�~���ߺ 7/=��ئK�?so!ܿ��9�>�r���H�~���i2W����\��|�A� z'9�ߎ�qwrvO|���}�������r��:1^��u'ѩ^_kr��S���_��xy�����������]��r�=C��h�������#�P�1����]K�89��A��
O����;��`�C�����b���w��^^�o0;���_�i�����rܽ���}f=��{G�����Ղ������%�p]G��7ނ���u��(o��w.@}��~4b;����zNY��ߚMɗ��N�oG%}�|�>��h�yp�����o�7��ye�n({�C�9��Ծ�=��=����)]���Z\�����%�2_ΰw�~��_���~|�{d<�pv��z B=c�ξ��4�����[����G�'����ɹ]�oG�w��%��
}w�)�=�����+�zwޗ#!u�nL���b�_e��:b׮������h3�����X?W���<x`̾訫�J���)�c�x��t)w�Qe,�2v��t��;U<p�E
�c�WfW�Hw�!�u�EEW���Z�X�)�76]��}	!��I�z_�A���q����u�#�5��mZ:8�`���Y�[/�+���ֹ;Z�g�!�`���>� �zǢ��\���?ގI�GF���w	Ӿi(7/�S��Д>C�}i��z��.w������p�˛����Y��ߧw>[��Ϫ�w�zǣ�(G����{�G}���^��>?}�=����}�J�d��ގAJ������Bu�i���d���Д>��δ���gy�}�2�Z�����_���.]��{-'W��'��]�R~��N����ù<:�Hy=K���h_ �{�������r]�Jto��ܾ�I���\�)�m}'7�����u�}"#���C�^��/^w�˸}���X�w��=kr>�#��:�r?����u/!�?�����^h^��w���|����~}������C2r���-�ū��`�=��>S�n_oa�x���/����$:|���K���#��z��X�W����'$܏���'�w��i}���޸:�b��Q��x�(j�{��G�G�5�OP����n]����7/%��>sHy#�αr^�;;���I�:5�y?��tk�����/���π�`L����n�V�""Dy�"#���d?K�d��t��ގOR<��K���|��9'���4����]ir^H}���φ�O'��ED���߾�k'�����CpP��2��d���hrNK��ߘ&@r~�}��N�ގK��}�ßZW��w�r;�u֗$�S�6onlK�_E���r�T�_D1{�#�<Dx�K��5�9=�7�~��&��d���C�r^^A��t�K�:�<�Ծ�z��{�~د/a���{��9b�����$�7~��y��O�G�G�~�>�!����=��w#�;�?`}?�~�>�����`w.����Jd��ח��_��}��~�����6on^o��V0�ʔ�rw���Ա	,�bR4"7MY�ӝ�qaB@�ߝf�MA�O<8����"���'���D"v��fߩ(&���u8ۗ��Sw��W�,�Hn�R	s��d<���
�L-B���C�� �©ߛ������߿ ~���:���<����zL��?o�� �u�?A��
ً�;��ѣ���>��;��������`w�;����{���\޽�v�Us]��y���s�{�B=�'�#��W:�~���o�4��������K��{������F#����"}�1���u�F���[y���R�}�{�w+����K��y���=���4�����u������.��������9/ђ���=y
9k��d[��ެ������u���u>�s1I��4%{/P}�?J��9�GP�W}���ܞ�w�h)?C��o��{/\�AL{��;��#���o��&�>�_[�l��߹�9/�b���.���~�~��{ރ��y/ ��hJܽI�{�?+��~���NJ����
��IA�|����	C俺�s����:��������ٝu�y���P���99#�ش������=�����%ܧ���wy/r����%�N��\���?oO&������pP�y�7�o5�w�f�oy��������?y��q(:���8�zR��}���w�X��+�}���w#��&�{����.�:���&���!�~��}�rG�2�w��:͜���Y����s����W[�/�� ����8{�A>ޞ�ܾ�I��4%'��<�^J�^�����#�����z��X����tw��;��wޏ#�y&�����w��/��ܩ���Y�{���_{�=#�" �)Ƚ���oz9#������Jt��=ù}���@{/���z�W����K켎�`?^K�tk��9���_���
j��3:>Yǹ}�#Ї��s�b,{ۂ�^`��<����@�$ް�~��|7�<�s��|��y/װ������ٿ4�/���,�������[_��_�21J�a����՜��>�����=I��4m�I�3�%�5��C�mu'{t�"���7��ʻ��͇�%�l��U�8�\���ʡ�'Sl:����ِ��@s�qV� �2z&+���[�t�����~�v�g�-b%�o�{��>�|�]n���#��ˬ��r?b}4����}/ ����7/##��;��u���u#�;ϴ�]���o�7/%��>u�w����G}������Z�|��ϣ�{���Ӓ��pu�S��/�ֱ܏�d~��P���A�y	�����d}�4������Ҽ��7������Ά'�R�HP5�ܖR��Z���_��Z]����9�����d�����bI��Y+��I�)���I�w9!ѿt�%���Jd����⏄�O+���N��Ė8�C������|���Y��zy֓%}���irOa?&by.��f	��sֳR?C�Ԝ�J�y��&��䇟<��O������oZ�!y�{�}����������y/R������پk$wK�:��/����.M#��>�%�������F+�����T��������ػuoN �����T�%ߘ�|փ�y/אxo��r=w�[��K�;��y/ru��H�KѾ�9#�?�ir
O�}K�#޶놉w���KJ��#�=�����$�����Ԯ�~i7/=�;�nW��;7�GR�#��r�=C��;��:��:��w�9'P�s�+�0��%��=�OmV��!5v�~���#�{��r�!�k ����:?b;����Y+���4�{/ ���w�rw��:���칧�������_ �}��{^��~z�۞��]S���������Z\��׹�9Ӓ�`�_e����#�c��i��^K�<���/Pu�w#��:�4w!w~�:���nMm�m��_]�>Ϣǽ��G�����<>ށ��ΰԯ$�}�r2G�����!۬��_��؜�r�-��#�=�=��G|=���CZ��W���#��^u�b�����q幀Րn�U�縪n��G��Xn�u��0�k%*��}�� ��}��9kd�$��Z���69�vP���GYRXR�&�C�Q��V�c��!�ڗ�[�1%�\
�-��������|F���=�YK��|�m~H��D����<�r?���GR�
C��IA�|����hJ%�o��w'G��r�W}{���x��X���:>��]�9o�_Ձ��_Og.ߢ�B<�<�zC��]���k�>ɐt������xr]�H{�h;�p�9o�Д>���?+�z��.]�ﯴ�w�����"Թ��W;�[�Є{�({�3rnG�}��z��9�{�<�����^��oAH�<ގK������w��v��_e����/ ;����:߻>�٬�[�z,H��{�Gޒ�v��:�'�>G��������z�s@k�_`伂���������u+��y��q�=�\��{��b�m�
Ol_���}*���=��ϽnK�^`�d?��:�)��^��c�_#'��!�����~�pR��/�n^FN�����3x�?J�5n>���O�յ�˼z���=��0���ι�䯗N���H~}���C����~��Ѭw#�����J���A�y/_y��w�#�7�W�u�ig��\m�_D{D{G��U'��~����r?<�F�|��]b���u��=������M�ֱO#������}����pR?F���u��L�9���#����Wꭿ��YU	��������2^I��z9}�;���[��y���{/��K���u��}������hi`从{���l����ۛ�����DP�����������2C�~�<���ßiL��~:揯a信�1��Ի�֑��/?bd����ira<�}�_s^��;��L�J3w��P��/�DA���= z"�u/��F+�?G�>�ҿ]}�A�wy)���]���>9����[׷��/�{7ހ�{���|л�����ב��0���<�\�Q�s3��8w�W��@���Y�jٵ�LK��F>�Wp��*z�
7�S�I�p�v�wj���޻��@k�![��4R��|ˋAS^s�:�d��}7j#vqἒu�4��צ�Et�DɚF�5�ai�VjF��S���z=�Uۚ�ĳ��B:��`���?A��
Jp���F�<��X�f+���ރ�y{)ٽh<�����%�G��/��OG�s�Q+���������p��{������/#�z��+�?o�A@���9/#%��>�p�=1��~��',�����I�2�^I���䯶�\;f2u�)����_Smb����X���{�[���C�����/�O��@�e��z
Wpo�.FH���%�2_ΰw�~��G�Gr�����]��d���x�Q&�IBW�������>�r9?I�sGrrW}�4~�p��o�J��=������~��=�K����7&K��K�}��cf���S���k��'�E�}�S�{%�����M��+��~��rNH�7�C�(Ow�%��
z~愡���P������x��:�Ϯ���^m�Ϲ2�Nr�<����$��=��u�'��S�}���^��>}�=������+��~|ގAJ�����;���|��;���;>愡�3Ӝ�� R�����ڵ�G��{�,�x��h�V���~��brW�����w)�xy��w'�{�<����f�оA�:�z9+���z9.�%3�{_fk_��]
y����rK���#���s"#�z}����^����w��2G��O��7#��:��7#�x{��<������^Ao����I���u�s]��{�~���w������^���ܼ����������K����C�0|�_��2Gې��5��|���brM��݉�w��:������~޻��>����������ގOP��������G��hܼ�w��u�!䏗\�K�����%�&��X���^GZ�r�FG��g���Ѯ��[�aWF�X���G�c+�
����th>S��h̋�V��R�9�Nuy���խ[�(e�}Ւ��V��[ht��v)[Rڲ�<X�w��t�7����l�{	\0b��um&��0OvM=�j�qP��49-oBD��$���""���RiŚ���	r��Ye�Xwk{)%t�^M��M�V՚���w�I������q�d��������h�:��3���B�c뫅geX:���s�t�9�kqQ�4�Q}��̩41�@�\t���-.�ԩ�Qyg�awU����QuīyJ0_
��
^>������g�3�\R����q���7M�zC[;53����D�pr�ޒ�JY*���Opv�k�|�e:�F��XsF����0t��Mmm���������+#��d����T�T�yS��e�/�e#��ŝ�Ԫ%�
	�8���T*���x�=����#X.T��Ӗ�n�d��Wz41[H7��4rҏr���$G��S7�E���U�;�E�N��x�̢6��b�r����˻i]!j��8�"�bGC�l��:k��x��qA�`p� sJ���:.nJ��TF�0]%��[ڒ+ݮ�{/�ُLm"�NF��UX��T�t̬w��s^�+�I�Ҍ�yOSXy�g7L-�AmpBWa�R�����i�̲��W�`�7�!	W^�����R�W�L���82£�/�U��{�\�/E���n�G�p͹�̧�F�"��ב]�Q������1쇄������EFv�=d�ؼ�%�IoWi��\x��`\"����y�]�t��"-�)�X��a���l�`�?�d��b����&}#�mm�r�*��.��U�)��.�ﲱ�#�����<�d���eE�Y�j�en��̢�����fM�_+�����_]�5�kxحu7�C����x�b9�kp�C��im���P�l��F�.;�c��R��'.����F�R�B���{R�9x�]xq�g_GOs#�SD���u�����Ff��`TZkm<�K�Ӛz���I�;����l�q�B�*�R��"�n�]���eRnȪ/C"�ӌ��h���.j7�tr`
Cg�s�H�x��ݤx���D�wq�:�&O�i�¸�"��ޭE��Э�s oyN�l�g#�x�M�4����Y�n�Y*:1Ɉ$6�Yذ�6��p�qvfҌ�K��R��Ok�ǹ\\={g��w�-h�+��|������ٙ0�9�h���b�-��p)��!8�8e��Tp�h�P���<	��o/�&���.��ݱ��_3�pr�i��rʹ{�T��-��R�G!����4]ֳ��m΢�q����c��⬯���R���M
��ԍ�m�p��A����ZC��L��a+˘�-��Im��J�W�Tg-i�����?}��4��2(2)�)��jl�ɉ*���,�bh((�H��)����f(��� �����j�
��)����������ʚh�b��"b&a�&*)��)h�!�H�rrf�**��������*B��&���
Z��(����f��Ȉ*�d*�� j�)"�����(2�&����"*�)���&��"�S(�(*f ���c �&�r����
�)hr\��&�(�� �j!��bX��& ����)��b����*&�J�������"hib�b������(�j��
�����(�*)�c0�)`�j��h2Ȫ
J
J��
�Ɉ������ �h�)�*�h��#��5-���{�	)oGϸ^�%�]κ�𾮩u�g�N�=Hl!e舧�ޑ솆2q]m��y�8b姳��ʨ��~��=��o�s���S ���u�n��:ߚL��y=;�@�A�kz9=H�N��G%��n���rOm��^iw+埱r^Hw�����s�?���-�e<J�E�?z({��b>�#����`n
O�k �^FHt}�$ܻ����d ��i�د$�7����e��+��;���ӣ�}�Y{4�W�1x�����R[��G��� Dp�/��<�	���tkB��Pr5+���7.�$7�t9'%����Jd�����qK��z��{�|���$"�].���--�����}�s#��F���{)٘nL��RP���ykH��������NK�1M�r�^]��>ҙ�����=��{�g�WK��y���c���P���e_�:��l�Sn��B��t����z�M�梁�b�Z��x�%��T'��ݷt�a\)�B�bO.�0�Ѭ�����̪Mc��D'�Ր��5�a:ۄ�m\;t�* ơ�V�ĆKp�R����{ӳ.%�y��vF�v�w�4�������M�;��3�/9c���i*T�@qC��[�.�n���s�U���&Շ**!8Y��	i6�+{U�󯸮v��(��s(�
佼������v:�`<N �|�3p�c���U��h�|o���懵��N�Գ�E��a���f��-٬ζ���	w[xVs��ļ�/q���5�+�ki��u+C��@{3�\�p���\� �[+A�yl����6.�w:����)A�_�ܑ��vj��^E~ǣ�����$�r�˸����(���S'*#�U�6�>�\�z
�%��EP�5�u���
SE��Uz���+�K~<}�X�Lꬃ�C��}�vgY�[��Tk��s�(V�u�ebhU�[���^���d҃�&�\r[:�'��n�N�B���M���&�[o�U�l,p�9}��qy�4�x�d�c�3=W�v��{�=�;��B*zz%x�ᥧ�/'(�iw��+J��b)A����	|�)|�M]��3�OP��3Q�h~����*�#C��'Yq��H-ݜ�54ի�ѵg����2?\M�Ͻֶ�m�!E�kU�s�(�U+^Md���k����r�[�\ý�N���0���م"�Q>�Vی3E��7��7W1����ӫ/��ٛ:h]5R���˪��*D/D^�1-��ɰL��$�F�Ict^�D��Z���\v��	Xi"1B�ud�uX�O�&<T�;�oq��>��yr�n5��a	l�ٰ:���<&r��~�t�:`Ay>��h�E���"v������彷�"׽%p�(����2��9�!�nY�=��oޏDz"#�v>n5��F�.��ݷ1���uD��;��˞9�榌� ����O�n��X�[��n=;�>��L���n��b�k^��F�S-�^�j_�i�R�sߩuM���j���<�j�q.��X��+��.k�VTޮWx�K��(Y��E�.����";վ��!U����ڏ?jP�����~��O�ksIҊ��`����>����'�Uɑ3M��{�.�d\�}��)9���[��_����<}�X����Gd�<Je{'L.q�b� �:�zP�Ϻ��=-��UO�|L��[]Ѵ��B���H0��ע�Md��M�Q~��Q��^&���Dv�k���L�������5�w�,5�%�uE`�nc�J�������ro416��t+�]jմ��i�/SyF�Nh\�6��hO���C�
���U/�U��`o?M�cpFl�Ύ�_*,�X��_�NPk���u����Z�/�u��p��^����]s��v�:�Z�	�rk舤2�7��H���A�@pkǸ۵Q� [[�����(���ε��`!D�rV�R9�3���6����諭�DF$�MC�]�u��ߔ�vyoVu��#TrU��m����&E���oi��B%�Bb��9�O���v>��K����]�ʩ3��Z�z�t������!Kq�|�}�n�w��uD:��;;
�ر^rw�RZ5�c�G5F9O��z����G�}��*A؎��8y�_,�߯�qM}��u	^}�zl�D�=�N�4�k�Z��4H��56�������ի�W
|�A��Ğ\!nF�
�bʷ,��ݷVr�"x?<�[3�S�(@�[i�ؿ:{N�)�S�+JZ����:�'�e{����[�|]>�[�nڿx9[i��Roiܺ�`C�5"�����N�:v������x�u��u�)6S���dTs��*��#kD����F��꾂*�X���%�d�퓀�bp&95	���S����Z[7O��ފ�����ܢ3
�0u�ᖑ�Uzl�\�=y����B=t"�'=0�"�"�W|��v���dո6ȭ-��ڗ"�$�A����؍$:�b�D���c]$�i���i����X��L��-��{WAD/����]�/�_W��}mB�9�"2R����Q=ԨՐ�Sw��EnR����58
r	X�YQ2���C^$�:��m0|����`=g_Z������X�w�k��r�}��3x�SG�\ArX�x�^��S�%W����M4��{�so9^>�nsWp=J��)��$��cMnE<�v.b�J_2���18K�)g(}��	��PJ;ag7:v9�M<龵���́��@[S�r�knͤ��ҙ-ץA��LW`H,y�w�����;!,�lM�=ջ�,��}��й5PzX�%�WJB�ho/�C��OL�`�P�j�*x�^��WͰ��Pم#f{����J��4��d���Z����j�t;��q�x��ֺ��5T�j"7��&�c�qI�d�u|�a�D�O��V�Ng7&���n��ܭ}�]�[~���<�m.��{S�w;�	ܼ8~�ϳ��Y{pN;���2�w�A��(ةO/��i���-�[5�xuOQ�n������UVĺ�ǻ�}-��ŕ��T���ȹ1ӌȟ2%�d��l]e�.,JZaTNʕ��f��Dz#�ꦵ6���o���x�~�r�37��M�WC�N�d*�`�%�vv��o&��֪��5�>��;#j�y;�jÕ��NEy7������ jK�h�*�>�����z��%m�7��Tn�&m\@r��4�Sa��1�C�V����o������r F�Ǣmx
��v�~��G,�,o����Aj�������U�2�O���Ŋ��H
Z�S�ū79���T����-<|��ud��#��L�
�p��W������\�r}����=G�����5<�|��|M�o�x�U4�oC�\���9{Ѱ���s[���J]]�Ш��nR�މ)Da�
*ǩ�lI0�y���g[#=Nm��S9�)Ҹ�N�꨸T+Ǘ�0��{�,�u��%����P}��!�X�\�f6���<�@/�9kK+_�����7$�I9���к��t��^o�w�
�j�G`�tFv�p����C�ϳ%���n�,\�A��������4�V�T��5}A,�p^8s�Y@�0*m]�ϡT�6j�;b���\Z�!�W>�������^{�}!�[p�����W���=*��Q.;�!5as��n��$�w:Fe���������j+�~�
Fφ�k �Uױݩ�r^U�҉��7Զ;�3��^w��������1��
?f���Kmف-j�r��Z�_%")N�})e���!sUo�˦���.�{HJ�h,Ӽ�6}���w7�C�a ���"���,OnW֦�y��˭�K/����ۓ�o�nͷ,kt �P�><�jV�0��o>~sMS|<�Mz����]�ޏ�
����^��j[����-D/CN;Ս�_I�*׹jD�	�\$޺-P�7LnDw�}=����#ͷ:'u�$�z���ޭ�/l�6�lEbr�>�^�R��i������k}9m �gdo����^��]�����-���d�����uk�9۶����tu��W���=zg8+@��sVĸ+5�Og��CxF�ƒUjt߱ұ��߉�e�w�RBw{�w�4��^�9�7��O��7�y��'T�X ��)Z
� �@ޭ˱$ٽe���}�_�;�@�U�9��꯾��Y���#V;�uc�{hކ��~]��58ʌM
�kC�3���q���\�����QV�Y���etNkpv��u���S�6h���k���5�
�a�&�v/u�f��ڦ/e2��8k}�v����W>[�����Kq�ؽM�1�%T�Qp��1F,�[
�$�;w\���q�p�-N��vyoVu�o�A��ၪ��X���5�+Yo�����.%Fϕ�)hlS��9>v���u:]F��.�ۄ�〫��F�Ԑ�c1�A-ץOWJB�n7����>�7��]��8m�K�*պ�w�BjF���`o!��i}|/��}�Kz�l�zs.�z^W-�9���S��W��]^�=��"u�اcӉ����	��IbN��CpO(�g�=ˇ���
�:��^�8�*-C�&��\V��>���]e��k����@�r��R�ٱ��m���o�P{�l�2�,�(nV��b�;Vţ�Ԣ�)ŰM2������3J[����\X
�p�*Vi"�}�nr�ꢥ[�@y�L�^qr��_s]ڲ���`���/�s*�Ɂݝ5G��z���^n�;>�����u�u�����Ok��LB���'Ӏ������Ju^�/��k{=�u�W��m�q9��w.���ۢe����P�x�.u��&oUo���-�C���M���E'#�]nN7�09�$c��\\[ަ,S�N�����GvӾ��p&95���W�7y/ǝ�.^�9_�Җ����T�q?�t�6T�����B�d��!�>���ѿ_}�+�W ��E��d��WJc�i�j��vR�-N�P!X�zOqz_|<<���>a&�uuE`����Gm���oo�8���xOEB��S	�8I�Ɵd���\�	J���	�U1�%�|��.�d��W:�T9�`Lw�ju:w��M=YX��et�&N�O=��c��ά:��;��F�LTv�,y�vY�nb�!���Y�k"�6q]�k7n8�.�����hIoO-�Okyr�աEzǞm�÷��a���}��U�MK� q����.F�Mâc�D��7Q;���t�YŬ�6ք� �m'rn��U+��������n=M��b���v��;h��#��z"�y�'����R�#l`j�J�uW��WJB�ho.�ΜZ/��Kv4y����Y�����7�ZT:0�l��`ku���-] "���w���G	R��*l�>�SӪ!���x(���S�.H�u��_?�����-}
Z�-�t)|�*��;n��J��u�'~�N�R�C�B����ȓլ�r��㗊��g\x'[~M��÷U�p�r�q�ݛ�����]�8�$��[����ڮ�M�j�^N' XY�]�ZW��l�zӅz
:���;"��D��X�s�U�����Wcf�-�J�׉M�ɸo��r��R��Y��5�
�J���#��l�,����W `���8��w��[rR���o������1bu*#���xt�I��ߣ�O'~iF�J�s<�G�|�������X~�t��'|��W�F���;�f�wu�XU�������%�xe�նQ	�S�8ƙW5Dle�O)���-mfӢ5-�Z)ҩ}�T�6^�X+$��i81ܕ���F�n�vV�Z�5΍K��R�ˢE��ܦ�n�����~�!wڴz��p�mu*�(�Rpe�g5
�y����@�7z�LIT�5�P-Q�W}��}j,C�q�He���F�CQyZ��R!�� ��i69���[��Z�T<X��F�v&�b�����8���ӹ6󭄐�/��౮ތ�H�����J�f��%��gp8�v�9O#���˗ם�옟%��(�5��\��m5�J܉����⯻� �F���3�t�A�WY�q� ��yd�p|r�U����^
8h����TVӷ� ��u���켕�w�M�b%�'k���_p��A	X��Ԑ� �����p��5`Ņ��X��I����\��V���\�5ڧ8��r��&j�ɇIM"�G��<�ܬ�FUt��0��k������4����̩�K�!����0kTà��wf���FE�+p�hʻ�|J��ɜ�����k(�vJxR&���T�اlk�+�٣pu1:��;{���+ih}��FNY:D���C`�C
�YK�l+!��_�����2Yn�ifm�ݡ���@}B�7��=���x}�oT�2������5� �R���&��ʹ��4Wb�W���I_�d���G��+�A��`x���1c�W.��/�*NJ�x�v�7�-a��%{r��Ö�%7����p���+�'q�,��V��D�T��r�b�z�|O0e"��rS��WR��F��@:��;0�s�`�}rHa�$Q�urkR�I��*\	�6v����mN\.��a���(�y��]'b��ݳefaiVQ�	�s���m�۫)q��@Gb��f��a�nK��@h>�2�寂Kx^=�+`(��.̨��:�1�f�B�>W��_;��7P��[�ډLg�Q��=�\��T�pQ�k4�D��D�U��2���H��7�d8�I�n�!��X�z�J�[��%J�{	��ӑ�^L�F�ް�n�i�m'�#:��]3;o&�#�jx�܍]*%N�GH)h�Z�?&���_[�X��WbWw�Ems OcnC5�H��9�'�r��y-���<nY�e���gv��D]�㦭�V�VOl�#�a�ކ�
��s�*T�\�捼��\|]���6�!H)�eui�D)��P�N.�F��oac�%#N��3�o(�ˎ�_(��t�e=T���I�����&.[�V-=��<N��g\�����/P��ڹ���ꉁ��Zs+-6h=�F3W;����Q< |�-0c�.��w���6�<AУ���:]ؓ;�۽ꏥ�&�p�k��g�Ob1�x�#�Rn���E��i�0�����M3L��EFfLAD�D�6Y5ERPTT�DD�S4���EA-%P�MTIQ4SL�4���-�2R�FXAM4�	NfQQVFS�EQIEKQU�4CQ3�5D�5R�U4LVY	EQD�MQQL�I@T�1SԔ�UQ�E1RPP1EQSAC3E4L�M1a�SAL��f4MEUUIM40E�a,TD�PS1FF-4P�e�T�0�	U2�TM.ELTP��5P�IT-Y�TX�!T�QD��a��&I�AACQE��d�FfUHRTQR�T44US�EU&CYYd���MADY%4�MQA1TIY�RT�ATE2Ĕ�(�� {�47c�����%,�M��Eb��5g�eS
,�@��W�F h+zI};z�kA�fɠ��o�o�U�UW��E��c�bL��� ����Ջ����=/�xD�����ZwJ�B�?d�Ș�˶�����:�w�V>�ν����o�wt{���^�\#s��d������_w��Jm���SS�)�:�h�Ʋz�F-�}ux�M󆹭�łC�-A|'Ԡ�h&+�$2Ct!T�;F�噧��ˇ���r�46F���qÃ�!�R�5�J�źxW�~Z'��om����F���|5��.�";�����5s7V�~�*��b��{���{ΝoWBauy�م";0%7y��������k����Χ��T9�3gj�S�r��\�u��}�����i������{�.��1[�W��B��1Sx�'�������Q�Z�%�ە����C�OP3�mw�D4��G�)��ͭ;Z$��f3B:T���E��#��#��W1&�շ <��́Q*��!V���$�߻)����Y��������wN[�AJ{ �uޜ!��^��%&�0�M�ǌ�u��$cqձZ�fh�Vv�x-�$>��;��n��~�������O%ͮUYV|����Oi�5 j�d^�ض���jʗϗ�~�q1:g9pݵ~TTBp�)7��]+�G\����b�al�v�n��K�u�y�گ���Z��t������d��Q�-t�-�`�g�{W�%7�,.Qvu��� ��#�BN~�������Z����M�oW��Z�NX����}��$t� ���zP�ϻ�=D�K���5��f�A����ڝ��6�÷���Ņ�+/�!����ZW�B�Y46zux��|Ǫ�����y��t+�Xz��������GX�z�*U8���;���W�wSN5���T�	[�U�Ep&��h��5�1C3r�]8�v!3B�X9�Z�B���o-��5�M�l��!e�]����7����}���Zahls��9>w>]��gS��P��\QV�fz���/�������-𦂮��*�#E�:�2������J���]��]u3����K�KN�\4�|��ܐ=C7m"��7��*����])D;��9�|��/�p<�b*��B�L�B0�#KZ6�(AW������y$�L��oÇD�jTN��s�Ґ������sO����WW��������J'x}�>���H���)�����#�����E7t���՛|�^MʮUM�U�9�"7���˫�c��=|�Q�EuT�Ǌ]���UMK���ׇ�p�}:��u��A�<�Bڼ�ə闄�i�,]0�N;�J�z��k:�u����t��% o�gg&X0
]���z��L�����U.A�v��r��8���oj!ܼZ��W�F�����]�u��g���a۬����F�a&�Bt����D��:������_j�kt>u�1yu�¹.������ݒ�X#��\�����Z'�>�^�uD!������b��@���: }��=*E/Ͼ�eX��>j�)A���Ua�jxEa�����
 V_��W�}����d�"���6��*��|�����l=��%�H����aqǁ�yl�+N�����D��B�j��:�-n��>�78�B�s[Zk�k�r�K�Q��|�M�N�(aj�ݰ+�]�N�PG��k���p�y����hjV�����r>��Ǳ�7��z�X����&�[���ou�W����I漬�5hT���.�]���jĨ��n.'S�)��$��O�S̯;hL�稓�e�5�]�e3���	��>�G`Lr��
t�Ú˄�������WF���ӝ���Jι�e��ó�1n:4�B۾�nk�콷�ݩ�<=�F)�9,/T�*�������WJB�7a�lJ��}u&z��F�&�w�&W���[��[n�mZ���:�ӛ����?M�-�L*�*j�<�	��U�kf�g�ܭ����^���*�\k�Y��%�-J�Q��\#�9���\ߝ�up歹*oH���Qws:��Z��˷Q����X���Wf��U�^޶��ݠ8{������+-@����������rV��
��6�ݼ�2�+v�rm��,,�orfQɨ�VT����ݎ Gn��횪VC��ԥWyǺ-��*�iO��ַ�3�nrZ����Icͺ̅�&�e�E����+�����e�ܻE7.k�x̻פ�Dɷ��Z��Ze�� �5ߒ��iμt����ۥTB�=���ޏG��sK�>�k��>���\9T�C��V��F6��?T��/]����އ�D5憅 ��﫜�k���N����W��D�}6�Hzn*{Ҟ�S��_(�.�4D�Iv���<���p�W��LB�ub�{c-ץ^=�,&�(nN�B^w;��v����OU螗�<"�OԎ�,C�r&�۹�0�Se�9ʲFV�E�Ϯ��ޥi���bhT[����X�nn�(��\��3���ǲ�
�1MO���\D�y�B�Wi4:&P��i���{�1�I!��Х�D��ϴ�C{]+)u�WS*zƩ�]�����jE[� ��OO�V,�4�p�Pr]�iA����z/V�ғ����AXz�R���o/�E�B�U��Q�U�]����n5���b���w�ho-�sI����>�:>R6``^o����,��@պ�=�Jom�4-v��P�1�e��P�i�R}����6�c61���$��JC��~�ʻ��k[���R�P����W!KS�[5T�Y��=0�Z��w�M���/�BB{�6{S7�-Y�`�Bmcۍm�qI��<�Dr�����s�\Sx�z�)��.]Dt�)n'��9��W����O��ZMxSi��9�$]'j�o��"m��+�7�b�gm��j�9w+���lN��v�ikt��:Շ="�^㏲���O'}���noݼ�'%�1�o�ݎ�,�X���[�5u��ו:�ϧ=+f7U��	YL���d��'��b;zg��R��u�n��1^ڝw�)n��/olK�k�G* �65�t֤�*Cvz���v���(�K��S!��X$�G�e1+ƘW�xs�o˹�E���MW�YE��6s!'pI����M'v�\'!)�5��*��}�jb��S�g���*�nY���
��!9�O8;���|'۾zL���c�P4�Ժ�� ��>�3����ov��ܩ�Gi	����8Ii��ٸ�uGE�:��,WV�qƹI\{��8�QMw^��xi�O�c��tg�ͱ]a�z��ЇgG�p�z��"M��ݲ����G��3֊9:�JfD�QM��:�un��7�c��ଡ଼��-X$��5��CWC��@��2�	�}W�Blj��ot�\',݂ν�.�"T�K���'S�c�9�fK�l;��p�޶�}c�#c�n��Sװh_�����S�>xz^�=c��U��\�,|}��hB�ڵ��ږ��Kΰ���+�=����w�ڶ����w�8�0�Fv�}���[��g�p�\�A�P(hLt���}L2����kq���lG�O4P���4z�$���W�4����:zcQ�ފ��
��h����$E@�z�N-K����Lߦe�t�^YLQd���=��'���˄�qr�z�\�2���j�u��J�t�9�@D�vx;�<��PJe�G>ڇ��!�z�v1@2����K�;�6�(�<ij��T�|O�T���LOeICaS���1{{�{��!���nInC:�����Q�9Q�X�<(zxp�f��P���n�z�^0��n�Lt�ɧ�LXv���95��b:�7�򐻇�ā>�$0#�����)��k�v�HI341v{����_�a��o!7 ��,�s�2��:�4+��v$��%�U��ҊT�Q8K��&�F����l%��x Y�7��C����QȸN���qE�8o��2�{�MO��EJ]�!P�7p�/z�r�k�ܜ�K�VL�S{����Ǜc{sn�@hnW��������T�9�q|B���-�z�\urj���2:��,E��ѱ˱�ɦ ��>��FCyZɄ���hb���F?�}��U�=�}�É��fh}�$��$<%�$��he���3c��'�e��������cn��^E�����ݿ�H�g�F�:��f�	����Kʥ��^
E.�ӂ���D���+�.%�&�⹬|��/Uo�z� &����u�[lٮ�J���	�����1�ZFyJY^�h���l�ū��C�1�V�p��Ց��w��N�c�	v-��f�p�~��e�Z�OF��sh��R�����ϭ��6����J�yLwlJ8Tqт��&�ǚ�]͎��2��Ms�ޚ�n&PDթB�
���xC��ڄ�ħw�XZP���l-s��:��՚�-c�:��n����k�V�`.��`^���`
[(;��W��OfeZ��i2��#��29Dd��gR����t���2J�3��EJ��
d��Z%�n��3r�@�Wl��f$��8
S�ᯂ�2���(Κ
��G�Ԋ��UN�(�VY,s�Sw˂���r�����F�*!��Ë��mܑ���PP� �	���K*�z�a�=�n{' ��u�ed�3�03�:c�;���%�١��׎�2��F�&����v����OV��
�+}5��+/{S�Ɓ칰q/9R�\F]�C,K�Z/2F�gI��TGD���ao�����a�ZW+�K*�p7�������~n%��K
��S�"�xr_��t�}�)	]�Ժ�>}�dh~a �yE_7�d�j:o���OO+�#��0m�DK��s�z^���Czm�0��Q����κ\)_�8V���4:�w��hMV��`8�%Q(6L#k��P�l�2�"��օ��Zm9vb������4�}5���	%��K��0�I&V�ĵ�Ü��{���[l�V�˚���2��:�E�]-Y���]=륁2���+�KN�a�+�Lj����ꘘ��g9
�YS/轢�n4�{^�#�68s
i/�ĭ 0�)�W��	�Q�/D��6e��^�����̸���z��t~Mb� ���P+�ĭ&����*!�#l:�eu�B���Q���M�R�u<���~��c՜n�5�'���'l�(!�c����oi�Ċ��׷`͜sph�]~�.�j��Q��P�t�.�������N�7�q�������i���2�O|`
M�o���ņ���m�K��sσ�0�";x=�-�����b���e���93��x�����aW��kU�_�5u��%���l�]�4��ٖ&\�[�ec9Z\4��A.����I�M��=�lǷK*Ԯf��}|��a�͕�Q�Nڀ��iP�M_=q�9��Hv�zՌ�[WV����ѸM��|>�^�Ԟ�c�Հ��U�~�;ǞIþӤ�7'DPB0̨�%��iL��PSɩ���%A��\�F��J�vD0�Ŧ���{,j��0T$&����`3ra@�q��o�4����Zc�\.��){.��
��c
u-�j낸��8T�%Iu���+�H1*��Z��
�v-����?)A^[%����b��,_����a���4R�<!Џ>��|�{�ҍYi"t��f�3<�L��꤁�czq��k�9[��7��b���ܺ(��|��u����d�iI(�����UAڪ���]��[�x(Y�V!ˮ�P�:�ў��m�e��G!ϕQ�>�ĲO�Ġ����]ឃ�mz�?L�5%w+|����%��z-�� ��{�X���`@���5�<�T���L�2h�����s����V4ÍN��5L%�3�b���tƻ�� F"t������`�LD�G���ہ	�g��o��;��ͳ :��8�6/�a���"=�U{���m��ɃY��㻕7kϊN�u�TD��Ғ�7.[>����y@V����'w-��iRl�v_@�-U���3-Z�������Ǳ�DJ�{">�xY] �`��r�Mꠍ�ʀ�Mhw�^>0c9t�f�qEe֤qWX:���FjT��ꫠ�c#m=�%%E@«�)�"���cʲ�XE�V\���uX�����wNW��e9o@KyM$��6���u3n���A�K.D�.�P�F�+�]���u���]h�;�*Ⱦ����u�yzJjl6.F#����'��Edj��?cX����$IqV_�=8�WA�!�o�W��n�a�����ܖ��"]
Dc|�3hs��uqֹ��)�p��Mr�7�qv�����'$�G+y1��u�qx�L��Є�3 &���Rx�3�u!»k!71�;G������4]�Ҏ'���;�I6�MIM�/E�9�m;��eD��m��=�컒���k��$��L͓r�=�Q�b����nu83sSXQ��q���8)����ehɐ����f�x&�ŘDe٭��V.���➣\p�=�t�7�]��_����5�e�p�m.twHgj�hk��R���D���#/�kF)�$+�Zp����^���V�SBź:�m[zRI��ŉ��Y������2��u�0�7�ōn�Mt\w
��{N��"|J¶�q�Ott�kFq捊�1+^�Wk���P ��֋��k-�f֭ύ�MF�諴zPmB;�b��ҧ#���0[9�O5]u
)d��s�u�c1�3��Q�dv/\�ɳ�9��`�[i�Em���AW�i��圝��<���H��9EN���wq˧6���X=@$��/���-�GZw*i��зh�Q��l��J](���X5��+o�&gKa��`TمE�"��K;��B�N���E
K"�GU��ԁ�YS1�%kW���Z��EecT��������y�,�8�L8�Mb{^�oPn��q�&�A��;5���vFeӦj��:qŧ����0��aئ1��JoQvM�ͮ����-�MO�Ä���GZ�k+�(%X�0m���zn�м�q\M����k�;˺�{Rj�����#��V;̜��FKU�d��m;�*�WM$r���9�����Tk������u8����r���r&����ώ�g�4
�V�+y�E6s�mwu��oF^V�]5�Z\�g3u�Ѱ|_bq�X��#,H�n�7;&+��g�m�/�do+^.�ѫ$wv�+T�eMs��&N{jHBg���]�%�%9Jq�5�Y'X�Q�]���V�t�#z��j�t|
�i�R*�B��U�T�h�r�U��B��̻�Z��7)�#oM@�.���9k%  ��jLKb���3���z��p����x������ιTc��-�d�Zld���w�_�XMUDRY�I�TMU5BE54U4�A1��Vcf4TT�T�EAM$�QPDD�4�DT�UEE�d1FYL�Q�a1FAfEE��1�&Q�UU3S0�ADEQUĳ5TنP�a�KSLa��Q35E1HSP�Y�SE���Q-f�QULMEfbUfEY�D�PISIKEQR�D4EQAU5A4�d�DQAC�M$�QC1UUE���SRDIQE��T�ETRD5EL�TTU1Q,2AEDPQQ$TP�FQ5D��SAEL1ADfa5UQQ)TD��D��DYԑU	SQADQIS��51�ET�%k�l��� �e�QX�����2(��A�
��%��n=Bv�+5�̡���T/�N�����).@.�IC?"=����M��9�٧�$صSq],P�ٰ�;��ĝA%>�"S�P#�	�va�t��NM鷺UT�|ح���vIè�01B�����x���=�'\&o
�<6g	�%+B���*�:�mkK���k�{L\,���UxhxӲ�����7�/�:,z��;�n�y��uVV�V��� U����8�N�k�tg����u����p�fU�k�h˳R�r���d��Pf��N!Z�(`��Ց��n�)����F��d"u�R�4�N�*+q����Z�pyǵ�xUtF7�7��A�J�gs+
Ʃ���:c�؛��4��^�s�#�.�Ջ��tӉ�5}`Á��QF�W�*_S:zpj1�uQ����j$IY4��,�!�W�{� ��}�fx+�@*YL^[$6��,��a�N�sa:{WǙ����J��d$X�c�f�0� iAw�L�WꂸUM�d������(ZQ9��g1Vofb�9���Lظ|'EC�1�D`I��u�q3�TEʢ��t�{�6�1�2a:�h��l��+9�r#&;�<�D�ogl���e�>�\���=�����ˆe�^�F?$��*��}�>7��vp��*����I�y�Fv��O
���B=�zs+L]�{�����!f�`�׹�,�ޏG�R�|�<]��ϡ:�����ȅ���s
��E��$h� ��ki��1�h׭ O�G�'�f\�}�i�s���5"��Y��v��yH]���v$	� 
[+7]eSJ��z$l�10ٯ<�P��<�N�V9��
�ð��:�X��"X3;o��K�-n��L��]��qrQ53�&D!��Ű�ulpA����(s1�|��9����r+� �p͉�E�o�nfm9�p�3�$��2-���3b���A2�X4�]������U�$ܚH��5~�M��Cx�o�uҫm���B�yT��k��A;J���o�^_�U�8�G0����e�m�j:a"Br����sPﲎW���]E�M3"�"*2��5���uv��iq]9g��c�T���#�=a3|�V�ׄ��u�xd��-����nQ�����G<DZ�7�W2��^V�Yq���X،N�7�)�4p�q�	����6(#�j��3����&R7~�CI�R�Bʧ��xC���G2{���^'�xe�'
bf��`4��,���vۆ��p���K5��Ձ!��ת��m��d2�4VU�[bQֽ�{\�s>T���x�-Զ\d=�
�e�`��X��-�S�M%��&U�Bx�*����w O.`��6qO+�be[��o^�]+����8st�\&~���ٷ�����J�(P�}����b��g .��;x �%~���sip�QN����z�3��c|xG9Ֆ��Ь����}��z���%2E�h��J�4\Mv;kΌ������\@R���Bu�b�jN�p���Ug�~+����R~̽�縷I�_�	�ں�j�F����Nyp���Gl:�8Q��I:!'��P8��';GF�y��d�������[�Pv���
��(\+��9���Q*	 �����xw�7e"X�J��1���U�X�8p�afӷ�<�u#��r|�(�޵�Q�I[	B�Τ���߅2oe�|�t�
�����je���~�{/!�1�㫭��1�}��U�n�=�N�ǥ��"�ܫQ��j�99��WT�Wm@r3~��2!gL�OU�!�ե�%b�wc�U1�P��*�"��&�$ƠxqS���f��`.�i�Ä�9�Y�x��q�@�R�	�D����0�D!]`Lm�]���/EwPɌS����v�#>��"���r�dB	nnjU ��[[��B��.ڡ��|�Y����e�'���%���p�9Ĝ�S��ضC��?˷M��X�ϊ+�ڴZY�[q0a�l�K�뮭�4zQwS�[�"�W�T��+�x�"d��<�����pMb��ʁIĭ&�΀�4$DƑF8Ӊ��7�р7i�e���c:jN�����4�B��1~\�4��N*bv��3a7�v����b���K!J��pp,E��hZ��,b9E�ͻaﯪ��q�$�[�	e���Sǚm2ǥr����޵X��-�	�3��M<�T&�Jv�{�]=u�T�Eso{�o4�o{o-���Ҥ���m��L�d��f�~2��M�eS~ ^B�1��u�-�S.�)s�r��L���)݆�+1�MS];���rE�Pe����E���*Sczt��Wif뾞���ãt*�p�On"t �!U>,aN���p��#RG:%�Gv[�/���f�L�;�$���	�V�a����=�R/K��L>�wq�%�#���ҫ���f�I �'�`�ٸ��u��[U��e�ȇ�Y���cxײⓩ�������!�	���!f�:���Mʩ͇�V�SU��S{�� w��>��]�碴5c����D�v����cd
˲��K�*q�U�(����V��r�zi�Nn�=v��GW�T�:�4��W��V�Kv��D{P,�oJ�Oh��8���j��鋈M��Tv��G{�s�ZZ=t��c���߫�;<���[K'0_��0�I�DS�T`Li�XP[���D����h���`I�j��2.�:-�Vދ�������Pt+Wƶ�^��gԎ��<5ʖv�5�%2܍�D%Q;�W�6a���:�)l��X�"��p�� Fq�96�E�c%cOZk����᪙���ޤ�C����pECsl�����Xظsm;�dDl7���(8UI�8�,YDu���£���.�gJ��s~�5չ��JM`�����88$``敋����@��Yυ�����t{S��f�(2�t���S���Z����zp��^��j����(��3O�ʥ�LQ�����&�BŐ�zu]]ri=��-�7����@����¦K�ygӊ���+�?Z7y�췙�������b*7]��^;U�]ǜ�ok#�_�e���X�]{�+0&:L�OX�J�r��J�=���u.��%��>V*��˺�A�.��L��S��,:�U�F@é���D��z�ͪT���5�n=��ݎc��V��MV�i�N*ʐ�,�cl�1&�0��af�9mi_vA�֡��ᵋe�(s��m�-qn^���y���B��cl�:˜��}КE	�sx��"A��¯{^��Tmp�E�,~���LG��y���~���컽�[Sba@��<Y�^LҧL_�:Xp4c9ʾ�n�~���iNy�q��+��սn�MGǉ���$�z?0���#���Y��L9�a��R�6&���ߛ2���Po������&�D�<����\S�
�U6H|a��W!�'�o�[�P��-���b��r6.	�N�Ƃ#ǉ�z��x-�TP}���3=��8E1Y�瞮�D�V���א���l��HD�CD(N�bee�HE��$�On��X���P��Ӑ�j3�!MF��MfFyۧ��Ro(*�00��/(�Ej�᪛��:֬ !�Tbcx�np�c��N�VC��0���V��r��;�8]1xx,j����M%�A�X�&9�d��&�p��c����<b�ݻ����Gm�
7��<��Y�%Z�gj��vU���O2B�ޗ<"j&`�l���A�ϳ1+W�`�l�l%�^���@U���n�V�#��>���s]p����k���^["��^lV������V��D��ͼ|��}����Q�[ˍ�wr$�f��,�x����\�Ox�O\�8��;��b<�ۼ2�[k2��x��3�i8�N���v�kgOb{Ӹ���S4��*��
)�{�3W��bo�2���X7ܺ�5���� W�� ��rUWD�ҫm�5�i`�^u,��gX%P�ZM;�`�E��#�ݰ��u�����ک�"�5d\ei7��YP�X��m�b
"N;o��v���L�/ӾUp�����#���i�g�f��+;/m�[�V��l�����K�Q)����BEd&&��%�	s�í/P�Ţ�R�18�밞�{}!��Z�#sȢ|�/���X�>�v:��0Ɣ�c�ur�\���Kd\-�`
��������w�o�B�ĭZ��*zX��	���7E����-]RX<�.��`]�B���R�i-��R�bQ9��������������e��������EVz������Qa����j՚z�B3����h�Jc8kk��	hߝ�N���O���t:VT��Y�5s�W܄K�|�c��o�G}�tG�S�/�Us:g�\=��|d���y�5��Ri��@q�O��4ux���v���P��a>UtzKu���쭋�/A�[:�6J�7Y�\q�����%N���ݮ��;�7(v��1��t.�Ύ��
�+�[�;qX�5#�_FJ���湇^�4�9X�Fl[V7���dxH�t]����^�w?������������E8�T���%�D��s�ɩ�70}��c��<��P�*jpn���iSB��d�mt���Ȯ.��G^D¨WDLr�'��<���T2��^"EV]KOW8��؈�.:��쀪��,H�	�Q�aҺ$�ơ<<L�v7{}z��96��K3��X�#�\n�\���J�x�D!����/^����׾g͸��P<�n�eux�1���]�s�&��EʁIĭ&��^4$C���M7w�owrH�]��W	^�Z������c3�q϶SD/�u�N�����CN��ͧ��^b=���r�s��,M��ʸ�?fm�}}T}8"�qQ��T��;��o*��k�5d�}8�G���S�	�g���Sσ�#��� R���j�������S(y���/(Qm�㾷;��I�Xp�f�N���0碩�c��P�����r�nsV�;�q3��9N�\50��j_l�}Lq�"�P>:�����C��#�PN�]��ԑ�����;1��ޝ~n�z{7�"�����V<K������m)��X���HK2�
�"N+K��3���tk��)Y����1!���Q�C���C�v�n,�$相��x�_M
LT����d�l�r�~+���խG%-Z��?L(aPU��D����A�*�i��ub{:ގ��#Bg�Br�d��Y�����S���0�\�����ɯ-�˷�C���Gx�-�L'큮�u����ػ���G�N
�RY��f�fzfDmmWp7cz_�x��UfvV7ssiGf��*�6�C깅X��Vj#����b��ӒH�D�J˜��u�l'��;���rm��ڱme!to��5�@�0��	�Ļ�{.���vf{�;۸2�0�F�i�^n�H�fhm�S���͎���^���j�B�^��e#�;7*�#��3[�iM�I���J�8ަO�q��.Uc���
[<2b���tƻ�#��i(k�	J�O?9a�s�+�n���;�Dv�6sϤ#w����م�R	ı�~sn��3i�'w�e����r��k���Iʌ�CL���e��Y���w;�Je��N�@ї5S1r�c8���Q����,��� *B�k<�;����tc>�|���;`�2����$X ���9��&�\͈UJ<E H���Ux>�f��yE�!�G&��e\�R�h�V�{-���U�P'+S�1LV�2�!fs;�q��p#ӻA}x/IR�!̺�e�������qX�.�"k�%�Rw�yz�_G�<`�1�B���W���1a��r/�tFJ�W��ǕK�&)��(dW��ۧ|��r-�-ՙ�C������"�;���s�o���Q��p�}ԯ6q�������%O�bsO��*(_��k��=6)b��&��>�G��B�cmX��z��z5?O��7�E9U�ƈͱT�_�]���S��+
Ʃ�ܧQc�5'�J��y����Z`��K�Ip?R�U�L(�x�j��R千Ζ:�2���Č.�y7ٜ3vn�T'��W�	��gE"I����	��`
��! V�ˤ�.���~;s���&HF�O}m��c�W���ܤ�aTM���8�:|��ҩ��V��$c�y2���V��̈́�oZQV\j�:��c�c��q�訇BchȌ�=�N��g�ؙ��6	���eSM��i4��-,�Ϫ&�V�A[ub�C�Tiܑ0�L�!@��MJ!��f�t����ӈ���Qu��^�;Q����DW&�#"�|o"=o��@xz���*L��c������lv���y�ݒ�����w�m�)�eH�b��}ȱ�ˋIv�'wA3vA�*3Vz�^�&�
���yt�^�������4,��5���.��?#xx7�ֳ�(E+�ɷ�N��t�K8�,9cE�ڥ�����	�2�ќ�Xϳ�!���ws��[#t�XMh-p�ָo��t���v%�3��4�-0!c����mu���>T4��-���ٛ���
����ǌ�k�k��.�f�Br�K0�EsX�ҷ�{�X[��fGV��nY���Ң��=�%��� ;/{�aU6���9{:�uC��J�Qὕ����Q�!j|��˥s���!G8�":׳�u���<�FerC0:HiͬN�"%�K�'�-����2��6J�6����Øϐ�Z��e�nΊ��;p��4����0��2妷iP�gvdw�vz��p��iƖGEaGۺD]��.���'l�(h���7fR��30�y��Ù��ܰ)����qX:�c߃�8�7O���y�L���('{B�o3�e"���ßb�V�9��>����֑�ca�re>�{$N�W��DY*}��7v/�xAvx�n�M�H:��Ь���q2oE�ڵyj��=�ԕv�ۏf,nj�XX��[�q�y��Sn��:me��O���V��5Ѯp��h[N��P}�q�Lmr��o�����-D�/hw�6���-&�t�ga�8�ʝ���<@�A1�f�%����CWT������Ү�:2� Ea�]��L�d��D�"�HI��SY�ys��,�8,���"��ã*�
�UD�z!�M��V��pf�c2n|k��hܤ��[�e���ph�W%B�V��pr�ݣ�κ�(;��ءp�ݗ90fLP������s5u@&lGHw�]ᴷe
�Ա���3���b�E��t�!����m��Q|w�b��^����CV��E9��!F�m}w/S�̻t4s�)��5�c�3IQXuΦ��Τ��쉄(�����۪(��ŝ�����wD�X*��أ�S�i�slOD�;PWУ�y���vLY�j������]�;S�^���5�#��X��b�˟8)b�i�
�˥;��R���s3�t������jd�3[�Z[��dٴ�uoO��i��]Er��U�o�^4c)@�Cy�q.�P7�[ه�cn�(��""��tq-ݐ�����s�X/n]� �.]&������%���7V0zDqκ�ˋ�tan���T�3���Zͱ2N0&����q�u�o��ެ��]�*�3�%�mۄ:�(L�7F�[]%;���U���/S\� Ou����$��V����];�X��[�[0s�)7��g+�uˤ{��ieq��l&��C`��/���<����p40���Vp�f���r����)EE�jڰ��+���JeQ�-)��r��  LPTDTT�S�a�EPRU�TPTA�MT6A�1�SD��UQDT�TKQMTPSUDU6f54QUT�QURT��MD�DPQ3ALDLT�1f�E�1EQMPDQM4T�UQE�DSQ1L�Q-faD�E51��L�UQSST��2EAUADDEQEDQI2�S�Y�U1�L�D�TASMMMM�NF`dRS410CUTSS3TTE�LCD��E$%DT�U%EC�h�DUUTFY�ASFE80R�VZ�QTS&�*"����*�bEEDULDQ3M1D�QE1D��QSQTdd�T�96�2�JJ�*b���� ������
����i����-fS,Qe��ɵ8�DQ�
�X�("��!�)")�*��(`�- RP����<uAޱ0+&5f�(��6�+��K�C��tg]�656w)�c��[�o�Y��Ũ�,f�k31f�Bj�v�@ }#�U�	��b�G�PӸՐ�L,b�ߓ�x��g���[��B]=nF�W�ӱ$r%�3�&DpɌ�-���#w�Sv�m)m�ˇ~���t���U�Ԋ;ʡ�y,S�$�9!a,��؉�>�"�Z�3@�Ne.:O8�Ƣ^��GI.aB��R�p������n�m�8=��O�;�u���̅Z��y���r��q�F���Z��iL4@L�2�+��}�p¾��౜.�;)�Rc�O[�ʶGf;�2��b�z��#TD:=��u��VT0���.N�'x��Ӣ%`+~�t��[sL�f�B�h�Q[Q��,`���f
>=-��#�-5��z��I}j�\xR�Dl䤳��%ᄹ��֗�gbۯP����g��]z+C��G���39;-h�/mU���t��=�>]:E�zĶE��`
�h���0��4�5թ-��7_�
� ޮã����VZ>7B�R��F��K��u�
��a��#���d�6�S�)�paWbe��(�e��ޥ�o�S�_C[:�:���˙�˱7o:�OL�)+�m�ȷ��-N�E�{�:U���=��^��P޶���B[�_-Fk���y����2�#��ٓ�a��.S�r_B�ḻ/���}<�\<�
[��	�mܱQ�遀ԳWKq�����^�{ַ��+НŻN*�B-N��܇�C�u"���Ӑ�KF��N�����F�w�o5�U�A� P�d��5�Q�Nп9/�ט˭��>�|Ι�:�����7	/OgZZH��	"Y/Q?K.���3�T��zt�`oMYe��DyuB��Pe�oUG�k<%�%��vK
��|��je����1�[�n����e���Q���ff��R��<+JEъ����L*�WDLr�5+}s�w��]Wgw��J�F������JO��:�-�� :�; �# T',Ey�L:�$��P�T�tI����X�>��FC�t�0�2�����a���"�����b$B������]���F�94VC�s�8�K-q���#�&��E@L��J�y�����P��S4��1{]�A�H�]!d����eU���ָ�9dO�u�K�7� D�#i���]�59֫F]����*�/�I���|U��@�<��Z�;q�J'��ԣh0�g>�v�3�Ҳ���^�[t��:�z�7�YC;���x�k�m��x(��������b}��%uD�y�Ć1��X�<���7�W-���gr"��Ձ�����btж
����ͻa��Pp-���oG.��,�nn�����b�$��x����Q��ƍ&x�����un��ziݲ�.+�=�jw{R���N�W��v�4c�ή�"Q^D���w�F�U:����Ҟ��+8�-!�	A@���7[H;����S\y5Mt��1�����Ȧ�/
q��ܿg]���Y�L#Q1� ���b�;D��΄G�w�z�{h[�-�<�-}�D��CvpY��ErXH�4�fB��1����'��R�!�,\AS�`�Gn�B�عf��qS�e��=������E��s3�3"7f{��1��9��)�{�/b����Y���,��Ͷp��
��6B�Du0tw�TxzrB�m1���z���'(��WQ��FK1Fc�.A
y��^<�.��c�� BS&F�%���A\LJ8��6&5�YT�b�t*�S���h�s46�^�����o߽m��t+UV�(ޅ�bΏǽSxK�S���p��\�lX����{�.�4�J�8�6s��v�)�`�2�Q�h�gSͼ�P�<�NZ1&�'�
��J�:�خSP��A�IQx��2>��N�Y��w��ɑƄ�pgV�j;e~��Tx��E/����U��rlnE��c�w�����R%��=��)��9�������'�wLm��"{�G�)m��.믞o);v�@�N�BGi�T>5����>����pECsl��ꐸN%��T��Ł�ys1o_s��5� �	c$p�5u�
{6Gu1w��	4���+��Inߞrth���gQ���߱Omٵ^��N�l�j�B�k�������a�]����>1V�k^�oxǅČ�v٭��cG����X���j�ת�<��VWd�6���]�����(�>����բ0���5;�K Ez�ZUw�i�z��-��1f>� ݢ*Ʊ��w{�Y�bC�5�Dl�y,8^���K0\bj��c,�lbY�#Fmr�=ݫB���rR���߾�W�Z��p�b&6�W@�q�E���*���XV5^�J�Y��1�%9��.��1z/��	��c=)/ ?R���P�N���ɕ.X�K^�]u'�<�dV�f��ǪT����:�:�V��e����\r�Z��=r��$$"k��;h�C�g��ڬ�����L;�{eN�moV�R`:.DN�&���z��q�Q�$�{f���������ݕօ�ks�Z�;}�[���;1�W�� ]6�C�F��a���qp�t9,���X���[���(��Ӄ�gY��%��n��vKFY�p��[~�b�{����W�|��IP���(�����̄�%b�6���v���n��!��6�Hu�c�c��q��BchȌ i=��],Rz��nRo����_'��ON9�b3TO�ej43���Cl�*>�6�����d��Hՙ�1%�j"2%�w10��7�=8�i�Z棄'��9ۧ��RӖ�d �s�3m��Ib��b@�B ��s;��*�G�i�b^sW�1ZE]�IZw��m�]V�����c���b��"}�J&�}�Ȏ1�[<��7~<a� *�`�Yn���K$�\��k�F�4_��Gb�:���K�I3䅆���b�ȶPkZjvs���pU���q��*$�e��uJ�92Br0�ݨY�n�݇}�ʓ�ZKBR�gCzw9�zi\��89���D��`S+�� Ts�2��j\�0��>�����x�i�M=\e��k���q|gM�]�0:�N��"ò��������gb���=�f)�����Քa�CzļaL��i�%.���F���R��fr�y}�y�8�{r"0f�-��!��&i�ru�/����
���N���-��'K��5S2;<�;7�x��nر��Aik|�m�E��2ͦ��ӟM�f�O�		Ԩ�Զ�8?,H"oMlL���1��wg��zʌ���Pb���NuR��Ռ�0�s�rL���V�V��N3]2��^�,,.â��w�}w��g�q�F j�������[G*v=tlU�Vl���\��N`(��-���jʻ����2��Q��P���W=:zX��	���tY��Ƣ$�r�bWUt��b�-k\����&������P���R���-��PНF��qs\`h0�G��L�E��/pij�ry���46�����N���r���Χ?�3�����\i\����⡢��Q�gU�O4�Iq���
��ש�B��h����c/��.
�^���Q[˩�}a(��#_��*	c��E��0D��6W^�ѵON�'J���S�x��ꐞk��*���O�UQ�U��I0�Id�L�Ѹ���LF�
�ja=�������G�j�s��r�����<�]��p�]�pal+�c����R�p�����Q�؏n�9�(�v��\�:�⸽91#%:�X.�9��1Xe�
W%�T�=�0�h����zu�P�n��k�t�����,}�I�^�!���;��(˾�+g]�v�����N�"ل쵦��ӵY���X�[�����qn�\��<��oE��C�t:^8�Y� �ܑH*e]�'�m��dut����ã�.�N�aҺ$Ơx���r�m^�N��o���jpUL����0�#���uQ��a\4��J�/ņ6�̈c�/�g5JmDӦ���Ի@���jKgj�1Ks��%<"�;��5�Vّa�P*�ZL*����QN�_��n$��hH�Q�Yn�2���c+o�Z㰻#d��=[Y��4�ٶp�x�T0W��o@0:ɏ�P���Z��B�/�����<<�[>�T0贷qm���f੭�~b�!�MZJ�:��'8矝�c,�C�s=��ˤ��(Ml]ݩ���3�?WR	=6'T#/=�;�l,��C�]2�e�|W�g��7���@��7܁�E%B�n�<�,��h(���n��w���j�i��j��ط��dNQ/\#��#z�3;����!����i�UŪ�k��	�%nt �S���0_����1w��Q���ۮ���|�_op�tF �a���wf8EzTLw;d���!��}�Ö���ޅ����_�m3�WQC�)ߢ�f����}�)�DD"�Ofl��"����u즟N��b��xJϼ6<�7�������C�lR���t	���[��Ǔ�nUAҦ�5�B��5�^��b��"F͊�jo�kt���:1��ƍ<z祚�_�*��'@�:8���.�dGt�@���)�s[*��6����N1þ�F���+0���¡rn*��q!F�3~����Z��^V���M�<�wi���9K�Pc������F�*5�@�.���<K�^=(+�ưQe`'q���Q惾\�&.w�J�����}�Us�E�5���^=/!�6����6틾7p�}�拋^ؼ$�g��%��K]b�u��ގ�.�e��-�1��i�"����WZ�j&�vh�rX5[=S0��o
l�>��ߚwTCsl��U��I���[�򤭙!iv����P�cc�}�p���<3�O�.�̛#��7~�w�fh�ITs��7�\�4��K�Wn���t��uL\,���HbB.�����c|:RB��Yڽe����i��uj58�4�B�P��:N{��5uL\,����ƕ1yh�7�O%Nv#%�ߨ��8�U���Q���0T't��;��%�j�3��n�4���6i�/v�M�OC�r��+����t(���}t�NEb.�$7��g��uT�J�ifSVF�9�*%t8[�y��Jodߕõjb=��a�*'��;�F��Ϋ�E:��j���h��z]%v%L�1a}{\��[yk���DU4�v�$o�5P�F! �f�e4w���K��V�l���p���R���/��t�a��d|<�#�2>���	�}l�m�%~2/:������Mg��S�������+J��W�
u*���ۯ1�Ij��V�pVp�
�v�%�'b�LO��^쒋*|���P�p��s/Yj�8��=9�Ƭ��#�b�d���RKG�S�}�/ 	T���t�){�)v*!X.5I�P�a:Z{a�Q�ؤaW�`i�p���!lD���,.�����J�ݾ|���ց�Oj�-p�xm����B�!�r6�y�U���(�'�x++d�9������6�4��%IaK��������W9ƂX��aI�rF��v�`s����h��kt����(Jg��S�PJ�=9v�ծj8E'�2�C�O�U=����$˂���E���R�w%��kY@0�/���ຽ&5�*��{K�N�a�o�@Op�I�z����{d&A��{N3sc��J<9�G���-.����~G]v��U�}Z�樃��2檠�M����Dhy�z��:zJb�f]>��r]�sw�s��y�싗Y��)ul�;��g�#��H��4��z�>�v�e�[2Q��m3b�+�Z%�Z�j�3����1�ڗ�Zv��$bx�$��:ro,�J�Wg�j�F��{=O���3��\Br(�\'P�ߞD��o����xV�ݗ�.�t+Iy{I�1�#.���j�����D�	��:�2\�r0ޫ��Q'}���Ŕ����^��w��tlJ�z�R�h�8=�� �y�r��D
��P�������A�
++��žV�G�NU�zp��+p�m�k��ͨ�sճ�^D)cA�T�X��,;+I�F���xM��;�*�K@�
�BX7i+�%%��*��n�kŰ�dV�c7�-f��sNi�-�Ūf�o����CG�̓���h�0��,,���xC��m��kD��tEc�;D����խ!�ﴝv�zBֻѶlU�R�Jǡ�.X����O�7*��W�y�[�ռ&x�� ��A�Jup��:zq�L�5jc6=7E��%��z��vlx��d�V�曯����H���Kdߞ���ހ�����2����^�T�ur6�m�M�ub�I� FIu�0��R��-N����CV�41~+k���z.r�ٮ7�ݕ!K�G^��ݬ��	n��A���B�Fi�����>�,��M�@�+-#@���xaqG��WT�� �N䕲#ƑB՝&�Q�ju�ϳ+Wq-|���L�"��
l{�ń!��n��f��W�t��YL�&���c7b!<ՙy,�Z��d����0�j�Ѵ��0U��^�7�O /75En�ꌆ�#��kӫ�%d��]�{�{Rj�W�����as�Ǵ޻�AM/hX�MaO"r�5�V-��f��-U�A�|��EGI�m8-h#*��l�l�S1b����Vt�:ŉ�;��$L��m^�Vz�t�2�]s��c�EO�ha����s �,�@�3�m�F
[}�j]A�f�tW���hB�02n^,�{�}з݄`�[Ƥ\����ݒ���v��7SN
(0��m3�q�ve��4����.��Y��Y��O=�T��;���[�D�f��V��n\�ײͽ�E��Yt5�I��[��� 5�)t�e��/EG�o3-���:[��X�'��IS�*�c���B��H�yf̈́��I���]�Xq#[Ǩ��V�4*}j���冮[ܪ|�=��V�o��N�\�>ɗ�9Z����y9�Kj�H��رFB�/�zL�%r�A�<
����}5�J�IV�Fe^@��-էwX�A=U>L!Wu�]��(��o	/M��Yi���"Qj�C�.�p��+��������aWL�](����g�1��I�j�ѭ.�2�>B�t�P��76H{+Pη�Ok�3��{s;��\D���3�YEQ��mX݋^K�xbT��_�5=�_���Q�]��|�9�2
��w,M�%k 6r˩�^��V��7��s��)��c���fC���>���B��سN�\�V��q/��/��Y��(�hk�^��C5/��;��v�!٨��U�Z�	: Tۢ�G�%�Ħs�$�`B��d�{�|_r&�"^�L�NИe
��&�Ϸ�% ɧ-���b�;��=k1.��#��Y�[�K�E�*�-����g��Jޭ5����YL���}��T¨�H��";}�[T+5g3�}#������'Ǘjӂ��V��J7�A�݋��S�2��С�"euÛm�)�[)�YjѼM���#�����ug�	�e���gO.w�]
��/+v�0�����&��p�;
��#:�f���͗O���֙��7Ku�͉uܭ�ƆW<�]�h�'�WV�0mFk�k�}V��P�ۉ!�ˀz�haT���4]�%c�����h�w��*�3��K]]Þ(G-�ݜ�̑ ���w�ʻ���[w�tB]��@�|�
Uњ�5�W�Z�:�d���}9t��q-���o^K ���Ǩ��["�iV�5�CP�5�{&���U׭�T%�[�GZnM�s���/2J�u�_u��u�UMD�TUQEU�(�$��*���*("�*��+S�QEM�$AU�E�3Q�KTT�̢*�����(�"�0�h��X��������(�91MPTCLUk�������*b�j& ���������4S5Y��EQELD46YEEE1%U�sȆ��������"��d������$��,�#Pa�aLęL5M������b�X�M5Te�1DDDZ�i��)� ���dDU�QETMULR95�	�33
��A�A�q���*���b$��*��&b�Ս�u�6�(�&"&h �(58�jĩ���0��b*��S�%SM��� ����&$�(*
H�"��5����"��Y��ʢ&��gV4Q%Z̩�V� ��j*��**��YPV�¥�*����)���i������	��bs2Z����()��������b,̬�1���#�&"(�*j`�����U� (
��.�u:Ŗ�u�'z��{��.�]��o�(=��{NL'�5k�]n��O
r�e'	���i�Ǜ��<��voB�1ɥ,�ڑ~<�2tW:$V�o������܇�C��	�,Z�;�.��P�mr���ؖ��8S� r%��,�'���FܾZ�}�ON���*�ZТ�;�7�,�p=�����w�C�;��7�X%
U&"Y$��Q0P��5m@����\��;g��oA��	w��sή�\"��9%ي�r��ȘT��	�RB&�%K
�N���]�|�ic�L.�ĬKިie��(4\԰�:�;"���w,EC��u
�	�`��3�k���ռ�-%��<;�oL �HW;�Hi͆�4�	�XGG�m��R�����i�&�r�A�u�1�G(�.��︋�,��ݩ���M��v���K�)݌|���'��2��"�X��d��^W%
��w��%=f/�ΣI���tӭ/�����8+�]*�0\����ھ�C�T�T�Ex^Ww�xyd���A)��Z���Y��>S�*58���.ZJ՜a9�������yN��~Yu.V=��Q��;�d��U���nwec�@�꒒\& ��Kw���I���QYR��έJ��/l��(�W��Y��Ǆ h��}S��-N��J�=s7�.V�KeA&u5+/����
؎�i#�a��DwHĆ�m]i�=&ᴰ��v�AB'N_�/�	D]eh�FWV~N�F^*{�wr�o�3>�L��&��8����=�y�(��<��w�Mԇ;�p/�4�M���;���B�Ծ٧���
��t�=�Y$Hq�i�;F(��l�.v�A��:UO��F
�fDӇ}�K���Q�-X�w�o�O�dh��K�EV�t��w;d���=���J��vWF^����Ė\��L�>��J��G����9I-�!Z�[���mdר_����@�#�iX^�vo[���F�	�#��LmB�:Gd�{md�`'|���O�旓�-��:��0��y=�XB�r�����*,̘x��骺���k��O���\)�bt:���w�{LF�nhn�R�Sc�<w|/!�+1P!@����qn��$����2A�H�:�bP��e2Xz���s�sw��GGy�+H�gz�7���Ŵu�u6]�0kY@1B�cT���z����M�}!�k�>��\F�
i��ɏaH7�B���:�8��(���cFc}ƼM�M���)�ΕWv`/33��F@�8�[�@L}�6���t�+�0����X�� 6Gs��H6��3�����RE����uH���U�V��ae*�+4nȮ��do���=^�46-L1��0�0!d�5��:'Kے_��~�r�Ut�.�Mb�sv��%���P�ڀ��t'@h�uLZ�8]�HbB/���ke��u�YSٛ;�d��)��|������u���GI�s��je���p��4�oNmB�uE���nv��t�6�����l�����jXwKA��;ǯ�v�/�+�9u#��Yy��E�|�����Vi���-��ޫ'���R���<��:��ɶV;�o7���שL�Z=Y�1���0�V��R����e��m �ҩ��6*y���(Ż˳/�7�v���`�~x'g	���>ļ0�SԩV���:�G����!��_cÃAF�!�>'<� ���x�g\u¬��&�,�K�I��~`����ś�G���x��[ۻ�i^3����L;	����F�~�*�L��$��{k޹1�k�x��~.Ta"�H�N�+uI�-�xo�d�i��IȚW�������5����OOb�Sy��|�\B�Gsmv��\i�%^_>�M�<�����]	�뎯1pug�@���ӀҠpoTɩ�tm��BA�F.E/:���@���:�w�;�Ô]̬��U��tC�ɼ{:��s�\ᮄH���շ��C��T���%ۖ��Z�j�KI; ��L�WR��j�=8�i�̇�D���hd,j�^9�F�������ޭ����#��0<�8�]�Lr����¥ONC��5k��K��糨nǘ��WY1����b�e �D;� ��A���	���=��Ӹչ)G)��it�|�9�\���p�iH�9n�D�Qđ̔Nze�>Cvح����6��Y�����y��CN2����p����iȣ�i�>7�%�D�̐����u��q�ڍ���ӹ�h=4���l\w:$��
êP/���*!9j�B�vQ%�t�����I��s�;��V�_]7^
E.׆V��n��_ڝ�iL4@�N% 9�-&�K��5{�fwo���(N�g�E<;]A7���͘�{ճ�^B�4�T��� �54����e=�N��$Mi/�P��dS6y_�n��2X�<=����f�k+"��E&��
4)�����k�p$n�_�e!ݱƎ41��'K���w3�d�]]�r%��Yt(^���F11�����.H���y�A���4�N��=C3qMK�M��{��=4m��
1y�uO��:fH�9�!�,١���Ir�aҹZ_E�Ѿ9y�L1oA��Tlm�4b�~M�g@�Ib]ϗ.�Ąʹ�8T�y�W.,,�%�ͽ��ٞp�7J����R�&��c�����0La�R�&p;7*t���׃�Xܼ�؂��{<zvPw�N�D鳜F��mmR���´�K��0�뵍fW;�8mʤ\��%2B�[%C�b+Х������НF����2�����V�V�RKl�xL!P#�����W�p8TxZ(���X{���u�ug��b*xA̭Δ���\Z[��.!\�����4<OU��e��du+D�܇�C�E��v�Zz�W.y�:�VE�r�ND6%p���/��ED��0c���awϼ"�W�^�|���f�.bY��OoKf�k£���]ap�M	�����70P�g����/w7ub��D\.0�'�:�5uu����ǒ��E��<���LD�N�QJ�	v�_v��{�:*�U0��j U�@k( �N��XR�Xtv�ܱ�ø�7{^�mkRJ�].�$�P:Ke��T�W�k8��+���TC�6W�"�q=�$wd��6!����u�:�kg�
�����mwR�ȝ�iHʻ��1+,69�U����8����u6���Jf�PI����Ryh����\�p�o�⮱b��Z�*��z&�MǮ��M�B��c�o_�"�u�;o8x���V�h|�7�9b׽�#Em�0�{	���6b�nu�)K��Q��28�(#sBpJ���.��7�藤�0H!�,¨�'n*W����ً�q�v�!^DfxAfoG#��Ta.!.���Ӂ��CO:�oi�"®���X�7�(CeTzޡQI��\IF�b����Vk�U�8Xś�I@gVi���~�Ӿ�y[&���MH����Apu�&�+��͌?tz�^�)���o]�J�6#/4_��k�3�y�T�V��D�g���7�4�ˢrg�ٞk����4��)�q[H;�N�f5P���T��k.�z.o�!�N1�ǫOe���	��4ϕij���<�BnÉ��S/Jsv+���eՐt��|�gqꛎ���Y\�n��^:%�s;E�R*�S]J�֮%�b>>.6�ۤ=ɺoR�1���`|y�S�F1�θrp�)@�3��4{�*�Z=>i
���]d�2��;�9��QF���T�+"8�K4�u�9��#v�T!�LmyU5zHQ^�f���Be<�{���ӄ�f�N���B��
�)�0V5C ���� ���@g&*���U�-���N9�#��׌�}錬;�fWʓ��7J����+l�;��M�j*��/��:�MÖ�W8zL�е#}T�MvV��3��[�nl�
�қ�)*ffꂆ8N�+uP�ũ�Og|�TC�p?5�d5����
��f�Ȑ%���
Y��.Ūd�����%]��wi��f�l�1�	���!��x�N;��dX��ե8�id���%�Tf�A�F&_�C�Y�oX{�u$�0)vx;�3��lOm�+��v��;�6㲀B�  Ʃ<		����ƣ��6rHF��;�,*|M.b����u�\�na��2��'Cb���wT�,B+ah��4��υ��wt}s�Ü�IjaV-�A~���nX�Iݨ	�GbӠ4S��/вN} E��B��z�uBw�w�/	بP�����h7�I��P��BX�JN��Q;�e���Mΰ�(:H�W��w�+Ջh14�����բ3ǆQ�������_�N����D�C6�t��S�d>�g�>L�����i�C��q9k�2��;)�15DJUG�I�mUڽJ)ۦ��ö���y��^�W��ڱ�"�ޏ!|x!n�ݒ��S!��߬"Զ�����oM�J���ޯQ�on�W��]wP;ʷ�;J�n�_Z9֙�Cx�͍�Ʊ�Z����]�k%Е�߰���^����>vMv˹*�<P���;�P�[*Hs��&�B�7�[>(�5r�[K�4̵#Cx��up`S &1�o�rg�)b1E:�������4;%�L��պ��/jU�|�v�h~!3�2(���:��J���-8,jȺ�#�b��&�'D��3��v�	J��-���
�@
��#�+Ig�7��t����Q�ģf`i�A8Kg��uFٔfs`So/���UI��N�;�UM�.	�����>�+!�r6�z�����7/�/�w,ҩ$#C%��+��*�&x+�TP�N��s��f>�'Բ�zp����'lT\LO�=�n)Zs��4>�]BQ;��R���×/a�;LjfcDY��,bC.6�bZNR�J��h8y���C�B�PT;�) 	�u�L�np�Vq����<�IYݍ��&x����L���YL�sk������ylX�y�;G2Q92�t���h��|j6%�3ϏHg��N����PF�9�un�d3U/�ȣ�p�C���I3�HXzi^�؜�9\�imWf���e�$f��t�q��^	�9�2\��5
�I�����P!�)�i�G������U�	K�f�c*�F��'d<�i��*P2�֊Qbӫ�(����+kEHY#����~j��ØJ���|l���nS̚�<��]�e4�2	rX�U)%��U�
���dG����7�ԓ�ȱ��/0c�oSq�G.k$���_�����𐻋�V��V��gz _*�z� '-�ۑnֹ�+���ص��{Ͼ��j�#�8��PX򭘨�ͨ�sճ�^B�4R�*���iOONm�O35b���/I�G*4����l�kt��e���D����d���}�מ��y�$�oJ*�.8���x��,`���:��,�Q����2l.����{���3ev��;+�t��3< �؜P��`��q.���n���FٱV�-t��z]�`]��g7��]����\G*X)���0���ҝ\,	�ӌ�ei�E����U�ɬso�oxf�����g�U0j�@�2B�[%��"���x�-v�/T��&�YB'E�x$�j;�͚tx*�����Y�ߨht'%��a�>�D[���e�ELM>K�f=U���bZ.����tK�POU�Dr5N�:���n�A�K�N(FRh�A׹�2���D�u��S:g�e��Dp�C� LG),��<��8*��0��n�w�_��3;4�H��Y��p���ڒȾ��L�1�PGh8��h1>��8�{�l}��'�)S��=.��a���4+$��zl���=6ͽ+)��Y�R���ksb��Y�n�V����:bCo �l��[�����j�<n]*� �׭���m�MRHT����<=;hX]5e�����Z�wf��J�R`O�Id��GYK+va���%}�%�Z��}��{+S�:��p�f��<�f([�vnD¥t`#5����y��WZ�RF�.p*���� :�5�E���@uHv�n�C��{!S�O\s���D�>�$��ɦx<��c�;k8��U+۪�wl0�9�@��k���T��ݴ�*�A��R�&tOa������֥�0n��JN@�/:CTh�ŏ:�r��!�T\PV�@��BB�,����P�9E��w���G'ĥ��wkuVi�˪4����;p-�i��`h��cE����E��YY�f��P�:�!�}Rv%%�R�Al_V�p3�N��\�/�M�9�x�g����/�ܝ�	�O+N���:��ָͭ�C7�YRp����P/M2.++Cdg����e⦁�m�i�J�{���S&hQ�
�$,B^�;�gI"_��b��]�h(4�M���;��L,1��<�@��D諾��۬ޥZFJyMk�7�I�{� �0��`|)�zp���ef<��9 $���s=�(:�&�٫Y�+T.����;*���,O�����^�ϊ\���T��Z�5S��ޗ,��U��{����K�q��(mG�sc��]�D�q}�\l�xh;��1�+(�*�ɝ.�;N���]����N�5\�yp:�^�=}��A��J���/Q�跗�Ws�M�2���ϦW!�V�˩����N�ʭS/N����r�QQ�����Z�1e��[��7�I�v��</� wYՐ������(e��>GUe���8W�'��٭�^븳��{C^6�^�l+���B�5�D�0^�b��Cff��.�;ø��./�G)W���xm��{�t@�C��k:�r��ظ1p+&���)}�@SMBT�W]�3/*���ˤ�2�-�N��ҵ�v�A�yVK��j�V�sr�YS�h��3gQ�y8��� ��αU:�v�_@�"��I�A�rgLC�Tu��J���F�����`��:/ �w2�Ik��N�w�A}wyϱ�|��<�k��S{��Hc(��m�l���S�%��Y�y�`X7^a�#4&]��N##x--�O��;9�+ӧnO�b<�����[A=ԥҢ^;m��{�;{�Q#abkhI�c�����}�!3Y���D'��*y�T�%�u��<z���>�kp�nY��2K�kI�&�4x ə��3��Tۓ�c����ިH���hd#ȩ��]�'(uX�ca/�m�8������`��#�a��Q�+M�JE6�"˫$i���G�;�L�\ą��yr��J4�
f�fm)� Z̡�C2,y�h]�ɚ���Uc[�LWܞZsq�Ѩ0`��_"b����Um��y�f�X�&��@Lo'�%�/��veM���U"s�Õ���r\®�ٜ�S��X�x(nf'�)nU�l6�̱[>�ͫ�x�j�6�ѱ$4g&!!<D�Ǖ��Kcq
��
���ە����w���oNh֡��<W��V8�85�|��i��,b��&�42�����d-[�Z��E��v�y�[7�H�v��(��K`��+p�Ner�^�.�++�n�����znJ�����sJZ 5+�C�s�o'V��kU��ON���ҖC�o;R7r��vD���]`���]��MIt��,��We���d�jD�Pʵǀ�+@��\�7z�]L��&���<>(l;�]7�N�v[;�kY�
}s:��dYm����o]!g!����59pWY�o6�]a�4i��:-��O6�7�t���M��%o_=ȡ�g#tn�t.Wd�R$��DR�2�[�����+�r9tA���Y�M��v;\��6���l�9S%b��TNjm^_۷x�u+{�oJ�9�<�W}�n�G}w��_u���j
*"&�j�����*���Ȭ��"����j��*�ə�����)�32j&���,��s1�02(""��#3 �"b`�����*����$�0ʠ���ʚ
	�h��(���3�,�1��#f�+3	��������*� ���&*�20�&"����
ƪ��**�#(h��*s2��0��f'	�rȲ��2���l� �,(��"
#,���&��X3���+,p�h���̫����,���2*b+3&����1�+
�(����0Ȉ ��3&L����L�'#&)���32��**��`��3�,��*���(Ċ��# '0�
Jb&s�2��+
"��p�0230�0����i*p�,,��̌�l��#2#,J��31(""�0��2�̬J32��*&(��ȋ,;ѯ�7q�$j���e�6��!}\U�����	Rgu��◼�Bgq���X�Xi�ҵ82m5I�[|�.��V��N�J88��>������W����c�L(������:�W*�u{��jd��~�$�6*)���ԑ�"�a��^ɘ��Q1�҃%O'kPn��0�.Ņ/ܬ��,\둇���;�8\D؞vJ"����&���q���۫GZ"���p6�b/K�YO[�r4�Lp��Lm*���I
*�5AvI]���U}(*.`�u}Tª��-NR{:�S�W���#va���!�&B襶���4�����F��P*
��Ġ벑.����r�nu+�pSc�C�w��n�F֫��w���������ف+��Q5'�똔;�Y,t=tQ�i�j�6��f_��z�O� �8���|�ď�'޶
@
y��/�G�u�]�74>�+�V2 ��o �z��@���h��
�q�'Cb��^wTV	��Q%u7�����r�S��kR���#�>�pI���)�(	�Ga9���8]�Hb�Dw[�ho]��X���*�J�cm&F��4x��46��v�m�u5��+(�7W5זvo �@$+��w0���](�"��M�Q��r�R��Sn�M���2��5A�:+��fu��b�"���d8�iS�ݎ�E��R�c4�9�L��q�4����WĔ{��B��u8�;��
Nm'#��5�T�n�)�A�v>d����ߔ�|i�U.&8*�߬�ɸ�gE�<N�5���XS M�Ԭ�<�]n��<;:�'�p�8(�(�	��i��kzh8^���h`�B5E�0@ն��9���4,�z����ئX�V����ke�i��B&:�R�~�1��}�R�Z�hh�r��	�s�ta��6�V�jX��6,?<�8���c	�A�ݕ���av���=s�A��6�0��ɕ.���Ζ��l����؉�LWl�*�tR#v::��m��ۇk-�= 5bP���+	fل�t���B�҇�H��y��������X�cT�T��.vh;�2ÿS�	L�H�>���օ'1��|i��Q`��2�zH�a�o�o^�	���������*�
�=9v����D���hf��͞�:K�ej�7�-��EQ#qU�
�Ȼ���Uu�PR��g%��#�K	t��!�O!R���S8N/#��� �"b#t+�ױ��E�L�wL��X��(��j�q�ʢV��͜G+�`Z�&����P�`n��9�Z
�F���UʊtT��&�qԛ�Uf>C� 9�ۮ2N�o�E��|A�#�,�u�'��C����)��ā1�H�0�����)����n��-� �3��}�IdC��0���V�����wLP�y�y�D*�#Ŀ��Z���~ȅ�Ճy]�{��U��
����L�C�sN�s5Q�ӑGb�:����"X�rI���V�>(��ͬ��m�8xS��V*����ǜt�~�tI�	��uJ� F@��a���=��͞�q6�{T��l���=��N�o�J�eo�/܌�G���4� #PJ�p��n��(���m{�mU�_L��j�������&c��r+g,�X�m8BJ��T�_s�Uu���?.�d\ei7΀����b��-�뤯�p�O�����5�V��1㚋S�^��E���f{fc�RŌ4`afI��g��̡��4��w]¤ܪi��r��WjDV�q~���oҝ�fB�5mS�mmpۣb�*�e��S`N��FLV��4��cz�m�*P6��S!-�s���N�'/
�a2�����f<�,yroUo[�C}�fr��[Y����4����ք֓��P�q��n��]��j�A���[��9Hy�۴	YBj���K�o�@٭�vb&(z���\W��Z)u�)l]��Fv��z������{6�@*aӤ̣ӱ.�.\ճ�J�C
��+�y���\�=�%2E�h�ɸ���R����x<�M`{��I��Q�j�n�jOȃ�a��%TI��2�p�h�ih��Y:�L��}�a9֥���,�����ON.�tH�uDp�tN���"���U���=m*MJ`��T��yS�&#�`���\��pWX��Φ
��¡А'��K"�T1�C�@mVl�[�vz3��Z{�������dN�5tՖs���Z�����:���������2����I&o3��~�xP/��ơ�7�nu�����f��<�f(\C�vnD�G����rlګ��\����F��!Q=,*��:�j ]��Ƞѿ:�ad@uHv�S��h��,��mKiOt��;�'�Ix�emOu���#}�]!\�!�6X�1Π̘1�Y|���v�}􋂃^�2!��&A��l9s�w�E�ȳ��<-�7r��.�I�6��O}"zk��m���]���00 G	�C\��=k�0�\\4���Y��+��R�
�:RL}���3]f
���-�a���̫0��V��.���zMGܡ��^=�lw�v�T�]u�`k\G�<Lt']��^�{���ǦP��b�nkM�����m���`%0��,�l�ߢ�v)�t�{����mDB�F���������f�o�����غ:����o�WRufr�q�j�g��x]�V�[9E@\pC�N*3�J�9�x��ph���6�c)��P�����\u�i��Ż�&8z�dᱯ.���H�����]Xs"/qS@�6����/9�s�L��x0��5�'��v��Ӥ�7�<"��*�5�&��q4�L��uBɼ��v�s�o����ʼz�/�6��駲Ʃ�#�e�2Lo���S
����� N�O�*:��ׅ���0c���x�,t=U��++��LdhuG��K�EV�k�V�����,'Z�*YֳH�]�<x��!��_.
u��>ΩbxT���x6@�qw��74҇�7�u2#�!Ur��^���,�������C�P�T:J���8��,甧�l�׭�]V�Dl0pc7V��S0����w��W�r������F{�2����6wf�(�԰;2`><K�EJ�A�)��i��nr�n{�_	�F�!5���\�Lҝ�5~�/��I��n���+JǯvS��v�Ӥ��+*4S��*g��4Yt,�n�A>����
ٳ�+Ur�}.�ˈ��t�̑`>�u�1�M{ڒ7��
2�w��Nc;�E85L�(�;�:�FS�uy��Fov�{�\�Q@���ouV��S�p.)�0 A��,�9�LJ]��b���F.u��999�-��k�3k�J���18G;�6�� �xP�I�j"Jg��q���M��o8�J.�	O3c��-�qƧpEy��ad@uK�pdd3c�uA�`����RP�RoL6��F�n�O�g!t�sa�>��߻��&��b'v�&B9���XŒp��FM��|8�U�En��G�#�gS��������s�MjqPi�����:O24��P�ދi��f�h__j�\Gd�;q
@�0�̉����)�Co����Q���< 9'w:C��$����V���i���-:��8gq���O/V����9k�0\��K�.�uobli�S�ؿT��,���j�>e��&`Lt���J��X\u¶��@;� �Dr�Ugo*S��E��t�~�N�	���b7")���4��>�Ixa*�k�0����������m�~�a<Y�^Lו;�2:Zs��Ƭ��B0Ȗ/�M�Pе��^�en֧v�&�c���]yy{�}�ť姒��S7�{:ɶ=M��MH�9�J,`fQ��.K�8'�u1�sR�1�����(��+���PS�wz��!�f�!]ʍ����nb��C��Z�ms^�؂v�њl�M��.�X����P�pr�s����s�������B@�%�of	���
�F�R0��֢�vV�T��v�JK`ipOȞ2ę�)�q
��E��x^�Z}�VC��ld����Y�
�w3�Rv�KxZ��h"02Q. �ؓ<�%�ON9�b3Q-�������.�}˗dՕxoڦ���:��~��u͚�h����>��V�Y�j�=)P��ݦ��X�JQ����̡����x򐻇��H�]ت�wVV��_xy<w�X����]0��L�+Jr�1(sW�x9��q	˳��"X�bH�rQ=o*R�A�m����j;׽�"d�7�+�[#�(<�\Ө\�Th�NE��N���\��r���4��o�5���ܷ���52�ƚ���A��D���a_��P-92Ҁ�4�u��4�Wݓy�<ҫ�[$�:�=e�-��u�K�̔8`tw\�\F�`�* ����פSOSU5�d]�@�@�W5	�p�B
xy���k��3���p���u�K;��&B��1�5e�_5tr�(�x"�2�+@nͬ+�Ol��jnKCsh�Ө�!�`�dU����}��M�8�I�`�z���7�����(���"��\�����o�t�#�Ԏ.8)�*ȝ\���s��{z.�2��8�u�жqҀ��ׄ����t"C�L�0)U[�^l[��I^7e��e8b w����@�4T���T�h�=G��mF3q�+�M��C�bX�¸�c0�/�3�o(Ȑ�n�P|1���\��DI-9b��]���8Q;Q�ܧw���ME�Lw�[\;"��.��/]��m��2��n�c��k֨	�X�ȸ[\ �A�����2�&{
�QsF���'Z�3�f)��>.�p���6�J^z�����w����\�,��u�r�?Re�ٰ�Ǫ��x$qq�5'�dP���Q����N���]�hd]I�w�|1U�q�-w*"�f����8�KFW�#]y�4:8�2tW +x����i�]�1Xr[������zJ��8;r;��/z|��@���tF� �|B"������IoJR�K>̺9�0�u�G51V�^QvX��󻎳k�J��鎅�����6��ob�h�."e�f�
5�jOeg��1������o�����r��d4��hys հV����vM��v���Z|pn3�´XW�u	-P<vP��=�1�]��gl���6(���Z� R���%�丫:�ܓ����^�+��H[���$�q,�&R�:��:4�mjQ�0
Ӕz��������^�U�ȸ��F�r�5*XU2�vL �vP͢�E�K�Rܬk3K��]��l��P���yQ&'P�$����S^��d.��n7U�䌀�V8����mM��b�8��L�q�%i�6�Ȇ a�D����]SyQ��bw�R�휋�&��J�z=ˮ	�Vّa�P����@mxА��!�u�z�O��xH��;{���o:dǰM��w���m�vdt�a���lbv�[6�|�[,h���\w�_��z������Z��a�#]���uӔ\�Djq1{��'�t�g��;={ǩ��Z۶��,���d�C�iZ��q�ba|Dv�{�]S�cһ��D|gz^Vxi�=\�t�6�wU�<ӅnK�W̲o��� ���l�!@�*��a��.����&1 �}'W�P�>���U>�������4�ĝ��
�����v8y�Qξn��B�a<8kUO�:�������)FF����=),g��Uh�8Te��%~&���z{�Mj��Y���}b�
ʪ�:Y�g#�9�G���ԥ���a��%�tyQ��837�e%=���t/[f��WO2aV2O�L�:��wb����{K��Z�Q�q�B3���sD-d�jb+=���I��ؗB���o3�-�Y{D1��,瑄�Lg:�8w�����(������@ou�ų�؂�IП�dC�꤁B-���If���vp1����B+΄ƽ��uעż�JV��⤅ �ѹ���2�*�Xb��'���r��y�Z�cY�N�V�^3شr�'KDsT`N�K�8��bPu�H�p�������V�s��>u̓�޲_�� #E��x�4K�}�r��
~�Ĵw��K��Ge2Xz�׎�(^�]��+��Tv57z; )vx0��鍿<��@1�ORS=WU�f��17	���k��X�!�%g8�4�Ӹ"���adT��q46/�a�u2�X$�B:�Wn�����S}����� �׾|�1s�����pI�7,A����rش�Z���[�L��z^�b����9�Q(8P��T�e�XCFIcu�%�q@��7�id�X��ۣ�2zn�Ĥi~wU��ےp� ^��*b��h!7yO
��Dg��; ���ek[+/��t:�5d�#E.�?:!Ր��K��+�6K�p��=�eZ�l���~�->	�hǛ�M�^�	Cƙ�f�i)�4�9G[5r+vի:5ۆ@�,5�P�\��� �Y\��ܻ��g2+���[����j�M�1ͻP�<��L��x5�ڊ��IH��1������iWu(�T}g�A}eeGq_Aһ;�(jpЫ#�dV��2V�;ښ�����*؏99�x��m|(.yh��%���t�o� R��I|��y�a��x�:�8��:\�s��e]��W�K����R"���m
/.�NZy��`p�%s	%Cx��b��Ĵn�F���GʯJ�j��M7���7�4��`#���5�WB�
>���Q
���Z�Bi����xA���.�^�+t)���b��!����@I���o���OV�YI
��hdk�xm�U݀��5��e�+�g}1ߒ*�c:`��)x"]�'�:`�x�9�q�6� x⫖t�:�a$>ˮ��ݭ�\�QyWΏ� ��/cס�#������ȫg�.�T�0A��5�V����#���)�n2�e�6I����$ݮ�Jv'W��.�Y�^�СJ�`�;��GTt��Y8�ުnBF�#����Q�X�2�Gy�dH�Ѫ�?/�T�?H�ٿcW=v��+x�9�p��wF$��fޔ-ҭ ϺLӵ3��ͩ5I���6HMdVa�y�f��/E��y��^���[cl^�`k�>��C4�g*��Y���i<+�`�l�t��׹t�,��F�d�xs�]o�k�H��dc�6���[ڑ��JØ�K�г6tZ)`'$$i��&t(=	�k�ӄ	���7+�䕜eM���!���J����܏{k	V^�>GF=�ia&�k5�.+چLEy�AV�,�
��+kZ��f71>!��7ף��8�t�l';�ܲ���0�"�*���R��$���Й�Ϲc���H[Z�\r�
;�.8�u6�ᕹ}h�܉�'s�	�ul�<*��� ���n[��is5q7�a1�d�ԕ��[�u�U��P]g^��+q�;�{Xn�}����Ħ���EWe��+�rL}z�b%T�S�g5��ņ��7L��΢�Z����v�l}�x�&�51r�fVu��;��V)`
�d� �I��;`j�Z�gY�V�fV_6+B5ok�i��F��:���|汽l$�KUm��\Uv-�/5� r��1��n�lp��-P�+��90���%e�[OY�U@.��TY�y���f�+~�]�n�O!:�	�S������9��m.a�����d�G��� ���n'Kc}|sK0`f�����ά����h����^b����ʁ�j�Ue6F�k"7԰e�[��sh:�u���\H8���ې'��d
$:�\(�wY��X;�7՝ֺw!�j�h�h����{uЍ�E��H�,��J�ǔ�us\���.�숚30�p�*l�̳��hl� �!ʌ��2���$���0��#1*�,"��'"#,,����$ȳ�Ƨ�%�"����330�Ɉ�&l�
(�Ƞ�	Ȍ�,�1�,���#��2����(�*�����#!���','0,�$¬��,��2&32���3
���r�ʌ��3�31�ʲ��0�00�"2�0��2�,k#2�(2�r2J+���̬���̰�,�,�X�3*���3c,�L�
�����*Ț����\�,��c3"��2�"�f*2���&��+��0ʲ��
�������r
+ɬ̣32��i�̰���2�*�,��2�"�12̲���0�#
�̌�3*,�2\�22*�,�(ʌ�(,�2��$��b $�"5tv�Q�YJ�������}zK�:k{���xn��H�s�.�%s�`z�y�$¬2�M�t�L%w�Q���7&���� �����r9N�Ψw�p�$^��u,J9ch�r/z�8�� �+���/J�L[�%X�cY�lQr�|z���ܰl�؆	Y�1ҩ+�y�Q��Kf��fĪ�����w�=0�Qq[H;�T����Zo�#r�`�o�g	���;E�e$�l`�)�J�.���u�D�A��c�8��7�U�ʗTƞt��l��"�����z�KY��Z��o�-�IQ�o�<)���a�:zİa! V��ø	���	��#�n+3ɋǖ�od{�6D�T<�t��}]4��uA\yU6H|;=d�i��]]L���9�Fg��mj����'�ʮ�V��`TN�� �e"�t��eT���s��cnѫ�9-�w��3{a�Uܸ��F���^�9�F��H�2`E��I<�0c�OIB��O�Ay��W[j9��qI;Lj�5!>Wt9㧆�Rp�b��}�HDp\ ̍��>�^u�s�}"y����o�DsOiy�ƬsW�3�|��;y�Ňt|2� ��L�+�`/�I��pvu2s�x%�θ`(,:�nkCo<���Ҋ��7+�|N��]j�ݴ���" �f�J8S�@yU���jCR��	Lfw+;�H��t�Q�st+��Ғ� �d(��O����M5�`Dq���֕�ផ�E;0�~��!I��6cs��Y�#vx!�۫w!���~��QظN��{v� `�\o�M���$�d�g%���Bt��^s����tI��aXuJ,t��}[�����H�>jF���w�I��h���yh�����R�p�Ӄ���tAjkU��6�ꗢ{o�q��>W�����. ?��u�:���l�J�Y���������v�Ho��~^��Ǖ^-]�w�� ��Ցa�ZM�:2ra��Zzg4�̡�yc�����o/76���u!=��Dxe�������:D�F<�;�X�Æ�63$�|�E�+44rM�鷚��oMa�("jԠ������.v���N�3<��Mzۦ;�ŭ��a�:�Ü��v�t�t��G���ϒ��ūu<�U�KdZ�����A��t��StZ���3fp�٣���a��Y���:rNQw끫�c�Jd���J���m�N��v:=7�yE�ğHFʔ�ê�M	�n�stx�P���1�e����&��M����:A��@PP�4vս���x9����e�\�[�]_�lЫi��	kU�<2���#�T3״����nPzx#=����x-E���ux֛,�A[�*�r�[B��R�V�Ȗ���p'J�݇�>u����Vj@k;�Y�l��%�i(�Ή�nX>��8{�_�Ud\�\%���d�p<!T#��Sû���)^kǚiȧ��ln��!�y�ⅻ��LJ
���� \r���1���W�6�t;�R�7����|A���
��Z҉�V9���|�(�<�"���㬫�#�x��1l��kQ5\�I��\�I(6w��V�W
a=��uLj.jpj)���"�55�stb�Z����vjL�ۂ�X�t`O9!QaT�ގڀd���"�F�]0��f
���ĵS�[Ҭ&PvtyU�`����"��T&����;�o��/*Y����������<��okܥ8E8鰂�e7�ĭ"�mÿb�X��=���kb��k�(�,�_N�=�&��D�OS9�s]���j1[fD9*���ro�	pF��U��ۣ�߂JU�mK����U?^fj�/v�!	:�%|���c7�p̈́4�;F���89�l�Z�ɽ��}��f�+��%���>C����/؝�o�<O\��0�� rٱ��0V��;�w\T�G����J X�4�YZ7R�� �Z�ܸ��/��݁]o�w%D�9�[7�ͬM����ۤPQ�Q�n�V�]I�ٵ
��lZ�o�<�ni�ZL��5o��ް��/��譋��AX�KݢX=� ��W,#�r�ρ�k��K���0�"|�����z�zw�n��>P��������#G��|o*5����]��d�(����a��9�h(3Jd�.i`�b�>�n�tW>Y�\JWc2#�B�Ծ�^��������(QvE�v�6(h���æF�pxk��V]㷘m�{�d�sh[z�dVWjH�D���;E��f�L��µ��f$C�Q1��("V��=��aŀ��p�Lg[�C��؞2P n�����滔j�I�0pc72ø��Q�Ip�c/NC�,�<]n�x1���0�I�a�Փee�v.ih��
��EIÃd�A��T��Xb�NR{;��G�r��f�ۼ���W\�	�|�YVXAѤ@��L
�ĸzPW���K�{LF�nhmԉvp��Ml{�x����%��z-������Vo��BF�$�GTLl��3����v�7˫�ݶt�������ڝF��7z:tts,V�n�w !�����%3ԣ�j��-��f7t�#�J��P���ݔ��,��=;:���cV8V�j��X]�W�<�)J��[��wLb�u*]] �"�� ;O6����s7�pff���Fo����r��xk��Yms���	�sC8ŵ+��w����;��1��\���|T���QlW3��#vӸ"���0���.8�M�sm;�_�	 �n�Td^^n���g�b���G��������7|��ܱ��P.���r�Cؼ�;����ʎ�r��Iè�0!B�9��������s�OF���B�Gp��;4EM.��6v���g�~����7�И}���4�*�)1�T���|�v����p�P��ß#�#�7�������H�����s�n#�X�Y�8�e*���7���;=ǻ��'N>$�d��e���W�2*���3C&��w1�\5::㳮F��A_�q��K��Ua���Շ����x,�ڄp��*��\(��ʧg�ӎo���q�b�oM�{��Z�t��s�N�����f�Uo�7�PP�"��J,�&j;�9Xa��s��!'p󎷙)sV�i%��}�h�tJ;3<Ӡ&:İa! yl�j}0�9Xwj%��4�v�
�;(����=}2�V�Z�0��OMrg��uA)����a�zO����C�Ke�V@���u�Tb���x
n�*:��q�)X/�B��<���*�E�ڕ(]W��9�4E��M�u<�+8id����c�pQgT�1�W�Nv��[�/9d�w�����F����n	�,�d�੺�>J��]�,�K�G��\v;��2�W,�IeN`��6.	�7��#E��%@�'Yw&x+��E�OM`#�5�G%x��K����S:�-^ȇ0��;�5L��
 �s����L���e3;���9�����ӎv�ձj8E'�2�C�O��B�� �yؐ'��^T��smqWj��[X����#e��l�<�P���/=�ƬsW�1Zo�˳��-��%�<�n�D���\��ݮ��?u�D���4!��/��]A�<�mջ���F��r(�D��e��yJ7I⮷�Z�=��g�:*!\�f9I˞5(Li���r����&X@Y$9�[��g�>��]���5 F@�R0�J���'���>�ז�˦납�\4`tz����phÎU-rg9n�4A}�`鄈��P���C�vQ�
������5���-CN��Z���K��v�ژ�.�r�g�Kj� ��MY���s�"}��_�V��9���Gg�aesq��&-v�	����Y�[�\g�j1��\��'���cG
�:=S^�a�g�_5�h�(r�����c�-�13_�k<d�u�ˈ��
yJ��%Je9��_m�"^���C9O$�m�k��������o2U��,+�y$�6R��E\�f�r���f�l�7:�mm5��s����:`�F�6�pt2J�L9�q��d7~�CI�Z�*uہ:xC�;Q��*wq��,"jۦ;��x������ʮs/�f��b�+6Z��V6��S�l������ҝ\.q�)�1]��7/���O�k|{��YgŊ�K�F�w.��P'�bS$Z�-�G�[5�!kwiaQ��^ӊ�c�Y:Bu�w,q�<`h0�@���1�*�\u�ʦ��	�K1�x��m�_���c�
��8�KE�#�Q��a<!*��!�[wpe�}��ܭբ��U
�+d��}d1O9\P�s����t�FF���@BTn����[���R�X�"���8�Y��i�3��,zvе�VY�{����t�w*�nnz�������T�	�șA�s�Eo��'��:�5uu��i�B-x�-�L���ʵ&\�3AV�#�.^���k�q��m���(4w����m����7k�$�\��d�8<���<WD��Ai/��G���5���Mp����s���Y;�ٷ
wo�^)­T�	���~ۨX;Ա�%a�m���n!wi�ʽ�%������X�>�F	�ljF�m:ˢ"�ev�uȹ��ph�e�Ƌ.��/�aVW��*mu=�:�]�t�'�7��z�A���FÙ�kW�ܡ��5v�rZ��żGd�jtB�6V� Zq+H1�dC�	�Q�H\]��[�m_�p1��7�y4�#�ɜ������PK�b�̋��P�J�o���pu�C]���J�\�{��0�,��Wk�0����0d��*S~��oS��^����l!�㝁���l�T0V	��?X���w�B�Me�,_���@z����3�f�5]w�z����h��vc���n����M�%�84W�1��q�����r��q�ba|D����Ձ���l��k+9u��u�幭O۷��wr�Z�p��.�L�o�GE1¬����l:����=��s1�$��r�g���S���a�}+�>��<��a��H�j��7��0b��ki��P C�
��x2�t ����x�Q���7<�#GA�,92��WS�}\�c�}�RK�<:�Pۈ�A�Kd�����"��e:�c	��T��5�ʡs:M���L�\ID@��ٙ��DwL��1��9��O[���F���aS�Z��ۥf�1/���|ꬺպuJ9�Ӑ��ّ2�z��)�R�o,[&��Ucڡ�h	����=�M�;��sr�S@Y�k�U�f�I`�l��p�PT7J�� b[FG3^pj>}�����6}�Q�]��G�1r}�f^�`Q턢��#d��8_�I
(	�����U\)�Og|�\���P靥�޻O�����&r�@aQ�@�.���<K�G�s��K��h����f�̙"�uO<�C�ں�c]\(&�ƌ�x��^<�f(B�0 A��%�Q'���꾧&��m2�I���T)�Pq���i�j�7z:ttt2�i��ה(T�5���yv�Y�:�Xn���o����^Ґ��l�0��\s���ط0ƺ�^�dΑS��v�_�����_n"��e�a�M��2�l,�un���	5��5�ځi�Gb�Q�Φ+5���ZWt��� ��+	��Z��#��63/j���h�~�tI�F�Pv^M���8o��UoV�c�җN	��l5w�[����@^i�C�T��g�V�|F�µ͏�H!�o�.ŏ|�y�_Uo�w3xiMO2��G�㱘\�WX�����'v�K ����A���5ύ��h`���Tn���vu��{�hL�����_�w���ry��B�{�K�;K�S`c7�իk�q�b]���Q�{E���&u�te#1J�%�9�Y�z�$�6[}��(���Ƕ�CQ�ʝ�vA���x��;�G�U9����t�尤���ͼ�5�ڞ)*��8���NI*ѻu��!±T�_�\\Em �%S��+��#S�.	�R�0@{��g5e��'�KY��\0���T�`U��<Y�^L�B�v�t����S�a���j�v�lh�qB��b�E\ΊF�3<�:c�K TvI	kd�A��d�J�,��w�\g�z�oO}1Q�ģeP¨�'�2��:R+GJ���J���B=C��)G�wZ�g�i>X�[��s����{�ñ1��"4I<J�D�-Q��@]m��u�9Jk��*ʉ�n�כX�M].��>�އ�γP��aQtH�UF�B�pO"��R�K������J��Cq���p���pu;cS3#�>Y��vmC�B�� �C��|�Ri��4�L�$~��S]�Ū�Ʒ8T;��{K�N�Vy�^����/z���w���z,�+%=+��\��IvEPq�$��%�S(GI�l�q���HF�s.i�.�j�C�oؓb�K:p�\�ڴ�E�T.7"X�w$�d�d��$�����A�u�| ��u���W�Q�Yj�:����ZA`���`��a?*ZJ���ښ�{Si�wPԋ��&iZ.V�<�����g�1��:^�}N����	��0�̎�@ܱ]Jݶ[Ɗ�dF��I\�f��f�X���.�Hu��V��;F�k9�Y5x�G.t-w(cPL�JGwb����Ak��yS����ذ��r=��s�<5�Ҡ��a]Ծي���4;�^��ب:u��X�ٱ:��)�1���	h���d��G[J�����Tp�Ĉ���odj�����V%[�o}ٴm�tks^�!n��[t7!`U�e�܏mTk2��� N1X�4rZ��')*��H�#���,Rw$�&�Q^�|�ե�([�*Ȼ婈b�*�C�ƌ�n�j�M�'�G�(�ݝhuҽ��%ՙui���7Z!X�υ��R���γL������%)_;p��D���d,��˳C�ХtN��W��B�cM�n#�a}�cK5ԣ6�����=ۈ�5g��Q��}FWv�sH~�2�p��dv��űvF�PLf.�\���F�]�x,���HTys�rVC��-"v=��JѫkA\�Zw�Rq �T�p䷝[{
�
�խ���9.N�&ǭe/'^�/�'!��2����� �v����c�3S���lkw�d�)�����%YF���� ��$�C�}ږq��u�d����AЇ��Q#�a窝w�QU3*^�S" }��e�ġ�B� Mv[θ�a�s�-7E)Fލ��}
�S�5�V�o�Վ +�Ұ�GE�x��
.��z���������s+�&��0�q��5Tyί-��#5��^�{$�d��Vj��W�j�_^i�ึ=�����J�tl�0��ۨ(���}�SW^�{��1K㸒�c�>�Fn:�F/���G��-ܩ�M�Ee�����m�Ǒ���N
)<�b�:.[ ʋ0֚�U)�ۊ��
ڴ:,7ت��xVh�(()��T�4�u�G�5Ϩ��u�N:�{×h��PEёI�LCd}w}��"�y³��'��m	V�M���pD	GC�vĹMO�e�,��g+Ɂ!Ӻ�ӹ�X�@�wt���%r���Y�^4!�:�a�|o��v�R-7s�~�l�,Ǻo��t���!�o��H#g��ɽz&`b�d�=ܠ�wboq)QU����d�nn�8����ۖ��Tv�ʈ��h�G"�G�0o:ӵEk��\�I(9u���E�(O<�>��*�l��������z�o[��G�=�u�H���F>gq���'\e-���.bf�x ���+�5g;�sp�2��]�����:�J"b�yYn�Z�|���$�B�͔�`���>1`tfW�}`��.�Ÿ'X=׸�4�Лnb������rk#(Z|�V̷Ǭ䵥�R��o�<��"����g�Np�
�󣿮���y�}��S5TY,�bce��VF5�YecF0Ue�5f65��I$VNY5�A���eYQYaa9��T�Y�TRՙfVa�a�eVbTCe�e�EH�`VYc�fNf1�VY.U��Y&V呐Na���Y�f�aY�15d�eU��8M&S1Y�YFE2FNa�UYd�VXUQ1Y�0NYVf�c��9fY�E�fX�T�ed��DVM�TE6aVaMPQ&A�VfNF0V6a�A�E��Q0U9�e�e�AQ�a�fYTfUD�LTf8Y�Vc�Yfc�EUda9Q�Q�d��faDfdY�D�S14daQdӑUEL��QS�&YU�Y��dQf`Ew�u}Ee���#�X�;%R�ov��U�L�t���v�\���⼰�"�!\]˙N��5�/�5�B��n����$CB�inʿ�m����9�T�M�I�������]�%a������[��~�]D��Ja�y8� �� eB��w�G+���Fj{V�C�rW�+oa�;�#F�Q|gM�h���J�C�MY��'����_��ehX�Z�X+�ݺ��s��7�S٫-B,f4�� �Qn�qCO@�Q�N�7�ǔ�v�8C�ۑ��w	
y?B�.~/����6��C���Z�ᄹ���d�x�W�,u�3�����"��
L��W|n�5˼�w\�]X;���F�*�͖���O'0m�l�����/Ӳ��.Le����;��5j�G8	S��&{_Lb����K�F����sꋨ/��$[9��K�aeg>�+�*�q���R���@R���hN�p�X�Rx��a�%T��j��3ڥDӹ�Oj�=k
���-�܇�C�1���w
��Z.���-�Wد}V�ք�V3���ע�p|�K$E�^�U�ԭcp��YT<�qA�޹�&%n��\e�l�^�8���c6���5����+�_	�a�mr&���&�r��{�˨�pc��-�tJ��z���M�7����t�u0b�O�蝍�֬&��j�b��f��8��N�Af���냰t�龲��Q#k�̗:"
M���OP�I�Q��iD�+
��z�+�8�X��������]2o7vS��Z�N��K���K'&Phߦ
1�j���S�csS�ƵΫR���)�����į(���b��\�7�0�]���,*��;�`��uL�I�F��[�*���_U��R�Xtv��k��t��1>�'��S���/&7�kn�1m�I5����HW;�Hl�C���'��,1�dC�	��zξʃy=x�������s*�����＋b�]��w;�k�d\E@��V�|���@�[���ٺOy�g)v�1n#���+��X>#e�'��T��S~�9�#S��^����f�o�#�P���R��X�m"��RB(<鱈/N���T�^����d5:"�S��0*��c�3r���}�r�껲[��x�,`�ɏ�VZ�k��Һ\�zW�
�W�VV�ȘR�4S�ʾƷr��庌�}�~�K�����8�vK�S,�⾣PB0̶Nb$0��n�6�p��b��iЁ��*���ûY�X�٫�wWJ��N9�e[*�(�W�b|t�����+�4+w6�Y+y����ٖ��M5��o�7ՊE��u\0�/&^J��G^�3J��Ӭ�E.ge�5�v��Nﺦ^�h,et|#�I�[¤t)q��)��5P���5Mt�8ܑc<�M3q'h��J�ls���ԯsT=Գ�ė0�AT(�%�N��zPe:�T�ެ�
���xԡRbطI,��Z��n&v��I�b*TLw;�Yf��R/����Q��w�:����#��\����"Y��f�3<�TȎ锁zFq�zǔw��m):�ͽN:x����*�?6*�T&6�U5��B��<7邃��Tª��-NR{!���1�
��x�7:���0l���0�ds���<K�^=(#�r�zD>쫭d*��:s�M�ӿ|���u;�q568d<w|/R�b�B�0 F�Y7'���<�=/���Z����
�=�d�z�9�I�ގ�
]��ZE��6�� �
 E�W�ҧۋrg>��&�/��#/�ؐ�s��z�&����0�:��<�M�a�9�&��)��dU�[�,m�C��;$1��p��2�l.���w�nX��R�yUD���c5�T|���0�}���\6�W]�%YnM_3n�@q����_b�f�dʴSO!plo�6m5wG`.�ޥu� �V��^��Œ����jG9pl�=�X�n��U<��1e�I�s���@��&�Ls;�
̜Eg#�i+vy�Eu�1p�N��H�r���X���c��'�ˌW{���75]�MA�,p�ͥ��{�4���J�Fϴ�0�Q�R�Rc���xP�=:,E����)�-ՙ�C��Z��qK Bu=��s�oݝP�7(��rNi��8*���oVIG.�8_X����{�c�Ȯ�&dX����ǩ,>���X�V��s{iZ���J��K
��lbxT^���!ˋ��ʧg@L�8Ա��Q&��+�h�O�s���l�����wh��L��ո���d�Y�B�&j;�0󥧖BJ�)�ͽ����y�1v��;��
�Y(��K�)%��������Dw�O��<��mfSn����I��S�[}5R_R�*�eL�l�%�~��
��.d%2�#-�_>r�S���[ւ���Ii��I�r6-��q��TA�$�%@Yd4�g��Y��·N�K��x�w��td*}o8�}~�b]W�s/���lФ4WP��Zߢ�z�=��f��q�K�E#�ZwbBf�ާ#�*¡E�k�I��jvނ�����>���Z�:Rew������K+m��]@�Y5��z��ЫxKp��k�b���dlE���ƴS�����Н'Sel�4�8���,�}���}����Y�;�9��	��ʳm�!v�b.���'��$�15V�F�㜐�A���y=cP9�3���=ΫL�Ͻ�-�7���zH��ն�� ��F���%�@�7��_�p�EЮ�/�h믻X�%Q��2�B�"��np�W>�t���8."NCJ�񸇑,S�$�9!a��<"IB���2�#�l:w�qd�S���*=yzY$4g��P{���=`oW�Һ�W�IC�;9�s�7*����S��دː��|'��\h>zo����vQ��h�� (� e+��q�GGX�zX�[�__{�}���i3K�k<ͨ�r+g,��,h5��+VEǃ����@D�VT12�P�éuw�������V�3��e��[���*'f-�E��Q��&��)�FN�7�NVˁJ�_.���R48E*3$�Te�d��ޱ���SÂ�FT����:�o�k+ �jo2�j�d���0�v=tlU�f�]��b债�@OX�ȸ[\Las啖���5��/%�ԍ^�4����&j;.���y���j{ T��7���3����/%l9&뎸��k�9�Q��]怠�љ1)��7w�*\P��&���BpG��P��J��uܻ�GZ�zw��0s�ӊ�$e��g�"�L��rZ5ĵW�����ӗ��o�tY�"Q���Ys��\�ȩ���R�j��,�k�6����/�"�N�НF��jO�:&��Q��[��)S>;-�p�f�݉�J
�h�ih����u���NB�-�rGS�#��t�Gm[iF��p���N@h�*���R�M��(=��C����t�={.d�X�ǖ���A��,H�/�H w�q �@@�I�^�v��$��a���O���l�Y�
��������g�j�����پ�,T*�yId�����Mo�ja=��X�i���
�o�Bmr�A���9%ي�ٿ<��J����$"J,*تc�;j T��Y�P6�n����	�f���^�7���@uHvAa���r�S��j����zT�ut��a�O_f�};���q�X�1��+��$5l0��DN%i�6�̈b��0���W6�oV���rh�d�#.��5�Y�t�o�	x��"���ZO9#T��.2�fRnY7�x�飮��C��p�γ��eA~9Q2�Oy��+M
2%`��˅����JWƧwA�I��v��J�&����-YZr6Q�j\�X*M����ɖ�[��.m6t!��4G�X�:�,Z�R^h�i
��H����ժ�� �
R_.j+���,��y�ës�"6_|�I�e�Գ���^���BN���Nso'Um�H�[P�p�)��P_�^�U�������.��D7�p��*�������rA��uq+:��'���＃�tF����ˏ��L/�ڟ:���\�ڷ�N�jX*lsN�F\b������,.�
�L��&��3���޼�^����ԃ�=�O�dt3O2n��w��ƦX�5�Oe�^��0-�3�D�V�9����U2=��:�N�h���:UO��F�loVW3(�F6,�[t֚䰑��t-�z"�E:��U��p�.��f�� ���S�F,{�{OVjo%E��	8Wh!q6'�x�E��I���2#�:� o��2����W�����Υn��3Z�Ye����|*��BcjQ�8������(;S!l*�G+g�p�Pʘ���(�n%�ݻ�|�c��r�0�� C�:�G�g�l�+ke���0E�m#|Oz(s�æ�ښ<5���Z	c���U$B��52��}�-�n����V���<3M�܊�G�D��j���.���Xax)׼�]��d�vɠ�e�W#/�rY��ڻ��̚&��#h��87W.T��CY��[���Y��K-$�
Q2�O�̍l�7�i�i��uM;��yJ�TY
`@�@�d���&v5��}��xf���R���Z�Xx���c9����K���'�tƻ������:Ȑ���JNݮ�=�<zKg��U�o	l����i�P��0�:��"���������lek5�Kx�o(���`���u�����҆��ٰ��3J;��&��b���)B�k͠��gQ��.a�T�X�^wTŬ���Hb�wΘ�ff����``�gp��e�o9�9�w�OvD�~�P�Rsh�9�G���/вNq�i���/.&�C�oJ�]�uMj�Wmui�]�\C<0:�N�5��!>�o���=�?��8��p�]�5.�q���\9o7^��^���d;3�^�Xq�]X�L��q��"��F��kU��,m��MI�N�ߧ��D����2�K���xE�ϡ�n�ܩS�� &V��j��麷`����O)��o6��w�`��Ms;EƓNtGX�P*#�J,�*�f�;�)�r���]�Y-��=��o��%�|w2�����#���҅��ݫf>]��P}�;�OqG
�П|X��y����ϟ[�uC�grGucŲ�.GJ�u���ײP��Z(�� D�K��|;�r����A�dSW@��]rY�����:7,.Q��ŪV"��Ƭ��#�b�MN�D����@OX� �vI	:,h�C$��� Y�p��'P�z��v��҅ƹ�C
�&���Z���ϟ��(\4m�H��[�<H�6���!�Z}�VC��l\>�mؘ�"4O��T 5�\�8�Ԫ��k_r����J�]�xy����������ō^ʯ*�_�#sf�(�z9ҿ������Z�����LL%Qu�X�T���9�cV���	�̠�˳j!�!sLu��&ᆳ��Q5�bCV$	JH�dCx�����1�ξA�}�i����5�K���ݜ���I��y{P<GG9(��B:MDCf7�PF��C�P�{��6��M���F�#U"NF�u��Ȗ*!ܒy���s�&�2�����Y��)b�ìŽ����Lr(s�@�����4�u@�fd���x�V�]�|�O5�J%�[���"CΛy,k:��$��P� Rq(Q��W5㲎Y�߱���4�/��|-nְ�I	�ьb���'�gL�U��T}B�e�;�ea/��o�0:*�&�})�-iM�l��7L�wéY�Wy�@�W�*4z��0(�}�nVT"z.�Sv��܀�
f���n����$p'21����˨�x{"�3j-�����X�j5S�Ebjȿa3���8�'1,���2w�����w�l��wJ������D����tS������ٽZJ��<��r��Ȝ��c3�?>]�֧��jݻW-Q;�򪌥U�d���{�.�n��N��+)]���"8�T^;���xn����mѱV�-tJǡ���0:�l���tW +U������V4 x���j9�N���f+Nz�Tm�n��xO
�b�Y�]s���y}�]N��=�s���i!��6刘R��`�Kg��Bu�Xꉪ<``0���oT2�/n�����H1��S��@�Q+Aa�C�!պ���V���w$u���C�J]++SǼ�J�����* B�$G#Q꣺U"z�A�y���Gd�/�e�C�]�U�NX�D��g�>��Ҵ�#UI�	yId@��A����êgQZv sShд6�һr{��ő��享]c/`ZkF�B�=����@[�	��?/� ����� ���� �����
�
�+�TA_
��
�+�TA_� �����
�D��* ��TA\Q{TA_삢
��W� ����D�* ��AQ|AQ�b��L���N��׿ � ����{ϻ �������>��U@TT��"*�$�l��TI(IP�
�*щ����d�
���{V�J�-3F��m����,
,c3m�fF�j��լef����[Z�X}*�姝�S5km-��4H1�Y�b�CFj٘�Q�l���e6b�[VJ�2&�V�lյ�2u]6�������h"�Z练�ўkˠ���z�f�x/��N�ڵ7vnU�K��m�����{V�Q�l���������U��q�k��w�N�e�\�]h���7�k���E���b�����6���"�{���8�^{6��zӏV�RZՐY�| ��ݼ �^��@P =�@  }� z�(��  p��C�_v׼�{�ڶʽ�k�=u�ݽ���G�q�.��n���j&�jٱ� �g������[��ݝ�j��������n���vt��˯y�2k�k�o^6jh����W��ݎ��:On���{z�\�1�ڥ�|  �|�+kg�����;�������ʛvwN�����/e�T<�����-���7oFU@ƻ Zå�5m�-4�-��� ��m�6�k� �N�ph.�R��p��]u�(�4��2Գ[a  	�@2�u`�Z�
B�F}S�
{�\ �@)����*-���2���מ���)պpn\�Ggq��� ��Wקop�(����M�ր���6٩�Ռ|�wϮ��b�5�t���Lr��A�т��y� 9���m�U�Vm�ُ�y�yr���.��]��`n��];����@m,)G3h�    �lU)J0FA�L�4#)�)RU0� 24ɉ� ��b%JT` � ���h�A���%*J0�40�M40	���T����"a10 !�&`I���4���a�d���O"�j~�%?;�~"�G��'����z�cI#�J�G��J+R>������tL?L	 B��%	4��HO�HB����@��7�?����48�gI"����H���$B@�$�C �'i !��~<���8�h���߿�� B<t\���E8�s_��?�?C��((��=�_��O�� A�۹�������ҫ�%�Ʉ�P�2�����4-VGN�ܰhm'N�<h$~��Ѐ�ƭ��F�[ z��f����sm�H5H3�E�93"zh,����N��'کe2�WA�Y,�i�zղD����m*�ꕻHK85^|�k`�Iˊm�8��6X���m��Kշ����ǻ�R�iT��M#Lm��hd�R��v�:�2L�kfE�>�b�l�t+iʰ�Fq�s*���W{��h�Y��K,l#v���n$�07Gw'S�4�Y�A �-O��6�٫��uR[�C�z���X��l�Ut�*�\��fHti�2Y�:�T�Ig�ea����"�n�if7,���LʔE��l�£�m\�٦�t^S.�Q�~�#xPgmV�mݫ��8 MZ9�Q*���!���nX�����낒���t�N�H��.���Q�k)�^ �5�@%�:������� �G�:۬�P�pe"�yW�t�n���+�A
ȉ,
��mF�6ۦ6���E����`:�f3n�79��8[��V��Xїa�.SUH)��YR�sN�5@��P�q���l�M��9DX5�/�����3r��$����)��n�6m�Z��H���h�zF2�LS^��־�ՇG5��+f�v/�w5�b���?j���I��p6U��xظv�j7�Z*�a����MT��!`�Șq^Q�����qQ��R��V���C��Mw3+^�m�<ˎ���ǎY�cY��T�݈-��qҺ�>5�0�v�3\p9��!j���̫"��C�m�dʂ�9�6�%�o5�@ӣ�$
�.����*�֌gR
�* 5��Ŗm�6����򶆋d՝�n�J�gC�cl=�҃7XG r�1�7�7�s�����S2�PEG�e'G\E�
n%ø��F�A3$f��(���.�;Zb�t��M]��=שAA�$�h���%�j��i/���f�
�YW��yP����Q��O].Y���oh��1X�`׫�k1�⸜Oh"L��D���b�1���k�R��7�Y�y��Gu��-Ϧ�DL�q��kf@�ݔhj.e���J�3	��͠��x4Deb%HݙD[�$F�ѡ�e�-@VPf��M|v��K�7O`C��K�i��-�.�o��[p��p %m�jX���i�����Wk7�+�F§��LjEJ�0M�7�]���u�[���x�y�
sdWE�%ƶTW��w����5$�rQm�P�	LB#�$kw7�	@��S8#Y���LwRf,.�:֞��sf]I�Kǲ���`ͽ�d�@XA1�鹺d���:��3��,"�����ǥ�p�(f��)����Z9oGX��l^��� GI�9�DQص���1���g�R;�d�H����!÷B���BYF?���,g)gj�ڵ%b�7M��u{��=7Eԗ��V6n��aRV^��F�42�\x���V��q���J��!�-ي,�s[��ѦK�{��M#����Xb5��'kˊ�]i�b�{��a{sr�j�(���OI�ni�Q��[۫��� MFfX7@s�3*�]d�Xu�iֵ��[ ؙ���a뙚l����!v��f�ͨ�D�͉�3EAEa{�Tf�V�١�jOD��$��R!��lf���$.'0���o>$ܕljKr�XQf��m2�Tڗv�Ԑc�slh�w37HCQ̖ݳ�MX������"�q��p
�!+j��(ږ�M�i�kq�PJCCڹ0Ԭ����dq`ɖ��y�*n�����P�z�`�+&
r�Һ�!�Iv������.���T�l�̶-�&3�BC[o���h�3Ekq�v��(�#��N��` (���D�hѳ
)ݠ��d�uh��X4p$�ӣala �;w�]�jĔA�.b�yZu�x�GrU��ܕ�\�r����́�2����MI.���&J ���y�f5C
��Oq,wQ�舝��f��vV�ZL�{QR��P��̵�[�X���s+���wrhz5&�-%lՂ%D��)ܿ���wc>�X����1��j�����#��5@�m<�V�{ V,��Z*�:jSt�o.:&�嬂�	��X��aE�]�t�vL�ҙ�R�����R�2�Z�T������5Q�x.
*_��LU�e��$�r�`��
���=�uz����Z�4�)���~PV�rlݘ�t�i����`[����hz5-�bVw*^Yn��N�x���b��u����U��>W����#q��(U�lZ��
1d��P�F����G/Uh��L"�ar飀��D6h�p����4^N���i�svT_Z��^9��KM�eC��0!��Mz�e������J:el��D�V������P�ݢ��L��)�۰�<��VP���2�P�]�;ۄ��,�wm��*�#�6������9,� *܇Nn'q�
��j<�N��h\�ͳ(����H�M�*k/L��(��vc���4��:&F��)Ekl���KZ�i�X2�*5���3@�C幔A!�h���MͳD[׬�EO���PŃD�i'�̵�F�T�	�j�v�]l��_Ʊ����앭��[݁Yx�+�,и(z���2+�8ko&[�F�ߝKVL�dP3h��X(n��/P�X8�t���Y�کcohպ��(���Qԑ�$+ !���-"��ݧ�u�0�b�J�
[��9N8ٶvf⡓^�)	gf�Wx�$Zi%Ym�V�b���su����Ml����B�!���.A�k�7v�2Be��c�3T�Ԩ��0����u�=g��6���v�%�0��{����xy��RT:�L�Xf�Q7B�t��G�G`0��' ����4\d���h�A4��ץb�7eWl�x���Y����ɔu=*�srѧ���uUa�)U���hIX��o�	��R����ss30�_P��0lO�J���C.�͏"�5e,yNӫ�q��/V� ���9R6��Xw`��V֥e�	(V���Y �b��(M�g\��VQ�Vɬƞ)#��`%f��d��)� �df���i@ ����ވ���WtQĪbݱ��X�.�fr��EeL��Q��Q�rH�P5��j�w(Rv32�����:�7M�;Ra-Q�0�ɉY[����5V�G��� �M��he-b^P/N]�[yF��"pGh�m����V2nD��v��4�{�&]�;yR�/d	i`��Ì���l8�9�ֵ���bb���V��-[�4.T]�.ь͓s����A<�5V#*J���L��<sx$ܬ
^�YV���9�	��N�F�$w\m���E�sn�J�4�[C)��N͈+~�F՗a�
K^Ǯ�Á�@�Xݸ��2� �@����H�e��&r�S��Ѝ��3�ja���{�E �m'��Kl[�(�Q8�9MMܶ2�	R�(�Lm�y#� !w�]D��*[:��/f�,	2,��.}w���5d=��53�f�d��Q&��3H�Y �)��D&��g5�k��m'�-���k�ե�Ě�o2�'�/NU�������[#�ȕ���p'qG�9H��&EI�hUu�[�}4H�$��OkqƎ�\u*�4�+�u�6Q���퓵��t��Ւ�ئ�ܩC~Y�DԶ�O�B3�1T���q �VTLfm�n��
:�3H<�n:�C�ݨZ9���o>����W ��9���Rˎ�)h�m��kw��#٢��B�b�	j�P�JT۷��:���9@�uf��x�ҩ�ǵhh���l���u�۶���j�.i*��C9��D�{j���iTTە0'de�M�`����a��n�@�0�(�f80V���$�d�m拦����^P�3"����C�qJ8hĹ�E(���8�:�vգWB�C�$B�<͕ec �CSo�w�r��3nh��h�ڃJee�MǇ4 ��i)l�ĦZr�vK�gU8Rp�:�MPǴmb�P(�,8��4��n�K�%k�J[�ںH�7QR,XV}o!����ض�4���P��cw�!�`�e��0r��D��N�~�O�}��p~���p��"}G�π:��>��_#�G�������~e�)��HHw��˻��z�d��x�|ɧ<�<�쭦ۮC�.���*��p����:�NV�"�t����L��<�9��*	i�����ħ��L|�ё8+�K��ĉ4��,�ܮ����<�e@�T��cl,�� 5.u&Q�;��*�k;HKf�\U8�:9�*�\�s!��|gY�fTU����S��\��&*	}p �Ѥ��GF� 8�R�V�E�8�ԝY�Wݶ��E��ꄒy�s�_fn�W�*}ǩ ��K�˖��r4eBg5�p��*�ӎ��ל�kS������+�qũ�E���y�2�]����ӥ�S:���[6�fލ��>�^,lZ�W�*ž�6cb��-�z�6����	/+�����[��M]���Ie�|݈�\��Cr\�dT�Ǌ�¥�{J���\�(M+uk2����]Q��v2EBM�xRS�ز^�fuu�&�]�T�Zľ��8i޺؅˂;��b$�Hv��r��3l�_���p�E.��,�1O]9� Zb���܂�bW%[��ޮ����4ƃ��}5�w*�u�����+;p��k仔;t 6�r���p�]�m�g>��q��K6�gD�}%���"_I\�	4���K�2���V���]^ЇF�s���[�λ4��:[Cn��y(�R�H R����ɲj ���W.��;q�H��8���"��y�	/kl��p3!�w}3s��Ԡ��nŃ��)c�b�Xl)-��n;�9xr>k:�9�gN��ܩ���ܺL��D�f�A2�r�dE�5�u��K%�������8 w�eeLD|E9�̥�H<��v��(Kw1���Sw���x�r�$�T���)�ٕ{�4�'��ۆ�ޔ0�U�o@�\%9β�jGˬ��3n�|��{XN�E�k���Z�]�ڏH�JKX'hb��.�Ttۊ6�$0urgD�u�;�Ot��7ͭ�|ݪSlQ�m*r�2���� (����L�VܺX�R����K(fN�`�/�7�5x�r�W!��h�}�,�@�J����m;.���[y� +�;�\h�CrRkzb�#G�۩Z�z
�-Jj��ؓ2��S�7	��Z�z�v��B���%�:ʏ�:���a�{&���{!�t61u.��W/�Rc&���Sz1>�@[k��gNԏ$R[��L���.��ɱ2��dWg ���k�M͚�Ut�<�Is��@t��sZ�u�j�K�!������]gi�.�7��\���OfAԫB
[�6�ʺKt摯~2�VSۡ�NA�TVq�wT�\��-�v��u�6ZT�Z;�:�;XmSGvGXr�'2����Ŗ��̦J�I1򛜫 qa����.�e��H�c~��o��Vho΋C���Ɉ[V���Պ��646[���6:j�[wn"ӓ��/�}�+����G4��q�׷RnA�A�c4q�Q��F�+t�U��d���f�V)o2h��n�����K�.��iBn�Kh���PӼ��}>1̠r��Mt��KB�)�Rsɉ�|]���0�fe�i���b����.-;�4(�}]�ӑ�يKo�4��s^�����N_=ڜ+s�ul�R���tf�t��{�����K���Y~CQs>�X�t���	���h�l�Eqv�,�1��c���V��âGxH��t,s�;�g.e�n�AC��E=j���-��6�2�N�M�6Ы���O�+�^	�\��V+;5�H�B�����.�8'D,�\�M6��m^J*�MM8�r��R[A��	X�^�x]��9GQ���U,R�C��e��RD-��`�r���^�3��hoB��:�n�f!���d��%#�7��V����ǒ��ȝ�ܻtV�Jfd��US�GE\�;.���Z%Z}�/�v�WRV_Φut�N�#��r��K��v�|BE���.��bB .�T�vn�oe�2���:U�wK30�$i��}�/ީB�]vM���Ǵ���3�]�f	VD�ю����ڡ���ws��H�K�f=N �����<ᳱ�2���t�\�]du�<�����	�N<�Shl�(>�+����[w��Y%*=c �z���&�.�1II:�q����f �*^�%��5��|��*?�!y�P��6��8�N�C��[76���N+/�-S�z�u����r�x�!f��B�>Eҭ��t�W���[�[�	�K���룉��@�+��{	ۧXȕݞ��Oy�(&��b�3iD��1��g��6�N5�F$-���R�p�zD;�헔��)R�_V])�Hn�>8�mܛ�p<ݬϣy�.s"i�b<U7���\��O���-�+�AЀ�� 5�a8c]�� �.Y�5�%�y�$��� �7.�3�]�7�q܁0��}�3�5�^�N���B���G.�Xp9��VM�`����q�~�����2�N�6�m'�7��e�=�.�H,��%�J�v;$(�]H9��1��Us�چ�w�C)���nг:�-���ҭ֧ݧA!�U�븝��}&���"=���l诬p�l[M��p�:q�Xp�
ܸPt��D���[*�a�5�0���F�Xy����ͨgC�\`�����[p1�^�sY�O�b-uk��N�iv_n��W��M:��̺�p$��t*)�o�2��k��Z��h�^���.��� ���;�`�����r1oX Y�eoX4'8�� �ݽ�u����GOq�T�S�ϑ�E���eZ����)���۾yƕ�jc�ڢ3�לЂ����D�X�<��,޹-ix����4���W%*S�e�/ml�Zz����_NPo�+u��R�z��K���K�G�9B�HF�����ǝu�붎de_<켂)Bh���k�i�6�^��*^��t�],�o�����W1l&�K.��fCG0�Yii���>EΔ��(Kw.�y�~��6���R�eh��b�Vxb���哕ҭF�j9��vmg��x�)���c�ϓ�>��@Me&�M���Tz�0oU/���8y��@ۘq�unG2��D�Y�W�"��Z��� �yz2՜���3��鸙�3m��շ�,]���vE��gT�򙥝a���Q`lyu�-O�ëv'�0غ��Q��!M�w�v�5r�����3����ZۛJ��d�����]#{s�=���+	���r�Ν�����r6�ƻ����Î$����R��3`��^,kM�-���n�&��(R��M�j�g)��e�L���I�l�1�(;�/r���{N�=�i�X�͢�FΌ�)���^)H��HKh�o&%��>��Zx�l(�þ��iqCU���Ls[��J�P]m��SN��4k�CӗK��)݉�K�ǧ�w��+��M5�5zp�L��)�+xKS�P�rVXwD.��2G�8;I�����B��V�*Ƹ�,�0�O��߄k�=-��_v[cUu�ڑ9NL�WJ��X箟^�	}��[:��H�XuM|�M�����G�pޫ�ȵjdR�����ڵ�j#p��"<\1��@�-6�81q��#�<O5*��\~��p���oWǒWV3�#��`�v�6��s$�c�o`A�S8;�w(�}V�p]�z�=];(J��oFs�朋`�����{tq�$�7��hfö:�Vt���%���+}B��
�Ѳ��� YVY�38���z�J��j����.��|]z>���IL:�����zw��f��Q(�ga��p�Y�ٗ�+=�ܓ��^�/Y%�N�QsFAd���ۙb$Z��):���<�P�1���v��5۹g��7Gn����WZc�#�]4l�4U�!u�eC.��
P�gWD��h�ߕ[���� �Z@��Ր
�gu�&��r�a3w{�No�F"@��RQ.]�����msèݾ	ʌmpJ󣹊Tr��,<�N-��.l�:áҺV*�ySvgsJ�I$�I$�oo��Cso���(7-���K}��n[�+�U�N¸ۣx$��A�ɛ(������ɷO_G4j�p+����VHD0��dnGǶ^���t:A�Y�![�*�$N�!�mbZX&��M�������|=H�C����?V�px%�pE��s��W9NtE�a��Z\��*B���N�uo,�{��E�31���o��ޔ���Y���B���d�P�V8�$���~��W�W��=�aG��HH��y�g|H$ o��$�N��<0! B�Ό�ς�>���]p�+�%���j_�ԩ!�N�r]��,Qm
S^�ufw�C\L����Q�^�r�F2y���#5C(�Tn^,�������eXʲ���C/�[��
��<.��i���Y{��Ut�x��@�],\�Vӳ���̢]���W�2��O�*0�it���jGe��؜�ߙ#���
Ұ��i�K���x'0)G�N�u����O�mtj��b�%;��TM^1��ə�
p���Ŕ9t�b��&'.��b�3"����(�F�*�*Z*R5yX�n�u0
4��|��ݔ��^�)��z�����u�6�$.:ю���* �c.�E�G2�-����˄�!u���o��F��u�E�^B�K}Kye�b^c��:�N���D�� ;T���mp�V:�^-��*�U����1�K�@v������؝�v��Fm������r	�QS^�.�� Vb�܅��e=[t+�P�|�m$9��2��p�	5����F��\k�T����:sי|����H�N[��TW�z�'rĲF,(lT����s�b2Vd_i�������|E+E�w$�FbJ�M�U�G`��@x�v	�ӗ���Xk^�W򶋅�P]v��uR5hE3u:���Y�f�m��[�P}b�`���Q���H-���h#2�H�A�7�c����1��3��� �e��K̐�=��k'[y��[��جD�_ ��:5Z�e������}�:+�Y�j¶���([@'`�������]��I�"��ydG�Z��{trT����'գS�VR��y�$�V���~�l:��҆�
�aC�X�X�,	�pv;1$������gm���N��ss��ܣc���S�y��t���RC	�i}6��K/��csR�v�!�5��8m����X�"�7D5��8�/Ah%K��QT�p��pmЭ�0�/$k^�ZY;�؊yw|����
b�Ll�-8���2��Z�!�H��[��]�	b�M��T]r��]nK������hMP�O\@nS��� QsD\vs'q�G�2��4)n]���;	H .��ۙ6
���YJ�֢�WR���ثΎ���,C� �E�b[�2l����R
j�WC�6e�vL�[��R�����C/2�K~β��$�%�-����ʁM[�EЊ��4T{oBeJ�Ͳ��%lcs��s:�tk'N"�h��Z�#�e���|���k������>��mT�[R�=�)5��S��b����뷝�_S�Bevu�RVl�Q$�f��S�=��V�fPF��4�9N�3���U�r�4)+b�{��wP���n���ؠ\�ۖ6��:)dO�Vm�RWA�Lu��=��N��]�m����R�f���<�X�<o	���:��i������^�V� j�k��=y���tW��ՇyVb,�ɓ�A�m�/'"��
�{{��[��ͽ�\�R�2���ǹ�Vt��_�h�� Ǘô�S��vN�M>j����g�Q4���X��LI�WX��
�Eb�v�u^�	��Ly(��������Ө��iWn�Љ�ȁ*�W`\.����20�[�wIج�U�9"��fV4�e�J�'G�����A50�Yp����86&�]���� ;7Z¡ݙX�!�(WU���h��#��C�GG��.����R�s�4|�d�Qr,\�K�9��(Q����K��|��F����j+5�dF*��mwe9Yf�[�0��&^��tN�5�p�+�wG�|�p��dx�HЈ;0V�'(18l�}��m��n3�pjkj�y[z�`�F�L�Ի�`��*��Ne��;�O8�ZYk)�m8v�af�]�z��Oa���$��2��B� �㊝���.�"e�k����˧35#��*_L��1j��,+�6�,���6*���ݾ��#�hGIP�v:��pc[�g: ;���
�t�iFٶ����ǝjXf������Px�A]s7!v�e!�.T\�LK�hr窞[�|| G�JT,�"��Xh2��w��۔�� l��(�
e<lp��q����U�I,TIM�V��u�w��2��q}bu4R�`�WY�^ɪ�-�i����Lӥ}QCo���:���6r��Mv�WJr�V�q�����]0o -�)V��sC�b헶D���Y����}�)Ml��̒��;�v+�ƬܽkI�M����R�����m��E�K�F�Ef���7� 犘f.�q[�úI`�����_`Tj^6qЃd�iw
xg���;��:�.ۘ\�/)�	9QY��Ks��j�s�_� R�&�*�[�l9),C�&��L> c����wDB6�,�U��}a��u�+���|PKA�"�t�\V����ɻl.��aں��.E\��L���1���4�]����~��֘� 4�Wf�z�\MX�xJ7�����.��5��،G]-��3C�dS%�=X�Ž��p*O��26�h�(s��'׹�Wer�[!So�WS	���ӣ7 #��sh�:3��h���-��S�)龺���8��ԭK�Pwoj��h����Q��fJ���ybW��능ݺ�-��B�F�AZ�#��Q������G(U�N��8�e�\���t�7G2��Yh��9�ۜM��N:��(L7��$�F���[OzZ�eei���p�uc������S����E2<��).���/v��Ee��r��f��+V��׍��ւp��}*k_Z��FM�}ղ�Ĩv�c豣,�uzr��F�uk�ɯ7�pq�~A�ct�x����R�.�HbCZW{���� �-Iҿ�r*Ȭ�i\��^rm��U�e�d����X,��옷1�#�$��fY,�\�F`�����-����7�AZ��r�Z�m�^�N���L�	����	�,��W2p��� Vj�i
��G~�ė/Wt,�@�Qb�
=KN)v͉Xr�]h-
�hG�ou+p۫R�y
܄\�Q��̔��~�f��C�G�9����&;LW���7�r^�-%Q�`��B۬��V����>v��b���յg���L�S��*�=ɉ���2��:][�FcMA�q)�o��6��.�b�z52����5;%!)*�ګ2��A��ڕ*�{>���d��J�.Yݙp+�6����M�Nh�O5�Z��-%w�Q��7�;�.Ҙ��ʴ���%��j6��uR��+9�uڹb�b��ʖC�}|U�eb���%yt[�-�-&hH5�|�d��f����/�wF#�V���L���<�Eu�8u���nپ��y�WРQ{uRS��(�l��=x����E)ڦ��6�0^e��mmI��ԡ7dh�x[�V��r��b�]l�w%ŵ+��g���	�1��*��(e1�	��ݍ,��+_ީr��V��L
K����Y�֭-E�wy8Ց-a�AcΊ�ѡoo#=����}�ˍ�Rhd:��٠�K�kx��/����If!���.��t����l��m%u��'W��v%ON8�F�_V `��,d���[h:��N�����q�U�`�iV3K�1�7��ۤA<�ik��$�5f��e�}c5�U��x̾�- WPu ǭ]�`�ծK ]����Ÿ�e{$��N����:���jˮ/]��W$�V�,�uǗc�7Ƶ=聶�5�{��*�s�U��w9Bٻ�U%�²�DB�u��wN�|�`�9�78x��h�jݮ���N��D�e,������|�"�����0�B���-��CN�OM���V:�G#�W��on_=w��iZ9����QA�I�,x�D*��L�rEK�27У�Mu�{�0X
�Ŧ4t�\�Y����0qu�6�W̸&������7r���:SÄ�,Cw:���*9��k-�dK_N�!
�'����pv��;S�']�8�W���5Zi�,;[Z���w���%e�Z#�Zע�m�2�Y�����T6��F�Y�T�d�O���}�$$�����Y|����۽��������`��p�>[��urVB�� Ơ��?���7��Y�8⠵�Gi�w
�Ý)%��}�f�X+mP�4��v��8�����|�r�8��&Wa;x*㮲��r�	VE�0=�$;�&�z>���O��J%E���9!�ń�xx(�4�����.X�2��9kRI޹����m�)<&������l��ˣrl��3mf�0����jZG:�q��ND�Yy9Yol�:��u��X/\��
�4H7{pl�������[#�k��Q�T��ki�KjJ�^up�)sLҶ��f^��|�>՛ T�"-��Q�u�E1��P�����}*dzֈI��O�(P�irZ%0�s=��U����wun'yX���30a�Qm̓ZF^J"�hRM��T��J,X�m�yX�VK�*#t1c��ù7�/�1���|�؂�:Ҕ�*+v����0�۝�Մ�_;�Xt�lx,�+k{(R��5��h�Y4G���-��G
n=���QL<�c(�<U$�f��a=
 x9"��#I�5�Ԝ�覞ү7�y�>��*���
!�J�KE����*�Z�Y*
�����*���E�P�V(+�SHUeJ��E��B�RT8�dX��iH(�&Z
1�RE����8٭Y1Y.��؍eVA`�6����
�ED���E�
�#mV������c%b�#�,Z�b��@,��,Z��œ�s�?q�v���5�k��LO4L�v��r�P9`���{a�ɴNSP�-O��y$ݏ�G����]\�=��W�?>�2U����7�G�J��|G��-̠�a^����rة�hE1�%g���o��������S�r��ɤ�ux*���7��og�ų����z�p���h^7��2q-���w�ȑ��M�F�#�JoE��Oe�V����H{��[��f���<�S�� �߫2mq�l��	r�~�v�,�={�W�W1��C1�}�����'����e�^�~��wV;'�~��~����#V��������e)�,9.��Al�XΖ�(�+f�������%�d��oE;���ʻ���ΜQ�Il]��K��8��()��N�Ư���F�"ƨ��ڵ-��服�2_�ri'�k0ׇ�;x쬽W�����MKJͱ�g�>��z�"�-��L�>N]*��_����N�Xm�<fɇ�V��h�|�W�7�����DSD��̆+މg��o�<k��c����{+X�..�����*�}��ma���o3�B�)C��d8�"Mh#D��E����cT&��%�.��=&�)-aa�}���E��mN~��.����t��7(c[����0L�FʝS�i��n��\�ue�Hnt���j�V��c_
�{Ngk��"� gZ����y�����$�K6�<�ObvCj0�t�g���WW�,Dk��b��H�	�בQ;/���E=,�5��:�\��Kv_����njpc��i��|&dTŪ	�&s*sY�Nb�۾��jȳ�E\���=�zUܗ;ڽ�;�\]���ҫ�2��K�;�]|�Aat�{���������[���}dΝ�^�Lj�����
����zTQ�]R(9�:qB�_��_Uȡ+Y��SI��l���t��oQ��W��Q�7�+VtO�v1��XR��F��9�G�OZ�e�0��(���>�K�/W	�A<�:og.T]��ԣ�2�v3v���=��(�/�.v]�	��$���^�6v��Vt�\�������Rc��â��Qm�W��\���Fb�{�)AE]Wߖ�F::I#r��e�&�����Dy�Z1<�w�מ���'M5�0E���<5m��9�-�W�*tP�w�(o���B�9H�9t�.ՉI�ϒζ>���v*��
gwA�����X������\�u�BX�9�m�*�m=�طm�',U���b�>�[lw'K������y�+ޑ�3㻙J��YK�ӕ7�l�Ԋ̫���G�ȕ���d��U������e���g"��]5�ķ��^��/���j��a�Q觲\�;��)[�5@�=�@�v6Z�%IA��<��i���Q|MW���B�uR��-po��
�/o��b�@���W�W]�d����)��ņ ��Fj�
��P�<�I�Nz5iw���r,Ĕ�g/Q�$'P�W�^��;.����s��iz�����:E$��E���Ȳ��R�R��p;Mp;f���}y'�'� W�r�iW�(>T��Tv���]��~z�͛+�}�z���g���H�aF� IɌF��nO��z���T�~��^�,$(��ц�FD��x�l.�fe{U�g)�#��*d�mN��S�z��Oz%$���K��s�C#O�]�0�-5qA�6���q� �T���G��i��X>h���B����r�[o6�U�+]�N f)��I�+0�ٍ�%�A�Oc�-<�c��t�e��0��%�Y��W�H�52��1f����Q5���J� �����sy�u\p��r6n�K�R�gA�����4�ס�gR��ñ��w��Z�r�v#Lx�v"=&:�D��o\��k<ˆ���{�	��������#��Z��$=^����c�˝)ӡ�mU�V4TAG
&�f��Dy.>&yDM.�f�.c��,/�օXk��ax�Ɗ�
���3Zk�r��Ǭ�� ���EJ�S���W��ix���{�ot��������K^�v��h�g�ϣ���	Bٰ7����a���}���Ч=\�X~tL
�����q���(K5u,�Y~�1��z�.��><)CXJ��H�B�5�j*~zY�g�� �{�|�}F�yr�.�����˨*�jx�G��a��SWB�ߤia���g~[B�<sv��[ά��S�'�׵RB�=I@�H�cg�AWͪxvE�������Nv̥����Yy}j��R)NQ��{�pw�%����H%�v�w_o�z�J2i.���{��|�$1|��J��K���/2���da�Fg\��cs���K05z�T2&�ȶ�p8�I�V,uf�s�~�^/�q�^�ˏ(�ӂ���A�4�8����ͺ�V���˦�H��+�Ј`��Q&Zmt=�:��sbI��"S@/jdi�XB��:D�("�3�Xם�ά� � �Z d�����h٣�,!Ʃ2*�ع�Wwt-2}n{��8K�.������#��]~�|Ѓ��6�/��N�k6g���6����*+j�\yKl��ѻ6��5���>`�Or�Ts��a�	Za�;�/4��pz�\��̘ī��Uw�Xɘ��i�����I��^�T�j�7��
�%���ɝ#�[l�A�5jr{���G5<�s�f�%�q�*0�����j�;��4�(�H���r�V8xn�/����f���ζ�!��Z; R�=#R�c+�1>祽JqWӀ���f����m/�
�T��s��.v�g��*z��ǅ[+��^�J���IVc5j�S����z��TniϴL��z���Q�S��ԋ�sѪ�"�7���pև�Ν#0�k�>C�3�ʒ����Tu#�F��Uu�i||`�P�Gŉff{QW��q6�yL�b6}a��A�b�+0�CV�p��ޜ�A�^���F���4W�YQB�W�%�8u�Dk���0�KL�* r��
�x��
�B��N�R�خSۣ�v�e׹b��O�����h�<���b୤-���w�:�� �1��6m�ʹZ����4~��V��p�0n�ӏn�k2�,��+�7 S��i��xN\��4��O��7X})<�Z�o���I5'R��@�-Ǩ�Ԥ��;�ә҉;Nsr�/��!z���7ע�Lv���C�� �^��q\�}ɍ��0B� b�|�X���	�%��D{OV��_3g��vK
P�W�V�����C��=]5ᴅ9wI�}.�Vt1^�a�t��PU�b�-:Co�΀u�%C�+U����U���C�Y�1`�< ��,�C���__�=7�����^U�*���zGN��,m|�o�r�5�|��@��;�������^�H����8��hW�dTKS�Ӽ�t���Qt����t���@�_C�R�XD��i���SH�b�q|ߝj����2��?p�
m7X��ed�rnT���$[�Id���غ��)\����D�}��m�棏6����{�%�~󿅝��C��ザ�X��S�G�H���i��
Ý�}�6hѳDQ����x�L� a(!��EV�<R:1�=��o�b�WwNǃ�/��:��Mj5��Qc��\��$=�>@�@�=$��p,�}��<�moU�}�i�� aZ�0�ͥ����r���+�%��Z΍ ������v"='��gn]������}#�*��{U��M��ゅ:���~�ǟ?X��EX6:95���b�`�!�qGHf�i
2%+#,/[\>�ccs���$tӳ^�z�+5�V��/����pU����<�+혦��<�
a���YBV5-{1z�N[�ny�
�O��쿩~O�~�����
�Z�^�*��L�GvA��pZ�"�t�{v��W�^au�Qز�Ґ6������Q�앑���Ǎj�
9e'XL�h��*Z���#�ỳ�QU˴��Z7Sjģ
(݁����u�+:6�Ɂve�*�7� Z�x��6�7�;kyܻ۹;%#}/$�ևFwi���r2Eލ5n�aU���]�V�^�]y�Zg���Ym�Ij�;S�*>�z/r�2]p	�N�MP�2��N��D\��8N�-�]�yQ�&��W��+}y�c�ڦQ�ݙ����u��qT�Z�j��bWY�`�Z��{�ϰ�2��	c;f��_=w}wcYL�nP�22����FN��H�G��c�Q.�|�n����ʻ����zZD[ms��Z��࿉�@֋���.N|Ƴ�sb|b3]:?F�MA�h��w)tkZ
��lN�ol��1���)���|Y;�cHfU��ӂ��c|,�=c������9�?���&�YI�$~��.C��G��.��u�M�rH,C�q�y�M7+!�g�>�Φ���h�vrV�h@���j�<�̵�g�D��L�[�W��8��/�3H����W�pC�h���ذ���Z{��Nŵ�g*�v�7gklڽ.Í:-�qa�|����%�1n�a,���f1�����+�`̛p�����H���)n�y�2]���)�n"/��B{���N�u��N��q2:��Xy��ʟd{{5�d������Y��o�kz����n�HASG�5�r���T�p�Xo*���0H�A9x@�DwJ1���Ҧ�5�kJ�uQ\1hd�#����RQ��%t���j��	>;���nԢ;�oL��f�E3O��
0ޗ�/4��-I���=���
�z۵�=�W[�?�����bTU
��,YYY�"��,�b�@��H��V
DE�Ƞ�Ė8��R,X
���RV�*E"$�VZ��\�
���L����X,�X��6Q@X
)R��UF�R��%1R�`�
(�0X���TTF�2�D�F
V��T��r��2��1�J�*�
�lE���2�[j�UVJ�V[`�%�+8��=�Ѓ��+���l���y�nӐ\
�Z2��>�Y��d����'�J'��m���H��.0�L�," ����a��ON �A�{�b1	վ��z����[\pU�ߜ����/��!��i��Tlp�!L�όu?2�h�(P��S砬�s��xԌ�������"H���P���>#ˁ���㬳6>1�}�B*�S�2��	u��eԂ^��ۺ���a��۫���2�@e1D�L�:GnL�����6F���m�6xjt��oqa�t���ǵq������r����]m�&�Z:����yx�L��`@o/DLi�z�{��]l��c���}1X��=�4A���)�Hq���*$�ͪɫ\���]H����DA4���U���2P�����M��p#�R�<�?R�X
��]xMn�σ�o��a/Xy2���a�s�ӥe�������1u�;�)1�`���BF"կ�ET���	$ɛ3�_[�����P��KP}���l�o)R��>>���}�<Y�����゘��Y�+_l4�O���V!tfr����:����ʯo�ٟg��n���� =B��o8��1���UJ�)�G�A%�Шا*V�h�)ə�z[�y�5Y>�����`�T!-�%��U���YL^��^+��u?�4�DZr��(�
�=S`1+��'6�A�(R�d�«H�JYCì�
v�Kv%��H_q�x�p~��xS5��L�ʅ�Us�xQ�C�||_�w��K�W��~�4��N�����F+k�l��
�aQ�+o5��\vb=�������m	j�;����a�ru+)#�Iv,�ȩ/G���(q�EG�a��[�t��\.��k�R�nHno���(g��k�Ay��#����,�v�'A��l[�X��ոׂ(�L?��X�o��G����gO���ҷ��V��Fr������%������
���⏸M�Ǹ�6���^P*���R��I�FʑB�W�5�Su���x�@�D姌r �hm�$��5{1��-\I%��=<*�k}j���$��ǀ=O��7Xr�I�IfOg�R��vRLG�u�������,ua�
��{fN�<~c
$�
��GB�V5-��w���h��-���%����+=m)B�#&��ݪ!q���0׺$���i��ǔ����P!���J������<1Tt��U�Zw��O��}<|3]��?h�����x��U�9��(���?U�F:�߱�z�#��J�yG��d�z��S�dp1�8��w��JQ����U�}�`OHߕ��f'݄K��r^��1��i�1^a*0��J���륆)ۋ6�:E�ʈ�������{5���hϣ s�*����GO
����~��b��y����b�3�:Lx�pH����@��%����m�߷'��ڼ��l�!:Y�@2�����<d$5��Az�7�*-�H]��/(9�:�U��iЮ3�N�Є�<��\�U��u"�/S:l�0|룍�pȎ@!�P#;C�'z��5�G�$����p8�7U�L�S�EО�x�(t�}~��7��xH`l���U@8�J<��,Dl<�Wv�xV�{��\k�MZ����^	rPύ	����<]���bâh��Aa��K�u�	�d�0p�I���d��Q����<��R�f�a�ݵfDHbl�N�C;gM���j�_?���{Fq����pi��\�V��:�-��!u��׺�n��M^r���m��g �dv)�%���RCڏq���%&y��O{9Ϭ���궪?�X�*^0��Kg��t����ܿԙƄJ�Eƭ�ɣzL{�$㬾�Y���ﻫ8�pe	��+Ш�U�ԡF��/��Z�8�B�c;��7��w'_G������4����,w�5<)�b}w.��hp���S��� ��05d_��F������HB�V]q�*���V�ʭC�#��T��V���"�]�)z�{N�6���=�a���Ǻ8��&�2n7x�u��j�_�����K:��n�����٤�/��W4�KF��ʼxSWM�떯�<���~��s�����
����^��Q�髣e�q��#�;e	�uq���^�6�*����^Y_*��^��Dr�g:'����C_5:{�k�V���!��,@��ax����_*f
R��7s�-�HN����=�5��E���RWG��cNЪ�NW
��׭�Lrv�����b��_�G-Hq�����z�5�����v�]ٺ�R��@�Y���C��2��c��T�%��ϕ�4�,V׾��U��4-�FU����#����O�:C�
��F�i��=$�3���R����{��8#�1�N�Ԡ��ڪ��훶	���>j����}����t*7N��;F��Q���M�4��ϧڙ��!{��aF�B.�G�J��a��Vڝ��H�~�ji���a���J����Vc�h�Ӽ���U�ԍ��<����r�R��x������0��\]�+b����/g��_b��s�f��T��71R���;WM厀� �"K��x޸����~|���p�U5�u���61��3�ͥ��U�S:Ùܔr��ڭ���h�>2�VCa���j�QM]{=�z�cq��x�w��|��x/�CPB:�V�S��l�y��5�P���b_x|0֋r�#����f�6�����׮�֫º�U[B�:O�Up� ^���;����BU��}�F�4�ܬ"hC��]e��N��^��pc�	SU�:q�p8	4U+*(@�؍�Qr�k9��M�\Y�Z|���g��(i��Ɏ�Hp��6�wi�\l
	N�:���nd�|�u?�������Ӈ���
a%��X��<,�)<:Ε:�EeH��3x�Pt1�AQ��!��o
����,R�5�,uJ2q� �f]�z+r]�:��0U�G�<�]�3���iNu�.ۭ�Kka{/�S:S�������.����4:�V5.�>/<�m>�g��F��{g�Uz��8 �v:b�5���[��B���/�U:�س���%{�n�@���������ԣ���-�^��+�br�@��KLJ�C��{�4��ԋ�)dc*�W��c���P���D�T+L�^3��΋f+��͍cԽ�g����X05kJ���+�U��q��$
�x�5nnʿ�4���&<U�!r�nD@mi�4,ð4�E�҈��x��HULyU������|4~Y��@˨��d���/��f��f���z�������^�3d�O����oF�,B �Yå�"�uti�p�
�LW�b�$��.��uݘ�Q��W���S�^��;!���)=�ݛx�Sf���Y�Q����2�{m�O�S!+�bd������v��������v������F��nA��-	Q�^�Bq��.3���24� ���,fg*��[A��D��1#�*`��%]��(M�S����"�7�H�}� ��		��(�=�x%�C]�B��wA̱�T"ª�x���_%YKB'�<�o�nd8�/��d�oe��uYHP�젃@��aB�u�Ş�s������35b�8�!�����Idqӄ+P��C�T����WY͸�x��6�� �F
A��3�dц�&=�i[1�/VfmC/�ޞ
�,OyiS�Z4W�c�R�1�|>��W̬}�-ɻ�����~�n�@�X�;:)S5F��vP&�Kk�K��qY��X�O����V~�4x"kiW,�tK��v��*U�ՙlL�($�X',RH
m1���g�T-�-�΁�t:w(1�����"$<��,f���N�f�M�����UUU	=;�������pP�5ʻ_�L�����J��t@�]���˱ ���ϫR*���C�}v
6�&�7�]*\
��<w�����?^����R�t_���_f���ͫE��Q�j�8�N�W�z��p�4���\|)�+�U�_�Ǚ~�������+/8@fR��L^�+�%i�\���U	if@a��dx�(E�>�@j�G�LinC{�z��ƅM.�K�<��8�Ř�� �G-Hq����7��;�<��2��{PB�����4|(���mH����!��q<(+��i� ���P :~�Q�i���e�k�'4 ڻ^��������T���f��}_~|��]�r��[O��_�R�R�nҏ�FveY��Gj�������k�U���� �l�5݇v��-�򷘠�VB+�!M���b�u�[���k	�ٱ��vܝ5�����:2��paR��
槯��i����ɻ��W28�PՎr!Oo@)@�ms��w(��S2ƭ��ť�1��T`��\%�N��ڡ�����uw�)7hګ�]@g6ˮԷ�tޖ���=�\���($.	�M�xJZ�F�y+��ܺb��&%FXK^ۮ�����*���B�l�:��mR���n䙍�����&P�Pޫ9c��o���
�V�G���2���L�xe���+U���i����b�r�(��=�z4��/7z��t��˽,�h,�__nj���ɰ�#�'-��W�At��b-ス-�b�,r̶A� ��5��&VU'C��Ю,��d��3��*K�ޕJMr+��[������T6���FB�u�����F�@c.��qb��p��2h��,�#�ӫZ���N��a]3%)y���OzT�u]�������n�"�SU��݅�s,����pEG��dÌ��qݬ۲x֪�k�5�u,s���Y?egu�u�f�۫`���]��mL�7oE�%[��u٪�-�:j���s�ؗSq^�ka�ː�� Θ�r�ŵ�M�������6 ��W�V�9̗\GL_m��f��|Yc"}z[��K�����v���x��Pw�ի�����*�֦���l�,�����hu�"���[��R�����a�}��=26��D�W�fʫ�VPkx�s�������N�޻���f�pڣ�)us1�k'#rȾ%�To���r�mM�f����r&���;A��X�]'&�n��A����������*�����`��(,F(1�R�A�T�+3)1VT�`���dF"��ED��
���ISX,R,�TU�%q�W-Qp�*�Y(�X��3�U�Q
�XH�H
��
�V(PQ��(�(�"�q��U,��� R
� ��fSX��)
�k�TR,V�d�Dbŕ�QR��J+2�
�dX��E(�B�A��ộl�9�$x�K�[J�pt��4`N���Z�z^=���< �n��T/��)D��NR4Yן��6�xwSE	��Ě��}j�r�Qh��蠠�\�B�-81xF=^3�픉~����T�ϕ����*j����C�/��^a��\���!cR��l��<[k�1���A�����s�|���vn���b)�8M$Mٞ��&0��H)8{d��0Ă��*p�y�(ö�I�钳�J�U�8����sǝ�~��E �l�Y6ʐx�Ձ���2T�ͳ�<��E��Xv¤�,Շ�1=���AC�t�gy8>P@�<� �ڭ|��7y;���{�g�gy�a�
ɰ��)��k�`
�Af["���6��HV3�餂�]&0�4����d�OYRh�H>Y*u�6���z��w׆�g��H/:C�,���°��ى���Z(�L*m�`Vx��]�w�R
C:� �HVq�p�|R
O{��z����L�' >�H,����0R4<C��}�Ă�Y��ˤ��wE&$<Im�d��:�I!�̞2T�o�w�|o~o��H,=������0�l�&j��咾&0�TR
M�Y=e@�_)
��B�;�1 ��"� (���C����W�]�~��~����*���U����Ա+	�Q�h]��w��7�0Z�Y3�FՏ�Q�N`�]�0ε%��p�S�Re,��d˳'q@�>��,�oH����ꪯ���|m �XbpΘbAC��g���TP�%q���<d�{��1��+��z�z�J���)
�(��z1| ��P�}1u����)����& (��:eC�� �'�E���1���$��{d���(��6��bAd��(�l;.a�Y�~���|�{�~�d�����I=����!^��uH,���IÉ9�1���{�`�R]�m4�{��;�=VV(
,��/~�N{�����J�Sg4��1��bAdû1�2T;�� ��l�� ^�85a�0����M$r�^��$�Q�O�����������P���u���a�s����U=g�b�{I�;aY4uf$Xb5V��0�Lgl����C���&3<d���V������=|�9��7��=�z͝P�����$�z`]R<�g��AH����1{jAd���TH=������ޙ^�<�����7�3�Q����{�`(��M�����S���a�8�H/��2vɤiǖM$�CܤP8�a�r�^lg�1�;B��Ry�>q����\�}���q}`�X
���sa��
�Y�s	�Mوm%Hk��vm��vv�I����v�P;�S�
�y�br�y�}zm��g��w�^o�ri�,+�6{E4�Y�M�Md�(�FXɶT5-#�!Xx�hbA`z�x͡�
)�恌;aXk�H:��:f�t¤3����y����y�Ga�J�+9aQC���0Ă�äs�!Xr»5`oT���Ɉ
�OP���ԃ�!^���'	'T��0�0}�����~�c���8�՞��s
�ޫ���Ǹ�T��A&S���p��ރJ�e
lʗc�{O���1�Yڑp�X��c')�M'���9W�g=���qǟ�G����<�74�Y6�8�R4�=��m;a�8T�B�]��٤�°ε�@��{d�(�Ve�$l��g�� �n���'�ݼr)}�U�11����R��1��o,�Y�N�y`T�������ɨ�����Aq �纪LH,0���%d���6ɐ&o]\3޵���p� i!��$RM t��v��t���p��OI�;�v�gUV���~o�x�[�Ͳ��1!m ��M��1 ��Wy0�
��T6���K���:I^��)��:���
öm1!�H,���C9��^����|�~��r�Rvũ�swL+;LH)P++�!�J�Y3vbAHw[%b�S��s@Ğ�YǴ�v$f��m�6���o^{��Hy�
͉�H/�*<d�%k��9H=�Ę°�)<�$T�k�� ��ݓ�L
$��2 �6�|^����g'�#����D{�IRERT��}����m�H*�Y�%g��6�R{2�$�\�yHV¼{d�4�Y�Ώy��y���M��t�ɳ�1 �t���m!S��ڡ���]�c6�P�NR�w���rΑa�;aXs-���+<a�SIW��뎺��xߜ�}�ϛ���㜓�<��=P�C�`k��ᒰtw`bAC�8�r��vi���1��R1�&'H ��,Ă����u�^=�=���߷sܲV,�:a�AI���q�� ��d4� TR��W�hp�I�:d�p�Rs�}`V�.$<����w@�fP�Fǿ:�6�V���y��`��Z�򣛌?mc{�]0���*��l�sw+�}���]�~��W,��s+�"ކW�u����$���՚���3?UU�}�W:��=��~	���Ǵ] (�2o2�`�R�^(La�|�PĂ��Vx�*�ZACԕ��T�ݞ���pÖF��2W^k�z;מu���ܜ���T7�&$�m���<C�ɤĂ���o(��*Ad�[ɤ��!F* �'gl�a�TR��q�o&sǻ��7�y��M��R�\���,+9=�b$�휡�
(T9�4�H.�d�^a
��L4�ݤ���*�� ���n$�a�|^�5�|���Ϟ�"Æp�ɾlĂ�0�8��E �L;f$0�Y+x����AIP�z�ՓH
,�Qa��
�YCtY5���T�<�}�e��f/���y����>� 1�"������Hyl{�+a�S�
�Y�w7C��N�X5�Þ�<�11�:�Ն�e�3�IP��o'��9�[��r�P�%w7`bA��q�I�XT��R;I�7H
)�u�
r�2�ꐬ;Mn�>�r���钾�y�S���|.�nL9�������`�a׽�1���Ho3,�!��V�Aa��1 �q�f�=a�;a]0*���vL@QC��x`V�����8Ջt�����׹���3����Cԕ�2VM���!N� m��q��xΓq5a��`�L@QHq��6ʐY��&yd�Y�xߩDx<ȏ���4�e�Tݿ��O��L@Qw�0�x�P�IR�P��i�l+���Y�%NKH����a�����4{fyHV0�_u�
AN�'. (��y�����=��`i�nwLH;�x���a���Y+6�*O��P��
A��Y1�L*�I���YA@QO=q �：zo>�Z���ztu�hጌ�1��y����敢S�[,o�b��Haw#9$ơ����9̅�^�h[6'�:�[j��Fa��w�)�$$�����<㝁��
��Ua�L�&2q9�Y+�'�N=� ��ى��a�P:J�Y�;C;�TR8�Qa�'�\���0�tq�ߞ�y�~]�ACԕS�J���uI����Vv��y�7��
¤7i�(��Xaݘ��Y;e`xԇ|����1�wdĂ�%��ٮ�9���<y�{�[�p�����c'����JŚ�xm�	'��^�1x��0��
�u`bA�h�L+
ɓ�1�Y�4wt��������{�z�7���{��8�7a���	�9H){̝$��pe�5��� �@��i��a���%fsa��=MP�A`y�;��ֺ�}w��r�Y1��W}��Y]���4qf�
C�J�z�8=��|d�1�:��t�_9�X)!�d�*A���l�a�Ro=�8�]���
Af3i���A|C��P��&j���OHbAB���x�PS�h��L
�IY�'��I�cXT�\�Z ��J��v^-�w�Ǡ�H�?
_l�@r�=�Oi��V�� ������l���ס҆Yg0\yÁ�+0g��b�^�D�@����!�m���ڑ�����;���?M5���#;"��R�噋�7���G�F�C��q�8D�CYSh���x�Vfoc��]�`�GP�LE]A��+�14o�[������d�˺�jG�m�+7�BT޶�'r��J<�Rӯ�0㝶�CcQ.*��+n��{�v�לƳ��؜�f%
���]u��P��g��m��'s#{k�9�1[����C�v�<ϣ��a��q���׽�cC��	�8ǭz���W�� X�ZĆ����뷝.>f��&�a�X%Yk��f�CEYK�b��:�<�����A��G,,Q�A���0�������" t����j�z  �^�$�{* k�`��_�e
"U�kw�
�=D����fϷ�v�.A1I�X��p�&�X�����9rʒX]��> � Sd�&#�:�}���`9v/�GR�����I�=G9z5a�hBC�=<7�T����b|�|�v|lབ���� ��da��u�Q��{R�NT�I��%���A���)Io��w��u�ާ���M����+f���+��m@�11_|�
����n7}�{^N�����}x�������̓Ǉ_��A�fP�j�_{W�]{�7�(�D�k�b��6������ܱ�#��m�ˣ����B�վ��y�>\W��q�YP$@���->��*5�ziaViJ[淳=����`��kz�m,Z�j��_O�D�U�d�ܠ}ؤ3<�u/]/:�VY�.	t����|���OyT�أ�be�����5���ǣƵf��/-\J���k��|ۈ̭��>cW���l��\0\s����vl����:�>���\x�����W��)�#���K�ncw@a���:��(�1��~ǳ>���Iۯ7I��\=���D��$DXAU w/65dN�{�ٿ]v�$p>��\Q/�k��i�/[�c`g�-���Xjʝ���C��@cS�l��r���l���}rYD-�d!8
��>��ﾦ��7X�	��$3��3� �C�"r���s1֍{ҥ����*��{�+`lo�{�����`�^w��^9�����	�d�uOY�,^P�X��+ 7Tg8����1ͧN����*g��*!��006E�hq�j���C���6�2�a���#�? �׼kY�)}f�,5�����S�]���4��i�(\]dB�ւ"��젇�x�9�F�{X��/���j{$Tx�$G�ti��fE,"%\���v��{�
���_�
2��g�`��� �����S��"d�<v
�[ӑ-�w����5�YЅh^/�5����KMY9Xi[��l��;���
�5�¶ߞ�f�ϙ��g)�R{P�(�]P�����Z�owa}��{�q�C!3(5�A�J����"�ݶ���$@�>�zt�n�yFrGF.��M�
�8�2[ӷ��R��'�}���������]�/��"��j�K{�����gp�M�z��ax���z925-�p�@=��"N�ێ��j���5 ߪ7��#L��da�D�}����G �������2 4+Rn������/���F<�{�Gk�d���͵�<�]"_&}���;^^���GV�=ks�8���(��<�]Y�Q*�����m	ody�98b�J����`�Gv�e��(���2	��f���PjH�yY�����3a
]��r������u�4&-��o'��	��4�d��m�?�>r�Ўˉ��^��>t�	ށ�j�@ظ�� oX]چzשv0v��<(bY6m��oJ`�W�C�]gS��_&;��c���0C�@��'n'��آ�(��L&i��y�7����׷ު�Q'��  	r�c�����+(�&�˟�p���e{�ֿn���y/��b�]b�q�4X�ƶ�̯�׽޿֮�n�ڡo@�W�_`�謯�3��Uzս'�ga^}��#2��Z�#���FÏd�"I��k��g��vl��s8t$:�h֮_Q�^G��y|/;�[�&ǳx4��q�|�DQV�C�>����k�?�</Mskmk�Db��Zc�ۣ� ��^�s��e�ҙ1<a��@8F=U�*�g�G�4�Ӡ� UQ3Zfnk����|��$��#S IP�r�4�p:ACʡ͘8�j��^�T1j��!-1�@�;S,�)�_��j���޿����#Y�q
s ���A6�Ff���oV�(]*�^�u�m�A�Ln��.�z���ݹJP�/E��ࣳ�E22�����C"��٦��
����2L�0�6��Ti(�����WfP�KS5���oL�����69��)V,�N�}h�=M^�1��U�b��Z���������Sq�\��J��z��8�����n�t�ufȿw#F{#zu��'vE��S� O+�O;Z�Q��a��(�ݰ��&l3��RV�,���ER�V;���ǫ"��L���3I7�[d-�F�������5i}s�>�Z�O���U�s$qw3�!���4�vt��^c����:a7jķ�1��,����A����j��*��xW\�u>�.����^�\�.��V<�K�H�fq���M��5�1�[�BN�a�nCs�|�~>ؕ�L��^��iGB��̒�Gۉ�*���\�o6��A��J]:�+NSϧ͙ �yuc:� v��v�(�r{��)ю��х_t�}ٷ�k3���/�bW��'KHLV�oa��edf�+�h�X��������ΰVi3J�f=�p �]���F�X�f޵�#!�Ju�I�c�z�r-M6c�R��K����l��ڽݴ�*+���OX8�"/�����9g"�4��)p��m���nՔ�L���Nt��n�8�!v/T��]r��rx�j}ѫ�
�7�����M6����x��"�]z��U����w�7U���:�\18q�d����C#���Խ%CPֽ�=܋��V5���]]Cbjq�Yg^V� 5�b�\t�։'��"���9�Gҹ�7�g$�:1��(���NR*EJ�%B�T�PDlEb�[d���[VEcJ$�X
Q,ee���Q�E
�PPE\d�cl*�,���QU�X(1U�$�JکQ6��V+l�XfS��PTQd*�am�J
�1�r�QAQQ2��U��2�dR�cmSe��d��,�cʢ�[)PU�`�j�T��11V"ԉ�
 ��b�ina+1R�[j�j��lU��+(��Z�6��F,J5-�q�+)e*"E���>�(���y(��*���h�ד1 ��s���هi}����܇nV�,n���X��}���<dEH��gO���6�;"R�R9y�Cr�6`-��n+�va��4�W��b�#j��&#�c��6���so}.�=0)I�k���{N�!@��P8g�z�c���j_;���·��F��kE �ֺ0
��/Ϟ��G����L�K��5H2�{�}uG!+n#�Z�m�V������/&�"twX+M ~(z��p~��PK�#�Ɋ��ե\���.>��P�[�󳡴<4�o�s�^kD4h�ڨXl؂�F
_���{�r&5��`��~��ؤ��H�Zȡ<'fw��[�N'�N��?X������:��EV~>~'?��.9����fl[�_��"��1�6��4����lD;��3u���u�EfTE��W��,Q�i܍b�=��'t���^R�w�c��e>����xRQɩ���QdI� ��8֞ʁx.;��8*������Wf��0Q����=r���{�>�͖��������N��a�APA�m
H����0�;U��l��x4#x�u9AxOp�@��\@�����պ���R��!O�Uo�!���#�����#��'�)\\E�{�n�/�u"%�r�v�M�CATbϳ(�+~���%(f�7K�b�Ǭվ���\�*�i��Q_V��E$�T��Y:�u�y�A�#q{�GG��8;5�[U0�~5�j�Kyڞ����ObR��@�@rgД�B�2��n�Ly$�I�W+G�y�/4U�0������Y��c^LP�X&z��O��-b�W+�.�AԬ	��q益��[q�cP�{wKx��S��m(v�,����ƿ�7�jc���YxAep��O��_}_}]�9�z�C񏙮?
y��A�1�Q�xV�ֽ]S��龜(�u�u�K����_!��-iy �)z�L�aV���sWϛ��Q��f}�q�X~V 7Myo���!\���]5�+�G OHQ�zvp��]G��!P��u!2_�o���z�>`��dp0��H�D\G,0x�^�!q{���0x��qz���^>4���FڑD�2ϡ%B&�^�D<~#Z�^��6������M���%��nv{޽�p�Q蕄a��D��ddx�f=��'), ��۱�2�{s�!ګxW"u�}���ؠb�E^�r��z��+U$,�>qQ&Z溲	gI21�o~��xZ���=(�K�X�H�j+�+W}�O�6ay�FW�y�ܭ��b��J���ΒY"����fP�fQ�㤝j�`i'����]/M��,�Ϫ����Y�͔b����#�x�Q<�O��(x<5�8is�_��{�?���
�?Y���T~�~tL>K��j�}��jc�������J|,�� ��}H���񯌘;%��k�)�C�>س*��,!W�����n�p���/n�ݽ��X A㥝Ň�:=��E���E�QS��WB���:�Y5��az�5��-���F�͉ä�0��B>M:�����Y8#�� �B�d��]oF��*υׅbJP�Qy}��L�k�����o��b$:\G0Gb�U���GG�!�֝w�ၯ_e$�����
у�Կ'��QEF�����'�C���S��q�c�B��<;��r�`�j���E�쨒�Kv� �E�R�.���\V��2a�9[G��y%�(po2����s�m�]~����}���>Sl�7�ٖ;�9�f��Or�8!�����X3i�7�ҏ)b#˖�@�dq��Q�ҭ�����N�^B�ݔ����QE�f�ϓ$���@�q�O��L��i�����C���}�额r�:k1A��*{o��DP���3s|��TD�(s�*���U�+C�΀Vn�~\j��)߼��ԾF�5�Q�]b�~��H;�����@e�b�)���;���.����^�f�KD!PX`�|I���o���ޤ�����U��Uh�0!wGLQ������~
n�١5�I0�<�	�p���;#�#`!�ոz��Q�wP�WU\���+��ȟ*�6=J=E�#9c��t�
�H*�C�U䏹�s�ڑ̲�/*���Z� ]R�ЄA���yj�l�x�R��\x��E��ѡ��C�/V���پ�-��^w�l?]�_������nc�5���h)ҫ�!���P�2�q�?�=n�����Ռ1E��A�CX�Tm,�ʴ���y�y�6cjtoԑ��1���ϻ>y쨆ܼT>�9wB�udip_�=t�7�_�)�����ix~|~�v��وo��}<~{ǀ�
�kB��T�ߔ�q��n�6�����2K�w��yк��q�����XC�m�Aw~�]�&-!�H�f#hPH�^�Bq;U�^�V8�ͷ� �ϢϮ������+ �*�D:(s��7�2O^uSg�|�ů�X����>#�.p�a��q1����9��܅r:X�/V�ƴW�*:�j
���wu�Ytzp���wm�t�DI��*<���.�P��x�u��>.�#T%+L�����㎰�)��7�wN�fC%��_-7�\D�����y���/kWȿ� ���JI��xp�aKT�������V�{�i�l���޸��my0����G����H��dRz�Ϯ(��b-�=��F�Mĥd:�g����m�D?"8u=�r�k	kpc��G_g��Pv��!g"��_�����lT(W�~/��V��?;��𴀫�0],�b2*���q����r��) ��Y��J�Tk9R�L�tU��Oq�~����/�HP��"%�!�8}er�C^G�b��q;3w��Ф� ����Y�{������ٴ~S��d�aL��BA����C��T/(�棖<tD;J�ꋌo�N����ɜ:t��|8�6DF�D)=�
�88-$5E�[�}�M.�k3u$J�z���A�f��5t-nM�Jډ�wؓ�0��aO����<+��MjQ\�Fi'�K�ɴ��屼�>�����W�ӂ(��L��My�ϰh��8@�M�Ǵ���\�6��j=�J�5~'�W��JM?���r�H�O|��{��yDřкT�%�g�1��x{|���w��z������U�[v!|�A����%�$� ��E��n�7�Y`��RЈ��Ȁ���>,�5`��5({��KZ��y�N��t(�����̈́(j�^���}=-�y�yv���C�ܨ֝����3J���f�y���N��?�gE]�����T��S�C;���BJ��o/=<q�5��*�����:}:������'�#�������F�֗уcÆn/�Ơ�ӁƉ'|���2<=��8&�k�K>ʹ��Z
l�vۘsGr���E�Hn7����ވ��mq9]']�o��%]����![�8�-2#/$�>�磌�&޶��/i'�PZ�C�+�6:R�����Sf�pA�<�=2���~b��T���j?/����{�c]'>�Ԫ��pȁ�̑ڳVc�PkN��d���ov��*|�����	��Nh�؈6cܙ�b�.N^�ݩ$������:����������R*�V���,�w��{�G��F�����j�l����8�N���w�z�Y�^�P�C��	���=��}v2�t�Z�����54�,M=_x�¤z�(��t��Qꖙ�^Ke���8�{�#҃`;%`j�F�9F�,qӢ]���xͷ��/Qm{��R�R�>����S�,j�o�=~�����5��f��<��=)���Quv,M�[�K��2����cmpW�f"�/������di]��>5����}Z��{ݒ���W�UT�F���˄�u������\s�n��n�R��75�������u�|MB��`���Uu�����tuB7 �x��9���ת!3=�a�r���C5Cox��f�`�(��UVk��"uw(#d�Ig%�Ъݞ~z��ο1+�#H�&iaP���g�Y�Gy��j��<z����|tۿ[����jQv�xT������{�ϝG��/�nD�Q�E/8���;�1�}�~��J�qM�9"�i�t�P��|�k��Q���0�Ɵ/��wk� z'/7����l�1ߔaF�N0��:}F݁Ĕ�|�z�ܵz� �!HQd)=Yg�F<�J��ʙS ����G7�57��m���<����l��:�쮊��t����.����vh�Ec���c����E��8��,���1�_bZ�4n-"
3`�4W;4�_�:�����V_���j��Gk�uF�\JM��{��"-VZҭ��kk�k�5QP
�	��u��a�����w��t����w�vwcX���S�.@��xu��	9V���nHp[�a�99�;%�Wi�SC*�&ѽ����;s5j�w'�	RC���=�o̦09�0i� D��M�WG%�ޢ�u�P�%oM�(D2m���ه�˲�uww��b[�]Ǩ�]d[��t�k��@��yi"��Y��5Ha�H8�8�l,Sd)��y��q"�BtJ�X�f��u�[yZ4ڕ�X�%��6�"z���
��!�T.�Co��E:��in���Ѱaq_DQ̵�(�t�Ɣ�+-\�2X�Z	���T/70�-�W�U��u�r�y�[Ynm
ȳ"ٕ+�T�e���Ru4��^�^������fG̱�yܰ��C���v����5���*�<���w#�D>�T���^d��9��7m]��,U�1L��W�Msk~I��[�ɜ��u�m�-2�3�6zs�:$Υ�%h���Vn��������7O��*$y��-��
����/Z]�y��k\��_�]��Պ7�f�����Ɵl9Z�-�)�)% .��-�(���3/2�r��uv��4�>1�4��6+ �X;�mJ����(��Q�{!�}�YԸ�h����:CO�Ո9���\ 9M��ړY�Σ��1�y/L�T��.�[�6I`�����o���ziܶԨ��Q��0T��3-1q�R����jT�V���X��Fұ���.2�e��#h�B�-��[m�(�ŭ%eb�j�YKF�l�lU-�Yis
Le@KE��J���m"�ck[l�Q��YYkB�(V�*-�1�K�q���emm����$m�Q�m�*$F�V�-)\̉�ą`�m�F��,(Җ�r����-,�2։j��Q���Z6���[j��* �Ȉ��Q�Vڭj(-k���DF+���33)jV���V(�[b����UE
�E�mb(����jڥ�5(��ưQ��.XfR�H�(Z�
��(�*#*T�.RQ1��m���8N��N���A�z��k��4_r1�b��%*��hOp�<u�W��~��4�'}?�����n�^���~�DB���ʰ-���]i{d䀦Ϭ�=�t�  ����!��d�n$uC�.��J&���oM����ykp7�+�ݏ�C�,r��k��{��p�q��R"zBq`|�ܰ�����2��X�~u_g�Pђc�m�8`�#C6�e�2u������kHI0׬����L��j!�#�As͢���6�ze���Z�U���b<�>&9P-�V�3&��%����d�e1�k���(~a}��L�6��Z��WZt6�j�����2I3y^�#Ձq��Lz�����v.������@Q�Ѧ�����aac�"O��݁�n����������:�{���`ᔕ�_�O5䶩�侻\�9���FGn4�S�:���`Z��e���#g��HrfV�^V�Uu't��{��oC�����>�{߮�>;��m&�S�G�p�X�B��XG;�P�j�畕��٨�0�KE��\����K�2){"��^�}h�^�j�v�� ����	?�`���PV�|�V���>�҆Ȝ��_e��A���Z�n����3�P��F�Ukʺ������@�XC���+�Ȯ^i6���N���R3��̪���8���z4Tz%>A\�t�L?!@�ۺ�{ī��a�~�J����
N�(�.��´�:���r����E->-�SZ��8�J�Zr���K05��2�([h����a� �gKjq�0G���%)"=ϤIf9	��F�%A�|[Rh��z�ݏ	`���Y�����eJ4l}�f���?P|SJEw�/����Ԓ��Z\�*w���$Å�5+o����Bz�g�]��z�s7��31Ⱥ\�:���t���w�_[]�k�5Rܑ��9�m�N_χ�H�_��fP{����+�ʿb���:.�=��9��f���'&F���Ȩ�.�`�^@���N@8��l�W��'*�gԏ��pe_�h�C2��J�%@l��/S��~ɸfB�~�|
���B{�g��Y�i��\{��-A�@�������^�z~p�P�f��]:���+`~�9Tgf+��=�t�y��<l�jVT`�\!�dDh<+���IѾ��ŝ��z�X>>��W<PWNP�u�8m����^�<�^LU�6�p�ܟJq��(jZ`R�B�G��(*�(`���g���N�=�{���{���K��Z���+��P#�[��3��ށ�!������Z}ۿ_\�,�Zͬ����V����̻����w��[�ӀNh�����+)�n�:z���th���J�<������#!Bp9o�)A[�Ұ���)��C�J/�x�t�g�����C�|ò4�?y�l/CF�$��'�
�j���k�,��!�Us�Z���ʋ���N� �@z��|�\��`�@V�����G��ž#�{��UY��Dp�8�B�{�z������X*���u�H6����.����=�Ӹ��Lg�U�ܾVxv5��'__ʚ�4.�H9�}e)!�>�8<*�ܦ��k���Y��Xc�U5I����!�ԗ[�]/|>����ϯ�%��ݠ�����&�H�MAd�!:�Pb�����<+�j���GA�7�ϗ]Ng�t�M���\th���4e��I3~����7����9��>�=�n�Xlܵm�7��mX��0ߩ�Z{��Գ�z��:����^b����Fd�-�Z����b�<��!�w-��̨��
dY|�]¦Y�X�Yy�;�C��hBE�/�}zR��Y�[RZ��ü�ǃ:��ϭ�yWB��|���J� �y~K^绿8<hP�ԕj���S����\�d��P���>ٟw_u�z���?�h�_I���\	#x�"�,�:}'Z�Bi�5F^o��Tv� �f9q��KBBCm"��a���@���r�=uoM7��5���xW�0mѭ�:?&�zk����(��M-3�:}�h@���������j�{�&��<�ܰq`p6=�����u���:$.ٷ5�v�נ�C���#�1��4,��t�1w,E���=m�}���Fiiz>�.#���8`�#3�����t�{(yxQ ��4��஻U��8��{�1[W��d�Ԯ�~�-��Th֥��H���Skt�#�Z���c���͔D���8�z�w@U�����HN�z�GV�T���?�Տ��ua��1憕�HP2%(�2���^������u�vT���x�xA� ��A3y���Y��MP5j��8��Z��^�T��ݞz����`����v�{#�N\r����8Tݩ�͸�\TY��A��ʵ�jC�F^��|���Sm� Zg��6H%�q�+��b�,��x�v��t� WS�
��hyd�^�C��#�	�-(��K4���8h�%{L��%�u^lDh3���H6^�$Ut��d
��}�k�2�|��^��8!ø�x^���0hѣ����¹��^��D\8�4�[}T%��iM
��n�y��&���:I�S��JFu��>�)Iӆ��p��:�DO-���@Ѱ���m^��V7ݎ��9V�0W1X׮�s5�M�@w<ߓ�{5��cEꝒ�dq����Xo�i�"����� ��{�mx�Ҕ+v��.8�O��9��x��,�k�@s�ȉ��:ʑH���DV�^����8��r�}��5�_�-IKC����N.IbYǴ�}�}��ח#�2[�Oz�;�;'x�7d�x0�j���I���v��Ͷ�������NM2�d�\�9z��K��S޻�T��;^���H�S��&��]�8��z�{Ԭ�������GPyso�m��)[�o�x�u�.�+�gi}
�/K�_k��bq������W�X��ߐ��yMC��}6?;��������(�j���	����E���f�<����a]q�q��/m�O�WA4{��G0�]���E����-I�qi�����&y�Ʀ��U'�\k�u�� ������6��!���c�Q�,E���rtra��1�ֱ���;�R�.Y9�_d�x���YR��Ղӳ���Y�*G�=��K΅�#��Y�lT�&��0^�����f�f���t�� ��;>�Me�a����W64�N�������

��?�i�n�޹�]8R�L4��{�J�&j�nƛ������9b�v��u񧃭�B�ۅɃ
r���t�c�ua4ziӖ7�2I%��0���O��������������C͜Jm��1uV68C�R�Q�7�2|Ω�So%`ǎm���$���8��]y��2�oGkx���8Sͷ;�w<.�c��?(�� ��u�~��"߅;y{y'b�\��W�����5�݋���}=�\�QT|�nnNB���&�9w�J�C[�tn���ɻ��6�g���P�l���(v���ۛڌ���4�8�h�z����isJx��5v�RfF �TenEڛ�u�}3z����X���i���N
��x��m`�J
���s$K�O���*bt�/��^]���̽��J��T�U5̛�:9�ؤ����ww������;���3����&�)*z���<�_�
חŧ��ܙ��@���Cݘe�ן�q#��w��]B_X�f��j4!��K���;�y��Jw8ŧ�o/_�W���o_���G����(mA�Y�:���~a�70��Umv(�[t%��V���۬G�D/��/�>W���^��*�Q�;��]�y��Z̾��^�r�N�,se�-%��^�V�f=��&y����,��V��U%��Ch55��%�S���VgcM�fnt��[ʍ��=����%=���X�1i�e�m�|�^/V�]�zs��Cc�S63��tg�)�w�띙ټ��f(z�۠������\�S�$C�Qg�,\��|\���8!��������_��7�r�1���Z͊d�Z��`�&�7:�B08%<��͘`�Y��
u��:u`��R�g<2��2�*$�E�m*4�EB�#]���3���`=�"�Z��%����o���d�����U:w%o-،L}R Y��V]J�Q3-gX���m񳔺VzSY�A���_Y�(U�e
�f�{@Ѱc�t9�Oa��C���5�@�c^a=D��)e����c���2�\��9�),r:�|��OQ�S3��4���0k��0�u�r�Xjs\C�J�TZ��/q�)(�<�>L�r�Գ-vf3�^�D� 4[�1m���]�v�<�Eٖ
���\��D���9��R�_h=�{I���r�ΆL'.'�>��]�������ο������x�'�n�9 �X��{FfPC ���w�!��'������֌뤳�C�)�:]�g�:~�e;b,�,.̬(P0�C��+·�Ly����>��;9-ܬ�a����8� �O�\���WMZ�{� ����2#�~B�.7!�.VU�s�*f��P���n����h59˫���ݎ}�9�۸0XI	�.e�\�T�K�*�>�L}j*�(s6�I��Ē'���B����ٙ���9H�]�U�&ռ��G$�/�Q�A��E�B��,�ˠ�s����&Z�7t��W���7��\5&e�j�a]����j�\�]HrBܨj��zO��7�C�K�y�Ǳ���^�2a�r�wK�q؇�g�tu���F�fGI��J��ѹ"W[`қM>���uő�hr���F�]�!n,���/-���n	�Jނ��˙]gGF)Hsъ�WmGr�ΐ�Me��	rf#�s�d�,��:���9�ȥjQjPm����U6V*�e�fE�G�#lZ�
Z[T,�X�mUKh��-J�naTTrʊ[EkU��f!����V��H�%eUh���e�DƢ&P�`������,QX�Ե"���kZV����U*TU(�+�E+*��+mQB�J�mik-��Q�[
��ڱ
�X*���E�����,b����*�a��1����R"��%�Q�,Q��EDUT���Ym��D+DPPmR��"�,��,X�Z�-�X,�Q��-�kF�-�-���&5E��E���E�(��2�-
ª�1F,Z��",X�U�A`���&6%TT(�������?F�=6�)�mMJ���dV7�S4���|u�_��<�{� -�,�����>��� �lW�r�.��w]̙�����S�$5�)#� ��^���_{�����T;s�zlG�x	rc	v�x�Gbx�o��#�4���W��k�M܃��x�G�m8�}�!�t��;ֆW}�����[���	'/p�iS�����d9���f����!��������8s�e�/]��k�FU���;�
����[�S�s�?I�x��&��ؿ�ܝ#���圙*�-Q<y\��G�7�
)���N�sNN4�U����umǓB�~�S�~G��^�8����)͆n�v�̉�jp�Ϯ�b�����T�>��WN���n�Vj�Z��iD�t����d�����J��bVKy{_d��6�P��l8��r=�!�6��HtE/m7֫+�g^�>��+���&9�M�
�X�#���S�<zcl�RZ��M�.0�L�6iR7���p�sm��4(�{��$k�k'��^y3�5h:{?�L�Q�(�;����w"�ֵ��I�ě���˜��N�<�YV�y��;�Y@���;�qH!�l��!�ڊ��Mx��p��N��N�JD�͊C�	�x&��^�f_�+�y�b�^3�{k�����sj~��[|�ή�+��q�n�Y�R��܂F������iPht�@붟,�j�wdA�ѣ�u��⛦(�rT]^��tdݾ�H��.#i@k+BK��e�s��9%�)�x��ɛQ	�X�i6���u�^�>�s*ܓ��(�a��ޭ�;��t9��{7rGg�S|
u:�;kޠO��s�q�^ث�gSwܡ����'�G�M݌��聨����8�ҙ���/��8M��Z��R�65KT��~���Bƹ:�ާ��Z�8['z|	8�Wu�>��44r�{����Z�̹z���`M�ԯ��=��]��2#�]$��Tۮ�<#v6�ᷫ��u>��,̧��3L��0C簫�"���ݍ��r�_W��G�yz�;(�Bc90��[���ѯU;a3*ƻ�(D�[�O��1oX�t���z*I�(���Α�L���J���q�� ����w����hw�c�<v�ܶ�,����Ni�Wgr̓Si������]R�7q�6���n�=l�tq��
�)�
vC�La�$b|5��n�Kp%��A��c˦�����@�C�V;!�ن�c���%��z'x\�Ҹ�V�?^�d��_��{�Ђa6�P!s{W�_d�x���<<jy�wd�� ��A��7�e����7��m�����}�9�v�
�W�C���/Q�Pà�����ZWR7~9�hd�}�Y��,�mU��wC�t�/Q����S�a���\X�'f퍘�b��>��I&��+!�D�S��N�taX�K\7Qr�lY;4X���̝�}_W���rm�a�y����w���K��/x��y���#�b&�C(1F�]����|5+�R�۳������I�ac�s��R/��\Qr�}�F��i�ԃz��S�]�y�HPj��T�N5�l���\�9�7�E*RV��u��ecв��1��UԙqX����O�����Z}�����rc�O��#�~��h�G�!cM]�}�����q¡7�u'v� �+���7=cf��Gܚ'�
h��

��z�ڰ�}t߂Y���Ԯ����sz R������h���+&&�}t��L���	��S�V-�A{n�4]=b�z\ޑv§�!���,��F�"+y�yS��2�Ϭ�^�:��;�|> %�I=�0o��@s�"}���~��qtV�y��Q�ֽ�z��(Ab���-�49]�C.�*QI�G^{+6no���ci��N��������ߖf3�����el������g���p�ͧ<#V4[�����u�cU	�@2��j�nDY�gDU�㫖Gl�is d�zp�ì2q'�A^�c(p��e���gbNo�Ɩ���ߜ3^GnTdza�����%�&��X�x^�a�F���u��]\>�,d1�F�r�_�TO{[]��n̙ȷ3�N�g�R�y�[�����%�+�N���zhڳH�l��=u��Þ+^����g�Q�0W8�)Υ/��:񒰅����~������U�2H�����n���eJ��=T�u�N����r|���f�j+�5s]����F{mˋ�b�:����ň����w�����1!�)r�%Y�`���z�n�S��{R�;y¤Z`A�f�]X׫~���踭���ֲ�90���[������Z���Wp�~����;ΝLg�ܖ�Ք�U��CҠ�3��\=�T�f=ٽ�jʞ!]����&eF��i�Wy�?^�H=��$����Y'ӓŴ�Nߵ���B��I�����Ә숳%vR����/I��-Vw�*M3T��!�������b��@�S��3quqO-�N�:	s�L��w?��۹������rh�s�9��&�u��{�}���G��a�f�)�Rv#�l�s%u����}���>Bg�mAH�1��,6�j6y��s�'tT���i�P����TN����w�U��b�z:$0�͌�(������*%Y[>�,G�w�ci�t��b+�-}�S�2��ε�]�rQ�rF�%\YHq�y��Xpxe��)�K�y�H�ԏ��ҙ!1��C�z(Jz�+F�0+�3p��T�L�	�{[\�B�*đ��a��I�.��t���G�I�N��1c�K��"�j�[3pނ0ƪ����Wy\b܈�˳���0eޔaK34���dZƫz�	,�IN�:6�I$�-�F*!sf�&�-�OX4�eF���ڔ��Y9f|j��w���a[C7I>p�~9!��#���)�B��3q�?;��?y�*u��bZ9B,A���!N�Y��5�S�	C�r/v+�+��`FݩZt^ҿ��u��(֊t=k�9�׽
�5���i�=/��С��#�B���qE*�$
>)�OٗXÕ��[����B�j�4����S�vl�Iv6�4��D��b�П9��H�� ��0ߑ��ֹ�tɴ�q�YZ+�H��M_*M�Ǵ���n*�oVj��׸��k��6珨Z ^��,k�����2���FN�r�tUaD�(6;\լ�g;-K#�RK�SvW����0>�F:8�	r^ܺ��}B��$c���]g�|�x�`�c�Q�l�Bvp��#Gh��
���hm�+:fgi�2�K��?�&z�L�T;�Vk*�@���Y4�6Ysz��ppT�0lyRF�P�z�O�4=��Zsz_��͹0+�9����U����F�OE������t��d�6\��Žӌ�~�woEj�����@�m9�^�����e�<йQ�}�^�WN�m���n�Ղ�:�
x�M�����B�E+��i��5�/b�CRv.��:�����2meH��JB�r��M����p-�Y��+x���ޢ���XI�C����f�Ob��p�|�#g�Af*Z��qн�����= _Llq�ùݜ:��bǪں=�U�old�|�2�V�����v+�:@�_m���Rp�V7��ԳƜ�vH���P]j�:�IEV��7qdo�i�U���[���)�1���<M���J���_K�ˈ��.�+����ۜl�aq2�*�(>G��)�a�0�&+��ci�q]i9-^�U��*P����*e�ض��M̬�]ύ#�m�rR�cm�������W#RȺ�8���ս��2���PӥP[e� ����X�qm*����ծp��ƹ��Ha�7�4�lf�}D[&u�W`��8���z� &�K6�%F[ԝ��������NR� P�Y�T][���˳*I��[n����_m�˜Y/FYz8+�m���l0���&�ʝy	���E,�f�����b(��+���AT�`SӦ�^���@+N�ʈ�:�����,��y̣&r�P�fB20a']N}w�(v��W�n���ŏ�p�d�{��XM�N�p��5+���zhY{��׺Enڨ��6<��v��+z�-���d6it��=���Õ%�-�5m�C�yj��� cj�!�� ���_a�h9�Qn�U��M�ڙcj_;�����z-��|@��f��%.g}�W�f�@9�Y7Mu�/7*J�k�O�O�eq��w���l�.�A^�2n�7HAk��񺇈5o��d0���b�_:�Ps�+��u���� uh
m��lO�n}���=v=�����t�����.Y��i����";���w�1��[�lF_�bL���Ԫ
(���[B�*�em!X,DAl;j*�*�b������-�m(�DUUUJ�)R��E�U�
1L�TE�(�0U��b*���XP������b�"
�f)�Z��UZ�+cikYiDF���Q��bVUX���ԕZ¢""�T��h�,bV"*�q��([cU
*����֠+QTV�QQ��QTD�-���mƊ*��*$AUX(�R�E�H�(���QEQm� ��"�P�*"�j*�,�*�iQQX��#`�V�X.Z��b
��"1X����e`����UQ��ADDP��k���9�<���nf�Jw�c6����kN��^9}����ȠcJe����P�(�O��+�c8G��ݭ�,����yח�t��ѿ95��J�'���^��i��\)��o�����s��w�_$�3�C������'.���5�}��ʏ��6P�a���?s�iO**TT�K9��P����:Ns7�F4$~��6+j+Q-�
O$o*�9�z���̈́4ux+�;ٜ��%G$�n���5Ԝ!y�=\}\&/uۣ�rr�����%:�E������k_��"����34����r<2�¥����F"������ù6r<%�')W4�� k���+ip�Z�"z�^J��T�^Iy�&�7%C*5���.�[��E��9��?^Q�[�1��Τ5�g�^F�A���}^��~Y�o��1�l�|�H�TB��I�>��+���L��]q�>g���}���܃M%��$��lc��7;ֻ��m���1�3Q�yd��OyͶ�H"�L�.ʨ��r���������\K�z��
@��V��4�m���9��)��8���P���"ˆ�%��*�o���3W�k&�r��i� GW���
/lo��w:��~��ӵ8�m�T_8�O���5׃lF8C��������L�M�F��Wq>����L���%/��W;��g\r�R�y�p��'�h��e�N:ˬ�D��*����[Rc��(�G}�h�G��&9��uΙ�G04�&�߈ȳ�w:p���}���s/��jv�<o��U<+����F�*��)k℡�I�>�<�}O��nH�B�<f�X��D�C��܎R��y�Ռٻɒyx=�F�z��uj��lIol�[Kn��&��\�o�ʄw�:�}������e��K3=��Gy6�,�EF�<���,�R�x���;x�S��R�S�15
�^�\!q���k�������q�s�'��ר���g�t-f�@	�J��.\(J:�%j�A5�![;M�{�ElNN�j�_AX������&�GɌ�����v�̴����)&˓`Q�/����ߐ��H[%/o�y��-�e��z�,�ޠA��SnL��v�s�����J�)�3J��a�c�ç��KZ�)5�=���o�L��"��k���n�&��'w���qu4Rִc��|�\^���<�g�h�1�"�u1X�s���d��ߏ>�
#�uP��#��|x�&Vl��[�B� ��޽��.��Wjp��^i����>��$t�5^�LM��n����\�����C�WF)"f䄛vB�̼9yX�7l��T3z%э 1�k>n���ѻ�<��S]_D�|��/��eay�-�e"+7�B�/��� �WxU4��y-}�9�6p�>�lUɹ�$x:W�l_{���`��qeJث�����ڔ-�ٺA*�7+�hy���t�Ϯ;�R�#��)�\���\(g���XcB��:)J���`"�أ�j�B���.�c�O{"���8�f�P���!���>���E��i���[�Wa������W�g���2s{�˝��s�Z�y�y1`��N�W����-�]�f��y}\���$
x���d����^38���4�{ڛh%G�!���3J_��7[W�Q��U��P-���|1���S�n��au��M���[����a��G�j�.�̬���ݹ2e>�e��1�����X���>�\��Ƚ�%ԕ�Y臼H�jz�������v�����>�Y���35D��P�=��KD�����ew�*���_����2�Jқ}oM��Y̦��_{Ga>��k�q���sjޛ��^t!��{�ӡ�­�<��t�[Jcie[
�\.%�^�Ɔ���w��g�m>R_��w���Ì7�x=��i��-�j�����e��{a�8�t��Mt�����5=�j��U��!x�9�s�	���`���{s\�vR�ߍwX�I
�Y�I���![�$#E[Z;.�me�HZ_nb��ݐ,�oj�`��w&ю�+��zDa�;mN门�u����i�-0�ᝡ���<C��M'6���W�攲�M���9�!�*P��g[�h%�����ڟ��-��J���/�͋צ�e�&�ݠ�L��werT�tO�]�]c0��<�
��Zƭ�q�9���	n�J0`9���cZ�K��F:N��F�0#��'b���o�%�Xs�.}�x��A�4��h@e��|h#^��4u=�QT��\U����������޵x5r+�9.�2��>��2OY���-�.&���ډ7�"+NuwI)+A>�����������\��n�v��S�,����8�z�2�Go�[���ջ��ڷ�5|�[`�<܂�>�+wsc���K����/gKZS��P�s�-;y�o&r���+�(T��!�4X�������SQ�����WХ�	Zs>j����)X��v�l9�E枫����7_g݆��P�C8G�����{�K)q�Չ鵇�{���@�^�=YV|)?gj�:B	�|�e+��];-�6C^�͛�6�c_t.a�3M}�]��`����9���϶��'�q2疵n�hl���_a��PjS J�A����y�]&�&�Xqxjv[:�x;��s�3�]������[|����|F,��4�+���j�A��TS��"�R�>X�V�֌l����4Dƾ*���M"��'���Z�����|��:�E��P��4m�L�^�1���<�D�>w��srNMӘ=\�t�D}��H�T.�<���#�q[�^Y���_��,!���m����_g#'�Ew��v*����t�c:���EJyy��=+:J��_���ݛ�D�l�on>�9�@Ұ�Ց����������^��YF]�	��11�S5j�� ߯�{�Q�[���ݧ't⵻c��X�/c���NK{(��U)i��}��f��^��ѧN-HSdo���Ƕ6#�0�nSo2��W��"{XVB	nu�t��)��S�xd��1�\�F���`g+�.P��={�����&�(w�e���F�9�^u�ρw��c�͑��aw�<k8�z�Bv!����%��#-�H^�fޮױ�S���$��W��F��a���|eeʒ'�������}ΞL�=�x�Oh^��j�˔9��J�^�O��(ZF:�F\c�Mk҂`�������9imE�"W��G��K>r�I
�{��Ve��*{�u���-�\��w�	�X��8ר��Ƞ�[�f�{�d�Ì�o+�~���2�vY�XQ��g���<�%�D�k����򤓯2]nG\��j����,�[�)u*{nE�n9_��W,��ѝ�k�)k����v
{�*�V�rcC"�iر��ȝj;�{&'K��s��(;vY1�����E+�F�^��,Yw$tkMȦ�l
/3]lw�9�ب�%�ܮ�j87.Yw���hF��]b��E���v!���ml��vpr�f>v��_*ނ�˼ݢ����X|�
'V���]ء����� ��1N�����pYN�N�<`e�Cd�c��*���Z�����<ڳ��"�J�D����ojWW$��R8��6�e�r���H\ȱ�E�����.��2J5��R���!�-�2�U�7yInjV��l+rK�(Η�(��Ay+[��ߢ�ٚ�d�U.]���«d[.-2�NirvSR�w�Ĵ@���W�{�]��1x��_�ה,��ll��Ū
gE���9F�����o���ؙ�+1�{K����=�,���a�����Q�a�G�:���}�lq"��H4��O�mJ��bq�E���"=�n:˼�({*�X��c5�z��S���FN>�tL��۶$�6;V�UѮ�����6�Q��W5������'��w�� җ֤yiTa�}��-�l�$m��K�n�R�8����h{��]v.� Uq\��Wc*�<�R%���U�u8�RtH���\�*�x�Z���ʴ��KtE�ƫ�(�Ƕ����G��~�4{�mvW]Kn�˻��A}��H�N��k�S�5WBP��s���٩�(��eؾo��1vK�N�]ŧ݈��B���Gevw���I�Q
�������u{t�q�F)��ڕxm�c-M@Ҽ�E���ةK�U,)p*VU���T_57�Z�/7���f��Q��s��lX�G�&���ꮑ1F"'6���Q�QYb�0X"��b�TUDAV*��E���`���(,UQ��EUDDH�����*5,�*����,��1X��UF"
�UQTE"���QX��(��ň���)E"0QDZ�Dc��X�"��UU**"���b�,eE�U��W� |�Q��n�u��L ����P��س�)����D�-N8f��tC��Q�n��+z��T�9�������0�c7]qvr�XiX�a.����u����T�}�V;sF(��h�e���pr0i���򧚾f����>����BP�f����;|�:�tQyǊ�[�n6ױ�^����>���L��1�).=���m���X�2����ز?Fe�ۦ�����Y�5�ߡ+��$M�[?l|��	�qڪF=ŭn3�����(1TkĞh�����tF5����_��'�i�r�GfM{g�lf�(���#�kcV���\9����vR��ӏve�\����~ϊ>���J�fV���}y�eI�@�¥�X:��Ru���FW�D+(S�1����edmG�3:7�z
}\x[��������YD��-뛰����w�\�+}��8Rq�poK�͕�e{�ᆯ2_�i����K�2��mC�.�"'6O?]ܔ{&xs�o&b8�|Y��Fßu�5��aGY�;��]gb��56�k�e�S�ةZ��
ŇA�!t�6�=�����t!�C8G�^��cZ�G��:t�QA�R��{��ʈd1��U�"ƛ>�^���ARA��R�뽰���A��%gm!M������&��MGg��1vx��jܣ`lz���v����X-��`�i�2u�{�<w�p�ҧ^����QL�te�/ aT"�(4�ס���o�O�8ʳ�B{�}���6������wA���M]b%01���6+hEw�:_x�ۻХ�V��z���`�}@x#GgY��#�xdx�"���o���bʧ����	���l��-[��Q���RDL��/]?ob}H)�זX�H����p���n������}S��1ǝ+m����.�L���5�8����7��(Do�]D;�:_e�\<��oV�ϯ%�T2r��r�E\<��g��s5�ƶN�Zi�wB㵝,�Ε���nkR�wE�t�֚3���-��YY�y'��Xq�X�n�r�`��f��՜-�4y,
:�o�"EK� �T�{io������m��58R)k}�U�E�kH��c����dL��kiX��ҪCl]/+��=Y� �nR�E	�}�;��<�t����訍����D�M�9���5-��s:a���_S�߭T��{��G-~M��m�2�m�5@��$�F_��G����no)���ٓ���b����ۖ�$�8�u�B�v���{��,�笼�dҗ\�҄�*Nm���	������&T�|#V��%y݇l�{s�i��zJȲ�](7/T^���镂�,M�X�9���5����5:�[ߨ*#Սd�z$��9x��c*F����ˁ�-���wDI�{�=��͘�V�E�ߍp:���v9sjQZ����k�㙒��㥫�)5�_��O6/b'��f�n��+�^�M/~���S������T�����6P��7�,�k9�fR
��qo��
�=����vj��'��6�=����M
���/X�]k�7�s�	an���]�z�����G�Aj�#<ceM��W�J�����3��P[��=o����V�G�&),�����'P����6q(��n��F���6[�6z6�T�A;;��M[����V���4�R�N���R�ep]���)6S|s3�����Ʒ��i�;z���Vk_���f�m\^gn+���6ʖ�*{7q�#�ӻ(��W��%}�Z���)
ם�;{�Pt�絢13�_5v>�1�u��5G�n��UsǤ!�#�GP|n��X�P��̍�����~b�}�8?5�S���`Y�5�\����ʟptG�1ERF�5C���A���m�)�VBmӴ5��(���h󇧎��s�L�zn��(fe��rL��:��zcS����c��
�,`�������w^ݻ��#��zϸ�iWk��`�Q��:�F�t69�C��T�箼�ZD�Wu֕c�{9s/����	���U�]��ġ��؛NqnR	�ֈ5��a�Y�'_Xhy_�C|����S��d'V�B���a�F���M�\��O��`lv�����+�C���{�Ob�m{�s]L�g�ycSx��~FŞ�L�\�7��s����ce+�L���wdt���i^�%JP�<��3���{���{�&�,L�m�M�[Ӯ�*��Za����W�jE�S�91���!������>IY�����v�dd��}�R�*|��+�W�t���l�m�أ��c>�ozǫd��ҏ�&��	��VhL�n�^oCO�zQ~Ƃ͙h^M��t<���G�.^d��E�3-�Z�>.��{4�"��	h��\dI*2���uR�:,��ռZoD
������	-�y���fn������ĝ^�;i
�#��W�L�xF���c��s8��]a�7�Z��x�Ϻ5M�F�ea&.� ��[<ۺ��]�a^�]e/\�/wH�~�W�8��:�]6����`��+����%��63�3�v��/pH���.����]ǭN�r��e�7���[�2(�R`��C�e�뎶QW�Z8s�r���JkpC�n���_�uįi��LwObN]�7��3Ǉ���:�D�dOxU2�']u�*i��Hzo��F�SM��6��9��;��+�>]󼬊tY������&�j[RN�ufK.U�U���**�+�z1J�>{�i��^ҼK�ܹ�=�^S�v��{<��{ٝ>W=������J��7W;��R����
���Ia�z�2�l䍃�)�O^.."6A�D�l���"uJ��m���A�p�����m��mB't,3���֘�6k��x�i������e�����~w�����kR�f{��c�G
M�x���:�V���c��W��|L��>�;�{�*�8�Dq��}gSW�ˑ��A�wY/�3u�zr�Y"?_W�^T��C�	V���׈X>~Wb�����,�)2\y�����N�6Ӛ��ǫq�q��u��ݽ����%���^L�ҥ����ޗ��'kq��n���jȺ�����N00�������W��E�Q��U�B��s�m�T�Q���b�ǖ� ��+��B�x��Ѳ�|��ի�+�=��>�]�^�L�䎔�B����߿mc_��4�{��{��Ic�n���vڏ���6�RyޓCż�l�����{����q���ۜڒ�J��h�^֫�1�z.��F=�
|�ӃR�4u�>	�V^<1z����I�n�3��b��q�����Y�ݵ�[k�Ƿ������&�F&��ը�&ܽ�Ѻ�8�
U}B�|aCE�6P|���m�����&m�`���cE�x9K{�of�����
\�.K�
��]���6.���L�Q��-e,� v;�����
ą�e�I�7z	r�7��Żb�e�B'�k��_1��;zM�	oV<����Y�)<�g��:k:��㔩e�}&�&%H�x,Ha��Y=�B����/(��~�t���w^TƯ�N�8�	9R.�ҡ��b�JS9؍+ܔx���}퉍5�E[i���	��W�L�Pd��c�P���"��;�=�e��]J<m�J��������:�Oj�r�i�哶Qz�l�7Y�$��r�n�|4��q��9������sz�^�nt&��2�g/���i����]
�F!�i?y���r�7[4�Cd��r��}��\�B���"日\p�ܡ7e����Or�M̰�mЇtZqQ�[����.�i�BP�	��̹�M�}t���ur�[;����Fd[K���R,N\�'�z���-��	���g��r��v��Ab�gWJmf>B�8�\;N-��B��\���k�tSF ��<tj;�Čˡ���FM�]��X�Wv�fX�������t�FEJ"`�y1��ت�L*��.)��gh�XCO.JJ�\��x��7�$9���`g�j�&~㶦`͚v����A=�}�|��}�0�_��KV�ڃ��;��ie�Z��[Z޵��� �#K�R���B�T)��uٷ���1|�8'����Uv��[�墌w
���F�z�,ٙ�WVq�Ѧ�ޥ�8�^\�5�b-ȑ�5L�k'4_YL���&�v���
LJ�s/d���k-��jt1kL<�z',L��QRo=��ߜ��}xy���TF1���� �QE/T�Xab�EU��,�֢֭��E���+�h�mb��-#J(""(* ��Օ+YFҕ0�m�bGmRKe���,P��U��"H�P��Z�T��Q���E-��P�*�R��x�"�K�6�s^�r֥7+v�
���Oa�d���`]98cޘ�I'ZxT��H�\�&+�ŹI�kʑ��k�E�[.���v&*z�̗����@�����z_o(��̐۬��%ʖ�g�)�!&�gu��y�Y�+��c��u�^uV�8J{n�2|��PU{��<掖Ǉ"3-|3�N7S%�W3>N�x��)X����v+���Ǖ2�����{����C�1g_y�e�΅;{�W��֛Xf�rX�^lU}�����#Wᡔ��]��tؽu�)#a�\��Ü��o�Ϙ�����Or�)��'W�h!8+��2��6Y���]�5��z^������Ko��rJ�58�hj�Fmr�j������v�P=���#�Z��� �'-�s�Ǌa�/��v�����Y	>��\�:n&��YCu�궻kV�!I�v2<�Ve�nD�����8�J))��e�lm�����n�H���5 +hA�߼'W��)zf�EI����PO�\�3��$����v,�L�b�>��De���\ݱ�>r��O�I��1���߉ua���7o��9�dM+������QU�>TH����!��̓��Xk�C/�����·��V����[�ޱ����|�0�l�;!;tE�c͛�$�u���htX���]��e⺅��[��=�D՛˔kyi�n�6�;�SQ;MCa(�RU��^/�a��s�yS����:{�9�n����Dꢇ4�ҫ]�ֱe�+\C���� �;|��OMQ&+��vz�*�f�^�a�F����]H�����QN<g�x6yE�+����\���b8[���瀞D�-�(՞�m]a�����i{�F���d~��F�pF�_f[����Uc)S�9ٲ)� ^:C��E���`�o �
�}�[��lKы{� ||+"���?z��74�����kw��粵{�`��S�s:�{No���])�dP�;����:{)�W���H�n���L�BGˍEW��#�/�f*�k���l�K���0��TR1G������g�R�#h�Ը������F7m��2^l��,��Qޯi���Q%�nfsr`��mVc��{Xc�f�ӗ�v�$�>�=�	���c�;�닳����F���ʺ]�R������[Y9�*���p�x��<%�3l�����FW���^�Zɗ�̋Ƕt��Wi;sꀊ��~�J��Rozn��N���ã��������G�w�j��-���q��3�T����5��� ��;�2�_Pu[S�6�]�d>��Ԇ
����eH�J�=ޭ�nX&��m��
���� ��Ӭ��z�����d/��]���5�/ԗ(�Ļ�(����%i��<K�^3ɨ�.TK�G���{�g 䕋Z�48����R�˧�r*��m��ǚ�5�˽��΍ؼ���>V*K�ѣ���T5��Ne_F%��Ԛb��(>�<:���sN�q�#�j}]�o~r>��1@�	c\��{�Q���Q�\���n�w!Dx��9���ۯl^��LĪ!���#����Ӷ%Z�(=Iޡ���`�x�j��&����+���3��M�����5|�Pڷ&�v�"��M��1���O2���+C����<V�EW�G�P͏*�ƦF�Y�O8�=nϗ�wy�y(B踅��G5WT[��'z����Lr�#�
�ڭ�Ȟ`�9�L<v��9�etR?���F�l�r��4t�L���#��n�Ȣ�ލ�E�2��TL��CM�>J�b�`x�������JB�u��3���W��*�f4�����	�;���_�y�]X"oI���z;����S��y�~��� �����Kݝ��v��F5*#�]ח`k���<s߉ǹe�Mɩ
#py�zps3���I��O@Cn�ע�|��[scs S�Z�r�ƺKy����s�-\M���r�A�]hV8�.�I�~k3^���J�[]E�6��aw]�h�{���4��0yʙ�� L{�Μޤ��C,�\R3�9[��u3+[�\0愶�<y8
�Imk.��=��EY7�`���ʼ3d���`����6
b�*��e��ul^�m���ų�3:�5f�����Y�O2��r��m̂�Iţ�h��f��z7��Ǡ��+������8���D�Rq�K�,e];�)�{�*C�c՛���fM���G��PT*]��d@��w��Q�󴦺z���o�uM�_b~�v��=��ʛk]��}�!��ƺ�V㙖�#�����m�����g{��&̿=�W���8M�5�6�v�mٴ�yf>�?6��m��J��qTَ�Q�mR�+5$*���Զ��7R
�=�����2�n��@��A!|gB�V���v�H���-�+�Â��ޗ���|�,����0ȇ@���A�੪��k�$]p�C%�;�:���.���DVDz��G-k�U函����h;w��~�{��,�*7�雕|��m���slJ��kbR�X�{�9���ZvXE�����n�xL�jvc��]"����B'C�/����{��h��S�(vǓ�.��tVW@T�}�6����H,a�k1V
���M�&�g��M��u>��Wa��iW�׊�T�d�����Y�Q�x����j�ErM�1������~��ˍ3���x|����v������a�핞C�{��ad�Y���L0�wk�,"���W�����=C�r��G�v�;�/��b�U�1��kM	�c�;���{/3\N�~c=��w��&5c��u��E���(��=�W���Q��LඬG�;|u�����aϬ�ϓI}�Et�ޱ�lIH3���g'E�f)��q�9�kT�ڄ߆�oĹ�=,`�sU���5�I����uYh:�Q���g��
��1g�}�P�.��f��^i���Z��xw{is����B�z�dd�{5E��}�ea��f��9��}m-��fe�ͷ%
 ֫��.� �e�v���u�у٠���S��b�M�sa{�����a��L����P��n�/�iY�`���O�2����Я�/I��\v�X�T�8�����U���o=�vR�$L�Gʐ��蠣������9>1ߦd��������o1;^�u�V)��ׯ&K��/����Wc�W#}�ov8� B�A�T�5�t���6�1�&n��q���������l��^��c��pl7;,Do�Ú���3�^�^�`�ʼS��Vˌ���l�Q��)�v]���ٙʧ�$�C�$�����{���{��7��/&{��.��X��> �1g3P8��fW]�駝ԅ\]�h.���Gi�n�.+�;�J�3��]��a�P�cbޙ��c;��g.+���ڱd�Nu��K��0�w��Y�W���ƛ<�ՁljnbO��n����񻹔�}Ѫ>�)󻷆�ڱQVӵ�qM>�/�L䦙���17$$�]�ը/V|�-V��3eZ)̏-`�U�9��	�q1�a;2����G�[lV��vL[ Ց,�#C���)�%�AwU��5�9�A>[7w�����,��UX�1�̽�W`��|d �$�K��L
n�ӌ�*�ó/2�PE�w��Ó�$>F���ґ�U�ߪ��wieLr�-^̽*+XG$wlCSx�Н�����oh�[���U���oiYjLδ���S�75�Z��wH��>�MԪ��|GPIˬ˄;\�&̬I����C���
;,e*�og�ɒ��xbY�ڮ�yV;3R��oqQ�̭���&+���*�[�ܻ:��S�u��k"0�/p�:�5�V���n������1KG~hq�s�%�T�������H.ik�h�}�{F��.Q��meu���rd4jV�݂�E�"�جvd�{��e�]n"z��T��(�fe�vW{/�wB"/d�j�˸�In���J�1��m�q�u��١�lX5c˛(rZ݀�q}��k�g޶�,��4��aZ��b";
�����}���S:25�����	��xWmҼ#k�u�^KU��sfΨڧ�ʺ�j�������]JMX�Xv����oS��4�%W�Lՙ�#}x�>�OR��i��8��}.�v�f�ē��5ΫU/��)���m+�ہӵ�y�ؗ&��©>o	�l�s�w��Y�8�**����Z�26��֦%eB1P-�Q ��Xڰ�Y*���[j-A�2�Fbb*)P�P*T�+V��c`bKl���QVE+m�UB�T-"��3*�H��9`�,D����
9I�9jT*()+
�U`Q(�Q�Ŭm�J*�ʎ\ʵX��E����@�|R��=�B����Eh�͵a��"i^��赔��ǉN涭m�Z���aU}�
������%C�<W�f^�7�RC�a9�}y��c���<"yq�w��xz*h��~�0�ƈ�z���L�*V5�K|'U�9���&\��K:}��[�^H�U{�j���q�{vf��o�VF��M����Ų��c�o��V�l�2�E��ԪM�l��w'�v)���I���?nt�;�M{Nq��lR����}��|Zߣ�W[���wC%n���^�.�+�l��؜o�]��'49�|o�r��t��ܾ�9���Ez�]֟����Cį<�=���
P#][� ��J�y�Xz���H��}ٖۙ	�Rv�s����y�dn,�t�6k����0Н��oX�̖�2d��ч��$�e:Y>g�(w�p��-��H����+��o����>�v��))<g����55=3/��䳤`.1��K.7+�׸ا|v[��b'gz��1Gԛͧ�:p�'E����׷%P�2>�ٖ���MHy��i�){A�:�5l�h�/���ȴ*lW�8+��8�������[ԛ�ɻX8���_����㶒�!ھ[e�ݸ1z��ٜ�l�h���w)_v��9�śj;͕ց�W��A�5&RF�Kcv��h��÷aֳ��R�nYy��{�C���Ʋ��w��u����h�������DJm�4��yos�H����g,�����&]���o�{�u~��3-ؓ��V��������t�y׭�Ix���$��	�it�.A�A�4�`�ڍ�u�M���_����x��ԥ�]ŧ�\�+�a����mh�[�Yng\T�e�v�u�Wo�xP�=�l{�$�QRر>j�j��᧣�擬��yJ9j,RΩ'�щC�+�MU�c���������ŧ��NE�����,Q���4���P�rG�v章�=�����Pg ��K1�nrUO\��zD,��Hy��E\��>~���i��cK���]Nj]�M����
�*e�̽i�vՃ��1�U��,��Nq�X�bEXw�y�n��A�N�p&r�4��ٍ뱈Z�UK�-��4q�Q��F��IJnCg��ub4����~a�'��=��$SfE��	IeN^��r=��ve�o��=��^� j�c3ކ�ǎR���-����A�sf��۾v*wvq��u�	#t��1���d��}]~��:b�b�r�s>E��Րi�E����\0j7��i�/��T�{.a�@��j$�-��׮�o�&� ��w�c�-D{;u����Jz�8)t��=C�kM����Ɔz�=W�&���n��Gm�Zy�Q�t�%�}2QV=�o]�Z�0ZDx��Ž��!t��]��Mͤ�/\ޙ/&���\�,n��|���VT��A�s˼�EW'`�Uu�±d��q��h`���-�U�w��QN0egR36t�J���+�|�W���7m�Wm����[7�F�&�~�4����j�&�by�����e������Q������#m��m�׻���}���C{ףʡ��G�dY%�:�l,ϦAv�����-��[��ՉΏz�}�	C���@�3E]�F��r��w�&[��m��ɝ+�=�ݘ��%x���{+7��G`�G��M���9��V�#+7�1y7��x�u�2,���Y7n�Il�a��:���}aُ	p�7&�E���6wQt#ViU���OI����]�A��5������wZo��<ۨ����82={t�ے�ù�5>��ls���8��hhԡ|����X]��9j���v)�ل{�;n�]ݗ˅��y����]7�p��SY~#8p�WC5�y���w��L�d�\�_����9�Ч�KQ�����<k�;�ñ3�Lz�0׮��%�zs'�b��z�����}���uF�i.����agR���*<�H��	��Fؾ��k+�\��-;[�w����]�&[{:�#ct8��i̻{��ҜT�i\sn��w��ݍ���Oi�NjI��>nWb��A�n��ܩ6�����>���}����)/4�]����~tP�\mnu�L⃂��nW9���>�s*܏����޲k�u��˼�ˇ�_�~������B�~����W��.���oq���ޟI�]���f=��iJ���b���Z};x��|�|��w���֡٫�����������m_9Z���)�i��q�8�S9��,}���W�yo�R�I�c*�K�	���=�9j��f��]�&�>��ᔈ�|����:�1�Z�=H�.�껪=[,�4^X�'P����N[���<�����n��#4�Z֫/D�|��rލ��tζ�WN]J���ԣ���+�j�qĭw[�2!��NKP�����v*vS���w��V6��s�e��
T\�~�.�nF�{����}����O3�F�>��R��d�Z�L�o�v��1چ�f�8�ɝ���q�;�	�����^jSNt�c���@�O5�Ξ������c�������c!Ն�f+���uW��+�yTYN�?U�I��ͻ�F��n2��I`�˽Waǒ���������	��ޠT��\1�Ţ�fb;��[����b}������7X��?{���O%{��4~�#�M�,�fYa���}j��\jt��3k;3u[Xq�`�]�۩Y��&�=g�\���d���O��h�YۺS��95�`���|;vX�x���ܙkw������ҫ��G)S���QjK\��}C!�7%MD�vBg�Gf��JwF^F���c�}Z��s�K�A���Z��7�&�C��#�B��y���d�8Z��'���F¤.w�����n�[�:�R�z[�!�~����B�8}�[Ndm��W�R`���2oɊv�!�}������ٖϾ#���`�X�F3�~S��xR��z�*�ߦ+����W�m���6$�wɪm����o»�wEVL'e�Y��hv��'ZO@@�zGO��4}c��؞6=#rX�@��-u��Wr�I��m��*n��83�z�#*����:O2rJW��)�#��}��,�8)u�uv����1��:�@Bԍ�p=HU�|�O�G5��z��'��Hs�݆h�#I��}�ݙ�bLr�+���ϟ����lwn׫��-���WS�F��;�rr��G�/��A,R#�m"��S�{Y4�����?R��SN��u�IU�^�@�����`�jOdC3�g���F�����羆��.9ǷS�[K�c6Wf��*v��%�&�W5(��Z�s{����q�Z��q���>������S�j�*�A�	1���� ~��K<�H��O��~���C0��Jg��k�;�m�J��\gL@�
�T(r���@:?{C�w�$�h,���'ɀH����/��O��{����p��w�C�\9�}Z>�i�N�߳���:��0�ͯ!�GG��N'\tk�$	?�'���y������(s�$$@�@��! B�!��"�ɇ��ӣ��C����O��?s���}��~���6��O��$@��������z
��	�~b>��1L���>^�q#ܟ�^q ��X�̈s��D�?�����ῠI���X�z|a���?<���` ~���C�t�	������~=pt��������$@���������}3�|����I��_4Y�d���};����'�~���?G��S���1�A�|}��@�!����d�g���O�>��>�pe���gd�P���ߏ�}��t?�������ٿ��O���}���G�~��(}�A����P����N�����dD@�$������@����D������B�������4��B��#��s�d !�O�*�}&
O�;'��!��N,��}���vxxD�Ա?[́�1�$�~�f-��th�]�<��H z`~?a�~�@>�}�	5���C���3���$����C���������C�O��������!���|��?���!�Ϧ�_W��?���` }��k�������C�H����Mx=��'�<�l���>$��f���N4�đ�?\�顈���ߊ���������<C�����'T�w�}'��	>��d������灇i��*}�C�z��{x�x�?��jIC�C��dB@���'�����S����u���A! B�'�}��9o��~�NC���v$㬳���)'�Ԡ{!�����]��BAk\�