BZh91AY&SY|!�;�_�py����������  `���_n     @   
 
���U(�� T�AJ�T��V����EQTg (  �� ���>�w���wc��v��J��3��n�'��7׺���4���wx�u�:�Ѷ^Ǻ��xwy��j�{]w���/�� >�Ŋ��k�)�eխ�����m��pջ�^��{����m�|��/�ݶ�^�]��{�{�a�q����;�\{0����}Q��wͽ�i�:�7��7�Z�l7x;�u�z�)��y��_M_��Z�۸��^�������G!�k��%} �w��n�����}wozg���{���M���{�_{������/-�7<�;�^����z0��
>�c1|�f�����;ǻz������]zm������swx^.��s����1�v��]s@    � ����@
  �@iR��&�L� i�� ��A��R�i�4�4h�@h���A)��&*�0& F !�  &�)Ub4�!�	�M4  "*��1M0L�i����$�z)�x�*$������� �@�4�ɀ>����}2�DJ�A��>��$2O ��#��O��H$tH�" )� ����[�B����(0�?������UQ"���f3-�����@	�K"z�UUB�r�hI$ ���g�I��G����?1�~Z�K�wL��ݕ�<��~�$ඍĴc�	�����:�[%�]t���tnMA���.�gL�lմ�p�앞�lI+E�Kp�ԵޥGX#X݁�"���K��d�n��Y��ILn@# e�&�U0r!�]��7F��`]��=~6HTHB�dSLcm��%���F�6�ݓT�V��C%��;�tL\���At�]XK�h;�k�d��N	�)�:�XN�l�d�&��4��w��zA,�yd�xI�d�4HB!�tI�ZMb�p�,�a��f���Tfj��M�)�p_�H/�I8�Đ���Δ���6��m��f�X���F��4f����b��M�E�qM'6һIT��!�%�`�:oK����KG,�M�l���ˢR��rS'Y%���I=E1)���ȦE2��A�%�Q�f�Jl�e-8��%�)YV`�0�4���SD�+�EZ2�S���ɚ.�4ɦ��IՕ6M�8P���K0�KM,J���゙5D��l���Y5�K����3L�g1��n�Ƃ�Ò��xUY,��Zg�R��8�-��M&�RI�X$<!�M��U�V��1".ʉ2짆��8L��M��V�8 6K6�',�I���ek7��PM����"�"�"�!�^zT�3p��wY���bV�,z��*r�h�-RU�D$�
VU�0�4��"�BbH�H�Fm�Oe���f�g\��%�Ѧ�:M�S��R�	4Y-��IN�-IZ�i'�,�S��RnyY)�&�̻��K�����embC*q#u����b���	u�N;��4��R�j�]j���uv�4��C�gL�5Ff�)��-�;�d礜E�K�A8Δ���6��m��V�T�S�)�Lњ7e�ŇrU2m��Nm�v��IP,P��0d�/N����Q,� �J��їe<8.˲��$�:Kԓ�V"�:\2�)�dS*���]���I�R�&Rg���PM��Y~�Ɛ��Yd�Eb1h�FCF\p�9!�pI�&�%4��*l�����!�,�a2��X��%n
	4t2e��Z����"�0�!�z^�U����7f�벖^�$�YJZaaJ����$�$�SGI�j�@�	zSgD�+o$��nʻ2짆��8`�Id�8Mf�p<*p�LZ��IƤ�
Z|���u������.��3K2�^��\��6]l�e��nΌòp=;4�=)�l�)lBY��)Y��X�$i2d0H�H�E�]�R)�z[:�g\��%낚6�Z��V��)k��*��I���SE��4�4Tn$�qIS��AVK�MQ�F�IV�%�J��:S����6�,�'
U&�E�c<�N@,Θ
�M�ĽJޔōF�#&�A���Ѡ��b(���� �$�L���Ķ�C)
`��`h�h�����jX�WR@�'�jM2�!�D�dO�H&R	�Q�S�U���"�,�M�K�u�t< �$�uiS�*�T�L�0�a��d�RU�,�K�V��)�r�~,^���)�x��4]�d��IM"�]JN��RMQ^~���F�pT22K����E!lY���4S�&�m&��C�L���L�O��ȏ&�!2Av�<)���V���c*��s̒Ʋ2N����U�+:�L�0�~f4{(�$�!ـ�/��1�R���������c]�1�[$Ț �d�ui;�h:iJey�C��JB��	�P.�%OJcvR�E1{i[���zV�}m%z��u)1Td14m͕���2�d�I��2K�U��S�۰X�(�h��,7�PsI8��t	s��I�T�C"C"<�A2�NҀ�-�:��X������$�,=;�(�������	d�TN�%�"� �@T��`[��Da`����b�!��y��0_��`��`�������l1�Wg&�w�����c7��uW�A^ZL�C��M���%䂆�,F�L�O�]�����U�tU�&�^a��#}���*�t�E��a�����	[��X�6�)�V��!`9��j*��K*���$¢��~̃I8 ��b%""�&���X�Lhv[��9��QHF`�/�&5&��HdHdG�H&R	�U/
b��Z�ј��eP�$�,=2����E�b�@"%��rMk�c�&À��@@�*@b�'&�d2d�XA��#�&}���6Eb},�l�c4'Y5�*�Li��KD���A:��S�=�š��w��z4Q/$0?$�h���h\��[ZٶV�]�1����vϝ��l^0X�X�dH��,.6Ǩ&�4N�,cm��~,5�ć ��-�40d5�����1��}2����ʳ|30#YS�d����`O�-7*'���K��v�|#���'�'?�O�㡫_�����1��N%�S�oq��ҕn(����}��1xx?i���Q�Zj�}����9yb;?�JA�VN�� �I����eB����f-���A��g�7"b�S)���2���T��d n�*�a�B�Od���Λ��f�3��V�+����=����Y�BFDr�K�f�몪�N�rmD��-T.ㆥ��~ ���q�{�A<�T�nы�ӏ�;��ۉ��	u��@8x�t���R�و�SE�E��JLţ�pH���ƽe��UF�r���s/i�
Ic����o"k��0�g�Ȩ�>Qc��i�ʍyTph�[B�;�q��j���6n�Yr����a�*rftS^����1�	�q0	0�K�Y�^�c�����@weaUV�]q�F����:�����75"�̐Z;7���y�o���|;{����8v�����[����b��w�y�h������;\�Ywob��#�f"�ĦD�s�6�]Y$�؈��ˣ��i�����C٧��]�B��W�F�d|��<}f�m�X��5j,��3S�3f	2�/��6�¬����Y�gbD�
�n芽��q�A8 �d+#��,�g�N��Vȩ"�a���˸n,Fc���Y�4/�Q3$�x��T���H8V�A��b:�.���AE�IJ�a�T	���j�N��C<w/��	�&�o"�\����Yaە�$s$ϖQFTv�a��>nʵ�`�5���謨�lt\	�4��ĨeN\e������ގ��P�~ܗ|�++��ط��,�Q�A�J���ZHF�䭦p;)�M���hA3�#9' �Me�C U��N\�q�R��0l�A;Տ��z'����wU���SR!AɑYS�/n&�i>ꄦH�f�l�5��1qUPs��[U��$�d�S"`�"LM1��6�f�*��2�9�Iyc7kb)�&��:�r2"��d�zf�0���ʣt�W@�5R�w:*�DJ0cH�TqEP���p4D���&���D16�l�tk�FN���ދd!�3�',�M VuD�"&7V8���;�9� Iú��,�PW%Yr��)TDݘ��a�ݻCnm\���S$�]Y�"b�vf����re�N{�U��UBB_Ed��3gf��?�����='u��̛6�B�*�����xlŐYe+�5g'*�duT�ƚ�SPI�:�l�,�ȱ	n�q+��Y�1��2�պ����F;�+/h�*��w3��1��}$���0�.g>D@�-����rEA���˘�8�!�p��Xjf��+Hin+�t���o�.b&"Zٕ[U���nY��{���w��y�/<�-�"!y���-��/*�M2r"YBЂ))An�:s0��sݒ�vx�;���.)5J ���o�]��W�ْ��-��g����h��j�d�!��f���C��DH�/"�!u���x�|�ж�p�W�$Ƚ�X�l�ut��F��C'���!�hc�������,�����3W�a��(7���υ��\�m̄�|�.on�Z	j�Jb#b�P��[jMKȰ�\�ȃ�l�p��ե�E�s8hAثҧb�^$j�ẉʍv�;�u8�J�i���[�ˋ��&�ᑘsL��ɷD"�$b��ΖkZٸ���b~gέ�f�n�I�z�N��?OgD���jN��LZG��6�f��Bl����`)��6`��<v�9e�e;zJ�k��͔��eƥ;��ߟOf�/݋�����MV�a+��G[��Lk�a�{{�g��"W�y)0�O���lN��'�Nl���b���H�A5�VF��.26n�8۪���F��5d��qc,+���o������K�L�,��=���[;k�o_����\;����oF�@�ڶ_�����Z�A�l�%\P��N��(���
*F�4���H��J���7]	o@��E��s��J��z��殴ф`�x�ԅ�O*,�E��0!Y���SS5���;-f�{U�^Q�X��&ט�8]`W2.��R)ى�QMf݆�qfq��UN*)^O�#ƌ3'eX͕6��&�wCK��'�Ih����o����Q�3�Wf�,������xr��C����uZ!�*U��"���s���j͚��-��S1nrW	I�|r���E�Y��e뿈7���~�W~�x@^�Յ�̌��ߺ����Z��;*�eJ�鎇0h��VUeQ�o��fu�]�j�g&Kh��.�Rᗽ;pe���(r�j��d	��|3ͬ]�_�YZ���ܳ����b��e�
����_�߻��yֶ�3$$aW�1vB��ղU��)!Q�VQ"�1��wj��ǘR��x�BE���&ʴ�9���Q3T�6Ɋ R�Z�uuUI2\�,3B(ҏw��w����"��{�7��9޵���c�}���
A�&.��32?�:�ɷ���$E�{%�z��(�*���m��J�D֞����3�w�<�����rQL���m��I�Yyr`��t�tޭ�n���A:u��%ȗ���	
���>M|>��3)�>�˓��>$��@�ə���ɧ��N��<[TZ#�����WRѥț�V��e�W��1�1���*c�,��*-i�8�Elu�K+�v:�Ee?�ʌ�e�Q�H�j�E-B!TR�2�r+E9�:�x��amN���zBb��+.ʚ���k�%�l�Y�EkU�*,�����М77�ŏ��'OU|�D� �[/��a� O*�e�U!C�u\�y5cl�E87-����w{(��D�b��Q�-�Ud��(5�#X���v�X�mʥ�%Q��:?�V-���.�7�,����N�MK�9��
)y(Tx�K[5�l�Vږ*�_kפWc�X� �Oޓ���Y��������KPn7������:��t<�o��p�k��sZ��`�B���L1BN1^X��N��V�xּ�knD8�$q1":�,��<+�����F58>8dN֬=��5f-�j�LMn8�nd䔶6���PL(�6�1W�[��QXBE8���t�`?�}ΖQ
[ji��MH�|�9r�IM��K��/�%���'E$D���eϗʫӤ���r�O���)*���[��+Ӽ����JDM��5"I���v�9����w9��#$&�_���ɂ��f�6�e���^��櫏\i��[���U:�ϥ�d��')d�K��T^��-Ҫ���t��#�k�i�Q��'�qڢ�
v�5�F�Bb��YA�7�7��u���Lf,�[�ڤ�PW�Ɋ,I˗:����2MnK���ʪ9��V��&�U�d�o3mƦ; v��&Xd�fV6��F�2�d�b(�"׷�����p�����H���DT�<��I>{D�G~���_�#�O����|�H@����k��A�F���ն�m�m�-���۶�m�ް�m����n�n[nm�m��m�m6�om�������m�޲�m�m�m6�v�n���[m�m���G� �x>����|U[�m����m�i��n�p�-���۶�m�ް�-�m�m�M�-���6�6�v�m��l��t�r6�om�ݶ��ݭ�[����m�n�{� 	TD�Q@ֳ�w���{���;�������m�i��v�r[n[m�m�m�m��m�e��vۆ�n�n[m�m�m�m���m�nm�m�l6�m�z�m����ݍm�m��m���  � �2�6�v�m���m�޲�m����m�nn]6��d��m��m����m�i��vۆ�r�n�m����m�-���m��m�n��7wu�m�m6�o��=��H����xwr�n[m�m6�o-��z�m���[m���m�m�fm����m�a�m�oYm����m�M�-��m�~m�ݶᶛm��6�{{�ww[x[�ۆ�n}�H x� '��u���vۆ�r�n�nm�l��m���oYm����d�m�m��m�l��m���M�x۶�6�6�v��m���ۆ�n�-��sF����n[m̐� �O��|O���EU$�"��>��_� �?��E?��O�W�?��M�6m�m�n��n�m���m��m�V͛6m�xv𧇇o�m���6�^���޻m�lٳj���6ۦ�t۶�x��������N�m�������|���6���m�i��b�ٳfͫ�m;m�Ǯ�v�m6�lٳg��V�i��m�g��Z`?��{�I#M�o�y�����?jq��,rep�Wo��YH�܊�H����>D�a!��Q�YT*��Z!��p�ܒ|�Yύ�4e�7Q���}r�1������F��t�a�;�r?
�����Ґpd�ñ�Q�3�����슔9��T�j��@E���lU��ShO���Ӓ��ʬ�����A$"����`:�w+r֘F)�f\CM8m�P�����o��+}m�"�����P��	u�I=��k��n�_{�5�6Ѣ�j9KX�Ьu؉[R�N|�G�%;�7x8��]i����JĞN���rNA4VD[}s^٭��mm���BLP=5@�
ֱ����'$����U
��SVQ����X�KTb��*��A5�Z���l�Ŕ�ۉ�aJ�����ku��Ό�%p {Ǹ�wT�����H }�����c7�-x$�=��33�;�]���=��9U\7���^s��s��������;�L��0 ���==(���~ޕ���H��y*�V5xEAA��*��L���̌��d2!D��9��9,*b�͘�h�4��bg�M;z5�����UQߕY �l50+�E0�<�ʙ��U�!��N$��M'��s4��Ru4S�7EV
UK��V�cm��6�[h�'r�|���=�#��4�x����BQ�s*��,-�� ��&����M�x��)=KL8�^�jRe-�I��[�Ű���d��r��!�
ц�����!p��e��;Y��i|��@�"'D!�,��2:�i�a%��{�Ӧ��k0���Fa�L��.��l�&&VZYl��'D)UUX*�V��QPɎ'ga�nЊ���M��0mU�	pܓH�f�j���aə�Q�eQ�����ư�o�mU���ڪ�z�Ǐ��9��w%���KN��JU<dX�R�T�,���č屍�8-�ĤޓI�LL�;���a�ٖ�\,�:)2D��ݹp�Wq��5:���M0�UW��&�k5f8���FH���m�iOj�V ���E����bm֘eN5���(��N�*Q�(�D�
�l*��LO+��TTNJ��Ȩ����L H��8�C�$U)'�u"����A`'=*bzjp�0L��P�Z*��h�<[��i�C&@�t��/z֬��J�y�X��`�ۀ ��(�1��;�;�i[�f�a��U�֘��Povu�8�ܬD�JN�m2tX����N��*�eCxH)l*�E*f�`��;9
����+iR�#$��ukBK2"��§���aa�B������w�S<�TV���6PPQ��"'sj��0Ό noD�XٙrZ@�;,�����6��ws�g���w�.v��	[9	ZS0т�(����fo7��n���2P�;��8�â�j<ju=���+��i��s���*>o��<̜c��qrrԖ�h�hq�����%��%$ ���*6!1�nb	g8���{>�qg���Sc��T�!}��>�-$ �M2 `Ҧ���+4�
�l��_SUʇ������ÿ<�����=)JR������i����AS���U.c"���"���iS��6B���e��K���ّ���m��ؠAK''nF�r�;5�1ש�A(�t]�`�,m�퀥�UT��6hY,�E9
�uV��
7��(���f\3
�s��7�j�MUR��o���\���@��襖U+��HX7K��6$���ü;��ʞa8�IÉ�BO4
u,*uh*R���,��=1�bK�J��ù&B�eM�N�Crz2���s���r�*1liqE�x�=�N'���	"U[UJ�9yyP �^#�1����6Xi=C�h��sP�\¨�(��.���)����NR�hQ>V��U�Ū��g��U��J�x�Vqq⸽����q\^׋�⸺_����&/f/�<(�Q��	�f�e#B#�W�Ux��8����<_�̟�g��S�|?	��x3C�>|��J+�xp�Q�<9=K�%xuġ��w�\�Z�CE����b,-�W��S��#�Ih��W<�:s/Lq�b�ʮ����M:{U;?D��=f��E'����x��^+����H�����)��y��)���)=�ځ���'n셊�ϧt�<���77��2��f���E�97G��<o^LLxr��MN
�Ҡ��`�ȥ!LI�9Fו���,��
��هU~�ܽ�\m�t�P"Ȣ��n0^��%�	S��9��{�����vǯ�1:p�)�R��UL�|�	S�{�wuT����%H��wUL���b<{�wuT������˻��g�o.P�wtwUT��Ep� ���`�-|	�ŖYe���UEQES$J	��&{*l`Rv+<�(�٘NĄy
 s
 lڠ���J�kT�LI5fN��%�HW�"��ﾱH���id�m#�"�G�ɹ*�U�N`�L��X��������*���S�&؍t���`ቦn:�-n6�oĠv�*�X��2���f���0C�3�QQ��.�B��WZ|z��H��J���`��i
w>�M��vW��M4�Ph�QEP���Z���v�(�ʵ���V���R:�a �	���䵙d���T���L�fhX��K#�I�H:�,|�BiV�": ����-2�bLw��)lR��V�g�TJ��$S�	C��m�N���{l��
e HCI1}
��T��`�-z	�ŖR����<�S�_�T[�o�I�%��B��7%���PF:�qV�����Q �fG$PTfWn�0��Y[�!�w�>(����j�J)�EJd$����tr�E]�K)��c2�+-��'��i���-4���B�4R>`�%�ۂƢR�49`�R&S%8�	7T̙r��D�fc1y�Rz'�l����8���"&X� �bx��G�E�5�V֣��j�O.0�`��͍YM\QV#���Ś�3#س(�G��e嫨�d��Sg����_�~xҔ�8&���W�5�P�htXHJ�j���Q�K�q��bv����|e;��!":�9���&�ܒBv�iN@8�)�tiM�K�[� �՛��&R�qH) �Dqt�F`�<g���u��`��20�"�=9@]��I� i"wƟ*��7�r4u���#��A;i0e-�P��Ob2)�t�ZVb���~i��i����F袊(�c\�0�
�,���SĀTG150z��i#Q�=KqΉ!	v��6Ĥ�C�G��b�*�'R	 ��ӣ����h�����T��蹼X�*���^JP�aL=�=2E�m��4�պJÄ�Y���)��;���z#����i��#�e�0�{ ���S�Q!D�ò��)�K#��h�#�M"�(O����0�@�k�����͙�Z$�).��AGd�j� �5�&��Ӟd�SI������P8)\p��0��֪�JkP��x��1�
��C�MF�4�~��<�y�ԥ<v�4�i�<<)JR�<<��d���1����W ��1�,�1��V��Qe��u[��q�2(�*87*��/x�8	��h�*�%�R��NT�&E,��JV�P�>=P�*�yLgǦ䝙���2�g��ŏ_�q�q�Q&ޭ�L��[��m�܁��#�����r����㴴۔���_p����Ǭ��\"�s�]�IX�J�a��OUUP��C�p�`�(4�i��m�M4�L~��2����4����FL�6�������g��o��I%o q�%9L'�KH���B�;=CA�OWJt5���	�� k��Q[ݔ`k�ur��T�]�6�i�܈x��>�>���>�T�>�ԵCT��4y2)��a�+Lvc��1�;���*��dP��R
*8b�*N=�p�K2��篍`
c���l�aY��ׯR'��٠=���%_+	�uX��v(�m����C�ޘ&@ץM�>��Q3	�za��	��߇��k!,�n���F����j�;�MF��+1Za�'��"S�,5t�����:�(S��P����6h4��Ĵ��|�?�I��~
�c�@��p�4TQG�
���14g'q
آ�cm�8��L�d&1�Zu��@4s�0�R"Ri.��(C�Ź��F�oҴ��S)`c�N&S,���T�.������:R%
<��Q�F|(�D|;�0��q�/�q\z�+������C�2?(��D~�G�<'�Ţ�Dv"m��1��/�������q�q]6�/�<^:c�L���S��؟�r|VO�|h��5��<�+�`�aH�H�AX"�Æ�Ah�;�L.�R��+�\�\i�4�^�W�p�m��s���8�-��<W<\�x�i��/W��x�c�qx�q|q������\�͚�-D,��vJKόR�*[��]F_������ �M���pV��a5�������F���{��~�,��(z�._�i��Uof��}�sry�Y�F���o�b���9k[B$|�殴w��[�6DeQ�������˙aHI�w�������÷j�<dW��3���TO�Fmq��r��C!B��A ��H|M��i�)ϥ�"q����y 7��r
�-P}�ۤL�xʚb
*�P����@�VX�6�./9�E5>��� ☝��ٹ~3�_{TS3���SRٿHV���AdҊf�j�ю�/֭f<Vq�E��(ժfLR������]|:Q�Ti��ɏ9	��U����Dc���T�W�e�uY�ي��)C���ʾ[|PL�j��>)�dj�Suѕe�i��;$*]M��-`��:�E|m �M�\����d����8(�j�1�K0�,W��+L+��QǷ��A�,��d9�*,�ee8�jJT4r��n����q�dm"<�.(�۶��&�����;����n��~]����uS<9�+�wOOu�L��Ȯ=����wSß"���컺�ܒg��;���wrI�8p!�z��DJ]���{�;��[)V��T�t�AX:��}x(�I���+kcv�A�(��bQ��-v�]���c��t��4ʬ��JRK�7K�Y����(�RA�����&71��Ⓧ�8*˕?,d���-1��5T�4L�f@��I��Kܷ�r�
��V��z�T�O`�D5��U�W��_��4�H�L�}=�,��d.:Ù��>���.,ZLlhj���jڪ�U5�n�^a�a��(1=;�AU�l<��O^�
�Lc�O�c�~}��_TT��Rv&Y�z�A�t��8�ӷl�l2�`���V@�y
��o2J��&��$$��������屮��J��:z�u��������ٹ��F��rx� O^&��a�i�ۑ�	P�b�s~���i��|AR��i�ck�d��1�֑o���4�����(���e��7� D�E�"I�y�%�v^�4��4���/~r�=���_���nq�P9\�m��Y��)��4V��%I%%�8m�]:���X|t�4�?XŢ��P���@o�����8/PL'
y�(�u�שO��T�QR�J����UK�'LCP��h2hJ���<<�{Ǹ{仼��}�kC��R	��V�aR����Sშ�0 �d�l,��1d�-��BA�	�&�뼂�m%@H�a���ڔ�p����g}G��&�� ��To����g��l��,��f��^�E���e��\6��;�w*�>&���Vf27�^*�w�حJ#~G"�)�!J"~
~:��_�В*��Wel6�nk���Zla.Hj�WXëg	�D����ٵ�m��#bɣ"���a�[�̰�d���c��U	d��sHRɫ��&�u-[bI��sK���i�cnR�l�n��Hv��PNd��9���YZ�(�4QP���-�2O`ճ,A0X�:�Kt�nI!�3 {A��۶��8k	���ƈd4ys�f�h��_݋�u	�fTQ�$��Z�?`�S�1,����갭4�;4�U��'>������JJ)���f���(�z����զL&Y@6$���H��}N���RPV4��eU��Kh%%��C�63�U���W�
�>'#��mĺ�,�>���A}��A��!���m���0]gh~v����j}���00榡O�
�Lc�M��i\�]F�H�����Pv�ഛ�P�*���C݁�7!��'�N�G���:� �n�L%�E��Z�r�o��y�*�-4�6�9g p3.�SB�l��ć�͐�A��1�v�0���3���N�q� f�y�7�Tw>�8CF�L�34h�d�ӊ´���j��w~��u��6c�f�\��Á7VLog�K���ZC.�\r5ǐʗ�WX�.�����vp�,�hz�m<OS@Zx�-�wf���R�m��Շ�n��Ĭ�N��Ä��pU6\�Hp��P��U�����x�v:tF���z�)`t�
R���<!�%�ӻm���J[�:6�L(������ˎg�2q��M�mj�If�\�JZ�)T���
"*r1��LatQH�����f8��i-�{�f��^�x:zX���0�wF��4������U�9=:=l�i����u(�N&F�&��}K�F���x�/N�B��i}}�:��l����p����j��z�juMV�<t�+���e���_U^pԻQ�;|vN&����j���2�B�i�w���>UT�@��w�ni��(�CP�+Ȫ�US@�^ �_�Lf� ���(��t��n�[bIZdH���i��@1� m�(���&r[��[��G��GL�;�xpE=1 �ϧ$�i��9G�8)�H��D|(��S�W��D�\���GÑ��=g�q\i�V����v��[W��Q���g�:(�xTA�����+c>����O<Z3�x�^��EpM	�Ԩ�Q�&����d����p/����������H�4�Ǭq�^2��\]�n1���=q�_���	���P�x8#��V�H<�nb�+�W������t�'r1I����ؠ�C���.�3UV`�{�59qwN�=�w'�.P����Mm�1��3�J������c�8m{;��"߭�!$�����Yۙ\�}s���S��]C~}�#<V�;t$��qdCܯH���Ց/�ٿ_debo�������wu�|��&{��{.��w$����컻�ܒg������wrI�������-=��=Ywuû�g�8ⰬV�Ui�W^S��~�[��i�7�p�䐩�u8�}3�M9N���|L{�R����I8��l�p�=��[�]�0F�h��Yd*�O{<mө�{Ci���Z�#i����9<��D+DhV��p�--m4VS	�&}��3Q�c��������N<V����<!�<7��`h��غ�RitM�IU�:w����=Kp'=;wVZRYE�7V��p��r�'�b��z;�'q��⌞w�y�;M���1�e=L��)�)ѼLNC3��}��X�9p�b�8#�����̍��{�F�m갬U�,ȉ��	���_�^l�F���[��S"�\b�Z�<��%����B� �gbx�5��Y���8:�4rQ��y�����ah���Ȍx1�_2EnG#M�:�'$ BZ�J��_+M��ӭ����heN�G
�,j[i%U7{$��<��_	(�}Ku:�2�5&��;%�Z�@txg^9w�,�6�Re��r2p�vx�0��Ԥ�2x�8r�'T����G�ؙxV@���.�%��7D��p�©2��m�L�Ԓ��q �3�J�>��$:a�ӥaX�:+G�'��Y-*�B��z\*s�m�RKK�n�/�MD��*��U�U^��C@R.�m��S�1�°��ᳪ��@��R��K76��F�nVDp�'�p��gxy�}-�N=�#��'�SԷ	�϶�S��h(:hJ�,�%�:vmwU����!�%�eEJ��ϩ&R������Zb��i�W󟷞�Z���O��e+�Xډ))t��8\9��t}����HIm�;����j:�Cm��Nx`;����58g����;�.z�:����;x�+��i�U�V�>��ȂW�W9Ը����F�c�eڴ�5�s�z�>�)M+L�O���i��;��jA�2�K��lZt��!��2��Oe����o�_ܪ��kUWV5V��%���)�ԡ�m��$c4�4��6��^�$��������_�BZ�/'�������!�I��vJ�����\��%$$���`ؙ�ⶫB8�UmJ"; 17,��Ӂd�ӊ�$���VT��j,�ug��X����a:�	�He)01�c���<��W^5�u:5Ҝ��C��I7�����UM4Z[��&Ҹ����$35!�a�Ð�(��I����>7
f��eCy�0��{D��~j�VQUJ^,�p��&���vD��������F�)N���� ���V���q��2����d}䝩*{�C��})=櫗WTVӍ��Y�Xs ���7<�^�EF"ߓ��֞n),箓p��$̄�㮲N�n�!8s-๜X�s��9�-�[am�UL�4n'%�X9g}r�3+~���h���aX��8P�5z�U-2MT=.>��70L'R��X,U�����SZ�����Ǒ�
=�I�=�q�ٖ��K[JX0��sp�ț4�=4;2��j���<M���=z�U�ie��Y���F���m���<�>t�!&�&O��Xd�	Bt0Y�(���1�����7i�4�Ǵ]��C�V��sʊ��a������j�=����ň��!���[8* �G�Lz���4�R�zh�R���L�t�tʤ���yi���<U��T��8�7
�� ������)��*�{.�!J�J�}����܈W�p6*��DТhQ࢏DG�D�|&J�Ԩ�D�/�c�88��+���8Q��GD��\��Q�z*xQ��؞����W��=;M�t��'�`~�+�+�xi_��g��Z<TG��|">�<d��Ʃ�84G�B�Ѱ�0���pJ?���
�z��Ҭ����x����������>aj����|��l�[�8_S�rV����^j��W�p�Z�q��8�^/P�������^Q2/�9Q{S)22��ƙpY[ʙ�ɻ�fۻ��߻��ȫ���U�׷E�ST�{�X3mTDI���֓w��٢�!��,���b�y��tǲ0�䪭��^=^k��n;oS�#ˮW��XE�OnvdފE�@�۝���"��T\zU��]������1\:\�I$�'lH���k�� !{���F^�����$Z�ǯo+�#A��TP�]����y��r��!�ڇΑQ�n�#�\�Ֆ�K��ȄT�izֺC��XR7a+�+z�+M7!��V���9yv��f6���7��n���\�)n�j�Y+�&,�ʜ�V5�Di3f�b�۱�N60��Z��jTJؚ���ARX��%j)-�s����~�J2o�MZQk����]X�|��^;�51� �Q���M�VMCV��3z��*�S39b�B�)ɪ�r51��JF�D��)�ɳ5n;��d�~�D%�V�Ty��J��1D��HJH!T&�+��]e��Ǒ����U�w|;�#�����.��wGOwwuV]���<����ꬻ���y=����~��s��}�q�aX�4�ǧ<�+$�ՠ۩�X-َ��±A��Gcu:�*�(�,���,00w1*�D�������yb)$��J��Q*����bɻ+#ȭ�IU�w���|��l����!�ݤh�L�d�*QN����UW����#R�=F�/���5�NK>f����������z����Qr��F#�;	 �����0&����=�<<z�+��O��?>~���G\*{093���d�g�������<�'��	���$!�&t��<8�� ���2�L�N2��{�*��꥙�ߴ��N�xP<�Cc��1���嘛�X�\T�Zt���5�5d%%������4�Z�����v�^��SN�!g�1^4��c����=E�g��$���S�Қ�e<4�$t4<N���Rf�����z��f&R�2�;?W��')h��"r�.��W"���x��Һ�L'��!D5q�>�;%,V�}2���B��v��"�)�l1�᎝��8���<�1�F`���^�]90��qc��5	RUIT{um(����Ξ���YH0�T,�k�CF#v�p�q�؞�-2�JC]LeÓ�D��1%UH�0�<}N>�m�y��#a����ܙ4��?4dy�~��H����ѷ�1������;�'yY�M�l�`����5�Y٣��m�#��r�0Yn
9jn�b�QD�2�(T�<��Vuvb��Ed��'FHH��jE�8��+ȟպ(	���Fq�$n䒹A���L�6dyJ���GQɻ��U��ϒX��>�Ǎ<.FL���ё��Pj�r9�͛����"d듒B�ש ���i�>�L�B�;U�x��V!L%��ۺ�	[񋴘N'WG��ڶ��y��?--4tx�b�p����:�?qv��U: ��ag���Mu0�e�������ެ�$l�����S{���	�@a&I�@�|KU�d���ےD�ud��!Rd�s�.�no�Lz�0,K��M���xz�h��k�aی1��U���|���X��cZ�U�
Or�bw.6����z*�A���k��j�Z�'ē�G���f�eDB���V�5�0�3p���<=�RgPߊX�Tu\�����@�2����_�z���f�ܒrSPǬ2�L��+����~s��an,}�]6ق	E�&a��G�P��ӷ.,�[�	C�j}��',8{�RT���h�Cg��17	��VV��6�(v>{(��sG��Ӑ�sϦ�,)�'�f��-t���r
~D�d �8"'��N����~�//��L����^n���lŸc����\a.B'����L�&����[�HH�X����̭��;5M�5[(Ȏ��̼j���4�PH-|��S�a�~I(�u��C��mb�J��m�0ޣ}�5���V��4��+�R���f�!�}�M�1}>z8-OYpԜ:��������p�o�͛�=�s�'�B�ʓ���G��7m�Ɵ�Xoce�[ 9H:z�G9�_{�����u��-�?�p;4A��_�&�kW��j�MYA��c�o��d�}�^�2�j?w<N!�����)�2ìv�����Õ"b4��~��f���p����*�����R'�
l���� %d�*���Mʕ��g>
.#e�Q|"3�Dȣ������D�UO�+�#�<t�����{^+����W���6���dh�*4x�|(�D|(�f�l~(����G������+���c��lq\V�gk�z|:<WF���G���<'�̞/Ʃ|;=K�ex��l�+�24F
F�ሞG�\������5��dpR ��<VJ+��|R?��e���t�<�z~gK\f�q�c����j�x��G���|> ����xۑË�Z�,*�a��/���91��3gF�ɩ����Q�m
�p�{�>1q#K��A67�^I���Y>&9���B�9>��S�{�U���Ng�v�":�DTTU�a��El�0�2պ=����3/��.�Ǒ����UYw|;�#��������w�wwuUe���'�x�wwUV]��{wwuUV]��'��1��Uvq�E���kZJ�o0�����:7CY10OQ��*4e9���$�T��?�V<���ή�c�E��t��9�;���'!P���!��R�"�!��s7C��2Q�0��S��J9.�N�����N��a�Wj�v�d8R����,Ŕ�d�UQ�iX�V��		��e=8��4��w=UUJ(&!��eM�sՐ�	�u1!��(9%�}�*1_������!���LMwj�룒r��æ���b�ꦨ���*���
>v���X�������-��o��	'qͮ�01���2]91l��Xӱ��<�����c3���&8�UH,8bjڪh�L�II��a 7u^N[)B'*�)�ä�@����q�IZϰ�bB�aÚ�:���@�/3(�t�v���]@�:��=dw�y���L���<H����哽�����l�R��7��w4rC��QZa�Wʬz���s�ֲ�:��by&�ns,��4��4`��ClN'-��e�v�<J�}CT:��(�����L�vl>�y��僮��v&���'0��a�s4T�=JΉ.{L��Pk2u�l�Y�:�*|v�b�Uc�C��N|
;{�i\	��w4�v�z ��KB&
603�����a��Q�!�{ж��x��^Yx��J�m��j芍g1x��C0����f!\�}��D���������nW���ON��I����4YE��ﳝQX���qtn�"�)D�s�	F!�L��]��EScwkb�j\75�J���;��g�~�Jw�jN�R�7��󰡞CQ�\:^㉀f���~E�F�F��u�Ñ797:9~�FDB`D�b&�)>�.UP��P��*T��L8��Z���
`�2��ȁ�*�X"8R�ؔ�Ed���TNF��b��"(�A4�V���*+l-�Eqd�L�MZ�8�nV�%%��ea��.�(��T���ø|!sȉG�
��� ���p�1e�鬪��q�Qf¤�2Lt����S?B�a�9��4k
�b$!-$ˉ�||�Mr2<{G9w��̹���t`A:'�J8"h����K�gÕְ�t�j|����w�iV���A�OM�^R{��XRD����)�g��ȧ���P��((��I��(i�The��0>:��6Ƞ�J>	{��~�����	�EOC���pA2&J4"p��IM��@{]C�n`=��ӓ�D�l2�v9!D�xI �}�6T�}����""��5m�g���q��cu���ˊ����ڐ��(4zdĨ�/l��&���:>V)a�n���f���hM��pD���Ŗ_xg49�S)��gĳ����-9S�A|�K��g�Ǘ6�����.��5E�%��}�:�y���t����~�1��x�%�i�d��M�aс���,��f&a�zL�O&LϬQ<p�>�ʡ؈��N�?
%���U���z���:^/k��v�_\d⸻q�m�W�ұ̶���D��D6	��^
�(D��0]�|9��>(���G����S�l|98U���r(У�W�����lվ(��_��pA��Y&������b'��Q�0���a1�0x0�b&��hޜgK���c�U�x���/���؞8V���\+�����*�Z�8�.mq���x��n���$k�T!^I���s5��f'��zb�������Q'�c6���s;5�����8��X�oe�H�����k���pn���|,��׻���z�j[�ve0�����~�*�t��&f�k�-X��"�4Ң�.[���3W{a�:�0����6!�Ǘ�>œ}4W�3�q�`����_	aܙ���s	E+�"%�*�����[9��0�'Q�֍��h�ҋ�����ڊ�T�-#jp�kٛ��Mmv$\�#�v#���w�����]z�8n:��^���ۛ�ł�cR�&��Q6ښ�Ø�K�H�4,]UX�Eκ�L0M���9��
= �n#*ժR���8;��z�;z%w�ə#B�c��#�N�K�򉊹H��(&
1B������lY�����s%NW*,��R��
��r�J��V;-k��h@c˶�ر�4/�5G$bo(�h��H�q�$�f[���Ϋ�,���7�8��MIcC���d�(�T
qD+�J�r��� L!!""P?)۽ڪ���������UU�|;��=���UYwø�����37]ø��g���fn��q=g���fn��r��)\WX⫏�9nl��\��j�ij�V杷���OA�&Q���B4cm1H�Z�#���d����+T�u@�;b���#f��V�'-��Iѿ�Ha]�c	$V���8q{�kҔe%;d�apܧ��q�Cn�`��5;P�
���nC��~Y�m�)���T���y�Y���ʲ�c���7�O�V�H�ue��ղ����==7CШ`��1H� �b%8g�qMV����s�99�=y���ts�.�HZ#�^`��6a#�����;���v՞�7 ������	�屔���T�쑃
i��r3�W!�?
�<�r`�p�E<���T�CSƹ�S���wՖ����T�+��z���᪈�.��$R` φ�pZ
�)�!�[��LC��e�ڴk��p�)�@����=6�B�YEc�x���۫I��4��l�Z��F�Ρ��iX�j5 �����T�N&S�<H�Hu���p��"zd���^�F)^+��|���]fww�]�P�`��V�8N*��=��3����Dj�.�ws�ŕu*pE�9T�M�8�|�xrqj����2;U��\࢔ĸk��S��RV6d��}f���J4���0i!�d--��ƣ�O"N�t)�+J<Q�(�|vi/F/��}�,hSZ���İW�C��׽x'M�"� �vŇ6ZZ�$��LLJZ/a8@�sr�g�f��8���!�M�۱��eaF��WE��0�p|K��56j,�Vv����C�.Qi�-A:�Z�h��0RRmѰ�NCԉގ�Gl�n�,l��[F�pM�j_1T���D�D�2Q��(�x�b��C�LOVI�Y�<G�4%}�Ԩlܗ5�)`��}P�Jha�1*l��d=��b�GŜW���,�_m=��a!a9qF8�r��P@�ߟ:�Z���b���~;I5�Q\����o�:�)\S�<cۜ��:�&+ �QG�+-CƎ��>�.U��J./�lϊ���v��Qxj�p%�LMʠ�1A���No[�od���Pw1��p�iɺ�՗E���I��c7�	Sp�/1�H��;�����u�ͩ�Ĥɘ�N��0���v.]��J.���bJ�S�x����6�+�=a�iI넣�BC���5&"m���O\0g��J)(��j;�0ziJڞ��1��+}c�Х�9���uTUM��n����I���eT2D�,����
�(��"j8Q��ƭ|u�Ȧ(���अf&b�.s]�hʢ�b�Æ]��K�U��j����g���)6��뭡�+�{3��R����\�����H�$	���g�gpLCE�B�0@;<�i�[E���a
UD����M�a���>ϥ|��؂lCe(����%���L �i�`�l�,4������RW&��f��|cT�)�����h��!p���*�W�*��ZDV1X�	)K�:é�_}j�w"�GѼ��V�y4���vvһ0������8qیq��6��mv����+f͛:l�8�O^��;t��q﫶�m~v�OXٳn�l�m���6��m�t���6�O�v�m�m�m�m�o�|���Zv۶�i�+f͛6zǏ<m��ݾv�m6�m�lٳm�oZm��n��ߛ���y�h�	�[Q�`�l���D\PV?���ɝmw3l�s�(ι��\2�i�^��۪�=R���)�}�K�k��{��޼�ے���ϞH��fb�y�q���{�CF�ȧ;�Ř0T�P�1�±�� �L̱^�	+��c���������������������������������B������$�~�y'l�Ѩ�:э�)3����d���1EӋ�eq��Q!�����H��xc��v�a�d�v��߅Ur�#5}�1�b��J~�$�S�WjWJ�鍱�z���j�0R���Ez��Cs��,U9	�N���V91������ЄuK�1wV7X�$!��v���Y̧ޣ�;�-Z�ry�p{��~z��N���Gܜ�T�!G��Ӥ���LHP��Ј�(�Ex��b���Ϡ���e�*l�#x>`��8�D�Ety����"m�C ��
,c88�ʣ��%���
�P��,RpGƤU�_��9�\�ږ������5K���U8@kW���8�s��Zg�
t�-/�m:�vo�	T�Rv��`�ND�$ɞ�S'�8үyy��b��Lkģ���m#�SIM��g��&a�v��(��=UiJ�U\clc�yg�^Yo���U� *ɓ1���K� �J.\P��!�cU=ML��yW��<;��"�;���`w�!\�s��n�JCT�m��wFJ�4f�J�=6!�l�Pg��gB����\�c�z��B�O�xB�'�"~!���[H���/��2S\�0�#�)�RY���m2�m�)��e���IX���*MKA�I�t����< ��Ok���V����:T*�q�9o�)��!i�C�;1�5URJ�-<B�v¼UV������.��5�L�(�x�1��ùP���\�^��%�]��e���C�o1��Ør\&x����m�0����q�}b��BaM��s�+#���!C�!�<=:�б-KFc!k�n:j�1���U��F��k�����pm���j��\�Ivʼ�������]��3I�X�BBU9U�S�\V�+���w��V؜�i��
8u��f2�󰑐�a���i�/y�Y7�I���"Z[f��or�쪻˴�gR��Q�nO���XݖՍO5;m�̎�
��V�����QF�f�Z�t���75
��{sO3�a<D��9�<{�i���������(�w�v���QxjO���ykҊ���#�b�����6�7�p�ۄ�X�xo2um&$��O��F��ª��+�Ux��ce2IHm6&a�U9�c>ʼ7(��8���dN���y���Kd���(�a����R�I��J2�B�����N�h��w1,�K�U�Rf�bs1\9=��ъ���*��>c�܋��
^X^n�MkpU::�x�����v!~CU��)h&��Q"a���k۟0�?
��8p8��SS�ƃ1Aq'����5=���C'�g�*��!�=�[���u���W�U?>1Æ͸�8�\V�l�q�m���lmU�f͛m^8���4���㧭��o��Ҷ�[0�m�m��m�n�|��=m�ͱ㶝;m�޶��o�|���6��gm�i��b�lٳj��N޶��o�i��b�i�f͛m�m�ӥ��:Eٛ9"�D^��*�@�Rt��y���}���ه��ܛ�7��fzt�zU�=mm?!֯�ܑ����&�%sO7�o��2�ݮ�-
�e�T�ф�H�\#*n+I}�yn;�=�ǳC7X��K4ݖ.���}�-nΫ-�f?�=�x�	%Ռ�y��=Ov8t^����̙�=d��;�uj��K�>u���b4�N���}�atq�&��}���e�Y�Z����:�o�oNf�rJb����,T�-��2ջ�6e���� �Y�,�ͪ�n�H���91�`G쫫T�I"&��u�$KB�M�ܡuQ�V*�Y�� l�MC�rsE���O��u�l}���t���Y���f�U���Y���F>ɝ�Q֛���4�lPm���]Z��ʱ��ЩQ����E���N-W�|�嬢(���Q�
9�Z��V�:���.�/7�w��uJ̬���:Vl-�t�Tm��X�L%N�LD�ETtU�,���X���)�T�ad�(��Ӳ�h�NX�2IaTJ��hܯ�337�τ���������������������������� ���=�=?����=�1Gn�]�H�ݶ��j��*ݰ���	x�q�J�n�K\aem�Tj�+������q��-Dp�rʓM�9lC��/��k��(�V�25�����0�Ý���:��a��Z�	Uox�3H9L&Su2U
!*��2p
L�����Rq鵃By���(�x���
�`�T$���e,l��c比�������dj*�c|������c9T�26�S�	�	F9
�1�rCF�q���'6�&��[l�r.�Ξ�B��������9��O+�UU�˧�p�^F�m�ݴwߏ��Ԧ�<��(�'D!�2QENE���u��p�|b��x����C�I0cf���4��T����چ	R��V	Rή(bոcf��R�ap�d�n�!ZU��}���70��N�9������±Xc�Ut���<��I�4�xJN������_�v������KV���ȧ�=���i*�QU�6�ݦ�x�USB�,��ۆ!�Es����\�%Cp����.q_�C>Ȋ����
�Xc�����|��Α?I�|>R����feQ�<rE]�ʫV��4T��~׸��%��,mZ:[Q�*���sl�p�y���G��NU��\V��`�
�!P��fɽ�z��x���^+ʻ�Q�>⼽�;�[Â[iz֤$d��f҂ҏZXR�9�W���LB��� ���U�RX��!�{�:�vQZ���{V��<;a�:UWl~QE!��*�ʷf������i4��ƍk�&�&6�Op�|J<�Ձðz������d���DU�QHJ���9j�Ʉ�c	��e6Кyg]#m*�%O�}����0�J����8�r���̨G��2��d%RR^�:�H�mP�<���9�%�a������Ә��5X�A��,�Ɗ���f+�>c*��U�|]���x���i���j�Q�-W#��Ì0ƕU���|{��}��u+�߮bt32mG�K��%PҒ���K��bb$^�jh�>$�*�n�!��'�Nڪt���UEpeQ�7�},j;�jj9
=>a�>UV��cm{]��_�ǄX(�N6Q�5e�:k�k������mU�*���i�����*K%�&۶'b�R8'UnD�Sd���J*)+#��Uz.�9#�2u9�[��#5.1kuT����f=Ý��3Wqz��Nˍ&0o5L����M�L%��qQ=U�����ۆa�s@r�8�:����+��'xX�`8��-i��}�A��S�vNCS��c�Uv���??/
˶�M�S�7�<�1QN����`��\��Ҳz��Cx�ʵL�<o���sy�����3
��)eBX˓0_�?c����ŎG��̤����Q.T�o`e<�'S�)�G�'����8lٶշ���u��޶�o�m��l�8�OOO�+��u���^4��6��m+g͔�m�m��m�n�m�g����<vӦ�m�o[m�|���6���m�i���Jٳfͫ�m;m����;i��b�	�0�..M�0p�D��j���łk!5#d[��AYB�m��B����6��	wn�U2�bA�EY����Bd�+�u^�s8k&\��}@9�$�;���W�'���t�XP7)h�B�CAP��І�m�d�̼�xt���陙��xt���陙��xt��ꙙ��xt��ꙙ��xt��ꙙ�Ըt��p@ ���c�9s�g#M�U�����O=YE��>��A��8\_������_N�1���h�M�{�����SS�8���F�6�u-�ɒy\��9�ꪚJ*�Fv�O�v�;a�<UV��c���[�U�	���E����>��OLCp�ȫ�I:���a"��I3N�=9�+�S��}�<v��,K1�ԔT�"m�	U��a�:x�q4fHCi4@�90r{�RE ���^i��z�r���{:m�j<�8�z�CD���}��b3W$+tgO1���5lw3�Ko���+2,�Wۀ��i�k�jM��U�ъ($����+j��RUNrK%X��*�7�b��W-���[n�e����FsDtI���2�N;i)�r�1���C��0�,�S!UEJ#��"p�i�xD�F�Ӥ0�p��%���hÃO����I'�}REbj�R^8t�����{_ط<r�������bpDO�䞶���3�"G�|�N�^'^5!��)�g!�>2R����#	����M�v����zc���˕�f�aU�!�z�#�7�\��Yx�Z��[�ԯǘ}p�(L�d�P;�q���?:�9�f.<�O'm��1��U[c���o��,����Y����nxu6���u�I��&�hs��I���~�'�"��(�+--���$��"�BZvu�l2�>B�S �46`�*`���ge5H��oԣ�~OsF�cp�>��~�Qd��Ҫ���+u�L��0��!{� M�<W�Yј��Z����llT5B�����+��O�B���Tf�v*q��A����bz'��B�5�,31tQQ���IG30��	s����:�<�#�6����d2܊�Ɖ�����s��0�Ax󓘠�&(a.,�ŋ+M��L��
Z��Ҋ��s����+@UE/�*5(��.b�fEbh`�РI�7R�ŗ��L��Zn�!1�V4m+̦�iԍ�ʒ/R��H�J4촴�k�T�2����[F\���	Ϻ���r8ڱ)m��8��"�� �Ӡ�{�ɚ�I��"'B��L�D��Ȋ��n3����δ�T��s�#�)��d��CW� j)�g���y��<�>�I��;��Ǫ^��u�l�l��МS�Qż^} j��8H�MѼ��O��RC���U�1�y��ԶI�&���J�#��eJ(ʦ�L�)��%I�T�9ǽ/_UD��F�H��m>�IyMq,��\���u����gL0Ǌ��(����2�H�1U�s&��M%���C���� �����?��8�� <�[
M��6�����Ւ\eQi��N�x�52�n�1��A���ϚH0��'�$�I$����(��������8`�x~����$!�
����D$2L���7�\L��IB�QGX>��
E$���*B�RE"�)"�%"Ȕ$U��T��J��*K��B��QPQdT����Ȋ((�"�"(�"�"(�"���(ְ�(��,���J)"���(�J,�(�H�ʑ�
*B�H���ȔT�,ae���1����dQh�E���Z,Qe��Qh�E��Qb����B�,��Qh�E�ưj����,��,Qe(��[��]K0�#�YE�X��,QGX:��ұ���ꑨ��b�E�,�R�Ya�#�(X��b�E�,Qd���TQeQe(�X���#%(��(�E�X��,Qe$��(�RʖQb�YE�,��Qe(��YE�YE�(��(��YE�,��QR���Qb�(�E�X��,QE$���X��,Qb�YEYI,QeQe(��X���,.b#"�(�E�YE�X��X��IeQb�(�E�YE�X��I�F(��(�E�X��*Qb�R�YE�YE�,��Qb�TQR�YE�,��Qb�)%J,��QeT�,RZ�b�J�T�R���K*Y*R�X��,QeQd��(�EJIb��X��,Qe(��)YE�X����(��,Q�&RKX��(�E�X��(��YE�,��,Qb�*YR���c$$����X�b��,R�*)e,R�,Q,�JX���R���e,��ZYK��KKD��(�,R�iie�e,�ZZYJ)%��E)h�J��X�U,R�))b�JX���)Tb��dR�,���JX��Y)b�J%R�,R��)b�KY(�(�R�Y)b�JX��Y(�)T����(�K%,R�I,��K%,R�,�Y)b�d��TR�E�Y)h�K�T��U,R��d�X��)(�K%,R�KK%,R�b�)EJQKK%,R���JX��Y(��*�)b�J,��K%*R��K�Qd��X�R�Y(�)b�JX�*�X�d�"�2"#`���"#�H���D`�1$`��R�UX�%H�VJ�V(Ȍ�Đ`���#"0FDDH#�dF�UR�UU��R,�b��RE����)��I�!*"T�	ңP�� �(��RE"��TE"��Y	H�JE�R,�C�J"��TEEF@VEVH��)��d�%��~�9�����Ƅ�4R�����I,�"ղڶGw�%|S5�ֿ�k��k�����4��9O��}F>���o�~��?��|g�������C0~$�a�w唡$�����_)���^C�7��ωg6}�����
|�S��������'����9��������~�A@?� x��UQ?�����������?���>ϰC��4�JT��PO���'���?����?ȇ� ~C����O���~�?��BHJ�����������V��SC���������F����:7�'֟��5,��)�fF��������� ��mE1TG���H�5Dj
���*( �{0�!Zf��%]7����ð�|<O���p?�� �J*�����T���Q�AADe�O����|ؾ	�8��_���g�9 ���d�`@�n�/�B?��>�柣�HEU��h�-~/�_ͯ����9�_��n���a���!�J�������h~'�	���2?p�?�|BK���_��O�~�?,�&��}C���}����Wڲ�ҿW�~C�6t���e���0O���UQ>o�+�?����U�]�P�>i��КH	FP���*(\�}B�l�[�tY�jrȐ$`RSG�<%4C"�
�a062��rSB|�	�89w�?#p0Z�ݮR����?�x  )J��RHO����_Ժ����}�����O�O��>7BP��?����>I�T�H�'���n��?r}�I����_~p~Ĉ�����������'��UTO�H�y������~�TM������w������������>��� ��i]$����~��� G$�0Yb���n���i�?'�~ ��>=Ȗ}�M|�-�ϘdEUI�	��~�4�I�O������z'����~����蟟�H�@����dR��Bx�S���?��'� AA@)�~p!��	��v�I�}8((�Ba*�'����Se'����O��
�d?�*�- 1ςo�����w$S�	�]�