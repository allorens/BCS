BZh91AY&SYx��ܨ߀`q���"� ����b%?     `                                     (  �{k���  
  

� E   
U P�(P  �P   �   @  @  ���T��D�H��*���$��R��UI �P��H$JJ������UEJ@����h  �H$��ER!
����W�;�;�"��%�
�`:��v-i�J�Ѧ��I8t�9 d�� � � : r}󇗦f�X{�:T�B�M�IY��ʥ��ĥ��k�w�(O��U��Ӑ g���A������ �| 
  �|�m�@YQE$JB��DD�_wr�T� }3��� �X/@{� ��y ǽ��R�� 6a�� q ��<��+�ǐ =w��J� >�����   �   7A� k���� ���Qx:݇�� r�� 9� ��(� M�� 2; �� � ( ǀ ����"�UR���J*�P� -�� n��� r ��I, �q w`:vt�� q�R8 ��@�J� *���tPH`� y��[�(0k� 7`Cvt.�
+ ��݀�S� :��  |��	>�RB�D��HU*�)K��>�9 d8���*�`6: ;���{��Wc��%B���}p(  ��  0y y��;����� �����3� �:D��fu@�@�A��@(=����UB�$UP���PH!_ 	 � d ��`�:*C������ �;�)Gt�@��4  P7� ���0Ǹ�	< d<@w0Cv w	8 �� ��Gv >       � �� R�0��dbd��"��LR��@    �Ѫ�aIH��1 0	�i�L�l�$i��2 ��  Ѡ	4��Ԫ��L� ԩoR�0$�h&I�M12z&�}��G��v}ݵ}��/��Z�7����j����޾<v��D<T���wB*�
!�Z�WڪD;]E������_���g�^���Q_���m��uR!�5z��-+�^l��>?����?_�����N�H��H��OͤO���ROͪS�h�ƅ8Ў1fE8��iEq�Uq�'Tq���UUq�8�K����q�q�q�q��U\dq�ƪ��\hq��!ƕq�\j����J�Ү1W+�K�GU�q�\e.0q��dq��S媸��C�#��48���j8Ҿ8�q��#�I�'�e8�q��IƾN2�e8�we8�q���18��0���#�S�T�Iq��N2xb��q�q��28�yj8�q��'ݔ��G�i8�W5atӌ�48ʮ5Uƒ�*��q��,�q��*�C�G�i8��T�)��:j8�q��)�S�S�.5j�e8�8�g)�.0���4�h��q��Y���8�̎5N4\aq�q��E�i�.0�ԸԸԸ�8�q��GN1\faq�Ɠ�N5N4��G�N2�5W0q�\j��4W����Rq�\j����yjW,��
�%q�\eW��*�|5ƒ�%q�wi.4����*��ݑ�Uq���W��+�U|0�J�UƩq�\j��U�4ye\`�
�
�T�5S��5`q���zdWf*8�Uvh�q�4�ƒ8�Uq�j�ƩUƅ_-q�x{��@��}��|C�6b0��m�Њ�F-�JM�F4e�'��;�ڂ..ƺ)��q	;p�����tCBa�8��#����y7��n��y�l��td�g�.�{$+u��-p�{��"ݻ`D�'X��Ĭ5<��
	#q�y�T�}� ���tV���,D��*�w�:Uߩ�٣�J�[Z�v��S�"����b� \��0��Y�8�WKڋ���;2�9��9��v�wn���5�ގ�D��ڀ}דT�!�Nn\֜��~[�ܻ� M��`��8�)�nrR���c	����jQrl=���֙8��\{��loP�dpy77��*�c�1z#�7`܋k�{��E���
�#\8Y�)i��J� ���v5I�r.�S��7��2M�u��mݑ$��Q�����z�Wv��t<;��)�_�;��U��t�j]�9���`#P�n6��ǜ T�x$ψ0�Odr�Kn�OX�E�k'j��C�zf�9:#w]��q̫b�]9�>y�_L���u^�V��1Kǥ�B%͝*m��R��>(I6���f�c���Aĝޖ��a�3�㛁w܁�����l�ZS�e�u<o;�瑞X&^{�;�w�K)�}�*�l#��J�S����(@��k[�2��Rsa�¶������g^�3.�P�6:;e1{�u�.�N��x#�b�6���U�WHZW�s����an�@�	O����f�&j�>C��;�P1�Y�bwH#08�]��"kq�g�X14MVy
�b*wH�S���g��G�}z;��2�X@���ep��F>]O'd���<t�p�V䇻7w�ko%7$m��rH-o! c�T��;�.�Q�����W�"�b]Z�J��[�[�.d�ƞ�]�4�;x]p��gC`N�m�藞,6����Ѫ�/\�c��{�H�;oK{4ئ.J*���H��v����ݘ�.�od���.�4$;8���fC���V�k5v��8��ڕW��p�yÚ�Z�߬�У�<���z�{�:v���{n���[����WE u�z�9ۢL�1�y쳓�/D!����6����Ҍ*�q*��uǃ7�Y�%��e�t���m���R	Ǜ����mO�^�KkJ߸e��mF�)+��N�oS�A�mY�7H'KɎ��N��z`��ۏ�Ly��;�Ӕ��n��1U��D�_#���Փ[/M�otÂ"�K�'��UɜV�O��D7ue�g{C6S����nlX�z88�c0h̨N�]�)wq��9]�ۦ�%�ݕ���9�ˮ�whH��V��A�=�ݙ^p�u3���7.��3CHf�Ml����#4�6}t�9�-�|�9oڪ����PY+:	��2�]�t�&��;��j�K�ov�۰L�Gn���eLj��kn'9��%[۽�%�n�oR)��Fi�=3{tf���޸V0�ҵ�5��0e�J.uq�λ˺��9�`��2�i{�&�k±;�,�;w��m�l��>�q�f�`C�c8��Э�9;�����t�.^�J�u�g8�;��S3���F��0��-1�Fn�[��_X�`���Ρ*���W+�ˤ�q� k��!�l��Z��0l�����)ӔCτ\^9�7W[J�Fv�6	zj���{���Xm{a�*8�`����wõ+�7S/w�|�6bZb����tTN:;�J��I[������7u�(uvs.� �������oz.At�8<Mf��L\9q�VN׏�p	�(�YU;��n�f;�{4�\5(�9�F����7�%��V�F��8Us�����ݎ���	��ڟ-ފ���/q�9
ǝ�Kp,��P�)Wwt�QvLլbUN�l|�$�l�.=O�����F	nP�rvRR�d��=7�g��+N���F�:F�!�%��������0��d�ٙ���,��po��rf�PA׻��E3Jӑ�o\�wV��'�ѣ�uB;t}!��7���[{s!E�4h�ï7q�l��RѽZx��>MEB�ָ ��h�F�ޫd��h�j�tgx<��4����<��xq�<˚0�dƩX*�ױ^�i�&���k�V��7�۷���=��^��^��u㌝����np� 2	��eD�����Tn�{��;N�X
����^��W=��X�4ȷ�;ww�PX`�h����0���C�s]�Wz�����gm[�"���sw�ӝ1p2u]p�Idt���Zp6f�o)�S;!��7j�󝦄;z�I(3t�#z9�E]+[��@C%�8];��d�*�� lI+��c;�E�,h]�ڙrĂ��p�.�N�WWc���
��E{^iir��L����zQ9��Fh�f��^1�<Y�םfo��'M
$Pݸu�uk�v���p1����㜅2&͡���.{jї%��°��=���������e7fq�Ե�EZ��6F0�Mّ9�@��������3C%���ձ�n��I�ػ���2��m�;yn�sx���ѬP�T���ġ���Rɼ#��cBD�!�#@ѣkߖ��N�i)S�\���%h�[���O���a�'v�����7.��8�b�^wR�0�7�JZ�MI��{\t���n�n԰�M�x&���5���k��A�h�m�*y�d����p��e����1�x4���]�`���,�i��)�1��ccr��eб'��˳C��d��rH���t�no����J�XX3O<��v��8���vg]Q���G�;��y��[ys�I��6d��*vyr��	����ed��7R��U�܅d����U�=ok1+�@,�=�WMȂe��ܧ�+��V�rEn�r���(9�U#_gaFbṳ
��}� um�y����9���$
u!�j�ywk�7On�2�{Þ�ٻ���k�{�Wv���j����1X�tXV�#Q��4�i���㛛���3EBn�wd�^����wCd�ےE;wht�Z����7����΁�.��O\F��Y���3�>yF M=���\sx�N��{��z����r��i��8���\��:.��jZq���nr�&Ñ���{'�2g^I�˸����
��`!ݥm��;gp�*��Ό1�Э-ֺ�8wQE������BP�c����<�n��liMҺZ���4�:��̀.�1�vk�p��[�wu^�f���9�Vn�7.�c�����+{���Th7�u�;4��aW��j.�F�AՊ���k��{&�[�8�ɛU��RnQ�20u��ۦ+ٹNnT�L
���7@�h�p�gQUkX�2xv�m .�n��9q�]����P�@7BZ��/���!�Qѥ�H�;QZ)+q�u*2ې�2�-��sA�t�9��L��h�(w���`H���<rM1t�n���v��)�mC;K��!��J$acW��0��e3q>�0Ϣs4��Ÿod��Z�ⷆXro��s::�ږ����j�}���	�����෱�Z��s�h�(;�oK}����P�a*SN9�R���=�u�0�,��76S,��<�g^9;v�f�ˢ�FnTm?��mc\���g<h�B@ -͛�#�w����1b��K�f�.o!�,mYf�Aq�۽	�N�ێ��Lp�XbpKWe{����7���xVF6�!KH7;H㯎�ͩ��I�{F�t(��1sN��E������6ϙ����1�{�ᒲ���,�xnv�/��uE�u��[�m���ii�W�����i������@�|�C9��{�wD���׹t��Y��RĚz!��0��ނj�9� ,�	ͭ��]{����S�Fu���ڱoh���8,BL���[�p�CV��@D���W�eӢ�gsc=�q
�Ĭ���Q��r�͞ޜku���`�ۈ��������5�.W^�X���9�./m=��g:6c�[�s���5r<��k�t.`�.y18k�xZ�^�[õ�7:�R7,�g����nc�_uF�j��:�L���JO,�p�Gz��3��ݰ�P	5�-�G�V�q�loj��NrgU�w@䕐.�0��Gvg�Z��K9Ѱ��2D:��E;,5�F�Ҕ�yev�q:S3�f�k"m/p��Tq���:W����7H����y�X+h-)8qcG��9�,�����H?U�F� ǌ-�-�O}��������i���oG�d�C��oF՜�vL7�߹՝S-�����d�L�MT7���Q��F�]�6�ҜZx��i�c͓@]��pF�Bhy�Rw.wI;�׌��s\����G6zx*79�7��};BE���Ǩ��	�8F�
"�$�b��r��� �l��	KnX�c:����on�
����h�:��ܝ��kz�j����ȁ�-�UNv����;����vs�KH8��+����Gf��Y�]խN�s�X�<Yl�{)37DM�+�)�,
o�v�xe�Wq���C�MN01�K从�o˧{&M�mc+�Q.�0v�SY� A�˴��֓�	iGꦯ�n�q7WO��*t�2{���y�ӻ��7�v��:�!��v�)�ط�����4d��Y�PԯMƷMy�[��c�_`����z>tr����R��%��9�Tu�-aD��������'v��>�`ד�u=|�Ks��7�L���I��F��sB�.cJ)>��"7����5h��'G�jǋ�Sl��5��n�V��h��wun�bz�i�/u�#A]8�`�RZ�ֹ�o=��G��{� X[��zu=�w77��.���]r^�DU���A����h���@�V��M�0�X칢G�n�D�璗���RS��}���oC�-��u���l�@����f�����RjxLŰt����%c�na;S��څ�lL����R&)��b�V�XP"��V�J�5���z �F���ܗ,���ޘf:��͎�K�����]��8�����8c�n��2���ˋ_�΀������R�T�7�Tư�O�&�ڊ,�6��ve�Z��u��d�M�*��ُx���˺A�����8�f��]���nYL:{:�E³�7�6��u��>d@�#I/�^�?k��3�a�`�Æ��-�N�A�,jk��Yr�(M�-��&zf���a� �p'�\{��=H����5�3�\��Y�2�[W=D�C�r�W�s�t����$��&w�#x��\�z����/�&�`�Q�R�R��Nv������i��p��S�"cy!\�fp������#�a�ˑY6��ڑ�P�ٺ�������풤�	[+�oL����b8kO�GFL���)X�te<B�g���Ѱ�1�'wy�j�"ɻǎ��[��p�׵��C���r����nIf�ɖ�A��v�ѳɏQ̪����)���{�(mI��`I헵�����q���u��w5	4�#"�K������އ75��9�짣ِ��$c�t$�ی�����9t�k칶L���i�_ۈm�<�n�û�$$��}�SϺj%vr��4����o{ͥXE�؄�Xާ��5kvھRkḨXՈW;8ax�x9�Q�����ɫl�n�̶Aݧ��b��A��遀����>�ۏ�v7)$d�:.u2�g&X��ԔxG$�o�`�u�b��չ�oq��;���s�R��E4s�F=���]ѓ���+�X<[���s	\�U�i[жgn.[���!��� s;D�ܫ�{7ssfR� mu��C���ÓW��n-϶�m˼�K:�S#��K!O{ʉ}^�����Ml
�Ӭ��:���}�r��!�`�»5t�d��)��l]�^ǜCZ�4�4A���λ�qQ@H('@�(���q�tS��(rq�@��:˄�:'��!�v2�ˏ�Ԕ�ÑS�-�̍��a{�2�������Ֆ�qq��
V����;L�5��q�Y��͵s�r�l�R�����J

��Q��i��+��|�E݁K{���,�ާ4��n�8�����%_g���_�ƾ���8s�t)hxNn�g17t�q�gL�ѳ\����¾\��f71E�{�p���Qn�P��&s����2�"���q>�g|��E=��]�9�*��B��{DO�mL�������3�7��K4�5���I6��m�����3����Ux�˻7��K`ĩ:���MQm�աdq��O=�sR��r���O��(��cGdǍ��9���~,g`��B���,z��$���sp���V�;��O��l֋���f���<�S5����ݺgw��ڒ���ŲPx$�N��&v=ޛ��ǻ�TV�5�{LTL�s�r�V�i�.�s�O�z�4��8�F��ĵg�j��ג���{_sЪ�ĵ~Nj��=�4�5ws��ڶ��G{_�*��|�إjɦ[h�;͡$,si���cԎ�3��qx�$Aw�׻ 1�v������^Pk1$����SCHՁ�ґ�W�#s�����^��dp���?C�|�}{��F_g,y�:�N�#s��;6^�l�^�<�|{���yۉn@=����?j����Uwo{Rg{X�wN�tN��iٻ�`!D�CYr��R����Tu*���~�����������}~u��㺒�ـ�%lBثb�Y:җZK�����+�UF�+���Kd[[AT�YU։��u�.�Q�Tl��:ʛ#aUlڢ�hWYki�T�d-�-�i*��"��[$u��jl�����U���U�l��R�%���]d�ZShT��]e)֒�iWZ)�S�Y*���֤��[U��#iKbU�ڪ��["l�VŴN�*���u�:�F�UmT��D�6�V͒lSb�"�e�U���u��S�+j�Z���Ҫm�QWX�m������ݰ�A�9p��#a��D')Ho�?���d<�}6z�_!��"�-43`�Oy�-W�|�q�:�f&���{�u�#�3�L2���K����ן͒� ��7��!�AH�[�x�z���9V�Kb�lC��<���3���W�K��n^�V:�/6C��^����O~z�FOBB/�Rd!X]����0�
QE�K:8Nm�OB00n� >׻�HE�=��:��-�����5�(�I�����}��H��������^i�{�*G��xz������� ���o�+���o�~�'���n�Ҕ��юn練��v�g����9X�ص�=��۽L㦻�Gh�7}���ڼ�^�%�~�]�dz����\ќpi�Nvh?k׼ǽ�Fz��&t���ί��e�]���[��*�>KۍǱ��N�"Oj��Gc�y`v�Oh�p����z�^�wF������Sg}D�>[ï���-x���E���]˸���H��)�O�ugsHt#�+ڽ3؇��j�7���}27}#�4�t�yQ�������y���qh|v͘-F{�9֒V"�vu,���:�v!|#����v�3ڧ�X��������W�#<�[�m��BMɆ������ޣ�Y@����uO{!���z#�z���iS���8��N���s��hv�ɕ��O�է$eBV�~�$���ߙ�����q�ֲ��y+z��b�}��=�e��T1x5��i�������9I��Y�>jd�]�1��^��u��T���xJ=w�}�����2�R����������a�HS]�:{�-k=���yj�B�O���y��gs������5,{�>Ľe=����6�ƨ8&��q6��Ny����ۏ�+��pː1ǃa<:=�jf�U�]��dr�^�{���С���8���z�x�'��{�X��pc,z]�KL���2r�_��w�6R�Y��A��*8���/g�gD'P��Cx#3�z���wl�|fi����?��o{�zy6};ˆ�[י�	��,�.����Xzo�/|׉_ogl�&p6��ü�7��8�.ֈ���
�z���$�Ӄ��#��Y�!������x'�==��u xym�7��o�<H�7�N}@mzo�/Q��N`�{om���1��y7M<^��s���ш{��q爗���{��AvP{����N�7�y������˜J_��y�KX�ٶZ�9�{}�D�����0gi�~>�]�r���$yxݷL�ţm�~<���$��^�(vh�f�Qtp&�H��>�/��+�w��o�0}M/7��j�5w���������j��7�7�>�C�A�5gpei]�>kc[�x��;�p�?@XXI���w��Ѐ����[�������˒#<����Trr�+���Y+���n�Ux#����J�M5���{��[�81v���YDbJi����65O�ɢ|��F9O��&�����T�3����z����I��k�H�%��y�hц��CG��G���^q���'�Ð��Z�vkt٧���.���Us��|<�o��p%v�%��5-^Ǵū=�g�'��_ ���,eN�}�$c}����P��5���]
��;���U`ǝ���U�5�ׂO-=�������i���b J�h+�+e%�>jĸ��[ًv`�2n���/T����+��P,�a��J�e����j�܅{sm�7B0�W�?K�3�-�0���o���x�ӆw����ޜ�~=_3�z�k�B�SU3�f/o��ݻ	'���4/q��]C�s�`uߏ��
��z��5,�#�ڏ�230�c����ϒ2��oq�|jQ��o£	&{yE�B���y�
���ʲe�v�R��&Zo�܏���sFm��8�ѫ|1zuw~8�t2�Q�c����4�kÛ���"��*��>0�p�Ji�c2�HE���Jf�h�{��(Wc|WnM1���yvЂ�/,3��\e!���G7�#^D��/3��<��垺<��i뵉�&����߆k�n����<�p�i\�wb�7�?�x.tr��f����`�޹o�/���u�� /�����7�;Gwo����{����Ȱ�	4	4����O=�{�h�r�^������Gpye��)�놀���gR�p_Dc8�7ۧ�s�L�t�/� ^՞6D��]�ӻ)��{[�t�����8��������]e{��rudyY���l)��I�����N��~]�>�~��58*ogrz���<`��XjT����m>�z���JÅOG���
�^�ڍ/�ߍv@�;�K��7 ��;�!�V�G���^(V]�I{�.�O+��ݺ����hC~���y1��5̤y�~���J
��]�/|mz�}�S�{:�}���M�s=��-��#���^�r�i�O������;���W�a^ �0�L���Mž¯�/ ó����us���/N�j�|��S^�z����{��-��?�\����Z)�N Zqx�����zg����r(�ǧ��G��tY���v��U�Ν�<z�y��'�����bS�%�!�Y4΍/VC͇�v`�i�T�x���T�:o�=��j����`��:dؽ��ٮx��$E(��N�P�5��%��gw�����{�{Bа
`�e��9u�q�5T����O�����3�Q��?��y\�W�iq8���l����e�a���ۏ]�	�{�������'K�4{����{�#��hs�TDcˌ5�GZ��'����}/��'���7F�^wcƽ
ރG}��w�N�F�����{����9d�,�N����wO�9¸�};�yy�?nT���Ӹwoil�u�NT�a��=���� :�S�?_%�ᢠC�;ó��>��UO����[<�܀lǈQi�Z��̽UWU��x9Ύoo�uU�����>�b����ݽ����a��>=�T�k̛�.;����}1���Ƈ3���G�Z� bN.�ff]�R�(�3�93A�4fd�W�N�g�������\t�<��#1���C*2'j�ݼ>}�N��m^���>�s*×wV����j�#�""����M��Kh�u,j�*��3�MC(QC����rgs�Հ��u�uX�N�)��hY�����ޝ��e��ژv]�O�D�Id\`��-L���0r'22,��������R��0lV���!-6o8�VU�|A��%�qP�.Y}USb���9�Eͧ=Y� ��F� ��V��Z5�9��iw/��_c�;6��"),|���3/%��R�ن�KO,V�g]��Y�	�����{������[ݶv�X�Ws���3�������EρW��Z����'�zxo�j�ty�J ���B�y3�7Ù�H�R�����\Kt�H��"l��3�ot6���8�J�(�˾��"wz�?G�������<�ye��sg�|�]� ��/c�_>;��`�nib>����,��dx�}z�M�����h{�o���ǋ] v{�T
A��y�J��y��w��[��M�s�!�~��X��K�}�{�K1�I��lNn<���4Io]v.wQybk(�w�)�׻�=�6�<���tjƤ��c7���Ӭ�H��:nAppP?^��w@��.jMz�{^i���N�������i���0Nzx<��&���wO���:�>hz^��.�^[�ۻ�Eպ䎗�Yް��W�퇟{�{&��#:3,Y������e��n*ΫZ9�Yͬp��i�L�:iZ��[ns[�u�0��÷���R��Z�P�A�U�9��z�ya����>�%�`��W�q�Q���@!�=���|�^
^Y;��wV5�Fc�@qW�S���Jf-E#Q��S:^�r0�x\L|7��C��C��w��#��AW�q\N�|�[���g\f�eS�v���B-||Ϙ{�.�E�r8��}D�;�j��f���|��F0(���s�TB�B ��u�ðY>���x����0?�x�7�粯/b�1�UG�)^�ʯU0�=��k�{�]o�d�td���ſxs�u��^G�#�Z��,�\�	`� ��wtlbvo}}'K��4�����Y�� ����nP0A�!{��1B$PQ����\q��<���gz`���I�V�v���/<�^�H����T;���Ya~[�ysZ�È��_x���0ܜQc٧��3y�s�u�����n�B=j�����_Q�f?8.^SϬ	!�3Ӻ�b�o̿5���m~�]�Ғ>��c��;5�|/��%Y�!]��!{����;:{�~���\���}�ڪ��X;���[����iZ�*�����������{���f_��γX;Pܢ﫛�[�Ex\Ѥɞͨo����}˽ux]���f�t�cg��o�{a�ު�YW����h]�o��~~|7����exT���־d{���;H��:m���Õz�T��o��MYu{�k^���O�.����&v=�y�ߪ$�����etDLS5K�r�����K���3�xg�\7��{��F�ݛ=�i����O�u���]��s�^Ku7O�bN~ȴ������4dOCȚ@��a����\�����^��t4x�
3�.+ӏH)ڽǑw,������<~���I��	޸���|��|��Z��FN�|�tq�ܼ�wF�q�~������ZV��y\��4�.��{$�&Pm��D�>��7�m}���|�4^}�gvKgi�/��N=vܳRL-���z���m#(��y��zT�W2!�]�,�f�31"�{E�>ޠ߽[�\�3���F�ݞ���������\����}�H�=C�9e��e����XУlm͙��� {fx��h���#��{��F����Mv{�����i�=ŏ_gd�V�����Owv ���������:�=A�񘳖-�q�O5�����u��{8�yl�{�|�6�-�2��Z�?-
ѣ]@U�0��.½���{&�����⣱Z:�%d��N�ъ�>}�Z.���Y%:ʘ�ږ�M��^����OG��=���Z��Z1��ތ��v]�}�f�g����Rzz!0��X��๢8�G���L��zg[W����z`L���݋�}�SÅ�<OZ���rG�a	����p�n{|_I,ܕg���=���^��7�.*�q1J��ޛ)0;W�ձ�ُ}�' �m��B��z�~�k]�����o��������Ig��#��^"n��0�d��{_�o��3�䴔���
l��(;<�%�L��P��������l�@纞��f��zy	�#��qJ��M��ͪࡿ��9�t��d]�o�E픰��Q|xo�힦�^��G�Ǯ�\w�6��ګq����&��]��3�!���K\�{��~�@���u>��7�S��.�8��N������}��ɳ�6�x�}�y�z�=���<��s��ZX��>���^�7�*��m�u�|sH^�߅�@�5�G��x'q��2!��w�;X����{��^#G�}[/f��51]��W�$�%�ݱ�ǆ���r&�S����Cd=Q^Y�ws����դd��%Nמ�{ʙ�
P��%��'��gU(�-a*��6B���eD(	*b�&(�8�B,�FQ˅1�+/�g�:2�:����䓒`W�5{�y-���O�ajŸ;� >�Y�n�y{t��of���nQ��s\���_|�B�`LÌ���^�$g���g��~��x�Q��-���|�{!�v;�(� ��P4thʏC|�۞��Ӎ��4dKe���D��4��z꧖{�9��8���}���x��7	 N���{|��k�K�-�kn�|0k�F�{�=���WM��d�u��s1)6d��]#�흯7�}�#��̾�Yʥ�*�cZZ/&or��9�GG\�pj�Fr�}���~o�D}�u�o����n���֞���`��z��=�3������'�d�Ͱ�O�N��'s�FA����ܒ�#:餇��W�#=�`h1ڷ��XC��*�b�)�M���_Y�ިSN�=龀,˱S�������Vz_pK�{.h�#۞�(8k����N��G��S����l�����{������6�(۲`�ynN�q6��;��v$.�Z�������t,��s��~:���&�����=���4�e[/�Gǭ���7���%�#p��Y��7�E�+&y��s� t�z��[��$}�d�+�`3�o�=���U�.߼�ԐDS�����'4/{�jٛ�S�a�ǉHwQ�{�9 �ݫ^�"�c��mf[��(���fF���{���Sw�==����ƲF��]�g}U2`�úp��'�ًn?=���_L���LS���S$^���_���xm�zOJ/�{�4�k���7���ľ-bs��'cM��~��+�O{!�n��{�ðG��['b�9�y�:�I�R�\s��<X���e�����i��)�1��Ь���
�� F7�Gfx�	,�<C��V'��t�I�jO�y�}z{��.v��o��{���|G[�{�7`�rN���.mmxｃ{��W�=��9�3�q��L�<�#�r��i�N�{����;}�{�<�{��/�)��~;���Ѣz�_�=����OqL�W(�c��{�/n�K�5��JJ��v�����'gbg��8�7K�g�o�Av�y{��}�&�;{,��+���n�6yW�f�k<�ne:�St	�ݘwf	���E�Y�\�M��/{�3��ߎ�c7�WFHğ�N��L]��{}���S��^kK��ѳd�u�Q���	�fyrŲ9�;ůwxn��(�rs���<Fo?a�6w��ߝ�A�a��o�_�^�|�"�wi�8�|�����V��)5+kK�:\�r{�[��s�����}��t[鏂��6����x�k�)<m�Oiѱ}�pq�Ov��~��!D>ݫ�~���~���y��?���c�x~3�~���������zzzzzzxxW���}��2s-nf.\���:�J�iT���3⥹�̵eG2�dq���ɛ*F5v���jJ���P%��9�v�,�K�ZVpۙ�L�]m��]��U��9�mV�LE�l�U�1Е&#a�7]z,��,�%�M�l�Ain���v�M��-�̱�!f�#`P6��f�MJ�åY+
����]��s�k���[q��0Y �Y���&ͩ����@`�P�������bR�7lF���cE�u9��#	h��5��S8+��-��N9�Y�jEGet!v�5*�ra��:��[����H�1������إ �W/.Wh-�5�3$e-0fq��e0����6l���X�(l�c�L*Y�5j�)"���2��nؙq��l,krҙ ^�l8\�-�IeU��u�i`��c���dU84ֱ��Y��5��Rb��.*]\i���r(l��8ЦU�Ma���B$��48�m�h���KA@E��:�r٢ L��rXq�J�%�!3n��F`�¶�T�X�3�eu�ō��y���Aj�;f�6t���%��n�3�e
��5�&\�h4PЁ���m0bYM�s��Qd�`��X1�F4*ڔ���s���E�m�ԖP�� �f�!�F�R�v���D�z�ܓF6-���=q�Wf��Ԍ�+fL�2\ћYk��bk:��)n(֫r.Q�V���	r���r͒�2�Ћ��fۄ&�
�L���6)���Y���2&���XJ��d�Y��t��qfX�b�`i5a1+t]62QwU����[����Y�:Z��rYf�[��]�j��ďKy�z�GlK�3kUM԰�XF&f��%��	���+A��AһW8]1��m�h�ͳ��W	6�a*���M��Rf9�.��Ke7eZ�.«[V�B�BQ�M)/Tқ=�G6ZShBa��*�+���R���U.����+eF�Pi�֖�,nV�.�jȆX��:��L+�(�M+,�xն��T�SB�X���tѰ��њjԭ����p�q-��i�n�uI���%c���n��h�*i��,"X��2ۢgUױ��h� DLM�@�����.YH��fc�K�i+������!�Ј h@cf��^�L�f3,��ФF4R��dt�뢭�]N3gAbf�dW-�b4�LR�� �p����iqI�X��˦,R�q�悆�J+�+�\�k	l��ʫ��m���\���L4%Ѻl��ʈ�Z.��P������l���!�� �@%���57@�ʵ��f���*Ku�Qf^���b���D�݌]fS@�a�,� �aڐ�k�"�YY/2�cv�p��(��P�й�ƍы�TbF�h�l�8�ET��dDq"����jkM�5Z���X6ݫ��Qm�Xt��fjL�e��2L�K*��T4�dU�k6t ��{]�����tb$c�9�Rƙ�+ �m��ܴM���l^�n,f!id�G�I���bA�,��[+^B;��kv�Ɨ9&��ҽ���)��tI��r�s-6��p��ƃt-�A3�LJ�S�)mЃ
ێ4�%.V�ٖ���F�����Ht f\��.�gM4N��A��H$-�r���f��v3cHksL6k�4Ѧ�15;j<�b7D���7a��)uffp�k��ҏKcJ͜.��pM+�p�e�4�����e6�Ɉ���H���V�SL6�h���KX�W��]p.t#uf)\�i��Ek��\9y�&i�P�Z��Ym"F�4stntݹ�6h8 ��Djb]��͘e���2�uv�HPKBY����1ٙ�in1�4��k15�Vl&���bhb��+k��c��f����kÝ���.#/@�Xv@�XCWJ��̚�2BVF!���m�X�4n�ef�k�մ��� ��3!2�3�b�E{j��jBU�V%S6�4�`�A��.8t���#m�iָM�A��.�f��l�hT+��ܲ� v�꣫��SicXLms��V8�y�f�Q��L^eu�P�6(�u&c-������Z\���.��3*��4J����`)� 2�b7W<���rnƃ���ı-@���JC=R�@*��,��ƀ.t�B�]]���rL$�n�a�v�#R+
q"k�5L��Q�10��,dd�F3f�����s���8�B\Yb
��C.�*n�Kq���!6�uX,e����;�vIq�0�M!A�b� �ZP��k֣(;���x5��j�a���cJ�q+��l�[(ڋ&�a���X�0HmP���z�W�g)Gtb@��\ꚦ�@u�*M�����BKf�4�7]G
2۩!`�f�ۊ��,$[���tl��.tҗ	te���4�f��ն<< �b�0+,c�\�M��m��F�ݑ�F��eu4e0,�V��V,Vmn���.n�[�8���ѡ�����.�؈�e��Il�	ș�*�2��y�%Kj����k&mWq-X�=�M���T��U�Ҥ͠��#2m�X$��Q-#(B�ڸ�P���l۫K��R�s!��*3R��p����Y��6�*�]̰ĻW/f�J���J%!c��4��c�� S!�j�	�ƣ�m\7[e��{l�k�Z�#��m�s]lf��K�mč�َf:�J	�k6li����Xʺ�׳n��bf`�Bd�K��#�-�
:�A:�ͥ�a�:<.���l����+�][4�"�Ġkmj���t����v�JM	�K�mlAeȆֶea���^���1V�rk�-��ky�4\�	T���t�!��ۦBf��:W*�Iv�M�`d�8�-�PR[�8��f�Y�c$a1�K ��Ը�(�5��6#q�l�b�V](�p�r�9�l��`�[,���ڢ�0��6m���=j�����M-�P��Sb0�\3�ѱ�3��d��6��	�*E-ԏR��cј	l�˥ L�B`X���Ks��Yun���:��	�le�e��f;B�kMSZ�hRXݳ�/�GZka0���n�Xc������	K1��J��� �H\�����Qk��5cq.�.�0��]Ʋ��$#+�8م84��ݦԩ3�f��GK��.hf�چ`�lJ��l, %���0&̀��&#�D�bɂ&�ԅ)T���Ť'mqNԉ�ѳ �ĬH���f��-�.^���b�Ҷ	��۝(K+!��Ѯ�k��Mi��`�u(�chZi��]��W������JѬoQs�c^�E44t��3E��j��k�]͡A�W�t.
Y�5{m4v��hˍ���^�Wd�j�K��m�0;�+L�,�$��B	3Jړ��Z�f����7Vܬ��"\MR�c��:͋���%��Y2-�*hDȅ��1%t[�*�Gl�&,��F���jH�F4"ˋ�5���L�%n�裐��M�`DRh���Yj�Q�28{mFl�B["2٪�p�-��LK�f����R1����k�X2��(�.{M���h��&��\����3�2�pƜ#)����e�ܩ[�D�+]X��#��R��j��n��4a�Tٹ+�S1�uq����ЌQ:͐���ʶ����U�R!in�*,k���`&���muKf�2�-�x�H��NƌҲ�#�mf��rkfɸiZ& ���7]��X嚐ɮiX�b�q�],fR�҂�7%Ll4���ힼA�u���2A�G�;��%�T�W#o.�MR�r-�(��f��+a�L��33���w-��,���	��-]Ԍ	a�M`s�q�� �pV�c���E��-�ƅ)�n�F[p� ����u�X��&�M5�9�AK{F��Y�S&��Z��B�n���Hu�0[ ڲ�q�i�/iu�I��/!�s[��S�/lC��ia2E�V��i�B�ن�̴�ǝ�;R5�1�Q�6��[��R�2G���\�-�����۠�]j�0V�ј
+���K,q��6E`@t&F�7W@�1[��,x���%W6V[�(b�Rҩki��eKGV�e���9Ͱ6�����[5��;��]�ׅ^]���٩��@.Y��J�z�;bd�@e0�&�VS�,P��噥������!6n��c�օ��M�3���8V�4-v���(7�ĳQ�gV��f��h,�Y��V�Q�qv�.�%#�;6a�\h�B��L-(���m�Å���d�4���)���K���kF��1R��-Z�pck-#s͗@�CX�Ȉ���D��2��[��t4n��h�[��l5F6�.����itH+��Vc\�9��ɲKٷ%&��Mx���j᠖b�iMDl�6�*^�º��Mc�˝{l9���ƙ��ؙ���S�6��MSIp�l���a��cl�W4�`�6Ķ+�E#3�Q.�"�n�a��㛪k�D�XY�� ��ف�J2���]P\�M�9K��Ս�h�9�Z������.�e��dYk4a�D��-�V`�G�e�:ݠچj	qP`6���7CG[��a�Gf�]��$����҉u�ip�K��K.#]�U"���]�Y������p˕UUUJ��يd��)��l�[�9n��fU5�
�hG,�Mc�fU[����)�ʥ�WF��eV�쪪��������6,�BVƦ�_ưCo�]J@��s�Ϗ_<��r�|Ri���-&%`�/)ͅ�����#K$�Y)�5Ʋ#���pe��T�̳2����B�LB�J��±T��3�u1��J&["�1
�@Ʊ\ZR�kXV�YY��PR��)*��q�&P��H�m$˘TZ�.S�V��T���%j����UTkaX6��*J2Q ,�������X��R
�`��XT�h�� ��T
V�C-��*ȭ�������E��*UJ0�
��������g�Z����B�Vŋm�rڗ*�jAJ¥�-U�R�[k
��3
(��ȑL���!�8��Z�)�(e�T�\1�B�A)r�q�����)��f4�[R�"6����$�lߺ咡�l��cQ�R�(l�����jP׆�M�PfV�N�L:5��[���Ј��jd�Mv-ѣO���XS�.9ˋ�pR5��3]J�a�����;*�Fmڥ�"2���v4*f���A�\%��.�kS5D��"��4Ĳ�IHF��.ju��[��ͣR��//g���uqlL���s-IcU%vq�6�� #����	��#�5j�h�7�%���,nM[x`�5���ڶ�F�������\��,4*1[	be]��K�i��َÐo�2�|�Y���4�ˠᙰ����&�1cy��h���c�h��lq4�,/3m�j��#�X-	@�r\�Y���7 �q*�P��mZ�]�BN"CKZv1l��D�M]]@�ۥa�a5ѭb�c.�������#<<�p�.�%��V5�CP��e��4É��ͅ�!�Y��v��-�-S2গ%����+F5΋+�����CL��m�4fq�	V!��5�b�]Y�Rf\�.)pU΂��6ׁ��6��";k]f*"i��Y�i�s�θ�WQ��R��u�Rk4��c��[��6�h��t������#*��H�z��"�J"Bmj��]�@
�M� /c�3[rkmYB�ݢ:C90�	�Մ��@v�����BіY�-0���f�s]���fK�+<���6LRgPĺ���)U���c�0;J`(Kf��3نVђ�.D�A�Fh.%�-��M�ZBS\�G�	����b��[4�J2��8:�	��c��-�����fa�ɷ�z�QJG�`��K�(��ՍkfRcVP���fR�e���]�kL�Zf��,6����:��3E��B4���k:��k2���h����j�b: �"^Xi����1���ob..a�iv�-��(�.U˴��XX��]�*���D}2N�����ib����F�X4�%���$%�X �,�,B��!�[�שD�	V�T�RƔI`ӊ�b�IZ�Th����*��U�x,!X�u�VU:� $l^���R�H�j�/	IV�����e��jګ(�4�60��������䪖��b�l�F2��(V2�A�ÛVU�5�����mٜ�ĳ��fP�������w\�fmxؑJXA%�m���hМ$�:p]�7�*���c�ɮ1�M��j�s���^1��I#3flК�i�1�0��L'��� �ĳ��Ӳ'Ʊ��I�ڔfZ��Դ�?��wv;O�#���O�`I1ƉM��j��y�'m�=��洰g,%�h��6ā|�Q��HN�Z|]�^ �;���n�w��ׂ	-�-�d@'�5�͙��Kj�qyw�+
��,�3%��:2���F�j°-jWQ����ӠC"�v���)�x�b�4�ۋ��N���$�Ak�p��)�#=
vfH��� �������g"<f�Ǐ��,O���6�'q��Y��ƕ~ҹ�p�j�֟o�gN$������o������o�����`%�	�v�:�9W��5� �H$k��I �������WI=���k���sQnSn�����ߠ�����X����Bݢ�b,H���A>-��#dpDn��gD�p�맙�^����WY��>7��I-5� ����wuyN(�$i��q�H�Ƀ�v-TN��W���{'\ݳ�fs��f@�	$�币�Km냰�����,`aN�Y�.kU�ZZ�X�	K�m���tD]e��U�"h�W��G��-�J�����Bo_=0	��{�6.X�lpKʉ������I ��8�!�q�H?�ዉ���í �"ٝ|k�w�
�^-��#Ă�{�!M2�J���J$P& 5�
vR�5�O �Km�C��<ۘ��\��rf������gh��N������}��4�B��wI�t����`Z��&n��2��gM'��T��O2C#�O�,H-w��[/`z�T���$�:p]��ʗ�e�b[:�X'��n\G��#��M��&&���E�þa,�ftK'�MmLA �}ǂ�;ô���ɜ}GF�-��H$̸	��qp�8��8�!�"�]�H2>%ř�\�W�ꀃ��m���rhK�9�4U���|� `vb�iQ8�	$W��d�ex�O�6 G���,!MPhM(�ռI-U��-.�]��,���,m�|c*���z��;�$�W�A�9k��	��W��3>%��O��U��0%�%Fc��-�l0I�������r� �|}" �������3�5�O%;�x�4��t�MW A� -�qA��قYVSX���ٶ%�ն*���^���>�w��'������^�@��yb����%����)������;(�Lc2v�i}��^�V52��YX��� ��׀e��h˵(;�l@'�]n($����׀hl����,c��u!�AD`+#�p�M[��L��f�K�iP۴��Mc��n�_��������þ�k*b$N�m�x8Ip�jZ����	�k����H����'�u��v�'��F��M�'ānۊ<?��p�L?o�-?Q����ġZ���	��G��܆�6�.)�B-�Z\���m��%�5���%jE��gFA{�y4������v�y�$Z��	!��V�jm�kSD��G��0�%��������|O�m��C�p�,��<B�Y�v�PI �V�|I|�pԩ�����E��#idO����3���B{4M��$o�T����z�<e�'�j���=���䆆d�Z�dS2&E��a�\%�y�Lu�ԳG	l�Ұ#�e�s.l�r͆�׋, ;:�&
�k�lF0fL5�b���q��0Ԉ7;c	Dص��
m�bV�ʚVR6S@��%Y�[�b�e�d�S]s` �P��؍Ҧ�k�F	�)�˦o(cBd*&����gp�2ܮ���<�y��K�XiXˮ.��&"vZ�1p�m	��:��K�]��W`�tA�-��.�c+M5��I����3,����QW��� lUYlŬ�٢�V�[�#�2Ņ��YÑ`Qb��Ns�7�u� ���<�� �^�^x�}	D�B3SK=(�C,�h�'�͍��N]9f�[S�Qp�಴�mJ�	��A>/�� ��YRr���T�	7�E�f.�8j����	ý�`ӂv�+��i��[�H%�f� H-��{>���H���Z3R@�G}�-�9��~���#L�I>i݋�q��S�M�f�{�M2�#�E?�%�:3�*5�A���!�Uh(d�Q�`�"�l�A%���x�,�)^M;�dɛݰA���"A1y-tmE�����6S���+4s+1\Rm\Xژ��v6�k$�_�Ά�[t�I ��o�,v}B4M�h���Y����AUp"N�E�Eˇ�ă���� O�Y�oR��0�sS[�߳���H�V{Hh,*�cFM�ю�vwR3qf 9�cӽ�1[�ۏ�ލ�w�`�{BMfݶ�R�e�Z���<�Y2	�f�P&FL3��l:��}-n���t��0p� 9��M2�B65��+����Knۿ���٨@�lN�$K�b쓆�J'Z���k+q�#�~��>&��7��ߏ��u��~�{n!L)�������TAc�l%>N��I����'*v �!�ψA 2���z#�t�r�:�%" 5N�1�c",�ҫn���.@ŨWXF#H)K"ڮ��������	w.L�Zr �,� �<�3Z��`�*S@���O��5A9�"�h�ē�	�η��^[@5�q�����o��Q �׊>e�m�%�oO5`�/6F���K�;�����rK9�;v�8>Y����0�R�N����\��)�:��_���}���O��i�����RcF>���f���-�©5oU�Wo��e�����������V�v�Y�����7RL�O�cl#�C�h� ��n4��}�jY ����p�@��1�HGua�kQ�rc���&1˪yx�_ʖ��$��sZ<I�/'���3孺���/D��|˒f:������Z�ƌs3��m�Y��d��X��K��Fgׯ�_b:�U7�߻� ��2�	� �۹Z6���>J�������JLv!�r�{���n�� �@:TnǠ�.����b�؂��� �/X@$��D�M�����8$�@"5��
�����:��F����H+s A� ��u����x��Y��l�x�Sx�bY�;�Y�ώݵO�v"-3(��.�m��!OMb�1v��$�͈�A cfǅ��6K�xZ���jX����*�.���<�\=t����c�:〭ȋ��i������*&�.�v1;���3�I䠽�FH��`��G���wf�:v.�8wg"�>$�>���^<�54������H�%�6 	�����A�vB�r)�ك�`S:�t��L8��bki4�	�45[tn�Y5vX02etX��r����4�����	�{�A,��a�BO���HmۏA	�!9#�wsR@��y~\ }v��S�mѹ�4��-uq�oc\A^HE�T���^gW� K�rs�@�ӹ�A��I>)��79�t���e�W���~����o�'�$Y�7�v�̦�Kv�C��z�jTgT�E|ov"�� gc\@��[��wDd�yM 0>�ٝ����G 9��p8]k�|7%�f
�@ͪ}� G���#����^�k%�ܑ�N�3'�����}��ٞһg�y~�bmЊ���Yx��״��K���^�{u��y.����Z��%��_z��^���i	�B�X^���Z��V��tͅG4�Gg�`J�k��Lj"��PI����k4I\i��3:��kfr�M
,J��u��\������E�J�m\���x
���������f�f�vIc��9���kG���j��Ձ,�]Y�ю����-c1nev��kW)X�Z��kB�Zh4��щ�&LL�ؽ�L��tb�2b�\�.�]��,�t�+�GX��	p�[�,]YFVW�y�wj��[�N��v�*=W��k��Lmk�s4��R��A*��@$Pa�	�;��4�*'_�[Y�ܱO{��2 �̸�I �׏��Ո�__�u�~J��ݤ�t��<q�\G�D�O��٫�P�^��\��'6= ��ׂZ!N�J0%�92�܋9��V����ǂe/��ǀ$��Z�v��N�T�%�[��vM�p�3��i�Ēm�tZ�\�}*���A>1q�րH��}؏C&���/+F��E�&J3S1d��Ҳ��h����y\q���j����Yun�pC0M���V"Ȳr�	g3�w)�A���$������C�IT�&�`A$�[��z�!�y�p�;	����<#�ۦ|��'H`ٸͰ�Q��ɶ%���M�S������р������+{}��H8�Q�$�>{점�����-d�4��㠀D��h��Zw ���iw;'�Y�W�=���$[���Q4��o\A�S^1���wm�b�X$��s [/b)��7�pJ�`<�c#^�f��i�¬h!�)��$2�r6=��觚l��ư�,�V<Z!^�K�dIgL�*3b�_1ć�Y7Z�#[k� *b��$��<	#_6��×4�Ш{#�ir员�X�b�͵�e[n\,(����;�e��M�ٵz���7��.νU��H!��⼐'�� �v���-�')��fk��%�������:�XA���.�b��o
.A$�Ce�G�>%�6 D����^���4��q��.����9.]	�������ۯ�\��ڶ�z|����yq�q������q���q�ww���>|�z���������Ώ.@�#&�{�����p_"[�r��3��O����
���Ą4<�	�����=�Vcу55�=8�g��Z:[�O`���_	ٽ�TB=BZ��!��3�����a�Oi�6�=�n�w��t�C��g��e�g�wɋ�|�����]�xc�ؗk����#��>���F�c�r�|��j�طӗN����/�$��\{�w���9�����I<��;�K��*��?L������G�m��ԇ����D��a�v�����zŗʅ��X|�p�7���u�vr� ��;��s@�E��U����w��[<@�ӹ�1UI�QEed�9׎�C�0eZM���q%u^�����(�H�f��w!�;�9d��v9�r��^{�v����0�`T��-�*���P/)�������ի���q�7��g"G[��x���1w��0��q�5"w�̻�]\7�<1�<�MsU�v�'���X���7����y��{�Q�����'�w�]W�Ѕ��w�`�FŎ�}���_<��s\n��O�^G[۲=j�|B��)#t{�3�E[Bv��y;%���;�#\'m�l9�p���5u�,K\}�qO�o��=���V�!x>��8�X=����>|'	�$-��r�:�Z>ZJ��u�گh1otی�z����X���㞮���zu���y`s�=a�)��^`>����"�'��C:�>��g.�I՟�07�+�Z�mb�h��e����5�����FT�\j)"�Td�b�ԥ�h-�mq+"�L��\��­�f\��H��T12�S)lc+
1j"N嘬U@����m������F0[ZQ��!Q�kW혓"J�㌘�=�r���
+E`ĩDDj6Ţ(Q�5�*�2ƨ�آ��m�
���d�Q��h�r��Qq�J��*��VE�J��E����(�Eb �V��e�6�֬A2˙
,`��Qb*��كq��%���Dc��QJ���Y�u���ju�Zmkn�u�R�Œ҈�m��UVjE��XbfX�
X,EVօJ=��#5�2�(�Y�AAj,r��QmPHV���P�
%O�Mһ(��Ecf4A*Z0�6��2�Pƌc�aX����̹�m��-�m �X[I�(��2��9�����%�d)i�����Z��3���8E:0*P�i�H:`���G�@�MtAh˷~n����}�����">���'ޔ(2VIXS>{ޑI�%������q!�n����|�VT%��w�!ćM���F���7n��!ְ�����cY�������ؐ�R�'��_`�(�B���GFe+���8E�J�*@���L�G� \]�NpE��ܬ)U O����n�SutX2�{;,�̼��U�ͳR5�j<݆�J,�������.��?���*g}����T+%�3�߹�,����-�߽�k	�����������Ce�ߟ�4�{H1Y�{�N�
��OK��L�w6��~{����V��s������|9w�����y�է�v�l�:˿���m<��N�
�M2�~��:�@��	�������ㅿ�u���}��f�� ��#�H�E��6拚�ć�X|���A��-�� ����q�$+D�J0+���o�o.�sۛ��%�g�U�uk���<����j�Ӯ���ǌ���.�z���m�Γ���p�CďP�qv�����.��,��恞6}�}�O���@�>�X�8�������HV�����z=�G�1���.+���Ĩ�8���H�Ğ�e��l��;�R�[pd<.�wlal��8�N�Z��7��E�.'س��Q��o������ ]�w�S��������.��ΐ�<c��ΠT(�S}��΃'PB3߿;���䟣��s}М;����2g�h���:�|����o�>{��Ăa��´��P̵[4x�G�]����p�z�r����m(�2�˽�����fٷ�Hz����!��B��Yi����ԅj�&&
�����t`R<�=�+Z�� ��7":�A��{d�0I�y���bJ�_?&��b���I�OT�|�@��T*C�����-].w �ஞc�|��"��a�0�|��u!��Ad�6���t�{g�(�@��y��j�+�r����C��r������@��'��
�(T�M���!�:��T �s�m\	��~�-�9N��ȏh>�V��翽޲v!P(���T�}�@�u!C����*廦7^��,.�� ud1��շ����H��x2�V�B��
�|��N�e@��g�y�	Y9Ot��y��vMd>$�w����g�o����i�ۦgH��O�;�a�a�Ad��~��Ǥ��ˇ7'mTN؊��H�B#�{|�$;�,���߿i��bB��Ύ��D������*�M�g�eq��)���13�����}�ñj�˱yXl����.�1'��Fr���uz�`��VDܢn�m�j�:up�����������X�h���/��v��n��:H���+���	w5�u��	ck���!�-���a�h�6YJ�m^M6�̔3pv�Z�Z�-�G6�ڠT+�=�������j]Z=L��,��2%��h�)�Ԙ�V�ٳR[Rf�X�*Bc�V4`1����P"�1K��V��fe�a�a]M�rnq
���=J:1
f��]5˜�O[<�e��5#a��(��貦u�kÛ��ԛ��Æ&���������.빟�|H7{�g��@�VJ�翶u���¤�)�}罁X#�||��=��3��|�+��"�VJ���bu!w|��24�R��{��������8�)'�=j']"'))�Z<Lt9�<Dx#�����<Kμ�u�gV�z��߉�-��m�7y,����s�y1',��fb�u�Ğ*g}���é�a�c%B����ܝf0(��R��	��m��,}r<,��x�0,}��9�?i2ԅa�o�%N�*]��+�,����:� H��vC��:��T����~YbB��7����:�,,IXPϞ�ޒ��¤�+<�>���s��>��vH,����a VVAL���C���?y�Ust���Ra�����Ial���/ߞ�YϚ�������)����u�Y؁YS<��yG�d�Q��Dz[��τ��@�{7h���E)�Y��B��E+m�R��G��i�sPr�Ù�X�#��d�+�����(�6�o��w�:�_<���yYyű�WYv��<<��E���{�d����O���d>��o���ZN�C|��xJ�>�|��e���w/u<�y�5�@��3f���_Ow�3���
��B"��i1nKeRf$s6��̇�''#j̚[un�&
ֹ{%��+
�Jf���&f�ܛ��u���������2u
2V$�)��s�IRv0��c%g3����A@�*��Kh4������lĸAG�w��\F��fc��d���C��!KI)i_}��z���d������.T\C�Svf�>�$��#�7ls��W�j�j���nsߎ�y�u��y��]m����x���L��2�**r)��{Co��x�I�}���=��
C���y�� �G�	 �����Vg&+�G�x����C�~s�	Y:oO����w6������k:�YP*d������I����H��7���{��>�G���ϟ^=y�h�y˭/sׯ��ū���>x�D?s�$'��.�7��6�r��穮����l1���E]-�M��Z�11h�p��Ek	��n_��׹~M�2ĸ���{ݲ��;��^wl]]u.�֞�^�sƾ$+�%L`T���xC��;b=��K��Gj� �qP<��S�Ld�(�����k��>O�߹����Mn{d��<�}{Y(�#�H/�r�a��B`|1�����>ĩ���{��dAM��C��R��R�����<��xJ�X/�O{��n�n���3�{�gbd*E��{���O#> //cz7�:hgx���Q�\�՚�2�r�\�1²D��8�U���+�JL-]������>-4�+���,Z�����Z���V�ڦ�O�Qg߷��o�?p�'�
��*Co�~�Y:!Y�D����Hq!�w�ަ-1��;K�>(�6�� bw�����,�m!����עB�Cȓ)9�p�S�
ʁYS>���R
kY�*�N{�@����3gl9�%a�����\��u�R���	>�}�O�,�O�zH��X{����؁�ć��o��R����:D�Q$�gt����Kn6����Yl��,�8���p�R:��.��Z���K2=�6]+�X��ō�m�Ϲ�|~a�nq�o�s���I�v$�I��f��'ڣ�����.;��T���%�O��$J�7�pf$�wS�
�����@uH�5�.�>�H��@$��dL�$<�-�A��y@$�̽Ӕ�����V����u�	r�SP)RWՐ"%�f���^��A 2#F����̀hIyw��ѽ�&QA%��&l@��AI�g�P�L�\�����܉��J��$�Iy$�:@i�D�[��G��p�ٝM=;8n����~z�!G�x4u��-��*MІ����<��<��/t����Ǜ��+m�gLc��&qd�����N*��u�N�"�f׻�G�7א'ҫIg�J��l}Q>�y� Z��~>��M䩼�'"F�a�$�/��L���r܆��>E�w�ebޭ�۹�)�'$��h��F���ˊ��CF���Ga�Z��ʚ�ګ>���=��0!;�zy&���I6�ؐ��fI%�-2����A��D�+���E$ػ#|�כ�C�c�L�K��'u�H	���o^�1����ϑ`�Iy$��ZR^	/'n�i�P	 �8���:Y��2R&�,Ē���cUJ�ėI$����@J%>e�wl^w+�F����4z@f$���Hq#a�q�N9LQ�S5]L7h7ښ���ͯ$��W1>�@$����BD���UqA�.�I��MM�->@+#tRpY�w2$���r�D�wD��O�1\��e��y�)!4����	/'n�i�PI��"	���l����n�ל�b��m�y��Ֆn��8D<0���Q�h�CL�{5 n�J�,[���A��M�f�N,؆�0���n#X2�}�?=~7��8&�2�aa�T5ĳG1��F�+m	�WV�pچ�a��#Y��,�#��j��X)p����K1���8I���h�P*]�����흌�M�e��.��X4��a�F2�*�fj�hM��D�BgM�Q�ێ c-�%�t��藿�0��`[*�Z[�`�Vl�Pn��eKPl�cգV6��Yt�.v���uk�b����[%Ț.e�3m���FWcM3����b3>�����0X��ao��[I$u��2�&	/4wH�	v��&��s��y�%�$�I�oZe(���ĦLĄ�A�����D���ɽs5y��<����J�5w4�32:��$	E$}\څ�un�����0v(�gPM.�l�J@.��)/$|D�7^(fmc�
5�;��H$�f�ƙD��;�L�s
��I,��5T��d�SK)��Gwu���	r���JA$��F􉐒	&]�.|��6�ݤ���7F� gÝ���'��ϒۛ�RI&7�!a5\�V�Ԑ����I"��Fl���H2��y#��F�K����)��aD��F����4���G^CQ�v���)�����2��1pY�w<+�4V�I%Q���)�wK�	��܆�m�^U6�%�F�	�z��C���2.�e1~�	����Ӯ��|���/�8��3�����.T�� ?))�w)p{\�����L��w'�V���.�79�r�HXY�
f\+�>��<A}��M4�Aw��}�&Sy�̓.���׹��ݢ5�T��ٽr�m���N��bə �g񪠔��O���I�f��I$����Ǝ<��ݶ�Iy �Gl���w�R��ݝ3�H�gPeSv�G����GDvma��{�TND��58I�S-�$f�Ə�[�v�\�T�;�Sw� �	�<Ř�Y�9Lj���VK�	$�e�G���Sю���.�e%q�"I��+�$�	�w�	�t��cO~��D�X{�ź1���b.��m�ή&k�e\��k�W9BX����w�6\���.$��G��Mk�$:q�']��)�q���|;��7ҊI�Ζ&lD�$���(QI��)��TSL��]�OE�e$�U�ϽM!$�L���Ќ癀�Ҟ�.��橇��D.�Mw
\��>~z�0�S>~>��nH����ԝ��][��X�7l��TdJ�A�U�g-�0�l���|�5���q��M;	��k����OYH��̬:�qR�p��>�@�H�����`F�I{]�e���7o�2�MP�bə �g񪤚{`�ӯΣ�'\L�8����$��	�;Ze$I��|:n R<�$���e���e�\����쭙��AgRd*n�i�����wE>H�ȞiW-V�>EE6ܴ��,�y���y������}qBH1�.�E٨��5>��K�Z�B�*����Rݱ�3�Ev�GK����f	�O}�!�%�wث&]�L��� $�O��"BG˶v�-⒌k����- $�^L�|�)|N��A�ӰLI�����5�@�J[�����l"P	&j�i���D=]�B���>��d��u��D�K'$��N'�i3=kA��I�$^I��3�+/B\j#K�]��I2��dH�����C����2.�d'/� Vz�gn�%�Lګ��RI$��	'�wC�>�0�o��>�Ǭ����i�F�2	5��4v�7�g��dm�n{�7���	�\��ZE�gf��J�R������������1�����)"��D`��?n�>�ΉK�L�LY3�,�7w�{�'Ȥ����0��Ǧf�=U��kY%-W-$�H'���E$�{�;��#�ƕD����s8�ڡV�:q��U�����Vh��-b���K���<��� ���<����J@$����I�%j~�y�Dx�dd��s�X���e�Q^H�f��%!^�9�\�;�)���q��H����K��
��=)�Oא �Ij~�y	 �^j���O��c�c��؟tr�0:`ʍx%{7%$��Ή��3{��f�^�4����jI$��$O���m�iIQ"�I�%�r]�38�vfz�-�V�^���L�d	|I!��������Lݼ��qV�OMPRK���D�Kdnim��tBfE�]���!��@$�vsO�v�Z���'_��hI��>I$�!�SzC2]�f���)�^�|���_/n��������OL����o��U�B��,/x��v�&Q%IsMΜ��&1˅5��7Y�0�X�a�X�UZ�{8{=�{���\oׯaj`��a�V�{���������;�`?
�B�;��6��t}�a34`�U)'h�|�����,tz{ir;��N��3/:��=1���ؤ~�%�򾰻��G�OjǛ�z�N�c^,�G��ov��y�>�6��&'�W����X��}����{�[ʍ{�`��ub׆���~/F2Dƭgxw�?S�z�{ۃ]t.׼z�r�w�鷅�����������M-���ڟ��=���r�3:^ǹ#�^�{L�ަ��|��8����Q+�L�$=讜��9=�e>�Huo��S��y��uD�W Œ�)4��s7���`���_��})k&�Ω��wvk�YL�{�l2Q4s�xd�Ņ]�|�y��syA�-�7F��3��x�_��5qf>��{/�{/���8{6?>���e���c�˚�ګH���z�o}�!繺��Q�w-*Գw��{/\JKGg�W��G{�gޚs��x60�W�ǈ��}�ѩ�W� �{�Eu�|�0w�vʮ��՚�����=�G؊�}� �����<����I��7�}L���=�� �'��f^� r�]&>VC��ޗ�3V��G�&���y4���5MѴ�ʚ���<^+x�#m<A�H(b��w���<uw{
u�Gwr����a����~��[�w�7�.^Ɇ����Q�,�7s���f�V�f���e��[�&4�z�UN��\/f��)@����=�&Q��맙F��(0T��0�e;�=�5�����Hg�_��3�~���y�\w	ш�\±-����B�h\��E�6�Y��F5�[�����mc� x������4TP��E�մr�"�JS]�¢&���\�+��uz�^�aK�P,"t��ݜ���Ƅ-�hq���:�,�d��aN n�9��EV)��+[^'����`�Yd�	=a�e���m	Kh� �F2/�d��y��[-l�/[aKP��X��ۂ�&Ĭ���3�#��,XDV%�P��[��2S;eض�KET�-i�v/��1%��@�Rq��rR�`e��iTQ��ip��Q��qB��ơ�X���KM")�����cZ�/2ڈ�e^�U�r*r�e���X���M�'(U'�0*�J��1RڤU�1��cV9w
(��V� H�bՔ��:%�(@╻R mql�k���  �l��kR���w`�K̝f�2�Uf��J���R1\reY8�6ngQ�.1EM�]h�X�J��2ңam��F�������W+�5���UEA��EDQ2�fs1R������|������gi�2eř����U�S^�v ��2���FM	@��:�M�6��U;.,�̱��ZE���;E��n��a)������ô���B�6\\p;F�ŷa��fh楩I,�X�5tV�vô���!X.�mئ ��ݭ��e����(�"ѡ��[��H��e�:��%�
0�� h�!wg=wA�;1d�$�MQ��Ո��L첸�V+z˝�6�%�ű-Ѳ�rX�s���F�ᙳ7Mt����$F3Z"���M�f�a��\�IM�<����ni���٘��B7m7X��S�7z�6��6�;M�\�R��Fk��Hu�*%%l6�l6Ӫ�%��f��^i���X�h�,E��m���[��f��Kԇ,�*J#.�&�V���oU+��ћ�^t�5��e�T�q%[���b���豸����Y�`$��nY,й̴�؅�0u^F4�X�	J���:��Z3^�,m�X�%h�Ԧ�6�L�)	fc��j��.DY�M��Dy�R���ڕ�f�	�]+0h�G%z��G3`ݰ����<Au �&�ja��[yj�E�h�ʘŎ�m1*��P�X�up�	�n�Z.���a0s�Maj���7$�n&�6e�,J��\K��[��I�a�L&h�aл��5���ݖ[�:]���GK2:e��Y�(`ԙ����e6�)u�"@�2�4�^b����+�3qM�����E�����W�W8:��� �F�1�ю�LB�v�m�fK�!2���Q� �B�sY�h�*�a��Lk��3u
�F�h�-&���F�FKH�A�vuLf5)�p3]�(�,���"IX�����ut��cBb$�M@�<h0^r��n8b�6��m���T��Ґ�(���԰�u�
#��U���1����X8r�Lƽ�hW4�@e�qKZ��5�me-�t8]e���6�˂�Wer��L~6`�Ϳ6S�ŀy��o�=h�U��V��jl5���1�s���n�.fkn���B�A6�Z6��S$ԕvػ��a���j�A��̰�X4�a��\\[��V5� V�$y��N`ީm���a�K2�Uea5&cM�5L���c���\3L��Cp�.���p]@��9Y7B�!�]l��Q��\q-��Mt'������v���Pt�e�f-p�:\��U�ͳ��C�l�l�:���a��҅�0gf�$ٕ)�&JA��D��Z�E�����1�������U�-w_��a&��!%�a�%�	$�osD��
�X�k\�fyGUH�e+�m� $�0sl��AgRd+n�i��4�,|�TD�k?��rb�d��l>ʐ��c)��}(������!M�>	���%�0 �p�1����Q��Jv4�D�����ط��زp�\>J�I%��FF'CC���:L��U�p'�۳�i�Wh�/%ޞ��F�%Cu�L��0d��z6|:��߶C��$'��Q28<��Ӻ�$�VL�4����_�0����O*>����21�}�ġ5O2���P׼�(��M�� �آf�a��m�v*����Ko�W]l6��PxWH�e�����6D]�lЋ����]�׫�4�-�a���W�&C �H%3�e�H7vȒ@>xt�������a��Ғ�K��ZeC�-LX�$,�34�Ol/�y�/�M��3�vB����^K�U
�Ed=��ݵ��I�/[�M[�v���Q�p_+��ޖ��M~�����us"Z�|k�SG�����i�[&Ҷ�+5-�m-����mSj��m�m"�*��:%�5�4�)/�}� �}*�mJ.^ؔr����$��!�Z�9)���׍"R	$��b@2�A#�kz������Ԗ$�Z�Z}(��	��D�K�[ioL)�9Ln�G��@��oL0��x��DY=����i���^I����e��1R�OKY��/8���	H�N�A��t�3I��f�A?S6r��C��S����|.�Ēz�y��I ���L�ڣ��$}S�����<���e�%�)��fm��q�P���ڕM����
�Ɖ����^��v�퍙�_$ϖ�/�o2I=�ă($�I[/>H��9�dGq���AU5O2�����D�U�]�tS�L�Ȼ�,u�2�M����r�t�-�na��3��)$�>���'�!���nlTsԤ���X��f(�Y�n��4�D�I�cba�X ^>^��w��r1]Pt���'�s�m�-��ˌ������:̻�~$l4v�Ԭ��=�����/e�;&�:2M��Q�=ŴV:t0��� {��zkm5[I����T�{ďx6=S�� �mߠH�P@%�c�rf�Rhe���P.��RY��M艭�5���f`���H&HI�-���$��1��@蹮l=��������)l��ɉ%0b�N���%�H��D#��l�;Ot�0	_V@�y#C�Kϒ%%��(�#c�!SC��F���H�8݉bY�4�d6:��j8m�ī�f�G�\�%r���t����Γn$��Gx�	g#bD$��J��e 2kLny���4^���(�$�dl��a�833.��3�I�:�e ��0�Nv���~��W�D$�lt���Izi�7���Hm��$�4�r�͈7���'p��"������ו2���"R"O�O�Rj��tм	/$��zX��E�w4z@)?�*�&,Y�(�r.��^{`�����#�ؒK�TĹ�)$��f��	$0k��x�����N���Ȉ��aa0l�"��۳D��),���-4�cc?�~�zg_�c�֬;�q����yu�?7�?�'�$"�dj�j���h�-�a����iS=m�u�O~�}>|��Ϸ��X�L�����mkY��D�$ۻd�E������.��Q�RQ���)n�i�II��D�P���Gl,dfb��^ieƪ\�J9avm�h[��k\lJ�MV�Bmt��nҾ.���������[�A�	 )���)�	7^��Ĥ|j�5'\�V^�6\���('l�h2� �%���9L��P*�n$$�f��ǫ�$RV�	�(:I���L�H��
�����*t'����Y��/Px��Μ�"��
)۩X�JI��'�RI"=U7-;zT��UV��A>>b�W���	��D�H
x]�.��L��|���v�k=��-xK���ʥRH$���4�zX��5�2u$���H�����Z�1f!$]�7w�i܉RI.u��@���l��2w��T�r�Iy$l�� J)%�������/)he�����s�^s����txN::W��t����VDn=E{���qwo���=*���}6b)���o��t�p�^ef\֮�B��BAY�mMd�V����7��h殰��m��t��0�7\q�^�/\�1�:Ӕ����c\�Z� Wh�դ�4ī��,)�����#	
3XYnY�ZP WR`	�\<�M+�6Ջ���
66騺kf�i��ki]�F��*k�f1�u���J���*�^��e��[�Im4�K�.�&B�T���pB��¹Uԓlp���2Y��y��@강��:�f� ��^c�s��a
�`��I��'��s�d�	ؾ���ި2%�v'�RI%���ґ���*i��3����~�"Q^I �sdH����j���.��˹��ڲ匄�����Ǵqv�K��B�^I$�n�2��u�-!"O���J�`Ć66gR��ts��ggL�0f�!*鸓)#�U�މ�Iy &Lhf���ۖjH$[��L��fK��,L�>�����fE3�c|�1أ�w���,��S��I�2�L��K��%��I���g��XE��� �:"��HW�%w��N�X�%�U]$�I����Q�3���s�^����4̤�K�%�$�O�ܠ�3��U�����`$=��/�����Q���kS����-�(mi�a��AУ�E�_'����i�]]�����oҥ$��[�.� �_�L���l_f�Z��x*��3(���k�i	(�G��L��X;�o�y`�H��c|`9;��B��I�E,wgˆ����l�l���E���e���y)�w�9ڻb	�����,�Zƞ�nohl-g�Y>���Ǐ��=y������}H�ŬJ�-���J�T�[QY�l�XV�6�h�d�X+W^�W�'o��%y?��)�PH�u}6x�F���&l-��.�×sUAW��X�I'��S)$�>�7�v_��Np�	$��v�H�30I(w�R%dc��gb���YA������{��n��a���I'�Y"R'���v#��c�@g���=����.'��t��Ok�RQ�;�31vLȦqb�4>ڟ	I"Z�bA��{���g���v@I�T�JK���PL�[{`O� �9N��PIl��2ݬd���s*2�3���j]��h��{]�����߷�{Z�j~�m�~y��32IG6�)$�M]�"R>No!�,�_IǶvΖ�$�H'��PdCɭdX�b��]����{bA����H6f]u)ȿ:^�3�-�T��@W�4Ge	�I>qGH��/^�1^謍jI�K��μX:/J��^�L�I6�ę�?��Β@?���Q��X%Ay���BE�l�u�q�N˸��Ƒ�ʆ��Y�K4��v7��Q���ͳ�c�ݖ��ۛ���t�;�wn�֍?��$F�S5«j�KYCZkUS4-�YϏ��>;}:�V���"QI$��șS8�r�d�˹��ز�	��Nٽ��	��[\�@$�y���D�H%��Џ�'3;i҅Ʌ����$��|�!K0�6�EˇwLɔ��U�p"RA+}n�@n�B���8�L���^iL��I��D�+��ϯҤ$}x�;i�~�����h���'�>�ZDݴ)�ѷe�ZUZ��\/30 3\�`d���{��W2Aآ�Ɗ��m"Q$��D�)*�y�tk��H��޿fm\�,�C�����(���t	�\��Q`�8bȗuT���e$��oC��&�D��I+~�L�+�h�G��WD�fw����W��Y.]����ͤ���[60A$�>k�3�Hg*y�Ҵ�3UP"7ju�pI�[� �e{_z`ϒ@�����μȺ/*U�m�{v���PeWCG��훊2J�T���	]��/G�o���$���!�Fe]LK�P�T��NL8�\2�ؔЩ�̦��	��g��5��WWǴ^��O��ɕ*�����Ji�,�ȏ}���xKeM�kM�5�[*[J��+b�6F�[DF$<W��=��ӧo���{����8r�`UXM��2|� ����d}��;���ͬ�$繁�y�!$�ml�>�|��xkT��=��.X8t	q[1H�P���Z���V[������&ln����͙����ħ`���2e���ͻY5�+�~���F�%��J@U�*�޻-/Q�"w�#��N�B��A��]� �QL�Rhz�2�G�2�%������$($�T����H&��R%�-��W=�: Ш�~��N�A�Bw��D	@,�3?4j��A�p�'ūi�����5+�H$���T���-͜�R���dQw�;��T��LΫ�%�OWD�Y|�$�	&׾S! �AtwO�tNc��Kt�3i$�d�J��2eb83��'E�O��z��y���]��y�rg���*BK�$���D��H.~�2���������KmR�c��k����\c���{�7�SsA�}�ƭ�9n�/���Ղ��6�Ғ3�����,�#�?sΘ�f_��{s�����wwW�@��[RkT�[�$H��\�.�ۙ���U2Z�F�����̈́Z��il��4�!
�.����̚l]�	fÇU���%�
R-��s7:f�6�e��PνV���&����j�1ReXaf�4Ͷi��� �kMb�L;,� ��e�-�M �@)�B\$�\�e-̢i]��[f���,ìKK�,j�0a�Ѵ�1t]��1�l�	6� ��JUXm��sR��Ff�p�ur`�c+v2��_ρ�ؐک���_Sd�JR|n�3>f�Kc��|fC���0�c*��hH�s��z,>x:rY�3&Ti.�{�).I4�5�v��)����Ux�~v��)��T�I%O��D�J`^��R��T�%='+Atȇbg ��'��S)����ϒ�b1v@�z�R�H�7ty�$I-~�0f�zY��!�@L��;�hK*��yE��$Nsu��LI,ϱ��D߭��~�U�5�ln�2Ƅ�]��ʇ�8�"��'vS4���R})�~�ؖ[��kg�9���&w�S>I�X�g҉(7s���6�dl����J`��%�.�t�e�C(V!���if��Cf
�3�]6Ιf`��&Ѷ#:�v/����L��K__eJ	/$���҈}��O�#��ԧ'�>m��R%4��fR��	�p��CL��������}�F1B��Ô�7ݔ��_"]�V�1�̥3<���7�q�����k��H��n�h�凶�;2��ۻ��U�^�N^���	�c]\?  �@��,�e�Sj���Z(E� ���ϙ�o�����r8��$Jn��T��I�^�fn{�g�X%>���r��($��թI���!�	�*m�֪�8�Դ�H���I��~�L׮qW���$�,]�4?Rㅲz�8-'2M-n@$�V<�'�A�+Ѳ�*BH����R�xhE��$tGg��2��ȇg�u2>�̲A%��sg)�Zy�b,�x���$���$>I5s�	$��s�)���z/|�����ۍf���ncm�6l�mb�׫t-��4�)+T��������S�-k�(�����M\�!JI$ݭ�!�
�� ���d$���͡%n;�7?z~;�W��1p"z@i�I2�1�S�yR���H�I���ɕ�e�S��JR<��M�햯$���m~�2�	L��d�-ɬ��a��zRye3`b2w!���7p�u�o]���Ϛ�n�u��yqǧ�����ӳ�=��g����{<���g���S�ʙΧ���8i�?Ǻh#�9zԴ�CY�0o@{@��M�%��7ٽ����;�; ���J�XfJ<5��Ob7R�d��`��mW��8��E���g��n>>�o�8gK~{���}�w#G�N��������Hy�x/)g��c�O=�m�B{ʻ���/�{�g���t�=�T����>�$���H!��7���^��b�
��0�k�Q�5����M��{s��#�X�3kʟ��/�,m�-�xMX*�,�pw]8;���^����Vx�v�<Z�<3�(���N^���tws+�|9��c:��{���E}�6ę"u�(/�ؽ��Q��%X��ٞ���o��Y�
-c�͎�ov��tb�O�^�-^��$��i7�<���)t�d��:גO�����v�!%����y;��8͵��|s�شeK�K��׸���87�b!�o��9V1����w=���r��5��g�'�U/;����Ǉ�..)��@�����x���H�I=��Θ_��.�Y��p�ٌ���9���]^/�[����eiY��3L0��7���.ɇ���ǝ����
�=��z;}yIq�&v���
MX���Ⱥ�ܖƳ��^;��۾�j�S�>��b��c&�٤�;�u��NkS$���^�K�����;��x��������S>�V��c� l��<�_z�d�X}����s�z3��ڹqT[.��{ю�'B�@@���)5���S�xg�_��4�i�u�ẇ����T?	phbX�Y(�q�P_����T��h�n9KH��b�.��]o֞TbR�QAX*.��"v�n�ELY��������r�*)�J��B���J"*!���Ê�Q�Q1��J��UQA�j���Ŷ�\�U������Af���RTpDF3or�,���TEJ6�iA��6�"1�(�]ʪ�r(�1Lh1H��*m
*��]���1��^YX��D��N%���i	na[h嗔�m�핁��r�Qg2�Q�,u(����T`��N2��媢1���.�Q�"�b#��E/mQy�*�������%�Ƣ�TC�]jjfS+LI�%J ��X)v�<J�UC-yJ�b*
$D5̡֯)DU��Pv�F&�1�1b����-
�iE�"�ܣA+3*�QTEb�j�j��a�V0U�,�9RTO-F*�,Ab ����$�(��"�`�b�)R� �cUA`��r�U-���b�
(�
��-��KZ�[�TE��\Q����-{N�f�t�y�e�u�Z��Dڈ��)M�Vқ�%��=���%��3y���be$���Pe�6Br@�:����_��ݛA��f��˳R	^�ȟH$Jm|�2<�)s�q{DH䩰�gRA�e��lZ�,���)�H�	����A"m��T�k.�Il��XI{q������m|��I,�GK���-�Q�UF �@�\����靂tR�P!v;fĩJi.���MW0���h�ˁM��k"܂.�3�ɐ�$�ml�2�����d$�V�ә���g�M�{-)$�j~�A�>жI;8r�w[�J�g�RLY�"�n�lS�k��f�~�5�$��1����)���(��1��I&B�#�b�v/*|��L�'�_d(s3$��q�2x�k�>�$��~��R�I-~�3�@!�S6� �N�3��
�VJx"���T�$��F)��I�3��3!$��swK~^�w3V�M���f-�v��;�3ϐe����`ٶ+�vaj�:�U�R��XiU��\����!	;鲋o�Ǯ������kTmJ�D[$���^�g��Ӷ��W��W���ՙ2�a/�^�)A#�SZ��C��A�k;<���s�)&RJ���)$�}~�j ����"R� �5�vgE�
!���6���Y�#vYH<��ࣖ�S.���h%��~���|L��]�)�p��y�� 	K�$���T��J|�����&��x�{�k�)($�=�����C܂.��k�λ�] ��T�mke��m�j��RH��q�d$�v�K_6Hx�Dkuf5\+��>P�Iٜ9r�����T��*W�I?�uz@��I��n��\�	OK-$�����I{����$`�Z�XwLQN��J�z�mb��aO�G=�Io��b�#%$B��e�"O�#�ګ�|	��m�bK ��0̔��we3`b
d�C9��ز�]$��|n�2�&:���.�K=wo�B�"��K�+vݖ��I'��S�G�����@̘.r�]Z��f�Ä�5����س����u��cIF9lW���	O"dNLi�l�c.���=�l<8q㈰�·;.�'K�G�w.ڨ�)K���$Rww@��:�'�|�2�#ѣ�SC]6�������G�f��(�a&�.3y�2�`Rb�M�.D��C�.F���z��`�Q�;d.(Y�kevr�P8-�m6De,v��-��l�P�@���d 2����֚Q!U��+m��A�@e�[+i����2��WM�R2ח�C�2��a,� ɡ,�i�%{c0�4CK�틹rrD�;I4k̮l�qC&�ka�L��V&�ܴ�p���K,6��a�:d7x~�wp�|]��>R��7��]1!�(�~~�2�V�[_#�v�������a����mL��]�)�Т����A&ۻg��jy�<� �J�_CJI%����|%��ڨd'�����}�o{1u�D�ݽ컷����Z_#G>r�%O�o%s)E�ksӵ��PDV��I$)��ZBH$���)�����ɑp� �檂M\�fxe�'�N7I��t4��3y�sd$����3�GuU�.&.z��c��{q��$��#Y����ʟm��2�I&�}�)�1)�w9�L�u%�OR�$�I;n�L�Im��2��k �ã�"\��V�c��1���u��\�������lJ�L��A4���S6� �L�g9�r��y��
�����RI$�oF���G$p+:��E�n�بx=䗂E�_4ʃ��c��.��(2���
PI����z�N��k����^�ss��{�r��:>�|��Owee�*{��0�����)	�����~>.�
.�g�u�x�Α�el�bچ�}�P�N#�w��ݢ����鸝M3q���ԁ�HIH&�>|��[mP������3x2^O��&%$�:Ϗ�x)��K����`�b�w9w`��R�{y	Kn>O���y�2��M/EJ�6�����D�훍2�	$�ѦD��O��.]�!�wQ>N��/�=����)���AM�QL@��O�E]�ߙ�%9P"A *����ǜ�/&w��"ki��DgwĸrgsvJ�{�)J���Oѯ�4���$���HI���ʿ&�{���%vb�]l��	�C䜐��j��
��v!+���GZ��m��`��='ͯ�]1E8}\�E�I$�e�HR�A)� ��4e*6�h�3����]8�!&�3�S�i3hbJfg�9��Xlȷ��H%,�g[3ϛ[��	 @7dY��H�36wD�	$��5�,���saՂ�`.;�t�I5��aJ	$���$�I#���sUH�yS�5U�o.�"zf��q����k������������}��r��Z��h�>J�޹���<v�;�M�5��$\X�+��{� <������I&����E��w�D�d�r6�ٙ:)آ������`qlҔ,!�[�$�?=J�P	!O�e$�����1��f7|��YdJ]�O��r`]�ϒ�lD�$�	�g.��3�1Wd�CэI���"L��A.�g!S�0)s�_<�|>�<t?x��E<�%�3T�.�E��` ��`[��J�{�+�ȶ������f��Y��|����T��[��Aw��%�� @Kve\�b�>d��K�I��ȓ)/g�̰v�v/H��kJlLM��A�ab玌j|��i`�	-�ȓ)�����P�2ӕ,���^���5�q2�Ĥ̟��0Ք�$I�h�IkVlG-�ֻ#���HVGD�H��w4BN�~�\:w��Mz�fn���j@�N鼩Iy'��I�@%���K�6�a�G����p�\(���Ĵ�E��Pѓ��拄�=y�p���ڠd/o9�%6f��t�8�Wuv����D�н6;������ ?�侞��L����vfN�v.ɝ�A�c�l�H$����	�7 �aؖ��)Ne�e"v�`&ތ2&��0Pz�3�����p�]ٙ8$1fr�@�I�M��*�K�����m�����Lզt��z���rI`]�rȎy�S2I$y��I$��$%������e�Lę$�(%]��zcx�f%��w=��Z�#��:��ݧ�6ncm<ZX� ng��H���"D��O詺� �vi�@0)�h.�$�^Q9�!#�In̉�Im�q�mU�I �^�B+�$��"|}%7�8�e��A�3��ZU��S7���&��n�I���	$�i݁�+_z$��U1E�U��	z�`����9wfTi+���)$n�x���-N�a �얈Iy?��g��L�$��L��0�ٻk*����
j��w����gv�ʏx�<��b���=���|}�r��G3��3��/zN���[�V�f�X�L)֝�	����k����f��h�(Z[�����*4��� �Ғ������՘5�t-!�Ί�F�$��cR��ր�5օ3t5�;���ԕ�`@y-�gc-ifv���dx��;&���)՗K�E��il�&�e�n�GE���F���4�1+�n�T���v�g��[T,  �b4��6�MnCbi�bD�;`5p�ft�ٍ����VZi�.��	�-l�&[h���]���ώ�:Iػ�w�Ɇ�s�H$םe$�I��$�S�ׇ���ie�D"�Kɯ�|&UAn��AÂXu���I����]b�nh�%{��T@$�ttI�$����c��覸J�vfE��w5O�fzΉ2��2=��	x������kA��ҩ�G�I͸(�#���e%��H-F�3k���N��QLo^�P3K�r3�$��M�t_��$�H�U|ֹ�݃>X�$�~W5�&Q�ޛL��H2O�s^�-�BD��v3��4�1��h��&�t\��$N>���%f�;2��M1���L�;L	�� �A8����n�%��0F�%\��7U�U���e�YuHؙkc؎c/�@{\��o�{��I[�<HI	�^]��;�Z����=T��P���<	/5��2d����3ЪJ:�!yz)�mk�d�z[�M4�SJ��)9w4⅙�Swճ��b:��"��S�$T�Iҡ�&�tL��oByf��"审�A�e��������#����d$�Iw��`��&�ȴ��VWV���[d�(8pK��Bw�y|�	$�g3��32B��5u��Z&��	 ��d$�H%���=MnY'��̒��ګ7�x���'��x�6��D�&�h&<�����>;e_%�Y�>fȬx4J��Z͎f�%݃$��ڿ%S�I�3"A��qI�X�1Ɇ�ؓ)�G[Ʉ�M��$	M܍n�oـ@��0:΁AN8Z��ʛ���Gbd�u�+�n+�;AB￳��o��,����r��y�g��  �h��<�K��N�*WEy߄�Sٙ猘�)$�J�Z$G=��)���Rg�W\���O���Xy�U<XH�`�&�hABmޑ>�I3�Kk\NOW^�y��cN��òfzIG[9�$K^�I��H	��v��l��6�OT9B��>��҉�3}5��ɝ��*�z�F���kl�����{��u>��`�H7p�DԈ�P?{���gg��D���h�	$�o�$JB��w���.:�L��7�}UR^H��@�@$�_t�f`O��&�(�\�&}��[���"�&�,����M݄���A���̟�^$$gL����p���Jr��K"�ye�3�kɤ��_Qf[���0C���j��5;.�c-�`��²�w.km�o]Ħ3d�v޽_��}��T��C�s���M�� �	$�n�I�%m�"�`M����.�h%7��d���8+�mfAI��j�_V<�	 �e��L{��2�+-�B[���� #bdL�"P���H
�7�?A�;vn�u��D$ ch��0vt�*	_eD�($���sĄ��H%���y�^jY섒E�:�($�7�L����1Iً�r���PJ:�n��fD3ti>��󤗒�݉�'�U������ �I"w��~�^oO�C��Ŧ�>C*���4S�M�:͙v�u�ϊ��C�ޥ珛{��m�=�P��ɀD�_�w�͇�0&�E0�w/�K�!ӓǿ< �����/>�"R�?��?��Ψ��x��	$�����@�c3	*�� $�A�$�I$���s�����?}����=z�n�ɬ]��f��-pl���x�b[�h�]��M4X/�p���V!��vx$�}��I�u��	 AosDy)Mi����;5�o�_�D�P$���IԨ4!�ؗNY$�^T��y��J�&���{�j�d����tI���@%���	S���Osf�A��Z`Ld��檖uc̀��̗�9��	$�N�1�"5-����@$�vK���(�%���ZK=��)���)2U�1�C��w�̳���"�$$�$��<�I�zF������ɼ��y��:�L��|���2.�fyK�3�I���GUF��M��%���!%�K;�RI6�H�%a>�/W����z���o����{=��G�����{=��l=���eg�y�N[OZɛ�"��{�S|/o�v!h�u�OasC�zW��Zѽ}�,w�>�yj���	�yn�J<�C�<���8ǵ��]�=ˎi�V67��'��Z�q4u�>���9Ȫ���,"XN�������ɞ���\��zc�\�<3_-w�iC�����o��)���[��o����{:+��{9wqx��ݳ�=�����&�#�F�$=�N绷�;$��0V�]7��{�A'.�>�us���N�����r[�3ٯ�w�ZY��"�׍�{�ϩ7���6�Sk�:�l�<�c����B`x�s�~�$o���4�S:])�y�꾡9!W�{��e������)��h������%��B\"5�=ιd#��O 
$�����iʨh����^+���J�d�ïl�O{�z��K��t�~�b���^$A�"��C�w��B�@�wcs
H���<Z|7���=�I��=!��4��(/�zAG	,^#B\�O���=�uC�V�3���Q#�z,�Ӕ�p���kԽ����-{�o�zwbMp��AL���U���S�,�[=�FQ�s������B��;�w����t�C�zl>n-)t&u�w]9d�:y��N(��(��wx���K`*��M�Ĝ��bs�°��x]GĒ�Y�O�J=�n�}R{b�a#��r�p�M��n��{�:Y�����T�"m����d��˙&�6&15L� ��$�u;���mOycrx��w$_���a�.�)"�!(�0b�ޣ���>~�%'�ߓ;6V�F1x�����b8��p5֋�|�xb.�hֈܓRh�rY�����J�2/����Ke�(�(�E��S-�m��UQ��Tf[��*�*�iGY`��±6�Q���\h�5�*��R9B�2�*TQjUAQX�A�#&5-PAO�`�(����ƥE�c���҈��0U�VcEPL��W4.\LLJ(�5��,DAxݥX�mM�`����e�LJ73e��V��1�9d�
8ܵ�,R,��יT]J��`�J�J�)mQ��8��[��0�9mX�U�Z1�Uk(֖��Y*���������b"��c�����X`�*1�b
)��ɍ�5�R����eֵ��]n��m���M[[Y��J�iJ�F��T�c���#l�Kj�#�FT�}J("�F��&�������V+�b)�ʖ6��֠�-�TX�����5�aA\��F
*�*�-� ,�s%L��)Q���UPUTDY���QGmQkU�uu��j���k�ͦ��no�znX<��~ ���ݛ�m��s�y�%��r�y̷����tԎ0,tM��3��:�y-'�\��e���Tڶ��WM)[b��mJ+���e��3����H�D&�Pt�Y,Qm�h�c��,0��"l�U�[Y"6��[h��
��b"7qM�!t+w0�uK�\,����|� jM�5�Ȥ�jݜ�Lݮ�WMkPT���4�����=nm�J�-X��b�x� ��m��3D�R%֎U�k`#��ma�#Tq����u쫝�f�V�Kt� U2�3Z�9r�&��4ګ�V\�Q5pM�8YW�fbؚQu����؋��"7n�5J�V[I��72��0��kٍsWd�̬�`L��ڭ����L���1���X�����C0�wl��+���e(h!P���@U�l)U�V��u��f�-�ZP+nA$�*�m��.��q���F��HbK��f��0��	`�d�[���k��Rn���u%�t`���u�sq�������RU���QKb馺�yw8HVٝ�0k(B�*�	�t��-	F��m)��J�:��R,����ZZ2�Ae[�fUslqV�7��� �B�[��RT(�.\�g�2�)ѕ%�뭭B�[��H�V:gW[h���[����s3ph�nH���Zc9���mz��caR�B�(��Y|�S\ü��d��5�YhCݫ
kj��Fr:�aJ[��%4��-J��i���5�Q���GK���1���V5�`��v�i�RiV� J�c��V㰦���h�jA�7M+Y��β���D�4\�7J�����ٍٗ\�:�fXJ�$�r��9���1�4�%��;Z�4�h�ae�[*�Q� L�i��&TiX:�7��EjS]�<�O;Ɓ�Л��SXUV]`.��,�F��x��rA�
��Ğ4�:j�h\���U^H ���t�c��:��Vb˩vTz�X�4ې��!v&��X��сˡa�5n�,MD��ZT0WlHX�!f��������nt���`6��2�3!����[���%�IjGB������8�4�[T��K�i3�$$�6��"j��Ў�q7-�+.V�+����mu�MP�f-ɴ���
�P�`��W�����#���&�Ur���V�l��u���n	���^���R`���i�Kq�1�ɕ�S����1-���5c��$�[�[���Piޟ	o%M3P�'bW����q�d%~f��k�HT���]ِr�;��&��)'���c<��ܵ�Ĥ�K� �9�<%x&��(�ӅM�ݎ�ix�$F�lvEӖ):/*B]:�a"[�"BR�$�F��53ٯPfI �w3�	����D�L����`���`�ޭo�1�f��Ѣ;�܉'kY��$�M�� �I}蓑0���������(�g=��Eg��3�ve'W�q �I���'���p�U�KGC�넗�N�@Iy$N��,~n�!%b�>��z�$�H4f��4��P��@�lļ�ԃEL�*@�Fj����Шr�����3ᜦg�d�MАI��bL��K���HJ�i����m׀��E �6^H�KG��N��t�L��'zn��$>�/*ͧL&�cF�C�=�,�1U=�Mz�Ĭ������ز߷�O���ŏ�^�S�̋Lm��m9o2ո��m��ea��2���h�
��?<<��m��"I@7۲$��2�{����$�X.zE�dAoflC8����t�̃���pI��'�IIs�lO�-�1%ni�-�8�y=M֒	/&��%��??J��o(3����"�*�K��k�1�9�a��?3��.��֦�K�%�}}���Ios,z����1�cI ��H���&+���̙�`�ve5̆H$�G;Y�i̵�a�!�fV�y$�&I&Cf>J��H��g(3�\�� H$
̃_���ቢ`����1f&�!V��X-h����Q���n��Y�1L坙i��V��*RD��t#!$�]��NF\͎�p���j4ϥ�l��ROCv�t��3<�%���$�C��h�J���($�G���)	$���B$��fn�GTfLm���7�nfS��|~z��HH~{���%�H��������@�wnB�gd�ȇ�˪:p=���m��[b`�Y,�U6��b��*�>,0��SkZccBL���b�$�XMXe���/��$o�t4�$�?}͞�Id&(�mfvb��j�$�o�{�"��ɚ�>�ϒIm���!�Iy�%�����͝�T㹌6��h�iK!Z˝�,����亹�B$��|���۸L�?nO^�$���Z|�I���@$�wG�m^���$��K|��M�
9��v����1�"b�U�f!���k�&�ۗ��GپJ��>����⬙��I#���f	;���O&2t&�w��l��$���*�i��"��
b��;2�)WCܩ�36C��1���ۺ�ˢ$:^	/$��ƈH��c�g�QA.mm�s����o+��!�udX�3=xQ ��X���33�>�$��ᱺ��z��m�3 &�Y�$���~���;ŝ�L���.��G%�r�L�I$�G4H �I����K�/c�����z	֩!�e�q�7�b�.i���' ��� �w�Rd�"0����I�r��J�%΃=�f8�KI���qF<޳V��{����/%��D$?l���,]v0(�J�_�JK�|�v�FK�AT�\��$K^���E �m�i	]��T�|�H�w ;�	Js֡+��ؼF�p�rb�.`�3(79��B4�S�n���vD��X��鶁��3dc�A$�:ކ���:�wwB�#�ҍ��E�l�n�!S�t6��1I?�<���ɐH,��,sW]WPA�>��`N6oL�N[)��A�2����!*����r�̦}�r[%1���4�^�\�Y����e�� �͛� �^��;e��9I��[��)��}�޼ֻD�H��ٟ	/��)零�;W�䁍�P��t_��3<,��2H?f�syq�'VCV?�>8ם�$���I���vc1�<�F�����F/�/�gnK�f�+������OS��4����]~{��D���*S����y�9���f��*�0/��.�.!�I�a�(uf����N�:�G����!0�h�	�6��)��kĭ����G[�LC:�T��H-n-[Z%p����V�#��Rҳ\�Z�B�HVYa�B�u��E��ab@�vt\�^�M۶�J�;Es�EeMh�et��6���pR-��X��̊T��G��t�jsN��5�����P끢ٴ�e���&���H�xlM��Rڰ��`i��@l����t����&�(bd�萱"�;(���{�O��~G&#��������	8��I �[{b�q��Ӱ���l{0{�Ȋ{���>��Zt�:�p� �N���զ%�_vi���kΉ��[�_�����M����p�&��.ɋ�3�ܑ$���A����]�p��k�Y���p�`)�g,��@�v�dz�s-��1��=m@��A��J�}&`$�"�%�c�H�F��.�.�L�(�E�	�UͰ���#&�ӀI"���|A-W�� ��Ϧo?g�{�|� ��ջ�l��is#���]��6�c�ړ(���k�VW:f���}?}{�P{%������>3��s�@���<k,�u���V�s� O�x�^�#�@o;�y�:	ӰgcTT�lH���a۵qS���？��`��2����8�or���SM>���Q���}��x�z��ѡ���[s�)��<6�暯]�X퉃b�q����:�c��٫� ��|0I��1I6	#�۶�"J�����Yp$��� �ƼŰ�o>h��#�	+y��'�G��Y�$�`�^���2Ѿ�'���<7�I�����,�����)]�FK�F$dtz�>�+FY�g,��P��U��>v�*���R�y$�<�@J����Oj�
���8L�)rXY�L�.˲7��6�U+�2����h�u��ƒ��΃L�`n��:rX�~��@ ���� �Wwt���vI�`Z/�������7�N� Βg�$'޹��X�cT�OU\�y���I���$�f32[����u���$Q����`��g�N��D��3�z|p���v�Z:u<i�=L�C+���%�԰���r�䲙R��h�q6.=�Q��3|�i����~s��\(focKcT��U:�> �χx����V��L��5�7���dK���n�Ƹ#;�c��7��Uv��ǻ��[QZ�p�B�v�$6IY��1d�A�kgrdKglz"�ꓯ�m/��x�u�� �Kos�v����h�]Lf�..Bf�[��aH��q]A�\��W�`��q��Ԏ�_^���E��r�1�8��y_^��I��^���8ަ`���_>��wt�zӲ��8�"4����^G�ǎ��L[�[�-҈!]�L�H�?:��+���lW*7^�H�r]���$T�S�(�pY�|�l�!�: ����8Q�%fg���[.6$H_�$���w`���+���q���lءӁ�Al��	�H��������t�y�dB�\DL(��2nZTR������j͘�����Kߓ���;��������_�,�o�nH���{�����<�>o�]��T\Kj>wLĸz�i����>-�6�[�ϛ�י�[]���>tG�sq�56u=4Ψ��$�����k�LMc)P�fh�\��ژ-���iZ��ىp�)�tޜ��i!٘� ��ә2I%�� ��E���V���B�V��S �|Ij�A�>P=�.��w)3�m�ǋ!p�@S����р�[�>%o?����5^��v�Rj����=.����&O"H`@�>+�� Y⊷�`�74M|H-]�!�B���������;�Qg��t�)=R�����DFg@O��k A>'�ݽ1��1�An�xo;�;�;;Y�cT
�n�H����f��ctDhk�z���A#�w�	�{.����e��%�V���P������������O����ߗ����?��2�;'��n�>z7�,�o,��ţ==��]��ɕ �A��T�]���/�^��\٬ɴYct��b$���*�2ĺk�35�PX�8�34
q�^�˜R���-[)��Ų�Kj��0�	��ݔ�`u	J��!�yڠ�If��ƺ��"���,��8%�:1���bf�B4G�Q����0 ޥ�U�U�Ln5bE3�6m�vG��T]aw�4(���.��2Y�E��6�K��k�������@�F�f�QlcN�\���a�u����>�H���k�x'�^c�>�����m�]�ַov��xq���#<�~��!٘� �>�ɐH !;�O�U�|o�Sg����y")�:gă�w3��,W�Gy��t�ӺI��m��	�u�I�8׼�L�~�U���|��D���e�p�ݜ32x�?R�1<](��*���Ǟ�>�7&|I �w3M�t��s���@�w�''���	���曽� �ݹ�x�R)<8�A+�zd	���,�6wr25�P���"Z9��P��5��uJ��C	�@���ŕ�5/��>��ݰ���K���� /f�H�|���:�g0ܪl��c�=�@�Ky ���$˃:Y`%�v4�n��|��?�����cUԽ�=4����w40Ɋ�q�"ճ�Y��BVoX��r�����!T�E��<&1���}� >y��"�W����|@$�_tz�O�l��G5X�H�V�dY?�y�ɾ�$����|��XpU^�ا�YF��)��'�=݂��-�d��$��z繞��/����"A>k}���y�4�SFdS��uE?^̒��i�p���&d�$���I+�;7\憎�� M�L�$�� ��D����M������Y�D��	d���gmGB2].� ��8�����l�ؚ�K�HhƓ&W��d��'pS�zʎ$�g@���-ށ&޹�����ܻ[�U@�B���n���r�'%�̕�o���7W�%򺧢H$�� �WoG��baj09O\�%��)`%�v4�l��A$���}�Z��5�wvq��������==3���{=��7����LB�R��e�f�z��9|��������a�{�񗟨�X���m�������U{�l z�d����(3xag��Ǟ�6�SN���t=��2X�j�%�<���C��%W���3��|�hi��Ύ���9r؊j��ુ^"�$�2�­�M�w�������w�K�zHJL�w��r`�@�>�プ4����L�'l���^=���.�C����+ �S��;��:����Y�bS9����۾\�~7�7|#�R�˝Гr`�K;����J�=��#�k�f ��k�慶�6Ҷ������RV�N��^/\��d�Z�}u�{�]�2�)"��i��9�xd�z�u��e�a�n̛�0���(ޯG&�M/�揌,谷c� G�3*���l�"�� �zi�I+��
�+O��<����7��^:7�W��������~Ӌ�-Z���'Z��.7�𹴌T�M�����sت�DeR���##!����S��c���*�f�-���׮u�-"�!v���Ne�c�Rq�_���U�єp��⽫I������=���<)��!{��v�r��;�gCw��5z�3�Χ��нEh��\e��~:��?p�s��j��%�9��}���Y�r���=���r�͐�ǯ���(�
��	T�i�xca"�8��q��e��&�,����D����^Z�v�3٪@i�3�l�e�G��M���}rC����1��4���{��hr�/�� #�������۰�Y�8�W�f���������n�'��sc�N��`��A� �>"�%#�U��)kJ���*���d_�UV,����(�h���UQQ&Z��U��Ak
k(���k�6�ugM��e���6�Z�Eʅ���H��F��T�\qR[(1���4�AT����-Ab��0�F&��\��-
?���iZ��-PX�(��:�T�m��kmk-��m[]j�f��]:km�����].����ֶي�j�e%1�X�1��E�FE
ƶ��ī�ESm��ٳk[W[�kkf͙��""�J��[�DƵ(��c-1
ֱU�J�EX�^\�b,�-�VV��$�kUDC�.������Ա`���DD�aV0�V�sf�[6�gZ�ul�m�6:몶mu��m�oZ��m�-�m�������3l�`�ZJZ*���VA"VE*T�Q�m�
�!h��Ԫ�Ɗ���ϓ� s��|�?�#���8H]�@�Vɶ;�LY�p���=ts�0�U�f���s��vc� ��]��K�%��.�
�n �ȵ���9r�3&������Z��$�=��>�d\S]�@$+� �{�d��d�g$,,��}ou��`!X[-h��cB�ۜ�c0VձRP&P�&������}�2��gd����e�O��q��|Hn��n,�Y(�u@�IY�<KȾ��;��w<�7u̐�䨻jn����!ed�@ݕ�TO���[�p�O�����9�~���NK��{��x���� �/��kq���J�=W�����	�:��2O�\���9����T4��6l��W����8�|I4��"A ��?��4h �����z�"�L�-�fL�Ow��yom�{SG�y/N�Sp���e2�᳎(;������&³�C�!ʻ�Y`\���<��}��%��&�Q���z����>+>��^q���4#�U� ���ɐ|��9L���_�~���:�`!��ňaX���;n�z�B݃9�G��-ݕ@��]sM_����$�q3R�qăo��>Ԁ$�?<h13��C�@��E_M��Pt��8gd�$���q�o�!�պ�	��^�	��� ��x�oUR��UX,��9E$������΋�A~Έ�����}۾�H&޷&|H$��D�w�DX`Θ�`]�P+�^G?���3d���$��{	 �A��CE���y�V��Wt�rb�B��3����J�ǂ�{��|��v���c�����H>%��<� h�wp�8&q�ɦf!�+&���C0I��eLq|QW�2�э-t�]�dSnk	S$�x����@�#ȧ!��3+�[>���J,�BX���|��x�e�+1�p�L��ԋx7bş�X�_��2�ipQ��$-��Ml��s��(�s/*�5���%�MH]ne��M�LH�+h� �/�Vf�Z������h��w*Y�KU��Pn���BQ6n�e�\��j2���
�5��ś3%�ˠ��S�eW�;h�wc2��,΍&3
��i���%�Tw7�Vd�R�YA^�qTt�Y���sv��lgbdaF�m�]�E�*�n�����5�'H30g�U�\�7w�$��cɢa�񥓍w�H!�!�	�:f.]�% I��xW��c�x�u����$��>�D H+�\@-��UVb(i�!s�x�vu�L��;��&�������|H=�g)�.6Y�{P�؏@ ��XH3y��Iݏ��)�᧲b�b�wXH1;PмIl�p#Z��}�qMOD�����vI�c Hukǉ �n͉=WW��%���H��>�$�{$���� ��V��h��ߑ���)�!YI^6��D�wgf���7T\f��X�,]K3n��=��>�M��>}�t�A!^6 �q�zkԧg�ܻ�����/�P B�{0Hh�-����8p^g���A$��Ǔb�����_��$Q91��M��|�  ��y���E���Z��-�5��8fw���{{�y�`�ffp�C��x}9y��H���͟}2	
�Oٯ���ٱ0�M��`�ݒP$[�^"	-��A�b	�gOkM�eNh�WkY�O��d�>j�H:g`��=
����޷��0��z}���7�/�I.����!�{���L�A&7�6��tȩ����pv���/�rȤ������11�2Ly"�:L���MZ���Q��#ą�輪 �#�" �ΆY���,Y�$��~����m�=�ꚉ�,AnjF����]�E��fͩU������d��v7�-��|s����c{�O>����� �z��3�Is��.|��:2G=���c���x��aA E�vȒc�.������F4�#�gc��O���'NHf`����2I>1���G�Ŕ�C�,P����8�ԏ,e�Ș�W9���g��q�p}��mY9�=�܅�)��(�"��c>�Q^`�(��1Pv��ooӫ�H$v?t�H��}�k�5���&]�%��z"���" ո���[Q�$L_t%kv�|���w�'��I������:��У����I+��ά����[N��	z���!��	��A��ͨeJ�R((e̓Ƙ�n�!�iY3va��@�:�Y��vZ�nS�42L��S>�g2I�܇t���^�d�I�͏@ �B��P���oE�e=�u���I>1������F�S���c����8)x�i�0�5�5�]��ѻ� Lqt�k�Ss,q5j��d3�$գĻ�Ħ�x�|O��2X��\�}V��z
��3�Lv�@>�n���58�tC3p���̩�'��u_a� A��mx����ѠG��L\�۝��>�w7��N���xB���=�����^��m8�F,��e�z/&��Ɂ�-R�b*��\5�����}�|i��y�p�:L�t�[*�`�t�}�4`����c�o�!Z�*�ꃞAv�t�~�����	�;33�ə�v�\�^tݘ�"K2�-��-��ٖ�cm�nWˮM����]�?7q�$��_(� ���� �׹jK7/x� ��*l��'|�đ������ 4N��
�N��՗�$�j�g�"	n��A�L];A�̺��~��`�:(8v2���A[��>^AxL�\�UKũw-�Hm���f	�M�K��f.�ρ]=��snY��Q�4@+�\$,���G?P�NF�$��t('+�md�wD2b�䗪}92	$�؈�U9�0���	�Q�|HW��>$�����y�v��fv�̝��((�x-J����5y��S���j����(�%�i�ɨ.�L�n���C8����J��7v��-8׺��k���`���B�?Z>y��-��meeY�FX�s�W�$\J���6Y���4sD�qsk���z)5�V��`5�ڒ�1�]1pmA�Mf�64�R\�J�T����-�,[���3����,M���J�a���.c)s
n�50�u0��
�$st[l�D�����4�Y��FiL5V��HŲ�T��H&�m���J�B]����Υ�j�Li���bn�*�u���"GU�\��m+k3p7$��������0`�:Lӳ%��Y_ �u�$��� (�,��3��6K�?��2�@�D_bi`]�r���H� ���W�|�n�,�$G�i��I�~��y�9˧�zPO��&.�ْwwA��3=�]U� �K�t� H+聜�wK��=�Z�<ImnD�I>/����	���tPp�b��n�X�G) [�z� �O��눔�w?�R�t�	3}3�0MK69%�t���WODB�l��f�|��G#�W�<T�tI��	]��GOkiI��w�R�eZ�~�CG؆).֓V(Ep5vfnL:$�̶��:hǊ����߇�-&���﷾ɐ	!�#<Q�>�ɟ�V����͍΁^$�g<z|�(p�&�ز�7��@�>K���[���.5��TA��\�M�f�7e����g=���_����~4����5Oڽ�l����Fjvo�;�y�R�����w���2���}�	'ĵoD[���݇����{�|�ѻ����3�r�B���L��@��t-����k�2{<A�rH[��	�N�$��˳�fyB鮔#Wn>C:�p	�fy���	n� ���;շ]��g����S���c ƶ�`���A�rװ�Y�LOtA ����Y��>;q��Y!���+��0E��r�LF�tl�Z�X�%-����5�,�e]�	�f�$�N���{�*��1���=�n��^ȹa"��Z���e��_L'�&n��N�LY��c�&A����7��B	$�:�`�^^G_;�A'<���_&"�z�A�y�XѠ:LӢʏ�+�k1�AƬ�A$�{"�&�qm�y=Ň���h�s��6�2Ե��j�d�k�%w���?���ݩw��X���Bق��3�ܴ]f���-:B�?��Y>%^�j��3��v�)܇g.��D�z�|ܞꗶMD���>1t� #�O��m��>$�o���p��'�(��k}��.~d�K�IM������>���f��¢:�>��:������/�[�Pnnq\3D$�Л�*���M��h�b�je۬�52��)���"Xi�'N>�a�S���c�Ƶ���;`O� �G�w��}�̯5���$]�s�$�69rIwd��d��Z{�c���P�D�B���&}�J:D7�u���uN�<�\n����'tC�,�y�S�d�I%�: ���؝9�dPc[A�$Y��g������ŝ8L`OCTn^�<��g�W�gp�.�� 	�!� 	n��>�O���-Uo�P�Q�{�*�������{�d��~�z�ߔ�{�]�g�09�ۤ�2�t�4�fT�[�ݩ1q+�*edH>�Ȗl!��/�}�2H }}�ʃ�A;�b�^Ɵ��cty!2�0�0�nHܮ��x�b�"%���}�1lۍ%ur}�!��3�NS�b�="��Қ���*��ָ	Ge���2�L���=���$Y�33�[Ul� ���%w>�'��sע�;�T�'ė���z:䃬J)�Iñ��S����f[���U��f��h���/(��	[�dAi�f��O����xX�'�c���vL��g�t�$���`�g�ʤ��KD�^����A�v J�}0	x��I��;��g�ʶ�*5�rx��7����E���F?�̽/ �/z7�6���h�������� �ɓ�	�I˖���ױ �l�u�$\���"�<A��`�|�߿~<����q����ǧ���q�����ݞ�g����z=��tL3F���J�c��h�,��Hy�
�����T��>^��Μ^	�c�o����+�{s���k{�Kn�<<4��Z�����4��υ�;�}q]>����m-�\T��p����<fSˡ�ǆI����[��Z��ve��7���	�W�����e?.9�u>"<�p�&�#G=6.�Wg�]=B��\c������}�����Y�Qq��Z#W74���X �qn�y�<E��۾��o��M,Gk�%�B�t�X�3�bF�{��:Fl�q�S��=�t"��*�� ���PR�Q��q�o�kf�OY��|;i�twy���Xi�p�mZH㾪�y��b��c��.�U9�Mr�i�α�\]�v���'��nx���~?�(f����Z�i��w�'�<@�'�>��*��;�R�m��j,�ݍz�n�=��Jq�1h.���y�a�V�aR�.W/uo��v���`�%|�%�q,�e%h����!�m����r���k�jm�H�ؗ0�m����C���"��|��pǚz��pL�}�n���*�$��MF�d���yؙ��9դW�wx���XW�k���}ǰbf=��߷��Ecq���u|1<Bp��S�����w�/e=}vqL7�VY�{�����71�2w.ᘽ�evu���]�=w9hd9��h��y����P�c[gOj��W;���\� 8	�$n�� �#YӾ�젬{��
Eea1��3�3��t��Ö���,V5:�mw����vW;o3c���UAAQ"�,EV"���ֱ��i�d*[kJ��U�j̴Q�
�D�,�DU���1A�TJ,UG�Q�*9kX[j6����+kkQ�5��U������l��kk6�Z�ٶ�+KN�2�����+UVT��("�E媪EP��b�EX#�ՅUclR���M���k���gmu�,�YƂ���������1Aa���h� �*�X�!Am
'YUS����ҥUF�r�KiFԕ5�ٵw�u��iu�Z�c�5��E���ъJ�aYX�Q�Z�2Ո��bVLE�YA_)���E6�%E"���o01�X��1!c���u�M�����l��gVv�;uu�뮬6�[]Zl�ֲ�dYU�"
bVAD@P"�(�O-=�,������X�����k�9�V��/���RdS0�v����y�\Y4Y�(�5H5晰[-&�)������YC��ש���,Km��lM��Wlɥ��31+k�V�+Ify��&��	$#f̕V�A@��A�0��]�]�mZ	n��&�aچb
��1nu\Y�)�6%��{u�[SV�K�Y�V(�H�i��(E�x��4u3�Z6[^`�WPL˱��-r�`�����Ba�k����J��e�Ε��u�.���	��RieN���x[uPK"�w�m�[���v`���[_���^����ckyLUk��K������ٮr�&]c�VS<�͕l�5��j�dj��+Z	.)M�Cb�v"�Š�ͱ�I����b\ͱ���+�,;Wm�l.h�f�5����=K�c:�!�5��e�Fպ �I,n,�Z&�&��+
�ʡ�d�j◚�%[���e fҷ��5�v���+�Z������رL���)B���8��"���Ƣ�,�7vY�)�E�pҗKq�V�Rb�CY�	H�FW��D�bUҘm]mD�-J²^�x�ڽ��Fdkm�6۫g��m�F�\��v#Hܙ�D�
Sx�o1�X�U\\Ch����m�6l���J��,"6��e�[F�"F;eүl%V�����҉P�4a���`���mI��&��܄�Qr$Su���6ݡa4���5����&S`F��ڛJu�a��ْ�6�b�LG0.��d�����Qoe�ѱ���!q�#�����>WY|c6���]n-��9�.Hf�ˣN��Hf���9��B����S�+�-�c�����\�+Z�H!r.��������Hs5�!�)a(�b5RۙY*l�k���Hfu�v��&t�Цط.��NJ㶍3]k�y�+4xv��ʛm+r�&��W+�Ut�	{ku�魵���)4))��\&	Bf-�3H�H�P��1��\U��cF]6a��S�����b�]y. Efr16���M��xk�mلP��Mh��̯X����A�t��n��5�L��qkeYn���9�V\�Ψ�� MCi�1`A�4��q��]�iRQ�x���xo'�n..d4P�\WuE�=�L8٤��!���T�V��K�B���!�ňY��f��]c[)0�G�6.�~�������߽mt��mͰ�$��{�u	�GCwn0N䳗g	:w	3ą�W"A�4��,��O맋qd�j~0$���>L���k�~�!栃�J)�Iñ�o������H>3sCCM�׮�H��� ��t�1�ruM���3��t�ڈ�����x �	�+���J�����ϼ0�W	��d�"�?�gpXԩ݌$������[{k���}`+k�'�a(��˩��m�t�\��J8�r�E�����N�m���6:�KXs�T��V�k�7g7�sߨ|��k�p=�o�
�܉�	]� Aj,�-�6Tˈ�W�O�{X�w�3��w� ~��#��T���ݘ�SMP��EK�]D˟���9S��e�ۗqḻ�*^�&���)y�e�"�t�f�-T��=�!��gk� ��>�H$����7��:Ԍ�p�{�o��i�ݝ;�w	�ӂP~��O�]{�l����C%����3^H	m�>~� ��
p�fA��x��k.�"n��F�LI^I��}"|Sw8f��n�J�*E��$��d�,O(���]�fv+�%�y׌x����{�+*���3�@!wv�e�Q ��� ����m`������l��i���,�3�i5�l�a4���E�6[���;p�_~�}�Jכ.Yl������� ��� �I[��gL"�b�<o{�t�d�$��z ��'A�9ffA�3&���e�9� �I .݈�oG���#�dK�f��~g�S�øg	��3�����H*���/ /��u�i�[���L�p��f:��'��J�BN�o����C���/�[}k�<u���@Y�2Dn�v�%� ��l��1m�7��%Fp�O��؀A[��	���K
Z��ғy�����_�l=s��x���	vt��'j�u�-�
�������PF&%�b�fJ��_���Ή�uv�'�>'�O �T�G���� �=�v��S� F�N�3��M�7U2�a��K]�.l(�iF��L���8�qo/�NK3���]7@!e���ݽ�%czդ��Q5�N#��u���]v��?���!@V7^L��ĵ�El�lu�����Up#ė���R�c�Ch}��ʂ�/��9L̃�.fA��x ��� ��{ҹ��+�S��}�M��$�i��@�d�r���gg�B�m��q�lp���	���x �	n�ɒ�����y�9�F�\��6�q�t���j\�I�O�Y�w���d:B��G-��궖=/'�c� �4=�m�8*
L��<[ٻ�uUH�eS�Mɑ�}����a�@]K3�gd�ܦw�Gu̒H+���#9�?2w���{ A�}�2x��otBb�*:1l)Ρ$Rߪ��_'��Y�WM[=y�m�\�Э�5�%[Q�.eͩU����n
	�����l�-Y�>H�����{��r5!x&��� ��ΑQa���fv0G>�~�"��YUM2<�$���ݳ �|Ww@�L��ٔ�x�X���$ M*��	!gl��+���K`~�0I!�/$�Q$��~���5�&D;�B��[U�R�)�#�� �����7���&Wk�f5����Ȯn;"��<d/l�Y.Μ3�
�n#��t�����=;���#o}S �
��J��P@�O�^�0m>���?Í����E�{�ݼ��B<��l�=M��)�/{�f����OZ�(�#�����7�ݗ�ݫ��ԭP^Y�)j>K�l��^�w��O"۱�����F��w^������˖�s�F�0�ĸ��7h�e4pV Y��� 𘣥�Y��*�K��7f���khb�f�je-
0n46�t�6�;L��Is"*1+&�tA��1��2���leu�YbVY��S�@᭸�m�5bL�A��pyn�ٵ6�Θ�P��B�Z]���3u��V2�lGJj�ưD(�T��a�J0�	Θ�3
6Y[;W9��v5�el��stn}{����$���Q�r$
�؂O����Q�p�Y��7D��
g.gĒU�@���-�$K�)��ĕyA�KM>�w����O����><|H�1m� �Iz�FZ���	����vD;�)���Y��A\� 1$sNeZ��z�0A ��� ��[�<	�A.�NS;���S�f�/���D����+�y��� |���y������$���s<9�&D;�BEb����o�� g�Ŀ]3Z��� D�D
�@�57B�[���
����=�Il���K�:�����[��"K�3&�SB�ˮie�h����~����+D3Y����]�k�<�	����j��++y֠v���$�Kv��m�v`᝝�2gyu��`�7�
�ؖ>ϛ\A]x��u{���7������ƯYy:/C6T4�WUڲ3n�Ųϴ�P�ό�"�-����yvMV��86mڙ��2��r5K�J��x)baۓ]���T>�D�xlߺ饟#��2�`�.��g!:ζ ����$�Ԙ��{�e�sh9#A��׳�>%���e�.��;oHM�̰�}Oy�ę�� �.x�]� �A~�a:6��I��{Q�[��.�N�;��V7e��3�|�	~莆Q�z�N޷&��T|g�z�{��+;.y^�g�zy�K���؇�l�3yЗ+�C<옸U��1�b:�6�GX���NRb]"���/JA�L�wt��Q�|
�
��b@$�C�t#1�DӨ��H ��t�"}�{@��,S0vgj�7V@��EB7/Rӷ��z؂I��ِH$�wG�w@S;�3k���˔Ⴢ��2gy~�ؿ'���>� ����Gq���._P���g��e�f�R2�ݲ*��{���*�kkS��h��l\O!g��=�d�����g5�X&��P2팟}��B}�l���}�<�!��"�fNBu��44B"���͙�� 7���oD@ ��֩�2g�����MA�"�4��vN��,��A��Aܳ!��n�d>R��F���ٙ� ��<|���̣Ec�{��=^S��tͪ壥�pr�qY��L$u����n�A��E�F^*�{����wVܴ���l��@$Fv<V�� ��|�u\*��Ȇ깒A&/:wp�]$ȇwH̃\�����u4����j懻�$IW� �-� ������O2��~<M�d���2d��}m�b	%Z�1�5�Q��l��h��A���b�>�z"�
I)I�����菧Q��W��#]�"ܷ�Oc�@��GY�]=)�����lv�����w�J��Cl�[���囜wQ�_]b�
�B��A@阥$$r�0'��h<�zd��)�<
'A��>�B�Kȋih�d�nf���l��{�ԟ�>{y��af	��8i�r��c�|~�݉<��]�(��言O�Sv�@��2j&e�;��UO�����"�b1�YJwb��%q��#m���Q�!-ڨ�eW�z�_�Փ��3��\t$��2|@9��3��m��]^��.W�x�QNBt�ܔ#����<�m��PI�-z�zF2�#��=v(rf��n�����k�]��wH���(����� �1o)��U�q�IX��lމ�>������fv��Ge��kE�����ַ�1�^H�Wlω'���\)�k�~`��~$C4R�~�vt�L�ӳ;ą�"I/��"�D�w/!�{%���	�k�$��;fH%��= G��V2T��uu�h������n��s!hVl��u�l�l��M��;�����7���e��̯J����t��ݓ���ܣ��藼��7S��ON�<;:�|&o�&.�%H	5Pe��T���%�R�J���[U�bj�a�ݫ]L�]R�*U&��e��fa�&b� �m�K4۝�t�6%��pY��!�-���d�Ê�Ff����V��c���
;@6j��(�;5�%�n�ō�]--  )�1K��mЋ5e6jR.��j�&��av�R���+*�Ì4a+Q���
�ك�(�.% ҫ���le�!,�,ᆡ��k�kXY��[f���1�e\CGy�߲{X���ٓ���g[|��w"H$��w�A�����ՕM2w'Ur�I>S[�>2&��t���L�ĕ�� ��lOS��UJ�V	+{v$>;� ��s���7l'	kj�|�+�����;�(Mw=Fx�s�Wdz	��UԤ�U�d�$c���7��.�`K��f|@�Q{�}��jy��m�H�͉ �LU�@ ��ܻ5�Z�9�N.IM=s~�zI'kj�wtAf!ٝ�X8�q��w@�,�,j�Nwl� �z�	\��x㹰�����!��{���eͬ���lQu��&��٢[�AW\�l2�L�����.&�Z��VG�x���I>\��^g�PӯpC[ީ�1�U�|�������8i	����%~>�_�]�a1ge9YnX��6�9�냸��<l�N���
�MI)�J��

�ҙM0��"	�H3Nu�F�VQ��w}� 2���ޥ�15i�ݮ��ڨ�H$���#ĂB��� �yfk���}LI�4*��t���L��-��O��x��_�L��%�o	 ���<|�����e�I��Bd[o\�����؃g���+!z$�ƽP�k���n���:IǞz�A�9�N�`K��h]��bIi���FK��k;{��_���lA%r�PO�{�2^�)nb��V�dc0�2w)�a�
�e��l��\�5�9u@�t��Y�
=��w��~�S�ٝ�p9�q IV��$����5�v�:�E����!57b�E�d�;�bY�ӳ����~A�/p��M};�HZ��@$ ם�>$����#T��]��0>vd�U�Wl�>'Ƿ9�ߏ-��vq��������ێ8��������{=��?���T���e�p�CLUz�F�餝���L��#���>
�G�wOHw��S�{��_s~��!A�>����N�7��fζa��q{p2%���o�I{��8-/�g�~����}�ӟ^�_�a�}���a�)x ��Ex���zy�3�C٣��N�nf�`HP���-�nI�%X�rg~�Ǽ��;73S������6w,��GqR��!�{���\��8��_e�g��_>�2+�����<=ஏSۛ�����do�L�r&/F�i�͉�7yJ����~ɛ
	��9Ǿ/���px{/t�Q���{����������؄�Iʞ��h���֮��<�������|��Q�:�Tg.��x<�]���W��U�9ج5u��U�_�X=)�\�&C�lV��i�@��{���������t���l�}W�S�D^��_w����=���bu���{�{�"(I���@6y���i���;��y��N ���yO"�i�::7T��ʝ�x=���^#p��2Z��k�t��jpS޷�i|�� h=�&yk��t�-]�Y�����¦�ֽ����dt�����728}w'�E���ȭ����pg���L�6uܧP=�%����C�6��c�jΣ=��-:x��<���g����cC�����}�qz+&o��+<,W�I��|s��j����)�}8���c4����'l��h{|`p)2Oo��^2�`���$0�̠dK^0�l8q1�Lڍ���><@����go\�����ef;"֢�$$ν� sS�33<D{[[VյmmlկY����kjX�P��+����FLIQU�m�`��+�`,̥AH��gX�H��\k�pH���LHX�j�mav�,���$7J��˕�J�31TL��(��-
�mT�ʐ̱a�RQZ�VT*Z6�U�Z��1s0S��J�k
�aP�h"��̭RT�%���h�\��1�JŬ
ʂ�;���j(
���*��q֢����\�`��G��A�%e�,*TU[KE���`��̅`�X,����B�K
�V5�I�+E�`���0*T��PP�u!�7�Q�X��IR��c>�m*B���,X)
��6�-g̳Y
��k>̖�7�����L���x����$���"h�[��1.�3�v
~�A�-��9�[1� �wz|���w�|V�g�s7Z�	��QA�t�ܔ&�mF~܁�m��uǳAjO
	$5��ψ ���v�^�:��̏ٚ�fu�Q���քz�k\M5t�ܮ��(��;��9�N�`K��{�=j� c⼀M��	${b ;C���.;��Y���=�t�WV�.Έ)Ögyt\�w.��y�"�90��C^^��ߗ��Yj].'���Eld95���^K��d�;�vv��ʮ�%��_l>$k�-+�!��r�I�]�L�A%������	̜4ɇ[�v��=��y�ې$	ّ �5�y~�������)ȕ�8d���?O{����3�#�j�%C��s�pNeY/����݊B�Q���\Pەy,���0G�p��T��D����0w,��Ao���A��d�.��fX<���_L��|Wtz=̷��p+h#��]U��L�,���I��USUeaU�Q15�2�eS8e�jJ���1��%WO���
X��P������2J�@�n8�H�m����#D\��S>$�b��A��tS�#1�]i�yף˳�cc[7rM9׶~�$c�^	�m~#ё5us�]%4�G
�_V�.ΈIÔ��(��Ǡ�A��� �
���JYGh�W���e�z'�_��m�ww�wvggi�=]-9�$��`��\z$��fk��z�.��q�@'ź:x���'X;0$;2p�^0��͹�\j6����`��}$M{ @k��#��u�8�)�j
�i{6$�y�OMLh5�q��≻1t�|ﳱ��c�}�<'r�/�c�?�-��%]������f�؀Df�;��A�:w�[M�-����0�A��
�Q��5ٔ�fyZ�t KIR�uЙ6k�^�sS�Hh���ב�T�[7S([^mU,��bh�eU[��Y�*��u�A�Y��.�3�\3=U��J��lcg6�M�H�@�[.-Ń�#
�h�κ��`v��լb��X�bU�&ʔi��777\4a!kMc�tQ�au�2�-��_
y�a�֒�������K��V]��D��NFmM�l�w����V�4c��?��}y<��f<x�H%���AW4pv`F��7]n|Dc^G�D�(��:N�Jz�Q�����M�,�i��=�D�t�Z�zgĘ�ں��uP�i��g��$ȇw(L��r�H�=�&�z���Ft��X$k����$ǳk(�gD$��gzk���y��x�8���A �꽙ѽ��Y���\� �5�͗wpX�wfvv���WL�@'�o�Q ��v�f�:���#�N>^L��L�k���a[�^$���|�!�&`�5Џ8ێ[0 �=��a������.���ʓ���}��DC�N���O��7bGy Aݱ�y��O�]� �;�4�
s�E;���fw3>�&��@�7�U
k�yu���m��Z�ݽd������/gn�ٮ�\X[��s�{�����;ܧ�W߲qڱw\��jG���:� rZ�[�x{깗�M}�� ���t@ ��B�xxQA�r�ܔ&u��d�D�����:�C�3�����|L�2y�F��w�[�9�x� ՍE:L�w(U��}=ãp���&��)���>;N��I�݈��܁�����GDEL�ۍ��	عL�A΋�@ ��x}�ބ�07�W>TH$��؀I[�	�\�:s�sX%��rc�+��Y�2=Me�X#�U˥mu�0����s�׿~����ٝ��v5VH�^�\A#��� �R�1�T�j�I�[��q:Y:LC�Nό>��sG*���������	� ���	�W@�}Y�-��nw5ӌ��$@|6�S�8vg3�����y��^H/���7tOTr)�O7=§aҸ�уyF�䄝�����s;־<�~�y�~վ�ܤ��t���X�����=5JG&��<<^*��I�nߢ��>� "m�Pt�;�����jh�QX&��<#<P'�	ѽ1��:�%���14r)�3ܡ]ˈ$�E�I�3�8�8�����U��s�$��'j��+���@��ڒŮ6bk����R�R�fTLє�#���
,�[p��ׯ�ϒ�;2r��Gx���-�^<I$�F��$���([�Qa�6DW�'�� {�?	�-����[�n�?����{���d�y�R ��D�t� �#��I��4Uh��k2;oa�F83��:t�@v�{�'��oݱ$�M?Cv}i��x{���\��I�wL��H�<�ӹ0vgT?kz̆}�ܢ|z�^<O������ݯ�����,CS�G��r�'B������sp���0��r>���I/?l�d&Bix�	+�Ŕk+.b.kV#�.	r�-�EKM�(���|�>�	�w$t�9p����	��#�V)I��w&��Q�'��}2H!ol������������o�C�/l ��m2�!��u3B�l��,�T��gh�c��tL����ϴ��jء��ˈ�$
|܉����e��q��>H^h��O��tgD;3�L�"Lz�nD��U�ʬlh�������>���� ���7����/-���_�g�� �t���hiۑ$������1!�F����2I ��A�3��G9t��E��\�
q�,�\�fAf]tzJ�ǉ�D�~��T)u���a9��@�Ι�!�,aI܄;3��,���y�뢄1�fb�u����H����u�`@ _�X�=/�7�V<�i�4>D[�o2�;d�Y�O�Yw���'x�L"��^�>��םI#ץ����B"�O{ً|7�����Z���F��� v�+k6!��B0�{M��kf���^q.0�]˂�y� �@�3j�82�J6���Q!�]"8��V�Zk�8�Y]�dj�6�g�Hh�b`����jӱ�).�Z�W��It؍jmG7a�����������qM.�D�e�[,����q��J�w]���ff	�]������(�5v�����=m�-�BkX4ŚdV\mrY��c�W7��=�nq�^.��O�F�\������;�q�O��l{����c0��k4e<�s��g�M��S�`X��B��E�x�=����(/`+��v��B ��vn��>0��O:l2J����@~���]�"���gz�}�!c�< I&�S�Y16�W`��n쑾�s���w�g\��L���W5��}�؈�1i�i���M��Ăs�w�Ǐ�u��H�=*�F����-�}]0SX�F��X�E��Z7^	$k��=}�ZzD�M�� ��7� ח��wD���o59/�� �L��X�Hj��@��Q�[��s�u�Ռ��5�4xbfU{������$f��}�!___ Yx�	����3�E��X���������!ӰL���[uӤ�����=���qdy�8{2v�&��fFZ�U�bQחR![�����	O7�0_f�w�4~@w�~�&r{ݯ���b7[,�}`^\ �m3QVا��}[]�	U�	'��}�$F�Sk!
����+�I�`K;��ڇ�@:��H%���k&�n����W@�G����M�^���t��K;ȓ]��9ܙ����Zz����$�T�l�$J���s:�Od��^��G��@ ��rΙݝ]�i���}ϓ�*y���	��O����2I �&����Hw��⸺`L3V�Z]�86Ic+p��Ɓ��FY�3c*�f��H�������b4X}��k�$��lO���Cwt/ܝm�%K{�x/�D�_<x�Kf�I��M� A�wx)��E��Z�ݮ� �ow�$V�?�Wm��tVU����6�v�ļI40���&r�	�y[>�Wn@�O���Ze�ul0p��6CY��l�0��\��k)甸z�������kF�	�X��ԒXC��S: ��ȳ�nIȓO�k�z[�� ��}�P$ǒo�Ȉ�u�$�0%��B$������R��ޖ�L�MD�I[��H$-l�r �)����eк�|H��	;�靜�w�F�. �g@b�(��M�/v�w��O����E�v�2"(0|���~�,�n�p	���Vl���\ܔ�[�h��,��jԄ��Y�;�X��!�Y���:�ӷ2x�ם$g��s\()3Ի��!�\�eԒ	*�"�y�vE�t\8��P���|Oܖ�}u�H!]�A>&���NW<a� �m�dn�Nz\��6���æw5EEtA�%�ܯ!�� �ou�����$��@�|HZݪ���������L���̿�r��� ��� ���� A����/o�7�;��Ӈ���!91)-G��+�b_p�����i�t��Q���T�3jY�o�P����� >�׌�H�܍9�t%�Z�����D��A�zg�s$]3Y�$*�ڋ�y�܉;l�#:D)�O���$�j� �ͽ�>'�sj�wbTy1�����m�B�g4�,���&R�Pf�o:�]��'w(�;���;�2-���vǘ���:��3�T�7Ί:�k45�D�|��x7����3�t�'TuE��gw9�Y��g�<I�65�A>��wL�M>1ꈷ�M�n�pc���N��\8qT
�����؟	/Ξ�־��aw������I��2L15����ܒ��fJ��%���ׄ��u|I s]��J��s^F������J<Oz'A�����'N�}7^+��:��_�f��e�Z�}K��A �WvD7�7�������ێ=��8�zzt�������z=�חw7hd=�W
�Ś{�"��Yr��\ݔY�= ^z���}�����o�20j�a�,���4t#�a\��r��!��/�r�ro��n��qk�6��(�顉�ٰ��1�q�)"e�$&�["�2���9[�=$��-��<���hl��ƽ@���~K�{����g��U��g��A!��z�4�fp~M�p�Lh������e���g��/����ĳ�M�����`>�@�};{���{�êY�:�1���kWs��o�c|�g��ｵ[�� 
�^��Zro���uwe��&��8t����������{�z�o����t{�\���<��0hZr��X�2t�<瞞��#W�%��'�s������c���<u�~~�ڞ\0��zn�o�ǲ4��g�a�Y�z��S=�7���Y�O��N��/P&V���4{<�.�g��x�O;ݮ��Ҙ��g���xù��8������s��o����i�i�|�r�0z����}���,��w�v�r��9��o͕gL�H��l��ӷ��;7{=��8/���:����ٻ�� �r��S��8O->@�3uT��Ծk#{��2�]�����;l�!���s���� ga
a<l_P�?. D�bw{����{���>��u]�Xf.03d�J�Zy^���q�_�f��7���7�򋧁jw-����~f�Ʌ��M: ���3��(�z|BkD�ֽ,t�,ӌa�b�O}����?� �{��ƌෟ�'�����+�J��m�e���=OK��
�!LMt��n:��7\�7y�O|�|v�O��*� �ب,�Ĩ'��b�E��PPāFAAխ����uu��l�k[0�o�+$DU!�dư���+��ūh�UAT�E�b�"�H�UU�\�V[Ab�AAI�Uc
"!ĕ�*ADE"�B��VLj,X�Z�"�aD��qF"�,�~�µ�o0*ZY�*,\���k�b�XV���Qd��jTF�U�U�J��r�M�Z&ZJ�r�*���[a��N���S�~�Im�8��b¢��b��W�.�d����`�̥� T��bDLu͢��j�,�5T.�`T�E"��m�ʁE@��Ɍ9aUP�u���?|���T�W�VԸ&�ť!���n�f�Ht[B-�=�e�����Fm���U�ڕ���MXs0�/�2��&�7D�@���m��f,��u�o&`�36ݠ�A�6r�^��#N�A�#MKP� �Mj�eJ�c�����ҡؙ٘m��Wdu�	�Ƅ��XX5�cR CL�v�5#��3�A�����D�J���]A�[�܆e�ЌRBchnr]���M����ҕŬ���	�j�E�5�\g5�2�-3�a��V�2k��K^Sm��Yq+J��Ƹ�I��	�4�cMU�E�3A-
s]T�6�(Bk�̼�@]G������]F�\�[G�K�H�eD���1�XĤ:�4��l�]�@e-.M���8i�-�K���5��M.U�uv"��ԅ�,U*U�.̭+ŵ���S[\�08�u�a�ܪae��(���65`��p��)N#hản���țj��41�5���	����"�v���d)íl3omc�4�vZ��K���J�6Z��Uv�f�˜��²��^S=hU��s�nh,2��0̱:�Z�t,Q�F5e�B��ҦX!��2�:�)��)S74Thif0�j�-BlBZb�^m��X�����cv�����Yp�Zm�s, ��nh�� k�]]�mֽsj�a��iQT�X�l����Ͱ[�:R�٬3X&�,&bf�KX��M��)ur錅�\�tpA�K��[��^���%^%v��l��u�Z��3Xj�=]l%�4 �L<�avk�,p]��7gX����,�2�B-åҹk�Bd�\X�E\�4G8�z�q�DJ�*�K,���)�)�2�n�[�x�8���˂h�{Ye]�:�$��	.�lp�l�ݪ
Y�	a.WZ4ZR�7�2���.�ګb޹2�;�+`�-����%ж�TaUլE-ѱs5��ܮUU(�kD�g�g����s�[X��V�i�a�⍱`�TѸ��iT��&bf��J`�% V���Ļ;K3-��h˰e�a+n)j0?���;Z�[��y40��U���Ձvs�&�b��	�#n]6��Y�0uA4m�0�WSC�`a.Xm����$`��j%��,���P�����lb�M3�m��0[ȱ��]��Ѯ�v�����3p���h�9�/,�$2Gh̄c3�J�X�1��9�J���r��.��t�S�H}�o�\1��gdHt�~H���
͡��	��n�#ċmΑ|��'w(�t��g�t[�j�U��M��� �m���}	��ax��v�Qu]����>��7�2t�8�ƞ�	*��A$x��aeQj8*���mBI��ɟ	>+���SOH��Ap���B�b��GP��G*��|	'��u�G��^�7>rSm^Ԓ�t̀a������gs
�ׂA\�#�y�Wn;llC�wL����+[9@6�J�%��AP��	��;;���pcE���5 ���:2̋�m6N��o�~��=�L�ɢ8�^���@��@��36�
����5��-� �_@��WΓ����Bsԯ�R�z}K�ݳc7�l��l�u}aO�,�C��0�Ü2*�\��S=���~��Ļ�L��/wZF��+�%�gG.���;^�K[���c��N��	���lA��ϐ�u5���C���(7&����3��5�q�Zކ ���㸦i�Ԟ��$�v V�r�>9bAfN��˦��j��2B���)4H$E�b�A�����au蛊豨ϐM���ߞ2ˆ �p�k�Bۆ ������eh��E4�z=���-4��3�u@$�]�%D{?=ϞW��I~}0OC��05,3xT�����CA�����mZM�tka��e����'�/(gsT���AZ�#�	-��2@��v�ֹ����r���Q�Y; ���
���$�_.�X0<�]��� �B֫P%���I���|l�ʙ�3'�t�9HD��ʖ �Z{r$	��Y�"ȝ���
�KU؜�O��ݽj(L���>Cs��L��Pc�:A��mi���r�z�3�K��{�Ճޘ�|�h�� �?�=�k�$����P�@m��%z��AN�N��;РtY�]n;#ׄϓj��<����wD�_�"[�7�D��b��K�v(�/��� �'N���m��$x�Uw@�C{r�Ut�Gb�Z	 ���H$��@ʅ�[��X�Q
)˳���|��y�6",�.�M�r!�&�Vg Va5�kWS3�w{�|�p��E����M$�{΁$.�7{G��ζm[7-��ۊ<@ ��rd,F�r�g$�;��T�Do�,�wS�씝� ϸ�2I>�d�oM{��q��f��/k�R�Y�N#��vH�;�$�v�	+�#�|H5�x��x�7�HY-7�2A ��A�����3�gI	��u��^�v�����IgzȒ$,Έ$������:]�`�z̖w������d��Cʅ���?{�p�{ֽf�sa>��6ú��=�_d�T���C?���>�ڨ��G���	��L��M|S���wN����p ���>U����ي��a]�3$���� 	�yAC]�_V�R#��~x�i��e���G��E��C]��1*쭅#�ÀK��su�� ��=�5�.���O�潼�>W{Ey"Cso(�~E���HSQ��`�J�؂3��;Jt]�賓@����a�iF8�u�ٗH$��q ����	���j�Cb�	׷��D��������fJ��9��$W8'����VI%Wky��T��~1�B�Iڮ����E�ܰ���z��y��ͥ�b6�7䙧�A�$ [����}i6�L��tG12�7sG��i<؝1o ��!#n�l|P�M��^flo4ř��.�#Ē;]��'���� /V�բ�����]�=��U��,���o��vph�^уٺ9}	��K$�������eJ�͒`D���\�ī�6:�[�ET&���K<���Q���8�p�q��nV1���^. �ohZQ��-)�����%%	c�V�Y�f�Q�B��f��X78������`R�:���r�6f�V�����\�Ң��.aҬ6mt�Te9��B�P����YM@XS�`�4�s4�4�Au��-/`�3RԊʕͥZ�i.R�G[9�mu�&�0Mw`.q��M���3n����p\ʪe�aJgK)�Z5GXi�{(\#����φv���6ߩ���{Y A$w��k�A%�{�J�ɪd$�ֳ���� ��l�B�� �L��N&Wu\ω���O�ܶ�m5���$����	��3�A9��\�G>y5�쓸brd��~p�:0	3`�D�O�ٶyf�$���H$Gwtɖ��3�Y��H*{s��8��V�"�s� @1��>�W�wBz�uaK��������� �~��� �ܰ����L��A]��y������L�� �#2�gĂ�@�۪=vË�v�L�`�!p4v�l̮�cK�U��`E�U��n�nKV;�Q���yg)�9��H$�n�I �B��a�mOf���c�-�	~�ɒ@���fw�wg�>���> G���òޢ	��}g-���e� E�1k n��;i���1�f?q�9�
���FFh���3���=~C�����E���hl$T���t�K�H$�f}A>}�@��@�`��f�b�ې�{16��:�RȻ��Ol�X$Uw@A�E�	�}m4/[;�	��2� ���H�t�3�!�'Fd����-����K/����	m� ��z�!���} "OL�&XGc�A��C&tfAS�	
�pd��u�]-�1>{�ɐ ��q��� �ǫ��~lN�7��!C7K*.�4��-ò��XW YGlŘ�kiF��QD�i����Eӹaضn8�W�-� H7�A��0�4�����3=4���{��H$�Έ���y���R&����h�YΪ�I�Ʒ��$�����|���s�o�R�Q5P�����gw	�wg�A���$���q$��PKm�g	�ǰ�9� 5�̂�SA�����nl4f�H��ɊJ�'����l�ة}��/��~_������	�{D}���ĂJ��J��|���H S"�S�=�Q���N��ߒ�}�A�� ���ӻ��4n7/A>;�Q<ϣ����9LΌ�1ν~@��}�$��nR�Y�f�b��AS��@m��j��,��n��i}�� �ON�F!m3�Xj�W���s�h�Lh�3,�bbk�&eW֋�.�7��dΏp*o��$�f<I|����d��c׺�v��؁���h����N��q2�����@�ѽ9��� ��@��xވ�����e[gC��0alS--��S&�ۖ-��$&Mmӈ��ۑ>$��i`�[*;7�$,��� /$wt���wwpΓ�8vz��Wtv��
S�ˢ�=�H7uo�ē�������?��oUgMT:֊t�� ;�:-9���w��}�"6�����A[0-�ʽ�N֣.[a!�
%�Eh%����>��+%���D��	Y�r4RI�v)��ߪ�|I
���=�2�0��X�M��K�n̍�@���a����܍����m������a�47W���Dt�3�9�w.�ƅ���o.6ͩ�z��=|L]R�Ӂ���I ���	x��� �p�Ɂ��l��W��i�Ē_�6'�X>�w!��C&tbJ��m5+͉��k��q~'����@ K7tz9�5�u������tpI�,ˊ��0��q�Ă�4%���ƍyO
'����dH��� �fN1�,[�3�HKz|��w81��v���A;�TI �V�E��$7o@�"�^D�޶l>�%dFL�{5�����t�������|�-{�g�Y;�j�mh��́$�}�[��<g����;{���b�K�Z�d3#0З��R�@�of:.Z�����x_u�f��R�^X}���䯼{�gL��䤚т������q��q�T��x}x�BA�\?SS�a��#6��GCQ6"7f�b#̖��]F�k�rd-3�3A�d�hqc��l
тǊ�@�0\�cE��Z̈́�+h$h�fn�i5R�J/b��"گk;��[KB�4�+	)U��(�Le�V��Af2[��:ׁ�5�'F
�Q��&)Y�U�ۤ�BY�[E��D4�muHOۛ�ywa�k\���&�]�qepFƫ��������^�`Uv�d��Xh2�������-V_���s>$Ug@�D�Cs�dԥ�纲_Geo�> o�����n	E��}n�"{(�b�6{�+���My� ��~"�q9l�o����Xd�p��C&tw�^-O��.����Z�5�-�{4�H*�"v�%�p�a��X;�6�]1'cI4ؘ�I��x �w7 �O�w�[��c��Z�Wy Z�^L�c�X��gp��񭶨� ���⦱�Z}���K�{zv#��Vci�H%�{�o�(I�3���Kl��c�e(�w=l�,����^f�7R�ã��ne��7=���ٓ,Y�n��r@ ����H'��wfM*�a�������yf>�&<�q��`�S��ߛk�d@^��Ղ�S�������YYn��K\wo�{��2���U�g{��ۢ� �GD��縞2��Y�y��)�пL3Q�|X�!y��hnH{�_��_`�׎����E���wc��s���;ۮ�+���vN&AQ��$��tH$/%�+z��;�F��w�$�T�Dx���>2äۇ+��2gF3�Ou�x�s��3~#��S-P�*����V�X�{7A����A#9�������0r�ø��c�L�I]��uւ��	T�G�m��H!os�6��w8� �J���Ј��K��hĮW��)@��b�Xܶ�K�8�Y�r�{��,Ȅ��2#��9��[w�'Ă|J��[�T�S�Ջ9��CM�L�{����wvw�=\�pJg��uв�7��D�>��� ���K<[1��y�Il4�z�0N�;P5��-]�ė��<��o���{{{q�q�/L�������������^T�@= /��y3�ח�8��7u��M������T�/"}a٥	j�d��ĝ����2a����=�7�co�NzJ�ʔ�&����%��;j�k>��K��7���s�P9��]�<ٻ�p�:�eCş@;5�������i�u��U݄��:�u]Bd�����'���ٹ^}��=�G�.>�;����Ȳ̝���B�Y�7}�hс�)�1o:� �ޗ���~�%P+H��l)��,]��#Ӄ7�B��e��ܜ~���^�=����c�������]�7��`�~Ѣ12�W�'��_�����k�s��w�^��U瞞�+E�/)�1I;���ph��R;O�^�C5r^c��7UOB��P���޾}�C4��W�y�����٨
���!4�zǛ;�x{���\..޲�{\��{[�/j+�_#�\�w�P���o���N��=6ٸm����i;7*ȷ�׽e����g��{�q	�hs�j8�>{��n���^�+Ŝ�L����ʖ��{�L��Q�Ϭ��-��;h�}�m�yq+��ݞ"M�X�����pc�jY,�bT# ў���.��ȱey�g��'�Q�\�{�;�)��H�ʴ�6o�V������=�9_3"���Q������K3>RvR��P�l˚��4��rr=�0�Z��7����>,�6*�{N�$�νkcQ]&�u�/=z�^o�o���2n9���X�-�}�e2������gO��K~�uמid�Z���n{A}�4߳���*�-����8�Qo̮�)��{��8�ȼ0��ﶫko�lu����-�fͱ�@ĳ�b`�I*bVL�R�<ۈ��`�Jŀ�SY`�YR�E��µ�$\�mT����2�r�Y�X"[u*EQAT�E�C#1
��
��0Ę�F�ݸ��J�T�@̕eH
T�Ȩ%Y*b\i
���R,Z�"��(��VGl+4IU�@����i[����lZ�j��!Z�*Z�冤���
�,T���1*8�V
x��)*"(#*��HWp��LI���[E+"�
e�Ȧ*�F���-7!Qb
�
�XV��\m����m&�rظ��E%E%b��.",�bc	�}���~߾S���v����Dyz�bir�/39p�����w1�re��*����vd-���M4q��u�"A>�=@�<���9�����o=�[�l5]ة�'#��x���3�A�"-��G�FV��r���F$ ����a���3�Iϴ*�ܶ-KE3������5eҼl�ku������d�wd�����]3�A �̀ [[�@7"�s����l^{k.dH$�v��ީ�M�����B�|����8nt�Fu/<�LX$A>n���#���_�I&�7sp,M�[$�V���ܔ��׫�H�Ի�
���B2���C_dz�!sw(�$w��-DP(	�qT���,�2�S�0Z�t�:o\�h�I �.k� �彽>����]5'C:vX�a	i�����k7��w��Ҥ�X�d��ӯ@v?����ޘ#�-Wp�i��`�>|	19`<w��_s����vN(S�O���bAWʷ�ƨ�$>uDx�W6j�IY��>6���q{��}�o�Y���xg.�b$���� #RV\-�P�i������[nY_��>|��5���Ɏ�S��J�yH!v�H��Wt��y�񺞈��ؠ�7��.����d��vUx�?L�Y���vDJ�PI+;zd���Ӯ:VMd6UA3I��3"�������3�|I .�&�+��	+Uj�H]��$�z���S��$�viN5��[_S�y� ���A>-��5�SU�7T��|ޚy�#|��ëQ
�p�Uyt�L�-Y�1��BM���� �K�o�2<c��?w@�#Ӄ,��Zz�T\�/�@�������u&1Ej�nA�v���;MP'��~���Lhg�==L�7��Qr�>�.B�xI�=��AotC���>�y���xsm�.Wi���Mu��"����m�u,�L�m��LO
7�J�i�<2�].��P;9�I��6�����L�2]�*Z�������1���996f,!�"[M*Zhc���D��a6vt$�U�ii0��1j�a��7&4jkf�X0��2�F�	�R�:�\��\����ޢ�+jƳ&q�B�V�� �	��]�+�mlgy����%�+7@��WL�c��f��ܓ(�l�_ߟ������2�g���nCZ�%y"I��6e-��SG!�!��A2�)[�H�r�ə ��A.�b�ԓ���m�>$ӹ�>$����;f^0e�:��,`�)ك�ĉ6۷"I-ۯ �E�2�f"��O�f_L��D��G�s'yӳ2!0t�	�X�jM�i�}^�$��� �H-�� ��_�n9��<�$w�xܙ�����9I�i΋x�]� ��8Y�ދ�q��j'�'Ē[w�n�:�0���$��u;�I�;������K�m\���btlɇrY��Â�����`V�H�P,�qܪk&A$���I�ޏ�y�!��Y���3�"�r�OyA|}�>M6����8NY�ǥ_�7�|H	�]1�������ɘ/}u,�8�;�i�����yqX���F�\Y��[7s�Q�OJ Q|ֿ�Wk�����ͅ��<`��_Y00~�3�>�I�� ���M�@�TC���~� ����V�H"�C393 �Έ%y͘�d�rzb�7^(DGd��V��D�;�& p�����r]�ς��~�L餙'I�Cy!�Q �*I�� �D�oLTj�S3���Dz����ٙ�;�Bd�r�$��w�13�T�3p�:�X�]�DW����u��$��L�:pԧ�x��ATO�Յݙ���ن3k(��s�0Δ����3J�j���L��r���Β~�c�A$�g8�I����~;R�*��lu�[n��|�Oa"AD�tS��kUt�ш�zL&d���x�{�>'�6=��D���=gMꋨ+_Z݂�;�E�8�0��>���;�#Ӑ�fs0��&��D���spI�O�'����ۡ�(,[PD<����k��V-3��v{B>�˞n��;m��{$-u����d�����~l���l�I%[��,�30q2T��a�$�z���9�$	���K�o)eW�V	�wG�D
�[Av`�1.�ze�v�A�ȃ����j|H쨁�@��ɒ�H��؇{���}>��X�ݩ�.�ƙm.U����NáJL�����#��s�X���|���526+�gq��x�$sVlO�%���Ff���:.G=��ْ'��!ӗd��O"|����M;�n�
i�y��ݱ ��ѽ��ũ�F9$��8;��>/�ޒ$�E8�֪�Iװ |�ujݏev>�$-�vd�_{#�B���`����t�&A��w0^���=U�I/ׯ��=��@�*yޙSŞ��NLͼ&(���������>����o���2}��n	Wҝe�;<r <b�/%�K�U�7Su�f�*S�6A}��?ftω��f�.�9	�8�}]	�$�Ƃ�Ⰹ�+Ў��L�A �؀I�v�=��r��B�Z*-�X
P'��3�eef�5 ��G
��5���h��#b��LAv������Bb]�w��\�!�#ݜ�`��ٱ�V,���#|�1���T���&!��30�2�� "r]ҽm�x���ݱ`��F+u�g��[�%ĶfV9~�w���A��2b\<�8�p �{u�ǉ�3���9ۋ+&�D�
�	�r="��Gz�F`�T�]=�uز����Q��	���	$l�t�>e[^��S9�'�;j!LS60>N�غw1 �SD@$��.�Un-�߈�� 7D�	Z�c���ͽ>�o��G]P�5r���nl{��]J�6���lou��4��yVfRl���H���w|����^Ӷ���G���9E϶=�I>���a�>��� .�)�����:9���*��Ή�L[K��-�,6r̀��X�:�[4M��	@hei-�st1��2F�i�K&���5κ���lK���,�"ktn��Lir�Q��Ee��5����dM����bRa�,e��ƙ܅*cR�<�(�B�T�l�TcXe��ݣ�8+sWl.e�@q16�R$t�V�b�8سGD��6�ɵD�U^���ll�&�YGQb��"�R}���ϒ� �.ў~qT���(��	ٽ2q�陘mpSϹ`���"�Q!^<%�w��9	�w>�޹��Y�KV[,݇��$V[A�c���$���oS�>d�"fqt�1�附ρʆ��@��Ή���V�_gc�l�$�c��@%�7�W�ƕ�t;%�Ȑm��b/�T��G3F��0��� ���&G���!�f��~Wyd�2�� �h�$Q%r����ʮ�$��؋��Maܽ��{��Wf@�Iy��I �v@�f��g%}��<;��~�]�]�jMś4�0����j�Mع�؅��u�K��Fgׯ�6���.��}�Ǟ�È ��܉ �	~��7���7��V��P�؁ �C��L���e���X9L��O��׀@�5f�Z
OB)R�=�k:�����:��k�a	;bDe��fǾ}��M�h	'	>�XP�|�[���%ƶ_9��ܽ�o�=�ԋ8��6��I>~�vo�">�\A�aD6���	3�k��ɉw*��rd�K�tA$��&;����D��K�dA�$uG��r��ft���7o0zE�Vr�[�]��$8(����x�;_�U�f)���i0k��8�=O��^��gb��y�X��A�>^U����J��1��`�\�	 �_��cč����nUy�$��m]��.�X�iP��eub�4HW/Y�I�4ŷW�H��`�ɕ�?FY>�Pg)ٗw����$W��r��$}�<g�N5"u]��T	dv�G�<ͦ\	�쓧s U���<-��kj�s��ĂI�Gv�d	���	�d5^�Q��01���t�8��[6O6c� �+ْgt�lCԋ���{�%+�ў��!x�`�+*�9�ײ��vnT��5�Y��"};U��ǖWu�5���U��Ɗ�|	�: �@?6��	�@�%�g&%�ͬ�C�����Q�}>KČw���B|��hz�J7��}�$���!�<4;�̃��L&�;w/�[k:�De�U�&�Oa"��#Ă}m[<_���m�M�|��dX[��ېH'���;Rv��m��F^��.&�v�m��ƣ�����ۛz�{��	A3��8~>=�y�|i��G�-��2�c��Dׁ��q��� U��O���ve���I03c��L�w�ē��>$�����'��\���$l����p5�C3;]�̀]�^%�;��D���1jn�A=_���� �Ke�L�@����$��2&L�hn&Ej�6Hl �j6^  �[��dF�n����l�11�K[a�4�e{�Lղ��!��q��	O���)�3�0�����f����S���s�ό�C��MH�����h��j�q���]��,K9����@��sЅ4��i�cz��u��Ż3bI$���ٝr����o���6m���m�1ݛ��򍠖��T��m�bAg�8ݵ�C8I�t��u	
��8��^$l�����k>�J���x��͙8{Ab�3�8x{"�@��@�w3�Mg"^�D�_22d�:;\@&�5KU�:��Kox�#|�Oq>�SN��T���I�"�dA���4۳���h�_+�$	�}�B�6܈%3:(���/��{��<�8��}��O�:�$�D�ȏO�_�_&�w�NC�Ѥ;�wʦ\c��v!��S�H�|x�B�)]�:͒	򉞙$�n��z�x�κ���{���?g��y�u�}��D��S�O�j��ą�Z�!?gU��חj�n�w+���Q�Fb��3R3�Q�FajFj�b����3R3�H��0�Ԍ��3Df(�#1FjFj�lԌ���f(�P�Q�#5#0�٩�f�fT�L����f������3S4f�jf���Y�53Fjf,�1f���Ś��1f�0�L��Y����b�Lј�S0�LŚ�a��Fjf,�53a��Ϗ����f�h�LŚ��a�f,ř,�1f�h�LŚ��b�LԳFb�Lњ��jf��.�f�h�a��Fa�f�b�3d�S0�Y�jf,�1f�43S4f�a����3a��%�f�������53Fb̦a��S0�Lњ��b�3S1f�R���,�U��Y����U�ViUf��1Uf4�;�tҪ�h��UVb��Y��̕Yۢ�颫;n��:J�Ԫ�UY��UY��UVd���~��UY�fA�UY��d�U�d֮��UN��Պ�f��5C1Fh�Ԍ��v��3$f��0�Ԍ��3Df(γ����f�f��C0���?������WW���r�U3B�m6֯��]q��������~��������>5�o���u����w�.ݯ�]t�_�����W�꾛�B�~�������%R���Z)�O�?M{�2��_���_S�+��D?���U���'���^���/����_�/��u����k�n���I)�bJV���)[3*�V���5,j��Y���E�U��Uhj��ZUYMJ�M*�4��LUZiUfA�J��T���_��#�W�Z�O��?Wk�_�R6����UmU7ʻ���]m^�_�]���|~_@Q��������W�|K�wZ����׋��z�~���TC����_����_:T�}��_}���������vJ>��goU��Uj�}�κ��vN�L
?������V~�Q.�w��C}/�}W�W��w��k�/���_?�����u_��}����}��j�V_����W���C���]Z��C뫿��|}�¼�ˣ�޺��U�oU����?T��W��e�����x^vm�����J�*�W���ڿ���{t�p���C�ں���t�P�g��}<?���������)��c�r �)l�0(���1���*�J�PUJ�HD�T�JTU!%U*UUUU*��T��%( ��)R�
�%DU)R)T	
\  �i�@F�( � ʔS��
��
�  Z �   ���ր�(/�                                    �      }   2+�z�*Ӑ��%�Hd  �
d1 �(d�7�׷��� �@  {�  �� �F zN  '��&�@��B�*�2@\�� x:U 1%Pe�"P��U"��gB�*��H*�   �        T)B���4RE�Х���s`H����3B�@E�4>�$��=e 3J��RE�СK�UrԥT�}�� y�P��Ct�r%OT� ^   y r4(��  H�b@ťP4:����� � @;�\��hPU	   <   �  h  $� `�S>�9NPN 4:��yj(�9�kRr��ma������ < ��{���U ��   7������e�k��e� �U��̑�6;X�g�ê^YsJ�������9;���s���'J�i�XP����Pi�   �        ޥ=5s�r���\��V�,��)��W9e�
�sr�j�\Ψ��t�� ݗ,UP&Gqh�@P7��
 }�{�<Y}l��+��� �iT���mä́u�����s 4�� 7N�/��VSK��A�B�i.�c���
��I   �        �J�]�FK�j�4r�Є��N�n �A3s�d+�uu��b�\� +�\�sj
n`p�B��A|   ��3���e��&� �Ү!�)��i��CB� �
de�@綇 0= �MIR�4*��RUI� jx!RTؚ� "{R��RJ  CB)�SM&T�@ 4 I����)0���~���H� x`��^��ᇎ�ʑ�9�@�$������$ I7!���@�$���$ I?���$BA��=�������}�O��#Z�m���fU{����>S8�3�K�!�λ�&7����=ثm��&3��<���ݡp[K�;�k��6�*6�7�����i�(3F����&�zۍqF�EFw�GRr�
��������rtv:h�X8j���-�B݆���e\wKM�P���'�)����HB3���T6v�;Euv�m�$w�8~�屰��@��₝�ssUǪ�8��dn&��fť�n�8�T3�.�u`̪�Os�\*�J	^ P��z���p����U����\zw\���`[:�<m꽚����}C���< �P��s}y���X""���̚��{i�ͱ���]Z��\�%����-�Flkܻ���oN�6�N��\��7&��7���+�\{������t��'ix��ݛ�AJ�,��!�-��*�V�,�X����a+��&��3�cy����f꽔!ݛU�½�pAm��VM��+h�)�[��.��9���7��f,��c���J��k�r�(�b�R�]Ά?�o+u�j-�1���9Լ�������'Lǚ�Ië
��)�ӶV�宺�P�=ye�5giќ�]:m�;
ڢx�j��뜃��b�A5�^d��F��3�S�*���.,+b���@��;M�ç榓��C��V]9�/U�gV{�P��j;#����'���!�w�n"sXy�����;U�:�;B�0�#��4Z��/-6-�ˡ�M����(��wLXj�Q[�p��N��Y�]��%]�7���.�o[GX�ɲ�m���n��n�k��r��oG����(�\�NM6���	t�HBwmP���6ë]���Xfp��o���?�1h����q�L�kF��i�wu[Ȟ��ɺ���2�c������- u�ڬ].������o(����1�8����T{�<��,7B;�ҹ����,!�3�kV]�i�A�V��æ��m�e��1o�m��+RI�\5h�r=�vر���vJ���L3w�����o��h�V��s/⒱h'��6n�f�P�&��P���!]^�P&~��J�:넡]o%@f��F(�L���ݏU�%�(�Nè�"��Čk��3&JK�s=^�^����ǒt!��NĎA����۝&�o$���,���=Vq��ly�Y4�=�J�n�0����7r�����~��4�1�bݰ��k�&[s`ݛ�SV���JE����x���wolx&���3��E�F���I�`�R�Y��.�e�GQ�	�$tR��6~�Lp��q�a����3{pv�i�9:�; �.!s��������a�UcGwWJ�ճ=(���	�hC9f]=�Ͽh���'Ú��|/���܇��&!��	FV�W�cw_�+$m-���{*�N.�	"u*X��d���X�S�+��
�0��O>�5R�0�]`�1��'n7� ^��x.�oH��sx^1��Y�����v���l��l�Z���븘 g)���=p�p�Z;r�C�-��r�4�
��)U�GP�qv���\ym���3),�Kͣ�Q^7w�r�֛��F�s����t��C7��8(�ڙ���=,o{y�G��N6���uMa�di:��0]�	U�qκm��w5�T'w/y�^����QJ.�]�֘�b�ZK��"-�af��'��47J��Ż�����Y��Ն����b �2Yf�<�@]�眚���+�qQ9�!� �H79N���N��]Ν6�̉/��6E:�Zyg�j5`����|T'w	ņ�Q�{��%:��u3K�C�Iu!h���K� }��:R�wk���U��#��������{��[q� �vmM��P��Z�t.���jȒj��8Y�uG8�nZ�'�"�*�vP�s���u��:7�
��{�	{�a�`��T�$��a�_F'GfÞ���opκ�ji2�,�9]�~k\���*������`�c�ۚ�>��]�Y���:s
1Q��U8��we�1�%����[�bKp��EO�2,S���#��{��r��YO yĉ��`���;5�M����P#�؅�i�k/4�=�9RR�]������i9oene�s"�#��ͻk:#����"R;jR]H�k]����n�C&-j��t�O8�pwo�r��vax&�B�9QFNp�ڡ ;�R@oYnڡ`%y���1%���ܴ��)#����w#Ows��9;��ͣm�u!�2��{�a�y�����:$Ŝj. K���\�(X�]�d��K�PS�
��J�݃�l�a\��ށ{J�J�#��Y���NHB;�[غ��F�S�:�6NN4�pG��<����	��)����o���<VSɋ��i�ϞI?S��#F�FcͩH*�GC4��y
PN���sz���zI�!3�
�3k�s�2u��L�31��6g[x0���w�R�ܡ(Z]B���%n�v���)�����yg�	�;*�f]����@���9�vM���]�BO�+�0�ǀ����E���f�{�7�I��q(��ơ�RLK�a�>^��}�X.��c�]�s���dx4n��&���ڝ2�?jJ�ı,y�w�v*�%B�8�W
�&R;_x��ip�ݡ'ݯA�r���e�8��΅�ʀ�w��7v�_ײ1�v�]°�ݲ��R(�M�� �J�l��ʆ�B���x{j����@-�:���#A��}r��/!�V��iŗ_�f��Ɔ�v�0gfّ ����ՋX��'�]�E�A�n7nn�o'Y�t�x�j|�uU�Kd\ ����"=�o��w4�;��NT$FW�>δ�����WO���VJ���C�����)an6���vҶ�Lܶ�\���ړ�Z���l	�(6k;�g�i}�f ���W�nGc�L�sF;[KV�������gE
ވ�r�8��[�WB�P������d���dY1ܣ�G�e-�N���'zK�K����L.nL�L�Gn<�'�n�pU,�ly̤f�UFs�ƥa�5�yͭwL��*��L-���{{:�S������M;������㋜�/ �D������q��?��,�3|ɜ�m��Z��Gv3�i�uLR!� ����7Lc���:�{�#�-<}�~���3�K$�,!oL9�	�[ƇIi�;8^�^�2�3��z�#g��Ņ��ড�M��k���Z�~u�\��A�+Y�pj�+*�8cD����5{�2���A#��jt��&Y��%��c��B��:�kBv�Dt^Y���pp}ݜ����S���͒`k�l�N�@鋉g�9��r���fA����̣`��K�D�P.Ӑۇ3!,3�UMu�&U�m�Y=��/VvW��k��hN���79A���!�&LF�hX�U ���~��)0v�p�cVі�{A�|�ާsD�f�&WD�)�"ٰv�P^�B��PɆ��b�F.�}1H��ECu�]N3�� �e0>Y���Cj�y8'B���1ې�,��z��˓z��q�ٹ�U��[^�f4�*�	��t�oE���s�e,pܣz��we��=��y\=��"#��^m����=�e;:�f�̊rmSr��y��n7F.��k�vX�!7zͽ5���j���0cQ{b�4����(�����S/JOE1�L�kyb}4�ev�	B(�D�w9�{��˚�Z�Fٚw\R˳��e��76�m�6�1fTq�R�Ѽ�_*�[�'54ږ��`{e�b�\���5@�LV��)M�&�x��;���Ql�Z�ԘD���^�l��"�Q6���B�}w�Z�m�V"�~�[/.��+��)��+vt�;@��*�Xy������Wd=J�ݳ��WVчv�C�j�[F$á7�tx���!f��m��M��oi���yvgUL���Nzh�vi�ȡ�,�N�)ǋ�ufv��:r��:W@��WE'-�ń�AP�w��(�a3�Ɓ)�b��Hl�ǵ�z��F�����D�"��;P�8��w�]ɷ{��������ۡ鮗g�[h��+��q��bջ�7��Y��"F�#�6{'e5�m�bTt�R��[�f��6����n��L�[�n,k����P6��єU�L`��\S9��
@�.�7��V@�,��_�㛝.��JO�Do��]�W6d��Hܮ���j���[sO@�SچQ�P�
nLӆ���'Xh@gLqU�҃��sX+�/4�櫚�3V�ʹt����b��Z`����6t����6Ft�������FX�!���PW#�{�Y�Wk
ekS}9���Б&��P,�9�I��:�F�7�Ȑ��,h�
P��ܷt�V��N9�r*�f�1P��˕���g7}�ƪ��3���u�l�<�X�gہu�qJ�F���{	����{{j;;nͣ,�r�e#�:[QN�:.@�i}��{t�ӲA^��2u#FMd��1Fs����;�,^��Ù���Ll����|���_K�AB���Yn��9�{���b�Mӑk}n�z�t�;${�<��6ol��n��
T�I�8��	�����T��OCɠ������K�cY;�����7�^�}/+��C�#�@�`���n``�CO�t���s3�T�.����ؔл`�BO[�-q����1��F4Q����I�w�U˥'or�ĎS�U�t�0�aK4��t�d�c^MtPY�\�ӔC�F%7y�k��b�#ɭ��Rs4h4<AUi�W*��Џ07�3E�qM4�ܽ�n��ywO���!��H�����{U��4�)Y�6���k:�3p��J�P��l:Q*�c��.tsįL�	��y���()6w9��^���T�["�,w'1f3��2���`�ȅ�ǰ��#chVo���s���4A׏4杊�Q�{�d�A�v^k5i64`�3ww�,]��{��wOW aJ4N���z���5��6�8�iɯx�q]�d�I�;s��
�r����e]+zX^��:�R��ҥ��x2�U��u(8������P�I�T&��x��5�0^�7���i�e۠x�G�X�k�NJdH��1��j��U�g4��)���7��,���e[�^6��S�9�:Y�#j竖��K�S��˦I(/)�ҹ����3f ��l�{��B�j�w)���Z��;�����n 8��hL�����	�*�5�h�ɜ0��*���˴���O�Po%�r�<h�}϶ۺ�`hK�K��,o��/�X�ˡ\��2Ɯ�"��f�껻�:g=���,����Tt��e�4ܼ�[A8C�	{̻��仮&�7m8�x��n\a#"�D�]��8����{j��D[��39��n%whRُ��;��F�f��F�
��n��t�m���-9nݗ9�Q�	�[;����j������
<��.Xf���l���p�TX
�2촁�gcx�\�\���L�i]�q	��n�78L8�J0򡅭��l ��B�D�`����eӱwcypR�E�'�P�'h�,#ovhۥ�\RK꜒�b�9N,�MC4�.��#��L�f�k�}Vǎ�e���o�\ʆ���,��^v��d�s�@qMw�ޑ9�E4�p�=�f��k��n\w���rn�b�r����L�9�̋����KA8�ӝ{R��P\�7v)���Z��`N�gnk�f�S��d=-l��g��&,�glђZ�8uJ����*k���HF��WX�1����E�N�\l�{D�ĞGW'k@�K��䋶�˹v���Ӽu�1���20a�u�lG;M# ��.��]I�[oQ��ܩ!2�=�]��Mբm�x��lM��ҝ��mhP�����\
g��P7�8�$(�^+�Z���f�gd�����S�ˬr��:^��4��I�4w8�4�1��a�v-f�Q�\�޽�u7�����apYLC'ݹ�:��[��M�,Vp��Gh۩$&W#
@��t��`r�U�5�l�s�9�٩7z^z�kf�3�iN@Ƹ�v���2a��	�$�h�D�p��R���*v+�͡H;*�d%a�r@�����׉>�:g�8۫�0�N?+��c���@e��z�1��x��z���lD\ݻ�f�$�
Y�e����PfG��7z�C
	A���A�����ǘM�V�ǇT��9�T�p=�w\�`���̰����Q��yPq4��S̹��^Ӯ��.6
j����K�^�>�N;}\)E�9��*7o.zڍǜ
����Wx��M��g��:'yf�󢃹.�rDw/��:c��8���x?{�i-�$�^��&����]};�٦��+V((+����=z���k9N$�]�,P;#��Eeu��7ZG�U����1sW�K��,��Gw!N�����m�wUb�D�&� .����W�9�_h�2�;�)E�ʺ9o�-ލ����!Y �$ �
J�!P	a �$%@�+ � �@��$ Y (@ �
���I Y B,,�XH ��BI�Y�I!Y
�$ �!�d�RH��H@R"�H Ad�H�J�$+	"���$XY XAa 		 ,�,E  ����	 � �
��$!P�a	��(@Xd@!P��	 �%@� �E$��H
@"�%I EB�V@
��$��$�! V ��� �"� ���E����$�,�� �HAd�Y X@��	$
���$
�����R"�I"� ()O�@$$?�B������������������5����jM㜔80]T��}�=���X7���wwg_g{����]640V���S�1�tMRںD�7/���n��.�/.��Y;�6���۝�3�x>�-��	����S����;�Ω�#sַ��w�z_{�OC�w��P�u��]�n��o�*��A�p"s���׋y�m%��J��D���{��t0q������h�����8�O�����g�6��gln�ͦ���n[�s}�-�͠���2�q��K��z��í8�g��ك޾+$������p �PJ~]��<;��xt�p����)f��{�[��E���ڹص��cmZ�*����ͭS���0+k6��Tg&�n�uh�a�����5�gK�_dx"	�ν'��M{̪���v�;����ȍ��G�����GL�c�3��V�${��N�|n�m�6��~���˭�:����=�"9���ʎ��:����d����l}�3�@���G�ͶM��n��8�����Fx��௷o��ô�����C�ð]��\�Y��͋������< %��,�V�� �ղ�bTT\����"����z%��+�s���[=�,žo������z����c^�0��A��=ą ��~�A~^�h�,�yc�+�107\��7,�[Xa�+��#��5vN�
�w�����>ި���j�Ɋ���f>�-��M=چQ�rb�<��զP�����}}j�����\���m��d��wG 6v�u��eE�z�q��Q�9�M���I��+ۻ7��
�r/v`��K��"BP/n�q��ڗk�;�]uq��&j�ڝ��z{����3V�W��=:�cr��s���ᗯ��m2�xn��K~.�u��-PH�J�f����W��n���N�:�,��k�Ԯ��u�~���ݦ�"�'do�����,��!`Gs��N�se�G��G���޼w �0o����C�	�O�n��7ח��-B����3v�k]��\;��9֛�K�f.c�WR,S�\*�׻�أYaZ�ͳ߂��nA��yw���oc��;_�W9���\IK ���<�f��CUN��#���Ƿx�h*,)�����o���cئʣzw�EH��c
v�z�{�`E����R���Y��j���'wF�X�2b�,�$ĝ�;L�'�Q��<:��;�m�3���p�����i`�-{�r�|�OJ�[N=}��=_+���DO��1Y4��=��q��r����$��=My�������9x�d����9��>K=��Л�x/<�m+��~����k}�\>��+�ݍ�[�|��(uu��)y��{Vn�����C��p���{Teb�w0�V<�lPļ�rۺժ*	�^�ʕ�n�m�s����G3@sS����7�q �ώ���H#3k�;�����{�|B8�3�b�_(�#���'q�+��O�r
X��{n�1������8�E�����r��9�	L4��������9Q�}��OY�9gd���x��;��gh�8ȉD<�!d�E���_)�=��3�AvOH3��|��k�`���ӡ�8��~�v��9����[G���]�V�fom�{{�t�g}�ۢ����P����"�$�?W#�g���R�)�W��K�/$I�/v����p�Vd��.6�Zî�����&�z(Y�[Q� =����n���\��ӫ$3�{�}��[�Cn����)�BnbcV,qFo�и���v�i~�G�w�	�g.��7E�M���:v���x��h^t����əٌ���_��7!�T\�^r���rɗ�� �p�sn��#XP����i��`�����l7 �,��x/N~�y��;�/�#���⳷����MMD��U��0��:4)Z��4�P~\9����հ������C��O������Y�%��ӃR#j��g�t �,#X��F4v�������,��y�;K���kV>���n���Ο<�Ï�{�@e����b��G�yw/W[g_w����� �/�3��
h�7���֣3�4hs�˫���u��sÖ�h%&{���v@5e��=��H�ؒ��M����]�=}e�qědj��{���t�#��:�+���c�U���#.��xxn���XW͝�f���x�Pj�o,->�]��q���q��2��{ۃ}ޝ�����;t h2�.�T��Z�I�n=҉�]�S�ţ-cx����'���J����{ˋ^��Kyg�c{�nS�yXR�����7�wa��ˏI�o� ��u��aD��Xi'(�����9��O:m��m����=�m)(�3�v��/;��K�ˑx{uE��Y����Z������f��3�W�gC�{����.=t��ɵ��;�΍�N��u�ݞ%;�����9�Z���9}��G��Ov{Ny��ݾ�G��l�{���b�N����qo]�7J�W�r�\�Л3�f �F��Tk�H9�,�1�˃F)|�<|}/Xk3�B�N0��c&z/\�Ǐ�~_��'[��R��}�>��\��^����߳q)Ǎ�G=�����5|9p��-��ڡ��sY��0;5+ug��8`S�n?Q/���ˊe��o_$��4/e���$PH�:ۻt����\�P�<�i�z���EX���H^�Ƽ=h��L/�/���;��=�mõ���`*����ƹ��Ԃ�,Y��g{�oyh� ����s�"�M�G�p۽�}�oc����c�\5��!��8g�����:�(5�p�{%�w��7��v�`Bt���K<n?^�i���{Z;�A.n��b����7&�Dn����g2��i�T`��1g����'h�O��i/;�|��F��U�XA�T����nY��3)�j�茌�cmV��X��cu���v���w�i�\�	�K����ϱ�l���h��2�	L�����g����b� �5���8=*�j��YwA����\ů���>=.�z�R|��č���P�#z� \�m�<���zo����Et�<N�'�<���	�y!�����:�a�(�e�Xշz�����7A����I�F���֯oD��o.�o�&����Z�=Ԩ��cggw�,�×�{�<rQ�,H���W�5&��;����^ί����=w����2W�����ߥM%-:W�b��f��yg�h����KZ"(:�����6�϶��n�flf�#rg�A���x�,�C}0m�g'p�^L&�qٝ���:�U�2{K���f�.}}:ע=���O�@;�����=x�dr	#�Oe�����]Y��ݞ�.��B��2���ɴR���sa=��f����8��?g�x#�ɦ$:��l��ޣ:�P�wxC��p`�/p(.���C��BꏎM\c�h��˻�.zoS�_A��`s�+[�^-�}���� �eZ�vɥ�.�� \�g�����AH�#�{ƽ��{3h9�˜J�CI6�v���H�����v(��������9��W��������ݸ"ݼ;K��5h=ۧ.��c��+�?Y��vQ��<"�t�3,�F�EPS8����-�ɼ$o�if�L*�հ���93unh���ل.ձS�zQ��ٖ�;o����f���M�y\�M����ۦ�/�{�s��۸�r3ߐ>Mv[� ;�����Y1�'U�S���4wOŌ��9���������B��}%��f�ٮ`皰�np=���}O{�N�=��&yxf�wg��}�OJ���r���78?Q����J����{rynx��縤��9��1Y�]_[csݗ�W�{:ed7�q����J�6�����w{�5f���hs���v_i6s�Y~���nj@�1�V��Lr[�z��4�ؽ �/[TS�ܨV�Z�d��`�H��;-���=z.P扥��o�{���Y��Մ��;����|��v5/=����;��%��۬m���+nsa�Gw807v�b�D�hw}I�=ḹ��mP�UPb�_S��G�޽���?w�Aް�o�Y׏�{k�{�R�_� a~�5�]�sܼ�l�������Ӊ��-��K�F��>K��:��#l;u5��'�jA"��ZJ'a,Un�F3)��G"�wkv=�K�W|8G�l�Z�5�Ϻ-@UU�|���2G��s�Ow_R}��G�+��"���9cx������ɴ�=勇��⺯����d�ePsɮ�u��:nEn��Е�Q�f���*s^��2ic٥q%�5�#�䄢���=X�����}���.D���2X�z�~��O^�(�|=�Ѹ`�##}��g%��\�<��垈�tt��HŞ�ٮ?(�C=�g��׍��c��:^o�¤76��nn��Q���F|�#�DwO_����o)/a����m8���t˓����Vrۜ��M9z�]Uv�g���o��i��������0�P�pW��;Gko�K��fĨ��wq�*[n�'�윉��ۋ����w�E@�J�,���a��n^����vZ�����Ūsǝ�qK���ewXo����!<?^a%;j�^>���rF��}�{�Sϗ_b�j2�ۿ�,w�.�]���X�r�n�[��k���N��ׇOQ�Π_u�j�G�A��F�^G��vyI5�����^���ߔ�+};��u)<�;z�
d{� �hы�f�l�$篼'3E���x�o��׷��e��r�L[@�L�����^ٌ_2���o��~�A�Mj�w��Cy�T�[VF�U���
��d����)�=�0f\��nr�3�����w��|\~�K���x��D�����6�y���-H{�D���έﷹ/n�8�xZ6���#�<t�+ڤ]z�׷w<���fm�Ç�PPG���9�Y����EJS�"߲!@	�q*��	J��W�Q�t�vӯL���|��y݈
�NR7�h�tbo,�\�W���k�ˋ��N>�=wC�(���6��Ğ�o�����+��c��ۖ<~#7���Ǧ��/�Y7w��|���9��6{7�V	�Iz��ܓ{Ӷ>�	a�=VOA�cڎ��0���	��>��N��sM�;�cz7�&n%7����������ln��R���2*�CuyH��G1�zxܜm�lB�8����|�+�K4��vž>{:����.�{�uum;����%��v�1�r���*�8_{������JW�Z����=~����n��<�t'f��-u3ڒ�pm{�n/'�A���G�]�=�yUJ��)����)*װ���S�[͈�S����gnu����d�]�����0A�4��0���=nڕ�d仇�tÖMN�z��R��S��ݔKq�/o�i�)
���p���Vve���a��`�g4ϩ�#��,���^"D�ekN�-���2}$`�l5uPn�I۵�%� ڡ�"h�#7sMHay���.���n�`^�f��������5���|!�wcl��DG�L��fJ|�A���ܻ��R/����	�_����<�_ݒ�_A��6o�otO45�X�T�Vw��vQ��#�8�L{�{��[t<�s�6���܇�\�jɫ�;ہ�H;�#ʍ9���x��{p�܋_N� ��}�F��/���mH�^]��'h|u%���R,oQ��rH/E�8�3�"��S��؃k�ڍw<��n�Gg��.�Y��_*�{�F&����M��yMtd��	F<���+�*��3��o&9����xoZ��zY��y;w7{���GrD��թ�趴�u��.�ZۇYn�N�O�����+�#f�������طf�����"�<]�^^����ʲ������W�Uٴ��L@ ߧ����FE�p��p$���` �{��Q7�⛊�ͦ�~��b�lj�hɛD2���������u5�ۼ������R[��*{ۯ;�}{'Y{ܮw�s�����h�^͓;Zѵ�k5���2繥����:���f��je��
ڭ��U�n�K��z�����f�{C|׆���_+�+9���`�H-�d~��<�u�gY���N���צ�}�1�%��8�궟@q�+�<F�s�d�{�HJa~���I�ι��o{�Bܛ)���2^M��:�o�uP�}o+�z������΃����q�
<�Sb�eǫAt>�-AB�� ���G�f��w)���O�^�{�M���ݕ�ֵ잕�P��wc�ޭG��)j�<oa�|����IxI6�rn�{ݰ#8�/���u��;���ak�Ȼ�G�1��u{|�7E�(�y~G�s����TgB�y�f�F-�>�Җ���>ݿ�s2䭇��b�6��$����7���&�x�a0�H7���T���o٦�6iIY��KN�)m�n.wo`��菵������pE�rدu7�,<0�5���uQf�~D�\�;���H���^���{���:}�r���o֮���!����A���u4bg7�;���|��X�!K����d]�6��^&}^tg���v�4ݿ�~Z�Ϸi~� ���>�fz����� ;�
m`�Y���6�ȱ�f��ῒq�jm��	���Oy�a���p�r��+� �ΧR��Ɯ�OϽM��Ԣ�wC^.'�i��x� ����(Ԥ�����+��=���ǂ���jv�|��|P+ʯBY�9�w/b�=^��)��%p�w�;!����+��y��f�����`�4F��q��x�lK���pH"�(1�Og�������{w����(��m�q{J�ݣ�L��qﹾ�������y����:!��nK�x��K�D�!��A1���=��f��%��J�������>�b!�ݍ��U��l��t4b���������{߱����:u����ޣ�5k����8��瞄�!�غ�6��l��[�4mp<n.Mo!8o
��@m��f{a8�k۶qD��M\��mck�N�ݘ�L�lVx���=�o/���Ҝvvl���gs�F�/��8�76y�ů%�/c��n o>q��v."�7l�Ui��ԝ\��]�3�[��rF���n�>M�{\r�	�ć9��sqɕ��X��q�ga����v�hr��M�={e%.g]�̭��ۋ����6�[���\�.�<Cz�Ѭ�T���woF��l�����mq��mܗ6�l�M9G����4�;��Ol���7NSi뵭�{=q��N܍��v�[l첻��=����`ܛ���r�!�I�nL���ٺ.}<�w�qo5a���vW�.����M�^ȕ;p��2놶Zh�]=D�!�<�tݠ͞R���gk&��j��v懱�y��l�=�pݥ���n�W� 3\D���(t�n��yW���N�q$\;���l��v;�ū��s69�V^�\o��Z��`:	���8{1��p�a�9ܝ��7�l�aof����c��3vۖ��=n|lQ���v�y@�y��[T6@�T�k�XL��5�^�+��X�8��Vn����Q���/�k\pp���Λ\�+�]�nsی����q/i��/��p�q#n7X�g�i�H��`{{ZE�r�բ�ѷe��]N��\��^ю�c��wp�<v�
�G#���Z���Iݸ��\�[t�s6�/u�E:�7".��k���uu�H#�e;�8g�vC<�k��2��:�5�N��[v�m��q��h<�Y� k7:sv�N$6��O<;�n[�M�n���f;<��ny�}�s�ó���8u���R]-��z�vv�a5����,�^��;���_!P{[��s��L��1��^�K����2�� +*n�d�E=[��	��&-�[̜�Վ{c����ӓ�ny��&8ޗ=��uu���rp�uɓ� �f�c]�7n艅m��3hw=�y۷eݵ�gl[ם�h䋒�N���|i�r6�V����<�����ni}����طL[��՝n	E\v�[/8;`�l:��3Jɔv]�6x{` {�۶�g���C�g��F� ��gC�zݴ���<�nwR�g�0�l�tll�gq�a;X�zwj::���������vTv/rш�<v:�ݲZǞ�{;��εN�'�Վ�˓�u���c�0�F�m�]�U=s������rbMɆs�����듇nk�n4;�3�2 q�k��+�&�[�v��ޭ���,������»b<t��&�d�c&��xi��D.�ʳ[jwn��(&��%�6Ѻ2�v�F۞9�Gjr�БŖ�r��&ղ��=s�����v+�ݗ;��gd�=����8ӝ�p8�۞;��1�u�]���n{\�g;���{ʼ-��.B�<�;G>n�]��G<q۞z��Ŷ6���n��Uq�t]ʝ����N1��lr�h��q��ڸ���6�e��q�u����mλm������۫��OtOiN���q@�vmŭ�FЏM9f79.�v��3u�g{/\��{j3�c<-�7c�m�By򐄚�m��Nzv��]�����=ot����.�;�tu� ������j���m������npc���d��mY:ͣ<����:�����8[����$x��Q]p��W��l�q�}�/f%6��Pk�n��I0��u���tA��<V;��y^�v8y��g���n*�˗�>@v�ѧ�mÕ�ʰ�r�c¸��P�x�	m7/�����Gg���q���M<O�헬v���l�d��U�Fz�z���m�a6�\==��Wm��K�V�׮�ۮ���ݺ�Ů�z�-s�l��	�xzd7m����ע�d���m�T[-Ԇl�x��v�V���[���8olu�m�S�{fk�
������)���Q�m���CN�p9�V���V탫�Q�Ҧ��۷\.�Hs�3������9θt�܊�p�[���[q�ŷ�������"8�<٭�qҜ;�f�M��({zې�����mIxSOdX��G.#l����9Fz���<�g)۶��HɸLQr�Rd��xK��x��l��r۲=�9�Tjڀ�JHTMjTzN;)��N;�c�ӷrz�����zX�\����a�.6��ml��2sŸ7m��$�^cO
�&�;�m�,T��n|d��<O��G�ݛݪ�j������t3�7��d�K��8���^���xۻ	��S9]���6�9n3���K�h�t�ܢv�ma���]����Q���
嘮K)q��{�\tv�t �N����mdϸS������x ���I:+��3��{�>6�m��1t�	8�M��[�I�}��MΌ�j��qS�8��\�'�����W\���]�W����s�w����r���]��tOn�;^�t�z�p�Q����v	��՞�5�c	����1��yݎDg��F˛�2�W<k2m��nԯ&��Y��.B�ӑC�۷n7/\��O�N�ޝ�Փ�E�	�gj�	�����;��e����UUm׬{t�Mۅ1�Y2�y��;	ポ�7wcǤ�D�pmdk�O�ڕ�G�Qn{�q��\L�����FL <����k�n�bX6[����;vޞ9��psp��[Ǜq��u�6�S�qGF1�k�7�����:����n&CSŹݞ���^޷)�;upS�ngR��x��p���;Q(u�v�<Z����;��n-v�\�q�����c���7�\��B��:+���G'G8��x|n9�nƶ�}vyƜD�6���Y�Q�u��j�8L&3.��`y�v��k�\�z��v#zގ[gjx����j���M>lD[W��p�>��M����8V�f�J<��M =ZW��m�����ݵ�����Rs\�/2q؛��<��ؑ8�ڻn��6{��97n��K��ᕭ�<��c��,]�vV�O��=�ubWn�&���9��z����q�qo9��Z�;/]�6#�B�<7��Z�	.;grr(u[�(���3�av/W\^ݘ�n#'(/ ��VN�[Y���dS�q�����9z�u`ѣ��]ۋ��7 �6�7k��F��ۥ�#[.��1�;snz9ݗvn�8�ps۱6� 2+\�w,��V�w+��ŋ�me�n�`�l���=#��i�8Lh:���!��F���S��n�Te҃�����s�zϬ3�r��٭�[pm��l�;�Φl:lkQ��Z7W��B��u�uk�l�X6��q�����zc���g��ŸM�٭Ѷ�CZ�j�{L;���g�v�����y����m��CNx;�o-s��qh�'�*�qi���[ ��n[���zpL����w�.��Z��؇����uٮMj�b۱�1pf�]uhr �60*�ʶr�t���m�r���s��:��vO\[�p���[x�p�,v��s��[u�Ӷ��<�5#�vy�'`�['X��]��nJ��/l�m�6��5�J��7q�Z��>۶9����sQ��G]��K;m(��Wv�S�����vY�#ղ�&�azN"���XS����4ތ�6�-�g��ӷ�wn#=���k���B�[�R#�s˚����6��Ƣ3��M��&�spvj��6�#�I�4Z1�O��h��[lnn���nwW��<jo7<T��瘸88��)	��ni�����v��Я>x.�Z���"x�Nm��넸-��tqs��)��>#=�c�n�k ء���E�	���`�=����-��mm\��\np�^�n'�ru���=���h�ގ�=K��9L�#ŷ���׬n���7�ް=�[�e�$f=�x�ٱ�9w�ђ��;�o@'k[�T�,��Û6U{b�u�f|n��<��d���u�D+<'[p(�'�Ya����5��"l� n:�v�8,6�㱭r��<a6�Y�n�]�vꮶ���:���qe�c���f�;���cs�F62�ݙGv�:o]I��۝P;%�J9�ۊ�c%��`�`"��G9�9�8�7k�>n7A^:2�sn��Cg�Z����u���)�ü�nb�Yvq;X�&��uY��7ulKӶv��SR�<�{^�uLӲvm.�=�޺������5�/��P��Xy��۝�p�P����x�;-ɜj�]��K���;˽[���v�+)s؇�aϤ|=��(�v޹�\Oc�K��x� ǝ{4�=t}v���h��z���ez#��(U������#۷.���7^1��������{GI��i׌aY��%�8ێ"碝ۄ�m���	�i�rܧA�kv�3u�,�V��v펼o1gE��Ok��Ӻ΍����Cn���(�������HX�vc���������h8N�uؼ��J	s�cn���Û��q۱�z�"v]�έ�����`��b�ɣ��7d�KÓgjl�'
,��)6�[�xک�S�&�9��L�C�j*�t��;u͋eͲ�u鶳�U�k�1Rn�[c�.9�{[��c8ᶸc\��kn�n�i�c���QŨyk��of;��2�bM�m�J�gl�<�8�iv�5����b�s��ے�ݝwc��;Y������[�6����֌��\8y���O6�ͻv-��q�zp�2���wf�z�q��<����u�)$��kZ^85v���)4ڼU3գ�=�����p�Ί�(�H����\�t��uh;qh�Ɗ�],�5�MKrU֭\��������c9cn�Փ�1ԃt�\�.n��e��#1ۣ=���ޞ���i�����?�ό8��۷��a[T5�FԨ�L��j��\��bY��fc�5��̵�� �6.Z�s&L(�K9��Z�p��i�X��,[Ke�JR�Z�j��"��[2�2�QZ�K���--s0�L�b1�ѥj�9C0�3*�k���-�P[J��ҥf\a��pT�ԢŹ�(��E+�`�Y�`(��+���\��+ikL����8�`��9Fʪ+mh�e�*��AE&2�����ڂ	�����V0U�Q�s-l5J,��ˍ����ˎ\� ��E������˃���(�VZQAT*	m�5*(�4�[E���T����0kk�\�)��.��J��լ��T�AD���
єUB�pk2�֊5*,s)�m�ʥ�0b(�̹1X�����\�r���ʩZ��fbʕ�eZ6����у�
�*����T4ɌM[�UQ
��+j���*���V�U�Kl�qiU�4��X�d�X��I#�Zr�C�t����{|;mpq�����Q��9SWj�@�C&��W9�]���c��#[2�0T�Q�On��q^�h8�ܽql�wn8�	�AtV�:��r^.+��n�;�g���4Q��l���u�ۀqvN��Te�V�`����q�+��Q����k��\���R���ss�=�y�z:Ď{{[yv8�ʮ;�e�>����v�۝���5��;p.�8���ϖ ��r�-ҹ���҆��2�v�'g=����m�c �v�y�c�mv�t������S�(�"����n�u�c:�,]s�9��z���n�Ҝr��8��k�aȶ\WK�;1����V�D��3��k����ڳ�����f���ny�k���.��&�b.�NיM�e�n��k�<�C���y�nN���:>]nz��k1j�Y�;[<{�q\���<8�.�ڛƅ���b��^0u���p�;w\;a�qӽ�l�;zۓ7>���s��;�zیg@;����b��֐��m�����zwK�=PMvz@.�)n2g�l�Tj:��]�wm�n����(�����T�sġRO\Í�.����|]�����Y+a���d'���cX#]�Q��I݉��:+������[�o'�8��N�Z�� [��¡탷\J[ێ���6�N<m��pi1�ݳ�űڀ����M��^��A��-��܍��ڞy��qi��˞�8=����m�[v�p���ȯm�m�k�d2-.�9Pc���2n@P渮G����)��b��#���t�<gn�uC�U�z�A��[˺�9��n	K���gvr�5����vn�܈�5ͳ�En�#���nwA���t{[���6��ݵn�뎋vZۍV��ɧv�;ط9I]�x=v�l����}u���6��k�k���7F�D:�7TcMi�m�0;I=�7F�P�Z�7`��o{������s��ۇEL���2��`\���<�q�ܻp�{n��y{�p�Ϸ�9{;e�ySx\v3�&8獗��9_;��m[\p�1D.
܍�32YQs2���3��*�W�nq�r)񞻳���S���r������v�L���Q�}��PN6��{l+q幒��U�k����㍼>|��da^�;�3�pn DZU9>�	 ���*odH2#(9�����뺯	��TN���$,�A`�����('�'�W�Y�}/��}^���A*s��A�����0"[��&πJ�IX�E �ƺz��AS��}��3��.i	�ު��� ���A�a�+z�7���p΀Hb��� �B��	$,{�F�8)���.At�����b���a:�nz\�A �y�*����j&�Q"e�Ux�|T�9� �V>��M.��:z��5����� �-"9�݉�k�r��Z��sPN+���=���7G}�Z��$Cl�8]��˪��5��uW�<�SC�s#Jo�g�;˞����e��ac)�%��0�ퟆ찿k�'��u�=@�x�N��+٭�b"V�)� �[@eK�^b��@��[�?��^�p�a�{��l���cq��]W��s`	�)��$���ULeWe��O7�*�7�����,�.$��	1�B�4i��n�g�X���}��J��$DFwU O��/$JA4�������FOA��#s�I�>��گ�|ﻫ�e��f��Af��Eݠ�`�`1�%9{�.�;�GM]Y��$"�O�&#shP%�wP:��wtz�;�t���n�TZ�'�$�ޫ��s��k\s�f�������3pZt��r� �a=��ω��Α^%�wU�ۑP�3	��r��TJ�MB�I�Bp�M��� B΅���wd�q�-�$���D�{�4I� f�Ը���&c�b��R�*��1���}�4$��T�&�%����!�T]\�d`#�v;�#C�O"��0n=�A����;�������c�4�Qv:nΙ�{�!*l�,�a����;��U�Aw��F�t�[E,�$����t��Y ��ڢC���?�~���t4�c(
��I�=�%��H�fb^ߦA�o�p=FP�ޡ-/T����|H}��@�O���'+�+������q�ӵm5���2�rz��H��{^�!�n(����"�)�p.�p�\@0��m���eUI}��D�	S�>���E@�쪯^v�׉�
���@��uF��A�se<�u��h�K���>!Os ��V17���n�8�B�I�Bp�M�e�|I]Z���򭮀���w��۽T	�WW9'ׂzـ�M5��7�����O�.|.�M� NbI$�]��<�FX�&�-�nB���\���eI n��M׾���B���š�=�b���ظ���ˎ�����B��ؗ�rȓ6.����TN��T�J, Z�I��r	�7����vn��A�7�gnn��J�� ��C�� �˂J՝��V��!���az;Q�/M�C�����n�8�As�<i̛	8:<��&�xD�!@/8D>ʠH$����A.3z��Q7z2.�U]v� I%ms�f4�a�@�l$�nA�ީ�q���ؘ>��ɲ	]Z��<}�@g��y�Xـ�2�ĊG��$�M��n^� �ct�8t�h�L�B/9��>]Ut��9��>�Bz�Dj$��%8p�^�]v�9��~$y�H")�����$�e�Ӓ�	k�ɾ���Bi�� ����f�h���C�� S��$����I3{�C)�SQ�31v�	U#E
��)R��
�^��������f竴a�ۉJ�F��q{C��;b��ǯ��������~:x�vzw:@���ћ��u��8�NCƀ���V�3�0�6� �����	TeA:�S���.6/�!�Ò��p�7=y�;ץ[�-�u�c^ݼd��x�V�#��A������kv}#�]r�n�i�����-�(��w'g(�ۛ�gq��m\��y5������GZݹ�\�웑`Si[�G"��\ͱ���899k�� ���WC<��1��Ƕ;nu=���\�ٍ��Fٗ��exl�t�W~~~~�?��y�� お�rI ׹TA ���4C�Q<3�ɛ�Kr��S�)��x�ue� H�D��H �c
������]x�I�y�^'ĉ��$�5
.i����:�Y�!�@�l$�nA���3��>����c���y�1O2��L�wU�C=�B@��sF��A��m�'ƶ���&{���I
{����6����➟I��I#pm�M�캠H���ɦ�+u�k�S>$E�e
&s{��'�)�s��&�'���)G�[�%�r�x�7��v�v�9���\�㇞�=g���pY��;y�!���fp*����D�wM�� �v@˳S"���dd�Q$�o���$[z
�h�i��G�_KjӁ�]�r����"D
nbY���z�F�L���]9�%g�oZ��ź+|���WVl�E+Wb}රn}
�7��
��Z��=J�� �m���=���6�������\�1���a�D�buP'Ă�9�>$�j�K����=��<A���|H*{��1�䖚
a&[rmO(��t<�א ��T�)�bA$���!YXou_8�;n����Rhw�ÈH�N����I1��Ff�ׇtm�W,e���ē�5� �����dڻ3S�7����7[�Q]n �q�W�̃�0��ƞOm��6T�:�������ߪ��۪�'��Ͽ�TH!Ok�I&1�M��>�5�k�+��uT+������
�f��(e3
�W�^�L�Q�S��#	$)�$�}��(�z�	�{jzj�#�f!�
�A�W��$���D��1�EmA����,_i�I�gK绮u��D�Gs�Y�U*WF�c��̫�"�k���x2�!5��JRjCg�n�U��=��c��W�xJ���#;���l%��
��I �I��D~�o���*��$莽�� �;����ZH8�f8��A@l'� ���׉�oMRѪ�sz�ĉ��'Ē".��|�{�����!,T̷q�	�P|Xz��X9�Ӗb��q��c�|��^�q]�v훣��r?{�! Sa9��bG�#3j�>$;��RuWcH���7v�H��ʠT��td��{�u^'ƕ�U�d$V���J����Hw��D��n���7��[�H����P!�fu;�A�h@3��*�3)oX�A*3����{��M���C�'�W��Q��*�v�$���P>�ݽT	� ��}2����ЃWrc��e~��wtP�O�-_e�S�I��f1.P�[=�tU�oS�F�^M�	�"Z��y.��3y��7r-]�.��ެ�З�+
i$�'����j�TOv�\g	�9TH%�wUx�
��� uPY�kq��"�a���]꼆۞{nk�!��L��l��YA��%8K�$���K� Cb�x��U{�I7���$�N�=ע�^��5��k˪$�gt�"���s��)��W��Ks�
�)��T�N��b�z�A
w���:�gQ�F���3ۺ�J��1��a��6�V�]Q �
��>$��.����T�U� �v��>$9�O�u3�e�
������s�"Q �s��$��H� -{Փ)E��*tVX�յD�|�8!@��p���>!s�Q�=f�s&h�w�B�%Ns �oNx3kpuy�>��.�`�{\��V*h����{N`V��[6��`k���\��.9�;V�bL�Slp��c� Y�ί��,a pb�� ��tㇵN��Hz{�f`��nϓ�]��ǳ�Mo;�F���qi�t�N�<v%ø�cB�M��s���l�4A1������\�{VS5Z�mok�����<3�;���Y �y8:�#�f���WW<�a2��ݥ�'M�%n}�f�}�O�ݧU��N�s.�˹�K�$�4j`�v�`W��/v�`�}[lf��՝�c�]�냞�n�m���H$'��Y:F�����_�`xC�P]}婢$�;�A$�J׽To�����&ܹ�B�� �c]�\�6�t��v��X-v�n�:hB��$�J׽T	 ��{�uw��@��G}���M�ꁽ�rI%\�M|S��1����>+k\��{���"#P>�I�jk{.��3����� �S�4	�'�����~�,)H7nA������-�S^)�eQ��;��閸�F]U��^K	'ʧ���+��}�eky�n��ڈ{���I`"�i���n�tZz��q��Y�&�x�pB�i����$�o��$}�4��7lVD�\ueX;[nA ��LG���V�"���O�L`��~[:������Kgt��!\�����潇aw}%����=~�t��{.�+NQa�5�lŤsە�2h�F�i|mڌ���������0�W>�J��@�5�C����D������m��{�Q����P$���k�a�6�C�d���� AW��@��;�pS�Nh����̍�pkĘ��$������A��������A!�nU O���#�m�����v]P$
y�A��w�M��_>ڠO�woP3�
b��e��F���
��㵋n�Cm�x�k�Ja�3����\[s� 6�P�B��=̰�0Xm58�J�ޚ��S�bK�Q��J�ձD�˪ �owUm�3	�*y��r�|�����vx��a嫋�ۺ�{��$�S�~��"��99��]+�bg"�WB�	@���P]W���|IO�� ���2"x�KF�2���V�a�Wo�W^Z�{�<�<�}ux	��u��G��_O�_G�E��{��wzvoh��Z�w=�H{���Z��)��{�y���9�#�E�(�Wn2�1��^2�3���c��5A�����&�gYC^�l�|_�cށ�}�o�{��wG�,B�Op)���+�:	ņg��Tw�y	��:}A>�"�?c����[����Á�ա~���N���2�q�ؾ���!���qIꗸ��˽4N!��ߪ���/S��^��_׻铴�X�?v�\Ք�s�|�x��2ٵ��7��~��T��UFQ�鮫��b�XN��=�_`=��.zJP �^�������"�A���ZP۠��h���m1#�^���&��,���L�E:X���w��O�����*�e#4��/�$��o�0�l-~}4��;�-9�����Y|篤H<���#��X��sub����N�}i������m�wsB�	iM���xԱz�)��~�vN��3��]�;���I�IG_��D��ߺY�jmy1�}�ʴ{*jz�y��B&f��++�N�=��{�f;�	+S�3�H4�'�@���فwC�x���g$�̓p)�sجW�&�g;1R�g��w!��f��Ξ����^.�k��&�����g�-7yju�&�:�*���Owyr{�zx\3f'�w�⣛h$�kYdG�����F��k�����D�짎̢xA���O�Po������X��C����ݘsY��wr�h]޼:��ƺ'!{�|($^�
�k���k�F���̴f��-�d֕m�eZ�Vi+�eA�kk
�[��U+Ke�F3M��h�,c���)\0�[X.%�
����m�F-abKl�TkV҉mah�JD��
�i�Q�9��\[h��lY�9h-eDm+iGV�j��TQ��L]S�T+�%W2�D@�5�m�mmh�չk�-Z�#��j(ѬJZبV��"ĮcJ�V֍�8cF֔Rڰ���j�fdm��\KR��Q�JԭiX�iKkV���щ�r��dJZ������)D��V�EĮ6���,�2عh�V�kB��Jң+TEjU��.e���K����-��im�)1�(��*�s��6ʨ���a2DW��i�Z�"�V�ʍB��TRѥs2b�YE��Z�`�B�Z*-MR�(�l�lY�mU�Ŕj�V��e�����m*#���2"��-X���T�fr��TJ�% ��h�-�����=	]��D�Jy�A"$��@m��n$�T��"�m�W�Q��O\�Mx�A)�H�Z��3Xʋ���3����go����Q9��I�
l'Tnz_��}�Z+.�Y�㷷yH����IOq��s� ��V�jvA���+Л0A0��2���C��%{�Ʒ[+�t�]��Y�x���?>�T4��mw��e�By�I���PHvV����m;���I%>�$^Q�e���j*�S���dC;#��ENfOxIO:D�A\���6^P�K����w�X'��*T�M��ω ���H�ʬt��Q���	)�9B��T5�@J�p�"�>��ɦ�>Ǡ���$I\�*�woFG��G�u1��2
�&[ƹ��FQx��Kɐc���cB1|��Ti�V�o9�"�V����fߏ�oGj�͘�}R��m� �f9�>�1g�����ĚꞡD��;�4(�g��̼� �B�{T	�͙0J�rU(���ϕ7-y�l��n����8�'aq۵�ٷOt��ݍVqÙ�����~����%۳F��ŷ� ����I{z�����z2��K�+rvk�������C�jEu��2��4�T���$A]��@H]��@�8�ckt���`�e��e���j*�S��� ��4I��e���x]���H*�vh
�ު��u,��a�(��������$�[�� ����ޑ�����p�MM�6g�##���O�\,��A.�C��|H*7�%ɗ�9���	gwP�IQ|��Q�b΅�>��R�nIx]ih�74~Q;;6�2wa��9u��vN*��V5J�gn����+A�=�`�>�$u��u,h>�����^+m��ޘ�K�����ۆ9�@O���s�{z�ڥ�H��w�nn��	��vrgm��,qr�Cn6�5�e�t�5�<����[]��=���6����Q����;B� ���8-�j0n��cGT69{`����T���kv�c{m�Br��'#�Vk�+����:OY�q�:zy ��!�m��vH���c���y�G#�]�:�4<�v9�"l�A�:JH�k�'q$�f�|lY׶��(q��{������w=U���{m��@!^�O���$�?jls�s5T(�����	��yB`�M0�6�\�;���,��J�����DJ��@�T_9 ��C��vd���O�v��>�I�jj��� H*3��	��|�u-s9Z	�1��T>*/��}YG���HC�j�}y�������}A
�.E|�6D�A!ouUOe63�^�Lf�F2�O�zn�e0�Ab
�i����>rH$���������$�uU�HQ��+��h��tbƾ �ƹm��TnɅδ^�:.6}�i
`�E�B�e��v�"��\��%4����� ��$�@+{�h�+��ڃiq�T���n9'�$Ɯ� 6ن\D��]3��L�&�;r*en�<>ns���9��զu���E썧D�5�~v�?]\���{�\@M��
:DũV�"�em���̩|J��}$����"�WV�1X]H< �i�&Ú6�\��|
��� ���wf�Q�t�Mi>$��rA�}�F�DF��0�NSU�uè�뼰GݱFHT�f���ꪊ�v�6�nH�TB�g۔z�PXB��A�b��$۽"�Bѳ���$�xd�O�>ʡ�LwoM�N�uF�f��(񎂛�4�nN�8�l{y��D���g��նI<1��U����߿����X��G�h7�-�J$�V=ʢ>���P۳�B�o�4:� �%cܡB�NG�
@��h"�w�?�A�{X��s�s}n4�|����s��j;$�I��J�����41 �����UL^�MO�vI�u.��u�"T싙�>��(���ó6!�N&���]�[9��V^>��瞅��ri��2�w�����*�����?A+�T	'��}�F*F��pL�h}g0��⡎�yZB/eQ'Ĉ�ު� �
y�9��{/Y�l�wCI'/��);DlD0RpڟUw]W�!<����EY2���A�W<��揂 �"<�����ΤN���es~k��Ș�}�cp:~�=�R�BL�kЁ�B)C>������kcv;5�n8y�8:+��jK=������n��Ø�u ���=`XԂ�����H=)
���o�}�8 T��{�'������>��ngFJ�P5�����u%a��<ێ�n5uMnH.~־�~bJ�I�����9s��w5��~gY(ʁR�]~�߸u�T���s~k���R�/٭���������:�ߧ��B�^��F"���:��5���Τu���W7������*Aa��9�y�ݻ=�Ͻ�z0�%M}��l�N�T��\ߚ�rq1�����k1ִ�u�4�ȕ��\�wyծ4WגG�#�R [��EvR�B��Zf�y�@R
q��O}>}�����긛�0�Af�Kݬs��N�E� ��/CS5PZ:���q�������m�f��x�B�1�����Y����؅��x~���d�T5�?���:$�.����>��.6�F���¿��7��
��S�����,Y��1J��{�&�o��;Ĩ��� u*A`V��=��rZ@R	yxOO}>G�'�ϱD�t>g���-�y�S����br�l��hpd�x�պ����˧V���������k��	?w�߶u:�R+%s�{��P�J�V����C������k��>9�=I���=�gRtB����{��P
��X���4b#�����4g�"���;�q��\�@OH����A�`V�����*Aa�w�ۇђ����߽4��C�}��C蒰��>ێ�n5]:�6Ã
��9��%B��
�o�ۇ;T���0QY�r���>�x�0��(�y�{��H6�a�y�ۇ�+C�:drP�!C���^Ȳ<��� ��R��;��|�~d�����2T(��`������a�°�
��~��u'v?~�����=d�ed���<�{��������5�sN��:�@����;϶�+R-=��s��ߝ���s5����
�[7�w���*AeM�Ͼ�:βVX�P��~��u�<��ɩ���UO��h؉9��8m�d���c=����[�ׯ���\4��$ލ�)���?C�c�l��l-��J��:�1�l+��W0��B����1�Є�Q$�!	�x�\R<�`���-�J𺸸�n�A�5�8��c��e�=���睶�����׽�\�3i���x˲l��j;u�8L�qu��v��y�N�w.��䎱�������lvnл=�.��l.ۗ��w=5���^[8�>����5Ю��tn���� �\K��#�X��?ݮwW]�p��G<�n<�s����قg�ь�.��6��h6�E���;hݍ�/����(ls5r�.h�=���~֪�Z3���
���͇#IP����}�8��ʐP.~��u�+W]�������~y��]�9���A�!Xo�>�p��`WW~�������k[�����Q�A���Oa��r��7޳�nΌ�B��X��������¤�3��}��:�d�+#�=ޏ{��43}f�6g���wm,m`�b1�P:��o��vz��R�5��~�V��AW��F۪IQ�䑴9@N�}���1:�R��7�}���u���J��k��}���g�l�1�2j�u�m�#
��ߛa�s���m'
��V��{��:�c*�Y�~��@�J��Xk�g�����������H)�k~}�q���;����s2浭b�:�I�o�u;+(�YY+�g~�C��������M��xEIXY�����
*J���l�N�R
As�ﻓ����>ӯ�֓w������W`]G&{���yx�7Pp����tt�W7�;�K�-�t�������7.�zi�+�w�l:=H)-=�߶s����
��]��18�S��8~ӭk^ߞ~�bw���ԂβT,C<��uĕ��z{r���\���:ñ�oz�a�a�(�I����7���à/��UE�rcQ8]�{�j2(�w���/vrޛ�nI;#+bjD�ȳ-˚f0O���wu��^�`�S��D� ��������O��@Ͼ�����X�
�9�{�� ��~�t���}�u>l�K�� ��L���bq'}���:�@��2VPd�T}�(y�DG���d�������uϡ��V�IDϾ��I�
�FVJ��3�w8~����չ�3Fj���_���ޱ<\L�u �5h���l�ii
�i�מr'*Q������ì���{˟�k�~f�*C9��l�IXS�����1���t��As�}���ID*K���9�>��)�9���#ﴀ$�@�>��@�V�9�y�� �/�~�|,���ꙭ/w�"T]anK�۠���K.�a�gX�7t�ܽO`�[v��a��>�D(��%��,�"d�'�e++%u��ݜ4�IP�J���}�u �s�3y����I�~���Τ����Q��3�������~�Ĺ�4f:�@�Jÿw�l;���N^w����~ל��~�-��H-����18�R(&}���:βVX�P���u���y�s�<C�+;ΟfS˭b�4�!�W���pa��B��V���γ��eH(��J6��d*P"_�!IO�&&�nd�Q��3��ε���2X�1���^n�t��v
xVA񜑔��Y������'������(�\��w�T�iK���ۇ^�
��~��]e�\7^���dY���\�X�K%ed�g�l�d�T������C�:0�+
���}��:����p��<�~d�ed��������M _�y��j�Й�5\ǇP:��o��l:��cR c��E�g)_�-�![�txQ��}�|�N*eL�~��u�y�Hw�(�dy�!v�Z2zN����~��+� �x��ӂ�F��pZ�-��k6��{\[8Z��?���ss�_\��ݶ+�s�i%��}��l�:�FT
�����p�A+~c����'�aF����懁#���#'v|,���-��
Q�h�^�C�Q/y7�F3��w���wg�&��J�IXS;���:�R
N��}��:�Y:�ɇ5��qߘogg�]�}���u���k�ј�8i ����ۇF�u��l�iJB��-F@F��џw�Dx4�����:2T*��l�IXS���B���0��b�,�X>���@~�7�����'"%�?o����βQ�Ĩ{�>��R�`V���p:���m}?_�jh䝭�s�P/k���XgJ��Em��J�٥�Y��5��6�H���%?^�G�`ۻ1�ȥ<�p�����?I7�A�)e������dxi֓�BMBE�.��~����@�����J�k���~��[�>�k���5����O�]��^|,|+
�����I�+%ed����ܜC ��+7����Q���$���/Ov�bnݽ=��v\���@Y�h�������?�����?�>J�<��l:=H)-?y��9�BҐ�����*s� �6&gT[]tK��
fO�o�� �g��g�J���&hƙ�Fj��+���ہRq
��x�u��0���ß��ۇ:2�T�g�}��P:%`Q�
�\�_n){�x/v�(����z��"i��q�|4;����m�1�f���:�f���:�Yђ��W\�^��ɈPIRo9_�WL=vb���i�|�@�"%�����:��T��Y]s�}�8	��tz0&�0�1\PdD#�u?} '��=.|��|��<H��t�v����`V�����
��J�G�ﾟ>퓑����������>A��P����gP�IXw�?f_�irۚsp����k��R
Aau��w2a�U߽���A@߿���$��\�5��xH)�o߾�8��V�v%�|���p�o��բ���}��Ԏz� ��\'=~��g*͓��l�l|i|cz�ؓޛ�;�xV����ܹX����
�A4���w�˥{H]d�O���5^O�znG�j8�W���zd|������[G��%T��b��T����BT�e�
v�n���<�;4���|�}�OR�����x2.U�Ew�{�rzT���p�>#��'��F���+�A}��  �^_�B��<���L�gL��佮յ���=�|�d�b��"��c{w�/�zEqǅd݉���D`��uu��U�4�H�܇}���p7��)4A�b41��Md���2�в��;�pxh�:��Y�盢�.N�߰gv�n���We����j���>�����ýWIb4���^��oa��į��~��۸R�]�~�0���giƹ�i/�{<󽻳W�T�˩�������#`�����;7�~N���&����9��8�l�dQ�H�h�3[q3����MT���՝�\ث:&�*��쨎�e{ۛ��W��xm'tx<���{{=�v�G���]�=�onL�$��[�b��M��ZF^��*�==d�<���X�{@��)[�ʒ��N�Q�ʇ�P�Th�凮��d�NL&P{[+\بR���:�A�S�z���h��]>�� d�5z����g4H��n�����"kp�8sxS��<�jz_)���ç^j�:=]p�3&U{f]��b�S8��S'C:���&������lxn��&ˮ7����2�Ŋ6�Z�ZU��)iS��U�Kl�6%��FZ�!�!h�*�h�hQ+��Z���*Tk
�cq��E̪cj����p�j�hե�-�Z���m�؋mm���n\1ZR��TJ㖍�J�j�\Dk,T�F��p�Z�Q��V��P���R�TK\0̵���t�������p0J��6������h��Q�alTQ���Yr� �Kˊ�b&f��4
��h�j9�f[T��6�6�U���)l��3m-��Um.���kj�TeT��f!������e�Eb�b��Fڬ�V��Ɋ�b�lr���&Z")�Z
�#mJQCICVhUI�Q�4��30j��\�Z5�eE+m���)i��.���V�2ТZ6�B��Q(�֩1��1���n&`�4ml+4��_s� 8;� o�8C{�˚�b"�5�#�#m�V��Qjj֖W-��(�Y+,kTe�a�����U5��آ�j�U�9dr�+�N9PQ��*�JURʈ��G�C)���#+�.n���@�^��t0�Ce�&��;<�u=#c]�䑑n�FY9oq�tu����:[��wݤ��Y1��pr��c�wUn7U�{�ǝ�^�\/=F�v���R���qnyD���-��M7B ���z�n��6�v�9rq�ڃc�4,l�� �C�[�u��x�e�
� .�xyy1ϛ� NqWՃ����ͥg��{`���Ē�. �U띛N�뵸���4k�8zk��۱^sV$�<�lv.�Qݳ�woHs���❖�ۮ��3�`�L>��if�r
���θ���q��j�1�u�[�m�^�q����q�nvU1n&n���1�5,���ny�h��\=a�����:9��� ��A�=��:J��}yb!�;3�iݹ��Ir�<�\�3���n��s�<=V�Ѳ�k�wHc����dAup�ɍ��ۺ_kn uk%�}���n<Jz�6=�ؽ���s ����"v�76۬��iA��t+�Daݥ����q�9w4���=��un��J��x�p�����
v�w[l�cGmz���Wšjy�-�*ŎxM��M���Us��Ik��O=�z�6�1�C����Z�D�_4f�t�<�3�<���鳍�>h�T^�Qcn�ۮ�V��Wj�n���ˣ7c�w����x܌����5=���l+���҅mm�wB9PD�m��rz�����]絗���Dc���r�v,�5s��#�u�ַn����m�$m�d9q�qn��s�	v�	P1��+ۛ�nzx66^�*vIǶ�[)of�+�a�m����m1�=t=���R<on������:�Z�+�{mӓr������٧:����t�p�Ϻ��.��n��W���6 �<N������m���ٓ�p�݋n�hM5l����m6�7
��wl��I�.80{F�胱۷.�n�0nݞn˥�<T.�Γ;b�����
g3��4ql̚���b+���{eѿ�w����r���㫮ɴ�}Q�Q�̝kn�ΰ9�=��/l�AEuˎ:1������YW��s�0v������b�1z����뙭��;�L!�uf�rV��^N@��z�۬og�b�닶6�i�c�-n��Ӱ6�pÁ�.��n�\�J˗j`��ۭջn��nh.��ۣ��p��_/�����Q��ۚ�6}wc7o�9ں��7f'��8����I6�n �"0W�����<Ñ��g[]�tw������u�:1�k_�O�'�y�6u:�YY++%u�w���8$�Q%aa�����0�>��xzw=��$�;�߾�ԝB�Q�����;���i����	�3U�xu ����퇑�AHg�m��r�~����H�C�$<@ ��;��bAN�3}���td��� |郌8Y,b����Q�G��\�{���0�殹��º�~�a�0�J!RX!Xf���:3���*y�__}�M��߇�D��Z���ہ��H[a�����to�`Dp�%^�7�H�>x,����{�g̕�d�|�<��M!D�
$�)���9��
�RT��{�ő�w�i�^�L� ��H�&*6���C@�w���]TsY���D�;���ñ��!m=��s�H\�W�]~s>�~~=!^�+�����*T
�&o�������T(�~�߶u�<��	����������8z��G(��N;�yx�v�bOk�Wk9�9��?����ϰ�ѣ-��>��>a_<�sp1 ���o����:�FT
%@�����@B>��P��Ɵ��j8��M�}�����f���ïX�|�}�7X�5sZ�N	;������
����oG�#�����r�����Q�f��x�}F�|n,v�(���>Tq1n�n�[}@kz�'l��(��f�|k���y+r��  Iǜ�^��d�(��RV���0�
*J����u'D+%Y5�~}{��?~�>~:�@n|-[)�D8h�B��'�gVH<��-?y��9Ґ�R��[�������9��*AN VQ3��p�:2VQ��D3�����tIX\�b{͈H����^|+�>��� �����~��s�q'�*K�9���γ��e@�P.~�߸u�XjAu�_����:f��x����r|,�>b���F��S�(�}�'�ed��%u�u������|����~&��$�/?{�y�aRT��}�Τ�!Y(ʐ]{�}�8	��U�LY�g$N�\��E�J�cͩ��S�]0dgts�/�$�n�=g�OF�O3�����s��W5�.:ύ |����϶z���
K@Ͻ���!R`������H����(�v G�����g�}*A@�~��C�J��}<��+�5m�Y�u�F��뛁R
Ns�>���y���x���w�3��@����è��������R
Aەپ��G1�Y�}>l �N���h�b�k�18�����:�@�����W~w_nC�*A`�g��ߍ�}�������-N}���*�(���w�ot�	�������mׯSJ5�|��s����Z��*X��u]TsyR*�)���x�gY�3�������7� �5��<a�°�
��g�l�Ad�ed������8�@���ot�hL�j�c���̯�@����o�c���#���I 7鿶s����k�~����q�P��O�� ��o�gL�}dR�x,滾nN�_6~����f\�����	��|�ΑDx5YC�S�˽HJ�{����R�R�{��p� Ґ�3�}��Ǭ
��i�ﾷ2�������^�>�>��Kt^�D�Ϸ�����:�ˣ�LBb	�a����B��q '�͜H,��������G#'
IXS=��rH,9�ߺ8�����?C�*y���Τ����VW^��@����UW5�.:͚@�������`Q���u���_?������ii
�i�{��q �+,L��}�u�dG���Dw���t�
���@�<���ts�[BJ���`�#�]?$AI�+�>�p�'FT
%@�������N�v	Xk�u�>���a�s�=`U��_e0ю�Ն��A \�}"���'�ǒ�r���I�w���N$�����}�u�c
�ID�|��H�ٷ�}���>ֳ_�*f��C=�Cۋ��3X�WR��X��~XR�6���vף҇��}1���ݓqw���Ż�nn������y�������?�?���5��8	�����t�&k5G1���a������HR�3�Ͼ�ă�u�߳9�{��t�:�Zk�߼�S�*eL����u ��%@�|��C�J�yo~�1��L�!��Ȇ�"8960vwE�[tX#mKϝhB�β�8k����������&��g���
�}��T�!RQ
�<���βQ� �\��~������͎{�]Sx�
��I�+�>�p�с^��]2�kY�̻���I�s���u����w���Zs���6�矷�
�T�}�<�:ì+
¤�3�=�gRu
�YY>����}<��w�ٟ{�B ��Z�\�h��8i ��߻�!D���H�x"<	^>=��o�߳���9� ���&y�~�:Ό��*C=�߶uĕ�u���X:ѡ	D�G���G>��zN��֧�y����y�6��*Aa�߹ݝ�J2�T��Ͼ���VjAu�>��s����8A�!m�~�>�:�`V�_p|��.:3W5�@������l�t@����d������2T<���Ǿ{���}�>C�%as]�XtV0�*g�>�gR'YY,eu�>��(���}��F���_E�F�株��]�7�m�S'`�U5n��2#b�7��#=����g�6�LԟmR{�JaWV�^�HBI��k�����f��X3(��������hc��G�f���nG�<f�m��볹y��á�ݏf�s�ln���F�i��c�gYE��n노N�iĞ�WX��/#�'s�a칑Mgc���Gmѭ���񄋋�r�ְ
w=hּ�=[0�n�+s�h#=�{d��e���Π�/^i,��^��s^v�V�U�d�j�c�n�`y�Aٺ�Fr�ջkWn �ۯ;v�7�C��j��\z%������_��nl��������o�<�v=`V��Ͼ���B�B��k�}�@S� �����~����huWl�YΌ�>�߶q��9�����]Z�&�Z��i����?0�*&�����߃���9�q �x	P.{��p�A`t��]yϷ���JB����Iu��<	�3�@P,1#��|��3�}ݝN�VVJ�]}�w��%B�*Aakc��}�<9���aĂà¤�g���ΤN��VW^s��ND�*���IN�(2 �B>���ow���VjA@����-��k���w�
q�@��g����Ͼ����=U���Y�� Vg�"��'��Ԝ�p��J ��#�������IA
�;Ͻ��3����߼�a�m�����k�~�g:��F�+W��|B!���}_}>l�U������_�������b���C0�<¨�t�����n�5�5�:��������ݿ�ڻ:�k��D����l�u����k�1
$��}Ͼ�8ñ�a�;���u��� ]~���$���eH.���
�����:f�&]i2����a��l�fπ@�<7qw؅�ى_I�'>�y$O�m�W������	_��I�$u9�Pj���+�u������Q�Vmz�reU��v���l�MX����~��� _�;�<�g?�B�B��[����@�ȁR��3�}�u����d�:�V7�r�;�S#��'��]Rw��)�Y�g!�a\��}���Q
��V�<�gY�JʁD��9�����~�~��ȕ �_s^�H)��}�q�0+gtw�.��j�Yr�S�L��wgQ��~�u�:ϣ%H/��\����J�X\�y�u�c
�P3�=�gw]�3�K��N���;��'"b���t�sYta��I�~���x=`Xԅ-?{��9�B�=׏ޟ3������*q�+*g�����u���T*������'���]�U��� ��)z0�%/�`��N��e��pn��Gm&E#nݵtw����~�h�Y�Y�8��}���À�T*J!Xgy�:3��e@�P.}�p�<	���h����ϴ��d��̤�e��}�Ǒ�W^�}*�C����kp18$�=��:�@�����_��\�}=�I��>��H�y��6Ã
°�*g�{�Τ���>ϖ=�go���S�}� !h*�F�L��e�èJ���A��Z����y��9�B�HV�
�߾珿0j^u	���s؟L��I��QӥVn;4xnү�ǽ($yr��g�ڙ=��f�&4H^��u��-����$e��{6��H�}��� T��>��jg#%H(T3���u�+
s�I�4[(�چ�xI�|��� ޏ��_���w���AI�
�^~�Gq���PJ�fy����D�
5�Z�m}>���R�خ�	���O�&��_ܘ(��m�U�,�#������ VQ���WW�{��&����7�:M!�$�.s�ۇpaXV;�l�N�R%�����p4���q���v��G��,A0be�B�����l�l
)����X��w<�e .��������eц�Ɛ>J�o����jB�@����9Ґ�����y� i8�H�꿗�\�V q�3'_�Q���d�PC>��vu ���6��k3V�Y���C�:0���y����T��y����p�랇�>�����:ʁR�S>���:�XjAu}�ہɺA���ˣ�Ǧ�����
_|�8�������L,tc�ֹ�N������
��R��>���hQ%B�J��wO�חG����x���aRT�|�ݝI�+%ed�����n�9�����`�u��
�����W����e(�����ԅ@�<�vs�!m!Z�����p4�� ��o߾�8�~��?��<�ڷ�q툣s���{�i˲��&/gq8��j�����FM����>XH��9OwUi����z9����)����s�C�{�˭f���w�@?���ђ�D��H�<	�_T���lbnxm��r��ہ��B��V�������M��>Cm4�@
+��@u+�`X5�����
A�����F���e˄v&DDߎA�� �7c���ۣə�1�"�୸�l��,M�۲Խ��;y0P14�N>�G�z2��N�T���]]���FM�bJ�IO���|(�W��>X��أ^�FF�2N���~�gRtB�VVJ2������6�K͟y��0sNh�W��8�����
4|(��
rW�\���s�o�{��R ��Zk7��@�p@�P+*k߾�8�2VPd�}�����׭�no�G�>,�s�CD8�0�0��Ϲ���i(�ID+w�X�}G�@�!U_z�ߺs�v��?%`Q��ߟn�)K�|�(��"����CL(.p�x"����E�7��S�>��"<	�׼���hQ%B��)�>�p�0�+
��y��8�������7��'VJ2���w'"m����5�9�%�vq�X~�j`pjB�}��l�A����o\�AH/�s���N T�a��}�m����d�T3�=�gP,<��R��ê>l�(UT��5p!\����=x\?�vX�U��3;n���;���j��VHI�Io�o�l�{���θ��패��x��e(m�^�3��	���U͸/c�nTIۮ��:98��L����h���F��;kf��y����w���tS�:�W����i;]�1)���-�9��Z�;���u���]�X�v����N�*À�Y7l��7:��1��J�e��^�t�ۧ��lM�.�;���_nntpk�,6��6v{'k��3���83�c�7f��½Mc��	qN�"�l�^���Hݺv�]N��r��q��Ӌ�|���3N���!��¹}��m ��
�_~�P�'#* ������dx�ϲ�آH�N6��w��&���k�y�q���ts�5�W15r��7�ؓ>���Ԁ��O�����E�p���K/$Pޒ	*%a�>�P�+
¤�g�w�,�_���������wm�tv��������6�e��}�fb9���W��{�u�?5!m;�l�iB���k������Ϸ�$�Ή���P�8�R
��~�Ԃçy������N8�#����d���x���럷����
LB��Vw|���d�� �g�y�� v%`V�+]o=�p���Z\�mf��K����Q��^O��CL(jp�x"����E��
�YY+��l�2isϏ>��w��=��Ci+��5�aRTϽ�ݝH,�ed����߷'���Y������q�����On�v�:8�ݎ�c��㇠J8�?x?��'��n���𕇜��0(ԅ-=��s���!Ru�{� br T��~����@��A3}�q����2T�����u%ag?so�U�6�����Ci������H�o�}��_	>�b�i��ȼ"��];�}��[:}W�/,ƯF�`f���t�F,�3"6MȘz'^^��ȋ.��K)#q���nC��Xo�����J�����p�A`tk�w���p9�A����>���Xp����4|+�X���B;�WY�Nę�>�ΧD
�2VQ���}��2i
$�Q%a�~�~��]{�^w���{�q�aF%L����N�VJʅ�{����֏|�\�9��U��>�zk��V�k�D�U� A��uH�$�����/w�UK7�4C�(qT��"$x�v��Ooj���{tp�j����H��4crЬ*���g1���&��{Rq<-����f϶�ە4�fs��p�������\�8mwWVUH-���wsg/Pˎ����"jVt�Q$���S[�,�� �l�MU��Ht*���G���}<	�ڼS�A1�� -RQ{�,��m�	��'e��FHD�lZQ� ��}2I�]�����t":T��� ]�Ғc'��D�}�y�z����l���6ޏ* ���f����S�����Y�/i�H�, z�ZY�\ϓ�����+NT�J �������|��r�����C����3X�X���tM̗�D���vr>@B_��jX�{(���}<���ކ�.�>L6���Nݾ��X�=�i�`�<c�ˡܽ�e�+�7*U��qk5l麗���ԡ��]��;劶�l����7*��m�RqVz�J�Ԃ0Ļ����|����E}�./h�^���{�]V�E���2Wz1����Ct�
4��b0ot	L(.�#�^Im�0��4����7�\=�og��P7U�]�<�]�=������ي�]������ԗ�lҞj\��57��sȯh�<�C8�
�"�ۻ����� ����{��<w���o�:n��j�V��s��&ݛIѼ߼,agap�+��l�N+�����c.��O�����7���������`!6���`X��z鶪J}r�ˁğ+���L�g��/w�O[����5�4��� �������"�j�o�!]孝����o2�}WT�Y`�Q�f<�;EW������j����Wj�ڦ�����;!�7���o��xoZ;f�r��gon<`��oH9�����ݹ���9O�NdL���<Z��s�ު��ٷf���ˑ��؉�ws��o����}��o{�{�Ӎw��˞��z\s�P��<�'Nx���,�%A( �8 ��Q������)bJZT�TV���2�d��(ҵ��a�f#��Q*UEY�a�WI��頊��c��Ym�bڣm�b���H��u�&#���X��]P��A���H�iE��E)lT�T*���qD���X30��QE��ab�q�p�.Z�Z1Dq�(����B�����k���J[*5�m�X�ڥ,B�ԭ����U�J�Q�LEDT�m���(,�J�m�6�EQb(e�2��b\�j*�J����rҶ��*��R�2�
��[�b��%�URM����o5�b�,P�Q�\�1*�j���Ed��#m��,X�Md�,+VڈV�,0J�Į0�-��,T[V�m,VТ"V�������������H�)Sb��]�YF4������mX�D̤F&Yb�7s*Ԥ��m���T`�ֱ�f6؃����.[YDUQZ[J+_�@�g~��oc�@�#�D��bB �2�P]=U�y��D�W1���fH�B�ީ��Ż���mTd�AlZ�DB0�I�Ӑ\wO��AU��F�}񇻾�>ڜ|dgc�
�ޯv�3Umds0�R{�:.ɍ�y�by2��qsE�ѴWk�@�%6�pQ}���ˈb1o�"eH1ײ���ު�=V/OF�u������o\�|\�')���&�sꝮ�@���s��D8z�&*��$���A�n��;P��8;�w>G�YADx�l�MU{Y I�����H1��U���6�H�Lvd�'�7z�K�Y��у���:��� ��>!VgH����+x�����M���A��^Ǖ�{�N�OM��s�]�rUq�w;]}����v�~�Y�\�y�y�d�!M\Лb��y�Z������^̂F���h���	��U�I2�4����XyKv�U�uP ����M�(vЎ��,�&"/�5Y[=����g�ז�4�g��=��<�OF�Nf+4��B��������� [y�^$�����y苮��і{)߉��`�c�xYi<E������e�v�+%L�Q�$����j� {|���j����Is���1�M6����>$��҉f���W{����:� �+�گL=����n��ʈ� �Z�wҼ=I�7ן� =��� &="Losa�p.��̞۪$M��Ј�у���U����oi����$���q}�(��d I�ot�1���N!�ߦH�	���[F�4��s���϶	V�E�P�s���`��+���r��x��O��]k�r�K�w�M@��A�S�����NQQ�[M�ZV���M�2͖y��,��Fq�Q!�q��W
	�<j�#��݇>ܫ�����`�e�]��X��nr���|��Д�����5��ph�O1tdސz�v���9'���{]���ؒ���4vs��Ӻ���#i��ٶ'�us\���U��9=�ɷ;���u�U�d���62�˶NӞ�nqv ���*�m��8N�ۛћJ�l�0*1�p[��۷F������;k]���1�p[�BAD4��NUP$�a�l�"I GwL���#�
���@�wdĝQ�P�	0Zr\w1W*�L��LE�;˞$a�i�ot�,s�.�0�zo�l]H}�(I�	�P7;du��&h����])���v��� �cO�F�L���p`7��T�ufq�cu�q��3`�!H�͙�$����5���Fk�����T�Q�p���ok$I���4�.����[S���y�3�A FvL�I[��F�^p�E�tC�1tވ~q�	�bF���fz^t]�YM�u÷u^�WYs-�����߲�$fi���[��Ay��	��꣯�����b�\�I��"�q�6ʈ�	���TI����]=��o���g�w|��-=�͉͘�rГ�̀���sIx�k����FA����Ͻ��|�c���lvC������� <=y7���̂A!vo�D�u��{W��C���6�|�DR`���$Unt�$�s��i����ω$-��MHw�(M�HDCT-�s�蝸��6��#� �j�VVuW�$�Y���Ğy�tG��UȠf�������L6�&�� �Lߵf���Ku���uU<Unt�$�oH��L�s�����qKa�sŇ�bH���Y�n{[�ۃi��kk��=b��������tki������IU��D�H��|k'A3 ���t9v��РUf����(E��Zi�Z} A1�sW���UZ2�{(
��$5�0	�ۊ��=��/�#9�6�D
*��z��>�k�`�I���쉮���\V_L�n��g&��|D\�ºc���Ì������d������P�z�I�o��
�%�5N� x�q����|����ď�o��K	���L���q���u1��C�;"� �qڤ�b���J�U��`�7��+մ%F	6�E�5U�r�dA��͓O+vu��rI*g��	$^Lb��h�F�]��T�n�/;���L��{�{9q���.3���x��$v;-�k�gKrZ�����ֹz��o��W]U�|I���	 ���
3^��$�;�`=u	�}��(b8�8��v�
�ȉ����sS@�A��@$�E�u
�|£Of3�'@$Nt�+D<H�Yopk�@O���L���L�徭� S��@���D����x q�X�PV��x��07Ѳ�'���mQ$����X�����U�����6�PF��������Vv�]��Z��j^'����W�^mHݻ��jDLY���Ò��ͽ���{��>�UR�����,��i�-��TI*w� ܮ��q��6��z���D_oP�HS��^"�d��{�[Qn _n�⭭��n��mٖ�Ąٺt���97n=��6��!I���G�2��T(��㲺f":���$�9�CY��Y�E���_H� W��'�f��x�6Z��ܓ�t�3l��k,:j�t�$�o;���Y�B�{�l��Mlk�[R�*����a��Qܮڣ�J�ޚ$T=q��[���&,�c��I>U��^$Nm�*����NņB�g���#&{+�I$*���L5�#�M�O�����\��4�I�QT�z�W�#���rg�6�V��J�ۡ@�*��H$kzb�'�L�x��++2�D��Gz��l�a������#̮�}�j��:-WT0ÃC+�ƃ��8_p�l�}��"L���_�o�^T�]�M��a�S� ��6��T�h����h�&a��`��ss9����<o�,��k�����Nm���l��и��q�y�\mc�݀����g�k[����:|���@6ݝ�GOv�����݋n��\pŸ�:��s��׭��4g�6�=�^#M&�m���jn'\���`c�����S�4�<��6�w]�^�}�s� �1�\e.6��۝�g��B�0!��wx��ٜƨ4�e3�yb���L��Yw�қ�v�Ž�훅 .�����?�ZD��O��s@�Unt�$�7���s[Oa�����$ �3��~�t��,$�	(MU��0Ap(����+��b� �W�TI&ޟ@%�����*�Mh3JTq,�Np�+j���Y� �/)��k��;��H$.��R���5�"�a�NqTw+��P1=Ӥ�	񘫩�O�S�A��]��[�䎟�jY2?��(��ee���`�A���P�Z1��x���T	�%J�^�o{��s۸������E�Bl����x�`�Y�Z����\]���.�sf�^�*�������&�!@iEpN窉$+vDO���d����K�J�*}�@�IR��	�܃�M�-90�z���OG�a��ۿvn y�~�U�I-T�{N��J�x�T
��\�t�"��_ܞ���F�{�\��8��E,��S`l��%޳�z�j#���<FUO�O����6����>;�p�����on�$z����Cj�ⅵ� �F��U��hw�:ap�����'�J�^��� �Q*4�X���u��9��V�Z�H1�zD���Y{���WB�͗Q��SRo5�"�a�I��<��>'�e�Mx�I��8�L�m)$�Ot� �,������W�~=�P�i�Ÿ�u���ۊ�g���7g�Zsss��ɜ�Y�������aHCZ+�cS�'ƺs���+/z�FҮ�qOol�FI1k�`�y�TO�X]a%B0QTު�ў���]-Ɲp�	��ڢIY{�^$��S/GNȪ���fT<�bz��M�-9 ��ڢH+o:EA�S�o��L������u+�1ү8bP�簠1;�"�p�F�U
xS����toF�Ke�M�:%�7�݀e��4���� 	ͽC����AY{�Q��+���&�%�ѹ]1�:m�{V� �����A!m�UA�;���.n�u]P'�Q*4�XP[Np�*zF�s��b�R�����>$����W�6��{��5�˹�[������;X��\�q��{\��&z�
��������gs<���~ev�J��@�!N�O�4!�ʌɥC���}UD-��]��%D&�"�M�n:,+�ʶˇ���	�*�:�Ē`���|S5�*�X����4���	(b �i:�������`�l�I9������fV������T	�w�2m`n!�[!&NA���l�=5�:B� �y�@��aOdO�7�J�t�M�5\9��ҫ�4ܨ��q�yndt��7�����${>�j�bl��	C{�U�SDYLm���"�RNR�[3�� x�/���U�Tih�0҅��96���?v�Y�-U��x;)u��<���=����;�Mb�Ӳ����cV�\�v�l��/c\��7<f�y����^�$ujF Ǒ���8�XPYn�}�묪� �sd3����p��>�|w��Aˬ�P0gr|Ϫ5h�`���n��� �]{{k\���O��S�#����P�r&�h����SC^m	p��MBE������I�gU!i8#��_tV�$3�I����@Z�n('4��P�|ef����ˉ$��٢I/z�S��®���+؛��^,�L��1U����l��-0�ߨV�t��+3�E��:4R{P'����
�ޚ/ϳ��/hrǉ*�v�TV�����sQ�Ӎ�HaG\$g�~$�g��C-�`׎z��[sݰz�[�}֝`�;=�.vr��}���wr���I�u�U���Yyͯ�猞r�g�F�tz ��r箰d�8ɻ>;+�mN~�ߒ��w@xr3�b���墖�Y���ܳ��ӂ�n�L�E占�����AɍŲ�;�B�S'<]�-��"�;=\�7��ޚ��Tnd��W��]9-=fu��8���a>>i�ft��&���ҝ�g���ঃu�m(�o{�mi��F����=Юh:�y�2G�wy��G'�V���t�n1��d����ۧ��X	˹���n��4�<��.X�G��Q2��&���׬i�v'�p�5nzg�Ol�
�J�Itd{�����N���{Z���4�[Ԡ�O"���PoS���f��3ǌ���g����ˁ�Rq-�D}p�BS�#����*R�����d���弮+`������>�`�c�t�4�`�f&a�.�f�����<.IS�'ρ��D<��Қ��Kr.f	��1:{$�*�z4<致;��9]���1h��?.~B�>����w�z�=OXp�����6W.�귶7b�n�hKP������L��.j�v.���W7Vm�WT/�OS��>߳��?�ʹ�G�3�{v��j���=���=�}�B�\�8�LB/%�Y�Q�eݕ\�N�}�P<߻����M���S�[��j���TU-�h���UTX��5YFҪȵ�"�)iEi[5IUʶ��X�(��U�b�h���J]aE-D[j�-�-v����U���-t�����P`��f-��1R�[E�m�i.[�qm�
��KX�-�5v�Q��)h֕��J ����s6�b&�[j���X.e-��Qb(�[V�+cZ.���b*(��X��h�"Zj6���b��Yh�Uem�ƍۉ�t��EQ���lZ�����1L-m��ەa�j�V�ڴ�V+-DR����T�16V����T(�W֚&5K�fj�n+R�kV��Z�Q����8ܴF�[��7���Դ��-�R�+��pՆ�V�j�J��2��kJQ���iJ��[�DZ��8.�em���P�aAƕ-J��E-q*GZ��c��n��Y�n��'c��G:{O9���������K˚�����])����'�Ƭ�g��y�f�x�v��p޷>�Bo-Ҳ'j݆����]�7Vq`��r^�Kq9����Nr	��t�����ۻq=���T���g/6ƒ�Z^�r5�[vq��U93vq��:ULi70Ϟ{n�8���u��=�!Ε�j�^-t�W'm�Vҏ;�jx���n{ ��әw���.즃v��i�-۲�
,ѡ���׷\;�ꇊ1Y��jP-�ҋ��w�f�[l:��c��zٷgp��mݜ�ƅ�]�Sd�����-����\��̜��]�;Q�.K#m�bݦ^�p�H�{���x瓶�4p��t��z^8�<G��=u�X�u�� ��1CL�'�nS5%�N�<8��L.�%�l��x;kOC<���6�]V�2�4�7����]��m���ه��t���go�:�v6��R)�႘.�ӘcpM��Ѫ�n&�V:jҝ�7pr!ۣI�Ãiɮ�eގ�mۻ{&n瀥6�kV���݁�t��ud�dѸ6d���v$�R�+76���s���۶�:��ヮD����=���m�f��yy�۶y���.{�[�����Җ���e�8`O/V�YB�"P0��B)6C���0���N,��'g�O9�7ˏ�5���vw	ڡ5�زu��s���|�Y/E�nP��%Hۇ����]en7�se��[�g#nx���F�msp�kX�'�q�n
\�z��xܗGv����v������+O=�N^���;��Z�M�n��z�����ѝF�v5�ۮ�t�\ݓxc�7:oC�z�:�0�TD�t�4�yl�{N�t�ڻp\���psF��R�Y�q�sa�{Nޭ�l��Ύ��N^9��>5��m����z�nz7<�U�c���=�<�0Wn�7�p�B\�Ǡ�ל��zS��� �^���@���>:C�չ������S��W�Z �j�7Yw	�՞�P�J�P湌Vɫnh��-�{�sB:�Ӭ�Z��ME�Í#ܻ��y�ʜwM��F�݃�GS��=<sŌ��튻u��ny��n��@�ٽc.9�.�`�燳n8�mR��ZS�bU�	��<u�ϖ����b5��8�g<c�@wf�"��f��g ;E�;�K�m�5�{;{\�E�.\�v��g�h�_'�ϝ�q�C��9xfm��y�7�ymrÁht�O=i78, �箜��:��+�Al�U�����}�F�D(4Yv�I:ﺅ	�>Y{�^�'X.���(������@��Z�A�	��8�[]S���}��Gp�dh'Ɲ�H�V_uQ �ܣ5�wH�1����̓m�6 &Kt;'�t�
�ޚ>���1�z�hݞ�����A+/����dK�TBj,���m�e�i��lI��{�� ����������W��8��tA9Ϫ�&W@GBn(':��P�Q��w5+s3�|��>YUB�
�:�H(����*;Ǥ�|�$���n(�F�8m�X�,\�vxcbG��6-ʔg!�I.���n��2�d$�i��:��D��sf���;� в�룘�$�ΐ���H˜��<i+���2ϋ��B{��P�����w:�r��q<7��J쳊޾{���ޫ�Cp�z�L5g�w�ɷ�	���Eg#���ɓ嬫�?�{շӟP%wgH���X&fECG�]{�TS�H��X�A�0�pC���A(�t��	Fi������|(���B�H(��M�ll(!�2[�;��x��y[�.���u4I%9�$��wt�r9kT#/I��
���J!5	Zn|Q��Evu
�xQ�΋�D�l�W����	[�U���]���f����4�����	J�v.ĺ@5�GOV޸�R�]�k��yq�\��������E@i=���eQ���$�LV�P�u�����9�ʠ|��Hb:�2�-��� �=TOF��{�5D��N���	]�P��w�O��.q�{~3X.#Aa�L�(&��=2�${�T|I�-��:���}�8���:���)-�wœ�u�l�/o|̙b��z����������CV�吝ԕ�f�����%T�P���=���9��x�g~��G����)k8&n�s[�t��q���;�I6�6��HY������|z�'� � ����u\[Ć7�<n@�j�!f�M�
*���{Z	j�bI���x�Y��@�8�n2�L=����sG�݆�nx;s����g9�/\�m]ֆ�>��˝b��R������ M*��e���٠I+'����[����؛������{�U�qet"4&�B��sI��Q$nM�Q7S]w�H�z$6�z�WuQ$��Z���-��;Y�FՆ\3�`��C}`Q���5�	���:�Y�5��TIY]�ј���8P`8��t�l�-
�5Ѕ�{_t�$���TA*U�ݲ���48!�|շ�(����\�ܗ'�DX߱��]���ۇm�R�}��}��)a㷅�sv��{"�`I��5�Q���������}�U�)k&i�C�__�B��R�鈡�ct��ݽʢIY[�D*�Ds���&
��e�p�p�d�Lޛ�tY�nƖ۳�]�8�E�uչ���z{��������� 0��}��J�ޚJ��AgzOq����9d+ɪ��$�m��
��ň) "���/�@7��;c;lQe]S�y� @^Ŭ`|��	$���#	���}��m%&=�J�*)o◫��� *���@{���f6�U�;�� {+��$���9�@.�B�JjR��@���.}�H�\V����5��� ��*��t� �vvfȽ�۱�}��/ͫ�q𺭉P�5
���kp� s�y���^���ek+� ^��ˀ *�k��^ܮ�	W�K�ݨt�,����/���n=bpj�I<��(#�{F����',�,��a^�"��
t<�͸ɕk����=�g�J^���h�ZP�E��p�{�"�[=v��cm���h�	��#�h1���4���X� ��wa�t�k)�Y:y��c���y˦v��q�Pl�p�ڲ:=�
}s��c�uq�ݵ�����jn��t��ٻ>ф���F��<7��cv.úv{ u��t��W[�fJ��q���g<��7t����ǣ�l')�u��m�m��50a�F�vv�����C�;^�D�2v��Ųt=�h�ϿC��`Q55JV��cW��	�*�u� �}ٙ�m��}��������Y��"5�Z� @a�t��6�ZA"�k�Ȟ=>#��w��  }WY��\�s�������j��N�r���$Wl+��S$y�<��ϳ�9=�}Kzo� )L��ݻ��N�_��	cE�0������ �5������0	��+�x�T��ֻ�0�y'�	�R��$R�R��@�ؕ�f}5��o�3�|�ϸQ�bU��9�8 �׽��F79�%�|��kg��a'2����l��؞��k$�v���%���b���8�t��UXj����WD�E
���U�Y͵2s�y�`@��r���Zo;غ�=��7sk���Bn�\�0��È��+�U�\2����rذn 5���꿸K�c����&��^��ٌ˕��j�d�t�g��^���d��,(a��3X����fc>�B�I%�_}vg ��ܛ	��A�ӝ;ʯ�"����C�1˥ݹ�~��^J79\�	�w�}�εko���ݙ�@o�6�uň$N��Yuһ�R�L���[������J3:h�Iy$�r:�5� ��l�	7�ݙ�u�Q_l	Q5P�R�AKy7� @U�k�V{sj~\���U��f@ D����'�~�n�s"c=~�G������82h�v����˝77��`W]{c=V���nn�q�����a�v."���W���d�+��� @W��p����>����w��2 �
�jl��u_`x�-4�'����'~;��P�&�Y �$�W�� 	8V��	uY*�U�}|�n�X�0�m6Êv��bs,
�W8t@�"U{q��'yx�D���r��z���U������mЭ�������6t^�=y�s�kp$����B=W��"^Л���y[�� �{w� ���ߓa'�~���D�z��T�1���[ۛq΋[9��Q)-s�L��"�׬p&vwf3w�oU	{���6�qb*��d����I�/��B3���wd�u96�	%Q������]�U7/Nc�.ӑ4�lU�����h�\=V��h����C.�੶0�e���#"��L�(wΉ2µֿ�L�����ɾk/��H�b���7�	 �j6�Ќ�`��eC �	�4s�tm)O�dfE��e��> �"+�sf�vf@L��s%��W�{	?�8�U�BA��c*@��vL����@v"�����]ٔI$���D璽��Jn�.d�d��in���^p�7Cty��T��f^�st}��{�{3  ��'Q�=�س~lef,g���Y�|;w�Ֆ���ˣvIP�=\zj��6�V��ۭˣ����=��$暅I�h�m7���G�� ����5	 vg�b���t��nmݤIF�9�N�Fg�j5��/n����k�2�7sy������&ÝI�
�任%TL¡��=�y�[�����1�)��=+�W�1ss�i���Jjgs�8R*T!	�D-�8t��瑁 @V�����p�����U���޽��I3#ڈn�P��[��� J~��U+��⠔C6���&�ns�	W˶�QY��:��0�T20�sI����I��٠!/$��
��S[���a�@ G{;�2  ��WY.#� 
�TET"����upB���n�m_�^�y$Wys^u�}��.lX
����'w���&i��)����D$b�D�W�|�K��+����'��q!Z�� !V/�
�>����N�}g<��-w�w۫��w���_��_���L�	���p��z�{os��Em�^��[�dbʉ����Ox5��uGM\5�.e�����r�ll����pc�ɑH�m�a��R��q�,���Q�t��ƭҽM۸^�A.�$m;���t"Z7[0l[��;���}!��@:iwQm۷[k2z��yLa�u�jı��Ez�<6������[l+��O��?�����NH�0r�R^px��6��Ԣ��ќ�Zv�q�w�Ռ�&��w��y�n:�f]�<�]nJ��۷��^;9�dܜq�:,qr�i�6\�~����뫮�����;7s0  ��u��� �k��=����sw3;���d ]���(�ŊH!
D*N��K+��9I�ɻ�*�7= ^��8ku�,4�]�������;ZvB��-�Kk��d�+]k��@`�T����7~ +�Z�Q33X��󦒩RR��P!7\�.):~��8������ ��c� ���fu{�f�;���_ gz���"5�^�
�TET"�ܦ�;��y��<ͯkԳ���f�y60 ��[��O���vfz��z�n)�ۯ:� �D#���n����p٧V9n��=�l��厭H���7"3=�t(�S)U$��������" ʍ�PJ�H^�u݄�5N컲f��^cC�]s&_�A^u��PD��H�P�a�7N��n��A()�_��'���{lf�����м�
�j��m(9�J�aї�E�N=3�u{t��CBRTr�mn�)�=/.�L�� ���e��@��c�&L��ݙ�@�=���s�s��j�����qb�B�Q
����ɖ��y���{��Ul�Φ���@ε��@#7�٘�Qu�e(��3J�P����Ws3�	�YZ� ��o &H+r��^Ԇ�Mu�$�S�T!��4�C �	
��o�# 
쭷YF�n�Gq�����`|���3�>��ܮ�cv�[����}���H�HE<Ic�t6�2x-�ے�	��N��vU8󋓵X�������t�U��{)��3��瑁�ո��8�Se3�n0ƽЮv:�I!}��d������eD�x+닪�$�Qn�%^��~u2�nwfd�nW7D�jo�ӝ��v׭�B3�UR��a�7L����i����BA$��ymq}��0ѿi����m��V��m�2���G�2X�G�Wd�?Q�6y�������ו$�gh��Ǭ�����c� �w�V��N�l��z�Ƿ�v�"��{��ؼ3 �"N��:&ډ�����׾�7s�n�"���lw��X���U�㲐���|yG�)������y�=�|tmQ��"�"�T��9�SzƔ�LB���C!Z֋7�}�W;��fҺǠ�˫3�k`��ZK˙KB�Y��v���jl��ұf_'���r8�;5w"eM��K��$ܷ���{�کtM�#���=����^O��IޞWs���"wg��;*�z+=��Q��<Sû��ys��7�����-�à��H���Z���0�H9k^������ۮ�:6?F�Eɤ���<���;l�ד��/��㮝��/l�r];���&��ۓZ�޹}��?]���� b@�7�k�����f]����Q���e�R,V��cKQ��,�".`f
�;�Z&�|��-��ܟ*i͚<���Yj���we�i����'���gOWO�{�J|�]�z�=�,�^�∸t��(�ժk��'|�U�G���uݭ�+�În<Xޛ��Q�J˺���9�� ��ݰy=v��
 �ڈ�s�w^y{:�ݭD>��mGg�;d�47�}n��*7n}�����4�=틮���׈Z�;t�{��n���>>ro��	�j�m�D�j ��HӢ�U��0�m�jK���S܄����{�x��u�,����>���z�*?�(��(Q�X�h�J�kT÷x�e�U��VR�F��bT�bV�Qr�"�R��,���+e�f�Z4ee�iQueDLq̨ʱc�0��\*��tܪ5j1ueM5m�([V�h�T�c�.�TEYmV�eiq*����;�f��U���V#
,cs+iUDa����k�Esy1�
���U�f8ڊ ������ޮkSy%MZ%�Kl�Z�頋J�Q[eZ���l�WN1��*���
���D�qDAb�*0LiZ&�;n�3v�Z�*al��2�X�"ҥ���sX�15J`��b ,R��h��
*��TՔ�j`�Keƪ�*��F�F�MfU��ZةmFڨ,Fņ�E��)sz4$PA5�[�2�R�)Qj.e�V���TQF��b�ZQ�kTTģi+TL���BOw������;�x V�sP,�IB6Ds.���t������^	/%��9�  Ev.c� ��w���/s�$�O�䷽���޲�h��*��R��� &k�k��K��f߯&�y{=�nk�̀�>+��������-�s�2��t2a��*E0{����q���sr����a�$�hN�t��9������)JbiA)9uw�� ��+l��V/��%f���Z�G�/[�p���W7A���t��M�ge;�@�x��N�yS\۞ +r��  +�~D�N�ft{���װ��a��NeURJJ�fvV7� �\�L�1썡#���� ���L���\#��QJ)EB��	4��v�<"��� z�n(" �>�k���ܾ빞��FqהWJ����x(�n']�+���5�p�
��H�x}��k��R�"�0��c��%5��ncjEۗ�C�4�4~��~�Iy}wU ��ň$�(UR����R��������
�n��7�̙~�@j�c�&PQ�T!䗷/���Zx͌ג`f��ݑc��/G#������S��3nn��ۭ�\r�;|���_��Zh������W:����w7�n�Tص�vp�{���D�}c�d���*&UP�% �u^\���81犴ib������X�1� }�����~t\�;��Գ�����"s{�Ш�1��2��{�Rd@{��Ӹ�I�hX���˴߀� �u�� �gvf@E��pd�%�Cl���+닢:����)y��@nofd�nW8#��v,�d����ބ���S��� 1�闹�[i����B�[��14XIZ���";;���>+r��u&۾��N�� �Mpy+���&��Z�0^n%��xw�hɴ��'��z������Zs�:��ˮer�.���_��'i��L^�Ө����X
>��!8�#��t��v�ي0vuxÎ��D��@�Y��<��}����cm��{m:]kn�v.�ܽAvd�ǋx<����I��q��[l;z.v����i:ݲ;��k�u���[�(����㧲�lsւ�k�L�*$�C��I�N0p60�{D�s��.���ͻY�q��q�i7c��<�6�0om�;v��nQ��l��u�wjzy�:�<��d����(�$6��u�+=�q�:��p3�~�{��B��B^���\������0 �>��̙��j66���&ȃ^W7D�Ϲ��"+޲�h�J��HR䭮�P@7x�1gV�� ��u��%䒍�tI�%[�cL,��َ3���O"�S��pjo�0 
��o���s�ڪ��` ;^�f@[��˷���L�TB��M�c�u<s��-u������y�%vm�^I�Q9Y:p���y%wywd�[�'�P*�UI))ۃ717 W��*.ԫ!+Y��k��'�n�@W�Sa$_���&�z1��g�[�߿�>�r̰���j�tG\��v+���lq�4z4)����^����_����\���� �����	���o��>
�WY2W�&���N{o���݄�$+�{?�� J)ER!+�Yu��ϳ=Gz��AC>م�c8��a������K��[�W'�������<�ր�;�Y�T�l�ٽ���ۗF޼��A���{��kk�h����&�H$�NG�B	 ��|ׇ�W̰=��6 �z¶�B���*[��[�̸ *��âPH�otet��Gf�`I$c/\�H�����FS���S��-�[��3՘I��2���	���o�d��p�o�vf�5^��y����[����(�U���	���q�@�}�0~V'���%͛�@?�������X�Ș��ˡU��R�.Q��ݜc��3v�=�W;^��M�;��(z-���/�v߁�4KA��`�h�#߰�����P�H�;+���]{"�zz�.���Ny78�D�V�U	J݈��� 0�:
w;nŤ[� d!��;[S�k�4��c� �ϻ2gV��z�����~$�fjd�M�76��i�=�y� ϼ4�����_����}5�=���r哵'E_&kjģ�b1��@�pnUv�;�3��6����x�TH֍MFB��Ε��P��=ח}=  S����y����
��+j�/�Se��m3�%ehI%i�T�H�7k���D���ѻ]�3K�zI1*�t4�D����4�-�x.u]�� �U�V�ʽ��E���v:`�{ٙ� ��a;T�)N�ϯ<�����0A^P����[�k� ������ro�L�s�������������ħY^����m� �>�`@�r����K~�'uw�8��I {^�f@yNN��UU$��n�bn �*}�{vǯ��o�v�@ g�vf��rs2�	l��l��Z���Kһ�*a���BMO_��c ���V��|T@q-�[!b���I�޻&�:���� �T(P��
��v~�%�[�[ ��y��{�n\��V�?
j�K�ɧ���cA�m���9�C���z�{�:�.��}�<AI����mo��/��W�x&���5]N���cst��~	!�ve�7�J�T�QE$T�-���f�����U	��ٙ�'�{ܛ	(��Pu�Lv��Ә����������sлZ� ��v�61��6�k�nz�O�9�I�U��ꊙ���e,⯟�0  ��� |�u���?v��>��Q=����|W{�`]?}=2UQ
j���1��G�
�x�o�#�ُo�� �+}��� f�B$�7ѽ�1І�����$������Sm�*h��X�Nm� &m�{��fF�.}�� @w�7@Y��7Is@l,x��q����Ix�+���}p�������@L�WY��fqosf�Cu��١���I¯yɄ��ƃ ��x�P�8���h�&}~�y���܍�� �ז�e�՛�p�>2��3-�8��wZ�;�̜�rZ4~|�f��Ɋ�q��������Y{���f��ԯq|\%^����¦��x0{��]�,���ؐ����#��(�'5ʹs�6n�����\�͹ݮC�v���Ě���gѱ�Ag��o�[Q�t�Õݭ��	bG�n����y�ܫ��v��me�2�pz|H6�\�q����hNF^Q���A��ةBB�'��\nձmXN��G���v�WF�t6�y�ۢػ,pB^ok�휒p�H�\wn㣵cs��'ܾ��PL9GO�ѷ�8�"��´�=�����b�p�	I;q��ͩ�����+�Q"�E�P��R�M�5f��ˀ>���̀˟{n;T�Qz��-i��O�*�kp�^MF�"�L��s�wi$: 3����̼�6��H$�Lg:`��٘�q+٠�Kyd��o��fETB���&���S m��s�@'�)�s��f����� ��k̙p�}ݙ3�+$������S�gf'�֫/�LWC�８&Z�"8H����v%(��N�,m�2��
3�*�)9�
�I��7.��;6�J��;�-�8���̽<�B�u�0�����o�7 ����k#޽Y���������l���nõ݈�,KR7ms�.�x�ˑrJjg7�R�$U*%	��+]y� _��F V����7=��}~��|�!r����$��
�A�Y�S�s�$Еf4�jՇV���%��n��M��eH`��39^v�zq����^�ה;���iPf���~L)�3q"�{ڵ'�hgg����?gj��������	����]ߒI%�9�&f`��$��:^{�~[�9�YQ�
&Rl�������[	��=3Y�����@��ٓ9�ɿ��`�U���	���>�u�A5��Ӽ u����d^�s2�H��t��3�p.�#OdM�$6��� y��BRRJ�H)��W� ��q���rdI�&`�f�K���݀��j�&�@
ܮd�eF��@�Fzi�K�-�=�Ol��u�Y,<rvx�vM���I�.T���S)/�%�Il&Ǎ������8gW�\��&J�\�g�^�IŻ�̙� ��M���ٺ� 
)B���}�f�����*��WS�\�I$#��ܰ +r��,1�8��Sƹ���rWUJ(DQP�S���~	�#�6U$�I�B�m#�$r��-2-M�4��Ӟ�\�m	�ktO�ӧ��ڻS�w�B�p6ԪR YN��Le��^oN�?$�ן:��H��}5	
����^i�[�
&{���Ti�94� �O��e�f-c ��ٔ�j�V�&=� ��&� �`ِU0���	�ܦ�� @k���e�S�m#1���|<�,������ 1�sx�O�IQQ��9�AP%G�e_o[f+�.:sa���wm��0��e��J�훢/3��%%$"�W|wcM�{+[����{ݙ��V���W��D�� 
���D�f�����,��f{���#�����]���ܷ��z ^��&Xc����*��o�����x,� _{XE�$�Oo�����	���0 �_��s"bNN���>�>�:�j�"J���I{Ɉ�e���(�6%���m����fº����=��� �^��6;��B%db�����$��=� ���f�,��1�0H��^);�.�e�ꟅԴ�/����,a��o��aiL�<�{�d�I7�mW�/TWB)��i�[�D��]��+�r���u�g�s�kf���\� ���I���4���#;�+��%LE�Lr:�t�n-��]�rx:��Ţ;SыuB�m�r@�d�(��Dt��J���e�n��&u��s�@��n_�B���o��L�e�$�}��|<�O)AI�S�w���g��+IU�Y�^�@ϻ�3�> ��M��£��و^��&ylRd�ʂ`0ܳ�ו�`@���\@����r����ǧ G��fd�j�&�[��
 R�%	��U���!^u�Y�L��L��}�0� ��[�  V�su����|����F�@7��v\�Lkl��EBUM�o&� +���?R[Z�\m���s���p<������3��>~#�@`OT=m���Z��rK�{۱���z!㓳ȴq��n<���3�OQ=���8������v��7Gέ�HE�5>��f�Ѝ�ݞ}���6gK����=��Ҋ����-q)F�uS�(ڭ[7�a��]���u/Py�~$����X�aT�l�L47t�Ny�s7N�U��,���:_��X���8�f���0�t�\[V&N�Uܧnػ���Ei�B��R�v�Kw�Х����z��{�{���o5���(�<�WP��,��o��r^���2��'�;��:��O�؟���&�ŝ��NLFrͶ��ygʸ�_=����,|xKT������-��Ԇn��<����%��>�2"I������+���ok���}�y �o��w�P3�'�MX��U"4�pS0��N�/nW�N^d�ޛ���Q�{6��ol��w�>�P+=?Ne�^v�\:�j����L����ƴ�r22�V�r�L��������(jz���,�3��wP�޽�5�ܘR#zg��w<����Sf�Mf�`n��'N/d�̉����A�"����c�j�4���;�Q�l��5Y'\�ϔ7V%1����	K
��s4Y�R����-'�א��.��Z��x��j�/Z�,]�cU�1zY��Fj����<{���G�Z��ܸ��{7�������7W����;�r�s{f{<'C�vT�s�O/i�b���n�i��@���0�p/x��{��病�9���A�����I�������:)��ﱔ���Y�A�VХe��Z�2"��PU(Ņ-�h���3#R��UD�k,Քb�)Q�m�
��H�Y;����V�V�bi�(��)elF�+"�Z����[imc��̥(�4�Ub3ٗ1v�#�3�̲�"*����T�P\�b�6�*�R��T+*�D�ܸ+��[�P�PE`�2�2���m�R�*�DT�,Um�U���d �Dr�Gn��һpQK�X�K���m[J��bb����FD�6�ī�Pt5���e�Q�J�"�J	���E1��keKs1��"����M�dT-
�"�i1�Z�F.i�J���)�6�TU�LI�t�iQ2��l]%RcUPnk1��Ӥ�՚�d3y���Z�X��K]e4 ��1k���GUR;hꙒ�ˊ�ĭF ��ҮaqT���Zl�Z�sZ�Y��i��"��ڠ���U���-�1m���h*14j�/�5QJ]��ض��$�W�,ø�{t��^N{Gj�;Zz=['B�+l���Ƴ�Ӌ��67.�r֤[���t�t>���V�Es�����19�v˺vwk�������bn�<��p�f'r��-�dl9����8�����3�����b�/^0���n��8����۱�	bے�ڏ85M���k�h����c����8x_j��7\�d}�����<��7 �;�|d:5*t\v�Wu6���z�;q��m�9�WZ�f��*�J{73ػng��{=6bh�x���;mX('��<|�%��;�w�qk�6�y��	�s�]> ����<:�
f7 �!lg<�3���mF4��fp�ͭ�+v{l�eF�h��D.��S��v�*sq̼�e,�ݸ�e���gBL�v�zٛ{,��C��z��[����=b�pj��j�e8�)ݛ�z��m�[��nּ)F�%N�v�Hl�t���{3y�RW���E�s��V��cY��P/n���>�][xsf.��,8�.y�4v�Z�:6�n�V�۶8�^N-������\���\�6�xL���f��F��t�<�]�=��糇��������͊�Ն�gW/3��X���h��!M�v��m�*&onz�lu�Xq�{s8{>E��c�o���ݶ��3��#v�B�����ͣ�\�;�<�]vz\���엨5�KW=�s�����m\lvoh��:�ArzΣb�]�v!X�'Jg˔�=W
�t�g�]�MgmAh��{NM�:�v��N�Ψ{z5�ù{nv�tS�c'R�f�NG�87v[�=ٺ���ْp\�����7+�����z�g%c�n�v���齶ax6�9+��3�5��q�T�(��n��a�` ��:읎-�ͮ��������}��k�hY�u�v���8.��6����]3�Ln+r��'7�v�����e��踭nL���/f#��u����]]0Z,���Wj������16ƈ���'�7�|sV��L�`��r�{)���c��w#������W��1��Z3���O]��ݡ�cy����u!{k�z��8͗�c�-�C��ϷX� li�մW���^����Ϸ=�͑ǫɮC�7l5�N�ֱ�5]s�;�����mr�vr�'�q�a��ۛnR�/7��qF� ���v2��f�[L�3�u����]l�֒w;���t�B�c�7K�pqr�!l��-�l}�|�~�SE�[[��D��9�W�[�>� �s�q �<b�K���^;ݼ��%-yΉ�V":�dQS�*�Oc;J��*�le���{L�{�nXL�T��Y WP9�r������^t��ZP�.U;��j� @>|�̟L'��Ue��f��]�V�@
�>n,!�d&�@,x�s��ܚ�2a���v�ڷ @ Q��8 ���P���s2��Z�����k�� 
)Am�S^J�˯$Nu�U��)�w��o��=nf\ T��S. ���̀�>mm�y�n`�@���4�)@�Ӱa�..{[g5��wܺ��sv�&\r�;~���Vl�h�J�d��}�O=nπ��o"��wO�Ü��^bo�� *o|���D��Q)EJM���gр |��u$�J{	Ze[æ�oip�(?����hts�g�,�R^Ok�:f��N(���tLˌ�%��i ����O_O9��I��N}L�I��vf@�r��D��{@���c�&E� �Ng&���� �>�� ���:�����:��>�����6� �}ٓ9x�<�$J�UT�s�չ��f�,�M�3`���� ���fd |V��؅ LNK��@Ѽ�"�O9H�JJ��P��k�nd` ��l!_z:�m�z	G��l 򽎜�/f��ݤ�IF�:����ۑ�#������`\�m�n��ܖ�Q��\�,�]��vƶ=d��JB1׻�C$�0[a��J�>�`@{^�Ȍ �+}���u�{��M����;���q����fg�yd^�HB�����)o&�}ϩ�*���yu2��{٘![�M��Q��}OC�dbɳ�7��D��J��I����̈����ڭ� | y�)�
8��Y�.�jʗ{3=�0�N��29ũ#��AY1W�b��F5i��S�0c�;�Z�\�B��(�܋<����y�W��?k��3 �
�rn �zLuDȾH�J��c9���ӛ���Ԍ ��Ȍ ���nfXU��ͣ+*�~�L���˻	/M�c�i&��*l�{�  ���}�_!yry� }˻�2  �^�l$�
~_I��Ǭ�����KM�Hi(��F�tg�1ɭ����뇭��fw.x���O|�>��А���f�BX�}��s�W�[	��X����ȃ��џnmu�6:��	8�sx	h'���l%X�����d�]�O�� /u�p'�?GUB$�����y�N1��o��}��4������o&�&@�խ� ,��Gq�9�Y�uy� �ך�M(�����/$<ebl¾�����}���ۙ=�@s�l�>�~^j�K�!���9���4��I�����i�h�t8��Cׇ��هT�I_+l�,�E��3���w����e�0f���բ�#��[�ϻ�P	���W�/�)T��c�m� @f����ڐ�W�u�l���� S���"�^��rdN�\d�ZXM"Z��=�s���
��b@M�'pP�]�ر/�V�i:�M%IQ[|g�M��<�n�>#���2��_�xg�ۚ�I ��6��O#�0� �n�;��b�K0�l���^+��$�
~�X� ;Ϲ���|꼲6=��U��fӉ�*��JJ��+ζ�k�yL����t�]�Z�� O��" 9�>���9]��m��l��iH%�����wY~ ���>	�y�f`Ƭ��rxQ����ѵs`������^H0x��������9f�a��bډ����v��� 罙3�A�97�m{��N)p�����д�>��ϓ�%��՟VOl�v����TZ����7ʙ;�/b��^~h�ϔ#GD����Kװ�vh8�}q�Zȇ�&�p��Ǉ�k����e�k��k���
��z��m]�7��.��Yd͹,l۶�&}��n��1���v�A�'���7N��_$�6���q��.:�c������n��k�u��Y�t��[��ᣏ]���خ��sf<{'F�3mǅغy⽋���z���q<���M�Rc�rz31wl�p��x����Kq�Tf�8�t��V��YRk�w4�C���nݛ;�|	�\��n5��==������^�E*�� 5�;s�yL��9\��6ǲr����ʾ�I>��w��'�	��RI���`R���f9T[uv`y�7�j�Nffg��tu~�
�UV?PE�k~QUD�
i���̈�� 5g+p�@G�K��g��Ǡ��}٘ �� ��sxH�o�J�}��ۦ�lf=ݾ� ��F'�F��r�d��W�t��#�oh=f�B�N}����r��@�J
�J�� Ky733O�l�ᢛ��AZp�j�OEk��E�����
�t{�rQ�d0�������q��۵���q��]tcs�]Wd��HY�������Aq}�Ϋ.ť䗒�z��?.c
�R�����ݙ3� ��%��}*�LT
U+>���j�{)��6�20p���:EA�Ɣ�ޅ���O*���������meۆ9���jQ�e#�pU7�IFyQ���9�cXf)فDDݼC���ן�  5g+� @M?W�Q33_u�1w���{� }m�y �JI!;pw�M� <�n�O���r%�����Z�y�	�嚛	�
~�o�.W��Q�Xn])��3ל�*%�H���$� ��.c �>�Ș�Ķ�l�����O?G �٠'���x���^u� k�n}��^[�$z�j �fۗ |W��L��#���0�E�f�e9��A�(4��	� bq���c�h�;�v�yn��G���Z��^�>��Z�%(*�*��R�M� @U�k�S$@�ﻸ�)��h�O%xy/g�a �'�[U��"f�X��8!��5!���w� �V�U]��j��2DU�s&_�vWuQ$��ٲ�tNŷ���5����T�@�Rl1�;&_����F��?���{"ň�H�\�C�z#l��dP¢tU�����R&�s=�-��{��"Do��B\���]����y0�`�S�߼<2&�ө$�Q?GUB����3 ���U�T��l�m:_{�c0�>gV8�S ���2 ��9:���u��@����{T����"�t�����H�o��I����//3gc/��kv��ɜ�I(��TM��nY���_a\yB>-��JA�m9�瞍�����N5��2Ƈ���IML��ّB�$()	�|�^p�� ׼� ���W39og�bu��3�� O�=�wk��M�Y	��m)-�� �xx��g���L���!'	
�= Bj;��Z�p�=��PC���D�%*�57ّ�vj� @L�2�W9������������ks��"�^��L��B�J�D��Mt9q�Mu_VZ$�}4k�$�ھݳ�?B�I��~��ޞ��]��|�������Z�{j+|�k��AY��-D#!݋{97��ld�j���e�Ľ��Q�l���ޛ��]����%{�~���m~�$M$��BN�|gcM� U�~p�1V��g,��q DVn�f@�nrnfO��W2g6�٤������\�iS�Vz0u����v|k�}��C���\��<(���~ۉ���%����̌	���n  *�]c����F"����)>��� 
����� �e6�`&�ل�����uw�{��b�����0" �+��ˀ ����D�Q�U��[k��^��I(SUR�Se-���@Wկ�u2�F]K#�w�۠D V�&�fB����C�ʊ�/�S(��Ul��g��W�7�� �+�p~^c�>���.����UoE��'r��,)�j�m!�J��i�t�k�nn�ZqJ��\O|n{-ˀj���2o�vf};o�[9ʽ1m�pGP��z��2��:��Ui�z5�x�:�}G���LnE���C��}/rn�6�f�ӥ��6�n>�7J���P��
)F$����OuTɞl����"i��Y�֎7=��v��<�eq���t��cu���v�����_��QC9,�7��P�vN��k�:��YX�bu�"����[�z����;e�+=�۵�:���v��<�sϢَ���:��;ӝ،	��mg�����C\�������W��b�`C����Xx��0���mή�(���5���۰�ʹ�4Y�]�7G����"H�%B��]� �m9� @U�m��;ϻ3�^A/f���1���bl$
��d��L
��
w+}�{� UEu�Ǻ�������> *�� ϻ3 �V�{=�� Dm빒�	*��iRv�
̮p�d�=�y�� M)�qq�>��` 
�W7Hf��ɜ��"��@��R�K~qs=�����^�:�����$�$���w�H��9�dGc��+R��I7={A�TW	|�@���M�Z�c��f�ڭ��љ��u��;y68	�;�{.�A#�9�!���-��!�A� �-���<�!�Żs�F���l��6�"p1.J$_i�0e�e��	edT��|��F3$j�[��O�Oʮ��?ucqI {ϻ3��I$�R���w�M�����*��y/̧�P
|�0��o�����3���^�u~j��c�����"�ҫQ�\d葖�`B&,+�;�%�.�}��?|�"u���@�ܭ�W��fjd@�݂]�F�R]�e&¢��BWn~��39�j�+ ��{�˙��~4�>�}٘ �rn �/��J�$�Jdv�+�\{������<`@e�y�a2��nX@?W;��c��%Q$�ٙ��E�$�)��*��M�L�](�y�k,VrH;�ۻ	y�9$�I�ԍD�[C����(O�2b'n��O=6��\�=C;���Lc�ӗ]�lU`7Z6;;`F�~m��.+����~I��$�	/�}J��1v�޺\ FN]�݄�Is�uA%�C]���X�ra=>Rd@__5G�}'�oOq0��\� &����D�μM��8����W��D^=���BJ�)Jv��6�ˀ>
y\�3ﾹ�����b����L�2��{b+4����6�"����v���n�ݩ��J��S��5��6Y����)xz��ɓ��=ԏuQp�k��6d������*����}�^m�\0�������_�����W�۬��_�d�GMػU5��7J�o����A��/7�MS1�I��_>;w���/��Ķ�@��3�W��sRs���N���m'\��a;�cԽ���j�W���Y옇���� P�l��vh�w�8�6�H��U��r�����>�ȁf`ʖ���P4�����a���t��� �n�!����$c�ty+Ṳ'B���8Q��l�� RQ5�M���)]]���T�Q<?~1��߼��y�N��w)�\��]��a�ٛ�2�y�B@=�L�8��^��>Z�����l�R��"�����j�:� M�O�yd���:Q����~v� hM���ތv��z�ع@����۳�{�Y�|��R�&�s�Y�O4�]K�p��~���>n�kî��p�_[߶v���u���cMt����!Hf���Z������f�Ѻ�Uΰ�Y��dU�n����j���;F����g<������f�$��쳉ͨ����m^p���Qs�/�w���u��⦭xE�٥NA�f�ˇh1�}-��#N̂�}���{��������L7��j��=�<cp�9�>��6%N�z�yn��ބ���S���h�g�����A�;����}���FG�,cڮo���t��%��O^��ަ�>KȘ�S-�jM���3�=_��Q�+ʦ���iDGV��5F�[r�,�(��V
��k�4�Ͳ�]4EDjUjo7���+(��"*"�E]��-T1,�\i��`��m:��ff5��[��"�V�3n��hR�EЬb��T�[e�,ER�+��eZ�Z�j�j���
:�D#�"�A��h�c�Qj�;��[�1t�H�媢"��X�Ln���ӧz�T6ҥ4�b���W2�"�9�Lv�)��iJ-(�YmSv�*:B�f%ƭv�t��t�E�S�D4�(*�Z�-
m�2�)�:ups��ʴƋ�2���t阥�.i��Q�4Zesyf��Y��ѭjZ��8�x�m��bN�g1������ ��i�Bɤ#PL��d�]t�F�7�.���;J���Ŵ7t�ڪe.�d�mM�XŚ�޴�]7��+P�*-M٧2����eݢ�)jkt�L����]Y�[V�QLs�7�$^���$ S�sqA���B�)��a����ܶ_����1����[  )��8� �ݙ��B͝�ǧ������ �&�%8�<�� ��x��xy ��r�&O�~�2e��y����=��H8��~~���֣�������3k-��#�#l�������R�o���}�jK#i?��ɰ  �ն05�7��z�}�R�گf��~=�G ��+�?��X�i�m�ebHW������G@"�tǲ�y^ <���|�y� $���M�%Q��$(u� �d2┪M�=�c���=� v?^&�=k�kr} S�s&fs�y����J�QIU)JU�A��o_��}OhGy�W> 72�� k�o �����*7�,D����<�Ŝ�N�b�ǥ�'t��������d+G�o�m�U��f�ǌ07~����v(��ۃ~�9�I��*�J\_B���� P������� ����W쭧^�;����@�{ٙ	^�9���j�OB슙T4,���0��{mv�ڄ�3���'=s�-�h�c�wYz�
T���)��i� �_�J���$����`|�-�[��zG^�`ۮn� �ϻ2g=y�*UR��*��)o&����(����*�*������k��� ��a L�>�P�Mv"���v�'b3W�i�m�ebl+��f` �ڭ�3�9�E��p�j�$Jέ�H���:%��@%2bp䚞��F�4Lp��;)/%;ݵb�	$�{�4i$������h�d͙�'~��ݘI��f��(��x�sf�F��@y\��L��>M��|�@L��jo�����ѳN/�m�Vs�����^F�(�LF�%�]f�C�����yQ��1K;�l]P�u�6�.��4}�k�ҩeJ9��U�A�E��۲��X�5�]��6'�Z�����b�Ea��۱�,�v�;�E�܌x�����{]����1j�Nʾ��`��B�����.�+v�����L�\��7^t���l�^f�n��ݛ�e9��J[[O6�&�Cb�f���K� ���ϝÃ�����=p콎Ѻ�ـ�d�l[!܏Y`����.�-�ۄ��v`�ԃqS����Ɨ/���,c�@vmۧ;�c������*c����C6�&�ົ6��  [�V��&H���?���%�ۘ�gg6�t�����e���I
� )�?��� ���{��0��C�d�}��}��e�_���$�i�ocje�6�M��{c��	�D2�0��)o&� *��é��W<Buq]�f �ܭ��~�o�ѓZ�!�P ��
:��ͮ#�lD�ڃWh�a��[� �W���"3��dl���u�nI3��y�/ �	E���R�@c�n3�{�#�]x�s�O�:��K�`@g��$�7�y�6Ml�S��7TQ)&�1�Y�)=�,Mζ'�H
�u�GgnY���a�qس/����uH��RQJV��i� 
�9�� I�޻'���k�FW ��]RE�J��!.3�6�&!��
w3�� �p�w�?:1����{y��f���-g�d-;��[�^Ѹu�d�1�Ӄ3�j�n�.�k[��-�u�{{����3��e��� @
�y�� #|��2 �o���馶����ݷs5IH�JM?��g?�����}�������s{��̜���I5��gU�D���݄�nz4�i$�I�&��몎vg8��6��%���y� �y7^c��=IJ���{�A�GR�P"��Sek�̌ ���V�&f+��;o�F�n�`|o>�̀ �o�7{W�ں,~��x�mJ��\Na.��'/3Yϊ�3���<8׷̂������0`�8�P�Z��s�KiuL?�g���}�� m�ۗ�{�]M��o�ә'��� �}ٓ)�U)"��T�(W~�:�n �������We�C@���ςd��a F��t{�go���ł�f"S�h���v�H���k� ^I�p7L�Z�Lck�B�Uv�$ݞ;γo!�C��^����ؤ�"h�r�!��"��9��{L�2el�ۀ��$�����.U��jݞ�zڙ���>��	��o�7�m��e�`���J�q�Z�P�֐�L�߽�0 &W���e�7�zۙ'<��2��p��ٙ�EnG1$�(e�0Ң�y�$�J�P�['�y���3`w{��� 
��7�H7��p؜3T{�9��h��G������
Y�ۮ'M�W��2�Mt�����P"��VI�x�# &k���57��6,�Mú��?f` W{Sq{8B�%%��[�2_7���'�~��{��73>+}���S~���"��M"�U�#=����۩IRT�R���f��  ���N �&k�����=�r��H
��L$�7�o谋Uډ�%5L�);pk�n\�(u�8�٩��м�V� 
/|�5�7�P�֪zsd�n��ŭ�z��z'n�������t)�yLu��ܿz9��b��>�#�a�����2�;4�\�>���������>�n悔J�J@��d�{�́���`�V=�n���{/���&H*or�J$��%�f��s;����'��瓃�\5�nkr���׬Pp��Eڣ��^���HRT$�AK96�M� �}ٙ�=2�:/k/����l<���H7�n�u&h �J%*����f C���p���g+� ��i� Dg>�ɜ���P�K��X���"�*	G�E)�M�d�n�@o�s���o�ɞNj]ן<�؀ *o�ݒ|Ϲ��"��Ԥ*�UT��'l�m8���[�3n���ggϜ;>�|���k}��w+�4��H�޹�JR�1�Sl��dQI�������
��[
u�j�p��AS�u� {_vfD������Ur�������'� �L�8s���>;���x�����{��˨�����ؕ*�[c�_\�ꢍ�k4����y�3G��oͷ��k\]n-W&n�4s���uɳ��ka�7[�p<s���:�6�n�8��D�\�n֓���6�&̧dM������dRݹ��l���e,����Kn\��;g��&�7u�p0؇�p�V�b��;S�"���<��ۭ˺"�eַm��˕N��C�1��NP��ۇ�w=�J��G����M�n��طg:+ؓl����-	�j+Ym���Ysͻqq����:5Yq���y�O=[;%go�����&4�`���*w<������D` V�����j��;z7<����K������;BI
�))P�����s/��1޼K��#�ٍ� ���@o�7�L��w;����7ld�`����V)T�\�c�	��j��تO�~�dV绩���}٘�[�M�����k͈f!�7+�fR��h�0L�+��79 @W{m�j�]jg�>��}N�f_w��g�^>��(P*�T(N�ͦ� �
�WY���I���3�U~H���+� �r:����ٺ�N.B���g�e�m��3�XJ�v��6x�s�I��k����H����cZ�غ�_�ۙ��^�+p� W��&�ʓ��������w~I$��3]PI_���R%P% Rt³+�:~��͕9qÙ��Tÿ_e�f-�N��d��H~o���n��P:Gv����T��Sޫ�8�O$�y�)_Op��q�spz���
9^�O�q$�J��` 	_���H���};eFwj������#JiRR���[��  }^p�����|^��P ⾾p +j�LD�Rf���QQR��+����o+�V��X��V�  ���0�3_u�u��v,GX#Io�H]�꼒ha�j%J���c�m�;���#7.'�����W.d��լ�pFk��w]�������|/SJ ��Gtn��t�r�L���'v�H"�,@�3���i�\��J
��(V���`|_�[����D}��߽~�u|��ܫ i'
ج"~֪� ,+^�;�c
Pr!m�ߌ�j�3o�� |^�1��ϻ3 &}��;yӗQ�L�3���ҪU*�B$���Vem�&s��s�|
��:��Uo�%�ymV��f?+�i�eWǧ$�~��f3�Cc�]}���2z;ufЪY�+Q�h�o��ek�ܹ6��������ZV��  ���&f^k�����-&�L����pбM�+]Z�� �k��� ���'C&z���ͻ���@��t�I���P���M�V�ّ��]�V�gRN�z<� ���`@���0 ��&�4{�,ظ�8�KT�m�8�ч;�������J��x�����a������o���T�)�[���v?���>��  "�:h��NGf�z5�s���2�Љ*���0/u*�(UP�83�Nfg�s�k	��I�?� v��̀>	��+iNun=�PMK���BB\n4\CfD�0�k˫;nŢP	Fg9�$�w)�YO��� ��}�� ��!'�q�A�/8����N�]댰���} [�. �����I�K�33Y-�y+|[��7�q������ �.���{��{2��k�Zi�Ⱦ�o���3 ��w�*R���GL�Q2P���I����>����0(IJ��]ɿ� �yåqk]�iʝ������� @n�n@>�sqE�_��d������=��e��[/[�͛���[�e��]CX��^�:�3v3�0Y���;QhC�Ҁ���m�g� V`D���e���&�#e�F��fL� V���9Ϊ����RRR����: -��+�#s� V���  +��虗���v��@٪��&I^=b|���H =��L�Þ�Y��w[� ���	> Vo:��j�UIMB%Rv��}���w�v) @_>V�� W]�N /{�&�}=�맖��
��l;�N�P�TM(JD��a�t����s��^w�]�9��F��t_+�2@��7��2��3"��w��n�.���x�6�7%f�v�μ6Fn)��uV��z,8V�o�S�^�;u�]����Y���J�W�5[����W�4Ƿ��{m�zz��Ί�� ��;v@/@+ v��b�{�rf씸 ���:�w�˪$��X��2�y�o���7d�"��G�>pz{�Ob�n�!Yc�������ƗE8�ݧ/w����J�H�f�Rl*��Y�ŧkb�꽲�Cъi��7s��=I��K�o��Vr/5�lL貫.��X���fM�xI���g�2��9���b �#��T��s9�skj�^�1S:����5�/q�̗whjV�툍O7���>��ӗ�e�u\ &�{|y���}�����u9i�j�'��͇Fz�ˇ7w��\�����|<s��{F!Ȱ�����`P��et�wۨ�j���`�O�b�Vh��������_b�Z�?������B�׷u�Nn^�{����=K�mjo�P^D����U3C�B����G�� �]zs.�p��nr�[�æD0"�dqhD�v��{�z��\5�5Nܸxo��8/bt��H���.&uSܳU�m����i��]���]G����������z��q�+����tM!��s�y�%��u��mV�ˡ�X�h�ѨZ���6q��Ýݥm���2�V��![���2�Lh�̫G`�|���׆��}����v��� ���֏%���4���-4���.��U~����G~�C �{u���[�SV��R�e��M5
�b�usW���٫��QQt���iZֶں�m��%�X�hQ��ȭj��cF�����1CMIFZQ���)DVZYYX�Eq�R��;pqF5�����L�+��4���DVZU#[&\��R"�.*Q[h�0����f-����2�]2�,�UX�2�V����������D[n:f6Z
�dպ��q8cJ�J�-B�m*���c;�wlDQ�W)SY\��D�۫E�D�҅bU˄U2��H���F1�
�̓-S`��UX���U��u�-
#-mb(i�Z�T�i�wqի[UWC�Ҹɬ��U@Z
cEb+1� ���B�ۂ+b�m*2�J���QUV�����&R�奥e�S�,-�P���[��BU�e7>�ݳ�n��;tK����ÔlX��1���Mu�P�e��i�\����W+��gy2#��5�����{V�s���syP�6��Ӂ���x݄���t%�[mˇ/0TA=���煫�;N��Lu�Y�;]�p���.ܮ���p]���N6�\�C�m�r%u��[L�S�J��HZ�k�<�m��הR�l*��d�&�:�lG3��w^�4^<�kì�e�p݃���5�ɳ�Pӱ��Ȏ���FיwLm�^'�1c��6���86mѰ���6���ݻp��['86�;;cq�cn1n]m�X�a�h9�nz�7v:5�ۮ�ś�n���[������ہ�]��b�3�D[Z8^��sۇ��	3�q�)�y=���x�;l�z��s��k��crݴݓ���V�b��l�&�S*s��k��+�==�f��h�OP;�=�I{tF��p��ǡv�n���`�I�F�-�������g�n;q�oW�g/W@��g��h�}n\��lF7�;�C����(W�Q4w^��[����h �xx[������-���Cֽq�۫P����c�Qw�D�ƽ�War����s��Ϟ������g��m���ψ@�)��j�8�N:[rvݶq���\�հ�
�v���;���h-���Ɠ����lE�铱:Fݏ8��=+WY��uìW'D�l�j�u�nϭ�f�s�z'�/��G�==3j�W��Z�:���l�/3Սn6�i�eЏN�ŵ�Q�ݨf��T;�.��=p=�e����ǵӎ�e�����k�y₷C�n�ps:{q��	q^�4v�p/mq"	m�99��ܜ��;،���J<��q��xz����f�v�]v���e��r�� ��j{{ld����=�G�vX7t�ln�5�2�wn_n�_���q�'=]�c��;vtZ`n�ܱ��6觋sC���]b�,7�ݞ�(x�k�a)�Na����m�vmɱ�3��NK��:x.�s���v���I�gN^x<Y�}q��&��4�mZ_�m����V���qE�!�
ދ�g�c�n���燰MGCC�n�z5\'��H#�A��[cd���\w]�^{
���q�������:Î}W`�:..[�ޠe؍{Ƿa8+��)�^v�N8��4ȷ��k�W6�#��v�mi����Y��h���HD& ��Љ���XioyC�uPʳ��&H�������XGxJ���p2
���A�9S�*���%SwݙL��ݺ�p��� � u��e���ٙ��b��E�'��~��(���@6�nBl5�� 6�y����:��~s�����;��>gsh�����πy���)�(�9�������I��,$g|�/�٘ ojw꬛{j��R�	Zg[�k
RSP�SE'l�w��@{�[���T�5��s۝ n��a2G^�fd��[ڛ�⫱2�(鑣ZeCP�"ix�c�tm�&Lhۋ�����h������~�?���f됗��
����瑄�[ڮX�;�+�h�{^E�E$��o]�J��R�)J��P�K�7 ���U��|Fv��z��0��������u�#�����z5��"�(� ��nc�d���2m����$2\{�ȝ�VҊh������ܫ�G�2G^�fd ��! �:��/������Y���#�'HAPJ�૽�� �u[� �"ԫ����^yU���؀����� V������Ԩ�UT��I�q��oN͜|Y2�Y�F��IF��	��]\T���d��ԐS�vM��OT���"SO�:�s,���gN�P��غ��5��s2��^:l_dA���ʮGF�%�&P%8P��M�̖ڴ�����Qz�J��ô��O}��*��D�h���_v�f ^�+p �>tî�t���`���o�����̼�ZjI��B�$��U�͠7S3��=���|��]��, @'����07g/��;�v����~!�)&���
�ॼ�� ��~SA"r�8��2+��،{q9N��&�q\��)۝ӽދ��E/���[{�8V�$y1L�}��ֺ{G��eA~�z�&�n��W��@ �ɰ� ��>o�ڜ��QHAPJ��M�A��YV�����L��V����L^Iv_u�Fj�J�J1��4<�	��n ���K�(�J�E$�s�~h 3s��q��7����pO�ˀ�
�~n�>_��2�f�F�ړs�(��6��kŻ%tǝlJ�����9�[m7{B�lR*J
��J���D�Z���m6�$���d�^���z��k��tj5E�&�fO��>j_˭m(UIP��'l���� W]Q{��e����+�� �� ��ٙ�/���Bǘ�sw����a��Yx�z���:zM$������ mR�^�ش:�v����T���$��w7�V{~!�)&��JU������\9�D�� ����@����� � �|�K&]�O�-��l�s�rN%�8�q].{N��+��e�ӵ-�Ǻ�!~�n���w�c9�pz�ڛ��L�֏:�I�4wt�f�W��@m4V��5��� +��+��zu�g��ҹ�ay�8 ���̀> �|��mv�X��#��+^٭�Kq	�7n�s٪֎�kA����o���[!�����v����;������%JW3齿��gw<�� 
����u���'�޵:a��d���7�9u\�S%"U�g6�� ���m�-=�W��>�ݽ�� Z��&�Tj9��꼔���0�!�a'!I�1�nf y�2@v��{��+_����o��Ȁ ���o��#$�e�����O��ؒ��~kӻp��;�0  +_[�� D7��q�.&�u�@�^y��)�~�)&��JD7^�� @T�yþ�yѾ������^#?f`�Sq RK��U	Q3�s8���mR̹�Q���B� hyC��ݸ�Q�.�{�dŞ���~��I����yH*�,���������34v1�u����:�١s��3�1��I�" 1���d��qa���0���(�������N�.Y�y��l=R�M��R/�|�|G��읟+[V��X�s͋���Ò��:w������v3Q�.O'���yv�.@�mۛ'l�FƬ]��]y{[����O9+uuɫ�6�nr��sh�xL.&i8�{�������u�V�8�cq��4mכ)�c�l�N�7{Om=e2OOI���߿����qԪ*	U���~�9 s�n  
/y��,��^�:�Q^�������'���c�D��	$�$��ͻb���Ǉ���0>��|�\�T��\��݁=x��hI�I�MC	P�M3|�l	������V�̷J��:��6|AR����[JU*� �);���<�rG\� �q[��d���4�d�����j����FXu�&��[R��(BWO���d�I�oU�S:&�@K���&�H�v�J)$guݤv�;�]�,��'W�q����<m�3�G�u<��]ح�T�����B�����ߎ��"%4|R�&�K�M8I%�����2л�G! ������YM�5���]�H%��9�j�^��Nc�莢&��q!b(Fu��Nu��b�0鑓��!�P�jRUZ!z�X�D��3���ۧ�	�@�{�SƦ���$��Z�`B�wfL��N%��++sev�ėV���e �m�ۢp�N
�I���Z$�3�8z�����%����d� m��3>�.��jdHO�m>�m��ڋ�@ζ���Du�{3 &CWby+�Ԩ���˝� ����"����(!Iۈ&���ZI����+j�dLm��4"b[� �����V�&�\Mt�]�W����v�T9��;�=<�����G8��5��p��9�v���x�+s������I�W���3ͩ�w��}��V�[��ۙU�N��͍�Ѫ3ʹH��̙�~߇3JD(Jh櫵_��"z�e�dYM�zڙ n�y @Mob�$�W�wr`�����~�߱��X�+Xi�T�����}�� s�n � /c�|:�w�)X��v�����]���h���(]@{�h!W���K�=�v����@�!�=�_���VL���] @�w�3� +_&��͏9RT����p�x����M8���6�1�a2@����U����M���b���|�|��dE(�$HN��`@g��4�y�t�[iWV��r~�̀ +���	 $��[��7�lE�Bq1�Ois�Җ{X��
��;�����u��1A�$�7��Ba�
�s�egm߭$���s@@@u��-�s:���=��<o~ ��ɰ3j[R�J�
��'S&���=�M�������g��: V��I��
�U	D�Fn)���8dˎ��S��q4���)�Cb^��57޴����yu^g�	�>W3,��ަe��G`D'�������9�,���N^{z���<���  T��	�{��i���xx��p�öJ�\m��r�
!DM�7�H�G���>˸t����Gj�`�C.��A������n�.Ep�Ƿ;�$l�I�,<e)cnBxOM`Oľ��N��ߧ��$���  B��F%��wiU�c\>7I�A��<q�OT�3�jt�����������N'�غ;��}?���QDH�+S�W� T߶�ˀ]���2��ѭ�F�|W�a'�7�5."�ѪJR�������3 7#������^�V�e� E�4� ��wi��F��ۛ��z��5�T�I*H�3mL��]��`z�޹��j��Ӱ T�svI���&�|���E��Ro9�=o`V3�Z \�6Ӏ ������>+_&e�;�^M��������q[5QT*J��U[���f}� W=W3Y������[W�T�e���{�3 ��n�����D���q�/u�m�ޖ;�Ư@���{�U�C��^��.'ޓ<���^�0��@!�'�~��W�O����w8�[CA'� ]k��[nL��/0QFǗm�'�^�����my�m���jW���î�G]�v�1c�q�;)��6�q7U�M���������r��ù�u�u�Y�Ξ���=V���,>]���\K��ўm��)�+�N]��<�.�E�4=m΋�^�wp���йjδ�-�'&ŭiYXV�أr�7fݺ`ы�l&٥a|�k���@Ӹ�ay���^8��^{[�m��o�_�2���X����,�4K�}���+_[��^=�I8�K��һ��d̗���π��t��@D�js�^�$�v���<v����M ����̀ ��|�	]ɮj�ER��S0�2R%�a����T:�s����$�W9�$J	Q�w�(��Mw<	$���fL�k��f�ji*I"�%+�����y]���"f�>�������� :���G��^�͓3���f@S�����)(�n�ɸ�������]sW��#|�ٙ Dy�M �Pv��ҫ�q+�S��7f}L��]��8��&:�[u����2��c�&a�L݈���8�OMI$�^�n��` b`o�@"﵁�/�nyo���-�30 ���l}��%(EU)SU	&�J�]K���wr�GGH�=2V��hD����b��͢65����$�PHp�?~:ۀ╅�g1��.u]��wOJ�Q�ؼ��} V��, >��M ���X[N��K�s����q+o� �rŲJ�$	���s.  ����� s������t�^�� Z�62:��]�U(�TIJ���&��)�a����v� 
�깗�L�[O]8�"��ٓ��p�ͣ]��.w�BO���$�m��x�P��� ���}��ͬ�l9ױ2N|<��,���|�$/}ݙ����V`B2�vw0F"�%Ţ!�[(n�b�N�u�ngbG.����p��\�������&�J&�7�K��� ���D ^��3 oE�[�M���a Mx}n�TeGT	 �%U���fF;����c�W� 
��t��/;�3  W���.�-�܅Zވ��9)B*�J��$�g�D�ﻞ}���4�L�ͧ�MءeB~
81I�m<Dފ}�@N�yŧ�=NAa*���`�*���s4oP�l������[2{:������7�םr!a�`����6ַCFKnV�M�'q�/����Q��
{������;�^��i�@wổn�B���<����EY�HFE�&�`o��^���Z U����s�.'�����}쑷��V:������n{V����W|�����j�U*l;�h+|��=X�)C����L�p�l���p��x����'n��H՞���]����d�uA��1Y����/o��|������3m��7wU=h�6�J���MMhDfE��K��g�g�j�X����g��p5Ǻۤ�"�䯮z�oF�zR�c��:�d��o����K�G�uKZ��s�ًx��}�ws�J>��ڶ67���ǵ�3� �K�Ӿ�#���o{�<�:/=���ys��7�8�h�w��}���Rmwv�<��|�Q�6F	��\G���_Q'��j�1~}��O�tzo��f�����y�}����@"��ۓ��5�L>�-O:nG5Մ�ދ3���Vm����T'h��}��ި����]j�`#t����c��Gw��d�G��ɪ�v'r�\\S��z���seƻ^�m�w���s�_��C)?wr�u�4�L��VlY9����⺗�5=��&|uH^���,��f-����b�#<�������[��"7�Y�s�ɌU��Z�K����vg����J��8jwD�E�B!x��PB(�������ƻe�(�q��R�Y�jZ�iPƳ��c�F�(�֢��fc�U�F����YX�Ңn�Y(�TRQV�MaD��lnf3no�QA�ۈ��Uݪm6�����]��4ۛe].]꣫*���W��UT�#6�V;ى�VZQժ���T�Q5VҴ�ડ�@Z�Xեt��b�5lMZ��V�.f(�J	����b�Tv���PFҳIb�D��TĹs(��q+&��t�2+7eĶ�M2�ALq�m�Z��n좪m���6�pJ���Re�c1ޮ�EuJ�Qus
�s(�m�T���V*��+4�Me4�G-�a��Ż�ͷC+��QZ)�kX�I`�����E�6��
�EJ�m�kQ5���.L����ƍ\j*1kr�Ү[ndnd1Y�EV[S(RҢ.YX��Ub�HV�J�2����ֵ�4P�W.J��U����*5��\ˊ�2�J.8�1E���T��"�K*�q¥b"��KJX��"���;���s�缂k�)��&��&�-��*.�y_6����U��YWV=�>fs�� �w�0
���rr�F�{':������6�֍Q*d�*�);���{����l=����W����Ӏ�>����� ���n�*|��i��sCG4�eDSB8a`����u�g�vvG���l��lq��=G
?��_�I4�uԽ]�&{�S'�y��0 �:�����:�^�@�|�$��wfd_��D"�lMMy7���TY���P�<�� "���3��
���e�|���t�� ?MC�ǜ��A�(���-s�Ȍ��5\ˀ�]�d>�j�.�\����	���M�>��*�J*J��a�c�K��B٦������<� �ͷ, 
�\ѵA
d虂Ȗ��E���eN��heߺ�'C���w�~Y>C_�s+�8MJ��6K���sZ��=�a��D{�y���{����~5�E�p�_Y�4y$"����Wd����	CE����	��n�o�lgt<��[}��L�vr��H����%�XT���Y��2M��&,�P.8i����BA�v5km��Q�ur��93
^�t��������7JUR��7�ێp&k���$V��`�[��9e���}���|]��'މF-6�O'�a.r�dG	���O��'=��y��@W��� +\uW��Ԍ�$Vl�v�w�	�(���^�� }\���@W�:�vޏ��ⳮ�� �����fe�������S9�E�IA*����g�*r�w:1 g�� �Ƽ�%�wfJ��I��&� �m6�=rR�E%�)+a��۩����y�)�^nLZ}^�΀!?u� Z�[�H�����UT��/����jr��	Fz����Q͝l�+r����Ό�2W�n���W3����'uBo�b�y�=7�2�rf���au[���]WȎ.�����B�÷E�:�Q�W*=��Ω���fu=�t���
�`�]:�)��۶|�x�M�f��v��'������K�LW9�yݹώ�����=�+z�A<���oQ�Yp&�uU���=vۤ��m�L͞.^qn3m˺�Iݍ5�e�;]fܸ�\u���nv�M��q����5�;t�c������`��\��a���9�=�{�����ָ��W��g���.@��ߧ��5@p1���Ǽ�n  +ιâ ��o"��i�7���|U��O���ַ�Z�̓����Nh�}�A�@oOk��/pn��W� ^k��/;�2g}+VA��]뙸�*���SR�E	B�:����}���w<�&@�87N$L�n���I%T��E$���3 ���qP!%�n����E]� >�V8u2@����LD��,��P����;eݽ�*d���U%��R�nf`���wG5�6�� �l��W��$<��	+k�����|+�~�;iڶ��ɵ��Ľmh���?��;���e��:�W;�����������u��Ū��ʪ#�����A$���$K5'mL�6I>w��@��K8��I��ꁾ�s�A[��&u��]�=u�&wm�KfLnc���[�RS�+X]j�{����w)���͐�9zK��!���4�ޡ�/����5q�r�Gf\�Q�uQ �����YW�5À�N���Ʋ���MDCs{וD��u�H%�j&�:�Q/3��Ims�d�S.m�P�*���JΝ������5����$		�uM��V�����@
�@�x�D���bI ���y禮��@$Nu�
�����h���O�亗D���۝��v�GgJ�k���n�!Ŗ�%�5�x�b^�a"�֏��È��)��?���
��$�|�oW�5UY�^��멍wYT>ms�g��Q2�L2ېjw��D����dn.���H$���D�I	�}&fw���3�մ��AQ��J	6���e� ��gUO�������et1Y�+eh�YĶ}�^U+06.r�ú�W�r�/DUXV��aF��ǝ���[��n�C1";��a�%�vл���$���~�By�TH��V�BM�Q��U�<��R� ��9��S��I���WF(w�����&�yF%���V%&�=2 0>�}���������"C�:�S��H���r��v�m�����D�2�Z��6�j�u�.�pWk�'/��͉��������f{Bh%����w&� =s��DGp�a��V*g]͗ ��}���2l.QQE���ؗss2�n�ܲ�G��;��-<�tI �!��Q\�uQ/Mٻ�JcQ�x��n�ʈ~n$�-�7=�B�#g���I ���t�1���.E�I���Ds��@�&�,Sm$mT�=]*NN�.B`�uP�I;;�^�����D��х'�����J|�5��Z��%U�cN��<�`�O��.Yڞ�{-�T�n��(�1K"����k�c���xJ�ӨC�M�Ux��icBm���m��yT	 ����"U�)��`��������V�1��'�;�T��F<a3��ro>6n��ׂY�������b�˃m[Y��<l�37s-��7"(���ns�k�O��H�â_rYq��s�D�rwzh���%I.h!&���>$����']��DN��UB��> ��D�Fw=~���5�i�r����Wn9�x˛�r���fE�oU ��b};veD?6a�a�܃s�[��'*2���$}55�I�̟I"oQ)�hL����]�B��-Sm$	o�|�� 	���t3%����O���> �a��Q��蓛N�C/��"5�u2�/3(8ؠ؆ƊS��=�F���������mx�����7�q���Cມ��;uٟߎ�����7jᇊG:�Ÿ���48�؂�X��g�{P:u�C�Y8�9}u��w�GG\����y�۵m�����-��u�U�\���ay�� nW�A;[ȓ�w�ے�.�0���\�6cny�	fM��|��P��>Gpo�;|���(�q�/��suv�M�Q�S��x}`+;d\�Gj��۷T�eS�v�`:F���.���	]�k��N$�u�����o8��WF�y�k���?>�۶�OeD6����	+;��|L>ު;5����9w���k��}l��@���W7�(��o7#�v�{�g J��I0�z��\��o7D���M��*ޒ�ᶁbjA��s�A ��ɯ�&&�z#[����Wf?H$C��S6J� (��B.k�7�Kq���q�9 ���;j� �{�S�|O�{�	ݯ@޼4��6`&{�v��4	:�zB���Oa�Yӻ�ĀI>���@M��M"�|c�C�sK'����tv<;���:����m�Gl�[g��A]��� ��Bh���6�A&�s�;Μ�D;ͯQ�}o{����i��d�̐bo\�I���^$:��&�RP����n /H6�~1do����gh���M���3�uYv��wF�ݘ��v֒�^n�pu�ʱ��L8���G�нl��k3��o��w��t�����O����(��M2"��g[vN�YL��p
n DP6�s�|O��ޚ���f�E��C�ʯ�m�uQ*�I �m�X������:��$�n��o{��!oc����L�1� ���hKzJ�0ANB.Ls���n99շ�[s
κ��&;����>+z�6�u��Ov`�h���)�ѵc�n]�#t���n���qŌ��tb݆ں�����5�bm�{s����+z�H*E ���2;o�;x�Gx�"󺨚�+�I�	�|�ω"s���01�����x�#7z�A%o[�	��Ff.c\vw�Q�
�lT7u�Ux�Vu��z����{zΪ90��7����l}��vQ��Vw��xgq�k�o�G��ux2;n{z�`����z'7s���S�U�]z9��^߇-3�W��p$��'�-�rH�k�������Ĥ�{{�w�^� U�M��AW�"|I"oR�\ɫr�����t�#bt�,��A-�/Ę{�Up�gDrg9�\��7�z�ĒVe� �!���K�uɿ[$�C��AbA����kaa"��Ϡxg%�hx(5ӺF����݇途��"�=����$S��
�{�RЮ0�t��>$��s�g�̨l�Ȇ2ېN�M{0���G�ja�'���bI��O7�W��������Te_�7$�a:�}R�	)�u
s��EM33������嵏�	Y=�('ɨ�Ay�
*���ڝ��r�$��>$��o�W�}�V:�)���g'Q�z��l>{��I������_�f���;�\V��Z��Շ7lN��e`�J�1�h����I��ٸ�����}S5�0g��4�F:����s�8���>ۓ��C��q"��{���&o���l��6�s��@���$HY��@�wL��}�P��NO{L'-�d����\�[&��������jM�t���p��ߟߟI�p�@�%�5ے|O�P �;�ꢸ�Q"Cͷ�J읪���b6 �81��=^�����gq�$���hP�!��P���,IQ=���b�xH��&a��eÐkv�E�;�P$�f�G-�ZWC�����];TO�+7�Æ����� �M�_ZP�7ǲsr���� �{SD�^��Q$�9�w�ט�Ivy�9��Tr�`�6�E6�ko���|T�1��U1�� �D�t�E3�?y�E7}�[~�$ I?�BH@�؁$ I?�H@�RB���IO��$ I?�BH@��	!I��B��D$�	'�`IO��$ I=!$ I)	!I���$�XB���IO��$ I?���$�xB�� IN��$��1AY&SYSEQ�Y�`P��3'� b$�
 ��B@( 
J� TTBJ��JIB���B���T��
� H(IR�
� qB.ͩQ6ʊV����X2(�ld��I@����*�l��1�kl�hb�D��Y�V� �i�T��ݪ�hӬ�Wf��Q���� (       �                          �         AH}�
�3|0Ѯv8�v����UN�����}���g�ۚ��7���n)���K^cJ�� ��
�������vUs�e�L�*�ig�  �R����l+��V׀�Sн���M���B�j���s�ޜ��;}� /��=��G������-�n��ϗ���ۚu�Vm�_         P �籡��}��C��՚�_/��j�}�{v���mw�枾��|�����S��ou/=�Q�>�{��fh�ox �^�nw}�v� |�4�>���R��"�    � ���  >�P� � �0�ް���= �  C��  ��;� ��4�}���o�7�  �z��1*��  �      ���>��` C�@s�r �X<��zP// ��A�G���ǧ-��}���y�;� x����wm��Yjڲ%�  d�Ҋ�g Ǹ ��*�c�A�2���Ğ�>�8 �,�$/g.���>��d���}7�F�m�T�  <         n��b�s;�ݚ�r�;�Ή��w�6ܚ"�{���1��TX ��r���\��M�l�f�V׀  ��al� ԥ� ���n�nn�,j���{,�9PK 4*�;���D�G=�u&�=�M��S5��J�  �        �=�q�p�>�s��U��^��� �=r҇�w�=�}���������p #/��9
�ܺ��P�.��ƙ|  �7���1��� �y�v��]>j�!m��@�c��*�z� rzU�w0ۖ��n�];�r{�x�J/���*(� "��Ĕ�@ 4 j��i)J�  ��T�i*$  �� MR� ���H�L�B� 1O�_��s�a���Ha�L��|��~�5���@�$��3?��$ I5!����$ I?�	!I��$�	#		����������i滗ffxo��9��kt⑌�k�С˵���5^F&oag��3�E��鲭Ƹ؜Ր@���鷎n-��$����u@`��$���:9AM�v��p+4�A�h�e��R�u���1�/+a��웩�%�F��*�g:`��71���z�p�Z�E�+n��ܘ�.ٹۼoqE'>	��B�1AEι�;a�IC��fm��ɖ��Z��КY�ٲ�K����)�����[�y��&���<��"�<�S�7Bo:�����1Iv��� F��1�[���<�b^���fH���1��d%Ze#Ft�v
�&��nW�n��xވ�
Y�y��+٨>�7/)���j��.�P�/��&7�)��R�\�q��-������9�e��S�D���ʛ�B���Y-Ă_;���I��2�F�=�uP+JK4q�*����WpG�cŧ�'+�^D^<<_t�gn[l9,ȵGQ�j���oHy�H�}�3rV���wf��{y��F��t��S�C�U�qf��&�cԸ��ӌ�>���A���Z���vN���H���"1!�)(b$��E�ͺ��1���k�\�2b۵�%�݇�fGs���^��#�7'<����ynsn�R;AP��y��K���7wMb�k;��:��D�q������m\t$�٢�	:>ʌTSE4j�Z!�5��n���g^�1l(6�J����!s�'J『��Ѧ�8�ƶ��cP�E�)�Vv�Zz�X��ح�"�`�`�z�ӄ�*N���)\ó�9��G�������>���{So�!��`��bǆg��q�R����3�/}�.��	�*V2P덃��`gygP��Y���Y�)MyvE��)��nS��T3��6���q��hx�ݜ�-!�����h���Cm�N�zY�{����tNs�M�vf�_.�:��z,�3u��y7�*Q��-�n��������4M�&��:
N�_f�Ӷ�pm"ٮ�X�<����wwz3p��Nga�edU�i*irP���:&���rx��ob<��3}��{F@ġieFw�b����&�Z�I�8m�&��;lэ���'F����F�Y��y͆�ɴ��(:�Aj�k1�oл6dybk�N��4k8�f��l����ns9	(̎���؃�ܓy�&�ɺ���$;rl�<��ӳU�"�Gy��=Y��ҁa��#�Df�&25foR�AgN��1��U��_F�a71Ý��c|P�N{c�k���e㜗4��ge{k[`�o.6�$�P��r��� r�#��w3݅q�������G`J!�@��������}r ��|��W�	{�OU�����8��0=�F��\O^o0v�ZX/ ��>�`�JnQ�N�Ve1���bޡ2�f��2�yH��E#�n�\M�,'���zl���,��Pv��]�L93�5��BL�%��GFRy����̬S0���P�K{�M�8]��V���M0�a��6��^�$}�i��+��Re_/��4u�.6��Q�7M�2�\O)�"�L���*^���:�q,�y�����X{���V\�[zn��'n!/ry���fv,l*N8���o�F@�x;�Viw��kk�B���nWv2U�Y��n�B�Е]����[����ַ�J���M��o<����ȍ-�jf����nڟr<���hԸ#�tsu\���b��/AM��#]M�ig;T��X��:�'0�&#�AF�6(8��%J���ж�̈��8<F��&��9����zld`l�JC�\͝�D�7�{Jn8���{�7jy�N�wkCV��r�tn+U�e��7���4b���*G\�0(��6�!�i����q�#�C���hЅs���Kp4�xD8�c��[fmLۘUر�.�v!C��pÙv7RX7�|T�������r7"KM�B���d@�0���y������ڥ#s���p�;T�2��n�6�	U^���pZ������9B$�5B�Ž�j�'p�{�Z�{Sp�x#Z�w�Jm�!Ō��\Rxu۔,Y��p����Vk�O:�<�̸��*��F�&�j�
�.og�<�>&L�f���)e9OO��P ڰ$�3k�wY=4tt]��s_C/i��8����v��Ե�ġ��fEpJ��]�o,�;
�Z�7��fC�7Ml�b|�-qS�&C�����}��e�Mй����x�P⹚�Rx��+U��eNq�V��/pN*�Ӵu�� {"���f�s�P#��,t�cY'{N�������y��٧�Ԛ�؈&J��.]2��� 0܊��ljZ�Jst�c�0őG����|WO���dS$'�kP��㹙8���Y��N\:M+Ĵ�DR�������&�˩c�����!��nճ��H��%��.`ڃA�mӒU��*	¤pm4hiR�o�V��w�)³L��g84w\�q�b)��-(�ٸ��O`do9,l]��N;!Y�]�ߛ�6��h�����g�#"܉
mc���%�	\�1�q���wv(�ٲ��bM���%9Æf�{B5�����Vo=r1�뛐���T���n�
O5��� �b��C������;��g��}۰���q�<#w��3:2�=߻��g�8��
�+0�[�K8bHhc�m�2�4�˚�3;�k�r��n�Ȭ[�U���,��*���}���ݡ��	�MR:n`���4�V�x�;%��1To"���$� l�L�2�S2Ң��B�p.:CsC/��Ksix
��*�cwQL�b�pk�b��5�j#tq�d	���`H-���3f凜9X���>��s�o`'R<��xI���|�X/1��L9���w�7�Ov٥L456@i�g콑ά�<Fތ��t�n�;��*x
n������$Ux�w�O���P���)�w��u��.1zK�$��R[؃�;��{2�5�1�ż�n����i���A~ݬPk�	��X876iu������^��%�'��&I�3�Y%m�I;Mdf�5�O2UH��oU;ЙZ�lS�bZ��Nj�ϻ�x�SxJ�Xұ0b��*������pdA��L��\d�;\�:3���U��:&&�SE=�ÛH�g܍l� KkK"v:��֥��l��_>�0n��ȱt�o���Є1
�'ȋ�j�z��RG�Z��W7$4x�gE���x�B�PF��72f�]@1�[�(]�­���GrY5�؊�N5���*�d�%�^��.���[�w6t웨wlU6sI�.�Ò��#�}����r+س�j��tF�������9��s���OT�TE�9�3��������d��@b���Lۥy�\W��`e�w\�|�<wt�gw\�6qj��̳+�{V,�y�]���3��H�/����$#8��u4"ךn�b��'(}�s�����t�;8J��Gs\���R��N��08��&v��t6c�����5r�v��:�g�N��8�n���7j�rvb�5��R�^��NΑ�k�I�F7�%peU
B"��!���O�S�H��q��oA6I;j��{�z���ŧ
X&QH�7&ف�A�"��"�5ȎSs^�a�g�mi�ŽJ�	����1I[ 1Jdâ`�M(��zX�6��M����e����niO!�Ȏ��D����j�-�np)�Fu=�8��7.1o]��=F�^��)Q�g��t9r��J��v���Y�0��q�̒3sB�H|��R��P��cn�I�2vcT�?gŞ��1�7���M�G8[-b]}�
��u��vnE_r�&��zb�ޡ�rv9�;���vs �e$,�_ٲ	L۬/*��ج�{wB]�6f�V���$� ���*�+�k&�Ŕ]{��/>���sh�P�V��n+̘mÜ ��z�c��db�� ��М7V�&��x~�1I�aӷ��ܘ
R1�BL����^�È�g' [�9�\[�>mCe%�8���c���&t����*伬C;�;�[7����T�3X��P�۳{Q�4��u͆3t�[إ��74�F�7n�Y"V�z�J�4 #�b�/
̓b[Y���cF�@K[�0fcYwi"-M{�����P_�����*MVB
n�b����ƛ�a3;Cټ�������^IfA:mS��6�ܲ���:5�)ls�R���[v���rM˚L35IRvNA{w����H�<�٦��<�7�ĺ�iN�1�5��Ң\����ϝ�z'*2���3��.�6�3^�wyX%L��Cۚ7]Òl�nd�C��D-�,^̊fI�AQ��1Q̽�m�� [!R}b�	6PE�y\!l?<�m�i&�ү\@'َս��y�54��nL���Q㧪�+��x��`��5���dw�?dt�&���թp�G �ȱ��)���i���A���X�w7fNy���]��
���;JU��b�gc�
��yΏ#1&q2B�����7-���M�x� �1r���C8��CP��l+��&(��L�\gc��1��@�W���6^ѽt��(�nK�ސ��QR�ŧ'_-���n���A��j!���&]8j� :�X�ثf���C&@�zޜa6���m��f7gUe�X��&[X I3T-��i�b:l�n�(#�ޅaٙwCTO	�֐G3$�:�s(���F!���3�B�d��us���Շ-k[�ʈ�,wc���թ�4=)T�+ݱ���{Nh4�6�E�ׁN�GM�ԛ�vgn2�x!�A��w��IH��{�z����˺2&�d�U�Ej-�XGp7Ahi�ך&�3P��X]���r���%�KH1O-��.�Y�xu&s>3�7�m9E�2��!��Ԋ�R��J]��o`yv�}�G/�%��hs<��Vy���k�R/�/�A���#�O��c��&���M���smH7��s#�@�Q3C�
������<%�����$�u`�X��#{��#����}ix73�\7��[C^J�r�Az�[���2(1�5�dx��ݕ��=*w�)�!�;*����se�f`9�r�n�`����Ky�ob/):-\ҕ<����qP*��&��ќ�fF�f5.Q-���:,ى1�X�&juk��ݙֱƫ�c�a��ꂹ��\eH�Y����N��	ŋ-�&�=���gi�p���-�`�Лѷs��7E�ޕ�}�*\�F�/���9�7�a���AW1B�5N�)�Z�5��i�,j�Shm#HX6ix��kź�M�	b,l廆Y9(y�`�Y�� ݫ7ݺ� �i��^�v5�ɰ�qG�s��n���cw��ٲ�H̺6�jr�v�y�	�w95��_9��nR-�H0�x����K#�ҋ�s���\6�f܆�S)���\�u���mϛ����]Q<�
��ǉ�Ҏ�S�f�Ԝu,�,ɺ0=(]Y�B���ų���d���j|'����:��9yz(�r�ر:�����c]K�4�xo*���.4!u�3p�Cͼ���ftKU"�rμs]�q*z�ՂZ�!��yW�d9�Ej�g!칻wg"Ld^D�튯L��;�������fl���w�����V^5�(�:��F�2CLi�Tی&�J���P�;i��ї�U�m��q�M�6Kd�g'x<=�ggoQ�
'ݹ���|scc{�wu�P�s�7�jw<
;�J3���=�vK������1A���t�"�d�`Zܠ �+${�r�!.�j�A��^��o�w5���+��K��ǹl���5�1����ȶv�h-�8N��a`n2���U�YI���P�q��r�pל�h�M���`���K�r��,��@�%�c-MdX�a˩Yt^P�#X�{�-Zb9{�p!�cG��r�2��'.�0p���$�:�P�z1�AN.��"ø�i��S��}3ε��\��4,Q��f��*x�ݢ���0ȃ[��VB���8�G���-�y��u�6���Aw{`0
]��^׻5���u�-�ER�Xx\p��O(Ԩ��@4��L�@@��k���$��z�����ix����3���8�l�ыG���}]H`�y[$|	��zø��Y�5�����9��C�Hp�J6ק��e��r���=��q��$4���51L�'#H�YxP9�'3��>}�����*��wd\�m��mI�h�/.Hc���u�q�51���&v���W@x�P��	�6�\�0�Ӈ��3Jο���t��6h�n>�WV���IS�����ꮸ;4��r�v�X�8�r[�K-��t�C��8m\/�h�u�V����s%��ئ6���4:��o)j۝+�+�:4�w�*����}��h����8D�_0�����ڳL���R���vj=���A��5Ǽ�݊��(���ڵض�4Q�[��]�0��OT���N��3~�Ѯ���u��)��ۯ�#�pk���כѩ\����d �� �B�BE$�, AHBH���$"�R@
�%@�,��Y$����HT!B��	�E	
�! (I�d��BI%d P� �E�$P�$RB(,� !@�)$ ���� )$ �B��J�B	 ���$ ,��� J��@ XBAd`�Ad@�d�
$ ��$RBJ�$�P���$��(Ad!��,$��BE!"��)���"��"��RV+	 ��,	$XXH-BJ�@P�,�B(d����J�B�B�BJ�E�AB�I$P_���BC�$ I���Կ2��L/��;Z���+/��a�y�[����YY�A4��2S�ͤufE��v�NV�s�w�M�f�fNi(�lx'��r�ױvZ=u���zƼ��Ch���
j˰|/V���L��i�[о&��jL"���[/LU[P�7yp�[���\|��V�0i�˛�{��3���5��qʹb�v�2��<���f�W�7�b�Wdmag�I�!�o�˵���g[�X��h1e�-�n�š�6d��ͬ�ݫ�C(���zw�%b����|�U���4"���^I�b��V)Ѻ˝;!i�/<=潎��~+��2�]�Ud�-;����� oG���7�܁7��P0T��u��0�ME��p�М>��<�Hƪ�/)�^Qd�-㠛�hZ2�w1*4[��"��.Y�%��_|���D;6����"O)Q���93�\N�\��qa���dV-{��ī�i�;���Ux��U�'݌�����E�
U�wa�o��V�=<�A�֘����*�'.@1hSiRK��ۦ��3mY53��P�D��P]��Ⱥ����n�N�91�J7q֛[2����_P�t��7?�����ל��ەs�]U�d���ͻfc�K����!j�^�E�̱�=�{���#��Q�0��O�a͇�)r���WJD:��<���K�&���j�(=B�K2��Q�G�K#Ów]�e�8i((XY�mkV<�[%�g+Rҹ�+,�sw�4��f�R�.��ѫu�M��/̚a��S�v"8�g��7��|��	7v��h�W�P|�:K5�&���I
�3F�Ya���X�hy�U�,y����U�{�Qǧ$\�Wk�d������r���t�j�I�E�Zo��{�M��{�`O�1_�/��㞚[Sz;b^�PĚ���=�A��9��6a��{,).�Vn6�u�k�Wv�������C=����VLp��U�P�1�M�-�e��v<�1iY| �k^�EF��G���r�]�\�b�%c���ܤOD5����+n�=��)�7ng�A�$��<��Ȏ֝���y64w���&�aS\���LʕQ�{)���Gt�:��:�D������X�+�鹨Z>�Yz�E�2��d��)"�a�ڏ ܓ,�T9`Z���<�O�`�j�E�u����>r-�l��Z�ǳ}���u�u	JsE��4�*�k�2���§ZJ���cki� �oK�$
��[|zp�T��<u������s�
��՚����/N�ֺ�m�w	�]��ϛ.����.�o�I�-uuY�`r�v��S�/�AM��5:�o���r��03�T
���ƭ��rV�
6��oz���rnLnK�T~��nf;ݧ21<_mO�zOP���Kg���[������7O:�
Űnc2�ޝ2�J���+�{\��V�d���Q�A^�bU��h��YLJ5Iμ<s�h�Q�ӕ��*#�VG,����$�'�v�>g5�L�sAW�?6US��F��c+��߆���A-Im�ͪ��Ů���v�[�v7I�7�7[���!��vt���2F�q�Ol��ڱ��>W&�N`��6�������=.0��lt:��e^�˥��\yzw6�Z+M{o6z�JHH��Buq7��k���;��y����`�S
�c��me�����^��#c���c��Mv���gv�AB�����}'&n&:D#��ض�x���,��H<q]�c��Y���pɬ�܆0�V�F�^�Xy�T'a�A���׊)0o��=m���M�U���	����I�'�y4=�^��!N�*Ζ\9y��3���w�{)��gox���Wæ�w5��W|1������CU^��Vp�t?d�������>�������E�䤷՝�b�^X���`ju-��꾧��	���2�r�$��=����oSޤC̺;��/���`�)���`*!�����x�!C��H�4�3�
����N�;b�3G9 ������p����l�Wc�y��྾���}�+�3&�`Y�V�w��ҳ��Nv�c�J�H .K�9[V)M=���4��P� ����!3u�,Zo0un-Wge���>3�3�[�!L~7��e�Ŷ/wb���L��Q�̓+�7�g����眆�k=���͗b:f��"�)ǵk��`��C9����m�����J<oN���R�"ee���#�U�7��7V.��EoN������ڕim��FA�`�&�W����D�yW��=���L��y9h+�pp�t
�w�m��2$Ĕ���d=u��j�Ϭ5ϏK������5�f���[Ȱ�J�Ǵh;�+���IK��ɹ��H�V`ݘ�L��s����{�A]Q�2��K���T�>#|�&���\v������^/��4��6��D�7�򃬕�f-�����:��^���DK9K%x����o�2�{�1�)�����hk��\4p��N��\�_���2�ɗ&<IgA�����'�p�d�e�gd��`��k�,�1�z��@����ܓ��W��t-����b��["�<#}�"�}�V�4�<)�Q�ic�����7m�zQ24�sݷ��H8&I�w�d�G���.E�}���� ]-���Mo�^���fC��=���p5#6](�xD1⼦ԇ=聆�&����Δ��xz�6��V�oP��9���r����;4,�1�-���ƪhѷ��,1�IC�o��Pa��|3ej���<�h$�����b��ۚ:*�z������MH��ɽ5�"�O�ߍ�e�8��X��=�
�h4�U���~��	���f!k���nn���Şu��ܝ��)�h��9�%���%�y���2mҖh
�K��n��OU6O{T���h��Q��L�2Z�ܳł�z�8�Y�J�,�;"�,��~���\\��SCB�R�zp<R'�������'V�7���n]����=s��r,Yw�ݞ"!�EU�z�Ô�J�#������T:My��l��۪�� ��Q)S���q�حf��d/Z�侥rK}ar=�y�zcV)�sz��"0K1+0��9�3i���=����n�����#¬�V�CN�]���Y)3!`M�n�<�}A���|��oy�1	ܷw�/!�>��̍wq����U���������1�wC;�@�l�{��xt�$�F*�1co��Y!}���3FX!��0�ia�5u��>��!�|([3�L�}1R�şt�f�W 4�#�� bP�.}��Jۢ�3U̯ٗ0�����Ϫs؄��Of�Nu��`/Ҏj@i���(�˪�G��^��-A�zڇA��`�{������{dR���&��&p6�Y��'w=N
׌��$Eu��we�KN-�-�mg�G��fmW��5mmA{z�nыؔ�Ҏ�y\�ŋ�����w��)�Q�������`��=����j�
�����I,��c��Fm�G���>��l��_iQCӕ�W���LDƥӏG���;ُ��Ѝ�*⦯k�m��5��(LB���_��2[B�9�{����'����;��������S�&ݫ����q��X�qXt�Ō��!��;�^�|3^�_%������x�4��]�1o"M�{|x���2)꺽�K�*a�E(r�XP]�Tb��_Z��[������KE�κ0�EG��r]���w3��ter٪_v�/ZU�Ti�!�t>Eu�.L�yIզMȲ��t�~9�^Tl��{W5J�?A����mӶ�f��d���@���OY����Ϝ*z��y��;�c���]��Yy\a}٥�v���lȎ�:E�L�ѻ��n#��CK`ܓ�=��"�e$�s��n�����T@�fg��s��Fe�wI�׳����d�D'w6����4�qB
�|��ʚ(+��������$��B5m}��MY=����p���Yv�<�Z��!�G8�;�|�w~TI�p4zw�j��,@�
��ib��n�LљBI�&��xw6�千ؙ�"i�I���BR�{x�T ��E9���Ӳ�4��n�������-K׸�a�3{����7�����E0�Mf���K�d�K(�e�V����{��B\sʔ'�1����b��&G6ը��<�S�鞄��q��a��(>�tMZW�}���r�s�)��	�*J�P�I٘78dǇ6VW��X{�[���՜�^n��H��BB��c�i�$�yw�1h�"���̪���D@2e����YY��j��Z����O;B����E�W����������Wp���!�(�r�f���F��<�m����s�A�sw6D���[���G�,��qP����F�meuL� �E�x�������ae ���^����>"�B ��.��θo����,v8\�Y���XGݏ W�J���W�twK�_t�DzfM=k4Ww��9��w�>Ҵy`�֏�$dA���m�̸6��r����+�[�M� oosw[�"ռ�ҵ�*<�G����J�W�,/�8r���<�&h���5^s��+98��� �q���.� a���r��)��k��m����)0��l�F
Y�+Z����T�I��\�� !6�^1	��['���	.]���͖��v��j��~TУ��u�U
�IV,A�U�uGyr8�%rS5*u�s��:�_lY
�m���W�xx�K��,��kN9N�ӼM��6�2J]>�
�>��H5۽M�^;IїP��C��pf���c����2f���]��cGk��N*˾v(�~7N	�=r�~�z�1bu���[�5[:�޾R�#ǏU��ִ���ͽ�jj�ݑ���`��#<���W��P{ڔޔ3�����c�x;�Q{<�����ih'ս6����}୏�<n����dal�a��Uf���^�^y��1��{ۗѢ���z�5�e��d����[r�
׀�n��q�^*�����S�*a�=G,0bҭ�OOh=���+�h���{}ya� �>��mS��:���%�-i0-t���N���E�̖�b|�f[#Si��o<��d}���yuj DrR$�AM;�>V��ﯮu}#���� �N�����˼�#�����c��_��ou����ǜ��O5W9p���uAmiiy��^�%?f�{c�V����ڴ&H�nh���wo]��9qX�����.1zE;���,����<BŐw�վSY��do����8ѽ�Ỳ/��(��Bۇ(mx��ֲ���޿(��i�#m�Ka��y�sѹ��4=է�����Rheoms�r��{C������]���m|���Z3 �H2��O5u���Aj����>��l$eV�EJz�wz�%mQ&�_gL�@gcը���9su�g�{=7vW�x$��=���o��<���k���n��j3W�
y*�oBl�7��kU�Y�T�U��dN��C�����^�F�.ߖnAR�̫ݣYF7�](���ɽ����<����������v�oN}jJj�õ�p�:�kަ���@�����]�aEՇ�E��V��/u�I�xv�:;k����!r��o)�fv�*޶�.=H�~<t_qu`�����Q#R�oۋ`��[Dܹ����1���ʸ�MP�h˃/
�ł��zXB�K�!6U۷�2j	&-7*�;kZ����{�z�QE������c�K�F�/�f��cPׯ0Y�1Sd�8ޟ�X��t�[���k�+,�D# #�3���ğw�U�-�;}�o��S2���wQ6�r+�7�;m�����/�W�����D���V3�U�B���|�k�Xx�PN�+g��L��Vo��*�MSf;�8HMi,b�}�� 7��\ǈ��Wc�C�5b�
����
]XW4�VA���͈�-��9w+������o��{�P����D�M��ɻXm��o�U�Y�V����>NeX�@ڙ:��3$���S��U����1	�n��Lbj|]'$x=�NI�	�݆�����7u�kc��x"5�������n��;�����w{��
Ν6����z�����Q.��oR���.���쌘�c^�HM��Wwܼ��}.��Uf����Dx�����˵radYO2�w�d�+a;ˑv��R�(��aZ�!�n���dc5nU�(�YW':�)���W�9ez�LF�M��Z��I�ݵn��02�Y�� R��whϨ�eCz��E�<7�S{�붳Q�;��K8&�7	������/�>�!����ږ9P����Oˋi��З�Yƫ��g��uy��3U�[�}�R$L���������0���{��������v9��s���}-�6Z�O��W�����
�G�#�r�cw:��y1���%����8*�ko^�s�uޔV��C�H��M��� *7I��n��X��p�����s���q��q5x]y�x��[M;Y�L�`���`�2�3L����3�q$��x����]�t���wa]&�|��Z���yw��r�|��j�lQ-u����K�W��O�b�R�u������V�XW$o�9#��Ĭ�3l���Ŕ�q�u�Z.G�^��ԗ��l,"�Pq���i����/d��lM�;v_��}�{]�;		r�&�Qu�|d<'9���ސ��$Tު`��3�ţ�=�Ƕ!5]���P"����"�&䯙"���A*�}�Pmnu%��^%^��wpX��J��-�hW+���+��ȧf��E8_s<ww�Ux@��G�o�|�|>�<$�{���ګ��C�ִ�uuK�Z�Β���#9��=t%j6�N�k��z��K�ڳ��ŋ�׃���c	Zt���n��u�am<..C��</�*��Wv9˷7oA{�B��;q��v�\v��7Qn�\�n�[��ܫ��mӇYq��ݻm،�W�\�(��/�uٮ�8�'�����eӜᣀ�y�l�7]��6���[ԁm艮��m�aMr��e�	{\��Wt��3n�أ�I���籞��n�ͣ�kι����]tuŀ�,����nݥ��ّ�Ʈ��W44kSAt���M�c���,l+{=[�/n���ۇ����L8]@g�z�q�ev��S��k/l��u���\���LQ�q��i�;bݜr�q�����c���nG.��n!u&2�ٹ3ԥxa�άOÝ�=*���ݽ�*E�|��$Km�l�k�Q�9�uvw	qk�ۮύã��qQ� �9�XíoD�:��{\�l���0p��
��ݦ�y����u�;s�|��Hܻ�ä۷׮�v�r��p6x-�c�N���kA����vi���j�a�Q�K��1Gl�W\��s��狵�w��<��u���C1�cm4���t�oe��n�7��d(w'`�0t��q��ܧm��{v�y��p��<]ȭy�1����\��W�l���ǛpER�G�j-dL�om�Y{d8�ga%�[�q�s�v��0v9��mr�+�j���s����§^�1un��c�M^t]v5+�7.�t�]���qg�	�Ӳ��-{�8�3ͮ���Fkzn���fp�.�/e�tu�uA���[��͚��piۧ<u�s����]ƹ�;���[Zx�:S�^�ٝ���n���..^�Xy�a��YwOgK6ހ�S9۬������jgv{�ư--z���U�ty�n�k	����۵��HrmYO�v�w+e��F���:�+<�hC<q�(��r�)��4v�y!��i�Vmd�����H�%'v�+����Sړ���{��l���g��J��E�6�v��{	�Ԟq�\�;V75��p�n�3�}��k��xgZt>�n[��`|�z�ѽ��pj�=;���[����p`���g	u����M���Y���@�2���pF���Ui��y��_lN�5���dX���N�vT����O&ٻ�˜l\�۞B�;	㮧s�s�nN�뗝vy��;�x�ԙ�v��n=���Q�5��u�v8n]��X��ݒ펹^]mۗ������{Kv9w<��,�1����(8F{E�1/6ǷR��n�Pqpgl4uv�:Qaz�l����k��q�x�-�Q�uvf�	s⮺�ش8��nv�,<CnV/$#����5f-�mU�4�5+��k����=v�c�8��Aɨ�ݞ���s�܍���v��]�[����03�f��<��:�B����;��p�x6��,��Ⓦ���JA�mcy�ɨ�ùu��@&�Z�^��U�VW������p��-��J��z8lkF�H���a��-�sz�C1�|h�:퓕�v9���xU��lTGT�:�[�Q��;lV�J۳�l��7T�n
CvzK��맒����q���h4nu�L�k��%�����w+n4�9^�cn{q�lǐ�WL�Jޢ䮞Q��+���.Imӎ2��[<�6ɸx|��=��v-=p7�-�0�5�w�F^OEm��pz�Ӵ��'�t�q����hį�e�ж�N����:s��/T����;o9\�riCv9��;m���	���+1����j�	�ۭ��2��m8:�C��֌�F�7l�:��xxK��ӻ��v�ܭh�v�7O.��k����<B����{v4�a���7��.��k5������b��;]���1�xWiwAZu�"�8��Y�=�q\n=�.g�bц[(J�˸กӡط=���;R��*�u�9�J����W�s �7�m�\\l��$���f�G�nۃ�u��R��K!@a�O�f=��osby7\�NƯ�Sm�]qƖ�\�{@�ֳ�g�Gc��[wU�le��:���W�v�u�����y��'���l�k����>����5�n�.V7/3�^�����d�Y�te�B��':b1�Ͳ�ay����Y=��M�p붶鳎��֡��(T�mw��{Z+nk�vt�R�ݒz��>5Wn��l0C�Oqs��[8+�[/Nl�]i����f}b�7��Q�ۄ�'�VͶۏ��������lQ��e{��'��l.%����GK�\��g�����Q#7-�@1���d��P֙�x�*d�V</1u�:ñ�Z�h�Y�6���n���I��������z���]���/*��rz�ۮ�ɺ3�DY��&%��f۟m�o$�ƒ:��L�n�VÐ�@֭ۜ��&:#6㜇�:��x��`V.P%R��,�ta[�=��y�[�^����RvE�,��#��nxE::�^ѳ�rmnS��HdW��۴�lYvڝ�=�{6�W��.�n���ѷV ��u��[	�=6<\�\�;8	s� �9w\�2`�c�8�����㫎�\[�v�Y���3ͭ�V�m�������Z8J28ήN�Iy�	Hn�n�����'lF��mqf8�3�LRhf�m�v\:.�G6c��K�v���	ݜ��r�m�OQ�W�s�ի���=�H76H�&w��l�7/b�ª��h$�(�qc�C�Ft���Q���a2t-mu����o]���]��屲{f1������x^8p�����{<�nw���uh���M�U�Xv����nhw8�/���g�v\�Л��\c!��һ m�6n��q�.'�G ͎6�p��g�[�M�lE�m(�>�xv8k������6�X��m�$.܏��jݮ��O	$bzA0�t<�)��nP��x��<���4���}�5�2
\땞@J��b-�g��Ϡ 9۞۶׷3ǐo\[��:��i�I��K	�`^�ɴ��x��nF�\n�Ի�����7�����)O<����-��z�7�����㲶�j#4�/]k�Sl�4`%�۶;rgQ��ۙh�뮉ۚ�5v�����YkrFۯ��x��l��ً�u:�ej�h���u�n�`�'�n����Ѻ�d���q)��W�;n�;I�{�c�ծ��8��{=�[���r���^!�\gt��q:3��s��2��V�s�g/��nF9�H�w'bջ'n���T�vM��l�m����ᮜa�������*P<���'q�s���x] ����۝��[=��y���\Q�vv�hH��\[C��ɣ�:��0��v��smؘvBl��g�{Ԇ�O]���A{C��E��[��݊#�{r��M�;��03��q1�>*I�[D���2y�3�t�N���A�t�{.]��u<m�X�×����.얝a�۞|�r��9�.�q��n�F�G�ҕ���:ϒp.�t�g�q�nجOk%%L�MoP#���s\�&ݻ]��QfYY�ڶ�q�9�W{Ss�V]���p���z�cpt.Wf��_lO];�ov�-����K��x����eu�u��#��I�z��z��.��֡�t��W�O�uN�%��F�۰�F��P"��3���2d^ǰ�̼zx&�M�w�;��M���]��՞���n<���C.}s��7e�^��uG��z:ې;C��;v�a5���R��:����ps�9���&�ݸU��L�]��-%�l.���;��ݘs�m�n,�wI�������l�rݎѷ��[����GW���ntt>Χ�7��S���;֥Kn_^��۱�ݍ{n�ޑb�xȹ�Ý7n��EY�!��M��fG�i�ˍ������xO7���w���ݝ9�8|{<��)����ѧ����`��n��6Ѻ7mv{P\Z���*l
=�K�ǋ�Sm�ۀ�b9�:��n16B��gc���j}`��@�X��6'�۱q��9�=�˽�p�k�x�{rE�]����l��:a����:�;]�e�����<wXm�m�as�Ujsn��.W��ݯ*�����GeVێc����v��b�h7k��Rbz�N�>�@��$*f3����n6J�ķ�ɛ�gj�,5y8��[�ln)����v�6�עL�v�ݭ��u�p9�<�O	<Ӽm�!��gQ� 9�p��JN����&�P��ƛ4�n��v��[qj��]=d;	��m����G'��Rw]������H�����خ���hM���$�c��#��rm$i�0Y�۱�Ӟ�^u�vNN�W�ÃI��>���玶�4j��7�[�k�ۄ慡���ױ���d�W8v�b��G;$u���"���C�ˣ�U�㇁�ct���=��pgA�n(n��cQo/&�ip��*C�\��^&ף]���q"�j/j��xnq��^x�&v
��zԻX�#l�km n-]xǗ���ٷ&v�t�J����c��ݛ���5�$��ѱwf�h,Ϸb��`��Yl���u�c[n[����Ó�ӄ��s�h���tk\gD�p�hn��j����c%r�a{;��F�(\�#�T���'�m��x��Su6�nΐ��k�9N۶�Qݧ5�g�	��3�Y�OE��[=����2����\�%��Gm�{Dv�Y��x�n��r۲���h��qy�r���ty�*�۞ѵ�0l�m��N��(��sn�e��w���]��5)CW��b���{k�	k���]�k�͖���G�4����i�N��[�Nvpe#�o<k�g�+�:�@��a�⌰��EݝHl��b{\�3v��vk��w��v�m�uF�bR�s3��R!h�J�Q�X�[J�l+A�8aE���.f3Z��V�E�-���#��b��m��UJ�e�m���cPq�-�A*+X�m�EFҩB��h�)Um���T�Es�ԱUPQe"�UQ��[QmQE�����FƔmh�-�U(�����ˊ�څ�U�J�+[j�ڠ�h�Z����\[*�h+UQ�kRѴ�j[m�X�m*ZԴDQLf1�bTV����6�UV-�����2�kmnS2¶�cn8嵍F��EJ �V��T�j+ik)U���ڌ��-KJ̦cB����jJ�[TTJ#��+[�6QR�kbڦ2�Uj2ډh+h���*�j+*��Z6"�Q�)m-��`�P�m�E-*j%-lh#U�l�AF�X,�*آfLP�
�PYmUR�
-�a��eFRƴ
���[R�m��5�FV#D��%���UZ�F*��j���j�c\�ԢH��cDU-vI$��)]]4�'`��e��ݐ�8�,G8���lG���w��?8�A���7<�Y�h;N ꧞,�ה�
�1��'���ƻ�r��81��'��P��:j���m�����ێ޹3����6��C�kӳc�9��z.�˳��û`{m�j�q�^x��|�(���Ə%m�l��ٲ��>Ŭ�{�.܁��-mɹM;�#�KDM�K�6�w]95]v�2r�rGv�kz���ܦK�zu��wf�y#�yݞ�5`�m�q<�\X8_c�*[�k�oA�vF}��e����{����a��D7�u��1�['���=�Y��a1�l��/�9��c��{iq��/==�I��=+�a�׎�v7�[�d��g���zq�dX8ޅ^��]��uH��9ɺ6�
b�6�<���8*��qr�g��kk��m�Y���]��Ѯ��O-��;�q�ێ 瘺}�.���s�7���]��*������U')�MM�]�3�>�rbMB83�z��em` �tq�	#u���x{\n�m��p�3=9�s��<����0i��n�ۧm�����ۖ�zt��]�u��v��ZGq��{]Dg�=����zCv�縹tpdg�ˋ���։ڬ8�)��[O#:�[ю�9�eǭ���g���/n��Y�%�Ĝ�s��Y�۝�Yσú:�2�Fp�-�oJa�:Ӏ�'i��Ѓ�[=���1`r�8;s�jDԑ�W����۫��;��$q�,�\m��mlj��s�۵��k��q��.y7�1�Ѹx�Ð���e����T��m��i�[���plK���p���W��!�nն燣�!X���9pgsv��D�M�l`QB�h�{�Y��]�d� �v�dٻ���ʔcXnۑ�b�4m�wk��үM����۰8�m���β�n}Vݜ౅狝������]j75��Dњ��Y�U�\pJ�3�����l1�ա�-3-fո����.����3UL��Tr��1�&�RʗfKk
�,�P�=��1��0>0���عr��s˘��.3m�����)j�D�Y�71�6����p���v|x|�*��{(�=���m���<!ȸLa�Sex\��*��{q���������ۜĊ%E�z��`�A��5 ��$O���sw�Xg�s��,��M��X����J�j�h�"���f]����Q;�`��������m�����	$�����sqw�߶Vg�Q��k�'�Kb>p�\�a��x�u�6 �R"1�leϱq]S/�r o;�� X�sq�n�lr��\��Hs�b���^�]\:�|�J+��Y$���kt�H#{��0}�N��\ �y�tl��#�6b���bO[>$ {����mi~��ى@c��@$��t�'7���kG%�S��Ȉ�H+z뒷dI�ݷ���w�g����=�Ǻ�/nky!�I'��>S10C&X�ȉ'o����u$@����Ts��1}��ߎuz�q,�x����J�DϮ��D�R'�s�ٮɓWU��)��u�\߲u���Ζ�w
���i�<ذK=@"�}kov�}\���ߌ��k23�]
�ڢ2����+x���Q�FyU-w�[�θ 7�� ��ի ����E���os�WՀ�aL�!���Y�t�/{i]����ffW���0���[�	��/�H=���6DN?��N���]O�}X�=�R�#Jt�����"�Fd��qH�������Ϧ�As�2��r��.UE��z�E��z�k#��w��w�Eܲ [�R�~$�fO��*s�dl{�z� [�A2@�J5�..�nv�'3�4u�9�}k�K#]����q�Ap�`p��8��D���ܥj��f>��[��x��Z�{Z�SL�� Fv���VzG�f�nFڲ©�Zv��I�6=�K�G�S�֪$ �����'�O�x���_��Zx�f r�^ gڨ��T�$�'����$�D���s����t�N��dr�9����;o��7�rRޮ�IKw�B�a�m�:�Y���e2
��B���]�����|k���D�S���$��vڨ� ̟qj¯Հ�LL̍8l˿�>v��a�nLR�N��
��q X�u��x�_�Jm U�Z��+aG�7
G/�sw�{ϲӱ �O=t�v�f]LR/o]���"=��� �}:��8�z2�/���ɗ�9^��S��.3ӳ�MY8[�C�L��G=�mz�F?~��Y�V�3w�~��֮ȃ��{�� �>�dE�)��o�'��B��H/zn�6M����`��aS�]�^����}�b�+6mD@ ��� �$��K i/�������wH�L�m�/�w�Z 4箙 �����G^��j� �d�d c��D]zm9��(Nd��=�v����9�;�n.n7�n�>.{:�����vڎ���g2ޥO�/t"��x�����c^���@ݝk�|�zfR=hҬI�}�����3��P�����)�ӎ�}�LN�����k�;�m��$<M�������OĒT��T��o=��%K�{猓QbE� <������jɪ�/�۞_���~���2���k���va��mj�3x`:�;;>����a�),|�����s˺��pv��wi�R  ��m]��\�\[6^|�yi3�Z���]�v�,Dۍ$܂̀��F�Èe�R��/++ޭ�|V >�t�ݶ�Y�����w>�9X�w��r�p�`pѴ�M��N���H�ᶷ�1][�/� ��n�D�vڿ����		,��m
W�J�_p���?n�~�@���H �3}��"� Ǟ�.�x���������䳽<��n"��Q�ʥ�� 3��`�����(�����$ǻ�j���=Σ�}����<H���S��ǵ*�!fq�ܨ{���|#�׺��W}��gx5|����ŗw��x�v�^ōŶ��h���O���l���c'^�h�`7���m�p�7E�m�'c<'���lx	�mq�1=��=�Ac���; s�����w�aN�ݷawI��z��É�������y��4]g��85�c���,�%�9n�����Z�6�8�ٮ���kKWX]pL�jiȟS[�q7�.�]	��U�������ԇ1,Qכι�8n��m\�OGݛ�nW	h��Al\0�u�n("c�	sqæ��ד3���z]�5[�h��E���妜ֵ�&c���i�J@ ��j� >�y�wh=.k�ϯ5k�w��@4c�V�y�� ���_����s`z�{}��/B8�� {;m]�0��iY�˱����]Ӯl�;jB���Z-�,*�yܫ@ C���#D��H<~�w׊]�I:���/�E$���v��ꑸ�jY$9��E�|�]�- �t�XG��:���0;[s>�}м�	]����]�X�[��		,�$e
X���u`|���m��X��W�rhJw�œ|��{�����cd�Bd��wg/����r(�)���7�/4dby�q�\A���ږ�OF]��������l����;��Z�@ ���_����H<I���K���W�_�@���{��U����a��Zƺ�$�DM�e�j�Hꊯ��ב���j��˪�qc���cCot~�7O<|�:�,˭��J�<j�`�̩N	D��xZI��}��"W��l�w�O�8c���g}������Ž߃��ڛ A��u��輊�ǫ�[퍴����c}��7jBɍ(Z-�,��9զmybP��j}�� ���X0=��P{�I�̳�a@$�\������R7G,&U��['��$ wzv/�#iǾ���� ��Q���|ǽձj�������擹]j����W.�N
�aW��z5F�Wh�ӓ��#�p�5�o7����_�[C�)��z�"��R ��{�UD��4�ôг�V���&����$/�����n"�"�-�6�g�ד��T�}�tw��@ �����7��*"���/Տ8����U�`0S̶ӈsq����@|���bŢRG���G��0�o����꽝��k_�Vz��yG��vM�q�uk���lW>,��>�8d���;��^
�B��U���W��pH���7@ >7��/����B�����~&n#Ǻ��n����:�R�gV��_�#^w>^׋ҧ��R�dZ[�l��ꐳ
�r6���D�Ko:����̐�Q�S~�q7��-Y����
�X�.�M�8^���:uvujmY=��g-�������nN�	�q���	�3����M5.Y.VG"���I ���]� -y���n���M��+�4�F���7@ �����f��	����
*���y\\]lz�?Ht�� ��ظ�@$k��vA�vV�^~
�TԦ��@wNZ�*����=�5�����l �FO}�;��u�L�G�h�I|���D�����3|�(����Af'4�k����޽��gj��$o�� i}έ ;y�.h��P��� ���ҤFG�^��ޙ��(��]�=7h=cP�.�$#�o �b��n�8�����t��<�*0��7x�����Ě-de"j�=Z!��I�Br���Z�PK��Lo��{n}{�vMYv�@|c��D�Iy���J�+�y�����DH��c��7M���W`|r͘oX�e��X-���_�����;\]�{ߦX�j&!��UG�9��Շ� �s�M�$ǝN+�}+�3!x.��s��k�"#9�a��Ö�P�̸�*̀���_$K�}y��7{Wz�r�h�Wٳ�.��t��>����eY�
󥚦T8P�I",�n�i�gK��	��/q��W�t��|I&�ޭ@�u8��r�9P�9q,�{&���9ٯ_�r=�>A�u�Z ��� ��oN���Y�f)|=�V]�~�K�s#i�9�H�K�7:v*+���g��V�>���� ��f�I$���m��C�0�v��צts�>�b�0���G��#P>�6�����z��n2�/�A�|s�&��,y5&��Lo��7K����}�C*f��y|���]���u���M���e�h뎰v�4�L�]m׶�1�'��]���7V9CGmټ�bK�N�8����灂42�ׂ�0<���'CTD��w�y[��=x�`���xg��O[Ř8�ʖ��8�йӠ����'8����T7����xv�q��W<���|��|n�:v�;v,�Y+9�jp��HQdj#4���v��	\��1lƁ�����CǦ۷[��<Y�q[g���c]��Ķ������nܚ��0�9����v {e�"ro,y���ب�g2� \�cI?vfԍ"�0���Y5:i�L�~�[%o�j|y��w}�gY_ �� ���Iϖv��*3I��#%CS32L���S��L �N�� :���V{q��QqZ�u��|gul]����	db��V�[�8~�򱚑>QӤ���;h �;¯{}YdH���4M�/ĸ���1�.�nU�� �=�z�w��t��W]g��Jۚn�D	"�ձj�Fy��gGe��r�o���@�xI?H�e7-�"[�z`^{2�n3��=�i����9lm�f���~�����>��Ar�%��I"o6a�a"P���v�@FqJ���5���$Jg��*-9��
�L�9�H=Ϯ�v|<�:`��6�8�6�9���o�Â�B��y@�}�+��x��um�j�^<y�X<w�y�G���X�3�)��s�n�-C��+�&G7��S$�R��ػA�x���=�s�}/1���%����b̀\��� �7^��`3�USm��ԉK;+�$�vN6-.SN������lڦ�_^�yÇn�����inϢ��X�kj/�S}�'���& �Z��%fP�B� "�Գ��q hv��J��os9Ә��E�� {v���0;[�Mخ�{�o�����cnWi�G<�ۥ���t��,q%Z^P��Md��C7wI�i�cHY�ɨ�ힿ��	c}��tI�ޜ�11]]�� g����S�c$��24Ar�c]N�_�ѵW�{�oC]~�u��+" =�]h�X�kt��oE��>�?��g����A��bs(sw�{�n�`��t�ڭ^�mfp^Zڶ�\boU�ۚ��`��K��lVjM�sN+��VOAN��5�>��W[�Ӯn�AA=��j�%]��zh�=�&���7�#�sU�5x'݋�����\��Fiߦ�AV�"!,w##c�ڏ��,算o=����kj/�Q���j�N��"	��v �����j.%�SE��+U���X A�倣r�G�V�
����s�a{��ݗu�h��Xz-'�e�;�ܜ� *C�-ɋ&]�M1'B�v;�������xU�̾Xd6A�uA`�ȥoT���ݑ�~��)��mo�w��'�A��=����ǧ%k����^�^�{��/u�.Lne��bZu��5z�e5��R��[4M�5��dEw���2��*}r�]Z���ך[�z�	�z�t�A�U}�>��B��ƀ��o_ X#���j�'ح�1��n9�왝X��.���c�Y:�@E���dQ�\ݑ^o��F�tV&g��Gd�P�Q�V(KR��ה>4^P�J�ێ�Φ���u�Q%��Ru��'�]$M���!Gwٚ��o�������N���;��aνάڋ\Ļ�.�6Vn�4s�Vu�r�ӆޱ�qt�]�7�8�~Օ��y�#P�
eQ1��&H's�3����W,��{��yr��P�U�����zf3�fq�
z��k����mj˛��I��x���Rgw��X��,�^do�\�ݼ�P��n>-�A}�$g;7n�c{"��N<8p�(�A:{:Fj�@�Ԡ-EYm�F���TH�����]%�5���Z�(Z�ʣ)[m����*��E�D��E��KB���h�"�HT����mel�2ՙZ�,�ѵ���e*Z�,D��5mIDs�R���)PR����kh2�R£iIPPYZ�q.YU-l1�Qh�P�T���(T*�*�+E�0��-�[���D�QE%�YiA-m�kmm�Z+*("����F�)jZ���ڨ�ҭ��m���k%h�)VՕF֕X�E-+[F���mTm�(�[mh�me��
��j�kcl(��[V),b�J2V��X5-[V���J�F��-A+Ecm��T�)kV�(Ū[EeT��+Fі��P�0Dm��J�ԕ
�B�([%��*���

����YZ�Z�J�,R�K[J"�UQmV�Th��E-��F�H�e��[X�Y-�-e�jX�)V���Q�kZZU����KKm������/b���7v�.� ��n��6HB"$M��W:��F�Oxxt�@ONYq y�ku���=ձ�=<�;�υ�H�wjť�q�p&�4Փ�~�Y�0���̛��׾*��i �{��|3�[-n=�q^q5}����PO�a�;��[�nz��S��q�[\s��3V8▮��ˎ\��_���}4i�C$�"�AV��Z���� |%���d�+���S����k���@���H��y2��r�p+���V�^�g�ٱz��g�$��n� |g��-Y,���{3��>'�{�=���#�e9q
ݤk:�H ^��_� �퉉�1�mGT�؎@y���� 3�[�s��
�.�C����>��NO�`s�
��c� wkb�,=;�%}՞''pJbW��u5��=���!���7�z�I3~�I8�I&�PYy�s�e�Uv�߶��d{�l�S�W�]��kt���e2B26�W�s��Z� �{֝�SJ��o�52�? �Ԫ� E��:�.1�[��F˓|,�k��R�mq׶�nmѭ���y����u[s"�B��O�4����2ExxN޺`��N�E��y݃"sަ�����}���e ���ؿ���\j�. L�H�-}jl�;�Wq}�yuG<x���ձw�D���b�'rV�"Rz޻���|��Ǆ���.F+�ݵ�v;y�E�m��S��{%�����4 >�����L��	����_�_6���\o�) ��s�`�_���,���7r�{s۳�Iomxݤ�A ��C��uu���C��Im��+�>�n�������`$��ݮŢJ���AG��[�]zP�L�T�
���h�����T|}7R��~l_3�D5:�o/X��{�y4g��۷���LL�]UÝ_��$%��`8�-�D7��vn�6�I�;.أ[s�v9p��k��l`��<�ێ���O=���pF�[6�z�ׯi��ub�r��.���S�qqh��B�n�c���tn�-��7:�29��3��6�T6:Zҳ�8���C�^4h����&���N���籱cDn�ݥ݊nVuu�q��=�:��V��=k��2K�����p<f�9��-u��Z�^�͊ru�Z��MǮkef��z�g�����S�D
b[$W\�tT_�"0��͈�y.��%�w�|5��k{k��� ?w���8�G���4Թ%�q|SW��_��Բ:]��y^���n�� 1�y�E��������׷A�z㕅s��KP!�J�n�i� B}/p�@�2��s��~��2x��� �7����]F)�Hc���Wf���̇�+�� ����b���I�|gulA���j��Z�S�d9���b9���{ �T�A��X��I�6��x�e߹(	 �o�N�M�.�v畿�؈y\�_aSk�b�;!@P��+�׊==�/c�}l�y���³38ZJ�2�r[�mU������~$�i��R��>ѓ%���Ր 1��� ��T�r������O���B���=��Ό�w��ɻ�^�O���W�"MzJ�<�
������ɳ9G��s��_mfY��1�[̘�U���.��3�;:oE&�j�����K3e�~N����_  Fw�ػ @�Q���!�+�{��Pn���#24�ڦ�[$����- �����|na� ��[� 3��-XW=q�T� s�e�[��wyV�>���"_:R =�[f{'��1z,x�����KrYt��3Ʈ������=��ǷO��s��6݁�F�N��A眨���^��egr��	p'P�W̰[EfR1E�8z��A�ص�
=r'kٶ������!��ħ3��r<�SqH ��صa��{�Z��6�Ϗez��z�@�V��c��(P���'2�5�빰3��Uՙ�^o �=� @_��.�|�>�v���
���]��+w�['�&mHh!�FE�W]ZlZA%�,���"H:> ��ڳ9�FXѭ�a�"�wC��*(��'�Čݍ�4;�廓/����;�t���r62�����Ig+�e���o�| ��ؿ��|���wgD�y�6���ӣ`*j���Un����_�P:jn*",���� c}��_G�"�����ձQj���D���+"(��S`Dhv��jڃsn=�ҟGD�]h�G��uh���A���+�V�IES���CH!�Hx]�rrD
]u��3;��瞋D��kg����������Ҙ�`���{��-XG���@��su�Zo���SX=�l��E| F��v��+ɇ0�71n4<"S��ibN��lZC�@s�k�@ 1����K' �y�b�r�����Ղs��
0��P��8�]�� �C<��" ų�3�~���x�y�E���7H�����A���b�Tq{xv7t}��C�l�D�%�,uh"7�n�v�lT�k�u��蠨���S��z<���*�Z��?h�����۴p�n�os]L�)�#��Б�Y�p�9Ԉ�l�+kN����I5��m����y寺���Fk1�UՑ�C[� >���Z�<�����'�0�"5&�<��cy������ߝ�>��#rG�L`0��FmXsѕN�t���yl`���e��n??�_��DbP���m)�"43�� ��$�ܫ��ceZ�Z�@�.��s&	�rC�L5v����E��.��rx��)� �����DR;z�-XPI������7���>���W�jHȁ8I.Y䞶p$�Y�h�a/c�$i�qeǫ���cy��)gt�Z�϶�(`L��C����R�{W�l@|���oml]��#_���"7F~v�t�|L�$�w�x� �������o�D�'�-��ŕ��w������#���iY#_o;_X�S]D�&bJW>���tqm���]R�ug��;[���}�l�k�B���%c��1z��V��V�������MW��ϡ y�]��h�sJ�Z���ez�2m$p;�[��(�ռv;e���)ۀ��1�\�u)�����p6�cg���y����pjm�P�ն�u����s���3�c�5�H�y�;t�p�^u[HuF��Y9a��셞88.=�1n���`�����a��uل�&��ݟ]�|u˝�<�]w>����ʹk�kZ���u���:��[�����%nQz�x���]�PZ`��\Zw]]���qP��v����9����$?����N��cn�������3sUW���_-@����wG�wc�wW>)U�nu��#��b���~��� s�e��}jn#����֯9��� g��.��_�������T���o M�2`qF\5v��ڸ��> <v���A+��bi��ow�=m���;��k���sd̸���Q�|e�����g^�h�o8*D 7��vA����l��;��ut�@|Vet_�w�B��19�9��8�V�#C<�Uן0.��W^���|�Y@cy���0���n�������q�]F����V��2��]i:�n��������*f��D����e���L̷
��u;�� �5�ZN� ��n�|�Qoo��tN��.�>�;���Q��Jr4K�K=���"wWU{�n�ݛ~��wm�Q'6��s��֮�9��{�m���njsW�%�u �̍�9��/�)���;K-*�7|Q7q6���Y�����Q�o�u� ��w����]�&�'\[W7Ny�����:zߵ��H�s
��~�b 43�H|{��^�青I|�$����.� ��n�@$߳$�a\5v��� j���{�� ���; .h� ����CG��F@f�w $���:4��ڒ-��0��b{���Ê@$����:�lTz�YWH	��i��: ==��/&���dͷ��/x����nD7q)�H�qmf�_q����Vq�Y��.�qҶ�������!�)�̡�p{_]�� �<8�� K:v+��m��i��D��Oܙ5;6�iD�)���\ZD���VW�k�.�7�}^wړ� �`� �=�� g�=�S�z.K��&���GN��S�jG	�Qqh�~� ;�ڨ���&Z����ԏ��/tm���H_}Z2���ͼ����n�(4#��B�W�xj���|�Yu�?'��]��ҊA��s�Gn�I/��k�Y��~xq��n�;���H�s�����g�}��UM�Q_} �ګH�F���y�km��/b(�t�2�%�9pH�ZG{n�-�s�[�DJ����l��x�x{c�=ݵv@�����s2�[��D�W�j�s\����5��+۷3��J�v��$�rgyzgx�h��L����RFa)�	sܴ�ʢ5D�MT�$U;� �
�}8h.G�|�/7j����m�L r�������g��^�Ϻ\���A �iw�H�D���t ;��<��(��W��~IOoT��X,��$Y���݋ 5�[���M�]��6�I� ��.�P6{��-/�M�d�bd&�77�^/SH.`�wyVI �yV���hp߽.�呾��>��`���:yxd:�������CR�=Q���{�˞p��B��Z�v��GOl��o��Ȯ=��|$�>-��w�m�����t�5�sNT�&���^	$��~L���[�f}�t�����A�8����`�(~��T-�W����21�4�.F�l��f�y�ug��u�ܴ�� �w]������"��g5|o��� �=�<U��}�����Q?_K���II4{���s��l�� Ԩ�j͇<8����L��륷�Z�4I�L�?��6�l )���3������[p$ʇ7a��v�@��)H$ SQZ�:O8콴���TE��8q=�����*�*�۲o���W�Av�������""=��V<�
yZ^{�a��W��x��E�B��:/|�$'�r���!�Ȱ�hHy9���������vR�S�X}����KG��I�ܦ(mtK�.VJ�i^T�}���أ@b RV��`��aMݸ&����C����6H�NXF�7���ºAX�=��c�gq8��%�m�嶝ݮA&��ph���Q�0�c�i��%�;�G��t��ѝI^��5��ŕ��5\:a����Db��������Ym�����-�/]�Ϋ���7[���F�`G����L����V�Ρ3�� :y�	��X��v)��nh`e��b*�Ł|���r{������솅�1o���Qdڼ�V1����Б%]�tm�������Y*Y����Ǹ�V����v��3V�dD�ʒ�6U�O]����s*ڄ�5�y%}3wD��^]���-O6ܵH������K�|1�rѢ>������L�{��n���ܢ6!�-:n�5�*�.P��ug��	�ʜ��!������Ƴ/,�''��0֕Z}��趵�*��R5��o�onF��{�Ѿ��4������-w�a�&*�3���nj,6�gU��epT�I�ݻ�=2?24/�����w���Ӫ��'��KTv�9��;��{DֳF�����vk���{&l�g�f:@a���}��������ofa�Ğ�x�Gy-��{9�������
Q��9s٢�Y��=��J]Rc��Hu{�d��;��Щ�@t1YΚ(�|0^���6�8͢�S���O���&�>���"ϓ�L��-���7��<���7��� 1�3L����k3J gc�{ �� �t�U
�Ue�*-��Tk[kZ�m6�V�V6#Xն�*(�U�eb�����XQ*����F�T�kR��TRZ���l-)
�Z%j�Ҫ�ʖ�ҵ�[h�Z�j����#Ye�b����j�ʖ�YZ��j�TmKj(�F����-h�T����+k�(ʥU�QbV�R��Z2�"��X�cZ�R�j��Z6��c+b�*��-��U*����lKJ��QjT�l
 �*Rҵ��F��(6�eR�-)m��ږ����Fڭ�"���d��KK��P�kl��(�YcR�[e���V�TJȍV-b����T[FҨ��E(��m+KIU	Z2+i%ZP��J�R�U!U����[���@�+"��6(J�b��+%�(T��`�eeh�eb�EVQKh�b�mQkR#*�#kJ��(��Z[Kl���5�hQ�Ԫק'.���e�h� u��uwn4����Y�"�;yv��z�a�;��[�y�=�gZmͮ^8�q�Gn�TOf��Ӯ�y���ըI]�ƺn4����j�e��^��X����Z;�݌�����
�kn���9��<F�+��Pջ]��v�s\��[�����-���ݛ�1�k-��l`���n,n����Ӟ{6�ќ�8����X"��4�mt[���\fw\��� L��(�fi�1+���q�UЎ��W��oO��ď�gb�vm�wly7���9���YK������n1��˝�oSۇk��t�.��M�c���[��`v��.�{�`�[ol�y֞8�d�t�:f᧫z���3�O��6���Yt��]��6�e5yz�b���lnn�ny7�A���v+=��v��!�=k�>ܜC��p�q��{c�qv�eN�����nluv����������]�4�������j�G<�q������\[p�� eR���p-ѣ��$����8Z����,�֬\�t�S^���g������J�7ef�kvТN��s��޺��-��p�Vp�x��v펋��tG[Ɯ[�^��Z��!}.l�e���g�;�aا��-<�=�]��I�\j^v4�緞Vq�l.�/vs�Gc����Q�gr�2�Ϫ��{U�n��㒼�fb:۴]Z���pI�v�!�Îc1M���^�k�smᎡ�p�¥�^Z�ـh/.���S;Z�0W<�Z�ьKs�N짥�{b�zN�X��q��۞��p��h#��#��9}�'mc2�{2ٌO<�xP3�#�s�����]�qj�㗑���#O	׮L��Ox9݈ꊗv�N�^wOr���R��ۧ�g��g�c�ދmpS���u�Ç�����2'r�=�����܍��c�v��*�愸���N^+hˇڎL ���V�'�]]�˧xN��=���ƞ�e62�SV�e�j��s_I$ 殝�Z:�%coY�8�����c�ۓ#�m5��T�K���)M����c\8��&y۞t��hpl��jʯN�"�{Lks�+�,�l�Cd�g"�׷ s�*���]ɭE��N2�w���:�<�ݱ��t�/`͛��s,�ۨ;uۚ���]5���{:���'�ܷ<����zݮힷV�8qAW��B�[ Ң���}�.��reON��u�V���n���S���x�j�����ܼbxN7��
c�߿C��Z��2"��ۿ_��l/j�H��ʫIi*��ۻU�E�9�}�I���S��A=��I�I�V��>�Du9���By{�z� �掀����dhDQ��7�_�O<��3.&�Q՛|R���ڻ ����6z���p�I�[��FÛ�H6�,Ir�%��z��{�9������ W�ۻ��Nq{[E;5M����#���u�
o��S��P�"k�[�� 3^u���W��v�J��"րc� �5"Ě3���J���^��	tu�m�mt��m�k�ѫm;�h�8��gF��X��M�{��&��2�'ǔ/<�D���ե`zs������]��ws���z��o��j�����b��s�����[���8U�Q2�s��ޮ���������2�G�t�J	���6�i,�L$n�Z-R9���ߢ���q�D'Lz�R��b�#Ċ>�%�ʋ�lq� ����� oN~.� �����	:��y���,$j��ۺ�� ����X	�j�={Nu����w���8���sjH�%8I.]���W�vƣ�W�iL�H 3�<]� ���UE���;��� 5�`��mCەLʇ7h;��݈�`����*��4�zq�>ګ���������z^����c^hs
j�335D����.n.��\Z������X��X۫��u����������t�W5~��@|�:݈"�� �'a�De��w��h�G�=��HQDrd��ׄH$4߷q�~Ͳ{&j'7�� ��� p���y��h�Ym��Y�\M�NC"(�w= �� �XӢ3��	z]9z���`�e��e�.a�ٗ;5�A�з?��(۱�����[�"r�Y��GX8���uW��3֦�f��Xp�����節���D���y��*����3am���q���7Zd�����wk8��ɎA�̛�� ��[���v��_'N�1�U�dP	L��QX��chh����_H ����+���S��ӳt�~�^N�㷶�3/U��,�>U��g�LD�p��n1�[�-1�5�����˺��GN]s�Ò��{w�0pܨ�3*���v��C5�I�;.�%�ʡ��e��;+�d sy��վ�*eC�%J�qe_mش�@����2<��^W�ߒ_|���r�j� �OD����~��(k>���T�5A�!6KKm�D�H�����F	��}<�1���D�OOD�D��}�����"�%%�DT�����~ �^:L�n݀�$ќ�Ñ�9}���m����i��G���[�rɍ���5|p����Ү�6�, �;�44.5[.�s�yw��xq�B-~%�_��Ww;��B��e�Ʈ��� A��=h�v��΍^}��̟��SL��@$g�o@D��	�O��(7��	�*�5
��g�m�GG1�G;�27h)��c���|�D���m� P�$��d}H��5|� >yᨐ�޺�k�nM��gh��|fv�E��޵7*%Lʇ7h=�,�1���aW"��	$��컴�;+��-��9k��/���X%z������0L�=��I�oY�,;�/������z�#> ��PI|�ޮ4l��1�Z0Bڐ�6���P��p�F�u*��ۼ�VDDwf�%D��??fBz��{/y>Y�Pfw]�\e��N��a+��j�H7�ЏG��g��h'��� ���� ?]�v���x��Hz^���B�o�n�2����wR�}�!�_;���Q%V��J_C�\��#�ywbPnN����#BrxyyO����T�а��5��ܽ���V�m۞C;��k���<��dR�{������p��]���lN���2�n�&�v�y�E\T��(�ݕ��#�7�J�طbth�;���/��g�{Zg�_Y�읞��n{n�޺����ݼ ��κ$��t�뷳��\v:���c-��q��X�	��.��e5�3�y(kk$���&n���օ�ܾg��ۅTAٕ��{X닟@�ں{��1��I3$���wm�� ��'�� �:v��]������߽U�O����t�+JL���1������{/�f|���^2z�� vW����;j�) �F�ر��vo��s����f�.�K�e�V�I�rC_ �"���o_F7p\��$ ���+m���{]�hg���h�.8�thOk�S��{d��.zv�b@ >�mPD�GOM���鵜n�륖7�B}�7i|w+Tp�0���ͪ��i"R]�5|�XdC�	k44I������j"���wcȆ�9���G��E�S����c����%0u��픽�uώ�z�T��N�"�E;�;�tfWKsK���w;h�3|����nFG�ׁ1�L�m��=�@UwM� �X�������w���ՙ�XQ��Q<��9�6�H�o�<2��h��m�m��Hȶ�K�����)�	3lo�^�����%�!��������mOߑ`D�j�) �m�E�^w{��>7�3OHM��n)��!&;��U$I9�ʣa$���v��hep��}�-"V�j���H-�˻Nl�Y�	p��\�O�y�1�)^��8�s����D�'��uQ 9�ۨ^����vL��'�Ѱ��"�o3�)�ӆ�I�\y��B.}���p��y��&�}���x/�Ŵ�l�G���r���I��7�=k��c�+���F��
h����]�,����C$���R�8�ʘ� �%۹V-J�;�b�.���F]����~]TI4�nv��r�aQ�L%8�D��a'�ڽ��+�0�i���� =��fDg��vzի @�>��	�rӣ^��u$�߾i�`�H�WIQ������kWĒp�c/�~9���s���\B��~]�X�)�����OQ��<���u�4k#��zf�Kcק%�DynRq����?/��$�s��"?����� #ַ߳I�ғ-��$�os���O~-X���$�O��'L�$�~�qR ߷@'(�ڼx�IV[oԐ�ًI�/�%�=�Z�$�&;� cBx���Qߨf������� yvҤA$�_�r?1���G�=|]l�&^�s��k]C�r��]oDk;��;E���9"���|[mu�ww�	�i�!$Q��no�<�H%�yW >u8�0�ħU�Ӗ����w�<�(.��-#�Gc����'�^ �,"��go�n�@/z��� y����q�%��a��.��K�o���!)�X6����h �4ΗH��f�t�U^ Ǻ��� u8� �x��*\̄�]�Y��q`u��V|�ʵ >D�����@4|���W�򼑚X�(���*��2ʕ=�7M�Wϓ�>xzx�D|-�а��G��"���i�����ۇ^k�<�w����I!&m��{��*�SӘ7$�%�s0�f���/P $�vݝ��З���i/����I|�^�rt��CC���c����k�8K͇�;]��x�<Z��VN�p��1��� �ekmڑam�&ﳉd7)��.{���6���z]  
������+�^;Ewm�����N) ��>s��&b �=��n��Kg{�N%o���v�JI~�f�I$�n��ylW�����:���Cgq�т�Q���� ��}�ńDEk�Z{����@|fˊ�~�{3���ȗ��x�E�v���VQ˚�4 ne�@$^���� �H�w�S���s�H[�S����8�1.fBF��'sٙ�Wz�(�ժ�Ҋ�LwT��I/{�}�"I��v�Z8ބ����rV��rμ��r��:m�>�d��5E�S���d�R�ӥ6��̂�{3i)U{v����wc�U�>�~`y�`�FT��WK�Q:�=�v�q�����Cnc{�; � [��Y���N�f�g�KW^�FQmn{[	u��l�v��̝&�՘0`�@�;�vy7O��Z�lM��;r��M�4nݹ��k�]��'���zMrz�ۧlvܑ���=pwg���[������y'ǃ�j2uǒP��r�XZ�<p�^�����9^�cI�٩�Y+�Kt^�(̖��:�cv��kv�V�z=x7;�j���;/�����,W�P�gs��"��^` z�Ԫ#�n�>�Ӻ�i/v�W� ��{٘'^�$2�" �l�v��]X�J�k�o��mL��|@ ;w������w�Z� ��Y��Qg�w������O5"��49Q
��=]��A���U���7=+#�6�Ƥ #پ�bX�	 ���ݤzf� h!MA�KV]��`�'%�I�w�� 'ܳ���:�-zJ�ݣ����:�ٙ���,@S���USM�{����n!7_��;�$���m� ��o� ���R�-�#��g�@6ɉ�L�v�*a㑵��[p�r긓��p[\��];�����LCrD�b�L���I"w�m��$���m��s9�U��tTg6i�l��'߶{4i/�ғ-�XM�1���z] >s�߰�r�ޓ���b�/^f7ڰγ8o�NT����Z�0c�cu��6��mԦ�f{�������8�O�-�G[�\~�����W�W��W��u��" _���v�,y��W� ,^�_r]������Rc�ف�O!�9���MEx �=.�D:f���-��ʻ�$J��M�-��2�3���+%eO&����Ӓ����eN1=���o����k�����Y+*�����o�83�0f3++�]��2�VT�30�s߽�}d�k\���n�����J��YS>���+<d��/���Z�4�4ܺ4y�J��0���i<d�fY1��LN}��wǱ'Y���3_[��	�q5c1<�7��Y�q�3��f	�w�6i�c1��2���{��âu��?~��}ӷ�^���;�����i��v*=��[��Ѫ���,Vv�Q��Z��\r���~��Zk���m~8�I�q���7�Ã��&e�ɆY�?g}��y,�LpLd�19����2q;d��ߋ��nw��,�f�)���w
��c+�1��뿼٦T�0�ba���r��j�kZ�W<��'bo���������C�o�~�������o|�ј�!��c�0���eI�q��f2d�s߽�}d�l�K��dǜ�l���Ǖ�N�u�G����C��۹��5�k^m���q��o���+%ed���&'�����蓬���La��B�}���U��
�^��_��z�5^hl�O�;9��]��ޢ&r�71g�.=�P��hZxNHk�n��-�2���a߱L�܃K��<��R���bbbu��F<���^$�X����+igo&��-꼈^�2�;W�1��Z��v�R�d]��/��zE$�VH��>q�ڧz��ID�Kp��מ�t�f�g�a,i�+^{��������mog�挅����DR��s̫wv��#�Vo���bm�e8�fm��U\v�y��jj��Cy�&T�wM��0umo����V�
Ӓ����=Ws�nҫT��1V��d	@���FY��5�g�9y���.wѫ��b��גƧB�82���;{��q&n�4�}2.<'=��ѝ�8��r�rk�e�ۯ��h��f�{�lrS�����b�/n�Y�5��������oU���U��S{:�g
�v;u]�O���2���~�nY�|U��G��}���}$��^B���Z&��Sw�F�|�����T�����D��z+���������׾!���F^�%+�֭�.}�o`7}]�����:�㳖vZmZ�Z��e]�\v�wW/����%��8r�[��çoc�,XA��ṽʷ���x�����zQ"�ȣ[�E�����m�O�+����I?Rۄ�N���ף������٫��r(�a%ӧ(���N�t��cDw]��@r.U� hgr��J�Bi��ֽ���j���������km
5*(��ZZ�+ebʕ��B��#(����mh���6��EB�X�
�JԕFE��B�X6��QIF*��b�P�� �"�E*��,�*Ĩ%QF�գ�k(ʢV��+
�mEB��h�VKX�%T����%���ҬQj��J�T�J��@�j,�e�V��F
(�+R�T�*�-��b�XҶ1B�-����(ȵ��V���m�ګ(ƴ,����`�FTU+Uj�H�YPѰJ�TQPT�*
J%�� *���#[*[T�����-`�YE*����m`�d�`��(Z�ŅJ�F��bԶ��
��m+eD@��m-me�Q��*Q%F�"����P*m�����
2���U��R�T�b2�6��)�EF�*)XV���ڵ˘���?Є�?���}���0�c0C�����y�L�x�f!���Cbs������Y�2y��?4ә��3Nc|6�$�q�������w�{^k|��g++'�f0�}��ג�d�1���߾�����VJ��2c3)��y��Y��7����I�W��pC�y�6i�<�1������[.an��C���������!�c%eC�����gc8��{���s�y1�a�Lf0ɾ��<1�'�3++%N~����'Y/l�LpLO~��w
�'13�>����}y��χ9k�j��m�I�9�n9�F5�kZ0VNx;n�f��8�^#X���}u�cK�MˣG�d���~�w���&3,���&'>����蓬�Jʘ0�bd=��=��N0�c;�k�y�{�]o]3�����P���1��d��}���é�c������j��q����19�o݇g0�1��}���~���g�7�{���Ɏ&2c����s�}�βu:�&&G1�e=��{�Vp9d�W��}�������:��{�S�1��_w�[�M\�ir�pY�pa����w�N2�VT:3���߻83�J��YX5��Û�\>��y�?��YRz�1���~��񓽳.Y�������=�+Ȝd��~�˗5�f�kZ�כd�+���ى�>��ӿ�>����߿�>ed��Y17����2q�����2~��{�+8�a��b�~��Pg�@.��2?nx�$��m��j�?�\Ge>�q�43d�~�U��e�g]���|^X_1lCJ�5JZb�.D��gr��}�1�O�>����?���Fc1f&������Y�3����s4��i�o��Ĝ�3����p��f2fY�?w^�fxY���r����?��q��������N��LLd�T��o�³�,���I���w��1�<a��מw<���>��s3Ff±���-uڙ@�Xg�Ľ�����Dh7Ok`4�=���#\��-�S�u�>a�}���u��C�c1�������c8�YXbc1�����Y+*O{���ロ��z����g��;����2~��YY+������¼N2b?o����iti�thߌ�8�{��f'����2Ɍ��=-����I�����蓬���Lc12~��{�+8�a��b�f'{��ٌ�x�f!�1���}���~��s�������߻���c�~;�k���j���1'#���߻�g�����Y�?w_ofyf2c��Ɍ��=��9|�����k�������LL1�?y���+8rɌ�$�c��y�Y+*y3^��\�SW3Z\��8�a����w�{׉}��7�{��YY��b�f'9����1�C#1���2w���eI�ęf2`e9��{��o�o��}�����.��Lr	��߼��^	�LL�{��.\�4kY�y�N2���}����1��LfL�b{��{�=u��7��{��w[��&٤�f&y���q�3��f'���6c+%eC���C#19��{���u����7����+�ǀGD0���a��\��
�t��'v��0	�m~������@S�t��ɧ71۵��+!�>E�ޟy�H_�I	&���B��g2�a�c�M.�Dv`���]�h�[�z��*��E��m��h��V1pf,C�Y������|1��t�T2-sѣt�T���vێ���������zǁ����.磶�j��s�%��5훳r���s���'[j�Y��������{eD���s�g�G��l+��h�6[1�[]g\��9�e��E��c��V�Xs���s��F�Pwku�v�E��s�,���Ѽ˰]kr�<�?�����:������l�'��3��o�G�J�ɓ,���w�<�1�1��LL��}�d�tq�����ܿ�o��M3�S߽�gY1����!�����eOc1���k�9����<ed������=�f2VT����.~�z����6����ρ��!�1��"c1�{���Rx�1&8�ḑ=��w�N��++%u��֏P��xB:�z����<~���c��X�th�88Þ�ى�q��d�VJ�����D�f9c11�3�ۼ����������y��Y���3++1>���f2�VT<f3������Xv'Y�2w_֚᡹���f$�q����au���vw?^�d�Y������7�<,�Led�	������w�N'\d�VJʞ����+;���o��>�'��D��pC�����eOc1.�޹ni5s5�˭�g���&�w���f3�3���O|�~��1�C�O�߼s~����x��3����eI�Ę8�ḑ=��w�N��.Y���b{��{�W��d�y�y���y��\♦�֭�O]�.��S�[͢�@v��*���+�Nu5>�;�.\�nhֳX:�l�O�{��ݘ�d��,���&'�����'^�1��0�bg�}�B����f�����OO���C�Vy�{�6c1c1f3������﬜ea�����M[�K�a��q�����ߛ�g���f2P��~7��h��l	`�s���Z
����}ݶr�+?s��m�x�QI�=�4C�;�r��{y�K���k>>��M놷�����]�HI&M�����3��L��c&8&2ba��߿��'S��Led������<g�Led�������ߩ�Ǉu�<߾sf3������F��0�U�C����'�}���:�Y�������}���g��f0�1���~;sZ��{�5Θʓ��J�ɆS߾������1��1�=���3�J�����Zu��9�F�8�YXy��Oz?}���~�7���H)���s*ψ�? �C� D!�v�G�g���9Ϸ�(j���/�����{��ϐ��f!������}a�:�a�����n.��j�xq���3�s�3���c&e���u��g�c&?wz��}�gs���d��Ld�������&2�VT����<g9d�Wc1�;����eO�3�"h�����&D��cr"B]h[c�vy�Œ6N���yQ����;,�&m���~���j�kK�^�g��a���Ϸ�tC��b�C���{�x��1��YXa���<1�����~�~�'�u�d��y���'��.c&8&'���C�����̢�e4�hcٟ}pQ�>��6bx8Ɍ�,����ߒ��$�y矾�ĝf9c120�b`{���8�'c1��c2	���6c+%ed��}���\ۜ�}�{������Ϸ��Y�2y�~i�3K�4��l�N3��sAǌ�&Y����{�w�<�1��Lq1��j�}��w��ny�|0~�볈�`̡ӇCD�B�c��1�o�n����of�Lk�τ��*�]��ޘ�{�[&���-TPUz3�g>!$�]���q��VJ���Lfe>��{�Vx�Y^	1�����ٌ��f&K��z�*a�7K<�S�1=���Y�'���5���x�+*f3��oݜf3����&3a�w��ʓ��0q�ɆS�}������|���_l�LeM��p��&&K��>�kZ˗4�.��q��a�w����tɌ�,���&'>���񓌮~����M3���3|�n�'�d��=���f!�1��YY*s߿}�0�u��?g�}}oU<d
*����(�!q
d%������u�f���:w����z�����~�ԯF���|u����bs�o��Y�'�02�a����1��_"c&8&2ba�~��A��T>��O�}�u�۹�}�u����9d�W&3~���f2VT��{Ӹ��j�kJ漂�'����}d�+;�b9�u��w���l�f��w
����a�Lf0����4�d��<�32e9�߾�Y;�1��ɏ��x���u�����_t��d>�f�]j�Z�`�Ͳq80�[׻4�d����d��߿}�=I�c%eLc17�����ϟ�<�
�2VV~C���i�����C��0f'=��w���c�o���jܺ]9��gr8�O}�l<���;�u�s�βl�1�,��u��yf�1���	���?}��|�'S�����&32������;�ٗ��כ��w*Н�	�F'�t;�P1�6�ǐ�q�k[���g����~Nt��v��+ϪP��:��Z�Y;V�3�B��4��$�c�o_��٦bx�����ZT�0u�<�Y*o��o��!�c1f!���O�{�vpf3�n�>?g;��>�7��L�8��a�o]٦bO#�Ę8�ḑ�������l�K�c&8�������2T����͟����z��V֛b�{s�k��Z1<ct����@�ҩ�,�����jL��[���1�9��͚O2c+%fd�������I�c�Lf&1���>��!Y�J����������c�>|���=f��s}٦b�b�f!�1;������f0��ߍj�Ź��l񘓃���߻��&e����?}W?]�󽕆g���3+�c&8&2bg}���u���11�Lfe=��{�VrrɌ�D��w���_��o�~5��}��of����<���;��#��`�� ��������Y���c1f3�}�vpf3�`�f0��c�w�߷�o>���k�Lğ8�I�33)����'Y/l�Lq1=��{�W�8ɉ���z����f���כd�pq��o_l�gvk�"���+&���&2�T���wǩ:�pI����3'�}�B����3++0N��f��}�7���fs�6{����4���b3{�߫�~g����҄I�N�L�%eO}�6��L�1�2�a��ٯ�2c�3_a����2W�1�&���|�'YY*v8Ɍ�)�>��³��c+%er!�wl�1<a��������?k��w'�*��"�Py����%]�[��!�ƴ�����D���b�0�ވ<�,�yv,�9�5�z��0�k}+�T ������W�Aֵu.��:3�H1�ss�ܦ73�;s�r���T�U���:�ᡀ��n��le�En���{Y9�-׬#e�u���u��\�v�h�[k]�u�ˮ���`ͤ�*�L��;m�9���	���β�B;���.ܼ���H�YGٷ=����l���y�9�a�F7=l!�7nºm�uƋFp�l���么�7-q�V�'�1��]m�Jni�ΕmgrfNg��Ҵ��9���3����F��W?��*1>�����u��C�`3�����³�J�Âc1�N���LĞ3}�g�^��x�:O�}���'{f2\,�Lq1?s�=�+��&&]}��Y�k�]kK�++3�y�L�J������������'S]��o��:�pI��Jʙ=��{�+8�c1��3���w��3�f3�c1�����'{�w�F�g�����0����ɟ�������f$��19�7�Ñ�q���a�c��}�L�J�1�1�>�}׼���n����ߙ=ed���&32�����2VW�1���w��3��L�{Ӧ\�9��5�q8�_}���5�������g?w�zͲVVJʟ}�~l�f3�df3bc1���{�LĞ8�d���9��{�2=޳��������;1���d�~sϷ
�'13�o�u�]j�ZsUכd�r8��o^��x��d�d�&'�����'\�~���o��181��<��>��N0�c%efA=�w�f��y��0f3����߽�Xu:�a���������}]9�p�9Ț��D�3ٵ��s^�e.�\�K˲���l��Bɮ����5n]�i�/��ԟG���͇�L�1����g}٦i��	����ɉ������N�c�����w�����_�2z��<���+9�&2�VW;�wݚf���L�����Z���g��*q�'�w��tC��`!�ƫ�HhY����� ����{�
�[{_Kj���&�fɺZ0?m����]7�u����wՐa����m&�۷�%l#l�t�����UW�~���*/l��f3�`�f2VV{�w��L�O#�Ę�1��?�{�2t��r�dǾq��Y����]��p���d�˯�z�3Z3u����*r0��l�4�YY+<�&'>��wǩ:�d���f'��{�]g�����;��OF�fc1�'��l�4�YP��C��~����S��^��N\tj�����bN8�O9����7n�}�����߫8��c&f0�3�ٯ,�&8�Ɏ	��������'��&&G1����y��Y�����>��w��G�d�+%et!��vi�Oc10�wӣ��nf�LאY�J���s|d�+?!��1��O~���+<A����ߍ�������c1�����i�d��<q�Ɂ����{��t;f2\�0�C#�z���g���������Oy��wW�8�nW�q��[��͋��v�h4��!��=�e�urܮg��}5�]j浧Y�u��?'��u��f��l���&2�T�߾�|z$�1���0�ba����!Y��a��}�:������8~�f3"sZ���3L����1������:'Y�<���8jܺ�\ӣ.ͳĜq��������&Y���w��u������w���?of��J�1�Ld���}�d�tq�#��̙O~�����c+�&3�qr� �ܥ^�<���Џ�g�A�o�k�f��&��+%O��~��Y��1��3���oݜf3�df3`����v��;ݝ��1[Q��"���6��]M�X���d�6�V��{�R/*bJeY]�����]v�!ܲ�Dx��mIJ1���/������	}������i�I�q����>���8��zY���b{��=�+�8ɉ��߽usZ.V�Y��2T��k=��'7�~�o�Z~{�M�	�Lfe�}����1ȓ������s�|�g�1��C��;�w�f��[��~����cسhq��Cbk�;��ñ:�a��>4��F��:�<f�+*o�7�ã��&e�ɆY�?fw��l�����]��^9��2q�c&&C�s��u����LLd�T��7��Y�Y1��&3�i��0�byï��u����׼��������{/�}��.��K��I�l+ؙCkX��:L��w����nf�L��Y��a������'Y�C�df3߹�w
�++D�c�4�I��1#�}�}��h�v���e;��{��t��rY�����{�=�+�8ɉ���t�9u��֝f�כd�pq��o_l�1���,��;�Î���_|�O����D�f8����0��<��Vq8���f3�i����b��35�/o�����ۿ���/߻kO�H��?/�ޖ%�sU3N��gq�b{���Î3�����w;�vk�4Ɍ����LNs��~���Wo;�9��2|��11�Lfe>��{�Vs�Leq&3;���f'�1���?|�l�f��d�<eNF�����y�����\�5�^���%eC���O��|�+<C�1��YX}���4�I�Ę�1�2���}�Yg�8��������'=L.[Na��"��ZH~n�^�3��W���[��5���A+��ve�v�e�z^��ֿ�}_}$��>d�ŘɌ����
�*p�}�˙��u�ˋ�*q�׺��'��Led���9���wǩ:�Y�����y�,�%eN�����NF�d��=��ݚf!��f!��b�N{���F��~���~�N�U�h'rۗi��sn��f�Z�ew+���n�]�5���`92�Z{�}��[���`�|q�I���߻��&f2VV���f�,�&2�W1�����'Y*{L���gx��{���y�³��LepI��"����L��3��::֥���s^Ag*g����?!�c%eC�}�^����������tf3�df3bc1�~�w��LĞ8�I���L�s߽�}d���YY*���߿ky���~{��5�o�¿�������Mc�Z�ִ�h�y�N'a�[��4��1��Led��{���'Y���1�3>9�����>�o��=�g̕��C�������3���0��J���}�8�þ~���][�5SZ4e��8�YS߽ߛ�N�u��~sl�%ed�Y�9�s{5�f2c+%q1��~�����Led�̧�s�w
���~�_����N��I��7�w͚eOc10��ߜ��ӗ+O!�T���>���Ρ�c%eC����7���q���~��Ɍ�Lf0��}�<4ʓ��bL�302�w�}�Y;�1��f2c*{�7��^H�dĳg5��>�w̧�!�s�����h͗,�x�Y��*=0k����T��|��8��G4':�
��R�Ռ���O.�=��*��W�6�?z���A32�v�4q_޵t�
��5��Ǔ粂YA]���<VM��.;�.�,z�@ܷ��멯��;ר�����3���+qmI�;e�6��Q*�#ք�疼���v������eد�^�6v�#�r���Z��|Ê<������z�ws�6���aH�->(��9��Nk�5�U�{�
�.�k�wW6�w�����(ޅ{'�z
N��+7 �v�}��}�Ѩ��9����t�l�w�K������ �zg?e�1��ў�ݯ�o��[���#3�����>Ǩ����t����ۺ�e�Ѵ7sl'zDL$����e��'}[X��Ӗ�p[rV㢥��}Y��[�f���q��Y$t��y���I���:]�l���`5�)P�V���Pm�z���b7��W\}	ӌ��!���P�����=�{\�lK.'Vo؝�l��o;ʗo�*���
	4x��;�W
��Ҭò�9��=��qW��"ߊ�3x;�$��v71�Vir���K�m!�l;�86WF���Ej=��Ä0k�l�`�U�8hm�m~\�D��������l{�P{)�:�DSF��R�ʷ���>s����k]��\�߼J�n{Q3[�+U���R=f0E��Z%�4�sw&�Í�Y�t ���;�{��N�8�SrF��T,�IB���o��X���(��Ub��*,Ul��m��5j�k@��bҍAchV,+Z�6��*�[J)��c��
�"+Z�S�J�iU���mF�R������UQI�Z�ie�mR�9�Q����Z��[J9h��� �ڱQRV�J�ʢ,*T�J��q�-S2�Ġ(�J�jX��Zш��Р�*"%�Q����r��b�*��J�Eb"�d�3S*��E`f�-)m,�FTZ��B�UDpeZ�m���QF$Ƹ�墑Im
�*�Z�[J���d+FJ�&e��j�R��C�"֢�j���5�V0*(TU+*KeX�Z�T1�IXb�k-ind�+%q.P��PPP[hۈ�IDZԩmZ������Q1�(����
����ҥe�Z���J��Z��*��DbȈ��+(�%Ƣ-����&e�"��������m��BH�6z�Wq��;w��:��H�t�m���<��E�h5<�s��kW<�Pn�A�rk�5�x��#��nZ�������o]�8)\�b;Qr�=���m<��,v���R���v}�̖�c��f5tt�X�4Fz����Om��V���).�wPP2mp��A��r�]6����$gK�{syem1Y wɋ�έ�v��m� �1�:�n�9��v�S��q9ɁnVRM7mK���G�{�[�h�笩Bn�:m��,�gb�\��n�Y�4��������
�j���v�`Wc�.�A���9�u�Ŋ�K�1�>d�s*���ݬ0�p]X\O��=��؎(�ݛ9[kn^c��>s�yp���m�a�X��7S�c����b\s��^�(�kY�bwe�s�%\��˞Z�-����2�ٷn�:;;vκ��rX�vv��,v��qv�%�w���0�vɔ0[m�]��E��#��j�l�S��0bp�c�M'g���8��n�U�Y������a'`��;�;�y�nm\k�S�q�{g�rs7�p�n�
��3���7'#�*웲h:ǎ�k!����N�A��N�y�-;��\u��;n�d�pW�b<��zvJ�v�y�+�>\��F�ԷN]��qsË�gڵv�n �vR���q/c������۞p���Uuls��|�8d 4�Y�W�Ӻb�]�m�\Z��<vzvm�V�����S��mq/�n���v����6㰅�v������=�8ڡ�>��y��ŋ��_�k�|ǫ�^6=�	u�p�D��.�b.��6�7�]�
��|�)��Z�P9zu�+qz����K-�7el���v6�c]Wmu�]=��N�0=o�0���>d;eVvqn{b�-��9���U���8���<��3��$w8r�n5�v�v�s�v���xr���..y��aٺv#H�������_<�5�ذ5�c��1�uu]SW1�kM�ֿ�BI3{ݝ����:1h�[Y��j��u��d6��X�q�	��#�������͎�]�q�1�z�e��lUu��OOn�z�pX���]���y��^�&T�+�I�Bx���<��f6�F�4Z�`�n.��*�ѡ��u�m֎���9��W�/O�2��%�Ě�m�<F۶;n3�^�׵���b6&=�[ti�6�#��K%�������Y�]�UFỐհC9�����h�Ŕp!u�.��������]5Ѭ�7+�:�S��Ú����x�&3&Y1���>���ԝf9c10a���߹�B����ax(w��~9c- �z��|EO߮�2��1��Fc1f'{��﬜ea��s�Eˣ+�:�f�q�by�o݇g0�1���h�;�g>ٙ��V����rY����Ɏ&2baϿ{�d�v8ɉ�2c*{�7��Y�%ex$�c��<�{��}�y|�vi�>�1��]�tu�Ks5���n<N0��?}����1��3+*{�7��1�C���5�?~���7�j��~��L�?8�I�33)�������VK��d�������9@�s�=��km&�$�{�N'a�_y��Gz��ֻ��;����Lfd������2q��Lf&1������+<N0�c1f3"w_~�f�P��\���������i3�c15���}a�N�aϼ��WV�f�֍|6�$�f'���7
�9�c&L�w=����Y�����}z{�y�}�̕��������'YY*u�LeO|�~����c+�1���u��6i�<c1?k~{�����wީ_�9R1D�h����D�"��"f�֚��i7]3�j6瞌b������\D����u�>a���~�}d�+:�3���O�{�w
��1���0��熙Rx�1'�o^k���<|s_}}�:�L�'�Mw��}d�l�J��\LO���w
�*sY��2鮍f��_8�S��מ�f��1��Lg�v��������~Y�K��~�"��"1q�	Sޛ��7^����%�L���ٙ��E���o�G{]�5�x�f5|�+���_��£����f9c11�3߹�w
�++8�3�w]���3��C#1�����L�2��u7����d�+g��z]�E�`�xq�I���9�v�3��������߶k��l��c&8&2b{�.���~מ��8��S��Lfe=��{�Vx�Y^	1��C��~٦i<�L3_t��Z��kZ���8�bk�{����������z��~d����>߻�g�1�Cc1�&3d�Z�f�+*Of2a���{��ɭgo��浞�u���d�_s�ۅx'10����X�ֳ5�74f��'���7��'��&3,���S߾����N��oǙ�{�3������f'�~�w
���3��f'��}٦ic1f3�����}�Y8�ù��w5���w���uf�ɟ<��`kwgY]{W6�l�L%[m��Z텔��3F�����չ���Ѣߍ�ğ3߽�6q�d����c�wݚ�Y�LpLd�VJ��~��:��VJ����������>�y�wp��,���Y\l��!�g��̆5��E/�j�,y2�T��;����V{1�7�ם�{��.~כ<��JʁR�S�����`Q�
Zs��`s��i
��U��/t�9�o�>? �M�����N�f��_ S�'��٤�����T�~�ݜI�(��<����_x���]y~X�]��ZM��F�B6��CX�nϮ���Ƚ�������x!j�������9$ֺ�2v+��������G��aRT*J'�s�ݚH,�2�PeN}��������0u6x����~��צ�������� kk��yHV�
�O{����J�X{����V|k������;'�?	*�ݚa�aX[����Z��kZ���#
��>�ÂH)��y��<���~~9��}�و�P>���`xԂ�����}�`x�y
B�~��
�S�������=}י~����߹���1�[:.��X��UԮ)z^�Y\ykn�ݸ.�,�Av��I\�f`r��Il/о�<�f��@��� �����8����n��*Ou��y���v~$�>�;��2x2�Q����{��9YU��r�%b��X(�;�ˠ,G�$>�}�����U��'�B
A~`T����|�ȁR�V����<d�Q%C�y�y���7��������i �������3.��\<�
}�����8�R���{<Y,e@�P<���~p�<�o���9�M0=kƤ-�}����)
�=���n�`T���e�]�e�� �n��͚O�쿑y�?p�+(�S>��l����+��?y�F ��y���������B��W��N�c�V�n0Rw��+K��*�]��w�ҖA��{���!9]��
����4��K;(��Xѣxwu��Ow��� N��7�{�`x�������&f�����Aa�7�� �;%�~����^R��g5�n�]���
�߹��� �
��|������D�����L<V��y��7�=��4y��5z㫭�/n�]�Az0������㫡���7Yk�����OM]je�ֵWY�*g�~�À�Q
�FV�����*A@�*�s�4���s��gu��HvZ~��=�9H6R�w~�p]π8;w���m2[�ˀ���� ��%f�Ϻ��:{�u{'���s�:��X���~��Xx0�(�IA9���d񕒌��t�e)�����'"q�;���t\և2�-��Aa�~������,-��{�^B����"�? �S�u��f��{@F|@�+*{��y�)�
s9��4���;�?{�����3!�aQ߽�����ה��?�'���U������YP*T��xi��jAHRӟ}�����=�5�q�_�}���9��n������e�u]j踾 ��'���l�x�YY*ANw��l�N!��ܽ&�x+���y��*A@����Ad񕒲�=���' #��O�OҖ���?U���y��Wd�):�[4��]��zB;�Ds��� r�T����Wز���=��+|��U��3���iǦ���|)m�\���֭[���[��������M;� n��[n"���<=s���1 �`ۍ&�$+Ϣ��z1�:�v_0l{/ m�����й�j2��n�vNk���v�̦λzc�8ۥ�i�Q��[[��-�oR�]�sI�nS���N7m�l��d�ɖ96�nql��q۲ss��^��v�z�m[ v-cm��y��@Z7�]�űpy�H=�؎�3�;��9���F�k��WW4��0��~��Mf��`����a���{�)i���i �
�R��}�ND
�gN�C�6��m���w�,�2T(��P�s�vi��
�ϻ�ӭL��k*�7��*g�y��1u�<�s��{��k�X*×�w6*�������_&���~n�7y��̳$	9����tA���u�?}Y�|�C�3����)��l��q���`JQ�ʍ��gM�x��٫�I?���`��2��1C!�e&Af���[�%�jH�1W����I6d�D['X�Ɲ���Q'=ٷ���F�s?{�뮪\�U۱��C�vjV�(���5��x�����!k���������-u��)�E�d�w���A���@�\E��n]��%�u\��R罆"$���3���|�8,e���$�y���n�ۋn�.f��8�-���U��^�q��0�K�F5E�6��T<��^ѻ�h���~�|>�E��	���A�I���|;�ɽљ��s��Y�	>e��Ee�ݒ~;��|� �ȕ�wei��:��������ޏ fWx�f'RE*�;��=���V־  �˒ � �(
Ew�d�������ߟ·�$�c�vh@\��J ��D�7��e�<�=�����ڥ@{� � �]��	߯͝�4C�]$A��X������wYs�iz�:���D�Zc<Ab]�:��F����ۃ��A�k����A �y_"I6�yљ=�MY����Iީ�W˟�ԉ�ԁ�E
Y\蟌��xV�t�7n]W���w�������sb������j���w��N�P#$i��]��{AI�}��L�n�e0�+�n�< �3�T�tc�g_s��߸m(,�}\���!�ӣ���4{�����{е:�w��l�n�Ɠ4�k�ꞟW��������@�޺�E���ٱc���WN�75�G0�}��n�"�=�#��M�w_"I#��I7��2���$����ɦ�3+�f3��$Ux�y� �w{���"�dZ���0�ʔEy_��$�{۷��JT(��˝�"q#B����%�,�0�˭ո�p&p��r�J���vz둯_���ߩѳ]�(
�{��@$7���&��j�=�����S˘��$�t>u�A�N|�7gz�Y]�GnP��������	��}��$�7��w�ݥ7�������W=�SR"�r�)ek�~$߻��_�`�O��t�t��\O��W��I��۳�[�2F�hDE��p��),/������ ���K����qZ�wA3u�{�_�Ě�yE���k���~;��۬�v--��מ|G�U�ݗ��[�P��vi�J�Ha�	�޾�_�磌���g��7�}�5�SM��G0�����?�~�{}3��}��I����${;v��6>�1������_d���ɰS#f�8��[�RnG�;b1l�D�L�ݲ�i�e���>�:7!��T�:$��ݷdA#c�U�#�9m����_: �@9ۻb�#�B"\��#%J �U2N�r���^'ec.��?H��۰I#c�TG{&���v��y�l	�9�d��v�:�r-�D� ����^mM�~${ٻv	 l}��\����F&�!�ϧt��kP����g�I��E��v���R��H>������]�dQY����E{L��]W��.p��?~��$�1QZ��OIUW�흷g�����8��wxȌ8>im�oQ�T�X7Ŝ��m��wu��S�Y^��U��9�W�s#9B�u��v���/�?\���Ā��e����6M�`�n��&�67(t�jUoO��{R�#w�,�3t�z��;���p������7���wk�}��='\������5��3�sn��4[�M�رn�8]�ǀw2V�k�Cx:�v��]��-��غa{W
����v��ݯ;�Y͸���ۄp�u��kv����b�0��{<碵���>Y��՛��@	Ө�yE� {<-�4��b�v��C���-Mԧ`�N��Ho�Ͽ����@��.�f�)
�0� 
Ew�BQ��U���2<�E����� h�^+�:e��=r��ͲIȻ H'�W���I����ⓩ:mhd�p���6#%A�]02H6o9��N���W�q<��zƂ}O�Q&��:>u�A��n|�5`�w]��U"Aƶ��H�����o������mWȺ]j�+�-���@�������ݻ�e�.�-���	�H��΀$-^�E�����?g����.B3)ęe�f4������q6�.��
�3I���-�+m2���>y�}��2�j",B�:0�k�	7��vdC}�(�.j%콠*���E�[���a*@ALP+��Y5Bt�ǽ���V��Oq-`w��0rOz�ɢswO�ֆ�Cg8��;�r [�Mo;s�����m�zݮÚ����Vo�^i`������>#���H<o:��o��ذA޼��2iD'�sΉgx$$.	�.Ưw�|I?��d,l��'A�Ɍa y_��$_om�y'��%/7��9\�Ň"�����@?wm��U��}w<)�k�H�^�D�׺�����Bn���U�~8kr��]Q�YM�髷D�}��B��Uv:[�[��oϺ���:���v�����]l��Y���5�n»���ԏe5�x��}��~��V�+]L7<��~$�n�X$uWc���h��SWv=�PyL�(M�v�uo��E���/j�ͳ�g��e��u�?@��۰O���D���ضS�<�~O�*@APQ]޺�A�]�P>�����}�֯zgd���~u��g=2�Btyh<W[t.N��n�������h�^��|J~����j�����}<��[��EZ����0/-����`M�{�[7�#ܗ|�K��ZQ��o.�6�Ѫ�b�\ܻd�Mu>po_�Q�ۃT�ͫ�I�vgi�5ދ�|f���K5t=ޅ�7ýn��B��_�#qWZ=�R,w�?S��|�
4���6dk�c������R���0kv�q����<�=������m���)���K ��hozh���S�giMn��K��n���e��b�:�;�ٸ�ȥ����v's3S��w|�R
z��*���	�GA����j�*�]Z�N�˦_	��/u�]��w�~n��.�YV^º��t��[�921�+N;%�9mk�!��*S�tþ{��z�.�x*�Te��d��#K�f��cf���oj���h��v�ZŚ���r����{Ҵ��r�/_Yk�iԉchOh{x���p�A��v�T܆.�w���Z�Q�P�xY7븃�8-�ͯ�T{:7�q�����{B�;�}��e���8�q�����1��a���S�;�zv̈́��P�,n�����;��ώ� �B���hюJ�����wo��2
x������e�'�����f��vن�r{���sl����ə���B�u��8]A;��p8_���~��To��^�=	����`~Z�qE���[J*�[j11X��UTDĥ��F2�L�.��DEVVJ�Y[j�h��U%e�¦%UF�2�ApF��F(�²��*��\�Q�Ym�ar��Uq�0QTb-�m�UeQb�1E�s-���
�`�[Jш�*�lq�ȰUA��TATPD-,n%�l���2�+U�"j"�E-�AcmLlm�5Ɉd
�2�����mL���*6���Z ,T���iQ�X��4c�̪�J��PPq�\B�.X�La��Ȣ�Z�Tb� ��aXcFK�"���KZ�P���)1����Z��[Z\B��Ur�X�`�mm�(��rܵ"����FU��R���������U*Z��Pb,Ģ�2�J�Ƙ���	��g�E{�~�b���蟜��J��p^�l?^���D��]�@2��� W�e�:��~�^��W3��$dE8�*8�>��l�s�R��ֆO��O+�:�7��͛��}\�qb��nzwXs����T�M:�Ҍ��u�ѭ����4_�۰�'!
�n��P'�X>�)�^�A�ktl�>=�v��r��_�ۉ(�`�D99��>������U�	$u�j�	 �ew�~��<}�9��{�C��/(��)Td]�d[��~8o���b��$�,��դ�:��P ڽ�@����A)�_��u1�2��~;�����.�����C��ާH]��+|�/8nzw{N��|�m�cuf��ڗl��Z4��";��R�(6rdp,
ȶ�ugN���9��M���S�ٰ�}�j����'��	R5#Cc�W��]�Q ������t�_��=n� ��^c�H$v��..�[�a���1N�^:�u�1a��a�.{<�G�F��V�I����N�P�#L)����>�y��$��۰tVev{IŦ���@�m_s�n�`(7NT���c�{}�r`��{������F��t���ł	�nv3z��Hz�`m��@�U,�tH'�}۷`���_+��/��I�y�P$v�ݟ�u�8R$�*2.���<4�՝T;�x\$g��'�{�n��U�g��An�����-T�@���?C!ad����t����㹬#ս�{���n:${7���^�:��roթ�&߬��ׯL�t��ݧ�__~��#�6{/�NVƹ�q��8m����e��?��|��eN���o@�of�<k�v얙����7]kE�i�a6����n&�nD;j
������y�lfE�-����J��\�ۊ�yq�9��<N;mk���:�N�����$��p�F���g�d��i3��<��:�,�nu�t����R�rR8|Q�l�#OB���p�pXi7j3����bۮ��q㧶��ۈ���k�����m�D7=�k���I���4��j�$7JXl����mk��,`'�3�۲�l�]&�w�������xQ���j��D���,����@�z���G�x��/m��۷����)I�l�����<-���ߦ�?~B }ܐ WGu��kʒ߯��%�L��q���@�uWuh#�s�	?ީ��K������s�!O��܅(�U�Q�=n��{ÌjY@�� ��H���Y��wMG:���H�e�8��*2.��������)�T�ʕ��S��  �K�蠏?]c;��v�^[�	\W|�}3	hG��:�&6���w+��b�]8aGJY�\3Cy�;��N��+�����=v,�	�՞�I&���|uL�G9z��?-�[��`�=�<�[�f&"h��������=Hg�Z��~N;�x��fIXp���v��D�a��ӭC-X�͓�4"4�J�JÚ��t
i]n�<oV�j��l��VQ�s{����z��
 }�~� }U��].NԄ��8�w��ts�ƁB���gGY����� �Gz(R>~u�8��q��&@��۾�]���}C!?>�P��yw��$�;kr�\���P�WT�?t8r$��1)L�D�E��ؼ���w��;�kk�|A���G�nv�a>�婖�y��.�O>n:A�pX��l���ԝ�':�;sn�px�M����Td{����A���G�=��v:�UG���آF��tHk����4Hp���v��A�z^�vI�����H�{�Q'ݙ�`��Y�m��݌5밠p�c-2�/<��H�<�
�(Fy�mb���˴���W>�{q�mg��zX�Ȋ{}�t�M��E��o6n���Uz���9�$Sm�5x\��P�WK�N�ʐ1�)	E�$q����ٕ�8[���[�� ����\_����ۿ5����@���t�)�L�ݝ�޻?G�=��=W問��@�>�($ί�����CM��w���$�u�S��۞ݦA���#���b}��X��Y^2]��go�y�#)H�b����M��زA;��@�$�'}Q�c�*$���3�� w{rB�b2YQ�:���:��kɝ�|�H'��뿉�w�%ML�m�ʴ�݋	j���h��!����d��ْ�$�X�uc7M��C������$��D���p�ci���ܷ�S�;Y�W\O�)�6�
��R�|:I�� ��Ü�Tu�0��}��n,M9�`S��!��$>��^!�glCMz`���_���zv忽C��+fl���1_,uOo'�VI7�נ���!�w�� l��]� f�;;p �������:|�I 3��@��ߎ��(|������:�*��M�D3����e�hcT6o'k6�h]kW��|w6�V���������)�L����y�,�G��BA��T��!K�fWu݂	�<�M�rS"d��B���+�Y]��n��]S�K(p��m���:b�(�C׽�bŢ��<�o	b�e�K�E����߀�MS*P�ټXivU� �,�: �s�T	k����4K14gm{K��Nu�������	�}��$�s8OQ��r��n� H�/�j�@�1��f��{hQ'ws�_�s���S��{!���@��: �O%;;>6p�]���޵䵏<�=҅���m:�uӚ��v�esӯ#a�[�!6'BQW�7GJpA��T<�`�N��
�TŊ+3�1�%$Y���PK��p�Cn��WͶ�޻m����-���cqú�sEs��ڢ\;��
v�]�� u<��uwa6x�c��ݼ�8�qcq�BFr���:PŻnS��^����Y�y��V�9�;�0X��,��R����xl�G({>=ok��=��:˷t�js�z���ZV�,�3��ͬ���ʬ�s��=vyX����^�.��%Ƹ0����v�8z��>����ϪBSQ�ڈ�8>��師�H#ݙ�XZޙ�ݤ��Kݎ�$ޮ�@��퀠�eHIp���{���^jx�Sm^��T7~�� �'��ý�U��5��wˉ���Ӑ4dQ1':�_�&�slY$�C�0��~��+������|Iٝb�e�H�1(�&2.�2�l����N�۷Z�W�Q ��αd����G������Oc�B�[���E�SaAFoW� ��o���U�B����@P��/��{삯�a��u�?���3� e��8�y0�Ƣ֌ݶ�d;=��݃%� m������c-�v���������u�d�Oޮ�h��0Թb�L�*��-�  ����2�������@�:4w��8�痨X�>m��LH��˥�mc��Ry��ޭͲ)>moV�x�O25��G#�g��mZբ-��^Vl�J�+m+@�4Ⱦ����O��nm��xh~&�k�����~���$[��J7vv�z�}Z�$��������	9�Ρd���h=�d�H����P]�ڊV��$+�i
� �o��(��[=x߻θH(�Y���W�h��{�)f1����K2[�D��p���8���C	�&L"���"9W�ڵ�s:`	0��04@tZs��UTU�8������r����v�!��m�P�Z�6��ˮ����R �������v��dn��L�$��d�!�o��@�1����}]B�%׺�M�=��� Py�h
����	9���7��z�|,�μ�%�%2�9�tE�l�$�ۇa�g+;�{zc�'^�5�#cz����F���o`m�!�
�)��E��j%�:t��ٲ��'�Լ�]���|m-h�6a�@'�oe
���4S��J]����D�%���Iz�_�v��@o�Z�U�ޙH��zT�m�u{#�k�Gl�$��b6 A������kE��`��ʩ�Eo�T��Z�P\��Ff�;D`��;�$�LA B0c��R1]I�n�Ŝy=�n��N�׃q�7Bp����ߟu�̮�uSZO=u�3���y�SbŞ~}�\�[�8�f���ʔ0/]�H6�UEt�R��i9��R���pOg�
$��o]��="���:��V�8$i/z�>�I����$��{�5j����h>}��  ^}�Tz�-�!��i1�ǯ��@���;�����]x�ru�@� ���ۿ�9; �F�'"{�7�����z��G���}N�%�1�L_����<�HWtW�������rhG�-O�	�ʩ��߫�ߐ]w(��~S.��鱔S��J7C�/����|o��^�Ly;T�$	�u�~;�w]�rs�@����u ����[��^&�קz��b5[�%��T�0Wla�\a5��9a@�7��$�܂6 C���A �{v�FN�|=2��I̝��A��u��#m��!�J{A�0T�8�Ҡ�H$G���`�	:a�Z��7�5h�7�I�(���u�mAO����#g<������1�H���	>�w]�	:a�C����c-(��W��[�۫ʂ�z��#f�]�A#v��~���x��U�xM(���\��/s�]h��ZsX����{�H���ADР|��U�r���H�7n�$7ja�I���W�>ȯhs����/� u����=lz�vc�b�����e0�iI�˸�pz���fq��.;��d���P�w�u6G����w�]e�6�,����6@��M�q�\zOJ-��ef2������
GZ�4M�$
�K@�K�"yrХ�MϮ��������f��kJ�N�E������3 Ox�H]�q±WZ�SI���ۆP�݀�vc��v��~����b�>�u�,B�A����Ą�4�p#^���3,�{Qx���hO��������ť$חr)�y9���p󞹵Y�u�S�Nĳލ����/��tN3���x7��{���v1(�ǹ�=�-��6����k�|Q+!���Gۛ��m�b�U��X�8lO����,h#���p�|։�K����b��;��Y��1y�~�_R��Uk>�f��um�B_l�f�nj�%w�]�+�xh~Ә3oiѲ�׷��jťl<T�Q�9��a�ќ��V�y�κ�;�ʈ��{N���n>�������c=fe̴]b�PO4�v���j����MxY�y��	�zD�$.9�ևL�I�ہI���wXڵ�[�%x��Ì񊴹��箯:&��w�=}F��2}2(cy+ ��\J��y�v�b]�&�}�+��!]�$�Q�����Fj,�F�i��BV�oSs��I�I���M�@��v���y\*ඹ�L�1ē>cn����}�z]o�{'>�l�O�_TY��vD�/qX;�>�)�s<����EU���,�d��iZ�G.Zb��DXcS)�,�3EX#0Ic
�����(JLJ�0�#R�cj�j,Y`�³)Lq�Vҕ�B����I��LD�m	R�cm�T���(�%He���
��r�+����֠�$�b�
"Ŋ��%f&2�e&0�1
���f1�X�r«�lDQH�dT`���F(�Ԩ�Xb[k��(��2�RƈũEE�J0mZ)i*��3��-*�̸��b�e����q�V��5��bUJ\�E��TB�UYU�HҋQ��ʆ2�q"0-�V��2X�c�eV*���i��qZ��%�J�T��!Q�*?3��4��M��q���k��v�̊th�zfV�%��M�hN�pxM�����R	3��m��:�@4qìr�v��n{kv��n�&c�Ay�:����X��#r(;�i.:1�bn�.�U�5u�Ukn��➧�v����z��2�n���ญ��۶�����<<qz��^7�";Wn۳���g�[��H����8�os����|/|��=9�'3�:��F�u������u���N��8-�E��l�^^0m^Jx���cN�k��ׇܶ��͊��!���8���r{	Dgu[k��ue�4���"Yz�N��\��Z�c\l\M��)�l�⍻x��N2Z�����p\=�u�u�;��<�)�-,-��ˮ�8�)A�NNj�_[��������f׮N�&�ǶQ�b���1��8�n��nXܾm�{nr����F�ڽ�a������z�lE�#��Փs������n
]�K�v�=aћM;�8��r<mn�xSeqk�6{y�+�v�j���l��[�s��u��D�;nz��v4&8��Lmɷ#������Ӹ�=d:;	�y��[t���*h�Qtcv�[�H�5�!�w�uI�8����`2�ɷO=<�w\gT�tq�w�M�u�k�G�r��#��#M�{<��h�u�|��_7�z�<\+��b�v��x�}��ۭ��f������܄��;ӣ�d�S��=d�����mi�<�yx��onۨ�Z�S�(��v7m������L�Q�xl�p�M�ˠ룞۵����\q�:S���N�Ï:�и0�Gm�4�۱n�Ӎ�P)6�����s�:����]��E��:�]�����F�&�]��#���3/���tS��:b�O�R�۱n֋��v��uF���P`:�]�g�����잹�Fv�ۆ�k� ���W|���xb8�H�z��������v���&n.���6���O&���1�B�X�78�v^�q�x[cCnۋ���]�7n�b{��̃�Z]q/G%S�5.��n0���u���;v�8�p�y�x�:�mԧn�"6�l��8���ֻ��c�,#���n 	-V�����]�y�w=��5����{�;�fh۝�g�9 ���g���px��G�y6j�;�7@��0� }2��<%��:-G�{;�u�[��w�.]�����"������d�q��%����Ӵ��xqK�s�k4��E�7A�'aoZ�]�^��L�����c4������ܾB��� P���kA�v[(�{S��ݣ`�k왂�o�m1�6A�#��(w���tl+�����4H${{(Q%�G���>���﬎��6X�	*���Oh�{r
$u���j��i$��h�}��(�~B�@ƐPQ���:%z���ǣ���쯨�o�;����%+�{���G����p8&2҈Վ��
$����;g�1p�,��ցR9��
]���ʭ����Wչ�2˰�b8L���/��ê���@;e��jz9�ûc�ճ�����}�o)i�e�K�w��A&�� �O��3��E����g�{��!@���@�+c(�`r4�n����� �v�=�y������۬�0�-�[|�f�0�,l��l�Bw-�ΝS�1�x�|C��%y��a���7.��W�	��BO��za	 �gm9������t��Ff��m��I�Z1_I��H��۲	>uݏ6:�����o�$���Ɓ��;j�w�$��f}�7z��8�������=��6�E�nݐF*�j������}�k*Q�D^���6�Q��6��IMv>u�{�r���h�M��вuWc��t?bzl��T�fư��!˗:���=X]Vn9��^{9cl�+i5c�???y���1��G�6�a�I;��W�j��E�Ua���,�$��ݥ��pƚ��\�>�c}^���I������I�v�X'㦻Z��k2ud쩧M������F�1��zﺬ��[��$|�u�7b�қ=���y�M25�͡��*�%�|;e\��;����嵐�����=�5�7�v�z���C�g���������{ۻv	 j��@�G�E M�b+�8�CjguXf�t$��u`�~�]��?.�q�-UE�2�k�N���w|2H����b7�BH9|��&���-+ȐOe���U���A"��ѽR{�u6uW���m�.�r�3�9wp��[��r�:���A�z��a��J����ݐH:kr�$��E��z<*8�o�����������o���d��J#v2�`�R�>e��:��ΥC��=� R]��>�ǧܗ�f��*�)��X�%��遂n����^-�h�]/	�>�(��N4	yތ�����1�C�����{5z�<z�����9L�@�A����u��Y,W�)]]�tZ�M�P������߹d�=~��.o{�o��&��iYw���u\�J_a��t�W=k��{�(q<��H�l�H������eM4	'�}۶ŪF3�/:}�-���|h��{n�Ngs�r�3���36�u�vke,���Y�����Ƹ������������S�1�>��j,�(�zh�I��m�!v"��ƍ]+u�sN��{<4/�n�8�I(HpQ��]X,�^U�!<�m.Y��kܨ�/�����e��� ��f.���o���d��J#W�S�T	 ����Ղ2�,�Z�|����]�p$z߱P$ow�ŗ�Ԝ���i�.��um*̈́��q�V ��~$����w�$�6�b95ߨ��岈�U������	8i�� ��u�$�}Kr��j���^�Hx6�HP$�ݿ��6�b�}j�!�z_�f)_�E;�u�J�����~�y����[x�GO��N��bz��6�r���~��=�2���0;k���p����"����x��5�c�lu͖,]v��!�qm^h��[���k�(u��8��c��/���Q�#�:.H^ڪ(�C1�@�v{(��I�勷��!&-��s������	��7]��g+�M���}w �hQ�`}��F,���3�ʲu`�d1��+;���n�9ܩȭ	�Me۞�tm�� �:�6ͻ0�v�hI�κ�Q�m�1��s����ThR�H�v���]�s�u�N�������r0c1ӝbH7ۻvI'i�*7,�so�N��8/ٻb�gf�#�3��	��O7�����u���wlXMv?�q�Bp#ݷ����!�BIBC�Nۯi���b>������d=)x��ݶ� j��D��~+0X,�8BSo��H����w��>���^�>�if���:�	y��;�m�j���8�͏�=�ɥ_<���on�G���=�K�7�� =�E]���y�|z�8�R��bb��n�z:z�[Ll��Dڷ4�[�Lu�_��۽k�{�������4�u���}�,���	o�W�~�q
�k}�0,�U���x�R&��� b�Y\蓚6���8X�G멅Jǘ�3Z��U��&:�p�w�Y�6f(߮���X����y֥�wZ�Q���Ak����Q�n�9e��j��7��	���[�Q6�y��#�\/b7��u����ۘ"q��#$Wf�����7��|H/C�dܵLçخ��@ ��D�~�{΁?;z��.2

"��^Q���{!B�0�mA$�j�_�o7���;����1���y�l\��p�ӎ�72�y=����Z t�r�_��*y��&�=h +�IzI?��;ۧOw��}A��==�O#.����y��^�m�;�냠9�v���m��okR6`Q��:w*�Y��@E�v���"I���R��Dj�] H��_�o*�͓�i��j�`�95ۣ2��WЂ��:�I���=V�u��u��y�9�cqH�b��,�tH��ݿ��O
����R�죔[{�.���밠,��.!������Yt0]7�	��J���-�TQ�sPy/qo]�й�܍�:�W�G�;~�� ��_��_��?gw�4�h�`C3
CFo<d���I���^� ���d�	���6:Ʈ$i�������<��\`�E�=��z�����4�}��>xr��������Py�}�����k���_,zA�:��eƍ9�����r��M��u:��nm�oh�+p��K��Ǘ��W/������	*p��z�� �ٽ�d�qs��
>Ɇ���$�� �(G�r�-W	m&p�HLf)���1�����uU��{� �~��۰I#�@I�Y�6���iyU=$mf��"q��*c�wh�I�^�dQ�w:�ˌ�zݝ�b�#9����"��3�Mv�����vH9��h�E��5�gT�4a�B�z!�m8]�Λ��!άY��V��en�Lf����PCxz�����ӽ+�
�<�^2$��	�;F��x"E�(,m��d�{&ο��Wk7.���g��)�%��� �󯈢vk���۹���W��L8�&T���`�f���$3w&��:�Qs۠�w����X&F@�Y��5�~�,�~9�xh�����_:�6�ᠻ_R����3���%!7��A�����ם��}C�*��A�L������>�ޙ}��}���d}))]�t~�ׯ ��@{�{}��O���'�w��G���ջ��8�l�;W�:����ù��	;��k�ַ��H7�θ���w;�Hog���98a�!	p��=��I �vm���U؇�b�1��2߯j����K<g���Z�/3�_.���S9r)�s�\��6�I��-uo=ҏ|�����O%+��4��_Y80�"�G�dkuv��im��
	0�ӷVTf5��nm��u��c�#ki��*�� �мn���5��vh���<g�n��������N7v��<�2�����S��k�7cn{�p��c7g��n�Wv���m���@\,�4����n�p�a�`��E��v[����;��nI,u��V��x��މ8�� �b�=��3�o;���]g�6�O�ȫJOV�Ѣ���I;���T6m4^�r�icm�v��g�����N��	a6Y�+�R���=�Q �nuXY4�ʜO��n�ri��:w�����&(P@�Y�M���9O|��10�u'�� o�~()��_*Y�8Gu�����N�V`Õw@����:'�~;�λ$w�(��g���: y{�ٱb�w���/����f��rf�̓�γ3ABL��<	���~$���,��
Z�6�9p'�]9�����1�`ƍ�;W�b�'�r��O��x��y�~�7�W��}��`X$���Q��ƪn�X��"�"B�!vd�6۳9��v��r�I��5ݗt�����������a���&C"�[�A �vm��u_�߂�����Թ�vX*�{�L�~��`hH�	���]�E[L�of�i���6��ua;����q��^!���=u$o���3t�'i��JUm�a�H?-�ꔕn�������Y��i̻��[o���+�
/Lۿ�������l�}�s�/�����%Q���� �v�e|� �ӏ�f=����?	���	;o�Q}��`��a)	���������ð���]�O[�T#�G��1
�&yc�;�}]��e_JI�!(�G1mPd���t�ܘ�k��ˍzL�� }@E~�@���^��s�����s��,�+A��!zZ����g����n1�c�6�2k+ф�&]��_≰cG�>;W�Y��7�_C�?<�y��i�;�\u�W׊�F���27��`a��~��ŋ�a�����$i��_H��@�	{鶾or�t�+}Y�ؑ�M��4]k�F��t	$���1{<������Kݍ����!Ϡ�kzwx�6��$��R�7z]:!;�Bh����ك=�MM��㹣��=f�l<��2��O����-��=[S��,�.BX��۾���&ip�A}p7`�2s顅���OV>��+"7�����7tR�%�U�w#��i��z��1�j+�n��f<�\��]�&�=.��v��[�����N��:�p��$ �5�
����81����N��0G���`���z%��&��˝Qw\(��u�B[��[������uќo���ҶK��.�,���s"��;{.a�/Wq���=�C����� ��m�t�e	vtWjF1��Pl�ׄqU��;Y��%%�z�X�X��:�<&���w��>y��^�{V�.��;���dRö��3.�!��y� l�v��P��{���_7�v>=O(�
��nw`�ѻ��q��nɓ�؅P7��U���9z�xe?UG���'N�-Ԭ�w/wv���>]�(:ph��p��
�WWs��pƻ�}�~L?)�Y^ա��ȇ���6{�=��Y���p,Y�������i	�/r<�|�����)�s��K�9:��A����U�����-[��z|Ǻw�������f_<p�;1kt��.����W)��R;�:����q�S�Bw^N�^�QR�ZM����;S�C���Unp&��%�;�㢬iy��!�r�f�8?��<��]{��_�/s��ḓ�P�������D#n3�PX��Q���ɉ���Vc3
@Re�TYEAb�FՅUX���P��s1@U��1�D�ITcm�J�B���*6�Ҋ �����q��+%j��`���hY%h֦8���K��˔�\�2�B�����jB��jfd�+PPURcS���"+LnPm*���P�.���* �(���Dr�r��Kj��[1�1�Dc�W�9�YlP���2�eİ�PDf5D�R�TAˌ3-b��Z��UTb�q��m�iB���.6�e(Ppjai�ʙV��q�Qa�h���[hTZ«��j�*���Y�j��.1 �e���q
�*)�p�*��%���X�k[EXԱFc�Z�������b(�(��(�l���-mb*��ʫ2����܅EF�E�
�[kmҍ�����5�j��#ZV��a�\�ʔ-�eQ�����A{|��ت<�y�%[��"F�2 �f��l��x���0�?9�PF+�u� ��-�ӧ�4C��Ż�E�o��!��PAXj��������}S����?�-��F��t	��αcv�sش��C�\-�iĚ�6��u�����b8;q�Nܝ��0J��K��nfgy�e�5�`�����8B	���I�����
��r�ʱ3S�]^t	 �W�葳t��L�6�1�v��X�K��ƍߵ�gB�X> pN^� N�_*5<����j߳*��l"�af6�!�ڠ ��ͱd����Ǚ�kõJ�A#��1@��ΰ,����$l�؂;�h��zÛT�B>�t	��ٶ,F��zD�j`�AW�|�8c��0nl�����j�9�g�o���pq]��Y��.�첱'��ûD"c������xݠ�[���=��$-|��@����D���I��ʔ�m3��À <q���9R�T�{C_����T�ONׁ�NAA#.7�e܎�rn�c.�zێ9�%�3�)�
M�]X��߿���C��������N�s�_�o��oC�G5]���p���$o�:����6�Q&K���t�UAi�������z	�{3:�	j��(|]U*=��Y|�	��|P&D�(ѻ�������撋]̞;@|��ٷ����=�$�����",`��O=�H.g��
�r� �*�R]o�SW�+}L�̆��-�@P�n���J��$L���K�FM���چ+k~�i'�*�!R_��5~��R��[���
�n��8����5��f����>sVb�53�z��v���BK����y��X|��λ��0���T��/�z[��N4LM���v�=p�7���E["a����dNE7SM�t�e�`�ؒq����ª;q�{�p��W�m�q�y��%����7]+��m8�ޗ���ζb�6٘�r,�Wݰ����98v�ݎ��˅�J�շU�0���*)khڐ����:�N{ru���V���`#cӷ&y�s��^�J�u��v�z3����q��Ű6�|�F/Sy�����:��p�Q����OOod���v?~����@���&��3�~�d���(BI>��v����{�ܑ�m��7�[�����_vՍ�8�D4�|w�)�`���ɝ����_sѻ[�ͲI?y^�~>7��w�B����|�wJ^��U���j$�b�Q� ��ZS׿@OS�(.���H��c�IW���� L�FX��w�;W���v����ăG��I�U�:�E�s�ν��K<Cڛ�ߐI���-�5�kE�f�a�j�nk��n��|�f�遗j.���Yt蟉�}��$_�:Ź<������'!�3�_n�����
�##��o6-�����Mè�����{�p�֜m�hu�Gnk�����j�'��|-r����e2������P�7�14	��|fu���j�}��N�[�~��L]�,\[�l�^��L]��ۤOlrg���xg�����]O^�֎�;|VfIPto��A�}�Q&���`�{�~�olJ�f�yo��3���b2�mAv2��� ��]��m�s��y�e��>���Hy0�Ē���Z���D�,32���K�Eޕ~=\	5������,����;���l�r;�n;4Oò�@���&�Jޭa�e	ǳ}]w'��<A#*��	 ��u��]�b_l�q��}7xWZ5�*�j��U֭��b3�2T�k-�u�* ��C�k�����߿Z���Ę�:��o;vŐI���@�����W�۔��s��4
 ';� �߸%�7�0��Ǻ2b~�#Kن�U&��ޞ'�n�ݐF��:�	os/�T�P�?<��� ��&&�f��b�$=�$є�Z��1�m���<yn�T��P�P�r\�ø\*#Q�;�Kw���v�̾�*)�f��pvJG��]-J��P�լT���v��@ wv������:����n���_5���R�m�$��j��(1��Iu�5{6��ͭ��ş����eF�,32�<{j����P��-��q ���� ���1�Ƴbl$5�o� lX�4/F�sI��s�s���jN
������_������������E�挮�.������x�ǯ�wzW�{<4oL*r�+�=^IG�C�]����c��!lP�S�~,kXo}��u�޲H:s��wύh�3A֍�b�����nB�I8�6\����H������ͅ�k���o���wӍ�ckē	f$[�v=�r1f�c$��u	?.�q�I ߷���:�5���槫s��v&w���^%�6�������/7���(V\��i:��ml��wv�k��֘�-���?f
vꙏnЛ�q�E�I�ߺ�(P�~;������z�h�~�/X���ܡ@>'�~���X�8Sls��ߟ���`y�\q�[�F�������Ʈ�=az�X�Ӟ4��o;�����W;<�~ￋi
�:
$�E��lAv��N#��yp$={�(��� L�4ډ�w��^����i��Z��(�)�V�O��J�P�=u�Vw�D�"��y�"j�j(�#�<H7��vIU!yՍ��a�(UE��@P>����PE�%$�2��m��V�v)�4��(A��v	;�ع!】*�~�2ρ04�a�>y�~	���YX�.�d��z�Q�fm�`�H���_|y�ǂk��k��Zk�ܳ��Py��r���s,u���H��'�l�"�ݼyRH��DYV���Ѻ~���c��S(����)�.��g�����F�\tY�69��n�e���gW�kqv5Y;t퍎��u�,�<�6ֵ"�#m�8�pd�JE���ћu�㖻;��<��ۉ�&�6[n�!7\p��c�7=q�-n&k۵��Sz����v�Y�4��.����#�����ku��J�Cu��\�`:��Jpf5!�-���I�k6o��>؝��Cs�W$�&���L����!oYM��v5̲X��]ی� ���f�!0A��eo��I ��:�A;ޘh��SwJ��P��������-Z�m��L��G{]R'��E������)�@����<����ݟ;ݯO���@�"e�&�J��d�o�WȂAŻ}����i{F�H=ٝv	;ޘhd�#jj(�'A�n_�9�x���n���A?{}�o]�?fzn�3a�ڡ���Nw�[��RN,R�|$��(�}�ٯK�>��rT���@ ׽�Y�Av���ɭ}�L3Y�]em�Zj�u�r�K$��$&��zRtv�ε���W��������<��~� �w�R$�~��P�����|���ALմ�
�<��'���T���p]���@�X�����q��}NLY�u<7�� �:h�9���sJ�s!&�]b�Gσ990��<������7�Ow���Z�*'�_O�~=��h�O�z�|D�9�딺��g�o���Q0S"]|{u�I7y�Q��5�BT9��w�;�O޾������.Bn&M�����σ2���k�O��6�(P$o79��w�~�z1�e>4HZ�\lEb������nРj���i�W�?Vt�D�כB��y���uy�b�{9z�=�Ɂ�/8z���Y�Mu�m.ûd�Y�y��n|��n�R~~{�E���.��G�$��(�A��꿁���L~5������A	�r��8�Ä���M�P)<���x'�~��Ă@��@�H7��X&J��:�3��h������!j�}{�+�H$��X�O���A#7������& ��j�ow�C{Zq�<;�ӗ
�7G��	ͨ�.�фר���oSN�,f�l�C|=@P����
Og]�����)D�L�tw9�ɗ��~��>`P6�}�@S����/d��:�p������wu��KXH%�i�ɻ��^���yAoU��C�ތoכ(�$�f�ذA?m��G�_QJ(�����.7Jug�����J���ۇg1�X��ڷ�=�w'o������,۳h^��h�I���N�L4iՐ�UF��ܔ,����F��ͫ���r&�H-9���-ܒu��3� �B��r�i�3�>����nnԁ߃�f���]�\34�~�~o�����n4�5\������:A;�λr߹{�Alc�/Ln�~��A����8�'j_X��~�_	�N7��x�뛨���7�mLtN	+VWv�t%���x��h~�߼v	^��n�Kt�nB�^�1=��%ԫ̇�$U����+{^��^_!Evm��N&
d@��s�������K<�d$���]�H�~�(|H�zqyEm]��D945��M�AD��cH�abm��vӵ�q7ӛqҜ���J�O�~��}{v��Zq�}����A�^�@�	�zq����<�� �v���u�r�Cטd�4�.���٭w^������<O^���)=Ƚ�@��V��P ?<���!e3�U_N߯����܅�Rp�B������=5�A���nT�=<�gmà|��בּ���xn��/���sǧ̀I�[��?7}8�$f�K�ֹ��/�����f��0�5n��L4��λ���W��'��t�����A �;:�Ͼ�w�ʭqے��k�2C��vpҥs��k�4�p��W����<c�[.H=�m)��k�3F��J�O�������{sR�%zm��Gv���W���x0m h0�~^k|��JӴ&݂ue�697-���Q>eՀ L+G�v�g[�4e�G%=U�C���ju<�+��L�&Mc��S��Ngo���}ٿ�᝚��/9��)S�y��0$"�O0�(�b���F��Y�éL!���U-����i����DB��f�yCR��Ky/��C�l	�N��Y�,ٮ�6�He�j���5��3���6v��J2����b~�4Z�W�5���h���[�[����;5��-'��#���:�+�$�X�.���oմ6�i�<������2oP� ���=-.8yF�ώWJ5.iy���������κ����=�ya�r��U���*��=R��)��ͺ�W��CF\]λ���I��3ԍm��������p�D}�K����^���m��P�4o��?j����$�e���������%�uh,����O�g{��<�ةy-6�Sy%������j����l��Y܌��a��v��,����6"���;@\����u�!����/�K무������ܺV5U���,�
cx5
�%���@���b�ř�ty��Z�g96�m�>�d�����6����	9r��g���38�9]��¯����p���C�z�V�y#��DgDc޳���u{q���{�W���r��w�3��e���+F#*��\aQZ�m[j�.1�J�ťKD��*����E���T�� Ŷ��*6��+�%�iR���Ii�nL��c���HZ���5��JG-k%�S�R�iDj�kKT���W-QEq�\Q��[(�l���+Af4Ĩ*�-ZE+�Kj�"ѥ.Z%L���*֪.eƢ�ֱiVV�b�--��f\��E�+m�����5m�Eq�e��F�e�e��\���"�#�W(R�b���ڔ�����`���cm�R���64��)�DTY�KIG,�[r��ԣKE�֭�EE�V)ѭq*`��Z�Z�U��"�J��EKEL\er���6�Lh��ZUP̹��%���h�DR%B���R��E�X�s(�m�V����l�-��*�b[��Ī�E���e����iXį�g�m�7�.I+͊y�rn��0n�6�Y�wav
��N�4c;���n������j�ɋ��ų�	��x�;Ӫ莗�d�i��8�T`�v�s�/V�N��i��8:nlFz���<�����ap6��Y�u{lq,�p��4y{p��4��֝P�5<C��1�N�ي;n;�(��Mr�&�7Z˖�tWbϞ�n�K�� ��YL�Wt���nۣ@6˗v��C�G�m��Xכ\�8\/'�:�ۭ�9�p��Rm��|c�s���ӹmSݕ��{s�ͻ[�<!1�tۡ�q㛬�sWe�m���`�����2�lxM��B�Y (���wdQ6磝�v��9�W��CQ�l
�8�LP�fCƏ^���ks\ɷ���]f��m��������*��v�ؕ�uǖ�"s�e����X�R�.-��Z�h�w0`c:��vD9�N9��.�%W���d	�m��;d�t���py����-�l��.4�\�����/s�`�t-�d�ey�9��P�<7gF�tW��v�|7Rsr\�䝗A�8◉M��[�8�p ����kX.W�Ef����Y�Ds���v��W\�����6�f�ls����	sh�u��փ��e`�!�\9��� �v^�햮�)Y�]�x������c��]����������ؽ��õnn��ls�ۇ�r�3��<���I��prE�;a�v�m����C����-����kYw[��v�SGZ]�Fx�ٜ�m��j.M�g�9Ɣ;v=�\�.�$o9k�����`ۦ8S6��I������v��gK<@Fa����z7WX��\�K��n��6��<���&i���'vqI۞$��"���R&�tkeժ�-�S�ؒ�<q�ݷ\�!�v^8��K�<�0竞܇;R��&��ȧm�<��nP�7f�N��oG�н:�5� ]��-�pmln��Y:�C��A����;�+�[^��G[�d.�$��q��u��v��P��\�W`.�1P�fwc�;s�j�u�;�Nr��m�XWt<e�8�XϮ��rs��ϯb�ާ	�tpc;7<�z1Wg��[v��<g��)m6�ۧ[��\���&5\�q��_��p�9�nJw[96lb��M�a���m�tg�A��{'�;k3C���3
Li.�8�����e�p眭t�i�8��.z�[�s���H�\j��n1�/.�6���u�@=�ow��l$"	2 E�;�u2	7�zh��>�ΫF��Վ}�y�TH�y�Ɓ=�X�	(P��66V����u}��ޝ�w^R<��ē}馁?�s�X ��9����/C�MR2�p���!BL�hH7��vA�Ugq�y��-;@]A��s�ʓ�r�yX�I8L���-�����nU�v>4%�N��"�R^�vuN�=@|���m��b�'j@h�������[7�J�+9��I ��u�`���ʉ�������Т\�`��ci�A��,�$�˵�6/M�b���m.�豧�C��������v�#"m�}��$�s��$���ʊ�̘����of_��벯e6�(�f����L��f�̪���_�_eײ�T9WbM{O��!nw����5���3F�յ�o�s+*B�*H��A�P�]9So�r�V��.�������T��{�ES�g=���t;sY����G�dO�Y<�K�����^�Y �m0A�=RGj���>Z	w۝b�-{�~}�P8\%���P��/*���7w����2��~�~�D�H�?r�n�<�|��~5u�w�ل��1��p�V��B�����M	�O�'�%���A�~��}�~�@��!H��{H���#s� p8�H}n��m�;=1v1gWV)�����.���c|�[��uj@x��złZ��$�G���Z�n��^�,	�~�@�=��.���+��	5܆�O�̴��Z,��~�@�~��r�@?Off�Sj*���/U�y4�j��B(�+��I�^�DFg��R���﹃뮧�/�#��`���PGU@msȯ��w"w5>�9�oZ2M��ڬ�dC5U������͈�G�@!^׭{��zoOi�)+���n�E�����~;Cݻ.�E@��6A�j���Ԗ|H*�m@���
zyy��aS��'~�u�S���C!-5B��u}F��nϙ�]�G<wVw3~݊����݊��}�]���9��j<ֵ�3C32:t�KW��;��bb�<nz4���\��ٸun;����݌�J �gqeP`���I����^���xb���+��;B�w!������@ȋN_��U�t�աQ�����s������2}'��T�n�K�{~	�\9N���@$��X�(����y"c�lOn}�w�*��x�A�nuڽt�`�I�Lf)�v_��=����Y�X
{�rT վJ3����ں�s<�����f0eA��J��lO\K��x�c�ЭwJ�ۡ�;a��Z�����SzJ���Eo�{n�v(YƄܹye;o�M�}+`!2#ʬ�޻ ����)��(���/��ݝ`X ��~�E�eI'�(���+��z�̶Cr(SE���sl���lC���v��m6:�J�Ӿ�?�y�F@Ym�GF�ʁ�vmX$��~�@�������ۿ3[@�<�
�� E�b���&]��j�g�Ǌ�ɛԒ�i OIʗ�5o�E/w�kpa�����=�{y�[t:�9sK��}�<����w�@��b,���zz�>/� �<�P��׹W�߂pFS���������o��޼��Z�*$�k�B���_�z�;[��=��
�Rm�!'!:;�����ob�r�9�W�	�@��߅?C�l�}NZ�/+/��p���ݽ^���ފ�;�D£���m$��=�K���%�z��W�VJ�s��~�����<�훒w�����L����[v�E\���\�՟[����(��[�� :Q��-p�X{^�M]��݌��';s3�n��{��og����� jp�W�L��;+���˴>��c�y8�kp<�y'n縯>��G9�Zv�lX���'����u�ط'��E=�/>�$u���v#�XFD�9���;c�yz.D�N�&�[x�V����:�n'�bs���s����7�����ڳ͞4��}�w���/��ֵ���~�BV讴]d��w�}����~$=ϱP��sui��'�7:�Ń�$m�b��{��d��$So�Q ��v�ݼݿ�H�~�D����;B�]����c��[l������`&�R6���B����w��O�2���{,O+}XAoڨ�z�G���e���&�/z���J=D�4�:�/\�~ ��<�F�|���G�F[�*���R���	p]�<�	'���q\�D�݌�t��H�ن���������)�9fX��Ⱥ8���x���Ƥ�Q�c�� c��m1�9�!��#s�wٺ�`�>JDLf)����x>߀s��P�V�廾z|u���'L�F2��G���^�|Y5�n�)��P�����M5y+��s\9љ䷆�����m�Hv33�v�뺌s�����}���Aq���Ʀ�wٔgg]�{�ʙ	�}��߯i��pbO�a �3��ТI��lY��j�=b�n�f��I7��H$�7:���(�^5�[�{�1�y��LCb��WĒM��_׊�̑�`��j{�p^�=�f8���\��s�|� �����un��b�o��4��ܾTB��C�2��s)��0�f���FGC
�i�]��;��Q�[K�s���Ok=�֍t�_�{x)	p@̄�3�޹�Q���H��߇Q}lvdk��~��[��6��fo�v�Άڅ3�L�C���W	���ɗ��[�ROr@|V�kE�dt���t9n@3>��s�a$�i|�~�m�X��k�A�A�M��ɔo;���1m���7x�w9����z��aoQ�l�n�'������msc}2��%���+�Dh.�۫h^mU8�w�q'�����'-�����,I�$L�}@7���w���8{,�A캻�� �j�A?^�q��Nv���	oݵ;;Ц�B(��[񨶫��'�禍.^����By�:�2��H'm�|	��N#���g��y?xwul���4��[��]�0�l6ͺ�`��5��'�j����~??~��]��bx���Y'-{�I�Ӎ C}-�P;�y`X �6߱Q#��8��|�%Aw�s���6'r-�^}d���#q|����Q8p�����g��w3֥R �u��U��$y�Ɖ#�Ȼ|��u/t�꿉�j�7��E}�U��7o�v۾��z�.�/v�����$�����馉{;�1���t�.�Z�f?y)��⾌�%/I� Nd�)��Uyw���-�vН�^�B��jz��*��~��t-�^_��N�i\�f?fq���b�s=��S<���u��Ɣѭ}C��Q ���n��oj�=w}�	��-�Q��~�9�rU~�%���0������o����%:u�t�J�:5����J�!�����ݴgR~�~}��;6����ꯙ��w�
�@�om�>�=^qmFe����}��U�e��(�S&�/z�XK�j���v-��$g{ ������߷�/�0�{����=�FC>r����(�� ﷶ��RλZ;���ۚ�F�
 �	ٽ�a�6�"O�p����Z�غ�l��yZ(Ps�ʐ�6X�?{�Q#_W@B,6�q�����߬r׶��[� v�k��гj
$���	#�o�D��ɋ�m��VTo,W{݋�^�~���~��}̛r�6<6��sݮ�/����l=�]�'��M�VI�b�9B�3,�ѻv9M*�P+L�Ijm���u�z���Y�<�����ا�m��\=m�bە����0�/K�Bu=���Y����;�����˷|���ëoo7�&2v�j���S��=�����v�պ��.ݬ�[���v�m�qû9Ϡ�g8�U�|��f�8��q�zNv80����vH�n��ź�ۍ�rtd��vv�����oH����guo3�[.N�7+��Y�g<؍]�@�i���k�^4o<�������3�4d&�B	>+ރ�$y۶,H��r��Y�v�z�+ݴ(A �om٬��S���N	���1��͵	��Ч�ϩ��
a?^�v|�E���O/��� ���
3�h| 9kܨ	Ӻ�j�������;��v	 ]W��_�ƙ�����,n����N���U5	=w�$����&��-���X�� I����d=���$��B��wj�삏{�����>^���$vߵW��o� ��}��9�Gn��<1��V�L���҂D�k�����x[���)s���)�\A߷X!�l��A���I����I��P��G`7�bGA~��݂	�~��#	¢l4 ��O��|H�ʝqV�"_w���{�%M�N�]�u�n\�{�"�s|_+uV�{T�J3*�6�w�
rز��8��
ú�t8j�s��O3�K�iNڀҐA��!
�Ӻ�'��[����/�(Q Th���Z����՟V��)��l��p݃MM�A �nO��~,5��Β���_y�U�$���A�삉�{��G8r���y'�� ��»���� �77(P�A���YU��B���;p� �s9xFVgق��%ޏkEϽ�i�񎵽E;��n�<���lW������_M����^�q��BH���ܚ����l��)˚�)Ǩ����c�������p��ymp^nA@�I��ۿ������#�/%�v�
�鵴��M&�r5�;w�V{c������Qw�Oy�
=2� ��_*=n{���y��<�Zfu49	���Aޚc���H|)Ueu��˭�(٤��NF�їSCn�i� js�ց�he��/g/	W{e�d�=�A�.�3�%�o'9�����X�֖yYsO����ɟp{���])D���w>v��O���uo�^�^я!�c^�Y���_9�6�ϭ"�pWnM'�k�ѕo�̛����z����[�&�L�7��}۝��A��os����>dM�zO.�8���H�m�����b��خ�k��=2��ۡY�������M�6�o�Z��yj��P�g�b��Fs⺤Ւ�'��ݶYw���!�=3���pqq��,��3y������&����ܰ�M�F��</t:)��m�y��풜G&(^�I�jL�\%X�rf�꽓n�y�ʚ��~$n��Z�\󦺭������oJ�ZՁ1�zi!*�Xh�pA������^Qb�{)
�,��K�R��6r�x��p+8�U�78��2xXk�s�y&�ɡ�=�>��Fl���w�u�ʭ�����ú5�Bh�-{r}��
��76���Ǧ�n��V�%f�M��M����Ki�m[��\*!v�cu��5��,�<����^� ëZb�*s�K�Y���{�ƷȌ~ԟي��q��Si�R*M��T�t\M��g��g�e՝�{f�W���C/�ݲ��Wܦ���Z�٪X��8R��H�ke0������΅{}�Y׷����g�u\T�O&9�|�k�.:0�'�ؖS��ĭ��⻒�`� *��^J� kwl�|�ܴ�%zil<��Uh<L���G��XG���J����<��\�r����)P��R�A�e�ƅ�Q2�TKJ�(���J�dV�6�QEZ���3��
԰��ʌjUK"�*+Z[�LUJ��F��QJ�"�B��EA�,�Z���-eeUm�Qe�X�V+U�J�
�1fS�*�°E�Ɋ1�*�嫊�c�eZZ�6��Q��J5��Te��J�Pc�kIX�KlPEm(�eZ�Q��*�lZ֖����jҖUP���R��*
��%��*U�U�[%1�im�-e�%����JUkZ�[��F-���V,+[E*��EYZ�jU��m�R�J����2��2ѢZҢ�hZ�FҢƥP��-��fe�m�
�m
�Z�EX����֪Qm-R҉V��[*ڊ3-U�eZ�!V��YceeKN��]�$y�B�$�yݶ,�gd)��l��p��i��}{x���y��s �$P���!A�~3��מ� �qmh]O�i�J(�p� ����#-{��p��q�=UpP����~�E?6�Ns�����t�]a��N��8���֞]�{t��x�\�E�b��,7k:y�tw߿�ߤƹ�] �}���D�A�nuY$��~���^��ez�I;��`Y��Q6Ip����b���N�Z�]��r����߈ ��ٷ`�}oܨ��	��y_o�{��]���-���cj���'-{k�Is�%�١��[@P	$��E���I�C��m1J��#�Ժ���"���F��ٝ������j�~'�oe�o�����!��3�L;N�zEK�SLv.Əzg�X%��vE��o�G�uԆ\�Ӿ·�,l2YF{͔�a��c��շޒ�����w.ȭ��S��ى��ؼO�s�|�Qh]�;����	�-�U|A��k��<-ߤ�ɕ�B�������dڮ�݄�i�Ȭ��)�����6��~���Q5ۛ�6cI�n��o��� D_�6�� ��^��ޱ:o��������8�|����Fc}ޡD��+�э�隺���?9_��$=��(�L��ë[�����Y��Q6Ip�����������U�͹���vЕ5�0�������G���u�6�h��]��{���ͺ�{Ԁ���&�e� N�e
$�����)p��q>[��C�u0�J�B	>��hQ?o{6�����`�U^t	$����9�۲�0pU�|"��ɥL4��_��V�b.�xA��n�]�L.�Է~넷ۄ�?\��*Lv�݂�nʸ�m�\�֬exU=5��*�볭���n����Gܑ��b�"N4�c����3��\=s�0v�ۆ�x9�ݜ�Ϡ$ݻ�z��'�5���wG\�9�C�8�3Ǘ�9Ⓠ0�m�bAq�n8Sn�r78^�lu�=�X؝ۋ�ktv��v�ގ]��n��8����8�� ��X-�Ϛ0�E��ݝ��������,�nn�pN:P��W��p�s��������r���L^��m�Ք&��H�皹����4�@��o�2�N~��ڬ�BOL�~�Oj
��I�@؝���N�e}_z=�m�
J(���W�/&��"������$o�(Q?�s���۪�L~��m����Zl��c&0`��o�W�w۝b�ėQv�Ƈi�ά]]�h$��I�ο����TM�Tn6cEJ1WvS��N�t���
���j��7����� ��jՂo�����L�雿����n&����t�|�����jT�Q'�~�wd��7~م���J�dWY^F�����m�y��<�3�Nv�L���gs3XR#L(L��W6� ��{���@7�� �k.�����v�H�<�F����"e��63��C��:M�J5�6r��Q���kwi@o4��]h��Y���\w�	���U�p��l������x����n+R��V!<�W��5�Tr�;��@ ��� ���й�G���M,���$s$��(��yi؂#C9�� y��h�W���Ν���gs9�f���wY��].�u7俹綮:�q����";�����7��Ej���Q�~�]Jiz����Л��%ÂG,�@�����u  _g�]����:�����׋���盤�=�j��ҍ���ڲ�C��1v\e;=�Y��e��-��qZ^�i���}]��<�>vR��/���E�T��%�����Ib^�B"IC��v��qԈ��f>�Ր ��kt�}�-��1"���v,Z'n��y���{�ޏn>��ؐ���7A#;:��AUM_V0�ֲ�z�wpF����p8n-�Sq@�:�E�F]�2��Lx4vn��^G.��mh��]��gs�u�Z3��3ތ�f�w�P{�ǽ���Tеî�������j;�ql�H�Z�st�@#=�j��N�9� �SsZ	�yXr�E;ǹH"82�H �^�]� Ӽ:w��}�mz<��7�K�FD��g�|c\�U"h��=�<�Kt�ǽ��;P���=~�%��I4�{,Q6��y�E��U}�=wŅ��r�D��*b'�.������\����B�5�e3Z�e˔�[�h�����%�9h%��eyҐ�z�DE���*�(��k{^<-o�����X�bt����l%!�Iv�{�읺�N}t�z܍)N�D����زl ��;ū ul{j��o[�mo�T�*a�KQ2� ���F� g=�� ��_']o\[�D	����  ޝ����w�Kr�p��1qeC���[�"�:�)]� �Ӽ]�p������o���\n{FW3����/�G���Z�\����ö�.�/.{aѨ�}~os8�b��A�lҼ�w�L�M*{)њ<I����[j����T� @2SsXO��V�A�g%�u>�{��0�����G� �3�H.���\��%�d�$��M��N��V�Ug]����<q x�Bi\7^��.I$KQ?o��W��Dq���� n�4���=�1]UKU� �=�v�=�W3#H�%�l�S�DN�ٵ�c؆{�B��	-~�w`�8t �g��o�������|��Ć�l%!�w�Z�y���<8��P�v:}x�#B4��vD@�yäV�J��LCjE*������L���ު<8q$��e�-���$ �vڪ�h�yw�
��;����8"d�\6����w���d���W:�g�>@}����8t F{��E.�̲�b���yx^;b���B�qY�'���vZg���D>݆u]�j���H�ӫ3��֭���t�@��Xv�`D��w�ϫZ��;l7 �&'��G/kv�v��������۷���u��϶Δ��uv��N��X����q�IS�d�����Z{O-�팠׶r=�܊��N�pn^7g\�=�M[T�<>�nWv�m�]b햷D�{6�.�cF�#ݜ���v�L��^$��['OaF�ǎ
�{{S���^���Q�g�����];�s��N��������.����rt��n�Wf���u��)j��oW�������07%��ɕ|�π��� =�j�7g��M��w�맪�>@x~��n�ܹ$d9	j'�{�-_�D^v�o�����"�*�h�D�z߉ �~�T��I���ջ{����mj��,TK� c&��T�{�J��@�r���}�u ��n� F{:�E��GI��*B!r�-W��5��d��W�=W�|,` aZ�C��=�֮� c���k����=g �͙R��E8(�Nfرh�|�v���s��q��H0�������� }���
��]q�=lW���f@Y��tҩ��
g6�uνP���]������F�	�����r�j&Q)�dw�9|Ȥ og�Z�@$?w��w̮�U+�^��s>dE o�֭+�:uK���)�Z>n�|H�2z�{�Kx4WP$�N�7q��3*Xg^k4
t	[W�^R��M����3�.�ォE)+�]^\��S�m�=oޚ������a� ��m]����dDU;���f;�?V���]��rH�r�O�h�^ڿ� �\������~t��UU�ݠ ��εvA����eU̲&�SD7v��u��~ݟ�E���+�H"4�y��[�o�#�����I���أs%$6�`��˴��yb$��a=/j��`Z,�ν�Kr�֮� ��d���*{+I�u��a����"#ea�as=�77cg�Qqo�n����+����npp�v�>���z�i�(�N{,Q����ۖI8�ctӤ��vV��{�֯� �#ǽ�Xg������y��#���7g����{3Ԯ�;�������|"c�ϸ��*�l�(�՝0G!H�3LY�̵6 x3�����w������-#o{�Λ��5K�,^��|�R���e���~i���z��g�7��B<'(����56�����ѦdBrLS���@��;V@��� �����#!Ē(���<��٭�E���w���D�x��X�^o5��}�kۙ>T�^�����o����bӼ��F��[2�.es�$@�Ԫ=��FLdrɠ@+s�w` ��� ���U�]�[�C�{#�G�%��$q0�K�G[[��W
�mױ���s9.���c���Ͻ��9��V�9����n �<8��֮�tKލ���ޘ%���n�A�:�ڕ-J&dr�r�,s�j�d~���T4�z����\�IZ߹�h$���X�l$�;�ä�<�~�3}�Gl���TZ)�����+� r�W���D�;π����Զ��=S3 @1$��N��=�
��x�6����H������� F�w���^��[嗔(ȷ��PU���^�4o#fлSk�)yR/��ʳu����#oB���Fm���9�H�	��ϭ���R\`KR�l�u��&�p�|�v��H�I<{�z_B�Z� ]K@$�7�G�=jՐi��vN�]�/�����?����r�����M����l��Ș�{ny������[c������S[���.&��+�|�> /sԮ� wy�Bv���؉ێ*��/[���m���z�lG�nK�L9��jlf���#y�@|�Y�֮"�F��wh��]/y���/^�t�7c�b&ܧ,�*���}j� H0���� ���ݗ�͙����=j�- k��v�����%�T�������'V�*4�սJ�"��o;�ky����~�^���??�H�εj�*ޝS3 ��IY��Ħ���g7{��!ӄM�!>̬�vA$����l��f~�E�@�$��H@�� �$��@�$�	!I� IO��$ I?�H@��B��p$�	'�@�$��@�$��H@�z��$�IO B���IO��$ I?���$��B��`IO���$�B����e5���>�� ?�s2}p"c�9�@     (� �   P  
    �  @ (         �T����%R%6ک	QQ�	P"���)E�&�!BE*����
�HUJ���h��vjJ�H�AI�  �(   ��   @  @     P  (            @ $��@��9��f���j��T�'T�x j�f�z�u��^��U�9C�� �:�ﻟf(��u\
=(�mc���  {�|�t^-�`��x נs��n�y�u����'����}{�  }����;�:�w=������N��*%Ru��  � @ @  �>�s4���|Zy�^�C������ ;W�9���O&������s�{�����}� ,���j�j着R���]�   !��}c�hR>�
z���%}*�h�y�Q|Ǽ�E�{�`uNv�|�u�03��^f���<@�9l�l�6��  � �  

���T\�_OD��u����C�\�v�� ��E0>}�TR���t|L�94��1�����))_. �
R���^�r��)�}xI+�  )G�JR���%JR�^�� ��,����
<�J��c�(�iI	/,��a�J�M�}��)%%V3K�)JR�l��nR�����):Ǟ@��(���I|  �     (  |����@��m ��� :�{� � H=޸�B��N�{i� ��� �t!�t{�WҪU*UR��   <� �9 W�  =�{���^y�7�q����� �w���O 7��� k��n���Q �Mj��   |     (  ��}rT)�`qd �d }p =f3�sB�� �j�� :{�4yv�AQUJV�  �>G@��s��꽹� o�/tn6��W�a�1���< z�2o{��z��ⷙ���`t| ��@
J�L���b��(2 h��S1R��D  =��FjRJ4ɀ�!��*R�  $�H)�JQC ⟧ߴ~?_�~?_��6����x��>d��.�����A��Z��H@�~�<����$�@$$?���$��B���BB�		�������������^<��Uc���p�CZ�2�ܙ�)�d�ν����u��׭�=�{IB�9pт�f��d�Ҳ�&o^&+x��79�����noNM2y���v�;A��}rc0r�qn��јF#)�'��vЬp��yct��ȮC��j�~���̀-��� ��:�%VΎ��if�dr��� c}b&��`�W:H����#�������ڌ{eŁ���l0����mq%��N�N���w,R�wfY_�8Y��1�'I�˱�!�pf������Fk֎PD� ������(�p�n�N �Xh�#K����'m�ţ�lgWm�.��N����d�X|��skE
����uv��l��]�� yf���4�xlo��ZR�X�ʮmOzƗ������K7q[Ds�թ�>4AB�
����'F�9@X����+�l譽ISb�BOz���y=��v�n:���op���P/�u�2�<�9(���c}c0�K�����>
��w��LO��UD�g�\�
��Y�8��[�wstȘB��N�n��5��M�[�7�F�:�᧧k�6RE�5��	�ۣz��&�Rރj�c����/;�V\� a�]Qۀ�GZ���ԇu��N�k��"H��n�g�C$,�wk{�b{=�N30�w"�Q3����j�)\�pïjp���4��$�#)�+�8�trI�ϧH_H(�sg0x-Ǻ��!+V v�z�^��"ɾN �M��ܐ� �dYrLc��+��+jM=̴8��i�K:ɴq������=U��'�;Jd�F�멕[[$ƤN�t��r���,5܇BY�E�j���f7�9���L�j7�Ft)���
���tZ3�< ��9ݐf�V���q�X:�1�:I����{�]�ۋ��.������X���Y��v%�f�5�%9�h�wh��/v�4���-�v��ي�ݰ,�`�"!�ƀ�t��
T��ZX�v������;�hzZ��Oe�t0l�~�6��]#$j�xQ��	j�.}kT�3I��u�4`=
:�T��Q�fަi�Ǉx�)FAc�� ��۝-�_�V��vXx���XѺ�˜�1�x�I���*��V��M���賀wfˠ����m޵���ۭnWi
c�D��م4V�Q��]���iY�I�C���]�e2C=�t�(��oX���~P Qv�ܭ�(�ܡ��.��m�V�TN��,��׏^�o_X��� ���vi�Zۖ3���l��ۀ��q�2���Q��'��ifF����Ns�,ki�l�][��p����p)�4kz��1:{�NON�$�3��[P�e�ض��PP\�!�]/��K��|v�4�O�ׅNa�a��VIӧD��-�G�/������]+L탱��17;�d]a�����^��D^��vӻF!���L˗Y���Z�Ӣ������ �븦��6���Y�.�X�w>��鮴v�C�+8E`�N3gӎ�ܮi�՛5�Xe<��<p�M���>��z5N�W��^I�n��q�U'DbM����}�\|8o}O-H�V���;��,ع��*Y5��e�5;)I��5���K(���U��t����&��R���� N��jћ3�N/^�\��tQ�B�Ʒ�Ɠ�W�p�N���ѳ�;����Ӝ�P���kǻ{\�,0@�xO9�%�i��#ZNM;
Z��vJ�1���;��⻶�'�#Y����7�`Z;#��$�a�a��ڞ@I�!���h8�����e��H���ǆ��Z�w,{N6��P8D��!"���K�t���Д/�$��i:��Լ�C�N�r��ˢ�7�l"n��\���Ϋ��7zcn�Ж����[Y@���hl�uW��%uv��q�ù$�+�r�l��#�YL��ζ<)�����l1��ѫ�a��'��-ׯ��</#/�!�
���=ym/��:�ymcM��Co7l�����v۫'`�.Q ���*���W�m����m�JOjS���\ۼУt+4s@�z�3f���z�܆v����Dm�b�N��0��T2��� u[�E����6-��[23�,���gU�ϮXE��v�@�އ~x��(+x�g^|�sz��w�â�����EN�Բt���}.t��	�	��ש{I�V���I䎕�pE��wkvhl����q�4�ဂWe��Owi׫BN<�'�L},nk;�p�X͖vA��qݼ�Ώ~��N��8M�Ȯ�͵�0�Rp��v��yS(��R(�y.���eҴT�HTt��f��)�"Mv�:.>�aNuu:���c�ͧ�=r����W[bȒ7�V���L��:tŀ��g!}⠏'y?�i�A�7��z4-Ŋ��%����q��㳜㬶N�Q�9��Z��o�Ɇ��>�EGZ5�)�M�޾
����&n���2��jLI|�;�����\E���
@��u�L.�ٺ�˕"Q-�t�����1;���<+��#R:���.��V�s��|kN�U���a�J�2i��X0�5qƑg��hD����l��,��2�+����PG�.ލ��VN�xw��S��5�u决F���Tݷ���y�����SM���Z�V��i`H�c8�!�;F�ﻣ��jӜ1�dI��0L���0�Y�{V���S =�](0W`X��3�+�@K���_&���-�o77	�>�.s�s�K;�R-�e#�t�E��#�Muפ.$G^l���c�&���n^2���8�m��"�+���bY�^�7.p��՝LW.�EN]5i�gp�����{�lhBSթt��;� '�^�Z��kA�h�tXA� ���s���4�(�� �5K�z�Ӊ��_N{e<�v��ݛp���Ջw�lO�U�^ޱ�N��T6A��t�$��lb%؊��mZ�H=�f=��oA�v�/^;*Vq޽Ďޗ�o�e�ӄ�jዃWz��n��[��W)#�4c1r�&��|���@��Ԯ��+}&��.�q�7�gQoQ:��g�EɈ�݃<����F"�D��ӽ�ou�����8�h�+��m���B�^�
:��d�o�s�8 �cM�7�bԷ�`����h�ߴ� Z�Y�K�������&P���2m5f�E�9;{a@���������&l&�]�Ŋ�5�c�M������q�[��n$�f��8F+l�n���*�u�F�_cc-��A�Jn++QB
#�w�ᕽ���;��[�u�i�z��	Y;:�za�ƌ�5�%�j��3Z��ה�e��+9��9�喢���:�+ޛ��<��cNv� tn5�@}L�W�t�N�7�k�NY���^{����]�Z^��;���c�9��3!�G�܃� ��*��WK\�p,y�Ѿ܊5�<�cq���-�gN���"c.��f��m�V�!�5�rgll��q�*{���D'���U�o5�2ц+��0�T��*�7@|�w���2RT-I�°V�Ю��ܢ���k��ǈw�3�;� ����_jK��9u��N5`D�92���1f��-�ǀرOb7Y�RI��G��[�N99[�Y�;w{V���p>S�z�v�"^��y���Vx�u@ r8nm[�{i�hnh6��I� �k ,�%�m���J+	B��٠]���&���Ѹ�J�V/�y^�V汿�杋��@G��`��d|;��ߟ��~��p-�άl���k&Ÿޡ:��{wA������4v3"2wF��ޱn�H��XRl�J�ǟ@���� J[�-3	�F	 `��9@��b1�{-�Q���u��(�E4�� s��C�'%L��R{s��iC�+����Z�!��!������p=׹G��n�t���]�Ȓ���t�;Ro�.iW:�9efv���C�:/��wyKa��Aښم�ۯn����@؝�"γ�0�Cj�����l �R�ȼ����l�M'���8"Ț���#Z�����Ѻ�����{$����՜�t��w�fҲ��wBݱ�*,W8
'n2�-�,Fz �ntO��FtuniN������'�UD���I��GS�m@cWS�4����pƎ�p<���I��ےh*w-8I�c"ֆ��b'q��sb7��{��f�Z{6���c��T�.pUm'h%m!Wp�ҧ*��L���	���Ou���w�I�������qs��/d�
`v� D"y:ƃ1�D�5��<}�x��ƣGa����z���;��!J�����)+Zm�770m&+�-�.�ψ�rqeޙp��zoL���#�5��]&�y���	�W;��Y�'+#7�-z����W��n���Ԇ�o��<��v3��ˠ�&��v𫻇 �mnΔ��D�Ï=���{+����PV��e�m���Kd��/��L�� 9�4G�� ��ʰpqΐ���999ުNgjXM�g.ω}�d����ΊA��:���-'�z)���+J�`�e�s��j�Y�Y���,�ɱ�����X�g2�g25�z=�qDֹE���b}�&���a+qQ{��V�Ӓ.�Hˏ8����A�=x��߹�&��nv���Rq���o([\�J-�I��료�O�:�kM��a+��o���=���4`��2�N�_�h�|�0e;�w��+X ��	y��D]�V2��{%9&��:�?%�fK��S&���kC�<��� .�ih�_���c��ǝG7!���5�1X�'�@h��|%�כ[�3����u}�A�\;���w����f	��\2%V��;����zjQ>�X�R�+�gTKC�ĜȎs�S�]s%�ۯ{�l�LU�;���ǉn8��
b�;t�1�4<�Q^��(�hK�sw�i�䩤�j���Onk�8n��3�87��Ӂ˻���O!7T�u�='=�ßQ�4�B�+f�p:dђ#����ـ��
^$:[�"������M�m�T����O=<)uŮVa��Ԏ�d�N��H�^�n� f�g|��3r,c��#��dn�`�"�=���`����>�^�%zT�m�n�: �p�8h�c��>�׶;���iZ��ʱ�!�p�t�'��=�uݡt���4�Ә[��B�%Zv�D�^�p$*�o|�&\��Κ�mCy{~}��s[�xۓ7Y�R�"�ФK9�3�K��{E��j���u�חI�4)S���0��\9v��M�1,vk�DQ�ΏqK����t�R�o.t�)�P�P�Wq�/�y�S8wa��s�n ����������M�����n�f�����B�b9;%�hO��.�㌻�l�YUq*3n���<�2���w�����w.�ww�8ON#��Ncֲ�d��p�+&D��9�H��UY��@ˏ;Z5b�����n��sI7R�c�QU���G�v��nیΣ�fŜ�4gj�\X�Dhڕ�i�#�03����n��SԎ&sf�.Y�iS�K�C���$�Q]�
�:���{ptz�)Gn�<��m6�Ǣ�=���s�/���F[ ,IP�m�}(w;/L�]�7�3n+�DRq��.]��-�U�����{F�;B��d'5�:�]��ċ$d9n���G�#Z=0h]���e����u���K���È���7�[�p�b�7m�`��(��8�q�ݻ��cF跷Soa�>�R�nۼ�}�BH����Vo��h��N�����a�CNဵA5�pp,�2����@
V�A�p?k��`aܼӒ��kp��iZ895PU��[�5;v��@�l�8E�t�}���ʅj�ay |V��D<I�٨��{>cC�Ie�I�z�s�m��b�x�����S��u�4<�5�ǲc
�)Q�|��Ѭj*���J��6���gI9�Z��u�O[��۫��w�]*�r��,���;y�Q&��h�	���r��=�M�-�p�͝���@A˼s�d9H.>��˪�)��V�{M�y���L�ż�Br&���cU�:�.������ZtL��7L�[#�Ů-zb�K�s.�].�Yյ�R�A<.mӵ���k���2N�|�ly�i�����YV���\ye9�д���ڰo`�� 8�&�м�w.({�D��0��v�ujљN��E[wY�n�]b{7������k��(��$��o�QNLv�S��S$D|�w�Vs79�Y�ݧAƱ)SV�(3��e��Zeo��VlF�z�9��E�£���:��{�K7)��Rdy�7��)l�F܅�Gd�n4��v8�3�6��ƝRאUC����m��A'�p%Ԣ蜜�fD����F�����)ӎT0fA���ބ��'��w�ᓣ)�~:ƶ��o����K��y�d��ȥDPVA*j�v �Sv< ����t6
\����[֒n1��_�����\�u��,u.0�b>�����J�(lg�\�{oL`��;�xo�rfʳ}7���Hs��b'���.�ώ����*4w>��{�.��~@� )AI	E�'�� �"�	�T���P��XB) T * ��RIH ���� �$����*I�aH� P���� dE$$XI"�@�,��H
@I�B(H
��R ,�
�BJ��$"ŁXBB@�%I$R@"�����@ ��XI$R 
��Y	T$�� 
H
d�� �, R��$���$!  X ,��V�@!*IJ�!%d�d�YJ�� ,� 	 P
I!
"�H
@���)!HY@Y)$IAH�$X�d$"�
 @RI?��BC�$ I/���������������7v3{��"�h�[����J�x�Kd�o�9k�x�{Z8�n�^�D׋�a��mW�!���R��%���ҐY�i������]��^�.��G������4nʛ�4�`J^#b��Ǔ���x�|��v��"�Z�Ａ'	�v$�X�f�nA1��kMZ����eJ��&b�H���r�(rt� �m�ά��!���;{:J��*��j�H	��t��͊�f��Eu�/��<��g;���ʝy_+A��_b�k�u�X7��_���7AU��j�N 3��q�	
�>�C��[揗�*�����gq�+�WG؍�Ռ�3�H=�WX3Z�J��� N��H�>�ӷ#ݭ�]�:�xܡR
%��6�(5�@���8��>�Lu�A!ނ`�&u�nW���vW6}��y�:sG�K]����yZ�����h����~����{�F���LJ�zu\���N�-�����U΢�R���nBv\���y�T�,vu]K�G}�3�q��U(��o�ӻ���򛞬
X��l��W�A����燡��'FyЃO�cyS��R�E�=��(��q�גF�,'7ʺ��ii��lؚ�&CX�Z9�9_����Ǘ�2��j=�����#��<Sw�
/�ʺ5�(a�o� ��fM��S����{/kh�Վ˞�h��|�����狞�0:X�CX=�poe����WZij��(qē�O����#�ڔ�7��,<L(G�Z�q��շ9����Y^��Sk��C��T��+SX]���s�j���u��Ơ���/;lC�����{���g���
���7S�Fn�J�J���O��Y�i�Q��r���%��d�rǱ�ޥd�<:�t�I
Qtո�o*U8�ty��x=}:���`����f��jK� �=ܵq���`��z���Y��b���W�\��a����������V��峺o}=@����4��f����c�>�#����|�>�Jҝ[d��ݎKz#j�s<(��w���\��l�
����1��u�F\S�^����ε'�?)�os�(mv��Qbm�Wz�n�v����V��<��Y�����A#�������O��F�����Y5M�W]��;�ɞoz��jupNw�L�W�[�;I9�.��<�����ҸPS^mވ�)x��;z�/,���:H�2մm���<�5$+O���7�h�����&�};|��N8�?%v�Ö�� _Tݳֹ�s��,k;O��7w���l��*���еq�z���^K2�T
`�~[/YW�rY�o��v�:��$�+��Z폠<�:�7��k��L��3z�r^�e��D�����ٶ�/s�(Hi`:W&�^��o��sr���ӭB��r�{�p�2$���zc��zm�ی��}��磎��͉p���Vޅڮ�M���L#�=y�U����w:E<�F�|^���r��tgE���5�A�wҥs��>��¢>��g�|�,Er�X�D�uK�e!-L���B�V�g���}�R�m����O>�s�sx�i��=��D�&ӔK��FOe�e�Y��%�-���ԌS�u;<��wL���r��Jj�ϡ��%�h�����w�V��h>��KsH=��Qe��^���s׶���\�ھf`b͢D��	�F��U1�bk;v2%��	/N<T����w K���!�A����꜇�� I��<'����z;�	_l�am��Q���rT�c1���ŧ�[�V�ތ��v��V�8*�!�����oh��f�]�Ճ��N�iX��zX`��K"��<��<ga��F@�����%u�|=�ʁه�r���kD�\����9���A�S��+̦�R�x��*�s�����r��gj�.�e���LTJG9ow�ĄH#��������8<�2S�i��|U�xr}}~k�ne��^J�J|�y�0Ne��_}�Wlfu� �P��<�`���)�n�vad>�y�fu>��Z�f���ݓ#�2�\�v�j��|��uSq��_��x��9u���p�����<u�1g	�z�8Ι�$�H�yarn��N>�%�4?=�Oһh�>�!xw����N���ۏ�y|g\�u�:7�\2+�Y��I�_�ԻK��z�#e�����t�w��ۋR�t|��=��x������/�j�£Δ��O\;hV4�&w*���o
��.J���	�����/G9�ٶ9�C���R��.�֙y��*Uՠ�{�չ�S��w6�pp�O��U�ԦpE��V��/�3���j;�B�k}������gA�zm�C쑇2g��̣��uSi�K6���	�N��DE?��I��<7<@����Q$���7F6�mQ����E_>û�%�ow� i����1�9�<�I���N|���:k�97�б2���PQ!��U�ۋ�q�z�lޢ��UKD�^�q2;�a�����X��}C�:-��ݦ���su4�o��pex�^=�yY�.�'W�g��|{N���iՁ>q0C��{V��Q��8����Φ��#��z��b$N�]�[����3q�f=���IV%��h$'k��/	���P��l���#���;��ra��ו\�s�(N��A��d��G�:3�'|���M.r��|��ɝ.V���=(��A�x{�ʦ����%*{�Q��w��vt���u+Oڌ�i19���mp��K��yv���O�^+���cV�,	1Bm�@����wYw�p*��$�p�^��wS#��!}m���A9�蛫�vB)C�.�fɷJ9��6���w�j��$�-���`�3�*Iح�^��<�0`2��ϑ������Z72K�=�e��|���n�y�J����Y�t�]��,J��}ֽ�v�\�9��f�`�uP�^鮷�Iz����=�iH0�$��Yq�6�$��OA��ᾴo���$��ɝ��=��1�Ȯ�s�����o_@s��d`��wg�sw]+�̫��N�3N⣹��S�Z�l<$�3�*~�4S_;s�F	��NļKs=�`�fwJE��}�̾3ᮑ�ͺU�z5�J��cc.M6T�-�m
.�ľ�=�ɋ�9����胞{�s�u�wz����e|���>�l�������˺����fu�o�eqǎ�3�z>~~������
��z��r]1AxDM�:%�$�P}zw�����5L9N1�L��U������37��m��J��v�[�/ ��>s��N���ך��-��魑���{�4t�������Uk&-��GWx�Oϳ� {�����6{�Ѕ��ILM6��-�me��С��z�4��8Fn����Y�p,:[�c&Y�����A�A�=W�V4��Q��6)Y��u������
� �#�́�m]V����Mcʘ���?R�ѩ�YAM��L}ĕ�Q9'fy�|XS}�g���qp=��~��Ƹ��C�쯲3�6? dl�z��s��}�s�{�煮x�wRTT:B0��X��/8&dvn9��y-˜�������"�fF̠�9��Eooa�~S��DI��5��	�۩j�8���ED�Yٔȷ�r�A�',��:�\d�̥OU�p��OP&��꣆�]G�tװ�=TMq�%v~�<���vn�%�s�lI�e�>e'%�WWܓ���C�)�I=��u[�0�p��>Oreoh�l�2�R�8r�l��Wu��}�j���d�S�j{���x!,��&*,<9`�|��rK5-�4�Ӣn3���]_m�b�,���z�Ԥ�/sۨN�W{��Sk)j[6��K�uu3]�f̾T�]6�w{�����&J=k�0�{=�4�ȒsA�D�8���a�$t��^�>CnK|j>>\Ǽ34���!�5�n����;szNK%�S��OM�1���3�����ُ��"�dԷc14{�>�7n��RYMQ��<|�ЮϻrU!���:��3꼩�%M��fy
�'�ο�G��<s���1��87�݉�j�X�A���\T�bC�Ee�ǹ�����o�h�Zu��,�4�ݝ�sVv������:��c�K������� u,,�*�Ҳ\����r����{|�͖����T/~�zJ4�f��5���ĵL��v��JGkU��])��]^sOo���;[I.2�Tn��4�̲�R�:�wFCR��17�ݨ�ׇW�5����w��l�D�A9#�[�c,�.@�B�Z��|}����*-o=�y�d�����>>�ډ�q�ONKۣ�o�{�2���ϝ�Q浇ᓡhɏN��O��O>�Y���~���.����{���F2�����ɩ�����>���D+�
��}r���������R%������׊�N��4޵.��H9�h�B�����<��C]���շJ��&�:�s��r�vf�L�*�N��*�	�GԎ�'k�#����ѾCF��z�g��^�&S�XЂ���<2v齛˹wh�����b��=�pv]�1�n���x�[��Cަ��a\�ɷ�Kn�l�{!��z΁����N��Y\���Z��j�m��n���z��գ/y=���J�t=9���	޻ҥի%�L�}]�i�����Ul���ֽ����9�+�f�92�c�o���<A{��Tn����zY�Y�]e��~'F���{��>[[,�}���e��fh��m|f�mx����.��Ǫ���<�5��q��^�v��&h{�A��O%�K��u;�2�/M�����r�@K_S��~L ��;�ܿ=�Z}��Td��UX��j�!�����yb\�	8�礃h��sx������C�skBչ�\�@�Ju�q��ыy�
`:��צ���)�\ʤ.����;��KR���z�7�^7�v���ՠ���v/\E���瞏�n���J��nҷ~�*0�E\�78X�n�H��X'l�`�1g[#t�;eV��ązAf�ܿC�}�ռ�N(�I"�A��)J�}�͟i�S��8K��X��������C8G,\w�iw�3�����{w&V�= H��m䠸������3{l�Q3��ǣ_F��6���=%s�ؾ���xWp7u��7�����J�b��u`Wu�]�^�*�*mM�{q�Qk�Wf�� c\♝��m�6v�־R��m�鸘=8�Q5���l峘���"���7�mmE��j���)�����_��]��M�kV��uB��6췑2n�*��w}��}y2�ܧrzL|n[n/#��7��Wr�V�8���w
I���h���W;�\o��(���:��,�r�S��o޻tk�k��d)�b��B�����V�~���g��olHNͳ�GEڷ���y��`Ǹ1�z Nu��4n���q��^B�ZԻ�A˺���Ż6�g�Z�Ő/���x����d.u�]\�0qμ��8q��[�a�2B�zu7�_y)71Ed�F��[aS�/67r�/5RtmK��Tsׁ��ƥt4�{\Q�ܘQ3�Y,��꽝����M}fV_4�we�U �;&9o(����ױr�j}�.����SA�Lm��s�ɯ��j�=M뛨�Ujٸ�fDEc�.�M<��e&�Pd�� !����mq40' �h,�5li���˾cYC}��Fu�*_s�*5�}�ut�JU�5WS�AF��r��2o&�nl�ۙ���WdƎ���w<2NS��(�}�:�5֘�^�c5����iwTjt݃������q�
سS�m�1�p�����};��F����{���7�N.-��uß={qs4����V��[m;׷m3��x񯻴��&a~��e�m?I�����nisNC=z��y����]�.%��p�1p&�aIU!i	{��<�"�PIV[2Tm�[��s�a����R�)�� 5��×a:0���C�Gc��38��ތ�U�gģ;D�����Y�P��eAv�Z�~߮�#.?9����p����*��{UB ��t� ºuT��Jr���܆���5���Ƣ��T�*��7�� ���a�Z�G}��4g����#�����v��(�p??^A�\���p���w��ޚ63FB �߇h�޾}��f���7�8ʬ'���n�$}CU�y4*��ß(�ʄ$�3x跫��Ub�43�Mëq]X̵#Ł��N��yj����/�B�}l���c�*�=ݕ���qh��N̐�b$Q���x/FI(��,`��C����uɛ��г���ʻ�}�.�L�^]D/)�y6X�la+u���g�Lx��Xb��)��6��C�����[ܼ����`�h+��6mG#^�]����.u�!��3�GU\b������-�\D�����\��P�2��"����b��2X&�W��l���xI'y�;{��,p��9_��]�*c@/:��Lu�|���Q�d��6��#)�"P��Qp	��v��hY����sW+)Va��r��]7b��7�=��oA�7��+
���c��y���J{��c%c>b����y�uH�_�h��<����<�u�l��;SSV��w��ǋ�|59��c6��W>/���I����NzI�f����[I�=5V�=��Yŀ4*{�{/�[ƻ4�9ggpC{�c�R��d<]��s�c��w�j��u����i
�Y���.<�k��nO<�fY�Գ^m����Y���xx{ߝ�{�/���c�H@]����M�&���%]:��룉���8�؛��b�潵�����*����`������n��.��n��ر��1s�Ɏm˕9�q������e���>a�1��Cۂ�&�V؝���vH��s���ヶ�}��v�rgܵ6��䬵�K�{q�V*\��N.k�yy�uu&�ӺѬ�¹��e#���]]1���f8|�=��N�#��Q[-�9�l7���ՙӃj����[���MW�;���:����Y�7�S��A�%5���� q�%΅ܰ�gk�u[m��q��]b7%�l'�J��Cz����>��7L�p�k������őj��\�����f��]��׋ �</nqu�݁z�ףQGK��n�:Mv��Xv��δny����Y��iR�kq������'Wt��e��S�5A� �m���<��۲����\��m��/P�C5��K]������ݲ5���r)ӂ�:lE��%ٻ/7��۶́��:S/+ǵbΙ�R�١�]\<�*^Z�M8�ᇆw���I����ݵ��9�^����vz��ܑʔ�"(��8GOg���AԷ�<�����k{�**a-�nW���np��G����f�5ׯO!�'�n֘��-���U���� S���[�E>U�����;�p^,wT��;]��r7��-��n��T�o�\3�.�&�ʡ1�Z�y^y7nz�y�r��wN些m
m��ц�';��
Xr���� �^�w:���h��m��X�N6gX^���<ݒ�x�Щl��n�2��ðn�t��3l88�7;��2�(�ä��2�f�y�<�OA�:�V��q���h6�rBII=����3W��m)�3ӡ3(�,��Ҧ�g��\e��a�!���u���q��d�R`�ݫi�vR�vL��v��V�P���=v��9Ӓ.m�:k��ڱuG�7�{ Woe�/�[�s�;V�:�,����k����ec�ܝ]�7lr�,$1kv}�=�3���k<��\��H��I-��ls�q�:�V��l׎�Lo'1����l��w<��9T�2����<��A�;��zP�5�y�g�K\��^p�>�{%�1UVෙ.kx��q����m��p�{���/le�QZ�\�s�e������r�B�����^��t���*U�t���y�rw�xS���w�w�nj�U��j�Vt���R.Mn�'���خÇ\a�\nuݮ;�z�5�a� <v��GvֻY����4����X	��Ӵ�!��]��r�`ۮ`�;�CƮ�r����n�n�+㳱�\�و���������L�1%���8ͷnK�D�s���ܫ�s��{��ˌ\s���Q�h���ټ�Y]�;c�Ka�vϷ9����k�/&C`�A��A��[cǒ�ˎ:�an��m�1u1�`B�<�a�l��5�97E��z��p�����p��5��ٹ�z�[>�5c+U�!�z0�N���͹ϥl�u��'q�|u�q���R�^rq�/���⥢7�zA4\�]c�puP�v� (��y�^6��c<���Ck�9�/hD�OI���6�=t����8vr�g����cB��C�^����۵�ڬi;'�y��csm���K�����ݻx�m��a�^��s��ی��*�^���ҧ�:\n��rF��y7n����f�5��듑�Umlc�������;s��O��<���b��W�=g�9�;��۫���Ż`[���v'9�Z���4�@=�"FN\�0��Cp��V�^p��x)��yB�T\���e7v�b�xq�j.M��Pu�=��n�@��@Y�خ"싲���ts͐���.}p��f\�k2݋qbv����,��J�vjۮ� n)u��n���+�3ֺ�n ������::�in�x7ez�v\m�'��kR�p�Li��]g���͸�{9La���n�}�[��SpE�W:z^-�k̶�BRg����B�Y}��$�v'uk��m�GY�:�{m��:vkIBA��hYϰs��\���Ky�JsW��a�nsF���#g��{]�ڂa��=�q����tEvy�7���q���n��>zs�h�'��z{�՞��;k$����t��gb÷��q��\ud�vˣňw\�"�v�&em�̰g�/Z�C��+nC�ܩee�mn���8ۍ�.�5�i]=����qX]y��u�w>냙�=Z�X��s�q6S��q{^��K���d�[h�Nǔ}�y�r��<��<���&W��9��[u��9;ǎE�`�g�x�a��ՋC�M����U��y�b{s��cq;�������:g���6xg�4���{WY��n��{=�s�n�݄���=�=�۝Nr�nƃW]��g����2�n	��
�{`��z�`����3v��ޑ�����!�{<���<�kb�H���Gn_`'gr�Sux*v�r�����N��MI:��K���:w��m��Gn�pp�J�;����`�pEŃ�ne���u��>�����T�G�V�qÆ/3��Ϩ���$=�pv
�e�����t�Y�;<�nj'n�{n^ޣ�v+��|;Ŷ^�n��;9��Hv�W�%Y�%7X^�gMω8��Pq�����vl�v�h]������4�hPF��ϝîhw%���y�lղ-k�ۦ�zXmvnm��nn4/8���t�'[�gT'8^˥=k��$ڞ�8�=��O���z6�^�s��#��Ags�Rq��w=r�*y}d��-��wT.�ٛ�����ɍ�[n���v��:գn9x)d	&'�f�۞ݤ���od�7�.��������b�q^�N9NG�]-��[�l/cG\����]A��T�S�e�\N��9���ɷG�͵�:���ˎ��F4����N����F�v"E�M�L�"l��vG���, !����8���8okQ��;z@�σ<@�.5����紮!�α�Ѫ�y��U�']�r���� w��c\�rw���e�<�s�>�������I볺�p��5n.�p7���t)����=���b:��7Lu۷R��\��k��{����/'�[���n��d��yNN�]qn�in����Ǧ�[�,r����؍�Vح�u"0n�-���ͮ����l=U�Y6�h����5�W�8ݸ�S1k�V	�Վ�WB��'g0�����\5u̇;Geݹ	wo%�ܷS�'o]l ܸ�u�ݝ�\��<J�7l����f�:��=�[�#!��݊�۴+�˷cK�cy���tx��d��o<��.�3v��4R�ħ)��vo;�`5�<6]���5B`jӣr��L����Wx�B[�mmՍ�j7\�r�X�j9�p�;˰�L0�;v3κI�b7n\�O<=��]3P<���y�l�n�GS^�s⫺�	On\�ݱS�8q�m�A�2�Hog�9B�E�@��,��o��۪��)l`�ܫ)��e\�7k����]���G�Mխ����3��͛���G7��\�����;>xPq�D�yD�qsػ���k�6�� ���]^s6�ø�N+����K�������>'����сIt{<��q���"�ϧ\I�]��5�/2���ۜ�Ù���s�n���M�׶���غY��q��\k���7I�A���	���wK�WK<�e�`wu[�E�םp[�[\���5!��lu����X͝!b붧�TN��I-f��q�g���P3�8�W�t����0�\�=x��ۺ����1�Smo���K�oG��p�m�Խt!�j��\h������a1=t�Scq�ԗ2�s����z��[���c3x�C�{nM1��KWgm��<�:ٮ���o)9�M�c��sf{������7'oc�v���\\�}T��ˍ��]ɀ�׎0s�;��vB�u�sltl����9M^�,o�ن�v��9,��G���4s�7nV-�N��̼���I.�غv�A�.j�s��G�v���>���b�p�aq�xG(�Zy0�c#�X�yȱ���J&�Q��.ڄ��\%��]���y��9꽫E�̼^�͞��K���+pd�v�)�:�Ff�lMdnb�]���&�NV�W�7�,���1n��(kk���qc:j:ذ*G$�7^.2	q�l^U��e�*ǰ��E��^v�N�n��hN,�s����m�V��=r�q&�.ݤ�T�<��2���ʒgX�SQWkq�]'���@a��H�Svy�=8۴�z�3��w'0>%�y&83��]Pl�(��m�(��.ݗ�V^�F�<�\]q�/=C�N:C�!;�Yxǘ���ۙ�<�y�m9n����zn��z֥^���qh;.䕰�cuٺ��K˰d�A�79�J'#��9����;��9��r���tᇬ]z�u�W[p=-��k�9�J�Y�뢜���q�v�O�7��"�bz����w7O/!������f��FўKb������q\�m�W��T]�ѓ�)7Wg���ۗsg���W�=������mr�>��.Kpk�qscC���㖳�c���qM4�Am�cY�����Vlz���n8���Y�ӝŸ�눢�[."�]Ps.w>{V���s'hum���]˯ou�΍��yx8����yc#���ڼ9nM���)�s��R�[]f��U�q�	tpmּl��vA�(t4�VM��c��m���t�N���We[�e��=M�]��zuLn	�����e�b��wnMـ���xo�;t2�״M��:#p=;���N3ӻ:I��]Og��;s�9w?�r�%��5%eV���j�1T�T�M��yE�T�UX[A����X����ayv(TA�x��H��Eb�J[QX�Q���j�b��EJ���X�V��EF"�Ҷڊr���˵���rmaUm
Z��ڊō�V4�E��\䎲Kj�QKR�m�)F�*d��ԣm"�㵖��o5��J"-��-�R�b����^X�-�1u�mJDB�Q���R.s3*��
Z�r�.�U�Z[kRVQ�Q����[]�]��5��E��Ni�*�������B��mkFט��*)U�T��5Jr�R��*V�VT�Mj5[
���Vd�������ղ���F,S����b�-*-x�[kDm���Zڵ�l����uL�Q�V�XQmU�[��j�\"*��殥�j�m�e�Tk��iΉ$���p��<Lt�Tmf箞7/k��5c���Bs���r�xT�b⴩�۶�"���u=�v	m�ص�5��<n�;�+����v�-�9NwK�[�//�)t��l�[r����3Q�V�]��.��֮�ڽ��K��uJ��4��z��<{$��	��Qŷ8:
Ѹ_���u#ć��:��&�|�=��W:՛��[�.��r�t]�)N+ܻ@�u�Rt�{b8�ңl�^���=c�ZfqnzGl�v�1���ݸ�=�q�ǃZ9ۓtNЬQ��wV��C�h8ð�!���g���Y"�2sR!j�Uۛ=b�Y8�n�v�ڠ�ޏImA����
���Q���A�]�u����t\p�g��_7|=��� �>:�Z7B]�8Bv�N���p���]��ؙ��;n3�Z��X�tq�H���H��q����#ٶ@݊����880+����N�м�듬�]q���C�ض[�y��'��p�z�v1�1����ϋ�����׭��7'��\vy�0]����ۑw0��8���Y��g�ћn�Ј����<���_��g]���Z�c�U�;T6J��x��Da��u���3j �y�5�p<Y~����9۶���X�v��K�I��v�bי�^p�s�r��p)��m�����N$�7K̖(C3���N��&��{n���gp�wn�gM��@=��n��6��tq=75��4��\q��p.�u�֘��t$;3�=3�ݞi��9u����ݛ�6�MɁ�a���F�f� )Ӵ�[z���K�IѶ\��n����n�w)���i#%rc8Tz������=�y�e�fq9�g�9^��v���K���ظN����ѭ=�Ł�k�n{
�X;X��Wku�]����S�<�l(�n����[�:k��r�xܙ�Muu�^�57j�Ef.+Ӧ碕�$�;{���s+^dչ��m[U�q�s�U�̣�h�"[�ַ)v�L\�f��`ơ��A��<�x5c�v�f�y�p�����"�n�yG���<�7�
���r�Mh�[f6�Ll�[T�"�]T���up��mQ*\�� �p2v	��;&���qqL�&�\����[\��svU����6�UL���@�;�}��)2\o� K.�Vm��q�O�3*b�l��Y�5�B޸�~X7Zf����<U!��ZQNW,�ճ��5�P	�n%O^��K��2����U�B���@4"!�I��@��/���5�¾wz����n$<;%�Sl���3����DM[��;@�^�M�o ^\Hx6cI�˪���4O�X�	ݱ O$B�����"N�z��+��OO6-��dT�)@��/ҙ�e�o���Ω&	h$�[CA0�+�:��E��vݵ��Xy�����6�R���{�����s����q�}��]�u^6^��0�}��	;e�YS���(Knj%s�]�D��X��T����3s��s=�� �@�u�)]�z/�u�j����+5QQNkq3P��P�ѳ�t�"�5�gt����;l{��d�����_I� �˪�潊2�.c���G��9l4'�&��ؐvm�*	�'�e-Ks��Ps�"�.���<:�C@+Z��ޛ�e=uPz��uJ�ݶ����[�/��M�p��.���	s^~1��u��%�VM4�\��ۄ����� Zv�U|�9޾��(��S �33?5{[+s�n��^�p�Pp����t3k�V?w�hhL�ɢ!����J�ۺ�=��o%AW/��^��ؔ�f]� έ#�j[$������W�1,����d]e�;��C�0#�n����n�2mk���Ϳ5�&'_}�h %6��e���y� �5����UW7K_��lL�w]~�7�S���R��W�۾ۧf��Y���g5�S����ø�b�����*���wۆ��� �o]״Χ�K�Y���ODHj׵�l�D�<�:����uH8޷R.�{�y9�+.���Y��)�R�G�qL��_LLOn���R��0M��Z�蹺��6���Mu/<��9�NF�S�d6�8^�t�\���㳭��kjq%ё���eHkk��_~�p{����K{�N>�����TL����M[AW:T��v�mR��\H�R�ԉ�6�}>�[5/ތ�J������:��omĀ"�同�ˎ��z�̡?lv�i�C�L��7w<����*��S{���؇�gF�^�^uĀ�����m���'(��ۚ����r2H�Ͻ{�� HYYQ ��ȲP�̺~ү+eubR�3i}*�fe9e���y5�鎼8�K�<��˴��f�'v�X�,]��%WܫI��ߪ�֙�D2�D�Xk�Ă��{wl�
CSa�q |'�Xچ�9|�'�!�U�7q�S =��u^1/l�?��N�n�C���U�ݦ�6z�l�OH=�Hx��G;\�m��4d\nj��a,\�ݚ!�q�
|v��� �ve�x�Y�x��;�Nox����y+��|���&+�HiL���J�����y;Q�?d%���� [ٗT�׫���&�x��6�L���{�m|}پ����d�D�+Ƹ��z�ʊ@���L�	of]W���[��C�x�\ϱR���	����S��*�#s�Sgd61N�l@��~=�|3�<̢"��t�+θNKV�BgTI�캕�����ڈ�Y'F˾Hh˸����Ư^�_8;�쾌�����Áp��F]��ۻ��,<f9�6ҽ̶���_THL9A�`n3)���]ϕ�����⨻;v;<���/��ۺמ�\�f^y��wnS��<��=v�3�F틳���g\\�m�bP�w��xa-T���JՌ���j���H�#���f��9�N7c��:;9�G��x5�^s�m�:��8�ș:������qs�2vu�di�tL�vxz�La����s͋�(���NsW1T�PH�b�n�\�O��fY8�[O&�.qu�3V����SY���(����H�׹L!nv\�;:�QW5K�v;�M/u��<��d}�5<^*r8R�ӊ������E0�m�z���T���HO�쫥���ʴ��\h��b%���Um*@��!H�i�N�&�w[�EKo��P#s�$:$<CÎ�ɢ!�Η�2�w�J���6Wx[ݑ( �Ǻ���w`s߮"�o.�g}\G��\K��>���.��S3kK�U���mj��C��P��<�B/��SK�۳����/o���&:�v�:!������<[\l�v����CI
\@�����c��D��nzR�ʤ���� ��E����jތ�1�kn���� �L5�h�
�*�O�r��]GCm`�ek<w��5<�����9�/��92z��ۻ��K�8�����+W�jWP�������=��hH�|����"�B6b�X)��le�M��@�f�<���)�6�<��}9د��{�>�� ̯L�������w[���rǃ�W1Z��om9EK��"��y@�x�ǹc�4I��F�-��m^�k��UM��}Q� #s"�}�=��B�qDh[k�:}U"�@��YH�S�c����]W5L�nݹ���.g�u!�7�名�˚+q̬�ڙ�xR*� ht>��;u�=��sfr�qzH�ހ�UO�͌E��s]Y��e���;DW-g�y��{��_e�"�V]˕����Wsܲ��o��hL2�x%��^���qDf��gK� ��d�6�.i�q�y�c��G?x:N1�h�w���)��X���^���UqS����[T'���7�����ť����g����x���w�:�ʱ�����q�����-�V4˓��ׯr�	�캩��9Rӑ�i$�N*��%�❕�cD�^JpW��4�Z���el���6c��Y��g�F&�����S�3�Tn�l���y.�%F��ÇA���m>ne�l�yG!�۪~��o���Y��`ګ����cd�x�s�k���r����#��M�[j�������NX���E���"�r�ԀZ���**ng�������@v�]*��k"�B�G��*��5� �w\����g�|�@�wv]*H=����z�Y\�sUM{.xܖ[�gbL�	C?m�z��yg��n���̬33.�[;^|&��12�cwsh�Ω��[ig�$��f	̻�sgkρ��ˌݍ���ۛ��e��7o�uU_9���[��ŵwЇ�n��۹��|�h���qU�i��"º}�^OO^K?`>�;���I$�q��v*�������Y鞈��PѕT�����˔�r}�U�ڵK�T�"@�Dx<2�`�{n��܏g��4�+���n7l͹_g	Y��������!�"%VD�z�����Wϖ�*iƧJ;�f�X�����"w�M>FsN�q#n3�w��M\T� ݺ�/�)���j�z�/)4M9���k!��
v����B.�j\�M����{�f{��[7]J9Ǭ������L�s_H�r�L��S�2��H⫞Pv�L�xoe�'~�5K��<�� Þٔ3�D;�DM"����Fv��p��ЭN�������΀�캡�e�t;�,'.�3��Z�q-I�0�	�ל�vW���}%��.���ZGR�9�d��*^t=��_o�{+)
�\��1�S>�u��k�8����g6��񞺤�[[��wl�M��G�g=��jHh��:��؜�y�f0�sh�3�N�SmۧG;j9�:(hֻM�t��Xݞm�9��S�g'�xɎ��;7���.!��3vٟ$�w7N��1��td�p�GS�.�ڇ@s�s��v���tP�w<u���V7Vc �/k�<��K�5y����-n���n������\�m��>fҷ>>;o���:����ι����~�f�p���k�y@.��i��TM������G�'>⽊*c���b�ʘ�Bbb%��3���@͒q*�u�l���� �~���칠�-��Q��h�
H�7Q��z��0���l`�p���u���T�K� ;[*S�"���ͭ�j\ˉ!��K�u�Kup�)�ٲ�@��˕@��u��)���%�
P�潗
��8��#̢	�n�G�¾݉H�3z�&o�6�C촠A��˪��wnĘ�*H�]Z���8;�Gn�r�]q��ۛ�:.��:csR���K^�uMuo9ͥ���O��!��e�����3)LDǻk&��wněT�{�M��[��*ެ�AZ�3���D<)H�ۅ>�h��\u��o���T�m��{++�I�{������-�*���ߥ
0u����Y������8���ܧ陘��ʠB�݉�	��Ι}�{*��%<r��PΝ<3�;Ft�����
�z�brk��ȒC�^VM!�܉'魉�H�Bjڨ�q^��ܘ����� [ݑ �Ȯl�t��w�[:-X=�J����p�tG��'Q� ��۟'�ּ��~�ɺ������;4�Ko�6�S��d��n�H���5���Ч[�����һqX�^�ִ���ot�P�:�&gDy�C�����_vB��ǲR�em7Ov��n��VU#�ݑZyӐS0�m;���(�P�_AM�^v������Ȑ@��{���&T�O	�E�Wd���iK�)m?���HA��s��:��L㑴�yu�����-�[�]
�W���ls^�~й!�cZ�*�?}t�/�}w��&:�~�.n�6p�^NѮygrA�9�xpM쇆��P<d����Q��m٠���o��dȁO�O{�V7�o��lR߱�N�Ho�钷[�s�F]�![c6��J���Gp��N8Wce����3�y-�_z��xo� �W��h���Ⱥs�w�q�6^�+�A��ۻ�9�'q1�|�*;������r��u�"v��2݅iˇ;t\8�	ۖ
��:�L����V75�j>��;�Cq�u	��3v�m����ȳ0t�r�dZ>�Ĥ�˅�lZ��9{�5}�{��vrH�(��Ԡq�
c��9H�(�:�-�����X����W%ǦtV�i�/{�</�4�/�R���p&0��ǒ��<���z��Em	�N�[E�3�oI��ev�Bn��{�q���^=#ݶ�问�f�(ۭ��6��8c~y,�+�p��΢�u�ͨ	|����d����j۵�s�wa���-��Ԭ��Ge��q�l�RA�񅍝N�H���-_x<.��x�η�:8e���og�T8ѷ:��c4���ڻ4�X{{<�#�w�2�3�d�fNeG)Q�e��6���E���H�&.t���Uߐ�M���c�������=³�^�W6`]���u�S�q�h��;�T��4�Y�o��{���^f93���PV���4������5�n�Q�_a��T�c
�Y,�� ���F�k-�E���D�nq��R�R���h�j����Rƨ�U�������E�hV�VVd�8b��c�șmV��˛0���R�T���m*d�K��͵�5�R�Z�ژj;c53�b�XV4�kTE�4lA�Ae��[mZҰ*��,FQ+-����T����X���`��6�[�6�-+�6��V�b�eAT�-Z�
,�`�-Uu�S �4mK�e�m�*��jJ�[Z�+PbU��T(���	�WYF��+R�QF�D�TjX�mVTh�KbуiP[J�"Y]ffA���Den����4Yh��,رmj5�9��.Z���E-�\�[[E�8�5�)k���E�\�"��e���B��S3j0�!��W�w��ݹ
|v=�F�c�(LlJ[�����s���i����[�d���ν��]1�V�ɏE#���!��Y>�[_��߻�]Z�2��=�Hx�{���Czv�J���Y�4���G�x]n���뮸��x[Tvl�d��.�e�Û�?k˗���^s�ϛ�Ġ�^��ɑ�o-]bS�7�% |�JU��4"<�!�Lݶ�-�.�1���q`/�,���2,̚������>���<�i��a��uE>���̉6�4�;OdL,���{��du�;�ù��g\V]QP6�m� _KԦ Uy� �����˝E��yQ�#ݓ���Vz{�w�D�����ɩ��m�ݞ84�^���T�0��j2:O���Ǘ���I�W��ǉ�L���t�D֊���Kws�n�#������\��y�#"�� �^dϼ�^��v;z��w�V��x��c��p�u��!y�Px+�n.�z5�n�h6eL������~��I*�{/��@�Y���]�1z��eQ
��}���}� ��i���v����3x}�qSWWLv�S�@�7�g�-����y��K���1��dhb<(��G}ؐg\J��x���ّW0�U����Ȕu���=Әή��D;��RE?=`ܻw�cb�U��" ���Ws�M���`�����"B�m���r�O�ݸ��#;�&��h*�z���)����l�H[�� +��Yﵟj}ԛ=(��dz�s=�P��%;X�	��^OQ��CU�C��I����Ot"�?��_�	���}�4�Mv��}\�V�s%	�.�0�Xv5��ip�@fh[�� viI�>we�mv�r��WkWl�8o<I���]Y&��-�7�]"�1�k](��ytvz�{�uZ{���.�s�<=s���n��C>3�\i	�M�u�ݶ:x�����7f{q<ۇ��g���8�l���=Ny�9{���,�g����[n�I:7.���0W�M�0]���9:ݎ��;��Ջm��9�=��땹������Qڿ?O���'��"�ߋ騔�ˉG�ދ3;=n^�yW��);j$'�C���#mTD��mA11S/��I�?sԛ���ٔ/j'�o=�ot���3eoC,_�W� �����@@,�)6<�\.��S���k�b^�Z��� �ʉ@���aT?{`CC�D<�ߵ�3Bf'e?Y�7��3�"f�Q }�]8�NTF�K�,�Ȑ�]\D33��w����^��Gnd�j�i��0�]/DT�I�z==}�$��qQw�4�w��-Q��汎`]�����N��ѣ�� f�bS�س85sRjR�����"gcԦ}�>+��[Li~.�bP�{��7Mc�BxO�D94�٩I��_��T��V��_Ԧ��ɑ��p�k���1~ ���a&s�%4���c��װ~:<��;��R{o1�"�^�B���S��f��탽��:kbr��M�1��Q��1�VvJ��usnKr�Uz��li��n=K!}���u�!���ER:##���j/ա���e0����Jw{v�k�.���?Of-�a�����(��G~�J�j\owYS,�R:%� V�L�/�q#V7&��E��3=��T�m��F6�6�݋ga�z�Ԥ�۪4�m'&�\B2�	�l�m���i�Q�]�x���$v\O�~Q�+�i��^���)�
��d=�,FD'rw��q �|�ɟ6��w�jy� /;&Aݕ
Jz|k�9ۡ4�<?sU��	�<A�=R6:��^�J@�!��KV�������X����ퟫ_���j�M��MCD^)�*�Y�yE���V5�9��1�P�d��G+vSzԶ2U��*���-칐{*$��K�p�i&9j;Z�d����&��L�̈vmB�.�z�܆���?���Cr���:hDy�"�;�`W�Rݵٓ|�7�hod��*% �x��r^qu�R�\ټ�l�ɁL�X�w�iɠ����ڰ#���y���j��^g�����y У��p�*@��) ]}H�y��M��J穙@	}Q �pǱ�d����wr_+��M��>KR�혮l�
�:��@<u�ܲ<=3\�;�K0��W�:��؇�w��n$B;q�X@��ż���5�^ �y���rǶ���(g �r�lI�����n�k!�|޹���d���ri]��V��Z�ncUpm����6��+��]1x���u�3�N�>o׵q�?d�y&�z��
�w�{�\SkP�\��>�#�'whw�q�!��>�
ιS~���k��+�$<	��,� ��\�1�ܻ�&H|䈇u:	�N�u�=�n2F�X��^
Ntv��j<�����q-��;�??������k�v{w��
�w�s�wfL��2�ҟĿdJ Ff=���ڀhQ�x'��l�H�l\���
I��j3v,RofB��,���x�B-�z�P%�ƽ�0����J[^o� H�ܙx����i�O{�����{�2<wfD��%FD'O! i�J�[�[P�׽6�f"]Z��Gnd�W5�?kv���js�c���ɮvzr xrk�F���8ܧ�4��yWf"^^I�;"C��}O#N������5�_�VN��l��� �Y)�B�3�]���o���0�����ښ77S��v�����_���g����Gê����ێ�6S���yʜ���ܬ�{r�%�;��+�K�S:���.��ƛ�wfƆE����d���-ڎx�|[� 89�0�{2'4�^+svc6��.K�iFl^���TĮ��K&9����Φ�t��!�C����)�Q���.�}0i��@,FA�.�$����^Zsһ�N�m7cc6�:�ւ[r���M�L��x*R��nmb�VQ����3��p�&+m����ܣŻz�\����u��������Ǉhg"�/���[�*@k_S�5���+YP�kJ�~�@*�ɔ��^��B!4y�⫙�@Q�O��(�����r$����ۉ�y�D�C�1��P7 �v�C�#�l)�fu:�,�kY�	�_�d�/;"P K���Pt�
 �(!�*�S��=q�u��鶡g�$E��:��]�l�A�Ѫ�Mu��2�Q�	ӻ48���ۺ�| gcܵ4�]��O���s>6�:�+�e|Of�Vk���ǑnY�Cd6�s��B���.�+ٮ�u���s���'��l�V��Ϫ�
 xrV=�zD8ܧ�WtY>9�1�;�8�����2��m�k�T�L�Jhb���'ϖ���=1lwڗ%;�~Y������(�����{����w��2v�T�2nr\2D�]���Lw���qߡ�2!���H�����$�n>@�/���M�"7lE��:�����b��r�'���s<�Ϗ_cܤǐck�&o6vM<�B��2�A+y�z��ژ�v�C���s��y�<��֎c��+m� ��A��&!�g*�A�m�ys�\(�Q�hx�+��Y�ܕ!/^vn��ִ��� ��J@��&I�3Z;Ƿ�+��������ˑ�0[3��,� �����wϝ�nx뎋����\���}�W.q����۔�@u�ܦ [ْ����WlV�qS��T���d�jq��B!���ϳ�D��x�twj�	�+q�_E��7�&A�}{�W,w��`?0�D�Q[����5�X��r$\�M-sQb9ֲ�YV�hS2Fw.��|���Qv����W�·'9A2Û�p�QL��L�]塳:O2T���ɚ}��+�y|��U=N��(��I{�#/����)2��ڤ\�N��P�xx��3�=���ens�l��F�ܱ�fol�sd���r��辙�}kh~� ��s�J����l��k��碅~n��@:�v�����6�TF]���Mhw}�n�v}Llحm�X^Ţ�R���Y���:����r�[Ȉg��}�'�Q�hx��WR���^�dۭ��V�N�;y#��e2+��H=�m�	�8���
Rvܧ�1��"	��+f��5�ۛ�Hsd��<�����=�ƦL㻪MBhv�"*�險�ͼ��&P��=��g��YݕH<\�6�P���� Ɣ��_J�-)5�䪼��[����T�_U!�M��u��k�tJՙ���߫߳�9�D��V��w�ه3����0��ٽ�]9{�n�~���v�r���gE�)�f"�QrqS������.�-����B�����C��⫙�A>�{ꭤ�+�jn�� kd�� :��[1��<?y��{c[Hv����Lp�u��N��SOW$WQǋX�{N�����GKB�O���SC;���v���u>[�d��i�:o+�t^��ʤ3�U�����8��`ۨ�j��ي���2��v�oC��xV�4�+yeA�5���W��s��������Ӎ�И���|�)ELv��f��AMU�Uz,6i�����w-��I���j�)7���6�X����1�f�V<���,� ��v���������⩙����0hj�|�m(���U��x���i7��-}�(AY�b���ڣ[oBˇ˚���u<2féXn�K��<|r����T��Z%��ɣ��,�݁�i"�Hh�Ҧؼ�@xR�7�P��Y���䂉��Y&�G���R��i�V]�žx���<�g�����k\���Dr�J����/��#�bvа�-�tS���h���c`N�W(w�{���<\�&ך�g\�[�D�ö�m
�x���ˈ��	����!�pT��B	ٵM��|Q�i�������k�B�1� ��z:�Z����ǧ{ݝ�D��{ݬ�9}�j���fIy�+4Y�>3�'R�IIw��i:²l��}�c����j:�0���3ۓ�+�_N�i��l�<9g;�36���Nf�t%��pp>(<�����-ބ/����\}T4B���'��Ao.� ���!&v�ш����n�ZY�kx!�'���ɒ��v�Ui�Z�{>�n��=�6��a�53;�QT�I�og�k�s���B!���0�\qG	��S��r�ޯ���ћ<��6�å��+���sg���W|0v����4�GOq�;�n{�!��=�t�$�U^����К��,��D#N�}X���X�|d��;U�d����X���hD��$J�Ц�˝��m2�ω9��,����ޱ�ײ�q��K�e<�zyy��<�0�b�Y��m�kμ�KW�����&�ZmRj��2s*��P�E�ʋh�0S��)T=DHD& g�M�=��Wv�HD��T(	�(K�,�s{�}���5?i͏"�ML�=w7:׼��l��DKhѠ��mm�b[U���Q-UK`�Q�Z�QB��.ڨ�m�cj(�E��-��7�f)��tZ�4G-���L�KUF��"�&����b��FV�k��3^"��e���h-+E�����,Fұ-ij�m���nm�V��ƥ�b�4lJ��[h֋V�9�eu������Q���m�iEN\���E�j7:5*�TJQJ�mj������64�����S!mZ����VȢ1eZ5,�')�)�R�4]hҕ���mkA��ƪU�)EKZr�Ղ�Ȫ��4��� ���6
(��i*U�T�+\�uKh���Ҝ�ܴtU��hU+�kqv����,r\���l�.�m���I[i]hj��:�UJ�,Uڢ��9n���T�����M&
.�.�U���;i��㓵��n2{0�����l�Ͳ�\.'��q���7Q�<)�K�àz2v�[7�:ue�mgkvjx8�&�:�ȼ�I�í	/8�q���S1�Tiu��������r=v�خu�����c��Sv�"7F/n6�S>yݞ�6윲�㫃eq�{`�����H8�N�붳�d��KnÉ�q��Ϗ=lY�4,'<S��۰��H�ݱ�)��y%�`�n/W\�(���N�i���T�<6��,�m�+�=	�ӊ�>^=N�٪N�GNãr��N��][v�9{T��ǜ[�G5��js�·f��m]���c���ך�6�9�T�;<Y#7��s����ݭ��OG�y�^z�j��3�ی�l;�ll��=uC���Ҍk�M�-�G;�\9���L�v�c/r��w< ����<����^ؑ�l�����ɞRwAݐ��,���]�/C�ƺYt�"��[m��TG�9��g�z��4�l�v�zc�rv�J�k7Y�p�m���s�,"EYס�n4/'q���$0`�v��px�m�ۤ2qu�ړ���6���N�]ɳ�u���[�)����F���h8N�s��gcy��I*6�ZԖ5�t�C�4p��b��wr�Y�8{Lb���Ѻ-�:q�^y���F3غr��]Ʈ�ȏ5��)r��p��&{r����-�gw.�:'mv��񶉬m֚wnzqs�����$�Z3̘�m�4R{%��W��v������ptp����OC��;hq�w&l�uM\l���p�sճd�t4�.{P�۔�;�8�[��ͳ�:���nkӞ u��"sۗ<]v:�N��m������G-wl���z��ƻ�yr^	�XYۮ�[���)o&��s���
���͆����3'=2�;\���y㌩����[f�;��G&z/�hڹ�N룗V��.��`ݠ�l�c�{n��.u�k�r�tV*ȕ�U��)H���f�^g:�� �5N:ǡ�9����u�\s�L'7f7\ɼk�籓1���͸`4c�Z@�m����(c�����O9��^j��U����C�<��ܗkp�C�=�bSo,�n�777lgZ�T�n�uѪn��u�^y�z�n힝�8wD��1+��E��{rbƯcs-۶2��}���z�u����>�;�F�ظ�N�٩y
��++X�xb�����y��\Eڳq�f��f��K	��qÛ�����Q��̛�����u��E?�{����vV��kos�ޭ���|�P#��Q]�@An~�е3/���f���:,����ڤ;u�\�̉T�yg�1�Ӹ�(p!���w]/R�u��P��g��bZ�����r�7�vh:��4'��O�_)�qE\=b����t�"��Y ����c�6��/�W��,-W6�I�P��"��٪T��M(�rH�3����PfnҤ�y��Y�.��[�����2J�!�Č����N[n�h��S��a�qu�>�^��Qڅ3�??O��b	4���q���AYݵHGcM����5e���H_k�@]��*J�ƪ��Bq�wq�W���]�����Vtg$3�֩�g��Y\��suّ�4����L�m�CT�r�9�7B�N���M�������ƣ�J�z����{��3 �������_>L}ݳ^����U��f�Լ�y;�C����=@#5��D16��n��3�$��wwm*;m�=�f\'u	�P����Cw.x�}���"�r�sʹ�H
�{i�G��<��}T��w����Х��Ogc����Z3��F[����� ,כi@��w=�Iڡ��#a����8��u�Oլֵ�ivW����u�B\T=g�\e��2�%��f���*hؽn��WkM���+z,�fL9L]�Tf_�����ϵVS�6�0h������R�&��U��eM6v]fQ�F�6�[�r�H�qm�x����퉤5ṖM
�K��A.��X@BH�[zo�Y��ݓ��6g���sƙ�Y��t@�?{ך�{}��u��R@�!՞[e|r�?w}g^��7yy��N6dݼ������K�W^�|�.o��Hzo�,�'�k�P46�Ɯԥ��Qwj�M�9c��gf����'��]}�Z�ץJ�b��鷔	FK`'L�'fw�'a� ;/2�T���	�޵��t��m�إ [}�T�{��ߛ����p�N�c��vG��F��^pj΀��U<s��޽��l��P�����?c��)�is��<� ��{���ݪF�#��	���zn�y@���r��h�èL��T�ٚ�A5*}X<�#y�������J�ݪ@�~�)��:#q�el�M`��%�Zکݥ�����kʐճx���/�����吁u����l�qhY�V���w��v���lL��y'�+�ݪ�\�6�m��n�tC썕f�5�f�-�v�)%q�-��b���q\�o<�abz�X�Ff�_B��v�qS;�|:!d��YE����wG�^����� >�z%=�rq�x��hx%xwﺨl��p~�ڙ��j�����@vn�!�ɷ�j���������(�yn�/7��S���.3�q�Y�\a�nۃ�Zs+yLc�
;�1�8���?_����1�1���ݥ@$�&�U�\.:�MU5I���_� �w��%ز�D4��ˊFm���\߸E_��x��@�}۳H�#)� H�K�՘8w��#G00K)i)6?/�S@��m<�uNf�M�cftL��u�ǕB��Z�!�}hĊ����b����c"��fh�Z��7fA!�����m<� ��!�+;����+�˪�cM�d:�!���T��1�$_cиf�.��lX{9U�G��
�{�֩�ރ�_Dŋ%y��T�����^>��/�^ۻ$�ڵ�}�/7��c�[Z��q��ٲ�AK�{Y6���)�l{�R��i���//{��Gɚ�����.d�i7	�Q�9q˦�ex���eg[�퇕'l<-�r�n�vs���ѐqi�<Y�dz�v%��ݷ8]�a������z-�\l9�T�q��:�L���Y��4��l�۶K��c��m��_&�E9�7�:Q�c2�^C�$����z��a]�^:�"v	��qӭ9�uK1��ȇb;������(*VzLѹ]N<�����@��\�rt¯hG��(D��o��Х�M��rӟҭ����m<� ��N��%��_zg �mT�ѹW>pԦK�Zw�<>����0����@-h�y@*�z�ކ­��]�{<ݛ�)ͩͪ�<:|�O+��ǡJD��K�<=�����+#)���)��*�@�B��"�>�ŭƞ�jt���S�72(��7�v��o$�ˁ[<k�D�4\DA:!ݢ!�ݗ�L+���ت�5��4�;^�̀�vn�{�R���������1�!�Xy�#�m�ͷb����7��'V�rj�[�d��gO��C��i�-j�u �w�S� ;�v�͛�f+z�:t�\�x6[��gq�tr��h����	���G]�Nl�����j��n����x��?!��l�q�'O��ͬ-�����0����Oy;�w6x=�~LtydǺ��=��r�%;�}æ��y$��Tkv7��/�'��/��ڠ�5Q�>n ��lA�ɡ����x�1��@u��P��#��S�/&�so&Rn�Jd�n��ޓ�4�݁��)���vڙ9JTf�.ɚ�/��ov�x{���e�' ���C����7��"In$@�ƭu���L�����NZ	~�%��ٻT�N�����	�nr��"w�5��Bn�����u��nQ;k��t��Pq�v�m������� tC�DC�F\����4�4e<�zgtO]旸�zw{v���Ε��Bd�i��oʢ&bs\d��LWRC�;�&z�;j�挧R-�j�����WP/j�&Ԧ�P9i�}��}�^aO!�#�㓽r~���Fӵ�m!�!�g����,H�t.d3��v;ꮰ��q����K2��֪�~}�;ņ���D}�S��B����h�u=sC��ǆ b*�S�3���i��5�@����@+h�yA�V��C��'"�<��ͺ�]oIۡ�Ρ����)���D#;��ut����mq�l��x����O�ܮ�#�)�r��*Lg�	�Z9�M��{(�L���X[u���T+Ӽbm�����������@1���MJ���y@�oE�1����Vq:�GUU 8�����2Q�����u�3���PQ�����SW�F����dx���f�vv���z�Kt�!����q� +�z�ǀ����mX��n�*&/y\�+�Դ�6�)�Njy��7W��S�>��U<��z(�-���8ϹJ[%q*M���^#H)M��u���l{���0�ۢ�~c�f以r�i���F!��s����H�=��󜯗�� �)��������w�Zxb!⨩��
���
�qv㨘j<
!�P Fg=O��}�4d,���(���ۯB�P�(!� N	��Ns��q�c������|�؆�e��"�9�uι���~�o�a�x`h!}��i@.�z��@��v��R.^���2 �_�����2)�"a�i"3����q6i\3��ku���2(�u��R@�m���}C)�j�fbjl�I��(���U�K�}��۹"�[J�7����y�R��ݪ'�ה�\�4�c�������/r��O��A���@������vjJ2w�2���g�妁�)NZsRs�<25�Ka�:����WHvvң�	Fr/����X���0�s�<�N�XA��^���mk)�Ιb�/:�d4�N�Kr�n]U�"�vز	x�f���*����W�=���ߛ����ߣ�7��vl�톷��CßO�4�:5M7�[��k�K.����I�3��.N�����@=�x�=h�>g� ��CSv��v�s�!�c�F��:�1T��m�Mţ77v�Q�w�g�����	9�g��@�6w�c�iL�3;]˷���,Ӝm</=3�:�����^٥9�EP���}�ghE+Tusg$p�j+����up�gu�r�R���@���㣾��=�9M�0m�~��_�IjS%�-<�D�b�L �۵@FF�h]��Ҍ{z�B]۴���i�}u){آ|'�,���W}W��� ���Ttc�>��90����}�Ʃ�T�������TwT�PF�
Px�AY{�O]�)A��ݪё��&6˼;�8DCό�|]������Bqт�[�SB�Ʒ|�ڱx���@tۍ��CEV�F�A��iF�t���T�,��%o=O�N�=�҇�3��!Ķ�0�o�iOmV`�SM��$;�2t��G[q�Du��W�����0��C��m���	29�@�*�%i�L?wN�,��$ۚA�p��ӫ�n�U�;�����.�^�*��sFI���_���]z�Gg��jjs��z}�� �~bnj�{I&1���쭕�Úǵt�α��/�����I/$���#�	*���ZN������Am4���;����B���$G��z���w�u��ʝ���A뎋$<����9j����&xf����Κfy�hEL��H:��R ��(�u���/�<�7)�,�},R�Ci-�m��k�&&g�ݷe���++���QD��ǩM�m��P�=Y�Գc�\�"~S#a�(�4�!���U�r�ui�s͛�2@u��Y;ny�t�~����ź�!��h�J�#	@+�z'�=�۵^*_o`��͈̈́�=/F�x�ǩI����&!���槓���Ǻ7o�Ein�R<V�Q(.�ݪl�I�&3N��1��Ǻ�WL��(%�wuʪ��{�fSnE�u�]n���𻯲��)IgE����"&���Q�ɖ=�t��*c����CBK4��8�<��x?]BG9S�[�WOk#�3S��/���\�Hm��i�^P�|}�g����\�!f��S�pp}	�������6
dz����j�N���������.�纷��,(�o���z� ���@�c��GS�b|�����0��l�&�FOF�n�HRHx�x�E�#N�
4o<NC�zI��n��:m�y���{I39�ӦS���T/.�k~]	�y��]�
��a�Ļ��i�����B��	��:u�A�����S�u ��l��L\�1�W6�˔1�](Ѥҗ8R(.wt�J�׉��|/q��sn.�����%ia�U��Ȯ�| 9</����U`��=�{Z�PAIKq!�b]���%��K�}^#�� s)��3Sbը>�i��	@�s#��g���GS�O}�j}�K�xM��-+C�ѠcZ�ԋs�*���ٮPX�y�6�l�n����}�e��5LK�α�r��#0K�;��3�s\���H��6�zmy65�)익gu粳,k!�:�W��J����Ǟ�}F�x��ۗ��Yh$J�Sn<��[�Ks���KC��)�7�Dn0�}vGz̆-.�/x��)Z+V39�����+L��U!�����Lr(�s(�ֹUN/u(�����y���ȳjs���y�o�k��.x��J�e�_g	w���޿��V�Z�嶗4�jRT-meh���AE8�
�ƍZ�PYT��E�*���Ķ��m+iV�:�F#Z�DRґK�
��Dmm)��r��e�Z�[khҴaR-�b��J�m�F"Ɣj��J��akm�JQ��JZ�5����j6��gu�kVT)j�l�Zж֣l��b![-�DC5���UVR�R�r´J����*Z�Z�H��lkk�[Q��-h�������TRT*���D�^XQ��Ū�UV<�,r�Ns^]��kZZ�����Q���UcV�[lm��,P�+E��)mA�"b͋0�
[9��U��ʭ��ڊ�J"�VEb*Ȣ2*"��iX�4BԠ���TQ�֔�U8���JT�TR�5,UkX�(���)���D\؂�(���J�����J9*�'-UU�D�g$QGYU�d��k32aڎ�	$���w���?����>��j�.i�Νjw�xpe���ɖ�	k�zR[�d�#��j�_LQp�gMqs\&��iX���������'<gK�>F[ �Q/	�m~֟3��h�b�-�.�[����g�^��isj��A���Z�ɮ���׵����: yӛxCD3�D9��Nˀu�mQ���%#�"G�ً�k܃g9�S3�$��vv�Rj�;C�D39M�JV�E�~����f�Ҥ��j&bp��ve�Ȭ.�D-�)���;��~�T7e�@��v�OS����j7e�V�mW�x���Q�u+f@pؔ7Wl�}-bw�I��U;u>��%B�n��w���4��xk��<9�tJ��-d��b�or��B7��eH{I�y̭�v�6�q���) �zv��9/b<K�����|�o)RƪL��'�g�O��"� g͙)�U&c�Vbn�ܥI��JZݓ��-L�7���7��P��1��7O:�h���<�;���KA�]r�ָu�6b�(�DD���:d�<3C��"�ji:^�G�V�cH�ٕ�DN�ɻ� ����kd�h�v�"!��;.�1ض�F����B��(S�+[�]xz��+�~��Ŗ�+~X�'B+��b�vK�O��eZ׎2�tgLQ(��ғ�jy�e��<���̪m���2|�s��� J��JAݛ��j��z���ۻ�k��O�ch�	i�
��������y��Y��f�]�y��D"����{{7j�=��ssd�.���O����F�ݚ�l�n�?�.�杢w~^�sF{�n&5�b^ @�2>�|S^hsÙ�X���?gok{'�K'��l��`���@���&�U�Sۣy�s�]��n.:-�=R;���ێ��q@��'�][�8�[<�:�Km��r��ۉbk�Z(��m�Y�
��z��M�ɺ�ֹ1ڋ=M�gs�ܛ�y툇8'�����0���rs��sm��Ws�i�1U���s)�p�̍�W6�4��q��.wG 8��o�2�;���ڱ�1���5�sgM�͞��s��;�jyu�чlN.��kz�ֻ*���:���߼.�z��ã潊'���l�����گZε�m��g5��>���@@�Be]��ؙN?4��׷3o�xB@��-�{�7j��{7>���X�����"!���i�t{�IP-2��e��cW4�Q��n2�[ٻJ��[����P��g�T�7Ro&�o8���vh��on��%e�7��¸k�N'��%A���C�(؎�T��z'��Y�3wn�0�P
��P��v����;��!T����d3����4G�xC�����J�]��qrmǋ(½;b9��v��6������?L49����Ja�98���4}1G�Y�Wj�2�<PW7S)��ݥ\�I�:���9+_"����W}V�XfS3E��^f�W��g���'[^f�2V4�ͮ�~�~���=;�`Pn�]�Fzk�D�n�NkP�jޠ������i��(��X�26�i���^��i�[�!}�}�^��(���|/5�l�(|���4L�gۛ���J��^�6����H λkm�5ٷP�}-HV�m��=�W1^d�m6Kmd��ۈ���Zf��0������1D�@���S5�����}��v͠J�-�xK��R�w��W�3�v7]g���]�[����Z�2b�H��/��^�]��`�ī+q��ĴE"dr�"RR4�)��œ��<6;n7������a����:�>�hr�����x�BFl�� �~���(8~U=����n�W$ܘ�I�r�L�KH�N��:��3���ܮL��3�gK�"+[�]�47,�f�}�\L�d�C��Rmȣґ��r����\n�ȹ���=��9S�{�������uGq������u��E�Da��s�6ws��i˗��]701m�Q/���mҏ���^�ٚ��3�'�\�\�)�����!���h�٭��g>�s����R ��-���ݞ��^��v�@�=��V�ΞL��D<��;.�{�T�Z���=1]8#IH#5��:.�ݪG���o����y���(q��K�r��Q��рcsc���gh�V�8+��M����}��K��CX��q��@-�ݪ��|�[���MD�ϰ�S��UP�ӑ�9.�}�H��ӯOR��m> ��ک�\Z�Y��og>��GKh�<U"��ZP��v���5�r�Ev���.ۮ_�[ٻJ���fu��ǈu)�"�j���±]<₝��΄�ݻ���R�e�	�Ig��0z*�Чפ��J�w��y�U�n���w��\;8�u� 4y�"m�r�Uon�?k,��ގ,>������&��S���Zpt����I����&�F'��p��)��i@��T�+�:�_����ιuݛ�L��y����Á��]�:ݍ���uƲ���i�ڿ�������x��-�%86�����C�:·��!�%ЁWomW��7*!�M�)b�;��b}�cީ��J��k�"��f�x/�(� i�e|�v�8�x<����4CI����/B�.r�],�Ox�9��=ݝ��<��(��̴N�4�)C��tu8̋����Bo!߷)P̗�PZݔtoC9C�Z&E��]�H=�T3;��x���?6<��x�l�I����l�ʌWM!9u@
�b�@�"��%<��ۍ���pח�]��jǭ���PM���c������)}��gR{��'�v����)��M�φ���꼏6�1�<t3�ʭU���r~����z�����9�S\YN��ĳ��8�U�y9ݍێ�T[C���vp��Y6�,�:Ur��%[U�m�۬w=av��Q�N�匼�h,�-v[{�S��ut��vR�����ׅ0����r����[���k�1��瑸�����:�v<l{`��n�5�0Q�8�y��U<�x���ĝʈ�k�t� {�<q;�N����u��:���Aj"9:՝�3�K��x2�qmKЖ��l���x�r�b��s��>���1������{5J�gK�)@�կ�ˋ�8fD�U��""3*�x��{�%���8��x�����Dų�d�mB%�u*d� QݓCK�FOZz�+�eD3�Bw!��n0��_d����L<�\��߫۳HyE�>���?�m46�y��^�NH�w&~��{% ���<���ڹV��P�L��=���Q3ݖ���b�1;��5�J
�wf��:w܌VU�:�)�*��ݚ@���w��}�l��r�D��Z��s�<(�w�>m����k[M��*���q����o��3��q����v�*��P ��ڡmT�
�o<�1$�<�ި}u�D�P�F��P�]z�sD [G��ˇ㿌?@W���H��lu��0V�n����{�/�)s-��A4�g���2�l� �h;ȦL���]4�g���I{���= ��ǐG�f�+��:�rsG���$,�&x��<CɆ���{f��7���e���xG�/1ԯvn��nTC'f��C�3���o7�͝����';vRP$ ��v�_LQ�/r����ƻ�W����0��|8p�i��S��_�s1�J�;���Ǯ��M�������ٯ�d�Ɏs$ ſ��Ç�sQX�1
ud�6j:6����¡�w_�5Ǿp��p?-�������C(r�� ���"�wj�����C���}�iشYR�ǻ{v��؇g�<@��V�E�te�1�茞֮��#3wf� ���|����{;q�b1��>���t:u ���4�ޚ��e�2�^F�mC� -����wF�8̳i�8��������i��}�mY�x��O�A�S.C��L�8<.����<�_�������/��T옢P!ndS��%�R�U>�|��y�l�K�ʪ ͗�P�V�Z�X����D�Oӗqk�{֙�41]����9�eD=��G63�U��.z���1d��\�r�ՙ�Zj�sC�c�p�$�	L�|�P[�����iL�����x׭�mZ�V��������������B��)���*����%<���=^��&,���*u��Lc�1;�tu9���f��J�;k�А%�1d�@V�\����Z�����T_ޥg9i8C�P��N}?{�e)�г&�9�ѕ��\j��b�B
��*:.�iD��̍�'q^�V��]�ș��D���u��su4t�F֛������Ǯ�������vS3���9�mq�hם8.�7`ɣ(i��5h}�k��	�Q��[- D�}Q?/%�����d��0C�'L�<Cɼӭ(�;j���V�NJw�i��˗G�o�j�c&����\��>�ހ�����[;���k�L�hF���giSHu��[g�u���o��X�I!����{ǟ "���	��گ#U-{�۞���ZwPx7n|�/]��
<C�4DJ9�V.fYάu�<f6[J ��ڤ��ג�������:p�\������⨉m�q/;v��%u�D�ͭ0�u��Fcm7�u��W�t�6�-8�P�@f���\�;qy32��S�=���H.h�WU�K�dB���i�U���'P��I�5J��e����S�%��+���R�A���^@і�G��J����=���׋���:Ry�:�퐝TA<��2��s��Sh՜��{��B����	�ys.#�@.�Ym	Ǫ#�rr�)K;��s�7�)BƷZ���'��r^ȕ�V�I��iT��z`=��m��V&cd�eQ����Ld�;�4]Pr����^��vK!�G]�f�z�Ѯ������|���s����wA�yV	��	o$<��/{� �_H4�Y�H��,�!�t%7���=���8o���G��`�v��re^���Y���m�h@��w���/9��F�O3����S�ñ2Ȃoy�pݫ�s��ԝ��2�f�Q����։���N�a�Gsy�o.Ֆ�s�)��t����7��߷��]��aOK���w4�"΂���4�b�#�B`�.e���Y0�,�Y^V$���(���T���F�嫕����������Q�,�,~<cdPOq�f���5��V�7��(�)�wiE�xw�8��^�ov�=��?���U=%�7�,�7��!��r���ɤ�3N߱���oE �p�焎KS�:�Y�`�:�Ӷ�9FɽfK'C^YK��{���{�@�K|���#��K~��[$�r�wN�%cU�,�]Udl�C����)����l0���_�7ޏ��L�gMZ|zǌ�8^a�c��Y�i�Laql���^G_�,�2�ﳲ��/�ڴ�	�Ӽ�����ٗ�T��4��p���F��M���M��4#U�*�	&�Е<���,�+���A�[`!�U�r�KM��*(
U��jE`���U+R(��e�
�	���
�"Ъ��s�:���skER(*�
��Ց�DEC�R�`�&aS[�J���+,b+s���U�B�(�()]��""�e�rŋ"��F ���
�e��^%x��UZ��-ZX#b�x�`�dR3����<��J�"�Z1
�SZ
�� �5�U�J�"�[Pբ�l)��jAdV������QK�H�%(���U���x��PPD������P+Ģa�eYn��Y7��k8�b[EU`�,**�l��UR����E�'0r� )QVJ��Eb6ب�"�h��*"�L�+U2U�֠�(��+w�ȝZ��o7d�����8��r/bR���8C�'��{;v��v+��c�h�s��:�Sێp1˒mf�놻�]��<����Z��8`m�>��q{v��fP����S������=��{\���{m���5q!��0�n62v�LXy;{D���t���ˀ�x���c���l ��n݋���:�����Z�v�
�t��/�m����>Ę3�y��9K�E�n=u�:i�z� ��c����p�۩ס����[�S|Κѻ6#kuw�q|�u���ց$�9˭��ܖ��i���<��a���GWnN�;�7��s�ƞ�g�;n��*puض�N
b���cb���K�&�zҚ񱝝�����u��Vk��q��͵�gu������Wm�Ruzr����WIj��Εd|���٥�9�ƴ������t����} �y��|�ۭ�l:#v"���0���c��c.�7��Â�=��^L�<<3NSsJq������N��mmË���Q��.���n����c��*�:ܓ���v�D��b��Ss�g�;^�kR�]c
��=�{vn�����t玚s��������=���[�D��ea�:�3�����˞sV�R;��=��,�vZ��cI)��`�&��U���k��E�����L]h��h�vGn^�{^t]�p�O=�<WA�'Z���n^;�R������@kp�c��T�![�C�vUݮ�Ӟ8�!'e5���ۨ�佃��G��;��
�v���öv�0S�K�u��Cn
�y�Ê��q���;�4�r�W��-�9��v�O��\Y� ]�9Pp��m:W���;����kq�^�v��L���n�\�Jr�q=W< 'nR8\u����s���d�̓5��Ul.(�2�ĸ��8�6y�\�>6����t��cF����� �n͕�,�d}�or�:[kK�P��<�ɩ�a�GC�苉�궘1Wm�P�e��H���k����g^Զm�}��P�8�x���a#�����X�i��8�8�U�9�����|p�F�\aN`�%�� R��n��%���lC(�ny�xG���Q1�;��AB�4w+2�1ES���-p]���"���'-m+j��/7m˹��9IB�4����1]����C�|u����{\��8��F�[���U�֛?ϟ;��qD��,���k��X��eB��Gk!{X���k�����<N]K��8�O߿?s��N��x���Ɲ��nvU!4e���9�T�:)W4v�o{*�
���B����֯}3��ӗX�*h^�Md3�:<7�)P.h�u'L��1y��vmS�k^�O�Æ�Cu��}�L�an�Ǣ�����ܜ���mB;�r��3�ت&c�Is�&ؓ�1;��iz����]�#w�+�xh�y��ꊨ�����VQ��J��`!�;���:��{ke5sT�5J���^�cGb��bc����$��s�8��a�D��i�1��=�^ۊ��MmZ�,6�n�ً��qTn��	�!��7�Wd�Q���e���־��]��a�f�w�9�)Џ��F�"�F�GE}Q���v�%`�N�EM8o춶�@��0�֫���6��O1�r=���J?.�i!�l�U�l�ݛ)C9������犾��5�i�(���}9md�ez��$�<�w阌q=�l���4�����J(�P E���Z��l�r ��e<�A�ʟF��&!D��튎����bDcπF5�<����m���V_D�:�S6���|�bNP���<s39۹wј;˶��=�R�0�ٷ4x�,+��g�����m����Kq�$W�U��j�<m�y�=41D�m*�Ӝ�Nr�"��=�U ����@�ݛsHYw.�-���1) #��y�+��!��*�횪�}�wZ��G猙 �}�� �������b�t��4��#�ݿ��	&�7n�:k��� ��<�������CDq��ԦXJ!�Nʑ�N�T�j���3��Hv��Ʃ�!�0�׋ѝ��=���59%�3ڑ,|�D��������[0�3317\҆��zɸ=u��h:�Q��?��m��X�f�| |�]Ų  7v�n��[��fFF���w(��v�{6U�ˆ��m����f�� �6�|�ͫ�q�F^������n �ud�� �LD?W�+6��=۷�JK��nke
�����㱻<x]����T����[]�7M,P��0�ߛm$�����U��;�M� Ǳ��6���%=/
�}w��;v�n��ű-5)��:��F�S3������E���2{�M\� {C$�5�'|��G^�a���͢Hn$m	;���u\��Ǳ�$Y���f2��{�o�̙�z,�I�1Ǳ�	��	_��R��3��	��״L�]����� 1{���,�_��k���L����53�:���O�B��M�W�^��>r=��Ԗ?]��" <��_4���c:�H�s�!<���;q���|�}�ߗ�^�3W?|�3q����iKr&���?]C  /��s~Fl��1׽���J��N�p	I��.���(�F���9:6��6-`��3�[��v$Q� wU����L�Ҝ���;8�CR���WD�[��%���n�\Y338n:���D��j�6�v4_������4� &x�:�F�aS���i��L��/��S>�>���u�9�|u���L���w�e)�pD�-������i�:BȔ�	����C���ɐ;ˋs3=�;ֽ�4kW�����	�Ʀfg��Ҟ�jiCq#i$�t�>����\�� %Θ�ٯ,� �>��q��D�;� �Z��}W�+�8P�jSt����jd��[�ŏI��EeY���S2Jj�{�v�du��{+��y�Rh�/~^�m�Q���.ե��5�ȵ��㗧l���qY�b�y�$rT̙������[���Cć<W�j6��5��a���o86� �,=\�1a����n�&I�ȗ-�1��ӭs�X��x�q�d-�m�uC�y)���&^�㴼�A����'�������.�6τ�r퍁��������v�{WA[u�����3�mp�)��ɝ[;g�"���v�b���p��^ݸ�]�yt�r-��͎�M��v.��s6�u�#�[��n]Gu�ޜƉ��6��כfݧt�"Aob����՟��߿�}��	�ۿ���_0����.��ɾ컰U1�>w�@Y�� gj˸A��]��y�r��9��s��O���!RTʔ�x���j����ix�S�2�;���a�Ο{�׽��2J�IP��O����yĜ��$�W��u=�N�j��R(ל�"V)s��Ե���<4^7�nw��%B�����!ĕ
�P�=���v��L�d�0�&FI���
_�������%`X�^d\�*��3y}�\yQG�a�jn����my����yÉ�>�����;=񟙐���g���Fx�T*2�����^!�!�g)8����}�R/��icT12�Q�h�P�+�����C��N$ɽ;���Zs�w6۝�$��f}�<g��L�9&C�'�~���8��}���κ����{��CǦ���>���T*x!��>���v�l�3!�T*J�m��GP�I�,��O���T�e}�����Bg#.�{�v[Jky�n9��9�����8��t�����_�p�ۜw9��:a��3������$چI�C0����;I_d�2d�7�����I�*J�7�~������ο�I�+�]s����\Rd6������T+���(�9˹��w��%O���'��Hd�
�<�~߷?M��l}Q�8���"�{J�
c;G �d2YDO5�J����:�w�������C(e��]{D�1�� I��=��<��3�8����a2�����{�x��!�T*M5?���*�JY'�I��!祴�~�����p�^q>�j{�"!���"���L����U�>$���2%Ov��G)��I��a�'s�ݽ�����v�y��v�OP�d�d32}����C�y���2'����q���v{{My�^7�nw��C>}qr����k�n%"�	0��Lyu}���g�3�d�2d�1����gq;$�T�
���=�����~�Ի���^�&�I�/���a*>�<�I���l��^[��s�v�i��Ns~���8�gq���g�sޏ#<C���ߙ�Z;k�H��N$��em0�x�39���}�GvuC$�T��3���{�<O�2n��~����zk��J�M�(�ɕ��=��kc����Z����7�)�M����������uvm���J�	�y�������39&C�'�~����t��&C$�W~��r��I�bN$�W���b����K�Оy���x�d34fC!�'�7��qӤ3�߮�m��ns�퇃��������$چH����~����y�^u_Y�L�IS&I�O�Ͻ��N!RVv䙘s�����x��I���I�m>c��|���R�\ba�����ʍ�<ܼ�:�Hv�D2~���Gq
��Y�2���{��g�q&C!�!�>o���Ͽ�u����T��!	��^b����^{}�K������[��A��O{p��
hp[��L�9b�Sü��\6�n�}����}_� ������|��X�!�cS���z8���%B��f~�sޡ�P/8���=�(��b")H�b�9���t�﮲��
azĘ^a)v^qs�~ts�N�ړ!�0�g߿��P��!�Ʉ2�O���ު3�k���������T8�̆C&O�����N!Xvy����Ss������!��|��<�<��q%B��P�=���z���&^�s��o�O5�=�'I��&M9�~��ĜB��T��������x��)2%B���w�U#�}�ީ���|b��~��]u=8�xnqܻ]������p<��c�n�T;��v]W:�\߿����r7(-�s�<C������G�:C$�Va��������*�f}9,%G��$�}�s�F��	8�)����Ύ$�%{fI���������L���ӯ0�qn��s�ĕ<0���\J��=hqyę�ﶫ��κ9{����z9�I�%B�0�gO?u�p��!�ɐ�fd�����!�<�q'<�q'��������Ղi�T�N���ϻ�w+��9�λC�9���~�<|C�6��mC0��~���3ę
��L�'~�:��Ϻ��|��~8���d���34s����z��xr�!RT.,>���z�x�0�g�?���n9����s�t�i���7_�8�y��-�*�S�p���$Ǥ�9W�\�=�CD�d4L�a�}�����8��N8���/��%@��)[xܞ����!��������>�Gw�A���"	�W	8y����X��˱��c�d�zA�/������j��e�~������ݯ��$���+�fI���s��<O�2`�~�����9�^s��$�<0�u�����&f�!�I�ݿ{*�g�y���B�|��Z/0������<C!�T+0�����$�Vx̆C	��o�z8�bt�a�;~��o��^1%*ZR��CNdlR�#@�Q��n_;Vrz�����.�n��כ��ޞ���p�ח�������3�^�Ρ�'��IP�=����g�x�8fI�&I�}�ܥ�
��^sٛ�}��Y�/|{9��y�<C�Rd.�����������2����3���k��<C��C�J�z��$yĜ�sȻ�ƍ}��y���G��������?}��U�y�IP�6�����q'}Pqy�<�󏻹^I��>���.
E쟏=9��6�]w:;IP�;��םVGę�9&B���߽��e'Hd�I��<�I����]�
�g�4�z����ȆC$�V�}��U�T+<fC!�'����qӤ3N�o%����
"�J�+IϹ�,m�(��j&�3����W�x�8fI�&I��Ͻ��N'bd���2��*m�׿/�����{���^q'v����a+,�q'�Gj{L3�v�����Hx�D2}���'b!�����<�N^?�*�X��_|ܾ����>�Ҭ��b\%��9�=��TyZI�-�I�O��{�ĝ�C$�fI����d�P�R/8�Q�_��&i٧�9cc����<��[��ޓ��x� �);�.���>6q��͈����cM�]H�j��E�+�V�N�π�U?ǒ�����<��yuz�c���͑i|f��Y�e���Z֧��i�ֳ{sz�<���o[m�^۷;�*t�����2ܦEI���x�.ڝyGm�={nmh��BӮ@� ,�cc�W� �gn� t[]\H�k�7>k-��x��9�Ѻc�+v�M�^���ـu��ǘ��8�ҽ��!����j|u!Y�F�����y扠�gP��݁wg9��ut���u]���8a�wV��޸��[��W������]��MW������:��3�>$����2{���s���6)2�2����C�8�)8���-پ���a�X���,��eļg�2�3!�ɓ����C���v{N�Tە�ۛ���!������I������gaX~�����%B���2L���ގ$�v�&B�������z��y�L�ԙKT�ҟ��o��*��q/��'s���߳��v��u��<�����d�B��fC$�W�����v�Cș$��9�U�l�V}�+�7yĸ��t3�2M5?^}�FI�����&s3��sޡ�x'd�Ǿ����׆!╋�$Ǖl}��-|���n�����d*J�������t��&C9�C>���z�hd�
��Y������Yzם��v�����q�fC!�����z2N!Xw)ߏr�r�u��w�0�9�����;C$�T��a���.Y�����#���$��	�/�fI��L�3I��������x�����L������Yd3���������~�v���y�'r/8�Z9�z�y��kL�+q�!!nJ�����ߟ��q��כ�����<���d����̆IP����Fx��d22�~���Ĭ�!Ĝ��}گ�^٩����'s�%s2L�g�߹�P�<�ę1�������9�Βx�)�/�k�s֋��/8����f����sד��{��n��Zud3uX^��Z��`	�n��Kd9tK����m�7:6;����	�<z_<��xjk���p�+�������S?���zD��������!��C!�D2�O���~�!�<��ffd2���x�K����I�,�\ʹ�nV�nns���<r���A�|C�*&C0���~�>3ę
��S�"�S�eb�UY�\�^�`�^s·��|������&Ck��}����*���Ϋ���x]�����;W�N��)��Js�e�9���q�G�Iɣ2������<C�`L�IP�7��}����<�a�!�mO�?�������K�Q���I��s�_�GO��ȜI���x�m�]��s���<0��_u����!RT*J�]�ތ��M��;F�3;���%$��Ĝ�'��2x!��*�'��~��C�x�ffd2L�^{ѐ�:C0�o�������?7̠;�E�sH������u��/U��.�����)�'��ߛ�߰0�S�ϻC�C>�󟺇hd�j&�3����g��$�T�4L�&�s��̓�ؙ&e=����>󴞡^��>������2X{�_~�!���q�������79���'��^OJqz��yq'=��] 7�_d;�v�����3�8��RT+����C�G!�T*Lj}y��FI�:��T*J����}�x�s���	ę1�|b� !<D3JE���/���c�>$�Òd4ԙ=����N�ڑĜ^a&{��L��K�K5���FE:��%��u���uJ�ۗ�Ys����z�\^�3u<}��Z����vn��.V�m�C�ro�����{��Bttk��f�}EHp�w��z�a!(3�z�K�{uqn�4����Q��u��&\�6��I��g����Sжg-����΢^*��;����l�hc�+`7P�bwfY)�8��5���8S���W
M�#���%ɛ��h+��r>㓯�@�K�v?������p^[e���?%��� bsjyz�-���;��
y���e>��}�a� ��ԍ�b�*e>+Ιzt-���ࠛa.b�<���D�(&�����pYԟ-��ADv9�Y��0�d�ݼ����a�CS;����s�������e�>��vq�-q�KYn��ӝ�rc���_n�e���B��ؖ�:&^�ۓp�VÛ��Ԃ��{��_,�H�W��v7\F1������"k��}�\�Ơ��{�^U\�DH���/��5C|��>�a�s�r�EJO�~��Š��"��,7��<������V�ְERI#!]R�|h�궶̛+MU��]���䶠J��X�Y�����}��Fzb�D��`��;��y������q�����h��>�B��3k!#�ؕ^��\�P�[�U�:�vƉjC�����+z��[��Jڷ����ɬ&�!���:d^!�������i.�v�[R�k��Y��E����B����{�S�����8	�����I���T��cr��T�-D`�-�jRv��lb5�Em�"DR��*�^Ib�+ �P(��eb�+F�����6U��1J����֎kȢ��U%A֢jX�j�Ռ�Qh�����"26¢��jQ
IX�E�q%H*��IE���J�`TZ�S!Fu��X�B�]��ͮ�f�bj��iZ�6�)mS2��Xs���J�F2��9j�@PR"mB�*"#R�ejTG$��%A�*(���e��ԱQU�*F����s+"�Eb��5�[T�Y�5��pр����Z�5�
1m3QH�E(
)�B�`��UUs`��B�J�#Z0�T3�	AJ��38����(��m�
��"����u����z�O���Y�}�����J�IP�x�?ן��d;N��7ݞӿ�.��m�s��<a��3��2R�ru��W����%��;$��d��]���W��$��d�2L��s���'��30�
�����v�^�_������\V/H�|��$�����XJ�D2���yk����s�x�i�9y�ތ��T�
�ِ��߹�G�<R�)���ȝ&k�*�P�	P�I�'Y���Cĕ
��!�T����;�I\3$�f|��=�'�ę9�������{������x�^q[�R��<]��Ľ���%�v�F]W�9�f֮.������?xF7+�Ϗ�*}0�������|I���!�&O���F����\�!�?}>T$��	0�����f`�cq)=By���uP��d�
�'ן{ђq
ò���}�w.�^q��~!�Ĝ߮:R�"Ġ^a&�����lk������{�C����2a2L�}���̓��$��I��>~����r�!u&C^μS�}�������{�C���t����������9�:C��C'�οtd����Y��������x�T*2��?z<9�p����9����Ĝ�t8���쵣}��;:��WFd��ϟ��C��8�8�ټ�[��")H�bLy}?Mg�}x�z�Ğ3�rL�ԙ=��:7t�!�I��*�����v�O2'BN$������j�Cl4z�����g�Y�@۸@D�x"��.��P���A꽾D�#�#�x��j:�B�I�
<��������?�_��C�t3!�ɓ��ߺ2�Hf�?���M�[M�9�w���g����A��I���T+��~��J��e�F�m���,Bqy��珮����d��9&f��sޡ�r� ���$������XJ�H�q':k�x��kjN���B��8�(L�١�B `�;E�6͸��B����0eAy�^��K��������p�]ϡ���d����;�t�ffC33!��sޏ#<C�d�d�
��o���Vy_�s�>�̛������C��?��ތ���d���3���~�C��8�&?�վsq�ܯ7;<H±9�{�l��,^s�8��_1�������*g̔��^�'�I��a�gӕ���C$�Vd����uP�3)9�<�N%�����ձ�uɕ����p<N���^�^]��u��u�$�W����A���q&C$�V}���V�X���/8��-��Wջr�z�L�39&fs���{�<C$�_)2��u���o��C>���+q�����*�'��_R��ng�}ퟙ���2��~��g�q�����1����C�C0qĜ^t쾇ە�Vf�|VW^}�PJ��g�����x�q&O��=;�r�y�tt��+�믺��fg$�`ԙ=��������~���wo����ӏ'q��NW��8�	8�M�fa=����T<g���3!��2}���G�'Hf_�����a\G�\D}sP(S�ި΁<S�.�'��sI�����|��,�`m��Z��C���xzz�[��B2��j�];5��~���� ���m�d�;�Ʈ9Ns��N��g[^wi�-��]Wo��-�s�5���ꎭi�5e�6�۶��t�y�Q&��fR`nح�z�wn��0k�_D�ny|Z;'�����i�x��[:�@;9��.sˮ=���Zf�7l퇂�1\�5;�3��G�m����Q�[��\$γ�pݛt�<s��N`.g�kk$��:�٢hʼ��^t�l6�g0q퇱j��r	n���y���kv��<�����қ���ns��d<a��y��{�x��cP�6��{��u_ �g3$ɓ$����tq'��373�\���q'��z��~�!��L�IP�����ߺ�x��!�>�疸���mw;��v�����OP��̆g>���s�;���O����{��3�8��P�d3���~�x��!�a�d�S�o�:8�T�N/0�^p�:Ķ�'j=$?�3��=�2i��[�w7m��s�ĕ<�<�￺�<|I��*ԙ>��ʊe�we�q���NM���w�=q�������=o�C�2!�Ʉ2����l�fC33!��L�s{��;���)�s�;����k�w�a�Iͯ��/��y�����	��K���95Û��:���g�2%Ov�ގ$�%gnI�������x����7
�1}Y�٫�$ҙyĝ��QW<C���C:o���xV�s���;�Hx�D2~���G��Hfa��̤�}�����@�A�o^kJ:yh�	ZL�a��ן��x�3�I�O�����;�I\̓!_?}�z�i��S_]�����"[�}�vzِ�@1��{gu�wm]�^m���pg�aq�}s�8��gO{f�bL𘈈�@���	�,����J�IP�ԙ=���I�*J�+Ǔ�9}�d�P���$���=T�n�d�'��C�����y���fh̆C&O�o�z8�bt�a�ݞ���9��m��s���<�C<��{�;C$�����,��e���C�bY�Y}	�"���Fx�%_{{���u������^c%���b��|�q��wZ�g��Y2Ƿ�?��o�@��0�w���?�$��d�d�7�����$�v&I��$�ß?��{�<C��L�ԙ���y������}�\C�J�~��Ϊ����mw;��v����:8����fC3�9��d�P���$��	1�lV|���S}�g������!�Ð�0�2J����GvuC$��d+��sޡ�x�I���y|���vw3�Ύ�T�0��u�s�<>�����>����T�3�rL�ԙ>���2J�p�!�����!���L�C0���������߾}�u�����̆C&N�����v�!�iO|�_�s�7^s^s��!��y����q&��I��fo�~눨^a�LLl3�ߠ^�r��/���@��2L�9&f���sޡ�r�!u&Cia�?�����a�����y��ǝ��q��(r�s&��4��y�p�'�tc�mY�t�u,!�sTp:��������4�W�����C'�n�tq;�t�ffC3Fd3�sޡ�%B���������%g��$�uS�����=�v�	h�.�\���ĜB��`̓:3?��sޡ�x'd�߿>�W��S��;8���&<����_����qyě"��O�qV�ӫ�,w����$��	0瓉8��u�p��D24C!���?����^a&=g�Iĝ���d��6z�p�^&N�q
�����>|�9�M���|C�G!������q&�2J�a����\C���3$Ʉ�2S�����~��|����[ŉ5��Z�O����B���N�_��}N�}�R3z=�ɿ�S��}��~���籤k�P	0gf���o3��ל�ǿ���׿㤜O�d���3G?��sޡ�)2���?�ߺ�>2�|y�]�x<.�]��*�L��*E�_iǎ&gxĸKRT*J�{��{����2���}�����<�a�!�mG��%H���2�B�q'���/8�<�}�<�'�ę1�{�W���^ky�nvx����y��u�;IY��
����%My��I�~���a�&jZ"w��K׶�����p���S�2�'����*�3!�T�o�z:I�+������ۿ��q���/�<l^A���-���ױ���u
�N2'\��'��l�{����MMח����IP�?���A�|C�1�d�
�����\|g�3�d�4L�)��F�)�T������t�ee��O\�����x�����&C0�~�����C7���o&����9Ρ������y�R*�8��Ly���}~q����������x�ɐ�h&C0߹����!�!�h�2M����ʑz��N/0�<��Ң~m�����#gʅb�y��w�V�C������fs����fg$�cRd����u�'Hl���[>}�n&�����C$�T�d32{�߿��3�d332&�{��N!XT񌸶Q3'wxx�����N}W)m��o��:��w�^a&�;$畿����;I_d�4L�&�?{��N'q2L��
���{�;CI9Ͽ}�m�����1�b�Z�k��&ͬ��A�-�I�uB��� ��Vԙ�"-��'%�.�gk�k,kűS9Q2�Y���>^�&�I�7����V�^��W|�mn�P���!�s}�GI�!�T+32����╉Ot���}�&����3S�@��ĝ���y�|C�A�d�
�jow��t��T��fI�����y�%O�����z�{��s|8m(R��i6ۂT�mZ����Dn���ݍڵ̭�����w-g�O�5�6��7>;IS��<���i+<�I�Ƥ�~߼��N�ړ!�d3���ޡ�'�C!������ô8��w�޸���fC32�7Ϸ*D�!H��Ee|'�b ghhh��a��_�~�x>!�MC$����}f�Y�1�B����Ϻ`�z��q{&L�%��󣤜N��2%fs��G��P��L/0�$�}ұ�6��_��ʷ��,G�L�Kc^�3�!�"";�I;�T����Ї(2����*G�I7��I���U[�]�2v�z/���*���2Ljo���GI8�I^�̓9��߽�<O�&M~x��Q�'�g�d��>���!���j���'��rL���%��ގ�):CiI�Ό2�����x���!�ɔ�I�:GݳV{�|��߈�m�18̆C&M�����;N��1׾�|�;�k����x���g������$ơ�`�3w߿���<I�����|���q'HT�=��{:I��2L��3|���C�<�Rd.)2��ف+,�q'+����1�yi����W}w�����y�'� cV��D���yyO�u�zW���LZ���Y�al��|�2�0������/������G��:��٣�[���8j�7Z4�\��ƻQ��WJF��+����^��Yݼ�\���z������O���j�.ۂt�=�۳�x��<ņ2���Vq���dE���^n<����7�������mu��mkdXty�/��K�g�a���;,��b&�v�۵���о�s��
�&�a���Վ:�ϡ+��/j�7cl-���-��tԎ�m�p�=On����;�K�ز�pny����sϏ���<��l��!�'�ɹ�{��vt�f����g߾�C�2J�C��f}ϻj��8��Z�~M������S�jo���GI;�P�*%p����{�<C$����y|mܵ�^���$��'<�>��y��^a&����r�ٽS��o���'��d2J�t�ߺ��x�O22�'����\C�x3	9�<�N%���_U1Q�����t��t�a�s��q���;^^^s��!��~����$ơ�T+���z��qy��qy�m��F��OK^�H�L/1�^s�9����bV�Rd*J��������v����q-��-�9�w��<C&�u���~�-W��α*c�yĜ^a&>��eZ�CD�d0��O�~���!�J�a��2L����GI;�ޓ?{�`�]I�X��$y��s'#'��~�-�:���g�<D��V'<��������9&CjL���Ύ�):Cwͻ�k�%��q'kg��ĜV$�d�
�'����\C�x3!�T*y��>ܩ�H��Q#�n/�h�~˕m����W�]����c���қ&�I�-����3����3=�$����;�o��`U��7��!�|��G�8�MC$ơ�_~��]>3ę�̓&L�&7��󳤜!8��;��ue��{�_�G���NRd.)2�����t�i*���ǡ�<��l��<C��!�s~��EK�R$��	1�|���~��U7�N��39��~����g���f��;�S�R�Ƭ�ɵU-���E�k�W��I�睚4{�տ�^��Ҿ��_�zĠKd2!�m����}!��a�!�cS���$��I\̓?� �Y�59�>ݎ�+qy�kh�{�m����T�3�߿���30�
���~��:Cb�!�0�NV*4&�i"�(���>���'�N%�!��/������3!��d2J����GHv'Hf	����������&���Ĝ��:R�t��͜��*��2Lj���|��x�!RT�L�&��y��N'i�d*J�9���O��7B�돺�㗨I��e�wM����κC�������q-����ns�t����M������C�303!��8��f�J��%Q/���T����͚���ɐ�4��{�}!��a��IR��y��N���W3$�f}��z����I���y����)���r}��ț���@)�;i�U�6nx喜��k�����[��E�����<0�"98�b��s���I���39&CjL����$��L�s�q����!���O��|��:C�v�����<g�2%B��&�~�;�3u��O�㹆ݶ��|C�9������$�T�ofߧ�^Q��1��ss'x���:<�2h�&L�}�gI8��I��$��s�����x�IP�&CO���>�wwȺ���'q�\��?���'wu��!�yɹ�{��v�Hffd332��������L�C&D��oם��YfM�w4�(��ې��k���$�Z�]�1W_��^r�Th�VxС%m �u�ۣi5uH7��hSl��lh��{_��n���%��	3��2M����Ύ�w:��W�3�g���=�!�T����owm��^a_���ݳ'�3V�Z��7E�g��jL������):CiI��d3���^����C&�9�B����W��,�o�I�a�qJ���}!؝!�';���������v�x�3�����x>!ěP�6�9���d�g�^r��>�jQ���I���y����'�2L��3A����z��d��I�ذ��~��x�a'/:����L�r�o����	� Lb��Xw�<M���A]0�+�S$���v�>�f���4����h�BN'ǝ�"����fC3�g���=��!�4L�CD�f�>���񇃐�_}g�?C}�T�%b���=�t��Y%s2L����=�'�8�&=�����qn�[�s�$�<0��w�\g���<�qyĲko�|�����s�J�e�ؤ�g0�g{��^�����Y��?���x���3!�}'����[n�:�UO�ʑ*B�'<�o�����Vݶ��|C��������IP�0j�������d(��L/0���B3�}Pѱܠ^�_��d*J�������x����]I��>��u�;IP��|x�;}m8m�nw�bP+HI����R�Z��xs_�X�|��;fC3Fd3��y�G�<C�h��!�~�}��퇃��2�N/?������^�}����)��b�Z��-�v��{u�ڵ�n�S�dў�!��|�-�U����{�x��s��M���5�ν��ة��1���$�_��%��3�3����!�T���<�6�4�^���$��&a�?�u�x>$�T��2���Gq���<��~��WE�@�����>����� &�P̬�$t䩝��S�Cd.Zl㣮R�F׎�iy���uӧ>�Gn�zS����w��ߪ%Ki�ct��y�o�S$j� /cU�n�ӷp�;�e%j��Yd́�����z��8�n�xZ���3ލ���^�@��.�� �����'�1�s�/��{���Ȝ6ʝJ�����7C��?_��Ԯ���: >�=�v Ǳ���72� �M5s<�_Z��ҋ;���@O��@L���T�r�S�Q���9=1�5 |�ճw CȶL��!�Je'j���@L�eeg۹�`FoU��� z�C$�"�,����nL�&�=�ɩrF1r3�YP]�цz����@Y%�}��!�\��]�	�ݞ9O�Z���K�_s3PT�R�M��Od��OQ��L̅غX���\Ϧ5J��o��)d��:Ѻ��Ddc�{^\���^S�ٻ0�75�W
�t��mnj���m�Ŝn�q�ZZ�4�`�8e͉��8�B$����]�a5�S��p���197c��q9�'Z5t��9�;��-�Ý-6��a�����g�a�3����{1���"~�r����T3��i����$����߇�4�e��.w���Ѫ��5�ë)P�9]#�t$����ñ-���Å%�Q�NZ|&zno� }�j�4����e%0(L�x�����g���6�W1����S����� �p�Oy<���)Ҟ��N<{#�������[�G�Q�����M�K��ܒ��vL�C5{�REmݢO�ڛ���㻀D���g{��n�x���D�3w\�=��9�d^����<=��Ou[����z)�\$I�F�����ۍo�Zw	�\��i��c&/+�7���>œ��\B?��=�C�?�Wr���F�<S���+��6]�'A�[��TN�X�c,����}�;�Yޕ�vG��]m��%�b�j����I꭛��z���3u��j�Pz��e�!5먧��x�����O����=3���͍�xcb��*N�l�ن�*i�+�w��Lv���*R��t�m�-ͩ��u��r����ZP�0�=�Kp�d#f')?EU5)U��\���Y�R������*T�`d��zxÃ͔-�"��[T���YPmFQ�TFҵ�E�IR��N9"ŋT�*��+��E����X,FE�3"�e����KJ��ʙ���UUXJ�*R�ȹ+uS�j�l[h�R�X���DX+mx�J��T���eb�X��0DD�b��.�0PʅjȰ�b0D�Ŷ��QDj�!Ym++*�R�"���@U�,��*�+EX�(EP�[��Ԫ��DJ�xِFN5'�������db%AAzJ�j$F0*,���5�uiG�W��Ö��V)H��J���^5�Pu
���PH�bň��"r�]N������\d�ͳ�=�Nt�,��;��7n���	lkA�o�~F��t�v-l����3�ܺ-ۯE�����M��KtÛ�����ѭv�{]sA�v-�/"أ.���U�t��4��98�u�s�ю�)"��=ۓl*��ֲ:��n74�r!��#�筺vâ96,ooF�]��c���\-�g�b���v��츼=���]��ےl��\����q�3u��=����3��^f���ឮ�n�;�sg����N�n�wI�\9q������Ep�:綹��69���t��ma7F��ݱהq�瓁�8I�qð����۷<W^x��ܽ�f��M��0��pcث�ݔ���h,sqx6��I�����.�s���d��ێ��p&⥹�k���Ɖń��[W>��� s$c���k����;�����Z��
^d�n�+yg.9������:�b���;6�FT��������Υ��}5��X���J���wϘ�8f8��t����vl������Ӥ�	NL�Y�"y�wF����\����2x5�v�t�q�Gz�u�����p�\vv�"$�"p.��Y{=v�t2����{]����;D� )<h81�xV�E�emu�pb� �l9ݒ�m��z;<�}����klCm���mv��˦����gʷF��r"3�ٺ�^v�|��q˷J��=q/`�5����ic���n����f���"��$����ݸ�kUsr�֬��m�5�ILW<;�Y���Ť�4��3�1֎v�n�fH8��m���������#ڝ�#���b�SZz��qץK���m��;�ۣ8vn���nݢ��m�#��-����ں}jI8��n���S�8y��^#LE�������z��Q��:Ԙŭ�pTe��;�;N�ܗp��5�8n8]���6k�:�l��G���z8��n��b�c�w��.&㵋��Q��+��^�c���6=�ۙ�=�Nz�J�p�Yn.�Ϝ7|uI���،��x����qon�	Ⱦ]�qhUչ��<����H�Y�:�ݴh�+�.ɭeC�ɷ>��u�m���]����O�z�[y���=��sp3�f�/�1�G��o[۱�����Kv�v�3�xiɌ�܈ tн[�[�z���k�j�N�1z�T�{-�癰�I��m��n]\�u��X�tl�0��nrE��n�P��G=gU;��u���cZ-e譊Kl�q6x��M[�(`�8��r�Km�����-M�hٷU��������� lr��������W�� 	�m��� #��,������lZ�D�-�u�w2Dn�}0��Bi��1�W �V�ֈoz(�������, �1m�@@oye�&g �u1�9��{J���a'����m����� ;<� ����h���~�@�b �!��h#7hؖ�Ȝ$$�sԞ��/sa������S7r 	���0���w�Y`@�p�=���8������}!��:f�S&D��Wa�k.-r�.�i���l[�P�+֦h���v�>��]�����IK¥�l�pD�4� ���8�&bP�;E�=L8�ٟ^7����K���~�����v5���2o�33�nR��#��3�W>���#I���z��g�˶R���C�ӹ�+���� '�{ݹ�ݧ��goR�"L��tɇ ָV'c����]]Cޜ�luN�qK4y�{\9�g�ڂY2��G8O2� ���=,�/.�$lש����AS�����{˲Ձ�ߞ�w�u�����Η�L*�)@�i��n�� ����[�M��/_+�΅������v]�H�7��v�I���$�L�j������ WȐ?C�� �y�p�}ǭĻ%'��͘Օ[9����{��Kn$Nl�:�ix�$�!�\������,��G� ���=���[�f��+ʂ��w����h��2Xvɵ��ک$֑�]�8y��Hz�t�o��~��o�0aFf�+K�V@f���" 㗭� ��}�'ۓ�f�[və7��w DWE�d�K���N��7C��uQ�l��T��֎���@k�.��[S5���S����|�R	���	�S�y���ɒx�u>��>uѥv���\?W��3K�"��n׾s2�ѣi�Pe���y
r���q������ŋ�����]��	m���NA�>���j���\�� ~=n�L*�!	&�cݫ�w<l-ف_k������d�� j��P@w���6�c�K��t�x�� �$�d�m��m��?:��@|{.�{B�;wfn"��e���n� ɷ�.�Cu�)�����j��L����X�A��V��D��ftl�RK����
���{�tKn$Nlރ-׋��pۇ '����3hՅ�g�]��R����@| x�u��72� �4��W���i�g�Ӟ�9��X@��@ ǲ�@cj}�&���1�~/B�-@O�J�	)��)��y�0 ;���#�>	-U�]��K)n3�@q��2ǲ��uN%r��	�S/��~�����Z���|nR� ;��^�˕��_��i6;�u�#z��x"������\���x�":��EԔQ����Na���]�B�ڌg�&f٣./V�}�)ϓ����|�Ǆ�I��1�W��m�Z ���\E��#`�ޜ�K����U @��,��7��w�*�7�g�#vN��[~��Kw�(/��Z	N.�u������#�if�:��Hs�j�V�L}���[r6�w���L �,�� �[�X{���ƶG�����@�����G�Sp	�Bm���[�., �ly��N�榀���_�������g��i�&W�X<�#�ne2i��oU�ր9o��ɒ��w(e^�8�=3�������Yw�$y>��p�%K���NՉ�=~��	{(&{�[qh��׾.�	���U[�k���x��� 独��npv$��J�	�s/Wa���y�xȜn��{r���y߂��� Wk�`@r=iO��&b߱�-�bJYA����P������#:J����Q���5�[M���owA��7b�f8)�ݜ��;��]�ǭb����a���ۿA���Nv��.����;�Fco�L��]�5���S�����)���j�8���k�l����Q�;J�G6� g�l���^��/b�d�uj�m�mە�˭��\˱��]��|����6}�6���M��ynPk����q��v�\�Z�u��#wc%j4�g<7e⎹�#�3��N�{8,�
ՄN�Y�R�y�%�sj�Q����X�
/)�n�>{ �j�zC�J\y���F{:�Q.�=��?	$�m��޹��/- yo���d�K֔˳���\�� ϼ\�2mL�d��m���r�|��ژQ�w3��ۋD��}��o� �z�2@=�o��^Gb��F{��)��bi�OR|z, �06�2d~��<��⯵V���}��@L��Z�`�pٙ�S &���r̞�Ѕ�n�Mo�T5�T���u�@�,�;wTz+]A'=/�櫊�+"��J$�Rv�H�Tɒ��:�ՁY�V�U��z߬� 1j�d̅�,�BW�J�5)��n�//��RuCv�f��ݣu��8�Ƥ��F��L�J�M�^`v�'0����+_�\E�@�Lf��Qa���]�<�5owr^²d5iMD­'�M�"[v���h�;rv�Gs$#���_r���`�\�daL��P�2qN=-�5�Ywy<�����	%8qz3vA�SlGN�����χ.�L�,w�w�37������W�����SR� L��
���}����)$���g������ �NEE��i���ߍ� �G�T2@�Yv�3^� �!2\��ݝn�sU�K�鋙؀�|� ^���s��Zٻ��U���4f*�>�r��%2i���YZ ��[���}���B. J�* /|���L�������z��)-YQr�%/p�r�%D�Y��F��b���`����~Q��aj��\�����8ID��~6�0	��Yqh� ;���
׵���A��Jf� ��m�i9��L��0f�����?}[FU�^�Ʈ2|۞we������7&=۝kؐ�)�}0���LD����[qh ;�|T� �<*���w�B�ȾX��%���55$�Vw�.�_���[9�������[�;l����Wl�ёf'%N��ӊ�8w�E6/,!����?��}���_�	����'�G��|]�bɓ�p��lm����J��9
9������������U�!ȯ/l1b�F�jڴ{�� �!2\����n��� 0+UC+,���lH{UQ3*#���&l��.�  �W�3�ŕ�_�5S��fP�(���|C`�/lY86�<�t�v}�?��l�˾m�&/����w�0ee6g��YE��p�����J���ث�Ċ���u� �~��z��q<���Q);WEj�L�"�r읞"���m)�/˙�C�L����/���yZw��|ǎ�k�fr�r S.�M��.,�����L�]���]U |s�.f�9�P�a퇒�LD����չ2�[�q�Ep5�S3/�Qv } jU�T@�y]S� �M����Co������l��߹�n/�ynSʵ��%��]���$�Z�V�1�T��d`װb9i]���O���'���p,�:.�ҒI7���ۣ�$�������� w����%��@R��v���L�'����{�{�}d׮'OJ�H�+�JY�㧬\��� v��l!.坎`ۋ��U�_>��lp��r�s|j��v |ʘD w��a=�:��=$5�g_�h A�U☶sa}D����Upֲ���
m��{�.gf,��4U  7���$�็*����fn���M' �Rt��J�*!��{U�Z" �ɝ�v�x�K2  EyS$�'����Հ��̊e����o��ۇ.�3q�־ 070�&Ov��f�#Wn+�db^���{��O�⯘L<�:)���mۙ����g�n*�WզV�ey�vנ2N�j ��y]�ȓ�9v��'2�c���a�����j;fպ�<;�e��K�R�~B�'!�~�ܺ�\��Bt���O�)7;��ј��%O�nx���1�ꡲ�1T�-f�/'�M���0΄���Y#�"����gu�!]uۃ��.�n���X����u�E0ܜ�iL��9�V���;*�r6�2�-��ׁ��<���]����h��d���c���p��nu�c�5m�\��(��xm��M��8�!ڸ��9ȱ�,][�����έ$ۓ���ы�Z�׃TI�=R��X���I���;�Xnϥ+�P穀`U����6�M���v$�j�u"j�㎮��u��/T{.uڿ���'G�lI��m���%z�� ��֏��5v�z��'w5pt�x�I |w����f�= ��sNj�WZ��&Uӽ+����Z�y���"72*����?m�W��&h��Ы9�EU�H��>�!%)��`+�e aۊ�� ��W�w^u	��� ;9]�B&d�ۊ����$ND��X�V�\F�VE��mo�U-��v+�� �U�V�̺+�W�n�_��]v�=Xn9��\!��f�/XySc�zП�.�" ���/��#V�+�x+ʡ����zY��߽������5��E��v�dz�#�#�c��^u�[[�[�G��ܭ��I��Li���9�<^�DǷĹ�y*�NT�l.�S��,���h� �[���œ&ܱ�6�m���C�L�ŭ�o��ڣ#y��l��xVKM�A]�p����S����q��Mý���&�^��q���7ק`5�{H��	�K���X����r��h���[��7�|������c��SQwϛЃu��$NQ	������S� 06�0�mFⅿ+�ǳ�նL��{�@ �Z�`�`���0���Wpֲ�W�����*����V��ɒ�֕|$�Yqy��կ���/��[x���{2�"p%'j@�Jp'0���c�sSJJ�޽�5����6�� 9�L�� ��˸B��"a;��~w����_�ǜ�㍗�j��g�1����1�o�y��5{=hٷU��\߿�OӾ����og�
^�+� >Z�a2oy�Ec�Ge���m盨�]ڮ��<����OB�1�2[t��V�֏��^��so#ԇ����d����@@wye�ȓ�����E��ˀ#�'Ei��4�m���C�`�}�� 3�3�]����}Kv����J�}Y����9�Ǧx�{]�;�������"UW���{�M�6�S�<�h�XEM"�o4�NS���K�c�hM蠦5�r=ڹ�VY�<.�m��C�!�rӢ���mg���-��M������3�
���'=�.t�O0G�33+�kU!p��6Ou�5�?K��w�ؑՆ��x ��&5��pܮ�"8�o+�s`�ٮ:F�hK�S�껍�5l�^Bc�r��o��]E�A��nrǻZ9�**�%޹��%n��3j��tj�>9��-�[9��q�l�[�@"��#v���{2�л���	ܱ�ܰOsR����z�)��#ϐ���:6��"�^� ��4Q��T\UL�CYf��>��e��gu�(/n{e�J�l�n���ގ�N�}7��?nM�D�����*q�͜(a957���,5�9"�L�p�;�/o�<Z�(��D��pz`QW|�p�Qɛ��޷6���1�.:6�k%v�څa@{�7�5��ޞ����[�yďה����q˵�"���#�+6�`4]Z�or�ʐ�Շ��/���7nޯ�`���hm���1�3��&{��;�/-����(��/b�G��О�[���靐웪���%�b�*M2;*�x�����2�
�W�G���c}�����A��%Lm��w�����V��v���d�JL�ޠ����>���b�8-��9j�7&���/[&BA�?�E���UCY+���*�(��T�����$��.r(�6�:J�X��A�ے�1J�əX��X�Tj,U�D�VDUAf�C2h�jT�ɅQ`�F*���%V
�����+"�bԨ"E�L�QzN��zaTԢ��bT9��FҦd�gR�EE�E9kT��!�Rd�ZU�R�J��� [�7-C=bΚ��V�W���iUR�Vq�"��)3QU�DD-���b��*-Kj��*�X^YYR��"��j[G�VAIYkJ�r*����,EEzkh=cDE�TY5(��աY�D�ձTkƧ9H<�G^��TAE�*��"��hlN��2���<��xرV(�lm+Z"�Q`�^5�
�X�1X#yzr�bʐP�)\��
Y�mR�j!��Q��Q̨�"(����N3��;�~���_u�ڦI���]��s�I&�Kna����V�[v�o������䦠 #{�,� �ۊ�1����땹�l���*�eG�fb��|���Up���� aۊ�ȗ��������@RUiT y�.�$��gD{�y\���G;��}?�o�>�m�uKx�-w
�E1�]���Ř�ּok��
r���Ϊ_���ߟ���.OD	�Q ���@˷��=ݹ�#:�}=*׾9�D2fg��*�vXȸ�R�JM��K���󲗕�P�.ט|$vs�. 9v⻀|>I9�
��/C	�v�DƘ�m�\�V�Z =��ə��٬�o%-���{ڲ��I Dj��v,�J�4�i4�m��r�lK[�w9z uymŠ >���v!���-g�B˓&�ڙ&:c7^]���I=��}҅��p�@�|ůt�iA�*'��0��߇����"%A3.��oe��J�ff۷��n�7�$��m�$�՜��\Y2ڨf����d�� 
x�ˀ ��⻀ ��z�1w���K��k�n�2�Ai�7,g��V�x�5���nJ��^2�1�a�z�qC'�降5����
�YZ>��{�X��zҙ��z7˸��;�e�Ȑ�]خf���-��'jč���if��+��;Y���2G��+�> �z�|�>	�vZ��<��Yx��춈�L�	9���{qz, &x=j���[ﻖ���� x��S6��T�c]��țI�n��:�o�a��*�y�;m\E�3&%��|w�^�&�~JéO@	{5]���-(M&�Wf��Ẁp���ozx�E��[�ā�=�}���1�P� ���.��l�{R��8/��k�3oڤ֟w��q?� x�Mu�]�����{7[ބ�uu q���+v>4��S�@�5�n]�ݥ�7��q�M���6�����۬-ۤ���l\����a��,p$8|[���@�v�Ç�M����������<E�>K*�#��5[�L�pn�s���a�ю�G�M�v��;���h�!��==�|�eM� ����<�3f�z�͑�V���ua���F���ݓ0 �Q��9��qݞ5n��<E��9.L2�-C����\i�Q�G;l�ێ������:n����]�����~�����NvloL�ڦ ��\Z[�wG�z9]j�x:�0���f,p��R�j�+�e�:���_Rʏ��, ���J� ��˸D�n�y��yz�aغg�h���8I�8I;r�S3��Yqh�&J~e�:g;����j6ҙ���+� 춈�L�	�����]�No������-��e�䦾� {^Y3@�q]vL��N`N�1�D�i4�m�L�ջh 8�⩉���(�zd��P��k�{�N�6�m��f汙 ���pW�.sX֧���܈�Q҆�V��6��nT���z�<��I��j��P�S� ���/��>�ۊ� 9A����F�)���v���s�ԇ��0�sw*�W �e�1��뚿M�KO<ڬ���X{�t&3z�}�����vXv��Vo�6�kҥ֜����^��'"�Z��� ��ՔXL�ۊ�f����7 ���D{��&,p��R�j���Q`@aۊ� &atS�;i�Z[ �eZ$�ӷX֍�!��8C���p$m���`3.��˦�S���{���G�^�W`@r=k<�V�Tn�J ����~�h���p�8n������M��W̩�L�$��==���	�=���	���U<h�.bV䲝�j��ْ�5voY�ng��:ݍ��;p�ָ�s����S."[����S"M&����2�mڙ��ۊ���9/ZUj��=�����-����������w��uJ�h���m�s����&qEϻN��#��9Uڙ ���v�z�C$�'{��J�۟]����Kk��o9�Hp؛s	'7pr��Sp�S3_����d��d�;�ܖڙ�7�?+�{�>/^���M�pn{�c�S�	��,���V�e#e��y���]oT��_ئ1<iw�<tɫw�����_n@LXᯐ�4��u�CkM�G�#1��p G{U� iP���K,��RA��@�'���y�ig�lƆ��NN��$m�� {V]����S�q�c���&f�3$��� m�Ա=�M�
�:X�:j�����;�)�L�S̝�޽���cI+����ces����S�\�5���)o���	�Z��}�,�1���[����~�v b6�0����(�SCn�Շm���X��Uv�a}��o�X@L�b]iW�@nr˴L˜VS�t�5�^��*�1d�6�KCI����~T� ��,���/��d\(���ų33aԔ�w�Y7�4MK��D$�ݝN���>�{����ft(/ʡ��=�$��z6ږ�<�(��\�켊�r�1�uRt�T������5�u�_!g?�PMl���^K��Մ�;5��낲=�<NY~�Egt��T0�;�HE�0%	��¶�\Z� 3��v]�����π���� 3�e�7��
��}���"�~��Z�n�]Y.TX����ήa�rw�|�lk�xls�P5;�\�w��?|6�7+/�
m�d��o�e�>���`8z��=�?^|T�ҡ�DＲ��춈.Æ���w2�n� ���x͙m��B��7�Y3`}��K�" �%z`�P���s���t(x�M!qϒ����K���+m׽=��,� �3ܲ�2w=���d�L+d�Si�w�ҟ�4���j��}�֮�@��K�����.�c���`���\m��A���&��I�NnΧ\\X�I�S8�);=j#��x��ɛ�"3ϴ��>	�=b��a˝�#gVs}?m�&4��Զ��]}��ZX�:7�w��tF�b��H��6N�a����WK�����w��>�w��M�'���1�v0�4x+�ֶ�>Z�Q��wk�5v�]����{Fѱ�I�	��󔥢��x�j����74S�I�ݵG'�F���l\�\뷒n7'un��4Gg�q�Wn��m�ɀ�G�k�	d�F��Љu\ �v�&�0��h�N��[��$DH�:����nb��M[&�<+!�i��<�u\�]k��.�-�l�n5KF�\�\�6��Y��ս��J;�`��<yn�j�Eᾷ��j컪˯7/?���R�8jKi��e��� g-��,� ��z�A�5�[����JS�up� �|�K�#����	�%�	'n�+l���ڌۨ��洷K���{���t�X�j��2+D/I�V*�G� �?8j	�SpW>�qd��m�� #�[Y�z|���~&t��.�	� �^��/�|�a�2ہ�U@z�o]�A�������V7�L����f�/ye�KoC��ZU��v@!��.��o��#��4ڻ6S�_0������-W����d��w�Yw�;'YQ��>/ye�6�L'���>�oӤH�m���M�H�v�n�P��u�d�C@�l��ƺ��uZ����~���!��9��O�E�@I�S �>��XW@���T��op��>:WY_0�sq��J[L��]k.������l6��m�	����f�$�`�u�g��[������ܝ��h���_�<�\�yOӪ�e�Gi��E�f/x� ��*� ���YV� h�����l����1[ߝ�@4����nɐ=�YZ" �Ӷqt�.z����i�%��繤��n�.�����u6W��6v��{�3�&aPɒ��\@ F��f�]ҟs�V��{	'.�{�pWX1j$����*��<z~�@��ʆ��h6K2 �Yès���|w�x��t������9V97�$cd2�1�����*]��v�=�@�uv����N��s�����>�~�3hi�skWG�@o��� o�x���آ�i��-� �8d�A��웏F?JJ�QTrzW����&�yw��=����59��>��ye����.f�;^h�=1u��Y���7QA��LZ�p�	K��v����yw�� +�����K�^f���N��VlIԲl��5w�N =|^��oՊs2K���]�]M���s�{��M�'��5���V�T:�.�<��	��{� �~���nb�ӏ0�	�⢐�����>��]}U�	��u�h� �y����G�w5nn�iL���շp��ڒ.�����w2�n��	�Ħ�c�n�uz^��g�w.��d�;��v r=���IDR�!�O��E�ۖ6���U��� V�cq�WJ�
�튼�R!�W��&s-�)�} �V��v�M�� r^Ī�Mg���/a����D��^�� ��D��P�j�C�L8�Z�fvq��U-� �7�^��	��zҙ��\���ы=U�q\]$�� ޏV�p��L!$��}>��mS >*��J��\\�u�Q��W�� "G�S��$��Iۛ�t����蝲�&{��n, �"5.�� ��YEfRc�5��e͒¬���Yy���*�OC���Y��	,y��ղ����(�w�#�mȖ�
��О��]�kв�;��te�<�uY7`}��|��NN��$m����g�eB�c�q���@GVצ�  0��3P�g,�F{�.su3�U�8D��6����2�����oBgk]]n�r�\ur^�ն�U��Bx��q�( �&x�ӒiΜ*�3On�@L���,���=WW���[�I�&��wȟ�w��1j$�����-�S3[-[�g���]ʴ�� A�����{�v9�a?+���r"�= �"&ڑ�J�v?:� @w����2e��,�Ψ��g[�� vr�&�cղ���BI���눻��{n�-GY;33<V�a @~��, #Wo��t�j�#_m >U��ۊ-	K��$Knn�],�S a��v9츪٬K�~�>��T vj˸D�.�+������m����z=��Qnf�eŽT�[E'��8�s;ɪ͈�S�m&rH��톞�js�c4�k~~�⦱�bx۩ɼQ���e��b�G�Ol]G�ݽEr��Ff�C�u�-�]�b�S�}����V�����B�g���n�d;��;�9{,E���N=���a�h��u*����.�d�G�	��ť�L�G�o����;ۯzb�)�+� �ҥ9n�i]�%�̛k�І��О�%�}�=���bod
C��}ᬠ�wz��&(�ّ�ήg�����9��Y7�ۄ3�x�2gf9
Fb��'��rj�G`��M���xÛ*���rm�vL��ʖ�t��n��i粧B&u��Ictdk�%U�=�K2�b���R�CA��UL�����)/{�d
noVPĠ���t`�;��zI)`���x�O*��aF��铳F���!�_�ѣ��;o#�o�1�5�"Y ���QQF�L7|'���xN�p��]P��	�j��iji�{�7�2�Z҈��ރ�J=�9xy`GA��%��/6Wn�z�gp\=}2s7��A���qT��X���I�}e��xv��)W�U@y}ѻ��Aܙ����=�-P�_W4�f*�7��;YaS+���&������[G�ظ�FL��u1۵��SAq|_qIs�,iď��馑�2�sb���:���i.�U��;r1���,�u>*�c�O$ߥsm3�*v����PF�q-�t���Z��.���G��>��kZ��TF;�ܫގ�y�tYX,���쏬�-����@׀��"Kmab���PV��i��
�d�i�8̉�ت��V'*��q��<NEޭ`�)��բ�
�8�QUEZ�
<�b
\�QsYS(�*��PF*$]iV����գx�ANl⢱a��u�0��b��a��-e��
��*d�[�+"��z��\�[8��J"��X1��Axʨ��U��TEF,Y�2B�):��ZJ�P(��J��֢Ȍ�B�:��V,��Yĕ��U���E[��⪱V*<eIZ�(��*�Q�1LQE-撹*"�F(�F,�8�F"�X,�X���(#"��
�f��
�b��lR[b����pʂ��2��d�Q�%�Xq
�L�6�d��)��5��"�f���I���#--m)S�bT���AdDX��fVd�0�"�m�$�-b�����[E塭N�X
��(*,�Ո��u�aame�lUb��,]h�B�
�D:��_�p��79�5�u�lnx������y���|�c�I���ݔ�m�0�Ê��r\s�/&�v\m��۱܆-c5�ݵ��c�h�E�W&��퇦�7p� 6�u�0�[;���¶��/F��w=��<�j��۴�phζ�k�,��ru�Q�Ge�vxS��]�����v���P ��q<��b����#.;�cer�a4+r6������=�M�z���s�%n�%�u������ۂ�n��[]��s=�2p��(�q���d�j�(x�8Ŷ��>{q��dl�Ʈ�uŗ�]\�C�ѥaǢ�՟e#��Ӷ�[�t���.Р��Y����*�۲q��n���M�$���V^���z�l������k��S40�g���XV�#;�[��['F�q/s��٭�:�8��[��à��=�r���e���]��t󌪥�D;0�u�ƻ�����Z�<��`�N�c��h�PRBrE�8;n"�O	�I\۳#�득]������ch\�h�Ͷ������p$sT�r*�׀핝�\�\gri�݋D��9N]�:�	��.���8�A��m=�����5Ȝpm9�Kr��^$��+�,vxv��ެ=lm�N�
8C�[����p��S�p��3��K�9��9��v^��b�Ep`�؎����i�㱝�n�h��� �S��fᶼ��N7eU���\ll�j�t�� ����S�S���[	�:�צ璹��x�c��6�@�9��{��Nk���=��ϋ�V� �����Hy9�ڙ�9�x���8��^��XQڛu��]c<��lZ`���y�s�R���0�R��W���v�����g*�.A����B[�����W#.�|0/�z�Ʈ!�{i�֍Ƌ��Y���vv�$�4(=��*�tj<���[�����:0��Xi�ĥ�$ʸ���R������M�sX�Mwn^��@�����X�N{�\����9@���C��'�]�������#�X��Uq�냴v[A��<;�4�]e����x��2���|��֠;���ۮĵ���`��\#<[�[n-$�AK�իZ!�p�;�/k�V��[���D����wi$��t�.����>٭йLm���ԘKO[��,�n;u��'I��c>�sV�uK���`�-٬�^d�9��M������¶���������T��ΪJ�|xߒr�i�I��̙"=�.��/w�̾�1��t���2|~�c!��=�� � �I�{o�?��~�����^T����ɒ ��^Yɫ��w W.|9d�l�=�^���"&*⣔L4�[mڿ��|�U37�v��7mC�N�Z� �=�"@9{����3�"f�Kb�	��8z�fj�y�H/� 9�e�h�#�w��� {��F��̨ ���v�v�1�-(I9��>U2M��6Z�U�u�y�Y{L͍݊� ���c�dd�Wu�����$�\��\t�<�v^{q/�.n|pƻ��1��׷-ʄ����P�Iۛ��Yv�	�;�]�'�A���DE�I�ݽ����Yw�$�<�q]��t���'.�4���FۦL�D��ᛓ���v��>��Jlr��ژ>��3�5������3�rn�^��<�9m���;Vc�+�<�x����^�}v�ƈ �݊�l ����D�(��B�s�s��m�c�O��p �:��Z�e��� �������7�7y{f@@�q]� �{C����(�i̦�7j�ڶ����*76zk �E^+�d�W[T�yeY,n:q���~��[$~�:p�&$�*��C��,���GU����]�L�m����ye\F����w;��<���U�8^]6�9��vymm�<7XoE���yI�gt�+�׶qu|���~��[���$������ '�Pə�7��� ��뜩�ո�{���&x���av^��J\7	(svT�� T��늒�LW[��gg��ɒ 9m�@w�]�� -{Ϊ�Ή�G���V`f̙9��i�IӰFۨ`~����I&��s��ٖ>Ub�j�	g�.�'�(1
��3�Ns]��2,+<������`���k٬�g��im�����ހ &x�u�$� �{�.�u�E��ȑ8ӹ�~�<�R��L�K�0 %��d����� >��w�YV�ݲ >��pg�}�"a�2�`ݫ�{�n"����n;��jU�;�]�L�欻�H��w ��eG���=2ba�i����z�����8�+�vz���OYZ�����x�\K`���s>���������� A��wp���˾�\χ�$�jʴ������$���s�w����f�ʿK58@g�e2D��s6�2�!И��0��6n	�pҁ�7`���a39��v �T����w�� 	��ʿ�$�\�*/!H������2L\�"x���wn  ���| {w��| q�b�wҧ!k�M�ԗ�}���/5 �s�7�sf�Cf�ޏ陷����]�
ˋ��X���g	Ӻު(��컋�f�N�x'�VQ7���["F�N����v ��f(����T��g�ݖ�w_�Ǳ�zy��x��"�6a��4."dqs=���=ۨ�ؚ�3�v���En\Ù��"[���G0ӉM�oW@er۵2}=ێ���^ƫ��Իy/M���B�]�� �oc���[�nR���v=jj�`��շh� �{X @q�jf�'wί1��m���Vr��6_�K!�a$��N�T��38n:a� ,�}9^:\��3�G�v+�� 8�55Xm�8nS����ԭ{v_����ڮ�� �/cU2A��NQ5��+ݕ�2�����%fC	8i;w ��L ��jˋUb�wU���Ƿz1ګ�]��n:���ye\!��uf�sV�5}�()7*�-(sh�y�����6�u��\�"����m�-�Xv���b�&��A�eT	���b��97ŝ�N�v�u�f"�|����v����V��nM�@=���t!ő<���/F2�+p��]u�������Na��ן�6�n�ǭ��Z�<���p�-�M����;d�5h0��]7��]Ԓ4u�v����+�H]!�o1�C7T�l�۷Z����s��q�1�5�=�c��a��4�C��[��;Xn�׮������&z.�`u�=X�<�Yc���{Qh��8�����K�G'���\�j�����v���(�iE�谀 '��P�g{�(�O�6���{�v��ӽW`| i�����g�0ӉM�n���^�D,��Y�W�}�V�}`@b�j� �,��L��{הՈ�z��t;�l��w�O���	(�.�8z��g�_ֈ�Wo�UQv����)zg� }�q�C$����,����e�D��SNnxOV�G��L�<߀�	�-�� 3��2j�b��B~���}H���SQu��A�r�4�m��U+�S a��Y�R��V��մ�/sU2���������2?q�&�bÃ��-��غT�Y�l��n:S��P�u�{�:�͕�&��h�ܸO�G�hc�&�'u�n�D��.-L�/v+��J�M�<NEbS4��M��E�&[Q-2F�s(��o̒]=/VW������ƶcfٖԦ�}�p2��~䔾���r�=v�	��rj؆�;��wW�F�2ʭ'���NI9mQ�ğ��m���&q��Վ��R-�)č�n���m� =تn ��5�^˺�X��@wye�&gN�U`.��k���
E���*�\֗���K2 �u��� i݊�  �z�/C�{�m���u�=�w���׾P�Zh_	9���V��fgmT0��R:��=��������l� ���w��?^�#狔��~skY��+p,^8ٻ�Zk
p�v�K:���	��v_�������o	&>���2�7-�J�������÷�|$G%�J�*��+��^�g@�݊���,X�I����T����v�^?E{=+�eŢ �5wb� '�֫�I����y+�T�غ�M�-\���pӗsc]�W` pm�� r����A�C��꟒��½���K||i��{�L��]Ǜ@#�63��ea5�y�����e`R!':�����MNmD��cN(26��Z�� ���+�> �z�3�q>%�s#h�Q��1������ 8εqa |%֕|���
�w/ٱd� �g���}i��%�<�����ܻy�|����<W�T��yj�d���쫆��݄�W���HZ����툯+k5��쳀�y�u�<�(�]�cW6�CN�����2�B�I��UM��֫�$w/e���Y��W�,���Wp #mW��;2�8m�jnn�w�� ������fSݣ;�œ'�Dj[iW�q컆I ��|����q���lX�I��BwWGb��@�7.-�@�wލ�zt3kʳi�WO�k= |�Z�I��컆E�Z�!5R�.�ƻ|���\�2�y�>
IM Dv�e�� 4��Z����^�1�u"I��,~�@]��/�bpm~~��R�����^`�{C���v��O�}j'qw�ا㍜O����g������_�� b=�_0�b��O�r����_��v�[���݊�<�{����u�6<j�  ��˿� �q]�q�ｷ�$���}ض���ڼ���ʝ6�r�Pcn��γù9��jaķ�o�F�p�	|����a @^��nfd�]��f=���/*��"���@_j˴��T7.e�)D�Nn��U����v���˹X���{����s�/��9v⹛z�Án/��5����#�-��ۖ�6�u�Y�H;qT�L��X�FӌR�R�Z'�欻�Hj��s7��R�-#�wRGS�	�]z䟅��1BI;�m� �>�݊� �>=o�v�_�� i�߶��O�0���ZB�Y������@@OmH��z�7��:��>;qT��zڕ��"��	���F�.G�IwJ�섊�tr�ѝkrY��VBF��v��r��2�EM=���ݘ3�*IӜ�����\w�J�3�����@�2�k�u�]wMӞ�ק�wI�{qˢ/]��`T���r��:
rOl��s�,n[g��l�U�9��U�'>66�۵�ܥ�B$��w`����mK`��'=b��a=���y���e�j���::���V L��׊����=�:��%����nG]5��ѷnWMW ���n��V��=w[��[uI����࣭�.�qkXu�����n5G�R�oL�n6�\�������;�
#�R�{��fx�b���>㗭�u�p��>.�m�37]خ��� ���8�.�8~t��.��Xzǝ�]�o���S3&/v+�� 8��d�z��<��3�>h��؟)IX��"&Rswr��Sp@O��Q��#3:��sW�o�@�خ� ���wS�x��n�I����"l��|gr��" � ��� ��,��썍����zO�_+���נX��)I6��Cm�0��՗kŹ�8�ϟ�� r��v��Q� 7����!o�3Fwv��(��RNc���2[uW[\���n���Rg���ƪ�kk�nk��Bxʳ\L�t8��t��`Z�� �����[JK��\���YQ��j� � ����tĻ� �ԍ�n��Z���]��O��s�Bŷy��+j�1�z�F�J���̨UU�"��q띺�j9ai#�s��ۡ���[/N�]�|��6���h�ˬd5v5Pw�]��=J+��]���V`�Ac���K�l��� @_j�,&J�g[q���*�n[��seÄ���n�{�+r7!6�#p2ӛ��N�Xm8�qޯedϨ	����  #��Xr�b� ���tĒO�*�O�U�@I� �����>�wh�>=د�&�Yn�w������ڨ 3�]�&d�����G���.uOIs�}0�DJx�ֲ]�sZ��s�K���О�yw"i������3�e�Bby\�55 w�e �/v+���Ϋ�y��u{k����� �]��0�pBh�	����y\Y3֖�o�Kk��u�&@75�7����<%;�I����.D�8
c@�ڸ�[qh��Wa�����[eL+��T�1�q�!����ǁכ��f�9��7��%�<����i��������6��	�T`'���qo��2��F�3N�H廳 t�}��Rs/����[�J���-��6n���
L�H�ta&��>��|����4�����铚��J�j�*�iQY}�H튩$Y7p��
��e�*�|3Soq��竁E��Q�>'#�v�Շn�� եb�;=,eSb>��0�f3�c�y�C�Q?S���q���Fy���<�e8d���|l"�U�v�$W'Eɶ�g��(r[�	��mw2ꤠj��ڸljGZǻԈ�Ɔ�U�s��!�N�}�|���5�F3čuսF��q�*�[Z=�FE|�B�q��<ѣ�X$gy������cʬC��ƸǦ2�]��SSv)�z}O!Po�<���)�M�@f��f���u�I��_�=^�,L&��|��5�˽��e�N�=�4���rt��i�Z�gbo7��D��KūU����~��\�c˞���s<���\d��n� ���iY�=�t�:�hcq-eK�yp,���r�sg�U�}�Y�<�v�haᝢ'J�	�'jP�2d�p��4L���9{��	�O��8v�z�[K�ܷ�m���`�D6�����a���Շi�[�$pܴG���k��f�95D>d{��D:����]��&���2�d�P�|�2"��UꬭL��7���"�k=_����h�v
�5V�ڶ�ʀ�0��&:ffL�d�jʁPQV#Z �E�[E/T3u�ʋ��"E��1R(���*��]`�"�����QgIǝm2F%h����eC$�*N���,Qm�V�R�q��d�%ӝZr�s+���E�1�Qu6mE"(�E���)3*DdX�%h�\21�k�b�E.��)y��
ŀ�m,X�J���/,.)iEԢ��,��m	F�VfB�VT��QV��%J�H(q3��QE
�"AdP�����aU2dXR�����X�`d(��H�$�FVJӗ2(�C!��-��+m���J�F�VJ�� ��sx̆@��dV�h�D�Xڪ4��i-�����kkE���ʨ6�m
�YT[e�N[2�EE�T*�"ŧ.�rܭ��)PUFU�L��ua��hZX��]IX,\ �X�T(��.�m�J<r#
~�H���&	$���\�}�.�$�݊�f��(r�s)|�����{ṽ��� b�D r��w�Ǳ����_���W��J�'{����{��l�j-9�9:�v |�q�2�v�����k��,&x��V'�Ǳ�*��{��މ�SI1���\f��5�{vg�4��pe㛮��%ܒ��h��;��lKne�9i���+i]7�v*�� �=�P#��z��7�N�=��I��Xu��92'�4� ͵[2��R�3�%u�Z�f`<v�  ����I�^�*�[K�&�{�/n �VJ��p�.����fx�ug�{���1x+W�쳢 n+� =n��u>1�l�Xujܳ#�(� ]��� ^�� � ��˚~�G�߯�����kQ�M`�;s/V���C;�+�]�,F/{o,6#4j������a�DA���lfdΒ]��up�+�˞�cZ�~=5���l����A�*�˥U;=q���K&���GuL �̹��x�L4F��ɯ��y�hb!��:q�Nr]Oi�l\�Gv����Od��WnBF^�Ǣ!��v��cA(ͩ� wf]R%lj���J['�|f�a�J��H$���_)����<��o�s�����O(�ٗJ�d�r��ל����[�X4B���*�v۔���T�riFsj�rwb���V�T�B�˪kjya���q)�+�v�J�0##F��B����ڟ:���x�m�������b�Q4�'-`7Y<�������u���ѷwD[m��@�s.���{�y���j��[��M���ern�a�|�(� E͞x*�"iL3qZ������K��Qs���8��i��&��^����.7"A]~�?�k{8�8	�-Ub�y���*����S��x]$�"v�{���]�q��T[g����p�/p�;����0���d�A6ݶ�vv�=��g�]d�N�&8��ʇV3�ە-�x1��s\Ϯ�dܜZM�:�=ǋ�U&�3�۰Wx�֯h�Y³m�]9����gzv�4�<Z�b��J�5���ݰ��V�L�غ�`���^�+��oJp�Z��a�N�m��V;hj��"T�*���֡��R���=�3)ۗJ��m��/�C?n�LD�8K���YO��/��nN�
"`P�U�1�(<3t������	�6%d��W�<Y�uH[��AvLr���6Rs��{��3�B�� ���*�gm��zzf6�B���wz�r/7.i @���Q<���H7���m�^���t|�xN>]U*�m���"�����1�����#�{&�kjya��"�K�u��A��R��s��.jWꪭ�^��o!�/�*S�̝W��qǸ��G��Xu��d���.q�:y�:�Zմ[1�ny��yI��;W�����AlF�+�����W�η�
��H���FN���}m�n����2}��GV_iH���*��z�^��OL�=���<��)q\��H!�����بX&�[�~�%�~]خ�d�}���� Gl��պ�g��З�{����:�@�ʗB.}�L�c��78���:y�Q!�v\��<V6��8 z*o��f'��4cg[�_��Oү�fSi�nZnar�؞r�nVu���Y5O(�k�4��˝�=4�f��e�ρd�mV�� �3D��j���ҫ�ʧ�VS:�㝃->����cy�?wq�<?���5c�V�Wtl��c3����=�.2s��l�w5�������m�f.���m���n\@ٗKld�\iM2�� �~x
N��%&�o�VҠ�y�)<������-���̹����޲BJ�NfL�d�bCs-��!��.$	{�*��l�w\:��q?ڟ��c��$z|G�S�noc���xp��{}�)�$��@NULy����2/�j �d��3��L%�Kp ;�nS�7�.������<U{��Z�jr��|�l�q
�2��~����XfJ�O5ԧ�ˁ�7JY����y� �)�d��ce��͸ҁ�ܺ����iA���N����uײ���7��\�\q�E�qp˲�c�W[��U�:��ci3�[]Tn�s~����������)f��� F�eש��m>9��EDN��M[.��캠�涩!�<:��
_��U��7���h��<�;.�{q��|�ޘw�����~��ˉ������n�y�����=��_L�C�]ܨn�}�w�|m�ve�$�;
����R�C�忘�S�ף��A�/�O/�~S7J��+��i
��j��Ǘ���wC�L�p��į2�Gu .�x���`��q�m�n��'��y�6�	���U;����>n���g+j�ar�Y�^���D2x���y֔z���ż�*�-U�-�vi�k��������o��:���=��'�C�;v�\<����On�ڰrdݮ_�����(�j CL{��t&�i�jZnaR������u��@y_>[#���Î���粩��m$v3pX<32�g��5᩶�A�S�io׻��q��P��s�B3���}̨���ԁkST��D:�Έ����M~���r�"�ye�ڢ̭�T��ٶ� �l�qt���gxf����C���X�7�u�"�����J7��N9����"U�n�'w�NТ�CD4���)�׷UQ=[ػ)=��艔k��};���}��us]�O�m>ͩ�uU�+1N5�~��ey��m_�X�����{\����<����\�e��u����^_���dhS�b�e��\N�&]z��dtE���i�Ѹ�M��ҝ���6{ ��J�y�k`�x
�V�����[���5�����,�{Go�ϗ��G>���<��<�W\�u[e�ö��4� ގ9sO���ɯ.)ڮ����{;�����m�㦶���7Da�=��l+���㔂;�p��[L��b�๸CE�;�����R������]6��s͋�(=�.v���.�Լ� �M9ٰI��[cMb�&�"�f:��^(�f�fA�Z�:��j��m��RB��o_\�^�t���(B7�1���l6�I�Դ��՟\���dc�)���HB�z�����#H�K�a_�^�x�fl�ND���ꆦ����κ�<ŐA|���Mt´�VK�������Z)C��:"��q=,�L2<44�<��UH���+�ܻ��⹅z׭)t���gxf����C�V��v�(}t�D���}�S����#��%�x��zns���@�"Bh�d��[Jk�p�&�n[�v�'#���i�v�����/י�U��V6T��F�]UG����������&�Q�s�W6L������Ux�}�p�4I-:��UΦbwxo��a_s_�b��Sq�pY��ki���ډ擾*�c�;EޟC�;DU&}7�ľ�Oϝ�,�qU�J����Uf�5T�6���w[o&��]������4 ��UH#s�$<UB��y��t�d�ċ}��xxw���<A'LeU +θ�@��ٓm�u�ҁ �۪�nuĂ���V��C�@�H��$)���_ nj�wu;�UqS��!>��Q����
x��,+Z������j��ٰJ:��ʪ�ٷ �Ƭ��I�ڏt��sI#ڈu��Z�wuڛ3ό ��B��n鄬n�(�}�%g�X����CB!����[Txv�O��㱫E7#<g[��κ�j�H��u3W>J�6�9�6T��eD������U��j�f�H ���l�����6�.h���:�lÆ�iI������}!���@�f�nޗ|���I�U˾���5A����Y�;�z���oO:J��RK}�#�9�m��oW:N���rm�k�鼥k��*�6�4���ڝ�%m�o(�ceˈ��j�h�hM4D�2��bf��'o��o�"��y @�k���-컭�듺�z]���K�L��p�4����K7*}�s6As1@�{bDm��C��q��޹����a;����CK@�G�g	^�n��u�85puX�m�O�];�s}��?z`�&�D<.��
P#y���x�*�A����F!�N��!O��m��44���̹D�pv��������]�v\h]���|{*�ƫ�nzS����q@N��.��4C""|v��:����足%eGK�옋@�Z�l��������#_E�?�x���;=w�f�IV�?��8+��`���.��2���Oֻ��{x�F7�G���
�V�J�W3)7G^,���Ma-��&ڇkx9Y�ޕWкHfm#BZ�tǙ�T)�}����8��N�~�@+θ\�.��6_'��Ҁ=]�uH�g\I�t���lr�6��E>�6����l<j�.��L Ph�Ix�oV��>D�F�BI�7�J��R���;F����#��'ųd>�<�,��R�P,���H<����<
�|�~��;@e�Ɍ��f������<vu �ؚΜ��:������gO�؈�6��Hݷ T�u��e�u|>�g����u�;:�P�-���l�m���ҵV؟3zej����m^����yE��;e6�m,@��6��l�h�C�t�"W3�` .�n|����9�bvP%Q=2!�q(�o����IO���$���!!I��B��$ I?���$�����$��	!I��$�	'����	'��$�	'�BB��BB��B��$ I;�BB���BB��y!!I�`$�	'�䄄	'�$��	'� �$�$ I?�����)��݂�}/�9,����������0쏏��@(I �T 
 � �(��AA PE*� UJ"�

(� 9Ф*@�$R�*��E   B�A P �!U(

�@���$P�R�@�
H
�T"��R*���QU(�H���*AJ)@(  T�Q�5@�D"�T��BAP
}�U*�j)V��*�&�ʢV�,:�wnIT��R�k*$WF�B��.Ue��*��a�O���I�O�QTy�*�p�⪻�H��wt�kJ�K6�U�I8�]j�R�mBIf�EYj�T�@}�ʠ� UT(�PP��I]h�5w�:�Z4�s���.�wr�]�ҽ����ۓ@K���z��`t�B��Os������C��� .�P�S��=��t]���{���R�ý�^�)K�Џm��PID�����A"�T�UE��7aȪ�c�{ =�Ѡ���z;��0<�v:(4��u*�:+�:��ҪI �� c��R������(wAU֥@ݸ��݁�u����@X�  ��)
�EB��  8tP��� �RRT**�T��J��: ��>���<������X��  w��/ ��� � ��{ ������>�直/����{����*���  ��� ��̀ ���(x�+�JhJGZUւ�\8 6���th������  ���'�
�UR��" U |}
��QSwu}2�&���@�J, �⤷`d�å�*��Ҋݝ � Q��@��w������R�0: u�uR���H�ݺ�9�)��SuUC���[��B��**݀�{�     T�"b�IQ�	� &&	�B)��J�  ��b?L���JF�dd`�  C�EJa)E#	�#  	�`&�L�$� 4   �  HSF���	�L��OQ=mOM#F	���R}�o����1�~ߵE�2����v�#�&f��I�"0���BI��1ABI!$$h  !`A_��7��'�������ǟ�l�����0�Ɍzcm�8�������l�;�;;H�I Zb>թ;X��i�������M��@���r�50�@�����,/���އ�?Á�P�bl�|�����>u��z����t�C3<edN��iЏ�L��QÙ��j�͘�a!(��k�7?�X���e)h��_aF���쥢]��62^su����%�d�˪{�N,[�U�wzjh���e3
n���5�3-*/5����#Xv+���؝V�3M�NL�Lwy�%׀5[N���R�Դj�T�ɰm]�R�t%4j��q�2*(�����hm��Z�˩2�n&5�t�]ԴQX��lc�����|��!�F*m����[�A�m;�6�wt�%�V��m�4��0Tj��3-�,J�1a��a5F�hP�b�Y�Q�^-$�`��q��`�0�ra�w5Q9wv��d�P�����A$T��fnۧLjJEU��W�I��4�P
s�ʵi�7�KJ��eMso&4kh|���X�"I��Y
�E�����[v�pGD\1�l�Yx��0r-�wZU�،Dm4[-mKl��o��7_�]^7 1�&��wP��1�� ńA�S���+d��B���R�G5�qUʰi�J��mطv�MA����v�JK��QYy"�a��:%@B!�C3T�2NʳP�{cv���*=8��ݲ0��Ds)6�<%e"��!(�X�R�}v��wtA��[%*V6j��b�Т�@�{g*w21[�<��-i[)�m�x-��O�<�A��y�e7��	�����:Z>;��#j�*�Gw#���d�1�	�{c"Ef}x"X����T�R��F(ߓP]����*���,%^a��%���^UF�j�K�V+&y��6>{t��l,mjw�P9@����5e�xޛX]�ƣE�*I���pLFN�ӰU����MYW����I;���]n<�emoҕ�/v�=�0))Yǯ�WB�9,-T*f<ג��X*ș
hC���W�$6� ��ɠ��6�X��7m-zѰ���#u4���ړfj�Ub��kE-[���f��<@�f�9cL;[�-�e0�ݵ[�s:����-Nj�����ͪ;��XJ�p�L�֋ME����T������"O�j��0}D}�b*�W�����E0�3�toPh�c�����n潊��h�졻�}>����Үufh��m��av*��k>�VlI�@��d�$׃ԕute7��j�59n�qg�G���5֌�l��2'M�6�ZE�;��[�]����[��l�f7�c�]�X����� [V�[�$�u��Å�md�$�R�2����hɤO�wD�2��l��]h"E<��A�4�^*�ݚ_YM܁J��y�A'r�<�pԳJ�;��n
e��z+,�u�#����e�3f��TkiΚ4��YJ�*T�(��n[љ���w*A�Q�ݦrL�!ĝ��*�x�{&��]�H�S�@�Y���K(ߛu(���0�m	�[f��x������ۓ�C0��MQ�X�Ҕ7j�B��̷ku��V^��ٵc�l㣱Z��[{�&��$k]�F���'Z�Q����>R]��R�i9t^ᣀ�j0��ABͼ�7*��J��YY��˦I�k~Wt���Al��j(Sכ��hmm�q�@�8��d��Ez�f���`���L��X��حL!���������*=�m��W�t[Ȇ�L�N��#Q̫Wkp�R�m��Z��82n"r�B<E=��(	�X����J�mQ���u�Q����q#w3pJf�t����h�{&��ۼaK�.�V1�,��qY&kV���nG��CV2��*i��62�Z�B��k�P'�*AnU��Q�X���SJ��A�,*���h��f�ŉV�+g&ޒ5h�7-0F8*R��Y�Ekp8�`�;�f�a	�*�$튭̈+��f&i��7B;x%_���z�e���Gj7r�,�:\X�ѳ���Nd��U��c40��i1�{����0nMv�J���E�xb��&J���m,ÕyL=s2���f����v���C�b�V�f�3���f��OsW5fe^I��
�:�op'��Ӓ��ڰ���a�e�e�h˕�c���l*�V����:(�ԋAI*A4�ͣ�6��{����v��p�`b{b��Y��� ��EeA���)��JTw��X�0fn�VBuf4�@��bV��L���3N�z�e��Y�Bk�[3��m04=֞��������e�L˚�˕.����;OM��g�D�Q�� Y�d��y$☁�+�}��Q?b�;�̫�ǐf�
�n�u��7��$�b"2x��P)�3xp<�6j��b2�x&:�0�[vv�E&�۟c�y���f�[�]�!�(|���A������u���\Q�dc�"���v��^jV�%�}�&tת�m�o�l�XFQ*�
�/�7�Q3hˎ��V��C���R��`^�w��GhTU�b�8b3Z��*�-�rڽV����?;-�y�Q���X�^�6�R���6[�0��r�{��Y'H�$l�t^�T��,�6�.4�7K��a�[ �x���<K-[ʃ2z[̕�O�����;�ֲu�Y�3y�i3�F���;�m��BBd�%�]�ܛ��n��*�-f�ۺa�U��R�ړ,n5c�m�y��_#��+�����+j�B)&�J��<;Yyla�oYٛ�ēX��|`��n�I�]ьջ��@ck%[�X�V� *n�����ϽF�Zi�`���ad��m�&1z�WH�U�	��Q'm--�G�1N�<;-v�YǏUCp��2�70�,��Jˠ6�eҳw�����4#(��ܢU�D�:��:P6b�$�h51�l*�M�v��Ù���Xdܸp�B��9���v=s�
ڵ�I3p�Pn���^�X6m�˼��c:�k;����-�B52�rd"5����J̚s^��o�e�2:�#���]2�0F�X���k#�j]*�6Ys0}�V��w>7sq��gv��l9{���ے��R�le%�������x��%�Hj~����fPs&�a��f��0.iX�fM�eiUy,ە�.���0b[viE)�CV��-�-��v3�M�ޔ
#ci���(��K6l�,z��Kc��v.�u��{[v��7�َ�\��w��J6�9�!�eDW����Pf�A��\Y6)����+Un]6.m��@ʳ��CJH���^ؑV��D��KV�x��z��(��$����Y�����IQ���!�b $@���AYsNdtu]�N����A�j�g���hI��MoZ�U��`� ^k$�M��k8��S��\ ��w.��B<s��`�i�~�K��k�׃զխL��s~4��%̹�u/l��༩���P���-�y�U�)�٭s�n�z���fV����u.Rk&�	ͺIʼ#-���6�dl��6X��J�+dU���N�似�bfI`��/޹o,�.�0��(c�c,9i�&<��eU�,{<���LW�>u�nz��xdp�b��Sv���S[�أ-}7x�+6���q��7f0P��GN&Q��cܲt
�VpVA�^��y��Q���+&�0���([�P�$�n����-7��������(ܳ�����щf���{�+b�U��n�\S)si�"����Xj]-�f��H�/P��n�ɢ�h�K� MP���f�NJڒE��nü1R���(7b�T��.L�`VX"�)��qC��F���T�.9��Eyb�Ě�5c)k�d�n��н�6�%���QE�p
 k�a2�CTxFMڌEtE ��w~�@�v��s.�j^,U��&G�V�:�@�����a(p�R�պފ�1�6����)v�ssv�b:��L	c"4d�K�f�����8*
T�Vd(�6�͊,�Ƿ�{�Ѹ+n�킵n��7F�%�*���U��;���U+m봮����dSɘv�J�L�[6n`x1��oJx��Ӄlma�v� �Fh�E<)����ef�	]�r�[�4�[Q��4��O[�9�FCkc�/d�r�J02MWX
��T�L�͏S~�Ry���Z$�1���F��e�z��E���#M�06i�i3~Aş\;ZP��U����k4e<�xpL�b�(/q��r��ä#����Bɯz���m��l3Vf/���/v�E�B�0Vh�_�!�[������6v�r�C��4���XN
�k]Լ���"�@ܖ%�ft�z���YM^��H�P�܂�&����@��Z�7%���a�i��{3nL��H�x\��p�v�(�Ԣ�m��b��<���uV�3&m������vCJ�:7n��˩Bv�C���oVk��
	��-��ˎ���S�b�yD�1�1M�K��݌� YN�,�;��ٞ�<єD�pd���Ǩ�f��L�c��@�)AfP�˸*E�{���2���-�׏q����m7�Ew�a��j��Fm+(���L�����Y�y���Q�:����'{�dn�Z�ː䅰��w&ں�OJ�� \n�%��5%� �4%J���7kHŹ�qXb�Űj�r�9
�ڃb�e �')P�+���ڽP�;�e�.(�^���1��f�[)LwW:r�����
���r��;�E�u$7�3!�w��-�sc�m��KrѬ�4�B&��R��F�/C�L�+��"^\�.��3ج۬�G3S)�Em�|�����5>r�0�B�CX|)�������1a�n�n���.]-nfej��W�/�s�]3!�-�EZA<�*4�,f�6t���N�a�����m�F���y�h�ytv��ZJL"�1��7pUE���RG���m:��W�]쫘����q�[Xv��ЈdP�"h3�vhޤsb;!/3�1�[2���(
�3D�gE��9tF޲[:ǉ�y�(WZd.��cX;��e�D�^���i+�biFd�V���A��T������_�Sؑ�V�]���U��aԜ�����Lf�&f�G �s0�mIf� ��X̓%aF�Ñe���U���@�ɕ��9Y�;���X�B!�{�2�R����t�z%�5c؃�Q�3P�C�����<7/7�*d⦳E�Z�ue�����˽�,�dYXrz���8���X܍ӿL� �Qcq��Y����V�D��W���(ұ[.��-)�5
tQ�N `ۢlF.�Tu�i�[�j�B)4lҬ�su4�[j3k.������T���d1�=�0i���8�h��j�f�sjY�G�]��%@����2�Kz���G�v��4�C�+h{�[��]�I#,�;�u��F��`����Ǒؗ[��D��*����,�UfUƪU;.S��TbY%߃f�5�Y�b�ZA.��G5Zy�I��D���TPn�mKݖ�n��x��wiV��n�`��{�Ea^�j�Ӹ��U.f,Y�֊�K�Y���ےk�߈ef�q���fV:�{R�� ��ո���
�̜8��n���p��ޙH�P5���
NH�dۚ^a�)]9v^���2�g4L�5=]���\A�A�B�#%��ղ`On������͂ײ�c ��$$�q�A�u�ԉ��",�@�{��N�8����]��ڢ����Iz�h&V�Ph�Zc��B�UՃQ���A �ktF�X��)P;F�l\��sT�WJ^^fU�Ҏ��@u���Cb��D%+OY�U[)��ֽ��蕛�];�CX�ۻn�NX��Bҥ�ĩ�k%Lx�w"nY���bRţn���,`�A���~��O1���_�uf�K�7��͍ۚ��IZ���?����8��4|��zY4�&���#�,c�lbeȏ�j�d�j|ϙ�(��#�`����! n Sc�Ɠq�i���( c`��av  \c�`�`�la@�`2��q�
m��m����ll� �m��v0�*�@Pv�Sl��NSӶ�� l(Hm��2��82���bp��1�ˍ��M�� (e1���lli�.���0(l� �llHm�P���e6�LӰq�Sm���cH(]��S�N�$�.�&���� `���'m�&pN$؄�O������WO�Տ�����Ls��I	$
y�q��$����/�y��p�?A*��@�a�Ƹk�cr�ç^��ǈ��V< ��$�y���(�Z:+�A�.�P��=���S�#F��Kk��6#��r���ӛ4MX��N�������4��:�^����y΅�o�����fr�6��S����V��4��,+
t�����qU��;!���>�\h�m`	�GU]e��1z=���A�^{r�	�:V^�O.�lI�E�H����R�����rж^^�e�Z7Xplm�1a��#��p:�k̚�����5������b�8}����7[��K�sW�����Mt񑮌��q�7T=G���3�<��r��M�n�%�+Ͱ�/�-wY�1�:;wj�h���h�z�*���p5������s�r��n���否x�3��֗�%e�YX�e�W��kv7|Ջ�K2�X����p\NT4��|9�a���.)����YJ
���im��L�\�*�c��6���1�yS]�w�������3e�b�-+Yͫ�4�T�9�5gw+[�I&�\�ι�O���
E���v�osսQ�M-ᛖ����٦]�
\;KwY���py��ʰҼS0\�ø�k��c��Yz+U����ZV�M�d�ʢX�Xx���-d,��d�5q1�ZK��j�c�W';sz��4UۥLCv���;��ٚ𪌪��&K��i�p�B^j�{q��a�8��xvA���Qu�:���^�V<C���mmo�R�m\���3g/\��𗓥(�9��f[����d8���7����)��#0q�s&X�ϓ���pi�)v*�]�ə�ܧwf��M�3H��Vk~:s)���,C�Rᕄ�i��4%3�L�ठ�Vuqj��Y,+��ʄK�D<�]rF7�r�h3��p1��!e�tf�؉�#�f�MX]�&�f6��$Þ�a��-񎍈1!YKm�z��һ["t��,s-�Q����;�ngk�ϳ9�rݝqvuX�}1�R{a�Cl��wvI�n���5r���߭̷!L�m2=��`�V~�C������=��z�R�`��^щ���P��S"Y�JJ�Ff�9e�a�8�y�b�]�z�S8U���k$s0l���\�˕��:�a�x5#�cן:���qV��J��q�~T4��k�B����붲��5��`Բ��˺
�6�����S�7޲'�`���D�C����um!�p����^eM����P����&L����7��T�o&I���~�N��I�:N��/rm�e
�̈́�=vr�Q����fa�[���� �޵q��nj,=/J�9����4ݚ�F(�Ak�2[��Һfc^J�9XU����lG������;`�G������͘7
�7��丯`^r-m�$�=t�Y���~�`ߘ�e�M����dr:٪�'\ϙÎ�b�,YV�6�U�j��z�ծ{�����Ε6�M�gvs(̓�jc��;��Y�R�+M�O��	��:��.�ߝkk#�6���,����f�7^����!��~�����Ǟ��,@�����
ȉk�]8��P��b�h�	ݹ�,$]�AX��Z��tt(��B�dnŜ�Oq\�wsv`���E�z�Vj̚Ѹ�!*j��ݝ�72��,�hަ�wDp�QY�ot��,�L�Z�괁���줨/Q�@1���V*՗�jL8���=a�U|����-�
\�v��A�a �Gu���������udBV�SdlY�&a�����[J���eq�\{h�}l�40��c<p��&�]���ӓ �p(y���WM7����8�>%��4e�/fñ�*��ܶ��D٫V��������z�픹�{Un���"á�Ӧ����R��d;�yWkS�����eL9�|)�[3NY��BeI���0�����ױ�цTۊ��&�A�җ��p�ݺ8�nC9�V��.��E�\�݇�K`���R���˥�)�e1q!p�z6,q+�� cb��u�ٹ;5�Q��3��C�r]֊߲\�ǆ�iCY�J�**��r�����P��x�,ˣ#˸�Z�&�/�b�A�k��eJ�X�͌�y�3�=z��-hD�f�	��`o
{�l=C��0n� ���qd���Z�b�i��e��\���Z]м�[A���/��t
+�l�:���JV���X�����_g{52�,��P8�vw5[�ޱ&�WD>�i�˴xA�P�w�r��mL%����j��1����9�Ek:��<3]d�j]չ�o`�m� <M�[���%;`����o�F�N�/��ِ��pȩ2U�3r�a�4�2�P��ؼ�E`fp���O�I������c��}���/����S7�^\��@�o����Ȅ�*�Vk��ڽm޴���v�8c#"�\�+W:v�G^�/9JI=E�j�4�8<M�`�U�6@WVVB��|u��s�k��W�g�Y�� }A��γv����<qiS!@�84��;�g�+��Ů�s�k��u���E��t���7l�ʁz
)�R�����^�*8��d�KlH�R�5����1s#l�1�u<��C�-�P�
ݛ���V�[ާ-9Ɠ'��m]r�QK�	E5��4��i��Uꦰ���*f�Fl�3Y̴3���Ѯͭ���JAo)�]��ޅȵ_S��qW��Ω�Zqjzn�7OU-v�x����}#��1N·��5}:��9ʠ�b�e��V���z8�ї1Z�,�U�J ����f+��zm׳)�NhÖ\�Z,��B�ك��y[����ڎK���]Kz���Mg�;�rb.E�ܞ���ř2��Lu�!�T��5��[�sjٗQ�n�u�uy�؎E뼙���qJy����U�JWsSy5@m�Q`��{j���k��#Q�|79J n4]	�N��pU�i��S�jd/P���;��h��\�*���:wQ�I��M�`����=*nФ�DM������xv�%1GA��U�Y��\͂L�'�:�Y�4�]
hs�ʷ��d��Ձx���[���嗒��S[KyT]�LY�U���h�7�E�� �g]��.���2P�&��N辝�Ѐ��ط�D�����
ؘt ��[��P��7譍�'͹sM�?{Vb�ve��^�W��+�˧�\���d��n�2�o<���n�c@�^K"!���/N=��]�|�#��ZH!���S��ܮ�rʌ�dۏ'kݮn�=v+�,��F9M76d�K�9_�r<O��/PfU����s�����JZ�Z(�UK�1��9�d6YǴ&3��JY�eE�ǐ����ͺڗ��m��sa����:n��ޑR		�)���TGVc��5};s<v+�/˂�;{ pc�XH��u�:�Dn����TՅf�W���3�P�6��N�Qm۹Z�,�N�n>���@'�N[ע�M`E�Z�����qܽ#,Q��ܱ���}F�7}��2Ջ�Y�آV9���l���뵼:��A�F�+�&��
z��:ƚuX���2�9tk_��^�X�$�	�PI���T��=�{-nc�i�"4�ګgj�g!w91a.��Į����y}f�
�F�;A��������-��Z�gQ�����u�x���-��˶�cKG5/7�|J�,���rL��
��՞�j%��}c�e�c�.鳙�y@�[OKN`u�&�cx�z�N�o%�b	������n�1FL7C���IS*���7jM�	�]�ofj��rs�k��ηGA��``W����כqps})W]�8	ЯgC�gn�4�Vȣ�u&�2[�Ƶ�H;�J�������f,W0�U�����y�8����(vTwl�䤁��h#�L�s���7܁=�U�G5�6h�tnd;�Ɔ	2�R�����'�[
Q�mwq][��$�(�Tn	G�:��*��mw
��e7�dLj��@M�BF��W`GE�_p�;���.J��K�C]�5��En�b�0:f�7\�_Ө�!��Y����ҋo�rn��3P�E׫M�#ҡ�Ib�o^+u��Zd$P���ˉ�����W \��~v��7[жM�������Ҭ�.��ɟ"ʩZs�uw���sS��OC��%&��3ՒT�2o:o0��Z� m�ɋ/��׆3��i0�@�{r�:h������<�ɮ��И����F�a;��}p�~�{-��c�E��Г��Jlޫz�q�M�������w���Y��v��tS��#vd�e�Z����U�>Ʌmn#z7c������xM^^�rK�s����&{2�p'�(��clUM�z+ތ�b�ɜ����l���bu�Uu��{`!�cF�Ϛ !��C�SVn�;6�Xy����F�+�ek>�.�"���/�E��"m���]w��^�έ�M�M2�����K*yX�ܼ�k%fe��*�<��)NW�D<tK�rGR*�]v��Y�t��S&İ3�yZ?\|`|������6ǻ�}�g�A�ҳP��2�d_d.��:3����PF�L*��nn����F�b*�������U�P����^V��,�h5q�}�]�/��1ϻ�٘:u�7�� R�(A���l
И�%�v%�X+\b��$�.�Y��8zne�8�H��e�fmC��EvRO�+f�%��x*	t�@7i�n'���I�'���~����Ӌ|����gݐ�Dݢ�u�*��' 3X�maM��9<�
dB�t�h�Κt����fn�Ŕ�<*D�ׁ۴*C�۫��U��[�(�%��m��W���T�fH�^(1�i��\��#-�0��D5&���i�ۆ8�����-٤g��3��(�6�bw=��B�dp�Y���S�ɸ�_P��ǧ"Z�g7V�#�=O��J��d`u��T�fU�]ǻ���u�h��-cX/N��	4���C���[�7�Sz�%��l鼸s3f��XԷ��`T;vgu-sz�9۲j�f�tj�&�`��֐p��+��Fӛ�e�~Y=���C]oS2]W�h�乂���������2Yd��:
�!���a�k�|����4y�̙�u>���L��f߆Z{Y7嗭����x��wFT��+6�ݕ{t�7\Ӡ��n�{wH�M�æ�����dUZ���(�W��zlp	�q�a��^��~9Tq۷U����L�h@�o��E��Szl<ݳiy�֡T���v�lL�"�U+VU�v�>Vﾱ�a�w2� p]���O���^�-	����D�E�b��i,b���m2��WX��wG�������.����	�F:[������;��5eTR�ܱ��"3��b;��|��\�����d��pv�jΘ��k,����:{H�N}q���
�� ��M� ���4�7��,�V�h�U�}�}j��E9�/>����ud޼��4<���H�6�B M9s��|��@*3�.�"��+����)��nj�D��kGI"���պ����L�vwr8�-�q�t�\;7:�t��8��C�GZ-o���Y!`���$p��\���e��<.V޻�7�pv�gc��lQCkoju�8U�;�J�1yf�y����!dXOQe^�RX�US�͌a�S��ll�w��zע��{�Q�K32J3.S4ܾ���*�]S.�ՙ��[C��;�4Ji���R���X�궅��2ɲ�&0�]�`�A#�n��OV�P�7��L�R���!�t�фf�;>QJ�-�B��$A�3����n�Smc.!)n��`�I�������פ�mR;��v��o}�Ļ���XոJwc:7��q��gJ{�3%d;<�6��]W[�OqЬ�Vz��/tmH-�������I�1��1�*��F3[7�9�� BI`��6���	i� �4<����`Ph1?����7f���b�Ρ����u-��v�I�v[KX){g\�]<a,��L5�;z+�����qݞB�:�ƄË�7i+\�5.L���dv�p�nk�m�]����&�9w'S��ٽ�'�spZm�,�6���U�zz�s��h�Lj �6�r��c���qu4]�	�pl�۲'Et�Q��g����{9��pqx톖��-�]���xVŃ�T��z{�ۮ�H�$����7Q�!�1��:qɳ��׵��g! �:�#ͺ͇
���'�]��sS�W���\�מ���4f���n�:�,X��ӚH�թ���U�Y�4sr8��1��z���{Z;z�Ѷ�vyv�NQ� |�<�{��e�-��e��a���Va�r�#�'s��>���a���.�ї���2�5�4&�Ō���e&�и]i[��rp��vс�y�J�'dE;c��Wt�����'/ku�]�x����ӂ*7mBNq�/��}��s˫�^܁��[��P�9�=f��8�Ԅ����:�8�j���X��2�N�6D�_j61�X�[�Oc��$�+J�'�� Sv�lKP����M�7�(��eô���U�.բ�v�����u�ƪͮ���&%�/�`�.p��yZ簳S�ٹ���X|�β
��Z�z�-.��\q�K{v]l���tq�f�K���z���^� ��O!�z�4��.hd�C/+V�.����)����ڸ�l�˅�qa4s�e����$+f�d��2)AH�ѤVYG)�%��2�3Q���!�6w&ɮT�t�jKN�����ˮ��Ύ�rc[gAa6������mq�B���I�v7WI��1G8n�`��M�(��F�]^�Ŷ� �MՇ�[�q��w`s�^�֗�vMݷ5ֱ9kd9r��2�nx���e��.3�;C�;u��h��ƣ/7mR��q���D���)i��Y5b��k��H����]w4v�o�\V���Άn��4�ŔT�ա,���/`���j� �`�+nzy���vny:�-����ri}<��S�z8Ʌ��x�x��۞���ˠC@BX��Wi��Й�nc+��t���6�<ir#Z11����������gK�nĖ��=���c�{(���`�7:��^�q��%�,�T��ء�}P�؀w[��n��[�T�p<�.�J�T�zۨ�M��rf�^��d�^���si���浧k�;����HXY�����5��X�zbv�6:���;VM��L����v�©윉�D��i�������]��똀�Y�{lW=���ܖ�n��!���X�S�`�tZ�8Dyݣ���Ϟ��箎�#\[9���z�������s��ۮ�[@�Cse�.:����Y���`�Ss��a�fAê�*�(��ŖD�:6�M4B�I��y2�䧮v솆7K/RVG \��ae��Z����cb·�#!.㵖K��V�+�i����v1ƪ��۱Cs7u��j^ܚJAl]a&�f�%�����"\3Ua��ȑ�XR��mF���n�.ojMz6�P%)���-�2��WK�&t��Lh[e�7\�B�s�[��]v^�=�M��[�^�5n����-c��s��i��q<�zh^( �k�nH��>Ȼ:�K�j�6+Q�Ms��hX���;u�k�zx�vعtt���}C��՞]u���{��hٍZ�y��ω�u�Z;m�v]�T\pܚ��Nq�K�[��-�AY����4i��z�GC�+�Sӵ\`:���h����M���3�z�����yl���w#���/��agq���v�n���L.���-��B!ۈ�=�v�'���Y1�jƓT����u��oHK�f�p+Ij[q�՚t�f9����^B˵X�Еy�����q	���t���ی�]Z����m�y:Ue�Zv�ԑ� ��Z���c\��]sѣ�&���s�8��:���s�6e��{��Cܥ����ӖכoS׶*���&lI�{/7[ϣ� �=Z���t뇳nB�R��Ood(�lD�77�j��\��[u�Ok�kAsa�Q�r���F�h>5z��Y\�9Ӷ���B�s�L�\V�-N�J�ݲ�Fn^v���n�ɱGhVv��mu=lʎ�]v58�<nɩ:0Cڒ|7j�]+���7*��4Yl".�62��n�[��b��F��j�ùT���V�g�֮�M��r�����Zb.����KV���i���aMr�r�@�bX]��Rj��s��p�o^�wn���Q�;&1K��P�#Kmr�RY�#��y���W8 �7h�]��FX��t+v�˃��Lr���r��M���[v9�Y]�5xZ�M<^�r��3]pK��:k|BNrV�r��Ɍ�Mɧ�AN�㧛��vGWe�t����m�v�,�.z
v��'Oi���-�����88������v)��;g�b��u�_I��,m�n�e`�2�Λ�%���ke�Y������C3����:5q�������J��e@�[Η��,v��2s����T�U��N�>��nv��r���f��f���%ǵ���ř�k�\dcu�C�8��x���۲�1�L�]=���ǋ�=����p=�FCY�{��OGnW�Z�͋x�j�Et�tyh�cb^8ky�	s�s��iI��Մy�̱�slM5�B(�]���ai�J�苜u�A�;�d�:_:y��=��n�e�I[$^��E��Kƈ//<�fG�����m-0җ�iPV�,�t�n��z�'f�����oe7ܴ]M��^�D�4,�q�N5���ɣN]�B6�e��CKt��a�K�ƞä3��k7:n�]��K��]��5����+�u�<ƷJ�*�UpB�Y��[�����v`t���qm\�,�$����nΝ��Y['\w!Vns�G�%x�a�� nvw�c��q�6�E(��Qec��B�K�m�m�m�Y�馱YcKv�FK���lO=�j�s	��꼈1��U�Ɉ�8�,u�����:P�h9�cTg�	d��^�Ʈ����H����\D���:��c�iN٬�+Ja��1�m4!6����b��R�چ�4��a�K/��v��"���F�X��(�<�6����P������w:�3�v-\M����`�z->0	E��;v���d�jvu����fS#/.�Y�����:q�i2�#u��/�^�s�q���ЗV���6(�l�+�ͬv�J��pc�p2��T�z�{<��-	b`|�|���ݳ5��ns�j@��6�Ǧ��cL��,r�Z�4�nQ����Vw�nl�Iص�q[�.x���e��:iY����	;Y�[q  P��y�������U���]���d��5�TQ���)���=.���	Ы���k�1��#�D\��3v����U�x���.��+�)�89-0
�Nz��9���t+-۳�F��س�F�ܽ�W�l��Y��IH8��J��"�TT���X��'GC��%���@tP&T����(�s��Q� ������s/F֋��Dm"u�s��]�S�Ud�z���/X��Dd��9E6� +.�-�Is��;k��\P�k�u�`�v]p�W[Z^8��+B�n_n�Q����W���$�H7.�Ѻ��g\�֝�\�+uP��vw+�*�>�5�z��\���r���mv��r�n�I=s$�mldh��Ks{t[\t��p�����6��/n����k��kf�낍s�I�rb�7�ll������]-��3H�T�:�i�j���d��,5U*�UT4ٝ���3Fj2ݝ���r��fKd�uר��Ӗ�%κqd��N�Gk�9���m��Ϭ��:��}�¼�u��݃�:���Hv�x	����V�ƳJ���lr�����a+r%�'�H�aXm�m�b ��e��Κ���91=t�8�� $㨩��sc;�\\6� LQ��0��-=\4c�n��H�&�3�e�cm�1�ґ�ӌc��ȵ�6ѱ���.m��+Gz�#����y{uہ��nen��<�im�Yy�����t�<��\b����.G��a�l��W��dR�0�M(�k��ߎ8�p���G����*��"�#�W���9���TL�����AL�ZQȹ���EˑG��9EEQU|����<(��*i,�*�:�O<9Ñ��J|#M��� �e�I*/4�\���r(�^P� �[^x�'0�Ѐ� Ut�E0���;�E�˔r��/]�e%\��
��E�VDq���C"*�H�E�y��;�W��2Y*U"
���W�y�D�U�$\�Ux�\*(�$�SC�$�p�R)�'.U�D��Y��ӝ�,X\�Q�E��N�Qmb4� q!����Q�9
�s���VD&g𠨳�Q�H�[Z�tBs>wI����y��.²�Ui���q��=ae&��S
e!.ʰ�o>�z29mv������Y���lvd���VA,�ܝ��5�e,�e�[ݫ�Za�b�p٥��2��u�
����q�R�顢����Z�X2a%Ŏ�S4��l��Z熸�k���:��6/�N6��ny}�S�����.F8����6|�`y�bC���؎[-6]f��bJ9�-�#��b�C.܃4���42��Q�
�[lsI�s������ڼ�g��5��p2KDF�Ό�.�#5��|�|ݷ|]���u����jf�JU�ưҢ�#e)�u&��@@��i����`��:.�֏��yC�BU _ƈ�q.�@Y�3�GeUE�e_n��<��B۴f��v���V��9��x�Iv�u���_*��'�D9�[�w��[������kv`I�˭mt�vPk�ie�l#,e��&`�eΣ����[s
ǫ����{F���KЧ%���n4�S[�^��q\F���؎�j�W5�S�){h�E��\7���Oh^u��@&Q�S��jx���;�l�&A)1����nR��C�/�x��=�x� ��c-�YH^f46 �@�σ��l�u/[�������:���uukJ�[yD����5�Sa����-mh��ێ�M��r�<U�m(����G#�j�Yl�%4fcզűm���ָF�]K�VtʛfN��3�S �,pv���V���s�盞�9��.s��BN``���v�TM-���Ƌ��Eݮ��-Խ�9�6���s�I�mu�- qe*m��8籧F�;�g]R�ն5�l��wi��T����j�`*Ԕid��)IB2�)-�N�DXKm���A�D,���ė�H-��!Ye�,�b,Ee �b�����b�c������0�#k*��#	m�h��z��k�#e�y󇲯��r�TP�/Z����45 �K[¥V֍���1�25m�������6����������RX�|�	$�5�İT�X��T[�� �&���W+�뀠�hFm�O
I+�^��6������z(���]���&�!�,Q4�5u��3��U�`d�l�a���S�TQ$�Q{&�4KGo(A��'�h����I�o��5��QI������^�[��3��.glK��(�I4=�I4{��SU��ĳ}��h��5I���a�ۈ�nЛ�B�I�{Se{����D�^��D�Ow����C�=�Wx��K[)A��/��:y�^1��M�I�h�#?!
a���,hf(�q5�J��*I ���D��˻	vG��Olm��f�4)�=ީ_$��Ɉ�$Q���OWUe����y?��������x<��M�Cv�;�W��x̮�K\��n�TV��#UG��6M��]�sT��uV1f嵾�� ���� ��kl�J�F�x���P��n�{0G.�e�Evf`��g�Sd�I���Z�c^�4�Geɟ$�I�޻���%�f�L�W:��=+�#=�I���b�MQ'�vz$��'��4�z�mX �=�R�K��d$X.|]ڛyv-�޿"�l}~�Ș�I�,D�I�tm��H��Vm�J�?�f4]�g��h�/@�>%ܩ��\<a�f�;�y�ˣB]�n����g�F�����) �Kw�Wi��/�'���g��H�w���D�7ѿ�&(,`�D�b&���}J��������f	�]$�Iwo��$I�|k�D�I�#����-w�BS�ꉕ"��$�am��� �:�U�E�{��Ɵ���1S�v2my6Px�9��wL�뮞�T���[[�����AI��R�����ʩ0]`�.?eӋh��=+7ݘ�$����]�E$�[��R[O��R*2�fա6��b�\&��ꍄ�K��Ʃ$��u���$�D�Nʱi
�2X��P�uiN~�K��!����Ճ!��j'u�o�I#޾$�F����]�ݫ��{�}	o�*
7��n	�X�k��p�s�\\g�Л��3����,>.�)׷v�DD��H���$n�V����/�ɽ\-�ri�I�^(_�#A��:����&=��������Z%�^�I/�G�*$��7jzLӞ*�r2~���Q�	���g>3A!��|�J���YЗs���ԉ_.ɦ�Q�z�$���L�#*%����z�+�[���h�|Oz��hl� �G�g9B��r�hFΪ�����p�[P���($�ܧ�~�#��W���{Y�ڼt^�^�]��ñh�;.e'��4n�v��A#���$>�z�B�Qc6�}$�D���锖gl�Oz�1h�BtX$���hr�E~d�6�]�g��z�j�y5s��p�a6�D�6���4�߯�`��9G�D� �]�0 �z6���^�Y�t}H��=��A%��d$X.|]�Օ��I�tuL�Ҽ��~$�Ib�I$���l��:tw'y����R_7ˊ�E��f��:��&��z&ɢI2��0�)bJ$�~��"����]���c�5V�s�w��`�V�	��)$�[��	 ���7��hv�Q:��R��ϔL��j������&����E+~1�-�'�O�{ѶA�I��	P�wGN&iY��>�Y6C�3J�Y��3���E�bnIo�����j娧P�����~MH{�.:�lcF�2�3�e�\�x��'��d�Wn�e����Y@!K�FҘ��=�r��n��a�A,w�B�T<�.��\�݌omY{v�>�6�ST'k��εX��u���T����㷈�4t8��4����i�]�]v3�76�m<y��E�;U���^��U��jy]I�D�ΑCa�W�噽�Wb�]1��җ���~}����������Y�$Mh�� ?�5;<'�i��5i�Cf�D�G��:d����]:�����D��̵�U}3�$�d�m� 	������Ý8��䤹mx��E����{YYh�s�TI$r�T������ �:4�D[��x�_4d��k�ueg^B��y��@k� �4I���)Q$�C�,�˭yjtI*o4�
������G��$���HA�Œo;���I$�� � ��U��
\j����$�8�����ع�6��q�{K��V���.3���ߊ�o.�̀E�y� ��UhD���X���l-V�_���I%纡����BF"�fա6��"E��2�n�4��f�"s��\�Cw0�{��P�0h秇eݢ�b�5�[��������]Ԫ�H$�K�ꔒHw�%���i��]�w&ѱY���`j�XK�E��I&��Ț$� �nz��S�����U�"��IA%�|���L'>.�g���ᢻ�=:��$�K/� �"lX�I/��z��8�h�uboبRM��B�h��2e$��-��_֎ɵU��m�ės�"MGH�h�{��z��ξ���~FL�
��\E��r�uJ�J�g��C��.�ݬ I�& ��#�0��&��T���$H�����C;�vM?6u
f.���I#�ꔒ�1%
N6��Y���wL��z��_h����$�'��`��ޫ��_�>n���Ioz���B�Xe�k9, =�k&�$ê��].h��A�ۯz`����=�ZKw=�v7MV��ꪾ��<��o4�IV������8M�Mp�vv���h�;�R�H��ޫ���K��*�ڵKu5�Q>(�~�_"I �z6�/=哞��3.��!&�3r�|���6
a9�v^VVI$��Aէ-v֦,̿�@�ʔ�Iپ���$�r�H�-k�X}�)a��P�i�-������Z�nRA��
l���
�pȘf��X ��k$�I���(�{'=}C�� TI�����4b�7 �YDa�e�Q�P�Ṛ�u��~z=�4RA"Vfz�� {�"��,����$����(R.3r�����I|���t�@$�l��y�a��׽9$����$�^{ʩ!��V��P'V�	�S̿.�J�o �%9�D�x�"I&��X�� ���9$uǮ����r����Ģg�=�\'�t�3�u�h^�J��e�ۭ��Y>�z��r�Y7�Ȣ�ij��I/���,��p]�D�=� �w�|� �="�N{ev��*A�;��ř�b&����!��B*V���]�HmsȲD'Ŧ�wqw͂�N|^�yv-/�'uI$�I_��W�[��r}}w���Kj�����\.&�:d�D��#���=��I }{�D��z��Kku��b�ʢv}y	�0�Q5X���$H���I$v;¨��ۭ	 �Z��&��II!7�
P��
&�]}w�.�4�����֥b�#}至M��y�x����P���z��T	�իBuT4>I%��Sd�?y�I��P
�4ň��&��Ѡ�`�+E֪��[_��L��X`��}4=륽[M7�QspQ}�d麌��:��_n|�F��Kygn����h.����Ѳ�)�O	��7l�uВ����U �=Pem9���w�l�v� E54 �ndU�.1%�:�M��v#�e+wl�y�wK^��s5�)����u�V5�d�u����+����VS��&�m�2�v�%���(B�4������^��\�r�-c:����T�M�:^�<�0%=�f΃�y,@a�4{�7^0;C��p��CA�p�x�c8&��$�I��F�%xK�y|��:����4MN���5���tѼ�[uG<��I,�6F���h� �,TI$���2	#���;�d�,������\L#dt�$Ooz��D��:�����$H���I.��ش}_{!�2����ݛ��4�0t�$�S{ȀI?zz6�$�/�O��U�H�$�2��$��4�*B�n0���m�I'�q�xVd�.�$���I�w�ŢJϹP�9=˵�ޥZ(�3`�Fg5���Tx�ٸ�MlBUIv�s(m��ױ�Z*�j�!6�	��U�$�<���K'+�����$?tN�4��B��E�KW�J	UoyP���w���_��ݽ��4.�)���"�Q|�ͭ����Jљl��F�1�9D���YL�3o����{��@$����I$����~&S�;o����J�z�	��N|]�Օ��	 �.�t�I,����>g�{k�ݽ�	/�Ang�Ţ�K�yCQ��B�23�������}�ڑ$�)�MI2��h�C�,��6���D��d����!A?�����wS���!��T�O:�	���Fr�5��m�H��x��k�d��J��2֋��Yv����B
��պc�pPƨ�%R`KYy�2\�l}����Y������u�h2@�ܪ��4I�b'�?gǽ�0a('��ݢ�K^r�Hwz��TE�իM����go�-7׷�̪9�D��5U������	yl�Ը��;���砳j�Ep�W^t�I$;=(̄����ikA5���W}������Ul$�8wn���o�w�L�EWe	�t�J=��*i�87&���;�5����R�״v�\��p��HwU��7EX7w�U�����N�$�r�p�7�k�o2�=3��hJK7r�8��w��C�iý�֜Yqi>�E���pg9fX]\U�@�F�`�D2�%��ɺY�#�f���{k(?Lw��b�,<�c.�u�i��SV-��ћ������Mf
�ϸlx��]X��Õ�sv�T�|�:��H@;�����C�D�Ɏ�� �.��z+�����6���ϵkw��{K;6����2�6�N�/�R�[�)��`:D����77z�4L���}3'��ͻn݌�i�7b����--K����kz��ݝ1񔮐��gw�[�A|;8Nھ�I����.�L��LǴ��鋜[�����Z�r��q����0yo�
�bI<�D�/A�e�j�I۬��q�]�1����"����9�Y�e�w�����H�8]h���麖WS!��ajb�Ϯ�`�d=���Y!�*����3��S�7����V��9�h��Z�������e�'�v�V��Q��E�/Mnf{sNb�r��9��`+�f=�,�6
�M��u��<�9f�3�V�Aǈs�����_���Q��~�>�I�xN��竘�iĥs�&IN�#��X�2�!YH؁ ���y�C�#�"s�te:�Y^8wV�'K�UN-Tu�	�4�F�"���y�I�V��D���d�	KW�F�C�7e��CL�a�өpHRэ  %)߬�D�eE�8�dY��ˊ�N�����KYB0Q8���"�D�6���x-h����%)Ltr*tR��DT��D��)$��˹VbmC�b#�5Nr�ǚ=[l�`2��Ġj3h�	�H[U�A�'��QC-!�:y釬L�iz��2:�k�G,YdG�K�z�!�w)�X����H�Z�P`���b�R���:����36�`F��+����v����������S�ė��44ERTT�,U%��9�x�@��N��@�"�aU!-� �y� �̯$�D�t�Q��e\���m>��>|}ʵE�ﯽ��ԁ��T&�l�%0����:���o�����	/��=N�I!������	 �g~�A/ԟ+4�\�b�H~1iC����$�\�`TI�o~�*��W��PaZC]��$���I$��og��V˧�O���aA#_?�0�,�ц,^0��t�릷5�v���E0�߻����r��R�R�$gzU 5��� �}�նe֜;kN �#dX���3G��`ټ�Y�~��H�"���8$��b$�&����T �2���J�.MY�%��\ED\MZf��_"Io�\�M*�������Z$�~�|I$���l���~�a���3��1���w�p�&��ٕI�K�7=��I,}���峨�Qn�+�����{������rˑ�G��i�<a���.K��+j�n��׶�8�~����!F�Q;��?��n�������N�BI<j��k�MzϺ�Đ�/(��$���2	"��w�+���>�״�-��6V��je��Ev!���ˣB]�nW����$(#��eU"P	noe��$�$�[~җ�ˍ_�s��n��X�A%����Y�+�� A?�e���wPt�	n��IA��)/�%}ݻ���I]����w��Z�o1ض�_L��⢉�Ӗmt��{�$�KV� �|�JS�Ϳy���fq$�w��%B }�"Gw�ZE@�mZ��ڪU�3����,D�=��I$��JD�$�H����g�'B��w��*�6m@�2(�ZZ�j ����_#�Vx�����R{�BMO_iH�Dפ�D�&)��`��� ���z��Լ��oGcӯ�1 o�Ǭ�c~5yY[e��*r��A7�=��vӹ��\7x[��&H*C ���g�ȼd�[�*	���8�z�=���s�qv�&T�8���G��N�I�GR���E�˘�달B�s�76ܘf^�B��g�ڎ�����On�=m��rq�x�O��=���b�'��Gn�7)#��FՄܩۘ.��z��M`�n;g:��e��q�NÍ�@g�X=s�6������A����e�A�O�^���B�F��з�_�?I��V�$��b�'�xq�o��0!'���R8t�i��4GL��7>Sd^��޻��D����	��7ީI�tY�S������8PO�j�*]�PH���T�H�U�5ƢE5��ĒF�ҩI�阾$��L?�m&��OJ뽇*��.��DÉZ '��j��{������4��P�w�XE@�mڰ��U
H$�3}��С�Pu/9o�D�y�$�Cw�($�Ig���ɳ�My��}�P��{ru뭨�rvgf|���gA+-�z�t~���ZuD`R(�9.^�($H�zU$�	.����/�Q�W�����D&������ ��N|]�S;��%�VE�)�	f'(�r�]��&,^�hn-�w�"�E3��*"3�ې�9�/t-��*x�-x-Q�\1�<����c �D��*$����B ��l;Cc���P���C�*�$_%ٽ�g�#D��o�{I�b��M93  {����W٬Ă8�Wa*绛�>s��M(�?���	�'��Gp�u��d�>=*�$���?�m&��OUu�$'u������2�,I w��"=7����#�G*}�2C��~	m���nM˞��QN�F�Zl�N�#
җ��WnĲT
F�.L��I�	{wr� Mo��t�n���j�D�H[ݹ�> ��LZ���Q\����*IS�i�.ͻ[�#C�$9�I%�۞��IQ&�� T�?��|��N�T쁑E��s������ϒ'y���U�f-��t<*,�̳65�4f���4v��S�kY��@:�����]͞��d}�}�D)��lm��Qt�����~$�j���l��I���
���X��h��yjO�{������%n��5ݐ 5�3,��5�!��H��r�<�W��Ă8�Ua*�RH$3}#Wf�����ޓ� �lr �G�����mvHgw,�(���3�Ò#f�ipaU6��������F �%�_h�j6�M��Z߾��j���$�&��X�v˼z<����{�"�H��({���Ɲ"ɢ��*CyN����=^�２F���qI4="�I$o�漨����ٸҁH��io��ʉA!��Q&��R��=Wb��js�I&��I�z:I��h��e9�v_m��Z�^��C���@$�,�:	������k�l�\Z��m���2�*o�~��¹��]�1�낗�Y���o�#�o�~�!Z�jM{*'�'���9�Y�˩#h�?��$v��Z=�*� �k���"R_�e�y	���b_�_L�	~$��}D�h��$.��'߾��ԏ�4N.Kr��n�[�:6S�tem�a���|ɐ��wܸ�8�Y�%^yJ�K�t�XI$�[=�Q7-=����y�ƅ"�C�z�$��[Q��nY�'�%Bj����a^u��I$��dV��I=;�$ �*ߺ������qz0uwH�XPGv�C�U)/gn_��I�gN���nm��p$��z��Iw���K�W��p���p��Ou�C�O�v�I-9��4Cs;=�$�I,釶��ރ(���2}]��н篡 �޽"9�v%S�,�S��_,�����	������6|w��)�;	WI�Y���H�PO�B��{e�p��s$k+Z��37�W��܂�V^�R<ՠ�bV*Y��dA���~?�#C�E�#��e�(���bwkc����S���=tɮ�tٞ����mɧ�t���[���[10��t&�Mv�kc��A�����0��L� Y�R�v�S���Z�q�n0�ucW�{\G&�Y
����;�%u\�c��tf�έ��r�V�t<�۞��f�.k��k+��:�<���[[1�D�)��b�rGSs�qY�-5��x�[4��}�P!����:%XOĒ{���$�TI�f���������V�I$��{d�M_b�b��-Y3�b�C
�����=��3�$���]�$�Y�
E��3�V��N�CՐi�I�哲���$Gu�(�$�M"�Z�պ$�I>�{}��RH,�B���KB,(#�;V�ک�����MQ�I����K�	.�TA%�ަ��2٤�I����U��P���S[^�RD��FB�)�6i�|����D���*D k�Ej�5��У���$B5fI�C�[t��n�x��Ux�o�	�i0��,4[�'��o.��==�"I$��"�N�*��-{P�F�^{�E$s�RA�x�A�D�6x���
w{�s[��E��&Ճ���}l�z�3V�F�#��K�<$��w�vz�d)�-J_a����E{��?�:�vk�P��g�TI$�2+D�����JU��8�ظ�CD8�WiW{D�4t�XI {vK�="�O{�Ioe
�IC��N�[^�.(-7�:>O�*���_waX H�I$���Q ��xf�K�{�Ix�`����Ɲ,P�U�I|���/��=�]�sxK�i�$�/*H�D�l�_j�Avwg�ޮ�k&{-mr��}���lc&fȍ��v՘��b;���u ��x��~���/кe�ù�dx�$�|6b�h�D����z�>f��P�R\wѓY{B����|m�9��$'�RU5d�цrO:?lI!��N�K�m�;�����rx*O��!��yZ$� �n��YT"A%�Ks{/�I$�������֔.�^�vvoUOcܾ�*Vm��wIo*��+����1�9p���Gl'��~^ڀ~$�Ǣ�D�G����#W�x�D8�Ua*�=���5�N�g�TD�����{�I,젍?v\cs���F�j��ŷ\(^��f�g��B@�ڭD�j��9{D�9���I>�v�	��-�^�sƶ�zQ%A&�U�)�Q��6��f�J�.�e3�����~ĳS]Z{�|�!S��� 
���!�28�i��UO����˾d�#f+���5��r�j̛�Đo�nł~��)�%�h�{*����Xi�>l-��~#z2K+��vk�]��@P�6�P�!�g,�A�D��}�Y��v8Z��(7U:�CX��}�`	������G��/���7:���Ԡ}�͊-�u�*��⮊j�- q���oa�Ow?W�@.��X�v|}��Z!�Z��� |?k�A�},�d9�w�7�@yg��w�ҍ�ڪϵ�^�Ї��!E��y,0`������J�WcmM��	f���Y.]�����A��M��>;W���t�d	޿U i�q#^�X�%�����d�Q5i��mWđ��w׏ל�:��� *���y�@	sv�����ҩ�oCE�ي���@���D�<��!�jwOLRO�V�CX��8���EPWvo>ˣ�R9�r������((v � ��AD��������Ӗ	 �"EU��u@�Gf�ؽ��Ζ���T��+��_I��@�`��f۷�,]�Mc$�%�n�w�vrf���4�7�մ���b�]XԦ4������f�L�/K9ல�t�v�przsuw����{��7�u�k�C�y�E�^�Z����[U��h^����M&N&E]�$|�^��C�V���ּˣ7�@MF�xf�d�Wr�ZZw0]#��9B&�T�C�j������q:SC%U �/(�����(�7����왃7X�r���e�!��n�+*_Lށtf�	�s����@�pQ{�O�J�[f�r� �|~�Ⱥ����m�8rZΫ޲�(knM���r�x;W�tB+���]� G�c����K[A�J=n&�8p���&�.���-A�q�Kpϕ�\�W����D�\}tp@^��ơ�x
X�y�������49Pu�uկ��q���sm�z�m�r��ӷ�d�ɘv�e�C<����?W��~�L�(g�?
���ur=�T�<"�,���Nu�J�����n
���zuӫ�eV�{���t�[K#�vV�V�SÛ�P�K��l�αV�/`��<f��2���Ù����-S�[Wnʝ��a�u[�4�WΦ�ա�9�+Cۗ�qf%�wtP4OBs�2f�w�e��6G��t�8����!��>�x��>��U��!���*��_��~�w6�yG��y2���f^5��tgU�Ǐz��-�;~���H�i�b�t�<�u�(I.c�t�:�e��t��R�1E��qiE^�X�+H/K�:R�b0��
�At��Q9���B�I�scaa! mi��I��Z��{�Ԭ#T�0R�9M*�,�{V(X�ZЄE ��� +�1+h�
�R5�m�� �*�"kk�! A�Ny5l "E�	T�%�V	:Ht��]��%XD��[kF[j!���[+	�Hbj�G��i%By9�TI����Ά�������zD���֝"�X�yE��PܼS���J�
%I�Y�EYH���m2IhZ��Sp�$=��$����Q:8�X��0�kd�2e�"ǖ�� �%A����$Ns)�6��zZ����@	��
�p$��u�)�p@��X���j�8��z$�|�9^`V�Lul'��'#���?"��*]P��=�Ѻ�P�]�q�s�{I�2ȉ�BEwy�n8kkU��f��3�4XmPB�'Gj#�5���۴&�U��'����v0�kv�D�ye,U�0�r��3���;�Un�W`�Xt�ú�˶'@
\s��N�nrGiٳ�M��Nuɐ�E�x�p���h{FnG��nh�5ϑ<�K9��RFkmu��p���W���9ۨ��39�A%�	�M�	��Y��i�1Z���]���Π���$
=	�x�!d��{1�۶�m�:�֞�"�Sd��p,��cZ�CvYKx���K���,9fG���eb�����X�3Ǒ���4�V��>�mx8�Y.���^�Fcl�ZPZ��,��8��^C��tvf$X�͖��ƷS9��`4��������UfA��[��y��E0K&�q�5H�m��3���O�B��%έТg�)��8��s/(3�����@�c��熑s�6o=,Ѥ�v\g3EM�0f�s���]zv��nw2t�\<;�Z����/.��̨�z�gf����x�̢i��E��N�&-���ٙ/n�U�a�����o��ܔ�9�N�m�{=u�@�uv����ԵY�o=�x���M<�Jc8�gq����6-��\A�i�ɦk-��Kx&��YX��T���e�-����Z����Z��V�,/2�-V��vl���d�:�����F��:��Y������t��].�Y�v�c�6�%����o�� ��u�.��9���Q�#��+�G���U�[ST�m��n�:9�Re[g)heoP�F6&���LjĦ��B뭨xy�m�I���3�Ǣ�]�<ۘ�g�X��c	+�n���yl�ɓ���sc��D�+�f�Dt�j`M�듁ƻt&bʸ�ݹK����=�n;H��r���r2Xa�Pq��vx0 ������s�����#�۳��@��I(�`7t�sa�Л�*�%�<�����u���Đ�+��Q�59�cZ��rmV�O5��1}���v�\�:��C�v�5'n���j,��n�r�BÃ���/�XE�Z� ���|?H�~��7�Y�}J9��g£}��O�������VY>=/����n�;
�5Ā��y�t>*�ؖ[{��\���z�\Q�i�&Ҡn��b�"tzWumɇhP�=K�@=�4�?P��uyYv0�C�Rmt�bn���D���u��.�d�>��d�9�j��0��m9�tvu��`�p�@�;a5V��@��5������ZS7�Y�@�i�!Dԑ��I���,������6/[]��r��� �d�����#ٽv/�����������$ 	��N�φ�
&q����'D���!Ƌ��y3�T|E�k;����H��e����
G�Cy�p˕�o��Tn�ck�c!9}��U����{旻�z�6����kM��ŨI�9��s�ޞIQ�Zi�VV���$�;�	 ����F7���,��ͺO�yC�m,	�ۊ4�}�m_��ۺ��F�(h�8 �9�F��<p��������7<� ��%z� ��{�o�C�C�󘾡�|=b|��O��*�b���@��%e^g��[:p,�qӷ?�8{t-��.}|{*��������+����}ƣ>���Ԯ����� H|l��~1��Wo��"���M���v}d�Iܷ �_�Z�7�~���6�������aj�"nA$�ؾ�UZi�j1Ь�l�輹��Y���5�7��F<Vh�ۈַ|Y��'���e�Z9�]�h�-�v\��U3oҿ ;��>��*钴���r�Uu�n�9xu��t���W��� ��x�'ݢ�?�9���"�d�Y[��(9�"����S��T��/ �7�U��K���Z��wel>�0�$l0̀�"pG"A;8�<	dv��aU��p-��������w�A��(�}�t��2q"M5)�H$w�j�V���l��cVg�Kߪ���޼.�� �Ԁ��m����C������_��$�ve�O�ݽwd�m����p#{~xI?{������g�����a�T����P���^��H#�:���v?�A��V�ʗuy����bT�{w6�#s�ϓ34�r�^>�����#݃D�gfh�3�nm�ǧx1�-2_ꯗ�~�_W�d��q�j]���VH#w'UBo^$
��k�'�����z���X�E��ܙw>��鶺6��XQғd�T�h��O}|�ٴ⍱�&UIٻw`�=�a��?_���J��Oom���Pb��F��tW�w
�WR��ʂ�����Bz1>=�gzyζp�=7��VI6T�0�k+?�� ����/��=�w`�I�y�8�W��$�^��"Y�E�J���6(
�6^P�y�]u���#��}�v��A���أaj��A ��e^���O�;���$����]ez�}}�
8�n�0ܗי:䑑H�p��[�=��/�\��z�]�5������[�tp	�#Y�1tK$r�4Q���靖ܲ,ϲ�1ċ�nr���;����:vݚ��0�F�u�֝�ur�V�ws�m1��*�v�+]G1�%��u���ɺ�-�׬̛���U�����.-��5��g�X�d��|�<͎+'Y��[��rt����\]�7Fܴ�n���7��1�&^�uv�+I�M`( j2݌�N+�Ih�^�b���f�m���X�c%�WH�T���������������$�� �u���:���>.�r��w|��v��b�'m�}6��I�����ޭ�w���~��������"����≸��۩��
$<9�̚����N�#z�(��
���G@��ſ}����s�Y~�A7������	 �ۀ�����d���T�Oă�޻����<!�"uB������Ԁ���ۗ���X�
�M(���p�\"�.Ƨv�򱤳�r�Ai�#�6������|u���M���=s�@| {�5^L���	�yB�&� s���j�qݚ��'O^aEɆ����l��g��q���n��;�<�jd��%���Wx����ZjҕX���7nk��g�G���}�==�@I�_�A7���X(g+�6?y׳:k�~޸|�Q$⍱A�ڠI �v��$�^���i����Q?o���+�M�(���ڋ�}cA��J�	��{m�]��<��\��
o���VE�s�;9�t
�m�$�;(�^���$��λ������N���"�#�"E�%����n��d�浻T�gKGC&�L���{���6���ٷB�'۽w`�����^�9�/W�*��gu���Q�)k>"g1���~6�s/,�*osLRz��皇��8��7���2���6���#}�BE]onvT]�ez`M+���(lPb��OZ(�g�v�7��3�����9��>v��tr�m`���׽����H�Ƭ�����;�`��T����7�.������-�aF��M:����s3f]O�(�t�n���|E��8�n+��zA�^J�m������ ��yT+�� T��췸	�zt���׋e�;���6۳L&��vpB��O�����CE����������7$$�Ou���s�J������u�{���y������� (fn������lO��O^|��׶���O>�eh$z6�r$���Ǿ=�e|~[5�ey�fV�"�_�oOU|	ܞ`�!M�b��� ��?z�e�H{�BOā��$o;��u����8�X��VFIE����+n�zd�#�I뫏~���|�n��ޯp��+�]�[�q^�ߊ޻��&�� ���ӿ{_*��RT�+���d��׵Gg𚮲���T�&�{�-{�s����z�&6Xq�8�*���lRi�6JvpW X�hk����m[~�ض-�h�(H>�(	�ޱӉ^��v)w��׹BA9{U@���Q%��S�(o��N�پ	�ɛf��|G��� =��W��Rr�g1O����@��w�$ D��򲾯�v��� �wn�Α�]�ϸ��J$nw�X�W�F��D������'z�2Wđ���'� )2mw���`7WPU�xk-���7ٝH+\"mS��c�:��=Y�+�O���,�c�8V��k�������)K�7�����ZV�$:K���L�oE��M봇c �	��:��mu� ʫ��S�_��}�?�Se�!��5c׵�D �#�)rE�U۴��e�,�6 �GM�Eܷ6c��&�tQ`�5��8�۵�����n��vs9�j�2�t��u�Q��6��u�L�Au�ֶSs��2ۤB"<�'�U�����u�ʸ11�ah��"Yi�S!�E�u��Z�� ��ԝ<u�ӄ��uet���V��h����KpB����i�C�����f�q(�qF��ͪ�� ����VA\2L9�X���mQ �{�ޫ�o�4��D�������C�n Wl�I�{�`�:�I�r[h���3�@����Z,%>�c�̲	��k�A��x�_l����I{v�X$���+���̢n��חNo�ҽV�@(�U�Y$�����{�V�=��:����wk䇣o�"MP���6Jso�e��t����z��I;��0f��҆��n
^���_�&'�I��[�p���ӵ������D��*8����[%A
�-����?�p�'zz9��JVA;�w`���@N�J$�Q�+��s����poc�qߝ�S^V'r��;�mn�7��m�L��يn����殲�l�Һ�]D\+�wF�U]�nѹ7ϥF�٭m���BF;��^Zcc}�h��]�� (P��}s�Zv{����DV`n*�S�$O�d�I���e���s��U�_�VA#�z��~���Z,%>��鷞k�]v^�Ě�����B��:�L�ܽ�:t�<{|H �%Z̩�|sw���mm�E�_��랪 �{������_3F��d%�����p�j�:jl#Lۈ�Uj���e���_8g�m�Mq�[���҉��H��vS7R����l�6���)
1�A�u`��T�l�]�礒�OJ��{�����5W�/;��qF�qF���x�H=��b�'����~�u����V��c��{�L][�ln�Z�b�s٦R�8���s�!��X=����������=Od���g���oq��Y���Q�Zsr�T����UW�V����NT(h|Aq�5�w6�w��3*	;���G��B���P�Qb_��u�@\
zE*D�M�5�.�c;�(>(�2�uƆ��眯j#c���l`����U+�9=�a�Ru�O%/q���0$�yP�83�Z8�}}a�p���IJ�*��7a3-����z�I��yY�ሠ�6��j�'b+���qV3�����d{ת`�8�\)=��S�b�ӏ~$�!����c'�T�x;|+��5����5r���WùZXwZ"�iE�t�<��2��W��-�)M���K�i��3P��t����cɧ�"^��vjN��<=�x�d�ԃ�o��k�l��v��ڡ�s�zB;�9r����G
n�J�ұ&��+c6=������ь����mv�9C�����q=Yj�VY�d��EGv�Dډݽ;ۜ��;�-�9��(���P�@��G^1Sm3]�=�s��˭kl���u���H�K�φ-��&&ten��uowd]���{��v��cz��0Vo���r�I�1��Gց��8)��*��3�ٗ�`/�B;�+O7�hߩ�PY���1�H�C"1Y� Q���5C�i)qٔ�#��9�԰HԎ��
���#��Uy��)��F�`��@�J_��C2a���iN�V�8	��2�r�"�IhI�k��;�A��\���W��D�DU�և �L#�Q\"�8���nI2�FU��I�r�ʈ��|nr����Hz����B���Q�S
"s��f�8W�Up��D�H*9�Ԓ�G(���i*��d���PQD��UN���Q���k8QTQ��Lt�g�i! �Jp�r����p��H�|���r�,ǔ��<���.�Zf"��	��QQ��PJ妁.D\�`E�����\�e2� �Ԟ�����W�2�:p��PR�F��>I$��3����dO�.{Y�7�q-�"@�V��I��l
�l�I$}��w`�H�iSRp�H�f��aY��S�(�yY���p���`�G�i"neQ �w7���������j<�Dj����e���Mj��l�8���nvu�E���F3@����z>{���$���Fn�زAvAA{{g^����I;ݷb�̯��2$�4=���%Q��$e$�x���VI N� $aV^�\�]G���ha�	�#.���X���O�#���+�y���y�w��3�}7$8�l��Q���y��n� ��u�$��$��~�w�Pu���g\n���4���X.z�v�g_,O9����(TZJ���U��1.w�u��|K��^|!$)ᘼ�4i�ݤ47h�q]�]~b I��R��M�l��o]�ē��A$�z����z��G:�Z
�1�n�u���s+rGY��f�I��ƃt=~z�Y,%>��闵d�;\F���ׁ��������ӹ�Ko|H �%]���c]c��:V}d�g�}	��Wħ=}2��S�ٟY>�����"HS(O;���,_
ƹ���w���	����T�}�ac%�	�#,>���:��] 7����|�Wwy̋�Ć����ސ쑢T�F��đ��/�`T_�>���J� o�����c��ZR�"7Y����b�7d����ߝ��׊�q���2����K�H5$�sj�,��>Ŵl##o޻?gt��{}>T��n �3�Q��R��2��Y��n�U�y|f0�<��Y�k\��9՝�Ժ;�۴�S���=�",g������M-Lq"�/m�qrjTp��f�m�&N:���{n<�m�7j8��Q�8ݵtT/~_�h���a{=�u�iʽc�ʯ����X�9qt�;Z���f���n�",u]r����*"��0�wN:9Y���[r��-����g�_�M���m� wVR �z:���KOi�/��#��+���S��XJ}%|zu��f�a����=��u����P}ގ�nS�Z�U��,{�|A�J�+*�����~$��]v��B� ��� �z&;W���6+3��O;�˴!���)�O��v���"vO�5dm�}�TOٵak%�	�#.���W�5�B�d��ʠ	���]�D�|w���c��my��0�I$YM�,"�ٵ�l5>�ӎ��vE�2���R2Kp���U@�N��l g�+�_�e���Z�J���Y����`.
k����Zu�x��w��X�a��T[:�N�N�2�譺KՋ�o]q����+�wM����q�/�����oHH�빯2	���ow��3�1>$qS�I���#����d���Jf�]�gk�|�n����v���߷}v	?N�!,u�� ��v���pZg���W�]g�I��`��X��C'��'��۷dL ���"HST���{&�&e8�����m��>����j�m�o<[7�i1%"C=�z#�$����uz�����U]#5WcϾ���TɢJ{��{�H39�7���[:OuٰT����b|{#8�d��Q�]Sk�罉͢���/;޳�&f1;��@�|��'}�T�S�9^�w`���P�\5���	#�2P'�A�g@�z3д��W��K�F�哰'��s��Y�Mn�'f�7G�5���ܱK�3G�1� ٍ�ۯr�g�WY�3�-�Y,%>��N��={��Q]ۀ�� �}6��޺��D���A�����k|H"'%Z쩀�I�޻�!fW!���A w�Т3w�����>{�ֺc��D���M|D�[�rq'jr֝l�e���M��&@`�� �ж������[��Aܛ(�~$v�]�=��Ð1�y_��2�{��X	b#"J]�6����fr�EW�G��A"�eQ?n�г��I�e��d:�d��Q���vv�t�(�{��m��� ���ΔW#n(`.���eg{ӻ�:��f�J�@�ͻ��yLs���7'4�i��hH�XU*�<�W�x�Y��23�w�ñ��C�坔��o��>���.3U�������s3�$$�F�ە@:�4	O���~��g�A���g.ױu��	�eQ$vw]�`�g���h�-y+Sh�_�Ab����+�fݵ�d��:90��`v�ߧ�Є�҃���T 7����P����������b��UD�/��v2%B�2���� ��|ZcM��<H�G�:��3��z�
�L���4w;hE���)\f�z�7\����ܽ�Ӡ�/ݷB�"{���ʘ����*6:=�B��m���{n� �3`���^�z�sFJ������bw�Z����n�}nA'�Y(��XJ���~����$�� ��m�o��Z�1;N���9�[���'�;u��b�,��֭�i�ͯj�4Pe���7Q�ܚ��>8x�K�5�1>�]�nu�iz�躶��V{k(�ຸ����suvr��Yg�2&��\�m9�A`��b/I\,h�iϜmq�l��	�ݵx�A{2 P�v�Vl9�K���jm4Zf�G��Lݛ����n���;�G�ٵÛ��Tu�b�^�,�jk!�Fn.�)L <��Ӑu���cuk��5s���[�#���L8?g��!�S�?�/.�f�I$���?a���rv�_ܫ��s����
Ø,ϵf��9$�������L͂���1oX��'%�{��Y=��B�@���	vV�$�Vm�0��jԢ���3 �������b�� �c��9g�˦^ԡ��$�VU|I�׃�*��X(�k�bRBJb(����+�O������ 9A�]V}�\� ��l��+�N�nBQ�$�b��������Rg]au�C]Ͽa�.r1	p��bO��P$7w���Է{4g���MdڠH�zM��,>�-��S�_.{�MŔ\{w���mg#}��j��n�����w�_�O3�u���|YM�F�����,k���|�.f��n�Ym���{Z44��w�8�ʅ���Z�IjB�W>˪�'�z�X'��\s	���i��A?u̡_f�زO�,1&�P&�u3�r����c������ͺH��:����ܜfL�	��x���"."�����&��>�t�~##b�S˕/����m�Wd���y
7w�#��'�$����L�Z�ȡ�[�E�v��
j3�b�M��JHILEu6�}ݷb���>���-x^Kꩀ�=��W�m�L�rAQ]��	5�&j���c�|��{s��'O�戏o�O���o/��]�	���/lT[2Ƿ�����i.�Ha>-m�=�S��k�$���p+t��7ڦffj�C<v�/��x�|>�|>Wx~$�~�w`�k�A��<I%�%U�Z�>�w� "ik���
m����K�i
��Ϥ���$�n��g���I�	�:�$�{6�[x�4�
;�l�Ss���މ!��Ġ�"�DG_��'���0�r٢\�M��3D֑mD�Dd�u����|���S?�{�Mf�$���%�-���8Dw�7ݝv	?
�Ϧt����n��_yrJ���9JR�=/sf��MwO���J"��x�9�^k�jfےZ����>'��ʂ��=�9��K��&U��kr}��Q=OA��e����Xܒ�u`�rID�\p�~>�(����7�)Ox�w�7^6Hm>�0Y-�[ᒖ���oo8[{%_e�u�*s��t�(�ġb�Gj��x�f1� 3^��x����Īl�kfL�ٿ�]^�hWλ`��O�ܒ�>��F�9lM��k�>'��kw$���.�4�\݄�lWSUj���i��_;�~4���bw��A �weY�Oz2^�m� �쪯��.�%K��]��q>��o:������A=�U_���w��ޞ!��ۚ<Ol�M�JME�uTI?on]�D�z�^V��I {�U_��˳[c�6ܐB�We�s�ǯqnN��!�lA��{/�������������z�Ld����S�ެ�d�Y�z��u�{��4[��D�w{�����X;���So�eg�KgT�ڭ�+��7�Z��f�nq��R[/c�yt���|v�[v�L�Z����e0(f�k�ոk��P�M�1�G�o�q"��XsD{�,�`:�h)~�t���b�L��Z���k2<g��"g �g���~�I�ch�b�M�i�EK����ͳ�YФ�/V��`[�9y���Cym1�ߤK�S�
/�߶q�����&!9��c(��\Q�]䇄��]ٟ*D�fs�]�+�É]0.G�k��<[ɖ��"�[���\y�VŰ��挕y��;K]wX��7�,�4�w:��Q�ʰ�Ե�ն����N?��mxY~�8{�(8��W$��Ӽ��]��jζ���j���Ш�n�+
-�}��ʀ��|w�
�s�Q����k��1����$�S�iZ��Gu�ljƴ/
���Zs�%^Y���6��Ԃm���n�+F�^���]�D��]wg0�Gi���Ў2��f*�HX��Mo
a���7�+.�S�@��u��k�HK���_L�!�uv�.�큭g@�Iְ�f���P\0g��<F�t�~V:��١]B�l���ݍ%AWt��vZ��@�u�/7�m��5��dMH��V��j�I�§�y���<' 0+Y�S�(��To�7G���FW/�.bȫ��#�YU>iG>T�Myp�OT�x���.Qa�qt��W"��v\��A�!Dv�*Ps�IЊ�T�bJtI��̔d  �#"H�'�$a�#��*�\.f
2�� 9�)V����9TӤ�9��*"���AUr&G���TDA(�8Ef�C�'�;缳Y��� ��8!��r�c�'J
�L�*I�3�<���ip΄�B�2�dM�\(���y	P9�����R��pѤr\��T�.QUEaW.�"�9p��Ar�TQ}z���"��g"*��H(�ҦST-D��ST������_�l�L�^���Gh)	A�@9ږRi��i�Pw3n�ݛiڸx�ϩN�w9�	��6�|�.�l>�+�fr�8��j���w;jmh�;=n'�t�'F#n`�ܖk¶���5�c=Gg���|��d�u��3ù��僴&�{OV6wG��lU���X�R��[��X�3b�n�e�MXa�[͖�������N�s��c)	��G����0���cuz��q�4`�dFԙMkrW��s���m�F*ˠSd+-L��ns�R^��Y���vV6.,i�ڧ�X5�����0�w)ֽli�}���׺NR�7����c��s�w)��#�)�v�h:�S��,�v�#�t#\xͼ������B�4��X8��W`ut��#\G�r�a����Hu���s��m���n���vD��=t�ծ�q<ݍ�h9���!R8��n�W[�G�B{h�9x�tưu��]��O,��W@`�]t�5ٱ�R˥��qF���3M�+�]�n3U4���{tn��Z:s�.�u���b�s0�6�bx��O���
��܈���v]�<$s��u"ρ���xcJ&n=�v;�'b@�3j�渁�r��3ʛ)�_\���0�X�M����cV�c1p� v�����D��ͨ��Ѣy�3��A�b鸞��e�����%��>?�1��ّf��8�e}�qm�����[���p��qۗB�[Etًe0Tt���vnvJ6�2�5��+p�r��=K�S6�T�y�8��X�Vj�UU\k2mRɴ#S(��i�&e�j��
��ܴu�],I�3�P��n��;���vj2���S�n�j��0�6k�����M��1�4GҚ�w�ގUnK�M,![1c3���.�M��^��M�ŉƴ��&6�c/3d�a.���,m�v��'<u�wͦA��G�kl(·QCs��r9Bt�v�:㮚Es.���&�g����;�"f�a�48���b�fpm�[��R�B�Ν�M`q<S��3���M��^�Ͱq���p��(,�7GMr��P{af�s�������� .��~.޽��{w���I"󠀮ީ`���eW��7s���0/cB6Q��Np���GEi��>O�� �N�v]�y�BA�Gy{Nmz{Ϸ���ǂ�˅9R����$_m�����91{����W�}u�y^�r�p�k��:�k4A%�ܻ$�{��v��о�?�w`]��S7$�CTG�H$z�Q����s�wTn���O�&{����~'e�QP]Vmp|��q?/�R�U�b����z�;h�����L���`�0�7�r<�h0T�Nӯn���	 ��/�z���z�<'_��ou���i���9*�2�Wٖ ���U��Jܶ%O�E���.�9�\������u�ovgD4*������Gv�k���v���{�X��������[?S ��BA#���@�=q�4�nY/H����F�Mb���I�e��{9�ފ�����A�}(�kĬ�S���7�4'�{DW�gƀ�yR����^[�񿦦Dܩ�܄��1A]~iP�'{�g�*��w��IXv��Rn�I;�޻';3���E���(d%a�:�u;Gc��[����r����7[����d���1E|^�"�VJ���<4*��ּp[Y(��d
��
�HufY��/0�K9C�L�Eml�A��B��{^���V�
1H�T߲'�{w��`��f{x�D�a��&/��yP�u�u��t�����ۼ�qݼ�2��F��C;x�l,!9�`= ���� �{w<66{y�r1����t<[���B6Q/�YQ�#VlA��v��P��&o�	���F�f��=�e`e¤�)vv��b���F��̭�~�A ���v0�(�uA��������t�q�d^Ӹ���]V-5v��@��J��W�a�w�9�!(($0pܗT'ۻ�,�	39�s޶xww�i�n!�ʪ���w*��♹$���!�O����D�{�� A��˿���b�p�U��ZH�"���O����,Y���BH5����m���'w�,����U���1H�TߺE���:D�+xI��]�dFNp]��پ�Yi�d7�q��N�����;���nn��������Ϛ�q���v����OD~����Y�5�����IP��Y��P�(~�؀��d��C��o�C������Q�A��^�
b$��1�E�0�t!�)b��k�,�eli% B2��;����
������H#��! ��ު����@�Uu����Xͧ��	AA!���(-�3.���� &z���� (-YS4�̯s;��-�iA܎O�1U�Ҥ?�w�H�W��uz_��I���}��QD41�%7�_f3�o�}	��P�Gv�%��^ї'�ky��/+�w'eP����|�ҧ�`�m� �D� >�{V�wc�	Y���v��o��z��\��L{_�ya	�4��Y����Nus]h���
 s^]��R�>��j,�����U������J���PF�-7W�ݴ��r9�����c��ln��ܰ�Y�p��6���p�+1㝸�#O�ь��JKIS:��b]2s;����ڞl$<���d#$�D:�ô�����콧c��������giɍ��b@��B���[�kWX6
��'��^��%��;i0Ԗc�&ك��w�z3Ϙ5����ghzg�짍	���s��8��%B�����]e����r��b�`���ު$N��"�R@��=W޻%�Q��ܷ�w� H$��e� 9*��˷d��X�d���
��I�v����`��ܴ�t���*�ψ�f��e�LܒO�1U�F�+�~4��*�9&*����(|'���Ϋڭ����j��TCA�2�YXH#:��=][��.�D��$憎���}��b�^C�G�C[\ݚ�9�&��6��z�Ԇ�f������}�\�W�n�A��ʰOğu�f��鹞�M�����H{�,Xca��~]����#V<��ٜk���TP����]ݠ]�Y�I��H�WB�ܘĮ�����uɌn[ܸj���c�	1K�$$k��k�m��{�ɤ����j��:�릵�s�j�&_��K�IR��_złF��	&�M���`��v]�Ge�#6�+����U��mf{��m��${��>}t����Ō��gu�oJ�r|��:���u�����G����˲A �[���(w�M+~o�����Z��xd�;�yc�U�zu��.��p��wr+Hi�`f@�����۟BI u��:L��:Vi'j��_��-�+����/��jT ��PK|�ν�A?�pv�� �T��󇴮r�Y�9��P�&Q��d`�ݹ�.�ɐ�KϹ���F���r�+w�bݗYu� �n�{���R�E���wƳ:iO��֩o�{V������_��/֠ ���TO�}�^T*H�`�_y�s�u��ě/�����}_���==ކX�&�҄��� 1�f�<	 �v�X�uʺC����~�!>ͺ�H$�쿯�]^Q��~��s��aaJm%��A�$]���]8�\�μ������8b�Ϣ�O��(����ʲt5lv�4�{�Q#��(Pi�`�J�^X��Ge߲��gօ|O÷�/��=�:���5'؇���-�J�nU|I ��d�<M��5��ܺ�I�ﷲ��f�B�F��3���{e�$��(O{;)� x�=�{����� �,b��5ҞEf�5�!����=D$.�i��ᎃ5���Eӧ��`�j�����oٵD���E�%D��'c�W����)lb�dcw������O,�q'Vl��gȖ��Bʐ�B%(���y|v�Z�r�I�N��|�1Anhk����U ��r��Oܳ�|o��u�>x�*��	9��bȭ�(;q��+��g��k�q�ڷ�$�H �fn]�I�PA�5M㝖o�WL��ꈡA�т(���2�>���]�Ǫ�R�齬X ���a�<��@��D���T�Y\����N��{�@}�ykK=:���l`$���Ő_��+�1�� z-0��؀�O�e���j�@V�ll '��6���!�{p�	��H�����*���d���yA�*-�&r�~M�FH����aQhߌ�Ih"-��n�n��������,���,Ib�۷\��Vv2vЫ��[q~e���GP�y6�O\��&���4!��k���K`V�{KH�o������p�k�f3m�`�L��j���U�-��3e!U����݌nn}s)�y��u����Avш��2��j�e��i�&�׶�4�f�ꍚ�WgnVZ�M4,����y*�he�-�.0��L���`3A,m�Ώ�>���R@�����݋ �������IY��!p��v/�;_���P�LAvʯ����p̖��,�w�����U!�?m���5ު��(:q��*�q
��)P��:�����~ �� ����Q(6�0C%�xr��K�Y�Nb�I#=�TA;����c��HZ��F��� ��%Z}�a��1�<�*w�]Q_���� ==�v=��guz_O���D�H��`�6ٌ$���� ��k�4m�e����|��xf5�'��>�om� �7��c��գ-�F�$ߺ�3�E��(�a7c����'ޡ�D�c�iWV#��7XѲT�31b����k�ӹ�0m<�~z�퍒dHl�C찥���ğk���cc���23��oE��M��^{�`${j��a)���uUy���'��s�m�_gCD�M�]P$�s��Y��n9>p�vf�s�zOW�$�R�$�oeYv;)��� a�H[2�/ΑF�a�.W�����{��+�|����)5!@?n�`�ج��Z�b���_{:a1O�g\R�4�B��X�-��;,ҤjT�Y�����=�>�D�7+y������U�ج���c0ϛ�$�n_�Afa_�G5���������Y�(�����m��zM�A`Og��AQ� M݃�}v,���W��P~�Þ5�;n�ԟ���D��:E�PGkw���R�vib�)�xn�mO!�n�|~��a�dy�6j��K;�H��Qs�{6C����b���O�%�\*z�W���/(M���9S��2��QˡN%D2ou�aPu�����ps٥3���s��E�I*��]�ܟf��ˮ;�8��yWe���t-�t�H�nT ��[J�s��h#6^�W4�I��ƢS�vci��#ƫ���L�W�w.GZ�ժV��V:���&�	��6�����Kj�^�q�A
��S^��<��<V�;ghkuRϯK��`̂,�pN����k�]n�>'���i����~��zA�j��`y~Jjsϼ����n]�fJ��f���A��.��r�g�+f<8��7�������t.��svW��ӗ�8��P����}�r��َZ�³��xB�o*r�n�?%�MX���w�u���k(�^�m_[�\��/A���!\;��2��Y��&ML��i�c3��G}JW:*��ڼ��=����њ�m+f^Yg`�&T�r�v�WY��3��`%�^=n�K �X��ٕ�st<��3U��Z��ӽGԡJ��>p�lejnVj�u,�I�*��+����s��Վ��w���+X�;k�z����M���{��_6W%��~�c�A�6�li�U�]!Q8���'(��ͱVY8$Rg������R�g8S*"��\�ƒȠ���C�sA�F�t�M�*8_�8TPS(���PQTʠN�p��!Ī2b�Rg!&$���M�PʻI�x���Wl�r�zv'
yF�	(H.5A;I ��&$RLH����:�nT9r]�Wbg(�YQ�H��������ӧTI�$�\¶<I���v�	� �	ȁF���6��ϒcǾ_ֆ�>7�07jQ@a)���UCO���qei�D����A��fz�ኒ�"��v=��vg^�����r��?	<��xT{M�����X�I}t!�Ϡg�ae��D1)�QK�7`��@K�iƸQ����ڊ:	�!p/z��� �p"A��<�*���J���ݿ��0K�YP�� oۚ+ӑ0Ș����>��T��_ r����s����p������L�ݹK�|!���ׇ��n��W?5K:B7 a̺7n����Ƣj��ڃ /V��>���	����hR�yz���VA}Rou�',�ݱ�Y:�_O�nw�`�M���:��|�+NVS�W5�ر�sZ���r�;�{��W� ���V-���L� L@������[��-E�|g��;�	��ܺ�I'=��i�,�/�&g�B�(�q5�A"Z�a)�f+)u�V�(6��-DewiOSqϔ1W���Nx�Pӽ�����d��������W��:E���ufX^�u����.���T?��*���uN�����N�Dn���ECq�Ý�@�A��k`}�{3nO]ҭʽ��I������{{.�f�%�G5�`�V��u�0(o��(���O�=� �3n��K�]W��i��F)M�ڮ��Nj�s9�h�U]�$�������
������x�����9�}���~����f��Z1;D�Ǣ�vp�Lǚ��MV�q↞���ǃMJ�i��UUx��=R�,s������@�3c:թN�(\���;����������tfղ��CL�����d}t�ɔeWWq�[�jcb��ֻ.�A.^�{�j�^�\9��=I����t�8S�匮�A^����K��*���q�)R`���n�C;�����������5�NKv����z^w˚Bv��Aɞ�WQSgC�z�=n�=��J�_!q���H�& c�ܪ� T�k
���#~�W'�^=ܗ�$��ܻ5�9;Q�>P�w��x5�ݗG^���q$�@���	���I�����z�(��L��gW��$v�@�?sҏowj�_�i����`�ؼa?P�9h�n"U۝���K��)�\}�W�L +OCY@s�^�Xy;'UՖ4�C	DH�F���I=�r�	�=�pn,�#�{�1�a���#G���.�aq�(�`�!���@$�v�l����&�CQ�Xi*Cw㣄�a7��[UĜ=������%���}�7��{]?���u��2D	���mUP$�A�=a�*U׃<^�Gch:�^���[F=km�{- eu\�2��ŵn��hj�1���.���ǖ�a�|�*�v�>�?�υy�x�{e<G�c+�^M�xY���ڎ9�+��d�}�D�`���t<�.=��I�󀃷�B�]"��f\�^u��)�y)��Dړ@��=���Rs�#��ǭA�J��'�ww��2�b~=������$}� ��vU����=�!�=M��Ben#e�6�t�N2m��2��F���qxx�'�DH�G���	�nQ$�w��N��o���У��h�o�*=�@9�໶�7���D��)�)�[;��
��U�si h�iw�L��9��2D	���ꪢI7��X ������>�$�	��v�9M�ص��֕?V���
�*jlˏ����zϓ�e�a|>��k�O��mТ?{�e�u�9;��>P�V�O���
 �L_ (zw�� OK{aE^��폒�쭪'�]D�A���(�yv �����|�zc����ݫ��������僕�G�F��9&κ��7\�k6�&%�3ЩfXІhz����!-�?���q$n�eX�}�p�c�5��j�#7�.�c	�p��h�� �M��;rg���ʲA�9� ���u7��2̼>�EH�-���}wdA��]z[�U�Au����v	 ��᛬<�/�LFMv�Q#A(D|H;'Fꧥ�y�.���T�5�8��o����pM�En!5�;b�fpXs�o&��f"Uf�m[��(������V�������CY)�I��zW�k�Y�=D�ٷd�r��� ���Q�3����h��$pF�Q�!i�Ԟ���\g�%�������-��$��0{�	gCa*w��^[�+_]e^~�Pܶ3�jC��������=z���:�D�D�O�a ������<��T(s���s�J�W���y�^����l��|��'{�|�52F7ǽ��W #������>�EH�-:��]��2nAr���ۼ�H
�ｳ��}���o_���&w�~�/�l�Mڪ�Oă{ۗN��t�f�ߞ�_@Uy�J������ܫg�i�l������U/k{@��1�u�"�cŝ�r�3���8=<��h1��V�󆜁�Z`���{���>��B�4*�,���'kc]i���]闤v�,���,�*�usa�0F�Ƙ�����M�]������V��\'m���F�7�81��K�G<��33ϡ�A��]�����%'d���7m�����:�l���Xk�T�v�k����;I�K3YҜ��]8^�n���<Vp<#sN�KWH%���WS����!����[��`�����8e@�'��J�I?noe�Ƨ�P��-NP	��Q ��,�l&`������Lv�DVu#O ��z�	9��B�ڞ��Ժy�A?f�j+���v�eQ �{w�쑛�E=K��@��\�s=�A�{*�N��$h#��2�-����*�gd�� U���L9��؁=w�D���T�Bӱ����>ϲ��z��o��_�֕B���b�$_8t?!�u�8sT��щ�4Ͳ�e�1ѷj3�H�먌�R�%��Mf�}~|�/���d���U~$�ܱ`�G������i���`$nnX~���1n6�+�6T5���{x}����njL#ʧ%��,;�����Gw���7I�j<GY�֜�ѳ~�Qܻn�)~A�U��� 7��?H';{.�#���M���R�[��v�,�l&`����X�H��9;����������}�ܱ`�O��&��G���!]���iy�	�����H��~��T�&vt���3��c	�p��~[���{wҌA7lM}�v	#�� ���=���D��W��0�`(��L3���t���lk�]7I>�ŭZM��b�i~~�?o�Dv\V��Û��b��]��
�2��_{�����/�X$�|�3:���ɠ;i%@P��:��C�1�g�` �x?L�T:<�c�~���:�r�Æ쎪p�}��H9������j�ZPp,��3�6�Fn���w�f�W�i��)�4g<=�e����V�����Oyu3n��c��|�����s|� ���{h�h60B��7<���$��!�@��P�~=����zRʍP��4�ω�8��_\;����~=����NC��޷B�.�* 
;ڷ��AB-��8PC�@�J7 L�*&ޝ����'�57XwE�s�2���fߴa<BF�<:} w�b� ������P��3�t{[��M�z�2�
���Q������%�Un,g�zd�@;��_	;��`�e�ޫ�_�q�?J�8�0�%w�T� =�k�(�~�+L�;{ك{פ�~���A�oe��8�-F�1El�+g�N�m�7h�Y��	��lP��v4��q���1-9L��*���F�S�Y��Y5*�{�:�v�g<�Zuz��D��Y�v^��Ay��]���1���!]�Z	�!r�޼�`g�O��7��e]}Q��F
ί&�4�"Hs��2�����E<��׌��{l��0��q�!*1�\1�CF,4����5���Vd�*�V8o�o�N<P�x�1[�b��Ҍ�{�d1��#D���h�M�8�8�nv������\�(�KCQ��J5}﹑[-��p��9
�Bd��{�yb$�ox�f,	�����A{�怶Z`FD��Dɿn�LCa�(�us3�cO�M�߻FZ6�&y�7Ѹ�*T11�[E�Fv���X0�!���h}���YiF�20:_
�=7w]ᶂ�h#�D$=���˂�#�&��E1�3���1DT`�a��^��3����޷��5cJ5�eg����lCbD���h�Db����te��?ޝ�:���F��Y���X�`Mk��.V0GR��h-Ƈ�j�#��! ߷FuG�V}��ٝ��-d�o���6[5;��)�l21F=~�h��#���z���t5���^�5�z�<��۹���.B���C�Q���a輄�:�W;H:�֌�ҍ���=ۭ�'a�|���[�O��Y��W�����f�b4��kz؃���s0)e`�Kŗ��2o�WN��g^����\���z�Mb��u]r'K����U��ٗ��+I�B���vk|
������6,p�r$��T�ݨ��`��z]`y����k�J��d��Sq�k���Q�:���U��V���i�p<o���i�i٩���z�g:�/R�ya�C�ԯ�qj�/2��8e�"�³�u.�A�ݺ `/WJ{���*W0\��� 7����v�5woٝ��Nu��2�kS;4I��3.f���eg5�y��۩�)��#
���b�y��v��Ş�<}�OWgAZ�Vm�kRO9��S~x�^�3�<B�ۺ���j��fAicSR�ܳ��%�[xy��H�����M��OH��o;������@����yԾ�3ᓷ��.���N�T�j=�k�$��eW�R�����ʍ�c.����p'72����贉�c�YE��0b�]Di���Jݙ�e�K��+��{���ΫY�:�p�w���mn�X/�_u��t(*
^���i�Aa�ȯ��sژ��s��Mښ±:�E�>w����x_f���ߖI�����O0��B�Ϫ�� �~��t�st�$/f�.�i��]�\)�r�,�4按��ӌH���m��i�:ybę��$$���RI	�H��I>wp)��Yqym*(���*��e�Ī�(�.Ċ��*�]�9L��&�Ӊ�)�S(NG;�^��-���J`��A���4ī�Nt�riȊ"���7]�R�� N�mÅp�k��"�/��Tp)�ӡ�M$2hp.��	��*�p)�<M��e��:�yJ���E�\L�Bs#�	���N�	&D���AAfd	U�2���NtȲ"(����iRy#	�����z��ñrJש�-��D�ٛ[�^���ݙ�h^�jqmXtX��8�5b�����6�����3eƹ]�~m{���%����'�0�ػ^���yn�^�<������Ԕe���e�0ל��̦�����v�YCv�u�XwU�WJ��m4v�$lun9ˆL�F/	v*MW�=����ɥjF&�)vZ8M;�	��q��x癶���Z`��A��l���c�Y�%���a�ltq��v� �'*�s�+��ptt��is#��q:PB��6Еu"��h[Z��Tj����Wd��^ׁ��	f�͡4�6��h�1�1v3��vk��0f��d�b��ͣ{f��[�.�ҭ��I���3x���::z�\�ev����(����d9p��*�\��6�sN˥���p��v��:Y�4f�v8��]�M|��sӧ¢����gu;�fv����R��y4��hs)���7^�Cv�����I����<X֨��r�(�\5�\���Y��7a�OWֹ���\s���>�N�k��/:�듒��I�7J^ݸ�^ۑInێf��K��$Uب���/��	�F�^����>re�*�(1q�]����U��Nݻk��2��d�44uJ�]�Yfͺу�9�9�YtY��!�&�8�ySO;;�bY1�Z#nSJ-�����M,��R�:��]�9�$8�f^[�Q�(dnãt��4݉g=;)q�-�v紵gp���5li�M̺a�L&�Zl6�\��N7��l�V���^��W�\
���ƕ!Ø�ƌ0��:8÷U�B�����q'W U����Z:��I3�G�9v��3�����L4���)"�RU��1�jѲ�GG%#��E�-���]�]�귱����ھ\��-�����g���+3W��2Mc�h[H��<Y�-��H�K�Y;d����^�l��M�e�A����x�5Z�i���qۗj�2��^d�5���^eج[���V�Sls7<m�x��7�%S�j0K���{U��������F�b�����Deo�܅��������J5����oy4�iƂ���f��o;�r�z��8���	��"�Zɮ��|"q�ƀ�[{\�L�5Q���[�ys�+�u���̞�ГN!���ǿ׬x�Ӊ4��3����KMF��*�������z��󚼋l�	K��$*�	�4q��=A�划ls��,Cz�6o��������W��u���d���Me�A�0=~�h�h�Y�$��&*T11�[��kאsl�oA�!��5y�2���20&����A��!���;�d�~��vLs�w�D>���{ޤS��FE�^LoEFV��wY�,�1�4�/��2Z�����m��ظс�4rb��SFZ#�����(�b	��hd7���O����n' AYy�ųŬ��sm���I`!v� �5�iB�߿=��g�X�J�4�yƇ�j�/,D$��wFt���4Ƃ2�}�lCg'ja޳p����q���"��J0�Q�a}���F��4B{�oM�&�e�CDes�̅�-�0�,�o��rg��zӗ��ә������	�=���߇_��l��T����v�Q݊d/
�2��'��D 54�'����"���a�皢Ʋ҃Q�/��M4q���D	o��\�b��ra��Xo��E>4��z4�D��l�*�yF��j4�Q�����lV�1F!�k\浿k����kE1�l[g��Ѧ!��l����]e�N�t"$h*��Q���U㍾������$�{���h#�dE��怶!���ɿn�Mrc�p靖�VìQ�a��Ti�Hh������&a���4�6wZ��8�[�Q����SI�2�|��,�n�ܚb؍)s��@�pC�M�t�yMg;�R^�����W5L\V�\생���kt�x����'Oc��A]ࡹ��f=�"�+�F/Y�,���F�j4�/��2[��Q�4F������2��^�u�f�o[
b�1�r�1������ȭ����_�0\�`�%cE��C�H�!�7�r�n����e�o�b'=��@[-�0#Pd߷H��ҌCa�g��n+�p9����hh���F��LT�cH�F��^��!i��F�Q��ۣ)���Q�l�ǫ
�*��f�U��S�f?�Z��H^�L-1a�Nq�l�U�qJ�7ƕU�P�{���pi����7]�ra���z��1��b!!�w�˂��7H���2�ѧ�'P�h`b��2�C��g�`[ڴҌ�j���+b�!9��є���z��4ҽo/{��b�m-F!�����X�`BQ����U�M�Ӎ����$$�������y�ֺw}��㶂2{y��bڱ�~�"��J0�Q�a����F�#G0z�78��5��ej8�:�v6��Sn����4��R�,4������{�@�6��#�#9w��,alQ�bC�wFZ�J5��;~�M4h=���j^���n��d1�n�w�#-d�=��Q���#4��ި�4��F�j���Wy�u�S%����7�aq8�_=����q�q&�$Q��n�4�5Q�����y�6��߳��o��d09�q���LS0V4[�=3�������te�o@�G�w3]��v^=��gS2�w�#e�D��n��hh�OtѦ�*�2Ѧ��篙
�μ�y������E�v���SQ�#o��M4q��1��}� W{�5�/���D�J�wB��Т�� ��AA�ׯz�^twtx���eRY[�͌����ˁ�R����d	o��G�s��1��5���)��i����4�6��Q�Ҍ�{�́��7o��<�}�	��3�a0��BMd������v�t�:v�H���h}�<@}7�w�?d��S�˄�Q��e�Լ�kt#2amP�::V�K46c�Y�>~�A�HʬBx��h�{�˦"H"H��і!�4����߽�lCgIy��1\�y�1[mF^=�F�iF1F��і!�h��>m�a���"�-�3�~�B��6�5��w���h��Fڦ��20=�N4b;�{�LCb���o���q\��F����ɏb�������b�Ti�lCkM(��̖1[1F�4F��o��ٌcY�y�=ΣCb��05��ii5��6s}�2�k]~xŹR�`�h���=5�
��*��6!�1���h#�����}�l�d`F�On�������k��ԭ����;�M#D��M��V!�#-h��{|�[b�#J59=�25M.�SW�����d`C�zɦ!���s��@���#�9�n����1��?{������޵M��[��p�dtD�9�qQ4��Q�B�\��ٺ7����٢ګ����&��[#x(Ŋ��� ���ҤP�Dg�&�i�vxL�`�t31���K+�ɵ��ub�{9�n��.��4m�z�	�.�7��� ��u�*⌢�]b�%v��۝�lYM��4����V1��ۭ���]�m��g=�g�9@�=�[g�ks�i�
�\�[νp�U[�ke����D��[��u^7���7gک�6v�9�պ�-K4��fXІh}����Hb�1��1[�g���Cb;�{�-��F(�Dh���h�Db��9�Xe�c=�z�4���(5Pj3����4���m��2��#A�*{�LD�F�f�eWk�ζ_}FvDb�A7�w��l�6�9�n���Ҍ#a�W==�鰽�tu���g܏�����Ƒm�������6!�zwtdj�Q��6�u=X��5��lCh6�$/��2���#G'�H��4�g�Ɏ∠a�l ��Gߺ��/t��S ��Q�4�;[�r�X�"h����4dh�Q�b��ߨ�K�w�v��1�������������J����؆�ٜ�m�؆����gPDz�泺x~[A�Ƃ2.w>ހ�[20#G��H�YQ�l"a�Q���G�+��^�o��_�%#p(�q�9��m]���R���j�n��*�t����O�Q�[ޞy�2�~�@���(59;�25M(�`A��]�&���n�{��=�1��Ϲ�.���7ǷH�ِ�u5�Hb�1�-�U���1�P��>�Q^z�?ԍL��c�l�fG��8����t4-��5-A�5V�9(Y�d��si,	Yմ�Y�s`�I�zr�*���*f���O��l �#Dh���4d#a�>.�(�KMF��-k���p�V��kz�E��`<�o��8ʬBd�Ch��h6鈊A�v�FuF!��Fw/�5�5^���m�����H�YiFb� ��~�LCh�y�9ƞa���-�l��w���}�㺮Oc���҃Q�s��-SJ5����}ɦ�C�Cb9�{���[�:�F76!�A��c��a堌�w���E�+@Fi���Ѧh`F!��e���K+a�򱢵�sZ8-�����Q���F(�0=w�2���iF�JFw��*�
������>	?߿K��p�2��̻�}�!k&�9\��^��@�u���9��5o���>���M窼u����]1�D${�ѝAƂ8�FN��怶!��w{��;z�s��a��;�F�Ҍ �A�;|�Mh�s���X�U:sH�F�#+��d-0�!���ѫ�z֚;5Tq�iF������C����-\�s����g�Z8�z������=�����6c@[�Q�p`F�iF�J3����ح��D#CB�on��g�^���M����g�ڎ�<����<{to����3�Lo��$��}���O��c2�ߺ�o�sW���s�><��h����{��4��Q�Q�Q��9�4���m�IV!4F�@�Es�{���|�
��b� �k�gJ�4Ƃ2w�s@[,`F!�r��e��?f_0�g[Kl81F�o~�Mh���g8ӧ�Xf&4�h��3���!l-�m(�h����<�'*=gJ06�	��Y4�hh"q���́�!��_�����ns:�r�9��f�6][��H�Tk�e�J����BE��2�۠�������QX�3����L���Cj(��=̖�l#h�Dh��R2�6.^;�^0���Mf���q�і��Pj4�j3�繑[-������+�U�M�4{:�dyb! ���=F7�>X��F�CbHe�ބi1h[װ4"o�m���v�]bC��3%b9T�̢���s^�C�-�&�m�`�k-(5d`Wx<�o~�u-�>�<q�m�b"���d.p�#�×�#,CfV��bm�)Sf4��g~�L�o���v�,��ҍF�g��w%�[1F!�E��#-#a��iQ�w=�=o��0_*��s~���-L��:-�f[�ܞs���B	u���9Ml�
�|,4��J5�o���'�~��U�L��m�����lC`|w��: ���Y�G�K���t4���~��Ot	!u���|�;�;HCa_�F�4�#G��\�y�`�s��#�/#��5�vI��t�j����l��W��Ǡn�~<{��:f%)�yh�Dgn�yalQ�i@j4v_iie����������
�o��19W�"H]���9F���##A�z���"��� Fhb�oTi�`F�ҍC�����֞��g5�� i��h��-���a�-�l_�FZZj4�j4���~/!ʾ*f9�w"�[ן�.�b�J��[���GLCb! ߷Ft�"��"��"�{Ϗ�����T�'�@�@�a>{���raL(zL=~�h�Dh���f��+�&�LCf;��C����cz|웿cŤ�4��h�R0���`FF[�w�M�h#�Cg9�s \��5���u�N�{�#G'9H��h#'y�c��)��lU��1�4�Q�����lV����`�}�*h��!�{�F�Ŗ�9��4��iD�iA����En����*��]��ǫ��܈o
.�9wN⛡��٦eS��lR̸O���+k`��l�Ztk]2�k�NiǏ�h�;��>���͚�`d�0ͥR�&�p:�ͬ�5�>78��\[])H�ٸ��BӲ[m��Z�v{����͝!4r�Wm\9�ŵ�1+v��ؠ
�ٍr��\,e����],\K��-ڪstۚ�[�1l�u�\��Ac�2V�Q��Xr����3��闥�m���k^�;���;KH�8�q��f�+��Msڪ�>v]�����O^���A�؈>*w��1�D$����ޓA�����@�,`FW�||݁��J�F��,Q�a��ti�CDh��������'1�[��k��q��F��T���5����r�G�!�##���M�1C����.��}D�g=֒�9ȏU8�}V%�������E�Sƀl�}z�LCkM(�6_}�d�+a(��4Nk9�s5ל�h�Db�a��s��M- �iF�J5�w��`^��独<T�V�bGef���3<�>�yLF�	 �_hΔ��A��怶[20#Q������O��5��	���LQ�����F�#D%��+�:ĚE4i4FW}�d1[ҍF�K�#.kq�5Ôs���#��-���6w��2���#F������Do{��G�r��4����� ��4�:V�Ն�\��aL�V�٪��n.�{���X�,�%�`b��2��iF�J3�﹒ح�(�6��_��1�=�v��g��b�S�P�뼣LCbKCQ��}̊�[������#A��ENz�#�!�<O;s��'sF5�Ԛ���z���:��#0��97�ٰ�T�9�1TŊT���'�9�֢nƗ�=�x�u�kwW��׹FX��7��Fs��2�l�6����)k#J1��9�Wq���Sa�і!�W�o	M�RsF�<�ۿ^B�b�;/�dj�Q5d`w�+3��qy�1�m�h#�D��=�d1�G�~�h�!V�3�"CH]�	���c���1;݁���Q�(���y,��lCh���(���F!�A��n�4�=�cS��/���Z�(��篞ȭ��ָ��r�T�VM44?gTO,Cb! ߷FX������V���Uo�:��F@�~���m��E1�l2÷�Ѧ�4F��l���W�����n�#-�CA���y��Xx���vn��`tjG$�h;�����٬u5_ޔ�6b�|�b�0�Ch|�Q���6��y4�hq��c';u��#�ú�!���^�S��FC^殡0�Sf4�ث>�bZiF�u�������{���0��#Dh}�R)�-�&���ti���J5Z�<��v�kl�g]�`l��rq�I��8=��������Ũ�@{���h#٤'��5��Ѭ+fV,xjPNO.�޼�4?'���h�\��,�8��Z�����=I=9��R�\�%>��4M����7�LL��Pt}k7A�3����D�iYY)��ZI�lp|�Ͷ*�+�^���b��l"<������Gq��!����zå�:T�4j���YO�.:��o�AX���U�;9�X�M|�f)�ri7�� 0�5;�rJ"�y��.�а�:R��̦���ʿ��8�w!�"�q�Wݴ9^F�۴�Td�y��]]CXtZ�[���#�����xL���jtG����EA�ܫF�WX�g�E�<�K�&R�z��j],̚����"��K�tP�ꡂ���g\��s��/�[��7=^!�����m����kX�X��+�=�������z�Y���m�V�;^Uɗ�gS&�f6���Q����i�N��F2L�"���j�wlC����v�f�g�T�T���x
�wJ�Y�r�6hu]e*�$ӹ��Ëniƴ{O�O�2n�o_I{�B h'��[��V!E���݃�o�;�X:��c#v�VT��f��Dߦ���$�5�-GMy����qF�]J�vk���|�l͜�uY{�{�Y�kTq�p��o.1�4�[�9Q)��T>:@r�M8kN)�����
x�ps��j�j�(��2I"�)8�N\=`�W�$���kH�$��"��"�|d�Yē9���B@L��p�P����N]"�M:t�W�-LyI�3�*����:��L ��+X����3�E�s�+����8W0�STI�Eӡ�Fi	�ywc�UN�ӄp��v���Q�K[�s�6Rq ��VEw8�
�VQT	���T9�ɖY!�aUʌ�*�*��I����/5
��Y������Ƿ׭�S�H���}�SYQ�b�#���bF����Sn���-��#=w��=}7u5o�F!�?w��ie5d`{{�bA��Hw��2qu;Eռ�.�!����"��A}���pl���@Fi���Q�h`F�iF!����%�[�Ng��ض�6�7�G�=$Є�������0�{���#������ w�����a���(F�<[s����]k;.;��ڠ#��;Jl~z�~�����+ŴN4>�TX� ����gPDq��4��;�he�ɫ�������CַH����a(�=��h�Dh�خ�4L���&�LCf;��C�alCiM�=����Ŗ���LCb���&�8�6!��﹐4�; ��a�ϧ����)�h#!|ޮ�
r��he�*��F��ֆ�j(�w��@�b�Ch�Z�=�N�{�kȦ���0�Pf�}�M-F!���́���9��ʬBh��s��f8�y����؍�""@=z���h#!|繠-���Ch|�R)��rj�}�=��M�r�w� ���L~�����U���m�ݻ~mc�|��I�Y��b^J��S1��c�@�]>��(�γ�2Ѧ��>4sԦ�S1�[��k��[F����2�ZY�(�u\�lC`g]߲i�m�b!!����pC��'/Ԋyh#*��N��1<�?i��y{vMP�v���i1��0^l��ʊ����-�Ȱč~ " �K���@�6�Ҍ�s��alQ�Dh|�R)�#Db�9-�T�aL	������iD�iF�=�{����z��r�T�7��m����,Cb7/8z�q�C^�o��@��tg���FNo�怶[2&j2s^�SYiFb�1��ޞ���V;ti�M����`ь:1���E4hh��w��X�؆�6��z����MF!�1���Dx7�l�A�Ƃ1$=�w���("80�ש�ɫ��Ӆ9Sf4�ث;�e�?f������]Q��Q��uy,���DM��̢��ő�b�;w�4�Ǳ�e�OI����Ce�~���[<g9�9U�G��ހ��{>X�c��hp'�U�زA��뾕�8���y깷sM�y�F�W���N�)��#l>[C��2���vSu\*xh���=`��,��S�9�P�M�7Rk	 ���6���D�SM�v@{ k�sۄB���ʺ8[1��#t*ٞ�r�C%A�#�5V�c�m�/<sc�)�V������w&��/$��X��CY���{9ٞ��2���ٵ�>��Y�[D��}v� ���R:m,�5�I��YmE���#h:�Kl�����6���۞�.n{Kc��&�,���r)�I�a�OhH�J�+gp�wn�&-����$�Ao��]���'v�|�#Y������v,I�����y�,1#F�l��A�9h]�Mz�l�M���}u���@.����H����V�a������#eA�{��Q��-Kq
���ˡ���b|v��lPl��-:/{ِ�b�y$UӟH쾪$}���s����,}��&�j̓X�U�y9/�����f�}"-��H�^�|	'��ʢ~$�;��nR���<��Lu!Ss�n#[�r��;��QV�\<�{��n��dE�2���A��?z}$��@OďovX�^�`l�p��z�u�	�ʢr��!�2L��M����F�=O}Y\�H��v�2�a�rT��<!�O&oC�/��Eu��G	68L�Wǐ�s�|���q+�}�[� ��U}UR�/�Ђ@$��@#�߲ł_�/c4v*RW1�:2���HѬ�t+�A�v�_����5!��/���R�N�ʻ������t������E��Ɯ��DG���H=ϛ���;ȩ^�����0'N�Kܿ��A�%��U����>$vuU|H$�3r���繊��N�*mPQ PO�$����ՖWGO�Yr�i%��L�a1���t��$'	
�����k�> V�^PN׳��x�}'�"I}��,�W��A�:B�ׅV}�ph �ge�Ă3��$��2��{�fL��(E֟l?6	����uXH#���A �����z�jW^>��eN!�ua�{OEp�a�;�ܭ�>D�|zk��ky/����N�^�����U?}�ν���9��v$�8L݌��.��,���rc��O9ɴ�s���P�׀�����jНF�P>s[y9jd��*�*B'޾���՝��@�	�߻�� �8?m�U s�]����xT1���"��#B.ѻlK6�,��W(�!i#���
�Ƙ�ف8Zb�o�w�g�0|�<߲�)Ol�2��G�T����j�H�Bp��Ý�D���~���Ͻ�A$��s��ނ���aN�3*��A�l"�.2�C΂~=��@�H7ޫ�JuC�G�ޔ8A��	=}r�9W�!�@L���wz�Zg�{��u2��<p	�z�$�;�L��!<C��s�s�V��g2��q�".��mt:�3v���Z�^ԓ`�/9���t?ei̅W��RD@��T]�\^�}��������g�H����Rx� �����ո׮9_
�w�Ny�T 	��b�QN�k���m5m�dm�	�[���듕ɡ_v��R �`��#REۺ��2|C����2�	9��  ��kt/-`(7�[�>��+r�2>i�	�S�'Ge�]���ݓS���	U��|H$wvX��.9��8}~�����!���eP$s��Ő�-]��{���׷T${w���0������~���{+�}�����n/�=��l ��6p����$m^�����S����ՒF�`��v�{�� �� (�ݮ� *�����b�	�Ώ�����Y�e]���'�hg����,�Cv���N(�`֫����ܩ-N޳�{w;
�ǝ>Ҙު��n
�����@�4�P)��-I�8�������4�,�7E��k�mYv�L�5���l��]	D�)4��F�V��YhC[�gX����l�H�1�C��Z�4�g�.�۫�P��������+���=l��\)=��\Ko����1]�m����k9�E��X⭵T%]��r���$.n�7�:�v��Ō7/J�Ԭ��b4e���df�~���nRbF��m�Wđ�����o����y\���ۭ�ٙ>�����������=�	��g���k�$�v�]�I��oj��K��z?4��)���ܫ�E�HH�ݻR��	;۹v����⒈�$*���������e|C�� ��=}t�}�]ehm*��3�`�w�I\d#@���'�nǡw���*�~�$o9�A#����U����'�*���d}�)c�h�P�\3��ѭ�έ�l�T�CO߿g��u�Ɂ��64�|>}��
>���
,5�������$�〟�݌�"�4{jOW�]=�[��9'M���%ó����,SF;{�n�'��Ç$�`�TEI�^�cw��x�W�{٭~�  ���$~��TE�I=U})[�埝�0�@̟��j}	 ��r�޿&Q�&�ug�$�s�A��$�b�pą�uء�c�ɻ� �퐂{�TA>���f���(BK|�5��m��zHW9�TA;�,^!��l�A{�	�۪�G��,]�7/�7���Yቘ�EGe�� �7VE����ɥ�Z�շ�x�m�����ʢ]HG�ٓ�Iz�
{7�����Ԇԭ�/;πf��U%����
_�6�js�#f��J� ���Ծ(Ow���u��<��f��lg\A����}��vX�~2��;%<3m��`���V�`GxzfuNJ��62-��;��ßq�$V�;����>g3'�)}y��̼���Vx�^��E�K� >��w�õ2|C����1�o��d��"�*W�OfvX�A��)�F���D������$,uN��O�^l�B����u@�@9ݹb���a���K�W%dj(~0G	Nq;�g*
���;�ӝ�����,��1�C	���� �Nwv]�	��`���Y� ��T	$����5��4�.2�FNy_/h�ecOϽ�
 ��kt � ��υͳxmT�T=�~�$T%:�묂H���?AyX���0�{;.�'=�7:��č�B�B�x�̽���Nyv�B�N� ~�'#�c��cwSvj�s�!`zC�a�ܫ1V�pvR:�ٖ.we^�t�빽2�[F����^�O��Ě��2��v�fO�r���O����{���I�L�I�!?��W�9*EK]����(���4��0iY�\-Y��#b�p�w9�qQ��__t~��fB����d�3�$���F^���3�^�����'��p��h�>w`9کX��q{'}LU�u�y�$O�&9�/���݋���(��G㾘> {�g���W~��N���_����?�ޡCn�d"*�ؠ����qu� (����)� 	���U}�I��S�"�4hv�� �v��H��������($J�;���|��w���z�U�׷�̤�w�_>�/ a�܌���� �`�=n�efLywLƳ�&�koMz_��6��JW`��͵gP}��b��-��׮��i�g8:ռ3&�κ�ܜ�9ܳv��53c��t3sz��J9�u����jQ�E�$TG�\P�V@h	��&n4�׽����(%�s�u���7T�(j5��v����x�����Շ�H��5u�U�e䋕t���ٔ�2��X���`�X�
��kY���)m�=��l��+��8�܊>�+,�����yb<��z��ݹp�Ժ���\L.(;��t"�[�z�Qgx�X��8�qN��+~vqe��["-���2ý��,Xܜ�Fr�]�5e�;�@jU�]�Z�%�&Tu�*	��Np�nQ�]sD���F�����M�"�jm�2�:2+���9C@�ٍ�:/�d��hǊ�S�Nwlbn�?�n�ڋ�t��+ώf\��n��F�bv5^ɛ�ۛ��&�Q(���p��楛d'��� `ӱ��ۙK���#o�O8}�i&�S�m�*�_&�p��qe�w�@܃�P
(����7�)Y�r�'�����y�}�z�&�v���Yv]�CB�u(4�B9��p����{D�ٚ[�;vv��N�{m؎e��=���#���qaUѕ������s{"�m"6㍦���C	���F�L�A
��+�*�Y�#$"�:r+$���,ʳ�b��v�eUt��
I �i�Gu.Ur(��TEQG3O���T�J��I	vTEGe�!8e�D:!q!iЙB����J��O��GjbE]�Nl�.y'9gD�< J� � Kr��!� h��9*�IHȫ^]ȓ*�:
�Uմ��iY���!ND	1:��l$�)Ѐw*,Pq8��Χ$ 3��It!3"�H�D����őE\���QI
rO���
�>������j�V��>����94;w�ǘ`�7j�6ͣ��{[��[��"C86���l��f��;-���I�".w1��c�l�7`.���\�T�\��@l<�:�%�lL�ˉsך�u����K�,���9���-� �
��qi�p3�t�H^]1a�ţ�T�Jl��u�텑�+ك2�\X�Җkv�n��Nz��[7F�n�ky�UZF��t�x���,ps�����ktbem��ŅX�s�s'�x��Lk)H��]]�$4m��ƈ���Xљ 0m	ͧ�).�g+��l�E-,�k%e6��Vٷ6���=��X��p�$/kr E�����e����ȍ�����%�V6�/��OUŅg)�0��[�aM\r\�]�:�q�Q��	�pJBX$�.��='&L���p!���s�����a�N4VZ��U���XĪ���Y�m �L틛[�:�hvn�5e�]���M�04����),��ǗZ��X⎷F�K���ݷ�զ�:��]t7S�"7s�a��F-�l�˩fa�a�vڷJ��Se�����=�u���3rkti�lI�� �q�[C���q��˺S=�)bj��#16�b&�JR1���[�V��T����c]2�J=��b��%��i�����ױ=Uz�rpK�`�,j��zC�$�Cv�1�0�4�.�^��9��i�T�U��r���X9�ҹ���{=n"vkpם�������y8GnyY-m���u��v�T/l�"�3Iuy vkl�lѩ�j�x��^��$�[e":��m��8�X�Sf�����G,Ù�6ڥ������n��z]�=��g��tP8�u�`�g���.�A^t+e.tr��ܷI���떡k
<iz����Y�(L�-#,�K��V��s���Vw<GG<T�:^������ݞۉ�:�k����t��iyJx�s��%�fI�⧉��uܼ��������)�-㠗���ú]�g�NÔ�%N�K�=��Bp���;[�Z8#,�vjR�M�ؖ8���m�B�<�Q�}����2|C����!{��_I��eٯj��~���繈	�{}T	ɪiD`P�]����:�q����߁$�{"@Bo��С�H=r��?*�f^�ۅ4CE��s2��H��˲H,7�g���c����H$�w��Æ�i\d#��
��R]�뽢J��_	&��.�$�{���m����gz
���d" �n�]��`];*�[�A�P�IP �s�r��G��{+|ᵛ�L(^^ݓT�,�r�.��6�V�ef1Z6���篿o���Y�G��4����0 z�w�x��Y/�}TA���u{�;P3'�9V�R����8G|���=�D�tC��/<��=~�C�)^ũΡ�F��s�f��K��Ӯ���`����9��gҨO{����s��=���X���f�na�m(23n���F{����<��u:���}��b����s�W�h��3�v�R�z�R{f�0 ��y�?E����r+n3�WmY�:m��E�B?,�C@wLB��0�,-�sb�{
����P Pٷ�����Ӎ�5����ne|GMD&�٘���͢]��2N���Cv��I�w�ѽ�FK������d�� ���萜����q��On��|*M��闉�bA5�uT �)}޲'N��u�`P6�
��U@|y�\rb�8��]���uI���v�E+�]en�{7sC��7��j�H�2�4�Y�H�Ct�!�U��HGy��-P���elv|�o4 2�#6*��p"VMu=�����O����W�6�%Qj�����< O9�j�,���f/����.]�Ցv������#l�i)�J|��sr���9��b�l�i�j� I��gz��}��wW��9���0�P�79�Fѹ0�!hpk��{M�y�[����Uq���$����ݽ�fOX�K&^_��I��Cj�d0�.�Зz6 ��p��#H�=�1P 	��v	��?x�d�η�ʶ�8�,H"b�����{w,X'w�9��^�[�W=�|I�������]�6."̟���OdTP��j��N�(��nU�~�={�>�sl
�l�J�k�. �F��c�w��9�� Z7��f� h�Y�~����4�Ӧ3V���3'��6���`�D�.Gwז,F{���t,Y�=~i  ~�kt(����ˋQ�����~Żn�t�˒�)�Ҙ�����\�,=m� ��w8��l�>7��ڢI9��VAO^��Vr�D_��POv�b�h�l4�.2�t��O|�ν�� �w����A�8OǷё7ث��9�x�����d�Kw`�wz�I��I�8�;�we	�7�,=�pD�@���A6C�֗������{l$w��Ɗޞ���"�>�B#j����ƅ�C���t�	 ��ҋ��វ=D��U@�6��I=��[���]��V��{p�����C����b�V�ź�;a�2�*xV�%�9^y�I�EJ�4����eV=*ii�2:�Ԗo)^;��;GP�L�v�	��u@����I#��$ps��hLf�{[h��a���Ůħ"�Ų��wUQjs�7l��M��[��A8ќuy��cWj�N�՟�����4-�9�5���_+���o0�v�v�j�즃��*��k=>����Ϊ�\�0'^oM����7Y����[n5��F]^��f�=�8���D��]Q$��$;{�Fc����j���(.��G��q)�.|n�^U!^Z��'*�$z��I=��;G_�Y��9��D�<i��E�B?/k�?��E�hB��_s�K$�v��H'w�Tz�c�1� -՚��[Jw3��{�h�l�	��~$f��V������sJ�8�2#cgI�A �n�������$���I��W��z��w���̝x�A��`�,�J�٦�pc��zg����2s♧������v��3�#%A$�sҁ$��ޠ������	�嬨#4��M@cQ:;}u�	��4鱣���*Ycq���V��9�vظܰ�$���\��n�ݾ���6B7��������L��f��ng���Rk���犅;�_R�@��g���ύ٪	�.|j�^U@�� ������{��\����P$���z��B�(��G���bY/�����/�
�=��D�n��KU��c�}����A{��e�̠m0���Us�w�c�^�Pד |;����Po��ܽY0vw{���Xp4�E�;qgې��I�1�s�5��L⦑���ߒ�qcMl��p�;;hQ$�n��rmߺ�2z�,ݜ'ٝ(m�$6d� ���l� RH����� �'��Pԉ��~43�U��6�h�0D�N�5�uD�]!��P�D��w9|����(nj�|�U2���ґF濦��:�s7��q�"U/	w��N7�Enǝ\�|���Fg��7��+���>$�t4 �t/>�n]��z{EF\�E�*@P���#w��=�h�׸��(�:U�MFC4G�O�������>O���O?]P$��87��u��9H��4��_�x���v͵��S�51u�f`�3;�����������mQ�7\�Fw]Q�P���Ҵ�{���C넿B!pA��U
 ���6�p��*��˯ ��
������>B�S�X`&8B
]������=+�A'���kܬ���H��	;��_��F���b�{�zn���Y�	#s�$����~���&�\�/��V��ٟ��yu��2���ם�h�U�X�Ҭ�86L�
"�x����r���y+�R�bw��[ύ�yy_P>��g��o*���	��	9��+� k�����C�mX�p�P�]mюuj:;7V�[���[��0���Ҹ��j2�g�ٹs� �oJ-;���H� �S�~'�=T����c@S�2���?:��ū}�@~'3=TA=��(��w�qwYu�q�35���	��u_P=۴(��}�6� (R�@�=��GguQھK��aB;��W�us�t/�{�(�I7��D�n��γ��[��
m�͉�ь�S1O��(�I��z��r�E��UOjH (I�UK���_}��{�;�i�R�������oT�f�u������"��9Sz�5V��Ң�k�X���WF�S�aC&���<d�Vj�Y�n�}�?_�,���)HJp�r|�,���{M�g�I�l��]�C�V�V5�^D��uЕ͕�{&��a��v�t޺c����v�i�D��'F�aR����g9�)�]�ڝK��n\v��V��t\v�3N�honų��<�Gb[n�:�-X��w��'�8�S@7Q��Y�k��Ғ�ms�mhພ3:�чgs�Xܱ�ǖa�"B|JŞ=Â����q!B��y|������]ա��W�S���_����)�B4w�Bn�󜼫�y�~�o� ���|�Pk׀C�K\��,o^�<�C2��V�
$���@A"��ƾ��x�@=۵@��1&\>R1�	���4����/�@�������V�U@)� ��X`%C
݂5��H>�zW�0vxt�C�y/��)y��Ho�E�n���~{&Ԙ�^�2�-�B�;9��t��n=���d�v���z]�!$���f嬨���=�U�H9\����5CP)6��]�D�S�>%������2����z�y�eX�EX�H+�R�i@v�5,�Ϟ�̱F9�J��Yaj��m�ea�Ż�A$es���ޔI���q��آ_(S(��!�!�]g���PBq��;�}�� <���ޔz���"�P$���܅n�tK	?�!$7��@�Oǳz�
<Iʷ3nQC�	�몢	�w%�=k;ȭ�VW|����O�z�o��d��߮jỌJ6�uZ��2[m�8%����
�5ڇYB�7��}_�����8�u  ���D�H�oU|Yf��d�=�|I"��B�u(IPp(b�z��ܵzȯcX(�
{"B�����Լ�䶇t�蟷ƫ�	&�s�jfL$�s;�Q����?;����������w�Iv:��g�������[��&����{.1IO���B��5O%�K-v�2i͋�>X����\hj�l�hʈ���Rg�6��s |_M��N��T�{^�����=sWn��总�.�;���U4NU�]���!v�^8�ؓ�8�@�U��aG7�B�m=7�/��Y�65w�;={�ɐ W�e�,�+�`�ki�]=�9��v�30y6PWu���oq��	ƟgN,[ĜZp���ԕ��9�ݓ�z�^�:Xcnov�pϦ�����
�������}�r�(�����Ci;�A��X�����*��NbG=�r\��ï+n����Pc�"USM���m��f��v��ٙ!����]��up��V��Ư�Qk�����2��Ӥ;=;Op�{+7�dD��U\��g�f���Zׄ,�umF������
�.lǢu�w^�K�?H�i��J�i�YM�g�܀�!k'����I5��|j%:`�E��_&!���ks���H�T����-�*t$����^�2�UݚS��Q�oD�r'�r�'=@*nQGB�mD�K�'���s62Y1\ņ�&��&�;[�Vp����,�9��
̭W�hecg���S-�D�u�3�rv�Ƭ��=u�W	���z)�S�ΔD��'لy��(�r'�"��Ώ+�#ĒM4x۬�Ug#�EPEQQʠ��D'�E2*� rk@�!�XC����ΑDT\�fH9�T�=�\��3 8<����Fko
�I�����AT^�ĕAO,wK��"<�^M�J��ÞG"/��8r��&<�̂���j�d����i]�9K��T�"L��ɸTG'0N���覨�:����V���!Ne`B�K)�w�r��9ȏ�
��\�]�.��T9�r�UDy�DD�6D��YfȂ�}|��e�H�Bw~HP� 4�Q7yb�!W=�4��^b;��n
 �n�
 �n����0��ŷ�h����#�0ӻ����O¹�ajE���[�,~_!=�T�P��x������\�	��j���(6���W3e:�#��[?�wq��2( ����Q��� �^�X�:�g���:wb���ϊD��#]A���Nu��$��ޔA�\o�T7��K�0�J�)�w�u@�=}��I�h�OE�᷉���R�~�x%�A%�\�ݺ��v20�-&K�o������
�� �}��xԣ���:�C�*K+��h�}ۜ��F9��&H�cV�^`���ccja�YQe���ZPR��H*u��$���n#V5��D�{ڐ9��Б,y4��B��� ����N���	��maަ_�]1xl�L��\��g�s�֛��$��On��u�`z��H�5�b�p��$�^��Āw���zv�;�C�S/��$A&��JIY��jH��]޻�I*/��o=���Y�I$kՊ�4I=�˻E$���1BX��s�]?%�|P�a��5ؖD�&Ojt�$�3{�V]�$=Y!$�����0�JCU�;����C���A!;%
'�M~{�m�h���Wl
�仂�/�R�Aa��I�\���+r�d����k����� ��*$�K�kl�D��e`�W���:5�������V3o\~�������Ebqԩ^3=���ܺ&���s�ƤuK��/{�{^чl�>�+jy{��^r|s;�Z�j��"q�F9.dm�x�Wj��UzX��5��<�]���v�U��\5l�n����6���ys5&q�1<�Bt�
;a{;�������Xq�Qc���e^����bh\�����泎�O\:��O6ƜoWL��2qڃ\��.�ƪ#s/�VE�n�5�"��zL�|k�W��dC���G���d� M;#�Bm�C>�2��R_$�[��`$�_v�
����s=�u���_$�;��]����7	a���[}(Is�eeW���I��z��I$�[�B�"�η��'w�oL	!/!�r( �ٵ��6I{:Q��	j������s�$��ŢJ]�B�%��Zg�MZ��{n���8�R&���I-�PI����{�'i��=K��eX���򁆍��+�J_b��āW=�7N_o^l�^��tH's���� ]�J	}���|g�q,;��\��^�8�m�%X�[2��̱���{�}����.|UpSonŤ�K{�H$�I|-�`,�mn�<����t[��A���P�H|��<�M��f�!��IQ~�W9����%ߡ�k�N�:۞�ϼD�m�^�&=Z��϶?c�Śˬ���
�)��o��5�Oğ���D�h_��H�|:ֽ��Y�����B1�P��'����!��h$�0E��+ڬ�w���I&��*�$_��I�3�H�PA#�z���"7|=��I'�I _eJI$�]�w��t��u%��uk#:�"
��a��'�M=�?���#�m�q�+ UD�y!4=�uG�^5�i^g'�2cp���Nd6h�j�5�vz���g]�)+J�^��f���~�E�������J4�_$&䆂I%��wi@�&�@-���V���K�A$�|�}I67Ȣ�ϊ�����I`��_T^�s�%�쐚	%��wh��Cv���v�{+�?�\jQ�����Ƨ�T� {��d�&��G2a��幾=1��D��[�x$t�V;J����m`�e�7����A��Va�u����,�e�U�%��_f�3�Q$��_T��I ����%��q��p�"j���g�O�f6�ε9$�I�Iv]�6Kw�l��V�6�UL1$w:�$�t<QG;6���Ť��/v�5W��o�$l�5$�]�wZ$��z�5���S�}��ς��Zĺ��B�:]c��s/h�e�|n�;IωH�}�]	�����P�I/nZA�I���eb�{���l����($�A{�wv���e+FWV�1I������]<B���WĚ��^���;���*$|_Q���|Iv��)�\��/�+>��A.ޔh�fx_�=ݣ&��6�]l$w_h'���D��*�tjy�
�xy��?i���;��/���3}z �`v�z_Yn&��Z�%]c�U�4����U��3S��9��z+ml]	���wխ�p1��f[�����RUݵW���$�-��gc��g� �-����4I$L�B�/oV� ���%R���H$��i�E$��T&��R*۽�k~%	I�˳.a�l�u0�7Zԫ�Қ�T�3B�>z����l2�.%�4I����EMFz,_%�,�{uX�nmشPI-�ƾ���<�"L#�a6��	Y,���~U�km ��$=ӍI gz��\����mN�֗��`m%l�a�藮��|�HN�@RA$�fy���].��I�k�_R($'zJ	.vN�S`��M���*�e��q�&��TI$�2j��"R����5U��D���J0�OH�<M��f��=�UI�]�uv��7��K��N�( �E��D���m�F��g��1�,��;��}����ٯ�ۨ�&�f~�Pww�U7�+63o���a^�v��Cmٹ-I������Nc�zM]���}yD��|�&�W�����IWt�#���h�"P���"M��F2���".0Zל�mb�n͸��MB]+1,%IiR,��!C�+���=C�Y����e٥�h�L�`�BV*Җ8͇g�sS���$\皧q#��ۙKK���UD��\�pF(K�:V�%tڨ�Ζ͝k�]ϛ�������R�.��>a�)tu��GvAƃ�0��b���r���i��߱�-�E�����^S��HL�$��y���x����x|�|�$���V"S܇2E$FGf�_]Ѱ����WJ�Z$�$���I4w�m� �R,��rG�唗�L�lD �F3j�AͨQ&��֐d�L�<�*`��D�>�M|�[�wF�x��Jـ�եy{��n��}6�$�옑 �~~�m�I'�����3��dݣ I|w��|�+'<�)0\��/++ ��I%�z��w]��$}uR�I$�w]ݢ�I.{����L~�4,͢q��L4LM(U��;u=����b��������S
�#��m�C5�n]U$$��4� �k��)V��lg���(I"@�iTv:��0勬6['��+����A�˻=7h"�X����]NM�cu����tW�Mt���]��)�#V4�LG 3z�l�+���g+^������<�I}�˻��%�׼�4���S�܅=���gl�϶ɇ3̶~m� �� �Jĩ���~Y�D��&oF��ǼU"yX��!�B3j�A�W5�B���K��U�I!�K�9U$J����#��+���Y3nť�n�h�0b����WΕI���S��y�#���D��&I)s�P�H]t�g�䝆�M-�N�֥E��E�f�ۇ<d��nL]"�՛��v=z�~")����6��ZI�z�t�I|�7]P���%���h���r�I��!�A��"�6k'�D��Ҧ3Ӓ�<{� �4��D�m���1h=�䌕���2Q�"j�.W��$�Cke
H$�Ca�č+�T��a��R�-t�@��i�Qm^`��^n���l�);=���c}a˝�$�&�=�	���7���I�����rm��N��I%�JI|���PI�����;h���ԡ�����	��fա����^�ʿ��6��F�b��%ߙH�� �${���d��]f/]�(�b�i�([�"KHr������c^�x���;ǃ%�fY\��P�G�HgĒOw��;��C3}��iW�UR �A�uJI}Ή�a�.|]�
u��։`R�nKt����Z4H�و�I>�˻E$�����/Z) �!�y�q��B{*� ��.�ʻH$�Ix�ԙ��|t %\�D���n�'c�ȉDX��'����혝���_$"�*D�'�L���d��vx ��c/���@;�%����3@y	�c�/�=�
�𲙣e\�Vȍ�ܧ�s3��Ǘ/(x�B��PJ���FH�0��A�~m�I?=|�O�'���HgT��H�fU�D��g�Y��mT��������ңt �&n�J�1 6��f��T��C�,A2�8

6�f���H$���U�I���r�0S`���H߻*�V�a�ţ�*�Js� ��{T�N�Z"��$�3;.�$G��H����V���^`=�5/*9l��ϋ�
m�Ѱ�K��K�Jo�w��2Q��ОIٙv-RݜaK�N��
�����q�I�vkM��/s�)$�7]R��8��fRG�r��Y�s"(�q5v���T�H$6�#���U�av�9/F�ĒF�� __>r������~��
��"�W~�BIx��������.�@��#�&�5���2�����AOS��(�hY�]�q�,0��1���ٌ�3%�	�H@$1�I!*f��������Q|&�J?�d2)؏�>l0�$�/�bo��sS�G�������Z�ux<��3L��C/�CX�-����&�͌�>P��s��W�ɀ�Q��ڠ����@����_?gޗ'��LJ�_j���`�`�$�/��DK�G��g_�������~h?�T?�����?�~K+���R���I [�H����_h~ѡ�b�R0�b0���x`b4�p(k��H2!��Ɇ�O�U���$����?&3�`�W>?�������'��_��I L��d���<���a���}��ƁI M	q:m�2(�@�|���`3��K>�R�x_�Q���I _	i#Cm(}kA������>�? _?�l�iQ0�ߺ.#!��a�/�F|/�I/����~G�$�����ÿ�k��|}�j ��@���k� ���|�z��}�����h���g��C�"+H?_�O���M}����yG�,�������>A�����������!	$�K�M=����	�_����6mel01����}�A�_ BI$	�a~�BH�������ZG�����qX�|P��T͙>FR_����$�-���C.���&�l_$݉	$�(��H,��hG�}���*�xc�Ra�G���,�uZҋ�@ņ�qX�F�w���Ȑ��ŀ�����u��?���I S �S����&E���_�4C�>B�x|�ρ�.����� G����K�'�A����#�x?�ɣ�#� X����W�}�W����H�~K韙�D��($"I~?�����@�_�!��=�������_���>���������6���XC��Q��0�����O�ş��_��sᆂ��#�_�����������}��� �$�-}�p��%�#?�1�}�x����63�>���}>��h�_/����dE$�$e�<6��$$�/�b_���E�>�6�G��U����o�>�������?j>hhШ>A�}�ZY�zPKi��������2hG��0i������������)�GRG�