BZh91AY&SY}y���2_�`qg�����*����b     �                                    T�
(p                                     {���(�Q(U$J@�$(*�%IT�$�R��PB*
 T!EEJ$�%D!UUUT�����)� RJ�B%JU)EP@m�I�p*�jW0Wvr��Ul�Y����������R[���pU�`��_    � ����T� ��*��)T�Ȕ���@^�:
%V��QD��D��w:��
]��U@]���n�B��   ���
�((���P��D��>�J[�;�{�H��
U��Z�JC=5��H;���j��j"���U(�o6�J��yH�ހ�u�Kѥ����   �ç��D��
}��%�Cu�>�R����݀�l�w���E��mH�V�t��HR���T�0   �|�%QD�ETA@QH���Pu�%R��ЂU��-۩TR�9g4�W-R�M	
��В�����m�T�M��UB��K�   �����A
��"EKr 廢�K��JT�vt"������*��*\�)
��KZ��-AJ��   ���Q$� �"B�*����$P\�*@\�JBsj�m���YhJ���T�1�(���`A����ԋ��Va��     h_,}��E#r�Ip:7w(v��wRZ��*pG@�����:m��   �  <��T�)JPT��!UT����H���Dd���*�rb(dj�2�Dr 38��t-R���}j   �  ���pgD��lrQY� �����w 8�m�N%)݃�,�2Z�>| 
�   5=AJ���a4�0 ��)*J�`L�10L��?L��!O��i�L���14���l�"d��h�bh�1CL�	=RTJzj@ � h   �cRB4ș4�L���<Pd2lQ�������\�1��P�+qO33>~�&�-8��o�=Ƞ��|����T�@}�{�
�ya�H�������y����N�O�vQ l���I^�
��{�䲧� "����7����s>@�p�>P�1�����NX�L�"S�`%1B��LP�S)��b%1	!�(S)��
`%0�	LD�S�,`�1�	L�
S)����@��L�
]���Jb%0LD�"S�S)���J`�P�S)��pĦS)��
b1,�(S)�ݔ�
`�0�!L@�(S4�
`%1,�i��Jb�0B��L� S6�i��L�S)��i��
`�0��1c� S )��
b0�!L@�S)����Jb1B�	L�(S)��
bF(S)���Jb�1�)L�"S6�Jb%��0�	LD�"Si����1�(S)��0��L��R�TR�""��Q)�
S�(L�E�
)LAR�(1J��*S� ��*%1����1J`���T*B(�L�%0U
b��)��*�A)��T�A�"�1J`
��E)��SD�Jb��`����"e�"e�
e�
r�Q2�A)�
SD��݀�RAJb��E)��S T���1UM1QJ��"�)�
S��0EJb*�!� LP��c)��
`�0B��L�S��(S.�
b�1��L� S )��#L �+L � )��
b1��1��d �
`�1P��W����}�4z�E���WZ�¬է�T�-�ze�Ģ���Uw���?�j��&���j�]}�Y�{dV��͍
�V�]�y�n�̹u$��M��9UYp�Qnf;4C�B���J۱��t���L��w�LXYgUG������ػ�2�z.9(�Ua��/ z0���;���"(K<�����-��xf]-ǉ��^a��9TGa�l5�ڪۧ��V���Aj_N�����gHmҤ����d5�ڧ����ּ�u*+Cn��f�7P�֫��5�%�P���6u�ZZ,�Y��4�V7���i����U�7YfQ�7*��H2�D��z0.;ϯ2;��һn�:��L!�#2�9l-�D�[{pT�B�[��F��� �P8�sq=2^�)���,N���*+6�]k��SF�\x��+*�^�#FV��/-����Vs2�κ�m���[������7r�#�x�O��R�����n��(�Z��A�46	h��9�ǳn�rL���s/&2�Hz����;]�M%�&�>iYhP��n�lGƣ�Yȥ�`��*��t�*f&�s2�U��)eZ�'w�cr���.�an�E]/D���(�G^1��$d��Z��" pӰsس/3o��l�4eU`���ۄ7vЏ,kp�4��rܖ�7��)�ѯ�wv�ET�C����,m�&�ҙõf��D�׶l�=����wtu�y(޶��[v�1�-�l�BZ��^�ة��O�Z'nm�r�����6ޣt�╹��ۘ�{P!OqJ���e�kv��ojd��p��{�(���/[�1A���C{��bZ���Q��`,���i���ܼ��)�����+ͽK�2NfAp,�uV��Y�g�Õf΍�t�ۡe�&5t賵n�Փ��6-XtQ1���q�z5�,f幙f�ȕm�����Y��1�s-e�tt+*�YU.;;,c@����W�+iR�S}RR���l�	��P���:j�Zk"�ӍeR�$Zi坽�4.%�Ǩ4��e�k�,n�Dݤ����p�R��f��jF�Л��"vs7E�w4��uf�n,[j��4%/b�� i�V�OSuM
��(��*�+��-雑u���9W�y��v�R�g;�2+������
���&q�B�H�����j�]�nm4�M���w):w�owɥ�T9�S%Q��E�0*���:r�9��dV������e��q�\Z�wa؅L�¬mfĳ-�4�AԊ�����+i
�&��ڽ�n���W���x07]���6��j��|*;��Ε��nc�fUQT�Ln�B�waY%x�*����
�5�!Ԓ��[/"�Z�BV���,h[ӊkU6��#��2�H7���.Y�Y�pPx�r=�j�y�b��˂�KW��nҖ�����]�3+5�u
8�$��"��:b)�.�S����$�X�Z�t�h8��n�$����z\�Tosd��Ǣ�=�v�]�l�Z�������^�����Plk�����K��Vkm�b[���=+1��:9�����ܧn��d]:MT�7OUGm֛��N��z���n�'0�B��Ń]�O:a(��%�B>pV;q%e��1ҵd�h�{W�
�ƱFr����IUͣ��cy�hVլ�"�t�cr�o�l�8�i��3^eF�XĖ��pU�:v�[gc7��v�oh�T��5]]�T�[�S�H22����NV��1ѐ̓7M��H���JƠ�sjX	���L�j��=���2C������4c�����[���ɻ���3I�j�ɔs29l��f��V�ҫ[�i�A%�wF�e�*����T�hZ�#+v�n�ƌ�t^ۺY����I�Y�����xhjtl�-����V��ɷdPW�#ï0]R�8�
�d�!�asp�����B6ã�*1�t�\�8�T�6]��)�,s/S��*F����FT&��x���+gD&Zî�U��f�a`�ܕ�̻��|�RV<x�"��)��#T��5��p�Xv�,8�T��#��W~A����k�Pؽy��Jʏ0��7�v�j������nIY���3%�����Z�7R�ӣ�)T��ݻ��؁�c.����ج,*Ch������pʼ�Ư�.7�d�v.y[��{�z5<���5M�V1X�"�����+`"���ӨMQ�K�=�T�[���{�LL��E5x�N8΂�cJٽ R�����rʉVR�˺�u�TmP�8�dLR	���"�Uym=�G����h�L�M*�͙@��[Z.������.�<�(�l`�e�Yn����m-:�n^du���t��*����M��̵wv�V�B�����G[�pn��@�
�c�5DUZ��ڰ���y��V��Z�e��hFi��VXY���5kbcA¡�����v�J^I��,�azu��G~u�`uuA`YkjyKw���i�A�ژ�)a�4�X&m�B�rm��";yP����w���4�l�*�Wn�un��OI��)kr��X�dK�hU[�l�J�N�����X�=�ɶ3n�UB�qQ�c3T��Q"ʼbꍰ��B�E�ɱctD�Y�s��I�n�n��m�������W�v��Rn���.Q�����`sr�<�BT;�F6�cS��[�G5��{~U
4m�Y+F��w�
�bسXQE4n ��5V$��r�9pe�#k&�b��U��颒���u�U���^�D��1��v��ـmޥal���b��̼үr,�F�����y{�KC�Vm<5���Ÿ�l�y���J��R�ꢪ�(�`��z(^��⃆�E�yR��p�h\�WWY�Cu��/�F�LGAȯ1�ٴ��B*���oem\��Y�M��(��-J�q�u��K�᫉��뎷)��]��6��ATY�Rsi;�S�\YhF�	OJ�Ot���q�"��r���)�7l��ct���R�4�V^T�(�6��Kn���Wn��4U���m�Bu��6��b�˻$��EǶ�!�-z�QT��pU�&���j�"*l-�by��6n�*���ݫtN$��n��ܖ6���z�-�u��<͒�-8�%�J�t(Tu��y�������%`$;�D���n<�2n�wL&���p�R��X7HPM��A�6mT͋\-x�Ԗf�͸�!�N�1`Tgn�)j���X#T����v}W���!J��gh���t��wIyY���o7���l��T�v,�t!�NY9T�_�ʣ��\��I���+!oY�P����^�N�!�t;�n����E.���BXY�ڻ]����L���v$�uk*��M�f֌5�+jѦD��˫T`��eZ�H;Y�F��t�0��
���AbVa�H:9j�,��a���tf#U����n�7_��N�#eA-X�,P����pT�ժ�,M�6���$���B�iW��%��!wwl��Ƿ��%P�lTr-�7�f&���+v�(�P3x7�m���=�G0�hB�Sr`S%:X�*ڙ�i�v��֩R�l4�2�Zl�,]���Zk�iV=4���fX��mӚ#u����uS �^^+��<�{�c�&�B�
�ƞ�۵W�w�q���U�FTm�ڪ7s0��� ��[J���z]��5�yn�Z�q����6�W��A�U7v���4ɰ���Tt�c��dbm�.��Ug5T�66�h1o!����a�owj��߮Mo/6�Ţ�,�g\	U�[�;����Rr�{�7�KͪL�p[sM۴P"�D[�8����w��i�oͪ�U�f-�<�1�x��9[�����!M�5DV�gl,{���r�0Cyv��j�v�僆�ȫf^a��w6ͅd�L�fUy���ҙ�̼���G ��ൌ�;J���!�t+������)����j�֡)�����nn=�5�ה^�[ʪ7���U?j�l�n훤��hXF�2튙B�S%T,�I�v�2�b��T��l���B���̩YB�Z$�����V�^��[����̨�8��B�Uų��e"�(����Zr��2���\ɓ1������E�6yH�e݉����3%eZ�d����;t��(ḍh&���b����.i+1f���7��=�!Ɖ���,�[2�m5x6�gw.n���F����`����*��i��_�pje!���Ν��,B2��UY�^R��Z��Ey��	�Hf�7�3��
����:{�w���K�h���6�4V�����P/Q��Px3.�`��i��h��j�*�4�Xr=U�7r��ma�j��ȱf�ۼu����)䱁w^iK`#(d�*��m�XJO7A��J��ÅL�u�yr�<���ѕi2-�q����]�A֙r��av��!^́�������Y�[�6�#.�K�{�j�K����b�U���C�K�2��2-ыk��KhV�R�%����^$�V*V�k\�ju�l�Ǐ7���{˕y�QJ�(cowV��D�-�{jˎ��l�Vj����b
�2�F�t1:1M��k�xt�r�L
�4�3q�����W�U'�H��őEM��iD��F�4��Z�lͺ����Xn�I[��T�'��i��H�m��B��L�ED���[Nh�9V�I����Pʕ���ou1�Y�^��*�f=�e����5�r���[�Z�NХ�۽����n��w�P]yL�̽��
��A֡�i�Ot�"�p�4woD��d�����U�z3[��T�SN�d�zn`ʎ�Q[T7T!ڡ��*�٢���SpUҷ�a�)]��3[���+�n�ԣt�R�3F�Uc"��"V�wi�S��-l���הh�x1n	��ӵ������l��3J�C�P�R��[W�%��;.�*����-h�O�m��vS�19WB��Ó.��*�����3]���,��2���;Ldx�^�w,gp4��S2�����y
Tl䳛�o(9�M���F�%Gh�B��(��չi�[, rP�[�Kn�k�+Z�]2�4�+[�R�qAY�mQN�u�a{�	O��#�8�Goi%.���Lc�6�9cB����ݩuk��AGfXh�.m�{^�zLգo�׃`4/^�A����J��ƧU�������طu:D"�qQ!h�vt�H���5N�PXi-Yo�	Y%<��y+
�V��jH�����[�B���dC�b'�Y���e� ��L�@���`�r��Q��t�j��L
��tp�ڭ�;Gk�ݳ�������22���E������r1��5�ww�{�wV�Y2�T�P�'Ԓ��챹=I�J�en=Ŗm��ʳLGpڭ�ͺu�����y����X7q��jK���6]阈�6ّ����@�FE��R�t�B�ûr\�jm�[�3wvU@�ӫ[�j��vԇACl4]��f)oEi;UT]��l���HL"\�g���@J��۸�VX�Ƞ3�ՏY�U�.]�.��N��#��C�^YAS�[zfh��sw(U���ܵ�+{�q^6�RO)�t���mfyJ�u�V�`�S*��f�H̫�K�XA�TQi�T35�����ɏf.SưZ�+c�+
���J�z�D��u��vJx�ܦ"�,n�UZq�ݫ�V�j��X��+d��[6;�{4�u/m�Ū�A{��J��5UG*�7J֘�"�;W�K�mԱ�m�c!*�U��c�T��K#����/sS��]=ܚ񦁂��N�ԭ�in�eR��Ԧ��^�U�5��4ނ�x�Ԕ�"h��֑b:8q��[�-��J���GN����5a&c4--��z,��oM�]EX�7�i�y~�J���j���+�w6��W��iu�r��A��m�5y��^]���w$;�ˤ0X��r�Um-+�qi�or鼼��zkf\l�,ckr��$5�.�a��b�Wb�5b�DUD�h��u�'��m[��EY����٥L��6d��8drWR�n��e�T`�5.������WÙNZ�R<�MYVi;�+,Xb���ĵec���V�%���g6Ϯ�q�V1ͧ+4;��Cqm��M!LZЕ���#�{���l����iTV�le����̠�&�P�BuB�!
*b��2�8FmY�5��Mô鼦42�gN��գiă�2a�7-���dYt,~{���zv�jۍ3��v��κ�ʋ&�
��seL�K�
lj6U���f�n@/Z���I:MnTuSuX͍�Z"��<�;��.�%�hU��Q��;v1�̔�Pv�޵�r�3^��L�XD:VaT�-�StЬ�W�T�z�[{�l��tUf�t΅�����H�k��:��ǎz�`ۑ���X�d�[���H\�Ot���j�'\1{L��;N�9wM	W
��"x*h�6P�x�	���^�	�fȗ�L7/*�8�R���܃e�a�~z�
�ccX��wF��t.���v�c��j%o%��zMjU"*nM�&������ +V�#5�ɯ&Բ�U��vK�i�n���*�\��K^]k4f�����<�D`V+���PnD���l;�.m[�h�,�5*�&�ul"}�����vf�m+Ff
�.�ؽ�+4^1ݴ�Mރ(ZəH֧�/+%Z��LD�`�7�<A3]
���RL�׬SkY���*�˴tU|�\�%�q V�j����Hg��J���<a�{ }7�߆��r?+I^���&�6�&�/���e'�0a����6��� �0'�K�A�Tkm%���\�%�b�\�UWf���&�'�K'/s���P'Z��+ʶ�+�=UJb��J$	���V�ğvê9ʹ.K��Z�E$�i�M.[�C@ݻ��\Iқ�Ս�ݴ�>�{,���[��o���J�b�K��Wf�`%%IZQ-KR��@�HH�@�Jҵ��,KzѮ�x�ޗv��՜�D�)U�WJU�ʫR�y]*�v�ԭ,J%�4�LT��TU�1*�����|���?*4����8�V�5p�N�(�&$	�kbhL���ZښG��ǿ���}������~����xA@�TEQ�E��Z�յ�X�E��*�
�H����"(*[[�kQ������klZ��U��V֢ն1�m��kZ6ڢ��[�6�5�U�1����[��ت�V����Qj��E�h�Z�m��[h����F�Z�-�0 Ȣ� )"�"*�� ��[X�QZ-U���m�*�ض�mj-�h��حV�TU�km��m�m��6��Z��Z-U�m�*����E�clZ�h�lV��EkcUh�m�h�ƵX��j�mkEZ��bگ>ͯD^ ��0��uݻ��@�#���ud�I�+����1��1M˗׻[���7�yX��� ��^)�/3���^b��ޠ�u-5*$���9��DE}����PE@<<<!;��r	���G��.��"�Q??_����<��N�^�[�T�aK���y��%��2�]�S�]��XbL���Z)$r�/m�P��Z�<�ڡF�w#�3����������mm�γ���Z�ڿQ�IQW����&�ET�aI�"]���%��pΪf�%25F�:�ܮ6�s����0:��кR���73S{;L���l�]	���)^��ZuN���k;ʹf�>��v[5���NbqJ���&�̡�eKR�7���u��9/7�Vt��W�vn�7u�z�6���q�+]����h�\�9�Au7Qg|�Bu����x����4կ^�d�;)��+[�0S�l!p�$�C�����0`D�us�a��53f`�]6�$��1x�;�6���;;&fnŪ�{_rB�][�yj��u�XF>T�Ƴr���EҘS�qe;�)��7a�䃱Y�}��(�:m><쭫��*:���zFǶ�VE:���a���OT��{�Ta���Ӷ����ƒ���t�6�"�f��黏)ҧ�K7{�k��R���7��m�iݽ�;��m�Qjrٜ&N��ۺAF�Cd4p�-��W�{�.�ݤ��z��82�92�K��YB�����8�U��:�V�TXQ��L�X����W�7F�VY�]@gR��^�47�kwB��-N�6t�qF�@���w-��<�S�����ׂx�H��6`5��i�K5���ެ�jwJ��|U�ك��`�Ue-��pU͛�g{6�r�b���meYӑ�����.��[YX}��������{C1�ܔ\�����K�c�Q�3��۪6�rbt�+�(8���VWHw��A���N��c;��3T���ȏb�S�e:�پhSM+vSı(�;*��Đv:E����jtʫ���]c�4��z�4�0;��B�Q�z����\��gbe[�e��6$лf�p7�D�.���a��=�7{jٮ	���]ڡ�9�Rl�R=�.#�:�
�qދ�_1#@��qۮ����T�A���
�ۯ]s�j͜�q�����ޭ{Ĥ�P�z�j��;���DtIT����wfʸ��x���9���
)c��w���+|r�6��iݮ��MQ�%R�ˏ1w�x3�ZN�ȩ��z�;�q��,�jZ"��&��g0^о�U�`��F�eҰ�h�fg��V���+�j�w=�*�2�O����/0��U_e�62�C�Bh@k�e�L�^L��+�V�nm��eUjG"f�*�ue�	u��#��:<�C���[�^�Uf�ʛد;����rr��LsK�5��y���/*��;���6V<��ol��R�#u��.W�W-�-��X��ln<eQ�1/�Dn�����9�j��W���\є���R��/7sŔ�μ����n�G�ޘ*�3���JQٔI���x�u�!:\S.�J���7�<�-ڮ���8ycיj5xoo`���:�{����ڏ8.� T���MӻƸ�G��O�7a����q�VJ��f���L�a^�зu�dta�ɗ6��L�C��x�m��t�V\�4��j�t����ҹ���^"H��j�w�^Aӑ�.J_-�}�{З��u���m�)�����m�٨�GC�*���R���r=ot��7v�Gh�o+�e�݋�Xg/�����j��~�:L�e�Y}/��A�1��j���a-���#1�xaWȜ�4��7k�wz�:�Y�FS����^�k�պ��2-�m9.*�,�]�,�"���wۇ���U��`����w:���{M�:j��tb;�{ZE����1��G��$�ȉ}${/_���v��;Sb�[�ʜ�j��glU�I�4��N�r�ݮ�e�wvՓ�-�j�.%�V�Q��l�S�7y/��=0�ۧqu�]�yV���*��ŕ��V�BeS3/70ځ� xQm]�y�HCE�kBS"�V�=zkmu��1��2�;���hڅ�n�W+۫��}��:�xZA\]7�;��ѽT������
���.kl5�7���X�E�u��v��*�y��t"ʙ\�MM{.�+*.����Gz�%`����[dǗTh�N�ܣz������o�u���+����C�#��ӫ
�r3����i�]j�W�����7�k�k�M�M�Ֆu�"��:��y��Q�+o��o*�/���4���Tr��UP���GnZ3��<$g��]1Rn��g]6�R9��ur32.�U��-k�l������;V�v$����fǗr��}��\u��Gz��ZԊڮ�R���vUR���6nU&֍
��;xqlq:^�1�F��V��/�-^b��]״���Q����8��>f�b�7�O���綯�-Gu�b۸l�mk{6����젧:���6q��ߕ����R�����U�כ�Ȣ/�e��]F�$'w��]ˆ�&������?7�'�i:�}�-Yw3��h��q�r3����J�gG}��&�v�1ǘAʛy�Wf��7�v;�wG���;�&�5�s�v��{]��l��kk;p��J�o/f��f����ee�f�Ѧ���(�J����so.�6�6��S�n����4T�'�;-_e]US6�k�2���^�H᝜�k�u�ZJ� �����י[��	+��j�+=yq囷� ��r�v,�j�rV�fU���7�_X8�Ι:�K�ޮ�Nܾ�d�� �������+�y�j�����ˬ�\)��+-
�h�=�,ی��Kѷ����I�6Q2C}�L7��=�9�K���}���uEY��t}܍aThE���T"��F!�W�5d��K�]�[U�p�ӃkWUA:�鷘̥���XFqu�v�F�U.��˅t�/k�ۮ}/vU�wY{��鶳R�8�ʢKƺ��(��Z:���v�cݐ.`����gE�{;���i���cU�i�ʌ`��v��e��f��.uT\�
X�1ck�,�b�6��v�<���c{����K�t�T�/i��ԩC7YT^�N��.*o����h�tn�*K��Bs�	T��W]��;6�	d�YϋX�F��<�H{y������n���FJ˶i�$!�:�dv���j�Uw]+�j����t�:ͻ���b.��U�|s�*�e�v�]_v�K۶�y[�+Edm>�z#%����Q�F�;�vr�S�4�wu8���FFԤd5.��f&1�v��t[K�1��\�n��-m�j[�ڬ�Zi��^*�9"{N��[�mK���-:�a˫y�2����ԁ�շ�|�YA�3����b�Vߖ��Cݶk��v�����U&�^�5�,ܺYF���T'lVNsSs�.<uJ�0��Fa�ܙ��X�d�^ƫe���^C�V��bR�����(JJ�������^m[�t�^�+D�[(P&�����0��\��*_^��ws5�����5��~��r����,�T��z�M�4��e�f��hVl!��v��8<y��u�
�\�J�ˡZl*	����{��Kg�vE�;C ~~L�\5%c����Bla��'=�R�ֹ�s.��˷k&�o^aQ���d��C�N����ox��;Hm�W�6���V�{3O.��۷��pa�mn^���;v�0����*o�����u�M�-k��>Ƙ�ؼ�LnW���e��܄�"�Q��k�ʧ�u癪�k�"�]W���utv�]�/[���mR�s�>y�|�:��HK�ٴ<���+�Q�'pY��>#�k�EY �����+:�����mm����W��s����
�M�M�hT�X���~V*���n���.横���]�;�{@�5�U.��oMΙ�z�X0qu�w�'�O^�YG�����BI7���W�[jb���κu�ugV�#u��2����u����k.bI#\p��=3��h�3E^7����������3n�WS���K��j�[u|��T�U���r���j��k �c{;:k3�����\��2���������PY���Ux��a	���#��R�k���Y�]ʮ�!T�X�K&]���pt�B��󫶗^����oz�;}K�*끅8_]Q��E�����l5[���]�3�]�rﭔun�ʩBɿ�z����]�ڳX���϶���e���[�EWY��r�W��֍��&�>T,��w
�Õq͝���el=�����ʹ���n����
޺aI[�`"����v�L9��6h�[ťf�7 �.�������̾����]��Uy׻U��47�Sy"sojm�o!��і�-��V.�d�@������t\5\���{a�z��%X�,y%��,�d,�+؎YAլ5�{Jν�1e���5:�H��]�^u��y5�#���;d}-�ξ�_	�L�Y7n���W�G��[�HQ��{V%j=�9����H�U�@üp脼�<��V��aF��rDߦ�ڂZf���ݱc�cU:��w�kCN�U�U�V"����w،t�aW������MJ�#^(5f-Ϋ��>�\��27Wy����l�&v�4{Z8��j�+�8iu�f(t�u�3�w�-
F�Ct�S)5zAr-O.��˝Km�uu���
6�.yʷN��״h]��0mv��Dh��yå���꼛���"�8j���o��	�ĵ�!.͗uW���sV�ļ�t)�v5��t ���DԻc��9������
����^6�N��4��ta��q��P�o��M�D嫦ssٵ9���U�vUf�����el��(���#��I礍������D����;�p>]g�n��\��Wg��S����P1�*�^�讽�=&Q��B�P��/5]�d�\�6m�m]�O�e����͵����Q���f�e���ڷ�ڎW �^9�V�nջ���sg�vH��}���f\]�.q7X\��!��!降��kc��;�{7R��Ü�y�H�(fw,��--j��
�`��Tzկ}6���wI/*yW:q_RŔQbr���Ag��BcX}[�� 2��������˦`��$�����hx::9Af�y��KP�#�4_,阏%�(j�ɛ��B�/�����f��DiR����sE�n��'��J���u��<�jO��n��s/�9L뾇��}��x��wo��C3�Y)Y�KAeMq�d���/US�jC��bw"FۛK�m8�oN�e���uT��eU-��vh3}��f�Q���m	=Ww�O* ���Xűb�p<��Z;4��֭���;;Nn{7ك6���٦�![X�mw1]��ܺ�[�ֳh���C��-j���V��&��"7�_]X&W��n��p�KO�.��Ku��#Rݝ�[�eVe��z�S�Ur^V�Ƹ�������:�i�}R���5^^�I�سX�Cl�+X�n��܈�O$����e��^\*��Ӯ$�W�ka�1/7}f�}�^�Y���\9���,��_`d�+�L��S)my[μ)_���fڽ��P�T�]�w-e�HF��w��Q���h��f���Rg�Z:P����gj���n�T/Z�r�4�2lc4��F�mee�Sk�Eu��`.K�6uI4�;J�l�sh�;&�n��:����¢�y�%z������h����j��w}q�y�c�W���M�n�eV�WJZe�c77���d����j�5�m�97)�m��a�1ʖs;6�;Y}z	(WN�Y�ٚ8�j��N�]
���L.�X.�Y��ω�U������][n�s��(��B�ʭxz��T[�ӕ0f�˺���N��SE��݋�� ��L�v/L^ݝ��i����f���D�^�=��~ꩺ��:�0�'��ܼ�����n�����xTX {f�ɺ���yx�H����A[z�[��F�]�z��b�'S4Q���oۣRu���s���Z���CW@�U-��)��2'B.f؉�F�7�Wʹ-0�rNP���ݵN��6��<��{N�eL�skr1���D�]�*��9Pu���ˌ���t��k��U{��K]�Gy�O�����tk��Y�Emz�����lkV����������3VV:�L�����|o�m
��7���\<Wkj�{��p#�eS�쮇�R�r�v`�{nW+�	�E�ݷ��4�UI�l�ۑѵ���z�n⬬*�.FҤ���#[�\_`�5�3�е���T.�(r�\�p��C}��!�;5��k�>��(��XV<4j�+$ݚ)�<y0���	M�L'\���б����p=g{Z�xj馞(%�9�6��]=��0�N6��`#��b��u֍ws��v�.
�KIwͦ(�-"����v�i�u��V�1#�-�9JDN���/H�F������@�=\�����@��c�򶪫��#��]HpS9-�/WnXxip5��oj�ʖF��8���Y�������It�eh�N�e:�^��ǚFJ�F��ab���"p��9f�[��[�a�}wU�!��V�v���M>�[`AY��ϙG�kU�I���w
	GW��R�Ku�-@�}W�%8��F��A�)�u�X�͔f�	uu�Y�q�WR����a{fuΠ��&����u���(���m2p�E���P�P�y֘XPc7l�ʺ��vWIق�M3��gR;�@����UOw���oz��U��M�ڵ���kE����vj�c�W�1C	�Zt�ه5¬uV�~}��<�E]㫃��Fx�w�v��[�S�p�¡�}Z���m҃�W���򯫃vw�%�c98�R� �	��{��.���1���u^i������4u�;���-j���gSWdʼ�k�d�:�A�Q��p5���}[�3����JP��8�>�\3*��O��r�2.�R�W��L�̢7vz:st�[I����3���]��B���S�Zc��9��}�j�[��ߙ��(�
�,�����<|���������7}���'��v�۷n�:t���ˏRJ��g�X���KL^ܥ�e����j��N��2|��v��o��|Wr㵹�B�շǱY��K��}_47VR����͌&�^�궽B��q�m|�1d��=sK��NWRY�ѹCëQ{i�k.SV,XZ1��VF@���A��t.�[ۂ�n�ݞ�N�9:C�����.��v�!䓔�s!�0���i�j�0�ňT�jHJ:^��,��.�=7[�&�.ňN�!�{�γY��L�j�2k �v�W���<%�Mfԃ�cl �X:b�!�� m�+�!�Vp��;����q����]�c�qf[(�v;��VR^LXmѺ�Cm�][[���ۈ�n]ڏ[G=����..!�t��q�nG�$�U�M��Xtd�ӷI�b^�Hsh��cԃ
im��rXd�1�>�/N�`��8͂ͤ��k�(�/��<�Cu��[r�t��t)�%0%Δ0�ap^��P�m���.�U�Ŋ�-�Уa7�V�V�ۥ�T�\�zUs�bۮ��<���i�إ�y}=<P5���B���hK�.eM)oZ�#�u�$���b�Et��M��n$�mM�uhԕ�3j��CDH�TG��n��9ein�c���$ؕ����g[��klm�X@�N�0s�[a9�9�m��m( K���>x�:2\����.�\/l���ȷ�N�q��
s�V雫=�Q#�v�3;I�ȼ�r�6
�'^J� �T��M3@J6��H�\�ɞ�3g��9�^���H̪��15)L�Y��A�C�K����M�m�;e�b�m���&yZkNL��-�J2�Ѕ�)�4XR��0�ږ]�9�����bm��]'[��ͱu�%�z'�'������j�:�x[Ȯ3w�i���|�����\:h"M*��5:��1�^܈4m�V،M���
��W3���h�@lW2�F�S4�T7c7%y����<�x�,�l��&�9�#:�c�vkZZ�m��z��n#�lwd�6�x��W;�w��rt�ˍ�M�E��x���A�8闛lm���" 鱜�+A�� �r���S�t!�M��Bb�l��Gi����.�仃�Kp�j^ȉx�L��3ɣ��)��X`�m���\S5�v�m>ݶ��1ϣ]Za1Ƌ,M�f�n@�\�۳�VR V8�	��b�uF�t�'���h˶v��o1|<6y}<���\��`��]�g*�Ml�4�z�A��j㙁�ۤ��Q�m��q�$�x�g���.k��Y[3�lҨGcvB�{B!� �;]�5=��7�=��[��V�ͭ�ڦ4k�k��t��=F�Ϗ΍���N
�C=�͍;�/4Zx���礡�@�.M�2#g]����aؘ!66&��`mDЮ��Q����{j�A�:l$mh�d`bܩ��iŸi��Q�v�b��vA�\@7�[n�\/fń�a�!���9Zkt��kv�w�L<��U:v�]^��&�0�m���X�kux�!�M�%��S1 �X���1�ia]ĠC�(��SK��ZKh,&�ЇD<��=aLv�a�y5�;n�&��ە�Q�IUƚ�)��d-���w�§]gt�ƇG6���ݩ\D��^.��e!6���X:�K����Fd���홝��m[m�赡KW\��d�8�8�z����,6�lmF:&.���w*����(�ɷ�)�����G�a�� ��]ڋ�)8:��՜�d]���N	��v9��mu���i�a�P�4Pjb��m��u)�=Z��í��<�9P����]	�l[��lC=U������8;���woo0nq����m2�uSg�v���]��q��Ξia�����:��8Վ�	h�̭���9Uu�t�V�ݵ�@g�Z���^ַ���r��z莄��i�7W�g�4�Q����p�X2��N1�y�z�d{`ݰu����]����Y95��k��t��݈uې�l�P����=�)�8�.]4ZachJu,#�u��6��뙧#��vFكCm�VYKĽtk�h.�mջu.��q�jKy�^[6Ў�ƽ)s���m�\h;g��k�-ʾZ+��۞��7c����&�v�D�ԡ�<re��҈�v�-:n�]h�.N��kf��_�f)�,�!Mt�J;YI4��эdV��z�nk{��%��	���'i^�:����e�o�\W\rf���5z^�^��'E�LRǆ]a���-P�ˊ$[1n��mej�Q��%E�&c�	����̰�	k��-�U���JR��2vx-�jwlqc\^���7WG�k^���nRKθ��v���];�2�=;�lsɫo-hu��;1O]v��ipF)&̼$KHs�p-�^�Ȓ�
��`�؛�'v�mjyӵ�\�.���=�.��R�Pl�DX�k+Vii%6�m�;q���GD�� 4 �YgN����rp`q�2lKtCBZAuL4!l2�(i3N�M\)v�D)7�$<��s��M�ٻ�i�����g]���c{Xie훎��䋚��		܎���lnr>.z<�1��1����;z#�syĘ�,-G�kOAc�B�,��u�M�=4y�	�S�Oo�	q�v�֞�5���A�������\M�H��>|���Ob�zM���j��z�^�Cb�U�X�p�5F�-�\�(��5T�V2#{%&�k*���R�����o(�Im�Fx����fUlV�g�=uc_dBc��[+kG�5;e�֚���"�I�ni}׵��n�o;n�WZU��%+%�1������ffIi��*��ԗ61�Ѩ�X��- �!�$P��f�Mi@��΍!.�k�l�����1�	ev�7@���Ԅ9��-L�iv�Q�c�M5��6@+N����A��"��� ��Y���K��k�[��Lkc� G6$�2ZgcK3f��ب&�x���3�%�K��cjf���q� �:�i�<����]��6�g����	�#�ų�'sH\&���K�l�5��r��Ȼt;����\sͪ�u�2�J�2F禎�7��KjC��������P�"�/.,Ih�rj�W�㳏����'#|�[;x�� ���ѸM��	�Z��R �e�.F]4E�G�$�$��;=�XL�@�+ .k�����-�8�_Ob�梔�n���O^ �7Z�.`;]�n��m�g����E���l=�æ�rװnݠT:�벸p��6kBf4ik4;i[����t�mӝ���>8��gq�T��L{e�t�wX��8�9���n�m�[�.&���X*���,��\�L;pg�t\�tGm�p^#N�L�݈��/MB���V�<��OY.�Jb��Zn�,b#n;M���uhF���;F佋Ѽ���񭡔�nދG;\<�GfI�Μ�n�{s��VShJm��,H������-Ω(�!qٯ��u�Y+1��1`�]Z9��:4��[]�Y��x�m�CSl�u��B2�S����st�o,��cv�hU����ٻ[fˮ�[h���ĮK�h�LFd����[A�ۇ����9�2؞wQvMӔ1�1��)��{%#�����s��q�v��v��ݬ�e�T�i�	�9 !���Y��[�1;�8bv�r[Ǝ�M�FÕ�(�̫Z�L��`Nn�e�`n��������F���,�:�<]ͯWF�c)��׵AbNiy�tÇi�!C ��.
褸K5��	��ѻ=m]'1�w��C���4�JCiYkbXB��Z��e	�\Rv��;�m�e���Ħ�$�0B�hR���r�<���U%��3(iB���b\0�F$o	sm�ur즫Ţ_j�3h&���y��ي(�k��2��m��4�)��`M��l�R�{;g��{ n���![4fl*�����XaVZ�I*n��q#��̹SB��K@
��q.sC��yw%���9x�^��]S���"X�v�+�Ї1WY<K\�7���=����-9�D�c��yn�979�1��:][�͆�h�1ƝkFܡp$[,�Re]j��v�̠#B��ٹ!za�H�*K%�.s�+<<]�=�qu�uݷ&���� 
e��`R��-�]]P��k:ұ׷vw�훮�.=6�Q[��,�Չ)���7��О�n�]�3T���&��6u)6b+s����k]4u����@���璲���Z���.�6I1a4����÷GO�jۀ�u[����y�ہ�<t�a-b�>n��n�=�u�����v*��xu]՘b�\
]c��D�IH;��<Q�mgu��/V���%PJ�X�+4m�����IrXaf.�r�6(Jd#C<V:���O����5{�y��.�nm,D�b�[�^���ٶۙ�1u���\o^'A��++6�B��P��؎@�O\큲�M뛫=u΋�jCM]z�a2��EFS��slr}oU��uM�ӗR9q��-�]4E�]���\��R�؁,L,SX�';{�s���b��˥��f�8Isr6�6>#)N7�<���k��1h�/fv����J��6���{+��]��m͎챻b�alف6��Ѕe���y�;iw@tq6ƻ��XiuB=t���npe�;='<N��"�}�:7<n@:ۥ�ǃ����7]lKg�Z�ƭ�݄b�� ��s�c�\d��8�99�K���î٬��#�%�לuIB��bmQ����8Lk�j�:ηd��u0�-j����̵UUUUUU�
�����iJ��K�L��A؎�v�ݶ��?v`>r�hR�(�D�pl����u����O<�6B-�6�%IvG��j�юM��B\�������X�3��)����2c��ۘ���W�qV�['9�w#��WqA�,�ç�(! >fۭ6�F$�M[�OY8��A�K�x8��"��|��0 [�8{��<*w]�I�j0(�Q� e5"Ơ�1���%�Q)��LQQ�#!��Цf�2�)!Q��h#�D*(#EF5�!��lc`�$ƈ�Ɛ�ȢѓF��W�b�r��ch�)7-�Ab�ML���vM���TcQ�1dClTTV$��QL�5�^����F��h���#h���a
��T[F���}�����K�2��;\7P�e�K;C�^��<�'<���q���&K+6�j�*��,�F��5fp�S[� 5i�Ӽ=���v>����S@!u��cA�笳K4����(]�XV鶶z��6v7J�rWj��z�6�w��̀p8��i�5,fYFW-�g��.�{�CO-������d����	)r7n�fS"	  �Z�
� ���K��6R[q@�X=z��=.cR�a��2D-&�X�V��%�<�n0k��e�G>s��M��RZ�Mz��gB!G[���S[�
@y�E�F�%�����\�-�[�yn	V��ͅf!�̴6��ͅ��aVuu.ص�ix�` #�n�f����Z�!��W��m�q�����M��^֘����QmHL���n� N�c�����5�S��s��N ��=)\��25-�č��%��Qܔ�#��ݎ8�v���cd;e���.��x�x璔&�f�BXhdРꐀW+3�J��îG��L��x��۩����-q����¡X��j�2���fe`B"����y�k��{qm��$L۳���#6�L�3�|�o�׶kr�Q��V�N\�[Vx:�9ۨ1�f�ג0�O��ט�#v%x$�mA�=�,;�݋�:G�Nrr�P��qǧLcs��'���hh±�MX��kH�S�i�����E�LK5�=�B��i6�F'��e��W���R����XLه4PQ�܍��L%�Gn��O�6]�p��kd��	���խ����6�f�,�t+-R<a���M���GS��ʐ�zl���P��ശU����v���C�8�r�Q�Ғǘ�������3hY�z]q���m��$0Ĉ�@�m%��͂�ެ��E��,ns�s�E�/c�t2<��7��pY.�μOF:��uY+s�ݔR���b�%ƪ���ZJ�E�ŵ��̣m���8�,�fF�SiGZ����������;3�
�^i
�F��K
6u,e������P^h��R���-�-��JaR����y����)	`�X$��֐[ X�,a�2�[�C���KF��QU�l�!j��X��� ��-b�����A��# ▁)P[�A����K
�/S�m���G%;ݢ�R̫K��j��T�]�����0�u�^͞���̙q�te�]��1�t�����3P�?H��6v�ܾ�q͒qݐ�z��ۙ>w΀�dbRHċ�$�ֽN�;���{w�m��wKd��̶͝l��"��|U�!����	���}�?;��D��Oh��+gƦ�mvT�л|/-��݈��v�$���ᨩ���pN�n���	4�Ŷ&o*���*�r����+���X�E��1%f.i��n�"���ux��w�_�O�I������N����Ȓ*�!�JipP;�|�ԇ\�P���b]6�hƛQ���#��>����Ֆ��j��P�Ѱ�6$�v�y������������}�ԅm��t\њm�rhƫ���'i�+LD�w`ci�fN�P�%z�����Q��O�EмH#tVfh��dW�a��*�Z�.�����+x��tV������!o�v�{٨��o)���y��Ѹ蕴[B<׵�����&������E^�u���v��]y�}������FĒ*U���Znl-V�I[m[(f�Pϕr��f�6�z�b�k��v���n�$^Aw|k���������:-6bљ��%����h�,W����i*��r�U����H�r+l5�5c��ma��.t���B��0ì��t`����P�`ۤ�>I�ܭ5������������Uw��cW0�I$�G\�)|�6f�n�a[�/.�l��-q9}���DH�r?�>��o��[z�>�	���_���]�u�}zA��
��*Z�no�Ɉ�e�n;��Hx�SN��
�V�����������׾'&�F]���5@��ľȹո�!1��uf�)�	�ࣗ�E�8�BI��n�n�_-j���7W��v�b���}�Ӗ�����9_��B&"��	�H�"$�m��
��".q������r�S��'[!&���j3�>X[
�ގٻ��n�9�;�r�QWZ	��	�t�Gai��4v��q% $�Fܦ�+
c:(�b؛x��Ѿ4���Z�[$�$�&��
�K��VU���6�m�9���X��4	�Z�O�1��:d��,nǏ�Ty&	0I(3ݪ�2!�#kmh���ɫs��x�c�`�$�w2v̰c�&���>0[n�<�ѝ�WX�����os��ӹ��b��oͶ�o.�����.�6tiW�i�G�n���5M5r=9���<�|;��G���p�}�V�2,�/g������?H�$�XK�u��bnՉL1�*�A��֩����������N%���Xhmݯ��� �h�4scF�1����axv�cuj���y���"�
���z����s�d�ۦ�����ȟfk=��i�v��������U�T�&l�h��>�a7rVث�sBv��ţ٘�@�(g��֧p͞���C���J��v{l��|9���˿�VQњjg'[�^����(	0R�մ��uO&���q�խ����s{{q��4eU��Uy�6�7"A�sm/F���z���v�T2r`&y�Z�f۩��u�dN���3u�L���[�b.5��.��qM4^8,K�x�@�w��Ớ�w��j��N�k�j�P�gL���RHN�]@���>Q��r]��7a��N����7���۝���3���f�:*��*Ji�ƭ�3,#��)�n��:�σ@�Ŝ�ku���"�乼Mmh��OM����G�8����l6�n\v��Yv3u��hm]���fl��ӴfK�m� �u����c�6�-�������c�:q��KY ��ЏAA��ef+������ub;J�^���M�cXZ�f,��X*T�L*b�VJ��u�Y��'�UQo�.i�^0��`ݞ�z*�B]����u�;Y�;m<�)�)o
�p�y&�+(F��51�/+�FI���/ay����H�@	#�G��p��
�S������>�̈�U(�٢�z��k�Am،9.�S{b���$^�1 ����,7�#>�:���Xڶ�Ӟ�ŵ����`$��6�[cP4�����#gh�/9�3#@��X�nl�Z&b�\�H�d��'l�@�.�\�[�uy
0���-ɪKj���I�bE�4�H}�>�p���$�o�َ��6�AWsy��W��vl%A�����o]!��|��j�?	���4X��e_���>�u����4h�^���Ir!~^�ظF��{X�3X���1�f��޹�kE|fwB��h���*5[z�^����\��v�T���gm�{-_:ã^޵[��>̭	7���r��l��;E�1wu}<@ć|�����o;PEƶt��g�`�$��S��]T�3#��.swj�w�\�{�{"���~����d��j������b٬H���ϖh���ҿ����g�^�#��ύ'��U��{�@$�$a+h�7�]��a���9R�sfF�Sxf�#����S��p)'R��,�\s�d�u��í���Ʉ\��GJjKVX��>I���-(I8ܻ3r�%��1�*�����\M��U�����%�$��$Yax�|�בwR�c6,�Vb�s;^Vh۷��d���Ԛ��m��R�:/H����E�I~@k�����8�P���N�̽��2a}X5��pM!�Xr��{[tiH]X�1�lhz��W�5z�����T����M��ɉ�k��v���v/��y�}��I��/H�X/�/�N�-����N�ܴf�n4��>	U5�����S9�J%��\\�o���q%#�/8)�J��	l�-���\�Q�v�����o�	H�e���I
��H_Q!y�&��OKy�컄Vm�f;���B�!��/&�5|���|>�����$��Jָ�S��D�f,}
���[�Ϋ�bD$^�>�7�_�훘���wݴf��Zf�_¦��L]��׫k��TUf���2N������E�e�v��59�8�S���NѺl�ݫn�G�"Q`��W�%q���o!����k��:*$���Y�$�}�|X,iǲ��^��Г�㌥2�6;��Q�;�ϭ���n-�����v�hM��y�b�7L�\o{�ګ��+3̫��E�h.�ך������y��#�I�9�U�����L�߹^���[����	�ē�ԕ�(�5|�n#���1ƝUU?畤�n�V�]� �kc�&��\�D*e	�"m�կ���o$���z��ؽ`��l�b�h�yF��O�mxI�zD=X�ҟ�}˳���ڃ�ٻW��J�x���b����T���A\����os��	0	-���:'`��)5yoU',C$پ�&e��`��Ս@���1�)��L�$͗����ef-�e�� %4>�2ng�
�I��I=~21"ٽMUf��
[�*�gn'[E��ϗ�f���V��O��7��1�^�]Z��U��*��OB�O2�x�H1�4p�{F�r��Ҫ�P��S3���{n�FohY�9&
�Y��I�Km�������َ�K3J\6Ӎ�ơ���\X��BVސ���hnm�v���ݲh�3��J�[�ɶ4{c��t��� �{[�eu��R�ń���\,��0�v��7a���F�cY�g(s���n|�p���^�l�`��.�����/�Ul%ӭ����\{+:7"��� �Ac��[R�Ц��B4W�	�]T�\n�W �Ӽ�}~o���T�TM�x��H����qCuRm<hn���nWSB��UH�,5�����ؤ^�=����.��)d]�b�],�*��d���fB���(��$w��i��f�d�V�f-�e��W�q���*dN`�oU��Na�7���!�c�cn5kͶ1�w��ٚު�*��$!���a�m�o�aZ}�Q�����l�}�� �����Ƕ�)�KI%��������b���['�`��en߄�<C�h���^�I� m7�ER6���Մ�kY*t�Ʋ�-�l�B^�?]K�g�D$A�m�k���t^�v�0�5�_����>Ϙ�zD����}]�նL�;쩶��Q��=�]�oI�H��dC�0�`�R�UdΘq4¦�S��T"����vWC��\��xcB�R2j��is��ak/,5��#m4=[���O�..��N�����ŀ�0��v����1i��	jRr����t��$���9���ٙ�tG��e�X�a��\8Ѣ�>]�e��0R��9y���h�A�v�"�o�n���
x�&_�n�e[�s��hi���MbD=%VvUf���޽?O�`�7�XE�xqP��l�:�.�*j�M�1+�(A�L8R�!�¢��$bC��&����~<³/E��;&l&�	5[�RlbF��-�l��M�{>x���p�N��������	 �֩A�%6���5��kZ�ִ6i��9i�]��۷n��r����g����!/�T�X����'ݬ`"�2�]��*iM�Ne�t�u2�4�^�ʉ�u��Э%Bs��5�Y�ۥ�[���jJ�9k���s,�8��P��Z���s��e�\j5oSU]Yg*�^����|�܋U*&��MÌ����V㴔"�E�9�<�f�҂{��:�P���я��Ǭ�0NJTPJچ���Ú��3.�	���}p�ӯtV觖)ƥ�3o��� ��m�]�;;�^듯9�O��Uؔ`������{r�3��r5J�"��+�)���ٷM�R��]��7o�k�٥v�vvg^�֦g�*��,n���Uo��2��[{�gVpX�4�]o\�c��7u �A[��6�����R�[W�WC(��cwL����=�������]���{�4�u+ut��+F���v,��܎^Y�%M��Ɏ��8���ڂ��Ws�V�9�;�WWt��+�ow��Y���{��p�/0ݝ*�4Ys!.p7uv��0��.�G[US���c��+5��N��q��4�Wӣ�u�5�K���p�[gV�vH��bp&�<���M�"aɍ�"�K3d�v�����U	FR2�X:b�N��Y�<^e�V�X��z������뛣s�.�����q�EvV�U��aو=aor�Պ;er��Gw8''����2�n�)�$�kY������8u��H����[��h���-Z<�{}ys���{W�Sq^^[�6�Uk[֚!�m#�7r��nVC�2�8��n��*����[��s�������F-�Z�Z��2F(�*�6K`��X���M���Qb�4Q]w��0m�œ,m��4sW,yt�Ѵ[r����湱s���s2ܓn�ܷwU��Ԇ*�r�Z1\ۑ\��%Ȯ��.멣sN�˥.�r��k��#S����+�����+�i��_^��x�r��u�afnm�ιA�V(iE|9�IOKsR��/'t���s!�jSnk�nN�S6��nRn˻�9n�%Lآ4��k�t��wZ�b[�]��;vĦ4��5�U�=uy�.ni;9����U�ᷛ^�h�c�X�\ֹ��n� VXl��S��hi�'[�"�� �,��{�ہwo��2�}j�6��0D�F�Ǡz���/Na�};�Vv�q��|+m=[|�������y����㺃f�ux|��`�z��UN&�z��1�ي�6�k�j`�s��P>�g�ܒSj���B�����D��4O����D�@���gX,
[	\h��ٮ��a��O�x�޾y���YO�&凜���v��}fh���y�0m��=;uu� �� 8�rہwu�6\]gl�3I�|��;"<E����/q����p����A��O$��9�`"�C*:�������>�n�D�P 6\�l��m�k[!�MO"Z*ս��4�1[����q�s��w=fϮ��5(%i~���]K�y� ���� ���m�њ�nj�ő���@�`�P �?�Ƅ��[5�*����TT�B��&��Xc�#v�\���)�ݺ�����\z��3u_<��%�
3[h!��W�$�����ÀF�РN�,��#7P����pz�������F��m��1��᭤y&���
�=Z�lΨdL��!D;9 f�df@��p�rJu��մ��Yt�Yi�ʓ���	a�`��^��@Å�A�p�Wם9�1�My޽��x�M����g<A�p��n�G�����m �n���X�ͫ�!�� �3��x�ǫ7a���zg;�`|R`��6�=f��c��u���p��΁ ����b�|`����6=�lGښ��kfk��7����s0����'���{�O�ڈ ڷ�7�����sQ�XY��A���7n�#�m󶞃Ls)�;�:��Q�|*�{4]�8"�b<Si�g �.���6}v�N���[D�� �������u]g:�a�A���>�v�x�-��S����͸*j�	���0s�#[=VJ)ޭ�8#|z�nf���.��p�5��1sۓy��\W�5TZ5�Kέ�e����>xZt]6�)�1c��#��u��>[�vx:	��{<��hh�:5�^�A���e�zwf\;$d���mL��˛toj�K�nu�D�Rnm5�D�j%%�֖[4���A���v��`�M�s�fj� �:��%��F㬝,m����\�	����a*A�*��u�,���hs�ј�x��G6S��VK�Hn�3>�U�UAR��0�r
����hJ���nMe0R�ٛ��b}���=�� A����w G���︑�}�5݌Ƴ��{^C3�3��z�����ǵ0A;���qwP���b����a�>y}i��"ym�����~4�� 9����=`����=��3�ܘ�~t|դ?��㻬	��h�"�N� �S&�ש{��.����� ���	8p� ��E��xNa\�����<(AJ>�f�G}�U���p����쩨��f3������||ɢ�||���:#N����@?��6@�[�-���N��Z�ͧ��2q�8zoz�>s�wn=fχUY+q�}����S���<�k�;������k����n�����z��M��~a���}}'��A��~�7v�̶񶥮'��gx9�omw�b&j�;!�2�H:t� ���dM��Dn�������_�X�Rʰ�7c�v'cb�#�m���x'+֊ܙ������$%M����f+�5w&.,��=0��O'�aO�Wg�fT���g;q�|@�׀A���ݰ/s�U�0�ӯ}��~�{�whQl��v�Ӹ*L���{�s�θ�d�t8���޺�Ec8�p����@lݰ��ŉ~z�[�A6���V���-����[�����3,�lp]�p|4B?�/j�ng����Ñwq �.��E�wo��ձ�,y�Cx8iͻ0����n7y����A�`�[���`�S����I����TMy:@�fw��Q��M�-n�v��kfx4�HN;���0ObD�g�
n��_�_�
��Mq���̶��F-
�Nd��6:td���"A���U�� n�AwX���[2�o+2[ښ�����wA[�u��fY��o��������	��l_V:���^�k����C�1յ�=��8 C�f�\�Û���S�eDC�����Ʈ�`i_וS�:���ݾ�����k8�q.o:Y�|�	�,Z��d�L�Q�����9+憉��c1��������C�v�A���n��6�s�b��OB�N�AR�<l����|F�x'#-�u� �p�����2�c3��nxi���l���ر���8C��1�꒍WX��8)v���+�֋��f�����7m�8�B��^���H�84��]~�,Zj��qn&�h�4��(��X��t��`�9�Y�:䃃bs���1���k��v���Ym���J�8����U;���1�����_;#�^g�ɂ	��^>��}��¥�wn.4T����S�)�����|o�o1x8ӗ�E����`79\�wo�0�/f'`��[���g@�י�.���A���"���b*"�{��LaW�}cy����l��n��wX~#w_�<������]3|a�(*�?�����z��he��^%p�-�[� ��n��>SWd#�<uCUPnʱ�����bt<җif7��+�k����k�{~]F��c���\�[T;(sTU䕮�wM�����6��1�P�2d��{�{�\�>?}�붣�N�3�ۮ����{3�����<��~�=�VFw�WB��[ ��B����=5�uvp�8�S�X�Y��@��q���]V}��q@�.4�f�%���7T&�-�U#c�=���#�^`�'w]�㷬b�Lq��[��9�<�=�Yhq^+?m
� �u���Р|wPs��	�񯧮T��6�#z�<����G/N��aw����u�Gk���`1f�]�TR��ù��� ���רa�����Yt�?��~�ʩ�W.3}��q��� ��z]�@��v���rS�l�����r	��#��޴6�`��M���7��H��2A�s�Ǣ�o�?�C���܃ ���F��n�ƎǺf褰{EC���i����Up��׭Ƽ[Ǻ�;_�@�g�>�� ����#��5��a������К<�OK;��ݾ����ܣ]�#���ۼ����ж�#Vv:]"��P�Q6���,2��%�턘X�*=���������v]?��LDJd��Ѧ*���a2d�f�n�6�lfa��\\[!�G�^�d�mq���8.�չyֹ�2�3鷯���|x�[.�j����sHf�2�a�ZW� {8<v�
�d�]a��X��ˣR��!��3ZU0u��爖bV�k���ʍ��*����!F�B:��0'�X�1�d�ݣ+���Tq۲�nD��zC5��u+���A������a�	m0C���c��:�:Y�8u�Ń�\JC�e7�k\�_ٽ�����<@�`�v������7��Cc�\g{6��1��*Km%L(���\z�����fc�>)���pל�T�U۾�X��3�����o8#o@ ]��o�����; 8#z�@ �pE�>w��f8�Jݦܜ���gE��� �JW�m�x��x2#�[�rx�m!�휂ݼf�/��ѝo���ho��|�(���>�a�[M����3�=U�w�k��>՗���㒗��"�#���������ǳ�0���$�ox4.!�,`1p��a�vZ���o89��� �6�< ���n��R��~�ƾ����U")gE�7D`n�i+���,����d3�ᛈ�6�h�÷P!��
.#����=�j��6��_h`�\��ȍ�a���7�y�3^H:��`�L�<wu�N�@���g�����2�#_���5�ŭ*(`Ƨ��WSPզFQX��2����EƱƎ�tHU���r�.��l]��2����T��I��QC�X�t�Kj�r�!�����ܮ�=�ؾ(��ͮ6Qr����>�{��w��L�j`�s�׈6�|v���p5Y�c�2/�}.�B�2���ps�x�8�vl�H8p���<Eݨ����鍾ۍ��A�x�o\G��C���-�EW|1�[��0`y�� �f�騨"�1���] F�hwPd���^:t���ʣ
�*2 
P�+���7�X���r%9�͞�M�\�z��q�g�c9�:�RZ��Y�oԛt�"HeW�.��9�7�s��[3g�K��jKA����bʟ���ߞzu�����n��;�V�u����;������;����c�>���#wj�N��<
�$n�{�իHT�[���v��ߖ�	�׃�y��[߻�jAs�p~?}μFhj�`�.�6\n��x��	�m���;Da��Ěkx�\�ug�5�ܗJxh�5vEζ�2��"=��+a���jp�N���i�<�\�mų��� ��{}�M}67x3��O�����A���}��Ȼ��x�k>�o*94)�[Z��d#����x���MC�{~���x7�9�����l��ye�p��6l���޻���X��}���ŗ+��!��}ṹ���wq|�m���c��>휂n���&u�}��2D?Z4�(*N�R
�S�V:�i��3�P\¹IF�[����_��>������Y�C��*u���%�FE'��F���fid{��^`!���Ox�Ơ|	�ǀ��n����F��H|ɟF�����zy�t�[���˽��s�^0���6@���N4<.d����9��=���Eۇ�w�-��Fo*UU����ң�������އ~S{�V?�[sv� �p#�Y���_���y�w@�6\��v�[V��wq,&��6�;��>���r�6��F(w�D�F�S0�O*��3��hW��|6���_�9CjH���
���O��ݼ�{CU�mO�Tpp�}~{��g9�نz��0�-Ջ�n	�V���Y�v�3�MYϤ^�to�>���n���tBv��y�|���x�8��ua����s��~6?ɦ�*��(�[�À͡Uȑiu�k�-4t��)ʏVf9�|ƈ�O3�39�x�v��Y[�Eu����c��n�b�;�I�����w�s=���s1��z탃v��P�(��X�;��>�[V�b�y����[g{6\M��c�wo��ój�t�ԃ o��~�@����7v�=�k�]C�m4pU�_y/4y�p|oy ]���ß����ѽ#b���r�9��&|Nc�މ��wu�7��'1<�n7NY�������=��;�7v����i�n�1M�P�x�����{�ݼ��e���{6z<	���wpx���3��OOg9v�����M4�ӗ-4�ϳ��������4��R?��ר�'2��Z���]i����i���k:qX��޾��܊����}��:|�gWeN'k�u�̄���ʺ5s��m�4k��p��덆qvk�a�lj}cDd��
���jN��r���h��M������j����k�+"���EڼJ��v=W�{'r��f���ꡚ�a�|��2*�Ĕo�Y0M�{����o	�2��Cf6�1��#��%�+�[���]`��#|��=O3��f=Vw"�17��qާ^��{Z-�9��L��ͮ�J��t�%&��`ԟV��2��~ʕ}��wF����\�
�]u��Zԙ�4k+v[�b�#��3��]�7�lZ�{)��Ļ����f�u�6qW�����$r T۹�a�����1-\^_aL>��K�{��.�sr�un��U�r��r�5�4�0>��ݷ\��J̺m:yc^�F�wR;2+2
DږPYT��=%����d��9X�u����-6�87)2���ʥ� xQ<pQYp�uw��]��y��D�i����ŕ�n�R��C�ŝW���[�+*�Q�����p���[Y������p��ee₆e�;��1���j��SWʑ�L=��wwe��~�1紎s�T�hv�U��wY�����}�p��L�^丳��݋�<h-3*�r���aD�����p����Z�]v�J`TFw[÷��ei/�d�:�X�ne�����H94�6"����m�V]R��Ye_oG�L�wv�2��n_�,�K����	;�x���[�{&��FW�),��]�m�[��*�
^F�ԟm����m�l[����E��
/�ǻXŢű��Tmsk��X�cQ��^[yh�E�h�̨�*66ѹ���y�V4�UFѴU���Q����f�k�lm�Z/�ymyRV��j�X�lTlU���5F��5�6�5�WٵnUFՈ�AdE$E$R�����q���/ih�M=�xi<�j"ͦm���0��uQj��d^S�m(������qųn��N)��b����t��`t ap�3m%Y�����l��l�V��G�m�F�n���6M0�l�p�v�ɻs��X�y��*:�p���:�R�{!�]��3B�CGD�PŹ��	pף��nS I���^[q������w9V	��A]��Z��m\�i�<C��>|1�"\,t,�ėVMnķ��df�ID�k�� ��mb���v�O���� �m,�����K����'V�&�spChei0��aˎը��:�oMg���h��qۮ�\VB΃�y����·�n@ݹ�{�[�d��I����7-�4ڶ}z9�J�uv�h��t`�po/Vo-�ma]Y�X�u��lU�b�6��Ʈ���[<&��C�nc%�&��1����w���j�pc6-fav� ��H�Ʀ
;F3�׌�i�6���k[P5�1���]��,k��U�<bC�g�ܘ�aA�Y��
6h#��D�h�3孊�҇&:�nK%��Lf%���JiY5ĳ:1�[`Z�ls�]u�ۮ�rIq�tF�YJ��惭��1¦�J�B5��i�ZD3x*�v��a�u��-�v,b9�c��t�$��r#�v�ri��:�\흸;'m;]z&4H�c#θ���U�y�!+��e��+u���K
�6B&��oWD�������;��Nc�����Pq>l^}v�<���)�C��wO��'m��n���������=kv���6^V����6b+�+lXs�ENͨ])6�x��Ql�]S�y��e�������,��/��c�,|u��b���;�.�6�5q��`ae�n��!Xf
�y��k�����{�Sv��%�i ��a�lM(�a���V���n�����-�N: �,3�;hЛ��LP�G#Xz C���7k%�\�5��溶�U��P񪘰<���n�[��q�{qӵM(ݦ5=By�7�f�#�duRQ�k��f����ӻ�9��/��u����88��b��=�YT��C��@Y��/3S���u�.wl<�=b��v՞z�s�1�����es�g�hKGJB�B/�n��ɹ�K�M��I������(��d�z�.���mƋZ��wau��A��nd����cRu�q��jø�^j���T]�RD�i�����R��͛J�G��1x��3ZSl��=�>���A��x.�w�vM�s��S�%�P ���v���hpW6��MQ;ߐμ����H �wu�޾�{j�y/7Ϝ��٢��Ól7���Grd����+���ºr�/�V���@�k�ۢtu]��hM�m�����
7l�A�"�>��9-�Og� �{w_������%&��rr�5uƔ3/�e�n�o�e���D}�����^>դ0wS>���r�ӽ�E6���Mݼg.{�O��E��p�[��%E�A�n.�x�C���u�F���,�Vۇ]�����^�zD�YσVֶ��MwwZh����A�C��x��/xCry�ZX#*����Ÿe㈞I�b3pF۞�[����i@k"[���'���}�����/���>�e"�?][m��v癇����� O%������U�G�!����9�G٘�A�<w�k6��~�\��T]~��I��,�z12�gT�]�񳄘��l�f�k����(��������a k�:�V�εo�EP���n\�J��BJ�k�Y�g�٨�1!��O��a���ρ�xv�oT��*[pra"f���pA�ۇ>w �a1-����a�Bn�(e5��pM؛� ��c�����v�8 �wn�))g��ɋ�`/�J �j ݸ~�c�4�?<��!y�|�qlop�Q�r�����d�z<A�`�휂n����� Ƒ�&Y�c9�q�����%_�o6��L�{�y����"�
ݏ{�{���0���'+��"� �&;6A�'O�s��6p�Rn#
�	�5�ҐƸ ߾���p����E����md?�U���(ڻ�	�q��h���<���y��q����E�p޻`��y�[�p�Z*�֎N� ��}��vֈդ��L�B�`��s��6_��Ffc��]�1��9��~3S ����t�wSۺ��yw�ܗ-]NP�g�zCݳeEf����oT�A�7����õ}�UeWR��ӆ:��A��j�oO{��u���;{���S��舜�/�� �j�C:z�Ļ_ϼ�'-��v�v��m�<n�Uvj�Y١\�{Θ�`G��;�V6��"*���:����x"|3o(�<Z(�� �l��&��	3�J!��&�Z,s)���'�ݼ4���53
M��6:L���r�w_����7_�����9I�N���%�̯��	�u�x7�˥e�M��P���B�:n���~�A;T�4J����p%]�]�/'kQ����y��������#�Y� �����An��En�Gu3v/�f?�x%���� �cgOr"��I��!�7��<��n?��m�K�,��ў=�> �R`�R$�|AI�v[/پq[�ɞFs.��	��S0��~�?���A���������yw*#��58�n*̶����?��L㫯�Fmj1��/8>7b`���; �nNL�T���M���.������ܰ�Rz�tm�eSى�8�_	ƚ�-9����J��h���R�=����{}��n��V���m��;���ئk�!�+�0pR`�$��	aI|c�ܛ��]���܈�}i;uc{������\)X"��d6o����D|��T��8�n7�t\H.�jznl�6��q�<��Ɨ���>;h0D��20��{�&;�L����c�z瀄sC�6������@w�c�zď��-�@�u0AR�9��/�'}&����k8���ћZ���G���q0���)0�{H�E�0E�v �H��!~2?n@x�Grg3�����{i;r�)�����dL�dL���ǃ�u���!^�T��0�=M�u�3G�i�9��~pAT��_�wu�Ym��7�r�x���0 ȼ�~fE �#%H(I��3�U��n#�g9�`|@��?�8(���N+�y�0N�}m��\e�v\���AS���]Y��k�[�X�$L�]��%��S��X��7��]��������+��g�Yz�����w�� ��*�\������-�[�y"h�T]p\X�Nv�n����6H��F��]��';v[������`���&Uv����|Q�^7g �F0�R�Iɵ���I3����6�6#�0�us��;l@IW�rd1>q��̼��a3cv)s���f'o%vy�l���$�K+]����sid:�I���k���7&���<�`���1�nƯ�ӯ���"銼˩4W�Q����d�'ε��5���}nL��j����X])��F|��`�r�$����G2u����'nX��E0��h�Gy�cc9r�}�_��L�c�"��+��k*3�Ϝ�"��oI��*�Ng{���8Yw�2$����!T�'�mqT���!'���M���[U�
��E 
�W4^��[���w����An�>�,ȃ~"F;P�������R��!'󋌣y:�ȊW�I�,n �M�ihE3-44;]��#�A��I��� ���L+ng��W�NѢk��Sۛ�1���3�x����m��s��ғ��l��>$L}�����z��:��#.�2�r�R�@�v֍2�1�6���e��1��/�Y�~���?����7����u'3��q1
�S���Du��j�`�`��A�<�u��F����y6�FasB���x*�W1\xՅ��N�n�!��93��3����Y�T�.ݕuo\��3��t(a^(��]V�h*Bcͱ�Ln�qw��ɳ�穙;(�h �{��	;����ch�K}�")ue!����r�&n��٢��so�Ľ~9Ȗ/H��@����&h�÷���c�	d�D[�VL����k�8�?�>��?#�F+ƌ��+���;��.&��g�ۼ'uV��z�9�6�R`��I;���pF�����|Dv0b�Dm�D>	dIb�M�g�/���yV�/�Ȋ���#�7��m��U�	7���ӧ5��\h�x�i�����b(�9I��X���b<���%�a�Dq��.\��a�f���[�)0r`��o{b9�"�D^w��8���vh1�̓�H1�0FE�adL�dL�Y�Fm]f�h@i3�G�M+3zN�2��o�9��Q�C��"�@�~�@�'�`O�`��L@��"@�2!^#ܻp�}m]��uUك%S��5i�I�?s��}���uݙ�dq��ź��*Z.V��
Y�2'qH�"��W�xx{ޯA�OR����ۚ�e���	�o$�A2&}#j�S�B�#=�@u+ ���yU��t�CdԨ����;x����Wm}J�F�E�y���I������ ��I��.2�Ec8[۲v��\����oJ`8�I���^'��ZS�g:sH�cU���Ś�\<D�m�Tb�l��;�Ք��*�) ����L_!���F����R`�U�(|���EGE��������[�,����؅x�L~Ax�ߝn���@_��[O�ei�D\L�����{u���*eC�w��8$jg �8r]��9c������|���dO��
Lb��wΡ�ۦ��Wf#.!��Ͽ��2��`"`�$`Ia����7���Gc^�^&Z���_gr"+��uk��o��K��Dd�,n�Idf�U4)L������"����#��/cNM�X�O>�;g��p|*�랾ڪ���Yyak�v�"���{��AQ%�c�絮��kog9�w9�r���.�E쇷�t#%Êt�c�ǭ��T=�{_���7�g8�����L.��sۿ���U׉ �"�2�D�%t�X�ҫ4�:��-�9+Y���|>��K����*��M^>L�k��;_V٘�{���8����&���0Gr`��#�`�y�U_*�ͤ���G<v���`�n�c�<wY]Ux�խ�F���	)5�c��;��+%o���>�l{�F&)8w��]�r%�5:�ئ]��{_������H߉���*;|ɪ��g>�ޭi�x��5x���l�s�\_y��T�G	R7���S�hr/ �0�6"Dρ�g�!�2P���7���������Ξ�"���GV�x�ܙ���^qY��b���i��
!�$��&�k.,V]#I��a��z)��6[���
ȅv1�DSEH��5��d��2�bk^K���Z���Ao�M��Z�%��ů0�G]��Vٵ���Þ9�]�����0x�5��O����M��A���/r\
�@a�KH���ٶ���f��ī��Р�icX�2�1����t� y�K��
��hĹ!�5�^T��e�*���3ve&��2�2��X�!����Cg�tb|dx⧍�M��ݰ�:�=lo�����<Ot�{����r�m�>�o�Ca��S�B���;J�u���1�cL]���n�6�^7Qgk�)tgJ`m�w��e��2Y}}c�{�2�p��3�4w[�\���{_��&�g[nw������Q��wP`șȘ�P��潦��X>�g�]���um��{����}o=6x�����Ȼf��ull-2�/�`IÈ�
L ���ݸpBN��&Ʊ��u��m�',����#�[��x�]�n��&�J\^�Y�g<3i��EK��	3�
Nn�Ǝ�|��{������C��c�*!��HŞ���to�عyd^~2&A ȃ��vm
;-sɟ0�,�qo{��H����'�1�/�{�^�t���X�	�lb�Gb���֍���o]j㋡s/4�ɫv����4���y�l���,I��nE���lv�̍�nN:�v=��Z���Lb�O�R`+�z����9!�JvMe������}�y��O����������v�"�*��B��2�l�
��JLX�RR��ke�s����=��*� �\�;n�!���c��]U�����7��~pN�.A�p�i�|�i�t��Y�A��I�pE$�A&��fM��CX�%�6e��7��>=���� Aȃ#�a��@��D�}X ^�>r����;%����Gs��(��Hn�L���ucv�����5�j����֢8W�E@�r`�:פ@D�
(��-�&ʱ[�S�.��+���1y�[q�e��`�]�����4w�l�@�g�o3ApCH" �Ge�=��X�Xq������ˣ�7v�o���~�o���ϒoII�ku�x�և�~�o|�9ma�v��1�Ϙg.���Qߘ&|Ž��]�YøQ�?C�~�r����E^N������	���Mh�V�8��#��}\��5l����g9�q:zzzv����v��M;v�ק���z�^�W�Z�u9N �'bPR��o:F�Ή��7��	2�������̒��moS��**���v�)p`����.�����Qζ�ZQ�M�zb�}|�ZY.JwG���s���M�l�YҠ�U�̕��6�n,�{J��XݓٕGM9�/T��b�nva�{*�R�;�vJ�{�Gu�
X���R�����חur��1�LEj�~wk2�83i��J���M"��g����.�ǻb��ۍe��2��첏v��x��:���ܓ���q�8�hݘ����ʸ�K/�vB�8��*�S(T�̎��豃)f�xj�ՖF��3jePC�m]f�A�UGv�&��p`�v�m�{��p[f�u���w��oK����L�������v��pL�t
���c���\���ǻ����5M�K���b� ��uB��-��η�)[�Ўj�s[g.�a�!�Z����|u굚�r}���7p�K�j����gtZ�p��uX�ˈwV�|^�ͮw�dفދ���YI���A�
VXx)m��37h:�ˍ���;cwW��@ڥ�e����%_
�,�t�����LT=.�e��՘�j�h֌S&
&G;�·0��K�Lڭ!Ue�op�+�E���{�f�w^�n��u�!�}LIQBO�i�V�L�xŧMǼ�v��޾F�9���Wt$&{�|6jc#X�ݨ�Ͱ�r탖�!̙ɞ���:���83v�)�O�w`O;^�3f�n	�=��P]���C�T
�&�n	�rvN�y%�*�qhd�0ö��4��x7�4B>��S@p ��Ԗƶ4U�To�k�ѭت���5&�h�j�h�-TlVƋElb��WۻTEZ�Mk����Z�lY5�֣FH�XՍh6�k4k_.�66�MQ����Mh�E�F-�X֨�Ze�m�m��V��EZ��-���Z(�-S���H��*�{�}�x=��}�x�˙�,���8 ��r�o@�.�|}v����;c���a�  ��u3�$ҳ]���`{�~X׾�������1쉨u�����0�6�����I;O5w��M� ���Wv�a�rOy69[p>ݯ<x�c휂n�F�[�r9ˌhbۿVߛ�n�1G��k�˝�F8m��wcG��Ea�CTi�ٱ�~7���~�~�ZN_�;wa?CS�������k%�j����F�A��dta��` �bg"U]����Z*/Q����'e�v;�sed��~w�L�&�c�~��L����R�K �`��B��Z�$��RFi��p�3����"� �'�-!��2&D0���j�����Y��8[����fv��)�����{g������a#��m�.0*��0��S�"��/�a�� ���Ny�v�g*.��7�����Ҏ���S)-f���+Ga�u"Ġ�&����_�Zbobo�)�Id��	�VD�BFAo���+�7���ɜ���y�O�)3�>źK>^�c���=/e�]����j�9^8r���3Ll.���Sn�hg�C���\�N)��l]j�۫z�X'������[vO��=��k�9qÎ��]���ݭ�M}6*�ϲ/>�of^/~���㚼̉�"d" ��l�����ѝ��������7wb�1K�h#k��e�w8pBK�A]׮%�xǁ�o<��[�!8	4�	I�8�<^k���A6r,+��"��n�l�x��I��
N6>�Ԃ;�(�� "�FF�?����F��/̮�Bn��[9
��Z���-\C~���L�$�p&�	8�L��kb��~n��#wp�h�\���z��l�5�������z<G���b;?/�~�)���[q�u�ǕF�y���/"�욮;՛��Y��}/~/�����I��Bo-��v���"��}��GD�~ ���l�3fZib�o�O_�����bz�T���.a��Lk
B�e�	Y����];��cv�At�bzp'(�ym�9#v�EV�J�-f���Ytl@�mu�GK)��7B���0�b\��:^)�w ۓ��ť�R�bZ��(�$K
�,�	HA�iQ�k�0�Yi+e�y;]v�&�(݃�]s���	��n�!�,���*�+(m�@
��,Xm綝�$xE �30?��0j��-�����m��.-��v����Z�B�6�]~���/K8 ���8��,־�cWDC����("v�؊�ʶk�)0r`�!&
L��~��z뺾�p�9���6�3w���Ŋ����A-�����tb츕���g{�I����I��Ek>�δ5����5l���)���Rg�-�gO㯣��~�jEG��wS ���#�M��/��Y|6[��6������<�ڳ�|m�g����	0r��'J�c��K=��G���s�f�?����i���A�[��L���}��}����3�奔����չ���GB�����l�+�s���Ê��S#�I���e��L`�C�V���tx]`|�\���evFs����Y`�#9������W� �o!��a�p����u��k-�4�.VE���S�*����FsWc����i�c�Dںf���D��)�.��Yt�.����R���I�7�g��λDX�a�	D�� U�M��3�Ŵ���f�z�v���A���fD柛ׂ��c�6yA�	-��#�v�uݓT�a�Am.��Wӡ���Y�4��	�O�l^`�1�H�ǅ�&X�V��2�8�o
��|�缓Z��k�)���D���!k���pk��`@?0dO��u�pP90��o��5;�����u���`�>^?x�;�2�0X;�NiϬ���h+�T�4�3�00\�\�qi�ٸ�zL��t�Qz�u���a�����c�]����V�U׫c�2k��4�F\7`���4�)����>)7�R�I���5�a�O`�g���p�2'v3d���͝�pA�E�A��m�0��V��LP�v&A��&JL|G���,��i���n�
�(ލsMff���X��!���kHmJ�����΍�Ȇ����U-�}T5�tte0��-�ݟ��O�$�A ���^�s��_g��w��;����"F�f�i�a�A��V!�|�X1<��~��vԲr��7M�z_�Af���l�$�󂹜�p���^E��Qz�z���s�ƅ��{��E�5�&l�\��A�E�����dD�V��P�ǌ��0X�0<�2Ok���Qn�3Q��]���E�󾿅�3���͇�4�)3����^&��C>,�'Hִ���ß�����Ak����$�$�J(�"�k�6��1*���.�:�?���js�+����u���q��l�r�(����ߓ�a�m�r ˆL��ȣ�r����bRg�N}00�b�z�Z�]��h~ Å�}�0ȑ���fD�v����藥o��a���$�-FwFDMt�h|��GH�_��z�v&�r�x�ECb�M/+`ƶ�8�&f��:s(|����/
�2�!�7N�<���D�r��<(�� O��"	!$`��1����m�ja�]�]���0L0�"�~"J���V,�����|>Q�/�i���.�Rn��pAI��&�;;���.ǲ��]
pS[�s~]!\,!�]��ƪّ�!/]�v�ܜ�k*�n�b�L~�����A������$A�\�\�ѥ\N&l�\�|��E���Y������;������y�I���9G9��z]�w��g �sG��S�ѱ3]�Zr+8V��L��Ra71��爧Sׂ��8#�Ã���I�I�>A��ܻ��DH���W����k:��� ���u�� �������z�?��	�{�ⵃ�.�<d��ʝ���f���*�8"\��:�t�85�7�~��@��μ�^�-?"�Rȣ2'�n�+��p�[�ƌS���[��cVp�n>I��o$�
N+�zQ����>��<��6X|yFZ��f�����8�S6�8Uڥt�]7��6�P�7��1��������c��e,6A͟n��C1�X$�a���(��eg�Ł���=eЋ��۶�氄Y]��X�.�Ȋ�N��iR�мhӚ]�攀��4[XW��,#2[��1]-R����CKe�m]������é��<�Axx��'n�݊�����Rj2'SBPK�YD��]	����ɹ�y�h�;�1u��\n�h�cs�/�˞yh���`�=v���wh7E��ݥ�`�^o^Z�|����,����.�u�@Y@ؙ� ����Z�Ϋ�i�n.�1+~���A7L{�`v�p.������{�*�:��k:��kJ�f�f8�$Rg!%��AH��z,� �#�a�\��K��l�|ny����A��!!���(��1���{����p���L��E�O���c�:����f���V�|Rl��y��L�'�.�����C�U�mt�|�hf�0�Ñ���);�#Drս�U��,�Y���U3��}����A9�ay	�@ȅ"��/u�7Wgg*\?�)��ʝ���K�{o���/W�o�0D����pK���츿~��6L��hPj� �f��(,Vh�FP�%%��,���M`RSg�t�u#.��~�c�e���3��
L�ԙ�W&�v���k(U�nt�K\��9�!D��3� �"F�'�&��d��2�{��&��qRh�њ��n��9���fS_aմ)����]��nfun�!����ԧE3���6�ETT�\y�������>>���|Fӿ���~s˳~ت�P�ͬ��})�����M[S6�{��.;�`+�d\@g�/�y��Y�˝�� �<��T���l�B�?�0���BM�	8	4�W@�#Yڅy3�O�0�9�g�@�;��lj�8�U�nV�ρ�v��a��r��>�a�#"���n}6��tM]Y�S�/�c[�ۑU�a)��ܶ��r���Ș �"ڳ\k�����-��	��+���d�(lat�u�˓��j��iP�յr"�����	�`���R`$���VfN��\��f�@�n' �Ք��o1�������� ���Y��k����F�։co�>���b�W�ⵀ�a��&64���'��7`8 � �F0�"�x�Z��a�wW��f�
Y���t��sY����ŭ�.�>ٗ�\['�=���f�9�&ڽ`�Y�S:���]rm���_� z��@�%wnw�3���s{�����3X4�JL�$�ٱ��r�S��L�p�|�'�w1�G��f[�<��(�=�Tɯz;��ZO��"#���8)3��&p>L�r�C=;��_^���^!ٶv:ݱP��p��/9EH���i���%�PTP)�t)J�`��Z��rM�2k���,�#�@�k4�3�>�_��a��ܿ���d���x��e'W�"�h�W�����A��)��d"��a$F��������6<x� ��93���z�[��B��E�"�Ñ&����~�z�w�R��/�`��2P�@�"�_8��πF����n�s]bl�>3��Pdo/C�}�dH��<�M��,���~~"(C��{o{�@�):�䛈>=l�?��J+6X|qV�y����W�-zK�q�{�V��+��/o.Z���]�hfp" �л�h�/v����	k�ǜ<<�G�'�	��"CDd~�;�������S����âَY]��Q���Âw�	�B�3��u��0&`��I�Q�	�n���Y�hy�ck�j���Wg����	�g �6��&r	I�����ۑ��X�>�!L��n!`�=�B�Fϟ�n���(��V��[��S��� ��p�,-��#��vs�����p>\�A�C���q����c-�KD��q�{~A�7P`� �#�MGlc��M��g.pt[1�WyCzv���HߌP�����::���/���kQq7���6o�.-����!b�po]�+mJ.���-`����9�`�a���a�$��ර�R��;�p�8�[g���p��frM�z�xs5��ׄfshΞ�zp�M7zv�۷M;v�M<�����n(�&w9޵yx�
�ۺ�v��Op�y{�
&��E֑f�x�HU������r�wZip[����R���U���]=�.;���(e�r��d}u^�<�	��e��j��!Ω��He��|�P�
�q�p�b�&��ofB�iۥ�]<鯅Uq'-��1V��{)�VI5m��Rg����F��u2ݎ�>��Q:�_r���J������ڭ�t�KN��W�F��S���7^v��v�K�F.�K�G�v�[�ޗ��5�Wt�|q��|}R���z+$7o��Uά�t��պ}�:����m�m%�e>�ݻ��V*���;uX��3�i]����B�P�v���c�'��Yj�\)��v�V9��H��#v��*�;z�)֪v�BZ�V�F#�)��ѢhPN�`*�WnF2�D�v��\杺:���0�f�f}�1�k��U^���0��W�:��JA�)�I}��aX�Pf�u�ժ��4�s���*���Ʉӱwc��lJ���(5��]�m]��Ues{�ݝ����C+o%f,o����q�ㅒN[�옍\�n��r�8�n����-.鮫�f�u�@�z�����qo�U�p��k k/�	'k�;�vn@�8�M�P!��j�ɉRʜ+�n1���T��;ĩ��-
�Gpܫ��L҂�X�_!i�toI7�<�Ob5��V蹣��ѷ�*p�u��� r`�ѩ�F<�KԪ�����%��L������¥O�vm�t~�K�Ψ��y�_�A2���%���N��^վ�i,X�6�bը�X��毕��[Eѭ(� ���h��)"�(����m�*�̪�sjŪ�BEH[Esm/�E/g���c���O]"��y5�(�nD^341c#�m��y�o���,��i.�ц]�:�EE]������[='d'tv
'r�q��b�-:�օ�A0�f&�a� `�s`�77:m�mp����v�n�-�,FTft�b:%v�Ѵ31���\������]0d��WZٶz�>8�u�{l];�'BW%fq.�lE�sf&���[P����\<re+���^#%��w:丮��Q�-jN���e�4<�����������7P;Stk���Ȉ�Gl�u�F&���2� �7CT�a���]M|�s۰��ثwk�v���:<,��!۞6���`�l�wVaqSv�-cX32��,��)L��t�K�.�ņ4^b��jp:��yKm�y�4�<R���)stL�읍c�����y#�:��:ŋS�&�0�vFa�ݺ�X��7R2Rn��tu��WlZB�	�b7T��PNv��@4���ٲ���b�^�,ōJ�v�M-t!�
�����)�.7��\8��q���q&�Վi�t�Ӳ�s�����sׅ0��F�f�l�`�ͳ��(+ǰ�8�#�q	�)��5b-GC�¼ M�G=���js�G����I��Y0�"z�m�WF0�6-�Y�:uZEaf�������4#F�Xl�ʚ��8�#Sz�Ɨ���Ő1�%�f��C�O��x˛7Y嵴j-��פ.��=��yī�s���5��av�U�me�7N�wC�2qA�tql	��H(A�Ql��� ��r�Y8�
m]�`�@���5]���q5�!c���|&��g��O[tYħ1���^ۘ좐C��m[���q�'F��J/	��+λ��v�ە����a6�bl��۵WR	4͆H�nCm�b[L�l���V��t����u��]�ܺ�F.��緕�n�N�B�J$��uۜ��� R��;l�9�����:���t���2�5L<܃Ҁe��q�m;�C[i8�°��j���iw������z���޼�>����T҉�%56���Z:�c�-X�gt��8�y��Gj�ۜN79�d�A��dNu��78Ҏ#ps�Xc0���6��sR v�Aaf����r��"!e�E3�]��%�]+��wg������s���2�E�TN���t�k�k���Վ���`p�-9������0�,�2u&#v+ڻ%x��(Mw�CE"僖H4���E�JWB�9�.6iQ�A�C���d��<��uų��� �?��9��>r1}_[<�7�[��k|�N����w��<�u�Ž�a�����;���!�dC�Ș!̓v�0�5Fz�k_��Z3.-��l�!bѩ�������&*x��5��Z޽a!�M�	?�6�j�-ꚶ$�>�q��i:�Y�I�u��o�)3�)7�i#kZ8��2���
��`���Mƴ�}��f�؍o�p��e�,֚=[�0�7��m��I��I�@L��R���׻���:.���:��
��M���g>"�Â�.AI�ߟ�z)rK>z�R�RR�:��J��GL�0Y�`�M�#�n	�o�}~2���Z��?�d|DR޸��'���3�7 p��4eTQ-�����9�g�ƁD"x�e�ݎ��߰e�E�����e{M�Pq��^���)M5}�f�!2GO����Tӳ^<g�Q&�V^�]�.칔%Wt���\�r�7���;��9��2�"�y�c��30��k��d��p�RWj�U��d0w��^~�k��Հ��tU;�K��$�v���}��4'7�zv��s^�"DH���<./�N�ڜ��BdF	S����n��gu[?� ���1�,D̖79��5����2�>2 �H�_^)Fu�;n�X���L���y�����WyG8&M��+\?�I��2!L���%��tw�g�P�.�����B����4�MGnuv{	�nݭ�e���W[����e�ﱖ^�Ov7�g��&ɳ������Q�Z4�0�ܤ�����h_�?�a����H�"D(����{�ϺBF�C�
��)��%Uv���.�g)`+[�)��&����U�N�󳷘Y��`|k� �"��a^#��Rk;;,��J:3Y�5��ZF�{^*U��Z�����s�IN�]^P����]�S^8Wsά�����i˻V���jX�e<�{�1�ۼ�c5������o|��Ok>���l�`���H��D�?g�����%�=5�*X?�&r)3�Y�Q�ܕ���ژq�`/�Y�,z'f!�O�}� ���$$^bF"M�I��7�����a=fSpmnM��Z�>3�����dL�dJh�ԟ��;�������Mit2��1m�t��ӹB:v�ݣLY�$��3�&������/�G���g�	0q���!��|1�\A
?1�$W�������h ���#I��Rg"f�O2�����Md|�Ԏ��~����Sb�V�pA�`���E�:}��tP��"�H�� �$a���z��7�{�ԋ;��@�o��1J&ۅ�FfH�M�oY��c)3����N�]^���4�7v� #���`$�����m[FF����Q�pA�Q������osB�Ułi"z��N����u^��];�K�T-��i}����zټi�UHੋ�C*���f4�N�
�h�OU����%�����*]�u���I��Rg#�n�A�jy�l��rN7h�S������{k�ط�|������A�"`�$a������ٙ�&!�#NLXm4��A�%M4��L�a��u��d'��e(��.�����~��7�H��A��4��kp���h�^j��k�p�k�y?:ϗ  >�A�ܙȘ>��L�2;��CnhyS�3�Ⱥg�&�4c��|91]�<&��f8JN��U��`;~�)���A���l��AKKq�җ8v熾2�c�p���W�M��� �y�?"`�#�H�"F�n�9�Gq�u�d����n�!2!��Vع�P��4c/;n�?=��1�7U
�^��0�p+���E�a�A� �Q�0���b���_tm>�掜�1[�L;�Mf8���	�������t�dسږ��S8���*��R]os��n�y�p�e*�sb��2s]�aA�*&�|/1j7�PW��wa��x��~���=|55�#�t�T�IR@���{%��L���\b��ۑ�{Z�sX�l�3Q<�3`�s��,]4��6��1jBź��m��%ce���\�;6��qF��<e^@.ȓvN)�e��a@��t�]\b�<� �g11��u�����@�h�ό���{<5�����vs��C��q���W��:���-�by�[ϫ�@:Xk2�e!S�A�Ri,5%.&:�U����ڴ`.��#�XK�}�㉼�7m��Rm�;�t��ShX��J�w���#E��l�j��a>"��+�H�H�H�x�������p� ����W���P�������m�+o$��b�_0#��F��W!�~A�|�a�$O�H�]�'6�u�`����+ݰ���F���g�l�S7��So��8"���f%��l\���AI���YӝEP�gEN:�� �E�*��꯮���y�@�������2�`IG9��r;'p�4Nk�?
�t�2�T���pFz<�G�9
;��A�ld|��wH>��8�~)��8y�&y�7e6�^�4cH��烍��3Ý����(0[>����~�A�A����Y$��7k�6�Ç"+��ܪ"[��ã���l2$�?Q��"~>�0C����^&=b�>)�Z�L�\��mҲ����Z��������ٝ\śd+|u�'�0��¤h���M���m^V]��$�ø�l4ų�M�_]�5�.�eBeY��z�{9�"�����m�V]I��Ѧo�
�8n8�F&pA�N��&��d���K;ԣ��D�ˊqx}�m��l� �i����|�9�N����<װ�AS�"���$�/d�����5�N� ��R��������F�+�;�3"`�DϤ^�DUT=��k�Jlg��v��{�J3*�Gz/������x��	3��p�a�r*w�_�֭��e���f�uP#3Y�N,˔��a�ҙ.0P�m�C��.��O���_��Y��l�bp����'D@������"�F^@����-�3t�1��� &���}"~"�d|ڋ�_p�2|��p��E�,�'L���pA�E����"�����пQ��� ��!2!�L�>I���_�Nİ��9��pH�g�}�����5���2}�gr�-Ս�[E��͘�zMY7t�
Hi��vᬱێqZ�Y��x��CZ�d�3�bP�z �0 �#u������8	K�wKĂ٭����k�p ���S"^�ۍ~9eK��6��	�g#y���İ�I�Blb�&A �LazD �0����vjp�)Qm����c���G��7�!Hj:� �~43�ߦkg�$�k�=E�Hx��$N� ���ہ:��n#3420����?gxw�l�}>�����y&u���l�FB�Xq�A���Y���_KC�A�t��X>a,�V�gLF�4��z48>n�[Z�6���'��2f�:-�����-���I�Q�wo.p8)�g]�9�����H ��D�w9�8�w[���Qev����]���?x���D�0�@2 �2&8�?�k[{���0~��ϓԙ��볇;�3B����9�~#��J�#*��w	�3��Qx�+u�?S?&Ov)o-!���[�`��E�d�<3�ڧ43Lȑ��+u�jO�X��̜���y�&�>u����G�^��Y0��'���D�:�$n�.j����L��(̓:��ɺ�����y����2��3Kr�up��~]���s�� ��*�C�N��+%�Yx9p݉�79%�^�E��_y�`���/}���ED�Á73��p�8�g���\��qԷ���p���L'�&��|���؈�YL3�S9��)�gvYÛ�ΝJÏތ��������	4Œ���4�4o��2�E�?�I������D�~�
���𕗛_~��������~�0A��A� ��?1��hnYk�t��3��Lr46g�0㩞c8>")���Ѡ��K�5�h�E����2&'"!�;Z%�ʤ�l7�[?��r��wD=����s�������I�I��˶��]?~X�R�e�u�,
�'����73A��U.ƍ�*����6����1��@�L���ىk4�}�T�x�e��e���>��=�(j�Zc���C��B|+V@r�le:6�ͯ	b�'k]�5��ta-%��N�<�vWy�nS���X��M�͓����om�p\驺�6\���1m�$]��8is,�t�F(��Ү��+��ܷgQ�k���]�1���F{=�j:�X^{ qn9�����հ�I���ƃ��-T��<�����*�9��)��ۍЁ�p^�X;i�'?��4-;48Un̦p$����p,���&�h�eGi�����k�<L��i��H/yD���#y�����ٵ�����b���C�P���wfoO�b�r�&DϤ~`�ȃ����t����
;��8 ��^1�W<�Fq�yܿ�[�b`�=��#&��*}��%l��`* ��O�"g�/�n�����<W@2���:���z�݆*�a��E�k �8�9�8g�]�͝B㷧vpA���Gs�l+�ԣzkb�ښ�v;{�oY�F�O7t��i�4OO�B�����ܘ>�dA�A�8$Ǟ������.�_`�<#9;���O�
�� OwP�7O�`n�v~X����4AK��H�IiW�,Mۣt�4���=���Z,�4�Jjf�=}�~�-���/���H>I�wn+bsx�W?z/��[������h#�A��&A0�7�HI��G���>9۳�,7M�E���{��̵�z����I����"�f3/�4kh�ۘwwB������������wi���\;�]��ڙ�?y������z�b[��D�n� ��M&c�<�l��P��@�y��3�`��`���)8P'E6(�aq���o���i��;�~"E�dA�~��i�S��wn��q3��Rj�H���b�}��y����x��m��y~pP�,� ��R��g���N_R����p���UlCsS����nz��g!���'u/�~�v�}���m�}��M�9Cgg\G��cM�Uť��$5"$�GDpd�X�ϻ�s�d���$L"WF���<����{�}�6!a��,3�p�(E��f��3"`��"`�W��le>�V1�oY�b�B�f�1W�?z�n�p/�78�oF����0��Ek`MLd`Il	�/~��==7zv��۷�nݺtӷm�v����m)�>���Z�k	ܱf껭!����7S�92���rwTfr��n����b�ޫ�{�.�M�1B2��cj
G6T��������"�\h��h׏V���C�ԅ����qM�=k+:7�ݓ{��[[��B`7��A�U���*�:M��P�S;�w�W���L<v����b��ڕ�4輦�Q�7-'l���.��CB婄V���{���撰_ul��t��2�q��:�si�I�]f���	"1d'�]3�U��ͺ4;xK��uɛ�|�!��=�z��t�r֣�ٕ�vK���2������}�GX��-��;���t}׷}n�L��~��z��uk>��Ώ���!�H���.�۪}�7&��d�Z�ufZ�y���ͪ��]�3y��&�P�0�P{�*�$&\��gݽ�����!�6�e��uur��е]h�mU��fv7���n�vwR��C�����-q]�h;��0<��>�8��K�oc�&k���!d�G�5J�zӹr͚��h�`芊�=����73j��ّ/J5��D�x�s�p^���&�r>	��dAu��e��W��t��I,���fE�.�]��[�o�L����5t-t9[\��l�'7a�[/Vs���X7e̢�t�Mw���x���Uf�b}�a�w�N�M�Z�cK�˩6���'�cX�uW�Qٴ��{0��=2�}s���ݿW#�B�[��DnK���U�L�F"���T�UUh:���9�bTCha-t�+��,��M�"
 [@��!�QGq�><���!>U�U}ϯZ梶��5�j�ռ�Z"�ѣW-�T[Ա��^V�[smh�5kͱ��[E��[y�sEy���U��d{�«���1��^^���Δ���-y��n�W��j�v��E�&5��6�6�k	�[�W5��\�[h�+�6��[y\���W�k�Z��5�Tj D$.Fװ�%�e,�6܄�y΢+sT;�i����n�泂5m�<D���oK?�u��|�M��wSO�z�?��g ���lccn����y���a�2�vM<��c�G7
,p�>5���A�I��&
L�Y�]��շ�L�t�f)��\��wX9s� �9�8�]�N��T�S�N�K� ��q�k��M�B�Ć�ɵ�#��3B������f�|��ˇ� ��������'}��m�?��Y�-�!��A�6q&�����,��>�@Ia��"�=bz�z�6N4�ӭy��3�<du�u��윘s޶a���pA�p�$':�H�$���<�R�5�dLv�����L�PD3{NҨѬ^<��r��3��o��8o� u�g ��8$�q7+��Msvͤ\�^������n8�Қ��n��>#�ɷ{�5�(D�x	��T��*f�/n��/ �cZb	���]w���B�\�uZe\�}��MV���=x�����2X��͌���忘 ަ����a��0AFH�T����S��z��G[�^���w3��n�9$�1����ac��M	7�MX�t�$�A�WC�^��;9�7N�)�]-��͉cՔ�M��>!<Am2;ܑȘ �����]���x��o�h�C��C&�w��!8����4�x�W����,���:,]ٕ�>�H߈�`M�y���kv?c����'r
k!�T�6L��[�S�ʕ�pc��#N�v�Ȼo"��a���ӱ'�=���w��3*_~���0M�>}�2$a��(C2&�g&~2P݉���rEc6g/��Y�Y�ea����Ff����݁�S�s��>�p�$��(��Rp��0��g�lÛ�w���St�ѻ��#��U��?�'�^c�̉�G����-�X�u��gL��F�#!�e���V^��Jع��f^l'm��C�Vﲰ/�Υ}����wKo�uGMQ7,_e�¨r����]�Wf���>���7�e�=�ϾTf4�	uTH�k���a�pj�ɚ�KD��3��)v�<����ʼ[��eҖ�(��²[e[a�]1�մ�� ]z2��t��	�M1�ۡ066V9�`Bd��&'�U��Z�m�F9�s�ƴ�Al
�E�X�h׃/n���ڶ�}Ouiŵ́�	Ƿ*:-�F�n(�99"�P��U$!��t)���UfTz��!��vs&T ���S�X��As��۬b:�k���*hg�d��۫�Y����o�þ�#:�+\9E��8x��uӼn'�!�V��ևd�~����i���;�dla��ȇ)7��ȭ��zꝝ�H}m�(�r<��j����y�6e
��p;��� ���E��2�-�9��� �h}���:"F"F�b�\w�cI��i�T.M�#)D���	Z��#��?A�?"{�E��ۼ���v��_�t�w��D�N:�޶���2V�7�2d�8a�&�1��J�6���;��������"�0�E��A��7�ֱ
{���1��p��یWG�AE �/9���WW-'35`d}v� �����5H%D��{o;z��9yj�g��C��֙�i��k~�����^�ɚ�$} ?�dC��z��9�G%��]��^�<�7JyO�{�!�wY��L�"��dA�'����=�.`��j�<*8po���Uܿ����Zp���Cn��&53c)�U�+2e��M�ɭ�j5�9ME�ӝ�HA]�+q�1����e�AX�����w��b��P7�p@4l��u�D������>G��{CL��2�ܼ��p�D�&D�^l��EA�A~*�Ӿp��wB�Q�`N� ��3,�#Kt�+?ګ��,�,� �����".�z��9�G%��]��;l�[܄Y��<�2�"�g���~"�@�"@��0��Aij,p�q�Vn�LVw����j>�a^"���&Dl�?3�)������6����;\;�������8����:���xԀ��rv����dH1�%K?��;���et+������b9�`j9���5�0@�t�G�a�$a�}Nd͖���d\�����ˌi���EuT�-�n��>y�{Y'1�u���t�*���F�pV0r3�n#�ٲ���=b3+rh�1KX)���=�]EZr�{�JI�S�)i�u,��������bM�خ�S��.��n��y!х�\
�Ѧ���'ΗS�ٻ�]�7з� ��%�E� ���L�pdL�3���R�\C9ɂ2&0m!��|7����Wz���㩃�76Q�oP�v+�3�]�x��8$��$�AIÐ��cp��� ��|۬wY7�	��P��f�xֳ�A7��&O�0)5��������[��i�$��.X;F4Ҽ�9t�na������4Ŷݬ��2����������` ���O������1U��Y�;η|���ڷw��pV� ����$A��k��	�g�Gw)3]�$���P|C5��7��a�Wz7���Ƀ�W8rf�Ö�>�U�(�`T�pB�B�rIÖ�J<� �¤����4y�_�ف9�*�A����k)7���5����aDN��Rp�62�ou�y���m��"��`O�z��ڥؗ��;?E-c4
ò���X����ܰo�2�+�j�EM4�N��ѭ����b���T���#/F���Xȭ��Sp���"5�Z�I�� ��A�2L -�9V_�GV���h^�:��k�y��a��`�#���g ��Z�=o�����2��h�kV#���.�`S�܃�.z����.1\ɖ��,>��2����Y���w� ��������y���B�v����ü�����e�W3�	I��"�pR`��#.;�@�T����������ld�*�\紇Y�ۜR�"��J ��7�OUmq�?�K{x��&> � �p�	�Z��y�0���$�%��3B��k�y�Ï&�Gj��	dH��	��X;�믘~"��Ĥ�Ź�s�4�M%q��������aGm��&p�o$�
L� �dH�׳8�O_�Ja�$���U���t�X�E�3]��B��"��D���2�J��ީ�U���^���׫�����g8����L���d�yft�u:8C��t���XR\�zl��%#+�W1�����l����U]�\|Nk�D"�;���u����y�\��B���j8�`�1���MZ�ut6��0���M9�[�.����������u-�	�)�c�\��z(̹:7.٥�7b7e<�O]�� �9�v��V�:�����;�8r��{+;��cu�o��D76��a�x���� ��s��5V���v�]i��q������ick��ں�(�埿q���,��Y��pU�N�s:��n{=�J�����_'��o���~z9�����̩3��%d6����kfy
�{g������QK���<A�s�u��v��I�BL�<X$����^��I��f�q�W�80sM�RO����� ��I� ���I�K]���'��g�n��o?�)8	7��8R�Oqq�qYT�x�տ�|"��e���a��!b��U�>�`�!��[O�G=CI�y}��V@7l�H,X�b2V����w���օx��㹟]��)�8����dH��/0)����!)���6����-���
M�X�i��I�f��۹� �{��0A2,�̩�V���0�ޚ�i�-���u�G&�
�U���l<YŎ��E6U;߯|�� ~a����^��+�nMn�jnZ�Bnp�A�"�KYS�#S�&�M�&r�{�ݡ�\�w��S���j�a3���BK�j��^҆݃J��1e�7o�ٛC�uQ�g�1���/+�J��>F�OԷ\�q��[o�&��P��~1;��!w�?~���ȑVD��7ݬ2*�r~H�d~~&Dق����I�)�D��z�v�v3V�g��&s�ϩ8j��ɖ��׌	���IÉ׉�[��7-Y��S9&0Lb�����X�I��"d3�%��dN��;��?�$F��h�u�B�����[�q>f�`� ����"D>��Vo`�H�@�B.~k.�3�#B�;[��+U��8;H����s*G��@��O�9�D��_����~��o=Ev�pF�g]'�j[���k7��A����8 �È���[2_\�o�n��.�<[�މ��\���Vh5�p|D�~$���'�6���g����L����]�q7l� ��>#��M�����Kt�ޙc�T��M�Ry����[i\��W�{%j2������I�[eY��S����;��aC���T��`.�o8 �r[�!&rI�J|�3�
u�N�����Կ�I�����]��.z��v���\����v�sS��>=�0�@1 2$Z����m.*$�"]Ìe3�"�b�v��E78$L���-8rw�4��=�}�}���q�yy�L���h4���:+�v����z�̺/ʒ�R*�%~6��ڦ*j0r�?��)3�B�p��s���p�E�w�A��?z}@o,�Ma�#g!��_��#\��_���N�'9��Xy{��7<)k�w�&��a>)6����ۍ�QZ�G{����W��`�L�9�8�}���*2z�l��5�:}�������~�v��X`���7�j�$E��m꣝-@@;l�7��&p����v��s���O���=�b��#��f��'��	jBn�-�J�}d�^ii\���Γo�izVʫ
��e+���{M]��4%\Zg-X�κ�$����W��x�7� ȑ0A����������=L�q��gq��.Z8U��p ��� �~��������u�T_�k���-"�&��O����.`K��u��ېy��R��y�e���>=h�XdH� ���,�;e놮�`�qh��8:2�v��3ꯁk�"���?"Ș �^d���1ܮ�a�4�\Ê�r��BD^�,��ZBЊ� �n��A�p�$�X9oXg�[�?��/��#��n���Ra͢qݡ\k�Q�>��i��fU0�*�#X?A�g���I>��W�˧�VG��@A���F�r	8�ϻe�F��a�1h�oL��4@2Om��x��m�O��8$���D� �"`��0d_2s�Ѣ;1�^�G\	s{��p|V0pG[!���3�FaJv��鳦��v��۞�_����x�}��W���%�U��	�o����>�B�:�m�Mfݫ�r���̫��'u�Έ�b����嵭Χu����t���\���X����;"���僴7����ܤ�W2] 늱�Շ�^��6��ܸ2u�Σ�{�C.O5c̾)\�JՅb��ꙓqy[�rW��L��o$ni��4�RU+{L�DҌ��k	_Z���e�bPe
�K�b��t�8n���LPZ��q��f�B�ن�	����S�j^}x�k���gU�}I�ܵ('�*�RǗZ�6�xe�r���������d��}+*�d��wd71T�3F[v&J�uه�Q`�ٲ������.s�n��qGy����ν��t]U��MK}bvQW��4��S������cS0k�����[�}������[��9�{;�����'k�c�&pk��7.M��Js�N�͵l���t�߳��\�*�r��4v�v�,�;2i��&bh�|(]�e�⼃:
��ѽ�{2��Z�;w8:�w�>_=-yE��������ߦYW�ܯ�*ɾ���DxWV�����@�T���m����������nV��޹}�#�\�Z�	�W�h��*꜑	�Y��U��Wn٫�ɷ[:�T�2Nס�AT�7�طYɹ��M�!�*1L�xu�;��e�sHnwK����^<8��cnÔl�=��kq"�;Zn�y�n���n���U�a�f��$1շ[3w�V&.΄pӫV
6!�('�\j�\�H�b���⿺����Ϊ�_Y�Nۜ{F+b�:�;��L�'�	�嘻y�b�"iн�#Ѷ����B��E��sk��[F̤����A��m%�8����nE���a(�Ɖ)wj�DE��4b�AnM5vm��b�������`�n]Ks���F���+��c`�h�lb��5^��&�b�2j�	XŠ�6�1��9�	co�]z�؄�b��ch�0	���F*�K-���fa�}��;���m7�!�k�J9���R���՟(�=�Vȧ6F MH�m�-�+�R�f`�z�'v�v掬����WG���f�.�.'1�Ba�.�5�Y�ĢR��S�Ц���u��i]\���f������\{�p��$�\nnnnG(ً6]eqp&Y)q�1F1-!+���b�̑F0���5�3hMa�
�,mX�@d��BF�eN3�`�7��n�hG�́]l��5`H%��	�t�q�4A��amdf�st�r�`����h1`fͫ��M���3`�';���aN�f-�`X'�`y����p]�����	�Y�9���Ei[-��fn�����^;FkZ�]��R�X���h����B� e��/#A�3G[	u5�� հWky1S�u�8/`ݸ�f:Ep':��)�L�λ�c��6*��Ϙe|"�
4�r"�.�l�׍��q�[;;Ea���'\A���у��y�	�ҕ��:!痶 �n%K��Z�f�)36pSo`�l��u�� [,�����9ʴs���g��!����g��%�?:8��M�h�|�wv����۷Y�e�c�]�B��EQƳ�S��!��wP<R�Żp7&ն��F���j;	�q����x���Wm�=�<7nlF��N;^.���p�Vۨ�p<��k�����.���'b��s�&$-�쑻{�X��˨��9�Bd��&�CK���D,ck�hK��if:�8��Ql��ԇRR�F�[T���!m&�������t-d�-p7��&�,s���4�;3���!ԗ�=�b	nkN�ݎ6�:G�I]A�<��<��� Q��������{���$E;��7k��Qy}L̳MaYy���7c��Vf��B���b;]��b̗gEpu��u���NZ��^Kr��h����v��cb+��7l�[�T;f����Iqu�	5�C[�2v6�:���E�aRj����g�=߱��Y�}(K�v�&��@�Ul̷�4����S�͕�6�5�S�-քN�x㮯L���t@����ũ�nbE�%\��T��.���W�{�\����Mv#���$%��xs�+\(��\��\�ix�Ÿ��Q��1uӶ��vlڃMv
B�c��r�ݣ��\벣v�ƅ�9���f��s��������c��O?��ҷ1,1�Xml�tܔ=<k��Xn�n���EuV6ݓ�t�����}�x��ߏ�)0b�T�|˂U0���z,u*X5��c�鉂	�A���3"~�!��u�A�@V����꘬��.�D�:O���W]��b�NüD�9U�r��*���l_���=�`��y�f&�FKU>��9�'�d����h�������ռ����� t���8��\��+*�;I�
����E������=��®����l7�z����g��ʵ���g>�g�8p|R`$�$��ne�dl���/�k\?C��/���;q�E?x8-�Ӈ$s}�%��o������;h�xK�02���+v8"�d擎��3���0��d#�eK�`ߵj�	�'��w�Մ5<G��13�\�e��ռ.Qѻ���l��E���$���	@p|B����s��K-m�a�^C�s)����"�n��i@��\A��̛6;�]�6n�;*������i�xM�Hg~�"���~�9�h�gW	��L�}���I��'ͺ�&j�'uۧ,`�sϻ���#}v�]�ۇ���[Ź�f$n'g8Ή��49�φ4?.� �la���0> $ޮƜ��Q�$�
�JL�P�l�[<�-�po�	�`��Y˅������c�$�8 �8 ��8]��5ӣd�mo��`��;B��aՉ������w8)3 ���������V��n��2�qs��{zBܽf� ��3�q���\�N���7���s�Y���`��H6`@�m�1+Q[{�F8��O��ujbd�	�h���Q��������dL��-���xf׳0�7��j����kg�w����pA�`�n8pBMtFWܥ�������~ �#��10�爻��1nl����楮5�h��c�M����̻���P����2��Y��r���Sa�r���b�H��[�s@���4A��i�e��y�~L�GF�vŰ�w��e�i��=��@>�ϒw�ji�s��y�t&�`?�H>I��LMp�+w9��Z)���,����]���.o8;��&s���)3�G#�CLN��e���#}{��Gk�Bw�������ۇ$�AI�´_�4�=g�h*T��e�t�$TK	Hjٗ*Ph�m�Jjmtm��]|���'�Y�9;��BNĤ��+0q�����ﶛ�Cft��{�qkSM������%&{�?��8 Ű��[�3E�������mM^�4��Y�@ʁ����D�9m���W���}@�5�� AI���8>I��k�1�ez���l�<�w��8>=����g����
0ɘ7��¯N}��5�o�������8{��m﹊�r��i��n��o����0�90���ӎ�c�m�C�wQ���7����hlѐ]3�rS��(�!q��[;Jo{C��)lUt��Y��j�[�V�hqߓ ���3�0|dA�}#���(��W@�yT���)wv�a������D�?�x�ۇ%�⥃��7 ���W7,ތ8{}��j�Nqɯk'xF��in�W�E�M����9��E*	��R��o����)�E{E�ml�=
����q�fMӋ/W�����p#52�2$@H�����}��:�9n�'��evn��.s4^�n �v��+��5_4�=@��3�n��+X@!&�O�>I��唤0�PZ�=E��4�7Ki��E; ���`�$��2 ̉�g�}�Kž+��/}�g�7��Xu���c�(LDo�p	�`�#j���f3�o\��I���9	@�V<�yLj�u�Ys��������n��>+�9I��)1�T����ubj"b}9�'���E�)��Yoa{_h�Mn�|�@���k�ju�v�[�e�+c9��'��0L��Q3T�,�4�TZ$�ʡEW��
5�:��%ჶ��bݞz3M4��p�9W��J����l2��6��(� �o��ko�ɻ(��@+������t�/1ǳ�ql1�WyY����m���e�q�t�5v����jjDҷ[�����k`<��5����v�+K\�@U���O�ͣHph�4�j�;I��e�.ݦu%cڌ�iG>����;�w�]>	���PiT5L*�	���%��y�I�:A]�3hBZ�M�]S���2���0�6�9	3�
N*fWq�Yݥ���эƏ����C�D��ϗ���"`@2&F�
���b�6�C��LN�q�J����{�;ռ v0rL�q�t����\uќa.7[�!`����,��{\^{��Y}`��ae�f���M��n��>=l������?�6n��t٨��\��x�����g �'�3+6�.;���Ú*88�*�Ԉ�:��'�"-�p7�~D�AD��F����?���H�4N�_>�E���o?�8#m�H����n����vB�V�R,�"[5���v�E܄ɸ�1Fi� ��W8fH�M�Z����~`�ڙta�#��Df�&�o\�h,���L�c�g�����;gu0)dL�["�g��3?~��~�������J����GU+w�������Ǟ�5y6��v�sp\��5�D��z�`��90a�1;�@��>f�J��"i���Á�3+侀��F4��Q��?���A	�t���Nc3˵Q�����(��A�u�f::4�4}��10���!�<Do�x8'q�q���BM�"=v�z<��?M���ڼ��GS����o?�L�[n��ŗ1�/�7@7n����k�!�M��}��|���0���	6�.�h6�U����CˇѵJ�^�3���v�4T��!�RĤ�����ƿ0�of��>	��Ő�]����������K�LLK.��4i�%�&(��%'��}���2'�)3���3��;���Dw�y�::�o�m�0�rd	dH�~"dZ��-��P�*�񃆫��s�~)�,���r7l���`�&=�Y9*��D�����>���$L���x����mg�w�~Z�����"�l��U��V=4�u��
ś�uu�����T�^glB�3Lwt�E��2�l��j����4ą@I_�ݷ���F���O�T����Â�~&D� �~�Y�������_���0��NS1O�3OT����o�ްpC!ّ��j'аi��"��x���"Z��ȅ
)q~����@w���_�>�fn��~)�,]:���9>;m�O�\�\ᦰ_ߴ�]���4( ��ؑ��II�n�K��.6	��S]�s��Yr�i���ϑ���>�p����>I��������iS���Tprz\DSBe���E[��)0���L�"�ʙB�[t�=�\����7�?Ep��n��>��������10r(�<����h�)�����13�}IÐ���I����a��x�n��q�k���M�r��8:�8 $�|�?��wf�2�!Ry��A���57�'.fg7)�o����>���D�8>躻�وڃ�"-�tK6�BRv$�rԻ���b��̈́�~g����l7������P�̾ә�n�5V�,�O/f�����z }��IÁ�����$�|�y&4��7}��g�teZq�f����#�[��c����D����$����Uy�"�H9;1Ab����۪��0��n�����=0�n�~�F7�,p�/�?�I����2F~)�B��n"7/��u�t�c��E0���;����u�*�'�B?����V��fg7)����M�>h�a���t�h�ː�y��X1-P�GO2�g��,�ɂ�E��A�n\��]���v�pr&Q��c7����"�������>���I���8!';f����)�@����?�L�t��l���S\��n>�ޫxȦC`���OY}��8γ�V���p���8 ��E�;��^�����DM��l�������FO�u��z|����Ԕ�eV1b�֊��%%Y�z
>/�]����;5�w6�9L^�o�tͽ�{�^���N,��[�t��X�";���]�s��+�&�� ��TZIE�e�N�D���ݮ���^�@��Qre�u��+ۭ�v9��̱�Ӱ�����)�n9��u�-�u�u�j5�ff��kY��=V3D���4�3�o9�qXh���ӣ#�6��m�M5�p8�bk���1�-a�M�J��ݣKR�c�6S:e�m��M���D��GU�0q����X����ն5_�> ;��_S��j��oi�xq��V/��z�.�l���&=lҶ�H���Yn�2�=�Ա�}�pA)3��M#��{���8Q��
��3��N��`��������Qr2�Z�-YO��C�1�l��'��d��n��ǁka�M�Ɖ���x?E�R�U�O�A�"�Y!��������۫���M��v�Q��5~>al�Ϙg�E��!��TDy_eyQb5i,;�@ƙ3μ�a4�fIi�cS�z�Jփ�8#����^�	0��.BM�)kE7sA��s�x���eۆ�M�qt�w��3�~ZC2/3"R��U�X��̆2�x�
=����q-�Qs�;�fػy�oC�Y�����~#�A�adH�;u��ǧGm����.�u�ۚlf�(@�9�X~1C����#d�?}����'�z�ӑ#�8Xpۇ"��pN̄5�\Y���a�c&�qF���f:7�vcFiCk������I'*�f�>?/��:�� �3��%j�Z~���(�0&�o"�!ѹ:^�p:`��p����	0rw�	��]bX*Sʺ۳���:l���[��[7�y��C���}I������vE�.�Q�LJq�6d��/9M�r4v�J;��o�pAF��l5>�>6���g��#m��#�pRo0dL�P�E���Y4u.�A��"t���L���1��x��>^܁GN�������sj�lҥT�6�ղ�m����)��g���{\)�`�ܝ��;��o��⋂/�9	;����Q�a��A�zl�eӭ�F�٦��Ú��pA&�v��v��P�Z���s�|`���8q���3#Gm��܍\���>�0ȓ#����fN��Y�+�3Uk���avg6��2ǧOM��;i۷o.ݺt顧/�{��ŋc��Yk��p5�vA�:Hk����y�G�]��4��Ú��b����4t�y[��1V��#{2h�Ώ���Y)�7h��k�Z�x��ʽj]��e�R��"�C�F�W�]�s֔Y�&|�KA�9��k�󾬿_!nfQ�ƒ����u�f���CE����^�D���ۻ��fR��2�1\����y�˂���؝<;RP+�ڢtΜj|]�V�mǚɹ�1��SEð^�]��*����[�CJ�K�o�H�h��sTw�uOv�,f����v�}�е�u��pK=�WSo{%Y9�ܳj�M�xʼ�e��brd�o�3�#����k���]��9���y���Kg�E9_�{e����RW�&�]�R�*�i�J��`&������^�pf	WhzZ��b�:E=�qD^�r�"����M�4�2t��9�/���]UR�Yj�m�6�a��JA]N��u�j���osMW-�p��Ѕ��6��JP�7�w����LPE"��crL<a��b�[S9�Vcr��d]oqkT�k�8��"�Ʈ鋽���^������gYvJ��	��^) �Ƹ��D�s&��^��.�lأV�c�Ȏ�^$7Y'O*ĩ-�z�]�ʘ��K�r���B��e���e�"�nb�
Y���e\�w4;ӊ��v滘q����V��z��!W³I�Q0a�O����ǳ��.��'\!Ԇ>��4�כ�I�<���}kJ��NU4'�t��κtc��G�3�A.Qq�݄�p�.$������lۢT	�llD#),D͍F2Q���`
��Q%��طYEt��DTZ-
h��kQDRlHhƊ���!FƢ�k�\6I�D� �R��i#QdƀH���X�#EL�ɨ42,����LdE��6KIQB�Hl��`�"H�F)1�1��l�Q�wp��2R��F��D�4ط:@h�_�H�	�HM��!$l��J�&�^��=�ѱc!��R)�b�$��	�{=C�n�ےڅBh�Gx0&�q� �}"D�F�/~�4}~�~��`��md8e�k�csq�|����pG2���阙^[Da�g ��;��7 0 ݰp>�pࢍ���9�0�X����6+6���zm�������9��!#~ E=�[,z{���}�_�T�]�Ml�[tf��CM��h�-�Z`����I7L(�DX��\>?b���W��I�P�;w�ۮy�T&�w�lT���N�.g`,rp��E�!&I�QpFS�A�cv����kiOȾ��n~2ϘV�7]7�kY
L��h#���٭P5���0��I�����`�\�p��خ~�g����]�>��Y�SnF��#G�Z�h���
M��n��6��A+X?��r<�?��k��}s�&����y��ផH'� ���_�ܧ�b�q��u����/�W3��'7k隵U��۾��F�fQ��87��v�~�3����V�DEN�_?;���������Ϙ%p!3��p�����z4f/�������!a~{�n~2ϘWN7A�g ��i ��6�5[���^&�T�TI�:%��@���2�M��|l��VB���	f�vk���{����$>1�I��'6&7_3A��	�FO�k)w�����5  �5��'6�3"ddL�B����4 �2��T/Q��/��Ri�Ο[���A����CsС�1�b�\8�0�oa��	8/XB-��������x_~�]O�S�+���{Zϒi ���x����.�/!���aG���Q�y'퍩�̝���}�ђý�k(ǈj�XK��ݐZ���#ua�u0AV�����ޏBk�p�Y�8z�M9��GH�V0���(��½��8ܘ��˓1�������������%rL�I7&�_YVF��ݜ�8k�t�/8���b]=�l��^t3ds9�V�������x>~�[�@4��9�驟g1���_��:�k���e#�2l�`6�뷧@��u�� ��6�¥Ζ.tKB:��!�q�n+ځ�ڷ�W-���od�����ی��XAۑ��=U,]��%�A�dέ���%4�=.�v�T�ܹ��u��<$����r���F��"$x��P�1�в����V�U�f���Jm��߯���K�`���YOt<'��W׋<=9v�A*�iq�I�u�<:���O~~��������Ƅ���Q��.�y�ߥ��)�1�7Ig�:;-�<A6��3�JL�<���`|n�9Ӕ�ٻe���ϭk���T�fN���>�h��lӀ����͚f~�-L�wj��k$�&I����oX��� ��U��/)��|���MẒ��1�A$��~��ոj�����|�>����8^�o6�#==�#0������Of��E��IHI%�ɁOA�ޕy͹��+��=�d���l`�DG�ho|�[����qrRbYe�U�ە��7�&�ζ�6���T�L"0QJ�pU!ݲ\���3>�`��B2c��f-�S�뾑=)�u)I%!� g��h&oC�rpc���!��oh�XRMU��F��!Y��;L�PqB��![C ��Pll��R�Hk�E�'q��]X)���T__���?s�US�z~���4`̍����!9�����a/�-`n>m�]�܁w7�/:�:-�u�8��'�b��{�r+`IJL)�2n���(ˬ�����Χ��q"�'�{°�#l�e�a��Zh�N' �'H��=�gb���T����x�fh������No ��x��j�.���������'\]���b[TL78�M7	Shr�CD;�����o����c��k�-W�9[N��^(��M���{���3�O턔�&	6�|��Ztm��.�'\��緞q"�g�xN7�RY.�g,�H�7x�0�����Q����j�!w,c.�����k�V)L��җ�y+,=��2l��v��u�f�YJud��G
�♪�	����(��}��9,W\5�	�n��f�6�޹`+����`.�$�EodC�M3/C<�j��P�����f��F���=f4�������1�YL��S�&�M�#�wf�]�W�{�~e�!��~���TMd������sz��6��f����>x�~��f�R���t����؎6�[�u���ISd�t��
|׌	�H��1��;4OKs�lo�r��T��J</����M��&jrm�vQ�����f��Mz��;��['�����YY%���sE-�Ce�I�OI��N�=���W�
��]����c����2ݜ=��v<��S�L+ȴ�/���C���hU��0	'Rj��K�B'��o��x�6��p��?^Mr�g��eLljC�Jѿ��/v�hN�Y �Ĵ�Pj�- ��ājg�Z�X]����������k����P��+6�_f��Q�9��;�YB������a��%��v��ݼ���b�O�v'sƖ!���N���c�]��p-%�V������	�2�2�iS�H�)']$F���Us�;;v�!� �b�^L�"�π�k�~��A&��`t�u�"y��n�i^�:a�%������_�2LI�^��s�Q�v���\)3[Y.{���q�]0޷Kscu�#���v������I$��_�p����y�.�`ە�»�0I�N#�8�ð@����О��d�Nj.�ΗȞp��[����{ɞ֕=�Q�l�3���I�O�%{���w>A�p�mY.y�1��[7�M��޸&�x�n���{�Ԉ�bQ����XPk���M^�j�T2Ŵ�~���ﲳ�q��$�+���C/E��u�A;ΫZ���n���o��]��ǈvҤm���<�\�n8���;v�U�K���i��ܹ��n�{�����/s���C����yéJD&,
˃1�0Ke�ט�b�ܵ�Ӊrp���CK@g���ۚݸv�h�7Rkl���h*L�,o
:�'mgg��S9�zL����s�8�$�r �֧�|E�V�����f���=�#�x�&,k�V�o�����]���	�WCZ9N��L儻gg����/Q��,��1V�[����y�K��ߟD��&lΠ�A�b�_0;>��m{�n	|��av�RIO�탁/�ށZ������Z�o��]8]�y���� N��I%���fWzSf7_:M>Iåj����<;b�k;%��*�R��q0�rLIJ�Sp��mgz�o&mޠ�[e��]��ݷ�Ŧ��c��$�&�I8	]�:l���U>�X_H�ȝq�=ޝa��'�KO)�U�Kē^��1��u�e�T7gg���s�����x]A�,Jöw7��Hh��m�F8�o$�I8�5#��\�OKZ���k�}�w� �t]e�M䓏$�+��7�I��y��m��pn�c���+r\5��qwY���ƅ�J(�(Bf*�՗�8"S6^��Ũ�m5!G&�[1���J�9?
�����y��B�a��_q'mp��d���t�͍d�{��˹/II�d��U]KH�1�H=Р��QM�8�'&`t�
���I*�:��d�^>�eOB`U�[�螖�M�J��k۾Mf�_�S���BHĈI$;��=�8X'�i��P��i�t�q:�|=�_��$�Ih����sSi0�����rOۯl�<�MkF��M���L�e�R�����c˒�I����R��Ȟq�=����o5������&&$��E�k��ǵH�mܡ,+7���������}�7>�C�zĭܝ�Iy�I��u�����v�Qש��
u��;ڬ��u6�-o�����NoK��u���a}FG[�Woc��g���ѹ
p�l���)WMW�l�}2q��F��q:���-��ݷ��=&ylܫ�C����v��k��f�ג�=B�*zw���e\&ۣ۩���&$�I�[���Ȇ֑����W�oe�w9��ߵ�$�ƥ��z�0['�tRT(W���h^Ups��;7u����f��X���:�������{m�'�L��m�ѯ��՝p�)᤾�8��o�����r�ڙEv��h�a���ڮ�f'�T�ON�a���(4N����/Dm�� 3^F�	]�6N�7u�`.�{�"Z3w9o���0o�$�^���0��a����ݡ�4C>�.5�-��oG��s����2e�D�Eud3�oQ�|��hf1�r��9V^�jC��%����
�6��,�7q:���[<����m�L�M��6b�>�$�I�I$i��c�n�W�).ꭵ�+ا��YU=;�Ӭ�J|���E��B��]5��Y�c�"��2�5H:i�R��G⤙����6&eF�St�u�mT�l��ԯ�����J}R`Wbm�yc�3��̜��)��:�����!"�1�ժ��~�vu+��Ρ���>�.5��>����$�[_���Hj�/��+ݎ����&�䣯#�����ջk>b٧��YU(uoO����]��$��݁YQ[`N�m��I�Y�o��E�Rh�С�-�4�Amm���W7�g��x���awoTښ#�	��ٶ��#�g���{�v��9��og��9zcN�zv�۷.�:o�=��O���2�Vf���&�6�9��;V��{ݮ��V�)�AY�6�x�Ӹ0�⸨�9�Z��
�}A]�2�sl�9צ��.�VK��P�(�Y.�s\�1I�DӘ�S�~�^��۠Q�r��؁�T-l����,θ.��%lΠ��4�vY��o6�٪n�ꛛۛ/$��:�ue��׶vd�y�݈��8��sW���rиQw7�ڮv�3.C�4���v	��{��YC�be��)��3��:�n^P�a��w��H�&�&�ƻ��j�;K-M���y�ޫ���ǔ9��zH�DU	�99vs8�G�+����T
���q9���Ĳ]i�:7����rX黓���-��7w����ĺ���3h���;��*�=+��v�%n0�2ٽX�_nm^�b�)�5yW��ZKpeB7��$�rnn ����+�;{��TUc��2�y'V���W�	Y4���N��*��&{k��M��}���a�y�PUm�'x�5�ĕυ�ݼ�E�&p���˺�lq�}���w!�.E��͹��C�Uw)ݑ(+=V�hz���n��L���GU�ę!����@�]�s�s+���Y���u�Nu�*.�/N\�U��>��l�����A*)X�>J�u�yu���Zw:+މ͐�����r�$,a)*^��}>�I�������DG��6d+*���V�g\Da�;�m]�G-=v���y�����wM�WY}����j�1קs�mY��QB5NlEcqjbM���nN

�2��s����Q�ڱDk�cX����)�g���lc��D�&LbD�4LL2F��Rfc�n�4�����FR4J	����3"�$�&Fb� �D�
R!	�T�ӹvH� �f4�c2fCvcH)$�L�!�(9vDa�	�"�u�BB��1bC �@"bD��SEX�j2$�3I�BI���M�01!� ld��I�����P�& ��E3%�ٍH�h��f�	B�2v�qH��$&f,G�زR�(i�J)�Mm)@�lb�Ke������Z:��TP#/.�f�l�#7^�l"`�(�cz����z��v(�m�Մ6m���]��V(���������/���k��j:\����ps�

v�;��]of�.�)��0��D�M����>P^��Q̡�Ԛ�ƽ�5Z�:�9릎�t��/�c�5{6:65+i�r�ԖT1��ɗZ�s<l�`�{�.��]� �[�L����K7Q^���V�4L�\.�d���A]C��ն����#q�]�b+Rcf�;uCܦ��V�k�/f^7OH�r�ڠ��ѡ�ۮ��/n��f6���)�a[���=tv���%(;ω� 0k�q���-;Xc�ps��!<����3�.m�鋢hT�m�4F�b^�^��+�u�mD��B��m�86��g��[����M�e�K����#���c�wS�qe�W]�-�#�b��.�2νv�����@������0��|����,�Gs��Fn�L������n��sX<B��7`�na.vS��q�
��wZśK�M%�B[iqj`�(%&f���tT8ɰ�U�;e�\�&y��x61�\2i�,&젅Kc&�٫]w]����;Qf�[AƎ��8\��N���)�p�uz@��Ɲ�/�Q��fr���F��z��u^h�����)�d9��Mu�Dݧ	��v�/��(��훆��t� �}���[��%t
gK��U���Y6�&�k5B�nb�O�J�f�ɫ,��&��c��,�@d\t�"�������,�,;RX� ��
��H�Y�,7u�!p�v�='Y�8k��x/;�o	��O"[u�h�*6 ��Z�k��X�l.-Prj7#�Ћ��瓫|���3�'�r�m��h�$BѳBn&	X���ky�\Wm4�k;�8��Wa�֫�a,quSiM�flK3�la�^���ݮ٪�9�Iq![[q���Y�;,�PE%o[�i>}����/�����.I�0��������n����n���u���ǧ�f܍�Kn�<H<V�'�<5�l[p�v�U:��Y{"�w]�a���F� �a��,��+�#�&�㴺n��5�ut�St�)[�	e�n�m�:��b��ڭ�7i݄���6CZ5Mn�t (�.���!�׋I�uZ|���Ż%���qb�o^�?2���-�����|Q�0<�
:&�uV�;�ʦ����s��n�%�	y�o3��
� ���-p�$�X���^CTr�Sӽ�C����t�=v�J��&oy$�i��jh��č�qr`Ww[뱺4�q��Cw[���.v�����1G�[{�_�PN�Uj��luOw0H,�D����W�5���5���a���B���U�n�o�p�m��yQʎMOV��oh��6L&W|�N]�K��I�I�LȑQBg����`9���`r��kj)=cnz���iF���Qz�t�����"E��ʻ=һ&���/"�K<�ȴݐ���f����îm����iIǒ�[��Ċ�ᩖ��Ud�]��*�7�}��x�뗸�&%��6Oq:��YqS�h���d�я���e�����6�NRz�#ib�T����8��'پCYY��t�h:{r�1a��!�(}�o�q�s{���O
���G&��x��`�Q׳.L�0����$�بqf�s޾�39z��m�JQX�P��y$�U/�3-��]\��c�Uyϐ�+o��೜@����T;�Ȥ����HI�O䠦����3�<�5���ר�&2g�xm7�RS����A6����v�p\�wf��u����Z�#L7"��UU ��? J�Ij�����$^G
a�^-~�s�JP��e蔨��i�/��$�'I����v�n�[��f�5����ki���+`�8|�`��.��'u��A�Wov�%����5�]G&�L(Ɯ�ؠ�Z$�Qz4��S�2_Z��/*�����ڽ雨d�m:�Gsp��-nPܠ�v��Y�?���	ތ�mx�{u��?V��ڿ@֔���v���u�
�ԒSk9k�w<�2��z*XMb���t�����"[٬�p�! 
I�g�iL�\��͚�&�`��s_7�y^�U&$�a�ŋ+E�ƺ����W�XG�16�e���L�R��;��OK�ۜ�ES�D�M�����?}�E�����U�O\��3�X��hD�̮���Mj��av�����!���w0�*���u	�&��o(
r�Z�٩r�}h�n�	$�$��b�ͬ�|�+�X���3�������k���P�%b>��7��b'��p/��♽y�f�����/�1��u4z�Y: �WWA���W`�;b�9��s����^�o���o9W�X2��Ø��k���~D�_V'���w�eP�-^�%C�f��ك���@�f����7�f�L<�)�QF6��)��ԆŵM��t����#}����gU3�K�5vT�`��u�G,9�K]ΎgT/k��&:��� u���#���-����лoٞ��/=X��������,�a_W N``a���욃�����Y��M8�����3ӽ��Ie=se���������uk�$��%�:��"�����ӭ��e	��������)P�$�m�;7��8���_vO�'�t�qhy�e�:sx
�Us�q����/73W����zD��O}�!�mmN�"M��2�Ku�Ɏ�����	'�J}^wmbl[��c�4����B���͢*j��)-��Z�uR���"��-��G2э�i��o��:���`�s�&3n�j��l��z��B��+���H:�JwE{�#�L�kf�4��ҁL�k�69�v�0o s�qi�?<������"ʚ�5�1(U�u�"�ڥ���uy7���;<E/<v9�]�5������������:�Gэ/�n'l�a����Ul	uϥ}c�q��6H�J똵�q����l�2�7�n���JS���"�ꥷV4��ņϫ	,/���~�f�Y��yv��y�9n�P�&��ɳ���l7� �_���av�$쥚���w�zV���`��I/w3�L�t�2�����ٛ驎�r���:s8��u�nN��!��nǼ�f��]��>�z�
$����b�K:���赶"U�l�9Dv��a��$�&	7��t�S��o>�S�`.�éf��l�=�]+;��9�qdMq]�T��MI@��I�[��oK��;�iC4�PW��Q��{:o8z��޼d�$��b�T�H���9������In�8p���i^g�N�b�P.��ͬZ{8��g/K���凫��o$��[Va�7Z9���}uQs]�]�� �y$�����ߵ�����Z�
�![Ud=,�̮��7L=P��,��y�7�vK6��t2�T�囵|h�qA\����	��ky}���!�~��ς*���D0>#y8Jz3&f�3�D=��kd�|��T��f��l�|ïb+	$^>�ݹg��~��;߷u������C$�I��_q؝X���n�	0����8��&Ȏ��w曌Brf�&ܿ
ġ$�O�e�Nni����_L��"D%g��`dw�&�Q����]v�j�&ɑ ��@��۩�싳:���땇�G78���V�t�vy9�-���}�־d��������wQ��{:s.He2���=wbM��I8I��`D�1���Y���E�(&걑��N�;����eq�\�$*��ĕ��%C�����4����QJ��؝T�R��8fz]wY�;+p�`��*��L���-�c
�sYO/�\��N��,����gv��]u��G�1q�����VH(]E�ؕ�B����xa��>J��$���m87�a@��&_'��K���ۛ"���s�]���0䒔�$�%a��^^�V %��6��l޽Xǂ:w�޼IHK�1=T��:��,"q���`a���ʫ�s��ul#Z⭮;	�z��"y]� �c�j�{���	7�Nf]�l��u��BC~ ��m�1x��s�^�E$bE滅��ϐ����c{�du�s���ۛ"����q�oU�u=ge�O�ǭ����&&�;�4���������豌�;ӭ�x���$)㢝�<q��+m�p��C�̼m��β��H^���oJ���f6Xaǰ:W�Q���Y���Y���2�+���~s��֯�P�vfⵗ�vR�,��\	��\+��ު�n��œ���m�Ē9gT��R�x$�Idg*�3�bXu�fGT��u۲-p����]��wq�ң��RMp`�Ç�>x1hR��˱\���Rf �Z$8����P���v���䜲<� ��n��ϑ/�s�c�w���ZRۨ�����3Rݖ�I$���j�m���<���l>��(����}�p.��WHݜ'�|�!�K���$�$�R���c�9,j���:��ҝe۲�pX����R�xְn/+.��	��w#�0kʾL���}1�{xm0�o�Ew@
ҟ�H�����ɻ��Mwl#<���e�3��k9���Я���Y�0���&.^o*��d�ʩ��6g��륓l���LE���M�Q�(\`����Z��gҳ{,��\߁CYB���؁���`�h����*�[�Fn��"'�-62V�Q�D�Ă̓Cuҹ!]���el)��tqx�)N�cu�gExݬ�c,v�:�^5d��ٌ�j�u���=z��Sɬ���&&u��bB1Ó��Ȏv�r7/:譝]�O�v�)+��cu3��G3�ד���\N����4����A�v���<;�b哶�"��N�'ٷξ��2W�CMU5LkK29�N�=�v.څ� �VoD9�ĳ��Ƿ��U��	���jOd���v�3����9~g|jfs�b>S�$�D$@g�X��Pb]��]�v�-�Z�"e�&��c<��ron����C���D�;lkxN뀓$¼|�tM�}\\�b��=s����k"ΩY�Lo]$<�y$�׀�VS�\b�]ڒ񞉳ѻL�7.��z��K1�U=f�Z�7�/�wr.��j�r��a��'a�J��q&#w�4VwN0�[�.�xz4޳�����m�$j"H�-���`� J�cR��[`IH�o�S�Z� -o]�I ��$WF>��L�4a�7Z%;���ew��I�O���d�:��T�u�*�Tܴ�ЗXa���Z��V�gWU�m�é�%�/��P)����m���iU-<;i��8퓏Vs�j-E?qөw�'m䉠�鷬]Q37��)�	#�	Z�ܮȣ���g�bfZ#r��4Vw8�1%!&�M��.��A�(�����?@˳}�ɱ�Ҥ/T0���m�O(�N���JG��ov�vb+]�u��ԣiy4�#ѹQj%���K�P��m�^�����;62��Tw��}�V����;%�R��p�ر�[Uqq��dL�E4i�~�m���'��\�~s�~��//��c��w���ܫ/�h�m�y���&>t�$��5E�u��=�a�xu�7��8�v[pn��gjI�-�Δ�"a��t���Y f2L�%�}��]��ONݻv�ۧN�=4Ǉ����Zu�b$�J.�F�Tj�V"�)Ժ.8�SJ�R/��G��}*�m�e�CEr�h��gR�c��qYn"�/Y��đ�լu�O�gY�ivлH���Id�}��w֮j��x����wT�
�b�g1�ζ1o�pY�읣e�i˯����
lQbY0�Ѹ{6����n�uWu.�ڽ�����R������UL[b��p������АtݬN�i��&�;��;�K8h�C3v�D��+#�ޞ5�<Y��jR������5[���9*}�2�����M��[͛g��g���8x�_:��.���hW'�[6�5�eb�43Y���duYhL�Ҫ��
�����,��$��Owv��V�-.��högQ9\��:�ػ*�h�5���3�9�Qt���p�s;x��廝@�=��9���u�3o�^R�s�^as��q�e�^��i�mz�z���1���ug�����tq��]�ŭ<w��x�Z9tE�+GKܙq;�W��=C��WV�HS�2�۽fVC8�����pSF�k���*JW{���V1/yV�m����X0�	x��p�Ɲڅ�(�z��c6,�:w27H�_��b�"��*��;��ǐE�Cy��0=�uC�1h���eo�"J���3׹7���ؔʝ�lY��N"�vv<�v�n�bWV[j��O=��om:=c��f�W���]L�׼!���5�	҄׬����74К"Ў�T9�|	 �O�#��W!��" �,@�B����)!4`��[�I�ʌhň�,a+H�CAJcFeF�S(��@�̂�sdd�1b�B Y���RH�;Dѐƍ�%H�-$&f#,�h�AQ�ˑ���DH0�Q���&Cb""1`�DlD`�؃�!b�Rh�L��!A�Ll����$RY6�f 1�1�����E)�Y"" D�$1���2	�����(K&�A4���k�lSM#T��ݒIB��1��Ծ(�#K3%%}[�6�a�k#(��'+��Qa!�z阉!�4H �A$��O��DFV�}��Q/�t�]�	ǖ�0	$�&��nu=��E�6m�	&6�+kb)�zt]�yqy����l��hJ�Z�x����)��<o%KhL��[�R2���兜�$�ށp�>�nt�$������C;�4�13�-�#I�.&!av56]������+�;h�F?`5��$��&�ue�k^���{5.y�_��%�q}�I:L�t��Ll�{v�jz�e�ENٱ�����f$�Uz�n[v�r�Vgt��&$�#�|a�7H�B]��f��!}���&�M���w��ov<��7g�����g��{e���]�T�?��㝍Ͱ�d�a����X���cŗ��ֲ�2��뮗D�(V`�:᪸���9��wZp˥Γ9��!�%�Ӕ 4�ӄ�oF�{��&,����]�&0]OH�k�I,�i�O�lq��۽�Ưf	'II���7br�����z��uT�Y\J$l*kŢu��n�f��xcd�`�I�GV�\�����t���[��*��z!���Ye���;5�2LI�I�c���0cx��s�wD�Ę��sw���
�V��(������~(D6��H�IO�W�T��t�����V�,M��]�������ǻ�d��׀˙���լO�9X�|��:H��^��s[M����.�Kx^�I�I�2Iwe�l��~�/�^)3�����״�z�8���"�$ޏ4�<_AaˡGǂ��]���7W�;�]^6��h�P�G��]�n��V곞�����Ҫ�GRkhX�n���;*zj����V�%�oP//e7k>i ����Cm�[4�q�#���$[T�l,�l��]�X���
��v�5�����Pq�C�=���9��t�J>5�pv����`�f�E��G�l�0�ZGB���Z�Ь�f) e�����;��Vz���u<f1����Ɩ[	�h�LK�*�pW�mڄ<e*�ir뵷1w�|����k��z�T��f��]��q8�wMq>���1���D05,BS.�Lp�o}��0Jo�Uvɛػ�3;w�����٦l1'�I�d���M��jR`�-�75Ƹ�c���F�z�{t���[ՊL!��,���)��^�I�)8ID_2;P���L��p�����.�N5%	'I���ܦ�bU�eR�	4��뽓7:�H@��ޭam��&���R��$�'I�U5M�!�y	�F<m����(F�黵�M��fgD���9v2��b��曧���BnGf��%(Li�G2�5dR뵮aY� ���5W�fI?�O�e��h����m.dJɱ��cV{Sz�{�'��C/7�M���GG�te�&�]�l`���F�R���/v�CQ���ܗ�v����mZ���b�ń��Վ��������4U�R�f�6LLm�;�-6 ��=��v��y>-�΃u<�H@������BI��5��mu�4�^���ޑH�J�̲��َ$/2�ާFFy�#|&�ûR��I�K�;/du��UX��\$�5�9Q�E�6��ipJ�������<�绵����cwX���ǣHo鿶oA��8������Z�v0I8�U��[Ye��y?&�kbˡM.7hV��4te땬�P�M�UN�RTA4���G��3��I����vM����F�-���a1;�=���I,	�ɦ��Ztc�d��s�w/�U>�k_��qɒy+k���c"�����I�`�q#0n��O]��3f���͚:*�"�y�,&�uY���-@�9zwEU*�}��V��95s���%3'4*y����ٽN��I$�m\ޚ�>�z:��}�x���JH�$����3������/6�$��l�gKg�B���bgx+i���Bx%���N.����JBL=)0pR���q�_ak���l)�u����j��Y�\Rc�R �����aYY�$�B�:uN�Ts��pYE�P=�ܴq��њ&j���-� ��������(�K��W���#�b��3��9�tH�����Iy&$�e�:�4\�:�+ӭ{�R�-��W�����}�������U�9U���cuH��	:.O=�rFaizˣ���𳒸	I���&	$���#�7�ꮔ�-�]��a�wffvp�h��O�{�Θ���k��d:3�2rr�(�;����/9L�̿@�#o�򷯲�]s���0C[yp�s��5���"�����/���7�IJX��_�[�J�v���I�_7%�*IQ&�ba�8��&�W��Dz���@��p3��:�!REUA�^�vk��sh��;��u�1i��5͊�+����G���N�L6$�$��&�O.�����V쥩����h^2I�`�{K�����Ov�0�`�yrՁ�'q�`fgg
��k$��;��y�Ná�7��I�d�9"���-1�ʜr���2�T�5��2�{;��� ]����u���ڗ���}s���3	�gi7i���R�*�C�e�O2h��+��]+���ݿ��^�v��Bq,��[[Mb&w�gnp�ݩ)�S��<W������N��zz2�N��hΤ���:�h�]N�ڭ���x�DW���`j�R�|���ɮ��
�<ؤotf�'P�6�Q��2-�jѢiI�N:�W���)�����\e7��z�@`�+��қ�8�<���q���nn�/pz{=5ۮ�q����O�M�ݮ�=[F��;lh�*oC�n3ڱ׮Sx��Ƕ�H�ȍ���piTx��.�:�y\l�鳷��3��]��W\u>v΃�d��I᫞�3��y�8ڝ`8i�M03b\Y��?��qbӣA��{kfp.�\�,��Kw�������^�g{]/�3Q�m�7#�У�@`V9�~>�� [�7�I��\1��+8�T�����,�C6W>��o��=vR���=�Ow6e�{���l^�Gq�7i���R�P���\����"���x��,k$�&�E�C@���]<��DL�=L���V0��O�$���q޶��`���~�M�qY����PcY>�i���w�ޮo$�����)����,�.�S��g]�ˆ����`�x$��?=o%��7�L�r1��X�5�Ciuڕ�f�Ֆ-�CP�C�3��,՞t{%>I����u�L��T�����~n��:��R/|�ܱ��	�0�^�ػM~�뎫�/���W\J��;9ZW�;�g�߷G�]���x����_��fn��JO��ٺ�cL鸦�v#eJ�eW�UW�՛[p��WƲ�)�}����.��l���21�/I$�;��1����z?��ڋF�SW{���V�`0I�Io2�]{���K�4��˹I�8�WT�ٖ}ɪ���x	�+)~�`t7�:]~c���[��"��ݻ�E��W[!�'Sg����ﮘwk�&.;�%X�cX��]�����"�yݪj�\!�pK,5�k��)�H������k݋�[�a�O�$�4){��mp�W{������h0x��Xk��I:L�N��qs;��e�[���RT�ܙ����V7bI��?|nh9��m��>!&�$ޏ'��g7�{�O#^>=�|�{v�[�Øv�-(K���&����)�,K�s)]�"�Y�{:v��R���j>�����+t��R�ԿT��&�i+H�Cn��^��ԭr���ḽݩH�LN�nH5Ug^�g�&FCnc�$�4-z���.�W{ʦ����p������V�	7�o$�z��l��ੋ��VUݩ71��fi�a�f��c��I1#����gM����B�	�T�`6�m�RWD���� ���WYa�ne�&�f?o���n�V��	'�Yw�?mW�ile.}zB��ne�m}��N6������5�9�cj�t�_8����.}
���{�v���(��%+T�t���
��
���y$��Η��B�S�d�m\��ɌqDfvoX��v0�o봠8/ˡX�X[r����)8Բ_Zs��v�ƹs�=uC��I��˽��M.�i��YN+ɗ3���J�&�ݞ�zii�E�%��
�@�,�Em���F����F��َ�`3$�&�
�:�4L���<����m�#bks��}��&�L�TW���NI~��UI'��%�ul���ǚ�+42�N��h:a�
J�T�(��I~�ܭ�B�8\F�0���p�z8�Q�QY�$�%\�p�uO�x�уۼ����/ڛy����m��JM��`��:V���L�xn7���'Jv!��pϮ��O]�Fe����&	0�I)9Yb��y� �z�+�з��3N3/;����潶�m(��{q(��0K���o0�Q���dS�<�[������:I~P����>\">�PV�b�(��?�� T>訂�[�p�s���y/o�ګ�-fZ̶̶�ՙk2�f�f�e��ՙ����k3k3[3Vf�e��l����̵�k2�e�ͬ�T�Y��R�e�ͬ�Y��*�mfZ��̵���6�5�5�-fZ̵�k2�f�jmf[fV̵�k3[3k2�el�l��̵�m�k3Vf�eT�Y�Y���kfZ̵���m����2�f�e�Զ̵��̵�������k2�f�jZ̪�k2�e�#�#�+͇�t�-fZ̵���k3Vb,`�b,B(�(��`�I"��b(�qel0X0DX0TX1TX1X7���``�U`�@1EX1X0U �  �@0\Xq�*�������� ���,*,�,", ��,Ų(�`��`
8`��"�(�*� ��
�"�װ�DX1DX0X0DX0X1X0TX�cE�Q�XTX�c�ٖٚ�-fkfmfmou�ޭ�k3[2�f�f�f��Y������m�k3Ve�e��l�l�Y�ٖ��Na�8��?�Y DcAA#��Z����~�������?C�y����Ϙ*�����O�,��������=ܟQ�i�=��������
���Ѥ����G���;�d��E����� U�{!��	���H��3�&C��a��� �����$���**�E@	dEAQcE�E��Qb�A A`�Q �XEb!E�0X!E�EQb0DX0TXA�H(��ŏXBX|��m��DDYdE�Pg���g����_?�`��3���� U�|�?g&?y��/�>��?np}Rpz����҇�<�a� @zQ {�z$�@w�.��
��Cz �*���,���c�����!n�&ܑ8/pp�8 g��{���C��ǈ( �����>�3Y;����<����������@Z3���J� ���0z9C��<WI�����>c��P8�&��dׇ ��!�|nI���Y��P.�W��n��T�0,���QT��0������{�y������)�����,�8(���1	�\                                        ��(�   ((�@ �R   �(  (	 � �P  �  �I 
�T S}�*	B�J�$�R��ID%HPH� ��T�R��J R("($�R���"R��%PHPU+|  �P
P�
R����+��
�vrU(�X�HW=�
��TF�U������
��yr:�����݇ �W� 4(O� � >@z y��� @/�(���
wY��AAK��{ n� �F���B�;�B�T�\��Jݎ��Y��LM�.S�[�P _ ����E%(%��A����R��w*U�S�T��4��=�t�T7�s�T�j��]���J�jP.���)T�zPK�J�7wB��7���*@�  ��o�c�Sٽ��B�ΩJ�:Q-۔�J7s�Kӽ�򐵽�{�V�G=**{ޚ�/z(�	D��)IU���E U| �| �$P$�J�H���}
�ݹ!;���Tּ��R�i�Ǩ���b�͒UR�eU��U ��y�U=:)��*���AA@ | c�J�!ゥw 7n��%�T�Kw�+qR�@�Ёn�Fa��r�ATP*@� �TH���A@E=�Er2Q\ةݺ�%��R�����gUE7n����W1��nܪ���l�  (��  }�pEN��T�P��}�@4���I�zPʞ�u !�*��z�O[�sĥU��L��	m� �(    ��P�R�*��AH�	C�}���C�qt��!Њ��t����O@�ۉ
Sw��X���հ�;�=z��J���E�zW �R���  �Ѿ�u=m�n��z���;���@rq��7����T�O@y��O{��R��n����U⡪~��*T   5O�C$�*   "~�U$dJ� � �d�R�  '�USڞT  ��MD��Jh���?����z?��$�jHl����e��M����Ѥ����$L՟���	'�V����ݭ�����ڭm�6��FI	��_������k�n������e-ͬ�lb�ƭ�Hͫ�B��.A�CUť[�����m����U���ֲ��Vj��$WH0�X�J+%�)�n^Z��%T*�;�tp�F��,�KX�$��L��o>�Ql��^d�ʕE�r�=��r)hb�P7%�z�i[,h[�����V��7����ʭN�ie�lb2����+�K'g��46�'{e�w�n*YM�݂���5��dr-��6�R*̱m�U7�mPʔ~�{{`�a��'f���oPaj=�U=���D�
��Y�&
h��e��e\��c���+i۲*��Z��$YҬ��+-�kp\�k4S;�OedW0ȓ�ʴ2�f�K���^mĕ��ͧUF�v�L�Pa^�݋��t$ܻmU��"�%%
��3�SFڤd*��y0U���K.J�R��7Т6��E���/�Ue^�J���"g��6��sA�휪"k�����ei{Y�r���ǈ�Y��Ѥ���Ъ�Op�j�y��^�l��7Ɂn���oڱ���Ńr�T���o*عz�j�G>ד)����r�r��s,��^����6w23�U���:;$&�Kh̻3`��M*��*`L��L��9U��Mfd�y�����,`�z�VME��JJe�9���z1�7M�PYܱ���������pV�M�7+�[u)ڗ�lr�5[�n�p��(���#ٺ R��W��n�mn����+L:��%w�ا���+ӽ6$ٺ����v�ѪäXaIW�,�:���B��m圫e���]L9t7a�{� �3�߲ԬR��PM�uP����c�i��bl�b�]n�.�h�n���й{�����f����ڍ�\*��:ލJ��4���]K��ѵ4ੑ��i��{� �ITn����:�
	f��wF�� D�� �����C/(˪6C��׌1e�VWa�5�^��Y,a�(���L�Վ� ����6������$��f����Ok�ϖ]�u[��[�2��;ZV:z�5��E[K]G]�TX�f�(\ݖ8��͙�[�D����w�0U9���W�2f[ҫ��CA��ꫂdE��%Z������e�7P��cj�f�yu���T*�$���7G^R͎`�wUm:�IV�V�rf�y��cz/C����Z�V:�]a�I"��;՟Y�u�J�;�ke�v��Yf�b���Z�^
��Xx7+Z׫R�Z�c+�rB�<�z%e�A-��Z�A�\z\��f�m�қp-�m�^�je\5�L'26��B���'T��j���QD�]�Z��4bWUNn�Ն7j��;ɘ�]�f]�Y�"��ͽ����X%�*L/B߱4E����s���%z֝���X��y�%!�	�.�ʸ��n�Ct�*3X �^YU��ǲ�.ء&�De��!uL�xݩU)�Ĭ�P�u���ɋ2
r��rb�cz�[��@�V�b��;i���-Uh��[�¤ղ����q<Y��2�n�.��C+N<J;9����ŕ�f]^V-�ƞ��4��Ē]5����d��c.�h�ڄn��ͻ��w��� �gFaۻ��q�ʳ����7��oX��VԎn�/�o���t[1{��T���m�u�tf]���	b�\�iC�/R��C0��o��*���M�4b��Q��)n`7gu�B�fHh#*�,,����t(�L��5n����d���F�ǻ���$+�{�O\���]�UMoc�t�uQ
�W���7�*5�^�%�YVlP���!���`�cF�r�*.�	���n����T�A1d�ܹ����q���Ʌ�}H��q���H�X��;���0�K�r�V]-'	5v����d���J�h=r���C(�l���M7P�Y(\)�����SUV�m��Fqn:r�RGEe&"r���wfd2n�8�ct���{�ݣ�E�EQS��	��h2Z�Y�u��0��9���6������΍��R�H+f�Ŏ]}�M�֏�B[ܥ�[�N!6j�*k�^�t2��,�r�z4���Mdjf��n�Y�y���f��ZN\ʪ��ꍡu3��on��K�ǡ�[dj�x�(:�Di{6I &]�3(U�D�t�k��h�5B��t�;KE34A4�1-���e�� �1{xv��b�5kuط�6��Jel�ٌ��F*]DwT�7>���V T�:�;kWM�7Iiq*A�8I�	ݲ�1V��ãv˙UN�k��U��VY��(-im\�BΣ&�:㭹z�[_T�z���e�bȳ2G�E{��a:NȬ��W��E�R�;�j�hvF����y	ݵWU�W�B���t�c:�Y�1#�)�ݟ^�4��"��˺�#��Z�`͎�<��^:M��,aא+ٹYWWgp��ySa�.��L�nd���	�zLi)����UL��JFlC�uE���!�
"γ�6�v�.�w�]�-�m�����n�EOn������b����!��*���&ޝ��i��wj�+�y�h����9M:�E�۹�r��DM��&�h�u5���	�l���V��l�0:f��յ�X;7 ��%֪�T��f���n���Xf�bKyVt^D�����.c*�;Y	*�;f�cl��*��ϰ#wj���d�YB��WOm]����Փ�S�ʽ+Q��Q���r��LÎ��[B"ku�V�
r��v˻K2�-�D�	�Wx�R�Ksl4Y�z(�(��3yN�h�&��Rįu�S:�F���L��:���Uu�0��[�����r
nJ*�3^�R8�e��5xj�ip��ܳ�w1�1;��؅�ow*�B��2�N̽����/p����InX�Ӕ�ҜTl�z��{ZUE�j鋳
�(yO	d:��'U�ٜ3���<���8v�P��e,�Ni�f��m���J��ß#7�iaz��N�cr�[h�V�uT�̬̽�U�ymڼ��I�&��/�`��M%�.%����6�ύ`��2��b���o(P��*<�6���U�)c���xʽ�yR7Y�Md�)�u���5z��&�k�(<ƴ"�+e@�2ݵr���ȵ�����Ŵ���1��n�ՋU�w�[��xlcB�SAZ��tMSU���.���w2�2��Q�	��u�Y�=;���I�jn�j30��ͦن����Wl��P\uYf�x�KڭX2U3��JD�j�֒v�J"�W�fM���RT�����~�K��/�iԝTwWҒ���h�ۢ�^���[F���a��*���|~e��Y`�f��s�(Y�+T�I��V�:��j��^��ڠ��"Nޥ��V�A�����x-`z��N��;��T��E���ޱO䵤�`�[Y�����5�3An���.�[�kǎH�#\��%	w3�cau�p(1�Wv�%�G�[�ckh%G^��&��+b*�h�y6f����ȍܫ��ٴ�XƜ��%�d��Q�T�ڙ��:�+%��m��A���AfU�Z�Lߝ�,�E=���h:�pm�%y�ڷ{�1,����nW��s2��n�@��1��-�PsI	
D�༃f���F��i�6v˨C����.�|�GM��r���ݪ��]�j�[�*�^�XQYPM9H���П*�����娆���1ne�Fj���Cj�*�v(Q�י����KͽX�3.�a~��-�R8~Ge���;ɖ��'b��G���:��oP��;-IF�8sX1ঌ��&c�E�^E�kvf�Q�����6)z�1[�X����Ϋ��fXl�n<��P�����Z�pe�ŋ[���v兎��R�� ��ưP̛Cekw���Dv�V�R���+weL�r��<n��	Z6[����lU]}�Pu��.���N�QT�B�6���w�c.a�b��P��4��A�7w�ܛ��z����I�i<,cPa��8���t�hO^�jt�S�E-&c�pRԝ̺y��	v�X��2=��T˫S%�J�Q�{{KZ���s5�:�^��G"M U���f��y�U�ɨ������ijH�4Z�f�
u�Ns0U��Ǚ2�[Ɉ��pʣ��*Vkp�D�+V¼��h����k�Ճ��'D�lVU�Xʼ�v�m�v����r���h��*�sL�aZ61a�4J{��I޹Wx3im��+��.�W��6%,�����Cژݚ�C�"������^eYq��p�/kie�7H��ݍ'%m��ٙPF5�M]i�X{���[�=�T�Yw���T��uJ;nXU�f���%*@�l*�����24du:�#}��aF��}%r����Ehxɪ@��Dk5Ec`�Ja3rW��kh)��'	�J!�[���I������$�&
���TZE�S��;r�[���L.�fʭɎe2T�n:ͻ�ٲ�UQV���uI����H�s]D�˽��bS��(�$��ķiA��L8����f��ۼKe�MlK%�ҫ`�U�Z͋\ͱ��Ƚ�T�iRb^f���ņ��ڢmm�Л�ƶ�d�Ww�QXmY>Û��V�GK4mfЗi���N/��ѽ��&Ջ�T�;M�$)�.���ee����lô��ۧkʻR���Ş�UU�*Uu�׬�T��1 �2�'v��7{��t,4�G6����f��0m�QD�5��,1�;��!�o��НIyyo�I�%uX��&�ᒎ�����]���0K���wt��YOQM"vj�$���/lJ5[��DF���'�˙�r�}G&�n�QY��y�h@�1�^�Ђ����,��C"ׯ#WM�Em�gsL��6ю�b*����$�ʼR���̦.].]�2���x,��((J��ժ���P�Eч1c����fD̸�� :Ujf7_=�P�7����K��4��]QFS��[L]k5���6�f;ٗDU@hk�*��k������3k��kީt/m�	�XP�*.�5I����ͬ�W���FU��5-�Ɠ���ٿ#6�lؓ>��5{cHגm��X�2��1���nm
9Bi�[p-�Ѹm�Q��7E�J�`�[�z�ͼt���A���7x�+\,�t�Yڛ�����.�����D���J��m����4�Z�^���Í�,UVX�J�il��	�V�h��X�X8%�m,/*���.�B����e�A"4eH�c�H9�+*c�"�$q���`�U�Z0�S/R�ٻ*�۶f5-۽יCcw.,mVY�˻�Y�7qJ)\�1*�J�N�f�'�t�|\��Y�jGqℹMc{#Hڤo&��ڕg6�0J�6�&�F=�Y��YfC��B$��p�#�*(v��l����DZ{�*����Y��WF�kc�薑�kN}���ȁ�]�n'�Y�r֌�r����h��4�0��(��է�B����l e��ܓ4���T�[�{N�^c�z�5TbYR��,F�C��S`ö]/��e�0�.��^�ZE`��z�@�I+4q�W�Td��ۛ���y�[��K鱺{{d��x5ޤ,j2I���n��΍ב�Q��h�S3x4�f����@�z��Y���b���F�2�A`��ˡ��������s*���NdH<{gr�ˌ���Zv�٤�b�d�&TڻwG���͗n���EO�i(�m+4�����G1��E!QP��&�׹��R�!Kn�u�ֿ�4�b̍歛P�SU��4�v�H Z��u�3��3FV�nѳW�U���Gf��JΛ�4v���L����q��7LЁ$�ff���n�:2����0��ޝ´Q�=��hT����k�.��s\ͅ�B��ں�^�m=7%^���a�ַ�s6���ƫ*���1����*5(k�Y��E�('Z�%��LKfݍM�iBg�v�%=r�Uf�M^,;�F�u���ն�da�[U%��a2^B�AZ)�t��%Э�utv�YwѲ̪�J,�8����RM��)�=�*^-�ۙRkI������6�jY��X9�͠����ܬ��.��N@�D�W�JhJ���mӼjRW�+VV�0,�D#�4Q�t�Q�����֙)d����:��seӫJ�-okuQ8��n��yr�mK�ȭ��(�ցK4Ewi�3c�W�&*���b�c&en�'Z%n�og/Wc'k+���.�����T��b�$L�Vd(^�f-���*z�C,-����k+b��Fh�l�W4�q��I)E�3x���X/l�N<1T̼�r��L�V9T�z�ɛ��T��:�A���ܵrJ]�V�ck2^IN�޺�f+BW�k��d �4n�܁�X�5�č�ڹ4��OBͼ�JV�P8��#MC�%-v�aH,�MF��3*�/j��x�V2A.��0ʵECK+*Se̶�E�m�cթyz�O5!s*��=wVZ�����0(��T���&�YV%�ߞ+��{J6mͭ����N�C���(Pbʫ��L9Sܡ��k^���`XfVD��ְ�oV��o�N0bܑ�{l)�%\�w-V�uDәa�Q�VR9&�q
ۻJ�n�6e�̣Y����Z���@��#6˼����wZ,��`�xH�^��D���R��m�ui4lF��Ӂc����1c�嶷~4�XkRuqh�r��
��E�M��U���0�׃UA��V�b;&μy����D(��VltC2��Tk`�F�UZ�Y�x6��˻�k�5S%7UN^n�6��ٺ��j�cde��oU�x��Ǘ6h��&GzlkY��c7),���B�Sq�������ݤ iV�nU���ł;���3(�ذa����3kL56�:��T�������ln�&n�
3���jYR�K�w0�ZNR�f��5J��n�M�N]�ɖr������˩g6���U��YJ��F��Vn�5<T��p	sn�J�lBr��g̚E����ֵE[X��-�Z��+kF����ڢ�QU�6�X�ձ�m�j�Z*������ѭ�U�Z�mQ[�-�Z5����c[lZ����Z+V�k[F�֍j�Z��mQ�����F�m�Ej��j-kV�mcV�-m��ыQUh�Z5��kE[Y-F���mlUZ*ѭ��cUFڣV6�ֱ��ŵ�-ckkb�kk��-kTZ�5i5�Z���U��h�lV��6�TU�F����b֍VƱ�k-jƫj6����cEm��m[Ql[�[kE�jߦ��	 ���y������4~_���r����'�dS�Y6[[zj���Y|�w����Sk6�ʳy��_c��m�v�E.����<짖�IV��e�W�cS�t⋨��8H��f�8�r���V�pƔj�q�ʩ�}�*�c�*޸�3»N�N<��X�Jb�P�yR��i�u̓�ݬy��+�ls]K�k�a3�er\.�-��m����J	��B=�c�2�Dm�����a32;G���r�-Q�[ۖ�f�Ϋ�t�k�1t͆��,J��bu���;7kJ=�����]����nV��Vt��e�Z&�7�����^����Oz�G�ڷ��wom��I�[6#�L\E�n��VFlUuٝW:�z�J��t��=�-'���M����@7F��_V&��Ư��ث9 �fІY*���ѹX&'E��_uM�j;�֊�zJ��象Kv:��n��9�y���+��훤��n"&,��-6f�f��W|����M��?s�'6����l�	�c�p�:˂rb�,��%���U��Wh�7Tr���"a�̕6����VF�]��W5g7����u�-L�YO%��gE��-Nw��:�n�Q�C�����]Ua�5R���W�wF�i#Ua�Ǔ���ͮR��",�'����76���,���<n�XjC�6��G%k�.�+�UK�؇Ot<6��
��)�^�n!,�������Zůi�N��ST�Dr��Ώ^��	8}��GE�Ƅ۸4�:���[m�`��z�.a�z��BZ���� ��ėx;C��leR��:�:�{Z8�Kc���]����a��Q�b7��4���#}Y��죗ֲ�7�!�&c���+*��}��o]�o��p�ɤ�I^o[g�K[�]E�]nWVjܠ��B���ӗ�Oj\���Q�'0m�&��w!6ճ�p�뭡�Ma�лsf�l3�]���'��xWh;,S�H;vn����3����f�;���-�����ٴ�V"�m�5���|#Ŷҵ�TZ7r� VJ�wdN���V,=�n)f����s+����w]��T0%,nm�zފ�yY�Z�����Sã9���n��8�V�ԝڷ);+y2�ft�ɬ����8QA��iQ*�u��&r���F��T��h����U����wc0�Ƴ����r⾔m��caӆ�������+��aŕ���C��s#�%��yz,�g79��Z�\��ʠ�t83kw.���+�ۻ��Kq��8j��	�o�;��J�]vf��cFB(�R8�7��5�H�z�@pdbc�U�(۝J���y��1���p-�����M^n�U�5�Is�6�>��bۮ�&���x*��^��m�Q��L]`;P�̬
"D��r�;���*����kG[s�1
P`�;Z����������\�J�Z���!�x51A��殲��]M���]L����wkZ[on����GQZ�
T7.� Jp�N�Mi�b�����k*j{�Fi]Ugo2����q�ng��U���B1p��k%���۝�ܫ�y]�0�ݍ��U����&Aֲ}//�E��7ɓǳU��rn�9�nv1� _S�a�T�q�|&�lZޮ�Jʗ./m���Č9�W�:��Xf#�A;y]Y�%���Pn�{u2K��1���yUJq`��N��è2����5��4CxԹ��9�Vյ��%�����!^�K#&֓�vN�z�
4�]Wv궶���t�š�^��+���=rv��:�W���)k~�T���uP��aZj�J�VnVq���
+I�(�Z鹻Mj���^�[���vl�A?U���m�Mj���g���Ʈ�����2_af�4�=ڪ�h�ݮV駠����ϕ]�A	�����������϶�i�r�F:�JI���՜�,Ӽ���]QfP��N�b����ãpXܛJH���2M,%}���n���V�̍܈��W�FSb���K��ͱ9T�v�e�,�I�m���wYq�j�~uj�M�p�5snRU�Y��3
�/�y�oNeelr]��Y}��9[��7o+��n�ٺ䋳�*a]d���*�PǄ�y��TAK�uEXvg(uY���N �.�K���j�钶���Ni�u�՛�-Z)�=�&J����*�|2�d��gx�t����*��|�H)�À�����dᩧ�J+ܱ�%n�yhX�b�_fg7Sx�u�ӽְ�[1K5���g�f-B&A��N���n��Z]E3	�E��CQb�$��=�XF�J�ju�9 &WY�3PR��o�Ȟ��Z�n�,��kBk�<�E�
�Z��h\UY���=�J]De�d�Zl㻛b[�[GJ��`�]N��E��$���Tֱ���s)��e�DӦ,ޗ���vy�*w��ߣr�컰^೽�u�~��3������踓62�n�ń+w�Gb�k!�M��Xb�l$���$��d�;E)��5lp弘�zm�e���m-�\9�̪'opn�kn�ne:C,5Yb0���TH[�Ub�-^VMk	q��.�I�̶^fc�Ô�9�Gj��u�TT9�P���S�*W.܈��r�ux�nf�pt�F&e�uuue[���[hq͓y*�A�hUʭSC�5�+(Ay�s�Y��u�m���Y�k+V�U*X�ܚE�_^c�R�.�'�]0�jSt ��"5lЭ��uP��Ut�3v�,�yK$��Q�u��5b�+�)�!M���r]ev�a����5�y�馮���30h��5̛�1�EUe�{��-;qo51�F=ܽ�6֋�R�"��9����e�u|�^%�3t�<���Ї���Rv��U�6r�f=!�+�oȞ�M��[�l����-c���g��`�Zrne���]��O�n��Ql©�X�m��Z��!"�l_��ݥ�J�G�5ƻln�2��ުc�YenZ��r�6`(���iK̪2�3!�������V%�h�5C�D��|��c�hDk,�Ǻ�˱k%��3�]ά�y��WY�R�*�3�g
ٲX�2�n��V�"�'m�Z��wk���^葴:<��.�p�%�0wLL*�CLȤ�״�W��i�өBj֢�䙷�s	}V�-�\��b�3l՛}2��r=���t�7��F��ܟub�.X��OQ9�J�f�^�U^�[�Z��Z��mޫms���\���E�=g�W�y��l�w�����Vn�E3�q����fX�,
l�C��j
�6�_�wV��:��4�+�ބHqEL��ז�rR�Tp^e4ٱ�yv8cz4����.���,n�]�2���,v��WbO��o�ta�����%���m���S���L|���2��⏩�j�
c���J�j�w ���x8ú֊9i�yqp*�ecs*ޝЩ�WR�
��Eh��M_֕2�ᦵgժ���w�9��"�ʫǚ����i������jU�E`��U^Z���X3]��l� �d3i�}�lp�Uq����:}f_"4�6���J���A�-���(�3ЪŸ��.����<�绘�]Y2�Q̷g;/.����o����R�ޗ�* ��v�U�wQw��@�����"͛�Ō-8KX�*��4�}Y��Mf<��T���v��-T,��1G/*ݺÑ�g���wJoiW$���S�eeQ� �W��k�w)\V�x��]ΛR������v�V�k��f��m�ww��j�z��9F>�5�e��ِ��8ǣ"��ؐt���܏�T���W�^\m�5AWĽ�4Wncۊ`��G�Q�Qp�_ͽ�Ys.�8�ޚ�:x;�W�G��h����}W�_nI�1�]��������-֚�[�T�G��T��)��q�����.b��eec6k�ۢ�nJ�������"�ٗp�����ݹz�Fܾ��f
�M�ʑu�/s�pGYo�P�*�nq�38��ņ�fd;���:d�s(�+(�V�*�KW\�V��΍���B"��+�ݙy��i�ʦuPܼө�%CR�S�%ѫ�j�K�����=m���1��Gu��UU 7ٴ�<7��0�0<z�E���ՇV^(S�և/l�z�N���؃;�6r�UG ]e�b	A��#������􃃱��S�I���mHIЖ؏0X�%u��4V�
P��wVi�Q1v�R^L]�Q,Uhm�U�^Sr��]՝;��x�D��=H�Y������闘����ܩ�h�&��ufZ�+�e�,r�M��b�%�F���6r���Gr!cm�*�a�4���b����ƺ�j�ʔ�]���[J���st=<�Lf���U��	�.0P�ɽ��.�+t�uf�j��vXx�i����K�2�ѝF�-���v��\4�W�Q��ڪf�%3��X�`d��JYj���괌S��5/�������.++91�wՂ�b7�w�Ҭ�F	�w�aQ�����y�N�:��!�WK��-��KZ�����m��R�8�g[�\ok`Y;V�f�cv�;`�<7j��.���C�m��Q'�b�+Ϯ�pΧ�FAλ��V�j���Z��C�rpb���	��IP���.���#\�6t�]�/�񌱖*�w�h�c]��Ϣ{�����j�f������Oo�n��*��#T��=s�1�m��^�v�������8�h�7�V��y�ef���U��]��c��Nh�)F�nT��e݉(�����,��G6��YUY����ZTC����9�-<S�ڬ���iTz٬ �,��x�#.v�m���T��&�m�����3�n�+µ������X������9��Dއyj��e]�^�ӕ>��Z�c�WI��E�Ս��U[��ژwt��.�7`᭻W3r-ɯI�}�˵d�og.2쿨l�;��n�1[F�MWt+��a�%Y*�\T;#�5)U-��{�8ָ�2���#wx�X���6���Gn���f�2���XK
�2����E��20M����\͎�ں�n�U��
�Vw�f|���<�I�͇Y�����X��M1R�Z��i40�gFf�XlL�\+�Om͸�U�Ev�e.��%�[I-�M�Ybp��DA3z���3{Ki��F<m���v�c��M��j��B#��H�$2i�8���3/r�p5��f��5w%�j��{u��y�un=�̦���év�k��ӡ�.*r5ð�
z"�B��W�>�;�j�;���pЋ�ƪ�ܻ37���[�Y�;������F���|�aw|ܧ��I��UC�sqO0R��IƔD�IT���;����sM�bM�d��w��j�`��H;W�����������,nn'*c:���4fL��x�q%Z"WY��|{�FQ�e�sUm��]f{`�j���;tL�_+��� Wq�B!Sz��V�熝<Ϊ�Z���˖w7�}6�$Q�m��2�W�)��"$>��qޒ�5��}ֳ��]�S1��*�MR�V�yVdʕ��7��}�8���5|B�f���CV��U,�dy�d,����mV"��*��
���:���=5£�ߤ�D�I�w7L�ܗh;[�͕�|��ZC��ͣHcB�gvm� ���-��7��U4�_@�]m1��2۰�*:tͦ��WU�x{Ρ(d�TB�
Re�o�)󾼪�s��`�'���㷈J�7������Z;r�䅾���MN؋�I��8���n4������8�������ڃ>�	D�9�k�>|���hx��mu��#Q��ݭ�E�5�%m��ʧ�3��oX=�B�*�p�1�\����mf>�7H_���v&I�)Y2�	�#��u�*%�z��{�[�0Dw�н�������E�/Ft���nc�tv�89�na�5"��7��B�.kF�`��He(Gʽ*�K������O��o��pv駘):6;�QjuE�CV�/C���^wb߯	�@��mI�f��yC7%���k/#FT؉�K1Ee�q��;A��Uu)CW�3�y��+��|V����ZRˇz�m���\����X�I^,�9f�ª�6�&*����:L�z�x={I4;�
<ms]e�;/]^j���;���Y_u�:+z�m�4U�+Gv- �����ra���?WeyUB�6����l���n�;qf�n�wm�6Lg!8ԣ����7�e����.۷"�o&�(�kR�kz�]�N�vq,V�.�rE;��H$���U�.�rZ����Z�$�Q�r���w2�Z�hW����[��C�wr��|OohHL�zW��\��T�bǰ�zfvHu�;K��u˭���զ�d�����(9Z�����������[�}.����e�a�7vi ���[U(=�kwC�ׅ-kq���eu�拨����������"�YA�E[4�<ųx� ����,�US�x.���E��GSdkp]kW�}˗P켯�4�D�6��֗�أЍ�mlt�;�:��ޛŊ����!�����U�u�rd������Ԕ	�s�Cn�ӽY1^h��Dc�5ʴ<R��W}6n$���ݫm�Q��Fvә�t�?S��O�6�:��b��}*��+LFʹf2�+�e�"�W;n���Xߢ�-�jZ���3O�imחXIb1�z�.jg^�󺩧�F2�wU�د{Kaڬ꫺�=�u��[��)Qf'�	W׹b��.�װ�F۩�,T˪�Xv���R[q��q(���=��t��'yLYWr�ze�5�
����Q&�u����+W�Y
��:�ՉL"���U���Y+��͘!���c:e6�+p�/4s�WI�nj���F`��4-�ӭ8֨�O�6���vi��^�9ժ����k�vz�l�J%�BPC��Ɇ�l��Ӄ����c�k1X8O��Q����w#�F���������>���}�I������Ϧ�L�meeJ�F���d�Z��Я D�{��b�qWq��BJpղ���x�]�:R���tbN�=��N�Ѳ����iz��ܑ0�٦�`�85t��]Q;4j�>7|��T�f�wٌ��%+Nu=��-Ȳ���#��l�(��[�����5�B@!$� �~����f�SX�LGT:�U9p]�rZ�9���[P	����)��ω�|����lt��1�	,`e�B��7-��:��(�i#��<7:�Ml�Jp�����X]x��9v�mccL��ga�ـ�HXbY�Xj�
�ZB��݃Y[2�Via��Ȗ��W��M��ܓѠ���\�`�ӢRP���渌�V9�L]6py9{/	��f�j�G�V5�Gn]O;�=�.��l'4,�O[s��E�Y��GC���n0;�`:^�ٳq3�"�>n��N���)������)z��Zh�R�$.�������uJhH��s����W(�t��Ł�;
6��؃�kYf�j�Z�I�.S���t)Q�T٬��7n,��m��3V�Z�6����!�R,(Y��;g��'���:�
ڶ���J�*�n��!���ѨDt��@J7L��n[�q��=rs��e��KBVX��kx8��b2���fNv���8�D�f��2�\�X��WXqs�f�ێ]�ᡴ\Y����C�;q�ϱ-�N�uhۍ�35ry�y�[iJB��B�]����3�-�v�	���`�/�-��EGnԴ���f�o	�`W-�%��JW�.1u�<�Yucq{���$I]nl�X����4Iq1�v월��=�����j�y��]��ǳ�2O�$|��°�q���XZd�&���沘f�CBD��a��,��6�- �j�h��K`�6�Ll�C
v4N���)�,��k��]E9۶S8̃a��Bikf�F�l��1�Pis3̸�j�$ZYpf���k`{rt�v�����u�v���2wG�xw�M9-����SetD�Fl�qt"�&��u]#�YL;V�61���
dX�3Q�j����C��-�a����!cW)��E��.��+ˁT*���<S��q��X7<�����n��N�6ј�n��i�ۀv���2fb^P�ɤe�j`�y���M����)���*�XYn$:N���`��c�@5�A��a�
��J�-Hl�Ws�9�X^�,\Dq�݇�}|���.��Ϙ�p��ҡb����C%!]�A�d��x�r�Y��g�`D�:�N5sb�{n�K�jI�!�N�^z�/-r�n+��3ŵ���\�-�a�\�P���� ��k�͈K)�9����-g�2ח`;��p��H2!��|�|Yˉ`C3\�K��`	4�칺Qf��ݮ�@aסИ3�v˰]m��Z5�鳇�K\6�]��T.�/`nx��@������tݝ�Ě� Ę{3`	-��	`j8쇬��|���-��h���T�6Ũ�J�]*�.��:�$.�֌�4k�ȗ1�l����љ&�����R���յ��nN�V��K����6���#AL	Զŀ��Z�\h�Ij�1����5v�5��ѫ��9O 6�cuj�'&��ܜ;���9��7Olp��YԗB\�.��^n����m���bⴃ�c�����"@|��\p96���xU�s1ρ��v.y���{c#����:7�r��AhS���խ���p�������]n�c�ӥk�9����ęY�;�%����n��;5�d/Z�1l�yK|�#�������.]i�ƀ�.t۷J:�����En�\����q�nӷ	��2�rC��Hm���ucW6P���x�=�DF��zlg6�j3m,,̽�DZ��Y�=n/P�4����s��YN�����erW@��.��<km`Ӊ�n�"��9Gh���m�xL��T��W�<��6I���v:�l�-.͔�-�K�z�Y:ok��s��=�X-�WC4���u��ע�κ6L�����C`���Sh�1�qn{!'k,�4"��uք�-��L��c�vt��5�)u�i&Zk��-p���FV19Є�5��ffܐ��e�Vf$�u�ֳb�6�6�c{R/<'b�C� a�����랸��t�����XH���iv�N���+�;e:$�c �s�m��nv;�k�p,n6�crU��H6�gV�QCV���[+��� .�A	�6�s���KW�Y2v�N��*���G1��A��aok�t���۲�.A��h��т�������6%��`�GaˮP�8�*W.0nƃvv���C�\�R�\��[k�5������b�����y�\�5��Qn��x&�GZ����t���:�ݠ�*�Mk�%�e�zʮ`�C^m�e݀K��8;fZk�!��ɋ,��P��M
݋56�l#V;^7���
�u�Y�2r��Z�8;a�^<��;�qY����e$��f�M���k�a���'��%�i-��\�0��X�х(l
���JY�ghY��XK��b�6X(��7g�|�ƚ��g��\�s&�݆�d8�ɉ��H>M�j���,\hf�eZ_7���u�5�u���˒��e�n,�T&5��d����R�-��in�q+��_[����8㕖.ys�&w6Gl��\Y.�k'mF�$s87h0�x�3�K\u��� �4OuX�ֺ��t�&ļq�N8�V�]�T�	��l��)��qcer�����7Iu`�2\vq�*\ �d��pnps;�^�]���1��63W�r��hɋq4�e%�7L\^��\���xn�&÷j�l7�;���-�'Z�Dt.��i��-X�۱�e����$�9�=���祺���r�:7$z�r�t+��k�4+A,b�f�wn����u�ӀM�m��]b{7��8��z�h��n�L��ذOZ�c���D�2�8,���'hvӻ���^k>����N,]�ln�r���qٶ�n �EC��9H;zV'C�%ƚ$�[��d����wAg��Z��<�Sq�b{c��<iq�s]Q ��c�z8"�u׳lA��:U"J[��[�������5��B��`��c��Rg����nuI�;:h�[��Xc2\8ۭ�����ݼ��k���u���N.||��/��LKi��fMlKH�ln��v���(�j�WkP!��y�gĄ=,���]��i�lvwd�lf�:��S���U�ϣpJ�a:n�7>ٶ��C&�=�&���6:Z�Y�2�l0��)X�j��ft+Κl.f$)5K���G�ݩ�]zbE��\\��n2�`פꓝ����ˇ�s/N�\��j��\�������.L���T��E�Ԙ���_/1�Yz��m�<�q0v�6�i�G���.e{l��v�=s��k^���@�wn���9y�gx���8�B�,y��n}�n�f��c�R�@�m]N���c���ɉ�h��9���6=A�4�.��)+��lr���W:ݹ*y�Ͳ�zLXf�M��[h�яh7�Й�A����n�9y�G�7k��7q���uE�VH�F�]���p/T��n��^��(�:��I��v���m<ڛ�`ef4U��]�[M��a�i��{`kh�-�p,sa�Ұe�y��M�&ݸ���-UF�tD�iG�S'V�ķ<Pv�+��vi��\�fN����.�F�d���v��ZS{c;��\p��6�Ұ��6+�,W%���uڀ�����-#���!��::�sn���.�8�]n�Pu	�KX,�LJ��mK	f�X����hv=^|�Pu��vу�kf�F�Г�.ۆ�S�s��Њ���f�,��a���n�sӹl��#x��冨��q��Հ��E�Kh��s4a�p�ؼ&�����g$�.7<���L.�P�*lc���ᘂg�`�Ƭ���8�T&ܽ]�ػq��=d��X�e5�=m�ٮ��3��E���ػx(�_>,����� ���j�;v�U��m�s�=u�&[�V� Ŵ�5��n3�Kk56R��b��8�N��qևCq�^:Ɏ�b׀��^�i�R��`9�3k���]�u���c�Y��ѵ3+1������_ט�:���vu:�h��\֙����������F>_-'�v��䘅��-is�����%^Ps�����05iqxFա�iу�	9��8�U��oc&��upgh�G�$Q�J�q�L��,Qv�0�nYk���Fic�&tH�و!I�^F�ֳ�Ѯ�8��1�8��!p�vG�"�^�k�na�7Q�:�E| ��.�l�ֲ��!dV���a����XK3&�%�z�x������y�h�vl%�h��ZH؈�m�fA{��cM���++��;y;v�8ɂ�'���\ZK�bY���Lbj
%s;q�9�0�nQ��9��g�����TyZ����n7�шv�����,��b�3��� 8���u�c�=���O4u��gn�(�g�����5�\Y����W=q�8;���4E�q�5p�x%]V�d�WX����W�ǜP��������:lK1(�\���Gc��x�pJ��7���kq�.,r�NO9�$�6E��m��b���m�ak�z&ε^ �&]I�0ܱ�k��Ɋ�z�&5v�k\z�z�l���$]�g��xv��I��%����m�'�l>.��;�MycZ� S�ݞ�N|k�Q�S��ڭrlnm��4R�@B��AA�F�Bh�ԍy`���kn�<���ղk�fыRG���DP�[��X�K[�1۪89��+�Ϝ�Ϙ@q� ��q����\[w=a]MlT�k�[lI:�E�c�1,"��}��Y��x��vm;pal\*L��my9�
N;&��۱'â޷|�#.�!�Ime�'Sv��7e..]�Du�u-�U�e3�yHd���݅�e�7Ֆ;JJЃ3e�4r�.�ZN:K��v�0�u�u�:4[�������S�/n�Mםy�:�h�X�Ci��6\�9����Zթ����cZ�:��u�g�b"�EF*��,���� Q�1e�H�2C�E�&d�a�e$a�`�R�c"�Ȉ3)(2h DLc1�&M�Id�ɉ�I�HJ���Ic"d��0�R���i!�DA!k&�F"#w]�Q�)F�Y�ĳ�$F1�H �$a�\ɐ�H�,�s��,���fF�QQ�F�I���T��0cL�h�@j*'up J&D!�m����$�Ad�h�3#L�4E���M$�(�I3F1�E1�ZD2�1��QHJ�:I$�|ȓst�f��Vˇr6L��]<	VM���u��񞝞�Lq��MW��d�l��d�Tkgc�ڞ��8{70�u���&�K�v��YU��MhLF;Z��I�,�L�b�K�4��k\%:�f:��a-�����V/g1��iv� z5Ĝ�;C�B��йuH0��MͩJݎ�7a�9#JO�m�����q��i54�G$8�i���//D����0��v�����0�wXܻ�(n�c�sɻ�'g/l�W�m����� ������[����{p؎+\{�N�ڎ��ֹN�Ɣ�H�Ĺ�F��V]������/t�uAt8������1<�v�n�����&i�1En4��"FR�Ζ�[��(�n��ۊ����f����rݹp�KH��c�|v��qu�5���\h�d;���ǣ��`k֐�;cv:�h�uj��q��V��t����1l=����r�p[GFzS�����x�5�cx�n�B�t��f_����󭙂����y��L��n��G/j�a���r�e��5�K��%�v�T2��\�nqV�|�;�j�9�p"�#(�	G!P���M�E��%��IX(�+='A��y��q�n�]�r�Nx�]F�˓��M�Wh�G��;�n8���� �'�/v�s�H���W<sV�y+yW���AaE�0N(�۷<��ט�s���.b��Ѐ�5��z8yE�y�Ӗ���z �8����'n��{]����[�SgR�s�����]�\����q#>m�'oj��l����]I�n���R���i�
!h�#��c��ј�j�=�i;ї L�X�[Ds��� �����ۘ��0L`�(&�Gf&��w[su�Am�r�i�bz��m���*���M�뷎��V�w^��nS�<n�S��jyȨ�\�fZ�JxT�5��=�=m�8�
��]�t�I]֚%��4B#Ռ-� �����!eo
�F$-����Д�J@���ԶT��G�q�Ʌ�"�;d6����6�V��5������H°�--V%(PE�U�i=l�@e�F��#c!yP�l@z�F�-��#B�HQHв�V�A�����[��u̓��<g0�y1MhW,[����J��uK��"���e�}=��{��z�Av��;w�����~5��ޭ�̺��;�=�W��@�K�ŖQ2��a}=�]�j�YA2^�G)\����6�}n|p$rw`���7�q��ƀ��OJD7A����5�LcB�4�q-�u��/��+��oYgܲ�{���ݶ�ݖv���G�� ��!|{� Ct�̫���:�����}uđt�t=���1�_w�/�t�YD�@�K���J�v�0xɶ�5Kzy���jW��p-�@��� [�n�T��X6��]ƍ�И���!�8Kqu�:�� !a��$L�3U���4m`���� >@2�?6���J�;�'WN���#l�޲%K���2w�<f�FǙV�v���X��{)6���\B�p퐁�)L��{׻�1��4����w+T���]Spp��p�&)Ϋ9����Z�X+I�(�^i�[G��P�V����~�CΩܞ�kc�m��p�O\O��D��kC�U�ʀ����� �Y@�A��e������+�d�y����z��;� ~=� �q�|Am �#��b��B�����l��C��9�uY���A���AÝ�J4m�L�3��A,��� Kt �鐋t[r��93HQjGdGV��kc�m��p�����A|e����v?;��ov��eag� c�X���f�i2:e		��iLbh7]2�a��U�K�ګ���#����w����g�F|��/q]��S��}s�=���y������!ޯ�m��_7H����jc�(=5T���OVj%"u'T�0��|Q���'v|E��=�k�/`�gJ!�|� �鐋t��>��h�w{0��v�G�5G2�9�����(��*9�\ˊթ�$ߛޥ��6�w��}�ҿ�V4�vf�U#��Ǔל��;��A�}쯐� �e����� G��{����R��=��` � �>�/�?�-��ۻ��<�p������	[�)��2���"�A�!|[�6�2ճ$}}��� �!��9zu�˽�:��0��A�_7X~e�D?-����=�t1��v����%!�.v�3�f��qn� �y���:8�@i�>�2���e�{���H�5rw���-��׹Y���:�V���i�� 6��@�,�����~��<r�̺�]L��=�v;3s�G{	}���p$C�!�b�w�g[+A|G��~2R ���C-
��������:���|=�^�k�^�@3��l_7Y���6�������u����@�wd<��M�n��n�t�#��\O�Z9�V�`�w�e|��@ڻǒK*�fҔs���1V-jv���B�_KՅ�+k.��Spj��t����ڦwν�Z!�o]�r5z`.1�C>U����>Yeh"�n�!\�{����`oul=ŎJ�/f�/����	��6wi��P:�v�-�C*�nU�wV	�r�,]�ل�=�cTk�l7�p��qj6�i�<�4|��=�i��۶Y��s�ټ�(���ʢ��3���-�Z�VW���F:�YD6��A|A�7�_9��Eq$R%����ǩ�;�:����u���e���쿐\��|���6�n���e�Lz���J�n:mbsry�:�\�>����R���` ���PV;��W��������qG�?&�B[�P=�0��0����O�n\���o��h_�@�>(�[��!�?7Y�q��W'���ւ�.Y=�.�-������i|A�A C-W����pE�_�7�f�}�I_Vr��s�+79=+�s&l�f_S��,9��oݸw%�_����]V��Θc��֭�hD�8Jĩ"�J���n�I
ܰ,�\Ʃt5u4%����̩��1��<R6dMm�z�6bYBÖ��7l���X{8v��8��x�࣭V�D����u���P�M��;L�A�Z(��;v*�G����q��m[�,5H1.�R�ve�����1�]��9ym���=���:��u�md��%lK����c�M����OM9�]E%7a`;����ϸ�F���P���D�I��p�7b��в�$�8`��p �����p��-��+���=��x9�I|�}�%j]��Ob�~���Q`� ����Կ��-���l?�f�q:�rJ����,��:�A0��A؂��T-�����>�#ھ_9A A�!|[��С+��B�UܜCe�kM�hgH�lI�@ӷ�|Ch"�}^ܥt<&yn=ƌ��"�AN���{r����V
K��qn �.3�J�ߩ�?/W��r��-���Y����{+���.��t4b��UE��gW� ���؂-��YϿ������׫���`�x�ؼ�j�Bw3�o���P�X.�� ë�����6^���n�M�����q�O�9�q~�~��N�z����y��-WŴ-��,�{{	O�H��.�Z���[�I�rA`ق-�XVz���S�c��%�>���Q3O۴K˫�L�^��=O6ΑY��^���us��
K��qn�A
���Y�v/uG�zW�6�2���i�B�2z�@ֹ�!1��������a]^?q�D�"� A�YD6�+���O^.%tn>�j[� �Ȑ;X�������샋?v׈ZZ���$��8��w �t��(�waM�d0��g_��2f��orュ����@������hu^�C�_��O�>�۷�V��n�Zb�y7^�G���\���ƻI`�:l/!Vx���?��_��s��g��h.�s�{�Q,��������z�����(��A|y����(����z��B0��"D�5��;�9���w�{b~#��4�a�������1���t�� �����,���\�77�K�`��A�{��Q�%]�w>w�2$�!���QTv�D3~�m�>���aP���XĻn�����/3g���1q��kӐu�l�O�y�AD�?7Y� ��e��4����ޠ�#�U�m-�$"��{�J�t���x��3g�Mp�� ߁�_#�Ch An�L�[�z��?=�N�N9�r7Ym��}v����Z����u���y�߿�J����d����逶��mt�lq�;X܄:#%�X1�V����%�w�e�}�ǯ�t���>^St焹��d�w�~���|gk�m=\~�V@me���G㮻A�7��y�6�gU|~����2K���$���<|?kA���]u�mӎ��8��5�,G}���mź@�B����VW�t��������_��>t�?y��e��͠�t���r��>t͞��Πe랝�=�Rbsa��>-@�EON��Q!fF�4�̮�Wwql��9�Ś��,n����â�����u�72�iRy�.b��E86e��S��9���+��{eU���x:D܀e�t� ���^w�^f�Ź� ����b-Ν˫�o�|�׏[�Ϸe�{�Gn��]��5�K�.$�T�%X�)ZU���Rl�*���Wj4����Ysf�i�iM�4�_c,���g����SU<sվ�Φ���p㾡�Vf�T��F�~n�n� �Y@��g,^r�+=a=H�3��n-p��w�'�-@��%�{n�݈��B�A���;ԁ�!��|~mye�v�vG��V�9l��:**���Ǐ� ��t���6�B�z�izٮ�&�{�P㈒�$��;&6�tgp�����o�}����\��H�;u���B7"�;��u��,���u�W�B�<x����=>�xV��N����A���a�НȡSs�i�n��#<1ei�\c���-T0g������6��ƛ���u1t�[�DD7��Z4��V��� ��C����~n��}V"4�"ib��$�є�ZQD,ݴ�i�L��N�/oGĈ8��GY��)w�]���x�*�V9����Ä䎦�
��:��u��WK\��.�a�.;�]F����[�u8cT��:��\�{v�K+���hr�m)-��zv�ό(�zㄗ���� ��mu�n�+���En�� �-s�lȦ��
���]q[��G�ۿ>𶈱Rq�zrƅ��b�[�t�/im�y<�&YF��+�>�ķ��>� C-WŴov����訫�_W�}K�F�8t�5�r��+�H[��.ꏔdX/Ԉ?wH�LV�/;��X�5l#Dq��f>�}��>��%��`��P ��@�H,��n��i�1X�V��-9����K�N��΂"?7XCt/>�fk��:�<���"<b�W���_.ǥɂ��z**��<}�
��}�˹jy}� ���|Ck��t �L��n�A徚H}�a�1!�<پ\^)�nV0��}�$�;d:~��U��;P�������#@��WJ�k�+r�j6�GQ��цShY�uZ�iL\���W�6X�A�K,�?_�~uZ��N������̲ڮ
�tYB�ea�����t��h���S�٪�xuǸ35�-��WQ]kdMܜ��lb�]S��j�ì&+�^�\�Y��˚0b�ʸ1���:s�*N�&�Uw$���������	{�s{��uJ��<~ͯ�k.yY�3�ƛ:Q��t0�鐾-�����u��>��?}��>�7�9��A����|[A|[��VT��h9Xp���Ǻ���L��з���#�λߓ���	!s9���sx�����Z�Z��-�!��^�t��q�r��٧{�S�C��i}^��x��Aւ-��Y^���z ���L���Ew �����晤:�e�3(ci^��ZٵAh�-t���2���Y~�lo�� ����E���M�si�o�s^�:��O�����?6�n���3�ZҾz��Ts���#�:Q��_T~f��/�~��<���?7@��_t��9}¯�X'\��=�X#��l���h|>�件�?kXc�CT�z<�[Ub�Xnl���3�'�!ݰ�FE���w�;$���ެu�svNMh]�C�![x�J��lp�H8S��*�,}(d�n;/$+_XMǽ$;/t�����m̭��������3� �ѫx�bjClq�7 �v��5Ũ	�:��֞��ڄ�m���ܾ����d��"�f�jn�z�f
+�0V�v�kj����Vһ3S����E9��t���Ov�7S*�m���Xq凨�vY�Q��]�]mA}}�ҩ͒U�ɦ�USE�{���:��\�,��]*�fr(����rꉱ��/gn�+���H�V��h��
�t,54DQ�.:b��fo\�g�n�ƨ�A��ϑ{�`p��Z�:���`�c�Y����|K]���Uu�R��]k���U����a��޵�y�_S�����ݬ�;/�C����8Q��|�-\f9�j ����t�U��-��do�A�h��]{�2�u���n�9�	���Q%�c����M^F�iKx�f��7A�A����gA���V]p:4'vz��>#m�+�r�OE�s�w�����-P1��J�����\�zC���Z��[w�RKwn��\I�
ʱg���D5�x�Z���n�s��a�V���}�{HLB�r�u�E��	]���*c��Ӷ�j�<��2��0�ȚS��O6a��m�q�\��%�^Sʔ5g6.VhԊЭ����x,q��N�,LZqK���'�1�������\�����D�/.F3 �F�A�#IEE3&�$�,م����@��a,���Q�E�CT7w`Mwb6� �`ɠ�X-���5PX�A�,Q�d �s�lI����1F��&I�clF��j6A-�$�#FP���� � d�1L�Pc&�0����FLId(5����5���#PE�hܸ�Ab��j,X�F4�������]�� �(�F�Q ���ZB���W���r������s���3�Zx@��ʌ���p)D��XV�ᤂ�L)2�I�
H)�ˁH���2�i!�������/�� �������Z_��
j Sr�l�%$(C2�$��_��\�|�y���?zH/+�0����)��P�M�����gh��{U���R�I�}p5tAH4T=�$���E��$T)�ˁI ��e�I��
@̢�W�9�=��ޣ]$Je:��
@�o���swU�4����$���AHQTr�H:��Z��P) ��g�%$)�4�XW�y��v�����2ϧ8�]�$	�Y�yP<��I`�G!u�n�IW�m��$�j��H)*!L7ʅ�he$
��4�Xi �Yp4]RT3*H.�������/}�>���}�������Y��/��~���W���JH,(?e�I�����i4�$J��+.$��2��� �(�2�H)>�_8Я��^�����G��d��ZAH(i��$=�_��������}����:�^W�ZAI@�0��ɦRA@�ݳI�����e��w����W��a ���- ���7��R5)�e��5RAaFe�I��Re�B�Y)��e�������7��\��l��f�U�}4��~�I�;A��AH(�- �Q
H-��$ЁL3*�%$*!�F�0���e�������^�g7�׼a�ꅲle$
���A`j4�_W.��	~	G�H�B��N�y(^ي���H�- �y��׮!�%'��� |�v�&n�U�,�����q��:Gp�e�gٹ�R���mU��۲q�_u�G-P=�@�i�i�j�ۇ�"�_K�߫m}��6eW�i �s�- �����h�ʅ���P�ZA�D) �3.�
h@��b���9���d!����6:V�~��ͬJ�0 W����~{˄,BouЃot����}�O~���m/�ۚ<�V� J����]����׮�Y��e��W�SsV��7�-6�I�)�*����XW�ᤂ�L)2�I��$JNe@��xw�����5���JH,9�:H)s:���f�QiR�RAh��$�0��2RAB�3(�Aa��\�FH)(B�fT- ��־�/�w��������]n�{TAH5*�$A�����k���{���?}������$P�O}P-$��¦�p�Aa���E�{�v�84l6�Rۨ�R�P|� �*���H:(�$�ˁ���XfT-�FJH(R�i~�l������gv��Vj�j��C�Ϩ<�I ���ɠe$
=�4�XH.e@Ѫ ��H.� fQi��+Y��s���}�W=&���ZRAa]ˆ�)ܢ�hB�%2�ʁh;~��~�j�Ǳ5����H,9څ�����i҈RA\�oN}�@�AO�
aߪ�2RAB��Q���R�A��I%Sʅ�j2�
L�4�XH.e@�{�~�W\��{���꧈)��T-pS����ϑ�j�U�H�	#��)����ZAH,57ˆ�
A@̢�
Ad�e9��9���lA��<�e�6DfTXߣ!_v��	8a���/���̹x1v�U��X�wX�{�+J5B�=(�ʝn�f��s��s6�r�v�{�U!wb���T��K���Ma�\�i����y릒,�
d���í]U��\�E���Y�����S�6���o�������U��t�v��� �hX�V���L��u�մ�q�ru[=���v�0ᗈ3G-��bۺ}���Q��
c�SWn�˒�֐�xm�^��j6H#Z�YL��� �U9j��L� �%���"��r߯��>��:����S�xtj�⛮I�yƌt�q�:��Z%ؘ2?����A�t�R*�ߨ���R���
H)�eB��d����D��'�LV޳	�{sVcT��#�J��y����3�����<�/�B�6�H(o�i ���p>�� �C2����`Re���YL�����II�}���W�������!� ��?r�I�) �S)wہh���u���׏c�����$��� ��H:(�$���H)�
a�P�}�w���s�㝓�AB�ߨ�Aa��Wް�$��0�T- �e�H,F�
�\�
A��eCI�w^�ۈ�؞����ȵ���|��G��I�){�i ���.H,43(���Y4�r��R�RAa�P����7�g����Qi�(�$��j$ЁL3�f���
!�F�O������3﹙��C�������
J��B�42�
w���~u�9~�o�_?k����|i ���}p) �����
@̢�H�R���В�
̸i ��-'>��Ӻ޾�k�����r��R���}*z/��\�w�|	�>�<h��$(������$�}�
H)�
a�P�j2RAB�̣I���}����6�Y��]���:�e�t��`�u�����[\�u�f�=u+[�s�t�Ζ�><�RtB�{�d�) �Wyf�Pi �Yp5tAH5*�'����Q��߼^)vUg�H�	#��YG���W.�&�V�!�%$w.H,40��I�B�%2����R��$�U�E�J!I����u��_�n���~�W_��q�S�<�+ؒU�!�z�y-h��4��/:�U���>.m������y��}U��n��^V�w�d�k��
x@�ꅤ�����$����������3>��u �_\
H)<�0�ɡ��P+ܳI���Ar��j���~�>5�
A��~�P�At0)�(���R����>II�eB�
A@̢�
AH.VO�A uo�=�½Wi�9{>��K$c��Xs�$����iTB�\��$�@��f�JH(P�eH,4��ai&�6~;�����~aߪɌ���G>�I������p5tAH5P̏��&�nb�Sw~�x��U��	 �-<�I��Ok���JH,3�~߹��~�s>�g����Q� s�ZMD) �S)�v�R���XfPi�AHT�2�H:(�$����I4 Sʅ�z��Y�����^�iA��'�_X���9�z�+z�_�H.W��
O!L;ꅲi��P(�,�A`hi �Yp5tAH4G�(�Qyg.��j�� ̪5B|Lk�p[^�
��o�m�[h�[�M�ĩ���C�?�q�N�$Td�+�I ��߮H,43(��B�
Ar��R�[�gr�{~������v�i!�|��{\|����
!I�ך�I ��ϙ) �HfQ���R��0����)�eB�
A@��ϵ�9��������w}?$H/�.�� Ԩ'
#�MV�(n�߼1�b�_�H����YL���p)$��·ۆ�0��-'�s����z����R&2�׮$���P|� �v�H:(�$+.$��2�l�d���fQ��Þ�7n�y�h�2�w��0ED�E�:�9��ߋ��f�S�����;�Z�}<��Gu�S�o%3�&�xQuXd���Y촱+yw��@��_�>C��.�����3���u ���?�H)*!L;ꅤ�����I�����E� �T3*H.��3(�ЁI�߾��ɯWs���U�
H)���\4�R
�E��B�
Ar��RJ�w���M�ٟhֹ�H,9�:H)ݢ��!I�_�]��o>��r$��T-�) �B�4�Xi�$+,4- ��)�eB�5I�,�A`j4�W2�W��o|�ϴ.R��Qh
o�ۺ��k�-]��$�;�Zx@���J^��ZRAa[��I��Re�B�Y(���" <n��]vW�f��j�����3V*�lb7�hs�-��=�]t��g�T܈ކ�ZAa۠�� �*���uD) �]�ZAM Sʅ�L��P�3(�Aa�[����>������~�:�W��<0�AI]�/,���a�T- ��,�A`hi �9p4j�)��eCI�0)2�MD
H)s.��%$~�����׸ZAa�)��i �j2��������uә�Ͽi�:)�;A�I �s�ZA�D) �Y�@���@��e~�w�oNj�$��P�;�i ��
���:J@���&���hv���R�kv���z���۹n8�}��s��X ��Ch!������D�~����LVVjSQ�v��k-�o�|�$�}��gf�'u�<^{�Q;[S1�v�PC�A����n^�j&.ʕ�s����	3LZ�W�:����,d��01�r��2���� ?h:���Yq���v�_[A�~�wx��4a�s�δ�$~���}�C��PD�@�H~m^������'�.*U�v�4��-v�:b�ڀ�Ó�օ�{l��cKeےg���K~�,�b���n��~�s�<6N�ט������|,��ʳ�����:�%�W�6�?�"7}�;��+s�D#���{�HF�5)���j��X�6G {�H#b�w�zҎ�?TA|^R �aeCh"�  ��vmd�f���W\`�C;7��7��7�wWϨx�q��|�Aj��٤z�ߒ�W��D#Ũ��ȑ����w��u��8�,�W�g��S��W�pO�u�,m-�DL��n���Pr�N� �z����l��]��58�6G|{�Ab� �-
�����v�4�U]������i�G�Ѽ�kD�ܭ��G�7ެzQ8�w{�LU⃫Sm<��f�`�ǭ�:PB]ݭ���������}��4W�7:87h2��+zݩa	�nD�$�Y�/i��-6i�JWL��c��s��mNiS�(^���<
[���r`xҞ�<2�s�mr;��tݝ�̡�-�L�u�A�+�� )�������A\c���չC�55��i+�c�2u���'6Z�[iP����`�1㮳e�Ye�%�X�,nJ�[[#5v�Lf#���}9���b�q�m��I.Ҭ�5p;b=���W��-U�F�H���?�?o�E�DYg��M�K	n�\7�,���%wuCW G��Vh^W��ܻ
��Ҿ�����JD��K���\-k5��S�x������L�/ؠ�/׹�<l����� ��B-� ���/Խ�r�z�'u�n�Z�5�o�yĐqH�C-
�����H�6w����y�à�3PGe|�,����ݔ�v���9�wx ~3�!�����Ar�{Є�����2�@��A�ݝ��YW��_�/dH݉+�\/��w)�K>+�G�t���{�e�y9ۣUoˏ���%��ݺ�`���<I������'9�3J�3XCb�|��e��Y�����H��
^V�'g���t�^��<(y��3���V]p�AU���n���Q�*������˕UW�Lʂ��MIï ȯ�,�G��vd6���Lp�XI:�l;Q������N�Dp�+T�=�nS������	`�9��o��ڸ�/,�6�o�y��F�B-����
�<P���",�	}_7Ce�����]����%7�ֳ���ur�q��~ ���݉��t��m!W��]�����5UCH?�B��;�\f�J릩���b�y��v+��On��|G�?-��H�Ye|Amu����l�b�[�a��J�������ّb���y���dH;��m��f�of�|h���(���j�8]�7Y�t4ћ������2�8+���$�<���dO���( e�����\��5ڼ3�}x����<֯F �_7XA�~o��@�x�w��O��")�g6��MSM�����~<�H?�D2��U]z��=��α}�Y��6���_ Yg��F?_B�m���z�lo�]�[��X�,Vsm�n<n��qj���W��E4�+k�1ܣ7oov�:��r;4e�;FZ��������
�c�p̱o��$�(F�B�D�AhPT�^%%P��n����#O�h+\���v�sh�>Z�� ��r��+La�:��J'��<P!��-�D�2-�D��\��P��ԉ���\��ꭶ�Zmo���@��h"k���y�V�āHmd/[����q�zX[n�kkTj�OR�u�\oKR���눻7�ݗ��n��T�pw�-��H�ވ��H��k&�V�t�n�!���@-�#W�NP��#q�>���#B�=�]F�F��v¸�Z���~<|~^h [��t5|���ٱ������{E�7[Kw��Am*x3w5�Z�Z��y�Z����s��W���@�Y�6�n���f=�r��<_�b��b�'N�O1R�Y­ط�|$��+���Wg�f�_T�Mb�{����J�1C^@�����z躩-5Yw,�P���L�N�힋 ��&/v����13Íor�^�6>�I��<?eL�?D۴�{�Fov$�_�����.|�s�wmD��2[���Y�?�nŐAӤp��qx�ϭ�����H�Sj�	I�2��&��̩�����]P��H�6���j���_�������݁=7��4�De6��h3dF��{.��^�WۑG����H�Ye'���4�/0�Α���z�0��]'�	�~ ��"A݌�;v�و�+�h"<|��|�Ak����ʜ�oҤf�C�[~��oJC�V�9]q�;�?G{�A۶�{���ϩ�U�Q�Up�C�/���!�Y�L:�ђ�k
�@ ��r���&��Һp"!�+����ψ?YD��ݎ���W����z�C�w4�[�����Z;��w��"ovP~j�9��h{�1�_c�wg2�
�G|�����J��%��%Tu{�S�J�p��l��b��=�W<y�(k�ڻ�HYV��Ј��/k^��a
�L�t�N�j
�{+ub���I��}���+�eNצD���ݥ���gT�m�ܝݮT3K�r��j��۪��n���w&��LUTA���7��}Wݫ�J��MmfӚ��:�UP��U�r���xF쀣}��d
�v�t�Lj����h���(��l@�ʘp1�0��W��`﵇��HH2��?Y�to��f��jn�9�JP�Nb.��J��R3�D����κ�/9��GN��Xx�w*�г��8�r�lڳ}Mw4i\���w*��U�Ә���=J{#�٢��rO_�9孖���<.�ܶ�ݱ��U;��n����a�����UPtT�3aV�G�{w�����-���yZ�V^gϱD�8�ެ�o(:j�0���$�wX_l�v�ap�\m��UCF�\E���$��!H���k��7;����sk� �z��)�����V�tQ��/����W(�8���\��2ڭWL_*ܮȩsޥb�#�h΍^@����r�S�*��W3W�+[w|�1B��ѱ�b����}ۙ �;yx�fUcF������D�Lxr�䷆`��הO*H�X.�!��eX8μle��˯A�B!�wZ�+��R#;Jy�2�O
�Oe�=sWU��vc̬���N��ϻTDwyvZ٘��5[��Î��Rv%;o�˙voCtM<͡}jS2e��j�+0W��=���>+�D�+�ѱh��J1�jKJ��b4`���E`��&d,A�D���LbŌd�2��$Q��Z4F��6��4$j6���,QI�PI	Ơ���F�J65�`�d�����6��d�.�sQ�r�C"� ƌ��� ر���u��L4N�I�����wk��Y(ō�
�EF
}�ڮi-��Juj:��&�(Xkq)qYs],*�g�gpZb�ų!�y
\c��\H�7k�l-K�;��Lsi㥷g7��p��l#6�ڬ�Y�q��a|Sѹ%����F�>XxK��pV͡R
�)w�f�T�L�R� MtJ]T!VǰE����4^$k����f��6��b���D���<�/3/���s��`�9;qO%����<=�{v;9.zy�6��XW��]����Xw�j�wG͞�ƻ۲q��Wh��l��`��W�]�i2h��e�Hѐ�R��v��3E��pKl����al%-e�2�\�1�x�0�LN,����)��LV�8��M�ڭ�L�T�rh]�	�:����4ׯc�F�tVƭ���bph1������'jͮ�i�Մ$�Nц��a1�C�b8��y�ݶ�J�1�CM ��݈�1��uԷ<�[�ٍZ��K��sr&1ۧq�\p�x�:2.�9[�ɭhd� ���X/k��r['8_5öc�=��n�F�u�]��y㛪��Ӵ�ҺlBU�Y$4mݣu��-E�C.���v��u�b��Kvy =f/J͢�9���y�R9Jk���U��%+�[���l�
��6�!bز�[��]��׮M��n�����Tm���3.r��$#,��IVbW�n��k4tۗɊ�]�9����C��xX�.�*�;�n�Q{Z��;-ΉpV0�n�ŔҰ�l4z]��&z�t0�.uf���aF<��f�s�0�YA��W���A·2����۠�{�Xx�^���[{k�+�IxS�P�1C�"J6�:nBS:#�w&�uH�/gX�cwZ�9u��6���#���.���x듬��p��<����v�A8,�l�9�,<�.�sd��ʳi����i筲en��c'�]��٬��k
�ب���#yؓ1̴�H�^��D�`HW���,3�T)ikS'aeP�1��\��3m��;�I!3��K�1k�g�<u�Rͩ<fn��^Q�z3�
��S��7�����ں^+a�v�%�7I�yyٺ}v�۠�j���Ƴ!ĥ2���5�&�s�b���`��E�1���n%ԁ��oi9�C�ݒ8�]	@�Fba�����I�]�����
�.��� }>�⛛�q���vr���^�;Rs�`s�` �g�<=��Xl�߯����l�8���OS�4�	v�"��v6L轱6��)cw4���j��/۫G�Yi�ձ��
�<�>}���9���^WѺ{(<͸s�@u��W��� � ~-�C�)��SXf1����}/d(��l�&r�Mi���?�D@���&���mR���{�Lt��_t� �C��Ǫo%����tt,]f�'��z� ���|[�������;6�ں�m�n�cA7�����!�q}�̗�.u��@�*Ռ̼p�z6�@|���@��"�e��-խ�7�S�}c���,j�/��n[VP�~=Ծ �A|C-|+���������������K��u$1k�!m�V�F�!��v�n�]e���l�f��-O��'��>��;����J����c�4�[�>�D.�7+ڔ��{z��o��u�����-�?VF;�U�挼��óN�ɾ���f�|sn��En/�p�u��|"�x�Lɦ�:�}��������f�]��:��̽Kd��[�a�8�*��8�����P��:g��R*�!��w�\�J._W����"��U������]H��ޠ-�@�͠�a^b(MF���U��:��[r���u�A��A���K��/�u���ۏt-�*�~ �r$�H$nĆv"p!����'��z����D>H��Y���U��D7@2��b1f���5�ZC5�_2̴��\p �Y�?~�"N�@�Ygǒ��}��gV���RV�7hƭ�,v�c:���e�8�S�ݕ,��k��:��u�)p���:�!�|A���䝾�|n)�M�A�"n^�á5�2"��"����H�Yg��g9"�9�3
yD�J,�	u��v>��A�	��ށ F�'v((�m����ƪ�̲�O.T�j�f�e�ۻ*�_F���*>��������lv{U����ǧ�;���3j������r�au���f�K��mdra.�'Yt����V]��Ẇ-lT�A�����K��W�6���Uj��̵�� gϏ(�۲$*ԕ��c��i7Ek�Z�!��<�i�E�U�z�:h��+�F�}���]e�Z����f�{b'=��R�<!>�~�� ����β���]lf�^��琿K��FFm�r�Y����7��c4��+���獖_�!h���)�IX��}�%�����1�=��|Ch/�/�ͅv~�9tڵҼEtV5Kvs?t��RYg�� An����4��������������=��d[�9(8߅}VA��D1�4�F�¨g����T+�?(�	)�J�&w�趇���	O���.=�ur>�^?I�P��Y!�SZ���Nh��d�#��%B�*�V#=|r�T�Q��Op�4�\s��U4X�i�^�ߵ���Uj�=x�����]L�F펭�\z�Opbr��xh���jT}f����/� �� ����E��fgƅ̢�r�/⒕����ODԔ�� pR���c��}'%�}VA����_%�v�x}��bm�Z4v�V(�tn�ʩZ8��s�kAc��ըuv�6&�љ��M&�W�����_w���U�Q�
(��۱1��}FxC��Pm�������"�$�4"D�@�"�G�v��,^m1]����r~���y[��#}�r�T�Q�� ����-����"X_Y������}( A��E�dB��{�RӵչՈ1��Zq(3] ��O�� �R�������(��0�m�P��b~Sޱ_�$�E�;NG�a���p<�H#:#����`f��E���� D0��YH�?Ir�ue�^ݫ��+����
�pe�ܩ�����$�IZ �*�ë�/>�����i�����Y�ˡ��"�7�mS�ْ�6h�+u���Y�攠ˎ��n�N�Z�S]ϻj�m�sڸC�ګ/i^N��������u��v֢M	�X�`���r�e��eoO��s�����#��9�)�XMx�ۜ�����4���ǰn��zG��lG�:ηlQ\��#gN�ָ�ڣ�q����,P
�k6�l���ť�-�7�����e#=]��MHc.�rD�]�;������6�IݎOX)77g��k�y�x� L
s�X�������U���#��޹�����Ye� jBݶ�m��.�]h�_�K/��?���S��H�mW>�c���i�/�G�YRzu�>s�mO�u�����J_~"JDe�Q��;F����<yD�	B�]	s�1�t�e��J���F[��A*�� �r���|$��Iam���Y�Y��y����=��W�$w��膃%"��K����Ό��O;OT;�9����D�'����-��6�[6�u���U}� w^������|��,)"J_RT+�vP��_�w� �����Na���/H-�y@�A���%8A�D������}�58i+�Jݢǈ�8WN�fT[&�lD�Sv��a�qǌ�S�^�@��EC�?H��Ib�m�扗��œ�q��A�Q��}�����`"Ib���A G��x�����g6w9��ʗ\�n��młL=�	�j�ŧ�Q��V�m����n
�k}k�h�,-����xu�j��qT���}� c�ܦ��H����1��mn�q}���8��u��AU����^����A���'R"8��d��U*��=�Rb/��%��.C���<�H?o�/��}r ��Pr��ϳb�AP@���Xͷz�{��٪�J� �ޤD�b����a�w�OW��%�`�d�� �*��*mŊ��«T�͑7-k�����ku��3\ $V>���b����3UfyK��[m�@�9�4�������7Qv��{5v���JGZ�i.���"=z�"}�ѡ̫���#51b]^�<�,�羡�,ʸ*^�6z<t,�6����"�a�IM|B��ڝ0Ӏ�e��6�^+Q��b�8�dĵA,��ZT(�w����$�C
(����,�PJ�H%4!)�te��1�wj��&�f}Ԗ!)��BTG]����̫Ui����ѥ�c��_y�T�1p#�݌�:B��N�V�$��Umm�`��  |'��vv��f�uh������ !��K�J߈[ۆz�^��4�`�s�@��QG�B^};Ã�vs�W�@�'	GGƬ��-�y�*�H�dA!�1�ٵ4������ՁF�p)�ɉj8���D7�%"	�į�&ģ�5h�	�T���A�]h����se�eV�W]Z�\��+G�!��A|D0��+"�O��{��Π�\�.����]?5C��B�"IIZ&W�6'eUL��w7y�<�A���%1w�Mp�m�9��$v8�%=�l>x����o�@�0�~VA�ϫ��ǯ+��Tw-t�t�Wev�\�CǓ�}�x�rU�Q�J(�	*��2,����Q��"A}�@~JC�}ݝkKDef�uk�q)�F:Ws��7룦o�y�AZ�K�UmC�Jzα�i�_a���T��W7��\��.�#]���:�^f$uÑX�;uҾ}�S������I ��9⣜��eZ!�"Ib̔��.�ߊYg�����7��Q�m���$v8�))��˳��{T�`���P����$.�dL�&�2U����*Q#���������7F75A�w�	iM9���JFZ[����t1�ĵ�"��f���6l��"���?C
"IX �A|G���b�j��Gb�!�j~�7�ON>w�oz�M�A���S@�p$|B*�.V?(�B���o��*�J E�E�P����kq����9�	�!�;���:����YD"�<9���|���S??��O�i����U�X�`Q�ڮ�[��W�>(������+�Z'�]"Ş?I4X&J~��E�o9<�ԬM@�����S�
F�iƠ�tRJ���!�W�D)M6�8�ڪ��<�� �z��ѵF�df[iDºrP�R��!��
�N�1�.�͛ǚ|*t[{�(�*wԯd���nKõw������I ���ݩwwf��j��b���Dꝳ�٭u�r�.�V����t�є���˘��X�,q3�'ۣn;<�6lt���q,8ֲ�g�痻Ԝ��j��&��,��]ٰ lMq��e�P�z����׋������v�� D�p�7M���;Dt��nOK�3^	v�gDz��HnǺ���Pܷ%͍�����K�h��9�M����e��������,�@M"�n�pi�����m��W��W9O����8W����fJDa�I�+��7��\-9��f���$�dH/�X�A|D1P?"�F�9�{|Fe� ��r�_Z���ݪ�;0�w��x�?J��M���⌅08o���y�uD0�$ZA!��x�s�_�C����r0��mƠ�tRS_G9�+�"�J�=�����m
8Q9ز�I�d$�������+��P��K�����UZ�|E�⿈�� D1
����~��#7�nKg>��]
������(���Q�|Y�$�
(�A(���2��5@��Q�M4^ȧ�i�ҹ�nh�4ȵ��\m-a,+���ѥT����"�^!$VD���s���T8�m���9W�ȭ���`����W�D/�% A0�8_�Z==^��oCv!}Lf��n���T�J�w�8v��^��o�"�7�Ni��{}���5<�oZ����֕x�u��8�w�>��MZ>ؒ	E��Q�Ur�ߑ��P�hxt:���ι�����F�����"�b�IH/���KN���U�ܗ�EV�y��G�[�f�eO��6���ѽ9Xs6���y�f�аA����}��K�|���Y'juk�Қ=��w�pw�.:�ivc���Q��QFH)*R��T���,ᑙ�p��m/�Nt���3��Џ7AsuԱ�e�Ds,��>�~�����uQױ'���E���!��,���Z.�����^�&���OW��ΖY��?I_I��;�^-��Zޭ����Y��*D0/��"��X3Ԉ?% D�2P@�巏N��ߍ�VAjD�nv�9ܶM�����H?jhWH��M�тr;����Yt(� �F�|�_IP$��L�X�Y�����;F���5�B:�Y�Y��I3q�r���j�J-�ewG8�U5<c6W���%\���;��r�����9[W.�GJm<
i������T��TX�$A��Y��s��XU�V�M�(T��ڠ��?��|���wc9��w��mq�{O6�-��������w.�k_#��K���.��;�T�^��Z=9�w7���G��7�g	��y@�͵�3��$,';�w`;+�:��S��ז9����0�[��fx�7T�*�3y},��9���T�������}�к���l5�:����'kq[f�4��<���^.���0aA߰ᩢݭ�v�����6ƹ��FN�ʍ���i֣�!�Df�7�j�ӂp|��{��sS���[�S:}�[�)�\2�vA[)�������̧Y���5�b���wͼD��C�����,�w�P�p��zx�	LUUJ����0^�k�U�7k[���h_v;6.K�T��(ھE77���{�D�Y�Z����Zq0��ۂ�J�2�Y�k����:�vi��R|����3;793Or�,�YX����]���cѽ�m�JXf��+�/ntME�P/*���պR%ӥb �1x�vQed��vr�����6���׺)�q��9xF9*���J��^��w1-��&��^lh��Yɽ�(r��ª�S��w��F��T��mܘF�{�Q�W!՗��ۭ�N���/v�f,+m�����m@�ST�t��c��Α-��B�6�Q����E���Q�n�g)Q��o� O�|ݺd�W9�WwZr�-�j�JH�4bM&�Q�F�h�Bd�S4&�E�YDbɨ�ر�(�-b���1�j��h�4m�mLՌ6MA�Ũ�#IRTd���m���Bh��)1�ccA)"��QDQ�:4h1˚4QX�h�܍���&X5c(,T��F��h��� ��汌�M%TbzBB}�ݯ�z���Vt�yTs���~�]��s2�e̻>1+��!䣯�SW�h#�r|D��㽒��|��Z����OR!؛5�Wox��+��;ʸ&fY��Qq2�����69�X9����|�\K�%��]�/�O ��D�Ibe����o���}cǣ�gk�CHE��@�fm�ՠ7	Y���������,�~�2���=���Jފ'Wi�}uS���ւ�#�ɪ���A+ ��L@�$W��0y�^����|vu�k$���_�9S�8D��B�Q��kz��j�r ���	��H))��==M��꓎�o������>����X �<��+�$�/�%}n��₲���T����_ǥ"�II�_)Wn�^���5��s�H"E73e�7q�^I|F�3���b�b������E�o68��9]8�8�BM>7؅��3�np�n;Q4XV�t*�ň�����k�$!5[����^�3���3,��f/�D�Bh�ә�>Rm�/d����9�۷���ԁ9,Y��$���&'`�:w����:h�M
��1PloX댐Wh����m(&m��.K�ћ:";f�����_v��A(�%9� ������p��mugsr����:w޸��{� �A|ϐ_%�%}��"+nT�D]��D5ħ-ʉWKk�!p�q:��:�A � ��鼍=x��Vq�#��?��>VA�H�?H��I,P��8��N�4/����V��#�H ��W�(�HJ$��
�����q�۱�����!�c���ӋouV���jk�m�n`�\0���?�W�F A9_!$�`�LgB�7�`VTu�'t������:�N�	%?)Aھ�ܬlkޫ�+�=�]�2ƗG{u*�M����[g[[�W��r��#P�,r�|��sz�s|mRF���ɀi��_ו�����j��%�K���g6�p]�vZ�rI�Ͱb��J�|,d��`T� ��8�ja�a���A�뜰�[q\v���m�eL����`���L�û�=q��&�8������9���V�f��h���c�N#7L�l��D�M��WF�ܦ�ܼ칺��l�&�j�o"�W��Ʋ���fK�d#��
�Cp^�u�:;0ͧv�:߾��X@��V-�J��s-�3��MHg�'�|�ZNp9tT�c�����̷�ߎ�,�����D��%�wr^c:��紟W��w�-ƦV��6�}Z@��"Ib�(e�"$�^���`�����gk��zg^N��vx ~=�Y��C���f��@���E��������3)�T����uLf���H�t	 �_P@��"E�>s�}~��V���<�??%�X�x\x�_��������DYXl�-�㯗�I_I0P?�I�|��ꖱ��/�v������m�W�uN��t�jh~]!����ǐ��s�IoS�`�h��:�j�	X�+6F5���i�E�k8�;ή���V�$�R�U ����b�2R IS�9N��]+ޣ+��	�P��o(ϱf��~��?��@��R$��?��/�A�L��Vy��>+4�fH��n�I1̝�j�Y��	ă#+VI�&�Xa�IW����p���4Kg{oJ��s{,��of�+*�����}=���5/�ޝb�<.<~���}^ ��>���E(�冄��Y�b�s�#ذK�?(#$VAD"o	�R��#�zڷY��F��t�[S���G�Ib����o���v$~�����A��$7K�)���cγO��T"��	!�WS��q{��4 7"O�H�L�X �"��r�?u�7�;C��M��[��#c�O���>(d�/�%|�0�s�-����G��^�ݡd+j��wV���eH2{����vV붖&l���3!/����~ �D��� ���}w�k�������8D���|/R{}9U?p}"@!�~RK��_aDd���N7e[�@~�ܧ\f�.?s�g*���x�$O,Չ�g����_Ū��d"!��?	%�~�&�`�J����v�6��p�����;Yu�ҭu/��w]�����ç�n��	��0��H͵��f�׮��RvK�� >�Pz�9���L-���� A0��
J� R� �Q�IU
ʻ�v)��P��$�4J��������c�r�w�P �F�^�2�.�=K'�T�{f��U��������^����.���e}1k�g1d|Oi�T'_���A���+ �F�5�mv�ߟ�I�Wj��62��vR-�-(���BSםu���Q���*]��͔�%����E��U�X�c�0K���������J�|��^m���R?C
"H��(	[;��t�˛#>+�~nv�g��+y{�Tj��-���t���Q����
o��B�.R �x���Ib̕�0��2t�z��ҫͬF�m���0��A�H#a�%%5�% #k��|�6��ݴ�+�"ŵ2�O|<%L{I�}��#�Aw)k]�뎤�w�EtM�����2��n��:-�/goj�7��>���i�D��Ɍ��E6嬫4�x��\���ՌǍ��˙�}2�.9�u�~:\�zD�
�3��{�^���9�>m+'�_?)%��yb��8*[�U�o�u���]��&Ŧ�=��X&;WXb{��q)zѭj��Suu��#=m�f�G2��Q��[�����-�.���;��R>���]��鐏��� �@
"AIM0^i[��i�0�}=�-�k%AY<<%K�I�x�>?/����g5����*��&����yT\A��H��A!{ȯ{���r���|������U�3� �jhWH�L�353+蟫��U��OY���#�բ(�=��-����1oapF�#��A����T��}5X � ����YPDC(��H�?��6Vv��-K�Z�P�[�Uw�����G��5*�J$	E��㽛�O-{+��'x��=����lV4L�7����[���7�Sͭy��
":v�g����H�)�����M�;O��}�ߝ��.�m��v#v��ӢYLj�jd�f'v�W�+��]�3u��u(�a+���=�{t)l0��
y���f���=�D�qt�31��hd�B��a��K�q�����N�֊ړ�8�ie�`�L�4@�ܑ&�t:�L�����*���6��)MKu��Ζ6���-;��c���9,��r�fn:�\�������iF��u/.�4�=r�7n���)k��4��l��7X�,���YW�~�<<�&8�̽Df);{3��{��M��V�9�-��3}֋�ZAƂwR������%��K��u��殞��dI�C�n���Ȯ[����WؠH �Rb���{\��.~�	�Ո�w��G2�Lʸ~?$�A��a�󈎛��ØJ����S�v���s*��,L��h��T֎��+hh ����+��(!���i��{r[Y����SS@���*2�(������q:�((�BJE������W���9r��8dg5�}DI�x레?8�@��$B��������A={�%'����FǶ%-�^ϲ�$��������Z�Bk	,f�i���e���ǷE�(��IP�����J�xgqJ��ָ�DO���ei(���=���ذ\�A)@�R(� -�6�̬
�o2�.�)8Q�4�;���S![{�BjL�	�C���8�Z��D��'���t:ۡ��⎞�o�<Bw��P�| �߽�IO�>nD��fv�7�����Wh<����t�!(�T��U}��У}K���	%�2Rd�x���s��i��{�����6�F�� d��P@�)-G�#���%��h/�����$��e;�u\7�d��5� ��g�n�w0�݀9��$�`�%"E�H�M^�ad�!��%A9��׽3�N��:�/���"J@�d�%qų��Y�_�;������Z쓕�Ǜ�����O;Z���R6�
�!"
��~yA C�!)~)@�r����[��)�	���C6n�b�oP���}�� �"�+�d���k��_cYW�r���ʅ}z26�TGބ��Mk� ���T(��D�s���A��,҂ �"�"�D�5֔J��9�V�S(���&�1��Q�z�J��v���9A����;�vQ���r�=���f��	
��ee�n�PB����&������*r�!<x��w �V��@�BQ'⒡`�_f�_/͏�@l��/�?(!�Ӟ���Bޗ�NHM��s`I��cУ#9�O��� r�$%�� ��� ��2!��}4�P�2㮎��^�}_x�P@�q}%o�4<w�x��=�2mY*Մ	��D�	����۲��]��\�+Oan�r,ʨ�dB{_zY}{ �D���IH�O��F�r�����g�^�e���ڬ[���g���I+��(�$]��<n"R�yy�f�|A��n��e�m.��[$&��9��q�~�Q˟W<8-j!�RS_�	!1�IP���8n�>��G&���ԫ/k�����P�R�����,xS�zן���A��<�~��4�#�j�+�J{�)l�;�h�T��q��(�������Y��h��ve�jF�}�G�t+�{3�Tͥ��m�Ҟ�Z��C��!	��C��v)�'2썻�fx{���ϺE�L0�$�X2S�W�=�GJ]�{*�)�K�<�ɀۑ��~�JJk�$�str}=Ǎ;����46��t�����v��u*�C��79�F�А�m�[�r�J=�*�u�X �A�K�$�/����</{R��9�;�-H+�Yw1B�(�ӯ�����A	*�JP�ؼb�N>�s��܉�dc:��R���_S� ����A�A�:�����{җ�6u�%h 9HD�Ń% @��o��l���Uy��V��n��}_f���P$��� Ȃ?H�S��^φ�y�@A�?oO��	*3E��n���$�/돸��!���ٙ�4�� ��D�JA��H�y�c�[J��M��n���;��*���3��O�����E`����%s�	*�]R`�7qy���DY���7[Ğ�#��cӫx���W�THȵy�ͣB�vm�YX�Ȱwnp����2���baB����hekx�j�hoVe� �}O�N�[�n�;���(i[]����l!�v�U�Ix+�lC*���բ���v�s�l<���fQʒ��5OGI�֮�[ka`��(�gl,�jb��'����-����:��V�?\���b�iD�v��E-6]��*j���K�:E����&�Qb�c���.+*�g@f���+�v������M]�h�y�T��le�Ә�k`�ٻ��l����ZW�>��KgE�]��LѴ�������(�Y�VlCmظۈ��WQ�o9�a{φ*RiQ�e����KZ8��.�vٜ����%-[���BYݼ�+wl.��1J���b�G�.xN�a�gOi惫���aރA9�%��Ƕ-v����豑Eu��yՅ���-Wv|���]��4�CQ���C.�ܝ�4Y���S�(��Tt���f��6�oU��AWesF��+,Y���e�r�k�����[��uu{�M[=��+hj�[���ݳ]�R�Ȫ\��U�ʫ��15�h;]��C�Iث�����0�����i�����t�%Q,���k߆�y�ԻD�+tc�k����F����k�Utї����WWi�"��j*���t�P��7����b*,=Uo�fU\D<_Cb��1_K+�̒�jC�fY,V��uS��0޸�Iwz�f�!�F�@��Nӌ�յi�"j�ٜ38��?|Tlm%��LF�U�])#h�4ccr܈�1E�d�J��lRn���-F��j�×6�sb���.�ͮAIh�$����Im��usr�d�1Fب�lk��ܶ��EQ��͹n�6�m���F���*��Dh�)5b��Ѣ��t
KX�E�mrQ��9�SH�b4T�(�F�رDcb4j-�Z�QT
d�
J��A��}�WV�U�+��p1v�X0�-٬J�����$]O��Y,����pr&�v��[�ņe��\l
�]l3v[���!�u�.ch�oh.��6�8�$���Îqے-u1�=k�l�ѭ�z�O��ݼu���/�q��,N4�����&n��1����1s=�����N�Ԙ����	��ܱ�ZΪA͐�a��V�R[���;=���SF�F��i���Y�Ė��c�儌��Wj��mD���P�,#�ݞ��tYF3kf+�(J�P-�m�0����mډl.�cK���G�v#8x�!����ظ��x��-��&[j&}�;v3�F[	�4�sP���������i����re��-���+u�.V%�%�������ڠ\��V^�����`	��2ӉIt���]�#u��ׇ�#�d�6���	Gg�jy޼�rY4�t�;=¤�^���[3��AΜ=�ӹ5ok����;�ti�q8�wXM�&��T��3v�1��j�%�-�\<�χɱ�١�^wr������VJ��n�)y=��p�s<���Ug����Gv�6�T�踶6�{]����:��gcGc�' �[t���ذ7��v�g�*hS6g���q��s�Q��v����#%�E��9�e��n.�=q�u5���p�X2]���T�:�[�q�c�M("�A���ë�$ku]>��ks۲�Om��V��:r{k7�Q��Z4��ꋡ4Τή���8۪ok`�yY����k����]��2rz�vU�Z���V�d\<) �M�b��� T�����{b4��&Q�5b�;�x'�8�.��[�F�۳ff����:k����:G�p{��n(��x�mj�%�j���tAkf��cM�n�&�vvn�w]tpx��+,6&%�<�m�R'��bM��;A�of�u�;�{>j����)ts�����z��U%��(m�4I�Q �:YM��m���O/�|SX!��V۷�v�6�t�n{j'=pz���N:�Ju<�g���۞�^�3@F�� w
��y0Ֆ��-��RE85����Kt��;Zv�ِ�m�,nj�"Q�v������!Y�'�N܉{aCp�׶��ֈC,�"����=]�Y�o�l��9iny��"�e��u�sz=��Å���Q���.=7N7��s����~9L>�blqLf7��բrVֻ>�9Y�i��l��A�s6��Y����	�H?n�
)D�P��|�w8�v�$���f�TC�3��^@Dt2y}bE�&H��&�&W����g����
��u�=u=�u%W�o\q�� �3]
)C��8yr�7�+��O>�A� ��	))����f]nK�����p���6U�y/�|'�jh��'��|D�Ń%/��;H�BUo�fj�J>�BQ?.��i�pN/n�O�}���{X糰�PG$V=�/��$	IO�@���"v/����!�hP�����nM��q�xL>?'���d��Û+o^{jߋ��ϴ��(ڱe;�ϬL����pݵu�8P���Tp,6�2qv�J.P�����y�D�B�+�Aox�tj2�nʷ�e�o�E���1�-�s����ȏ�J���(�?cPƱ����ۼ�f��c�Nؘ#qܮ]�i1��u,vF�ݭx�p7�mVu������&Ǩ�� �Yk�vjyؕH���h"�;��2S��8A����D+����z�v�[|(�A�D�"�<+P��ʵ�I�j������ D0����zyKh�ε��vm�����yy4���>!�_I[��
���P�c���˕� Y�,�s@��#\gN�-ft���f� ���Z}V%��)Y�+u@LP"���F�~?"��~IP�R����0iӦ~I��7��Ïd�����{�u�D��! d�� Ȇ���J�����D�`�j��Ϣ6]y���R�mR����� f�f�vn%�gO����K�$�T��)�y�mD?i�Wv���!�A�WJ�]�����+��$�>(� ���(D͌��6�U��#NO+���Ao���LE�w�b�P�7����@�2j���]
���2�fh�ʸ�q�7����e	i�õ�˯�򡇴t@���!����[�7�1�Ŵb��������s�����ѥ�)hrv[8���?V����n����Yv�Nԋn~���k��E��"�b����Y8+my|Ǣ��%�K1�����ۗ�N����Ռ�w
�þgݻ>�r�C�V�!fJ�d��2D���k��̱C�	kl�m�y�����A-��.���%�IaZ$yծ�ol�˷�W��"m�x�,���B-����V٬Y��Ut�3�V�J�o2�h����&g4hs*�BQ c]Х�>%��dmH��\�k�ŎvOP�A�󯷢߈"D3>�A�M�c.��Ă8܈�>�W��v��}g2��a�q�_@�A�
���v�X��Q&���ʠJ�A)�JJ~J�M�F4�\ٶ�����"�8a�{��YyD�I/�+��#f�NU��C���� �R�9˺���YkVB���sc�VWl��&�UA[�nA�mA���S��;Bs�ɳ㢳�(�8���^�V��,�闇Z��K~��S�ّ��\b�?��߁���r�)��YPDIH�?��ne��@Kt+ݽp]x^Vջ9�8��PD9�% A��C��YUWᕶ��>z���k��خi��\�����	�\Q�I�uZv�tHjdB_o���}~#e� $�> ���vt$/m�oa��yC����|󰼭��4�9H�_% �O�����iˉ���8�A����l�uY����A�>_ d�|�Q����W�`!������ �V��Ic=V�6-m#�Y>��O;�����P_�B�2W�� ��������ٝ���@�A���A��A	H��غU������8a�q�h|EdQ"���F�$�C���@ ��P)D�1�s/�p$^�-Ov����H�ްN��ϗ�"�A	H߅�]��t_Vf��'q�b�c��μ���tk�nf�ޤ� l�߳3��gOP��z-�TW77f�WT�0�#��/�e���;�����h�TMZ�0�K��I�ԛL�k��t����KPjZ��@�v��+�#rͣ%�i�y�uy0/�1`�vn�픵�f�XB��h��af��['��Kp���6��m��jt�QN�rq�C�;dۤϞ�8���x�۳ә8�H獰���ˉ�bVm6��l��[B]��T{�Y0+��i^�mtX9�3nm9�:7M���?0?k��:���[����u9caݹz�u1�N����)W��E��"J_��K��n���͗��_W� �6+���ҵz���{����A0K�L�#��z���uG�y:A�����d����1e��+�t� �S��u�}W�K�'2��C��b#�Yy��Ds*�c�|=�:���ٷE��zۃ#l��1ο��_K"�m}���(wo���ۯy}����
��,^�������ï��c׭�����ڻ���Sw�̬�����E������NV�g�f����*�<pŗ�	X���H!��"�ݦ^�uRF����m�Is��1�a�a.$�U��C^�*�`�;���~d3zE�A���.=���z�Kl���;ݹ��.�V7U����g/�D���H���n�ZV�{�N��̘-N6
ر̈��KZ��S�*fA��]9��UB0�<W:71|3G��7o׶�i���c���	�w��5��9���n�����ï��$wD�F�@�u�0T�wD�|��҂�(#$_\�p��v<���_9�U�y�8[��h�	�R�Ib̔�|��g3�.ϼ��}�W�QFF�����s��,��F'¾́ �e�}o5 9ܾ��f
�8��( D1���Wy��!ؠ�o�,����~g��ԨP)D�	E]AoG�?z��߻�\�0ݫSk/;��)����J�%�d]��l5t6��)_'�޾����FY~��IM�	U���r+�ᖙa��#��g�l�O,��1���ʾ2K��?n�c�{o�ZN��}�t�%�g�k����S֣i�WؠH ��~�*��"Cy��� �#N���%D0���:^]�F��1�Y���m�M�XꊅJ�0R�EB�Bv�a=t��e�=����V�S7=�Ͻ����=���,��u��;��9��P��)y�ۥ|��>?/��,�H|A(��K
%#���D �2q9�A�)9Y�ܲa����6Ώ���F6+b�������!fJD%�$�䡃�V}��Y�k�t'M�ǎ^�dl�`�vPD����v����}M=�!H{-�oSJ�ۋ�7�N^E�m]��W0���m-�1��u�KvΞ��<���t������
Z32Ӊu~�[���8�T'��;v�Ive
=�?�FHIP�~2PC�6��+r��r?���#�3vh��'�3��ܲ\����6�򴾝C~"o�Wxv>L��|��Yݯ�,�IP��Q �QEk����)��=V����}Ӗ�ދ^26r;("uFH�@��*.�F�d^��zo��#A�����,X�cv�W%��UV���A ��_���o7�3n���}W�����h�]��DR�c>�q�7�K���4�"�z����ۚ&���fW��t�%��?�z���D9,�@)P�\�d�#����*�AK��,�*�����s��J�?Rr$�b��
�񷩮�~�CҬ�*�\O�b�^�Mj��u�����@�s�R˥�,�ܪ�#�6'y˙��q����:Mtk�jsoH��S�Q���!�[�$Q��%*S�Ib���/�.:~X��A�������;��r�[�N�qH�޻��.�k������JI�)31�y�
��VOe6���V���^��A����BH��!%R��*�%�{ޏ�H���E��Ƽ���'{�vm�mos��["z��	"�IRG\�$/�3G��|�,9�e��i�s�8��~�R�K�����GH5c%�W�\p���ӡu������i�̚�fD��]c�q{���ǛBs1A��Qp(�y�&�Su{�r*����:�`��ں���Z��"��l1,u�'��r��SOq�Bǝ�1���x.4���[�yiBy�-�i�[��w
Y\9�<��mm�C՝nh0\�b$#��(�%�	���-��]x��)�t��'$��n`s�w��61x�e$��6yø$����g�k��7Y|�c�K�»Sm��Ln$�zn
ܘ�@�N4&�s��{�V4�YrS^&������n��m�֠R�llR��8����::%i�.-k�`��D������ ����]��&���A�����.�V�ڠ1Ʈ��������ԕMUv2��q�������*��Of�y���e}�)%<^۫$:!qν_N���$��V�ӛy<cny�쑒�:Ms�0�j�'���R������κ�A�(<��|�����y��-ᲃ{������T�!')(IE#^ʹ���lZ�e[c:y�7yV�_|5@�u$�(Vd����0�E���34M cXSS�G^�h�
3`�f��RSJN�rm>���������$_I�ŭ;��ھJ����ߚw�ɎK*�{"r��I6@�r(�L���K�;'��'U���u������TMK�@��9��u�k��T�q�@����Z��t�ٙ�ݑG(��c�@�R�y/��e��s����a2�8,S�pY��W�`{�~Ͼ~��H��$��a��w��h]A��9l<�Y��ʵ��j�7R�H����tZx�z�n��K�&pړ�;&��]c��On�72rn���IHJJRR�&t�.�z�e���e�;	���b�Z��P��R�1~}?OG�i_�dpM�)�ۤus��=vy�3Zʹ���+DXF��H_ʌ8��_!%}$Z����[�py�k5���,+wq:v����$�I�Z�,F��"����ŭ;S�o�g+Y{��C�)f��Qq�S��!�%))	?��ɩ̶�VG~�/#��ⷫ���;Y%��˫�Ş�Ώ+x�E-�vk�*����[9��G�[Q��M&����ڷ���{�t�t�nŞ�-w]`���@�Gi�]a
'*�jr�)�ɺ�f�;�$V'�9l%%��Uܘ�X��C��&�T�J����]�]������CЦ�ټ�[Շ>S�g}Ym�eM���&6��7�9���h���S.�UTM�ᷚ)C�s�u��ȕÍ �ܚ�^�KEl)Yuk!ӳ���0���p@)���0f�
��o�`�W�����/���bz\�Yq1n
����l���o�!2@���ͨ�w��Q�z�*�5�ͨ�s�M�ݻ�q�R��Hk;)�6�|4���p���X�d��J�Y�c����3�GM�jgo)Gq_ώ�˂�!�9�=y���Z�7q%�+zF)�Jgo��'&&�����W2�>O�����(-��0)�#*�m�yYΙ��Q�Ƌ9�d��}�q�e-�pʖ���>��3�W�)p�m������������������E8(PX9��*����W#��evԱ�]���J���;V�VΨB�o5X�H��uL�5��*��UD�T2�w#1�D�h�;T�`�R����[�O.���Oi��7C�u�̨��8%�2��%���ǽ�|[���D���CA��:�3��x[Ӫ1����٧�1�	�7G.��.���H{#���_;uf\Q��՛|�9f����?ݚB%S�w�j1�	��wm������љ�n��\��S�sQr���k���#nl�EPks\�&�h�nW6��r+t�M\ۚ�u�EEF��sF�ֹ�,[�n(���Dh��\���u�ms\�Qsnb�-�v��r,]5ʮb�ƹpѹC�W1�XNv�r��n�j��Qs�wr��ձF1�*Ṅ�S������X��GJ�Q�ͮ�Q�mr����;�޼q��w��X���-S�JBQw�y�������a%?f��(ʷ�%��M�}���y��f0�P�"D$�$%��;-V{|�\-7�շ�λY{ޝ���RP�H�>��LʛԊZ��9��]g1��P�Ğn���My�gH���=��(��i�0%u�lkR���nM�\����/Je�p�K�E��}�WGܺRR�����=ڞ�uZp�Hͦ�d]�JW9T�_�>�j���Oe�6�D�`ꁭK�?���S������	�����ڷw7X�>�;T�����h�)'�ڲ�-��H	@7&��|���K҃y��{" � �ym{�~|���5x��h%�"�TE,�U��8��1�w[5U���),���H`�qv��y�V��n$�i��׺�L��M��!�E%|$�H�,�N�S<�����k"�%�TeR�~�9B8��	8��M����5@�B��6Q�,u�B/#Zڸ�I_ 5T���)XL�!Q���c��	�&|$�LZ6OԼ���c�[�xCR�s�*��@IHIHJ^����Ӝ:���ډ]�=�lK����,{{О������t���V/_�y?W��_I��F+�Hj֓�m��+���֍��9Q�$��%IZ+-�I���9}��o�;Rw��gen^>�>��Qf�D#�����R����X����*��U���9���`���W)�rJ�H��X0]�j�JrGP�S���F�i����\F�\����+�W:���]����A�ԅY�Oo�*P�>;uoC�|;ne�����U:)7e�ט�Ƹ��[���� �����Z� �	I��	\�^`$)s�&@2BT�-��N.�ۇ�Pn#�lF�u���c��'v�`��b\�obY�f��e|qۛ8;�j����Pd/6��h�cp�xǱcq�
�ARX3�4�C.�Cs[2���������#Q�� y�k#U5���X6,�tE2��Zi��y��	��������mb���.��4XWB)���%���:��KY:x��y�PJF*O�\���Hʕ���ڪ�9��T4�/��"H��$2瑻n}q���@[�kN�}�Ƿ�[u��O��?%���s��=���Ԁ�|�����3}ֻB�y5���f��g֗_�)IJY�e^d3�<ϓm��%���o*�&��	�y��̏�Û�w��P�3�d��	)	)�%	,�m�gO�+��jG=S�׹.�.��}#9O�@I$�In����&��
�34$��xa�ˮ]u B]�&�#��jd..6�]���m�FC�>Ώ�z�X>J��Χ}�;/3m�k3�󦪖�9���߻��y}$RW�H�!t��f��P�.�j�8���n�T,{����.�TT��JZD �a��Èy��]R�~��*��-ӻ����8=v��K���ǽa�v��>Z����^����Z�k�t>n $�A��s7^Y˷�1)�(IO�$�8�Q��QR.�N�aۧ������	@I$�UK��H��6�(����r����bZ��ְuV������WU����wJP��R��%$�.�[�w99���e��p�2e�������I�sܩ�U�*��k7��~�z��#�v�'����\�l>�����st�[qT�����D�E��$��}n͡����w�n���uvw��֝�RR4��n1�����n>�7����{3wm�ks��R@It��/��m{�H^��	"PJ�2��s��V�.]?�H�[���6��W���1�хӋۈ1�����խɔa�E��I���|�UQ���s����r��l#n��f��vNZv�c� ��nI6J�+[�)����w�+ދ�$B��!�O�Yol�����/Y�ۈ�}�Z��y%�(IO�'���� �7ہC�{ל3�~��I�E����:6��A��/��^�Y�፝�,VR�v��ݭf{Sؕ��%U_ʎ���k�I3S���]�]k�w�������	T�I:W�^u4���OG=�H�ʩ��&z�ռ���O���!!}��VD@�j���Ҁ�/��IG�Ak���E{��Hoͷ}��~��IE%?1SY��č�ϛS�K#U�^Ou�j�}���뿺����=~�Y٫͢�����<����WTp��@�Z�ܨ̗�����c;v���-u���krJ�t�4[s���gRЪ��rWVd�������O�����9�j�ېML��\z�ݼ���O��֕��TuW�Ubw[�Uԫ���
�,�M]��ڀ��B�f��G8א�v���.��wLJ�}�����=�����U�p�F9�λ-n��D�$���uл{���$���R�}WL�d�O8�dj�ד�mڷcj���ܯ��N�~��K}E���LϾ���T�}$��Y�:�5��y���4��	�C��Q�IHI`�r��uH�C/'����5�wS�c]��x�?\j��ⷐ���&����$��"��Fo�TG�9��M�r���ƶ�m�;�����"H��$�uy���殕��⣮��)��o6�/��U�2�ع&k��VB�Us;�1�c+��r�m��0z-�����͏L��um�ER�)�?S��DeSa��cp�j�.o�%�j1��!����h�j����˯[|0=U�9��B&�=kK�u�ŭ�ͤ`B�ĕ�iVVlVz�����Wnh���	5���]��Ir�� �jR����˂	l"��^f��޸g�xxʊ��t�������/N�1�nF�1�mn���Ǯۙ�;����((�U��籬Wz�[/�N��JP��.�0`���6�J�����B��i�Ņ�q��w��������>|��E��X�윿^g^JM>��@�Vb5�*!���r����	"���Y��&)r��it��PsY��lL.͋��﫚����#�M��y�����)(�6)�;�.��ݸ�|�m��4�=�T����V#OUlb�|�b�Gv=�%?��\\ĺz��,����'Ψ�����h|�����R��<E�2.�dȑ�Or���]0��}\�o@IJJ��= ͺ���}@���UF������s:kSqw)F��v��FƮ�Wb�Y��_�f�'�	(I��{+}���xm�f�;ّ3�8���IJP�����N֑�C��z��X$P^)�V�(V޶}�����8z���7��!|.m���̎'Md�(���*v��U��v3k{���-��x��"胬���'�w��dN־O���LQ��,��~�ڟ�� $�䔥���\
§���6Jx�ݖ�{�\�y%i)Jxv��\M��7sz�R1R����-���Z��l��C������|��S�P���1���Ҍ��6.*�]�WN�D�k��Ok��}$�����W�ZgQV�6��M��
���b�m(q�;��C*��$�`�L>���k����ku>+D��췻�E`�+/z*��5i)J>IL�Y�&&8l>ElWr��%?f��=��n���.����$�2N� T��|2��'����I3�'��o%�6��*v4�9�w��B���+hA�c�FUb�1�rűfAQ��y������6��$�i�bpM����UM�y�{�\���ӺQ;:���~�r�|����"��\����r��V%Úԟ�u�W���r�7Q���@/�脔$�	"�����m^�˕�L����}v�x���	"� $��Oxɛ��D�ٺ�����Q���lLj!0���݈M����J�Uɞ�m��t�����I,�7Dgk}T�ѝ�}�9Vn���^V4����R�s�,^�'���>[�>��R|V#ۊ\�7�¹�ބ����o��u�t�#䔥	.7w�'��i�禺�gx��|�$RE��H<��E�����d=�����3�}7WՐ��x};�,���]̵��,=��u]��e`ɧJ��dZ
��0�>1EVDC�P[�c4���
�I�%��K}v;[�����t�|�w$��������	+�"�Ud�5j�Ɂb�5�Tly�\�����r~�"�I/S���<�����-~�Ե�:���a���S,�Sgv�bąVԻj�Bm�G:��K��O~����קϑ�JFm,��;_,�u������0����}MKi+	)%S��ŵ>V���8��wO,����O�'y�����^]�ܥbz��I�)nXau@�B/9�M!���C{��[��$�$BJ��9w�a�z1�(I��d>9��֗��O�݁U�	�r���u{����g�E����<D�Ɵ؏i�5h�m�];�kb���`	G�'��p���v�2�cfU���'./�<zJoH��j����0fv?,*o�^���5>��J�v�w��"�7v��Z1���a����Afn�)ּ��qN��!$�xlU��:BT+6�}��2�p�y�E�6(Y׽�ѝZv�`T���3���U���j��/S/���	fU\Ь�x֝m^5�|��ܱ���RoA�����`;Hc�i��ؤ�㚹�-Ֆ*�L��v	�u��!�mɑ�W�_����Or2�'תR{v��:f�^��{V�Uk��*�ur&�ks�Q��ثn��]W�'V
�g[�����̳¹�ݬꝙ���fu���h��w�39>�Dr)Ȳ�M�ܻb�G���3��ر\�,��Sj�ō�o-qT�e����X]!�����̍�_M�Ր����Mͧ�0l��؈Q��K�"�\�J&a����7wk#4 ]��E����;Wxb��O{��)s��n�t�p��G���u�i���x�M��0�M��qY	�����e�e*q[���k%���-F�F�o^V�m(�M,�Ϸ6��U-�z�,�y�����aĮ�|�9�m�8�v�f�X������YћX�n��e�!u����"no3c��q�:���+�;�i�Ѝ���Uj��c���נ�]z���#>Km����YR�k��\[�q2ާ�1�1-��l����N��C(՚҅��]�:�F�N�f�hK
�q�����N�t:V'��`��\ud�k^当t����\�D,�paV<U��ɹ��l�֌�{y|��c��K������5u��4�Z�i�3+ci;oE0E6$���U��z��u��A�(��Il,����T����sb���]�ʣE�#m��ck����(���Z�n�"�E��cF�w����r�sc\�9]5͹�����!�6wnr�h��r��sE���nb���1I�h�sk�m��;��1DV**��5���wr�I����wt��X5�5,mN�Z�Еr��ܴich�A�!Q�tM����nW
ر�&ƹ����hHoc�����q!�ѻQ�4��T�xb=���=�|�l6
;g�+��@���פ����z�������rA�^)�4�k���Q�X8k�ml��D��O���ˤ��*��B��c�%�`�}��2���1�:8uL)i[5��E��AW��:�������`dy�=fgݷnfz��}�u�Rh3�oR��d���T�\݂�y�$����Lvݨpn6�چ�+p�m�.�kk�D�"1#���k���lu ���)�s-�m����GC����<B�.��/&�=pV��ݎ��ێ�d_U�Y.�v&�e�m�&Y�%a�v��㹝��3��Y�rI�l�-�m�k/p61�ݰ�6�k�k�����2�5&��Αj�ꫣ�DbS�3��FY�u�w&ls�Zy��X[�B��=����e�s�\I��Fюxvv�f[�m-;M(m�k�K�r��b�����	���,ݘ�糎��\R�.����D(��b�2om��]�RZ(���]iu+�m�D��4����;�ػpQl;wT�ֽ�[v�-�E�ݻ-]z���ly��,1�!qKm#�H����%Smu˸�m�]Jvg\&���N�d��.۟L�b��Ļ1d�6�:�2��LX��R�"J�q�6�خ�1 ��Դ�,�F�U�L�푷k04���S ��Y�h�h�:�R8��m,Мp��Z��<]������6l@"�cY�CV9�1��o#��::�}�b*P�G*k�=#����6��Wm�8��/����p6;�����c�cI��٘�[1�kZ]�l`R�-nA8��<^_3lf�����n$����(��s�Vͺ�ܑ��i���;����'��-����,\n��L�W3\z�B�s�c�.����E����	�ZnZ{.*�����m��X�%����s�n6n6�v}��7;x5y.������ܻqr��&,�s0�r�(�ɶ�U�]%U��'���	���q��Ů�s�k�(r�u�@;�v�Z�2!vS�Fj5�p�8s䲷|�pp����.�l�ʆ�1�<�Rv�t��g�F��k�q��$=��W��Z[@�hV���g'��������k��&"�,�8oV��cb�×��݌�3n{vv����>���=���t�]�m�r;��F��[�X"Mn��.��_���6Z�t��ܚ������qw(qu�Yh.v�ٽ� �	�V���֒XV#���˒Vrڜ߾V6!.k���OLI3�"�t���-7��WI��_{ݭL�^�����z)>�n�$����W5���>y�1t��	"�Ic\8�w��7QS�Ɯ�s�n�Zع��'��j����I%���:T
�����H�(�.����H+V����r]�Q�s/kED������I����u�B�Wϲp�r׾eM��H��E'۰JBJ@K�Q�Ή|�i��@��FP%�7[�V�a����r]j�	P�Ib�b�A&&��U�!���	)	-&Ĝ~|��P�Y1��B��w��Ba|�wZJRS�P���������,U���=�+`moT��}M֋��
<�Д&H8c�	t��q䓁�|��u�Fu��v����dl��w����ŉt�O�FV89�o�+�$�:E�%<�����������!%$�gu;����>�t�3�������$�������3�,�_nF�?|���b�>�sT/Lc��O���jQڻ�ݞ�Q�sI`J>E$\��<[��]�u�;���ܒ2���kx�+�%#��֛0;nߟ�`��N,Y�6�U�7 ]=A�7H���z�@�`Ղ,�����J9��:��vw)V�=����Ob�#j��?�%!%"���dE������lo��k��y�0�o�}��- �d�ٯ��8��_G��6'������68����l�D�l�9 ��x^Y��mJ�h*Z���K]��2��jԞ}��P.UXfr��k��&�Vj��}���{B�=X5��:��;I���|[��4���J�������v�z�����^8ά�}����S��l�S�=ݱ�t�P� $��*H�n����{5����
�����UV�ny�'��i�	G�*r��	��wg=�!UDA�D��& 1%"�m׵�'`�-��L�C�"5#w(Cj�>������߉`J,ES}ѯ�sb�������Ȝ���"�/��$�玷�v������f��o'�1�kUo�)��6ڔ�$5mb]�}݋5�|��!%I	)�r��H��x��n��y�>�6�%��R5e�]�ԚmK�!("�Fs��ؤ���>���ܵ�u,ө��_�u=x�Kõ��b��̶�t��ܱ�IZ�y�XA���u^8']�3���m�3Օ�ƗN�̎��7i�m����j~z�(	)$�"�!�T*�Sֻ/2�*����V�<�f�ۮRS��y�E���o��a(�A�vE�n�S!�Ӛ7��p�zs笙6�n�\�:ٶh�;�^�g$�~����~��J�KT�|���zeë��gl돒R���}���nm��������Vێ��'p�xom�����.Q3�Ճ?7kr>IJP>I3��F�|��ӬŹ���'�n�Ԥ�|�$��ݙ�ȄWgN��p��Ib�s�~��J�KT�'����:|�`�8ԩ�v���|��R��&L��ԋ�aV�E�o�l�zw-��v5֒��E>�H��Ⱦ�'W��)_�ۧCm,�`-�o÷M�P�V}c�BR���-VE�;����I���y��u��6�[�MGcm�p�`ax`�m�umt�L����c>e�ơ��g�h�S=Yz˅�qnQP#Έ�rr�<�����π�ʎ��q�F;kH��6�,�j�����a[9s`���0n/+�l��Ѧ�ۧ�����&�̒�P����p��\��<�m�� Ղѩ i5�!m�pҵ��)hH� ���h[m@n;��w�W�}k�K�[m�3��X���j��vЦ�qh���GX�p��i�ѡ������{�����Ut�/�w���'�d�v.���!� $���	!��En���x��R��;ѽܶf�*��}���I#Ʀc~��:��O|�/���"E�x_W.7X&r�\殝�M��x���?еHH�����ޯkK��������w;�:Ұb|�r�gD��'xsٙ'd�}$_IBI�VTt*�v�˹l�ZUQ�� �H����|7���>��_���ػ\M��b�͵�4�c�#t�����t���Gv���&��}���T�����R`�>M��kx�ٌہuU'i���_�%)G�.����<���s���)�jm)G~��Ǩgo����Q]X'L#��R�TE��O��ﴍR����.r㣴J�P�i�
�|3L��WgC�=���;�:�Z#����"�U%J�A�5I�>�dC����&��覡���˞LթTv�'�R�RS=]�Gu�r�N.��Q�
]�+tuQ���5��
�r�^o�[X;��>BJ�H��}#�r�Ό���'�5nm��fgoS�ذ��܀S��?$�	Q:�p?[71 F�%"�&�Ʊ�X������pdEѳ�	�1v:��zI���}z�/@	)�䔁�^(����T���^��{<!Ay�9_	"�/����4vPS�&�_H�b�ȩ���ݸķ����UY"�Y�����!l����J�\�G���W���Ry������K��۩�H`X��1�)�!�D�Wb�!��	-u{sݡlդ�!������6�WTX��v���v���hƞ�S�����ر���r>"�H��J�/�T"�S��)�k�s"R6`���UU�Vv���Q����q7����"���I7֤<<+E��n鼜����8ķ�����IH��!z)U=� 4k�7W`ؿ��D1���.x��3Ǚ�HP���y+�x�p�?__��������$�y�_Wm�g:s�,c}���,����ߢ~�PE$���\�{��veߴ^-6���b����JR�F]U��&�;~����s����S�N�t�<�ٕ5S��)�q�o}���J~IJQ�˸����uNj�� Iw.̾����n/!Xz��&5q�5�.o�W�b���v����G��������·�V�P�Ī2�[H�ݫv�e3	h����qN-�H�.�%���$_I�I�o׸_]Kjձ���޽�p^��_sʪ�
���t��R��H��.{����;Ab��F�آ��5F�#G5v�8�u�"T�+b7J
����a��d0%���}'}��)J�ۛ���b#��q�����]T�w$�% $�̽Wmݞ�Y���}��.˾����n/aXz�^@Z�$��̆=���3޶��}%	"H�e1�5�dob��]V(Vv� ��|���%��gy��_d�C�n);rʛo�"9ڗ�p�G���kk�n�H;��hW�D$�DqZHQ���gt/X���ޮ�����H�}𼏒R���I|�G���GG\T@�w{�R\{$�=�͹����=��F�î���ߏ�;ku��{[��ؑ����5�Տzd�l(*�Y�«X�
ŋ�dTt?�<�%�X��v�%ˋqQ�*Z�WoEW��ov��Fb��2�����>6w��z���i|j�$�"M�'`֛�o/�{'k�vy�8£����<��1�dݺ׬5<�Ɠ�"��a�0d.s
1s�͍��Z7V8=�dç����;�/���m��B#.���;���	��q�����hV���^ԍ�e�5�h���RX_�����-���gu���\0�Q�եK�9��$6+��E�u�)�r�������7���ۺ�Pc��>�CE�t���>ɨ>���!$_I�{M�־�V_>k�+�d9�[��;�qigo9��M��t�l��1X��O��~BH������^gt-����j��f&��/_y$��/��$H���I_���}_zy}$d��.�B����A�{o��{�,>��|RI$�M����SqE�ڍ�pOKYN-,��_�)�$��F�x����_Λ:�Kbv�jL�aݯ�[u���\OR˙�*�Ղ�
л(#T���A�I�H�ˣw��/"�&�z�霘Y��:ʳJ~�wrJ�ID2zf♘Q��x�řU�l�*��^�VfR�6�k�ctsX�Z�D��x�&��Y�/�;7/��6ӹ���F����%F�"/��]�Zu��?|="t{t�}]��B��>ֱ-Uօ����S���	"�HU�E�pd�
���|88Ʋ�ZY�y�\���J~J b#��������:�䔾��}9}�ܬE��/#.aD5"ށ��7$����@�U������OO�!o�Wb��P��	�R��099�SS����-��A��N�p��qo
u��W�2 Z�w]��v��W���a#y/�GA�RE���2��-!ã6ݹ���e�b��r������$�鵵`��M�&X������n�<�=�';݇�{�t�I5ka���z�� ��������m�H�sT��λ'�����r�o���fR߰ӷD��6�����R�rI�2MTs:�F�q<�7���$܂M���n�]����D���Yz������]j�VU�eR"N%m�f΅Ԭ����]~��{��A\Ӣ��}��4{�<nn�H�-�tn�]���6q}���FȝX�W���u^[y�y��G���7���{�s�!z-s����Y�2�g,f�X8k���[�b��ຯ:�^��[ӻK�����t���܎��Q��q�k776�]Q�yԥ��7�蹺��v������P�Gkirù���Z6�u��&v�X�T���U���v�WTʺ.Jˣ��)���ڮ�b�!4��B�%�UYu����2�et���x����;8�l�{[�&>Z��ŋ���WuDe���X9AR˫G)M޾�!X��l�Q��g�e:2 ��n�u�.�V�t��k^o�M�X��Yk����q�����]7��V��X�
�nf��ۆ���mU��[yU4�j<.�[o���U���n
���l��7[>�_N����l=Z*���b9W/���C�TM�ed�ye�!����;>����6U��H��#��%�ηU�L<0ᇮ��ܥ���ۯ�:����NU��A��B)J�ή��]I�;y-���yu.bK�=͍��A�䜣q�6^��m&���	XZ�	�����A]��R唔��a������m��*�ױ��]�9��n8+0<�ܫ��t=���δ��������Ȫ,�$�)IH��ch�v��f#�A�0�����h�J"��b�(Y���F�t�B&��$ssF�	(�2��F��H`���f`Ɍ�ĊI�j1 �2��AD��2b�:EM̑L�"M`\�MJI&�J!��	��JdQ!����(�Ȱ1F�PɄ�e�Ph�LE"S��ad��AjdaGv�Q�$�Bi(K&��4�C"����b�ĵ3���%w]� �BR��D	��Q���� ��H�S34+#����T�D $�\ݘ�$PdH���/�4��f��ڔ2�|�Oͩ	G�$�9Q�1л����������QHp=��9����rˋQ������0���w$��	$�w����˞�_��7/��Rs���|-@�����XڋΣ�}��_��6k�h!Fݥγb���|�x^��,*;�����I]HU���_O�� $��99�t��ڝB�_}�Yʕ;k�-��|���S�P�]�=c�9��u��N��r:�J\I�iӺk{y��䓺���F\1Y3�\��XQ�I:���\�wY�ܫg5)��"���ԧ����L�oe�<t#�	"c����kו��;ʖ�c��*�t6���g�ىA��������/���~\"���g���(N��.ݪȄ���s(��n��n���U}���W}}�k��!�I+IK��#�\Jak�z:��҂�$�4��%�7���RA�kQ��(����A�1nc��֓ilř�jx x��;C]�ܱ�l�5Q&hЩM�@�vH�R��J_.�����:�������Xnhԧ� �F��I_I�EǽAQ����ܳ�uo1���֡9/������:�#�Ԟ��k��JRR������o"*�k ���M8yIo 7��BJBJR���Hr���P���%#�͎���R���9��|�-T�ﶯUO�j�t�$��� �7}���@��1=�g���{�nA�{��_zE��$�vVc��K�ń=wWږ�]�9Ҩ�u0<X$x�*��chf��u�]��_P��C��S���]��ʃu�v(��\�Վz�m�(MбF�U`݋WdXԹ�Z�f#I��ո�Q�	��:p&Hf�n�k��ƛ�u���Ԝa7u\7Sqĳm�oc[�,��凷V����S���E�5a��Syʗ\�-��hKK,X�1,���vЇ3Lj;>����fֺ�5X�8�"�kB*[�g����10����֛y�p���Lp�N�r�]��7�S����.f@e
B�..��	�B�U�g��ͫ,kt� ��]L(y�z�t���R������G'�%��w7�,W{�����Ig�@IH�G�6����/z �R��ӝ{ӭNZ/_%�g�ͺClYqϏ���{"AX� �s_�	�5��Ҹ\gi���F��k���^i���𞏗t���_�A�۠r H��f�)����|A��C]@W����3�|���1yNW�s� �t� ��ໞ���>��j� �K�D72-��n�|[��jMC�me{K�����f��G�oz��q��t+�t|[�R���A.b-�����v>�7��!�&�jC$s=k��nKl��y�x��Nf�E�K��i�U���،}�^��(��s@Knh<��zj}�cQR�'�쬧����:�z@_7�(�n�m�Kq ���㢮x^��Z��H,$1f���;.�MK�T����}�Y���'K4%d���kwwt�gz���1��ͯ����mn�2^x?�	uW�zD�g����NM�y8Y^mψ%{��/�$��˼�a>\*vh1L��}�(�܊-Đ[t<�_�Wb��o2-{D��s��/5�b����8�n�۪���H-��4)�⨛��t9@��$��D�nh<��zj}�xO{��z�D�%��u�->���V#3;�Bq��q��۠e����>��"G�w�?G*�̏'+���;�5���Q`�̻�|=׊���՝Ӣ�ZoAR�Q��H�N��!ӽri��56+�E��J��~~����	 ���J0@JD�o�ӕ�o��qG�ox}A"=�;f�^Q���I�?X�}%$S�y����p�JD�ӣo�����hJ�	�} �W�I�JŃ%U}���(?Q�7� �ذA��A�)IP���y�pZn��q�F6��F\fR�[[�lv�pE��λ�q�c��0�r�(�W�Z��o��V�T���Z���+i��zi;�j�^�M�˓.��'�ǀ �� ��%(�	IM|BS��/t%6{P��7P���$��N?�˶����sc÷�}�>��8𡶲�������D�R�?$��)
QKGN��X#~�SB�^���D�)Z�=��~�W�(�R�Y����$����zX۝�u<��b$jܶ������%hӵ^�l��.��F�6gX �� O $�𿌒;)o���+�q��ry8�W�ݖ���}~��Q���X9�s3��s(��_;�r}��O9�$�$g�o�.۞ۏk�͏����Kr$�[�צ�r�vr��*�s;z��3+�#��xh�-����{��MO"u�xOxH �G%_%A	H�T�:!���_�vD}��IJ�|R�?��|y�ҹ�q�>N=��|�!g�;)�n|��ʛ������5�%�jk~2��(
�Wj������n��ΪA-�NmYg��-!�e�h�wG6M*��imE㝏U�\_ICL� �,Y��K��~���D�Z^ۙ��͏��@>q$7HIP��R1Lx,S���M�*�Dk5��V.�1k�V��w|��7��X��Z�I��l
D�]�^ ����<����$W����?MO�:V�'�E����0l�,��/� H�"IvJ@��i%�]��Ƒ��|~]"C�[!��ڹ�Q�>N<A�����'�2�U�ᡕ�h�p$�$����a%#a���7���K�Tn�+��ع�����v� |�H!�%?`JD��A����oIN=�z��wdIn'�	IMm��/z���`��xOxH'}H�}�Y3qX,��{�H!%B�)G�� ���rX�t7���"@�~�ةd_����q�A;�4o�IJ'��%;�����ۋ:���&�f)�G��&���Xe�&��`��;/��x��tşq���K!�Ŧj�<r��^�]l��J&'��tqcsd��B2�F������]$OS�rݵ�\�gd�y�ɮ�bM������hIC	u�,�Y��k`^�{�2��@5ܐ�Q��0`�-���>���;v�5�O�6�������И��R�j�u���ї�3�68�ܑ�]���e�t[�՛)0��;��\�ju��H�ۚ�MfiaQٶb�G���k�5�vzU�{#ݰώ�D�t�D�h!����Z�Ѱ��q^�ۯJ�c��b�4S�6q��Gm��3pS@����X����g���eX�̲����wq�3���xv�ERû� �H���j32�ʱ3/Q0����z:������؍� �� ��sCobߙ��z�l�ׄ���>;���(�뽒a`�]=�w����&��4>ʴs,����	H��b�2�;$&���E��c|�z#���7�,s*�.f^�fP���ܭ���״�� �["�~� �"Fz��ov�n��7���ޠA�vf��k�Q�dw;������$VA�d���^��������^�������	�]����fhәW�<}�����~w�w�?�_y)����VS\;�9���d�r�ϜN����m�b/�ϯ}�����gߌ�,�	H쥲��+�~j67��wY�f�d]x�ܿw���R$�A$�"@�%�M��Un�En�Be�С.;�Z��s+��cUvtd5՚FU�ٮ�N	yU��a(���f���FP6�1D�q�e��Ǿ ��"FK�;��w��/k÷�(��H!8$�lq/霂8���_X�}%}�������L�[^��+��ڵ�z>΀<T(�~ ��O�-T(sv%zu�PD��o��/�24:{�s4皂��ǁ����.��=���A�ȑ.P@�$�`�R��!L�捋�?*a��zk}�..sùH���$���]�~��������qj�ň˫quێ�'.��x�� ��3���N��^Ѩ�Lqk����"~)D�JJkk!�=�/�<K�k�z���j�N5�(�����M���t��DVe�Xd{���)�뷲5��,�~j�7 ���D���Pw�7!�=I�0����"A=�BJ��H �!�j����U���6�ֆ�ʭ&j���&�<WXU[�!�,���Z�9�R�D��n+�a	Ȋ�ٝz�Y)b �iD��W�6�zm��S���ܽ_y��AJD�BJ��O�(���d���F ��YQ�(��j�u���d�x�b]%�� �l	Tﲗ�eR4���W˹D���% A "V��"򐰾؁^��n��W���:������s��>J �����6�8�q]���ĕn�9�[�WF�m��G[&��9�ڔkvu�h�31R����}�������AJD�8����7��0�M�oz��/=M{��y�"�H�F�U|~JD��I�$VA^��?,���~Ԉ'���[y�vOQ�!�^�	����B�(,{�Q�����P'T})H�BJ~����-�c���%z_Pqt�(6�R������G�'W���R���RS@��H~�{� z�F|}��R�#���{��ߗ��fo<;���F-���{���ne�fu�
���rtn�uv��ZF�"�`VNwK�	�X��I�$�:�VP*�Co�ϒ�ar:��өs��V6j�X66��̿|}�_wG�E�~IM|AJD�R�ʧY���Ǒ8Ś�����;�}��ly����w���$|�Т�H �#5��G���svj4�
��dޘ�ݹ�SYLպZ�6g�%���GW��ܷ�Z���}��JD��DI�"_�����G=MI�����ӫ�����ھ�N���Z#���̲�e���<�x�W���y;�$N�q���^u	��xw/
��$����'+1<���"OlI}?%J$�RR}A�s�����Qoe:6�/�} �d	 ��Т�O�R$��AV��>�
*܉ ��_�WR�}��G=Z�5v�_���U�m�������"�d�� �%� �Y����;�%�`F�ޗ�ڽ%�Uy�ܼ(�A�T����)��sY��=���ދ��S{�J�{wq*���f�����ݶ���x��U^jٙ��욡�%d��l�K�̈́V	�R+�����j�A��;���kȞϘ��Od�bM�{j�X{]�+�jh~73_�$�W}j����b[��Y���b��*�T�I�ӏ��3As��"�����Ø�c2��{�H�w�k�	��ty;���t/U7c8vRˮ���2#F�T���u�\��V�+�6�t�V��fBպ��^�`������1P���{I��5Z��2z��jmu5����ff�w�Z�����Ϧj"\����w�q`�V�Y�9ީ��D�F�*��]VҨ%�+z�=��w![g��UfE1q%��8�� &ќn*�XY�K�
����n%O'eŜ��^�6���F5�mkB]�1����v�����3��d�gCJ����{��w�ҖA�c��dim᳄K�3.��9Q�<�gk',En���v*t�+�:+rJ:�g�;l&��{����b���M�F1	ݕ������P�3I�J�*[w��f��U�c'^��k+׏����\��n�[ڌ��[��ɸ��d��q��3��%��h1ngu���K*�	��̱wRk��A%��uB��\�P�$D��#,��ʺf ��K-���[e�[32��ưy^t���7׵T*b�M@�8�KzՎ�h���8��C]��D�v1QL]�9�b_�;����B�H�;a;��O�s�%u�§Z7���{"ʀ�[ec�K��%��\�@�e�Y�wz�����<�@���TCh( ���#&R�M�lh�R
{9F$��,�2$  4c�PQ���R�&�CF$ȃ�Dd)K�����rH��d�$H��Ęl�A�J�`� �!Dc$  �QjA"()s�3K�(F 1dY��P"h�����%A�0@��S�]�I�IH!%@R&LF)�YD�i(�C\�"da$E#4���E���Ʌ��)	&0��A�����dI	� h3 �Q��HC � �!ŉ31"Q�&Dh)�"I � �!)�	II%J@�F#dȹ\�4��#Ϗ<�z�8^�`����wa}� v\k�ݭzxw":�	��Z�Z�:�P��G���p��%�����"��6̠�3�b�n
D�fYv��65�8�H�q�]����N���ڷ3>f:�x.�K��!�����N���!i-�
b;.٬r�ٷٶ.�����:X库j�ו�ڂ3�q��E�z��/�A!�{v�!bY���uЉ��E,��i�!H"�'W�k�Y�>x�%Ʈ{6uv���8�Tv�ՖWN3��l��v�r���]�1�-�!��x��2���qpQ��R��dܝ���V4n�k)�q0�h�Fme��A�F:��f&�����Wa,HI��D�sGB 1�u��$�&�+���	�,Dt]����g��;6k>�up.�5ڑ����F̉{�h��Լ��v���&j�j�t+،1˰;2�j6!M�[���K�S�ee�$�C7(X�Xsn�)�i.���)u�=m��rŗ�M�Q�/Sui���J��U{p[��X�<�  V�.�.�4F{	j��DBCGn��Pl�;\��kv�&�hL���-���q��; m��o�^���*��V.�L��B�v%+�c���Y�,���1^��� �y��sN;�ї�mtLJi�x���(m�c'd��[�Yd�3e'vp�r>.�)D���Dئ�3@�]�;q.�jq���Z�1����E7(�:{mө{Mۭ��Z��a��C���	sgu�NS�w3ۻ��hFx�vC���h��/d�YL�e�D�H�4i�H���@n��ѮO>Z��];�n�f��`�H�h�.̺��D&Z�h�v]�§U�`N��ل�ņc�3��Xa!���4ѩS[ %v���Q��tV+��n�Gs�DqË10M6]4��mz�,=s��vI�v�dv���p�m;.1��ŗsnI�v3�Pqq�ۺ*�Tٞù�]wg��hwE	ٝ��L�k�0J�Z�������s)+L8�q�g��(G�zB�ڧ�9��ݻ[X��������Ktn��M�3��UCCX���^��1�Ynܷ������n�`��68�b;d�7)b�8Ԑ�`p��0�b�s�8z�����I�"s�p��7d&�K)e%li`�Ch�^��M��CWi��ë�`k9�ۑ�.�GGU��#������h�M5��Ҍe���/�g���dvc1i�[��߯����rcT.Ҷ�%�\ಆ�Ѵ�|��GYd���q�
Q$���܍��뮳c��4�W},���ƺy����G���Q���d� D��%"<;�~Y��wu���	�����f���V��^����O�7�Jk_?g��W�,�1����IP��H ��u�$���S���)'%�u��ܽ��I�RK��P$Q$NUclTn{��~��q􂒚�����u$��	xG@����;�M�_��z�{�Q�r$��@�R��H!$3��][�}���):}�Ԏz��j���uzk��H��O���ʆ{�_^��D ?��:ݠ<�Y��n���=�A�Z����6�k�-��>�̽~|#a����!)�מּ���%�MC����X����k�4��D����JD��H �RS���e�\�_ɺ��VM~��nbУ��WN���/w9�e0�>��'/FVY�oҶ��ڰD�[8�[���"�J����!�wϣ�N?L��S��'|�K�w�� HZ�QJ=��+b�B�ސ�
���%"A	*��JG��}����cܔ�}��uy��F���;���U�G3/I�G9����'GUC���ە�Q����/�Ӟ��i�u�÷����#���eT��A�7_�H��J>������(�ޮq=B#��V�3�5W�g�t�]I;�
^��A�!5_%)HVw|�G��o�fﯗ�ϳ��Ɇ�F0��2�r��,�bуm ��#���M&��Z��~���������P���|~JD�j������ܯ[�����`Y���BWW�X �h ��2E���
P$�^�(��F�U<�~ �H�9�o��=+��P�3÷�(��O���"$���|^i�{�:w)/���Q'���_{ˣ�j�l�Y�c!I��kl�V�v1;cxR[��v㫷4nݼ���V��� �4]^�Ѧ�}sݤ&ᎎε:�Iڸ��2^Z%�3�v�;���Ѡs*�9�X"J��"n��W�<�2k�}#}"A�?RR/k�L�fO��z˭\�x~+�k�D�5k���
9q$}�4JdR�$��E(Y=Q��(Ǉ1½"Dc��v��6�:������<?j�$$�W�)�����U(��c �B����[xY�v哚`v��<�HvHZ�!(m����;�lx�W���D��}?��´n��껒s̔�#�to?;�a\��J� A�
:��J@I`���{���c�Pd{v�㾑"����<��ܯYu��Ǿ?/9���#%4�u]��'����A!%B�)D�BP+|l�E{}�f��b*�ӂmo��Mjfxv��A�"@!%?PJD��~"8���/_����ˢ���h��q��˒s�D/
�O��$m_�ٞ�z~�ASɻ�t�o&jY3�+�;s!{���ɭ�`�1��=b�E�9u䩷շk��f�}��ۋ>�*�F�:�ܹ��	(� WD�} I6���DC���_�U�f�	��N���<��ز�e֯7 ��4��2R �"����~�<?&�X����'[�sn8����ڷ���\tŲ�12�\�uYM����=�'��QJ>��O�,[���)�9��nxr�}A��B4h��4�G�����2 ���"��B�
�CN$�sU�7;�wN\��{�+� ��AZ�_�D:΋����D@�=�_hc����Yi��5̳�����K��ݪ����T�:K���y�W�IJ$JJk��"_e�=�큤�:�}BP$g��~��)�+\�����W��2����E��O �����(��)�A	H�R��z��Uc�������uVL��؅�]�?o@�A֫��	H���Ji��:�"��8�KDx�B/*rY��*�_m�K�vn�ws.Z[�y�S�곢�8tٔ��3�%��U57��z0a���I(�O�%���|k��D%���sq��گ]�ˋ�N�H:n�݁�v�E��n��U�c�ݲD�!4�U����N̻+X�4��<�@/�SGc�s]�Xѝ��Z��op��m�;=-V��y���^ÛD���r�8%2.n��	�j�0X�n�8ܖ�{����\uYE�rF�s2k�)�ۍ����r��� %u���.������r�r��R.�2���a��Mӹ�n:�k��n��Cz/^7����U�L�f|j��"��y�^]ϖ��:K�ǈ=}�9�kݫ�o��x߬�{�b.f^�f\��Ia&u[˅�(dj� c����ȯZ��g�.�}T���%�qv ʱ��{� \�&tVPFJG�"����}�J6D�����ˎxaxW@�/�'�MW�F�	$�Py>cX����y̮����7���({y+�^M��g�]%����W�����<r'D�q �
nh��	 ���@�C���tN[�$Tȑ��]<�<1l����?�R ���]�%
�`�1��W��HU������Z�N���|E|�V��x�l�6��TP�]�ʀ�^�?� ��H��ї����.=LB��y�kݡ���A�{(P:�@ �"HIH��O�j�̾��9�7o��uz��W�����ZEé��!�un��晋2h���,��Wu�*��;\541"�7�t(M��jR���9*��@���]��.w=>��W��J� ��
Q�e�0x�̔8�S�nH �$BJ�J>Ĥ\���V�EB��e0�u8���{��˼(��3�_$���@�H��/���_F�[�RSU��_
su՗�%xW@�~�?��t�[vfW���w�BI�d���/��G������}{�$?^�72����]j�q� �4/H�
Q$RS�+e�S��}_Y�����ml�]�+]+����xzܵF :��/Zժ��E���c��}�s*���H�K�������xr�]�����xtE���A=뿈�}%a�d��P;��C��<�;� �����m��r�չů
�H ��	MP�R��ڜ��y�e��oA�{�b32�3>���Fd���G��=�wq�;�%*Ȅj�]]&9]
+�VH��v��y]�֫�۷c����(߰�'�K���r�\U�
(�FU�]�m�Y�T�H����\^mj��/'�����/O�@	)�{��{����y���g��=�\Fj��*�oF�=gZ{�ù�����?=��;w�h���yB� r�%(�A%?RR$��mX,G ˼��{ˍ�:�N�K�+� �� J�B�)D�
R���i�W���᪊���h�D�	�h�Ի&���&�`���g�i�������_W�\@/���I,_�D2r�ݍ;��]fy���R���a�V�1���>�"G9R�̽&e�2��u���~�ݯWC>�A��7�_r��g��Or�;��c�T��36~�uk'�_�\{ږ�<��")L�d�Ȋ��� ��U�ɜw}}p����/�'�Z�QJ$��X(m\`{υ_.�A�� �j~���n�5ۑ����3���/M!�<`��ݙ�[�w������{��B��\4�tW���K��I�o�ْ�Ok2���n���v�9���$�K���v��Mr�=
k<4���o+H�("$��*�7��_��8{:D�z3��Ͻ���ܯ�G��Kr$��W�@��"��n|8�f��U&H������;��va�c�WY�]�WUC�:��>'���� ��"~)G�
Jhm\5������,%�]n󻸨���~����H?% $��(�6�lw��Ï>�4W�p$+�Ҋ����Iu������� ���?�=goB��,ۚ"�}�G���49�.fYwL��ti^��{�KǓj)c��|�(}蟈#��$��2 ���#��~ِJ�-��� ���?��W���=��^ސO��P���ʙ1�X`�A5 $��)D�AJD��1���k��}s�$;��,���b>��3����R�� �IJ$L�`}�r���woG�0�O��9�Q�cx�ʫ��u��qC�Ʋh�M}]����j�Vc�m�ϫ3b�+p"�v�������U�M���V��I i0����s<�]�n%��3K����Wm4�[mJ�rad,X\q8���;\6��q=�m<p aƎ-�ڭ�2i��[1.�%�v&�Pnݭ���e�QM��\+\)v:�:��xw%�}R��lb�&;X�X�f��қ����:bV��ȵ�8�<7�ǵ�-vn�!_��~�3���-pr�c�k�O0z1���q=���n����ma7�����}~�'~�H�R� �����}�;=�ARǕ���7��}���6ۏ�d�#|���	IM G�K���A�j$@+���h���ڞ�̉A/
�} �t	 ��Я�Q���>���zw:�I�P?�H H��h���,��'������5��ٿ~��w���;^E�����ˎe\����DU���giL@d�(P<��JD��,^�=ّ>%,y~��}�����k���֣ܲ�2�#̹�2�P�����]�|�9sC���c�j���/x�v�>���,��U�s,d'�ϟ�C�ye��,^aeE��mV�#m9�j�[-�c,�z�!1��	����m��[A;�_�>��Y���1��`D�^T��?Oܢ�"��$2P�P�B���hC������%���t�(����,}4��)il���F�e��Wrǁ��(ʳv%7�˳����wi����>�R<�K	Z���5�U���|�@�}��H$����ș��M��� �?W�H��I�%-���c<&(x����\�P������/��}b̔��I	*��գ ��}8�H?zD���|R� mZ����=Y�}��R����)ߣ�Dj܉�zh��A)@�?$�P)Evr�B��t�_	H�9]��t�׉��/����>�}!z@Jm�D�~�x��Ts����o�x�6ȴ��c���R�hj�������X�Y��އ��ڎ��Q�&'��W> ��H)D�))�g٫�u��z�d�+ºw�+o��f��>����Ѩ��,̲�34jfU���|�}@��W�5#fИ��V{b�+3����K�@�7�'�>�{/���o�j�'בּ�3,��U���~�{���8�>�̆�b�e�^6�ٙ���a(�ՙ��sh�#,%j�U-��=L��]��Ŝk������z�iH�ζgU}�-�*��;�Z���U��m�͙H�^�
Cb���(ũB���s���tỷ0�������2�/�G/u�3@�h���M���q�������Q7yu�����Y�c��yXU�c��H��l���WS6�%@M:����/-�����wv�2�f!�{O��W�F�z�Eo�����	���N�#R����gC|�-a�%e�E�,^a��]R�rݸ;���V��OE۵ʓ�\]Cv�,�+z��Zrm�M.7Z%:;���rY���<��-N۫*
�r��t�e��)�Vo;sV�kvE��7��X��FV Rv_e.��y%
��Vb�"$tHղj�)�p"�2,�WuUTS��Y�kY.��*�W5Yw�nه�:e�|�P���g:�l
�Hyjx�ڻ^ȭ�푚�.`p�2��܏�j�A|
�rɖ*��fLP)d�+���j�����R3�R�$譌�rm���-�BW@����ח,vg��mL����JHڔ�؜y�p�7�NNS�RM�Fim7�%��rL��Ԍ����ˮ�]̼��v�aW�+B�"Wd�_i�*�]���n���U���1��j��Q�]y�i�Cz]�`u����Y#4�鍻�i��f�~�
wNY�C�#ǩʷ�`���adK���*D#9K	�O���&�+u�nfԭn�e�k7[Iоl�e�CNQQ��V�m%���r�`��O-R:�*Z�����L�$�&%�3Bf��L�a(�L��e2!��a	��&E�ȓh&���qJe&d!ih�d�P�D�I3
(F@фD�P�E����F�d�� d�b&D̄3P�1$0�bM1�@�fYC&S	3$"!1��Bwr	!��% ��%���H��,&�%�"��#1L�I#2�J$c$�P2$�В`�$M&!�2���D��&��$�I�S!H҉�$��*2��A���`��wtcJI)B0�FI*LL�����*4�dd&&�Q���Q&)$����&1(��A"����_�����>p}���}��A��H+�J~ĤIJ$�����g�U}U:�VG�A�"	�+�����u�׽dd�+»�	ށ?T� n
e�ıq��D����)H	/i����ԉI	������Y�}�D^g�h7�,ʱ�e���^�e=^}�ИÞ�:�Y[�5$�N��[����ٵp 6��V�ZִP�֊/����9�Z'��LQ�BR'ȬN�]_�7��x>�|(T{To���ո��Ybg{���YneX�Jh/Ǝ�ww�_Os��]����ru��]�P�R��c}��:����)D�"$�/�(V����nT��1w��B�ȍ���t}�צ� �H)D�	IM����C��4|^D ����ф%ȫN�u[�ᓍ�p}~�~>�}���^\��-e��%�vJʕ�y���+�b�Dz{P��]�\$���73��ٶٰu�=�ң�r�;k��_�&��5�Y`�U��e�FfYq̯~(�S��)��0���S�;:����P7�,�H�"q�ﲊ��X[����-ʑٵ��N���N�pv��z�J��U����_ ��"I`_�PARɏN���K�;9Y��)Y�apԻ�=��.z�3/Bf]�s(�>���D׭�0_��x��ޑ<���W����ח���@�}���ȒY���Y7��'���,����O�E�JJd ��7F�\���1�B�wٳ��ސO(;�B�J$BR'�BJ���7��
ǵ��H#�D�<��┉�*^����=�y��=� �R���o��Ozeog�k�F{/BfXX�e"ff�es��4i�(��J�.ϳ_��W�}�[Y~�>蟈>r'�U_%�o��t?f�ު۶�FFU�v���f�A�]���J��z&�|󄷫r��ҧ�7���b��W���8�ͻ���
[Ţd�g��VW���}��]gRGW�fř,݆��s	��r��.��5ݨ`����&d�Xx]�7dd� ���m�8���.���\���:$��Q��:v:��n.n�v��vԋ��4ل/iW�<�Hv��ˢ���F���K�5��׫mۂը�ё���afc���(`��lZי�u-�7���F&�B��Nz� mAP#s�0�Y��&-�P�iZs����k�ڹ�ն!Z&�!�tf�K1�Ȕ��y�C&�Y�Z� ���?�'�Q�oסe�eKs2��;�Us�.�齖���ε��˗���~��/�"�"$�/�)Lʭi��ս�|E�����D���N�(����^]f{�<%/M�H�R��͖�}^cAN�n~�O�A	)J$��R^X煑z�/DiX�c�W�n����<(�Ar$����O�(�E�s���ʪ��΂
�{�� ����8��L{�ݖ��]�'�p$9��.�������D���+�$A$ʧ�(�몹�b�_�KE8�:��Y���^����	)D�~))��'�#=��xol�Q;Q"�Ms`	5]�����tۣ��^<Kz����ͺ��7��>������JD�V&��}y�8��x�~��_se�:���#=�X&w�+�H)D�JJ~�u8��*�e�]�Ḧ�E�ڗR�%#�b�b�6��]�jt�ky�:��K�U�zU���r�N�3dd\bR�w�QյU��i�����r�u>�:<A�M!�8��&=�e��+� ���wz� R��r/�Ȕ#���w�J_�D���"�޽x��گ���4ƨqMM=���tx~)zh���D��A���J-���#ٝ.�A��
)D�BR%��7���=p����.�P �Ă2�d���������IJ>�RS@����1)�k�`2�п���ǽ���w������Q�%#uv@}���&`����_U
�����u�\�yl��X%�^��I.$6����~w��}@��$��"~!%?RR$7n:9�O�ʩ��g����2�Vy�cq�(qȐyĐ@))��	L�R�${=Jf�N��|�8��Hh�M�~�f�y�a�]r<e\�喙����ws;�,wڱ��@�� �A%9%Ǣy�ǽ
���^kK��"_��,�@�ϫ�+�܋�}q����J��]�^j�+��xUۤt;�2chZ��.��cB����*{���w»�	�H;�_%!)�!%T��"�.��6��� A�6D���|R�>v��[$�������tx�R���y�7��~9}�P�ρ	H���$�|�d������M�p"��������᧭a�}r=���"HIOԔ��>���#��5E�L���$�L�i��K�v��<������a�c4wEܐ6��L5-����( �d���)G�RSZ=ߎ\�������w»�/�o��X_���:�E�HJ Ie�J$;������b�YU���7>��>�+��+;�<A��鯈#}"JQhW?`�؀q)�;&A)@�
J� R� ����1ۚͿM��z��;��KZ��}@�|���?��_%A)�o���d��� �� _W�����uފ�|�5����	"/-GE�?i����Y���{��*�[����+S�N7H٨��ޝ�����v���uǋ$���s"�r*������;��p,��@��})H��I_�l�з��F}�}7"E+ݗ<�=^�M�U�� �S���
Q������P���Cޣ}3FSI��Pe!��׵q�t�)�f{da؍�mZ֍^�cz���G�绣Q̫��"G��T��fᕭ�y��Hκwܖ�*�x�I�D�ڪ�)H��Q �
Jh9n�eu�lP4�~?g9�g��Wދ���j;º>j�#yP��Q���tU��4`��IyU��>J����(s��:/.�.���nT6V�Sw�~�~+�h��%(j�%��<ɦzWl�)Đ�	h�[i�G�v%f����@�8����9��ERc|�� s��� ��� �?%D���m���~�d��sQ��<y�������A�D18s����~9����&����t�g<p������k�fg�|pG�F�v���06"y,�b��:��Z]�,C����5�U�PS���WwV(�1q�v�l��Ѻu�&�	�v[�y�)PHh��_)������/Z�����nc������񃦷�x�ʹ�Ԏ�j�L�@ܘ��qc,�tt�B��i.���z�XOG>γ��ͼ)�83s�m[�@`�=n��V�� M�wMv��c����a����vԛLp�gQqܗ:n�7�D)�3lp-o	4����?_���==I��pe��H�[�q��n�c ��Z�5ٯK�" �~
S�@��}+�$���A)jߪz�S��]�t{�=Ad����`�ҮT�����v�D̽&e؎e��>��u�8�A��+1,,{ۛH���>ؐ>R'�F�b����u}�H }���}	FJ@�$Oo'��'jvoE��yD/|�5��8A�B�J$~JD�����M��(�7�1@�W"H�U_%^�}0�'��o2����	[��lMv� �>�������D�A�t�!)�JP$RU�P�k�
��n܉�l^y�p��6&�k<l�|}� ��"HIU|~	H�����3}�1fD�h00K�+�	�a�gT�QI	�[hG��33To%�*�5^ˬD}�ޢ!��2�"�)��;�+��盪3�w�zx����r�����j�|
Q��"HIH��Q?�9��f�����/,Y���˚���iΥ���<o+y�0i�ṫ&��+��t��λ>�a/�+\�;��޸��������z��a0O��:�e߻��
�M�D��,�ب�iQZ��A����=(	"�J��@�����LD���-�i�-���=��$�(%���)�)D�B���λ]덹��M�|�H;� �IM	�^>u^��n��
�>p$���d�;g=Q9�l�g�"Iv	��H�"I~���8y}��]���w��ȝN�/���+}?P�H�R�����{eT�2�>�
z�v*���t�
bx#qvr���K��4��5[��V�K�����h��4i̫���$=*�[��]�۲ڿ����*.�{���4#����E���$V-�#��ϩ��nh	�~�9�x*��wT�w��8A�_%��^2�o��>L_��A7%� ���H���"�Ĉ9���{��Ⰲ�[q�DN��pTE]Mf=��9U��aL���jd~w�[�.��<�i��F�!�l�N��vU�	�:��GW��Z�3=�x���_�����%Cg���/e�0��#P�yGҔ�������{3Ֆ��>�|(폐�"̩Ӷ��I�4��U�nD��~ ��������ӧ���s.hM�Ź��^����} ��Aw�P)D�JG�P�����DG���I��F�\�5���k*݊����{pp�s��F�Wv��
��{�`�{�=�"Iw�D�]������Uk���tx��wV}���g��v�ff^�̹b�PWn�ѥ�u�īV��돳zD��zۺ�f`ڲ�/��+�dH ��"@!$ �s{>���f~wY^��!(�(�))�T;`������[*�b�=�R�_zA��o����IA D������{Z;���_H��}_���9�cy���X�3=� ������mD`�$?d��^X���esm�w:�QV�ӻ���w�g><Sy�jzN�+��{�M�B�-S"*�2*#=W==,Ѻ]�$�W^}ZϾ��N�?%�	J ���E(���^��$^k�Wz��j�t�g���D���@I`��R3�7�	�����κ��7V�� �����o4s�!ֶ�8Nn��v�v�SZMU5v��^F;�פL�YneX��5��b�>s��S�{j����v櫳��WM��_P�Z� �"A	*)G��E�eUgN�Wq�ǀ�\+��"{^8:����Uc���t{���Oվ���'��]�����;۹�Qq34i̫D̳��#fߠ��G֞`ܰ�>��P'�V#=�\L�֢fYne\O��>�m�~������<�O�)����V�|ͽ��K����{�5�v�=�"��~ � �O�$��)H	%���/���G�2sG�S6� ����}�#�V��w���I?�B@!$�RB@!&�v��[n�ڭm����[o���km��mV���[U�����Z��[U���U����j���kj�$�BIR	&�	 ���涫[o}����嵵Z�{�mV$�B@!$��$M�H$��b��L��Ə�e� � ���fO� �'~}��   @U             
   
     
 P@ �  .� �T
� �@�U  R�
 E
(UP$*�A@��@($� �@@(�����
�H�QTIT�QIJ���R�%JT��J����UR*JA��R�*!	
�   �TRDR�	J���@;@@�-R�� 8s�"� -�@/����@�.�:���"� �@v�UAB��B�  `׼�E�΀#��C�(��@9���0� ��@1{�z

 � tw����0P�砠���w� ��@P
�  �HAE$��H*UϠ�4�gCͨ  w���9j,����!Nu*�w��92��!�䒇uJ����nm� 
��| {�{�8���󠓝"DΥ35 7c�)n��ۈ�g*��UvuQFM
�6���b�P(AA���
�*��Q*P�	*P�� jGR�9���&UUwRM�9%r1*��P��ܪD9Ҕ�ܨS,�T�PUP�P}�ܺ�}�!{��W���xJ�o^�[v��ʼn�U�wE�ۅ	F� N��w��Ww��	[n �z�OT EJ � π�"A*	R�@�9�����TŒ���w/f���o/fT������C���&�"񷬥J�n*���H�*�ǽn��o^� ҅IT�  �}���mw�yTUWq���=��V�Wz��wX:"-� s�J;�@�2 n�q�t�݀�@B�$   <�%
EJ�QUR(�)>���b(l�r*�� 0꤫�lq ;�8��h
Z��qH8 NȨv�@��(P�   0@!� c��p:Q�h n��v��� ��^<$&��z�(��ѯ{����|P5O�I�*R�  E?M�&�  =��@  6J�BR��  $�IU54�&6��MDS�%*���  �������W�	$�Hp����7��~���~��$$ I.o��$������Z��~��ն�ն�m�ժ��W��&��I�@������$J]톦�#�CkbK��j*g^^sH�Y�P�iiY�W�@n]�����gm�!��FU�ͬ|�U��~���:Q�0��L�m��U�gE(m�!pji7-����ǂU	r�Yx0*d`�����N�<�lh[�n���r��WyP�V]��4U�)f<�l����K1.a�YN�ʊ�Pڍ�;�����-��,0`�����Y/]��ٮ񜰮�M�%��f�`�9�
��I0�R法�a���-�nHl�C��D:��X������KW��������Dn<��!#�aYf��*��G^]'�Ww�e�6�n�ݡ&�2�V|�"�J��@ə��:�t�v-=�5*��܃ J��ږ7w�-�M�If����;Yq��s@�C.
��b(5efi�2ӕx55hf+��E�b��[�1f4ԑ����ښq�o�X���t�k�ic���@����j//K��ڙg	�^lj��F�Rm謚o��b�"pf�vr��vUݜ�zY��L�m<Bb�0��.�Yy�/��Y!p2�i�;�j&j�eHVU�y��2�j�TvF�fhJ������.�#-����{e�le��j�Q��潬I��Jf�6���i�.�n�Y2l���ɭڧKtٛ�P�,�"��B탘.n���-U�P�A�u����p�v+iŚx�{��U�QZ��j�̴�n�J8�
���^�/f���ʄ��2�F��XZ�V�&c!`Z��]ʃ%B7�u�M�c1�]�h�&^���r�9�ZZ�&�p;T�1�\4�h�����T4�E ���{�a�;fԔ5��4��5h�E-�F����Ym���qM_e�Q�	[3*b7r�~Yxj���2��+DU�{�����׷nХv֭B���f��nƋ��;�u��^�#�`	J�aؚe���3o6fyhS���mJm�jh�N9�e ����[�Q���LXh��K1��n[�M������ރ��T�΢��zrXڭG6�l�#kr�m��(A61�e�ePѻugs�k.�1yu��R��V|K���&5xP �Cv���1I�*����,e�;I�ƞ1�9��n���ZV��6����J��{��$4� ��]��+���hл6����YA�)�ᬵ�� ���1�Wm�9�5ĊY�5[�YK~0't��ҟ�QF�ond�9)�@n�fଋ1ۘ�J�0g+0��Si^���ҍ�Z��'Cm�W!
S��xi�,h�������1�.�VǕ��x��w\���)ǔ3Fi�OiV�Fkkn���їl������	���Y0"\��K�{f�$�@fᱛ'{���;Q�Q��K��VK���h^;zwt��[��X̧4Xj5��M����jV5����f��-i1B�����N�N�5a�t�Ӳn9�4�/�k���,�eC��ښ~Gp���5A�5�P
a�`���E�)+w%e�{��h�\q��hψR�Y-�V ���q��[I�����-�1��U�\QѣX��J�v�ۦ�dvwn���Q��3 ��+�G[{u�	x��V�V��[9�]��f�y���l�h��Ʀ�Ӫ��b�,*�#���c�Zv��(��@W�%u���欅���sL��Q�7#!f�R���v�k�ٸh�Zv�$U�%�JՂeͭ	���*VI&;�\���1z�B�45�w0+u$BK�ŋe8��yf"�cܸ.�s2;rX5� ��7�D�����Y�$�,��򆿷w�k���������t^m=.��Ŭ[Y.�cEf��"���"��p�t�[Q�b���i/�ol�6�[�ϤI�mnX�Ml�p�y3rcd�<���E#�V��C��xZ�\�5g]7A7�K׻��#���3]@Z�51�{FɁ�PM�Ѻ��ڛ�N�N�5�dg1��.��֓xS!���+P��Y ;و��˷X�>F��C�˦�,�ѺnT�!��Ӹ��x-8�u�B6*�S�6�P���-e<���o��I��L��%�̐n�W���]�aم�\��̽ɚ&=�ya�ō�2�������{LeA�5�{c+m*�zKIɮ�۽�?ԡ�G-��X�ic��;����$RRq��ƺj�V\��Ո�K��+tˣ�a��h�kmU�۬/.)�`ݷu�����R��a����@���l�Ǹ�X��FZS٭pb���(��X��Ǌ�OvCn�j��}�������&�^�b���m�*�%������h��&�jش��4]�2҆�����˺�KF[h�J2[��Dцn�e^��*�´ӖC�.�Q
�.:���3B	��nn���uA0��ҶM�<0��c7B�bה�ض�T�π��K�O�g��]���E�ݐ��`,uIx��2�n����m`p�WWV67zov����,(T�V���٫7�c%9˛w.3>���mKV�B1��N�����@�B�F^Y܄�l2��-��h���!�i\{�>;0mգ�yMM�y� @T,lGm�+��9�����sn-�Nej���5�5Y(�������h���9Fkڲ+e[��[�ǩ����k�oUJǘ���Dd�lffAƷp�d�ǗWQ�Ҙ���N���X��TEH4(uc2���V�E\ە�F�nV-�NS1T����Y+b՛$u�HY�Yv���r�!l���gN;56V"�J����3US^�V�h �Y�tۨ����c�{��c��e��,���ܘ�eAhٛB;�jj�c��t>��Y Z�H�O2��:/kotF#�S.�51�j�Z����3L"�M��q��C6e5�Wp�dp$f�WF�X�M����1�K��Ѡ�����D5�{m��h5+*�]ȝ�)j�˷�v0w��^���R���]�se;��N�һmf��v��''.��14i�Wʰ�-j�x���GA������4�+��ֶ�40ℋ����̵b݊�vf���b�㠮��Z�%@[b�d�$�
���I.���VQeֈ��1
�ٲY��w���2��M+� �r�&	��R��W�Q��J��lɆ��{*aI�TZ�b�p�L�	d��ŉ=��!QZ;�Ve9�b���KEZ��Ȱ�w���y�iƠ��ժf��W�5ª��jf�A�nQ!68��9uu,*t��&�pc-P���S`�ɵ�6%���L��'0f�e�^�IF��LQX��4�四#�YD\��PH@4Z���ԢSϤ����n���b�û�Un�R����3qk��i݌��  �YN��Pl�Ւv��ǚ�����lձv�k`�DV�f�E)���+,h+r,�E�ٹf�0a��*�P ����KpT�9C�N� c�]n��l�cXH�u����u����+t�zm�b^��I�1Uޭ7!�ľyw��ܩw+q	1��#�&.�c۰L��-�#d��Feݺ�%ǻ6��,�em���ZL�w����Gv�X�Sj�BNǡ�q}�PE�OY���u�(`́c�v�Q^&V�U��Jub���9Z�P�w��e���K�u�t�v�!������b̛����%ݽsD��+,mn��x�F�s#f���R2�hj���XNl��/bڗ��$	W-8�:����C%����jӭ�e�Ȳ�ḧ́ɭ��Q	W��Fѓ&����Y&;�i8�d2�_e�6�b'�������18A:w	��S��nKw���kl:;.����v݋�m�����u3M6�^2*ˬ@O��$5��2#Q[ڼZ;X��[`��0��Phv��wl�5�ah;�[�2�-��a�V	����`ۙY��hG����bdKT��]�0�6�B����Gĩ��ЌU̕�U���Sn��2���h�s��Ƅ�ӏFQ�*�/cww�lU�-��F�œ��RavYʕ�+3b�f�*��qm�%���M5�:��s5��M�b�YƊ˧�B�'dF���'h�3ue�B#W�]�(өI1Y&݇�!���cN�Jd�e�I0%�Y0m��pkܸ�QS��[vT��	{vf]%��ݯ��y)�r�Sf��[�.Wy5�QS-����0�ᖾri����ԄB1�m�r�Mx��-"��I���V�M��Cs/V�a�R���F���t�jY��jT��`�6��9[��@uR� 7.b$�#��{U,Y���7e7�0���{C7J�6���R��jMV�vҚ�Óz�j)�L�;N�ɹ�.fϯT-�8��KB�*R�dX�1�����n�̱yB�^:wq��ĭ�(�5p��`�����Y��y�b���w������ne���Il����Y/3ܢ1���+�wR��1U���&��jc3iڽx���5�^=�U���ї% 6�qhA���@�j�Q�շ�D�㦂��Wʒ�,-א�J�4�%鷑[�h�BsN%YEؗ4��㨳dfn��:2��@�FЖ�j��\�˽im�RLGU#���N�cs2���^�&�ͧ�4�	u��f��[��+�H6fl��Im;��U�/.k��,Ն����!�0謱l����(jt£u�(�3;ݬ{�'ow謅%�X`=y�to.݊����`;ys!IEY��Ys�NV�Aľr��)B��ւ	\R���i�ו���/U��2����&n��kf��Ѥl�j�a� =ז_�o1V:��xud�ɻ P|Y�N�b�n-����+
!��`�a�{�u*��;�J��f�E�8&�2[wgbz�^Z*=lL1��ͬ�w�
EQ����ڑn�͊�,AM;��b�X]-�+�i˵�K��XRc6�lԹ�2n4�+�7��6ݛ[5--�����~S�6��4��RM˺*č��ѠCc+a��7�ʌ\-�Š�,�r�0*�w��u�E&VoJ֛biiIu
�S��-O�Q<
�`[����H�Z�?��T.܅ͽ�l|�3����<��Ц��e�J�ǈ L�;-ؤ���ٺ���k���90d�Ԯ�.!D�ژM\����[���I 2J�L� ���kh�h[�^��ɬ��p�g6�n��y㙟b�*��B�Oj�Ex]Ϯ����B���L�a'��43FډT�����eY�Z>����T���f�U�M�d��A�Y+A�t�
�3�T�V#�zX<�Qrm��U����6�L��X ���0w)'v�X�R�Ez�M������Mj����TZ�4������T�j<Z��P�#�Z�hI�\��BT(���̭6]6R-h���{
���F���٦A�l9��� �ٙZ�EK��.�ū)���]�0V6� �������nD���aKv��u �5�g-T�nc���e�SТ�	��wt3$�v$^�1�c����CZ?
dۘ����z��n�����W2��0P+s`6M(�tF�N�
ӹN��7kM�����QJ������
������	���f�i��)��=ߕM�r�^*�Z+6�;�b�{Y�H>Kg [o.�:X�n��{�%`��m�#�֔� �&�e���ۥ�r�yf_�SJu�������"�ܱ�l���t�ѹ[&�B�*چX��)X �����3U'C%�]é� Kwba!D�6Yrfue��Xs�x��v��kX"�V�g6n��-gS�j8o&��$�niMl7�]�F�nĚ7C�x���y`
�+٧��黤3H6,P���<�_��Z�2�&-֧�}���QwV��yzs �R�6fe̢Y�!�v�ެ���z5 S]�}����ĉ|ɸ�̔4��3(�;a��Ĕۄ;����K�5�B�h+^�Mȅ��/�����t�]�Yv�P�W 2Qܤu��у+hf�#�Q�Z�V��4�ek8�f��5��b�l���Iff�oB��'y��1�N�����"5a-�y��m+w���b���4]n�9�kB���1�vۣ�j��[�	�ɝ����mܠ�)%��V��N����w���s!	��&U*#����iJ�m��i��:���	F�,��ܬ���*L�����Z+f�n�`�b�혋� ��\��[��yRkz2����u�W]�յy�PY�`��6���%����1�H�vUeỻmi:0�yFD*�/IXC@�i�,�*�bA�ɬiz/�֬_�`��l�6��٪cF��Onڻ��Ma�b�#%7y�p:bn#Va�2ؔv�e:�FK��f�eBoR�Ď=
�n]�P��ݴ��h�;m�MyjT�vN�g4216K������B�4fY���j�`�Q�&��6�ܰ��h)���`Ea�+-�A�*8o2JV�5��*%w
��F[�u);G&�*����A�+Q�uG9��tl��E�`��!I��H3RfZͻ�Q[���B�!9}����d���4�����O�0S��X>ZQ��Zװa�YLTt0+
�XG�e���'�,��5W�й�b��*�[t56�*y3o,^�ϳtT�#E^���/v�h�7aڨ�ۧ��n!�q-z���͟`���y#FV�b*�|�`��U�f�m� 
�d�7�o
�)愝Bl�cL�T�0%���8���˃)�\h�	�M,v�42];&��Zf��FT�ԍ�b�L����q���6�O4����6M��F[��	�a��gC��P��t^D`Ym&3p��K2��d�r$1]=�]�+�9.�7���d�{�i��lж���2DxF�kXP�]��[����������W��y��u��N���|�￫��C�@�H[[Em���X��mX�V-j��U��bŋkhյmF���6صQ��ckEZ֋m�X���U�Ej��5E��ŭF��V5kX���ըڪ5�m�5h�QV�mEc[��ƶ����ֱV���Q�[+Z6ֱ�m��lh��*�����U�mj�m�-mX�����TmQm�V�X��m[�V����[cU�[F�Qcm�m�*�QZ���b�5�ŭ��h��kj6ֱm�-Z��5���ر�Q��*�mZ*�F�m�'�I!!�$$ I7~��/�y�]����kjnǕ�y�j�ӳyBĹ�{j�m&�wAJ�?-��&ū�v́���/)�ٕy���K���-z�]�жM������ł�Z��f;�Ӝ�n���<I�Jӌ��3��2��X.�˗���nj�mn���B)�
�[';Q��;z�̺n5'�y��}3�W}����-KG����i��:���b��n�t9Ҝ]��ΝѸ��y�#�q0�e'[t���4ƣ�p�5��A�����vtm�س���ou;��pC5���z.�y��Q�����ŚS,i������j���葢�ˣrPz^�ou�C^�^�c�Wb������9�w�*�m�ܼ�i��]d/fՅ�{�Q��κc��
<���鹴t�S�z`�6��!{Ĭg%͙w|��yբu�!�(�'���]����^u:o�����7���*�K�ws�n�'���wk��(;�`�v=�N]�����h_m��i����e¹	u!��啀�wwty��l�|V[Z�
P
�㢠ŢX�����������O^�+��uiy:�Xv�]�X(�V%�i阕�g<͏��J�����:�����B#E^�[n�l�p� ���9>ѩ��	�p4��x��v�L��5S��1!�S��{�e�5}gw+�^\�w�8�]�BƟ��6/'r��uLgm�N�����4�Jl�u�z��/n\�^u�(ӾN�so���#M�t������iW�A��T�8�О޶�̮҃�2uk�����uu��>c�9ɮ�[ʀ��[+,�V�WM.�i��94�f�uny���[B���Oe���݁QDSh<�F��g*}��՘�Z��K��w׻�hn_^f<�/�DP��;���o�w��X�Nz�:�هgm!��I�1�>se󛒁G�7�3�yB�8���cN�Ct�r)i*e	ʋܹ�ST��K�wET��Ϻs�K�����"V� 8�7��_g2Q˃��#s2��wy�	 TvŪ)��ٗ���YX��f�O@r��͔�)�X׮Ŧ2��5:�7�pt�[�IJ`��]��;�,�k�e	����Z�.����ݡ�5Z�u�����V�ZQ�*���T�n��hX�������;�꒍_+wM]a+�7|�
��b�c�r���W�lv�iP�+�X9��ӂ�kx���o���tK+"ؾ�f�F�U��+1�V�]h�I;�*�����Y���G4���w5��Utu���o���ڛ�=o��u.��:�<t���2LI��`̽��Xy�'�v��َ�]+���r�苦SC���n��O:�6�r箑"��ÂcK5u�B�ړU�Y��k�z�/�{�(�<�tc�HK#HN�S�cw`mgS��a��㷃;�nҭ���!@м�+���y�m�i{��<m 6���)Y�okyU�i��,�;�{\+�S�
O���:�	,��xղ��Xϊnm�Zn��e�ǆS`R�/�{n+]�X6�I{37�*Y�/7���,��Y��G89�Vlw�9�OZ.�ѩ��X�rLyF��
�C>X<��z�.���@m�A��Q����;���AΣ�D���-��hG���}��)��xQ����t��Kd,��,1��`Nm��9k.�]�2�]�:���Q�Q/'��I,n;<¬D	Y��@]d9��Q�yM0q�i٥�Pj[�H`҃���9ʊ�N�H�G@�e����VA�+��.��H���Y��%ż���zYq��탓��ݛ�>̾��l,��4J���1ї4�3	g�(���%G4D�ŵ�)�;���Y-�0��v���oK��̤����c�b�7�l����/q��$r�]!�t8�H5��L'��u4�5�O_��Ju�b�&j�z��{*��;ߝ�Qӊcf���AfW/��[��ނC��E�כB��Vy��D{�F+��[ʃ��n�h����^�̝�K!�qWwS � i�z�u�����]�pM�Tv��^�A�e�hOb2��bܽjr�%�*�yv)ي��y��@o���[j	�h�V�_hE��Co��*2n��I=�Z�yr��M�xj,{�4^�:zs�Sӛ��xQoM��MY,y`���ly?<�or���v�_���/�֢ͫ�b)�D����guӽS���-�c�sS4�Y��n�����������ğ�or�L֜5�"�*��]y���<�ĳ���j��e`�������dA}�r7��;�*� ����%����"�	���%�j��vP�#���b�
��fQ�����w)BE	/w	ͺ�qw[�Pcv;��}�f���F�S��J��/9G�0��Sb����k�Yg�l;w��s��6y潸�k��+ەf<؈�XS�3kR�Ԛ��J�s8d��:����UM����A�B�C
���ՠ��<�a���h�G��!���5�0߶S��2d ��ۼ	!SQB#YV�`�T�����C�����l�U!)�Q����Z����}p�V�a޼�u�!8�k[�l5]��t��Սإ�+E��ͭՕ.���8����U"��G���[�V�8�d	�j�Ԉ
X�>ʽ�ݳ,A�w3:;O�3�ͮĲ���D�bY��_=Ԑ7y9�Ӥ���o;���wV3���r8:ַ�6�tu�^wi�$xR6��%X���j,���m�ұf\νٔMv1�l�k���ٲ*�V񣙸��V�yK	D�LC��[� ���&X7��!���j^\�+H#P[ϳ`(��mQ��b
�n��5��]�1@}mnI��ל�� �`�>��p9Iۯ&�L1��+��vSk�V݇G�f�㒖��ښ07�Jz�c���Z�z���@��)J.�e�������מ%\�/���!�*7�~��z	<�ʲ��\��]n�VN�t�&[�{;ep�-�QL��=Jc6�XUۗJݧGVf}z���C�k��2�ozJ�;��f��̉%���tƅ��}h���Y�0n��5��v���[�;��0_�����ހEY�y��Bmqٳ$r�.�f4ɭ���e>�u�frs��K71���E*�d�L��m�k4m����jq}�� J40�����ĵ���y�v+|p��e�f��o%��gW.�ˬ	��gN#/I3[8p�=^$��S��\��f��%�����zҳ�t��ě9[�-�m2��L����H;��:�˿��ǥ�1��`9��/E��HD��<��j^Q%^{���Iu^�U�����h�;*��xD�G[���zLy�X�
Y^�om��p��3(�{�����%=��ۈu��V.�5ݶ�B��|�PJ;�:7��⻷F�0Vmufi#.`1�����`�:Z�M��u��0����	�	{�AY��V��zB�{2��s%Y`L�ma7; {����.+{1u�-~��xD/r^�S+��1�X�g���5mS�M���--�2���Y1u��������U�}/*���1a,C{�:����1�:�;+2Nl�z�L���#:�U�AYB00��oT�������R�!��)8//?V�Z��
[���a/����4��w�WC�a�p�a�=�:,m�Z�D�v�PeJ{�����ɇw��2�8ݓX�ހ��/B�����yۻu3h�̼F��3��;�&�\���y�V�����4-��(e�|5á5� >�r�����Y���'[���n����r�ȵf�+�����#2�fpz!"<E�`畣�1�0�	���j0s��y����B͍Sn�Br��٬.iPӛ]��).=�Iv��5S1P�ۥ\dS&Ν���)�d��N=6^�=�hT���M_;���F�1�v�VY�l��7)u��� �{�Θ�|N�b��n�U��j(�R��=�j��2���h���p�X�ތ���0f@	���x��3l��
�k��ܧ/��1\��,�k�U�Ź��ɹv,�wLNwKWY��a�h�S�5
0���z�,�Xݔk���,fX�����<bkfT�y��"�g�u���0ЬT�噴p.y�0�<�箉[�u�Pc�)
��Unͽ�a������7V��6(�&��'�{�{�`P�D� ���,��V��TeăB�i$�ź�퇂�/e�L�u�2��67������dSg-F� ��Z�r�]�ݙ+uE��O�킶�R�J�R�Ӥܢ�U�
w{�g]���
 �x��KN�
�p�n�lV�H��+���`Uo[�v�HY��(9lj����k�f�ڸ�Qo.f��źǵ�hy����S����3��gmi:J�o�
���G%J�e��,�xf��ݙ�,n��f%�Xo�7yx�,ܻ��v��gF���[�p��X6�eC��È��!fY]Vt���륥�M/�H�r�z^j�Vo�ku���6����5��fSZ�g;�6�)ˌwh�b�'|J�û&�� ��:/��F��7�! �n�+.�n���.�l$�;fe{I�C�X��z������r抬28[�v*֪{���Zز�ⅅq����W5���͕�ʥ�̚(�mn���C}�yyKZ�%��l��g�z_$���21=Y��T���47h���6�Σp�tR�H���o�a �vB�/+j�<�Nw}w�zj�y�ۙ�zfX4E'ձ�5�c�JVT�؏s�+k��wW�eJ��:e�7wLR�}J�w���y[��:Nv�Pc�Z�����5F[2Ŝ�%6#ܲ��n�M��.�3��ײ��{�7E�V�b�H�T��
�����@��{R��0��M7�X�����@ɵd�Rps�'#��[�V�����4l�Lj}H��yy|�8{6�ve:�O�6�jiA�}�����G��G�Z�YH��V�Y��P��DV!���F'�k	r4���� �Ve�$ŷ��FJ����KzG
��
�PA* ;�iM�����R�3�;�HfǨ��O��}��i�b�,�u��	�����G>eZ����ګ����R�X���1>ޓ7�^�o��9�PaG��m�5�����j�06���rM��;S:m��ɂ�=	��so����zm�ZzOq�Vv��J�/K��������I�$46��N�8�x�EQfb�7b�X�~����[T�:�x���ؕa�6�zm�Ni8<��4Y�hpynY:���g��.V��ۭ� �I��N\����I�0�����d�n\��]W��*E�e�E��=�NPk�.[b�̝*jCKj�n%t^"�.���2o7�ua�)�(��;S�Q�H��;0�.�1�h]��h��+U�5�j7«5fq�� ء���|NJ�ak*
i�V�goXq��VK�t�9���`�Քw*���TJ��F�ƀ�j�o%mB��ka�w:<�{�*"h��5�E8y��0�G�f�C��闂�����]�VI��Y�N��ٻ�=�w�I:Q5�m�X��eEu�f����ҳ�)o��UӇ�*�U��f�ﻍ���$�?^*Y3�xKըv;��ͳ츥Mk���]�m��:=l�84���|4P�N�@��� v�SFB�5�����FD4	1�`x�/D���s�ܰ0h�����Ĩ��@]vmޗ�m��ͫC9� o9]����l���b��k(Y\,�{����)	]��f��l�j���B�l����Z��.��V�[���˥�����C`������6��r������{;��θ�}��>��+7���̊�Ik��x�H�&�������/Ҏ�L��ŲDv\�p��:��L������	�D1���:�Ƒx�'z����w:6�������c�L�U��]�[��X���9�`��7��bU�%h�姆��v�ܣt�@s�Y������fV�Si�4ފcI�%rF���(T熻�[�LmmfY��`b٭�8��xs#Ko6t.����Ǉ�pɯ����϶1MX@��uX�x�y ���S��a^e�|�oTm�������v�Z�������4'3���\ô�V�yn[Ǔ	B�X��Pȃ��m�I���{H�U[ڰ�l� �v��?��p}��]{/�X���JoM	[�Rue�̒�!a��2z��q�������C�z�rI{҅�:�ޅR�øUج���c��J�� �⬫q�v�@��T#f�[w�t��L�^��I��������e%^��;.����E��?�{.�љZ�7���`�%�v�_n��]z��������	�o�M�$�[��C.�����#�vl�DrI$*�I}�
�=��-��Y0�z-]���m'R���#	^�Y�o'
���<K�#F��hjDUp�⋮��y�jR9��	�oG�]�i���W���l��95P���y^�ƞ��%ig�fLMT^�K7AP^#e ��IU�Z����tm���m���Guw�j=���:d�(���w����s�;z�En�X�����5n��e�ˊp�0�a�؞�v�_���*� ���k��e9w���(>�TR��ZmR#[}�`�:�t�'+6	 ���,��d�z��2U�ب�X�cd�c��zM髂Kqҳr�����崵��餛�^![�v���~���ܨY��%�5��VV"kw.w$@h�oj����Lԅ��Tp�Vr�D��ң�L|�ur?V�x8m䴊>T�%34���כ������蝴��b�ρ�^L�Ǫkf}æӚ:�Q[֫u��DueX���o*önE6;��VȪt�N�Y���SٝsD�)�:#��jx-�����Փ��kv�g�%ZY������vN_����I��t�I���j�C:�e��sfsi-�Fjf`Qqo�w��g��l��i����iL項Xq��D�4�@.jܞ5���[�6�*���4'�Bz�V�ma�Vkx.H[!Hᮊ���U�F�-�D#���T���4&,��4�؛Jl�Y��"���k6I���j���1i�ˁ-w]��]i(Ӂ�\�Иuif.�l��"i��v7kXl6��M�X�kU�ֹ����S"%Y\��S\�d�n��+��L&�u�fԉ�q�v`�L�[+a*�f�f*hm���ڬD]6�ϗo.&�Y����2�6����* ��I�Ԭj�Fj���������F;P,T�eԳR��nK*O�<�J9��C	f���VfW]����� �mA�փ�u�.đ7jR�]X�f��ͱe\�J�uEsk��V)�s
���;X�LKm�\�+)B8v��ٕy2��c��+@��B��י��Mhd�� �@4e��e�TXZK� is5a˭t[�Ktf����1�Xm� ��7�뱌�n�iPB)r�m,�h��[N5�!L��TMn�QKNғE���.�)V�-[n��c�6��2]oYa��J0��3u�l��y/]
�0&tc3��`�8����T�)k(�ֵ����E�����YZf͡�X��Ћ�m�.���L1a����Z��k]r����L�fB�Rf렛R!+n�Y��[���KuՄ�eb�˙�pv�5�5�ME�˝z�\*�i�z���rg�󆬬5o�ťV�f�]������&k��L�Ii�˳cFQ&�I������av�����hjF�6�6P�f�{`�ث��)5.ʮ�0�1�Q�'K�`Y�n�+b�K�y ۶Л2�1X�WUlL�X.�����!5n��طF�)6�T��V�67K@,t86x�k�UWi�{X�6�Wi�Ķe&qJ��[SmsE͘���M`�3ԍ�wZ-i���I�b8%�H�eL��u�2�3WX�bgQ+rթ뚺.�#4�Xe֌n�sD��AvI�Y�m�VYu�=�6�j���ƍ��,ic� ������3�n��Y���T���,m��2�;����ѩ�1��Lݔ{L�MjVV��ʴ���Z&��YH�1�����!L۴D1P��2�`�C�^�kcu��#�Ck��Y�J#��&��6�k����X�*\Ș�[+{1�wf�\���hK�f��k�6uw1c�e��B����Gi^��[���V�]ڭI
�a���V�<�B8��f�[�5Jk1pB�L�ݡ�u$��Lʊ���6 ��Z�U��JF��4{\�{CGqMPڜ�ae�P�l���f��mK� Bx.�5
�D�1s�M�V�Ju ���2����+6�/��u�hk5r�/�������|�ĖTv1f|c�,|�X�[%�,�e���^n�����bl)0ѥ��*a�[2h��d���tI���&�-��81Z��]LKV�ʅ�aX�n(�*���X�0��Bݭ�1`�Z�LFYi4���6�t,+2�+���.�.�I/*R�z��vm��5Y3�Wkr��� �e��<� ����̢�]�K�:�Q�I��G���3�L�ٌ�1N���k�t�,SV��u#`�&��ˡ�,�@.]&au���5z�W�]�,���(Z�X5���c���\q64�[�3K���xy���K�M.)�1�7SLLÀ�0���B$E�	��%��B��R�fPJi��I�qT7�&��1۶��f^VK�8%Gc�`�mכI\�GFS�����̈́
RP��k+
�D���f�@����-�-�:V�[>ȹY�4s�m:`4+r,x�̷D�M#n�.�.�+sX5Eb��4�6�F���*���Ь��l#H����̸��a����g��gih+Pᦼ�6���uJK�*�#lѹ��4�.�cK�V�x��u��@l�548P��^b�.�\M=i�|���[�ד7V:��U�n�fɆ,����HR��������Zj�Eܺ���mK�f(��&�RƁsd"�%��W8�-@�R�8&ѹ\X̧Y�&	�1`����lҔ�yԥRh�E*�2*=�R�f�h��6-�+s5v��ۉE�s-nu%Km,Y]J�9AK����-��ұ6��\i��HY�#��Ļ]+e̴Y��l,�SSZ����u`�r与�K��n���6;����v]��-΍���X�ݝn1*9�x�X���m�)k��b�9�l���B�L�ؑV�U\�	,&�V�]v�Z݇`�e�z��4� B�a�pr��,�tX�E��ku�XU#,v�UlS5ҙ��V�,��YZK�"�%����h�P@A��`贻Xn�mk*�D�@��K�F�]�cZ�u�eɷ-�
�]ۦm�-�J�JL�*��7T� ݋U+F�
:ˎh�l*���Vfۭ���Q���B�a���[�#�,`�7mjB�&�l4��$�����)iu��+� �]�b�J��5���Q��ʭ,mcm,kSm*��1��ub��i�����U��XW����Bum�;32�nJ�e�*hV]Ib3�3̡,)\���&"l��7&���8�0l�sM�2q���2��g��E5����� �e#6"h L�ѼQp��WXFjX6�T�fR-�Wf衪��ݡ�q�Fj�Tl�tr��t�m�j�l�cB�bĚ4n��MQ��J�!B_Q�q/m�آ]
��`�۞�8mTr�+pn+�ID�d������宍Nu������FWGUq�%���k+]K׋Wf�m)�a�y�u˖��E�k�X�2�u�my��V���ݵٶd�	B�F��ל�lâ�813Ju�5l�"B�YIXء����٧��5-�e��m�Ŏ�4�ڮHf���"�.A��aux�n�}kt*��@0�B��&5X	2MHi��]���`X�k��v��]�M�]e�R�e�n��b�-K��mh���#��Е�p��5&�r]��k���`���#B.:�\2�	k��`���W0���270�-f09��)�����m
Y�6a-� ���8��Mk���!Iv���cnM�eց�.��
���V:Ŷ�X����!iZ�4F�Z�L��p�l�::^��R�#0�Shm�H�����m�X��j�FŽe&5�����CB"�X��5ʘD��ۥ��l���Pb9�� ��ڹr���F�;D�#���4-�`\�j�R�v-h��Jw�X�1�9�xA�s)�q��]�䄭�!�!�!��������hظ�.�e�ˑ��%c��q\��e��3%WZ1����V-�����[
L�Pw<:c�n�<�!,c�Չ\S�r���54���<b�!�ķg^�2\IfƆXB1-��8	Z��Y���K���-9�JrV��� .ʷB���,�*�1s���XZ,S=�c��ᙷg1Xk-��;Z#3��J�9�&GZ��!	��B尥�H�b�«n�4H���7��d!U5�%{R�6Y��H�� R�+��Y����q�����.�i^%Bb%5I[@B!�f��&�:�B�a�����TU��*W9�-�]ԣ�!{;icV���l�gD��:Y�.Xtj�V�����(M�Y���X�Y�Ch%��볥��A���u)���.����`؜��n^������x���:ՈeF�iP�(���@�-h��lؗ�R	1�h��cK��ݙx���qm�stJ���!����l�JR\�g,�kRьBb��T9XXֹ��f��,&����c�C�(�Զ��%"�f+h�vKe�al{����L&�)�b^�KtH��1̡nF����k5!��Y`�3Y��fú��k,kP v��SM���!��$ʚ��xƵ���&.�����e���G�F�f�l4mr�U����"Ü[P� U����Y�t����n�`e�A�����9���V=
�I60C�\�:� ��5��!�k�n��MMji����D�P:k�7涗 �Ij��5�k����Ձ@��S[3�w;Q�uu�潒	G���WRd�5�5��Cm���K�Mwj��l0�*�t,�b�5f��LrS2b�l��v�ґkY�xc�ee���*���@��M)e�`Mh�n4�VY,M�Z��X�dh8G�SW5�#ak��
�h^����ثEf���\���ltk\�:�-��v;uv�%�����	�-��k
���LT�Y�be-��<�YlE�����f��B��!���Gg���i�Ɩ����Y�-��\T����3jJd���֖L�4�̽`�b´{L��й����s���p�e�ۗeܲ�D�fJ[X]�m��my�貑Yt"�GEȚm��GBM
���2��Z����is �m��)�4���\ɮ׭�rR�e���Ch��tV�k
\$в���&��8�Yj��)E4�KeΪ�m2"-�0�c��j�G��c��`�e�#z�.¶R,]�6y�uVBÛ��ڗ�+�h�l	VqX�A����haJ�[m�JQ�mu�[B�t:�Xᱤ��4�Ť]h�5iX5�Y���un�5��ڑ�R�ѻ+5�F
MJ�4�e�5�Za]L˂��0FCK
�F����\ґQm�Se�e�
�T�f�jE��s���j�<�����ǷcbR�b�d[�et��Yl��.q,�hFث-��ZZ��,��9�K�X���4&�f��0\b�������6�s��T� ����l���:[4�1l�u�ˮ�e�W\F�Y�#A,,W�SM�ڵv���n��e!���h�Ұ����U��l��E�sa(�����itV+�f-�E
յ� �e�3���i�2�@[k��)�m�]�CM+2\�d!�,5h�e�j�@�rP&u���me�n69Q\�UȪ��XՕ�}�7��� �%"!�l)4��R�l����@(h�i��jP��q$1b0B	��L�����L��d1dL��E�\.�fLI�6BJ�F������)���h�X�e"X�3�����(��	�ɠ�D��4hM�RF6���d��ILcwh  ���iwnAI�T�0��!XM�#b�M4l��IATc%�Bh65%E�f4E(F�I�Q�,��h�ƍ��sQh#H�Q�ѣX��1�llc&#d�H�Y5��F�	Ih�cPh�4hLlF�Ew]��Q� *-��&*t�Iy|��J�����3Duq���ݵ��D��t:ԅ]j�Q�Y�.8Iqm.�dV�Z\G����-c
����qtR��6 ��`�	�v�͙]S�׶�(Z
�e�%�`�a{h�*D�����pe3�9�-G�
hT���:�m�����5d�T)�YKt����R���8mع�l��et�X]�a���j+��R�ad�gK�5m���\�@`L�Q�M,cGV���#��e��+`@ss��9�ZЍK&�lѰ�V�h�`8v1�<0&��-KYP[�k�Rf�/m�F�2���-����f{J�4!M�L�D����k0Ҁ���amXh)F�J�b`�BiB �-[��.#{c��he,��M5�ףCAm�)���K*�����j�f�j�͝@c*��e��!�.��k{�v��Xk����PSA%��K�M6�=�^VeѮe\����l��l�h�岱����.uw9Ƃ�;�dT�u����.�e�����f�,+�7[�Mԍ.�g�m��U"�l�\���޼-�[��,U�:�"�2j)��0����h8��L�a��ufi�Tq+
�J�����d���yLf,�A�(��� �gV�M�T��n��9��̝�>�L�h�rJ�ke�S�,.�0%�U �X�y�Y��!2����{A����jfh�-u���SL!jͥV��6�I[k.Ѥ\��"U��e�"�p��LU�#��G���SHR11�M�F�$ֵ�\����ķ�-c���8R�c�fy�Wlz�hi�[
�j��u�4�TA����m��)�urb:������YT�YK�ƅ�s0&�Qcs!I������J�����ׂQ�*[x���ijK��\�V�r���@�WRR��U�f�`Ai6U�[tUP����D3-0l%��Ghb���auB�4���$��ŋREKb5�J[m��a�V�e��S�`Ң��aJB-��i`�k!���
�60�W�T��RYe�Tj��+���qBF��mb�i��z�E���`BV�h� 0��ʤ�/-�b�  ��P�cVVū��1���,,Z׬T����H���?[�_����kB7&�P;fSb�d�A!V9�[�4�<f�)XWb�1�@-���_�HN���h��;��h�Y�@�Ы��=�`�R�An�!�b�-�[��z�sv�"D3�T٦��jt������j�b��҃��v�"� ��3�@���_6�Yn��CƇ�PM���O�)��S�B^���V!��R��w�/�m�����n��b�k�, �ҷ�_�@��|A���������ywױF�S��=��5�~/X�]�^�e  Πy�	n���Co�!Ԣ{�;�.��{s��6��m�|1��q֬\A|Ct��ַ�����a���z��2!Mt��Z�Ք�sb�K���MtZ�H�v�Z�k??Yz�_	�����HAn�{_9}�B[׭���ǖ�	�;'n���P����@��	m� �7Z�J�r>o�����J�t���q�UΈ*i��Kj�M|ߵs��+�/}07�jk�I�0�٦9�n�X4Emhz�Vת�O�ǛW��N�K������T)�@���n��[��tY"��O���Dͻ+�[��m���-����Բ�ꝩ��^�n��/�Ǐ�ڰ�A�(KmY�j�;||���W�F���r�2�Fn>[;��AGr
k�������4�������"Y����mYg���od�n]�����v�ێ�V���!�b�t��9����%�:M0B��!^���A+Z[�iU��HA��h%�	-�)fET}G|��d��:�"v/�A|��������a~><��ږ=���[�1wn� ��}Ǐ������	e��vj��ǡ�_n!�2���3�n>Sz�
�kr
k��m A����m��Ġ����}����r���e�A��T��>l�î{wV���!�P]�4ܖ�r�#i���߯s�B=�g������u�[������z����X�_��D���c�Ao|�e��[�`�~m|h#�{�K0ӫ��/��F�7A�s%���g?/>���A=�F�;_k"�@}��X7A��-��n�ï���T��E��ַ��P��[�S]`�m A�_ Cm}m��T3����g�B��\��+i8�kf[)�j�ю���jif5����G&��'��|��"��A���a.�ri��c�T��d��ގm�	�~�$��О(�k����@��՞�D���g��=�b�?H��L���9��<�~���F���ź�(��z��G���؁�|�m�e�D�_`3��ɔ4{�u2���7���2MnAQ!��Hw�������ź�����L{��/�w ���[i����U�9ly���*i�|*�١_�\Ovzϭ���C�],�{�L�D;�$��n�_^�]�U����6E�T����l��yG�aw���7�4�a�3^�N_ Cm-�����afz��c��B{��e��e���{mg��5^��}lA�A���N�0N�Ju�����4,�p4R�
���.uN
����h���#+P�ҿ���n���O>��ϗ ����]:J�B&� ��X�D\�.�t�S �Ȏ�_���@�AAm��|�R�f:Ɇ�4ܠ�&8�6.vGw[��~��[�u�ȃ��b�n��Q~��R��\_ G�.������6���h<����鯟��ݳ�z���5�~� �ѫ ��|�KmY��=j�WM=��{����ެ ���|g�>�:���ɺ�
.�O���Er�>�aQ��_�F<��u�-�@KmY6���A��j8�Ԙ<e�^�~�����?ly�-��u�#[B�t�6��"��M`���o�:IZ�R�t��˽7x�6~׻Eޙx�%i�F�4r��н.��G�Z�]!Kj�Yƌ�y���x�yc�5���BР���mU̳TXԚn����P��f�Fi�d���H_綞�����:,z猥��(ܺ�Mx�p���7��1:�RZ1�M��e�-��a.J� �\�$�1��u�[���L��sj�	���a�5,�*	��;FQ��Un��b�6�3{;�Pױ���K�,��5�"ٮ�M�m6��(L1��t{Sc��fl�-owϟi��B!����a���q�MTژ�`�ͱQL�ݛqY�"�UF��_�+�+�|Cn���#��SMͼ�˾o��w���9w��_X|���?6Ղ_/���x=�=��Mz��2���_+���t�/B���(�ו���o���-ڠ0b_c��;�X ����A�i���\�z�7~{뭧$w�� ��@���A[�e�@��m|�!�v+Q�/��m߲����3]����A�$��5g<���?z��{��FYP��[�|�W�C��� �{��Ch|�-��CnŖ�^�ǖ�W~�|���ӧ1z7�E�X'�K�k�m��[C�����}���PGƯ뿕ՃT-].�Jff6��6��)h�lA�c,Kx�v̮��OV| ��d�t-�a�=��ת�H�G���C�7��7_2��|Am|y`�[���ܧ�+(lS#!��c�����ҽ۫�st�pU��8��A��s�A4�yp�)�KH�v��n͖sf`����Xkn���#���h#��Y[6��_{^����M\ lA��-ߊ�2����x쯐 �݋-����&=���,W+��b��<r�iG5�!����E��5W��-��׫W���ź�m_͎�f��n�H�G���[���T߯�=�q�K�A�_"w���"m|i{{���5��/���[6�^_^ů�C�?w5`����|[j�Ugk4�X|�|%59Z�B6\F�0��&V�u��SP[� -��uk��35��}�|9�/��t���$�_Y�+�z0��c����{��'+�
�����qٟ��ý���j[���G��Q�xz�{(�cs��{/eg8��x���Au�n��3�{�D��}�J���H������m�D1����G��e|�͚�-���ĩ�h
�����2��敥��¶�=��ѡr��k��)oR�,��>liØg�4��;i+�����{SX�WA�j�. �i�Ci	���uwy~-��B�����|[�{[o>���'9ԇ�E}v]^P�,�^�CF����@����� �RBv>�
��W��u6?^�Z�^��{�	�"�݋��7Mz�qJ;��C *�"�)n5���@���d*�7B�B]liB�.5�h�2�f�KSl���d��!����_��ٵ�Oz��`������ʋ��d	�Ⱦbjΐ�_7���m�^��=�霧BB�<i\S������<���X?m�C�kqՈ�vbs~��yY��j���׀ ������v�.�����~�d{�'C�#Amز� %�ۿ�uwt�\m����u0Am|����_{�o&��܌� ���d7�ƻ�x5��Vdț��=���ɮZ����ŏs�X����}�o	�KH��EKJ
�{��އWQ�>�&�����4�Kcۻ�b4;��A A;9_�6�?��m����_w���8ǫW�L�X���y�7�%��>�@�9����_�My����ߚgM*$�T����	n���&Q�i����pUz�5���֔g�g��v���(/�t �ڶ�>~����� �!|W�=rؕ�}�j���z��)m|h`��������)|��˿�M*g&��:���(�l���z+��n�\��E��}�Q�5#H�|�m�e�D��a��qX^:{�{����z7�d��"8�!�b�-���{��OYJ��.W����"���j�N�߶�99~��AN@���^�nk�w[��6׶H7㎑Cm-� �[��!�Zڗ@�׿�*ULΜK�*zf��}(Y����}A|Ct�����W����ڛ���g{��U�o�&�4�;����S`w�f氰2;:F�o�q��ȇ��Y3el���){���e�� ����(Xi�l�C�\R�u�9�#�*�Ի"���^#Y��3
��msMJ�ViVf�hll�e*"Tenck(¶�2
T�qfE�se�� �MHA�X�v�"!u#v�Q�0�W[�bQל��1l��	[������]1�x�7V�T0Ue��V����Dv�K`-q����S*Zc!��2��m:�q�Z�bWy'߿>�/�Z#�kQGl��rhb-�&) ���(s`�3[k�y=AnX�[���V֎�����o�-.���׻*�9	������=����D7H�[j�"��ዄ�}o1�E� '�E�/yng{%9~o|���1�_�B�u~^�q	�{�"=%�Ө�ۿ��H��z�zUu������A��	��d>��n����
��fQ�d���8��!`��~n���v�h\׏dk��/��U�ݬum�wc���1��!�@�mY�Ե`�pxyW�ib�=�Vwi{ŝ�n_�� �	�"5�,� ~n������ZNa��S[KJ�CJX�*jE:�&�]	e�c.�IX�e�3��R�,��b���~r�6�����@e>s�{��pS|�W&�w,����<� � ��H��_7�Ct���>�4T���J��U��ٻ���F��i
V��}�G��7I]��I �L�U�{h���J�S��ΦK���1c^ׂ朘�"�G)L����s��hOk{�
K���"	ޠ���m袎dX�A AȬCh Cu�-����m&�:�/+fU�u��o|��8�� ��ز� A����V܆�W��,�Ԁ?fP@�}`_�6�Sd�l��qSm�>� ��VE����z�dM�A:+6��h_ź;Uz�,��h���W�c���Й�f�]���"	ޠ�m���mZ��d��2-٢��_Z�*�Mj�ƹC]A�&V	)c1�eR�z�f�*fo'�~C��VAq�!�@���Sq�|�޽��j�B���˶��P��BoX���_]2!������������q�}br՜��PشWM����';U�_ �e���v��^绶��|��Ծ��D݋-� �d?�aԈ���C�k)Go�������k�`����n�R!(\�QU�"��/�gJ�a�܄��oK&�-�N��Ѭ������0Pӛ p��c��׬yT�ݦk{�d�}��v-B��`An\U2��>�����kZ��sc��Wƻ��7&'&	�:�g�/qi8kvs�L٠VIf�����8G<5]؄p��T_�|��ƪ�W^gK�KLŶ��[�<QLȧ�ŉ$�VF���]i`��c�p���uշ�i��)�=�bX���+\�e�o0V�؄7Wk�,����f�sL���f�������A��.�h|2�]B��![o+�Y��vL���Y��y�� ��omm���Yެ�:�N��w-����#z=[���7Y�[eu��:�Z��1����+;"7e:��qr��ͣz��a�}Y����|z��7*\v3��
��WBV%�Y��ƯFv;��t�PG��Տ�-P�hu]�Fa�Q0|�d_[ԑ\�R��^{Km	ml0���"�jXT7�n�޼ݺ����ŋ$��f�)8j�⬏���W[M�%v�#y��
Ș���_��9���WZ����\�͛�vn=z\#�79z�ظY����Cv.]�M��7<q#T+����0�G#0	W}�_;/��>������O�˼뮬�nfQ��x�)`��e�v����1֜�5�R�m���c��$<��g�6P@5h��ԥvۈ�2�̕�ڸkn��pe�>z^�yYxz��ۭyX�cYڸ�ނ�|�]�}���(��b0XIe&�4i�F�L��R��%������&F�&�jLl[D kh��1F�h�a��4$TX,BA-���4�+RQ��6�(ɢ�T[I6�+EEj�sh�b�QF�i0[`�J4��5�DF�-�QA��h(7.U�4Z47u�J���lQ�Fƍ��Q��lh���F�����L�b��|H$���Q�ly�&d�\�X'%|���Cn���ͯ�g��=�=w@׫+�-��,���WM���qM�9���
w�����t�xJ�r�A�!v/���B��ط�����Q?gͪ_q���&�J�~�;�a����c�|��P�\nN���_};���>���,A!�5V���+��uU��K�4��&�+H�3�m]y��z�{�-������n�I�*Z�d���*��W��:�����k�����A-�`��o<�*w��a�0e~��Sp������e�~AN� @8����,�^ۏ��	�Ɛr/�yb�2R��k�����͡ݛU��������[f�Jl����}A� A��ՀCk��J�3�,纾�s���|_'Y���8�6|�s\�X t�# ��x������u7�M��V]Ʋ�q]V��e�!"曠(uM��K�y>0�B�=}�l*���=��S˜�F�ۂ��GG`_��h"�|k> ��n�+��*��uh��V�t�z�y���A8 ����ۨ wiF��D��n<��왌�>�@��B�V@t�]k[[[�`�qq!`X$7hA&L�k�;�ǽ~���v������Ñɺ���n�Jl�A[�Xt"X�%����� �[k��Ct��W]������δ<?*���d��R>�9�
��-����w�c��~�d�_dA��֬�_7C��ڒ^�۷���V{f�M���
p@��_"�b�n���6�X���Vqq �P�@r/�8����I��ǡ]���~��`�������Ư���CH'5� ���_/�m�`�L.^���ϵ��B�����d�S�s6}$�\W�-�#�|�m��Ch%lf�f� ��u�1<9	A�
����q`�h�V�u��Q�`���^��{A	t�U�j�E醛�·T��a�{�k�y/�MG[Ύ��n�EJ�����m.9���JU ذ��,��M*��m#i��[�d%�v��t�Y�Hh1��ml��j���:Ĺ�eum�h��m��f��ð����M)�t-!0���i�m�#+��C�ɛ��5ve�33+/S0�pGJj��#hLf�XR[�(g�b�3�3��&��T�b���͙�L�������.{&�� �,�ɝ��B��k�QVn�4O�'��>��ADn�E��Sp�Rc�'fIm�)�!c|���~2�>��Aז,)|Cu�!�b���H��P�^����}d_m��� Θ��^�
����P�=����-��p����ei�Da��dv�J�n�n���ȉu�<2�~�JtQ�z��c����_!"�6��-��n�7Gֱ�gG����=��P��V>���y=�c��B� Aݯ�N[2�/����}�Cn��Kt�n�D6�6<#+�L�]��ɏ���U�����VGu[�m����<�]�o$���o��7m�"�)��^�f���x��IAe��,F�f�5����e��Ùg�/������f�����������U}b�
�.�/�3*��T������_7C��VG9y�R�z]�o;�B�Qy{�d�+��S��z�4����knIO�^l��m,T����-�lgff�k�}�{Cc8��9)6;x�}���̠������U���L����;�_ #[���S�>�<���k����� A����_[k�f�|�����X�^�[���~=���;�E���VCh�����d僇�}`������!��}��ܫ�w?P��5�Q��$+�D<w^�<z����_^�-���__ͯ��M�ꂌng��_�V<���y�ys�F�����|��Yn�!��r��O�5��՘.�M�
�a��
5XcQ�ͣ�M	����4$��ܩ!f���`����/��6������٠�}n�q����J2j�A��:�"-�d6�@����b~P���+|��(d?!�iS�s��s�l���Uk���A.P@���)�f��q�W��|� �?� �֓}	xG3�q��A�f��UiC�y��)ו�;��/���y�9a����L:��-�2���[˙��b��d^�  o{F�<�<��#~�B���#6�����̷@6��x#J�t���@@9��c����73+s!5��l]��;U�4ӱ2�����H����@��A��b�-ҵO}�����PBE�U�)��n9�_X �G�( Cn���� ��?!R|���qò0q��wV�0�	��:ku���u�ȍ(0(ީ֨uz+��1��ze���KmX�"�'��27��\��㾥�3�8F�X�u���� ��`����\z�OS����y{7���Y��{������ � �!��؁Xph��r��~,�$(�����$���H,�2Sʅ��%$)�H�~�u��o�Rp�߿;���Ξ'?w3����AK��|��%2�s�@�RA`>��A`hi �fX7D��C2����Xe�?%$,���_9�M��m5����II��T- ���s�MFR@H�"�� ����}����e��27��ﴐXo��
B�U�n��$m6��޾*��]���3I�5Ҽh���p��!<Vڂ(�Jǧ�P ����p'�ae.�y����윷�q�e��)��������	~����ùP���X}v�X) �fXlCi��)�eB�4��XVf� �4�AL̰;�Z���U�.��0��XVT- �e~��Ϲ�_�p{s+���vϠ�I
�)>�l!�%$}��I&���v�R
����L��g�?z����������5�(,t��=�Gb3e�M��4mT�.����Yldq�Gl��t��'� ��P�� ��S�����͌��2�hi%$)�f]�?s]�sZ����No���}$�݇�m �}������+��Ka�ꅤ��u�i��I;��7� ��3*H)�@��v�FJH(RJL̰4�R=�}�y���~��
N�s�l�I�R{>�������垹������~�>�=�Β
A`?�v�R
AMs4�
Aa�P�9�����a<�P�a\��Aa��S���6�Y)�ùP�	I�R�5i������`l�RB�$���ɵ�sA0��;��d��j��?UW��5�l�2RAB�R}�l!���XT>�ᤂ�Q
`9�l�e$
JL̰4�R�:H)
��{���������`RAJ>��i�����ZRAB�Ve�@����m�\��w�d����|		Z�Ci��Sv�hJH,k���{����m$�r��肐Z=�$�0˶hd���S3,!�%$�p�AI�
`9�l��j���j��i �RRk7`i���s����oY�W�~������Xo�GI �ݻH.��
Q����͌��2�hhII
�+1!_PW��sr�៍ğߤ[3^<�읯.���yO)� h��πc�)�L���"o�Z�f$��{�I}�������+9��՛�� �8O���7IJf$G7vKn��R�GJ��jL���f��"�������k���Uf�m2�,-f����VgK�%G�)0�"ˤ-�F�5H��j<L��x�;L˜JV�pոkA��jF1V�B0a�f+��]3U��P��i[���
�%��!�A�S+��71�7)�!Sn�3q/T�6^n, K��ƳW0J�R��\̻ͤ~���^[H���SjGee����V�C��	�1��DV�k���4��z}$޽`i ��P��) �*��ZA`hH)���肐ZW���/��s�wox��+ 8�Yvϙ) �]�ww�_^�}0�O��H~RAa\��I ���d�2�
D���L�$�H)U@s.������G>�ߵ�k\�n��62S��hhR@H~ܑ~��Kӯ���1�
]���Ci���Ý�ZAH,O_�I������`s:�����H)��uP�AM Suۤ��P�II��HlII�Lˆ�
MS+.�4�H(�� ��Q�Ko���]�G3ը\ۼ�˼�~��������I!ETݻR
AH)���i�)�eB�В�2�H,4) �fXlCi����9�oo�ϵ�����ܨZ�JH,
��ҐXi �}�����]��P�AOVk;�������v��<���Y�d���	)>�,!�%$�g]}�e���;u��$�B�˵�L���S����cI�e�������jAu�R�3@m �c%0̨Z�v�5}�\'�
FޭH,;���������[�~���AK�XH)��T-蔐X=�iH,$��I �3*H)����k�����}�?�@�/�a�l4��F�l���+wRjۣ�&^G�Ҁ�Z��Xf��I-���/qgE
Rw��H)��޸i �Ѕ03.�M2�
	I������������_���v����Xo�H)���Ο~��yZ�y�@��jAq�I+���Af�%0��CBJH(Ta��R0����a��JL3*����X�W���}w5��խZ���}�<�ͧ�VN*�������U�p��..�e�nh��t�7����?ޞ��Y��
�j�f��/U��5Z�v�u���9����AOX�RQ�������g������۾k�y]��y�Yv�ᒒ
$���4�R}P����S2�d�j�ۯ����o���H)>���F���I!UP>��H) ��fh�ld��H)0�թ��v���kϷU�y�3/y������?w�}$�Ձ�����a��- ��{ZRM$��f肐Z�fT4�SH�̻Y�JH(|}��^��q9������
��H)5�}v�i��� 
"�� ����?j^�yW��G^ߴ�Xo�����U@�۵ �������s�^Ă�FJa�����P��3V�aI32�bH)�eB�
A`k3ZRM$���v��g����
A`W_G�������v糲��zS��?Yv��JH)>�,!���X{ꅤ�B��k&�I��3,02�Y_~�f��>�Z5W.�ZS �����7f���4�k�5��tE�~'@�A�t�R*�{�jAtF$�����Af�)�eB�В�
�KD��?ߩ�����+�y��$����Ad��~埓��]�-�I�G��) ��e��� �̨ZAH,˵��JH(P��3,!�%$��׿g�����AI��0;��ɦRA@�(��� Y��}��׺�U�y�׽�G��ߪ�RP?v�H.��R��4�
Aa�P�7�?�g�LH(la��Ԃ�Q�$���hm �P�a�T- ��f����S3,n�)�3*H(�����o��$O���0謆m��ն�\�x�{H]@ǹ�J�Y�L)+4l~w2�����Q�Ң����xjG
��V������ʝ"�wfO{���w��`V]��) �I)>����RAa^�ᤂ�B�̻Y4�H(���`i����:H)��<s|�
�ڐR
AM����6�L;ꅤ���fj�����^�����G�s�È�-Z �AH,9ʅ�}�5���;#�)�֒
{����
Aiʆ�
i��k4�I �fXCi) ��2ᤂ�PB��k'??��|h�i �q)3\�4��߻���u�g+w������Aa�P|:H)���jAt����w٠6�Y�Ja�P�4$���0�թ��v��ax_��G��f�"�uV�]&e�kcl��dY�KFĆ-G,2i`��qlUf��$��XH,���r�h�I�Y�����S3,n�)� I_#�H����}ٝ�~�;� �e�ϙ) �^�>�c���I����Hr$��ùP���X}v�~����@���`i ��t�R*�f]���
{٫��ϗ� �AH,=ꅡ�%$��O�?��N��w�R����~�qE�@~Ci���ý�Z���������H)��O�gR}��o�AH/bz����)����i��
AL�!�%$�p�AH,˵���H(���`i�_{ǵLv��?a����f�r��W�����I!UP9۵ �`RAJ;�h�n2Sʅ����fjԂ�L) �fXlCi��}7���7U�s��h����T-�RA`Q�֔��R
w=`p7D�Їr�G��cߧ�5s��}^�;� ��Y�%$��}�Hm%$�s��<j���Qp�0e�zj��O��s���M^m�� u�3w`�c��Yu�W0_���ha�ox��h���1��\4�`����Bɵ{`9v��~w�����=��~H)��v������}�I �̨ZAHp���v�Q�I32��Af�Ja�P�7�ܷ���g3�����]����������|���g��>��
j�a�H)�{P�RA`g�Ԃ���AL̰7� ���$ޒߎW������{���0?[lL�@��-�!��4�R˦.%��6 Ga�Қ���͌:?�O��~V���bJM����6$��»높
MD)��v�i��P))32��{�뻿os����������A�� �/G;����{�m�2�]��$�߳@m �q��g��R
a��I��
H)���
Aa�P�%$���W~�>^�9|� �:�AOgl��
Ai��i ��}�?sU���s���g;����.���I
��}���II�}P���B��˦N����_��vq �~JO�����H,;������W�I��
Vfh�m��fT-	) �3.Ԃ�1�����^�^�۟��M��?|8����X|!���C)�v�h��פ����AL̰7� ��H)� S2�����P�9Y�?�����XC"JH,(3.H)4!L�[&�I �fX`l����z��ǟ����}I����� �*U@�j��$�n�g�^�w���[�� ��*��%$)�ei ����a�6�Y*2�fT- �eZA`~H)����������p��^}���
k�s����}�������<�˫g̔�P�%'�e��6����i&�)��V�R
���偦��5_~K��m�����'ޡC�ײ�0Y1�p�Otj<�e�v�e���z�M�?\��m�#3kn�1.�I�S:◚�Q�Z-ye�/J�c��Jڴ�2�fn�;��y����fXE�)�쭼������;��`tLE9݇F!ڲ>%��3UJUjf�P���[1�(������Cz�15����]�zx#��T8¢ķz���{��p�����/�MN����)x��ۄ侱�P�@tU:8�.]��&]��Q������ޝƳ~�z��|�LK1�wu&���#*Į�,2lcJ�Z�g�Y&yd�r�:R��b�E�n��MM�EQ�We��*	�Lш]�Q��x�X�N���q-jmw|�q�[h@�G���M�,�5��'	eT,�.غ�X��V�7=�*��ͱ�\���ّ�����{��M�:��"�7Ny�>̫�Pά���,K 񥷢��a����1��湎�ձ�v�Xl�]+T��$p��v]ݞ��9!���-�Q@��Oفu�/0݇�gv����6�����F�ѽ{V�ye��C�#/:v�=���R�_9m���}w��s���Cyȥ4nX���	�%m�5���X�d�D�ı��*j:�ʝ�Z�o8���C
�Шl:�ՄJ���������ɔCQ�ιG;���d���b�a)	LZ�Z+�_�|k�
�Äe���Q��Q�DJ�gxF��U���7�]a��J��F�n+wj͙4�go{m�8Q[����u�sw��8S$�*�	lD�b1XƴE�*6��5�ۆ0FѱEb���6��F�j�cb���JƊ�m��%\�h�T�Lh4b1F���4F�BV�hؠ�6-QQmr�%&�Q�1��ԕE�+
*4nsDjH��h��ب�I���Q�MC6Ʊ��!�7+�I�EId���Є����^��
��F��4��mtp«3k�����J�����W�[6e4R�B.c-�l�#{B"]�c�����\M�"���Ŗ,m��|aI���i�4]R�lز�p�uk+��,�PJKZ�7FV�+6�+��5f��<KiK�q�bm�����l�wXT�5Z\JC:��L�eE,"��{cj���Q���i�1�l��X�՗M.5I��<Jrٲ�Q���JҴ�f��˲�]�o.�2D��l̶ˤxv�mM��K�rK�`	��Y�J��v���b�ҹLlU��6 �B<�]��m�K�Hzn�Tf,�Mu�D7iPa���P��3���BӒ9���ib�8-�3L�ݝԚ2�=z�CCs�4n;6�	F1���hg[vϪ�_ yb�\�c.!B`ғ[�Z!��F�,��7,�l6�̦ZK��GP�
icc(�[���(g<r�9��	[e��]u�K�F�3�`U�lP�����w��֨2��U63�V����X�b�ر��;62�%�8��ats,![-�f��tSVĹ��h	��ד6+(R�L�&Kۅv��;D���@����ɸ�F6[vqQ� s4�����^m�Hƌ���v6�X�,�lڑ�Qdt��"m��/8�k����a6��%qm��WJf1�lF��dSTλ��!����Gvctff(�	J�eNś�Z1�
��;����5���,ڄ���|5%�y��
J��!�+i�]�T�+�l�obTl��Վ+1Z�K��3A Me41w`ƙ��%�%b!&u��!�ɌMGA+��4V�K����b_"����S���`��1@s�2m�p�mL&M�ˢ�atF^n,�Z���F[��t)5�5�a]2
��c.u�%U��/0���4��)��G<Z��;��IMP�FɬU�6�f��M4ښ�NK�n�Q�X=u�רךW$��������L�L�Ipƪ��Ũ�iN�e2MV�ԥRf��Ɇ*�JmM��L��Eg�N�;����o�m���YcM �����n�B`��hY��Rǭ$s`�$aK�S���u4[@����T��M��KtS���Shk���5����^2(���z�"Ė��L��X	lX�vh@v�[��h �Ҕ��Qw,ة�n���[UT��27)�t����%n%J�*�\)�g2�YK]�#�āX�:�k�j�C*h�	s[j��O�o�2ڕ��:���m�h�4tP�$	��]��KnԱ�k�.��h�
Aa������Xv� �`RAJ��h�n2Sʅ��>�>�����m�#7:�Ⲝy�;��5z���L�7Ϸ���U_|a�La��-�I�G2��Xi �������]��P�AM�̫H)D���`i���¶��~�^�ύ�G�}$��)��U�i��R
}�07=�������}����������AH,�� ���;ߴ�62Sʅ��c\���~��'�0�V�
AH)�zÐCi��L3*��) �+2��XH)���肐Z;��b��*d�C�)i2ٌ��d���9�|���|�I �����RAaY��I&�)��Vɡ��P))32��m$�H)��=G7�j�~}���V�^�$�������Ja�T- �40����?o|�G�o~7�#�G���|	z����ùP�A) �0��������7�$F�
}���肐Xg��SH�̫f�) �BJL̰4�Ĕ�XVe�I&�)��Vɟ}Η~��w�I�I߲����ߥ����7���RAa~��t�RU�V�]F$�������Ja�P�4��
�2��X}��߽���+e��Ue�:խ:hX�̬;JM .�	ͬ�����;k�a�cM_�>��O;�����Q�ßT-II�A�^�
AH)��I �̨YC����=���	�����~�Ғ
�ߺ��ݽ{Ĵ���H)���ZAIȅ0=괂�P4	I���i �̠�$�P3*���I/A��������~�u�o#�.�����C?;�~�9�`9L����gd���B�^%�&`�7H���y�n���n��#}���� �����w���̔��ZII
;�Y~����&���$^�`i �|�aܨZ�������M$������Y�]���R�=�����)��U����JNfXCbJH,(̸i �e['�RA@�)32������ϯ_�r�~9�;����ԐX_��RJ�ʴ��`RAJ��4�7Ja�P�4��
F����Q�$���m �v�k?sO|�̝aܨZAH,{�����I9��7� ���$���y�k]�~�5�����y�۫g̔�P�%'��I �����;���ַ�yH):�03�l�����II����cI�e�$�Tʴ��R
fe����2Sʅ����_w��mU_��ACl5��Aa����__Ͻ߯�3����H)�j��6�Y(e0�T- ���zH,$��I �̨i ������]{�]_Vޚ�B��Tl�)�v��1i4wh\��G��Z1�z�Z�j��n��d���	)39`i �>��I&�)��V�R
AL̰4���߾����~9_��{��H,/�:H)�����T�:�`_���`RAJ߽�6�Y�Ja�P�4��2� ��
H)��Ci��L3*�R��?t~ϝs��߷��ߒ
AH)��XH	t��W���,L�y��ٛw�H��`eդ���)=�XCi) ���p�AI�B��l�o�����k���>���A@��׽`i�����i!���ZAt�������4�̨Iq�e gK9���oX~����X�T��vS���շ^�	Hw�`l	z�ᆘ�7�{<3r��3;	����9�AJ.٪���.4�m�������f��}UU��Q��qA��&���5���]݇�";D�,!l'{�L ��� �h60��go���c��e]Uk ��a8��p�����A�{p}�~�V���~���/?|�P|0���PKN_3����n�oޯ�d�R���~�/�C�H�[4��gXTy�=�mzf��#�<��Jݠ7vW8��͜8�%|fQ�_#J�*�M#*�e��6Ս�0�@�A�%�*[�a��ٮ�~땚���C3�m���/�'��uU���Ywҽ��:��H�C�n�׻������������;�@l�7l�`���uu���)���a��ԑInE����{5˿'얽]�p{�賍d�9h:%ߒ˩n�q�L���������}��}��]�s���\�q�+	���mo!]&�r���w�T᳡��Nb�A�j����Ma����y�2b���$��ǁ��2ؒeo���}���W�����i��I����!�JUY���s�y�{��oo�w���b�Ԍ�1�﷛�2����.�J�%H�X.am�6�"�%b`%�ĩko.�`���I���y'�G|�y��v���s�ݵ�k�����i5�Ǘ;#�L�3wwwE`D���'{��8{�ng�~��~&�����Z�n�׈�~μ�?W�����%�����c��]w�7��].�{}��!��tU��]n�+����{�}@Nk��x彻j�m�;��j�5(d&���ݼ�O�!��"�mm��cw_<�D���{�{˵�M�]��}YM2I9c{@	Y�9;n����n��ݘF:�y�~ۯ%��*Y�����c��bO��i���n�F�ҵVq��M������ꪭ�K��B���*0ʁX��%45�+��f�eXE5�@:�5lH,�a�`d/gY����k���ŀ/(B���Ŭ����h�p����KF���5	h�i�[kl0�!�!����#)�[,����y5�ԙh �V;B���#��1�Ͷ�!u�:�b�5�sS���++r��8�ص���R���崕C���{@[a����֩�us���߆���ƚ�555��pŲ���6���J�-��٥J"���t�,?�.�|3�v����M���vKw1N��Me3�N�/�s�}<jCRE!��R�׋�@�����e�W3mp���I�%n��E�tv��z��5$��Rk9m�{�u+�/v��-�]7uv�}�C4ԑ}!��/_�������+�}�w|���S���-��;���Ck��Q��߷�<d��5!�?@��ׯtuP��'�ӹ��|&��&��e�$>��^]��]WF�Ih�h]X��Zv��Mi,���46�����4�pAZ*ϻ��^���~��h|7knl����mM5UFy������P�n��CU!����a�i*�3���o$��Yx�����;i�Ej	�-շM\E����!��J1�MQ��!�v��U�%��_V��&���� �/f6/�����i�r��b��d?v�%C�F��[���j�?IM��;�U���)}y��d���b�en�ۺ��ˊ���8x�tmk���.uGbkn���6����i���UL{��}!�R@�{:{-(��O�V�0���$��\�ͯ�=���ߞU��ɰ�
}��g�-�%�gѮl�bحͅ�A54/&!lm���[�-�&ͥWD�l������L���T��]m��0>i���g��{/�7c���Hk���ee�Zs���n�Ӝ^�ꉘ��4�w����܄u�Z��Y����CROr[�c9y�]�[�+�Z�G.�FKԷYpξ82��vc�x-<�[E]d=6���i�`\��m��U#'�����F٥������E}ߎw7�}���lR�9"�ZL=�F��f��7���fy���s�p�4>y�l˛3,����n������NJ�x�2>q��;��Gt�	>��5SL�DmO*�<v���hr+���ٱ��.�U%&$C&�ʭ��2*Rg�ac�(�6v��6�����}�%�RLr���o��;���_����r�E�d2E!��v׎v�����UO`���a�s�훸�ݝǦ�r�u|�����b�.�ķܼ�q�5;��|A�S�l�Ԇ�5\�ax%����;���h|7u��9�U}�2Oze�6�{e~��"�PG�
ȓ>��D��G�kx���.��l�9��AI�u~b��{c,��xh�ᕚ�v]���ˁ��k�����gm�GYJ�~������]����*�ԆID^~�����1�ٕ�WIX��f�9���R�I�o�r��"	<���ںV���$[Cl���Ëc�Ԣ��aX�a�f���}��׹Τ5Rz;���øT��\m�Wv��j��Y���Ԇ�H����k�/�ƫ���L�ް���Y��c�}N�z/�C*�����w{j^�R�?Iۨ{���-��b��V��za���s_o����,ݧ'����V��J�o�[!�\!�5�r�p��lz��g�ԑT�D�^1��_���έ����o}՝��>󆧢�Ihѩo?23�Dh3]�Sowru\Gr��v,�_fm5*�m=�G���Wۻ-�o�v�n�@m���Y�A_�2'��y�dO� >���ܗߗ�X��!j��Ʒ����ch�C��Ҙԛ,��U�m-`��:���p�Rhj$p�:Z@CS[XT��[fє����0кf�i�`&kcV)h�6�][f��v8�S1#YAP��[5�n����%I�z�E���y[ͺ����)e�p&V8H�h�eeDZ� �+�ܸ�\,�Y[�l$q]lA�V�JĺY���0���Ś�Y~Ɓ�TL��ш]3Hʁ�T"�*\�+n��:�ث�B��+Մ�������"�G�=�VS{��a��ݼe/�ƫ$U!�G�//�m��bo5鯦��עqN���n�]���}����Z�u�{�}x~��I%��nRK������Q���o���������"�=<o#~�>�ow�۵��v>C�����l�扮:�ao�n���?�3"��*q���Wr�wW�&�f]�� ��uRM(U��~n��0i {�7@Z�2]�1��ٹ\�5S�B2�&�.iI�l3C-��ϒg��J�>��3F��֮ԜrOzg��8>���;u�>U��!�I����]��͙y"��}���ą��fnX ,}l>�`�e�L>m����ʌ���L��Ճ)׮-�&Vi�5�qMu�A�^�_�I ��ټ�2��睿7��]���4{���_oI�e��7/�q^��?IH~�'��7x�x�cRr\[��8et���O�M5RER�4���o���������%,���ھ��o���5׆D;��o��"��2�&�\�3{5���N-�=��YsC���7vzg�_���񫏈-�9A4���q�fI�CW�t.iqLKAT��+47tڬ9U���Hje�K�9v�pM�������_v���Hd�:�{=ݞ�x���"���w}�`�o��W��gI�x�ڹ�2����毪i��}&�Y�W�Y�3%��*���Gv0��y�[�4nd���o�.�OA�̻�*�^-s�w�ۺ2��
���^@�����[�����ne]]3�K��tL�	�"��#kY�ț���oV�C�����;��玓�]�H��x5����3�#���n��܎8���h#H���ھW���dꂆ�Y�L&^#��v�g3��Q�z2�Y�_+$`�ycY�U��ϝI�6ȶ�;�^k}�n�� �V"�^���Y��pI��]�&s��,��5�1}���#Nv8�z"�44��N����[��@QKt黬|yY�p(ȏsT�i��T	�OV�5��fUӷ�Q�V7���@�u��Wndj�U�4�%�%:F���i���qVR�v�旕�/ ֡K>�-�0�ٺ\Z*.��D�BJ��u�׷���wr��!�j��]����G��o��z�b�s�չ9m<��I��b=�� v/
ؑ���*�6P��Qަ^k+E�w~G�ś��nT�v%v�q^�i�dkp�`Zc��"���z�yU[L�α�0��I�dҴ7U�3����IYЁ������w�V��ݗ7�-4�5f��k���9�F�Q���^[��K��5�;�׷��(㕲�F��j�We,:(�G+.omĎ���+[5�u"יS��B���d&8UE�;f�wy�	ڙ��qT�Rή�o�]2�'}��W�o��*�&P�t�
&X�ڐ��]�~c~�[0]���7�0�S�B����jf,�(� � (���k��Z*#Qcb؋m��e�ű�Q���FƋE6��h���mQ����Y��F�E�$kEb�t��*+ʹcѪ�75�%b�h��ݭ�(��sV��ͫ����Z,kI�Qj�\�[QQ6��V��#k�ܭh�Ť�`Tb�,KI>�H�����b�毬��?.'7ln���X�;O�L��"}Cv��{��:�xCr7P��zPV��T�/>V����7kv�݋CY�)�����]Ws�K�����{k��*��z�f�u�=B�J��Ep4��[*6&\�����b�ԭ���{�p9n�2|7�mG[���ct�elw}g^�VX����7u��d�U�y�m	���{;�k��ނ\�����P��u��$�㓦l�j{���װ�=�T��?I.�U��;y���K�\T{�oc�s�8~��_H~��$_=ݿ;��Ԕ���~#���v���Sq����x'}./�;���������Z�~�2���k�HTW��:�N��;.�������w�
�/7Q~�����v8gPFX>�ӿ۫�B�5�L�,9��+���s�W������~s�N�6V8ڇ��{�]�_n��k��Ȼ�F�bG�*4^���X3,Mi�z4B�1ݚ�Rg\43���Gʾ��ԑdC���{���oN�s՗�)��p�����:*���T�x��z�q�gG�f/��BΩ�����-��W_-������ )�]�?OI�P�m��e��/���o���윷�>���jH��2q���^f��|n}�zu�2˷��v����s��lZ*J5����d��?T�Ou��&:��.���g����7�=��L�������ۻT1:�B��'�_wB`��=w��uҡ�����2xM�`[%�\��9��+�D���q��Q�{Dp�*���I�;��|��z*��x�@�Z��Xئ�F[�%���a���!Y,��f���s�:뮒ɓ��9���ʜ��ΈZ1��(��W!J��%q3��\ּ�	�2�*���X����A��WZdvZ����p���v*晳8��H�����Z���+*�G#JU6�KB�:W��O�ue��lJ-�7�ġe��&f볛4v3�q2�,He�$���%��WW��u��щ���e2�ejB��R��6Y�K���w�D���<��焥�3��}<�]�N�şP�<���YV��=��C!�"�U�]׋8��b|}ꩼ�Qk���]���{��fr�n���Fd��)�U�j�?IT��YO���kw�7zf�=S��r�h}��nС[w������۴v��o{�u���Ͼ�{5u�R�_�q}4Ԇ���C��|�A�ޫn�gf��Qk�ooJǷ�9�������}�a�r߄��TE�c�b9i.���v��I��u"�m4R�AlQ��뉐iYJ��i����x�$U!��{L�=Y:����]{��+c�E�j󞆤�mn��,$a[&��^��N��0W��t3��ˮ��r�U���q�5�*����wv��vrW��5x���|r��1��U�����  /8vW��Y~���O��56t�Ϫ��i�`s:Z{ۛƽ���C��"�xj�%6�v����/�s�者fs�ԒG�m��<��L��T��T��3oHYޭ�Y���2���o����k�ݑ�R�"��@q�5��u����}���Μ���<k�H��j^�ݏU˻�#R��\a��kh�eGF\]1u�����QWE�U(:�kY�]T�Ua�.�}��ޜ�z�7/�����5�~��UH{B�GX�Bqw]����+F���Nxy�<S��W۫e��C�E��c�{�����G��
����X��쾼�ޣ�+/+���m1D������N`}nU2�w�h�pOb9�y�_��P��!��8�j��v����J�)A�����ˎ��F�{�Cӧ,?��񯦙"��K�]�j���#X5�^�����㛵N;�����s�Ym�͗��;|�����$_H~�H�AxrV���3Z��w��S�\C�7o�݋P��Ԫ��Gh��e��U��mYe�q5�b��Հ�l�k�Y�*�S3��~���C�/�������sya~��F��{}k�?J��I���=Ѩʵ��v�{��2Q�T3�Sѝ��窲�9H7:1�u�|����麆�-�5ن;d�~�CM��gxw��S�\_9[����7k$��ܞ~��[�6V�|2����S�2�O\Y]�#z���Jk,}�hbKݚ���d9�"&�ar��i�y��u�񫬸']�{���
v�m�kv�����kN�j�ꯪ��w��ԇ金C����?kpw^�{^��ș���ѝ�}{�!���5%�ˢ�y�*���x4�����t+�,;KG`�d�(�n�-�Ė�
Ԕ&��H�f�ӕO���#����V��L��u��۰�tY��n�h}��n��oj�����z��P�C/�`>�s�di�˾�c���]T�!K�gP��_T��?T�E^��p�9�ߩ�����g�_-�}��O:GU$����oF�qY�Ȫ�5O�X{Q�s3�nY�}�ʮ�KO��\��ȷk�C��C6������k�n�l���9^��w���W`����7���=�4N��E�Xx�+����VS�[r�]S��u�n�eՊ��Ƿ�4V��^S^��X�����#	~�y���/�}J�$ך�V�hG�Qö5���]�B� ����
HZKk�jm��X�m#��貚�Y��Z�6��뜫u	�Σi�2��&1kD\�]���a-��Qt@�T���x6))Qh:	h�ݭ��
Kh�3�9b�X=��U��U���z�drX���s���`�l�Q5�W�u��Z/]���B�Z���e�Gvfs�ۢB������ݳM ��Qm+V�Z����4f�p�#uU7-r7��g�����ݭ�[�g�t�[�&�w�8#�jKy��>����T�W��{K+����Wݚ<|��`�V��S��	����.�Y�Mnl�"�~�N��7n�U_��m���#�#RT��9��wP�v��W�w�/�-'���#�1OW�����]/���4j�d�Q���H�CR$ ��Cݫ���[t��/����2�p���[�7ty��4ʧ*f�iZ�ԶP���!^[
B����DЖF�&-U,�Q���@�Z�uV��#Cv�ݠ/=����zJ��us���&o�7��N�����(9ʾ�Ԇ�I�Ȏ����n�{�إ6�fJy�7�zOU�eê��s$�*��b6��ta���9NM{L7N��<fۻď�>�M�����w����.��z��j�j��Q�=�O���Nw*��!�*�ݢ��}ä�Ϲq�p9�X�}~՜d?T�HiI�L뀔��S6x���]N=�����S��+�����}M�S���"��i�j�Ԟ�������o=��ﯥ򞪐���CR]��:�I���AW��jJ��7c&27S���f��,k��Y�\L[���k5[�#��5^j}��ų��`r�{ᓲ����mtfC��$��!7�̚��Z���^���8�}u�ڝ���O
��uŏs��~>�URIT���zEc��ݭ,���̛�q�WG�M��Y���iU�l�D�W:����=��oM��-�F-�=:ܻV)Vh��k�Xsx@�>���ǡ;罽�s_�~��4�UHj�?d��73=���z��zD�	�~k��^�K�նg����P� co����R}$��{�/�_�8HWt�.���V��ڹ���:��7my}g~�<���>�!�N�kcG2��	J�a΋M�l�x�9�ZB�6�ݠ,ݐ�1)F�O��/��ӆ�|�\���g�}���=�2Y3���H��CO�4O�Y����ʃ��~k�������,�����n��;��hL�.��z��v��^T��/:W<yAA&�N-u綧�1��!�i���*�#*��~�"�9M\l�s��d~��H��?.�����!)3S�LbI�Δ���swso����Vs���;ɀ�=�[�퇻L�Z`Ǚ�.�1�}ٟ���3}��o�$U!����ٲ���b�ܺ��<<���?j��!�$����m9�k��7�8�C\�[�]P8��P��ɪ�F����Zۦ�c�f�+�%@1����7k���AAݽ�Ů����9��e�3��=�#�Cv����>�����wjֵ�s������z��Rs��Y���t����O/����T�N~�#M�?r������q�X�U{5Vq��E!��)�b��T����7��!d�uSb��s�J�=��]����*���C$R'[v�n]�&��-�\����jOI��ݯ�"ݠ7`�w9lĽF��.�����hr,�SGzi[=������J���6�w.�а�����������˝���E���5˅d�/�3[�g�Ӫ��6-Ѕ�历z�t0�Ñ:���ʆ�R�;7{.7{hܤZ&�0�ۙ�4�1�j;y�ݮ�[\Ы��+�2ӕ{���;��b�׽������/���s�xQ�b���MA���A�%��r�/j�.NI���쾙��q�U����.+���S\]�a�׼�ٝe�b�m;t�C/P�3��{s�ޙ����F^b��1g�OJ�݆2������.5�syn�;5��%��ܷ��[��cp�A�f�uݏ��Y��z
���7��q*6s�MK'iI;Ga�H�B�؎2���<�s��1O^�%���:���ÂV��̏��|9$�v3h�����ϯ�J��a���T�Sҕ����S(J�ln
���2��>E�߲�y�Cu�z�;�$���G�O�f����x�ל������6�K��¤{��[�{�r��;��k��KfN�17ba���i�n�����I$��J��m⭔�&P��ga��uc+���mk=e�_(;G�;������y�Vƪ������':��m��?n�@X�1Q���813�Z��E�B,�{G��6��f����j
�u�hw=�K)Is��d��y��N�v3[;�KFН���]�{e+O8�q��y�Ud��NWF�F�؇�H��-�X���J�}�0�e�u��8��~镭�(� �@PXԦ���j����W-p�Ak�oO5�\�W����5�Z�nh��p�yU��[yo^�r5�ݫ�{�(�������W-��ͯ5o5F��w\���5�^V�nk��j��ę6��\�1\��6�-�%���\ۖ-]݊�o{��cW-ʣh�wZ���k¾z��f{W0\�)�R�ݘ@d6�]Am�� 8�2ݢ�5��u�����$��%!j�j�e��V�M43Ø�n�nu�ky(�f�\q�ֱ�CkPe�qβ��-�5���`��X+�3�6��*�l�5Xd"F��eChcUJ�����+[kmc��P,/WZi� ��K�s��)ɭ��̽�B�.��3�n��u��� ]��bX��ȅfM(���r�u�hd�bM�i�0+�]te�U ��5��E#W�d[A��A��<Ͷ�����Ɩ.�J�	�����3m0��ԤZ\�et0K3�c�-�:ۨm�hƚ�ʊͅ�XL�-��U��(껐���P�mض�s���k�j�&�b��-A�HPΔ�]�7�p�g$���Mc��ٓmf�� ����MoXYH�YlEǭ�)r��6�VQ-�L�iW�*�SeZFҷsX���I�pl�qin�8�F"�Û�.��È8�����HE���%�Is��J�Z�	��]�^������4��kT S�ְ[uɦ�zA�6�j��ؚ�-�s."qt��@�{R�\��
�Fh���Z[E����l)���6���Q(��h�mD����I�[Q�ZBܒ��ܴR��$������.GGD�EIfhʑ+s���a�sj��
¹�\ƹ�������6Ku@c�͉k���(e��,f�+�ԩ�f���Fm��cbV�Z2�[uCkH�%l�\�k�SZ�[V��f4obc������AK6��l�TiL��՗��Ė���F�JF�ˮ�t�l%����Ҡ�W�MSj:�\�X-��WG#H��*ʙ��5e.'�;��:��ւ�(�i���+*:�usK��f�. d��2����hQܷ$f�d0uҪ�j퉱6`)i�v6`^��뜶��V]0�ٌ�8ƕ%fr�CJ`�� ��p,�Іl��4�+�ڡ�H�w��l%�
V:g@Vգ*��;c�x<�(��VS����Z��E�`f�2i�b�F܋D��K-����U���+Il�&�S��.��DK���������k��jJ��X$\Q(�Z��S)��ɍ��n��������Fj[G\��D��c��+x�Y�k���J���L�Ū���zTxG���C��фHӍLke��۫�vbK�L1�n�6����Z���G���aI�GTn�`�����m��J�ch���d�o?Ο~y����>��j���㼱�Wq]5�~���I$uR�'��_�<���W�(_�B�ݦ�K���t:�wd�u۶D;S�a�9T��2DE��R�y��w.��sݩw>�s�!��#�I/�3��ˡ�_��7k�o����=/}ye��}=<�Չ�T���9��ݯ�u֡ePw/�e}������ڬ����5Y�I&Vz���y4�4I�RTn;@��F�)Z�K�kf��@t�5��Ms�4��gJ���|���!��&q�}��nnr\����6��)J������y��d�?�C[�-�{|�ð#<�fc��D�N�ԭ@�-e �
�RTʼ�Xj�n�w:�2�*\u�E�&G]wڷ�w��\�'q55��Fٵ؆��i���vvw����]L�w���~����ƾ+���TK�(8�Z�<k|~�H���:��c�RM����,_&K��L2y7�;�u�:�����yjTMn�4�vf-z�W�wP�(7�׽�����s9꘱���)����IH~��Q�u�W�񥏼!|֧��z�,O|�����=��f�1_�~�����}��9 �}��� �\���[u�i��Ħ��[#�ܚ\	�w���D���'������`�kتJ�jw!;��(%�����T�C$Y��e[{`_L�k�/� ܞ��{ڽ.I�\�o 7}�f�O-wj�uѯ��C$U"��LP�]*#�i����U�����G��1�����~\[��V�m�V�X��BW�)�G:�@�̣n�v�'[�(ҳ�?�S�F�O���;�����U�K��E%z|W�m=��i{>�^t{L��o��xѾ���d}�϶E_n��5������=�nɐ�'�v�����K�x�|7+��!�[��؊��U��2��b]f��*��%ҙ��&��ҵ҃�W1CQ���ne &ҵb�Ы*���~��*�=�e6�k����X�k��;=]�����T����޾^��sN;���m��룹��=�����W���X6�dux��K�MUR��*�I︿7�׹��/����W���$����P׉����u�NE��e+�᪺�ɨО�=�m���{��[CpLm?q�[�hNT�mI۽�x�Z�M
w}W6�5X�=�<oު۷���m��jp�P�|����w�v����׉��2�ӹ��$�O$�8d��ö�έ�@n�_��'_z��H�@����MXBel�,�͇����Ev*�Z,�f�Rۼ>I��O][����˅���o���$�������(n
ﳵ��CwW۵"���0�t�7�_N�Я,F�]����(l[��YY�<Fg�y���5^��H��ԐY�������ҙ��:�r�k����=$r�#t�7%�=9p��vf���[����w��,���_M5�?���!�2`D���́_�=B.�{}G{�s_dݱ��T�/��ﺹ:=�ѝ�zE��:�̹q5�ѭuu�<o=�Fmդ�u��\/C:���3:<Κ�y�pj�\Bo����8���ӻ�|�On�UĨG��.F��V"i�"Gu���Ŏ�#˶P�VB�l��MM�H���m�ͫ�X8��it�J6���d9E�Rm����R���0&����f"b��;���n0\�\!@ԍW]��d�1-ML�X�j�b�-(�躴[�[B��!�r9w�]=Ba���5�k�MalR�s\B���:���f�6���'������]�����fʘ\���U�-3�����77�[Y��������߯�<��q���ݦl^~S�sf�Y���gw=�?W�2?�5R���;���U������ևo\.gvcw�ל�o�~�����u�Y�A��Y��UY�I#�j��ی���׆h+�w.�yi�dg>��4�~�ջ�
�R{o�a�V��P��q��t�i����j�����ō�@z���I/lq)IaV��l����y6��w;`^�k�<�CR]A�ϯ������dje*}�	���Π�V��IM�Ƶiipe�+������N|�i��)�粮��Q�p.���Uߡ��ǲ�6~�d�C!ܲp����x�3�G�b��aa����ʊm��4&�J��Y�x"P������ܕ�U���PT���F���Z�]�w����h�~��Ͼ��F?:���!Z���jl^~S�h�ݞ��> �����_Hd?I/^�՚������r�7Wp�}�/k{��2D�[��u����F�&�7_d����E�X�
�K�����z�����t&r�C!���Lңn���9�o+3��B�nl^~S��Y����,�>�������&���9b��5�ֲ�(�G���ۦT�hh�*�X�tJ�m!���n���<$�_ck��1���8���ݭ�_��J���/-$���:f;����W�ħ��U9�U�dj���L�;!��?T�}!����G�Ы꺶�Ϫ�(�w�h�ӕdr���yE`�mO7'\��DW=UO
$9�_�o!t�<}��	z++�J?,�W�,����u���ξ��__����)���](��h�����|7u}#�%�����Rf�����e���'<R�~�i��G!���7����쉕Ӥ�y�隝*�����o/�J�v����5i�[�"	���(t��<B�`]5�Mr��`{[v�&��3*Y�Yc=}�k�_n��v�FgoXNx<�R߮w����AP��ձ����/�2���lh���Pp�{BdR9��]�i���y(��ӞRv�Y����3��k��jI#�� �M����н�!>z�}��8�$��Iz������T���?Ir�7���}/����WF���^[(�~Wҟ���bN��2E�`iL;�=���fn��p_�2u��͎dG���T��O�r�-�7��i*�����䞠���;��I.���T��w���M��aw,|u��ۢ�[�=���DiW��߾����&%1�c
�Ķ1��+f�LCW[��D�F�mH����	�{���z;��y���2-�{��\���C�S�;�r�3�W��?I>T*E�BB�S:�W���_?�H~]')f��V���z��5��m/�#��ݡ/���oTy�]}y>@���)*B�??c�Y&X�=H>�� �ړs`5� L�@�1���n��ݯ�4�V◖1c3�9-a�P�T�R�HUV�5<m��^����p׾��=�h�xFz�q��$����	ݯ��_ F�9w�I���>��Ah�ˊ�3�-�1�z�|?�� ��;�)|$7�M��I���5I��f�CM�+r�C�X��]�t3�-�	ʠ�;)k8e��]��5�uw��dh�M¬�WVnɮ�p��#��Th�BU��"�2�p�v-мs�� j�B)�&ܠM.�f9&���"V,�����1���m]F�i]���PJ͉�vt�ҍ�SJ�A�:l�JZ�(�	l"VZ.Bkn(k7X�F��7\�� �-n��K��9��4fYYR���Jh(��VQh͡�����]6]��0�TfI��M],/!t1-)�͚��2�z�3J�i`m���>�L2�3\�14����6������6!4�Į�3LQ'���~z9������Ϟ?H�B�c7%ܛ��!�7�7ƹ�^����?Vx��_Hi�B�|Ǫۏ6��FT��u��O}�/O5k8e^��� �_n�]��<b�#A�
�|�!�T��]ק�z���eL	OU�����.f�� ��� � �;�v���*o�y#��u�� ��z�u}9҅ƶ�nK�7��fR*�w�=��Tee{v�7�H�|&�_	*�P�!!�̌�����������}��vw�����'%|� ��#�K���Yr\-v+�̪���sj�46`ԥ�@���A	��k�G���l����� �vj�4	�H������7Pp�ܳ�T���lׅ��W�s�a(P��٦�
B��H�!�
r�Q(�ԥ����F�)x���2��{�W7t��@��{+��H�+-��
wo&Y97m����]>YAU�^�0Y��ɷ�B�:@y���ڕ$[nE�7��@��HF5���G�w���/���� �_R ���v�?n�V!C����v��o|TίU�86�9+�AƂ;��#u|��/�.�W�VU%��|�ȇ�/��ڱ��b�!��~��K�@�^��/uiv��60e�� F���|� �J:�`�w�������y��r-��"�����P�3WʅH�|$U�߾�i��z��J��#�:��+��	�h�Y
�iu�*mN�p9�E��=�e����zy�}!�����!�}������R������f����_�/��Fj�n����#����e���o�z~�4�'�n�.1{�=����@��j�Ђs���He�𮊩P��B�?HX�R/�X���y���鎯)u�b)M��n�?e�t���ߚz�jO��Vc�/r:�@��b�b��������VA�{V�	]4tI��䞼�\IJ�h-��ǹM���G�]�5���Ql�}nu��*�`U�Þ�����OJ��y7��>���x��d���]��:Zxt8eHN��xu��ٽ�Is5n�X�j��9�j�N����v�+۲F_^�˾��fNY̫r�1�m}��)b��j�s.)y�����.�z��ٽ\���H��74o^�y��k����n^���J,�̐e�o8�׹|3����� OJ`�xp)ڣ=�y[��e����#�z|�*g!�n�]���pY
 �Y�^d��{���K��e��*6E��M���
8(���&:�;om*�V鬣K�ʽ���ok$ioSΠ��t������xa]�wx���a����e6���[϶e������ջ%�J�iC&Q'<򓘱��/d��>�g��K�r��7PY���K¡�.f'v���]w��Ժ�_5]�ĕ\s�j�1�ԅ����;��Q3[���w���Rb�q�UK��5Q릳�TV�=��gg{8��~o�v�m�X�s���/���r�`���X�!�C&��Kj���������[��q{��Ҋx��[�ۆ����x���j��Sx���d�%\4خ."*�ݹ���5�%�����ӟˈ�]�k:�]AʏN^��#-��]2X��عvc7}C�%�W�/�3�N�nD���5��߻�Ѫ7[�m �N�E�[V*3�k���4F�k�R\��Q��kp�V�s�Z�kw[p���뛛sV76��Ur���*-͢����[��+�ڻ��*�W��F�v*�b�-�cr�ܫ�^nb��k��AW8h�+�T%d�جZ��G*���ל�rᤥ6"�nn�F����(	|I@Kmm6�7"�7r
�T��ؾB�T�*_	*�S焑��7�b�BCJ���<�g=����9��-�#�6�@�fy\�WL@_���bs�X��S����0l��g{e���m��b/t!ǳޠ8�_Gj�4�P]������"�P�*�U�!�4%ȵ�4.����άĺ��\�����i�+�@��|�( �|���Nv�M��q���3��|������鈞���#9 �#u� ��"F/PqMo�B����A A/�G��dy[���u�+� ~3kౠ���r��A��L_/�\J�	���ꑯ���d�=@�ޗw��vs�Z�J�_�p ��@����G��_��𩨼�өW�����vR�����)��뛹W NJDvZ�!I��n��5�!��t�]�)>�yI��:�}.�ԫ��i�˔7���,%�\�`s�e,���ږ%{Eу�m�'�Z����J�����$_Hkd�3�1������/7����6V�@���c���U�<��*�;7���,���l��+�K�3b\��g�v5��c6^� �M3,5YbT6*�p�4��!�T���焗c޺�9�c�����΄���ww��s��D�!�4�}!B�K����2�Ξ�6��z�j��7��r�_�-ɾ�w�_�V"N����1�����i�{Ֆ:�,eX�s�9�6"9^�]��7滏.��ly�����݇� Lu��4�HP�R/�
�*�
�E�]@���*����!�|�W�4n{�r��������}��*}ݷ����� F���ݯ���	�=�e4�T/����Wo��^�G:�5�~[�T���}�z��T�q���2M�i�^����+C[�n�ŁPC]�Ùô�^Ũe�,s�ӗ���{���YMҶ�Vf��5��}b�Mv�5���������'8$��J�m�%�F�'��_�lZ�Rhl�0�˥����f�v��ȳbW����R�S6�=M-P�eԌ��<GM m+5��Ρ2Ya�`kT��]�Y�7ڲ�E`.&:ծ���U@�c&T�V,��!�)s[U��0��+,,��L42l�1�v�sPz�&��!�.&��8���-/w��I�bS�2�B���--�5͠�k]�Z5�7RQ�P!�:��Q��'����6^�~��xH�����Fo�B��/ԩ�H��;����=�,v�9Si�Ycr�{�z3�z�_`�Ծ��&6=�n�������H�����+�u�ńߍ󺳃]�Nv�9R�'9e�9V#"��������c�u�����G:�� A�H^����v�;��6]�yd�����4��=�H�l�ޠ�ᕷ���Ա��~���s=��r�3�.'9B;��;��F�~���0��r�=���OÌ�s҇�m Aj���sts��u3^B1�*�'�IXV,P�3$c]t5�ƚQJ�0�]CL\���h�Yu�EYZU��)P�?�
�!!T(T���u=�z��7��Ӽ�1f�wXA���!�BCT�HW�*{ջ{�l&Nd��u0M�h�lo0k���
ACU�oq�[o�9muiA�H�7qճ�9��ك�	%���:'Y������bz/��(�ٮ�f^i���ov��	��@��}�^���@�tX�.'��v�9˖'9d��9f�[�@�.����,nن:^��|k�(�P�]�b���R*T��?J#�����u���A�_!1s�Ƀ�{�ɱ�`5�/���2woU�xN�r��D�T��HHi|(	
>�R�!��O0�v���T�i����}��C�� @�?!C5}!�Ⱦ}:E�l��8��*�G�����J֬�Ql�\6\$�ЛTr��#a[�u]ۘ�Ά��>����~��Þ��?�f�����*�I��P��k�ɬ;�3՟�3��e�U�9e��T�����uF�l�p#~���E�����6Ok�p.R��&��#v}�w�׻7we�ޢ���bs�[�Qq�������XH���XW��s_H2\Я�U�*j��Vj���i��)�:��W��>6�;��;���oz ��1˰���(mo/V�~�}�܇�c�� �h#�_!��@��İYo2�&��ڪ���D��� {Fn��=�0�by(q�H|=��c(�,��g��T���:�
���IU暷n�U	��^���񩾾�$s5�|����_!R�5�鎱K�=���U�S�����6n�bd�eۉ2�	P#H�+2Es\���i����B������X��9~��q7��3;|C�gVM�?O�j�ҨP�|��A|wi=��:J[��:�O�_�n/x��F�bq��A��� �A�
Y5�~ϼ��@�[H��n�u�B��/�-����ǚ�׷��_�H��� A��c_"7W�}�_n��7��ʅݽ��"�v���Y��{�togQ��p'�u�!^�#��X�Oj����7���P��-!T݊�-Nt��N�����w�'R�LcZ_5�v�T���'U�	͘�z��P����*$?/����6k�p�u7�V�^����^'� ��P���P���Z��N�V���z�nҡ Ɓ��䌲ׂ�Dw*GvM4�RW)����	�)%�$�B��K�r�B�P�HA�v=����\6G�X*��^̧�-�����x�/��7i|A;���4cB�GtPo�d��ޤlޣ��7����8�'L!q���`c�q�^J�~���P����ƅf%��Uvʣl߮�u����	/ҩ��-Ӆ��m|�4ӥ|A;��#u�r���A�}6��֐���o�1v�&�}�[���V�ʮ��D!�}�ӡ!!B�H��׷Sm������գ�yӨ70ʝ�"�Ӕ�׾��cA�HwW��Mq���ז92�]	7$�!]�3uo8�;׏�s\45�;ˬ�Ժ�b�Wƌ�PJe�ѽ�co�Ws@H7����k�{u������n�������+^	ڽf���ѳfuPx��Rޫ��@#
9��d�6^ح4w2�dD�	f�v�`;�YH2��6�Tj�M k�T�ٶ��R���ClF6j{	n���1�pg�$4�%�iKU ���mdֶV��f�1�\��U�	v�Y�$���^�s�B՚�zв��:���Шŗ�LZ��0w�-�~���e�>�v�GQ��R��V�6�6�����B靨P�3���� ��ȍ������75�^%���ކ�{D��BVZ�~l�0�СBC����r�6)7WCa_ ~־By\��m{���c�X;�[��k��w��Q���5_PG�)|A�E􆘡���V9�"��妳�.L[S��\�r��P�8���HH~���"_)B©�1;f|(l_/�n���EQ�A��'�Ox8sh7��;�A��WM���U�9v/9R�C���Cq���=~>��i}<oZ����q{�����H�_"7P_��Z"�=��b���2��i������h�4GLla����"�1 k�3��z�|��]wϺh{�b�@HVI�;2����G5e-���{Ļ����w��B����W��*E��B�������}/D���m�.����{���g;���=KVo"-��7V,�f�}o%�7����J!5���.�߸x�����՛k
�&�9E��?K/]��{�Ǽ�����=Y�K�kT>�!�P�R*T$*�	��+�[S�yK=�v����]��PF�?!R%�R�HiP��W��m�i��N��(	I�,�˕��!&j�zk�u�!��O�/��sO����w/��n��C�!B�H�T*M���!�t8�i��h,���c�Qo%񽯖4�CT��1��O��fi#B�th4���e*Ҷ�q�5���gvm&��0uE�,�3YH:4�z�Յ�;�K��<�X#7W���^�]aw��й��g<�}��|{��&��_!Sʗ�T$5K�!���oz�"ޯ	���K�@g��7�uL�}=ƴ[����A�Gv��1=ٮ�.�^��[4ǡT(H�B�K�"��[�s�ڑ�N�1Bw�clh�E1V�ʙqՌ�����2J��#������r���m��O۴>�d�����I0�ޭ�y�����l�\I3^�	�6$2��C�ה��~v���J#�߬5yo+���P�]��P�~����y鼰W?�2�f;�	�H0�;o�*r'2��,��(��h�X�PԠ�8k��S�TW;��L����i�5�� N����;������Eo���������y���Z�h�R��-��i��y�Վ���L�lO���/_��}y�7W�|F�o��{aL&��)��8W>��Nn��X��� ��A|_P�� ���� CK[�Տx$��r�k_MY}��V��{������ A�?=_�c��ށAD7��c�A�EK�!�BBV�����tx�>�ڶ�_Hi浢��u�@cA�_wW��7hq����7{�A��{���!�{yS�'CM�8���Fr��R���	�c<��H����sj�,��(�.������h��f��p���*�%jZ��[ŝ�ٛB�`�D�P�������j��*�"����"�$;|�7�S�Yk�K���=M�m��(w�� ��3W��R*_�TA��>�QLIE��r�T��9�H2��h�9�vc�V����V�G�.�j~'������e��2�����w�˝<ִ[�
����'��z��ߨ���h�����b<�Z_��齓�V���_ � w!��f��+���i�8m A��_n�op�Y�e	�
�R�;�ʅ	!!B���W�Ԇ`�-i��Ʃo�����g	yJ�P�_*"_Hi	*��r.S����)�:PFuA������[w[�:y�h~�:�%<�4m��W�*|Am|��A}�H�_/��{i	y~gO�&!7k]z��L&��by(p �m"�P@��D�Y�w[`h��e�[�������U۶E���{u�-җ�V|]�]G+qV-�:#�uI&��賄��;8omQF�4��'�l;P�<�4lt����+]ҷN�)
Tk�����Yʲ��֩[��umA{�4���7���,�f�PS��	��oy�;s[�n�b�42����N��Qb�Nm=�/ �7X�2�t�<6���9��j�6�d̦κ���b��W5z��f6,��K�*־T��n]̭��W�_r�K�.W`�b3� ����6�>����9��_!cXW�W�	�fS
���Cl��[1l��w6�����70����$�q�L����j)^ʥJ�w��͎�����.��`�1?TV���ע�T߹��t(y��Cj=�(*��8|7um�yoC��<��Aj���ٗ��v�fV*v��f5��#WsyQ�s�ǘn���*���+;z^$-4��x���pQ�/VCg�U��a�9o޼͍ݓ�{3l�S�k�]9횆�	����t�)�/�}>��P':��[�lB@2Tw�vXz���J��WfG.W>���>�4k�Z*j�׷�|������j�>V�^,ә����!�Xb�f�K��Y��^f���z�6�Ҵ`&N��B�e� �a����u�x�i���{}�Ǧ�=kJ)�ӻNPT��ε�P�r��mf�.&�&�hm�s�V�F���9[,�\�}�Ո��W�J�\���j�Ds3C���z]�(����enz�,�w��z�6Շ��Q�N�i��[��� ��%p�PI4bM��#a2{���lE����ɑ&�*��X�s\�6�`�4X6J��y�21��dE��(�4������Mr�����<(�hƌP�,��Eۚ+�"b�1��i���� �(<�k!&�����ut��]ۨ��=ۑ�Ow4���yɂF�$�(��{�JH�"B�	b��Θ"E	H�),��릉���s�w�9t�T����,'wb �p�B��o^T�)�ز����D	��mv.�8�:&i�RJU�Ѯ��vQz�*V���6Z��#�j(�Xhmu��e%�f�l.U�.��%e���	��c�-���ᾏNˢD�BŖ$P�f�9:�L�d,Gil��y�s/T�T-�f�Q�g�.ڍ))D��uN:�!��{L(�fm����P�e��g�ԫ��lF��DL�˲#� 7#����u��f(VС���5q2F�j�@���ےݫy��!�T�b˚A��E\��ҵ�)r��lj]�vj�heY���K���rR�Q�l�3"�8aڔՕ-��؇�WCf;����4����R��Pep	��`��fv�nC�/VX��\�l��fT���9�B�`�F�=��rm��jr)XZ-�ffZ\Ҏ�n�#�nmф�رsc�JqJ�֛ZF����U�lR���f�f�J#1��k�����ֹ��Y{G*S]��J��[�sB��h^�f5������-.[l�6�����,(C7R�.��;4Ĳ�.�h�6h�vDI����ܭ��mxG`2���ִ�J��)h�7^��l�ڰ�(:�fkpb��[���-��	��0��h��GK���V�&G�J��6 E�(&,ٮ�H7��֩X¬�v9%�f�#X���j\����J��s��eq���T�u�+ns�2�&�#4me�Ja�Y�/	ف5̬I[`�7[V��&*6!��u���"PVc�ek2���μ�؍`,�(ݘ�n!d�K�o[������I�q��[���ֵn���6�vZM�ƁrG��]���L3V�+�1af��B�A�4�ѱ)+�vK�jd���CM\gj�4i,c]6��EʻR$ph��� ����M�X͆VŚH؇d����[¹m�K�hw���5���.p"�ii���+�f&�e`	.��14T
F`%�������16jFͩ�*��CQ�av�
��\�n��E�Vh�+�'.�8���RKn�2ږVl��[��j&�Jr;�.-��uq5�T�V�xCS..2;],I�d\����eiaC���تa7�QI����Me`"�uSM��ZZ�B�V���N�L�ZA�Q��������_KH��H�N�uf�U��&F�]��`��3�Ph���Є4��.�Fb�q[MNs����+���ӈR�5�Ib����3��a�v�[n���:Q��#�VR�KD��=_ A�wi~�_,~�;)��콧st�!�,�	�>�ά��Z{�\y�-�(���U��;�w٬�_Y���A	n�v�;�u�=Ч�և�u�1��;�6#��a��}�7��,��e��Ù<���<9��Da{V��UOK�B��lt�'���sk���6�� �_�@{"��wι�ȃ9�}HwW�d�y��e�w�P�*&��ډ�6��q�����BB�
�R�Fzz϶�}�/Ǧ��7j�'��������+�R�������m?`%@�Dr6+�8{8��4U�f�!�mYa,m+�Z�[�"Ô8:���������5p8�]�tgH��C��nԇ�}�U�%u~��R%B������}]W���G4gbl�i���i��5�%j��%�*�͖'a<�ƃ�Y�5U���i����U90j��!պN�r���סRqENַ���\AE�%Ǟ�ioW`֦���~�~b��N�l�}�f_Ƴ�#r�c�ݠ��A;�˺���q�U�w�����+�c_n׈ݯ�#u$��P���������A}��N�+�lT�~�8�m E�Ҟn�{8<�_R#u	ݯ��*�!c3Y�s ˮ��?)����R����)st��_F5�n���u}�<}�m�q�}}��3�4J5\Z.��#���X�L��pd�]	�h������d�|�� �_��	ݤ�����Ot)��+_�S�s�N�
�����~T�x�C��T��	
,�Т�I�7�=�>_k���g"�7<lT�~���W|Am�;�=�S�u��=����|������}"�BB�!��k��.�=��e���m�0S�{g}�^[߰w��e�er�P	9G缷Ni�f>�w�\�]
O�����b��d{��㩳���K���@�2������_n�����X<i�Wۘ�:�	Hw�dW:?p���*�ׇi�
�'�f��{�ߞ�8�R��Dn�Gv� �/���AG".�i��SG�k�U�L?/���4�!��2�����K���!]�s�6�GMB܃�7
I��wX����n�����s>�#-������ wi|A��������w]3�\�pB�#Z����B��ʅdT�*_	!���^]k=����T(�d�z7w{7:��h���� �h#�]�эSgy\7�6�텈�j���\��.�R*]
��
"�������{xP
�P����:B�T�����[_"�G%|�W˵d���>E�/��;ʀ|W%g�W�罇�.��z�7·^Z�7w�Å�f�j��6V��x$����@�^��{�кY����h۩lMɦ��[(_�}S���r���*�3����(���~0�b�3��Ҥ3���wkgl�s5�-����Dh#�H۫�B�Y����/�+�ҡ0����]��F/J������M�j�n��Gby?$�����,��̳���A����0z�7�s(q�:�Eg��ݦ�}!B�J�P���-S�6��H���
��9��3�M�|f�9���A�u|���w<�뼝�D��\��6�eX�9eǜ�� �C}�:�B�eoDSz��3���o'=������(f��.�	�T��_T�S	�f�z��� �����ݡ��+.�Q^�M���Pw)�F��\���t�@�����H���Єs�P����=�ǫb:��*���_d�#5|�#u/��U	#��^s�n\_[u�Bq��v���ӹR�l�2��w�o<Ȏ�K�c"�I���=qi�"�.�CH�����sd٩��n�M�dN�AOӥW�}gK��c���30�؈�-X�JǐvJ��m)z�d��%,Z���8�))�a�n8��E�i�nSLs(9�*p�l��,e���"�Tn[Y�s�5�ʶj=�6#kQTmf�/jv�c�IZKL۶�*�Ըl���X�W0����gUQ!hj3u��: �a�,�Wĉn��t���Ts-��IV9���1��p��/��_�e�Lܺ��u0�ch�b���Gb�e�f����n����F�(�1�U���9�6"�i��V7�ϱ�y�<��
V��"�J����P��Ht?)�T��	
��a���G�"_�ւ�fc�Ga/X��B�(w��"ւ ������h�ʺ�"�Ti�
"�C�ק$�+7=Av8����K���TqT+!�
���E�
S�F��w^���cA|7k�6r���s�lk7g�[�}%|�5鏮�I��.����@��_!R*T(HU
H��6iYc�������A�\;�f�b�q���;�3
>���	*��4���ٚuz��-���\�Yn�]J$"��!��LY1.�\!ɳb4�l�{����~z9���e���BE�Ï�陋վz��;Ծ��N�:�Q�s^����\����\�(،y
�y�yzJ�x��W���u�03[I��C]1��E�e�w�s���
x��ke�t|�lv����;u�%��w%����:���+�{�#�#�TF��젾?>��kLv�<�n�v{B��P��+4�r-t�g]�Y"�����,G2�#9˖���g9g홿n�s����԰}b��-�C�'r��SU!!���B�"�G@*��}��zD~�4<��_/�{}ܼS����U=��@���	�ϥ���~�߼+�O�B���*EK�!���{�P���Ҿ�����7[�=�o K�� �h#�HwW�ۤh<	���P��*�"�T3J�ۓ]�.��2��ae%l��nЉ�/���!����Ծ#u̖o�ۀ׊�Z�|C�y�J�V#q�i|(P��#�B���+X�y=�:�����=�mx�"���r��_��j{��|:(H�B���cFz�y��ʐ|j�	�P�R�!�B�	}^�'�̂�ȯ)��)�&��w�.�j��:y%�e�΃ި�N��b|�#NZ"Cv�ۻx�2�ހ�
p�b�q{���*��E7�ڍ��$�/Ԩ���V�HH~U"�P���9=���B�ӏ�Ⱦ#u�{�.��W>k�?m}{��1�Ϙ�cA�AAޯ�| ���n��ݣ�.^�-\�w/�����{������B�$_T���M6��g�7��N&�ixmK�l�E���ft���fS4��Vms�"�qS3<���g�]~��=���\̙o}�^���ܙ�o��ݱw��H�?S�E��(T���
�*�iP��]�]>�:�ȟ�r����s�:�7��+�NFk�P���T?fnW�d_7^tH�|�;�#�H�7W��ĺ�=k�o�׺�eyd�oM�3�
�P�?/�_T�|*EK�!�B��oP��~P@��_@;��zze���sx�Lз� 쯑c̛~	��P���mV7F�r���ӨzM�:��u����׶��yjy�lyG��N��Ս5}���8Bް�j&,�4�h�~�}B����R*_HP��T�^��eY�Q���7o��oW
^���Z�AͤAW�b�P��!��++��I(�j�X����Ū��pꬼZ	W��Ø:ۣ�٥����)P��T+��!t(}"�Y�� [�����#3�p����8Y�XA��|����u� �ݤG���]=���u����/�������f����_"��ݦy�;;;�UbFU}�x�P���!�Щ��"��e�|��[޺�N=j7��A6����J�
�!B�J��4�X~b��CaT(H���/�վe��̭>T(?N>^o煏*�3��������v��@HP����޸�{�
�
�S���8u�;y3B��vWȉ�t�B�_{2<��NǨfcɞ��ybV���ݷ�F��r#��7V��g�e��[���������z�\��p#���:}wHa��Kg�_)�ZT	T!�ɱ6���&�l�M�lM.LBʕ�k6�D�(s�;F�ԃ0f�bjư�ʘCZ�[Sg�岈4�ѥ��&�0&�]��P��-�kU��b��ff��S cU꺘��F������A�isv��,HK.�aT!�ט�)T�n��"e�
�B�A���
]1.�ś6�ҍ�sUZ�LK�"��a6y/Ͽ��]u�p���&ٹ#\�A�7� ����
D�f�I+���l�"�':�[��7R��{u�b��׻그k�)�	�����g�>�T����B�H�
��S��3�oL�/���qT(H���</=��0ؾ̠���Y����T:���|���t=��t�R_	/�
b&Z�����}x�#��{o&hY� A��dA�H�.\Nr�p��S�k�y�q�\��]�$T�z�W;�A���SoMW�d(Q̅?Pr<z 1�@��_��۵�#v�v����.e�����VO������뙀� O���7P_��몿?t�{zl�>|��k�u����6Ѧ��t�F�nh��R�J�ʠ�]]������l�sA wh#��1�ӯ;���{��S=��<�x����z�P�~R/�GJ����[y���]y����~~t�c���&��z�^�N��U��ˋ�@�����4�n�s\��C9�vz�ʜ�tȮ+����]�@�ؤxz�Z��y}���f	��>���z��p?f� ���z7�0�ߧ�=+��_>��u� #u}�r�ZV��������>�:K�x�OR��*i��k�/�����W>����D?#u�uzPG��cg��;��z�{�/����z�������&��(q�"5�#v�;��n�ȍَ���x�kP��`ϨN����bϹy��:A6�lA�A|A$:�̾������N0PUd� +�5cq*�u���s��J2&��ev�U��X*m��{�4��J��*B�?!z̯S�c��a��c�k����(��:�tFo�-=ۗ"�$4��+��.��'��.�(_�"	�H6gu��ey�s}����?*�i	�A*b�[ʾ"��Ң'9r��,��9f���G]����%�^@�W�uH�����v`�/�`��Xܫ���'�,+@�;��(V��^�]b��=HV �w�3$��2�ҝ�u��$e�}�̥�_JGh[Bٷ��8�^]�\�h��4-{k;77o�
8Gqշ�t/Uə+'sSk�\��^V��g�hk�^�nAa�/F����;�{��ROD����i,�a݈�_m��\�M�z��$̫�u��dY��.���s�]�ΰ����(�2�;�y�o�nL�N��5�D�r�5c�+'�)�ҳdo������8iS��&�ǆX�K����-E����F�&)n<���u}������`����li��U��¾��Ѽl�G/6�H4p[�������i�n5�%iɛb�Yjni�x�<�'t)�]��E2�wg��kX̋UN�g�N<�ּ�����|o:�0q�p[�R�sp�k���3�R2��y�Y~�
^�P^J�rg��U`��T�1n����D2���<�0n��q�5���ҫ�&�uۙ�a�֮�qO��T�\-�ֳ�ž�F*�yn�ԗza�����If���G�����P��\mئ��t�]��o��A��gSnYbX�b�������=����=��ƺv��St�C�������ү���ս�׫��ku� N��_i�[G��n�^p���� wr}�
�����X����Z� �������M�\�.�{���&n�[�ЩzY+O����y��c��|����s�+�TWwf��m�i���B�0EH�D�\1�r�1Bd�I,��&ĘB���S3	�ƈԔ�s����W9��4;���L�7eK����I4 e@�gw$��b� ���BB��r����$�2i4R!Pd����"5�訂@�B�ȀA+�[�&��3�!CA0�E�"���(QA$Mwk�����RD��L�DcB�(���h�F2�M"����E�H!������ �B�"�4�(�i�;�Hh�@����rw\Ć0�+ATPR,E曾����:��1{��T>�P��j�BCHP�?f��|��?**�R�����{gj����ݐr�2��*���-L����Ч����T�Hi
$?)����ɪΌNOxU�;=��a�|��7�@N?*+���*E�WZ�w����U�I�c]3yjpi�"k+v]�ذ.�S��(u!��,.�c%�O-�^_��ϛ�=�T��ҩ�t�!oi���|���ɍ��*�4����\;M!@H~�ҡBC�#���f_�}���=K�Am|�7.�kw����ck���2/�#t�_�ߜ�����wá�>�(T��	*�@HV?v߳,:y�{��0���yE��y�-3�[�U��T�9�,�^�7�zw�u� _/���7PCp������WU��yC� ��H����;3��(VԻu�m����dSΆT�`��Q�y�Wr��;�kI]�z	ݻ�~���a�:�O4q��E�T�|�ɝw�=��2�Nr�yʖ��M�ϔ�ԏM�|���3{j�r�&���W��w��r��*Xs�w\���������>|���+,�h��P͎4h\̲Ѻ�֎�,WKR��#���>�!�����/��W�s��w��Xo7z,��J��f^v���z�� ��"� A�u|�#uv��M�U���t_�E��}An*��Y���=��רPB�O�3������"���_"�A�����`ʐ�K�/sh����ٷC=T��K��|��K㺂���DY�^�Jli'Z1�����C�7ӖI�8#�csV
�;��P�/h�.��c�P���*D����E�$���Dp��r��+d뷶��{�52�|۴�
��HHi�/zu	1N>k+�(ՃnY�<^�f��o�Ƃ���=#ĭ2{�u�u,R�+����4A�=c֖��^y��*R�^�2���μ�[>Or��H�ۜ�B,[����Z���V[l�F�gd�@i�ѳpRЖS8���,�E�� ˵MŅ�4���S�c����M�1S�����ݥ��p�X4�֬��VFf�6T;A�S��H��+��bA��p���;��#�jʶ2�P�I�b���H�%%��e
�e4rԴ�X�� 08/��Q���[��5ap��v�C8�֛~���J�s�e���� ��f�%��f��b%X\��;�����9�����e���e���7k��c����z��܆_�;4��U3��i�ܹ�T�(�r�Ln���d��OT�t�����{iA��Y'��{��Vr�W���ݥ���@�k�y)P�P�R/�
�|�H��H����䴰i�9��k�C�
+5R�!��,T����Rz��'�?z�o�Τ_*�}�������>��_N>Bz��_e'�v����@ wk庾ݡ�w=��>�f�v��7����s2I�b���_"Ȃ;��;��X�aG���6۶6�jj�ĸ�h�i��Q�@CKe9�e���P�������}�;ϧz��|�R���z%������^�^ر�%=��]X���{�X��U�9e��.%�s�Q^��X����yl�ˌ�~�S�sn�iy�L�)��Ek�j��^�s	��y��B��P��ve�{�RU��<^J��_R �@<�s ��]v7���3^�g��y|�T��5i2��We����D�,��(�^r��v��1�����r��HV�@���,�K�!B��/��[N�J{꺶pVm|��|�u<���{t;F��UzPwi���1��wTu�����*C�>�R~�9^�'���<�C�M��:]*��.<���9Ԉ./�o���<�����3���;:l	�d�q3�X٘��6s�h�Y���lڳ-�J䂹�2�/��O�� ����x�mX�3��3��}SvM�+x!�)�T�2r����g�� ��_۱`�[�Ev�ݫ7���%G�o��2�:�G����w�;F��UzP��v+ ��n�r׽o|��%����� �݋�@���}X��Ww�=��=&�v�ס�2\��g$���}0M�J�tg�mV���^����!�visd���, j���";�ҭ��<�]`�s�C��Cn��� wM/���q�g[aE��U
�R���ڿ��v8�˸��&���m|�]2���J.�>>u��_"h_ź�6�D6�TX;��޲��ys�ow���v�}�������������U��|g�{>O�C��c��4HIP5;��c�@�Z�H��s]��%Al�T�o���@���	���|��|ff��w\��^���qp���ڿP�{�E��u\?{���_�6�-�D�mY�kS^�~�Ս�6=����M�2��ྛ_ FF���/+����� ]_a���:�n�t+wW�[�����xO��'�Oo�WB;C}������b��؂-�ڰCh=.�c���A�v���lX=)���5��ΕW�۞~�R:��U�~�̕h\��o���S��<<s�*[�2�m���\ع��ͧ���t;���쬎�˶�{Q�Ӗ���y����"Ib� 8���mY�źߥ���La���Fl��ޜn��&R�8ͯ�cv,�7W�X47�v�Xvm��$X���t�-e˫@ Q�R^�ŵ (٘����V__Q 3i Aq|�m����&�'�v�����������(c��g�y0A�E��	m�!�����_G=�i&,=�g�� l_"�u�oB��1�Hqޥ�WȆ�W�b]u���	��A99}a��t< �׻v�x��K[~�NUR��*�o L���݋��_&����^���U;s���_h��K�����=5Q�hv��yG·|A ��E�ػj�͡|4�+~�A��VCh ~-��6�X-��wJ�o��_]�ɼ�Ύ�̶矁ԇ�HC��Cn��[B��Wt��M�ܕ���ج�i^��U�fo��2�n:�X�q\!��KvS�c2 ���Xj����}m7��1�F_�/�g� �+	BcYk�0M4�UG-4��&���p��m�k�X��64��0�X�S0��pݜp:1WXZ�5��n��s`�$�!m��1[2gWD���heY��p�H���B�^4H���*�GnN\i\,�n0m���]�Ep�X�\(�F�,�:�����Lݪ�ř%���yBS)a��%��Ą��4`Pԕ"��Վ�s������`�	z��w-h������De����;�*,.�ۻ)X���P{ج_ ���[kz���s4��;��n��ʉ��y"��+��}/���{�[_/�mذKt�oL[ (�5������_t�[\���%��8�syX ��"��!Z��~��K����k�x&u|�݋�D����'��gCr�pN�A��=�z�5�_�Ԁ"J� Cn��[A�g�w�7Mf�$������m��y���3��㘬V����������'�N}+�_���D7_"y=���A�f�������������A7��6W��-���2�.�n��^sB%bmq�����e�nu����j`�gYD�̋EBV��@���F��e�D�����:��~�ny��X>o;�Gg�;jL���������A�m�"�����̵eNFn�0����>ty�{�:����P��:Ƭ�vD�6��R�	��F����ϊ��_)�q��s�xa�%�eA="��=�0�%��1X���W���n�a�J�eX��DzjvR7_"v/��h?y1�*��_ml��g;:��G·	��`���n�@�Ր�B�n=�ys�>���#q��Vk���Ƨg��������� �R 宂nJ��?�g/�kA�%�����-��o�mpч�S�.��7k�t㘬V�㒾@�1�[����؈���7Մe�PI)G�]\�-"�Қ��a�:m��,"3Jc��bKuZ
���5c�N�@\_ Cm}a��u(�^K��x�y@{�r�eU�/�7@㠁�v���;��<����ү �ϻ�,�t����?9�ڝ�{ٍ���ޤ?H�D6���f�+���@ܠ/Z�mt��m.����?	ޭt�]
AP̬�a�+�X��JT�N/r���!�=hC�S�f�.����Ij�g�`�E�eV.�-Lv����VDګ�3�F����6���ʑ�V+yJ�7b�n�6����{����&;�UeB��Ȉ���6���B�^)�E�x��C� �syYs�R���ܮ���}��k��`-�Ȃۿ��SJ���[$_!s1�w;�$�f73|K��u�w�[u�n��x���hݚ�E��k���	���Ȓ��
#�-]FUᚗ.�Ef�*�����~���mX٧��l�>�{��ўT�4�-��
�K���HCk����Kt�!��XM������}H�=7R6�)֝��	�87��6 �t:mlx����@��`�����B�n� ����z�����(�N�o�	���.��}%}�w��@v�E=��QܼW�w ����ڽ�/�͞u�jI&+z�Ϗ�U��j}��C�Ű�s@+��Y�z����V�]���@M����S����xU;W6�}SsU����c��Ѳ��@��4[<?o�ޡ[�u`��"5��c�f{'��=ε=��u�Sn�;���8=(7����n��-�%#�Ix�]T��EE�T5�1��e�^#ns�`E5↋�sD��Pj�m����_$w�u��_!�~�o�����\,;/�س��դs��������h"�A-�^ԂŮ�㾌Yn��8�x.�͞���I&���+���n���ӃZ�@on��Τ?6���|��^�G؄�j�FY�Oθ{� ����. �n� �ڱ[���c�j>��k��]c��q�7W�|���[΢��7�1u�� ~�y�m�}����^E�Ⱦn��m����k��M�k=y4=��b����޾T�b�I��o| ̯���_[_>���ɼ��&?=n� q[��|�oN}�w:@�d�5��\Qi,��Blj�]\����ʮZV�Û���"M������Vr���v�6Xǃ8isW^k���h�y�X���K��wfJ���`˼C���P�:d�vh�`2��-w�;�'����\�#�th�F�;����b��͡0��Q��\FI��j�;	��Z�i^�Z�<\�;1d�an�;ٷ�����yk��h�W6�'n���:�v{�+�5�+N��]�j�|��f�ڗ{lS�v�>D�me+�P��7մ
��f�n�j�4�u�q$ʘIQn�g1Yٔ��(�����}�t�f�}�_t�dn6�gs��tَiK��gv��񳘩ďù�廬�zn�����޲ѽ��(]d�$�]w%=[�/H�2!�6���#�Sm�'F��3%�g ��r;R���m���.vC��ĕk��0; 'gr���jv=��K%1�,����ޭ���sp|�o����b�%�'�Ռ��j�Cˑ�[$ʴ.��e"�����X�5,=�5�l_.<�w]�{�q��XM�e�������v�+㺚w ���G�N
�ݢ��ξi���S���dR�F�r��VK����b\�͵�5mA�[�^�4�=�,���4�M9,xS����21��/���v��G03+h�Z��m���F��:E]+!|+p�\\��2�P���9M�Y��O%.{��]v웹o��� 	��T�/���^�Ƌ8��׻PH��(��wpL�C�-]���f̀�Dh�NCb1��f�LPJDl#�Q���I��"ut�I�B)r�A@Ț)!` ��#I ġ�A�H��l%	�@e�d��71"Y(��wqwq�0���A! E�D�&@с�%")$CDS��� � ����@�H�1#s��C B���La�ŉ�J���
4�
"5�rcI�P��bƒwW ɀR�Q�i�2��n(�"R�D�E��t�5w.�
)��Q�WwS$� ͙Y�b`�M$����2Aѥݹ�W.r�Bd�fIA�H�)�J���̄(�D\�Rh!� !!�@��~z���vaV⽵ut��"6d�l�I�AB�n�ޒ^-�)�fn�7����`X��!*.p]��- ݊p�lf�JD�k���[0%���\]�`�3+�)�h+��X�5����X��1lq��%�ųBl�,ͅ�g���tee�Ԛ0���#4Ɖb���8�T��ˮ���m8v�lSu��7�bN���Y��GD��݅�U��HW�]j�
D�J,���m7
Gg�6H)fq�*jS,Ƞ�oZ�Sam5�U�Y�(M��m���DJ�Bb�-JFL�u�J��̮{d�p���f�U0�ݳ�K�\���1�X�j�2�+�(bԁH�	������#f�k3�c��J�ʌ2�.��bn�F4��Ř�2­
�eñ&��WK*M�'���)�����v��e�r$��"mD�efv&��Q�fŜFmi�jܬrWr*\mJ�ݪ�ƇcL4���,��B�\��S]�X�)hi�(�pF�ۊh�R��ޖ*�Lmu������ማ �fu����hĺ��@��]��խ�Y�SWx�Ԗ5�\�lR��]�1����Y��)m�6�[d���Gmuk,h��l`��BhY����Lt�d����BѠ�G���푛[�A�h���&�ǒj�A%-�:��Sʺ�d�fU�L��ٷKD�,v댦X�JK����h������(BmmY���W`�r�q�@N�n-.	�Z���؎�VZ���3(�1҄�],�����u��f��=��� ��\Mnv��D�ٖ ��f�7fh�*0�f]�\䔗��ͨPn,v���"d��k1���HW42��� 8s.�ݙu���9l ښj��V�u!��X�̷�@�-�V6�-�h[a�`��5�(�ݜ��n�[I�u��ictp��hRe�&t���$Ѥ�m�]YlM��$RnЍ�6����k.6��KG���
0���6	���3�kli�ȹi��-��QK`�6�d�,#�T���K-��u���1KĆ��hL&�^H,�A��8��v�`���"�V�)I���k�Lږn%��,2��L\hV@�E���jT���\��x���"عe
Z=a���P�[��-nb�֖��,n��2�4&Ti�#R���:���Pݴ�Gf�\ǛŬ�aX`�^�L���\
��mX¼��߿�?K(��������`f˕c^��)G]t�fY�IF�5�	v5u����뙺�D�X'{����_Ü*�p�c��҇*)s{��=*�c^�Fr�A A-�`��@���~��,�՝�畤�r�o�����Vө��o�ć|vW���|�m�1okե�m���_� ��Am[�� ��Y���g:`����>I$�b���fW�}�ذ[����m��9��w��J+�� �~_"#����p�B�m�=�_��@p;��}��Ǒ=𿏝&N_7�^��
�u�"��Q��e�ӿO�_)���{=�E9����1p��;)_/�!�w���G�����4�b��P��3�5Ԗ�jfR�Ѳ�u�Pt"˥�k����|ꡠ�f+�/�t �ڱ�x^�q-��MV+y
�Y���$�y�W�Go/�� Cu�m�[���m�
vޟxrT�A2oU�ٙ����p]�7N��-r��<�n_+�M`N�d�^<��quo<T�a=�����lM_A��q�
��p�oT���C� ��V!�n�v�"��Z�����ޯ��݋�@��k�&矴n_e�6q��_�#_golt9{�i�o�Ȇ��ŵ�t=�#����\w&A�D/�"Ŷ�lG3�R�9�b���k�G�C�T���s�H{��w`�� Cu�m؆���o�i����z��v�^T��]������VF��A-�7ܒ���P�Vi4Ew@�*�!L�Nma
(ʹa�oj�-�u�1��4k��g�ւ���
;�V7J+u|��[����ίzI�b�exbݮ쨦�}�������t�mX"E�.]�]�Z�>�4���h��n�+8E�dڱ[�6�_���I!��g�MO��B�ƾC�3r��A�H[_ Cn��t2����W<���b�g,�k����x��q�#`,y�Qoe��'q�tnX�fm=���3�G�O`��>�Wxn��"���8���Ŭ��w���U����E��6��=��l�=_Yx��ԁ��o������6׼��1p�Kt������VՌR����X�؂��VCtn�X��qUuW�7�����p/p��dڱY�6�[�����a�K��VX��G M��W]�VRܰ�R[Kcr�#��@�J�iU,v�쯐�@�݋����nXWt.]�C���R�Y�^�a��դ1�?6Ր�u�ͳ��P�s�n��`Ò�r���͛;؟���$�b���C��ޟj9sǈ�O>y��?���+*�PE�|[k���1�~�q�p��ɵb�� ͯ�dv,�Hk�Cn�v!���\��P��Ӳ��[���d�{�BwS�z-����+#=�M�~��>^%��� ���ʬ
�h�؞�w<�-evRGE\�1,��L�a�G-퟼Ԃ�պ����P����ج��e��6�_ź.�.��H-����ol�fߕ���b���A/�"w�[��w+k7XB����Z@&AB��]K���X��-f�7d+��e�j��Rn.��}"���@7_x������6���)�ɵb��*���;t��Dƅ�vR�m�`�K� hWnӴ4����C]Vm�W�t'Jj^�n���+l��n��}�Z,����!��۱�An����\��9������.��D��6��!��=^�y�P����}������W�����U�T��ڱY�&��apK��?N��si���!�b�-�[�tlk+�|��y��pU�oӺ�S~�\��V;D7_ [kr$hő�"ڂ+�C�z��k=�z͑�U��'����]b�ڻc]��Y���>;g��w�,�]��d��lJ�[��>G{����u�Q���`�ΐ�Űl)qa۫-ըnr�C�jᑰi	��f�U�Yx3���gb���
= ֳ)�r�fS�hi`=�ɮ�&�]���YMfQ�DY��)V��a�B�T�WYu�jRU�*l�`����.f���"�j8�rC�ZR-q���R�+2ҶW+��.���m�l�)���L�Wbv�n�HU����Y1iX�&��F����%Ll;�W�:��L�����m��{�4	����e�@�������2׽�@Z��ۆW���3��2uF�`_Ŵ7H��VG7���v��X���V�F|�C]��nzU��;�&�@�2;�-�,�]�Rmg�P���K�	n���݋���OG����Zk:Q^��x�J��u�wܯ�6P_�"-�`��S8�����G�pJ��wX�vR[��3}���_�׽�@ZC�yH�⯔��u����׾?6Ղ��n����ټ���+�_�vmz>�]�lnd�܁"m�dv/�� A-���U���3_�8�>�IJ�!q��1�n�ܝ�eX)[^�`3.&hɐ�Ckl:�fW���6�_���CZ8�*���]-�;Q׏Z~��j�$��ڰCi�v��X���ۍv�����dO�&�NVc�|90J�K�����@�]�Ξ�mn�RA��XTZ��c2�k8�3��#�u���c�_��z7����@���r���ݳ�?e4���_[h������znϕ�9*��*���\�V� H�A�7_an�m�~�]��S~� A>������Z���y����[\A��ngIUr^D�B�h���y��y���/�6�X��=��ވ@m�C�/���W�^�n9��X%�"��m��6���mܿ5���6���P�6e������3j��.U�Rj��VQҕ��+�A1�L�q�C��� �[kGY׽�u�-��J���{g�P���4X���b��_"�m݂[�~Y#�2��͝D�C��#A|�â��p������r�6P@���2�َ�e)����yC�� �݋t����w/hI�����լmZ��ڐ�9j�`�ڼ�T�aǨ��F����T}\r�<�s��Z�W�{w.�G4�eW���F�n	��P{[��þt���rK���D_P��m�#Fo v�b�e5(��@-��"���ו���J���D��x�6k��Rƀ^R�(/�m���[��!��\~�k�pz����������-���W�( Ct��7uN��OC���i� ��?%@�.;fg4:�n�����f]Q#�)`D����s��f*=(�/��"-�O�}���*�����ۿmX�����
:�!�`_Ŵ!�D�V�=Օ�m6���� ~����Yz������s%x/p@�D���u�\�l�\�����#s������Cn���͡��3ɏu��|��l�[��k���U�F����Ր�Ag��<��z� �;�� �� �=�7�?:W���Q%^ҖJ��X�G��l��v�k#w`��2d��� �U�ܑC&إ�Z������[��h˦'��t�=Tr�'����O����2X.����9���mY6�!��mƥk#���-W�^���x��9��/r�� �v,�������Z�u޿{���.-Ż}�%s�ʴI�����T� K1ic6�J�i6�V
���PP��7U.�'P�{*π��v�!�[��iw�D��j��!�nW�������� gPy[���g�+���ip	ܯ�u�"l���͢�>BD��ϕ�mYeN����y��8I���^y�G2V���#����2o�{ؕ�͙��2"l��C�=���h����D*��+�F%��P�������Ӡ�֬�@�Yd/�-�����XxK�eO�y���<}����lq���r��������c�wܖ%9�y^i�ˈ�$�V%�+��۹v�:^�=�4|n��f83!����/�ϻ���.��O[ך}�sĮz���~p��Btv�M���F� 8.��%�ա�j��f��&Pc�Ye��#B�H�J�=F�7tX�[A4d�����lGu#������M�XƗF"۱�+o.�v��2�6.���P�bYlMl��&1�Қll��cR�WZs�=s��Xh��J�+m�r�YK2��c��m������+���H� �L�*�n�љ�њ�m�������:�2�馹��DBl�B�f��4j�i[����&��UI��O|��?}#�㠈 ڱ��c}�˳ڲ9��/rU��=��fKy�������n�����ȭDuO�N߯��D&ָ+'�gxI)���ݪ�lA�vn�J��ˈ�A{��> ��X-����k�^�`�y�wA֮L�ٽ��_�8�����@���6��A�";�}�N�C���;K~ �����A	m��9^}:��}�#�+�m|����ơ�gm_�uyWm"��hX-����y/�^I��1܂�|+g�gx�����:�n� ��m���Jk�t����}����ǀe�yJ�m�%��K-%
K��m�Z�}�*>���WBC���s;gE��ٱ�U��\���w��|�j�N쿛��t �[j��y
z���U��R�l'��+r�J#i�jc�����|1��\|�U��l���k:fNؔ�u"{�s�$�N�����e���J������u���G2V�f��I�WCt�N���︼��(��]z��~=Ծ!��۱���5�/_a�������л��F�������j��:�_�"��Vn��cUa���o���t�-���Y��ݽGV,��]`��_cOGϴ^���=�wP_�A��Ch"����M��+�9Y������f��f��q��n�M��qκ�=O��:}��b�M����f����42b�����U&f�A.�(�n�.�3"-*�{)|A/��6��n���c����v�ц�*�R<�7�
�"�%���u� ���|4��l���[���[Y��':�lq����/� 8�@��k|Fex�z��V�7��u����@�A@-�>���O��w�/��G�5�]H�z�f+�%�lye��i��6��W�摘GЀ��]M
)���8q� �M���ӶΡ ��Q�a�D��ڗHoT�m��pj�\�u��\�᳸��\�]���:o>�W�=W��g2%$v]$]��P�{{��+,��C��$㥮xo���g|��'����11������j����[�y�� �ՙah�(�{e�̺gŻ�-O�-KU��L-���h�~"�U���rdb1�ǑQ�m��M�4XgF�nU�O���˲*L��q㷋�g�ՙr��<w&I-�V�ĵ����)�ݸ�r�l��!�>uݫI;^T2	s7f�
���6�H�A���ҫefn��(ĩ�v֮kw�M�D8��I�`�O#kj�9+�U�#�9p�[��SAv�^1y��0C�ס�^?Y��F��� z���M��Wٺ�2��Iv���{�I��*[��u��`��\���ņp)߇|魤T�g�Q��x���,Ry���$\���1�F`�f�|�ܭ3*����i�.��4�=���Y�;oZ��<^U��M/�'���x݉C�j��<��Y��w��pYחN]�ڙ�:��3 '���ԙ���=�|�w}��ݿ���e��u��c�y����ƬX��8���wa�KR�^	gz��=�M�d�\�4/�2���Ǧ�y�}tKwB�i��^Ñ#�o.)�wo�f]�H:��˓���Oc������֗�A�am�J���v��ٚ�y}8gG�p���b���	DX"an\��"$a3�"���H0P�!���("Jm�d������LI��J	07w!��""�!(�P`�Ms�&d��c�%�II�BH��2RH�@�A�t K�fRw]fB`�IX��D�dX؄dRh��L���b�Y�w\�@��P%��HC1�Ȱ`��AHhL!D���ېQ̊ؗ8� 4 *D ɲ���h�M"a)�RJ�2Y���c2,����2&D2,DIBTRY)2j0(���ɲDf$F$H)JL�`���H��CF@#0�I f		"*)���13L˝�4aX��h13`���lA7u�E&K�B%	\�_}�^��Ww2�nnׂ�|��_ A�`�H���ۻ�W����[�!��_�����V���N��}�;�[C�?sVA�G��# 4�L0{h"	�ՂA�-�Ȃv,�A{Y�}v�B�wvfN<6�3c�@kz�ܤ!��v/��=�k���=yTO�B�#B�a%3,\(�;B�g̲�`�J�������2���?�	��V/�������m��ʯ>�e�ڰ�BPZ| bN�z�_s�ŗ)Ck�Cnł[������S^�{k�~`�ͻ���)�\ԖwU���Gx+hq����F���_Pk�1ٿ/���#܂ί� ��X-�����f\+��_������͐ް~;��|�@����~mt�k��'���� ��:�m_�2���w��r�/pTC�a|a#�fuEh��n�����f�E�t������eq�&
�h��)uh�۠�#�M�xn볷R�fǚ��v�lm^L���!d"v,�t�e�}�����}x���5%��o}أ�:~�}�����~@�Ի=ٷb��WԍU���5ն��Z0`d�,r�Q����X�j�f�ų����ou�-�ɵ���ly7���������BS�ma�~ŵ#b��ؿ����� �Ղ1`ʬK%�`�J�M�>ٕY'�~]�6o��� L��F7b�n�k��ܨ����U��#}�`� A��!۱7A��
���%����W*:~�}��@ւ,��?ڲ_!�sܵ��~ުF��وYr��L�>�~ٽP#����Ծ�WW��,*ȫ�#A;�q�e��m��6�����.����������ٹU8��W���f��/w�&������x� q*�*�ջ!�ɓ�v�h%��������'��6�����;C{��[
�{^��`N�貄l'�V]�mѝx��ч�q��n�Zl��D�}����-�jʶ궻v0�+�ǝ�3�6�P��X��c.�-m29�Yj���%�C��:i��X�l`���#S����ڶ��-��-a�Pk��n�яŹx��Z��X�VXZK�殕�UĲ��な�a�����6s�2L;V`K��M�n"��r�6�VṴi�=]u+�fӭp�5�h�CP�ֺR$M�K�@����Ȑka����2�v0�[Q
-��@R�UIK4�6j��j�,gX �A2P_ۻ��
V㚳��i�V�ǘ+k��h�u��b�ʼw{���]q�VCh A�D����QԽ���� �%}{�������H��z���ۏ;�����7��D�F�������wQ�ٔ=MهO��&���:3t��D���݋��_ [���=»�Kty�w�~�@wL��m:��;ذ��}Q���++"�굷�n��Y��7A[v,�[ǲ:ܽ����믦�j=���̐]���H��Ak�mo���}�'�&�?-5�5����bM5�α�CC
F�WF��쭈ێv�U&���}~��/}����[j��J�<���js��갽��v��=(0Fv�`���n�6��-�"����o/��~;U�{G���u�jգ�b2��ig��_h�`�O:�af
�5�������]ރ��Dj\�/pei���~���xˈ��J��C��w�BV�6�v,�7�T�`����� �5��g��~�0��`�����nł� ~n��:�5&Wk�q׮l��W�������������>��{}�6����|A �e�A/Z����vΪ�S�l�U��p����i�z,������D6�X �C�B6��bv������ئ��w,ͣ���}�Q�A=5Y( Ye|A ��[��WM����j��]�IUa+,F�������B�&k-׵cH���l��y߾@�g�@����e�D鐾7���>����͐V���0t��i�	͠��w@7^ ��_{�5|+\����,��W�W
�Uv�:ٞ��������1�m���]�3j�˿�R�Ȇ���6�"���{���K9�<�K+69Cw���M.��]<�F��N�ƻ	�1݂k��Ʃ�f� �!ebnI��b��3_i|OffksMl;�}��8A�� ��/�t����Ct���U_7���\�n�@߶:�;�~���͐V��AyH6�G�,���V���f˿�h"� �Ղ��-�۹ZG��m�_����1SgU\��갽�/��ȃ�k��� ��=b�eu�8��*lN��,#UCq�F$Yq�c�#V���A�t��`��LJ֋J��=��?>_!����n��N���Y��0�h�zw8��h�V(�� :�>-�d7_7_��m!���+� �_ o��I�|�Cu� :�� �����!�j������RW�ۙ� �A���mY�n���m���_�zD�n��ˏs'�܁m|�����Ȇ���J�~v��b�euܯޯ�r��A}5M��y}�����ᆽ�
�/���/,� \��ْ*0ε���	T��xz�@��-T���[�3���6�O;Q�õf0.��V�����[�<�.L�;㞠�?8��Ciu�۱`�UG%O,�]թhU@d�=�d���\r����R ���۱�uS�e���8Q9ugL�i4�`�h�p�;b ����	�� �-�@�u�WJ�6�q��_/���Ŷ�|g�������A{�ú�>�O	|���@��,��� ��D6�X%�_u~-h�;L����#2/�NA�T���쳛��{�[C�'�Ղ�-�&��ӵp�U�doP@+�A�[�6��Γ7���8��\r[��/)|A�y|�m���t-�DC6�Ge�I�Dh"�%���p��b�w'���ͯ�#��S�7��:G|�s�r�w����j\�nZw���"�7=���Țt�g_O^7�{]��-���	��؂���^��Ǔu�����Yr��7�z��ev�(�;�rF�l�O6In�Ys���sȹq�Zr�����n`&��/���>��Q֣Cpl�PIB�E�ʗ`5��1u���Lݥ]��TB��Z�7:�A�͎����!��v��f.�@��"6��0����K4�M��`�46���.h�qm�^5V�.�!%XL�&�:�u����n)(lT,
����H˦&��7�15i�j���2�K�K�Gcgl7aP�F���aW������.���)���.�՚�f��.s����Q,yS0"8t��6'ğ�����>��B�"k�}�Q�֕�ɮ9��k'�^�U�X��������t��VmwzVz,��e����+����������Az��� ��l���~ĉc�Y+_�����6�@ۻ����S���E��j�ݗ�L��ץ��=G|��e���Z1�{z�������N��1���A3�X�|�m~�n�6�n=rH���}:h�������w���{�Ŷ��A�K|6�xʂݫ�aI�˨���M3�U{�&m|� ����[�����[��n3��xz�D���-� �k�FvX�Љ� �2�JWpȗ-�Ccz��l���l�������t���S����0�'��S�y�.�x�z�I�gWӨ{�~m�6�%���Y���*��y`/^ָ��Ѱ�>*k&��y^�	��ݖF�R�5�o�!Hf��p��۽mi��'�-X�_�:��	�ΤA��@߻ �`\�n[rH6��@�7���̏��R'�}y_c������6���AKmx4�E`C�*�}مu/Q�����_t?5ؿ�n� ����+k��]W A�_"3����h)��ٱ]��k�z\��8��훫��cRқ� :�"�6+!� �_"�b�u�.�B[�������K���n9ԇ|w)|A�_ C�_�к~�{9A��[F�������d�P��,�Ҵ�.�����c�jcmq@�T,P��Yt_7C��[j�ʻ�QLp7���(W�-,�[q�$���b̔��!�B�t��V���OnQ��m�"ul��j�uV��E<t���Րv/�g)��]j�fK���v O &݋�@�2%m�l������^���Y�n�>Ɏ�mN�j�;��3����Ԗ媘;[�*A�V��ب��l���=�P>��Q�-�Wx������zM�;NK(n{drs��*�q�Zw�֢�νv	\I��Y2gS�5y��Q���T��-d�R+�8��𧆬U^s������6��-���"}�Ӻ�ڥC�;�Y^V{��8~��j��;׈ ����6Ǹmf���_������+G����S9�,qD�b]��)Sr���n�&w�����[�A-�ֻ6�K473dr[�X�;�T*�a��erX���|A-�`�u�sv���)��wR�Ȭ�>~�����(W� H�Aݗ�u��&*�z��TUF<B��H~-�D6�ẫ&��<h�f挳.H^T�a��\A�� �� n�?6Ղ�{�b�ޙ-�(x}%�;)Kt7su�r�����z����"��E�R6��Ï؍ۙk^�*�^�3Wp�.�4NͬN���¼p����9��W2�5^L�-Z;G3�ޭe)��;~#��w�����	m����7[�$9���#�3������^��;eF�W�D��а[�A�]�8GP�q������Z
�&�%d��s���q2���z�ʸ�ٻ
RmVb]S�����=�%�ۻ���=7T��u}T��ʃ�\G��hݤS�6��U�A�A� �XCiCu�)[񚶕�,ͤ%��k}����5�b�:�9ԁ�PD6�UǴ}� ���~�Ր�� ��O,mn*�#ǜ˿IW����*5B��C�u����t!������u���3������[A g���M��g�T����Ղ;-�Ԥ~��7�A{���@��۱`�G�^�6v��;ق��A�3d�F.���w�W�0�~�s�8r����	'���֭��U��m�=���m�kkV��V�ն���Z�߾��ն�m��[o歵�l��kkV���mh��HH@�zHH@�T���$���m�{kkV�鶶�m�{kkV���mj����ն���Z��e[kV������)����S 	�o�9,����������0?�� ��EH���Ti���i=E��(Qm�E()J�%-���<�J!O���@)TT0 �&    &"��AU4�     hɉ�	���0 �`�0����@�� 4h &�  J��i��jO��Ҙb��C� �4zAACI�O�@��ze4h4�i��m#��;����DHW���� 9tE�( 
�%��@,+��s�'�J� �@��A!P?!`(����)�
��A3�nj���� O/g�����($Lj�k�頁��J�����JJ
(��ģz�m���]�[�kkyh��B3kPY���wS��MmB�rq��Ԯ̊�5�W*)�kc<�V��9���m�o`���܍�ۃɔ�D��c�x<k+m�.���1K,H��E����̩H���c��mސ�dM׌.s�u�1[��U:��7%)�V�F�
�˩�B�݋�����L�̨�6E�P"J�;�/VȖJy:�����q�.*�<ٹ���]f��fS�iE��Q_���y�-:E&���jT�$�.-,��VEf֗���݌�C���[�wj�1^�P]isK7f�z2*���Hj�Ā��5Z���gϑ�� �gm� ì�g`%�p����f��	VET$UEB���d�pqn<ݘ��" >��V��m{�
�ti��C�v=�`T�44�8�]Rڹ����-��36L<cᴌ%M����e��z\��uJ5+%�Mć6*"����%slD��p���T�G͊�˚Иf=	�MA�(f3�M��UU7mb���Ľ>aA͔����d���%5
]�QPK8��Ց����owj���扙Eº����n�hv8��!lWl�mPX>T�B�J��5�c��S��˞mNd��p��,I�1�Gq����)��ܾR��r��E�MT��R����J�����!�2��K1n()l@][˪j4d""�2*a����!�D��qb	lV�8@($	"�>(rC�,2$��]x�ҡ����܉���A'qIjXHJ�,�(�%��R	&LL �[I��                  6�                   0        m�H䙅  �!ĐȖ  �58!��r���a-�&L��&\� �vD�Xے�R��'!,��&&�Cd��0*��H�.$�1��Q#Bw�7ܲ[N+��;�t�.r�RI	$R��Q�rm����;����\)(����:��N��HA@�X'��%���r��R�"B   �     �cL$@�@1�s� $�b[!B`$����m��-�������R���I��yZ��X��h`�g�/�p"ő�h���&.n�ec���"�*2�C�N�%�s%ėx�t+��-�RI$�	�r�~7ۛ}6#z)����f���+/E��i��O#�J�dѓ~���2]�YF�i�4�W5t>�y��=�]��  �;�ޛ[.�Y�otr�{�L�I���b���>���v����/������F+�9@��b�T�/�}��1��")�6�& BBqՔ��)[N��X%f3x!��(�⧚>A�l��U-+�}k���,4�t�ESE݆8�Ό���  �7���+�����9��f���9���n���q_�G�%�U,M髺�hxJ����u�g�'#Kg��C��~���#�=�9����}�o�RI$�I��)�nw}��!���:Q9/p�����_���}?%[��#���>T�A�ך�_Z���*�2v�q�>|p� 9��� �ϻz�&Y�EM7e�V)K��|��m�i*���Ę2���B3�k �@s�8��t�����dM���A,2|�S]R���80        �����nP���[!K�9l�ύy�** 	$�9r�s~�8�v0��0\�٨ck�� �a��� 6� �1����!8�*A|m~8GD�X!����*�$y^��I�I�IE�$�H$�H$�H$�H$�H$�H$�r�t�|��I�I�I�I�I�I�I�I���I�I�I�9��D$Q�}��lN96v�"H����x�ˋ�\� �/���S0�-�C��q���6��$�I&N�gS{�#�A��-7��z*	P���Ȓm�} f#���焺�m�iTi�.8�M�ŉ6|�.v��"��a���p�)�;G���.��{���m��)�Z�ɂray�.|���B��@�  lu��üA%�i@D�[�S`��\ A�0�|p���d�X��!��4G��M��}���<��B�����i�T�͛!�o2���#e�#Hs�"����Q���	�I�A,	aI,����Q��^����(��f]�Ԙн���p�l4�#�F�MD3����Gp����U	$�I2H���ߖ	>�!1Z��u�V�uί���U�lkN�C ��9bb'�I[�k��I���.����
 ��@^r�<ő.�`�t�ArO�����4\�Н$�I$�"�un�~4E�,��p�O��u]�p֌~H�H���T� ⟾ħ���2_ğ�C�S�W��~��ˑ��X��\��㥛SZ��0��B�1>���u�a�V]]���ɋe�:�yso��E4n�#�y���8^���4Q
�YPIf:J2]`��Life���P�c�h@�        �H9KM�bY"�9�ș!�1HL�z�)QP  ):	+�͟;�h��rH$3�;��<��¥
���'H��6D��G(Ed�)���8����}a��TQ�L�E�g�t������/��}�m�gT�2�Mg�wȢ�  �@�z�OM�>G�,$��Q��o�q�z��q�g���O	�W8b"��z�1�>��g�P+iś6|���V��L5���rǏ�ffax���Q���O�>=��q  ��{����^�Z�S$>��T7��_�ZXl��d���!�&�?��m鎞�9�8[�R�S�w0��]2��x�Z��ʕ�A^2U�VZ-r�=W{�oYBm�xU2jT���~}�/�"��8o����얳~�b@��il�z_��� i`�̈Fu�#_3$   `�g��}���U�N[7yT�w-���^�,�Dt�-M	�,�"��%]�å��z���j�!^l�.|��=z����H  �3��M��бK
K[~5�n�eG��z��V��Se�FzcA�J"�i�'t�������ʑ+	cT�>���ssqa����λTYn�-�˝�qq�˻���J��狔��U:�U6��I���          �")��AJ��3$H�@ԃ���T�  	`	�w���GEV$�*2kb�c�	���F���ɵ�}��J��eCvEFeA��D�;��9]%���L�"H!A���q�`  	c	a���N�V�s����Q���N�xE�g���M�R�����P�l�}q�VZ���ur?X��*f��6�s||��"�9p   �9�Y���̳4	�v�T�36m����\������~�O��=�=�2�n�ܥ�&�ܵE
n�P��j���fr���<:*�A��x�T�>܊%0����ˆ��= �7'�F5�C@������   bf{���/QST�6_f#9�^���w����X�,�p���<�?�������6Dv)��3�k��[�Jr��Q���rswn/�'[  �I't��}��o��lDj�Z�'���sE�*VP�-�hTMU%O5 �Ⱥ�S���q9�u\1�[��FӨ����""�2��-tt���@j\�E*���N��&��!�X         c�@���*G0
e�CP�!�@�	�3��
�  Lg;�^���=����˞�Wv'Y�ڛKQT��a5P��U&�S�*�d&&9�yIw{�3�2�L�wUN�0  �[����[L4�3����{�r�Sڷ�˥n͟(�Cu=ޛ�	*��"`��3��0𣓷�#x@� C
�w�s�Q�("X.U�L���6�v�����6�ns������P�2i⡞d���e����[r�9�V	m�˜]������$�1쪂���:t!� (Q�μ�����E�P~��2d}S���~ܝ��@�y��   �2V�9ڟ-�gI��l��;6�lcC�@�����մ.ƆkWV.#o^3y�WHu��Q>���x��w����{t� "_r�b�W�<�m50��C��]ч0�	�c�Q�e,��//q�JT�L8�ؘ2b5�7�f����ǎq�_����$���}�z-1�$$�Y*�PIj��䂂{|���PN�$�q�-��(*_F�b|>��/���F���~V�t�(%���`Rn��Pox�n
Zڃ�=1E�^RI�il�Oοd�F8����ߍ���Lc��؄��˧穮��7�P����!� ˛�tƅ��E��n]����"���"*	�M#"`ZB���jM@~ľ��g��K�)�-�<(�������򯝃������y ���h��Ӹ�j���� {�*�-������s􎓕�=��^r��(��m�^�pyY����V"l�H��,V9V�
��tàz�-����AA99�+��8�=�gQ~��-���	��.��S!Yۅ^��Z���0�sK����������NY���;�C����tbS������w��r|�a>�����*[�|�t�Ô�|�8z8�@�}㮡�����=9XB�D�N��AA>�{�s�>2����_g�W+��650�#�aq�� ��ruZI���b@���D�AD�\R�Ѐg��`�l�0�*T)��eCl�[.sG�#b%R{�.b��|����	�`���� hK@PL>#J���7օ�w�u']9�q�Ξ���hէ3N�q,.B�y�`'AbQ�=G
z{`(%���Q�X��I��]��pN���w�+��:�%����E��$+,C���r0�a�����ϧ6Ϩ�z?�?_�Ҍ���'+�8A;gM�v���nUۜ5���C�`��7�!z�n+�3uh>���2�"*	��vѰ
k�Y��O7oB*	ڽgp��2�!��C��	��ԃ�-O�_Ȅ���a@n��&MܑN$6�-��