BZh91AY&SY<ƒp�Hߔpy����߰����  a����4       �   R� �_0      ��   @  � �]�RQU�ǅ ��� �     �p 9ֺ��[��Yb���v�e�q��=�� �dJ��vh �
�d2 R��}�A�"�P��Y$�e^�4��  � 4�]��JmI��%��D�0�EXunU�]��1Ω*��¢�*��;ۙ�v�٥%v��Sp  @ í���W�UpSZ��J�l`v��R�ek8 pc.I��p3�����:�cp�sW�w���s��@  � �V�m��j�t5{��]�(R"t�p1�o{�[gP�ઙ��vh�p��E*U�@���K�S�;5٢�*� � =� �N�]n��`՜:۹�ss��:���m"��8Z�-�s����oa��㽽ƴR�ٽgZ���    @  �U)Q)TR�  @")�      ��A��J�= �i�	���
J��	�&&�  L�����Q#j����4  @  I���"i��4204 	�I �&F�`�i��L#G�6I�����Ti�� � 4`&�4� hm�8E��%KXir\\RrH_cEE��˸EF�A� "�����)%B������U����>R�ౄ,��?h�F2�A���E%����% UQ*I�nTQ����A1%�BI$�I �_�&qGJ���z���w�^0�ޙ���GY90�w��aɜ͊ĸ䵟y\l�(������R�c��6m$å�q$хn;ʜ��ǳ��G7Q(��K:P�%��m�Ѣ��	������;�4&̮Ty%�:2X�X�J6�D�0��)8hM�O�y>A"诺djp��U���M��
؋u6���=s/<��>���v����u�UMF��l�׵+�&r�`��gM��DM��Ʌ���T�%	D����t�'�d�j�a��4q�[4"lu���Q��F�Z��k�_Vqg<ά^Ru�QT�*��*�	���>F�&��bpʖ'u�4,��Q7ܩ����UĤ�v�TYE�R�^	�jpN[u6tܜ�5\����ؔ�9iI�قhʉ߰�f�ޚ��5'��57q:l���g�飆�MK�����i�E.��c>с�{�p7�ܣ� ��J(L��P���"pF�Q��U0L;����
j}�{��BP�&��"-��f�0s�6t�:Q�$�!��;uSe����6X��N���""art��%MO�G�Q0s���:ttHܖ9#��Gd�5)�C��	���M2|�w��$���*&	�aX&cQ,饩�0ؕ&��ȍ�D�Z�h�.5,�C��$���;�K��������`���Q,�j|�j�B#]����=���iI Y���CK:5�X�e�	�p�t�*D�6#؜�Vd�:¸e��h~��樤NP���֊��Ml���tA��t�O�c��=��DKp��E0Л��Ygm+� �p��Ϩ��w⩓���n�%7��B�H5ڈ���K�J�8r%"w�#�(�B˹.58ɱ6$D�q�e�zU��S�撑2ږ&�DK�&7Q.�U��D7'M�|�$j"Q:��zʔh�6:�!�ʈUϓ��J ��>�S�uU*D��(F]L�S�֧�ɇj�uUcq�S��D����N���pG�b�,���(��TDnA2]L8o��";�Y���D���Y�5"?M��&�ʃQ�D�6u�C��DM��UD{>�j'Djt��b�u,Ќja҄�D(Fr�"hy;f�M:+D��d8U%"RA,G5T�:M͈'`��6t��%h�̕E�v�G��;DY��6%��&�Y��N�~Iҝʂ#�X�[�H�j���ҍ�)�:"]��9�	Ӄ�J��!_?D�"i�'�H�&�y+���~Y]+DM5)8"u�H쉒k�	�	� �3%&�8��#��D��҂?:����&�RA��s������$��Q��bcr�����R"tyBc�]4V�$nR%�)���_M��d�����B&��uԤDF�+��hk%|�}�U"iԧ�l�H�YT`��tzM\��~Y]+DM<��bp�J�8#����\�O���{wSǏdt%&5_Y�DЙ��P��D�*�$��nJ�GJY]6l��N	�r��㒑6/��Y������_K��q+\���F�_lM�y#��F�`�U&���TG�����UF}Cr�DwuI��Ul���ܲ���)Ԯ�q����U�A���Gb$Z�3�}�UjpM<��Ή�-et�e�D�r���2�}�h��~j�d���WȲ�S!�\�(J#����+��5_P�'��	�S]��	�C��YT��Лm�N��UGM�ʕ�M��:�Q�0х�Vu�tF�8Q�R�-ܤEԮ���_?7)V�飻�b"s�4[8QO�:#��1�p��lM;���
,~��Tj"P�"gȐn�a{gJ�{+�H��h��JDL��_#	��Mɡ4i�&�؛YT"[�H�&�U'N�n�;��{)�RG%��:;�����+�����B&͍�	ҍ,���*�L��"`�UI��M���NyK*�.�<�tge|�P�F�R�n�&n�9(�r�&�!��6"]	�7��ѫ��%��`��֒�BX��%�8py�4&���T�A�	���i�&	'J�D��f�B��D�0w¸%n|�`J�H��b]%"`�P�4k����q8h�F����4�(�':� ��NhMIY�P���.T�8#&�4��K.��K9Į8$N�j��R�g1*��~��i��M���q�\;�\:X�ߦv$�J��+g]������nHf��L�pw��%�hՒhM{+I�m�Nmehᬨ͔,9TrG5hÓF\�6�#&�4k�Dٯ��&�;�؋6Q��N	�l�'��v�6%�*��;0��R�NN���ɀ�v�eg�Bt�ϴMΏg�=�����ǰ��f�s���F�0�ϥ��<j�D�U����~�4:ʤ�crN�8'u8Q��3��=��rWMȏu+��%X��`�DG����ڈ�&�"iܯ���lGQ��ٲ��r���D�2�h��	�",��P��&wR���W�?&mܤ���&�s��R�MgepN���&;�����Y��N��[,�t��f�9���U���f�?D��y),LYX&��gײ&vU�:;�h��`A$~y*�FN�6P�ӃSЎ�P�&L�D~D�H"?r"9.��y��l�m�ʥ9��z�)}�޳���bz,�t����>���%;��lK8���f�%���&�Y!�L�������6&��L+Ü,�2���Nl8jh��u(�ýd�t���Ჾ�o�N�4^�E0��䑗'��h�k�d�T&�u܉�T沣��#��U<��Q�N�j&&�jt�̖r��>�p�]jQߓ�Q&xݭnм(�R�5��M�Pft6z�(�Bo�<���:m����K�!phP�@���l��N���1����������;�{}���.�XE��n�j�?i�[M�
�0�ܩb��'}��f��벘{7s�����\^���\��ƁH�{��p��%z�;�{)ʘ �l��l��'�NbO����7�O0ݚm��p\��͏0p3���u�a��.Vod�}�~�;|b�x�m�{��>����g{oe�tS�2_˛�������M���sy3'�uw�w{���5���1">��-�ʷ�ʱ������'�R�͞���N�ܻ����\��@h��N͜3p��ؗ�ګ6or<��u�i�M��3�T�of��'��nd���p럦�oo}�w��ϓ�$2�쫼���r~�๺������5uw�t�T��L���~�ع�D��OA�~]�0�g'�rwq�*2�M�ۗ�F[�g1O�x���۱R�����8��̼-�O�f��vչ��Wyw�ۏ��L��{s3������a/�щ�c�J�;X�Nk'o=��;~���d�ﳛ����g/}�d�^�sf�/rM��WU{$��=����žϲ��ܳ����KHD��A�x�{��\������=��>W�dg]}�Ё�;eϽ8���n̉=~�����k^��j�y���;;�U�g5>W��8s%�eKx�s=ٰ~�N���}���%�!�)��[�vpJdr�9�LUr%8��Js=<olg>]8{�P���
\�(��v&Ł��fK���78��x�;��G�����L���Yw��w�Ӊ{�X黊��W��ͻ��h�%s&��w�-X�Sʡ��(��������oY<C����|��{�^e���'��t�vi�xQ�ŸK���|��������fvi�pwv�j�OM-���9��P�;s2�o=����a��;�JG7G$�8z'�\���"�'2�{2�F;��˛�d�g�vs�˩�7�fx�a�{t���zrK;�ffn_?����0���9������gu����3ٜ�O�9�Μ�s��]�,ЛD��h�pc���gG��IV����ݻ��72ahFJ�$"�B��qM8)��׹��6�2yE�7�=���]�Ӌ��-�����z��]⌙[RpR�=ə��(|�>�ӷ�n�b|�|����h���7r��i,��������Ǖ��Ki�Ӛw=s�p_�s���s�g��l�rd!�f��gK�2�O�$��^�Wʘ)�U����ry����S�y����N{�,�4��[��L��zw�ا@��Ӽ�݀���=�;qz̳�޹q-;�f.b��Զ+9ޗ9?s�y��Է�}����=�Y_w���7��n�oF_6�s~�n��ߴ۞��o;4��bw;)ї����k��ܪsn?`KO�8��,���rLo�[�b�x፳�"�yh/q��m����,vB��	Z�o.��ӆ�����e�tng�7yy8A-���ɠw�Y�ܧB_va*&{��2�����=;{;;;������j����H`�U�7sOT���̛���MW��x�O�����X��,�fK� \�[�����9:[�8q�g��i�����s�3�N	w��?g�ܙ�OOI3֛̏��d�t �lÏ^NI��X�yd��4�--�c)���Ҝ��m�:�er��:s2Lԛ�3S�d��R�˞�޵<w��r5.s��c�70�&c�;�z�o3q-ޝ4ٜ��5ϻ��8K4���GM�������f��)m�d��q��h�x�94Q�bN���t���9��1Λ�&���Ǉ��9�{{����1��-�ٻ��<a
v�l�܅:>��
��*~	6_b����&Z{8�T��h��d�}��s�;ɝ�,���l�$�Ç'�s��G���4>�l���'b��z�٪�͐ӫ��������=�fE;�/}���e��W#��wM�'�^J̷p���M�}��g='}>��%�arwfն�ؽpu;�ԋ'��o`.g�ם�-oc�>����ѝ|;��iڳ��'s�d��:���1^s�����rN�3��n,L)����9V��g�c�;��%��o�/���>��i-�/;5��s��_L��^9���\~rC�0}��\��K6i:�ܟ���{s����[�^i�[��>JL9�sFLO�Rq��]��ow���5����}�x�ɗ�;�K@��l�5s��=���z0�Ӟ���[.�:qs_�J�\�n}��7�\f�(�c���}|�E������g&<O�G����;٣�w�e.�5��]�*���WC�㨿>��\����L���;|uu�������Y�g;��i6�-�����xDwI4Ss�����!�s�gK�=.}FS��Y)✘~Ί�=�Ls����7f=8;�̞�0�v�O�'���#�q:�w�����^�.�v�[WsM�R������o��	�6ns��/:a�-�sg˾1��ž�N�e�s���[�I�{ٸ��w������`w�״�k\`���sPzÛ�Fp�K �y8��e�;�=�Rv��촹$m�8k�[������j喛zݴ�g�͟s{��{;�7Z��*�{O �Q����7�[J�=ɹ�C�y��\�ח�Y�>$N���zr��ff�fxzқ�>�F�^���.{}�=g����|�#Ӥ����縷�ݳ��q�_X7��S�s�*���j߶���I��v[�ͳ!	y1�wss�ݜ��z�8���@�C�!��Uu���K㗜���䓆ڭ��Y��w=9���c��N�2I��+s,��^�0r�v�^�s�8p|�]Nw��3�-g��˾5��*����/\��o���8��ϖw�����ػ�V��m�n�G��s9�����w��ӗ�v�{�x�䛹�?
�����ww=6�1��﹔-�ܑN8<�~�NsV�/qNsw��p���v��{�0���m���.�|�v.����1�_�ܓ1>�^���]��rXuN��*�!9�ƹ�I���f�o1�,��s�����ݘ~xz�f���wy��Gs����Os�?)ӳ�}��ͼ.��u>s��G1�������ܓ�d���x~����w�xbY���%󼞜��qu��aIJOcJt�yٟ6aӜ��Ǎ)��O�b}��N����s;�8�߲����� ܗ�:�����뜕q����������?xHy��c�T�w��ݻi�GD�H�{ ^��nG&��p��Ic��v�F����v������u�pN��"F�h:��_��&8B*$���62��Q43��X�9�5J�蝬�:Q�%R���l��E[) �	+pc��إ�A*lc�7
Dr������~;buN��U��8Ixf3�dY%@$�$��4ŢJ
I�B�Z�N
�%%PB�O��\���gN�$���"�;�%�[�h��N�d��A8�>�+
wTT�8���a�wB��SJ~��g��&Z��H�A"�����Z�4��[�nk����(6����^`�)=N!���8l�k�[��\Dhp����m�H7]�#M��e(�H;�Ru1/���;�B��Sǃ�|���������3,�C��v�����.��ƚ��-8&�ũ�RW��nd����0UM��NSyf7��Wv��GYNE����O�`�ǋ�I5�x��x�|Q��퍢6ꂬ_UY��PA�&��7xq�N�0ܥ�Y.��Y�TV��QL���m����>�X�v��hS����%�`,}-����%`�'����`��Zbe�37LɁrF�t:9�%��q83�̝b37Ln�	sH���ރ')̴�gsF��]S���un�8԰c��~c���gg�E>��Hʥr��Jp5g5Ls����.3c7���o��MX+���7�۩��@fo�Mj�*�������<�TB��菨!c��-l�ͪ��VI�S{թ��a���y�{7�ܭ'%"�A�lݥ�k���֟7��w+!ϩ�T�p���Mkz�v�.��Q�+r�7����vh}x����,���ULeM\�B0I^bϊ�|n'�~���b��'���Y5�~����B��b2�\���o3s#V�ȣ��)b��5��
�r�("0Z��"�MX��D�0x�L�'��Ԅ�r�,��[M�l�1�18*�M����D-���iY4:O0�;��kI�/wCc�Z�Խ��|����T�?2.������&�6�f������d�&0�&w���7��Rq�c�s�2�g��=���<gPXN�!�r��ě�ͧ����&���kT!�m���~�9�c
� ����Ĵ$:5�x����6C\���T֧��bCuT��ޮ�)��]���~� r�DP�167#����_���ڮ�W������-�*�v��UꮕW�ү{�s\Uz�*�kU�Vת�Uګ�iU[X���������s��H���R����qmiUx��iU[X�����kK�^*�Ux��U������]��Ux��U��UU���[��^*�Uګ�iUS����}��H'�B}�X�����Uҫ�W��U^�UU�UU��UW��zw��U��Uz��U�UҪ�UmiUV֕W��Uv��}���I��}�߈}^���{�^�W��X��UҪ�Wj�U^�UU�UUTUW���{�\EUUEUW��U⴪��������UW��}��(`ABAa`b�I�R@I�(@Y$i���zE`BI#��ϗ�����5���a��C���\B��`s3111332�`�YӇ:'؛��e�4QN�BP�4"'�`�h�P�F&	f��%�tN�(D�DЈ����BQBh �$�lD��0D��J���un�:�:�L��ɱ!8A(DЉB"&$�A��bpM�	Ԉ�`���X�X'KÂX�hD�':pND�"lK�l��&pN�A(�'�!�{>�Q��f�?��B~��5�i�S+��"TG#����Tl�8�i�fH1����`�2��e@!�ʄ�Dm��c���[A�_��1 N;�a��>-�����
(;H�u���A@A�q�,h��G*rʆ�T�T*��꼘��"U[d�[U��+P��TR�.\������euY@ ):�@�����9
%##�QR���W򐵫('����U��)i\D��F��B*}
��U�(J�	��dj}*��t��[�A�ci�~j7G~V8�Yq<��J�l��&���.�Z�UNJ�b6+J�j}+�Bcs$W���$�R�+KH�cR��m؂&�b*���+�HK�X� "�"�"yU&;c�_��1a0��-(�n4*F�$�J����F�2�d"bm7A�_�	$7qYH��P�Q�*I#mH��-jT�
���br:�-[�E���b�����5�x�e�4&��+*m�W�����?�j�R�,U�P���Iړ���%#r*�HF�F1�I�)+ c�¬vn�,�+c�Imj'!�W$>+d!#r�WY]h����5���9�<i���Z��,�+/��2�gɪ��v�U#UX�U��i��h,�D-c+�qL��n��2����#r���Щư��6;$�O�Q	��V�j7_Կ��>1�����ߐ�Z*�U��v6�}e�5Jъ�/���}�LA��!Z�TC
�i����d-r�'ʷ6PbdQS�Dԑ
P�h�u�+rJZ:�91����2�t�jT �2}��*����9"i��T14���Eh�H�nIA�Dǘ�n�A��Ƭ��W씍��-��)cTY�D<���bt��!��m�V�F��A���`��!Se���i�V�P��i��J�fcu��ъ(�h2�),�(��D�-;�%-��Ȥ>x�'[��(��U�uQS���M�	�:�(䠝�g�P��do�#��k��S�T�Q����
��g�NFQR[��q?�1�����J*UJ눶ߪ��(Q�6�ʔL#�4���Ԛe��de��F�[Q�4G�J4��YY
��N�$��S-�?��U���ۣ��q�� "$��*�P�'֫d�VJI ;,�������j��i�T0�UGcVF�q�IZ�r��+aU,	 >����}����>��BI?}��}������|||��{���뻻����}�W��{���}��}�=�T�U�y��8��ň�Y�:"hMa�����鮡OF�i�%n��RUAV��d��
���>�f;jtV�KSCR�T!�61Z��)Zi����-�Ͳ�`#	mf&��u��
�Ie��7Pi��M�J)�>S��B�+T��#V�����+&LDy,�%��	+i�����l%���l�降��,w檍���?�+m�㉹(��P�LFXbv�J�K����n�9�u�JY~#"v䵋"2؜E
��6�SQ
���O���UR���V8v��>>��.-��k9��g{Q9����	gO�>�p/W$�8�&p���{�7���z��f[r�/���:yW�xs2�ɾ�n�a��C�n�~�y�\a�L$��y?����l�|S�!���x|h�;�nSG-�C��B�$SZ���e�V�FZ�qg��{�_a��<�&�;ճ:xMý_�&͝0�,�Y�:"hMa��Ӄ°��32����<��}5'�_}�U�Sxd;�;��p�ˍ�a�>p�'G��S��k^0�>�Bl�sRqK&�M�s�}��u�Z˺ن�sA�f�0��2�����C���l~�l<����ԃ7���0飆���(�0å�ag��Ή�:ì8�N:�}!�I$�vW%�S!��K�)�og���FapS��l��8�������b�����!�j��b�+�u��J�f
E#��|��#>S��U끸%��`j3Se@�髿�]�a�q����`{��f4y�_4�]��^Õ$�;G#5ŵo�lśa��0�0��tDК0Æ	�F�QD)��{=�}���6�,�¢�ĭ��mU���w�fh��ޫ��F�*�(�Oe��E�V��d�8l�����CF�3k��e�F$���kkNS��㞼��~��c���<4`|f�u[�5U*��ێV�i��q�uŝ�&�ц0N����YZ�n�[w+�Lk$�.Lf:	�BՑ�6��f�\NKps�Ԡ'!BJ��(4��
H���E-U%x�]�Ƿϛ��(E����B������i�{SLO�7�^�"���{c�\̹h�pÜw���c�D�K8Yz�|�{�ڼ����*#�`�Dm�&*����' w��Z8ڬ����q�@�V�z�uǚWi���x��;��ɽG����N�k}�\k��U]������yv|�B����!Ȉ���&�T�Iefm��q�q�4�N��za���Ӆ��6�S������."�������`����3ꠇ�I�g�<���������M��_�\��w�EUĬ̘�t�G7<4>��ዲD����v߄>X�JR�a�[qu&�����0�d���*4�[&�m-�m�q�q�N��:Î4㭾����t}Wƹ��:v4zXzx�|HN�DؕdQa:����G�5�m�Ǎ�s��5
|r�L�`f�~|��Q��E,qk��g���o{:jZ�y��&�YK9�ԛѰ�ӻ���˨n�Ɂ�7��V�Sfd��2��<0�6a��K���׷LQeUCM4ӯ�yǄL,��4&�0�t�(7T��I�:���P)����Z�\iR�$�2[�1/�,��8�����|��R�!�&��9[/M�����&�t�AM0��|�t+a(�w0(��Xx!���Y�!�&���S�Te��.�XWH	�G�DL<"ag؉�4b����W�68A�ۓ2X�t��v�9m����e��Ɛ>ٕ�2Kb�&�+e#��B�Kd)b�:�����~���%�Ś����g�L;�Z��	�i瘃��E��c��kbp~��[֙�=�V���S����jo�U̩�b���9M�4������w|���X�P�C��C���4 [�{�������y�OYa�)��!`z�CUND�Gp�Xs��t`y	-BI��^�W�q�eo񍶚�(���� ��ח�o2�Rɐ��鸗�J�5r�m�n>u�u�af�؉�4a���T9ҹ>kw�hf�U���s�a�JlJsףa�J�k.��r���>���:��	�ֽW�B�H������O�
v!�=�R���E�p�Q6Q%Ik{�ٗ"W��5YUh�{���U���%#$�Y�ɓ�t��MiO���m-��2�W�i,�	���x�5�a�~=/���Ɨ�~4]|�����\���<z�c2ǚ^^_�^�����yn�]y}'���y����<������y|O'�Ǜbӯ.4�2�'���y<�3��a�����y<���+�m��<�'�~u�<�L�_��Q~G��O�/))��Zy"y����k��%텼��/����by~O<����j��O��������~y���|��~~q���αח�����<��<��_����ky8�<�I�������7ry��y<�a�O/O/θǜ����<��/��mw>��������ϒ2��Z'��5�����/_����s�2<�9{��˸���?���Wgou�����6ss�����;�k}��em���]2�ë�Y8��eG]=�,�:�7��-��Ny��t}s�z�{�i����܍r�@�/^^k�X)�[����<�'�����55���W��Ւ�����}�?�������O{���뻻�3������{޻����匿����e�����Q��y�|�μ��:���y�y�]mן1��s�o)yϒI*6J
MFW$Ї�$��P�hC�h6ui(��8��?���Q��n�	*ጎS�l�R�f�[�%S�:�Ȉ�ZUr�2�H��eJI�M�6"iS�?:���sc�[��5�,���X��!@��<*���]ROzKaZ�0��O ��O`����#r	��j�u(�7�3&�D�U|�Y���K*3Ut��y҇ ɱ�����O�K�V�SC�p$�d�`���Ht�~�ļi���l��uDpXY�&�a:!��;�0��`X��u���^q�uǜy��a��u�����S��O�U���5���C�׹��MN� �%������7QB;�P�R�,Ϗ�p$�F�����-Ig��y���M�|Â�Bb�J"'�	�H�<v	��D��T��"�%~M1C/R�P�XdCg!N��,&�oʨ��`���w��[��>~X����"	�)74#M'Җ@�P\2DA{���pa22pI�ȲƠD�N�SQ�JJ�4ymk2I�)O!d�I�DHx{N�f�A��!�'#
�Gμ���~q����<�O<�/ʯ/-^_�"/��_�(LE��j��K��JdA�V��ƂѬ�4�b�۠2L�L� � � �y�@-R������I"��A֢ �i�� !G���{:!�T.qs����ӛ�pZ�S�t�Mf��������\�ÏN\�'�˯�v�/�9ȴ�[}~����D؁䌑�)�:<)4" )��i2���~"M��,�U������)dTG�U�ZkiY�\�᭽�C{���"$�&QA��1 �<�T�P>�&���ہ�!����0�0'�K&���i2��[�R���[J�%W��/J"�2���C�9�Cѓ��6"&ꔘ�	��{0�Ј���2�ŵ�p�)��.:&�vxe�c��� ����,�Btdb�!��aO�D�!=x�{�>��d�'腃'6)_���R��*���ϟ�~y��w�|��e�e�]u�^{���ĒI ���!�r�'�@� dd=]��B!��)�H�Ld����P� ��N���?Ca�!���N���D���d<H{�(�$��d�|xSIϵ���)(��C��iKL5 �+#�"v$7V��bM��MA=�;��{�P��gdME��f_��TLZ`CV!���Hq}忾�����-�_������d��l`Q��'ǥ��&�9?8pD`���偱����vtDO|��I6�	6S�&"�XR�&?����$�\��Y)wG�.�$~d���u���m�_-�y�y�]m׫*bU�R�Θ}UU����V��8'�'���e�N�tDM	8��0Ci(( �nr�A�DD
�z},WGȻ���-�`��:0�JL4"%�2N
!���܀���,�,*M��"&��~�)��4��l��=�0�y%���d�x�!���J���l�I�2GE3G���f��F���VIӰ���D��ld��D�L�|"=2�C�L���(�6$�QF�����T�8R��n�r��6CbM�Y8j�ߞR�D�7r0�=�&�&	�?om�!�QD���ø�>_��#$P���[��y�y�u��u�ߞe�d������[V1$�=����2�A�	��R���d7a�$��j��,����S����&21�Q3F
_�KmL�s[�&��'�xbc�h��:��P8XFR�����A2�4�B��!�d��h�����v��dY�C�a;�!�d��}�i9 �öNAR��F��'�W	�5�S�����=�Z���Ry>T̑:P�CIA��NH�Y���Z
w ��ՒjVD�	0a4�`��F�!�����A�'D�a�A)m�yǟ�u��mռ�4x��c���^�Z��ݛ��zUs�ȥK�\|�%V.^)��� 3�'���gN�N���ߘ�,4t,b��`�*VМ�Q�T�͒�� !.M?=����?&�W߻�Q�s99��xJsC4��[%.� ၹ7v����͌��竸
?�$[�O݇��C?+$���i�6hFT%���zy�q$���/ޯ ލ�f1[A�"Ţ"hŸ�\B�Cb+,R�J��߽��9�J�6y&��T�b�Z�y*���jJe��S�.�`M	7��AI%4%2#JCĔ;ա�C�!��	d�>a�a�2�����A��h�X'�ʔ���'�XK�d# #�@�A��R�D}��/橑�ʪr
C����̭�P!>�@�`�$6!0���_����MB��qgϜ<�n�?<�6�h��-�y�]u�Qr�}*@���i��*�0Ĥ0�dHÉ(�<�:$?�C���<3$�j�],�E��i�70Q9�A����uϤW�6S�����d@���@d���� 0�� �*}�ኦ��n:��	)�.)6�D<�(n�6D�Hr&�!����&�<�~-?+���:�XҎ��&m�F����Hv�Ij��3�bU8.�λ+��/;�#����0Ȇ��aD`TѨS"C�� �w4�m��%C�d����4PY2X4�)��m�C�p�K�j)��>�-U�IÌ4u��:���6ӧ^yo<��2뭺�%D�]$쵟.��n�����Ȕ��pn���a��(S�\�9yZ[DH��՛>:�0��(�V�6�~:3'�G����B0D��6�*2�6�*]���>��ֱgQ�(f̶�k��T��˓+MfD&�>i��S���y�r�͉�%`�#4't���ˣ{���\4��ֶKVs%�5T#8Ky�5U��)����a�W�+WQ,=��DC�'ߥ���>�a�C��<������M��G��A�@�&�6�"4�]1���2m�κ���N�~yo<��2뭺��E!����J��O"O��~����Vi�+�qB�|R��xW� �ŭ�u&��3��&)V}�߿U���U�ͫqnL5��I�Hq(��a��D1i��93H���hEԥ�cq��/5���Ȟ|˩G��q�;�a���0N��K����)�-0NFzxa��-�CF������6�*�a�5��K��m���Q�����)؈f���oȓ�	�ګm�1��bG�W����4��Y��8k�'�'�'�D�	XM��o/��m<����|�ak'�����יy���_�^�_�_�'�P�I�$��I�x)'�~q~m�q~q&���ח_�[O/�/�-�b�̯\�/���-�<��y���_��c��.x�_��0�0�0����UtT~>���|h����0�/��W<�'�c��y�<��<O�<���e�O�b~~7����c��i<W���'��y%}��V�s�4�;r|��N6�=s,���^�\O#�\��y4���~y�Ğz���~���Yĺ��'������Mb��G￑V/ϯ�K]6�F3����k������3n��	轏�yT�9�M	9ys]�l���U�uܸ��x\�5����uc������"����g�k;=��<�����&���{"���虩�~{�JS}��=�o��{':���#��sqw����T&��6w&J@:d]��>e���a��of����F��T�<��k�E n�_l��Z9����z�í�v�ٜ�\�k�����z�矲�_K~�oυCsۗ^�Oe��������9:y��%���:�.�6n,����Ļ<��ǖ�&S;7sϛ�cm�Ky�\�ɮ8/m��9��Y����-9��};�x����+OU����������p��Nl��8?��+���S^�[$��ٴ�����yI'x����c^Bi�?��;����oҩ�`�[E�%j1��Vܱ��Q��q7Y�F0���?��E���M�F~̙�Qz�Y^"�g2f�"u���7GIc������܀�F�1d� A�NEDZ,R����J�4Y�h�a�O5M7��U#UK*%s�УN)Z�?߶~ͧ����7�o���}���;��{ٙww���{����̻�xUU�fffg�*�߳339��ƞu�:�6ӧ^yo<��^^Z���'��إPq��AaF��p��jb���[e�ۤ�_�b�4' &+U�r�4|��RV�$��J�dW�D��R0pv��FD��K���@NF�Ɗ4
���$~`�r��vș\�R!�ʚ��A2;H늸�M��QF+c�g̳%vV��c�[��M9��;B�PV�#�IJ�k�8�	m��!B��#ት*O�,�Q8TV�F����ղZ���Ci��[�(��AX�ϭ�V�� 	;��ҏ��f�<g�8f�*��V(��p��&͏jk�Ն
s4��6꬏�ܵ6�B��[0��@�����<��<��h�3����4�"{�O<�Ν��o���e�U��gh�H\h�*�n�5/�����|���ه��nMA)��"��=,8tӦ�*�{߾rQ�+���������Ǚ����9�y��p,b�ӧ���f�|�K�f���?2�4ێ����6ӧ^yo<��2뭺�3uȞS��w���5_t�����D�f��:��Q/��I[8ZK/�ɷ*G�l�V6ɾ��+T�K��i��ˆ��?i1U�ilն[�p"7�K����;r��P�fB���>;��s���x3�)�M��}��r����l�~q���=6&�`��ҘYʹ�ခu�GZ9��!�s��~eם~y�\m�N�<��a�u��g��ȑ$���nD�\�֕U��?h�O��:g柳3����e�a��M6a��������ϙ��n�Z�,J�Y{���t�iC����_�7�T6���i����\ю:�[l�8>�=��U�����,��lI�p5Y��C�a�ls���5�~\�<���Ǚ���yԟ���FZG��!>�2�y�V9�6��ze��S�i�|-����qǝy��\m�N�<��a�G��eR
������Mu�ت���ȧ���7"P�@����6k�����8t�Cw��]]h�BZ0���X�Q������vL�:��t�j��V�%:w�����F�4)W�$�4!�Xa~x}�<ߧc�[��[��3$h�o���bO>��������.!��>��[{8t����̼��Ι&�~��ߤ���u)�?6ٷ?8���N�~yo<��4뭺�������Nc��U��E-�Xh�@�K��l��Erh�^�����$�jn�F��cO0O��*�m�7��V�k\�Gj"aDu��b���;%� ӑ�� 	;���?=j���fWG;0��p�]�{��f�sWW���ֽ�[���&�!I��nL$����e���>���9[1H�-_R�1�ORm��fo��]:�[]�H>���j��{�����a�{�ɔ�J����=�u��Ubd�:��uT�,���籉x�V*8�>�$�Y��c$~��Ѡ�6`t����U_�sE3U҉�ٍekO�<�|�k�N�Ɋ�㵧�m�5��}.��.m���<~0L:pA�<l�'D�<O]���U��؆�,0��s>��ۜ�s4�%=�y0�w�vŘ`(���O���!>�j�2�-��όRe?S��r�h�Vڛ;O�wܷ/��N�OA��'�ɨn`���Z�s����z�wn��Gh�Z�ipѸxos~�L:}�����$��'����g|�m���2a��zy�TO��[ƾf��9U��W��y0f���cM�q�o<���6ӧ]yo<��4뭺��F����Z�7y֙z*�!Ҍg�MڜE��!���I������g�����c���UmS4���NW~��3_S�;���%R$"!;c���E�߇!�c���|ȌMI�}���(�xt�>?}[p�5���O|^��͝_SIM�t��L����J�٨Ɩ�z���l�F6�-�u���=��׫T���y�^~q�iӮ�-�y��u�^NU�]������ �˃�8�Af2T8^`c<9ǜ�*�!��g�?O������d��u��U5I�������7I�Lefk2iZi[]�P�9MW�.���1���k��4JR��?���!vP��hc,9��^j͙.C��za��v���㐺�?v`�PL��!����g�m�Z>m���yt�S�e�|jT~�Wn��xp���y�V߻�e��B��~J�0m��u��\m�N������/-^\���ch�2��+cnH�1�]�8�n��8�$k���90��rX��C�"'s���E�O��Bi� �.z�ܜen�*�x8^J*f����^�ync|�t>��F�x�n�y�{�	M�"GN��ַ��	��K�U�ܤiƘ/�/��?]K�[��f�Fd�t�g̉��ߏ&�ѽ����~*�i��o�/��d�Gۧiš��ۆZq�CWmZ�����8��P��p��>�����ϟ!�8�jV\�%0`�������s�30Ơ����B�A��b�Ӕ��Q�['�.�O#X~1v�:CǄ��x�X��:pA<�̼�.�ۮ:���wV.��]4�UQ���7�N��.�[��Ͻir���u�q��7r�8њz�mۺ��������M�Q��\��u�S+�V����'��������6yBɉ��?��R`f��4�p[�����ڽE�1M1ګR���3N��-�ǚ�Ͳ�2����yŰt[��؞G�뒽]m�}I�5��F�_I�帙u�4�|���m����ט��O"W��&��x��4W��'�����|�,a���o1���=�3���ƒ��<a^"z�V����P�s����<�y|O>|ǜ_�/��a���;s˷�a�=�<Ǔ�/����e0�,Zx�y.y~e�<�؞_�y�<�#�=�SǗռ��\z�yu��Z����h�$yo-~b�����[��y<�ͼ���^c��W�i�x������~j�柙�����~i�<�uzv���؝_��ǖ���<������_�[�/����1o�i��z�O=s����4����O�1�<���׹�v�/��ȿ����0��]G嶖��s;g?0����/Ė(CO��5Wr��̦Nn%���v������>�|�P+ް㌔�ovn��	�������!#ڤ>��������7.�h��z\�����z�����.�H*}���87�䫙���m��{w��y\���=ȟ-�j���=&��zE��aj�ۋ׬���o?!�{�y,�^O�}G{�g���fff~��Uoٙ���UV���������~�����<p��&	�'N"CǏ<h؉���mUQC��"��r�����d�P5�_��o��zJ`��U��Hn�~ag~���s.��]O��<5���C���8BV��Y�i~�U��?$��S,}���un�6����2	�('߅X�0?I�SB���mKC���ܭ�{���i����,�M���~|�<㎶ӧ]G�y��e�����q�i}�*��`�־�U�S�:�\��:�o���=Zl��Ӛ��N�)��p�c�qƙc:.�ra�..�)�G�=k�k��̢zx���<6k����O�B�S�0�f:l?(~ؾ�P���iCr��0��I�rDi�<���a��-\�T�Z�ɺu�Xe��O?>}H��&;�C ��h��i<>:a�<'��!�Ǎ�4l�^K�t��,3CLm���j�����ł�X�ȬMkzك?��	�y81g�|#2d��cm���6��0LL�-$kL"�S�H�MQ�kq�}₃��[$--�`![Wk�� �Ź��+���� }����w��;��n�x���_ϋy�tz�a�Ӳ��U���2=�_V�r�U����wѫֻe�If^F����/���+g�b���]��7�M�ST��d˵m�&���-��߮�9\��m*y�)�}K|z���r��;��ɚu�}Zx�?W�`n��߅�R�N��h��(:>��ÇвR�����^V�t��]�wf���Qj��:}�^s��vS��dч���m��}�|��#m:���:�N�uy�^a�ǧN
bT+��UUc�������~|�F���4a��W�y�f]u��9�3��������p����_���S��������]�u��}_�!��A0G<�up�s�ɦ�;��o�ʁ�֭�D�?tQ"u�+ٓ���S�����yL2�s���a�q:�:`�)f�4IS�S�8�||�󌼏ο>~~q�[iӮ��<��2��}�2���j��UD;<�}�\�g���L���7�Dl���ۊ�L�HC�q��Ǳ3�5N3�VU�Yg�CD��_1�[��n�?C��O�o!��j�Uާ�a�V!����a4~=��f_�̹���0B��26j�n����ý�l��3�j�s�3O%i���������u��:�:��GƏ���=<�'#�[`x�V,�X��y�+	�oy�⪢XSP�q\3��u&"�P�������qb�NJ���?���ޮ0�]y̿2����|ʹ�m���9��/Wx���]�՜y�w����2��a�8�/�~��Hn�yw�"O�2��b���93LJ�ϳ�\�[v�`�-��˕YWm��v��]]6���{�q���0��%a�����y��GϘ~?�0N�D�x����Y�+D��4߅$��ۭG]"؈���ܗ,Ŗ���"8c��19!�aU�"�e���l�"?�-�XJ�W�(6��˗� !/I�&���j����=j'�<�+MsZ�>�Ӣ�B�s6c�3��L���gfrCۊ.�߼���	~,;:w�M5�|S�<(�M��C��Jֵ�ܐ���1�k�D~����SԺ2��)5U����z�|�}^j�j��]ܹ��e�Q=>����{0�!�'�o4���@�p=$�Bz�_�!���|(��b�!	5��Un	�$H��5�;����h~�{�&���w䜣�,���:xO`�8 �y�^e�mԴoXĄ$o7�ETb�ު�$��=���w1&W���Z��ʅ�[{�L��J�Sο|�i�J�3]zc�[3Z������d�Q|�����}�K��͹ԋ~v�βƤ��w�y�i�eܬ_y3̬�v�9b�$���'\�SN��w�bIO�|�qk?V_�Xa�*���_��r�q�kq�h���"a�t��$Ǎ�6x��==ߧ��e⸪&9����UD>�>2����9�"�|¹jJ��7_ϛn�3X?SUn���S$<��Q�z:��������Û��̹r�e�����-�_�F/g�k>m�j���ӎ��O����f���a���!���)�>�������]C��F���'�"	�������5l��[٧{&]yպ����㎶Ӈ]G_Ǚy��m�km]�wKl�%���2�o�wx��UT��}��x�ɍ��-�E�z�n��u�R����_˓���?���(���MlY�u��'��ç(���D;,�N�a�=ۗ�H��B���q�����O���O�UM~��)�m�E�m?o��m�����uw6hف�Q�4h��<4P�<��Wr��l���d�c�UZ�k�ۓ/��bO4�ɷ�q�'y�z���4Ǔ��u&��k�������yymxexyq<yq����c���#�4�|�+	�+�%hJ��O�(�f�+��_������4�O/�.<�_�|Ǟ_��/��+��LD�G���///�<Ǔ�/̼ǘs/1Z<���0���ˏ-�+K�5rZ�Dy#�����.GX_�/�/��y{y~O<�I�0�yq��Ǘ��~e�K~m����Ŀ�~q~|�b�y�yn���8��'��x�r���<�+$�XeO���$���&�Ǯy~O2�&�{�q�Ǘ��|�|�$aq듋_��)�O��|~2t��<���o������v�됷-2�W|?��V��}ڷh�����h�bⷸ��{���v����}���x/H�|Y����nZ�Y;�1�E�^gg���.���q1�u�{b��܌�g7��x�6�g&��K�6N��\���g�أ��5BȖ\�v�V
c��Bq4�R������fe�svAdS��H�ܝ�c4�ƶY��M�k_�E볧�Wl����e���xH}#����y�C1���sfqd���]ok�sC��a޿��]����Xv�>[��^�/ͽ[gwר��=��lPyr���Q�˙���KoJ�CM�Ǫ{�^^^ݓV�#:��Mw�����n�Í���l�O�]�7TL�h��&�;��
6�Z�le�aSp��ہl��Q� SE�uW`T��)e�O�2��PϞ6���KK�DS{iJC��9�VQ���ƫ���[_�[
16	�F���3�0m�U�TƵ��IPMW(�q8��V��1B7H��!@��q�	U���f��K��y������ޞU\�fff{ޞU\�fff{ޞU\�fff{�8x�ŉ�a�tဉ��g���W��oHI?7�)S,j�5  ����]�;h[J�n�	��j�cQ;!cJ��c����*��]uX��uE+"�H�i�X"FE$���4�V4�U��Fղ;m)$VЄj8WT����qH��+�&(Ϝ+C$j+iZr��d����R*�O���bj([e�I>%���H �rߪ,UJF&��Ye�A�qB�j+\r��- ���7K��j�~� �P�9�f[{�b��C�������w5v�O󽷼�w�x,�MB��m��u�w���x��'{է�[�3.Z����*l�h"D�ٛQ���O!���Ð�%:1XS���ɐ�1�0|����8h2	g�)���P�}��x�a�tE���4��������0�j�E>������x�y��\n��XZ�� �������s�(K�*Ϸ�lS�S�,��bn���r����N4�ϖ����q��p���2�/<�j�߿~A�q���	� !,���"0�/����??a�i=�7�������)��J	h���f��䦾�F���,��!����l���Ft��6"O��~�Z�}��7�06I�
ʋ!�
�Z80Ԛ��	w���Zۮ�]q3��70�)�qOJ�C�Olx?z�3�pC���]����VЕ��&��1��a�]mo��~y�m�����/>=8p�ѷ/V�ӈ��Y��Ӈ�UTC�ԭ���y���P��������Ȅ��-֘3M�`�&��mQ^�)�8Y�"���!��-h��%*ܖ<\-�[��މUJ����e����~}_H�3�幆6F"�C�C���5�������CSڼ�L&�~;Ŷ�i�>[l}>es8����-��+�Էi�k�4�+m�<㎶Ӈ]G]y��y֛u��U]՘J^"�TA;;���N��a�~��}�n�o�/�0m��ci���&�C�#9�������:I���8o�q�嬎e���Q)���1x�F���f2Xt�iCE8*%�=42%.�Y�]e>�om:��%z��M���0��~�;��M6�N��Ϟ~q�[iî����ʿ/,Z����U �}-v?�v�ULw갍��T�/fn:Cl�n��5V7K�n�,3[ͲWEm��(���
�-ej;��FT�v� %���v~'�	��每ו�7ƹ��9��{4"����d�seo�v�^����,�=�a������n�/f�vl$��5�b�<�e���Gܿ���f��})ã���|&���䒘	�Y���??1)�y�|�i��:kѳ���$\�rS&}�2�A�HK<u���v����Օֵ='�;M�l�&:�9)u"B�Q����UKLʙJ"��V#���a9;$������e���<�ǌ0N�0 ����g���2����WO�D�6�r��UUOFZe�3M-�S�)���1'�����h����Y-���io�MK~7N杤h��wZK�O�n�k.�v���g��em�O��]n��Z9��.WF���0�῿V��~�[��\��g
�L	|�e~��߮��o�[�����8�m8u�u��^e�[m���5��ba��*�!��C�!؛6o��3��q�l�2]��Ј���h矏ǖ�f]�i=��
�����|�a����_��r��kY�ŷMԮkZL��:�/��Jf����6�O|�?98��ҝ�����ݤb�q��D�a�BVY[�RIQ?qm?7L��Y>�%6�1L��T喒Jٵ�]am6�μ���H"h��g��,��]*�!�?�s��ne�ޚ�A?ԛ�����6MC0����f\��aU6�噆�T��I�p�j{����ո������1�9\t�>v�M��~���M^�5��!�KC�]�)���a{%8�[Z0}���&��N8ו�~]2��S4�St���^�ƹ�p�ST�U
����g��?-Ǟ~y�m������_�_���-W;��޿������Yn���\t06�n�&�F�%�>�ev�>��Za�
Y��)�g�U�9�RS�qɩ�v!;UTNL�,j ��#%V�Z��d��� JnsI|x�eB�q�w���i���u՚x�j�nb�̛y��N��9���՗�'$�6o����|~7�ٱ
~0��~U��L������!)�qu�������\�Ϛ�^���D:��h��k�帇��MS+{Q-����>{4�k1����j����)���Xa>w�3R��A4�>�q��ˬKT����tX;�����U��\_�(�@�H��tgo�ձw$�9����V���q�[iî�����/:ۭ�K��r��c
��y�~Ώ�UTA��aOO���F�p�U�QB�	qX{�o�JT���w��u#�i?ch�!������J�>2`'��5��}��r��Vl�2�M�\��5�qU�M,��֕���fAC���zw��<�4�W�2z�y�[~�_;�m�OұU�J�w6�%�c�i��e��x���dN�0N�%	�X�!�8t�8&�2h�F�AH%�: �gDK'K�:%�ӌ�%�6hC�"A4"tDN�0E �$4"'DDN4 � �A(�&�F͔C`�$��
�$�""p�QDO<l��<x��ň�aD�ı,K�Y���bX�t��f��DM6�:ai �gN���	F� �!�]t�k�<Ns�|n��n+aӶ޾�w7�,�2�؝���M�5<��<j���u����)ra��nTq��g;�3��^�_V-��������(f��:���>�c�ʗ3/x��W�.ьU�K�����߻ʘ��5y���ޜ��ة���s�e�X���]~ɝ[b�2l�v���qW��Ųx�_w�ϯ���É�4�������Z#�y��^��r�]�ܮ���̷33=�z���_�33���ʮe�33=�z���_�33�l���,�a�tဉM<l�:�����I$B~�Q+���#�Í��i4�L���Xa�ܦ%-��I4}M�6�UXn�j�u�����M���}��������8,��2�)"ymvd_౬��qib���b��q=H��+�q-x�\��.�JA���ԇ�f�j14VC�L>���\��x:zP^p�Su����[ͺ��8�m8u�u�y��m��_nݟE����]j*�������t�Tb{�:�OC!L��������}t�B�kj����csg�+���D�Z�7�e�]w?�#o��,���>��n~����P�)�'blt}������iR��N�,��kN��T��4ӨٮD�f?LF�{�g�7��ߵ1�\�������p�����j:S��<t���������	��$]^��eZd�d�T�LPY�˳�k8�sy��dG�D֭Ve����j�2GK#i�[�V�Y-N���Ɍ� K�O��/s`4_�W�us�v�w��Wm��s9������釶g����`,B_^}��a��5,,8O�"13�Ј|~��ۙ<�_�)�x�T#F�Q�ӕ���N�?a���V�7R1s-g���u�閩��&~��2��-���?S.��IS8Y�w����0��F�<<�M�� �����-��<YG�Y�D���H"hO<'D��n$��@�|UTA�����C���w�Uɇp�Rݦ���w�|���Ĵ��|{\���pɹ�~����G߮�٥��]W�#T�6�Hj��x�0�Sa�B�f�:t���0����B'v8�rF�q��}S��1ka�a<4��ձY�2a)S��q�wy]�N��7:����l.��[4��	Hޒ�R���M-���.�a��x�a�tጉM	���:&�|��X��>����U���k_����k�.LLqtlCPL2	�L������d�u�����:M�?Otn��!����i�z]�7t]کE��.\vc�<d2g:�(�9��kw_	c	�*@Y�<6f���f��bݘ��8�.��[g��/��|�٦�D?m5�_W����rz��󏜾Nm4|ul�=���o��O�i�E���0N�,D�&���%��
0�c.4�.\z���4j{�������Y����I�?vLpC�[z�L&��@a�a��R!�'!��a�����N[L1g:z�<2a�J_�.B���l�G+�^��Sm�����e���?7Z�4�$�ޡ3UZ����~,�X�"̵�^�li{��,6��ч��a�t��%��������8G���X�5����U2�Q�℩�N9��q��L0Lĸ�y@�v*�q(_�j�P����j� �z巽���ލQQ{}����a��;WV�x�r�z.��x3+��ŏ��ܒ����s�<z��j��=zd{��cNM�T��}� ��/��>2,�
�Q75���$Ⴆ�xk�-<žݜy�;L�����i%y9[�����|��pօ�!6)�C|�����ޘ ������4P���=r*�G�6HAʆ��ce��ߺ�_�����-o��u䫴i��l<p�gN�?'���(DО6|zzt�~�R)�Xcks���r�a쟩�y�YFT�v0���Fqmax���U��]~e������SRq4xX�y�=4nD1�y����Qd3�ݧZ���H���;*��Z]q,�3D`<3��-���=�I~�\��&ҵ$eq4aD���#�Şk�c�Ld
�U"�R����z�)i��[-���������0J4'��,;��Ȟl:Eq��^*��  ,�=�fW1ٳs��隓��-4�f�~���Q�k~�ȼ�Ma��f�u�9�ϪȻa��u�y��t�\�}V��k`�2��W쑖�Xj�4�u��q��W����x����]J�D�����ie���d�xvѯ��C����?sϋ6'O���b~<a�Y�0J4z|h����������]��IPt:�d�!�+���Vا���4�Ԍ�MS(�����R?6|sO����K?cX��I^7h�T)S�rO����O�ͷ�	N���ˑ.��Z���]b��Wi��WX�h]~a��ˆ���z{���67d�jSp��a�u+�T6�4��GnF��\~�x�"�l�)���������ܟ�|�F�??�tB���<'�<'�<�4�M��N��Xih�(��P�'M	bpЛ:"pL4"&d�N%	�:q'ç	���&�L8h�4PP��DЈ�0N�(A�A(�&�F͔C`�$�&J�:""' ���6x�g�<x��a���`�X�%�b%�P�&,K,K:pЂwdDN�t�0JΜO��(�DHC��N�����&�6<�O�=��g9�>���d糦w�8��3{;���ˎ�{9ż�\�	TAve;��}"-���lVs[��$�W ��<�:}@`�=��b=���qC9���;��m~�k�Z��R�Q��y��N8�.vY��Zg]Ǹ��P���ڱE�/��y��s����3ί`�l�˗.�.�a��.՘n�緱�3���w�9�N/8N�W���fI�T������C���o1��Gv����g^n���_Zމ���G�WUe�鈛���nrc}�F��������y�Ao�ݽ�X�-^���}ˆ�ݜ6�>q9�a,l��|�⢿8��>-��N�,UA�w$Q5�]�`��n&*����Y��A�Ek��GP�N�X�WT�/�g؇�el��Z��+\q;�DT����t��$
KQτMxf1�j1���K����4���ܥk�f`���m�qG�>�[����z�e߳3=�{��f_�3=�{��f_�3=�{��f_�3=�<t����%��Bx���	Մ�5J�j �n�X�ʝ�E�$��pQ�ڢ�|�J�@�4�>�5�D�+N����g��7,��!��1���Ҩ�-cؙ�ȕm2�)gѱ��M�ZA���R:�5\uT�(Y"j��YF�W%C���46X
��4E�qʣ��%*P�/ҁ)��UF+�+R9�ND�QW,�B)~n�"���[��YBڥ���"�v�n���7YD�߂2�� 	;sf�:�oM�kG���2���K�/F�Z�7{%N��s�D���y��j|V5�T���#M�긞"��2�'Gp��^�븋9ܒ�>�`kE���&�竐�����}Q��Z�5LW���3�符�N������Z3/잲?�W���rV~J��iu\�Y1��z�/͘C<B��:�[$�-P�����Am�����w�����)��o��Sr�?~��ӏ̿4��/μ�>u�V�8�θ��s���R�3�q+2K:5��DJ{
zD�8v^�(�}�|�ŵN�~�,#T+N��.��׵V�Y���(yg�u�����2�~�3QtjlcM�"aa����w�N��(��u��l"}���\LU�R����@P�4w�F��=:Ŝ�ʯ'�7Ŧ?9h�eڟ
��C��o;�h���r����i��~u��|뎓�l���ga�D�**<H<1x���V"`{p��)�Vr:lM��|"zp�=07��h��2�����i"1�仗s�K,ӧ-u��Ʌ�(��+�C������"Wμf�tn���=��>F�<��2�즸Q?C�Q4j]=O>i|�:���Wc������x�m��iL�����2�n<�����8��\u�a�^uǟ=�H��j"���O�,������껇J'��D7��+�mg42k�l2K��y���'���G�RC(�Å?5y�Y\�3n���&�"A(��?t��gN(������C!�����/�K���p��<�0N�Df������%��Ȉ��~�����]-�q�0���>p�7���N���BC��2��/��w�̗u-�Ϝi��~&�0ц�<a�����9�cCQU!����Ƨ!�?e�9#�r'��-X��:��i�b�0����S��r2Ƭui��<�P��0�I� aP�� Ģ{��� >�1�����6�፿�������u�/qsw�z`�����^(�./N욲�^�r��w�cY%&f}K�!�;���s�A0O��+?x�6�y�=]�2��W��Vbm/+C�O�iO�I�r8?.�`�}����ֿB�6
�絷����z�0NJ0p���j<�a���C���6d��I�Uh�3�41QP��8�<F�,-��x���?����a���n�`mwX_ɆS���8x�tM����ŉ�&�4a����
�xSĘ��iq�{�U��+��<�#9���h��x��̆C�
'�:{)it5�L�"|�~9X̷p��$��L�{X�..���8�7W�W�Ͷ�,�=Unih��=�&���k�9u�������.�̇f�C�Ο`��9H[�Cɩ#���(��)�a�g��Q�[���޹6�;ruūuRR�ҕ�r�F�|��Zuםq�θ�8Ì��>OJ��Պ�|�/V"$�сp������ZDn��T��2��lSQ�{�7�-w1~Iq���vֈ��q�h79Lϗ�|ޖ��f��uu3���9Ƌ�9�a��?O�a�RS��D4S[_���u�pE�a��JZ#�r�Q2�i��e�|����}�)1L0�ke���Zu��\y�:�0�.<�ϛ���H�"��Ub'�C�t�X}f�#S�y)D�ϋG�3)��	 �V����SX�"ɑJ�`�̯�О<�0OBHY5%H�*������S�:Q>�C������b�O�[/Skayf�j�i��iƑ��K���V�DJq)�w�ۍ>r-�Z<�z��q�m�L0���x�0Dц�6a�E��+���ƣ��Л�T�~gƽz��	�$�㕺I�|�Ua#9��d��̉����t�? �����~�屹�F:�S��k��9�i�}�"��K�w�k�3w���xj�7^uk>A���J%��i�ꑋi�}%���՝�u�ʍ"4�]|�(�;ש�i��NH�(�W1&R����H��4�O���k�8�:Q��r�ٳBR�����.8�`����Ƅ���Ru�4O�Ƅ��!�,�UQ
�
��'$|��]���o�>���'[��[�:'��0�b`��l��-g�`�h�>��VH�[��{�9%=��s��pИXuXkoggZq��o�=U�Z�s�^1�/u ��8tO�w'��:�W��[og�O����|��E�kG]��^K�b�B��u3�r(� �D�Y�\32�hm�z0��OBI�|_��ut�'Y�~e�H�ݶ�#���Į2Z>z�ϖ�r[�-�"E���8p؞8~?0艅	�`�uŷ�:�<��u��[/0�����D�P�4"lM2}�b`�a�0ؖ$0K�	bt�0�4CDMl��"t��M
A�H����գ�#�N�a�V�N�u(�a�(,DD�M�B&���<x�ǋ<&$%���,D���ba���bYӆ�䉱0N�'D�b`��Ή�	�`�aF� �B��g�Msom��vG�X}��?¾v)͍<y옉�sZͿE�v�N�\���NDk���=j�w2 [��˅Y�y���e������Wc���k�4|+�nW1�O���������?w�Y�����}~�\�M׻���z|�od��޹߮,�5^���?�sl���w�֗:�q�;v߹Z�;�f�%L���u��K��{��y��,�nffT�h\���w��������*�e�33�����f_�3�����\���f{d8x��ǌ8xO	���a�\yǟ=^ԒIQVku���u������$�H�>��=o�Nȉ����<�Ϝ���ޙ֖l��y�70<6I������=�S��_�ځ��DW+X��߼����yf����6[��(�a��a�e��F,8|~�0����ZQ>�O���FHCIM���ę�Z��؉̛���T�>u���R2�F����v���<hч,��<&,L4a��|x|vi%T��Ts*-���Z��U���߇PM7�&�%6P�D��9$h�Ե�{��ڛ���0��>������F��'NO�,�lF)���6h?��~O�/΄նh�!DDn��Y�D���q��6�U�.W����FV��u��a�,0�"lD秊����$䨎��ڔ�ѻ�f��>mǜ<'��ŉ�&�4a�x��_��ܧ�g�OfM�谘V���#u��cA��I��m���C�<q�`&�]��:����(�PH$)3,��E2��$��3>���>-򆭼������e����w����U����4o8���q�7��sQ�M�]�r%i~PO	����m)�Z,W��.���~�p�^&���2lͤNC��Јs�Әh�	��xP�G&�����u�L:`�g���[M�t�h�e�at�rx]8Ԝp����&��3�oۜ�J��rb�w�"�Y\�&h�6Ɵ�vM�_OO'����<�~�3�h�ݙO�`�h�_��q�_�uǟ:㮘xa�ç��G�M��J�2��P"���4��(��>��D��{��2�_��!�Z֌2��ff0����!a��?��D���D[l8�ъ�0�hrn�Ŷ�8P�����XDG9�]�p�����Tj71�-��;O ���}&GU�a����M+NR-����8b�SB|2�ϼ�gQxl���8�\q�_4��N?<�>u�]a�e��<��"��J��T�H���e�|�&�]3O���9��A�[���+�|�h�t�k�y�������".2��d0�?oB'�S}�gi��f�h�V�t]e���k�Ð���ˆ.����-���LEr�e��D��������rp���4"h!9�RQ���ޭm6���g��mS
|kK��6�4"#V92�ӕZi��m��6�θ��_:���.>y��ĺyJ���7q����UX�bS;�也B�vȜ(��g���^C�fϩ�>��7̚i�0����N��a�F	ц�]j0����EO�8rp�������Y�鰲&�~����\�̥�tM���p�2"iLRa���*��[�=�֗y~��;N-�^u�X�V��0�-4�κ'�0�bX��4a�<x�vS�UTˏ1�I�T}����c��q�e�al���V�Ғ"-���$%S�X��dr;e���X�	>�Y� �B���ӎ����!yȨ*������6��oyf��͢��lዑY�^hV�2��̼��p���<�����Ќ�)�0ay�J6��D��񆡽f�CYy
�M]p��8�f�� ����;�������~����=i�}�~�[��]w�eX{l%#�|a�`���;&j�L5ng'!�N�2��f\�X֌ŇL	��#�3R$�Nu�,8��mםq�ıBh�fx�f'�I�]��U5D�UX��tԜ���L1��YI���לe�(�a�~����7=0K�TLu�����p��L�\���cg�6�$���ZG)k��葤�~��W)�c�B���	?��v蘕�,�'2�_q.d���p��D`s��P�ֺ�ש��G�[L�L?5Ya��%�b�J>s,�?:�?:�����0�bX��4a�<x��E��h�ejV��N*�D�
z	�f�[^��t��80���vh�-h�~����.U1+���?C0D�I�����Q�� ?
�!n��8��p���5*�����u�n�J�_0�4���Ft�~]�u2���q�q�8���~��0�����t{'��<4_ҙL�tٺGX}����o�����N�S��)�����ӯ2��q��y�|��]a�e��<��%$z=)�U{�I"'�J���3b"y�Xd<�/}�q����#�&�U~��3��H�q�&0�����r�G�ܦ��?4�LT~E�D�2�naJQ�|j	�<��O1+x;U5L0WJc�&��H�߮�4�"��d=��08'Ss?;�m1�����F��T��9L��4��2ˮ���n6"`�0Lå�8!�8&6y���2������N��BP�"tM��hK�bt�,K:'��(DDK0M�htM�"A6&	�,NAB	D �	�ѣelD�L �"h0LDA6&�����Ş<a��&�"aBa�,L�ĳY"aE��ΉӅ�D���	�,��6#	�	M"��y/!�>[�!䥝����9vn�ys��B�z'�v�>�f��7sq{h.h�#޵��
��\��9y��.Ns3����'[o��)0��Q���k�y��ȯL�{��.c�'��b<���%ñE2U�����>6��\�:hk�7�V����)��xN,y������uo}�>���2�)���W!�'��>o*��r�[߽�Ͻ�o������f`le�}/O_�em���m������C�򨟎{��a睱�yv�;���H�v��=�܁�q�y����6E�Ή����y��r��w~�&�:c����������=�W3a�g�2ceH��HȎ:�'7�oW�,W�T!.U �+,%���| �χh����V�',��/�G�;���P�h��Ʌ�\��S�)[�����ϡڰLvHܭW���C���n<�BO)D�"��$m�Qɑ�V.]����uF}�^�[�r((�핦4&���RF⬊FA���\ח��_�{�[�ݷw}��O{����w}���{����ww�{����-���������<x��O%��F0�ǋ?���&z�V�,�bm��[cq2�
��$n� qY-��-#��n��P�?�P�G"���ն|�S��P
BIωm�J�:��C��dc�RU`��1���b�G�1G��K\HG)����n'�a��e��)~a	j��G���Ѩ,����l0��S���-�����b��J�!l��m@�&�Y�+��k"�#�S��7�N(�j���$�¨�mt�4a]U�CV�>jY�� �B9�2j�?;q��$���	x�a�]˾n^]�^�q�s{];��fZ�W]��l���9���6�u����h�G9{��Á�M���Xh>��J�~B��<���2�O��0��D`�����~VlD�x����3O�+8��������ܓ��|�8��˩�q��AEr7�N���G��V��@�æ�8%�:x�x�,DК0م�>:gd����1"�)z���;.�����'�%\���}�iϚ2�xƘ���M�e�m��}Ӣx0�rS>���>\mmkFG���d�|�D��M����~�u�1��b�UK_�v//���-�Wϔ�_�[d��R�����2|�KZ�N�|q�N6��֛F��Zq��N8s�͖Y��0蟄O%���2��|�k�\�����X��I"�?x��F����������4�7H�f�iyM4�4믽%}�z���|R���#��g<��R9�#�B;�}��nK��y������jd=�M	��O6xjw���<ِ������:Xh�<���K�Mu)�n��7W|�i�����)O~N�'�a���P�6X�a���D�g��L<4xt���,�ì����2��=��O4"�kե�ц��l�d��h��w|�g�Jۮ��&4uM:s}�Z#D�����ߦ���D�3����Zݟ|��Oe����e)��?S��|�a4�y��.�q��)����I!�Z?�D�+�~`�7[��֫�i~�~}'~�~3���D�ç0N��Ş,DК0Å�<Yt�*N��ַ�r|��eʕ�x��tPY�b5�c�]�2�����V�e)��}j�����MбK�B���B%�� |!~pu��5���s����6g̳D�Y�����Y7��6�9���J�'16��9��Ú���顬�\.�|]�N�?��a��;5�G'�?B�����]�!DN�\����4�	@ܧ�{"$�iiI�<�Z[LF��ĕT��~5ӆ�lOu���<º��0�RG_˹W�'���j�]�.���rn\����~��>u�o�m��'�<X��4a�<x���;G�~`*��D��L�0`���-KM���8tM�Q]C��S5�eG��4�eh�-t˝]��7'��q�N�]�z���!�D˽��w-��W%�E�VֵO��(��
�ԓ��ט�6�8��m�$�a�Ms��+GI��t���8pDN��Ş,DК0Å�<Y$�,��*$bq5+ct >���S�~u���D��8h0�Q5�DD:zo_Yo�cӞ2��3!�O��q����i�3�����O1��G���#rqE%Z�'�x��_�m�mt���i�vK�[�ϜFz�8h������=�,5H���l��<6fԛ=�0O`�v*�Ch��,��?	����"x�ň�Fp���ӆ���`T�b���~�Ub&Cg�|㣇���8z%������е���k�G[)[e��јb���6Y4r�M���%����y�t�0�}��p��b,���.��$��Ə:�;驳BjL6��~�S�s_$�,��'����ͣ/�#�o����<��ζ��Ş,�Fp�ǋ3�9�ueɒ��&Wʴh��5��sk��ĭ�3*��4CtԪV��ͲB�cv�d�;S�R;$b�| [}�_�9���s��i�x�[���x�a���xN����þ�}o#�yȟ9D̃����][������i{�1�w[޿g7���;�h}��\}�n���%u���3�헼��꿶��ݓ���h�'�����ݝ(��'d�����.��yg7���kg��'�p�S�lO!���Z��2����T�⟘��Z>[_}�5��-��Z�f0Djl��)Ȯ�[�t�3I_���'��~m����D����xM	�8Y�œ�W�/��t���\6���ؚ�L����߷߳Z>ͫ���{,=�M�tL3�ᙕ�s7��᪴4'ƙ�0���Sb%�l5�Z�Ԝ��y�g�����5�n�1�,�'M�&A���}��_(ӂg�����S-���t����(���8}$�����8줮<N�u'M�4x�D���0L�	�q�l��Zu�hˌ2�t�H���<�<�O6�ϫ2u�]d�0Ж&	���l�N��e��Ԉ��bX��P�A
�%��,D���D��ӫGY2�2�N�:v�%�J4$�4A �blM�<x�Ǐ�0���,ИlK��,тaE��ΉӅ�DN�N�gDL:pNAHP�:Q ���+S���������|��f�&�U�.ȭ�\���3� ��_ԍ��{��Z�w�{��RQy֚�M2��0H9�邶��m ܎>�������{p"�F��wh���Qԛ��v��|޿����t�z�39�E�_9�G�<,Aрq�����yܡ͐1��Xr_C	�u�|�.�i��ɘ�;��ެ�3��gf�=���u�ǹ��lq�W���7UWu��>h�����~�9˾����{�n�﾿{����y������{���������}��O0��O:x�g�a�q�y�n�̒IQ�!a�q0�䑊�6ˌ2��_��٧a���Х<���������كs&:�kY�����z3�Ƌ�~m�&�m]��p��$>��l����`���(��CG�����}m��O�Vj?e�]m$��f���I��T�+�}���Иp�:x��g�xM	�iǞ|�zconI$��+ڒ2�������W55���Xw�Ӣ���by�&����PvpMLg����iW.,5���8tMɞ��%�5>7��ţT������[N%?zI]�6�8�:Q76��D̸3a����LS�p�G!J'�O&׶��}����4�b�û���Dn��8�5���8Y��X�g�K<x��4&�0Ⴟ./��?d�$�"�
&ۈM�a�f}"�ƫC�m�.&��1���2�e��9\q�5�Yi~�U����$T>� |!E�&~�������p�#q.3�-^�ι��,DƵ{�_MzwmO6n&\��/g4�Oq�"��33�湞�����t����ְ�ov�9�~�DMK���=�И�����	��S[w��5M�ìS����u$���5���c��Lӈ�Govv^���t���w7y^r�<�����:}���jk5	�iآ%�����"���e8yg���ð�ϑ|50���Ӧ	���Y��:xM	�8x||t�Yoٟ\��-u��W)q-�V"r	�?Y4'�\��6zh(��������Eq(��a���������p��/�>8��k�o�v��}DF�y\M��0�HYv��]��H1*^5��QG]>�	񢈘YfΛ2z�����i�>97������+�_�2G���F��o�i�|��|�y��u�XqƜu��M|�$��\��Sv��G�D�Y��g�N�q��>ڙ��=�.GMQ/�BjQ���oS���0<��'�7��#��Q�ڕJ9eUK^սD33���,�<ό0D�4|k�*̹ӲQ5!�h�I���}�Z�t��y������E`l�~H����W�Y�S�?2��m�'���%�<t�Fp�<YOM\g�Ռ��j����/��ù��naǾJf�w���5nh<9$[�,��,<=��=�����CFN���v��!�	��ae��wj��^qE�S������ti��80�6��x�f�(�0M�����%çbn�iaƚu��_<돞x��4&�0�t������&�Z�V���-T�3�dشM�Lex�����
�L)\�+l6:�Q�d�90$Q��j#p�\fc5���;����o�.}��>�*�)Gg]��7��Z�bd:2���&�7;�t��~��q����{�g܎����ߟ)�ϝ��-���>�O>���&�]N��Tm?gy�~����2�1�霂xt^/�����M�a�U`/�����om�����ʆ�ll�!/~�{�#��+,�s{��fg��Ά�N�����������������i��q���:��m�u���g���g��,"�mm(��Cb��U`�C��ဘ3�x[a�s���O~�ڶ�^�}>�nv������)�)�n�l�,���8}���÷�-��5����\WZ�<���s4�OO���<��&ϧd�����t�,��e�0q�nv.�!�jL��:g�P����>8z~:�ξ~u��<��0�8ӎ��\]QeI:�e�2���N���a��q�\r�.�-�T;]e�ߒ��|����ݫ[�d�nXQ�*U]��_�mS3��<��gݶ҉�l:H���o�u��p;��u�5��aɞ��2u�����������m����Į�8�p��Y�0L0L��ag�<���8�o4��ܕE�H�UAd�=z�n���bh�z������lԧLa���t�=�vb�6IKd� F*�;!gس�o����b1��5����ZaS��1O��`��I�4�r���}ܥ30sx'�y�=������pC�Y1/3��0ͼ�|O��I�0_�*���"�{o����&M��b�>�Q�ňf�F4�%�P ��x������k�L��,Y&҇y��T"��"��*T"�"��5B��$!)A*P��B��	HD"�JB!Q!JAJ�B% �J�"�)B*)�%!(���!��%!P�JBJB*	U!(�T*UBJB)	HJ�%��!)
�����"�J!	IL�!)B!*�%�HJB*)BRP���P�BJ�TR��BRP�% ��"��%!JB!)
�JB�JB��!)UBR	H2 ��B2"0DF�E�#""� ȉ��E0D� �2�d���DQ#"�"#"DD`�����A� ���� "�F	��#DdA��b$F�2#��D`�#H���"A�ADA�����$"0D�$D�Ȉ# �"D`���0��""A"0�DdD�Ȉ#@D�$F	��F�2"DDdD�A"0D��� �`��2"#""$FDA	���"�"A�"0F1F�� Ȉ#dDFDD@B �D ����� �1���%J#�bF$�#H��$"#D`����1A"#��"0A��FDD�Ȉ#A�D�R)D�A��"%"��D�!�!��Ȉ$"Ȉ#H�`��1F�FA
�k���0D����F	� �D� ��H""2"#""2"#D�AF"#""0DD� ��DF�0D� ��`�`��`��A"1F�"	FD`#DA#"1H2""2"�F��A�20D��A"��X"�Ȉ"#""0H"$F#D""$�Ȍ��"Db$FD�#"!�#H���A�FDH��$FD@F"0H$F0D�ȉ�H2##H�"DdH #"$FDA"2"DdH$DH�"0D`�H��$F�"�F�$�"1ȉ��2"	�"2"Db$F�1 ��)DDD�A��"R �UD�A�RSQ�@FDH�DH��2"DdH #@FD@F2�"0D��F�0D`�#"$FDH�"0H$FDAȌ�0D����
$��I	$�""1
$� `���F	�
�H�V ��`,+� 2 # �n��fJ8�`���	P���"���!VBR�D$"�)��"B�!����A��A�	bBR	P�J��7A��A`���0AT�D%!	HT�"��U	D!	D"��D%R! �"�"�""��*R�T"�)A)�%�Qt�!)��dA"" �d �����!)
�% �"�"�"" �2 �2 � �A�A��"�"���*��!*��!�B��BT"	UDD! Ȃ0�T%!JB!��ʔ�BR���%T"�(�!D�2 �DA�	(��"�B��0A`�# �A!(�A(��"�R�B���%B!)
�B�	P�J�D%B!AA���A�J�JA��JB�P��BEBR�T% �B$A�	A"	QBT�!�� ��!���!R��BR�JBJB!IU�BT"��"��"2 �Ab �2 �!	U��B��"�JB*��B!*�JB�B����T��"��TBRU!)���T% B��A�D#D �!��BRBR��B��JB �	A)�5%T!��BJB��)A)�!*��� ��J�JB!��!)A)
� �!)A*���B���JAJ�!)�J������J�T%!P��� ��B�@�BR��P���%A�JB����ՕhJ�J!*��J!J!��A	HB�����!*�T��B�BR���*!*��B!)��!	HTBUB!)��P�D%T*!)���BR�B	HR ȃ"� Ȃ �D��"�"���2 �2 �2 ��P�!P�BUB�P�%T"�*�J!��`�����!*�(�B��#" �2 �� �!�T ���D"�"�`� Ȃ �	HD%!Q	UBR	HD%!��JA*��� �B�B!*��J�!)B�B!�!*	HD")Z���!*�B�P��EBR�B)�"���-	HB�	HB��%B�	HA�1A��AdAdAD �FDA��0Ab ��*���!)�A*J�A)��D%BR��R�!	HTA�"� �F �*	H!	P�J�TA*��"��JSʁ%Q�_%�cNlL��,%�J`�p>��9�Q�P@��E	@/��T+b_[
�f�,7i��qM{C�~�-���\����r�{��̼�.�u��]�0.y	��2�x����9l�MX�
/~Z���������=Z(s��3���D֔;�3�� hlEQ�T��j+��/X;��<�" ��%{��(��J��X�?����|�����`�!0��JK�)|�O�l�Eu'C��f0���;�N�܂(��=s�<����A�J��,)ߏ��o}N����,��L���"RRz��]
i��!��L9)��a[<�z]�ؒ0�/i����������B�ZY�P���"�,R
� 6������D*��(���	v-�ރ-�QFP�S`���+ہ��^�_�S`�:�@Z�"H��+�* *��"�j@PV�B��  ����&!�]\��P����1���Rz�qy��bf#���`QI�C2��U�?���@�"(��'1�a�d6���L~�2�U×�v� ���ZC �W��̏���`JqA���)��� ���|a�+z�xi�0>���&�E�uD��}�K>��W����f��>Ѐx��*P;��� ��^� �(�a��R+����;e2�S�a�_@�6�����,d���(y��@� �ލp H��L�q$��x�oR΁PTiB�x�������<��a��1?�R� �LԽpi��h����b	�/�����QF�0>22M��� N��ï�����`����<I��+��t��}a��{�07��B��)�x�yj	�=��Лǈu�=�@y�E�*Y!�{���nQ�(�5 D���+؂(�����{�=��_ 42���6�����K�����!r�2 �$X�HC����������,3`��
;�6�!rA;j��&�Hˁ۝�Y�&��l^-�l�� �(���z�U�`]%2���q�]��,+e�p�v�����0�"�D������0�Q��<c�/ӷ`�D@�����%��Ft
qO'��8�1 w��.B�@�:�)p~�0��A�1�z��S֒0�% �`1CX�?����ܑN$1�� 