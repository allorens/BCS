BZh91AY&SY���_kߔpy����߰����  aQ�|    � P     
        �                     '|�PP)AT��R�%"�ف@�� {�P��B��*��=� /��7ׯS�wv��9ݍ��ݬ�^�k�e�K6�f#�u�.Z@  �����W[kK��P�}��g���k�SId��j=�:�����P�=�Ƿ���,SG��ڍ�L��܀ �Ey j�����w�*�|8�G%$�UѤӘ�;X��`��]�nΤ�/t�̽wb]��v  0��i�}57���j��.��t�Ws�7+[f�-������[�� n CD���=*��V���k
;5���h^�s'$��JWl����D�����=�j������  ;A�>y�l}������r�6�QD�*�j6��v֑U:2�k��z��    nH�o���*���{�W�n��=ڧ��8��zRq���m^���g�ѫ� �|㈥�[L��ô�}��Cv��t옓x�/^.m��m�[Si54 = �hh������ ���z�׻��
ngM�m���v�jۧsݎю��Mve5  LJ|�������5v[f&���w;�i�Y�\t������n�Tz�W�                              DF'�R�J�  CL�  a��S�hdф ɡ�0   6JR��&�        �� J�LLa4��  ���M0T�$	�h�4�ѢO
a=CFM�I� *�A7�J�##CA`��20&&&~쟿��ާ�/[�^΃ݷ
��Yl��rq�n?H���^�:}�6l;��Fw���}�=�v�6��c�����ſg�6��6�]�������?�i���Gӥ�9�¤ù�ٛn��O��r��W�~��ٛ�����g����Ǜwʪ�����rl`=�������b�����K�O���-����8����y�����予��&5�E����"$���QNTD4��G��2�����"**�M>Zb�E"#qH�I�)�.+h�EF�LGQ�mB#���F�H��1�kB"�DGZ��(��Q��GȎi��4�1���V��"��6�"+�GZDG�DF���H�DD���|��#�wdq��z�Q���1������GB2��#h�#"�բqH�"5":�4��"">���-qF��q�b6��#(ӌ�8���}h�\DDE;[H�)�DDu��*�5h�D��GQ�[�DDG%R""�Q�:���#(�����!�Dj""9�Wh��9Q�8�*#����"4��'ՔZ4��":�;��-��#��˱բ"�"#t���"'*"4�]�DD#��Z2��#H���>�R�|���:����:�i�j8�Dq��F���G�3�DD��Fz��Y|�����[(�����v)�Q�����][(���"�q�E-z����c�DDku��U�-v:�Q������|����"-�EDDGc�ʝF�����W_-���#(ڢ"">��4�E���|�GwQH��3�)>R"7���F��b�":�qE�DDDG؈��DZ"9+���E�*""";��2��q�F�DDgUi�""8�e�Q�|��F]GɈ�Q��ҩ�sQNF�ߑ�(X�| zH��lY.'�
��ebr���FY���mu����:�H�UDDG%Q�������Z#��v����#��YE�=��-3]ELqD�E�2�����i+�DD�m�5���-�DDD�S��Q5Q�Df�����DDj�"#H���Hӌ��DDm1F�I��"#����	ڋO���j#��I]Z#mR8�QiĪ��"'�ƈMT""9*��R&�"">}���"v�6�"&kk��k'��k(@6<�zχ�����<N���8�*���>�����b)�F�ꍣ��J��2�DD�G�M*�Z�MTR#)��N��j�������{oU����<���*���������5D��:ԪDM�DI\��LDNV�D�F�Z��Սb)��U|�E��N�}�ȬDe��qO�8�8���GQqQ�T�"+uh�+���e�S��%TuL�Q�oU�q�Ti��Keo����'*�q��Du�V�>Lj�6��km:�b>u��DO�#�]DF���#��Z)�TDq;Q�SB'*Ȉ�r�.�>Rc��v�"8����b�E&j��D�|���i]E'*"'k�D�DFI�۱��2�"/�E���ָ��\���8���+��H�#����GȈ�눴F�*�%uh��j�"#��R��"�R#m&*�""7ʈ�4�DDG%|�F���������}���m��G�y�:���7U��m��DFQI]ZeO�L�D|�U�"9V���UDu�D�R""j�"#��>���%�FQ;Q�W�D�FФSi������#i���>Du�V�ȉ����U�""r�#H�Q�G�U-D�DDG%R""}QDK���G�e-7\DF[LGT��M�DF�MWYDD���i1�Du��5�Qڎ����Q�D]�Ȉ���l�.�""#�T�������ΚZ6��TGZD}uDDfTZ";�GV�"�"8���O�r�|�ꨏ��JD�DNT!���iU���W�3n.�9\eO�8��U�Gɺ���b,똎#hΛ�h��G�K��I��q��G̣z�B��-J�u�Z}]O�J㭴�]|�WT��""">�TE�5����R""7����x�����j#(�]b""#uQ�F�Lr�8��nU8��q�\��H��1�7Q|��<=���6�j�!uc����K}�cX�kZ��ʛ�9H�6r6i�4�W�Do��DD�R%TDNWȍ3����DGb��B"n�6�Rc�_3�ۍ>�q�WE��~���Q������h�)ȤGL�#����ԍGi�2��p�ڑmF��[L��GR��}Cn�u�����ƒ���Z#.�̮e1�G.�>jV(����T��DD���j8��[[i��DN�|�c��NTDi�J���4������G7Q����wJGڨ�L�}Q[m7����j�LJ��i��"2�Tt�7�DNTi�TDr�P����m5�Y�G�!�����q�I��i�ʥ��TDDG~LZ��TDGQ�٬R"#�D|��8��""7��"6�;DR"8�De�V��_"""/��[Z#Y��l�����#UQ�GU�DB3������ȍDDmbb#j�DNTG����D|��"�GQ�DDLGȊD2�DF��"����:�Z"|�GȌ��IZSL���q"&�FV��f���ۘ��R"f�"#��V-%un#��sQ*����i9Q�����"�n�i��"�Fb":�L�"";�#+D\U"":㩏�e�G���6���2�ӱ�:���u|���6�8��Z�����^ꝍ���2���#nDui��h�+m�ƛ|���Q�m�H�M������--��-�D|�:�rF�c(ˋf">�����7�|��>o�u��m�H��2�R4ӱ�{_.���a��-�b9�qͣ��ӌ�*�E�����neKs�cK���VP�9S�΢�Z��ˈ��L�ng��>j:��qg�բ:��t��"UV�;Q�SDi5Q��|�DD�Du�E&2�/KK��.�����U�)��n�|��i�q}h�E���|��F��6�>�F��h��#YE4��i*�LգP����m�ڥQ�b��B���R�V�e����ڈ˪ĪDZVj핦�H��J�m���G̭5Q;Q��&#H��DF�*�	u�mH�v��j�MմDq1Gj��#V��w*m�TG_'j:����"�U'�h�L�"�9Q�T�"�"v��qF�YVQ��YDG%|�Gn��L>���5]j��8�h��j�"#nJ��DG":�%V""#[�����DDerU"2�J�DDGϗ�E#�!��uh���n-�#(�V������Z""J�V��r�4��1U�D�DGD�FȎ#�]Z6�&�""9�f�"8����%�DB&#�������1WV�":�9\i�8����9Q�V�U�sH���Q�ZD�DDG%R|����|�E���N����2���w�랺}|�g6�W���"����+|\���+N��U�XJ�9�DIzp�7�l�����n���iY���e��Т��0\�@�u�^��V50Ϟ�����۹l��p���=�z,����^�sZ�@�Ņ?rܚ߷]�:;,�>��^��o�8���O���xٽ>���Wq���$����7[6y�2洘�4�fr���:6�����w�>o�*�{�S)I�>�ܽ%#�-��Hf�J=-����#:�v��1cC9��������/��r&D:|sF|�;ۯ@)ެ)�#`�.ێ9�	����;__�����{I'3u��s3fr��p����>wj}�m�g�����Ň�޻v��fQO�`������峒.�a���{�b��5�1�m��N-��f�%���XLҏj����x�?�e�p���(��9Fn$D�f��m��q�D��W���So��b���ћ��9����篅�z-0�{����S�Й�*�#�%`xE���c�r	�d��R��}��=�f��h�S��fj������̌(=��'t�e �v��3֏XV~�ńl ?^Do�}����ٖ�֊�fAв1���Oo�q9}�w^q�grҥ�M��ڮ9=l_�>嶱ko��H#]�7=����ɧ���w���
������y��4{��v*d������-@��e����l�.FJ�N<�eɶ�vom�Qɘ1^�Y����s��<q����m���'G���s�g{:;�$�M�H��������h����/�u|r�^o��ǎs����ۧ�̲��Ζ���/�2;y2;~��~�9�i,����{�]���g��#��=�X�79��{�yK>fLq��b׏��"9�lK�|��o�\��*��.��?>,ů�B����='e�ʿ[sb��^~��?f��>?KaR[�`˅ÇI�������݈�i��^��vF�+�~r�2�"��@���-��_�����/��%���e��!��9С�۞Xl��^��g��j-'f[�`و ���L��=�����Wv(ڏC�nv�?K`m׬���|n�m}�c^»#�3�5��W׋r����Lq�f"���C~zI����|N�xWt��+O�v��[u1���8p�Y�W��ߵ�����?O�|^����ŅIw�ٚ���γ6sg�N���ň/o��Y����^�?^�{���h��@�վV ��7F3p��<xOv��O��y�钱�q�3����¯F�yht��6��%6�������O�/�}��vy��l�v�l�=�{�
�%��y��]ݘV�!R�������|�����M$�a<��6����k�38��*�����ن�㻝�I%��喥�ܲ�kLLX����'3��/�/�����SE�V��V�x�_+;�pل�(ç�aJ*c����ϛ���;מ�%��:zv���ٷ����R:8�I����}1�9٣����8�淗�!�
�fL,���z~:A>��>{/��HDr��3�o�����k�j+�9j�?w����>>+�ׇO�o�H`3��ŝ$�ϛl�)vHSu�\tb�+O��Y|�e�4�[�f�YQ=T��e�>M�J�g�0�X^32�Z����
,�f
�����\��R�A	�b�-)륌6SR2D�dZ���o�,8g�������}�]�y���%D$�
99��L�nT��Y)�[�g�a{b�� �����3P���e���N6rG�[�JCٲ�R��IZ���m����=?Ld�.K�={����P�~�x�k��6�M�IY���[��9��"\�z�qf)�΃��w�s=��=V죡�����]���松c7L�����a�v�?�o=��hVf��1�>�!�7/8�����dk�6��G>�G�g6H��#[�b����V5�����o�oY>>>(�z�"��<��۸��=6qXI�^����q��p�}ۆŝܝ��%�,�Ӻ�M���:�#��[(��˛����4�!�13rX�� S�c7E�.���'����\���,I�I�7�w�n1������/�54�������[0���}���h/HKGD%zQ�sr��� qY��l'�­��K}�o,��cm��.�m���.2^u��ˑ����
�(����[�&�X�l�U#��-)x�x��9��$�)�=�%�k�zv�����.>=n�h����������\:���WF���b��*z��i��s�wn�Bzk�vP[���=
� UL�s�xaV^FI�ݗ���I��銜�O�T�S�Y81i���~q��f;}�B7�珠Z_g{z�Ee��9�輲����7�6l�e�/�ʶI>�m�ꍆ]�]���ED�	��;q�,���hb�eB~�Hݪ�@�0��<�#�ww�����'���p��a���kW���g�D[�y��<-�r;��<��8%��׍;�/���&M���B����oYW׻l��d�q5����;�S^#���J����D�E�A�8�<�")���q\o��Zz+�ޞ�~��vd{���[�w���v����=�|pލ��V�H/ç�<��a�δHHWa]��z����sY�}�d˳��>�Wg�J���?ZG�/�,(L�}�[��{<a��V�M[&��|��nE'8��8Ͻ��%�\N�7�3{1E����_13��~Zw>g5�L��^�}�C�����e�����\*y�%G{�~.���a��/��f�9p�����C�}����}{h��3���X}�DO�/�#ȭ�R�I9^"����wۈ<vO��������e��"����(۾�ؓ�?_qH�l���I��l��:I�}�FX�џ���ǘ�m�ْ�'q�ҞX���-��D��xc{��6���c�Gd0��g�'B����F:S?F���%<m�
EaI�L�͆���I�#6ˎNd��K�]��d�9�r�1OJ.�D�~��	����wT/����D~:p+w�K�Cݽ�sr���Ϗ�5�j7����7J�!�
ga�Qb��dS�;�e�{v�l�w�/�z1�¯Y�qL�J��.[2��7�m�<�%�xR�=�~�r����l�Eo�_�E�V>�����<@�?q5>Ev����Yܓ�e�����t[>eU����3����E^:֝�f~ύ�7�9x��1,���r'�3�w,��n��.ý�Rܟj:N�'��R(��RA���1��ǲ-ouݷd��}�	&��z��̫��������e���so�þ�o��6V��Rݱ������}׷��s��k݃�¾����/2�9&�%��5g���4�FIȤz�Z����n_YS猍�{1t����/����"��BB�qf�� ��{^��w���O)��&�Ώ�V�~2����n��1�s׏����̭�<E��\�o0�w��°�$[]����m����}���o�>ri��D����~n�߲����_�fv���=�ݪ�&^t[�'��!<u��Rù�׸�侻�f�G׶W��Sv;/1s�ooo��6��g����7�C��#�/���Tw��ݗ�[�Cq>�ge�C8��m�sXP>m�'��+��-?z��{o�՘K�U��O�ii�{q[��&[;xK�l4���\�a�8}�����U�3u�F=�ވ3��Y�8oPX�cϵ9V�e�:�d���XS�XwD�C?+�!�f���.-�W���Q�aK�bI��aj���9�,���^T�KW����_3!��o7�	<NL�y �������3w�O��v��>�_�u���Կ�_��]����7�ܼa+㌛��g[��,B�9���ѽ����Ǯ�x��w}��377���??svr��g��[;�Kₙ�\����N����������S��N��~�߿���������3w�n�w�}�o���kç�N�C�]����lmYQ�ԄkA�v��f�u�ݴ]���&��]Ԯk����k]��;.;�ڰj%���b1�l�F�ݢ2�͈�j��)�!�S�xtp�5.�vl�ª��u*�׶�9��,�S��F=����j��:���b���ę��$)1�4G-\b���.�U�f��`�`�4�p��J���LK0��$*�5�Z�ȵ ��b��2�-�v؁%�lr�]š([M,e�Jj��5�\��\6	�tƳZ��d�Mc2���L���%.\6���J�Ch���fȺ�:������M��l�dS�li�#�HU�JR��[��ʕ�(�jL�:գ5���4�bc�f��B�b�l�X��p�&������qmY�Lp�:]fn�#n��!/�z��i��mk"j��]��v�$�׷���1x1���;��bmt�s��ݴZYm��F&,V��M�d.��AI��3]m)sa\&����Qa��JRdʕ>����X|_�2�%�q@���S�w������c�<kR��:-*�E�� e#�Sie��0�����i�h�6ɻJ[n�k�Vh�v.nƣM�����븶||�u(����p�-������)umє��bAmb��pi��Gb��[l���C[CyjW4�a����Ms�s�4�.4rZKd��iZ1��������Xy�hҒ��+��0���nast�nʩ5ݣm۰�R�Q���SoWo� K�E-����[��)mld��j9Ɖ6Yog3�� ���Ṃ�j��5ʅC���IY����i�$naCR6j���Q�\F�lm�t����9��)���ؤ�Si��������MrY�~�P�I�p��uH�Y�`��Ozr[!t+(^��R���5ic_��;�\���Kv;v���E����q���n�2��B�G\BMh[��=qYm8"nR��=����S#[#$��{�$�h�@�-�&��ra���S�S��%'N/#''���0k�l)N�~��l���RZw�_7����^1��y�[��Y�eaf-e,ɵ�ɢ.����W�t��Mҁq��a�϶��+Y�m��4I�f��yθ��'Zn��iP�V�f�Y&�]S{؊�rM��sM��u�1O~��Y�-�ӲJ��tSY�(i�u�W:�#5�i6k�tU�|mNr�[[#�H�M�!�v�kB�&Ip\+wk��BjG���x�-'N���-�9:)+�aS��L	���;�:�0�5�l�H�<�����U�&W�Z�*�l+������#�J7�t��<S�e�曬���R�.�e�;p"N8����e�Y�K�1��ާW�EO�����#a`�g�ϝ}x�ڿ����Oկ��+~���3lϳ���W��u��ٛ���oOG�o��<?��]������V[ڙY�k�3F͹3m�θ5��e�j�mX�?��������h�A�⅂� [  xt�@8;��v:ɜ� �@^���� �@�<:I$��.I$��y*�Lb�Xٜ����ې�ճnF:�0�cs��mX�Y��ʪ��Z-���h;�@,ʀY�P �@��4�u�G`l4a�ִߝ ��ð8�� � ����j��g�Sf�5S5+m��Y�W�v<8d� �@pv�@l4a�4�������]
 [  ����m@�<:��@�4�V3�cY�V0�+�J��,]srī���L��S��YXV+]��oSn�umɪ��[�j�S(�;�:Z������9��b���v��;vvv�����o�6f�-��?�������������߃�?�~��~o���l�eGȍ2�QH��">|��8�GQH���)DDF��DmDFQH�뮢:���H�DF�h�DFQ�q���6���)�!�DDD|���""6���"#,��H��#h��")i�m��DZִ!H��R"#(��!B���|�#����������GYDDF��S/�>|��o�"-�DeDG�"�E"6�q�V�u�[��������Di�F��-DqDGQH����Dm��9��G�S��#���ݥ���f�v�k��s���Tݭ��,�pl�h�q6���#�2fku0�J.$pA��ke�.H#��k���ݛ�&]wH�a[Rh��^mv����N%t6��mf�
�*��u ��H��q͗�5�[�n�Z3b��	yb9��X�R)�n9�ԛSk(e� ZApL����Vm�t�GWh���X��6����ڛY��\��a���k�l���b���Kh,�D�h�Gk6�Ԋ����T��*�kX&�,L]�Ң�ZM��%��c�-�yVq�Nlܑr���k�9�8�
����[�V�m(�wa2b�J�,6+h�u)�$W!a���	eX�:R6��aճ3�I��ʬkp7BY��n�F��cY]�R$�#&cE�SB.bMsY���X�j�6�[�-fq֛k��q�l��R�]j�Z0f��X�̀��u�X��Z�m�+��̝��n����6��8.��
mse���
:�t�H�g�dc�V��n!D��#�o!)k)n5�5�����h[#n�V"�nAb�T���%�ȋ[߲z�z�ژ��p���%�]�c��&�6f�]7rm݊������V���p�k�GbW�[�JM��йd����65Y����]���b���"�}���$gz�<��։Tطv�U���I]��cv�Ae�X����
WKX�J�f����N��[Z��]�$76d�3��u����� ۘ�M3�ٛb]k�k�]��J6(1�'
��k!X�Eض��:5�TfƙΗ8"�	�����eҏzܠ�M5Eҗ��]���B��h�EΥ��09
��͘Ǝ���&,ln�#���. �Z�U�quu��KջP0Yt�`�.���� Erf��3J9єx0T�M�۵���ڄT�&�+q��ˬ)�st˳@��[WcHߥ7��Դ�5tH��6�K��cb[���s�m�t�Y&������5���M�:�E����`٘B�ͦT֭5�l7j�T����vŶ���		�z�Y����6sFbۜ��.M3�h��k�6�3�\iVYB�İ�Z�q�����M���`���UU )�{G�~��{����}o{J�c�1RK�2H��}o{Lc�b��&d�w��������1x�yR�ˮ����G]GDD|��D�)�xxZu�4�J��4���iF�PrA�+� u5�v�`�l-��@��6"���v�����@�{w�G�]n�v�e��˺��;jh�Z!�:l���5�ZRV:9Ԧ�����n5H�LT�n�v����q�8g����q�͘-m�c�f^���4�+�eaًnܧf��b�F\�$
k�l�e1e��R�`�JD�j�t��M�RE�t���@B�I2� 0}塆�>+��{2�nL�&��-�`N]����)��n�Z	���������A~�$����m��+�*���X9OHC�C��Iڣ$B��E7U��9���b���mx�Q$����1�s�����h�꼲ͭ���ϫV�ob�n�ƚi�R�|���Rz�ќ�K�f���^i��2�Н�h8�þ�N�e|�f�<m�~����<���G]GDD|�qJm�YiN��W�/]*��O��\O2/noƲ�FF���.|\�8�ۏ�\����[ �j.p����i�!U�t�����r�E2/�BM�x/N�>y�s��Ka�f�Ru�\}�F��m��l�1۷�!p���X)a6]��U��>��2���ׄ���,���<8� �mVoV���Qlu�����*�庶۪�G�k��Q�䍡u�OS�)^6�8����R:�8��"#�S�Sm2�Ju�Ֆ�\�2���I�'d�n����d�����J�v||SC�v|'����`���#<4��r��SܥϡÇC��4��5�����p��C�t��J2��ƠpF�l��<��re��9�Uy[�G����_2��۸�����k3G�6/� ��s�c��_g�(�Au��L���竾*�p�ò�k iÞ<Ļ��U�#������_2�_<��^q�QH��#����N)M�R�'����Y�\�t��"����2_�64xem'Q�Q��A���9��� G��@����Z	c�2�3�?Z3S1��tvr�:,4��>I�a=���S8�8���]k}�nז����-�a�gsi��VZ��OV>R5���4$�@�"[R�%*���Y�oh�zÀ��iHj$;!Їy��V�N9X�iU���x�$�q�g��k�8�|�:�#��u�q�DGȧ��e����U�*�H��� �-�AF�۵q���Hi��9:r;��d������Ƙ�MiƬD�6ִ6d��cjŃ-]�]�h´b�ȷe*��G:��
��$�:=��4��)������|޳G�����ƶ˱�c�7��|��m�n�ލ����2�#,6	)�p#c�h<3�R��%|xA=ǿ��"sN��^�)G4s"�e���aO�c_)U�n�Ӹ�=m��� XtH��5c�:�D�8�mO�V1��yG؋m4�V2��W~hs�/$"w�Y�d:�/2��j�F�<3^�p)�iϲAo��%�MI�(�Wiմ��g`�i��p���/���9����>��.'g��ǣ�͙%��s�~�(��:�8��u�q�DG��8iJh���=p¼s�l�3�ڌ�����|�G�8mxR2�O)N��b���Z����lm��gƍ �|�9����u��Y�^�m���NULE8�+�wTYQ���vR�<[�ng�>�4N�|��z��ۻ��ղ�F0n�Ǳ�B���0<��/�ؔ��H&��)��롚��1<P�1�^��2��U������/	�Zu�-�>qN��":��>GSm2�Juw��(�n�f��N*�S����қ�OGȩm�4z����uc�����{u+u�eϢ�����44�f����ș�B���ҊJ���E�
S�'NFUЃ�Z��m��\����	�>W�m��n���L�����}����C���ӯ�[3<8fg|9��`&��y{�SOtJ&nyd�Sr�W��\�i�E������
wUW�uL��my�����"�uDuD|�,��e��3ě>h$ŒI|�����
swY䑐���3z�703���56�$�9�!=�:$�f4v��eֺ1�K��}8�oD��|�z�	؃�O�%*�6�c���A�}a&!=4�_�2��4(v+׻�Ȭ���������C�r���!�X��UP��!�R�i�E#�?���q6�+B$��_&�;� �a��=ǛV�G_>��;�+���\|���^~|��")�Q�GQ�\u���L�ҟ#�����A�vca,[���� ���ݣ/[��Տ��͊s��xC� ������]����௙)id`��AF�F-r��1'
tq��K���q6j�EMt�����ȄW�3���m���������yݷE��9w�H%�BArE��_���$�����K�n��_l�7��;���$��0��"J����Ck>'`�[B��M {�g��vB��;2���	��x|@:G�����a�'���)�s4;s�g���7�ľ�u��\�/����;�y�>��v�)HR��t/�5���B��P�2��4�OHp;;��Ҧ���	�D`k��Mk��p=j�F'D�������7!O��Bt&oK�w�)���f�1ƵΪ���i��yN��":��㭬��e����ּ��T��u���܇�ﲜG
e�����}ʻ�1�WT�u�S�7�g�]|�9���q���>���S�.�<���J/gbA�[�M��c�h�A*�V%�K��X��/xc�)�r�	I��-�I���e��D�G�ð�-�2�0ĵ�ZǙ:���c$�c+�=^oL!���P޲�Ό��Roq�i�,\a�Msǧ!��=�?�S:z������q~~_4�T��W�Ǘ���ח�������o3�g��u}W]_ϗ�غ�������<�<�y~ym<�>y~y||�<��_�_�_�~Z����������EG�ח*������#<z����3�<�+/]WT�����y�^[J�SϮ�o.�]2�*�[ʷ��/o/���ٯ/��W��y^W�_�<Ϟ^�_�^^^�_�_�[o/�<ϕ�����׶���W�y����YyjZ��yo*�_��e��X���yZQj⢼�Z�+�ڼS���f��yKy~~y�ϗ�i_?/���_������O*��_�y�:�<�<�8���6�,�D\TE���5�k����^y�>y֞W��i��������\W�u_/�u���U�"�U��U�Wח���V?*�.ָ�ʷ��V�~g����^]<�?+*�^W��/:�>e~W�\x�<�<�=u�����6���{������iq� Y��xz�^kܦP��w^;�f��/����~a�C�@%�F�<���7�¢�������d;��!���F1ƽw~�3����s���8Z6A�	vܵ�������w���飈�[�,��z�B���39�9ɯ+RMI:��<�s�k���UI<�u$~y$�;�'��c��<����yպ�":��q�q�J[l��M������v����s���cힻ��d�d����m7�:S����[�3��<��ǅ�I��܊N3;ـ��r!���n�L��!��[sg��=&汻��׮O�[��v���t�[�6vM�nl$[n��o����ޖ�t�㾘�iL����&@�w~=O�n�'��<�_.HjG:�:����y�FFyG���	�Ї���t<;z���c&�>����������7��]�2�!A�;�2����tç��ֹ���3������F�_[�X�ʝP�c���/9;��,`&y�o����M�"V���L���#i���V@�q��L���d�c�S��k������齷�����n���4�:G��vS�U��q���e�y1fJJ�a�uf��8�&~8@ʀ<�ngũ�2��������]|�κ��\|���+)m��M6�\���H(�f�	&S���u���>��r��ߥ��{M�c���xM&���m�>��p���͜�I�V-���Q�G}:ck7�l�!���9��v�\�E�`6[Kk�����}�|7z�:Kɼ�~;>|9�8���c��w��1�1��d���h����CϺẏ���o��}y�H�[�<^3��z&qGs3P)&a�ғ�
�t���g,;ۖ��dw���^��vWm���<�;�C��ODγ����[;�S��n�\�ΒxGvn��囼remN�Ӄ�<��w�l�{s�E��6:�C�gӦ6��g=���]�>v��!�a�_�'{�a ����#N�2�u��t�Zh�������]u�7��͎�z��]���Y��AU�╈�̾y����_�[��#���y�VR�e��mN��ޏU�h��6��j\Mƍ����j�_R�Ҹ�m�F{²�2�bHn��iX���mv�\��H�,}!����K�U�\�ulb�&��JR-Z%����{�=�iM5a�˵�$܇B� ���R�3�l��Z�-������S#��P��#||�����ݲ`���PW�ф]o�	�~���˧���N�gZo:n����1ӛˣ�f��s�$Z"�� ������p?s�+l��xX�3u��9�N�����{[�vz��s��L�8�HS��0��^������A��a�C�m��xx����xM�ˍ�[>��Xʛ�bn���;��n�Zε��C�C�}[�g�t���:yq���m�Ｚ<��o���C�w�\랝��u�u���l����t�n�+6��m��t��pw۷�{����m�n��7��:Ѻ�ח9ٹ���-��єL�B`���lm��.�j2c��F��}b^6�-�wF���G��U���f�ڸ���v��d� �������A�6m��3����wl웻돚oz;L���Ke�|�����Ȏ��q�|뎼�+)m��M6�[�ՅW:��Т�8~�h�Di���h�4���n�mC�uË��@���\�-��R�M����o1��:L������u��8�D�x-�w{|��gg��89��/�[+b(�cVT3XV4�/���\�<�s�6tX$�{'P[e���}}.:��շ�����)X��~���ꘊq����X�o�c�ߩWziH�c��Ec��#�����Ȟw�6���\�@������Ff�n�&�ay˪hXM�-v�u�3u}��4�;���(�yN��z���ѭ�����.w���m�s����yAs;<:d�j�s�3
a��8~7
��ə�4�!qñG��d��u�4L���G�8����^�/:㮣ϟ:����GGθ�oR��l��n==m��ǍJ�7m'�ێ���D�K��p򟜡��?�VW�
Ŗ9�at�ګ��ڰ]]��g�W���۷g����
E0�e�;l�qٺ��0�#x��Xc$u��:�m@�39V�u�G���v!�m����.�ct�Ӯ<��ˣ·�<<����D;����?n��Ke&ږ`S�#R�_ߪ]28�2[�񪣴��!A��&v[�|G�w�۟>�\�Y�qηvݞgl��[r>-�N��G���۟oI��m�;x������St�[u�=�r:ss(~�1�1����7�`م>Qt���Q���2<���Y�W�~mӷ�7��jd�<��D�;��ԒO�L:蘃��zG����o^v��Ӻ�d;�/w�T��c�[o��_����?":�Q�GQ�:��)m�1b�/o��@!�mV���������p뻙�>���8���'D�C�0��
L��a�qa�ps�~��7�À���	oKN�?Q��2D���G`h�ҪVմ�͛�ڳN`�u��Nc��ͺym���YվT��[}zp����)�gI�ys���V}#���l�t9�q��D3��0� >����q�&���7�-t����6����-I.�;-���C��Y�M�B,�O��v���l�D;s.X@?w�~��n��ўm臛:��Nl�wϥ�:�֜Y�xG�������ݫ��gm���Vp����[Ͷ��g����n����g6��x�}NȬ|�3X���U[e�mFm�μ����?":�(�#��:�̩J[nS�p�=�:|�miI$6�	^�p٬y���Zo�MK�Mvq��섣v�+Y����u"B�`ԁFY�����.��讽L�4y��Z�:�f܂8b��`�j���7ve5ɖs�EA��?|��z 9��x�>Y=�i�}gɪ��K��Y|ϗ�����'|`%�]��oW-9���O���"�^N��ǉ�$�+gž|�ˑ�����s0Sތ���dc�R�b-����3xou]{)��V1���]��x�<��(uC�Q�~8A������^�i���a��^�Xb�g��W�2�%�Vckx�އV�S��s�'M�m��{���ݼ���z��o)�jn�pw&wt��S�����q���xz���6p�$�w���90�۵^S�-�0��Q�P��JKc��5˓�8u�G]oe���w��h�z!s30C���b��y��^[*���U�°gy	�C�}�����I4��������W�i�G^y��~Du�Q�GQ�\u��(��i��ۮ� p*
{K�3q�S�=��*,)ێ	;��t�<��\�w[xyp�7�n���q��<o.9��Ը�m�c�VݓwX�z�0�	��(@5�:�L�TNt\3��ÛI����}M�=z]o(Dgo7mr�[t���m���w���/[��%0�<�5��>ͺ��;����w�V�8�n���L泄:kn�I�7�������ޓ�yCջ'b~Wϫ��1B�l��k1�L���4��$[&hy���i0<!�ՌrZ��k35�4���U��K�������:SxJ!���Y'��[n�v�-���l�����\�KbM�"����N;{q�|��uίk�ia�v�&���E2�G��|��#��N":��㭼�KSm��juƽ�*�uq$%QEA�.xp�[�g��=X�yp���淋�Ǉ6^������)�12BdG�	�t��=�t�Q���lvH�{�7�o>��㫮����h��8�[q=�t�,ݷw0��͝޼��ޓq>�<����^k�EV1�������0��M���k%剤�a�U��y.՜���b�(����ݐ���#Ιׅ9�ۯ�%��M��\�u��&��N=O����ݖνq�O�gŴ��t�U��a�����<;7g����������s:��;�g�>�ϣ�����z�oN�*iX��q�V�-~q�~w�!B�X�]�.f����g�K�N�L�\��T�^~|��ξy��Q�qF]q��d����i�;���=N]q����R�f���3p�)8|��=J��i���D�*V�i*��R�K+2�����Mk�r���G��6�f��v���s�ǅ��7���Z8��|Mؑ���>�k����.�klH���U�K�f��N���v�����	��G3������,�8�M�B ��^���v����g�]���=�\�<O)������4��ۜ��5;��ON�m�ә��x:�>��??_��ZEh46����)�Slj����A�d:�S�T���{�������ҫ8eMS�(<Ǳx�89짵t�m�{��֛�l�N�3�^g���1.�ͻ��>��0�����WU�W���q�<����l���N��?+O/�y�y�|���^u}u�z���K�����|���<��_��y���������3痧��y^W�_�/�/����K|���"��>y�<��|��/δϞ^�_��y]W�����ު�٪�W��\yl�ʊ���o.�t�4��^U��+�y��^y}y~W��W�g��������^V�_�_�^�^�_�\yW^_�_��y���f��8�����6����QzW��WO/ʷ��4��_�~V�ũ�_��W��k�UM<�<�*��yQ��uZW�<ϕ��|y����_�R�=u�yF��^y~y~E���u�z��������?j�yy~y~y�~y~G��+����6�y~W[�W�c�-�c/-�[k�U�m�iT�W�KZ��>R�_���g��������<U��<�*�y�*<_�[ȿ_����痷�������٧�A�C���%��4	l�E}a8Ea_�Ңl�IG�+�Wy'�=�5"XE�Y�MK�o�6���EN��`�p�56�6I�����.�n$%�H$�R/��Ԇ-��0c�z�d�I���v��cF�)"��Fj��e��T�B;$zm�Cn�<r�3�_��H��p��:�X�C,�Ļ1�ƹ&>��x%��4���P�����jҜyi~��(rBJEm����lMC0��������^�i�G�a�v�(g�93.n�$�9e0��r"A%��0���ά�޵�J�Y���ѸZm�l�v�1���v1)C&~�1Ð6Q
�I���e��O4`�ް�-�f�a� ���1^e���dZ(� ˱-�8�ɍ4�MVH�m���v.�jV�.�l�zc���gI�jH.�%�mFU��q�p�x��v�B�j�#�l�oZu�|���0��:�O]����-ԣQ�`L�Jdd�Kl�Y��Eb�����ɭz2�6�[6#�Kx��u�(15mH����d��"��[�殻5�U+�2���ݵ��Z�2Jl��]�&�I��ȑR:�����\�l.!�.�l5�v�v��GZ..�[��j������WwR&��kR��-�Ci���՛��A˴iEf�GH̷,ݺ�i+��%a��ټXqD�e�"E�Vkp���0�ir1�D�u7MƘ��E���O'�1Q��gG?� ����7������wn��ُ3�}��rMI$]����*I��$�]��s\�<���Du�Q��Q�G΢�q��d����m��iR�2����>��Ɔq	f�ں��v	]l6;S[7]ۚ�2̎���V5P�dc��w���\�j4��S[�9�lUںY3U��f��[ccIU���6�=�M�Ac���JL����ڴ���qAKo.Ҏ�#X-��X���u_fѮ��ثGL̦�Yl[mڑ�BZ&�8)E��4�[@�Vm[,ż�e��J�E���d�6�'B� �/����~i��~����s��^�����f`�-#\𻻹���x�����	f4\"xD|ϧ\����<$N��p ����r���a��U�Mc/�1��ff�����WUlҊ��-�p��ͯs5V��>Yx��ʳ%m��|����\�.��������c�>'K����s���ǝvwG�c��q��bG�^ys�Ƴ׃�%��vN��ּ�xO�>�7��A=��0/gAN��-e�;0��A�;�Ss��i�.���0ZRztu�iA��z�%�GM�jM�6�U%�Hoq������ÿ8�}�U��qX����o��ݦo9ӿ����w�y��D~u�y�uDu뎶�%-���m�m�a�RU��w��R��K��k�b�X G��_�d�<i���V���O��dncx��N?wuZ~wܙ]]^3f�����k�>4�Uqռ�QB�O�wYn�2�(��։������S�Q���u�O�ò�:L�t�e۪Fj4��5�k(����c졭e�6���Oz�8����ڪ��Y��:��b	���視�ʨ=��>�Q�|a�h�忥�ŶX�:�ܴ˘�<��q�ߞ~uמy�]y�GQ��o2R�[m6�y��y219���(�u�c��|vs?���Ǵ��\C�|������=T��ÇD�ߕ���1���4�;��m��ݱ��^�>Ҕ�!�f��4:gگ�n��'8r��]�v#�b�X��j��T��ᰠC��hGԕv�����t@ ��~��~oǴ�q��dȌ�/�.Z�� ��E.ĕ~�ղ�mdſZ�H���U�l�3�.���τ�k�o"�#��W��?>q�u�y�לDu뎶�%-���m�n��^�Wx�U(�O:󝊥]|�������1�==��/ޮ��T�r�������W�嵈�Z|�5^��6xy�q�~=�Ҿ,$dI~�\7�n��nUU�+R�i��lw��}֫9�~~E�jf���d��ϜU�uJ�=���s�*�3�6+����~m��fT���D��$'��g�i'�α�0�����&�Y�묿+�N�Q��κ���"<�#��\u��C�8iÁ�l��*��n�K�+��R�z�7�o"M,7�J�)ƃʲ�fLÑ��YA��Ұ��7�fԴ��Z��9�7!�+��yK�=�c�[qi��sr˷^o�k�G T�C:ц��V��!C7j.e�7��A �@w���wnͦ�6��`�N:�j�V5`��X-b�gr�ݶ��D���Y��}�JQ��I"
C��|�U|�t�*{��Q�y��4�����+J:?�mo٪���,�U��b~����t%(L+�����������_=�Z�զ?c�u
b�Ec�&2���E1��ݙ����NI�`R���Fgy߄��C�V#|,h��;�� �����-wT��l-��n��n�3n�Յ�x�ZGΊ���w{ok)���9�e��U~~q�c���?>u���]y��q�u뎶�%-��i������f>��G9�*�)ORG
���s,�E>?|w��[���`Cj�Q�QO�뾪�>��3^�}��W1��8n���8�e����S7���:��7�{�}n�ԇG��L��PL�+�*?0�v�nu�}�L��=��$4A2?�9�����t@L���~�R�A�k}V	P��7B�u�d#�G́�s���������n�ڰ��gp{!���H�HU�ѣ�	Z,+8`�a��N��ëE���eZ����WWL߱����_��ל��O��#��κ���<��#��\u��)m��NY�I�a�(��f������:�w����i���$蠙��u�q����N�:ɪ�'㫵ez������q�xvv&��:}V��꾩�D���}�l%�lae4�-��a1�1D�Z>��d�rg
�@��=ڬ���ج,�&�j��.�׌���F93��	�V��+���)���0���x_���\�&�3��ۍ(�5������~yQ���]w��f�r,� �U������[K�EW|��`����0�S�lb�T�4����|���:���<��<�!�m�K[m��f�k�>C퀴��dPA3��hyw���-�ch���c�����ۋ�#�1 &C��wel�5��Mv��!u݆��W����q�w��8җ�z��*���8��cإҩ�����)���/����V|��[s����,)_��@��:&C�F�z���ߒ׶ߟ?ix�Y:�������?^2�)�}U+��e�%�+��m��S��z��������c����f���)�1�8ʱXoi�o���ϝG�Dy��:�m��d��,Ab������5v�mYd&�)"�䧗�O���=��%��=�e��mv�FT�ni�$kv��n��/�^}��@�Ggbeys4Е�^v��-`�v.�3$�&Ĭ��n�ͥ��8(��d<3/��gɍ�v�8��Ɇ3.m|��?�.�0�z�	�{c�i������X�3�'�n>6
<�U�������w�l��^4�ֲ���V_G�;3��:���Q�|��ϒ�ҿ}U��؏g�N�(!�A����6WFn���N��M !���2瞫Н�g�|׹O�y�3UP���>q�i��O���nu��+�;vzz#��:���V߾W��_�x��>m��Z���`&��@;������m�.Ɇ9l��[[��IM�^p5!��ٿS��[=k뺿��֢�ϛM��0�ꔥ]]?&4�o/n8�y��ϑ�y�<��u�[y���m6�ӣ��S�m�(�
)�'}'����2�����}&~CA�'��~�f��b��=�ɲ�Ţ�mX�;�z��v8Kv^S�|N�N�T�=[�h>�I!��J����#�09YU߷kS���S柙y�E9�߫�5�	���v�){|��7�oM�c�/�7��LR�)��V������O	o�<��"u�*Bc$�z���S�M1����l5��8����~[l��yי�+�m�ו���Ky����̳�g�/�������~yo<�<�>e�|���~y~Ty~q�|�+ͯ�_��m������y�]y~W�_�^�ڪ�U]m�Q���y�����������8�Ǘ痏+J�U��^u}W��^W\������]+JR�W���g��8�5��^E����W^_�_���g�_�_�^��i��^y~y~[����^y~e�b��8���8�y~yyVU���yTy�|���+L�����U�mLZ����y~U��*��O8�2�+//�Z_�_Wu����W�y����R�?/�����me���_���:_Yu����������խ~W���>y~u�|�Lڼ�2�+��ʺ�+����N���e^S�.��席+�R�E/ʶYgʶ^e꭯�/�]y}y|W�e�VV�^W��^gȿ_�_U����y���/�/�<��yu��V�~��y�������I��
ˌ�-pa�Ox�H�:fe��/��Y�Fv��q�E�=�x{5Z��/˗��/80���IYe6���^e�Xыqz�猣j���z���y{I�ك�C��$G:���ns�HW̬�����A ���s\�$��I�/Rs���@�@��9�o�y��<���#�<�#�:�<�[u��-m��m�q�U*���u۪��I�9���]�nSx���-����)U������)��(��Qd�~:�βӰA:�|77V����L�;	?f��v�.ԓ�`@�B�"�/[j7�4W��v-�~��.�Zy��~�2R��~iߺ�m�FDHx"�As9��mh��'�CX �7~(�4X�=�ܽb���������،�����)�QVDA��y�N�����F���u���<���μ�!��m�K[m��gW��r������]炊����{=J�sN2�o�i��eJSV��~�G\�إ�?�G��K]���"�#a
%vSD1�*��-�R~��BM^��S��'GE��F���B)å�J"'Ɲ�{�����ci�)J��[XգkF�io����xp�H}߆�u���w�ijR����q�[�ڟ�eJSZW*�mej���ۘ��R�S���8����ⵏ���|��:��y�y�x�N��,Ab���7��E"T_e��h�h��#[�v�����b�H`8�ĳ�'U�C7\���*'i�7��sJ��:��8AMIjk��k��7���%qY��`��T��,� ���֍���f���"���S����HA�ۋ߮O6ٟj�@��Á�
��_eLLK�;)�q�����*�`����铼���A��Q(��a
�ϰ����!��$�e؊�����0֛�H?�;?|qd�ƞ��'�b���pC��Qz��?]��c~�}�㘏׋R�2�jR����k����2�i�(����4�������S!��M:8"nI�1>����>&A?cG��EV+@
��[�-�Uj�Lê�m|������8����Lm��}v�|��'4ӌ�+U�[c_+�aלe�^u�]y�y��Dy�:��B��N0����^�PA&)�|�����y���ecm)C��ҙ3���SD�3T�=��}�m4��h����z�uQǓ��E`ƻ�3��eJ(��d�m��֒�`�F"�n�7U�^����k%���*�8����_a(i�f׈��~FJ(�3\�$#gB$!�&uť8}��p����i� ����щ2���.��;�S8ϑ�u�:�<�<�<�ȏ<u�[y���m6��>G�	J�EC��'��xJ.�`�����ġ��,�a-
QX���m�=UHҖ�(�k&�S1a�=���*m-L]�P�����jQv��ϱ�y�)�,�?ui�᱅^���殭�䧲#�%�% �NR$�]�P�@�6�����m�V�SO��q��]��������`�Bd������9��N��uw�q��Z����?�W>o�S�'�||�����g6��u�ϔo~�������V۔�H��]c�Z��u��R��q����u��G��G�x�:�2Z��ݝ��[ү�n-��JQ"%cۺ����1���y��R����c*ǅ4+P;������$d�dk]�n͍Ҕ�GIs!�0:죣����N�7�Jm��!ѧ~���jQ�߾o㮦:����g�ʺ�j��i��ӫZ�W���q.�7��v�]��}�g��\uG���)iH!Ô���{�m���oZ�;�Z��y��>S�e�\q�m�yuy�u�yy�4����C�
p�xs_����$���l�V�(�1ie���g�ُ.y�~���̤�!�%٥P-�iGjMl2��>ޱ�n�m�)Jpd{�A�&�B�R� �#���1Ĥ1nP�kS�0Z�Pȧܶ[!�}�#�G�������eﭰ4�Z�gOoI��27�<��Dw�b���ZiOu�6Mde��/z���0��_��Aq>1>λՐ��:R����o���qj5yU.��SXi�1�ǶGγjQ�]E�L�j�tC�:)}�ؖӁ�� �5�z����/L㨪�kʤÙ��0G�°AV�4O���I��յ�j��Q�~e�_/�t�6�Gqh��<�:�Lg�4���&�.�U�k���#Q�,ha��� &�X�m�v���g�c8F_8�<�|�o>y�^y�מy�y���OJA!Å8p<>�=���U\���@ �)�%p�:-��n�Zz���?*�yωW^>#J!��앖�#�a���������kQ����G�i�����b�U*a��z����(��U��c�4�qe�9��Y_�u�h�[uavFIL�����4��ѣ���}�֝�6��E6�_�]����m�c΄��)ѧP��Iñ�R�0�!��k?�����*1��m�#�������#�<y�i�V���N� ��':PD<�}��a�/��1��Xy &��CA����oVJ�ݳ����wqܑ��p��6*3����}̇����;?v~7�O{�9d){�VT��Be�&5s-��1��n�X�Y��O�[�8��n�-�J����JF��=m?<0}@�W����'κ���VKS�V-��3y��QT�1��,稥~��1��(,
�BcI]`����5���p�-cM6ˈ�/�8�����"<�<�ǚF�2�-��m�T��ͼ�u,&S��?vx�{:f�����W"��J5�i:��\�����W��ϭ6EݕdI��.ںk�#�����F����k�V�|�b�-MUW���V*�u���:�8���e��_f'N�n�x�%b�_��������Q�cR��m�$�~�__�]R�x�b�פ��	D:��7.���JLH!��HN�[>�G�d
�/c?m�mof���^+�ekqn����)����GH�2��DDi�F_>|���FQ�Di�">G�DCH���"#(���G]iu��""��DFЈ��#h��"#���!(�eH�"8�":�#(�����DE�,�DDZ6���M!���-��eH�<���T�̭��ͼ�FQ�Q��":�hB#he�|��>|��Ϟy�y"-�DF��)�|�Z:��6�1�-DeDF_"�֖�""2��h�"-�"#�E������*�V��Yy��l6r��n��M|�|ͨ	Q�ʺ`$���7�F�em��a���#P�D=[�t ^ͱ�[��جn ɇ��OVe��[��"l�M��C�����Z�EW ��~�I��dj�Z%7�}l��7���W�nݼv6�V�Bو�Z,l���='�x�K.�VE7��"�DA%_��5�{�����H\ �`����4��rx.aDi(ev[5�r6�n"�䍌����њ�Աb�l.������v�j��CE�*�.i8��El\��!2�]-˂;��ǌNN ��G��VSRb�l�+� \�ė#h���Č\��ǛŲ4l�hܻ�^h8��v����"ޞ���G ���]���,YA�,Y�-�p���ݭ%A�����)��<��6����m�i�ntֱ�m�A-3��E���f�Ů��t�����%�@��m�ɶ�oV�E���DNJF� �Ƅ�,pYp3JY�0ک��i��\��ū���W'?{�������u��YZ�2��ěIGr���`�b´*�D۬�f����Mv�Uj[X�K)��@K�	�\�	��z�й�3>�������`K�T!�����ѱ�Z� ��!4�H��fm�{�����{���s���v�ܜ�99$���I�Ns���8���<뮼���"#���iq��m��m���	��BcJ0lj��ķ[,aAg�֕W�_h�y��F�*ṨX�e�G+�Z��3[g���k�LBn	��wM�n���y��5V���dr0��5���j9.�[1kD @͎dŷm�)*�lZ���n�T��٭E��uα����[����ec�v�2n�j�+j��/1��FmoWj�&Rm�eF�h��Η^K5n2�^M��{޴����t�t�|�QA���c����旅�O^O]ܽ�R"�(���#Vi�-��E�O�!��j��\*\b]�|���~}��I ���hє�` B�B��
�(4~D������%��-nc9��4�eGb_k��m4R0_�D+o���?B|7j��5�V�]Z���(��Q��h��DA��3���&����&��k�گ��Z����c-7�uq�SE��g���M��=�M�)K[
BC\I�"�� Ć9r�>�z���9��mE3�ZwxիDFz���i��:뮣�#�"#�<��6�:)����8wϧ�XIn�$J�TR�1�e�>�|F��z�SL1l��($K��4~�M�'�@�iៅ�m�j�R:�o�"RWm����a��֦��V?+˂"�k٧�� �A�r�����C�/�cF$)%D[jA-�5�FM4)f�~;<:�~Ӈ��9N����9�p�~wU�Z���J=��cL���k~o�:r�U��Y�������[/6�<���"<�Ȏ���<�4�+R�m��uKڍ��EC��f|ts�{	�-���)D��G�+k�|���u���i���XbR���w�L�o9�m�[y���W嶥1�7�u�eh��}��5X�ڼ�J���\a�mnyh�f�4��7��Ju�3O���^��(�A<?nzoe�����W����{<�ڵu�v�yӊ5�g�I���?bwi��9	�?b�p�w�vKz4�v$]R��q��|ݝ��n�92�ڳjfJ�+f幪���ߍ��d��A3n+0��~�T��?<���:�?"<��#��<�h�l�km��۪Ms2�Q��ʣࢂ �}�$�:�3�6}�ju�SL�����`�O�忝�3���4r��qsF�H͍���i/���rp9+���ΗN����.i���KHh��cڹ��e_����Ђx��S�΍[���mDR��S�ӏeƙ[��d�}�3Ӹ��>%Ϩ��j�����'�z>��:�朠� �����t}�};V�T�o�s���aCG}��tz4��贤9���q��mu�]y�G�y�u���c�ņA�c��my�]��Lxa�=��_M�(]��5.��	0nٍJ�J^��h4������mY}���6f��UW�%�RWT�:0�j��Si�n�JJ�i��A���u5����y�qxÑ,n�ug���AK��F��WG2_���OVbS�wzN��Y`�v3v['!R+zak����""wRF������f��;���j�s�~��v|y絛��Q�]�cZʿ-�3��n�n)j)�E�]�6�x��ZǛ|��A:U�74�e<4��T]7.hX�tztt"baוf�(z�2v겧�ڬR��Z8�N�|��~�Z�ҝƱ�p��S�m)G'��4��r�hE��dݒK����#bp��3"Ǆ����Lj�w<#�{!Vj��K����P��o�6,���&(tP����^G]y�G�y�u�mp�!!Ç���m�ܽ�("	�
vi蛞7(�'�!|��'Oo<�����e�mi�eG�s?<v~�|;4�O�!��dk_��?[o�p�&�z�4�!>!�UU�c�q��-��/~�T��ju���dx6���n��RA�KLJm���e�3�O�|��o�Lq�<��J?Z��W�9�}I4�?WJ!�'���1\��Jy��L����Yn��̇�p��>|��|���#�<�΢<�ͣm������n��j����fQY��je�gVw�R��P�!�B��>us��74��f�ul�8�V�����<�H�-F�m�׌��1X��<�]��O>ƐH!�h�g�f�4�DD9��}<A��{�-���1)��l�P��MH�8�I�>0hکV8o���{&|�g����1�J�>ƛk�U�Ω\st�x���(���xir�D)�RW�gf�;�|$(�C��|�VG"�{����A�n��1!Gզ�~��I�t2�ۉ�G�Gy�^u�y�u�mm��m���u�m[M�{آ�!O1�z�sD�b��TegYWj����ܬm�J~���ß�n���|��6�E����곝5|�:�M�������8�d;Li�u_���|�e+_�x#{�������0`�AX5t��dgGXxBir�LNc�$�t|www|��;i#��zҧw7�[�rŌ~��4R	��<��LX���?4��K�<��N[�6ɯ����FI�/�K��y��	�G>ƙL)�ו�\[�뮣��<����Ȉ��6���ֶ�ZŎ�x)'�6�p�!(���a���)	qbC#)MQ��Yj�$C�D������7���kbB���F1A�RF�v��X}�Wg:�4�H���H�b�#r�+!�hD�=���m�[��}���svuJK4�R+K7dkIj��Y��3�؈#m��	���>PD'����$�\W͝0�v��W^�H�hHv�4Y�Rǃ/�$6m�1�[�Zy޲H��gΡ�w���6�(�Ng������9��w���8ps�����0D҂A��\s��|�4s�Xd �dHC����l_�Y&C���̄�pD=��.2i�(�F����~8�ɑ���u�@�����y�:���􆛟H�Y�?vvpN��2� ���U�O���JzJQ�s�ܨ���7�WJ:�Vd��ʷkYtr���w!ô���r�4��4Cs�p�������2��������i����>q���:��<����Ȉ��6���ֶ�[m����8���e�#d�Q��(���̛ۘX���\p$b�آ�&$)2��.�|���KV�F���C�}�x�����}$x͎���ov�s%��Ҕ��a��x#����:?^2CDDC�j��z��x���?�I���Ya%F���	��U�,`U��J6
�X`�nf�"+1P��7�A���H�c���]�)"�m�!�·>74s�e4H ���;���<�W�mݹ\*�[Lm���TuKQŴ�q���\��dҋ1x�ߪ��w�s��|���i��/�cV�[SO?:��*DR"�DGQŢ)DD|��O�>|㎢"#h�"6��"#�������e�F�#���:��QE#(�!2��#�Ȉ��qHB�":���8��)�����h�+DDDDDD|��(�m��kZ��meh�GF�[/:��eo<��Deu�":��-��!DDF�||�Ϛ|��/<�<��<���"-">#��E��|�l����4��>DGQ���ѥ!Ɵ""6�"-�DA������T�,s�����B�.ow9��l*�1ȵ�Y�=hK2%+���=$�[�쾵��D"- ͟�9�,��&ލ�fZ�Y�H:�)$u�@��#H�ܒz�N�X�b�8H6�����At-�Mk�R�?h�ˍ�� ����n�{��|�Nm��e�Է��bx�͕E-����$d�t�$�E*$JJ�3��j�м�:6�m�Ao��x}#�y��z�]�G9�NI;b�G9�I� �w���%r�J�����t�J�G�G�DG�y�m�V����m��)+}U*�Q����*mq+��(�l�Г _���ȘW��ۭ��Toǖ�Er�T�y���U��L�G�-��oߪ���2��g��(��ߟ̎�v]���e��ʌBG	��,ҹr�m��p�U2�-�(���[��ں��X�Z��=����6�SYT�c�y�5�e���FU�m�^cьUU1�)[6z�,�]��+zvG}���_��w�����is���*���pB�0�.3�g����8뮣��#�#�"#�<�6�+Z�mm��u���7Pwi���'0�t��E���.~ C�֐re?����/�X����$��� �]�ȃ}�k$��f������hO�0�/��Z���#M)��eY�Ww�wq��ͫ��W_INc�R-j:1N��9uY�����~ǹ�oen�|F��k~��E��l��P��G�eoͭ��<ʩ�1�^N���,���9���g�uN���s}���.�����u�yDy�y�Dy�F�ek[m���w5����9�-��O��x�f\U��獫m!��l�n�$�n&�(5�I�����@�-�˯4�+`�[�f�s�!i4�,����4��L�
>ͯ�~�@ ��{�m�v��r^e� �ӻG~|�ڶ��^&ɲ� �`r��vl��ۖ��Bл��1��G�]��)�<�/і�#.(�ex���d!����C�����.�ٟ���xs)���p3N�4��V������Rk�vt�3�O��D�����6��KE� `���7��������ʎ���z�M������,���~��8�٧6�b7���-@K�H���̸�h� �Eę	9�`��MKt��y���ӳ���/������s���ܪ��o�κ�����G�u�Dy�F�ek[m���:��X�s���E(�:ȍ#�}U���?`��"�c�g�CmM#��+��c�	����t��g=U΍��)),���L>�iG���汼~ž���qߝSyi�L���]kZ���e��:���7)�;�N��(����;Y���0Fk%�ݥ�u�������Ū��>Ɵ2ڜm�T�X�F��=��݉�]��v%N�D<Ύˆ�[��j���*�}�ҫ'R��T�b�[8���s~q�^u�<���#�:��"<���m�hC�����_z&[;Ψ.��TR�Z��V�9�]ߝs�Q��}L�Ҝ��j�(�b;��qH���j�ʔq��ǟ�8�/�gK�J"!y���RA�6�m����7t�I,���t�{�����=~|וZLS��⭢����-�/�O-�B�]��qi����Bh�xCuU+da�9�"��Ҙ˸��W����b���W�xқQ��o.�mﰷ7��R��V���Q��uWn���ƽwz8��፺��θ��Dy�G�u�yy�q�ֵ���e��ϧ���h�z(��oD)�;$����qv�Y�+�(謁�Eg��8��ut��DCz�I��l���&�`i�p�� �BKcC��FL(���!��.�3��G�C�x ��4�+��Lw���h���n'^k'���.L{�a�/q�UWV��m���g۪�U�j>ňxi��D�Ϸ��˝g�8!D��O6��V��n�qO�Z����W{~����3��e��>u���"<��μ��<��#����m��-��\#H2y�rmز�i]�g,�,�ovo����T�]m)�M�����@MBr8��92Bq�U����"m��O:U�+�!�f��Sm���Y��,�-�`�Y�v��YJTݗt�� �����b˿��9�$(.�ݻ��I>v�1��v�Y&�8V�Ij�[�\8�7�Ņ�K]��;-�10\f{�3�s�����v�6��?mag���Q���Me���TYj7�ϋ�v~G����;HY_������)��աMI]Wtï�>$����vv ����.y��Ӟv�(�oʿ��k�]�c��ʎ�Y4s���#��G���w|o�F�M���f����ꈅcM얍�|�c���捸���|�G�S���+��vZ��Le1��QǑ<��"<�<��<���m�k[g����1F_�C���qO׎;JQ�1��D�>���j�s։�~?}��C��S����3y��c�(�g\V�6ϱ�Tg����?oq�v�Ɛ
�̂A�t�a�Ӈ��t��
���ݔ�ˣXD�7lgfi����.��I��)��2?����sJ|u��Y�H���D8g�N�Y�S����v!��:?��v���W��3ڮ��7�]V��y��u��"<��μ��<��#����m��-���\�I�B��]��Ϣ�|X���r%��B+��K�W�c�v��S��#��U�R���2�:0����l�X/xy���b�I�[�j�uݽ�˶*~!�������]g�C�ᐑ���e���8�㏤�>��7��Rcg�Ǩ%��]9?6JF��߆����҈��S��^g��$;�{��Z�{���ұn���<���D~Dy�^y�y���Zֶ�p���o��um�(��("u�	���-��3����⎮�x|��)�{!�J':_~��}�u��S���`�)�Y.�S��v�Ç��8qY�-=�w5�ꮳ�i�N2��{eH��W�6�4�*��?<��7�̺��x�|	��eL��	��IX����,1��D�ޡ�����N�ni	s����6���^o%y[i��n)Mm���q�3���}�̭�~u�R"#(��4����q��":�����Ϛu�Dq�iDDGQH���D"�Dq|��Ө��eDFH�DF�D|�h��iHB���)��-DGQ|�DZքDDDDDDFP���M!����e��"Ѝ"ԏ����-�yN<�H�M��G̶�"4��m��|�ϟ6��Ϟyg�<�"#�<���-�l�|�H�u�m�b�F�DuC�Q�!�DDiDDhxxh��C��
8��ıg/j�KL��`��l�2!�aZy��q�2tv�˽-5
������Րꀹ��1���:�yȅ��|�OK'3��Jv�������31���N5 �q�,7]0n�Pl�B�wn�<*�۹vY�e��6����A!#W�˶^f/80"6�{i�'L�m��J��^�L,��q� &{raw�˝ma�99��eA�8aW��3֟���:�Z<��f`k3ٲ2ո��@�o^E�|^�N7YD�2d�-��uۓ�)����y��p��_0���&#�f+Fk��b�V}x/P�3z��z2���i�� �X�o�Y���D�b�-�q'ׂ��_�񳻭D؅)��"��X�)��R�HŘ͍+t!j�'E��>M���l0��Q�	a ӷ�Yj�135����*$�uv��,1�Jq5�Enʊf,�a$[�q,��v13vSK�#��/�y�F^�[iY��縌h���d�d����Ao�#C���0��ͩ-���Lh�c�N!�j��l����b2øn�8k��M.�&�\�-B]0K��
���Y�� ��ˢ����#jA��Q6We]b�H��v՚�n�m\Ҳ�i!��]s�tkn�.�0ݭ6j�4�<Ժ�֒�$i�m�t	u�٨uڂfa/T����K��i
5�4��= ��t���77]�8�$��MdTn�i�M�m���F�ݡUk-��is�4D��#�j��v�i���vښ�J�[����O?>-�%��IF�0��'y��{��{������~��.�T�{ܒ\����9��s<��]u��<��#�:��<��<�6�ֵ��l��ܕ�x��]kQ���Y.��ti�b�-.����v�n�MF�wk�c=�:�ā����>��O7U�P��k�
4ւ� �SM.�J�]�#j��DݞJ�[�WgJU�-)B[Ee�J��n�]�-����Vf�- PbYJK[�R��B��@�a�b˵�.Ƥ�v�e�.�!�p�i��Yh��aJSD�Q&����֚�Ck6JۜU�Ff��b�g��T�XK546S�E �}���蹌p�v��帯w�׍X���s6�^�G��h��:ÍKP�M#g�p l��X-Će�
k�Sf�~�e�uY�ӪR��Wt�|�������B�JQ9�B�G����:ӂ��U[�33����:�6s�D�p��2��"�P�:��?���[��O��ޭ<�n8�v{�v_���:�%^xC����3�:~;����=��i��]�M,�#�ku3�ջ��Ð��;�����q���1M�ſ2s��>�UU+�����Jy|����Dy�^y�G�GikZ�m�[ur�_��k0���EO�G�����gV�y~������ejek~ǽU7����Gs�'z���d�J�3x�����;U�{w|qJ���������]�'�k�߰!��Cl�}ڟ�����T�����w�0��dO��P-�q2�]t �02A�Z? ��u_�>���V�v���uM����οc��2��m�p�")�Ė�`�����\u4ۨ����u�G�u�y�y�q������e�q�cV�˖�o*Q'����w_O��yaE�-0���Ӭm�4 �.����Ӥ	�����{<���h�w���'�ǁ�}�k��*$�L��V��k"�����ia���Uy��������2�d�T�p��@�}��ł8en��.������(�T�ϯU�g_�b��>�[S�y�TJ�$EҤx`�,<Ki��)�r]_���q��^):ۨ�בבyמy����Zֶ�mN�2�q�fT�*�EG!�p��""xR�p��$�F~_�cm�k�[��)��Yu�܌��K�v�G;8@�g��go�=����3����%۩	����{��4��?e�C�Í�^�+�y�0����cu�q%_t�>��8���e�SX��ںr�U��)�9�>Rz�z՜g�i�����ã��/�F� t"~=4����pۯ8�<��G����μ����<�6�ֵ��l�������ޞIq��%\�|��Ƨ1�Xk�ڛ��rU���dWK��T+�a�m:b�I���et5����si\"��a��\�h�kQ��q��x	 ��c;�n�Xo5�k0ߔQ�CC�}��\��f�!H
y$"�f�+��c�e+#�Ο<G�<�JD~��ߖ'�㲈��3���]<��$=�ρd�}^	���c�	��\���-�����X�)g=U�m[w��S�%�M>��Ʊ���(��!�+��=���j�Gb'�L��D^κ�$�����znT��<>�uڱ��hUxC3��߯]�Sj�%�M1;O#b%Q9��lc�����0F�~2��VU*���_��u��u��u�^y�y��#���!8S��Z�fk8̒'���s��(���_-��sÎ��l�0jf}�e!%���g���2������D�j�l]LA�uݗw���-O���5�q��e��c/߉C����.�?�Q-��he}�(?�ü)�>f�d�s�N�ɐ;�z�����3]�]�tm���Sz��>�6���,��)��U�O�UwMg5L�Yl��S)����m��fy�a�h����A�n4ۮ����:�#μ���ϞGikZ�m�[u}�ׯ8�ޮUUQh@��j�"�h���A�Z�4����,-a���I3�#�|�ʻ����[��f�4T��6�Y�Ǟ�<)D<�'#��ݭ�WJ,�cbJiAE:4Ӈ�~7�>="��y����8�u�4Ϊ�n�8�iI�𾞷~�t���,ۖٞ�;.�'�7{6��ӽ��'9������Ӥ�U^��>Z׌o5*���)��T�:�~��GO-�����8����<�<����Zֶ�m��ü��j�n\�Y�ɛ�m�a�j���UX�7N�Ϯ���Z��� ���v���x.�~ "N�,�ߤ�\۠ ��.�=�ZY�~-�/���m�)�8�Ebk)E�ٶ�X�F[N�����i?���۸���G�y��"��	Q�ՠV������ A��|��U�
x"?�����z�$���v9ؓ=j��Je�2ұ��xq�u�#�먏:��#�>ym�� ��X��t�=2V�*iFB�!�n������r���
CS0c�u�G\��XT�a14I#��kE�#��B�Mt�˶
CKshXJ5%�[�m�MuֳT��M���ߕh�/�x���ȚC�l��!�v�V��2��r�{�f�n�\&-N�Z�%�x#nL�A��=A�~���S�/��u���Oz��%�/I^E�V�k�+�tI0 kt?��
�=ey$�ǧ��6|�m-���Ӳ}a�;!ó_�dO�u��!r��O35:�}k�ޝ>����x�}L�{�u,��ӱ9�g�7���'1:�v3�����CM>ǂ|"!ć�Jx{e8Q'��l���$B�$�ѠAQH�I��b�����c�ł=����Avv��ߑI��8? 8 ��G^|��#��>~y��y��)C�p��7ī��n�׊�A�fL{�UڿLm3\0F��K��Z���c*��0e�|���kBM0H@��`��I~�h������]]Tr��c�x���,Ab}R�F�����^����$v�dD��k��#6}���+q+��ϯ�[YF�GW���?3��Df!��߇���!����$��6��Ǜͅa��Ҕ���*��*��^5�)�y��p�ז�DFQ�F��8�m����8����ґDGƑ�DDu�����""��|��]G]t뮣�"""">DZ"-�F�">|�#�E�B"��FQDDe�\FQqH��hDDDDDDDF���m�""ֶЄF����DFQ�Q�#�"2�(C�)��4�6��G̣�B#H��qy�_-���>y�yO-�E:B#�4��<��)�_)�e�8�(�")F�DuG̣*B"">G��":�-D|��W4��f�_S5�x���)�E.J����N%�Y�@��������Z�4m3�\�n�mBIĸ�9� l�ԁ��س.��8Ð.�Ѕ����Q$<�G\psӽ�f_�=���/I�P�AB�#D�(�Cv�nuۢSݞ�+�q+���s�cREz�X��ER1Iܴ�zw���­���n+�ܬ�I6׹��b1Jkf�@� �Vq�l\�u�_:��Z�}�vϖ��w~�9��I.d��ʜ��$�2���No{��y�ϟ>|�8�����yyǛF�ek[m���{_UUb��\Y_c�4�-ƽ�5�=��f�)LyOqY���N�����u&+���Q�vh�7����?�p�H'?rXW%�].�vQ��
}�5�w׷y	��]VQ�q�ʹ�=��5�{�j���k�mQg��V�|���p��~oj��ו��8��5��z���Ӈ����n�dϻ:��,X�f]m_�D-�|�j�N�4�<���#�먏�y��y�m�V�8p�Zz��6r@�B`	��/�&��#���V�)�d���a�8�5���`��ţ����-�X��<�H�c���A��	��A��h��N����eA�(z��>�2~���J��C��Y�USR��ocm��p��W�s����4&wGxy`�WYL!)S�Pp'�`c�rI����Mj),ߗ�Ga���.9���^/�{��VUO�?h$�gUZ�㌴�ͺ���G]D|��<�<�ͣm2�����n���sv�k.����9�lRݬT��
&C�wgMݢ.a�h���Mc�jB�*L�v�����L�m�m���-�Kt2͖����-)+F�Ԧ��S��sd&ۢ�^(���y�a{9�����Ԙ��9	m��a��!�AZ�\�;l��	����m<��ͬÜ�#�4˰ff�8>�7<
5�|0:��J��X����DLE:*�j�r�8����Z~S��*�Q�\=d����>��uO��3�NS�ꬴ�g��ґW�}�y^}�p�b�{��UWy����i�Y��V)մ��u�s���g��h�ҭ�۩��m4n�.��Ű]m]�������'�/��	���QN�Kl���#�u�ȍ���>G�yy�� a�a8ml�~O�%��^���wO�ͼz�:��O[q�p͇��VY�}��S��[����&��R�|01�j������3I��6��x)�M9�҂xp_Nh��������%Wq�L�oC�q�zն��U_>K��6��t��tX& }�����U|��w�؏�-�f���Wq�ʥ8�جb&Yq̔�-���}T�Z��w�;l�/#ζ���^mu�<���ͼ�6�(B8C�Zo!�Ӯ*��t<1�k�)([l&�+���`�#(�i���U�Gq�s����y���&A^���UP@0wƏ�7d�i��t}��X�Qܞ�cʋr�G�svV\��y�H޳��!ׇp�ǼO0����sO���o{f띧�,�eSos�]X�=�Z��mU�+�^s��z�]���z����wuW�߸ʱ�~�Zi��S�Uv�E/Ԉ-���#�U�:�43��qw��1L�2ڜe���u�^G�<�:�#�y��y�m���8p�ߐ��O*�	���n���kU#�GJ�G����@xfX��8;�[Ȓ$Aa��X���ݫ��6.�R�xI6�ESMl����g���<�Y&-e�{��wU����S�6�Xkꭴ��~U�-0���}����m�mIu�x�d���UU�m;��H�;�?�7.CVCO����f���G��w��d�:;!�SN
fx3�����l�ӯ����#h먏�yy��F�ek[m���{��jQ��Yj-�F�,h�C%���晪�9s�|{{���y΋��e�F�l޿����1B�3oz7�����Dif!L�#kp���7b�v��XRn�[��¨��imEn�d�&��n�*�,��۴G	N�_���`���OFi=��4�p�
K�
6²G)�~c��{|$�*���A!�~�1�q��u�s�����=Y:�8�;ǋ��fݓ��ᛏA)Ί@K��Л��4�����ɽ*�b�WY|�Xk��2�aW�i��5��^�������<�J�=]��U��&���?:Yߏؼe�MU}�m���֟��K�d���
���D����xh�V;g1���F~�6�:�XP���>����n:Tb>|��ȍ���>DG��y�8iHB8C����~h���,�O��+�%w��`�D9�x����>�xn�$�ܫ�ȟ��{<8vs��(Ƨ��!b���ޜt'��y��<h�V�}�ti�?<�a�0Ӳ7�u_&&�vI��i�8����j�!\l�}�.�[�y��Vq�?o*io�����P:E��E~ʱ{Ȣ�z�f\Rr�꺫��ꩋEy帎:��Q<����>DGQ��h�!p�<;�<J����o[$�i$��Y�����?�^����f6��Չ��|��S稶�+�4ۮ�~�J�.���u�i���±�.z!	}�b~l_!eѳi�m��GYcEbK��zsk����~Լ��ULe�Qo~V+/�畤k�OI��}7FA��D���C�0���,u`������A��bF�d@�J���4��k�����oɽ)��y��h&Ĉ�`��1�1��,i��y����#��>DGQ��h�L�km��ۨ�1��0v��.UT��N���g��C�D^Ar�P4>�r��W\����F�g���D�x[�Y����طdmn�����˻n�w]�m�ۗ����,���?�X�h_�`1��!��p�~DH�F����N1VɗجeX٧�i�)�ܬl���pe~��`��ÃŠ �$ݻ��X㘩�/�|�H�WJ)�g���ԚM*�lS�;�-�b�繛��S�_��h�!�Ho��-�N8��y�Q2��"#���#H�DD|��q8�D[H�����h����DDDDu��#�u�:��"":�����F��GȎ�u�m���!H���"#H���":���Duƚi�mDDF�����eH��hB"-d�DFQh�8�FV��G���ym��">Z>RDDe�De�]u�/�8��|��y�DDu�"�e�Sμ�GV�̺��2���eDm��he���8��4������يҴ����M◘p�Y���!�0]��!<�"Q$�u�����=�V����ѥ
*!�I8N:�va�M�K�B��d�		k,�n���amcK.ɴL���Z,��;ٸ��nI1�s<�|o0r�wH�F�R%0�e��)��ĄvAM�2�eǌ�$�7�bSrY��Z��۳��F+�UHq�[� i\2 �g��b{�^�5�B!�ܲ>�=�p׈i��J������kq6,�5�=H��j@�ddW�3����M�Ze;I��l�6	���HR���ڶJ�Lz�A;�6ݳ,b��~9x֫>s�ə�G�8��iñ�F�/��O;�1����y*R��D]�EK
�b\)��!'�)F����eE�70�EǱB�� ���/��&��.{�6u��I���ǄÍ\V�\+�ܱi�"^[�7(<U$�w�ں�WSR�0�Ɖ]��+(�����n'�9��0��@�T�;oɆg�>#E�M]ħ�阁(���ǭw�^;5,�n��u�:�6�9�#��6��������`ݗ,R؆c�i�5�֘1W7u��uսi�lQ��R�.V�itci��c|=�Cx�CY�T0XLܲ�������k�]�it��̡�]�a1�b.Л;ˬ��n�~o;�Z�1Qŀ�C[�0�u�껷EՉ��h�7T�U�������i����(��ηSI�(�7M�(�qٻ\t�GM7f��k5�-�H+)v�$��g.�f룋9�L]|:�DBHZ$�
N�|���{�}�{}����^�$�@��S{��(ww���y�q�ϟ<�#��>DGQ��h�L�km��ۯ�W�O�U��܋��һƪ�l"�ݕLg\kx��Ri.�]�+GC�[�6Ьؙ���B鶼*U���fc��mC�����e�l�P�	�- �6�Ȋ^��B1:�g[�q��:�U���鮰+�A�S-�!��PéuK1`GH��릦��lj���v[�k�jm�*CB��ٚ̐f4jR:Y�':���b�s��.��E��[�9��L�b�C��U��vq��������]Ww��w���3��O��*�$�g�1�zK]�2��h߼�9��
-0ߨ|�#���R;�����>
�){�[.��x���	V�<)
c��]���|{n�~T�Ǎ��ה�8�w�ݨZ� Ay^���Zo�U�Q���Y��L�����֝���A.|��I"��gg
~;.hA<�����z4�G���w�q�VYvGjn	�X[4M	DIrf�3ǜ�v��t�ӡ�����
|���*���ߪ�z�u�>~q<�H먏��y�<�6�+Z�mbŎ�gR�y�%�$|
4	���T�D;��JR�d�AI�d�v�W�ѵ���΄����߷N<�x��}�|�նڰ;}^W=U�Zq�&����=����5���
^�tLs�w�������J&"���t�� b�M]	`�"1�5\G\dR�fgԿ=���ۜO�_V���K ��m�U]�o-�u��6�Ob�m�)�-і��<m�/S��WJ������Z�|��Q�u�4����G�SͭM-m4�m׽�V;ʪ�)>ѕ��?��`\�n�u��}h����[L���/m�[}W��z�����w~��꫼��SϞx�Uy���XF_����i��>0���v�/[��6]�Z��L�$�e�:8!p0�0̥7���}!l��l�IY�<�sR�[{o��m�b��ӈ�ls�Wv�=����6⴩�u�1�`O�$~�������5P/}i�b�*qd�QL����:ӏ�ϜG�>Diu�":�<��Z�Z�iNg� *]��Y��wڪ�#H�Z��<%xS`C �g	���	}�OMi�R�)��5�d+,�X�`l&$��OeEc>:�E
v���z�y�U4�K��4�ke0��"�|�j��iJ�;�0����.�����1/�4�3Gr\<����!وy�~�:�6�_��F�9�unr]�O������b ���N�4���L�L�u�cX���^y��#H먏��y�<�����KF�[���W��U�H�+��MH6]�I1p�T�V��h�l����n��JV���m�����@���r��h�s�k�S!\�J��ڰe���G��k*�m��X�i��b�fr$���>�I ��wэ��m��m���ݶ�?���Io��s�&8�ۼ֊X�\��N�����\�Xh����R�>ip�{4��4�VW���I2>����<� ����9����Z8|8X �m�m1٤$�|8[��`�E�8M�o�&:����]>.	�D�]��i����u�����͋�QL��>@�`�k�Bn�Y'xT����f�T�S8�R���	vh�1�ތ�	4�"�?� u�z��;��O�U���X�ʗkƚ~�q��l���u�:����>DGQ��k&���CӇ���|˳#{�U�%���u�YI�����6J�L���s4�S��O�6ѳ80?v�$�e`ښ�&!H�V(����T��4��4ixH����s�JbG:g��'Ee��dm`�m��&�eղ(�_r[����g�)�3N:0�N�q�P��t"7��.i�q4=4����s���c֏����J����Т�00tֳE9�o8��|���y�u�q�y�<�����Ku�qB��>�ڶ�1�g�՘뷯5('��C&Rd����ϛae���W1e9��)��J����c*��wz}�ږ���/*���+u[�m��S���u���Ռ`{�Rw���Z�;Ⱥ1",�"���T�a%�Y��̜<':";�n'�`�\��>�ec���|E��U=�V���:�V���?���|<�I�TpO�%�����`XZ<�(�����Zu�bV1��y��kk_�}������T��m�CN#o�<����:�8���<��mJiki��ۮm�c>���n�s��TN�Y�S��F�i`�ͩx�/w��nz���t?#ݭ��m�5k
�FH�8�٨�o�rc$NJttxS��V�8d4��{���)x�Z{5�s֟��|S�Z�Z4�q۫���R��?k}ey�=�]SkGp�N6��j���b�Ug�R�y��WU-U{6R=�*��O�b��Ŗ?
��U��ki������� @����m���1�)�#����euDDuy嶥4����p����"��ٵ�1\��^KT��E��=}����4���+S�0G%0KQr�ݤ[�Q!����)|Qf�Û�+m�6m���˅��Cf���=p���n���ŷ�sRJe,���&����j�'��u���{�u����~�sr���{
���i"�l�nH3D���gn��Px]�W��~�JtA�8���G8i�Ϥ�� �ށ�Ƅ<s͑��}��2[�������;�!�B�߉�� C+k)��0J�`<Lc��	��ʊe��iߚev[�x�s�Uf']M6j]����}�᠞�74�=�3(S^ؿd�I�el�l�M��f��Lj�M��9�����ec4��74T44���L:��tҟ�]Sͼ�(��#�-uDDuy嶥4����m��������U=��O��Yڡӷ��I~�dãsre7��@�V�B�{�Rd~h7�xD]Z$�V�Q��++A��޲S.�/�%��\RhC������t#�h.��!�{�e�jW	-6�b��6�I�#~
xhܖ�fn�s�NT9��[x�kZ���[���6�>�~�0}p��3~)|.��X�e���䫪�]��[q�IV��u���庅">eDG��FQ�D|���G�qDG�"""2����4����"�:�""#�\DR"8���-��h��u�GͶ�R�E""#���""#H���#(�4�(��2�h���|���H�m���Z��E"2���DFQ�Q�>B8�����u��F�y�<�#��DDe�Sκ���>q��<��<��6����R-h���D[�yn���y�8��cǑH�4��":�G�BDDF��R""!�D&9�V�Vsn���]�Ρf$*���q����0�5È��ap�{�)Zޚ���đ�7���C��uN�Bx�I�nh�Լ5�5OF�kX�ߥ�a��A�}�/� ����>�	��g�f���i��f�c�� "�Q���V<�@M�'+uVR:SD�Nyj<�t��TE�F,e�ʼF(�0�t��� ��/�bE����7c,E��a����}j���U���ww�3��rI% .������$� ���;��5R�J�|���<�u�q�G�Sj&��4���mUA<��N�o����#�qޫjhөUW�+ư��U;tF
`|vA;♢�:.��8ҊọN�_m��Ø�k�]��Yz�MH;Xi�ݕ�Kֺ�IhA���S�@p0u�6 �;|;;��꧓��7h�8�tu��|�.v?le΄�����|<���ű��Vv����[ެ|e�5�2�W'�
7"��K�LC2����m��Oc:�W�/-��Ϟy�ȋG]GDy�6�4��i�]L��ji�S�UT��X��Wx��qh4�(J�,07�~P@�tܽ^[C �	�,�'��A�n�d�aX4S��5p�������,H}�Ф��}�����ujm���=6�2�Nb�s�W~��1�_L��2~�O��R�z���j��\�[�4~���j�S_;[��7��[N"�]��=�&�y�qX���Y�_6hV+���u��5^�r�����Ǿ['T�/ݪ���|��m���8��Z:�8����<�Ԧ��-2��j�a�&s�U>مr���k��R�q݈�b4������I���r�@�eW6É1��*3�/-"�#�`�J������m�v�+�9:���䋆�Dd��tv�q믫{�=-��}�C__��a"��Wս.�.���Hksl[Q�V%wu`�����](��5�6�Y�0�n���*H�m�Nr�Gt�;��Kv>ښ��~o�og�o���~W��u2mƞ%#�E(�~iő��Z�����ѩ˼uXS�:!؇���r�V�}�� G`�X���m��u}b�G���^<��2�^6����}�Ѹi�|^bAiN��}�k�)U�:8\�3O	��p�CD;Ɩ��W������+�'إ�uW�ct1�L��E&_0\�Q�S,��d���Iî��u���<>�5��UUV>�xu���:��>y���"""#�)�)�4�L����k�~^4[R�d�@`�BƐz��a=[^��]8
@�/j��=��$s>�D�{*U�;Du�c�CFh�I���To(�Kuh��c�}�檚s�Ü��uk�[�L~�wݽL�k�ߝ�F�z�ܶ���5cv�ev�V�Sl\i���6UqZB?����Tl&��)��)�hRH�c�W�Z��1��k�6��-��4�<u�;ʪm�;˪�+5ʣ�h�SUɜ�:�1�Kwi��#�<�>y���"""#�)�)�4�L��;��ۥUQ�M�T!�M���G�Q�-�:c�X���<����ri�V8�;�������4[x�j��~C�9R�|�`9����j�ͭ*��3j��w#����Ey.�W:{>���=4�M�s�������v�����M:<<��������c8q�2�qt���e<뎋�D��>Z=�r�xd����cH0j���Zx,~.�z"��b�����6��q�����Q�DDD~yM�M��Z[���{U��Ԏt��a�P�`���p|� ꃆ��D"�*�?;��F�r�dX4��6�.�fۿ����+���**�8y��tx}��O:8�iw}m����<��qx�<��Qױ��u��w�������^�h�i�?eViCG��И�����4�7���CO�	Fk<#KgE��� ��%Ėp:Dp�i��Ŵ��ȏ8��Z:�8��"#�)�)���Ku�g]�kZ]e��#�x�|�#<�7�2-Sĭ���*�4�Yc�c)�l�a��a3wM�DPe����bGK��6ˤ#(�)�!�"���2Ԍ�d������!��ƤV�"4�%.w�/I�[�A\����C	]iyA8���h�|�88.o-Ih��@oN�[��x�gZ���_KR�E�i�Nv9���Eၲ�	����W�]m`�cF]_���[\��@PZ��Ql��8U����c<e�����_[iŹ��T��ᤛ)
�~�X�A�їX%!���q�2f$Mcm;�]�ZgK#+|�l���>����E�T�Ywwb��"l���8��c��vY��y��e��3�]��ڶ�1O�iO�ش~ծ����4��yǝyH��#���<���[--�[r���e7X�$�hA��>�^�	Z4`tH��R���UŲ�;�+co��%����Ie�`�4]u*�>���=C����e0�m4?enc��OWՋ��F��9_��>&X2�����:�C�8�[m�AX1rW-P�,���%��6�M�����9N�4 �<	���	IH|=P����O�)N�|Yd�3IOH�S����8窾e����9��o-לG�ǝyH��#���<���[�g��y���jՊ�Z��^��=��9b���p�qV�F����I-����QX��n&��{�θ�s�;UC���xy���{���/��e1O~���[~qʪ���1�&>e\Y(���2���A��zC�2d�J�q�+�ja�it��qH��f�ݶ%��Zn����X���x��\��� ��)�̎��D�2��d��Z�>[��cjywKi�������s4	��8�����4��u�)��4��:����G]GDD?	Љ�JSD��L�z��$d�)�Ej�C��Pn~�N�e����M�z'Q&�w{��Oq'����!� vu�6a6HF�v�Hl�p��ZS����
�H@���3��tȔra0X�y�q����cO??;�>S��ꪴ��?^?8�V��UR���g�3��NH��Pᢥ�	�Ex]0i����ʋu�r���_|�ӵ_7�{�T�t�sr�>�{���������7�?��)�,��R���lٛ8��~g�o�zv�+��ٷN��qm�cn�0y�;�{�}���:ӿ�Z빷�[6��fu�4D[D�dMD[i�h��"&�G�7"-��mD�2&��h�E��DDZ&��e��,E�B-�"�DB,[hDE�M�4D[D���&��h���"h�"�B-�h�D�mD�mm��4X���E���К-��4Y"Y��B"-�""�&��km4DX��E�4D[E������""h�&DE���["h�,�DE�b�DD[DȈ��E�X����D[DE���[D[h�h��&��""ȅ������h���E��"h�����&�"h��[D�b"$YC�3���h�!5������&�h��-�-�E�""-�"kmmD�4[DE�5��DDE�DDY��[h�h��,���b�DMD�mE�M��"�&���m��mDE�MD���DDYE�D[E��DYDE��b"",��DE�DH��DE��"�"&�DD�dM��""Ȉ����"�Km4Y"Y"D�&�,�X�H�Ki4��"[Y���H�-��%�Y�[K$�I,�f�D��KI��Md�K$��h�D�D��f�Id�i%��Y��,H��i4��%�4Ki4�l�K$%���%��M-�I��,�%�	m"[I�%���bBY!"[HKi4��D�[I��4�d���[I��im"X�$��4�ĉ	l�,��-��im&�HI��K-���I,�-����D��d��[I,�,�Ki��ZBD��,�Y&�[I��D�im&�f���Kh����K&���KY���KD��,�H�Y&��KI���ii�d��%��,�-$���i-$Y5����4��ii	i	e�I��%��KHKY�D�!,�$�����D�d�d�Yf�%��d��H�[Y�Y"Y"[H�-��kH�H�I"Y"Y-�im"Im"Y&�Y&��H�I���e�%��m"I2D���d��Y"Y"Y$�5�i%�$��Kk4H�I���%���ĚM-���D�X�D��H��%�Ě�4�&��im"D��f�&�$I��%��M���X�,I��iĉe�Ķ�Ki�M,H�M-���4��&��k5��4�d�-�%�4I��id�B[H��i���D��K$$�,�$I��id��E�ibD�&�,H��k4��D�-�Ki%�4K%�im&�$X��[I���4��&-�ƶ˛c�#ke�l�����e��C�;u��N$X�K��1����f�e��[e��[&����!ۮa�X��9ÂАM�r4B!h$-�Sn���(kk��ZBAhD,�P�m����hHY	�rZhZBЈ[C���!4-���4,�n�h�Md�k&�Y4��kM#[F�i5�99-�p�ɤ֍&�i4і�d֚i�i�����M5�dM4��&��MY4Mhɦ��M4֚M&��Mde��5�M5��h��i��2i���M5�D��D��DdMd�5���Y4Md�MddM&��&��5���Mdd&��Mm4Mm4M[Mmm4MdК&�h���ki����M[MM5�D֚h�&�k&��Md�5�MY4Mbh�Mbi����[M#[M4��[MX���i���hMbh�i��De�Bh���Mbi��i��m4Mbi��ki����5��Mm4M	���k&��5�d&�5���M4Mbi��4FX�i�ki�Mm4�[M4�&�dM4�&�k&�i�Bi��2d�7\ۍ2kM5�M4&�2&�kd�5��&�i��5��i�i���&�kL��4і�L�i�M	��D�&����4Ml�i�Md�MdК�Bk&�Y4�D��I��"h��h�ɤ�M	�k#$�-�"ȑ�"l�&��4[D�i��扢"dDY"-�i�"h��D���!1dH�dDZ&�1hDY,�"&-$Y"E�LYBE�dM[iBБD�"[i��BвؑhY	D�D�,��ӎB,��"E�E�k[��DE�"ȑ-��"ȴ-,���Ѭ�DD�e�����D�h�-[k!4Z!�,����E�"E�E�-�D�E�Ȳ-�H�&�D�dB,����h�-�"��Mf��""��&�D��-E��m����m�"Ț�[D�dMDD-�E�dDDY����DDY�h�m��dDX��"h��-�E���",DE�DE��s��Ȉ�&�DE���Y�"�"-�Y�E�D[DE�k��"&�h�-��D[D���&�4[D"�&��h����dM""h��M�b",DE������E�DM��E�5�����&�h���[k"h����&�h��-��E�DB,D�mDE���[E����"�&�h���=��|��;������͜g�1�o������m�e��m����%m�o��}�}����>�������_�~9���o��np��~o��_�������~���>z���ov~������wn6��~����������b����W����׃���?����;�c��~?]������6f��������������������G�~����܋H�����kM��M�������^��Y�ϳ���g��o�M��������N���O݃����lͅ���������*<xο�:o��3?�m���|m�ʙ:�~y�o��e��g����v���n~^<y��<��g����W����ǭ��i�u�*���G����ׇ5�m�n}�:fۭ����c��n6�g�c�ٛif���cr�lDm�ݼ�8�}��k���S9�7_����g��}������}�ݾŽ�M�6�&�y�m�H͔$f�62���`����?���7�xm�~���v��[��>_����>�>א�h���;��Yo��w�uxߣ���6fÙ�n<]m�o�����m��m��[�oH�7���}��z;c�w>��;_�߱�~��ݏ�3�~�Y����������o��?��>_�����~�FF�����jw�?����>��_O���s~fú��cfl?��w�m��鿏����[���c�=�K������ϏYyɳ������`�}����7J��b���m�͇0����7Y���<�<�]ۦ��O��7~���ϭ��=��]n����o��L�m��ޛl͇6;���UW����o{5��Ǐ�6f��S�?�F��?��~���L~'����������{~���u��6}C���o��7�u��v����_�o�&���~�o�����o��g��fl>�a�m�o��������Q�6�������O���}~������������3��޷���m�Y�e4��I?ɻ;�eK����v�����~������O����C�׮��������>ͻn���u���<<�������s}����g�~���7�q��[���o��>ǭ�>l��-����ݳ���������M�oٟ����������?�������7��������y��=����9����/.g��[����~�~��|��#M���������]��BC�|