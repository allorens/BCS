BZh91AY&SYqB� �p߀`q���"� ����bF�:�   R�U@�  <�$�	B�JIQ*P����E)@��TP*T�*�"���R�RR�RRT
 ��"AAU 	%(��� ��%)AP��*���T)J�T  �R�*����UU(��H���UUB���  ��B��D`	�J�U*��Q�)U�l��U(���T�T�����J�DEJ@�%T��*�H�
U%T�U)R���	    ��1)��-��ţ[M+cU%� 5�Qڒ�b���E��)&�֬Pڕ�[[j����K-�@��
I!$@\  �@d��P)@!˸ �P�2�
 ��  h'p j�:S  �HB��԰ EBbԐ �ʀ*U�Q��P��C�  &ۨ  ����J�9w� �����e@�� +T�]Npt��n�֨�����#��C�J�F3�t��
;UEPIB��
�I�  g�P'+�҂]L�{x  ��M4�\�@ +���'mPs�h(���� ����l�ݥ�S��J�UH��R*���  Mp ) �_pt \W���R7f� Ҫ���p@8�9��.��TQk`�Sb��5B�	р �6�H EP��	   �@T�Φ�)@��  N.攠WԠ�JtpPm�b�  �XiBZ`�]�P�'p�P�R�UJ��UIDTB�8   f�P *� Qe` fX  �L V�w  s� �*�a� fWp :0@�EJ�R �%Q!�  7@I���P��@�e� �  &S�� 8�  &0 ��c �IT�TTJ�% �  Ӏh�� �� ګ
�ڋ E� �4�, YU� XKh t`@�aTJ�
 �����  k�(`� bX j԰ �` Sj0�` Q�� m�� f <(�   
�֕O@R�(�  �& S�0��Q �� M  )Ji����O56���h�����S�A)IT`#�!����1��UFѧ���M�b2h �IH���@� �� ^�Og�ۍq���|o�MoV㫾q��=\��[�v����[�x���7���"IZ�z$bI �������@��Q=~=�u��$���L������w&��D�C������e�'�ć�F�Y��Ndy��9��^N`y��y��y��y��0�Na�Nd�N`�^d��2f`�d�`�`��y��y��y��y��xd�e�e�`9����e�d�d�Na�l����y��9��9��&�Nd�Nd�a�Na�`��9��9��9��9��8e��9�c�9��9��3sd�d�Na�Nd�Ng3���9��9��9��9�<�̼��<�̜��<�͙9�2s0s0s0s/6g�s0�2�'2s'0��d�<��<�̜��<���9�0s0s'2s'0s6`�L���̜�����c�3'0�'0�'2�'0�Ù9��9��9��9����9��9��d�a�d��9��9��9��9���&^d�Nd�Na�Na�\�Ù9��y��y��fd�Dfy�`G��Ty�ȜdG�Q�y�^d �e��A�Dy�^`W��y�dG��9��A�y�eG��y�e�Q�y��D�y�0��	#L� ��1"4�df9�eW�D�R4Ĉ�4�H��0��I���Py�e��@y�aG��d �Pt�H�	#L�4�#LB4�`G�aS�A�y�a�T�Ay�NaG�D�BeS��y�NdG�A�E9�d�T�`�Q�E9�Nd��Dy�a�A�y��®X�	a$i��b$i�F�#̢s(f@9��2H�#L�	#L4�L�)��T̈�
<�0�1�H��0#LHe���aG�A�y�d�A�@y�`0 fDy�e��y�a�Y��E�Ey��U�Ta �&U�TNe�e��y���$�4�1�CLD4�0D�aX4�C,�	1�aP�Ay�^`&@y�^aW�U�Dy�NeI�^a�Ḍ���U9�C� 9�^a�U��Q�D`�Q�@eW�^a�^y�0�'0�s'0�/0�9�a̜�̼�̼�s�0�s'0��<�sL��̜��<�s̜�g�s2��<�̼�0L<��<��2s̼Þr���^`9��y��i��s���0��<��s��0�2�!̜�2��<��<�s4�̼�̼�s0�/0�<��s�<�̜�̜�̜��L2s/2�̇0���fa�<�̼�̼��<�3�0�/0�/0�!�9��0�̼�s̼��̧0�1��O�}�c�[��)�ћ�7wMdU����:��t
ib����1�Y�hϲ����\�7��i[�[��P�4M��%M�lغI�0�e�JI�����3ws5+ci��HH��z�l�<��aF�����R�ak*���h�Ǆ��&nc)<n^S�[�ZgwFo�[��wU9�Ŭ-oV��#4�f����sC�q�4��f�Z�P�8jۂ�������bL����=��9�BZ�d<}��[��n�Nj��%�fiz�G@�P;' ��̭�N����.�.��Βe=A������-�zP��)%��ģQ��bKuux�d)43�J�	sY�;bi��
4h`��m���n"3FG%^���-�h\�6�Z�uNd�ܦ1L84�D2��*�\�Wz#��5 ���˒�!ݏAGrF�^���l�O0 ,��ޚ���V��b�uekJ�J��+�J=�, ��ӯ��]�Vr)��'�[�	(41@0�Z޻�(h�f��j�qm%R�(�jZu䣲�Q�D:-;v�R��!���p��B�.�h�5{*&@���&�m<���E}i�wF�kmvRU*�w-m�9xhKٟB�,ݡhR���Vn�HN� ��#U X\�mU��5�Q �ZX�!�(�!w�t'WB�a�,Q�ZA7P���e[����D�KP���Ѝ]j@Ӵw2��x��u�elm,�ƌ
Լ��*cB裥��g�o5J�GV(�\�[p�\��%�-�x᫽���Չ�GC��t'@�K021�1Gw�Bi�кݴ�K�B�ӭ�6&�B�EK�LL{F�ڎn����� �L��(�M���xB3Z�k,p���!&�dl��3	'!�FM�k	���%�U���-`jģƌչ�*��͚���k'4�L+�8\z3aO
3*��k2�-U2�LY����ˁ��Af�a�Y!pk@k:%-�1$�А��&^��),�.^7�.��u�@�n�#zٙx/�ܭKZ����u�jRl�F+XɎ��IUXsa,bw-�%�z�Ŧ>��u�51U�a�U�I�F�|��N�Yo$r,���Z�j�����d��p�Ū���&E
�0��ϰZ�@^]	��gp�&�V/IB�xoH��M��E'���-��d��aj�{o$�|��P%��-h1�8��Be�c��Ѷ/�;����,�E�7����a�5��aQ�%���)d�з�!M8�+{Q�������۫�hH�;��N�83\�`�n��^�cy��t���Ie�0h�'7bx�:om�m`j���y
�yޫ4�h�4ΪfEi*`Ә��h���S$o��c�����#a��^���d	�mwu)kZl��I�[�ˤUi2�� �bm�jWK2,��vb(�S����֦��r`;J�JRWHO����F�SM�u<�腻R�M��y�apj����q-4��e�˧#N�^5i|RL�B71m�Miy.�cM0�0T�X {�'kH��5���Z՜�n��⡦�խ0Ũ˼�܍P8�����*
z��D����]����M�I�(���·������Wq:Ni,m4*e�4��ɴ.+�b*|Pɏ�1  !�9AU)+����=;-;u�$���[[��G����ի҉m\���T�)*�BM��ɓIT�*�S�A�/6dt�H+�l�wL#e�A���U]�[�@��hw#�`�XB�# 6��bZ�e]]��+�WA
V��bS�+o�e1r��Q)��7i����2�Aq��U>�FҭJ[��2�. �檈1(�7�CH��-�яUd�E�#5�S���[w[�-�Lw��Q�����%��+N�]V����J�(ihV�bh�&4-�Cc �J������&i����:�L^��+mO� �J����KXf�)n��J�;rJv*KS��ͣF��B��Ղ(QuB�j�N6C�/)���`̭J�`=$ �;y?-�L��em��t�[��������?@)�hBU[�s
Tf���h��S�Cv��T �-�Z�g)Iww������G$׋�K
�kjE �v�ٳ�Z���b� Ѳ�w+V�6�+��yYO �j�� !����w�ϵ�Z�Q��le��s3)�P��M��z�Y�R�����kْ�`m����e5J��xC&�9��K�Z��z���j���5��,���Z�	
��0V�jQ�ya�-`��`ź�ii�c�>���z�^��Pr�����:ÇZ ��LL%m�����R����+`e]��F��
Mqɗ������^�Æ�+f淘�^�:�*b���mԈ��/3 Љ�,u��E�{!&�ٖ@v�̴�[B����[Pj��0�m�(���t��S��Z�R��g`*�M�Tޅk*2]�g'�`�b�n��]�@\Z-PX,��ک�+&�K4^���s�i�r�D
E]K�n�fU�B�{ѵV��[M�j�s�V�H�3.a��-R� ��E%�RL���.�n"[��o!ytD5W��cr��(S(��LY��ixi��כZ����bڳ$��Ix�*/�ϐ,mLf��iT賴eG)%����ی��.4n�;9Z��0f��n؛�r�A���`��v$�v�	!��,��.�v�;������a�m����_���N�L�rd�^\d�w�cY)����Y��ڇJ(�H�1mḝ���0%��3�M���!��$iT�4�{q;�˂ӗ���	�Kk*k�z&0��*"��@M��J3z�����Z3f�[n�4�Y���$f�$uk��rT�' �(�R�à�{�+NU�����朎�F��U����m^X�wN�,��C��C7Ʌc�p��$����Ʀ�L���L!&ءJ�n��1u���Fo����ڒ�zs섨�+��u�f�Ph���1&�:lՌ8l]@���b� "���&挳�QQm��Fv�����+wd�o�r�Y+f�	U�L��.�R��x�����w���0b���мj�)XF֛�+4\{u�N�h�$K0�e]���Cf|���q�x��5� e�iH2\ō�Y�E�Ӻ7nX4���A��V<vZ��e���6(��u���V����p���t;�e7�J�V�.������Hы�!xd�aՊ�AOb�E�ź������L�O^��%�Sf�:�[��3��f⥖�PSwĮ�zJ݄1�3wOv�j�b<L��˃��"O6����gKL�sE�X]��i���r�$r6]-T	xY�^1N*��T������g5��[P�(�,,�y#�$QÎ;ې^��M�X�x��ztе��:� ��ꦗb"X���ݐ͚0̌�F��q��P�r���w-��K��������nU��m�z��aJJZ�2�h�5bl&�7t�f-�^��*:gh=��c�7%�K���GH���Xmڍ;6�R��5��8#�ݔI�ݗkS��X	[&�z��+�x�M����mT���U�Ol��"��Kj[3E�ȋcm%�3dɡ̙@
�SK��q���p�0�WF����W�!�.'��q��f sV�w�2�՟�x�Z�
6�̕�=���K��!��T��W;�(�̺w�O�{uLֲ5�
	�4�Է��Hz�fm�f�hܒ7��saW,lY�٤�@%�'-%�ʬ��0�s��бl�/&]4�N��'�����L[���T uZ̑�r�Je��]��o�U��1WIX�C���N�����32�K�$����( u��*ല������fE7R� ��*F��`�L���r*�?*�.��k0YL�	ͶX�;̡�������e��)���7��;�C�.���Ժ�ěۼ�6;D�`��n)�d[�f���^=�m1�8d��ܭx)��fX� )2���MJRˬ�/f���.����q,�H����I��;5c!u�DQ#R��6X�-��X`����f�YH�͕{M,��qͬ��!cyy�b٨�;0
[%�P��usV��f���X]j�*BE��wnjvr�dō$�͚6�0��KMVt���U�1Hț��%�����cXld*����V%J�r��%Ưr��ڤ+^��;F�v8]Lf�M�V�#MCJ
f���X%	4�C��&-m�Io~�p]3V�M�跶�j	JWWxwa���tFJ��
��*�l�h���v�U�X`�1b�Sq�Ʃ�,GM�^��FY�im�%�-`�4��^,�$���%n���p�&mX� ��^�Q�O�v���l�ׁ�Y�m[�
�E^;%���I�&��\�nU�[�*��Z����nd�[���2���p�de������*C��0�@�v���7{V��
��o`�5vm7kx�(e[&�5�ai��em��%�k�s��M�L�+L���+=ֈV+,PO3l¡m*����J�T@�
�]�.K&�-�zFZ
����o57/Pɶ(
0�d7,Y�v��H��cv	>ƥ�b���#X���K�M�sJ�u���$�����l�L�ꤣɷ�J�
�^;6.i��S1��x�"y���ȼ�"��A"e"򭻁�}�d��Y���֫4�!�`��m���@�&����5*śW�m
�a�5�������j�X�CO$�n�;E�M�"�ͼ���Ň���_�+�Ǣ�T��*w�V6����h�N�j���VvU�E�R�4�M�[��/!�a7t�lͦ�p ���]���x��)�-�V�i듛�ǷA��;XÉ�9�dFt�y{Kb�+BP4��xأ�j|k/7Q�L�aې���E��$6���fl�7S���
�B۱A;4cnT!nۙ+%��Vrm�����u*e�[���=)ltJ�j�{�n����;w��t�* ��|r����V���n�m��Y�c
�\��I0�`ֱ�^ēaa{S.��̙y�����A(�+t��w���*IdV��k �+2,�x)X*3�V��Մ��� �d\��Ж��դ��B��sM���Je�']�T�O
hŹR'����+3T"�5�+*,�y�N���"�-��J�3r�J�jP7Y%�1�n" ���)���8�o��ev���r�4��ӹN��C+N)yID]+���[���`o�R�f
�ɢ�-��jY��8r��#�{���Q��B��Zaca�f��w�JX(U�Op��4h�[F�e�O]il��#C�)�e�.������;�1�n[4�95�T]Y��X�-����� U�0�YE�e-�����"��im�&L�N8�CYe6����nQl\��h��[�P�1�Kd�^� ��th����͂-�sk�YZ�	�6e���j�м f)j�ӐMx���M!q�Ļ��d��n�5����%-Ԩ����d��a�˘k�� �t�,6�$e��&��_����@{���fC��D<� �]�۶˔\��2�V�:�W�$+f'B�Bᩮ
5�1	�F,�U�5-����V<{P�claG���7[��q��srm��)頲��˔Tz x7F�6)���)�ۖ��7��!Z�y��ov�3S�RQٙB��je#B�k�0X�̀�TV��b����ͷ<�#Ԧ5�����g����ܖe3��Kf�U���'����4�#2 �9ocQ�X*=�^6��d���!�≡,F�UŻ`���޳sk!ƕsѺ��S�y̗K�v'e�N�O!a`�m
�(�æ�`�j*aC
f�ٵ#j�T��.���E3��
R��f<������b"���4]�3�V��Sbu�2Dl�n��	�̲��z�wq���SD�[Y��RPR�OU�2C.B�w2	D-����)��G2�y�J�N�A��en��R!�i7�Xc*�6��{�� BJ�1�n�"�IV�B�V�����t7��s���9%��8�C&�%��V�h�:��3�f���T[��v,L�����BN������U�����]:���i1)ן3b����Vf��D�doYwI�ܧ]�I���SI�`��tn�KV<��]9#[u,�ԯ�(]�ixk�Ka�Z������a�°sjK*ƀ)�;c{ke����cX)�Gvl���N����tf�'.�!��`Y �Qu��Yz�^e�wB�B[�6d�2�+D�¾�Oc�&�%�ە�����m*��Ώ*.9��X�X%2^NwRWB�^���:%̻�ۧ+e�VL�(��Ê$K�$8���D_Fb6��L�OS
���[8ѫ��E�J-�d�v;��J�OTR�SY�Tyr�^
�Y��&:@3A�BY��m��Cl��zz�İ���Ǧ�պȍD��-�բ'c�#�N{]��I����m�K� ��<�k�̺�80�C��(Q��`A$+cx\U�H�;Cݶ��j��8+ʃV���>�7��t�&B.Ү�*g$.V�aL���ձP�M�t +;��]JQn��s-�����c�-k���*�7>�5��f]�{�E��>�μ�l�{L���yjS{H	�E��yt+(�8rRVĽ�V�w�4n�+V��n��M�O7���yb�uJyaLyt�4TJ��N��xkV��o].�c�W��J�c%�E��1R�
�k�CAՠ'|��Y���i	01����Dp�4W�8kq�82����8����[zܺD`�x��5Y+��!!�ڰ`v�$B�vJ<���ol���T��a�D2���$.��]0�*S�y��"�T�tc5��*v���p���X�D|@�����/�?GwO���я��׻6+vo2���]Ѭ�<��X�Tt��;�;�Χ܅�j��+qQ.��]ܔ��J��k�J�u�ç��o�t�ǎ��ԅ#�������,��.�S��k.h������gp9Sok��5��ii�GLj���iQá��G����icJt���k$��FGW�\T��?�M[\�#�^b7��]Kl���T(�[��.��&-ξ5��];�LP�����.k�ۋԞ�<��Lv(I �p�&K�f�)�iγ�2���Թp�[erY�`�z�H�Hf
7p�T�N��݉p%Y�כ�Q�[j�J�L��]�9�]	x�#�<u����y偫�2k��8[�|�;ոuG/��%F;Р�N����`�g�0+�H�=��^�o�N�X5ʐ�Kst�|%A^u���u�X$�S�L�oV�yAu���y���#��>M��M[H�c(+�sM�YN(���ƴ�!TNܫ}�m%��}��Nv�u�:�5w4�qM���ќ��܍w[�]=Z��]��/&�J���O7 ��њ�Ա�DP��D���(8/�����;��$�����Ge�DoD
�����5+ ^��*������792�ڸ�}�;Փhu&N�����5�����Z{-�4MB2��rZز�������ą����(�W�wZ��؜���7�+��@:�=ў`t�0bO��*�jjo2W�3s*��dSRI�˦
����V;0k�1�vu�)��n��l��xuL�r�N�˙�l� �gF1evc�FRUӕmՑ�-�~ᢺ��Lt�[�������p��ق�g�<nM�a�<ηQpPG��;N�1���`Ǭͥ��(˅t��+�+��SWZ��F�^�u�`JU|d{\{bb�X��84�g�V7��0���s��k^���Xn��/�lYs�[�o��Z�_C#�í��1�ŭ�b<���'r�vs�W�u�_\Tﯫ�JR�g��]���Xs��t�)h�W�q,��Ip\x�*�9ק��	����.0+K�Bء\���\�Bvgoѭ�W�I&�j՗ϯ� ^"��r��jԡ�n+.���pbA�
�q��yx�� �,�]s�kq�)�-�N�Ѓ\�5[��.�n��'l��Z�S�r<��2������w�5�(�o_\�Z��\zc]f!,Yz��;{��F� �zl3Fe^������]>ו.��f�ؚ�ʳ&�`w]ĭ�Z��Ón<��Fs��w��BF��Uwn���؈Nn��}�:���Ὕ%���e=�A1�\pt��܏��ޞ����CF��PI,J��Ш�I+�#�� �s��9����|Eb��20�g_�S��e�},3�Gk0G0>ݷ,I��3KE֜��eȏW[7F���֮RПs��r��|���&�m
[�Y�J�s~��Mc��w��C;bFc�\�;Xc�uw9un���wr�X���]#���ŕ)mU��T�Vzys�CYw��Z��AQ��2ǉ�ۘ[�o(ؔ��a�gj"�kM�R�㓯����M���������������3(Y����N�C�F���UǇm�n����]F��q*�%6�Q���QҢᇍ�w��t��Ȥ��oe���w��i_^��%���ޤ%�v�M�Z��[�ZKM�-��C)x����W�t�����m�s�y8���g��E����F��N��k2��U�˕����-�[�r�.�������q�vA:�\�Է���+���-|��y"R�b:�����Wm ˔P���G���.��K
�*�s5��l*a	������ً�:�����.���Lw&�P湽�Q�����G����u��Y��H蛫%�{���g)[�J��
R�r��X���-Ǚ�Ż]ԫs i^q���wi�s���D,�Ѣ�Y������r����3�����K��c�fCQSB�&S[�Ɨ>Y+_Q��CPN�r��b�+�N��8��W��n��Ѥ�*��f�hi��woUֳ
�f*�NԷ���3{e=��Z�=�+���rf�R�3ɼ��A�nP�H�ԝ���l�lN0�� p�G-����joc�i�&�-���PR�MTBQ/ ��e&�������=�s�b��[@w]f������g�E�)���>�dV�y�U��Y�M��ƃ�G�h$�^9��׶
咹��Z�/mRy���"��g��u{41r��Jة����nL�+Mc��uZ��A�gq����V%*XЊɣS��t��=Ge��z�%�P9
fr�]��Cm^��"5q�N����#�2h���U��'ۆ�hˣ��>�pV_X귤*m��lȬ�uxs �B��]'��f�t6�=��2�`>[�]�F�t���xҧpnT}0a�K]�e9��^5�y4�YC x�G�e�+6�!�~�!gh��5�FQN供�t���j�,橌���
�>p��*e�]�LE!�$]Kٛ+Ae��W�۴�e�/ ��{��A4y���0� ���]3d��윇�3^j��PZ�[Wȡ�Z�ϔ��6>)퍹�ٙ�'5סlR�W)]��a\[&&����֯e<�gd}Y0����V�\F�[ۗBA��Ę�WtxiU�s�4e��L'���[���uH�zf�]��~B�*��e�T�E��V�����C]J�=°�ͧ�����oqn�#��}��tX�c֤q<�h�x�
�Ѵn�8�ʡG�ATq�`�N�Hu{��uY5)R=zk��%�2�#�t��iY���y3�vYV�˦�t��A�̻�^�y�A]�Xd�b��oE<���2�V4RΛ`tt������wR��)']6��G��qye�w���� �_�3�eD���q�-,�z�1���|�6�;X}��:�Y`P�	-FN��V�`3Z�]}ڪ��%iR����7X����k}�Q:U�S=˕'J�Zச�	�4�G\�W|�]��X9���ܝ4oQU�x���6�������ݵ]��:ΩI��X�e�N���)0,5����R�����u�;"o6�|�]]%r��ٛ�r�����{�	�5�kwv[�r�3G��x%],��-�*��ekSdIˏ�V
W��*��+q�wO۹��][�u>Hp�l�I�`�y�6�GT�&fv�j8��ie�Wi�����ީ���o�T�V�ё���Δ(�-wn���nO����Ҳl�(���A�_]s���֒Pste�=Lu��}+sf���R����;�e�۾��eqҰ�8��CWA�:��h8��Έ:��	���]1]�����X�\�6I��d R���wA�-���F���n�7뢅��8�����������%�b;/�d7n�t�FC��j����U�7��mw`�o�Sò�𜑊PL��׆5���{��-vI��ʱ��v�L'MWz������Y-�Z{:ݻ]������{g��8RF?%�L�a4��X�n�X����|�ZϱQ�����3�Խ%i�!Z�Y�e��c;�ݵ����i��Й�8��ݮ�1���;����|�+D�Cj˩�9q`�m1��&%>#cZ��F�Cl]��C��Ѹ�	HR%r=S���[�v�N>��$�,oL��T�qh�u=��0�&ڽ۵�(����T�WmSX�V��v_L���k��W�%4f�y�`��HT�F�7�/�y��lv�����J�L���
»�����X=�ե#���f���~��V�Xu�T��)<�"N�v�rp|	 MGإt"�m���9�*Ww�����x&pbc�wXm:[��
Zq�Mv-Z��Q,2�Y�AĂ�u���)Ky.V�X8�8��{v��gB!��HU7F�45��Mpͩ�Su�C��#9�غ�Q�C�l-��G]0���΃��
�3jb����b�tݦU����O�ժ+ޙ�)�Q.�.R�n���P�M�e��:�`ꚤ��OD6t[�sz0^4N��"��Ȝ��0ɸZ�`���Q�X@�;�����Z�i�uǕ�޺-dK3�Zt#�]Wh�8<��e�c$8Gy��9�,c���b'k�n��zN�խ7
T���GW����Z'6@8���W�N�a�2��~�{��ԭ�u�<fHX�˚��v�ʎX��������gf�U����Y��)S�g
����k�ʸp��y��E�&[�З�>�=X�٧��󷐐Y�g��hHh�X���6N�gir�\��fp*"����@PI�b�m�]�-$m>{�}���N7δ�}�.��{a��U'��[�O,�p8EX���o+όJ9M�(o�r2���m�K5}�K�Ef���i��`����',s�F�����t�^8뻩�-�y!v�*
��О+"q�ol,��C��hJQS�yK~̿j+ۖĽK��R�˫�:�%�"��"F���^��8 "�r�F�Ԟv.�e��`wp�4��lY]���Ub�$�
L-�������d��,3a.���b����=g���n-fIC�J.ᒲY��[`μF��m���e�F�[��Ԃ�O{����uuv�<��׹�T]��q+�>S2�B�O
;�:�Dэ�W:�\���ȵ��ƖӮ�.{.�u���z�pW��H-��2H-
�8�D+����N�v�7pwV�� F6��2t�0������	�fL�/�ۺ/U��ݐa���Gi���W>�\'�`ı�_h�{�(���TӲU����DN���*k��r�ו�:we�V��d����^��U�K��`Q�S�ز u�髕t�[P!yEAbmcih�����cJJt}T@�r����t%�Z�%rdFؔ�g^�Ζ��k^��.�ъ<�%U{���f����T�M]�u��Q��k���.�f�ӽ/>GΞ��&�vx���s{���u��F��傜̷]�7PTl�YZ^���݃���u"���o��]
�G�;�f)m������pu�2��;D�.�J��]u$����|���շ���g���S�0���;�G���l͢�Y.��3KS����zL�u��WA`�tI�,�t��
�l�Z>�q��Dr=v�v�'W6��н��F��8��Ɋ�;��"�f��%�MTyvо��|�L���kެ�X(Z�J�����+�uż����0��Z�8��+��&R�pY}oWm�/a}6Y���;y\Z(L���V$���6��t�����BO3��^$�V6>�k�"�BsQZ�+�S�;Lw"��Ul�$�(E����U��U�í��.]k��$��r������-2�gA�M�M�[M�{�4�׹L�����ʹ���R<0\ӓ���+
1'J�R��0Pkaʎ͛����AЌ�k!�6�F�DB�$�}]A=�/;���rO`+D�We�9һd�r2�{f�Wkht���(���o�w\����oRׄ0�Q���/z�;��:Vt��R���~��8��l�4�պܥR�qGUi�܂��N��7]�{e��ocS*%j�f������@��m֍��4�q�j�A�h1f����F��rpǻj%��s|�+
���n���έ��d<�s��"��-�ΤM̆�Ժy���#�E�vV����F�ClR�cXʁ���H�.������^�H�@�aOZ:��_Iq��n�&��s+k�e�&f�\��
w'WY����ט�[I.�G��e���������ӵD����1ƃ��ٵ��8��\6ӥa:{d��v����-�7�(�Z6d�Z�ml���\�Ln�k�Wyǘ��h�+����yӼ~ں��<�.�c%��v@v���U.ʔFu��#;n/�K�sy�mô�����~ׂ�M��dJ.C9�������!۹]�z\oU�L�kQ��v+	(�N�oT#��v�=D5Q����ag]�g��I<K��*�T�\���¹��(E���8g U�nm��'!���[%N�WS;��uu��'���ǵ����J�m�r�Cϻ�%dm�{����Et��e�2�7���v���Y�<��xl���]��PQ����I��d�]7�#f�6[���R*W�  �Gc�@���$ �+`�O��ög�[(��"QI�;�*���*N��@��L� Le$	��@�P`�9e�HҤ�L���qT4iRV�u"RM�M���h�( )!h�4h^�������K!DZ8�>����m��\��~ �aQT�n��4I��Ұ� .�J�n��5��
�Ֆ��_CC@
��������
m�A4��^��y瞼�m�]��
��5Ӣ��PJ+� 7R��>JJ*V�N��,L�n[�K���j�Tq� @��S/1cN��SX�E�hڡŇ�B�3u�J6�$ѧ��t��h�F�A'�'�qf�ʆ�*Kk',Qb��Z�&�IR!8S�ҰY��&�II܎o�&�J��@�]St[`� ��J)4�f�'�E �h����P@���GEK�)�  �)N��N�-�� �M�
�l�M2)�h AE3H�h��
��h��e���lǁ	��Lm��
t�q+���l�hP)V���������ĒH�I�߯>�||�}�"B?O�_)7�_o���9�ٌkǳ��y��8�ňxC0��UCK������B�z���;W��/���5�'��^&��8|ĭ�w���,B9����yq�(6m��T@oe0e���t�\w+s���[/��7�FÝ��˚���&�ރ;B�ZPN3k�-�S^���瘅��ݻn\�˚yS�\��֖;.�L�E���&��t�3tn!�^-��%�-<��z7���R����ѕ/�M�I�wn7���b�S�����@$ຮ	:�Wa�6�g�Q.����p��}H=�-cժn6�NR��w*�|�r�"�(��Κ����<����81Q�Ԧ�ߡ�uh��u���OV��!�]�nQ��ܠ@��Y|�ʷ�--�,a��x��ډ��Sp�}C,�h�yY]eө�GCz�͜����͈&ȥ�#I�ǔy���6gn��*l�9(�������u�ح��n�k����eU�u�C���w^а�P�6�tGg'}����I�^Z�`�j�I���a�SLv�N�QpK�OWV3y��),|�|����q��n��f۸i�e�{�d��V�O���Ց�3Ք��*�i�WȤGn�-��ݢ�	��c�f���ҏs��C�s:�k���k9��et�Wa���q2��A�i���vӶ��W.\�ڪ��UUp��Ҫ���VUUU[X������UUUU[VU�UWj��UVYeUU[VUUUU�aUUU]*�J����UZUUUr���UYUUUWj�����UV�UZUUUt��*��ۧm��m��Uګ*���U{ֱ5I�J&I+�#cqQ,��'�Bb��9j��Dy�)��P�SݣA�EՒ�r�m��7z�{��,����3�����;��;�W��u��!��k�,ΐF�ke56��mLq�u�1]6���Rv�X�(c5&ְ�[+X���ѷ�ו"oI��e���ł|;�"\wD](�	�UUnpK���Y�������Wشٝ��u�Y�J䠼Gzn+�Ńӣk��������W�մvs����n�+�.f��)0ƢF�'G��:]8�c��mQ��e]=k�c�ʓwO0�hk��o*Ԙl.���j��)u'��s�I�z:���o�M���xW���mdU���ﾩ�}�F��ݠ��Ӧ1��I�6�$ƺ\���4s�Q��=� �7f�9}�@7ݚ�w]�u��+{C��a���A#�8�C;̼�}WV�u�Ͳ����e�����H8'��M��=|�J��]W��pG7A)�2�])<d�UaT��N����8���e�����w6�C�U*�VU^�E݌��j�;��Z�U�L$��>�7R��5t��ѹw�]��]tɼ�a�vⴝ���wmNC�;*x��n��5n��]�i�8�=��=|�U�S���6]���Ӈ8w�UUUv�ʪ���UV�UUª��UUiUUUҪ������XUUUUmb�4����UYUUUWkUUUUV*�����UUUUv�ʪ��UUW+�UUUV�*���UUp��Ҫ�ۖ�a��mUU��������/C��W�[�����-;�h�EL1Kxԣ�J���}��[\�ۂ�Y��>���X˚m���J�>���@����w:�K��܋hX\"�^�F���_^��u׺���G!�v��
����Z!�(���,��+{��T6��� ^FD7Z�!K<4�1�XAQ�ժm���
#M��
[�qr�]yի�]�;$s�Ju�'J����kklj�jJ{��U���M�u��p�[����3uk.�Oi�Υ#3�i"�.t_�MY��l�o(�}4�&�%��6�ZDuv�T���`Y�Ջ��uz���N�eǆB��Yu�tE��4��]��*�̷x(�V��TIܰ��*\�wa����Sov�0B{���]f�j���F3'V�:p�Ժ�69��K�,+��ټ!<�NU�]k���OV�W�k�ڮ�Kncp@T��;�;�7fqtLZ�N�vKd[�[�_J��hA�,t����"tM�=�	"���Ϝ��ڢ��-7�j�e�m0��M�Bn�S��ܘ��Y�r͎]͉nosp�,t-�}j�u�dAxOee�-1�T�#&��g�
��aU5��*h��ٛ��`	���N�f�6�"6\Z���G<R����w1E�]�<���ZͲ�!H7a��3X���}�Ģ�gvS}��]Û�`��7�g?���>�w����~?/��ʪ���X������ګ*���U�UUUt��*���UUp���UUʪ��*��UZUUUr���UU�UUWJ��*���UVUUUU��UUUWj�ZXҫJ����XUUUUUaUUUʶ�M��m�mUUʪ�~������:$��;٭��_7��2M"��u�Ն;���<CV1%hjJ[;V(.�\�v���I0����T��դXN��59t�n>��Y;.|i����5hzђ�H	���jYӾ����.�W�K@�{˗KOQY�s�{*4�g���;'4���|���W�n�b�[Kn�nЃW7-��v���=V^q�q�Ӣ�tq����b�M��TU���9͍�Qw��ق���=B���/kevPj30�3n�B]��
r������f�u��l�U��Xp�õ�F��U�v�sc�n����U��j�L7K��u�m�r�
��L K�v��o,:�a�ʗ.<U�HɝV%�
�*��z��Cf=�._NB�NG�����p�.`��ڻ#h�@�HV�ݔfbw���.��+R���`QJ�T�hڧ��O����
쮙��֎�Մ�ǵtt�y����[�^T8�[m}�eޣ&�2Vh��Ӻ�'V����`'3a�I#6����uDܵ]���˃%���n�*�J��P���LWr����^�ŧ ޮfPB��N���L�ύ�(<��FU�(��J��bY��:�մ��8������mt��vv���`����Oy���.�Ԙ���[t�:-��Tj:�U�1�S��9[[��7HX/��vL�:#��F��@5jݖ��R�gJ儵�A����Z&u�����6�}���F�2'�[c3a��=���
+u�����wإ������$���d��&�}Hop���S���t�L�]��'�͑l��L�a�Ҿ�n������	>o!=��Y�J�+m٭=�Y�+0�A7���-��*d�k����4 t��C�RajQu�Y�@�(��=@���ҁ�&E����N�%o�˥�!�A��.���{����:�eMGl�s�#گ�f
�(L�0���q��U����wSQ����n��!��q
��9����b�H���;����R������ʏ��զ�l�x�š�{Md,�a"r{>&��Y�M�\�"���;�����i�m�{�Ѫ��S���o2�'+�z�eÕa��K�ç���\��/ u�!я�ț�r��u�m���}4��6�L������Tyg��}���u�qD�;�]S��#�Qeu�8	�
������`��W�q�U�ha�"���X#��S���C�e�t��u�g%�CHǈ�.Rs)��%ۙ>����t�S����H�u��^v�5�8KP�N
營�t-s����/8X<+���"��*v��Uf�7Gn^Y�i�:�������� 
i�4`�-i}���+���_$�Yڈ�T�s5�B!�9��//'�I��bp�oPݧ��_5��&�ʾ�<��|�K@�݀��=Ŋ���ӶR�W��s�.W�8�I���s6��쫂�ЫF�;��g}��8��1;_e+�Rz�Ӏp��YٵVڪ�I�r؊�n2��X{U�,#s�T�^�,wwP�Ի��+�¾���,y��:hu��� 	viS�x�V�*��z/���f�
'�Rv�������cs�#�j�}��g�R���jƮ�-���:�d�5.�}���x��v�.��6���Tp�3�P��Ͱ��Z�ʆ�*���b!��m�Z�r��\Pb��@�9oA9�Q�-��"�Y7.&��\�r��8�u���������ٙʚ��v�]N��˾hX�2���u:�"��v�ȫ@ɟ5�=׷���V+8���iRA�B��ocWu��F�[5�3��9	}���JJ��u;��坆���)ܕs=m��ՎT.X������oj���Ƒ����gnK��WNͪ���{HCZZ�62hȺ%��n�hf�:k%�Ѧ���4ե�4LV�R��6p�w'��3����`�Y'j!7Hߔ����{T��۠��k�����]ԯ�W]1����XA�Vr+��@����_�@�z�ݗd��
���&Q��b;���d�=o{ ջ>�1�+�r�Xor���hi#+��w]�������ƈr�A������#�m��,in�j=�7w�_�(.D;wb��'C�BGt\Ͼ���kM��h�ǯc��e�ܨA��UZd��/E�1�o(���*ouj!�n����h��"O�85�P��Oq�r���%���f���n��]��,��M[��J<%�N[q��,Fݨ����dU)v9gE�3�*��]�j����7�v���������Fr{��r��R�kJ[^Xg~N[�*�����Ŋ�pp�D���v�"QM�V+����Uvj�M<��\�U&^v����
�6h5)�y:�Y��r�=J��ʙ�m�w�Xz�u���&#d-��WW\�r���֥+0*{g�`�+z,
�����ʽo[�<-����� Ⱥ:�Y$O�i/��������{"�i�ۡ�8�F���+��]�$��B�W8����ob��o��'�p(�Gs�Rp��'ڭ���i��<]���ݲ��:*�O������5ڃ���е�\�`�L��&-ʹ��#	,�8�g�n!Vz�%@V��p�t���B�u�A%&��Q2�pY!�r��X:ʾ�ܦ�ck�vʪ�Uk��(e8gƷ]oU��tӧ"�������D:��e
���6��\]�u`�Y��
�+2oe9e��m*0}}i�Y�؜�Ē���R�VS�*�휨�ySkmZ�ʽȐ�UMu.�ôc��B�a֓(^�N��l
�j���R˧�f"j�6�u�����r��Æ�w)Z�go1�D���'b�p�5S�E0���WR��u�ۆ1�/�֣����]���S�"�����D�
Ź`��M���:�Z��`��F�R�c�Ǒݚ�I�"Si�v-�/h	���l]J��ޤ��##��WZ�z��s�-tޢs�
}��J�a��i�]*��p띄9MN_g
����[�PvQ3t���s�:�УF��Kr���;"�D�Ӗ��¢mvϩS�"��rߒ���R�}�[�4^8��ɇp�6핋���'}vW�m�JZ=�(\W��w�5�������蘗Z'Zዘ����zv�qivm��/l߇;e�nm͉�8Ցݷ��#v�)�x0m��X�čtӝ���XŁ��Zoie�ݷ�щ��b��}�_W<OTdQ�W)���U�}��;������Wv����s_}�Ɏݭ���#u�����&��������s��S�
�&���5��YB���,Ǔ�i�<Xx����ݙ�+���⬥�`LU��B���� {YuGHjVEgP�[/$=;�Ե��e'j]�T�rw
�f;Ӛ�)�O���(��v撈�RT�k�9)t����:hNZok����9C�R����W;i5�*�_C���c9�8�_Ni��M6���� 	��`9t8��vEm^|r��<��ِ�	N���z�;Z�tf�9|�p=dM"��@��Ź�Pח�+p^h�n9r܈	S��57P`!*�C�r�l��"�>�0�CqT�dô�7#ma@]�r��d�4M�A��g���k*�f8P>�}A "�E^m�]�Y�S��_w���ם{WY�V�s� ��1�]�_r�y�f����Z�Su�
h�J����Y"������v�U����r��:�Z��5n���[�~�KqD�W�����a�U-�*�sj���6��ǆȠ�'Gt����t���:i�zp"��VZ���e4�5OhE��տ^�+S�d�@���L�Mv%E�v�{z�;���|�j
n�y��6o�W�8!��&�6������EW�̌u;�}�W];�FS�j%ysK�)�O�]��>x�[�o�԰"򬢕`�����.뭰Ĭ}�0�;���*���|�F|���76�oi\�\��
��n�t��6��
���ᠸ���dV1�,�L�(�R*�p	bۼ�����h�9A74:�5��OL��z$�[/��ٹydb�@��f���ЧR�"j4�vCh��+x~�]�.�R�-�&�=SLG�b�	��:�H�ǂ*��]���M��u)�ٛՂ��J����7��fb�x��Q��%|�"/@��@������
{hcy�M���:[E�J���`X�i�=�E���`�wr�QQX(+��)��X:uV�#}�:e!�]1��X�ö�K�V�5ܾs���c�u�+���e<A� }D M�X1�f_>��W|�Ǽ�m05N�*mh���6;��*X�bd������.�M�ѝr��n���Tyە�A�SA��=YǻK��[C)@���[]+:���:]���;�\��)S7O����f��Kngfõ�ok:���*Jl��O�@���$b�Р���w�;{Vr�{�ЬPQq��(v�bӐb�֧!7��(����s�B�v����=i���ƳJR���t�9b� �H೑���E��3D����J՝h;���<�`�N5!�������7�\N7�7��=k�1�LNy��}?w�DI x��k�z}~�U�O\}�{1�<a���s�~,�v�眔�F���(�M/�����֨8�)"�(	��*̨�E�hӔ>�����H�㷉g���=h��+/l�虸�G���/���6��{�J��
V:ɮ4HG"��zfT����\�eb�D��S�x.C��-B���lԸÍ�W�R�k.Z>�a�yeoF{p-����÷�?�Y�Q��l�5!\�6�K��vĦ>�
m�}ٯ����X�ڒ���'����̝f�w�]6G�U�R�m*%HxI��KK!�Oj�e���.-ؕ5%��$4t�Y��Qc�.!-b �,gc׽�:���O-lM��;#u;��usw��x�3����5bKQ��ҝ���A��;&�Ӷ�e�yS2ږW=!1����[X(�m��ͭE�r����.��:/�+���ٶT�to�+�2+�{�V[�����jV�杩q� �ovB�\j"v�i1�9��2���^Y�6=��t��v��';��3/��W4J|-�Q�nV�wÜ�wڗ<��4GՎ���6eX�U:6�a�p�;�&v���+�z�c���=z�b�h�;��}k�P�/Kk��w����i�l�Xv�%h���Q^�̄�$U�(Z�e���һ:�kz�۶������.�P5�����-�Eb����\K`ue�}	�9���s�I!)Y�A��UM��:��C�8Je
*V>e��~��I�X�E6tX@ � ��@�e݅���*�i�I�D�@-�����K�L1D��q��ߌ�SM{6��1l5��IF����EQM��0_��;OcT̳Y���}>ߏ��������3���J��Ν�C��S� ��h�Z
v�PUEh�1��~w<�|~9�Ϗ���������������45[�*��b�m�ɭ��Qlb���M�����O��������Y��~���?~8��+�z9�������,ly�QE$Lt��<�U�w���=i*9,5݈;.4��=2�W�:�Ʉ���n������֮����뻶#[e�i�v��͉(�dZ6�� 6ŵ4�Uv�]ݮiS�7wUΡ������CF����w��+��H�c��mJQ�v:zS-�܇���jQQu��mK��n�Rv�U-]�2���V��͎�;y���'�W1�0�k��,��`Ʀ��~]vq9�66%Q�nߜ���������0k�����լӍ���g����M�u�ݭ�cZ3v��+ltb))�vεc5WF�j	)*�gASy�;j����$���檽l�w<j�b����C�`��v��ט��Z5���ƍ��*�?��SLI޻�w�>I�>�G�
`*����J�����z�V=��c�%���h�v��mq{���vkeݓ��Y��v_�?&���4SE| 5M�����}'�z����(>;�^Ω�ͥn�l���+T��B�� �sh��;'��v�-j��]�:���tzz��F�ע�j�v�HQ��I���9�}�.�P�N�{�ƫ�7:�&���u}ѱ�0EEu�Nkм��Σ���goª�I݉�h�ù����ۻ,y߰E�Һ���+����&���l�-*��k��R��v��<z����Iܳ^��+�{W"[�x��ʮO��3k˚�>�=��p����>��7��7�6�����O �z3u�dnl����f�w's��;�-���=��G��]Bd��t�x���OM�ث�d����{��g�c7����2GV?���}���L"��X�(�V�=�k��(�@��O����:K����;�ٰ'k���7r���
��m#������<���o���U*������m�C�n�}�}�uϚ�a�sI.���P��^Qhlye���cZ)寥f�tX���Jheo]Q�f��>�N�Cח(�ڞm�J������4k�����<6A�n�4:�|Ps���4j��ǁ� �DL�w��0ч�&u�W�x<B��]ڃϫ���9݌�׷�{��Uκ~�j�e��*ygg�KKމyv��ug���u��R�}΂�V�C�C]l[�w?y��E�����{gM�U�pz�힊�o*��1k��P���|!�k����`������}�������c7o4H�5�xn�r-�[6�Y�f'�݋+�Ws���_ԞuMF8�T>\�h��'c=Q��L\wM���w�{B/�*Z��∪���U�V�ӳ��W�����u7�_���k77<yH�A�ǫބ�bs7u�ŧky{��T��>����v�$�^���ϫ�Z�w�&��Y�a#�]qF�E�gʏ��4����wg��� ����z��_;�H�׉�x=P�p}���������ct�ݑ�;Fwd�z�wOgW���vu��g��=�����Q�R �`xj�5{�7X7r)��R��Z�U��k�>�p�L�0]�4^vR�\����2��;L�����Q��޿����a��>zk<����W<z����mEm	ɇ�°A[n�^��Z5ѥ�ԕi�bʮWZ�Ι/�-u�r����1�/4޶�����g;�������ϳ]���Ә����U����<ZFmKW��x\m�~���3��֌��W���5�-3�v8��0��T�V��f�^+�;�)� W_ݴ�x�ʩ��zry��u��#�1�zz�7c���K��/���`v���1�7o?��tm}�g>�%�*��S�ݴ=���F�pU��s�{Ԯ�jt}Xj|�B�Kί{+����T^�	&��6�V�Э�w�V���^�t�up��}�}hf�.����l�{I��C��}�;�/.}�^A�ۂ��4��Gr����ʌ���~�n��|tA랗�0÷��GE]7����f�s�[�]�}��zߏ4����eX^��<�0}_yTiX����TwY���=�G��A����FZ�]����g{►fy:S�'qɪ����Y�}NZǭl%�MOM�<[��A��2ϼ)H���櫻����>Y��6�Ĵ���n��-q�.(�q��Z�~�K�&�e�դ#���0BF�Pu5��j�5��M{�6uR�]��_�YX���6elҲ���i1=ʱ�Wо�'}�i��wR|����bs�+<��-k�5
xU^�c��Gu�x�l�cY�����~�n��-`}�,���e�N�E�q��Ǉo�9@| ?|�������d���=�+ޓ�k�����s�^��;�w�9Rx���!D�&��Y�+n�w/w����V�$�K2��t��������{޽�!N[���?]K��i�^�=����kqZ�}#���V��j��R�Ta[��q�~�Tz��Y�3�).��I����/�x�'�Im�uޫ���A�y_���P{�rVzv����5H�ۏ6��Լ$�~�7��=���^�rb��}�d���t-�7C�5�og���$w�m3�ñ�o
>���5����D~�vR��̟g�-�H�Ȋl=ݜ6.7��vG+��s��`}��y:Z=/s�eT� �.���
`�� W��G%Bn�t�3�2,����㔴�")�6�����FB�դ��w�J}�g ol�(�d�(Q6�M+'	 P�Ki &��$4RAVhСN�ڽ��ۄ�����B����C�Ӻࡲ�l2#s�wDr3G����Ox{��n�1�/o�9��tw],���&
f�R)6�Ҡ�������j�}_2�����'uK�5�����]{���B��G{�<�5շS�WtX#���.{wU^��N���)����O��LU�ƻk)}���>��>*��4S��9v{���#�]���nl�*�9ʿ*��k�\2�<xb�*XL�!��쯨����G�z6���>��g�>�������3�V!|�7��j<��{����z�Cr��}Nu����2�-��؜ƽ��6�rj���.���oJ��2�[��=�>�]G�d�ޝ<uD�W��_�\��u���v^\��ː����^&�z{EN:���|�s��]+���2����8��^���f',uo�{�}�}�k����{��{�>ۼ5l���vQ��DRIPB�40��zc��@ޚxG�:S^��V��� u�oa���Z}�{lw{�t3��/xͯ.p�g�O����븾
��k`Ʒ�#ů��v�m��7�@Wn���Q,����/���Z�����R�,S�]O�[�o��C��tF�U�wF�Pa]R���:p�$�gb�i���0�
�6�N�����撫*!�n�;��5g��$N*��*�Ȳ�ɽkr��F�}�|���:�����{X���Cc��+���|�tc���MՎ���-��恵���}�r�"�_ӷ����{w��vd{���Ȇ�;g8L�n�y|�q��Ü����ק�bv�Gvg]oC�j5�{��ZN�n���;f���v/���io�%���7W��_h���7`��w�w��&���Y%���|�me�Ϯu���
���}��J�:���3�&w�f,�ft>���ݕsj|�(S~�U�~���(�º!�]���Þr�n�um�@���wk�iϳ������42�_�o�S+� ��KO���ﳤT�Ұ�&j�=�ϫ� J�^~(|s�ɒL������퇋��}��[3O�#��K�p����;I!d���w��O}�5���-CM�0>���w�獙��W�sL����
䟣
�1�x#i���Ǆ�Q�zm�"���ۀP�eܒӳ}�s�+LJ-	@�C��=��6�}1��Ր��:�AҞ^"i^4;;�wy��e�qQ�J��I�c�]X�Y�W_I�?'��:o[�wj�]���-�����s�%�ش�A>�y�R������U��|j���Uv,��=�q�96���~+r��6n�F����xy���U}U��U�,����-��&����xz�I��������s��f����ϡXӿ�}��t��8�#��:p���,������?�;0��oG^V�p�{�/^ۊ��[��w�S��%�����W���[�==B������]�+�'yyJ������V�yץ�=^�mZ��+GJ��뎩x�u��ρ��޽�?z��Z��{����۫5Nk�YP}mW>U�M���	��sC���Ak������78s�^��z?�m������]��}�Nڬ��;����[~�^;�rs�}]�>د�cg>�ul�4�^�{٥��(V�<��/Ofv��d�{�^�*����E�~�;��u���ώw!E(�Y��i�_L�3�녂�p��C�{t��Ңs��^+�c+�wV���$X��![����*�f�	�Gh���
�T��&�T�Q�Ы���c�7%�$����\���DZ38��92M���e��.�*���R�\�;{;��~���IL�� ,CW:3W�w�-�=��ЋmS*�.����'�w�X���C��h�uS�]�uu}w3ӲP���u�{<�-�)�tg���@5�����w��U��#֗iU	���/�ɗEs��ͭO��{Sz�^�~>�cη��*����X�V1�:��3�{#���v�84���^�u�h����{S�o���hm�"�޼tx���]c�'"��֌��I�Z9�v:����O}r[*m�ޛUi{{�Ms�����v{����]���Ɂ�� fwd��쮨�=�M����w�\��/B/�����b��f�_�;�74�g�m��~8��C��f�-����jh�%��0g�����-Y���l�S���ܰq�ּΞ��G�~���uC��zv�Bi�]6�m
~��3 P�'t��g+_��6H~������ZM�������k�@U��b��[�Ysd#8
!�<��;+k�x���z�'P_�dT��:��U I(p�	�H�}���(��F�7��!�X�H���W!���E�v\��9k�A7��Лʴ����+�O��0�A�E7mK�>@��}_���{:�����L�Q$T�{oV�U�b���{��9�8��½h�Z�������Ww{��q�3÷" ����ݻ�73=g�֡ꔨ�~��~Z��)��<n�ߜ���ٽ�E��������ήp'�z�Cy����ޣ��(u9���kw��[�y>��Mwڦ���k���,׼�""ݧj��V�.��X����|���\��j�-�8�.�Dl�5�(���o�4߾^x�:���ư�qK/��b�4f}Iy�����9��D��~OW���z������@=�o�	��臭���k#)�^��-dM�켬�����O3W�.h����D�=ޛ�����w�oWm4��=�+�Ow�R� Q�+��Q+$�����J����z!y��[��w[>�,��~�ރ�݁N�lE��y(�q��T}��7��t�H��|�ܳ���S�_�{z���������C�0�z�х���j�i��b��H�6��$���F��w��׳�V{}��L���s�N���J�,.�`����;�b��qN6��4gw�u �{�����wܜ���W�Ff���u���"!{�����W���V�������w��O_���N��:�K�%K�]��Y�纍9����<��)g3)�ԋ[�������+�ͮ+MR^;c����2��������9t;{⬸;��=~��T�z>Ǫ���:��_��a�X��{����!�;��_lG�?.�g��{�%�{��k���xJ�n�����hs�Vh�`�׵�_���u���k+�����D�kH�΁�ٛ�ۙ���+��C�8q������贺	����4yQ��>��?X�����6x5<s�L�K�w��|?{�G��K��y��S�����b7��}��߂��B�����_\/����v��:�F1����k(}_�⇖揞�a��r){�[�\h��;6ӡ����Hm���|pXX�[���{��x~[|m��n��"F�5w�c�lj���C�N_�ƚxe:}�y���+M��c5�.��淟:?�;��a�T�F�.���:�L8v�Dlt�]58F�4��;;��%sJ$��n^����ݬ�i]���(-�{���[]ݕ���H;x�����j]�� �óL4�N�X�+ާE��K>�r�t4��40�>��$ܤ[��@/��*��A��봭dͮW�{[�>,U��D�|P��Dm\\���j�6kV����D�Vo�*��~*<�ʴx���M�oq=�@�o�M�|k5��G7�.U�R�6���)˪�:�m�{���ʔ�����b�����JVpe����2�Lp��k�,uO,3�k�}Hh	��Y�����
��)��9��MS#b���xh�KȁB^��@[cm��w5��#jn�õa�Hu���v=Ju�o�>v��wb��g.Uӭb���3��H�}g��)���n��ݮ:��ʖT�v���7y��\3,׉�q�ɕB�'F�X�.v�;����:�]�٬=]�V����u
ڊb!S�i��-��<y�z�no<�]*ᾭ9Q
�ݫ+�M�0�݁�Y���� i�G7�PW��,tr�@:ɰ�e��8�����,_�k�P�K��(�{8��S9S�4n3�٢�I��c�~W��6�1��bɗs<�np�b�*�Q�v:C�:.�0�	4aXg�0�p�pZ� Ы*v�D��-����Gv��R�m�5�ʛ^A�l�]Z��!׍��ǁЛ��T��P+����(z�\iv�ؑ5����Q[s��톤tu��)-�xdi�X��p�=�gj-NS;͝n�I��R�$�R
yY]|un�+��c�"����1�C��.��dԱ+�\M`����� ��9�����>�I^Pk�@�ge㾶���7X&�5kB�en�J>H/�\���V�)��2�T��'�Y����D�8��%�7��Xk�lk�Z	3=�tw"�_�{�f2�-p�^�l���>�����SsAͷ�D���;EE��y��W���>�L��ou*��5���[��ڝC/.<�X�:��|�U���4�rf�j��<ɾv+k/���O_6�)�B���v	p�ݜ��l!����ޡN�Tpq��a���y��O�m*���E>4��Ru1]Q�}AWQi־�����BK�fΤ��D^M��iQ�2�1�P{:��.+��άJsm���me���i�#L2���}"M]��⼂�m��w3lQ��i�8!㋇+����L�'[���v"u�@�	�b�TقV��2��}g\i5Ґ��G:�+�U�K�Oߙ��V���SZ��wERS~��^l�n��0z�h���RvsQA�>�o�>9��O�����~?����y�?*�d�Ս[��S?�i"��=؊S���|#������q1ъ_�^|}<�O�����~���3���ԓD��i"�������tQ{�MR����g�}>������||~������~�T��O��+mQ�Ŷ�lRU;bRѢb�h"*�*�ͬճ��b:3��D|�tt<���o��T�-D�Y����;��kX1�:x�-���]b�wc�'^GED��tSC��tր풎�T�3$M1UT�A]:^�tPh�8�)��������1m�������:
�i� ���l�#��D5Eh�֓��5C��[� �+>Iv�JJ��v4E:��-��T�Zv�����㠶�����tb#�c�CHo3�> q����@���K"�������lta��p�9�bv��յ��u���绳��BƄ�U׫��¾>o
�iX/�����k����m�g6�����G�	
*Q��@���@�A�q��M�o�硳��f���nn.^����V��]�x�y����@ێ9;��y��!�\O��0�A�ir@�Q��\���=ٸ�g7�9�}��lIi�O2��py�����!w��L���'�w's`�M=u9|5���q�2�R��O���6C8�hkp�N��y�mHF���~��)�p�`����*!�U�����{����M2
^}6�ݐ�@�z>wn0�\�����ƚ���8�j���Ze��|����ε]�������6�-N��"�Đ�I�߲xU]�爠%��>��I���}p,�]��Z�OLr���(��;f�xydP���մ�ד�V��yM�j<$�򋶪��	�v*d���֓c&�X��l$=�2�h�ކ l�o���|>'�a��
��'���1H��R�,�3�p�[�|!���!^u�K�i���쇅�<y�l�S��־�4+y25�o<�<�#��ly��M�4i]��Ŧ�! _�<5z:�9�o	�����d,@�^��c�8�ϼ�~��6f*T=���O���y��)���jV���}���
ȥtׂʋ���pj�]���®7؄�oռs{ukw������"�{�Q�ug���`���/���w��u�Ӻ5�n��b[�@�'<�����*�3��ߛ�������?<�/����3�>��Wn�ڮ�����p��r���GH���Ф	~��!���ձ��3�_��S�N �6M��!Jͼ�n��;l���F��{z��/���.�X,��Y���0ь"�hv�&�Yr�
{6���t/x�����'���D]k�?�W�]}nWzpϥ!|�~i�t�l�X���j-��g/xx����0��6Ӭ}�FRl�R�x�O,���!H`�!�H a������̚�uW�8��={<�<�1J�/�$2�R-ǭ)"}�s��n�>ѽ�0·��#��.;�VuNvһ�̀�\����c�7eCJ��� ��u����d�H�<�ѹ����1��^�-�؂����j@ nX;(޸��P�C���q�œߡ_S�3�%�Uh��5c����m4�tp�}�����NMB 
���!r�D�W�\
 ��U.[����i����]��p���L��
=���I�uz��D����个��}�v⁨�`�"H��Ѫ)����Ɖw���J[�R��[�D����;���r@�/�ԚO�N�[Q@����)�*��jw��2��`���َ�"9�*10�N
���+)�e䜅��y�P�^�7yF�
�e��v�`]�i�Y�5 �(�p����fέ�r�P�\[uwuܪ�ąs��1�EA���2��\��	�0��,7�;���cO#ޑ���SN���%�b�6�F�9�rz��WVM����׿E���[y���a����������]X���2yV��ΠD����n�vu���7Y�*�S�}�+7�9V�x]�|q%4i��YMy�8;m�s^)k�[%����,�vSd<y���E�8ǫ#gIfQ��|�/w�e[aޖY��w�9���@t��`�]��~�Ʀl#�C��~���vz� ^��/|�v7`��>n�̡}"W�S/��A��T$�	��dd�T�Ed<�[HLM�(�m���k.�*��jDd�\����r����2�dF���c����_��O���߸���.��������8߰~x�GnлA��i�{tgf� 	z`3��yf�]�&���a�eF����ǟHV�}&�l�ݼ3�Ƃ6j���L��קx���� �����{��O��(�o��L��|�$V�" �& ��Ogj����� %eF���^��>�?����Q^��v��÷���׮�N��}��
��Z����7��d�r�l��3Y�w+_2�a%
OE���A���3���1���fy���Q��@���`�)��>�y���ʶx l�z�r��-�?	G��@���@o�F�i�$�� W4�Sa�oEs�be�����Eȇ븳h�dYD��6����w/zRˢ0�*V`��ϊ,%�Sx��w������us{X�d��[����.�\DI��;���L 4EV�F��̖�byT��K�lg`��&-�o5y(�O>�|+�𯇈�f󧺡�u���a�aZ�}�n/[H�W��I��]���c)w�8-�����5M���T��ɛm��C�����o�"��f>�i������%.���ӭ�+ϮK�9��)��M���ӧ����Ƴ(oI�o^��Q��恖�y�i8�*�k��7�H�r�DE�jtL��ux"j���>���ર�.����E:~R�>���ހ�
R�m�ͻ��P7���[jzZ���E��Y�Ǚ��ަ5��n�j9��Tx)���N�Lf]�7>6��i;��]���8G���D�+�ځ'Xv���M��I�2��;��S6���D�P��y�ɮ���^�"�����q�^ޙ+��8s��E|�ϮMY�O>f�Η�w�Ec^!����f��ȴל[y ����{S�i�x>��"-*�9�@sB����'�h��bE�|��!?5;6�Ze�n�1��'op(�N0��Wl�5b��ϼǚa�98@{e)X�j�19G;b���%������X?7�f�?��[ '8�X�� ny�>�S>;�u �������,7@�ooZ�!�,]�_�j�F�W�7��(؝������`V_(�>�h�6%l;KV�q�����o1�zw�)N�Ԝ՗pi��>�m
`Wf�M���9c��Qs���6�Mv��� 4��/�K���.]w|�~~��ͽ��3����߿���>�/[��?����q�y?<-���o�?��}zy3�p����F@kXG���"�ⶮ�Gm�k���`�@��^P�;�]pM�y��@�Ok�t�l��E˜9����s�Y�0���./��"Wg7oI}���{�şH��%�tY�o4�� ��~�1�ހ�[�\Z�
4*t�1䊍�R14�xGSΧ�Dvma%5(G�޷���ǆD�ϟ۱������m�3 M��E��Ӊ����b��ӄ1d���������L[�f}�}!�j<(�8��}�=6|�G0�HqY�K�s��FV�����wc����>(�0ô'���'��{DF��桶y�(��� P�%��]�P����Kj�9A�]�0Pfsq�Ԙ0!?xz j����p����cs��gוG�G�/�.5l�_v��FJ$YISG�u?w$����!T��jU���G�<�b_�}��arG�rIETG;����Z׺��;�m���:(D��:�'(m����w��'�k�@v���ddr(�u'�iL�J��U����e���4徃��s�Fs�_z���q�]��W�s����rx?�V���z}��ҟ�-/���;_�o`xXs�2&���p��
�(>ӭ���n��acdh��M�9�_!�̓�������D����q)��sz�K�r.���ㆉ�kB̩EF�b��+��:��3����y�������^�7���_<�O�Y	�7o~�wUV=M�}�����I@��um��[V<�����g�~�1��(�歀ld�s�u\m�	����ʮ�K����c�|Lz�� J}������:;֣�k=Jl�7x��8lv�����G�j��Xޒ�ܖ��
MI슗g�#9����s���^�<�(�3\��5p'���,��_r7��jB�	eH�ه"���5�^�u>נ9!����ɜ�cu��.Lhmk����	Gnn̲�ۣɟۍ$K�ٹ�(1��ȒU8�!�7w���g`���>��K/�Nwc3�-�o>��+�,Q��G��_~�����$��9AQ��S��o�bc[e��-
�V��]��[���#:4��|��}��\���~!��h 0�KI���ύ�Q��;���Z� C\��iL��+1�0��G�=>ŀxw<��z�]i����5�yy��f&\�k1�2�ᶛdS�o���iN8{yԷsq������[�V�-�x��S�OBZ�������8b�oZ����9����<)�:&����:��2 \B�bm���V7�>�=&�F!�͢�W!enՒ3�+�"\��x�����ٍ��}�bx~�kR�:ฏѠ�׊�m�w��S.�uܕ|�li�U�%�����RByd����=׏�!e�=|�b�i]^����G@B��J�@�Pt��x��S�[#�n=q�����^W���^^r�;�l��l����i�6tO�H�Dy���5z�w���T-��{�RuUwn]hn��TV����>ǟox>�*�c�D�vi����Z�=�&�-��u�u}�;���@a���K����ө�9#zZ��ת)�k�[u�����_x)eɔ���Z���O�0�-\YT*j�v�<�J�M��"yeC;l֣y"�!O�H[Y�œ7�Qm5 �cx�9�ڛC������d{_���V�Fa���D��K-sml�%���9
��V��=ce�۶&��xQg���݅(�t�}l�32�~sk�v��M�y�2�P���i��$CS��,����y���	9{>+��)�ow'b�`�u��S��<�����l+꡴#b�	�-�\C"���+Y0�z��k3;B���Dp�V�j�W�C9�m�	2�Ӊ?[��XhƦw&sq��0�<,�����!8��~hMO����oJ�#.�\R���U��;�Y�p����;����IT!-���a�Fh�޶������g���U����ӳYz��}E�X�ƈ���k���t�en�enĴ��v�x&�iƽ��X����v��}J��w�w.�IX6�O��5�+�3��;�B�΀��L9k����{��u���ÉE��������j_��]��J7�D�C&���au�8��ڶpg:"������U$:��y���8��,�%�'�i��h%D�Ο#�L'�c[�q3b���^'����r�Z�2;���_1�2�J�*5��ྴ���������D�)l��ǧ�:�N�o>�����zS#�*|Z#H��Qj��~X)]2�ǵu��i�m��L��z+��g�w\Y=��k=UEڳ�u��!�!�fb��P5��blia�5�4�`�N����l'[����B�/���Y6�t�uB�����V��#S����㽠���ͣD@v��H�zT�l#i���v�����lS���?s����f��5	�]Ɣ�o^=�L�=��i�3L�����Fzw�ay�97��÷;��������|>���a�2` ��`�i����U�x��q�U<�i���e�C�ٹ�۷�-���I���0}��w*f~ȑ���"B�	�1Q������E�f�*h͢!�]"�kI��]��[�T���WQ.nv���� f�J�1p�F��7�;+�t�ATE
d��a,H����L�'�.ƌ���gsq�����ǅ�]v.�:�+��ɖaYx9ŦuѪ_���󞇫�����^vtCf��E^y)��V�Eg�l+�")=l:��h��r8Ψ�Ȼ����
���&�^�@��Z׮�̈зjQ�O2١\Y�݊7#�E4�H���V��^=n��UN����O���ӎ5��=�>;�ލ�ΊM��m;(�f�5]jFyR%\��i)c�����;�a��3�Ti��V���\�SPd�mH�p(%A���-��~��;zـ�!l�֟
<�f�8�a��DwdCfת ��A�+K���st�Dd�fr��h�҆42I�K�8zB`\�pM�a���y��4�CF�2��45���q�=�.n�Њ�����>x��g�{'�G^���-���5���`g}��(��-��}SݭJ����$�Y1�n F���&<��.���6=Go�)����x_QQ e]���~��1�ţ*hkv�9�� ��Îk��k=i�X8⍙�}�]��:Y���g�#r/h�p�]}J^�l�'v�,0��YS�r7���7�.�ϙ]1�Xq��S��v���e�v�F�E�3��+���!J�Z��ݶ��-Tf�weG˖T�[� ��@���;�zs�3iY�w�R�eQ-ԧ*yBp�ҏ+z@O�+��]=F�k���/�hF������3�Q�� O4����Hg<H� 7w׽�Tn'�Z�W�T>e����ȹ��]����1�7*���v9w�,^�;n������2T�@�	A2t���Q��H���g��F�@�V�x���*��8��k/��y�EA��W��m>��6����V�?x�d5<�W,Djzwx��z��ݨ�r�3�i����Lj�ڒ�ևc �Æ�
��<�r� �̜ĘtN�|N�9^L�T�]xK_ˈ��ԡ뱺����dS�/U�!Qn��f�,�OZ�-6c2����~Se�ɎH���ɤ���!9�E��l�lӪ�0+|����۬ k�|��P&��g.�q��et����]qp�����-d8���79M�O��lk�D%;>jã�GwI �9;���%�f��s>:z��^JGT�FR�k�@�y�z��N�����ȶr�
�����+�i�R������m���c��ٹ�YB]�38v�(�^��Ω�C#�Pl��=����~ˁ�2
t&����N��Ce��!�'��ϛ��y����W���[k��E��~D�=���+b�Mp�Cy�3-�nD�t�}PhWjuGʢf[5|*
]���L�.��p��W���끒��,U�ܬ-����>��M��ld�B���sWY�7/U�Q\m9}ҍXf�y��|�u�X�+7�%Y�5��n[�O�,*��8}��SN���;��o`����^t]��0<��Kî07�`�>�+��6�ֻ�;N�m=��Θ4�wt�,i�"��±ut�c-���kLۑ'+p ��nab�%���A��UjV��M*���̷MI�2rzyҸ�����[&�5�nB*�dr��
ά��X�k+�j�W�(�{b��#Aκ&�=�6�e7q�VPHz;��ޛ��XM����_�r�%]�S���.x��/�$������Z.K}*ZZ�7�mth�qY��R�I��f��&�#	�p�*�N�nw>�zc��oU�WdM��*�Իj7�]0!(Q�],�ǩubǂS���1�h4�L�g]nh݂� �E��u=�g�Z㜋٘���N�+(��ѻi.�`!��s'�zI�-��;���G:���cv�@i֓�[n��Yp���=@*��c�{]��K��Þb`�p;�������.�nb��S�!8\(Ztk��c�^���`*%�:p��[�^EZ����P��U���K�B�)�}۷��#X�,:�,'G�pܝ��q͒�Ƕ���x��b�����C�U��^�'���>qg|+�����^Y�]�}]K"��K:����L����������@a��Vn�Gz	��ȓN.2\��0ԩū�� �?[ۅ��Wf�b��ʲ@N}q�u,�z���5�v��DS��0������ݷ�K��*�ܶ�����Y���y
��J�=q��\t�'��t-����;��0����T��q��T��n�A(&jJ4�\��a`�����`Җ�ʍT�`������H�gAŋ�\L];nP�4s%Ԓ<x__
2����NǇ�쿆����v�7���?1�ɣ[u��T��~�*ǚ���tj����pES2>���Ѽ����\�qM��C���X�HowJ0�Wx��t�7.P����mU�]u|+��e��)�zp*�<���:�Z�}�܎�0�1,�<ySp��V��ޫ�gy�lEɮ�2`�h�;x�WR���+�fnQј���;�0���\�L�ܭ��&��;��+aH�9��������ƱU�]���_mE���,�0�,���T�X���*t���g�ek�mX�	��<�1{��0eԬ�Ҥ�*S��`�L��K�'�#�{&ܖR,�^Z�/K����T3UӮ�0v�w��M��`��e��Z�mRu��A��fp%�C��T�Er̂���*�2�b�H֞��\��sf<v��Z=\fC�B���@�@�'RC8d�d�b��V�q�'7C�R)]�q�eR����A�ŗ����Zn�9{@�6HwG�Q���`J'4��E�*�e�-yszNS�D�5������Q
U!�!( i�� J�(3I�����K�A;��BJ	M���N�H�.S�(���P�LVLE
��A::f��������c��������f!��~�{������y=�4�l�`�n��Ed���F�(<���3�Ϗ��������}>?����?���]�Q��r�bzր�PݳFں��48��o�}<��~�?_�����}?G����?�~o���E�&��cK�t��1D���RQ�������Ϗ�����}��o���~�_�s�������l�h�TP�UQ�:`����V�z���I� ��i�,Vhj�i��bո�T�GF�������"z�A,ZE��HUICvtQѤ{��ATi4MRUM�Ǹ�z�]�ыn���w&����wO�jj)<����Ӈ�vn���tSTcR->�`��Ƃ�l����b�$�mlY�X5]��S�k`��:L��݃MM�7��	n���]�4�+I���C�z����?;�d��Gaã'l]�{)+��
���.�}t״^���]Y9��iP������â�����28�ʮ��7��o,S�w��o[m��Ϡ���eO=O�_��x�����T��j��e����ⳠL�Q�o��oY4����[���!��u߿dx�\X������� �E��̈a��m�4>p f?&^��g�`>{#�Keyi׌k���K(s�)-L��6@�k�3��<�_8;*n�S�� �#	θ3_��P顼��1QT�u��v�i�Sy8��g��K��8�����=��ࢬS�h�z�y���` �7��LĬ9�^B�����C����4M��͝,�	��B{!���uC�P����O��&�k1B��N�q�o�a*�>i]4̵�u>hƏ5t�4���
�T�u�7j�c�<��װǫX:,�ݛ6�Û��)٠b�v��ݝ<ެ����3��r ��2�S�'��%��Ω�ہQ�}�^�z���gő�*��c���uQy�'�����ݒ�c��F��a�,��$'��Mᵌ�ɟ^:=�C�������+�C�ʹ���v{wBP�l*���r+�m�����"�6��i���B�<����/ܯ��b���a����Dx��Ӥ�9�?��ߍ��*��f�ŞjǶ���p�vr�[�'�Q��z���@��qTs �pD�Z��3�v&���zq��}�b|����W��qp��Y�͉_.��U�=tQ��K_C��߯>{�����?�0AJSC߿������Skq��Q��U�7�j�b��i��|d�N/Sٷd�f�p'L��gC"}1|��q2TwGCH���sWs�\ܓ�4Jꡕޜ�z���[��Q�h��gj��M!�EN���a)��d<���)t�tE�:c��[t� ebSǫ�հ�O����k�+s�&�n�&���Pt�M�q����n��7���zTmy��.�+��4�M'0��Gt�ݭ��n����?�I�����D��>}<�����&F(��?Z��w�?sY���a��eX�8w#b����S�Ta�lN(g����j渇���h*<�}�r��]���ݸ1�Ԯ�V�؃$]]K���/r��h��W�������y�cW�O��l��	)1y�<�L�R�޺43++���Nc�S�����0;�;C3ǑQ��N�j�ig�)��Q)�;QkE��/F}�$�e��,�ҫg���U�?]�	^Q��]i@��K��húX�2҆+�Mۨ:����4qɫ�.��)����3{�68�u@������0� �I�s���3m��x5�8p����-y�Q�.Gt8���еB�r��=i3@c���p����]���T>z���uxk�k����153c�׫��HlT;;3bj�NY�njHQj�:s��%Պ"������Z%�OK��j!u��UW�cpC.@����S���߯�WO#�-5��2!����'"^�ޮ\m0s�oǝ�2#xA��u=ԝ�=�z��v_i�
%��2	T���f7���_��ž�L0�0%E�M���]�G<+L��ٶ�fF���l�d$��6��Q���	uT� �A��;RyV����=��3��"�74��D�8|�KAU���ܭ{,]�ܻ�S������F��sT��I����w�Tr�V�X`�b�%b�ߨ��5&�����w^S%�V{�f�^)����ȟc�������<ON3'[��zZ�N��I��Jƛl�.+�xb~֟k�s"-&��K*�W��ϳ�(�7A��)��̬a�<�-E���A�M8E�n�h�XKoF�hMg9>�w�+2
|%��>Gf�oS��2�m*5��n$��g�Si�c��K9Q*4�=X�C��M%��!����'��=�̠v7&��6��j���O��~���j����Hx�HՖ;�yAث�}�g�¹8MϾ�r�=X��<����	���0d2��G���[�[�NȰwv����"}d�pR���m5 \ϴ�6Uu8跮Z�T�'c����Ǘ��O�Gk;������P%sϬS:�Z5.�
vV�S^i�b�lӗ�43����8Pb�5IS�C9��מ~�ן��?���p��� O�*��f�\"bV�??TIĜVV�W�5>���g�}�h�C�"�iVܨ�{�S4&�M[4��gj�e�sH��f�>,����r����~:}>�H�꺈c�~�������8��{p��ں�-�����k���=�O����� c�qķ�̶do5{���sT.��wǆqLj�ը��ۼ�Jr���,�۝p���Fߚ��\�q�'2�=���q���-��w۟�bɊ�W^�k��֏�_̲t:%�}�&3��~5��x�����b���.���f�D�b�'�rW�L����.����ǀ>�M'�-��@խM1/�x������S����"'"�u���s��7�� w<�P�^��w�if�i	Ibc	wq�Yl�ɚ��sYyJv54��&������v�3�炍�W2q[���|����S�S+]�UMb�9�/����.-�"F���R�#Yճ�sa��m�)�� I�	E[V�����b���lv�vR\������h2m҆0)��C�O���
V5����ۉ��t��ֵ��*�v�ɛ�Er_c�֜�`U�2d�K�-��&C�kA�FX�kE!�&�T�[j�I�2�:�Ƞ� 4(Q�PR�+��{������J�ú���s��p��]���eX�9f:PT�SNFFUʽ9��Y�3���]LZM�(�����y��6�W�u�O��ɕ!�)�0h����S������߾^��Ĵ=5@wx{v�%6B3��L5������~�Q��Se�}&��2�S櫜��O���*;-חY���a���6uH��������K�	�Za�0)����sc{KeTQO�[CЙL@C��G��7[����M�A����r��q��p�4�Ȇu�y�f���g���^��JP#� V|�O<{5�6��)s�Z��ue�܌{fb����.�E�-��؉]��A��6�9��Kiz΁>��)=���y�o����������b������>>&�o&����1|�~�W�ݻL�K�ÕC��<.�Z�g��[�O�̄�e���Ybv{�J��dt��a;��/�ڰǿ��ߔ�(h_!�_5�σb�p�G�?U�X �ן^*cr�\o��L�"��(-۬�>�m�v�gޔ������>j�#��#>z��`5� S�I���Z�:t^�T�r�6
�x,�)����$��f��"��ʡ	�K�Hֆ`3��a7��BTI�M��v���;�'1l�7��a�m���m�I��Ȇ �)E�T�G���f\�c�]�������{+& ���:!!yA^]n���{G6#"�#Wym:��F��Ӷ�DeP�5�Fe�㥗$/3F�νajbN��}�W
"��T�U��[뾣<�U*г���â�x
%%�i����Kj;bu]�I�4�����?�.P�ҨP+J0�%��~��|���������b�I�U8�(c6�y�Ƨ���nVŻ0�)�J�mn=2����i��"�d�ܝǩ��i~��N$Cl��!&R�v�
��\��S(�����+����p��Fʡ��%ܽK�dɛӭ	GߌF�����:j�=������.���+�[b	`2R��B�ˑV�qc=>Kчn��4%E�7�v����}(�[ו|�[���X�.�Az���^����SY�;
3�y��l����pC;<vD�WE>���W�pK�{�8嗢��k�
���W]�GE���Z�J����||�n�7�z93�.Zeى>D���2���\��Ј�َ;�zъ4�
�Ht�\�n)�����.t$>(�L�?��.^ΐ�kg��4z�@�m��ԧH��8�<�D�Hq���.t�e�o!����U#X8�T���<��|�l
e���N&]�Ɉi��D�����sWhg��eE�����>G��������z��������|��g5D>&�CAMo��4v�-��iq�;���d��pa^�R� �!�^1�o�gU�4U�"�ڌ�ޒ�+8��
���+`�XٵP]Z�x}�P���8bt2�!W!�s��[G����&�r޽ͱ{Z���_p�~8����}Ύ�,��kݶ���a�~�x7�<�x|<@M�U� ] *��|������/�W���߭�E��cy�4�cCy�U���sYT0�����t`�+vo��Ԉ�/��ϸ���[�j)�ن��
���{˗������ҙ+��.���]c��RDu�[U���w������Ss`p�` Y��q|���ɀ�Ohs~��`�7T�_��s�QL��ō[,���*�d.a>q���-���b�|͙�<�p3?��}� hI䃯�Д���d���(@ ��TbY�lbX�N��::q�/woB�mS�3��q�i��f�������*����st��h�u�q
S�c#?]ş���UO��h3�v)�"ⷵ�^�7w�9��²��8��R&چ,0!eC;F��Q&��56���3	����έ�e��z���4F����^
��$j�x+)l��}���%T�9�]���� m[��z�QW��n����G[�s(J�����IL��i��r��$$|�p�*��f��<QE��Y�w6.9�!�aX�m��E�@��~����̈��4��_��?������Uꆅ��O��8��h��e�t�_�w�mp�r緹���)�;���߳.F6�4�����^]��OL�L<Mͬ�@�&�|  2Cq�H�{�9����;J����]�:%�+ܧC���s�_/�lB���C��PZ5j��3h���W:����o���*?���!� Щ�]
$�*� ������������������&fQq��G�^B\�u���V)P�y��[�Sa�KZ����	�ϔ��ü� $�s�6��������fM���h�3��&��]ļ)'~~@#_����7`�eh ӳG�������{���1�OU��]�Y����Xl��I�p��K��]GT�_�m�u�>}��/����(I�n*u�2~�Ӫ߃���r0�C8�o̙�&�e�M}�L�c]K�kG\2�l=�6���F��`?��|D~�����
k�TW�˄R�s
�[�e�m������-�3�j��.�_]�O�:��J���}.�Rxw����=;]+�~��^?���n"|�8q�|�mg�Z��=g[X9��wl>����r�ёwy�{W=:�;�.D
؆.��>�z�MC��[������6�b��镑u��˫w���At���B904(N�^��y�M+�>xO �↿���j�~�l�x� �1L�+Y�s�����C��Hނ{��(���~�f�|$��x��	/M�����m��v�����V�XV�S��kvh��,��a�5�^����ʗĨ�x8X��	��ee�0̺�B�H�,ZT5'�_�(n�Wj�o+n@*�� ܝ�:�I�X��譠�r�U�.��!����W[�����Zd{(�.���h�)Qn���$0C �y"��}�uhfW�"W�Z߳��&�3ΨϿ�����Y_���O�&�b>�
7��ӷK�y}����z�O�$����H�p�I�T�v�2(q��d�%�&@�������d�6�Srֆ@��5�j^5�<��O��/�YgYմ��EpK������W}�d]����|�x��a�d����b�7�ݥ���ܡ�@�{"��a#C����K&����!��Mb@@��OM�����k�_�U��U���t|��0S����8S���Kr�\ή:�7q�gE&��K�ڟ��"���0�0�L��ӏx�~Q�݆�D�P[}�^rO��7I�t{�^K�{]p1�c�S�s��Q/㩒�X�Wi�gdg?o�uj�g<{����+�A�l�+jF��G���VZ׆=�1κ��#]eH����7C��v�.y������˚���S�Z��z�'����*��;��e��Y�]�c���5J�0�^�\�<;�/��7����<�l�C��at;��E��)���F��F%t�6_�<n����iVf���4�������X�2-��Wx;�=��k��`̕�d6:$y:�Z��<*{��`��աV,�7�|��wxWr���0�g#��*Z��c�t����B ��]�1Wf��{���^�=ߟ����>_�~��߇���_��: (2�� ���Q(�$yC��\�"�V ���M�� �ĖMă�16峙��pʛf�ɽ�-P��ޛ�b_cw�LK�Z�ϧɟ�xVu/;��O)Mq��Do����?��Y��NEtd�(.�V���S��91�7GG�El�jm��n��iW?İ��D�� h�IVfW��D��٢��S�Q/ǵ����b��
	��m��M�R{�%�N��ok1�˧��]`���y�S��&�i�f��l���oǝ�S�qqp�-�w�l���T��=kmF��.���=�����;ΤJ��Jg�u����Y���S��"�ga�������[W��T�&��OU�������m����h�ڛ��׃2��G�����4emkR��H ��d�CoT��7,��E&�̃㐔W0��ںr'��Vυ˳6}9o&��Bd@#fj�]��O��6|;��<����[��lGo���]�j��!]܎���g	��J��< ����O�]�ٯ5q�gq���P�X�s�4���4�����9G�<%uP�3�-N��6�o������3O�;��Huf�]�,R�V�ue7b�:����W,b�,��@��,Ԙ�Z
S�5�Ղ�O��Z�+\�t�P1��@oLh	g3W5���!pk����,M��Hf9�黛��e��F��i���ܮ[Å-T[�T]���8�\Â���2�{+v��Q)Yga�4
!�Pސ64��.4p�:�VYe:��Me�$�[(�LQ�h�]�1�Z/���ycw���M�ݢ�)��:m�Q�%g�!��W����0^�E�X�&\}VXަ(U�9���j��M��)���عL9p�Z2lS���f+�`kK��:�L2��(��(�a[���3�������md�R��Δ%c�p�+���}w���.0�A��G}�oZ�:��Vk�4M�.�7�֭��C�u�i>gL��z���I����6�+������]�z.�*�Ź��U���p�V&�U��t��ӍÏF�b�ZJ<�B�����ˍ.�t��ڪ��z�I��x�n�Y�|�"��{F���
�W>Ԣ3����­>�i���vl|*�E���.�^�7m��5/��tl_E�i���WP���e�o�u����C�����3�LA�D��v̔�kI��2��Ǥ����4s�Ry���S�hM�]��8F��mm�I����9�]��4ɻ��Z6��Q�lXt>�j��d�qm��]i Eu1���k�?: <HZT�c��U�]�%�[�Iɉ�/5��k���x.���{�q繊I�7^�w=��n��X͜�,gF\z�
gc�Z�[�X^�^6�î��wX;�Sx��R�O>��L㈣|�VI����Jy�FL���5=z���R��m�tl�.ڇ�̰4��%.|�!��i�mU��=�ɑ�d�mg1�B%U�7.�V���.Y��ӿ�U�΢"����Vk���݃�M�o9��,K�vh�����F�ȍr��kX�#�p�&Q�'e�T�a���Nk��q.Zp"&���Y܀�r=�p�)͡�fr�ТudWoq��7C|&IO,�`�1l��Y�0`�������h��;]�ahH�C��Q��akkd[(��&��s��_:Go�v�N���E4Ѷ�r	k8������}��9Q3�Д.U�X�E-�o0R�4:U�7F�9.�!ǯ�.�[���>�����X�P�h�#8�[�4[<;^Da5k{1��k��/h�GJ��(N�X��nf���v�Օջ �J�Z�3)��yV��М/$�1�2�3)F���v_e��UXnՉQ��|NZ����ָ��V���t���m��
�uq�{*� e5YY*^m.�&�V�qv�3;ubE.�ލ�#���҆�X={�=�{ߟ��߸�Z ��EAQ�Ɠ�Dm��Z�lwkq�+��><��_����}��O���~����~��tk}�8��I��3�LGcR���)������G]�b�֑��gǟO�����}��o���~������툨���mN���G��٢-bi"t:1����U1kGF���@P�ק�><��~�_O����}�ߣ����?�(��7�m�
*�I��UT�Ez��LxeЕAE%hė`ݴSQ�����V=lt�Zv�#�5E4�I��[A݆�w�no0�J(��8`�X�(��Qy��MP�ۭu��N�A�;�Pt��EumA�d�]T=�Z(.���b
� �*:4LQ\Zf�O��˧\[�E�k��b�h�j�cv�N6��M%�
�Ut:h:8��Z���]�=�A��Ol���[�W�;41U�i���=�E��'-��Rw�����V{'r\L�X��i#xr�<ŷ����1��;��&6�8��}�z�����T� 0$B�0��J 
P�������{��?��k<�~Ce�/]�} �J"v��W����Ӝ����ij�	wR���iqr��E[S;��gӎ�Nke�&��.k�y�t��%-�����aQ��F��6 -�u$.Ndn;3?��%��^�ϙ���wM�����q�&}�7�n������f���ن��۵��R�DZd o2�iT-�H�㌱�f���W=������_���.���y񯗶ґ�f�[H�p�摼�_�i�9��x_GG�<�.���ؘɸ�\N�����͘�����\�s_�O��K�J��=t)+ƹ�:�A�~�:��ōg ZԌ��ww���ђ��SX�tls��<R�+J���j��޹�<����:� �Ǚ��m��Ynm^w�Q͌ȅ��}L#�N���ab�ظ�u���k����}�4�lmsƫ{v�U�����&Q%��f�%�\5G.���Ľu�a��\e�v*$�׾��MQ�����ދ�Æ��r�G�ñ��Ɍt�W���pO�Py{˶p��l�g2T��qV3�}��X8�E���M�
B�F��)_f<����5��5�JJ�5��sG�q��w^�v�[�~U{�>�� �B�:��qBU���ܡ���ĺo8Jĕ]��Ϟ��ן��~���UaC�$�a�t*�7��ߟ�O����������~]"<=��#�\=6�.;ݕ���F51��X�1�Ύf$��2y��g�j
=%�:�2+i�x*Ҋ>�J�P�r��[��Z�5Sd(b���jOղ&[U˾��j��̸)ړZ�cn=n���B+-)���֞NO�+�#�MC�ښ��
%�i%f\&�t�/�Ue�qX�t�q��>Q��_��)�wl%4tLe��d�k�Nl�(�5�%��>�V'��N�Ȧ�KF���~
��F(Z��O���Z��ڋ��vf.9����,�U�=�Æ.+\uO����_���� ˲�����.��6�]oF���؇wom��!��<�W�>���e�Ogo�^���0�2�Hx�'����6S6s�T7#{�.�����*1������k�d�};i��@V�h�x���u��w|�o��3=Z���?�L��?��X�T�g8'�����h���d��!r��a�{�n�q0jf���֪!��U�Z%)��39�5�q�i���C�N�����W�eb�o��-1%u
%�=EcIU��o���"��n�4�@Y�U��F����@�W�!u�񌕜Z�&L�]i���'˺�^F��E�D'�0(���WݸhU��M}��,��OJ�r]������Jq�c�%]���׋K��o	SgH��Ӯ�u�
}��-*�C0�Q�T�/��sǔ�Q���`�".R%(BJ ��ϟ�?=z�����`ω#��;�N������8	�Χ_6[Y�_�Yca���*�}�]���������dk��G�ݍ���c�1�U\����v�����X��p����a�=�2��(b=���BQ\�G<æ���|2��3���"��uB����+���ڼ�ٞ�^���w{�+����0C@x]Rɤk��s�2�I�G#���C�/4e��Eşw,�_���FMdy�)�j�V�D�JOӻp�G�b��f)���*z��Z|Z�R:�)����;�*\<j�mB��y��V;�d�+����w�]����ܑj�v|n>��f�C)�Ʋe��a��
��
چ�+[Bkg��8��!�鶯�5�xa��(�j4���'ُg�FG��M���ŷ�d�숛!F�{���1���Q�w���0*�L��ӊ���'GzґW����UF���� �|������LN�u�cFq���؉�����g�w?{��S^_)Ut�����A��G��X��p�nq?_S�V1�%�٪�քu�A^f!CZΆ-BGc.��Yx*;�K01@�(�Y��&��q���g+��l��G
#jZ�9�Ó��|qt(�w(�.���N+�т���7�4�f󳜍��V.��,��('����ЋB�P R��ϟ����W�����0~	��+��
�l�g��;y,vƳ}�]�$;fwk"�N�iqm�*x�۹��~��4�{��F�Rq�|֚ڄQ��8�����e��=���^���R ���v\����XtDFy��CH��W�"�F�sw�$�M=y_�4����ߖ�k��!g�0�J�b�<Z����C�`,ް�v��/�Jn��pU�Uf`��-��4��p"f���z����|��b��k�j�^���6�?��vV�4�ĭ�A-�䧆SSq�C7O�+ͻ�$ft+n:Ec�O0��~�'9��#�,Wǯo�g'*����Ŀ#`@Nq�!��D{<�|�>٣�5�=�⁀�G�%�ivlE���IY܍ٝ������7�E~�M`���|��|�c�w��G01d�%N�z%�5Z��V����/�b����{}M0�L(Ϫ�cR�5mǝ�2��~���_q!�	�9���n�ْQN�+Z8v%�!�T�_�T�z�ߏ�s��u���]�G��������;DH���@��:���<'}�7����ِt�r�0��:z�ⶥf2����k%At`��L�[,g,����|�
olw��g:�Lg�`��_YZ�ۙ��d��X8#ZK�˫�9Z�2�n�}���#��~k�����'�`�He$T�@@>�������῿/}�f~�e��Q�AՌ*�˷4k���n��}�3�S7��M�vV�;��]�R����e֓|�{Yn<�ʵ�1'�a4���K$~�
�ʶ+�{Ƶ͏ϴ�~�<j�z��Փ�F�c�@�w�מ#���T+U�ȝUm"�٠������ވc�KY�pU�L�;���gȔ��Ϯ���.&�t6;j`;�
��9/O�j:�e��]���<�Ӫ�2��m��ʚ��%̂��S2f���{Z}��i��.+�g:�0�ڎ=m~n�G(Q���;�1ص7.���B�������\����.�
Kq��֛h�]+�y��R�#(DfL_������* [ڳ�y��-=:q�݅�Yڇ|e�"!ԶЗ�9�H�Y�3����5���B6.�{��W��l���~"����X���]���Jcdtz(D�&��Zy���4����Q��}�E��)��<;�a�7���q �bpH+�8�(��9���^�&skz
�������8e�hŶ�3_�=ѥ������$x���!�GI�=:u���;W8C��<�d�<�y;}y�������
o���㎰�%!X3!@��~��6$\+�x��{���JU_!�_PYݼ����Tk�f̰�W+���Tݣi�D;R�Jk%��v��R�,����k�ￜ~z�6���z���0��
�P4��� ��?�Ѿw��dc��M���X�O5�cl��~��\���Pf�O��~����`Ha��r�;���v\�Z�ٽc������pÄ[�i�6��QW��i��B�!��rC<��$�b����#��J����~�����s�(�a`����*L,W\NP+i{&�G��#w��˝���ċ��N���K���v7�.)���_���V�#��p��c�]�灘���;Ad������z9�0"�����DQ�b(z*��
��?/�&�y�lmF �xTş	�ܽ Q��0y��}	�UE�d���UZ�p���M�󦬽WT=ܪ�X����JݭR�qR�#Y���
���+�^<��r���Ч��R/���/n:��m�nS���+�� 	,(�*�-���#��]����ͪ���r��X�b�a��,��E;Y�aF ߞ�*!���p����P����ns�Ե���3�X*ul�d�o>���<���'_����_yS(~:'�B���M�Og�{��_��/�ѽy5�Ą�(r�ɸ9a]G)QMܬ�1����ΧLE"ωX��PՁ��) N�Zh��v��)�j��$:eKb�����b�o�g,���NZ�P�T�����:�;l��|���:�z�3Ï�<�z�n���X�/O� '�`@�UeD=J�@J y��{!pC`�A�g߃������b�J��F�V���}-����`XäC8CS��l��v�^Ms��5k�b = R�'�4ְ��/�>�X�w�E��P2u�9��0|<���K�r����6����i�4s"���x5̧�]�ؐ.��>�$�L�*mb�s����;U���b4ȃ��w_r�;!�n���m7�#�]-U�eQ��2���>�un��Cw�vw�I_w<Tb��Y���
�c�18����l�q"{�k=0i ��Y��-��2,���p�U���Il�tE7���Ar+��Hg&�`�Ti�`�=�n8�nr�����Z42�Y;�2�Xq�]�u����S	���gUN�����)�t�ǀ��ա7Wl��D-�'�z�=������:'z	R�p��RɧX�E��C�5(֖�í�l���R��&
��c�że8�����W�\�x�|��O��ϖܹ���N��T�r���J�r�Qd�۬��<�iĴ��.�5�m�����c�pȮx*���~d܉~\�~�F�'ۘ$�,�mVS��z ��4��S}'ؗ[�b��8�w��Lvp�s����u��797���]��S���ZW
�X3�&�H���㺕�U9 vۂ�/+x�l�λX1j7קc���K -���F���<���^�@�S��a� �< ����֔��ϒ�vs�޼3Q���3wKߍ�=�q����z��
�+��K6NP�zK*󉾆kY�I(nB��j49d9�f�c�w��f|� Q�hJ{#s�V�2���J����Yw0�|���doZ�7`R�#Φ�\4���D_'�79M�w�o�nu���e�!Y(j�K�s��S~v��O�Sd%
���uK�u�l��'0�`Ի9N���Ͻ}:�t��T����<4��� �$�R$GL-eg�=����NϹ,�>t�dn�ԙ�+a�Y�(_�8�``l�g\��@6����h�V (�ѭv�Ws�Z�txԞ�2�랭��z0N���e&W�|fpl{"6:7���5�T���Α~� ��.@��ɓ>I`a��GU]_'�.c�	'��!g�W��7�� ������)���y�O��>�?�����:�u��ηR��,���o���}�E��	ͳn5�y���ؠ07M�^RO�c�]�Z����v��d*���i��[s�����(C�H�r[�óJ�t��B]��<)��7�R���ߍvAMBw2FjK)%ql���+5b���LԚ�h̲��u`��r�WW|�<�M�+��r�yѼ��c�AS��M滉X�l1`�q�\p���&d��m����ϟ������y�y��_��0�샆a�D=w�߿w�߿�=�����pqoy��nLz٠WG�3b�j����8�4M�٭��&�'��{�;c1C��q�Fe�)ʟ�
i���Q���9kx����q�x=��-By�4ޱ���J�[��(f1tx�<��h��8�&�T�8����6�y�u:'���a�n���ɩ]�=2�K�ݘ�ޛv:����������ϡ�Z%���Km8f�nf31u˲�b��������֪�6��7��l��)�;A��x���X��/PM�lخz�WM)}ˊ+��2�g�&}v�{Z���)���^Ot�f���oU����o�^��'Ա��n۟�4>]��n��y�J��7��@��(����J��J?w�C�<��~�N^d�b���~A��7��z��?O��&9| �:=�  ^��^��� ><jj�W7g��G���P�Wf����^��
�W�adC�&-���n;�0�kYF�]�3�[�*R�&l�/M�s��ﰻcV�t<�*4��N�
xv��ǜbFІtrD8G5������+�y������֞�����s�V�Ўұ��C%.eY����F�a����T��Aw�!�w��б�N����|a:�Sc7z�^��b.��\8F.�w��Dg=J�
�YW
Zw,����n�0��;���W��|ۼ��� O���p�FXx��x1���R�ܮYA��X|?Qc���
��<)j$V僥4��'���t�Ʈ��a��e+��}�,Ϝ%{/gSƤ�}�\���Bc�X���� �w���;���W�R��	��\#z��0z<�4��R.��Z�z��g��0�4�־blx3�1�T�'C<5<�r�ƨ��~"5�x<m�ن���}��jGti{g����b��V>�SP�>�@��A���%��l�	s̈́G�0n=J,�;�60��m�LL*Qޞ�b����x�{���~m�Z��� ��G�( EE�	�~Md�N�����i��X����S.��5ݣfzAVer:$oE�w���f��g7 ���q Gz�ޞ���ά�Ǖ����`D��h�,�7�]�A�� \-�v�aȬ���3��,�`>��K&I�t�u�09�nAC�OC�Ϣ�:����B*���O��D�X���<�BP���uCc�W��t�]��������g��Ě�q���%4�Py��bJ��>ğ��%�T��a���=;;4�~��6�sc�ذ�� �g:��U7�u�LɏJ�靁nrK��U�#�s.䛼gPtdPJ=��!t�_`�[���8��'^6�Ҙ�|0]�ML�׼tQ篃n�w#7q�����:c��)�+ڦK"���66���Wi�bcL�#)4z�T%˗&u��ҒWS�W>�O������g/���%�u?�U��ħ��P�2���Up壮�+1����X�`O) ;���V�$[5;�^MU}Z(p�� h^�t����hw�m7m�wc��O�'<�A#hg�%D�|9�� Y���B�ݶ�%<ú���9�9o\��,��oD���u{s��@��u�V<��Lڔ��aĒ���j�r]��kT�N�qf�Gc[Yp�{)ݱ�9_}�g:��$���e��M�>������WI(X'�-A396D�z掩R��;�E��p�>k)���o+Օq��傸���]%
�}�u*4��9B�Hp0ul��0�\�A�Gd�����y�)P���]跴���������qӺ�ݻN���5VVJ
�l5;6;��������W�͖���[z�����gK65`87�t*�Z���o��:)o��p�ݷŪ����ݤ��X�t�������Hm���L��X�
�8jM�j]�����:=i�'-S���G�EQT'%G�
���[G�LQ�H�)��TKl h��I$��&������V�<f��ܺ�ghw]���[�e,��&Vb���HƦ��ͼ�F�8�k�)�;Z�Z�J�c-��,EI�t�C���|�R�6�J���2��E
��;�t����j�g����R�:��)�
:.ε�Y��#+��sgvm�I�8�e����z1���^���T�B=Z�4�}��|c`m�����l{G�.[U��������M�2�$E�0�4����NXFY"�l@���0�&��j� ���MڸAۨ��2wmetq�����oإ���g\+s�����湝��+�i�"�k,�E�է
�wf�9`�^�fΝ��v�"���:
NR��7[�����X#f;X#��.;*3Y��d�F=����"�v�y|S<_:��&�"�)�ۉѕif_c@E+/h�ᒅ��^�d�:F4o.��=�������2���j�͇��,�mr�ru�.Ҋ�ĂQ�H�nV���V�6�K,wU���Ѽ�̩��V5]Fظ�)�Mr�[�Lw&�SC5��ت����uc�۔{a!�y2)ٯ>��ӝ��Vo[��Z�8oU⭋�N���\b���wR�N�r��8bwy��x��1�9\�ѽ���[�/�PW�p�P������� 3/����,!�3y��)čIsj�����>�Pf]+��h��*h��Q@�(�D �)5!	��	F�T���$0��H0 ��b�Xh����v1�I�IN��P�i-Sh��d�I{����)kZ��h4_�����F�[[��{*+A�Gl�<�����_O����}�߃����?���Q�S�d���:*���wV��Ǩ�5�jh��>>>>�������>�o���~�?_�[���Ɋ������z
M��j���I�{~�Ϗ������}?�����?_�����O����=�`�X�Du�Km�����]�h|[]bXص[Vm�:
�R�
6&�ѱ��{ۨͱ��j��u�ѭ|��F6Z�5[]v���&�u��)���e��J[�q�Ê�^g�����F�VԞ�vh�t�l�Ϊ�U�E~��U�P��(��M4��uX�׾�$�Z+N���t�n�WE���v�j��Q��SC�i��c�GPKGj5�l=^G�;�P[
"J����F�I��Pi��G�����Zn� [�^���7��ujS|pC���@7��>9�5+�L���b7�����e���jd���K�k�h�a�?r��� 6[�<��~�?�
�$0���%�FF��A2�	:��!��&��-&�ƚ	���`�!�����J�s�j�z��kX�͖��x{;oe��,�HK��Hnˬ���z�[0G1�)��Z�ǇI�ZC3�"%��r#!�찵�2�dlE;-3i)��oNI�=�ӆ�`e�����E{E"���V䆛W�*@��x��Iߝ��.�	�� ����j6y�i���z�.�����c\�V�u�T���<j"�bNң0��t�ZJ��Q��l5�vcJOs��]���6G�3���0�ƫ�ui�*m��w�vb�N�[]j��l;��*�`R��Z�2}	8ucۧo
�@���f���'{��z�����:��o_�/q��?�i�DY�������{Y߮<�/�0�e��r�f�JՆ�mH,!�A­�1CX5��0�|�)�����Vqw�uW����1�Å��P��+�I�k��Dh8h�~�?;�;��2Y�ֆ g��]�w?؀N$@׏_=[I���9��H{�g�z۾Z'&�8aҙ:��}s��#��";��oH�!����.�������33B�U;oV���� ��N���M-I8��z��ځ��,M�!��d_uz����*X��SۨV�ole�������RC���M$C��P�xj�2Q�ֺͰ-�q�X\O8�����`�����֎ɂ�'�q��{s9��*1eV,KZb%��
���ˌ��NG�Mx��������q��ݬ$X�*��z���]��g7 �k9��O=������2붟S���W�T�de��<�����ae*gu�,i���m,$�|
�/U��i�����E�w_�ƾ��<\��(�n,ilÑO�ۍAWJ�;�kkXڗw^M,Ԛ]��᳠L�@�R!�s@�p�:��v�2+�
6�îǇ�QZ���%Nj�5.��併�U��g1�`W:b�˷�v�}�ͳ�j�.;�1#krc;u�VS�Ӓ˓ζU�@��Js튷c4�V�G���FL�(,�M���י��SK��p�#� ��E(��C�#�[`��BԊ��)�0��qp����H4D�(�<Y��W+��v�쒌�$�qv�R	��g��5s�s�k�IP�"��d��cqÏm�Ʋ��O.����ZGCv����Q�݆1Z�G�f�_�?�נ��ry_\���3;w�y2I��ױ�[.�{�ϓ��8��QH�~����т��gZ�6&�5�յ�A.��T�j�W�[9s���ԩ)W���F�BoΆG
�Y�0b[l��.�τF�~��ӅԫD�ӂT�]��R��.�.����e��/�֋�W(_����;E��jbm��f��o9E];,ӥq��1�����w�m�nk���M
L�9�-k�o��{�x_�C�0!�
��|X�?>�����>��������k��0�����hL���T�"�1L��`�<�x�#��Q�Vze���^Kc�#�4�s���x���߾wy�^�}��oa�>|����gUnOb�8�SC&pl��s�3x�wl�3װ��<´�~y-����16sW���@`� ��6�5`7��'��ov!{>`6uȜ��n��+����GE}m$��eo�Ǩw���!h�g���BUߨ��K�K�c����"Ǥ'�#w��P;���D�t�
�<�%�eP䳚%��5g"��u3,,$�̀��x(�Uc�q�/��,+�����|��p}%�U�#����4��ټ�"�a���rW/��u_�?NC���/~1�f�J�n�_��V|=��Lc99�5v��tGP�V��7/��n��7��nL;��P+|�s�&���
�hS���Ռc�]l��'R[Q�P�䮬�U�g��]���0ÞX��`�oPnx3�a��A��v�(����9F<q���[u4&��/�H�l*��ӕ⻲Yَ��ߖQ���GCv�̫z���[��/�e��:��os+H"Y�T����g�t
����;�:8u�����׾>{��q����"���s8^ԫuWWcݾ�׉s2�����S�.ݢt��,��W
��,�I6��]ˎng:�����W¾�� � ��	�
A?}����Ͼ}�ԵIo�y��k+���M�a�'f!&��Q��^�V/Z��@�U��ۅsE��==��p��8�*,��&ٷsx"��4�Djj�y+[lr�n���Hd�*���@�K$�g��5�1�?8oqh�_ɉ�hAZ�)�zހ����ڇ�so4�/�S)4��WuU��2��8��(V��Siso���FІ~90� @�i��h�.�>˦iEw=�8�hշ��fa�v0\�J"�tq���~�"=iX��I�F�
�GX#O�<~��o�tVk��;��H^t�dN�\�k�4��u��n#fЩ�Z�����A�oX/��b�l���ܮ��H��YƷ�'ƭr���͑�o\���H��� ���Pް}G�v�gČ�m��w��4to�X�F�}Q%&�!� ,�K~5{��0}��ô��;f,�����R˭&cJ�8���;o@�Ǿ���#�b�X�?����*��N*o�}pa�'5n>�]RB=�\%sFF<�v�c=�<b���?�<(�̟��c�i`���O���MI+jS�NMn�]�P�'*�����/�0�YZ�Rl��eΙY�'Z	d�x���Ό�ԫ/}�g�����8_r�Q}��9d�v(ի�! �o��IR�E�w�������yf+���w{��Mm�#��Ʒ��N�͘��W@�M��$H��C���`�"!�z��������UU�w�ܕ:�~d����A'�Sa�$�i�v�%�ɧ����O}o�{,��`���P�/z��l�1m���o:�o�-�N��S��d��v=�r"���c��o{8�ܮwm:�Ya�c���f�vǜM�����J�V5�́#�/:��EmmV�s^�ٛ���i9���Pvfp�?�׹�L��Py�
炮��>�J�+�����O#z���ũ���9	ݻ����F c!d�pz�����k��¦��=���F�֨�([WYJ�����cV�E��z{q5o��(3S�;�VW����V��`�Qū.�E�v�ژQ̈́$�8�oD�r|:�ʐ#���p��aF`�Z����dw)�<����N�*_cFFq4xD��b��O���Cs�k<�Nh	B��B�.;\N�/�>�ɰ�V>Ԝ��o�m>l�m���H�"�F[�3�ޑ]:D����Q�����<�-�5=ͬ͌/_�b��jt�1��� xS�����V[�g� wG@�bEt1+#L��'N�Qηna��ǅ��{\���S��δ��?B�޿d� ��ϓ�]��S�Ps���ў�oh)�uh��]�pv,N����Ai���9�:Yc���D�
����-�E�wHb��
XS��D2���zj�ڎX�ɾI	f�����Yǅ_t������{��
��U��C�BxUK�I΃�n���Ả	��<�tZ{@���$ݥ�1�ڟ���L���ز��B���r��hp��U�w��~�~1�<�a���z��}���-�{	S���?�N{@�ϡt��K =Lt��b6��hr�౰��ck�`����Z�Z�gE�����s۠��x��^��.i�� tE�ʨ��t��~��W�/ָnkc
g�c�9F(�t�1��'%D�Ϭf��Kk�/]���Ȯa<�������Ag��\�`��S�{I�w+�%�����yP��N����o�3�rw��F����[�@��:�i�� ��o�΢$���ߊ����PǞ�kH�LK���������扥�i� �a��Z�^��֝0�����W��U��c�>��x*�j��W3��.\$�M]�����`Z�V��Vl�]s'(od��QN�c���>v�C��g�>N��5�26���C��T���Z���CS��ݍ˼�ؠQɵ���د.'��?r�����;���
?���k��/j6�K0�u�WM�P��=�H~U�J<9��a�&��ŞrVph� 7�o��+c#.�,����(v�U�.��]}Q�UlN���;��q�Q�kV�ǘ�lZ�_��"�Z�i�v�κͽ���1g�ϟ����{>z���?�!�R��Cx�>��fnN��������k��ұ���Q���M��u\=˞��Aj#��+eF��X��j{��Z�	z��%�-(�>�q�z��6{�#L*n�:�9��k���t�5�tA��4?k��r��"�a�nZ������kӮ�;��!�����v�����N��;
fy۝�m�o�?kH��npxy�'bq�ZkjE��P�ܤP]��Q��p�uV
�5b����n~+��
�I�G$�ߞ���]i����>��ⳡ�e���eJ��]�{w�M��Z��:hW���t�"�ͷ�m���(�C����o�+����=5*�X�C�-�O�㉹��"��Ǖ[^x;�y@||H��̐�}&�R�g/�Ok���O� 6�t�d�+�p5���n�;�O���W0��z��K#f�e��dvܮ�<�2�)��i��T
rk����}sK_4C���[��y��Ż�V��񗹡���^kPQ�XE<<{��� H�Yk���u�����9No�����j�5:���H���K��q���Y}d9]�!qG-j�S��-�*30���)|o��9�SE$���!�X0
Eɽ���3}�6�-�ǭ��9Q��]v�h:ޠ˚̵��@��ݱE���f�2坫�B�3d�_Ϫ��_{�x��G�����n�I>\�D�L�i��qu\��?�z_�������|�W��),���E��xY�=ߗ�}4��?j��	?�j�ֽ;5��q�͍��GiT/�"\9�ieC�D:aQ.m�թ��vVFi�,wbyRo��[���i�tr|�H���p�2T3�k�a�Ij4��k���E'�.�����Y��}M�=��h�2=���)�-0��J.�«֮\�o5r�RX�7z���˹���d������N�sO���@�DG&��Q�V��ƕwr�5Q%<�i�Qy�I�0����{,x�ۃ��ڹ�/6���!�4��e����x�����0��^��W�clC�[���V ��2z��9+���y��^
̈e���B57+6�w��vi�����R�_>��%l%B��4խf�/�#U�x��_�L��Eߓ�����3	�q���mU���jt�:8��Dp�]����+ǉT��`��릖��ms��#{gt�-����=�im
�}�:ݓG��1�֨�"И�;�ŷ��ř��3b�Y�����z����MJ�Y"�ޜy����4�Z�5����b��0�+�mIP�XT���baHG\Ɂ��K�\(>�� ���ک�ͶnP�O�iJ[]��w��қ%m4��;����΃��� !˹� &s�))R�P*IB}�������  =���Le�:ym��L��|���y��>��I�@{�>�_r�t7�Z߭�����a����QX�.�ӐJ���m�i�0* ݯV��<1��ǳ��{��=�����qE�8N;�7�#�Wtg6�i�U�n;(U���=S�H�;"�,�1���u����اWF�.��jUc;�������ю�3�ʹ���N,��aS��z���� ��R_b��9S����5y4�i/|����-��+(���B&|}��L������q"�%6A�x,�6����ϫ��+��uf_9�oU-t�{z����H�*�����a~<�:���g�Q7߮��05�3���w��S��zTCe�k�w�
���8̴t��VpxF ~��G;�SZ�h���1:0/PT#�.�<�����^� �2���?��udVti�s�V�;c��^�m��q�w�9�=�h��K.]ډ/�l�✙4`;bj��U���~";��WB*�v03�f�Ov����ʧH�rz�
�Л�gL
��Y> 9 q�υ���0�b�EO"0���>�e�����<e�\)�;s�J��3l<��>v�l=�������V\O��l��)�eێ��u�_p��{�t�m��Vuh����:��E�$�{aΥ�4Z���o�����T�h=n���&��η�+��|}��<� xz�RZ���]��	�9���jQ��qSɻ�Fḉ1E��r��0C��4���bF�N7wC�!G���k
�oF�Ss�l<�NjP���'{���i>19�����-��i�B�l(G3�g�s�5ӧ׫!�_yFsm=h7@�iɄ�G_���Rt]ư���z���O��[B��wtsh	���O��A��� i{`�L�a�c�t�c9�.�ګP��m���SË��Pڀ�0��9�o3��E˛<�$�d@����u�f�=�&j�=�����W`o
��|��_�᱙���S�N��o�m�4 ��l�n���{6b]�MZ����"L�30sP�(��ȥq�_}T(w6	�>�#
$�ď��4ms�������m�8�Y<�����S�G� ��N6�wc����#��P0F31��rm�u���;�o�����tE>7�T0���[��#ۻ�#4s�8Г�0�y�M:�ͅRK׼��C9�\b���	���/z�pFT�xz<��ѭD�{�%r�ruA!�*h�>�oطo����қҘt�}%��7�3���,��nư�����gQ�J��;ۮ�ˬ䷺h�gN��:�@���د�f`O���'av���7�v��k(N����C�<{��X�379��J���rgs
2پ`�ϮV�b���Nz���9�ˮ8i��klv�+S��u�����6)�\�-:Ñ��=�RO�=��5'l�b����h��m���
rs��n�-���)�m"�ˮ��&�r��Žgbw��YHr���:w=��HS�4��E�%[V��(�F��26�p|�n�eV=�;�m�X-���QP���rcb̙ÝI�Vf��i�u`[��rsBlض�.�v,�*f�Ƹs[Q��fWh��H�R��L{����6�l{���&n�R�P�,s1��(Vق.��s�æ]��m`T��\kl��b��ooqr�F�QEK,�E�g�0.kU����۾{���Q��OptaU���r��M� ��q�#/��$݊
� ;��lz�1�,u�;���pg)�*�6��g.���aq�ZG)���*Y��sZ���M�⭮�	e�gb$Q��7��|y�(�b���I[W���O ����ڏv��:]r�v4�ݛ��7t��\�k��U��;E#�*��t�vekt�4�{9��8��;V4X��REaX�1G|;A��Q���&��J���Bյn�Uy%�'�riu0�B��ۆ�݆�kB�+Rh��%1�炊RB��x!7p׼�+Ҍt\:�Н}�K�}�Kܟ�Q�Z��lH��N�g�v��gz��3���SFB��b�=���[\��JX�Z��&��Ӈ�)���:@n�u�S�}Cqv�������>�ʛWt�Mñ��uGi�;�.�И�K�t��X�Ы�0�F�	�4�pn*�ƍ�[�T��S�A������렺l���L/fSCTۭ�W���]��]�:�N5�y,�Ν/�ZTnR�9�7��R̈��7hH+k9�R��BnwQ��N�o�2ۜ��/z����zm�8Y: _A�{�R/gݷq����#�wY%_<ŵ��ux^�8}�[���e�w.��z�ݑ]me=0�
ܕ�h� �O;]{�mA.V:3N�T��h��=�ڦ�23\��ޥ�ڊ�ְ�u���'i��R�6����ȇ4p��R=eLx38.;1#�n(.�/r���[ ૔�}Χ�K��/~�jG7�J�3�w�j���kyf%Y�8��:8N��ڳ*9���ᢲ�>�}�K�i[�2��o�+��3|�E��49x�U2�j�Mv�m�#VٹRa��uj�xR�.�ǣ��k^��okz(�fr�ސ��˫qu���MQ��>�zu������oG�������מ��3Q�
6�Mm����X�"�ѵS��~0qWb�ƪ �cR~?�y����~��O����}������~}��'V�A|�'��t�k�:�[jӣN��fv���=;f�*�w+~�><��������>�o���fO�E��g��Ѣ$���:�h�gF�|��E;e�lU%5��U4:��\�x�g<��}�_O����}�ߣ������_2h"֍i�ښ��0F���4Z�itk�n��Dj-J(�v��EZ������Ƌj5q4��螴6�-�{�3Eb�El�5��흰h5E��i4��������S���PPPR��6��4[8��j�l�~���Wh�N��F�:=m�:��l[Ť֍�V��5�t�Sm��1F�����J�$�W����;th��q����&��!đ5�5c4��h�f��tX���S�Q�V�"�C[$l��_��l��VƃbΏ��h�ʌQ�Tƍ�1�U]�����Z����,^��tEIM�ѽ��;7w��]��<���͛�GÉ�{��������YGw��l=x���ϗ��W�)�2��C(�@=+V#�K>��$�~q��I�=?���#��1Zy�w�(�OA�������Q�B�ܵ�t����Y���Ȍקw��I�;���7(!��v�b�G�&T�CFI/�b��1�˫�ٹ�Z�D�s��y�C��9ڜM��A��k7T�!���[��Q�� ���w[x�|yT����Rǔ�nT4��������*�ݕA6�ɣ��K��L%�2�
��^��֖���+�ࡐ/雋"i;o��S:�MA�0�w�Dx�����j������e�c�z؞zV�	���!3���7H�K�[ �iN��3W=�ZSb��i�*둁��-�fN��ʱ���R{� 3~��O?cFv�~;��}�@*���}uCʇ�g<��E��V��}�M:�Hrܡ.1� J�pU ���s���C�{'����9���d"4gc�WDw���u�7a��J)˱�<���Yv�p�;X.��D�����@|���x���E�B�E�)�l�<�3cH��0�4��z=�T������w޽������5~~�_^���n��_xٳ�(��-��?9J��X76�j���k�	���ٷ������\lJ�y]3��{�V�o��U�����x�aqn�\�k�K��OV啤tf�/,�,PB^H\Uv��;@�7�y�V�4<��
�:�f��}_�`a��U;��������������o>oҢ�+���-�0��äYೠ>H�8a'���CB�@�b�<��3v��v�9��bb�p�m�NǲmH��K�\��~����E�<��1�m=��EBp�P#}�/����F��_�dz�)���2�SGe?�2�FQ׾i�g���M�b�J)�noE��)֔�佴�d��T�hg?:M�kMgʃ�\����`7�Y�Snׯ��:��b��.��vVl�=z��,�u�q�� ��8kd�=4�L�����ؚ��;Y�KD��<J\�i��5�p9��.�vh݊v:����98���êw�q#y���`Q���^\̂i!�:��dCh�trR�&mlYqeC;l3�Q�ힼ���eV=��gL����Y�J}�qL��fX�:=�C��6P��/�>\��JCy-����r�>�����Y�/45�E�Qc�g��xJ�4f�6D�ס&�(�ε+Ʊ���\�
֮���t��>�]⛮.E5�	0���E�(�Y^��쫷�Uz��A��[��G@>K�]k??D��t�ej�n'�����9y�*:6���x�o�$����v��A�޻�~�?r��Ϩ��v�ѥo=�"pT�����"�\��t\7k�Re��"]��\�7�<�v��m9�Cf[�Wg47��΅�w`]��8A�u��q�2�mɲ�.��6��n;��yy�^]�m���BG�� x4�K-U����>�9.�����X+��V�H����p�5yڋ��Ɛ!��6�tk��f��FT��2.�t�t�:�3���2�¥��v@J��pA�����_�ʦ���3�A��ڌ��c�;m*�Ilx@��0ޕBZ��ڠ�"-=3ᥛم�৳��Yp3�!:y��Ԃ�f�LU����;�^�_`T��.�(�"И�#X����l>�yǓ�')�!X��	v�I�!���\�q��"�)�n؟l\?c�y~�YSfXk�8%��D���6��g\2P:1hm\IE�Y����Fk�#Y��P1(]��1�uKM�?0�p�z���'@Y��2��_���c^N�C�z;)��{Jg�f��̥��5R��n+Yk%�t���9���K���W@�����D����sM�ͬ��q�,CMl���2�Si�S�q��8Bآ�-����lh�lSi^���W6��*�V*�=�.�t.]��	�������tK�02.VŻ�U.D��/��46��������p�5U�̭Z��gF�egjy�2<։���N�xΩF���Bμ��@����X���_7[fof��(]R�O�rN�y����:�z��b=�'cgbm�U����� �ƣ��+��Av�q,הFW*�)eq����,0�����������ߗ��x��0Ҏ�5,��<��W>�F��%�P0�t��kq�55Զ�������ɨs�G�~� M�,X����Di����>���'΢y�1v�<��eeI��2���29oK�S��0�@r��U缺wi�Ǒ�ɱ���u�W����+�z�䉭I�_N�^���j�w��)%2{���;J�����܁$
�eNH·����zf��-b􂑭��?���tD����N����"9C�x�i0�:���^��@�q���ڀ)�bE�n�QeU��3;���ο(/�4�R���Y�[y�[���<ߓ��r};!(V�j�/��km���Ōn`gOe�L��qn�̇�	�/BN��f-�4z��@�}��<��/�')������S�f}���W���y���R����H�)���0M�q}�LA��(ec���
BM^��O�v���Y+[�m��������?B�P&�s�K��2�|	L�����N�Ύ��z�����U��-���������P���ұ��4q5�Q�t_SP�t�4M)����d9�νc4�ݰ7sjep�	�o6�롧 �'��W��x.��w��Z�g=�;��;�-��w	�u�+�V�i�0���YY �3��[�x����!�i�ӄ�$C^�nU����8�S��ʥ3�V=[o��ڭ���W�����#����ԫ� ��_y���=R�n=�O�w6	�*�>�Qi
Dc�E�wƄ6�p�V���n�1qC�7~>a��[��Qؿ�dqF������\VtT�J�!O�Ԉ��4��B�mj?�Ka�"�5�DK�.Y��%����lM��>�du��:�H��4 %<��<æ�+�z^�b�h��_��n)�̂��Є��xz:�[�=�2���N?@�����H�Ux�����HSѢOS��z���o���zY�P5k���:�
�U�������k�>�/�x�<m�%�i���g޸r;��]ކ��W34��(��D���
�X�W�0��F��8=ym2�P��^�r�%QR����+_��(_�����6.�j��f���@ු��=��^J��t+�'���<���I�J.��(�an�l��.�8Y�?q�߇b+���*�(.6�Q��F�)U�Óדg^)�Jl�2;�.�)ɰ�]�2ҍ�@���n!�sǈ�s��4�K�ǁ/iF�;�\�9�5�y)O��l���x<���Z\K�S�@�jL��32�Zq�ϸ�^�6�r��T��G���(q��Y����~~���~v:j�>w��מ�h�Zp
a�Vyr���?v��;�Ǽ.�;�ݔ	�e�IO c�Xr�Շkr�u.���"7�B~����_<}�#�
�\Clh��}Rǆ��K����N���,���Ҍ	݆1Z�Fl��訬��ׁ$�|�j����Qq��F5;rtq�K��ƃC�:��E���X�u�"��t�qԘ9�|�D�3���y��7�df&.���_���r����Qh5mL�|�`��D��泗�\Ɖ�/�6HWf+Sn��9@.������ǟ9L�y�Ѧ=\��	��w�\z�j�u���cΕ}�zCAAa�<z�u���,cɅ���(Wib_<����ɡڹ�ñ���^ȭr��kZ7J��}f.�E{z���A/�U����h^S�s8��])T���"�)|����͛��ܪи�ML���ePҫ��_Sj����u/��x<�I}�ຳ������3��v,ֳ���E��y/�;�.�����"(�ڌ�sa�.����m�<�'{d�B�`�?o����I6�;��Nʄ��b���]ߓO���Q箾�Z���]�������b�λ!���q���x�G�;G��ia�_�������{sϏ��byB����&��t3�uY,�ʹD`	\�n��v�bq���]L��7�pf�=4٘�e�Ċ�H�LIBj���$�\�s��)K�fc����>�T+��Jr-4���J*��a���vT.r�=�/���
�K�r�h�V
T	 ���� ~C�<G��3T	k3�T���s�%ܐ��<�c����M SI[�5� zk�J`EZ��$ϖT3�l�c7p��x;���iO[҃�����g&�6�3�&@z����Y�^SmZ�>��/Z�𠞸��yq��#�����O��ϣ�CO��ǹ����2��(����؎M�(���[���&��EY�Ű[F��J��N�C�?��ل���=� "�E��k�i��N�̉;�>F�L]�wV�L��n��؇(��U�Rq���F��lf�R��� �+Z)������v&������F�oG�w�ۣ�(停�%��uL!��s���i�^��ή�O�4�)ۛjy�*�!2��I���q)��fשN�T���C�y6g[Y��Y33l8<�{e��wa?3j�
��y�������t�`�Z����R}�\���!��f��t�7�]�@L�)�0�#�IM����0�Uzb�w���Ⱥ���l!��q�wn�;�d��k�H9I=֙� �#����tDxK�1-cj�J0��mL6���
6�:Ъ���<��ۊ�
�ɓ5R
�7�3U)z��ܐZ�>�+��'s
u�YS�8j@X㱮'�W�>�
��c����;��t���'']�0�#z~_-�5��T�+�@��Pպ�U��N�5ձ�ۓo$}�s���G����<G���j{{C+R]A����ߑ�w@�;#\|��3�O�DǾg%5�t��e��"����⭛�-�YAL@ӕ�P0�s�>��.h�k�){�+�L'�����C���/H�|ʖ�{u�S�N2�)��T�^��y�����O$��ItN�h�d�!�}�q|�$�`^;g��#�|�N�x�b]��([�w!�[q�h����X[�TÐF��p�<Nd��l��s��L�h0e�����y lr�8�������6����¾`a��(ϫ}G�M�TM��������ྮ���J��8%^�c�=�Bca��A�ی�zJ�4D�ŮT�RJ,�~m{�n~�0k};��l?�W�0kG�.S�/�Y��j\�%�vy�\�i��r�t�\�i�M�+�"}���8���eO,��t��`��{ŕ.�1�Lݰ�Al��M����sJ`4����m����OtS��@-E�y�+y��Zpe������ɧ_�]�|�k��M���Ӱ�uן-���9�~��Zӏ%�X�U�n�?ڽ���R������W<0�s��D�Ub����n��Z9��Hv���:�Z������h��MH��Ҿ�q�7K�z��v8ㄍs�54un�U�R���Ǟ�x���^��x_����?>]����jfC>�:�<;�a�Bs��T{*UA��W@x��)����V�q�͛���u�*M�����F�0PMl��6ŷ'-����r�l;���"%���:�2|������.��t3����B��`fۆ-���^�K���1�������&�k][�β_9^�܋z\m'��S�3�����:�(`֕`_�E�/ߌ�xg��z�y7:ڜD6u?v��$�f[g�/*����M�o?�u׮���|+��OY}��V+�W�|�,��[���دB-ncn��@P/�db2�4�w��}�G�Jۏ����)A��H��ݼ�侼��f�P���l�'C�d�Iё3�S�睎WVHc��(q�7���K��d���Q�;��ML���������և��ҵc]c"���L�/zB�@�M:����≶���Z�suĊ(%M�-�קff��F4�`����/$b��щ�9��_E4�qƄ��c����.�r#�ӻ׵����8߃�-T�߀�m�Riw�×��z."�Ⱦ�1�%a��̓w�lPu��>zYq�ַ6�7�2a߹>�b�����SV�.��$�S+->j��)h�Or�����&ݒl�षHJ���ްq��V�o3X��֯���솰L��� �G���_��o;���!���￞�o��!��'�i�~Ms9F�.YTv��i��44��획@=P)�+�1.b)2坙+�$�X�lk:���EkR�M�1����5�	�ʷld�)��������u�v��]tF2���C��x�^>2�m���ԧ��G����XK\),{z[yj��'����4`.��S��6n�9*���$���f�{���6P�Kݑ�	ğNk�䞇4��ܻ�gY<�o1��$�,�~���:�yU��q�}C��(~w2/S��C9����Y}��)饖�r?�k�}|9<�+�]�{ba��0ʠl�gZ��dw���J����cu��MӜOB
���&��⌄�4�<��hQ�\��K>B�_��<zl3��@>��x�Ԝ��}u�ی��5��(��.kc	�e{5�s��:�!|��#��~ɬ_�mV:iC�>3�@�j��h!r|Ɣ�z< ����{dY����=3���~c��y�0/6�~
<ФD`��qN)�}O��-H���E���䴎��/<��&{��nC�V�X��7x�愂^5��f�d���K:�U���`�����v����9fL}}�bK_5Leh�M�5�h#���@�D��N�Ǻ�O��jt�$���g^wdR�=����2�\�z�
�*�Hc��ɽ/5��*��Lp�aa�L2�|jpW8�-h�e+�>�mꙐwX*��@�.�
w٧%s%�#��6�(wY���f�4������
X7�Ϝ�K��ڴ��ٸ)q�7�+��M̮,FLʐږ�ofڥu�N��Ʒ���[˶JX�N6�WʳU��;9��9�R������ʫ�}�V��,WZݎ�~����91�J�K�odi:��l������kv����Cn��0<��"H�5\j�|tmA��n�f�
Oz���u���K:J�7��0�z��\�l�s]���Z�p�C,屄t9�z>�/{)=}��ǲ�۫R,�;� ��9�i�Kz��@C��.�V���ɻ2*K~��V9:
�+U^��qalD���y�-�7+ ��80ڦ
I]L�s���ku�0yd�mNv��%�i�SwV˩|��l�
�"l����n�L>C�Zfjh���)y�r�v:�%�'0�
�9c'9���P���hh���l��mܮ�3����4hv��x�m[N��7w.�U��ko3�T�}���T��**X��mw�#̬�p8���=���X&�X�	D��XtR��bp�N�V�����Y�|�Z�`�u���:,
[v,��v�&lD(c�,T�Z���Ԓ�ѡ�)1?�E��]("���ε(�$����a�}Oq���j�p�Dr��`I���]:)YE��#}���p�un��z��W[\�0˩�͗̓ctV�K�ko
}SXs��N^�ǳGuڑ���WPv�%zTES�����pJ��1["��|Q��mf&"YKz�]��Q�Ş�tT������,���/��V�A8�_R���u��.��wN�LTL�֝vb���[G��/�͖xv�[���]Ys,]�3�R�w��5��h��dܲ��'F�^a�Ҙ��5]s�^�.���-��8�E�#z+jm�C�i��t>����0ndSi��Ӄ����M٣�ۚ��w��.�E�)�Y�gF�8�<۷]G*ŦqV��g*2�����\���2�aw{��fa�0s�m�5�mq�fB����@�.��pR�j�IJ��_b��/:|6���wr�A�gҌ��e����3oN�9Xov�;F��Y��s��/_e�VԼ.�4y�py\���*!�G�u�ϙ&�"�:���J'7)���qȫ7"��G^��<���KBX�)���y�St��ۖ �;�Q�ϧd:[�)+/-��t8�):�q�W]Q=
���ᣳ$��N����{Ik�y�Y,d�O����y���
	���P(�G	*B��?���uɯ����A�?�FW9I�`�C����f<�@��(�!Q��i�7 R�P�A�Q�P��H&h���Rgm�rxy症p�t��qlSN��E�[SM�тcZ~gE��ѱ�6�q��g�Ϗ����}>�O������g��~���N�j�
�M���T��:3��6#��tuZb�_�����}�>>>>�O���~�<�~��1���f�3fJkF�յ��ւ�Z	��KM���������������g��P|4X�5h��i�k���j�m:��V�<�v��6�[Z�]�� �"<�䘨����M�Vڋ�㝳��o{T�^o#�����-����詨���lU�E��1[Vj6�f��7v�&�-�EQ0N���w��⪭^���D�f4oSmEq��z��'V�;j�E�1߼d�'��STzَ�5���yZ��ڌUNڬTm��T��5�l�EDEkED�֨�DD�h�h�wV޼<|$�E���w�cDm���N*(���(�5��A�=U��UZ+-k�]	���v��۪61��zخ���ǁ��5�>w|��U:���֕t[���������!u��v��\9�ɾQӣ�=s�KZ��=�QQ�ɵ{�
�`$��ۧ���/?��n��)ަy���Z���f����g�q�2�i_ʈUQ��x�a�T������fs�0��_t���%�;"���|X/��
{e�h1��3�J������֋9�I��?�V;��)G���`Gb�����a9���?�`$�D��yfY���t�-sߓ���
�De���!�f��
���=�&I�Ǐ��d���|{��iF�4�N�:��������6!g]���kTza���5���N$Ct�	ע!2����T4�l#�@��#W;�E�(��v���D��+	YW��P-֩-�ހ��{��0�,2k�k��zM�k$e���u��	'Z���V�)}u��k˲\��b����%�Ӷ�q1*,��}�]B=y�cz�z���87�t�&�T*ۮ���&7���l���z��V�Ǉ��	��z��W�s4C/���|��A�H6���v��N�u�}�U�C*:*���f����.����P���s�;ޭ�i���6:f5Ք�Ӫ�(�/ǭ����s���L%c
�H�� ^=;C�у}�K�8~;���R�A2�^�/"�ը��X5n�"-�bN�n�RN*��Ј��M�`��.�r��{�)n���½�}�_S;�sxM�>�|�kSm�vI���x�F}R�����٭�H����Wo*�������o)d|=> {�#��RҵA��p�M6��O7�V��'z���G��S�#'�c5��c���3+�]�2J0�j}���1ɶ�����"db����R}�C�q�-6����n�n��k���]2�&�G�'������jg.T�F�U��H��uƵ�<v9Mz�^U��z��RS7^���S��9��J����U�2�� ������͸����W��ޟ���=��-�ƺ`PO���OCD>Vs�;G�{N�v�<Ç��uYSW��wr�wWG��0|c]m������s2[��h~�]����&v
!vX^��/N�P��TG��x�N��-��.�`oK(�+�ո�u���M6͵�~�����|I��*�^F��g���t�;_��9z/ک{�c��:��yBy3���i�m؈�j[7�4�YwB��N�n���y����UC��ԮV�(aY�����O��c��5��M���
0�d�t��W�sy}KF�b+�tj��gD�y����WӪ2�C�����7�8�.�e������ zd��˗�3������9�FV�0p�7����F����y�(���Ծ+�U�V��M�ͷɍ�3�����W���M-����-��2��MR��6(9:�%qB>7�{f��shg̍m@-~W#�%4��o/]�)��*3��D�Agh��{5o+���e5B���'qz�=��jK֚Vm.U�+�͝k��hR�Ԧh�[M�&�e�=�2ࡷ��[��Kb��qᮥ`�	*�U����ݭ�.v��<� �f�`�ro�'�6�pʖN!b�_?��~���Ӊ�I0���̷5.n';ʷ��. =}�78<;�,X.�j��w�M0K��͗07>EU^�I�+/K����&�G4�±�oC�%0}�^�Ӷ1jƤ��7#��<�̨r��&����K��6ۜ�珒�W]54Y����k�o���u�v�w-ʳrw��Z�����o���e���6մ5�\Ԁ|��H�����V��j@9{��O�x�֐�N���,Ӓ���L"P훇0��X8�	.!2���T�';��Q�]�U%f���@x;��
ʓ��^��1e������C�o/=����r��2�|��[ڀ8����%�W9�~U/+WQױo%Q�����o;�ndAg65�����r�y��I`�;�P��!�v��VA���J�:��G�n��B�b�>dB�ƙ���憨��6)���2od���5�����v.<�D��j�F��pn�5`6+��U��真+�Q8���g���z|�����+5�8X9������G]2^Z*��E���.B��.>�L��\�>#v�G�viY����nȪ�@���/������R�z��.ԳR�F�%�1��q�r�1F������E�r��ku�r̞��]ʲ����M����걛���o���j%7���]�y���Vܘ,�����v��̶[6��Kw�חU�>6c]�$O��,y�Ӂ�%qm������Ux�ua阸k��ݎ6v�_e>�����,�H�b)�������;u��2���ѻ�u%�ۙ��7c;\Tx�{ ��oҮ�..q�����x���b$׊������v��zAKŇ3�<͆�q�|��#�m]�ܽ���r�V�Ѻv�9X�5F���:J�;�!J�Y܇NV^U�>�@��ɬd�X��&��4��Z	�ʷ�Ǖ���p��r���s�{٬P@Q�� �@"@*��A�@+���Ӌ���o��1����	\�vR��Πu8Vf}s���U��z��m��x�;9�h^�P��c�mDY�5�T7SƑ��+�\��y��	w�{��2��Bw�;��B�����o��H�6�]{��=��v��<�v����Oo�?��m�w�0U�kpZ��U{�������'3�-����b����F�N�ؤ��Z`	Fx�ߩT��S=�{q�(���jʪ�����+��t�k)u#\��ƹ�:����j�[�]�i�>]dݨ��.���=߷P�5��	S�J�*1P�-ucQd'������5UUk
��I ؐ��.B�b��,���m,&ǻ���h}��S���T˯ҿ�3=����2�;�A���G*q�1�;-�w袲�f�8�^��6�M��MVZ��7D�r}��)�M���X�@|\��_ 7<ox��y�7I;��T͘uf9u�y����{]ܶ���ٚ>��=���O!���5!70����+��}GD��r����ut���[W��sI\�W4n�K�s
���jI�,Gn%�K��������;u������o��b��ׯ�������y���u3WL����x� �ɣ�U.
ה���-z.f�y��7ݝϷt�2�r�֢���~����gƯU��ׂ�2L��8���]�tf�b���\��>��9C�l]x����Ew����i�������8�H�L5z�f�9�vqX�����T�k2�>]ֳ���0���5�\�&���[�NWy�i���.�=�͕X��Z�v�m��w�R�	�Uֵ�)���:t�P�P��ͷ��k>J�Y�WJ;�)E��s�ʄn+h�M5�'O��>ЬMa�"���(���ur���Juy'���*�μ�=�C����j��`/�u�c�惊!��بI�!��j��Md]Vf�&�Y�lj֨ݬ/͔��0�'l�3j��M�D�~}�K�Z�Q3�U�[�b�WG4q������N�#���U�0~3-'`�_��G"�p4;q��y}�M=
�߻J^v�o�+��wV�5ɠ�	k��R:9�Vʵ��x�ü��zG��H���	�f��kp��M�2Pn����ڹ��5�8��e�׋�W_������-�d�u�z�jޑ���5�;�~;�4Hp���ޖV��%���Y��;�-f�'nV�G]���>k��}H^�+v伱�Fy��71O.�OBjk��f�s�=3��t���Z�EhL��.���6fd�`~�eP����޶�E�3>����puK��B�y�ԥ���=J{�1��&��Ft��Ou,����H5�eh#>޵<����ˊ(r��Y�����yƷ-�J�([>�z�O�S[Q�,��o9OS�}|s���,ν��`/�"����}5�Ρپ����x���&���]�7���|�sG�:���͜��Ѯ�`�N�f��cMU؜�c9�3�N�4�d>���6(^;¿xAw�eΎȘT�<uz>^�n;�d�l>��p�6l;�חƔ��֨ߺ����D�����8�'�Fe3*P�m�$�������т��A!b��țZ){�0$,P�Lv]���M|o���,�^y��t�s��᳔05�o�c]�)�Ǐ6�S4r�.���_k�%i�;(�b\�B��GɻUs7U����>�W%ظ:�g��{��˻�����س�?��!��kwEy�����̕I:�U%J{�i���ۑ��',�҇��\o����*-·�z?}ޅX�7�̹ȠE� �6O��=v�F;Z��#U�n�]c��m�`�7�I��׈2������A�Q�, ��_>�a��T�x!�q۶q��}v���l�j��؛���z���9��%S6���b�X�z������ݔ���(��֪���ú��0w��+�`3�fG���:��~��%�0�Cb����d��fn9#{8O��M�m�)1?��J�������
�s4���Y|q�C��v�X9�y���T���=j����G'�u�f7�gFgms�j�Q�����5!�^�UJ�e+�
�#��!�0Ǉ;)��ȵu/�K���zֽ,�����d���W)�	]��s92M�^'�s��}Q�r�s��ss�压 �Z(A4�()Y�n��Y�Y���ۻ!9̬�'�pA3��'�^]��=���^��=��<RV�0�_8��Ô����on\hc.��dz\����^��(�~�y�m�\xZ���0�{<��>z��9V�L�4h÷��~�͚)T�O�*ּk�r[�O�����|�3���绩t����vd
��P�� 9�0:�\�l����-q�=��;�9xڕ�}��&��h4	��+l��=:��'r�r��0!�g����8���29u�n�p�^òّQ��!ˑ������p����A���f,�Ԭ�����y�SVƽél�<ݴ�3����M��mb��?�[��Ef����������N����ƃ^͕�l�K['�dS�sݥS��ꞽ������u<=�����y�ݴ�0��r�8��)؝]���ѻ)�r$�t�L���j��L^�*n�G��Ό�a�[C�m�D��#�-��Z�2sc�E���ef!�]�BmP���,ij�ug��c�����}��'� V(P��S9�]p�_�U.����t�@jžY�1��W0��nu�����[\X����w���w�N�
�;�3�0��!a�ħd�R�s��,3ժ���WR/�ڻ���U��ƺoW�|<A�[g��tB�v��G���Yַ��W���t�q`g͋Hv�'��ڽ���f;�n�Vd �*���a�щ����i���F�i�(C���z���3��-���/G��]��13��лО�#��W,����E���33K9ey�,�/
$ˀf\���lJ�`N����vn�5dzT���1�v�/u٘p�ޞ�%8�8���lӆ��v�ذc�f�3R������n�7�=�,��ۘ���&�en�V@`%f$Ke5Ol��b�
�{�\�`T(�}��~[�q��v�̡ܶ<��$?KT{d;�.�.�H��=4�;oۦ\Z}�jWԻ�7�7��W�Ľ�#R��Zԙ��l��R:;A��4�v�:�پ�+�Uvt�,R���ڈ"�se(��K�Td���,�Õz�	�ܥ��b����u�5�z�%����H����^U���PO��5�,7�FT�P5(��Zm�r3�-��,�����1v�c5��]��RX����=��vz	���:�mtkX�2���f��\�i[�7���雰U��e��u�vI��}�ra�*��E˥x2�@�y��E��ಝ�]s�_ݪ���s�]J���x����`K���ɗ}��֓�+������Etĥ5I:pr��(��NPʔtfē���9�d*tk-p�*����3v(��x���y8�����'Ee��5��2
}1��m-��+�_-p�XFL�EW/����t���`�����b�Ѧ�m���kqd�T���%�s�Z�B�� ���;M����K-hֳ+�y�1TI���wr�;xл"�Ȳ]�;���1r)a��Z�w u)i��H�B��KY�vy.��_Z�4I��Z���[|��'Y�\�������^�J��H��YB�O2�
\D�e^�o����2����K���E�aݬPWM�Y��z���.��p��ç)�	L|��#5���w�O�q���V�%�<��x�#u���|:v��w�8n2�c[��e�F:,
��{��}a�٪>�����y�iJ�r�s�6�V��&������m��%7�e�����yl�s�HvZ{��m�#B��뢪|���+���{IQ�Sc�U�HP�Z#�@�'f�M:�5,��b�Th�����R���b�
0�����}ϻ��̗��%sBA�mY��c��-}V��\�����z�! (B))S|�����լ�ˊh;=mvT\ga��-�������Ժl7��i����-�9��H�{�lf�FtZ�.�f�t�LE�����<�w�Iu��D(w!�l@.I��y��k��z��>8U�g���a�u�]\x���p��9�|�1�E�]��V����q�=-k]���%�,et��&�����^iV)mC%�݅}o��:���~ds�e�t�_0嵽�t(H$���{�l�NN���恗o�N�������m#1r�p�ź.�R}Xz:�S��m 6�[z��!�U���T�&�I%̏(�;���l�O[��XΓw���oeH�Yiݓ���Ac.������r�E�{'W:�*����Y+$�-d�[/�Qk���ݻ�S�7R�yp����T�뫎����$צ[�ե����U�Xo-e,�;��bL	zM��Ǌ�o(
ʾ�Y���J����Ʋ�W'O(���L3o]j��60�����#_ ���`��Dv�;�j)�q�WSJ�i2����+U�BS�W��z�+y �Kk�J��7&�{t�c��m��}\.�e]��>f{�<f�>3�N̄�yg&��z��U��=潼�k.������  A��k�5��kmՠ�W�w&���$芫F�<բ�������������������������Ql8�����*4(�U�0����LM5��;��wu����*6�5]�q^��������|||||}�����f?j~h+��cDUAE��y������ڨ+kn��1h�ε��Y�FH�������������������[��qd�n�l�6�ǐf*�&���j�*�ѩ�Ƶ���h�b�<�D]��M�1�V#PTD�X��kT�T���z�h�Y��X��)��ǻ��
(*��~]űj��V�U�X�6��b�o��Ϊ��H��L N��[Xō�b��9��&�;Z�lO�b��v�T�TSDO�s�0[b�*�j����3�}puz]�<��
�6Ɗ����MGl[$h����=�Yј�%5U���U�f$�&.�*��"#�um�v��A1�*�3�i�TPN�*'X* ��m�譬V��mb63X'muB����,�%�SOH�ʺޞ &����.��J�����z��YZ��iqW�I7�G����k�b�W�С� �����5/�_���>W�^;_�L��c~�U"��}�jٔ�xɶ^'7�6�>��ʨ��{5�c�_�҇Zy�0�-DJ�1h��>�����f����~^����cQ�1�]�QwƲ����,��u�j�f*�j鮯k�v��h�Ƹ�MZ�c�����S�c��Q�((�)��N2֚��/��z��w��г��Esl�̪���v�c!�O}�%A⺥����ro;��$;Z1e-����q�F�v6TW��S��d���율�=�=���W���@�wd�{
5��.&��sۼ���Kh
�/��V��2���t5S��O�UuhzJ+(���ڹ�z:y���@d�G�sjY�B�$U��8#:��g{�ѹ}�M=��'�f��t�yB��S'˼�5[��NK�����}_�b�/�A���!KUv�2��8����ݻ��\:f��Z�_���[\�9�r���{�������A#�uؿ�d�8SRbݭڈ�S7�Ҭ��	O������:�R��Q����E�,f������S3
T}���iזג[�|<A��<j�J�W��r�v^���Z�ԹB��V{��6�<�U���9�dnn��Gr��m��G\	��Lb[��l�K]sͅ��\X���.g+�v�D]{���[!�S�͖p��	V�2e��nǅj��0�Ó�\��sUUy2ʌ�fr�K�Cr̔�`v��^�W��̷�|y@��4/�\�����//�Ӌ�H���KuIY�a�V��S��c7�3B�^:�s!�n�6������S�Vmq�������m������[M5U'|}Gu{|����^~A�ߪ�~F�Dy@�u�]Ư�����˭SWO۝'�����Hq�X�]\ҷ7:}s��ݴ�R�o6᎚�ݶz�ќ9�2��C2���dK��խ�X�Ue�\�r���Ξ��/Ѡ,��4�Ӟ��P5�\{pkY�t�3Ϊ���[�J�/O˼\�-
����}�p��jQ���w|I�+��b���\�y�>P]�PM�`O�~�S�x��a9��P��T�@4��X/q���W�����.`uz�!:��D�E*4{��ʏ*���>!�f�wJ�ί;���فV�N�7^M\R�4m�[���ʎ'�:�iB��*�5���=m;�#_��<��篾���}�{����v]����u�wwtd�*JX�@��߆�V?����~��dg�9�A�/1,S�^�972�s�ԅ�s��������5�Ifa;7]h^��K�=���6��v�ƥ6$]��v��.|�ɟ�	[f�������hSx�m\�
���zĬؽus�J���-�n�W}���־�����1^��j��eb�)`����!��x�}/W�u�NȇJk=��sT�=�Z�ْ*m{<��������S�F4�/]�����[w��v׏O�^ZZ���ayF�o`����!��t�;s����fu�N��z{��/l{6{���j�Gs %����nAQ��U�?����1g��g�X�r���m>ߢ�1wy��g���oY�Mga�T۷�x�̈�����>����>���˟hM�FH��nw�w+V矡����^:6�n�6��u�ƞZ��c��:�m㵿u��"�(�_
���S�	�l��=�Y&��]���l/!�7Q'������uw]�]�62}�{W8�݇N�4�s��Őt"r���0�N�Yn��S���Д���/��&F�mk�Y��*;�:�̐��֝�1A��>��ua��ٜ��{w:�"#�e㦳Qi�X����ݾ�lA���"԰S���Z��Wm�,r�����Q�ὝS�������9<3��-�R�<t��_����N�۞e�y�ͦ��0̺X'����*n��rMs	��ᵅ�T�ӻV��O��%	����1�./��o�(W�+�d�e��k�s��>se��y��ewsN�/+���<UL��v=tg�$Hw�u�\��3x9��1gۻ��M�T��7C��ens�WL>�>:J�_��>��3=2�;/q��s�
�?��ݲ���"KZ�r+�WK�ݜp-kHj���h�ά��׾�i[���j�^J���eb��U�A����\3���mJ���2#o1g��n{��o_r]��Z��UQ�����ͦ�z�>)YY^z�W�%�[����!/���]I���j'iJ�
9z�n�eH�sy@����u]e%'ٷ�ѩ�\hcy�X�����|�s�Gpa��ݵ�k[��-:`S�����+k�H��bu�Q�\%^U�6��R�"L��x����|~���̀q���г+�j���?K�kOPdXv̈�������ܦ��-������K6;{OB�Yxu)����
���TgnKZ�kX����e���ݺJ��6;�[B]ڢ�X}WQ���N�v�D�\-������x��ivd�cqY硋y��3�ɗ�y��[�*tli�b��:;9_.�hFh�ư�4�3�͉ú�����2�j����^��i�2�ݩͯu��7��mϛ�1e��z��uC�z��;o��B����n����3z�����ݮg����8�p�����
0u����9�"��#롍�c'lf����.6ֵ�4�v�]P=7�ZM�Y�o��:ħ^v�]�ۼ��һ��u�/P ~�������y��tV�k�5�Pel(!&g��ۙ 5�w=�M���cm�����e'Z�Լ����<�$��^ܰ�t�6W`� |�Ǜ��%Յ��C���2W3J� �pv���]'NN`nmuq�\�nZ5��u���V3�sRX�aٲ
=M�Mc�}U�o�vl�:(�ٲ��l���D�9k��������tck!1xT�8�g����/w��i���+m�ԥ���5S�SQ/c.׍Ʋ�{�k���#o�$��5�vzy�H<��ȵL��A��%e97tSs�鼗��;�t�6i�@�a;}gϽ>�J�r��V��u�)��������pd��'{}����zj<˖M�a=�k�1�R��Vm��0�����������  9��p�S`�>��l��ޕ�K>%эۚ�O1�i�2{#���C�Sܥ�����������X�dђy�j�Mw}X��_�oUs̻��p�����Cm��{"��gg�*��`;�ݒ�{f|��7��'t�Ιw#����Դ/"�*)Qw�8�d�,�J1b0�;({̹̾�`u���!��{ِ���e#nZw���>��t�F��F	�y�}&������Tz�kX4o��M�)=tnl���ީ徑�f��ޜ����.<�5k9	�wu;J�^�#@>|h$k1�au�
�8�X�H�ŷ�n��ɻ���A&:lp���D�]��'n �ˠ�{J�&��dt@ô#�!nwuwWqu���߷�����}��W=�E�̀�[�����ߵd�����5@}�jĚ)�o���=��+^Z������^��+���Zg�W��8� �8�g�۽��og��:�+��_�kbܰUă�-}ي}b��U���5>б%����,ܪ�����f�c��ie��kE��;�Zw����
�Ⴇ;7[k���奂��)X��Ty*b�
�6�N-�#�:���ऎČ��͛O>�C)>�3n;)���ԅX�z���@�L�6t艍�j�+i�V6��fu���#��UL$�DK�*�t�t�B�*���Ό������ǋh-܎�zZ��{��R�Y>�O�FjY!\+��[,klf?\\[�n�3��,ŋ�!f!ʮuKX�+ ��u\7%Y�Q�-n�5I�����*��#[o7va>\����D����+ُّn�S�F���h>C��m�m��y�Τ�}^���1�+B�]:�V�}SR�*:�Ӵ��m�Ya5	Ek[�Q,毢��eAo��x���IO0��f��&� �9Ff�KvJv�>̔N����T����Gjwu��Z�ז#Op��$��xЏ�7` �m��z���'��̔-�wP�^W�w�=:*�>�������,�1z�N)��7�$BA??��3ʅ�,�g���.�m�v����2���;�g�]%����1�����ٻ"�^yDz{:�>����Or����Y�C����fFp̊��r�;K��޼���yߗ>��Ҵ����un�G�}YSqhd�Ӵ6�h�~�ma����J���M�6s��T�u������ۉg���X�
1���7�����->;����0��Ԕ�Jޔ_�ES[:Z��'"mpkd�o�̯j������@;�|E���.5���AN�uNێ�pe���H.363L�@���7C�y�_`j�lf��24�!������x<V�>7b���:����%3��J,��u��(�Gw�&�L���2�@x�����F@��hą�j��䥝��u=h�M�G`
�7�0��_[���,nG��Z���/Թ�C�;U7�ίC��j��4.��E'.�����]��Z�Vac,�U_���\o�V��C%]��`��/n�E�>�v�fw/k\�:����m��y�u3�\��+�F�ϫ�޾���
!)�_�S�n�!Tov�K���i�6cϻ/�+mOd����d W��Ǣ��@�\����ݥ����0֞5]��xy��=��m_B��[�ޘ��e���j�&����l��d�)�+�/���s �Cxts޿F6�o$����bi��-SG��h�n>�)Y*D��cF�|q��I�wrht�"�,}R��)ԳT�\�u\?e޹J9�[�to���8����ඖ��J�g����m`�}i�Ƞ�:)��8V�X/��1�����C�Ͷ�e�'���ko�n��t��w������vN�^���i��!��c��|��߶��E8ɪ/O����ܫ��Zϣst�mR��V�d�o�8:�����;�ԱP�?μ�9ۓ�8���f=��v�z_������ꂝ��h���ŋGD��XTo�j7cv��N�Ѣ<��u�p���埚�a=*�<�\]��.VN�*ۺ���/�7�*C]�{]�Le����-���o7�Swo䮊u��v�����^F�,�]Y]}�_���_��}������@��q��s|���yM�{���%� 6�8��D���l�n�(6�Î� P�;��ld���_�O�,fڸp�]�4Bu��;w����4H0L�[�q�?_S�(�ޭ�Tn���yΚs]�]'��������Tk�Zz$��l�.�����\	�C�!:S���C���sTk�-�/rC#P�$���Ʃe�6�3��aMgEH].�M���y��v�i�`p�3R��%s��ȷ�ϐg���`y�3�p�1�Rg�K76r����k&��;}���[��)�XE��	L���p�\�UV�}�S7���l�Ҹ�r�6��K({�J�xs���yD��G�65�X%A�Vi�M�L	rO"�'�k]�����N���lX����lM��-QS�;۲�� �G)�y�(�S�m,�d�m�f�\�t@ǉ�ޗ��]�;��|hI���d�;H��������>�!G&f�+edh�65�%m�v;s������[uy]�i�3k��B�ӣR�c2u�4���n�.ݥt���puu�ux��^��`�BN�ڼ�_k��N� �*�w�1sΜ�����O�������{�7���o�0�p�,7:�b�E
�<J���7���D�ݾ7�M�ϻC��kx�s�q Gzl��i����wY<�!�m�t��e>0�ׂ�R�ŎZ9�;{�)��<���)f��l��&��9Rv�"7��6An,�����Y,���zNB�t֞!����a2w1M˕��[�!g��Q����bm�Á�oAԢaV��|����ڹ�[�B�Woq��^m���տN�ռ�ī�0zb4&����xl���˳j;<4�bK^�7�M��o*j2㔈w.�oH�ʵ��`�:&eޥ$��Ӻj���PÃ.,���v���8�������|�v`�y�MD�
�Φ%���yaA�eL����T/��c�n�<̝EJ��Kn�	c ��W�mm��52>��i[�m��냺5���C!�;����;3��*T�_��}��,m@ކ��]�n�h��Y%��.'�b�X�q-3hi�w-�^թ�S����;:(�U�M�&vѿ�v�owT}��-0��Z*ɰ�Ā�t��U�u�K^�LM�+M�#�*V�h�l�HTgZ�y@����$D48�'*]���+-��}]51�'fVP���V%J��Ȳ�3��D������]�ޫA!�K�����ޤ#�v����gg͵���	��ŷb�7��ԛ/:�JO]v�Z̦v�Xu�m*
�Ϋ��(T����[���K�ޮ�ի�&�P�l��:���:�n�*�������-���3:�ƾw�y�蔫�N4�Ρ�Q&q�Ȟ�L��5lLڝ�0����������U��6�:��+�0�F��ע��N�f,�[h�*�*>4�s���-ؠV>ʷ�:���3��^�Ü�,�N�z4D���L|6K�hN�ʭ�Uϻ> '�>�hǛ�e���Ęm�F�;Z/��N�ͺ(7�p�kh�\!H�	%n�֕�oeՏ�wv�)���O��o]�	����K����쩳{$ �s�/�<�[�+z�u1��WrTS�(�@���onî=)M�xf�F���}ƕ�����U��ԕh휺�1�P��r����{�&�9q�a ��(%��G��\y���G0&�ɗ��&Ii6R����R�\� �X���$�F`��6�@�HҮ�uNrɳm2:��N��5k(�`�A��|�$�E���Hda���)qQ�)�(� ��m�@�4(�I�L$��Ii	R#�i� ����{�ػa�JR���D:T�l��%4�%:tAI �C���-~�1ۮ��-�m��ĕA��Q�RMlb��߹�K�6��E^w�?�����>����?��g���c�ն�E�t~��)��Z5z�::{mT[�n�ӋmE������������������+�:�4C;m��Em��wˎ1���i���j�5Uzƨ*(���P~��<��~�>>>>?_���~�?>E�84?q�Yh��>[���5]����&�Q�Mh�[V)������/[��5��"<,�Gm�y���N��b�A���Z#o7��116ƍ�D�x�ƜZkA�(ш��`������yƎ6+X�AZ�k[���[�A�Z��ϓ�Y�*=mǮꞋQ�-&��u:��V��[tNݺ�%i�5X�h�w]]py���~��A�Q��1�Ꞓ�,b5�=m4]��M�[QDTWV:�f�솢����󎃨�cCA������������
5A�����m��w_`���΃Zke��X�(+��������]����t��,N(���{����`���ylts���T�t�J�"��EJ�! Ǫ��Y�}�#��l�T_����gh��Kl�]sO������L�}>�~�}T ��3��E����jnZ�{�n�y^�L��;b+��D��e�d�3����R��#]��'������̤�i��L���#x@�Ul&v���l���k.=�d��}�>���^�_*����\Loc�0�עp_<�e�kC��2��#t�+z���8k���/�*#\���(挳��������|��v3���`su�s]����k��2�݆۪᭔�׻v��`kHe�Cx[�2vW)>7=V�&r�x+��Sp�P#n.��ʭ�9J�in�sh��5��q{�طe�۵������4E�{�q�e��p!��%,k�J��ӆ{��C$tNP�1v�_{[F�Ow�*`J���x��z��^Mo9,�j���{ԓ���p�i�U����r�k�ܭ��0$`��N7�t�ӑL�E����kP��J՚�#�˷��*CǼ��}W7 �|>�&���++�U�R�u8���epY7���*\�6vx��;�^jvL�S�"�rDW꯫���^�c��M�oiSO�ltb)�SR�Ϋ����+�x�E��nU�ޒ�L�AʸS�x�-NR͢�ƥ��4	��$��9�P�t�sUP�j����S򶁙L��Ί�I�I
��}��5Ie2�W���m�vV�_mt�	�Y���&���n4:YL:ș�v�3�#tp{�؅��:���ڧ�,=�>�K���'8��k��zem�����TS��t Av�t>:�˰��%�^��j��s� M{�9p���M��r.���pg��+�7lꈞ͉��)n��jژj��7��!Z�� ��Qjr�)8�
]@l��WыP���ݒ�L��[���/7~ju+�=h����v���b��]��M��u0�
��M���[F�Y�ڪG^�����z[=��o}��l*k�[���l
��`�6Vɼ��)��2�R6�L.��V�$.�tK���x�sj��}׃��Ŋ�o���>��EY���i�݀����=�� ���3k1ّ���,Z�:rz���l]��m��m]�oF����0��Ѵ����.�z��DttR]o⧠^�F�u��t�������6��&��!Xe;In����v|��ˉ�:�:��[���t\��ԧ8�t�^���i�N�{�:髋�8{�=b]���N�#s��ݽ�����+��V�9~e�&�˪&F� g��ڒ��ک�n[���hă��PW�'�3[e�5���nU�ע���b�zY���jG�r�����h��IW;7+j;H{��q.�C����	���F�B�~��������S��h\S�7�����-��=��du-��JE*�J�f��EY[5�D�1y�0_V0�:w.�&�v�!^Ǳ��?+�Kw�ثb�hj�sh���\"x�u6u�L���l&�����u��Qqk���#�e]��]y�k���S�\��Ƚ�0�����m�Z+���Iyt���Z�~RΈ��^lG�e�54�K��I�u�M��'}�m�׻5�%.�lWy�؍(O^N,Ӥ}f�QH�۔�����wfΫ>�|Fu���ʌgrUq�RП.�ΚVi�5��^R���Ks��g,�a��Zl�����霛���3�s��뜌���#<��n���B���{��~'��c�������K{�y��Z��4�a�U�;dz�l�5���;�'��̮����`X����v����W\������3���:�Y��S]u��	����}���͝��j�+�oi�Fnیާ��{5�CD�FS��^aP1>��ތs�EJA�VǅG;*pj�{��[�b:���mC��3���'n�xs#�DI���Hg�b�@�AR�_��"t�]اޣ�s���������.h���@en�x��{����ݎ�g�z~�#n�i�?PS��oޗ�= �G{xH|ͤg����<�gv<�(�4�+�����:��9uT���"�-aNw��6�C�pv_�Z�1+�ks��9�w�]�)Y*����{�.B�g�T�b[����Ev�}s�r[�֪�*</�A���79��ܱ��%]zZ��T���iU���S�l��AVS	_A*Zb�X(��x�u����s�(�VU�R%Ĺ�7�@S� ���ƭ
�7��*��ċWB_Q-.���yLRt��6� ]�(=U�$�3�^���5�7��(�����7�h��tzy�U=�w�\G�S4В��x������^�g1��ת -5��4�Jα�ٺ��o(��Q]�2�v�����מ��	.�x���/C�i#S�dފ[~��#�%c5G�+۾Zf�)�⻺ojm{u[�ꊀ՞G!�ezw+t�Zh�F��*��x?D�n	�t������Ԩrݏ$�d:�~��k����ёY�p���9y<��Q�v�)�����媇���.��o�O�,,�;y�ZLf�MsQ�ݽM5�w��!�u�4	%f�o&ķUpd�Q��F򹙬_�Q���&��!�q���6rw�Z�iTKe�;���=��q�T�Xo��������߹�{l�2���<��tT'}poUH���`�W�;���u��S��=�܊`{��G�+�]J�����m{&?T,�Ng��.��8�����i�x�dP��m�A��]�.:��;ަ76G17ao]]�>"��ܸ���UkM�3AS�C厎r���}�-��}ч�~Q��;ӻ]g1�����Ɓ1q�zY����MnED�]�wF��Zy��Hu#\ʆ8�,�l��D��AS5����wL;���׹냋��H��Vs0�W�qG���o�ϲTq���y���a����s>�e�,�22�B�.3_�T����O5yW�<����wB�?E��hi��*�U��DL���aUz9�!Z�VK&���� �l��}Wv2u�1�e�:M#Rs�iɧι�	)�C{Et+��hR?�H�q<�	�y��f��~�V�_����f޲�!B�ǫ���9������͹"'.s^���SrWs#�3�4VA��ʽ���75��,�����zc\��$�wzP�ׇ%�>�����]�fE�/���"`C�>�u�m���ݡ���θ�Z�s��	c���Ⱥ~]��l���f�ݯ�v�|^轁pF�c�.�q��𼅚5%�s %�%�ْ&��M0���i����Q�S��,+��34.œ���vr�ݧ��V����T*�4FT�6�o8���}}R���R)�t*�}�T�[O����A�:����\�63ۨ!]5Ŭn��ں\/��݁�ee��}a��M�pč�_Vlyo��m�ɮ& :�;v��ց&26�>�v�p�Y���t��I5<��_��6��|�����9�m�oCϡ.�Z':e�k�T�����Kk��4\wuNn�Z"ޱ���������m����ۈ��٧q,����/�����]XV��}���b�o��8�MG�ZY���{k�z�Y�1v`��9|Ӑ���lZ=V��*{ޘw:ۧ�x���yŹb�9�af}�z�4�}���n|�r�VԬ|���]����F5nYbaS�I��Cݩ̮g��n�y�+���j�X���v�o��"r�n
O�����/��8�5���Q^�-A0�N� mMV8�,"����;U����ѯ&�Ow&�\�K�2��>�=�:6��`��U9��u�>�trF�����ݼ1�uyd�Pmmk�p���!���×9�~?�Y�Q��^���H~�r��'�$[�^�B�;�t��d�qLsBP�鐩���)�(X�^q�|��n���w��v1^����ɋ��l_K�B���-h�ۑ�[%o��W��0[|/�O�
��vL��@�����˿�W���>��ޓn�ﳎ:�]���2�J�t�zW����Û �V0Lt	ު�u���v9���}�;.6��t����S�U@�4�C5��������Z��oP�Q*e��.���Evݵ[�ϞlOy㏪}�2�w.�᫔�Zg$Nv�\�B3��[tS�ɇ]we�ж�Oq�J��=�H�e0�^֞����=���_�{�τ�G���#�گ?R�cT��J�,,֮ʍ��;�5�w)�Z�]a�\+���[�u�zů�Ȏ]�q�;�0�gy��Mm�|��.�:��+���ve*�.{B24^��,N � j;k�eM9�Ӹi��mD�Dp�vj�j�Պ-r��1����R�>�S���k��*��kH����ޡ;�/���
�YU�1���7�����U0�FM����W}g��3�ՠ�=�w���*�*����_o(��&���oT���¨)pa��n���s�Ǯ�.�������]���6D��6xV\�ά�`�c��/�$�iA�IU;	ڰ)>���ѣz�tI���M+-HTi����b���Z��Ԏr茾��y���:�v�Qv[�q��DՍ�ؔ܏Y�%���S�c��T����miv@�\�Q"�HM��|�~�{r��!�jl�Iwwc�����ν�??��T�vk�i�p��S;W�oFh���F7��sׯϒl>AͶZ��9Ƌ�In��ð�-�܆o�������9��{r�(�܅M�ײ�v{�_j8[7D<�FT�	��^�rז�W���K4�}*��ف��'J���Wf�;y�x�TQ1i<ָ�S�C�O:���Z���\T=N\%'!���hL�*j<ݴ��M��>��r���3F�3���Fv�s]��9|z����-Q��d�=�>|u�zL���j�ʁ����;*����4�m.]K:���US���X����98:D�t�g?���{.����u�>���{�;��|��~j���߭�g��{ %H���H����x�mh�sz5�K\�&�3V6�f�9��]r怯��rv�]���gŞ��~�����~���c�f&U"kT)�ʵJ��K9P�gv�{����qe�OP�X239Tb(8�9��E�vt��=�zzG��*o���;oeZ6�v�YD��mr�6-��K��TT�3�݅_�����C�N��r�ڡ�{fS�1���L�,κn�+1b�˶�<%۹lgF�f�#�,D�)�,N '�eh3ZV"1�� �*���g�̤�ך��)tuĻ6h~��Ǥpi�I��tz�8k��]\�f�m1\������h�~��5@~�݀w}t�+�}"-uz`,���u�0�Euk�F�#�N,�}ڲx7"�6A���=o>,�U�j Kd�VN�lb�u������rs{$w
�z4��p��Gh���ܜM�����	�#uן)3թ���E���r�T%L{�����,"�ޗia�����M��;��L�=s;�e���4b�ps�g�T��[F�¨PW�L�5�G������F��x����w�v
�IMRӻK$c���d3�l�*o��{]��(��r ;��Ѽ�6�U8*\�� �=,��ߣ��x~�w��de���}6��yN�������_*�T��k�6c�˞�H�2qd�h�pe���,!t��%�drL��H��Yړ�zo;X��q̙2u]��ΛЮ���,P�	��Ӯ�|���uc5��8��$��[۔��+��b�f�qk/�i,��1��n��:�-��m�خm�\4����ӻ6d*��d��,?�*��ܰǘ�(:�C X+�������ئme�_f%@�'GЌ���\�*^�5Cq��s���a;ֹ��uc�ډ�år5��RW^j���k�,dB��&�0̃�^��{�� �J̤���B�\��e{����{�EV��\�R�E�٭�ͬ�4����Y�sE�N��[3�������Gi,	^vag8�t�1r��&2��Ц:T��+����eu�w�r7��Þ����;N�N�aw@���8�pa.��ۭ=^�u��'2�����\0IvރήrDF��n^^$d�c�'T�t���9A3�L��� Nf*閥W�M<�;�M�m;p��꽒���vhTPq4a�!��jigok���w�ma�RӅ�Ѐ�!�ی�PSu�\���l�w+I����u��K:^]LLJ�F��[AEF���;D�e��ͮR1��xN�P\]�zf�9z�,�,S��P�{r�.YwZE*$'�\�c�\���6)cJ���F�ZW(��n2� 4�����`��yrZ�u���m:���kU��+h�FP&j<n��r����W������P:,pk�9לj�S�զV��T{��2��j�X{��ы�"S5�i��i6qz
�R�ܷ����^ݣO��ά��{��rsܑ�4�)���+,����?���ш��yC+��Zj��\g
E��K>��<�\o����ηx��+��p��l�Z���ӑ@�qķ{�o_,8���L�o�Mu���Dn!��q�oy���r��[Vwo���J_JmIv#��i�(T��n��յld�:�ɰ�Φ���AqX7�6W'{bֳ`v��_VX�	�1�6K�>��]n၅�L�L6^k��B���U��ͼ�H��r��x�hIT;Ic'�ێAn�j�z#��dq���޼�����oM&Rs�Ճk1��W�ճ�&�bd�E&�ύ �s�S(�noEA��id��$ܰ�����M�-���Ѷ���-ȩ��[aȶ�i�h]��K���Ԙ&]�]
-��GE��h=�m�ۧ��Swi���t�Ы�س���n�SV(��you�@�v�n�ٚ�[��l��U����o�Q�l���c�nhUk��q���~�E�Ƈ{��{���b����yyn�u�hI[�7�b�<�<��}���������ߚ����k����c�&-����yW@m�u��D[u�Y荝x�g����}>>>>?_�\��ϑ�~v���4|.n����Sֺ׫�z�Nh���(����-DE>[���
4�
��|y�y��~����?�~�������Fڈ����j$7���X����bjf(�%��f���b�l�A��a��tw�;�<�+F�h�6�9��R����+g1kAV�X�֓�kTb��5���D�TU���Z���qW�Q����j6�&�c���TlU:���Q$�4QD�F���vԛ`�=F�!�m%�(Ѣ�Dm�+�=5N�-�U��cPF�D�m�Z4Q���D�c�Ѩ�H���ٰ�*��5�qq��V��b"H�дAE�w�MF'}v(�ڪ����`�U�(�$#gZí�h�z�QP�v��_����X�[��3��䱫����X��ӊ�m�T����@�t��������nnP5K��궒���UWתX�����h���\x%[<��h��0�@O�C��ۗ���ҚsG;�v8����������tKvk��z�#U��v0�Ƈ���)����B�ᾗ�I�[�%
�t-�WuV��v�_e?qŏm��wA`ܫA�[� e��d�:��B�T{fρ�\�6�>?_+�b�J��:��G���*��x|�ΕlS��ǥ�{: ����d���(��٩�xz�>�ܟ��ǲ����d:�f��ޛ��A�0���5���;�2��ƨ\���+{pW��冿g�u>��$[���ܧ�̳�EFG�_wVn)�u�tc�z[c�|o���9�,ҵ\�n�nFV���[��*��o:��o}�^���na!��C�("���S=��N<uq��q��p��U"{�
����3�7�g�����䨰����ͷ|z
��\�i��Rؠ�է�;�9�2���;��f+M���s�+7$����-=��╦�G��C��ok{; �b��ݎ�E������/�ͽ�w)�� ���?Yύ�M^�׹�,.�ώ��q���?Uv��]�mCcL�ut���6.�n��;�)�^�Me����׷��p�;��c��ާoZ/�g���)�ʷz�����Ƃ��[y�΃���.��!��m1pqK@�5����C]�:�K[�;�S-U�E������%����oB�t�k�6{-L��Y��9������IS07M��E�cf�md����X��-.��[��}y�*��5u2��d��s�mEޫ���y+�R�w�,
5�/ҧ��X��T�$�Z��UZr�-;�>�3��3;[��T���t�W
����]�j�u]��ڋ��c���
ޭ�a-
P嗭�/V`�7����Z��M]��l%��ZF�D�H�^�������qU����ʗj�Ű�i�`L��X�������m2��7����ݼ���e�p��V�:³��>��]F0t2�1ۦ]=O&z�jfұ��>*�Ru�����3�r��E6����e��x����=zǯP�5Y��m���̫U��Z%K	^թ�r�óF�;���T�8�j���ڛ]H2�W	ے�b!�x��;q;7������}���-�*#k��LS*�m�D�LA�1���g��I���ٻ^�g�)d�h��Wuڤ9p���@���r1��L�3&�����'}�~P��ջ��ȍ�$�{�u�}�|ާ�}E^����u�ø�{����K�q���^�o�V��%>�S>9���&H��'���&*���S<�ok��h�G�cx�;et
��m�V��W0��R��0SelQ���*P@g	��
C�?��gu}XP�׾m|ԞVK��os݊㽽 u�7��6$?t��>u�p�˖�w���\:�uK��ݢϧݺ�%�Z�ys	�Cx[�d�f�Q�}��c9ɑp&�[�hw6��ks]d:ف3��EpM7��������L�_��8����/����5�8,�;�� ��I��r��������u��K:;a����F<�Rw�	�V@��Ȩ~�7�h���I����`6��N�{�s�!�(t�׫���o�A���J���ѝb�)���!YX��~��޼�S�`�~;بL��2�P�<�`k�� �{3�i;�W0�<-̽�&�ֲ=!LA����A!�1=�*C�;�.�U˖7���s~�����ۛ��Q�"3}��fnz�@�Z�Va@/�澙�6��^���W)>s��V��}}�-��� Jͤ�"U\n�<�S4���Э�M� ��s�LLU���C�*Iipږ�7^�;
�-�IV��~#gr�`<�=�v�tk�k����:�����>�
��>���Λҧ�g�9�*"����A�x��;Z��l�T�L�
Oys��J[��̅��:��T���ڽ���V�\��췡�w�{��唻p�g\5�f��/wyt|]�5�	�R�lv	�z���e%}��P�5�O�k0������Ǘ����*��-�;�@�$�v�|]�S5�С:a�'�K�_FvsL@���n{:[-l���;�c�r����7��y�h;K��ǃw��M�����d\SY�8l�o\��^���T���ԟ������&q]m��9�Ù*������=�nV"�'3��v�Z�l��K��5�b�����3��G�^�R	�f(�6�9���ZN�%����B&���������&�����G��2� L�0�}�x=�Ǳ9�S���9���E4'7�!5���x&�����w���i0�7nZ���M|4Z�C�85S]�犘��]wZ:�_����\�u�Qw�z�f�UN�^ͦm�fT4Q �]5>�O1>jT�m-X���z��ˎz|��io+��nꤳ�+�C�H�u�^e������ࣳu�`N읞��=q� W)�J�yK\ݲx�oG<�]Dmʉ�έ��r�7n�z�[ ��ye�K��ޚ�*%f��븁�훙<]�3v+���o�L�ad���ԕ���]G�^RX�d_;X���/j�g���m\x��1��CT��q����������l�p¼�R{�n:?���ɓ��Α�C�56W��w5�8�;���H�Klk���k��8Vf�[��9�lU~��� ����|e�!�'r���+����i���nc��վ�aYKP�fd����6�ށ���K�v>��L�����d>WYM���Q_)�Q�փ�Z��jZ�&NFƥ��R.�پ�÷��֧�o���u���zy�j�3�}�k�����WS޽�㞑|+7ۦ��t1�К�.�u�m�]e�i��؎t�H(��-�@7ʀ���r:��:1���=��"�2�-��3�\l�N�}t_�����D�~�<v�0��V(���w���:����Hkf��]c6���Cd�ڽ�l6{�%�qO�!F�ީ�ئ�{k�S��{}�\��r=fT�)d��>p�v
�+���ۖ�2��W;���bV#��4~�<��i��3y��i��=�������%F�����RL�^����˶�b��`���M9��S���f}PϮk����� �iΥ�3�佶�ѷ���k�iTz�i�W�1Re���[\ײ�Wsa��L-+c�S��7c�j@7D���R&����d�]	H�WJ�f��VMk-v,��ޣhv�>-hj;����Uc������'۸,J�[�1Һ�r]�-N�}I�
��v_��i�^�_�c�K\�vP��[w�Z�/�%��
2qi?�T�Zh�F�ȕ��Y,�]��eķ��CN�$f�F��^F�]N��� :Kw�����]��s�qs5�Py.���g`1,�M)J
���/q:���B�V[�yع�Ј�)R�tV�)ҍ�T
�0'F�a�+�T��ދ�����x����O��a�X's��1I�a}Ei֍v�OU�5W�vLE;\V��:���B:���CKz�����B���v/��W�L�<ϓ�{���:�cw=&�dywRe�m��u���,���&m�171���;Sۏ����{%���VK�,h�1^W����r�[Y
���/t ͫ��\�[�+y�uw1]r�"6&pZv��N�u�N7\�QvnGn`�ѣ�,��y\ ���+v{�F��u~�j��W��Um���#�r�{蕯k�����p��N�����j�כ�>�1����MR���Y>z}[�N�ݘ�L�]tP�R���趎SNf�m����^i�ʭ,�N�4�r�.V���L�>냼��.�'O�N��Uyy'5�H.7x��w�h��o��eb�=9�����Z	؊��t� jh�֪�#������+���wZ�c�������:Q�=��p�9QU��k:�j�
���فs}(�6���V�]�s����Qju��c��L�r.�[ ���ki64*<�NZq��zm������c �l���k�*�w�ۼ��.��,.�'�\�����l��l�[1��y���k��{��_x6�Z���(�K^P���Y:�.F+=��D��d��O��/��f�������"�uW�m�NY��W:�ָr`A�o�7emNlC�R���38���̹٨lU	0�}z�B̭�'[���us�����*=�T�o�M�MᩀM��K Z�
ӽ,�:y�)���f~�v��n�*S�����݌}�8�!�,��[
�p�zKFFm������y��J
�U�q��1�4^¥�n�]Y/���Ni���'�PWOo5]l��r�2	� >�����达l�`����;��*�:\��gt�ʊܞ���P�7�v��� C��S��`d�Z��%sn�u��6uh�wj"��vڝ{}��!��)�O�����|�_=$޼�U|^!6�ͻ�=,0�SV9���R��&�q��Տ�qV�Lݔ��*DdU�@�㧍-Z��"Got�x�W�%��1@�\�F]�ݽ�h�7�;���=��ye4�!���F�e��_����e��u��@v��#;�l;�/l���}S{�t��j�h�{��y^� ����9��IG�����B�U#8l�~357��P�ͤ7%�m���\���;�F�G�tߡ�h�M��8>���w�YJ�v[�����߫��$dT���`o��}`k��b�S�*�����Ul���w^���sy�:{��=��r>���M�UsE��ͭ�odfέg�k8~N�k�ꃒ8���^hS,���wzgv�q�xv=�&��f�>9��[��Sgˮ��sv�=�"'5n�ؖ�B8�}m�ez��l���aK�LU>u�`��KB���ڻ'\����Es�'J���n#����+c�`T��_����YOb{�w���|����W��V�����r���fpn�}n�ODI���/��v;]Ͳ���y�ވ�Ktk%�r��o7��W9�0^�U�{)���d��q[gF����F���6���Մ��ȱ�`_$�S��)cu�L��˻�M#h���Zw�=�`�Q�҂�� � Fr�\Ѣ��G�����ڼܛ�-;����\p�bAoc�vC��q\j��p�v�˙x]T��{xO7eJ�=h��)]���㰯)+�1K�O5H�l3��Ӽ;^����6����	kpܖY/�buaW���Y#G�&'o3H������޾��l.۟O�9��B�we��[�)�ǥ(�SY������]c;��ncs�;�ofn�jufn2�{_�U�y��2��h8���Ӓf�r,up�o�m��7u����k<qŎ$6��ma�K\ő[q��������w˽X7�nz��F8���F.���/����n�-�f�Nh�#Q�#zC��\�e��1{�p��<m2x�˺|�����h-���qn���#bT'���O�������S�0wg�yL{�_Ӿ<j�}�6�>f�>�iu}�Eߌ�����oB��$ݬ������D
���=C(�G��lx7�z��~���O�=����͜��$���$HG���?�d>�B3�jMMN�$�Ru�S��3� �B!���hf���HB a�d�U!���Hbd�A��YP��Y���II�Z�4I	3�L�"I;�C�vP�+�V ;p��+�!�@!D�@<�c�!�!(�B���B �!B �$B �$PBE �"P�@!	�@!	D�ep��@��"H!(�B�!����A��A��@!	�@!$B � hD�@!	D�@!	DD �%�@!Ta�!B�HB!D� B�HB B hdB�HBD!	�$BVP&!�I	P���H�HBA!	�$�!�`�HB!D�P�"����HBD!D���HBA!T�`������{p׳��ܩJ�JYd��e�N�M��ͳ�﷛z3��~�5~���{~&�����٦��z������$^����Z�T�zv�$X��s0������#��I ����=oT�i���7�y&�CNN�љ�U�J�a�%�	dBBD$ B �I	��HP�Q!$B�B!� 	�%�e �!XD�D�Q%T)��!H�!H�D� `R �
%`%R(��JQ$�H�HA%�&b&YTc(�Wd�RhU�D�
EA�P�B�H%�P�B�� �H��	!	��D"A&D"$�aP�	$BHP�D! BdB	�p4f�����|$�K1Df�Ic���(�L�_���LbK���ċ$�'~���H�ߙ==����Rk������e�I��b}?�{�D���'ʞ	�"����Uz#���: U���u&"HI1$������p���_�0�����S��8 ��@ǒO������$9;LbI׻��O���j�m:OX�2yv�Ţ�Uk�'��$�<���d��N$��ߢfx�c2v�Fd�珶��rO�7�0���DI �f�0�f�\�MC~�9���sO�q� �<GI�=Nx�B���ן���is�1AY&SYD�H�4Y�`P��3'� bD��^�H��"�*��IT�$�Q$)J*�D�������D�UJ
D�E�"�"I
�UJJ���P�DS�¶��ZJHBITEhV��P*�M��B�5�J5�����U
Q%B̊�Sl(U$�$�QJ�EI$}1P)*!$E"�)(UU�*��J��T]���� �E$*�URIHi�Ɩ�ID��@�UIA
P�B���  3GM�6�b�j��jvi�[JV��J�6h�M:6��6��Ms�Wh���Q5�֐����+J��,��*�kV!m�T��Ru)B�Ji���
�"�O  �y��"�
(=���ӡ�B�
$H��p�P�B����o+�gZ�M��4wesFm7v����fJ+��F�Fj�
Y5*Kiݵ��ki�PR�aU�
UT��(�O  +�����Һ��T�Il�s�1�]�vƪupm��j��r��ZC;wng*��*ѫwuv�����j�5�ѹݙ�[h��VҫLݝ�$����)P�i�x  0�!���0���X3	Tl[i��Ҧ�ڢa�UZ+�� ���F�U�@4��)UT���RR�*�JRR*�  �JSe0Q-���[6���u�U��B��)�UT�NA���3ݝ��U�� ��ZL����EU(JKZ��   9@TFb� 4�n6ٕm�Q2`���FmV��m�lJ�S�]J�#P
�kj��A"��MU*P0��UB�IJ��   ܈��*a� 2� L�` 4j�  u�  i0�P��]U���� � � 2QD"�h����   6�( �qԮ�S���;� P� �N�@�˝  ҆i@a�PX �R ��@��J����   ��  �k� ���:p [;g 4e0 :�S@��p �ҩ�V�0��*�X  ݚ�����T��x  �� ��ۀ �N.  j��P �  t�� Y��  6�� A� �t;� ����U)P  E=�	))S   E<��yC�  O��I�  50hʔ� �	2��U&@ �T"$ �3��2'CuT�܁���51Rc&J6�\0S�Z��b���������n�����0c�vlm����fco�`�1���cd��m����������R�$��w,V�t��U�w��>`H�r�2��wJ���]�ڏ
n�U���'.ȏFf���XoY
V�W+t�ʄ�чhmВ�m��ˁ�b����m�tDT����d���r|D���H.�ә�XC�^\h`a�1�Ϊ�`�4��8���K)	Y�&�*$�oc-f]1y������le�'(�V��n��{��BC&)%��\��vmY1����@�B�;�����q=#�/��f�]�t2�	��z���*�u#U��eD�'6��an�	�K�!tb#/n�` �N�w{L���L+������˦�ҷ�/j���v�W<c+N�~��ø�D9m)A,v���f�%m��)�zjV��Mջ)e�Z�,-Aڦ�̈́Gt5�r!�kS%�S �Zm�*��lEo@�ۅ����;�&!��9KI�k�b��I��kmm��Y��mbA��m-�ҥ=�!n&��b���U���z6aܺYR����<�[��Z&HTaP`/+2cW#3l؛�o̉�[��q���YS#�FԈ+�Vr�.����l�w�nD%�E|�մ��bˤ�y�q6$���A�Nb����v�JHJcդ#��UmJy��hh@�N�k� Yv� ]�&i�J�m]b����i��eLt�5�B�A���7�b�&M`әEY��X �V����Ұ�X-�*�A�`W��!��kMG2�,�z�J4 C�m�{* �� �]�9%��T��C]��[kZB��ع�K��mP��t�Ne�-�+M6��gj=�TA�u�(:KBX�P�8 �$Ѩ.���u�
#691f�L�Qe-5Z�OI J:bUդ�	�e\L�J	c)�[����w��3\ƃ��4^4l��a��TQ8�ks	��U�Ѥpl#SlM��I+��=X��]#l����q�7�[�j:���Qj:�%K��ַ1Q���3A;���&�p̛P㫊�Z�j�6���@w�V������	nY��i�Yk*a��on��
u5��r��
�_,�rZ:Sw�����R㩮�b�)��K`3{krX�Pn'��Y)l�ױ ̓��0t]���4м��E��uV�B����U�.ш��_=v��AK���蹳v<G#�l��X`�x��F%NT��9Y��)*o������ӸΠڠP����U�Y�0�@�VE	�[��Y9!� ]���2�G@��
����	�D�.�c������-j3����mc��\h�u��X*Ki	Z�ƳM���u+��)��8��
ז�z�Gl���L��7�
���rnir��GU�؛�g!�u�q��繗l�tV`xZE�7���
�;41Ҥ�0�rHi�SI��A:FۛFbM����AT�N����f+7!�@ku��2ܺ�32Y�K�eɅnf ��@+�G̔2`3[�D�1A���)@n���F]H~ՌW�U�#��ơt��3 �\�6f#M'P!���Z%�iH�Ԉ@�mU���ih���{PhTE_e]�A��,��[���w0٥�� �a�r�*̭*`1���3/bڵr���QM�n��� 
2�v��LY�[�B�����U/5���Y�	PV����ٔH�7ie'`���)"��u��j�q�ű�77J�٧XE��Z&2-yX�G^B̊^fEH��G�kXa:m��%B��J� �3]9�+N��e��J��'�i^��Ɔ� t���SV�g��-�12K�V芠$�+p���U�S!�F��tҘd���5yu��S��IabLjB$֬��,�0�r�%w��ݶp��KL�̵C�wi�(R��t*��W.��+(C(}�����.�CN�,�U�R�#t���lN��bJ���&%w#@�f�3{d�)�����҂Paލ� ]Z��#��7,E.��̛�W�X����^��t���R:+*!L�D�z�j"xM�Cbˠ�(p�ˤ5�x/b���d�����g�\�x�l�`�he`t.��i�ݽ�6�P��У��0� #6�W�6�"ڷIe'GI�H1�"�۴��s}}��<�x^PX��\͎Թ�<��T�d�Ȭi���xqQ�G$V�0@��ʗ
��}�fM�z�D�	L�fI$���2¡��+�*�n6v�з��n쒦-��[�mL����ӪZ�iQ��Z�e���e��Z8n��
ktf��[�I��lSv��t,�d��@���kC�B��w7*+�Q'r/&�ۣ�bL˘S���.MslcVL� k]�Ғ�2	�fm���CS�Em���=X����h��m�XM]�HJ�j�m��L�Mi�:6���5U�GE�=ci�x�-
ڙHk1�J�
�d�2�.��2�������YX�46�S�r�A��6�:�ue�1S��e�p坖���ˬ����զ�f���7�.��F��ӣ��p�M-�aV��ll͌P�2Ȱt�x���
��6(%F�I��w4 �b���R�V�2�ZQ��)���`%L�y��b�w+OR��M�rZ��¾�Io#r�l�h��Y�@����J��ɕ�@�wwI��,���T���*Ŭ.ҤL�ϖ{��L����� ��Ub�c�ALj^3d	�e���6��/�]]����hԕ�.�HrR�r�[��Ԓu1ڵY,+S�BƆt5{����-*Z�1�e˥Yp��إ��뼔�LLZ��zC�������e	&�5��c�.���8Ym\�t)�ǲe�
�dO36�^�����ۛN�3HS�@�Ư%�b�;�	�o(B"h=!��7�5wy�=��-�)`�֢�tJL�f�
�'�v�-\���];=�ѣ2�ߤ���<��,a�XH��P�w,P�׎�wl����^Ħ<;@%���a`�H8��^�w&�J��$�5ֽTۥff�cLp��u�@Y��*�إ�m7�*��B�(��z&���z�\���R�ѽ�����O7��S)�{�YE���V����q�h�j]ݙe�����bNU�<���Ж�P�K{>��;�Qd�QIb�[���N�s�+.h�lS0,��v���YT����;hT�(.�B��ߖ�{J� T�w�Zs"l�q��v�+�ܷ���*+��oAr�&���x�jI�Ů�=�cU;�uh��6��!M�
�Vt��yX6%�)� ҪI�6�����ڐ���ckUұj�1��0dv�n�ة-ɂ��N�9un������,�2 �$冚ͽO]is���HX�1��2 �j���)!�N�f���E�B�{�jp- C.&���Ԓ�n�2S�ʫ:QZ�x3	�Q��\�r��!]�Ӗs5��ԁ	����w�����c,'w��b��"h�-&�Z�6�K��M����f&"�F=�0Ve�S: �,V�K�y�-�r�B���|�*^�Yj���-�t�B�eV\���ZF�Wq�tb֓�{�x�Nq\����͵�
_
qօX(��P%텷z���6jܚF�ò�fCZK[7Y&�J�3�%-d7��� d���,6�qRR�n��Z2��$��D8Z��8 ���$8ol<�1m�ȅ���cTX�V0V��QP-Sܗ{��o4!���G�E�F�),'�m�.K&�@;V�Q�0�cSڲ�X��2�-<s���%Q�־�8D�t��Sc�5�V�,��6w�j��p� rm�V�M,{�\sCZ=L�o�̡d^���6C\�c4�)V*��z�+^�Al�n'@k�0
��i��v�چ�'xe��ݳw��fDYgk\�R�n�c9�9|yX Eݷh�w�J'W�VK#� ��'dw��ǖ���j����M���G*��8�rU�O���t!Q�f.���;v>#^B����V�`��=�e�������j@�ى^�엻��q�č^�E7�&Tͻ�D�m�k1
�2ab�5�o3�{v��Vr�Ì��"Y�T2f'x����C.��f4�AF��o�?, �dWO1;�>TA7B9�� uX�����؎�Yu� #X5f6��Z+e���v%��X���>N���y��f�,�Mĭ�H���E)�A;���M�6�LG��K
�i������0��ͺ��U�e�I���
onC�)�5�{�7�(1WL-����۵�"�&C�U����2�Z]����Q��0�L ��D������X���j���o-�_M�l�íX㵴���3 iU;R�֐8�Z{Z()�hV@�d�L�HX���#i�Q[�HK�ѷr��\��5�,�r�M�t\z�,���͓h�"�����"wDTh��� Ж�C��X���5|a/*l�*�< k���*(��M��%�����s�f9��<�+R��b�����|EJnXgD��@� ���̈́��*cl"-XD���;Ŵe���Vv� ��C-���DQƾ��Aۈ�b򴰦�n�ڑ�YN �5	HɈ���f�.�/IT��w.�1�(T�R�$W�`�+��i \����PKQ�T���8�yf���t�2�"�b6�^�2���2"�㣰�r`��ݛJSv��M-��HFŝ"kw�N��D3Y�W.�v�JѬ[��2�e�#y0�,;�FjBėNb2�2�K����p���)9a(-I�a���GF�yF��D�sA3�W+m��NБ:�b/I#]��,ڍ�K�Z↶��ZqX�%.�d��[F��V+��i�� �2�VTR;Ov�I*Kko�&�ȶ^�s�[�j�%J�ۋj�F��3&!��\Ur���HSݠvʹ�T�s�wZ",VU.�g2�e�ZkrQ�ee�д�I��ۢ�u<X�8!�,�HM�b]HA�R���K��"���ndJ��l�&ᣂ��+���$#��ۼ315uB���������m��hlE�i�^��
�7�m
f�\ڊ�"YE�V��p�y�"(:i;!
�3l۽�j��+Af�T�C����6��ӦU4�C�����f0~��k�QS0�RJ��	(	� I-���{���l'q�uvй-fmX�;��[�iS��s�����LV�ab�5
"������q�OF-4)��'Z`���d8fi+���Ƶ��W&�enJ�8.ʆT@ժf�������o��j0� ��wb�u���47t�P���S����i��5fm�Ww��R*��5�0+�a�KzU�2��kR���ڡw4���k&��[-����l��k�wW��Ϊ����մ�%�Q�_5GC�!Զ��"��I��Vk��� ո~ NIwVJ�i�/vY0غ�n����v���io.�oD�������`��t�E�VC�Q;���T���86�H�4&2���2��zR�֭��V*�`�t[C\�v���������
�K!P
Ě�L�+5�-��^��T�\�G�Gt<i|���FR�,���I�DF�����),�Y 9zV)��h�{O [.���xe���tQi�i�Ô7��.Һ�/uJ ��b�g��Į�`ںY�z⽪z&¾��Ҍ���b�l�/]�	I�~7sp�sC[�J̭��v#dk�TmZr�;A,cCGj����4
�+�㹶 r�
���u1�TQ���`ֆ��v����U.,X��-*�8j:�
�D���{�C̢JKF���#�qR$FR.�����
4��eD��0m�#�vD퀤1^,One��^������f�Ҽ�E�#Gp���*9쬽u��z� �`'At½Z^�r����"�B{n��N^�� ��B���F�)f��KkhH#�)�ca�R�3�hn4Ƥo�QpVEѡ58�Z�RYVZt���	K F�W���=�H�����{��v��,*=I�sX�i����
� f�llB�7�:�U��w��jג-��XE(%�'^��^�Xq�4�#H����ܚ�V����So
��!�pR�gp�����f�1}3F��d��&ۇ 5x��7v�5�4�jȨ^=a�rں�w�h�.�ӣ�mb��p�z�T���d�S1Qv�ۏ4=TL�x�pV���a6��[.]��:G�J|�7����|� %ab�(�w��6�ئ��2Z��R]S�e��ԣ�. �U�In�)r��d{�)�m�uj��[��,x�
��X�ke�L

��nylGp���;8q�w��FhpP�9/we;y�'kH�����ͦi��yH�!�S�Օ�lʊ�`���իG2�$S�-Fjb��tun��r���IdZ,TJ�\JFp�r�eK�&!�ܫ�>Lֲ콚o^?����1͎\�w�vڈ
��Җ1��\�hܪ:�l˖�Z�	��z�7����#6�V7xn6*�jʱ��堤���1in[i�]4�P�:��ZDE�	=F��MV��Հ;�켱[�R�4
*��r��(\)��٦��0���b����{�����Y�C�NA#����sw{��r���6��@�4�"��:䷕j�_M�IiV�*��G�_-yQ��b��X�kh�m��U����OԺ&c�\M\��,�C��֙��י�V��
{��\b5���v�%"���vطu�/6$cV��Ͱ@��f�t2�E�T�-�,�Nd/,��.��+��Z���V4��鵷�(���f�bb�I7C)k"T�&�{�j�+"�;HY;)������-vN�]�{2�1�`�U���WgU��År5��7�X��!���[6���#f>qp�J,�Y��Y���l����ţo�gK=b�N�#���O�!ն���E��>���ص�R<�8�����1f���J�c�����Z8=�֮+�l]�G"�Y�&C�u�;����0WAz@:�; �K��`��jw��%�]=_y`݋yN�kl��� �XRڒ�{�&�y���aȺ�^��po�w8���M��q��R��[�s�����+��#
�ǟT�+�r.%+������8+�tr$�Xl�FjFh���d��-��u�1��{;$���kq6����O(����Q��j޸'MW�M�2��2�}l�9(�zz,It��{zl.*����|b��.�R11ƶ�������[ˤ��o�D�˺��l���l�]	c�K�+��c���!��,�����p��N��ٱlk;DeW&�et���.3�o��g7ćK �+�h8DmL����q��ynf�~���j{K@I�������9���EY�=}ˠE�B
d�T����$[��f�9蕫o���wHbGv�k	7�c|31�:��:����=�6�\������r�u*.�t��[�v+`���)ŷ��7u��&��w����@�2�,ۅ*l	��s\�`;�]ʰ�F�����JXF.f�Y�ή�%iຑ�	Mt�M��WV*�B5�N8�#�b�����֯�p(ۗh��#��qI�7��u����Œ����� k
,�G7�z<H
V�]ݖx�]��zt@����=��Y���5�x��O3�.��sD��SR.�yۻ;��f=����*P�ɏQ�$�VP�R�,��� �@����7�ƅ��Wg�����zέ-
L��k{bE_$����Ӄ�=J�d{%��
mk߻�;V��ҡ���_|�T�9h�TZ��l80�5;i�Ϧ��a���ril'Zfe^F�#ޥۘ3@��Y��i67}�)|1�c�6���kEu�$����.�)�����
<�r]&�L��S������S�U�:78H���ܷ��t5u�6�Jq3w����G+��������lɕx1Y���3 ��	._��x<�JN�%]��onVU֨2-A����E�]�v���� *�.��NB�U�I��݁���&n��Պ:�y�>Ӛ��OkM<�,F�¯>r�^@��p5,^z`hf�ɮa�%[�=u���#��y[T,��8�R�[�n^�q��Y�Whf�z�ۄGe���w20�O�GW������KXk�<#{�4$����w�M�F������+���˻�sh<m��ʌ�M����VO���{�*4���;o(@rx�!×i�w�k�sI��F�@��ެ#���7�]�m��]z��݄�of���.�� *�ר�u֧��\�;d1�S{okfG\�+��m��R�ͺ_: �$�wm\�M��K����s+��89�q�ܹxE����N��I�K�x�̱F�Q�M�3�'�\��=�[�܆��YAEL���i�R�2u@w�����e�ȹ��)���x�6����/6��su�J]]��c���6�Y�x�� eL��[���%]IӘE�����e�ovgRS.��S�7Qy�cd��Λ�u��t{`�3"ƶ�V�S�wy�����Q�4���K��ވ���4j��wca��kOTwz��9�"\k..ٻo:��l�L�4L��uHt�sY�*�u����S[�6�K{�򼐒:�]��* eN��Z�S*�y3��"�W�ɸ��#�An;O;�.�4��*p��,�:�zd:�Lx��cz�II�$T�
�ܵ)w�E�0-w�ف�(Jђ��v�igD��Y���n�}�oU�9[���j7�JG�MypR�l_г��ӷ��`�9��㙰ԼwO�%��N��}hD�f�/�����M��/�%-ܥ�6dP�ڸ��=p�!�Q̮���:��\��� J�I@��ek��4�[tH�'x6�v���]��9ݻ�6'�(���f���ܝ�q�"K[�;�D��ڢ�Vm�u<^o����\�2N���Ģ$��E�سNfn�!�V��*�
���irڊu��^DR]G
�vi���|���{Jrv;���H�7:� �+7[�r6��M��@ݚ[�V���U��f�<J�U*�3!]��n����)����|�sS{��]X�)R��[{�\L�:��:�m�+'��L%�QЮ�ؾ�	����i�-20F�&Qu�\����Tz%��y��G A�p[�xeqn�2����iw+�5ڠ�!J^��zb�����0#"�$��ة�R�+y�G`���^+�!���@ή�\��l��������XJ���2����b5��S��)@Ms��F� �ib�F��AI�v�������^���a��w=aZX����1u�;���ti��ݛC�"Q�8�Z���*��I�]��ճ1���vtaj�r�1�������cKE5wU]��Gs,Lov��ԝ*o���.�re��1A|]�HIxzRWf:��*w�U�J*V�)�s�iGl*q��a��l6x����%���X���2^�j*�Evޑ:Z�5',��`�y[[-�5i|��Zj�=K�������˕;V��ԧr��H�p�r�Ge�pbH���B�Z�>s��[OLͪł���Hf�޸A�f盬esldȮ�\{i��P>ܧT�QP����:��cHil�Sej�ٻv�;���^cH��%��8M�-���!^l-j̡��;�<��a���W�:VM�:B���-����݃k5һ:��x�j|���Х�c�mWu]�F\P��[��t��|7v\��x�#�|	�[�þ]b�0C%�=<�MK��6��9�}u�j]	���J�܋��j�֋4!ys"�M$�Ə�Qnvi��2䨷���6%g�Û��\��I�f�p;�"g�.�μ��6��ں\Bb]t�*�!�t�/�]���F5A�{M�e�]Ku�Y��K�d�����Q�3��)V����r����~Я.|�ݣ�cS�**�;�ըM�e\|O',V8�9�$X��[HL���:��{�7VYqu���[�hTz��yw�2�tRN[�Z]�:9wYXx�{yU�{�ܔpnEkG�!���r7h�{��]�fGF��ȩ:���YɇiLns�L����J5ڲ�\-LU��N;�/a��u)F�4���6$5��uiocֻr�>�](hsѻ�u���TX�Ruۇ�L���VV����:��v��\yR,����V�0јvð�:�5X�4A�v�jd�y���PC8xv�1)�N��s�澝�u�Mn�ܾn�#f9�]�Z��V"о��x�wec%_��Ђ$q�艹��7*5J��١�p Z�|m���S�;�n�%�p.S�F�ɋ�"M^:�s�^س�H�(jS^�'��c~��ݸ��u/�tt9ݲzY9X9���K�#KW'��#�w&�|I7��ti`{��Lc5�=���K��u��xntɻ�C���j��w[`J�ʲ:��ɠs	|Y�����@e9[��"p�,Q�D�� �5��ۙ����k��ʗ����A���Y\17y�23Y-�l�:"Y��0�|�2��t����0��b�l3��#yŉ�i7���X��GE���*��ٓD[�U��n!1�U�����mw*2n,����2h����S��جN�D���
0���u�5wY|��7o-+��]�4�zm���N��My�lॖ΀����	��1JS��H�Loo,��BG������C0Ds�nP�ܠRnR\��^,�S�^)`���*��U�8Ժچ��:��_P�Gk�Q�zd�Y�An��B:��1���r��9��v��c�I��k@��ɚV�[��u�#�a$������5��6/y�����]N�����Z؋����|�KU���9
o�Uii�k%v�2��s��z�P��M���92����z9S<��::�Z�9��_XYi��j}�w��ty�xu�z8pK�7o�lb�����2�E�����3ΰi-޶��ۦ�q�x��o���b�-c9b���JU�5��) pN뙏����/�kz�P��ӕ���х��6ĩ�ۦ�ڇ��I^��[G1�G���<t�&]����=?j�zK��s���5;1����pP�J�=D˗!2�;�3���������S[��>͠E�=���m��ʍ
z������{]a��h�yH� Bw˴�MXDe��7���7�;�p���@�R�{Xk�/w���b��!��r�K��,_]��t�K�)V.�b1e�hۡeܝ
/�y������\�HA�Qr��m�&�h $�����ۍt���of�1X�X��SD}GԹ�p�w�C0�O,���Q��Pޒ�5�ĵ �7�<�s���7�Q�&)YB�(�L�
�#C�>KO�Χ��s��I^S6'���'���]πk�1�R9ӕ2�&^fu�u�� &$z�3{��b�a�;�ǻ)Z&a�3�̧����|^����(W+�ҭ�A�t���E�O)��<�fք��X�r�<��f��um�}V�j�(V�s���8�J���,ۍXu+q��)��x�E�7u��-v�@�m���ں]�y��,@�n�]HZ5k��k�\ңP�v!|��[+o�N	�a��]�S�w6��rx��9�T�[�� P ��}6���ݼr�acy�[¯1���Z�e�Y��ѤŨk�F�p��>��M���W؋9��n�����[�M�h0H؝ 7��Q!7����\F�#'7p�<֑��5j|7h9��ݥ�c炮Pf�8F��i鬞���HT�o��`O�Q��p�\���|��*�<sA`U�Hu���]�1�	-��<X�ˤ�^v�>�M�@����B��;�jwuNw��\���m�F���7F�k!rT�}}7̋1�m�������37�t�{��U���]V��{t�q��č+6���E�Ž�Z�<u�~�Uy~�j���Wv�p8]�$���FwWv�k���(�m��nE��<��O"�]������!��8�k.`�Rm��q���"���|H@H���d핋:�H^��l�:���̓i�HfD�k#�X��Kqv��1t3�*{��N���l=7���^����^�X�!9��'ϙݜsD�e�Jmor�Hj����ۭ�)aw9B�Nx񅕼2����6�"�_+�7�`8�7�a����J�c��}��2�V#Z�r��+t:�g]Ne�*�C��v[���)���Ãw��M�C+i_&l^u�q|��2�%�Z���4��wwv�[X�:V|RH����,�7�gsB�t�D�����^�e]���|Δ{�z�s9C�U��X��M!Pʂ���xݠ�A��hVj�3bKN��R��>�Oq��;��, r���]^lH����ÝE�A�Xi���p�������)]J6�T�G����Ӧ���u��Yd̍ԛ�j��'M�>��9Gst�+��U�S��R�{�Y��f�HV�%bË�!`�ڵ�Y.� 0rW ��P.�F�҃WZص��ݣ|�9��;�גF����Y�Jh*�����n�����Le�ڄ��>FEY4��8p���/�u��K.!%�CY9n�<�u���Vv��X�:��6JV�E�"hG��iK�y�7���jWY�.�P��Cr0/:\��V��Zt��}�n�����j=�4qܤ�E��U�*����rP�pVv�\.��3�a���Z����/[:`�A�ж���m���#}GnZ�_}����z�c*l\8<.m�n�s����x�j=��X���<�\s�Aj�����;t���/���c�ɚ��m�[��E˫�s��*�
�x{��to^lb��|�W3�uYj�z^�]�
.lU#&���3;�Dt�&Wt��\x��E@��%[t��YWV��l��!��������m\�4�C��r�o3h����k.�GӺη��r�)���'����E�����1��N���CL���%X��ao+38���x`zԚ/e_W�Q�J�R쭮v�i5	�I�=/��S&�>[Q/���ep���T����4����T��H3n�mH�����!��Ȗ��W�qa�pG�s��@WŜ��d�0�-��h��K�Ŝw��{wQ��|��ۙ�X]*I���V��z��o!Yq�9{i��Υ�H�8�Jl�f� .�sy'L�mi����.���0���6�$D4�<2�� �[V\u��j5Vo9�>�kM�;}��$Q�:��ls�Bz3�G��]��u�L��h����[�ŗ����c#(��;p�X��$��P�0�.+o��I��<x���J�,8�o�^���^���	H�W���^�:�̶�ub:��i�:�?c��%���C,�ֻ{ON��L����Z�z�ö�[ت���%^'O�+�պ<�P���ݡ�O��8��ksqr	��G&3�l��:�����'Q�&��́�b����uK9�-�3���ru-�\#�r���n��Q+(A�uDS�P��;�u�D�D0[���i��� �.VAʢ��Q�^ID�9Y8)�<�l���L/f;�KE����WZ�e��@�X���7�l�|�Ռ�������c�I�]q>�57C���AX����4`n��e�B�3�bc5����b+ojb1�&���0f=ή&�u+��2'_���,\�is`r��jf�Wjٝ۱�4vt�TNW)���+��\f-u37��:=���_o+3�m��ms���y��ajN�4��c˜K�����ﾏ����D}G���L�<�Y�/+,�{�&��8WV=�NtZZU�H��9ٗX�V��5��W'M�P���Ý� �yҜI�!�]s3	3�V�u/Vaڶ�!J��#6�04؎��ݟ����6�Z�hh�}WW�ؾ:�mKįE5��uXK�@��r�qe�X�c���� ��G�N� \��'#0n^�gs��Sz�T���n�]�.�ӿZ�7N�,��:�7]��A�x)'�m��g6����Z�N�y��dsx#�|{,a��� Ȱsz^rWus���s1��|�C9���r�s�R\�Y0,z-��v�3�����3ivU�%�O��f��7�s����N�3���|�S���wL��`eu�}�����!�������S+0f��Lވcl�c��q>ms��]�=����,���4.���T��{h�V2��@�z�Jk0�x�C�����!��/qf0o�
WS!�������C-걛r5�z��2}*���J	��^�R� �\�Y7���b�щ�l`]�k�g��M�K��}��$��5wfo%4{a��;����iG	��V.�n�Mh#���c|fL��טQ�����67�֍����-���m�=y�1J!�`��l��y9�>�F-4�M�,��m�es���m�̡{�n�(Jᖛ��Zhݱ��2�d뫽�i����n�{��C\�v�_pM��V=�4wr�%wT.V�[Ϭ<���`Z��ՌE�H�l͛�=�K�T��u!�iwwF�PΠ(1������Z����Vh�ДP�u�Q�wd3�(I\6��#f���6��q-@�ǣ8��HP�O�;]�`��z�B�جi)>v�^d5l��]�x�J�����)�ݬf��V�K�2:����Pvo;o;m�p�(�t����-�.�ںcdF���vfMN�:l+���hu�Z�q�2,̓�R�j���]�9����̭`Rk��j�Zw���0sWk2F��g�*$��ܮ:̎�y�+N��l�Y�{�|U�'�u<9Օqǆ�|Ӵq���p�ݭݬQ+t��xQ�D�49&tSGE6��OR*��$��Yj�fd���������AcQ��i|�Q-��ʞ!#6�k���T��^�f�N���$�i��XV�;���ՋM�K��Ԯ��^u�ڕD^����]X[�4��@uq_'ǥ�u�Z����p�za�kN������M7919��X{�W�A@�ۻ�7J+���б��b�_D�1��ڮ�|%$�xr�Ǡ��Y������n���;�;_
0tyr��6����w+
���	;�Y:�}��c����\w��R������hLG>c���:���]]!�A^��36�7DTj���{�+TtTǎg+[}X8���M���kl��G��1N;hS����ڭ�}û.���ʆ�7K(�M`�ոڊN���p�ɸ��{YQ��o(���5�Xj�'6�_Z�z�oe݀�L��t�F����0p4��š��U��7"���,�h8���]��7	AA4��97DY�n�ֻE���+y�7�,����*=3��`ʀ��+;VDo�o�l�z��[���XډaײSq��wJ��%��uw+I��c���е�4��)�ކ��=+6����m�R�����J�鄅y6��3�_u$�S.�9��Y�MV�0P'R]d�c��Ю��F�A�j9�{RZ*Zν�Nk1��"�kF�T�_X��V�1�E�
Xl��&��-�w�M��U��լ�ڎ�',�� x��1)ʈ�i�y��d���ŬulW}���+z^�Mb��Gnwp�����ܢ
,�5�����Q2ʘ�ϖ��E#�����ϫ��R�-|.��X'D���Β�q�h�
�3��ȺiN�G������E�aS��Pu�w��-�9=4��"��qsF�Va���$��|�)#޳��Zh�vNSR�T��J�?,}ܑ��Mmp����rmu�yє,���GVtk�ar�$8�̽��Z�48f֡H�A�Al���<�Q�s��)Ulf�u�4f%�uC�*\В�ilޭ�.���T� �E��x�[OR�IRN��\�eYڴ�C;h�ڵh�+^�26k����N��[yF��L��ɣ�W��H*���]��1����
݋1R�Ox���g�����a�=uYmQ��³v������ˤ�{�����:�����{;�U�`�R�|��,mB7qEk�e����.����&p���5�V��AMխ3tU��.�D�]z�	.��p�ۭPӒj�j�J�YCsz�Ǚ�Ƶ��
�{�{��"�[3�v�3B����K�5%����d���ʂ֤�+��[$��]=<��Z0V�\b����qV�)+ۻ{��
ݝ��9Вg�y��V29+r�-�	��v�a[`R�Z���X�Sc��:�n�n��W׋�ї���+/E,	c�{�1�P�ץ7�:÷�
���\ݕ���s��[:��ӷ�wv<��(�g��_P��C5���b�R���W�y]��ח��4+\��ОK��z8T�Hk�u���]\Ua��;����,�LS1-���eMUF�|K�J��˻�ŧ��2[�`����� ���B>�����]�y-�-��٬R�;Er���)��.��6�{�wƴӕ��F�efdz�u(h��έ�l�I;�m�:�Y��ކ>'�{�t�]�hA�vt���&�����{ݖ�.�`�)�R<�v�pCv�ƫ6��M������i�����Z����wIM�Ѳrj|���ݍ*��'<����`�X�#ĉȷ\�v�	�;�Z�8�0�o�6��i��;5u�1/GYÖ���mܔ�Ug�Y[Ζ���u.��V<�Q:�Zz7���^ݠ9���hT�fV��5�D.��-R�o��c��.J
����oGt6q����)HwK.q#U鉷c8��n��ԭ9��3^;��"��C�+[�n
�'�cA�5[ 7���J��h��o�s�����gtK���9�P<���k����ܰoj:E�ط�2!"�_Dke]^��cS>�n�������l7e����)�%4X٭���2�w2��_ˤ53��5{B`�:�wf��+F1Z����<�����6�\���Ye��9��4�m���m��vm��kr �oE��v8��_,�0,^ͱ��2�Ff�(D7����w��B����U���Sb�_=yN���k��Ѿb�Nغ��.����z�M$�M3m���F����\)��gdP�c� >KMBs)�6�ˆ��K#���
�4PȦ���hhMcPnS�sM�Pa;F�|0��aqN�Z�p�݁P7{[��Gdɡ"RݵI%��)-��Y�*w�(�u�N+j젝6�kMp��º.;�ܴv���csdF�3;�]���b�`w���TE_%���,��(Rݼ��E3�hYr�q���Z�D����2��|ҭ�Nr�F�_e{�s5��OV_=�@VU���N$پ��R(�=��c���/�]]GE�8���i^[�)\��'����Qr:ZY���2[�7!y�XN;V�Y�I��(��5�a�o?���
Wn�bw����nP�7�cU�ru�Y�c�u�\�����>�j��:U��K$�k!J�`���Y<�Z7�r��R����P�긱���e����8N��lǴ��E��qv=᛽dg�El�8�ك���
�=g�*�S��C�t��{�ηЩ�_]���n�. ��ܮd�T9�v���5��y�l=D[���K{ZOb#h T5��]A�C�ty2Z�������E����:���v�"��Ў�nIF�T�k������R�S{�ᬫ�1[h5�߮صQ,U��h;RV��:��Z��Ż�l��͹n��IJĵܩ�Lv���FQv7&�JU%�J��G���8��l�#��V�]Jʼ��l�{Y�˟5f`���+o(�VN���m��g
笟�[��t]2�ވg`���em��{`KT�\h�7ك��S^eڠl�!�y�\��5G`��x��.���g��Ƕf5fE6��ZU�/��͚��'��Õ�ܰ��/b�qu�v�_t�K�fN����F��RAh,Z��>@������%Aݍ_ں��T���c�c{8uKٝ[af�^�ڦ�&��y5��!���Z_WfC,�����n�6�`�QnD>#���w���G;�e��u+TE��`Z��t�,Ԡ@�w�;�#G.gq������ZѤP�Y���hb$4iQ1w}jNn+�!8��|���h��p�L��`8�#W�u\8�We��{LZɤXLm���jw֗5�^�'�	gcd;{R�<k�k/���,Ec����<Ni�j���	pF�	�f��yy�i�W���]-�R���`VRœ��,�����5������)	�"n�)�8l5��f�hD��C۵ik�U�uyMۢ�56�);W|����RamY�E4V[��GJ�\�f�w���G(Vf���aJ���ĕRƈ���t�����QT��:�p��`Ա�ޝ7���zEf�� Q``��K���"h�VӰ��@�)R4nt�2V���bhY]r���u�˫����m��Y)�2�����⁠�Bo�BHv��]X�
�4�P�O�b��R��+�`wjge͉k0%wC���t.�]�:tY9ѱKu�b�pIs��"��e���<�����u�-��9|���aPT
��k��-�+�x10��������G'��p�7x깴h��-�,c�U�;f׆�	e��4����A_:�0v�����g�7V�$.io�L�,��b�X��NQ�Ͳi"��`Gy%6��yG*����b�0M�Ѭ�t�'c�6����lc�m^k=�������5�w���k.g`��AZS�s��a�\ڝ���`^wR�.�aˤ��׉��h����q����:ŸԘ����n;�(ΐ-e�'7y�����jp��9G|����B�6�S���.��ai.WI���R�g�i��F��^A���qu8�*��1��H��gd5�7�F��m��4�w�����Ns͙�w�YGo*�DlM+$B;{k@9Z��nf$j$"���؋b�w���e^%tNN�	���F3W��;�As5�ևX=�Q���v�"b]�����L��X�
8�CW.���U�&�൮]���o@�=+tXm�=D(mhYq���4�G=B�I��c{/�*�m����\"R`j��Jd�1�n3'9luI���j����CaR� Z�}y2��p�B�[��u��S�-�rriܭJ�0�#i���
3�ͮ9;`�oztY©�ԷLajET���Wg]D*���ă�U�K�ʔ�'��:��oL�GmJa<��9r@!��D/D��ܫ�ޓ�0ں�e'�,-�H��{�r�+s"�p4&�%;9�%_£���Imvn�]̉,T�����z��J'��S�5�λF�؁dܨ�/ ���x�Cæ,̝��0S�����z,�����*D�X��+:fʸ�=���"w�Z�l�	u��]��E��>�du�uYPA#Z�u�2f\�x�5�NZ�9�֎��8P ԝe#Gh��wK�4k,��9ힾ�����*w/D�欬gyA�%Ϲn}@����y�;�s�/
�CB���O�ݹ���I��^}z]-"�/L�l.*]�s�t�f(]*�W�6%�U���2�c�׷ܝ�5��6�[�������g'=�E ���XhK �k'%C�N�chG����f�����E+}nK7�+���؄�c[-cCN�հ]d�-�ΰhm�w�,FF�&(u��g]<��D.�}���!�v�rp2�	��&��ۡL���k^�] �cw��ڢ�_dKm-ğ_L-v����t�5�2��cRwk�9(&ٲ�T[F��� ���/����on����iw�aZ�7�F�*��.do�(K��`|r�j�p�6��&����m�������y�R��F�\�5en���z��mY۩|��:�&�cE��I���Fҷ�*ct�+�N��egCh�jm�w\Y2��־,��zov�k�C�w��hT�[y�Lp�2Rm��c$%v)�Ƅ�ods���Y����ꎅ�ݵ���7t��'c6J��法s��t�mif�%޹yַ�3����YN���Y���-�w�1�t�ƚU���ɓ�sLΈ�`S�i��ұ�3[�J�)1򥅅	�%�d)8샻����x(<
�îY�C����!��� U��03^ء�V�mv����w��d���E⭙�^��;�� ���v�n>K��nr飴Յ��t���턀�{��t�:U��:�g"۰�۷j��WXU�Z�H*�I��H�B��mڦE�k]𠱸m�ٗR���ʇ;�ɑB�h:��h�n;z�V�WoS5[ո���5r������Ԃ���)]ݻ������v�I�b0LEM����Ѯ-�wS4�������O�hݢ�z�i�ݾO3��9SP���ս��V��B]v�*��p幗�����Jt�u�����]v.�p�!Ty%^�wʙY���`��NS�y�U˴��b�P�V�
ʄ��ڠ8x3#U�閝fZP�܇�QV<� �:���R���ﮮ�[�XX�:�{3���5{)A�t�qGyt�}bc�:��mZ��.
���5�[ň;)5����8�]�v�>cE��.�ڠJZ�U�n��D�w�ak��w��K�pT߅����{X뙜������!��,�ۧgE�z�S���Cձm���Qx.��l���Z�ӻ�k&����
��[��/����������t��WQ*]���d���v��ؚ�,�k�ʵ�[��٫�ˣ��i���a��+�fw_;�6e�@[��/3�;�Z����Y`��0P}����JԅK���i�Sq1f��۶�ׂ����3�ٰTH����c������6�إ�ҥ+��8�[��l��k3��T�ZM(~��9r�*�[��`�r��v�r���QG��d6�����gV\�c�l�j�b�T��\M�p�8S�o���N�<��o��tW3�*:���+C�stV�{Rv���SRl^�cN�v���,��B�Ұ,��rg@9Rs��ܺ���bbN���2�?f�νĴ>�j[]NmsNhB�E'Y�KfUNq��v/�27��'+ó��Y�����n�`�iw����$�2Rۦ-��,-i���Ѣ8��J��k��v
Vɉ�õؙ�b7z�0�m��ۖ�98y27-�����4�/M���cZ�l]���j놌��������u���/�1�"��+����{Ê=]��Sv�;��J7u��y��`^*y�v�>{+��9��a1�(����&�S�y2u��r!z�:7S!�Vd����V��B��2h*r˃#���tȶQ6-r���m\���,���(�P��wt�bk�=�?��V������I`i��$�v�c.'\�b)�,WOn���Ňpf���D�Mr�£�Ü��EE\��$��d]!	9�*��#�N\HMYʜ`r�Z�(�eE���d˅B�PT�Q�]2�啇#�DDU�9¤�K��eRX�ETeN'	'p�<�j@d����ʪ��\�0@�1J8TQ4B��.RI�
����ӁUQTPS)�QDU˙%4�\�(�W +$�QfQHdr�G+�ͭ&Qh��$M.E�B.Y�ʂ��s�"ȍIU�����(�
��3�]�����Yȣ���E2�"+�U��r��U�EJЊ��eI˅*:I�eD�
)!�(�*��QW5#��(��MŉA�!&TR�ˇ�rT�Ȣe�UT�.D�&D] ��ͻ���޻�����akSi�΢���7w�aYW�"x�+�5�%�淼{}C3dL��&��w�J��Z�hR���z��{�8�vlH�/�@�.�M[�ٱ\.�[��8�uָ?��@U�3�fr���vx����@��`?�5�%\7a_p60�¼w�;e�� �{� )2{�gK{Q����K��7�@v�R�v*�����V
C�8��g�ڵ�f�����J�2���s�u��<��Oe[�e
1k�΋!��KS腓�-H�.;d+�(v(|�by9���WՋ��1ζ&��DW���{�>�F���X��S�y5yu-�G�j7�~�O��p��\��A�3~*����(uS~���hn�vW������h�]��{(�ºĒ�=-]I�����Y&�o!� Nϱ��N������ޚ+ʑ��q񡲭��3��8�\._������r�Hw{=D�ef{ :2X���F��ٛ��1���h�\����M���{=r�9�j�l�g�6��"�b(f��S�!�M�Kn��<8.����p-�Љ���e�N{�����W3�;~D.;�>`VJJ �i�tL]��U<�7t,����w.���	�o\=�wQ�-�ur��ƞ;T�W&���%��/T/%.(H�6�́�֩��.��˺������[돻�X=���{Y�и��EwP�w;X�9������nh�v�ݞ��r��.r1l�s�5��2���3��j�{yg����0s�S���8�ѷC��sn��9(���f�)ד������^DpBi�=O���\)?+����5��2� �oQs�a�mi����t�7w�����6z�C�.�>�0�]�6h��S�f�L33
/m
����H�^�����O$��J�XT)�Q���.V�2fR���۶+���b���uRT���Y�F%6�bW��DG�G�PG����>�p9Ya˜�W�W/�1��u�|+�U��k�8��D��� OGD��i�J>�y�F��؜������Ng`�������1�]ć|��Pn|�x+��u��?#��Ѫё7]m��,K�|����꣹�a3[
��t�@p�o^L����ж��H�ϯ��U����#"1X�h�tE8�{��Qb�R��EvkҭW����S�������>ԯ�x׉��y���z��Y;�������
���*s����������{��| T#���[��������K���kN�%5�8YSW���"�Y��/,�\"˾P�y���]#6���u��f�
�_ǫ7+vӝuژz�m̙�,��F��7#LR9̫�ds	3{�0�k�+*�5�Q�Z�8�L�b��e�[eG��:�Tد5��b�A�!y6������H?�����5<��C����+=�1T����ʓq����8^�b��zz�������j�`~�hf�<x���ҭ,�{c<�vFa軵�G'�U3Q��"���s��~��ٿ6V{��R�+��m���ph�����u�7xZa��j���}+�aq�����
}$�\.���<���q!E�a�|%+/�յi��[�כ�*k�@u<��ĸs#mQ�z�,K��=�W�У)����Y'����#�<�!y����8kت�"�P?.���|y���Н�%u�C�%
pO�jzM���*2�)�d���pN��$���^Ƣ?EG����A��pߨɿ9y{}wS[6����\���P�g���9��	]���@�;�r4����jP�fˆ۾��g�97/e9W[��#`tBh��^���~�� O��x*4pv���׍��z6f>��}]ݤ0x��5xe{ygCuJ�ɎuYN���ĜUn�	Kiw$現u��3��ӌWB�EO�,��9ʌSg��;.Xj���F�y^[�'zԱ�N��Ց��뭊�����b�]�b2Gc��n����jz���xQ���mN��`:V���@��6b�V�37fm"�8�is�+w�ӝǸV!��{[2+֕��Ӎ�"�������Ήn�Ug�tC�C���_����g
�%8����d���:b]ݷ,��p����:ڛTVۃ��GM@pڨ����i��D���p�����VS�܋2�Ɉ�j*zB�q�f��������;�t%R���w�.w�q����Z�����by�@�N�"����n*�Dχx��a�saY���a��k!��%Q��ZT�����P$��Cuz� ���N{d���nL��#�mb޴�]Oy��+h�7�n��üp�Ʃ`n�k�t�5Pu��]�7iN��0�{;�0)��6�q�3F�ON�3_���@O}���*үW��P�;qDE�U���L��5�%H}��P�=u�i�W�Ӵ�Q��fGd�G\�ɒ�&\��P�s˩����(.���3 k���|4g��N�\!��R0o"���U�H�.%�|w��Fq����w\����Ҽ�(��������\��Y>�����! \�/\�T����]��I#vo0=��3F,Sh�མ�O\;�!�����W��˔�.o���VO�����vN������T�Zck��S�3{��_r}F��ޕ�}�ZE���bT�3�d�T�0���c|��|'X7\Օ�kM���tX2�ޤ�V���	��yj�h����a@s��?u�=xP��s��-�.|�����㜉�.��qW##���|��!s
��>1V�@A�;��))�
\����B2�$�����5�:d�tfq�3o��F��l�J�!��k�s �T�j-D�6��,��X.Q������tvF��_3��ω�5pu���	ژ�C��;;� �dV̈�d������Dv��Fb����<*����!�bc�N�4��[V���R :�������}2X�ʠ���ӧ�RU��%ԶG:�爼=����V,�1�22yoq��B^�7.��^� ��@{�|�ݏ��/��~G���+x[���e5M�\��S(����b�.j��i�}��K�a�[9�����988�٨�R���TW� �zF؟n%'8s��6��;ۤǬc[�x�^u�~�g ��[G���OrvG1�y�s��7�3�ٕ�mѸ;+��Cc���.��m(���"��� 5}�Y�H��aw�uZw����ng���΀t夳]_��G_�<5�/��f�œb*���j۴3j�+����
��m7k��-���7n���+�Y���ox�G�W^��\�h��- u�p�MK8��Y]"������Y�nK��!g]ޱ��+Xl{7�7捜�o�6+���`������`:�\3�ow&��5Px�8��vǗ�Ѽ�x���:����O�CW��oOz&���$�J�e���Ğqvx��֌�y��]o���Ν�����ۻ1�ׁ�  �GX��wEkm������"�T3=�)���hlt;Ts�孨�SaZ����"=��x����_6ƻ��j���.Tg�S����F��0@���^�9�������4��Ͱ�s'���j����Zj� �-���-@�&��<�ɇ��Π�g��|X���D�\:�&���S>���|�o�	f�zKu��˼�M��J:'LF���r̩Ms�@�3�v��!
�i{������)U
�؟��:�3)N�^q۴��.#_t�\�vW&�l�O=Ή[��~}S�:��:�ˋ�#�c��\�ħ;���7�,k4���Fw��i�>������3O���`l�z�<� ��;Mϔ|)�"&Woe��9�mNo���a��Odyf�f�s���J�t�K%z�=y&�'�~���oO��Mޫn�Do��J|��[���gm�[s��Q�o%u^�*�M�M*���%kMMZS�7�9��_r�}��K�����!��K��M]�yqE���f�S��乛���.���nOIbf:�Ňʝ����g�dC0��-m:��������PR�=r�w%�6�[�cle8ڛVxy�O	�|��{�����T�8,Z7:�����;k���}��vU����nx�U�B�2C���v&�W�Ov[�U.bà�x�Fz���=�3��8�)UM@`����b�I"����_���PA�6��|#�f���__Bb�Mk��N�Ӷ^0o�f^��v��#��y"6�V�\��䭖�͊��Sb�����3����
�k�o",z4���/�/gd�+��`u���a�5cG����}��t�_�f�����cS�֫,��m�ED��N{�\:7�r�g�d��f�Ox��Uj{��J
��5�_����j�J#������bjڝ�^GNE��\ǒ�+Hڳ��&.��,�{;�0mX��I0<�x��r�2��j�
0OS�����¸D&Z�Z��w33�刡�6�W65*����
�`9�=b�B����7�hY�_�3��2n�ܑI��٠.O�ֹL��'ف��n��\�ٛ��z�:�C���3$Y4p�d�f�_l��i���F9��
	y�r���{��N���\G=80J����8f�xGe��΄o!q:^ED���5�v����;lr=׃]�q"{�z�:���\�5�Ǵ�;��\ �>Ct�8W9zv�R2fy���sZxu��S�~EV��1)�b�b������%= N �@y��e튾;N��>]j`�������wXy5��ۡ�:��\g&/خ�H��$OB*v�]�	P��K��2����<�S�f�"��믚�5��+t0K6�q�M�	�����;����"��3����јs�}j�ɑ@_m����:"�F��w�a���&."��N���A�Js,�s�C�^�)��p�]yV�|����
������/��2��V7� ���OeQ�٠d��M�fP�qjW����Y�wl,m��k�A9�S�	˚T�1�.�w=:V�w�=�mq�*�}�y��8�3�ߩW��t9Hׅ��8��y��W��J���wfbw�y̪Ϗ�5�)��#S���k�ٲd���a�GF[E巻n�K	�[��K���@����Q6�L�؝nҜ�E`�ܙ�@�Sɚ��J-�OS�<���4�|r�ܣΛ�;ء�KsD4GZ�G
��2�h��c�kr草����=G#{�._z�A��YCP$����S������t�v �.��_5�v�!"�>�����.=�-W^u&�N��O�!u7�J���R�v]�/r��Txz��!S���w����d2�[d��C�<j+y��*�;!���O��i��k��gC�_���\�!��kǲ���$�������m��ݢ�}��2O�{�Z3~��ςq����`��鼪q�O*�n��0�������ܗ��T�>�n:0
�͛��D�W'�o+�l��UG٫Elh�W���1&��������A�88s��S�)�����|���X���[۫8'TġT�NcC���'���"�K��*+�Ĥs
�1mx�r�>��R�
J_
����;A�����Y䐎��=f��W��j�S���:=�{�����gab���ىc5��(���U�#v��$OCڥ ��<�+�#c��&�(�����=bJ��{��&z��x�(��D&�&,b��/��9���S�x'�k��\+7�x=�~d���:���Rx�u�9ȸ��� u:z %%�X?hr���y�/a���p�>��,ͱ��cz[O�tW���پ|�`�w��O2+�k>�
�L�X�^t��t�.�,ٹ��[}*󲺭�AQ�t�� ���x�V޺�3�����YmC��U�θC4'W['tã��syG�je):]�,oN������� 짉ٕ����9N��z���Gz[�wwU�;o�rR�ܧ/9-�;J�(&����*�~-�F_=���^�B_{��ۺ��V	�b���@��:�rl��z�����ٚ�bA����_�fz�P�"�h]l�Ta���,�Duͻ��+�%H��v7,�NrQ�6X�RS0p�U|�����+�=�`X����\U��N�����s4�/7v��P�{�ExGJ:���>XVlˀ�iDPB��X�{�!�v5.����d�.��T����پ�.�l䤾a�+n��CZ ���^���uL��Z�ܽ��U�9�r���DS깢��]��u��/��é�V�ɚ�2��S$����%�2�v���BU����y��]{ˆ	��J�@prPp:��zW{նʙ'B�[����i�ǘ21���q�J�gt��!�����xs��P6���CXJz^�gs��u����=Uk�C�����T�o�݂6�Ƀ�����
��b�l��F���Y�F�m%��7��4��V�����|y��[T��S��J���9g�U}���<���V=��v����k}�uጾ����'E����7`�����n�z��f�;�I�V���.mZ���q�Y����z4�XH��W�u���¦Ve\�.G"X��H.�� Ïq��.�Z���Ĝ�P�JC���Tv�A,�{��Һέ/w��em}m]�\�����Y*@�>�5�qq�O8��%�΂��_�#rM�!L���,��|xL�U��)�Y��M$�뎾k ���h���
��u^bʭ������)�D̄Ԯ�j�Wf�
T�B��T����#���O������:|7v��%Y����wZ�8�������re\s��[N��Λ{��S�X�6�+�V��Int�̷��u`T��&X�[8]���&Cu�@hܷ�;qmC���X:��Tڗ�L���]����r�٬Ŗ˩yW�Jw�zH��n���j�ewM�O+xڦp.���҅P¢��7��c5X�hs���J݃p�@��ld���%�^=`n�ʝ�4)B �k������W�ʄ�jB�(���\ Ldwh�����j�f,M#c�R�Mm*����&1G�{��+�(@m�K*G*��J�6-u�k_|��A��񩕆�f���k��0��u��އ�{E�a;��{���\�nqQt��Kw��i�e<��ެ�cg�޶�W�i�8�U��D'��x���yʺ���=-����y03�]Ӛ{��]�Q�oΕ��_}}�MW�ǖ�y�H��Wj�\�G �*�$��n��F�PI�J��s���(
d���'�NW!!�;��A�Z��#+�.�Y���+���.��\a��C��(�k�$�p��ǔ&Θ�=���,\���}����	V+.$���H�bŤ�Go�e��V��O��;��������*�`�V;T��v[�u��G�`w1t<K���s�R*�h<��flu�ك�ū$,Z��]����2�i^��O(����]�q�8vXƩ�B�]n����[���u�;�v�b�]Ĩ���p��i�yw|��-�'�^Lm��Qc#�7��lK;r�0D�K�e�c���4��ձ�IV����;}XPw�z#��T�u	D�<toZ��zȃ�����֦�c�v9-:8�&k��ݘ扩���oU��v�}��eh�Zb6w�<yeM!)��FQ9"gMY
�ŏ:bF"3���V5C(D^l ���{��+�NLtx6�#��+g��%*+�J�/fBIկc
��nt�D�X��b�ζ�}]�Y���;9VS����;2��4��U���)�F�:|&�-��Fg�=�B�,�/��@Q��cx�]F���Q���[&�YG��e�t��1�W��:/��;]8>��@2�!��˓��k��.��i���rθ�6eh��H��ˎ�nWA��Xbj�O2����h������Flz+���\�����\��1X���O����I\���SE<ۭ�������z:5e�[�$��T��Χ�<�����e�V`�WH���/q(�v�{2�W ��0;�s��={��Ͼ��	R5$��.�"�+�W���Qէ,���;�U�"��9�ͅTQG
�*)�Tʢ���\�Q��(��
���s�$U"P�(�Q�g)���8�rSs@��QqE�D�H��1���*PU
#�HQwW9�܈���N<�(�x2��J8�<VyEQɑ�]�#�y��7#�3�҉�A\��3l��A�;"\���H�(NEL"���vraA
.*&f�W*"��#���Q� �r��Q,�*����Uʢ�94���A""��\���Ҧ�ȫ�T��*�
�/@��'wf�F^b�	�K�k��y:�N�}q��Ү+qT��n��$>Z9�^u��2us8�iF!"�`e� w�]u�]�������˺L*�w�l��~���r>�C�{N��$��}G�x����!��7�$��=�=&�>���h���� ��SG��>�DCk0�:���]y��'j��\|�F�� ���{Bw�kמ����z�箱�Ǵ����ĝ�@�B����v�=!����ܾ��zq㽧{9DH��>����">� ����w%5����,S]ݵ2M�~� (dr. ���7�����o�I��o�^���J�;��@zM�'��u�?��q	ރ��ސ��8�pU�i0���� }G�Ea��>�����\�\Y>Pq+�=P|�DF�Ĉ�Dh�'�p���w�}��I�\z�G��7�N[�_������8��<�|ONӧ~{�s�F��]�|��]��i���	4�>�xǢ���X�� ��ލ����<�v���ڷ���>���d�X��	 }�����>���{�������}��G�8��:��Ӹ�_��u�M���wg�\ۧ���;���z@�tE���P��DA�v�L��w�揾����}'� ��{q'��t�I��ӷt��4��<�����~'N�OE ��k�!׻M�	���Ͼ��88���u�8�����6�'iSu�u`� ��X�m}�I�[�Ng��>���;O��e	=8���8�w�~w��wPt�U7�����hq0�������m�=|��t��q�9L.<qw����	7�B����3�D��NǠ{�g:i�ia�ߟ���
��q�����N��&[�;���J�]���r����Π�8��7���0��n�?q�ǈt�U���:M�oGpq���8�Ǥ�F����>"5�\::{bƩ��>:��&<�|��ݫ���O��ޓx���]��?x�����<��^��;���8��Ǌ�םp�7���S�}{����}�~�z��}wa�"���H� ���:��L�G �q���J�D��N����!������I;=����!����I�P��O���}�;L/�;�u�Jo_|��I��|v�=tc�=��Rq�M�	ݥ�y���x<��?O�g�p�1E��rH4�^��'Tr�U��<�\ܝ�������<��p��7���Ai���O�/;�s4o��#�Jm'EĨ��-���bu�h��<��<1
�!@�lJ��5=�)W�R���o��}A�s-����6x�B�GU���Y�����O�R��*�U~�u����a{�#�n�v��ݤ����~��~On?8� w��=!���7�����w�>;�}�ϝ�av�����'�8�����K�Ă����G���&Vu̥W��-돸DF��������~M�!�ě��ogw���|@������&޾��>���뽻C5��U����`{�cW]�,�����Ͽ>����q�L/�Ϝ�N�}BC��2���8��w�ސ;I�w[�\�ɸ�S�v<wH~M8���&���O{>����>&����Î�3��N�s��!���">������X���j7G)��>B �|�{�q���DE�����y������ۧI�>���0��?S��L/h'��}C�����Ӿ��9����t�\}qu�#E�� A�k��7W5��үV����=����y��e:C�i��{���
^��F=&�	��뾶���1�?'��8���H��N��$�+�僉���S�q�����}q�>�>��0�"�gpk�SD} }�n�x|��:L(u���[�C�~C��-�ۉ�ɹ��'v�����ݦt���s��o���8t�q?�X8��)���?'�ӷ�i���]�]�+�s���ۈ������7�/��;�}������z�������!�s�&�	��y�:@��o�I��� �㷴��~w�z@�N޿u�ӿ=&�a�y�[.�ɧ|�<6@�w��:���"�}B ��(c���n u�8���wn����o譔�P��:�������;���=s��ۿ#����?t|v��n;�w��� @�
o��� �>����^�3o˶w�g�؈�"$DAD8����:w�}C���q�����[�Ѹ�A럐��һ�ӽ{��:C���>'�X�0��>p��I�!?�G�����D��%�����B�}ۧ��{v��>��B��q}#>�ں>�#�^���u�������{����>�}O{����]������4�S�V<wH{N��]���Ă���� ~D}�w�,��#�၁�����1y�3Ȟ���N�v���̀]�CN�=V2������ՆDu0(���)]�w]�ӝAa�(��ʀ�X��JohΡ��[եR͓4趆�0��6D�������X�ۏ�C{X�sY���o�v�ߪ~�T\N'϶�s�
&���Ӟ���N�y�����+�G�p:M��o��On	|x������aw�v>>�x����n+���q=���ñ5]>��;��aq����"Cٍ�v��N=��Ӻw���@���v�һ�k��7Ht��'����:����w��8���wn=��zL)���ǳ�s���ݡ�t��������O�g�����S}U�n"����b�����ێ�|@���w��O�v�_{>������@����x�wN����=��U���8�hq��:�q*�^�� �C�i��z��5F����X��_�!@!��ӁM�n����{pq��;u@||zC�����$��~tv��P>�����x�8��x���>��8�ן}���i�ސ�s羷�i0�����D��sXm�vV��hG�>"!B"G�}sn�Aw���VM�u�t��n�L/���:W�	ޏv��N'����t�Hx����󝿜�i���0u巷q]������[|��w<{�NZП������D���Vׁ�����;׾{M<M�	ǣι��۴�|x�&��=�N8��'z��N:w���q����t�������D!G���p��c?p��W��%%F~��;����k���C�>���I�=�y��zW��'מ{�i=?~~�x������u�;�k��x�U���u��zL/�;9��U!UV�!�W�G�>�*�i�qp�򖱯_o��<�@��U<�������ݞy�����8������C�i�~��G�n�
��zW��p:t�u~@�ˤ>��8��zOޠ8�|Dg�} Uz�t>��z=[�efc\��PC���C���?�������|��'i�ߑO���HC��t*��H|O�sߞtc�q ��;��[v��I��q8�v����ӧi_��y�1��N'��y�G����[���Nz\}""�|DFqF0E�pN�z��>�⾻��o�_ ��x������_p��7���L>���S~}&�����p]�I�[�9�+��ﮏ�uW�ԅUxQ�qy7O���n]n�6�J�Hd�;��\�*�+�/+�ݲ�tYb�g�gJ�?~��w92Mo]�7�2�;��:�b��[�t%utjӥm[���c��|8A��:�Q��	���Ge.�t�t����.���7*¶�db|�93'j5�:۹�`��{����h����?|��~W{O]A�n��|N'�>��n?[~N�v�������|������ì���;=�{��7���Kޭ{1���yL�Kn�
;'��"T;[����&�g�7W�����D���Ozf�Sf�v�LXɥ [�=�o��SB���y��&�.�U¨�P�ǱG��כ�ሶ7w\����@������t�p݅}��O2<�k�k�==���D�n߆��Q�J�l�#"�qA�'�����j]eD����q?
�(1���c�r8FZ��͔�!����kD�zta�����7�_�P�"��C/��w�x������٭�j�ؼ��{���N���ҍ� �w�a����&�Q݌����ҭ�Oo"�c��{
����ζ��h�fr��ͪ�Ǭ��aYuW��\�����~ g�����^c[;Kzux�!t�~����v���`�p!��oJʇ�41�����[0��]o���um9|.�!��gl��5u�q�{�~�$nvv���é��}_�x��y�[y���yx�ݹ�l��5Oj�Aζ��	�W��o\Ñ���yPTWs!��?V�]�,�[�Dԓ��ێ���v��xбUu�q�b{�ьͤ���[�����=gr>����ܹ�u+��nq+y�i��Y\gd��l��e(7Ut#�X��ۥ�d�94��^��}�t��݄p�&�o v=e�{�����������S�ږ���׹Vj����p��N��Ӭ�ص7�Ϫ��|}�ɚ�'=��-'���[�coRP״�Q{O����Y��ci90Dk�I�ٰ����Hd�j���/j��6�����+˘�@.�� '�|y�c�I�X�5vϥ�/a�{�i"���7���g��w< ��`����K?w6�K��<˹�2�h��u���6	�+=s�����O���K�(���\���&,7np#횅"� rY�e��؂����R���v���O� Я\1iŇ�t���bx��c`^<���*�SWTg�J�`O@qnm�\��m���d�w\���L�&Y���{>S���>Ҥ�W�J茵U���vL��Sՙ]�+�Y��C�Y��n�4���&��N�>nlu�C7x�Pީ����ȵx_J��vg�ڮu�-ՏC��<:��[�5ɕ���mT9i�����Z��邥힊�\�t��g4ָ�ׯ�<K�b{=�����0�A�ko,����8l(,�Ӌp�Tx���s.,�j��2nLr�35A��*uM���7:�0[�`����C���@g��qe�e`��PCG52=�ׇ�!����W�t����~�&B2����z��╘p:����}km�;���=#�o����z��#�J�gC8��K�~(Hw��n�y׽�Y�//d�!(Z�h���u�%W��X`��C� A{�G?��f|�p�o%i�lZ5Qg�"kI�3��?l�\����P7�q9��	^�U��a.�Ö���+v��ٝ�p���y����_N��C5Tl�>f���p-��E�3������N*b��TG]a�w���l��l��q��h\(��EN�ҏ+��޶��Ks�	fWN���Q�~re�ʕ�ҩ�mgS���M��(p�W��SpsǆZU��ᾼ}g����WV��^�;:��:ߊ��sY�g8g�z8h0r����檻%R�P+�����K�N�}"�9g��,��_{��ু� me���j6-�8ʞ��]L7Y2����ԥ=�y���2��X�yr#����͌�_�;JO��
�3��=:p��t�K(�(��9�헗�=��/�mh4Z��ɯ!ĕ^���?Qg��J暆/�ۜ�a�5����
�_�K�.����+K�,��>�7�Y&<8���A�P7׼��g//��6����aD{�I�-ӹM\xw��e���+�{��u��gI[�R����J��D����#JF��1;Zdg�(js 4�s��魗Ӎ;
2��d'�I�xk:��;,?o��zؐaȝ�ڧ2E�
d��#����˻X�&Lt�`n�Uy;��&����{��jtH��3�JvD�*\ȤhTw������8ڷ2kT����c��h������ёV� �x����h)/aͥvKxO��ѿ��'����'4vV_[���Q�ʁq~m0=�R�~&��#Ƒ>{�P{��]>�~F�$�̊خ����V�@�롛<��Q�UK��� t_��0����b��2�d�C�]�+����Uq=��:�z���7X4Ŀ�uRg����w��y�8"?{�o�PK��O��Җ�����P7�/?��W?���ϯ�5��^G0�]lOIK�]������T$`�i�:cU�s5!��[9^h�����Q;<'��L;���ɹ8���g�Dﻔ��E�Y��9��5�*FxA1+eԌ�ڠ��uʋ�_�� +�ؐ�}����o���H�z��.Nm�_G[��P�[%s������Zk��>]��[��Ԃ��zcV��,ଊY�]mD�h[�U��Ձv�[5�t�nr=����
�<j}RK�`l��۠h�k�v%ƈ[��ܫ�����#��g3l&Ӕp�Ѹ��?v�[U^�2��;�9{.W6�L\)����3�))��L�����Id]Jۅ�ʫ�5K3�:NG��0J�6`w���~��\��ڭ� NN3�����o^�yb� �ܥ�ȑP�ޭ����������'N�E���<|5\@�-p�&MEڋj%s|!��t���з���:��w�Y����I�R�fr=��J�=X�ZxnkLSd��I9=���8z�e� ��W9�&UeGY�$%C�����UUm������%������P���b��/d�̅�Ȧ� �=p]��`L�<�+��P�q��Q��3T&�;:�R�jo��Gv<�LO0�D+�H�Ȟ�u��@{�hT�VY�k��UӼ6���&��JR�*��{�[��K��~eW*�u�\ ��ބ�p۔W�-�2<,������bV'x���f�:�`�r�L�Ȯ���y3FH֮!�"��
U[��z?-M��V;n�uGΑ����)�FP���~�Kf��ٚ�*+����&к����a�jfr,�!;��@�����m��۴�t1BV:�"v����:�����njW@3lnz���1�Cs�>�K�q�5h�u)�n��/6�D/(��r��
�s:b��H��]2��<̷�.kvǗa@�N�i��tsd�:r�ee��k�n �V�����\y��[��ۑ���]�}Z�x�8�d�bǟ�X�Y倫��7x��lU���WT�Ψ���W���Wk�1�}�0׫�٢+D1W��xJ�|�(��/U> U��dJN�K�����Kx��~��=����M��g/����g��\ �>�Sh��La���������j�D4��ǵ碗��4Au�˻އN�V,�C�e��b�����=�����߳�g��Mh�6H��D(�N��h8�!߷f�o:ݚ�E����G��V�Og_�Ixn<�T��V#��f��Y�}�u��ٰ��������9��#�F_�k�o��)L���Ѻ=d��Q���~bPMg�ui�--�g?����!�=��:}+$e�<&�;q�t�m��W��*�X��O���f�v���
����c�J���Wl��ap��Sw��:(���Q����6yc�78&X��h`=ˉʳZ=r��m�R�]R�d���	�2.�%{�[��ژ1`C�Uݹ���B�p#W}W%;�#������	z���醹lT�����,�T��F�e�p^�}�ԫ��@�Ķ��t^�$��5H0M&����'�\K��"�J�e��G}]��̘�S7Y���yՓ��ݭ{`~~����N>�OmY(��q��a�����;�jwCC�q��|�g��������kwn;�0�g�TG�/�]	L�#|���$J�&�So1]��{1�#�x���e�ަ�X|Cg{��<7�IQ+��tFZ��O�I����,�/��I�.���Uр]K�}���FlG\H\��:
g�f��ry�>��)jl��O��Ƿ�p�ܩh%]/�V9��#\,xe}���f�O.�V]��q�Z�[*������K�����{���>㚣��k��W�uN���P�b%vl�:���mlFdX�Ii��G#����g�?��N��l�g�{\�^{�@�8�3H��u=~Z��Ng�L��k���y������2j��ub��T���8(҂�i��L��QoS���l��=]7XwT`ݔ ��Yq�K����Vt��͍��3u�'��{9�)ۢ�J3���$h��؏蝞�if��"�ebU�y��'�!�q�x��O"�آ�j��4�\Л:�!tn��ڵX��}m
������ ��o�>���
W�T#�m�Ӊ��p�pP}���@��rТuYc��71���b�<�$�"�h�k`�K�י�����S���]k�C\�i
M*�n���Yd�%�^;=�%+�n�&k��
����b��r�`��(��5�l�F�[�n����©�ˊ�z�CF�R���;cLYk�]J��f�+_]a,]�S|�cvZD���O����H�#�����M�N���L���������z+�h�+i�D\�\A9��YX���;7	L��S��
����W�x��gi&q!(@�B��}B����u����z]NsH)A5z��u-0D[r��t��9w�t��Z<'0��e�[6 �� I��`�QV�vR��άy�ܫ��ν}έo2˚�����7\xZA6 ƌn����*\8��D�n�,�x�6�oJ��0��M�ˤ;���Z��l���m��Z��T�B�Ή-�VhG���o��v�ԵC�%B9ō�C@u.�S��cr�a7/���o��K%���yZJ��w7��4���e��tJ�x��"	*��e\��&��Y�
4�bT�sF9CB�ܶR���V�T�&���alLi�>�zP��#B�_�J���2�l��Z$�VuwRZ��J{#��݂L��(v�f�P��x���Z+�m�1�u�r�M[C�⛔�f��)�Y�F�$��	�Ӵ9Zl�P-VkK�Z��l:kkfgX�\r9�8)Aڭl}����:�L]N���4���N��=�MnL����V_JC%ui|��Ra�����kw��e�8J��#�9r�o"z;�K�^�:h�p�7Uc]=a`оZ^$;��8����9����5oMm���]rm;��n�N�?'���̮X����u
��'!���T�[�?����릻�ƫuh�{�L��嘛�
7�>�9��g�7�l_K\���V�l.9�y	�2�>�sZ�Zޔ�cEDb{W���Dn.�KȐ�K�HB�u�gF��̄f���im��3-ۘ9�.���TƵ�������󲖊|��lU|x>M� �_7��v�hQj�l� ��(Ըz[�E��ճ�1ۑe-|'r��y�i�G!�f� �õ�2�m�{iЧ3���ʶ+��#h� Z�9��� �����	GZ�c�2�!�����h(Q;)62C��}1���I`���isG+�<f�XwqpUʭ�A��iu.�m��ܧn��]Z�ِL���\�ٔ!!�c����nX��� 42�� �W�k�B��r�hZ�je����+C���[27��(`�%hm��0<��\���wd��6J�Z��H�I��8�K�g,���d��$�高�-\%�';X�Ԟɳ���k@�f
Q�&�;%��'���i�&��J���A�X�]���J_]flU�pN�r��Oz� ��t��#�.Wwν~��=���{���'e ��ŉr4"$�aEAEY��^3�	\<a�

%I����Err�E]�s�Q��P()�]P*�Ă�&��.r�Z�s��r�VB*,�B�<�����t�Q�(�3ds�*48\���(�Q*<IPP\���p.D�
��(	S��UADp�"�*��)��Tq�*���r.ʢ�����%ʊ�죓�����T�H.șTY%ȯ.;��*����EDh�ITW
�QP�J)�Wj����9�Q8�˲����\ ��'��vb�UD8�@QC�K_g�V�K�Y�sμB��@
����Q<��fkj�7[�i�M]l��C�s9��he�Ի-Th��x�sQK�(���ctr���	��Oү�W��I��g�	UiWO����T ��WB��Di�ݯ�ά�{��~5l�y�
j���Z����K�Aw '��x����[צ�/Aoڈ�>;
�a�}a`�V:0�N;H׊:3���
V�8�$����ƥR?G���h�����@�X ���{]�ǟ1;Ǹ>���Q�v'���EHnY@o~���\�����%-ީU:�*Mj�s�垀ɕ��z^�T��>x�Kȋ���;�u�Ѹ��VԘ}B�����4Z���zUq��6;[�0��:'��YY�y�w^j�҄c[0�d<z@Ld��5�1��+�
�t�EZ�|��.��n����Y��;�aޭ�H�n�r��1Q���R�7�=wo���,-�of}^�F����m������5��	E��8��K�p��7+��m���ݏ�xh�G�=q�o���S}a#^��+-8���v	�s*X�ѡ�7�N()]Ӝ� �����*l�8^êaa�s�a~�^��x�^�A��{Ks2���a�=�,�k
�[[��z��.�4�v�c>��0]�]$.�vM�(��L� ��{쥴�Z3�-[ê�tuw)��;j�n�����nA:h�,B)��I�'$(N���t+�#�tiާ����:���:
7bN�Jߣ�|�Ŏ����&�W�e�B\N͞����+et����<� ������R�wrϫ�F�s��+��僀��Wf�g���[�
�<��&��eTm�֪��'�ɑ~M�g�"�b�g�ߕ0��}+f�=wzߦ�L�o޺[:x��_�orFڭ�a��*�!�tJ�u# t�]65�%~3����d����k��IFWI��,Ջd��wF�g=�+�a�۬�_(�������:�N�Z��/�y�8s2j�Kڣ	OB��R�XN������+E�O��-��\Z����Z����.�����Y�w�����S2*��������N���r��b<q�S`V�����>�SQ��P��o^ +C<���hY��]E��F*:ĸ0�w6[���U�I�����"�*�+,�r�����v��Fȗ�N�*�Hi;㰎5���p�1�Ç��5�/O,h3�˽^O=0�^�܈�R��̅�Ȧ���[��W"#aܙ����~Ϫ��/wJ=�=���&�d%��*D(���2�c˯(����]�@e�񶼶V�`]�B����Lf�6f@eN�tm:�t�������Ik�B�;���`4w�5��lhq�X�!���%2�2I|�ꂸ��6S�!]9v�D=T�3z������V3�z��O�����*����A�6Rۂ:2iHUWUD=��@��c��\�t��qi����$�iCo�x��}�`�z�t�@JJ�n�Y益��n����]=ޗ�8�m#Ygg�R1Z���X���� 5ڸ��"�V�N��5���;�V��������Qv�p���gt/�ZF9L]l��w��U@#2w9�5�k��-�GUL�
}�6�H��q�$*�Q�ƺؚ�j"�v25S@Gm���^�ᗧ���9��7���̆*o�(�ڷ\ �B²��#������[�[S��R�3�7آF��zb�1f0{7�'��L���� ��簙~����v�<���� �^� �^����r�	^���Z(Z̽���a?n�bf_Z�|]|o�C�~�w�^}#��b9ODÂu<s*6�q3^��u��5���辻噈#^����f_�s�KF�M�
{ezZX~p׵V��\"\3)�ra<�b�M�ѩ̎��W��[w�N���z���W&,]��BR���Q�0��j	x�t:��N�r�{�:�w���{4��:��,N�AY4P�O���e��/+xǻ���\6 6���m�˞��N�6�0B���[[9Wǖ>�Mx�nM"T64�W�UUc����$�dx"H���Z(����!��<,�����x�>���=ئ�p�#���(^��g𒼼���`���QJ���f��U��}��V.��X�<n�nDb��gB���H[\o��-Q;� ^%kЇNB�q�%6R􋺃IZ�����U�*��lpӛaB��JX��C30b¾���'�HG�0�P�5u]�\{[���Xޥ��	��۽�\����'o�/v��v�y[ܞLlwS�y��Ǐ���kS��w����8��R1N��~��:����)�A̕7S�}Q`9g&D;��U��I�w��ͭ~�z��`	�%|��<��s�
���D�6'�$+��D��ي���WokL������9t"ߡ���Z�S5R:���6+N6��Ar,l�67�&TD����v�;)�p����s�rh1��!�.��V�&&)&"�ɩjw=�~�q!\iey����t 6�Q[�.������,.ɱ�Ҫ�E�r�y��@�y�GL�y��*�r����~H<��N![ޕȬu����6��ٻ ���щ�Ha<��]� �A�y*ܿ���i3��k=�3{�_��C�G˪Ѥc:=�Y=Z�Hv���ݍ�C���8@֜�3q�9�ֺ���5*��-�+��y��wX�����
p��������[֦��M�;���8 ���Q�U[HN��2�_��dᬯ$F���PWK��:�;�:����{�^+;^;�>��Q���|������O�`:j��fU�5�w�f��sC���aX�>G�8��3:�0d��6J*$�I��FA����\���Q�hʃ=�g��N'C`6K,K�!�8uD������R����O�nK�\>zDI�;kw:�aS�nN���M�������U��ǔ����Ǆ�Ү�\7�{9������O)�R�v�a�ԇʭ���"r�{�>S�檻"�P+��lzg��t������}������:��](g:�/�xn^zp�<�	�3Ǯ��?��Ƴ+E��y��/{��V3���B�Cr�m����|��:� )>���j�`��T)j3����/)ķ��l.U��Ə�䦐T|�MA\7�J��.�gE��vM��lԙPVƼ��M�iot������^љ�aР�ĉ�GzJ|��ģ�l��W/��h����NƆ\U%z�w`�Wmȫ���ocaTN�A�K�ӟr׳�[��y\�6��E�DsF:�Պ�;YJ��M��F������ԨX�Нfm^��Y�/kf�b/Z�Ys�K%�����M�:I�	��ا�������WV����UW�`�hzW�x�fU}΀�wbmM:�����^7.dg�m����;���V���զ_U�.:���[�tn!l���7�_�](փ�[�"õ��KXeV�
sQ̔��t-�
k�8)/V<z�G�!�j�Uwə1A�r�g���iYgc�R���{���NW5���S��U,��fng�q>G�D�Jec�F��q0���-�o'��r��H^�ޑ�+�6�0��Ѳ��U��;��k������N�T�*�aA��:�5s��
����	���V�\�^��P���>��*뒫3W��A�'��:��{�0as��^��g:E_�ܙ�cL��E^�U�(�����W���4=����ǭ_��U�כ����!�����۞�e�^�G
6��c�(�G�\��Т����bw��%ۭ�S���GA~|��t��oy�g�����Up�;)?�y��8�P��f���x2j��~���yT����,��9G���*�͘.���[>�0 ���������x=c:�]�/���c�� *=�L=ny����C�ֈ#==��уz!�E�w�[�=��I�Y������~9-����յ��on�.��y֠�lꍳ%ԻY���w�a�+�	]:G!8M�����
u(��muw�U�UW�lr�P�O���n���Α�P����*��8Z|<+yI�����#4�r���{菛:Q�W��
�@vJmu���:�G����x���+Ή�e�7W�>{�͊�P��3��.� *�Hk�W9�$J��0J:��~J�N�a�UDl���3�&t���ޑ/�;���?��l�� 9t�Gl	nlH����H"ga���] �K�u�=��ۃ��4&�߱ۇ���gb{y���b.T����.��\о����	�ڎ�o��"��';n�\��' ٰ�r�q���rem�r�`�x����W����~BÛ���Y�M�}������x6���Q1bwd���y\�K��M��u�>]�)�ً=Y:���U�S���n��B����q{
uV�aI�����Y��4�Jc��/��Ƨ(��Q6�0#S3Å��i�mxl5vy�V<)�y`)����>U���߫�O��eNη������f�)�rd.b+�碠tl �a��e�|�(��>PC�� L ]�|��|���?���Fuuobܛ���=��~�:[����o0wW~�� �xk|���/vn��w+��[���WZ�G:�[�	>�@�ݾɜ��y���<�Ü��v<oo|�n�^����'r��x�"��afTq���]
��7Sg�| �ލ�ުK�6@y1\@��\��R����%���^��F�E�� �Z��?v�G��.�i{1�U _<z ��_0���颟�=J�`>�]y�v�Ӡk�{�C��4�>�)U��z�H*l��DC�#S�2�C�y��t�s��k�h�hz)�.��zG��|�r|����b��n�U3ҺZX~p׷��Lt���9]/$s����R0��lu��I�f��`��v��\w�v�Q�I@SY�C�<7�KG�s����6*-Y}�8��������F=^�\>5W]9^�?C9s�(�U��|y�}��z.��<߫|�-/���x������j���pK�2ի7�Fxǒ�uHC�w��wg �J��BRo<d�Y�fx��K(ycaŊN����(��=��!ڪ��s���"� F�¸[�[���X��9�hənt��8�gb�]A�BY��G��B�@[˘
g�b�+���w��17��5��Ӗ!�(h�:>+�t����2��&��u�.�K� S6���8���]"~B`m�Iɳ�u�׮,]�)�ܗ�3n�;%A��p
F���p�֖��0���yG����4r��>���4��^Y�n4�:Ȅ�z^�����F�N�eC��叕�rC%�OV��}ێ#菢"$������p�ڨ  v��p/Lg�OgH�Pc�$-J�e�C��F��R*8��};�rú�	�
���%#Z/)7]r�Վqxb5֯��Z�1Gl{B��۞k�����ڨr9U����L_1�p;�����r����g���Ȫ��ǧ15�	��Ƈ�Pp���������<�����ҫ"<d�gNU���>�3]�DR;��xw9P��ި����λ����V�u�=�����i� ,?��UN�T%���31Ov9�{���L�Rc2��f��g�@.o�(A�ӫ"9.L����|x����]�6��ݔ�� ���{NR�c�N�KK<�g+b����i�]`���B�����*�IXSj�M�7��>7=.@J{�͘�!�v���W�Z^����0j�4o��u9a�D�y��g�Z��p�n��mq�>:$(�)�V���u�Ta�
&\)Ss�'���î�[હ��SP��U� 4�b�J�
����G�c�g����Wd����jM-G�R�V���]7�Cu�C�\uL��4Z�y�˨f��*�Y�7�3�Գ�ǥ�H�;��Y����t;u{�m,9��1�U-��T���%�:��n�j����?���ج]yRA�[���Wz�{1�DW��x{�J�÷%8�[�ƒ��^��l,�V:0�O�{��l'�Ì��J���SӞb��^��z�G����hf�����}�ܭ;a)������:� (=�W�Ǐ]Zx�g�d��#���yMͤ34����H#��j|+�����l�wHRi����&��LH��T!1N/���{�}p��ߑ�+G|h��ޒ���-�PW/��h���A�nbR{�n�)D��=X���Fq^D[K����}l���� mU�
�"�q���n���������	�K�Ϗ!�R��zU ����co�q}�k�������_�W�z�N�z�OG�lW'X�Xu��|)��s�9!<t� ^�3ƥ4�73/-�!�qY��ssR�!J��lv��v�$	���
Wt�r���a�8y�p\�+��/R����(���5����6Wm ��Lp���^�'ӑ��38"/v���]W�bN�f�US��#p�+:�+�5U5>e�)�L��S�n��8
�qXve_!�R���J���Mv�JvV�-Qm�F0����U�#u�A��3��	CI~ʿj�r��=h<7Woo@[kzޮ[ѭ�9y0�-b������X�w]���J�7�	���W�4+2���r]�L����/7Pn�@Г�'�q�q�M><�;��{f��Vi݈�V[����@;=\>Q�Ŵv�2.�V�UY�SJ��8�����v��c�}D-�{2�9���'��+����������{i:�-6�EG0I"�/���Ǌ�΂�pFp���wG�+�aU��J��j�i��� +y-�rn���C[�+�����&^mnoYP�v�Z�rۈ;G>�{��7J&*1.닝�Y��[&�ki��f�Z�ڶh���٬�Ѭ�	+K��p�V�F���E�H����Ot�jv�#P�Ի������V�a5p���ث��	��Z5�-��=�)Mӫ*gE|u���([�x�U�VG^��.��i��wz���e�ӥD��4Ռ��<t�A��.��ݽD���g0 ��J�j��VQ��B䮔IQ��qgn��ˁ�#�����lvn���]w-�i�w��L��ǜ.f����n��=O���<�S��,:�Y�5Tq��~�'ٶ�yл�X3V;T���<�|$!���޷��w4IX���&�1��h���9Q�T�ű���[��mP��Gt��Fb����Y�T+�K�6��orIۼ����k4!]�b��f.V�#��:��꽭U3H��oҍ�C��]� k:�u���7��F;�NY�qƅl.ZFuc�f(1��O\�s"��f`��]���ٿo�-q���R����s��H``��93��C�C9a�̽"�u�Pjc������]>�:�ĸg(�V�y�vp�z�:�[ؐ��5�e��h閃�2��U�XY���/38�|:��4rB�����
�>�WGأ��8v_)P���6_CFȭ���hj�-�o"��Gtj{9C�e!PJ]Ռ�|)J��E���17��WZ�i�o�nG�N���L�wnξw�U�~覕I-����)��H�D���SoE�L�m��[b�bZhf�o�\-[\)a�2ƊL���Qy#\�9��:ᩔ�D�+��kt��j��!�R�E��x�f*��^,���f5�mP�ɵ��뙵O7
��1չ���0�/���gbDRP�ɬ��lJv�3N�ۧv�,=�*��/7An$aIV�5��*���С2].nJ��Y�^�*Ƭ�5|W� o�J`q5�R��df�k���:͔D4��������"q�M2��z@ΧY�`j	���i�\:޽㍽Z��i��s$-�w�YW���䩇A}P�+K�eF�_q�q��*v [��̀*�E
���
����J�"��duC�T�	ʼd˅0�+�ʈ.��PPT7K��"��ᣉ�AEP�����4��ĕH��#'8�IʓKD�[d���yU.\�5�5���^3��5*9^S�8��!�)�8��q�x�)W.bR�dL�.Qs�LȻ(�"�E�@(���ED���Y���p咄I)��rpi�t�؄�.K��D�\I�Qr�knP�x�NJ�x�3�O�d���x�q��ĐP���L�V�pTpT�r��G �9��+G�®	�8[/^r�2�p� ��sp��!�9'�T8k���p4��Q�4\K<j�j<���[,�t���Y�ivc��
L@N�w:�ݟ�J�g\��Q��Y��C8ggk��-l�;���꯾����t���X����=���$5u[�Fa�h�����U�Q�.�ł� ����#9�ٛ�n��v!3����{�J�.+�sF��쇍Ava���l�������H ,��#9�����nX;Q�U
{Sǲ_;C���y~1����.ԉ��<�]o6���f��po�U�O�0��U8�<��Ѽ��>��uK���A��]@� �t���贎S��wr!�bB箩3�ˬ���;tϰ�>q�)ˀDK�D��w��Z��<�e.�a]�Of��z�ۺ6%!|�q]V˹��)�u�&�fQN���k[���c��i���6*z�'�fB�p��Qu3H�K������'q�ռ�t$�n��n������HZ�`=�ܕ}WՓ�6�9'QUlB�gaߖ�ͅ�oC������K�T�]�d�J�c����q绚��]����$o�S����e9�%`�oV�Do,*gwFW��e��M��h�ۻZ"I���L��	�AC,e^���	�����hfS�j'��|�D�d:�޺E��ms��t���rx5^�¹���Mf�k��1��fҮ��a�����k���2�6uw ԼT(�s�+rp��gAJ-9;���(�ͩ�'*��=jt=r����W�U}�pP��K\}Qd�CR�-P�h��=+�ݔ�8�۬4w^gR���14�%���r3��]���qhǳE� �^޸VT���"A3��&�m����D���O�(?=���W����b���W���F�}&^�f�.�g�s���0tvF�Q��O�o�b`�;��_��\���jh��|��o"�>��ܷ��9��s�.6��A�� �﷧���\mL�`�X5�
��^>�oX;M�rly��?%i^��I��OJ��j��*�I��C���57�O<ݶ�mر��J ����1�����ͱ�� ��=zՁ�U��� �W7᭛M5�RH���50au�(]�Uɾ)���W.r�Ӷ��M�����6�����gVM~�;�omVr�Ӑ�a݅(vR�u/��7�C�S��F�d�iqݛBj�yf�V{������a�zX9���u:�r���Rh��}���G[�TJ�/�Ab�y��%�(:����L�ڭ�G�.V{E�@]���&N��&s"�L���gtu�	4\ ԡ��*�*3����Ρ���U�fܢN�{������ꄞMP��ް�[l��`�v�gPH���튝�3W���e��O�򽛝�cN�Wp��	�64�1���Kr�q��[���$K���s2�'�e��ߢ'���������9|��v�|o@D��Y�����˻�q�*���U���`������eo>x��ry��bu+[���n���e��V����<n	�o��iq�)��,�녙�Mv'q%,���n�>�%�z9X$4\�L�;6��	V1�׊.�!���^��&9Zsg�JQi��}�Uc�B1�;�;;�Q�X��2s�V������!�e>{RJ��,[�;a�/,���D;�{.!��zf՝�c�4���sk���F�)l߆��m�S�?oj�L�l���i�;����Q�ƕ:���*ϲ��b�e�@�+݌�����qz��e���U�f(8�Su������̳�f��=힝���)ׯաYx�Y\(Pk���۱�jͬA��3��i��r��G!�g7b�H"z�����4��3{ �Q���m��܆�CPE,3[y����=�f���g*�z~�����f��T5�H\�^]G�3�w����������\Ȼi��9=п5oy+�5�J��<��7���Dzp�涠���t�,��r�����z����W�1݅E+U�NV	�@�����pj��cG��&�fۜ��V�
���[{]Փfusbd�s����r�R��׉5��w!�?>ڷ�P}��έ���K؞n�S�v%�j*��C<�����=\�`7�KG����l����X@�X���u���D����{mڦ*��� %B]u=By�`��0��>��x��o�s:�x��7���}�fx��V�O`r����$R�rs
��;I�v�h�F߂���z�g�AW��ȿ)r*X]��k��ii��%����[ۡJH7E��&��}o4=�]n}�]/�?���]��W�87u�լ�7��Y�%�%�y�ě��\��h-�\DN��ޥd��=I1�)P���n+��
����~��:T	�5fKT�L���-�1uE�Z�#���:��p��Æ�NPЏӚh���;OV<!�.�h܏+�4��4�{ �y��d��yR��EuЅv�����������G����}��ϔS7�~]�(�.sv�A�3t���ʕ\��&G����U�9��<6-)v��`����}�������[q%nz^��n����4~���;���]�`��h�Uk��j�T��^��0#K_��=�<q�[��6���[^ˋh.;T|��R�^Ѩ&�c���7�e����ø¢�5'%��I��fך��T��^��U]����E�N���}US �x��	��y��{�~����n�/v�Ά���Ly�7:���]^W�3�I��;X���G�>�kŽ�x�>��+�9j�/���h^��z�0kdvź�oY��y/�T���\>���U�x���r��zk�^��]1\ΊW�H-�V	��V�, �z�tj�(>�]Y�u��]S{x5��&�_��-�PWnP[�����}�V�4��K�q1~!�������z�L�eM�V%��u)���XD�</�n���՜���SǕ�N�ggƴ����\�~�gc׬�oM�x��q��6h�n��U�꼐��;9a]�q)�2����F���w��U��1�����{H��DN��|�3�����}U_|7�*����v���@����`2�����'�7�Ɣ*��F�e����u�9iB]����Oc4[�"�n�X����3���n�ϼS��M���'����%]��*��C;����j���[
�gN����tŅ�"��',��t�&�����`�o:�)�{�!ve�iN�J���A��M�z��x��!guJ rsvA����d�A�n�S���"��`��=U+�R��z{����Vn�ԛ���W���C��jsd���τ��DP{��>ܝoh������3.��;�^fKzߜ�hQ���icu,[�:�T���#r�G���1�#M�&,Mf����7�i�ݛ���hY�|��]��4�/��<Fvq��{��a��*s�m1���D�|d��=�(Wb/i��k:��LlBW3�<8����"�,�1W(n��4/E�Eoi9�{K6�M��2H�W:��U���"��C�]wQ%)��[ƒ�3�	��AC����"���3r���+�2����Ub��u�����w�:��䉔�s{f��|*�j�=K���q����/��W�U}#媘�[��Wʉ��g$��]�9^�=�n���yzn�t�w�!\~>T�Fc��p1�u`�V��Z��$2_,�J�[2.��ƽ�qB�J�o�����z������>��*Ħleo
��!ss��#�!�n젺�)\�b
}�j-syʳ5��a�am��O� E�Λ��Xk8��P�k(�~�U��݀��p�h7m�NBY�!+r���!]�MvM�R�5�VX��,ch�+�^�O�as>�&��Jiӷ=�zɳ�g��x�c�p����j�	vg�q�:�ԧ[kC8�Bp�n�iGQ�fPG{���Z`09�V j6+�E-g!�8#Q�|�����g�;���;�i�2�)h�s�aK�v�m�@�Ƭ���X�gj�wK\�E0�x!��M��[���S�XF���TJ���tɬ}Wo},c8u��U�6�䨞we�w�uv�5��Ȉ�/,�����W�=�8E�Q`Y��R��J6M6�w^�[�1ē����K\���^z��-<��.	�bu�|Q�����{��/36���/��}U_}G�I^�z�[K3g,�t���{�F"�q������ë����TZ�s��{e����olM��f5�,s�;m�a\Q���F/U����&���|=���Oy5	��r������GAh�WE�_r��eh�c��l:�6���z�Ѳ�z��ǌǯf��\�/B�����^j�� ��YPv��.���Իa�N���-͛-�/
����k�K��~���9sy+�5�J��Tf���ZQU zvR�2[�8r���T��|�3ϋx�«�X�TR�g)���ژ�v}K�&�&�ph<�[�+><�>�ڱX�_/���턯u�:إ���i�:f��~w���C���+勯y�؝]�|q��V�Y�±'��E��g*(����*r���15�WP�X�X�ڮ��62z�^P�[�X,ct�V���^쮥�l��KS՜�IދorXA@���h=hV�Q��{���Y�yse����k!h�uu;r������-77U�~Jdݧˁ�5��]շ14�unnEP]��O�f��X5M�r�L;��������F|]���������],�s�[��	�'�������N��Y�E��U|r�\I}lޕ����0���&�[ȫUҜ�z#~�4���Ļ���8�Uo��s�5T&��m`��'��!v<�i�>��	ո��cq�[q]^=,�Z�v�>=���K�4�V�X`O�G���Kݙ�.��-/I�+W.�[Z���$i	'�V��]h�k��X\��`�X�X7�3���56�ٽ��j̚wM�M�ÏF4
14q;�{��sֲW_Zw%�l<�yu(�UE��u�f[���|�7�y��6_D�3����.�(�rj6����f弌:�i��8�V}�V�
�l�	���Z����A�װ�og����Vr{�$A��(��D��L�q]��L�c��i� ���cJ؋�>O�����u�an:&9o.��T����v��ȷȊUy�Ұ�G�wv7�Z}[�g,
c��V�024^�A^�?x�B9r�B�VH�lmZ΃^L�a=�)����e�����ڮ��P��/;�u�c�llŠ��/z��0����k�|9ͻ����Ojƽ�څ^��x������R��}I�*U&�e�/�!�aa�8�C�׻�4�\c�Ʈ�9�B�b0�:������k�`�h�d��T��L�i�>x�������f�3�˝�c��T'�%s5��c�B�%�4��]��܉����s�t�&˭��.���o#am��ڞ�϶Ov]4�R�y���^/��l�V�O�c�p �����0�GW!pО���]��I�=\���2{��y�}�]�4-ڛn��0���e��~���>6R���5���{&�Z�gc�&B�f*�)I�;�ta�a�9Ðu���%��d���5}��m���NlJ�Ǧ��m��u�Q��}��vD;Nzx>9�M�x����K���������Z<++�x�\�[��e���!भ�Vz����F������U}�Wچ��l�p�13ꬭ�qdS\�ԡ�s�J)O���t�1�`c�So�t�Սw�p�ujPWN�qpv8l�5�r��XZ�ѹ(�7�\gJ�V��b�9�u��}s����3�:�vt��/��4f>��F���һ%�������m�Nۣ���]��U�A���AqI�e���{5��	oN�!�U*V"��E[`́��f�Z�������a�QrU,�۾�.4�45�giq tc/[}}��EK;���qK��nSmܝ�ܷx�
�L��ҥ�m|�����{FB,́�"]V�\b�v��Vd��i�3n�f�n���ZZAѠPj�*����S�F=����6eu3�� 3�.47��^��Z1<����'y$l�Qv�q[y$�p�Ms���j�y�-�(�4���v�9]�]�C ���\c;u�+?DoX�>l`�r��}$���Ff�V9x���2/T��J���&�j���+~�OE�6RlHS*^|-��������۱c7ܴS�w$C
��i�h�Zx�w�۫��]n���rw�m��g� �h��wvSeY{�fgR��s*�)�X�Wm_Q�yf�v��qd���,.w�*e�����ݵ�m�X�ZOm�����oL�s8�
Mée�C��b�.X��u_c�݃�sVNS�s0v�Yw5N�D�U� sF�j�v{_u�vʭ(U�N;`2.ؕ%�۾nX}�(��{;;��H�[S�]�4���\j#w���񏫘�]YnȘ�Ý{]��l��g�R������$���	v7D�&�{ɞ��Ev�M,Yht�/6�۽���Z$E�ݱ�����c��1��u�Ք�5�y�4�hN�z
ܥN{#x�1�� ��Un��D^����>��F���x��yS]a�+�pA�"�!���{Vۂ�-�$����ï9��N����}Kd������k���y֒��=��ŷ.�=�x�ŋ�&NJ�ц��V����C�ǹ�S�v�(��]=��|wl<��+�F>�ɋ-f���?�Uk��y�X�wƉ�U�:ˢ���V�d��Pyd�\��1�pp�G(���[���k+����ZO��	u�{.>�k���Pr��
6�K�7wxn�*��U�.�8��tgn.b��ł�[�ԥ	���H��9�}��Χ{��rQyQ��o��;6�``��oYۦHY��%u��vR��@ۤD�ki
��K�o��j�u��5rLW-ac	��l��ŗwtju��O�ޢ�[��"��O�9���ah*WRɰ	1Yʙ��x�gAA��a�lǭ�L�[Z��56U�!��¯c�+�Gr�N�:��ޤ�0sQ�$��t�b�T�F��W",sܰV�t�)k9���wep��T�%9�!>#6�=�]������a`,�/V�̏�gkD�ϺI��6֛�YC�;[v���Y�N�0^�F��pʕ�������p����Ǝ�V�'J��a%��/{Gh>�2h��:��rX�+�)|�k=����
��RȻI�L�o�q�N:x�t����3��7�Se���,qۉi-	*N�5�6x����).\�TQq�$P��]*��AE�UyUEQ���Ѥ'B���(Y8�s2e�E�ȋ��9�'-Z��G*8Qɖg.�L�b��8b7�J�T�T����\�p��	!��r��T$���qJ�hYQaY����B���^D���4��Z	p��qI�"NQP�V��q �G(AW���\��Uӑ�X��mh Y-��$�fN$�pZS�#ōS�P�i��R���$�4���8R�*��q�\'�f-*@�H��9i�(�,�
*���Ӑ�r"q�83%$Ƞ��+%T�6QF�&qUTuB�R��KVkN6�)����4vT.e�}���f�B��]c|Ga�X1�)w+�4ő%q�ܣՃ�)�W`��)��v�l~ ��L�{�;puL���B�Ž��5������{xJ�a{0��b+.K�����X���o����,Xz�oɛ�h��b7/Σ��+:	/n�f
�0�3ģ����v���ٰ7�T;յNy��ޜ����*y��t*fȍS�'�
`Ky~�=��A`��3J-c�mk�ڊ��qO�Y�H�[C�1��+p:&; �k�E_�K(r0��P��{��˫�d�ddf��`r����r@M������J��|�U"��֣Wp.���j&y̜���oH��ʯV ه��VbR6�c������� ����3�Z�s2��1����n&�¬�X:��l;�<͌�ۘ���n5P��Ů���mu��J�uy�^m����ڀ�CHT�n��gr�zxC�(�b�L�z�حu9T|�]D��O�� {�)m�;�:'����,�{#ܼJ鍩Iڮ����~L���Y��t���k�,�o7�4���؎�h���� �u�~���s'Ƙ�-�Ф��񲝳�]�U��G�ܝp���Ƌt�#z¢Ѽ�����ǹa�%�ԦU6�'�������� <<=s��H�v�N|:G;���uW�>̅�0��$[��&�CU=���$gU3|̨���J~3x��!�j���������ą{�\�=����펼O�{���~ru�	du��-K�}<nM�x�iq�=۸�{;]Nޞ����G_g\���4��v,��.]��ZOe%����=k׳�n̽ª���B>]R�͠��Ǟ�b��>t�iZbM�!t�}4�%u�'p��V��N��j���Ԗ�jY�7kR������f?E��{�_|'��%3;�H��Ic�)��;Bգ�5V�f��/Q�~LF�u`�#(��`�]����S���8���ZNwu��ٿT�Hk�=��u]��T9�(��!yuS+xHֺG��&��{�[)��u���#y	`tLt�#:ҽ��y^����~b�پ�:<�l�K|���)g#[�rD��w8�i�X;p���*���kM��i�{��
��[��Zu��ѵS��ĺB���r�u�>ڈǢä�hsE$��>wȆ�����9�����6���.<:��%u�͒����ꯩ��OU�����1��߹���oHx�¥�Z%r%R�JQ����^����]�W8ݥD1��%��K�V!����!��U�����158H���"���gw']�alؔ������X�����\�&Q���'���t�y2������Њ;BR�M�]B���Ҥb���l�|F�l���-&A�v�v�w�Wwӊ�.zj����^���[�|r7o_	�Q'T�����V;�j��pӡ[�ւ�=r0�yZRt�����Ъ�����x:�y�'��7�XǑ^�NE�x.������TV���z�W^l<�5g^�Y@w9v}o!��%]�K���,H�]+e�{�G�Ew'�� -�Yu����|��i��'������/:}A ߤ�Ѯr�ޕ�����p��:3C|��]�W�.V3���p�5O���4@r���^x�@�s3�Z҉t���k�9����H��=�uSWPk��I�鲲��b��C�2�b�1C�F�Y�`���e^�355`�]F�vGŝЖ7����iXf4]r�(�p�F�͑:�a�j8[w�>�F��y]l ��f�����ꪼ:�u�HeA��>P�O����̵���Uf׹�+�+��:�L���xh~�7=�f���X,ܷ��k���8�����Vđ���M�n�+�@���e��Z�I��fo�j����e�m��Y�1H����i<�/�]��W�͝�,qE��X��ޘ��&�S;{�f�i%�>��l��F��cl3'���C|���������<ݾx�a�+)�p�KnVr��E��	�e�a�~�DN�=<i�ujy�Zm7�2;j�X��y����(�1�x�["��f�����K���V�M#4e��iv���1ݩ���ظ��A]�An
��H_sU]�HZ�޷���넲.�cW(m%�5E��I������o���*yle�6Z�1��iL�,��4<^�O�t����C�'�e���-ږ����ޒ(��5+�S�[���JT|�1�-+͊NI�K;��Y&ݑx��r'$�[���`��C�ϰ�<�E���ׂwҁ��F�f�/�5�,��o���+��|�k�Xx�7�a�vTX۷u���{�|U����'fV��\��n�ӣxr��o������Iozu�[7?z;Vd>''۫F��Ȇzap�y\X�s>�_��&C���n���+e�ZNL���y˰�[�����F�a-�&��ں��<�W�.x>�ѡn_��������6�p��G&��s��X�|!�	��Jo*z�K�]d��2�r�+�~�r�
��}����7iT�\$ު(vDB;,J�bJ��.��u�ȣa�W�����{6ac�<�br�o{z`�my�=�Fp�ͳ��츻�w�`�Z�I����l�z�ũ���'ݖ���g�)��-�dٲ�	ݰ�4�Ӳ{ܸ���	l�G�W��]w��0�M!|����8�ͨ�Am����"g��ogy�/v��(��!{iuN�<���{9�)y���Ϸ��[��{�f��䯸�%p��z��y/�:��L`4��A���<�ŋ�!��ף��&�Z7g��U�����ƭ���0�Ƞ��0*^Vˌ�����{]�1�fHH���\fiوcϷ�����pz� ��$/��h�7�7&�'w���8���X��.Ɯ;
L�j�T������x�BVʎQn����ť���㍘|\JS}a��S՜�����92��fo,��xj�~�L��<��
����������r��3yU��v�M�D�+�bݲ*�j���l�+�
wk~t���%�x,���m�=�����,T�K]��º��Ou���=�&2��k����Gw��&T�[̆��u�P�f\sN�{���[b�;��=�i*����[Yn��s�Q�b��F������襯�����R��h�U�:-_NY��7v�+���F��ԨOc~:nM�x�}K�hT 7*p,�|�q�)�Rf˃��2v�CA�D<o��Y������4�k��{��eW��ݒ���^y�#T'��"���,�
u���F��LG���.=t��	�7ᄫVޭ��S��.�bީ�������Tc( ז�%�SWu���(g�[�OQvs�ǽm�S��ᕧ�+�pe�Wr	���}M�M��[� U�A����S0Q)��<������!L��k���9���7ԛ4��q؆ӣ�8<#�۵ �'���P�b�	ی��*���ꪯ��2�t�{}��M[��{.-�.'ǝ�Wy���w�?9�=Y=-Fs��9e���oa��{:��f���bP��+,e�1Ѳ�w���12��F�lN���qv]ɻ^���fy�n��l�,�s���Q�ɚ�*�������j�A���`�Qcg/��cD�&���x[���<˞,��Ե���rg��ߧF9�O3��kO�=����l�v����PD��*.�ފ9씳z�Ua���7=�͞�B7��I�`[t^j.)��%��qO9K�S�Kb'��𷒂�т�-�Xiu�^���A����X:��ΊA+�OƯ{���	_���NB]bh�+����]}�oMu�Y��\ip��|�\�i6�(�n�DT jWHꣾ�o���&8�T�1��+4{�Jo֛�Z��Й�� P���5�XtR��=
�g�kd�O�Z ���	G��7�O�5Z*7]D���� \��V�P��1`󂻴��M�|ҩ��f�������0wnr�^+�e�ǣ&��
5D1�#�gwRT���;!���F����if��W(�3�����W�Mv��]��@ɏ���pCTn�U��c�mhO�s9x.�x�.�+��][�b��w2bk��H���s�~o��4`U�����\�NeEB�zuVj�U�a�5��la�Bْ���w��8�m���1#U��xydmk�ڶ!`��T==6�������N���Тվ�ˇ{�%js9ݢF{�˔�GX�}��w��Yg_�d�o���ɞv}�L|J��]��h�cK<��`������كcX�.c��Yc��EӾ�����k�l��cH.���VӞ~��nW���W��<C^���KhYn�ĥ��X��')��w�x�]K������yy�o�����\iM���~<����B;o�6������!;�-��Sg��^n�L+���o_a���Ʌ�~�:����
��߈��zy������`�����g)rߎd,V���*\Pj��t��sNh�z��kF8w{D�P�*���ǡP�����>�T1���I�>U�z\'&�n�t]��p�E���镦�m\��2a�{��:�W��&�[X�6��;��������GҎd���7#�NsR}�UUn7'i^���3��tq+�=�RpV
�-�Y�I�V���]��v-R��7�rE��R����a��X�t�-�

� ���$b�N�6!-ƹkE�I��5*��m,�n�3|���8�Xd$8,����a���Y{�׋�4O��q4�f�}��/9;
iڛ�n��Ș�[��jzX��w'N�͞�jU���mܡ�]���}�gc�����ʕ]nVe%�Fp[s��a���j�'Դ���
��r������6����u�]<��Sc{C�nE�Ж�,#:�3E�=9F����މL�z��E>Jn�h>Sa�,S���}�6��	X�S�T�C�����=xU���j����9��ʾ�vI��]Z��ɍ�V���׻��U�s�b����Lnn�ڶ���%��uKT��4`ޱ�P��N���4OgOH�}�r^��9���)~�/*���2�*�]g�)ϒ��xjV�ՙ�)����k��	�f��Ec\��N�0�J�U��.�\#�)S��k|3;�ғF�N)v��\lt���g=7����rs�}�';�3
}(<�:���o~����;�����^ٟ�{�~-���iw����o>c=�U���d�mE.�Z;�z�o\S-��N����z���Pǣ]&��C��,����d�z�Gsf���V��Lm����tLv
G$��]��+�ef�H�e�������Vk������Sk�w	XT�vX&��%aR�zk�=��3I�Y������޹A4֗�l*�5���ĭU��l](��<�J9O���rW��oӥS��o��/ہ66�<�Ѱ��,<��;w6���[ݡ��>�DQᖹ*º�l��]�
w`�v�V`�"�ʭw�ޛv������TQcdoXr���!.�1s%w_w,��~ljM���]��;�\�l�R�"_��f�+�%P5)��B�5����o��F�� ����zK%8gc��W�"�R�c�5�Xk�ik8/�%節wz�_iM�Q�U΃t�L�X�[���*�0�Q���XJ)�U,m�` TVK,�*��E�Yk��dyث!�Iچ���pp��1^{�<����+e ʳH�1���j D��$��/��pC�q������;ո�S#q'݋�p�nD�M)���ڣ�5�7uq�,�"�����3�k�H�����e�l���Ń��.R�&�����ެv]�C�n;�z���l���ۧ���Cu�ucf0"�zk0�=�.�L�2ݷڹ��yr���黜(P}]�\�sE4�k�8�ޢ�Mz��]���1�X,Dq�J�>o�/ЛD[��ǖ�ީJ]�t.��{"`���܎5��YI������E����4L
��ܢYV#~Ε�������LOndVV����<K�P��]�O]^S��Z�N
�#�l�r� ��y`?<CxNd�y;b���-f5���з���O��fУ9�y�ue��J�Y��	OVc��X�P�X�������K1��n��U$²u�K���y�h�8Z�N����Y8E�7Y�U��Gw_��^uZ�CWr�Z�����WE�2���w�F��gZ쥳f��Z\z�4P޽�\x��c��|���
X��vq`mn�
�%RZV6n0��/&��]Zk*-�1��eA	� (V�b�#`k��c+A����4��}�x�e�3k�[/����S�sor[tWa���-|����W��W��E��;��ӻ�F�P�0$�F#:�S\ح �r��kA�ˆ\����2VJ�/��B��1�XY=�y7���3Qr`F�H�8��F�ea�uիF�f4q�	�o���# \�+zCWDF�:��eꙵ(���yMxAF����� �����u�a����[��J�#��*齀��f�n��W/a�]��]��f�V�wc���Zp���t��Sl�.��N�H��ċk�2��\mk깐`b\}���mh��]��`�6�+��ld���R2����U��t�G� O�!���݁�*Ռ�*tφ�/m�֢#��6UpU�݅�w9ZSo��nWw����h#r����[m�d��yB��be�&�j�K�����j�+�`_,i�zY'hJ�ߜ�[dR V; �qV����P�c�J+CU���+VJ�c�.ax�$8�L;Öq���\�4�n�fR�歂���<�6����D�P�Y{]�)�+|쬼uu�XV�\��e#�8Վ^��;uLdA���(T��U:6V��fl[p��^�M��ε�8 B#Z�bY��4�b���^������`z�e����s�%�R|��Ŗ%E�\m�f���a�珖��9xb�Yհ<Z0�[/,�r���K�-�Bl	4W9����+���R���Wt�Hܣ6���צ�������;��߯{���yr>����a:�^BD*�� �$QN-d��p�k,头�2*I2�0�.�Jp��ek������%K�j�*����в���B5��ar��rT�3P�"��I�R6��g%eʺK:r�Z$E",��EA�7^
O�S�TPN�n<�N�CVTI�i#�t�#2#2B
BJ
�6�4�3�RC�NDT��I�ҡ,��X�- �(TvQG���+��9B��eDr���*��t�
�T�H5**,�%R
��AI����qЧ)�d���9
\`�6�V"#��f����d,��U\IA%P�
�KK�DDh��$�EC4"Q�s�E���5*,s���9�r��JЋ��B+�*�*���%fI%5ds0L��%:A�$�U�9V�QVHQfE�� ��r'.�"drI5dBP�J�Q9����Q㘑QTT�(��-}�<F�=�����kŽ�. �)l�q�w;6��P����7�mP��zC�mq`�8�uM��)
+�Ӯ������q	'4n�_糓X%���7/�[y�8'��h��'�yM���C��/��ly���f��6����z�ʰ0�5Nv8U>�ˢ0��ۊ�,Zp��f�.�Y��p�U�h5L#�����6��}��3�m�[�F���jؒ�K1��c��N�ϗf��u�^u�	�RZ����&�1�G*�2���lC���3ΰ<����2�w;gC�ӥ�kY&�:��.����Խ���'\bM��3�5��P��`�}}Z�����e�g���ը�y.�$��O=#�|�.w=��˼گ����Esk����J�編��*?V;�w7:)��ټ��d�[���M���@*���;FG%��g�ɾ./�vH��%�X5�N
�"����c%s�h���}����c�"d��
��U�ڋ�v���f4����YӪ�3�Uf%|���ж�X#��L�V	�մ��_Õ� !W17E-�5��{�t:��6a�e�<�k=��5���ԭ��W�է���N"���,�üÚS�ͱ�.{����s7<0�O��_UhJ�<(ff����Flm$([�Ɨ_��]��!⦴���^�n=���)a�z�瓾���.���K��h�\�i���bI��/�9�l��X�,t���K���a�OW��c���4n�_v�U��T�{�^���-}a�;	1���SҬC���(��ۛx"�v����sv��۹�6N���V�Q�;�ЬcȫT�:�MLK�6�vojM6�68f�Mؑ]���B��Ξ&���n�vB7M�Y}�Y2��e�S�`Co&z.W�[��ٚ(���׻�S��x(Q�������-�7�|��:��Uc�C�^Jܪ�]>ܛf�c��F&�Nv.��c��Z�����fu��Pv�T9x����z�r�\y__����X*��e���<�eMR߽��hTK��#�������v�77���m�!���Au�@�����b;YAթ���_����ʳ�+/5���jŕ�=�7�3Ej��¡#9�� �ϼ,ף�О��V�_o�_V��2�EE�B����Z{����%��kk� .��S:^�����i�C*�2�v롦��ݷ�N��`|%�xj��S���j���UUm%ی�q��3�x�{P=���=}S]�ڮ�)&�����V ����}o�m�b��G'�y��US]Y�(���_^�U+��}O{Q��Q@��Y�H���ؕ��r�7���Ꝯg9�=����^x��r�n�㾯,��z[{��W(��M�V2y_�_=R�b[���>�~O��_�������vlDj0���RpV	��B�%�p�r�	��%W:����F�[����U�����a�G�Nٙ2����7�lT�7ګ�-�|�Z��bN���	����Y/����̫�T�zwV`��x��բS�i��,�o
#{���٭�)��Q9��L �#z�r6+����0B�sНv갫[�!����e=��Շ7��d���j��h5�$3W� R�pBd�����-���f3��C�L��52r=Ŝ��-�
)�Ϟ*�o�����z�j�>q
Ș*R�v�s�T��7�E�>�g:U:�^}�u�Žuu����|1R��Ɯɽ��k����Z�S ���]�E�I�ӿUUU7�b�[��I���u�zZ!`x'ԋ�~��)e�|/���X��K)N^K4⚁�S�����7�CL>Sa�,ӎ��}�K��seBZ3mA,#����4���ɝ��؜�`o\+���w����k�a��V�К�Eͅ4zV���u��v���bh$���L0�=i���F��;[P��AY�3R�v��3bN���~�F�Of�	�e���)�k*�6:�۝q�ϗ$�~^�O�2Ԍ6$���{V��z�i(Z��vж{��[|3�wwe0}|�l=1�9��E\5���.��T�=̴�v�`�>�׵�g.�S'�n�h��u�L$�2;E��\S�f������J�N6�\�0��J���SM��[��s}���ՉI��x�]���&R%�pv��kg'���CS�a��U���!m���N����G�v:u��s��ۅ������:D���W2��K�Z:E��J�MH���<�+o�}�� `Z�%[�������Y���n��ؾ��n�ӹ��ʡ�Q
�ܑ^�hL�ս�7�����74V��\T{fT�zS���S����=e�#gzru��Q���k'Q�=�~��6y��5�趹z��On�T����%�su;��B�tl���yΆ�T�%�qs%w^�)�q�Z�J�+Re��җw��e'��hv��t�g���#~���Y��x�Z.62��O�o6�f�Iƫ�0�BL%B��XS�)8j�����)k'f�t�d��;�Ӽ`��vX���k�]o<�s7q].C���1�+�k���b���]��+�_�I���;xe�ӛ�&��c]�ri��UU�NZ����:�6M�%_�l׋.�Y��p�UC�A�yUcK,��^kc�b�\��ש����p/G'eK�<�}y�u���ڏ�h"K��n�F6���7��E�~U|Y0�;���и���+���oځ�Nњ�3���P^�9���a�iy!��=Vυ�+���>}T%�f�;��U�
�֞J�x�Jͩ��Z�)4�����fۺ��S�/�lO'���%��=As�r'���Z�e͕x�A�ͻ\��o#�����2��TL��Z+�\�����2)(�؞	�etN�Q���o���ՐԙPu;��������=�z�: b��U_l{$��V(���)<9c���X}�V�����*�s����z�CrP}ڏ���=�ާҕ��V�å
�� <ݶ��~D�T����+8lb��|��b�D=q�.s;yh�|�em�͜������b.�Up7�8K%ꋏ�����w��p�8{}>ΝO�_������ܞ8��%Oc���-v9�Zؕʐ[��RC�H����S�e�#v��v��qx\#R�]S�{[ݟ0�C�!S�B�nU	+6t�uY֚�y���K�j"F[���iX��,f�v�g��V����n��s�M��̼O���ͪ��U�_P��aV������_9���eww�׬���>�B��_r�����#~�Wz6���79����>VR�^Q��.�E���e��ÈW��f�E�oX�k7��l�|W۾>~��J����CA��7מ�}Z����PJ/�B�l��ӻ�
eڲyq��h���5��;�앫� ���^����W��cU��<��2��k4^d�<�we*+����Č4n��'��]� x-�q��Q��x��ʕ���UfG�� �Y�:�ju����M�ܝ�~0������.ܛF��
ْQucQ�ݱt����{ڒ���l���z��C<� չUR��g+�<
1)��J���O�3��>��'l'E�"*���_�Z˃�/֪w���Xh�3>��X���e1�bh�G��<�%z�����y3so�(kK�YB�b%�����g���A�d�xh�(z���B������d��A%�;�m��~�=��ǻ�V�g�,��^=�(cj��u
�mW&�=��!�y���s���y'�~o�RV��\c�R5��YﱎW�oSf��p�\+�Z���)z�-~�[���3�Cγ������DN�==���Tw%'G'�XR���*���<�H֛�-��o��ζ_W��9D��]0����BZj�{-Y�5q(=<��6���-�r��5Ԑח�Cl�bعY��BċO����c��EX�9/#]�����N�(|�tF�L��4-���7hI�[���3�4hE�X��AQ�q���3���5�6����!}����7})K͵~K#~C�@�7�(B9�VVU�� �Q>��ܭt��'2����.��w�X�j���ej����-�c�K=���_n�t݁3��e�ra�/��zyn���BWS����ـB�
��[)�7�	��R�E�<�p=��eHx���J�F몄-y����'C�U���[M^t޳�n�i[iWm<��M��`2r"�_�<��4��'=�W5�;�
�%�Ǵ��qU4�޷��s�V��Z�"8-=6��p���&*rw��}����j�r�엁8���x*��B�A7�3�{_�Ι��Wxio��7��13������&�~t7��uKm	;�t^�g�l�~u�K��߅�I���ɵ[5������ױ4P��o ]�LcQ��;,T���#^�L��Z�����7%���xh�)�ޡ#ݖ��=brE�X��
3�O\�~2������EjxΝ��Y�=c]��2S��u�T�r �u�����.
���� ն#��D]K˯��Uwq�Q�"���j���qP���6�=eQF�}�8뮯����w١a�9��i��X�{NN�����u�j��)�hҽ�ݺ��-�"n%OF�:R�ZV�{�3݇XB��7�����l���!�^Į�Y��pߕ׽�ġ��ūv����#F���Q�Ӌ��^n�h��ՙ�*&;=Xk�[��ۮ�y謙Iy�~}�#j�%=���|��=^��M>+��V��2_aqJysd.��a��;L�V
|)�Z��FcS�a�M��{1].�,n��w{�򲢵�n��P[��)!W��`uet.� ��W]�vE�&���q9i��?C�{\5�o��ݵ���/o�\��Ȯ���K93zG�<gU_vtŪK�J`)=��2E;Smҗ�BW��Tϡ=avZ������sn�vky�gc�6
�� U��8j�j;Y,=�
��t�ԯ1��֢F��{ys�Md�Z�����J\��-�ˌ��u����O�c�$L0)#Vy��t�G����{��9J��R�b�[5֚� �	Wiȯ&^�ͬ�9No>4�k���W�Gj+	��:�K���"-�c�[���HcV�2�1[ni�-���Jڼ�Wi�tv�!T���NԞ.8��wn�mv��"��+�b��岬��-p�n�	K5�7}��5=N�o�YwS�8�r�qn�1�jֱW"wFo(�Us���;J}*�L|*�ܛF��]��(��f��땰o�z�Ƀo�����8F�Ok���nc��}�O/1o��ձ:N���|�������xB�A�u�� [tZ���#o���rV^2�a�~)����M�{�y��ޖ��z�3ܧ�z�>}��̓^Vs��m����~8�����Ã�U�tUr���L ���(v5�k�zM�C3k�[�!���O*�!lU!�����|)ْ��Iv
^�:P�we���m��c��̾�����n��I�:���+����ȅ�����l瞦�����bb	��ț��n��T��SGu���)�X$V�y<�%s�X�ѩ����	�C��wٮ���S��?np��,���b�%�+D�H[���R�2�����w���B3-L�~���Ňۀ=Z���Ӑ�	Xr���1Q�������cw�t:1١����i4W+X��=��"N��/3�ֲ&�A��+�t��P�s2�M��)CO�t�l\w��Ņ�9p���Ί<�z�DGj�orK�25z`خ�9[F�Y�=D�4�ٜ7^Q*V䔝������j㸕�:pNQ�C���#�ח7�f��֮�����}�q�<O�dڂ�v���j��];�;��T}�yd9׌�icTF�8>"� g�o�{/��F�5�փu���e���Q�-mv=�2�*?fM4��)H��,1�p�N=��ASZz��)� �y�ﳡ�5P:a[V����	���ɤmjݎ�6��8,㸉��+����v�\+��hΐn}6m�ʾ�}r��X�+&T�{��]^H�U�v�cZ����:��W�ӇJCP�$����!�;yƈٺ
t��޾ݲ�V�
�A81ϝ��kj*i���'�0.ޫl�H��A��CXv-�vg}k��k�`�ԎS�;����Ϭr���u:��t�B����=�EiJ�_;�AGuiIz�swX�T�4�;�emn�Z:�	�̠�晕nn��"�;�5+)�pgɰ݇�����]���U�P�,!g~�;uٽM5�����+�7(�\�԰��B�qM˕�����mV�B�����EG�Z;�G0�8��]1��m������Nc��2�Tv@^˛�`�'VfQ��z�FS���2=�731�0��k-�WN��(3�=|��ڂ��,�c��=ia�{��å���:���'!|�]I�n��
�*����"5���D�m�T5+.��R�15#�2I�Gs:�ʧa�3�N�[�����y������\CA;����x��=f�;uư��O��-�WaS� �6���Tp���u�"��2Tŵ9�	[��5��7��M�����<�'~sV�	G;�ޞ�(�0�����_k�l���������}�l�J���&b>��"ƮMP�N�S��#n�t��!�� ���{����61�'&�(s�Y��ټY���J4���W�ׁLuvw�d�p0&���*R+%WLv�m87�-�(K���neA���ۇh3oI��#��u՘�-�[��b����s��*;N�]�I�c�KE�����[�ߣ�5�Q��Ĵ��9j�ɶ2]��Rm��Y��9��S������4�(r���ʂollT�RW�Ӕq��N����S@�����X��:\�ɏLΣrvs:�Aj�+혐�@��3t����8�4�z(H9ʘ����`ن�o^L"�*z ��+-�o4Vo*�ӑ�y1QJ�̗L濻�nPI�3}ؾ�o��=i��V��m�����	�	s�V�qփ����0�_��[�f�gr5�5p��֩3�laQ�(������ùw$���� �y�U˔2���X��c���!Q� �y+�tq,��쥍��-ɝ��߲*"���:r�ED�#"���(J�9E*\��i!����A�0��EiT�d%d!�l�����IB�a\��EGSA$!-��rq��TF(�K2 ���E9ZЙ*	�Ҫ����\��*�(�"��E"�AU�r9T�9��"(*�&�*�*���ED��eq�UW.jM�#�Er��$�"g*��*,��ȹr"*�I%Mj���#�Ȃ�Q2�<���*���!Q8M2�Nr"�9%c(�J$��DP�UE\�]D��AuB**���+�˔p�����ʇ��ʪ
�)j�A�H#�t�UD$��#�DAA��r�Yp��&R�ˑr��2EB�˪FdD
�����*�" ѥW*(��șQUL��
�*"���ӥG+�C�H�JW����p��%Y��X�9±BLԵ),q✊�
�L��!*�D�8�DQAB�
!����|(+p�3z�8qQ�����+���ڸ�5�.��!�5/���SFe1�=��)a�j�u�m�j-� ������j��2���)P��y�ҲƤX��,e�`%^���ֹEὑΓڔ'J�%���W���k����/�����y��p�js�Mr0<ڥ
�k�(��ѐ��ϕt&����M�.:�aT�a�hs�.�a��J�˔
x>9�ո�)i��:!ew9w��[���OT_N���]p�1�o7��X6�l�Yn��y���F�«fh���B�X����l�ud��ji��ݲ�h��wE�ʬ�}�6͌%^9�݃����]O�-�^�Clz���x��~��t�S�c�*����9k?Ve��e=n;��:�3�뉯x�>��u0>S�Zܬd�b7"Ԛ�zsk�y)��~�_�ua�%��m!Y؅�����fog*�L��<���y���㋙�o|b�W�ʃ�\|���<�溕l�� X>[��U+6!�V5����c��D���� �W*;}�����@9�g.���Xp���MΰӶ�q��iՈb��4���HǛ�g[��#�F@'��Rz/�~���%a��x���7�q��%�7YM���:/����J������<���s9|;��������}���g�-�Es|��5�F:V�j�K�c��(�6&�4�w��j��V-�֛�\�>1ܴJ�vV	�j���@�Y��M�֚NU,�)ƦSO��-U�An8�AW�YM�p�WNpȦ�Vs��ײv�2�/^u0�$�.85C�±��O*�q�a{R���0��O����7�mv�@�k����gx�_Z�EW���X�� �\Oi�r<v!;w?#W�fpLg�L�5�77��;*5��n	�.�G
�y�x����ʅו���|���//AQ��B2�u�ic�;~:�{���J�^�,�;�M�Y7�B�����\s<&5�P����h�TJ��wy��V�6����h=�� 
���"�U)"���2���ǪQJwx�a�����o�4���foL�j�{yM��&���̤\�t��N����"�d�\�!�tC�O	�U>�[{��sO$�o��|V���|���6�=��T���|�ӓ�}R��!>u$p�5�3��?;ɑ�����"�ti-̧�[B�"��7����t�s�ݎvuJJ��a��<}C%`�����00�ځ��V%����;�;Y�k8�=SpZ��;�IS��F6��\���9�:�W(\�p��P�5����F�Y(_غ��6�NJ�q<�?Fน�+t�O<���v�v_T�w�N�v߫0ø�e=7�t�� ���lyuT�.!�);wBees��|+Һe�!���I��Tx��T/�=�W��xS;;(��V �N��.�"��ՙ��G-f��_
��o2�>�BM\��|/�"rP�ǫ.:�/�o�(s*`ǝ>b�����7��o��q�
~u��cw���\U��z/�T���YXz*�ʈ���ړ�zO�mk��7�d����頷��Oԙzs���-ի��koQ�a�R6�V��ܦ"�����t��^'���ⴑ�%�ǡ5Mw/B���ye����N���݇/��=��������m��W����Y�O#�P�گ�;��F}���}	�ZuE���]V����<]��B��z�?O����Q�-��#/���jV}�yK����)
��^�^{�ܟ�wӐ�b�0W�۶=>���	M����������+��T�������yU���U��-��q��#�T�~�7��V�kYK��ٍ���+������I�nMa��<^ܻ�'�k��7@�*""���M�4�c�K�ɩZ�)�_-����/�i��3]���SZ�k2I�����!ؓ;�t�eG2�w �j����R!w�ckb牧�+�-9�.7'E�W!��%v#f#�S"J������b��-�f�K9���Bh����^�C�U���I��7#
�#"�R��Ѹ0x,z�J^�[�ꡱHצv����v�_�����;+x=���u]nc��s���X�?\z�M9 .�a��-�zLgvs���:��3/�V��YF�����HglԔ2�)�{>���	*`9�]^�4��]vo�5�../�WuT���zs�ǝl��+���coX�/UQg#7���r��gC�����M0=mMP�>/(
���>s,vo�l<>�L-�e=7V�90����,>���xq��Zb��{��b��z�(���q��4"L���x�������KX���
״��t9�.0���9Mk {�|�t�c̸��o,Ḏ,��q��˜�<[Է�v�UdoL۵~��(Q�{�\t�7�9ӡ��Ր=�����ꍸ{�t�?�5bI�#6�}ܼ�(�-�����><,�iq�@ŲC������S����kw\2j�}��>��ڐs�֋����ҳZ1���ƥn�X��R�E�c������q�7E���%(c���d�w���m��:Z�U�J�/6�WJ�hE�`\
��>c���m�S�e��t�H�1B�n�l��	��B��n��׹Y㕶��M����<v���p���$\�x����{R���8��c�FԄ6�;xu򦎭�1�·n��V��;��/��Z=���13Ǥ�]*&��LV���y��(s:�a]^�$���)^�碽�f^���)��lh�U}h{��Q�Ct$e �v(�	��\�R�oٽ�x����tɆ�a{�\I�]� ���Oiq�K�q�uZ=�@�j� ���G���{�2>���י�3Ua��85�u�`W��c�����q��n���~�EdĤuҌz��������0�V���ꈙ�+�3��Dd��{Z®�erx�L�U}n}q"�V5P��sݜp��8N"  �3���-��Į9��(:��,_ʶ�|VS�{Ccy�����xo�,� '��z�<j蕧:d�������Q��)��0��Gs4å��<!���E{N,;~{=�Z���/��� .���\���am���߲�U���5VD�Y���������uG�!��Vj:�m�ٸmP��UW���z�-K%^�sLv�E�g��$��s`��7�5��쎻ن��F98�W҅K�sc�
nK�G*��+����j��y�[X.O�P=-	Q+O��7y�HT��΋��:�� qD�y����b��:V�]�gh�{�D� 3:ݴNf�ˆnH8r.1�Bk��^ν���	{(a��<;~뻅k���[�:mk���=����������:�d�dԮ��������j�W'��k��9�_ޜ��Jk)=��{�Տ�=�>�;7�*��yg����}�9��nZ����Ƿف���0�}RY��r�}�zX�d��R=�g�������)䎘�	�����;t!�����'�����ت��^��Wu�o����1����=1!u^M/z��^q�-�Mj��_��
�q2�;�uX0��C��W��>"U��:޿t��Y��.t�C�=������=��t�J�=��h
Ḧ́o�^��/-�ǁL��_����zn�ϲ�,�%.5MT��9L�8�/M«���(�Dc�)*@YW�؇�ͭ��rs�����O����r��.=3�_��¸+�b�]��$��V���fpF	8=2�ތ�U�>�C�6T���G�e"}}<ʯe!���1��!����@b�d�l��|j���1���<�쿧x�,5:N�YqU#�O:�}�T.���J)�q?Dre��j�~�l�V��ُ��w��w�.QJ�4]p��ѽ:�p�3��]��9�lJ҉�?`�Ez�+��bf1������_�b��P�̽�th��e2�R7�4��$`����#WqY6�@�)B�}I����e���ʹ����͞�(D{��Br��w��^��l���W"ӧ7�d57��&릅��@\}�0����[Y�dϋ̴}��3��(���Q|tN� �^�Z�RE�A�-t����?����O�>���AC��DSFa��E|T�\�D�P�����q=@.;�C����]��叆�*���<Le�ϱ����[�肯/���YK���;6��+�)��%Q�&����4
M���~�u?;�a�l��Ǎ,���p����(b�.��mP���41�Ƿ���y봵饾+{�,���'|nJ㾝�{��[짦�\�3Q���n��%w,��F�U=�R�y�)Fl[�~�m��LX��B�˙�8}F�3�/�,;u��
Q< �d"!�E��R�r��dO� ��j���>�'M�<ˑ|�
���:s�DK=T�x\��J�?������Q~N�@M�3�˗R�\-������}ߡ��_\o����腒FḇӀ��T����@��_Y�^{0z�?
]ƜGL�1x�r�?dj~`��L�g0�}Q��Y�k'	H��ʀ)�Wf���g/ߺ���G���0�O@�Vm�H��-�`����Q��P�\�R5��ֵ�GN���u��v}K�nي�@w_Ϩr��˹�\:�����I=�S/@�CuK�F�����_���pA*���hˮ��2cy�z�hk�m�W���^�.#�8��e�^ّ�v�,>R����f���z�P�\�B�Mg�b���(z_Ⴛ�O��*�h���jw�瑿L��eY@bu��i�ڸ�z>�d��7�!,��8�����|���vn�o�j=��=}<ʬ�\z�T/U�+��2B�/Ѿz��+W�<��8�>�9Ӧ.z�eρ��� ����TJW�ߥqx����Kc>��z����*aǼ^'P�Z����q�|�N
�v�@���J�@H�'�?ne�[���=Ь_��Z�y�4�7Ϩ��o%�W�P��6x��'���GK��S*H�sѸ��g ��uyoc���:�6K��u�����y��z��~�s.%Ϡu��X�DBYː���צ��:���I�D�;麎��2biue�R�����2��7#{}��9.��O{���b���a��
�}�7��&_������
��d�X]d��BP;P��3�8�֔��q�p�״�9�d/Ht�C�c��7��I������= �|��
-]��ձ�y��YF�����k�8�'YWg˃�w�W�,tk�g��'�OȞ~z� �,�\�Ϭ��nq�2�nV����eX��[�M�#D<�DY:Z�����n9����V{0�
��M��t*�!X�ۣۋz�n&'h")�\܊?�����$o�D?}����]�2=���~GX�q'��Q��B�ΰ.��؞�77�ӳX�\�u�����T�����ƞ{ֽ�r��@��S��e��7�p�gg�aО��Ja`�uX6�^��}�1:�{���zX�8��(��^�ޗ�8�[���J�Q����يYۙ�i�w%j[s����:��L{�p��zg�R+ڐ��- ;�/��?V��˓C	��u�轪�����\9���x��	H�:��{�P��{���L�>%�Y$!����#t�;�q�����s��e�˞����ѐ�+�b�*{�S���j<k�Y3�ߦP�\+��<�wr�mk�2a_�s�Jw�|�2��ֆ������rQ�n����N��I\�u���ܠz�7�O�w����A��f@�]���3�|�V��^v���� .)ʠ�!��nE����^9r�y��x,6WFJ_^m�I:l���.!��4�\(w*�ރe��c��ߪ��ޝ�Z_�.�F���!f�d����)�g�y:zV=ޮ�\�^����ye���;��*�w��[��W"rj�r��v"��X��E�)u�V`�����aJ�c�HA��xGg^�j��[�Y]Ef�u;��x�+G[[�*T�к�Sw)�s.��ڣ|�e�N;N�n�ن`=IwL�.6�L%ލ�e�[��=��rT�Z*:)�Uq1Ke��+�d�N�bҾ�Q���_�u�K��-B�Y���u`o��t����	N�&@Xjؘ���|9��^=r���/*]oWn)�O��.���[>-P��� �o,
�z��=Lv��6��Q
��\{�w�5֡��>�yF��];��}f��:�6�;x��UX��_-�%U�sLwM�"�^���t�sճ��ǡ8ݤ&�xa���è�{��/B�sTT��?|Q���B+��_�?~J��O���-`�\c\��S��0��N
�q�X3Q������Cʵ��V���L��^�_�nG8�{�G9fu3f[��/��"r�{������x�w����Z \o=��h����������_���5����F%~�>̯qezR����v�>����&�tU��llU�����j��V�hu�*����љ%�u\0��C��^'���()����yT˘g���m[���g�!��t�s��}C�\-�)Z���9n����q[����j.L³��y;.��{%*j19�]h7����@��բɋ1�=�#���CN7�YWP�Z���.hȺ�VvNyqnT�}\!,���e
0����@�Xt�ei�o�j:���pӜ�׬���)�P��8ݔ��U�6��	3R�Zo��gҮ�����Oĵ���T�����dN��Oq+{�49$����2�����n���w*�Θ�.g������r���ӼT���پ�Na}1Ty�M�)��Gn�eow�R��ܑ���ld��nEiU�ʗ¬'Ƣ��Kt��.���N9�;Ře:O���N��/�)��Ŷ�����'	k�A��������U�/A��ǘ�:��R� �o7�m\������In�ԵX�
�i����a0�u�8����Թu-��%���I�Բ�����u��<��h*صP��onf:���T���6Tu�Բd����ma} MU��v�R.��"��]�������n�>wn��^���@������;r� ��J:)�+-*�ٕt{�D<k�ւ��F/�^�����ۦ*�Pc�]ƄC�ƍfq�˨+��)��z��n�0����r��(�=Lg�����je�l�殰V�{&vc";�R�L��&�A8�]&sܿ��,&�t��Ft��5�Υ���Q��>���&]EΕ��V𻂯�.�̗��m���@^���H>��=(�lw�a�k�tC\��4�=��n�u(��Hin�X�7E$��Yi�2\�__L۵۰uV��E��Kh��kfY������U/f�>�cn�aRAXa!Y9��ً4�܌^[X�qAyQ�����edE��G4�]\���%
7[f�O.�5����m�mO�闕�����v5�(-��MlR:;��Fm^9��<��\Ҫ�A+MfvmvJ�@wV��v�6Z�z9�i���*�*Q�)*���u�VZg�gi��+�z�6_�Τk��ҪV:R�ܴ9*�
������2)�?·��ꮖj� ��jlɒ���6����	@V�m�Ė�0(���ݭ�7�p�2����	t�Lk(ձL�gwi�\�Qq�)�_w|4�O�t�B����!���+!�>�綔�N=]([�Z��(!�n⦟g��\��HfY�9FC˽�Ռ��0])|��S0�zG ��u�j�ӡr���V���3�Z����K�m��������>�#��.����K��ۙك� �t�ZAg^7�9�i��. f˶>���� do"�a�j��2t��xr�j�f^��Y�E�o̅m�d�A�I���[2�`�Aw^��eG�����;ŎW�¯^WV�5�L��NLU���ʶ��bG�`3�)qj�YY
â�[}b�����& +'$�M���FX!�M�j�����a3�QD��y�Nh�\��7%��\h��wT�O����றՖ�&6v5R�umt:ͪ�kfs�Ԩ|(P����kY�DVds4�ȫH�r�<."��.�t�I�TEEF����%u�J��Eӥ\�+�.�V��^$�,�$9Ts$��Q ��3��\�\�P�P��*��ʩR�4J�TZĈ��EU�%��)2�	Z���m):\�9\U�$�H��\t��:QTTr"���rͭȴ��B"�D*\�#S�A�8�*2J��<,�D�*
"���)Q��s�Qr���g,�R
 �(�%49ʮr��qD\�/$DTQ��A�P�"�� ��f�AEQUS��
��G*�*����8�\�B#:�H�TΪ�D��Ur�"H,�$�UUW*�&]� ��YUZ�p�j�a�*��%��Q�9�G*.wp��aI!�HQ\����\y������!G<I¹r�Reܲ�r4B�(-J+�*�TEr�:n2��dRu0���Ar�N�B�.�".XYt(K�bQۊ�]��ҽz�߮� �V�V�}�}T[�����,�¹VZO�7σ۫�a�t�����.}��1hb�rܬ��V��k����zw���Ea=��L�S��4�5S���ߤ��Y��.��\f;"�ͽ�j�=~}vV{ݰ{=�`f��j_e�c}3��K���ء�i�'/M��nY�����[a�:wlZ�$���{���,эn�u�T��b*�z�R T_O2��HuD_;�ǡ5H_��u�����G$��<=��dK������2��в�D�����󞳐J���]W[�?tv]cI�n��®V�S��+�^{d`�J�d'Nn��jo�@�u�B�����W̌��.۩�(q���Ê����î�6rN�֝���� U�D����p`���!�z}DֲbG]�[���1��}G�8�aY��F��}vϠ��\��@�o�}���s��;��Yb����Q��oh�����yLo�=[�.�71y�a�ȓp��z��^���5�[��#��NQqu-��B��^zX�5�p��oU�����R''�^t�}$@���d�S����*��A�	�u/��v��ǫ0¸�SӬ�3�H=����ؕ���tkxﻎ��b���!)�ߠ�ػ��m ����)2���T8*vF_l�+�I��j���K�6j����M%-[��9�4_T�~	oK�mӻ���r3+�k�]�gjMw3���������r�Ki]wa���c�ܝ��A�����"��3�d���]��xdOՂn��=� W����~'[Q4F������a��`�P��̋��1:oeȴ�V�yS�\�㓒���k�yR�]��^Z�I�v�����~��4���`w�����7Jk�qV�,�ۮ���obU[��׬�uJ~�ܠ��K��gO��)��G)��!��O�}��;������ϲ�����p��i�.��ך���+K��+�Ux:�O��^��ّ�2Z,zT��~��#=cV-���kcw�L��q�c�u�cH�7�N�x	���}ny�>�����~���gZ�pb�nԥW��(ۇԆ��o�>
�7!��)��MG�M%@T_O2�&�^a�a%o�:6.���c�G7;���nݱ�}E���������TJW��E ���)��\��E�[�4��P���4T4��C�CN��؜n���R_�" $}�#�n���f9�֡;��<,Ec��a'���&¿�m�|\���7#
��?Y���$�ձ��ub��**A	{��X�����bʘ�׫�^߆�`�Sٲ���O�Y/�=�K�n�xǕ��9 JH�2"���p�̴Z�Zz�y8Q�ج��4`w�S�g��GE��>�4`w�ː�V67@����{Q�ܻu��]���0~:���?R�G���9Y���h<�t�f.O9�T� J�L�L��ys�熫Y;��SvI��������d��.��b�7}%TwU�B�'V�S�sq3��H^�9�/�\r���e˅S����k�����Xv��4+�~كX��g�W�B�����o<�س����$=�vx����Bf৖�*�������l<7�ʅq짥e�f3M��ww�}U
h�qQ�5��Cк�Y��Bt�3��ʛ7�O\:�;	Þ�)L	�+F;�W�<�ʍ�z7rg��ɗ�=�~��Mk {k���'�q/��I�'0���s�t���6�W�l����u������ǥ�Ì�9�(���ާ�t�t�>�\Wӯ=�P�њ��n	-^nl�������F�u��n���-,�g��zV���m �_SE��n:�~�q^}{c�U���~��Ķ��f	H�+���U����#q�c��ڐ����[�����_�~�gl]^u[��֩#��Ʃ���߄���F��ʧ�)�MG���p���}�[�;ߗ&�}<��'�ӛq�:�p�:s�R{���=Z�ͦ\Y�� A�,��HF��<g~�Y��9]:T/�4U�&�ớ�p��r��tu���b��U���!�IӃ�T�i�+;8��c�*3Cx�'Ʒ���ʤ�1�J�:@��� ��m����{����?T8�T���eo���._Z����Y��N��^l�]Fz�%l��vp���/�4׵
�j�㈆w}ei��y���VF���!eo^L��W��S��=�k��Ꝯ�X\_��C���.N�0�58W��HC��׼�8ʶK�ɛ�����R����t��6`�yUH��g��<ϰ�Փ�%U��o'����>S;��6��>�k��"U���S7��1-���긘������Wd�����Ry��7G����Ǹ\��{ɿh�f\xU�f���s~���&'�[YF�0�wP���!�q:O�k6�x���Qv_6i�Y�� ���^ u�y`�y܁Q=Lvẍ́2��e�b�k��<�_jU��.4�
�z{wY�k�M�@z\��
��\�ҋ�c��sٽ���S�q�9_Wy���=w,�m<�MDaA��fd,��T\���6�V�(�6�odm)5�LkIb��o����IL���Cn=������1O�f���o�ǢV?@}*r}���(��R�A˗~�]�j�k��Մ���j�>5��F�y�6�.���Yʶ�WJ�1���W7f���pd,v��}l��rޣ8��X�x�VY�Ϣ��fT]�j.���y�Bj̭�µ��d��u�`���ʰ>�J���n�����Ξ��Y�]�ʈn-�vw�?�_��d8i8|uT�9q9P�~���d�� c�@_z�6��!��S[�{�~]���8n�ی�CC�	��xkt�ԟ�ET/NL,�ζ��1f�3�;y���yF���CG��*�c;X���k��G��
�p�(��uX0���_{��BR�r����c&�uKӐ:J�N�k�L����i�[ޓǭe]�l z���1u�g7VOp�N���yq���.=.��FB����r�\s��zmU��{�Ye�{F_��	T�\��}ٌ���Rc��1S��+����3zؓ���j�=��X�q���g�����oQ4��w�D�,쀖�T�W�)*�y�^�C��`b��hf:�2xN�}��ׯ�!�kh��nߡ���x�@؄j�:�}h�-O�톢7�˰��YU���t���É\���9\
�΀Bb���9F�ߌ����ɿ���[.ʶ�_��ehK?y�έ��Z�e��4�۵
�V�d?N��׀��,���R����.h��.���DR��~�l8}�r�Z��]Y|4�8к��ѹ�f��W^����s\�R��kF�#R���.�rP:AH��LU��7;u�]������F�><(H��c�4�{y0�s��J��"ӽ�:��/��[gz��N�.��1̤���Mq���_��LL:��������6�����QrqרmP�;~�������]����;��������n�eǺ�Us�dTF9�w���9S������S��7F5g�M<7q=��E��/��2{��u+���^���ߣ��ɯ��3W���$��.��=]\ό��[�a_�	�q��cV������6�_�ӵ}9�c�ON��ϥ e
E��Dߦo���[��p���:�D_�iI�N�_5�\/\I��Tx���B��څ'��Z�����w��F�Bקh{��49mp~~�w��)�C�BQ�Ǚr.!���I��ɜ�NJ�X�K�39�~��p'gێ7vz����7����@u��9MTn��^늸{�t�rʑ�p����9�,-�qo۸b��z���2��XU�����S�����5�Y�9Ҹ��ŧU����x��4���ӄ�\�|mW�������o�/��Gh�h��MSGa	l��ay���@�sޡ�= �7������Z�ƽE�13�B��*}�W���@���n=2�?m/52�߻hѾ����N�sK��܅��P(��T5�*�y��
�l���x�;\k�6;������,�Vb��+�`fڞ�U�{4���g_N������R�����Z�Q)Џjr�Ou�t�*щ�;Kt鎰����]�@��E�r>޼Α�����g���;�M�k����Ю7�7A���e ��Q���辞eT�Q���٘�%�j��fO��X�),K����Q	۶+�TW�BSp�x� ����9.ϐ�����o9���^d���{�
�;�>��u=��ڹ�9+ц@H�]�"6Փ�wGS�l�:���D���{���}�%3Q}�p��:,n�7#
�!���ꍅ�.��}���H��`�yq]dLR�g�.{@B��ho�u]nc��s�nE���{*札���@O�ރQjk��OD�;蛨Yz�11K�(�/l������5&��;�M/}��ս�t���ٿ��:��f�>���ML/g�0¿:�5��׶�4|�¦�>�hΧ���,R�Qf�@>��j���Y@SBO[�c��f��~̨J�������w9���Ӷ�l�)E���3Q�	�/z��ܕܲ=�Hw�|+WQ��	�x��>�Nz�S�V���#_�����=9Y7��ɿ��'�o���@��zo�m����!����8?v~�|��׈����>L��\5�v�otA�]u��J]�!�$���뾍�֌�}�W���?1�������E�͙��O5���V]�W�~ؗ�{�f+��CE*�â�ǿ!����g F��ڗ���=�f<���N��mQmVP��gZ����C�:�u{��D����*��	�]ݟ�鷟�����k�,B��)�d�=�ڽ˷<�v��/}9 K����ے��[Ƿ�c����l�[~ea�Ϫ���Vy��kC�MȀU��^Z������wnpco��}�����)#�S�u�C�Q�B�,�V����n�(}�P)\�6������T(y�vJ�Ú�6w"��]�a�:3�1Y��D�	M�F�5��wRug���h����֬��fp$}��
ƪxq�g�|�lh�Wև���w���!M �\�-�|�T+3.��ں�����2�Y�R�d-8�c�ګ��v��9��N�����z���cN[Fj=�:�wg�m-�`O�ˠ5̑~�t����转���-qը��� g�n{�W��V�b�HpOT�Y0u����{_8:�hkK|`�����ݪŃ�,�Ѷ�:8�@��ū��~�~?�z_�ʈ���w.�Q�𖍘(,���bim<>%q̂��5 �:��7�%ޓ���WU���ܝ�
��=U�f�\OP�-�Hau?Oڱ��_rZב��[�&��x}�{m�-�Ĝ�f�#R�x�^bޚ$3�w@z���MŧE�]\������r�Q*�3us"<:�+�z��<Xͣ,=�A���T�����c)�v����DZ�}wu�*�t�S�a��I]�Ky�]
d~~��ly��7�}@7�S^ u�y`T7���/�;l̈́5���9Ǆ��ݝ�����By��ka�7^�3	s����@>%L�{z��j��U����)�7�n�y��WG���%��_~X�f���3�3�����Ժ�\ǚ�8j�Aϫuۡ��X��owtl�e������S��;?�Y����>=�5����~�O��)[w�b�ee�B@����f�F�`��R�fU�o�|c"5����>>�W�z��/�5��H�P8p���ͨ�F��g�/0��R��=/�F��$l<�X/���l�~�>U�^Ac���~�Gi#�
��yayֻ�Uv�0Xo*Bk:���*�v��mz�h�C���ew���QC=���oL-����p���qo��=��\F�ٔ2�S���=��n?\n��w����w������}(��������W��{p��<�<K�=������e2��+�_\fe`D���?yV\f�s�*t�G�$���Ҡ�"��LT�Qr��q�:XQ�i��W�3���f�꾖K���)�C�d���oy='��^3�nhZ�)�����h���.pW}�)U�B=�J��PRկN��֐�D^��S��,�����/f�!��e�u0U��{,V���Z;Ԛ�������c�T[�V4��W>�
G���������3�(��TY��}U#�2��/���w׎�1��@==������׼rw��������8܁���1�|���!)`/*�*y�x�	\_���#`�w�U�{0s�躘q�?���S�[��<�푂�ڹ�6n��CSpH�g���}Ʒ������Z\�s �G�&��}�g����� W���T���}A�/�Q9�27�������O���s�QJ{@H��I^5��;���|\�.IW sw@u8k��W�z�������>���C��3���ϼ�Qs�dTb�g}e��7
Լ��|���]�wMt�W\ұ�h�
��|���F�ǋU��y���ᨺ�,<~���B���L-*:�=���^��|�H�������"��p'�mԾ:va��z�+�SӬ�3ކ������d��@7��ds�,��Xz���!P<8���g���T/�څ(�bH0N^]Ov77J��9E��gg�޵`^�dy�!:q��#"�X/�yS�o�͑xW�Oأ{�YƇ��pǊ�ɯ6�)LQ^u�P+�>����R�Ѵn�nG͌�����Y�rΨ��훵�u�9b�U���b�-V�f��S���I�Q����ys;z:��wψwl�[���hf����AF�V����Z�n^�R�GQ�������u$��6�e2 ��q���`�����R����0ԜB^���ʝ]D�w}�㺼�ָwd�I7�uG����Iml�b�y�͗|akFW$6�n�Ӗ�b}r�έ�0�ĳ�<�؜�b�d��IО�{}�`�n\�+��<�ܙ�u^v�?�X��5N�ev]W�რ���7�]��ze
N>xΨ����k��y��W<��Ʋ�����(]�*�G�3n�P���K]\�0i���Yő��ǚօ��Yմ7���Y��/�
<���a�4�{w��rs�p1�h������7n�T�|�ep��ج�r_�\ޫ}h˼�KI�Yi���S2_����� �x��"�Vv�����]^d�*cg���ĸz����ɟBy�J���w%xOR�:���T�R���h2j�il���@�U�-d�srn��z>�}/6��Q4���n��'j9z�'۱�}%%���z�8��{��ROe\��ڮY��O0y�I�Ԥ�ZBn2j��M�ڀ�}V��Q��9g|�p،K95|�Q.�ʷ�e#���t�u�2�|��vc��|��mAN��������0k�� �o������r�`+���+l'��t�J��V붹�`m�m;�N,�����M\h�M����0�\&����=�=�PR*M���q��b�0dLtd�ks�4D�Bo9Q��@�T��u^ѹf{/�ʂ}ʍv�.5�ƹ�Y�
�N���.�u�wU�6*�,��-�dP�9�ۉ��ʹ��y�7��t��Һ鵸
k�x"O�ms��eV<��bZ�o���՝tNJj� �vbI�X�}�(��A`�.�;c�ш#ۘ��!���1�շ�dE��]���2oAO������^�6��/VɆ ��U+�j:! ��|����xg��VP�o439��rSu�ov]����x�GM���oKEм�v�S|Qn�5��Gf�i�n#%A�f�}�5�e��^��������^��2���xM�K��XT숴�k���	���x�n�߱�(lL[��n_N듏Kq���ג-v0�et[ ��K�#2�b3����ӎ��i�d���j�5�]ϭ���M������Y�p*}�)����Uh`-ԟ3ڦ;$�zY�mnr|z�[�3�]K��9�.fŷJ�φ�=R#O�G�I%��-�u��m�[�o�ɦ��N�AK�ؙ:�h�x��4[0�u޾�h��.��q� k��N�$L����%aA���-읕��m��׳������d��%J"��h]����t��d\��r��J��}ं��!Eա���2Yɖ�*�BIS$!!*��u�HU9�ۋ�H.�QW� ��*�(�+��Ft�N<Qr*����
��Jb	��U�(�E"L��.Er�ue��I!�˔]2��QUd$Q��Ƞ�s�˕!kF����:r��IđT\��*�AQ����Ir�es�AˁʢQE�
.Ur�)�H�
	*���ZU˖@DEDUAF�Erщ@P]�@R��
����9A"�Ae�&Ȣ�GVrW""
���!Ȫ���:��Ql�WH(���HV��h��d".\�r��3��F���"�ͱ+��M����e��i�jʬĖI��K0�ÑADy+%bDL���28Dh'O@}A�?b�4�˕��rښ�|�Wsit�����V�ʜ"!/dv�u`���#�Bv7�|9=]�U���-�3�wLI�z�g�fT�H?��O|k��;���o�.n*�ʱ�����rꍷ�}<nhxg���Ν�~�Ӛ�������:����q�s��=�C��S��Rgt����<��>���S���U�h����y8JG���^b�YC��;��z6du@�h�Zܙ%�p�c3�ܺ��<�����?+��Ϩ�y�]���EM�h�N���#q�9�m¦����22��ޡr��<Ƿ�ю%��Ct�ګ�z#��\o���Q(�5�1IP�/nve��ˬ��۷"��VL..�m�����ǎ��M۶=��z�+	M|�x�]��YKʳ/{��͚��#D����Vz#*�څJw�}����n�ȶ꜔�}�$�y}{X��������"�@��^�a��S5�P�!Ww�9��O��"�j�Ӵ������~��"���*9�H�:]W4�Y����C���Ϋ��mf�y�ʽ3�z�B�z_�e�*|[d��5�LF�B��"���_L���{s�o��Ȫ�=k��Cx��S_�̘T?�%�;�dCUj�a�d�;pw�ޱjη����'#�Y�;�v&+~R�0u�f��	+�vc��t�DyRU[�B�D�,*]e=9�����!Hn"#f8vrd�[�yW�b.3���Y�6�Xnͬ����*��e.�d�T�b#��QU�"�*�w��I�a�VU��h�ꚸ���� ��{wi��k:��d�a�Ϥ���)�f�US㾉����lW�R���l�����4��.G�vq��,�U���ʄ�z��7���ST<�^�龇T�o��xN�͹��>�Mb���;��2�ʆ�Wt��d'���N�C���:��7������n��/{�c#�\�C��
���d�aA���%@���p����.��7�.&;�c�n�����?vF�4w��/�Bxe�S�=��b��ؤc�w����S�:�����Ԩ�u���\y�n*��{� _~�>[����X���Y��??`��8��ĭ����.����W����v��s����z�e�1k0RG����y*�g/��ZY�+�|8K�s�3�Ƥ��jC>V���h�C�1�
��e��ތTiM��S念�bo~�O{4zS��G�q����9���q'U�Ñ�K��F:C��u1q>���t%�l1�(NL�v�����!xّ`:θr�J��4׵
ƪ�>��{O���n�팱���%���dȟXu٬U���6f���a�9޳��K�Tgb3��*R���=P^���a�=Mu:�EG4Ʊ�z��CU�'u�s�@x����f�=��!�]�_S�c����N^��Hjl^�VFâ�e�/rT��>��Pe���7Pp��.�1FgE7.K�' s���}Le��9T�UH�J�\���(wD^m�I�Fd���9�6��&��5�u�~�$��{p�K��}�H��
.*�u}3���G����c�/kB��%@��ɷ��V�w������=�1_�~�Q��bG�0x,��c�Ki��Į9���ӧ�>5^�ѪO�^�a|����-�XN����6���BS� -5�ǳ�����j1��ۄy�{���9�w�	��܌���[>��@>Fl��X�n���c�}�+(,��WO�ȥ�h ����$�x]�+Gu��x��||۠�S(8O� [�����Q/,V��u��}')����nxe�+���3Q(a��޻�X��\���:\������LW��}Ր��B�YF���#�X}���:v��ޜ��1O�g%ߡ�C+&p�r��w�J{{���Wճ�O*���>1P����勞kב�o�=g��X~k���A���K�� <Uh�m=��V�{t�{����V���9�W���{.�~\�[�N����0e`��e�JDS�,n���m�ی�j��������ZҘ���n�Pqv-T��'����܍�d:�Oܗ^���=#/�����g���m+P=�M_J��3u�,E����͕�t�LM����3�g��G�o׳T8g�U=j�ʬ��_�_��F|��l:�zFj���9G�q:��^���{��t1Ǻ�3�㝏��ٔ3S����;��3��z=��3ȸ�bL����<�;�O��_�����S]¿L�L�s��4��V��2�Z}��� b�1\�ӻ��q���ǯ��dZ'���V�5;�T\�(_�x<�ap�\pwo��ޕ>5�5�Ƽ��s��V{aq����f�(�e� ,ک��R U��*���*��d�x�V��閇��������l�n����B�2��'�,�#��y�x�s>�������:�x2i<�J��K�wG��p+�l��\��N��/}�CR �7˽;��O)�;W���޴��\�f��j��������ߴ ��b�ʒ+�����k�.:��x�b·`�z��&�wx�a�l��}��;��L�S�\�Oz���L����.��^l�8XŪd��v�|s�t�y�n{��S��=�B�dr�70'T�P)���w�QYet��q����n-�ۏ�n�����-��f<a�/a�:�^S�����6p�`��t�`>���#mtԃ��"Os��r��KĨz�w�r�K�&��X�茨�+ �������������^,��e�Ĩ�1T��|��nv W�Ys�Z��P����I�P��PY�i�L[��֮zM�_��|�ӓ�}�Ծ:ja{=Y�_�����3�����}UZ������&��.3�<� ��:t:��jF)�sX_�� ��p'�n!Ծ;蝨{q��0��e=3VTy��5�K\�UAt���<�.��E��'m��"��
�q�$�����.r�x�k7�Q1 ��v�/{l(��q�#����vn#i &=���=<�n��7�w����\sʝ;\���\b]��ק��#8�|.���/�oޗ+qX�X��7q�m�u�{�����ע}[:�ѝO�H~{*B��e`=�2��XU�g��)���yF����m3�_�]mGl�m��Cʋ�+'F<�]�\����J��)����{�Ux	��P�L�7�|V�;+"�U�θ��ǎ=w�Eޟ]=��=7
��3�Cye��be�T�>��S�@�sȊj�c�������+���Ac���E�:����盤7�ݡ4o����s;����z!�z��̪2��6cs5nC�=��0�W^��|m��؁ʻ�(/NtF:Cv�t��+�d%9���)���!���T�X�{�1c���RҨ쐓���������;�V�La�j0_��Pi�l�wWS�ܭ��K�j���q\n��$��_J��kdToW^�6�.���VT�&µkY� ���uz�O���Rw(����>Ǳ�����-GWǜ������-n8}`����z#*ݘ[��#�g�u��i�?P~Ev0|m7;�ѻ�4�������	�eL���z_���)��ڄ�i��\��4\���s]��m~���'���d�^�*�S��1-��ˊ�&iN��3�>�P�F��8�A�S��Oo5�e��s9���>�3M�̐.6
Gn&��ަLLE.��q���'��ҧ��g��f�8��>�������Mճ��Ҥ�`?\k昮.��:Ee��ovC��ч#�4��w�ǝ�)pۚ�2_�}�U�o����}���m:�����r��T�=n���')���#sw��M {á��_fTm�)�+I��L�^���]U,�����Ng��#�6{j(�L"��'�l��U��:/>��ӕ���0����y�d�z�Q��R�
��{
��.2|�_ڲ����}>�q9Hz������Xn1H�7����[&�G�-@��I[F��&+������\kO�Ȃ�~cd��A����Y�z����1F�˳���:�\�������vj�V͍�q�ѱ4���S���	�i���A��ح]\TTD
Ij5�N�F�s:���\�n��t�]{��SՑf��Ag���
ч�� ���T�ќ��-om�z�ƶ�c�mZ�s�bg�"��k�D���t����}�N���d�@~��hO�S���:6��|5���Y��.O�OmT<5���	t*lm�%������T���|N�mHCn;x|�SGr!���5\<1�ý�U#*����?���ޫ�,�� qo.3��w�,s:�aw�U<>�<����4\+�B���(�'bt7�/ay��nU��}��o��;&E�⓸r�J�d�\om���S�|�g0��zp�e�U����=���7��d��O�U�6����G�U *.P|_��C�g�N�0��46A�y�f���y�/�5n������0�nP�*��B�T��d˥��6����9�#SN���=�A�6^7T��*^��^�"��#q�Ah�A���kw���M��_�o���d��	Qz�>��K4k�|1�ç&����=\y砋R�@=��L��􈓋/¼yr��G�K����Z�bxH��+�wO�Lw�*�|�����N�|�n�	����)���1�#�?t�?s�6��Qj�Max]Ұ���j�SE���*���:%PB=v�9�1�o�b��t\ahT�������ʺn���F>-��R�<vb������Ғ��ĺ��jS'3�\l괁4ũ�:���{��ǝ�1TW����X�3���RWO�F(�2�_<t�ZVI8�����뿢~��_�J�x=*�~)��¦��(:��{н�]˘�=�h��9����|�n�Y3�NQ�Q��Ea�'�9�;_�ߧ0���8��gc)���q�Um:���h�vH�q��γ��>�;7�<�m�1z�N�rOL+��=(_�k�ED��L�5��7Gj�Xo��*<��@���`_�ϭ���=�ޏ,�8>��)v�6�ˢ&6�_z[ӗ�^k�ܞ����Hcٸ��<�ߓ�qz�h�>�\-fQGR��]�own��t�oh>n\E^wp�N)߼\F�e�]?�)��Q�k�O�q��G�P��sw�ٔ;vހ�s����lUh��W��yL_���}�h+��x}	�eq1�v�pٚܣ��r�ßnu�}5�me�{��F�R���?T�W/���x;��aE�^�Q�-���Uϰ�8��
��r��ҝC�)Q�r�)�����&n����"�ΞeW�k6Uy��ڴ{+0�<�:�!p�V��=�IPݿC���j��)D�bDpʪ�u��e~+!�����I��T�:�+��o6�Ƶ��o]޶���h���Nٝ��ȣ;�
H,>�z�����Ozq���K�-�:�tUu �)4�Aj�>��������*���c���5�2��uΔ��^���!mw�$�[�xp�O��Ynv5�F�p���k�c��׺��J)�q�y\
O����Y�W2��~.sˉ5/{z�=/������W���g �=�	���P�V�g��h<�x ��<�=�99�cK|s.�O�J�R�$,��@����"b�����>���Q��n�U3l�\�����Σg�v�IU~~�*7��RE��CsΈu=�Eb�g|
ޡP���ُ���������#ʧ&ض��rn��CWNOQ�/�l}7P��=Y�\zX�5�)�f�A={:s�؝�2�VO�}e�<ԃ�\�p�D��Ox�,{;j�s���ͪ1,1���]���'��t��v��k���oiIۆ�?ް�J�Ԏ����s��<�v	^^�>�q�-�wʬ7[;7��޵`o9�GC��+O���"���DD��f�M�q>9�u��տ��RU,�k���+=�5��#�@�gP}6���Tn�c�w�8]{��J�{G�qO�nY�'�#t�V�ߛ��V�KK?*��;�iC�J���ž�R��@F�iV�B���^���R�x�l��ɁF�Q�A�u��A������k_o8�v��L;��e�u=����Ҟ��ሖ�9~Z�LT���O�mAA�ɼN������ɝV�	��X6��]%_faA����i���U�(�S5�ܟf���ֺ���0WzwM�~^�~�q�Y8JEO����x	��P�L�7��nעF�:��S@׶�]98����JZ8�V����ye��F1T��h�ت��N���x<^�-D����Vzf��'s�ix�5:��q/���6�]�C��Q��qN���PS+��S��U��y*2�32���'�U�\j����T��FO��܇@x'N�͟Q���03fz��������7���{��t���l�"��T�|���ѕ�E��"�w��q�^��޸Z�{{C�����q�ٚ��r��%^�:�I"ʗ��C��ђ��ݨW����D�N_&2%Mp��]U��N��~;�?]1N�I�X�����e�U��)�px��9�J��~�M����ϐ�x/�v��/+�Ͼ�>��߮E��$��\w�7P���Ɋ]9D�wϖ��m׵�(�\yЬl֌{5%�̲��v'g���?\K��S�Ʀ��)����~���k�g�ot��OIxVW��
ޱHj�,�j�}�5C��
���'��>���K3�
��?N�Ss��M�Ց����ǫE[�:����+!�ŗ�O
m�eqC�˴��E�y�Y�LJ5s4�3���N�v@�8��h6�_(�~��λЧX��EB`�u�Ne5ΰ��%Z���wA�n��#��Y��d�����yH�3sq�:UҖ8�yd)dWy�KFα��d�nZ�%�uB޾Y����]ʣ Z.�SP�����?�����_u�`3)wS�-K�S���k�^g5��SA�zc0c�t0�5v���Z7��&�v"�kZSS-�*9��b��O���Qʚ��*�=��s��;WB�x����2��QF�q��UiX�������>�4��{�W���=���}F�e\Yxz����ZmV���9n�D��ᆭJ%I�i��G rn��U���Y�fvDp��V����]�y
�bO�7*�vӫx��=�N)��.川�f�:�C�EhWgiv�D,��X�$�D�rU�L�2 @���Ho{���p�X��\���VM��.����w΢�����!)��}/n��]3%Y�K-�w�%�Z`gH�4{H�N
S%��b��3�cyq-�=l�J�u.�Y&b7�ќ2oʲ�M��Nߐ+U��Uj�J�\�Yk�����Z��XǴ�A��8��X��"�U�+u�E���RX�fh	
zk�.���/�KThNޛ��QpPJ��]	���Po����;c�V�Mz��n�룘�Y�F�������1֑D-q�b�V\6�h
S��q�x���e���سM��,��Xr��A�:�������:=h	��A��;�&�;�*2U�ζvݎ���Yf%�Ot��(Qt��5Vu���Hk������z�����鉁Wj��Lع.�W,��-��0����*:�q�L�+8����otq��՛BV�P��֗cD{9� Q�x�]�E΃V��������Q82���]J�Nر����R�Cm=���W�ުy�En�Q�����\���ԥ��<P�Ր���u�j=�䨾�{�@S����O�uq�1RpLY�Fib�kTǖ�P:��XȈ�7z���-�K��CB�+/j��t��B�u!�s:J�63Wݝ���B�t�h���*ƶ�r�+8<-�i�f¥�tup��8�7�9������v^Cy�kH�B��G�V������͘`��G[��� �Vۍk�*Ó!�%� �����S%��R�s��}ۺ��w��NWjcvu�n���{���^�\����ma�]��3cSO�%�j����QA���|����99���qlM��ƍ�	��<3
ۨmA|0n��l)��w���퇱v��W>ş z����t���a;�	]�o�U���\�x5|6(�	��[�{��v;=*��8n�����Urӆ��&`�EG\��b�Oz;�{�b.�I�NP�=��:�s�*��{Ҥ�u�)������Uwo2��E��uϸH���U�STݾ��K� �����"(9E�i�ITL��Ad�"e���q8����4ΧB���Y��
�(�TAfr�t��q"��˕�i2����AA]P�����E��C�
�&m6U�8Q�	'*I.Er"�*�)2#8��(�jTAr ((�����Y&Eȼ�;q*QEșEE�L�
*�Z�I"!0�eBEU�\"-����UDR`�8$�0��TUʪ�3�ҹL:m�Ȃ숹(�29�D�EVIG#ē*(��2�L%H� ���(��G)#Np��Up����h��I*G
�H�UQSQ".f\�X�UuH�U"��*���V���� ���)P�*2 �R0"�"���>�=�<���o��D�g���u}�K�Z���������غ�H���4�U�mv��B���LQ��{(;�yu�K���ns����7�oٕ
��Wi�+I�ʄ�Y�[�K!��[�k���e�kV���j{������ma�7�E��>����C��Tnvv0��f�J{����d�L��OR��ih/��M9��f\M�yg�9g�x{')_����㑊F9�Ҁ�E[��wk_��o'�.��<�I�]Q�^\�X'p�:����C��(x�f�8ǀGy�w�7VL�(��#�ep~��S���ߛ���C��xJE���٘~7��d#R�V`�8^:�=��7��X��ڐ��˝�/T�8�ˑ��~�%��u�_o�ņ�4�bW�g3��;&�2��a�K��b�\;��|J�j�B���}�y���lh��U���tER��'�y{"T�
�<�"��M Ϣ���J�T\�R�4���z���b��it7�*O��c#L��]��N{nC�~�E@#�z��誑���P����x-z��=n�v������O�Îqը�#�bݫ���衆
G�.�GTL�=�⧙��9	����@4����q�%�K��TC�nv�ܾz/$h�D�]+�n����x����T�)u��	�n�����pX���8��y�y���p3F"���HM���������A�h^�`��9J�I*B6�eV�-���I��4�v��Zy8:r�;-4,�W;re(�G�0oB"ݪa[��e�{<T�<���������l3�4/eW����潖�v����X\A;�3�%��t��&�Ee0y:����A���s�N�+ɞ��z�:�t0;���11K�(�H�l|&�w3L_��[>�j�h v�j�/R�����{T���Ϊ�N�A����e��d��
���^9�f�Z�sf�@><�5�!0�������:�� �K��b��>���2��X�)���0��Fo{ޅ	���WD�z�c�kF���ő3��wz���HEa����v����~���O�g.g=�EL���<�O�k�ڸAU��;7�J~�����u'�_�9P�~��E�.&=�m��a�L�r��1�mpޫD�{lGϫF���lH�{��\s�[��6}�{��s.��}�x��7;0����7�WRˍ�Vj�gi�_>��C�>�\+�b �O9����I��{����;���F��Ү�ɟ9��j8O/�;x|�S=�����G+�2y���~����Q7��ZG�Ն�|�l��yT�h�����#H�����xCvg`�T	�g_�wM1X�iZɪ����z\E����9-�|��B�K�C>M[��l=y��^B�]�on��b�ҩՎ5����v��o�����X��\D�+��_ﷱ�=�P�����z۰�ҽ>��ʤze�FB�êޜ����/uz�:�.�p՗�q���^����:"���R����MN�r���x;�b���^���t�9�2^��:�)���y�?q�c}���r�����H��s L��"�;N=�g���S�AW׊�1��!y.+t�'@e?[�1P��%#d�,n�,�ش�Non5w�˗c��Vx��Wѕ��t�r�wCy\
�=�0[�R2�n�n|��O;�6�j��[zu��d��M��
�������3�a3��P��U�����z�w�s�^�~~f!��i�~��C J��F�������"��>�3�}��f�}v���Z&�Nx�fil���p�W���9%�J�����R��z�\w�7He�y��{�Ŕ��=(���1��K�Wk��XqN3U��ǡ�@젠=�'��˒��Ծ=��\{/��,l�w��s9��{�wz�@r���59�P�]E�6�NO3#��YV��7�|wӵ|�J����.oI���fV���V��o+��2��R���:����ӈ\X*̠��T��c�^�;}��z�j�|�Ek��5v	:�:'T+{���.�
�8��W*�Y���u��v���m`��X�b���F�H_1�L��Ir��ƺ8S?���o��%��OPc�ݱ��Rȷ�j�y:�E}���(��~Ti��|Iu;�Y��j���t�V�ǜK�~7ݨ^ɟ�)����@	���y�2;�Ԅ�y�#��}�b��֨P8.o�VM�7��=�{tZ`���r�J�Uk�E>��3���7��V�S���z��~�s8�(ګˋm��D,�����{�U!�3�dzg���o�2E��W�n�eU	�i�ꅚpx�O�q�K�����7�7�q���Y�,XO�n���<��-�|%��<�����H�=��C/�27��\|�ِ��\�Դs���6T�Tz���3��R=&����2)OrmϽ��+��v����7ҸߦX������b1ľ;�鍸Uw�t�+��t���5�.;cubn��5�SݼC�3\�zgH��<��FT.5o*��]�ќ��]�X0Sv����(Z�������f�8�27������������/=P�����N�����QI_I�n]s58͜�|{l9/�nG9�Ev#f#�H�/�C���d�j"�j�v�v��b����o�MDﳻ�@�W( ��9i�M�YA����ZU�NgT�y�<�Ȯ���vet�y�me�ȳ���N�YW���_fmc�V
��.8���ff��}H��M͠rsTwR�ݝI�n�����ՠ*����Q��q[�#oIg�c����~܃�gP�UJH�KD@ཟUq3�Y��.{p�xї�-�V��՞��JO�1ߋ�<���Ә���M��%π�oރ�Z�H=��n�eǩ��|:��}���
����6kq��ј�OwMIcul��=�U>��)�f�}UO��U����C���wdWG�9BY9�}9%���um1������2Y�j@n�MP�#� LPqblF����7���v��ۅT��D��oٕ��OMƕ��FT&j����2�約�^�[�[����y��A�Beж�TٸN$��#�r'%[�W�7�aA���@L{����v��W9�W������-���3�Q��Y�q�A;��	�9Hz�5��=,VDy˘qbH�ٳϼ�������K�*����p��qO}GLo<5�}�:���=�8P��њ,ũ��,Y�9�٭{E�H�6�vnR lFvu�-\��o����W*E�T[rG�[�)P���%��_G)�q8\G����3q�9{jB���h�C�1��=�x+�O@�G������	?Z��+�*�8H����V���6:V>N.���Q�7��}��#�N��(�䓭Q�����V�F��Q����ԉ�v�Mk�7;i�u�sb�T[w/E+�� P{�N(�	&b��:Sms��4��r��;�f�9c7;�1��eO�Rf,V��~3�ߦP�}�.&�U�>�y���y��d$b��'��ػ�TL��k� JFx�E�)T�^�2h.:�atU�z*�^#�VH4��_�/+%ܱ���핦�u�l{�QEz0�	�*�[誑�T���P|_�P���t��)nV��j�U��W섮��'��dt��Q�G�7n���Ҥ�~������UH�y�����ۦ��}�}��*h��������!Uk<=�qS�F+�����R�GlC1-��,o�u�3������;�q���>%���@,>;���Vգ핶�XxCWLE7d�p�Z]8�����;�g3XɞL��7�ǫ���������f�o���-P�� u��
���㳹0|�'3M(�ҹ�z����e�-�I�+�q핧�Y��sd�_O��������-C)��/�J���V˕5quLwM�~���q��^�Q����#j��5e3�)�/��ةr�]���*���ꊝ7�uX��6~!!�۟߄Y7��O]�?,w�A(��l�h6Қ�ͫ9dx*D{��Ʉ���RҺ��{�t��L��S�{���ϡ����}]so�ʮb�Y�]�ݫՁ�OT����p��c��[S���h��AG+�ß`��'����=��m�ב��2�2��}�cT������9�1k�
�>�O����B��z��Ii�o�av�����8;��ru��~�U����`y�h����������g�᪺��a�oL���<kՕ~��7�9�Hc/qX݊����\6�+�N]ľ�����_�V���[�H^�(���uX0���^�W��q������2�_ڝ�/Jgs���acc,V��w��8�W��o��Ւ$��W��U�&��+��)�����}��aF�a�{�\��^��w�f����)�>~t4�T��d�Do�1n]:�{���\�9O�.��pam�8=���]Z9���_�:�>���Sn����F7J����R=r���#e��i���7Ҹ��SQn�1qͫCѮ'���ݿC����/}d%:��qo[�k���wnmP+\UH�ͥ���ʅ�}}�*t��5<
yDxe��5����ué��~�v��vON����pH�n�h���Į9�	��څp�m�����r�c�N�Z�G\xb�2}KK����6�Y�)_Zi?[�]c�_Ld�,��UX"EX#y`|2�1��%r�v�<���W��m1K�VU�h�]�sr�4�#������e�p�dS�nw	mP���Ki�؄���_eӎ�evI�%vˈ������ ��D8��S�-��f��D�R�Þ3�|J��sp�x}7�{<sv1	~��mj�ǚ[��5&���߬
�WNH*@\sf���}s�dTb�g}���O�%g<��q�H}e��Q��9���mP}*M�{�^�5L������mG^�V���,��<WtG_�����4�L��t���4J����5C�}	��]d:�Ox�/�:�=�d=�6���#�~�&$)��O}�3Ҁ��.��E��'o�ꄊ�k¸3Mbn}���=�s�3�Ϻa�6�j�8rcl�ɇ~���)��٤ ���V�2-��+��4jӹ�D�*v�x':q�={���$�ˇTG��NJ��G[���P����en+ެg!�yT*��{���⽭Mw��+��t�������t�,��β��U!��*���9��1H�"|�9vOF���cFٓ|7�AF�L>���}�z����R9>���V�1:��:�i_�v������zk_Ql�2��#�d�X�&�����=*k�<ߨ���EI�T�����z�i�H���N�U�6�D���Y��O�����"H����[^�W�:��؁u��������{���i!��5xy�[a��Y�z8��� ���]�Y6��a͹�#���p�Zhh0�:�vۮ���u��j�uwA��Ok�G���G�������}K?0E�n=2�?F��B��w�5ľ:�]1�=\����yo����~x��E[��{o/�KӾ��:��_�2����
N@�<ʥ����Z9Wq�آX��;�D��3�:�f�Rh!��ǝ�j�2����� �}FG��J����/=��}{�
�;�/��E��,��}��q4����v�G�s.J�#p`�r�D�/K����}��L��С�slGy{r&���qJ��9���rp��?Y���$��%�f��Dҝg�an��W9��T���Wg�4Z���9��1��g���u��A��HiΛ�[M�髣��/{gt��0�z����Ӿ�=]�rP��[>����S���)�f��_i��W����듴�ƅzR����?l�֭�8����x��D�
j�gѠ-ͬ~7�=�²���_Nn��,ĝ>�T�o�3a�fT+�S�q�i3�	��/z�]3,��=]\y�ߘ��1ؚ-�VǦh�t�:�;����ς��V���3�n4�6>���zy�%�_?��Ֆ�����*ҦºJdjס��� ���"z�=BW�b�\��!�J��6�r ��t�X�d�#�VOh��s��+{�il�:�]A��J@y�B��X����,`,y;���CJ�*�\�q�G��t_;����=˞]��Ԃ����q��WZ}��TM7�p�9��Bxa�B�g÷��a��1H�� x_��f�oK���c.pp�m�q�X�A�n����u�[ܳ�9����R|s�T������7�fҚ�o��8�{��锍��@�q�!��Z W{��n�kw�p�yY�-f
Hף�mD�֧����`]g,�l}�a73�~wL_ޙ�|K�jB�����R��?Sq�w�m f�.se�Yy�Ӥ=�Q�6�|�1`z"��+���C��j�B���x}�y����	�������FU����G7��
W�@-�Q��@��JY4�m���@�.�>[7�[��^����9����V��FϨ�x	r��$_�R��ŷ��p�fVz\��z�L/?�hW۴�{�qը��5n�¯|]9(a��0/tUH�6�������eGe�5u�U���/㓬�ђ�U�hWJ��2�E�����WpD�:F�}�1,8�+w'B����c�������&&�+��2����q�5���u��~�pL#1���1�m��1�m����cm1�m��1���0c�Ƀ����1�m����cm��co�0c�c1���1��`�1��m�1���`�l��co���cm�L�6����cm�1�m����cm���cm��(+$�k1�� :k�
B ���������<�R��֪�*�*�)�P%%fjD�*��"�J��B����Q@6����*D��E)T�UP�Q*�4��z�6��[f�e��Ѷ����n �\B�
��E +�� t Oy5H�+�"� p;eUD����*�KI5Q���d������ͤ��PK���[*-q�$�s�QF�]!�-���ZԪ��v�[�ԃ�(Wa��ƪY�Nƻe�q�۸�L��M*���, �ٮ΅�����4*]2	(!i��I
�s���miV�AU1%l���dR��:Vf��4�0�����6BM�4� .�%I[5��Ͳ16ɱ���b�U
�:�f�D���А�T-
[c�"� 	  ���T�* & L���R�5`	���4�����	�@�hѢO@�=L&�jB)� �JH� FL`��L��0# #	��14�JzH�54=C�&��4 �LL#\�r9r�n�+�,e������5PN���Q@Ux��"U�|�����@��c�~�?W��Xr�:���\AT��� �"i *�$F�P�0�M/r�>}g>���~J
��Q^�+z4�DJ�q��H�U[��P�/�3=����_�kr�m�- �әy�Ii� �IOj]HM�GXۻ���B��4��`��L0u�H�Y�l:�Z���u{5ڰ�[E̹1�)P[v�)���ΑF��Ղ��w���Ƿ�ES�0��SlJtW�Δklv�!�ѕ��o3Ve�5JBK�m�CM�k���n�Ӽ;&�u�t7��Y�3R[N++؎�si�GR���;L�
��v�5y��
������̕�M�eռ�-�-LW���jZ
��X�g�S�
N@1wN왺�38�R@���I�(�^�m�v��"t���o,9��ʢ2Cp�C)ǆԔˋO�,��[j�H)^��̒�X��mȊ�t���a��JR���sO�M�����qv��0�V��ʡp�M^r�IdQi�T&�iU��H��*JĪn�{P�6�3��脣�dDeZm&�Ф�*m�S�������	t���r�[���x�4w k��Y�Uah&���,$Jퟰ-*��QWfmؓm bh6s&32�Yқ�$e�F��ݺX��+2��7�ul���e�D+a
�G���f��]�r�5sdah�s/F�mQ�V�ڻ'$+ �&�NM:�&dpU��ͨ��r+	�Y�h7�^Ĵ�&#wo�u�n�u��Q����h�%"�tSj�G���%�[H�ԫ+6�{��ِ�3C�rk�vڎ�4�h�˵�L���m�.B����m��KU�Y*��t�E�f�L�C2�.�� Zf�WE� �)J�f�L�P�dw�f� ;Ah��DK{WWd
m����#���*�Ҹв-�ud��3U�O�� *閳]�&���6I��e�F��(e�h����dhoj��b���'b��p�S�DQ�7Wa����]�L����=�1��I*y��0RW�Rb�K)a׀S��su2,'��Y
�55��Liw��M�8TR֪�q
2��Ӻֺ
���ŵ��k�7X����Lt[��;f�wr>�d�������]�)DPA�\�e+)QUy�S�f P�r�n����d޹�z-����P���i�4�[������ح'�l�q�;L
�(��"sJ��@� �,����X�´�o^�QM(�8�T��K�.�zA۶1�e��\#w C��K��"����f�4A�)80X�y�ۀRZ�Xb���6�l��n�^
�S��L�iRb�R�(�ȯ&�K#c�M&�2��j��c8�X5��T8%��6��mP9#������V�͝>�I���t���-);#
ǿ,[�LdxK7�<z��X�r���6�4�=ʰjF�,�d�ܣ!n�R|h���<{�̄b?�7Hi���I�):��$.�'@�bH(<z��ѺΙ{�g#�Y���KJ7��tr�#F�,�WP'�B��|j����F��ai܌��DQ$�o)|q����2��<V�AǪ"��{�Dǆ�����8r�P1�P�!�vCW��/s#���꼅�ZpUn��r��E�KT�B�x�CV�8�}w,+�̷{-6Jx�5'��M����a��F��Y��`�����r�LZh�T�����"U)QdZ�n�,ͭW2�i�?���|�]N�is>nZ�r�	h��&4�W°Tb�ջܛj��(li�)�`����%ѓIT��`TE�V�f�kF��JxH��oQ�	��
����՚�M�E�^��e5����KV5a�4-T�����3h�ʗV0��Bk(����95��e'�e��x%C#w���!	 ���L;V2�.�̆D����R�c�i��-U��@4��������h���JX���t�5��`��+r�:�j�l	�Y;n��I]�Ϣy�j�`�@�R��Ѳwt�q����N�kcF�h��D�e���.�Uf���3��
��V),҆ԇ�L��.�#)��PX��H�b�]��1y����-�T�+���7+U�Kj�Be<�3!��w,���R�X�E��nR����:�x�B��+-b7a�T�R�������Y�
����{����4hެQR�U=�"ѥ��6+ڠ6��T��w��c^M�IkX��ücVEz�MۢI�A��&���j�tV&���Z�[�g0�aE��7 4�f��J �b![Gn�[M���!��p(��(2��&�t�o��e4eK�ivf�e2a��l\��ah<ƅ��1/B9Ե��25����3	J�I}�4�ה/&\�������V8���U�vP�R�T�̘�X�y��Zh�5���l�/��e�kY� >�4f-b�Y�;���[�j�S�J\Z[{�)��Lp�s�y���1�_7Ͼ5����:���S�� $<�ڡN$??�?!�R~���%�}�sH���\w�A[�Z][���(�@L׶�i(�n������;�;93E�f��+/��X��t�]��]�����Q\H���f>Z8�/d��ő��,t��P��'p�}��Ҳ��0��]M��w�=P�Z3E�G������qw[��G�h���nwǂ�9Ȼ�*
��.�<s,puoM�Ў-��x�6��$��W�ac���q�g��]
��ܮ�Ρoi�6�x�����p����5�u������gY,~�ӥRH
�΍\՚�B>=@ˡ��m����Q�I,�W4a�Z��#֞t�E��zڷ+%��<x/u�F]�k�ņ�e"��.=����Ђ�&{�	KJ�R����ܩ؎=]9����&�X;l���ZRt�N�K�l��a�S3��-u7�0)B6��7{�u�r�cᦓ���l�pjnf��V�1�ĭs�����6�i])W�V�ܨ�al{/�@没G&L��5d���Y� G�N�4VF=z��i1#:6�d����Xn��v�-l5��V�GB��MF��˃b��K���}��*틴(^-�3����\����	{����R�Π�@�]]m,�b<rk-��q�i�.l�ɷ���!�vS��ju)���^�N�!� �ڄ$�V���:�(\�UC1�WHTt�<XH�|D���ԺK�}}�fv���@���í����j�M���'�2��-o>����;Ɯ#l��ˈ���`�6�����G�yZR�oH ��	��k��8T�gh���F��=]{ok�걂s���^y���e�Lٖ�i�]�+��XA�8.���U��l�i����}N�g^-uw�;��vҴ�N��uw{I���nPm��(�lv��n���דy+Nz�V��_X�.��Y]���^	��bzT�x�مVj��[��k��A]W���ܛv_b|6�*��G�Oz�)R�7C7����y�#a��V���Յos��ӏ7m����d�;{�/�� 
6��]@v�Wm�w'MR�*9t~�b���h���׽K�@$�I��~����ݮ�z�bQ��<�u�0@x�,�tĬ���ʂެg�Ʒ0�:q�R���[��[�쳣�T�q�jz�)kK�@��i��緣A��;��;f짣��r��t�H;O.�O]n�}_�4*�9�uМ�a����˘fg_w)F�06�1�M��,袐hm>�ׁ�p��c�٣�7��l1,X�W���_M�"��ܴp�F���]���*5�XC<�ƈ>C�;ݘ��u�����P�>/r'݆��V��_p��#��X^�w&��;��Tn�k�����I��ɓ6�nLqgQ�����ۨ��H��g��=�������q�z��Y�`�W��C1��:j�m���˷x+<�L�ٵ�(\�{R
EdS�\�h�T�v�Ζ�V
߷TR�w,��u��&xR�]^m������TE.���;E�� 8*fj�(�����5W�d�(J=6Om��LWZ��V7�Wrx��%���	D�}��"�o_g�ƙ��f8(��­[�z���_`���˓s��.:�ɕx����<ѭe�wG�T{;���+t)DR"�K����뫡�%�G������iƧn5NJ�c �̼כYY4R3%Ho,����M����- ��mm�&�ɗք1��Tc��T�@��]G�D�M���L��Y�ۦW\����qv��."�7ϻ{;^u��2���+ȓJXp (a������� ����P��[���h��of�:ԫL�:CZ~V�S��e�:����a���_Y��}��}����ζI�&Շ[ �[���`���j��� ��4ڃ�M�r׍3on����+zi�6�Y6��\���j���(+e,�ܶ�̓���*QVU�ܩ9�P�w ��?c�,�mwP���|�fI�/�qU�&8 �qm��pǮ��jYz�T��On�䕺��ڷe9h�o_���{�#-r������7w��U�Iy�dK��I���y[ ����ךo� �P��JF� +������9�FE���7ƌ��|��ت�嵓��ާѭ�J�+�S�\B�&�wl����u���(;jeF6іk��n�S;��u	ejR�/���*Ꮺ���|�S'����4�]�~DV��A6v�Փ	k�͜��#�Hq��p}a�R�h[rC+4�Tn$��`uIMqȞ�v����fg���ښe��y��s�*�X�}m�m�C_!C���L]�'%B�����SS�E�4�a�j�֒��s�̡�	�d�E>&s����x2������3~g�ӏ$��c��1���*KጧNێyf�����k�*��4�V�TD�
�E9����s�"�'Q�#��V��kkƛ�mץ	j���xg�7�B�V�R����;y��Ol�]3z��%4]%�}��1��+�Ըe�����k�����sfp�9�k��)'֦-���ڹ�лfRoۤ��-�S0wkK�����ȜZ�]��ӫ:�/L���t��:,��d긎v:c���Lx(^�r*��2k���uphGMc���X�y�K�������nX��]I��yr���mt	��^�����c���f��ZH�ۣL��e-Gt5`,�&vVݎ�Y������A%4�"*(�	�N�U���X:�Ѡ�9�*�F��ʋpVaC��m� �.�W)��g�Ӭ��+���cC�%��= ^�w��ow�eu&��)���/s;zi�c;y�l7�A�2�5D�b,$���Wa�FK}����u���V�ݢ[)�WL[-
&��+��2���l:[H	�
ik��)fӜ�rG���:�q	� rⰳ+�B^6�@ԩB�%�e�<}�oY��ʊm_2I�W��L�CG8��|��f��37F��i�!!S��AI�jpu�oR�E��qupct]:BM��4H��θt0 ����Cr�vg`���
�IvUK�����p�D���P�h�$�Fp�C��������������Y�[/�6a��s���r:V�0x�k��,.�{@4U�����b�A]��#M,TsA�n�'Z:=�.�	���4�za�O>����������ꇥ�B����%(���<!#rݺG�OK��Ԭ��X�W�5�� �P������1̻�2��r@���:��6!�DVQכ�6����=�r�����%7���X��U��u7Y֨���eK4&�kp����L��e�ӂD�o2�� %���т;[����^����Sv�H����h�G{���-��um�Yt`es�G�ם`�*[�/y�Y@�����A���F��M�C���� ,�l����������p_g�b�`薪�2p�͂�
��خ�n��E؝�w�v�cz�&	i$�o<V:uϔ��������ˠ�9�@��1]vn�/F�{����ی�#;i�̸ӹr�ha�$��:��%��B�|�j�t��\��Y%�.�uh��C2�Z���D���<�8�� ��.�4B�=��,gv1���:�N�2�˂�`�4 J\d�t��ǳ
\���}N%�Qx�<���.iՋ�eŋT�G5�%�.��Y�Q��%�q��7�Wv6��*���Aܗ��X�a� w\��U6����
Bj1S�F
�9�6+��Ou	&j��GPʘ�r�t�m�8���� 02����p<��wb!�԰R��#�c�7Sx�K��E˓%�d鉰)�{���QM7��%������_+���kV��&�x�F���&eay�Iwm��a¦[���q
0�Vܓ��C<�� Ie�a+��[�{�]�u��	n�H�-%�Wiu��m��3M0�;�w�lpT�Ь7���d�kӺ��U�KzҔ5�i:���9�;$���˝��!W�sso��sMQn�Rϋ5�%��s��";����KΗ;]ۨ�%�7ud�>]/UƔ�M�0�Ekf�:3G4�-i�,wB-oBͰq��\:���q�Pv�1op�]p2�L�QO7���p6N���Ԫ��ɦ��MI��.,Z���9��hG�U��S�F�:�q�ӸU�;�dmIŜ�W�p��tW�& Ov�Qz^�$gc1I[0�Er@źj}R�f�������(W��U�}D�R��/Foc�C^E]N��M-�����i�Bp����bW��w;�F���z��J��AnZ�3�NP��ēcX�p�(=��w[W�f��6{9Tcr<�Q�����F�R��ۈ��+�t���.��7{��"Gu�w@SOk�"���3��ه~��]�'k�'�ƴ���mތ܊�R����7v�Á�Y�8��.߅]_Wih�Z6�8�B���F������|�&�Wn�B��:���țrSN�9��m �jeE�+�ɹ��OkSCM�RˁEʌ 	�-�Hy����|iqQ���(s)�ڻOW���
D��8��u7��^.�s�R���R�]�K��e�cN�x�{M$*.ᛳdoi Įf��@S�'=�Y�Jإ����k��.��{��ɇK6�8�nvAě�s�ݬv K�];�#`���F�P��I��}���<�6?��t*����ζQ0���%/v������c���)#�؅;A�c�4��C)�J�M�вQ"��_W!���M�ִ�+�7/��A�48�Bu��f;`с>�J���σ����8�����3#���8��W�UAB�/�(5E�O����֍U6kW��?X�-s���_�8͂����qm�h��D�B��v�|��3�	7�RC�Svi�����+�v�$,��*Y�mN�G@�^�ط��|&�!�C�V�	Zgٸ�I
!�X���W6�f�*2�ej��A��҈�
����c���2�Z�	�/�2����IP�R�o�+[�H3H�tՎ��g@�j;���i���	{�V*��&���,���9,-v�R�m)+�.F�o	w/7X�׸s�������s|��Oh�J	��zVws�W>�i��ۡ��7s�������<Ͼ7��\j�$�	$8n�b�W�\h#���p�2�5KKMbE̘��"a�[PV��DQV���0�A��UZF���2���*�mB�h���R�H�FH	�5#��.)�Q3+6q1wmRћ��Z�*� ��)��ih��������R���v~��r���#s���̇�t*� �s��ln+�̡��9;��ɨ������K2����;�Q��Z�7�S{\}�I���.kQ7W�Ӧ�6��N��ѹ����lh㬼��}>6\u�}&Z�p^�CQ{9et�r���m$�8�Y������Ӽy&��������O���{�S�=J��D�Yܻ[ң���ز;]�l�����t���uNY���Mz]q�t+`ɝ��x�ӶӐ�M:��M�Ā���ey���b]��=@�^���;�,���Q��Բ^�H��3�0�r��9�hʻ}�5$��"��y�̄yyǨuL;�T�M�����9�דwVW���^�0�QVtG	.�C�Qu&6`�h�I�&NL�Cv`=y"]��ozfq��9W,�4�6�R�N�{�c�a��u��W'�O*�;3CUR���\�Å.EWm�ۛ/�K��H���{d9yiT�Vn�.�������<�E������:��mB&��>�����x�u[�i�t򢫰�y��kn��eV���_�-$��3��M���b�}�ZL��Z���J�ހ{�Q������&my�>v�� �ezi��y(�H:��2�accboga,�x欠�-�'���M�uL�t��;�"4�X2-��xg3��
l;9�[u9su�V��{�J*��
�-O}��iCǁ����K���T�˒�W��!��s�R�w>D��w
p��8&�J��	�*�XFh���D��e���g^���Sr�0�y�I[�G�M�I���}v���&"�a<��"��ĕ�6a q��X�b���%f5�	�v�Y�_�F�]쾼�=�q:
�u�|�ؚ"�wi���q�~"�m��X�6[�YY]9�(��R��k,�����'�fl�8���f$�J�^GwLQt<I��Lw4�k�e�ۧ��N���E1�C%�s޿/o]y�E�Z�T[biM���p�#9�P��t.�tv%��=X�Gj�g1�GUBru����'��,,�3P���{cΘ1Khkgc짙�����|�_�5�ꙫ�	;Ь�{5�j��X�w�ξS7����v/� ��[y�[���W�v��ګŇz�i�OMq�H�;Ɓ=�D4<=���B�`|qV>�S&��\+�	x���u8��-��ggu��poh��RB��<�����,�eW�Pl�ti' Q��؇�9\��5������%�\���1��ɒ�������R�K�rO��W�2>y���Ϝ��sᔍ�;{*�!�3���(�L�W<��Nr���j�.t�R2��#�D�k��n�z4O_m�#	�u2w�u�7�}��3R<|W�<���u��O���L򩈱Jy&�������j�˙����Dx�F���������{��&�-�V�����`��4��b�oW!#T��w�W> q1��I6S=�N&���.g�a���t�24�{)/��b�
Yw�u�n�� ��R�{m=`���������e��	�h�����`Y�
ħu+�����&�̉�hЊ{LH�����Uѕ��������&�×���'H����g�'i�M��]6��4� ��@�lB��1|+���8W^���avbT�Tb��.��p�ы
�rKe�����%�0̗ϥ��]A��`��+�K1-���T��.��V:�Q�wi��]d�{e��,㼅wnB*t�Fj�����ʁ��drO|)>^z�ٌ���y�0#�0�"�e���<f<�L	�|�m=�(fSQ����cu�kMfft������=��u+`�6e���YȔ��h�ҋFzYVC�K��ҭ��hא��T�Wè�;0�N�Z�XR]�\;�&=����>���G�:�/V}��{���Fk�X��h��A�A�40nǙ-�+t:�:���Uց��Yw8�5�7>��e��Z����d���Zi��h'1��q�Z�w�L<���=�2�϶=�D8j4 R;A�ұ�#9jB��M��
f�zn� �r^a��v3V��2*Jwb=�⵽��*ܠ[���uv�gy��Zv�u%��(���D9B�tCPDC-M�)K�'t�`��l�ҷ���]�ɪwdN9+�5���PՀ�-�kO�S�h�����6��~�}^�?�!���B˰	�x��0F!�XM̤�.��ȝ�&��;�,1c�12�*u!)�o��o�+1��] �4`�ܵyo⃀��I0�f��b�k2�,�]L1�I���2TL4�?d�pV��YE�P
6�0r��¯(�@�#U0�k!�s$v�p�7P��pTA|� 6j^
���/)�a�E�fO��E��KC%1W��4IT�0)j�Z[��&c�p�Au+�@�*ШР*�)����H��T�)ikiJP���H�p�*
ZE�V4EiER\���T0�PQ�ť�jbb���iQ�����J*���D�Ej��V!�5KJ��D��� )BM1~��|7������V�rc��]l%��Y�.<Ćp��� �3|�5���U��i���~{�C%N�����,���s��iu�=�5nI��U�'��t��~�����þOq���9�,�\�
>� ���#���$��PH�ⶍӖ��p>�-� �J�_#Ғ-y�M�&�s��QAt�}�C��ϛ�@����+�>���U�W��������*���~��wYPղ��,�E��u{���R�ƃ��j��U�E�x�Ӥ�F���w	�W�F��g�v�Sė����8�U�ٵAIM�;K<p��ȃu�(O9�rI5�M�����d$r�KZkO������(=�=ZW���y��%z�	嚹k����5w�M���j���Y��=v��.'�[�HI��2��b�KNw7�oM:[f�{�	˺Hz��ixLȧ\P���w�,��'�M\ �e��Y���u>4��bno������>���Ikm �k�]�����6_8}�S(�L��'(��5Ӝ� ,��R�%���yqR@�h{׀S!z����;T �"��2��u�9�]�5�ܐ�Cw���!@�@�`bm���P���ׯ� ��������Q��S�<�֖5{��w���k�>�}>���xLz2c�J��T�V\k���o&0b}�6�4VR���&��Y�@2�U�D�+-y��Q涕��Q���g>L�� �
e�p��`��B��B�ˏJ+h��A�+]�{�}��e������������%W���El�UD�Um �B�ho����-�$������"ȴ���m�8�_5A�(����
��g�o�Y��s�Xj�W WR�ю�ʢ��T�Tv������H���UQ
�UF�3��ڪ�!�}
�W8�q
�|�h�Һ��e+h�ģiV�P���q�1�_8q*��-U�8�h1�
�Tu�:�u�$B�}+hQƃIU]B4�����8���a('�
�UZG�<����T���WP�Z��GZ�����uA��إ�x.0m�T��T��Tn�)@�T_�A����{�~��w
RQ5��c&���y+k�������Ƨ^��+���Q�*<�糉�����9�m*��ˢ��*� �Q��R�v�� i�y6�W�GR��{�;����k�ߪ��i��A���q���a ���%V���A��(W�����ms��;�5�R�-J��B�J�{�R�q(5G�UG���I_ �zoOf~��W�R��
:�DC�q����\�G�W�*��A���TB���Ҿ��ϯ��ª�)j��h>�kM|��J9J�@�Tm��Q�%S�s�}�y�4�M¨�mW�^J�^j�%M���Ua*��UD�+)U��'g}�~�v��h�Ҩ�U�@>C�Uh2�`�QGNZ��UԪ/�����gX�J�4jU&�!�87��ŐS8�x��4�Fڢ%h�a����UQ�ʮ%V�j�r�:��IUXj���i�_%q��^���ouԪ�VR��Ua樈W�ʣmV��j�Y�\@�EW�YJ����ϵ�o��}�?ƿ���4�̩o��:��pN����r�Mhڷ=�����i����+�UU�V�*�����A���(:�҃�N�JUa��Es�����%�uQ�� �*��a��Q9(�A���J�
�A�<�B�w�׻��ێx���}(4��
�Tj����(P��뢈�P��Vڥ�{�y�
�WP+	U�h�U[TQ��4T@�%q1�V��ﾝ>�{�D��
���w�--=���b�޻�e�TWR��R�tMjs���C��z�-�+����Kv�0�;�fd����o�ePN� w-�m(ޙZ1vU5
Y1��)����%B����c81���:�	�vD7��]�*3��9eFtZQ��j�J6ў���8@Y-��io.���0�H���@Xf�c'
�~�B�'��d]��yn��@w��O�R����p+@f���B,̇<��%pr�[J�A콡9n���r�ޒ�v����7F�N�A�I��ot�ȼm#�|�Ct�b��Fo��k+�}�-ؿ�&}V���q`OW��/;��&#��� �3�{}x����������G�ˇ�)��l��J����1�=rx�Ӓ��.(��&�V&D�յad�b���4�c�֒n ���L�+���XN�Oۛ��-�Ya�Hwf$�l7M26��3��U�4�׆��Q�R����|�,��WN^��7=��][�)�Fa�ڋ6����F�6m�^��F�1�����pi.D<N��K-Z�͸�[
;Ӽ���x���g�{��dܥ}�	�� �S�xo]wtͼ�;�Q�Y7;Mtot��muPl��^E{!'-/9����ޭ�6"�K!M��Ĉ㓌%�����"��5��Ju���h(*���Q�;� ��٬��)����:�Fx�i��H�w��ڇוW�*�w�ط,GA`ۡ��RB�-����#������(NA�}�9���;Gp�V��$dc��V�(�0�㘠��z~|V#n�;.����K��b�`u�뮟�x�^(��'�����i�'^���A�m�hH�+��k+�gc��i�"*8GF[p����䳗����Vm6�>�}����[˽���`�nӥ]+W�&|��=����T�t�@'���Q��E���l9���t�{T��o%ۚyX�|�ݚ0��A�!��̩��v������m^朩;��.s �<��$6F�,��-�_�IA�j� �KFS�ߑ��+u�PH7!<��l<F��s3Es]r&P�j�8��;�yZ�ӻ�T���1��6(��Ъ�H-m7{ �Ҝ֟X�b�l����^�0��=�Y4�>6�YY���}�����k��խ_byl��+��j�3�ˢr�I�j����3���K��P����>�Yme]K��'�t�T�F�[��X�ʓ!1��VC�v�:��vY��E�4q�9N�"��bY�Va&R�*�`��YX�K1���l�(�ܲneȪ�t��aKB�I*����k.*5UVnS��ꍤ��@Fi܎f�}�Y
�#u ��T�q&Y�Ir�1+YD�c�Yx�:YqG�r'xK�1\l��7��uj0d�;�kvcoy�f%�o7���_�'��A�n
#�P���J�ZH���LJ��a�!x�.ڶ�nF2�,K1wuH�E�*�I��m��D���B��؈�AZAEp�q!*!)$����R5�B�%ZܔK��bLD�5JA�H{��9�sx���g��;s&��g)�P|�g��R�1�g���Ͽ��E}Qg�ciժ���bq���õUe��j,@�H��>ha�g�ʾ��'d�#����h���tȣ	��5|��u��Y[XY�Cg17����E2�7�IĞa�5�ee�-׼�nZ��B,�7�Mb�ك�}"�����Dp�J����F�0[��K0H%=u�s78�˃��wY-7#��=ڿ�F��*¥���91S��Gak6Q����E��[Ov66�{���f����B����Q;��8Kel��d��}��^86,f#.�0:Vv-u}�a�ke�٦O�c�����vc���p:cnЊ�H�7zwF�÷�w3~n�;ݔ�QD
\|�L�%���$�q��X�VޥZ���ׂOM�ØAI�w��K��&xx˵�����:�$�g��N=�wJ�#���|Eڄ�8�d���-Hi8�������#�1Pa��y4"(e�Y+^��}��5�9�zFG1iVv���.��jS�0�k#�Ý�Ʉ^�Bޗ��$����#��*�Vt�����mE�%�>�NU׉��V��_9���s�W(�j��ۛ�h^;S0%:Y��H5ۦt��s��sxN[��p�{��D,��i�����~ߦ�n�NOT7`��W�/P�ջΐ�Z�@�v�m��0�c��'�o��~e�;�Q^M*
LdϠ�65]�����;�$�����ƵxG�ұ�"�WG�
:�ћ���e>K����߂��j��ɮK�s�<�$��p�<�a�w�v.N��y�K+��d��VR#1N�30+Q��Um+���o�.�+q��ۆ'ֲ.ԇ��+�{L�Q����s��/��f�������vǝC�Oy(u����_cr�R)�|u���L��I�Mg��>�X�#I��o���:I(���P6p���Ba`oR�g�jƓ�t���B��\rr����xQ���MN�:M�K8��7�U��y59R����E��-�Gj�SY�Z�iT��Yj�I6�u��fh|����A��W�9:.�S�Y�/�kt�\(����y7ӭ�v6Ԯ5�����Sm]pxz��7�v�pe>(���� Y���t���z�zH����U��X����m��6W:u�IK��y�+������K�S��"����SK�:Hb�ٻ�`.�"�֯�N<�bYXOVL:��kj_Z�/��EA���r�T���rS����G+�{�舌mWV�/�=E@��!m�^�hd�;]/��d��Ac�Ήr�^����<2�#&�S�dbPo:�2����s=�W:���W��fkm���|�G��Ǝ�wMi��8���Q��:���wZ�	&�x����,fL���\gg`9@RDuǾ=���w�Yٶ/7���Վ�.��FY@F/�P괩&slΰ�y��{����4N͗l��UW��L�P�S��<2��}�DG�	�W���&9l�C&k���V�yDe��j����k�����&- tIm݈]=��s�&��G۹���Ҋ�o��\Uq��i���u�J$`�{y�����w��0�F�ڍ7ޝ"TZY!*L�{��N��V��;��^U�1p�����vfW���n�x�^�mp�Y�X�Um�F-�
�NҌ�ZF�D{��:�_�c���ͣت#(�h/���9.z�n�>���Я,�Qk�%��!�a�C�-9��u�Z<DT�Y��Jm��%��:kvJ�$:y�õ�����Zh`1�����eu���'Lů�z�w&ݶ��FgW��%���[�r�@g���;޹iև��zt� ]{OMD�t�r�<�r��̨���m.���_z""#��>�?@�~=c����|6:v�K��%��T���Em��e
��V�[.��̅<K)�]�;Ȓ-�������a��MW���L��H�r���Ćy����b��en�,�4X���[H��]f�.;f��f�w�~嵅�6
՚���J �7|c��0W��Oh��x(��*�Y�ʑ��ӫ��ŷ�]y�u��ޭ�}�v�K����q��w�9d!�\�ma��%sL�oLU�DAu�pP��]%�g�R��Ӫ�m\�(%��ݘ8�0Li��\�3���֋tU��m�ֲ����Ռ��a+��ZgBА30�e��6��HΫ�mu�.5kR��P�����,��Cг��U`�+�.+�Z�R#I��}��Vt/k"o@ȏc]1W$I\�R���'u���S�w�i�[nF��������5�
�ǮQkM��$���d�U�tr],�$PɌ/�I��l��J��P�3L����(�A�a��b��]�KcE�b�\V�����Xp&�T�Ҡ�q���_َ�2�L��%L���1RT���",�B��fb��Tn�^S(�D+d�#o>Y���T�N��ZCU-ap�C(�Y�&Aݼ�(a�YV����p7�����T�J���ݲM��`���T�E�a�H��ܢ2��(��YZ����t���F�*(�4A�1	��#%DP��Qdؖ$q(��i0˃)��il�UUiX�QiZ�#PY���ҫ#Je#� P��{�/M�O��s/��B7$o/y���}U��_%�����������=�1��5ڠ�����+g]է�DAfw��a���t&����a��ۮ��Lˉto`�隬SF�`��c��
���
�݅y*b�3��hx�<����ך���%����z<p���IF�<�m4�e;�Okxy���Yb��,h��F�����=�ў+1�d
��_���i1�ymH������	�N�r]6����̮�/8L���We�Vz�N�ama[�Ǡ�5�j:�����,�[��ࢊ;�e��������5���y�X�V�X;MYx��HW����0`	��h�!�{w��:�&�-�O;����'i�p�Ǳ�ç�RD�^$m<*�^7O
׋N�S��A�W|�Y����M{N*���Yڨ����Ӗؘx�sx�{��֕��NC=��a�҅T�vj�;��C��T��+���b�ۺR_=u��"�|�4�E]�͏
���?G�b��X�a�B����B�
��շj�d/7��*�}�smfK�j��3.������������"�~L�W�J�{;����3齛��1�?hا��/�k�-�os{�yX�4��ĭ$j&;�R��nېY7�y�6�S<)\j�0X��~JϽ�"��P�4��AN�්�L�U�_@ I{ܸ}[9|�p"a��c�Ƴ�U��>�#���h��C�**� ���6�����4,u��^�@S6i�R9m�2C����x�L۱�=v_�Ә���ƍ:5�n/Z�-Z�r�6+���W�Vt~?;�<7/x\�|��kRr��'e�a�/�L�\�� o���R�{X���A?UW�W�o���O&�8��['��z���f�k�];h�Z�lu�Z�69v���{Tŏ�h4>���x�=4p��#��>�{>�hV�)�~B����b�w������Sה�i�{<���:�蝫�o�]��m���;h�^L�ͬ>v��k��{͗�m�P��Y&]Q�.N`U��)S�����ɇƸg�ѭJ����w3��I��YD�@���U��[َ�X�>�,|T&��}�ɡپ��6�G��B�j�ٖ%X��F@Y�����ft\+�pwGEj���._G�=�:���>ԩk��ڵ<�t�r���_�s�\G�@���Ы�����0X�;�J��-K��䅇�U,���Kױ�gq�kոd�n����N���Ǌ̗ۖ>�8(����a�8��6N����-�L�mF��8�3.�<���9�㷮�-޹a���DܙE0���k~3ɿs��Y�V�秚�4#Uճ��3g��͏�O��\	�ډ����Q$C�	��EG�b�X~J����hwt�7�D5�wm���`6�%պ�k1�	N�����ɖ����;�.���W�+�v�ߺvj�y�1D%�H%c��:�H�y�}AUF���^=r׆��^�;��י����*����pp"�c� 9G����P}p�R�W3꘳B�[mT�!b������*��a���#
\j�*U��*�Q�:�6`C�Y�����_]�V� }�=���c��KɗML���0��{|]�M��J�m�Z�a�Ǧ�9p�N�x�s��ѐ�,���A¼�Nɧ�7O�5��1�&
�*��X���|of��g�4`����ę��FI�5*�l��O:p=o�ުcf�C�6�꯾��9ᒉ��2�3��X�>��|�_wg�Z�E�]��ڠv����@�º��V8S��4u�QN'�&�4����b���.��c�<�M뿈�
������u�Q0V�����x*�5�*���V��Y���e�!�N?����b�U���<}��w�����q8�s�X=j$�
GǕ��{s�Y�f����Mgf�z�ɜ�&c2�������l��9��]S����CY��dy2����Ɗ0p��QU�n����1C>�vy}�s�Ѝ�OK]��0fԫM����OB��!	Ǎ�0��ϻ�@<�y��ޡ�-m˧�R�'f_����>�·Mw�WP��a
� �a�W~Γ^���ۇ/��=6�u�]x���N�(
�4ׅ�1X>���0'qLw<��kO��K�j�ɱ�Cm�:�l3����X�~�>�]n���� O����r�SUXc�A�<kX4.K����]���]�0UX�43<�W�I�h�;�`��sR���ha]L�+͛��#���ê�yj��ւ ��HV
c���������d�&���˳)9k7C�q��O+{w{�: ��:���_V�X�=79B�����֯�xg�Z�O����L?o6r�t��^��8w.��-{� �8�s��N<5�b��pq�ZW��a��r�0f�3��>n,T3F`Lr�7�=:�21�z�z署�5s7ĳ��P�� `�Fƅ��n����`�u
���N���F����oS׍�9vX��wzGO��f�75�d�㻁����p�_�߃�޾���>�����*]�� e��cV���b��Xj���`���ʮk����"���63{��Sc}ݧ�k��8�K�g炎U�y��Q�Z�����[]�=/����M�hӗ,I��y�:N��^�@���9���-T��v~�63�o��P`��~�r��-ƒ����F��1�4�j��+��1KMvz��;�{���-��mht�bi�wf}�9�F�Τ�<q��NML9��ʙ3�좪�ԋ���ZxUv5LW��b��c�т�6|K�5��|���X)����5¬
�u�zi��CQ��r�>�`���RC��{+�9*�z�!`٭<6#��X� ~���6	�Z��葝�,o^��|s�GSf�6=��OK��e]��u�ݮ�\j�,;�Qg�ݣ(!ۼ_��k �9f��ɒ�^���:1��O�1����2�?��sn�,K��7Y@ۢ�ñ�j��Օ�q�p����@������D��ҩi�hp��]�[=}MB��efv�;W}&��o�ua�!��4v2�l���`u�#}η��uq�&e7͗�W�O�%�L�ڔEj'V��u��%<�z.�[e5Xf2ܹ{eb�뇃V�uj����.aR���Wso�b@<K(���c��bT)'L%p�BU�{t�2��Tԝ��gar��I.�Ye�����
�K�+8�A�c�d�8V�^}���t�6��oYU���.� 4H|1��r�:�QT���}d��ɚSM�}ګ9���tE���+O)��]NB��V�X[sv��1H��T�}��*Ϗ��=�s;�9�Jb���;��ޒЛu�q�7FR��9���Wلur����J��i��ɜU"s����w	4s��w]���R��DA�SK�RHƅ�פZ�hUQ�R� Ҷ�R�!)U$!�-#lh�1�"����Ҋ�M+P�b]BIZQ�FITIJ ��E��F�H�0H��F�*A�#$Ĉ�[1"[ZE�Q���"��*"�J�D��H �����ׯ��^��6�
��ڛƭ�磌�Q���W���:X�#^��A����\B�U�.6D�Dnv�������
�D|`
�P,ב�����9��O�W?���|�¶�����m��9�ty�pr�J4�\���tΘ3�^}S9�9���㦧��)z�w�؆};�wP^z����'�V�����ge�y�����vkPS\�����&'w�X�x�N�xֆbh�����¼=RGLW E0����\N9��_���&^��>� z[�5%��2���:���2�L��ӗan�륪��e�M�,�C[�����/r��=!�,;x,�z_�?��}��&\�;;�V�[�&h�b߭�@|Q����@T��6,UDl_c�Uͳ���؀t4���-,M8/Q�{����}��tr�;�e�e��9z���K��Xv�L5�
��h�6h����jc��}ޜ$��ϯ�sܵ7�q�B�j�7�}8��N�rm����{r��9B�h��/��=癵�����Vl8(q�i���ٗ{�o�x�x�x|E8P�4��P�u�X7�����y���P ��R?Rg�N����ii�{:K�ߪ�}�ga@s��O����W�չp��).v�m�K����k����&�y5���ǩ��������w9��i����E%by,|��ɜs����|pxQf� >"���4Nv��DX���f�
��0}E1=�9��qu��bǮ�;s�OJ�!�۪�'Yw��
���.���ߕk8,V��.�ǗPa��`�����lךV��=�
�4z�J����Xb� �_'������XlT ?�,x}�y����e,x�|��:Ǭñ0�d7����F_L�0���]ɚ/��6ᮼ��������\x#2�C�[x�%��s�o�
̽ﾯ=~E8���ʼk:��o��w��]��S��([^Ore���ӏa����e� �OJ�q��t�����SI��+��C`��N�P�a�͆���V0p��*�X4!T%���7N�|݌�S�
��&;s�V�M$����=t�s��[Z�^4���(t[�32�Rxp`3Z BW^�c᥊�xz��ja�#��eZ��Y׌׳�7��U��o��P�Q�T6���a]�.�E�*9��cif��s���b�,;���)J�Pw	X�ɜq�mN��"��}�^��Ӵ���y��!��	i�ɧ���7�ڶ{���=N\*��|��)�p�ʧs���F��v��o��a�K��L�	��_zJB�i����Ѭj����h絹�{��]M5m-��K��W2��cÅ���ADW�S�&�i�y۷��,�&�4�C	�_�c��T�b�`�5�i�.�@kMWL�nſ/����~���޵H�:)�k�D�^v�s��μWnNA����/%z�ˤ>k��3㹶XR}lua��gE�͜��S:r�0w�_Wվ�w���q�����eS:�nq7��?C:�3���0����^�L�S��{Z������o�x_'9<�y4�.�=kɌ�]{N'rw<�+iԍ��-�9̊ul��;}s�iJ~�.6}E��SS���;�������1��>�]�Ʃ��ϋ+��w�����g��D�R�'a�5e�&��=�&�=�V�#^��k~��br��8�:�6�0�#��R�*#@|�i�񧸀�)��B�� ������z��r<=;���s}�p��W�pE���۲����"*h}T�Y���k޻-�w��&����ps�i�V��2����q���h����wX���i��6�<�0���μM���)7��g�4|~�����Q�K���n'��c�8�9O5�2ן1��L`��OkBޅ��:a:�uL�򉉆�4ǅs{�o�lup�������U�����ex�M�{�wP����-�!����kƽ�Z�ʚ�U��/j��>�5¬z�H7���b�C�]�U�=u;t��#�w�QƵ��c2�V���\�t��E��
V�-���л�L�$�f�b:G._DG�	��>v����,r����5-��7x�e�p�sS\���W�4�2l�x��w�f[֢ML���Nj���i�z����[_AZ>���ШX��Le���2G؄uY��,0V�LA�E[��X��"���V~��^G��0`�N���`u�Z͂(���(���#8�}(�����W����-4�t^8�;y�]hNvy��W��m8�nI�\��i7ɇI�TK����1���* ��w�a�Û '�+���*�]��Z��P9k[eHd���(^�&M���#q�/w�S� ��}�h���N]jV��>��Ԝ�7���sg�����A�.!�f����=xN��	lr�Jȇ\'%;u���u���r/�P��b>^5������<鏱�)V��5pa��Kytk$�<�SN[�-�5��2�k	��Hy2��[k�Ֆ֮U��Y����%��������?+vm��2�y��3�u�8��JP��gRO�}�g�}�q���V���h�JB�<=����Λ�j����Y�t���5�|F)e�����K�Yݹ���]���o����۳��H{P扤�K�5�o�}���=����u���5�~cE{�З'b���A��t��ʶ5��{��w��/:T6Ѧ���\-��� �]���n��[T�U����̢���{�;�iϜ�����t�� �[7+)MӶ`���r5�j�@ Ǉ�o%�m�@{�_�b��をG	�>Ap���&]�z����슥��%��H*��;<����:�X�)iѢ��axՌ>�Bqؽ���5^���e9�͞cr���X��>/�[!��ǲ��`��u��.̕�Z�qs޼1I�5�-@9�z)���\�D3e�Af��5���<��	v����n,�. 䛰v�VFV��j�ַ��u�WLsS~J�Z\�n��eIq>���nEHl��]�mY��Yԙ��M�3��YҒ7�q���;Gx낙����'GM������YX]^��EК�
�r5���N]��W7k�gJ8f�ѽ�N�K��K���=�-/�s���Py广cxPuؚ#��Ȭ�'�pv��]�hO]㼈\�4v`Z+v�9�BG��|a��L����u|�l0�U-b�oj�+/�B�l1+�+�iQ$��Q����O
��q.@��&���dj�V�͊��8�a�w����;��AjH���r���wj�	�9�I��-Nf��Yn3���0�A�����^$��.��Qo}~h�7�S.��f*dr|j��XR��ٳ��E�V]�@��¡������vX��sC����3�M���(����o���̒�<���ջ�;��.�������2Ev�opD�DF�U�""�TAEd��TDc�J-�ؠ��܍��L"�(��8jT��

�b-("ܫh���7iEQ�FH��ZZ��EG	
Z��T��0�[�*H(Ƞ�A[H4�KmTij��H�[F1�U�Z*"Ĩ�)!0�K�Q�?����q���=O���]트�J�G g|����rI??�[M�O�<��Hm�c0�k:�w�wV�K�;����,�\�e�*z�&��������ۇ�9k�]�iM�{c�i6C�
���a�#G�;/�+?p�� (邮�F���bY���|�\�SHud�d��a�͢ׯ��13˘���^$��؇fV�C�s��2eۇ��Km�mk�������+��n�&��p��0�=\�w��f;�f�>Nvpk��氙E=��W�_�5X�����ڙ��&�M�q�wo��jd�O��K��j�'�����F	�WԽ��3�y��/w�0zw��&��ʵ7v|�:�r�5�[�CLx�9+Y��s^���������cC�T�±�v.��~ٷ�Ֆ�\5�0���K�9��v*q�2�W�Tw	�O�`NLC��}Y ��w:ʘ�Uθ�Cb| �g��z���9�T^c梮*Bp�'���ne|.��o�}حL��WFMn�d�hW��b��>b�Mg�	�y�)���*B�8~��*���f"3\Q���J�eR�Hh�O�	�1g��B�#g3ѵ^*��!��7���)L��WqDV�
^�q��}��.�Fʚ�/����׾���Yt��,�s3,E�h��\_1�������+�M��VV�����]�R�6�T�ۺw���p�w'Ng��9�S���j��'=�.���v-�>��ǂ������Z�o�[���v�j��y#�N8p盳�����y���G#�vȜh���[���m��X,nZ��?���J@�ʼj
��}e
��e
��5PW ��z���p�0xT�|���<)�>`�~����՝Ѩ��UM�����"��"*0(��޾��\�U`Hꊟd�x�՚�jCN����4k�8�bnJ���cP�Xr���{K�k��&���bmJP� ����fyߡ��Si��6`B����¤����Ռc��]��8�4���s=x�x�+����!��q��p�!�}�N����W\1��̭z�g[��{%�bk��xy�y,h��j��YXt;غL��k1Rf����C��LP�;v�;&�����`t�<�|�291ǝ��cO)_�����ۛA%�p�����#Ӣ��1�������r�?��bg����|���|���>՜L��>O��\v��N�w�ii&�����;1�{�=�u�{s�~R��Y=��x�J�+ۅ�Ԓ(^�o�sl�j�kA� +���g��3�)�gڀX|��\��ʸZ��=�^�愾�z�]���X�j�D5���U�[�;g�w^sʚ6-�+��Ps7��%�aX�n�ry�}�,T��n�'j���߾�67��Wu��k��$�Y���m�<�U�nv��VR~��-���R�zF�u̧���6䖅�tdQ�0�]�{3�h��<[�8�x���IW:݋Y\f�r�!u,���t�F�j��x�Iq�P�p��0�a;�ٗe���^�����T-��ǜA�u�<�ˈ��w�mx��9��� �Hi�i	�4�����>$�U�}pgK�bR�������}�ν�^��[�WӦ�3+#�ؔu��f��[�c��Qf�5	��$�	��f��q�x*��qx�v�Jd�~M	y���l�X}�뜔��,��뽎*s�6Z�_2��Ms1������~Hwݹ�x$�j�g6B������l�յ����ݾ:�!���=#t�buo����Ec���5���Ja�P�Xm���h�st�4��`�����! ��v�7ɀ�u��4��#sS���
�vW�_��$�H�_�m�kˉ��A�(�m���l�n3V]PS8�ܷ��.���(���Wx�J��Xhg�_�Tڊ��8��]Z����Yb��u	���s�L"��ݝi�̽�k�h�_Lc�L�2�E��U}S7��]�w�U�wX2�\5r�M��}������L>�pe].&�l�4��n�fL0Ԅ'E�l��z�p1>����Z�Rnف�ĤmIt��{-�r6�a���p��3��
A�Eո��FOdWA�<�<=�N�je�[�L���(�h/Xkq$�RC�y�D��Ӭ壱�x�t�`PN����E׽.pa�]꯫����ᰥ��.M
�tk���������.{6�3H`���n)�U���s+�MN5�_F�x��Wu�K�Q�L��WƦS�Զ��$d���
�tn���f�����Ks���S�Q\�x��
�弮��s�Cz�����4:��$�VnC��^V'���Uo*�F��5�9�z�}�A�\uK<v<р���]�8�/�;���qK��g3�9��I�����kRs���CV��h��shJ����Sv;&�B�1���LԮ�+VOY�`��w]��\�Zy����ۄ�V����+����ڍ!�kb*8^�x�^�o���M�
�Z�R�&%��-�	ɷ}h�/�I��g+��7PP6��'���M�q-; Jav�0�2�k^�Բ�$9*��d���e/\+j��V�ڨZ70B���e92�Ǖ�cv�t���*���H�B����w��uWl'�/!�n
V.^U��9b�pڔ.�È3�&$�
�42��*̧*�7x��b���gӰ��dVER^I��(DI�?�"�Rh�%��K�e,w+N�Z��0��D���[6Kٻ�����E��`UvN�
����X�r�!H�\)ƩLwX�*�!yf�o:f�r�UUMĀ��@Qq��B�ĉ##.�"*�+��V�bZңKH�i-�Э+r8jbTY�b۱��iTQ���Q�H�w��i.��Ш�ZK�*$��]ZR���bD�]��.���5$�i�AhI,�[T��^"6���I-��[l��wm�Q2H�F����[�cS�˝wBv�.`Vh�NH	;{iC�&��Oz��^)�ἤi��R������]�d�����Dr<OG��y���Z��F��^;�a`Y]�I�<�*ۅ�z]�U�O��:�"���&��ޗ<i�LY��5�J׼�'L�>�.dI߭+4i��<�ԭCj�%��\���G�^�K��J
Zŷ����z����s��{��o�$/к�qz�y�/�ڡOi��5@�.i����?��j��_ڮ3yg���P��U��[�U���|n��ҶV;e[��f�Ǌ��
���v^�Ð<��7�n�
U�Ќ�펹��L��Ui��_a�05<��{v��OSS�W.�fۻ�y�6��×���ױ7��2�5�K2䶜��7�1u\e����x�C��uib��9��Ut��BF����ƎQ(wj�"9�]ߎ?ދ0HV^l�N���!�3&zLMP���D^j���8���{ya�3�dT,ަ]���I�������Rr63�tj�^�i�H�9�:Y^�0Go9���H,d�cU�����s��}6� �>Y��#�}��+�S����G�J\��a��5FT� �F���D?��.���$��(��9��wt���9٫�Du�$�Y�,��u�m������ik�w<*�q�*d�G]��c;T�=�/����6��`*���l��+�׍�Ïtu���T����TP����@U�e��Ǒ:"X�m<��Ա�]�mtLЬ�ۜ`�|�������{�����Cn��E��,�ft���0r��������@�Hu�Ўq�e������ϢyJ��c��tlz@s�OG*�2w9��8F=����T�[5;���/4�#�E�C�ؔ�]��+��S��ǭu���,�E������`�\e<4@[�Z�����
��DSͫ���A�.,�g�CQ��H1���iЫxp��#��n<n��l�pd�o)kL�>J�B;�M5Er�Z�y���{פ��:$JԷ+�,�7˗ވ�MwWg�bݎ5��u@YVQ����5�0ŗ��g��^���T�@�f�&9�*i�����5�҂��W�X&F �x��9�c��E��}1t�aH�����>�륳�(��^,�Y����@ނ/�]5�6*�w<��n` ��i9"
yH_���Z����U�@z�֥�7���;��os�WK/��y$�0C��)�,b�n~��㳨��]o�@�.�qSC~�蹌�3�<��V���K��8Th{���I�K.�v}�dߞ���ە�o�R�r�+�p�[�Q�٬*:fK^��īz��raA�j��z3UF�b��������g}W�3��q=�z�p��_$�|W�{���x��MӶ;��-�X�BC�g��UʺH��d�+��}m8�?����U�|o������۾�ؘs�ֲ��X$l�M������b��c�c�F�/>M��nN��g�r�"zn��Kwũ�>[x(U������.�L�2�ʑ��f0���������`�������p�u���~�r?Y��΋��4=:�i��^X=ʔC2��P\�m�E����(0� ;���o��oP�7L�ƥ]� ����k�Qk>����QJ烈�-9`��m=WL�)g��wX���:�Ր;½O��-e�~Ѿ^�>~4R��|�Gv�^*�M��yq}:J�*7v=�`RH�$�%�Y�b�0J&P��ӜrWSaȅ�m�sC���W���&�^R۬)��a�뜘@,Tިc���C]��:`KmRW�0<��A?}UU�'��Z{Y_��"��ݘ��c�P4MU�kE�=����iC%� z�i��7���	��ˑ������q`z{'>����y�ذ_���zG+<��O�30,@�:]$jz׹ ��lv��	��z,8T�HA\���Y�eC�����*T$���6���o��7:p��e�C�,�A��[��M��q�A���W��+��n�xdn+����M���z��tT�����9��M&ǳ/<Sz@x�Z���8۷��{e��"�`^�oauo�[�6���qkK�իa�;ƶ@����6��-��޸�Ȑ�cY�G�p�,K��a,��|�'@L�1�-[꩛�f]�]2���M�wō���~%��h�ݮ";��,ctH���-� Z�yWH۶1$b�Y�B2�U��b��M�0bF�L�ı"��fY�h�VVZ(��Um����Hb��V�T����YF��Ѭ��?p��]��U)�Rf�I�C^6��7�2�i�x�m�ܺb�TqZ���@Х�TQO���X����@�����t��%f�0j����Y�
/�D�I���0�ر.��L�Ӥ�YM������+Ǌ&��a��|k�(P��H}T���l�]�ȳ	h��P���J�Br�2K�P#r�\�6]��%���K4�E�1,ĹKlih���e��kuRE���U)n�V�Ս��r"2EZR�R4�Ҩ��-F��B�	0��F�*+U�]�b�iwDiV�c���d!6��Z��D\Kld+�R�1e�#D�H�>�*�D��([��wַ6�)C%��p�s�:w�������R�da������[�qx�Tr����Y0�V�t+�*r�v2rT�c��<z��F#L���<�R�����dz����`-ػ@�6n��Q7��d�l�
��&�ݿx@:��ȋ�� �u~�(��:lU���[�d�c�!�5A����h�]�B����N�}��$aIԮ �#yc�]?'{A��� T�i1��S����b:�{>vZ�ˌ9p6��kTb��#��/2>ǑV��Q�n����6��̓5-���QEk�/�������RF�ף�)�v��(S*D��ZyْK7=&Ͼ"�F�k�>���&Vi~e �pz�}��2g�qɹqF�@G�m��{Y�tQz��nN�:�ڭ�����{5����f�==L M�Aa6�p�@^�4�e�ҫ��e^�U_%�#�G��8+P\����v"_�3��VrP��fZ�=؏\~�Ԭ(}
��vjܱ��x�ąTU핂��3N�m8u���/i��4«Ί�u��_w�s�S�"�9�c�8;���!��^�Ǆ��چ�n��F�gss�P�{�.b�YҴ�R��s�wZ��29({�w���0�9�Sx��¶T�< ��;/J��O�Lb6�q���xGv���þ�N���+�u]{U�G�g���pT�k����7�-�o����
�)�F�+��K�Y�=[%�����e�%6b����B򈖌�/,�*��N�k6:�/A����!wtu�{v����9��ع7��0%-�=�>"��~��%O:�ɕKWd�>x��=��חn��q���L�[�b��-ŇJ^������q�F���'[�څ.˦���iSc<yV�q�)��0����,���\�[#t�A�WP�5���J���fEd#=͑�kN�=�WV#E��Q�8��(x���
��6_��s���`P8�'OJ\�2J��DrR�����jV�y��w$k���,!��'*�����:xR�.���%/�4^`c"���L�ӡ�F�C�U3a���\.���S�Пx�A�*^�����O��%�����A56](��X���,[��=�v1�˿�af
���f���W���mU�u�Ћ�P�l��[l�-� .�qV����1�K�� ��ywؚ�-���E�8�[�ԮF����.Xi<��r^� > =k��\�)��PB����v�!m��^��6�N� ĝ����΅hi]��4ܘ����=��^�T1Fx�y"P�NM`���?����_-�q���F�lH t�u����J�����(V���IBf&ɫc5���7�v�'Sn�uf�Mn_w0�o��S���R��ٚ����;+v��(��8{�(��|�NQʵ�I�ƨs\TW�(ޤ��-�l��&4�}�V�ۭ-dtd�[�G��˹���s�w��[��ߦ������z^}���nq�g���������uBW\��ۖ>i��^�%���:3Fѧw�2���ܹby�l���p�aR��\i�)~�������͹:d��	��ʝ-��(�2j���aZ��^4�̋۞z��V��^��������/��F\��{$�r�9�aK�Y�>rևOY���S��Ƶٙ���5���0[1a��^r��e�1���e�z��6f�Wc.u���n	�b%���Odݯj��]�v�ٺ�N�Q���ȓ�5�jم�а�� ���g���ӳgyk4�N�Fⱋ��:���;���hs4���"%3������{�լ����ޑJ�[� ���I�!�w�b��&�T�����j�w�'1��|h��Ƨ�f<��]z�O����Wo��5mze�D)��B�;��	]�<��#��ɞ0Vc����R畜yE�.N�o���J`N��V�e����v7��EV�#6�)]���r�j��4SWN̻V,j���.��Yk�E��+�8��z	j�=�Y�rΡX'Wj=��gգ3�"h�MO�ROl�ѧaqY�Dg����M�p�s�oٚᖱV��̕�T��G#�s/^#���r��ϖx��iX��6NA��h;�:%�����5o�Lʕ	���/M�+�"�vp3n��)��M�=o*�+���1w����{3�W:DU�g	}@\�)�U/egj����t����N�&vmݣw@&d����by,�\��`�'I��!�蘧�'���G�,�`�[Lq�*իM̺�L�,��1�j1�ѹ-Z&嗋(�K ��WU��� �π&���гP i�"*�b��WvD�\��3�)B�,����]^K��Q*�W��H6�:�'q���+ʫ���V]]�"�����"�ln�CPq%�0�x��!�EJ�F�R�%4�)ie�D�Y.�V䌨ܻ.S0��2�J�(�Uq-�[U`�4Z��
�8���
4�J����2�B7.�4�+��d�+�"�����Z�UY�DV�R��e�KZ0˻�*"�iQ"Z\j*��ő�bh�U��$�����<{Y���*��:��'_�����2�������L�tکA���ѡ�o=�����{y�]��[��)>���y�	 ����+�B���{�����F�խ%q���9xW���SW3=B�A�w�k�7C�3Ez;�ZA�x�)��G݊�����=gl+���l)�P}:�`��0�sGXKiV�4��j�Bvww-�7qj�X,�'8�Ro[ ���������]/���x����c`���a`W����q��׶F�νN^�9E�}<�vס�����"p�ޖ�c�-��޽ױ�	��F��AWמJ�hm��<y�1Re�P��m����\�5��q����O�o�ѹ]�҆�	�N���\{%��kOZ���,������w��U\��["�����<h-	�]�;涴��}-J�E	��y�uප��^e�$��R�U�7:=�=~Csw`L�vr�Ø )W*�ս%��
�p����^��m+t�Rj�ًȫ�&�w����v�����꒢���I)�����.���aFUD^��d��-��^��(�my֏����z�Zо��.nc�����ǭՌ<�������K|�&��a�5����4�eG9�HC�+�S��^��t<\���4E<J�Q�wƧp(��ת�2�/8��J��-�o��F���{Kw4^̩�z��N���`v�N�:;�e7��W�,ѧ�#r��&��z9V�.D���B�����Zc#� �����u�����2��K];"qu%�Z�#�2B:��9�Lg���/t��	��Uw�z�=�ù���wb޸��|5��0�:�����쪲�9�V^��c|���#�ѳ�RӞ)h����>[l�h���������d!�٭Wa�TN�vÿ���vl3.PB��{ ��7Fc�f�:P�����]"6�W�h�]f� ˧Yo|�m;S��7e��O�h}�BWNX[����Ǚq�Znb=�6�{ġ\�{��+"��[�IoYJ�Ć�x��-�k��f�Mr㽕�+�@S��ͯ[���4B�&?#�'cBkI�wo=�w���+��햓�rK~�p���Dn��/C��4�{�^5d�A�����{qu�q�)���.u��X�)��q�>�bI��
��j��GY���r`�]X��'X3%�;���tb~5Q.�.�ً]�/�{1}L��v*8��C0m�m��u�ټ��=s�����$Z7��9�YI�N�FR$�"G��������暿T�1��!�*�����.$�
���;����gF���t�49;��Y����m�h���'�vm�z�ɜF`����Moq�=��h��umB�m�]�P�8(d���ڔ�0���� bq�%��{]{)�1YO��x�FhiD��6����=�
v'��V=�׊zN�}�~U���Y�N^��%g8�.ShV,���H|�s�~�5�b�4M�Dsn(��z�ު�	�,7B��]�NaQ��r	����Zf�ī6.�1�Xvfb���V.��#�K3�r�6�n�W(���2�}Ҏ4�=3�wd��*�E�=������+�%�y�l�(N�[��7-I�I ��-�����d����s�M��Im�(�UR8���f�ˍ|�_,�(05Nu7�Ե�.�%���rΎ6b�v�e��/6�5�8���m�r:wa�D��Nsp��Ε��p�~�aĕ�D �V4gX�����r��X�$u�̮��|�&�_�JO�(��No��~&l�F_1ݨ7S�<��50�Fp�d�E�8�S1sm�[<l�O��:�P�w!���9%�ysA ��C��̕~�*�9���<����x�rr�e8E�X����46?0+�Vos,�\�W���!�@���֣fi����eG�*oV����E�r ��`
/o6ܓ8���PF!wW�m>#�fʺ���.������:�]E+L��][$Y��K\��t��|5�/Rh�хҶ��i#\(�9�s%������I	T�+J��м�E���a
ƝwqT���slQ&�����<=��R��w���F�ڽ4�E���`�]t���8�y�N��V���rqw���y���'�k��>]�Sy[�U��L���U��i>�����3s�%��|+.Wf�u��C(Q�2���4C���|�d�]�I{`��(��c�3W1[�wϛD	7s%Ɇ�����\z�@�a�X���n�N��_,�������DZ4��M�Z�] X{%�[ŵ��U� ݼ5e�t�R��b�9��d��=n��D��К��n�LuS�}(��1�����;�o0L����MTϑ�Ov�>�v�.��B\�gy��s���YWK�)�k-�\\�[�i�ЌL+k��1%�C1*1����T�*�c+S�a��$�B���0�V!v��XL[0�ZbCG�#DH�K2��)�īm�Q- �#J%Tj�d-��C��X�5�ĥ����V�	��0��b�a����ADk	x����vEhZi�D�Ss	b�N�Ø��\��qW�*w��b���>։l�Be\yz��6��^����I���y�t��M�_Μ-���DZ����xQ���۔�ST�v�f0��-ͪ�c�lp��h��v��y�\k=��8��Rl}p�r�Ot�^N��h��>]��
�º:�J!��ش/-�)<��!כ��x`V=I�����\2���c����y���](���m);:pT\���[*x�����ԉ������~�.���44��� ;p�
�%ɢxd���XpC�!+���~*�m��t�Ⱦ�-ͪA��\^�k�z���u���gm��	dN�uٻO�I8;��i:C��:v��i��E-X7��ZcsP��;��gw��N4[ނ�Y�Y}�%��UI�R�`����Ce<�\���+^v�g!�7d�n�;�H��{=Y;8>��=h�)7��>��O����X���u��fk��ׅz�AA����joؐN����<��b���ت	��`��Px�k)� I�:aa���{���^���Iഒ�y��;8���dJa�{#�e��G+�5\�/��^��t�4�u\�@D��wu�R�v��pΜ�������M��]�l^˫.kHK:�ӧ�L��v���R2�gY��M������p�'s�c&�~	Ԕ�
�S)H�)Q�Xk�A
{�8�/���>��k���U���}g!
n�ϞX' IG�|�(�h�-,�d��=��߮�(�}@v�� ����/�xi�e%��\\�/;a�s(�7"��'M�u.��L�gkK�Z1��z�iͅb �k5.F��2��F��F8b@Y�s��]zBq��Y��35y�U�RtB�	a�{x�Wq��Y��aۧ��Ú���))���pm�[���i��w��Ǔ�i��u�&�*zB��nn�[��>�x����1қ^OU�o*Y!��!{�
�4�gDiB�3��B㼩ڻ���)eq��9�A�IQ�Z�@�Q���$�9�%x�۞y���.=$S�6=�+݂�#��0u�s\�]�u�p�����tA�	��y����nK�\�\s��&|=o�0�^c��Di{"Na�g6��;�T�4�v�y)�8��5ޚ[�oj�[��d�u��+7�l�tqqj˖�0���y_k);̳]WM�y*\{�%�wr���N����Q��uy����;v��/e���m/z�v���N�]2�j�t���RUp�x�V'������P�o�=G�G�Ŷ�bg�
:[�"�}B�eX�zy
E��
�OLwf��ij9ĩٺ�b��\��B%�h��&R
�Nv��4�}���+�ߗ��6�1'��bމ�F(Wh�a���G�LY����DG[�M�,wcy%�Iz����_'�)s�y� ����wf)��@9P�m�;QK��P�yGC���yJQ��a�sӹ�)��f�YνMu�R`�ы]AGyu�x�y%�>�<����6F�S���+�-�mqOßS�}+}W���[e���W֓:�=����ol���{����\{9�|��c{+q�+�k�ڀ�/.0�4����w�O��c��]��(�5�h��������o�.)�k�e�� �<���"���2�!��
@�
y����}��g+�g�X��~��A��Lkۇ�/�����킭���O��^�>3��W�ս�L�#���⮤�Es�ݝ��d����:���EZ��]�o�os���5	��\�@��0�|�c���,Wi�s������W4���U�Iw6��J�f�cY�z-�kƹ*疕�4�A����b�����sE���d�oD��0�!�s�e.�YK�� X���j��Α��N��3Ǚ�Q����U��X����EUU?}%A+(s�(*�x������Q�X��"��$)*`�7?!�?����0gF<�N��*���D�*��,?��
ĵ�X�F�����Y�MqO,h:�k���E���7J�POIM�1�sw֜3�n} �xqt�|�S��ؕ8��x�s o��4�ާ�*�w�����A.Tt�]����5PO�^󙞻r�g�;A>#�T�^ %�i���:'�H����������z��B�װy�J����&_P<��*=]�d��q���
�߱�����f��f���)�Z�JwW �w��G)��Σ߀�
W���
�*�L�5E뾫S}�eq!. �	d�B�P�ZI��B�/���4�}w1�٠},hx(*�kpG�a���k}A��d���d]�f���Qo$�}�Q�?3����p��k��AT��T	Q7��6a��^������jl6ᾕu	@(8���N�f]��Ip7�u?!���eu������{Gq�ATk�@�2���d���p2�n9T��҆� �#�D6 �"\eG�AT����([� �R]��UC�r1.� 4.��p?�E 0��B0}�թ7P'���PHE�(2lhܯ��c�}/ޠuq�(O�wE�t�?x�J;�91˪���Uͨwq;��8'PIo#�_��f׿h`g�[�`|G��Wx 9��v�>�@�7���ӵ��D����nJ�8�V߇�PAT����|ދ'��@~�xd�� �	E�.wɩ�y��g�C�?f�6���M����� �J'���� �J��s����4�/�03 �.z�^�*�����wˈ*�v���gڸ�Ⓕ)�cȇ�)Bs����Cq]z����(�.�ݢ��EPO�@�p	�y>����ǯb��'Z�7$\��^\�8�����5�W�ks 6�^K�D�5������"�(Hb@�(�