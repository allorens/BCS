BZh91AY&SYz33��;_�py����߰����  a�N��          (  w     �         �x��m�eb*�B5`p�
 ف�/>@(H �i 5M��/�tӡk�.�ޚ�4�Ό�������h 3�s�BT�u�w�y�*��eJ ( �Pi�K��%/{�m�W�5Zn  y�`�4kI611׮�(��m�U%g��];��4 pi7*��-��� l�U�E��{dQ�t�� GG  ��s���$���������y�IB��=����0�c&��Ppa�ݎ��N�W�W��z��;�n�vd-����0��{ `�*Q{e��z�k���!+���aǶ���T�Ҷh���ӲI*֔k����<z^ڢl��Y:� ����]g`��T���[{�ӷ;YB�s�� /(��Q1�D����I��.�#v��l�gG�8    $   �(R�P�  ��T")� @  ��O��J���40A�L� dh@�?%%R��ѓF  &CLFOȕD�P        	4�T�4�`	���� ��1%4�&@���1��=M ��*Pa2hh���h��v�điJI)+Px��qqD����h��7�ׇX(��ꨂ	�@EG`������(J�*(�8"���G�Tzja*�h�"d"�d!!! �XM��V���MI		�����C ����
{"�� ���C�̼�'O��]�ܹ�w��5*vvK��4aI�Ķ�Ai1!8+��*G�|�4`xL'���h���p�eD��"]eN�㼩�>��{>��TJ2��N��$�f����u�Գegd�&��Tu&�N���v�ʖ"`�1)0�Æ�M	Dd8��}����$�D�H�#���u,��ǏTه��K8l����6P��
:q�J䉜��%�Q�c|�����x��'٬jo$��sU>A'Ɂ!�E}B%�9�Tk���K̩�ӕ(z�LƢ#��F�|)>W�h�$f4`7���?"I0��2���n���w�0�r��w�*�),�t�ؔ6ԣf&����,�i&�/��]D�&�/>�d��$0ԇ��42Q�4wMNdN�<4Q��'D����2��.&̅�6k�0�9Sd:�����Nn}h ��\$(���kUb;�Dϰ�0�L0GmN"fڝ�l�:��Ć�H�ڛ6Y�셍�"`�S�Y�jP�;�Gn}�E��p�E��D؏;Qb#"^�%MNA��0sUgM��Q�7#۩G�8�J����`��*&���O�GuSf�DG�Q:'9eY������S(ؒM�ڑ�D�R��D�f���a"Q�U/s�N����,N��"ax���>�P�֪'.'EJKR��+	Af���N�]0wҸ'��6M�M��ja�|�"hseY�tu��x$�V���m)����e�ɛ�r%4R�e؈�D����p�F��	�bWnCN�K4QGI֤HN5>A��5�R���yʈ���'^���ĤN�&���-�6ԶM��"&�I0�o��J����R#mK0E����ԊH�~�L(�d�����*i"hե&�;�T�f�M���RP�jCd��	�jQ���d���:�&nD�u(Fr�	�ʈ�mNdÆ�e:$M��LySkQ�SB,�(�Z�t��D�e�4?"Q�X�|�܂d�K8=�:";�Y��j"&�����G频�j"#�Ĳ��DF��"aē��6�"5>G���D�N���AyS��fT�,Ѭ�P��DD��6`�h��K(��%":�LUp�V�˪D�t��!IPEeP�eK%�\��ag��I�&ԮcU+�;�PD~M�g^JL2pN��B�Nț7ܔ�a�C��Jؔ4����~�%:��o%"X�-�0D��gJ�~�%5)4"q�I{"2k�K::쯐~̔�d٧R��#Ș&�>�(A5D~�,�H�70��[4";�y>����F�j'D�r�:jD;�H����&7*����ܤKfSS���2�j����MMJD��{)o���X�@D���h��8��艎�#���J��>F����R'�ؕ��&�R&v��>�Ǻ����(,a҇q6X��DnlMa/$�2|��Q���hM����JL6[��v�`�w):`�UF��Uʪ�h�+퉽${ڈ��L���Vt��ʈ�4#qj�ϨnB�����6=j��6Q��Q�Ye:��N"<��J�H2|����D�U�ao���N	��U��4%���l��"�V&�Tޥt�@�� �r��QL��IMA�V�ha��TA$4��lJj�Rj�_Q�&���P�%9)6hMcUF�,�hG�BlM�+y�uj�p��p��ٲ������"c�]��V�%�[+���=��7ȉ�p�?D��َJ颾M�L�e�X��n��"A�Dϑ!�R�({gJ�{) ���h�mJDG�+��?	� �F�%	BRʡ��#ɂa�UbYΓ�8h~w))�G�c0M	��K67$��I�e�M76%)et�2�D��0L{U��o��;S��8A�H���!õ�L�XFB�?Q;R�N�&oR��iepM܇�3Bt�a���$]JDL�ִV$؈�UF%��,؜,{��ᣆ��T�>�	��)ܤ�!{JL6;�|����
8��L�WD�C�+�3�R':'m)��K:k��*�q8B���Y�6CI
+���%6�����#wQ0N-J0�$j`�w�HtN���f�&͚�I�N�����B�Eȯ������Į ��_�Ș�RieY��l�2��Pٴ�A.��S%��h�$�6G���#r��)eh�d�Y>�r�A�pM�u>~Z��$�J'*RWé�(�*�E�Q��M	[$�>4A�M�����Uf2��)�;���$�	��I��(/�Ht�g��d�ML|j�#uU���]��"&��aF?DD�Du*�DG�(s�b"<j��%ԫľK(�I������C�&:�d!bh~уQǱ4?����o���*�D�r�3S�n#q���ߢpur�E�:j��D��R#rM�~L,ӹI�oe&���åT�gelN7),Kw(ʕ��)[+���6&��+� �g�ʇh��oe'D������d�)��J��3M	E�W�'!tFN�6P�ӃQ;B:�C�50G��� ��Ȉ�D���Dn'u�mj�O�h�Hs��|��	pG%ޑ��}����O�T~y+BhK4�f���&�8�ķR����?Cg>��6��4?"aX&�g6ɜ'J8f�'�3eցΥ6^�>�iD��p�aZ)4h��h���O�kE	���	¶'4[r#��^�p��	ҵ��D�Ԫ8n�V�KDt&wu:l�N������5mJ/�;�jI�?O���iD)�4\i�2���1�I���?������g� �]ޛ�K���?��zA�L�9O�w	�D�����{�[
8*�]S5Ŝ9q�MM��8m����O:w�n���c��%�������W���a��Es	½�*��t�~$��?n2}��@T�N�x[��V捖q˻�l�{�E�l�3d���V緾�j��o?Ͻ��R�G��N|lⴣ����:~��W��9i�{��B3is��C6`�uڱ��9-���P���??��l�}F���pU�s��E�@;�/M*���~�γ:�g�(���øNg�"���{�x�ӄnZGB�5e��ßM0�7����fE��s�+?݂+^���4�?��o4�0�݂��,����;1U9�˦�{��������ҙ���7��_V����u��s����*?Q��^�Y�7�/#���'z{1�b�~��0�]�L�p�	��e=��>�f��rUNM�t�FN~�[{�[���K�
!$jm�2�8*U�"�o��}>�Z$�߻�sO���;�YKY;9ø����_8��}�}_��]���l�4z�D�XK&�������qe]9������7Qh�w�xK'�z9~���rc���҄����7}�d�٦�_>��J���Hp&v��p��o��+���ݍ��k�\�f�a��f<ǤZl�cܭh�XWn�v���F��?:}��J*"���C��a�f0���u;�\�6���m���t~(�i��TY��=�'����T9�LW�͐2ܙ{��\'v���@0P�~s�>0�rt�w�T��ψ����=���f����y�ĉ2c�uR~�Jє�]R����ʸt[T6;��2�dˁ�>xd�����Bx���a%r9���{��4�ެ��y�6�'O�Y�~㞬C�lZQX�3
*c@l����J�}�`A<�g���ӻ�����5q����m��_{�'iV��V=Ɣ��ڏbs��}n����^;K��X��\%��;�W����x�dj�pb���t�6����@�I 8ke�a3NC�v�$1�.�O#��4_g�Y��p��e��p���6�߮���U
�Y]��Ge�)�8zi��[x�$ΒW!H�:܈"$.6d�%�^�t�)�b&4@�u��=}-2�x�߷���9�,���u��c�����-����yb"-��hk�y�^�/������4ýJ���&q��#�q��T�_>=�a����u����������@i����Z$���1�2��t�i7��}M����lqvv!��#����*1�ͳܶV�/[����.�o&oy�╾:���P��r��%^��O�l:�ssn�����ŤR=cZ���)*�H����/��<�a^��������2u���疼u�8��iz��	^LZ�������fa��KA|���z�8I����ϟhY����榟M��q�◛W�-�[˔{}�����C��4�V�#N�[B�il\�;pi*�����)�*�=m(��$��ouk1�H��^~�o��d�?:�쭠��G�$�n8t�{a��m�v���\s#6k�k�zi=sB�7����n�'Z�	��ۯ��O�8�����7��#�!�zf�L�[��`��<�r��XFi�6]~տvJ|���>�M��8J}����O�oP��5�iV���p���Xk9v�{��g^�������^ˉݾ|��ш��֠��N�a�fN|�¯>9��$@J�_����f��_�d%L����+���{�W7�]2Z���8t���ޕ�H�;�}�ѓ�Ѽ�ZB��C�2B���>9��-����Y2݃��YY��Ը1hC}�2�@Wۋ9�=�),4�d_Z�{���{T�C2«|s�������Ϧ����'��}7�|�b g�(��g0���Nz^-���᏾�I��7��7����c�θ��GY��W��>\��f�����q�{|%oݐ\*	>3y�ݜ~<��>�S����>+q��ן���~x�g&��%��ߏ���?g�����/qߜ�S	)�(U�Y���ɣ�}w{Q�K�]7����㤨�a�}j$��dǝ����c�jUJ���ٯ��tѦ����t�˖���oW�٭�(M�����og�o�P�ݢӇdg7v�	Fwh���C2��J���s����@e��%\��n1�����rr��@p���qΔ�&�wn�~ �Ra(���M翽��S?�ۅ����(��
,�L�����g��I�ȞҶy�70iۍ�#�Úk,���yr=��[�]kdɛl����v��$�NͺnA�M����\r"ɵ�bT�wt����}�X��\�=[�b�{��#k41���w��G�a̞��'#��i��5!�zWN���J8Y��(���Վ��v)�<O)M%��l~�\��r3_���ߖ5����L�^��=a`���n_\>>�������G��@0}�2��W�n�xa/=�1=�Vh'�PP�'��p��&��T_\%W�]����}̼�y��������#��{=�;�M.�&�&4����$⧹���!+�--�iQ�o�d	3;3f�d��zz�a���Q���K�)�[�/���d�>w�_���+�r"���3��y�*fY�،�*C�qL�ݏ�����l�	nY�����|�y�#"�_�/�^J�y�ۜ,����y)�o����E���8KA��p���N:0~Y)�߯\�����a�x,�݇�'�<O��sj$�ca���E�;��o�U.홷�BH�ݫ�i8t�<,�.F�]�v��l�d��Y�F��]|q�ܙ�w�;����gL�t-���1n9��k86����]���ߣ[U��dxFn�ː��jF��u�􇴟��=�Lw&Mَvd�{x�.CѺ��{�n5��kgu�"��x��=;�x�*�����o����zI�"�P�G�o;/;����g�+<�������׉ꊸ4��ƌ��_��pË�Rv[��uI����C�p>��vB����$+�=El�1<x��-�#�yy6sk$��!��?L8/������t�G2�]�˲�����lC�Ϧ���HBSB۰�U!��`�P���`3X앎0����dRh܂L"$Hp�I,FKq&QNBeԣ�]FڴŁ�R-�]d�m�����:�}Y��Kw��N"���n�H�[�@�#�۠���#	�$nD�2'��w��c^�N�`��L� O�:	i���v�ۙJ�$�)�H}��0~}0�*U �`D�!#��ݥ�nȉJ�ԁl��K2��c�~��'#7�<��)J^ܽ`�)=N�R�}����A(0�M��L��!:�櫜Q��Z�Ű�����8�*/�������D�)����0��<}f'�����&��	��}'�iH��A�MƾL��oD4�>m�[|�4�l���X*��%:�,��4��6��V(�S��R���U�q3��&��տF��z!�
z�U�WJL�����1)l��]tt������G�`�5�k����$@ì�T�$RO� �����I��{'���hI%c$�*�%�(c,͈���Ux��EX�yL�S2`\���:���:N�}���#3���\�U��sC'T�-:����I�2����$$ʌ��Ƶb��[��Yg9�N�GYڽ�`q6T���E�Dy>��.3�9���s��C��
�G)����>e�j �`����������y��o�f���kgqU�M*É9��6��W*ʚ��p$yR(?z��	�>' ��EH%�\���Gu�1�:���V����͛�ܱyh���*1�nUg8b������^���J?vY���ULeM���fU{���[ݬ*��J��r��CH��W���*$@F/�!l�a�D3R�nZ	0�P���Xq��Fߐ� �!\i,�Fb�`ͣ5o����T E�����Ne�Q�@�\�>K˯F�Kb͡���Sؑ�q+&���g��?Z��痾P��֠v��s1��� q�s5�����C�nXxu}I�O3^�q��|��&0�&w��Yg3}�:b��λ�t��k<}�ܽ�^!�;A`v��!�:�8������n$�	̤��^��u �p��V2������o9�6���M0P
li�j�0Q1?7w�hC�]S,S��u���-�p�DP�15��sr��Z�ZֵmkZ��ª��������Uڮ�W��U^�J��9�qU괪��UV�E[^��Wj��Umb��"��S�`�ā�'��}���>���ġUŵ�U�եUmb��"���.1x��U��W�{���v��U⫵W�UV*��ok�x��[]kZ־ֵ-kZְ�.0UYE���UWU^��Wj�t��X�����kJ��1U^��{ޫkJ��]*��t��U�*��Ҫ��*�v��iP�Sﾐ �W��k�����V*��t��Uڮ�W�UqUUU�{;��WUUQUU�*�Ux�*�h������U�}���ā�ğF,�R�,4b"$�k5��EE��B����|=���#�g�8�N&�p����N��6K,D�0N�&t����6&�d�ɳEA�%	�B"pN��	���%	�4a�`�lN�bYgD�Ht�0�(J(MA���:"X�bl�"A(��a[&YDd˧N�:�:P���DL�h�"A͉�8pJ�"a�""%���t�0L8%�f�L!bp��t�B$bX�e�0��p���u�;%Z:uꪴ�t�r���O���i��2���\�[���jJ!i4ո=�!�^�G���hҒ$B�u����Dp&RQF�MH_Ĺ!(� D�(�Iz��$�kOe�ܔ�Qج�P�����sVS]XR����mtSGi�n���޽���.���#�s)]�C[�vN���a�t� P���ε LݍCe�bKR�����ϥ���}}W�L��.�l-���[m,ǨRi�fu�.�Ƽue�ҹ����ʷ̫�sA�ݻs��Yry=��Y���v����j��C)pĒd���eԝl�gЃ`'�X-y��J�ć�4��:ʬe�fJm���5f�c[u�vϝV4���_��$V�p��V����3m�5�հ�DL�iR#B�nf 6��si����m�z�U�H�P.��a6���-�]��2ᅱ��%��Vc/-%D��~@�I:Ā��&,"Ң���B�0��dvl[m���!P�u�j����-+�D[l��ˁ2��s�+���e�%)n�um@m3m a))F��3�8��F���XN:��[L:�ՆXLf�gk���[�3u�fXQE��t��Mh��e k�z���Fϵ�Gż�96�Kn��i���N�̩�[AZ�+XFh�C1#���cYq�xh*�,
����5�s,�k��2�7.��w�=	�u��8	���``�bfB�e|ZHF͛�/�Z���K,ǜF[A@�N8�n
����)�?3f�$��d��V^5D��p6���n�F*I\&�R��m������sj�I��ԍ��4��@IvŦ1�1;��x[���5��)*�R�KDfm���P��wF���4SX��(�-(�[Lɱ]]`Zjz���ܹ��W	,��	�qu����K����z��Y�e��LG.�!��n��R:bc��/؎#��[pG\'�)������gGm���r�Ŕ�]1Sƍ��������^�x�
޸�ҥLg6m�,.��aU%5�K��&HKtt�Mi��1Z!BYa�
��)D,E�� �9m�>�"�-k�Qk21
IB�0��"A$��&22���4 �����[h:�q�I���њW�Rh!�Y�b\�����.in��v���BH��}�����}��>��{���뻻��}��W��{��������^���{�wwwy�
�4�Ϟq��>u�6�&�ц0N��ݽ�5�uTn�7�e�t�1t�2�j]}��}w���8�gF�n�Ul�I��1�
�-ivǕ0���m��M�v��dչ�o�[�j��Ҫ[5��P�2�M����k6lֺ.���������ܱSc�<�u��\�w0�m)���*т��L��hI�X`�c2�']�hRGBW`�eF�2���sKq��T�ۮ�:ö��*k�����	���$CMw��ƛ�7��?��F7��;i1.�	�t3�p�/�+�)3������Z.k�8?���̶�._�ÒtwW�xu�mj���gT�bS5�)�j���q�M0�����K]n����|�6f�\y�����[-�]ܨ}��2BF���N�nvn5�̮�Ð`��_a����֫鷺��+T��?C��ۏ8�Ş:'DM	�8`�'J��ffX:��'�Ϧ��߾��֩�2��p�uљ��<Ð|��'c�um��>�0�}>:�8aɲt�����|(0��cOH�E|�H�nf�fC���z(d;��Ӄ�a��w)�,�8ҴóN�!J:YfxL,�4&�0ᇧG^�kU!�<nl�FDÿS������#{������p�N,���������}mD�>�Stzl6w)]�t�Sn	�q3˖�W�zz�!�t��������063g
�!ٷ�3��1��:|g:�����&�{��n�{��}��U�h�f������l<�8���L,�4&�0�t��T$ IR:7P�v�ݻ�M�F���8����AB)2�H�A#)!��_8��\8p�����Y�X�m��]V鶞��4�|�X;^0f�M��،Is��֜�����m"톽e�
g����5yU�H�aN�g�>�N<&ab&tN���p����A�:j1%,U�P���uT�!��V��n2%�pޖ�.6�-���$$2�i�B���MH�Ed�����He�*z$&s��*�$a�=�B�'*�����=�_�-��/�1�M_��Ԉ҂� p��������C�(d=�<8`�Dm�&*����&���\��8ڬ�Xts�]F�|�>I�>C�OO��y�	������C��Yd�<������ �9�+bI	J�!Y�ތ�n���ò�
S�(h�ӇL0�&pN�Fp���6ũ*Tĸ�2��a�˗A}�C�>CÇs�p��ۛa}T�����xp�N����=,�G�A���ў{�QUq+1��z>� ��b�a�aG�"=\n��S��@��=^>��d��==4v%��UG�N�4:�hN�`�&	���&��i�[}YL%UH�����s�4����.��r$yT�����.J�,'iQ@)><4�Mʶ����rt|`SaO����L������/�i�	DǥV�6D�Ѣ|�'����}YK:�vNi����-v���`oC�鲊�*p�̙��W��S�����Z<����,��i��u��8���Yu�a�q�Ѯ����0;QZas�M��;�t����s-2�pW
�fV��g���OD4O ����4a؇�=p�N����|�j�()�.f_.�+a(�y0-�Jq"�I+6�x��"+�O��Q��h�{a[C���D��&pM��Fp�:w��L��9+����`-�"Od��Y{&��_A�m٧u�X�N�k��JS80��i�e��[�g�3!k�|f��	�GQ�A̟0n�_�n+A<��)4REDi=)�c	��<�9t�q	��gx�!�:�6���7e��(�F�_�o;�'w��L5�p�4S������ [�{���e��b�F&Cg�����P�=J!�N�w��IM�M�O��R��6��3�-π�Wk��r�gX��l��'�7�̴ۜ�d0&���ѿT��(酈�""af�؉�a�q���u��o��q��u��iV9�㘗�s�SbS��=K���Զ\:���C%��0��i·BÓ;<����!H�S��v1>ð!N���Z�-����%��>..۾vx{�L�=ri'�}��E[�"R2I�̙1L�IO4֨��5�2�&V���/��i�<Y�j�a�a^0M"a���N�m�ؖ�7ry�����������'�\�c̯�///�/i����8�[�:�N����y8�y}y}O8�6��_������k�u�Ɨ�^����O'�q�p�L0�&R�1�<��/ɷ�c���/μǓ��~'�����i�x�&R&S)h��D�h�T�\��^ַ�_�ɗ���/by~v痷�b߮O��O��?0��������,�G���~O8�y~i~O<�#έ���Ǳ'S����q<���q�J�����=�%�������؞^�_�|ǜ^[_�������Z��W�>)K���v�	�D~ן��^��~m��ۼ�������eMb����tL};�>NK(x�-
悃�HV=�g��"�!�4�f�t���j���8�8��)S��� >�.z���¸����/����|1T6vv�N����>h���������߆�^��}��v��]�پ�D,>^����������B{����]�ݹ���'��{�����ߟ}=^���{.������t�o<�ϝyמy�_2�/:��2������9<��mѻ�
�DN��I���4C��tad�J��xq��֒�����	�0#�G�Dz����$��29OͰ!��~�-0I��v2�!FO�h�"uB0d>a9���������G9˜����*,�8(!�(���!֥�!���e��wJ����F���DJSt� ��!�K	�N���`0I;"5tieFj���:�t�\������k�~�\r��4{�A'#$;�$>A!���ʍ�V.[e�]��#���vR�R�C)T}O0«�J.����?:�8�<�̼�<ˮ6��ȧ��}UV""�07)�:���ܴ����$���,�E �W�CIJ|�֪~�X�%��B&�a�l`��",�ҫқB�B��٫DGlV�" tx*�2RdDDbNT��"�%~M1C/R�ӕt�!èS�����o�yU�&<����Il~����b��$DH,���h�t0(������"��~0�<�	���'Q�d(��8�'���Sc��4��kY�NJy'�L""C��}�	u��JJ=Hp�ԥu��^X���?L,���4l��~��#+#�x�@e�dq�4�K{���XI��k���02c��% ݆Y��A%$Y��d��2� �#J�m�H��Q#_RH$�A_�xz���,ߠ#L7Fߤ$�aܿi3�0�:.N$z�מ��{Շeg^���8�d�-�cnF/�@��)�3bp@�FH��:xRh����I���ɩ��8&p�R@�<;��D~��Q%Wv΢�}%�����p2�%4�"O�a��P,ȅM�*�eaL?.]�ҡ��m������$E�aJ;Hy�;�	�2OFN�C�s�Y%�#��]�bQ���#�a(v2t��"r�I� ���'�
M���\�P�̷R�(�����Ls���	��&a`~����r���> ��Nby�������O�N�)O�R��+��~|����?8۽���/<�/2뭺��}�I$���~!1KjUv�b�b�S�%/J!���h���a��Ld��Q`�
 "'�N��wk���u82y#	�i��*DN��C!�C�'T�$�%���MN�܇grRQ�
���KL60��+#�;�U�A5��'#	Г`����h��<�癅�~M����#%��t��,�ON����t�èo�0����i�d��80(�d����Y:���: �%� �`pC�~���0�b"{��2I�PI$��aK<�T�2pDd�	%)Y(J]���I�2���y���u��y�^y�^e�[u�ʥE�w�Uه�UQ�r�=�h~�h�U~��c���|������H�AAC��fA+	���-]>E� $d�l3������a�D]	T�l��߾��N'�!d谩82`�����qM�cKpM��G�3'�Y(6MO��!؈��P�~À��N��)�{mOVl=�`:QJ;;�&FA	���Hh����	��#ِ�:e,�	D	�%�h��O��#p�!Bu�<L<l��"(�tl3	�<����r0�`�����ȟ��ܐ�آS���a�"���p��,���<�������6믖��/<�/2뭺�+�t�j��#��� ���gԵ�Xu���R$P
��@�d<�pz��2Ldc$�"f�)~�-�2��Qni7�D�sLwt�Bv��P:,#)d�I�A�`"$d;�4܅%CA�@`�~��FI؅d��2� =:�	��Y=['C!���A=�vN��҃�#I������q�����������XI)<�*fH��<ԇP`{�#�C�I���������A��M�� ��LMM`��F�!Ȑ�*��R�$��iO�%#m�6��8��ۭ���a�y�]<;�hdm7���sW6���մ7j�C��CY(��U��Co8U}�_��C �p�Lh�Q�Kā	�"!��
��s��I ������j� �����Hi�VZ׶�.�n4�r7���:i9^fNB1�4c��`�Hk�c4�?���?��P�����&�2�,�O�}�����
���웥j��uL�"22Q�>�� h!��d)�!���ۻ���<<�x��ұb�Z�8"2(|2@�Z��C�u�7K�%�V���4CRAIM���!�J���?t0R�@�LC�,;�!�`tO�48�#?�	���a�	�����D���4�c � ���hq0�D` !k����>K�Sn�[�DP!>� `0�Q��
Hw����6C� �)�|���6����:�n�����y��e�[u*GҤ"j�n5��UT`
=Ĥ0�dHä�d�A����!؄�!O�"I�.�1%]��R�En�e*�z`�E��0��Ʃ��-�)��82L�P�(�A������/F�ä��S�\Rmt�y��j��E�L\�4%����b���Z~V�6�S5��Q��8L�mC�!�<���܆%S��벹��񣾒<����0Ȇ��aD`T�aLd<����Pd	;�\8����*# �E�M(,�,w�<�[�b�F�Z���YoSKUw�F��m�?8덴�מ[�0|p��ӣ��Q��XW֬�iw�5������dJ~��]�DS�0ً>X����a�V��`��6�a�ã)�A�m�q�v3'�Oy�o���gT�J4`mT�_�\}=9�b&�D�,ƘT��0�"JL���5�ry�O�<O�)��\ad�|��w�@����=�B�.0���Ф�ZM�d@�M����9'E�á�3�a���JOD��y������bv��4���<�����1��T�N�ɊAʌ�6�"4�]1���2m�κ���N�~yo<��2뭺��IԈb�_�UTByxD��hl=I�ٲ�.j��ޥ��Էq*E�\z� v'YJ!�w��r�S4��gߠ���-܃(���{A'���89�5X~ŽA�G?|�L�.6ZQ��3	S�}�NA6~"y�.�D"y��Ն���Fߟ�׆i�H�.�Fش����-�CLߡ�:�3���`�d�|�x�R鶛a)j�O���ߌ�q�F+��"O�%�d�G����1#����e��a�־~_�i�<W����4�)�%a6N�ŕd�<�O2�4���2ǙZ��x�����^g)���c��I~G�n���u#��m��y}y}O8�6��8�8��H�K��ˌ�̼�����αi�W������z���2�i~yW�yט�q�b]_�.y/���
_���.�mUt��"z�z�����^��0�'����|?���Z}X�U��_˥��~i��ͣ����<�:�y~e�I��a<%}��V�Rx�M��<��N6�<���>�����yz�cɧ�����&$��?<ǝ[�t���E�Q?��_�(�>0G��(����a9���|�l�W��Dra�4��]7c4��xK{5����r��Aj)eN5�en���֜�Sp]Ye��'m��_���2=_�^�������\ܯ�G��YE{{�����~�xYstԆ�r����@BC$���k�B��jkl��.ͧnnh��͝[J[`R/i��%($]����8߫�83���JL����nU�s��O,cC�zȘ�r}Yϖ�J>�f,G�dxIeu���������#�v���ő2���Zs'������n�yܾ[��Ha�&�-7f(���Oq�������W|��[�n��$j�q1g�s}e?O�rQ��W���0s���׎��B�m��2)*�טw�����Z�Hx��_�-s�l���|�P�5�R�X�2�3o+umu���I�'$9i��ŕ|�l�i:$�]��="�A���nH�QG��UI�Z�ƣ���	�+$BZh���,2ۏ�1��龽5thK��5����P��+���R�6�8��T&�/߱���M���o�C�@�~s������ww�>=�{������w�
��������U[�fff{���0L:pA<x�Ǎ8lD���
�	�C�'$SL)	�(Y5�ƚ�6�3��m��-�y�3FЉ6�ḱ��}qr�4��\��7�d-6ijv6�������CF``�6�D�Aٴ.u�]����0`/�`�l2��"Wb��41�+	F�*b���\뗍�<�PE)�j�X��\JMA�%+�n3M��\��y���&�<$YHL_)�����fU��M"Vmn��Y`�ί��a�Ԛ�Om�6"dH�$�AKې¸���j��T]78���'�t���Ǎdi�)�=�u��`���� H~e�E|����Ŧ?R~r�C�l�j���cS��'���Ƚvw
�ge
y'�FВ�8BXS�NK��Ɇ��Ky8�i�}X{\�Vi�-����X]=,:;Fvvic��=��ԟ�&(\��N�%���q;^d7�w��R��ϟ��j��������/��/�p��,�n:����N�y��4ˮ����"r؆���d���UD?p}:;�׿/��r��]�i/->�|���&ܩ��IX|�&��|�S�.�]��k.c���V��V�oε�a7[=�g?�RY�H3du�g����I+�}�1p��[DkT��b/1i���id����zpL:`��j�Y�\S]���7��D�[�1�7Nq�̺��8덴�����<�.���(��f�*���.ꪢl<��8S��������F���b�8�~��M��������ϙ��n�Z�,J�Y{�������H+v숁H	�K(a8���l���b�~�j�q�����0�fd�ٳ�U�I����o��r�?O�����}�R~��i���,����X�$ھ1��2�O������o��q�u��q��:���y��e�[zp�$CY!���M��*�!����9H�<�3�;a������=�Gd��~�v�h�J��TO�1@m�p�!�8Q�{�U�_��)Ӿ�0Ľ6r5�)'X��2��aI_��{5\�_S�[��[��3$h�o���bO=�"�OCl6l��pA���Am�tvN{�R����Q�vdX�I�X}�J��>�R�c�>>q��^~q�iӯ<��a�u��s|����Y�I	�ȓPI�aI���&����dn�J��b�S?�}��R�5�� �!l��Ѐ�%�/��YIY��޵�!�t�\�_�Q�$����I$�@Zv�Q���d���2�9ل7�����]w_Tp�8y�9w���V:$���nL$����e���>���9[1H�-_R�1�ORm��fo��]:�[]�H>���j�奻��'?I�kV�b�O�LF'a��κ�n���yR�|�:��n�~Y���ļ^+r�~�uά�a��?W�E4��8`vuD;�����W���L�j��ٍekO�y��opN���i����Ӛ��>�w������8���N�u�o<��4뭻O�X^�UTB��q�d�á'&}Îu�6�k(��a�ÿ﵉�b�0SC�O����	��	�Yl�6|b�)��]S��E��p�g/�n^����'pS�.���r`���Zhw����6�q�/�<D�����i�xs���L;>���%�Ѻ���q�ڧ���ܸ���:�tk&��=<ƪ'�{kƾf��9U��W��y0f���i�>i矟�u��t��y�^1G��0~$��cAQ.A�	&H��J����~�n$�O6����9��:2�%?z�
�2�hr��w�r�q���5�0��s�I�2�(� ��
F�I� o�ĸdE��ġ�2#d翾��F��ӷ����޹w�)�8~>[��l3Ĥ�gW��S}�3��if?"Ҳ�j1��ޮᬛ3Q��Kn�_�|��b���/�L�y�y��\m�N��<�/0ˮ���ʳK���+:a�1$z�8���1���z��y�O]i�����xu�|��뽞�VN��1'\~�uST�,�o���|�'1����U��k�%DT!�SU�K���E�~Z�Cy�JR��~:�<�P�(s���Xu��|�8d�8����m�_��v-��Մ0Ԅb��n�'������Z>m���yt�S�e�|jT~�Wo�ܽ>��?m���r�a�!�P�1��Y��6��<��6ӧ]G���A�1��	��W���a�x�1��	��m����oVɂ 5�6��ɕF�0��9��AaKH���XH��Xl���2H@ss���+u�U����QS5|����9Uzkr}�Y;3�]�r���r<%7|��8o�rZޫe�'�~7�/�Wr��`�[��\�u/m�n/�X8ZS���V6��Q����&��9��"hw��U�ӓa�ԓ��d�Gۧiš��ۆZq�CWnR�/�r|P�;�({up��}���oϟ>C�qLԬ�LJ`������<Կ�5TMA��?�qY	E�e�f���2�"�=Qt�y��wM��󬶏�~q��u��!�Ǎ�4lD�%���UBI�ϭu��UTC�<�ч!�������ك���Z\����]b�r��ܹN4f��Fv�.�b��qi�h�eW$0�|�T��յ��6����k��i��9M��#�O��Sd���i��kk(-�{#+�1M1ګR���3N��-�ǚ�Ͳ�2����yŰt[��؞G�뒽]m�}I�5���_ɖ�&\q�:�<��m����ט����u����2�O>}���nI�W旗��+�+���<�Z��/3��O1�������^���y(J�u0�x��&+	��5�
�Zi<��������y�<�O<�>_���a�X��<�/��^c�=���g����8��D���o1����^Z&Z�k�F���<�����i䞓�]����<�i�O-��O1��+���T���??/(���4�������q�'�^������y8�un<�'�������_�[�K�8����[�|ŧ���\�����<�>{�zO/��u�1#/���������k~.���KO�ݙ�3�ߦ����n0�8~xP5��VP%C�����U�7��~ȃ#��5vE���r'SE�w4��0O��K��  `l���(4���}3%��½��|����[��$��O̎��7>��}��U������*�܆f�nqT�[��<�-��W�.�7q�,,b���c2QH��HU5�g�׻����7�~���V�3333�ǕU�fffg�yU[�fff{ފ���333�myǝy�]m�N��<�/0����龑UTCa�ǜU��:�?�aLQr`hd�P6	���V�Ԧ�auP�����w��K�p�8b������w�?x+����V��,�8�L��~I(�1�3�k��'�d�'fA0�����?J`�S����-�6���ܭ�{���i����,�I��|�Ϟuלu��t���4��OON�O��_��ت�k/�ս$�H���F�OS�q���j�N��l,�w��������2��t�(�	qt4��|M���(��'�"O�cm����(�<�9�i�+�̬���Vi�����[��
�4��$F�C�?Z�����5Na5����]e�]o�����{:�P�L�A�{h��i�,Ѳ<'�����!�ǈ? �<0xy	��)� PE%RܨLD��/��"1,�X�!�bF�� H*zQ�~ ��~�I���x�+�2�<~4�����ձ�k��Ǩ�RQ��mm2!���b�Oa$�A���E�C���'�r�凴��~���1��w��FnG�b>�/rꈌ♺�k'���4�Jz����1���'O;����Ss����iM�r��F]��7�M�ST��d˵m�&���-��߮�9\��m*y�)�}K|z���r��;��ɚu�}Zx�?W�`�-ω�~IP����ΤCI�����Ӹt}%*`y�~,�규���������TZ�;�gߡ�뮡�ܧC�d����m�b�󣒞+��~F�u���u��:�<�̼�/:ۭ��HĹK�\m�$�!)�u�m�|�z�>y�N��V�0��+�<��.��u�����sT�}M��VVv�~��Di)���`�r|���:����y�j��Ќ>�e���Ia�������/�$p�e��ݹ�ž���駓�_���ã�J	í4e�����i�v�� �Y�eUq����n�>u��^G�_�??8㭴��Q�e�y��x�-�����-_�UTC����[���r�k��ߩ�Skon+M3m!�a�g����8��YVe���=��c�[�he�c��Dy��?R1mVj����L1��:٠N'�ѥ����~�˗0q�CZ����3L�H�u��w�m���p�W�����������~|����:�N�u~y��y�[u�b7S�wt0ĕ�:q�z� ����fx����aȮ��)��Ɉ���S������vp��m�llj�E�8j&dQHW����A�!D��)�ӛ��w�x��޽YǑ����ΘS(��S�����>t���
/gf�~�O>���c4�����[v�`�-��˕YWm��v��]]6���{�q���0��%a�����y��GϜ~~~q�[iӮ��>4��㇧G�o=v�nG(��33�q���j(C �d`�'���(�Y�[�´�{�km)�C�g��΁�m���a_R�Ը&'��R4NYĒI7���+_����w#�6��lA� �dc!�%,�ݸ�x��w��ݏ��ϲ�x_'��E����vw����|S�8�"���w���~fH��k\�Lb�NԜ[\bIOR��/���d�V�B'��e��y�i���wr��͖�H���MR;X]T5H�Mc2]��A���RWVW`_��cE�*2�+á
uî�L���`;j#Y����D�a����!w�{z�9�r�7�t���t�㎶�Һ�:�̼��:۩h�3S��`�Q�Z{ڪ�K;)�6O�(������rrCȅt��l�eʕ��~����2��f��$���f�WMS'uVɚ���󵝲�ޗ��s���U�e�Io�����;
�/�;�h��QE���'\�SN��w�bIO�|�qk?V_�Xa�*���_��r�q�kq�i���]q�[iӮ���<l��:#�j���5$�55��s�UD>�>2���ގr��_0�Z���������a��0�:G����7X��^�f��]5^�����tKi��i�	�P�l$�b�>Jb���-gͳ�]4���q�I��0���M}OοS���А�"}��[���嬻9�nvQ$��`�����vM[�}V�i�ɗ_�_��un����8㭴��Q���_|ztt{:9i����Y��3)�����q$�Ag۞�D����|F^����q��+}�ϱ��g]Ix�5��^�Xf㹣sI�����N�"!ܲI;���ks�g ��<��_8�Q/T�}M4��uT���r��٤_������K����[�}&�L���Ҙ|�+e�Y�9V��j�S�I�ѓݎ�]Uo{Z�v���/ؓ�/�m��k	Ǟi�����N��I��0���_�/ͯɔe������ˏ.0�[�aǱ$z�c���/��W�:�:���u��>p�:�>���|��q�8��I��/�.<�^�y�<�'/Ǯexy�-<���k�����O1�����1幉���U����c	O�~*|SVp��iG��
|T�����u~-~a~O=s��y~O<�I��y���+ˏ/�����&�����~����/Ϟc�/�<ż�^+$�d���a<L<wRy��W�������9��q|��d�ˏ\���y~j����<����O��8�.�[�_�<����<��[��Ko�������Š��-��TId62"�L�Ɯ�DpO>�q1��{�G1�N���~y�fO߰F��\9����_��vj^]%�lE�KWЋ�����=zD3�Ӕ"���bejV�<�=(�*�)�]7���$�/�c}-�w�ϳi�Y��)�
]P��A���?%i�g$�"��Q�A�����İ�2��U"ώ�����m��I���#�9���i��Lrۉ�jd[��$+��5�M����ü�~�ߖ�OE�d��d�����KG������p�Y,�3'+�v{�����U���CϞN�͛:cx26�"���Oj��㻔�j��<ן�1��E��@�	1S�>!���ED�h��b�6�j�u�Ht��!Ad�`�c��D��J0��&Sm~�C?65%��:�/}[�5���܄��[�0�b�K+.��i�֔�f�Cx�l@�B&	F�kF�fc4�)*�b�rSj�,��H2��~ff	�a�w}�߽�������O*�_�33=�O*�_�33=�O*�_�33=��<Q���0�:p��Qמe�^u��o1�LLcO]�&4MG3\2�J)I}ak3�a�m���%.��,u��5�Q�O0l�Y�R��t�R#�.B���X�jBԴaie����:T}���f�6��cٴҕ���[�*�kfl�S�sץO4��Y�3����e1�Y�c�j�FYM��[o��-ٱ�(�ݽ����_fk���A�ҙ���f�6T�	��)C>��!�I$g����N�`��go����'	#3.���N����L�,<pO�D2vOr�pw�����@��m4��_���*p�h"D�p�(�o3'�����t��9�T����,1oF)�TC�a9uq%��l��Y�[�=L3O����\�����!n��d�0yk3rG��&1�&�����[~�߅�\n�9`��t�*.~QD�����ﮮo:�9:�2C��s�;�4����a�:Ӎ4������u��:�:�̼�ζ۬J���I+7+]wQs�UD9��∘i��;��d?��pC��^Fhx|Q��~���iJ	h����'���;�ӰY��C�ߣ����z����s�$���;{k��'�0�V`p&�+*,�*�&���d��������v�qD�<6��-,Xj�<$�����%ӻOvM��m^�^�v��O�5[BV�|�wl��-�u��~u��u��:�:�̼�ζ۬�1{�l1�� N�B���������	����l��Y��~�|~'�D��06=0Uv�8��ge6�uC�Y�0���6�F�I(L�DF"��~�!HG�/�'�����l�3=�[�aÄb!��>��~�M�l�������j�"�M�略�G���tgof��V�ۅ�������[��5�u���Ǟq�[iî����̼�N�N����C�UQ�w����j��W뮵�$�8�Ȇ���lna��b�(��G����κ;���ߑ�ʬ����^�����Y��rr��ߌ��?[��d���fV�H��:ɦ))uXB�R�)�8�{h���i+��m�u.�R�Y��iq�>�&ߪ�-�ӫ|�矜0N�0 ��g���D��0�S@����0)4��i�[k� ��r�Y��ɘUAR�dy��|(�R�pLM�`�Y\%�F�&�왕�]�Z�.v�TC����g�}q�v
�l����확*�����~��X�Ñfj�����\�@��>[�H�G�lO�`��#�Ѫ~�������SK�ם���m�*��r���u�{�um�Jh�x��	����IL�*�>�����uo�'ZCt�Κ�l�et��I*�0�ߑ��2 h���z��v��.ZQ��snӡ��>_�{�Ѻ���(�^eGl+��֙je(��QLLnf�����e��_���/����y�m������̼�M����R�~����E���nv���zp���a�a����t;�DN����`~;M-���io�MK~7N杤h��{����:�Ja�/��?r� ���r]���.8u�n\2��,>>0é�ϿV��?I��s�ztΊ�&�q������ã�J�����:�Nuu���y��z^����8#��ޕU����i���3��q�l�CV҆�A=3粵ӯ?�-\c�j+��JB�?.�Қ����!~Q��!���*|����R���O�|�=ʶ2Y�-�o���S󓋻m)��-�-�F+g�QL63M)���X��
p�u=�M���#�
*΃��4Qå'��0�:p�D�,<�/:ۭ���%�I$�b����_�#s.V�oE�w�rC���8M�aC���̹��aU8�e��	�i1Q^����+�q��5n0��s��3�xz�`0�{Tp,��.��W��eh�fR��Wi�|9�X^�N-��֌f��ɇc}��5�n��L�{��;��53w�q�r�:��-�B��m�Y��/��q矞q�[iî�����/:ۭ��~�'/���X� 2��&*$�I%qс�3��51�S����&Nm���ڳf!�֋gk�;���b���[~#%s�#����X�d��&�pILA��E��q$�A��.x�U~��Uٜ/��GV#�����7-�y+ݧ^=��s����M�!��~7����a�S��U��L������a�<,���!�����;9��g�LQ�٧�{]n[�~��g�hxCJ}�i���+�|�i��c,5�)j�% ��a�O��|v{�����A4�ЖQ�(ƣ!"K�mj�T"�5%n�h��S:~�A��y���ߝ�b�I&&s[a�̭��?<㎶Ӈ]G]a��^u�[j�*����&9��@��C{���� �ధ����Ӂ�wUfTP��\V��Ƨ-���>^��a��}M!��mD8�U��Z�mr�4�� G�@'��w�	�j��#n�(J�y�
pQZvi�P���iZ���8b��M;[󯸙W������OQo9Ko���y��i�V*��S.��D��i���m8�/4��o<�t�(LĲ�D��(M�8h�L� �$�N	��%��a���0M,��'D�bYӆ�8"$B=�:l�M&� �M������GV��:��YZ2t�vD�d�	D��:A(�"'�6x��8x���K0�`�`�9%�bX�&	�K��Μ6lCB"&��:Yb�t��П%�D�� �!�b�'Q����+��EǤ��/\�∼�X����2I���p*�0�.옑��u�J�9QY2�O3w��-����-\0e�տ�Ìh,��|�ͼX?A�qF��;��:m#�	(S[<�K8iUw���`(N�s���VE�b��W�*�¬\����|1C��)ױH0��^�f8�&X�lOv�?Ox7��ʵi���~�A�<�b~�"E�$4�_U���ݮff{��yU̿ffg��W�\��ff{��yU̿ffg��㇊<Y����]G]a�y��m�����$�!�T������?��a��]4�r&i�~�0�nS�������>�ߛY��7O5L���x����.�L�_��?����$�5���8[
�u������"p���~�P�O�d��4�<��ņ���D>�{�!���(f��<�gfs�s.Ud��ՒmZ�j��?���|��tD�	ӆ$4x��tN�;ꞽ�0�dl⪢�/v�EQ��;�v�O���v%�%��p����ZϮ�����t�7УI�����q[bw�}�����K">9O����I�&j���n�����s��9'a��2�(~!��Zi�Dƚi�l�"J3�#m=���R�ژ�ɌGͥ0��v&��ʱ#4����m���:�LH"hO<'D�zуf��sgg��0ChD2-f��V=�h�76�����R�2��?"�d��X͖�jVܔ�h�1����$�H z���#�A4����_�J��?tl���%����a��O��v�x��DaW�ܘ�4�hf��H�L�4D>?y��̞�ã��b�CĪ�� �"d,r�:�i�'�2u���&�F.e���7N�}2�4����ؙ�W���2a��{�x��n9�/���L)���9^�S�R?�[�;]}$��ɺa��?ag���	ӆ$4'�y��i�'���o3wrI$BSK���gOF�}�\�q��-�k�~��!�q�]�s[�\�1�������s��D~�f���~95M�l4��kKܟ0>��G�7K�vv{��P~�o��p�cmܸ]m�+VB�ѳ���e��}d�>���̚�40aSa��{֖��o6���l>#����rIl��%#zK}KcK�4���,����~q�[i�ȐDП��	�8?g�B��BI>�SUTC��־�3��<>�<�11�ӂ� �u0OޮA�����-���0�8~����gw����HeT	�a�,���i�Wg;��/}��9����KN����8���L���vb���4���m���ߩ��f��e���}^���~����f��>r�9���ղ��Sm�[>y��|���:�O�uu�^e�[u��e�7�x���ˏj��3M�������à���b�,��z���ɀr`uᕷ�Z`�4���ڥ!�J"u;�O��r�a�:��8xd�լ��H�Rۦ�l�G+�^��Sm�����e���?7Z�4�$�ޡ3UZ����~,�X��۞�li{��,6��<��:�N��B&���%���T��k�{R�%i}L�Ca"�)��.|��eoq����B4&"b���Q�Lg���@A1�	RnĒI�K&��v{2Q�L4<&����ɪ�.�A��"�^�8ǽO��.�5h�����=��I����MR	|Zņ���9ů�x�~�a�ԋ~��H�����P�����	�0�N�4�8��%��/���>�i�S������|�C�'c>az��àHN
|P��[}���w;��N�L8Sa�
���Q�m��c��\ѭ����ya��]4�;J�d;�y*�it�4���a��_�q���Bx����Oj��h���S����j��u{0�O��z���*Z<}G�&�9���~��Ѯ�2������]��il�n2���%{��Yj����֍Rݨ������s������f܎�������-���a��-�y0�qSJ��Q(p�d{�Y��&=�c �V2(���Q�}6R�6�[i���~q�[i�YBx���>�i��&�j�U��w�UD,�{>̮.cÇ'F;)���G��i��d�io�N����M�yf��H�<�*r=�Kg�U-0��z'[�sn�ӞCߥ;mlfP�*�=�2��[f���n4�4J��+w%鏦��2��w߭�빹�����N�;�k��'Ѵ%��|��m�Z~i���~q�Y�0J4'��,�y��{������*�����G�!����:1OS��iǩ���Q�ﵫ�H��vp�R��;�r��Nfm�v�M4�73'�?~_�㣮���~֨�=m��%?w4��W�������к����.�'�r|��}��/Jɚ�����i�Ԯ�iP���~����q�y�4�ᲄ��*���ڤa~um��o̿4덺�y�^u�O<��#N�۬4��e��A6A �4%��Bl��0L0Ј�'�P�'D�0��b(M��8Y�4h� ��b"""Y�B&�	DA46l��L �%""tDDNA"%<l���:x�g���,p�%�b%�P�&,K:p؂wdDN6"t��H&��0J�A�3��Ӄ��$�=bo"������cw@'���^����{��ϙ��}�T�R=N��7�m�&c��Z��6�[QH�{Q�B��1��bd��~j�%+9�������ܾ�VR�9
��!��Dr["kֻb�0�^��-�ӭW2��8��*����vm��n&u-��xĴ�m�f�Ңi�C�i��ܾ�k�-���Iݡ1��<yXzA�������5-̡Κ�l�@�GF����1�y�;7y��B���Zi�,��Aynr�n��<�,.PW����%\م�$=��9�4��z�es=3
y^����z%.�Y�<��x�]|6��:G@�,�͆��s"(�=Vb�� �P���p��"E�5�$1�LP8A�"?�*��H�6}@�4V�|v!��V=k\i���.�f��!~;�VTl}�uI��6_Xo?N�g��K�;�s|5]�>�]���ۙ�~�����kʹ�~�����kʹ�~�����kʹ�~���p��ǌ6xO`�pL�M	�ǧ�a�ÎB��]��-��j�4vk��鬭%[Ef%��n��mX�pz���[�B8#��>E���Aˁ��;%h��<��Icsl�bd�k�Q
���lQ`C�(ik�k]4r`���/�p�f��R�SP�*,����V���@��z�.,"�M*��d�4��Bjh����B�]�f=��ٍ5���a�keõkW��.J�\�|K)�3I$�
K�/�Q$��K?��`F}����,�c3��Cl{�0&fbWH7@�F���ݗ�[�ң�$<�i���B{�i����Ρ��(3�f�CNC�ʓ����{�8��D��i�Ð��~��sw�G���x��7L���'�����)�'���_�8Y<�����J� `�8;Qdm�L���q�4O��N��2�L��?Ci�it���ܥO߹.�4��/�?<��8�ϝqպ�0�<���~���h������:m�_�+D���x�����e�j���ڍ�<�}�4�L9=?f��&uպy�ϰ�8�~���t���8a��ߓO��4�u�GX<㭦#�`�q1Tf%J�'�C�iߦ�a��uU�^�'GpNt���㣨�O�Q=��-�:U���ۦ_z�bn\�6�M6��/οa���(L4a��a��U*����,��x��؜��т��%n�|�5x&���Um�JO�5�.�0��2�����i"1�|mm�Yf���i\����asا���a�8������+|�o3���W1'���v������H��J�OSϚG_+������e�����:�h���S4���0�ۏ?2���<��[�0�=<>;>�O�=�Z������'���z8z�!�D�Y��Q�'=���,�'���Q�f�0���,ba!d�n�!�"�?� N�?"�ǐ�`���X"A(��?v}ys|�����xí�LS[^����K����_m��9ZaV�%f���=����DG���W�4��nӏ!�~��)�׶�e�_,�D�Md�Zs�}�}][cMY�0ه��&,L4a��|x|v?{�+�.�a�U͟���)�5�Q�e��Xr�� � `��)��V,�n�q�c��[ST#Pa�*�Q��aD���Q0#0��,���I$�Aj3�_p{���I}���
�G�ne#�ΐfb�UI���ϱ�]y̱ORw�Ǝfk��&Z2d>8'y���;�	��E��ȑ.�y�=]�2��W����z��O�iO�I�u��0O>ΰ��"��г�|s�.������ZRa���4��#
%[O�}O�쩳'��L:��3�8� yUt"�>-(\g9̬�ӵ�]t�����St�h���U�FɌ�YÇ�âlD�u�]a�eǜy�"J��6�`bKm��a�j�4�J&��)ׇgB0����5(����R��i�)�O�~@O�U��y��u"'Ǿ���Z�HW��\Z=^�6�T�T�U���Y���Z!
ԅ���h�B���ZZ���{	�Q�BߪMIu��F�M1MS�<M2���}��ɷiۓ�-[���^����[��4�e��'��ŉ�&�4a�|v?1,
��Ľ*�DI�+,��%勘u�����<���~��TF�����K]�_�F�|�yiDN͇��C��`�|���5i��ܭ]�3ۍ�r�/��z�Od�<20��p�Sx��Y�0�D�xdzQ��{�զ_��G]�b������0�-����i��q�θ�8Ì������q`*wlH����D�(~_9WOSgՂ�)�rSU�c� �m!�d2bL�e�@����1�kR�k<mG9Va*�rl�"�X����G���D�����)D�XvwM>�Eayf�j�i��iƑ��K���V�DJq)�w�ۍ>r-�Z<�z��q�m�u�q���|뎺c� ��p�4R��D��}B�̼�"9�3�ŋ	p܌�o�ıoX7��)(^-O���Z�'P���ّ��&�I$�A�'�I$��>�z�EDh~��:C^�AC]��2�����ngN��86�xb?z�`��ns�HŴ۾��[�����:��F�~��i�f�����m�'$i�i+��)H�m�]e�i��s�����z�-�������(���,;���\qt=�{��%$,����i?�������T�f	���ս	؛{Lט��l��0��8'�	��M8Ì��>hj]�>��7vg,`��9����D�J{6a�J�th�Xv�7�s����z!O�I�)<��˙�/QD�	�؟B�O>w���m�Ϡ����<;'�A�]6�qu�y�O�0�����b� �يJ�ݮ͖�AVϻ��j�Ҫ�krx�:�O���?2�$a��m�T[�bW-=[g�\�-���we���2˯2���bP�"ɂ%X�!��<&�yl��KG��t��L:�.���DM��a��D�8X��,K(K�Y8a�BjI�"&�DL:tؚ4 �$4"m""&	�&J �A�hѲ�6 ���a�(�""p�!�(M<p��Ş<Y��"P�	b`�"X�a�0�bp�,��B��GN�X��a�:A>L�(�A�����B��t�;TmP#?g��-��AU}]�N�'�ỳC���{��qq�I�0���FX��b7����@�G�a߱"�n;V@�D�%(D����W��؞���D�;of����;x��kd~?y)	D���}�h�[�E�/�ݎQ�Z�fP]T��]�ݷ�V�.�����S n|�o	^�`��bԝ����W�nc���f{����\̿ff{����\���f{����+��~��l�:x�	�\y�:�0�.<�Ϟ�jI$���5��im:�U�s�w�Ӓm�AV醞����#\k�}�s������1��֕kG?��iU����G9��cmLf������88o6��9�쓦_>��L�Xa-��U��b��2�kD�WM���a��e�%��I����L���8~ޯI3,��ӄF�Z�ˍS�֏�IH�-���8?l���4hÆp�&	釆x|x|w5%T�F�Ts*-���Z�Ҫ�D�߇`�p�;�+Um,�D��9$h�Ե�{���z���˧��8a�ܻ���NΧ��v��J~�"����z�FU?'���D�lҝB���**�Tu�S�6Ѵb�ir��>�Z4�z'S��ÒXapD��ߦ�3�.nL��=1?C�ã!��6|&�t��	�0�b`��lǜy�~n��gt�\^�Z�7��51�3yn�s��:s�FEY�v�D-.�A,��BE�>��D(u9(Fd[ ]���D�ͻts:�Ub&g�>�žP�oT$!?���'��wJ(��7��q�st�9}�0̽h��
�%�
Z�!W��q��5KE�����8p����\���?FNĉ�?rM�-:�O��#60ө�}��̻����J���`��ݺm�Z2�L0�}�<.�j�h�>afF_SVp�3�s۝Z�{(�L\�DQ�+��/G��grs��zy>G���y�;�?bc���ޘ��0i�[/��8ӯ�:�ϝq�Xq�q��>MԍD�R�̽X
Y�����*�v��d�����FOӳ��h�-��V1�J|�~�<���i?G�D��a������
&N�0��C�u�-����%0�2��ς\x q@Q�AM��Y�9O��)=O7N�L0��T�ϩ֚NA(�����tb覉��s=˘��\l���8�\q�_4��N?<�>u�]a�e��<��"�0����UF��!��">=L:�f�S'�s	���q=�V#���Ѳ���N��]��+N7K��D]J���0�6���?3Z���J���	�F�PT���3��~f�~�"][K��[}[h���4�u,�����kU���t}W��4DЄ�ꤣ%�ǽ�m8���g��mS
|n�[hۡ�(���|�0��NUi�i��8��	���Mh�fx�g�ԯ�1���ڝ���N�V"X���~K�z��5*�kF����|�n�i���}���Y4wZ1�����vl��`��7�݌9��6�S���FD����`���Eύ��"iOԢ0߸�13)r���5E�\2��!�p��d�'!O�=�֗y~��;N-�^u�X�V��4p�Æ�~	���M	��h�?B��A�Z�o��Ĕ'7�ϒ�s���k��ɝc%�)a��.��Ĳ��.�J��vh0a�DK6�I?G[����౒�M�u�H�rQ>YJ�f	ɰ��,�K��_8����M�{G�"B0�F�k*�ZJ#��>�7�xg�#'e8&/^4�o�(���>0�sG��h��}L�ˆ�=���xi���<�6w���GF��R|ܧ6�L0����:ߟ-Z뿓$��'�|a�`���]ɛslL6�ΧP�'gfC�?L˕с����!\�u�q�jD�I�.�e�|��a�ıBh�fx�f'�X�z��m����P��7��7Xa��YI����a��9�_:�cq����Da;�GkzN�\��T�5�_/�f��:<�S�~ӂy
Y｢���>2y�xb"u�7����w���]9����j%��H�z�N�
)F���i�ֺ�ש��G�[L�L?5Ya��%�b�J>s,�?:tч���<~	���M	��Y�����ѽ醚�Z���S�U��!OA0L�յ��S���:]:�}L2�-h�~����.U1�Rtv~�`��'��'ޮ��>H��4DN���p���9�;���.mr]�u�n�J�_0�4���Ft�~]�u2���q�q�8���~��0����%�O��#�L��q���b�ži�GX}����o�����N�S��)�����ӯ2��q��x�x�,DК0م�<Y�O�C��zUX���T�!��8"G?$�)�I�z�|������l[/kDa��1AI<��>��<?��ეޚG�Hđ=`��1Kz���'�:�&���y�X���T�a�XC0EG}L8&����mO�1N�'����c�֮]�3�1s,�5R�h�5�Gq�d���0L6"ɂa�͜�[uƙy����x��O,N6"tN���0�0M�&	�Ĳ��,�6&��"""t�0M�lM(�"AB&0N�AB	D �	�ѣel~d��	BP�DDK0M�AHpDؚ��<Y��,�%�P�=%��Y�X�k$L(�8X�t�D���D��H�gN	�$4tѢ� ��O�޵Z���V��ٙ0o֫�§ܼ��T#H�g
�B%L�0�⎃���1Hu��6���$kݷm�?!XQ$�Hn�f����r��^��D*+N�Nm���-R���P|��I<D"�<���u�����zk�30n�)7�&l�0�����2*^����خO{�����p��#�:�	C�މ��[�	n��g��~�I<!�1�q�JĤ��;X�9Ėc�܌w=�*���^;�%<6����6�{�%Y�'�?o�;1��ly��b/��j-��6�l���)x��\s�_.���E���o�wXﱄ��]��(/, ��ٳH��XHZ�[�R�o_.��Gb2��k�Ʊ���O���e���
�˝]1�dM�ÇU�%�tC�Z�~e��RQ���E��J��%W�
�\�AH�ȉ& :�@�ٖ��p�?gf���CQ����03:�Z�d�ԣϟ��~o/{����u[�ݷw}�.�?'��{~[�������{�[���߽�{�����w�}��N�<a㧏	���M	��Y�ş����'��1�9	*0�d�$�&SML�qh�� kv�uخpE���Q���Y+l�F�1�6_,���[X'�eV�c��l��FɊ3MH�k�^0Ye�m|�V�Ԏmٖ�J_l�|�=�\�u��B��[���}��p�N�N����L#�6�ݳ��me��qM���a`4#-��M��+:��XyѳT4_XІ#���u�F�XM��hA ��EQH����$�� %�$��O�Q����j%�J u�g�sf_N�u<��R�őzr�c-���'3Yy���.�u�]<�����]��t٢2�_�a���B���?C'G�w��;���|Xpa�^CJ#������g_��b�>q�i��Eg6��Դ� Xtu&	��:���}:�0n3=((�C�=)��)�{i�<�^�c߃�K4Y�,��Ǆ�ŉb&��ᧇg��fw&���ċ5Kګ*!��]ǘ?5U�ONJ�}����ӝ�ޘ����	�̴����;#�O�Jgն[�ˍ���hÈ�gA����a�O�D�ߛ/����i2d�Ⱦ!O�? x[r1�C�R\>4�&�B��'G� ��gN�jm�لz�~Ӎ���u�ф~�V�gtēM4�>e��[q�u��^X�"hMl��,���
��UVkft��sQ��U��l�:�l��ݹ��>:�rm�C����>8zzw����C�0N��"*~���;>�y��z"h�:�/��ے��z�|y:><;�̇���w�0��������i�w�|�H��>]2�9R�^̞&�v��:���-�aà���4ч�ܟ�0�{�ġ6l�0ç��"y�ϝu�Xq�<��%|��U\�EY�|t=�Ub'�"�o�Ka�����{4�M�t'|뙞�+n�WQ1���\�L��-�}������pxQ<��^�L<����姄v�����e)��?S��|�ayE��XuM�`� ��Z~q�J����u�[j���������M֏�W�:�n��m>q��<"x�ň�F0�ǋ.����hۭ����v�Z=��Rw�`��̩�	�Ԓ�
U$(���}iZ_m0�aé��0C���zI$�A�*-;PbC8����|thx�
<!-
ʶ �y�Rv�Y�Mqk{BA��3�_;{������h�e�t�����J���}Y�%�b�Q���LG�ף�D��D�2������:��N6��DI�8�ғ�y�����!��J'�(�a�ta��{��$s�����ì2��_��a�.���rn\����~��>u���<xD�g�4&�7��ǋ�=Rt��U1�ݪ�D�&w��0D�疥�!�y:;�TWc�}5�eG��4�eh�-t˝]��7'��q�N�]�z���!�=洞��TDܟ0�I	"�<È�U��~�����������6�&5��^Ns�sm���8"'D����"hMa��,���V����L �1"�3	%b'�A�>)vvw��p�M�F�M��No�[�X�u�,�����?/i��wk�=��ϜGߣ������|䌒�oC"Sp`�/��{�m����y��5��v�t��o�!ѧBu7��M�ȉ��p��3�N���%��W�r'�4ӎ?:������κì;>>;:5<a��+�X��?x��!���g'�8���$.N�D�w�!�p�t#��v�������v���f��*-�Å�N���d��ry-5���O�C�S��m�;�b#<vx_�	�"�?!񧝯g~�8h�&�L�?V)�9���`�I������>m|i��~�6��_>'D����xM	�8Y�ř���+���N���V�E�4������퀣�I�)C�@@��T���vf�X��j6��$��#'�g���j��jAU&3y����f��%�_>�0R����:kS��v�e}%�pp�&�/g�;�3�:���^���zHMz�e�ڦ�zM�W_-�#>�.�{�����u�]W͵OS+Dz������ò��<)�w$�:��.�������ݹu��_��mʷ��9OԶ}˹v�2����T�⟘��Z>Y���k��\�滷,¦�N�ŷQt��G]��i�J���I=O8��oο?6�κ��<���>y����}�|�yNr�+�Ï��=��I�t}�������k̯r��viɇba�/FfV���2ãj��>5�ɇ&p;N���\J׳d�K����	����}��n�cTY�N�=�L<�'�ƥO8����g��Ș[��-u�S�;3
To��p�I~���!�q�I\x�ȅpؚ6xâ{�Y��8`�&�6pC�pM�'6h�Ӯ��0�L<�/<��>���q�6"a�K�btK6%���!e���"&���EP�$4"X��N��Dt���L�����N�	d���DD�,MAH'D؛g<Y��0�Dقl�bX�&%�f�
,N6N�(D�"t��tK:"aӂpJ �$(M(�HC��&{�=�ΔVv�=ߑ	vLՙ�M#�m�;��%��$r\�����>�bZ�i���xy&4���@��B>��P�$��H�A��\�oW<�/���Yײ�/H �&~���Űyx�C�^w�E�\�������5�(�J�K�e��5��dg?Fu�3K�b�5nxv4�u�a=a2N��zy�������k(Ybi�3�Rn�&bM:�
��^�9ww}�����{�n�﾿{����y������{���������}��O0��O<[Ϟu�XqƟ<���;�$��7�B8ü�a�7�#�m�en�a��O���~���n�U����F��O�����n�f_'G��g�/�����&��o���D�Je8d��tL:�B����i�'b]3��[q1S��͆Oƚh�t*��6�����7��ǫ���q��8��:��<��Xu�i��>b�1��$�TF�Iv~�?zy�sf�E,;����Q�8'�$�JN�*�á6c>0�J�qa��y=��brL��Knf�����=R�����)m8���%vH�t�O��Ѫԓ�Dc���8D�	�Ӑ�N�J'G�Cɇ[��o�{�w��p�ޗ�dD��l��xᅜ<%��xD��O	�4a�O�Ϻ������r�����
�O�{�l���46׮��u9˥�sݒ��ҷ5���>�w]�Ԧ��n�Z���U���7Ka�^o��W��[I���L1��o'Ԕ4��`��.8��Hǔ#+�39���ڽX�v�������gUX�1]�W�����A�����;V�1��)����תFu5�k�i��u�q��n��ҜF��}�ax�I�q�-��������,ʹ��ۥ�=��a�䈉��w�_�G�`��!8�(�2��3,�G�zlxw��|������2�n:��_�<믞y��a��n[�g�25K]�h+����J�:�{�Mޗ>?N�D�����Ljz�R"����I%1M��n柟rII�Jv�}�ǟF�5�7��}R>�#p�>2>/P�4(�n�V�˟�u�V�ޚ���G{>�	�0���b�����i�>97������+�_�2G���F��o�i�|��,��g�<&�ц0Od�
�ȹK��8>�Ub&��Z���z��/#LV�?f�N4�?Q�)r:��4M�D�!�������B�K�l���N$��L�{�{D33���,�xό0D�4��:U�s��(�!��I��O���{��:��<�fqG�h��~H����W�Y�S�?2��m�����]|�ͼ���8�����Y�c!��U���]�w&�%DO&��j��s�U��W����sCé ulR(�{l���h����w�Kz�p�i�����:0���O/��t%�m��m�&sO=#S�:���i��pa�q���s3�
&�%9y�1%b\:v&�V��q�]~u�Β�:xM	�8`�<w~�lɺֶ�%X.A	H��߰'�a	'F.v�*���牍o��r���+��&khDenq�*L�Ig����I?F��g�W&���"� �o�{�l�Ъ2L�!@�{aձz�/WG������=��cm�|Y��㦂�����D'���u�q&S��*�ͥ��>���%}Í�Xa2[0x<��@"q84h��́'��U`/Ժ��7���6�����h��[]0C߷��w�s	���\�+��g����N�g�'rt=�vl?+~Ի��jM8�Ϟu��<��0�8ӎ���ܩ)R$��v�V]WUV	��9�jpaN���y�m��O�C�=��j�5{�˾��nv������)�)�n�l�,�X����2!����K{:�t�^��&D�~8��ntxp8 �L�i��/ko�6]<�.��}Lc۞����6&~�Y�7�㳆~|�ξ~u��<��0�8ӎ���:]�ʒv�e�2�יִ��%����q�\r�.�-�T;]e�ߒ�c>�����%�""����m�fc;���}ݶ�O���"�=�E߰pFS���޼ݻ�u1�j�̝}$.$�����}[=��q>K�L8s�ؘ&&	g��Y�ͼ���8�o4��ܕE�H�J���z'6�(�f��+�zn���)ٌ=<������O�p��%�Z"J��S$_���P�>ù�d�#:�#^�oϕi�MW!ٞ��sȹ����{��w�R���9���۞�ٲ}a�@�#
�%ᝤ�F�P���/k�9 �E/�Qb�UT"I			B�����@��ȹ>�XG�h��HX(P�t��B �a�<�����ȓ����Qd��<:�$��!��!R��J�D��,��B�!*��!�EBR
�J�T%!�J�!)�D �!)A*@��!*����!�T�"������BT"���B�)!)�D%T ��P�U!)�%!*��B*��*JB*���!(�T%!���!�P��J�%!
��!)�EBQ�J!%T*)	HB�)�B�TR	HD��%!��D%!D%!JB��*�)��FDFDA��A�H�""#dA��Q"0A�H��0DT�Ȉ�$A�B0A�(""0B$DF	� Ȉ$"Ȉ�" �`�H�"0DFD��"D`�#"0�DF�0D�ȉ�$�dD�ȉ��A� #A"DH���0	�$F��"$�"#B#H#@F �H���`��D�� �"�FDH�����`�#@F�"0D�FDDdDD�Ȉ#"A"0"0DA�"0DH0DF�F"�"$b ���Ȉ�D��$�"1$F"#"""1$�ID`��HĂ#`��"#�#D`���1 �"#"#D`�0DF1Ȉ�A`�")HDJE!�JD)�""R)�J"*�dDFDA �FDA"D`�#`�D`���0D��2T�p(Ȉ#A��D`�A"�A"��"#""2"#""0DH$b"2"#DA�D`�#A"��F���� #`�� �DdF0DD�2#�" "#" �`��$# �H�D� �!�%� ����"1"#�"Db1DA�""A����ȉ�$F"DdH"2""0D�Ȉ$dD��"DdD`"#�D`#H����"0"0D���$FD�2"DdD�#"$FD�D@D��� #@F	��"D`�� �`�!RK" #�����#" �`�"#"$F"D`�#�%"""����"��JD*���"R �0�� #"$D"$FA"2$� #" #H����"�`#A"	0D�#"$F�$#" �dFA"D`�P`����I�"0I$DD$b$( �D�0HD@FV ��0�a #�D9i�Dj�2�J��%!���BR�D$"AhJB!)��Cx���!)�Ȁ��A�
�X�0D�D%BRAu�BR	HEBR���1c"@A���!dA�!	D"��D%T!�1(�!*��P�J�D%!	K�]!EB*����$1A�A�� Ȃ2 �
���!"�*�JB�Y	P���"���@��"�"!)BT!
�BR	U���B!)
�%!J�!)B*��*�AdADEP�P�%!	HB��at��!��C�!	UD �dAb Ȃ�J�B�	(��"�B��JB!)	HT�"�(�!(�A(��"�R�B���� �� �"�D�D%B!Q	T�BR�"��
�JA��JB�P��BEBR�T%!(�EBRP�%��EBQBT�!�� ��!���!R��BR�JBJB!)IU�BT"��"��*�P��B!*�BU@�!	U��B��"�JB*��B!*�JB�B����T��"��TBRU!)���T% B���	H"�R����%!��BRBR��B��JB �	A)��%T!��BJB��)A)�!*��� ��J�JB!��!)A)
� �!)A*���B���JAJ�!)�J������J�T%!P��� ��B�@�BR��P���%A�JB0�/(J ȃDID!	D"!) ��2 �� �dA
�B!)	U�BR�P�J!��BR��*!*���BJ�DD" �A�A�A`�DdADD ȃ"dAdABR	D"�TBUB dAdAdA�DdAAD Ȃ0B������!*�(� �	"�DAT!	D!�T ���D"��JB�!)���BR	HD%!Q	UBR	HD%!��JA*��� �B�B!*��J�!)B�B!�!*	HD")ڬ��2 � ȂD! ��B)�"��BR��EBR��!	P� 0@bA�"� �b�"�" Ȃ �B2 �"dA��A����B���"�T!*�"��	HTBT"	HD��$��D1A�"B�B!*	H!	P�J�TA*��"��J�� $8�ؐ��,��ɥ¢^��	�D-��ň��� "���(HB-�JjI����,vg��ޖ�g�%q�y�P�7~~�-�S��>��!vi��?�������-w�Ad��W*h��P��i����MCv���SYB�`�{|��ʪi)A��k��f�QE�M_<����q����z��?P���lQQ�% �� �F4���x�\w���È'���%�J/�	���]���:߳^s�b'9��QQ��y��>A�@� `%pd�G,("m������u(�$�*��L���"Q(����.�N8a���À�T؆��o�ޗB�5����`i�(�8��.�eQJ"��TQ�J(���b -`�tQ1���b�!X��]�x����U���nE/��U�G�Zd��Nh]�<���t�C0�Qp�U	�U$"T�@@YAZ@�QISi�C�tp�b-�I� �< G���;W7HA�b�p0(P?�X��>A�~�Ef�D�EQE'�0Ĩ���?��z�Ç��"���8�5�Ap:/)`�N���P����&#�$_�������P�|A�D����mQQ؇4T��/��`C�4�p:1,> ��E6�耂�^u��(���>�H� O��uJ�S�P��a�k��ǆAS ��(`!�.�(({z4�@�#$��7K����*�EF�ǀ��7�s�F8����%'�J!Ax
8XK���@jJ���>�oJ�L�I|���J
�4P�[o�Bl�<F�rܮ�Ew����+�7;Au��� }��-��S�©�	�x�iZ���h�����x���*���>!�v�l�
�(��O� ����W�DQGx<�������9} �<����i���.�O��B�7d�H0�R0�8v��7��7�!Q����P� W��!��a{u&qH�׉S��0�%�R�n�>!�����A6��]81�!)�l5��`����5Tv ��NI�9J(�z-��+UT���Z����8/�^��"��?�1O+W�
��L�P�ެG�K(��6��P3�~�.�&%�8�6�^��(�;��@��i��v�w$S�	�39�