BZh91AY&SY�����ߔpy����߰����  a8^}   �T       ��� �!N@�  *BP
 ����Q)E	(�T�ҟB� ��)J�#`�hj` �� ��T  �R	� Q@���q��^ܺ��7Mws���-��Zc�w9ǯs�9W��{g� =����liwr��w���נ���)��w:v.���� 4�`]�n��l x �� ���D���>���=�
:�� n�����t��m�$v�� =����l݃�� �7 �{�<��v{�� 5��(m�������\h�vᓹ�:-�N� �x >��=�* �<�dV���M��7t(��m)��WE��t���ݟ 4�m��g�xh�l�{Χ�{��/5w4v���� 9{�w|� ��k�����k����x��v�(�ڎ�΁���7w> =\�6�i��85݇v�۴�ڞۘ�v�kv��s�ݨ�����燷*�νٶ�Gn���[8+���;w&ܺ,
�w> =^z�u�J�P{�Q^�q̣ua��@�4�2=��j�Q�        �RUT*�P    P P %OI��T�T41 &#@ɀ���S�%J!�0&!�0F4ɐD�*�jh       =	�ROS &��@� ���$@MT�jz�D�4OI���S�{T�eQH4ڥJQ��F	�M i�������~��m��I/l
��-���?y�$������C�Q 1�i������Ap ��"̈�\9B"��H%����k�?��?�
9
����=$�$r�* E���Y)RI:�2�* h�=*xb����@I! u �� �=�~#�O� ����+�?���~��,�vs0�\Ώ�c�4o���V�擸u=eI��4��s��;Eѱ-/�S���t���� ���ɮ�u�#=&�NT�t��,H�6z���<Q6C��$�e��hq95�L����{Wӥk�{ ��ra�Gy%��;�gQ1ܞ,�WND�%u�L�${77z���S�:���U�c���uXp��Du�'��DD�5�'�*�<����OT��{)0w���̮�N�DG$�AЈ�O��+��:����i�F�D��������7��D{1�2��z�X�nR'[���+�ʸ�Қ���2�l��%p�0�CZ����R#�=��i�H�[�H�uܬ8;�:})~ܮ	oe"Z��'�]��i�H�})���L8;��:Y\6m�D�H�ܬ6;��i�H�nR']D��nU��V�>���nW���-e'K�+U��"m��N�+��u0�f��ND�m�d��N���qʮ��2�u��R��܉Z�<]O���ܪ/H�'G�T�=�WO�W�ƥ��$�o��7�=�VɯI%A��:Z��%�Z�oQK�JE�&c+��"9���M�w��M�Q; �Ovu�x:�rt��Ïe'�{U�<ʤغ�D�r�1�XeDd�l�Djx����0YFE�L2�c$0�΢-U";�d��NȍD��6V�dQ��ع*�ry����4�1yyRN�D�,K��ˊ���0�,��ؐx��+���9�: �A\Ah> δ�=�ԇrC�p l�(�8�:��a]E֤���&���L=
#��=�t���D�Y.{�]	�+�����1QJ��%Q��x{�*�a֤�h�����x�]g���:����Ea%nSuF�n�bq.���'=��lA��}dpg���n�O�w^�'5�ORO&q�Y��"u�=�1�wg1'S�d��Q�	��*�MM�v���g�aΕ�&��a�I���æw�'6I5z��I�ؙ����$����m �y �$�u�l�����Vcrgf��r¦�oB���ɴ��ry2�Ol����-!�i�Ru�<���3]d��2wY1��'k�+y%��pOq��=�8x��'u�ȗ��"Y���,G�O��l��N�e		�&i���&'�ŎΙ��l�4���9�t��	�I��M��E�H���	�9ӆ'��c��o�sp���6�o���<��2�cFk�J*�znD��%��1(��Q�Q5eM��"{��^��s='�Jq'z"lH�:l�A"&�=����D��Iq'w�">���s�D�x��D��X��DLD���"%u"L���N"&'
<,&��"'�"l{�1&8�4��H�"P�t�:X��DH��%�D�v$Do	�e�"&q"tyd����ćQÅ��H���DLzI���Y�N��҇H�<v�%�i:l{	�D��<C�G*�H��D���	��H����$��
�#�Yx����GU�~��r���DK'��u���5�K���8!��Ї��J0�N�"ba{�D��'N�'N�؞N�)�I&"U�˜">ʉ�0�'
���Y�COT��"^y�-�S!�j#�D�<2`���.p��p�&D��Q���t�9n�fMl��D���TG���	��p���}<'2P�S���vH�Ǻ��uΜ᳉Դ�'���V���Ĥu���t޸ar"<�D}�B�J�ZRDD�yᲷ,y�$Hf���>8�S���w�z#��7ڜ���jp�'�SO��>��매�תa��TN�S��A��d���r�r=�n�x��;�zG�Q,��j�t���yQ,鶪QBP�u�����\6tF]DNzY�]UJ�R�G���쐱�^��';�$�TN�:smM#ڨ����.�#֦X�6�I�b=��DٶA ��">�DK�R��GuQguB3*X��8A��#*�(o��D��jp���DEʎ�/�J8W�G*�	ҞT�ڈ�I�
I4�$���<$D_T��Åm��{Uu0��j"`�N��5�!wUǼ��^��R�Ʀ�AȞ6�J:3���iDGd�܈�u(F5�m��{U�	�p�8t��G�Qje���tݥ'��ã������t�`�����ID{<p�	�|�J�0�k�	��w�<�2�u�6Cڳ��F�t{��DÆH�TL�S�=j&ډ�L=�<v5:^�Y-��#$�u(�	D�7F�j����}U,{3�p�L$�=&�D:K��i���h�a֊��S�%�NyQN���GRҒ��9&z�c2��H����9�®B8N%%y),�Բi�5�5�4�����
����A,D�A�/@A�p�H1��Z==��֌ƌ)94g*G�#�H���o��F��#|��*7ڍ��py��:$D��a�Ҹ$o��F�Qr�9R�3(��z�=���h�b=-�ޣk�����cSލOcS��/	$9��ݡW	�\p�5��npBU�)�g�E���������OQ�"�j�C�C��H�j����)�̶9�t�N�r'�q�̎�U�gp��".F"�\���}~�{R=�R*ɣ�QS�{1�.���t^�m�EDY�w�Lԏ{	ȉ
ɺEB��(�Y#���<���M#�Kl��Fش�8g�3���0�[6��ţc�"�TG����{KZ�͓�&G�f��a\8R4�e&�V�y��c���H���:�N,��3f:�6;ܭ#�(ۨ�5G���'���D�b#�%eJӯT�m�L:ܤE�]6UΈ��V'<��΢#��Å�K�����L(}���R�6ܤN���Xtw�Zt�R&��\��D�����[+U��H�})���L8;��&Ȳ�lۨ��r�1�Xlw���R�6ܮ�"yԱnV�V�>���nW���-e'K�+U��"m��N�+����S���iȞ�Vɮ�N���]d�T:EIwiW�Q�xgK:B�~��xX�ԸX��`��X�`�g�Dx4a��rt�D�[&�$8H �O���j���ڭV���%�o�"�1��w4��JÙ7�23�=d�� �wÑx��s�{~����=T�$L����'���q����Ӓ#S�$L�Ba~j���<�9��gf�f���̃��H9!�;�rA�L��v9��'�/%�tsG4^��'!�D�'����ʢ�TWj��ຒ}I>��iJ�q��eZWt������J��Jv��R�4�0�$�$�$��}ev�J���� 4�&�����{Ma�`�h�HW�B1��$7�b%nv�`����)9�'5��[8+i�l���Ya ?�L1�Њ=dY�|1��&���ROS�Z�<:�K��W�]�S������W��z,����<)i�)a$�[*D��+�Ng%���H�ׇH�uu(���a:l��W���t1`��'>Ѐ�a�k��G�J��7�w�ǂKu��7�;��|{regM�/o��)�����{��f᳅�宀 ��&�$���8opT���#�(ܚB/dC��.�c�!��QHBޛa�N�S
P0<�S�	��k�>���gN�i����O�۪�d��0��lc��~�&yE6f�WS��P]E#Ǻ�ʔ�K��n��I5����������%�|�����)'jt٭��P��"��s��y`�٣d� 6���Zۇ��s~Jd��M|K-��[��*�]�-ᓞ�'H6n�'��/e�D �L��G��ڏ[�Cww��[:l�f�ZÆJu,܆[t"g���g\�9U�9Ѻ�Dup��]�x���E ��I{E-�gn8Q�3���R/�ک���u|��V�Sg�U:=t��Ǟ$�D�n�[YT.�c��
��Zl�s�m��v��Y�V,��u.�Ǯ X�f�3۴͒I +Xn�� ��Z}GwuKJ�'��G���e>xٮǅ
XQ�śGԜ۱���U��Sgw]�#��Ο��@��f�p�7w1�G4��l�V��S��p�E����Q���8ʳ��8aE�||:G��QLr��xl��=M����=�装
��(�e4f��Y���r���-����ag£l���[.�gJ��q��{��xQ�O�N�1zkM�G�_o���7f�=!���tc>�F|E��O7Y�o,�/]:h�|�xٳ<p���<t�&����x���:1��
3��`�b�<<=�γ��'��|�J4lW�8EU;i�<Y�0��G�|Kk9<+1�(�c�����g�����!�"���^OM9S7�����iӳ��4�@�8C�@�ݏ��b���w��Ã4��{S�LC@ �l�k'��;X��ρI�
>ӕ΋(���q6�y%�m<½��}�����8�݌JW7�k��z "_��͒��Ul�|,�� JO9��=����<5b@Qf ��j.�$����A:ٌ(@�M���YF�{L=
�Gw�}Ǝ�|�6Y$]�ZY U�Ei�'������ V,8I�%�<t��H}������F�4@�����|��l�#{#����h��F:}W��: \Xa�ᇎ�@��]Q��)LUk�Q�d1@!��OFb��y8$���&�8�I���eV�"�m�R���ڤ(鼧DQn�����F�J�4Y� �Vl���F�g)<n.,8l�Y��O���h�mm�G�\��(��!tÄm,=ͣ�#�ki��-���[�
"�ΕK�KrݟƦ�>l�b�N�a5L�4�L]9l�z�_aמz��� 8��u��D�eL�`]�5!k��\��K1Z�1|^٦A'�/ӆ&P(=<�V�4�$錆��5>o3]2�v���^� ��ڧ	'�-�A���B�8xtK������ㄐ>���HSv|4�'�� TT��^h���]�\���a(t��V�0���@D$O�2���Si�.��0�9�(����"U��>�E^�(�:h�,��ҫ��t����I�٧�'u��3^�{+5�HQq�g��WVp�u��,,��~�t�ϳ��R��0����'d�D�/�9�݌��`]�+p�0��sM�h���&k��'�=F�o6�I��Rոx�T�J�.��Tb�wZp�=�nca�m�ч��
�qz�z��Ż�at��8��ᇷN�������sլպ{H�_;)J,�UO�>��-�(�!FN�zJ
6p`z��������I^ms�t�gz���Տ�8l��:x��q��h(g�_N	ig+�|�Ξ|0g�4��t�z��(g�"�,)����*?��x��p����'4I�g�i/&V2����V	VaGL��8n�H�0��n�G��Ś;��aF��Yf�*�����qw>t�����8Q}�B��.�����i���:���t50�|3N�慮��{
��0ѫ+�4�Sʣ"�;���.	�i��=�o��əD�f˭q�e�p�ne�Q�IcU}o�4I�B&$�G���a��{�:t���2��HpgI�{��%p$��d)�4Y�1a 0u�.�ej���x5#����ч$xfc�g�6@��������������$�O���'�I�zr÷�ѐ駥'~�����`i�8h�R��KÅ���:i�{d(� .�<Q�����g��p���4==�ri��ݞ�4��}��c!Æd8��9Ҹ�h�'_:�����I��Oi�ӆ�x�����:Y�C@��C�� :h(��p'�3e�vy[7ώ,��*TlR��њR���FO<���F1����L�- �H]� pew�
�Ώ	8}�����-��$�,���%<4g��HS��Ѫ�OJ<8pĩ��NI>���@4�t�<1xO�s�}�pd�4Y��:nS�*Ο�>�Xۺhg�`�`vJQ��zd4��փ:p���o���G6iF';=�٢G^d��xz3�\��=��W���|d����i�O���;G;Q>�zY��k�x�Ӧ�<r<I�QP��3�����㦋�˦i��{Kt�4ă�o���<�ON�xVBy�Y��Ç �������6�xS�E�>������B�O �����Q�NY)�gƜ�����z:Ue�Q�5Yp�H���Kzx�|�<���0�M�$�Y�Tpʧe��f��,j��;��ZG�d���<I�.;0��S�Xċ j�(Çj�M(��˵	�U0�,#����c4pA�t��P.8I}��KL}tџy��~��u�}������Y�p�zS�?0��!ۘM���>2}�dr��y��n�$�0���z׼y#������ÆW4���o�����l����a��mt�>�2�: bZ�<�/6y�ss�6l飥�v�UQ�٣�T܆����O�p�f[h�'��f��o	b�bo6r�G�\��l<Hzz��xSW�4
/�^uYg�j���m�S'�ݫ:���!�8�r;q�F�Q�GJ��ZF���� ,��2a��8r��n^s��n!��8x���tɋ]�:h�K�,�ӇH��aV����M.j���s���d��;\�_Bh��(��������7_�)�l���N..�h%E�I����N���_��T���� in�� �{�� �|8m�H ��R�z3ã����czt�޲�񢝲�@�TI�3�\8`��\�Ͷ�B��}P�9er��7E"�>#Hޜ�hxdx�IE�I`�G&=p$�U_U�^�.Q����4l��$u�o�<^���qN�;ƽr��?�>=\��b�����(o�_�g�"���~���O���8����'��T��@_�� �J�����oZ��v�n�G�Sbi9���W&��C��3�$s3\����WI"j�c��ZuJ6R6ڶ^�+��ĭ�P3P�ЭL@�^��̂�Ļ?@����:�Ɏ���h5V3�R5E�A%�A�Z�!��(�gL�mw�R��N�bmF*�+�A�H�fH�ɶcZ�����I�ڒ�;�mj�c^2�y��X�ە��5���+�^��Z�hz���&��g�Z�T_T��͔�����r���������Ę�KD���� ���H����/�E�f�C)��D�g혠6�0�\��^q��LIJ�2� q��P���D�1<��I��������8YSMĨ�u��k����1*b��q׉y��S1��01��S���)���"�13hX��H�tA��)��,�uG����Q�J� ^�<W���j�x!V4�]����ҺȔuŕ��l d2
�ڲ��!�IP�3!S�҂Y��1[ #K�A<u�C8v�k���	oZ�J�z��b�L�vex�b�E���4��ԡ�FkOX�#I7f.M-KkJG�H��$R(��^`���AA�
5��W�c2G�F��4풦�)$���2�M�

�H�1��⭅f3Rŗ�1Qh��zfzyG��#�k�L}Ο.�G冨t�����b�.��y�"Tηl�g�*���w��D�A��f����J�Wtw払-'����Ȝ׮�{yy�� � ��T�	�A�1`�Irc}��Td
 ���v2����E֤n�F�;��)ȟMMG�+p�A���)��*��-
�A���������p{�.2�c��Z��C�h��}֋[A��P5�LK�T@��V�WK����-�n�s�v%@*�����M��SU���&3�w@J�A�G�0�������C��?k_���YEU���K�o�؂���gn�̇���������������"/�5?�P�D�����������_|��ZUUq������������]����Ux�j�U^��Uz���_u������1U^��V�^+J��U\b����U�UڽW�*��iUU�*��v�����UUUUb��"����U|��54j$C���D��	�
�E�$d��2�$����! $�Ȉ@# ����Ȓ�Il<��H�E(E�CR �MkP��I��hַJ�����������J��ZUWȪ��U�UU�Ҫ�Wj��[U^*ڮ�W�ү�����1Ux�j���V�U�*��*��iU�W�Ҫ�EU�Ҋ��ZUn��V*�⴪��v��X��������T-�8�U�4HiH��H[Y�Ҭ��"ԒZ%�X�jK,�h�XKQjub5ET-�%����&���T5�M��4���v��V�U��V�[Ux�*��UUTUUTUUq���1UW�J��[UmU⴪��UW�{Uz�]����ZUW�UqU�Uڪ�Wj�Պ�����9�<UmU��V�W���*��iU_,Y�։5�H�dE�h�H5��*��HK�>���+j�W����U�U_-*��v�ګ�iU_+J��b��,UU�UUTUUq���]����ZUWȪ��U�U����U��UqiUx�j��[UmU��^]�8�UW�J��1UW�J��[U^*ڬԚ�3T@�UHUNQ�%��iU�U���$[!>�F�"�gt�Ȅ��EGd�*@**U5CU�VD�-��bN쐨��$�$�������C��@�X?�����?���� ?
������?q���,�3��l���A�D舎�DJ�'�L0O�p�B!B �"Qf�Kb'��a��`�&	�`�&�N	���DD؉���x����6"'DD�8$�tKĳgM�A(؈���p��B"pDL�O	�,�f�ؔ	D	D� �!�D�AĂt�IbQFa��O��� ��"a��&�'�	��A8pA����_���Y%�1;EcL�l*����	"U��GVݵ4m��Ev�z�	��:��^ Zz;9ۯ�a�Oa�-��x�n{7:+L�t��v\�|gzMm��A�n�d&�M�l�w;�݊�#��l6��[�%���㋛<f��m��d���ń��������=в񶍽s�nl�w\�Iآ�t%��9C��BFB�D6I29�[�M�v.J��s��u��S���;�s��n�5�y��v��Wrq����[4-94���2ۋK<��g��ѣ��۞q�4x�vU�ώ��Om�`��d�Ek��6ԓT�H�ˣqʝ�	�
��Դ�#�ձ��m5�ݞ��T�n���iN�v�8�:�k�6P�KZ��D��%�FZ����M�rX��j㴑�Jq�Of�LnA����7;ٍ��gsh�
�\�Z�mFmvV��ɻO
�}|��r۳�9ݺ��Y���q���Z�M��6t������ ���ە�e�۵�s�W�y5��@ڭǞ9���<�6�S�ku�����k��08��
��V��j��ρ9}����m�����Mō)/m�<۶8��:��_�ݓ_:�ɷc�e��ņ�ڸ���`��=q��\;C��|�v��W#�����玞�7m�v(��=v�[G���l,q�y���V��iy�n��P�
��s�r��=d��v흽��xh�5�LpBX�Ҩ6�x�n ���.��_9�8�%�r;�:훚�6�[,f�P8�᝹�kkWv`	r�\�d0�ەQ���q�l�W9���6�ssѤ-��u��)�j�*%��x���V���������+��.�ȘS��5K��V��tQ�H'Q�f�'��ǝ�8�}3�������d:�8]�*^c����CV:��;f��9>�X�φ���{m�X�n4���9�T:*F1֢�$c��L)ߚ�9N�c�3�i�u�p��n��96C$�Zr�`����Xn��6����q��S-�y,�7 �;ѷ%�lp:0n�n��<k;�v�ý`�����nͺ@�iOY�۶s����=��tS���7e܆��ëm��"�=v���(��oc��^I]������`�89�U	�7h��pj ����
M����k�dЏЛ�M�m�O8���vz3���*nn���"r���Z��5����b�ƣm���!��m��O:�q`���da��E@%P���u;�M�q^�`NU.Ǝw�뵧�����A�+:#���r���쯀Cvݷj���;;���b��Ƨ1�;{e�rq@�>����v�ӱ�r�n�:�<ヶ���ޛz�5-^]yc�&�8J���v�e��^"�Z���歰��v�%����W����mVB��/e�#Bm�����0[�7�}��p\����L���{K�6ٛn؎�Q�u���'N�.@��!ͺlu��Yq�Ű�D�氻��nQ編'�u;�^;mvܼZ���3�h�ջU�
�L]9�nLlZ�U���'�&�5�i����vH!�ֺ�y�ׂ2�$�(� ��1��8��������i�<�"uSvq��n����LLi�6�bw�Ӕ��E8�G:�m�>tv1Mr���jռ��9��g��<�0�dl�m�����+Y�X�H���#z*�9< �p����8�;I`쒍�*Fע���v&�	 b��z6��uѱ�F�m�n��nµ�q��#\=�m�t�ת��NP���omZ�@�ӌ,n��i�`�U"R��O ;�{����.�|�g�u��㎰����ש��6Ƌ�-����,�ɷ�r�tcu�RB�����j������j�7g��n�b�DG�jR���z��k����}�tKG*����%ex�q�+[�j�^+	��۶�rq�uj�-�r�E�t��y�������_'��04�q��΃��l=�d�4.V4�nU��]�Zۜ����b��"�wwn|kZѣK�U��Uq[��s�4kF�j���*��*�wv�Ƶ�kK�U��Uq[��s�@2Hh�+鎘�q�8�Ɗ0pcF�0Xc�{��/�Q�ё���x��pk+��m�\�5���֪ۭ�E&_j6�ݭ][n`>�A�.�e�TH��r�p���!T<[<qy�u���5���s݁�A:��-�\�D*"C���z��f7vD�a86�x���Z���0cͻJ�^.x�WIōz�Nrۋ{��e��d��ڛlh�֮��Y��>�ύ��	�O	��Ŷ���@tq�fݲ� ��n#<�G��/3��M>�{w\��,�����k���M�5����mʹ�^�W;�vǺ���^�(�IMT��*&�&آ}�	�Vֻ9�ڰk��1wm�DN\��z�<m¦���Om��zx�
�rc��+����g����މ��F���GG8�.�ݞֈD��h 4� ��!�[TPq�>����]�,��Z�i�7�V�ҵN�!PI�ꭃ�`�d�7*=�������rלXr��%V:��6��'h�t��>��Vku%�P� P8.��p�޿c�y2থʕ0�������p�:䉄����~��zA�M��{��p�H�iWtnCfS�գZ�U�d��#�.$:�6[A�xM�6a��4���M0�G	�M�%�4
�����L�'h῜vssI�c����q:��������Lt������|���Ѡ��-rIV�	�)�:�@ �� 1u�?����t���0��F٦/qqW獾B»R�|�H�l������{^,z�x��T�Q�z��--��w%���Ihu$�B?�Z�wPK�*/������o�^ V��qo�C�p�ܟ/\�����I��g�7s��O��]֨�6x��b|'DD�0N��0���.]¦�a�B��<�bbZb�Q&-b�@ PPO�{[�(質k~Eϲ�}�Ɵ�*�-!j��g<D�%7yG�I�.L�D�	�e,K�%,D�[Rq�Qxff82ӃNM|��Z!M�`#XL��L�(6}9*S*VS�I$8�u���te3��z��l0d��_}�����\&\t��u��Gwr�
Cf͞6t��舘&	��Q��ь�1���S��m:��V�WF�m�i �ɍs�{�1uE�km1�&�,W�s*��[��٣��իa6`N��dy�	Į��d?\1VMdǕj�����;�؛z���f�vIR�u�0�!�g�i�l�%�ԙ�.�P�ZYq����z,ޞ� �6xم�	��0L,`���`�����aB5R�e���Xʀ�n��,b�1ƣ�ѕFख�ا�9i��J�2�%IB-DA�I$�2���G��Z��.�"�-9�-�6(Z�\��X�v�2�VvK�v3k7:ҹ֝�s�;8ƫ7K�(t��'�o$ZƖ�krg#�L��T>%P]E���8դ��ݥ����0H(5�d&HL����ܒ� �	�b�a- �:D`�����|��-�wkRF|��?s�� r(����0hhM5(�pМ�X'I�̌t�H�Z������̝L94��I$p��J�o���i�ydyg�-ڵ�E�b���Ée���#|%�^#��^�H�,׌ %��!g��6%�0N���`�<%a6{�lhv�-��)� .��Y�S�8�p��]�-^,��*Z�J+� 7�F�&�C�����!�l8Zl���*���t�Ԛ
ry�c`��' -U�7�2�9���ģ pŜa��a.��8�2Ph	D��/'�Uѿ��r�^C��f||'DD�0O�B���I�
��T���  W�dd��Z�pLt����m�/��5U%L�"*��"�D��fj��f���̘"�Ň�N<6XΪD���a:e+T}�U\������:~n��r��0��l����x|*/��-[�����\K�Ū��2�4Qǘ�9&I��,�Ԅ���Fi�dӲ��*M�S���h�|l�gK>>>:"&	�x��A,0��8p�4+Ub�y�xE>$�H�
��f��%ɦ8_��׉�^�s߱l���o��n���\���T򲻔+���M5����dɼ�Ma�e�[�N-����p���$�ηF���p9��T�TJ�i�HM%6�6B6����Sw��~ޜ^[V��,t�նcl�=�bCFFʪ(��:2���Y�ϋ4`�舘&	�00�:l�6�bf1 ��P����I�X��g3�手�������!P�-��*�v�$�E��J^Y��L8�u�n�FE3Ej�����__9����,�Q�Q��ƪ"����x��:]�k�ms���:�*ՖSJG���b�v���zz��cn\C��ΰ�`�3aO���]�*S7�V�����+���;�K�"��		X�� n!nh(�r�)���$]}��	$���m8c���.HȜ2�&��6q9�U���td�*�$<[��j.��,�ɤ���g3������p>�3���B1����eR7�y�w>W�����t��t���z酟��<&C�M����#Z���C݊� s<εp�i(�O���l�Vp;�-�|G]4Y�祤6�J2�Kԏ2��Qu	v]Į�a5�n��G��!�4��c]��\%QfI(�d2|;U,�`�^�!Z4�4�6�L�#z���/$�QiU��� ��d^-���Y�`�g�!�D�.�[̒q�2hm�pHk!�RL�JpSßt�s^�m_,�b��/��X���ս�K�j�X�V.3Wf:���z֮5X�.:k�q}cX�3V��qqƘ�V�������j���UcJ�v����-�l�V,��w��Li������b�cF>|���N=j|�^.8����Ŝ\^./���c�|�v���/�i��k��^.ߚ���_��������x�.[X�X�^1����z�������~_�~k�i-~k��\x���5��ǭ4\ZƱ�tƱq}cX�^4��q�O���ƽ_^j��ݸ�LV��㶭��t�YXԫ���q�\Z���e���b�zV/��c�����9n�[�t�e$H�Rx¾'�O��(��|W����j�׬k�5n/i��o�k�x��ƫ5eb�jڳ��
��U�W��_��J���[�1q��g�d<���������ᱍ���A�M��fq��)/��Gb���R�tyU�ِ_C��*?5aY'
�u���W{q-�q�o
�Q��E��
X׷y2�E\CfL�G9�G��2Ƕu-�^�W��@�K8ݬd��鮡�wpp�F�ǎ��n���d<^��}!yK�H��!&o���x���h@�)�O���N_���"cx�{��{��o�����������w}��I�h��ff}�U����Ϗ�]�{~��������V�~�����{���&�fe�f}�U�U���������&�0�l�fa���0L�`a�a��5�9�6�m6�4%��u���19wR86B1,������.Χ��Xi]*O�=�ɓP�X�K�C����� ��P���-:�h�H� ��'�EW�70����jb�EON�'����)ڗ����N�����B8��'�G�ޝ2��E���M!���a��NE礆��
"x�K�����$Jt�b2��]L/��JxT�Q׫ƭN��Z���t�$)���뫪��%ۄ�����|e,+ܞ���I�8 eH�p��Xei�Q��^4ΣGK1��M���bl�Y���t�xæa�Qu	|�H�#Fr4�M����7!!�"�0(zt[�җ�6�w���/tsvX�p�=�$�P���Y���m��j��#��StId&�O�Cd1
8u��R���>"!ܒ8����W�咗N-,��!�	���b�i~ɒ�P@�<�)"8�¬��:C%��l�$�MvI!!�
N���ַJsR��J�TomC�G���jưP|E��~���� ``��)pF�Ⱥ�+M�];�ȧ�,���钡UV�6�l���SY$rY�نτ���tDL�`h�pCC�
"ldU�N�Y󲵱Sqs��噶RT���潰ྜ���hC���M���5��r�	B� �	 �[�{�FKV3{(V�ھ1�#�*����US̨�W<���n�wf\����#H�UV9�Gm���V�7����������L�Y4�Q����Z]����zgu�k��̷�����TꄀP�z��).�����ja3G T^H@*;)4@�G��%OI0�"�D�r���bJ5��B�U���'H�rX�T������Qܫ�^� [�0�0��h�#�͡Ơ7
���LK���'�w}��tA�0�#��H��4ѓ�"="�����J��$�d�[,>`C��$z�s���ı�!�u�H���*@�
IT0aF�����TTb՗T��ƈғV��J	3u��Dc�b`\ `b�!��DXff�����'�Y���l�	��0l�Nx�g�O4"&��00��<l��{���ֹ2L��[�6�m6�hX�P5�Y�e-����T�F��z%&X��c��G���%�����A�]�UP�i�X���D���z���+�(B�F!��)�dC	���)8Wt�IR��u75��F�8�g!Je�Hl��Qq-�A�!{)1L�(���)�G?7ϑљ�n�qe�W!�pdP��A�r�D�oĵ��a��p@��B�h���!����o�j���Gr�WK6��m*{��O�/�{���g�Irˎ\:�i����H�=䛵�	�4XdY�-x�jO�N���Ο�>q��D�a�<Q�������l*>�e⩦��6�m6�hJ섡���. TZ�h�5G��[,Lm(���%��u4[d@��#�
�l�a]5�ғ�G�aC�{�����t�)�.�-UY�*'"?_l]!�ɗ��0	�!�*�����
�D0���P {�)�U�cY.�e]־�mg8��\0-!�SN%-���C��W1�H��)tC,��מ*<Y'���Ե4���]ĔZ[��011
>��+�C�,��0���,�(���af���4A9�I��g2Y�0�"Hn��a�l���#VXTB�%����k�{6C�e�,��?�0DO	���a�^˚�u�m`DtP`���1CwS�8�(�����
 ���B�&t<QlLA�������A7����)�-�FC�E��4�}LM�6���/�뜲7��Mk��WVݶdXj�VE�VNG0�m��C��ɢ�iD�U
��`�e�D$2k�U�"��l:@��C�%'~�UbZ`��m)�k�a�.H�4�Eb�6��LQ�J r�	C�$��[��i���ѯ����i�:Rʖ+�ՍRض:SUdR�%QJh!e%D�f"e�~���I��6@�aک,pC5��m���J�1\W�]קn���Ll�����tDL�`a�<|x��z?87j�jz�i�1/]���䡓�()e	��*᫥TE\�M[-`$q$�UYt)Rd�!��I�I �v�'������X*�mQ2�*�]*�+�`�BS�pV.yp����[��A�B���m#4Yg��������`U��^ܦ�Q%�fea���]Î�sm��m�( �
uVQ_O�^�IRJ,ETL_��w�}|Q�����i�x���d$Lǐ�eT�C�m��!!��+���抉dB2cD�"�f��F�
��Ym%@����ƒ�$<^����ra�BC��*$�u�QI�Y)}e�%���wR�]�ÆKi��6�t��_jz�g"�Q
H�K��h�I�oF�7�T��n��H�(vl�p���e�>)
!��-z��h��6@cq(��L0pB�Re���%�^�/��}��eb�j���*��ayҐ��:(��J`�����TC�O�sl�t6a:l�g�8~?D�a }�5��{����{�@��ի�z2bH�>��I���`�r����)A��8m,�����bS�p&�`Zv>rl˲ˉ�p�I�r���:M/�����Kr�3FҺ�t@2��)n�s�M���ǩ�A��=NS��Y�������0� /������N@~���:����R�Vɷ@��-0�.g�W�RB�0��F��6vvo禂����4Jh!�!i�杤�)>��m�:i�ؔ������L�t����%%�M[x
 Y�>,�gO?����"xL0���:}�4����*,��כȷb�0�	$Qx��v���§U�o�O������t�WIIf�!o%(��yK:ZRYԼ8r���� �)�xl�/	M85E��Y ����Z�O!qL�[�ч�vj�!}�(��]�1$PLB1��H�U-|��Eu2-�w��M3��@t��R�Ķ�Q��1č�>2�-��{� y�~9RITU�#4�,�%%��z��*��$B�[���!�-������գ�66� �W9���=�����_*�-���eڙ p��^�8m����!���lD���舘"'���x���^�6z���`J��o9h���:�1�chI~Fs>���d�ޒC����'�U��m5�T�$*���聽�r]��/>�tC	���4o&;��KKm6�+�X�SF���HV.���}�&�$�s��@6a)�eiI'�ܱ�9�z��t�}�'�&L6ق������ia ɨI%�2h���i�I��i��8@�Ѡ�f�F���`�!���Âݐ(�R r����H�a.3�!������%,���u��M�T�n�|��vƧli��O��
�t�5f5���q�f�4��cMb���k��\tή8�n��c�����4��=c^��z\Zƪ��q���[�L+%����b���n�k�;cN���b���W�jb��^/�n���f/i������q\\^./�/�5��{\...1���/�k���ƪ�qzc]��Ǎb�5����qX�cN/���q{oW��i�������Z\\i�~x���/��ƿ;k����5X�./Lk�1�/-��_��lk���N���qzcZu�>0W�ԏ�<a��!<BI�O��W�U�l��\Y�ұ|\]|n��>&���Y�%#Q+k��5t�-cX��^1֗�5��j�Wi����z��b�²[r[f-V�W�j�-�4п$(�a���'˩��9���:Ub�@Ex���t�.+N�udfJ�լ���ʓFnb93'��Fr���E��׷��!5SF��g[uc��M��v���a�f�-ԗ ~߫�'b^l���hе�{��i��w32��wZ����5=�0J#F�Vo艙�� �v���/�Y=�c�y�h�3�b�r����wf��+�.F��7��~4�^=���+�[�ߪ�z���ZYi�oSՆƋ���y�Ý�Q�2�BE�؊�N��2M*P͝W.���i��6��_��'����q���	�JϷ>W�~������O{��C���ڧ��RB��!H�0���1��a=������nѫɮ�V�H�vw��������q�:Rd�7$�	c�C�eֆ�QwϾ�~�xNWS_��w��~���Uv��O����{�������}�]��V?}�/{���32�3︫�U��~����ffe�g�qWj�Պ�˻���a��6a�����"'���x�����JA; �@Z������<�gvĮ%�]/=5������J�"��n�z/R�H��4[�vY�{`���/���uD��q�Z�]�Wv좨Q����!��{Zص���d���
��,[u�(�˹Z4�:n�U0t�Y�-V��AF>x�5����F�]�M&�g���@r�]��_;,b�Ek�a#�o[4�uE$�r(�����0*���`y��%#i��4#�AZ����Z
4�`�:뵸�@�t�E��Ƿ,�Ow�ȵ����4Q9-c�-�<gpVl�IY�s5욲�^
���K�i��r�N�VЫeR���`C�ע�J6�YUʛm�W�D��X+��A��"�����aka6��Xܗ" ��y#/�ш��(�� �Z�����~E�4��3W��g4�;��Z�T/m<�ҕ�<��M��<�C�𔯥��s5Ԯ��:���ڌ���O��e�k�<��#����ɜ�N2����n�g��#��.��:π�Lԝ�-����Hk+X�j�L�TYo��(�.������4�Qɧ	w�>�j��ݾ��Җ)՜|Һ+�������~q��-$M��ҒӔS�<��w���%i�^�h���/(��+�5��ل�<3�!g�FH�|���
t�JN	e�a�����ْ�M�$&�=%Wؓ�6���ݘr@�)�ɛI�4Φ���*������q�f��P�B!7�I�MS���by!�3����z8��V�J~n8�����S羖���%���
{�)��G
>>6~6~����&��00�><@G-���UM�n��eJ�*T�@6ģԐ�Yt�|g�Btk)ad�<�~�(��{���z��.(�Ƅ�^��� �*h�x�-ɭV{�bpB^�H0>�884};�l�j�Ml)�!�In�iHd�ԁ9�]�UYE�:���q'ٓ�rY�6PB��E���\�C����H�����P���:km0k̋��0+%'[�Y�j�@��ROLm0[����!!E��씐����4�� d�vSDv�ES�|�,2h�.H%�d�����V�$���R�6��4Q��,������O�L�`a�<|x���o �By^DG��y���q�pc�1&���K��8���/�ESu��$��N�,�IYL5��%& ��g�&L��Qԁ�qSA@p��%$p���)t��(��Ɋ0D�iE{�RUB�-�R�2�i%� �ěh�B�-.�[T`�*%@�HBG=��ۑI�ĤAM5q&�Hf�-ɷ�*�e�HAmD=5�JR�@�zD�i7�$��fKL�b��`ŋ��(�d9�W�ړK%���V�}f)ڦC��ԨP�:C04@�����I��Xs1+��a�I�8Y	�0;��w9EUUUe��)8���~ц�c��i��M��@�05��8E�4`��
��LђG��<��Ӧ�>v�ߞ1���D�a>����[$�$�g%J�*T�@�
"���E'ʺ��M�7U\cQ��hܰҞ�&�:�B�a!��\2��%P��g�ȠGR7ϻ8�֙��3{��O=� )�P���x�4RZ`��
C$�y�X�a�5$�c��d����FaA�4�+If8�	�ђ&LRQ�%�4��qst4[l��{��Y��4�=[��RJ�ۼ�4QdN4QL8�.�Rh;`�r@��80L&"�%�GE&� ���!�Vo�[�D�%Y
�kg��D�6�6Y��4d���pd�dt�GGN�4��:qǏ��X㏜<&C�O�f���k}�9go|�L��;��Z�US��Q��sm��ou�EMۖID'2�E��G�� �1�bM	]��Ų|�~���j���.�ݐP�X�j�ܗ�m�[�vgMb�`�ggU�ow&�:���=�*p]�Zco�5��C�GXP�uG:u���r��	���3��lC@�1ސ��Z����4-$迀�����ڦ�9��G'��"q�3��51���p�J6���"�@� e�ˉ䬕m�0@<�4�td�����S�j��Z i e�e0��Jl!�W�⩭F4�[�u6Ə�q�j6�S�c�ME��9m������o�QҮ�~����=RCLN8i�B��VMu-�H ���R�rG�%J�h��'�p�f���if�����z�S����T"m!F�j�9�j�K��oy�]��M*r'm]�Qd`��yxO�k��I�B�䣇(06@�@,���g~��X�^xeߤ��&�ç����Ο1����>q�q��A,|���H�"P9�l��5*T
 ��6��y+�Kd��@;��2`9�IV�ԣ�,�gk쫩�&x�������8�B�&-��u0�M|RQ�J��D�;,�DB��e������N�;��FG�*ŖN��KV��a�Ձ�)M��b�y<}������(4Ӳ$ q C�:QTR\2F�ĉi���ϧ��ŕ��5���
9?.��tY�?p(��޿��?D�@��8M��!K�p�Jh�.�����e�t��(!��2�0wVy�ԩ�q��:yz�6C$I�8��²[A)�n�h�m���x����q�80p�4h#��lf��<�~5��QcĚO��mG2�����b�=��;	!������h�p�L�ԛKN䪷#� ��F���IG�Kɖˏ�u2��E��=�U���M����5Fb}
.�d6LȓiT%�_~��F�Ks����b��]�j��_�w>H�T�u
	��K�p�����)2C���l*�p�6�a>��]��Z^��H�i�ta�P|�g
L�l�d#��}���1� lْ!���w�Ý%�������{�K&�X�;X�1e���v)���<;�%��d���,�e0^�,�q�0G)�6�5I��gޒI	��ؓݙw����ݸ��1����0p�4h#��mz?D�蘕U=��\�D�vI�4c�1&�X�	����dj:V?-��\�6�ݴ��HL�.�ι*����:y���BD� ���Ĺe�z߃��)ן���)�p��q�I!i2p�K0f�4@��7
"ccF3��6�ن�#���Ɣ�(��*��2g�q!ԇ�iK��F������b�X�b��|N%�7K��⌇n+�UL&�Tv$�bZ�QFl��&JB�@�F~�%٤�O%&�����mn�� X��"e7��lM���*x������YA�K0��b~8~?>>D��@Ѡ��?at?A�رR�E��1Q��+210S�,N7`���j���"
嬖�E��{)�,��(��,��L߻�	�x�n�J�Э��h�-ΑI�*U�����l7�������f�'/ff��c4�h�z��Z3�9�m�N}1a^Ƭiv��K���u����L �4���NQ���Xe�0 ������6���l�Fa�O�SfFV�4�(=f�����"x�E�B�� h��&;x0�e��x����pA�#���ڮ&SDc�`x�!� o�TVJ�*]u2j�l)8�E��6q0Yl�^�*,�$�%ٯ�\ V{X�I:p-�Q2��-�J^�Nf�O�IF�c�Zl���]�M$N2B�.
��>�@�����Mk���~	��IW���/��ܣ�'X��HQ��Dh����'c(�yZHS:H�-1ӫ��������|��o]�c���c��q��||�[b������j��mE�U��»HF+c�*T
 `�IHo0�u�퉿J�K\,,�|�r��D*�c�%W�&J�c#�Sj��G�W�:��@@���-6AN'����|4�hfs�C%)q��3!���x�@�Х�:K^�ͦ�v�rI����Om��؄#6e�\��Uݦ�dk�͚q8|S�6@�Ԥ�����4�8�)8�n�I�u�z�11Dq��������VMj�!����%6�C��G�N,0��d6Gl���I��YtRm��'�Զ�L�:o�fH�L�6E3l��A��\M��LC:7D&�nSP0@��ia�'5Yr`���B�Z�מ+�1^����S�xƞ/k�]��ƫ��Z�ή5��������i�ZƱ��1�./�k��Z�Ʊqƙ��z�^��t�-ƪ��̖���Z�m��V��[1�S�4�x���4�zƦ.�o-�+���X�V8��i���qq\cUq�b��X��޵��X�Ʊ{|�..>k�vƪ����1���./�����b��5�o���m�\jx��[\_W���֦�k�5�[�\\V8���.<kK�kN���_�~_�ϝ~\\G�|��|���|�V�@�!E�t�.;k4t�1�cJ���jUū8Y�U嵊�tƵmb�����b�q��?<k��:��/5�9��iqU�c5zc�\_X�.9���k���jy�t��z���njڬ.[j�j�+�-W�$�	�BY%��7�oݹ�W�߸v��԰��-DYTK���gH���"��Tޚ熩a�Gec�Wm>�G�5�oF�ۡ��y[�M��EJW�6�l'��V��<ZH��w��V�h����:;�Z�+���U��YJWi�"u\ɏ�X�Z�	j�%__��N����j�Kd�Eקf$m^���9�b���t��P��=�ش��O�;
;������!+�|����֫�U��~����fffs3�U�W���ܻ�����f}�����Z[��^�339��֪ګ�io�]�f�0�Y��Y�>>:||&��00�>>�.����1�m�hK�)�$"bc9r�L�ݔD�R�(�i��F,��ɂ�B�$�L����&�� x d0(��XN}��$r@,���M��ލ7׺�@GMў�����F��,�	�:�Q�Tk����i*��5W*����^ �1��Hȧ�v��,<��q��NF��5N��yIh�-��|�C��51T�pm!���e/�8D�4T[ L�������r��fJz��Ӝ��8C��;ɺ*jUUr$���l�k��^��?;O$��� q�ߡ���9��3��%U�	�S)Iԅ�Zb��㷮���?=c|�6�h�F�_hd+,��T�OCwtUQUEU%��%%�'S�#�K�f�h�4C^�Iۨ�-0hh��3��%P�
��1�H@���ru]U�N�Q7^b������r^<e��#�I=i������,/Y�J��M�d6�Ӧ�RQ��I�$HB/HƓDL�&*��M��1�2�)4VR�ۨj�~��ے�	I�.�Q���P^o��7�4���z�%�[�m�0�䄐�>;��.�\m-3��C���&�o�m|誹j�y�|{�cui�ĩ�W!Å�:`��GO�O����`a�<|g}��Y'�M����`A��w[$z^0*��X�U��p�y�+�X:��Y���06�s]�޴�M����#'�;�����5κ�3ئi�˱W�����u�ٯ��goс��R	�ru�x�e��V9)�&x�	zPO��J��#�맧dH�5G.]ɒU�K/ i)4D��t�
BD�$&��ɷ	��0���k��
����hx�e-+�ʴ�e�4�4"�p����[׆�O��d��!!�ʫ��uT]\���U��i"d>��sɧ���^�$6gI Q��&>L��1"d��'6���)��!�Q�b�ˉ�	���4e>�D;�2v����6�L>8`���	D=X�l�4���`�,V����g�!�)�.��j&CD41/t�Rge�*�mi�穝���+æ�4��ӎ�����6�1�8�n>>|��x�$�u���	)lc[޴�M���Ⱦ�
�	����9>)+E!�I�u/	���I':4۴���IX}���*������~��P��Ů�{����	s:z�4Cئ�u�f �9<��B��&T�L�M%ԧ{�a��T�ɣ'nmi�@�B:����D,��0w"�l�I����HI�a��NK�F��F���N;�.���R}�Ͼ2�9�B֤�$$2�����I)<lż!��F�0x�e�4|h����8�m��ϕ�7�+Z��I ���۹�֕�ҾMi��i��Bo��r�tQE�yٿ��S^��Ӄ�نwą�d6G�x��X�4Z]D���M$M�gj����U�*���	�O���e)�%��b��Q���|��o�z�M��;�껬�wl�9_r?f-����ƾ�?f�ޟKL1<;��/��:8Z!�MЙH�{�.T��]H1�Q
C��a"q�M?4�`�ƻ�qt�r0[���g�߆�����:�G�<M�C��8�L6o��	��0{V`2Q���,�g4x����><&C�=�Ѫ�
�ޥ������*�(������Jza>z\�rC��W36M&̴��D�4a�2�G�(�6FOx��`���!���.���e�@�I�OY�L����&$%0�fZB�a�IgL�	���Nl�iI�ű����Q
���z��W��xD����]�tTm��l*�m���?=Y������:���9�q߮��&��r�l����G�S�+��

4YFώ�tۍ�~clccm��ϕ�p�TrD �}'Z�H�J�Z�KF���$��H�$�9��
[�5G~�0�	 ��@��^��6,�=�<��J�u�XW4�Ww7�% ��B`ٗ����@r��O��#�$!Ѯ�V��Vji`//'����7%�ou�֕b�]�D�ݹ{vQ�����&�^Ԫ��_*�x�.Hd2B�N�L�G	�ࣦݾ d�%'������h� �J9	F�J�l�6�i4�g����Q�c^m�qw��������X��4���薝M��l!jI$&j�޻�\$6l�=:!�zS���z��v��RD�(� ��u1�������ة�b��t�z�V�ҽdv���ӵj7�uwg��|պzԦ��t�o����q��1�1�6������}�:���5ƪj"�ab
�Zj�Q�o�6�i��x���Ϙ!���4{E���ĞL&ٔӄ���d���u�:!F���N|�MHf�6a,���8��B|\m/��N���֤�d0nI$�Zt(�!���̌|���h`���x�ڼ�1������	6�����?���޼>�X,��-�t���J(2C�G�0Y���Y$)tcyܪ��e۳&((m�x�6�������8�8ۏ��x�Ԥ���_F�m6�oB> @D'�sW3�5����n��&�	5e�!AD+��s�}r�O�Zm4B5Ly�}��F���"�S��i�k�&�CF���1pÛ�ɍ��
!Ĩn�8{�p�ʽɃ)iM:&d�aj����c���Ɗ�[z|�]<�=� ���>�59ur�����51<Õ�YvIrTJ�\%&Nh�çO%�KJ
!�h��K2d�&B��۷���x���6�1�1��m�E��i(#�d{HQ�g�P����N=�Rbe�dO�kM��M�M������o�yx!�)!g�,-���^W�����V�(�W�"��[�:h����!D"	�&�ZQ���Ȟp��;N���"g#֝�+��u�����|�g�D"c���x���]1���ץq<��p��>����`Q��ӛ(ӣ
!���?\�!��;�ǲ[���id~�k&��f�#Y l�M�`�S��^1�����v�_��..:ή��..>k��]����.:gWǍb��nun/��q�S7n��]5�^����W�Y-�
�m�m���V��]w�kYom1�+��vƦ+i���cG�j����b�Ɯ\^1��jc��q�_6�k������b���\\|�X�/j±X鮘�/���t���|�.+ӊ�qX�[��O������v�ұq��b�Ʊqq�|Ƙ_��5X�.��.<i���/ˋ�k�5����k��Ɲ�/k��t��;k�5-��ZcJ���iU�Vp�
�ۥ�O��(�x�O��M�(<t���:K"mܪH�?�_����T'����W�X�..6έ��c5n>i��OmƽxүK�aX�Y-�Z�,ū�U��W�]Р@�'z����
?!R����6�,�U���%�ݛN�6�
��)@��/�wv�Ne8�0��y%:ʺ՟������lKk�>|i
�鏳c�e
�+U�U(���V%����T��\�;��\*R����oU���W7��
�޻�����}�G"��fc�2�Ƨ>h���l*��P���(,0^�p�C)]+!����CA|��hsP�ٽ���G�x��G�R�TZ�u� Þ�H�1Yaaq,�xY.uUT��R��sv3\����R���Ժ�TͥY-:�[�D����\.2�Qq�71��n�y�p�˷���Y��鵖2�R:�c��Q[�X��7�R6�[��-N��*`)[vڛ��	`�wë��Xx2���#�H���fu�w};���^+K���י���Ͼګj�v����y������mWm�ܿ�����Ͼڪ�V�v����z00�Y��;|��clcc�f�W�c�Y�[���M �q#�T��m��hhT)G�w[M�����\r�2�k�*��H�RE�N��*�`�5��*�-�
EԪ��+c�n��pM��X�ΗP�{M�@v��a����sO9�p����4����6������z3lX�����#y�Ż�絋tN+��ꓸ7!�l��K]�.��s����ݼb�-��z��8 }�fv3q��ՒƊMzI��l�ώ���Ξ�^;z^O	�q �	�Z۪ nV���*����{D\m85+C�IE2����[nx�h<2S��[s�&8;tq����+�zݩ�඗��Uwŭ��T�P׶��T���v�Վ�A�qNe���GgQ�m��KQ��pϤ������A%�����@�h\����ʵs6�m^3/V�%eìBw�/*�'TX�-�D���r�TI���F�ͦ�tqڛ��Z���eں��ȁl��]�һ���Y��`�P�c8s1z����5¯�Wr�_��ɇ.�2���	���b/ۢWM�tѰ�:o'��#�T��,ó�'�SfC$,�����1�]��76���iE��)Ic�� B�h�V^�!ҹ��|j;�m[}KS#ز�|q:S�����sD�x��.����c�*�,�je������!'�LF�b>:���!�xYlɃ����fͼW��;|�<~m��1�1�m�m�׭���u�u�]t�5u��պ*������X�FH�pd���!Z�'�6�������auR]�zi4׭)+Z���$:�!�O'K7�+������;����!-6�2�|xɀ��y
������+���Sl҉����\8t�ٞ�W ����Wq�0�c�J��.�;c6�=Rd��Cϰ�0�f&,�_00�_��v�lc������6ك� HHiWm��A$A%��?x��W����W|l_sR�"ZY�'S�:�끰�<�#)g��$�UUA��&�4ם��!��   F��B G
E9���߫3+�2��q�M���U�[�X�wc|	����0����e�f�^>���ٱ�A<��^�(h�u�1˔�5&ڡu�t[���^!~ԓ���e�p�W&*�5ajI|�������

,�L0x��O<l�1�1��m�z�j��Է��۪�D�dϞ��M���л�lcC�cٓ�۫kR�z�m��qc&�C��`���vV
���x_eK�Uպ>��HI	ԍ�4���݆Hy�L&
L��f��!Ѡ��\�L��=>��<�x�=���A��=�j/66�h�M.�w3��.��u�dL��ɃyiGB�!���Hg�I��
!VpN<0Q��
!���n�{uq��C�`��1�z��lccm�m�מ�>�]��T�5��1Ie�]�J%eDiBN݉��dѶ�Ɯ�����~�A$A%��U��_�?	�)�}|��Ů��(i<TX���TDeY�X�Օ�j�鯥����R����	!�K����VE#�H�$��l��0]ϤR�����_!�Yp�"韆nجRk��7�<K�� �U��]���A��94��J�v8!�H���1�I��g@�����'����TSqeI�yM�v�m��FL&
~N�6?�T����c�n���̝���,ᒎ&~d=I��x�SA�ك	�ܤ-��� �8�U�|ʣ]w*��Uw"WWw���4�Ot�]H���L%Hm.�<_z�,ࠄu������ }���n0�8���SF�+�o�����[~m�c�c��m�z��/qx,�y+�QS��֛i��x������V8�<Ur���Ϲ֚j:�t`���:���&�x�5�c���v9$6��qx�ϙ�D4��B��	��S�h2C�}%Ue���LN�^v��if�tw=*&��i/:����Q�Z��0���0�l�{��Ԭj��$�X��p�o�#��-&B��0�?�xc\���H���WC���Gj�Uޚp���/m�Z=4�_;~v�n1�[~m��X�^�4�rH�ECk�,��m��m�hW���Ěi�2>�IÆ1� d4@�FvQ��Ad>/ϊ��yפ$��'��}���]��#!6��
M!�C��U�Im�*�;�G�!�8�s� IަR���}�M��X�|�l�gDl���i�oU���S�c��*\���&��:�'���b�.\.�&O�m4��0R{������6Ch��̽GBM�ܩ-68<V=x���1�ߛc��m���.'cr 1�b�3��n��*�(������H� @�S��CO��c���Y^h��FcGa!%F�<|�8��C;�C$-,��l��I����Fɀ�^�d2B>�GF�'SiN�)���GR�6m6�0q(6C�ͻ���r�Q�Sx��O� �,��x�Zn̘
 q�u�SO�N��LM8Jc�8�H�C�Ïc��k���G�Q�<;6�^�t�l~~m��lccm�m��~Zg�H��u3G��L�*.ţsw6����l�_s"��ab�����}��I��>?|;%l|��r�Wٔм�ІK�j*Yt
2�WƲp+]M�dХJ�[�
�7C4C��Q���@���d;xDI-�gN������ �m�Ҝ���QkR;�dPf���U�#i�5I9R��M%�b�"f��-��N���#�I,�ڽ�r+n���'/�Ռ�7�����h�&ݚ6�!AR`��R��KI�;fd68M���y�����1�ѝ�#������kElь����Ox6C���]Sw/R\�Yf0ɧf����Y�6a�e���"|�ћ���>/ì��cN�t����cm��q�quuu��-4J��G������2E�mQM[
{޴�M���Э6у)����� Q$��[��0g���C`I$
Hȵ��y����e���d���}�a0cG�fB�Q(,7�*�ܕ���l̚m<e�y8q�N�6C��t��E��_"q�ݮ��v�թo��]^A-ś���V2:n;�:w��xt��Vw'���:���+���C�0��Y�Z{��l���~3��Lh���0Y���b"'�OD�"Y�<X�""xN��� � �	�e�,M�N$N��O	��0O	�`�""a�<p�
�B"`��b�M�b'<`��pD�<X�:'K+�i,DD���b	bP��'D��Q�`��X��bP�%)�H ��Cd6$�J:"aۏ>|�8���c�L1�i�ag���O��<'N	�AAO�B� ~�ݍzO��;�Q�IT�y�X��HSmʌ��cR�q��}^�uq�S#�1[
(&��Euk8X�{�<��t�ګֳ�J^@�G���U��\���&P̗������$��!g�Z8bL�Vq�a�`��^���o�F_�ȧ���+��U�zR̝Bv����i��jPEm�W<���j���f�x�����M[�>�%�fm�|�W��������333;�}�U⭪���������R��V�v����ffff{�Ux�j������a�0��<|���6��c��m�����p�:��I��X�"�9�4�c������Qzz�N�5�d4�U�e2h�S��(��D!��0Z@�8~nSN�$��G�4`�(�Z�~i��`��������5���N�J�$ag�F$("S�ep�9\J69!�ܒOp�ɣ���0B���C��)�fI�錭��!L��1���#̞�W���6�I��Q'�- #��Γ&�ɒ�i��O��c~m�1�1�6ۨ]Ms;�gF.�D�%����p�9EUTURQ;2f#�l�F�v�X�a����I$�~<a,�d�˲�@�2�����x�����V�j��}�{^�*�b������>d�0!�:��i�'�.��4!�̢C�Kf^r�i���d���$�F�:r�4�M&����9�m��%x��
<n���/���	$�Ƀ�a�r�����>�$�6��k�O�M̿?{���j�O�<~v���ߛm�c�c������2���$]�\�*�Ux"��H//2�uG(bA
M�i���U�RA$A%���7��>����L���Lὂ��IXNY���a7�w�$z�>k�pTX¢��˲���oon��r������܌Wu�Un|�c/z�RN���p�wۀ�~͛�����pYO&���wͼ�������Es<���]��=�ii��y Y;�T�T��d!TN��l۲��Z�=7�Y:Vwb}2���M:����!!�4B���gMI$�M��L�w�Ԯ�p�8D���=#Xg��v�5'�w�8�m�� &��(�xg�1	V�*]�n����ą1�B�N6���8�lm�1�1�6�j�k��}�QsdM�\%��?i�*�����Sg���2jeE�Z�#��J�^_�h4lԑ�>r�d,6n��BJ��%�:Ӵ�-��s�̪C��z��BӇ��m���M'�6��-6m'
9�$$�v��,,��ɂ�O��ނ���1���;�Y�����w��r�pM�ܕ���'S'S|&�M8�H���}�_t��a��D��_%�>*J���반�N�Yߦ��?F��Wm���������lccm�ն��!�k����Q�Ppr<��"�֛i��iG{UA��ܨ��}�&8���Q�F�T�&'	�[
��2��$�<KSUL��8���!_ˡ��@Ӎ6���?�*�S~~$M���zxp�m=���t����^.zL8i��p�N:��M��s8���B� :8q|����m<0rϪ�����FCɇƌ��2S�a�䧮�IY�"^������(,��8lå������8�8�m�m=��;�VtR��X�Mݸ�G�F�i��x��%��n+�V��(���FB���|[�x���l���l�g����+� �Ը�KfS��Y��p��n�4}�B�����g�����n]��I��#^;~���@#��E��I���G�!f�rh��ϓ䲊7Ϫ�m8�,ٔ�po�u���G�{���m���d�9;=v�c�Lz����������>>Ǐ�Gu��U�7U�F����%���u~�	�4ɭ���VN��-����5��I���@X�i�r>_g�ΫR�&��������3P�	��6I��	؋���U7&��eE�H����;v��Ң\�lb����B���Ahu�=�wU}l�̑^��֤�bL &���������v C|Kz��-~���N����S)�0�O�'p��&8N�N�!�Ȇ���>�9�Φ+�),����&�r�%��^��t�y6x���x)��b����D������[��L�nۅ_󝲷9�ā�l�5}������d6i�ra���|NzI$Y������c�~i��O��m����lcc|�j�O\y���:���J�����[u�Oy��M��M�MY���6�욛���@��߼�h���m�KY�>�w>�R�x{k�$�ܐ4�`���ӿo��>��6�a������N��䦏�M12�M�rLvI$��4Cg�C�ˈ�@�ph���i������On,�3��Xӓ�)<G���������$7�A�)���֗��a\y�&��Mr�Q۳�'C��G�|z����lm����>m[i�5�Ԑ�a�r���qy�4�M���C+�il�H�JFwׂ��~�2,o�|}UTMU��Q���C�xi2�xPh���S�S�=g��Mǹ(���N�M��k�:>:���ދ%��*��7$�o�'~N�%
��j'�^�:�$�3�Ѥ�%�7$�#/���kV����kNG}_K8�8v�^W�wUuP��)Ɠ���<Zp<��I�=��
8A(����������cc|��m��uƳޝ^��]z2f��${��(�Bo+J�X���Zm��m�j⋱}�n+�ʾO*\Xv�!�!�IY=���3�!*� bV�*��4~x���T�K5�p��v��ɉW�2CO���|�݅�g�;�4`�|`2`z�r��ΐ��:�5�^M����O���Ã�y�ܧ�C}0�8�g�D��^�'��CI�%��:��f�Ο�M�>Oo{���e��0h��&0~6Cb""`�(A�b"tD�����6Q�A6AA�lٳl��6"pD��xL��`��0DD��x�B"P�%�""& �"P��tH"a�<pD�6%�c�p��,DDL�"A�pM����Ĳ�(J�lAA�Ab%"Q��ݴ��M���1�>i�1\q�n8��1�1�c�z�1�N8 �'��Y��ײ��p�>�t�Xj���X(k�.�Wh�X��嵙�,��\l�0�Y�wj����*�5��c2A�%iy
��n�u��R�*Ӎf��x{*i�X��M
9V��wa��]
�)����N��v1�.���7�
�}���O�ϑ�W��\j�v�8A�<����^���yX��]I�L3ى��6,3VUA8r�WY��ȹ�@-K�����ʼi
�N�iv\��F�T�3Ԙ�lt��'I����>�B�+�Z��	0�z�c4�	���<�d!�4�>�UÔ�̗I/ٔ�u�.(I��z�pB	E(C�F��&��(*9c��JD61J�LNV5f@-�8��۞��Ɔ>r��Z2v�H��R��&#+gtwU3jp�/b�W]ٯWz�+��s=�*��v�����ՙ���ﾥUz��[���陙��ﾥUz��[���陙���}U�Un��ײַ>W�>|�󧯟1�1�lc�`�F0!b����6EF��H���^��N�nf�S�q�u�ώM��y��Wm��q�sA�r����=�M�E^�<���ݬV-�Ů�ۗF�W�Bis����4m�U��qYU$��*�n��n7�X:(�pѲpv9v	�r��9�.��Ov�m(>�m���;�a<�<�q�ru�P�n(�ˍػlr��M���v�d��M�*���*PW7LQn���F�Ѳ��7�n�s�8[�5���pg�]�(�k��+m�a;\=�89�#�ݸ�+����!V7]�=��Y��rm"�w]��p�8�k=�,���&��s�v��3�99�����d�'��X�[\d:Ҹ�n7lb�U@�s97�g���`��ch��/��Wi(��FZ�� �a�Ƥ��z<i�Ś�瑸j�|�6�]��	� ��-��ƛi$^N��?q�T>�|���IY�0֝=��Y�.�fqu�f�'E��w�d�׊���Ҙ��}j6��zO9[y�L�w���n��B�#NHf+`רL�&ќ���	�f�=޻Ty�2��N��<\ϐ��B3��j�`�¡R��O�S߰UbI�?�
8�,2�M�1�!��rH[�ÉEPS�ڗ.ʢ�?Eu�IӮ��!
 ZK#��	��.JNvN_���q2h�p<=�I����C���^�LUJ�&�(�UIhCQ]&M؍Q~��/R,l �Rq�^����~8x���Ο�=c��lc����^.�u5�=��nƦ>Ƴ���Z� �b��`��W�֛i��x��<��P��J]�X�`#ă0{�����lmr/-131�f/[� A�q-8�;$%�ncܗG��U`�F����'/�ifd��&��fCh��^lX8>�e����aV��������v]x�z�A����:|a ���U=vp!�O �Zta:t�p�ϒ��=�&M%5e��qvV��M�t���o�6���X��|ڶ���ޭϚ�W���1M����M��M�M\��ClaP���>G��8�+�{3�T�8�j$rx�&��Nm۳)d�:NGT0�Ēp��!һ3�n�U>3�a����U���Im9Ou46��Q4i䇎��2N�'xb�'�s�y:0��5�&�p����j���@�0,|O1����~�Z�~x6�i6SI��c݅!��,��q��1��1�1��6����5�# ��Q�
�H(&����a�UQUEU%O`��;.q>KN�tl�4�?cW��ő|�&� ���3��'�iwgn�9�wy��8v��pud6��j�B�U�t, ���M�]>0Q���,r_y����M2Æ�^�o��ur��UB��<zs��S'�+T�$6x!�>+L������0�U$ԉY'J�$���GCp�j����h�z�>m�����X��|�#3-���XD�� j(�e9�R�IxT�,8�65�'D�ݠ�Wڄ��M���p�|���sA$A%��I]��	��bm��u�����<#?����N�9�n���*��`���K�#�X�Ʊ��7(^�5
������g�2��=;��Z��)�]��\���=yWX�T�Ж����r���Ȟ�a:Ǧ�%4d��&J�FB�Ԑ�i�e���a���^"{&���ԚJL�no<��(�2����	�_�)�l�I�Zoe&�dɐ���g�Y6���d���z���' �����/t]��X�P���u׿r��:�џ4�i��2י��+i���I6(��4|Y�͸������1��>V�z��N	*, � ���P�1�m��0��	 �	/+�|7���h�,�G������т����I�&�?|b�؝R��:���=��	��<咬��H���+��>r0i�1&��i�tb�7Ӂ������34��_��ABq~W3�9$d;��C�
h�1;�^��_�[o�y�[r7��q�Mxmg�G�rz���������W�=m��N6�c1�8�8����O\�9���4�0�ۉϷ�6�m6�5�����U.d��5�X�J�a?/SI���,�6�x�%�](�^�d^�S (/��(���'���2�
�{9����5�Ƶ���4��K><����$��K�єŹ8䁳<쐓F�08zyF��UZCGɗe�����'�U�3���s��ڔ)�t�<N<2�ɐ��`�ㅛ-���m�����cm��|�֯�{��A"��}-�I��<�L�0�Q����T�?6H�ޝ�m(<#�Z���G�]��(.ІYưzBq>�-�0|iB���$j-f�I�#-<�a�)��)2GV��0lƳ*�E�����
=����m2mBW3���Y>Z{��v[�,
u7�.m+�e,��Ϥ�$�z�mG4f�!e2[n�?>co�|�6��o�+枷�U���!I!TҌ�G�k�����TP�3
b��XM�Sm��[
�F*
T�Rڑ�_�Zm��m�B䯐ϥ�l#���k$J�4.oˮe��*h��*�z�*�4/-_Q�8`촊�ʽB�N�k��H���T���fAN�a#�X��}��G-�:0o"4f1�E������Ғ<��x�iɎ�%$��CLP�8x~�g�;�<;)>L�[}B��!���F���OO;���J=�6�rQ�p��䅞%J�M�i3��	}K�:m�������p(��8�Q�F�̫����m#�,2}�R�Pb����ɵ��UǢF�1D�!j�8|i����t������IY'��J�t�O�ϟ�c1���8�Ѡ�X�hl�Q�!�D�b*������i�i6�e���;9�2dɧ������B�N�'٘�(�q���:��0�2��UFag�:2FL����0�F���~���R��;׫m|�8�u�x�W��_eȺ������j#�6�����йr�$�Y�5.:�2��3=�0���_��J�볦�%�4y���Ɠe{R���?�Ɇ�`wG�)֯�O�0����Ĳ�?	D�0O �D�:"`���pN	f�B�A��P��M���'D��`�&ؘ&	�"&:'"%�"t��� �%	��xH%�"'D��%�bY����$,DN��'JD�"X��艂`��L8'lJ8P�%K � �AJc$H=� �^>i�O�v�l|�8��0�+%���D��ç�O�
>�p�ÇV)��Z�9��|�y�uݍ��i�1?#-�<�m*�	�6��A譵������0���v�k-�yJ;d�w���r�N_wd�������-��D�!��;��*�l��A���,\3* �G^4v��_[:��t����Nm
hP��ה;���
���}|�/6�@�|
�ߕ󸬑�B���������y���F �^ni�n�Fۓ��/�}U|������L���ϳ誫�V��ߌ���ϳ誫�V��ߌ���ϾEU_-*�wv�k!�a��a�Ǐ��>><'��x�a]��ˢ���*�Gﾒa*2?$9��o}�!Q�m��6�~G�઴���3��`�w��Ǔo�4N����L8wi�9�K��~�e��-��1��,���\�{�܉��HA��!^�f��u9�1�(��6�F��ѓ�'ܓ<%%����0頤��=������~x��ϟ8��1���8�����m��޷��V[����/�`��1�bb��Q�1Bw�����*�0z��JJx�tM&Ϡ��(������짿�2�*��s�n��~�0���,�Ǳ���UY��m���ݝϠ�@�2!Q� T�uo�p�8w��㏂a/T��n�,�Ÿ��y�����<�a��C�ɗN*)��}�+ؘ�ő�ƌ��I�����S=�O�N=t�����>cq�p��A�m�d6�4���,����om��wJ��PL��rA6�%r�U
�X ��%��i��A%�/�	M��e�(n +9 `D�B�6?��S͎���ڭݷT��k7+G�Zw5�����,Q�)����椞eB8ڍ�uo]�.�ٹـ��>I�(qD����8��P���^��J�I��<a#�d��l3着ݡ����>M�7?p�/�Zs9�\	�rT������Ã%.K$ra6i����{����Ī�'fξ�L�)�t�W'�IIf�r��H�@�N˺�6�M-�qU�ML]KFI�9qo��u�'��!ҍ,���~c�1�c��|�����XE����Wά%w'�HEiW�r	QUEU&�7��t��9���mÓ��Ɏ���	$ �e��>&�ɏ�AVd:k�Cy���	�W.nI!�e'�=����/W��Xc��ʩ��U{i��]'�8�Z�n-]�swŰ��M-J�{�|����a'$��G�S�#��9gc�/�ϧ�>��|�oΛt���6�������0�Wd����n��.�h��e��!{�i��i�����5r=�����k�m����ї��RY��k/O�	��&°ZGF#��|�3R/����w^�:&9�lN&�dy	��m����'�=&uuRU���Y!�qk���q�Is�4�Q'�3���.� �yZ%![�{��\ c��;�����Z�.��M>�SA�D,��6Yӧ��<c�1�c��|����w沾����Z��Z���|i��i����Z�1s4rL&�80p�h�M��ú���a#}O�~vk[��1T#6���#���|���azd�����{�`�y��Ď$��IU��r �U�C@?�lڪ���U"�*����)�1�~:�"s�W�LͬY���4�0�4d4p���į� �ٞ�m���s̶W�?J��J�N6��O������q��o�+潷���;1��%rA�Y����k|4�Vqsy�4�q��(��L�D1��!�=u�Z��+% QF�1�u�^��	 ��R���ۿ���>-Y�e��s�P��+lm��a\z�0l�r������L[�g]��3�ʋwl�}Ukq݋�+	U�s1�'e�B�dQ�n��"�Z����
Ƥ0^�2��n�������W�.�.`�gr��,��1:��K�s�/q�᛫�|b35}�NOa������G����gص!�#�pY���JN�<�06��{��|�<\�Y��=��0�Ɯ�Vͅ��>�:L':HI#-؞���1U�r����+N�a2Vҹ��Ʒ�J��Q�Q�!�\�Ǔ��%�t�;W�1�OΛ~c���c�X�4�Y?|}I!&KͲ��4����O���u���B�I	^��b�Cg�9�m������2���I�⪶zI&
N:�9g���8}�%6t�n�)��T�;�&�T�c_�|���8"zT.#bJ�PeQ~t�1~���u뼱l�k/%~z����6�t><�*Lz�vy8�j�=����t�[�v�m�q�n?=q������6�^!x��x�G���&<7\�Q=;��H$�K��V�2GN6�q�c�GM[W��0��-�kn移�����'�ݺ��P��^�;��m<x��S�ܜL�M�>$q�M\*K�)u��s뗘�U�MC �Ģ�]V��$���F�Χ���4�2��0M|ɀ��Qo���c�5ݧ������λ~��d���Wz�Zv��O�1�c�1Ǭ4h#B�GB
�#�B)H�"^9�QUEUT������!`,N��-����u�:�7<��`�Zː��?$N�C)ƞ���0�eBIS%e�YE��#=Ǉ�;�!�eǾ%t���}$G�BEn<I���J��<�7MlC��� ���`}��i���?VM{~�w�~#߂��y��>5o\t�<M:x�!�""pDD�:P�$�DO	�"'N	�8l�4�!�K!bl��'��0�&	�`�	�`�"`�x�A(DN��"% �tJb"tDvM`���X�%�d: �J6"'DL�"%��0ؘ'��<X�Cb&�P�%K � �A"A� ���8�Ӧ�6���c�i�1X�,DD�""t���ś>���a�aX�n�|k^f��u辕B�\B}iڷ�i�#0��N��Y~4�ғ�q課#���VD��d�%0�Ωt�����ʶ�����O�c
$wq�^��>}qL�[���j�-t*����7�U�1{�n�2Xt��G�G,Q�ALq�u��U����G��5]�_f1t�.�1Q�yyY�������(�In:2�K3�*��������R��F"�G�ⳋ�\p�	�(��,��d�5&iR���(��9�m�i�e�Nj�])=�᳌]�b�"Ս[l���0�j��UpYylv\�dfUW_Q0� -�|��o���t$��{Y�yp(\*V��m�74Z"y��h-��RX�c!�mlM �9#��q�,��Wػ�kپv��n�su�o�k������Ȫ��V��ߵ�����Ȫ��[��~3333>�U\b�wwo�������UUq���ݿkXa(��l���c1�=cm��|���)�{�L�0r��b�VA;�O좃�R�棕@��ػvv�cnXwL����.�omN�V��DhnA"���5B��Y��d��v��͞;\p�ˑ��tڐ ��1�YGn�x�W�=�-��^�wC�u�z�m���n��S�lqv޷�[to:�ŉ)'[��]n&�'#v�=u��{5dk���s��u�uu�qmf:�un�:6:[��Ճ�۹��Lv^�o<R����)�yX�-�B�׹��i��
��1�Ϟ �+W;c�7���a\�V�E*����H7W+(r5e���E$�1�n���kZ�/��:뎻ܕ�[r�i�6����8��m����t$u�M� �d➘M--�vn�f���>�I�Ix0˿��ܬX���p��W�Zf��V�N:�֬�-�Ogs�غ����|/r��;W7�.���)7j�x�ab���'Ohp.H��x��r��;�UWtA7��;W}g�ɾ�Y���Y�l,�(�&C.�AC���2t�d�A�王�4h�~\�ɔ����s�Ɇ%����p�(-�Y=BG���YU��f�ݗD���/��>��Q�߂b���M$SJXё�f<s�y����\�
���M6�7yS�Tg�R$.�Źy�W�vfsX���o|�)#�A�'�nzC�T�p�l�z(�͖t��=q�����m��|ۧ���_��q���S*\�w&�y�r�F{MD��I�mRc	�%Xcrm�>~N'W���ϰ1�R��I!I�-�!:U�%QIf��	$�m"lbYFC�m��aZ�?c	�:q�F������|�{Y[�.�������/s[��`�e\��G`2W_h�5R�O���M�2��L%�4�I��b`:cA��,0��6,�
��,�g����c�1�=c��|��t���,&$Dԏi�� �W �p^$ RH���X���Y�Pp}��}��Gj��箓a��f0�P����c�X�XYX�M�U�H���Bx��|&���M�/y��LT'R&������L;y��RVWAi��$��}��Ϊ�X-6L&�\�D�]��}G�u(�R|�o�h:Ҷז��?>q���c�z�4�]2%ԣ�!
T�Dy�nիV�Ѧ+����s��c^U���{��}��qI�|�#�n��7d�����8fw��vNj�+��a=�UB����$�K:e��|���G9<�G\X�$I�&@��܅�I1r�Pt&XP�	�ڒKuq-\����^0�m��M<[��55+�q4уFpd(�V��͘m�z�1�����>Wͺk�z���WW�D��9�H���zE�X(���|;ݪ�9i8�� Q9麤��@�/�=�y%��ʮ�+�X��ζ�S�[�B�ˣcP܃6�0�֮nwZ�U6�.֑f��c�0;9@���c�8�!�"!��O:�ui���s�3��2B������5ZΪ�T���x6���O���r��|@��N��!�a��^�ޓ	���ݦ��8?$8�,�2x�{�g��f��TJ�%l�p��O'
4GGP�h�4��I4iu��@��
�����o,ʗiZ��X�����=��Z(Ɇ~<�ː��2v���󧮞�q�=~c1�1�m��/TOW���Ʈ�ۛ�Ɓv��HHH�����X�B�L���^�{zU;J���6Lp���I%���j�Jץx)6f�H������®I$%�
�J�V�6�0`x���J#�~������jQ��(J����	�O$�>l�X!�d�`H��0��f�3u8�6Ku���y��b����#^b�ZkY�O?}�'�tm�c�O�?;c��1�����6��mӬ�WZ�kS� ̉�1��� @�q�I�QTUUQA�I$!�ަ�oS��l��<�l���6����]F�'���hƎ�9�����_���;�G思6��ٕVEkw�in��݁�vRj��h�>�qz�XX������u�]]kF|a<��i�F:%'��0��.G�l�Up��٪���QQ~�C�����mȵm��r;l�tۧ?;~|��1�����6��mӽG���4%�1���\"4B�>�7���<������=$�a���aƯ��F��M��]ʨ����1�P�� E���V$�$�!׼4�2���-�S����m��N��q�?8�#�O�|&�e�:y�NE�:��P<N��`��&\�ZP[o�ERQ;��`�,�f�8y���c�z�|�_6�u���κ��5 ��s)��<ܑ~x%�C<W�MS��X���<�ŗAn�U�$	�+��>��~�_�IS�3b�����;:wc��,N����������&>��w5�2d��9�\9��hS��	aWI؎n:�UN����Mܦ;n��&��x�7;;����3-��u��
1�^(�i):ͤ>JN&jO��l0�"��}�I��5g�%%61!ҼUIU���)!�y0ZD��ĳ�Q��у'	ϝ�,ޗ��i�Γc���̆��^<>���`?�r3��]m�N�6�ݸ �ἧ>۹�d>.H�gR.a'R.���t��tۦݱ��8��c�x>0h�F�X�>D��\�-�cR"%��a!!"l�I'-��C���2Ca�!9��UTd���Ή����h�|n`�ٳfʁ��N���y嵥�r=�_Gm���x�:��o��a s�L�9]�]ʔ{n�Z��fu
/�]Ÿ��+�|�y�4D�F2��b�D��LQ ���{
�%I����u2��0;���%���?{,�X�8p���6aG�FDD����t�D�8"xD���8'�&�AC�	BQI6"X�,���<&xL�0L&	�'���D��B"pDD� ��6"'DJM�"tM�bY��� �E�D興� �"P����tK:Y�6A �	BQ� �t �D�H'D}&�i�ϛm�m��8��a�cLa8"xD���8'�!��Y�a�=WƘ���{޳��z�w޾�)���r�۴5ؽ��	�noG�����2>��usK5��;�2��D#���<2���ƍ�M��UyD�{.�^��ʖ����WE6�v��Eht`���i�/w�*��^oY�F��IY���&:�Ⱥ�wrÝ�گM�U �1�<>��n�G����Y�ͬ��*^�;�JDC@�.�V���d/4�Vf�
 �^�h��Q��Ȩ�oF��_���=�eң@��Wݵ�u�y���;��\b�wwo�fffg�"���Un���&fff}�ª���wwo�3333�b��"�wwo�0�a�����=c���q���o�+��<r��?8 @��9��8��ί�m����{��ӏ��v��e�Gx�qɗ��ڸؚ~[I��|@�z��G����7I9�r�J�L�+D���N�B�ټ�B��UUe,��?3�ç&���!��'0�'F��>��� f�Rj��i��!A���W��E9/g��i�x��6����6�1�;|8`Ѡ��Y��4Q����$�2�j��8�O��z6�֡�c�� f��m2���"@��F<�L� �-�i�<Y���XT�?&iɌ8t?zM��d2vI!�T������to����}�^�i䅟$�%t8*Ze�{��-��+���u�4�G%��`��,�g�>�||'�τ�����NA3[����1_��uTc;�Z^EoMFS;M�-6��P#"{J�q4�[+���� #�=�� ��?%����N���ɫ2�;�4jo���͋^���z�'W4V��S�{�L�Z��j�3wkT&pn⽴��UO4�K�8	�-��#��޷�fTt���8�;n���!�6~���ӿjW��u<�CIІ����$ʧpܕ qݿ���@�T|&M�l�7h&��Ŧ��&L���Û���E����WB�Z[C��	Ϩ�Wl��޻���"a���vBM����pN�ɶ�M�k�(�M�z��n1�X�n1�1�<m��|�)�/D�C|b���w�kXe^� �y�sqE��<�ʲ�_�ƛ�OSۜ>�! � 4>���{�%U���)�i���nL6N�#Đ�4L�a��@���=�0��$���� m��Î�3�����w/�4ba#}��r�%a���g+Og$zZa3��c|L�Oө��N���q������u�5��ՙ{�m���dZ�lWՍ��iks�;q];t���n?8����ccx�����+����H<`�� �ϣ"D8"�_g�����}e���q�QF	�Ʉ���IUE^���	;0餚5g��D$�Utl�(���*V�P*�*� bfx�J�\;o��G�L�s�Љ��Up�B�Y1eHB4ji�(��r�D%u���h��g�zl>O~���J�M�m���=~q�����C�h���Q�[�FHj�ҷݶ�X�u&q���ɑڹ�b��G�|�@��_R+Q��)uB&�IR\NM%�^�c��'T�v`rZT&���lH�0��䆹$�-!�Nbp�&����U+3��N��Ml�-�2V<eM:~"c�ի�ӓ���>�~�N�����"r�~�css�l;�V���c��?	��>��0�6a�t1�Dr��/��v�]/Q�W=��s�o@[��K9�+R':නD0K��d�*��I$�����;C��T�8lX�S.$`�TX�n֖������(f���t�ԝ>���jU�������so�=�/#h�f��F�ˎ��]��t����~�#�]X|�FEe����wz�m����g6o��l�E�!��w>�O����l{g[�|l�>6��d�S�$�.M���B����X9��Q�=�Vn5WEܟu6�'{�Ϥ�t�
9�Fe�$6M�퉖ͧO���>�>oZ]�B$a�l�K��f󜙒�$Mb�8�:Gz�����d����p2`�t�f<h��g4`#����]v�vލI����HC��l��e4l��@��D %����}lvH��n�����cf
����鯣n߉`�+F���&�)>"`����1��z ,�\�PDH�(p��@ܩ2�ۖ�P����+I���A9���f��T*��h��OƊ��/����ND٢�ZD���4ї��7��.2�'�2t,�,�g:x�q�q�����m많��\�| I/�@�W\2���^� e?��"¤R�=�;�B�>���������e�٘�98wdz�]�$;9ȄT�7(�h�<��+0�:w���o����GS6�.��/�9��I!~������4}w5�&����/��7S\��~��}����-j8�R|0/�*L0)s�*A����4ڊb�ix�_=t���qǬq��>c1���WC�4�&7"l�t �M'_Q/�R�2e�c�2����Å���:/�id�����S�P2#����Orc�P�Q$~�!��8��5�UQ�!�zy2d�m2�et`/~�A#��`����ʂ�;x,�|�R�e5�FM�Rx���NRߎ���ѢΖ�j����?��Q��A��I?T�I$��X* QG����Q������������ܝ:^hѥ�t���!�����iL1���h�����J�
7��"w-,�YK)e,��4���e)K)Ue)j�eUYP��T�Rʅ�-,��)eUYK*��,��,�e,�b���K*�,UU��4���KUd�T�)e*�UU��,�eU,��RU,���KURX��*��,��J��UX��T�UVT�J���������*�U*�UX��*�T�b����,�ieQ�ZH�R�UUYT�Ub��UX�U�Ud��U%���UER�U*ʩV*J��Ud��J�URUYT�J�T�J���UVJ��UU��YT�,UU����UUVU*KUb��U����T�,UU��V*���XUT�J��UUU��Y*�Y,5DҬU*ʥX�U��Y*J��%UY*�UUVJ���R��UQUVJ��T�,�Ud��%UY*��URY*��R�UU����U%U���*��VJ���T�VJ��T�%UY*��IJ�UU���UU�UeIUb�UR�X��U%�J�T�UeUX�Ҥj)eK*�ʲ������R�X��*�J�
�T�Ue*�T�R�YUVUU�T,��T��V)b��X��J�VJY*�KUeR�UU�J�URYT�UeK*�R�ʖ�Bʪ���RҨҤjR�YUVUU�UU%��X�U��Y*��RR�URʪ���*J��YJ�)U%����UVR�R��T�U�U,T��*�eUYUK*J�)UeX��Ue
�YR�,��I�Hԫ(�,�X����)b�b�*�X����X���)b�b�*�b�T,R�K)b�b��X��U�X�U����)b��,RģJF���JJJJJJ���Id)(RT),��j$��RY
J�%B��%�%
K	IP�%���R�Hh�"��ID������Id�-��F�5*�UY%R5!Id),E%�)*%%B��RY
JIIR$�E%�Id�H��RX�D�*B��RX�J�GT��Ĕ��%��$���J���
K ��)%	IDRXE%D��B��RPRX������IR),%%D��
J%%�)*%%�)(����JK��RY��RT���II),�$�RY
K"RT���RXJK"RR0��0"�	�%%��	IR��IHRY$�,,"�(��,���(��,���(�"�P�Y$��(�%D��
*IEH��(�#Vj��UZ%�EIE"��E�EHQdJ*%$������� A�A���0`��T�T�	R�R�R�R�T�T�T�T�J�"�PA�A�`�`�`�`��! AH�� A��R*P�P�a*T�*�T� �H1X1X1RD�P�P�Q�����b� Ń �1 �X)K*�T�R�,�U,�*�BX0� ă1`ĉb�R���R�X�U,�*��)ևU$�R�%T�R�XT��RʑJJ��R�X�J�*R���UK*�� Ń1`� �X0�JT�R�,�,T�R�EQ�A��a,A�bT�T��J�J�R�X�J�*R�X�J�*Y*X�J�*UK%JT�)R�JT�R�K)R�J�J�R�Y*UK%J�d�U(��d�U,T�K%J�b�*X��F�E*X�J�*R���T�T��J�U,�*�*�`�`ă)1���d���"�)K�YJ���)e"�K)TYJ��"�U*�)T��K)JX�R��J��U,R�YH�YJ���,�R�%R�*�R�X��)H�J��R�(�*R��ևTt�U,�)b��)T��,R�e)%�QE%�Q,�Qe)K(��%��YJ���T�(�H�,R��JQb���U"�b�K)TX��*�e*�)TYJ��EQe*R�%�R�e*�R��T�Qb���I5(�YJ��U,�Q,�Qb���,�U(���YB�(-,���X��%�,RK�(�E�����*�X��(�J��)%�,R�,������j]h�E%�,RX�X��K�)%�YKR�),RKX��%�K�)(��IeRYE���K(��YIe%�T���R��K(�QT��K),�XwRMJK),�)E*�eR���(�RYE��b��,��*�QeB�YRʅ�,��eUYBʖ��,�YK)e*��eJT��T,���UJ�"����}W�+����H�:
S������1� IQ# �Xz5�$����y�������?��ӿ��P�d��_�3�����{����������Ϲ��O��������� P�����?rx6~���Q��.~������5��+�_����?����2����� ?�C��O��o�A?�A�?�
������* �J#%�G�	�������~��!�d!�҄J���	���A��?���!��o�!������ԏ�?�������<��܎�����8g�-
``�ؿ�6����%%'�I���
�B��ַ�A�������!5��2���d����������4��x-Q��--� �ES� *"B*�Ă����$H��~+�Z�o����`}���?��G�� 
T�U@��!�Չ$��,��%��"!h�$P$_�?�������M��~o��?A��a���#�����P���?؟�$��_��N&���V )?{@r�h~����u�����k�q�^�?��ƿ�9�=����4��?���[��p8�/���}���~u��������g��~�� ��G�A ����޲��W�~��z����O�8
� `'��@ ?����Ed�����e�� e�a��8��x�M��Bj�@((���꒫�:���We����@@��m?�G�T�?�@������JJ!�����R�'P˼Q�6F����lR���:���AP��?~�����~g���H����"�pAg�'��_�X����������?�Y�W��-"+����~������C�?���g���� ���G�������b|�w@�����_҅D������(����������;�������@~�? c�g����;IAd#>h��1�?l
 �̟��.+��?�������������?>�K��5�\7�p7߿h� T �����Ʊ%$j'�_��`�c�ࡰxa�����?��_����<�E�А+z0�[�����+��𿤈��1_��g�Cd�������?c〠(���a+�'�?�.�������g�w�e����b�J�K�����o�����.�p�!3y/.