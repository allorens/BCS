BZh91AY&SY�`��٫߀@q����� ����b?��      ��
�D��(P�V�lJB[l���M���M(*����J���fJ��R��e6[m%1m���iKg��� (�EPU�XҋV�i��X[mik56�ղڶ�-����͋aUh�i5R�J�)�Փ6��3TRZFf�*kl�cGf���^Ҡ2�<dR�J�#���%�VVZ[aV���j�[Z�P+4�jDZ��
l�kl�d�1�mm�6�ckU,[F���5XYe��[j��p��e+m�M��    N]�O��� n,�ݻf�����]X��jޫmu���������G�����U���j������ǫ�P+�y�6��k
ي�j����  |�T��+�tw[i+�5�����J����E��*J�E/{����(�{�^��z%*����w�e�*k{��zJ��Tm�w��z)[j���7mIV�M��J��mDBbml�jAK5�  -�>U*�iY�M*T�{������%J���Ͼ����[{_O�>����'�|��J�R]�^9�٨
��x��O��V�v���ىI����B�{h-D��YF�m�����  =���P�R����=�)R�u�y���%
μ��^�ӡ˺��JU@���W�0�aGs�m(R�&�*D�v��x�z�T�Q�Eh�t�;{M���3�dٚ$
��  �[��%B�ϧ��TI��ޥR{-�wJ�:kh�qA*�I�x�T�*`��U-cs�ݰ=T�Ns�rԪi���R�	��OZ֕Z�YKݎfѣ�  &��T�B��f�Z\�z�ީJ
�oy��ʤ�:�x{އ��QK��wM�J�í�^�w�Z��fSǝצ�%)���M�=�=�b�O(T�����kj��Iel�Z�"Mb� �w��R�R��z�j�����*��=6�G:���=��SZ�й=���;�c�z�g6mܠ�{����==�@�{�[,�Z��J���3{� �A�w�-��:VWn
��[�<��u�Ax��� �' t���mƀ����۪��ZwJΚ(5^�,��։T���;-f�Zž b}�[P�OxQ@;�����]�9�U@���{�
��zo<�O^p� �w������zW�@���:���,�kfJ�M���j�lm�  �Р����	]�n�y�\ 7��V 	�\z�ѪΧ�t=��QރCF�z8�qܦ�և�        j`�J�b`&ɉ�a4�Oh��)Q��d0L	�� �~&MJJ�� h    U?��J@4     �� �J��Q4b`@ɉ�M21J�mJD��4M� M������>_?��%�����~��������yw�J��2�N^��>�{޼�=3���w7~|��UQ_� *�"�*~`���?����+�C�O���G�/�?𨪊��]UW��UE~�|	S��
�+���_��='�e3	�L�fS09��0���&a3	�2!�L�ff�f0��̆a3	�L�0fC0��̦a3!��fC0��0���&d3!�L�fC2�32���&a3	��f0����&e3#��fC0��̆d�3)��fC0���&a3)��s!�L�fS2���&d3	�̳	��fS0��s)��s!��f0�̆ĕ`3$��s!�L�fC2��&d3	�&�f	�0��̆a3!��fs$�f0���d3!��fC2�0L�9�S0*fLʩ�@s($�f��s�aA�9�S0��TȆd �Ds"�eA���S0 �L��U3�`�"3 �d̂��S2�f�#�Q3 �dI�0�fȃ�s�e̠9�G2�0 f@�Q3
&a̀��S0�fQLʉ�3 �da@3 �a̠��W2��G0�ʉ�s �d�*��2��E\ȃ�VeA���0�f��@s*�`�2"f�#�Ds(�a�
9�2�G2��@\ȫ�Es
`A�9�\Ȍʃ�s
a̢9� � &dP�̂9�S2�fL���3
�e� 9�0�L(�̆`3���fC0�̆`3Ø�f2�2��&`s9�a3	��fC0���&a3,��L�f2��̦d3!�L�`&C0��&a3!�L�f4˘L�fC2��̦a3)��	2�̆a3	�L�f2�2�2��&`3!��f4˙�fC0���&a3!�L�ffS0�����O~��8�����G\�Ȃ��4�ۤJaÁZ�B%��'!!��p�Nw7����=����u;�%,�O��N�����F��J���79_
�;sFbC�}U�����gC{�ReƩ��
r�w\�'�T��irP)�(	�,뗨d��P+yHh��_FPv�0��-�rC�b���R�!�C�H��Ah���{�7*�!���4��s��FD!��*�˺֫c�����H�\�ih�{-�Y�j���]�n�9G`~�õ��խ ����S��pO�q��ٳ쇮��qv��k7+�؊쏧�wY��E��5ro�	vs+���|�ݍ�4w{ �;SG6$�Z�7끅جC9��<h����gh���.�:�RV�ӂ���2�U�Z�W�u�oe�N|�A�����q�����/7ы����B�P͡LVM�{�1�F�$V������,E$f�jv��7��ɨ��ܯd�膹\ł���ol�4�C�yO�:��W&��r;��R��8f�4��Ft���J�O�<��{{	<�����Ly"�U�0J���:��3�M����]�ާ�4V��'M;T��9ɰ��nqʴ}ʀ;b���`3�lJv(u\du�;�ʊx,Ҡ��)
u͍��"�����B��b'-Yt�CssA�i�B|�wB���s|�4�$��f�&7���W��}!�4�O���I�����̟
t��wh�p�FQrk��Wa��sU���/D
2$�X��Ywm�ZJ�J�s��8��%7���%2W��(c�6�ܵ�J�v��vHw�"Q� ƛ�Q�����ug��57���R#��)����.�0��Ѹ&�ub��� �@�1��h�TḤ����3e@�rf��d�E(�l���g�++������4�z�q�(Rw7rW���S���1���(�ɡ=��7:��]�#�hc4��t��`����ʑ�i(�}���͜;Yf���
b��1cCq�x��4X^�iمd}�����i�4�Z�<[9�x6�]�'���(�y�h��]MӺ�^S���+2�n��R+�7k��rYk��I�5m�����.V71G8�4kt�s^����Dr$y���FP-ίt��͎wd�N=�Θ3��Ʌ��I�f^	4��ܽ����n8��CEjg/I���c�8�la�g�|;l1�cdS�Z�*>����j<Fn�ׅ|�p��]�2=�s���n�ɶgl�-]�{焛W��xxeѼ1-��C���l�qH(#.ê
)6�ۮKq����ñ�K������Yl��ֶ��X�kJ}Y��ū�Ah慨�8���=�D�1*�No
:��ye���Z��3L�6I:IC�Ђ2AheL�Ͱ�	�ٲ5 �l�S�C����]\1�	;���j�YJ���6�+�"�6m�at*Y6t�Vp��U�n'�{:��mȠ\"�M������t�:�����t`�*�v��*�%�t�t�r�|\�1�<v�Խj���r����H2[+A5F�1;d�h��tis��vN[��ڏyCp3��ۏ1�2�[.��1��{�v�f��+�(�{UInI�gw0-�h���f��j&tw��\�)��}^g�n��ݐ�t�1aq!H f�-G,����nݽL9�ޛ6.�n�|dH�)i�x�e`[.��ɟ�Jƶ�M��*��ٺ�Q�4j%��]Bc:��gT$�����<'M�+�07����Z��"��ݛU�80c�+0�F��	����Z� 1�"�)dd+�1ӝ�
�|nq*�9��i�v��	�%-VAV:p�э�{��
��"�3)իчeL�B.no8�v��Ġ�1%2ӳC���
�RP�c32�e8��@���)�����xFu6������x����Ƴ
��!�$����{�_�%�����R��V<GAU4�x�7�D���:B��+4鱂����i�{�ZL�IV+�q�\�qk/�A���>���n4{�^ӦZ�ܗD���D'9��PNs��wT�_:NV'ǘ�v�K�:ƅ��Z�ؐ�Gj8�n��.�#$��������o�<�êv�����9�
{�Mӥ>�M]��!��Fzu,�0Kٸ	����1���P�l����'-�׃X}y�G��9�Z����Jȷ]`;T�x2E�l�pp=`��d2�����n�ݼ�H��i�y�ʺ��(����y렭ś��d;6n�8)���R�1��L�Z윂A��^�0��o[��"`H1���K����q������0eu��_,Th�Ƭ�Nq��w�bs!  ��ܪ�pUͷ���Mt�.��5�M�d�h�XÏ�`؇>ѓ-Љ�1RK{�Y��jY(�-=����_6qiI(�ͽz*�8VV��R��Z��9'8��:<X�}�r\��1Svęov,����6�Y�Y7�p۱1�!8��:�Ad,��;�d�`5c#5C��hoc< 2��P�W� �6��w�VptxY";����M����K��-�x�аW>�X&����e��G�͛�@�쵙ϤR��YۢC�q"���i,�OI�i
i������m�NK#�G^l��t\�XFn;�W1�}�p���m�����'t�/3+��S����T�G�FvH��za�'���h�N�u�y֍˱�9�.
��q�r"RKK(�Τr<�����v;��%S�N��-L�'6�\L�K�CZ͏vS޼�x�}�������m��'���
�M���-W6��d2C��z�T[��܃i�r�j���u��[�:'�5�'�,�Ƭ1\�vl�
7uj�ؠ��l\�6��*A����I�p�����I��Wl:��DָAAe!��ZV]�iu��n�,MK.��	/A�,(Z��sZj���!�B%4jO5�bd��;��e�YCyJ�n�=j�b���Bq�7/v����FSZ&2���Wq�!��;�1zDn�X;�с�fb�.�f�ralq̓���;��
��fN�kHiOi�5I���֕ܶ�!�P�Z5����
[�X��B}f�:[�gf�%�m5��29��}s�����{F�+�1�ͺow�sfDD�2��1��[X+�ti�V�f�%{& ^�9�v �ů
S� M�{Wl�e�f�;R�+!+fݑ�6�f(fMVM(�]��m
 .+@�{�iN�c�vT�roT~O;4�3"��{�a�%��5�n���9wC��%������ͬ�"8�5@!ȩ�Rr�����&�5g{gT�
ؠ�ɲ�tB�ѓ/��� �rF�E�%�����l/R�w;*���*�o!����Z�͙$�J�t�dFQ��5�q8�ٖ��q5��`�!ǣp�qu.z>�n8�vɺ��U�8r@H8QwY�#q2�m�S��X�v�,tR7D,穮�7����C�Ú&�.l���\��*�C����$rQ��ZSQ�x�9�L�VJ�tM�Gcs;U�ֱ�s����j��t�YЊ	WQ/䫋yż���u�FŖ�(��6 k(�Fb�s��Y��2�<a7�f��G�A����ï�v��`e$�n�H��m۫�j�-�V�	π;l$L�r��b���Dyn�h�`{̓��f�0���,�L���۝F��b.-ӑ�=���A ��1ȓ��+��t�y� gf���Nʥ�A�˚L;��E���_J8rp����뜑ng]��ZL�)0��tmQ��o�P=lh�x9�:�p�kkT�[�_��ۗj�0u*���K\vA9+w�d�A�P�`�谺z�	�7!�}9`S�]8��Յ��Kf��.;�
��{ysgjr��t{�8���ŕ��i�jG!Im��-�-��EVW��:Gט��ԑ���h`2b�p�xʏ.�V����*�j�IR��#خH���i��	&܁�p����X,��\!�Ko�� ����8%Ѱ*�K�"��yx�NĘ6��,kN���דb5��*b�T!��M;��#�B���9�;�6"�-v+��r\��]�؛����w"vÚ�A�X̫!�x��F��f���}Poyo��X�ZY7��.�<l�yw�+1��۬�X�9�:d�ɴ"�1κ�kif��K���4�ߍO{��(�ͅ��c�4���nZ��h�ǷX@QN�b�:�c�rD�nȮ9�_vk���ͬ�ז�QJ��
)�UXȱ��躁�4ޝ�)��sf��@dr��V�av�4��Ѻ
$�"ƮK| �{Zk7S��3�����:Ē爂�g��d�vS��AS�h^XY2��a�T�S�2L��X���ʍ]�a2�`/b��S�*i^MՒ�澙�K14�oa���D�Ԙ-;�<n�R�n����jjYfI���l�6ⱕr��2�hK9��ge�Љ��]��Fh�GJ��d��5�Lgw�����`S�ɬ���J�ѯdZ�UT�-������V�N��\��p��gw�j���1eÕ1�##��<�zF\O!� l�	z-���9n^��K$3�דs��s�s�%79��{��}��}��h�J�����:��n;�^!�o	ۣIc,3M[Egc8eƴ�a��ƫ���	ǯ4 |6��X��7��{)"=�� ���ω���
��Ɣ�k��R�r=F&���j����O:4���uUf<�p�^�����=�jrU��Pӹ�{_=b�����ݬt�n:�F��l4�\�KȌO(� �1%T&�ON�� ;k�u��dí5��H�CO
�`}��d���x��ps$F�ŀz����7qs�#{H�-3:%��r�7�sZ�7�z��M��*a�d�u�H�~<!:�������Ř^��:h=���H��b�n��E7B�4����a��ę�Jn�8�D(�2��j�T]!o��`�.�ɠ����sfk=.(�uYa�@��@��atù#"�k���]����e/9��L��KK�Yհ|��n�S�x��Ӡ-�����x�,Tӷulh�u���6�{@���Z�Aêj+����4`���Hd0�hMK/�]d����{A���r�Q:�������-��9�R�#�U�قlveM�C7d+"O���/�rʧ|���B>��wWfv��ѐ�U�n�J�]1��4�}��#y�p�j��k5��nWF�bh-���Hj�ª�5i;�w��wl?i*��P\�(��K���6Of;�tUcA�-]��2I�c92�+=�k4��k��$*7�gތ{�gh�h�̫����M�]�#�a>�ڪ���)�5�(�ʤ���=)��V��Ō�P���a���R��T��Vj�5���ې������"^��hڮ�ZG�ס.�p7���o>�3��e��^-����sv���<3�yƈ�V�ꜚzUb�8^��O���mV�T�M��P9��/J| �];�q�G(��fE��$��Հ���[�v=f��7Z���e?�����'��G�sXr&�Y3t��h�������,+y�1t��UqO����,�p�Gfn�Xd���?�.0����2%b��h���QM�E�0-�m�����t��M�t{oiR���]t7J�:�P��Bp�q��60��ӂaA����?b�4]���(PS��N �
�f��t�j�-]�d�(O��쎵�ܥ��B�%�Cs�z*ڙpV^۸&�Y��CPj��tdr�R�\�D+`ԨD�e����/k��skIrO	x��`��]�r�y�z�[v�RQ�#�]37v;�%n�.�%^���bJ�2xRGQ�Z��oQ��U�|��lk
�mi#3�l��h4_�qu�[�f��3Z�#�n�s���U�#[�2���L**MC�����`g@�n���D�a�ԚB�g@�ql������6nخD�w���:���ҥ�N��0p�zˮJ���AC��Q�ć;U%#�g!A����{�E����:�E�z�ᜰE��j7E�"b�î���wR��P��(V+S�a�,'7���#"	�f���?^锰r ���.�
�/n�n$`�u�VѝGBwq=�z��uK���s�7`�v�WQ�vK6�(�?��pJx[�0T�xX9:^�I�P�2�D�S�Ōa���c$A�J�	�Ⱡ㼹��ں�*췸Jv���[*LI�*�m �-Vi���t�v���p���a�����Hak"�
x��TH'Z-G��Y����\��֭����'w�~M"�~ٞ*��K��#'�D�Q��M��!��3�%S�".;,�q?���f��� 6�����YY��]]��:ϤX	$'T1 �E�0{'͍-1���6�s�G����N���y���:t�s���-�őx�4߮�T��R�F+���)�MJQ��㶭#��a��$�8�սU��x\&7�r��� ��8)	�ͦG����IX	�8��.�ĉ�%�RQ%�uyz��I�J�0i �rP�Ý"�W|�q�<t#t�c$�~ѳ�#�;<' H�ZX�\	ѠcCC@�!F}j�U�1�/���S��D�4� �%��+��čQy�L%��^��F��d��.�æ�����x�ff1�	(TTXoN��'z��),�x��]��0S�;�f�N&���)B3��v�(r`jIv��OF�Ք:��`uc�K�u;�E�B�	c8�wZ&>�{�Y����~{��V�~�?��җ��$�w�.ߢ#�~~}�ͱ*^�ЬF�I�d�7{r�h2��G+b&�%��	�R����AL�+�F��H�ȯ��
U����c�b��Vr�/���)����:a��X��9�/4�IbԦ\r�I����dC���<��W/0���wT�,�a!=�6�7�{��^�}��q��v3vj2��m���M
+�J��3��n�T1���0��Y��"$�3��|�o�Mܥ6q}е�p�V�f�ȀL���̔�NfK���K:y�M��
�e1�$5�����z�+�9�mejb��P�p�y�`�c�^��qEH�c�����AV#��&]Kz�&SR��B�����ts.Y�N��qs�'�;tM���W����.�0���uV����*�d�1ʂ!+T��i��`�������-�
�s�N	
5�Ү3ft�:�QO7��5V�qo�,��S�Gj{Î�n�ˌ��%t��i>��ʙ8V
>~��뛾�i�ŔqfP��d�l'�o_p�J��^؏}��o�w��ڸ"/��m�"3���B֥gF9�ĸL;On�!��;2��ٕ+�ҹ�k*-��@ۮb_4��]K�1�oy�0=܏,K@��w\����ͫX�U} xmu��in��zݳ�B6���vB��{}�m�l�ăg�����lPm)wec�j�c]`�K��1lb�v�t�S��ek1�$]uu�[�^'�V���VȻѧ�����{���z椩�����*�<5��`A��)�:�qMed�kq��V�s���۰\��ʘ�>����M�\�vYY�kF���aR�Y���ZP*H'b��y�W����:�WD`�{�ז�s94���WP�^=����J�ﮜg�vnqEg-����+�	$�Μ,4���%{���HdL�;��J,N���l�:o���M�0˗��L���)�I��Q~K��Ia[�K�$Ȉ��<g�}o=P���f!���򈰭���V��v�ӉK*��i�7B���Ü��
��9!rҰ�;�z wS뚶����t�hߗ���w�r0��e��]����v�ij���f��%Δa}�d�����2�7������ރ�&x�tU�W*�@���w��h�Y��n��Q��K0ԾD�ݝR�Kڢ�8W]Ff�t�p��4�B�y+�,\6ܥ��@��5e���$�C�Ī�wMRs��6[�_U;�0?r�Ϛ-}������E�X*�R�N�Xzscp��8pnI�|;��x�l�Iڱ!r�ɳ�\4 ��v\�2���xV��vQH�uػ�Ĩն�p�b�H}�#2��Vs�Y�E�E�mAw4׹@�e^���C��CO;�P籹5{KF"%�\���t�F�/2�sb�^5� ��p ���n��c��V���PY���"ܙ{ٮ;NLT����G�����ɅoUov��P��c�7E��wWdÒXqY��Ht�� �1*˕�J�6Ţ]vN���XG���!-������%C��^� ����g�+�������I�k��G��ْu_���w�\����2�y�z9ѣ���ƄMTխoc8�U������K%E�"�i�獕�J�]B�z�jE=1on��u�<�C#��E"� ���%)�>{�lc�>K��eY�@!w��M�� E�@�]�+y�Yo�Ԋ��s]�����L��!��0}��Mc�v�c��ꅭ����p�u���X"�1�����%e�o={�3��)i��֡���7��n~�e6^o#����|�C��GT�������_�6���p��`�\�1����t�h��3�qT��ާ�w=ԭ�)�l�>R�J�jX��V�[�т�|��T3��FN`�A�whS�Ĭ���qބ��o�k���.�;�|x��^ė��5����=㚎8��*��u���+��{��:�
�T����f���=װR[I<��������`��d�W�Z���<a0�w
~r���"}9M�O1E�2F��<�D�� ���%�V�.�G����\����s�u�eɿ��tY�Y\6ekPiNw����8zy���<��k��撈���ۢ@x��l�>+p�q�˂M�.��[^/������porߥ/\w��ì>�ͥ*�۝��b]��^�mԇ�֟ۛ���խ�>te�.�g��ҥ����"�t*Wfp�\m"5��*7m�9������0NKO��*8�]�f.f��sS���[�����-��y�@��x'���L�����]���bq���k4�!{'>:��T.�>�kpr>�A!miv
Qu&G��.��q�lrnQ[z��'v].�{(D��E�AZ����C�yW̫ۤs��o���,`����<'d���y�n�Qr��pl�r��O��Wn�ps�Ź.�`}��M��ww�N
XW/�ia�ڥ��B�
�b�����j;!�B��	e��DE��qI��b���ڐ���>���xq����$wh)AКtb�E�2ج̝t/�bŸ��wBS�x�1�����QF(9��I�1��8o��M�+����^ǆ�=��8iչgGf�5��V�I�c*��l�
�	�t�e���m��*��g$�J�9�m#������XNg&�$�� �R�O��Շ&_�s���BD}�'k��*�$_��x#�3�'�F����k˓f�c6�4���7�-�[�;+Z�-:̻�Md���\�}�@U6|<o�蟲����a]�3r>�g�M��3��d��M��y2c��I�k�4��:p�{R��M�V�d�y�kz��Dɋn^8>A74����xÔ���=8m~&{:Q�M���W�Œپ��-˺�M�|�9:���%B̖ )�e�/B�.q���iIP��J���ڮ�xC>wv�F�׻ۑ.�a�QԳ�+�7K^���f$%u�q �+�R�9i��XM�AnV���t
ErmU�B�e__
���lt;%3�����e��f�q��;�jl:RGV���\z��ѕY\��J�iw��cF$��z7ᄴ�j�/V���s��z��:l�o
�~�\]7N��,3:��9�3�;Q��Լ�D^iwϝ��.2��55��'Q�z_br���d�o�N^�sΓz��ws>+���9"!o&4��c}ٓ�EM��S�l�M�S4`��v�բ�/[��n��疞s�,3���K�܈ie صƶT���Mh���ޜ�0���f��L��4�QފQ��ve��Q���	}���q�P�&��t�w�y-�n�4J6xl�04;z�J�u��.'�h��X�w↓&���~��%=��,e��z7��[�����+0NΪ�����T����@ǄM�j���ds��2?w�5�h��&h�׽R��}|ᶊ.�t6��c� ����p"�ɌcW{�3q0m�\U���G/���b��,#��49���f���IOX}z���e@`�y���_LG}���܊{s�{�|R��Ȩy�����7��@��79��3�Уr�q�dZ��[}5(E��On��0s�l��b�P?k�|��n3�,o7��N��ǂQ�s�=����~���f�c��,$/N�;N���ss��p	�Κ+�sɹ&,�����b���p�M�����8uI���%1lӸyͼ�V��T3�n��X:��N9����5ݼ�:�9o9������;ICFm@���|��}W�G��z��q��:��O-ި�𮫊�t(��28p��ԩ+��I�RS`�����GE�i�]�D��]��4�:�h��q5��d������Ҳ9,��սJ��gݧ���j�R%� ��h����gt������ˣ�QzdJ���̬wI�s��n�}ƃˏ���:���A�s�"����"�h�5����.�we*lr�טP���G��v�G:m�%�N' u���c����_@�\�阴\u��c��G�433e-��9���p�@�q��識HJ��G�<B�������W�Rw_'�(ۯǄ x{A��au�V�;\^�2��u�2�>9(X�hgot8y�j��<�L)�4r�3R,Й�ONܧ���>. ����%g㙠'�ơ�z7_vW�e븡;锈3���rj.r'9�,nY�]6��(�c�e����p��˳�ì��Lc�L�a[���49Oy{Zr`���u�xr�`ۄN���=|n�f�/W=���C�!.�f�pp�'�ȿs�py�{7�j�gn��<��v�:w���ʑ��I��Ig:��Л��WF�ҠK+�I����f���;�xc�D*B�d��P�zn�����ɸ���wr��n9����ɼ��fg
�f~��Ou�:Ծ�5%���z2�tӂ`F���Y����+r���쑮���y	뒾1Q�8�镟��QIh轞ѩ�Eg���ޓ�N����'b�n1rw�#]��<��}k�mMn�et²{`/W83��A�F�5��w��vl��\�1ۦ�z�@g)vB@��qǫ��j�Պ�� ���3O�{hg~~oSL�{��n��������3[��[�ࡒ�fsC3R�|����������^q#��J��h�kJ�;��xR ���'�D�_٣��}&UoDb�8��f�!��m9$�1T3�k9:�z���އr�s=�k��}��
�[�l��j����>���L�2��8����a)��s��ɾ��v&+޺<=x_����waӒCLvҠ�nD9չX;bc	�ݻ�'�J��g\x�y@re��|	��ct��7Ԩ��9�O��x�E�.�S�J�̝SkzH_���Ѫ�Hz�@M#��|&����
�M��xDR}����w!Ci�ӗ�vx�8�l�t�]�J$ʹ��WW��:f��Qn��*<���s����LC</�>z�wŊzNG!&�rg~���t��G8dǹ���*��pU����E��*9(�qNěR������	Ll�W������(sP�p!a�'�x{�G��k5�b���xԨ�K9CK;�(b䇢��c�����>!�Ul[ޱgZG7Y�C
Xy�h��W>x�q�)7�4a��ىV�#^�6�Z�7�m.�����c��]���|g��P�D�8�tf��H�ʧ|��qN��,N�=rnK��O=!��-~����Vx�#�!^�ü3��J��<H�ӀB�U�n�E��zS�u������_J�PM���%
��ݺ��0J�폈Y��֫V��-��$���I�f�s��kW�#��]4��>���f_I������h£�j��Ҥ��\!�p-�L��G+:�Ng�*/��2���~��|/�L��I0�wټ׎M�gj揟+��Ra�����A���l�O�w�^���9�������^��:��qъ�漛;�kد�o�.�`Zƽ�����\��%#c�sh�]Ŏg{F�<�+�TW�(E�WfD�0��/2C�<];��'���2�Cs�-͈0ѭ�Lm< �=�OwېR��K���Jv;��^��U�Ӛ���;�L�'�1$�d��dZ^3��ޚ)�2V��%� �t�N���Z��-#�ӎ�'��>,���N���e��'���l;�xC�k8��=�����x�j�ѐ|Î�@oN�\�_H�jS� �$iZ
�k�0�N���"h��9��	%�M�������|��&uK��m�qf�a�[i�Aj[O��0x����?hS�T%�!?bA�gq8p,�����é�x��.�ɳ׎qY1� �H�a���^��R��M���Ś�33T"����w������ҚÎ`�
��q�5 /z�`�-�ui���Z�JHLB�Z֌��f`��M�a(I�Y���ͮ�|��nً�0�����T !;h�Mg:��홙9Ĺ��us2�Y���̄�B�֣���\�X;7X�5��u�o�,�vVZ�����F�[�{eZ�/xa��D���D)���Qt�ݪ��ޖd�N';,��^�^�l�{̓��N�_�d���UtB�YsWe�,�V�Ëj#D�w�[{�ҳDu����7��M�\<H3��z,uW�3�*/���U�ʘ1�yh�+9���5�Aw��Q��ڵz
��p{���f3��6��qg`��P����J��ǋ����
��y�k���Ue���7�=K-K�z��xQ�{�5FnT�U���&j�6���{�q��Ӂ��ɺ}� �-��r4�3�z=,o�ųL �b�;o8�u�3dY�I�h>�t�����7a�!�Q9�y*��t��Jj�4�C�P��mV�ʂ��0���L�A��֐�p��i�Gj�s�.=��/8ӆ�
�A�/d͛S��i3�u.�l�k8�bRf6�*#��&�J���T�
o�Օ(��A�jhC?f�x|3>Й�y�f5�y��ֆ.����wT<Z�3f���}��t�C��N��b�[i/�;آ�a�H6�C A���5��5�!�����f1���|~��g�gڵfm8Fg�>�&~�`���I���p@	�c9%����
^�|��R��,�,�)  �Z?��8�����(�!)��֛0R#x���U;?~�yhc-gۧ��AG�"�fi!'�	�%�k�;��U��p"����������*����?�b���¢'���������2��o��%�}���^����bߠıu뤮f�$7�G�>�n\��e�U������ٞr�f����<&Dz��2����bqխ]�m78U���y����	aY�'���{�Sr�K�H��=��w����gt�T��ХWt�֮ҜA+� �FC���x���؊1�M9��j�mMT��GYZ&�ыK�T�7e[ ���b��cGm�*Wno�CUPًc��7F�q��s�B��H��ŗjU��!-qx���۵*,d[��ʐ<|*��p��9V�E}��ծ���,���p۾rJ��O�A}��0I�����cwV����R�5^���u�_vh�����V�鬼}�*냔�nf���sv�f}Ki��ʕf#r��Y�^쭟V܋���5�w��m��u��f��2iL暕k#��Phe]^�!A�p'����+��١�x��4N�����
m��ܐ[��V{��Q�ܻ}�X>˜<t��:d�r�vs5v��tíd9��ZU�[��vc���q2���qE��V���:J^�]�3sz4��{��eo;R���\ݡ��ۈ�K'���`�S3�3/��a��f8a<�hk�礿e؟�
��<��=
�LS�-���s�!=}}�.xl���vm�����d�cg*��7؆�^�Bj���|�>����}�����{�}�������x��Ǐ<|x<x��Ǐ<x�x��Ǐ<~<x�<x������ǧ��<x�����~?�����Ǐ=�x��Ǐ��<{x��Ǐo<x�����<x��Ǐ��<x����ǎx���x����ǎx���Ǐo<zx��ǏO<x���Ǐ�<x�����}>ϧ��\�L�v�yT�2o;�+-^X5��޶��F�W� [Y�-WGb�c�t�A�繸vd�Ť>��1�n֖v��w�����х60u�޸	y�N
�4�ھ�gz@w���pQە��{�h�S��:�Ϙ�6����,�oٹy�ӂ�{�6<lT>�� Gq�2	=q�yn �{ܞ+�L���ۚ�9"�5���C�@�W����ΰ_p4�;qY�
+�D�C�Y]����&P"�"cn���=�NYW�4�O�rwgkJ�m����޺�ɒї֕vQ��J�Ռ�A~��4�Z2��أ�S�g�i�9��rb�H[�n��Ǧ9��9�'�QB�t�w��s�߬�ou7�wY��g{��8sG��'����mV����iìe�G1*޴�"u'����y��1r�4�P�������:��WF���XJ�;u�Iz��"&&ڥ��V����2��v�te��Ac�p�#��R6=�m���Ұ�]�d�t;��u��C�Z�gW Wg.��o7=���=ټ��/���Ǌ�Y�
rrY��$C�T��2��a�x��L��Ԑ��"�m��XY�����C��)����z]v,����J��P�Gjv?p���$�"Hr<�do��0�a���.b_�����ǫUs��������0��V.����0oc�����O������{�}������zx��ǏO<x���Ǐ�<x����Ǐ�<x����Ǐ��Ǐ<~<x�<x��������������Ǐ��<x��Ǐ<x��Ǐ3Ǐ<x����ǧ�<zx��Ǐo3Ǐ<x���ǌ��Ǐ<x��x��Ǐ<x����Ǐ<x����Ǐ>�d�sڟ�r�j����cz�ojh�>����<I�#�ޝ{ۊߴ�:P3���x@;�[J�F��0S�cnQ���odH3��|�b�x�I�S�Owa{�>UO��G��ޅ�
y��PJI�Mfp�n�v��X��BadXY[tZg��]:JeSD�*]��fmv��mδ%�1�4M*ӵ�iJ���ε(��0� �z�|��p��}����&Z�cE�����ֆ��������&+��O�:�n�;��0 1s�`�Nu�u7z�rc�HvxP���.�]�Y�9ZGp�P��r�����%5R�㓶
��t��[�;�U^�L����c�eʳVmi�\]ZB�\��j��#��
n�1+<�5�k���H���јZqfj�%[��]���k�)_X��`q�6���Y�|��Ш���*7 �>8&��Ղ�a����<��:�4��-B��9Ew|C�r��J��ű���L��ߒ����K�P�����˹��}Q3���C���Q������0�5VP86K���!�0pH~�ɝɇ�8�c�\K������h�����]�S��n`��'h ��0��;�`��cF��\���Evl�&E��S}�r��y����.����]�.��Y�7��B9��ٯ`�pf��8�m�WZ�b��=ބxl�{ΪBRZ���FZ����ŧK)n�ƀ�j�Yqe�n,�Z�ӎ��(_=1�(�C�s�Z5kMXa����2�=@��ڵ$=f!mD,��ͬ�y�i��.�;��	�_L�8u9t{f�^�g��+k+w����^"�ZW}��c�>1�$�,߁�^#/d�N��^�GYH���9Lr@x]���buJ�\�͏����o7����~��=�5O,b!`��70J���hQ8�w�-}}:��B�JR'�D�#��}�`Ҋм���Yˬ<�����u��Q�-lpѽ���Y|/�̋��K���Y'Vb�*gX�;y("u�0�;)>���_�?1Υ<��'Mݾ1��� ����>`s���k�s���ͱ��~��/�b���+�a�w3P�>�|�X3�W����ɨ!`��˔�z�j�9�=�ws�>���&��b�� �v��ۚ���M̕��N�&�;ˆ�]tx��5���ecBx����=��^P�����f�pr{8��7���S~�����y\���L��+��X����|�ѝFu�g�����ݠ��x�8���Y�/v�+��zl�neo"��Ի����!�}�,��c���@�o+j�Zt͕x9N�u:e%�R�0���us���t7k��8�������z;f�^Y�K�����ı�{�%����8;9:���l>���w�Y��qZE6�Q$i9¸����uN��o0�7	�7ʰ�ǽ�G��8Q�!;l+�x	���cW4#a6C�O^Y�Ҿ+.i��ؾ��Ub�lw�k��&��K�ҧ�f1#�TSHZ�Нnn1\�ڷ�����t��v�����m�&���^b>�>0P�J�8���y{� �|W���e�m�a��G`�osm����rQ�%�iX%���Tu�*�
�_���ظ_t͋�6j�ƍ�mv�v�N�v��1vK�
��R�"���whΙui���}E�rStd�F�n� M2����V�|ðFŗ,{�!f��鈲��K�5f�U�/H��S�� �e;��#ѦN�"1�ۯ��r��A��8�c.й��թ%�sX����j�b�XU~���O��
_&�M��J�zHu&��)�lD0nӪ��#Ï[b	)f'T�6��,�Ah�y;7 �eMv��fw���i6���ۆ�ӴT
;�I���tk���x�͉���1�k qR���i��Rز�0�\�L�x�Z~,o$r��Ꞟ�B��ܛN�9d���\//7ksD��M�J5<��+/�ɦ���g��3�����{`�5v��pZNԔr���ɱ�3/�R�Ո��ZA吺v#~��t���zG�����M2 `Lޱ�虘ثۗ�K
ؤ	�<��a�_o-��� \0.=�a.�4M������|e#
���X\�e�s+ti��dbU:c�PΛQ��_Z�M;���C/:yڮ:B�4(<����F��^#���{�a��{�ݩ���.Ȳ+�X�y��t��2{9=��c�I��t��Ls>�������acd��A+��E�%u�32/*X�o�^�V�"��o��7��\#��l4`ѷ�/���q�^<_��w}96��s9X���]��=����3�)�V-�[#�^.�Ƀ����D9�D�3�t(�婆ް�a^S����;�0`��kZ}�fvN�N��g���+�������|��&���ш>�{��@�3����[�9?r�3�[6w�!B\�Z(z�^�{��ֹ�$7Ow�Lפ�Cê>���|�=����,�����Ѣ)5>g�:�|�D`L!��l��������}�H�&O��s�Q�-�D����熜��{�̪�4�狆T��m	��q�/��ŧ�^�[-B	��F�6�̬ɯ��y-A��4־�[]9�c��*b�3�L7O)&iub}�ʾ׀n�W��ܾ����³���"�%�S�ef�!�����*AtG�0q��F��<��W��ˬ��<�u�,���T�k�Eb�	u[��e�S�騃�r�}�Kq��1X��'7����ڈ����
�[!�;�.��~=�OYОShJ��i��j���%�9�b��_@���g�y@%�1�ݽdr:����r�� �������D��YPc��	M��u�L��8CrXܻ�A�ld���n��HD�]A��o�S�E��]�E#>k��A�h[�[ܷo�	�O�F�2'��M�����p���S;�c��w%J�q�f�.1]X��76�N�.˜u'n��ژ e:"����|�W��l��v�wA����Z7�hOo۫��R����Y�L���t�^�1p�w���OC&'�I��I��o�)��쫫C��{�[]�gs:�Y��'����ZEdp��m�� �v��P�q�܇kȞ0�G#]'^���w�ŋk�����K��i>=�;�#ZF�ܭdm�LRE`��7&I�>}�pohΘ�D�~LC�w���eK��ۓH7��~��i�WH�;x =]b�ޜ�o���6r\�nv�sR��[��*��z�!-�?��߷>���^�҈���mI��I����H�|� 3]�q�.�����5����헖�3�E٤�9u'^%y
鲂U)��8��̡�l̂��p�m�uS�>��A�U���!�������V��6���1��\ѯy���f�J\�bB�	�H��ydr�3���C2���sN�<�	�-n��|n|n�ԯ�i�m�G�����<�J�|�*!Yx��9b�����>db�C[\Jxvh噯��K-ޙ���c�� �s�q����\׏���V�b�8�Z�ȁ�V��_0��#4��P@p�c7�@�UA6�����)�ڵq���0J�Y��r��IIȃ򽑝��/��u��+B� <riC\�*���^E���m䪍ޠZ��oC��D���\�-U��G�W�9F0�UK��� ������Mr˛Otͣ����X��ǧ�2��_�ꨜ���>Fb ��`	�x6>��7��o=sf�L$$����yj�Pþ�#eyv���V�p�U�R|�^�2v����F��uj�/� 8v�4;�[\�0t�����K�J*�=����Ո_e�zPɫhB-�q?�VdG5���8�v�=�<W#�s�F!CU���R�Jء2�;{i�Q�����H��gV:�i�ϗD���Y��!�������MM����U�����:����ç=���z:e7�}� s���@���y$��NUm^��ۘ�/��h���	�-E�Mz,�aw�b/�Xv��k㘆�E�Π��t��:� LM/����=�)�SXY���;Wgd:w�=�<���Y�o�l��O���J"� 6�ۍ��c�:�v��M�ﳧ��W�c���I٩1�9N�]�7 Q5�v��x��M��=���f@��;.8��F���^�r�&�%5j'6+��އ��,�:#��e�9��eq,��A����6�VQ��F"�z"�|n[��.��Y�o�q[^�f�\Xհϫ�f�G�6kr�r��i�����iдF%{�
�������^/7A��v:���N�s��U+7�4�.
����wX��zo}� �sz��!i:z�rD'�'���ݾ�ι�/��`Q�\ ��P�������Th2gg��ݽ5͒��fO{'����5nA�/�L�����Cti�ʡ�`��X�u
�p@
a���~x��cʙl�"ŝ��w�o�j��7�^�6s�u������UN�^�W�.��_)$��:��K·pG�xzmz�x�IW	��
��9+�3϶�mj�S��/�ҸfGg����v��9�dЮ6NN�������7a/h|�U:z�вo@�3�9q��*6���c�Ϻ�RձR���*��u�t�Iʛo�-O�������c3�����RUc����`��K���A$�/,ɶ�DC*)`���P�y$gw[�j����b�C�D�S*�vݭ�`gⷖ�'Ÿ3�ՠ�$�]���$��H'9 ���;)��7 :������m��\W{k ��lP��@�=���¶,�t�W!ӣK��4�*��٫�x�e��U���S�ˋL�	d,�����J�T:ڜD�O"	��u첑��ta)��lr0M�=�p�ɹ}��w��α��Z��e�ogF_M���t�Xƹ*��;t'*�FcZ*l&~8R��ޟ��౉�=1�^�p��^k�&v�u>-�<�h�fW�ةT�G���\�>�G͐�:�Z�pti���ݟN��<��c�Dł������������\^�����XM?�MИ�η�w�nN+�>�s�wh=�|2�7��3�i��v�C��{����0k�:��C�s/K	n���ZV�<���t^N�f�p�[���M��W�p�%'��B�g��x\��c��=L�^�{G36taPg[�t��sĔ��S��i�.-2��;)vL��
���;��Ò�v=�%;9YW�|�nػ&��F6U�w������K`>��:1��1.�3�����J�̎9괯{g�y���5�K�7��ctb}ÕY�.4�ڻ;r��S"n���B�T"��Dݧ��^���>������{��G��_���/��=����o�
_s�q�	��̃���@��	���!b�N��?�d6�5Q�\l⍈�,��<��n�!B�F�H�D�"�%d�V)���V!�d�E�!1(4�0�L�����^�rw^s٬�cԈ
�HY�%��u*T";6��ǅٌC�[��薳0�Ƅ��V���z�MBU���~�n{ր�'{���Yd�<qs�N�"L`��v�z>�HbśW��\�G����0�h���+�2p��W��Չ�~��T��ryn��';�l��x:;��d���B�SnȘ��K�a��ڂ� ��q����;{�k:+�ݓy	�o�=<���~
1�8��%�Y|x`���	�!Z�H-pRp����r�h'{��!�l����3ƍ���sԂ�n�d�Ek3e�}v�S�|�8s6v]IE�ݘ(���.�G�C}Q6\��ig���=|���>.���N;�$��M��N�R�]�̺�ך���F�[ۏo���Ky��ԫ�������&x�`��6�f���]6@�����i�P�VwFt2��8�Ib;r��Y2Jj�7f!����n�ݡ��FB�`c}�N��o���uq�
fL�X�nV�����±ԭr#�9���w�G�Z�gܝ�*a�j]n|Ye�R[��Y=��E���Rw��L������W�Y&yâT�M������p��$��ճ����h��%)�Z��pz�7ۻ��M��?>�ޜ����R
]O���&��4W]���N�<�a�#��oz�����d�``�I���R)��p4�$m�Ap�Lq%�C`���D�C.&�,IMR� Re Q8�GTt�'�e�e��L)6�Ft�!M�E6�h"�Kp�.XND`1�,0��Sfj L��%�ߠ@��q(��e�D,�$���-鶒1 �"8�m�q!'�!�	F(�!F�i��-�L\�В�C�[;��� ����s�bI(�u�蘩���ئ�L�P��}>�������~?<g��"�%��:c�v�APEH�R�"H&.��5F�D�V���&x�������~?���ǃ��EP�TSLsh������(n��Z'X���*��
~G]cg4�IU4��4�E1@EM5S�3QAED�l��h(j
("���������4�y�4wb(���h4��ij�l�)�����8�����*�*��b(`�*���z��j�����f��u��RT��c��ELAT�TVf��`��`�/[DRQD߃�]][b�(�m����Gx֦�E�b-�A;�A�Lk_Q�kDTĸ����c�Z:�c��m:��tQ��T�;X6v�UZ�N�ڰv7���è��V���6q��(�[m�c+��z�q��X6��1�4m�6�huZ#e#lh���E�dѱcZ��E��A�"����F�,F��jm�2kAS���q�Fv]k;11ڂ��F���=v|�h�"�
��B��A�>�'�K=����8�w�����yG#��
O�C�J�� c���d3���zb�j�;�z8Dw9��S��$)бU�
��)�T�J� 7��l��������ϗ�j�D�a�}���2j��[Eʚa�\��2F�����{�oF�yXo�=.���z����4�9^�x��1��7�z��\מs��;"Z��f\�)�J�Ϟ=��R3մ�V}G��!c"������{x�Ӭ{ >��r���f#}+bJy��z>66/*���Z���������$*�Z�.���Sm��H�V*Q�yJ�S>.��\����_�~wf(b�s��s6����{6�
��W[�>�<��ټoi)W7|"e�V�W��"���:ĸ��=���� cC={'�[�]��g�T*w��	馷�=�Y�nE����73�۪�<��AuԔM���5���f�M�`����E �/�C�𓶤~�S�nM��v��<>�=�*_J{^$�bϺ��S�){ w��<�����??\o�f?y،gi"�E5Z�����>�h�`��z���qaĽٱo.]7�2�g�s���D�BV�uy�������݇�wݡ��`U��$��k3�ڣ_j4�SU�f.]�xsKaNӶK+-VéI���yu%����		���*�p��A'@�){�j�|��K
�,.�Y^Xz�>+��u�����Ι�I���q��Q�i���tsY���W�:^���=�LY�Z�;B�03�t��| �<�I[%J� Ȩ�Ԇ���+�3>�t�YI�Gk<�b�Y��汯c>3�y��8+{`�����૯j���-�C�s�\�6{���ɨ�٬��H��t�6g�[H��/s]G4��Te�z��_��g�
qCzD<l�͓C&7x��c�z�xrYD�l����1r��v��S���~=o����87�+iy���Gr�xSx�&����Ή��r{x�ʹLbi��:���A5����,��~�5����p��ng�;5?/��CK�7ޞ$.{|G��b���R��E�g�Sgv���S�Tϊ�����A�O;�-y�����]Vk�<�Y�A��ͳ��M�r�\�Ё'`���K�F�=$����I��¤�im�����$�9ڤ�����ם�ؽ/��"w-k��xk�m�lh��S6\�I�bH���u��>��4_M)�<�{3×�ͽ��,oC�U�]c�K��`s7��{!�V��r��_��N��K
rs�A���~�GM�=��� ���j=w+E�_�����|E��G���kK�lf��]=���`M�x�Drѡc'ne��f#:-�W'E��� o���lv�7�x�qw��z�r�������o
����%��~�����>*/��t
�km	�v�E%cd�(���Y�����'�GQ��o��bW��^�>e;���y=n�{|���ke���޻�実9�~���V���S��!�\��V=~�oV�}C��C��~��V�J���dTf���;���<��J�>��]��	^�=ㇶr_ߋ��O�վ�m#�7^���q�vw+����Tמ=`�*�_�jv�y�p�#��F���:m�^n�O;���U����o��<�Y3��a���d�~�~4{�!�TAZ��ܟ�}��^	-���
��!䌹yE_>�&�i��õ��P�g��=rE�,��	��!���fz2zWQ�qt��g)�6�u��n�+��[qq�#G^�oj�s4�4(6�K����E�)2U�b'8uY��鍱�{;�j�:|�H����Wq/���F�O�ݟkP� 6�q�#�Lw/��d�����I8`��>*�v��7�
�7}o��A�:A9�@�V�{$�����g��n��L�Ox�m`��7�^O���C�x��^]���L*�Z=�$�cčy2	���u�W����b��\�����xh��p���]n{K��^}����|�}]���*��?8�=!z�׶��}^J���3�9�WOmU�`�-�{g�P(.���}̵�71�)0�W�L���b�Am�����������Z�|�z�>y�=��q.zi�s3�ۓ�']
_Ɠ�1�[(s�3�p�{h����-�r-{�=!?-�ȶ�ڷ��K;��jÂ����2H��_�u�υH�+�TE����kҳ��{�x��V�P��ƎY�(U25ǆ��\4S�ʭ܎��i:�1�[$3��K�:�1�쇕��iճ�T����/�Pf���
�19��hV˚Gm	?p�{"����H'I��ws9j[�!21]z���ZnW����!�o) �����͞�g\�����|�\�L�A���>tz�Y[L{߷�Ô�ۓ.{|������f~�.�J�{:,�3ߺ��4�s``�+�\�e垣t�IV':�n+2맴���D�;���������V�2�Ϯ�V���p���0������ϫy��o�A��llS�e�X�	�ؚ��4�b�W�ikٽ���mW����/�@+�:�݆�t��d��|fCL�T��B����>��9d��@��d���<��׶q����iVg�Ҭj�k��`ʁ����o�O��<�{�xN/$kx�; >S�<����y����[\
�E�p1Z8EoFlnfi�`̙7��]�E�t���R>�z{~�^� �_�p�����6�9����:^�N>�j�o}ѹ~�:���}<�!��9WJ�<<-�۵�y6�y��y{Օ�k�H�����EV+���\�uq��D�Ź��3�Co�����\%~�s��;
������;���+̎�P�E�������K.���T�Sx�l�����w4{$�zS�xz��r�"u�2�ByS�d�r[���g��y��m��z[�կ�T]|5�|�y"#�{J�z��-̞��&��\�����m׹̺x��L���A�SA�3`A�#QV�솬���9�������=��30dG�ji`�u_���J���e���(h�"��f6-��~𚸒�wZ�O��^^��O��|U�S�d�.|laqce�f�NHl��J��yV��v|�,�#'�\1l���9�VNf�g���=Y�N���i�WgI��)��c��I�[l�[lix�l��~��IR��H2*>cD�>�&2�{d�k�j���c���&�J�;� ���@��Y9�.+d�X�9�4wwpz-���?q��{E�}��R5�o�t�<*u��^�������p�~�V����-��P/+��;��E�	����e�s�%�V7I�lc+�B�lͬrL��¬?vv���ձ��N6�tW��t���|R7�����0��&0׷�O�s�3������Q���2�C���f�;4�'.�ը�z8tR�[u���R\Jm�J�/Zڒ6�N���	K�4��cZ��u�a�	3&�]8�b�����a�%eR����3Շƕ�DZ�{���w�bf�OU�>3�ޞf��leN��J��^���<�<Iι8��*��� s�����5O����̍gY®���}�-�sw��Vz�T+�_���ݞ&��I�������:6��-��<��%;���{��F=K�w���E����GH;�c��%��4�K�2�uZ<� �~�8ȟ�Ѝ�xi>�y�h^������G9�֊�}��vIe��ל�]n�o��'�˯8��^�z�d;���A�}�.�{n'���8kk�^���3�5w����~G8^��yv����O����]<s�ڿ/"��^�*[�l/��R@�/�r&r5�va���t:���0�?y˯	����.`��u�n~k�|��ߣ�ӳ-�P�3��}�t{|��Eح��j(�}`<�����L��=���+�"GK� �F��S����	�F)V���Y(�Ŝ�nkm��\�8uaB�n�^��Rܝ`�%�ҘF�K,�51F�tu��������%#�Rn�~����������������M��IS+� ﶠ�!��C^QT�z�=<K7�,R�(�����/7W���$n��h�����XeJ�cb~N���t����4{�[oc�<E���蚝��d��g�#^#��p��Ou���E2��t��"��}�o�ty�3���(�p��?}���I�K�R�~���̭���A6�C��֠z�@��;F��u���Ȍ�0[��_C���L�ۗ�"�����v��8dў�9W#f��Y���"z���˻�3|:�� ���F��X�[�#\�A�WF�d��� |M�e�w/W����~����D�g��f��vI6�x�y3�t�����#��u����qVZ<-���lV�A[Ŋ��kͻ�v��&��#���H�ow�	�0�-�{V����y�Jl0�Bլ�xd�y��-��T��u�E�;E�	��k�V-a�aTpA/���ۧ_Qxo,��{K���]�ٛ#�+-�v�:����0ol_n��wXI{��e��뙠�:h^A]'.O.X(�y8r�ϛ
Ko=�g����<;��R��<>���I>��QOz���`��Pz�>�=&�M���,�o�v��w>�I�{C������&n���~�i�J�>o����}3����~���;~�����z�j͜�%�7�z�>�N�*�I�[�:���=�v�?��t\�|�`�~��=�Gg�{%��㻧�֜�^��c�u�%��z�V�V����'���g--�t�-�ѥP�UEǃ�Ma7~��v��V���<���e�O7d��Uo��G����柬��e�l��bwrc���1�1�{�`���>$��=���p��v���^F3�'v�ރ>ȹ�Ouc�q7�ó ]�;|6I�p�����{c�PO��*Q��+�#3�h+�.��0�8�qz��9�uS�^�d�t�v�٭��s׉����������Փ-�'���3�A�<��9yh�%�d:�k.썼�*6���������Ot���j��e�[�]k�&Er��K�m���4aZ�d��s¼gG�e���}:�F���z$��K�=�oNb.���B���U2�5�m�v�+��k���J�ygB$`�~\t�û���.��z��[?�0n`�[��i�� �g<r(Sa=�x��U��2uչ��ء48�D4z�Q{Ԏz�R����|%��0�^��L�qw��=�l߫ޞ�E���HVT�����3FS�:��淳��٭�7� WI5�O���:���1�K�k���=����O�I=��z���Oa��4���x��5z[��X�ӧ���[S~�y\����>�oң5�=��M�8���|��k~����^a���%��S��L�^��]�?e]O���X�����<��+������T�'�������mH2i�7ͣX��q��T^��'I��1�:��N?{r�S���z���;`;�A��`��_S�ۋ���6,�P�K��w�,��=Q��ቱ�/Ӌ�l����W�${�4',8���"�;0���C��J2���*�O��$в��I9��]�5�$�=�&7'�_��Q�Ф�Y��U�k��������UV����Ū�@��\���8�r|)����<�V#E�����-j�n�lwZ�ku�Jue���
y�D���M�5���=�yv�_/<������?&��}���X��$�ȣ�+Nh�1����{��eu���6��{~Jx����y��IJ�ۦe^���mAS��V/��e=~�+>;��y��R2]8��N�M����x
��$l��:�s]\��͂��裏u�ν:��\F�5��z�5��Q�8t9�>��¶{�[&9+�S<q��	�t��28s��@�R*�;��i�j��k��²WWvq��E�l��&s�:P�H��@�ww��"������c��e ��ގnf�[�>�т�^�:I��X|e&��kɁ(	BM�u�	f��<c�Q���~��=<i�Z�p����Q�P�£�ʽ9"�k���{"L�9*�x`��Qt���$S��6;������ONpr;�$��w��ϳ�~�JFn�n��� ����W��G귫q�����܈3rm��+�0��5b�k��f�H��W�,vľ:����[���'}\��q�8���K�����Q�̳ظ�.y��:!�"�ư�9�_Q�YɎ�f��MEf��s��rR��Z+V�챣P��V�����X�>���̓��UAO@�u2����� ���ۡ�^y�6	`��U�Eo���r`:�M:�[��Ѩy)2�S���2�/;�U�;+ :��cp<�4�f	�5�F�kz��Ѣ��ƛ�y�(]욕��
x#��40�)�m��։����k���Y�᫺���R�`6��v2���W�"�T=�Ycm�6[�g�fmm<���N��:J&��5�{�Њ�9�K��B�O7����5�^t茋:�jf�܎��gV�Цe;�6���vWps�} �j
�ia8�Z��M���k��6�=� ���U.�W]F+	m�h	/E �@Y�{
k8��o�w�j������:����b���l]��crGoB*��B�1y���O�D��E����VvaKk.c�2<�9���G�����Җ�(�^FHvxO#�={�����gf�rHp=b_��F?[5��+����֒Z�)}�v�N���Β�xh��R��[	���4�wy��cf�Aɼ/��R_�-p[��<R�Jğ���#���9�aε���;8��ƭ).�N�+�H$b��
�ºԋ0��4�Y�F!���&�s�{�'�F���#�wv�JW�$�PC�vc� X���SW�`�k�7���n4a$q���V셛{D3�����b5m��N�X��M�V-Am�*a��ؘ�}[�Qlf���vLV���������~?�������?C��$TUG�Q�u��cF�1kD�}���{�N���H�-`���=>�O�������~?�����<�ܑV�F�*"��X��*���*��(�@�A����(���u�"("���	�0��"�����*��MM4��3�DE����1PQLACSIQ�0IG�$TQTBM1Z5UMLG�a���mh�(��
-���f���(f����%��b��(6�TG�uA��EALT�E0�Q0E|�UD�T�j�j �3DMCRUEX�U1Q5AQW�����|�^�N���hlB^��E�w4V���%h��w�{�%�G��G��4�z�W<��}����|>�d�^��8G��7�{NU���~����;��h$�0�1ý��*�d9\fm����&%�g��ou��+��,@�P��ᔝ����^�� %��,:��W�2a����y6�F&&{b!>
�Q�����Z�,W���	��e�����O���cW%L�ge���H����&�9�UX��|p�^�Z�J%6���(/	,$.��-��
�%{Q^��!�m�n����Wr^vJ�"rX���s�jj���@3�་M)/	�d�3?�sxT��L��n����b+�t�ț���n!�� S!��F%�{)�V�Roz�Dm�5XF4'�T�8����N���,�h��T�"���zۘ/D�/`ϠtD�I�?-�`�O�Fwt�yM��`*ie���0�r���9e��7Y�n%��26��7���_Iw�e'��NV�"�ʱO0��e����e�w(h��m�-yg���80��q���j�����yL4ڄ���-?,��:Vwg���H;���be�u�{r��c����#}�=j�`�Lx�>k�����ϵ�Shز\?π�������+��X�F4�K�0�����ځ�w�V�K�
ˣS���1�IO�d��8��WvNv�[۹�GX�,e��腛�_*�eL��˽�J[��&�m.iC��	V��*�Z;kLe�ˮ�!�6�s������5Rt;�1${yİ�!'��$3S$ct���1��u �śBg�u�zzE7��fO*���215���+�Y wUޙ�����;��7�,�e��d7�x�F�[%۱FOl��=�Eml�ݽ�;
�D>����,51� u);�m��ƫ���� ��-�6�9�{5;�4����ww���<��)�]���B6��R�ә�Šv�b����X�q3��km�Go���E��ǋ��R�v{�e6�D1�O�)D�m�2�X�0�	Y�s��v�}7:��?j
y}jZy[I�^[�-�2�]L�&���b�yxMF@xo���h���S����������\zU�Յ�6з|�xP����C)i=��z�(UŖb������/{nq��!�.p8@_B��梲Hj(͕o'�S	 -O�P�	��#G�a�Mk5���l9�߷��>�>�D�^m��	���0�z K(ְ@�[�^Qp�ߤ;G�P1-�Yp�jՅ�T����{aqm��y.�cY��S�v�4�e�?�)>�S�)L�<:K�4����Wh��:���0�7��nl�=�7f]G�AO�g�#v.0�*k��H1�{C�tI�H��7���r��չ#$J�c^}�m-E\��TG��P��7S7��mh����j�б�;�����{���O3&���&����f�'"�+s޸�O��<�-���|};�bN�̊m�U3vϣʡ"k����<��K.�k�nH'��GD&I�9�Nl�^�U$��gH�f��/'w:L����J��:�[��8�FYo����"؜���X�dtq���L[�fˣ�m��uVHk��!�.2�c��ǭP�Jc���qfD�e�h�4&</7��,o��:�{ ��k�Jn�3Q����yZfا`/�V��Ӭ����N��{�i�h9�<��f�w�kp��uN�֓"C��l���հ��UY��j��Ic^Gj�Sø�g|RTm�B�i�:*��_Y)2O\��U|G����B^S�ƅ�����/��F��|:�|3��R���(&�ہ�:�s�f��vU�kp��	�B�M"�ʦ�^���	��@Z�T��%G7���:A�˸��נ�1u�+*�x{M��^��%p�7��ႮZȞ���>b����yW�ȽnC���ETn�5tF,#G��Y�x 1�\kS�`�=?z��G�p�o�z݉�tU�6����T3L�d�{�걍1{��O��6�k3���0��8��Ç0w�?�?*"z���Ms;�]E�ܗ3P�Yf��Y͜p�uN}��*��ݭ|1��v�M�P�r1���te��SS6��U�	Q�WX=� +,+�o�2@�^"��lu ;��sW��l[7Q���۸LK��C�E�r9�^fh(���v�v�j�P���x��Zq�.���Ĉ��SZg<ć�TxXd@06 tE�����:����e�Gm����B�ZG�*;@p�^�w������H<5�Ŝ����My���@鋇 �覈��Zqҡ§�qdvp��i�F �2�ɼް��&a��˔��gaV�|$�*��W�mv&�+ g&�.���p���Jn'(���f��v��b~��t�C�5y��M���P�xR}
�j�|jRƩ�M���m#������׬z���H	(�`$��Wz݃p�9��
 �RZ���N���r[���6���}u3L�����2��J-]&�J��ËhN�|�0o&�_u�;At�Ч5U�c�����.g�� ^%�u��;�c��m8�2���-�F�:ޯC���K4?�K�K����z�*Çٷ���/]��Ns���[!i'�ڔ���"D���n�mj�WX�N�ai����
�>�ۼ�*���_K�cb}k*��%ߚ�^�<��K�!�_�R8{%��C{X��e�ng`g����wĘ�om!w�Q��Q��`����f�m��&���P��y��A�I�����#1m�{N���#	�_�Pg�-��+|�T�ft�L�*��u��r/��o7F�'`=R�Z�DA`L]�vFE�W+��Xs�Ó��G��n�:�"�Po*kbq�%�r�aj�����L�/�{Fh�2{ �)���
��cy��t<0�v�[+	�aD��p&��2��EvE��m��Z�!�^i�]WAiWR͵�!w0A�8s	��`w�&k��Nڈ�p$���dN�<��m��s'��u�̕N������F0��Ó�5�u���J5�a|Hs�'��y�z��4j�o[r!�֚�'OB�k~]r��{)?Yx�����C�W�LZ�� c=�A�<s�nj1��}(y�>�C���ü������qD1��Hq��MCI}��6"���V}��;Ǜ�3��N55��!�z��^=�ޡ�Y��.�5�Xi	]��}�՟��u﵉���������4��c+�7 >n.��e���R+/����%��;������;�w�����|Р�w�@���m1��9,2}\�u�DmEm�V$k��S6���׃�<���r472Xf��tk���Q*���ڢU$�9�*�b% Hv�#��V��ޮ��=9y��Z�_��qdĲN�@ȪG֛0l�y�"���@E+I���"�F���Y��n�F�毙4fB�z;8=��#�����=
��۝�R�^1�c�>�vr]�WZsf��o{b2D11E��3fq�Z�eN�+o�Č� l����Nf�s���3�_0�͝9{��T����\d�*8y���>oV$���,C�ٮ�p�s��H"}}+$ܸ���ܲ�����2@W-��4��n�0����P��ŵ;�#x���o.�	��Ͱ�2Å�;ެ0���E9w��.y�S���79���v�Y\�S;�>��S�.}>O��0�Ф�����u����y��8�cV�3��e��<�-�Y��q�ՒBv����룚����C����|u��l���b1�&=j����Y���Mk�t��8�x|�.�w�<X�¬���b�Gs�O��q���5Cp�㘧��e�6@wn�[7l˻G��K�u<������5(�B;��݌���va4�"j�(a�f����hP�&2�&sG�HI-�^�d�E�P�`9�è1�e�c�O�o?����<$z���d��t����6o��+�5�W�-7�T����u$�1�a��@��+���-x}yÝ�U��_�˨�L�y:=��C�1T�c���"�uaf��µ~�y{!�h��Q�������7����������e�����O)��2S�h�q�"&us�No6}��$M�1t����O�I��(��Y/��xS�/Vq����oqY����t%�J�&Ή�rҬz�*6�3��~ͦn_��a|P�zzJY�i }̌�����뫲�5�(�OXΩGz�SUqZ5��xx��!�v_W����	�z�Wr�:�����;if��Bɧi�������{� �n+�*�Ă�S�vt<F�;���N�=�F#��l��\J�<��m�q	P�85�ZOj�� ?�33w�Ε��bR�g��_��=B�[���\�[����粢���xS	+�℘	qAw#��l#By�ʻ�\ge�)ۜ<���ߘ(���%��B	��a���ƁF���c��<��h\d��P�c[THs�E6�W�r�{!a�Ш��C����M��;����(�:dN/*�����Z�d����Q��l�F��t<M�f{��䠳��ރ
EИI��<�2�SsPȄ�=��Js`�Z��"�Ok6'L��e��gN���=淒 �;/����y�}�B5�~����{��=ԩ2t�5C�`�f���g�`�m��و1��N"�f���lz��5�r e��=�e�.���O8��s�xd�xμM�|G��;-����6Ⱥ�������P±8AIa<s$t��G���̞�g[f͡ǻ!�k�1�'�[�%��SZâZ�1d��~�%� ��?�&�}�b ��&�U_'�o��/��e?e����.��K�uSƅ�s'��oF�{����aY�R����(>_���g_?f$���`uMY=�����<ʲ+cy�V�@Қ��%���������}�u,V@|��o�p�
��Pn�b��g��>��¬~ӓ�f���z�4F
u%t_)�Y	oU�X�n�޴���}_ϧ�///xGU���'����дې�� (Lj`kdޚ�̜q���{ �:�ϟ��`�{�Z������n���ဖp�/po�[aq�
�l �Oe��3���A�2�c=��pģ�G"nr�j�P�s�e�{R�ǜSy6�1���5ä��L��n#�I�ܻ+e�v�6r�=����94P�=�z��o29J<3]ظ�'cIZ�Zt���&��S�S�oK��~��):������Hz���Am;Ǿy�� ��
��J��0{C��'I�`�	X<���;��d��o;�����p��Kߦ���65���[ő�Z1`�"�W���-P��;L:�'C	\D�J�d]��h!�`%�dh=�KL�r���"����G�q�A�xZ�ֹ=Ƹ~��ő��4�?2��I��za0�_lS<�scH�0Y�?=}�����R���BlЌ��Zڟ/�6�#�?sճ���c1\̂��5axLf�Xh֓�6��a�NG����qa��δ�j勃�7QC��E���x�|�n;�ǼϽe��Z�M�@�I@"Oz�B6�0o[Tm*S��fÆk��x�{�䨙��U�s�����q�gq�d��M4N��*���	6���C2{&��%3�R<������:���2��wa�'V�2�К�'y��Twݸx�ܘ3�uoW!$��)}	Oz؂�DC��΍��xf�����?�����x6^vl������`����z|L�N�<2.�<S#I�>���{��U�Ky����/T�	t}Im����ۛ(z��l�\�2/D�7ҝ��(�#9۵wMb�!�kd-0�6�M:�9"��a�S}N��C�|��a�ZD!�&�4(��P��Ut=Z�O�~*��0�х���]�T�5=�y��	V ��{x��v��r��@|�F���%-�x
�1���(�s-�3L)72�e�E�m1�������������6S4+#$�o0Au�dƹ�����X�f�Ղ[j8��R@�=�b7�����}_?>���s�N���_�c���&���X���v뾵�N����E�v�c���Zx�}��}:�8�4��f%�v�W�"�5�a���n�%9�"0N�B�׻({-��K�s>���{)?N��ꁚY�\���'��i:vM�T1�-v��r�B��",m��, �#�.�~6����p�*�b������$�4���o'�)��V7/<p�2�Q��S_�ar�6�d�*|i�'7�sf�i�}%�RWA	m|�ܭ�iA�l���%�j���_aD�f<3��"C�r��C��/� ��;})1j���Le��-u�������:8��S����3�ex"ٳ��H��ݯ@���80�p��%򢐔'^�+�[�I�Y���8[I��޻T�>7��jޝ�;��W����z|��?��x
��������N�/���Q��1qi�a>��֎~0��T�?�zm����mz6YI��`k�������S�=T�F��PU�r�J%7G���P!�H]��_��>��>������e�.K����y�O���yV�)�A�LV���ΰ<�oL�U�-I?aOA��v>7��=�[�mgd!�a�:��VJ�j�qDĲ.{�g=�ЇO�k�gʡJL�v[�N9�WV�����d��؉�VFt�p���N{���:��q���/51"Q�����$`ꎮ��"��y:�{���	�3�p���N9#�N>�#z�$��)��yf�.AV��e��^���NF��<�/+�Zc�>�q��{8ו�oћ���E��r�&�,a-�#a���|�� �Aqy��bX{�[��dz���05��"�ڮoJ=���ڵ��m�ą^�v�-� ׺&���Y�˱w�~lcc��$_=(���7s�;'��B1�Un�Wѓ׻�ԅc�r)��j��t���#&�eG�����7h�а�<{�� ��Xzm�`�_�\+y
4��R����v,�+�1ցl�L��ìݚ��b���Y:l�)DK�P�M�z�ԊtQ���_H�{�0�.x�Z�.�_CK��ۻzȨ)6�6�R˫��b�wPs~v��2�Xw8��.c�L�CwuS3�)��F��=��bc��q��k����Օ�ø�l1iÂ�d�j�����{���q������eQ׀�<�vr@��w�֓]j�;�a�s9����G8T�^}�r�(�G�o
�e(q��f�f �f��W�T'o�e�1iN�T�C,���vWE�Vv_�H�w��<y���b-h�c͎���]*p�q� �xߦ�߽��IWc�i�TwZY}ƓB�'7>X��b��;�Nz�94��+��H��ڠ�4��b�=�|��0m��F89��Gn�@szm���0��ҫK��!�����Ϝ�{�*�1��	��zb&�8��t���Y+o�Į�ʎ�0r�Y���,��ܢ��	n�6�:ј�
�'8w(R�[�� ۧ���#�<h�>�Ә��:|@��T�
�}�d�Y�������H*�킃O�)�� H7�kf��0u���:�!��*�#��m/*�г�*c��+8w�(Z짔n��.g:=gF��p��C��2�A�h�/�+sz�7s
���3u��:�Gv@�ov�j�Վ��ͽ�Ǣ���M����.��/'6N�@6���`��q��!6�r^��C11�I�n�*��,ݏP��wbGӅ��9������{3��Q8u�_����h�s�WG�{��9y����AS�
0d|hE=-��5�}�YT���g�
���3x[iK�$����L.	4��o�
z����W��2uQ;��yv�^�8򄧪(s�{�����Q�-; h⫻8-�ݜ������f��U��y��)���U�U�B�,�ئ��EY��0yy_�A�.����N�n�<D��<vs���"��-z&�/]����t.��b�nJ͡��搶,��ʲ释������b;�J��h��|��K�}FI�!5u^���;u���x4���wGNz9���ہLЫ��h+������[�/�-e��o�7k�Ȼ��̗+-x	�ܼ��� ֊�{Ϸ��;Z��1	�{�p�k:MP���FR���5��|�/>:�R��)��V�㬢�`����E��Ǖ��]��f��ſN�9�!/O.�$�u����3S���	��S�xeq�:��v,���Ta�6d�% �{���繤�1��#���n���a:o}��닞avV�"3���-�X��e5�-��$���p�kw��{��q�3]���
#W����_-ՙ��x��� ��������T܆dL�UN'-�8�5��e����	�#&�M���A���j�ߐ!��*����b�/v*j��FM�툂�n񣽨""d�������~>>>>>>>>?����	��!�����"��8�)"f����*��5?_�o�������������~��9�:")��	HQ��ت�k�DS�cQ�1D�MR�$CUEUT��AT���PSsh�J"�h(�
B9:*���&"
"J�(���{�@���""�h�"��fOP說���$�''���/[ATU4M������PQF�M,AD�����4PUw�DDAU{���ЄET�D5�	�%-RPU%SM^��1QL]X�$��b
�������BP4��AM%Q>��QCCQ���_���$!1�"2� �<����cA̕;���f�A��-���%�͟g'L�	����s���.�v�n7�S��oh��@����p�2K,��7W�
	�U$0�(�Cn�]�w]积����s�"�X�FuYI������7␧�Y�42ˎ��A�u�dye(��橾q=�k�5Y�Vv?��>ק���^��ut�B�pi���*h��%p��p�-5����{/L���q)=y�Nf���sA1\ѳ���SL-�ֽ|&xA-�ļ��RQO���ޡ��2�[Nu[�jz�f�3X�e��/xil�C�s�=��E��aG*��b�:\E��`EE'W1m���g�mP:��T��E�A�=�hJAm$�J)�m���֮��o�,�`�-DH
Zj/t6�vWZ2��eU�ܢ��q+��֓��q@� pǻ������U���a%rq��H�Vd�)~��;��Z-"U�����ب����EchF����'+ K(ֳ��Re�2ۥ;X���>�dc,�<	�
�\fLJv�Ӭ��as׺!Z輧Ej�IL��/F4�1ͺ��VK^'�<&Ys����nq0�b/6���n8lc7�>Z��ZD���f=�����f���k�#5	V�FJ�݃��ưQ�K-�-��^oȾ{��K.��]	�6L�Uc��ͽ�ѽa�1��YQPe
���yV)��z_%������Xw^Ɲt]�XƷ���z�֓΍��.qc�u�t�k{��Fh�ͶOp��-[oo�^`�=��n�����#@�4�&�����}U_ϧ¾��?�   Oe�L�A��Z����s|�^fN������O,n@� �cL9��O�h&D��ţ��wp���J��P�� T��`r�d]axҷ�F����A.+��Ax`�!�~��Ֆ��6̖[�W�(�n�B^m�oH���ŦyR����/6
�Ƒچz�G�!��c���=� ��J{�'��;�,91�z󮣌�:�N8�Uk���Ҭ����o͇�h4KnM,펉�|�ԁz���BÅ�kq��Sz�:���`�J�)�ze|'�n���%�(l�g12`?�%��^(6�<1I�
�lbz�n4�1Xt��R.�URsSs�ׁ9~�o+.��^z� ���Y��m�5����H(���3\��	�d�W�F5C	&���ElilCq;6�k
ė�v�zfa��D[�VkF�JN8C������&�Fp-yݠ����OO�T&+6]�[�<�t�C�PiD�4��-�tM�1�Ҕ�4�#`m�w9}ѝ�4�J�Eļ0ݭO�T�Fev��FSh���p�v�/�Z�q���a�uȃ�DȊ晘��n�3J<����{��d���82s���0O������L���kI�OPXD��8v��Ŷ�d�&��a��:��n�y��i�J	�8��l�dX����I��b�E��NVC�ݲ�9!�}Q=N�łq�q͠���^�n�����	��u����?�\�~��9��D�sE�j1��*���r����Z�K;T�����C��|A^4�����|�/A�L�q�1�����n"g�$v+'��z�#��K�e�WM�`І.��9��lxs����+������mz�h��r!����,�D&T9�S��2���ށ3槚Qy��O�iZL!%�����X��a�d��4�����8Yb�S��):��,�ƕ�kYj�U`��^��W.ڣU��{W�5�U��ĺTFR��������i�.'5q�t��cڜ�$Tu9j��0����;��Gq���-�����!�6�W�n��B�����W���z�S	�����K�#q��F�z��T��sإ���-�>-~^� ��
���g�͐X�nD���ñ�b�Lbk��jTl%To��O<)����䶐å�Y��p���%�7��ֲ<���ה�z �=c��QԱ���f�,aY��{]J�^�H�l;.��(!e��=�<Y�6�pȽ�đ�$�Z��t�L�&����[�@eK;�.��0H�)�ٚ�͔��g)���ԏ���X��KW�����h�}}�/��� �>�6 �D�0S����<�]{Al�����]Y�ȅֶ���+Q��y4(��fI�rKR���F���a��[��RVI���|��� ����+��QW���~?�[�	�5�)���n,�/S������rv�����`���l}��OMQٯW[2:)"سS��X#<&�uf���c4�ˁ��>#l(:lL�2:��������59�[�Vwd6�w���i��mj�n���ㅘ*�^d�1�B����j���S,�V�Z�;��S�K�e<-����@r�)��'�6(�����&m����߶�|�X7��x���l�����8��'�y��S��7�6?�2	�g�#)͉���ׅ�c^�T���5��&�{�3b҃*Xޜ`Z�9A�6g������І ������/Q�1LMR����X^U�(BlЌ�ɩa�[��hXh��1x�oV�m���:آ2h�d=ʤ����"!�a�d)�ވA?�x��@�R��Y�j�]�u�5�t�ג&]$�^�r�[^����0k�|g�M@v�:p@"�����>�Nlj�Li#I��m���=u.{��;�*b��t�\�ʫ�~!��a�������_B���	�i'.�,2瘘�s�ѷ�]����y��s-��l	�gZ�1��c������F�1��߃>���{&U���p�=�Ohe�@������S���-� �.ҏz{�ａ�-��g*s�Wf\\:l�눚e��c+1d��vҥ�#Qp�4kc$�ڦI����>c�������r(�Q�oJn ���T�&,�soa��:�Sy[������ �7�l��o�5mϹ�ڜ���慉7<KՂ�9�t�^�I��qyK����z����7ܬ�-�OZ�;.�W����~�؂1]�����/�R5�= Tw?He�k:E�5Cp�����3(߮UWEu\��ve5���P�)�z;�L���,3]���c����*�$Mձnn�S�H!�c��q��;$u�ҝ��ܡѵO齁=+_H�Z�R��Eϟc���A ���z��*�n;XRM�:͕[9#���,-)�4{��ި�}�/�Dn�RU �Nf�P��;m;�D[曞�YM\E��nsf�+=�BC
)�Y �hr�A���˰�����8��&6�'�Q�j�CN��4�%���hA������C`�1�A������̠ӭ~*jo����SO���l޻C}�G]�yڼT� �36�֞�<����N���B2���&ʙ�\[�>�m�DO#���\٫�M�������A�7�쪶���a%r��o4����i���}��C'R\� ~��!��oI�$j��xgF����	���e�\�L�Z�iYQ�/)1N�s�*,EÂ�:%��YF��V�s�5�G��{�%��`���Y&C�rj�A�.'y�wO��d���k�i������p��0o�x�����x��ǽ����^�.evB�������nB9/6˜��� ���Ɗ5e@�*��M�Iٚ;5���'��^=�'��l%�3�ψ��{<i�b��2״b��Z�RL�T�lݜ��#:�5���r �CI�P��IL�w��Ĳ�헲��|p�������9rI��Q�ڲ��{t�{���d����a=�%���Ƶ{��=b-��j�RW�<��E�P�;;w����̋8LV�G�j݌q������LC��p��\;�	�w�V�ΫXڻbu�z�=(]�Ƅ�8W-�0���l���x��-�qq��+y&\��Ⱦ~����渖��B�"�9]D�w�i0��+���iy����������(�g0��F�($7��S���`�D@M��^u�q�E�qG�Uk���ҭaH(�pb�S�t>Ea�]���A7�
�됬�v�v��y��=+_i�~��OZ�tZ5��tfe�����Q/����A�4�`�\�W00���v'���H��/
�e�t�i8DZ>�@�r��R�w�(}^l��b�ޭ��i�r~^��Nњ�r�tڧ�Z����^Q|.P�F��{޽���T���t0�Dt��m�ѡ��ӗoZ��qtʏeNǛ�om�}E�f�IA}3-j�B<=WȞ�u�ꪯ����  ^^^�� ;�֣�'y��3���KŮċM�j�o	����?�G�o�0��oج�@��U�ݓ����۽,���K7��me&��ő�Q����Ϭ=�$�V'I�`�>tȶu���������N^"�;>���,c�ay�� ��T�L�tM�1����x�@�%͖�2d	�/�ڄ5��)ᦔ��k/4ۡ9���>�K  ��4��\�S?Q�|}X�#�L��U��
j����A�U<R���c'��{�}�)�n�٩m'�ķ��f&�p��l��<de��^<��Ϫ�!�P���.4h2�l�buϞ�u{"�KwQt�=M\�;�>e�� ��9��Wtm���z�^��S�d�5�� ����Ay]m��QD�fE�Wtu����:�Є˼ħ6
�Ì}���U��ܠ�X!&`D�݃��,o6��)��j`^oD'�ʽ;� $��"�x�4F��^�C�L[é]���b���;��Gqh�tO�n#11�r00n��ԧ��3����5��Q�n֎@��UY�����x���'kΘ�7���xu,"I�4F��胃��#
��`�[==�����蕛4�|��˞�d+9d[Z�oxl]�m-L)Z�Қ.<7�r�w;����	5m�T���n$�yT���Ľ݁a��+��K�Jc?$�����s�PH��ϟ���V�K��~@�`���lMm� L�|dI9:�L
9J�����Ҵ�94��6��m%�rr����|e�5I��+��.6]�5��;>����4��r��R��hT
��E�<�i�k�>����;>P�g�� Ãa�b�w��Ķ)�ݥ|�"����[v��B1V����{*	{��J9��3nt[��Wa1����s��>�W{6v/��q�ʳ�dN�qo's���!T�����Xon�� ���	|���w�YyB��Wr9^�P�Y[���>��_�?���-���H:"���g�w]�E�������F�n�|�zB���A���:�����W�$(qWD4�A!���-�se��w�%�b�=�į>�C.�g)�����KM6y���j3^�{Mi���f9��Tԕ�Q�V�v����>�"x	���=���'j_ʿr���T)��?��ǔ���A���Z�>�p)�xH�2��|\�l^����$r��l�|�=[��%�"<������U3�R��5��/o��[�n�r�X}
1��Df�\i�Y�k�W����7�A�oH(�XϽ�*@wmF�31�u���'�]o*�rd�����bZ��h��4����7�6������V%t��,׶�8��Co����'-�\��ڨ�u�_����N� ?O��o>��{�����������E���&m^$��FϾ7rÍ���H�Jc�Ī�&��S�ѯdG�iD��ڠJ���ccu	��%�����٣��%��̍���$!Y*�����N(Ƚ��4���W�k�FEi��m��-C�2{�U�U.��K'�qL)��g�MG���y��C����;3��U��	1)m�kɮ�.�ׁ`PP�D�]Z��2{�t�M(>c����q��n�&����+�u	�ԃ�F�j+�OT7=30��������3�d۩fp��:*���:�/+��Cp������G����<�����*s��ڮ�]7}�����^���y<�^�\^O��3l%f���M�^/M��qWR��D�wO�63��妙g;�yfEk���<�β���Qʒ�Αa�U��peាӏٹԡ���P6��M]����;[^�]P��M�wU��BU��0��y�J}
�FVŻ�~�5��\�7�^b.�I�h�@���i�v$O.�]���Ȥ�,cYc�otzs��2�/���1�[��'��@��4s΁�x���h�ef�C��r���p+#���^���x��7�4fș�%�O��[y��k�����G�����fy?G���zv�;�G����p����ll,Q���{&g8 @T��uY.r��;}��f�_�6���-S��n��b5g-i�1��r��/h�6�m�	Hc��F) �E���yX��xg�^^�������s��i��Y��{�[�:l/! ���aE�m.��Kg�t
��V�	�n�s�����]ښ�̺��,�g9:_u��q�7�IF'����n1�+
eܸKu��+�-ӄ�U��!Kirr<�/�M�<�TS ��L�M����y��]�(\<�0&cyQ�8-�J��gm�vќ
� �Ľ�\�����Z���p�Kh7��{*[��B
�֝
�R���J�# \���|Ǧr	���e�B}na���(�3�Ur���i8˝��x�\�Q��K*��(׸k
����M���2˭ZZ㠌Ru�ǖ]�R�lم�t!�s4C�w�3���eQT5�0���ȸ�rp<����&��K<��bpO6����#�f��n��Mk�$�ZS)8���`�)��@ǣ�7|�cκh=�2a�ʎ���a��eF��_Re���|��Jp4%Ɓ�8]�)�ۄ{h4�`�¤��~�	&��VyS̂z��YU�چ�}RS��d]g���q׉�Ƕ�1BXV+�ر��U���N8�h~�2�ȍdg�T�C~�sG=|�k�QwRA0�:�
�siVq��%��I��s�·P��A��2�1����	u�ݧ�!~So����̕���c��u�֩��Y�"��Ҕ��2'�TG[�\�޽�^�X�5��Ĝ���vJ��.����wk6���	5B����tr:U���U8�n��s\��홷C��He���25-���@��F��)J]{o)�[Q�6�k�='�x��[eC���Aǧ�֗*.��I/K���eJ�0t��9�S�������B����������ˋP�>!�lƶFW=n���щ��N�܏1�	�Uq�0Sx����M_m�Ṿ��n��S˲w��*��Q3!�9�}����Nj��Fxְ��#���Kx]`z��I�1'Dh]ԥ����	�E�1,��P�
�nD�ͷ�a9����N���9ݔ��$�͋��G���2��Em�
��*!�3�W���l2\)���;a�<��-���2�r�����P��/���یn:�، �_vi�MJ
�/��C�[N�*�fv�9P7y2�u�|�d5ڧ��/��X���P3-�iگ{|�6Oj�K�OF�=��5���u�т+�6nIgxiCP�a�����[�jh��岧k�p��i�������<YAH�$*$Y��X�{�ȱ{&:�Vڼ�f�u���u{�pgP����;'j���V�L><{j�vj��~We�bE�wL䈮T��p�6�:���-�=�`����}��'�0|�]�?ѧ��\o���0
in���gv�ѳ�
3����\*��l�kgs�	[Y���'���7��X��E�	���K(�#,�ե٭�4D��)�e�ce�Քd�E�Y���:�0�=Q�G�h���G�8w/�Cj�O{9�^�놔bN|���5xh��{���:�)�:��YW�wݶ�/�����.����ݹV$@s(�0��)�<���3h��C0�q~�ȗ���ol �1���u�ӁWl��3/���;�,js���7��^���93�b�s���BUd���8���!���f������^e>Р���g��R���W�zH}ۓwV��8A�B���Ev�ڻ��s]��k(c��Nn ^�^�'��x�R��n�⒱�e;$bU�˧f�=�1!�a�0��:�vӕ]��<�����	7{�8�X�*[{$�<n�(�;}9z0�/����cB�73������X,�+�چ�'z*<7�֢0j�<1g?�앤�{q������P��8��E��l�� �p��wzN�y��C�۶>�5JXFf_o���W�7���:���fB�}qT�J��)
�G���*+p3X�XC�o8�`��C�g���=B��sQ�1u�3ے��"���h��1b<I�t�P��1M�#TQ@��O�����x�||||||||x�~�&�
� �亢����^��b*!"o2i9>��nz{}��<|~?_������j����Z��������ii
�"j��i#ͦ$��(�))��� �l���CE4$E1%%Pz-R4�AM4�����:�PS�444QJ�T�4�^�Z����������))j�ګ�SEAi4�TK�tMIEMQ������������F!����.����=B�����CԤMUQM �i��d���QU0�-4z�yuDI��@bh�CG�UUE��Q%RS�{R�h)�������4u;gUBM�[;gTPPW�&ty.gb�{�PWښffک�҂�,��[ӣ�S3jk��W5ݽ,�-�P�,*m��(5�̭�������芞��ʋ��PS��~��_}�~_��g����y�A�=	yM��ƅ�I�P�+��j��Ib��0얫٭�uyb����]!�����,<�!i�fsT:}uSƅ�d㋱�*�
���g���[[*n2UV������:��0���J �� �pU�Xa�0z<�y�Y�Á̝pd35M�7q-uPnfߓl��ν]X۪L�o�Mx��g8`$`�,�C���l/��_-��'�:�?
k���k�}���FRb�]di��;�f�-:3a���	զ[�,���5fYf�ȠК��4�ͮS;+���v'�tV���Tq3Y�G�Y�5݋톓�1����:>Q-r�$L�H�졙{#�vX���[/A�}"�/"��wH$=G�fZ ����n)v�J$���{��{���c�ă��p�Oܤ��Rf���-М��e��܇,�jf���9���>s�̆�R�]���4Ai!w ��2�$k<+3�3m�!s����e�7+e�	圤5�̡Fɣ����H���:��hB4^����bu��Y��vpO\٧�(��k�os8�ĝY���E،�1[v�dx��aa^~�;���8�l�|�TM�7e��O>��`�Lmt��j�8� p�	���mEu&J��ʍfʽMN��A3�K�9,����=W^sνw�~j���8@3��we&S����~ �D��	���r�ѷwiX�y���k(̒5��N'_�(���~��'������Fl�� /O��%2,��R�&�)*��'}��+�������D���-ӟB�����h�W{ԯB�C������v�7�Ru��K"� �c^H�`���F�x�)���o�fҍ~lh٭z �\�%�n�|$J����E�S�\�QL��ň0yi�4���cr;��a��6�;4���M��Y��q�����I}�'��]Tqy찈��wjh|�7��[q��}e��d�m��� �ψw.6]�6����H�Wu���vI��͆�z�{�Ў���ùKUz�1s�8�X:�a}P�a��
��b�k��wa�"�mFΝ��M����Tr���ekߒ�^��R�i7Rͼ����81x%����r����#b�G��dv�NS��l��V:�9���f����9;ZAGh�qCo��EwF>�ӗ���L؝��
�Hty[������~Ւ�����.3Z=6çG;s�{��Ь��"n� �.�Cc���'�N��S����h�q���no�8(���v�v�����_Q11�ҷ�r��4ɯP���A�y�gLg��ZO�J`Q+�Bk�2�+�v�a�3��������'��g-�s��Ͼ�}�������� x\��O��N�7G�A�z�@^����A������;99Ĝ��DЫ�@�����W�﷠]*�/d�z�5/�bd�Y���ߩC��/��Yd؀����)��Ck��6�e'�@u�g�p,��g���R57�'{� ���=p0�
�}���ג��r���T)�|a�>�ooC�����T�lJ}Ο߄��}�>_�q�Y�JTͶvPcB��ԑ�^�z�E�7V8���g	��m��ke,��������&��hU�
������Q�1b�N��0��{�%�=c�v��츐o3;j�Z5!��� |�,.bA�l7%W5�A8%�~)M2�J�Z�������՘%g\jz{d-I\������'�MD��GM�q����,[�~M�RnX���4�w'D����Gf;�Ԇf�kg�y7����u@ky�K�c�p�p'����C��cc���I�1�u���]�f�WՉ�lWF8dn5j���$G�po7���p���#�7w���e]��,��s%�i�ia7C׹E�����Ժ`����I �k2=�Ýp�1����佂���}��d ����F�_�9�Z}Q�'�	s�7�N�ci�%�ߓBߦ�����7��9����E�F�_KN�⧃�c�_�X��禁I-��M���Y%Íٚ�m�o�,F'H�|�9sQ��|���
��6�����y��y�� < �ҋi5V�X�C�"��M1�g*�{�1�E���#���f(�!�5�"��"t�t��M�y��D��S�8��ɡ2'�W��SuGu[]�oIO�~��y�K=^W07Z�
�O���3�vԶ��y2&�؂���5����26�T:6�o\GZ��0j�V�J5���Wad�j�}���C{��N��ly��Ƈ�?���<��t���K��j}��)C�!���v�:�(mv�F8!i�R�)�6Z�6��ԶC���x`��WM�vtD�����7Pr�]�%}V��2�Z}�>h{B�..��lg��\��}�_���d�Ƚ�qݸ�y�L[*sc6}]#{��QLC$L�H�ִ��6�h�@mx?T�ib��&w�%�ߋ]K�c� �ܞ��Ϻ��8Ҳ(,����IE�z6m����0%&]��n��-����B8 �v�ya`D܄o�QX�A	����'+ K�����ٙq���"-�X���+��U�O��,��8E��s
�@���T�g�e�gLS�b��2�Zj�S<S��5۹9�7F*�|��}�IY؛�5��)u�+SO��m�}i��
��2OP�[���xr�N�B���uє\6,�"�-�`���Wg����)3P�`�(�L��}ᷓ�=����n@�RqT9[2�4`�����f������z���x �?��{�����8�F���4(�U@&z��z]v���p�� ��"��v��V9:)�,E�ָ����˾�筚�OnbS�)P�aU$��FͰ�zhYӍ�cD:A��w[��PP�θ=��1W��CO�T�H�I�����I�� ���5�<�Jb郿N�b1��&����V

YC�/�&����Aۨi��)���E�x�i�.iv'��Y��^&z9��&&��$��+O{Bi�p=�^�_��ƅ'ԘQ���Z�E�ʓr7��Ԙ�z��t���l(`�vJ|_#��JTo�M�fsTOk��`Y��N8�������v�L�q���uB��Վ�Q�GZ�Vr�����{���mnl�	�Ll� ^���;۪�y"%T]$�|��Ю�>Z��۠)2��Fۆ��y�3��+�)�'p���"�P~ڳ�������hr9uDa��� ǊS�Ƚ@����5H+_�HpRl�8L����d��j�ެ�w�6j���-�V��fIa�bK׸÷c׸����\#Q�l�|�&�6yd���1Tr䵵{(%�A%;r�s���`�7�Xs,'�nU���h�b�{<��ő�5�)�T�exv�"�ӡ{�}3��8-�T�$ɞ�^|2z�f������{}��خ���������5�M����8��� "�c�j�����9��ϔj|��ӳ�f�F��w�Wt�C9Nm��&X�&�k�/|���s���	���hi�Sw+(u��Y�P�?E����/�oؽ��;T�M�d^&=�(vNǋ�-��ǵ�Yl{
oPm"A�BCL�jgT_,
�sG:�#!jbr-F�Y�ۧ��@��!�Z�o��:����m�71P��3�Bli�	��#����9���*�wit�I�:fa���%6�2%�D��Gh]���Ɣ��Vg�P���qۭ���=�ḭ	�H�{^!��ss�	�3�~EJ`����]�M�׵���E��^n^k0���/�C�cG���������^�7�Ru�/Ⱥ�x� �e0�mNb����])��6za[.ܳ���M;6�ءփ�8?N>�br|󫈡���t�ZoP4��S�~����ў��kd-0�O䠰��M���a�}�+��7�JS��Rkp�Uj����-׼2�6�E(�Wx�ӱ���A�a�
�����<�ِ�NC���6Ӧ%�g���T��B꜈3΂]�S�x�k����H�QZ�VkYN�:�ac�J���G��l�2�nr����r;���>�=g5���D��#u1Yǫ*q��k��`�tvǛef��	7OS��Ag[G�Y����)�&o@�2���y�<�8��<�u�m�2�Tٴ���&'u�ڱ���=,`[�.ܡw�Q�y������Q���AFSpk#$0��?K�l��8&'M��,ٻ2���P��kcpMcz?���{���d�s�A�N;!|l�W��j��*�6���ס\������r�+I��1L�/z9O�^�q��10�p8�����e����&�������j���-����RV�i���4�oڲ}��%�@��*雥���;���#�ہ���	�gI���0��PM�:�����D�!d\EO�s��.�z��g+�Nחz��4@��b��J���i��K��M�=ʼ�%F�S-|�]v���m���u?l�gϗ�Y���4wk� �i���m9M!���ˋG)�"�%���Yu�3����͋���l��C�f�=(2�����Pz�i���o
�E;�u�� �5�2�wJ��BY`s�1q�4���W���!6#1d X���Tg{�,�͟F�jc�]��L�^�hU/xS��P�WV�B��X\��`�o��n��bY���)Uօ�+����fN	X��{=�n�S�m<}˚����CpF�GpEVF�gw�[�1�M��fA%�
�F�7Aλ%u�C��O{=���G!#؂�[��q�^T��Λj���h�E�KT$�*	�;�-Fjuqd �o�4�G-AU�V�kNn�16W=�
��=���<�8�˒-s�qe}��o��++��i0 ���9�9_��������<��	�vȺZ"�E�Ք��x+r���u[�9�;d���eC.�o �XIv�rn���9q��w��j��ʻ�m�}�L8C.���ሤ�g��5���a`n4ꀩ���I8po0Z�/���^˩�ښ�MV`�R�b�l�Q{�]��&�z�(���'�Kח���i����F�~�Z����9:ͼ4���,�>B<��ri�xX�^���7cy�O8����b�r��?��#%���ª�EN��S;0;̹�C�~5�:ꁢⅱ�&���ۥ]'-�o�m��~�~�|�g���\����_v�
�'�p攉�� �8C�plԉ�ژ�S�)2Xuy�k,v�}>_<�-�y�[m�7�FǾ]���{^��a�5�Տ�X@L�5���ʦ��^K.'��,�m{�h�r�qkf��;8��A|���$�
49iL�V�����v�̈��[�k��ք��\r�S�>GG�	��懧�yqt��`�?��5���H����驹o$���y�#9N��+m�r�����W27�}6uge�X�ʚ;_Za.��u�ݢb�;�$7o�� �������z"3iN�b-�d^<�S�`gx��b���=�JN�dae��/#�c��<�^p���������i�J��&4��1m��y����	��'����A�1�{a֞���d��W�#7��(�w^# I���������fִ���KZ
�A���!���x�zt���٥�b�k�T�\gǐ^��r1D�QN���s�q�>�h�ظr��0�|��� ���LN�g�H��wqeG�_iY���]Xg���T�g�)3nv�Ӭ�!�=Q=�$R���v�׳�"˯��ͅ��+
�0�����CK.�j)�������v�F,�vTõ���ً�V��I���r[���I��NyA�Uׅ�2���ٶ�Ы�� ϧ��(Ͷ��a��,Y�:���e�Y���bt��E��lq�(q޲�� ��8]�)ᆸ.����EⷳZWp��#�cOK@��0/' Km�P�����q�e�E�sv�i����	��չ@�W`VB�k�ұ:
Kv�à��R���\hU�L*�.xjU��=A,�{�
�u-��go;pWG�3�S)D7 ��ø㼠Sϔ'�,`ۊ��
�v?Td���7'k1�a��J?��>���ԕ��_�z�XLpG��	����{����mΛ=G�Y��~5��?��~��"EI��H�ԙ�sd�l�#�yw�-�v��tR��n,/{wK�B{���E0(�������Į�+%�kt�)|��{��<����ꌮs�]u`�DU���C��³�ShPЬ��0�a��Y5�"$Wth91�uw��osҟ%c�~Oҵ����Q��p�R�@���+E���Z��Ј�<:br*�&r�A��s�;N�a`VG�6���Ĳ�v�2/Y�����@r���%��,��b�Kb��Tsn��?ޠ�C^w�O ;����mD}tg�|����r�γ���4���A����H鈽��%:r�p���5bp��Q	Ԟ۫�DҜOY�7E��y����jN�-��A��X�V7V71�����$��5�V1�>
��o�ew&u2�ͪ6&�t'*d9���οz��5|�6eg8��u]�����N����=:�����Y�܃��L�jhTg�xoBx��;�дA��E���B�n�k�DL�W�R
����l�AL87g��!��sѐ͉i�܂jz��2�@����*��[�����h���eb�Фg���y'�oR���CY��^-{=���V�V���Y�2��!���� ��9��	O�V�'6T����J�Z#f�׀`�e��^�B`.|[v_ߊ��jY�]�H]�ܘQ��?Z�E0�L�S�:!�QC5�Bt����Y���]��B��k��g����-�KT2�Wv^�JaNXtke^K�\��v<爤r�B�5}�m�uY���z�\�H��z�:��w��S{��� ��׵!Fiy5��{&���)����1�m�]e��纫�{}�>���$3hӣ�⃽����ǣϖ��6��^�ۙɅ��nm��;wQ������6q9r4���_\�JJ�j|����̽µ>���+�Wg�
[h,|��K��s����{L�9�ՠ��*1�f�]�#{�ͽ�̀�ؒf|,�nn,�ֈ.Z�'��i������{�ξ�;����hVgc�t��V����kS�1Ȑ9B;)$���o#d�jf�ixm�!Yȥ�
g	���hK���8ɕ��]��.]فf�i����pc�����%>�Fj4��'ޏ��W̚N��T�v��V�S�L�C�fi��'�Ug۳.�ms˳p��:̓���E�+��K{u.�,�g=�=���:��Y�Դ� I/'9p�s4�d�a�jsp�n�y����A��^�ڇj>޳�r��od��H.���N�b�H�FZ"Xo�V]<�;��	�h�e�ɉm��n��m֡w�B�o,k�}��h�k_iO?T
���s�.wXY#���Y��~���I��{c�ǘ�o$��8����rx)�6[�,@ol���hα�7�L�������9���B�3r��9[ڨ�hy;it ���!����t�Gp5 �k5eҴ�d,�r�x;�l�w�ag�^�j15�+P���B�*TY���+X
��B�˘Yǃ��J���R����.�(�V=˺y��'x�`Z1W�Ѝ�\��PF!�ގ�"�kQ[�͡^�D�4׽�ua��ၷ�OZ�ن���C]e�T�{Z�>ݓe��G�fJ��qm����O
�/����˓y�s��	K1��&Q�d�8ڥƄhX�X�U�S�l�"�3e�B�K+�oё�S�t���6W�&�W��`���`��]�㸃R�wVN��b��Z��"�bmic�F���;QT����鍉{[Plz�+�Æ�Ǻ��:Od���*'�}��a�v����&�gx����Q�$��u�WEE6["�T)>�jmq�Љ�6�6����6Ntv�Ð�[��E\mQ������&�\f��:���1����Ս�F�U�hK�d[˖�+�	�!�*�=Իr(.�4m�]Ҳ��Yِ�kD̊r�q�A��^�x9ۻ�b	�U� s=���J�yN�Q���a�2A�ږ�A��t2�[�
v,�1�BJޙ[��۳�F��Wo]oNͱ��h�.�`ľD��F <9�3bϧ�� }��SAEi�!JP1EH��OooO������||||||~�_�}���!Ӫ*�H����UP��R��j���"B��O����Ǐ��������������H�H���Z=�b~l��C^@�
-�Э ��˥"
iiS��
h�����*���!;��V���E@D	4w�R�X��(��(
]�Zhk��A��B��*���)�h�hi�����Z(
)��l��
(���]i
%�4�B��h��&����(���� �LBD�EQJPSA@��LJU%	CQERSD]�ݡ��������
Q�&�!/�$"cy��W��r�y,�9=� ��h]�w�RM�!��"لӰc�YيIHlqEp=���d�ԍ1e����A�B�j։`�I
?�N����Ez6�޵��]]~h}L�
t�:��_�'���kv%;�m����I8amC���B`��8#/�z@ޙI�g=��bh;-������{CJn�i��fKu��SN�L�Z�f�@�&��P�n�!e�y��Qt��k�F��섿'Zs�{�~(o�0�?/B.xM� 6�%�bh�l� ;8�7}D9�iȈ+��Iz��FZ 5��^9a�Xsm����&�l�!��B�e�kv4Ҝ�C�(�M�y��M���Yr
h�֭++��rTa��w9��w=*a��B	�� ÃY\b��6oTS��MS*̬T#|A�Rɍ�Sჼ۱DF�?kز�I/��)A�:ʆm�b�>T�H����C��v�77�8e �x!rvG�I�S謟A=-�w��M������4L$ϱ<�x�x�z_Y�4�bAG_X�8s��8��j�G��ӄjm�Vg�7�Rv��6�M9�}]QC�ݻ<&xM�<\m�s�2C#��.H�
����~y�.��t��+�ݿ-gB����<�.�H{D�I�.5X����C,�L�7�6�<;��l6y���|�>��}i��ZW�a|�����6��J"��f8��j�x�i#��ɞJ{�k�@����9}����M�e�Ӎ审�'���fso�k*ĵ��]�(fbp#gm�r���#�+gm$��ɍ���ΝL�q�{�;��q�htn����)N9?yul��f��,4�K,!iJ�"�o�z�1X���)���×��m�h�=�w�W��e�ߦ�Ҟ�F6�⩛l��Ql�!�͛N�cb��W�k�S�������u�S@���F?�`UZ�+��W�y	M���Ɉu�6�=��ΰ�#z˫�R[z�(�|e@c�_��e��!�2@:&�c���l�(d���'	�d_3��T^��b؃�����3�k�F)+S��52��]t�� 5zc�)��}'�<�lx=Cr|׳ڢ3f�j����6"yȿjoH�)MM��8cʚYto0�$����;`=�C�f����d.�g��xa�X�É����?-���6���9�ƝP����-$@!�ջ"d!����W����ZҦc1{]�{
�i�	�?���	����r�@~�h�7h�Um��6Gi�#Zˆ\5dǭ5�9��gE����M<�β��ي9RC41GP�*�9ܹ���gӦ5K�o�;�à}>`�D;)�q��ŗ��"��������C�o3���e�zx}��\�;W);ER��^讵����/:.�3f�?l���9�1������<yU�7�؇���ݼ��(\���Au��ELfa[3�!Q`5x^¯3Z���[�L���X�:�Bn���E� ;�D�J���[���g~}��y�*���ɭo/mD�8�זǱ�+B��/�y;#k�C�����-d���|W׌�&��)n�E�����n|:i���H�[P�������t�+7��ʷ�]���u02%��D��:����K�+Nf�W���\D�7��
Zt�HO�1Ma���9�<��j�Q�x����������|B`& �͠����P=���k��uc!�j���6Ÿt�5o%�]���q71�3/!��hsCV2�����l�W�>���@wI�j�Sl�W�37��kO�}�[�!ۗ�J�,�������$�k��V���r�z2j����pB�p8c��A�J�H�p�R�9������*�ԡ2Bl\��zeZ)��C��k1Q�=�Y��?�G��:��I�������0�����# 9��z+U�ʖv[��ØK�C>�P��/��x�'yi��q5Q�Zj��_���I�@p
l�Z�w4j��P�j�0�[Qf�o���U���"z:� �<�LՁL6JvW�D�-.�_K1��M�]�'b��)P�aU$��b�u�z�Wt�{�K��V.+�]��WY��=\�-W�!H��U7s0���H��ݺ]Ky�[�?��5���z�8+�~\�Opɣw�O����hpG���c�+.��wP`��֞s�s�AO��_fG������U���ҕ��K��m]�Υ�m(�=����<���*Ĕ�C�$C�c V�2>��v�oR��x	��y^�.6)�,�M���qq:h oz5u�0@��!��'�pG?{����P��<�h=�{S:���Xb�tO�9�|�u�{��P��8AI`4!֝����П�	�B��&B̮xi�vh<�=���b��]�ؤ7�6�;P�Sø��T��ې��a�5C�����'c�2��J�a��6$���K�C��aB{��E��³�ց
�x����ۮ�/��9�І6�\�)�V8�/ҵ��A/mr��H;Bu�ðy�2�l�'j�Z�C�ԭ����(
`ұ�6��0̲E�՜�l���¡�t�����,�j�fܥ�4B���Ƈ�~��x��_�Lp�pm��� �:�3e�V��Ê�OEC�c��e����m�d�幦�O���l*��J=�X;�Z�2~TBu'����D^E��wH$:�T�;�s#f2���[�@~����P�-3����bO�N����΢T�E��^�δ�C­���:�V��ĺI�h�'ΔвT+����vQ�Y5;m�MQ۫��墊*��S7��5a7�zl=:�j�Z������]�9��\hF��n�<E��z�y����++��,�x�B��
9ƫ�>�|(|>ա��[��~��2\gD
,Q;����C��Y!
��[�l鋇U�g�`���$���h�W��AƨuN�v�����<�������B =��A���'AU���x�C�v������l�R��a`�A���Ȯ�rģ�t%ė�|b�mT�3q�6QqA2Zf��iȫ=B����cռ4D.���V�qFH/�1S&D(��Ϙ&BE�x���<��Be�/��R�&����{d��9����f��S��Z@��[K-1q
s��\�(b�
Y�J/#��5l"7V�^���o�u��s�ʜ�����;��}�XS�W8�)�nQj�yƱ4�ب:�q����.��e�������p������jOy�&��U�=[!i���L̍���I-�&n�Is��2+Wm���wV�e{:�8�ʮ��Qi���,WA����:M��[���8!q��F5V�ީ@\>�GUgXP܄ħU�=%�j�r���� #������.�0�t��yY�- �a�]����G��A�^^p乡1-�6KS"b�2LC7Z��9F�{���n��Q9������U�H�����繀�i|�.ҽ��a�y<�0V����f���ɸ:Ðs�������u�3�t���}z�Ź�}6�*��])�0�ʅ��bh<��*9K%{���"�Lj|�Q7.,�]�o׽�]�������>�}��J�����6HW�!�� ��5;?�Z���O�'�����n����i�w�h٥é���VNs�T99�
;�5�aa�ݭ��j���p|�<�����4������م��4b/xZ��.P��֏>�h:`���y��.H�
�g�Lb�v>�Ac,����� �U�F��7Pr�]�n.H~D	3F��^�-�dg)�6<)i��ѕ��Q,%E<�Z��'qKv�����hkN]d�'H��#���N&�yF'���9L�Բ��h�U�,�����\#)�Lz9�^�4�rT���#e5jq�j��3f����ݻ�͌S�FO���1�c^���[U����U�)7X[(2j��4�m�h:�WL�S-Ӄ�����TJlQ*������v>���[ ��U���' ��y����h��b�Qi�C7��ߕ*Mw���1I\��R�XQ��}D�.#�ӁƇ��+�n����F]dD��| CD�3W�@����`�����Yt{�0�_���t�y{�s����%�0�u4�C�w���ϺN������;f^ۭ��R��5�`G�P��g-�I��&����1Cn��b'9X��N�D��;H����5"$y�&Ir���n�T��B�Z�}mn�'dCkmc�X��,�����cֹ��m�5	�1BvY���+=0 o:���1���Ftacۍ:�/+�ZH��;�2���y�	�'��ay � �צ81�{<ԟ
�n�	��g����zL���L8��e(52[�+Y�o���a���KYp�F ��׌�'9��ֿjc���:�=�ى�mL��Ȩ~���ի5f3��$yiDW���h��͇���%�ݚj�oJO�=]��ұ�5�HA[���I�)���iH�qlA^���p9�k�14����=��Z�bb\�3y��;�كY��[q�.�WA��+�r�dF\[l+B㦃+5��Lj6�OvӲ���x�|~˹�:�pm>���\{5��V	[k�	t�0J1φ�.�+z�v닺Ȑ�'��[�q����}>����C��v�Ŵ>hA���;U��eϖԾ$���Դ��CA
H���ߦ�6�+n[�59�q������bf-��aJoI�� t�^�;2�Ⱦ�-	���!&9����2���xo>X��=k�!�_�ָ|'_WM���ox]s�71r�w2�ê�3Zf��$G]<�6o<�qfM�2G�/,W�/]f��ˡ�gϿ~l�ŬP��	ޓ�j����l��`*i�
r�˱x���TP�����;	}tЖÄn�S'Wvۍ�;v�����o7��� �f��_l�>k����S�$�y���$s!:c�u�·�쥯���]�O�5���Jy����A~�;c��K KY��[�Pʋ�5p� �\؉.2�'���كK*��ܢ��]Ѭ.L�c��� �c�hŧV�B��U&Զ������g�[���Wk������L���0K���"E��殈L��xNx�*�2�I�>�0˦��Yy`�������d���ַ9�a��e�Hޅ)�����(�.̀����Gb�y�u� MBe�*T����9�	��y��H�6'CO��O,��v�Y�����f7�����'�m��R��q��A6��t�"�У~�I�B�+���]��&���a,�y�i�T5b�o2���ٰ�?&H7��Rt�7Í�bڹ�P�ۉ��j�N������+]��QaB{��GE��<�|P��o@����0��pPu��ER�ڽڻ2)kt8,P��l2q�ҵ�%�Ts_��ؔx�]�����z�{�����wAo�}��k3�A�[��=7.�a���ey˾��{���x/5t����{���cJ@��ʨJ�2w�Ga��������ˬ�EPؘ$�I���CY8�V�Fj.D�v�|k $��Gp�����o�h��l��G
͒	�e��2fY� �����.-��6�]c�r���C�Gx���0[��"z_�Q�i�� ��6�\E�5-�G`Y{)߱��bݖ�ى�'f��W�����7x6�3T���Or3H3���" �g� f�9I�߸���4tNGw;�.Δ�M�e����0Ѭ­O�O�H���x�j�~=�f�.���nRb�oo�w
͉����ٌx��fhvt����	_<�
��g�iI��[�eM�C��-ٝ�{r8��8���d�!A^iK�v�VX���#��������6`���1�����v���&�j[r���:P�����͊aP�tlS?Sn�}��L�
ۄ���tH��+<��q������D��FBeAa�
Kс�p���KC=���5:Y/�S՜�P��S;!�bذ��]���]>!�ʞj�B��(���R�&��Ȗy0�eNH�d��~X�Β�>��SyP�eyAJ�p8���!�O��@"o�zw�Ru�v�j^z+f���c٨�۬ئ䌦����v��i>beٸ��6ա�C����mػ���z��LW),~Mv\��73S�k���zv�er_	�;*�b;{;�Ļ}k���?H��oJsۿ��~��ә7ӛ��7��̔t��sǽ.�a|��S5���#�ūe�9*ͩCNͷ˩�50��7t��c�E��؊�o7���=�����
Ȯ~a�aHs�2�]^@�J�	i��Ñ �q����1�AJ��Ul�X���)_mq6T�?'���,9~��vo6� ��`��C{A�g	Uc��y.��GS�b�`Su1�`吇����j�q�|U{O�c�����.��;ClgmTN�}�/�� ���g5��CfD�9J׿�ʌ��l<C���v���K��ƒ��;����NG�Z���N"���78���b&�q4v\���J�W]��.K�P
2���c&�;+5�<T�n���w�4����Dt���1-C+" ��vb�+�x_Qx���Xh8rF@��p8D
���@uHu8�7v�6i����Y��2_x,��F����D9!��MCN����tE�x�_��T�$}��s��E�S�o��(��[��JvE�0S�Kǳ���J� �q��i�sͼ4�_s���:�j���15��8��ᡨ�}��������y�ױ�4�rT�@� �^*q�jxO�n{=����s{�I�p��u���s��j�.�l[���������2�K��ۙP��yk/2���S����.����#�<���4�;fNZ�vUn�D�ݨ������h�V��VV�"v�Y�C��Jӛq4����Q
���MZP:�K~#&^�t0Y{�n����x�p7�kޝXW���'8
V��u��ǴLk{����A}Ƴ]� n[�Y�;�Ӡ5ؤ�N&x_x/[X;��]Ĺ�=�\�ݗ��[�9�����z�h�,3D�-���=~��'��:�>��<��dI�(���:ê���G7�1�ھ�/h����}���5z��Ǧ)}���q���F�[Wc���J�ɔ�9��q�_k�Rs�;n_iF��@�P~7�Y�:�v%;-�4���+k����A�V�V߼~�}�<;�x�rF��<�G�ڃ�E腾#��i\D^����aQ����#W]8�$��2�ni.e�4Q�ۥig�K������D�Ak�P6,���у*J�dM�&f��n����60a��U>'�sjhs	rf����v>x���YF���I�$�dr���H���Ānv�՝wd~=��j\��/�B'�^S�{�~f3�2�,{�V-�vV��޽ �(�^��m�U����o�K&�!<.�<=4��S�;<�!��ٲk����Ԯ��:wl�[X����<aq��b�3l��i�h�`w��6�tHޯ`���NJ�Kc)����<�/��0ɫ�����Co�����I�d1!����ƩV]Җ-�+N�^TQ;T%5��hη��Nա����]�5�'�F.Q����vA���+���w{7�����/���j����oMzB��w�r�vB��w*V�\5i<����7C���0Ɣ3(k��N��E)�hft�k/ҕ��*��(h),�Ehն97%�6����Xf�s�����	V�Q��=�[���+��R��w��um��rq�Je�v-k����}�	kTm[��}tЎ�_eٮ����e��(��ڡ�J7�F�
������*f:'N�=��ˊ�R�J��u��-n�����g�Ƿ6Z��)�6�B�ͼ�ؠ}�Su�7��@+���e��6����p�ƌi��j>a���|r#�gc@�7�<wܽ����k��Ճ�is���!�ܫsG�F�S�=0�a�g�g���.NxS��7���;^rn�6�>�I@Wr�Re�UʜB��o[�Φ�mL�%畳5_
�߯�t��b�'�K�,?_k��+ǅG{ӣC�'73����q��������3�����R��r|�n�1�d5c�I��3Ck7�3pqע�E�Y�l0�+3LXP����L���Yj�Jb)��+n�{P�'~�PD�dh)JW����)�	�� ����}�^>>><|||||~�_����!�)CKT��V� �Z�"��������Ǐ>>>?_�����D�-JP�KHU!M��!�Ί )�m�Oq��
G�t}��=I�@�za*��t�-(z-EQIHRWp���)h��)����5@RХ�P�:�OP�������;2���)iH������ �����@�D!�4�����JhiE#KHb4��@ҕM �1	JB4�%+KW��� ����ҽ�p�Gg�^� ���]L�;�R��]����'���笌��5�8W��1F6w]'�����>�%uMl1�h�彳�����E�$6�᥼���k�v��G�������4S]L��5�8��ʾ�]5odFw����ҫ҉C�0�	���@<v�[����e��Qt�cWg"/ -ؖ�{)H���P�Q����{gN���P�M���n#�����+9�|������AW'��Bd��D�68�z;_���>SK.�	��M4�{���;}z�9pD�̜�D�鹐��4��!?���<�4Usj=^�#�˝���T�)|(m���G�-���ۇ���TI/��?(�����.:�8��6�_�9�Q%;��[���`���$7�cYv\1x?�&=j����B�̮x�R({���-�����MqכT��ܙ"��J!�
a~=�|����=���r<�3�J��%�<�h����+7q�k��#��¦�R%�t!�+�쎮�՚~{���冪.��r�$m�bZ�%������3� r��A��k � ��ǉ�S۩��_��}���e�v�a'�V�XC/Ir`�9]Dvb���E=�ֵ1��`�!8^5޹����س�1�/�'P�Z<[&}����`�Q�>�g������,n��H�h.�l]oN��zx��ius�$Am�$��Ptꢀژp�v�^�gk���`��y��o$����*�n=;�s>�f�7X�ғ�a><�0ˁ�ф9M�R&)��y�;�P��лUXV��`P <A���Ot
�
��V���}F3]G���ld7Ұ}�0(]Oo�H�7��K�w+�a<%a����(3�dU���=fI�j*BBS�����ӭ�΋�\��j5<��������H`���[T�K� M=��սDHk��I�I��L���5����*���`ni��a%r|P�	��.��T��-����(��Y8���37x�/vAO�a��
�K�r�N2�*���
ϬD�H��\�[����C��g6�˳�..�Q�l�L.z���h�eK
V��
j�ۜǲXd�c�9Н\c�̸�D-ർ��R.�8�M�&�Kss�e^Q�b��Ĩ%���6�&j�\�o�sb|�U}%���3�'�pU�^� ����,�o�F�)L���_<�.EO�:��j��F�kd��2��&"e��#�'���#�{ K.�0��>L˘���EgL�xk�8]ޢ����j޽gq`I��k���6G9PsŌ�n��*�r~�?4���hrY���՞D��O]xԛa��=�<(UI靚V�c���x-'f�`T��ݴ��Ix��]ϋ�N���e�O0��F!�A;����F;޾�w=�f1�N-C��������bl����-p���Z�m�c�����˱�}�>�)�i���>z` U�o ����R2�{:�9�#_W�9����s�;����XZ9'��BO�F���C�d���NB؅��37ϐ;Қ��zR^�wTI�~���T���DOc�ט�ܤ�q�P�k@��*7�Mu�VeH���MU��#��5��]0��rL�Z�@8�E�6�NK����C�nُR��lm&M-��hދ�p��&�+(�A�̏EHWG�Ul�k����������,Y�;(���5rv��+<�j�V���(p�	����R�C�=�i#T�F��g�j����D���ѭ��/n��m�8��+U{�Æ�oXU��$'P{o�p�l�f�0�I��)�3��x{�4/u��H�!��0�C�^�S�tSW`��:���roFԡ�@�����3:�Yu@�Q�Y��"�Ȉ�Kװvɗ�VH���6�m:�=��#�)�xG����r]�^��k:����rE�{��*�a��ˌ��u�dE��ho>�
�����C-���О���T�R�n����r&c�w��/$ã�:�d�o2yI�x��nRq�e{�:�q�*9+{�;e $�9�D
�|D�j�ɣ��[��r3]���vjڵ5#�6�ϊ����I��h���G����tfI`}2-����ؾ���eq0�!�a���o�(->��B��J��Xw��!6j2*�XhR{
�Щz��g�b
���(�G��J�L\@
J,i.12�x����y���	��Js�kU�5�$7#���0�B��g�Dσ[�(�)+��g�ܠ�ʘ	<���H"�v޽پ��V�<i�3o{�o<�U��]�ڮ��j��惰7�9��ӈB�v� Z�˳qj��S�4;�hEfF�.��A��w%�:a�as�7���+��2��\&��8�)-��^�˸�FgY�N\��akJ�	��H��iC�����r�O�Rӻ����}��]Q�Y��$F��;��<�Y�7vKY����.�ip���c�s_�DqTa�:�RU��zY��|�ȞjI��VM��}<�ì0��}�����/\p���z��#�B�⠗�}�;
5�_!R�O5���w'��H[l81
���26��dMJEw�(ӏ�1�FH��S)���Юe�{����j=��W�m��� ���`J1�лR^VgU�G�ݻd�n��/���dĝ�Ytd1%1YZ��3nw� ���S7�}c@1u5z
V�\o\��f��a׫6��Q]{	Q��Pr��ꚅ��h����d��<��}E��bqsNB�ZVF���o��ݯB"{��������~�͒�<����>��nN��ǥ�����H�2C#e$�a��6�i�t����u��j[����!��m�7�D9!��MCO����b*�2]���ie�f��fٞCN��A�
9���z��zY�����3Ot�H!#&M�Z~�Ž��_���wU��~��Kߞ�~�O$��`��)SO+goX��^Yk.;{`��A����{,�6�5L&6)��~�AvC�mQZ�\BM!	,�ܜ4������TW�."S�����~呚DOKon�2�:�+ʹ���f�[զ����LHg"\3����vD�Ս�]�E]�l���w�z����$�ȿ{{�s�W�r�ႹP�)0q�8�E���ڧ���b-���
��D��\��'�)�P%�i5��ۑ����۪R�rՕ���F`���s�3�T����1����P��ܨi�� ,�(դ�����/1���z�����4=���L!��	��1��͸}P'9ѓ��X�<��rq���\
�>��j[\w����T��sb����:��]�b�ŮZ��;Կp����l�yCݴ����x*Ѽ5nI{1#O������>�Ob�-�r�Sf���k��dPֹ��FU6��^�a���BJCZ��G��P/!���9Z�%��o��x!�,rH~=05�C.?j{���	��������r[��􃬶��.�W��`�]4��*H7�2E�aE������<wk`��+n3�{���!��o��k�#�6]����-hғ��x�خ7��@���KH���d7�+�쎺/hm�l�%i��Wv�B�ܫ�\��(��}h���W��|m|/ZC\��x��� �X@�j7�ʵm;ד������.��}z�m�I��'����C�FՒ���gU���Ĉv+����n��~C��<�M���Ǐ�X�sNf�e��~���Q���?���%�P�5_B�"�âU*�V���Vy���y�����㇬��Fp�E��N9���}s[w��z�c��b��6Ÿ%z��w��)i=�}�7s�]N5�Tk�4��Ւث;x������>�{\O�+�J�k	�M`�F�ߏ����¨��i��i���*��%�}na�ncE�r�He�Mz��J��������gۮ�f` �Ґѱ��eaWΐ���4oF�pd�f�wOJ�2gv˖=��u�7�KL �8�w)�>��Soތi�X)���6��f��)t�q�Cy%z֫�_Y��.r���ܾ7�K�1-[I�uV��%��|?q��q�7���Z>�k�̡��J�]����|�%;W�N�l�\��!���	��"R��ݕ�/P씛j���ݬ��hl.j��!7�tt�,T�>�4O�����	�v/	��AL�����b�������y��@|"(��'=��!>�-�؜/`�~�<}^؀���������	�c���tf���*J�2 �a�<���#���Y��P�t���m�Z��+����G:��z����1�7�6�er����0��u�e��(�9W
����F.TΒ_4�wV�!pW��0��(�5z��OeF��_l"�$2��!-�\naS[j�v1@�/�q��W҅��B^S���V���Ϥo����ϣ��~Ro<�(Kı=�}u��gsj:�~�pڙy�>�������oMV��	�u-|*������P=Bo��;�\�7(��Ul߰��Y�����J፥�Z�̉�x��#ܤz��O�c�,�Kg&{VưdJ�b��o�������(�˹�3��,��C�J�v'�<�#O�΍"�ߥ��۹�� �������8fS����;ٺ{�q�Y�Ho=f�3�z��|��%׍��4��І��ڳ�gf�w�|��<���@������$w��ڕ�s8u��w0i��D �\Vo��N�zc���I�'��Y���s��|R�����z]�^�;����v0��id��9��Z�2~REEE�-Xb9�C��Y�y9[LP�N�
�����C� .|ǁ��� 5?{C��Dۯ 3:�B,�x��Z�w)�6m-la��z�q>6{z5�^A!���Y!�nǋ�k��=���ŧ)�ff,Ί�\:��0��\=TIu��l��G�-~ � ʅ��h'={6m���G<�#"t���ʡ� �3ǈ�m6H��+c+�t»���|w�.�.V/]f[���B�#+^&b�k�9�h/f�ҁ*%1�%'��O����Hn���h/9φ=����{���W"ǬP�z�kHv�no�i�Ͻe�敘+�z���Hqm:!�"�p����]
�ۊ<���vv�//e��:�Ĳ/��xolq��˷+"Cbeٸ���&#���i��4N��r��&k��5���L,j�E�s�2���u�r��@�`���~*���\Sf7kP�$w�D����P�򳲡ċ*zzO��S�L�zL?2ack�t)f�rķ��!��&�;�h����</�<��\]�;/vq��02�_ro-y��[�b�����wu ��^��ٗ����ޚD�+w:8B�š��L�`;9hG*r9YX]�Ձ�T�s����t��ʒ�Cj.�6���x4<���(�$������P�ϡ���t���F��(]���V�X�C��w ���8&.R��z���u��o�w�J	��`������`��Xɍu�zfD���XN�:�KṅG��Z���B����0=R���[ �+��0��w�\\2&�8�Ǔ�u�8=��i�"�*����"�4L�v���~{n����9 apQɶ��7�7jF�j9��ned�˥���b���q�ݒ�y��Y#SzaE�,|��?����ǃ��BϩD�`�ʴ��
�֝���[jp*��=%<62=�A�:q�6wA!���	5[E?�lEC���9�U�
�Z[,�:"4x���$��O&�Fy�/��{���,:��PA(�A��n1�n��cѪ��K�T�ǽ�ʐ���`eO-����Rkݝ�>JF�p23	���3����n�Yvr��D�'�s (�y�F
��oHBKHt^D\zeL�o*+ӽ�(Nq)�<A�9V��!Y����X8vSb��{!�j��Sj�(���\	�JCp$��c��˃���pẜ�C����X�{�^b�����M�d��o�.�:��|fX��o��X����*|[�5v���.݊�G:����g�z�fŘ���͙f��)����N���=�G�W2/y�ۙ�9�^T)�+�߻k+W��w�2�_��|>��ߩ�=r��ֵ��F%�r�K"�P�=���r��R���b���O�&�'j;�9+uٮ'��9� ����C���{��e@����R���3��p�ie�^��N<��c��\t���P	 �zš'�q�vX8�rG?����*I���sH�Еs\ޗ�Q�3�T��{ ��+�7��"8`o2��n�y��'9�yZ{��Yċɾ}�Q^�W'���yyD��m��1�� ���5�e�E�/x�rr�U�E�SQ6"j1v	��gs���+���6b�9RA���-m%��L-�]��.n5�2']q�?j�{��[��lm�#�����N��/2�تdel[�4r
�$0C�B|F���Y�r���t��΀�L�_u6�aşY[�����`啥��A���8*��+����b⯯"F���i��2Ӹ���UV����Ԥ��(���o�Z��r�C��ec������7��B^�X�����V�~����A��ga���%#�h����5�
}���%贖���V�ݪ�U��R�3�,����+�ܬ3*�<W`�)�yemH{���X5�0m����s\8��ri��`����;W"Or5�܌�9�z�v�ަ�����o�˓���G�w������k.��a�װm\ڔ֘I�Po׷aÃǼ��w����s|��l�̺�+�jz�yi�6�zkslɱ����(�v����'	r)�2����:��9C��6ɫ=y1��ȭ�`�<[�~��2D&x�:G�g0��JE��o��Ls�;�d���������Ǖ�S�����TG�׹�,,� ���r���5l�"U�X5��G�	}e7Z"��;��.�՘���A���[�=�hu	 �v�voǍٛ�U�`��뚟��Gb���/x���\oڋ!��T�0�ph�.����X{fڠ�j��F��\���o[Ʋ�ә&�Tfԍ��w��2�<����`׶'�7��`�q�M��I4�m�-��O�ށ�l�M�gO�/m�OӍ�%�E�[�� �%�����-�Zrˠmvu�v�3H��fIL�r�X%Ԅ�]�x��}�T�)�y�|��W�Ce�����x�Y�ך{�7G�r�s�xy��/wa{������MĦ,RC�����X�WVe,(n����3�e��Mu�������B�#�+�{�������RX���vA�����B�j���g D��bt͂���7��x�^��a)�n�liy����vB�H���8��齽���2��5�X�f��%i��|�k٬�w\�-�S�N�\��ʴ��#dcgr��u��e��^�ͱ��R5����A(5���ݭ�\֋���f.�)S���.��@�湁��afιPi�/�<�	,�X͂E_#��(�CM�96��cUPGE�ҍ��Jc��<��H=|��E��.�6S9v��:�N�0_.���f�W�2�6�.�p+����Ӯ��6f���т����I���듄2U͢��Sg�'3lP�S3����CR_-���GXat�їOXgg'��Ć=��{�ȯz|��6���Lt�=���{�I��"���* Js&�!��>�Lk�������H]���˺+��2�!���A6�s��f���U��Vm܍�6 ����Ә�<�w�[��^���4�1)Q���<ΐ6�1�sgs�L /Y%�i�aq�(-[�#�n��ѱ�謸�5Ɍ�ov�&��Y�4 7/j^��(�����>��(l�5�Kt>Y7��?�/ ��U�c�=u(Kǡ���=��9	�myfRپ��yU�o�}�L���oF�\3L~���*�� J7�ne�T����7K�G M��H����m뿟m��3���W�S�\CX��nT�mJU0Deuj�r��G��׹�&��"�Vj�F�c�Wg�~�o�|��h
T)j�hS�t���}>�o������������~�D�'$]PP�M ��HOק��<||||~�>>>?_��~�����B�#����#�RQ���!ABu�(�IJ� UR���:�(
)M	��*�
�B�J(Ў����h(t��-�����J�˨J��))����
: 4	��4�% 5I��@F��ӈ"�)i��S�i�� u.��B�JZ�=�Rl4"@�C��5!�j TQʵ�ך�,U����ՙl)#S37VC����2�L��g���*#��ToG��F�/+�u����|���^�"� �K1ILDbb6�R2��F@�Q4\Q��(�8 H��}���������y��q1{�+�~q�EU��P��DZz�u>��8���[����2�<�j���u���n�'K�&lo��۪m�{2A �0��XZm[�P���4��ZOj�<K�5�7 =\*J�7���n�k��M��ޖ�o{@p^m��!r�P�H�$.��-J4_��O[�c	�+�y6��g6&5?5��O^YX�g�[%�he�C�_u����b�]q�;�hY��a5�����Ǉc����^� �uρT&U劅"��&�n1��M��O�ETf5-�]�Jk�C���s����[��M�]�'�)͔�#j�2�̑)��t�>!*���X�1Q�
K]�e��Ź8�f���l\q�}l�WN:��y��ԛ˾bxRq�f�����3	��B�hj(�,d4b�_@�B2΃~����[�.�_{w}�nC��h=��ba��]�����(	h(-����Z�6���MD��~������ݡF�mB̠9�֮R{�N���D?&H7��R ��a�'�a���n!���W_�h��͑w��**=�Ͷw3�oM_�MSA���p}��������ȥj�۷�{"�Vw�$�����ðE�{-8���z.�L`�Ϧ�������d��s�uO��*�~��@�Q�::m��>��o�c��7������/���-~���d�+qZ8�,*�Oc��U�%=�4��8F fR��.j�z���� ����S��\(Mu01���Bչ��(���e?yY�>|C�C_��^�ۻ�%ں�n���HL9�R���!���OZc��pȜ�Q�q�Y�� �<Rg>�M���u�N���Ku�Ɇ�t@��9H+�����,7�3L��b{��C�A�ރBY5R��36{!_v�`�dM��J����a��c	+VK��B���)�E
��&y�.ӹ�:g�ak�Ӱ�ȼ����������S��V0O��>7L��=O9^k�Pk� ���+�L��@ڤ����C�Wdr���4�m:j鋇�����}@��\�*�� �I����{��	��-��@Z�*�P%A���Ji��íY�URE���
��{��g��k坃���l�کf=�Jm�d&J_�K!���G�(�?���H~�ȁ��JK�c0���F��!��f��}��s�h�0��0*Q��v��5)�s��)0]�ܷ�"���G�i��]	��ر#����� d8�c
�v�˧]5d�|%����m�t:9Z#���Ar:G��]��ӭ���y#4;�^�˒X�L`��+_v�f*��׫��aJpf�Oy,�D�w�ʫ���!�w}��9��ב:��<�Sԧz�S�(ԕ��IT(��B��I��{RB�����4��@���e�~�jRtBx���TSL!�l?8�e۔z�^a�L��<�wJ0�ͪ�2^p@i6�eԹd_@��)�G��Ô�j��&��]�25�V� mcI�=|�p�m��Gjh� �0�B�逛d^�
Vv�8�eOC�zO����4�L?4Y;&�n�Vn��vOs?��n��R���1Mne�ɱt=�����^F���0�a�N6@����V[9y©]!�K��e0M����/B�u	�lU;B�P�����Z�'�.�'n�
��R�Ds�w&�A
�pA{F0a�f�dmqpȚ�����stԔ\Գ�d��su]Gv�y��U��[�J�Y�K�� ��@�'��hn�k�Vsl���&2�L�IMʧGVuk�v_O��Ǔ���Xܭ�_����]a�޴��d�f��j��j��.˛ב#���؃�}y� :������!���$= ���_E��//�3�<�[8jC���g�8Ux=��m�vQ��mS3��t<���*�[��4�g�z�~��E�^3������l墵������k��W�V�}�u;�($B�"U(�ݝ�>��s�
�[�wa����M�_9�^�5s?���W��}L�}*#��{\����x CG��#�a�$�%�ލ�נ^_S4�Aa�T�&<�k�����n��/k��\~���e�g*���(�4�219�MO��_F4��S6_w�H:��N�E�rώP(���;u�1�Ψ
����RW8��HB���IףͰ�o�3� ����ݜ�Qy���m�)����ɩdIz(ΰ��Ƕ�x/�ݙ�Q�sb%��g��£7*������ٴ��$�<�D�W(�E�Q,��6r�Rk���*��sgu�efB=Q7����f����C8HB}fQz��9w�犑LJ2��Od��b��~�9����5d�#x
�z���i��pg��f
Gl�8��J�|1	��9�QҴ	i���VZ�f�?<^�{�,�5r�*o+RD`��>`�7��>p*�>�\��i��đ�C��哒͝Zp�ʾ�U]�N4�����m����6@4�9��-�(����<��w�I����J1\4��{�Z9'�+�d#̷�b�))#��Q8Sp]��&㼹�Nod�[�k�lǨ����e�z-���� ��K1��8N~�v�_:��9� Y�li��{�,3��!��r���� �,�(��gz{_���OH\�\.h���c�^�%Oy���]'%�X�M�+�MآRyV��Tw	���>'f˫l$ڟ�x���A��
^*�q�#`���� Kb�Umw�)8�Z���*<��{�n�jDȧɻ,cq]ݷ���&�Rc��o�w�?�U�:U��D\F���p�9�t����S�4e����e�i�Pϙrg{���B~�a^D@�����;s�~}�����z�:]�R�LY�ҋX���V2{��*YY[3Y����.���-3-�����#FbƇ�{C��VW��y�pA�X^���ۭ@eyl����T��W�Y���&���q	��`JB�Y�V�5�%<�ط���4��ZJ/�ecw[Ɇ���9\���%x��q��!�{`�,md��⌆��e�����	0��*���a��	SѓQkf�F.�^�<\[������Ej�GL9G4x����Ex-��O����$��3��PU��s(J��]�=�B�ǐ6d��=�5�a>sF;s[=�E��]�k��h���$
g#Tq�]o
ո5�J�xD�'�Ds���Zvl���V�상�������
wcq�J�9��9*�y3S��d�{��b�Z�O0��^�&���݄�'�CDԕ��ָhrl��*_P��Nd'���\69����u���n�_1+1��
	+
1����c�^\�������|>�1���6i׃���w���N幞̑ty!����U�z��ʚƧ����6�$���'7{,�.*���Dϛ+EK��dzd:]"��;^df�3�� ��枂P�+��=�\� ���@��<�Ux�7;�˫��!�X�F��m�*k���IPp#2��ٴel�����-��cK���Lv�����\�ֻ�B��z͐�b�+�I�M���6�8��󃞗�b�H�4�&�j�;��Wc�fE�ճI}"�y�4�@ύ7Gy�"�7��10UܯR�a�v�����������/��v+&� pM�D�6;�5��3��"Uq�}[�R�[��#���}j��<[���`��i���W�H�3�-�~�8v\�������[N%�Uv���|�$O"A=���Z����K N��Q�L���U<��w�:���u�qk�x]��]�����tS	F�{��r0��<�A������ˑ�j>��2��M������5,鞗J��]m�.��6Ӭэ�z���"Y��]f��bi�l�_��qJe�Q�|�Vr�ޝo|������W��]�v��l!��Qۍ��YZ籑�s��Ȟ%�MC:��eb��[nu'�%�l[����@�{�5>��Z��:��E�u*�/�֦��=���;��e�^�
��s�-ī& ![B���9�Ub'��/:z�d�٫4歭p�n@rDj�&��b,�ٝy㙡�[�$f�����.{G���_*�Y\�8�fr#g:xS6����/M�����`�XVoJJ��8��q�qM���v�� }�A�sh.h�ӆ�DЫ��>Ƴ�W�B�6�"M^dnj`�e��q�j،���ܚ��v�r}�ozMO���L�����ʁ׏ԑ���n��7c����:�l+����ק�=wv�,�Vx��{k��7�8ǰ��3�m23f����@t�a|���-��an�ڦ��J�خ�8���^�9(*�e��/�@�a{��]v��77�Δ���6��|�o�{�<�*Vcw��r[�K���厭u<q^�x�9��a�Ӝă��ŇC��oA����5��%�78�T��z���� ���*ћK��7��?��U�uU��:*ɳ֛��_ Q5%q�@��O��d8�)�ѹY�	0%K�uN#���������9���{���l#���
½c
��XF+˖��k����BD�:�5�\���pׄ�r���c����m^�d�]����a_�f h���(xXk�d#W��γ�� �p�8ӓm7�1x��s{0�CwzZ08%�0�wPǚ�r���f����h����x����T��g:{w`���et�}2,s`|>^w�F�OOP��븘����2.��X[y�����R_l�Y�Q��@�X��������ޛ�us~�}�g:l
������㧏b�^\K�U�"":歪�i�ڭ0Z����9�\-�o��́VT�R�AOL���j�[��#2�StM���2��\k���O�_.��$Qx��*���"�ߍ�
�ļ�����{c{'��iz/�5U����¶E	�F�[�Ƭ�&���6�������7�e���xo��L�[�m���7�S���;屝�u2�Jr�>�Q�3hUԔ4S�Oz*衲�`�Z�	�jQ|��]A ������z��r˼��J��X�g�1��b��)i���'Ô!�(�T��x�ԝX�[�51��}C��od��������!lF�t@ݭ�"�3H��˽ȫܺRx5�z1zԭ>��θ]�o��Awy�1qw#�]͙�S;{�����Cfo�a�9�ؑE%vg�e&�B��
�#���ѩ ���k��>Ӹk^�-��*s�T7��)n�P��FX�`�=!��Kʪ1q�a��5тU�,	(F�a��~��]��+ܻ��9&�s+y�p��C�ξ�|��{|�oC�#@@YZr�-!�{iZ�^�tN�D�R@���a����[X͢�-���X¨rtd��7~���A��*�b���U������!�w�׺$賒��C:�:2,<%>y�^�n��v3�f�oL��W\bw�;0�Qs��Q���9���!]��֕R�������#�g�����O9t�j�����a FU�u��s���Azqr��m�v���[�6������khɞ]�##]n�>C��b9�ڮ)����������ʗ���#����3��{ky���+��w��E��C�L���z��̘�c�#���{ދ��Tͱ�u/t���s!a#�v�
�$²�V�zXF���,���q���љC7�yD?&��e%��/��4�Rh�� �@�l3]yUA<�ۈkΫE�^Qu��P�m��#��Ȋ�F�����x�3�fNI�<f�<�L6]s^Q��� +��4�M^�t�������P�DD8���0ãLކ̧��T}y�&8�=��n��2$[��\�!@��]H��kzc��x���6rE_�<�H��el���f�` Fǝ_-�z���3%z�ov�Cʴ�>�-MмM�V�_*Esq������8a6��!���[��*-��T
�=]�U+�E*J�]Ӈ�'i9�W�֣P�qͦ�e���`n�锺
ٴn�x�k��+uMʀ�Ī��5����X>�a��}�M�#�H�7�V���'3.���g��V�Yr2���6�Ǟ�l��qő��ӿ<-��;guA%�۔1M�&*��7��0�z�k@Ү����z�m�GovgG6K�5Zdu����,�yd�ۗ���������d��s�6���@C�x�kn�$|F��r5=�S�n��'E�˽����

i�<�٧7	𣏕&�lA�F���V�8�6�M�I��y�g�w���=���7=��;w��GC�GoNf�����!�-�fv��`p�r��/����T��،7�ٸz}��[���}M6Ov Sګ��^�	�����v��6�TF�z^��x��U�f݋i<ʡ}}1$
����c4�bݸ��V�/�(6y-�8e�@3�z�탓/D %�z�d�у���#��N�Y�����Bʃ����,�6�76��g�����>��p��p�17n�����{|��>��&�v����\����q����F�C�n6��`x0����T��Ŵ0��=ä��t$ko��H쩴�fȖK�
����D���IOO~�PMf���MYc��<6�Kq��9<��e�hp���Vd���8�ScX��Yv�8�֟Pm��b�'(��ڧ��;7�������Z�,,�ClV�`�̜�uJ�����w9i�/��c�!̵����'[��3by�!�����T�yM䩳�(tw��R�}/vl�o\�<q귅��*1.���4r9+�BS;�bWt{��V-B{���7�:�M���E��+���m��h��e�[>q1:wl��'�������hX��I�Z+m.ݮ��i �"�H������?�b��DNҵ���7	�8&�1�^lU��wO..��:�&ׂ:hl#Zf� �T�����ƻ��%��_���A�N�2b����z��.��.~ܞM퓽A�q���!��p������
8�[�X�F�A���c��9R��Ft��N�f/�XÁ���3��q�`���Ntl��,��^��򅉦��&�}�u,z9�p#��^�yNrz�GtE1S}M�v�n�qX:fUG��˷�v�
餞&m�#�Mf���9z�NY4�7�ik�,�i���N�k?37]���hӐ,X��a���2Q��ޛ�tQ�$^G���ʽ�:�f�0�s�>���~��?][��~o��+
Ȱwh
��jf��l���V���>����F�'�����E	[�F���t�ŵwWk���{���pa�u�T*L�	�J����)�*`*jM�޵|ú�����w��`y�%��-�;�䮽���Wԑ��h��ʜ:#�ҔXd���$��A���C��T��Q��3Y��A�e�\(�9�sާXYd�7�
hu��Je�)E�pܸ:��3:�&�1SJ�eM0�*�:L�zg�O��!�@�J=��
Jbh��{~=�_o׏����Ǐ������_��F�(>H'pP���I��}��o>>>>>?_����B����K@�F��ҽ���+�t4��t�]!H|3ܽàZ�;Bu��I��4� ���P4��]'r��QABw i{��9�ԁ�S�X:�4�Bu%
Ӊ�1�"F�M-�Z u��y4���B:���4���n�P��Ĝ#�g���5Up�	'�m�Ӥ�#���O=��u~��փX�:�W9}�ud��r�
�8�qY*
7l��Î}�/�꿯�������Y3ƛ������}Mў��oG�)�p�rӝ����ʍ,�-��o]דt8�Ϸ�{6ǈn�0��M�^�������=��������a*�ɞ-��H�����ᤍ�ktoR���X��c����JVz�klz��7{���"A%�ח��;�}C�ګT��%�ی��@�c�ILm]vnh�$GY�U����F���kb&s_�u���
�x�CP*�~v�/�������.��F�����\5(8�mn�7��oi��,�C=qa��q,���#��n,}�y���kyM�*�RrAڸ�����x� -����R��u�/.����nuwGl�B�; �
F�]^�R�%U>U��(��y%W^nU�W>څ-xz���x(�u`�:W�IX/ױI�<U �^��1�(���$Y�����){9�W�H��I��V]�pVC��,J��^��{E�)�jN�ů�ՎGM]��WKG8l�gl/��9�
T��b��Y��qJ�H��ZK}��r�U��A�d��OSJ��]�gaղ4�w�C��s;_,f5�=sɜ���|>���5�A$m�h�Q��RB�\
��3g��T��y���mڝ�\�7�Y�nӸxkE�M��!�؅�#V�����V�4u#z�� �MK�f�E;pG��eU�F�0��tp\%���ۜ�����4ԉ���}�s�\�X�fݸ��q�B�Q^�$^z�B���"w<����U���'2�V�/��||�iP▷�� L�#*�>g�t8��C^q���pf�
f/ot�+�b��b���J��<v�`g5�ݝ���l����,lq�?^�qX�&��1�N\R��=�R�k������'�Ɠ���;19@Cz³Qi^6`����$H:6�P���o�Y�]�-yX�?bu�0"0%��wt4K�6�&3<]������cl�49��p�<q�k2ȐN�S�i[LbF3{�#ڛ��kRD�n�n�T [���풪^����ܨC��ѿO����\�n��k��C���6Q�l�x����
�~.����6j�k�p�U�m-ݵS��-�I�o/�]ɑ��f�92�@_.���e3���Y3.�H�m��{w��-��C�p|||G�Ǣ�OV��F�b��_�b��;dl���4�қ�P6Z����>EL���ו{�ba�{b�\����d�Aj(.
㧏b=W���4�[p)����h9�$��cz�]�nκW�w�=x�(��O�H�ؔ�絡�Eu%|(�>��NjOY��w���"��Y�_.�k�k��z�otm�
tX�!��b�ɶ���1��W��'S�7��?pj��xޔ�������5���\�QU�6	�[N?Ѝ���L.WFN����E����Qnў������{���]�|j��7r�T��O�ؽ��\:�-�"��qک��ƍ�x8����#2z�/�U|y��Vc�Ra��ɖp��3l�*lL�1�����맆ymVd��?�@~�U9�O�wLT�
�'i�8ʚ�i�����n��8r��sz$f6�VT��O�|�d��JK�ed������|9�7&���v�bz`	xp�~]g(��V� ���3�߿v�2^����v�n�4ry��;E�?��/�%�{R�a¶<�F�Z:����<�,�vZ�Pr��ݎ3���)�ܻ�������^��-��0��4_� ��{`�@�7��E�8o���IƂ��Tz��8Bٳ˫�vV�U[lY�X5�kVhژ�q�m9 �a�0�V9�t�6�ߏ�۷����U��IO݈ʐS�T\d�mRx��G���3����N%c���*���{��:��1No{Z/�(���x���s#E�ލ���έ�q��<�{:�&��B&��/qC���U�@
�H͕��U��M�{G�ww��~�|=�T�;�h��W%�/�3EI��3�b��F��?^��t�FUC��.ɓ�+�2[�[�c�F���y�YA��'�u���j;�n�@�l���y:�Լ��>k���F}��G��%�YމB���Z�KYʨ˷c��sQ��|ԒRc�S�)ܷSِ�I�!V��uЭ���3�=Ιߺ[�!yQ������*W�&B\�2+E˛�t�O��eT<)#v��Ɛ�P�`��cpm*Ƚ���	tkz�s�z�X�μ����c�������{CD�j�;#D���~��立�n��h���秀�<���7ay�����%�����N�Q���`��M�D.-���B�������ᙂ.�������hB38u�9^��(�U�W��3�]o|�m]$��+��|w���?S���s��@����^��Ԫ� \�)REwYֵW�\�j�9W�x�J���,s�#�;`:��	?��]W��HM�]��RƠNͽu��*c]�kl����	�l⺽��^�U��ؗ[�=uY;}�O\ہ�QOR"C�kL�=��>"k��1�љW0C��r��3�k��mu��|�W�.���.w����o��	`G4�k�Uބϴ�R�{���� �V���\d���r8�{�Oi�9�4������S�oV���C��QW	?�[b��=��'܉Ix:(f�]�~���u��*��dQ���Y���ѵuٹ��`�r�;�e�a�}�7��9vîs�6�ϭ������%ow&�c�V\�޽�X���M����h"!Z2������N�>���g �ʅ�Q��휒����x���1/63m�}�����o���wV~���,S<�N;C
�H'U�����
����_(Ȅ�Z�[��5���FmS��m)�|�o7��ѵ'L�h�s�UUn��!yJ�\�G�����n%�3,d�=�̊�]�g��t�g8��$��)�#6�j�L歀@ր�l՗H�W�5v�A��=Y賽����wO:
t�.~%*RUW�*���:�'�M������LL��oz,�2b}���ýВ��%�I�<w�㮵�F�*ƌ�"Fp�ތ�}<�G��&���(�-6y+�oH��U�:1�5�6f�M����@��zæ0����A�5l������V�n�o��c���ţa�z�\eb^�[+���k��6��GSx!��;ޏ5fa9N�\m,�ö�����y���>8y�s����i�c!��a��'U�U�Q�qu��8�w�M��q���pV�Vj(Js1s��g|�t�)�����F��g���T&ˍ�>������|YW������pm��3��R�bE����(�h>;�a����*��mt(=U��n;�5Vi~m�hYA<�Z�fI=�/��R��Y�S���r���+Y˖�n��F�{��)�����9Å��a��������<C8)�8�%YHf
��w4���զ"��:�������"j�KF����yз)��dy_������hw�����z����m�ѮuR͎�2���ƒ�k����r�K<yP}�޶__F�Hr�N�v��x�n�U�-�eXmT�(G=�,Qd���F0;�.Mx^�}W�8f��/����6�rJДK���;�rYŎ��E\�4V�g�~62�7y�:��Vd��2E	hl���Q��fݪ�[(�%�ӷ7�-D��g,�9��<����B-�>\D�j1�Y�s��M8�N>L�k]�g���m��t:���Y�V�pk�UR� T�RQ�]�79�׳6ȫ=o�4i[������)���o�����t�n�5�Ķ���7��wb;�W�j��P:�֗�!��X5H���b�.a�z�RV�`�/G7;0�x׃l�N�oP'�[��]9f8i������d�t�g��9�������T��Qq���K+�,(�ֻ<Kܳ���c�u�^ԡ�lѩ��Wt�G�
����H>�k_o��(�����+�2K���u�AL�r��ɏ8]>��(wG:��[��@U��x�]l��Y���V4�=�o��O��f�}�9��mW-�j�j���g�k�0Y+��<�� ��]DF�1������UY���-�]�k���9�إ�>��>ٷ*�n�}4�g����ۂo�#m����XP�W��䦖鎱EMEa���9�+ͬ�T`���e�Y���'��dۏVU��=E�e˺�k��n�i�Z­����|�8�mHRh6��|�!t?b5ei̾K�ɇQ��ᝁ�oR��*:NϨ�Xcޑ�5�)꺄rI��2���@�L�|���Rԭ��~q��cߓ��jz���Զ1�p����+�ξ�a�m�H�R�鯄_�z�h���W�N��D��{(�z���s�̷yX*2����F���vS���^yb#��YY�W��M� 񧻜�jw�9�+s��9z�Q窞�k�d�ϗ%�/�3EI�j;X�3S��m�3��z��_ޖx��tݙ=/�	9����XPS�k��yWٴ��9���/�x�j9[��%�;\���hX1��dMh����i�
��h���}�y���(�Z3�lm�Oh�C[4klkN�Ʌ[�-͛H�es1~]}7��KI��gz 5r~9"�_51���L��F�o7�Ҳ4�.4ܝ;-���E���O*�z�zi�M3�z�������
��[}��|荹�7�7zN:�'�hIIY�k|�j}�n�ȑnB�8��5ʺR�����cA�=�|Nx����J\w�6V�U9̖���MHq@�����Tk�I���6j�^�-�UR��#k[	��W7Y)��w�ɐy�����i/���!��3݉u7��y�*K�>ę""�Y�m��-�cݬP��*r�ltYV��՞ˊ�ʧ`�$��s�`K�w�S��{�=z�B�8�A�y���3�M鯗n=�9�ܜ�|y�����ݡ��M:3s#�?f��dk$PX6���W8u��Nd6����/3+#�ȫi��Y��|�Ɓ��=���ϟ�ڇ���^&j
�v^�ƺ!s1e���U����j��mZ�H���O,�'tW�b�[n��]:���b��?�u�&�y���u��B���OCw���#2�atOU�:zI}q��k8e�of������k�����29�:H������ñ�$���pT�VVx��ź�@��i�&��C\�[:pE�ےxX��k�y�x�m��x��G# ��%ݶq7!��L]\aew45Ěy|��QY��J�n���Wܽ�͝��i�Y"�2}�E<�,�������u�^跷m�X�A+{�-�/<����7#�0��#�m���#�ᚂ�F}�+�]�m)��9�6Y�B�׽�d7�o�/g>��̍h����|A�JIa��Od����sV�'%����Px��{Mn�RA��ǈft��B�D�|�G:�Y�0�)R�|�����}�L9�-��:4�0�b4*��^����{���I`���4%���� �Zu��FT�a=El��q�.�б���k�Q��8)�K���ܥ�Ɯ���n������a�kr�6�8;�d�5l������=�N�F��[����I�&2���[:?H�XN���K�O>�n�w�~�x8ʫ{ p� rT�`��4�צs�K�'�Aɜ���M�m�revm>[,�W���w���}�m�S'�]�]١#��-{xj5�����9��]�:��Jd!�� �%����&_-q���Gc��fX����L���]<��KaYq�ty��R��I�W���|+���P-y|�bI��<�R��)���̜��7�Y0d���Ґ�Ck,�T
���A�.�$lY��.�߽;m9�&N����h��e�nB�"����oZw8b��x�Y�\x�ڬ�2�oP\NI�8�n��iN�͕����	 _���Oot����z�!�ޢ�}`v�"^d�z�,�-�����tg�̒2��Q�=7���+�S��'���G��1c���i�r�``/���oi��i�yC�_����3��M���7�Ǥ{}
�&�=�n��9�i�߰�l)���z�1<��x�i��.��0 j��)�b!�:�M^��B���6N��y����v���\���8{���pK}5OO�w#�9��"
c
J��1:���ㅵ�,��n��k��]�K��zf��������R��;s�O�<���U�� �^��F�����r�����i��ք���,4�
�Ǟ����>��y��uAӛ����Gp��|�`�i�Ӆ��&��j���lx��Le&;��TG`%�Z�Mlc�Oq�9榘c��gr���{�����߆�h�AR���N�超X�E{|�S�	to�l���{g�2^�ɍ��U�Zu��_If��Đ7�����tz�HfŚw;}�c�����z�E����x$%���~P��{������ϛ��qޓ�ޕ���4ý��hz��{璘�O���Aժ@�I��;�2~w�K���L�m�Գ$��jq[�r��*�]t��]�4cN81���@[�޾��22����ve;N@a����ec�����W`ӈiۅ�r��j���%�����@��굺b�Yƒr�Ҡ��yi ���oxu!�;�s�}�1=lb�I���Zw[֦���)�q��9{�]\��1�m
����n�����\��Q�rV�$Xq�����r�Mx���n+Z){2d3��\֛���Ҭ*��d��*�Yt�3��,���Qt�t�������}ٴT� Zz˹ҊD�i��C��I�ה��t;'!U�ԛ��`Ͷ�#w3f��O��F`��G��"�n�.������/	a�왨k��8�)���FT��%��{B�)�yv?�Ա͈�2l�y�3r�^�0�5b)��'1Ƿ4���� i'���������]JV�32�kL�EͮT��L�����Aѫ�gv^\L=B�e��A��}�n��w�G��}{7缔)���>C�0m�t�㭴��q0d������|~?��������?\���- R?`7vA��=K��߯�������~?�������E'�P�)��i]�E4�uݠJfO����ɭ��OP���(t��Ԇ�Q��ӡ-`��'L:M!��uBѡ�A�률��=�Ut��a�.�ҥ.ؤ�Z=l����JP���w�}�QAA@hӡ)�i
M�����R�:��CCC�u���iiz��{���)h:����CHS����ؓ�K�V�)%&��H���v�*N�.K'LS��4%(�����ѨԾw)"���	�s�G5mŇ��;_θb��ws
��((:%:s�p�0H$��D��>n��a�l�ʑ�	m�1�B���� c\��	R�}i���<_��d�7��ݴJ�&W��:�-���a����i����\�kb^�9TJ�K9��ZA�S�Ư x�`N����5F�j1�.�)���DA2#g��iP�+J&c���Sy)�}�00!#3'hB�؟P�.	N2�՝G�n���Ҥ�=d<���]t�J;s<�}���S8�Y���f�]a|�/Q��~�͸���y�\*>��;�[�S����H�Z��qy�x�ՁxVhE�7��{}�4��̄}�H�v�/��7�\Csuxv綅��	p�`����j��X*w3=���\�Is��jw�wyux�A�YJm�k���H�n̞�Z/9��Y�i*��=��õ���%G�?��rBz���h�m�fҜ��^�f�O0�|�X"�j����{A�{���ɯ\�.!f��
B���ثǯ1�oc*y�hٸjg���8[=ы�/������g�j���һ�[��K=��b�7U���mk9f��_^��ed�ö��(���n!_t�7�a��)C��׉pF'�����+Z�@��;9���ZG�[�j����d�{�
|���w������)�f�u��*@n��\��ᓽ<�j�R�x�*6.��i����y��n���٢5[�[\�NjD"�^�|�}��1�/r�t�4��f��{�:p��GR]L�]�u`i���@z}�j�'(��QH=BY�,��h�穌�#������2ُ~�Ab�l�3�25���&z��;<8�GV�Z���r��f�vB�`�n�L�s��f�˝��A�B���9�zz��r��)(�Wt��v�O��:.m�1\G`X;��Z A�����ORQ�	�Qʍ�42:��R-�i�������U�Wf��/5�d=���#���G��-��wNJ�>����ei�jv����ֱ����u�ށ�rFO��lo�;0�K���"���JB��*�{�Y��tY���ג�!���џr���g�����&�vg�sf�_{k�F]�1:��l��8���Y�w\��^�����u��F���Ez��v�k&��+q�.-ռ!Ҳu�Ħv�ۧT��b@��\��v�v-�"�#�t�L�{�S�Ԣ|V͂vQ�S����\Zpe6�O�Q�ǤoIr��tq��p���ᓱ�ٛ�����|� ��b�#Tt�6������Fz���k@��6B<t3Y�F���|L�����x�^Y��<
 ��{�ڮh�:�DЫ�/̈́d^T�ն�&�O7�jE�[�y��E�nk/<�����:|U�WF�Kә����3���X�uM'�ҩƗJG! �U="�՞�����uaA8�-{v�?#Vl����\��#v���ԓW�!�ag�+�aߠ,�k%r�X��3�];�ns�ڃ�ø���zM<��9�f�&���
�B��N�Ҹ��ޗح�ˍݤ��.xm�����YxJ�JA��R���_Aَ����S�˘}mNɬ	A++T�(�<z*y��{=
�� 4arӥj�z,�f�$ p��O�F�j�WŠWIU�R��ׯ#>�ͥ�_���g�7������ч�1ڟ�-�!s��1�Ī��y�I"������d��oX�-S��ZQ�W��-��s�ҌN���p��g{(ڧ�TF� s)�x�o��&�`���z$E�vOt*��s��ӻtؔ$��i�r�ap��/j_)ݮ(�V�r"�n�'Zګ�������7Y�OO�����F,V�l�e�FSyr��rF{��^%ܯ3D�LE.eE�m��=gZ��R��1@Jݕ{,�l͠k�t��A��lͼ�D�+�-��c8l�/�˨%�J�eW���cXX��[�?l0���o,�Ce�[�5@��gU�uفX�v-�kWjD.���.w�;l{da��T��dnf)���a�U�ׯX�����Z[[���e��-� ql����"1Ae\�TDf����C����:�qV�f��[߽��'܈D��M
��j�:�Ո;h�؝6�L{���l>z�X���c�goz�!����e��K�v��3(��<�oiH�z�v�
B	@{�5��-e�U6��j��;[�@��k{H4)Y����V�	�; 2}A(�X�*�=���z���2b;PYCJJ��*���;V}sR�_}����{q��]8�ՙ�"fn�[�<�Bxk����� O�?baS��6?.���c:��4�1���{C�7og�g��B���VPS��X���p�z��s�����Ő��^��/�P�#�N
���W)�����
[&�g^�Q4.Ι�����o�AH����|>�,����I��{4vn9���F���
C��� i�$_.�s���{�P�R�9����������n�as9Y�T����k�c�c��	Epr
���t�	9xK���{:�D��$����щ>Q��O�5��P譠'��\xW͎ITk\:�$٦{�j�N'w"���ϯ�g��Y6�8��5��赲/zHS�ͷv٬3/3V?(���}��;�gS��W�F`�ly�t!�j�׽;T��1�0ot���f%Y�*����K9��=��e�����%���cf�[	M8���|�q�&#���m���mLԼ��iqQ��N2I.xx��'�]{�����8%H��Y��I�Ϲ��m�U;\zq��F4�a�2f(rz^���#�7Zj@����5]a|�{G���g�LFrG�r���]ۭtEd#�Vuk��0��<͚֔��܊=)�+��!�%��9>�~��]��0Ou��b��8�KJfl�i!(��iL�ni+�f?�9�E�����!
�Y[���­U7�# �ԁ����8ׯ�e��	��=\Q���M^	,��U�W��t�����X3�<�{ �����#S���ҽ�xk�k���䚰]f)z����S��Anb|��=1C�C�c,��5�����:���U܎8�������Z��YJv)����-�e���n�t焐ѝ�J�B�}��Z#��0QƟfґt�q��4E���u�װIm�c�T���,������,H��+��=��;L�yxJ�U4z�nb^��0#j��}�a��]�d.�s�*�)F2������w��{��j/לܿ�{�����Mt���az�/�[���Ym�f��͘�g�ѯ4}�Q))�>�7]:��bA�t�bk�M3�5]59�8�woCwed�x�&RV9����uq6u�6�.�r�I/R)%s}62��G�#�ե��9R�~O�k��*Gsv�7��V�F3n.�l�c�/v ��������5�_h�*_�wH]�6���oze��5uOH��(��R���βXJi�O "�J�&o�}�s�s�S޽˽Z���������z^C�m�h�x�y�wU��{���x�P���j[Oh��oX#p��\J�wxi����÷�M�cZ�K�Jd
��y�����gLh����h��2"}8�4�VG]V�SKt��8���z/�������7\��h̀�������M�~��y-ɌT�֝U�o��'n��sf���������������uÁ��zA���ѺF��q�s��.��Gd�1��lϺ��C?�s?����R�C�SwL=���Y��De�	@f�śS�:w�L�Ǟ�P[��{��u�M���e��ޭ	а����Syחу�0�A�� �x+mTfa��{&M�f��b��0k���v�D��̏,$uv��+�c鶧�&Ԩ֨8�Cn��tW���7�,�1���	C�I�D�vC�������8��OӓU;{������3���{�,Ϯ)�D�hAd`�w�Yh��[`�/��N�[<����u�y�Q�&9N������בx�0�
��E5/U6u�۸-�8�[ߢ�0����� ^?g6���f���t�B�1 ��j��`%�:+�99d-k���0����_��F�%�N9�1�H�u/���(��/M��w Q���/�;�w�]v�R�
��L�#!Cud�%����Ͽy��n�.�u��p�Ѕa��P^).8�=�y0��{3�}P���[E��sy�;{��Ѕof7BF�Ҳ����{j�y��4�u��Ra��j;t�L��n� ����t�mi����t��q�-v��#b W�Pn��;�ݷ�e��ЖO����G���ؕY\��������-���������ԗ��e!C>�g�|�dy�oTASJy����־���u��^,
������&����7�_�Ҩ�z6���3�s��f���O������y�����4:�?��GȾ�>f�)9Ej��R(U��z[�	�J�R4u
�����wn9�a�W&��]���d��7h#���*�Ǚ,Mp+���&@�^�GE{�#35�f�Jk�����/�ĻWJ���C������{f�_��N-�Y_w\����ȰIº�7��P^�]LU��Æ�˶�v&8�M쥱���[�ۄ�::D������v�v;�g�Μ<	1m�A���)�{bh
8�e�JbQ.w}+��[�xJ<�Ѱ�sa��*���S��xgf��(�G�}��(�(?����O�1Q�F�[����q�3-���)�h���s�k^\��8�,Ǟ��V�g7��KT��{�/�Nbh�;��B	��ƈ���yK�^���0��?2	@{��2�]T�p��Q+f�V�K/eh���BaJԂ��}x�m"��΃P��3Ҝ�w9������
�d�i
�]ձ�em\����cTA�|׸!���\2�����9M��F�"}|�y�S�W�)*��uG��GVD��u��}s�T}T� �g�p7��Jy��o�x�t����������;X�l�J:����Шv��s��H��EqhC����FM=�h�ͮ�{+��y2���mt�-��BCpY1�tx�-HKl�(�Y�9=�ʕ�a����񍍧
�jzM����v�ٶF1H�ic�C�����40����F�\K{ysϨ�y���߾�Eg��`���WkC�LYj�u�4obI�[�uC\->�|e����ɡ�ƅ.5���t6�e	˗ms�:�+�I���c,]L'*�b�Zc���J�Sjn�ˎ�z���| ������������@��o�t_��o7�-�4�;�'������*_v���Q1��'��nKȻ�q���m��vWR}B�����Xb/l���R�[��ŚTf�o�Z��sʱ��._<KG���H´v��
���U�L�c����4f]󼜞�k����6|P�$f=���J�;�*�����b��U��Z�F�q�W(�H$q �<{�Q��O�2G�:���/[-�]Y������^��5=��*А�sW���ޛ�@�.�I.�N�bM�>���0�#�5Vc�/qrB���	���(�^J��s�4��n��3�z�;���B�,j���
m��d�!N��� ����L>VE��Y����z�����s��yq/��M�s��j����c0AOWY]��&[�oE͞1ч*�S���@.��������"�����
��T/�*}ݲ�.��m�y7��<~n3�c9�WG�Q�K�2YW�#7`s���@c;cU�H�ϱ�-��'���8?�v�a˄�����\'��m,4�*��т�v���Hn����u�A݇���}��-��=M�눟���*4�ӮX�b��J|~�|�JԶ=�t6���O�������F&�e�h�)\�����f�Y�uL��hf7\���%�P[f�DȲ���]n�G���#����a���YU����#5����u�Z�����y��s.�k�@A{�=zb�N�Ovw��
ו�g��ŝ0�s���ܙK��2v���G��gk{
h$Cbv܆�a]vڊ�uo�<s��Lcp@�Œ�:1���S�J��T��;B���nwk�ot�ͼ�C%N��\�Đus��tZ�XˎY�6X�����̴��w�P���>@�<���� �S���I������n�7�:^8�����h�\d�9RU��3/A�`Ǽ�)��O+��!��e�6�e���[x�(��Z��w;J�7�4iNΓ��0^ 5>���䕀�"t�lΦ��z|�Ko˦�?wIV����{Y�w�O�.�1m7�e���cS��-���E��{�A��K:��iΠ�&�2�8��ۏ7�/�2��ԏU����\����|�p�:|�|&���4A�~	�#��җ��Y��t*p�֜�9��җj�L+���ed�y4G�ŝ[��,�8�4Ƕ�"M���=r��C	_��x��4�P1-�rJ��>rS�g��i��l�;%���w>�31�SI��-����T�b}��fSÍ��ݰ�S	c���:!�t�"Jǵ.�f�v���r�������j<�㎮����n)ņ�6͍p�+�z��{������Q� �0�<w��Pf���{4����G>mt���3��D鸔���� ,vT��)��;
mK:z�J���VI�z����$�	�t/�Gx�<��0#�=V���g��{��7p�de�]^l���C@zB�>����������O76I<�Ѹ�{��菬<DN�Y� 롪wg���\�@��]�������8?�a����R�8H0����:'FH[h`��6<Kz�Um��=��C��0w��RR�4��v��h�Vɧ�R�B��#V��	sWE���!<�3��;}$�0!��bHNi��(�	�����/���ϭ8���}��w�b*�[xM��A�X��Ñԯ-.�]��w���ַ;y.HO��-�**W#Ub!��ݝ�N��	K^&���k+ɿ^�WrO��i롷{����A��J
�|02�y�R0�]{��k�%��G���`����`N�
�wV���i�FR�7�28k���f@>�m՘�Ar@���)� 077�h�����I{�`4:b��q�fg�k�X"F4q�"�I��a����)u�����JB��<{}��o�����~?����~�K�̆�����4%�X���Ԗ�h�g����x�~?������~�_���>�f4QP��
4[h
M%i�1U��)��v@}���v�P�IIN�=$i"�۬uu��h�TA�:������Ru�UMPF�CEI��G��n��&��qG�i���4Wx�MATڶ�Y��
tb���g5QOS�#�Rf+F��t�8��*����j)��z �*&�n��ў��tU4�DD�4�QAD�s�(��DU[i�Z(��������T�IQF(�*�V�h�����&�"�hj���z!ӥ��LT�4�3@MTwvA����"j�`�*"�O�@?�?�����ؤ�y��ӂ�Ak��L�W
��kq�����*�2B*f���Ej�r��d�W������OD�����y�Mv��&�w�Ꮫ�7�x�l�@����]r��� �e��.�yUW�z�/c{gX��zRWθ�l������� ��!�n��	���a'�u���S���w9R�~O�k��\�{�vynM�s�6��A��T�-�ޞ�Q��^�J8�Ƙ�.8����5T�-�[c9 ���cdy�G��R#Mw?S��@ƾa ��=x#a��u����PNO��8�#X!��E��VR���me���y3|�[�w� -� �%�Nv�vа a~� 0v2���o�/L�/�]��+Vt�zOPc��ȋ�7v v��06���Y'��h�͜��aeiΫ7�q���c��t�o68���G��(g�ky����ǤA�f#��L�	C�Rh�^t����AEy�ȗ�w�?�l���瓃�����H�)��\Fʊ��V/.���=ǚ]��Zj�&����'M\�h��s�^g���w��X�j+%�:�[�'_n�1��v�jƧ�̾�����|v;d��w��CF�w��o�3���[U��z���y�;ZK�7s�䫋}"�("�U#�5uyx���;�-=c7vl�,�w��z����dr��X�{�A(z��=�&"�������0��9�/�7�;����&�8�[��%��gA\Y�a�eXwj�̹]G�r_�Rt�5+3G��Z�u^=y~��ol��i����$n>�5\���LF`T����S��E�))8�y��[��J/t2�x��͗I�\��!
�\8G�z3a#c�"���&<������L�_��諮�������H8��F@|�O0FǫH��H�R�+�3i�Ṙ�Cq/�yT������(���a���WbSM����g{Cj�X&�0�+1�����ǭ��;�囯�t�F��-��e�jmH����l�Gob8�,�P�<��q�[�����Ɗ���1��őE+��R�R��/`�Is/�1��0��!1jˤ�.G�{n#�� O���;5�<�m-�~f���4��jY���� %𝚩�{��zv�d�z6�/���&��{% ub���i4�ɥ�N�[��	�1�V���7�VLɡ�,�������5��cv�gS��$C^��6��rnOj�{�_�o��`����b��1Ӈ�9�X�8���¸}ƻR4��j����;��	M�̢6�6���ZV�����}+����'��&��f�����=�L�u��f���$n	�����>tY���EZ4km�/�+fuګ��,�x�;�B�s(�:'Z���Y������M�	�L�}2�revӭ��r�H��M ����������dp��B�i��j�K��&b�2�+/	K5.p�V��l��"���ge�-�.4@ڤ.�i��Ұ��2��d�i
�IPe�*Rp�գ���*���D]�����ݒU����	��N��^�]#�#L.�%.m��^������q�ʺ6�}����M]��J�=�"�}�{�%��:�l�V�Z�j�OT�y���E��>"��ttv)�z������c���ڃܴ���$��\y�����Mւ�WS���� Y2�y?D�����W�m���1J�V�v�
�ٻ3�����{��{ݴ�04��d2f��U�0������ }�>��<����_��'��y���N�0)�����0+�gÁ�� L]���w��N��(�h�-n�mt�-��B[����%���d2���^�:�L�����ɮ���+_L�Iw ��H�{����ӗ�A��=W�*3S`� >�ͥ�Wvqʮ(���y��-k�a��2%��#����D�
�8[�F�����]y-����D��5�Ե��������dm'2|�Ba�# C6]gJ�жG>,ȳ�b��e�u5V��嘆gA��`g3�G3���f}]�E�}�����:��MC#G��E{�w��Qћ�@6K{�e��j�Vֹt`M�8�}1�b冠���1�����R���%����SǺ0KO�gqS+n���i�ǔkK`�.���^���{�Q=�qT�6�޼�#b��@%Cd�A�[j~���O#����`��È�{ۛD�㎋�n�0�a ��q �>R�OO�'�j�:���Қn-��F�:�����>��?��`g�i%&�mxrS)������8}�j�M6��M�fޡ�������{�7�Ҏ!�Ų�v�Å�p.�O\Ӆ=���:���h�n��sa���F�l��wǞT��e�PW�{��6Mz�1q5�U�>�7��<�-��3��P��~2r��#�A�
�?]�<7��k!W��jvpi�n��c�]��\f��P��VU�Y�@&�oEFe��6j&��nu�;b�u�t]8n���c�$��"Q��RUA��uө\@7y�
F��y��Xܷ�f�k7�b@���hzJWθ�E�x�\zζ����q�`ï]]�K����
<��t6�l)�4
�TP�K�����|�dA�SbZ:�4niП�in��C���w[�7��v)�Er�^�����3�ÍT֛T6�l�4w�έxN�mt8f���2"1O�@5���N:���mًTY-/�ݳy�� �ʅS�,3�^��
7���0����\
a��\M+�f�-9YZt{������@2�섮=��u[��۬���Z�sժ�mjI�L�2�"Ż}�q�b�쮑8�[Qx��!+�j�7�3��74���B�
��k��j��r8p����t :#6w�ϯ��	'�鞧�g�_�e*O�+�uP��d�f�m��m�ճ�JS�x��X�n�*�P�M�nrG�-����;���x�d��lvZ�Íwf�1�����
��qq@�
�#a��^g���,���Y�1��i�8��tN�=��A5L&yd`���ȸ-��P��g*��Hׯ:��w
!�����(�79}���s�/(�Z*��Q����qWuB�=��5<�̨.���.]CNc����T|/}�<�²�u��,�����G����[�J�~���Wk�J����y����U��:yG"�4��ED����W^��8���r�v���T�x��*�Dr
�"����h�Tz�@�z��m6�����*Y��mc�+x�Z�s�i�ދ��ư�)+/�� c�S�.��B��v1���	y��2�3d+�d���Hs�!X��V�k�ts�W4��U
���;�M���wZ/��x��;j`@��j����'f��c�򏎑��շ����h�N.���/f��]��M�Gz����Qq� �2�M"�9ٿ�LP<��&k��O��!Bbf�����U��C;�;�z"��z��ĳHUx3WT}{ڮ�^�d��� p��}���|rt*�W�
�gm�����9}�S���FC��l
�*���}%8ަ����߯D���ow��iz[�Ȫ��@�n�к��tVE�OT U�>�[n����V���葶\bP�/��ʆq��7�$>����u�����U[���wLf��V[Ǖ.�*�6U���`�e�CEZ��ׁ�m�i���;�=Vd��g*N��{ac�=ԮWB���1M��-��miv�6�Gϡly�,T�r�H��8}�3@���'/��c�;[2�jQ��۹���R�l1��&|��_P��
������f���jh�c�j�j�YG�1�Np� _E��¢�}�F�Z�#�*9y(��Չ���ϖ���'�	�D�ח��!fޒ="��n�\���H��"#q��5 �܀5`e}9�cYT;��.�/	��������.���ӛ6<���:����+&��p�����<���ֳ(U���Rw�n_?b
̤=�՝��e@���I�ZELb�Mqڥ��y �r�O����F������n��n[|���ÄR����I`+V��y
��������F�`�h���Ee�Kl����}��>�觕�Q���С4�0�j�f�#QNǄ��zB��#�?�b;HXy$B�*�����7S[�����o��"��U��q�7.HՄe�������^���6GT�fV3a�;Щ\�Ux>W m1�j��	�ꔯ�Fz_�=u72w����ϜY�C+��8�Tk���N���譎�
>��T��z3	g��A�hޒU�U�ɛ[��]!�h�A-��F���B���Yۛ��3��!{�t�xV��:��~�M���e���b���CsZ�74���Z�ò�.d�3o�p���.���!�t�}�XSK�BY�(ήа��l3���w�G_��a�[��K�)�Lj~�Ͽ{�ǌ����đ�5K�8�N�����s�� $0��A�	�*��n�\�v:�:�Fn��l���a��l�:�է���J�j������V�O����1[��)f��z��.',w�6��'�4�AV�!0�1M̜��A���Ue�S��c�˖��.�9�N���Aj�5�d�;:�im󷫭jSh�ѯ�{����v߫��~�|�T��Ȏ�ۜ���B0;%�7ip�v���9�f����I��>����Ӆ���m�ѽ�{�5{�|:��"�:afdK�l�{�4�q�s笃��׍���A �s�	7�OӐ�+dN7��h����C#��ETUʡz�uѺOp*�D��+!c){�&g۬�7շ}�lXk�0���p�C��T��Ge�@\��Cw����n���=θ��,�MЅV6��諊y���r����	�(�����6��x�	��{:�Ld�wk� U�ϻ����s4�*�
� A�]����-��]-׻��9/r�JP�lu�4F�uWa����C(#&"C�ힷpڡe"�t�k���&��F�J����u�.��'Hg�GP���T5�>}8��͋�E ]^�(����+�R�fD?X��扖}�s� �:\J��H�L:g~�6j�7}���}d�*K{��D�-�E&� ؠ�* b��@t�]-�`�k��'|�2�]_]v��rv���|8�f����˝*M<�)v�Ks+#m�����}NU�{IaX��D�����<�'ph��k�\�Bۂۅ���y��"�=ZJ�R�&�y�7�#U�9���ݚc�߈;*In���vXP/���^6P��q֠�"NK[��A&�y�d��ղ�yv6�Ͷ���4�3
{ ��<�\��$w��jC^nd�~�qu3t��؀F�8(�爜��i�j�����x�#*��}+����r�;�vH���_���r��6�է�V�Y�0uvoP��,�9\��1eR3��1ǧ�s
�"��/���9lj��������~��%�۠gY��ֳ��2�m.��޵w3�c`�B�/o���+�E�����	K�i���n�w�����P��uQp�%KgWn�*�x�.���ng����B�]��59y��Ug]�MӍ*�!���v�>� ω�$&���ndj��ލ��~�������{#��*����DD���?�?�[�� 
A�}�b���`aXa �!�a�a@�P!�`eB@�U�P!�aXe@�@!�`a@�!�a�d��P!�@�@!�a@�!�eaB@��a� !��C C��2�0!�0��C#�0�0�0���0�00�2##��#��#� ��� � �� ����0�0�0ʰ�0�0�0Ȱ�0�020�0,2202�0,�]z���2 0�>� P@PP�G C
 C  C
 C �C  C" C
 C C" u�@� (�((�4� � .!� &�Pi� !� &�Pi� !�@!�@!� :�z ��i�&&T@�&DF�Df&Ea�Y�Ev\��Ȍ�Ȭ0#4��2��C3LL̂M0��]�	�C"�r!�U�P!�a�eXa�!�a@�!�aV@�?����׸1��?�DI� � d��}���>���˳��������������������u�6���;������?�QU����_�O�}xʊ��{0����� d�O��S��?ȇ�
*��������������H���O��_���y���!���X�рDXAJU@ZEP�ܐ� h@ 	� " �@� "D �@	� $! a  @	P�  HFQ@�	B%H@�aBE�	$VT�	@�!V$ @$aI@�V@���������O�DDAiA�@(
�ǂo��������������y�0TW����߯����������v��v��O��}c�?$���訪��a����_�;�S�EU�QETW���C�?<B���_�~�װ�UQ_@@g�����}��{��<������?1��?�����QU�b�����**�����������C����`�ϡ�� ��O�����8U������Z��+� �������)?U�y�ӣ���ggA������{��<�$��zTUE}'��~|?rd���>A�?������\
(
�����^�����g��w����2�?�1AY&SY�r#T8Y�pP��3'� b6�����Q@z�C�A`����))J��L��+CT&ک�TUdٴ��j��ښQT��Y@SLUA**QIH�+Z�Y>��ʩ�Q���)���kFjյ�f̱���4����Z��m�i[TmCm�V�-��5��[0��ѭe��[l�:�K��ۺ�[5,ٓm�jٲ��VM��R�4K&�4U�ͩh�&�a��̫#jF�E*m��!��m�L`mm�e�!If�e	[m5���l�dU���6�,��.  j��2hS4�A��z6�Q[Mk}�iyp��{����Wn��C���t [t�N�t�hdw����봻��8��顧uֻMۡmC��V�l�uv�e�E-�Jm��[�  -�B�
(P�������B����Рx���>�(44(P���p�>����k�k�s�kf���ٺ��C�։�n�Ҫ���+���S�{sm�5��{���J��oZw���tr]��h��v�+cMg� �ж�n�ܺ��:mK�iښ�wnnK��:V�t�+iv��k���}��ڞs�q����N��oZ�@t�75һ5l�ڥ��͠u��[��MiX��lB�kZl��| ��a]IN���v���c4;�WU�[��m�wJ��m�{;�Wt��tk����ԷNs�*��v�:��N�ҵ�ū��lh�v�kKej5���@���6ڴ� \w��v��*�͵+k[j*Y�Ε���\��C����Y��m%��;��[:mݵݭU+�;w&�D�C��*�b�TQ�+cjU^z���k����:�)�;�� ��uP q�qAEl��Q�]]���w
���wuYAJ�]F��.Z�[U�6�jkVaXE&�|=Cց.�P�iݭ���K��:�[\��}���w )R�w�y���^��yHUH^=���
R��nz�)J O9�+cdcCŦٶ���	���J#��l�Ky�x��*^��QW`5��q���N�(��)s�qJ��L����*�z�`t
Hѝ( x�m�A�V�����3aV��� ���*{�gy*EQ�+t�ĠQF��<��Q%�e7n)/{���;OoQ�Ij��EJy�7����5�볏E(U4�H��R���͵�j�Z�)_  �}�
�Q}����4�����R��L�L�){2�S��R�݆���8J�w��J�������j�N:qВ�Gz��UUIU> E? 2��@4@��0�)P  �JR�  )�CIJ� @T��fUR�� h B�4��  b~?g�??���j����};����`���.��������z��;�?G�f�o^~����"���]{��E DW�UE?��"+�� ���PEaUE:���=�?�a '�u���f��S�>p��Eeςm���fһ�c^�&�dy!f�Kn�e�I�[J]�N�ό٥^7�+o-����U �CP \X�Ѽ�/̂Y�V�Z��u������:#���Ǌ��-z� hQ�C��L���Q�0ңy��U��ӧa�!%B�H�-���D7��d�$T��oK��ܙ6(g��9�6�d5�s�ua�VrZT7n��/T��#)�-V� �e�������7u�.k����ԴV�҈��&�;�%��*��Kws]���(in+If�7]h[�B�$2͊��KK B` ���v��{Y8iX��2�]9`RܩV�e10�(퓔v�R�
�.�Kb�k1őy��aur���Yn���\ͽ��\�cc^�z)��1	���f�_ ��бhW#(��G3I�ojl;ni�h��)�ޒ3]C��#l�9�ZՓ2�vY܍֍�krT�f?��N�3�4����) ?��H�Ki���7[���ov�h�4�R�h�4��cX@���xƑb�n��^��
S�ؔEe�.�M�d9��lc^�S��Ih ��Fvb��ˊ��m�	�l���6S�4��V,	^��v0eYb��I��,���Bǻ� �gLk�ҵ�
��(��
^ 9�edWy��xn���dm�$�w�u�v���Q��r/� ��Ab�DK��0P��]@���,��Pz��5�a��E_�T��@�����u4�m���#۲f,�J)A��� �<�Qh:1Y�7�J�T��"31_�Cn���V5QkZ����q��nf^��by��nf��oq���Z�)�NKB�%Q��U%ꉉ�Y��*	j�	��џ^Z�j�[��f�/j�`)ݥaIf[��&�ڹ:j��dAV:�����Z�V�/q��j�Պ�uj*�*�A;L�5ͨ /UM*ۊ�ё`gZz�l�K���ib
�姯��kcd��)9���0��+I�BZ#��c�&c	K�楻����o�ݛ�CS�*�	��Z�ǭ$/T�,�F �n�����z޽�܉�����V�n�LY��p��dH��:k�MXF͎��`z����:VF(-�������� c�#6L;L�P�[��mՒ�������P,�$���&LL˛����wY��᪛0�FIMnK��5�J#P{AQC��`�I�%�c���Н͹Cm0��h9�Aқjκ��Ԡ�x-�oW��!�\�t�`P��=�ֆF���Y�2�zڱx6�hlYR��{6�mf��lf�[Oo��2����l�N�w�S����v�������=��� vQ�P�*�q*�hʕ/!�Z�Z�zL�݊�,��E�V����E�72�{ź2���'��I�Ҵ;�6����8�c^ބ�^����0j)*�2j���ۢ7�����u�����/]  ����puL��&�|�E�Pl ˵��rn*������X�I&�ֵ�ɥA�&�:��Xf�4�k�,r\��j6A���|���M��Va��[�XqJɸ���b׏-
���ۑ	p�K6�ieHո�v�r���+�Re^K�Ze�V��.<n�����l�߱���d�7Nރ(���͹y>�p��;m�1���W��7x�x����mMTb���d$yJm ��qI�Lܸӎ;�ܫ+ ��,��5]Xjb�jn�2��n
F���K7v�/Ll���bH�Ԟ��5e+���-������i�7�JAN�ix-\��R���m��Y�b2�f����v��ʖ@�wB��*B��1�RnE���]�
;yj�ꬒ%	6=�7oEޫ{�K�զ~�e:�u/�ѣ f�e2�f����� �#�Z�[�&��#�!���IRe��=r��ZtR��Xz&m-���أY�W�s#�.�ږ`���<���u���VR�L�vR%�"��)4��0�t[�e0��ٖ��#ӭ��j�DV0��E�R䛊=[��:���'��L扺�9f�J�+5$YB����^�bKNVi]Z�rTZHg�.�Utӕ
J�s]�[�å�T��36��7VA���y��&�f��{
[�3j���lEQ���D�	&)l��9���,��נe�1��231�)�i��6ԫ�y��NU���:t��xe���H�@hhmJ[!Ia��R��4ne��ds
o(X$��ʋ ڛ�^*{�����,
�%����j�R�l����4�$�r���i䗮�TD+Fi$�P�"F��<^��]v���s:��/�QHD�C��9�I?k�%=�oi��ʛgN̙%����J�̍�*k�VU���ˀ�v*ђ��n��2����:,S�ݚY2�˟77-M�M҉5)���8�I��ܻ%����m�M�!$7Ld���ӺR5�P�f�P�e]�1#�</)��-��\2��%q�hv��=�F���(�P�ٸ.�u����b!��gQSȶiR��5c®[�@`�Gk++kN6��$V2���Q6^Ұ��*c�&��x"�V�4JN�^)�1�G*,ɑ�����%x���쐐��J��zd<���LTP�UB��V뤨�K�к5($�Q�#G������Қ���++l��*|^qtB��ʼ��7�G
5��͋��v��+(͸m�賁�^�+�0 h[�r���;��/ظL�u)'I��{u�^M� Be��G�P������VK�{Ir�ƂC��;�t@fo��koa�cn�.�������K<�x���7+1P�d~�F[�/@UiRZ;�%R����G&�*�`��He�AYp0�B�"�1�BM�w]��<�;Fl��.]Ŷ�'-�i�pPe���<V��"YP&
P��$�*UB-�?/�N��*n�����K�j.ޚ*Rof����!^���#su3>��+X��4%+��Ν�LǴ�s�٦�~�<����@�(�)�$ɣoi���)X��i�VB�l��blV����	�!k���D��B"⧠�R�ɉ6�Q�-��d0�͉޻7x����%��*�\��܆]̎�����㧛)�3����䫊TӺ��l ����4A�1��us�O�#��6�}�z��X� ,��7i�" ]j���N
Vh2X�(�6�'yI���QU�&�93P���<wQi��DɤVlV\���
��ja�1���.���V�q=�j��;�#�ieV�2��0�Sq�̜uO0Ji�2�/U-N��)H����V̌��,"��,ֻ�cU+Vk
N�ʑ�,��u.L�w�v�@�e�	�������1%<{C1�H�>Ǯ�J�Uifun�^�r��j0�O/�T�x�:��69&�
Y�P�u��{qd��8�������f�`
���r��ܓb�7��Ѥ����2��yW�1�4�m�L��k-� 3 �i9�ͱs"��E����e
�ԛ&�fV���ņ\��HB��"�Z�-Wx��t *Ѧ�VVM��J����`��eܬ��#M�v�9J��[�N�w��8k�B�X��*��%.�Ga�͈�r)����1�*�j��s�@0N޷GE����B���wM�ajԋ�V��N�����s"i9�᳔���Y��@(�ܥB�]�`��Ȫi#t�FK,V�3*Bբ�.�n���.f�t�9���덓�`�E�l�U��)�+��kv��M�4�HڦD��E��jkpRkoF�e�+�['70�YU�Pt�,���Ղ��`WW�[��l35^[5� D按=F���Fhe:Ո��I���,�(0�ϓt�1�$hb�x)G�k[/.-��y1T�e-�R^T�z���rT8���Nf�n�1���v�LTX������f�)]������%w�l(�0����mn�����Ӽ4�:��^�١�r�� �Hr���kBw&����_ �H}w��*�Ye�$aBۻ&�%X� ��Vb���h�X��t#�sP�������2�[�K�W��M+N�tc�#ueV=0�6��Wy�얠�c��J�M�N�W��ϲ�Ò��lҦ)����u2q�b��{������2k���bn:�e�`����gM�� ���u�������.�I��6��6��H���_tI�P+�n+q��u2��yp�Xfk��v[��wfI�Kd=��Шq��!�7&;�UmK!	0¢QY�V�a�9�s&Xq���ӈ��ݬ�VV�:�TmP(��k��L��mn;x���ݬ,廂��Y�+ص�b�q7�v��ʭq��ZHiK��%7�*�K*�;:soh��-��չ��R�1CWeP�1fʦ�m=�Ow6���rf�΄L�J衺o�$�\)뱂�(��cS2n�ڼT쿬�mb�*�BQ�؆Ӊ�۬�*�R�jܫ"'.�&2�gX�������i�I���LV�Q��m�( �C^����^�4k0V0�ʫ�
֬��g�U��v��Vj�f�PTNm?��n9W��u��9�ky���Sk�m���+u�<�&
Uz���P��ƚZ�c���]�(e�f���Ď�(�Q�Wz+ %���	)�t���*��{k�l����5��)0���r���Ag���N��n�CIr0����sZY`HM�M���CJZ�Y4F<|$u�\/�"��鱌
b� ��4)�n����0naA�ycC0�*��u�W�5�S��n�q�J*ĨZAT&R�PY�+He�r
���T.�iW���K&<iU�k�%mHϘ�he
�p�9w��b��V��E`���&[0j�n�]��*=5�I۫��r�B����O.&��e mkp���`,��G��u�d����d�2L��ͧ`����Q���)�`jY��tS���%�P;���ס�-�:Ӧ6��f��Ka0o0�����,Q���KHϙbK�[���b7�}�޽�{a�$��WJ�!��%���;"%�����0���K�͔)ӎ�ծ�L�ZV�⻭�^�$Dٺ���Zջcp�!�$Ј�E�8��ݚ[H����d�"uhٙ�2�dxh�p�CN�)��+t�&]�@\��7r���a%�5^����΍���X��t<z�#5�KL���q�$�w`k�����k�7F���|��+(s�`�����Z�:2"�[/f���+Kذ�]��$�ʬ۱��G����P�#XJ�L�9re�պ���m�!��$�K��W��t4���Wa-kt��qAy2�Œ��*Eu�R�I�(J���qV�X�Ev���Uj2�˄��-`(ҷ{�q��bb�3[f
�pŮ�Q �έ��鵰e�m���0����]&幉V��-�C������Yf��b�к,;�yWQt�0����S)�J�n3.] �7�J6�[�i9������b�������Ĭ;�A���(��y��n���i��J{W�"��jh-�U2c�5���ˇfl0�4�r�Wu̶F6Q
@]BQ�ɶ��x����	�=KV)[�m�1�����o�a�+^7h\�Q��1�2��>���պb]b�i�r�Q7���k��b�p3��Vܠ�5�����j���D���cTb�kb����B:���w��D��u�`��$q��F	��r��8���7iY��IC@:H�{ne�%�+���l:Y�,'C�d�n��*�[OT���7�n:�x���Z-�e>�_2���,��U`ZC����v,N�VT��@�ڸ���0R3ʆ��ŝcjG��S�X\���3-�cI���h�ѹ��U���I��[e�lF��dR;�Fn ��Z��`٘�Al��݌ n)��.���nl�.�)e�iz���,00&�ڶ#xP_+��1����Q�A���=B��B�)���p�z6����v�e,����i�q`ج֍��U�F��(I�TQ����l,�V��d&n2mlB�{�����u���ǳN�9A����$�yy\Z�7�e7sdu�1(���ۺ�!����.*9�Ay�[�V����iG#��J�����X&�i8�]�d Z�z7Q@�C2m:6>�aX�[�3C�Х�)�ai��8�5,�X�6BX{��r�c5A����%�xl�BH��#B��,)V[7J8��6h�[1�(��4۱�U�!��,�J�%5��E�2���wu��-\Y�4�E<�d��J� iRX�m�fȂ+aP���D��ai���BJ��1e��R�7W#�Đ�x�d�o��%�)���t�����h�w�.((�W��'j��k(4]'m}R�O��*R��Z�A��0� '�j ����7���X�Y�T�r�GV����U1EM�R���YF�;�����\�Et��A�[���tl:$��2٦,�×�":j��U���w����']m-z�m	ic�t���X1�X/a�&�V��EU�0U��ʦ�ɲ����s*se�7BJ)Bg5i�3Qq��5Ru���ϐ�Z0 1=Z"K�dC��M�N�\��:O� 5ա�t�kp;!�6�<�v5b��dwcRt��1�I+a�� *��Vf Ӣ���Y��`H1��Y%\�-JifʗZ�^擆��ӏ(�S��#.���2C��n���� �[Ku�Ӫ )ưd�#��l�̛��lP��ZH{z���to�з��S�^�%@6��d�)ϣ����\�j9)������'�u���o��l!|���^�9��;��W(��^*�BU�r�*9d�|�J ����<�k\ŗӁ��vfXӭVUl`�b��&kbv֎��h�
�C��u���⫺"YY;EZ��5x7���A{��fֻ��s�L�)Xr�0�A�yw7�u�Rb�Y��U�k4XX��o�b�U�cp�Ӭ_9���G�3F:�g4��o�5}�I�34n��4�\E%�@��ڮ�mp���K8V�,��^cz��a����Z�v�y����B�t���C1Ѵ2�dR���H�z���Q�Fk��\Ӿ�"a5l��j���5L]�0�9c{�m�t���H��Ɂ:=HdܓMr�,�x�l�.E�^���m�s�o��P��h��0�V��ҥ(
�{�b�JD<o�!�/�V����u��H�2��Jjp���;�l�Vm�y�yV��J�N'��d�5C�K6��A-	r��AŸ-���R��^��5.���C�{@7;i�K����UiRWSAڏ�U�p�j�X-p�X^=��,�ǵ���7����,.׸�]����u���J��['m��Tn�(^C�T��@/�y��R�{�e2��G.��l��o+\X��������w��U�[�dqm�P|ǻ��J�+��nZvrv��R�*p�5ܵ��o)J�}[J�7���'���l�ߜ��d<�܁�&�)��OR���Z�/8luM�Q�w�~�wa�&�7o7V�y#�TՂ��HG$��ޣ3��B��e�2�T�&�xh�n��T1>�9A���0c���/���%$.��Z�mr��Y�:�,eJ�o��,v`��"e^��|��U��/�65`+��tyq�I�i]Ak�HRp1I�q���ub��i�}�,�/�љ�Tz+�>��$Rˠw	�Z�v#��Nc&��.6	Z��nv]��}�7�$���S�9��_9e�1;��Jߘ]�M�oHǢ蹉(�Y�><^���Y�����!t����"��}�����^E[�Wp�sSX�R�����,v��wMO�Z&�x����l[��^�Gt@��jݩ�R�خ��S�+$q���TN���U(�wH,��K�Up>����Y�aS'ef��U�o�%���+$�kT�fm#s��X:����xQT��L�Ȇ�v�Q7�]bz8`;N�ȇ1�"-���!l�n��O3(�*�A�݈�\��0iz�k�l[�E9�>*�Uӥwb��g;S��[�y�odu)�h��(Vf*�]�t�j�]@�]6gV��ai%F(�ˎ�潝�N�떨�"��i�y�/`���B��i��1��;��>4�ؠ�����8��!�N�V�:�����xj�t.��4EA��h�iPv&;�qN����K�,��͖a��)�T�Z��m������G��l����f�(�;;� f�Sv�|RW5��0�~ح�Q��a�D�q>��(���'�[�{Ųm��s2��Ⱥ�c4V�������`ݨ6��O;6/��.�� o	�r���'S�᭹�m]Ԝ�R�,�
�﫯���wP�1��ՒPT�Ѵ5U��&��k�c�]��&;j�ģ�lpz�z���+R���<E�}���7(���*v��j'Ϯ�t��ڻk緱#�J����/-a��1C��s����y8��8m9��xb�h�t�3�Ȁz��i����_f�*���m��,�t���ӫGo)�v����GnhC}����+��gr:�[�&WQ]�Y�`���� M	M��d5�)��fd!�ý Ʈ�, 8±�72������7C��y7g�V;�mE�A.Ƿ�M��.��
;X��]��B�q�7��pN�A!vB��Z����7���#V���O��	��V��Ū��,��I|�h�4��:IX�x�����~��mʹ-� �C<�*��Ne��s5zS\���rd�z�t֕6�-<�:rj��=sTO��S/w����ۭ�x�Ng�F��g�m�"&V^ec;rb�0Z�K��7��\'���[�R�p����lor���J|Ʒoi�/����r�٥݊��u
���nR�
���lu�%���әbGG+��Ep��3���=�bVLC%藝�^�zR��H\눡6�S�� \[Rf6L�Oz�]sEJ+��z��!��RŴէ�3]��ShZ#�0���p��C[�o0����c�Ϲ���fᴲtR�S��R3h��8��j�����|����?90�o�v����H�'���dR�8:�ԺZ�T�+cܔ$�O��w`ү'>8o�Y�'��K�ݫ��G2,V�d�Ȝ{O�B�Iuѳ>Ў�}�;�tc�Ģ~��sF6����l������4kX]ҕ��ʾ�6��$\�u�JAa���S��Y��]S��9e�Gv�W����u�]2�ۛER�Z0h�7�sXq� e�q��Ȃ��Zۙ�e��E>w&��lm�)!���iT��<Z]]�.�;d�j�\�����F�z3鮔�_D��H�i�Y����5p!˴��<��`j�lL(�@ύ�~9����c&���5���s�"mH��GV�s%�@肶-!X�R�'da|k��Z="���X��]�����*�T����E�V���ya=(A��c�[|W��Y���T5.�L\���X�&�Yl�e^��a����S��I|j�ָ��H�+���F����qNΦ��c��s��Sn��7��k�%�ou]I�Z;iٜu�P#B����1w��~I�5ԣ1-̺5y�a�v�,�\(^���oZ7j��ѣ�-أ��p�2+jQ��T{e-qp{��R���"j햬���].�0�.����0���__:�DJ΀�r��V�5���)��7§M�ЩN+�Y��I{ۣ�����)�����B��Z[1�+�h�Ы�{��;K�y�Zkh&��ʎ���J�
����j*��5gV6�����������{�[�m:D}�D�g@���Kv�L�l�t�n㽟n�ݽBNG={@&��[��]��r���@XX�Ȇ��L�,��opx1LHd��*n�T���X�#�A�j;Ql��E��nl:S��Uµ���BK��~B��o�j��o\�}NFl�	#��q4p<:/J�
��,���L�H��e۽>�[�	q��$���{)�\kK�V\����J�I�ܓ0\��cӶ��d�9�Q�]�\;��7M���Å��n� ��\�%zS'����n�Pe��U�w��p��)���̼��WxJ���;���\���C
k�m���gٻpւRy�a�qN���1)Sj�uXQn�ҵe�e������&gl���t�,�\�ƖvF�X��g�2�fi5tHv��@N>��l����#A:L�S��ޙ�vS�ڵ�\�d[��\�i���#o{x�Ȳ�a�:��0\��\2��-�s�@��q�^q	�.��D_@E_ ��O=�*>�c}y�CI1W(��j�J��S©�Wx��q�J�-k�0�E�2�F��&be:�Yy�a��e�%�̕��q��U`��Uր��n�W�FV�˃r�N�'���e�7kr�p'��4Rv䮡� �R˳�]�^s�7�T���NR��_z��Z�YҰ�q��̇(����<餉��S�1
D��,ն�4T�����\sA�����P�`MV�\���>Y7����r����\Br\��t�u'z���o�C`�t���եa��.(���y�L�w����fk4�
֞����	�A�sk��f9����(S7)�3t�8���Y�|ZA9�AY.`]�N4�����v0X�E���1�D��#���޼Z�tU4,��iJ\�5ٶ
�� VpU�]_�^���KtwCco�����Jbܜ��i��Ƿ�WTX �ٖ�"������s1��o%:��J�E���3S����&7a�K:\�M���w]ݍ*����n.�x�J���m椨���9+k��C�Z]f�]�Ú���qtZ$)֧ī�v0~�K20��bZ�ɷ����H�z��i�˷�hhS5Z�Z2��Σ.�]]R@Z��
u�0R4W3�¤���
����ãbم
7��l��ۘuA��S���Qw�����D+Y�F���{(���ܯ)3P<��LyC9��[�����P+T+&��UG� �**�%R5R�;�����I
�����dB�n�V��I|�qN�g��y}A�h�H����^\ж����s�q<�[��-�9�1K���� i��m����U� &o9�﹅*'2�I�-Z�Hj!��mpς�Q�4�=V�X�}�.��R,�E҂~x�f��f/Xj�y���7攈���A��m���Aŉ����`��;�'`�'E]�}X;1ݴ�;Y1��&�Oh���E�@�i_IW+`.1]C>3�c���Nt��b��u.]�6H]�6�r8��z�1|�]'u�C�9}��ta�45������������	*`O�U�^S98�Ⱦ�U�8_j/�)Xʄ�̼��[��7�d+���`�����Ļ׊����$��eH�)��K%U�Z������9�G���J
��܌*��p󐵠4]������V�ܥ��:*����e)L�a���e�ޡ|Y=�U�ԥ�# rs	��홓��9jdN�����4Z*��E�~z���ۨ�ƚ�[+Ȳ�������L��m!Y:��u��a���K����c�TS��˽��ۧF\���������ԉN�b.���b{w���B���H����%cՔ'up��)�B��TYg�j�+����s��sd�ǘ/Q���l(�^S���Jp��y��\�Cr1F�l痕f��ۭTk�gK���J̤�n�9y@̎��rc,��;�X4x�v�Ϟi��핚]�|KP֊I:x����iV��wm�0a]�{������*�s�ٗ|:`R윑=�f�xZD",<,¾r��dI�}i��udx��<������>r*y����1����X�i��Y_U�:�!��]�����η�SJJ���n�[P�1�A�Z|�]@� '�* p`���~��k^�'}��w5��k`�fR��n��G�_/.�G*���[�Q9,��v<p�L�QV�������6"�uz��/�q۴	��Y�m'�vJ�ʮC5�+s�p����=�6n�mӂ=�#�����s�e���������E���8g�)��'e�>�k��ʫ1ip���":�L����X]�n���.�Yu��"ݫ���4��P��/�=��:�����ݝ��Y�u�����G�P�/���mA�.�fʰ&�)�i�JZ�:���]諝M0�Q5��M՘��}h�k,�{���[�Ghc������T� |�Sk�m^�����Mv��=6��[�v��Ln?+%F���B��-�P�	[���7�9Y�;*���/v��u��K�-�Tcb	��.5
���WY̘wUc�b�rQ���3��)cF���+9}J	J*ŬV�ɽ�15ܪ��ُ�5Zh/�wG�]C9��\S҉[)*�s,���}�/�2���]8f�lf��%a5�;u!��%*��*���Al�x�u�֯0�Rj�sR3(+�k�l�������^�<�9]�k3$�9��(��Ԋ��]4	Csr�$v�T|����z��n�P��������^Y�@��
/&A�6�YH�AV�쁧�A�qثZ�8 K��
oS��F;��>М�Mau�ry�&�<��,��xI��q����$��e����6�:��E:Y�S������9*��T��nM�yѬ���`:�Q�׋-Z�m9��â��n ��S���x���q�[�֩���.C6S��l�@3� �����tA��<��KT7A��oe!k�H}������9���	�g+Z8�vK�S���nf}pX�X�m��	��y�q{O��v�T+�v�VNE	7�xQ�)�ʀt0.�ү�����fcjl��Y
;AB���ZɻR�9:r��1��9�}�ceb �;��T�ZPp�#�����N� t}�������ǻ23Vc�#ܓ�������+ �z��ΰݤ]&4t�u��n,���#�rh�D�a����4�'Q�����o`�2Rw��mD��2
�ڸs�9���l��Nm�vA�3�놶�p��C�N�Ă�W�E��/�C��/�,Ց�h�LѠ��4�l���x`	 U-��|�Y&`�9u�����ˣxj d9W�tv��P�$E6��7�S��oS|T8�?���Q:�]+��o�M�*<��+S��qV�#n㏾u�e(�&��2��X��޴i��Ս�9��ũ-�xi�C��{��mugJ�mq޺�`�>�;`�f�؜r\u0�"+�鋧.�,9���d��7��٩v��
1�9��ԩ[B��VZ��'�8W���Kr`L�������}:A����ne�F�2���s��M+����*@Ses����`;�P���ֺ1Q�x�>��]Nu� �w[F��i��r����K61u�ɩۀa��b��C���ٚK� �E(ee5�9q�jԑ�}r�)^a6Z4+5r֎L���<�*7I�U6�so�(r$U�5��Sj>�E��f�J5�n�
ɳ(�2�JZ�m҂���0��R���k��V�P-Ꮡ��vu��-��6�^|�	���Ӫ�Zr�Z��:��W#�kcXk.�q2J�'E%��s�k�AU� ���[�>��:�:�]g�W/��sG�u�F�~$�5�	v��i��@S]�`�0�ox+ٷ��=c]�IM#�Q�I�;[A�{FM����bYg�X�oaw�4�����m��ɕ����J�C��&���G�F3�I���*R��vnSE����g�v��+��E.�l.&�r�"��W-��֭lL��fȦX�ڲ�vjц�����6�ܲ�%��wz�N�^��+�M�y%�ڦ�hU�jn�Xll湶5�fF��+���Kٍ�G_3\Ǵh�#bto�a��Y%^���unD��5kX�q�T��fb���t�Kv�m����A���5յ����X��$j�Y\��˚wɺ�l�dá9���;f�pΚEeL�oQ�E=Ȣ�Au�K9��M�PX����]˫&��@���H�e*�9��N��5��:À_	+��Ķ;K��r���t�V��q��0�8�I�tv��\#�c'Eג`_.\1S�����Z�×T�P��b�/��f-��ɗ���T�ғTJ}v�)�\�_Q��:��Wy*rѴ��C�qRC�1[��|;���M�c,f�R鯝sc����ۘ�4wK}YDZ�kS��Ĕh>��`�!���]	[�L��mXR�ԩ/�M��t[nf(�8#�k�E�� *�z�
�t"����Ƥ��z��pUrR]�#���� 8а9Q���@Uv�5��m�Sd7���B���:P����/S�h'F�,+lޥ���Z����.И����Z�LV���S�|bwHCn ��SyR�ko��3���\h�']�2	%��C>UwA[[�DLq�x4�Rf�Y���(�,�H������6����>'�>|�^컛���6%sU�����"��m�C������R.��yY�I��nho��5h���r`��e�wZ6�FK;}�@�ɛ�X�,r�}o{�u�u�T�J5]�y���;B£%���e�%gE>��8�..�m��K�y�&PT���k2�f[��$���(�x��:�L�ٶ^.�xo���eZ�Zc鷺U��K1���Z2��b���W �u����;�{y�ʻ8��y�K�!Y}J���l�vU��^w�f��c�h��Px�_����T�pd�\����"|iѕ��2n��zĦe�4o�4k] �G_a�fPZgma9�0��R��s��1}�q�Y�_�8��3�
os����Q��XZ8�P���ϕj/���x0���7.�+]����],�7�ˑ�1	�آT��ޫa�З������&����,�x��AQ����t�������H�����iZT����l�O�ۧm���Â��Ǚq�j�F.W�\2u]t���0���Fv�97e�X��t��nrCk�9R� ��g��FPt�h���sCd%b\
=�mFu�9�lWM��m*�h�����-PoKl]:�Y��u�{nJ��z��1W+����.��Ʀi��19)��W΄R�r�@U�oEn@e��y�su�5��	u:�<2��;ά��QEQQ>ڐ�ՇY{ל�/��\��	m�NM bBT2	qV����:�q���)�q;�����E]t�vok���Lh,�ì܎���`)�Һ��RP,*;�t������.1K�+ �xn���q^���a܁�5�q�8v���gv��h�6�����%���U�-��y�RwR�1KX匣��'=�U>c @�.�R|� ����� 9��d7��Qc�F���|�Kg���K�0G6�[u���u���sz�NGhkrd�l�tS��X�L�z�@�����^�W��xu��k�*ne�������l���W��%�̔p��3� ��q̾�k����oT�X�
�g�a��қ���"�2������-��):�ͷh8��j�~�V��7�!�%*4�R��1NT�f�����x���V�qZ�K��p���]�x
�xi0���J�/l��|:��u���7���� �p���Р5B�U��N�sf��ki�J޷��+�jVroe�ïl��msM�Ʊw]۷�V����l*��kJ��z�ș�v6��oE��*�ӥ�s�����_e�L���)�
6���gU*옲[r�ħ.�s�u���0�Os�t���t8�oX�N����!�ik7[���+��?s�SE�~&CE�]�Z[w��Z�`�I��9�)9�ܳj�SS-�Y��0޻,��rၡ!�sp!|�[Ok6�Z�vj��W�&�HU�ji-gZ���yвu��w,��-ӓ^���z�mJ��m_�$��F��{Q�
�Kz0R��Θ�h��'3먀1Rْ�;.�s���,R5h-�S1�������pw���И���++�K������=$��ym��P�s��İz�;41Ƶa��9�a���<t��ͧ��"��Vݥi�
s+z�.���Y)��e혬7���ӯd�� �Q*X�u���kD�G^�N�C&*4&
i�b��X��A�٬��4��4���륶��4"ژY�k�(e�VL��� ����c��5�}���f��V�arE�d�<�����V���N��BW����6�,��\�8��k���D޽[|2	9欚l%��vKTN�d|�b�m����c��g��e.ى޿��m�[�Iw�.L��R�]1�����y@l�&�ם�2.5�:��N�k{L�me-�:�7#�]���6]c7I��|5�p�l6,^���Iƙa�D���<�n��G&��F���+ċ��J�a�ł^��4`{B���ig4rS�/�7��{�m�V�wIQ��ge��75qiP,����9j�j�`�C�y����DT�n��M�l
D䭔l��WI*P�J�����+hdZh޾-;���6��ԍ��b�7}3�nP�HI.m�eB0�3��k\�yH�]�Vv�������%f�f��g*�-q��f0,˒���
K�km����g)�$�AU�<i!gv��c�do�4��a��ք���@(VYG��.t�Oy�\�7��4����>pJ��mva�8!Vل��2�q6����w9�'F��K]�.-�t�I�vKc���V�%�,�s�B&��Lk#Ů9�$ 2.�x:�%���-º��	��R����#b�u3��W<��8���)��ڷP|� k[���}p����Wy�"�aw�{�@N[�n�T��w������(:�+z�,�CWDY��:��T;ff2�N���^��v�d��� gp����V�����ٗ����5}��=�����#֊=����e��W�D�t0�:>����^��W:��1�����N�c��J�����=��(ӷ]n!K�N�P�
�EA�B�S��t�ۮ�\��*�)Y]b��3u�kQ4�*���S�*+9�U�:s5v�+!Uw1�}N�
��)�J�ϐ�C�Ɩ�w
�v~�.آ\w�ǝ�2��cY�մ*>l���+;��Oa�:/Qh=%3hJ�0(h�5�d/ ��,e����6�Ѭv�8zU�Y��wo�P���y+��h_+#;.��=�	c�h�u�R��Y�7,ʥ|���BqpKD3R"C��]�2﹡H�����EZ��ޫ����]@��+����@���v7w.VW��JZ�[���C%�ǐ��gj�IE�%��DKNc��*W֫Ó)�ksS[x���Gb�~�{�8����)�q��n8�X|�m��:��2Y��)�T;�չ�>�*�J�/ ��T��U�ͧ�kn\�bJ�Аb�ͮ��
4��A/k62,\T��^ѝxH7���Y�Ѭ���͕�[D���cY�ʧL�y+}rݤ"�Fr1ٸ-B�)I��򔞜bp	��Ν"�
��;N�ia���uv`/!'`�cY�4��{2�uZ�g	���7�)۸k��vh=���!n�-;��,�@��R���*
j[�����)�	��sR��5 ���"�,�u:�R�gK�k�\g2RA�q7��
ͼ���Y�wzg��)�i�üp�A���K�,Ŷp���Q��Dڊk�a����7�����=�bPX�0�"��%ژ�,t��hr�*eɅvl�`HeZ���%g��� �Ι}�����V�6;L���Ɛ��r#{���1���Q}{c��V�����i�77J#-d�K�����ޖ[�9��u2P���a���<�̔�m]Jfȧ���v��*�k�56N:�&�]-���N�{�|�Ju���r���)�z�(O�@�ז��UʳRJ�E�����4)�y6�yVٹ�^=��ulsT-8ge���F<����|�Kn���Ԛ���wf[�'il��D>�Ҙ������Gj�z���#������=S�v<+����N�1�-	�iJ���;�9v��#��v7��X�S�H��f)wX!jW��73��Ζ{��E�(�f*+�r��3uZ�����Y�2HY�	T]��RL�p��k���A���[+��uyh�+n�z���k2��K+lT�R�j4���6-�gQ59X�W$��*՗�|���#�4^Sc_\�Z�,��c6�+�/Xfwov}�%XQ�U���w����SݻZU	Ϟ4-EC�A��\Dq$�[�H�.!�i�t�����W��Ƣ����X/���Y����WIg&������ޣ��![�m����3HI���L�ڼnd���;un��{���+�%MARma�*|L���_8�Aume�
�bQ���qG��:��|��]�o7��u�V�I�S����>nV�ދ#�y��6��"��%`�L���p�Mc�\�ٽ�o�,:�N�ܳ#��GYɂ̗k��+o�-̤6��|&H6kEo#������k�tA�N��1WR��Y�z����[ZޙZ9�^hT�u�a݋�X�V�:�{)��`�=aSa�$��fN�Ć�-P�*htІC�����4�:U&�9b�(-��rk�g2�p:(��&Ȍ�KU�ݝl�j�^���mqs4�ˍ(��`K�����W6z�%kwHqm웻Ҥ��편=�B�]�:�O�v�T��}���C��EN�'Z�1��������!����=��%�j�Wӊ�W&�˥OOH͊��V*����v�	U�t�˙��s��6��tdY!"��:t`1�/����&�.�ݠP�t�P���o*F$uNس�i��D%�.�ٶE�1ە})5�>K/]�M�٣h��i�� at&ޙ}����x��'H�V"ٮ��<�� ���Bh���)��5W�6^_J�y��<�(ye��35�ț�s�ǝ��)Zo�����Ʉ:�	Y�(���[54pfkU���V����5����M'slM2*}7�t��x�qDɽ�4��ż�r��ڪ΄�1L��{5��y̕ɭ��G�*�YV¹��3WlJ������M���M^���5���{�ĶbR��`�6k�o5lJ�AM�ɯ4K�jl��޴+%^0i�bڮSm�T)���i+Y�����M�NP ����%�t��2F�v��P1��Ϸm↖$v*�YݩIQ�s��nB*[sb`]X��,����C0q��bu�0Nׯ%�R%\�\�,YU�;�o������'lPvH�DP�0[Z6�W*i5�/.�Y��+�!���Be-�3�����n+Ĥ��E.�l3�.��Q��9�ʹ���vU�>:`�"W]KtD�[�.�ۺ'��Av$y�nVUnh/QOE�H/�`Q�8; �t&M�MְE^��C��m��E3+r(Ŝ���Zsw)-���j�S-�� ��wl��0Uڰ�Zه~ӕë��)j��·e�Mո8S�[;��c�e�|*V�|����٧��-�v͠�P�G^���!��B��3����eL�AU��=k?���׆5������
�(m�˶3av�e@0�,Ǻ���m�0e�u �p+,���8�be˙N){xb��Cc�� ��W,�w�w�,�����/{p�(U����0 G(�S����մ]�F��Lv�Ԋ�Mq�x�}�h��2�pK;t�0����G	*�|tt��au�
�7��&�0��y�cbjZu�,:���C
��t��1�m1{z������L'(�S[�T@U�ǽ�V�Qc����ˊ	�_��
����e���-F���������`�As=W�^o69p�anͭr�e-�9)�ǲLuލ\^��9��x��֒#dӶ�ty)��T��IP��Ů�ulj�������0XU�եb�-��'2FP�Ugr�^4n���9K#o��Y]���Eq��C�[0�V��}X��$ìC��b��Au�eҮIP]�4����A�X̆J7�tU.���M�	d�J<v`�u�no(��JSV��2�w|�<�kQ�s��ݶ��X�*�R��1{'N�#�
쭼�%��ǇE�jFb0�N]��;�3��n�ln۹�qs�:J��p$6��m�pvR���,�����Qq��'d��9������	2��%�����{D�VN�U*u!d\g�)h�38F�/�LlO��ͼ��P���Uo2!{t��jv� �ۨP�H����*�)f��9��]nYQυ�kҤ�HSA�՚Z�&���7b�t�*SGa˰�V�j \�a|v�x$e�܎�s91 �X�DF�̈́3\��~���Y��	�!�hc��҆�>4wta/pa�7E���y��p�*�0u۠���]U(��&��Y�ץ0��3�K���>��������_fB��O��M�]�N����_9Vt)�mQ�ʗ-��� )�t�����&��غ��Bf��S9�]Q�0u\s7 5�z�̏U��y�;�Je�Wj�B����[QYh�P����y��y���Z��u�!BM���5T�](�H���e�56�	� �%¯O҆v��f�|�p�š�R�1��Q��ỵM� %t�l+��{U�ooK.�I��,_a��/5¥i ���M�.�>�.�p���ѢP#��hɃJ��-H����h^Xij^N�F�a����v	í,��DY�05�yjd�oa��CF(I�j���4�O�;�2_&��pe�(�0c���K\[�T��7
��j8�uw��zf�j5	؞T7��M]]���v����ծ��R�V���x3y<��9C�E7�P����^Ǹ��tk����`U%p��c�@�A!Ó���<�@�c��U�Y{"4�b�ݒ�
�:�Śc��tN���\R���]W'ŬRdmhx���i��R)D��VM�3f�!���:���h0�i�4iJe�39�a<�+�`V\?�C뻗�����%�(�!��ye�"�K��1\�}��=�Ƥ�u6�₺��Cw��Z[��_��M.�,�Oc��ne�S��/���\�ݻ��rw���8;��Z=y����mH'c,���-J�d��,����UE0ETEUQEUDQSQIA2QQ%KQ4QT$�3DPD�T�5A�1T�DQQHD�DHTQ4UL��KTEDKQ%11D�4�4�QEUTd`IA5REAMUDPE0IUCE4YQSTP�L��UPf95EUUAMSDTLMIDCAf94R�fMSEVK�UDP�Y�fSf�FIEQEM�eR1T�E4�D��AT�TKM�E5TQL�SQ41RUADI0�4TE0�TEPDD����EM-U-U-S@TE4U-U%!UBPPPPQP�@UCEEA@��3U-5QR�QP��
���N�|A+�oe�I�[pF�oAg3/t����: d70Ǜk��9/�����
�0��s�jږ\*�������x�:��c�@����J�טr���ASz�wth:����޷���Eu�xs����D�]g��c�~�,����M���

7�Zs��#޼�m��h���C�=eo:ɱ�P��on��7�a��|mxJ��j��T��L>�)^1vZe�&m���W�'}[���q:7�;�W���F,5�!l(�r��8�o]5��R?8����뀮R���o���:�m���r㸇AWd��Z��j=0��R��	~����f��b���_�M<�9�Χu���!�=7bh�w�-s���\Y���,��|/�`weP��
�ܑKg��ה�)ۑU�J=��i��s���A8�����\�'M}'��*�����P��W:zg���(��	�E,iҍ�]q�źT����&�q�I֗ ����iq����"�������WF�̡B_�վ8��_�!���p�f�|�B�	%#����#=���ң[�N��D�����5Ռ�;Q��$֋���oo�_j��m�4*��n�Q=��o��l�u|g^�yӐ�W��n�!|[���$.��:"ɲ�>�(�a�z%JZ�w^u�R�b���1mԔ�&�!�c�H��x����w�k5�\rm����g��n��r���H�Rt��2X�)�Ժ�U}��B�3����7��J�>]�tTH�Ӝ�]p�-�����t7]��=w�&\�	S;q+of��Wj�K���"��,���]F�hy|j]P�I�C�D��c&����=ц��ӝ��73�z!�\M(҇��_�Q�y��zwR_��pu��׀��87ãI�奯#Ζ��
`g���K����{^
��L���Y:�G/��I)���4�Mgݽ1!ڔɒ��5��_LY)�@�ȗF�����d|�dÊ�̃'Z��X�XZk�ח#����~d���\	ۄ�l��p�q�:b�.U*B�1����Wq�g�+�KT��N��Ѱ�9{q�jt�{?�V(du�NJ�����n*wFҼmJD��`�rc��(�9qր����e�ڧ���e��s;8�
�eȋ9���FލL���~�Y�j�=�6U	� ��J�<�$a#��-�U�Ɏ��97)LN���\���V��,{/�����Q̃�.�����OV5Y蝬�}طi�'�:�Ԕ��X�uՙn�K�����Nj!6�u+��ͥ�{��[va]�p;o-��R;z�xgg�V��$ܕ�Y �G��s��sw9r���iy�/k��+m�M0�T��ێ������\5
�Adz���)�y�JQ[úTNZ7����}�n�c���ۆ��Μ���� Q�6�����H�i�`��蚜	�w#���**hI��s��)@��6ܦV;w���P�5�< �U�A�2�:#
TB�ǽ9��ME]K�c�}�Υ.qd�	���c����`3�	���C���ۺ�V��q�$/�3�g���'�R$aqߺ�]µ�(),X߽�
?y�!�����ĺ}F,9Oě;�۹85|#$�>�ᐄOǺ�M�y���}¡k�r�8#r��)���f	X��IJ!k;��O�'�U���erEMG1" CJ�iy�~\k�+�U�٭+&&m�{֧v����;Xn�uX"Q$���%t�0&xE��'ڴ����vVW��?9i�tS�cr�rn��Ys����P��#���>)T���C���h�Z_�Q�KGG	��7Oa��D;s¤�BIٓq�F�&*4�2OGO����O�܃)��Y�?�����O	I��t�7�kVp/����b��x��Ч&!K��k��{7vU��U�fX���0ؗɝ��8=�gt���  �T3�5��jaq����B򱹗&W,���2I�WwF�ǎ�<R�o
B�R��wF5p��H���1ϥY�^��ږ��?���Y����{͛w�į���d*���G���`��c�v�2�	\*/^$>�y.��}�W�2�X�2�t-t�F�t�l��F���qw.T����QWR#&�PL�ݨS�ђb�X��L�Ҧ.�=�t��<̖f��/�"���h�CWQ=oۜ-d�[.P��.r:�*�lTβx�
�^Un6N�ih���Sq3�\<U5̲v�k=i�����6"��
�rp�O\VO������z�5�ac1�vd���n<!d�����x��N�?b���PW l!�W^�mƗJ�U_�Vn��L�V7�
����=q���k"��
��LCe3������z�^q�[�Ӗf(X�*����G��{����+V��,��އ����q�B��L(3Y�ý?g=��`�(�:I�~B�:��=�s�˱(�Wz~��죎�1@��8�^���x�8��ҷ�F'U�`�*��7����L�:�|�t&�d^W��ɟ�������%��b�f�B��X9��N��5�H��1T��}���>Y��Vt(IIoy�����^�w�$�L��r�& �5;��=���!�E�>(�Ҩ�C�J�p\��-F���1]q���.��<V�(9���
��|���rg)�JȦe��vN@��n��wV�_�P"��4�I��_�y�'^��{;Q妇�.�p�T�𽖊������m���\����*A�u��jA��=��HH.5�x�;�1��T�*K��1�VY�F2S�d*Uy_#)#�3�9�%[��>����$;LMGm �+!�����|��KȀ��amH�[��f��j�F��TD�d��C��G�f	HW�u�}���STz�^���T�I*�M��g�nKJ���\g�?GK'����M���jC�dc�'2��������蟳&�[\���jt�p2���݋�/e`�
�M�	P��5o��~�G�-ҸW�O5ҎM��x�/:��jf��W2���W���h�iD�TA˙���7�;8vSNw����vO�J��Φ^���K�qT�;�ʬog+��G/��kJ�{�ٹ�Uۿ^T�O�_�0p
�\_SO>�����3���f�'!k̉��.��^�2�7'H��U�:����/���h\�+5�κ�p���{�z��:�N�R�ϑ�����v%+���Y�Y0$��>�899pM��YA�C4��F{��W^�:�->�W`�� ��LI���M�Vh�'ajĖrUA�>ږh"R�3��4B�,O�mP	`��\nH�S��D�d4}��̏�v]9�-���UTgr�vi'MD�f�ʯ�L>:!@(��U�"�o;���H�^�JG�rӇe�>� yq��3T�����#�p��GA'I@X}P��Q��# �z����le^�j���	��V��RY|r h�6���Ͳ�   :��Z`9��{��s���V9���6qۯ��8XKwԝ+^��B���B102�n�[+`��́�&H�%.�ϸ�Q]p�ڿ�����Cu�M��q<u�n�u�@r�]�k�j]���4�d@}Bt�<����cC�	r�4T$ա�]"b�UѼ��u�t&�5VBO�Mz��(x�����D��r������[�9{Kv(<^E�y�q�}�WB%��0V@t��L�{����b��P��إ�H��!�B9Џ�=�\5���=݇ye|�Q"�JdɸM���q�I��G�aB2�kI�[X�/;t{q��g��g�}�7 oQ� ��eƀ�U��>���t�')%�U,i_k�nKʛe�{V�Lɞ���/u�a!块׍11jN1����)��)؈V��hur�6�Wx�'��;�;qA>sH��>r�<u��;)��eLâ�""�ʲbX�[=����v��MB�˅����~d���N�YGc��8o�عd���x��tc�e9�ʖ��2�k��+�+ wh�b�>���q�g㶪��Y]�@���~Lɻ�({��c�$����7��h[����gAj^���74���B
���73y��H�ok�Q6�i�35�!�_*,ԵD��*�pT��!EFg�����g4�����&�{�5n;�j~��i��ep���)|��ی��U����\��W�"utmΕ��t>�蜮kd`�ɯ�O2��|ƨs�3m��+:rN���LI<�����0�ck5��Ja�_P�g�6�+�)�����x�=DS�u�V��_1�yb�% ��ب^p[�qyeWb�����}o��3�gk����*���u+�]�=�Փ.q�4#�x���A|H���\z�b^��g
�c��ь���<1�W�@y�hRd�FNqה�a�T],nFIF���8E�^&�'Q�ϸ��]��O�Π��)�;�x�΁U�.V�ݤ�Ո��	�U}C&��VN�iT����e��dM�H+�m�Oq�b��͋p��/��d
�uc�W����kcɕݮ��BW5r���:Er�	b��i0[�j�,y{�m����}�v����f[N�����S��C��`�4�IS� �p�����uX�x��ϣ|kE��yF�t��g����风gD6r�`6۸�y��$OQ��]@�0WZ� �9���q���w�摠�:���mB]nKf8C��-	�6>Sh�J�
?Sb������"rm����g���A���/M�:!۞&)$�ɶ�#<낧X<� �0�~�h̤����T6U��
'��D���*^��\5����6���#�w��D�.�����#bڐI��S*�]6�[(yf
�͗��;^S��TeWe���<��#9Oro�"_���9i{ƕ��4n��}a�x:�������n����\�ff�%.7�=���ټ ��KJ���CWQ=p����Lu�E�4���僖%�ek����&�RA]��.b'�+���k�d�Q�g������SC�lT��"螹v�T	��U�9#����5m���G*��bT�p3��))�0S��/3�f�};L5���A�䞷վe)S��)γ��-��Պ���cā�]G{�'�{0y}�xI%øT�Q�V���8+�$��k��2���zfw*�+���=7�²}�`�c��J�=,Yݺ��/�M.G��XRXOm�D�M ,���m)G����#u�.ຈt�$���TQ�CJ��
�Z1ܦy��|�Х����t�5�J5[s8\Y�#d�̃҅�L��,B�V��,�kw��0����c�_�q��I)�nsߡ�uܮP0��5�L��%�K�|j�_��{�ٚ��/b�rQy���9(��c��{���]���� Ȣ<�ʾ��ҫ��n��7�6��.�q@��z�1�r�#�-�#-�Z5q
d�FD��>˯bana��{�4���@�xE�|j�p�N�1��-��0E6�'-��4-L�o�M������p�"��Y"���_#����?*������i.�e�,�c%\3_C�H��3Z��9�U���%�3�U�&a;�Oa�492��A���'撦K*q,�T�Ǭ�U�9w�`n��",����X7�:���Y�|�z�N8B+��s_#a� ˥�v�^���;�� b�9`ip�����'�OP?D,��wڐ�#b��_v1����]·"�����[8���$�i�}[��P��y��]N5�_j���҇uc�Yn�,��7
������i�?5���+a��뎋��--	k��=��@ ����f���2]�c� }��ˍ;�ε���� �޼K�E-܀��6!_�������&�E�����]C�K.�xTτ���EoH�Ȣ�S���\�yJ�&Oޔ�����S0��N'Y�]ī���4�X6j��Qef�cᙻ^��F׾�������#���U<�J��>^uLq|w9U��U�%��EQp
t�n�g,�\}�@f2�+��n��t_0<,`@L_+�E�u4����ٗt��F��{���sa�}(���/���qe������'�m�,T��crFދ��b��cu���2i�7I��J�k�7��쿟Lhmխ$�"x�\�hנX+����!��r����rL�si:l7ON@�<���&b�*crV_��4k�X��������u'�3�sq���GVo5R���&��(MrV��RY|s�ڋ}p��6��F�P@���:d�큙{ES�\� ��`wt��2�T��p�--v��jN����}�R�5}�T�dx��Ojq��`ð �����E|O>��P�Z��m_��7���븑�����k�8 Ӂ^��e��ysl�V�q[�ug�4��2��\ U�An]�Ĝ��V�5�l��'.�<��`���L��%�f)<�D�V`�Wf̻Ho[y :r�
]B-���N��D���S����B$����b5Í���2��:����[����+:��`!���)sĎm��W����]]t:�J���٣��d�W]г,�-�!+�Q��p�"wk��[I+�VJ՜��Mkz�L�e�[R�P�B���3��Z�:�T�uʘ���rZ}K��,5R��\��P,��k3-P���U��$�b�X�ۂ��nw̾գ��8�S�����Ds�B��G�T�sյ����1Pڴ��l]�qaz�EX:���"p!+����Gls�rZ��Mh�}�/.p�>v�y�/��vk�r �V�Hjtr��+Z�2	d�]���9V�Q=��&[9��q�O&��� ����J��+U�䬒^u͎!�^�Q'$R��I͚�&���s5�T��\\��s�$d�uҘ�]>*���-[��D��oe���C�ùvO$(�'�f*�m�֥���c�r&V)�T�wtA򳉌zcW���Q0B53l���r����m������b�΀MV\m��8��.k|e��p%��y?�Y������okƓ�aj�\,�d�궲]���aPZM۝F���T��;����꽲�iO���R��	�É�(�!%�}qf��J�����G�����vY��jL��)�Pu��R�����+#њ���(V��r΍��,��80o9O@=�x��2P�u2C˻�}��egt���8�!���v�.����RumY�;3n�	�ci��!n��u��oY�.S�MkK��&��땵��٦�c�Q][(&/�;;��Q���ԋ[w$�C�5�3������}�o�S]R�p:�F�*<{�b�8����<��7 Y��s9nf]�ؾ�Xs�$b�����z���.��h�m%��P��0�6ƚ�FѩP.���kE@��D�Kݠ�3:��6N�����]��	�0�R��`��A:�`Y�mAwb�6���q��[���T��a�{]��I��:��u٪��t�5dmXr���$ߎIǊ�Z������"9*�[Tb0=F�r���@ﮢͰ�����kb������>�C4��cJ���N���\����퉫��E�z���p�i/l���e;P��}�If�n޼e��ϊ%5�>�G���s{b�)�]��+6$�{Һ�;�@�U��	4\�X��j�'E���N�d['h�1��*��ۏ�Җ�Oi�Pw�ܱ�gW�P�oy�WVӰ��H�o19����OS�Y��E���*'�[▐�[�3��˶�J����l��ʡ���)���b�o��2�]`#@��s8]]_u��x{�x)+��LI��Y��|�P��+�v'D֘�W{�J
(b*"�(��
B�b��b�������$������*"���(�)hbj����
� �I������)���(��������@����hB����
������Jj*)"��"(��$��")hhF���h(��)
�&*�h��iJ*��)�"Z(����h���������J� ����i��H��*%)��"�� ���
j�)������b �����&�hi((�B�i���*"h�Z���
"�Z")���$��)J

���ZF%"�F���Zbih���
bj!��b�*(�����h��*���JJZ��_|�U  U h�����gL�m���ŴCwn�*���5nJ�X�A19\	�2��e:��z#o"�F��+7pخ����F�#ky����	N��k�]i:��p�G�dPd}���Zr~����w��5	Z�~�߸=A�?=`��s�����.a�{9�{�%�##��K˩�D?[�Ք��/׏s�>�"8!���~�4�?���u��>�N��s1��Jw%�?Z���T�9��#�u�'\��7C�jz���=�Q�O��P�O����y.�GT��ig!�T����#��s����R����:�e�c�?��]C�9.{�w�h
��������d���w��v䤺,u.C��59ɪ��ˑ�n�ΰ���{����e�c��%�C�>�b"�H���Hn}����s�m��*��ﹰ���w�o�?A�չus�_�rd�_W�;�pd�Ǹ���jN�sp�3R������#	3_r������F���q�}>#�|D}C�e߸��U!k���������ך\�C�:y�{Gp��Oy�����BWﵥ����5?~���Zrwy��w�����5?~���A����=�q/uo��E^����DC A|Y�8DL%���n�����>����\��^�9W��5P~�P������f��2~�;}������	O�9�׬�婡��4�
y��.������_��&:������K�}}��1��X����j����5&��<�փp�O�m���O�j���ᯣ�uFkA����5��;?{��yNK�>~���(~�#�����^`�:�ﳯu��V#�3��y�r���}�
@y�7=K��Ƽ����
}��Q�u���}�S��A��ѸJy��Ӭ>�A�%S��������A�`��W��sz�9&I�h�V�~4=Gw�����+��c�2��lz�b��W﷦��g����y.�<�#�q;�ϒ�����ػ�T����ը}�;���7<����Xn|��)�wF���5!�۹*��z��7��}
+� �� ��5|k�!��i���5��/��j^�y�s�غ����%Q����oA�	~������y.K�~�cq�]ڟ%���>A�R�5Q�X���2�U����^�0g��(�z�T7o4Ե<Y�?�f�s����^x��g\��3,X�..Z���{��}|$�=�,��
1��@�m�w6��
��tz�J�҆��o��r�����*6�ʏ�{Y�є�l�kL<n�	�2A��R4h���5|�Ds��d���׾{���q���<��7�^^��+�a�w�;�4���.�(}?sA�乬C�oT�rMG!�����>�Q�}���J����.��Ht�(�"��>�>���2O�����w�y���=I���8k�-����l�������hr^��X�u�sk���i29��=�����I�!��1�/o����\�ZP�מu��}��=A�J>���A�l�^`�F�`��;��d�&�֏oe�:�#�X}�K�jN�{�pu	o>����g��\��3��kk������<�����}">��zxuM,��w7�^{�9y�σ�:�-C��X\�2uv��y��~��)����ܚ��P�PPy��Y�K���m�r�=^K�������.�����i��o�6�������"s}<����|��>�z뿗�<�$����:�K���O��p�^K���lMÐe�:>ޓ��`�;�������n��NK���S[3�(0>Ü��|�5���1>��h{ e��wI]��s�S�u&��9��7	A�9�ǫ�rK��zw�C_G���������5�g�k�{��2r>�&��2��a�ܺ��.�éw����a�)����;��;L�]��]��@��t|!��?��������ZCs�N��<�a��J|����os��Hw���>���Gz�@o��j5}�M�w&G�1�wr]C�3�惸wj~�>��hU��Y/���|9oB�}�"����>�|�����p�/ӓ�r��' �qN���4����{}�aְL����~�$�w�������M[�Pw���QA�}w�i���vh����zT�m%��`b>�C�Q��'�b��J�BS���\��B]o�=����������_֧���JA��{֎�(y\=��^���7>��1yn7��ן��߿n��\����\�ڏ<�BP��u��ܹ���;��Rj<��3�n�c�;��� �%;��w~�����t��C_G�~���};|%�_K��u�����{�6Iv�1�_��X�X�M�Ջs\�������~� ���%�	�n���>9)�>�V������B*^�)�4�a�utY����;�^�z���͘�ʸONCn�vr��9��&`�S����\1�u�b��=���T[�=���뙒?�6FK���߷�����;��v���rSԹ���7&�ʓ����j5�:��x&O �uA�n�^�c�z���j~�?LD|= d {������<{s�����>��`	��<���� 8�o{MG��u�����>�+�^F����P����N��\��a�l�S�ܝy����/��u�!�y=�".$ǄEi������o��C��Fm���<���u�>yjNO#Ru�n|��Ԛ���4�Z(7��l��_b�y���>�C��u�Д��.�þ}���U����x>��L����O�s��@}�K���ֺ��x{�����s�<ߝ{�/p�^I�a��HP�=�ܗ���.�]h�^�����y���\�]�m�*����>sS�sXzs����Q���Z}�BS����?`�DH��`co��L������k]����s~���R{��Ź���#���&�9=�Fk%�<�-ƥ�ْ��ZyQ���0�sԹC��}�䤧%ˣ�i2>���L������}���xw���o}�Kʪ���pwo�D|}�@`ML@ѨJ:�{��w?A�;�U&A��l�4%���a��w���7&���u'nu���C��^u�C�	s=�>��ϒ��뙽s�=ޭP������ٽ-F��":�h����è3����gU!C��j׸���0L�jN�I��5/��S욍I����*��:�>�`�%�N��S���u{/���������.���|ߝ�|<[K:.�C�>����@ G��u����59��a����'a���K�����=��w^O>��:�
�,]˨�1�f�%����7o ��\��a�sBU���z�5�W�Ǽ�^�}�q5^����H���z1^\}<�I������;����}��{�jӛѺ����<�_��lM�C^�]��׸FO����w�%�=Go0��\�d�o�JFK�p7ֺ��g��X�����YK{X���>����HQ�Ԕ��=����jNI�w�����5\�ݏ^��>���}��>���$f=���~�A�����O�d�?}���������;��PFu,�X��r�"p6��3V�8�]G⻆SQ��ZƆL��c2"����<*����t@�֗6��-=L��΃ʭ���,�H��T�6��� ��|&�]�p��I�|����ַ�qʕ�j����;���ʝ}-	oyි�B_9��{����Ur�wk�5���y����Oѫr�~����+��fF���xk����rܼ��9=��C�~�9�����*B����}���#�g���MOИ�0f~>�|	��6���F=^|�����o��%R�}�����-���S��uyy��p���'y�����+�z���������a캩���惨FG����o�Թ�dzU}���� Dgyܦ���=hZ�����?{�^��9W%�k�[�:�e�����:ֲ����o0>���=�!�5>A��u�'��MvkG����)�0�Mǐ~�Rxu������Һu0Ժ��¨]}v\f����Y#����~����~k�z��?s�mz���=�����>̀����?A���k��g4��r?FA�թ))�?{���5��:��HP�<�GZ��;���ϯ��nf��~�𿊏~kuw��n�a�>ncE^�GZN�NF�@962���ݎ&lC��ܱΣ����:�����_q�[�����{��~>&�I����ޝՓ��Cj�����'���O��{�X���)�S���a��#�}'�'/:���YdK�qG7�Uc_�=��2�J�⏽�ON�{ٌy2��>(dU�a�4`@M�]G��|5�w!6���7���:��z��	;��[�w'|3�B���
�FvP��
sq�J�'�N�Ǟ�<;6HiO'<�X�_:�nJ���eH۹�N�H�Es��5�FWx�"O,k۫�,��zv�W��^R1��i*y=i�|�x��l ���axM�K�N��Nv�ZՄZ�z[�r�m���5I���.�n^ķ�+i�0��}]g	α�v
����� �w(�T]!! �gM�k{���sjw:u�1���QU%J�ʱ�����f��o��!���;��9R�tD���ba �~Ѱ0�0r;��fyc��ѩ�Y�ĩ��q�Bk�J�jK/�@�m��@3L� �(�^r��u9ܽ���Q�`pN�!J��?_]Rg"��i�0%�����,}�
r���j�	�II٫ޓ����� le��H�'�NdGB)k�2%�\3zX�"0�EW���E�ZȀ�o���g�UƇ���ZM/���3Z=�*�t�D��W�8�}9]����g��p8�.�?1a����wF1<~H����o�uh�-}�w峢K��o������AϤ=LTm�*�M6�x0�5`*�o���U@w�1},x�:ͷl�W3S�� ӽ�n���1����Ǒ2_ɺ�9�{1d�0�N����U�C"�jY<�8,bG`�Q�����/�v�����
�����U�}Vq��1N�~8��y���c�h�Z���U��װ�t�=&��5p���a���>��N�07�`w�٦��ʅ���7���⏓��S e�!����<�H�:	�e�Uu���	(��r�����{��Y�FY�>�敛�xҵ/;1���
'K�r�]%�+1�n�X�K.mK݉V�*Q
+�,�gvYHR&�u!*#��lj��E;s���b�rz���������G!���g�,*v�y��K�wmc�b��(��\����>Б�\r��jW���=��Q4m���3��@���|�,�TI��x�oz��a&�{�=��1`�g>�9��E���i���5����a�� �%P8�}[|��qA�4JK�]Nn�Ք�˘�͝�X,2k��/�-��s<"��Μ���d��4)ι�c�za�ި�G�s(+���:��0���jx�+�)�����tx\6t���5��ty�4e��x(��|W��¸���Wb������|!�`3���*;r�͹��f�ꅸf1?��c?\@���:I�(	���_0��]�K�V��%�1�\���Ӿ4v�+��9�
���pN�B�%��7��()�s�y���5�s_]ݯ?RT
�e�ȧn��~��u��)���:C���0S�J$��� F'�!�ZL�*�Hc�f��'�yM�4���Y�~i:H���rlm�y���xdh�YlOx�R���R��뭥��9-%N>�k��]f���A�6�3U��x�ǎ�v{ڑ.�K�=P�m�zD'Ơ@ g{:����+*�[����J�s9����5�O)؈hJ}���tS�Wa ���k��,���5���ט�i�ntٝN�������
�	�KӍ]��ú߰4�a�A�mB]nKf80���K�F�
�6���Op��kۙ�F/{=��Bju�<��\t<&sWi���#�Фca$�ɸ��#ZU�&���T���˛+�q�~r��~�V9�T{UKfg��*YI�}/�s��~zB5��ky%���;�>+�Խ[��E�UK}m����1�t���0�t��z��bػ�ݼ5��I����W������p�Rk]j��PS�71C��D^NW��^ژs�c�T�G�����Fz@�)�o6ձ�d�T�4q���wZ7�s^���%Y̨�a�3���0�QHmd6qf1���x
̪ϩ�N��*�L�v"�k=&��jo�|"��-�j"RsH���;X�}Y���y�-�tp_Ɲ�4��Q�:�!]r=�X��@��>���yz�L��Nsb�P���Gp,W:P��b*#iPEg�51�φ����?
�6�2��M/h��b)8rVg5�*��iq�4��31z�����
��+�V��*���Ld=h9ΘGZڹw��4}����iS��M���X�q��
��-�w&�k��,xR��k�=u�	��b�d%+b|x���o+�������Y�uåpv�m���F!iRs7)#�V\�w3�)kYO�̾��Z��=J��}�edl�e�|�λ����o����epY$�_#ĕPg�!�$�x$��hw7<u�8�~�]a1+g�*�jK1�h���{�#S������ ���1W[[�~��&XR�4����r���|������f�9	��ݑ��ѫ�2��0Ù�AmD�N$�r�]i�@�]|* ���q�[�Ô�l�6Z,�����P�sH'\t��8�S��� 1�j"��T�蘺�ʼ2�ҹA������j�'�,��:{��O�l-'�5🶺��'���Y2������A�˕��#[8�t��9��1JK��r�r?=n�*`kQDE�)�D����c��+(��
!FN!�{�]�l���i����[Q���a�5EF b�9`ip��ߋ��OW������G�����V�S��/o.��.:�GyLh������ޝN@rb��S�}�e��
��;}��U�JQ{z M�Zϖ�v�=�|�`�������e<1i8�ekWq*�6�4�=�.���!6���l����^�"��Y��rD�^�W�����Yˌ�F!�N�r���W�����C���\�Y�ǋ�ݏd�"t�T&5�j���	�F4��&m��:dI?k�դ����������ܢ���[M�t�/�Z�Mi1���i��;}?���}U[퓃k�w��`���ET+/M\2��F!�D�����@^�pt�"ʛGVӇ�Q�r2)�jg�xRp��1qyS��ᢽT�<6_0<.�}s�53��l�u�&��A�6��!%�*��ف��m���t6<s�f�L*,O� %ґ�V7�pp�e�k%s�dX�%$<S��;�#T:�nD�*��6p�^�@y|��S=[��8���X�Qvc 5��w8�zr h�_��1p�S�+/��p��tw(�v��%Z��+��t��yP�*e��ـ�'���q(�/�ڋ}p��\�/ZB���;}s�v��79��n ��x�RS�T�g�v�鯜���Z�#�ԝ*c�g��ڣJ��t�}���L��@�]��'���!k�:[WUJ�4�������[2���*�&�Z�'�L�����|�IO8��5����q�殮�Es�L��n�e�&c&��Z�����D�����b~��*5:�	���MI��,�-�r�hs�ļ.������p�'|��2�``V��1w<��OeKZ��9�֚w��ӽ�G�V�����e`��ڳ��.&YҦ��Ь�,i�h��P�0���!�i��=]Q�J9W1�{�ȱ���J�3�b������}�}R�,n��-5ƫН��B�*6�T2i�\���
`es|���*�;ĕ-ŴV}�y��䫗^��U�����7�t�6����2:-JdɸM���}1d��Ne����z*��d��Xuz�,ꇅ�_T��q�cB�˯.}����?2]{�-ˣ�S�DW�����U��2Ng���GTv�Fo(�߅x�{Z�i1�Ph�_:}�����Tnm�/eQ�V�|+�Mg�ms�}}O��T���_�~R�:��Ơ��9c6�"5R�KBAoi';�ݗ�PB��xҿ}#���S�0ё�{^��52+�'3L�¨{�ʨ�-0 x/gz�D��6�fx�Hm�)�� �j�؞u�����p��u�zw���[��; N��k�g$���ݴ��3�V���\P��S̾�w�nxFm�\!YӒt-�D��<A�)j�r�-�$���`'�즔�����_GC9�7\�q�7�����{�]X�s�}�z��y��%�%�G����(p�T�p]=���>��&��c�|!�>��iN2�T��P1d�N�]���u-9/f,�|���dR�ԯ-�fE�Cc(���
��r�<��E%�qS�V��&����LWV��DSz��Ѽ�؅Z&Z1�6��ˉ��C�y�| 4���҄�6r��-�y��
��T۽Ь�jR3Em����n֊��u��]z2и��ر;�V�u�-�	ԏfv��Ƶ�U����nQ���n��mɏ���p��F��&�ܡn�A�2���#�ƋiGݲiH��M���F`�ص��zP��J�)��q�B��r�i�Q�0�j7�n��v��q�i�:��E��I��G{n���sVvR��((U��Iج[:�Gnfn�WR+ZȾs��scVpe��gH�tE�����՝��s�h@���\�`��D�[�pr`3n�[7��m�HL5]�/s��7$��ȃ~՜�����G��1�i��v��]k�c�kYN���E��(ƙ���V)eZ
S��H��֞Ŋ��gk8N�x�-�j$9�\�
�rSܴ��.��D=�ӻ}&v�F����O;��c+�1ήf��v�P0�f���ss�|vƓM�1T�Y�@�����[�'a��Fk�D,Ʒ^�u{ԩS��h0h��IZ�gr+ecX�u�`��-�"�0�J�}>�ھ3�ne�+�ղ��ș܅�	�` 0��Vt��Ĉ�Q�|n`?��Ba-,�j��$���N�Z��.��MUê��鄈61@I�n�*����֞ ��n6iC�]w|P�Ӵ�.9��i'+���Y��N�����W"�aQYK	;��:Ks�9�O'eh�Z��s�c[��5�ʁ�)�U9{��!O^�ӰH�"��&iG7I��4]��<����WqWP�9�f^_ǫ��S�񁖒 �nNn�v`�1�A� j� �`�^��Ô{��ض�s%,t�T<�����w���{:Zgt���Vk�8�t��fm]b;j��-�(��t�Y���Џ��P���b�+M�FY�"܄S���mWr�뾀+�[tnsfs@���xoN�P��|"\�������sa�E�<����9���c�
t̓+O3��=\��H+N�\��J݀��s���4��4�;�D:����l�å:+E�c:gAr�3�17i-@rI[�/��j���
�^Чu+t�!%L9c��h�.��V�&� �z���	�d)��0�0pvź�����Rh�V�Le�g@�>�?y�wͪ�=�7��Y]�/�9f���;�x���Uv�]���L���R@5W�.��"K�`-�a��v	/!�f���A�h\�+���kT��[�>�������o{u1X��YL�����;�bQ�!�����<n�����9��dv��X ӕ���Ջ��֮�����iga�+T%�l�)��vZ�FF:ʡ�٫�7�ν`�*$�!(hZZh����hJ����
Z�V&�(�j���	����&�)ZR��%ii

h���R���"J��)J��b
JR��hh"
(H�"

D��i
h�(
��d(��������X��"V��X�����������(�hJ
)h�)�
��i��J (h���h��B�)
��J��)R��
�����hZ ��*��)Z ������)��()i�Jh�H�"�h
j�b�s�x�ckoX�#�|%+7zԦ�]�ִ*`��#oH�
��
�4��6��� ���9�QU��4Wn���}DD[�ç������W*���y��,W\t�\BC��]�K��w
�p�\�#Yp1L4���:�-&θs�;w,�t}�PR�&��e`�ڜ�N�	�y����ފ�/~���o�*�;�ܾ9��M�yP����� q�B����xo��-vF=ĝ�}bxBo>����I�G>s:!��v��hf�OO��o�m6;*/4n�6�l�K& #8�%����S7��6��rm����\�%��� o�l����x��l��O��Cw0Q�x:�WҦ�A���+������E*��0D<,�N��^m�	M�H��{B�K�;h���~�c�R=�����'P�^/�[�����Ѻ(�S��C��d�!̶Xy��T�ۖ�	}Vr��H}���F1.��Z�֜v����܁�pc�勄������5p�()�lč����EFNP66wj��\�Fo����ܥi&��7����;�T�4r���� ��!��5߀��aVҦ���$Cr0&ۙ�j��ľ~���~*�g<�}��o��'Z�J����C|��`�z)�K�h	k���^������5	Zѽ�`���+ށ����\�����N�6�c'��ƣY�宸�6����RK�h׀҄�U��}}�}��F�Ʃ��>���v�X'�	�T~��u��"���g�Vxk�s�}����6�Hmf��6��b5'\�_	��L�8����U����A,��|�,X��uW��K���f/�8��wQ�.�҅�ng��lۂY��j׻����$��p�v�Z#x�:�t.���5������ ���iHo����|��W�Kf�ojnu���l4�FC�0�=�t7=7++���Q��$�����]�l:��si��S�e8Ӄ�����ن��w��{g�R��r��k�!�臽R6ӻ���V) oOC�ͺ�t�j�V��N��W2�.�i=����\U��{�&�=�ru}m�p��##Th���*qr�`�q
G���_
�S<"�p\j!oWȅN�1��-LX��M�S�;�C��]^&�k�S޻�X��$x�h��������1z���R�a�Kb�d����a=�j'�d���>uA�VM�Y��L;uA*���#G��zNk�쯨���ܺ���I٠��{z�E���������oyE�cY1A��%�
cm�~ȗ{�b�>�C�ެ�����	;�wv�`7[Z��&s2a��l��-x�vh,yG�'o��؁��q2.���Qe%i�kI�sS��O��̙8]��m5���1SUz�Ι�>����#�B�M��ŻS�h�����IS%�,j(��%:����+!��J�7�m�0W����^�ᬼ�6��N�ګ�xX���f�\Ax~,���Gх�������&��vz�*�{6:aՖ+d���N`r7��ˣ�I�z�9��d�iհףD���A�1xz�/�ո2�}	�a����L���'�_�U��YXjvZYf�-T���QQ��Ə0��u�î-ã��ON\gR�Z�c%Ӹ���T�\D�y�z߬�!z��z�?S����q�w�ua	��W5��*��� ��}�UBPi3�U��=8���o>�l�C��t�7����ڞ7e������������lN���}�d��@W8����9#�O7=�򘎷U��ȃ���b7�� `Do�J@i^��:ܣ�T��*A�]:��Nꆘ��z!�����LiW\&9Ql\�]t��=��tS�,W����m.?5��.�N{���Cp��t�Y�hMv�����ث1���@��r5�/":��A9�t���@(Ǝ�6��F1R�n�&Uӭ̤��|\X{�k�k,�t�]���mN���[�,�̕6�]�B뫤{rlƏ41�ō�e\t�;�7���}ߧ�������8����^Q����(�'�B(����x���,p�p��H�����L�q9���!:{�����u2x�J ltPU�5�Hd�E��Ю����t�w륮@܋խU�w|�F�cS��z���t����T"�G�ZM%<�7T�h�0V��s2���s��t��]o��)&��.�1a����Z�Q"1��b� ���m���M�?�[ǦE���_pp�
��U�m��� �p�X��<iL�b,]Ƽ�c-ڕ�A����o{�����bO������L�6��9�2,�M��lb�^Js��m�a�b�PS�p��T����a��|B���Ǫ=��^ϼ=�A�5^��wQW}�T����'��\;�=�a�����Z��`�F��s��W�(;;F��N�ƹm�Ǆ�����7�W���|)���-�����3P���9��L=4
8=}Vk�ѳ���u�����e�ڧ�c��}���(�O���3]�{�÷���\`Һ�ؽb4z���G.Lҽ��-̈t�{jY��]�Z�V��tR���h� �� k8k�4����.���	�y��1�R�K�4"�!O�Tk�<�#}'`�#���m�����]I���ܨ���Gi�}�x��?iY����u��u��#��}UU�|0덟s%yIHw��@���.�.y�6N|X�}7ܶ��^��E�l�@^��m;�.a+棱�Z\ڇt�����h��X,2ye�����\9��T!=���냙��o�����F_�z@@������UK��]���ρ�T8�nS(�⣷T���
��
���4W(�稃���\%Om�r��T�u�����X�j�C�O�#ـ��Cj��Z�EC"�OW�e �(�����X���vm��M���:��,`���h�D>������v���}��a@�)V��5��{Ns���E�m����s�5����[�q���9:C��s eC�J$�� c]"y�Y"-Q��`�WӭtC�������?>5���$�#�9��g&����f�H��gF �l��@��O�&FI)K& !��*$�83>�)��ƥ���s!���-M"���ͼz�9���Jzn�Y�~�����k�\x�^::��M��G���h�noz#=lˢ���R��k4�
4��Y��ִ�ц.��[���ⲅugS~��!{N
�g��a��t�[��;��[�2���h�R�.ҼH��A-( �&�>�α����Z�uk�I�J�S`�zؽ�b&(-�T�"`8��Y]Q�[�9���}��_UW�P��������ʥ:��5���"\<Lc���h�Uc>\���*�R>��-����!�{�S�=��|���p!L�r��P��k��o%��2a���!��{	w�4�������L�ޤi�p����U�ꘋ���5mS�{Ɛ��O�<N:�x��z��VL^u6#��:��J��J�����8�Tfڶ d�5LCE�������n�����ˑn��%���W4���/���Q,�;�8J�j�l�:�����&Dc;ɫ���1U=�.���'��۾�� ]���M�Ϧz2�g�G"����D4��5�*ط�b����S�u�,�!1	yޖ+ԁ���1�e�t��T�[J�+ l�j�B�crh��+*�_0�~xt��L�G���ϊ���Lk��Vh
�~�T|-�l]Nєc��֚�����0m�{���쁭ތ��a��{D=�����]pYpA� M�%wzk��q���2��>�
A�q]TJ/�Kg�*����qh���L����p(�7"��]�O6m����z�]CWceD����K��6ó#4ܢr�l���e���O��	��R]I��o0�$�M�U�;Pˊ��%-�˦u�%�t|��9�j�&�����u�bEZ2X��@(0���m�}���)8�M����vk3�����Sk�_}U�}U�p��yz_� d_���������:|e��p�a�Ӑ��Vݑ� W1�k(���$�h�$Az�d!*�P)�p8.+zxoB�m��6Z;3Z��a�EU���^ueש�*8���[�GD��CQOD�>U���[�-��F�n�#J�7��*]Hpj[��1����|:zD�����Y'�ɐ��؋�A$������N5;!�:O�	*d�e��Q`L'QÀ���}�����:������'OC��]c&�.��t�}5E�`)9`ix���/�c����{P��n���Y���8=@�Y�Z��Ս�@�̥{{6#�'w�#S��E��on�][b0�3��X[x�y��W�e�٠�޻��_M�=+�ӚS.3��ȘvcRq\ʚgp9�&i%�蜚x���dO8T3���4o�2��S�d�u�S�~1��rj�O=ҽ|@X�!5{D���WJPʫc`)��I�b�K��PU�6)�C�ٜ8iPl	SU'_^�Bɍ��rV�Y�dC�ىM�/T4o�k�2�%�;e�|)�/^�c��vu��4;T�0���Bہ��`�G�p[��eR�AW]�voT��,�wvP9�Ⓜ�T�8��]��,.̏���o�N����UW�T+i��<�`{��:Zw�P�=����m�L�0�x	8g�x��G�{�r�0�s�V���^��%j�烪�nH��O7=�)��u\Ү���R6��t���P�L��Qy��u�u���I�Ƣ��Y���qt�����pًt��ȕ��D�7�L��64�s�Mz	8�/ �u�����B�`bk�j������ƍ�(5|��N�l
�o�qQ���G�X(�( p�%1���jiO��T��n��r�7��|�\+,nڜ�|���Z\s��\d��9�B��(���2�I s��;Il�<�r]��N޹�3Ã���������u�K�Q:xU9�ʭWڬ�N�j�������i�޽[�5o)�BS����\�&�]"~b�'[u�_���M,���%�����e'k��oNv��R�q�fC�G��.B�n9T2ju����4!B�@ҩ�̑<ݞ���d�@ŗ?I�u)��}Ҹ�Oo��Ď�)�&��`O�}��PK�'Vݫ��k3k/D��;W�A�G��u;�b�A_���v��0�uȏث1�Z��bF:@���tX�K��ml�C�mw�<^�h��x��BO)Bw��(��N
	�]���+�[���H��r۰\᧳j��ǥ�F6��Ϫ�����}�N#����7��Lg�aB01a��=��Ŷ�ڸD[�M?n�U�K�5K�)7�^?�g%^.��c�a�]���*;�1�W�\�I��6Pc�׮]��Y�{�[Q?.��/�&�h��+����'j渌�c�WO��`�,F)��qu��\��� ۊ��FY�n��a�#4���FUԋ���b�	�=gΠ�+���q�W����q;1¦e�=�a�&;�.'�Cd�+�����u��u�Qx�Q���v�����`������ʵ�%�ֳѳ��+�Mr�e��n�c��̈́x�P,F�]�R���_>{ˣ�nrO��I�8z�u��G�#]��9�=S*��C
��~��V�E��|y����p����/�#�
5[$�(	�X��}�oϖWb�����G��X˅����u1���6�aU��t,WI���2�+,U�r��1s�1�gS���"q·�(_ʥ�m4cI���85	۸y��,��7�
���F �E�oI�˹���l�y���s�՛�N儃sX��*2���r��+�rk�pY���JՎeZ%�v.��9�\��;�_���9Rr��$�P�(�Nŧ�F�֭�4Շ�&9ȫ���ND=X�\�:-�|�ΤiV�zp��b����}U��D�U�#y��7xO��g���T-}qN]G�K���I��1ד�*[�v7"��kew 	�"ڦ�+Ḱ?.4��}I:H������m��;*� �ṹsKX�j�r޵{|"[�'�C�/�ɀ���+�+Nϴ�f��1��]nM�s!��d�X�>�.疓�&�p��!Q��>31��V�1# 0ȭ�� ߰_��,m�O��<��$�*LbJ����kBb�K�$�D�Y��4�tu��/a~X�����-�8	n��3��9�dCк��/����S)���B�U �d~U�lkr��+��Y��Z���(C�޴4Xʹb��1��e|�()ٸnb�u]H����uh���=�K9�`��ͧ�VSF�f0FΔ��m�c	���!�{�������܇��Hġ/'�qN���v��a2���X'|�65pԙL�\Q�g��Ȯp`��n�Y%�J�5���9���oi��2YЗ�����Q|Ǣë�롮��W�����xk���1�H	R������;eN��ԆvSX�$��$G�����(-'ٗ��� ��sQ����V��'+|�)h�3YdY�q�ċ\k@ Ծ�T��D�-��]�M�9	w�|�3[��U�9-/E�ђ�d�02^��f���9�[d_"Q5'|�̉p���4�p{|��XK����9M�%K%fAF�Z O-�:�.ڠ%����=OT-fLN��řmݭ�'��7|O1�ܓ�RmCm�w�v��Ӥ0�@&�gk�tWBù �ʂΎi��r\��D��D)ecS�`�}���cJ�o&W2��X�����e_8�'�r@�5���	�\n�i����x�h����PWr���촰��(�,��л��J�m*����Z�A�iӝ�B���Upa�6"�S�w�]j,in�*���ۭ����.�r5�9{�k�#�D%n�OjK1�K�i_
 o>yJm�yѸ�ι<:�N*��"�W�)v+^�c�K��řPo �څ�	�w���fƕr�3;"�>���S�n]A�*>�O�ϊ��g}pea�8��kH;(hb^�]�2ohP��i�F�����Qw�|UhES�T͵uu�J��[��en��dZGVC��1��6i���ק�*Ɇ��/F�[*�BfN��$	��x?���Jƀ�X��٣w[�4�E��|�*��d�Ջ��1`��w��KR��A�cZ�V�6�^� 25U��)ŗ��4��G�5h�0���̹�Dy�T`�'�3CK�G�e3C#��d�ʙ]&)�_KЖ�oV��
@���͙]������ζY��N�{i��Eu\��FR�Ɔ�ub�X�mӤ	�Z�Y��P+E\Y��R�8��k�m���?-ˮM!��{UŌ�n�e�7�r\6�M#���2��!5�^��
��Ur�ek�v�#�N�CV:����:��<;�h �v_+�uCJ�e����@��4�c�4���e�}��[�(ܖ.����E��3��-�V��i�; 6*\���n�5�zWܥ����z�ugRT��l���r�@��r�ٯCy���x	��*^+�����rX9�o(��D�RN�j�<��Y�[EP�4��:'d�d���g)�-��+B����2�bte#��\4Kޮ�F#����Z�o���&@B�P��hTk~��n�N��ĆzeD{;M��q���
��#Z5P�J{�v��tȧÕ��{
���������Q�_T�9�"P8������~Aux<�:�/1J�P���9�<��/�c#��4�{����'�ן$lv��@+�X@r���_�e�jk��p�](��Xu-��tQ�;
c���mՒ*�oJx���y�)�h�S�����ﵫ�i�.���|�#�艙h��� �M�v��[�v�]��QN�C2����*�qah:�P�@PDPPP��M STH4Д�	IAR�@P	T�4�R��4� P�- RīB4P4�P���@�4��)J �-#A@+JҴ,M4P�E!CJ%QDUE($J�%)K@�
P,TH� �KIKH#@4R�" �%RQB�4#H�ʔ�-R �P��MQwU]nwe�5�mn-]m�,��e:�R���^���Rk�,�\U�4QѩӉ'&��uK)���4Q�Φ�\n���g����""-,�f��e!5��t��%�=�
�@�Cj��Mؗ�a	yH�]a�|9��m`����<�M9u3{C-���+��m�g��pk>3�\�;f �&n �R�_\�j6�U���Z-���h�/�TpG[�v!`��F>e���w��q*��%�4�-oxżI�8%�Ǽ��(V��'��컉f�-��!J��!�,���!��Ćw���^�2ư��j/3�5�� ��$9����OS�A�{��U�4缈�Z��̯d�
��!���������HJQa uw/��
g�\�Bޮ���c-R�ݹ��՝�x����]+N�!���N�C��X��H�u\�+I��L.5�p-Ol\���+Z�H�_�ݰ�-Qe�1��!��%R��I��L�;�=����iTux]sv�s|}�;�+u�Z�d1l��%L�����Gy�*���T
������t��)U��%{��[��"8\��1����mUѼ, �Br���������N�4�*䄠=�.�]4bW
�Ou1��^�x�����;���#%k�x�Q��_��m�����=pvrw���e)A}%v�y��ƭwuB���xWq�)Cm�#]lzOn�m����J�m���4S������OE�ݭ�NJӼ�N������g�ԛ����R>96��3��|W)���rN��{�#t1�
ڃɿY�V��mS}2���yz#�3��厸?*��<�����/��@+�( {���Wׄ�z�PIZ빅�;�'-���]c���TB��j���ȍ���~�J~���!��J�Y6uW|&t��i�s��.;�uAWd��*_�bY��<LT���p�P�n�p��b8 �_SO>e��!�}�m������,������mt@�؜i�˧��#'M}��Y��p1�"��s�򘎷U��*��]�#xs`�{Ip���5G��}	Λ�d�}H�Y^R��|�]��.��!�����S�j�v��R�}$����{eɯT:	:O������Z�B�O��~�=�x{@H�f[�|LnԣY}Y6_B�8E��;�.
�e���J$����`4���L�_L�ks������ś�Qx��9o[GZ��_ؼ>������x��D��ʁ��C&z,hb����f�,R�^��
���k�ͺ�]��v.�/
+�Ȁ�����AU���Ű͙��뀐�J����m��Ω�n���m���卅ghr�"���f�Fte�ZD�i��7���q�����V��6�8�H:s��e������Zt|�#l��suÆJj��oK��q7]��ߗξ�C��E�-&���Fv+(��97�W=];}E�crᚆ�u�)&��.�1q�c%�8�:ǑW1Wӹ:��0�IY�B�ѕ�tߌ#	[�C�������ĺM��� `B(
��-���c5g��u��Y�ޙc�\'�b������2ԪE3�n;�q��{_ͪ�jS&L��}J~��S7��#w��Z���P kM3�G%��Ň'���8�ؼ:��u��(;cy��I'����r����"�@PY(D���~�zV�`i".Gh#"*�
0-���Ͻ�z&h�ˣa���}���b���mU�׈��h��Չwy�\�p�d�[ݧ��J,,��| ��U\|����5O��CSCx�k��&�E\t�wi󺺜�����.2���&,��՝�os1�=�	� �Ĭ��u��X�})���Z;b�����Z:	閤彈י���2�ѝ�w�:�n:�!�4��a���?5]����U*ޫ��u���:����޺��0�*b[�/2:�kS�NQ�0�0D�����k���;2R���{�� ̕jt΂�˵c��5�LW7Դ&OD�����9!{3�
��1��&s�!μV.Q%����vB�[XNV�xoE�[.�8����}�D�ӵJ�p��Eg���Μ����D�TLD��iz*��F�����ۉW+�u�����ݨ�q��+��B�Q�$QP����my��^	��{���֌���u%�[V�����ϡ�v��p� ��?X�\8i&g�W �	��->G3'�,/�6���GSmQ�M�n��9�}t$f�*�l�|�D!�f�&1cU�����wR��dtS�(�ǖ_p�Z���N��9�|u9᤬s c2����S����/�9I��3< a��>U��+Ḱ?.+�~ߒt�ϜΈl��`�򮌼B�5}W?��9�v����Ru�����@�0S#�K��W�b�Wv��<�)����o�ٕF�f�=�l�D��sK)T�Џ\��<&u5v��!��1bȰF�Oe6��Sdc�<�I��$�ɿ�HC�X�Tb7O�#���AVE	�V�8���f{�����O5�7��NM'���jf#]?c"�NTb���V���DޥY1t�e]?.Bx��G��+h
�"�8����Ŕ36����u�O�燽�留��%w(J��k�#iw�$�/�k1r��&�t�0Us(,�x����P�\dD��냥6��S;�#�
��]s_��0�7#Z�B��������g]��ָJ�}���}<��}���*��9}q�ׂ�\q׽�V��

F�L��	��r�Ʒ�~��+�ru�����q>i�;x���o�]���߻'�pj��E���U�r,�Do���Gg�Δ�l!%Ѽ�0ȍ���}ù����캝����:��9�;R��W���yRM���^n���F�U~���.����6�!mV�۹�UaM������@�ힴ^�*��R�����lR��\Ci����_T.§@�)�5z�L5l
7�����&w��\�>|��W���ݼBi�|�XT�L��E���b�V�:��``�a&C}�tZ���)Ob�z�<�fb��T��<@�\�y���W�q���ے����K�M�M9}�[�]k8�Q7ԟxjp��:��'�r��l_�ݡ�����lfg��i�{�z������gb���m��y������Q����b��2n�J;�w�p�\��8�"�k�^%Z[̇�Ͷ�w�	&�j�V��]xh֘Z�]#��u�˻��[�7L������PI��NtX��v���ˌ��7�!O��"/'����������3�*gjS�D.!v@�~�Ϧ�k�Kd��%FwpUm�ܰ�K���%�[/�����9�����mŸ]z�r�]��Ow��Z;�ͼ���P�Q�}F�I0����Jw��}�{ki��\����I��C�$Iؾ�n�}2�8E7�4�Mٹ3]˗\���JE�[V�}�g��	��^iç5J��m�'����aLV�uo�*��N$['+����j���gx��T��\�3�y0�DŽ=���)$�{�W7�uOL\�j��EC�nNE���\���q��M�mͪ�fnk�eJpvr���(Y��哵Bv}W�##L؜�[Ƴ.Ojƹ^�Е�Q1˅GK��G�}��֗}�_����u�Y�V��K���_sR��W����ɫ]zuZ�N�>c7�����Wׂd\�l��Pr�<[/V�P�:�v�	�ư]/Q-��Y��uG��ds����������8������/4�ȡǣ��Dα;.�Ւ䇅��E�D�DS��TdR�p�;w,j�j���@�bݬ�u@鴄�m`S��#�V�ﾛ@9�%ru�w��d��T�ȇ��ꀫ媕�������m�ݷ3Z�
��]���Q��Ŏ_v�������k�~� O+���T�޲�I���W���n��XS�ࢇp������=���J��q4�#˺T��[˄����:��꒱aO}�1%�%���6�'�������p���&�������k������uNj!�;���6n�o>�wv�-���ߨ{�7���H��=���öw͹��i�������|/��ܓ�3�=·�����]��ۼ�r˙��p�u4�]N����������Cu�e�yGP[s�)�kQm7�����QŹ�O3��ny��3�{�5\#7_k�9�kh;g�ͬu�T^O�)!]|<J��s�*r�9�թV�pʇ��'�_k�u�t�-u@�UT}%ef�a��]���I��{n��N>4@��Y;ke���'�	2�u�� ��3�ͨ�>�w����x+p�:��ը@Mg]��F��%Ś�ƙ۱��͔�wKL˂]�y�ٮb�n��>ĆC��/���ܻX\�f�$v��
B�D�fƵ�[�Dȯ.�'����>�U;վ~�1>�J
m��z�D�^B�zLo���������S�[N�L��汪޸םQ�f��.5.p=�$���t.������nr�����b�ć����kzd�K��u�=�9���L<�	���v:^SWC]��
�6*9sz�����O`��=÷��_���C4��X��(/���Q��
n��>��➘<���)óG���m>�I��U�|�
��4/�-��.��9xi�3�º���]�yߪj!k��>e�����n�XS@�jRyל�Ɨsw��K�hq�ۇt]|�l��S�kZ������N��2Q��g{���5�={r>����~�y��8�q>�m��6�n�;�B�r��4�e�#W˾�ih���v9uD-�4�2W��Ԟ�������ۖFH&mtEK���D���)�S}:vac+�Fu�d]W\:hU�4#YƔ�`�����b���Y׋���r؞�"�^��ع���I��ub�4�Z�6DC��<=b�66ܼcf�;m��P�s �5'>�?�-���=Jx(��4�~y�6���|'�mdD��u�^����hA�M���5Z�ȿ���xǮ��*��G�_��?����'���gz��q$7�w3W!s�9N#y�Q	�I0k��k�"~�DO!�-m@w:_C{ВI���Ш�M��bw�]H��9=i�5	�;P��F�"b1���|�
��a�(ю�ŵX��qy������9���18f��)�oj��ܔ1$U��G�y8��ᷚ�NUE�WǥŜ�^�;�2�\4��|��m����-f�\S��GS7_s��w?b6p���
cO{*��^�!�b�I�it%�Z��V��Mos���}�eAW>�=�~���]?Q�Z
�`<�=��Ԭ>k�:��s՟&�������.�0�	o����)�oa�uXEt�kK��.Sڥ;��we�بZ�[i�uϬ���	�r�8sj���(�OԎ�붭��%m��2Y50����A�9V��5��mB-�̱j��V��|Ӭ|[�����3�u12W�s�<W�͘^gWmV��}����5	b�3k)\=�	���Xv�����Q�U�8D���ng}�7�%�DmqkT�������X�OB�IS�kz�Y2F䗋����-������R3���������3���΁5Z�B�)����XS�ࢾ��Q���}=���>V�q_�C���8�������|�s'�Q��v�C����6R/���ld�]���=��i���Xp�;N��"�к~	��	�#s�yO+����SjSe��ܚQ��b�o#>��g��l?e���|QK<���p�v丝ܚ��t�Z���a�q����P�څ�MXB�7P�U�=[˒�n �
��a�s]�k��mL�E��|��t�{v^Ǥ��KrqK����������᝞s:*�O{�`��|Q�K�	�����S�WF�؎�ܲ�5�c�^�w����6�7�+�MT�%O8k����͑��
N�!��{��-:b�6�]�Ɗ���f�s�*g8��F�2�c���8�뼈�+;�e�<�^��3bc6�h�,���I��s���B�;��AeNZ��R��Y�^r�'�z����:BM�k�5n�nXLtA	�չ@��vD[)�� ��!�y4��[ΓKkwq��:�QS��t�*U��B�j���s\ڸ�D�u��S��z���\�vr����}��B�2>�J���*4��sF���^<�� )Y�we1[��X�I�Sp)�L+��Fzѥ�w�+'��ns�p|��pM*�
�u�%���Cd�=g5v൫�(l��;;���#L��Db0������|Î�f�rá�Q�'h��C�u������ek���742���6y�6��ܮ�st�&�`��%{B��bk���]��0|z��yFc6����w��A�Q`fm9@p�1�Dܤf����29Wak�����4�2ea���f�r�1������E�aFٴ�W#R����yS^���,��=�5�����{�Z���j�LR�t�%�]��h��3uz�<2j=�
�WUʮvU��b&/�ɎJ��/�+7
G�:9��qz��p�V��G�#�;V�ZJB`<c��E������4=7ҺTq����@nԾ���=Ʌyr�$��@�uKw�rX�ܷ��l�R��bD����F\�;�ӄ,��<SȻ�m���Sb�G]�c�^�TӖ�.�o�g��7�J_�:�A��n��kq���Y�G��J�Qc�/�z:0�х������>�*ك���6�h�j����:��tӀ;Rb�!��+���Z�����N�	�vbT�Uu{�.���^�M� o	���R]����2����u&�qZ���*}F���4.�1nYk!��g���A���]Mh6�	����䎁P�zy�T�[|1�@vd��X�Z�,�^U��:�X�����'�y��֌�n�99̝�N���=����bePw�Wu�<��!��Rۺ�3.��T��c
���ws@�mة{��|E^�#a��n��j��[��`��P��Y�a�T��{ӹX�d�w�MhWu�X���϶�n�'�S�^/h�s[k4v���z�e�ذK�=w0@�	.�&y��w�P��Q��\-$+i8d*j�5^��*e��[�.�����yJ²��SJ
���1�x�vm���i�����G��1,���:���ײާ������m�ԫlI�ƪ���͗v�n��:i1xi�!F3��	XyC�����'��d}ŭK�K 9>δ�wZ�vw���T��U�t�oNL
*ۤ��\j_�2��[sf���:��ӎо�Ln�*<�>�f�����x!��ǚ��ً����2��J�������Mܒ�� ��s"����PAEPSBP�HU--!@�� R�
Ѕ PP1B4 RR	J	H�!����,H�+�� P���IH�!H,BҠR�(!E#B� �"QC@R�@�4�A@4 U ��P�E
R- Ҕ"ЉM@W�@}����/y��w��S��M�ir��ث�drQ�bIy<�	�Ѥ��!(3fӕa!G;�v�.Ū(�ؚ?��ۋc������a��OV���f�C\PK��"�o��~ӱ�UV�lg��%Eb�/���8����>��{�yL�z�[�ڡν����z���=}�����E����U΂/K�Ϫ��]^�{�d/8�V���6�q��*q�{B�e�����Fӄ��P1�Q��t��]�!qsY�������-强�����I/Nt��J�Ku���Ƙ�<gU��!�"�#<��O�g�>�ʻ@���zsF#�k�^��y�����\Urd*q��!�՜5+
�|��sm�

To�L�mlV!c��Aж�˷}�kcU5/f��<�����:��)�W�ﷲ�!m��NB�R��EU�|���-�����}֎6�W����>~��wo�mEGI�h���]>�s���N�+U�Է��M+�u���OZ����f�O�B�	�,yf�;��ޠ��*��4|i�B�ٌKȦ$	�.R�%跛X�nR�}ܓ��B�6����S�o"����7��7��K2g,�R���Q���Σ+�X�$����]0�'\�$��ʶ2Z�]^���%��v�ث68U�H����<Ԝ��xX���l�����Ȏ�M��xmB\�Bo����`��x�Re��/*��q�������f����<�՛�سUd�r������cR�[`�&�]�71���7 Z���پn��Y��OS�Sc͌����o�t�W{S�N���O*�ٟ����3:e��B*�F��)���7���Fo;٧��}�w�ʽ��tKSm�ʗz(���f�]���͌�q6�����-�)�����t�ܵT��E�d�d&	~^'d��ve��eAۑ�MM��n�蟻�/���c=�w���q�R���)�X�,b�&3־c��W���gx!<��Ə^��E��~�%�>��Ꚋ�3h�����U�����%��x����i���W3,6�}�ˈM>�u�tc�Sp�O@�|~��/)M%ۏr���Bv�'iX����7�Y[��7A���2��L�Z� �W��I�}�M�<Tf�«�*��%�]Y[';��h�"ӫ�=�WoZU+���r��/�T�A��1��$�d૥G�Wb��FN
�5H�N_J]VO_��T-o-�o.���z�ES �����&ӷ�:?qO��O��v��
��D)O-���z�M�E�yAJ��l��t���Ϣ���*ܗO�E�寧���b�bw�:&�w^6z�)Ó�D7�q:�9O��
��=�=���=%f
����{�0v����ɕ�\q��ӛr�Y�W�A/Lĳ��!<�h,�q�8?y���>�[��c��6�;�<a_��J�1Ԏ�<�j��8����\��FM�Ep��RN�ֹQ	�I1P��vD�tD��l-�L�vr���ǭ����y��%)�y:5i�5�n6����DM��8T�n"[��=V�mY�=ݿb��4�[�r��S�]��يʁѷ�<k[XJ~zN�	|�ŷ��Q6�����ru{Iڙy>MSC�.Þ���(���o����F��az�m�iڲ����kjd5��emK/1U���v��d@����B3�n��f��Ӭ������
�d���4���U���z�Z4�v!ض����O7��!�l�:��mj$�\��vk���L9u���Q�;�(Ҏ���
���*���;�>�)e�t�yxf�~�J�L�=f�<�縥�Zw��,��h��c��dN.vRs](QU�@n&;N��-W-�����r�w}ih}�ۤ�˦�Ԫ���8o�Ch��q�����Z����Z�\Ci�uς�ߡv�p��X�%%xO=]tq�ݐy�D��R�=ո����oSOe�Ԏ��y����'��h8!o����R�.O-�֦$��t��o�U�p��y�v�������������>��7�;�,<��H�I�u��rR��j�Y�^�le:�Q
�c�<�^���h�+�����41�(�3���V���6��Ω��3�Q�Z��<�]v��e2�����	����s�q���ѕ�rj���8��Ƴ�U15���4v��T.��֔��/J�]w9u �7d��-���Mk���kC�Jl�j)෼�c�6��\�q��{�V�]my^>?<����#�9 *���4G1�whG�j�v�0��������TJ�l0z���_خ��Cg9
*�ު�����{���o�����q���ӗc���1��	|�\r�U6�XOj�vP����������|ک����]���wˡ����ZH*�]=ZU���[�χ���簬��e:5@ �Y��h�>��ܯ;��o*��c�>��"[��FL|��� �:�6,P�A��7�7)Fc��Õ3F�N�܍r8�^����/��4�rAf_tU��{��V�s]NiJs��ܾ��b��S�`I��^�@��؎��ss�'__�L_._6���f��t��SOBs���eΧ;e8�
~
��Yݞ�����cv��#���ۖ�m��=P�;\5��v�r)MQ>�K%��\��u������1t�`�����OB��V�7>*ʰ<-+]�jx�j��vOb]����<Y��۽+o��3�� J�{�{���g�a�(c����]�q��!�n��ݠ@���+��V��Z��;96����!�z�Ťv�*釪��'sb�r78�qt ��3�s��>}vTsS|n�Պ˺���X�w�R�/��lMto,��v����ʄ�k4�|()Q�%A������c4Qx�U��m�?�.�����JS�KZ��:���t�����﷕�?
yS#�wzv��w0���w��B���q���E<gi����֫���m��Ws\}������wqW-�>�ηثӧi}�e��ه�3y����V��Y����I�j�v����s7���)��-�fd��g�tYSe����C��Jy5�Lx��ˑeC�yƝ)�ʥ$���k�nu���[�U~f�cx����R9�f�q�x��kjU��N�ӆi7S�ȍvg�c�lAn�o����\~�g�L��4w���&���������$�CYU�f�0ot�~��V��c��Ԟ����`f�2���>S/E����H�Y4�<�S���-E���`�����p����wZ���Wj��^Y32�4�.ȸ���=y�̰�cct�X:#k�oTcAߜ����]�W�_ɇ�o�t�Ǹ��KF�t���)܅���IUjS���\kV�9��9)��F��Ȟ�勧wl�}�&�v�UC���Z��]��L�;�����.�ܿs��M2���ky����8^��8�l�P��ڬ�`2���ֹ̧.�]���jɺQ�Z*�$���O.����6�!e$C�Z�>�s6�ېM�kӵ��TUE?�����	_Bi�ç��j#�Uhf7���oL�������T�`of��r�T�����zsi�������[�(齄�[<����6��~	Imu�]P�l�Х<�i�z��9Q7p���&d���y.)�1OP�g٫��D���us���^>�}㞛��v�'���<��E�z�v^d��!u~lގn� r�[�]�|&�'�7u[����8��gp6�~snP#�.����=��B)�\�=�+}�˴NK���%ξ��a�
ٸ�Jz���t6�vu��&^3��)f���qlɐy�[[z�M������)
�e��"y�Fi�8ԥ��̈:2��ٴ���K*Q-�a\�%�Z����#�P=V�W�ps٣�����q����iv[���1����ׄ�f̂)Y�����*���Ua��_!^;�#�TH���g�e"�r��y��I1_Bn5¸NH��7
��(SX*2:{���;�=	ﱳ�\NU%:s�ѿrp�&�i���ؙ(�9�<�擧�������khc��έ{�o-�ں�S{x�34�Ik�u��v�qw�+�'z�bž���m�}<�m���^�b'��;�]t�M4�]�+q�G4�N�{ٵ����({񫓃��4C$�G2��k}�j����թM�����N�n5�VU�[�%�w��$�5��2�^ns�=��Q��L�l�UMqw�Z]<^�v�;������Tv�z�u��U���閬cb�jor�i�=�UU��k`�=�j��9f�S�b3��_W�J
���kv�5o}:��MUdN@�kT=����ֺ�XR������k���$ɘc�U���Ex{�m4����I������os7�"we���JHq�7h���×x��VA�%V<�;��,Ȥ�^�#6@������'������;2��PNp���
�q��.�vH��{!�xz�}J��\2��]�3AsZ�N �Cy���v;��>��Joi��SW!֤X�>�.ig-��aLB�x(��p��Q������M��~����dS�.^����V֯��le|꒸�}�&����w�u�c�w{Y�����T^j�IC7�r�ʇT�D.�t������Y����^�߇��ơ�c�bv�i(�_p�1Q���l�4�9�Q�jȷ��e?'��ě���P�"�)s�\��r�j|�n5�4��;(��j)�-5wЧC�6A�QnJܚ�y�kQo�ߏ�ޛ��!��no?3�>��FsAn8�p��k�'��kk������S:V�n]�ܗ��5�d.�s=9fMc�J���ᚇ��yZ��k"�W�1T�ɵڕ�3�(ąb%�ג�)�.u��[�r��|�Q�ǕJ��!|h?E��)H�����8�ﱧ��<_�(����3������]���P�I�GfQ�q��)���p�������O3�;y�:�ݱf�(�m;�oh{�]M[ojbU�d�7�/�/�bK�p�p��K<�8-M�@�C|�Z��Lވ`�!�@r����b��)gfö�-��ܖ8�a��g��vۋ�Z�����~�y�	�}791���|�W�����:��Ѹ��sZ+���FI�L��ݖ�*����l�}���G.oot�y�k��A|l��5���+��M��[Z�و<��U}%�}:�*Z�+�\03�0a�0��s�<��5��M��I��U�.§@�*ʾ��oGS ��%�H�ŸX���j#y=����p��4��M�b�����Elp�oa]t�T��Mr���ú*�-�R�\5�v>��^�t�P|xc�i>r�j��h"�^y�z�*fz��G�T�q{��r���ۍ�������6��gvʋ����S(p�]!�������Է��M+���冫0�s�:�^	�����Z4��0\Ǒ�֬U	�Y=H?lN�c�sǙ�����ߋ3�G�|�W����T�J;�@�+\�-{��ۼ����jR��,��'cQ��"K7ђJ������� �w�!<385e�9�Qr.(�Y��� ���=�ɼc�O�!�:����Н�r���t�¸S+Sް �\L����4�c\l���e�`����Ea��.�D7"Y�(�f��`�q��9)���6ˢ� E�!��/Y7�4;���1�h
�{^�zҍ
�S3DbP�<�m\�,��Lxp�6gTK^�׋x��90�0Dœ}���C��WK�뷣��e
���c�zXM�Y�ʹ�z(�%i�� H1R}k1L��[d32�׃b@��S��>����2Z���t�4U�YZ��"(��]$�m ,r�S޺C��z�K8�BgLdۇ���6&E�Ż�.�ݱ,�㜡a5���>�1\߻![��5���>�V�]V�Q��D��(r1�8��ol�[�]K��E��4eΦ�ʴ;���G(��ʰ�E��1w,U��+t�dJ*��#�L�QДΐǈ�w�+W �\���ّWSt�n�2\�0�����ts��
T�:V��m_V�#�ztW>R2�s�D����A_�^q�8N?t��|�����ΒY���_c�ۮ����a�)�6�S��1�2������T,�H����[�|���ZOrk����\��֊Ӗ�#V<2��մ��#��u�����zeXj�52��K�_ h7�z����t��h5���=3>�4�H�Nt��[���2�4E���m��a5Mݚ��{�6*�LO�`+�����NF��u�4�@�fg��x�ӗ"��'�7����65��q$&��v���w�t/�t��z����3aƩ��6Y��4�k�)]|������<�5��x���U-!�@�s���p���+��wP`Qގ@��F� �s�i��%�k`�1f��K��Dlٔ�R���LI�.(�x_g�{)�Õ8T� Q�WӧmB�<��e�>"�`��Tˑ��l�fV.r1��}rˠV��	,}�r�r�v�c�v���b�Xy�l�4��b��{��9I�m���d�Ȏ��$/9���gL(ٝ�1�]օ:-�\��V wo�������������Ij����z��u+bd�Gek�
{/��P���\S�a*ګ]��ʼ��3�E�����v ��:�����ǈ��Kv*lr[m���������$҇���Ӻ�vf�0�晷���w�H�J��
��i]�s��V+�p(h�ַ��dTu�A�����͓^�oK��r��Q�}�!J�[suZ5Ȼ��Ÿ!����b�(�P�c�)����qs���	����,��M��B�.N���i7�D��;J��K�i�Ix�S�h�F�<��S��j�X��{��t�Rl�����hՉu�]]���IT�@�<r��0rϸj�OMg��v���V��V����[*eB]o+^w�Duf��C�R4�H4D����ҁK@�����B�%
�!J�B�@�H��.IJ4�H9
HR"R9�dy�����~�5�5�~�w;�>�������J�`]��|kU�Ɲ�P�B���̱w��<z�e��QҦ��㫷82������r:�Vףy�P�T�BI�_6�]�q1�ȞAWE^�%��MB�v��cdI�.�Ŕ�V�˪��tj"ӆi7Z��vF/[�c�3�=���o�9��c$9�z7���[�r��T<��\�p&'/�dp���̞��ݗ[�Urr����IX2�9:��M�kO��F���L�����uqM�]4j�ʂ�C3k;�`~��fS>�d>\��!�y�8i}�ĭ|���y�Vr��ʂ�A�ז��X2�<^!�)ʾ��YO��a6*9sb�Z{p��m<Y�wi�z'eXS���U�x�y���)�����p6z����Yp�}n���|��w=V|��B����oY�g���'�V����]-R��[�zˇ��Ci한�Q�!!/e���/sc��>U%.��ԭ��)��A����ܱ���skqx;,v��j��Q�R���(�"��,���n\!`�o������^�A�+Խ�y��iV��O����]����"�T�����x��0�P�R���#j,�{%qz%:��%��@k��0�K\3z�1E#�6��r<E���Q@�-���)�}�T@I���W�Ժ�>�r�������mȣ�C3%y�L�I��i����)@.�8GCKE��.���y��ݑ�"�G�)\�[V�kLe�o�_��u�ʢ|43�zd�iу�ܮ��]��])M�t����&_��^YS`� [�����f�K�����,�e.��s�v���	�����\btBɲݠ�ov�,ڠZ���`�Pw1w2��Y5�j;�;MQ����ڞ�/r���s�W�af�s���C�򓵕|��Y�g��1y���[���6�g����6�\�ѧnzs��ݪ~#����:�f���ⴔ���ЂX^����\94����L�z��?Ol�7x�q���
r#3���`��26��pۋ�z��B�S�����I��e62^��N�__v]���3�ރ�/%��7|/�m:�'s�	�Z�1�n���*�brㅈ+���n!{�{���Q���Ի�����C�K֧8j��P��7�_R�+�������`������I�F��Eњ��F�J�,�@G�X�+�Z�R�2P�5=�5��r9Ӳ��Įr����U��gՔ�w���MquMiOs����3�j=J�=R��>W��F��
ډsմ�+��2ՌlW�S{->s�H7�G�K��\}�H�O��C�Wj��*�/�iAKT��_�Cx썾�tc"eG�����oo�*�_��Z�Pb�_II�]J�L;�Ȗ-	3xbF�A��}�^*q�=���<�^7v}�lO� T$�%��m��|޲����9:��[��B��J_e�Z�gφu�/a�%}�oLp�-N���I�z�J5r[�x��"��������:��uNj	_V��ws�U��s�����8%�-�	4�|��1M��7�HHb�4*�ގ�zի.!�*�N��V����;��!rQ˙m�nY�oF\q���zk5[�K����P㩎cp�m��5<�j;V�GsƷ�<ʿ<=�x��T����b� ��g�qM�0/G^:z7v��{���q�x͑T�G/�o`N�[y�D񘶍쫡[�lΙ�ۥR?�����y���E�����T�K�y1i�(㈎�갆�g+��Q������%����%b�Ӻ������ʍۙ�m�_&�]�7Q�����kh;u<N���������K2�O#�<�U�W���'������r#^�c��`�3�8^��սq��p�"�>����[�r��8�IތyT���؆d��4x�e��<���lfۛZC�y��r�vT�b�]Y�����K.��d�J��Ҝ�nr̿���ˢnr
c��tE����a:��{�9Yt�G��Yܼ�CX�#;�y�W �{eC�\*���mlݻM5m�I
���ZV�6�Tgaڭg��`U%�}�/��5O6骭�J��m����M>�I��U�B�*�@�+�˲	���ͳm��u�����(u:u<��|��1����Sm�Z@��zT�5�|���wu�]Q
��)޵�v>��br��j���s\��[����{�'�΂�1�#§6g��oz��̔F�6�{��z�����X�宸gf�{��
��ȍ�Vvou'p����5?r�����xA�Ҩ�񽎴LE*�Nt�69-g>V��eɢ�zG�%3:���u�W&_G���l�rwY�B��8��E@��G�_MC��p�>܆�E*
�OE�K�n��b��WM}�9��H`��T��ꅼ6�K�z����9N�'?��H���ǑP���"����h0S騕��9�%�m����֣1��w��z�k�M�M�p�ЍĪBz�ڀy�U��wo �o�����R��{�Y3/�{���C}SQ	&Cn5�Q�쉎Cb֤������l�[2c��\}������ߧU����Zp�&��CYZ��uqJolh�6��U��w>A?�Z���"^a�z7��׵n㜽��8f�Q̔�nV�������F��,����L澬�.yF�'p�^��{u[U�[휝�w��!q�������L���֨{9ҵ�O�Ϸ�g��G��R���p�l��NX�/}S�>~/N�;O�M��	�*������MD٩����V��9�̺�i	�H���~00�9�v����}1�R�0r�F�/�
B�Gj��8����8iXv�l��0�V�䯉�,���LhcT�ë���o��`���̏��/��W)t�h���7Wt�T.)8�F67�|�-x����3h�z�T'�?Vǚx�'����[O]zuZǵ}%�7!裏�W�����ȃ�C�L"o�j>۲3<�Ou}�NR�+��=�z�6���T)�v����f�]ؓ6{@R\�}%.��-��)�ڡux������b�,Juй�N-3�	Sw_oIP~	1	v��.��>�[�N�����V�Zcy{��`���Y[%��n�ڶ)|V
�������+�-S�J��q�3����RҶsZ�gpSl�C�s_"�H]P4vJ_<P�Z��:�If�IsV�������?M�)����۬F'v<��V���v�qn`�9/�r;S�\��O��I�l��ad6sr��[����N�J��֍������=��6�Ŵߏ��]=^'�B�v����F_ޡbI�L�nл����j,\�@�.񁄜���F�*epG��n5W�?e^�g(�>�6�\��!�J`�e�7E	ӓKn�Վ7i�}��@y�����"F�SWJ����P�tm�V�纋��A_��↿ymr����杨i�_��U�WkU�'p��i8���<���,]b85��e���5Õ�t"��)���*�@�z�������~�{.fg5���m�[���9ֻ�2���~�m:F�9�ʂ�?�Ft�r�"��r�1����|�qu���]�bN��lg���=�|�?�p:咾m��xzNw�b/��z���v��^}fV3�����
�v�<���ܤ1�b�ۓ���V�N�[PU����f҄�L�lR���O�Y�?\���N�SN���y}��u�d-�Wk���7���&�SgZ���^t�)|�c��V�t�F�.���ۂ������l�PC�_II��tRi�s�47��]�]S�Kr�_�m=�\ס�<�^7p,)_oIP~�b�_&P��_l>ø���_RJ_K/m�����g[b�!�%p,)﷋��tNl�*�����PŢ������\�<;P��ʥ�����ۊ>P'��)9�]A��=���r��3�J؄�d��@��}��;�"���P�7hhO �M��h���	��-Tk��X!��摆m��Nm��o]�}K_u��b��{�Z6��9����gYb)Jt+��\��T�-��Z�]xm$ҿ�|�8�	������o*��\�a��Ɣz�j��k�ȎjO�Q�Z��.�4cw�Y���4��1F�F�b!1�l�
un`�8�Q^oÇ��EsƓΚ�O�U6��7������H����̣[v�n�5Sq*�ٽ��[���|�څ�j���n#�k�x��D7���g��e_GJ�:7�tI<qz���VDC��sS��{�^�'�>�Տ*�Y��h1`H��q<�	t��n>/�c7ۿIX2�9D�e��
����ֺ�a�o����`�|�y's�xv�d��ݕqʛ�����o�/� %o"���K�>0Y��G��^^o�,�	o����f�>:�W��^z��uS|��*$�Z�p����{��6@[�a�h1h��ک���mLű�#C�	�w��&���a�;�m�R��!J�
��*�5Q��-�e�0��e�N�mM+��ƕ�+7�҆.Z�4�5-B�8;k7��ؐE>��D����Z�q��72i�9l��yg����~��[U��f9�UD��9\�y
�̥�}w��
�����X��C��\&�\:Mp��2&���g�W�E{1C���x����Dn��Q}=3�ͽ|���&��Mą*� �0UT�sK��v*�1��!�ߺ躅Kf�R�_�k]��u}o��p6�yV�T��n[��蠚�z`�!-�_ܵ�ӗ�h�휥a�y��,��¹�neC�#=nZ��̈́�T�"�ˡ����]�����vpEپ��v�7z���h�jX�m�W����3��Z��y�"�CW E�Lt+1[��h_h9/�Lmr�S|�pu�\�(��	��hi�*�[��JZ;���ɯ�V�r��؄���Ш��dLr�NJc�p곣���A��]�B{�x��=��z�Zp�nl5��{��A�\ё=�����x�9�-�߳�u�J5��,�����
6�6��Ю�9bm���ux���m�0/\1�-3~{�l�K��uc�징���kuy]��[ 6��'n�F�fX5XY�}I�x��3+n�u5�dÜF8���e�8TG;5��G�[6���[��������f��K���qsG݃sV�Qw�����;O���LY�b�4\����#/jV"�h��3Iw���ڹ�G�mB�7_k�U�x�&�*O1�gA�0�]������n/V�
g�/__ɭ���o�K�W�<���p[����3syj�q'au��Cϛ-=�]�p�*�õ�p�6�M�s��Q���{�K[=w�g�ZB�Yp�}p�]���#�<Q��~�Y�y�1Us �ݳ.V�T�[�z�z��.��+�=Ikot���Zu9<�p,)ZIP`>U%.���R٨R�m\�C��������xoc]ig�N�����
�&(%�Ժͻ�]QS-݉�Y�϶T�����ۉ�u[cʜ�D)��xD��dG�v�7�=���q��zI%lt��'�T�u#� ƜHM��wqЉU�F�{YV&(/\�lD��%x0f�}G[���3����,���������ko�%8���pGE�5�������S���g���ʝ]�:4�v3r�B�ee���157�0Z��`����}De��klne0M>Ԡh�G�D]�a졸��t
%�
i���f��_�j�Cl���t�D΍/K:uu�_�5�K���+��LB;υ�A�m+	]�4�4�(qU�9�I!Ͷ�*HH�n�[�̊�x�%��F�Z��_jyѥq�J�x<�_m�ǪB���ܵ�ʹ#fȹ�ݙi`�0�����s�$��$�m=��ǖݹ��QV��z�#&��hKܛZ�ى�DL�&��2�]gZR	��*�ݻ�ػ�=�J���P
s[3��@��V©�A�gkM����3�<X1�A.���L�4��9�x�
��`��A[%&�b����	nͼ�9k#4N ����zƮ��ND�:�<����v_>�E�}f[�C+5# �]���v�Ws.^ͭ�_>L�0�5�����3>����M�!��/y�����<5*Kػ��+%�&7o�r����:e���MZj'H\N�ñ�o�S��uș�R�J�r3�U�b ��0��ܵH��/%�M�����jÂe�)W���I[Z���{��`���F�k:��,ej�5XNB�n���l�.�l)�qPv�2�G��b����N,���]��&�T׷:��')M��0�L$�D;5֌���ZK�-[�VnG�-�j���m1R���ktZ��}�t�k.9���8rxÚ��)�q\᭘�U�q�`�,�F�<��2�¢3�8��;���h#�]�ׯ�tt��Y��S�<���f�ƸT���,���9J&��tL��B]��N�;N��\�&��s��a'7�����uY��'VN�s�@~��ҷ����j�MI�0o3�+8Yҏ\�;l��48�:�lU�5�����jA���Gw.P���)*\r��2VJ��8��ۖVxnb�n�R�=-�:6�Z�G Bs���I��������j��k�c#o*h�a�aǜa���VnD�']-m��h�(R#�zԙ�]cYl��KN���˺9�0v+T�����6_p�6p��}[d���+(�C��
��I��� C5Zw|!����\#�L�Gc%���}J�t�M6�2����쇹=�-`��5KnU��鹡����پ�$��G�U�Б�Z��E��b4p���G��4Y�n��Y�pKU�������BK��3���Jw][؆<�b@<�Ƌ��n^�o�\|��&�t/z6o��b�Gb�q�8(���$t���th�|��K����Ghe�ݺ��ۤu�U�{����$���Ӈ��ͼ��G]e�@�'%�r$b9�ZG&(�k�+|���_n��q%��n���펡[�n�"b+ �(jm�$ӯ��:��G,�rE2(Ak$@�T�
X�(JT��L�hV�����
P�(�i �i�iJZ��rJ@
�F�)Z������qlf1j�p�౗�v��l��U5o^�ƭK)b�؉�(vkS��fBzrXܨ�U����&��*��E�%�y�,g�֢��-�����+g5�gpSl�C�s_"�<���ܧ����ғ�����591&��i.j�����
�f�aR&6,�U�+iR��UN��|���@w1��Wd�v�_.A��w��q��L���mK�Y�����wmU�8{DO1� ���}�þ�S���}<���E��-z��Q��(�p�.9���\]������3fu���"�>��sy�8�����)�oj����:E��ųo�Mj�]�*aZ�m@�Ɨ:���D��i�5����{�:F�9����W�\���%�糩`��OOT��\Fs���iڙM��%����_geQ͇U��#��쉕�]Ыp]�}Q79P%�}UfS1ڧ�K��sZL�ҏ S�L���N<��ke��'eU�7=�~T�+�-X��-M�v�k	���U�I��]����B��%ƶ���W#��b���x�c}��=�4�M�Ô�vt�ۺeY2�Xp��>2$���q%h�¥;�E�� μpƹڕ�:�db��eZ�r8�(�.����a2Ȃ�n��(��!�-��J>,���	�n[�6�'8�%Z����ÛX<�JE6Z����h���r�r��(9��o��{e_+�7>*Ȅ�p��=[���I����S[����5�C�y�l�n�XS�ޒ�@��f>��(�C.�Hs�;�޾<������e���k]��u[c*RQAP���+W i�oNXm��|W�1fz��G��w�_u�ҿ��{������vs�P�jQvj槚g=�o+�y�Z�TY�Y��B�P�J�|d>�Efʷ�O��&]-C����n�R(3��)P�~+\ԭɨ��P��w�����99س���\F�¸ƻ�n&!<����Cn`�ɩ瓯sc�]/7�.8���®��{���j-&&�]�7Z���:`Z�t�P3"b��x��S�|�����k��k���N�x��7�_k�z�X5����E�Ћ��,�S��YJ�x�.��7n�V6-K��X*��\j�+N\\�O\�8�������ٵ6vV	$AQ���s���ٓ���o́���۲���;��sZu3+����ڪYJ�Ʈa��M��EHB�̅���Z�*{�o���r�\���yBf�7"m�z�fw9Pv\��.NE��GK�oQ���t8�_W��3F���w�ޖ��^V�T�i��w�(�kz�_f������뫝F��p��$gy��cl4��p�ż�/S�zY=o���a=�c�[+���e�Q���䤰\K�˛�|����}��&=W�y|��4�� �a�	����z�8��Q]+�kb��4�C��*�R�tH�xi�^�w2�,��k�Z���.���k�{p�5�C��4�*m�����U�9�M.O����O�%�t]D*[4�<�kZ�|3�ΥF5?^�Dn6}w������})��'�P��^�[��#ؼ�k������ui���[����q�ڇ�{2a�9UO�/����]�r��}�����b_�;��
�5"����N�e�ґg2��-WmES�lX�Pލ�jW!�ۗ�8��8���-$Ws�Q�f�ծr�oz�H�abn�o�e:�9X�𐑑�|��cWE��ze�s�Q������Y+z���g1�n�l��4ru|E�kp�܏+R5���q淁�
m�T9�4���]�@�E�RB����6��s;�˵ګ�W+�)�:�!o����7����Ѹ�HLu#�8؝�s@{���t��^�-l��/�j;^�0�ٞ�@���kB�5��=�,eN��wS��.j�1֫��Ove��{W�WM.NK����� v0�R2j=��3R���~�-���mY/k<N��?\��pԽ���o2$�t�u��Z����؄[�*�l5Sn{�W'��:\u������v1�J�9����|�4���鋓Vz�_f�9e�������ljZ唅PO��OcN�L�c%�����^����1w�U��C�&�;/5��o�=�ҧ�$�>��8��bb��b姷�͸ODFv��\&�n����F����2=}]�5GB��G`KOT:��Y�Yka�XV�0��*!��cYG������38�UC	��K�:�M�t���i��U����n��3Zp]�H�/6��[8�(��+F��xF��!}L+���U�+�Y��h7�����a}G|hV����#�]lJ1{ ;r��>���VoL1nች�iɇ][��H�R.�j�S��0*�ݳ.VµJ�kyp�7�����v�c�|i�5?�7��Y����8/�-��_]P�l�������v-���[�C��c��8ާM���_oaPBLB\�wE�W*��|+8ۉŅu�O������}��q�m�s*R"e?�υ`�o��e���:I�t!OD���7Է�mKJ��k!��_6��:�5��4vQ�YÜ���k�]���5���h��|�|�x¶o�j��{}4�V\3e���W�Z�Wd�Gjt�I�I0޾/(���W9��}��^:��R".W���C�l��BV׼s�<Ϫ����~�ٍh�>�ڽ�t�Nޤ�Gsr}�t�ޯ��SQC]������r;M����s�;[/��w�{�x�g\yf����iz�,,	;�9����%��E{[ܸ���3���Q����·+��P�D�>�w\' ��b����Z�Ύ�st+#3��j^@�r�mkTEu��a�r|]ײh�#��p&G0�3�����N=J'v���M;��,�
U��R1��җ�!�������5��U�.-��nv�NTuyu9Ԯ<g]n��۝�۬m,��b�s{L��sQ��t�:p��siPjL�!��s)���Q�����m��N~��W_���MAŘ�-���@�C�S�tI��scU0*/|�<2S�x��'걽�W���oG{s�9�˕wi)�rϣœ���Z>fp�r�@�`-t����r�g�.2+d�V���]��5~�h����mO�,�R�3�>�Gz� �	��������;�[�4���Hz�e��!��<D��-��w<I�Q%x����{�\	f�+}�iV'�׵W:�wU�m�O�i,�^v�ϝ�q�%e�!K�<	=Q2��)�����1��ی;���{���̛�ܺ�6��b�������IG���-�]y��AF�1Ӫ'��d .g݂}ם\��<�5�=ǅ���n�)ˮ��K]�>}'ǯ�}n��
v��=AJ����̖1�f!��FA+�s!a[�Zd������_�l7]��s�hN���K���讦%�ثd�C�|�,O:�3K�h%q�����D�{�*'&D���^2(m�К-`�E�X��|᷻��!����#KrQ�������t����������˼�.t���'�O���	�5k��e!���eJ�)��{x'Z��4���G7(���	2[�l�Z˙�:��cAL��4�)ڶL���e����>�M�N�"�x�M2�z��$l�+iѱEi�^�d�F>�s���wN��z�������'���|�� ;��`�o����`e/~7F,�hy�`���{�G��S�I{h�gt�9�G�UTtgKdɰ���x5Q���2kM�:�dM�M{�=�3|;���W���q�V������P���ϡ?]���I�l�O_�{g��͞r���#B�������b�d���kC��i�t�q=�oSΪ��н^�����<�Ĭp88���nf=Bu��w�>���w�8nd���z��a�O���.��L �<��"U;�'�7��|���N\e��h�0OqW0<ӷ
&ޏ%��'�=����M��:0��Jngތ�gmVm�����t�I؏]G59ΐX�����vOQd�g���@���U�gZR�z^�u�E��k�<�c��/|-�L�
}cہ���4�X�I�=B�׈��xoo7�1��~����RT��󫅑��~�����3��a�Y�B�,��E�u��������zy�Ѷ��l�K�{4'r�S���jLnp�2�E#ͱ��@�6Y���(�m��#Z`Uh(�B��[+��-�cS�T�ON��t�w_N�"�}Y��R7Z-F��cu��GR�jo|��r�Mn0�[&uZ��|.�s�����@H�Ir�G]ԣp�U����~3�!�c���;&�=޼��G�4F�w׽ku���d�Ӥ��eDH��LP�jqe�O���-�������+D����#(Nz����t��^���[��2K5�FoAE��I�y���Aq���Qk��#<�ދ�����u7��y�����C�����u��ثs%�B �x�r�p7 �>��t��g�Wl��ox��2�Y�����[g>������}ՠ߽��.��j�S$���+���c�#�g&>�Q~�󄶖hW�w�F猦_!1�ڿIL�%��d�qSh���*v_;�fmv,���ᱝ�=���u`�r�hX��j�ii��s��}wD_�'fM�,F�������93j��y�2O��]�]	xb�������7���j�	��B����=����|k��Lz�.����
���%�,_�mH5��U�}bwL+��V�R��lr��y~�������g�a3�s�ְ���a:�؝���������ľ�uC1W���H�`5*�ơ��;��"�Sn��5��!�嗛X,��H�GjQ��d�h���l;��K�o{�x��FZ���Rs+[��wy!5Ҝ�΋]J�����u2�$Q����Ku0y�Ք��5�ֈ����ܧ�6R57�A��O��ƹ'e�kO:G�>>���W����>u1<�}����I��p|}bea��м�]�̊�04'w�<��_nV�^l��W�diP:�q�
���O�γؚ���Y�����_9>>𾼳B��Ә̽��c�&xz��ttI�S�vX
ƻ�6�K���W���;W��z�j��R���e%��/ҍJ�x_��,I>Gc��e�頬c����Lk�����U�z��j���a&U��]�o�gI;@�L��z�]L����
x��y��z�b�@v����+7����+���{�Ǹ�K�AŒ�I�2�������{��K0��nV��v�]�M]�M��vS��S�il�9���n=��m�]�{>	u�)�,n\�=����n�;���}}���Xl�+��W�#�zg|W~��\g�dm��F�L�F��¢�b2���Ͻn_-�OՀ�+��>F��;!׭"09��G�9��6v'm��5^���F�J��%�̟FԐ��QSSB����#>�+#�W��z|��������Iΐ\��j�3�Lf��<}�\�(��JSd�K����������*�E]�������l�r�T�%�Ų[��!�SV�m��I����WF
j ���k�6��u-�\��'OmB��YX�Fǅ���	sWo[��ov����65�r&JNk=��tǄ7}Bk�Rv���݈��*WW��Qkf�u1����܉#�_���z���_�u�+Ȟ��e��>� ����5�J'j��e��}�c������z2*�������V�{F�5'�c�鿟��q�4+�u ��{A�������[��Æɚ�U��G,�=��k�m�ӛWP�?]����_�ۦ+��{�����g/���G'�M{�j��#��p��>ƂS��ulz�u-'N�L�m�I��h1K��y]ī�����<m��h������x��μ��{�CgGI�:6*Ux�ϵS����:���;�z��g��c{��=��D������}��1��T�p�'v��{(O�b����t�l�:�@��\��p�o��9pf%��3�Z\�^�ׇqϛ�B�V���R�0���z��W���rj#�P�hs��U�le�=���9��Y�#�ܧ���1垻C�t�5�#�.x�ƢJ�L<�/��흞S�bL���Ѯ8[�e�9���4�~/Ie�:	l��S��Y}>���ה��K�w�x17�o���ե�W���n����U�5����� ���.��B���+��g��S������J;�r�.�S9/T4��
beg
�9z��I�Ĉ��쳼��.vK�Y�jóU�;f�Jmo#�5����r��rs���w)�ͬ��#f��CP��@o!�;��lʖ0�k�T����-]4rN����4q���_�`�X��\�)eRX��D���n-{��ݳ-��s�ɁC����|�α��N:�Y��D�[`���h�C{K� ])�h�{\�:�={�����1�#eauk� �8��IeY�ҡ�@msT�N���\���0&���ig�o�-�ص��$;�t�҃*��a�0���͔ƅt�իQ��
����� +rM���k�Ц4�-��-��z��8T.�5'X�)9�M�t
8rI�3Ϧ-��q��i��%ut���4�5��]�n��)ٕn���+Mp챴�k:M�J��R�X5:�1�&e_"��v�9�5��jkg�(��|���ss�S�.��Y���;���wzN�n�Ҋm�Bmefj���>�ԩq�L���bIy�1�F�NC�`��\�Ʋ�EY��7v�uҡ���ZǅޭE�8m*Q>[�[��B߼Ҟ�����.�&�4�!��6fR3��RD㽌d���u��n�ltS�vM��Q]�r��;&��J�h���Է����*\d=5��,�Fa�vb�2l1�;�J��>�	����Y���J�u���_�n�}lp��^Z�կt�o�����D"���Cv"/9�r�4�ʵ�-��u���N�Sm,Js��W�"����jʙ��{��蜼N{�s��\�I�J�QU����Mc��v^���Qi������L����z;�@#�A�>o�_ƶ���G9.Ԛsj�y0�H�Tn#]R���rCf�췥��}�Z��˔�vP�j���
��$��}%�LV^u �Ho�\旆���k�/53�+oc�v[�qS�ܫ�O�(���妚bK{�(���O��|����KRlc�l���)SxT����t��i�2R�k@q։m�鯡[���VHe���f�X�I�E��b���@����n�Q �J�ʙ�+�N�d �V0rԓ|t25v�����E��n��Q���=��.��˷87���l�#��n��Aýʰ*�7wi��V`��=�ڜ�:��F�-]iꚡNt��+kn�=b-�kW�D�@k�er���4�����B���nJu4T{F���"U�Q���,�������:�拯f�E���R!���9J���,�wd�⸑X��b��kHD�K����%��J	�wF���s�%*����dN��V�����2zf2��Z���)B2��Q�͋K�Ejd:G�fw:X�@;��e�����k���V�gu��┅PRJ%{d%(Pд	H-B%- BSd�dD��@P	@RR�!@ي�T�%4�B�
��IBR�JčR�%!HRSM ��	E.@@P���P�}��F��1a���Qu�,u��s�+�-��η'L��68����3�.�f��Ǖ����T|�-ˎ���F��l��r�����3��.��Z��\���%��^%0��Üe�r
,W,񖯶k׮���(���@EA�=�bƻ�� ��E9uу��[G|��Y�T^�Je	�X�3��S�/m^'ƾp@�PdL�IJ�ϑ�����D����Nu�q��'ELm��^�}���▒����c�݊���k�D�O+��d>>�&>XG�k1;��w�Vr����g�r��d�f}�m��[�bh)�3�a#`옙[N��Z}L��"��oˠނǨ�bc}	����{ԁ�W��f�
wL�,�f_��bnydS���V�I:����N3�7�+M���>��61Jd�M�G�j�4��<B;1W�Q��d�v����lg�*V������Zo����N�H�&)ɷ�b'l��Pt�q��Su}{��͗�I��2C���;���,
�ZN���J�ۼ�^�����#���(�M�SŔ�'&���]{D�7z,_^T�>'v�3	��wL9���u��`��~E�\���Z�ۯŕiU�ʏQ�j#��Kgt��rE����SqR�z�йꄦ��K��:��^^_�p���)|t6��R���w�XtZ�^�<�qD�*������Le�:�F�ĺ�n�h��e;�v��p���N��J���F���B�\��t᭍��ܨ����']ⱪ��s��yR1Nf�f ���VUx٩L�������%���Bmw+�`л�ȸU�^���]G58������Ʃ�=\��6�e�=P��U.���m���Z�3�˗x�;,B��O#̿+v=��X��kqG)�����=Cq���«�N��3��2����9���@�_zh8�O�y%����/�z�G�Au���M/z/:����7�=i)��k�=|��b��T���J7
�X��{���#�z��t���N*��}e�l	��ޅ�\k��dv�(���'�Q>��LQr�N}�u�v�t�z�����Doa�u�<;ϑ��:>=x�����۰�FIf�0#z�2�)V�d�=�Ƃ��r�4�m:�-l�O�t�Ξ�W�����ב�~�8����m��ث�̗4��$\�\�Ǩl�ﾽy���{�[ռ��~f��6�����;H���ϋ����E��f��,R�h��[�j�C����=�~����{��HU�Oqѹ�W���*:����M���,�s����DP
m�הOH���-�;�=·(��Ũ��DiN���2.N�:{)j�X;Z����{B�����K�����0�R%r���GX���\|�/���ԌeXgs�C���j�cc���.:tԞN�odO����X��8����
�iS�G�aɗ�[�I����2���X<����5.���K�G��UF^�'���z��|��[�z�O�����l{�=�IC���Ʌ�%኉koF}Z��o7���j����u��S롶�ˡ�UFo��g�:gжX�	��{jA��|J�0��N�>�ñJ_-�~=y��kʶ��J���e���5�<�^�=���	������;{"7X����P�'��x.����Cq����;zY8{����Z�
f_��ΜsS���<���rNipp����pSuZf�Ϝ?kx6}�=�uR7S>d��v}��a��Q8)Kg�&�og;�E\ϣ��kS'A��vd�{|�L�`%F�O��^��8vX
��������9�~<�Tf��E���MFl�o=��1����Ƈ�K��e<X��g��u����A\t��:c|�3*9���c��}����p�҅Ц��w�Q���'h�^5eS�L�n:�)�<yb��[�9��#����z;5�1�'���a�j��z�(�:I���B$����2�V�������튝��3b+��b��;C�l"	G�c�ŧڋb^�Ӎ�ʛ]+Ƿ����W�^/��Ҭ���UJ����,u%�k�(���+��]{�a�Ӻ�ckU��-�"�,�6=5����:&K�ku,�n�1��o�6��/D�T���
��Ny���HҢ=��m�]�{�]C�)�.#��:f�V���Ep�>�ٵ�,8�⚅�S��V�a���������썸�ճW��뮇{ӻ3m��s��]x�;�5ׁ��|��T>T�)t�	϶�>s;�m�bvv/�^���2b��[3�}�׾Zhz=2Q�T��c��SC")�x����#_�ڿ2=>V|yUm'�^{���DJ������=�j0GR�88˓�"ds��E	[N��Ew��S����0�^S�}=Ǧ]��.{y�1��%`�.#Z���\���Q:������R>՘'ԇ~�Բvzx9ks�'����k`�7N��a55'��@z_��i��\w�����P�����{�W��� ��v�ڋ\���;��yiyח��~�=%��b�#�찇�f����v=�8�4QV'չ�{O�?�:�)��U�'�oK��w�S^��~�^/|��W�՜}�:?G�>��~�V��ױoK������;0�)7'#EOS'��`(�����t��}9��^\�U+�#���=y^�͝�oM�������%�.wB�1:ˉMP�k�v�)Ԭc����0uD�\F^NchE̒n�Kv7lPO��e7��&�é���tr��eJ�K�}vUbV$���p�4�pcGR�Z���j�rh܈ǻH��l��Ν"sV�=�
~��Y���Ӱ�'v��ʁ>E����pi�Y��`R�h�Q�g͋��L���i�hR��G���8߫�ǻ�:n�'�Vp��V)�q�r|���y���NK�g�0\6�G������ϣ�hx,�����#��'��%x�U��G����7ۏN��n��ԋ˟�/]P^�/d���A���W�d�����<	={�4ו�^�u��=˖��ʇqS+҂���t�-�~,>��ӏd���Az�(o��xn��s�d#
�k8q��^�h:}� 6����PnPWR�W�ԅ_�ֆ�������o.����ث���Tk/5C�Aު�c�2O�|��ʌ���[�"�%yN XI��2'�v���n��9uQ>�dKY�~�{2��?D7K�{��>�TKfK5�.I�����g	W��Uk�cg�Wq�\��|GG{޶2=>�O���2o��lE�n��S.g��F��1?	[N�t1��"����:w�ޚ���Zbcy5~�~����z� �dC5�:�)�3��3/�.�w���Ƅt��򔌺�4S[`җ>+x�� �����A<@���� s��We�7e���z�S���N��*J���SW���GK��vn���얅��������f">�CUG�颶��8s�����4�{P����*k��;
59�����Z������o��zo����UG��/�ɿ��@w��j�q�L�V.��s��P��>Kч��8����ԭ:.+�m��ex�]yag'w�`�b����O���!뽑ᰭeEu��溳���C=�p�"�U&���*}�E�'\Of�(w�m�C��Op#�9�n*������Q]�jW�j�J��ދ�á���az��wY^�%΃��� ��\�o^Iˌ�ܠ}�}���^{��uN�n��/|�������8��\������y��Zf�E���n��8���
1Ւ�K {��j�Kޓ���� ���/T읱r������(X��]��{��F�c�}J�OQ�e�C�Y;�)�^����Y^W�����j�����O\#�Ʒe�e�&v6�L�9'�D�*R�W#]86�E���g�*}��b�z��	7s���7^��g�gM�Ƀ�e�\XʕHuT����V*�z�8dG��1��=��V6r6�;҆�ϊay�[�V2�Q�GI=DX��LW��]8;.���o8P�徝�T��T�;��z�$vU���!�h�4�C���v���݊e��m`ؗJוo���J#ǩ��݄�X�e�W֖5��ׁՂX��Pi}h����CQ�Z���ʈ�#����M��Ҧ#n$/��aqwr֌y��'6�B�փ���W�rK�������^'�ПR�[�GJ��:�>6��#$�A�FB%*�l���Ly�s6�c�v6�k��)�����V��t`S�|w�:��m��Ǭ;�b�%�� ���H5clֈR�ӳ����v|�3ٌ�|l-衶v���}������dF��f�L��&WpQ³ק��Q��̩�A�"gUxT��#=�S6�������r��a�d�&��x�>9>�����C�r��f=�Y���j.���v��߻�v�"�m�̕P�0��Gt���T�	��%=x�F�񡂺{�\Y;Q��쌕޽Z��ozX�]�b�EC����G�VOGU����ܽ#��L���N�/f��b:|J����W^��t���~���=6y�I?_N�({�	�o��y���P��ՏWK��Y�#.6Y;Q �~7wj���Z�Q���=֥&��T��>8<瑿�֭��ts���5t'ly�6�x6\:���q껉���j���>���ɝ;�L������x$β��R��	��9߸��w⏸~d���>*7of�=�ʶ,f�κ�㊱�x�U�r]��Gu�|��]��O��7�d���������m/P�V\�QV�G\]Q�P�` ��˫�rw[L��;��0�/]쎭b�w�v��*fҼ�gF�mj��`�ޞ���>ܙc��'N�L��OeO���yO|vX
�k�'K��%R���nl���|�����"��m{�X�>�2,w�tݔOu�eFW�gJ���#u���#�@�_�k�B�E�B'+̓��+Q�}��:^+>��AͣmK48�3Ơʦ.�R7w^�;��v./c�%��nT�֮��"�<�z2Ķ|�L?pn�=8%z��(��%Q�p&�Cי�z�}����+�"�y*՘m�e؝6:�ثT���jKS��Q�~�R6���`8K�r �9�b��^��sj�����p7E\b�G"���w�Y8�x�c�n�zú�k���ا�+�X>�Ô���� "�2���p0��KF��;z�1����;�~��C�ʞ��gN-[3��_NW���wp�u!TH��Ʋ3��|v�aT-�#m%l1ߢ֯}�R��|��{Wu�)x�㳾%�1p5ۨ��F\����/X��/��n�[5.�=�9�9���ޤ�[�>#F��m׉�@���C7�ԃ�Y=P���>ʊ�}[�g��}!)��-�4a�P�MLۙ�����A�3�B��:9�@�2�o���T��:�� ����kT� ��݅E�Z�5��rծWH�����R\G�3Za�ʹˮԕgk�x6�Qȵr��"T��ua�n( ��<'���+BQ�u���Ftm���\��j��p��Oo��\��~�=/��4��o�� �)�*����a-�!��ȓQ3;�+6=ڡu=�Wi���#����˄�����~�=&��LWg��b�l�p�	�ݕ��x�[@��*|=@����C%K�|x{e3`fڰԙxF���ex>����3�Q���cʶ�[���h��fp�,�������l�w9GE�T��N���<��t��ixS��J�\�c�7�;��xw����W������|N홇�'ȱu�Zn Ӡ<�m0��79f_�7eVu�!���M��;�����J�����c��7��Ou��
�:�2��oz�n<�f�K��Ҋ�n�C�}�"�����/�ǖz��K�B᭩w:I�BO2���
�'�ͱ��k������6�P�f֫��K���_��;�yNG�ׇdD��@8K�i����𧻓O�g�3�O���]L�>��Y�n�U�ӿq�)>/�}����p�u��V�}�a��^��k��E{�p5�@�FX����
�_������z�э�������Ȫ������Ύ�gd�J;���JT."%	)۫�qd��ٮ]�"f\�į�e�FQPv�Y�Y��Y�VQ�O��e�+^c���NPѼ䦭�;�e�zX3)i� �+#}�N}�����Hh�[����ۖ���e�,���É��n�L�66 _��^S��f��( r� z~��,��9��
���=aFw���n[�z�Gk���}N+q����~v'M��݊���k�D��0W�����:u��T5V6o|�r�>��N�ГT��>�Kpr:�����ؚS.g��F�ɏKu�����~lM-�G�s�j�u�f�b��W�7���@�>�������(ә�5�=�D%�P}��8]�l��*pT�բ����o����^ۏg��c��d��ޠ;���CWAe���v���2}c����_���ԭ:'_W�����ˇ�'�1��>�5��s��߸����(U~����Ei�7q�*�L5:}S�:.):�{#z����x<=y��åZ��yg#_q|�+�y7Az^�U�W��b��Tḍ,��3�wL=��q���փ�,ߺry�k�JW!>��w��3�U��|���Oάr9�{i���)�;�a�S�1��|߰y�8�nڪ��ܼ��Kd�LX��-W�{�v=uԿ9��{m�;'��ġ��h����+R�S�7yv�����ƞ��c�1�6�o��f��fe��f���v@�q8��{ʹ��Mj��y���7��14X�x�ð:�z��z���w�H	�����}e
|-�JԮ��7wە)Tګޚz�@p�ͺ6���X���®U�p�1��63!%J�V)�V�b4�Z1Ӌ���n�!C�,���.9yw/�5���;]4��'�о�vS2��vX䃲��>���IP��՜N�[���7��K�Vؗ�8)��w-[ֹ�g:�7D����Kn�*{(�P���V��śX.�)ݕ+k\���RZ���qo:;���#!�w�Je�����'xr��S\�WP����p�]���U޳ ��̹���u�����JY�̔"��b�]"+,���L���U�����|���+%`N����#���U��ƭY�IwT��ֺ�CbZn���-��7�N�AM�i�|S����Y��h)>��rz����m��+xl�\����\�P�F��g�:7 ����& �#��:6[�Rf�.wu�R�2]�2.�S��hO�i�\�����y��r����Q��y$u��s�wfQER��)H��D�ͻ��9.��zvA���]�C< ��ټ��ڶ,[�Y��sz��:�E�O�uW�����HE+f�C_3�u��ʏ�s|(�*��٭��yYO�i���*�usi���[7�!wy���;�� ����6!�Zl�Be�s�`��1�O�n��wF��GRv���jb����D)!�����Vo_U���v��{9٥un�K+Y��\q1k�E��f�ԇe�!l�H�{$�ju�I���qѐ�2����2uGmB�b�و�+#��Nb��UʕC�C�&ֽ]E:��()F��k{3k�i�a�A��c�l�ާ�Dn)�+Lg�v������\��l�b$M-_.��q3���a`�8��o[S����ɲ�y�Ȕ��Ch����یޫK*��A�#]�Y��3d��d��빖��6l�9c��sx�wT�H���ޒ�m��Rñ�� ]j�YA-����X�~�ұ�"��٩��v#��ZֹiK2�^���y7Wp}g�x>�S�Yy�	��i�F$�j|x�bd�;�Ԍ�%i�ٶ7z�W��;�]�h�v�^�׷ڹ���u3�|�T�}�r'�p�uI�0n�qu�r��=�����mt�:�:&걲�����3��Flē�!U���q�;z�v�X��(�����V	aq���4����;��b�eKw��,��ڌ��d+GG�Z��O�1YkL�՞X�˚,�͑�gl�V� ł���z��Bfŕ�ɩ�PwT�U~j*�6��Ȁ��ݵy4c.����
:7[]����0�'z⎰��v]79�����1�L�@�p�y�h�w����.�)�
��i���bH�(
@��"����!�i)*��(���)(������()�
@���*��������)���������(�� ��, � )"&���*$�"*�����J�J�J�(����
��i������h������)��
"��**j���(������d�����(������f�&((���*h���������$*���j��)��}���eH0�Y�m�Zޛrc�]�)�)7����@\{�ﻢ�����=W�������ѤV޶P��[7!e���G��f��}�*��=>��o�ĦW��߮�ϫ��{<��u���ψ��*U���y��֤����B&v�S/�N���V��Y����,�nS=�S��;j��+��6'�{�:��`�b=�Q�{&�Q�����*z���K�nhWC�_��ϻ��q���e9Ѿн���?:�j��<c���,�3ĕPe�"E�Kjr]D�P��ZzpQ��3ޅW�g�l���~��}^eo��=�n�K>���2� �ZK�f;ook}~�4��z��;�Z�h$l��U�}��>Nv<KΦ=n�ث�2\�|��su=���7�I6�<���ݾ#��Wp
E�@UF�!Q�߭#���Kf� �n�a�c5�<Z�l�ň���Q���#�R[���H���
���g��L�ފa.�&ӗĳ�8�{gݶ�yO��㼼����~�F��cnT���d7b:�
:�G��x����}Ό;���6����bj��\�v��k2_��B5b40W�/�C�'hFH[D�1_K[z2+]{��oS�:¼}^����� sE�E�7H����!�F�B^;o�j��]F��mJ�Ok:�U�<f`�i#�.���%��0�Di!yKe=��5�{Y��\���l���i�NZ��2��8#(�jHI���Z�'��K�x�/'u]ƆSX�� Sȍ3����/��y�p�w�R��i�s>~�=k٢�������=Q���'�#�S�x�`��D��w�d�7Q���{\Z�x�v�b����52��}�5~ڱ��~٠��E�d�p?rۋ�!<�;�gsy�*��~�U��T��>9�͌�V�L��yˍ]-��;c���p�rN,��G��\͍|/n��I�K�����xh>���*�l�D�J@w��ԙ�Y2ϑ�V7��|��~�陔�o*�����o&Xl�9�,d�I���)ò�Q��'K����?��Z��)���gW=>�+޿\wg��1q��:n�'�̨�J��_mT"��١�"}0�7F�-
�~3j�*�{�r�N=��g��u��>*��]�(賤��0�j�b����_rG�O=岎��ºކ�8���o�g�;߫��	���{��u��Ǹ佤Y,���80f� ����Yic�F�^��W��Y�XV��XT���Ijw�D=6�Tǭ���������Ellv��[]֩�7��'��s�s�[*�[V9�+����qD�=��'1����X{zq���dxތ�o gj��{������U���W�Nn���N��[a��z�V��;u)�c�L��b^j�ق��_ҏn�BD��w����u#]B�նA,���d�g���X�#[��%ݵ.3�LN���D����T���Ǻw��K�L�x��qD���7\��C3ॣo�!���ُ��>���&}�"����7���u����F��S%Rap�1�O>��GY����V����np�(Q&���Rn�ǆ{3v�v�
�-�Gϙ+4<"��Bk��=bf�Oa��}Gh��OT���<Ufo�7�/Ez9z��~UR:u�}�=>��A<��](��ai��4���U�l���.����Y+�O����^m��p����~uro�M���>Ϡ9���ːj�����k/��zB��,�ώ���ñ[+���R���ח!?]����\G�����,m���]^��mt_U(�U��ν{3^�<
#
~:��f�*|N��)�͵a⩧�0$�s)Y���m��z�=(M�,�qu��^��Y�F�g�?���χ�:���J���j�E�G�T�9�"�Ʀ�|�(�i�>�[����ہ�����ʟQ>��!`/��VMi��:�se�9D�b�����}�{_�/�^^���~+=t�qϽ�/V������<5z��2�o���!~���x��O�^k �V�-��!�k2���Υ���8�����wGs�Iy��.��)���(�����;�γ�\��%�f$W8*�7S F��$�t���WV�܍�����:]��wS���k����Wf���ֆ��W�3&���ν��3�2� ��:�x<�o�d_��{�޹c��iW\d��E�t����$��\�=�;m�Z`܏:2��۞,��v×��{%�����}8�^���v�Hq�k��#�gyϰ���������qS-φ|��Y������r��>}%���,�sf�c�����8[�ƿ�ed��P����(��.��z�HW�ԆO^���n�Y��ӊ�{�ݩi�Nc�|��d�k�@�돁o���W���.fS�7;o��:|���=�ο��<����
�FJ5�.���W����bH=r���v'�ż���?x�N����V� r�x�C&�n��_�&�ϦU��͡���-S��z�x��W+�WOQ��{��uB�M1Q��j�&��R�=^ w���*�ϲf~�*꫼'2��ϵ�Y3�`��6��{k�W�Jg�lv��w?Xxj�"�2y��zV���[B�٩Ź���_�r=�'�9�4rX����Zt]k��ާ�������g2e�JU�9TFn�6nM�x��{q�$l�kSF��)='hRl����yȷ�.�o@�޳㕒b�O:~�L���.����Yx\�"󳫬m��S�k��oi�b�n�;ە���Pa�!mA{YݦAC2�;��$�R�=ͥmN�]�8c��R�C�/�(D�W�7����Old��#ա�O�踤��ަ==g���S�{�r��X�w=���<�>����N<�ī�E���*p��D��ds�!z�����ĩ���'c���R�-�9ʘѸ��c���9�^^��uc��d���b>'3b����ʽ�ꊁ��=uz:�=�ގ��1[U�$�'���8����Y�y�7'c�Q�K���и�S�z��TWu�s���2�}�워`L�2�m�N����b8vX�q�L���{�n�g�N����k��o�>���G�[���~��`�W&:K���%����)���up�5Ӄa��/�X�kJ�kW%ӥ�!߮����Ze���H=_`H>E��T��O��C�V+��{<�3Y��rd����!��,{�U��>:����V2}%I�|eDH{��e.�}��o�E��G���n��������(\*~�}^elG�*����~�Xy�d�h#7�F��
.�W�8.�k��l��/�q��F��ak����w�v��l?RO��#=ULS�̗)sy�)�����#5�[D������A�^��k{�HO�)�Тo�^&vJ]��w�lJ\��V�J���A4ė��&�Cu4�k@`��'����[�/\�UQ	��u ������]��<E�k3��5�$5��B���\�^�+��"=O:�Ee.�͏�`��RA�>��_P�|��w���8�}�������E��*��\n7s��/%^kƘs$�Pu%�Ɠ����i�{`�yoE��[��|K&j��v�ݹ�6�L��쬖��c�dEt�&+�s�`̎v#�"�N�Q,��ݴ��ùч=u�Ү����s�����j�c[vd�	��>F�
�xd��N�2B�>��މ�>�qԕO
�cƟN���-���A�����T�}��=3q��'�{4X���RGO�T2a���0�џ����W�?_�a���zW��ʘ��o/�#Ϋ���P��ՏWNC�U���R2�Y;5�������.����)k��,�P��\tT��>8=ҙ��j�)�xO9q�����c_�;4?5�}���1�fb%���`pp�;����+�^1��%��j��S\�'�S�g���Z��O��eET�����E>U�໙��Ib� L�W�T����4�yH��K���$�O�N�d;�N5y�����{!ڸ����b�mO% X��3ŋ���=L߇��=���=S�x���H�TШ�������Y_��Y�r���C=�L�Lo��[[:�E�ٞ��t�e:<�\:����ZCف���G%V]�5�nM�7e����uYb�G���,������#�0epIjs>�w Ţ҃C������ �ŗ�g]*a�ꝝ�s�p�0G���xn{��W�P{�Y�X]�j4��24�(T��}��7}���J��>˺�K=�������0=�l��0��v���^����Q���O3�ۢ��U�����"�G0(γ�uBYЭm��Jߎ��;�΢��ڪF��߇��?Z�[�w������3Z��ﾏH�k�>b�x���mXh�+���z�9���a�F��Vr�$'��/�B�"r+��$��w�][5jdPGQ 9���}�Rѷʐ�u�l��^��\zc=��YIv��\��;�o��;n�٨D�|:���c��4.����3���v��^ƙ��K�=>�Q��,ǘ��r��8�|�X��)ۨ��rz��/\	�0_O�Υ���T�}⏘�|���k���CN��~Ws��K��>�ȊO.`��D�2[L�F��Ӳ��[x���v�G*��{������i�}��8� 9��wSp��+C�98�����P��F0�t��.�/K���Zl����ޜ�~�=&��LWmQ��U��r+���zk���.`��"�T_��	�v��_v��Ա�v�v�P7��bs΢6�� ��"�e��{yA�c�O"V�[�)��.��cC>t��W�[�l��Y@��j�0���☈�l��KU6�;Q�Ǉ��{���E����h�Ε#�?�ϼ�=3� ӓ�N��Y^*_��ޗ�y��=����<�S�f�C��?"ͻ�*/q�<�tz��5w�?z����3����ۙ��CgC�����W�w#U0
�0��S��U39zq.�{3����<�;^��X�V7���۹�(2s�yB|�Y5�Vp�m��^�ޯB��o��u���#�S���g��tn���WE�w�t�2{��<(ۍ'^:͌�~HuFz�WJ@�P:�x<����q�W�=��c��Hxj���Y29�{F�ΧLvO��_��$����tg��"Qе]�5���K+��9�^��������I�=���{��'x�$�g�Hj��}S-φE��˧4)�^�������鹀�5+ӣ�Ƴ�'an�̱ b7��~
P5 ��C>Yt�}^�)^�Fb�]�~�M紾�G����[���|{�sC��BJ>�b7��C�Ɍ'�Ny>���1�;k}D���F_��޴����6�o�u�M��btۻv*ђ�D]��� c�q�7��|�Z��5�o1R��Y����V^��El.ĩ�e��P|���:���*�]us�k!X#��f.�:���޷\D��n�q���R�Җ����i�ǁV=)3����T��P�݊.��V��ӭ����^Έ]</�p�XD��h�Z�wʏ��=�5w�����팀���9�Mע-۱4�\�8�x��;�p{���k؞,옑;���Xɭۅ��W��=�R�=^ w���7��2n�6U���5`�;��{�F�e���S����/�h�.�����<����S&I��Rw���f�#�u��2/�V̚�1�ac��Ǥ�|���[������u�r�gT���/=ôn��1�
r_�>���o�/�p��|J�0֍�O���N���3y oZ���uyޮK{`�����x<2<�ݑ�k��{�V%\o�E��yS��K�f�Ni�E<���.͕��ٓ���F����n�2W���w�?���#��C*�E�>'v�7���	jh�Y�T�Ѽ}uTz����f�ȕ�i�15Dt�R���޺�j_��佶��!�=XA��Ⱥ
4'�3�#���\TOY����y-�U�ѥ�Q�Y;�S;.a3�ٽC������X���OU����?�Z�qcK�����|�.+�������ޯ�Ί-�*.6�)4ۗ�Y4�x�u�E�~w�e�I�8����FA�M��t߁k�{�O[���A�[Z.�R�s묛*WoS��e�WI
��X�Z�KE᎖i,h����;p�{Q̓ ʌI�
� �6���=Y���뵲z�O��
��Z�����r�VG��y6�2��7}$�2���XʕHOT�\�ӗ��/3]����&�7��;mS�a�v�V�V2FIF��OQ���"ߨAȟ8�gۗǢ�RU�.�ۗQ<��:~�}^eo�Tt������Q�$��2 rm�	��z�e+�^լp�S�&��=�8�|V��]����;^G����o�����U1S��.�S�X���W4��ϾD�@�������/0GP\l�=`$�#���O�t��A��[~��`��mks�k�W?���X�\t�(Wʤ�SpzH/҅I|pgG~6�
��m_���ϻqA>��N�f�n)�6O��+��Nm�)\�ٰfG;ՑBT�59���KL�=�ǔtص#n�xZ�>#|����ͷfM�,F�,ivd����FHZ�YX�������z⚵9���{�m��j����c�L�~�<�q#~��Y�DTzRVwY���?l"̕����R��qJ}�˕xh}����U�q��x��jǫ��١��f��T����C�&A��W�/{�t"�u��(���в�J�kp󺾢:u������Q��mq�K��`6y�J��ܬw�
�x�k�I�y��ڢsF�ai��sޞ�5��}ٺJ:���,S�g^<�5o�5.��J:�粝���G])�H��m\�v��2{x���X�o;(�T$�r�ef�tﶭ%[�u�%s�p�F��Ɨ*e�2�VKlÐ3ÿd����ed6�R��:�!RB��h	rt��4��\��5E�^�v��h}F�7,4"�-�q���S�gN��}\"T���%�1"��ϣ�A.񏻮�����Fn�w�w@�+ٜ��0��4��y��^j!>�W�X(i	�]��Ü�K](�a�x_=��~J�幄���U��X���@�x����v���Tl4+���ռ-$�ЄIե̄*�mZ�F^�~/������)_�H�l�&�[ ��/#��dl̅�}vd
r*�2J�O{6��J�V��Z��3/J̙�����r�N����J���V�,�t�;�N��ާ�"��N8N��v]Z��BJ�\]�f�z�T��)-�������j�-���%�d�ݗJ��ë�hC(��l's�0V��&ۏ33�Yr��@*��K�e��E��۳о�f����q�#u_L��-=F3q��j��cpv>צR%�ƬN�+VMz���ԙp&]+Hv����Ѓ�tIjc��6A�fV��:KG�86�=�e�̏�@����C�+�KS:�m��`@��xۣs^�-NX'Cf&���h5�%�+����s����eH�Un���ü�J�+7)��
�K%�^G���_Jgi�ن���y%8��
�sSt����Ky:��rEK�͔�I.���Y�}s4Yn��ʳ�B��Ob��81ުyC����0Y-*5����PD�%t���/dh*Lű(���#A& ��l���l�6��mŷ&`ဵx\�|�����7��t�T��-��u��]����	�M�Tۭ[N�9�s�9�\����UG��2�Ch�:���)�W}S.-�h$���X���hzѫ+r��8N�to��&K�S�Ҭq�?#��A�xeY��t��b�}�h�ŉ�.+�ګ���ҹ+�=t�U�DJDs7�D���ֆ�zm����5W�A�r���`o%9[�*{���:i�˻EJ`g_q�V�b�)\*gS�e�׼��n�]{������6I�ۋ,��8:	᳐4�dʕ��H>2�d}u��ut�n����#}{���[!U˜�Fu-TcmbR#X7>0\���g�2%f�C�@���Y6#���*���"S�vE�k,jޒ���x�������X3 �|��ߙJ�}�
��r��'�v����a �����_[쵈��ۘ��ou�~���k����Z�"!�i��J&&J����I��
Jj��&�������&�*b�*"(&

*�����*�( ����bbfhi����**`��h���b�*��*X"�Jf���*���*����*&""b��H��h&/�$UMDPfUAQQ5IEQQTTTSQT�L��ASEPDQEQ5DDRED�AST�ATS�3QUAMUQTE%TLDRTT�ETUMTUETQ�E-!D�1,�3TD1$��1TTe�EM%#EEA�PKDU0QQE�MTU5TQ3A���~�bNӸ�:۵F�܎��2�VM��@i�b�'�
��� M;�4-*}��d�҉�=on^Ұ��R��w�n�w]��?�*���;������+T�lfڷ����r�_J���:&�� �󦠅eM:���g����a�z�K.��Ч&t�<����P���Շ�*��Y/|\�ć��->7��878��k�+����,��GE�΍��:t�/�'�tlt<�i`'~�_N˷�1�>�ٯOUc��7=t�
��w�;W�׬�ƭ��CĤ����ϑ]գ���{<���%EW���]�������r����}�Vqz�t��BgǕ��~�ծjj�7b�W%[��$���wt��|�e�C[��{��=�m�P�佤@�,��Z"�a���Z��ϰ��dh�JC�2�����K6�m���[��Ԗ�s΢��S-D^����4�Z�����'�H�Ԗ70 .;���q�����N��'�U�L�uV�^�xTWH���/gË��#<����s ��(�=΂�����o�ʐ�^^���p/<D�G-o'w��w����mПk��j,)��}�&�'�rb��O�\,s�������%�'��<k������ז&A!�;ܞ�w�ٙWkM�~�oo�4Z�%��S!�zz�l������.諔��&M3�	((�
-+Wa��'��X%ӳ��TR�ܹ�t���W��p�"{&�}�F���n���2SP��觩ٍ��[����9�2V3C�)[������=�&:�f���@�0��)�壼���{f���øi���۟�=>��E���p)K'�c�v�z�@_'}����QQ>�n���ڿ�n����ήM���~�������ɬvc��뚚�ֶ����]|���\}N�M����w�R��u��O�Zq�@rr��A���>*]��,��P���)��l�������_�_?�_����\��h�f�~k��0�#��U<��/<1�D�)�TO{���7�l��|vv�g��|6t;����J���O.��gI�~��:o�������K�쁑.������CW���neN�E����|�s��E��4���|�/U�A�@5��'Hʼ���>�����-��w��T鿅�Ov2YB���/����E����Ӫf�Py�������q�W�=��c�=v��dK�Cz��wS�~�"�:=K��9����.O3@�PWF_��J+ʨp�x�V1�a>��{��	�&�%v�������q����R�}��lw(���N��7)+��[W�����8u������<��j�h��u=�\3�H�uN�N�$�*��+��8k�&���F`˻�C�mn]-�>[�����V��7E)ΛP�'��`\��x~W�؃��v	;�"PRJR<+j���W��ƭ0Tr��x+U�Og�QXw�g|�\>�����8 r�aJ�7(dB˧�va5�beM�4t��«74�ݖ��ӷ���izN��z�ه���( r�� z~������J��;�V�kz��U=����ւ�T�9ͷ�����N��ثFJ5� 5�^���t��;�W,���I�O�u�)��5o����*CޟR'�=:<Jnr#]�;�2"tg�]��;��;�*q�K|�g�d6o��"g�N���j��6�E��u�6ۮ���t�#]��3,�*�!X�㛯�_����w��]aV����L�S����/�h�.�����{>�����u3�
��@�U3滺џj&O�]��}>ɓQ
a�5��c�zpz��Zt\V��ޗ�_w��F��]�^og�2i1�]�<��%��������a�;��L5ckC�����^���Q^����X�>�O��Jx;ګ{���J�Y���񟴫:�[��#_&|w�K>��U�M��k��^
��ֲaL�K��[$S��'h�h���~�9t���/�WK���h;Y�T�ͣS�i�w/653�[�ʉpG���R�fLT�c��:�Š��*��e�3��i�t�ަA��iY��C��Ll欁y6q��w��O�R�R>YgsU�Q��~����yz_���;읅��*c�v�tO�Aj��{������-�묪�S'�=J"+9+0y�?Iz�5�~sâ�ټ*���q����ĕ�j�o��]�.Q=������N����B8vX�q�L���{^��W9��c|���M�����oq��5N��w�I�������'�*ߥ����P�'w�1�qw��)9��θ�}�TQ~-�ί���Y��G�e�`�p_$�@�c�����Fk>������-�9>�g��Z�~<�����g}��ݐ]c!�%#���eD^ԙ�������N�����\��H�9��]D�N�P�Oף[M������	۰Œ�/iY\^vjM��岱��k24D�|��`��fq�����*ç�ъ}O��;M��FN(K����L��L����������騆@M����AT4n�P�����|�}��3�g�I}1V''o�r���W^�j���2K
��7���_�
���F�/�D>B���>� ��_��g��	�e��2K��^�}�������j(�E}�3�.+i���z�A��+��xf���v�Gr�w��)�R6�sZu1s�b���ɖK�Ԛ*E��>�o�U�6)�����`H��=h�Zk��;�	J�f��:jΛ1ۙ�}]�Io��Q��/���$TB�s�pfaz�*�Q.{Ƅ��5�}�f��7^�[^w.���Ol�T�ImU�N̛��40V��$��Q;Q�؉xA���\�����/ �/)ꗴ��=�l�M\f�i]��ϡ?]�X��̈́��N�炣]���K'kپ�������ѱ�,>��'Y��;�iK����8_m��g�u^G!��x��jǫ��MDtޒ�b.lNN�󫗛�k�?�0ՃnK+�N����� 5Jg�.��9������K�1�mTmo�It�|�����ū���,:���t9ɞ;2�J8v\
[�q�4;�Yu7;HџT�~л��#��Ju��V7�S�`����~#:'�U��Α��[	�򛔷~A��E�c��7�bs���g�����W2��t��v�;��Y��[SƇ�K����5�Q[^Ń��8V^���ϣ-PG�:hy��_����st��w]��8�w�Q�:I��bq��y�[���5�)�J}��r���|on뢞�.���џ=�l� {F=��1�*^��PUK����l����pD��f�����iD�Re�R��._a!�p�����g�ȡU�w�^�	wdF�=a���Oe�ɘy�F�%�$O�Y���]���O��m�_Sܜ7X��f:\"Mi\����+��u����y�U�1����meH��L���gǣI<̆"HY�H�]P�uZ�`*V�p5%��΢��bX�W�J��{�N�����.B�C�� r�����uG���Xh�+���z�4��)m�z=� mP��^s�>h�}�#J���#n=ul�$T�(��=���j��5�)Ӂ1R1�F�q՝-G1��1϶�>s;�m�bv�ݳQaL�zI�ލ�9����oo_^xm��qr�X���t[C��f6�]ng�_Yg>s>d���J�	�F\��3��@�����´S��Y��)�>���Z�c�:#�?+�ۯ������O�p7s���re�w����"Ѳ��N�ߨ�v�3n����Uto�N��v�4��{>pB���(�]������,�P����w�z�L�|}�r���.'�.h )d�YA�=^<g1j�B���|���O�����g.:|
5r|�6t;���6�>'�F��žP��D�{��ݺ�շ����a&+�O�������ٴg�g���&|?P���(��}�vG��t�ɋ��iCeM��C��*��6B)v0J�%ȇ��k���\.�����db�I�ƾ��;
.ị��(!�ky>���*�b]$U���ɇ!�^.����ĝXfH�wd,D���˪H����9Ll��l�p����2a��]ۃ�r�&���׀���<3�O�%�3؝X���z�m\Δ9��ȕ�&�o��b�{���\����"z@� ��N�"�y{<���+�(n�����[S�y��� <��������[�&��aa�����L��n�o uP�q��������e1��<6U�+�Q�9P;Tz��Twz�Է�z<��*<I�I~5�3�ї����V���F�~8�K/�DW����]q�J	��2���yϾw����h%����2����C��nbzd��_U�^]���,�b���ј����z^�ϸ?u���b.
)�@ʈ�����އ�/��_�#��WQ��J�����HS�R;����߼��V1����BJ>�b7��C���bX�~Α��[�o:͒=�s�����ђڵ��q���&�~v'M��b�%�9	���Q��3��R�}� �	D���Q�/�܈F��|����>�%�r-7^�cb�g�'E��5q�o��	c�3�*&cI��������ۅ��К�I�{ԁ������ԫ��k]���c�c�믮O�U:���.����l��2�:u��sL%�x��(L�*;�P��<,�ǽ[58b��u;�۰�_S��J���t�.�CK'	����_^`\���K�*T���`�R��Nʋ�+"ڽYK:+��.b�֝�$e�vq����� v������o�<.����}Z*���]/�����Τ�f=d�p�N�.��GYl�)�_�:��}s'aL2��KcӃ��JӢ��}~Z>�(/+V ���o*�X������ז'U�8y1NK�b'��QZ^ð�\��p�"�P��vN�����`ST��l�5�m�C����u��
g�7��zx��9����$����oJ�F���1����O�A��lQ�wᎫ����u��{�V9���Уo�z=�'+Wu)�f$�/�+�Q;��YC�YU�$�O��rVb��nK��{2��ۘ�$O��>������l^��;b���X`��N������v}��W�μ=��vt��Y��)h������Z���=�.5N��w�I�P�	��|�/�З4F�UJd�U���Uz}���S�8=�,�<��c�q�Ȃ���Ze��A�X�b�)�F�������oѳ���W��V]l���Wk]����(��,��j��*���2J4��z0Ǣn��"S�!�0P���Pd*wWf�nEE�\�;���q��iSn�jؕ2S9O��h��5�p�b̳G�Ԕbon(	��u�&�q&���L)��"[}����riAo�得�f�`�w�]v���ֵR)�.��r��!���Hy�>��Iq孁�t�GҒ�Yu�N�P�Oף>���+cʎ�q�'M�_�=j��k��՞���k3�U�'�2 %_�@��u��<�fƂ�-}b�:}�����^�8���Dr՚n��_�	ux��ݡH���D�5� 7\���0*���&3���C��%��V^W>Ǔ>h�>�����z�oƶ�,)%�L�b���F/��g�N��}a:��}^�<ƧnJe�,�\�%�F�"��d�W.zA0��V�x��c��>�V���e��z��9�>i��������%��y��al�2M(��#$-��Ƙ`z�zY��j�r�f���ף"�+M\f�%w���?]����O��'�{"�G{*A���k��%s�W.�A���K̗�p'tßN�}�ݽ^=�y~�U�rz��{f�����9�^�-1��Ng'ՙ�
�d_��v���;����#$��8�Vm�q�����{B��~�o;�1m]>j�%\>��o'$��O�Ӷ^��t;�������(��e�߾[Ӄ�{j�٪ٚ�{����BN��'�7R9]�K=�y����d�����G�T���	�h��5�V*7&����t�w�f�Y����N@2M96�aqu';E��L���\0�Gz���)"8����1�}����g��R��)C�KY͖�^�1F]��9a�{��[ѹ�kU5���9�{ MX�Ư�o�ɝ�t���Bg�����4�����^��}JU1n}}>\���UȨ8�����n�X����N��'�̱�>�m��^��,�hfN�����$����#�6j�v�Ņ��ǰ7I����m涥�oqI<k=���j�VI�#�,�S�'��������[���O�w#�D{��c�r�0<�`m�h����oۉBFI�\t���b!�Q�:��w�n�\U��ߴ真9�f.vx]���}�H=Z\F�|�cJ���	t��k�,	�7P(�w��E;��=�Z�Gt�伨g�>�3�}��%1���7f=a�Z5aL�F����C	N���23G�w�y���k�l�|�m��u�nxo�z�1����;��M��O���5�J5�&\m��mSQ��:�q��j�bSC�WO��a�}�cm.�
1��,�q��3C�)Z�48�_}T0��T�#��7n��-�qv�T�S�qE����T:\��.�"�T��w5��vu_�@�� DW� DV�j ����e DW��"����eD����� ���"����U DW�@DW_"+�_���E DW��"��@�J ��� DW��PVI��J4��(���@���y�d���<��<:��@ @PT(`��J;	U$����( GA�%@)E
  *�*�� � k	R`;�Uv2�D�iFQ���1U�e���
h�)J�vQ*�R�N ��  v�  "B�+-L�
���:�HF�)�5�,*�ұ�م ��RJ(IH�p n��&�Sl�5�:�R�g`�����ԋ�ҩ�PN  �ā�h1��;��VԴ5ѐ�݌��gn�4�Zf������j) � U K����6�h��Ƒ�ں��l�);t�`"ХdTEB�6-�]�m��i))MU #c$٩P�ɔV�EEE@�8�J��12[B-6�m�P@l�`3e�PR'�0�! 
�4�V�$�L�(�`3-�TEG��I*(�fP��%l�Y�i�͍Z�     L�RH��14�`&&�C M��0�)%F�b42@ 4�4�ɓF�� �0F`��h%IT�4 1 2h!�2hsLL�4a0LM0	�C`F&��d)���4�b=FM46C5'��>�~>_��>��y�����HH�`?�S� B@'��D��q � }RBI �q����L��	�A�ד���?�?��?��u�!�$�Hd�	 �(��C�!	 ��B ᄐ�	�C����g p	��<|~_g�܄	 ��u�f9��=��p}�wi1>�i���}�C8
�H���7���{9�g9�O���L��$��q��1�<�oԯs�V#����M0�,*�$AWcJ�ۥt�}:6�U�/�����ʛT�]�m�VW%%�{�wk���A[��GM��w����.�&s��C��(FQ�������
y��ܬ��՝z$�%��E���z�5�����
��X.��6�{Y����ܬ�^T!�b�>2�b�^���%{��n�s�	f�1eM�Qf���3	t�7w�Bq]�nD�����ܰ��wV�.�7�X�h���R S��e�iڳ�q���	]�� �Ioo>�c�v�EE�іr���9T0�m��j^�X�U���*��E�
�v�uP*�Qr�2�� �Xn��{ Z�i-ݫ%=�Jۭ�lU�TM�(Q4i��T����cz]gp}��;���f�n���S��2�ƛR���h�e.�͋?b_
	��՘����:UX"[�6c�f	q�r���fS�ͺ�D֋�u�l�1�%����lmѵ�3Q���Of"F��շ������8�K����S�����x1SPl:���C/R�`S��mk�v��=�E�b�6l��23�n˹E4�,Hd��l2ӻE��
���V����jG���,&*j��dķ	+n�U�BA���d��iQ�YT�1Xr�=�]�k
���d6�lǫS�r�q�&ȉD���f\�Y��;[W��*P��-��]�Z��Q[m,c4��,�e��մ�&��Ӥ��ye�w�����+Hff�+�ҕ[��1ja���
��fk�m�*^eC�ä��m&�{[xP���Qj����إ�m�-���S�Ҟ�[o*�d���T�4g�m�9�2���
���u�)�U@_\y�K̢N�<p���(E��`�*�A{�]G��jJh���LH���۩q�n�^&����x·�G�:`n%*��XȮ�Vh�uի2�-]��\�Ҭ]�kf�ݻ��!X��,��rQ9���d[.0]�h�h+LׄۗMIz��[��I��>3eE4����*�Wj��ynYN�Z3v�;�	�2��ȭ��ӓO���#i�ы5U����N��;�6�!�-s�Zv�P�}m]>��u���2�-\�oV�S/)�~khc̙�ѽ��E�&�b�رm��Qܻ��KU�0��̬�K1��m���֓v��WThf�U�v�^��۬C*���T��fk�*^i��ّ'��:[-v��G1b:U
M9wT�Eû�`�|�F�fS����LGt6��mmnQYݨU��t =\��j���c�!ֶ-Ŵr
���8��-U��j��eL�0�7i��u��%��:F�a$�٢��V��֫��A�qZ�.�;��kmm�J�Qm���na;�6b���aZ���۲��3����q!��z�9bβ���;[@�ݡy��-z�����Pe�k�/�T�]V�*ӳ��iJ�.��m����όeb2�L��&c�z����b���3��q�[+K	VJ:�ۣGL@�����[cѻw��1�1��K&Ϫ"ζ�Q;���n�k6Sª���K���Ɂ�e}wXi�Y�jT�n�h�v�y�41Wz��.��{�{F$������sj#�*�8C4ifA�<�Gu@�����^�l���Ø(�Z�n���%��L�!��V*3�Bc�t��U�e�J[U�5V�
Gn��uzl��73bZm�B�� �d�����ٓ)��A{iыE`Nn�����X7�u"�X�Y\2��*	[<����<(�UUL�㼫�y��]�Tƙ��e��3U;�+���p�'J���M�:���a�iJ�B���SD����H�Y���)�Z�+�&��RنH)]�F���'d��o";b�Nڷ&���U�ƓŠ �8��kjU2umB�ح`h����u���i�ECi�Dv��I\�{�ʸ�����:�l#*K.�a�i3n��LN�sp䘬$�b�oM��ZV�In�U�wMؕ��nXu��':��{�vSF����ۻ�+.l�[y_6H�Z˕E:��Q!�c/u�BJ�@�hX�����5tB���ܩœ��T��ǂ���UJE1��k%���B�K+�n3���.��f�ɛ�yZ��|���L�)�p�ὼuYp)wf��b��0�hn��^�!��*[�R/L�+/0ۼ��V	q��$�U%�ۦ ���z�"�
+I擶�9Ԩ�l��Nڼ�i�HXN�+����빊Z�����&]'�ä��ֈ��ڦʫ���뻠�j�C*Ӻf-�`���P�A�6΍KL�.�X\,�oT�"�]��N�ǵ��o�/QYm�ҟ2G>���q4�pS�ɤ�;Lҫh-��m=J��[Ҟ�q�x�(��4�3{�w,؋h�7P����U]Շ�Eʱ�R�O���׷��qZR��顳i��J>�r3t4蕗�ÃO��!uU7E�a���G(3~&�in�2l:2*��w�\�YS1�	�u�tay�F��YUt������9��a�^?��<:pvN����{P�6��).��Q
L4�Y�C(\h;�Mku�Լc,�f�r�GP$���	�wj�����I��n\֝Q�Q��3��\��W��$L8�*�c�ʸ%MшȦ��k��EZq_ץ�Ac	R�Ka�c�/#%�1��d�N��^�.�5��j�M�Ӷ�	�^�u�/�*�G��xI/���&��LjO.�+j�d8�`���5���ֽ��Ȯ�U[�W�K�G��T�t[�.��6U����e�wI�O1���Ŧ+ShЯoME3�{0MwQfV2�&���D����f����>���Тq���SPH�O����zv�j�z��Ld�{=��M0�y�<�%a��}!�(��z�Hyٌ�D�*����q8�v�Ou�5�b����3V�;.��k㔠��:�D�D�cay�����?.�3��&����W.7�	��6��OUb�p�P��W��i=��U�@��w���<�+q�1QN՝!=R(�|�V���΍�ېfd�*n�ls%Y���Nϧb�F�51�d�Ƶ&	�Q��w���Z.�oïo,���U)�E��YÔF�+��ʔ�RbU����P`�Mv�H��$��oo�G�F�;��6�%nİ�f�.f�ʹ�hOoH�(�7yz����(�j���E
�spL1��۽ڻy��S
���C��Zޢi�;P�Κ��b����Y�!�n�My�Kɛ�A]��+J4e^�1F+)q.a��s�R���AyT�h�@�&u�ih©o��@�m;��9���o��\�rs䝧ׁ�H�;����v�件�Jԩ�"*j���T��kdv�V������v.n�{ϕ���I�F��Y�����Eҧ��u���yv��yk����Q�]�\�qs����j�>�QO��O/.'��u�U<j���S�m	U�;x��6VL\����lӜ��MݱGL3>�{�,D���]�j�����i�]���"e؎�����]ԅMI���(��"��{����i�xؾ�Y�撆�V`0� ������(�-
��gv�j�r��s�y�j��o_�IT��Tl_���G:OL��u���oH�˹hșȭU%V�F��N zfҾ��B���楒��;�5]@�d���ꘔ����Ae�8HW|!Zy���{IǛ��\�<�+{�CP�yo)�.N�M�5n�:R�ulܔ��b��]쪮��Zo3\3-��vmPK	����2��XmO�JY�ذ�6��«���ೝ=�f�٘�T˪��Z�j�g �ڑ��wn�TtR�][+#���nA}wb�m��?v~��q��-��UT��nVg�6�9OP�`�QK�*�2�^�gW�M��X��źga[�:%U�f���l�=���z5v-wI��5-���;T�@e�ea���-v^�䣺$�?X��#f��+ot�yrS��9H��}]�v�g3����wA�������F�+MU��5�:��s��-�*m`���·�LխwE��xӶ&��{�����\8�{a��!�����oN
�4;��W3T�Sb��.A���V�R�.�仞KG6��ʕI�9\b镏Ha�س�����旻]ksm��55���5UIG2�+�bۨw	�qUeDg%�6_J�'t��4p\�\��]MTQ7�ҙ@�X�r���Ӟ]Z_�oڮ\�K����v�d��кm�Q�{|���Q<*���2�E��r!wI���7�[���Wt(%a�W1g���Fr�}2DHǨ�W�>�hn�*�l����ZO3:;��Ѩ�ܛ�\�ɴC�$'��M2��{s:�_�tvO&8���	aS.�[�vn�����+V2��1��!��s�n�fv�KA��8�R�m�)hj�.��D:��}��;޶�C	��U^���%���¸-�Pș5����s��]i*L����]i���xI{�e^f��r��t�Ʃ��;S�Ù�zPٰ��/h��e����"gn��E�+iO/WoGY6�U��,f�uf�V�Uu���5*	�i"�aҷ�iC:���J
J���D�[��]��ְ�D��=�b�j�5��9���М?N����E]��c�)��>��Q��H�4�KY�:G:��֮Q��&�\��
����o|�����|��Wڨ��R���x�	���K�8�'��@;�!�9�přZP\l+�NN��(���@���*J7���w���ԄϵBo��s&6���:Mّ�Ҋr:ȝY`��ޘ���D�v
=����<*^E�LFU�Zw:]nKX�JL�����[���NJ��HU�ųfdJR[�nU�.��P��˹]��R�Yb�g>7��yJ�Ԟ�*³X�/�������I���XZ�PyG�;�3�vU�5���[7���jUj���MAj'v�mu3�>���YXm����sN��+�V��l��mq6By�Q˝`��c�27%��$��$�I$�I$�I$��3u;�8v���R%'v:t9�r^3��a��=�6?��*N��Pެ���ު��zi�+O|ȳa�*m���e0\������4L��%���Er��lnQ�W��(�:�9ݵig�p�r�`�hU�f�;����{q�:���]ݛ}T�P%��{wf��Y���)�^�P��I6ݘ�4[>�V!H#��꾾�$[�D�z�P�$]wFԇh�N�u�GU�cP{��Op��M�2HT�|*T��72�A��Uj�'e�!�[f�УqU+�F?����\�f�(�_iD!e����3"n!�(�Uwu�|���J�M��٫�0�_թ�+K"zm�˗R�0@e��F��i��������sw1w��X:�u�&�cBZWLV�>L��B�@���f�/&Ө�#��1qƇ@���c��U��*�]�w�nB�{s�7Դ���@��ސ0�j��*�5��Iץ2�N2<�DC�?Y��چcvi��f*#�����?#�+�3�ѱ�ux�*x�z�q[�	�W[�H��~W�7;�1$~'�h�j0����Aqj�7LH/r�f\֍+�Wn�Ξ2=B��r���W�ԐwV���ܔ+��H�oi�tPCSP"7��ar`�]�s�����o��5:���=^��^�L���ńH���8�!!!{9����zլ�p	 ����w}�������`��}��q���6ku%��������2u�q��C+@]��I��4CTQ�b�㊷,����d�	!����Z��)�T�n�h�n>лX�5һ�tyY��x�B%c�54�&ɥ��p��YN�51�}��M[A��4��S��f��4�ؤa������j��?D��]!�V7`ŷS�1[��W;vP�������	�rއ�[ ;�����c���40���`�d[�����hWmm�h���2/(:YKe��ۥ]�z�����l̤,�g�H�\R��'Ωbܰ�+�n�y+�LtK���wN�UT�I �m�ɨ�!1yyP���<Ә7��;e�4�T��I�<�ή�� N�g/��Y�
T�q�B�)�6D�:.��e����g1��B�iw���(�FA�ȟ"�i�M:�z�k�˪����ۃ\�-ݻ�vS�$;��0U����_aJ��ݐB�������|hP[�#%����G�0L�&�Խ"���+�+=�N'�UӢޫ7�(�j�.��t�˙P)c&��e6�JB�⪎>�̨�z�]���S_Q�T��RU�U$zM�L��7(�>�/0uS'1�n%Yf��:x�)�|H���;-@�5R�*�,���N���*2N�@�xnu��������!vW^μ8�����j�.��K(ӑFp�Ӓ�����1���0�(aJ�LYb��"�U�n5��Qԙ�!պ�"���7w]�H�N�ӵ��th�����uql�MSN���ܢs%�K��3On����0F*_p՛��.��b�+�ƶ6��<}Y�R��;��UYD$���Yݯ���i�`�Lh͗�rݛ����Y���c��_;�Cע���Β�ܸ�tRWYi����+�4U0v��e.��#J`
�v/�5�!�~��Ը�@��6�42o8�d�Ǥ���\�ןf�4��c���u�S�K�����e>�&%(q,_�T��{nVQ<V˒S[յV�+����^٫��Д���R'��=�wP��!;W�2,���˂�"�?@f*r'ts�&m訅"�b,�-W(]rx��XUEw�vЬ�s�\5Ծ�tub��A��v2e:�/m�,G�����s���8U�؄̄�/^j�e�U��"�5j,g�0���Ӧf�P/2DY
�v�`-��@8��}��ae�=BN�o�]9ͩ}C/M��,�h�+U�N�ʔ��H��!�b���ba�W��:�꣈�/O�:i9���8Pޙ
̚2?�z��M�t�,WT~lC٭<F2��`��z��'O�h��]R��ثX��$]��7��rw(ˢ;VUn)�L]����M��+b��8��w+�/���@۫���	4�Q�so���E��f�G
9IXQt����(��·�۽�Z1�9ï[�PܩG��@b癁���B�ŝT�0�pΣ��T���#�w���b�7t���X�eVt�	�X��,Za*r���M�E�Ƃ���mu}UCU}UTSDWͺ�#Q�Diz�]u�Q�mjv�5K����Բg#//��Uh�[�E2>�E�,��Ya���!DJ��f�F��oO_8+�'�ғ^��;f�Z����ʍ@�(�ަC#^CWS�x]����F%�U�Q|�ӷ�YE^X�V�gA���7*�����ʪ�j�_L���%^���a��w��:�K*V�!�V_]l"��kD�wF�:4�6���0��{0��0��-�]P��ѐ�UL?���QG����d\c�x�LG���aA��9/� ��[̻Xq��iZ��R��~�;c��0p�#�-���zC�n!_��fݎ9k�o+##�R�L�����/(әt+]�Œ0R6�V`�.e�v�A",�U\w��t��I����dt>��]�ؤv�Ut�#���GqM
��Ӧ��k���oǳ66��1֯P8+�&���X4:�:�l��w6�D���?l�1GL,Xt_��UW�We��X����YjV��*�]�uee'�v[v�z��*�n}(�l4�뻯�1ҏm+��t��Ծj���
�����o�V��	��aeb�ǘ#�:�l��<E������B�tfl�MKw���*�t�"�Үn�l��_B�����rvMwo(_�b�.|9E�	Vi �l�+��W��@��u���6���YlK�U.yXgJݹd[7��%>y��p�s�
�.u Ӱ�Գh<�a��3�����J�1���R��b�w6��Q�2���$���K�jqO���wp��N���wiWUyr��c�ADI�+� �س��)�ֱ������ʧ���mkT^̡T����3q��t��wF��a�0I���/��Ż�tf]m�:��T��u�%}P�_X��։�wm�j���F�*����fh�viuа�k�^��d��W��PdU����U�3���gsWT��	�O:�fWV��"��S����jP�Z�i��ZS��8U-�^��9�U�kRƦ�����r�I��Ky�ۊ3�vtܫ��H#J ����c���$!�&�)҂�������z~�*;�]B�J6D��N�Z
�5�j^bږ�-M��(���#tP�i��B�	q�YWo���>�)�C)>s��ʴ�X7e8UuI�ױKӤn#m^�s������-���0�{����[�M�1:J��LfU8��T#	$��W0�p�cP�5�]��ƃ,��|��v�Z*˝�&F4�gC�>�� XE��9!��$��迀�����U$_�n�n=�A�~����i}�ӷi듻�D#���%sy/��L3E�-#��sSo�w�c����&���-�&:l\�Jq����e���U�T� 5�c�&��.��&.Sq��u|Q��;8l�t�%U�e�0�i�$<Ӏ'γ�����=T7�fQ��0�3�q�;�}q�]L���w��	�����Qj9�>�����mn����R]�{��	!yܻ�s/�(dU����z�~��bA~5~�5��/zt�h��fJ��ǜsV6x��>�U�]_2���:���QT���R�����c
�����ŔE1�(��E"(�p2���X�+8�C��UR",W���UUUb1T��TA�-��R��"�,DY0��Ȥfg�11>�聕_��m�T_O=�;��}�ec0=M�צjJF!U1�i��^�ބhmzx�* n��\O��\2�mEn\��v&���ٷQ!���Vzf����7�~���9�Mz-�J�=��p�Jr�Lf����y��JC�l#�ו=MgU����yh_hMF\ϊ�[���ƾ$d��v���{
A�,������ǎ�p���f�FK�}���Oz���၍\a��(3��U������N�W)���4����z���w�ful��O��ZV������P�tBӝxP��78֮���Ƌƀ��dy4{��z�1���/��db��n�'3�����^�3bZ�UN�nA��r�*�"���p�����`�=�)�e�� ��m�b{�+�5Љ�/�2�VM1���nߐ�ᕞ�y�|��R~\m�Ry�qj=�^ñ�e�^nﰦ�*����x"&�s���*��=�X�g ���[@��<L�q��R汇��Nƫk��c��x�&I%���·i*��M7�'ofy݇Ȟ���N5-���a�;��U����f�+�6)��^U���8�$���9�b�杨t�uV�ּ[�U���Ng2E����<|A9�K�v�f�7����$�����W�0��V_��4�����Ia2��"��8�<J��-V���%Q�6 �'W��b�O�t䓈�ԢtzD�ev�Z�$�=��^jd쫔!�zDf��U	���k�d�%nX���=�+�
���rMds�)��%�$�Y���8��+~`�Iy�c�ug��&Ue���V���`�pb��&/]��ԗ����� E�$}`\���*˃U�g.���	Ms\l�c���t��o����=b�Cj�l\N�{��z�ܮ������H�T�qٟcp��ǱS�b�Z���$A�*Vh}`�Vb�kd�3w�&r�v�O�f�2�R��WgC|r�l�ks97a��E=r����쒰��~�ރâ�"��z��L��usC	�ח{^�����)J΄�0��pwP'��Ď#@�N*9�"6�y)�h�W�{ˡ���;�QF-%t�n�?oQZ-/r�P�T�@	�-��<�D\�J���`��T���"r����/f��.<�=�����S�LT㍜�˄7:�J�Tc��u���}�PX�6/i�Ř�u��)Х(��ț��b����85���1GØ�c��uw��z��|c�3���I��2m{6s���8{H�5�%��a���{�thn��]6��.I"��*��p
��5�^���k��=)��h�����{Q�Ȧ|P��r���k�!SXB➞�[�nQ�Z�y{7e-f��¼���^;]C�^�v�9¯i��%=^�U� �ݳ`B��	@��y�*�Cp=���Ӝ�Ԝ�S	�[D�.;��FN.�%���s�O�3��P�3�_[J�[��[K���5=���46�%���=�g�-�0EdǙQ)�J���O#:��y��rf��~e�v���ƘxN��2�ލĚ�Dߕ�M�1�uԍ�,��HZٗ}��~�Z��y�g���+|+�T+��7�}"��D��3bg�=B�.1���UJ�~����}u/����Q}��Mw;q.�����tkv�o��F[��ۍ����w�Oӫ`���x��Ͳ�Lt��[o�$Fm����4'�9�k6�B�K��*�c��k:W �H�B��i�܌�pq��NG;���&ּ{�uәd���x
�t�b�������Xm>���	�;�x=e�jo�|�D�b�`�1��;��=�b�ꑿvz�`�&��o�)k������tg^-��2���<1��cca{�6%��n*�\[�tƗ(�2+ҝ�+�r�b^�M�KAk��n^�������7�:���x�s[��Y:M��\�;k�����|fHD��׫�"��7��&a�*���h����f1ĳ�H����F�N�P�8S=xm0ps��s�9m�Z�;gC�b�8�A�y.+.EZY9>F��n��l��W^���l�� �����24�VΕy�W�y�����_:��p�y��R�8���0	�)�_JP#��it�9VOd�y%�XQXi��øf��K)��V���tNq���V����h�c�ׇ:ㇶ����$��G�G���Y08��9�1é�Q0�_�.�}���[�[��U����e���|ԇ7pM}������X��}�t��K���9��(�g�@o��P����4���֝P�:������*}�>����Aؕ,���p^#J���e�ؘ�rs�rŮ�H�u�F���(���^(��Y�2�
�t(紗-��s�ֶ��-��v�t��+�����u6^Va�Nc��N7O�hةY��EV+8iL���1:&�H�O�o-W���c;�h�,Nb�n#��=�hH#�Z��yTbe_WP� F�m1]-
\�A�>�{Y�u�ZD��NTSv�Zp��[m�d��M��]$����Ǖ����|`�f���V����+Em�yH>˰ΦNV��� �i�#�����X�L�7�fee��&e�%^p�������&`������)ug�m�A�vQ�Ӌz��X1�U��h�̅�J���W���V�`�u�8a#�<Ws���KT�8�ۮ5��k�)ˆar\лY��%�8z��6fk�X�	R�����d'U�Z�&���g�̩�����A��+���VT<��V���q�-�OnRWnWi5�8�uS.�K����Wt�J	��U���Uةj�����4N޼ށ�L�#�9:��%v�:�4-�Ov�k����RUQuD�4�e!N!�w]yg�uB��xٚ�*��Ӥ����̃f�8x��<k����v*��I�E��`�B�KiXBTbE"�"B))��X,kI�`�$X� �Y!X
E�!�E%B�A1l�T�c���PFAg�T?��Y�cU�b��v�3{v�9S֛��s�ty�^��_����OP�uf�U��2�g|ސw�������}�_����#%�O�3���ȱ'��"��s�
>��rx��M���_ hx��j=�s�ko)U�Em��t�'Eoz�$T��Zy���FqBY�w���Zz"H�0�{��̤`Տ��.���)�P��٪L��O;����y.v��1>5��z����b�n��m�̗'��yg�LJ��Ed��G��Km7�_I}��7ߓ�w�*��W��W�׫y�y[��x�2�ºف��iMv9��	9��D�xGN�O}�x�w��2���+��
�]�zqu��R4��s�^��c�x�hѽ�F�ڷ�V�G+^����<��O��K���ǒ��m��58���Oyo���6�&G�x� ����t����+D�Y"�7�ƦmFn�܏����c��3�*B�n�oG1
m)V{\Mj.f�s����V�J��q�*����g�N�!!�<�B��9��sp�B6/�YǷ��g�Q�>+s������p1<�W?_�0a�އ�_0V^�|����k����y��ٰO���mN�u��3�'�V� �)�Γc񜯠���[�C1?D�M���wn0=f�յ�oJ�Nvfg�G��ا(n#�-\v�#!xQ�~���x�L�x9����Eֱ$r��w���ݬɝ���bT��߆EE�2�楳C-�̑PHp�d�]A��E��GID�f/H�ls먀��v���|:��I�����z�ö@�t���6�@�9d�H(N�f�'l;I��x�7�����p2�m�Br���$�n�XC)!�'�@��Xt��
v���8ֺ�>t,��t�����d�VI�j�L�i��	����2x������r2�^��5a2�d:`g�C���2`It�&��r��W箶He�hL��l�L�P�M����ǖp�����Ch�x�>8���Ρ2��Y&ٌ�C	�m d��m���i&P�!�Sl	�L&�d���<1�����?��9wsĈ�l���Z-w�m�k���e���/x�]a��	FГ�rS��S�FO���٘Hp��
�<<�e��!��0�8g��!�:�w����{�,�I��N�L0*L $�)O!y��!�M�<d8Br��Ǟs|�y�{��t�L')�'I'l!Y$�	�62�I�mL��(x�3�/�q�s�x瞶Nv�S��@���r�!Y&1�&Y&�	�i ���$�'�����\�ߚ�Hi��&�8��i�L�9ՒĐ�i4�e�(��8�y��$��Y�a�v����L�!���@4ɔMw@6Ɏ,4�8�y�x��5�}��d2�02$���0ud���:d8-�i��͒��H,�4��z�x�x�:�L&�;��
uHi�4�9I��6��4�r�;`���	�5�λ޼��6��v�w��!�I���NXt��m9�"�.,��w�r����z�Ͱ��C��x�v����2C��ov�9a�I6ɤ�BgǮN��~�gg�=������j�vv�p�Bm �ܛJ/T�.,~/����_�|$�3}{/�K�=}�	@�������~����2�(NL<d�tʄ4�Cl����$4�l$�h�ks��x<���Z�L2e 0��Bt�e�$�Xy�$2��Hv��$��'I0ʄ9s����s�!˶M� ��9d8C�����t�e v�I6�*l条�0�^��7�li!�M v����2���I�6C�	&�L��|g�ws�|ﮎ!��;I85@:d�T��6�*I;L�He��Hnɔ;d5�2u�wq�\s���8CL��8O���:I��a'�+ �'�NY&R��A��/|y�nHx�ެ�И�	�O�
�9N�CS���N5I2J��L�,������{ϝr��I��4�:͐񀳄�����sO6�q�$6��$n�K���>y�A��� XD�4�B��`x�L;Bp�:C���r�aj�0Ƀ<�ӏ;��}I��8d0�X�;d4�%a��a�@�vC���6Cl�a��Hn�g������|.9vp�g�^�鷲���� (��
u�{@��D�
���wf����kdu:�>���x'�� �Xr�:J�NR2���N�*�Ci��i��<�m�s�y����2M���ON��'i!�!�I�a&�Z@��0�����ձ#��\j~$�N�e�9��C�Wt���O)�9�}����u�w	b��%�y�N�׸��{�P���؄��<�Lhq�F�ٌ�]lx�m<��`��Pj͜�zgkR��+��ЮץWk�ĺ;yl������=0;��S�7��S���u��D��*a�����b��p����y�������:w������ӕi"���������/W���V���X�Ѣ��zb��k�5��V��맍��F#�����;�P�]�L��yԗ�n����)Y�+���*�����!����n� D;�ru� r�#0	#E;��vý�:q���E.<8��W��;�����ˎ���P�EVb4Yo��^v��=r(G��3��D�־82�����UK�n�Ý��y��������ǧZ�a[02˕�v��-r����[h�q��m} ��1�7`�LJ���s=Z���"ю0x޸)ŭ�{���_q���,�t5�}g�;uά�s�b�qX3\��v��Nx4Ս-�3��n`_�����1�b|�%ѓܕ���vF��4��-&/1�Ό�w���K'�P/y�nƢ�U���^M���-�Ϋt��Z��wm)�,ӨQ�{*��٧�I�/{����y�D�w.i�~�k6y����@Z�p_�����%��TĮ;b>� %a��p���_6�2�3�����S�0r�69��|����2o���;�I�vub��Ć�6�����_s&��l7xʹzGk�֍�����NЁ��jۣ��v��9�w�1��*�܅ħb��Q�s�*�_��7[Í�v����U�߯Ğ����U�₻�B>���\u��Ȼ�n��w2=��Gq��qw-��	���Ϟ���vpT�m`��bܻ�]̫�x��u؝��[�����	EtAX���ͮ�Ԥ���U∬��m���3 ��?�e����"��O&d���σ�˜��qN��c��S�P������Q�w鳥��Юy
΃�uW��ĉ��ປ�o�2� �}�)�{e$�@�]���amN��w^���t䦡9�_Hkj�YN�ټu�,Q�*���`���1i�jU��3W
�u:<�O�!Z�)�x~A�i%��ZM2}�?~�Ert?f�pn8Zq�W:7�n����Vh�Ք*��L���!$:]}s���s>«��,G��ᯍ�}f��q��۴9m�^b�)̥�܉��V��傄+���5
Ê�喕E�	����ھ[r}�x��:���s2]�ykX�k-O�ݗz��ŕ�%�)�3Z�dr\˛ȉ)r.��8���%��s:>Y�,�zw�{����]��mr��I���6n�k9\�pjY��WI̦h�����J�ո �w}K���͗.��G��8㇎}'�y<���-�C
�0�V
���C+U��*
b�`�� �a\ ��B��Ѥ�Ke�C	1���"b�(#"֪A`���0�I�V(a�HaKj�*��8d0�aYFQ��+0�"����DDb1@Pm
b¡"H$�!��:��U���j�ff��jj�9�Fl�Z��s�ګ�꡸�~����0V��V�&��c���߱�����X�#�]e]�ގ�n�s����ؘ�Tkh�+��	~c�Տ	�q�;"ؽ��;'ܴA-5�e�<�x^��4fSSh�K����l�'�k״7(�?`TAϩk�a���N��o���n.�7�b�Ky�T����޵ݡ���fr����x_�7*�(7�>��z*���ʹ��%~j�R��4�nm���'��G�=�E����{���ږZ�R��+(�����
�j?t�;���\��D��}S�99{�R�t~Y#�T!m���O��u��5�w�W�:�u邷gsv�J��P��\9у�>�mB��ȷz�nn�/���H�*��੄�u�E�x �
�n`vS�P*2��Ʌ�6Ƒ��}�,n/	�V���CP�0}O�e�i�vx��|�S�K6�ʑ��a�(�$?ʯ�着��v��:����@ϧH�/6����p�ةi��U�LQ۸�Y��P�V"B``�T�;P��7�5=�Q���p9�0`�b1�KPW�@3�[:���Ǽ�ws�9�.���q,�zrq��Nu\�h������z���WwT1�C���+[�\il�L�ȓ4�d�����/���ʢ0:��Z��e���V�C=��soy��P(r�N���s��JBK��ِ�+��l¹��}����Pkuѱ�z����ϝ��(q�]�PӺ��呷z􃋕�.}���iGV����c���Z��q#{=}�.������2�y$�Hq�X;\� mZ�W�!3l���g�A�W[HQR1�|/	��c�u3�wo2��A�+&�yI��{-\���^�o����>��C���[�"n�:x��U��ۦ*�o��PeG&�ڮp��v+����wG����h���}�}_}��I%��GՓ�������W�G.��oP5��^T���4���;zv&�_n
I�U0{�{�l\�2�����uPY�������s��sE#|�"�H��w��ZJ6fk�J��|w0�'2̽�Z�u��OhN +���ݢ�����%���ëby�v�5�Ǥ���Q�`��/�����7r��`�v�f���4��@�quM�V#��v�t�Vh$蕽	�I_����H[��Ƶ��o["��H����)u�QcB9P$��.�)�(�����8y��"b�1���.[��ݍEQ�Q�����Q�y�caa\ �+h��nƖ���lwQ]��W�����	6���Y���Դd�/(u�V�V�b(���nJ�aj�_*��)�](ma�.T�f�[vM
�bw[�7$5��-�rn�5������w���Lj�Tӕ�I�k��������{co�g�������K���dh�� k��-�P�<X�ӝ�@B���e5�d��K/{Y��P<]D=���S��Ǻs%�����l�KY�R�#^�&YN��fۊD�A��b��=��BT��>:qKl>1�v���Y�S�b���SvQ�f_z�zC����.�EO@�Or��+s~-�n�ļ��.��$����r��\$[��6V�7gݕ�Y'��U�odS�5F�r_z#������&)ѾƉ�K�k>�S��Q�æw�g���2�o)9�o2�C� P���E��H�u��Y�-�Sq ���
���0����[���v�k�S(]N�Xӄ����v�V�E@�r��ZN�&R�'m�.�F��|�j��^�U���Y�Na��m���O��q�8�Y2�bm��j���9r�쐬/�B
��]J��2uo�gH��M���-�	��Y�{���7������W���5ܝm[��~R�O��\�O�xR��/<�'���݇HU�+��:�����-[����)�~��[s|��\iS�-�!�Pz6[��n�g=�N<7����/�I���sW<�V�iWf,�s��vs�q��2�*籼�VT4��>��Z��v×�JO.rU�x�|>�}��*g�ʕ>���)Y̭�`IJ��qj#���{ރ[Ï�n��/~��U�93�"~�]�ی3�tM�U}ُK�[�"ç���g2O�;�w4�}�W��6w�݇'=6�(��zH��g5�,�e'����7)�^nZ}�����
 ���ޠ2{6g��#����N�P�m,n��g����7E��7_y��c���8��]���[��
ď`���h�N����y���\���������w=$��2��|m	��޳F�y�9N��6�W[�>�s�d:��W%*y ہb	��U�h%t�%X�"�y�Å�i���|\L�B���Hd��[�f8x;�K㙊)O2rWQ)��ө�.���d&�>)$^�^ތ��$.�櫨���;�*�M�{��m��Z���UF�ݚp>����ʨ5��-Q�a9��r.�����;��N��U��Lk��� f��cL�+����sn؏�{R�2g"��\�i�����S�\#5�5ͤ"tx���f��+l1�*�F_�ʪ���Q5wO�py�sw��R�I,*i�%�ʇ�f�ٮ�N�����V�0lf�����c"nÃ�V7�%F��ꥹ�5\ZeA��l��y[�6�sz���&���o6����1F���}Y��/wnT���[r`=S)�춪ễB�Sy���OI3��f��l�Ÿ.6:w8�e𪄉z3�h��jaǑ�\��lr�].RF܊H���7����ȓ�,H&��³,�����T�$2H�9�"�h�]���w��UT����M����U��+��H,�V(B�"�T�V�qJ���PiA`-J�5��ɆT0�Y���$Z�l�(���E-�J�(,P�0�-���B�Ke���XT-l�k����$��\[S1H(�m��\8b��j�S
����eV�DC�ū
��(�ōp%�0¢��*,,���E"���B�J��6ѕ��U�EF�h��qkm���aP�ieTҶV�J����x��=��Ƹ��Z��x��;��}�J�!+�2/��U}Uh���?���R���=�,iQ}7ą�i��t�ĥ�m�ٹB=�hժ�]�V"]���a^�����@d���T1�{�Kr�}Ҵzƌ�Bč��S��l�[�X���2���Y"���X��.���b�S�YFT�y�WQ��� ��B�^�n�wq�ck�<`p=2b�N��P*[��AR�lg
�_���ݕ��e�wMެ{2��"���<�JA	9�z��G�70�kO�̜'"�p}kD��[@�	k�KA�'o9�Rr�wQ��T���2Y9����k����l�u�+./Ք��b�u��y�:A�r;�mV��t�#%D�̒��J1^/o���16��~��<��oG��-�v{9�����=/����_E7��/Z=�B��)q�����$�D4o�x��N�s'�VZ���]�Mk*]��:�+�]���������Rc�?��_�����\Ji���^m�}�B���׹�pq�9���.zI��p�^H���u+h�@+%8N�+�6g!� U�L�)�]��k��/���j��z��T�xT>�7���v$��+�Z*OêI��fʏټ�w��	�Ti��U�Ǽ���b����kv���R�;�+��a��2��g�������{gUr@�TF�m�y[��Hs,��L�*=!4ކ�ﾯ���b^����=����}G�]9�4��e�g_<w�pQFY���zP���o�{���}��`=�Ypy��}+�k�ΐ%��\�w�{~�==��bR'ӍEf���V���'��k�4�l��9<C���D,�"�ͱ];N�ɭ9C� �WKa����g��d�� �G�z��U؊�~��U�}���H����i��s��'>�HLA�eM� މ<���
9Z��Њ����Ά)�_��GTP�V���	�^S5�B9��6��"i�V�)���+G���_�����Gy���t;yM*r�3A�|j����o�؂�e�%�sL����.wO;t�N�}l^$D��!<��W!@�-n7�����<G�hS������r�<k}��ǱW/����Em\eӘ�#j���\�g�*Z����Z �~�D�1J���V�{3<{�;��z�k�N���HBO��K˲�d3��w�D0���c�,_LAb�k��Q����e��7t��]�����ξ�R�bڗ.�<�K��.>�t�l��m�Q �up���{�����50�����tn���(Q"ʬ�)e~�0�)ٴ,�Z�$<����d��v�w��wP�=h3�C��㤛7HC|���g��P΍�,�Fj��a�)�Y�xw�r��������+�X���p�D�ҧV�-���t����y�ˏ�v/����%��q�Ӆr��Z9��w��x
wp)�q��k=�ת��驼SoIު�e4��������s�����w���ZS�x���:���F��^u�|:~�_Z�@O!Qx�<��T�L��.1�&�D����}�U����%w�Ӎޛ ��fɖ����-�\���O�:�����^ons�~T���1�^�ꉘUw��Ya1��*�d{�f�yq�COċ>/�ާZ�'A�r�j���s?,B����fȢ΂"צ��#�Z@�6�_R������i"�H��5��x�A���������QB�?M_n����,����ʈS�3詅>�/=��+H(}*g6��*�\��UV��7��pr¦��Y�קk�B��gn��4���;�^;�]�'k��=�)H묯
P;�,�S���3D�
���.�qf��!%C<`�݅��l���:A�]����]�n]��IV��90y$�ozM'n�הͱ��uzq���!��h�&�Vz��ڼ~�/��j�&C#�{�:u���p���8u}����(���E��ɻ���%�X���C���h���P~��P�E���)��w�S�u�V�����_[��h��~��!�"#���<���<���f�wN�-�U2�}t����+���[b���Q�U�Fr
��Ik��������ڻ�hY��E�Q�.�O���d�ο=���Cڸ�x���*Є���)�93(���ЅΣ����嘴c�ͽ'X.Q4KmV�-��v�fѦ,��D&�p���������7򃵥�Xp�����p�ף�)P����C� ��(�B�p��8| �Ǯ��2e�&������w�E��C�iÇΕu��2����D8~۫�.PUG#����x�뮱��MSL�l�9��=�:��I���9}@�;zw�m�	�;�w�<mo{�|��3Gx;�W��.�SJ�.3{��ﾞ�����YM���`��:��V���!t*��5'�l�҈E�BW6E�v19�6
���u�ҳu*�XB���^;J���-6�ɔ�=y�_jׇ�����;�=w8����ncv�[1<3�Kvmǐy8�������%��}_��9���ߌa|���}^n��d1���wT���~�V�t���r�� N�a��t]�We�o�6h��c��q�Zt�~؅��/���z��e����z*Y�YB�
�[0f$�;���A�1�N���T��9������<@x� 3�G꾃��$x��w��H
�P��:gx{]v�"ϋ�jA�P���>c�3ǌZ�����w��p4~6��{KH��!Ah��)_OY�E��"��\�K���O(;ӧ�.󖺜DJ�~����Z�	4>��u����,צ{Mi�E:�_^1����vI���f�A�1Շ��J�ozB_;�c� 5:����Qn��DE�4Ҹ������/e��F ��gJ������a��iCn z����2GnM�	g�-keS��Ϧ Oa��gj�0�rrk��Y�&e9n���bܘm�������C������,N���,7�(L��qhq8łწ�b&0��[��2$�gGn�P�y&;���Y�Y�b	��巴R�}��N�n�Ve��U�����ap����GpB�[\�u�)�Z�J�n���<��4S��� ���;Nb��i�Etg9� �.ΰ�[ZrcV�[�v�*��N�_&X�,*��m˻���ub��W�Kz�C%!�I���ᵜ�E)�SX�׎�v�Q��%M,x�F>�\V��UO=���K�s�x�F�gWa�����Ì���7 �mJX���E�����2�9,��.<ai�:��kw%�2���ue�	iӰ7��Y���;�*]1f.�7#nG$Ml�9˜�\����Nv�)�_���o'F���G�uOF���UN��n���Qĝ���Kv��c�8�S�<��,[h����P�V�Qm�0"�a-J�UYmEjZ�"�P�T���mX�eՒŉY\R��6�(֢�1YF�"(6���E"EQ�E�iF�+ZE��kQ*U`�Q*T�*�1X���UUR�Ţ�&�kX�5,�+PXE�"T-�#XV�F,TAB���"����XR�*�5�b*��dQ$FA�)V(�)Z�,U�0DDQ
�UF(*�jJ�iDU��

�5�(+�R�1C	X�[hT��F�X��*��*(�*��2VJ�AKj�e�U�U#j���(�Q#RV�ŕ��*�XEQKm�eH�QH�����@UJʈ"�b��`����h�X�KaeJ$b)J�*E��
�**G����~�s9#��/R픱ۛM2˔���$ڪ�F�/���\.�Կ!P
W}]���KQ��)�:{Vʟ\���$���x�x�O�(�[�]>�L�F��ֆ�@&K�c^4GV=����+������.,�_0��B/���^����%�="nK�jg!e�LwW���>\�C�`�s�"�'��.C���W�Ӏ�@���;��>J�և��0�1;lMC��g���ܪ��H�x��1x�Zz!��\@�:�����e:�ݯ�����D9�F��ؾ���������6>���%�,�?G5A�~$0����pw��(ZU �j�eվW�5�EM�;����#�@�n$��k����$���3nW=�RR���T�}����秢��
4b_aG�`�����������_m,(�㧹��)��o^d�z��צ�����FN
]3݃��&��0�l�$w-<Q��ؽʞ����#M��x��g�S0��:2r\.G��>�t�����F��͟��9=��ҷ��t��t�P�
~ʏ �#\7�>��P`��+���B�����ߗ?8�!�D��|k�Ǌ@��shiG�|x�lq��<C6I�[t"�O!P�1�i��ǖ�F�dk-9����3Z���k��v�kZ\Iv��h��w(k����ݙW����Q�� ���f�Lx��^w���iˍb����Bݾ"�i;t��v�K"ȇu(ߗƔ ���VXy
�z>s�=�Ċ�D<��t��bk�!ľ`���E�d��4p����{)ۺo>3��A��>7wW�R��0+��~��{ی�<�yGV�xf���M'	֮%�����<�ro��U���ҏb��F#��N1N�d#������ۤLBE懃_a�"h��;����J��
fPw
|��aJ�k�1��(W_���u��"�
v�pV�|��������U�hCz�P����RL8��X�e��&N1��T�ْg���\�2��6�|��������J�������l>Z_k���M�b'N^��u}�a�!�lNTБ|�`O1|�Q�^鶢'�"�3�!\U�r&�VK�R�c���X���^0�V��~$O?��t���4Jv���@^h��F�]�޽�����C�Q�a�𮝓< ߃�=^8�X���]����c���{?���2A�ݸSQ��n-�Y����B'䚋6~��^=B�A���&�����mi�����uR
L�,ۿ���W����>�9B\oO�_�>-#�l��%gkwk��Z���-m_t��Q׻�g:)T$�nWm������������1kK�0��j�C�������y�5���.}S�tn��3`L\詑����͟�x��A�����<t45�:^����j�N�T~�TD_/�r�����w����o��t�~bБC�x��a:��x��e���1a����T�]��Z/�$"�<�j��H�$<C <F5��]y�+��Z��N�nޙ�3x����f�w�&-��>��Z'Z�����g�+͗���l
�Cpko����s�MZ;�}� ��]�6�vw{ϵѡ��W�cU��+�M�ݙQf�/�`;�m�S�)	��g\�ʫ�L���{~?
(ܷt+�a�a�[¹ы������2(�0�Zj��Јh4x�T����V��5��}v�Ed!��XI~��e5;{���M���(�l�-Y`��'�rP&3�U��R��e�go�2�管���1Otތr���l?y���S�9i�@Xj뛪޾R�ρB�C�礑ma���ykA<-׻9�+۰�.��B�)f�������#��<�z�M'/)��x�yŌ�N���ݬ���ʆ�[~�<��E�$?�
�,�l��֣ʛ�4�K}�.�{�f"P7��GY^�Ʈb<v�\YEز�S��j��RE��r2�=��N�?U��=*[��¶ͫun�1S*���P��*%�M�"��Iڣd@��Br�^2B?^ �\o�`�a־>ǆ�3D?(p�/�y�8Gy�Z�ٸf˳ztyQDY�f��y}���)�$�y:ҷ�y0�-�?qG��Fq�|r�.D�U����Ru9\F�rg�p�'(A�a��(Ľ�~�'��hC�C��D8��a`�����8�F���)|�ן�k�㦳Xq3�aq M��u�|H�Dk�N��G=he!��=�މ��y� ���!-a�g-6E���h�v���n��37f�=�8�x��`�f
l��1������������Gk��r\����ܚ��������WZ��y|M+��8Mꬦ̦��X.N�̃�㦅�|G��#�Nn&T�̱0��ɼԚ�fb�Ap�R��O�|�d��Y�V��I������{3��k7��^��v��tR�c����o^��/.��;�u��R�yM$�,g]�>㜀f�+Wj�@�����5~���I��,����B? ��ʚ/��;�T�\���"~��!��MF�;��L9��ј�L���
���ˈp�Ϊ���雱��G�͚�ո�'g�{���&��SVa����Uo�R���scv����;�{�Eʤ�i��$�	�% ���h��47\dL�}�Y�^0��_e�>5�zkPg�B6:�s�T�3�u�����پ"�xV��;��"�?a�Xy���SW�]q7�'h���7�Q|h���`S����Ű���L)���f.H���5"U��
��n�ʡfsk�>�(��*�
WJ�Qq��Ͻ�st"�b�l�<|D:x�4��z��{;=wބ��n����&�����Y�{o0�,��
fJ�T�U�0L��(�(w~y8���)��*\�TT����US�x�\�: a?z3�Pn:�n���+�����ǮZj�����G~�1N�~�}�����<8�mʚ2Kt>�Ϩj{�}d�v�sv�򻸴�����p��3���=���}�n/-�<�8寈d_Y���.��;�Zf�95��/��v���g����������j�~b��1��r����!�֜��"���q,"�_.,�&-���=w��蔒�Y���ȄC���k_�)��˴�oD\�/����x�e�.�(�a���}+aw��{�r���Gf�6A"�7���=׮5]^���a�kOTzv/��
0�_w��m�:�c��d?>�L�����q|�O5��OX�@���	 �ֳ�m���#&��$`ʮ�Av[�GJfȢb+@�W�ʃ��7�7�\5v��]3�%]�"{�c���-#�&�c]]Ϋ��,�����B��qT���<�wX�[G�P�}T��u����Se�᪸9����qo=��n���TT��l}v�Of�v�V�WVF)Q�g!Z�����>���N�P�=��K�1NQEE2f�L�V�0�9I*�:���U.8#���*���3YG7�&��CB�yMn�A#[ӯL�E�ǰ[�B6�zt���qq��[�E�J�A�E�S2��0�Sk�l=�)[����l����יB��@��I���ᢆw	�Ǧ�N�w�uJ;3~7�u�ڨ>>��a�Z�Ds��}�R��������i�K�m�p���c����>Ed��[kQ��$/-�U����R�.�t8�Mu�sL�m��OF�&�t^`\��V(�hh0J�[�	�����ܨ�T1m�_Ӑ[*�>�o�f��V/]��97Cn��Q����!�z\I��r9"h�c����Lt��{x�+uI;u���3uq<ٓ�%�"I<y��9*5AUQn�����gQ�t�y�4�)�*(*-��V�EE�J0R(�ֶ ��Ac(�`�A�1V"	+(��FF��m(�Ҭ�QAQ"ԬTe�D�QdD1�Ql�E�C�k"��Ȣ�jT�UD`�Vj���(�X֋R���B�ADUm�����*�-�UdPS	X��ył���0�b��U��QV[DQ�jh�X�j�H�bYib�Z�X�!QqJ%�m��a��g~�k|_�N��[8,5�h��9VH���?g���٧O����9uդ�Ma?W����ۉ)���(_]�_�t���Z�٠��KϕgN�t�����r
������W�}t�A=�Czbmu�%�Hx���"��H�1j�8d7Uuu=0��$��Q���p#O�K
쏮�m��ƾ\�*8AB�&���&�>m����ތqÇ���E��Y��u><��|쪛;F�:xr���\�ն'��Hx�B�����s�'�OM(�C�C�>9�F�ʝ^n�e	�x�ˍb���'8�������"�#̇�[�7�qb���n0ǵ֙svC��*"����cf9OZ�'I��Q�Z�ɷ_�Wz�W�!�ByD8~�(ܻ�άU~����b��*s�ӓ �-���Pf6L,���4�!eT*Q/�8p���C�fMC���5�x����K�q�Zr�Ma��|�����C���C���a�*c�]W�ue�4�Ó�
���C�q�7���i�؝Sx]���z�|����)!�B�sC_ab�	#��U��"α¨_����Xw^�p�w4}*�Q}[��m�}�����1�{�wJ��]H�ؖ�_ՄUK�$T�q��l��J���Y@��'u;i^c�Z&�%t<��V�Ґ2vK.���K�J���ܷ�lr^�z��FK���Uá��͓��ȴ��?/�*��B����veM磇s^�~�g
�P�~=a;~2��`���j�_TQ0y\�[�QSc����T)ٱu;�_]"�/xUw�a]�sپ�ތ�#�ޱ۷o/{�%9�}kNj=���������湯��a�!�h��9a�B��S��3ڂ��z¹��C����'��윑^w�0�=��$Yӟhy�t���Yoo}����"R�&�/���r�#�Y�u�*�=b��M�,��1~�WJ��:��)�钆�KD���2��S��mge��%�\�?��C^Y.z�Ž�w�{,�Z�g�F^�s���UT���)=HYq!~����x�7V��;E������>�P�{xî�b�B���n���]�C�D}�p�؂��yW��=Xp��S��^YR�[��ݩ��wp��j��I۪�1�T���5$Y�Õ<z�����#r�yiR���<a���6Ww�?v����,�}��v���j��+Zt��;����̪�	��AYf��?W��of�:tR�H��-�e�^,�1ZC��?]��o��DQx��yZ�׼)զks�
$W�t}p�p��K��c�hɣ9~5�{�/,ǶaY^�R+���A�*\�*y�%?DDD{�F��l�>�߱O��"�� �Yч��8�k*���W�)�n��Hy��Pd��� ���/�����dA$(���9KR���i�m )z/y���#�]���<�jÑ}԰���L�Cn,=�z�Y�G_ʮ����k���ßq�y&Ȥ�..c�ϲfr}b�X��l��fa��lI�S�� �*�T3*z�ȟ"m��Lt�Ã];"Yi�m��3�Sy�.]�G}�޷2��S��}q��z)OL(���6�6�ˉ�i�1���Q��T�wK��	ֺ{����p�LZ6�m�'W� kԬ@�w6����ɏU���/�	�`�AY�8w�BQ������ތ�x犯C���$؜syQ���h�����l�P�OI�L��R�N`��^"�̼�"����$ÄsV@&�Q� ����q��޼<}�s�Ü����
(�'� ���M�*/��{P�@C��a�X������6FR�*��V��:����2�򞮙[���E�X�Е>9'(ɕ0&�ާ��lX�=TSL���$��x�,=h/L���ݣ��Tc�Q���_�^���Σ��.�1�b�͛�e˦õ���Hz����'�3o66���C_X9�с��[j�g�Xʂ�m��e�����z�:�=}�
@���?}U�T��z����t,���rֆ|��X�R2k�ڪ��e�!�{q%�)�s�J�}++ݪ�&�<c`��T6�*���t�fOM`ۜ�f��I��t�!^�0���N�rs�5o�����'O�ŧ)Y��A|��M|�ޮ�x��CE���^D��* ��*Ϟ�ߑNn��)[��U�n��C壐@������+vYDz���g$\@q�V@'�˱{'�P�VU�4۷k���>d���A�'M��(����|=�������;>f��xY��*�m]u�:��V�n�9��}�/N��t��櫄���72�oInÛ9%=���y;/C����Nq��4�wL�ۧ�`á�M�%�o>�M�⚇A<`Y1�`�,���wr=ƓL�!��}S����Pj�|r�#�v����nV�hy�<is�QY��Z�r7^�}�l��rC1�V��8k��gO�Ck�U��<Y���F��`A��1��g�J$��Wnz������0�=k�"DO��^[[��-!�G�#jç��C�}�l�wM �ۥr	u�H[+��� 琙Ӳ�>"���ťZ�<x=>�֦�)<0��Y��Vdt4�#6�{C*i'���IM�̇sRǚJ�ԩ���PpI��eʲI��N*�&p����De�5��X�Ghy�x�澲7)x�{�{�",�T������A���b��G�ݳ4k����/��1)�B����J�ґ����3P�i��(�"�����ӫ*��n�����$�プ�h}���l��sCU:o�>$֯��ǁEfȳ$�7�3_E���Cƫ�c����_[B��׽�۝�#;�R���ա^aZ��Я��ۇ�J�˶}��Μ0����\��A5�g]d���սL28��L?2-Xa���\3��{�d��c�N�w��px6oX��)�Ǫ0�;5�68�b�V6�83�j��`zӔ��Α�;n�(f+Ww[�b��N	u.�
���+%���x����.�`w���T������d��-�y\?2���Nb|L��7�
&�� ��Q���&&$��W!d�	U�q�]���_�m�č?_ ���r�
7HV�8C�	���y�kǅ��O�e�_�Vj��ٮ���w���͐�x��>?#m1���h�Q���3s¶L�P��kB���"�?	�6P����.VF�q4��"�����6Q�wtD����q����t��55'�"��E��j�D{��]��)��PQ|��X�V�lWt�>u�֧n(��c�mf󆴙͂�	O1nۦ��
{�,���`�H����K��qiܹ��|��q��XYFL���݉��)h,.u�s%J{dq��ݙZ��lb;m�a��L�[N8n�>�Kiu7e�u}r�{nfRŦ`m�F�6xdyCU`��Z�.��&��m<e�-��Ѓ���Ň�Mr�8�t�;e��l*���nb���q��8gYˮN�cl��+P�io%+��Ρ�����an���k6�����x��LLN�BuMW�y��wfH�\���^[wF�|�&S�r�(��|1����f��̥�	��ճ.�G{\���Y7Bήy|�rlB�d����k6�i�|�1�6k��3L�X(<��wU7a�Uk�Ɔ�L˗�Ħ�ݻ�O��5 rs��Ds!�娶T"y��(U�6-/-�X�ޫ̀�\S���wV��U�ׁ�zr����7TJjM�9�햀}�pٍ�w���	�:��w#.&�i�$�=\k��o����a��6ۑ�:���s��%��7fn�2D�#sgt�5|��{y�	�Ύ��'N�z���I!	$�b.(Q��V�-(�� �Ef"��Jb¥-�YkV��VZU+DT�J+Qg\P0�R,R6����,�"�@1i�(�B�H��$"�8J�#$Y8iYY�����7GX�75�:�qucr\��,���xl�WY�����dqDUT�^�4p���,�n�7�Cj�����D%�x�-#Ηk���P��./�Gj���F�0�$�2�*�ܑ���C�~b�՛Pe�黴�9{z���:·5q�q�PU15���**|f4מ=��ö�b�2q;�z�f��s�Naʔ������`�=�Ђh f.��8��/� }�B�����s<��O�b��m����y*	l�o�UE���g��zL쉊����esA�W��bji�Jc��[�+׌����0B*!��j��ڞ���t+X��FqC�_v�H�ۨW;�#��j�F��k�k���V�2q��M�IR:�������w4m�(ګ��z��%�+�y�����=�}�.�g�&9�QǵY����l��	�G�Z����bT�;FVA�JRa�G��"`~_
��.��~��Y�r�WF�C���f�d*�1�a�DqCV4�S�0���u Pm)���F�%���������{p���u H���9X�!���3��u~�C;�Fӆ.xa���/�5�+�%t��F�W$1����.挷�˹�I��m��;����6S�O��jy7uR]v��B��f�����U����S�ع�V�u	��,�����& W���G/[�1�F���v���f�U�P����kV(I��e����~Tţ���W:sX5�2f��{�֦�ü;��}Ή�E۵:"�_*�k4��"�2뱁���gvn&I��J�+�{�f���5�����g� �{���{u�J�%�S*�6)7��F���t	���T�'3��{�-�� c�{\#V#�|�Gg<��|�u��n3�yZ�O.f���NX���b)����ùO��M��)#9Cqv�v�F��ۿ3Wsy+��a��7fw.
h�m�xK��b~) ��"7�S�b�P���%������.�+�|ޫ��g����8�)ܻ�ϯ���^y������3��F��n�&��g&=C�L5^딮�g��B�p�%o����]>���F�Y���p���!u��yˬ���l�2ͳ��^S�ӚDY�룲w��!�����時��%�^�铛��1I|�3{�~pR�u���"v�4�'���z��a�8���Mu�i���c&)�&+׭���i+���;QW�a�sGA��[MRy���\x"�nuDk	�OD�F|��y[���c�< !|;���^uB<�7��4�ʼ����c��t��
�- ΃4ǘ�n��L�+�Q2���"�5�Q56DK�in[+c�Lv���v̡Jq�E�.7P�Y3m���e�Y�.���q��L �\U8�K��A���I��$��b=��U����E�du9��}Чי4ӤM�ug��T�Z��׻�,��{�ȹ�����ܸ�Nk�ʡE�')����#:�mnAow���c���y�e]�%_��!��-	no4�cR5Y��H��z"k�w��wmjsc* �Kݺ�7ʣ��m�1@��@CΌ��®*n�3sq���=U��<V1^>q˪� am�x|���d�&�:�����:�"��W�(�$�/WW^�so:�!�;V8X�kVp2=fjY�#�s��7�<�ؼ�Փ��|6���c#�U��l�Gl:�B)�z2�Pi./`�K��kr@W���OQ[���ɥ����:ƨx�k7c<s��۴Vpac|MG��|U�o�����i:_6�t�v�[���c�stN���Syspq��K.�1�λI�x�4|<�z.8�i�!�i��]N��I�Ƌ�B:凎;�*���i�Τ�dt����+L��e]Խ�2�!#j�͍�k�\
����a��s���T����V��D;n���w"�7��ۭ/�@��zf|l����|���I"_�(��(��.UM[�^k����m
h*c�dB�뉰{��m.� �aj5�\�i��se�cɶ��ܥ<Z�?x}�*��L��q�p»����X�X�>��hU��<�BX�I�Ψ����!�ҡ޼҆Lr���<JtลE�1��7o�U�[���77;�؍�p�]s޽�Vz2
�5�ڄ�fY<S<���2�p��Kr���������@�6.v�����H�KPf$�4��Wk9Ka��l^��]~oe�X�,�Z�kD0f?3س}KN͒�پ�|j��A���&�k�-��d�ҾW㷤�G���o���M�70��Б�;ԥ�L�@�e�wb7�3���gt���ky��KSo�6�������hTaG��p׷C���:��E�~��P��T�A;�n��lָ��1A�g�`E��nmc��"��+�f�W��
�f��sȃ��k�U���D��N��~cӺk�{1���r%�ʣO^�{wO6����S�4`��n����=8�\����S�<���<w��U�w��O����ৎc�KFTo)d.N4	Gt��+u��ݙ����WƬ6��K�R:#N\����g��]��h���p�������ip����V���Y�ܮ��������N�ڝCZXҾ��̨#U�C�v�����ڳZ�M�i�*�W�T���ԑ
V檕�3:��:x�*�e��_�
�]:;Zo��G������o���9�Gq�oge�y,�|�V9���Wf5K��v�e<�K�'|5�w���-�ilPnG|�\�/�z�un�]2nRg�Y�f�S
�Gb�⦵K��.�2�k��;/�x�r�E0�A��ki��v�*mjeR�������sR�N|�,θ��|W ����X��^3ݰa�W��V�f�ht��2rZee�S��wz��3�[�M1QKY�(�Ⱥ�o&U[��c�U���顇K��	�;;2�Z�w��o�5�ls��v�;k]X��2.���-����H�}���Z�v��r'��K�{�@/(8�+w^�����;v��Vݬ8�#St�5����l=i�݀�<8��G��9�$�,͖͝�;�W\��(���7�g�����,�J|'����w��N��$��d����7��3�8�/W:�y�ʤF�P�+C ,#��6J�E��0Ŋ(��kP��*,����
��Y.)
�`X�������J�@����f���I �7�t��#�]���T��+�ґP4�h���7�,鷰�^Es�z�(\Fh���C[�qkE�����A:ed˵RR8��K�]�{�1>�]���ז��>vʴr�e"�+E��%�8�B�tj�پ�	�,v�(�F�W�>���\����ST{�޺v�4%=��}��T��2�S��V��
�%��=���9է	��8���w�껷�1�'_e�� ��z:顱6T�L�Z�q���+;��wo��NT��RV����=u����+���(�~���= ���@����)�72���Wg{����]f\����֕5 �k�=*�c1�;U	���[8���c��*�gOV�d7NX�B-����)o�:u}��=�_�o���u�N��~'Ǡ,j��7�0*��2�w���v �̓�m�-�����Z�G3�ʟM�����2�bH4�K�4�k771�b�#�5ʟ�W�+Nw��:�
-r1z�^���u�r�d�[W��U��������{ 3�:�*�1/��ڑZ�8Qu�[Z���HV�epq�@j�E�����+��؞��y.�0G( �nכк�7�����:�R7������M�i�t��5W29���W�g�v,���R�k�����MxR�U8K��;*�Ƅ�T���d������[����*����s7��ir\����2����5�r
4�+<�9���PEX�>k�a,��s8`���ݾ.�!���w�JC9j�s�.m"��l�001�#u���ޝ��-�X#W���l��٧�Йg��3gS<ӓ�΄�Y΁W�b���T��Il��gr��D����7�Y�7љ;���s���[\��-����m�{:JΛ,7{�p�3!�n��b�㷉���V+j*y���`q�'	�`�zZ}��S{���d���W�"�4�ɬꀻwS;#ltɹ���
2���Y�}{æcuά�v�0yتz�{�-"z�4��W�^�FS�̲�a'�g^�sGJ���ˀzL�ݗ�T���Q�g�4GF*�4c�� ��˩4LG�	Yt:�2��Q\��D+����~Q���j}V���� �����*����m߽���p`��&$�_Zx%��A����]�r�d�DL��6%^tq���6�r�S[#��&�|�q��z �
�s&t_`M4�����c�H�����#����v��'&s9�mc�oBRc��н�(<��eK%x׳݃[�/ֈ9=o�h�H8�=�W���{��k�������a����Le�)3\�\��o��1���˕u�j���˝���I�%�8uof�#�ލU8�*q`�5�1���9��N�%^a�X���G7�H}O:t�\�z��e��;-�ӕeup<�/��x�u���0��U�F��LO*� ��u�Aרܭ����/�lV�Ӵ�>��Dvrz�s��]뛍ʎ�ͧU%[���m沵�#��3=���l'�s+�:N�.�:g��_{����$1�2��T�sݻ�{s��[d��>��3|��[�O�#�8�y��ߥ3�<�fO��sH�؄����q���cs� �N���+�$��o.ă���l��������#��(��-�\���L�k�,� ��OJ4�=�&q�=�ޢ0M��#=~�X�Y�Mv���&r�,,:9c��z�˝�!��9��?(3�U�+��ہ����$��f���:�DH�Yi�;RU>�v�=a퇒0`����e��fڼk#md��T+��1j5�@ji�c�&�q�xVQ>�Y֩_i���I]y�w.x�t��,Gk���j�غd�ػcD��sy�%j��J����Mʒ�%��9/*�E�͏Z�3��dT��E�1J�D��-˅5)m_b�Y��v�:{Z]���"r׆�♎ж�G��$�"���e�9R*����B��ہ�x��t��z���et$*֝f�r\�P�L��}�7n���	W�}g��c ʘȓZ�1�����"�a����g3P�yK����C;�iL�|o6 �+�VT�C��ogj�ۚ�UL�����N2Uż��Y�.��S#�.E����JN·Zn��5�P�pns��:����}[<�����f<����O�i�o-�4zd�"���~y� Lh�p��8��,����Owwlu�P�n1o;+����7I�j��U}9�wڃq5��a�7Q
��2��j��IB�"�����,f��ɢt�ʹ�Z����d��D�QU�^��!�'�_ �S��W�o����:zV���&�i~���eO@��sf,�T���G˕���>ʌ�uN�5�p��y=G���Y�QT��Tvs&��vR[�h�1݌t�8�w�
��8+�ܷ�EM��_�cX�.RK©�6�z�x^fWi���N�63_E��k��`S������݊�A<�p��n���g�i�ͩ������
���#]p�hKv.��:�ԥ/�w�B��.q�e��bJ��\yZ�RVV�WK��#����
��U��s�8������G�*�G*IR�	�ئ�QJYt����	uժ��[rs�lCF*���93�j�ը�jp�6w+̙�v)S����L�ΟlٵZY�����ʃx^�"�}�SA�M�\9��0f!}9�/>X��y�B�0�m��ޘ3s#Ŗj�n-����Uӆ�B�kz�Q���q�Ee��ѽM�u����sWhE��m����������nG$k3iT�F��Uj�������N�.}��׋�ƣ���E͜��ѵ��P�s���I��uF�ux�ɮy�r��(�ÂVJ��A�UX*�f1**�*�JʋaZ�R�\Y�b�RT*(,0��"iZ�T)l+ ��YP��UDm0��w����v��b�;Ɛ�[�M��d��(Z;|���zʏ����^�� �,�t��xB�DT��Y��7ӊ�{��yu�hVFu;b2P�ڬ�p+V-&��?A��p�4jO�WV1S�D�+�ʓD��wYu�����Z�ʩmT'�� 265���uØ5��-�{��7�b�Fk�-q�&�oc��iyM���>6Ό�S��Z^�8Ͱrһ"�=�X����:�R�x�W;�?ȋ�y!x�t���Z�nmD[.S��RH*�d�����X��y;���9}��v[F���bwXH�M�эr�&2�*iz!syJ���|d\��{}w
�"y�\��W�EF�����f�÷�z5�ʺ��S�e.��$��{�/j��n1ҽ1��
(n�C1�rh���Ή�.�7B��i��T��T_d���;��;��ϸW�L��+m`��CQ�M���Y2�nMh5F�E�폋�! �lu�y��Ԕ�@o\܅�\�-蘁��WI���]Z�:o<}�N>|&w��Y��9l�&�c�G��s\�G݆(W��ϥị��g�0�LNwdW�.U�%���r7Ej��/���r~�I�qr�r
v"�iq���)��^�3�l������1�֩�Z�֟얇oC���R���:�+���U�n=��E�R�н�_�\Eb���_c�+�=���c�&pxz.V����2�o]�n4�A�wRnP`$�F�����+��w��t������{x[�@���y�&�^�)\ɟ<�`�>WoE�b}���5Y�/���P��{d;\E@�7(�;=�\٫�M��.�@���x�&��9)��CE��<}C�L�ˇ�ew\I�ek��2���$^�,.��XJv\Ig��$���k�@f{@��
u��_���x[έ���~J��+�=@[���4��9���-	��q��$μK��F�'���ڮ'.��&X���9��4���������yNq�پZ|-�X��M5]�Z27^���M�4r�}��y:�y[�W
;����D��r9�\�vy��k���2�>�|��׹@��Q s������ׂ^���Uc��nc��k��m�]����<�^��r9�F�j�e�aŕZ�d+ʃ�R����1G�Ji��:�쒮�,�(�r�m$�%
ѭ%f�>��!G�v{1],<_ZEfm���v��nk� ȅz&�Ô�yƨo��K�j��{��k���j�W��r�R���%�Ҙ��f����"����j�hVX�bLf�*ۂ�Ø�P�>�C�D��s�����t�BU늍#ER�1I>�ڰ�j�8�t�\������9]���B��I��U˦ɐ��:������au��-U�nrO\�5)I�re��}w�^����w�r�����������¶�8�܍�����f����.���|`ĬG�d%li���C/I��J4�u�nF�P�o4�ȖNˊb+���C��v^�V���~�3���&6f���]��w�\F������t�M�RD�U5B���Z���/��'v.�óC���U"c�z _Q�T*�Z���_S�V�e�ѷrAxj���W#o7s���g"�,�9^>�ގIˢ��7�[�AF��Lv�q���U��/B�=��*Lc-��.�z��*�Suݓͩ�mn��g��Q�]�k�Fc34t���}�U�J�כ�Q�
���3W��i�4�#=�-��5�X���~�7���i��h#z����ø@�Tr4�b�0���y^e�l���}ڶKsk�|s�Y?)#�g�<�L5�S��r�|4�0���3L���Q-�I�B����ۦ���]�_�֯ Xy�X���\:�̂�:2��~ʨ�;$h���=dis�zp�Ouy�z�wչF�'7�D�&�BR�}��lrP���.EɎ�1�y<��wa�s�3��Of:o/vs�PFdeZ�o=9��$�7�u%��#Gq�sOC�z���q�i����v}���������pVﻸ)^�v��f��u�vn�El��!�v���W'4���=��E�}��;�c�z���v��H����O���+Ut�\VU�甲L�G+�j͍�dFy��8+��=��F렪�/&���M�D+��=��h;������*F�1X�<y㒌�!�v]��G+gbf(W#ƧN�cK[��pl��+%2y'�Z80�d
�jҚ��>�d�{��=�'~��!F�U��t�[���lV)�ԫ��4ӕ!�U�k�rn ��Ţ�v҇Ej,)t�<��d�W�gA���[�4��$�t�ag#ǲ�,�f
j���K�8,m�L�U7��Ҩ(�h�hL�9
Vdo#3�K�	����G���p�t	n���T�pU����Kz��V��ښ�u�]+�iL�)뜭�#�8k]s�I�����7v�1	�@6MnY�Z-AZK��z�a�`�t�H܄Ν����Hk�D����T�<ɯpBk�O�73~�WH-��þ[K�*.B�/��k;4c��#|��S\굣r���.�FU�V�7Y�{w���2�A��+�&�uc�qLU;�vA�������6��T���g�ҬnW�w%]��#GP�Xfɔ{�j��ɢv��F'�1JڼKA}�B6^����P�xD �f�&6��\��&��.6e�����"�z��W]x[C.���#���\�C0Q�;��έ�P9�o�]Wp�f򹜍dnG$k7mT�E]�F<����ޡ����=�"r���遻b���LZ���޾<�|+T�]�y��q�8�9�y��c01T����--F��d�jV�QQ"�
�ьQ1p�0kY��b���#q� ��D�DUqJ[V*�����	dV*(""bѶ�
���(�^��y����:O#�δ��HI<NT���Fk�K73�X?�7�8�)�(<MuԍOO�@oS�W#�{6����T4k0`A
q9�[U�l�]�f��h��auq����3�6�m�1S�0����+�J��y4����ݕ�Qm[����,�:�+3�6��л��]��qM���!�j�3�FP��Z�ܑ��W<�J$p��fB�V}l5+N������]^��t�~�U��wU��(Ѻu�����;����R�eg}��9-� έ�|���v�.y��6�,����u"`�Şu�'jĨV��Y�r[tH�������bF��B��T�3 e��m�8�E[~fHW�9����q}њ�A��|c�ȝh���
p:�3-�є_J��A~����Yy���VqY���u��b65�tֽf�p򞶒�j�zmx����S�Iܮ9�_9����](�{�s�r7�S������K0쉔�q2��q�]i���T��5�OT�_NL���4��x���	��[��t������v��[��ZaST\ы.���3�~��椤G x]��c�O60p{���c"�����s�t��Q���F��I�u��wt��#,9��Dm�m���	2���X	�j)~M�M���q�˰ĕHө[:���7@}|�ַH`�K�j����Dv]�������;Te����v(�h6�I�ʚ5�5���[����p������BҠ�##)�U��V�R��8[�	�v��P�᠇�H���f�uƅLxX�|��t�¸�;0��{�:����a]~�V�#=ռ��s=��i�=�2��l��|s4�J�u�Z;�z�|>@��#3;^�7�=�u��*��
���zzɳ�ۦj�M�:r�a�mV��7C)^ѯ:��M�BAos ���挥��V^&<o��"I�u-흜�{��|��)ўN��}���7�v2�#��Rmu�xI��-��M(��ΞA�ŵ1�1���"k9�aaɵ.���;�=N�8�=���-���OP1�s�ľ-h=�}д����9݀Jt��8��8�CO�d�C^=�5M*T�>gM���D�ۋ۴��5R���t�۾c�o���+ʗ��x{�I4GP/g5��u��1ptΰ=�vuN2�z�\�~7�/+��*Y��;�.]P��P��L-%P���1U��Y1�m+b-�<�Ƴ���"3����{�ų�V*�ũw�@_s�y�+B�/c��/�6�,�����6�1�a�+�D��slf�݋\�������Ld��>�f<�G�wk�(�'7}u���	-��\X˛�u��d�^>�����vOom�NY���.Lv�5��Gl��ZNײј��л!j�*o]�F��E`�լm��䈮�M��l�����H�r��Js:�7���Z�#1��sc5��aTov�S�u}Ž�s����Q�������k-&��Ob��&Gdp�D�y1���ΰf��]~&gdM���&��p1���3ƍT��!�5f`���xi5�6"��M-3��c(�s{��~�v��6x�w-�[t�m���'o�U�̎6 e�9���?x�|���{c]����u���N���3�kP���k!�su`���^�|�����!H�l���0̮Y�x*шB�1e�F^���8]g+������=�|Z��i:���[U+�,���(�L�X�KQJ�]vwyeqj=�P9�Xsms���]�x��*t�{��(*ɇ��Û�_8��47�̘}��\f7�hS�_S�&�fG.m:�ٵWT����V�3b�{qVG9�����;�E5[q�lf,Vp74���۽��n�t����p��n�U}"g�D.͒�ӄl��j����/�o'[���?Us���Ղ8�+}�rmҝ���PWb�shH��/l�"�o@�`dc�Y�E��;Z��%��U�R�E'��v\�vs٪W��>������YX>�k��!|Z���f�h�ː�_������Sd���hR����z��D�w�b�r-���z����뎅^=S$?=���������H��{,��Ǐ���U��<ԫ*�n��rD�,�[�E�˕mv&�n_>����hѭ�ʅ]�82qpd�D�X$}Zr)Ϻ��h�]��8o3x���壌�ѥP�ӏ%��'�~26�*�΍+���hk���>�:�����sx+�ɓ�+��Y�;a�qyF�y���S�
Z�(+؃��̃��v�W�c����c��@�&;��?�����}�`��j�����[!@&|�"$~?�
N�@�	�qa�F�C�8`���,8y��=g��3��bv'IA�	(I	 qd$$�!��dcs��q��),5y�X�&�Ґ�����s+�a�Y/v��!��	 �x�}N��>��}�s�����<�����?B���ɓ!��C�pP���7�R��Lx`�R��׋u&���80w����k�H?�C��|�}:��$I4�@�	���D$$�| ��`�C��׏�B��?��y	��2S�z`7�!�|��I���>a#O��B�M�������}A�" y����	!��~��Hj`%9�g��2A��)�	!ǎ!o�c�"�{���|؆�O���\�s,���JB�D���gq&z�������D��	 �C�q�aĒtUHrK0P�z��0���pC�s��?���>�$z��C���S�r8Й���@���?xC0�F?��Y�2���=��!�	�� �? �����~~!�����#)$	 ������@��!�9>D?ԇ����prp����>�`���4��"�������.I�!?�>A���=A�I'�s�����4{�=`|D��_�D�C���&͆Ca��@����Q��qꐄ��`?Q?�?q?�A:'�B|�����Ȕ=8$��	�0�!�2����`���NC�=�D$�L��!�͓�D��,2Y2M ���ɐ8��;��qZ������B$1$�g�&ZC��3��s ��|��� ���G�|ϼ���}D Hx�>�O��!�?X�~��������z�$�t?��{H`$>��=�zR?�������������C���!�����!�q���R$}G�{s�=��/�BҐ����7�!@%��d9�������{C����~���!�=�L�w߮�k�6!�1�Jp1�L?3� g��@>�G�����b��R�~��!�tv�>�>��rB�L|>=�9�(k��_�9lO�AD��A��������QB��s}�2C��L�g��!$	 ���~s� ~�!!�?���3�:�ϗ�I@'�O��	�NI�z0��i9�<�$�`gX����2s!��A|��Ĥ���Є��5?�.�p�!�U�