BZh91AY&SY\���_�pyc����߰����  a	�                �   P      P 
 
^" �Ʊ�j�a��� y��      0���}�������]�ݵ�wQ����x�z�˳r���C��j.��t�����h6��r��8��(v�Ѫ]�s>�Ίك���^8�m�`��;�z=굽��ڻoO;=�n�#�z{��;��"i��f�݋�ko�m� gr�g]ڲ�{�/yu�unۚ�U�F�pz
�b�w��{�m{4{۬�<x�oF61�s�Ŝ�{i�/f�P�ݵqf��ޥ��+sWN��u]ޔ�x̵{nit�׻��D��*���7�ڻ;��][�˯�y�v]{���O��"�� ��s���׮�`P�λ�����z6�k��y�����玏ym�׷S��������T !���u����u7z�������k���,x����,�Pts�k���]�C�]��ӥ�Ekzn�yG�z�uγ�Ѻ��H        Q% U  )EI`  �    ��iJTHhщ� 0b  T�B"%*��ahh���h���JB*���� �   M"@�*Ca4�F� L�0�I ja1Q��L���MM1T�	�U(`i�  @�i���H��
�"�21i9��9*��kDTQ�T�D$Q����@QQ�UA6���>?��
eJ%J}�*�5�� �ߥފ-�ڴ�1p ~�2 @��H��F+r����CX��RI�nATQ��cLB	`UURI��!XH	����I���+缝|PՏ�=�l42�PQ��J~k��|�1b`�4��2�$�K���CI�X�>!����u��bdq���2��K(�̲���\� D�33��H)�)�!�c,���xD�I �xf2I�ã����{��e�L2)&>�"C�aI�^;C<x=WS(�2�eWaF\).FS�H�q��\��&D/u�LmQD�4���Gɸ\g�r���p�ѝK���(p�1�3�.O����2=�O=	���兌�X�,�ǎ�:1���F��@�23�G
|�QHe�	�1�>c�C<I�X���S����dd������4ҡa�����$��|L��z�<>�1����I�# gG~��t|�p����
�x�	�F$�"�B�0v���#�H�C |I�a1�B��&c�/�8L�dt�E��������ux��/z�re���&X�a�������x���1&[RX��d<\��`�H��$d$�>R�X�1���A��$�0��LIȊ�Hb��d+�G�g!"�1���I�#3#�����0�L��'.�@�B�X{˞`��]8RL��k�hJ�C��g�W}	�|f21��c��G�$P����L�!2S�,,�����1���aDÅ!��7�I#�,	q�	�1�i2�.\/ C��2<�&t���j(e��c-�H�\&{�I�1�²O�1�!1�1eBe{��0sP��j�P��dc�э�+0ļ2S�іO\.0c\\c.f���ބ�w	�e��Θ^8Ta:��8�N�	�X�e�C+Y�L���YT�<6��g��@3�����#�L��g<vg�ZL�dt�Ҩ�0"��1�eu�c�B�'e3ô�x��<0<aڢ=�1��lf�D)� �&!�/8](����K�PX�a?z�1�M&"e��e&C0eΦ3��B�FX���%��|Lc���wO ��p����')>1&N>)-��ҡP�d3��L�{i\L(<y)iq�l�@��d`�Ld($��
�2%rI�P���a���	��p�!���<?	H�i�7�X"e1��B��mYdӅ,t�%�.teє>�1��ĈKŌc���L�Gڄ�X�=.�B^�5	�fs�,j%1�t$�a,K��1��欁��\�1��	�c�C(~AI�g��Q#,q�D q�Lc��G0gN�#�+�2��#�g�3��"�#����j#�Ώ�PǍD�!X�,�R0cRY�FV$�X�#TPΒ9�`��P�0�������3�xF>�H�u�a摃,w*:2G 19Q�3�<�C(���F1��Q(��d��1��C,�I�2�Q��2�:K�F2?&`�<8⑐!�S��2�S��c0g}
 c�P�֢1���S�e��ut'��c��mE�W�F!;P�[TAO��1��G�H>bT5�Hd��+�tf?50��P�u$�'Fy�P�[�f?b�`Ɗ C;�\����da%���c0���4c�C4�p�Ь\��Ə3���W�e�%4.��FZ0a\�Q�	!�2Fu�C$g�(f-�3xo�0f���8W
D#	)&Q:x~�L���!�M�ae�Bc�BfZ`��A|���8L�N�!�)�i��Մ�,��R��i���fq(p��Jy���u�v�"IK�%�"��S�æ>,0fJf�c��UI<aa�B`��C;)�� ��0�!��	CڒH$hGFAp��$1��F@��qA0�r�+�~L��KȎ����"DY���Ν�L��я�I�Ptc�ӧG)�e�P�^J���x�b�[Q�G��]/8P�G���c&1�eG��Lc��0fr!1��C��a��1�DE��$`ڣ��p���H�i.>���I
$��2Q0��C,�n"�Y�KĞ�2���Ƥ��3��Ύ�TKJ�Pt��c�w# �(�%���p�g�`�u��w�C�Q��q�6��z�C�0v���P��>�2���u��֑=c�2Δ�,d��E�2�cȌьm�d�P�(�F?LC:I��L��>� c.����\gFA�Ld��X�,|����H�$q��t`�1�P�}!�t2YC�#��H錒�$��d��Pt�>L0|���(��($c^���N2��bp�e��
�Q$1�X��S!�%�C<N2)��{�R3��C:u�H�C�{QNH��1⊄&tư��<3�
9d�C<��u�6�pO#"9�_`�j��ֲ�\�bAD��@��"�(�A�!�Xb\��.>>�s�㨎1�A�@�/��$���c��J�j�$�H�WᝄΌ�W�t� çZGFF$�#�A���c�FJ,q12�6��ؕ�E�Ƅ�c���1��Ę�1��Dy��]"b"�+���,d�Q�G�3���:2��<`�1�:L���I!�	�~Le�$�B��y���(c.W��1���ڢ|L�ͨ�1��	|^C��2Ң�aT1�tC��H��&�O��;P�o�,��x��$�mY�R2K�(�Z>[QEt���ڥe��agK|\fo�0e�%G�t��H�J�0g�(X�RA�QюSڲ���t�eq��LdWD�1���.F?&xc��*"$dq��*8���HQ���rJ-U"�NE��%樳U���>4kB�Ҡv���\:�,��2.�O}mݻ?�P.�5G��;�l�N�˄��R:�95srs8��%�dgy8w�`t�揙��t.n���߈E���}�����3�vYV�?�wg����'_���ܻ�7y�h����N8Q�����:p��u�=���l���Ŋ|陣�~�}��6q9͒d�d�%�Ss�C�����y7 ���2[0.F>ݗ۲3vEs�y��9���=��hL6��G.d�E�s$ʫ�9��]���99݄�n�v���yy�{���=�6.���NZD�H9�Nsf>l���Ϲ�����0��e�c��Nft������"�e!��v�L.\3{,�9S2����sf}��M�˞�����9�
�W0�!�2wt஻94e�&�vY= ��gd�������2���+�p|���u��嘝S {7����8��}��O����;3�s[��˦�@��O�gw�����͛#3����w>�Ig�ҵ��0f\������)|̐�>f�u��r���`��3��}%�oy���`��ŭz���Kp0�N�����rh��al�~���>߈j�~���2��'��(~���8�,wڹOvz���<�%�N��1�IҙL��oƫX�a��e�gc�o.'�Rn�rN��ܲq|K�b����s���������}C�9�b��iy�y8>o�fL�y&󙃉�׸8^d�͞�-��N_"%��om�Ӽ�|��%�]�N���}_)_R}I��[�
�򼙅V��"xcX�潺��EGk��k�U�o78��89̛��W-�Ʀ2Z5_|�C���T�QNUԝ�w���fWy2^q���v�l欹r�V���2od,�9�l��˥˒�I��|0��)!��9��Q)��Cئ����b����l�vk}�h̓��`� D�����GG�9�=7>��b��dRz=1�ǻ�����n38L�盻�9�仄䘱�~nnV���nn�5?۲C8���Z��Y�+������o��1��S��I�-�9�7Gb�q>;-�fLm,�;�9|�2N�R�N=�����Ӹ���]���8S����=��O㞯{�9�`b�跚����rv��̒W��7ӷ������zޛwx���yɻ��3��l������1`y��t�֯����J�>�s0��zZΝ�̙ο9���`Rl9s;�=2�ge�Fi���{���]���JJ�A�:]$��vX����#�zd�Ou�I�ZUK��l4�:���r
;nl����m2Id�)
�'���K'ʘ{�Wۦn�1s˖�ё�zxg��Y��⅞C����[?bü�﻾���|n�}���k�7/7ϳ����'�0e�wߧ=t�tɯ����lz��4�<�ec3D�i �����w_k���ݞ@�7@�YM�ʱ�ǃ�K/=���;�ǖzyV0s���)N�g�80��&�2?QG,�ɺ{l7'$�Jnb˝:V���`iQ�2������SEӍ�
tw���'-�9������j�;���9عO����0?�6?�O9��~�\�����9 � ?s� �Z"zzqf��Y�o�}�?y�2��w&,�Nf��>A��Mm��%��ۼ��fn����>pKz�n��oӓ�y�c)���Ø?g�����=�-���g=��������{!7����3���!��y���#�̙'�����t gKl��e��M|�o�!s���r�f�\i����}�ϻ���q���m��Ha��}~r2I$�ߺ�гU�<wUṈT����<2�G�{{�J����&�d��ziܙ$�V�*�:�qNXfK������s�{�N�ư�Dc�92l�Lܜ���O��vHw����]����=�9��G�N�Nfhϯ�]�.?M�R[}�nL�y+;373���w%I��'�Y=�6_ɜ�q=y/;��\9���C&�z^I�vY#�}��	�����=�rH=���e������B���i0p���w%��Xt|�2q��wsw&a�6ɒg!�\��y�U����7�E���f{�b׻�!ܣ�� ��|�|�&� p���S���Ϧ�fQ����|�ts���8�<���3�X��rO�kfs3۱��_d,��͓7��;�y^C�H\���Ҙ����m���Gy9���-պ�\�>l��T��(P�Q�7O��2�-G�D�3���i*]8rl����I�d̐fK$���JW�d�7/2FcD���9'2jk�9�C�����gH�ь�l�2�>,����a{�[?f�:>S�y���Y���Ϥ�3��ݝY���/�f�W�����i����.�:����9�G��|�ܜ����g(s
G,�%Yh�r}�a��wa�k�m������80��ٚg��ГI��>K�'�e�t���wd�wB�W�:0�sv���eX-|�|���{�(�v3I$��$�ܞL:3���nh��	���?�������')s9�4�t`w�GH����q��ܐ���(vN}/�N�m�^\�0�F)�r3
~8nh��gO)U'��˘󿦒jҴ�2���Ϩ�Z���}�;�ꯅa�s9����o'b�/~�
�����f��Ϥ�'{�;۹���p��y��ۜ�{w�ɬl���Mɧ׷s���'d�rv8e�9���{d���ǳM������L-��$_7w��{#���S_��.��)��볜�>�I�76��uIѧ�����g۲������ |�g������K��gw n�%�{9;�KI��)����V(샾�C�͗�M�dr��}���#9���7�0����2d�rB͗�
_���3�v����V�Q}��/y򐣣�����n�ߧ#&w��X�g��>�Μ�e�����O�$)���C�o��a���$�$ч{�w�g�pG/;���)�����8��fHb�ᘤ[>쓖p��P�/9 $�fnk��-�d�9�i��y9l���p�9��	vlM��~n��58��{���S��cw�f:�&�:w|�wN�9��$�i�]����߶k0d�;0���$����=��u�T�",���{�'3��͓���W���Y�L��6kz���1�zq�0'�E��p�}�2�x�q�Y�=8����:0>Ӧ���sHs����������;�P-	�%��ݻ5�I�09ިɼ���rn/xtq$��H���6�%�4�������k�;���AL�֭���y6���,�{$S6ČSkrv%"��lg.�嗗cf�6�:̍��Ǝ��������oM�b�`�K.�c�լ,h��ڈ�\�2�2���C:Y{��̲���ح&w��2ԓ>Ηq��E	c+�:TԌ]�pK�{�uw�D��G]UQ��(�#3δ��k*�c�Y(�
�������"��G�+S+)Uq�^�$�R���M�ݎ�:/�Z�}��/|�o��`�yե�v	k~��N��BBĮGJZ�l�������bakn���ݸ�K��Y��h��f17�`�u��T��
������/��\1K�/�	/O<��>��q��\jZV�Vء%r�$�@�ܐ�Jji�V�v��"zЈ�Q�@zp+~& L����E�
vΏ�����d-n��#U�	$u�� �$d�Ċ輪���s=͈ȸ���ip˥ݑ�.{�
t≳�-��2��0(��D
��'��-M�3l��^%^O%T�Lq8�)l�K�^�'���� �Z�l�>�R��N���.�+t�;6_�����b�[h�&Y�#X��z�@%�����3@`C:Κ�{l�uմ��鴥��\������[��
�l��MW*~/���X%�L�?\�%g��nA��x��xb�P0X7e3����x�T�-qF��;p��������s�5U�
�Z�(x�"�O8h��PԘ��hm�{W��ﶽ�����ɼ/C2�9W�����8Z�q�2��V
wo��ʇ�e$ٌ�0])���	#�(Km	Lit�79t�7܋�LI��`@�^��!=fwI�v�)[d⒗ڗ}3��}c,lt���#�V����0)"F�띃Vj�3���93@X�]�g��{ĉ%��9��� %1�fϮ��\I��T�0G/m�S"8ཌM�b\E�v��E��6����俗��z��]�g]m݈�9�7eIN��_\�P֌�Vq��>7�|�8�$pb�}>�J-��.7X�<ܱz�bi��b�(L�.�ҕ��r)٘U���!���v<o�
�=UpPU�kI_���;ipUF��_�7呑�Y�	���s��f� s�ETf۴5ɷvɐ�����ᙾ�*��
(�}�md?w��zϏ&� p�$Y$#$A�VEI��G�~�����_����Y��1��m�M�ߛ�nm�lm��m���v�6��m�6�m��߽����v�m���6�m�p�r�m�m�M�m����{�����UJԡT�U��
(�H"(H
� Ȣ9�q�m�6�[p�m�cm��-���oͷ-��6�cm��m����m�m�M�-�������m�m�Lm��m��ߛo��m���6�m�i����(H��
���2(Ej
$��89o��m�m�m����i��m��m�m�m����m�m�Lm�۶ᶛn�s���UUU7m�m����nm�m��m�p�r�m�m��m6ۣ� ���8K�����ڥ����M�ۦܶܶ�t��m��6�m�p�m���ۆ�m�m��4�m�*���m���v�6�~m����om����nm�m�-��	�P�R,�dU�RE�- )+$� (���Y(�6�r�<E`���������v� 5�䛷;Ü6��9Q�BBf��I<tc:3�<bI��f��33 ��2O��'�HΈ�1�d�1�����3���@��,e2�YC<a�Kt��c�a� a� `�!�gFX�X�XΈ`κ��ӥ�ɖ�Z2t����!�d�c�`�" `��C#$���ь�F1�cc0��2L0f3a����"K(d� c�3��1�n8��^Q��=��O�~]S���3�}kQ�a)��;ABd��{s�-�y�f�e ��p�+��^h��o$��_Ck5��l֓ �c���f�/Sj�Z�5�ʼ��6�j����0�)�l�u�vv�f�^х��U�Δii�݋�]r[��f��&#�u�e�?Wh襭!cS�� ��[4�/��{��a��Z��o{�F��H�,+���yM[��u%#�m�n�b|\><H��lYcRNM�\�"LkA��
"�3tڕ��Ɩ��]j8]��L��I�����C�h��h��m��)SF�R�Z�:�	x�����ֳ�Wk��,!dK4u�pR$��j���)v�3�bd��g2�UYK�ǚY��%�e��n�!Pt�h,@�
Vɬ�����;5��Fٸw8��ԥ��]4Ũ���FՄ����aKXn��orYz�L�؍�gF�K�,[���^��̌�Tc5W�q�4h�^-k]����N�՛Mv��f�!!j�.u5�:2Z�n��e׳M4m�J�4$V�A�:�j��nxI�i��~��ӳ7�þ��x8�e�\��Ffe�XSp�6h���
�RLh�Z�G`��]���׌�I)m��ɡ���nve�%�ғ7 ��GX3l����9.�]�H%`X�]��|΃��������h�V�&���
�m4��ֵ� �&m��/�	��o����au:�K��P�S[-�����0;���ڇ1�R��.иMa��3,6jI��hWR���Y���S$�9��S&�Y��ǳ|��}fE�&�L]H4f�jC3Â]kZ�����D$vnJ��n���L�Y�]M(a`�l�D�P����S;a����m4�6�L�
Z�l��ڗ7j2�s�;#ef2Y��i�)j.�r�;hK�!�[h�V��e���R�JY���JY�d	zʄ��Ycp�k]��[Ycm3f��l��:٫�u6�o�Mg��#�sZ��:����_���s�9�C�k�n����x �n���m���o 9�V�������ևs���������ց�49�i�3K0����C#$�'�2�UǚJ��zV��s4δ%�i�LR[�,�M 2��F�w\��%K4�i�Yn�(��5�ŮK
R���s�v�[3ff���q���J1�;ZD�Te+�{m�@��2�v�Z#��m��5�\�pƆp��N���4��A�8���Y���{v�טvظ��45]�0͙ZK�f(�E&��(������`��yS0�z�=�*mV�~9�Y%�M��hn�`�el�?�'�Lr%�L.5�M���2�1p�m���L���kSӸX`���i�<��4ɞ�r�T#�����Z3Ki���C�:{���Jd��U�tʒ���)��ꏧgJ�A<̩Z�q���i��>y�|��]q�C(c$d�a��	 V/2�p�VM�G�w<���l:�O9���%d��I�ݤ���gҚj<0u)�ia�g^���ީ����0��/ܬ�6v���HEc��O���vmO�&�sf�옦-���H��Y<:���:<3�0����C#$�.T��C��+�H ��qv��&��C�V��-4_xQ
S �xyO��ͿWg]"A�	eJ��|�C�>'��R�O����agp��>0�F� c'Y0;��Jw���n��k�'p�zy����Ni�4��+�v�S岔�,2��e�X�ae����a��:R�<���L0` ��e�u��UIKX���ͬ���+�.�4���%m�b���Y�[�OI+m��].���8�g��Y+��"1O���n���r���c?&+q9FQ��M%�rEe���Ip�
���<F��,f3,c0��(c$d�a�8����+܉�D���]/�+ ��1i-�16�Q�cf���1�H���9'1b��-�[v�(�D�Mr��

X�fcbi����Mf�S6��I@~��bQf*��JJ7\��.���(CޛL����az{���mX|�ٮ�6�uR՜��S'�ӣN���g�M��bY��;O�M4�LT����e�af�������es�.����Eg}�옚��m�]K�(��S!�şa�˹�ħi��M��`��(,(��(�����Y��:Î4���Ɇ��Q�i�׼U�;��z^��S	�y�rrw�32�ԡ�|v�;��I�9:�t���T�;�����
�q�B�����v����M^���]�JH�=�-Y0�s�(:w`Q2�)����.��z��K��"���̃�N�x�L�0f����a�q�pG\�fC�Ҷ�䈚h̉�F�ڤ`�t��s�G���F������q��ߤ�Re�c$�ā��%֦l4]��N�w���]��,=4��(�i�;�u�mb�R

#yl�3���m��w4�J��ߚ2Q�q�c�`���kEQ&�^��;݁�/f�;/)�M��bu^�pM��ރ�wCڧ0a��pUY��HYF�X�i��`���጑�a���,d�V�Q�B��M�@K->c0e���c7����[���fGMT����8}���߫���k_O�Ӹ�;'��p�it�,�#x�t�3ľ$$��S4��R�^�<��.�Ɋ�2�3&��9N��Z>e��u�u�\|ѝ�&x��j�aJʎW�";�F��wn;�d�ԍ]�5�H��n����Q',�^�^��l�V�z����p�F�,�mO���^��O%��G1è���|Jio��,+mUU��qc�K7-���a7��'�W�5r�v�F�k���4�ͳ7���Qk����UǑip\��3���ve\<)F�X�ʢ~x�1&�39��3�r.�U�}S*�8.sy�&?P%�YÖ�a�㝜�7.[W2���N��O��w���)��K�6��ͦw������#N��z��L�I��ifa��,�Όd�Î4�U�G�(�4����]�o�COӒ����}>E��O���������e�0�B�=�qi�Wȹ���IU�[f�F�oym��Z����j���<S��_EP�� 
p;WC�����ߞ}�wn�gŶ�I���#�:�������.����]��'R'��i�������iF���Y���#D�!�F�L#L�P��JŢ�'���$�� �gfe��VO��~��_�_///�/f�f�h�Z2$L���4Z#"!�FL#Ef�NF
ť��3�`�:F�6V���h�fvE��M��B�BtH�:i��4�:\-#FkN'�E��<���]���QvtQ�4h���Q���W�t] �$�GM#E���4Z���:M��E��O'�_�?/O�ۭ?3�?,���F��4��F�M:NFA��3H:1��d�bѐ1a���F"͙QD��F�F�H�iDidh�ZH�Y�e&'�9��
���Ɛ�%6Cd�����>ȳ%�S�~��J����Ϟ����)�\��?$���~˻��Æ黻�����wy��7wwu�fff^p�7wwwos332��4(�L4f�1�ft�Oi'M:3ӣӳ��EUa���{J�!�%�J�uD@�R�����`���	9���cIitj�E�R" W�>J_cȾR�T���	�ٽ6j�7sU�~�螚�H������P��i�Tͫ�Fi�G���"=l�襓�!;���?�b'����"�[EjR��R�Uws��r$4D����U�
"y(�l�$7Ɠ�͇e�q�}�i;f�؈��(v�t0�%or]Sԏ��e�ο<��,�N�i&�:3
0���#RI$!�>�Czg���2�t�@����A&@Bv2pBC���?9���pS�c604My�^6�����D�--�)D̹�?N62(jb�@�T�F�Cb)�b"�tX��	��e8 �B6P�<�ڗpA7쐢��s]:`t0��� �7��&��2u�R~����FJ|�(�QG�UZB"���Ԕ|��~�pU_��B¤�OP�����O`�=,X(�`q60��i�4���1�Y&�x�I4�ь���$u.Jk�u뾩Q'�ĵ�m�/1}+�ibQ"��r�*��p���g9����f�G�Y��v�m��a�X����dœ�YES�)[�2�R(�!j���z ��&��Ų�ܑ��W��d�5��Ih�$
Ex���Ky�U_2���y���<S�s�6��@�a;���C>^�>a<�(�4���OV�îBz$�Da���C��=�)`d�N��!DF��Λ�p8r2L��=�'4�n ����4���<�qD��hM;�4|�:��P�`T��0�DHt2N�!�έ�$:&�@�Da;���!�	�$D���`jq���,�qv�9��)��˛�{7�
���	�$�ya�I��&!2QLH�{O!��������)�6�N<��`�,�M<i��x��P���_+Ԓ�"!1����2h!�h�""T�Kd7��Q�����v�d8 z"&0�2Tؖ"�=>��vJ"'^R�/�Wߘ��멡K��%m�о����f�VWnYna�uЩ<B�{��7'{zI$�
��A�FFON�C&�=m�6�39p��L�uG��9P���DF�����5<9���+�D�9x�Tf\/I�~0d>�i"R���"C'�
r ~�p�yZ� v"$�!>�D�������3U�k��9������x���i�Ƙ3
� �N�i'�e�[u��=�b�H��N#��рy�6��؈��3F�0�Z<��"bC�
��'�)���J�m���+��!�0=�
��DK��ξ���jTܪ�2_��Ne���jFRߓ�!8���y0��T��9_U��DA9�`h���2),,2�N��2"DN{�~�'�����1pV*���JOm��y(n$<�l�!�a��Q�)�Q;��D�$���2]��2��a� DD�$c ��8%d���$\?�`��?|~3
� �Ӧ�I���e�t���g�I$!O�`dI�'���N�ZCO ɂ"I��9�B�`VHQ.w~�g]6�Z��naZ�[T2N�JS�`TPY%�����DDܖQ�<�fj��R�\G�Ɂ�v��ԋ� �S��کa��~�|vY&���@�B�`��I}~���r���E��PB6f��N��J�rɐO�5pHVH�JP�e�M'���h���}Y��NA<��0B��2��S��a؅L=:
4��M>0f1�A��4�M<tkի��~�g����U�q�W3-K+s��D�1��z��$8��
���y2
|x��Q�_4A���V�r��!`���bq�%�qYD�ȿp %�Q�u��~�ゕ�Y���˱��69�u��r`�_3k�%�<�q�:���(*X~��(��#`�2}`~ޅ�]�a�,J2 ��!���I��H訟!;�&�(�C+�Z?C���pD>a4� @�e�{C|3���������������w�w���ɪ�3��)��vț��o2��&M�ΞW��=��s�ӿ/?D����ђOŲ)�BN����~˖��+�莼�G2�I���}:� R�1�(ot��&��C�r�?<���n???8덺���/<��2뭺fL���9v�X���ڪ����ia(�xZx!B��D82��N&b"!`X��jQ
�����D����T�Q�bd�Uz�� }|��	�i'�N��ޡ:����Hr��F�������Y�)�jid���p�!a�>N3�1�!�r�J��7Wz&�V��i�(�E��)I�# ܠ##JO�NN���#K��UĢ�Z�y(���ld�	�3��؆	'~����j�9VJ���5RV`ۏ�3��aC(di&�I���e�$��UF@D22DD��(~"����W�f���9%2��P��E,�0:�-��`J���뙻sc����!�F�� D�Ru���~�T&8&$0���5�t�m)j�j��۔���^f.-1���@퐳߇���؁PY=Hu�-%d�I�S�b
dN��=ffg8	:�Y8�����oȮ/���|�JkRt�<q8(s���C��.�:�k��$'�J�|�ar�C?ks��&�+4H#>������*�==A�DHpa<�(XIKEW�H�O:������N�4�4�O���I$�sx��@��A0a� �$6 yC?I�c"���s���e:����6ŀ{�_W�m�|���Rd��ů1��,,�ک��]��Ct�Y�iU_��J8��e7F�ZC�O׶;3sxd�v�pHKR�0d��D�J!��'�����4%��5M:s�\��&��R�.(6��`f���œk?yam��J8p�=d���&B%��
���,谘�� �ߣC�'DAG�dD+"����`~�xu��*��/�_�i�phߖ��FG��KH#J �x�4�I�H��'$�����Ѥ&aa*�i��m��k�K�m������I �t�4���]4�D��	1H��1h�$h����,Za+�Fa6*� ��f�'�|i���������a<��������N�,4�A���h�'E��Tr>��7�~Z��}Qt.�mUr��6�z�yh��ˍ��_�[����y~O<�'�+��VW�ai���駉�x�>>#���_2Q���H�H�h�0��CD�Z���dX�4�4��AQ-�
M'Dx�4�4�e-6#������6~���G{~��R*	<w}�b!{_�dR���o�r��Vρ+���x�M�Wx�����0�/��'����_Z�r�m��K��$"f>��z_k¶ʶ�VYkT��L�o�0����~�|#<��*`�U/��X����0�n��`W"�A�6؅�Ac�:���2�QG,�{	j���X����ʦ'��9����3�7*��|����D���ݚ,�[S7�L����k�n�g<�㺠�8�F�q���%ƛ����t������r#K9� �㗙�5V7�L f5"l��vm�6Q��d�z{�^-}it��٬5#|��	RYi~/����y0��,�5��Ys6u�Tu�:����jR�W��_s�0��[v�pk`a�eԲ��J��h+ipZX`d&G�<�*���S��MLx�%�����Ħ���6�Fi�Ս�]j�v[MPsI[�����t<�����BR�Kk'����b6�)q�F`p�.�pLs/8#3��	��ٙ��~��333/t���ݽ�����[m�{�������n�333,<���yǝy�\m�N��<�/*������d��:���R���"�׃k-ƻ�����e!�y���{��6���dV�J�K��f#�2b��]f:ͩp����\�G`�h�*a�K�V-e$��շ�J�\�#�q+�B��׾{k7qiR�V�Ms�T�u�����6�`��xl�17��gˍ�}-��-%��#f44ɚ���Ci����,؛d��[OB&
)![(�] 	\��E���U��ҝ����ކ� ��2�VU����9KA�N]Z�u�W�J��A~0�p�E��B��4a1�%��9��&��0��JC���a h�Ȍ�����	=����:C�0�x!c�2{1��S$:���X�p`��h��1|Q�������i+� �Ӝ�t2xЗVwcy��Y��I�}�}ݝ�y�Ɔ�enJ���CO̽��I��K���c��]��Jm���]u�y��\u��t���2�,��n����\��$��󊪣��&��~<����5;���C'�"�|�d�������)��H"���
�gS��Ǉ��Ӆ���a�:�t~�.4��x���,�"�vAj�<��˾�ٚj�1O��~��S�F�W�z�$��;2I�ؘ�󍷗����M�c���8,K��<3��3
<0c��tӧF2�}b�G5��HA�x~�Uw��_V~��*��#�'e2��]f�w,���%�i���Y18�P�����y�՞e!=o�)+�q�u�Ԇ�}�|ŚFK�����%jT�J۔�1�7����y�[1F�R�k��d��}��#nW�֦mRۻ�)�ڇ)"V6潉��jKn�Tm�����|����:e1���N�Iь��!u�%TB�s�W��S�FE��5�,�q4Ҭ����'s՛�GQ�\Z�s�.����
p� ��,���{~�${2���=�~�p;�4Ã=ɁCɅ2	C�����,���d(^Fxj����:�)�T�9U�ϷM6�H��Ƙ|`�Q���4餝���S����eMF��Ey�H��^f&L�L �7k1'dMS����NMt C�{�X���12���7�˘g��Z��A�<�$�*�������͛-p�Ύ�h��?p %q}�iYX��m�sw�d!�U"sh�2�s�\�1�\w�l֪�����c����*�y���=����0�?D��q����>��!���yj�#��`o�~3�y�pNÓ
i�Z��[�g�y�e�8���&��Sٽ��C��vO�W��� �t�}��������h���'&4�Q̶[V���y��N�x	�{�a��ߙ�~]���6È���~q�[x`�#�M:i'F2��!�D2�.��p�oZ�E�}8���2g~��㜩��
�s��h���,0�gP���;mފ"_Js���'�|����û����4�a[��׆%}3�4����rT���'\��b�O�Z1�b�=Y�8�W�EL<�rew'�
x������̹X�~��3̓a�����i��Q��eu�qw�ڻ�=Zwq������ٳ?{
t#���̷1�eM6�y-��~G_>u��G�b>4Ӧ�tc(�� �8I*�Y(a�g���2�)(}���%��Ѵ�V~e��^���0f�I�����3ț1�q�VZmm��g,�%����`�i�U����a���]��%��8a�]a����r�M�|����x��1Y���l�< V�U���@[���5�k����E����;?N���EC�{^J��m�G�U��.�v0�O.��d�d������+�k-��]0E�i��e1��M:i'OON�쾬��ꪢN�ѓ�������^�(��J:39�n�D�:���y�ie��)[�1�n�'�U:�Bv5G�S���O�'S@m�86pTOߘ�|y)�R%�L|��'���k>ܗ|�>v�.���t���W��ɤ9̟0��~��)�����a��r�IS�J��̑�.����%e3Z�.6�>q����2��3M:iӣCŞ�2�����L��JjZ�Y�?k0cəTn�ʞd��Q9��ѱ(($���go+Z�ڣj�V�,r�.5�� �7j�OJ 	-�_kqS�4U���Z~����1�kJp$��9��M��]�]�*�d��)�0�Γ'���\-��)�u<�0�CJH��Z/�V'}�.�"��V~X� ����Q��,.
�=�.e8�9?V/ˋ�\�|�OE��0�]~g�Z�Ѷ�H�y�%�^��L��M�/�N:x�
L�e���'�b{C�a��I����~$�F����L�<0c�4�񦞞��h�"�檪 ����1Q���/�M���i�o���p�|f���=�
�BDW�";�Ƞ���r�D���몓�V�q�|���y��d�r�u��j�C��v���W�eP��؟�`��H����+�G�W�ѫ��]�28}ã�_��Q?p�Nx|/�x�r	"�:��+�*u&�I���C��v=K~^��-]��ϗo�yk�QDx�I�h��	�H�H�FQ������užOi��O8�&���k�k�y��O1\yzy�<�|���'
#E��#Rd14�-�T����iiL#K#Fa6*�DM�����>4�tZi|a����/̱i������+�y����_�[�/��b'�/�y�%�*}Y�bh]҈�'W�ˏ.'�jK�K��yi�O/�/�/	��i�*y�y�'�	�W�œ���ğ���i��t�X�XT%��a�3a&a%��#�ёB�H�H���hZQ$ȴ�ZD�C�#K�4�R���\/��s���|�BE���ēC1D��CP����3$��5�����m�a�#�'L>�8��$�9I��R`�a!�Y��yi�t�:@���Ɍ�YXC��`w��x����Q�����������<�l�'ޥ��;����ﾻ�333wV��y{�����[m������խ��^�ffR<�ͣ�8�8뭴��Qמi񦞞�<UU�t���Wj�4?T]C}z��#�n.\�}L��n��km��S�ǟ���#�>>b&�n�o��Y���^k[���d>�$��&xY<0�Ľ��̯�{��댑պ�Vy�U�}L6}Uşe�U��U���Dš�>d�8��T���#��e���G�~q�\u��1�f�tӣ<2�;�xD)$�C&�{��f/�L���>;�P��5�����k���	nfD�Y�ϙ~i�sϩ�<��M�~|���j1Mf������m>::)�Nѷ�_��w�(|~���y-G�(����D���"ϸhd�vP�i�Z�ݙ���a��?:�-�0�??:��;��N�b��4駆Q��&!E�OE2B���;e�K���
�)Rr��]�7�g,<_�L��f���B�Y����10�X(�;dG�;]�V&�+d�GcR�zL�� �lX�~�Mn��/�,�fY���W�|�*�S�x���]y�\,P�p�r��)�&O�g���ٶ�~��:�FzIQ����a���X���v����Յ����0�\���6��-�]<���k�M�q5Z\[nS�|��Y���R�E����≢"B7�h8���fFL7�^Vq��l�Le=���9���᝕UGi��|��~q�[iӮ��<�̼ӭ�I*�wE�IR
H?���QY�B�(޲2(F2E��# (U@c(
�e!��I�J�"�L`�0�a	Ē�@FH�yq�RH�"ő@�3	x<��UD=~�?�tpD<���'Y}��'e]0���N�pޡ��p�?�I8�z�������r��a����`u�Zϣ]��.YZ5����~]qbUV��.�ۦ!A�^I��e-���㽹jj�qov����&	p�	�mZ'��c��e�=T�z���Ƕ��}/G?c��,c��9!�m�<M���R&�d�韛��F϶mi��@�Z��ll�Ue������k%�JZ�;fc� �6�JX$T� uǁRZ���j`5�Ah� |6��$�����<�)Wf�Ε�ŋ�Ub���.��KjuA�kTb͈Vť���e��[&��;L�9�v��F����j�Kw90	�4Mj��5��Ne�Y�ЉepV�\-YՇ-e�Ʈ��d�Zj��-n>���Js������㎖��<N��K�Y��2�4�L0e1�gƝ4駆Q�LBI-�I$�Ĵ�T�=WX�#&�������!�n�6��Z|a)o�)�HǙh�^\f0@
6(4F�p-qW� �<�G�����\zInSs�8q���5���<`_-87��.3'�ttz}���aA�,��Gb,��� �t�4z�^ޏ�i�m���q�u���3M:i�Oʈ]��B�I$��0�2������m�RݬGpЧ�e}r�����y�S-R���*�hձ:
y:���=��j�_�u�~��~m�����ό:a���#����.�3\m�I^c��5O�W�$�k����[���Y+<�=��L�˛ӕ�4�9�$�x��h������1�N�tєw��z�=��xE|�e���J]�"��5e��X��x��ej�X&o����M��:A��*4�E0��:��Ń=�X����.��  ���+<֭��;6�j�y�X�hy�V�R)kTS��/� jf��Ff�b�s��flT���$��]�M�1QS2e�\m�����_�b\��O�*���N|>^v�j�,�ncsx�ϰ�%n�f��o�m�Ǚy��<�4��9M�Ӯ�w��Mr�~��Y�[Z7�z�e�U���C:��	��c�h�djE�Ҥ+0ݗn!��7��2y?n��ߤ�xh��e�A�3FP��!�Ӧ�4g�Jjb��I$�#�R���U�j�Ҙ���'���T�b�v_��c�!��~�;9شo�[�w6d=��<Ι���3�~�5�~~䇑G1�?)F8۳�e�'8�Z����,UbSś�q��ߔT|�øo���.�L��E����q���|����q�(��!�Ӧ�4g�/��z�RD.�KC�j�2�}'�~�ټ\.RG�\ș&
KG��g~�W=����!�N�v�7ک��x#��§�$-���U�-թ��/����}��҉��&&g�Q�q�-rG,�z�+���~?uKgs��OEi�h�Dy�e��0����'�s{u�3V�r�_[�F��6�Nt��> ���0f2�b����y֜�I$C��5�3i�b�t���3�(�w�#���ਤt���m�G,��q�	G�/|���N��y;GÓ�Gd�=>e٤�`a��	'	^i��k�U�{\��!��t�t:i��Or~0�|X�4�kt��a�f�W[|���.'�?�S
S҉�h��v~3��t�Ɲ҈�Y�t�a���K4f�i���|��'�/h󍱧�i���k�[ˍ<�yq��o1�/���(�ZE�F�EFF��b�d&-0�i�ZFL ����&�I��_�Ǘ�i��g�/ɧ�b޹���XZx������i��Ϳ1�������<��<�=W<�-�0��\���MX�;V�t�O�̧����ѥ�k��y�o�y<��[��<����Ǘ�<�&^�����ҍ����2>��H��>>#�6VB�6����L�5�Dh�2<d-#�Bҥh�Y)J��#at�t]4�<F�
�&�#E�b,�Xϋ���Z����m 1�MИlB�,�7b��_9���k.��ܦ���\��`�!ג̶1�U
�]r�.5�:(��:�-�b�2w�:BDYp1�Uwp�q� f�8bmye/���V}z�{�2��e�%��y�ًL9�*ua �Z�x�Zx�
ˮf6g�#x� �c�o7 �Wn#��4��Y,x�3-�f�h2�""r���;�o�S�o���r�g�דI�I"t��	B��|�����e��)<�����&�Z
p���_I8(�k�f����8G�HF�ڌ�j�X����4� ���Z}�m��X���J�����?L�o�lQ�+�Kkam,�M)�2���lC+࿬�ޕ�6��K�ff1��nE�6e5�1\���
���@5؋�t�	S-�Wd��_
����=�aVG�S�������mf���cT��Z��*� cl.Jb[_�iv,�b��'�K%h#��J�֮�۝��E~�sݟL�����w���_ٙ������˽����[����s33wV�m������<iF�i��3G�1k�Wʯ��u�I�6(y(V(�M
ؒ�9�˶�����!�7Ri��[bh�����)�T���R���w�a���m�X<DѲ�1l*�)����ֶ�CI���3��7�ik�tE��P�5�b�kf2����v�֦���[�u�J���ჶ�B]	��]� ���X%�n���m[US�  ��
�<�:7��;O��#�3$.l�ʦ�fAX���ӊ��x��m���������C����Ir�綻��Sm��NӾ�rd:%��/�e+|�gb��0)�)�~���q�wk�ð�O&v�?Ci|Y؏�����?�N���թ��&�8~��6�'㩦�^S,����r����N<�ߜ~q�u��:�:�̼�δ�I$��}+?	����m��O�~?7Zn�u�[0����<�~�]�u�.绉Ne�5_�Yo�u.�孋�����XF	���me�H�g�~� ��$�_�sž~�'}��~�e��p�V�͇�{E�p�RHb~�'t�M9҃;=cj�-��st��m�?:��^q�t���3N�tћ��2�ĈiUD��{�Ym��B!�X~;~c����!4�{�[a�u��H
~=�L��gt��;��e��h�����3��3a5�`�z���cx�����'�O�W��ߜd�T�Wk�����S�LRi�隹M8}��К���~���c���ۙܮ+���Z]4î��ϖ�����8�m8u�u�y��|srI$EakepH�[%Z�u�b�V)�G��|���%���A�cB�1��0�by裦p� �d�|U����ܩ�w7L�J�.V����:��U�y}<��<����K?X�;c�^1m�g����	��|�Ye\�7�_;R(_%g���=�(��4�Ϗ��4�Q��C'�Ɵ�x��˟1f)ˮ��P1���y��;fƘ��m��u��{SMҁ�u�XIs<i�Pm�d� u�m����hM�rB� $������T�#[y<��c�˳l�s�nd��B�m[�px��N("5���|��}IKi��[������$ϿR݈�2�L}!m��wu���V2��],��7�3Xh�M��O�n�������͆oR�)a�f�4�=�ŧ����Թ�AƲ}$�t� z�����tv3��l���:bfw�-��ݨ�-�i��[����8�m8tb�4Ӧ���t��I$���V�f�|�5U��S˴�C�%[{�L7�4������4��9K�)�fHut���c�~6���!!aJ�?1�L�૕�W�k�fۮc���LE8u��a���SώIÆ��ي��"�']�����E{��$F���J��x�Q}�*Dm�mź����8�m8u�u�y��s)*G�i"7$�D#�:�5�n�����y��}L2�c�����ڊǳ�P�p�M,K0:�?^&9�L:�1͸a��,�s#���D�����SC�B��7|cJ�t��ϼ&xrA�1��Cn~��0S����;��SJe��w�Q��J�Xex�4���ڵu���#���b{
�i�R��Rm�wĘw�[F3X�ڦ4���eo��o6��FA��4�Q��C&�t�ӽ�t������%�/���~����4��J:2P�*�æ�L��]��������éaa��cM?~[(�z��^~�_�S�8���]�!���f��=���#O۴��Z����[z>�'�\��F���SC(�p���������<Nw�>{;\|�	�<"(�� c4f�`�<`1�c$�N�3;Ղ���y��3F�ZK7,Ć�+�@��T�kX��ʧ~�zt�� w�ܘf�0P�U#��B [�\�,q��H��'��=� %�����N6" d�N܆dȰ��(��X�]�(h޽������eĻű8V���M�Ն�����q~e�]˵�P��?|����3�����(��P`w8l��t�a�ȉ��M(u�2�j����醈b�~d�:��V��������e���16�\r�>a���8iCD�=��?7�r">#�p��e�x��4њc��Ӈ]G]aיy�5I�$�"����XZ��5k<�0�"]��/��^C�C��ف������Hm	�b�?S8)��b
v�駇���M��ykO�7��k�]�͈l �}]Y�J�G�[���.x���,=CfL��I�LFp�Jd!N��Om���zl���,/���2Fߑ����x뎭�tc<2�YC,c0f32�P��çF!�$�"iq��bF3���3�0fH��<Y�3�FX�c(e:0��1gGI1����@���C#ьc cd�44�!<y�"0x�n��ɔuc c�c0bB0`�2�ў<3��0�F3Fi�Qg�Ic0f3Y�Fa%���,��Fc<`�xc,��1�Q��y�pȸ2_����N'�W��9X�mu��6���0��'}n��2?���Nch�<��8�|8��kS�w9�r�������`�oS��3�37���ub�{�\��MU���s"���2��������y�������o2�s3���m�˽�Θxҍ,��4�Q��C#4�?i�$�B�\�K�ɘ��>?SoS��;���Y���f�O7����r'��a0��)A�>��r2:<�-�hMO)�8��3����1�ii�یSŘ!����<���Hq;6�����Ϯ$�o�X�FKa��C��|S������%E,ﮗÆ����3>4��A��4�Q��C#4�6�d�����HA�Bʍ�
b!G�����<A����T4>����w����e�&e�%��/���5���C�crwT��3����n7M��<�!�j9O�]I���(����7ؔxJ�����ϸ`I5O��U�3�?;$~���E�u��a���e�i�'ƌ�G�1d�Ӧ�^�f��*%LlԚ���W���6Az�y���������d��[�3q�w1�8Rw;ze�Z�Z+��Y4��J�L��6QWc����+ :>GYW0�+3":�� JL�������򭵊'yH��ƺ�m3��6]%�פ�`���ʖ<�S���OY���3�����^DG��B�(6��a�jI�����$n}#�t�Bp;�~�`�����c�㙆e��C���]�gi��n����u������/���Yc���6bm���g�[_�s㳓��cD��:�ɱŶ�.8���q�_�G�1d�Ӧ��3��UTB�I��|y8����|�ϑ��X%��sR$s�v����C�!Ƶn�3����´%O4�k`��97�¨ E5�N�Xz񝛝�[B��������P�'�ut��t�Ec������+j,p�Y��:���8xtD,��	����yU*��E]B�êuнC�Dgp�x'խ���6�r�{�֑�E�M.�Q��#�#�%sD|��3Fi'��4�Q��1d�Ӧ��;��1al_n��ǘs1犫:���y=� ��	;;�Iw��۞$��YZ��>.���x"d,JtCMTW�!|���݂��������I�巳`���_��h|d�B!��a����(}�?"���[��v��]�?7M�o�JkH�C��;�p�G��8p���~�
W9d0��Ěh�0��x��C#4�.��I$��xEؼB\Af[uD5zEƩ������խc�˞�4l,U#h%�O���B�N�i��~�����n���8���|a���~2~�4�Xi�o�fغu���>�/s3+���skM#����!�P��3M�D�B��vwZ���FjYaeƞq�~y�t��0dd�Ӧ�܅؊�2(��^ډ�m%֮��_��>�G<x�p�(<���"A� ���g����w�uy�����"��2ݝc�1ql�� !=�Ϸ��s
K2 ̮,*��Z��ZWr���_k�eٛ��<�Kᇑ������|E�F94�ө�e;)���(�$�M�rq4b!���,���mq"�f_���"gRM���MUמ��}L��r�oZi\N0�M>ܙq�L:�	8��~��I���~����?����x�"�{(��2γ�ۆЮ���۬��֚9�����"'0>�#e
X�Q�L<X�,���i���0dd�Ӧ��qq�J"<�x�"c�o�wT�h�Q�ɺv�H��+T���Lr��HL>�w0�x��牑?t=Jt&�W��*n�Z�[E���挾��e�>i�@�QO�jx��!������ò�C���f.tt{��k��-�[��b��0~��m��y��ԥ
&x'c=��,�fc4馚a��xf����tюx�g���ݏj�Ģ¢���(φZK��f�b7�x��d��� D��s�^φY� F���.��}θr�����ty
"t_z�RўV
UX��e�2ʞU��-]�CD�n~>8#�rH~H�g������u�
%/�+z,��p}[|�>k4���w2[(�M0�y�<x��i�M4�,��#$����̗UV"l����N�m�S�Pi����vTL�<"K��==����k֗�j�j����:�4�ykG)�u��"F_DW��=��:�}O�ʜ1>�����x���3��/�(����o�A�	���q-���7ӗ�ҿ����}[�;Ke�4�Uԑ���[�ţ��<u�V��m�Zu�J(e�f��`�I%�2�2�K��u�a:iӮ���묺2�xc f��tc0gK�$�e���2��ф�c��1�(��$"1�c$c:1��]u��:aӫGV��:�&YDd���#ǘGV��u�]l�1�<!�c f�F2�3L4ь�M4�K,b(��3��aјIc<3(�у�H�b��Y��1�Q�G�t��;��	F\J,��.H�ߦf��t"�d��:f=@�Y�m3��#�]�eYUP�T4&���D�Cc��6���ˉ���G��K�eMeI��ʛ�_\�u��b+���۸�p�4�f��WnI퐛S�����@�Y5��a�%��)]�90�D�!h��W��	��ۚi��.�U��D�q֌���V8�����KU���_!L�P�� �fZ�4[H�tMq�f�G��*�Nc��sU��O`��h��m��=��1��UH�6EUĳ32�E�S�hK�دj�d����5��fR�k���5�]It�R�R�������v�v%,K�[�F�`{r,�bX=�4Q�^��nf��G*`��Gj�4h�])�cVf��M�}Z����r������Ȥ��;[^҄�cn�}�K��7z��)�^7���ff��ζ�f^�fn���m�e�ff��ζ�f^�f4��,�Ft�M0�K<3@�H�4џ$a�~}�ʸiei�ՙf��!h�s���`�iK�]^%�0�����9�\���R�:�ٌ�B\�V���F5PmʛL�[b��֒�W�!����37].�h��L�mt���±�HJ�VR̋m�2��͜�,���k��ʨ�0��p��&G��շK�)�pbW������	�f�~F�+� RU�]-��0U�퐂q�5�Y�b�H�uG�6+��|��<s��h�x��6�Ild�����)�HB�?C��|���!qp�ǵ�Q9)o�##����ei?.&iĦZa����9�k�$��E�R��~�X-u�W������ۦj���-[nrMS�0����.���������(\t�a�њ*xy�N��6u�n%㤒x��L��M��3A�q��q�s$�TGj�u2��>=����dvrN���4���F�Xa����.�ߛ�4��0���b���ӡ<�'F�iD�����$q@h���<O1�~���=��)�=������J��%>j�???S�����l�M5\i+[.������h�4��2a&h�>�B�>�Ub%���)��O3.L����v���l�?Rب�^��b^=O��iƘGt�v���S�S��[��+���L��T;�("�JeD�d�D�ᄐ"��������c�����ԋF�u���\Zv�����~I�-ؤ�����?%9�-��&M~)��;?X�4gO�4fX�0�	0����8�S{��;UX���;��Q�[��E�,:�=[q%:������f����Oz�2��f��ʏJ]喈�$�#>����I�@��S!�z~��Ju���',��mimr�JWK��~)�l:�:O'�č�����(C��BGyT-��e�y�5V[�;_3�-����Z|2�0����>4јic0c$�WU]_.�kY� j��"c��j�-� ﲟ�@�|#�	1l����+R�QE
GǞNK	�/ĉ
:�V��6�ئ4�<rU!��T��s�����bZX�M�+*����J�HX	x5��tn��C����9����-�|�=���be�t��x���'ᇦ�������i����u9�D��V��[Y�&��K��*����>؏�¾�����&{٘�ē�b�ZtE�=���~��Л���U�v]�%.ʴ[1�]��oŴ����o=i�ԎWΨ���Fi�M4fX��0��i�ڻ��d�I%�!qr�"�-�xo��m�O��+4�#�ߩ�k?Wԇ
#$��k���5�,>)��R�?s�"J�	��#�)����։�M4��$�:Z�j�	i[J�Y� �A�_{"R�JG�ϻ'*��Ke��(_7Wk����Q�>$ь��Oh�4��1�a&x|xu�*�D���,�*���ٔ[�5X�������"?;�]�!�a~��7"�/���F{#�7����&����µ�F�5�Dc���铇��}�<��A>���G�0���r�[;��-�q�H�.��1?9P�YX���K�W�1e��eb��Q1.�#�J�-ʭ!����Ǩ�_��,���2`�)k������	kpK@��ťF/��^=�3����T#���I�o�]����l�O]RU[H<�R�J�P��T6�6���vs�5Nq�V��i���Z��2&֘�r<Tl=5Օ��Iˡ\�J�v��uO6�W5��x��%'��.=��&q�j�]0�km��������{�=�vʊ,,eUP�*ݻ(�!�׶���3]i�	�rR)\h���L��&//��hN(L������c�0��1�7 yc�6�.m�?�=�c�[�l����5�|²�@�6V���3��wfl�a��'��T�6��5#3�^�K����7(�%|Z?b�O�?a�m����8�1�4������e��R�|���uǚy�q�θ�8Ì���ĩ�RT�"@X�
��)��a�/I%@b@�(2����,A$�`���H`�$�Y!��T$E5�a�Rc!Y@P"��((E��A�ERH~�@�I�x�������Q�Q�a�����1;<T�'2~�po拜mn�i��Ƞ�9��ήp:�$��vzyҲڵKkI��FzŔ���i�~�.��N�2���M;:�N���{)D�u��gCO-[I؉�_����uG�׳N��u.[����Τ��G��:�o�|��<��<fX��0��i�k^.��(��ڃ%�-�8'W���⫱�΁�̚(ڈ�LR2��t5�2���:��ͽ���k`~*�Ds�[���[ļ̶��N`�O�[ŚDMhq7$��MW�e���FLu9�K&�Dm2���n]�6*����v�y0����Gm��-a�)��њ��~~;�������{�3aɅ0����t��G�kt�i��V�=_�*O>7_?c�F��5�aR�đ�OVօ�?x��~�4��h"�#C�<��_"#�^��<����͸ێ?4i���K�&a�4�Q�G��$��<��[`�<�.>F9�f�Sf�쟺X�Y(���B�_��_���RD�T�\[�C��#.�OR0�p�:�U}qii����(��&Q���転�����L�S���j+���tQ?h��S&�}��%�������`ü�[�^FXa����G]G0c0��҆X�`�3�,��!�2L��d� C�b�F3�C*Rd��PΌf�c0e�c,��)�GFH�IX�1����:2I0c�H�tc�`�(��t�Νa�e�FOy_��0����1�1�`�`���#:0c(c,f�h�4�Fi��"��0��f�3����0c�ј3��X�1�z��*�$?�Hb T�7�O��'HjOoT�O0X��k	�=a���I
ȡ�`IƪA��7h(
E&2�+S��@������|�!1R('�SR^�\�-:�a�W�3�	��8�1 ,�d��%�Y
����& z�XE��%C�A�q�I�8�1��$��h2h�%Ϸ����.o%/}Y��W�g���z�2�s3www���̽̃7ww{��32�37ww{������<iF�Y���3,fd�I�L,�9��Iq�z����qD�9��tΰ����w�>�ȏ�����f���q�g���M�iZ�_/W����o��|��]>_5.�	�Ͱ��-����=D���h�t0��	W�nH'蒸_1��Qqy,#����˕v��8ӎ?<�����32L$æi|BI$$%x#檬Dp����S�P;7y����[�����~�!�{��`�����m���q�qؔ����z�|�<��ח%���u�FXs޽��0�'^[N">�SlG��>���L���;�SLV��>e��h��ND�������Kk>F�����i��M4fX��0��v|d=�[��ۈ�J��nSq��gm�;q:d��� �El��m����lBZ�9>MSb�a���,�,��iG��G����)闅�l���3)��� p���oK�g�n3�KNY]��c��!�����"�����f:��<�M�'G0�������r�çȋn�V^g�6��)�!�ߥ��a���32���������a�	��xg>�̷=���b'�<<:�}|e~��6�Dͺm�r�X��x�.�%8�����ݻ�	��+��H�i6�l���^y��3,e�d�I�L,�Œ�Iq�2Æ���uG��ƥQ�߄�V�����;�H�|�5�[����~q+�[�	Qo^\8ӊ��vt���v�Q�C�c���tXyX�x�|y$���Vm�m�<���R��>]7������HG�q��B������׆\�T�*u�U���j|����ne�V�mz��O2�>���%Wݧ��q��u:�/�|]'�|;<"=�ϭ.Q����F|3�M(�Fa�����	0酚V�1Ub&�`��w�ê���K��?u=�q�S��aߌEAg!�D;��~�[*~�sa�v"y�s����p�[B�k��S����O�ϩ�ˬ2���|��˻��z�v�Z���9/�����!	��iaGxj���H�����S)M)6�4�0��F�,��M4�M��2�2L$æi��]�����,��~K��ˌ��z��ʫ�R�F�C�Sȣ���]�MԒ9�lK�0���҉����(�]�Y��ǥ�Dr���m�eo���a��<���}��-ߩ#�j���F[n���a����mך�km%V����p��h�_nD������(�ΔP��јic,c$d�t��*��b!Ҥ��&{13)R�9<�^<��g�b�U5b��h��P^Gǲ�R�,-Zj����9��4�#q7#q�KpZKn�_>�͆�6��O!���%a	�@�
�,����c���I����L&y��6�T�1k��c��ӱXʝ*���T\Z���T�0�t��/�Ώ����.�h�[H�I�{�6�#���<~䟩��<�H�ֈi�ٺs����������d�D�n�y��9�9��cʯ�������[	��5T��Z>��ۦ��_�2��m�i���|P���2�2FI�L/��"3RI.!�<"�3�xFUz���k���Ȼ��>f����%��?{�����B�~8pO;�����%mb��-�b�uh�s{��[r�����g�`�F:¶�[3.��mL�m��v��qݷ=�a��N�ON:�OD�%ZH����"� ��AD�ٺ���'�~����[Tӆ�p�şx�4���3,e�d���Yz�IqgO�z����g��.y�h�X]ar�W����u�R#�[5���j]#M�N2��7='�HU��CX��#�Zj�m�[�hp<;Tf�0N�{�丟��v��8����ب�O��e�.��q��Kw�;�4�?S�b�4�Ry6a+�O��W��}_6��m4ن3Fa������a�"�Gr�S>UX���Q��'��Cñ`�*��Q=���=���뉭�de��BpE��+mnJ�{��4�<���t;�_��;�ӣa`��a�2a�r�Rii#5��^��DW��_̦R�az[H���6�(�5n�mi��][�0���U�[�v��Ÿy�el?0���պ�_0�]i�(d�1�36�f��(�P�ш��N�!�4����H�tc(c,:3aь��%���3Ō��Yc(��P�1�e3t��$���1d�c<1�f�,`��0`�<�(��=^���<�yn��]1���c��1�2Ftc����3M4њaf���`�<3Xδ�E��c,�Č�2Fu��0�+�,�9��׳�6�<�2?1\���dqXH�'2�*�-��0Y"�jq��"��v�KP|u�K�n�*s�!O,H�rȟ3;uZ�f5���>,�xғt3����K�.cKkUi�˫g�?�64�N���CT�7��L<�#Ǒg"�dyY�q���Y�Eg&F����`��kuD���=�<��i��gGlBղ�c1�:� �6FU"��f��fͼ��Kr�әg5�؀6xUkJ���l�g���A���2b�VWk?O�h|c,E�~��lO�U[�ȕ�W�!�k�Yu�\�ƛ�mv��V5��!1{�`�l�㛑�6�6��s�-�l�f�j:Zd`j�ͮh9X;�������>�{v5�SX�m3NF���2˵�\��D�<�O}
	쟪�}~ۮ�ͻ��˽7ww{�������������������k�����A�x�M�јic,c$�E�WW���Sj[��$���.�m�F\�%�t6�%?V\����4վ�R��ڣsp[.�U����ea\���UƢMpL�%΋6�b��GK�����n�u�b����Ŭ&�B�t� bѬ��.�*9u��-��k�m�e���f���*-�|ˆX�\�ڸ����]3Y�U�f�J��j[�5(jٍ��$�T��I��<��I�D'K�Zr߿ �������7�� o42
�2?�F��,���`Y�L�{4V��l�'�tn��f(��NZQ�8/|^�<L6S'����))ò�Ύ��i6�;�>��У�!p��	���R�!iE��#�p����㲉���`nIF}��dC��>"�5$.��o��,�x�1b2��������Y��1�uţnT�Ǻ�mڲ�(��||i�ь��X�H�<4��^ݿ*�DO!��狂|v`��J 4��X�B/|i�q��x`�y�J��&!U?iN�O�2_�S�2s�}��	K;0�]��~��U��ƕ3��p�Ls]��sv`��t>N�Dg��}3�i�dJΈd�+��e�!�	G��Q��<3�,��4��h�if�1�2L:ae�ũ$���4���NS�������KD��^h�����]9�D�va��0G���k�'4��q(�5�k.�ѱ���3Z��8d���'��>αp��K;�4D���'�ua�,O�D�l���8��ۘύ8Sx��&���5�i���]��G_f���j�4��:2�4҆h�if�1�2L:ad�u9^�kX�<�Ng�*�D�㇧C!$:,|ҹ�0��Z�&g����q^ �U}�4o	�S$YeR@��J,G�+�,�����#�2w�����}ñ4��Q"��~��=�����s}�;�Y)ʋ[�>����Y�Oy$�>a�?~�_p���l����7NMs��0N�ϿLn��zv`�D�cc4�ì-�sD�>����ǩF��SM>q��|�6�Ι��X�H�0酝~��)�:�����i�}����I�z1ĬAh�~V��D�Y��s(�t��#ς�kLd6�f���I�V��&Л��qX��w�-g9� x![1l{i�S7 �ԉ²T��L7w�MےLwJ�nW`V��2�eݸn�[Z�E�%,]���=>�}>�Iт!�SzT�����ܘ#'�	�g����Qˋ�����Z�n��ϼ�u�ю�ᥞ�=�O��
z`~NwC
%�ف�����K��	�����1����`��1)^X\�Knۮ׺�2�#�֕�m�nrM��ie�f�3F3K4����az� 6/V�k���> y�ԏTD��4�T�����#Y�˔l<�m�y��O
Q,;<ؿ�Ouz4Bu,�1j6�x>;҂0��!�)���Q;��>}��p�Y�H��b ����)Zj/TiLz��%"6cO^�l[���='ϰf�?8��B\�Xe�q�a��P��,��#$�8v�)TL�Ub'!���s��v{L��!�[�O$C<L��m�q�"��>n�v��c(�D���yT�B�X��j�,�ٝ4�]%e��dm>�ml[�u�iGÇr`�"��t,�q��ɶ��i���8�+7�b�x�웳ɉ�k�B7U�Q�y�<a���4M:�z���x���3�E�ߑ�����̅��Qf���:|P�4��3F3K4�N��8���I�p���I$��k�ܟ>�4,�B��`�}:���cT�G�m�Ά&��u�����_�/���
:n���#� �3+���,_Y��߾{mH����S�Q�C�]K~Z�Ѻ~��ԋ�:��G)�S_Ivj�ah��K��1R�eż�M>y�μۯ:饚Y�$d�a���L�*faz\�v�:�b|�G:�儾�����_v�WāM-hzhݝ������$.�
�9�mi��z5�F��| W��z��LM���o,��Q}��1�9��DY�j��jk"~<���s02	;����{7<�kv����>�џL�>0�6����}-�DN�F�
za�wݭ-[�}��V{,ONCN�4�tV('T��˂��á/웥��4���Xd�k�h��s�_U�R9\~�J�O��t�cj`"Ըۆ+cE�:X�=2Q�N�?1�p��$�Fa�E�if�P��,��#$�e��I*�I%�!���X4�a����,:�g,�֖��S�e�4��i�BV-�ڵ�],���S�m�:>Vi�h��<G�]�%�E}~��߽�(�M���qH�N�1>-Sl+��B��l�������'���[�_���bv"�5L>�a�Ն�8�ܺ������]6˴��ah��<�##+@�D���3�0�3`���,��(d�2te�$�Ӣ0c�$d�1����RL�2�Y+�,e2�YE���0��1���d���I0c�H�`��`�GN�uYӧY<�(����C�1�3I1�c$d�tcD�e��ƌ�M4f�Y�(��3��2�P�%��G��1���xe�0�����mBpB���g�ꬶ�럟T��Nx8����<���}�ّ1D���?�s۷ww[{�����wwu������wwwU�����ݻ�����Q��iC4��1�Y��2FI����w��O���a��7�w���>�;��̅F���4�6�-�ֺC�-�sk{,$f�++��IX(V���Q�r�Ku�Z%>�gR"�m��G�u�o;���b��d��#��仧�i���0�v�ܦ�}�,�:�����.s�P��}�Q������F3L4�N��8���I$��i����I�?y��=��'��SF�Ɔ�s��U3d|b�y�F�7!?��˛����Zu�r	��øiF�3'��~��]n�LUa�%�z�IYj��7^�y�Z{��;o���8�e��{��O�F��xy0J(�%���&�E���˦[i��a�Z3�Y�,ь��h�&x���WӘ�@ܳ�b���#����Bz4����G���3g��O���獷cے������CM���UE�&e�*O
�ZA$j�]�T��F���-��� !	f8(,��"1��,�`�x��`�m��xm�	��s̐u�2�l[�Ct��P�#��`X��u��D�������欞(�����s'}'�6�j��V����"�i�i�0�'y�	�!�G�I4�]aW%z�6�i�G���PNC�䡓US�M���������3��Y�]ք	���]7WQE�`�a#�S�V��,�Y�,ь�M(ђ2L0񇳱>UX2&H�����4�N�}��M�0N%"~�d�|f���ڭ��L]%8v�����]t�B������$ܤ�S��N�ܚ�XBEBq:�_j�B=�H<�&3s?m9���"�eb���k��S���;=>��'!�F
�b�C��JB#�F�H�,����g��7j�Y��n֦��a����d2�v��qd��y��}�4�'OV�%1�a�I�VҞ�7N0t��`�,іh�Y��h�&<?~UX&P�Þ�n��aOV1&":۴�Ԕf��ʴ�9*�S)��o�Z_3\��p[8��n��vy:0�iȆA��K�/�ۻ���F#םs&�#�N��4���}���U�~��ڑz!�΁�Vi��!Å0袆i��2��4ҍ#$�Γ��~U�'p�{3G�Tˈi�Vb����[ŭ��4���K+݆�k��{�r��kz��0���y�57���˚�����0~�V�~e�4��EW��^�LO�m���},�zi	F�}����_'��K&��qۗ.oQ'5_c������:���,��`�4c,�J4�FI��}_��e��pRG�ט^�GȉE�e}j����帅1<kE	mśnk�F�,�BfڅMf�+�8�]6)5��� 	
n�5��Eh>���m_	$%tC,����n���!��ጌq+�|����E�]�9��3>��KG��}N-�#űXcˬF��g'b`��#;�~}V�����"�\��xt�𠄽Δ;�\�\ȑd�S�d���w����m�
ˎ:@�\h+��t�մ���]���*����6�����Z|�����Y�0�M(�I&xü�̈́����#u�˙OᇫJ��adfC�{��XN1C������l�J�ɑ���rvl��N���gge=�_�~�d�t��;K{j���[m��G����='���pϴ���F�ɇ��囫]zئ����>�wsYf�V�N:Ì���:�x�,�J4�FI�0f.l.r9�gCƫ�V�+
�a�igqI�Y�?a����מ'\��{?B�	�������\2���{K���z�cu�Mz��̩S���s���0�`�����m���xW�a�ފ�/��'�t�y賩��Y��ɣ==6��1�u����?Sl��u��8���Y�0�M(�I&x�-�2�V�z�b���5S�`�mr��h�LA�#1R����(Q�#7R>~��S�[U�Ӵ��6z�b�\���ϩ��1�O��Xa�v�S��B�ҏ�?N���2f!�*eJ%
#ܒOsC��{�ܓ
?O� ���rI$�$dd	I���4Q�y�)�W�����#�M_X�,G0���Q�
�PA�_���L���ٓ4�� �
Bj�b�JB �B�	H"��rHD	HB�RP��!�P�BRP�%!	HT�T �A��b!�1A,eF!�J!�BR	HT�!	HB��J�B�Q��	P�B��J�D% �%BR�D1
]B ��B!*�)�T"H"�D% �J��P!�D% �%B A�T"	P��D%!�A�A�ȃ!�`��`�D`� ��"A��DdDF$�IH�`� ��A#�� �H��Ȉ"#A �ȉ� ��" �b$FA"Ȉȉ�H ����Db �DdD����"#"$H1D��D��D�" �b2�D"0DdDA �D��"Ȁ�
�QȃD`�$" �`�D�2 Ȍ��D`���D�"" ��2#Db �"AQ""0B""1� �""0H�""A�EB)������!
dA��1#dH �"1F"Ȉ�A�#D@H"1DFDA"�D���$F�AdD��A" �"A�$DF�0D���H0D��DD�#d�A"0DD�#" ��Q$�%#F���� �D�DdD�$FDA��A�$A�$FDDA"A� �F�"DD�A"2 �"D`$F�DH"##" �F$�"� �#DH ��F�F"#A"#A@,DF���! �1#D�DA""#b0H""0DF��$D�D�H�A#����D�D�$F��	"""F��`���D� �H�$"�Ȉ���%� �D`�#"�H�#dDD�ȐH�`�� �# �2""#D`""#���"""A Ȉ�����2$� Ȉ�DFD�DDb""0DFDD�#H�#""0DF	DE���"1Dd�0DD��ȉ�"A`����D�����D`�"#"$F""ȐDDD`�"�B0DFDb" ��DA���ȄDDDb0ADD#" �"0b$FD��H�H#" ��#DH���0D"0B��"0D�Ȉ�� �	��Ȉ#"Db $?�aDdD�F�"A�" ����"DdH" �" �" ��H����" "1$���Hi��!G>6��B�!J��P��BR�	CT�Ј\HBud ���%!���BT"��"��%B���%B!)�T.�% "#�	PA �0H�!*�]B!)�BR	HO��+BT"	P�B��]B�� �A�P�"�2 �� ��6�XT�H��HD!	UB�]!J �P���!B�kPH�"� Ȃ �A!R�	HD"���	HD��P�JB�BRBR��!	P�TT%!%!�A��D*!)�BUB �2 �0B" Ȃ ���BB�	P�D%T"���stiHD%B!��B!)	
�JB�"	HD"�Q��!BT"��B(�!�JBR��"HD��	HD*T!BUBJB�A�P�%T!	D"`� � �"	dA$% �A
�BR�T%D �@`�H�ABR	HD�%Qd%C+��RBR�TA)�T"	HD*R�R�D�"	PD% �D*T"��"P�A ȄH�" �!EBRP�*ABT!BRP��B�	U�T%!D%T!�JBUB*��!	HD!	P��B��*�� ȅ���1H�R�D% �"�B��JB�JB�B!JB���!	U�!�B!R��D%!�JB!��JB!)A)�JATBR�!	H"�"	HJ�JAJB�	H!��HT ��BUBR����z�U� ����BT!U@��B*�JB!�J�AR ��� ���B	H�BT"��A)�����JBR��A)�T!	U!*BRB!*�	P�"�%T!��b�H���1 �D"�*TB!*�B�	HD%!(�� ��TA�� �"� �0A!R�EBUB!(�!!	P��J�!��!)BR���D"��J@DD �B1�A�$%!�%!��B� �A�A� �#HA�A�0AdARJ�D%!*����%!R��%!JB$A����2 Ȃ2 � ȄAAD ȂD` ��D�0A"`��A#H�A �"�"� �2 ���T�B�	PB	HD*!*��" EM �#��|`�f�S&�	{�H�Bg�vǝ��F(��HH�*1�_ &��&�ƾܰ�c�O���6��[�T��Z��0
:����ظ�/3��r��sI{k��Ѡd	�y��L4�J�+]�X$���j��"�Ģ� �|`O����.��)v�������QGޮ��55���^�����S�Q�sW��"�?��b��ӊ<��x	��#��~��~�bP��/��6� ��Os��^�!�!ܪub}�"�08����,���b�L��"X{p�G�>���P.I"�[0��_��II�&/��*�l�[Ŏ99��e��E�^ aF��気��/cbHD<Gᓛ���(��Ġ ����6�@
Dn" ���p��"UP"�DP�P�PB������I��Ӕ �6�伸�Mz)���`�:�AU.P���R��U%Q ��$�@�T-(HI�!e�zb�r��'�a��F$z\qN@�@�7@3�b�x0(����{�x�=�S��;��O7  �TQF��i�`w�u|��/�	G�x�Ā}:�W ����^��D:���3 :W�5'�L�G�)�&Շ�>p�������b|��z�Ew!�b�5��,���W�9ԛ�tL�E��9�V��nR�
�H���"�?rs��F+�����^�I-e<M���(6���%`h�S�aH* �ލp$��I4Ē�땃�6t�"�@��C� 7���:p�D�/����%!@����jކ84BA�m���(޶`�1$�B{G$ED���B��t'.*�̢(��-�^��H�@��p��ԩ�?c���z	��`]�`m�+`@�M�&�C֜�x����$�y�����{��gj:p���Ҕ5�>E`D������QQ�X�Jr�����a��7��ڻ�r��u����!��܀2I�&B�!!���e�7�Xa!	!qAB��h�7=��)rE:�� wf�E X3nvw�d�}x�:ļl��m5g�\LTE`�	�p&na
���p;G�(lpj ����r��kL��RA�@O�p.�Z����$f�7�R(��>`�u�`7��� ���1Srk3Qr��(4�����a��)':c�������$�<�AH�jm�ݟ�]��BAs�w`