BZh91AY&SY�d^��ߔpy����߰����  a=h       P  �  o�t 
�              � ��D�$ 1�@��     >�� h � p� .��w=n�M=�ws7Cѯ����}�;��dk�5mE�غ�/�$��!ʋcv�@#` ����S��*=�W�S�卢��z-�:�j���Um�.���=���{�;������Fk3<`�v�p�ۻK����h���k���ݙ�/+*%��  ��޺]k�@��-�s��mu�������m�� �#�+A��r����쮮��8��]n�F��N�F0  a�����k{�s�n�t�uf��.����&�Mp{{��Mک����8{�����ۡ� 8 =3�� {�������m����<{�v^�a�b��8.�E�#����Np0V�.���;vӸ�]:�Ƕ��                    �
M�4�%S�3ԩU 0  CLM0  ���B��M4 F&� i����<�T	T   �4�  �H!)R��hd4�4 ��MSU"d�4�h���LM	�zm#��h�iL2�� �)�����I�40�� 14a�z�+�-[�\�Toc�߸�;���ލ��f�SNo>�O���f鍘�z��f��/�?"���clپY�H]�������MS��p8Cl�0#`ߑ�3f�3���s�8���nm�f�ܶn��L�UUU6u��l0�lv��~y��������ݽ�w������xv�����t�����O|����0�.���&8(�$	ߓ�A$z#�	�gL:�b�,��GI#��RH0I'*c�1��p�yv]���z]��8��֔L������'N�#̘����3&�L\3[M�QLI�F�c�ra8'G.a,�� �C�va(N�b�?�|>���8p��nc��v�b���e��$~��"9ل�g}�|��`���8X�x���L&&%���1"@��a��L$�'k&3���1%�@�D'G�0�.LYB\3x�����F(��x�"�B3鎉W0���3Y⭘�!�31"%�f�L8>�S<�bp̩��Γ#�E�\�q}a"$ag������j�1d��Y2p�����D�E���p��)#�	�$�'�~�� y5�'\%L:Wx�Y'm&�I8K�?I�G�>��O\�$�8�c���|Ǧf,N�1,G�Ғ�=��Œw���	�HD�3Ig�"d3	�=Ě<�X�^$���b��&r��Ygb8"A��D�
"�S���
*#��Q�>��"�"I���C1�53�$K b�(L�9�c�b0��&�Ȅj1ɏ�UF#�L"5	�8�H�$s�	g��cS0����G�rc�\�H�K(y�(�����>DF�a��ơ�����'���GЖ"v�B"�I:1لDf<tGЈ�,�����1d	�BH�va�J0H r(��8L���$��L�L�g9O@�,'�3"r�s"d�˘�bY\	�<t�<�JP�aD>��(��D��(��ba�bQ,���&b|IC�D�r%0N�@�:5Q? ��d�ߟ����BtN���xǱ4X�=Ȟ'�X�0��+����"Q8&D'��' A�OT}g�b!<X���������A���% D�D��z�Ȉ�tD�12"3��'9�)�K�H<KQ2"%=��TO�p��P��N	�x�����	�����_?E�&�B'D��)����K(ȟ��$��5	%�剑0E�O��Q}I�dO�s��>$�)�JtD�IJI��(g�)�أOiޚi�'��g�P�"s���	g�����IV'�~���y�'\�D�F	c|��\�fZ���fG�0��4#F	����O&$~��9�A�za�ň�Dؓg�/��A�f�D� �F}�90�r��x�
p�Fg�r��b*����"#���'�f����fj:%=��G��-b|a�ߡ0E�N���I������~A���ȱ$���|�53�1�?3=�S�Y������C�����ܺ�*(G�ÂtN����3Ӥ���H�	�<�g�&�6x����:u��O�%�D������8[H����-�K�"5�c ~D��Q0X�K~� f�	��(��0r�l��}��<H��'���6Q�Ģ&v:O��?Br"���"�J�&DKj%�`��OD�
���CȔ��Dr
�35	�+�OJ��
�����)bl��(D���2�`����bh�BR��@���G���뉂�#�FzbS�"Q�>ȟ���0�{��H���fl���B&	����II(K��	��Bp�(��L��!Ӑ_�$�$�DP��D"YbBx��DIn%���0L.���bIL��0��)�)�\��`��t��	�1:Q��8�tN�1�v ��q�D٘�$$�x�za<"��pL���	�U3&J'�Ä	GD�:u���'q&OH���f8aǓ&T̉ڸ��$����&?F	�<,e��}�>�VQ�;��?&�`���14p�fxQ6DH��g��8��	+3S��gP�67��V,1yg���K�4$�3&�"A%��^L�B�	8�/��"���B@ϦR�#�D���p;�6�g���ד��Vq�eoɣ�K�!{�(���n�T\SH"'�(�.�:"H�Y"�&��fDnb|"a}�$J�L���'.,���!<{������>�8�)�����~~r%(~�����DG�#��"za�"#�'�蘞�"y��K`�?<�Dn9�DÌY#GH�",t��Љ���'!$��L85��J&?G=0�T�%�D�	�"lKȟxx��NK��N}�$��?BtN��Kb�qbpN}	���'�x��DH�3�}�H�A��N�D��!��f0E�$����<5��0K���#p�s'��#����7�d�;��>�پ3ө����Օ�T�d�3��ugV�*�a�Y쮴N��?%���R�X��">���Ʉ��DG�,H�8s�N���10��0s"<A��B	��ýb:I!��0Ba8I_��
<��D�Ã�Ό�G�'�
8���L��&��=����Q?*��b������i��ǎ�vK;E�'�ĝ�:�X���F�}�	��N�+�b���n$E�Ş8'�:t�BpL�-":8zb8��1ҸP>��.�྘�fM�ab{�����|L�(J~I|�Q,3َs�(f8%	�t[����Ö�pI(J!�2%H$�B�(Z'�@�Q2%����;�Z��O0�i���:P�C�d�'��$J��8IF}1'D�Y>,N�d�D����`��'N���ML���H�~D��&����tb�̘�KY��3_��;l��p�vbfYTNy�����^�g��/*�����ad�{�I=Ԕ���)Bs�����)������M$|���{�t���|���d,�+�ۤ?��'�H��_3wh�M��Hh�Ӷ�gy9V�.rhﯱ���4��]��mn��!���t�ӏ�!Æ,~]t×Қ<x�4��݁�����<z��ǈiC���;~U99�X3�ɧJ4���x�>�^Jx���9� �g���NU�~����!���Y�2���q�d��C�!9�CO���k�͚��Q�<SB�aL��註����O��a�����'��}ӆ����0z�83�0����Q�8t�e;w����;���j���O���.����;��/5� ��m�A�@�Ƿ�<1�91��d�8}�zB���t��J!�﹁��x}�}0�7'��x��Jg,�Y���ݧ�e���ɳ4K8��L9�$�2<����|Z8�2@�����g'y۹��373��;����=�{x@_d;� I:p��p{:]��n�^(�cM��,�.�v�����I� d�1��)���N^I����gFϓ���|���f���~l�?K4�!g$�9�H 9!���"z`�)���t���h~�p�N�/rg=:���vp�㦔���0`�/;��)L�N��}�{��p�G{(�9��'d0�H��_��!.Hp������狔CV;�<Ja��8A�$�T�p�
CW_t7�AѰ��QӦܳ�i�S�
@8x�4
��4í8-n���0`~�?~i`~��`���(���ϙ�0g?~v�i��g����ǈvd��?|3�0�����=s�t�@�=��9���?�Ӆ�(x� ��0~�+K����:Eקɝ�Ɣ����<SH3�<�;�ӺH�?������C���M9���aJ0�`�/�)Ӈ�S�;꘼`� �H}�4Ҍ��.b�(i!�
Cx�|��B�C�ȗ ��.�s	w��Cƞ)yg��<z|��N�08O���)�g醚N/��@ &	���C� �,)�R�Os�-0��<pВQh���^�]���׆Yd0���N�Zx`i�@��:|����h��H���iM4e1��&�fS�
L��(�8P!H3�~�0U��3��0�Ʌ.Y5�6h�e:�a_s��8t�aӇ;��]ǧ�p�CN��s�"��zt���>A��4�3;8�
}��<a�)�������%0 ���!�ts��pQ�B�`SO;���8CUέ��#��<xf��y�E�~5�~ ��Z>s�y�ܳ�=��n�:I���ӱ���}i�S�����ru䧎�{��4�f�k_�M���`��;���ӏь�Y�����ɫ!4#K�E3mt1�g�L7�5�&�4W��É����ӖΝ0y&����$�6&�_ܛ���}��a���L�}4��{��<qW�Q�=�;ݞ<!�����=�m�5�#<o9�3�O�{��
a�d��m~O��u��;�yq�iy�N�L3�%>P� ��_O��M������,�0�?M�ӽٶS��ty���f�i�H���S�������k^��e8~<3��<�vzS�0�lf��G�x��d����yd�{;���4�Ë�+�i:iҦ�O��z��}�́��d���g��s%dy)��:�ûe��Hi��>ΌÛؔ�|�m��L�3e�B�0$�4��D�'��m��O���Y���'� �o�9�q�h�p6O�=&��|�O`����U����xӅ#l~w;17�7,�� �&���>��Ivd:;��O�;})G�z�W��w��<:Us&��ےq���L�Ns��N1�{'��hä^p�ngwc<j�ާ��q^w��gvM�O���c8{ݐ�g$:}æ��������Ӆ/2SG��b�����}�ht����峇ٶxwc<^u���6s�p��	D�~Rm���/q���o*|�q��l�~�wM�b·��?f���~YFs��;7����{��yN��:`��;����y#�'��g� ��Ƿ9��̟���9��չ|rrv�G9��&Nn`�7�{{��ʦ���`��L�l/L~�s���͞!�l��J�û��3�Z�1�:�����IÑ��Ų���씇'�{��޼�	Xqz���i��*l�`�t56a��	N��^�\ɓ ����ldv`�|4c��R�fE�㥻�ǃ��H\4����N�/I�@|Vt���g;wن��T���$yg�k�2���p��rO��8>rpͳ2I� ��+�xT��6���?z�!�7}��K?N���a�{ S���f����2uq��a�T�|
;g���y��7;0��퓸�C��O��\q�gw�I�*-(�go&��%�O�L�s����)��@{�:3��m�g���̖�8gG�e0�6,��ۗ�㻱�c��'=��Ý�{8����٦	���s���~~;x�%қ{�9�;���Je�H|�63�O�ܱ���ڼ��F}��00c����G��Ty���l{N��w�Q��rb���1vv�L<]���:Hՙ�p~OG�Q�Nw��{+��2O�f�����sf��-�l�Ʒxɻ����aW;�O9)���G����o�<��u��6Ӥ�x�>L�;��[휅E���}}��>Le͞�G���֛�yS���ʜ��<�4���C��B~LU�;�u�
x�n˦�מ��{�t�xx�{gO��g�🷮��)Ç�
1������� ҇9�1W�ӷ�f�ܐ���+H�����0g������gd���Mޑ���xg퓇�!���1�
h~��0�óg����y&�/2x��za�Kִ�[�$<t����5׏��*�)�^@fp}8S�(����x�����_\���ik��P��?��q+?���J�K��_��>�zz<��ޟߣq��?F"rfe���*��kg�G)������twx��;���4��O��6N�!��&)'O�;9M]�:��I8��י�)G5s3!�bI&�z�kq�I@���S�(T�t�QeE��bNb���4�y"������A��m�lu�k�|eya���&vɽ��i�S���-�M�'��5�7f��J�S�����:Rw�:~�Oq8�Ӽ�>M q� ���^�]�X��qiMXo�h,�H6����k3E!�Ks��s�&�����b�Ɓ��l݉�w����m)w�4N�L!8���ׂw�MQ��tT�ZA��}������xa`w��@񇌄��(�T�N�;�t���WY�W-�I'��oM�Sb H�'`t�Gk1еI���5�1�<a��d.�R
h�D��	�1R��cm��\a<�M	�j�Y��*�ru��P��a�{=�_y�S�8�ܤT��`i��^fNm)&�.%��iE��:�+!�E��f�sX�udK���Ȉ�&�3)��YĘ��8�e>�ދ����4�09����13WN�t�H"b
i��[�˱�1��7�4�k�E2n�5z��Cm�.) �f؈��4��CD\�%a�tȠ��H��#�5|pt���2c�sJ2',`b��CC��7�5�$���`��Cl� m��J�,��"8�5�U�H�Shm�i��!�Gm=f���w���)�2�N��n��'���Z�ߜ�(���Pu��K�B�n�73"��7�(�ͦ��\�n��S<�yu�}�h�a
}���"|�1Y*�s�SM!�:����O��7��ΰ��x�oT����4o����?�׏�{�x�m�q���zjx�uه�����{Ӌp��mݟ���/�?��yn���m��%�jm��^�9s��=��wnݻv����۷nݕ����ʪ�W��^��V��ޯ*�U�U򲪭Z*�[YU^��U��W��U�UmaUWp�� �>�����">����#���%�qYUV�UqUUUmeUV�4�Un���ު�Uz��W��U�UmUmeVme�W�Ҫ�W���{��=�{~�rHIU��Q
���4��U�*���UmaUWUUQUV�˻�V�UUmeU_+J�^�*��*��*��ª��ª�V�_Y��DG�}|}�۲�fwwU��*�Ux��U�*���UmaU\����U�UUTUUq�U|�*Ҫ�aUWUqUUUU[�����#��#����cZ��g����7��f�ZZ*?��~��~o�=,;�[�����7�X~���u?3�]Sk:i�u��%�d��	�xL,I0�0��bY�N""P"""abH�% �%� D����pH�N� �pAHN�$��"H���HA$K8'D��O���"%���Yb`�pKĳ�YQg�	�D��'���xL,��A,�
$I ���'�:'D��X�&	�a��<'M��a\ޟ����|��T���li����h�d�it�3J�m64#/hY�u�/j����K&iX[��4Q��m�5�Z�e���^[�5I����ri�1XUHQ��q,H[�&�o�/�<,��#e6���\�4�R���ͳ��X��f��dc�j�m��mڔcD�:4f�݉c�u�3�[��4W�5`l��5ƙ����Wv�S,/;kW��b2٦����)<b���!4I���Dƽ^����@6�m�nF�V�и����.�z�WBU�U�������YInɍ@����C.��mQ-���x��-�gmp�5x����lh�-�:k+]F �"]fݭ�w:˒�5�%���u����`Ѷ�l�Ӌ1i����9�$$ܕ��C%t/�cG�Av�jb6���f4)-\:Z�`�f�k�����t�@��Z�e�LT˳A�t�o�m=�e��s��kXRb6�]��YP��W7Yf�����ʙ��D2��-v+�+)���v\#��f�5֗KV���.T���[�M���Y����Nц.Ě��m��~�n҇{^f�1	f�*��֙&���v&�62�΍�a�5��1�LL����4���������k(!s�� �����CA2�XX�n��ߍ�$8�f�������nA.6,%�k+i�&b'ቫL�g�l�9�>�ef<vz�Q��|q�IvjW�6ԉ9e�3���]F��aB�u��VlvIX�ڗk1kF��cB�)�ciq����&��]��YumHeȍ���ilؗX ���0Ku M3:lV��%e,e��Xڹ�9�cBW&����V��Aא��"�*$�Y3���+k��U��kv�����3�Lٰk��e�E�[��rn3%#��Z.tl���͚�;X�]Ve���O�>	�e3c�wW��GWB��5��u�+-�� ��+[�m��0ۮJ�d���%��S/c��M��&��$��.U���*�hu��[���,ږ��"�m����DP�Z�ֺh8�J%̓�Z˫�ê��BYX�,�[���.Ը	-��CS �[��ћS�n�I	�c>���!(>���m�uo�������㊖�cv��]*r^�jٓ6�kP��Yn61vu�1�b$�t)�i��\�(�m3+�c*6
R[(H]5�
�H� \�j$FЀ[G�f$c�$q25mk\���%��]h��xB�urM�Z@�ek�AU1-�X\�s��,��D�:4���6m���R]Dn��+�\�V��Z���z�L�ڸ�"�lk�L,2�K����l��E0Z[���0C�Fj����1u�JY�JQ������Xml��m��4Δ����
�
�lq5h�9��gBqM��NT�!m�J+H@�U�U*j�ڑخ�v�:��e��k�Q��\[����I`���͗[\S�la~}��iQ�[���R��b�t�M���շ5�ds	4�V8�F��j��W�Q6,��4-9b]l$�aH]qwM�,7kc׋��e� ������[�����/d�lF#e1���B�4�m�6M���H�#���h���)�lѕm6���M11�t�J1��ZVK�Q�m1���Q��4��E�MHc��l0+)�-�g[��W����s���+�}����[[���݇~���wwwr���݇O������ܻ���aߏ����ܻ����߾�>���4�h�if�tJ(J0æ	��-��~T�8��� ��n�j���ޔ�o��F{Heu�v��lDn�ir��Zg;xm�:��u��K�%�"`"��-�s�ݏE�OKC78��+1���x]f�z��m(M�94�����P8&.LWe�NZ$�LǦ���2���E��G�h@��˂Ԥ{l`��{}N1��W��JɁ6���½�fW[�2����t��b��j�������ɶV;�ޛ
��m*��Ϋe��0W6�U�4Όy�)4:���B�^n�XkohEe�K��O{].�'|�ņI�k�K��hD'�l��)P?��/�BY��?� �)��l��?�M4b����zS��r��HT��n1���h�[t;�tMlz��43�TY3z�XB���P�2��w��>e��~T��Y��23P�a��;����b�d�W%���U.d����*�����C���j�y,�
����"������XP��C\Z?w����r���LΤ�Y�"if�tJ(J0æ	�	쩙:NFf�E5��,�*�j��c1���C眭}���q�y�0=�CPM�,��������0�m
}���ܴ�Ρ�t�Pb�o��^�i�uiL�3[�F�x'"r0E�b��Rʋ6��U]�qŔ�+q��u�ı,��"P�a�L�c����X�����>ȇ�4�t.	)aB���]��o����Oaɥ߁��t𧦈��<u1[�sU�<߹�4%*��a��i7|q��-�DK)'�'���N�q��������' ��S���<��-��Ç4M4�Ĳ����:`�=���-�-2�hav���Y7�8a�ΛM�}f�/�m-��&-b��墲�N'kw֤E&;�W*�#Ɋj�&��7*�������a�p0�����&�������dD���6>�������֭}��B�c,��5���0�Ӈ,K(J(J0æ	�	�k�q	�&*�;�U׍E6TM��SM�&(�n�em�	l�$H��{�3Zǘ���UD���U&fK"��gs���\ƘV���Y-0ɔ�h��bO���Vr�|�<���o�TR�vՆ� �5��!��a�e5��8��'#Qx8�V�-kU�xK2�����w���^�)i=Z.`��(�A�/|��s�~��n+���K $Q��5�-C��F�`d�s�Ѩk��j ���r)�N��%�%�%a�����`����H�t�`pH��NOpS�A��=h|Y�	m���a,߆�`pMO�>�� pOy���S&/�P�J�'�S��>=�Ҵ�_��ץ���X��D2���m�n���7ޑ~/a�vL>�xv������p�Q�  �AX�<�i��4PrR�����4D�,�(D�(��'�<o�m�F5�-6`�i��!�sx:��PqlԠ]UR�1�F؋�!����n��ؑ��A�-`91G�̰D˾��ه�A�j�� ÎŻy݀z��c�,�i~�֩��Pks��o��=���S����ԞjKKDih���n���BP�BQ�0Ox���J��c��LW-0
&N�8p��2OD��]�|'0$�H?�v2�Wr�����X8��a�3'�v��K	'�P�E���5J�V�����q�V�-�6����F
Z�Q�UjN)P��Q����$�Tff�i��u�u��]�(J0æ	���c9\��*F2[��g���v5��f4�[3.&��R���Ԗ(���L��[�''j5�b�26�� ��Ż.+(�^m�X�3�����;פ�={ud�Xfa�m4�n�{�\��j�}G^lU�&N"Z��j��F2A�j�<�<�sS�xy��Â�Jt԰���0��6���3J�YC�w�������L���G�ӕJ�BÓa��d��px;=9%�g�̆f��յ��nEQ�M�V�kr@�G�*04O�l%}�g�Å:a�	��K$J(J0æ	�1!�TDI�.QHhdײl²5�t�GG�5Oh��*d99ܥUd��nC��� ��>mu$�	g��x��
�߾BW�zI�ȯ18)����f���톍�>�h���b{593*�j1���V*)��NF����+�}-_�˯�OGe3�5H��6cI��+M �JF�OM'L'H�4N�&��� �'(��D�0�8NM�8F������Bi:�׫<��[�y���^U�[˰���t�$Ҵ�:$�#M��t��sH�8x����-�ye�]o���VUC���(�(�pK��R�ao�xa:T�iF�'Hҍ��t�4�QRG���?���0��G��8~/Ǝ�������Ɠ�~+N�&��h��L�N�)Bp�! �	�0�0´�xa6Tƞ*H4�#J6�I��d�s����
t~w+����?��+ˬ��Y���*��yVyfZ[/-��ƕ��bJa)�a�J�$�#��=\f|�C��Ӳ�o��_�m}�2I�Y�����E�|��z����K������m�6��ռ�|�Lb�q��!�(|>
*�:w�_Q�N�/�z�|�6�{Wy����>���L��p�����ʮ{����w�SϚp�}�r�Ϡ��뗸��+���~�+0&Ob;��Y�R���μ��@��d�s�}�_�H	��9��6��33��l7www.���7M�����������l�ln���]�����x�Κh�Y��i�%i�������UU�P
�|'�Q#�QIg�����)Q6u�dC��J2ZS�s�622�7��oQlE3��U��G~�[n�~T�I��D��j20�'�#=��D�/��.)�j�"��5�sK��OKMı)1	�T��YJP�D��ZmP�����(UL.RqLк���K�"^T%Cs�Y�cSQ7(fT�)�(eB�ZIu#Y�ePʅ��Gb���0R5�*��)9��ZC>�vD$�~�g���[���,��hR%Yb�!z�d����2��|�Ϛu�^yg�]����<>8|pϾ�U�eiZJ�Z�e�.���^%.k��ܨ��]Id��9A(��M���'x�g���u�˰u��ۨh�0n��=�OC�%F��(�%�4Je�HJ�����S*qy5I1�D^(�T8��U$ʑj�J�Q�br0�"$���}Gi����K{U0D`����@A
���ʁ��mL� ����I��4 �0�FCG�&%
Y�e>�R���ɛ(~���������xMC��%���`���ß���1"�֒]��q�_>i�����Q�N�O$�EQ$���Q>����!mH>�+�'6h�k����>��:�y�Ne��Ç3�4�0��h�����j��v��\��w7Z���ٜw3�ܖ,Y?Gd��Y�|DQ>7?k�����,7"}s����pA Z�9kO�Jv�ƮG�""������_q���(�)2���F����~�DC����dM�� ~����V��FAd�h��Oia{@|�p�?C�r������{�y��0��f�9&#�����*�&�2�5-"�*��k
D�E\��-
R��Ī�&��x[D���nb�}�����
��)�%�Ҍ
	�1���+bQ:!ua"2Y??�$?z&����6��g�CQ��4"}
J0�!c-;��B�"�,�n]h^,�/�?�֭%'֨�|dU5��%���kWY�F�5T�����"�<d�,��l �����,	���?lN܁���ޛp�!���G�<��u�4��گ<��.pӂ'��Ƈ�M�{��g舩�O�V�zQTDD��P�M�&e"*F◽�e)H�T��]K�)ʬa#��w%�2�TmC
��.�E)K�:ԥ*ͦV��R��HR0"���d�1LXZE�ZF�в�UK
"3m
K"e��?-�Ȑ=��%i�""vI��IfDJ�Е�)��`&�:|��s-6O���{�w��[֍&�&	Җy$���A ���9*{?B�CB"�;��4&!DDܚGs 0�AM�
�1 �&��/'e2��g�*��%T*�L�O�ȽD�y��*Ib�qP�Iئ%=�T���2ӎ��x��M$�J4���if��p����n˚���UQjdK$���?2F'!���j�~�!O�2"Y�:ym��78"vRO��$�&褧�̐d�2)�"" T�d��Ro��[��!�"��d�Zb�sR2B��?�Iс��H�d
���Aa>���������jT��Yr��	������ad2,����H�S���'h�?0�a��(,��|*�!9q�"Oe�I�P���ȓQ
3g���PDdA=T��
PDOIdpa�qiр�"pd��P�~���rd��0�0�Kd� 19=�S ��*C>��,&%��݊Y����-��P�!�xy�q��<�: '�I4ҍ:pD�Y��.��������j�Aw���5��B���ꪢ"2L����s������
�!Q�-�bT>�---&eCJ&��fT"%�z�����avG{ӹ��.�Ӗ�ٮ��~��pd�&I�Ov�CH�
T�����w$���v���I��N��;
N1��y�a:!��I�)JL(w�QvZ+ۺ֦c*�X��?mi�h�Oa�(��m6bX4�Y�M���}��,�'�Jj	6$����ڴ��B�Tp�N頛��ԧbq<��T�*$�ɣM��N:��tM4�M(ӧO	��x����P�p;G
]�Jȉ����Vf�O%�QY��zC5ld���#���d}ǽ !I��	����̈���e��R��<F~�����3;Ϊu>��δ�9��vc�r1ӌE>Ȱ�rE4Ń�Nrg:��������L�Nʲ�k�'T���Zڿ��2UR�uƔ3>Y�U^�)�ybɑU���9ed0�"������a����b)�x-�;�cr�.�Y�ֵE�s�`pO����!�'��i[k���)蜂(|{<`�ё&�)ު�x`��Y�72��%�.̤�$f����}ѹ�)�L$O"$�'��}����d��Å��?U����ϫ'���n%�-�i����˥ފuPaI�Yk.��,�ʊ0�l��4��4�M(ӧO	��x�z9U1Q_T�ˡ�CX
�����UT#"j�����POK!D�&B���6���/
T�{2'@�&�������~�L4'҅<����[�t�R��CJ/)򅔚S08�'D�(��=}�͝�)`�p%%4J
(��2DdL?�2�1�}|�����{\r��K�n�f\nf�:t�"<(Yt�����)9O��I��������),�J������q��VU.��))5��s9m�U����m��K���Ze��i��>i��^yg�]�Xu֝y��S
��qImU���k0��s���sX��"OO���)R�)11U[��2��Xmx���S>�l�6TP�֘�}95��Y)�Ch�SF�`��FC�wW!�{ن�d�aM��C3)�;w��Ѵ�0���c.:�����a�E2��쒇��b�SG��n\ѣr��=<�8p�p�@�f��5��(�$���0�m�&�gG�a)�R\DJ�)�T��)b{�M`��𝘱R�RZ.�aJq�i�<�"	��i�t���4�O+��}P�S�󊪂$@�E*T�!�a�v�.mI����S�2�ɂ��%7B��6t}y���Ͼ:���i�)L�G����� $�(�'�4�����.r#�z�1-)���E�F��Y,��O�����vR���K����X��J��奅
8��O�t.��U�3��RCX,���=�d��/����1U�*�jf6Rt������#�����xa<#B��DhG��t�|Q�it�Zi4i%aZBl�t�#HH�:A�I��RF�:a:a=4��	�I��&H�	�4�zi����M#I8T�1�	�:lĚV�4�:N�N��i���#LhN���I҉ҋG�@�b���;�UvT~>��d�t�2i:I=(�"�'H4�ƛ����~>�����������t_�t�v���=��O��i�(�V�N��N�I��ai(�P�p���I0�pل&˘�OM&4�6b�(�:i:Y:Y���P�d~?L~���E��`���G��Z4-6b4�4��㦔i�J�I��+'DڄғIҍ*�&��?��~����~�3q�w3�>���;��{؂�����e7\j�&�s�\i���^u���tO�.��<�5��n��o*F&���s*h�N�HH�z!�Fpj?N�H]�u�ײ�\�w���3�W'2����mb�rtS�s9|qk��k3;?g��Utf���ؓY6/FS~�F�]�qi%����72_��,q����;�����I��{�w�^ן_YKٞ�{/qKN>�E���7�q
����U���Gd9<{;�8oj~)������c�t�F���E� �õ��տ3�&�G��C]���Q�ב<��vA�~���������R����~wk��<�]=�k�)Z����M�VQ��x��ƺ���I���ss2����U]���̽�UWs3337EU[�����6�xD�<tA4�M4�N�<&�i���ύq0+i6p�S��l�[hZW`Yʲ�yB��׌�e�b���j�i3�e��pCZ'�E(�k�[4om�����|�����B�,Cl9e�7T�ȭo>�+2�s��m��e�1��ƍ���4�M�@��\c6��Rf�cHF��I�kh�fv�#��r����cq,�]be��bJ�����k����l�nRXTB�e�Q��5ϖ	�wle���������V��d�ͬr��R� hR�V�֎��k*mMM�K�.�����җ���b�8����z:b� ��[���>ϰ�s1��nZAa��` 	~טCk�p>#"����j���h�2lJ��M���U�ue��ֶ�T����@� >��#�ms3sw�� *ܮew�e�7��>��oU�()�᫽f����t��MF{`��:sa���:�3;[�}9�ǁ�?�,>6^Y�����7\��Qye�G��S�y�O��?	4�c�X��4<��A�	�h���xr5'����<;.Ǜ:�a;��m*���a>�C��,a{�S֕%�3��|�6)Z���NKh�����|�S�����>������2�?|p�Ɵ�,�ǎ�'�I4ҍ6h�����������Q��UX����S$4;9�{NӁ�~�?J'�{���{ƣ�u贞����F�n��\��p�L����r}!��M����c,>Y/�`ًGb�>�Ŀ�>�-K3�c+eA
^F��7k�.�^���G�D=
�m.Ćo�g9��m,���qvM@��T��n��.A�j�za��u6˭����2���,�˼���if��#�gI��ɎADD�����V �?~ga�8?�Tү0�n��ф���E܉e����Sg��f&9�ޝ�a�!H}!�hO�ߋ�k�����skh��F<1�G	3����>8a�� �#W�����&x3�D�	bY|�@�F�rn�g1���>`�S�vX,n�x�^|Ѡ�?����0��6�����ᢝ�k�jR�x�O0�Ϟ|�.�|i&�Q�<&�i�Ȳ6I����.�FW�5ޞUU�0M����k�N?�&>
]L*wC�p�4"���ʷ�7u�G�34oz���ht)r�L�l?C	�A"Ln�Jɭ2�Ź����*0����'s�R�>;'&v2�І����1l��O�[���5��b7�9����Y!}�(��Z�tM1�QZ�j/ul��m,���<���O04�M8iGDO	��x�n�;�i�n�r��������ϩvP�hO�#b�2�Zd��uȮ]����ֵnBE~�����QR"�r�jU[��!x >��0zP�X��c������<�Z9���q�T�G�&Kc�����bۓ�E`&�a�S���1�у�#�܂1Ņ�&�2����O-R�X�k7���ծ��i�51������,]r�ew�3֥V��*1��%�e5
&��[����l7�GF�e��as�h^��k-��܎�B��%�S7�/�b�X��&��J�'�Δ�?(��,�����>Qb[�t�$�8Ҏ(5"pau�{�\��V�SG�.Y��bf56��NM��2�Xm�<��\:��y��e�Zu��iZͭQ�����yX�19 D�$辶h q$A�`{?C!�s�ݛ���})���e4
d�U�T�ȝ=c���g!��J:�K!�0?u�Ѹs���?6߱SW�<>��ѐ�&�8r�Ѹl���X�?F�|�n�R�ᙚ�b�>�V�>=�n	�a�����6��p��~=�j��},�]��1������S�>�җqO2ۯ<��L�u��<�(��4�Oa���O�90w�
�~�){3r�Ø����|f�~<���U���ީ�;�xzA5!�
j�3}��33Ӂ������N�L������nE�;������f�mf�h�Q�ұ�*�{����{.`^Ɲ��*��F�F;*-���0s��T�0�2`�u�X�v59�U��2^u�z���QxQ��KO���LH4�NQ�=8z|t���^��Lj��hZP�O0f*�Cp��aɐ�5Gf�Pѓ����a��9k(��b~�4��d�p����.�\��b�K����/�.�IN�ye�sU�4j2a��(X|t�B����bsSc^��{ᨯ�>T�=<��e4j-��sU-e��R����3*^)G�Ǟ�/5����;]vn�L���b[L��Ͷ���2��T�M8iGO	��x�=p$����;���n�QQ�Ó���p�>K������%K�L�a$Y�� !'�V�U��)2��/�rЯ������n���rݕoPw�>�j�p=���}#h9ڳ�7H��eQ���w/D��2 �ި�B���(L���w��ε�}x6�Wx+���-{�֡��K�y�}�"nPO0CQ4gtA�C���w?
a�0OH�O҆DW�p�~6
R�����G��z?��&��\�Ա>�x||l0�m�h�ɏ>�n7�棑u�sB�o�̷0�7J!��&�	�T��
O����b��~�h�����Yf���3m-�?'���O���n�)CΞC�܃�����i�����0��~�LH4�NQ��i����L�֍\�G.�#��4��!�)�E��tSE�!��}>�<��za>a�Ҙ}8����E���L,WiJ)�h�i��������_�k
��>�����q�\s��*S)������j=��)��\�uy�[�ҧ�y0�ES���O!J����S�g���u��xzh��L�2������]
T��)�S��R��K��ό����	餤lBO��	��&p�R8i)��a:Y6Y�Y4�L1�=j��y����eo+�-yU����&�Iӆ���i:i:i>4�GՏ���S�0i�S�ϋ�f�Z]�l�;�S��R�[_��O�����y^W��i��W�y+�-�ֲ�W�-�|�f�6��|��Z�|��L+H�'��F�}�	:F��a��A�M*�4'D�'�I�4�.b��tڏ�M��h�t��N�N�Y�j��=�ݭ�J���>0�~.���h���??C���Nx�l��YFN��&��N�O
0�#H�
��߽�3���xLFY��}��N�o9�S7���m��|����&�j��o|�}�*}绗�q�2�s)�ŝ*��x����b�r�+Ϩ�_�^Gz0{{U3�v:縦rM�F���������I�!�>w�<>��NM�����;ڻ����u��ڦ����|���������/4��L|�ٓ9~�?��������������nfffn�
���fff�ª�{������J4�L4�D��4ӆ�pD�t�햪�!�я��!��wlt�0�{�"�L��<�.Y�0؂�����)��fA,?Y�t�ݯCAf�z�cR�sћ����)�;���D�?����b%ġ��*�T�*^">�f,�Li�I��P0���t��6d�a�a��0���0�pN�.��9C�wMAÔ���mv�i�|�.uO<�"������q~]X���Tk����h;��b~ܜT�IӦ��K�y_�����O~����\��fV�e�n�����C6f2��f)G܋��q��K'�����j�d�}�C�Sc8g��LѰ�)D����[�������̠x"��h�{^/�E�}�$�i�Ͷ㏚e�D�M4�4O	��Mw��53

#)~�7��n��rAi�G_ڏ����+�u��4WV4>p |��a�R^�+��H�A)آ�c����' b���������s�}���3�̑b�u2�E\`�c������Jbp�5����K^
��+�ͭ3��f��8�}�pT)qSA��8jC't���D�ٔgMK����pC���s���$�����N��0�c���W�de���j0Zmx��U]�>�8a�a��h�"��=p�DN� �<�i���^�S���L(�Xk5�Vc�﬍�\�Z� �W8���8���UfLŝk���{�aɵ����(�bh�~<t�D�M4�t������͢�)i�J����0�3�4\ˌe/i>�Vu�Ӝ�ѹ�K�炷��Ȯ�|!�)�L0����a�0dA/uU���KZE��kh��)G�{����۶����Lq��h�]�)�`��7
	L�_���X��sw�m4QNţ-6��d��
{�1��.��<��Ϝ|�.uO�y��y�Zu��Z_�e�ieEn��D5MKn�9'�ɸ�%=��=h�ŜYc������ǣn`�$�7��9���җFS�d����ݛ�Z�[�04���<�(p0!�a�����W��e�ᆊe�g#�:�-T������e��=�X"q)�"�d3�֍�����PK=��o�6ly
WƝ(�ĳ��0 M4����=>:|t4���!M�I���oB����6���`����ݝ����IR��}�����S'�+�������6}�l)��9�{ޫ�p��q�����G_a���g�R蚥6R�mv�a���T�*��Ye(�P���4h����,��08B�����4��F_�N_զ"���	C�$��$��N�<&�a����&�pӆ��if��
{��k��Rr�ػ���M�L�z�j�n�f�sKF�"�J�XuF�g� �Ӈ9s�Lrg��c������lT?��F��Y���O��O�{����m�[��ɒ���٬{{V����
���o��3���'�O}3�)MmM?]Zx���@����s��IH��,޳�+/F?���Ryϒ�}��v:P�
r+��+2��*2d��xƪ���'��G��lؔ8M��xV0F�_����E�?[MW�U�[��w+\�s�'��L^���҇���u�L9񆡩
�ʪ�<��<��y�\:�y揍�8z|t��������YI!�O1��>L�zң�e:kuUUT�喎��|ɓ����������j|�Qe��R̨��Z->�w}��{]�&#g
aC���v;��(s��*ew���ֆ�k+����lٚ���|)졹D��~����2\���8�Iڒ-)r��nU5��V�c�};�\|���|��<t�D�4ӆ�4OK4vI���n>*� ����8h���b�Z�zx
t<�E�"��4{��?!��e9�<��F�8���;I��TeE��z�֬\Y�k<]k�겕���i�L�q�!v�|8}mjXy�$�:Cӿ�f�;��f�/��n�����0��Z^6��:�n��%�?N��Yy�^|���-�uN�0��ӇO���=��[\6��n2湺sF�>*�!����l�����Ç0A'����Op���O���/1\�f,�ئL jY�}�XrL�!ga�� N͙;?t�F��}��7��c𪼡���)P�EI睊�d�ۊ��G=.a�s��
|�n��}ܓp�)�2PԪ�Aa�%�>���~�����e��N��OM�G�4x\|%�||�<��fV�y�V^_O)o<��M�0�G� �I���h��F�I�0�0�,�,��I��|F�O��͗��y^eo+�-w����x�M$�4Һi=:aZF�N�N�eG1>*l��>3�>*|S`�R�bn�(��O��K��ʧ��t�t�6cI��i=��j(�4�>����~���n�??���o�?��RTƚV���i����N�a��"�4�4Jȍ&̘�*4j,���|GHУj4�#N��M��
�I4~0��G���C���>L.>(��>��h�O�p�]?c��?U��,摆�Ri&�	ZBi0`��_���{�^O��<�� ��p�j-a�q����Y�٢�;6��.Nn�9ݘ��^n��o3w7��u�Y~�Ӝ����z���O�L��b��&�"01h���ߙ�a���?>��TS9��r��&'[���Fv�g���;ۨ�;��7i���~N	�{�8�Bff*���N��e{��zĎ"kP�k����N�3�i{�k<�!w��>G�.Luqw�����غssՐ`�p�.�cT��_oy�珟�U��R���;���%�^�x�3��[��a���f5��F�dMG��L��ݽY��Y|������Tj!�0�nH�0�31�����)�7$�J�U�$�ɪ_���w�n.~��������������*���������������� ҏ	b&	㥂$	��4�x�Y��{m���̣).	�6��ͳ�=�x�6z�kn.�6��o:�l�H�`uX�u5�oi
Ks�M�Cn�aLm���c����MB�e5fJXL��ݵ*��eڙ�pmM�ML�{V[���WP��704�B��e,���J�nơ���i�5����k�cV�^5��2]�%�Sd��)B����&̺��p�Zm	X[y���hEĬ�Mn�La�]�t��i��cb�5E�«$�J����,�|�Q�A��6̦�jakv�̴�8�m�2�\j��W��X�j֛m]��7.�&5uXg7�T�� K>]�s�ۙ�P�1rBA����歃S����~�SQ�����F����.�sy����7�����\۝/M�]��q��p��֩n|@�I���Uz�8!���zaC%��~q���ng߇a�܌���d�w�Ƌ9~��J��x�pau������.�A�CM�'����{Z،΋,ugn�,C�YF[�0�����x��g�&��W_�}>�τ5y5ٸa>I�\����>MB�	(�i��	㥂$	��4���Ç��O�Ǎq���4��UD9
}����-3��(������=gtR�xSs~���U9��0�d��7&� ����>?j�.����Y���FW�sc�9F����I�?G�$#߂*�̤ٶmg���kv�1EE����˻��/d_�gC���0����01����+F��y��>q�i���Np�<xM,ә�Rڶ��UQ��v���{��7ç��8d2�rMM!�M	fj]��^'�.^0�,uQgj��0t#�=f.4j.e=�>�}�o��W���L���C�J}CP�	C�ѣ�5
j��>������!f�ݔД3���T��
d����CR���mm�C�G�MC�&�|����'��"��hQ���8aG�M?~<t�D�N>=6p�����J�i�f���T�����Ϊ�0?s.��3s:~�ܞn���J!�������S5�u���s5e�NM��!����C���¬�=MՌJ��%L5�*�G?/|-my�rT�0�)�4�5-Ueq#T�og�y���v0�D=�~���Baӟ��X��h�~,l(���B�/�ߎ�F��G"�ҩ�51�iM.�o�qǚd�D�Np�<xM,Ӿ�>d����nIz�l+A��H3�R-�F�ؓLb} 	:xN��a+���<����r��OB�̊��s>_�b�)�JRQ��Ϟ��Ej*�����pg�U����u�Z��#.��
+�.p`vg�M(4B�&�KU��n^�O�0S�2XJ�٨j7�Ӧ��n�>��^�ueS*rYQ�e�T=EX�'bL4;[kL<�N���GS�4&��GS�vq?wp|����Y��&��~�+�7%:SQ����k�Ɯ-U*�72r��iѰ�*�A��n*��f�?W�U�UT��6�����>i�κ�]|��<�N��o=+�*�J�U%ڪ�Mώɩ��JF0���[gd	�rxPDC�W0�a��ˣ�χ��ۢ�l��(`y���Z�����4d)�xvq_��������T�qnr��,�n%r�ҋ�!�/�<3g���O�)M����W�SB1�E����ˬ8��|�-�uDJ4ӆ��<if����������GєюXo���'��9RɨXiv��}sR��|�X�0��z�m�ᜥð�(y5<��9�g�$�M�(ؑ:�nHJY	;�Z����Y��RΉن��RЧ(ӑe�����v`��)s�����!�N�CR�PO��qZ�)��(�3�,�y��e�e�i��Ζ�"Q��4O	�K4����r����)�]��m�*�ĳ�cl�ai4�~RwX]E-'�}נ���字l6�ɛ1m*��N��8&���Oc���:>�va�f����Xw���1��p�!�P��~���'
y'�?C�{�ɚ:`�2Y�Ї0����/yUT�IS3������G�pK��?�4���$�i��x��7�b �T�=Ҩ�r>��%�tr<���,������k�����m�U�����^� $����H1������al�jǊ�m�^)e5g�}�8�U1�m��S��AQK*�s{��^V��Ϛ�-%���L#����us�ߜr�..V��OO���)䰡���"��6n{�+Y�ǑS�.�J^�Ge�)r��*�����5��u4�L�P����b0�z����d�Ð�>0�0�p��p���M��!�J?�T��n��-BBE(��w#Y]�amR�i����D�0K:X"@�F�p�<'�:|{�������(�OLq&ښ�E�UU�S�҇��=2J\�'L��N�A4����[F�k�p�8Xd�)���t��L��4�l�3���?٩���D�K'��`nf���o��Z�ۂ�40�?��P�eL,�<[C��:�;�Jx��cp���6�fYG��2Z!ˣх�2����$�i���P�"pD�"X�&����,�%�ǎ�Y�>J�@��"Q$� �D�8%<"""Ye!B@�@�	��p���pD�$I0�$� DDO���$ADҍ8i�4�"a���	e�b`�"Yba���btL<x���"�N$'�-!�<tA>D�0�I A����N�J,�4ML�	���+0��M��ف�ɳ)�WD�Vu�]s����#Z�i���'�;�����&���j2r�p:mm���;w�����dc�#���sr�ً�ݵ潷o��*ɫ����b��y��.�®bo:���q�Xu�oZ9�N�ǜ|�z�S�v��>q��S��}�:,2=���p�&�����Nw.���s33wwiU������ݥW37337wv�\�����ސi㆖"`�t�D��ӆ���g�O����UTA��)�~�K7|^Ot5E8<�X`�����[j���4�f�]s�����ۣ��.�\�ҩ�;��&������y�����d���{fzt�j/�ل�N�����X�x��h4t��O��ff�pD�g��,ᆟ�0K:X"@�Bi�D�>:|[���Y���u�3���UD:y�!���i[BΞ�4C�6��R��[kZ���˘��7.*��釻��$��C},�>g�W�|S��b�Co��{���J0��N�L�S;��
_�Oy�*���\m����~��x���f�3�J햆Y��Ӝ���%�#��Q`��a�;��[<5F�:~?~,�`�%	��t��;cbg�#�p��T��
�ZR4���n�0S9`��t��5�1���\rdbt����`2L�� !'`{]h����
�Pn=SU��>32���m�Z�s@����೒��ͨr|�8�m�9�/��P��_<�؂�
���: r_���R�(�T/�J��|��[S�M�Y�pA0�}˗,8n�q�u�*1J��0�|�'WU��Hˊ�s���1���E,m,e���!�p��uY8X%�$5�!'���_�1V��6M-��4��P�?d=����0��� ���՚��XO�e�6��>m��u%	��xN�Y�ߦ.f	j*�3X�5�*�ꪢ��������ˬ$��<���%k7�Xz�!J�Һ��x��B�P�A�����~����pS�Q,C�-<Xl�fC��r{�"������&��㩛���!@�C{���4�S�v���zYxuhף�4�W�.xjG'��zh����Lŝ-�H(O��t���~��A9dH*f� ���Ô��7a���u��Z��?h�_b�� y)�N����m���`��O�+*>yr�3L����\�����i>,�П�r,��.��T�O��R�3��`?��_�nS�çA���{�5v����T���u���4�o6~0�Y��H(O�,饚vn^���k���7��ݛB�O��C�jp�se��L\l�r�������e�������O!�{�{�ML�T��aЧ��`ΟM���v��lC���kV�8'd�|�aEݘb-��gf�rL�i��*��i����w0�5m��<�ŉ��Ή�H�Bi�DK:if��kM-�&�±M}�ߛ�ͧ���춌
�J�ی�R̺ȳ3�X�e��)+c�� 	\�i��S��f5%�G��׉?<,��h�|)/�ߡ�W�{z�f���}���N���͊k׈Z�L��ف3ܘf6w����G��<-�e�*�k���e���3�|�k!�;���r��Q.�Ѽ'ǁ=)����S��jtU��oӆ�(tNçO3rC�/�r:�+6�y�
-0�&q��QC�\��^z�T^*�\�X��A�i�S0ŴȻ����a���ZΤu9���~��'�J<h��a�Y�0I(M8|zzt����:��+c3j��j���!�MC�+������&&���E�xkn���K�:C�K�:��O�cN�љ�O���h���4���|b�l\���֔Z��1����]��%Q�K����>&����5�#�/񲇽�u�ӓ詇�.�ξm�m�\$��&�4D�Oh����&#�G+�V���s���vkH����g��m��t75�r��S�6>.͟�>ٰ��������wV�H≊)�S�U
�d���8�|�a����j��MS1�MB�נ�gcؚM|:5+y�L�l���� }2,Ѡ��W!�>;ϓa��~,���X�"P�p���N���^�t�V��4e*���mUQ'������ٰߑɓ���,�}~a�z��T��L32�+i���zc��G��`yJ}�U)��f7Y�wLe��0�M)�����3�|�[W�^�!'f�R��/V��ˬf/�U���9a=�W�,XK.��NFx��0ɦWewI B"ABP���%��a��0I-��0K<%�g���:Q"	���"H�"Q$� �x�:%:""`� �N�uN��N�`���YL:$	$	�	"H""'�DD�P�"I��4�f�x�K4L0H	�	b`�`�%�pL(�:X�x�B�����xL,��$	'��I�F���t�	b&��`�A��
�TO.f����x������������d��B?���\��>�#yΠ|+5������+V;�*����i�a�鞼���8qcL�q�q�U�r�A���̪��Ow"����ͳ�]=:unw8�i���r�q�<���u51��}�Rw���^�g^.cS:�D[GVxVY�n�=�s��E";e�OG����p�;�
=��:����n5zl�Lm]��J�|���f��<�}zX���7���������˯�wW���]�i�G6w2�;i�q�fem���K�ȗ4�-Q����3�u'#�BE<�11Rř��24{���K5;�Y��O���-�h,'�s3�Yem)�9��w��_������*�fnff���s3733www��������x�K4�a��đ��M,��[>����"\f�-�i��]�4m��D��ư���9&S��i��)��Yl�2�	�l�n�3	eV���m�˥��)���m�#��b�����,35��U��H�֙�Ese��b�mXԥmX�.���v�hU�u���\�nm����WJK��w�o6�t֫�����n�$�I��R�k��[5��cl7MR�xu��9ƛA3l&�pA �a�v4���6t,Mke�	�v�-�%�Z��ktu��1v�;XGA�An�W��&�����Rb��jd,��k�Ee�%��tf���)Gr���Il,A�[�׉fvm����jSK23-N)n����+kK�6m�]�i� �Դ_�{�ǖ+�/A�|����#ș0�w��j/��c�|�ONpVaT�"�d�Nm�d�{�<d�ɝ3�l��5��v����$���H�"၅;N�m���M���~��Ǉ��B!��'�<j_9�sK�P�p����4>�[�>���	���>�v'꾘{0C3j��`�%�3�Ѡ�k��S.9��j���+QU�d!������*��F	�Ue�M�RθӮ<�ͺؒ&aF���ig�:A�	�����8���	b*E`W
�F\�Rc����i8���L�)��%�D�V<4P���A��:�6p�~�ܛ�C����0I�U|�,b������?(s��e�#lM�Q�}?�&��L�㌗Q򠝆?a0B��05�i�7!VT�o���a��=1i��i�;a��,I
0�D�K4�K'�ਰ�c�7�UQ�4X#�*��*���Yx��~̩��sB�-.��2�)�N�w�xn	����߮kE*�1Mj��:j�����N��O��̱Rqv�I�ZL2��(�eJ||�y�*��^9�϶⊣�mD�8���Kk�a��Ņ7�K4K4���ı�(Æ�>:|t���3�uJ]Kq�ڪ�ZTfL�ٿLQee��L�8�*5�����<�b�v��C�̿C����-�>��D��O�C�eEO���-鰤O���ܟ����Y?O�5��:P� ya�Z�?F�J���Z�o6�lKϞ��!dD_�tN%�?�0K�J0�i��if�6�zI5UP^'�t�%��3G1��<��q���>bn�;h�q�T;� ��lO${'��շ�;&�9������Սꋺ�
��g�'�DLH��6Mk�9go3�Z4���]�w�3\z��[e˧.a��&ᇦOCL�6C_'&��j�(�T���Yye�g7u�GU�1g�V�ɕ-YVX�4�ڲ3⎒p��)9by<����<�\?�L.ly�qde�7~��n�x�z`����U�u�u��L4�,D�
0ᆘif�i��T��UTC�g��a���`�L���֯���Q��qK�_�Q��tC�ёS�G���<�5�^>{�&}�)J�b�*QK�j��������A<��h���ѻh�ȯ�ܱ7���\���|�%�.C��;_K������ޜ4!������؇���a�z9(�p�}$����p�0�4L4�,D�
<4x|x|t���c����5n"�-fuUQ!��!�b�����kK6N'K�h�x@��ډٟ��P膏)��e����r��k����|��3�j�_ѧYu��,�N,�
�ڪ���)�`tOg���oh�,O�ף��yT�Ygηjz<�K����~�;�IE�Y��L4�,D�
0ᆘif�iM��2DԒP\i�UgJ}�~/����tCԙ��!/����]�Z-bVf�s9x�)�`�S��d�6�>DY�AA�������6nN��~тiVq����کUx�2�/4��KM->L(v���l��Ѷڛ4}��C�O�|L���Y�&�~,K(8a�Y���GN�n|�o�՜a��Y��iEgm�9�ɽ�!��13Pj�%�d|G�U
�-�x $�X��8K"���o���1�o��fW���Zq���';�"��D|��S�Trw�⏁Nͨ.6��w1B��z�o73Q��5���O�|�.{��Z\�Y7�)~��|�Bd�GD�qƋH�>K����fm�u�]a�Q�:�iy��避�0����nᲓ�
u�JU��Q��n��͛mFfV`�`t��~������dC�?]��P�<S�R�r�֍�s�%�luK��x!�#�w"���FQ�å�0�i�X�"Q�p����������خ���(a�U�߫v}9�1�!x(�L2|p}z�9�2	�b��;6������T���0*���06	oW��l�g]���U���^hY�'��;l�BO�r���r��"�	�	<=6=��y1��q�^S.2�.,�Oi��i%	B'�$�&	�	鈱(�,K��bY�<t�D����"&�xf!(�DD��1":""X� C T��t��au�`��T��D� DDK0N �$8&�4��M,�K4D�(L(K:%��Y�X�a�0���bY�����	�,�"Y�x�H$�B@��H�pJD�`��LD�,�!yd:֧�j{�G��7�������P6����h�;ۑ��$]���f�|�/ʢ��)'9}���,ζ}����z��=�81��?	��
��.)w|9�:�,X�w��Ξ'���g8�c��9�7��4�`�ճ|���L���^w���o=xU���J�|�Q�s�1�I��]9ɞQ5��/yd}��q�5xS2�7��s{3���4�yPU��ǜ�9���33www����������W33737www��ff�f���&�i�4�K�J0�i��if���UQ�CD��>z�y爵<eE
�4�Ԥ˦Kɍ�������C����0���q�u��2CrpC�za�~���s�mR�'�xXU�QQ�h���`�R���l*Ho?#
��b9n���*Ud��Qzp��Ӈ�f�0�ı�(�������O��:�f	k��hL�2��f�UQ�����a���L(#��V��5��&�aQY����Z�3,?#�5�xY�f��.z)襁��Tl���o[�U;��(~��a��6�����f�`S�tҚK0�\h����(j_��Q�O4O�ibX�Fa�ç��O��N�k��t3�ᨮ�t�rH���DF�n���h��Z#�g��"'ѭ� ��l<.�]N�&���\ʾ�)����W��c�o���*jJ�G�B�PZ2�c�?��W>�ABG��M��@�%����4u�=�	}�2�|!O!��z���m�}0�|;3Ֆ��/:��Ii��1.E�T�i��w�ϵt��䐍T�(��i�2�����54��EE12����(��{��>R'#X���m%���r5,�e�jL{�{جg�aL6��MK�J0�Y��if�,:��S����C��x���E����a��:q7=�!Ц�٩�ȵ�S�a�w�9�E����~��=�f�]��;���խvxz������p�NBS�a�M^o��j"¿��h�j�pL�;>8��hJl_�<����ߏD��0Jhz��inܖ����DA�J��`���X�Fq�y��m�����zU�����7W�*�D��=;68Q.��Gj�j�Ѧ����^};�R��xw�V��:'O�y���f`��0���JT��*�2eNY8^p0�
'
cm���a��蚄������W���_�������v~�)���&&�ib%	F0�M,��*xv��f �UV"'<\5��K,:TRzn�eg���Z1���%�~�`�U��VVҞ:o�0NC��{֮\�B�6&��5
z��g�?��9r�I�)Ȋ��a�����F���y���)��R�]��=
���iL<%�~?i������/������)x�l�j �� 2H.�PN�fQY���ܥ�:�M�`ڣ��nH*�L�L�S2I� �B�\���V�ڥۙ"�m_��&Bdեx��y�2Y������#[7y^L��g�7�w
I8\z�v�Ӽ��;.58��5��&�>楋{"�`�L-Zv	����"p��ã�m0����|0З��h��vr��<��:1���d�a�8{�<�O���Y>6l���lOO��&���-j_�~�7W�s�Ri�i�>��I�~TU.�R�%E�,�qfu��u֖i���Y��if��6㡥O��x��� B#�ЛڌU�Q鼬U1�ئ�ʗiMF��OG<�12����l�7��X&	�'`�/�M�DJyO��aD�!���>�Lֳ.E9�X�����u~B>_�(�q�~T�m<��ԧ����O:�����G�8I�,�����xD�(�G�O���><�Kn�Zho�U��~����<�oOM7CP�7<��a��p��.|xv�N�)���oB���ߌ;j��a��*fX���"����)�0�Z�U�6Q��N��.�O��p�YO��+�0f�Y��XS%-|s2����4�ζ���yכy���Y��if�V����9�I�n���F	���(��/��>���P�lB	�����VTA,W��P�ɲ�L�:S!���(�Bu yC��n=�����2�����ߒ�`�I��R�fffa����,��O�rpa�j�>�V�d�R�k,2���0�l4�Ҏ8i$h%	"%i�4�Di�M$�L0KX�'D�<X�xO:Q""H""tDDN�@�@��"'<%�'���	I'�ÅI�AL I(H�(� O	�8&��if�a�lF��0NpK��,��L$�:Y�<t�D��'��gDL,�x�H8QB@��P�pJ:'K O	"`�&�Y�:$�=�y�\� ��i~ȡ��^{W=�Zܳ�j��5���n����JV��ֿ�@���l)���W9�f��-,sZ+�U�6w9�������7�CAH��8Q~5z���s�/?�>N)r���ًwb�����ݺx�J������o3b����}�Gr��k����=�Ϲ��po�}6���¦���K�G״����r����w{����s�]�Ug�2\�.r���k~�;̙��Y�7��5=�I}���\���WV�-{�>��RO�E�
�,n7iT��HOlҭzKE$R�]��=}m���ie�K���5n���uW��Z¶څY�m]n����О�5@�1���������s����gww|�ww�n����n��n�www_7ww{{��OY������tD�Wq�y��m��x���^���aK��l��Ф؎��)u�5�5���lv(���f`���045��v��6���M�mq[�Ƅo1M�Y�)̰��Kl������й�h�u�l��mEn�F&v����P�+"D���٬�7#(�уB���j�Gh�M5�Z�6.�K,�&�\BͲ�E��^i5����B7�s.�0-\��m]��9q�0Z�A���vFmh�@��aq-���,ea�@k�h�j0��]�����rC[l&��Z ��r��K�
����f�m��"�涍��Ԣ�s�3��Э.�B7�,���h�z������XBYnu,v�%�i���Sjn�	+G< N�j�/$����l�wu�m����b�j"�s�X�}��S����͐y�li�٩�t��;��w�NG���]FK��sW}��O5��kEsM���CPч�J8�YO�j�J��Jt�u�-��[G=��	�5��m�j:r�*���=��:�M�.�	魫6%6?�nC�RlO=4.��n�n��r'�[.q��]l8X��C&}���	�^l�~*�H/�$��b&���tD�(Æ>>:|t�燲E>[,&�����D���&I�>1�V��G�	����g'��Ζ���K�xa�&��9�g4�Ɇ	D�
N��M&�o )Ƨ=�4�r�X����6���r��k�fᒟ��p�>�L��ܱ3\�>���50�w$�LEϯ�}E�<Y�	����t�(J0ᅚif�i1��D_(��&y�6�j�Ub'���{���s'�K�*��ZSr)xե)�8�궳VY�:G�#YL9�)����|+[�Q�2��
j������ߖ�"�};��M�5��uI��d<�6}kof�tI��n{<��D����M�Rh�����"&!��z'�Oi�h�Y�M��Y��ig����	�T�e�y����>e0O��8{�D����k
���'���	l��vY��i\�3W0SN�S��C&��?	�52z<�?��-3�ч���|����tJ7L��g�����O3�o*Tu�9jM)�/U�[�R��)T�/4ږSk���/֥8��8�4M,Ӧ�BQ�,�K4�E�����JPi�\�ʁ��r�Sy���z_r��a+b�;C����t >�ff���䥱ګ^��m�4��_�?w�=���3�Cž��6���ܕr3#����ԍ�y���1��o�~�dG�73s�M^�U�v���V��	��'���䶞I��J'�bQÝ�ya^O!�������R�v8��G�\eO�aLnʶe�R�Ih�8q_���Q�g0bZ�R�R�>��3�VלY��M�6��+o��O8x�4O�t�(J0å�if�i�>�e�f�7��M08%)ז��%�SQس��>ٕ)�F"�.��y�v�Fc1���g�M���3D�!Z�<L֫�1zƜ-nM%Er��:�����{!����~���ٲ��[~W!�ѹ�&R�)�;l�׺S�J��]q��"i��4J�0�f�Y��z���,�1@�jLiLޅt��3���3.eI��{�nΉ����k�3��TC����S>Q�g�Qٱ>�ː�K���gBn}�F�#O���	���g*��GA���aO���9E���Dн慠C��8�]J�;9����Uɖ��R�D�)J�f<Ԭ�f�
]�{���x��p�DDM0Ӧ�BS�2��6�o(�R�JR��e�U�a���D��ֈ��L�	���!�9��a�<�N"�[�7�3Y�Mh�F�K��P���4Q;�u��O=�=UJ�����-YvȐ�"&DO��#.��B'`�u=�U����k��2ffC��,�&|��Uɕ�]��yםyǙxJ�0�f�Y��M��rI�����5	`�"��U�ܹ���S�2�f5�bx)1���P�-B�������d2{ȳY[�_�#psÈ��D��Mn�u������o=j&- �5�E�إBݟSw�ϳ7���{�P���r�|�Zݸ�6��VӐ�|�C�>��ڧ=ZtD��Р���p�;�ݢ%��T�橬�t��˳p��Oa��9kZ�G	�&��F�B�,2�)��`l�a������q�6��b?��츰�o�دUM
V؎ʥSk.��ϟ<�8�:�采�Ξ�>:|oJ�V��k��I����0�T�O�=�.�}9Rг�h�3�3v��Й$�a�vj4���ie6��kS�:�b�w�1�o�/K�e^?�2��h�)`�?�>�=П�p��nJ&�����+�cҙJ%��P���rfi�i�e�a����Pp���O�%�&i�if�܈�K4��'��$x�ӄ��#��bX�$��D?$$���K<X� A:AS�)ӧX0a�.�N�;:��$��$���X�@��'����M4��4�L4DK:&(K�ı,N!bp��x�"$���%�tD��x��A� � ��P�8"pN�g���L:&	�'�<+����ܝ�u�����*����hZ�1{=�Սp�k o�6��G֗R�yZ�>��ֹL��e�AdJ|Q�REZN�r�c����S��n>w�Ŝӽ��jyޢ�!�4F�����tſ6��F�U]����E��s��ȺL��+S��\�F6��8�y<�;�\]��u�f�L�swս���Ne����ۻ�������owwww|���������wwww���M,�MDM0ӆ�BQ�,Oif�����"n{8h�N�f���b��$�zS��pG��i�w�ӊ���F}X����cTu��8��*�jdQE�'�,R��z��������Zʔ"�2�z�i�M*=����(]O�ӌfBdy�6s��0�X�e��^e��u�]y�[y�4�(��'�4�OT}�""*h֚��O%�zA��s��Q*�ɦ�5	"��"n9 �s��?	�h�f�����E��v>��|RYJ���7)�i)g��	��V�v�CG����z�4Q;��ѐ���4���4qȈ̈τ���6tâx�DD�M8i�	Ft�<i�����r9+�ہ� @;�Ȟ�Z���jUn�2ܓqZ�0�m�j̣x�3 �F.���֭���
dk�&W[�ޗ*�efP]�)r#0�5��f��f�|{�L���51g��w�4J�_r�i�܆&�d�c�p����+n�=)�2y�{�?ni_��8#���٩A�3�(�zP���Z�K�������SbO��-âsH�=5�I䰤ОD��e��l��(��=9pn�O�^��$��-��׊㰋!�Q��d�Nf��b�����݈��`���I'�:'���g�NiBQ�<=8||t�����77J݌��Y�P�T�foZքW4;:����a��'N�Op5H�?��Eu`����9�ތ�kF/N�䴳���'���3��&hS�&	�XQU��O��Bޞ�\Hi��[�+W�bhV�P�33%M_��/�KW�C�d�R���%��T��<wƛR�*9�*�s4�buk��L:�g�4K4ӆ�P�a�LƚY�\R�A� �z�@�~k�!�3�!�����m�~��9�pK�p��Љd�'Gļ�SI,B�+��^��!-����A����ʋ�2�S��I�^����L����1غ�+�Yk-�Z�N��v_�a�ڔꪚ�a��3�*��6@g�'�r�$�O4L,�NiBQ�0Oif��1�*
�*K����&qUb!҈��Gvh�I�uQNʜ�^F�{>�1R��e��L�^<���JZ�j^ӈm���
J�&!Q�C~8$��bC!�Ƣ�SJ�c
�-0��)Lk%(����B������A� ������rRi�?���"af�p�J�0�����~\_���/���Dd��5V>���ؤLh���� |!wL��#\nEj.դ�����j�Ŷ�fG25C��Fc��0Y�M�	л3��ϧ�i���2*�v�SΗ���ESzTAn�^S%��Koj�s��7��7�����~�C�(xvJ'Uvz~j��>��OO!�B��o�;�˘���{� /�I��az�V�Qv��QM�>��U��b'j}��4O&���� V��߲��	cV�����_�'��E���j�E�C����N�6l����0�M8i�Q�0Oif�����)0ˈ��5s"���犫����n���\���=�W��~9z�b�բ��V0���t���>R񙖎7(��q��r#V�3�"˗tۉ{��俿�迟��o*�/=�i�R��*�j�m>*��<�ͼӎ6�o<��.�燆�N>9�J�R�������h���h�p�X��CP��{6�a��2�>�¼2�Ɵ�g١�k���~���n�Ωʫ&�:ڋ�jM��ܔ�����m�>��J0Td��}&�vM�!Ҿ?M12a��Ɖg�ĳ�iF�a�LƚY��l���*`���dC�Xc
�Z:����/������74h騃==�!臚t�KJϫKiU������QO�S�-�9
��;'������v�UnmhӾ�U�5�W<��v1z�q�n�m���p��}[�y�4���+*��6l�8~[ᾷ���G��ʒ�?u���u��e�n�D����Q�����1�E�&t���q����,��h��$Y	��b,���3�F�E"-�D�"Ȉ��B�!m�M�4Z"-�h�5�DZ-�h�h��",DE���dh��4Y�D�dB,�����"-�h�$X�6��h�,D�mE�Dr���h�-�dL�E��5��E�"-�m�#B,��"h�&��4Y"�,DE��-�h�!�",�E�DA�4YE�h�Id�Y&��,�Y$�D��d�,�$KH�$�H��%����m-$�I�D���%�#�ی�Y�&I,�e��Kh��Ē�$��I$�Y,�2�X�$�$�H�d���l��HH��"X��%��ĉd���%�id�2Id���X�%��m"e��bX�,�%�K&D�D��-�Ki%�q6�,�[Kid��Y$�K$Ki%�id��H��K%���ɓK$Ki4��,I��&��KK4�M,�-�D���ĉd�d���K�4��%�L���D��e�id�,�$�I���i4��KKd��,�n��I����D��&M-#K�	bY!,�4�,I���[I��X��!-�%���g-�8[Kd�K$��BY&�d��M-�Ki�bdK%�m"Y&�Kɑ-�Ki%���%�,��	d��B[HK-�ibBY!-��BL�Sn|�Ě[HKil�Y2im"Y,H��I�ɓKi%�m&�I��X�4�M-�K%��d�k9g�3YHk&�!�6���8��3Y&$�L[L֙�f�6�8����ɶ�CZf��ɉ �	Z8�n4�L�BѴ�k#i3Z6�d�E���8-@R�(�UQR���Ë�V|�h���DE�DYDE��$YѸȴYDE��wr�rm�m-�e�L�Dh�-�"�h�X�dDYDG.\Y�4DY,���4H��E����h�m˃�94[D"�$L�"E�K8��"E�H��,DE�\p�r��Z",�h�D[D�h�q3��ȑm-�E�H��y	�"ȑdB-G$8�4[D�dMDE�#sp�	D�D�dL�h�E�h�E�[D�"h��4M��$YE�["h�D�b,D�dH��h�m�dHZ$khDZ$[D�"E�n�8B"ȑh�M"E�4Y�4DM�M"h�E�M��DE�D[E��b"-�B&�4H�!D�h��,D�"m-"��",�-�"�DYm�mh���m-�"�"-�E���DE�2",�D�-�E�dDY,�ȑP��",�"�DYD��DDYDE�M"E ��,��""Ȉ�$h�h���DE���,���""Ȉ�4E�"Ȉ�",�dh�DE���H��w�F�H�Y,�"�-�h���dD[E�hE�"mE�m�h���Ȉ���""Ȉ�4Dȑd[DE�dH�E�MDE�mȈ�[D�h��",�m-�dH��h���"�,���"�[D�dhE�DX���m4[E���4YE��"�D[D��h��D�""�dDZ!ȑd[D�""�dk"Ȳ$[D�D���,��D�D�#[E�E�"ȄYE�i��",E��d!�D�h�dYF��$YB�mё��"h�$X�h��DE�"Ȉ�,�"Ѭ�""ȑd-�AdH�$Y�h�$Z4�"E�"Ț-,�"�"ȑ4H�H�iD�"�4Z,�DAdH�DF��Y5�σ��$Z&�""����d[E�"ȑh�DE�4Y"�[#MD�2&E��E�Dkl�E��ȄY��&F�"#DE��"�",F��E���4[E�B-�L��["m"�B-5�"Ț,���F��"&DE����[B�H�",�F�dYDY-�Dg�AL����ö�ѫӺrgv��f�7����a�-ll�J1�ҡ���q㗫�q���~�_/���s�~�w3�c��p�=����?w����'s�x:�;sh彂sO_Ov8mG�=��vz:�.�O]�qx�/I�{�9=N7yݷϗ����g��'�ro_��=����f͛7�g���8�M����^M���������oͬf͛�g$BY�����Vo6�.o������o��p���t���#�o����ӹ�)�f|����f�fo�����"H�g���m;��3=}���q��x�vrʌ���������g���s�q�7��:����<��g�;�����[wg9ݧ)-�ۮ�����8<��p�1W$��eA$�//bBKZ��!<�$"/A ^�H�cl���,�X�'�;H��K����~��L������?$�~��B M#�H�Q#l�F�$f�A�q�Q�c�O[�:�;y�M7�΍�����o'��7_���7�oF�ާ~�8?��w>��l[����{|�lٳq��ݸw��V��o����[n�?��V>�O�����3z;�v�o���+����џ�>n���O�gf�Ym�Oa=���Y�8���ރ���W��o�3f�叚�#]���6�?����|��ή�����>��g�ɽ�8�a�i:>�f͛��m�f[o2��������G湘y�T���L�;��?"�d3�'v���ǆ6�t�ǭ���nJ�o.m���[����n��J.?V����&C�4.�6�2�J�Y*?���~�R&�:��z�`�3с?�;	�`��"������ٳf�c��{R_3�x`��ݷOv3f��9}��߱6���yx�\1�?���y���vY�OQ�&r�xw՞�>��F|7�����o��7�#n?Fr��8o뾦����f��f͛7���g�dM���?f���lٺ����<���{��y���,�<����Kg�����������iղ�O���������9�8c�^-��G���8�ɟ/�����(�H��X'�w(��-F�F웛r���::c6l�~��m�m���'g�<��z��\7 �zG��zۼ�a�rr>�ÑH~tU,ޘ&R,L�V�G���oNz�&f��l�7-�C�ή�{�~���<���ff�y7v8;�{���ۣ��Һ�7��u���������r�ѷ���_�|�.�p�!�ȼ