BZh91AY&SY�'� ��_�py����߰����  `\�� 
�@�P�۔H  %D�22DI}��
�}�R���13[R;�NU��
P[iD��8tI;�U�`e[���w`9v .���v� gnV�S��q�����w`t$t�2�l��n�@����hT�w(J�]�֛�\�-��%�\f�d   h  �� ��*zA����& L �&  O	�JT� ɐ4b �$�?Jz�Q���z���z��Ѡ   ���HL	�L L�0@�D� F�&О�=M<��iOI�D��R��2`� ��oo��S�
{��D"��TBȀ��"���@�cP��*�w����?Xj B � 9EB-�`�PoTQRIA?�u0@NQ�E�I$�I?L� +��#�����J�v�~_�n~/����p�I���~��N��DG"al�C�H�u���m�K�zf����t�a���|G��I�����v��[�t�^���rӺw�|w�o|o�髾�՗��0�.K�㒽y���j��K�XȲ����9+q���a*#ș�g�"9��ܢ��)�t���"G�[})�}.#��2����_�U��g�3^�ް��G��n#��\�+�*��+�����2�"eK9S�H:jRS�I�ܤj^D�l�Y�p��ŕ�l����(J�w��N�*��G�r#�V��u�9���eP�u��2/P�ʕ��<����uܤ���H�c0������5��ʸ����Z�g�8Μ�u��������1�c�$����h[�DhVѫ�l��<SjRy��ґrV��,���W,o��ήز�����l&�B��sK�i��5���t��\Ӌ�}/:ދƫ�U�%_c�WOnX�����B7)��%9��U>���U����7�m�xw�oV�C���z���cy��������ކ�����7*�9��	3�V[T���l�:ň��3���	z�x�<�Mxd�$J�D�Rx�A<����Rx�p��I����,��
,�(���A$4I4�C$nQ�j�yE0�CDd�Ӳ:Fr���\��5�5�zνf=fXh��###!��tjxY�-JZ����Ƨ�'�c�3xoa�f��i��{��/d�|�2��l�����(�VvU�N�=�dg�Fp�Kʧ�m�,�9��1h�Oj�m��ӗ9�}�ܹ6I��jRq�{/������Y���n�Z�黐y��D��D}�L��r����9)+Vp�<{l�<�[ٵ�y���L�Y�Ѭ<�q�|o_����Z��i��:�:_K�/��p�ա�8m��8�'I��a����7��|{Oi�7�oCb�6�z�m����owڧI�0��t�"�V�7��4��M�d��%:FD�p��V����X	��'eD�~�&�w���m�Q:��~ �,����Y�S��,��7m�D[�+�'t�ms3�Xy���79�6�a����ɷ*�����P�K��ɎivNDAv��9�y�Cݭڵ���0�����FC����Q�~��{u��#�r�:q��Z����2�x0�K�p6���t�5�l����z���c|�d$w9'�m��d7!<ߝ��q_)�����+t-�ǧ��ae�mc�i�m��{�A��I�Ǧ�x6uXu���.�XɅu�l��i�㙫Vnn�#sw^9Ӿ׮w���Y3��6	1"��סI��.�{'P�ce.�:�hjiq�����N��O�3dzC9�Nb�U[���9�k��a{04F����s
-�.��s.moâ�ZñNj�21P�	�$��n�Jq��紐��9��S�c�ne�1�2���S	&�BS�p����ٕ��/A{=�vx������.t�L=a(���M�O�ю�c<{{�mٻ�1�½܎���ִ�L���`�غWA���N܃C~<G�β�[�ko��F�r3����F�[�6V��6���_��g�T�X����Cu���0�7�6��+>��0�`қ;�b&��]��М�E���tC�_xe���i�dl!0�L��up�}�������jBk����QDӜ��g$Lac�2u�|�0�	�)�ɃFA�����9d�+d0w0��X�2�����,s7�?��^�A�;G�iv����
%ȋy/������h��aPˏo��+���O[j�<�z�8N�O	����V��8b7&�l���Ԋ��0�4�p�匳�yֳ���vL�(g�d�"�-��W @3n�dw0˲�m̾|;m�D<����!5:Ͼn�Y��q�.����-�n7����K��q������ݬ�j�L3�oF."���o�Սbj>�����7ن$����G�!T"�8޵��1��fdGsZ��s����׈K����x��ِ�R+lYn��fD��n�����G�gKMlf�R*{��������}�
�E�0#���}�Jo����[����g�����-bQn�篳Λ�	�S�l���c~�zQqE�nޡ@�p�?��A�Q��(8�g$�����L�T�D�9H��"D�-��DY�M9����q���[$q�Q��Ř�*Kl��(���V���-Z��_��S# ��19�1	H�&c�x��:�UӜg����p��a�Bn.#�(��[u���^7��5q5r���r��9��^���QIn]���b�:倭Z'���b/f��0S�$0h��|�A�
�E�U���a7"o"%������0j�)�5 �kR$��
`91�V���Y��c擂2����`Nz�g��m[���u�.���eΐ��M�Ec���q�5SQ���&�ҰB��&$K$���c\�0am�M��^΅�x��p���Ҙ.js�:���??!?�N�3nm�گ4�=������������Q�򀑄H�=��{�_���>s��Ҫ�Wj����UU�iU[W�F��� ed��3|�iUQq�������j�����U|��v$7�M�R�����R�nnkC7�xUUTUU�E]�{�]���W��Up�2TP�H���)"Q
 n%@-�@[�*��*��*��9�U�UmiU��(��ր�G��%0$�j0� B:�[�&*��Ҫ��^m�)U_+�UW�f�.h��Z7|7�n�$�R[&����ՓK]�������U|�/9��UV֕UUn�5"Hȓ4jf��#����k���W��^���9�UUTUUU���։ *\�p�֦�ւ�QK���Uz��U�^s��*��*����փ�К�"
�j"T��ZY�HKP����Q�C��������0�3>�x|�����B$G�1 xTD�����0L�8 ����b��N	�6t��}'D���:'JbP�%	C� ��� ����㌲��$DM1�jf�(ը���nD}u�q��:,��Ks�1�!(c��ƒNW�˳$@��\r�l �H��2a�	�Y�2��LcE��.O�,�`�*��N�E�.
Ӏ�6�R�V��#�!	F�Q�� E�o0d �ZِH��Shq���S`Z/��a9�Y\lw:�Ϳ���9�pHs��9�	��kZ�	b�ֵ�k@!�kZִ��ֵ�kJ�kZִ��Ԣ�͖2?/>��e7n[����l-ۊK���)$.qVH��L��V��dQ�iUҁ1 �����}^_-�7*����Q%N�y�e�p��?�\N��.>���=��8IaF�̖|B<
X����c�⒈*	VTq�$�\/B�tcm�C��M��"F�)r�q�M�6p�p�*k�Y��i�����-uK�3g
���;d,e�:nw����%��:@iG�ĔJ8��&�b�Fa��&d��1�&���VdR�J5z���v���k�+J����0�xEee�e���!.��˲Ȯ֩W�Ԫu��޶p2Cl.1����R��y��Bj�Ƙ����m�N)����|�ϕ�0�%קe����4��ܥ���lq!2�NK�(�*�U(D-�G~T3N�p(������aٳ&�#ƇN^8i{}��kIb[E&L��x�.�'7y*���R0�C��N�9/��$��������*&[�n<p9ޮ�U���}�n�"Q*���F/�p�8���'��A����K�-�@#P\
"��Q�4��wam��u䱡[`�����y}W��򗴌'���v��̺]�r�ļ�u)�b� A�9"wa�k�)�V֥�����R�q֨$
)u��1��q�I�{(.j����9pى��\�^O��&4B*�!��N�G�0�4�N�NN����!�F�M	�HTA����4v=G�ȣ��G#��7�K�x�>#Fi�=>#Fi�8FFI"����F�$x~(�$�9����q��o�w���.��V�$:0RO(�eD=�"�GfY׽Զ���<c�}���EGt��o���K���9h̜̔�fNfH��m|����m���qa�XY�6%�gF.���1�6�B�n�.�k�;K�&�&�&0��� Y�_��P�b���D)㣰$_H,f�T��
�(Ri��X� �IkP77C㦄����NJ�Q*UD��8��-��^����!�W�%]�jDq��S��`՞������P��t\/�u�h�#!)�� cB`B{=B�����|C��n�]ی�H��"w�v�S)�i$�9 ��"M�$h�����*�[�2F8�NHػg�6l�z�1��D�X��lF�w	f����JF�>@�x�#lw���jQ`�9�kp�I��Xt�h���!�$�W�IR��l)��d@� 8C��zCQ6t���9�D@�f�,C��:�Z�i-�4_�"&�X�] j��!�&u$�X��'ɠ��AТ�y�5�1�6�4D��<��.X/HY�F�!ȉ��\�*�\������B:j�5(��R� [Hz��'�-��!i#�h�e�1~�Q��
40zd���E�=
pt�N���kw�!])�0�,���4B�ڪ��RHT[�(S�Ig\0�H&s��"��6�\[18����i|&K\g�$�/	kC�w�-b%�Lwgq�����\��h�"I��lC	o(���l�lp�5�W�m� �6�d����M��>@�L96�㣶t6�I�
Cx�$	*�d��bA�H0(�l�$�}���9����/�DG�L�t�E��D4����$|��M)ä'(��-�qeJ��RRF.�����a �J���R����,,Ìq	�8%cp�p���'�Ku��_��OH�$�7-iJY��$�L�*�S��2x�Ƶ0�C|��>.�1,�8ÌOw�=�+MB��C`Yd��r���a�x�U�2���yv���	V�9㤱���pW�C�� �@��Ł,>�iR5P��|?�ѳ�g�� c�>��H�Dx�?��������3���#H���DIC��#Gc���t92���	��#��~�>'�>4�G��h���Np�,zL6h�4�zD�I#��龠!����Y���Y�+B}�Bv'��`Ù�S�G2$GM Ҍ:+�=�!)i�=�<�Yc9��e�扞�Ƃ[����K�J[ V�<f���e��]�Q�������(���"4��[c`�rV�+���s&�!0�!��Y`Ș��y�'��	
d���
1BN�W-�\˅f'l�����2�&��2�D^]��:�����-�Z���j��W��W��W-�Z��ܧ�A("�0�� ^1�P�F�i��jF��8�,�Ec��Abb�U"Yc@�J:u�Z�G�2��k�A���ˬ4G�t�j��f/��S9�.H�֣��Ɯ ��|V�C~����`�M�ې�`���L���Pa�)AHa����%>4m���,)Õi��:g�$��K"@�8�*a�yPP}�R.T%��)ʅBJ�׉��wm��ɻ���RC�&��4�����$�O�,h0W<����^I
�<HѶ�`�6C��S�.�MC,#>���L#��ѷ��];k8��F*��IIi�Vl�8�\�Ӥ�I�W�:m)�c��ŀ�(~8�f ͈�D��*ۈ�}&�)�h��"�bvg!�࢔��(���A)���+�+W�Y#����\6y�%T,;^<�t�+�-NG@�`�P��]�Լ�������f�L^ ��d�x,�	X>Rr���jJ^�����ވn ��!;R��6t�a�����s���.H��|�O�ta@I!�E+:x�A�e����,��)�2Z|a�(T�-�k�H�u��\s�O��x��q8�k��ɣ'�+���PS�	��0�H0,�sɌ�n&[P�X�pr����A������a�Ô�����e�m�i�u��)�h�P]2�/��.n��tX��I���%���n�3�q��!	�'�AM���&$c&&@�����±��Pn�N����-q�	&B�y�B�Ԥ��(-�u��RhK�k������� w+�b�ժ�BԱs���Yn�"�Ym�b�]&,�+_AgX�W
�;db��"Ҁ���6J$1Z8�7@����(F����g�_
��(�v�Qᅘ��	�>�Ͼ<C�ل|���(�tzi�t���T=!�C4�"�MB�dx�,~"�#�<p���0va�<<A㧉^4�G�|l7���>M#��=��H��0��hzI��̨p:���c�PKk��*��fM��C����-Ľ�.غ���ޝ�W�:����oF��Jh� ��ws�[m�ym�)�۔�m�@��o-���m��aD����AyB��"��>^�t��n!��ps"M>�aGJC8��\<̛�w!o&���U�:�R�Q�%�3�i�*=gh�_QN���6vEL1H�s�4gi�(v\�u��Adt��pۍ�ڔbܐ�|1�3
_̳�+�m�QiTx�n������rd��!i��(T2�e��8Z�-ډ����LM���#�G�I�{���S<PT�;Ȉ��!��p�+&���j��;FWnf[���E0����4g� �p,�8@��k�0���yNê��v��kD���C�q��aAӊ!q,)�z>XPb��&�8i'�y�a@��ޘ8���r�LL��PV�h���pѓv<��!$eq"RK<��y����P@i��(F&�R�B�1�:I�ae�y��L���
{8��ڣq@J��m|oL1��<��H5Te��qd*ߘZ�PB�(��]8||I�������.����$	#L"�i0܆�2c( �!49v�-_U,q�Q��,�S\_ōJ��vH�yqD_qt���(�z�X��U�Rd�1Q'N:؁�8!�8u3$Sc��R�F�Դ��Ĕ�q�<;�\E���I�����ͻF%��}���0mp�|��m�����Ct��a�	�4�x\,�<Q'��B(���L.ɡYjO�pp�#������줨�Q�,<o��"a�(��0��%�+i�j	��J�4x��Pt,�y�0l�.TI�ŭ8:⺬�k]$r�i�$�*�������Q��\�����ǹ6h�I�������>����G���CL��8ɾ���I��I�a��hzF�!�F�O��H(tii��#L ��x>���:;8F#���'����=<A���=<F���e��ő�a�|�#�0}��xj���2�Qh*�u�9��>�z����c�R�$}U23�Wqb�p�=֏���i���36W2wy����	�#LF�;�4�1���n:�)LM2n��"H��՛�菨>�h��	����"t�pETɷ�P���s�Wf޻��P�Uӌw7hsݴ�d�s^�O�{wFf��y���U�L��H"wa>���lz�;&�!iF{�$��un�1��Ӱ(	�ꄇC�6�])�	YI�$�9$d�*A��°L�"&BT��
k��`&����DV�RÎ�

d.�Pm\�~OOgז�m�n[m�M���m��nr�m�"�P0�-�v
"�e�>�D�+)� H��P�I�T�N�8�	�b �_R�4�KN�\�C�.h�P`g9���r�`����J���Z)aXAIA�g_;��Qd��pp7ǻ&�xk2FT�NF�Y8u�$���(��t
�!␄5}g�8�`��8�8�R���C���	0,,�=o�y|B$���CA�8=k	,���RQ(�(0�J�9G�/��{�I%4wx�fic��׎i%��s�X�^G�G��j���q�_7F⅊JD���r�G��ۈp�W�E�x|`���:t����ی�⏋l�!�Frc0�̞���&>*�4�yL"�dD��q���i⶘7"m�E$q����YHI5��Ej)�)j
D��wA�<�:aм��X���]T��h�a�c��]�X�U�č]0��h���.Z�Ⴥp8I<�Ո�O�z[���9��e���q�w��F6a,s���	i
�K��J��d����>F�,�U]>:t��g����wbc�%Gۊ���
TA���'�H��~�މ�H�#����W�zG����Z\Zb$��:�k
 ��,0,&�s]+BӸ�b����(�B�%Zۦ�(W��E�/R������V�Wњuh�YkI2E��%/s�0�&�g}�z�̐`n$&,x�ԋ"!Y�1L�;�y����c�v�d(�N��Q�\D����PZdL�Z'�YJ���p�D�A.)JiZ٢tY�7����;�.-GW8>��|I�ae�2L
��$���V�m�%"�RJ)|H,E)R0����(��$��(�N8�������E&�sL�E͝(ݦ�:�'�N$p���D�;���A�|?F�#M:N�F�4'F3Hf���NF�v:4�4������g��OG���<p�7�Ğ>#G�4~<G����4}<t���dy�!h�z<(�tG��W��}����t�:�Fĺ��^�=+8(�zg�v��m��m�m��m�Z���m��m�P� ����N_C)`�<(�֚,�OzV�zt�4�<�WQ*Nb!�I��Oa�I]TQK��gJ<Ia�e��%��a]v��e)��Q$#%B'`Ha�]�#V��ҎB��uaeW�ܥ
�C#\�Y�X|�PL1SR��>0��'��u��<�C�$�*4NBbq��.EHG�cimDVi�*5�72�8�)ɍ%K86�Nx�4��ۛLFk��6pD�U_~����L��\$�"8�� �L>�Qh_['LD��Z�0")F$�-�,�s�w�����*��Rp��fݶ<��(�ۯG8
,<�D&����pGD�)�qk���R�E�A�PD�}H��u��q8x����K=���p�(��j"U�g�8w�lAb�(a��Q�r�%�q-b��P
�h��J��1�I\�X���h���I&�08c��q��H��xd`F�03DB�%�!
�ڗ��,��h����R�bd�E��*f$��l�^\(�����*;��j��-�,�T(L���qù'�9��G��%�̎$�_u|�8���6i0,(�P,!A�q�#��H�!*�ce����m��x8A�loOC��p�T�6�I�!Ǭ.�u��N�4��pB�r��ň��̖J�őf�����>��}Cה}SU#�p�{��j:���p|uY�҅mWV�p�p(���Cd��gU�
����(t�b�8s�:�4=N�2u�-��0ݽ�m���L���Ԧ�=pNBX��2Q8J$���I�~4�8l�#O�'&�i�F�4�6�M���(�4t=cӄX�\7�txt����Ğ>#�����#���h�t�����A�=���:4�'�O�N�o�Y�C@�2aA��f�Ȧ}�X�z��"Y��CչT$uh�d�R�!�����0"�E�/c�"q̆v^bYD��K�/�js3	�^H���f*��e\A���L	��fuG1B��s�V�<b�Q�"�RF+�F\��-�mZcƈX���HDIH	v�X$�4�Q�)%Ʌ6PP��_����m��m�嶻k��m��m��m�Q�`�'��L�(dB-�m�\"Wh�+9C�q"�-�!]�F�0��I@�}��	�a�I+�S(�<�?x�CzBk��1��*O���<�T"J<p,)>\��C�<Ik�딽��֭}� B\�U��6B�,��)��fjZM�#�p�6qO0h����dw�0t,(�N�6��H��Q�(�#��}=sB�!Ç*zy�qx�-� �R	1qH�*�ב���z�6��IP|=��|48���q%��k�v�t>���GF�p��w�����vx.$p�0�,�Q9V��'����G�{�I��X���E-�orbY��[d�V+�����b�Z�hBh�y%�iԕS��xm��{��CI��u�2�=��T���t�|�ͯ�ѤD�"����xň���N|Ky�`a�B�d����E�1���(�N���#�a�E!f"�����y�G�)����8p���RQ��^H�qxɢ�����29����{�&Y�Ʒ#&��ӷE��ĸd�R5L�|Y��I5q�G�O�J���0��ׯ��ƈY�rD��So[����b&'�<Y�=jև��)�.�h���	>��9�iݜ�dd�IC��╮IsQa�_#��C���q��d��V��E�$�0*f&I��@B�
p�$�ɿ.�KWT��"�x8��ܞV�.���F#��QA�$�淐�����TO ���n_���&�S�S�2rB1t	�|�yQ���0:R.��e�!�:>������I���4�����prhF��G4��K"���tiY:�ig	��83�Häx}<GO��#����f�O�����:G�<I�#ђl9".m�qv�Q��5����ӹ��z�z�$7&����6���}��^�%�:���/w�om��m��m��k��m��m��mdP�� �9����R��j�.�;���;��8�OG<�i��W�M�)a͐�n]�Ρ��F+WG�N	0��-R%I�s�����sD�6A�GWS><�U��|������κ5jf_lT|�B ��J�Y�L�1���;�Т���ZE���b5|R�����R���MF�����q��K���V�m#k+����0��cD��8�J-HQ&g�6Ϧ��IF���	�|M�Lܱl�#��D||��K��Y718yqw��1�e+��ѧ[c�3,�a���2C��m��"�
\���t�GȤI��j*��9]��b$qӂ �R.�4�q�T�{���P�#�޺���U��|t8w��zLX�m�S�*Ŭp���{����᭴i��iԔߎ���Ť�m�X�:�F��
��Mw�'f<$��@㈂����)�dL8��8�m��%�0m������>R�ڂ�k��ڒ`m�Ξ�4�$�X����%;Ki�QMD��L<!r��S������Zg�UE���2A�<�Z<4[�������*����$��I8a˳������ӥ4
w$�!sE۾&���Φ�;&����UD�EBGé"kN���xq:xq8���&��c��ӉFA'�кP��A.ti���:?.����	�V�W��vz����q)�s���:���D��vv����6�ä1�}<I>��i�I��9���6iG4�l�
؈�F�F��HTa<F���<>�#���f�F�G�>4�GN��e�A�H<ܑ�ɰ܏O�瓇{`�1֏|��	6�Q��4l~�U�1���w�z�٥E���A�3|^e�5K�G�\E`IF�g*6t��OL�b�����=]�e��Ը���}��H`O���W0�;`�����4i��b�^��qc<"'��������_����]��7$�Ka/!�Ta�ёv<��H,�ɻ�����挴��󑈻W�9��K�2��8)t�j��喂+��ջ�?L̏�CiD�����2�����T��/�������mv�m��h��m��m��m��� �?���i?pD�[wQȘ���(� �[d��⺰��~�_g�8oy{�q�d������j���B�p|R�tT�$�,,3��^��iP��O9�B���X6;c��I3�xZq�RJ�q�E�t/���7����|�|p����&���-C�(���
����[x���0K"415���X|����J`%�MQ�N�xQFL��ː�<l�R�X6�u�]\%w�R���K��ǀ��5<<ZZ��G�>\K�|�nPT�� �"�,�lA�z!n<�$&p,30�3!p��<ar��%�,�F&Zi�4���XȈ��F|�B����-��qi���kk�Z����6���߀��"���409��-#)R�ѿC�ǻ��_��,`���2��M�H]3��8lj��2��e4C�8$���zqO��i��hb�\�������p�e�7ˀN"P�Gms�E%�0�� �г:�!uj	��ȵ�B=_*'�u�y��OU#�8p8d�/)��/(�+Z�_��5��{4�qiՔ�妡`P�V�cr9¯[˹."CP�R�ݻE�!�?n��4R�V�6�5��ŉg��xɬT�&��iӷ��v�4F����Q'B�8?�
3�K�wbë�J^���ūN���5�31S1.a5��k����k���$h�h.��p�Ç0p�:A ����b'؛,��,���4�4���O������a�a�A�A��3뉝�;��)�ud:��L�y���������ѹ��j*z���
��
�L^"�T� ��2gs:}C���xz�Ǜ+�p��$��vޞ�os|"4:�}5:�2�ժ�cǏ��v]��m��m��m��m��m��m�"��G�+�q5�oS�zj�N&;k��x�@���H�.
Ǝ��x�z�Q'�����R����}�:���r�\�f&�dp��Gڥ�6�C:G.�(�6���/.�Y��K(������x�lfF�I�I�1̎8H�"ԒFA��m�,��d�
&G�t�k�&�qyF���ZG��n�I�č�����P��D�i�8�TA%XQ]^lEAc(�\Tm�$�N�u��4�.��6�,��{�q�B��ҳ�<Q��aD���-t�p��fXQ:��M˘kE��O�Qp�V�?�f�L�Al�0-�Y�&��\�q�u ]�0�R��yQÆ$�Prm�h��������0z�ۆ4ڥ�FG���$Ϗ�o�x�x�p�pq5Э��Ū+J�Iz�P�F1Hԍ�;4�؅���[�vSN'Kl`�
���o-�V���ח߭|�Ł�����,F�ի�Ŋw�')�2`�P�G���Ĝ
DϮ`~�<xY�%���$�496CN���"|9��"�P�E�J<��]�l��@�>$�Q���)5���)v�"�h��{o�z[�R�QLՉ8�L�p6�z�KޒL3ʕ���a�PQ&[!�ԑ1��i����Z�-Z���j)�I$u	�Me��Ŝ'O��X�]�����a$HD��I$�H AB�?���~a�F˟��'�<�KbĄ8D K�08��o���c%�l"TD	�BD$P�	����H�"���AB����rC!�����0 0�0"�")
@��(��"� � ��"@! @�")+ @�� 
 4�
@��� ��,	(@��@�0 � � � ��)!��)@�� �+�+!!!��#$,Z�����RY,$�S�^�e�E�H2$�#! Ĵ� FH`^�� D�ĈT�``�h�b5�� H Q )� %H` ,`� B ��H H�M
 �
TRBB ā B�1 �H�		D��� H�H1��F�!, ă1��`D� $!1"�B�+LB$!$Ac0�"BbAcB$!$�H��"B��0����00!��B0B$�b@H�`bA�B0��bA��h���00	0��	 �B%�% �F`� B��F`Ā��H�� 0�� 1��� 1B$E�`@XX���! �X`A E��T� � 1RF� D`EH �;����+ы��	Bd�9�z���
�1"	$��b>RW�'��k����oT�fh��R##C�tBj�,��=O-�<X��?P|����\%	'�~�"g�C��=/k��y���XѸ}I����.��z��9w�Ξ��(�~������p�������� u~�"��{�ra0�8�n��U��XF"��A���),�����8|�[�H|����!��9�����=�c��|���?V)CܶḴ>R�f'ʙ��Q))?:k�^(�@��9�ܚ���O����Ϣ˄�1�����߫_\m��u���)�  �X�!J�T	J�@ x0(� "�*B(���E¿�4��W �jm�}'�sA�����{��C�� B��@�d@E	 Q%�#������/������3���@�h�G� t?���G�	���Yi���$*�'���Y}�ܿ�?�?�q��'�蟣�1��M��
����~c |��z`?�L�!�����bөZ�s�j�K
�y	 �{G���O����W��9ޚ8}�����>Ȉ"���R(
����Ϸ���QV��p��d�p��L��}��t(���׶HC�K>ۄz%��Q(�`�t{��� P�!���RQܔО��dM�f������/���-�]��C�)\ψ�'��pF|�ފ���o��hAFc�SӇ!1J8i=�`N����>A�S�
Op��o��??"DO���#����}��u. ���H���Q�&�ĕ�$A(-@�rS��>	�	�{S�~`�����6�}r�RA�!�ܸ!y#�,XZ��[W��,�������?���.��p%��)�bݶ�۾|�(e?���G�%Ғ�>	�=A�qC`�'���;���;O��)��HV�\0�@㌝?���h������i�~ !�����dr��M�����J�ۿ7�K���f�O��:�0���+�!��R�;������w$S�	B|p0