BZh91AY&SY��W���_�`p���"� ����bN|         P     �   �}���K[ef�Plֶ��Vj����e[[Sf��6�j�6��F��Hٶ��$Эe(4M�e�j�D��MD���ٖ��6kM��Z[�蝔(,̚�VMYj�5Z������$��jJ-�m����j�5�fd�Dh=  d(�x�k-�l� �-����� q��eF� wT�3k`� f�@s5&��6�l�M�ٓM�Um��R����S�-�����Zk�횖�A�B퇒�H   om'�^�Mۮ��z=��͹��uא�;麳ӕv.�����ܻ�n�v��K�jU�k	��C��6��=���f��Nme��r�m��(�,cmF;n�̠ϒ�H e�ѣk(���z������x ��ם^�] ��� 
{���Ѡhz��}���hO�����y�< J�[վ�{}p��|.�l�Lb��֕����D�$�@ w��[�6������� :	�}���@ ��y���i�Q�p{�z ��ϫ|��li��>�z��U��wW��=�6�]��������{��x���-��@�Z٪�cEl�/�$�� �|���n�y�  __d��o�׭PS5��}�(Qz���|M �M��)�@�3{�}�U�>��� �����Twٻ�(UOb:V��!��Q�Sm�(^��'�I( n�>���D�o{�>�S@T���{{��W��]ӎ'����@t;J����Zot���Ѡ��ڽۅ(T���ધ�l{K�h�wg��ZԵ�Sm[JV[l=� �}�
 �}=Ǡ �N�� z{F@s�� -�� z{�x 4^��*��p@]��k��ҧF��j5��kP֬�֧�IH=d| >��y��s��ֽ�^���H=��c� �]�� �ݷ#���δSN��yx �2���{^�*��Fj��iSf���IH e�>�>g�
 twv^^ Cά ����t��� 7�O�# 
{K��l7=>�� 7�#@�Q�m%�ٳi񮦳�%$ 鯀�g� �-� h��7`�=vy�Eɽ;��v���m�E�mà n�^ ��� ��u]Q0Im��%HCϒ�( ;��G��,m��I�á�M�� �����ѩ�(3��� 2l� 4;���` �E @ 
  ��DH�ACL��JJS�'�4�`@�A�bRU5@     O&AIU=Q� �    S�$�I�� �    $�$	)T��L ��Tz�?�R����h�=H�Phda=���~ŏ��q�~�a;��?��d�,�{lK�P7޸8�<����	 $�ޯ\���$H�I"	��@�b	$������G�������'�BI�����m���	$Փ�Y(����C��?��?�ԫ$��?����r�,r�9c��S�I���Iʓ��)ʓՒr��,r�)���ʓ�NY'*r��)�$�r�,�r�)�����r�,r�����O9Rr��I��,r���r�9c�9NS�9c�I�V9c��S�9NS��9|Y9NS�NT�9NY9c�9c��J�ʜ�NY9S��NT�S�9S�9Nx�I�',z����r�)�r�9c�J�S�'*NT����,rʩʜ�,r�,r�9NX�S����,r�*r�*r�����Rr�9S�9br�)ʜ��%Y���r��r�)�r���r�ʪ��ʜ�*r�*r��ʜ���ʕyRr��ʜ�ʜ�ʜ��r�,��ʜ��r��r�,r�,r���',r�*r�/,�c�9d��9NX�T�9d��S��U9c�9c��T���y,r�,r�,��9d����c�9NT�r��I��Y*�)�r�)�����V9S�',r��,r��)�'��)��9NS��Z�)�r���rǋ$�r�,UIʓ�')9I�%S���9d���$�r�9�
��r��)�r�,���*�9NX�r��r���9d�r��,NY',r�9}X�I��9NX�r����,��9Rr�9c��r���$�br�9NX�r��NX�r�9S��9d��r���r���r�)ʜ�,��9j�,r����NS��NS�ŎX垪U�Y')��,��9d��ʕ\�NT�9c�9NX�r�)�r�,r���$�z�)��NS�9c���,x�,r��,r��)����,r�)ʜ�,�/,rǫ�,��*r�������*r�,r�,r�)�x�c�9NX�T�9c�NYT�NS�9NX�9NT�9���X�NT�9NX�X��NT�,�+��OV9NT�T�X�,�����r�9c�9c�9}Y9O�NX�X�NS�9brՑʓ��X�NS�9NT�S�9j�,r�9Rr���r�)ʜ�œ�9OV9d��9Rr�*r����rǫ�*r���r�NX�T�r�*r��,r�,rʮS�9NT�S��9S�x�r����)�r�,r�,x������I��,r���r��S��,r��,r���tX�9S��9c��Y'*N_9c�I�)�r�*NUT����r��NW�',r��r�9c�9Rr�����9O9NX�r���r����M�6 lI��b,���9NX�9c�I��,r��r�9d���rʱ��,r�)��*r�Y��)���$�z���r�)ʜ�*r�,����z�9c�9c�',r�,�d�<S��X�9c�9^������,r�*r�,r����*r����r��ʞ�*x�)ʜ��r�9d�X�J��9c�9NX�9NT�T�d��z�ʜ��r��*�)ʜ�ʜ�,r�+�V9NT�T�T�NS��r�,r�)��ʓ�r�T�NX�T�T�Y9eX�S�9c�9d���',r��ʜ��)ʜ�r�,r�,���x��ʞ,�����'*r�*r�=x����ʜ��r�,r�/����*r�*r�*r��ʜ�OVI��*r����ʜ�S��NX�S��r��*x�ʞ����9c�9d�9S�9c�Iʓ�')��Y'���9d��9c����r��ʜ�NY')�sǒNX�=Y',��',���*��NX�r��S�=Y�)�$�r��',NY=Y=Y9I�����Iʓ��d��)�$�S��#��NS��Y')��,�J�NY')��,r��N^R�NS��9NX�r�,rՒr�,���Y')�r�9N_9NY'��NX�r��9c��咬��I�r�9NS�I�$��$�9NS��r��NY')�r��,�����z��9OVI��NS�Iʪ��NX�9NY')�r�d���I��NS�')�$厊r��,��9d��D��6 l@؁�c&�M�dCbK606 l@���US��r�9NS��9S�T�Y')�r��NY',�U'*NY',r��9���r�=S�I���g,O�I���������!T�9a�Iʉ',C�Hr�9Hr�9a��)�"NQ���NT�9Pr���NYUTG��I�$�r�9a��Aʐ�Dr�rĒr�OI9a�z�$���RG,���"9d���9S�9S��O9S�I�r�*r�,r�,�����*�X�Y9c�9c�NX哔哖9d�Y9NYU�r�)ʓ��9d�T�T哖UNX�S�9NS�',r�,x��ʞ���)ʜ�����c��r��r�9NX�T��NX�9c�9c�9d���$�՜��r��*NS��Y'�x�,��I�$�S��9d���T���9dr��'�y����',r�9d���<T�Y'��)�r�,��9NW*U9NT���r���r�,��O9d���r��NS��9d����J�,r�9NX�r��NT��NX�yRr��br�9S�I�6 lI���běd�?�B�K��׍���f�G���QU���C]B��&`�v�C]%q�Ajɑe'Y&��*�L������*� ,j��7a�v���JU�A��ahs����4@JP�sL+8�cf���ִ��2b���T�֤���s^e�Q�V��E^��Hl��pD��6�mL��Vt�F4"�����3"ڨ5j*!�%5��9pZ�cB�PǶ��l�rɻ�7Fi9t��٨��L�Q\�Se��-ƨ�f�$D���5�e�+V�zo3=wLZtC�^��x�Z�nl��`b#�.n6���љa��sg�"*
Z����t�I���9i��w-�h�E�z��7-V������r��3cu��]�h��G�Qja5���V���oT"*j��6&���n�]��f�����z��OTݣ�4��[ya],� ؓu�W�%�l�`�a=-m��eݸ�Ӳ�����+yKƎb��[�S*�ذM����#�Pb�;CL����$oh�c͘n2i��)jyu5FkF[�eIt��Q�,Ű[Hp�mp[
���vļ�5�Bs3ו��t�E�s&M�-�v]�e]����G t��mK�1֛ܗsv5=.�f0l�r���&�6���5� Ӷ�Y�P��YG\���;"�Sh`�
��w���E&8v���]`���Nٷ1�t��w��]��nbzК0p-JK�O5�!r�`cT�l>i#Y�@.y,Y�M�����cz�)$M�U`7/�L��L����Y��Y��hj �^�Z��G�]����C6�
(Qwr��"�{p�ݏ`�Ʋ�nk�]�9TLD��_�˚[��薍�V�^:ńaL��x�]kU&��n�we�p�y��,$h�%ƥ�n�4����7x%L�k��q!��2v�,��k���ͻ��Ks64]��vMUz��B̸$
�۽����"6�v�H#&�P����3.;�SAG\���RwE X�+kn	Q��Ӷ�dm,nV��e0Q,�J�{mZ����QIn[]�)Jd껑<�����5*1�E-����k�q��,F�'m]U
+/l!�0�i+��'qv��l���Ƥ��x�Q%k'�m�{-�cvL7B�,ZyB�`�t�m�ŀ4R:%͸��u�K�sp�Jضee`���1"ƠV�
1ͬV�$�oN6�<��%��^*j��8���4���
lR�t��u�˅iȵ9a˨�ܗD�F��5��U��e���6�ɀ�����v&Dͨ��1LIe,���vUdz;{I�Z���U2�j�LÃF��y�!���x�b�u�X��J�Y@Ӻ�w2^X�JZF�tAj�S�5��k7eb��M�y�FL�Y~.�aVK�XƳ-�2�Ȓ
��&�èQ�(�z]� � R�ԋwE��B�;*�w�*solݫtpH�n�CXṸ�I�����W �y6�wM�G7om2K[����V8��Y+X��el������/p(��kS�e��d���'���q�U�wS[�M�`'�Z7ff^؏c4۪D�����*+��ԭ8vQOn'Ǳ�SFn��wH�j����'n�
2��l9�f�<���mf�D�b-Ïr�lfV���a��j��bM�ma�`CMGb����y0ڼ~!��ÛV50�Nиe]���*�������e��qH��L;�s|�V�x*nJr9���W��f���3L*u�F�h��e��0ށ�bc�T�A��
�,Ӄ	T��jR���ML���uL#�ee�-8�;"4�l���,cm�p-Oh,Ua�Wj��gd�f���h�5Uݷ��Y�M�Q��s2�%G�+��Hڄ35<ysZ����^N�TLlÛ��I��H�J�`���D5��P�q�x��/��	�%Y�a�om	���HVq�Ԟm�I'Y҈{��'�W�b�ݧ���ڈ(3nC!����&�TE�im����7����ss.-a���%f�Ia�I��-��ÙiGsWFQ����2�wP�����/��.mq�I�2
�AMV�W!��n�vؤkln�yOs'�n���l&�*�s@�,MJ�m��um�v�A��n0��JUK���	���3W�Wx�=���� QZT�R�6����r"��wvBG�ʲۇ4b��oI�牆T$���Xx��j���,��p�F*܏1ArC��3,�(�+E2�Y~ǢΊ44)b��n+��ո �A)uv���H��	V���bRT�Y����n�E����
�F���О�W�UL����p�f���&�.��V�أl�Z�oD��]X���� ƅ�i�꒲c1;���ȊF�˵X7r�:l�r��$�tS*�]A6̱�W���+R�W�{(T˔�&����R�S��F�%	���t�x2�K�6H�e�cn�\f]����X̔����4RK�Y@e�y7!yxڤ�Ѱ�˖մ�QK!r���[D���A7.�X��8+]��N��dswB�5�慍'�3Uj1�Ya�Udܱ�ܬp�4�j�hą+���%m����K6��.�*Y`ɬ���ٱ+��)
�{�N��zJ�S>�H�U(6�r� ��j�ǧ^����o5i�v�7��6��S�̃f
QwHq�U=x�lU5�	�ߨv9�D��1(�ɉ���rܩs��Ҩө�$n�A�U�6�me�i�E��!WUu˧#�Ƭ0�3$	�ʱb���l�CaY��fU��3&�t�qJ�Sf�Cf���i˩5f:0`M�����ijf���{G{4*�
&�	>�ޚ��t�)�夝;Z�U1�۶yf�$B�*֏��kX�z�̧w�5�-4�9��{��h[X4V�Px[n��#�^��l�-I�C�nV=��՘͜&�XHp�9�:2��5 �^�+ab2ʔ �EPڿYKj�W���Yq*���V�6-B����bL��:�w�'2�KZ$H�$J��
[w7��F¹);����@X�AX�� '3[�呎�ڋs,C�#������Cj�B�H*�eln�iǔ̼����q4e�j��+��&j�U�� �V�y���Ap�P�mV�&�P�)L�Ŋq'�X�n8�;7+A.Š1���+M%�2*���L��ً4K4�o�5���˽aQ��n��+%JfSc�t�L��J8�2��V�Ņu��V�w�qm:v�)*�T�xp��+�H�יaF!�ɂ*�Y[7,^�&i����[*7y�lT1y���1��{tLu�s^�$Sǭ;�7i�a��qL�a8FeH�e���QیA�C[Dg���Bb�k(�⨡���ʈ�N�Ma��ی�{��҂e۷YP�rő���*��f����B�c4��2�CY��� ��Ӣ��/%j��ܘ��ˬ@�R� t�"���wD�7w!��1-li�-�B5�ϐ���@Q�d��^�
x�落���*��V�!�@+�B����"�D���c�ڇJ�}@�q�ַ/;d��/F͖Xi�z�JT�#�Zܚ��c��Cm�rޣR�<si��U��<c��0��[�޲�j�#�Jb��b�&�)~Ҩ54�[t+[�d��!�%+c{�VGbnnC��A	eM�nY�cl��Y�t����5"�UW0I��*[o1�34ݬ��i��ӣ֒�n�+�<`�I �yz�[q�I1���Q�S�Hhػ57q+��G��(�ۑ=�81�X��*BQ!V�afC�:����w�]=��4m@ė���ʭiZݖtT�\�8)�(�Ǡ�$��4�ˤV��Sfn��d-���Nkئ*�D��6݋m]��i%R�f&^,N��kV�4n�!��Kt�B9TF�6¡pǃ,���=���M��j�b�+fk�l��f�������B)�L�qC5���{�Ue�m�6b��(��#U�YaإM�i\3 �J�ɥ3�d�ق��fk��}!3�T�֜R�;��2�*�����Qem�=�_��(���9-�X�6��M�ө�n����a8��+ �f.L��ҋق-��l�UK�r��p���uf�r�V�����Y��AФSی9ZQ�����OZ���(CVL
#%n䒚+4�p�"c]Ó)�asI�,sfK�$�vfG�nX6A��f��r�꼁����b��ܞF,���i�g��TbJ�Hv�����R����kx��^��F����
C	�i�NU)bn{W`e��7+!Әݦ��HI�ƪ{K)cȰ�D4e�h���D�+,-�O��.�Z��z�١/`��<iP����K�oA{H�2���j�cL�ރy8�;R��̫,�Ȥ{iw��"����2�J��9!kК+f�K�4�n����R�h���,�^C�G��]*E:�m8�@l�5i�j�M]��o��o,fa���uǫ�0�x��hR�V��-	{R'[�j��-UM�C4�h3q�X2��V�.&j�������yW��M�F*A��+6��N!��Hf��f�'s+bh:��;s#��;ۼ~�'r��%�5�Z���v3�i[��ff�Ui�ċ�ssT�
ե�m��d&�z�͂,���kQ���VƑz����7(H�
��5��ϳ.#�a��}rEۨ�M'jĠ��t2iE\�Fe�͕.e�����⼔�n��+�E��2����ȶPU���1��ӏsv��	���@�ЊZ�2h.�K�PsQ��"�ƱіO�@��;%��9h���p��xr����b#*Y���0�6G�yޭ^��[hݷ��������Q<	�&������8���R�l��r���P]
��B̯A&��ܲ�Tۼ�cQ�lQ�sv����yu{����k(I�������ne")�]���ע�L��Zv�I�I�8m�UE�[�ެ��}+V�CtQ��-wW'��%��m܀�ř��̩BX���9�'T6���A��sA�xl�YUZ�u�6i#O7�Vu䚪ر��ݓ�æ#
���/�7q����n���\b���hc-$�$&�B����w5CB��6*�Z�F��YPae�d�-d���sf�iX%�5$��F���k�ؑ��1�9���.�Xq6��4Z²&�ٙv���B�P��D��t�ː�$�<�w�n�z�M6��8(�_r�`���(s���$�'��3CV������Q`кW.�K����*�@m�I7��<z�>[H>t)3�u8�^�����b,����͂�u�ޔ��u-�1�9��2�z{!��0�K�jF+oۑ�n�v�h�0���k,�鞕�Q�}ƚ}��m'��i���˄����ҍ��76��+64��K�}�1A�%���v���#F�,<�����������a�4�1KFN�kZ�11�:�*��Q�^^�'r
rݕM-oB�G�Ro�fmՓ��=����B��ܬūC޵q\�&��r��4
�`��z�m,7 �#�T�nq����x�4Z�4n��h���^��mm��P�T��P���ED�N��B���G6՜N]�Y���+{�@S=����/�3��H�qx�r��V�+��8��+0ڶ���1\�Q8k��=�=4��䠩�zc�Y�A��aB�P��d�4��P�!ij��Mr�2#U�d�� 1��k���5{ni�7G��Tn8D��i4[�콨�M
��%G�d��w�A�%�r	��j�Li�<)*,��<�,�)@���;FS����9�E�6�j97�G��2�Z˸��E���sj�yT]�S�AG.%���2(�Ѳ��S��
6 Ϣ�TK\��uB'p?�B�1ebI��ܵ�;Y�,8_�V[9��{��k�a��2�Yt6ٹ�+F��r��m��Ǥ�Yu�׊�E&���N*-����f����X�/I�m�P�+�"
�4bh�-����{%-��,��k��_s��u"���8�5�w�9��h��UR�V��{z���Ջ2�ʌV�f��[ʂX71�����<$����{xĚ�?M��+������[gw@�S�g+�B�ҭ�����-��xU]���O�1G.��9�:��M;�@�"�.�T��a�b;Ȥ�"���%�v�����w�>���N|��*��J����`����X �w�yu\���^n�
�U4	B%1����/a�䋻�T��J���J�w�3��5q�	Z��b���aH���Ó�*�bn�Z\�i0v#�כ98�'���t���A��@��n�wM<��z��ٹ8�]J���B«pXUd��Kh�gۏ�g0mڷ͘A�zi5GD�CFeX�{�h����vGO)�uLg���RO�AJ�D��m�w�ޜ���$�y���Vps�#y�"��\hV�񦅕�ػl�GHF�Z/�aךqtʒ��j�Yc_;K弈��\FZ�$m<<�
܈�R~������g��TE\x�-�}_'�^�ӆ�%��0S�yi�����q�n�s�(M�|�tId�q��bp�F��1���9���ⳃRG!��6�v[�\6E-�׫Y�$�Ŋ��F���aj=Xi_k�u�m�fڸa���
�ku�1��k0��;���ȧzEbu$�78b���]�q$m��E���;��ga���E��5yl\�pڼ��]&��o]+��Ó*��$�+!Z�[o��_cH}1�=�O��uu�g&����;s7G��h����t
I�!�g���5��S�w�sCx�������	�����Z��)u��0�üB��Na��=IK�ҧ��M_R ��i��\����t���^4�a/d�#ۓ�7N��e�KA�	����� �N�A4��C�w���TU"��r��r�#�s����~���h���t>�2��!�M`�M�e(���У��"�?�>�����頋o��PA�~a�E��^�w��33333.�=롁O2�TX��ʤJbշ0��E���36��茶Q���i�������ub�쮶�<�"v��F�f���0^�.�J�]��
�9a�Mۃ(�ꛉ����۾[��p>����}�����ol�]�; ��vi�P^�Ǹz+\���-�s74�o�]hR=e�ܢ�����y��JF|��Ζa�j�fPy��+�)A��\����r�t�f&^P�N�4���`�Ո_Q���tL+�`GB�8Dӻ�H�9nn�h;[Wy��c�vmx���l�Ib�p��'j�'.	�S�8��R�x,1�>du�t	�Y�ovS�����٥<�;9
��;n��Uֺ[��]���°�t��h��Gx�ꊂݍ�����s���Έ�f�)󈎛��۝���z+����/���*�"ȼ�@j�[|�qa�P��M�b�0�:��Č/��&�Tb�!�7o�!΄L��i����q�6;�ŇJ�f5�G�Ş�\�xHi9�24�h�d5|/Lݗ���(u΍(�s6��&�x�����לkCn�ee���.s+��Y�L���u�Hnɍ0��N�
�`N�4�\�pd����u}�K�z�����_N�prx;˭ҶЗ`�J�N��w�J�2�δ(R�a.�yW�eE���Tey/���p�K��Pg�:�2u��}��S���/wm�3��M�Z��;����mn
���y�����G��Zw�+OX+c|�����Q<�����5���ӯ�9d��d��l垂q��螴����&�Y&�!�2�S��wB����i�r���������v�aC5�i���y��݃Û[u�h�ʔ�n>�V֙�kv["�
�]n�Ǥ���>��ͺ}���i����̔s4��h���+ZZ�r%�@kf�]p�zt�u��s].A[3*���x4b	X�4mgQ�gj:��ue:�{ս�p�i񋂓���ѺZ����2��	��p��-��t�7x��=�1�xgf_e�fL�8�I���q�w;t3����7o��wRвl��ގu���Z;�[6�fѽ�,���7�/�[�C;kqU�AdWk^�;H�"ӇS��m�vŊ�v�.�;��{���]�0�l5��}����D�Zӭ�|n�c��u��cC������4AK��Zy�E(�76��M4�;&ԛ���9]��kܓ�qo�=Eԏ��f&hmK�q�3�*m�N�a�l���ѤA�ײR���j���27u�Ɔ�V�g<=a@K��S��h�n���A)���ep�G�����܏6�jb�|ՓWt�Ucr�HM�r�UDsf멢���q��c�p�һ�K��YVkx.{�S��dbgon�4;R	D�V_`QԳY�a���k�h��������^a��4�����)�\d��(���6�{xt�.���ct�MTv�P�?Ll[Y��������b9œ�k�D�hN�1�GNӝ������V��b�q��&g.��FѤ*_4,��۩e���5���a����ZeL+$��Zq<]L�f�|�bV��U�-�r�k�Mۼ�ڰ�� @ܦ�e�Pz�� 9w�3(��XWNɺw@�Nw	��	t���{��9�Me�n��v;cr�(v��ޫ'΍Jp��Y�|S+iN88.��ka��5��z�ɹ�Ӎ�79p�u�K+d�5[qoMA��0�Z.�W�맜�}5iن���T�A�޸�y�}��,���us���ԕ�����	��+�c�(gKs�v)ٗ���p���j��R���կ�/�s�s�Nm���KSX��8�hu1�up	c\p����z�P2�j͒�{���UӖՑ4ͧ\��0?gq�����kF�{ ��ʐr)�b�yz;`t,>Ф�����N�O�Q-݂,�o��5ݻ�=`N���wo���I'��wf� ���νW��
�����Y��u�s���h���Z��yJo;��kJ��ɹlM�Y��Ẍ́\�,��#0�k�Qypâ�l��ʖ�UD�n��n�j��x�)�.�]��/cUEٗtsn�o�K{��.�o3�-�WG����2L��Lnj��j�r�芡����f�@����>ے��n�����B���9n7�v��]v.y�he,��(7B }Wg�q�yH#̹I�fg��&:��t{o�2�[�Eu`�n�R�f�3���%�L�΢����7!�QZj�fX��қ/ �Q����2��i�Ș�Ѷ�A�8ktt7w0�#��ZI��'V���-�Ļ���n�1�s���7��i���#2�u��Н���L��^�ݸ�)������W��*�o�������F[�b��w2��v-;��K=�5"g
^����m/ÜN66;�9�8�82V�B�L�qk:�9mH,tK��U��s���c�)��
=��KS��B���r�Ϥ���o\k9H�z�v+��gF�S3u�˲k�pǝ�A	��B8���c��7�t�&h�Z��#ث�3MIk�z�[�̂ub �tq�v�㗪�ɭ2����VF�4�^<V�1�������]���c/���we����mVT�U���hɔ/�cBv��A�$���Ή���މ,ˊޮ�9E�Gy��y���8,�L�ָT�FOv[ ����40���v��{\��x��6�a�ܼ"d�����T��>9��\�������Yk��l'M-_f��Ӎ�ts�&��Z%�ȷ34[p�c���k��'a��(7���s���T�s�������s'm���[Q���%B���T�/�;q�Lv��K�h�w7�\�PՕ4L*�i|�W�-J�|YG�h�Y̭x�l�ht�:��/�Ma�W$�:.�7�f�@�ʩ�����W����FT:��=���ę���L��J���h�w�­�4l���f���34�*@���Rk���v�9ű�e�b�˶Ivs���f��Cb5�J��{-,�8к�r��]`7�=p3��S��z���g�$���J6j䖴X�]Yo�p�m�.�9S�R�cg���'i��F2��'����kMu���K��K�.ю�p�P���o��\��*^ѿY4��{eL�;~i��H�_.��ՙ����h�έ�&�`�5X�"}nef�����3-���Mu�P����]�ذ�Vr�$�,Cǖ]I-Ѧ6s��W��V�,��I����R�}��0��y"f����x�uJ�sfࡌS#:@��Z��N;\��jaz��*�h�Z�&"[}xp�6�ENK.C/�W*[5�[R�P0�v�j�-���X��*LwoJ*ogY�<�U0Zތ���:�����Ge���IY�2��;���.��@�M���MҖZ�bZQ�+�2�6h�ຝ�?L��.�3�FT�j������̺h&ތ�R�Qg`���I/���������AfK�&�A��,�@�W[�q��WQ���<��U��tX��	�l�RoP��n�XG��l��u�J&�����M�wx��"��I�M�������r�𠌕%
���|��b�=�a�R��}�	�+��᧸-�`sa��v�Dg^��K@��m���Uv�U�召�����欫�)8e�w��G�J��k
�R�,����Zx��#�Ci��ZFV؛�zԼ��!��fY�e��c4��Lv5F�����)�u9p\UG�u�_q��IT�H�Du�fҹ����z�:��ӡ���;����k�y��%ݻ������6�n��9���ntV����󂺰��O6#�e f��6�J����h�S<p��9��%����0s���۹�\�R��U�:�X�Q�aMm'Ob#O������|d���
���*���Y�t&���
�c{��؎m��f)6�������f�Yǃ_3w2�a��U���r<.�ץ��e,���"�.f���	n�w�S���2o`���qs����&�Y��4K�M>�x��`���K�Co/�]d�M�ٻ�_J�� ��avƋ��f,*�&��T�[�W�n2�V݆ΊL��]�=�����P�FL�����ukuS�D����8j�������[�|�}۷6v3K�����o��Ɠ�շ�7���<�o�*��̳'N
�n�Tս��`1Z��m>i�j��Lns��Qf����ף0�:+�J����C35���s\-��"��Ok���n����Xi�Y�]���]�hz�G;b� ޾��+J�o��H"!9=���.;��XKr�r:��^-mQ�֑���6�!k�ܤ��Ut�i�<��'Ѝm�T�°�2gomG�]�냮n6�Qf���k��-���U�p�L�Ls�ݓ����A�@	:6*�h�*j����F�I�w^M���R7$�D��3w��F`fƚ�j��*� ��EM����n�8�OM���=���;euk����Pަ	x�V���Z� ��8�����Ӹ���=�]\EYD�xM�y1nJu�D�ܾ{��syP��\�{(�Hik���f�t{�3�c�d��ⷙ<���}x����v��6��E[���"�i�J
���>	����$v�(��J�l%{�xĐ١�臧�!83|��iQ��kK��gSժ� �Fuv�ۗ&�����s��j�'U�Felќ�>=+�
Y�0f�7�z�8�&z봌0KK���ڮ�l�®[\�,'8st%s1)�.L����Qp����u��32��X;{z0�nnb�}'jw;��c�Jqu���J˒wa�v>��sd��,l�k�gN/.�7�d�s�����u;�_Ʈ�Q�β�v�")"��Ý�e�:F󋆅%�TF&����ë��N�w-gY�B�R�o��{�������X]Q����k�����������*GM��N���o��n;R]r��u�淺\;mŠ>G�o�<���G��JG�3%'61'�i�s������H�W�t]�dM�ຯ\�;�G{���{1k�6t.��wwwt��������������9�k4�u�^�`��*��W'���c�م2�N)�R�u!�-���Ǝ�b3�Z�:�ԅF�n4ږ��֪bbh�$ɪi�C"ta�B�)ˌB����#l�zLd2��eT�AtȆ3�$1����DV%%��� d�I�p�U3^�2�0*�
�j-��1�váV\%�>�*���
��|�sj�[�̺��J��]9jQzj5��A��sч�G�1�}��ل�@�-& D�\��
R0��}0�d�@;
X4ˁ���q����n繛B�M��a'ܔ�>����E�V:	H �n d6`��`Ҷ`m�&�������?��A򻉂�VB�7�{,>)��э���U�Bf�H�a���a��Xp��N�N*�����RB�1.6ԭ�L5��%�6"%�F�2"N0���I�%4^���p6�x������"�i�n,��Ai�L-y�H���e4���Fɖ�.���	D�Z@��F_\M���c���B��
i�(T�HM��7v��=ID�uM8��I������A���̆�m)��#�^I(��Fڀ2b��)eݔ���7�	8���*(��j���j�nl��׋q�	M �q\EH2�i�DK���JF��Ø�ؘr�&m\.��s6n5�y���M޹s�xV�.��Ҩ�b�Lܦ8Ko�܁FT�C������ʖL*-�F�j-��v�Ѷ�%V�WJ8���@�`�����pj�c1�R@�-���DB�0�2�m�/@jZ2���U��72�a��;��(YF�E�'F�T���B�n4ڍ�Q����g��N4Vͺ�8��a��S��I�!I͖Lˇ�F�#!b�M�\�y�� �)��8g���J&l0I�ù���]��9�y��2fKTM�p�Q��/Ҟ�Ȥ
7-������&�hJ
4#���9�i��	#���3j-Wx�^f2����j���oG%��5����V,�R& �p��T�"��%��X$C�S$Ѧ�QZ1(�t�$�`�8�H2�jېI#1"�mC>�EP��8���e�a��Xp��	�i24�?*��(|PE3q�6�1h�i+7��_R����HPPC��Er��0C��%�YAyN% dD��/����I!!?�������	O�����33 ��30��ٿ�o�鏓����n�zt�C�5����
�@ަy\��31�5L^��;D%:P)ڮ�0 M25�y�m��`�8����)���4���/ �/�ԫjă/�����-���WX3��w�fn�C����N�Sg����wS�����R;�Nթ�n<��i
�����wsVwW�j���&������R���&�-��Q�3
!hE�ܰ`��9vӠTx�?f<�^v^q}�YX�d c���h�e	����ȷ]2��� T���eS6%rr��y}s�4 �u62���v	������z��P�!l_�U�x)�6^��~{��6)��خ��G�pa�Xt޳J�9�H��N�������w�� 5�5" n�m������0fƻ����֦e�����{e`G�tõ��ˇ���,W1���v��y�55zS��l�f����c{��n�*�-���+v�3q�
���]���z*��7;��7|��e]XkIVn�T��/�ia�]������qb=L'�k���A�tpٴT<��}��g�߯Y���l��Y���l���ff}33=fff}�333홞�33�������33홟������333334ffffg�+3333?YY�����������fx���϶fz�������̬���Vfeffff~3<ffg333陙���Ϧfg���϶�����fg����ff}333>���������љ���9�϶ffs33>�������������Y������Ow����y��^Ǫwn��n�V�c���L��5���S��5��U!�K���Nvŵa�WS����������<ԫ�YhT��(���+��Q���ˤn�����c�u�(0x��WONj3F��`�4��;x�i>z�����	��,u�7�N&�6���)��7�����l���_N��EG\�ȉ���j��B����Ŵgg\�e��� =#�p�l�^1L9B�Ie��.�ȵ�A��;��Q]\�hk���n�7��ї�eBhB[6�v[0���iS�оǼ�G7��a�Il�6�t������cWvےM�4��Rf�*�m�������T��8Ɋ��4��U�"9gK�0��ڵ���xq����Jd]�����枋�4���U2IM�fKԫ�{PI�2�O�bS7��7*�,�Pm�F���3rˣ��;o��(+��'�sn`��g;8���ol�Rf��^b��^kO*���a<�v�R��kHʹ��`��v,�V�0��5�6���w�kG�b��y��o������'}���z����홙�l���������fff}�3�fffg�3�ffff~��333?�33=fff}�+3333����Y�33?��333?333334fffffh�����љ��������Ϧfg33�fff~4ffffg�+333>ٙ�3����l���������efffffVfffg�3�fffg�3�ffs33>���������Y�����������љ�����������g����p�{9�	�����vǅI��V_'�U�ٷT�7q��:���EP�:og6�r���-�}il=^:7r����M�XA��C�����E�8�m��<F�e��u4cV��0t��*�5LGi��G	]���2��;�ڭx@��7w�:�ݲ���܄ag����Glr�F���ɨ��B^�7��� m�\����#7����R~��[q��k3�����2��M����0�`�h<��A�	U����R���b�/�La���m��ؼ�-�/Nۮ����/�2�ص���󶦍����S��To6n�� ��s����-R1N�]MT�[L��F�A�����F���H���X�U�c������͡KHX���k�jWV�MwB^�>��ٱP^�ݓ��=`�[�޽b"{����v4n��H����K���1�1�e�s2�]�<�����2m���8Ѯo6��<����(ݽ�^ɻ�%��(o<jh�{Xx[���+,$F*��&̴yV!���E��&0.bc�.�*�����1��9��Zm�JR/Q�?/_�z{}��w�����Vfffff�����������333334ffffg�+333陙���Y���l��Ϧfg333���������L��g�3�ffg�3<fffg�2�333?Z3333?�333����������љ�����3333?YY������Y���>����������љ����������fg����z����������񙙙���񙙙�������337��K��b=ݻ�]Cخ-�Q}�U���=�G�n��|�T��p�B)6�+�8�9�!r]Z$L��5`Q�{�8���w�ƴ;�:΁ �&���;m��U���82+6��X��ՙӍ�_��e��uݚ�k|g���Ez����	c���ZR��>,�
DwK.��)��6��[�pJ��z���6�ꆆ�W(���`�O`q�pazؙ)"^������%���@���zh��k����Ku�@�(jJB���Qe������);�%��K���	R���s�V�
K�(ZB�,u���4;HA@�mr{��sx�[��Z9��s�Z��+��x��)���5��4*m�Tn�F��w5eA9tvPK9�<�iVm'�B�ij��r�(툆����Oq蕘%�~ ���A�;���5ƸC�7�ډ��6	A�C@�	�� ��*����6@m>��P��s�go�f`�9ڛk:�J��nJF���z������
u+&s��k� ��.�<����CW��������;��y{���=���~�33?Z3333333�fff~3+3333����333홞3333�3333��333>ٙ�3333?YY������Y���L��fffg�3=fff}339���>�����effff~�fffg�3=fff}339���333�Y���������������ffs3<fffg�33�g�3=}�ffff~3<ffg9�s32�333?Y������ffg333陞33;���{���/w���=6hL�:i6��2�i�fD�=�a��橪��y�!!��܏�����:�R��< ���/�2���0�0��,+E
6�>��8��`������}q�N[s��wk��`��p6��9yq�^�:I���x<=x�خ�ޑ��Px*����+�gu ���]��_-J$/��
���#t�]$�����m��aj�MRᇕ[���V�Mdf(�������0����^�'�nv<���i�Nj��#81�e�I]+�jY� �n��t��0j�-�6�IF��>g��4���ro����M>}6!�M�ƪ�r���E�7s����6kw�EhTü�}�U>���s�j��\��m;2�jKT�B�r�{�t�㸒�+;'@�j���u�S����M\�%��h�%:&K7weA����B���^q��1.�{�����^MoP̢Ӧ�s4�TlgC{\�ڗj�숴���DH\���B�v�������n������4t]=۱t瞍�9�&��)���v�lxf�BM��[M�Ǳ��V1���״L]��r\Y�좝L�8<��wr�|	��cE���%tdvQ#"> �Q�
��_5�^��@9t���m��h*-����M�AF�e_I�f����5�8��&#&s�{��'��Jٔh�N!�2��f�y��4xt,0�O{��t�A'}q��u�;W��c�I�&�A�sj�*岟A,�k�h&
i�{��j��ͪ�#7�4w{��SvT�:���r�9/�NE��O2�{t:�"D˅�!&5�q������ EgA�+�j��L�ֆ���׾�;�4D �C��B��#L�����vw�αj�P�t�c���Z�*���щ��B�L#���ʝ-ULTo�Me���8�f?P��ӑ�9v��Ȝ�1$x[�R��AY\C���Z7��G!�֯Y���O'.�Ӑ u`�A�TwB�<��<�wQEN.�Zn;��("�<��-뫹7q���3�����qۼ�'VT'o�M�0�_���(s��Q��͐�7s�e#`p�A�c�	NK�o��]w3 ���F�5�s2s��Ʃt�$ஏ���}9�s��-�	��+���VCOi��;vTRV2����J;�H��v?x!�}���l���9S��MB%�Z��9][`q�B��$�&9r�׀32�Y�Nd�_7�{�i��"��OѓE,%�W��Bɝv9n�K�xN{����������eQ#��^����saUP�9]`#ޖ��e!�uݮ��>������uq�Y���>�w8תG�r\@��̔�Ff�tV�޾]H�t�a��fT:�^׵�e%g,�m>�u�}�_���»5ޓ�"E���	�e�s	��m�Cf��4�;g�- <;%���GXm�i�B�E��7�m]���;��K�Rޅ��ؖ���:��K�^���,�.�fq��m�n��N�-����q�C�X)�v�I�'*� ��c{���f2���7� %�ԓJ
��df�7T�Y�T�wg��,�閇��m���5���S[on&��d��bf�/��L.&�L�v�����@xgb½��'o9��m��бЫ���ll �����+t�+��w��+�4$����c��ö2�"��}��նK7��.U�=�L���,Y�gS3T�5BR�/�9�od[��<�=��$s�c���9�N4��|�=T�ܝ��6Ry�`C�$ֺ��A4���h��Ś�Kb}$�U��t_T�����f� �ˎ�:�bڄ:Vi���� ��^�ם	��9�X��xL�c���|�ES�j��!!�<ԥ���ug`���Z�ʾ��7��`fjړ�X3��yݽY�y,���g`Y���N[�E�=�>��=��D�Hl[�w���t烆���o��ʍ97J�蹝6�{^WPI0,�/��7�Q�F�"��\��m���7sʌ�$ⱉˈ��}�86��e�li�ܲqLW�y���@�W ����>�zt����WY��dag��Wo��x�H%μi9�y��^�>dI�r��cyf��p�HcF�q�6�;y/P����Sehj�֣Il���n�پ!)��ӝs�-@#j���04��X�誋��B�83�|1��wH�Bǆq{z��:��Ķ]rY��I��[aͮ&���<���dU�*ÿ=�z'.�ȅ�u�{8jx�J�;�N����,t����1�rJ3�s�}֌�w�:��#��_K�]ur� �k�a���.e�U���N�pӽ�ӧ!}L(���dٓ/I��:�����Ļ�:ǐ���K �E����7�]x.�z��+}8��^U�amq�kZ��<�m�=.M�6�_u۬'?	�z6Ŷ**��_u:���������.��9����!�R��57��M��i��:VW��Wko6�C-hk7
��z;��@�Y�!�F�I�l�2�v7�Vo^�D��Ep�o���-����A�z&�~�N�!%c�ھr�Ws��Ѹq���z�8�s$��g*�{)�}��Zӕ*��β�n�Is6��ΐ)���(L�\���R|�J"X*R���y�Hkh]Ta<��q�� !����< ��<�4y�F��F�=��8k���[��l��Kv�g�P���{i��]٨����X��ݦS�4�\���u�C���hʰy����w�Z>dK���.��!mfE)���,��<}�𕧩�P�M�oy鵖��-��Χl�k��>��ξ��[qmؽ��lTh5�^�"Yx-�`x��Ѐ.���)2�m��3�<�1��6�3��7Ŋ���톇��]�$v�]}��[�6V��o���{�&���92��t�L9k�ޕ��|M&��*�s\���+UGq��I��c��:�.°��N�ޑ��]ٖ2��b�9��gu�N�\���*b�z�ΑRj��j��*V��/}�!��GU���h.��[\*7e�⥊]!07�a�Y�̛�O>�	��rCeѷi�H��Aݯ�Z�v��K< �;���.�Ă��Y�S3���عw��x���3x�(��l���3�Wv��W�\�#.4P�����W�8,�`̴�3�C�:��lB+��x�AdΘ��k�������
���&�p[j�W���9�Y��Z���왖�֣�.s�[�I��}W���b�lo�����8������&����Qu�|{%s�r��sc�7w�W��Q��u�p��*�����?U;ɑ �v�5�Y���p��4b���th\[T��j�ڱ�I�8�U����-mq�͡I�$�X��c�s�+�OS���_�ݍ�®��V���DڒL�3^��d��a9�2���{�-��L����hvs���S	���C���v`��2�Ö�c��7�CVc}5W��R�ń����x��KBM���Ր����~�~o��������	$�l���>����Y�����>�������4�Q��M���UF��DC?�� HN~QG�D����V��O�7�+))Dd
!5�e� ���P&Z��O�P�y��u$��BG T��&�z"���[���q�`��a�Nap��#B�+;G)C�_E>_X��ȅwJ)�,��V��pGn5����QQ�o��ȥ`r�{�;7[}�g>����J~8,�Z�����ĆjUx��AE�B-�Rw%Y�3�#&�TS��ת���O���	LGǎAw�u7;��N��t�MoWE��[�����̛���VsrY[Qo/;/{����wu�U6nJ�c!gɎ8�W��=ݒ�v�-��-���pU��������懯6���Z�b��n�HZ����/zu��N���͘���v1��y�h��Iy�6_-{��ҨS��;	W��Uܩ�.;Fަ.���Z��r&U_��+;OX����fK[{�\]{ء�UK���4d�F��npu��Gu)kh]K+z@�kv�*��N��3s��q�ӱ�7��9���wV�L૰G����>׽�^���]�eM�X�4�M\�5٨�Ja��9�d��3*�(�/7{���õ���_S%���t���c�q�έn�>=���k���Ż�ڻ�p{ʟN��j�nIt� ����P�"���UmA�'�E��aax�E���,R��8:�W3MR�i��tS@�כ	�L�#�BCP*(&����$ф�T/ɱDG6$j-5D��"��4�,��J8���*2!�#"��f	%�������i��q8��q�P���"��z[�&B�� �GΩ�-4�L$TF6��	(��i$�mT�79U�Yr��k��9���v�8ѽf�h׎`�MWx���Am�5(��3
[�YT.2�"�g��rؕl�`�u�z��g�?Z333334ffg9�s?��,��_l��g��\k��+�N4�^:1cVF����Q��S�Dq=�fOg�����fVfffg�Fffs�͛=��#�)m=�FcQA8�2ж�(#%j[KV��Yj�e��e�*�z���g�2�333?Z333��9�}�TA|�96���*�Q�*��b����Q�f��E\��=��\��3홟�������h���s��~|����}�/��$�f��L��qZ��ک*��aDD˒L����d2�V�ɊaJR�B֕��dr��K|L��c�Q��2@�l���Y��dpl��X��c*���TE�����33$X �H֖\�bX �F���1�� ��(�
8�Ud���-Q������R�(ʄU$��.f 
c��$5ԑk�nG�B�8��D�Um�@
�Ad�"YZ�
�R��\HC�[R����La-)i@ ���]�A�E��R�[)� ��JH�1Lˌ\hA2�űYI�X��6���
P�/�hc^����Bȱa�d�2fS=���D�i�"%jX���R�UԷ��Y��ض�;�Q���lf`�5,)k[nV�A���=]-���l�as28R˘�,��3�ݦ�Y."�a�-���iq;eQ1� ;M�P�E5�%,��g{qUX��t��D��*�i�m4�S '8�r���1h������2�r�]W2��L���[��O�n����'!��ٕ���`/�ͯ���
'>��_�/b��fz��.sm��K2���J`�j��CQ �I���C,��3�dA�1�L��T�^4��9�Κ�J\˖��^����#�O9>�U�sb�Yf�y/;�ϟvQGt�I{���;��'�ɼ�2�A�0/>)"��~��4/��`��&U��V�d�ܧӷ�x��9q��G�� �9S�o{�҃[��;{,ɥ��|��m��D��2��d/}N�X�����o��~q��/Kݑϯs�>��nm��Z���x�}��,E1���#UK�毶n��Gyw�{�;��6\��u�1��2���	&
A�:<K{�}7�������vo�>��ރ�}Ҵߨv�N(����"}����so��V:w�u���~�c��u�I�~.V�߄+�N!R
�}�ԓ��9!�0S�Y	���� ��>��� �nE�~ﺧN�\����2��Iϥ]m����{;���}]�� �0�̾���+���j��,��2L��㍼o1��q�'�QO!=���S4[�����B<�k�Ve|�|���B����QDO_�c�US�/ �AB�n>�>f��B[��Ϯ�J��k�1�T�2�o�#�����#JX����ʳ�qu�y?O
���X�,@�z���Ȣ��Ǭm�d�'r�̽���_�ߟ�1���^H����ɏ��]��<�Eu��K���y�s���6�k�������&�z}�j_3�1l틯ZҊh���L}�b�9�߾��|7z�Jz:}wC���x���8�w��R*���+9t���!��L��s���,��N܇�p6	 �Gac���@vp�ع^]i��߳s��<f��0F�������\���/��{��5w�ݹ�[��}�|�h�B�m0W��G֓tT�������|��}����x=^�ؚ�y-'�}����IKU��\����r���N��A`�w�b͏{����:���ޟ+O�V~��F���J����]�1J�ʊ��Y�75^��DW��j7*��sޭ�,�>r{BK��(}{:������O�XPR�/���V}8S֜Y��틑��=Q��t�o)�d;��tm����Շȁ��O�����E%>o_ï"7���ާ}([�wjΚ&$�-�8M߮�s�T��OZ��� W��T��`�۷���Z������=��}�|:�>�JG��$	�W���N�'����ȈY�d��0[��܏^��rH2}>�7�.��-}7m�Mq�����%�y}���9=�}�S�bns�����E��g����>����P�mRƁ򰁥�g���{~���or�}3��2�\9��;�IkC�a#�&�'`��3V{�2��]~TY�����m+������}n�+�>[���w�CS�O���&3�m�? � U
�k~�s�x)r��R�O����)c��K������z$e���o5�c�\�e��W_}{[�؅)��gT�z���W�_|��~�b9��}t�rA`�~��I9�ɱ���37N�=99�����]zY��A��ă�f�u�<{h7���3�yyu��&W�R��j��.�,��޽U�*e��<qd�$ne���o6�����Q�s����	 fieB�Ҕ�X��*SX�yg���*�U�]�O��]��Ӿ�m��߃�q��;��f�ĺѩ'j�;�}��t�>�g�|<<=�
��^Kr_\��³�h)���tLK��o��9�息�.��']��W�|f͹.IiP����C�]V�J�X�6��g�8 ޳���	����Ȃ$i�����R v�g}��I�e�ʁK�y{���ӗ)�>�3����}�>��)��|����1�8��Y�?�VMϾ����9�_��(���۞����}�,O���MV�jH׈��G�����C^y������R��}��}�/�� =Eyo_N]�u��y������$���_�{<Ľ������D#���X�~��m�'p;���[,}A�{yM���~v%o�Ŀ��J!�N�7nFihbվ#.s폚j��*�
_�=�}|(?����7/۝��T��҃4|(?C�U��j���N������ף]LO�|�v�NS���w�
m�Q�S�m8
o�w�� �v���{>��د�q(�RG�����<�'6����@`v���z��7��>{��u�H,�B%�'U�d��	�A��J�]�+H���f
Y~%�5f�筺=�̷Ws/�����w˰C��hEf�<�_���}|̞}�a�i�A;��Fr
Ĩ$@���b��T�nh:�cL.�6�K�S��sc�;u4jO#�bI<�0L=u[���ieDڄF�&�!O@k�����$���#Ѧ��w,�X=�~���~�Z7� ѓ�"�'o�٭o�ͤ�=%'B}~1uC�0�d���K�K��ҽ8d�9�ܬT��ݧ�@��kd�dYc���ا6��©؉@�n��6��@���(�!X�jѢ[~�7������lֵ��b� �o���o���}�b�Z��clM���~��.�;'^������WﯶwuIo�^�s'��~���U�S�������}���C>?J{�Z�bTP[�����]:d����MuB��{����f�]�;��Չe�V�bg��/x}��թ��W���^:��h�G��4�}NF����7�{{�@���DQ�э1[ zK��'�sk��|`�w6�9�P�D�w��X������x;�����dϾ7Z ���_W��Crڢ�} ���d�!�տ=f�a��}��7[os�p� ľ�pE�O[(��y�8�[�e	����[�~v�ʎue(�]1�7[瓵����#.We�}�lK�j7�6ס��.���罊u:�� �s2��_��M�/s ʰ�e�mFT����қ-�3��ړ�d��e�m��y�� ���X����Z�Z��n��v�v��4��zy�F۾��{�x�m
��)��k'b��s�@���*��V��-����çgy�@���݁^�����i��R�嚧����|v��������p��:��M�`���P�_�_�o�ٽC�O���rߤǵ�� �/�
y{������ZG����f�4�Q�ݔ����ƿ�:�aSt�� W��'�6]{�����=���{�x�o)�����w���s�}缾R�MO_���<x]� �_}�T�ϸ�+���1G7���_%��p] ������u���]�	O��BU܌�}�]���dL��ā�W����ϵWg�qp{�{<���Wd;��ɫ3��ߝ�4�H�Q��Z��W7��!��M��&<�٥EU��q��r�.�����t��L>n�4i;�I$-�ү�ַ!��h�V.�OT�xxg��������w��f�oY�}�N����G�MGAf���Q	+�U�^��� Q�>������_��^N��w�,��#����?���٩��7������<N}�o����r�h��}2��y�������׋����z}[���ہ�ol7��]��Y�2�k�+`��^�����A�(�D)�O����&�ݯ_�r�j�����j��L���?k�~��Z����V]���<"����*��~��:��,���s��vi��o��y"FP73�$���ר��@�>��{[q������~p�@v�m�?is㚁T�.���`+�k��z\���y�7%������~t]4=���WҦ�����wfm'hq�����ҽ=�}�~��^[~���N�|*�U�S���O�n�)q�)s�jU.����3x']l��N���b\������3q�Ke��@¹�Ō���)�zv�����h�tah�f��"���14e�-Xpf×u���e�Ƿ���x�|||@> x��{�˅�9ϦK$���;#ƺ�6�o�W��ԧ�}����� pt�(oTg���cd��s�>�C-�p�c�L�UP!Y�2/<eN����l#�X���X�b��^���Ŧ1�������� 
���E/?��+{q��w%OUR\����WϗRs���?z^�l�ϣ���h���O�png��!�F�@��c�ܻ	�5xg�	p��ܡo���o��9{|m{7�ӊU6>6�Z��n�2�|��g�K>&��fAu:�C�z����ﻧ�꓾?z�۪�K-�3� ���տ,�B���)���>�Z#�����{X�A�Y�}�����[�ۺ�>u^P��࿫�5O��?Q��J���C������/�Ȣ:�+F[�yk�1�#c�,x]��]J�S���j�._A8
v,�X&+�{̘�e��ֹH��m�9�Ɋ!I���r+w��a�%)RG���`���Ū>���{�;�h�tαD�+�͙��V�%
k4�H�%mQ��ɷ4[m1���n:�[���S2��6򛙹�Wq�M��X�1� ��S�����tԑB�=��~w����_���}����C��,����S��V����Ϣ�f-ѹ���l�5��fa�����8n���g�DV?xkw�o�3�����jy�V��|�204���`gyPQ�ʿz�(��}�3�{Uh 
��}=^�w�Ua�3��{�����[������s1����w)��w|I>h��!�?}�p�O����<���W8�{�S���*�Zˌ�H�	��4��q��o�~��3�ޣť��w���|$�#��O�'=`�����p���jw}��@ԙ9�2�����wѵ_OGF�WҩC5��.����`���4�}b�ܱ�X]��v��Ă�%�h Fϔ�^�
��h��z6��۷uK��V��w��|�,ݍ&�}�[��AϹy����#V/�}1�n�Xw��w����vZ�&��[��s5��:r�&���ZB8>�~f�,)^�������{��:�?��#�g��.���FK���kq>%2/��"]��P�t�wL��N�3-��v�u���|ÁbA�@c�w[ӻb_d��_�T2�N}K冷�;�%�u|���s�*K��o�H�۵�v����1���[�df�b�T-�����!����Vx,��Ƣ�^�v�	jT�}��#>_8�#]�k��/�w��yn��{=�Z�ٶ���h�*�^����W�� ��~�?��}�y9��_���=����o��
}��O�_Sb���s'��06lk���S�ڥ�_��=�i2q+g.^l���0����!H�I�$��>L���Ꞗ��jɲ��81�����h�7&=l�����wz����m3�Ns�^ƻ� �vJd���{7]ϗ�3�:�$��>�?�����i��й@��f*r�ۇwT7͸�N}��{�w{�~��I ];I"�5z�@h�#i���3 ~�������UW�9��?W�O2 �i���t��n�1hf���|���o�LHf������Xsս�C�����$�YY��m�%��ن2̢�a�	q�w��}�g��l����o��ppX��谴c�2�Jo�d��[�9�QD�t�0���k#8'��u�q�<� Lݸ�H�[��<u|����-AC$���4����.��i�Q��I��+0n]Vd��w���[!l2姊��L"�=�u�GM���l������.ws�ٕ��B5��*�ڂ���:�Vc��|�wN��k��q�mqsos9.5B4��`��M�<{�͘�ox�1v�޽n��k����4��&O�X��G^]��W�+!����V�*2\�Jr����X���������1ܞ�?}���e��q}��0v6�֬�޾7w�����b�R�]����#��J�xv�Br!�¸�mާ��G�:\�ڤ(�CK��j�&N����g6�8JD���*+R�S���c+XVQ�5��4��%��Qa�	%��Za����9�tma���R6:�=��% {���9rb�J-Ln���I�7JtA4�k�� �*0+kh/��I�A�b'c�l&I�Y���hN�f�_d2�����3pv�
���AFp"���[��؎��R�������I4��l��?^�s(�.��&�&���Y6T��\ū�8�Pi��s)�5�ϝ�U�A����
�Am�sg�����}t�ES7`�}7~�<��vU���l}Wmj��S.���^��
�A��vؔmR�%�0��U�J���c�:��g"Nn=�� Z����rghW#��op�6�m-��Y�2̋�g>U�[���;]�0եE^�ڬ��)�٪-|P#͐Wa|�,���l�;�j9����Zvy�w�r��`���2޽��l*0�A����r���s���f������k]0;<v��ӵȌ�4>�z�kΰN>3E.����5n�y��Ӝx�(����%k�6K�N�]���3�`�=L.����|T�e��⇠ci�Pe��=/����]��)��Qd,k}�ηM�nc��R�+AcPx�K����x�=�!���F!���oC�̌�fǠ��jT�{�����6Q+K��(޷�f��T�v[�5�����OV�S+��_K���8��b��!�-��+᳎g7X4�ў�H�I�Pk7��ڝX��Y���k����FD��&z��z�s��w;�k��*����7����e>k�+ջ{���;���I�����w�S���[�Y."㝙������b^��ơZ��mk--�vi�h�r�C�jcE֑��%�<��?��������g����>>>33?Z33=z��>+��Y_�}{���E+�i� s֡�NaZ��"�����ĬD�e�l��g�|~�>><|||||f~4ff�2d���t���`�[e�X�U����KJ�-�eMK�~����=�x�������g�>>>=|||||||~4ffz���|~O�}��Y-��_/y��km�I��UVĨ�
���j�ҥ��m�O?�z����l�������ׯY���~Y����}�y��_s&"[dQDU��*��)iJ�yq:p�,V��U����"�lY���S[��)D�U��5)Tz�T��b�eE1�V&9i���F�K,TDQAZ֣e��°Z�F���
��F�Ȋȋ���a߲�t�z��abD\���*���UA�j"Z�p��A*	r��c�E���ՠ�WY�Rk��
e,x�-h�0�=%_|s��EE+�;����Z��\�P�Ė��9yۻ)WCOwOۻ\-��#���|.�����3���),����X	a�"h�����\Z��\P�(�����s|@�},U��ʂ2s�"���o��fw? >!�ɂ+1��!�����t����_yĖ������	��Ò�^����⦧�:83̐8�������|����?�뉑x��EC[[*�2*r�A��nK*�q��{ng��7ń�ozWڀ&������b!��	�Y���2���L�RҪ��f�����l�_��;>��!-�y"�0��~!'�9�O�0��oJ�>�^�������;�RS�M������v%{)���`{�/iO���k�Y�/�<7�m���ǹ��^����"u��L�|C�J���������}�f)U8��ҷ�37�|G������c��<[㷮ۿ>�z[z �\��n�#�8k�ʰ���=׻�� �WL�[�,���~��=�v-���6T���k���������Q�ǯ�t��{�x3,�i�T�cy�mG��q,���|-� zF&���1i��GhY7��^�@i��Ԯ���3�l���j!�V��@�
�	���:�1^c���(r<�v9�5�3�5\��$�aڋ��y�gr�?^����ޱ\��2Є7��m|��6~;O��-�p��ϏȀB>Dx&pn���y�}��&�:s�B�ƕ�\�o*��%��atL\TNm�X�V��*6���y֟��� R2Ƒ�4�����o�;�W3, ��_�㞯��.m'˃v����u/�����~����Q<큄z=Y~�w��V]�G�n}�j��ݯOu��2��d���Y!@Ր���,��I�k~f�ߗ��b�g�����|l��/� xxL"�耿G<Ok�!��/��5����z�76�M�"�N�x<O�+oX0���R@������^bމ�h�~�B��<@�)X@͟E�e>�>���IS�W��[��tNgmp`�L8>?��;�=(������D�t0�.��V���h�mU��<Ni��� �}�����c��5���{y��(^�����u=�#�,�@�??P��V� �u�2��oW�c����fu�������&���^4ؘB��@燽?�Dk}�����ĉ"Ob>����{�{l~wWo1������ ��C���I�D�'>vo?�u�4���j��L�}��^-$I��uQs�y���W?|��Y��B�Y�@����1�L����'�{�tX�����v����k�+깯��`8�VS�������,'P,`4-�����ϯ�=oѥx����_�L^!�?�	V���eTw���H=�.,��6�3�E�/��I�R��Wb\��0�Ҫ4��Z0�tt�b]y�ڨ������y����j!w�O�Ywߏ��R<��ë]��.��Q_'�h�J�Of��d����3qH.0��/���|"�IP`�D����4ۆ�9T�\4�~#>�#,e#,��� f�����e����?O�h��n���P$�@8��+���Ě�ϔ�5���
���0j���r�~�<��;��\�cT�XQ'/��Jh�p(í��x�,�% �&MS�Ÿ��f�� �9���z8�H��y���d�ʠ�R�`��d�} YG�T��@q�<���I��>�2����` �*-G�(7��3	$�>n)���p<�Ad'ș>������eG܀�I��b)��{�g!�[�����@a�²�p,�6lo!��`��Vz�/2`X���d^V�ӑ����#�K[@
T�8��5�E��=������G�5�q��f��P��<�>݊��� (�7;�&���e��o#��	�+�x���y�s6⥱�e�(����GЇ�f�/s:80dI].�ÊO�Z8 �S
){ ƻ�Ey�o�i0��>Fxkz���.��]�sL�0��d�a?��D%6�!y���p52�� ��	���@q��3ͳ^��d���h6�Ƀ�<����^+���]��6��2�2�^m�`Y󠃧P'�~�i�����<�������h$��PHO��~��� �A��|a���e�
'��Ӄ���!Ε�3c�\�W�o����'0��=`� �9�RM w�Yx���+���k]@Aǜn�-�-Ŋ��ZƣX����˔l��|ߥ��=���)Ie�#,`g}����������!�3�H�C�\nW���9 xb��b�p�@��wOR�\t>�.o�V�ZIm#�Q���K[�,>J��!�X����8o�������ݾ=���u��t��5��
դ#��t�c�3��0T�-X��&|��_D��Ǝ��7�-/Z���� �c���c��G�ٷ����K�2���7פ7;�|�6���&>r{�{�"
y펟7��{T��ג�����Vk���ǗL;�,�I�K$<yI%���C��v���|s���r@]9��'������30hfl	^��-~�mL�{���	 g-uT�Ł=��c�vY4��A酳\a����{�����
�&����N�N�+�k]�J�������$���:����/���m��>=���q���z��}�������׳������p 4�c���#�Ӣȣ$���N��!�1SUJ�2�z��ם�ןN���f��!�\0�>#s��.���V�h�f�S��9Y}L�ݎ��l��:���z�680�����fx�c�C%FY��~@f���l�o5lC|���x��������Yp�(<p���]���;!�����kw,�e
��G;�e*]�u�B�³6����,V=WJ[�T�h�>��]�
����)���K�wٓk������"���,)���3ǫ2����
i���{�Qe%�RYbHϳ�y������f�u�1�d������:�e�Zq4	�"�O�!3�ݿ�+�ޅ���6���=�{�P9����_���;e��e�(c%dX>��D�ӭ�w��nx#M�����b���\�b�,]��{׈�^�sV��(=ْ�e��D��Q�Hc�~���r0�������!F�b�jx�E�f�eM���vq�p/�ͻAx�a��ޫt؀��`��MXX6��`��5������oM�Csi�o�I(��Re�{�����:@q�°��xkvC���e������������rg��}��|�Y}��3�7�z���| 9�ğ��*�ϾqP�0�����,�Y��������O��JZ@$P3�4�ϸ��P��=�!�=z���E�p��Q�����F�K�Q%�ǟ���e�N�W@x��J�	�����y<&���0�7l7J�'��/��l:Qn��ҳ�"Ȇ�Dg�����W�5���O
G��6׆�,���6^��W.�sw��P��81�i��|7�����lQg.a�xu�
�]M��կr��~ψ�Qd�6RB���nz�����huܘ��s�n���wC�ޟ��z��(s����h�ҘN�85��ҁ�V���ּ�"b<��kx0���T��V�A��Vj��S������]���O�<��V̙&L�	QH*��������������n:s�<�P�9�)��S�7�ig?��8M:��7�n�G����z̽��r��>�mY�P�D�q\�s��h8z�`�=��ìXS��|q�ݞ	Ň#Ġ�j#';ҊM��2IĈ�#�-�d�:\Ϥ\2�OE�gH
Ʉ��G�ۢ��[�
�sʪ���=(��;�w=x�@i,1�slU�s�Ö׮' �"C�y�����7�����<{���<��g�'	zͫ�����,G�Q�����oo��.m :�$�5�q{69d���͊�<fv�*꽡�4Jǻ����L#���u�d�-FRH$�$@�p�{{<��o�D0}WƠh����P�6H:��� �+L���ߐ�vz�iζ��@�6v�� �Ǥ���{;�Y�8����K; ��R_T����r�B��!���M�D�}:neVfw��q���go Ȑe�
L-ʣ�Gm�����W�ǚJ]�:�Db���0��x��ft���6�nے��K5[�6˃(��X���9@������	���$a��Ε��P��� �(�#�f�0�ʾ�<1e��J$���$�/�p�o&`�5�y��ۯi�GAKa�VȤ����9��f1a�s)/3��;�N�Wފjg�پ۷�d�v�^�=���9�r0hǧP�#�x�cTf���iL(��D2K�,�	�FU�H��$Ċ&S��=Ϸ�cׯd��د^�ǯ^��ŖR@`C ��T�$L^t�� �1��~�r@���J�t_����CZt��a�h��|�e�3�)��Ag���8Eb~�����p��
B�y�Ė���f�:�5{RX��j����*���u��x<d�wO������mwaP��E����F@����C�"ƺX�U{3���͉����rgw\pZ�x���
�H��<���(&�#µ�8���G��&��'����,`V�;�:�}U���/g��w/#�j���\f
����,��������,'�$�O�����֍��^�����4�Qoc�7�9)X�^�M/G��(C�I[RH{1��n���ڸ�`��ʣr{O �[�m��c�@D�d��<j�� 5J;�)z[	\W�<1�Qg�8�]Fm��5\�o��C8��n��z��f�/Y�1���0�i��ꍶ�E����\~�zL?�����l�3�!�JD�����+�~����g��3�A���~~�z՛���\�	�tFZ�R���������i�α�#�m��oD;!�N�ny�o�P�����޴"��=��]�0��z&�Oq���Z����� c=�Nj��.A� ��*�P<�#�7-,CEY,��Y�z����� N�cZ����0��\�%<3��kq�z���b�=­�WI�G��e�ǚ�+����R��!�/SO�@'���w2Ba2d�T�
��Y�	�fL �@H�H
y���}���yH<���x��")[�6���Ӿ�Mx�y��^����P���(=C��&���	�$�'����X����y0�|�-#���E{KO(b�y�~{ʨ�x^�ĈN��귃�4�càYk�AG�:�9��� +C�?�O5��~Ժ��I�񞮨@u}I���_m����\N(�;�R@�T3���Kc�XS�)�v�bO�,��yAW�}�1��I��ͫ�	5� �A$׹�������!T�f�'?W���^hy����ܦ��,�`�y�$�2��)?* x%��0?d1�Pp��)���v��]P.����V�9��	�?�-a2RY���ű�s|�<<�8HFD�&O�⬂�2�X�$j�k���/�;k��l�Ñ�.�z�;.��J�h��$}��,�b_|D���s���'an4�C��k�e\v��[�e�ߝ�}��%d��Mw�a$�`�Y�?�;��bJ��p ��{�:�+��"N�w ר�ڼ}V�!��`������!C���K�Ft����Kr�K{7���B�&eã��>ce>�CZ˕eW�n��X/��}Z��h 賶�d1Tgs(�b�[3�׀A4�$-Eъ���������C��d�gt=W5��u�����G;�{�]vM��#t}P�Y�p�	fL�	fL�L�2���"�R`�����Ol� �i�}���,>�d8o����=�Ȣ o8�zR�~�r!�`Ψ�{b瞧O��\���)� "J�1me�K\>��tк#c�M-}�7���d���<��ӳ�g�2���n�x�;pv"4 �0�q$��i���^�y�|4��͌��R�oK���l�Mv����T	ᓬ4`=� 8�浾i��e����16;q�^�ǻ�u���Ĝ"�9ek܉���th);�C��3���<���ͨ峁��L��������} A��[#i���ے)I#<ko{oc�j"n_�-9��q�=F\V68&�
m�5���'"����f�9[Tn�胙C��p�wȘ�n� �0�@�Z@�V��_6�犎�t&�DcX�H��l�:�z�XO���Un͞���yD��\C�+4�|l-i��k 15���Y����$��O՜�v��vz�ֽۛ�5��ۄ;�sΪ����X�;��ATG[~%���%�&}��������;�PYQ��!�� Ţo��ƽ�� U�4��8���K!�a&x�w2񋿏Q�]�)z�����G
��km;#xK���=?r�&�ؽu�?�Qro�>]<8�a�2^�nRҾ�H)[�dW�箶��푛:_�3*�v��Wb�(��K����� ������ת����z�^�{,�W�d�� ��	 �{�{s�� �+Z
,~Q��%��$1�#���#{�]|w�#�'y4�����q�.c#2ǫٹ�@i2��	"��݆f�UD��� �m��I5�iڎP�bT#��Q�����XG��l_ﳶ>���m�����ڴR�6~�}�\�W��򮯜7��E��������H��<��3��b�����/{�\Ǯ�+����7�����	o/��{C��>��!��f�-Ә��V"|Z�t�¿GIٻ�{\���%�p�q�+�J��}�Ŷ���3�޳0_��s��w�M����G��ķ;�@�$9�/`t0�Z�y�!��Vlv�>�I*/ �a�9���_�����Ǝ��e�zba붸i�D\밆2i��v�c�Y�B%�ta�3�1`}^ȉ�W8a�]]�0����~�~���wP+�:;��07!Ԁ�⏠�,6��ΗWV; �U�%�[�-ŷ�3 g�Ĉ'��"�g�DY$�:?'�5�ol�O� g^N������]�qL`L��Nt�rD��v�>�~�_O?ltr�  �x���&��0��w�~Q(�z�'r�>�\��Q��	�7�������w�m�)(�[��d��i���6��՟�>cf�2tC��֓��cLp[Iu.����̼�[��XD�x������QS�Y��fɇA|��ClvU�i��m�e7������ǣ��;g��l!*{ݗ�ƻ��2�[��ީr��kv����x���fh��n��O+H]\�����C3���V�2�C�(�M��V�l�`v:�kj�4B�S���p�u7��m�[}�{*�%6ξ�-�N��):ꝿ@���WFk��o���r���Z#��Os��N�]�D��ⶆ�/ojH.���2��V��Nf�vxl���ن�!f��G+�AdNE7�*'��/�>�YO�p\�y����ܑ�����*@U���1�Yɽ�{�ܻ{���h�{���l��4����u��^5[��L̕g/h�3�or:8�늻Ms�Z+C�6Q ���noy(5e����1�2�R�P��;�O:�:�e�I�ܬ1����۪�\ԉU��ܑ�|z�u��rV���<��O��$�O[~d$t؊�U%�ɹ<�4n�*�U��7��	�]����4TV�Z&��@�e���l]��!Y��$P�]�D�r��Ӫ1����X�*�B��r�D��0���Ae�3�K�*����u1�͗�$��H$}�b�(;�ﱆG(�.��U���Lۘ����z���Qy�9���L9�����~��_ws2-��O�!o׸Gt���0�TmV��[���n����-�U���8i��e���TZ�gnq<볷�FS���L,��H5��㲂5}��h��4��+��\2=����Xf���v��H->�$'�֟t��7�[�����"�WN��}M>����� ���Fm�g����Y���!��q�����Q��n�oem�xW�>��ξ��}l��c�1�K�V�ǆ��f��}�Fxb����咑�5�iC��{��Z|:u��`�����+
D��З[{z1��[Şd�2�\u#�>��� ��TY�F�`�X�	����V���}0�Iz�i��,����X3�y�:	2.�YP7o������ťm<部�J���(>�S�ιr9�w�m��ck�Y�����;2[�)��
��������L�Ǽ�̔k��OA�M�k��/�����4��2�:m�TG^X§�3FS�����z�x�,T����y���*h@��]��lf��nr˧�R�/�Y��ҽ��z�E�TթZK��ٗ�7sv�n=]�T��I<�j��b��)�c-�\�C�R2�AVRB����₊�6BE�EGT�R9�D��D�II��Q�c.&���_��>��%�,�Y1��e����$6b�#�HI�P�#�faK��3v��qn�]��t(B-H b�h�u�H�K)c@�$��a��NH�d�-��MD�C#$.K�EJ��s�$zt��5��$����o��@��+g0̊ -e�ڰ��{d�ʲ��>��׬��g�>ٙ�3>>>>>?_#����ׯ^������%OӃ�v�ej�!V�*�[ݗiaH�6�fDTD@Oo�j�ʷ��ǯY����}�3�ffg����||||z������~}�,��=j�[_s�,�]��[lm����%jV �6�(�q��r�-{|��$�l�O=}��l�Ϧfg���϶||x����^�>ߒv=�Qm�b[
�T�=�c�:j�-F(���ŋ�Y/���G�׾}_Y^9��~3�>����33>ٕ�Nz������v5�
���eB�b1J�QyL5�ŊDb�h����mh���,0�&V#iZ�+e�Z�a�&Z��[X�E�R�EE^2bb�b1DU�.5`�b(���X�4TUEcYj�b��LEQV,^YӉ�*�Z�1{�b0N�)YTV"��Q�$�0z����-�mb�=�0Qb1NҍJ�m^��+PUX#<��j�����UҌ���癹�].<��wv�Ҏe�7
Tn�[�-6A�#ڊ���wqQ�BWsN��]�v��ƌ�5���k�p�`�,I`��D��cS�~B���"�8�0�DNF�e%A)��-��M�-�u��8Z\u�n��)������W�Ԓ{a��z�Cڑ��z�@1	��d�� �B+���c���s�<�@��Gߠ&qL���K�΁�_F Dy'9��b=Wm@��X���|�;ci�dz#v�^�+�h a0��[���!r�*5cz/|�Y _!u�HT���"�[w��^D�GMwD��, Y�K:��~~ "�5Ç]�O�����P(��k;�<-Sl���_U�}���r�Nc!�;��&�t������ei�A��a�w5ު���G���a�ʞ���xN����]}�Ym� �v���������y1���@�>��־�����X����=���ķ6�g �kUH@�gQc���8�hm{l��c�K�S�a<��u�����Ov��K)h��s�G҅G�Ưc@\��}�g\��ȗC9T�6���T-�����{<"��È�z-t��Đ��+�_�ËZ
�'6�~�~��'`�|G��u��+�}��GPIڻ�����$- �)�p���J���Ì����Q�]��0����	ZCڝ[�[ڝ����{c�i�a���!2�w�" �� ��Z�x��H1��4r
��$S�1u2˾+���g��/�����ۋ79�	�Ő����ޙy��W�4��U�,�s7��{�ʁ�L�R���S>>�h1�����K�Z�s�z+p&��r�L{У�2K��`�/F�4�����F�_u��2�&�=����sؑ��z�G�U�؉<z�N�Y�1,�F������i],��6tl��^	��^�z�$<ILm�y�J<MՆ��!��,M�T�>�Nm]�vnxp����}z�; ,Rڀ�Я�]�7��I>�lET?���^d��𸅅�c�{_=E�!Ln^.�˂���܇H̀8��97����ۮy�`��A��8r	h@����r�_J��>�*ṙ�Qܝ��yD".���ކ�8��d{,-�m���lYʈ_���D��ۑ8���2>N���`��c��	���y��zDWE�?Ư�i���������>�pe�N8{<�o��$���J,C��.*��/ <��X�t	5wJ�n��!Uo;�V��*(���<hi�����c�������xj �&N�8���@Y������ayN�����ݞ����N(�8Z[L�吅�z���J^%\$�=<��P/�g�z��ZLM)�qY�U��<I.����
�; Q'�ɠFr-6�gF ��b�+<��a9��>�;��6�	S�&��Y$���SF9��H�Z��M;�����7`3�X�t�������H��Kߋ���_N���elݮ̀��r�مM�w:��n���n`�:��!�U/�2��$�I�\�*
p;�Qr���\�s�D�����0�Ӟ��Uc���2�&��]r<% ���Qƪ���{�� ���,g& �&K� ��x�^��=W�PObT�Z��[U��28�J�������y"w :�́�öآ�}�H/��˿DJI�8��1��ަ�.�����:�z�@�q��gO��$զ�S�^+m�E�j�Gy��-��63_F���� �XKBƜ!ƥY�(j��%�j@�U�@��lҫ`D�_x���g�4���s��>��y�7�/��D��}O����y��=^wE�ܐ:0��TC�Z}��~�V2�dx�ӠE2�+��aߞkة���a?��Ja/7�:�.=0�����80�	�վ��:��E�p'��C��L7�3K���h��������L1�&j�$��ӏrL�W���M��I�7n��o��ou���^����Dmu�g���8�Fl1��O�c��cn;��0�]��.NԻS
�ۆn���g��)�n^�p��p�X���Kv�
X�2�N�Jń-���}�bh_@�W�5Q�;��!��ޮ�p�����b�׳l@�Չ8{qE��2y� ��_�q=<�\:�f���v� �X�@�.�j�Y���m�cV� &��U; oW�r8���Ҽ��7!lpc4"꨾�w{�^o"����p�-���d�!��)W:!��x2O����� �:��)�J���q�&Z�x�Zȡ��W0���Ceeah��v��&g\ͣ�(���?��
� ���x�ǲ�װ�lO^+עI��z�{bI-�	��~�������� g,�;�<s1�M�zL�� @h6h��d�� E���%��� �؏wN�KA��c��7�pֽ���1��S��c!�e��g��5&����ٯ�O��qb�	��]��ɼ�tHì �ep�t�Il���<r[�X���;���޷�@�.��g���q�0�87=cܴ�5����{oc�O��C�7s���J�~��ǁ�o���~�h�L�5ܸ�4��N^��~.7�'��/&�1��8ؒ��lSj@J�$�Z��N_����^fa��2�f�M�Ϻ ��>���#@kX� 42y�4��?���N��|BF|W��aS�c/�YxG�4E�rP���3W�Y�a]�1vՅ8��K�ñ[����ON�uS�t�1����f��ۼV!E%����C�����y��hix�ހ4�l�;Y˘�ō��Y\<oz�n�5�������>�w����#0� 3��w���ڛ_z6W5en�f�E-���fhiI�����rł�]��cl�1� !� !�cI4�8+ 凳#+���z��ɩ��lU���W���X^�P;Z�L�d]��� j���l�e�t4?�t"�O躮��`�@Eb���!�d�@FH�'$�X�e�3���kcux�*5�������w6Qb��]�n�[�F��!9(�]�>E���D���rU��L�$�b���^A��AY��13�&���XHV�7-9�� N�2aHD$�ez�$�Ǫ��ڒz�^����0 2��P�����OiL�8x�C�G��Q,���ӎ��vG���ރԁXD�ن'� Z|��o=1�ф	����%Ѵ�=�k�j"�p����sj�vφ��{,2�/_�ԑ,�����d(�-�j�/S�l���\��L�Ž�|�Ǣ�[�e�(�f��c��,� ��4I� >3���o;Gbڵ�*��^���q܀��#!�sbuNK��Z�����m<���I��hU�Rr����Ez�v���C!��[%ڷ˛��l0���a�>�D�4��C�F7�� q`�D�x����*ܩ��.�34V���KrVčVx�k�@ĢTrU��k��
���<�n�ls���/��ڽ��5�gY��h�dзb����`S8]K[R,F����n�	|�Q�Q��	��7�SK��Ic\'���w���@�y	ɬc�,w�����H���������`(O�p�z��TKȂ����s*��W����7�����!����7�@(����Ʋ<@�kr���,.=�x���S�v2�@l2Ҕ+؍�D �h[�q@􅄽� [Z�w�җ���g���/�]���LjSS3pʕGٕ�!u+�'}+�����}��uY�1-ά�P�3X2��5�ǃ߉$*� M�N�(T�_n���MdSu���ţ���ݛ�>A�r�^�H`�~�2b�� �׊��'�,�$��{I��z�$��$��E��Z$�o6�> ۩��o�@y�zP�e5��讉b�a�~(�/����W̗���;9C|4t\eTuvf����-�pӯ����(A������j�Vyߗ��T
,j�r�<�=�>]���;�O��Ks_T;�8��"�a_-K�if?|���-`���A$�	b/��Ɲ�/�_үj�����=����b�nّ���n���@�5�x����u��C���%����d
��������wk�m7���po��q8��!ك~��Z��E1���Łdx��{����}~y�4�@h!��:���u���Pz��H�n��Z�^����%d�0�ҿUX�c�A�o��9��c��F��2���ݛ}�_���S��L��<�3��F� m����U���A�9��#i�xX=���7�<{��H����&�#HM��G�`<Aa�9=G� (�[�kCx������Y�y�2u� a��������C댇M�:� �O@���-��W?R���k&ZNz�g� �T�\��y�~�A��h�-�űic���XаU~2�� E��~��>c�+h�M�=܁���/��c�]�]r`��dkQ�5���;�m���WU
�{����()�oj���ۢ���F���1�ʺ��VP},���ۦ�������QDy�-�����߼Y�"x�^�	<z�^Ȓx�^��Ld "��`O�����>���	5�#��f���;���c�H7-u��1iH���t�;|��]�ҁ������L~ր4�o�]2Z�Q�S�
ށ�~=�3Q�K�{x���	�Z��J�����izW4#h"L����$�@���{������H�2�d^&�z�6�zT_Wef.���0�;�n!��wI�ͣk��xZRy&�����	���cFl[��Y8�S>�ٿw��A���bM%4�b���k�OM�� ��y�z���筷�P��p���"�;�dS�8gE戍,ЎgLN{7J���v�����̟95��
����M�E~�ck"�$�u�u�$���G�L�s���&u��C9L�����d`4�J��<s�R~�$�1���:[��5���ҟ(xݞ��{�o;��Yvi@�$��o_�6���<��F���=h�&T���DR����M�sҀ�Cͫ�lZp�����i�X@s��G
}�����=|��yP��o�Y�7�V����c�W���O��r�g9q��d��3��;o`�co�+8���s^����h��4��n��hK8��;�z������\���;�.
}�Eəgoc���L��$�^DFz��.LΣ89��]�ijuPO�,������.sQ�Λ��Ϻ���l�p��f�ns���@��3��&$�r1��IǪ���ר�=�e�`ĳ3 �v��� �T6 'ɥ���x7�᪦|��V$]�D_Ʉ�=x��ڀ�+1o>�ދ�}�u9�8�n���Hiع��q7��s�� ^Zܐ8�u���al��{��<6:kA#eS�[�y�an�hyuFT_�p�*��	ø+f��`��;
J۹��a���X@2E�rp��Թa��x��{yO_��en>��p�.$��~-�}(5�V������peVw4�V!�^��f]}{���_w�����p�`��v����x���O�[9�= E $��lN�����3��.�N�m��S�_�"�T��_*������ ����q���/���?���Q����g�:фm\�и�Ǜ"���r'�{���,�y��4s�!�+�e8ù[����4Z�mAb[��ɼL��'����>04!���H���VK����W��FU�^�Dm�Xֻ"���V���^XIE^�d����~���Ζ��7��u�ԓژ���}�{^����w�T9��]���m�&����D@���cHCX������'�������]�]��Wщ˙rv��F��ܨ�r�z��3�f}�gO��?��unr�;��>|d.�Zmg�yk��V��Lf�Jj��ӎ<E�5u	f�ʺ��v_�";�Vm��8�n^<]�w��^;��T�/����K՘wʧ='dD&�6�j!��Î�~F_�R	%<�a\�5Z.c��q�g� K��BY���I'�U�ԇ�U�؇�Ii�� f`G�����Dt��u�d��$�B��Q]匳�}Qe�n�M�+�I��lV�a�.��S�
�/����9C\=Nem�q�8�C3�BRJ^:���#�j�G�|@:x&�|�u��N͟� "z����6�vEs+�/=�@�p�z9Ɵ~��L�s�@�oC	c���75{�b.�2:�a��Z���Y����X� I���G,�I`�<�`���3��^m[�����
���W����5��-�����ba{i�z�jB����sP�$�h}��dS�½��񱞡7}���x�!���c�U�L@��o��n���"�0��Y��J���Yւ�����²f�n/_C�;s+�vp�[��$�	��Ÿ�[ɳ"@��Q��2��ܨΪ2;_�73==%8Z��\뷱x�;�m�����ԙ]c�A:ĸ��r�}^�HRw��ެ��e�fkiN��pK{L<������l�On7�Ns���ZY�+ o/
�oF=y���f1մm{�f��6�����q�X����an0�X���qR�\�*��wWӫ$K���]����T$eL���.�uV�ͽ}���T�4u�B3q!O�M\y;�8���_�f�z�Q�C;9Nw��vS����N��C�n��I�.V��ڒ��D�ܙ(ǝ����پ>���$��#90�2W�R$��zx�^���$-�3 w+f�����0��F�o�p4+\�:�@�0 I5�(8]+<%�n�$�y�g�w��"/1U�s�����-���pِMp�hGSR�=�ں���%���qsS4q]�Γ���<�`�3����~c��߱���
$F;<:ϗ��{�I��>�����3R�8B:}�����p�H��C�3����,@������W9��:�1�Ի��Z�����O�jZ��"
*�]��T�����hK���,��sԚ��w��5|g��.-Gj�kBnhS��#]�x���Z�pT@��Y��)J���ߝ�L����l6�M�;{�CElú���r-IT":�x:����P�v�}es���Zn2�vY��#Dk�<��f�y0��W��b��GX0��E4Zb�	0�g�I�� OuE��S���N��ۿ���� ���m9����G(����uEB�E�$��@����.���
�ºNw�p5���Èww4�ǯ��Nڣ�ZR�M:#{�+����i�X =����ѹ���a���>X�(9qLt�&�����3;Dts��u�b2L�n%Ntu��u\�;a��V��'�r�s3��L��<�ҷ�]��ne��\�NOGrpj�`*ͦ�T��l�uN��<E��$���vrK��Ȇ��oB.�0�(���9�*Mf�=�7Sb���
�t��o^�&0dn��5�5�	Yyח�wX"�ӽw��2b�MY�f���/����͹;no+�]�"��)���w"�v�h����\���#���8�$@�96�B�Ly�}�N#��#��8l�6^ڼ�Z�;YNwg4�θ�I�[�˦V���x%�`��%��)��N�w2Zyr�9ż�ou���d��8�(^�3��f1�'`Uy-��ћ<�\����u�M�0��
Nlv#��N���-��B:�`��U�7v�f3|7-��P2�!�AoE�v�Ѫ��hh��;#���q���X�IveB�#d]p*����İ�U���I�xFAuX[��k�
���7:pPI8�|���.yW��n^lc���2�4oZ"��z��PaNmS�����*�T=�t
��Zt��%�f�ZYi�)g%۲$ �V��%��r��4a� Q,�p�F�=�"���N�Gĸ�'%# j���"���y��6��Ӌ`��;���5�j�~�����D0�*�JrX����|Q��u��(��S9e=}�`��J���9�R����|�����뷼Mй�t6LWCrm+7Q���z�D�˹�12'FɈ?3U:.�ʪ
����ngm)�S�qÊeUN���9b���(�*��m�Ԉ�P�}���v_r�[���W����
�U��m�
ћ+�]\�`X���w����v���7ܧ�;5"�v�������E}wBj�|[��0me���,٨ˣ&��讒mΗ]4*:J����Y˵�r����|G �5�*)Ip<"Y����mĆ�y[�H�:��w9No�����]��w+��z뤙S��pΊ���ܑͦ�_W^�܎�l�F�Rmq�dw�����f�	\�7�uL�rR+����K�.���c0p��<.h9�;��V��Γ�\ɴ+���R�,CP3�a
2�t�<�\	��
��Z%e��1���Qs�
�G�v� �巹�,��Bd};Yg��}#�{3wf�+�����AJCIYE�9�k�<����[U��y!���m��`��H
��+R�
����ȫ}�>�}_j��x�|s����Ϧfg���϶efg�Ӝ������{X�XIi�J��b��H�_�N�yJw,�������|}33=fff}�+3>>��>>�oŶ���y~���/�y��QԚ��������Ym���z�~>�o��ffz����fVf|}9�|}>�$�g�ߗȢ,|�QZ6,F{Jvʊ��D|�1�F/��������W���}?���ffg333陥��fϧ&͟N�NҌF9q1�j�i̗�k�Nd-�eY�)�Y����E��x�q�)�e�U"��ngPp�E"�
Ո������Q_�EcQ\��h��5Q���5�-�TQ�T�

�r�EcF,�1�)`� ���)��{�u��"�hZVUkX�����Ȣ�D5|��LaW�VL�,F<��(���1T��WX�1M�R�QL�Z�F�YX1UAb1,�3yqQ"� Ei�[g&�-�iou#��#G� ��[-ޛ�1S!T�u�ST����(�Z� �E�s?�20 �,gs ̌ɒ Y��{l���{ ��!:w������,%�>z>c����;(��!�~��	7�!q��#�7tu!.�ye�vkw���}���0F�D�XOB1�qj�%�r�@��:�n�c���DyI�����9���:����|�O�z?}�mͤi��o&P��R����@e��?_�&~`o �뷻7���/;�D���V[&�X�ò���Ŭ�i�bX���s_J�g9<(7��8:�*�X�h2��K����ED�mx_�G��c�u�m0�;� ^c�a��$�e�xjQ0��)�H���P����3��Bn���=�!�>g3��<��@�^҄�a�5�"βMF����LC�h�� ��>����x�K9�@<#��*H<�h$=̫����)��gzH'�B1�jmG8���U�K��?�9�Ǫr��S�O*��	HA������ixh�qEn���'������'ڣ���������&�w͹��X�u���Jw_�G��Ui`e���o�\��{o�N_H=
�hNH���, Z&��6�%��&뢱��#��z��.D��z۽|�R�ȍ}�z�zc�0����§9s�Ic�}�7�����m�|&wD����$ǭL#���r� � �#��
��b�yj�[:J)b�F�np�����rJܕ�=�WS��ɯ�ǒ��u����*S!�s��N�����`O�~�x�	^�x���*I�3�g`vvL�3k{��~�opoΰ�,��6XC�j�݁ kȑ�p��b�YixC^]���}����;�;�5�U�n�d/�Zi���)� �c�~�@0~#��?%��H	k���·:9�<�ق(����P?|A?b�1(gZp��?���^�y��lQ�z(�����ᠰ�{�Uw�UӒ��=��4���qv�sъW�Kr�wባ���J�''k=ۙ�֙OoE��4pa�K�o@c�
�Í!x?Z ��x��r�v��@1��u�]��y@Q������ �9��5K��sm�I�t0��u�r���O�����W�2n�c���i`�v�r���xl0�P7�ȍ@ZN��`�)b���0�L�����\�ׯ����&7^X� U>���ᝢIs���0�>qR1�K%D;e0��t^2��˺�B�y`n��}i��	TGF��=���N�Dޛa�h������Å9��mnӻw$��{m-�>Pw�� =���K9T-��⚟��W����j�U�Ц��紬R_����\�����,K�n��{�EFq���t�R�JY���/v[܉3Ɯ%���	wq�^!UYh&�X�%��̋�+�%�%4�(�z�����{x>"N%�'��u�nBݮ{�+iĻ�q:od����i��
���$X��Sԋ"6c��È%�Kw��o�I?��ܳ!�^�{+ׯ�+ׯ�=�R@'�x2�*�'�����N0��e$��ks�S�Ϩ}��W�ڡ�?`{e %z��ί;����q'�j�:w#F�����>��҄�����Ak �-ɧc���5�{��<�3��"��y槏�v��{,,D�F"�8Jq�>hd��"%�;P���H�b�' Tk�N��oD{a��~������f�PcH���ۓ�b$Qqz�73����;�U��5u�w��Q����~��MS,*�!��k�%�^*��Q>;�>�ɂ�I�	&݀����<��Z>Ѿ�O82�u�x��B���	���!нN/C�S�_�`>5
��ϼ��y�#lu��8��wy��MC�`��X|/�Y���MMP/��?g�q� �v�ǈ��"�rf��<-�z�љfa��*��p�9�:2����c����z�[��oKHV�ݏ��X�^!���mv�w�*��93�.'�Ȋ�AP�" _�殺�\sn��[�����@N��eZ��h1�~~����{M�w^�7W#ܻ/�����.��������T�0v���,cP�0�dr�����F�z�H�pH������K�ֵ��Z�K��ޡV6��<��"�͙0�T#�pN�:^w��m1����v���4���^���ggN���sfAoL#��C�l��s�������1I�nod�M$I�C���[�W3�@?O���L��Y��P�^�{$J��ǰ���?��m��y����6���Ï���M݆=�q6�ƵY�`����
�I���4�0f���0A􋹻��ׇ(��C��y��nqU���٭����P��:�oK�"L��m{g�*n.�/Kw�`��J���3�c��I��Y��UdxOF<��,��� �#.o�� �^ھy���X� ��^����`�.��)x2�)����%<��S�09�|�Y���|�i�b������"1šn
��,J�;
uԷ�]��{փ���1��� �Iǘ/_e�h��pX�g�G	/�����ϥ�խz���tV�v	/�>]�����	�0t��!�M�����vp��@X�8��=9yw���	�P����r)�������MoN_����֙1��b��@�J���It&��n�yDC�WOO��=qW���c
�	��fCĒ�/�lU�Y�^�Ϙ��q\� 4y���i���Te��O]�o��
��u�D�#,gc��m��+�xB|���C�8q+~�y�z����C8_����ٗ?Zx(]0���h�i�!����]���s3/��`'n�(|f�8�>�7��NsHޫ��'Wn�y�F\���ѝ��&D�wU����cR�K��{}�w���$��N��$�ɒ�!^�x���Ǐ^=�B{��o��o��������=��t;�����-��ꏕ��p��Н�A��QRy �Cc��h��e\�W�q��]�e��]�|�����Z���k���=����,Cמړ�_��s��A�om��;���0���&�ʯ�=�����E�����+���b��ɫ���/��q|~�Q.�b}d��q���wy�H���Ô-f�c���[�Um�E5��F�g�7��2a��$	�����2a�	���>�+��4�H��{m��j�Ɲ7�,�Y-W�N��T�c��Z��O׈s�^��K�����q�Pc��~�<{�����i����N�:N_tq`�y�̬���!�
v*�@�rz�yey�`aD5t&/àK�W����f�WS��rP���@{y�1
���l��)�c�G�,dS7�aX��OK{kcv�g9v#C�Qh���9 ^��	���^@�\a����w�Iwr��K2��P}+{rB��>ٮ��#vvl=�q�������]��+V?->���z7��>?O�jE����)>�v�)仮�����sv����=���>v���̽y�`�F̗w��"=�>���VT��ce�N=ޫg�Y�m�FVmX6�`�Y��o:\�P�c�9��JZ���� {�����1�e�,�$�̖d�2Y�I�Ā��̋@r�(�i��$ca���MH�r����؋Cl��}L3�M�ܝܯ9J{���.�T6_/�ƀNjo<B�gv�ǐP������TM!Q3�(�N�������3���y5c4L��H���c��?���on���=�D��5���dn�^��!���|^�8�E>�b+���g��瀲;W �b�z���>r!�KF��@�Dvƿg�%j�Q�~;3�D���^�f��et�+���B���t��Y�����J�w��/�:�;>E�K�~d(nr�a{�A_u��:�#���@�=�@�.��L��[�ű��=^w@YL��~�^j�ev��n��J��f��gm�5��֝�B��np4ޯ4� SD���^��@�1�N;�+dׯ1Cj�K1���v\L8�s,,LR=�V�6�G�r�w¶�f���6k9?x�_E�7�v�:�Q���Ӑ�0$oE1�2Pv��Ws�&z"s�K�G{�/1�Ҹr��ؼ10�͌�Գ�\f;X,�ZC�d$�I��u���~����#V�H��^rH��k��7�fr�I��C�Y�\�v��0����O1��m��^�c��hg�Ux�Qi22����dَ��;;o��GTU�ա2z��z:h�=�����nn�ܺ"߯oA�lK��֫N��L4�6\�UT��H
�����j��q���6��o�HN��̑+ׯȕ�׏Ez��О��"�M;��O�ovO��rI	9D� H�Ia'u5� ��r��a$뀻z5�շτ@� ��RFy�<�ƺ:��K2��a�_����� ��F�J�* Vs�n���t��:!�@�L	�$0G�;��W��y�y�ǳ��i�B@q����~7t�s�a�2���P06T�?���V�<����� ��hg4�>`i�~�'�� 2yO�*ݮ��p=i��S��X���[���M]�[Ά�Vx�2t�\��2��� �9������a�p�&!����v���ǣ��;6�y7������8ec�-D�����<�}���in5(��+|��xg��ν��ni^�9E <!A�	�M���+]���Ǚ[`-��2k��jޯ�L��&hE�{���C7� �m�r_,~9�W��&�G��1��>�a&��q�������"'�)	�R~1���U�%\@�$B(�D"M�U��4�\�
�~�P[ܸ��ן��M�H�wʚ���OBrm������Z������b)xo�4�~#�82t)�b\l:o;=��ZF�˗�����7��m�
�R�!���z5]ٔ�󯪪�z�p���"|g����]d�Զt�y��B�^�lU��d�ދ�1�n�)�>�n)X�&��w�x��E�� :���kA�m��?���Ǳ��ǯ��=x�E;;&v� 3�n�v{���35�Ӑ>l\�b���#��8�An,8��E9��Av�:|�ʳ3����8݀R��l��NH�@Q���s4�,�q�@��&_�W3�bO��n�u�<?�G�MO��Ճ�{7֧��q^�a���@@��g�G������_���꣣��/3�W�"�<Oc�5��l�-�q@�����a`LmyȌC֘�"�I"p����x+چ�=�y�K�h���heQ(�;�<"�T�\7r�4A�O~��J_���w��}�E`�E{�U# �J�w��߻����!�����4��6�L5�@> ���xݫ;�ᦱc��;��.1�𭼮�C"R ��NX�q �|HS���I�$\�F�:ym)�����	�8E�����9��qkj&3���<���D�u�sm�'b�I��B���[�J�P��#�'�_�-�]w��<͸��x��큐��ͫZ�D[&��Zh�� \б�>�Nj���[뛜]Y����ww��~+p Q$.1��k��sy��# >�p	��d��dә=w	ǻ�)��{�|���g#��J���rs!XV�'�gfr�ҭ7FY�~Y��Vd�	�f�}ׇ���.}lV
k������5- m��|:�q��	�Ǹ6�n#�4i˖dݫ�4��afyC�n��y�����sǱ+ׯ½z��3&K2�HM޷��_�u�7���ߩɢCU@g�� ު,0��#щɄ�- 3����N �ּܱ.}���D/Ï�}=�~�D;�Y^yts���Y`М������5����]'����%�����+Tk���8q�X�Ag�P��E�г6����y�
@G�9�X���#��]���(-��|��(��?�ПF���7�`�č�s� 9�P`���3�cz�~P*����o:�߻N$J�)��l�҉�44p�Ê�V{K
bw��3ESR���}t��卸��t�^�b3;��3µ�Sw<4��X��ˣ���B&$qNR-R�c��=p^K<�� ��^��R�țަM�(o����Ę�p�}j��v����wf@��j4!I��������z�\�c��sn���s-�H���c�@b��s��{�����s,	۳�� �f=G�a9������}�>�z#��r@��ZA2��r�̸��,#��]�E��\��=r�����9�O~�ܜ��9�^�8>:)�Z�JC��ցń:�QRGg�����~�Ǽ>��	���t��i�E�@��Xʝۗv��vN�]M���Qۓw���Ǵ�w��{{�9��{�dY�Rq��Y*P� 0U��|S�S�x���;%����΍�=x��rr8q��]���/fJ���c�e�� ?�w����ɒ�1���d�YfK20�H`3L�^�w�&�	 	+M6��aw���a��~�}5�eQ�6B +p6[�*]�u�QW�
�v���ㇷv/S<��ڮМA�$�Q�M�ac������]��޻�p�sT�y[:��I�<�M��s0h�] \��LD��5�P�k�s�S��8ƍf>�Q1[,�g���R~���0Z�,xD��8�1�zb����)�HS�2Mx�v�\��ࢰ��`�[=��\	�;H�:����Z|�T�-(�O[L$$�:!ǲ��Z�}���\�w�r�Ǐi��}����{�)t�����󓪴�O1�����z/iY��I��374R����y�8�<���SS��+�`-P+�C\E�������w�".����!X9#{h�������u�QJ������C}�^r0�z�%�������.���=ש�ק����K��U�U���4� @���Q�Ϗx  �/��\bXp$!���>�Qj���U��)�;�����y\���H5Av�s�k��}�#ٵ�t���0`�ۤ�����tH�%�2'���qIQ+�e���ݶ�Ǿi`��qEh EwU�(�n<�R^u�N��h��I�7�����Ýf����齮���,��m��VZ̡c�H�jm^����	�M�7J���%rPKv���0��
/h��v��eeen���T
F�Kڝז��\ze�VĽ#]�a�7#IN�;&��zMၬ�����j���;+q�M�{̬�X�J	]v:�b�_@D��[<��[׽�O�x��t�(*���Y�W���Ԗ�!�|@���൘�B�Y-h23Dm�'���ˇL�熺%+X^<�>L�S�c�<�"ɼw��%<�=a�e^�jtWy�՗I���3N�&w6q�O�sx2n�_S�/na�R�˃s.����")]f6J��/�/���$�J�:�v��Ίd6��<��쪠�ﯯF���v���b��ol�-E�����(�t88�gtN��p{�\Q��׽��4߹�_��Q+��[��|(v�n�
챨��{3�V��M3�wI��D:�y�8*gXvŻ�]��~쿉�'�b	[����+xU	�	��ݛ����ժ�btǹU3�Kq��Cu�℈հ�f1B4
�S8P�{���n1*Q20Z���}F6i"����U�j iX��Q�N�ZN������̷T፶R���Ӑx��a�ا��)^����$4�k/E��J�T�Nz��7*0���%��y�_=�R��+j������,`��[�>v�QV\���TX(�Wf�����`ޱLG	�e���>(멌�CUV��2��Q.²��4��$�ue��;&X��pcy�_uΣ��#N�u2��@����B9{e�5l�k��S%Oi7j�ݼdv�ԆZ�s�C��������n�FT��W� �+"Ji��+%��]�rp�9�K�T��b̳)J��=:ە�"MXǅ����<O���[��v6A��ֱ·b՗�P�=���<:\ ���ros/I��us'�X�L:r���Zc7#��^�
˻!�Q�'�q�( �W6�v-��.Wʥ�L��{���G954�rԫ_^�|#�iL�5qfE5�t�s��m`#3���b�{d�h�"�r�	�Ù��\����U������m�\��G#�&��Zm�t�%�}R��Ԉ���G y�lѼ>vʺ=�����ַ�&)�Ǌ!��sx��"�z,�t�u����$�u:91��v���Rn�4(8�5o�:\*���v�:�'��u�����\YqT�
��|��u�Wc^˽�ݮ(�f&`̎��-Dqh���¢��Y�G]l���*Sr���;�p;���v�W�Bf#�źn�_-�=\�8y���w:^���3��g3A
�����E��U��i��q�TƩ���7xY{ڤY*D�j�bE��y�`���W�A�����Z>�H�6i�#e�I�a�J ~I$�-�-č�����fj+�h�hѫ�.&�9��Z�)��5n���^f�2+��7(J-���f
L�E�q�fnW9�L��4��s��8��h鐑 Q"�M�@�l@�F$L�	$��qg�<!Q<ٱ�#�ܺr`ㅯ6[�<7��J��*Y�I�Y��\�8��1ao���e���׳�꿖x�s�����g�333���������s��vȼk"$U��N�y`c�ٙiDE���V.ڱWٲ̜�g�������ff}33ǳٳ�ɳg����iE�PR�
��\JbV�d��m��U�S�Ul��Ξy:���>ٟO���㙙�����fg��s���~{{G3�0S�aZ�*T�5(��b�-�~!���d���}<�lϏY������ffz�s�ɳ��~���}��1�)�j��-&9K����6�y�Lu-h1;N���V
(q����B�nm*�AB�R)���".ڈ��ݕX"��>��t���-&L��`�V�a\n\pTR*��X��2�YYX�R���։]�V`�� 	���e8�QdQT��e'."��9aQS)̨β��ID�R�h'�A���j�xy�̚����m�7[bev������/����w �c�����b�3M�qҬ�s��\�Y ;Ofԡ/Z�QH�G-Mj��eD�l!UL�����=�Z�i����w,��%�A�2Y�3&K3��N��m��}�ޚ)�I�s���^�䨊	v��C㞻��Vysy\z=�.�~���R�ZAfH,h�x��w���8o=:i|t��|<]{Ͼt2�b�|Ő�3��ޗ� ��>���=p|�
}�^뽅? ���g������{��ô��@��ft4,+�i�&"�H6l3 ����苞�4��=�!�'pR��ޡO[��K�G���fпX�� [�X�'	��>��w�|�$m�b8]��/c�(�ǻݤxf/G=��'%�'�0O��S�f#��l�r�p(�.9s� Ƕ�r�%�Z�M��|�g��]nǛQ��ȑ
\ξ��р�)q�TQ�_�.�8f~��%��.�-��P�ISuՃs�O��w�X����H�)�*2��
������g�S��{�5)��6���y�?�#��K!4��M����� �$�sD�D���C��;�	*�j�+��O�@uz��W���rƦ#�}sz���{;bk���s];�@t�g�:�={;��6�g�E�X������K翫��:�ay��A��;���dk x�]i�]tU�W%&u�ݨ먹��J:��Ex�Ykx�:VX�O�ԑ�|�|9����B�qHóiLOَp�:����qhu\�[�)\�+=2s$�(�t���0�4�gŝ����׏cՒx��ǩ������~|�O1���>z�.X���
m�Z�F��*$�^b�hΞ���GL�+�N��ty��M��Z��Hпty�ҝV|F������>�b%��r�ݗ�;ՕY��j����1kHoL7�A�e���j�������w�K̙ﯳ-�i���n ,`U���Y���p�	^�:�[�
��D(��=�P�b�(w׏�؇��s��\3ک���.����0���#׎�	��_[��m�#���	tB�$��y���}�1C�ΟL��]y�}��7+��M�V�{�Q��GҀG���,L��a�\�G�GtNd����fg�ۅa$�Z#����=��)^��%����-���Q$��M�;R|��}i,��ҽ��Y�3�;��l�~%��6�,��x6Frъ9KQ�q `叝�����E��M��)�#im\l�OF`!�."���<���=�2��ܬѪ�ΐ{���C�^٘�|�G�#�<z/���	�`�*~��1�O�/�y?Om��d��kq�9ʬ�HU���UT��޿r�k�����������-W���ۏ��e|47�-��L�03����'XGu�h��˓x�O3�����Gr�C**���+��(K��E*�z�0�
�-J�f*�h�������̙,�Fd�f@fL�`bKi���~o���\�}��c�A�R���"�1��u)��j��M�>!��)һ���v�:bz�Ҿ�C�({9)rk$���.P�w���/�4��s���1��5a���_�` ��5���Yq�:Yjg ���,�n��ZdR,X��b��5��"!��6w,fx�y�w5l
 ®��]����ِ��',Є���|��
;�1.��6m�Y�E��L�"���U�(¸�{��3�#p|����t�+���ό��V3T����0����N$����CF��������I-v�>�6�Ё�Sr��q9Dњ�qd��^ͮ���9��Y͎�ӄ3����_��_����zI;��V�<�(�7$�XZh�p��k�/c��k�U;t��3���֔{y���^�u�ɪ���˧�qP�yx���[[2;f��b皁օf�
�ޮ����l�6Ͽ2��/D�Ɋ��WhAv��R�׹������+��D�bN��0/9�P�Tu���JO<TIn�z7�,w�ם��m�̨�=��)%��w�B��*�(���r����Ov��Mʶ�[�._q&�_� ����j�XgF�v�k��Q��N��^�oK͘�V�D��ܺ���Ax􍰍�p?�O�����W�^=��z��W�^=���aћy]���9}�����z2atۧEG�H�x�R9��<=�t��T�$gT\/H��z�H��Q�Ȏ~wI����D��|e��Rgl��Pv�bn
��=W���<ѱ}��X�,/]"BL��Z)�[z��u7�����u%�K�Z]�n.;�����Y�s���<��V��w��;��'e�\�兕Z��49��F��1�o˽�����սTvn�==��w�4�8֖ย5��|�$A���zv�'��n��u��\�}�7��s?�s�G���B��{�<(�|�n�g/.��ä��<ph(�ie�1�gn�h��7A觴���z�-���u�2�䎇�v��A����4,����B�;��ip�̭ǽ��4��:k�z<�^�	R��Bf�z��w�X�l��w{>W���P�z��	M#�q=�TS�N�Kw��#-/g�ق|�l R�2K�ߗȚ�y['�5�����5��F�(*V��چ�>1�${��C�
�[��#h8i��wK�<�~.�Y�_����͑]��m��%prB����'|;���u;[Rn���C�!��`�[B�#̢�7�!Ő��.�$�
?Q��BT�U��B�ML����>�v涇'�qEBs=���y'l�����*V��.�U#ք�bͰ��"1���6!�2y���q&����-)W2�Www5�*f7��~�?K3e�,��%��2Y��yG���r���L�
I����N��Fc��m9�p�K.�����T/�8/�?*�q��յ�X��9�3j�)Wb��ͽŘ>_޿*i���g2GP���EO�}8t^�:^Z�sKI7;o�?v�u]��~M�o<V;Mr.3�7I�j͗�wu���I+���񉄽+�=���p?xe�-�(�0�Q9c���`}�Ȱfu�&��;���cw���p���<��o�h���t��o��H�厏4���0E�M#����0�����^��vz��9��I�ܲ=DsǧCҖے�l^�$8��1Q�p���ĭF������{��^�����6Kz�aO����jrm��#+ş�+��t1��UI4��zc �>��ِ��/����C�u�W�zx��:��{c;Y�C���"��u�=�~5e}[��ߟ���)w�	 ����ڴ�.�&=�e�Otm��\<�.;޸�9���>�ĕ!8*�V��?��m� �d� ?n��3��jvև~1~h�~����{#w*���� ��lb�z���E���[��P�TRol�G�xkT�l�8D�:��i��2���d�}����d�i�x2=� �$�@$JJ����[u��3j,S%�蝃5���0R(���"�3C�Fԥ �&��,��o��i�)�;�w���?���?��J��ǲ�z��z���	j{�}��?|��[��G�ɑ5��P�%�@��a*���j]��xL
c�o{{z��1�5���h�4A��QvH[�|m+Ь�ڼ){�<�4
^l�vi��.ǉ��ǔI�lh���O�kŇ�(� �G��FV[� 	g��]��t��j�[��|c�!ڕچ�c�:_�����Q<��[<�yA�g	���XD�������XI�'�ge���}�t�j���Q��|6&4��|�0D����Ȳ�_�������a|��q���2 �SE�ނ~\�^��7�0�u��"Q'-�{6���PLRp��#;�������8��5J��k��ҟ��Q0��þ�uי��9���{7�u{'�G�����=�m}�cV��|XɌQb�H��C�	l1��F�.�y�=}�z���ǶMu�y��WSz�39j���pߟ��U�~�����l{��۾���̒==����07}-��n��4�z.})�.�M�<�-b�wٛ>^���2u�׵{h�cu�\}X&��z�|H��8wD�����G�p��`��(>���mC�h�{3��%��Ee��L��y���q�ǽ}��KZz��:�RiV��tرT�:���.o������L�`̙,��%��Y��3�r���w�9���ڸ�j׆" ���b���	���g���N�ޗ�]f���&/:(�S
���_����Üܐo�ɟ8����,�hc����l	n^������/��r-����z#�мG�Y���+A�!�-i��nmȌn�y�m�z�Ye:��ݚj�p.q'u�Y����!����	q���$���Ʊ�n�K�<���������������u��+��,&S �,wrGY��hng�S*��ǚ��HN�d#5å�I�Z�i�c8n�A��w�-�S�]���#N��Nށ| g;����_S+��_R������y���)�r��nC��}���݅�}N9���4v{�� y[�lY}׳��R!i��9��9�r�W������EG���d?p�9�&�����U����s�,�'-�͵qQ�Ղ�l�X� ܸ�^����gV�y����A�|��Ӓ�<�p=���{���5�c��3��u�8�� ?�3���б
�ż��)iU�@�4�n�to��v�^ã��6�*[�Xܔ���b��P���ݹ�l��e�^~+ޯ�6 g��9="L�ڜ6M��7f*�yގS�/�{DcNVl�S4�֭]U+'-��nU93���� ��P<Ӳ����tQ���͖b�ɒ̌ɒ̌ɒ��g��=��e�_o@{ n �&�c�i�zW&���^'埧��I�hZ�tK�+:�_��{�+�����Mn�vy~���cX� |q����[n��&��=�>J��_h�D�_�RI��<+�j۝T�d�~S��/cA����2�߷����F�D�_���߭�E6"����ѻ��z���H�����1��xĐ+�Flu!3]~r"Q7С������Y�Oq�-�Xu�j����I�y�;�/7m���k6!�\��c�(��E��冀�Y��|�HQ_2�^c�㵽E˚�v6�d;^LN=ђQ+c�\�=k/ga)8�0 5Gg�f���:r׏�~�Z��!�h	ab+ �Z�ǖ�Mԃcˈ.�FA��WGvno;�=fit�5{�9:�����TR��;Bw3��!���|���X��n�6���U�F{�)j�������^o!c�zx��6�l��%�T�:$�Q���ެ�B�x�r�燼q��)���b��C���?�Ď�Gw����a��~�i�䳍�4�_v�ؓ4���R����}sG�$%��K�O�d�fV���X��(Zx�J�f�B�Mx\���ftRl�{U٤�e]'v�q��-V��E�7�x�+�|Gl��f*��z�#F��%IJ�uEB)�m�I)4���J3\?N�R�챙,�̙),����/}eko�S���������2S�B�~"$n���V)�P��=F	�o8��m�DE�E�c�>~����؛��5Q��+��>()q�u�l�6X�I�m�I%\G��Ύ#�{R@�S�S�8�g�ۏ{�����8�HI����;�?���v���iT	-���#�b��Q瞬��@5�ۻ�y1��?7&̳��ǒ������~���B���/P�S�/R4�Mz��Z��;%�8Sss�'�U䴱���ٵ�5L��X� (��@|#�|�g��lPUS�[�"�\d�t ��P�4��N���$��$v�X�T�Q9�*gg���ϰl��r{K�y���6�&�4G��rD�lp���u�#�N�P��.���g��U~��n���T�,Iŉ�Y헫e��M�T ��`�^� �jXw|�[;O?�����A/����N�G���2b�%�	�dm}�����P%v�J��(�/Hf�,�M8�<d��\�ܳ9��v���T�5w��v��\8�*�"2��v|)!�7
n��A��oZ��jg�F�U��}z�ù/�ӽ׎eB%(S����2��I�sr�Ȇ}����4u���N�\G�α?z��=�Lz�{��n9`�:^�0��H�[Q�\,=Nl�,�u�r��Y6�9�%W�
;8�u)Q_�=�C��ɾ,��&L���̽�zz��d}X���)l>���'[�o9��+���"��t�@XV�a�s�龫���Rgl��z�e�׭Q,�'8ڂ���W�O�G�$N�/�;�����˻���vx{l�\ʜ���_�i��y�l��^l\w�'H���x���A��~�~���'�T�l���ҩ���RÐ5�s���\a�J����泞@}Ɓ@>������0=��5�jpJlB�u.`�F��\j����A[�e���y���DV^<����tm�e^ֽs����l�A��"�.�-
�j�^��Щ	�~����	�Ϧz��=���M�������4e�'��?tu���w�|��ҭ�;�ܶ~~M��$��8���F�eD6����
ovy�8��j;ʅӍ��È��Z�9h��F�9l�ϯ'��Y�4>�~�1�/����!�P��7��1G�4��}�ř��~����:3�����Hxy=�P�\x�A�1Rپ��J$q�C���O��R��uVHa����[6�A��Wv�����w[o�9��/��}�E�Y�PF�&c2Ӻ��R��㱐�2��m ��{0I�[�P�9.H�"u��[x����s�k&��+�Cr��*J'�J����+=j����%M�2�( 8j�	��.�\����Wa��//#�G��t�sۣ}��X6����Z���6��v��X*s0TٛBM��֨��6�v\�Zs��r�<��@VK�ǰk˩��-��$+�h%�/
�xN�h+r�K�R!�ٺ1e�����sv�&.����ɣ����.��L�x��l�WI͘7��<���Ls�5����%j�����#rٙC_$��i�$D�,l�X�)݈��蘭mn����'��iڳx�;��&L�[�z��*�\�!���6�EL��=שx�{�1�#}��� ���)��Su#v�oCd�_	t.�#k�lue�B������x���-�/J�����1KT�sn����3Y��c3�wN)�Σ���8�|A���`��΍w]o�V㓫���-���BG ��$�-#�� H���n�^�xڷrX�%
O.��,�t.��n���ػ;n;�"i����a�2��E�*���C�N��$k%�b9(�D)n�!{a���zu�q�6 ��D0lٳ�� e��8彯��+�G�"i��+]�;��a�_B+�B���<
T�r��U�\=�@:7_}.�^E��2�v��N��a����3)La�Ld��ON8��Q1[�����)S�;ۮ\ݺ�9^�r��⚱Z�QS-���v��69>2�TU´�hj��;�p�Y"/�CN� ���0Ez�CЂk��]�)3He�盉�6�Z��b"�s2�է�(�gi�.��z��\1Y�_N�TZ��{ݜ�f�%�M#�3�ړ̡X��"��S���SWՒ�C�^��sZ��;!���b�1l�g0c/n�탴V}|k�ʒ��dv�k��-Y:��N�y/��^9Gt�oA=):g�Չ	�c�TAۮA�pgڗs�y������54���;sL��\k���o;��)Ç�V��֧n-7��{x����N��Y�
�n�SN�ڱ%�����;'KC[�PuwL�ՙ;��IvWwZ$��1��������蝓qf+���r�b^Q1Z$p���l��k/u-3����>}ӛ�V�[�2rv� ����Sc]��t (^<�)*��,Ab���$�VU:�=�~�z�~3���||z����ffs33�s�N|~?/���[лf0�Z򒳉�!m��+�g�������%�g�^�o���Y���L��ffz�s�������n!��H���jKR��,�VK,I���9�l���3��ffg�33�������>?$��U;kX�>��
���/2�y����?�뙟��||z����ffs33�s�������[-A|e�ا�T֧�2ֈ���ze���"���st�N4E�a��
ċq�/Y�0�F;�1"'iE�WX=@�1����� ���<gdq:J%B��eW&�rƶ+�jIY�5�/tܠ�PX��R��2�M ØҠ[J֧��)�5��rb�Jue�ܳR���1��Ƣ��PFf,��=%nN%�y�Bd���R�bM��\�	p�*p[��k�w��ɓ ɓ >ݪ[�cZr|9�	�Z�l2U��J~�O<��}3�-i�2�8I�-7�^���>�������-M�5^��ZN�bS�(Ƈ�~N�z`kx��Y7Iy؇�ۺ������Wk�C��IXȜ����4�Y�1�̿��8�/Aއld�|�%K�;P���@;�G�y�}w���U��E���o �Xw�����UV�T����	�b��Z�t�
��xJ�l?~�י���Ei��$�K�$�C�{H���\���
�z�E�8���t�Ŕ���=������ �ܓ���s&���{�+X�鸅��t&�m��4��H7����k�ܟ��U��j�M�v1���ڳ����X�b��V/��*�v�g@T�j����Y�S��}�t��lR�ʭyapKM˾�jv{����挭ׁ���1���{ky�v��.���^5�e�#X�j��H4����	z�Q,��t��GFnH�y���n���"�I`,���q��|F�n��S�����"�7:�y�uT �}/���="��Z�8䟵�y�a�,l6���>�4���F�u��Z|�� >�S=��r�O;~}L]䚮P9R�K������I|�s�W�GS1����jÏ*F<.��qO����),���,����^��w�t> #�na޹�gh����GP�+�~8t ��uz{���mT2q�^��!���_V�Ԭ܈lȖ7����^��G�jl7���~��M�� *FN$My��1��y���l�:�{��.si�����W~��׼��n0�Pga��9ފb� f|���Ie)��t�;J��jj�
>�y�.�k,v�����*��aw���G�=鞽8��S�ڕA��/$km�FӺK����m��ўjo}r㟠��ٱxp3~�}#21�2nv�M;�Y�6��|؞�vy�R�"+�Ȋ���}���k_#}	e��;� ��x���;Fk�n�z�gL7���=t�a�{*Gwm�ˇ�;��^��!�aq�d%c�����{ c��b�wG�aLt�]k��F�l˖��=�W�m�%�7���^^����~x:�nRQ���W鵱�ݝ���*�[�N��l��� ��p��s|�]���vY�!�ؚ/W����]�|Ճi�� �͘�V����rs��e>�r�.����E���4q�n`˾3S8�xn��U����rތ�Um�*���e+Lu�֘`��`��2!L@�By$�N��>s�k���)�g��%%�Y,���3�՗�[r	�Uw��oF��c��l�R-BJ#w}G�ￅol�Q�:U�x]m	%�P�]�A�(Rb�)Z�^G{&�=�|��:2;�娽�wx?xC� �m��S��k�����ȩ71�x����={��k�!���2�\l)� �1�5^5kc���=W�����,\ �<��;��G�{�v�TC�G+=���zwC3g���pm���.͇��+��U�tF�DՒ�]Er9�.iӝɧ]Z�S���v�ss��c]u5@����O.
�c�����9��8ˁ���#Z���F��l��qՐ�UQ�GF�UG;��̼خ����p.�j�Ƅ�;c�q7L4��� xF���z�
Z�98��b��eMI;�6B�e]��՛R|3������|�r|I�:��X԰W�D���5<���u��Ӵ����A�8�C���RQ ,�x2�MԶ��n�4������,O�cF��s�D�+�Yn�e��>�yg�u7a|8M�UF�"c�+�=DU{����g�7k8���<�.�r�nY�Ԉ�]";��]>�=�j�\�?�<|k�����3���2ny��������B�.�C={ِ�6�``0=M�|�l��H}��n �ל�����\���]�U���ITM.���m
3S-���_�79�;�r~�ÿ-k3q#�>����c�-��G�&u��X��=\h'k��tl��E�p��C^�{wg���+�{h�[9��Ϲ��g��}�>��B�[2��{����ԉ��U�Y��!� �a��Kf��g���~��w��PD�;�H��*���Sv� D�F�Vnw��9̹[h;�~�(������,�lF�Bx�'.S��J��������R*[�}}������(�D�_\ǚ�{�4�\��+�#��F��[<���GS��o��}�v�p<��܍��x���z�/N;�!z����R�����Ր�+�(ߣ���G'2�9����ǒ�izb6C&���xN߬� v��t�~A㗥fUz��ۤ�Ŕ�I�Iq"���=���sy�v�*( �$�PꬾUc��]�=���|�>�Uk�C�k���u��7�^񫷦Bυ�O8�S���t��T����y;��t��^��
t��斆M�ggd2d2d�;�����Ȝ�b�i�S��^kg���y�(����w�b�^j���`u�j�I594L�5ͦ��R�AD݃�Ax��N�|�*��g����	U׃��N�fHD�����P���_*���g�O��b=�/��e�GJM ��'��LA��c��)�5ੳj�!��d��I�-�i5!���0~(��B�o`�.�bz����0���;m�u�הU�����銘���p4l��1����ۙ�
W�����=	��{��"�/ٞ���;D>�������K�)����`�J��w���^�=b�+�~�Sݩ:+�5��Ym�v��ϼ�'��.Pq�{lǰד�)���9�n�a-Һo�X '��6G<�A��闶q�<�y�^���w��u����&]~|��;i��w��W�p�r����W���̑�X䬰��Hשk�N%�/��l�Lpb��vN=�b=җt�#�x�P �Ħ���[��̹ZUd��2�X7������3�Q�3����ʒU������j5�*��B���K��v�A�&A�&A�&L��z��R���uk6��hG	��I.Z������u.��!��VףҬA�$�ŉ����r�St�77vn�ֽ�gh�y�N�	��[��q9�=���X&4��"�O��܊�X�APA�H����e)j͌�g�z�t@�Aih�[��_f�T�/zc%�L�jZ7fۚVdcgU���)���vR���L|��H4 �ڿw�E�/Ӈ�}nq��|v���諝�^��fnM�����"!l�{zo0�L!�Fso����N�њ��W�-��kR�]���++5�V������y��yǇ����i�[���W��S��#oe���0o�l5����E�:;�������|��|���z����X�B��V{b�ۂ�{<�z��o*�Ҍ��VD��z�kׇr�-��',uoE[m.b�#��ǰE������j�=�O[�t���6_ԫ8v���Nƫ�^�;�ㅅ[�|����\틍C�=x���e�:�W�@��t���5T(Tx�C��!rbQ�63�*}(!�e��m�A��8���wJz1��G�K�%�4i��m�4����b��,�L�7�"(6dH�$��|���t�e���Ԥ��K,�����γ1{ÿ�Ͽ������wwZڪ+�o��p-~��khkpV�0�7ӛ{� ���댩��̞������"��||C[�h`d���g���l�����i���fE�	��,nQ檡 ����x7���&��� C^כl�GS���ng���e�ژ��w&��-Pz,o5�X+-���}`�3�z��������峽q]��cz�wL��b� q�{���H�z[�o�R��UW>Uw�_2{�e�9n�ݻ�7ˋ��|�8Y鞠p!��w9^�֜���������H�퍽�U-��k�4��=����|�s:7��;ݦ�rjv켏v�� ��pnɺ��_��#�����?�Ӂs�Q�K
�%��� v������j�z�=��wL]gyo��2�zhz5ZI{2�ocS,���in�t��� �i��q�����'_n�ߒ�ģ�O�_.U�Fus�n��G98vv�)��9¾Up|UjU�NU�Uj�lf������Y]p�X��網��uՏU%t��wЃ��Z5{��rKޓI�,r����w��yyyL�L���޻�eo*$ϝ��鹾�2��,v��wvU��M=���	zf B�Ⱦ��ޞΑ9~~��|��* �Z���T�$�����5wxI���x
�ث̏>��2����v0_{o&4 a$,��>Ή�O���U��op}ҽ����7�A܏B�/�Ȧ[��\?~[�G.������R�5�z������ΆƐ�h+����ِ��?oL�f{?}iP�o��ͅ��C]�-(wCΈ��s�Ty�V��9f�n<����"W#�S"�I�!�y^�����Jn��^�y3���ݮ�3͋�^�G���s����vy�[|���u=�T����z�=9��;.j��YT��o�vMy�h�ni���6ڱ���ҧ5I����H�/~�z�9����t�[����l�gaz�u�6���}�8���'���m`�N=6b�Q�����ZϺx٘-]bo�d�k渮��{w�P��|��&v�g�t����`�Գ%uZa���MVⷅ��Ej�U�̽��.d���)����2d�2d�2dɶ=�7x� �����)�㔛&/<�m���@ad�"{��.y�٣�/���86�N�e�e��d��,l��;=χٍ�o���,�ދ��Y��q���b���M��,�y��o�%8����4���/��2�o:�
�4��l����,���f;mQWX� _v᯴�94����/+l+'f�L�`i	EY$�����WP��*�2 �"Q�-�-�^c�}�%�:��i�&�7����S�s�?�g�I��c��J
�"�l�;Ď���s���h.@L�h{y�N��&��z,rox�)��By6��[��sv�/aP]�v��iΖ�lq2���ȟS���w��M���L��54�މ�A��2%g�m�=�S���g�@�k#���*���^EYݡ�Bts�� �Ҝy�Zu=����ϸ
Y}]K3����NY�x������K�	���w�+��R�iH�2��ڔ���43Y¦ݮ�8��
�>��]��^�����flo�:�g8�X3e�M�c��r_i�z'3�M܄ŵ5�!��[�{�^�zjg��:�,�fL�K,���E�9�/}��]���45��=�-�'t�C����߾z@�g����j��K�U-����B���u��n���;� �I��,�y�?h��iQ��6�����vdyӺ�O��	;��3r^�m��i�����7P*3����#}չ����R���\S����U����#���]����_��g�<���߽Oٸ�i��z�N��Pg^�&Mu��": n��c(?X� ��ˍ��n޾�*Ɍ���y5���s׏t>ntk�uQ"�9S����6��Aǟ��"q�nfG^rȖ����&��}#�:k��!D;z}��y�'����]W�p�5z�!�,�Nv{��עg�T��>.�f����k���_U�K^1�k]�k�r+g�n7��Ij,͏{�gq	�74��zL�댭�&��ހ@�s�!�����5�v��+[^��}�?:E~�FS6�Z�sT�L���d��W���g�_[��
�l�7G�)�N�*=�b��F�z��fm����^�ґ!��u~�>���sǴ!Η=OΥ�f�dξZ{LP���[�[pvr�GH���@�X��èsڪ�r,��g����l\[�4��x�w��wX ���ã{cg�y�A�/p��3Pf��$oak��`^�C��R�,Z�n_C��=���EWAH��]l���O�`��G�ތʊitq܇���4f��e(����lC�{/Q��r��n�.Ϝ��¡��xc=���g��;O6�\*�!�d�A'�Ku՝�w(cF��h��3��0��V��5P����m��镵�Ժd����=�sc�m(�v[�]k����:�9!qLO�&;'�ͺ�\N�u�F�f?b{��9��"<�y{�d�Y��R�1`��o��8��#V�m�܉�O�H��I�<�a��.���bP|�W/�Wú#+su�n=�x���F��Wo��ǱDu��;79����+�)�<*5�ܳF�{n�+�NR+����5��WJ��|��]�A�hJ��Z�A�
�
��p�6%��;�k�*�����`��+Վ�K2L�*H�bđ�ZE���;Ӯ�:���cؼ�=�,���|�HY�Ix�rSm�S�sB��2��v�/;���YwF�ߍ3�*��F�Z4��Ro�I�ڻJ�ȁ��R�
�%�l�����C��0gB�6�e�U
%T%�zj�A�+����U�+-T�3JFbۥ��rU���v���{����C7����yS  �
'��7r�62��uF+ �vչ�:=%�R�U#��W�G6�mG�6a�����w��W�("���-�˥KD�έ#Q���j���j�1�}8TǴ��w3��N ���1ٯ��ݽ�r��e����EbH�f�쭊�{��V�/r9�w&H
��tZq<@��n`���싆oJ���v*��t��Y���qnW��ۏ�tj��٠�j�l�scY�_Bn���i>�7��#�-�3�������sy��=\.V��s��P�1p��^�Ծp�XN��IԹ�J�Q�*�fd�����c0ɬr'^�5�acY�Ȝ�.qġ����Z·7�ms��iM���\�q):7U�w_VW���:��� �m�L��m�X� � v�5gz�jUvM�jF2`�����d�Yu���:�u������)"55���4�.��E؉dRV�J��j�]Mޞ}������]�<�7r�����'a烧3o�e4�4+z���u�hw-�ӳ&�r�)v6Y&�$�b	��)Ⱦi��ܜ��9��$|)���9w�(_�ZC�B��L� �n(DBV���\3�X��g�)u���3r�Z���-����e7V�]10�&�H�%��Cm��()e P*0�a�'A.u�$3i�R���"� �p�j��T�3�FY����T^�@vĪ��,،��R�wݚe«��m���d5���$��q�E�SW[373swn�UѸ�<���di����}mj(m�#�P�<���q-�����������~���33>��������>9����E"̥'nȆ'̾ޘVt�+#מ[m-��O%���^=}3?_��|x���϶fz���s���|}���y�P֮^m�~�18�[W��娏l>C�E�D��ǯ_O�Ϗ�|x���϶fz���s������u��c��g�˜eq�(����V�e�N^���>����||x���϶fz���s�������α�~Y�Km�<=f|�/���B�j]��"�S�(�%N$��Y�Me/xoP�84/tu���v�c\L|B�v�6��fS^h7�*�CƳ���'ֲ`ΐW�w�P��f'{�,.�-�mE,�+@]�Tז�6�w0���++1���N����7�����Qa�O6���믶�$�4+S�dzL��e��i�N-�!e�j ڬ���GcY�����z�K�G_j���x����������q�L�:dx��b�nm���$�
%�bQ�;��Қn[�i�\6�Z�n`���tsMܮ�;�Q>��RY|���������vk0�_-o�r�#
1��P��V��I$~��o�ш�����ߝ
�+�� xr��-�D����i��W^)ޝ���M� l�
5�j�q
�&���uNw�y�YS����/��s�}����EsC,鬍�5eK���w��DJsb�E' .�����^�p�VXb=u��9�P�C��V����H��Ɓ�I/`L��KK�����i�U���)ɜ��|���'ѳ=X�Av{�V��w O����3�0�>���ۍZ4��2��k]��ZO[Y���-m�_���^�:���x@�w������w!*�=Sw��_=�{^���ޫ&�Ft��=]�o�3Lc8z���H�c�Ig��#]�6/RdV�3?t�:�B]:t�
7�W�}|���<oTn����)���9��rF�pǳ�/#�֌�q^���ym�݃����8Q9���M��y��[�	�����:��t�����δs��v�y,3r����/ES;��o.��S/z�O3��xQ�P@��:�A`;fecV��y�4�	$�}�PʦT�UG��M�*�K�ӻ����x�Ü�{74�2��GI�3��E�Dv��L�~�5���^>L�&L���]5�;�~e���b�؛����Y׳`Zڷ�6�m��_���z�s�����S43�3M��E?���%�{z6��~<�s�{s������� ��t�Cft;��9��(9X�v��cOW�&.k+��I�]��-] �`��g78�M��&�<��g;D�T�f�#��I=�ύ�ll&OZ�d2X\eh�!1�he0(v;<4�����8�z���^�y�S���wm����-�->�k��Ӝy�Wi�V��K���}�s���Y����0�PxW�>x���X��w��Ty���s�ee������h�B鰾�EM�O�r�!G�O��8��*gf_x�k�v�|ǋn��sѕ0��X��&��ݚ�S�@�	1P���)C�y�g4��i�"w���v�"��J� 7��{��߯7@���y���30��iY��խ~ʸ]z}����}\��=[ϦŽ"Q����W���g^s"��v�Z�v2���Wų/���$m9,����@�����;z��0,an�,�m+!Χ�ʻ���j�_X�ēѪ�5fN��{��2�s���Ie��YIe������V��c��:�h�o4���c�e�z���Y�x���Xw�{�}��u{��ݞ��m�����'z������
ה��w3�Cގ�X�]�	���7˨�i��k�wr6����Z��&!uDb~U�/o��*wf�q�
��M��c�=�-���Y���Q����XI�8x�\�{v�<�"��H;tp���~�hgC|�����q[W�v�ީ��gh��_n�f��)����j�l��}e%��2�04�EK�}&�f���i�k3bz��[��kh�x^�/���s8;�{1�� av.)v�����^o�LN����i ��B/߮v�����{V�v�����8�r�}�w��F��km�g]V�ǳ�'��N��3�=t������g8�|�6���n�!Ӑ��m�7�CL��zA�ꂘ�w��8�����,K�m��kU��j���`��a|�	�:Iu¥T˫����������3:	t��C��g���u����^�+V/��gj������#DTut����a]��wK�g��,�Y�3&K%�Y,���w\��q���1 h�Z��n{��hV�pM'�y��ؒ�'��*�7�cr�u����	�Ϛ���yǏy���B��ݜ
d7����ɿ��@( ,��VIV�����7Ǟtn{�צ-bϘ�K07�犍��Mo�%gK���P��r{�7=��OR��1q���p�f�8�K�����~�g.�ķ1\�3���󊌈oX�|�<��Ms����j�"�i�����^��F�s4�:� {׎�R��z���y��{�6���وޔ�a��DTת.�s�״ݭ����`��:G�|}�w����4|�V�|��4��q ����Swe��������aUQU�}�%�x��6��r��vPY�z����i��a��y2Ԛ2��i�Ee��5�G4���v��:��}=��+�k2 zoVm�uӵf�m�"j#h�Q�α���;7Rq<<!e����<!n���eU�W�]�Ȧ�-�-�:�7M��~�Hx�W�0+�w����=!ؘ�߽�Lk��qb�^.VL!
iDiQ7�|ŝt�[�C�X�a�"
�"9&�v�M�ݙKC�|�h=R�9MZ�������\b�����
��xk��]���2-.�v��u�5GS�2�����%%�XYIe���'y���w���~��U�'Ϙ�&=�}�fu�p�U٭��͵6(kH�e�Ϸf�3w�:++�M
�6g{@Bg"���8cj��l]�j�*����o��:�xl�mr5o���"	�� [U��O��z� �Y;K�Z)y��]���F7(�G����CZ��E;t��^��V�g1wE��UN�{��:���㎶������h~�Y6�]��%z�2�#f.�׃����بk�/O4m�7ޖ�5��T\�����7a<k���5<�zyVe��F꺫e��'
r��W  ��`�r�{\c��T�zqv[�9I��<��p��3��l1��љ�����p�^�`8��_���W��ƈ-��e �E�_���nn_]�E��-W�K秳|�4Mc�S���ӱ��|����s=������r�tS��'x�v�ݶx�0���R#�������>�����d��V,���v:7�5�{&�$~ς"s�x�?��.��'�<ȯ�t���̿�L7��=���qP�y��߭�Ã����=��bOx�!�8b3J���W6�9�eJ�����2�2�2o���#ޞ��6�����������S���?~{rN��ɝvo�_&�unc]v��o��ޓ�mx��]^��U<A�����yUf_Sn����y��E^���Q�2�~�$�i�����`�X����W�yu!�0l 7|���轼XE��y�7����V]xt�FG!�S�ᕙYE�uK��εO�Yތ���Pپz��iS��C�-Ve���-�o�� ʹ@�ZKdڨ��w��Jށ�^�~��m+Ȓr8��a×�UM[�7�H��BZ�lE���(�{��1�v֮"�'�ֺ���
s+�z×@��U�w���T{)�۷����-�e��c\��[U���]�yB�^���͑=��	4�gN���l��0&w�V�mdu�Bs*.��p:�g�̖D��]S�띐�}�r�E2���F��C�z�+����fsb4�6ɨ�O���e�ᢉ�t(�;�����x�)������}b�$<H~�b��D� Q��p�~Ϲ�Q�d|�l4�ˏ�y�"9���ô��wal�&eNE��+L��Y?��^A�&Lɓ ɓ&��_n����5S�����<��m~>mv��!��=;�Nl��`�/j�%ǰ��^� �{n�x���8�d��z���S|��w7W�Xwz}۷�ޱ�Z�oJ��7.��D��.Ӿ��"�yǹ�!�NU�v���]9�o��=Y�󼓋���c��o=zc����K7˓���������������
qiQ"gɅ���=�(�\տ��g֓����o�'_���{*"�j��/6�㵮�Uzw�F�=��=���:�i?��Cif����( ��'3�jm�@��;�)�z�ed�|G�z�P��;}&����/
�z�V�2+2�5l.�=xָrą�-T�$�)q6���;^.���%+��c��]K�r�Vr�xg=���h��~��#�n�tP��������w�E}7�r�r޴�7W�4�O�=q�ʝe��]��Ѻ���aQ�7�)�/���I[�]dT�鹭w׌��Ю�q�̓��1^n[�z"�.����;����>� ��$1����l�j'D���u��;a���&�;�ć��`2��}���Y S&v�T�G�����������d2d��[�������Vcf--�,3ņj����2��������stpBR��C��bO�@��z�f/�We�v����E��˦ Ы�7�g5-�tJ�~��g�.��Ⰲ%�X�0���u�9��zn��u�46k��fKnA�������`ۊ{v�߈��8���8ʏow3SI�t�#�Fv�bA�E��9�AV+�Y��"(v���r���Y��H�r��5y��x��Fs]�}�Sǆ7g��q`��U����z׫?}f�������}r{ϧ�pg�}�O{�H�q{�/<��:�Ȋ���m�(@��׏g�/�.W2���mD����ۄ��h��^��p&Nw�p���
&�ʹ���}\ϭ]�C~~p���׻7���i=��X�z��$Q�1�U���4�w���]�N�}��l�q���׼0�.�������s�]M�ᨃK���6�����Oo�(*���O�
�2]���T�I�Ԇ���L�GE�)�Pb0���ǕL}z&��hii3�[7�r��9���m�X���P��+�='gwRŻ�x�����d[�?�	�@k�%F�EF���m"�l)U�iS&��M��s�����K?�%�P,���,�N�巫�.���g��'���3eH�T�&P ���[���_y�� ?���{m�=|7Ԫ,'���6s_z�^��<�MYr�X�k͜ox{�< �91����{$�>�k:kw^���-f��}Kvr������Wo��u�^j|��q�Gm'
l�t�M뫺��7�];�vtk�uQ0��A��s��{��(W麳}N�o���}��z@�"����jk2��������QJXT�����c�.��\3[��O�km3��W��mx5T�S������Y��s=��iyDf�@u�{����#���U���酏r~Sϑ]s�w�^d�4�]��@��B�2���	�v�YVv�.��{�z�Kƪ����U�� I��:!N��|#ag@����J;��驠oy�B�Wk�q���:i���@����y�h�Q������襫f���%n����$��.��X�f����ϫs�{7[���ȩ����q���9zЦ�S�SO����_;z�^�-�f�ܻ��yd�_�Z�u�0�YC��cKB7+yID���}���=l�&L�r��ɜ���˲%���������ǀ�9�8���:8��)t� 0�
��~���p
��@�tST�D����W
�&�H��0���e��j�6��+����E ٰ�""��6^�����R>E�l��M����Q�ٿ{�"�k�s�9͖��H#ۛ>v�.���Y�fa9�Y�N�����i%�,"*�,UF|޽�}���Y�\����w@�UqRG2���UO^v�-����lfOTzbS�y��}�l��7����P۱�2���R��%�fN.��z\󛆉�W�ٯ��HFHM��,�M��~MP��76�U^��ި��[<�g�Ot'��Gf}����Z�������= `���q{��~�O�NmT���ه7`�1�4\���{���o�����e��2�
�����W�U�}ʰ����7T���\6ߣ[.À�ױ���/��_k�Dә���ǵ�4���=�����=�q��B��W�Ax��M���T2*۝\�-@mn�5%���(��{�h�i����}��l�C�r�W<�H�f�KkH�{�
]�P�U	��Y\���û��v�uud�$DjL|+��9�A����3�y�z7�]��E6�b5�lI�txH�N�J@���U���Å8��pT�f����F�=���O�[ۡ�����!�C�gQl�������ۥ�.�n 9>�j؊y��h����1�2���۲ft��iY��9%��y�1���b����Y�S�����zsj�\���Ln��-,k�͗�yԬ����r9��J��u�66>ƦJ�4�q`��ͩ�N�Mv�E՞钑���>]ڄY�dg�����4������Aˁ��%�Y�
���]C�n�,��f�*���wu�1X��s��G����*�կ۰!�h���U�x�4V���S�M4 <�oEk)!LL��i��L�n7����h���k\���wC����T�DPB�B�uu��jCS��Ǖ�<X�9�B�5z�楎P	l솖`L�Th�X��^{¡dt\R��B!;X��o>�*�����`}��1����	ʨ۾�:;Ƿ�oBN`�ٱ�bt$YD�����@�a�.�۝V-D�f�vZ�ڹf�������b���5�׽S{�����k�F�Fa��|��ک�o7��%,lŝ�r���7�*�~����tu��6{$��Bugh�}�¯u��_ڝ�\��V4`��k�W��YL�y��4��O�Ѵ'o��MTӷ�Hq4L�Ĺ�d���vb�b}�fQ*�e����W���o	���G�'����݀��͆/7���-=�IMRy-S����njb�R�%[(����L,�l��&B�܃UM���E�<�{��_u�뵮�^�x�����o6p8�X��N��=�[k�8h�����f�E�|MG;{�]�AǫVt�[8!W�v��N¾�6D��v��r�r`� �;��|�f`��I��K�,���������It�17:Y}2�^f[�6�k��oS�d��W+�qb�����>�L�ݦ�午�qǖr��{�8�L�wqZ���WڦEY�f�@ƭ����57[�E|������rsWk��>��!��o3YOZ���ޡ���DYU3�J��u���K��)L�`k{�2d��ό���fffg�3=ffi�f͛>�O;���q�p�qS�1��E
�J�j�~l2�FKi�c�qZ�&L�6}=�O'���333홞�33��6}>�������O�� {q��J�m�����*̡R(V>��O^�ٙ����ffff~3<ffg9�s��������-��B��|�t���/�y� ��o�O'�K|�O+��Ǯ||g�~�+3333��339�s����o���qU��f�㐪z�����Y�@Z��Q�.*�jV%��~�۸��!�5A�,R"s�LԡX��7rFҫK`���qԩ�Y"�"%��"�E�j��-�� ;��u�h��**����;��5LeE���F)�q�e��l���1U�J��Z��QE,��/C\
�&8��bo2�eʸX(7�wv�`�H��:�"��%h*�(��8�8��:�l�Lv���Eo�o��9�˥�f��C_bA��-�lN=�nj<HTm��z��+���C�fL��YI�ɒ̝{wu��W�y��~���*j�޸e���@��;��ڑU�}���W�y7}��R2��g0��H�}�{�Ef�\Ha���s����ٲ���/`d�BGg��c������=>�8�p��j뀷�0mK�6��9ѯe�(.��R�����o4p7�����l�~��-�4GgC��D�T�!9�@�f�8+�^������3�unn,VK�r ޕ.	foW;?iTӝDQ�l`L�{}������ۯvF^.��b����%�`(�a��畿�zg|ܫ���-�aRz�>�Ί�Vu]�j�<����`s;�e>���m���O����K����Ϙ/:^��J̎z�y���w�oz����ŝ����o^��/M�D����k}v��v��~��_�U�X�\��Ι�7����E?��w5XzA�l��t.S^�N���v�#�Uc��: g�mx"5S�Y� �#͋wzXc�_tL��Þ��"E	�x0:ɛ��$��B�,٭y��[�ue�1�/��'��gd�vvA�&A�&L�s�^tow��k�4حe�:A)�[�vv�n�FF�G�+�P��Q^�{�>�>�C�)�TVt	�:=���;��uv��ދ����8T˻�ߺ��l�# n9P.��b*|���՞:�(+`��i��v�cMDB����ך�n��۶�>]{g�y�i$Jc��oð\�������z���o3��$�l0��c�ֻ���>��R�64d�̕4`ݩ�Sh�[�n�9�H$��_����v���Z�l��*��3S����X�{g=��cm4�Ƴ�|��M7��5�NU{w��#��5����D�j�8Q�#NȞ窡^�jκ��z�u���������v߆���0�D�(������z.�sM�^�=Ǫ�F���|Q]�j�u�����c��<��x����z���㙁��ge�'4�����/��A�\~�7CS�I� 3���i݌��i=��;xTӽ��\����V2�	��2_wK�c��s,���!�.�Kx�&a�.�U��x�J�R\�G^�|sq�u��L�/j�n�I��c��1l�Bh���]v�Ʒ����U\�U��&?�ӹԡ�2d�#2d��ɒ�D.�8��8w��O�(q���DF�*C��@�T�А�o7���}�+����=�B�u^�]�4\�p��;</_+�@�./h	h�����v��tc]�!o�6�㙢�nQo����lEi��7�#��XM�x��3�}��
���@�O�>�����dx�Y��:����);�y�7a�@ܾTb�G��͌���>{�꽔��r��e�r�s�Ƀ��H�U��{�|�Z�{.�����D���lS\VYk�	��5K��Ώ.ª��1�����z_ͭ���|�m�r�HD���}����c�RlkV��l�w��N׻�6�Y�]���.�ިȿ5wu�P����Źk�` ��:�����C궅o>�W��'tH%�tM��MW�����--,����--�^V���ћ�F�E?���3w�/m��CC�vxF&��]����.�ݱ^�ղ%�.����-���Q}�jt7�
ܺ�F�d��u#��7/6[�a�{n�ؔp�i����UE0�5Ɯ�A>�ߍk%��9�0�	u�=�[Q�i�.��
mӱ��4�U�EU�����|}��/3����;; ���g�]�}���s}��[e��GwC@}��דY���7["�H���>}�����WV�f�[��k�Ed�ޘof�q=^Lk���U]����Tl�>B7�+(�y�!����yr9�r�}�w{z���9�#���C#�s�8́������2�=�۲�ϰ�_�.�n�c��E�@z����ē&e�Ԍgݷ-�>��+p��$	�bA�۪����Vkӓ���	�v�k�`B�.�W~=�A�|�H��Ы�x����1�	j4�� ������3����ܱ��[���;n��XFk����z�33^�ͽ�w���.Q�;w�F7�ѭ���9KDKRU�Ǵ�:��b�vf��g`�1�\Z%��vx̻W���Ut�vy��}���۫�K�7g͉�+�woӛ2��u�i���J�!��7>k�>x��O[��A��E:�ץ\��T�X�o�rjR�W�V.���[����Te�c;���YVE��F�'�����d�7P��[ꊦ��sL�+]b���|]�)u�?������޽x��^�{�׏d�Զ*W�{�����<�������$�>���l�
�x�MQ������������z�/�N�q~k�K^�]�X�Fq�q������wnJ���v~>[��
v=�j%����ۍ��_y��ת"* �oF)�NW��|�jh�~��rjD��b@�AI �֝�>�6����S2���~W�4��7/c�h.��de$D������Ͳz�z�P@�[�'�;��@�Oz�h��]z�ۻ�~�s��vξ{3r�ƤJ�=M��{�iW��wݰ�ՔNn=3�F{\,�5�-��i��$����� �Mhf �!/�9Oy^�ǭ�V5߇�D����}��צMyS͸��n�E�C��vka���˕fpgy��,oc���]bD�ϧv�#[�L�aP ����׳�۽ꆿ	��[���C�z�g[V��C�\�z2�ք�W�!S�[�XQ�b�]-J��M�+�푈:��2>�9|V�75�	��M ��x�E����e����c<�\E"��HTTc�g�w�jޛK>��'M��Y�p:�q�懴d��<�*Iʅ��*��6�2g���;vvA����g`C�w��}��V��6�m��� ��!���wSz6�����y�Sȼe�&�����F�7��9�ש�|���"�\�K{�������I�$�y���Ϩ� I"�K,H%��ձ�LR��F]v�4��6Ƿ��5sS�����?>����f~�+G��Et��&�����=��[�}��m�Y���gd��֓�i�?t��-�q7�������L�/�h>H3E�EW���G6��n<^�sJ�f���6���o��x��8���^�ǿC��mj�4�j���֚��,�l�5=(����Cb�U�E\�������{���N#7�Zw
�˱�?+:Z��k��>���\ގn�h��Ώet@Ӥ"	}�s&L5�UNHp�����_����l͝��>���G6�zo���v�S���������kܑX*Gs�II�9EX��X-1>��������"1���3ޫ��vy�^��D=)���ʋxe�7��7L������h�TIM"<b���M��Th�E�i���ȡx缃����m�F�.<�7h����++�\"A�gMˬ��ҏ�:ݹC$umDK	��&h� �c\��M���Tk�kv�v���\Ĺ��?����d�fɒ��%�\��^���}ϼ��yq��R�f
����������'���{�W�1�Us���G^���|�~��w}��][kH�a�KV��J$�.=<�fG�Y��|a���=[9U7�=���1�tU�5PV�˽p��D�dOz66��������=nCX{�v�oK��6�>;V�m#�Y����v}v&����]�����,��f����{�3��:�c-;���ڗ�]�%��#:�h�{�zj�Ew�>�hv�ڐ�f�T�\��M%�ڞ�8W����3�?I~�i���-O�{�����m�u�́UL�x���i{O�������boө�����C�����%�ϣ1J��횇	Ŧ,DiJB�q�!7Wvz�������dn;Yd;���z���W��`8����쩽�oe�o���2��w1+�H�w�������P[_���~�`��,�d��^`��b�7[}�w��P�W׷{�Ձe��=��,k���yY����8���^�˖��E,Paw�T��=�Ú��qM�s��&��ԟ%���VV�����2 &L����� ����]�־���2���T���lw�L��"����ܚ^��z�5m!��������.E\�X�@V�u�lFa���Wuj��^�W�g��64gN��y�����*��s�"Ȣ���W�Ooq�J����嗦�M(כ����F/w����w�;�6�|=5O����Wzr�(��;Ѣ�]km�H�m�h���~�g�ij���ކ1=�=���~S�i��	=��Gg�[��l�MN(,ݛ�D�R�6�x�j��6j��D�!�f���=���T��& ����ӯQ�S�	� _��&�=��ݵ��:>����Q��h`�_C	�8 VK@�d
�Vh��w�!��~�������¶2�ڹ�/�D�?�^�ڨv��B���ޡ�[���d�fO��f]ik�g�y�Qs�p�ꠇW��s���,�n��I�F!��u�X��Y��h��.�'I��#��6��/1�({���յ_-�#�C>��m+��Yچ�F	�g�cSK���m�ް��v��ܮ����GUc�6]*�\A?��<��|�����&�ggd�H�,�ެ�S�]��}OS�c3?�^k̏C]��M���C�V�m]�:�z�f�stlb-�mU�6t��Я���O;f�ء�,�$L���^{}6�:k��@ݝަ��5m����[���ߩ�l������w���h��㶁�iM;g��
}q���d��H���������R��G���>gU�C��C$-o���~6G��=2Z�,���E?����z�|鑹�Q k�J�|����Za�-�	�ž�^�$�p��om{*23�j�P��|O�������
�姅�P�:�U�׮�; �9ہ�{3ٛ��T�Y8�g��d}�5_�,��T>���O��M{~�W5��%a��4;�ٛ5��o�FO�9\읫5Mv��5�=�'r���H�2�����Ǧ >:�3&�7�- l]&���m��I=�8}��Ƹ�Ϙ��V���KM�u�z��yͷ�RƐw��iAr���+�ڭ���ie4�p�O^�]Y\%�y�DX,L�۹Y}J�ϼ/�ǤJ?�����u(*}�+�s��ip\�c�]��ت�ʈközEZ+S����ޟ{�������^�x�RW�^=�vvL�!����󟦟����"- �j�E�-n�o#"�<./�V7��*;� �����g�����̺��} ����2�@a���f���%%U�k���� �+��B�%�b��>��ٺmv��2���ZF�:��{�g3s{o�,}�W�/8{3���'��ݘО���w������Q�s��Iݺ����R��p�"c`��(���cj0��oDp9�>Uf�V6U�ed��Szs5��% ��	6�tN�}n4�j���ϴ��UѰ��L�ae�[�=��Mp��҅� ���/�}�MM+�����7��5��	���/ON�,ٍv��*l����{�gfq�/oP����EG]�J���*�oc�.I%�t����V�w�����v�rn���߽Yp=5yT�i����of���P�_؇o^���zl���)q1�m��^��o�^jO"A�
k�;o%����hv_s�ʦT�ݳ��P�mP���X牓V����ӕ�3b��@�U�Ue�f*�V���:�Ɗ��k&�Q�j������{W��莠Rw�%���z�u ���32;[�0kȸ�ޛh3Ws3w��j�y���k�[7s	�T�MQ�5��8�p��	9o���S��+9Au���h}:���H�w�ӛ��p.���5�(٩���yuB��Ä]Gځmqp��{d]Pg^S��R�Nb�`oʺI���cը��A��N���.����Ggt�n�ڴ�[�}�̴���H,�ژ�Z#���V��[�i�Y2���{>{P����~o�v�qL���*��.Z{\g]��53�g���sȳ:��:�C�w�wP�fn.N��c)�;z�>Ų�����2�v�Ѕ��3�U��s�C����&F�Zkk�����,�fRUݪ_[����)=��Vx��t/��*D�y���f����V����x��V�������b޲r��MI|4t��ղ�r����S��mX�c�>|�*�;�UJx�R|D9TX����,��<�,})��n:H-HC&\�n���gZ��}*���ڣ6�Jwl��2S��UR�cn�ͻ8=��3�Ե��wE�B�yb��T�pG
M�<]�f�wq�zU��x0Ĉ��6U�+�gRMH�JE��W�e�iS�ZC2�Dr[��a�nT��,v�}�/�,��:�h�0��"DB2*MYպJ\�K�I�1S2��\��j��,f�;�gk���g�@Rw@�h��ۨ��P�A3z`-�Vb���솹&�l�]y�����;0�z�;�e�0
 1��0�:m�����#z��^�xɑ�9A��vuWRRa�����t:]8��+��������:,m��V�����C|������X��Lޕ�pO5��$\�֧�p������;˻,X�Z�-QU�V��ɝ-���J��5-T�)s�^�w^e���h��W�{}��緈x���]#�u՝R�)�|�������2n���j�����0-6�|�m��V�M��l����W*��,[�.Q��V��s����#����8��6"�+'V��ga�"I�<w���H/�cI'P%���ܮו"x �g˩�$}{���K=�+K�v�j'y޹\keJ~V�S�؟!|�S%[����{��1:-���6�_o1ҷ �y��%��<ʝow���#��;��)a�η����v�H�n]oM�i�S���8ux��uw]}�=��pW�˗R����\�\�#q�K��[�֣sZ�K�nUsjcQS�PJ+���E"o�۞�	%j.f��"�[��2��ew%�nਔ$�u	0$n�
!L�HE*h�]պ�{�k¦e��_���1l����5<�8���a d�F$��H�䨋I��+�H�0���E�ATݯ($d��D�����k̘��:=j]8$�d��CS3s?���mm�6ō�R/V�����PZ��){��s�c�<z�/�����3333��339�s������o�-���/�=;J��V��Qd�����~�_������������s�������ʾ�'����ٖZӺT}��q-UEEX[+�����+���>&K2r{;��>4ffff~3<ffg9͛=���^�**��ኢb�C�A�A��E��'�b�TN��"�}>>>?�3333?YY���s�ϯ����.��l�O-���(��f\�y	�ե+l뛊��64N�d�"[UZ3�(��M�Xz��&X�S�mQLs*�ԉݨ{oT�DTFtԬ��-ch-J*��E�x����"V��fe��՚��Ղ��YA�b*�s*r�2��J����E�ԙJ"#�Q;�Jq�`�b%j�2Rڠ�IVҶ��w���k)[R�����\�U�j&Z��2�K��*��p�+UU����7��c&D<RI�
��me��}�N��y���jh>��7,u_\���:�/Q��s���5�������x,�-����A��VG ��(�e��e�B��E�2��H�(����n}<�R~fL�c2d����"V����0_�)JM"i�RG_�}���͞�5�4fN
�?Y��xGz.�Ǽ�}�B�ܵ��av���������z���`W�`gr��>��on�v\�u�7����W��U��� �M��P|C$<V���� �����m�9����B�}���l�{=���	�����[�ᾆ ?��2o'U1��t_S�EN�Y�s�V�Wl�@�T�c2m�G���o��lOp�Q�hJ;��������v5��;�ݰh��xn?��j��������M$�pK�4?~���e��+vcц��"�/���4l{����gg�l��v!�����������M���,n�#;c�x��*�l���������~ќ+�`�����1�>(2��-�߷��*M��o��g�=� �k�����<%�y �9�H,�Vr]��ia�|�x���m�ײ)��q9+���;���ٵ)♨�δ6�F����*{c��Ւ	��i���1'F�óBU��t9���W=uH#}�.�3AxB���M��t�DA	����=�	����x�x� |Y1W��3�k���֑�z(>wz ��^�n/=ݑ�,�zr}��;>Ƭ݉I�z�'��nho�� vḱn'�2D��G�X��W�/�W�w��f̵��C}���.���ڶ����E;h����>�`�3:��}�m.b�225�o��ڦ_"��s<��.�=�7|�{�(���|�B[k<�U�{-��Ӣ�y[�J�ԫ��c��/�)k�4Tׯ-u��0:k�5��nvWz�z��q�Oߴ=  *V�����
�<�?��׻�n��\���!dI���l���n���_BU����컾�Ի,ۊ|y�yU�唼X�!��p�ά�oxTtI�/q��\u3�Y�C��s�;3ria���2��C-���6K��~�����.�q�u���w:fH�$�V2�6�cm՝�zǸ�g�xv�#��=8e+;H�����=��C�ّk����n|&S8���9��R��{j;���ut�{C*�j����'SB��
�V��Z�7$w�{��X�' � o&���:C�63���)`�<���|Y1X�,@@��{�����n�.x�ש6����-(�H����Z�L�,t�k���;���<=��']�zXy5��"�i���4���¤?e]g����h����Os��tz�rV�]�{�v�1�}�>7%��#��(�>�an���@*��ˮd�׸��+��ó�*s�^�<!Eff>�یx��萋�('���u�6Vʡ�k�n[����������I�u���={2�<՗�{���"xg;]�[O-Fz�KJ����ו]��6�S�_e�u6{��S{�v�T�����MU���������b*�O��s�ĐI@���F�nv����O��x�����)���<��N��C��X���tP �l8�^���xs���r����fo����^f�&6����W�����yy�I
;����?Ot��{��?K����ժ�E��y�%n�:��y��磇�������e��B<�c����~��:;E�� �Bv����JJ_*�wu!;�yY��W@뜾1w �d�D{"��7�*y[�36�ͣ�I�g�,H�Q�2�KKN��z�x�$�o(�Cn�����Ӥ��$)p��t5�({4�u���c�fc��i�i$�v=�l�ɞܫ�j�)�"�ج�F ��_�d1.��H��v���4jx��UJ��O�}>�>��*���̓��t�)5��n�m�S�y�;+0�U���"��w�u��y���A���"�ص��*}"w�	��ʠ��^���	�v]�B<�;fk�&�ۚ����q�H�ߣ�O��+�
�� �쳌m��r:���o�66Jz�;�>�Ϋ��z����;\Ӵ�9�8|����a�ｱI:*�x��������89����G���>��H�����X��}�W�ߑ���R�Z#]m�������_OYg|k�*�s�v$�2���0^�$�P{ν��)�/Uz�^���=���l�/;�ﯸ�kmu:��.𑞜#��?߃gt�G�v���gkcb�����1���;�
1`�2fTw��u泯:Y	l��:	�Z��:�e#p�P:UJT'���*�Bz�a��"D�'.�X6��,m[�����)��:���Cq��se���x��dZsVz:�uEe<�"�*�,� ȉ��!L&�$Ё"�e��H(aE��g9sm�]7.�mwts��DgQ��2�,B��QNuF�>����~��iIQI���E�ez{^�Vo���g��羞��/�_-���={0?�&w�N;��������JT�/t')�ocb����B��y�̯u�!>�Τ⦎�Rg��f�zǢ C�^o7cs��7ٳ�cכU���>����ɽ�KϿO���_������=��rW�_�� ĵ<�77~θ��e�o[}�ս�tq>b���� q�}��D�8�|m�X	�����^}���]�Ȱ+m��[]�o\�9L��eYݾG��?��^ߧ�p3�ڲ��!��J �=7�-G;@��
�,t`��nH�A�����=4\u}�kӑ���{��k�A�Hp�.\�Y�Ы��&��e3
q�n�F�fW�_���/߇g��#�|��D^�foO��/65^�vm�b�Z��mcn���gln)�l���
�I/����>��BR�eV4�#����SI�+u.r�o{�	+?u�ϰN�F�߳�:��$
wI���4.�b]L�2J%l��R���D��Ku����'|N9ɮ�D�����#^�a���'�9Te����!�Ų��]j���˚�����&WeuO/v>'޲���kj�$t�;�]I������XF7��u�������*�e�]uJ��vr�zcS׷�<�⽼�!�y��ǝ:(Q$����W�5׽�u�p?cs��PG�;RS�m���RP��|��.F�dNb �!tnE߸�_k9�+@��R&�W��[�Ρ�3eCw��(wN���+����,�E ��-������˃+I���oT�6'���*��$�M�~�?g���m�)�%� �`��Wh7�q�L�Zq�9�{�ծ��q`���U�}�g�rS!�חR��aE�n�n�}�ݫ}M3��A�˸�(����>ެ��[�N��{kѮb����-������|��1�kWzv�Å<�m�nɛݘݪx�'p�I�t��d˭Δ��k/{�@�����~�}wm��Q��ӽ��;D�N:��=h��5��^U�ni�Hv�Y��:�j_-�,����A+�}<(��N|� �r�N�:خ|-ƚo�P��n�wl��E�Ҳ�l��ε�}�-��N��L'�?zx�x���d�1bȖ ���ѽ���z�C+T��͎�ʼ��>����k���͛|�Ͼ�ׯ�gR� D`�d f�^����bh�w���VS��fgĽ��^?��e���rzZ��v��9B�[�-�L_����.�%g�'鸥��gl�Lf�5��|�)fnFy���a~G|��l��=��ar�Jo/(�h-�o���ȴ0�E'���)˔	d� a�s:dWuk��T��`c����1�O�����|���5(jj����+ɦmqE�$}��)�f�"k����˶��eaMV�P�\�z���$��8��Qr�ck{k���9�w�vɼ�~�ԩ���P���n/z[&�Zi�Ix�nBw�k&�B�=Y��Ǽ5��KT
q�}��[�pD��{�����"���5&Eb�y}���zo��~c>��s9ME��[��??Ϋ�&�דnRM�8�uFb��u�.��.���tO�ʗ-�9���BI�����s�͚��\ß?�PE�W�3���aD��ܫ�v�����mfK|__��3Ji�o�Y�����2�ϲ�<1f,@o�ɈbŀW��]���M�ݕ2G�C��N�.;#++��S���dS.�TA��E�
�Ws׮�g�,e��R@�n��k��rI'p`�nM�{��x淫����ݬ�d��P�� :��p�W��N��^n�9����{L�!e盛*}�WX��|��h,K�����o�űۺ�[ٻ��te=Ϣ�]a�܋Xv��֫s/y7�:m�/Ҽ��4��^; ^(��=��fC�r���U��z�(�y�.������2�a�-age?�Ɠ����+���P�����Νv�ǘ�l9'jݍȜ��!�gT�z��LL)����ުh��zY�S\o[I��4��!��s{.��ڵ��}���31�W���Ȣ�v�!�yq�%A	7;��9�/"�� i�y�/�E��ϰ�fj�|{q��n�~#d��Rp�r�鈿ZhY���3)w��w��~Ǐ�nA��:�#F��;Ý����$٩ގ���,��V�Ǚt�u�5�q{�Γ�&H�ߕU+f6����Q����}��} >b�Ej��";/I��;[�����K�`v�ҳ{1��Wu��w�B_j�W@�B�õN�ylI����«���⋠YEF���D�F�r��QM���uك�FF21�̐�
�v�����g��o��谘`��o�z��EAǤ��c��0��'f ��x�����z�7����𼍀/Ɯ��	�ka�!S{�h�u�=;ިO�V�6��sJ��C+-�M䩆�X�=8c�{.���	��VZ��YM<
��h��K�/;�o�2�tƈ٪����j �ǯm�;��{4Db���zz]ǚ����]z*�Ш�-���sކ3��蚚Wu�p:�z<&-�B ��OL��n��u��;�)8���$�f���C�N��k>�i*$�nʎ�^��{�v�[Ykk�$�5����#���@X5���X��mu-#�N�-,���p�nыC�
5i���:����&/ܧ?����=�("��3?n�[�	�釶��Bl+;[ه�M�oT�j}޸�c��Ζ*_с�\cn�j�	�p�R��I4G�fJǜ�.uԭb$�<����^��U�A��,"�j��� ;nl�9t���Ya:-�ɗ��U)�f�Sw2�ǽ-��T4%y �î������b�X��;�z+w�{��@罷צ�>߽��2@�l존}^F�0�˛~�<vdl �"Ny�G<9�Ť@�c�����x�q2OE$��y�=y�U2Ѯ=�F���{� ��M4uEY�e��c��ja��oy�x�=qqOٻ���;�u�N�!ё�q�}y��%&kv�u^_Ot�ܟG�!F�=|�(�q�n׆joKݽg��w;��:���=�}n�/� ee9�PU�t�g�d���ꕕ}��ߜ����a�cA��65�YU��f�|�`z�3��{���5}C��7W2�'��y����}3뗣�;���*��P��f�G�Nu:FҿE�EVU,���{�͍�񋅋���:-�m�ߘ�6�_~��w.���-�/K�����[Jcx��-3&-�Y��?e9]�gg�Wݟ�[�k�W3�uT9����nR��9����v�Gr��Y���yS&!j=��y`��Qw�G�Q����}':5�f�3{���d�2L�wWU�"�h�YHGR��,ԋ=lJ1mc�x·*����]�]���~9E1��63��>�x�z��Vዧm�ؗU��{4;������(����3	����]�#c&���!�m�s�������V�>���ʮ�:��c����e=�������Y�B�N�U�6�篜�H��V��^�-��ܖ�u�
jd����SL�mX�Щ$귾�r+��֊��6yX1K��EF7�S��c3Rç�D���O72�1��l˲�:�i�ï��y[X�ƛ�_`v,5�&.��¾P�
�p�lgL,����*�-���&嵵;GӍ�UA�P���s��L�*����a�����]��
�ݥ1ua��1��������eÚ�zv��{ډ藵M�8q���cV���"��#�Ǜf�ڮ�1V���m�[��ę���}���_c�Ws���a1p�p9^��=Նr�PTb�	uQ�i�g��7\���52����������%�����iL(�����	8AUlW��%B�@�;���|%u�0����<���s�#�>GC+;kM�$m�d�����j�6���`���*�g=  $N;YK;�KT���A��i�p�i�g|isM�I�P�<#�D^j��~��oP#/������fct�l�ޱ`�������g��2��y|�x��E�/�f��F,{��v���� �o.^uÍ��;�n���l� �gs�]�Y�f��@�j��u!}jJ�|�Y��!:�ۓu��WK���ڨ�6���ݴj��Ky�U��[��>c
t�ds1jc�U����#�ڬ����f=:or�HR��H��g����N��G���ΙE�}����e�`��W*�)�����l�:#d��5s���.���!��6SCX�yN���g7�/
�8l���cn�Q=��jZ콹X�R���݊��t��S�)w;��}�x됰,G$��<��l�î�W_gj�����f��wbR���°m9�v�˾e��]K{c��O�FRv��b��_ޝL�Ou�f1Wݸ�iܽk��q�}ڏ��o':͏G_��M�r�x�e{�Rr������on���6��ٱw�紎w5�����=�}����3�=^\�9���*V��q�X���U��x�ݱ`�b��el�V��?Y�ό�љ���������9�g���j���س���Q:�ޔ�U�#�VDL.a-��E����dٳ����||h������Vffs�͛=�R6�,�+E��LGq�sK��ĮP�ڥj)Mte�Nښ��+��K,���{;�O�ƌ�����effg9�sN��wh�d���T���!��6���ҫ�¾@�em�QjTf����le�=��g����������333��9�C���b�Xwg2UqE�A�0Q��R��h��WiS-I\N9�TUj��R��d�q�W�m������h�J����+�ؘ��Z�F4�m�=�X���(�[h�fK�0R�j��X���1W[;���u�"�C*ٍE��,���O-0F
�.NҎ���qUX�ֵ��H�b;�d�U��1ʹL]��(*�h��r�JU8�QU]�Y|p��#Z[Y�)���
I� �@)"�f�i�q�U��X�����׏Z��^����y3JS��=WU��UQ��k�޹.%)2gށ���e���*H*�i��wߛ�?��������ކٙ޴��d�8�
���0�{��Br}vk��no8�1������ug�GF�Vt���j.Ц���mD����U�m�����:���ѤL��RC^MnU-��m�}~��m5�+p���3"��^�ٱ#ʴ�3��:��g��M��w��f۱Z�:��~����ݺ�����y��;8^�0�rZC<s���_K���r�-������_�=~�Oz�T�#��vM^��z��������>UzGC������-�&�b^������l;���ژb�(��X��~D������Lʥ�����|s�{"���7ޖ��ۜ�ٍZoɎf-S;�N�t*�l���EF��m{��)��S����Vl\C8VN$A>��\Rꩬ�C<H~��ݞ�\���S��ZXX�_���'��r_֟�5�Ty�P6x����LWZ��q={r�]ћז؄pL��Ǖ19Rb۰Т=u:�.��Z�f�[��T����K�~Q��;D��z���� �ِd�K�Y�ݩ�K��=<||����"X�`	��ѝ����{+�X�^pI'y G\V�H��=y1��묧��]wN{sTk�O��l51���r��Y��=�O�ۓ���lw���axrvJ+j�%J J%/#������諧�����|��w:4 0�^ܽ���7w�vI&�W�[�ܽC��3��{�9Y]���藕t*�tu��&�mN5�r�wC&���S�<ם��@~˓�Q�/��k�s��~p��nr/���@�y�gn�з��%�(*��dWY�������t�M�Vz�F�_�$�7�ß��]���ܺ|��#��:��k\\�S'}iuHȞ�Eێ���|c�_�[�^����M�^��ogG&��N��;i��i:�d�^�i�dW��8^��z�ۅ����Ά۷ܫ��O���5Rׂ��]�7�[w4��]n�,�����ng@����D���Տ�&�8�X�/�L/�O��2��V�8pD�(�Fh��<��"�^��V����+6�dM���8�(�SJ�0�]K.�H��L:�oe�w�t��N;��pF��:=-"��J�i"]�=H���uE�t�m4"73/V��#61�chCs������}������o[�m!��y{���@;z�7��1�[#3�f�U&�9�FO�d@L����� k� ���H$��Q��6+�U�Y�'a�P��P�^�����o�y0 cL!*B��-v �ŷ�䪆��},��>��~��ݒ<�L:�{޺tI�-�kgo��4ճmF���k���*�ʮ�����O�Y�Ӽ��36N@�q������g#6w�DeDﮤ^�����W�퉢�y1w�v�~c6s�o��es]w��㚵<S��'��^
����v��P�e��$N�������:6��^���E�(^�M��έ�Y�Dkls��{6slV��|�.ͻ�g��0,V�cØWUys�:��r*��*�(���~�� ~��Y�ot	�g����x��ҳ��3��闰76R{���Fd��@� ��Րֲ��}t�jB&��$�}C<����9K�n4�^_�m=����eKe�W:�jm�����l�{�3��-`������/�&R;o�v�(f���IF����X�L�b��F1�����}�m��o��w[~�`3��fU�~�;�����ƽ�������v#��!���ߨM
����Cm�;������l�� �,���Q}4A��sSr�M}P����}�8􌌗�͍���6�2ZZ���Սة�����8��rjv���Y�;����fX�^�:�p��z��U�ɺ�Fz�f��dff�z��}S�;��!���G��߸�����|�z�a�y�U��mu{���b��J7��[x�����}�z����o}}S���Yt�8������ݜ��*8�qZ�_Ee��hd5e4�Я�f9­���Ş]�&'[�{��o���ť7eG���B�\I)�;x%�=������s�z_=Y���e,�k����m[�롸s�oX���Y�O�-�`<X��D��N.�\yuoc���j@Bc������Ս�������,�eesu�(\��]Ny���4z����prcS"��oeǩ��z�V�\-ͭFww�Y��&~I:��"Ǵ�*�|7��g����|�F^�d���8
̵�u��g/D�ރݧ|��9��_�� �1����{��=x���|_K#R�,�>�	#�<7͚�����k�ڬ����.v��{g����=�SӤz=3��mk�k���n�Q���}p�����~W.�H��SgI���^�~�����+��+(7u��3�Y{h��΍�f�Oy,�#�������z}|+��i�^�o�O`~GnJ!�<�w͚Ң�2�pgD�Smz���9�%�ꝺ��eW�>���� {wC�gVX=��ι���b�D��5u��Θi��o��v���z}wq�����5�&,T\��ִ^�o�dM[��u�L;_���B%����3��~���	�"���V/�[���9M��j���j���]o�<�s�Y������ɡq�cQ�b�n1Q��kܚ$��9�w<ov�����SVp��ͺ�nzl�n-���5'���7��Q��f���j&��h�B`?@'n��e�DÙ��.�MK�\������idD�LO!�8���xgF�߳��՞�j�HE0�垕���>z��:���qu�7V��9G�Vb�����@,X�f?��ܘQ����N�eW�C��׍C�����鿞�����Lnm�ݼ#���v�.��[0=��am-�rpeOf�F�\Ez�z���{���R�-0�A���`���-9�hqӓ�[t�o��<�#�
��r��Ť�{\g	��˹B�l`�2�>����{���"���%����OJ��R����W7+r�^�>�<�p�;�Y�L���������XW�/�^d(������	�$��r�4t��l��g�'���D(�A����[2��ׂm�y���W��}�v��F�E0>��k����q�E^���Y�p}�y���+|�i����͍���]>�5ۻ�fs��/8z�xa����j�܌[;��i�\k�|��o�\��v�
���T�+�nl�� =SFf��n\c���G^ƽ����B�4 ������tL��7��o�g Z|Y������.�pX��ْ�N�g���aC��-Kڬ	�j�f�f�;���S~�&����qf�_ìs�<��i2��{}�����I8V_q7gfզվ{qP�:�I��[��R'�8X%$8�E��n����i�F'% T�{X�X�,X���Ԋ4�?G{'���\YTQU4�ƛH�1ve8~b_u�i��H:=�;�9~����,�C9�FEe�t�ϧw�3]��v��=����`m�D���n6���7m�^U�|����7}��4���8�dy���W;����8:�Z' N����~÷#�����:s�|�E�0׷�]�3��B��@|��>�۳�%�������L�-��9m��oU�t�dd���_�T��{>��t���`L�˝�e������ɺ)��6>�@�cm@�,�o|�b6
>�,������{Z��A�v kq�z���u�/9��c�r{��lI���O9m�/^T���g�^;����|:��h	���^�!�u�e_�,C��4�)�܌����b�7�g���F�4�<9:���v�����O�����7���c�F׮�-��J��)��J�lnr����������AL�̌���G�X6Ok������\�q	�J���� D�O���aWf���6K�w���͈Χ�K���V������wS���D#�sb�{�k7�f�G�ZǙ��6� LX,|�1»�{��>�UN�W�W��vqcoF���`X�W!�qq�(���S���}\�k�\����`��u��V�j �tU��^�9����Z.w��u�v�y�_x����;L�w͋�~� �ȇ����{{"nm��ݎ����9��$���ҹ{��{�Q\o�f+���n����-��my&&LL�)��֙�S�c��^{��n?�<�M�����g�q��:=�}������!�����G{߳O׻�S���$�;їy]Y�Y}�������%���H�͸/�Zsw'���օ{�n=}�ՔI|I$���t�h���؛���!�b�޺�[��{����K�/q��.w���w^Uڡ��-��	F�T޽[niؿm�D�����x�@���4=y]�}�sQ�^z��Ћ��y��i!dڏ_��mh�n�[�ݖ�c>��>��5�v�5����=�+8�8���7�1��Y������K�x35������[��C���	�^>>#��1`X���s'�m��G�m��Jc���t.n�z�')&��������NB� Q/Wcsٹ�W�@�X�y����%�e�ƺ�z~�\�ɯù�����r��}T:q"i���//nn	#(e	nB��������f�n�H��CN�h޸�
~��f���Y�4�Z3����yk%���Xz�,7ƿ~T��M���뾯.��6B|��S���1�w�V���M��|��3YS@s�9�����i��^�����=��^va��h��/��0`�i�kd)Gz�@ƨ�q��X"o�K�[���6X����+"��r�{k�8�p�`�Z����X&&��V�ї�ӼW�f��n���֓��rR&��;k�����4LTV��S�6N���'�������ђ/��̴4�=Ӑ2��幃��8���T���+/�M[م?�����ܫ�2mwf������0s���X��pG��j�S>fŵ�2I#F�o[�wI`����3GyM�i��i��8���+�e�܃���Ԩyz����ŋ,@f��ޝ��=����xu��@�g{�͝�-��7�ǣ35�pA���嗭�}�~ol� ?S�a��aK�{8���c㙉�A���<z�s$�˱ 'O�w)q����پ�U���@�|e�ێ��v���=�0Dרz:Vb}��v�&o=|���]���ջ-*��ȩQ�l׽�^�Ǐ]�n����α�>��E�@�<�#p��q!6�1���M<t��y���O�t�9	�L�kkh~q��9my>�ܤ37#hEs�X���_e,�Ю�G�������{[ӪE߮��_da���,{�Z&鏵�y���v�9��C�>�z�;�ܺ��p�.�ve����������j�7
��K�e�:"H2�d���i5ڎ�X�;v@��6�ڟ+H*�-3T�����_�� G�!$��� "B���9R�ȴ�f���S	!!C������H�NP%H��J�j�beZ��$�,���ūV	*����-Z�H�b�J��	V�T�c�1�X� �VX�U�j���%J�lQ%�$�bI,UZ�*ʶ*"ū*�JE�V�BȨJ�lT�K�"U,Z�D�U)"ȩ��)"�BA�200 ��	,��T��a<Ij�J�Vő%�`�jرȤK"1� ! �c �d �@��B0��HA��#�@����#FBF@� !�B0��H�� B$ �d�# �!@B0��B$ 2 �d��@��"@� B$�#D�!D�� !@B0��d���# ��$"@� ! �d�ȢK"�K"�K"�O~�� FHD! B0��@��"HD !@BF� !B0��@��#$"BF��Z�#	"� ! �a���#@d �I�#F� ! �I�"��$"� B$ �B�"� !@B�@B0 �I��"HD! �I�� !@B0��H F� !@B0!@B!�#F@�@B A��@cB 6�%$ �� D� ���$��EB��JHA$! � Hpd�%I� a d�B@��! )$ #! #! -�JI  D!#�a �@�@� D!#�2H!��R2@B1�HA� D !� )[$�ĉ  D$P�D$��� ������$D� !FH�I2$����@"@���!)�A"E�D�F	�E"H�D�E"HK@�"!��$"�e��b�U�e[$J�e�H�eYb��eYT��RX�?����+'������ЂJ��H�D���d���O>?����W��@P��W���o�_���?��߁���w�G�?�q�C ���R�����I$���U!$�e����%�d���?��O���?�!$������O����Sϒ������_���Oޒy�2Y?��-���D$D��JH�$XId�@H$aF���B�$�J�,J�,$�$�dIB�J,$�T�R��Q%�"QQ%D�D�(��b%����`�`$��	 D$��$H#@� �[$�lYd�l�"BZI%�O�JD<��$�A$V� ,!0��a ,#0�Ē"@2 �0��0 � 	2 H�$A�� 2 ��"@A�	�@I�0��,I,�Q%Q%"RIQ,�(J�(KJ�J%�%RIQH�%��O��K����r�HKBH�l�$��$@$!�<���������!��??����@�O�y'��_��߯��?��J��O�����i���"H�d��O�������`I jBI��z��ro�X�H{��=����@��Y'���������0(P��/����3��h`��H����?������	$���2[$��o��}�I�;�O��$�$����d�����@�����$$�?�I�O���jC����_$�O��O�����?��I>&�~��o�BI�O�-��f��'�I�Rt����Od�����|?�$@��b?���W�O���������?П��PVI��cWZ)AU�6` �������F����N�Mi�!�]��H��
bd�UBӶ�ڡ.���*�ؚլ�KV��i��UJ�@�]rUEJ�%J�n�R֧fD�UG]Ɯ��wk��ں��v3��kv��vWL����up�ݮ���l���Y�r�u��wn�m�����n�[uV��W5v�sk7W[n*�mҝ�д��v��ۛtG7C�ee�������n]5+js���k]]6�h$WXv�swn����r�w+Vv�[������껺Vwn�k:�FΫ�ru�u۷wu�w]ݰ�37wq��ɭ��d�gn�[m�l�t���ܛ��;�   oo}Z��F�xv��kc%j�k1\�͖���<�{�7z��i�l[Y�n����Y��֪�U�ji��\�ʛm�Z�5��-�����5���̨��]gs�s�m��n�;6�
���l�   w��!B�
(P����|>�(P�E�Ow+�3m�s�:�ٛjڶ����i�kT����KcZڶ竻�mY%��<۶��Z[l���m6j�kmݶ;�f������eV���7]������]�w�  '��iBKg��(R��[�z�*ڝ�@*�Tׯy�	A�Y]T��U��Ȫ��7z碣�D��z��V�Z�������a�w;�ͻ��jU77VwNݻ�  }��(U_}���T��=�8�U"�R2�QU#��(��F�*���"�]�ʪ��ۺ��1ESݛ��*�7=5�wf��w�t�"��]ݻv���  gS�7���{^9�B��=��EQ+sǼ�i{f�U
��k�w[f���y�"������@�Q��R{ʈ��w\�正�5L�6  �>���4����y� ���l(P��r�@�������  ��  ��� P���o� {�sY��6�5�`�]m�渻���� ��z>�k���jP u��  �w��
 
�8 )A�LP��ۀ��  �@ n����� ^����kvtv�w'v�uL�v�v��Z�  ���  �S������m����׻�4(3�8 �=��y�  �޷<��6�g ���{p ��{�����]k����6��w\w�   |  
�� ��y碀��� �=�x� �x` ������ ���J -�v�JMdcu��i����m�l��9�՗;mҵ�����   ����� ��p� PN� ��q����  u�x��{��  z�oH����
 �7�{�(
���fJ��  "�ф���  )��b�JQ驓0B)� ��@ 4 �{SɊ��F@ I�&*�� 43S�����?���{���<���O�*��M�vʃVh�~�T4w��-X�?�_W�}�cm�y��Clcm�6 ��cm�m��������1�@6�c��������̴��<woq鬺M���V0�%,��Y�a��x���˘7`P=n�{s�A:T��+��X�/M���i9L5A�vH�u�ya����{�����鈬��\m�?N�kC���=�|C LN��p�<�ء��y��o"�$Ӣ�
t�T���.��z�;�b&���{讯�F rU��ļF�L*k�Z��3s� X�ܭ%&Z̋@���z�FcӴN��sX�)�J�B�bp!J���]1sL��p�0% �Kb�t�У�w�[��2�.���M�ʤ�F���,C�y�u��.d����R��f �a�<- �Q�B�&�U�c�l>���v�Q_n��Z�Õw0@s4���lˉҖ�H��&0��U�ofS7w�Si��)�hMtr���B�}�:�� F�T�Ǉd�S�YI�(:B`ϮK:\�tu������A׋�@*;IU��vr�ЧR�o~&��)��^ȁ"Nc�뉆^��7y}"�!|@����lL����A[!�[�ok5�l!�������v5�@5�+n��ǗopU��H+���-$$"��`�3 �i��mڽ:��������"3! l #�I�'�D��&�2,vm�=4X�f�N��ئ��,SV�˨��R8�&ڛ�Ӧ,J��1n�e'�ci�$�۴�^����YN���<.6v�2�zJwOl�����6�Z��ih�u-��w���w[zemeu)�!��&��6��T�m\ݔ`�!�N�*'�b7g�F���ꌵ��n����*豢U2�4u���ދSuiF���qe��6��Z���-� ��U
3*�]�Y��Y���L�II7�O��!|¸�鐣f�''C�mE�\S��Y:l���%V�I�"��G*�W/bV^�@hkD��V�	��!b?^Ac��i�c`�4ZI�Z�+c�5:n�b��@sp��s�$���ժ���x3���'0K��E�gт��a�!�p�//6˕F��z�m�H���S�Ĵ�lm��8��H���U�J�M��VrS�%C��,�.)��%��@��9��4�f�e�f��Z��9[(ĖczF8����0B)���;�c�X�MEf�Ӣ�:C�Aմ�l��(�V(� �de$�^�5�Q�x2؃n����GS.�%��V�y���S>|:���a${'#x���1a����N�d�`��5���:��z�Z��I�֌���E:?&�n�v�۔��m2��(��3��"�� ��{CT�����"=Ѳ8jЭ4(��ݼ	@p�$�E�����]d�F�
b����j��m<_J*ȅ�1�~;�j[!�C���b��G��]0%�q-�I��{ Į��5�t��6���l:�u"�;��GL�2�\y�:I4��z.�����M�9��q��F�S���l��"9���[�ehVe�|�� �P�{�Xд� @���Ţ2�9�c$�LQ��k-%�&��Yէ�wmР��"y�
Ն�1�V�cE����9F�U�<x��FZ �˨+,*[��G0���V��鑑)��̖ohS��KpC41ڻ�Y�R�T.��Q^%pdHI��'4*ںY��L�S���(PD�b�@8��"!6�\fO8J���<%����PD@<v�q�'BX�]��k{g�d�-��j�˩t)�Ҕ7�n�^�9�WJY���׫`-�`��<�sD��J�jVU���ڋ�
�׵��EP� �U.�I�c�V�p�kJ'vƊ� ��������7a�'D3�H7]�&��+N�H�S�A���öZU�H����M�q��9!��ik���Kn�VL� b�w���!�`�QD�Fc%82+۳$�A�sVDR:�P��	[��q#�E��2e�S�*SRcͫ���4�ST��U�u�[�zTXTO% �*Fk#���n��u�a�"������en��z Dc�A̹1������3)�L�H���iXj�.e��CLu��9!�Q[�p��5�j�[Đz!1n�0Ȉ[��(��X���,�B'q���a��˼����m����������dѠ)��M�����v��� �Cˣ��x2��'n���H�h��!62����xN��XɌx6�~��p'9���ٹ$X�.]T(�Up��Nʔ6�o4��M�b��
�Ǌ�-;�>9��r�oa���$te;�֞$��wo���[1/L=�d͸֚+Z�Ayd��چ^7�c��wQ[r��o/����`/
���+N���7!�>��-hv��x`��Ttk�	]಴����nZ�����L#Z���x1����������	�F&`X#¼�k��	`M9y7f�alZ�ۋe�CT�%�I
`�{��N���X�8�d�W��%_Ш�8��=dm(j�(Zb�D�b��W���wzs����*Z4��wvf�J�)\���U�RdwX��Pt�7km�V]�H�:�^��,m�go%�j��YB�n�3"�f=:3W�m�kCn�Yn�!Hj�6*:��ʟ[81Ę"�+ݬ��*�%�m䉱1���FK�u�4���Z�I�h��|"�E<� �֘G�;��}2��̀f����O�;b��Mځ���;4Y�����E!��m�M,0�S�%�0�u�ܧ���.�u*ˋf�S-[�yX�L�-P�U�x@ �������,�a >����=�t�م
b
�Z��zIۉ�]k���v���v��o-ּ5��B㭆}�vro.�+KB��!ױk�N�b�7���{Q�Ҋ"���љ%�8U`e٠&�	���T��x�J"�0d0A��]�gHȪ�W����g�I[IS�M*���o)��BS��)n�����ƪ*���Y�cJ�\�6�@M�!�Q���{p�Y�b3$�H)� ��D�ϔ��v\J���|#rc3)�"��ȶ��w�g�%�AWYLs���d�J�$�ipi@9Z% j���@ˇ)mK�J2ރ�d���7l�u5y`�� �mk� ��yw�MsY|$���N�5��!�e�����l⽕���VV�+�z^���e'�#���b�7h�L����Y3A���8�b!��`��ס�[4�2Ε�,8����Ϧ[�,��8.�e9i�ƚP�Rb�[�^ S�ER=/0���֯��#�ᐿP}�qǣ=�"Ko����0~�SKt�Z4$�I��#�&d�F�Y{��#�x��l��U�"V]�gV��`
��.:O&�*�
�*�`��X�Ч��F�0����w0HD���lź�8�fa]�$��K�x��N�V]�!j
��9��EU-V��k.�+q��"u�IV!�����m��Q�PƐf� ��]��=��'C����H�ܬ�2�6������ݹ�1cpL P��X9K5���4��s!�Z��m�����	�[�Z���G��W�+
�چ`��D?�c)�jN�>�X0����[j��&4�0N��5��;�aùT�K���3�haL!5����D�,����h暶E�M�U�S��j�4�Q�G0+VN��#�!>1�+u+�mشԻ�7���Re.���"*&�U�kn��m��'jҧB��aDp��ot��a�_.�1��r��A��5ÆA+t]F,�@��K4��f��P�8�{����\��nMݓC�)�r'���&�}�2-b�dU���w(83��[x��`C 8JD:��чmk��:�8x>1��4R��NK.E[gO�t)V��2h	M�M�fA$yEVVAJ[���S��m��qb�Q�0jy��T�t�E��b��ߣ�=vo$�tT �0�,����۰�BjnG-m�,f����jb�;*�(�mT_8cC�l����m��!y�lrV��x@Wmin@5n�h�*jw0��!�[yVc�>pl�
YD�Z�[�-(��e����o�swD��}�Kݢ�I�N�����`V#3v�F$A.�dU��z0CTv�6����-S]k>��lSךۭV����^Pw
\s{�q
,��YJ[�̊=�Y&Ѐ��6�MwD�ME�<�6X���!z�������z̼P�;V�!m�ԳF���U�CAzT#[4�\�m�B��"S�f�:�@�pVQ%R `���Z�y/1l���� 0Ѐ�(Y%�Q����r�a� �jwK�e�#������W���ڶA���if�d����[�t�V��L�n�V;R#*]]@���X�ڕ)H���-��Z�<�YCq�61X�)T�Rk2D0+g w�(⥛6ւ��6\����_���t͞�熙����{1����O�Lh�)'�m&͔lQ���k���$� ���������ki�z��0آ@�MV�,�:��+ T�n��*]�̌�kF�n���@�����ZS+VPp�(í�ɋM���\�C�j��q+���X�+�\���6#&�tX�7���š�̠X�!��-�e�uʈ,a��&2Hq�~��D�� -��E��,J(�����B6-�#�#���{#�w{� +H<ppd(�� t��&�E^�Rj�լ>�Mf��`e�Y���2o&3ݧK2�CJ�Q��	��5c;Y+�l#	{+L���)��F=b��Yؘ��Y�E���K�Z��S��e�i��ul%����30�N��h;o2�ȷL������%�Xsn�Y�1���˚��F#Z�^
�7i,��m3h��f�l*�����ԒFe8�Z�/n�e�^����KP@� �(���&p�gr��fϣ7Z���x3�2��E]
���h��,U���m�sv-,�R��[����*�gn%��U�+w�R����E"���Ӈ$��;v�)�e@�ҡ8rj{C�Ю፛��C6�];�[*cQ^�*�h:j�Ep$���#6�MM+t�-n:oDp؆i���K,:¨V*���p9�
B*�kSb�a[c��7A�V�u��*�U�T�����˙�U�+c4�2��"
�T���^��ɎZ7�(6�I]�n�'�S)^�-��#E�Ґ����t�����AJ�a8)�NL�.�p�u��,��l�唲c�%��ˎ4kt��Q����M���A�^'Lٓ&DH-e� ĵV	hІf�$[&�9��%�񓎰��YS�0�����<�2Oa�R�eX��2�����
mY� o(�Y���ifWFh�(�o*��G�2(�A=Srn�e�X`p̋f��6�7t��ɋ2��X�Y�nU1�n��
����X�L�ߵ�_M9���K��K!Z刮�Q8Rm�8�di&�i�AeB�y37Vk�zf�:R�1f���c3YMX��� n2��b�{cjZ�EMu��F�7lGIn�,,ښ�߁��/-��a]^S�pQFb��SѹU�BME����kz�%)"�f�#��WP��1jw�1�ּ��:a=z
�v]��1��(��<IǇpG���L��ʵ6�ft�[��:�N���
���z�[xn=�]��6h͑�VE��aXi��@I2՗{F�rg�t�n>K
��b�Ξ��Òh�XW%(�҅�ۖNj�����q!�~�QM�m�b�*�V�Kɬ���/2�Q�V!V�:���5� �M�E���1��a٘2�f�� ��bHf�6ސL�Y�d�5�fZ�U��体
ri�V�8X�r���-0��Oo&[��v�(K�J0@����*��-�e���fŕq�V��0�յvĦp��Q�X
'���Q�LcŰ��B�^��i!˳��&K��v�ܤY��m����̨1�r�������VEDK�F^a:�ilGB��W�����:�4�]�AV\t�`�,�ɏӆ�	���lH�,d�M�_�ǣ2vr�����G�0�pv�8uݬݷ��u�ܔ��r`Ne��lR1QZ�WR�
���#�S�U��D�̧n�P<�2��LQ:�q�Pԥޚt���U�C��V�8(U��5ݭ�pe�:iA*̏iCB�ܱ.mL�	1ͽr�:�+\W��XTj\��CR����˫*����?h2�!���03shmj+L�?E=�=�n�i����ѨL�2X&U���b��U�hnVz��P̟�r=�[�W���^X�UcJ���&~l}�o9ѷ�M]��IB�0co*�зS�\�b
�aҭPñ�a/f���E������x܋$������:)(�ÍU��v"�*��k�$d�)@ �IŤASQ��r�<װ��D�B$56�d���u�`��6��6M��Z��S�p�^d�3#�*��6�[�I�b���!:�r��7[t���L����JPA*E�$�:o7&�[b|2a���qDq�8��á���A���F\0�?&�;Ռ壺fӘ���pD0�z+f26��[��6� {���:X.��(���oX�L�^�K�c1��ΟO��aGZ�7X�^����WMR�XC`cJ�&�����2s�f���sӄ���^Zz�fn.���R��'KUf�bc�� \��_=anP rҤU�w�E�ܓv[���7 EA6�?<fv���j�V�x��腌;�f͂��� �԰h�7�P쿕ӫט��XڕL�nC{ET���3��ճE�e�1�G������P/!�ua�Ė�7i��4[ҭ���<��Y@#�.�i��d>9#���H��`c�V�������7��z�a?{-�����k��t0��j�G�s���R��Oԍ�mlŻ&U�)`���'����9��=��2St�ךBKT��nQ WQ�ߊN�-B8�V���ު�(n��\��&��)�f�v���:���
º+���֏_:{�Z@�*r�\mVus�o���f�e樺�`��)'{o��^en����:�h�B p�������I���9d�֪�&B%X\�f%bOr�w7��%�d�j�$[���c[�of0R�F-t��\�=qY���u���9v
T0�$G��TA.s���Xn�b�(�'#�ׇ%*����$)��_#��]S�H��]n��!u��=,�sGmzБd'r� �#�8�����W�x���R����¶�Nbj������7w�r��<ן�GY���
�u�*��A�qh�����хON��Y\yܝ�����[��ݨ��V��X�޸9@A�~+N0|����<����H죑�;Quo(���+}SW3Yՠ�䴧-$�@[�.vz�M/�Ј��&��̍oq;��G����I�v�6�t��*v^i�Wv����۫����x�z��g�]�*�r����G<	��EQ�B��.��I�����s���*{���z�Z���%i;co���WhY�{��7)����#�f��.T��E�W�Y�N�̯t���������zp
�|����RW�撗G��t �	/g��Ȕ�%�"Ͳ6tR!�<��
� 9bV-[]������ΰfv;e�q,�Imr >�\km�GS�:iX��g!�Ȝ�]Պ)P�;d�2N
����]\�]z��W�u�H"�%p�>��S�w�G ���o�,s�@~��rΛ�2!ۜ����O�Q�̫��IK��2���h�s*@o �#`��R3��dq<�S����;��[QS�[L��w�m��,�ykY-�L1�=z	�������y��Kun����g@Wf�<������n�5��+[|������9���!��_� D�(n�zz�,�gj�mUՇW�Y�V��ST��>}�RtV�]��v���M�F����,��	�0��@��G�)�7��l��Z�?��@n����#b:�].�y\�g���<�2L���	�V^��˺�w�zv���2�(+.��1rh�^�(F�y�6i��Q����f�nL�+C�
�z�ӳe�,b�}�*z�ͯb�{΀�=sq�.#t���z�ȝ�q�!5���/�#@M �9����	�i�1�8v�|�^��4��0a����]�n�M�xS�=�Z�Hl���l��8V���z���\�*~=�^�"�Zjtw�� �*���(�t+��>ʧ[b�e�!�d�;iy��+OU28�?5�1A��0�΍4�=ŗ�údzY%y�
�|%5�|%}��C{69�l�Z�8�1��#P�o����Tw\�hѮ�;_gwd�n/W��A��8��^�>��>��jL���s�(����"��X5��.D<��~���䤠ޚ��;�!)�����j�|@c)�x��O˶�8on=4}��wX�t
�s��1�՚=r�
u{f,Z�GQ�Y�9��`���=]�/�;�Fd�G�7�ŎX��]���r^]�cl�g5"��3�S[�w�f+�\��ڇs���m`Ǜ^	�r

96��M\'Z�Y#y���X�� 1�g(ۇO�C���ؽ��}���+�|��,inԦ����E���1׍�s��cv)�r>�lf<5(X`֡�q/��L�{Z��r�(�B�q��7$)��)�[�{�Y��zՓ:x��{!�h����d�'@���b��o��5F�;P�B�\�~*-8r!��@�gG;�^?�F�X-]h��j@k�S���$�`����d�t�.���
eq�@���s=ſ`|�j�w5�Q��m�#�z�n>UO!w���c�7��}ϔ뜗�̔V��mL�X"P�Ⱍ+=���3�
C~*>Q�/��6U4cxڀ�Su�(���7<w��eT�
�Ǥ�y&M({��Pl&
T��<&�e[��hql�!�����|p�w)Ʀy���f���7Eӣ;��)#��Zz�=��:,o�W��2�E��:l��Q��D7���uז�"���M��ƒzo����|�wf�=N����]��IrgQ��j�R�S��Q���q� wA��իYB��[ʙu���I��+�Kٌ�;�QT�eg4 ����و�p�|u�*�-��]v��7��Xa˫��)˷��yԚ��'vB �ΰ����[6����5��|
����Rv�eX�t��/����|�[L����%�QۆV���t�z=�Z�(S7��Q�V�o�\2���S-�̃��GPB�E�3.f�CD�=~����u����m(�~3;i�ҝʯ!r�xBOe��}N\C���o�4Kw`NU�кcqWn��\������/SXL[N���W]�x��nT�p�lK���s����?1x����|8R���k�h�x���S��E<�e˨��D�t^݄
H�ר6�Y���3�N[�=�z'��b�Jq@4D)�2���|�o-=�^!�e1XG��um�J��@�Q����l?tyj2&�&�⫮"�Տ�;�+�3�zY��vۺBףp�D���0�ǧn���fޞ�;_{wuD������
����1�dn7��:7����������A��m�����<��/&X���/��I'2�ڪZ>�{4K�xN�ճd<�����3U��ń�(/��m�Hcau�{�F�	��B���߶r޺��ʒ�]h8�)���jgsҩ�|mHt���jk�u!�e��R��d
��m��DT�t�V��:�j�h�5:�
ס7�մ�ܭ��ĕ����c:(���-Kͦ��W��q*�'U��K]u�.�^�E����7��/:�j��a��6v�����wv�9؉�݄�z8k��6+�5ى�OE����Z0�K��7�����Rx�$|��Q�\�"����:���z�%�Q�8�� s�����U����gfd3Oy��n;Q����K�Lk_������r�z��/n����a�/
S��sx����\�Y���E�[Oq�W�����hM�<y2��v����%#�懈q�,�9�c����f�wI�b�ͥ�"��h�@We3�0��,:FopH�:S%���Թ��>��;��qs��{L}�_X��vG�Am�^�XMy���ޖ����ǈ���b9z/
}���e����Ʈp�M];���R���`�+t	R��o��������B��GDT�e�c|���C����s��_?V�ќ����-��Zb��иb�����0X�XO�k��%m�@��λ���Ў]���k�:d=hs���򃆹y��6�e�{(ٹwJ��ŋ�E��ف*9ʭ_4oVLv���ώ;�)bC��!cH}��<V�
svO*�Pw;,h�;)(�۹�2p��*b�˦����F�Ǔ�Z��1�����i �
����9[ַq���İ�7@0E:�6F=�ᩛuZ[��.�byC����*�?wFU<�t�X]�p�%�w�U���ڀ.J<wR���S
��Sˢ�����X�U%���p�����d�������|�}��?p�~���d��q�]�}lD�g[ܥǲR��d�A��oR��I�<�K���V�ӏ(ʈ�v��/3���U:�J��B�an�,����f uՖj[G� L2M�^�B5�
t���[�)rgC6����.�B�)�
L�^�%�t��C���2�Z�Ub���]=5b*G%��35����Ч�H���ֹnQ�L��R@����2�%�{l�.����h�E�HI��z����O���P�.�ܣC)�g�=c���_L�Q�_b�]��Gٸ�hF�a���g���zW7b�tJFBBq�3箆����6V�ɔ
9��U�G]��+;]x��:g5t���E��ş]@��ڐ>,��](N��t���b��f�l�7��bw-��y� ڜ��a�Z���q"ʦ.v8����Pb�R��t��\�9�W�N�+y��{{�C�C���=J=�O���0w{��f�!Ya�Fwq���L�V���-t�b���sb���Z���4��\ZӦ����L�)�b!{��q�6�e �N<���{��qG��)�L�L���r�y�NN9v՚�w	[G9͏����ӳ[]tD�E0���^J�,��7a�n�/�З��<��JW��_$�������R��rAx�!?�_nx��q� }v	�˟k���.���8^����R�{7bm6��7���zYvgE�����v�s�͝X��ykl�t�5p�x�3����>�vՏ]N��lf��h�*�����'������t��a�z������G2�1����ݢ]盇{�{�Mࠩe�����]W�${�x%�ʝ��ze-�{M�$I��S�C�'(ۨ@�"��s]V4��oA)Vu��V��vNͣ�҃Iv�7�Wu������me�������FE7S��s�{��;�۰y�2ÄĲ��7+A\C�.�5Ƿ$���3Yp�A)@V���Ѥ�$�AK�poTCE�xz2b�Y
(K�v�XZ;2��9��n�
R�[���Z����b-%����l�R��Nʴ�.OM]4%	bL��x��<0�_g0&_����_6����p4�I���0��Q�9V((�}tj7�~�Y�ǀ~I�"�ց�nL	����W9<��r�w�k���oxr�ݣMkNF� 廅�W޶��%�k�ţ* �»a�&Kᗻ��	�s���6��C�Я�c�	�K��f�W�k.��ok��c>����:���I9���|��!�����[Y��@c��)�R�V���&X������o4�(�Y�+��{��xZsӯkv8vx�:�L܌H�xk����l�(Ӹ��aV�H;:���k�[����z��/Q�;
�NL��h����(���TA��ia1�Is��;P)�W�[�f��7�x�C�[#��`͞�x��aީ0�����d�%d��Ȑv
U�V��W(՛Y�>���]
����\�B��SB��4i����ذ�6Y��I�o���C����E�������M.��as�F�r�
9��XM��	V�1�ހ�
��D�U3Rj��e
�^l�9Aq�(��c}����-:��/��q뛯8L�X~|��W�A��4MԼ��&�	]B~ɽC�E/x�}[|�n�����&4i q3Y[�NM�Rp^�)�&˅�A*`'����}���٦�&��X�=��E;V�v��K;��	��3�/!�jRxŨ̞,��d܊ZJm��r��hٷe*�IV5�
8�ب KI �]7��i5k ���b�գ�+���#��nݎ��6��վSigv͚h}W4V�b�Vɰ����=�G� �xج2H�=��	0v���F��ˊ�ɗ�7��Z�w/u�7�XۉÐ�6�8.�8�8<="
�����pY��CK�­-�t�F�S���|k��;p��\�E+r�.�o�uf}s�T7�]������\$"@����١u�ţ[�w�n��IC�u�y�/e4�iJ=�Nxw��N�m���l��I���#��V@�Ҵ�!�8^l�����*��55���iP���,��.�p&7sa��E@W�}�[.y��q�_p����'��u���������nų½��Y�Xs0j�Ty�d�V����'�Q����˳�g�����p�p��G�ktK[�O�$�5pg``c�۝uOgwn��pQ�h<�-�p3�ո�C ���V�DK+"���w)=��%�o�����>����О*wj�e��F�:�������A����Y/^�E�蠝(M8��h����Ki���j�F�F���5H��l���_Sr���iʃ�}�i}����w�ن00B��BdK{+Â���ԅ�b����J��Z�����d�t q[��5��:�sa���vZ��D�]@������ť�a�鼲�y�l$��*������,ILKqe�"�u{��v��B��S 7���WQ��F��n�3�0p�*�W�z��Rꕻ�
8�́��+�N��{�|v1�V
�S����7�ǗN�QU��\a�J�f��9%�5>P�\��L��	�e��I<��N���( ��Gl�w�ޞ�6B�uh�°��{M�\\��޹;��[sO"ܧ��ű�?\'	<�(��_��d���떬�bY�A-e�p���`[�����}���7q�O���Q_%t�mx��9!c�g
Uͻ��Rݺ��w����NK<&[�]�'V�[}Bgc�zq���VK�5Xtr}�׺���gr�#���8�4/:l��I�r�U�˽Z�U�4�jo�^��f��ho���z�+G��RX���h��=���`W���}sލ4;g?e���(Iҧ�|r?<>������'����+C�/��{�T\���)ZZ�KP�>	 ^��*	�Q��U^�}��n�E�U7g*����.�2a�v������=��Zx̸c�Y����TO٩��DG�}��G����>���|?��K R�2�� m��zv�9�0e�Һ��r>Z�[rh���][��f��h��6��m#xy�#����|���{,5������su��J��c����>�ѤL<��v�[��6�K}0M�����j�;;)}�;.�^��
� ���[��0U{�<�����4n7��jص��#���,��ba^�潞�2ꃹ�su
���o�L=$�y͇�1��^��� �3Wv��:�f�f��b�R'��|����E��7��S��8�m��@���T����}�9�cֻ��!�����p,�b_���<���Z�R�V@�s��r&���yB� n�	�\�)�w�Gx�]|�;2��7�#h'�m:�t�j����>CT�� �{�p	�����ťnf>:!�9�Q\m���Q�^�6��K�9X��a6�Y�(�^[޸�+��WZ���=IL��F�Z�>E[�.T4��(�;�U�ry�Vv,>�%_v*�T�T�u�x�I�'����"��GnZI�4脽�3�z�{ٱo
��<�^�n����¢�Oe�'/tr�@&p�d�i
���2b���͊�@�W*C���-wg�w�a���S�:8nx��3�^��,�w����HJ��0��/��5�(�ꇴ.�1�I��s�l��{R����h�o7�����	�k&�hf��ǣ�72�i3Y�X1�--�
�
V���ź��?!m��l����z|8�4-�U�E��: 9OT��F�69�qv\��.��Ł�WW����vB�(<G��1���8�m×f��M���Q+{Wsr�7ح�jt�>�+n�4��zVb݅K6��1ҭ�C���*����^��B�o7�rU����IR
��N*<#�HC��D^���܋�./s�݂���(KzCyS'�> �IY������͌�|P�)�:�*�(�������"9�;fK��}+�SHq�������Ծ�)�ث� ��Reɲ���#�R�i+�z��z�8IEsS6��x����w��U�=Yt�E*/5������R��;p_l�G���*W�]>3�ը��A_'F$@�Î�g)���h�LsfU�u|j�#��:���O8jА�l�\�i\l3
���v�>/�����R�A������Ý����{��n���4�+��>��ثy�5�A"սS�}��Q,pxol���Z͡�5��������^l� �n�4v")[�J�w�SY��A=y�j���o8��)�zG�6��,���X��J�o�!%Ǆ9\~î���\�| �nt֡$V��tS������e�Q�d!d��$YH�y�K���e�z��؄�~B"����P�i�ͅ����{Jt�L�Z0S�u�i�zu��Wr��������[В/,_	�J�X8Ĉ� ��h���#��9a�僦a�?s����qP����2�	k<2ٌ��y>�8���qd�8L����J+�6�}qs_��T"���׻{�ho���Dm���8��'r��h��$�����%x���U�h�F_]�p:�镯wf�2�@�u��{��y��������`ⳕ��.���3��I#��>��Vu��X�>Ά#S��i�ѣ��;Z�+|5* �!,��]�֛�7Q+�j1�� C��,Jd�O�����1�8���s��(��[J�xf�ۡ9Gz�⧆���H��� o9�d��۫�Q�2�G�zNTM�^����iov��Iw��n�>��y@����^��y4x����Ji����^Q��x��6楁ꖪm+\iw�"��h�}F�&���um��9
�v�=''�>�L�E�[g$� �0�3Q[x��]pӑ�ھ)[<e��#�4,<�D(Df��.[�D�7��J]�����x�p�����&N���{���-f�m�凃�,q�N�|�\��6c��=�i��Kk�S�=��,��s��Z	��a�fg`��o�n��[1�˻nIW��!]=�Wޡ�l�9h�O+��5���&�lc�V��y�� �����2� ����&,��1���i�K:%�d�[�t�eF��`sυcY�[��+{�o���ᚶ�l�� �;��'0�o�Y���`��-
%�Q�)�O��э^x=f���Ò�4��2 ��7r��1��Qڣ�@�啡���ֱ��_�K^��*���6�X}+Wf��	Kr"�2�ۻnKj��u
�IW��s@ۛ��SW*�H[7�����i\��2W�z6|�+��`��yT�]���7��mFg��h��R��z5f����עW�՚"��S��ܯ�>%�vJ�F�_jG�{[Q�g�%%ة܀��-

����P�� ��%�%>[wy���-.sm,�a�k0A�xr錱a݋�ʕW`�-�mvB��sV.#�Mcj[�y�PQ��k�M��>�.��kUښ�}"�u��NW�,Biɱ���a�.�)�=�BN|�!�/��"e�L�E���M��H�e�<}Զ��S#�������8��ޗ(�<�֖-��;F�]*`wN�n�����
�\��^��@rry��N���e��1����Aך�O���p<����ڍ
F��um�f���%a=��P������KDS�Y|��O6w;G�;�[�%��-KLJ��i�g>���f�D2����[g�1����L�"�X.,t��j�!��l>�g$k�=u� _sw�*
6ү+-���/����gzZ.�3�1��}���;UX��� |t����ss�ھY%�kx���`m�R�uѕ	�ν�Λ˄ij�r�����������jD�Տ� ����6gnod�1uU���r�e&�sfY�Ellj��j�/���V)�K���3U�#6j�u	3���������:T��ݪ��FJ���3��6�T�|}�&Şُ��g�(w���	%�;;�AO4�p �65J'vJ��SEb�;2�7���v�!��W��xٺ�T�kl�u�.��]��ج؆!�fQ��7홹�ԡ6S�gP5�z�,�ή��s)_n��HiP7X�V���J�E�"�:e°���#z!E���c1�YB�a�a����)��m�=�`�׈2�8Eq�.���R�2��w*I�����v�	*���0Q�y��*1>C��]���»>WA:����3�VZVPs���+N�:���U8U�jԠy�iZ�n�>�q��
^|t�7�&vk�Y��I^^w<����"�ɒ/g�4w}[�wq�^U�'9u�(�v��P����u��79���mq���"��1]B�=��@9��n�4蝔s���v��G��y��7.�T=��x�b�d<|7.m���e�v �"`7/���@���81�֕��|��u�oHk���yN�ξaWC�jޫM���Tyw*,i �)�Ճl���Һ��=����<�	>�o'�\�ٛ%<�g�X�u��n�sym��h*�u���`�UaM��9�Q^w����1���|!b�kHf�'K��2�_p�-֫��V�9��XQ��6->)�n�]�d,�<��C�]���u0�_�KӉ�i�J!}��9�h�{ܮ/l&i�	ʜ�+[��:E��$���3�r���]�ĨW��+F�n��VRi6{kz��&3$U!��G����T%,��LD�8\���]ڪ>W#�t����Q  �{+�ꆼ���37���*�܊yl�Etȱ!}�&=|�.�^�2� �Ƽת�v���͍:�h*�.�N�(�ǩ+ ��93����~���)��q���ú��ś��<�����4���G�H��Yv�˺3J��-���`��'���Y��>�.6K�ug��U��L��[��[
MS�k���Ж3u6���� Ӥ��Ҡ����s�k8_Ev\�8���(����-��<Ӹ��G,�`ث-�V�v|����Tj��v�NX��ξ
�U�"�&>S)x���ɧן�3s�(0�+�٠_����V���i��sD�[1R�4�3��/��A�S�,�u|lQ��2�Z<��yB�s�h�#{�n{cq=��fpO�c�s�{�~ɖ���N���>#�Vq�^3�����ìh������{u�4\Wr���q�vҲ�W��M^���)�#�ד.��YY���E,a][]$�K����^����fmzf����x���P�=������4����z5�[-TB��-�Zج=����pX~H��LY{&u۩l�v���b�W:��盜w_��J�{/����SV3��5��с@��!;U.p,��W��wLKc�!7�rpϊ���|�oA�[�u��ٷB�Y�(H���z�jq�/�W]-��Gtjv�<n����m���S���,��k�9�B\n���r����o�N}��uٻ����L壣*VC��'q�*�q�$D��%�3�ʻȰ��'�ϻ���5lwpM0ظR���q�mV����/��&����:�.�j��##n��^�=84����U+�ڴ�xj �~n>C�C�&����E���_{��^�I�Q�{4�]��R��sJ��f�O`���S_��_��f��;�p�}���p��A��v�{`GP�ʟ�Kޙ}�,��$�ۛ�p���t�O~mr�^�:�%��e��`��k�HNn���.�����b���^%6A�,eQ*B��$AD�n�>�-�Ƿ��]�o�l���[{��)�4�Nq4Y5�^�BA����Ӗ'��<�2\_j	ǩ�ŸCot�b<�c P��_,�<E'��͏9ڽ�Y�?\hǀ��Z������egW�-�0#�.�D�u��*y���}iҺ�c�G�(�Ҩ��/�5iF Tg-x�7u��&H�'9�!��Z�M6���-��}C�@3�<��)��dܞ>s"�87.��Ĩ�u�꾆5����!Kd�f�����AJ���Pd���<�;;E��ۜt�%1�n���*�P��a����g����*]D�9 �(�к��|��*��Y�\����g�1��i�ڣۊ���c_R.�)�ռ���e�=r����ym��;Qp�)���qRGz��>����vs�+����A��w9��郥9�;�{J���l�<c&í�K��z��dX�eE�r���c��Z�c�J�2��:yx��ՃwkG-��~.��V���$re�7P���8nC�U�����(jg5��7nb�ڟt�SvJ5ս9��pIy��k��:QYK%���s:���hu�mMc�|`�.�N^�\E۬:�]ml��?�,Α��uzr��銗R���.`Vk�o�ݣ��J��t^�x<�3'j�����3h!y`�vd56��~�#O�V�,���3��E P��{�[�P�z��V���{�,�� *�h� ߧvm�q�q�i�d�T��\�mi�RGS�AN�!���H�����Mn�Uq����h�k����꿈�HV�=�8��,�������=�+�x��r����=c�h�����iQ��7/�C�w�P�O2��,fK�WN�i^�9���tX*���3�jWv����\�`���,��x�=�]��{��x���:c�� 3�]x��%!��gw`�>���|�]�r*����&*��q�~����=�D�{]h�,�&�1�x\�Q}F�83�fJ]n�4����)Q�!�,W'Q�<���Bxt\� R��^���ض�L�����!�(iA3/Y��, ve�eҪ��{<m|�/9�>�Mʎ�V3ْ���BE�`��S�ub��b u�c�l[�ں��u���M�kA��:_��7F��z�v��@�-�:"�cZk���-]	S%5-B
�u}Luk�;r[���
ԛ�P�հ�:h��
����ՃY1�Ŝ҉=6	�Vmgr� ;!sz�v1��7x� Ҩ���	�}�!\:��.�T��Mz�;Ӷ|7:;���rSZ�Q�k 4pY��j��`�sr�59���Q�Xr����
�+�WÆM(�{u �7-N�B��*���s��9�t��=ȁ�N�4]V�CHl�5�L��v�4���sS̊�*�tKHw�Vm�4��ͪ�+M�R�4��5/��E|o	ķ�X� ��*��g�����f������jR���C�s���UH�%(����Nro��
Y{#���V�����eh9��.����;�o�(�t>�]�'�j��..�"D��(��-pj��<�jX<�D�#U]���t幨Պ���t��n�-R�n<��uy%J�(p���� ,ëA݇3E� �E> �;�;4�r����^��[�f�Ň�`ÀwVqT�&�ŵ�L�@�rӘ�.���l<$����A5,fӴ����x�'ue5ղ��H�gX]�VM�}�`�7n�h���ߵ0����u�n�#��1i�4�Ӵ�T������B��0-�=O ���7�l3�ԠȡLPtH"V?��$^I�:�Ws"�@����sY��j�z���Kv�ںэ@Ѡ�S�8uns��bz I��Cp���x����狷�B�@0=��=X�1���sՑ�0i�����{7w�x9��B��}W�.�+��WX�m㱨�`$����dܼ�>�U-uN�䬥����щ])�k�(��2���|0���|3l
�+(��d�_�tٷ�a5�U[��2��?�������>�����~���~���N#���<u}.�kv��#Y���o�D Y���5Q�?et�G�6C�n����Kq���$.�,��/ZnN�ݦ �y�Q(nn��td�!pO��u��%�����x�֭�9׭�b�����`� ��9�;2C����y��r��k���q����-y*V5��;S����h�1�Qx��h�M�΋u�6��h	`�%�ŜX4��N���u�sut㝢�T3��КtNB��}�����Ś�;twP~��Y��d��H�2~[m����f�{v��:������혃�|��&U��>��|;'{4<���]�*Ǆ�hӐ�cumD۰��jU���s!oE��=;!��FN���&ȡ̝����P����j�5�t�#S������������s�4��h$��~;P�1�Q�m��8�q��4�� w����� ��BC���Y��]��v���A��s��H�!3V)i)Q��P	����Pm�����k����V��3�)Nj�݇�˩$O��=�3u[@w6��'�# �m��m{sν��5c: ��z�Y�w�V��y�>(�N�Y�'�P=����O?� ��|cz}O�����%�m�C�u�"Өl�+�qSDʲ�q�Y|���՚�'��}���h>�H���-_��Kێ�SY�#
�RГT��"�4��)*�SS��k"<fJt	��.���j��[���9˃��W�
�;QQ����N�H�QNư��#�
�zʎDDQw&%W21*T#+���9À�UUXTDQ��hE�(�IQ���U.U�$�W��'Qȋ�&�������U�I�8˖t5��TQF�TE�2"��FN��"�QȎ@Qr�YUG9�30��h���Q
*.TQ�<�9$�T�5f�f�)+�\�&Ur����*�H3P��\�N$��"�,�#�\(v��U�K�	��u�PI%AAg�$���qĎ2�t�E:�(+���N�G*�ӕ��eʊ�\�ԅAP�dS�aW(���r���I0�3�Q�I�#*��L.p�R�8ZF�*���qⓧ*%1e�Ll�^8�kEN4OR^A*�.�@�tDeQJ��:sCYEV�DVtL"��YI(�p��Q/[��J��U��2Q#D�&a������?���^�|A�N`�ܝ0��5i`�20,���]mM�o�ْD<-᜶�}���8��z�:j�</���]	�����}��f���V���;Ā�>{$�*��W�.���nՈ:� �w��U�]Xd�$�/j [�ɺ��H����O���˴�$s�D��
7��s���j[�kp�s+1��t��r\�
u^, ��G�eR�<~t�7=�uv�ɭ1�O��W�@�%�˒��x�-3l�_*�T4��4j�w��t@=�@1�=�)%^>J�=\Oz�Y��7�Oj�#�M}�9JዄA�*\�M�=*�� ���Z� 4^"F�w�����}3s�۝P{�� 0Y��
/�:�Nc�|�D�Q���֧��3V�=��o�57�׽�%��N��:���.�py�o��@��<ga�p=�^�V�f{�7|���q�wc��v����8o�T�[��m����b.�P���y+�p�z�[����Q�T=�3gͪ��Q��r��9��=��tᰰ����u:�z��)��j��o��}�Ѕ��Hf��n���tF:��C�5�ˡ��v��y����ݭzS�R�-������D]{e4[	�������me�L���sG���/ww����M��`�^M^M��7�����oAU�Н�j��:���#�e��.=����	`Kӧ��B7� V�y�9�*wvvX���gZ�`c���W�pi���ob�]w����]��ӌݱ_�=6�\�E���ʆ#\L������}~{{{�)M�+l"62��M��|ˮ :��ʳ�4��Ǹ��__a��;ʽhF8��O7�n�Y�=������]��%c�J�U�_�E��*��Ѭ�M�:��G���k8�[��`��yKS���{EcHmE�.
��T�����5X�@�K-W������W��" ��I�jd��ǵ�ֳD��e��*/��>(r/܇�	U��p�V��W������
��	W�����d��:��P�L�̌��_6�C�0@ Y2��0��b�>�i����Q��r���y����u��?n��Z]# }�r�: z+�oȁ)u*��G[;]���Ȼ��~��go������$]P�zi��n����E&B�������@���h���ϖ�~!x�3z�M�y`�U.�vk'c�_+5\<f(8O���R�[d�a;��yC�)����?g������:��i���)^�S���@�+	��*S�Q�����'���X�(9~}��;�V?w��u4h!3r�@#K�P]�?}�ܻ����'���ˑ�VI���&z)�9��3��ǃ�tu\�.��X�z�
Q1jHT4�����pH��<^�؜��1fͬyx�<L^�N�N�h�aB�]J<��9:p�c��@{�(ߡ�J�0\@��>j*�x�㺣�z���β+*���.�g<�z��ȟ�Uu���Q��_w�]��
�	\�����7�Qc:�*�h�o׭�̋B�\>�t5pw��u�3j�-�\��5�q���G��dJa�~`�p��Bg1hZ���C�T�oҶU�"=�X�"�}(75v����A�6�����rV�Nv{�V�>��V[�%{�!>�u�]V�ao���|w�׮�I��'�NL�;~��JήROG*��0�J檻'����0�v��'D1�V]0���Pc=*��(83�=��o��~��2eN�Q������ߩ�!W�p�*I����ǣl�r=�7;9��gէEhs��:p�>�Ht���4�4�oՋ�������^���'�).8t���rm9�MJ�#A�Tۣ nٔ=A_G�t�z�Y��Y����\������9��+�c"g�
\���B�wq)˻_zVw4/q.^,nW���orչ��S�L�v�{ܢ�*	]��J�PZ�#�4�%�˳����]}�T��O�Rv�Q�0�m�N���!��z!,�4`�r���0�p��S��1{��&_U�AȖ!��nmb\`�owm�׫.[�GpHI�2��$��ݧw�["�mS�G�<&|k¼6��x����W�����E^��^�Kq���n��r��dA5�x����E�B�:�"P� ����0��G��W���j�gвX��3�DW�HS���Y�u��ؑxj�j����p�����^�(au�����Ʃl�+!mA�����dt�D�঍�n2P�J�ޝ�=�Wy��w�.o"��_���$e�9�#���[ܢf)����������}���48d�)ֵ^A�Py�x�7T���	Z����yߝ�)��2��F�tvV#G=�.�ͩ�^d�}�X64����t����z�_ 3�߮��Dt�U���9�����m��׹�A����X���<"z7lʴ@����Ǯ1�J���_�o�%�IR��<K.~�9bp?�pf��66v�_ԫ��S�\�!SK�8�bZ)�g�LX�ۦ2U� ]?C�^���+�p�B�vd�}�hVϯ̇ҹ:��t�zt�}j��(������R��C\�te�]um!����w���ٶ�E��N�r��Y�z<0�	ӐŻ���3�w��z<Ӡ����|w�;�DK)O\�F%�5=��y��W*�D�$OS:�m���/n"���iN�$[�+t\Zط�y�a����c\V7½U�d��oi��¯����Y�n@׹�Lz�0;����]x+��X���mnk�]�t�ږ��\�[~Ϝ���t�}�LxL��o����ٶU�b{����a3!�+WNpm�v�1F����9�"s�^A^���5k�߶�\EBe��q;��皊
�P�7�Χ��+��1�sV ���5��2�C~�b,N%Pנ�Ĵ]F��Ux���Z�-� z�!�"7�x�3'�^\ҵ�
�i+����Ul�8�P��l\�|އj�D��ǀ
���^�l	�_p�����uwq"��i�j�Ef�I�yF�q�7{GH?=�}���w�����~F-C��D��R��~�Xp`����A<}mw��+s3Ч�j6�|v`9��+�L?@~�(*�� ���&�P�M���j������>%X��G�Y�w/��AZ}��^~�;�Kс�x��Qf�Y)�����SҰCjL��𩯰�4Ә�e�����|��(k(�ܯ0\���������U��9�摙-�����T��3��u�v}�{Jj�z�n��P[�=L8��~Y����]��c�A�O�����sצY�Z]��n�^�����b��},rۜJ��OY��r��*�ek�����鸑=٬Vʂ���{G:�����; ��c�{��1^���pyվ Vi}{�~7Ԩt\$�;�D�`1����
�xm�L|���������n�������]}g�yM�y����
�J�����3��@q��b�|ew��	U�ƴ���G	^J�X��H��\�*�A^1�C)����t�����P��g6lPZ���ݚ���}x�\_>|(�7`)|XY=g+g����b�SC�1�la�*�B�<G}(k�ZW���L!p�U)��y���Q�/�#M=��nF��$�m��bpt�;�����>ʵ��$[���ַ<��W������Zz����4O�vM���_dUگ���-�\+�gvo�GC1�
������gK��r�Ew�k������B�؏LF�7�h��iZ�ݘ�z����I2���Mp�J����6�����[�~�?{pY��g}C�(���"+��ޏ@���f�1�;�i���OG�����l`��?�U��O�N��J�\ ?[�����ʖxԪ����wv�+Z~)gJ}Wj���`Eú_�8��v����$��l��h�_�[��#�Z�1� +�M��V9��v978�ɶ��S���	WxkY��"_Q�vK܁�F�x����y����u�F�^�L_.,R��mѓL]���^�;Ʋ��\_��*7����	}@�y��ʡ?o��z�C��0v�`����u/���iq>"Ưj�����z�@+n�	,x<<-֦O�F��N�a�F �=����:}��ɞ:�|��n�X"C]�TIګ�`������Z��}�	���N��ڴ����T�*��7_V��d�CG.e׸�,��WAv{ī\ ���|5ǹ˜k�N���<��\`J���!"�ʠ����6̥�~k/n�t1<xX�^C���۪�(�l�{yVq``��_"�1P�銸���ؑ���|F���+;^ZX������v�ҷ�zO[nTbЯSE�>5yS8�2��u�1����~{��R��{V��w�p�>�k�����_23��P ���e^����2�1��}:o^���_U�
{����#h�KQN�Ss��Օ��Բ}6Kױ�%v7H8�����E!�Ą(S��^�j��Y�CΜzu$s�ϫ��u���+��앯렫Ӯ+�3-.��������N�s�ȹ_SA�����s��e���q	�EΫl�U�=�����*�hȵ�K���l�=/aP�w�����Ĭ�6�E���h�e���ظ��bW�}�+��s}��5��J��2��g8��uh��s�z\�b�*{ccTT�g����H[�� ��μ�<�*rφ����yN?�cF�w.�����9�^K��SZ��غ�U�%f��C�+����{�n����1�x�L1�~�g�lz%eA�@JtN���x��1�n��|�����a�9�}�G���!^@zg�I��=�UԽ=��<�����φ5�8:͗���y��T��N��v���tn�~Eh�tf�����!S�����!%B�����NQ	�~�f��>�KdVȰ��PO��𻿂�c���m=2�/rR����Xʟ-��8�wٍJ؀}{��T-cڥr��ەKa��wm"��^�+h(c���t}JX�Hz��	�<�x� f� %�Ĉ��9ۃ&�,9^2���R�K+�;� ���=ۊ�(���,�	6}��h]��z�[�\��Q·J�&8z�Շ}����Y�o�Y�J��{�{���Y���P���۠g���U~o»�1��A��Wr���Z����N�-�|��{��xvh��0(e�Ľ��\�R���	��>4���!ׅ�ǰ��'��9p�5"B�5|3n�.l�%	y2h8u�W#[ql��^f�����8U	��U�L�z��c1�Q;�W4���w�1B�ߓT@v���gm����$��:�it���v��C�kE���Eo���"e���~���R��)��H qE�w;������_f[���N?W�q`�����ÈR؝�h���7���o� WY#�vy�������#��b�7��y[\�n���^��ޮC]���g���hC^��er��W$1��7�p���u���퀐���U�D=-I���b��x_�=�������I����W�z�EnW*Չ)m���;��Oi�|�=�9]�S���KnO���Om���jT�@E
GX�݁���o�C�RW���`�cCQs�v�b�U�vb�:[>Zc;^�5<%�����@�Ԧ�n��%���X ި��k{�	�ߟ��^�������f�6V22j.iLC��J�u�bO�"����Y���}x��s�.�]�O��p�0���1�`��͖�g����B����T/`[�?WQ�J6w%B�Uz{�œcE݅\)_���O-d͎�ogb���]�lz�,���\ �z2.�ߣ ��o��<o�#5.ktC�$�ih�*yL�<i��A�����__|ng�������%�o1���6O��lQ��
�啤�4������G�d�`Y�OΗ:��聃r�/^T�I����1�?nL6��u���@�7��u0zu��Fb����c���"�U��s���p\�7�toՄ
���>���K���^, W����{�'��B���y�(vw����zj��(�����F�P�T+��N���L?D��
�$H�%��{mH\���|s3\S�r:7�̤���]o��	5�z�uwpŢA�XYfܗ.��7D�qU��y����%!V �z�d�e��	�l�
9��Z�����`)��?Q��&���I�G̣����`�sZ�y�	ۃ�9��7����]�f _�> V��Of���F�?_�w�(���{3���o�Z��ѳ=�,�d��j�<�W�S������>�mKGn���5��Ϟ�;�m���T"�)�O�1�N��eHB�d�xN��d[ڮ|�j���{�B��D�����\>lƽ7�B�,P1+Q"԰�@[�1yQӛ~d>3��jgQ.�	*�}��}���� �g<��n7�īJ�zdw��ϭ�v�+��ڤE;����w�*d��s�����WH<��܋�w{��Հ�xϭ.�S�>�_*�^�w�}_xG��VJ�W%%~�Tt�E֦X���Ygx��A�V�╈�)�0��=y�%#I��b���٦�F�4�wU�Ymh�:�m��k,A���2c�91if:��vt.Ȳ+��;��9���ٕ��D]��wC�����)�2I�ڲѧ�:�fթ:�r#��{�
�Уծv۷Ie����,J�ιЁ��*�]�[&S�`�[݂<E��)���uW'r��m<����Fu��=�J�¨iٍ#M�t���\�wd�M����/��J��2T[��r{�r�����sD"+����3t���s�`jbd,E�m���)��p"�M��i�:�.VՎ~�,x7)wwz˜��&�ʯvޣ.�1
���Z��u ���|��%�a�m��{�묺k+{E�������{���3���xs� VhK:�&ikl�+�9W�ꖹL`���x�9�Z�͝ZT�Oj�n���
r�olԂV��%o8 ��dO�r`���n�(x���8n�lN4�6�����XS�<m��gvV�M\=v˝T��s��Q�d����,�'��J�;O��� {���FШu_
��BUɋ�	��[�5]���U�:�+B3�;�7���9��1aY�74������
���zuö[�,�޼*��>��I]�:u�/�xNnގ�A���W���eAv@���k?Jt���;n,뱡�7M�����clMĤ�gCf�Fv��A�Ld�ĽlwP�h`��dp#n�u��<�)c�-��s�8����7N͐;��}@hm�EB&�6��WÉw���Q+��YB��y�yq�ܔwq�{�N�m�u#�c������1�J�]Nu�"�P0�	e[��Y�nЯsJ3@��ŗ�/�O��_|��\��+#}��-�s��-�r~�cu�V"�@��~ۮ~k�en�N��U�����c9J	Hx����b3MRN���r�,�����`�N���Pf�וK����p�m�j��3;=����"b5��}o�������:����Z)��R�����vO�m���ݛ�Ьp]8�sZHS;����[ekI��x3���L�F�3Q��8
�v�ѽ����ٺ9HhP�.�2}ۢzqe��+�؃�G1�澀�����΅j�0c�ׁ�A�<I��ێ��k�@�E,�e
v�g�2.(R^�.�Qf���a��}QX����)�g��_ea�u�h��*\)��ꆔ6r��B�:�϶��l��,���'@�0V����;����YR��$w��s�q05�due3	�z5�F\�����	���IҶ]��rp�փ�e^��IT�k��)J�]Zt�66oZo�W�2�����݅L����i5��������6OZ�.�f6�\i�fZ�u�H@+�բێw[/ &�u5W}W/�[�/�_�v��*{�_c��g�\v� ���Wob�-��E{�̥���x��r��kP��"d�Ƶt�t�����k��$�;������ �K9�ʥ��9r"T(�k("�tʌА�Ial5 ��Rd�q DaHEʨ���+�b���A2*Q+2ɗh���m�f��AGE��I��a�9Q)̊̍B9��$b�&E+$$B"*�BB����J.	-E.S��A\�Q.ERKI"���F���*N�\赒Ir�+�^R9�"%eйs[@�KYQD�r��E��-��%]��NDL���d��W+�����B��"IY�+��*���AADp�!0�҈�	Q�)0�ͺʂ(�x��EUTT�"d��9���"���,�E\""�U\�Y�H��ES���*�˯U9"�"��#�IDQ�C�r�#��gr$��L��h��%i��AUDQȃ��iȊ��UE&E���,��&UUjDPT{bAyB.�BPJ�eL���A\�r��N2
h�$� ��ek�����I�8��Rn��zu��'�zN��OlO:���%}ٱ	^ydz��bYKvᶖnR��!@!�xA�J��G�@ E��͑7�븛�~����}���\= x����G�8}w��$������ě����R�c���8��|"Lp��!}�
g����]G���a���Q�AD1tN��G�Н����|pu������q���0��{�sI7׊��pU��}O�����'�{?�������I��A�v���u����a�I�:{�8�����o��g0�tT��#�1A���v�~'{BN?ɿoy�Iߝ�|=~��<M�'}�{���|OG�su	�����2��>������W�i�޹�^����^�|���'��1��ކ>��#�B�奄<w��$�L*��$��N���~�~N8��}��Ϳ'�ӧ~}����Nރ�y���i4���	4�O��O7��.:��~N"﾿����S9~� ��{]����}#�B:"Oh�7��~8��i�V�q���Cϖ�G��ߜy�;�m��:�_G9�����w��ͺ�@Y��������	'�����;�qI>}�~�|�@�0��Ǵ,9'{��|BD���èq�O�=��-����{��C�i�uۉ��H{M~�<��8�����s�q���>|��㏧�aw���I7׊��{������Ψ��ݵ�>���RN<#�DAǏ�篽:O=$��}��������x�~Ro���y!�=����}�� ���C�S���'����8���|�$�P����>���>�ymvGl��A�YS���~������u	'�ߏ��<w��
�z?w׆<W�?|���<�bz���:�?!��o���>t��]�7Ǐ?�zOi�aW>���M�	7�'��q�jbM��b$}�C��eh2��Yۙ�����C��n��������o�OS�=�8��Ǵ�y���<w�i��V��N�J�����Ou	����y�`��'�|�c����]���R���`�>���7��:�J��W(��_>w��� � @��P���O�1 H��o�x�$��G�w�~C��>]@����Ğ�����O�z9��q��N߾�C���=�s���@��{MRz��ͺ�Bw��7���y�/�b�&iǎ�̬�J���Z���}�֥;��t7X°Q��7ލi���\x��o
�8�ރ;�j�=��L�8�K6l6K�.���F��L�bK�G�:��n��}�q�|�L��=O���
�Y;�"�X�J>����N�I�R����EYj�b���9�z���V@�ꬿ��~G=�}|z�_��~v�I��+����L/����x�Y��u���~N�u'�^s����������0����n�������8�]�>8������~�*�
��Ώ���M>��9�;|C����n!����o}�y�>�?����m��}q�G�|w�w�������o�8|v��|&����&(�{��x�}C�b�����u7�$?Q��o�����\ސ=��;��y���qē���1�C�����ߐ�����u�I������ .��wO������&�>��FX�,g�����{��OUm������ߟ~x{��|q?o|����aw����v��8���8L"o����L/�������C����sώ��㷯wS���8���p�!��?^uo����>��E_�Sگ���x}}>��I���=���<@��ɯ1߿�1�o�N�s���~��>�}�N�}|z����}v�M��������w����=�8������.�{��Ou��ŗ��}O�>��F��L?`���>'�8�����$~O���|�u7�$���]����N��ÿy��o��8�O߶?� �q�$>���~�ͼw�� E�.����P�n���O$A�1�H�Ծ�!����Ճ���P���������z�~|M�>'��@�I7�$�����8���z��= u'o����~|M��}��v]�>�����Z3*}s�75UWܖ���#�4C{bq�oI��zzEw�i��ӿ'��w��S}B8��=������u�v��:�_[�x~v����?&�S}{��7����|���޽��=����U���h�DDH�؏�C~w�8���S�Rq�?�n���=$y}C��\x�w��8�Iɧ�{Oec�RC�rщ7�'��=�w�ノ�r>��8���oe���Ь��{�s*v�-Y� ���">����S���w��0��w�0�8���o_��I�a�o�|w���]�&��|ǷzC��8��Վ?\H/�?�ޙ��H��"&ы"�P�\���c��W��7�}=�{�Y���w�q�Ex�\�f�vܡ%�p�y�%��~!��y�j�~�T����L�:R�|Ena}G�
���v�t���[�X�*���xMy1��["�_�m*Y����n�7&T��M�b�re�CX3m���!�)!��Xy�3.�rju�H��~��)�ꈍ�@2a !����^�&�����9�30���*�7g�@9�W6�{~����}�\�a�?b�^�Q�����G��ۍ"���i�v�7㝌�G{7��ۛz����BՅf}~^Ԧ�}��/��`�_�ç���=l�xZ�L���ݩ����dS�^�6s*�"������i )��R����oR'+�t�ʜ�kެ�[�*b���<�X�^n��\^z��eg +�,�Z4ߍ�V1ꂬ��6��������9�������7���,�ٿT���\B$a��cT��P��
j�=����^�j�hC�hTb:��0�V���z_�>�2O�;�Xb���UÎ٥~ͯq�<��O�#ss�t-I��[]ݙ{fK� D�����;;BtP�.�X�r�5/Y(���I��ݐ|{M��*��O�}�gƘ�?��驽��oXU]�mx�Źî�vqƖ����d:��B�B�0:F��d��V?���3>B�f�7#z+BSlÝ}P��6�D��:ei��t����1���>���f�~�bcح�Ne���kȒ���9������U��nk�w�n�E�yk����r��I��\sU�j������$U����)8?,{wL�]���g��iv�4�D>�A_�vj�e�eڀP��4�gN��N��}^�5�t=��}�^���{J�U���K�ur��!��
��Y��az�7o��TECʪ��{�����y)V?_���x! ��TYӄ���fk��,�M�R�M|� mC�됥�:��W~^��oR�D=��n����٦�x}D��^U�ޘ|����0)׋ {��"�k?:%�s�L��3jǣ±�l��4��~�{� ����F�xeB�_ـ��:�UU1W�� ���ĉ}�e.�<��Ԯ���ˍ1���~�]��V��X
v�y��J𜂪_q�f�4��U1�^�v�ٞ��Y%��pE�]��'�mK< ��u|�(��4卛,T�Fl�;D�B��♇Nz�窽!�`�6�1��~�x�X����ץ������ +�{2�@.�n�ڬx���;[��I��b!]e�3�_�����w��"�Uע"Ŭ_[�3��b�Ɍ�e;�SN�z�"Bn��x5f��Θ������RR�\(1�n2о>��bi�^����F�c��k;����T/4	�4g%�ȅ��>�<�V�t��J��
�@E^���#�u�<,L��z^�J�����k�r|P������ThH�ڟ�U}�?R�[�:�}*z�=Qh���x_]�u�}Y�kL��aTL��E����y~dw�6w��u��[�?T\��o�_Ŋ6V�E�a�
L�{�Bi{E�	��aA��#��;}3s�"�/�-,Bkz�}��)#�('2�k��צԧ�]��<.B�n�͜n<�M�V����n��3	�5�ac�eg/����o��f���K��7÷��wQ��aiWZ��z}*����.��l�`�� �W�qp��p�y�]L̓M�/��|�[��Aoh�*P�z���!Llzb5<?W�m�T��V��]ى�6w�g����v�������+�Ϫ{�~\lxS���Ƹ��#�G}��p�5R��DЃ�0�I�u^O�V�V�k�G2s�'�/��:/�{���`t��p����˽�.��BI���������2OI\��U���X���b�p�[����Z_V�vL�\=�n�t���x��I�cJ���h�唫w� �;�a"�p���𷩓���7N��q�a�Nuf��4�zP�m=xAw���w��*���%�`������N��d��&a��Tx#�oz���wt���j��vF_jC�jү�I�tŊ���L��㠾�,0��Xy�� �{X�wJ$�x�W�B��.SFܺ�o��,���#�J��a�'�.�^�7p}�|b�!�R�n�]�.�t�:$���&���6g�7X#Qt)6��Y��9�vW$+������A:���-U[�נ-��V�W�w�̆�*JYr�2�f�h��gG���B\�!��
ە����`�����[X�U�lk�4�@-5�{�7~Y��u�y�ꂩ1�l(�q�c�E��1M]1W���ΉÂ�±�}�������)4��^�r7o˴�EV���5O�lV�����W�L���5u�1�������������+.�Z�X�P�oj��������#e(�I�̦>��R��Pw�;^�s6=��3jc��;%vɯ�ާC���n��nv>�����B�߱��T���N�{�)���=���M:��5¬�=�K1�(������� �ُ��Z\+��;��/���2_�xP��S��e�Q�͙���=�='�q�Z���Y��{�{���;)��^����2
]3��z��Gvp!Ӿg�:t�^0F�I)�;;|��8�[�H�������m��D�gn�Kƽ�̝��(!dR��{D��ٻ�y��y�}rKT�@>L�f����{:H{�U5���~]o�����N{/
<K�d�zL�5P�u�[�e�۾c^Z�7��L�D�zplZ�
�̅�}G�z��IV\����b�¦�	�]ڧ׺�/=�#Q�_���7�:TE|S�u(F'�R�{W�}�u�����YPR4X��h[��X��Z"�����q��K9:o��GPS��ݸKD��LЧ�X.�ug�����D�&7�xx]�\-����z|z3|��K��b��S��;;��pߩ}���:��=����w��"�IGa�,,*#G��C�/s�96�Ю�Xq�#� %���sqj@0�bDT!��Sس�vW�q�T�j:�{���?��Ӿ�PUr��ְ�:ԏ� W�[T������k�D9�_a�&Ú��z�qA��^Znխ�=��r\l��'���/:��(����t<��o�b��d7�3��OR]��:OH�� ��ۼ��=6ϼ��t 1S�U��ʆ�>[�^t�:S4N�K,��OC-]x��m��w.���Yگ[�|,�:A���+��Z� ���K}�F,ݯFL�H��I��JS��o;-i�C��+�U��y�6x,(_��fVr�	S�^e���P�c[|c��Q��7�Wf/x�+�^m!q/6�����`����o/�1�3 ���mO�w����zr�+{���C"���G=��-�����u�t�V��4\��Lx_<P��o��H1Vǹ�`添��:n��i|M���#ﾏ��8�l�1W�����V�3����/��w��,��R���N}�[��m�᯳$3|؞[�=^����#C\ꓰ� �A[���2#6<�E+E��J�X=y^1~}nξ=ὼ:dC��*��Z��Y��#UدKnO��g{��Uo�����C���qi����{��3�ݐ�}�`�6�*�¶�����l<�����B���+�;��w/�W�9=��OA-
�*�Z�*������u�����+�l{4�dGmϒ͙�n��M%~_�]��ڼ�t�4��:;6�#&�bb�*}j�z�b<�Hx?�zk���ݳ�Z9��bS�@%Qoމs�!�J�e�銩��~^D۠�HM�Y��S����n�g���c�T�z�	J��>>,D�#��H^v@�����'�s��gn�r����qO-�s�/N����� _F�P�e'�t^˹�k����%W�?""�<~k�y�E�>�h�3��֎�S;�o�j��3������u
�������gIaò�g̍�Ka�Vn0
7��h�iĻ���եrųg%�u��}]8�y,�Ʋ�]����D[Chm)f��Fd�:j�9��^��X����q1/ϴ�*s��'��������e����A%`|���k�Yǰg�i��W�b�<�;�X��B
�����諭��J>����4A�v$�x]�bǧ��˭���bο:�%^�Ut�b�'T`����`%Ec�̟�T!g���z�{%xJ6�� @a���E���Z���+����\6�^_���\\�).��������E��Yg~�G�O���׎�W�� �?�V��� ��-!d龻��!��a�)��}�+���<~?%�y�Ә�pZ߂ןmz3��~���{|4�'����n�n���r���lo�7\�/�z*���ƴ���x׉�>�������L>���W�J��x���0��*��Oo$%_/	T7M-���=� ��ٳ:�N���{��tg�2l�F�J�_t}��%ňM`�Vg��Oz��_�dap����06����]⿞���K�,@vut��[� >�|����5�q��_�=�/'��b�;��W�\j���\3 x�O�ǧB���Z��e�sdcD�_d}v�����K7D����sddQ�Aӎ��|�57��b�攠�P�2HS���~��v9zڐӿa�*+��J�ĕ�Α�tോ=0��o�p��\_gE�EҴ+\�$]���箶��t�Y�9�V��Ϗ���ʻ���V<s��U�:vy�׬�γz�.x�h�q�T��R�5 �XgW2rJW����� :��mHsi��v�i�-2��~���ﾯ�9ֹ9�z^g��w׵E��8a�ֳ�v�<�"��Ԋ��A�^��ꕺuòQ�P�d[�<^ޖW����T����&$.���o�K�;��wy�ү�zۤ ٝ��~/x�O��r�v���\)`�*�u���x���5��P�R1s?k�����Lc�l�|���1�t�_׵� T����c�� �Wn�E�8X�V���kQ;I�Y�;�i@�Ն�%x�L:6�̞2P���\G�rM֋Hk��=��b����ԯD1b�~t69�kہ�ٯ�6���D1�#��=����v9[�נ_cl�~���iuL:����~��70�k0��| T�*��X�,Hf|����DEC�#}6^S�6}�������omJ��c���N��Ȍ� �Ҡ*�l�d�X�f���Cö�7=�E��wF���Z7/���[�z�,֪}��a�u�҃���B�����ᡚ�[�=���>�<��;�vp7F�!���p�m���,�C��V�V~�GV�Ϣ%)��Z�Z�ZXL]-��S]����xNWs��{r�@��;���{O޹���GphOt�9�b�OGhp����\I�+E�������;�;�u�%9��,�,�F��Z���+1o=�fl��n#�ǑՇ\�-#|�x�a�����w"����;���q_p!���$|G7�G�(�z�C�vk��W6�J�U����M!����ܼ�L�h'�C{�%�PÝsȌ��|�L�'|'gS�U���~]��]i������
8�w"�[�r|�>�v��svVJ�������&=��i��}�{�"oǌ���Y��ܶN�I��p8����3æi����"��Ϻ_A���	嚝jǆ
`�i���p�<������8J�Z�,eѴ����=����Rn�i�x�ٽF5Wh,�1�5yJ��9:ď�qY��o��֬�*���iǜ�Mo �* �!;ā�ѠaƏQ��F�2,,��IT|]�k/f����Ӕyp���]����Z�v���N�"p�@{���p6���05�k,��&���,��<�5����V8A=I�s@��9�6�Wc��7��ٷc����
C�rkR���V)`�(��rM����x��P��� W��s�b#Onu��у{nk��y�w_$����Y�N�9UڲH߲I�y{7�1��E�f�g���oe���s�i��e�<��w'AY����{z�V���(�3S��RJ���gܗ�c�Ǥ"��=Y���Q��t�4�ܶ��(�l!�|F�x;�zm,3{(�����;?d��a��6���%��ţ�g�a�O.rC4A�y+D,q���_+Ky��>�O�:�zq�6�\9��F�ƶ)�����<3�p��1{�z@;�?E��;g��|�73�b����$���8p⥳�ʹ�t�jS�W}�F휬t7r��������[ER���)^�����ŝ[+P7�wc��q8W�0��ҽ�7�.�F��{ۧ�{R���)�5on�2��c4Ǩ��t���|.�^s���]{*N��\�����=e�&��(9�n��i�{�w����0!ɵbҙ���{:N}�/>>Y�"�T) +n�� �Uc�ⷳ�r��Gb����.��lT�i�6��,�}$�0�)]����F���w�Bz!
��t�z�	C�w<\%�-��x���V��V�-<=�'��um.��U�G'�Cֽ��kF����d�n%�1� ݾ���[�1��-�Fj��n�#F��t;;N݆]G��(�Ա}�`EjTɈ�jF4د���^ޤj���N>�r��i���gy��-b;ٷO{A}R�^}e��r�TM��I�ݚ��������ok%�ag�1Bӷ��Ğ6`�����9g�ho\��6vv��.+�M�]����<��om�}D�F��Ed�$V�\���I�q�
�F㸮W"�����]t*q��J1�U�"��vEJ,�"*�q9BU¨���XV�d&��T)�̒
�� ����U\2J�E�UJ�i��U:	�"�2��!EG(���&QE�(��EW*��R"��+P��2:I�B���:bF�b&a���
�r%�8DY�T�K˩�\�t�r�)D�d�PU�Z
$DUU�ք��EEU2�fAȂ.ʮN$�<I2�E2�r*�
0���TU\��bȪ� ���*	$� �,�QE�D��³"�A�Qª��(�Ȩ����Eg*��Q��
*�#��ȫ�TE@��\%)ĔA"hP�( ��^��{�K�|���w��[�h�����-��t���v���[q��q�Xƥi�)���-z��}�BK���}���>����e<�)��j��ӽ?1'���z���ʮ\���������O �]h?A�x>;��=�v%��u��vus55VW�*߹.^d���~�xz?vv�&�?}X�γ�����,���m���uv�xJ�0F����O|��Sp�}."��]7[JN~2�y�w����*u�'��HaK[���y��t��qlȉ��7��E��y��چYS��9�b��wi�"�c�����WM����`+��MY�M���U����+�/O|'?<J^����w.��7�p�����m!]�k�x��I_�z�玝��$]�s�]5�$���r�mD7pb�9���ּ�����{�&מ��x��k�.��<af��Q��)�mM���xjW����k~�5eK�o���CZ���^�֬z��2� �g�궶[���*y�oL�<'�I�h�Y��rwR�5|1�]ye;��{�*��9�}&�q�[�x%��*�$um	5M�,&&��ˑ4t�Ev�tԝ�&�|��9�}8vQYx����� �É����#�����zJG,w�ˮ΃˞�q��3�>��Oi�m�o��_��{O���?<������^[�w����2.��yʗ*U�\�:��{[���?���i��ƾ�S:�����_�vһ˕:�Y�Eڽ3�O#���ݖ^�vv����V��]K��Wϫ	'�5e�a�f?G��%	�_��N�6���M�ڇCL/V���(Ցu�;da���V7z�V�z���'�P����#sӱ+�ګ���{3�
��T���+��;h��{y)W����T�I�F�����Z�D��+��ג��Z�u�?�g���;�}��5��ׅ-���硯���JȠ���Ƽ�1~��~k��!Ss/��g���G}�S����/��ǤD�u /U+��+<YJ���n��7p6i��註[5mm}~F��? d��o�k�|z��s���N-Q�����˥Y��Vk{<���z�������Wx���0��S���G���x�ĊF7κ���}ݧZ�]�-�J��x�)v��(�x�bPn�0�N�r�{�5gG��c�(�͋a Ηyz�zg'|n�W��6��&s>8��Z֑�pF|����<1���=�:i�U}��US��'?��P���;�n��v+(�5T�Ƭ��.]=7�J��+Th�o��㓦����)n:��ڀ���\m7�U�b����k^{�o�pMu�Sk �W����͵���&?���j��!՜�us
�o
&[^�y�� ъ�:1'�N���v)/L��9�?�ʕB�N5��m�
�a/v�u>ko�Nzd����.M�1�!�w�	�����ɻ���{2ĜT���z.�v8�t���K��wj��W
~F�+�ZA.��,̳;�O]m��֣��8���Ѫ�����~��;^�^��yk񴂗p���^��3C�JɾǴ�\x��������[5~���mx^���m�����㛨�t����,הyVK�}���r�׿:YQ~�����m��g?,��E�ovk�F5Ue��x�N4�7�S��w��[-�}�u���N]�o1 p� .Յ�]���h���K�c���_� �]��+Qq�"���O�~���хY9'֮�K�j!z��n�3�w��t��q�LTVYB'�;��TC]����M�W'�}Qf:��ǝ9ࢶ���PQ݋��Ώ�����T��x�끞V�a��K�,�YٵDt����{�N���5��=O4��;_��?�6��{Ւ�O骲�|�~�6����%	������s���s��e�&�{��w�+�kë�����J��
��9�,��`.q��}흿v���ϗ��:���5u;���{q!E �Ӌ�ɉq�m�u�{Z���R��/=�w-CT�/��v��S���k+�+k#�FR��i�����|�o�.����m�rSi�5.ő�����&|�VZt���ur��A*�7^��;O	�4��5V��������5���+ͯy�U��VUolr��{)z$��<����HW4S2�=Ggk����ǩB������Bn��D(zbd��D�y_Ͱ2�r��U�{��d�������Uz�eVTzFJ?6[�7F��O�W���~d$��)�pn�{�_u:�<���v������2��#�[�:���|���.�31�����g�K�vg�D�N�mj#&�W�Ws��W	h�ԟy����A�����vl�����5���κ�鹉/Y~:��in���\��1;�r���&����п}}�E27c�ޡ���h�퉌)�lڊL<xYN�2��� ��W�^B��#7����3�;�ZAm.���*b��ƫy�ٯ��u&���oL�S~��t��=���Vu����i<�]K��'�;<;��"�K��Erǅ�}�ؓ�{��<���v6��Ҽ����V�U}��X�WU���	��Ĭ�d�����w;� �4��A���(�x����>��@C�	�+XZ�:�Q�Z�kY�s��zy��G����^ޕذƷ4z�<�"��ޯSҤ�E2Y��{��۔gz5�^2�v7Ҳ��S�	uw�V��'-��N榜��z��T}�~;�N�U>~f?=�g�R{8��G��D�S\��S��s5ۋi�?Y�4���Lv���q��^��k�X+ǈ>�:�����i	�+ݴ�>f���g�6zW�ėm���D����x]��k�"������t�z�g7 bcCN��LQY��;B7υ�S�����,T��xWoW3YؚZ�#y?�1��c�Z�_��@g�8v�jE݁���iC�����HVk�W��Xy^A����J�A)кpL���g)���߷������2k�^8v�_o�}n��^vV��ݨT�5�+YD�&��y%|y���8���^%���Н�e���6��f��U�������?jH��8:�ʅ�w6w)�IN����1�3����S�)�0չ�;j"d����i;���-ë�3��N];}����dz;j�ؓ��6[�Q?�;6G.�r��d^����ޞ�Ax$G%�i��]E罰_A�L3�b���mb�
^Q+�SaeZ�h��;��W�񳫥�� ��4�7��G��-&|q�;�H�^.�P����큧^�/hs��Z�m)��������z���C�
��P��N%ת�j����o��=�V��ؕ����rכ�+j��]¸���}��xyo9Y��%'���Mk�W�&�lnC�G��Հ�T@�	��=J�fz��f�GNwݸ���5	'R�r�<���
n����ʤ#��D�p���pE�%���,z{C%V6�t<#}�ؼN]{���	��Y���활)b.�뎭R����`Ư�Qq� ��2/��z��/R��Y�k��P��@t`t����r�	)]M0	�)q�H���91�|��N�[�X�������޹��v�X�������#ak��J��kq\ʧ�/�n�ǧڊڲ�[��Ci�{!\8����g�i3�~=�~;�ڝ#�EavԾ.���~^m�a���qB��ë��ů9V�O@}��Ϸo��R����>��T|\$�~��eI����_�k~����Л=^ܬ����/��_tP��/7UO����bP�۱Z�-C^��h��GpW���ҹ�n����uqO�eO{�Y�,u㰚��N��R�0�CFٯ��2y��fwf5ޫu�Rz�N�e�f4��vkQ:�b��R��į����'3�+�Swa«ڽ� 2r�m?,�}�_���<&�bc��'�X��=�Ğ^�YNy 7��>��b\~�a�>v3�ޙ�
JV�a�۫�!�ߊ������O��k��B _{��ڡ��B+�֐[��1i�o���^����a�+T5��G���2K�UI��u��;����N��)~���P��z4G�.D���:� ����l�6�*ٺ�Hn }Rb�G���2-�)n��H�qU�TzzW���Ɠ �>3��>��e���źo,�.N�>������;s����~�������+�s�{�~�����_����k����v�f'=t�X��T*�N�B�Zu��N�Rz�,�C���oyN{�k��{��j��T��AS��^�#3���8�~����km/R�O�}S���?>5�紽݃4�{[�)�sZךFc�x+��˷,y�G�9�����k��\u����j�i��k-���R7�Y���K�����)*�X�z�<��������놪��6ىm)��|V\7:��٪Uק���&;�
Yv6EqY��=�����^�t��'{��w+�}*^��Da^�p�X�h�Ჩ��q��4�OQ��=&���^.�w�ߗ��!]��9�.��R���/A��?v��L�M���Ԙ�^yW<������'JN��8ݻqt����y����]�-o�	�f:���c)'	�"t��7	E.���rz.�͘e�ʮ���!�@bR�]f�:�̨�jӦ�sOWj8}�#�Λ����o�˰�o��'oV�[��j�@,e�""Z��)Ьs���ղGq�Q���*ݣ�΍#�<���M%�b���3>����E^w��m��u����e	^���+�y;�r�E�[�ʫ�{%�+�gz3e�q�vG�U=U�C���V�^��|�����I����p�Y��(�V���/W��N)�c�	���7�s4T=���~V	�^l�-�����;���n?�.��3��u�[�7U���p�Y9�z(���&'�N���x���}K����ٵ�a��~,�'�{s4ҿY�+�����⾈�"��Aj�/k�5��}3��<�ݗ礞�0,���[#�9oN3��}����f����Z�m'�K�s��Ꝟ�z�O�*o��m�^<�8��䯙�bW��\�qycʋq��?d9�o,d��/�ZC�=׳Q�X�Y�����[�����kJ�����V*2$��N�E�,ï�~�5<[�ON]=+���/�y�w	\�MT�~4�jg���|��O==��=c���m?N�5�x(��`3�ӱV������"�eD�h�/�c�o4�����hխ*���*��0˚,��t{�uZw�fg[�G�֢#����w9�r_����sȿOe,xĨD�w ��6菾�ﾎ�R�ok
�?yy��M�KqQ���=���m=��e[p�W��e0"�$몣U庞��|w=�"�����IG}��J|�׋�:mה�eևS3H�YƵ^m�q釾�:��ߞr&��G�}��w/����kw����g���z�j:o��א��K�e�����'��y-��&+BqR)Xs6��WY��:�5�Un�VQ�u{��T�4��<uU��JxP��+8��@�̚�������cY��pP�6�n���eCW ����Զ\xTl1:�c��F�ˍ�n\�C1��X�!MA�����ݟ�:�}�NQ��]9ȷ�%<���]�}�_������{�ҋgk+�-���9�xA����@_��/ƿ6��u1�/�;��zǲq�ѿCMVa���ī֋���� Ү-~F�"��Aj�1��L�Sі��6��n�+�>Sws�j�h�	P'w�n�e�fۋ���f��`��Ǉ��₩ꐁ��w�6%��#1�O�諾Q�
6�8c�gz�,�ym�q׌�&qЎ֣���r��S
V����-�O@�t��l�����3�/8�S5ȱ��f�!k��w����z#Z�no�֘rJKїc8T�'��cv�����'�`�'� �Y��^��G����7���r=���M�SV�ݯC�d��84�yQ�	�������ss޾:m�6����R�S�C��R��Gм=7|��]��U�-�ba�fq����b��W�e�\�:8��`��������'mZ�������s��u9L�<����n��U��Nm�sh��#������5#���"/��l�
t@(��-F��̕����˫��(�N|x�$r����+B���	�go|�0i'�����Qg.�	�sN�K�۴�-�U�e�j�SKO)��E��U�$�"���u�Uv��+ڃ��8�b��*�ξ{Q���Nt���6,nz$��۞@�1n]k|M��*�p{F;���^cGv�V;}���:E�G���꛺	2ňc�3&��k%���(L��ދ��+���7�I�����jq������$��0���ղ#t�9�D���g�Yz��u-�9�Id�{�B������l��)�*�Z���@�P����ځ�L��VZ{�)�OOJg�]��ǣ�NwMbw:c"������6n�Ӏ�(�c��v����)
���6�*��r]���,p��	��<���b������L�ǂ��i�!X�7.:��ئ���[���k� ָ�"Ȓ�Ն]f*qg��u�yW�S�(;�ڼT��q,�w�t�N�{�}����+Np~��(��fS"󑂐�\�M+3aLV�f*ХM�h���1;��W�����dkéd����ͱ(?�a�CX ��C�G5m��:۔/6��b���8N��Z�e
�a��y]�̂�^l���r�����B��x�煫��n�0_Q|�f��P�%-�/����)3	Aˤ���e��yB,�tU!F��6��Ku�"6g<*�y�ȯ�k��Wqm�Ѳ�R�m��r��c�w	r��Lh`�h��cwL(g�8wǇr��"P����\�K4!��߷�ֲ�<	�G����Q��"�#���Y�.����yc�w�3j�j��`�:�ʞ����Ͷ������%�lX쵗��s��h��-�Y���M�-�'XbEՒ���],�7����2��P`y{�����ϵ	��T8���k��E�|�TE�i%����a�ҵ�W��R�{�T!:3��ئN�A^>�R��^�|��Kr�V�j����"� EQW�*�EȪ"
M,�L$ȎA@D�8J,����"
�(�W�"�"'M���"��A��9r9�"�SD�) ��ADD�#$4El_Ԡ�����\����*�b�UAt��Es��GIVU�c�yǙ�*���UQU&DdU9&TUr9E�" �EK�,�,B)���:#���$���$�AUr
9Qj(�Q�#J"�^AeT���[H�Ȩ�/{�l�g"9�k<u�\(�^P�!Y��'��<w��U&rL�bDT\��9^Q�B"�*(""�G(�Q�B��J�""DUDp��U���*ÔTr� ��W9G�r��(9��R��B�Q8�'��* ��>��*�n*��1��L���l�=վ�2ȿ*H�/vs'��ħ$X.^�s�,�e7�VkҎ���"kqG�E�ﾈ�� ?y��Oq�6U9o��ƻ��^�k�e�|�UW���)�����u��������ە<̬�l�9�����k�[g�bW��\�字�@�/������I���럘��'N�]�w�ߗ�{�\��J���zN�f�=2/ys�>k7���q�;���s�=8�_7��#��*�Ol�+��N���8Sj���*�K�H���RU����؆�Ȅ��\��Ӛ����o.{���ߜ�{:�rxk��[TL���4�f�}I��x�����Π�N��|��;���:*v�uy���^r����*!�	n^Y~���;6ճ=Q��8�t��,�K~�Ƭ�t}_F�!B��՜��7��w��&;W�}�ۈ���]}���j��	g�I�x�o�3lj�2x�S��Dّ%~8��jw�54������05�
3n���B]8��ŵ��Y=����B��7Y�1��
�f_ �8%ϕ���qqf�i\0����7yb�Y8z�2@��1*$��I�L�=�m�8���I�]*��7\����wmު�C��FYх��Y~���K�s�r�Ek�������G���z��߆�����Ua�%]��_eR~��T�W���G|���7��<q�Pl]O�P���Đ'ӗ�i�eL�Ϡ�g��;����A�9�,����� �W�����<��z��]�^>��W��*mo���z���������{-���d?�6�V��n��F��̝z/��J&�[6�_���?[W3��e�J�o#/t2���/`Χ�m�T �E��,�S��5]�P��᩼�{޸���#ms�F�=��?-��ּ�X�WR�~)�
�<6�˶��y�I��^�	o���N�{:��b�g�ȵˎmrǚG�;�߷'N�Z�W�׉�2�V�%9�y�{�F����)��gf��ƞ�>W�Jó\��;�22%�Nj�WI�Y�I��^��X�J�T,��Av��DKw�\#�2�[�Q�no%�f�+?eĖѩ99��e�-_���k�^~{���l�T4VLɦy/
�qU�L�u��r�6�ڦd��'I�P[�����fm�(��q�[���}�:�ո�p���m�Ԋw̃�EWl>O;�齛K�}�� ��(����+XEu��j�����݄7�U������}�&w���l�n��'~|�y���N���}�^y^���rڛ�`]��e"�95�w_^�li��u�������1���(v��L$�r���i]���m����Է�2"~��6���h�ּ���{���ߩ]��^<�^�gBrx�X��t�*ryD{}	�=�����B+Lg����1{aa�2r7V���Z��<�	]=u<��YTO!���v���[��T?S^�Pi�F������qcr�(�m*���[BW���������$�Ϗ/gOV�|�S�4�������ok>gB�JQ�'Kw
n$��QP�	�~��*����:5W�Z�Pۙ{�$�t��K@~��2�n�����������P�Fn��"���U�5i���g˨<���]V���f�O����{�6��[xٺ��9��98��z�����H-�Խ�������ڜ����>���EV�����읺��:V	��K�mҵ�J)�9��!�e=fl�a��,�S�;�qT:2C���}7�z�Z<�Xudl�U.�����t����-5�]y��-d���;^97�f3������]{�����>�����|/Ry�r����i<]G���o�W^��{nk�M���I)��]�����}���z���J�\3�dZ�G_��q����-g���l�lK�e�4�Jq�G7T�'�Z����	y�v�a��J�r���S��m����x�3�zC�����d�́)q��E�weB�86��������Nw̠���יJ��^�}�YӾ}�w��)��6�a�,�h�'K�nd_��Ff�*�yV�3��IG}�Ϳ�/(�/�~�8��l8y>��S�{V ��U׽�*�j����r&�A��6���<؞^�KN���Kv�{3��)�yӮ�L���W�53Kqm{<�oMu}㙊<���ک���n"w؂��	 �^��e�V!7�v�Q<��xX�=�p.�}���G�wYO����jjk���G��N`l-`��N�oO���ߎ�G���F\�ͱ]��f��^BX؞yX��ܨ�$$PS�b2�S�:*�W��������
�Vc/U>�/Xɽ�DΌ҇��%<~3[ͥ�f)=���&��K6j����ʉ���\.tТ��=o���`;���b=�=)�����ʵ� �OJ��E��}����"ȹ�;ޞ�*o�Z�����^Cꞕ��VE���3��8.ğ!���z�@�2q/*�ی̙1��&<�����p�m��L��r����y�w`?��uM�v��4"^?���uK�U<����}m#�$[�nN������0��FB���3A�����ߗy���2z���o�9�>��6�c����3Bϟ�����j��^�vw�_��3����D�찀����ͼ�f�{�(N�����>T������D	��Ak�T��ڙŭAn�5q��%�����4����ڥ��rW<���p$2���ۃ|�x��z���k�6����Ŏ�~����w{GH��w8��8��]����G�w�j�j�
�
�������#��wO�i��!���QzN}OA��q��t3��5|����������YT�*�&x���=���27�9��G�ı��[�sy���t�!���S�~�1���V��r���Z( 賷@�%�s��<��P.A�ho��w\�F4���*䊱�D�;�����i�奍�+���ͅ������UU�N�_9ݲ�Q����q���q�+W�aC�F����m�n>�2/%k�̤{v��+U���o����Ūt�+�ܯK=1�.i`9��CSwN�o�I~Ȭ�q~j��D��?�J�AT�C[G .u7�|@_���s���UG���D���{�z7��>��M��V�����1=� �:N�ٕ��j��Rd�̫O2{HGڀ�^ʖ,�]�F�b��Ng���i�`�T%zmP�/���I 3��ٯ�#��N�3��ٯV�.v���lNT)N�M���fKP��N?	�Y{O���yqrٕ���O���&���G�d��[B�ۙ���o��x�s�rX��{^�ơô.�Ԑ��?0�)��1z�^ڞ>^��� $}����x�t�Z�צ]���~�.f��D��]K�O�N�=���)�}��"�{�o�] ޞ̆]�b����SI���6�^�G�J�H\2�Y�E���!��kW��v����1��+<�6�^����2�	Q�f�2yG�ّ��k�֍]�3}���=���_�~������֢�1"��	�����T�Ϲ ;��QI�v6�*N޺�U��J�?}��}UH��'I��_���Sl��Z�~��|��d�Wي-ra'�}鍊*�f��Ε~���̯$���+�X{_2�6�g�ˎr�zqc�����Mr���5�C
,�7�ǫ����3�bE��d�Uǎq�|��YL|�4�X�1�6�ͣijZ��Y���rӃ�*�6���]N�=ʽ^%zvE2Y������4~M`���w+�j�:���5�������8O��*߉�oǺi��S�5�/���J�]����C�&�ů��h��Iғ�3��,)�?Y�6��}���s~����;X����s�M�Xgo�c�Thv�^��
|�Q^>D՞�+�6�d@"=�L���zX�x�Z�G��`��6��B�0bZ��Byf�'���H�s
��֏.�}:��}_��K��o�~�N`l=|�a�?$@ߎ�F�|��V�{z�ty�]>��ٿ��m�<(Eז�Wn
:kXr��.���m\�lZA^��j61At��+_oY[�W]:�$ i�}gB���z0%�v�z]�ȸ��W��\�<��ܔ�$Zʞ���o�`^����O/x�����x���34���d��;OW�D�kefg�$�]8���R�c��w�����-�WUnfv��������CU������X��K��~��X��*��_lڊ�0ߥ���Q�$�nK[w�1���a�@��Ù�Ao��WRx�eF���z�˙c�5n*w�&δ�=��ͪQ�rA�U������c�m.��Ly*��t�k����o�כ�7�Og�^�mrW�����k+���Ǟ����EL7�C��؞f�=��~�T�'�M%�q�n��Y�7�o�^�k]����S�$����U���Q����w>�SӗOO�:F�%�c����]�yN�GwvOw.4�ԵT>5�{!�/{�������3��,>��v)�kCT��\�����ru7iQ3�h�C������͝>��y�r��w�x�z�$�ս��X�!� R�&&�#;ފ$���Yx�S`Ʀ�1-��{5ğ;Կe�W��*��'�{@~�e�.2�B]�H �l�3�[���ܱ��ݾ���B�5�3��|� ;sgy4��KZ;u����@5u�w��U��V������N�?}�5q{8�ݿ!+���c��=�BP��I~ ����9'+��ǥ���v��t���]�a��Ƭ�P������V(��3I�v���襛�*e߽�>�A�eD$�U�U����ߺqνw7K�٢AP].B��?{�Y��=�3I�H�U�ؘ*��}9	Rq��Q�c׊�
/�^+7���ӛI /'W�&_?X3�=�	��^R�Fi���.�?w�3��*oh~K�ߍ6�ϗ+�����.�_��"��
��!V�B�Ӧ׭۟+���sˣ�h�5B%������auy�_Z�ҕ�J��L��6����>�͞G~�@���G���"��.�s{��y��vFFE^�U��x���ů3�<��;��������k��"����"��@�u�-l{3b��'U9����Ͳ��[g�bW�s��ʒ}����K��'r�S�N7,W;)3q=�F���ur��s�f	L�-o�C�@��G��H?^�l|1��w/�f**�",��bvI�+1��F���˖�82��T��/:��Vmg�-*7���Z�u�U���(���=��;��	D����>��Z��v����[�sӆ�c�v����5�O��7���^�D�1��9�wK�o;�Xhx���5���d�X��k�4�n�ƕ����p/1��L~罓}��5u�p���U���*��6�����ڙH�����m�z�6=+֜j��,i�o]�0,�n���L����Gg����
�Rw}KV��n<��'f�or��?&[��Z��	TC�.6��
�-v�,���[w�ל�r�m�<�����R�,�o�S�W�$~~1����+���"�,s��=����̀�zQo���߯��ο*�`²�`�`�z���ܳC�~z�FO|E.f���<����v�/pY6���Qq���r�������JV���È�+�A�����'�f�{��j�e�S�H�c��h����=�{��ޠ�=��v�R�7�1�_{W�$��t��_E~3ޭe�l��B��f�*��]n�CRо��SO:N2�ut��3��q�N]�tT$�r:�y��M~�z�w�m��do`����
�䊗pd�%5`�}��31��˖�
�v�6�k8#�I��n�/p���wV��;R�R$�/�S,wGV6M���&��=�7s��F#�t�w{_���	 F<���1��F�wʸu:N-�t4�4-�c+s;lK:�#tͦ��m^	�ʅJt�=��az+p7a��NLr�sh�U	0�|3S��흼RӅ�Q�g���W@-6'�_QlbLˣ���q����<(ߟ/c>k�	�����r��<ݝ����3�M�xJG�ښ�) �i�v�n��g?t�3w�{پx
��B���w�.��r���6_zi�X6�}�Z�[y�8ٴH�mY�h|���gu�WX�k�������>2q��[�_�=w�O5&�'��^k����h��xx(!��j���K�3�2�&6�r�1�1����M���"��+4��8� +�<�n9�cv�_9���#��r�c�Ү�v�5�=�/���୴!F�Ʋ2�d*��7�;S����"VV����>p��&MgT������c9V��jO�RA%���>�]\m~ЄU���m�:��LW���޷D�W����Ԫze!/,ٓB�ׇwμ�kD�R�ǒ�V���#E����3���xZJ券��S�� f��� �̜s��,v�Y�gg������Pq�4���aW��Q��!�,Ng8.r�ٯf����(][j�����VP7�o������3�d�R��9��xS2��̃8�7/]��nYgh��t��i�w7{��`b��OmM:���2���N����C���$P諥���'잴�����C�q})�b��-O�n�L���Om6�B22n�̍��w��++(svk��l��Th�����m��I���8Z�f��0��'j�؞"�[�]�e6&I$bjnC�3$Sl��0��ި1)0��JH&
7�L������w�^�ʳZ�h쬨���,�h�� ��$�g�����w�Т��8V>]���YK��v�+*u���|)�6M�\�>׏���7�3k'x�b���������-��L@6����}���gk�ỽSf��/6�Ύ���AG]$s���ėh=Ю�$j���F������.n��,ڢ��h8G�{1��2I��������ga�A�u��KG�9�+�����s,W !b-i���9&�I��eY�wQ���,p��\ӑF5�!vz_�e�vU((��\v[b���Z��q��!��K4~� !9�!%'�,�{Q;�br�ԷzT��1�'�v�Ӹ%��M���k7��yǄ�n�O��a��w�|���Y�¢��WN7����t����'���cM<��B�k;N�o�%� ����m�B^����<��W���;��yӊ��eTA��AՅң���D��x�w"2���r9L��.DDW�(��TB�Ĺ��$f�����S4R�->�U*�<�j%F�q�0�2��qs���Ȣ��cu׎��E]�n+đEQ�W"�I������]�UQ���u��I��W�A��Qˑ�9˼�)�,ʹÜ�r��+�%9f�e�U��6�:�)P�IQC��
�M

���w0�q��I�ȾPu�U��3b�H�dsw�;�����)�x�8��p�A
"�Ak���I\5���[2X{p�ܴ-*׏Z��s�=wU�4���(r�C�.8Q\�$
"�	�H�fQ�iÜ���S�
��*��6�Y\f���:V�m��gy�PT�ي�.�y�0]�Ԩf9���dߟ��`�����Ԃѻ��QtȎ��U_Wв}W���|���Am]�{x:����.��Oy ��kΤk�3��ˣbzY��3&��/�a0�6[�St��g�@�TK��CF۹V�K���c:Ej�z}�^��Q1[�N5�癸�tbٜ������Zg��y����Z������^����:p�n,�I����ӑ�'q��k�eCU�g�<^X�iu.w⪟P�<#�]����.����M��N��W3��'q�o��Y\����m���9��[�W)l5}��}���$�OWy�
��oa�ګ�\��c^5C�s���J�yb�G�~���#�o�U����hK��goݒ����C7e��(��ѳp��5�ν������;QG���:?���^��T��t׷^2�Ӄ�)���ڙo���h�M��վ�u������z>�8�0$�+gmz ��ǅg�{oS�4������m�ئ�Z�轾Cqܙ���i�κ��<��w��,\.��F�@��3��ڰ�9R�浟�XW�c7�tW���ɲyz���
'��9���lSS��^t]�+k�*b	�����}�}\O����_��MB�?`+眉���zD���S����z���2�%*���p��6�zj��y
a�Kה]x�ބ��gͿ';�a¤@ȷ���/C�n[�U�b�am9�y~��^����W��D�̒�Y���]~�����F�	S�q�:r"�212|���r;W��
�F����ۙq��5�o�iưJq��t��G��3*����|<.n�ɚ��K7}hM޸�ɓ~|�ڥ_l�~��:r�C��GD77R�s��o�"v<���/�]�~{@�ƭ �w�e.����V�bOS�R��EbU�E�箾���K���]_�R�^��>�ԫ��;��a�o�n�s��{	U霡�>ͤ�*��.YԝgQ����V�ͥԻlS�����e ������oz�P���x�����'W�/c>�ۇC����U� ��j� �!�Y5*�-���4i��8inmo�c���#�ҳ^�V/p�x�O�-�y![r���^0_�;yo���-t�6é��s���ݘI~R�������NktY9��}��잴h��X���`�TV����]�}�}L���Ou����݇��8�e|��}-%��O5/dJ-�c���S�]����5�f�Y��:;���1Q׫ֵ��s=B�K�qK`��s��e�I=�꣊�5SUeq�[�{���);�J�1Q�Os�y��P T�:73s��bM��^{���iOW����`�q��3�k��7���:F��u���9*x���޸������J�kۋi�"l�T}���o�5�Nt������WWn'qW٫B���~�Jk��*�0������z�v֥� ���}$��S�ݞ���y�e$�[�a�j�c���=�����^-��7�T�tDّ%~'�3���&�>î��+Ǫ�����bW�yu9��/S�q"��Wk8'}�=S�'��a%*Ǯ4����nwd���~�Rm���/$��.Vy}2�*��jF���bu�F��� .��[�/�a0��]�i��8M�.`兑�U�)�SqV���b� ���Ìx7Vq�'-����<��:Qұt��&Y9��Z��n�.����fnD)<��儆]g-S{@�
�~�s�%��>�����ץ��z�װ\������M}�G�>�\N�ϳҗ������6;}^�OK��I{�gz�eʛ���uO#�z �\7��("�դ-���=��a�y��/{��9��=O�t��n+�A��f�?]C^��y�yQ���ݦ�0g;������{6��s�M�go�t��S|���{ܭ�W����h��������9g�k��7�Vx�~ժi?*Or�/{yx)�	��6�]^�{�}���,�X�h�Nv���޽S���wEﶝ�S{"Rj犓ƽ/����w�*߹.͢:y�q�z�Z��ҷ�wQ�O}�ӟq��<j�Ͻ^���us3Ug���h�eo�����X�4�r��{]�Iҥ������L��m��F�5q�|G�ݮ�ӎ�'��>�|{ű�FzmQ]o��ٸ�ǜx�:S_&YW鄮>T^xZ�m{Uַ*�kx�hB����E����W��
H��Fq��ҳ�ɸ�8�o��1}7T�������
]�w2�G�|���&���O�����x�@H���\V	�A����e�S@#�U�!�n[���_VM�FW�}U��[��:w�����[3���j/��ט���F����:�Z����R��Q�,�e��|��� [�{�Y�<u>;A50Q�Rǡ=��r���Ij�lS�;�gL�����]V�*-<�U�V˓�꼫DH��i�{]U�8	B�.'D�n��l=3'{�^u�zgW�Q�Y��N��v�-��Q�!bJ}��q���\���&x�Q��zs����^�N��H�z�vJ�Q���tߡ��n�e����6Nz�G=W�����Ͻ7;�;�5i��u�'Kz)ǣPf!�٤�n	�{r�'�NON���-���.�A2�z�RϧP���oyBuK%������kZ=ϸ����~��lzJ�3��>�X9��:�R��Ե�i� N���p����Ǚ~bo%}�+�����\sk�<߈����s�bW�S!Mة;�N䝨�'VY�<Ҙ�j^�u���e{��@5��i���s�|�����A�Ƨ�gN�-����Z������_�y��-��j�<Ŏ�{(ٽZ�SI{_��0��m�ꅣI��n�+/��x;�˾��i����S=P7�g��o9��kT��ĭܸO'w�J���Ϡ�-7Mtr��71H��S[~��W���X�����$�K�w}+-�*�EB���J�@�?{�81*þ��{�ѐת�^ʋ���)��X|�{0^jn�nJZ�<����e�{��R��6f�מU�Oxm�ƽ"��+��R>����G�s����7�=�{i	�B���)�5�ů9Vz>��-��^wIH�dA�,��|q�:֋��F*��U�v��^��Q~>D՞�+�c����^Ǭ{��%+�6�j7F�*�`²���F5Զ�<Ez�>O���{Of!���$8�,ۣ���;���ڀ�^ˍ���9����M Du�ۺ�b��wx�{�̸���W�ʕ_;'�ĺ�e��Sp~j܁�>�-�y��z��|���H�n�>Y�'��O�?mR�p��gaζ�"��4{xᲥ������O;\�VS"
�E�.7��^n�{}@b[�o��Xf.��2謫�;�%��|�L�o�\�.�űI�F����%>��5E�M4�2�~���55Z�_��ÉvE
*��d�'6���n,b���7m��inmK@O7	e�8��K������ǽ��m>-@��B�h^����cг�Ǽ�����}�k�;^w���]PE��ZAj�^��y��~��]�^�o3��y�o��g#���C����˪*���\ŝ9 �����N+Fr��Q�9�Y�������ON"o��No��"�}��J󝳑�qP�~Z��K�Y���%{��S_Bk�^����~T!J�/�=�,سs4�7y��p�<�j!��a���J�U���pa2gC鷘:JΩ�OIg|��a���[[��W��F��'�-�G��� �hｭ�FuG��~�3�q�j�f�WnׇW37�<�ZL��=����%s��'��8�$m��q*�/��ܸ��+�[���w�5~;�͜+n�Z��B\�N��6�V��/7UJ�׃iCqN��{Ƕ��{����m]u
���E��"n˩�wO׾�aR��������+U��P����Ub�o�q�5�5�v�||i���~���@wBwu���D�P�k���l�J�{�9ȗ��ߦ�IK��3ޫ؛ �G��չt����8�������]���̬��^N�
��^ʅ����x�-N�ՠ�<ʆ� <>�FШ��5U^oVF�z�׉�UY����~�J�A��=�6���8v����g�W��=�g5��~H��|�_�|�`��Oӣ^r;�n	E���VZ�@Ïc��z,.s�ߛ@:\�e.�}2��j�V��n�u��M�?�`x�)�p_�<㖀�#B%�_�_���#'DN;�.Ϥ��G(Ï����e��맾������'�j��+s��'\��2S��ɬ؝*;qQ�7�g�������ًG�.�L%����]���ҙ��K��US�;|6�|�g��Ձ��J���[Ì�W���;����ykͯ,x��O��~�S���.�W0�7�s3
���������k��1�Ɨ�������:v֒s3Vfׇ[��H�x��^h J�zh[;�&��{�3F2���t�D��`�{���Z�9;����>�^*��@�#b��I\=�zGܼ���u��Z��S�A]��X�%�0Ȣ�B`j��C�+�5�:�ŠV�>�~q��o�U��w�JK}ض��U�݇����xҮK�H���|��dm��פr��>ހ��=����ܰOO��3��^�����U�3ʯޭ��}%��G�� Y\��������>�Qyd'M��JW鄘P�3F�nf���n��Ej�{<�~&A��m%}��n/yz��������ש��t��qZ��}�E�"�g���kzWx��|��תu�������J~�G��2�r����S�~���|uY�I_�y�hG�"�fS�r\pt����͌���esCԱWoޖ!�f*"r`��DeF�^&�<ˀ��/N���7��1��l��d%_N�l��q�+�j���{W�$sm�s>`��{�`�{�%���nT�@�|�K�io״��3�uzh���R,��u,U���+�͵�'*1`�oIw��n[Ȯ}C�����*���4����p�r��f��Ε�G�>*V^c��V̹%P�Rހ�o��S��Xً���/U���S���`v1��t *�5};����5/j���η���O*6�	�mՇ�,�b�oӨ�f�e����}\|5V����Ue����H-^�T��L��L^�����)z���������#�!��X#Ar�����Խ�>���{=��a�1�-a6|�*�N7oM{}�Ռ�������E��:��N���V^�*x��5H��U�9�)U��o��X��8���#}6���U�r���&�<�!	�b�v�2ue^�r��ͣ�T�i�ä{޸���oa��Q��rz{��V\�>pޠ��Q��V�)lb�x���w���y[qZo%#����9��F�z>�{��d1W#ٷ��zy���h��w�/�0|����v����p�s���#���W���}��r~���W��^Tn�#߽�J�=ͫލ��m��!#�c[�����kf����X&q�����e�)�Z����`vᭋv+(��W�i
��-����D���ez�~@��$���
�F�trmk:
��q���*fC|;R�g_]2���f��k�ϻH�Ǧ�pev[R`K���>��h7��Ht�T	�=T��B��k�S
�o�ƭ��Y9�K��&�,�:�A�m�!��6���o!���%pZ.��6�L�6=�a�Xmu岯����U�l�
���;mIa&3���.�t���䢐�`7Vt��h�`cY9�]�;����'�m@QWx�6A1&vh�;2���e��Jqp�&u�u=1+��t.��gR~Ҟ�J	֐���f�#�T�NG=n�dŇpA}�0�4~��s]�n�Jک�����xNQ��7	D4��\��yԴ��v����Ss��`-j�TX٤N�f�TN rVo`s��xض�/�1�xMs�Z(���4������d�g��@�9Y��"ꫵY�=v��g7�,�}B�g��!��<�ٽϔ�d�{�{��
	^����X�S�hb<�&�άG��^K0ň\��ݍyH�(Ցp��*�����؅��oa��Ow���:�V�u���7
V��T� 8r�S�*{9g��s
u۝�8Pu�]��x��E�@<1�ԾtFb$uLB��1"o��^�7I2��|4*�2ݰ4S:Eb ���Fn�Q�ْ����^>[�������tL�}�֠��@dU���y�ɓw������<�ǧt&���P��b�w�*�>^ʐo,w�W%�Y�\V�qI��Y����΀�7
����VS
�{v)��S��v�#X���b��b"`���K(���V�P���n�B�<��5�`�if4\ᵼ54��]G�q%�G�̋a<�@k)��۰(\���%J�k{fHm[tF[���wc)q\m�V�n�`+�={�.��w���M�d�`��ښ��Wb	5m���\U�W��=���x0�GI�ݴgg>�e¯�9��\�� [�{[Et�W�CUB��w����!��>q�U��3}O�:%�/.����Zs��m�a�P\�qХur�e٤�B+�a�q�!
��A�z�Z�1ܜ��Y���=�
�|��Ь�Kh��嗗��|�������qW��o7��	~���L�EU��*�Z:�����-��6�7��.��6����Ɲ����3���<��v��`t;���&U���sM�n�/DT������L�������>;Y/�������[��r/�_l"���uU��jR��ݪkut'1N���}�`�^�&�-m��a��f��Rw���},���+o ����LWys8H�w�����)�sð�iu�N*�މ��Թ��Mub|hn5��0�� ��5�{ľ>�y��!�>�$��օT�v��Z/f�a��ݤ�+��j�N��9vz�/X��*���ϙ˄W/�K��9Y��2��|�fL�U�A��W�#�rL�"�AK�����"VkT�0�2��3ä%e�I*.S"���{�*�Re�һw�kpz����/
E;�**��N:��-P��.ˑQx�r���3Z�(��,��`Et�^E�q(�B¾$�.Q�;y�Ǩ5(Nn<��Q�0�q	��0�QĈn�)ʙn�x�%�\]"�
����Qǜ���Y$�-T�D�EDX�E�\����<x�!�9ơÔV��.�s�8E3r���\E�#��VT�UE��q"��AE�Ȋ\����Ȫ:t���b"t�"�h'���NX�.QE5Jysqyˈ������1K���U ,я���pw*�)�ј��Re�ξr"�q�b��\��q|>�7s�Q��d�-:�t�P�x�oX+;�s�"J��_}�Z/��ϸ���<ʉ�T���n�n`�P����Q��|k�x�Y飖���vN�(z���+1�1�;Aƺ�K���)S���z���jo";\��܋��C���9�ޙ6��+�i�[�{-Ҝ����P�b�=ޞg�V*o@��`�?6.�OIW��e8凞`{m{����~�'���;�T� gu{����BK�֑�}�U_Q�^�ytS}6��[�,�����\�j۶+��Q�Q3�q�2�m�̛���ɸ�dgJ�bQ5�J���^�%
Ԝ��;��@z`9{������;=��2ovs�ϧw�E;��e^��W��}Ewkӥ�w���Cs�O$@͸�!e�0�;���W�W�*��,�G����q�9oR��b	m��!ﮯr��>��{롸N��v�{7�ǓT�Q=��j�c��4���q2j�Ίg��n�R[�����F��dGc�E[�N����]>�%���ϗ�=�(p�.t�&�����RW����~\��n�z� �9Y�я`���uƇ;�v�+��2�zA���'�Q<W`�=���V�ɗdv]lz+����48�Ov�+<M���|%���vB!A��׉Ö��҆���:#�M7l�wnٶ2|������+bKK٧���vw�:�M�@<:��瞀���v#�C|}f���{��)a��lr���^Gz�KS�Ol�n�\J�/ю�w=,��U�� �)�oŹL,+�=~���&�^gH�q�{��]��ɨ}}q��,��cцsxU ��wC4�鱑��d�%:��2�oi��{�s��m�d��ӧT����с˓�����`���P��h\���9���C�,�O�S�@����N�g)��8'n!����$d?S7�72�,{h�ys�^�s���ڏХ�乥k�~�s0~���%�fn�f�e� 1Dd���L�|k��Kٍ-�'�œd#��43�W�t��fx��K��}2�5
���d�Gl��ωP�yR��+�ϰ��7@W��\d�*(L��}Օ���l��������U���bɟ�]�׹���3�)ꊗ*g�oOe�q�Q�-��\���Ӿ�5�����dK̝�u�������;�;�OC��[p��:�S=<{����]�����L��#c���?C_��;u���kO�o�Y��ا��`9�;�"9�i��m��Rwgx�A��^e�ֱ�%���	�
>������v���7^��e�3���~�v�����P���N�;�.�����J��Q�=_a�]6"��S9&��z�\�%�do�>������ڕ�N��O��(a���0�9��\��g��S�����s�[^,:����'�?���_�f����n1�3��ٮ�)��7�d��u��}��cw�OVb�܍9��W��[�ﺫJ>vde|���W�U�o�9��'�o12���F`)9�*��A)hio0��Ů�S�ݴ��<d5�k�	k����E[ʭ���Rs�Hl��c���=��h��d�C�c��+�"Է��J�|�l�^�:�S�l�Ϋ���S����p�1�[|
]ͽ���L��o�q�Ŋ�wu�����_A|�:�*��m���}���˅v����3Y��{YW}Y��H�/dߊ�W���si�B�5�S�<=�>��p���p�Hl��;��c�zr������kw�}�t0_ʖX�Rn<x5q���ON��Hwf֌}nȻ5�1?c�힕5��U�ў���9�I����L��n<cn�s��.'�	�6:�q˦���[#Μ��.����H��WT���a}�
s�ˠ3���x'܎d�L�MgmGB;j��ֳϲ�g=�y�&�*��27)�O�u<���[��d�P�6�%���������+�(�lL�m�殠�7�qm6�V���^fy6fo�����RsC7�K�CIj�K���s����;��%+'&��ۭ?p{�G&����}~~(�m�5�_n�艟)�7M��u�����0=�W�~;�w�l����N�~Y� ��ד!�Y� ��oWC���3Q��N�`9�=�t� k�t�A�3$�~λ���J[�ȷ�q^��8����L�φ�m!��L�_":�����hwz��
��"����z˦�����ԇ�����C5�^]!������8*��"K�:�$7<Ϫ����W}����$Y�}2�^�)�E�	Ó�Qޝ9�~�ro��}:n6� �����'�"�'��~y�Uޣ'�y��ʧ�����)��|��M�=��u�����q��yc�&�ݎ���E�c|����g�6G}~�϶���ѱ�2�ݜ��w�u܏W�*�j㲫h�9eO����G�?m�k��Π�����o��k�O�g��0=�~׮�/ċ{�Co-;yQ��8���Yۨg�T�"WJ�i!����ǓT�P�O��\w�T��~�T��Q�c+�&r_�z,{�3[������&���WT�e��h5/Y�_{���r�8<��VK�ٻ����Ozf��!�&�5R^�㐈k�=�{s}���vC2�wf��1�<��3d�+MNv>���A(�Ⱥ�U}����3N���5�҈q��iG7Vc�h�ݘzt��\��V�RcB�9A�@:�p@e�XĻ(�oI�f���W��i�}��E9N�(�ugﾂU��կ7����8�5��ݖ�2�M�x��m���迓<y�O-���W�j6+/Z��]�����˞���k��>�Vhe�O=�ާ�o�G�1�unɟL�\o-і;�����K���N
�[�==��/�$��0�Nw�uC/i�@�(��G������ʌ���U}�*��Ģ�eO���W=됦Q�7���Ϣh�{e���_���e�U��znݏ�3wui.�W	aW۵����b�%��6����蚇�]R�T���ߪ/�8���� �\����C���EǼ�l����xT,4��z���G�w� =}�7��G{Þ�>9'r��}j�1=�4j�yx��Od�^���:���"Gt��N��q{��^�5i� �ZVD���=)��Ŕ�d�]~݉�U�})]����G�����z}c{BW�	s��n�Y��q	e_u/'N�e�~�aÆ�_L���u�Ϋ��v�2�Ú�i�ih^Y��I�5L�ߣ���[��YDυ�P�=��2og����LDUq�Pp}���r�2����:{�R0��^*S�FLzM�f��;c��Šk�
fn��p!1n%�pX��]�/��X৳N��+�c�׵�{�-����^�w�:���c"�a|=kl�H�}k�B[��'�u*�ب�q%�?��G���y_�9`t�F��0.y�������/��ݟ%;���@[��>�L񬉜ת��� �]OFq���X>N끴{%k6;3���(y��ͱqezu�7��ثW�_�zg{.�rks�t.;*����@N��c/z�Wɪ`�=��ݰ�]�PJ9]�c��c��j͞���:�"���KPj<���K���<O�������{�f2ݯtmV�Z���;i;���\�Ω�!�`=>�Y�;�����^�����	�C�>��=1՞=;�e�Fέ+'#Q��h�7	S�H
�^�f����� ��9?{��}L����ɛ����ښ��W�\R���잌��_w_\u�x��0[�ô�G]��z��e���Sנmw�^����`^��T�G��9��ѫ��7d��pFC����������Z���/Η�M�^6��C�*�D��z㞸ӻ,Yݮ3}8'i��ǻމmNT]����@MI����֯��G��#qH��D�]�^�DϟȘw;��Sr�i&���Hi�?�eA�o<�E��\�!������*�s��ɣ'�#���xՔ���s��K�����s87����`����|�>]!qA�H���.�m�ˣ���zD�6/��y�$͘��08A��SA[��_�¦�4g��Bou�o��~��~�X�U@J#�W�&��ݢr���3Q�y=��饗5ô8����91��Rw�9���{�g�ʀ*[�;\�\�\d�:(\A5Z�2>����ݭ2j>��I3E��S��{��E/nj\GP1�L�n���Up�@~�'��\����9�r���A�̞ݹ��vϣ߽==�J^����JtI��@�i�p��A��=�n!q�Ū��/L��v�,�w�x�3*o�Mm�����[�^�@g���q���`F��Q���-3��^Sp�+�������w����ʃ���&����M��5����;ێ��U7���{\ ��@d9����.�眊�}5�R�%^�Nﲐ����%J;�dc�ۊ�Iʝ�p���xe��@W�q�4G��Ȟ��Ǹ׍��,{'��MO�{h���ʐס���W�:� ��=<��1~'�8߅�NE퇖����~J�ҮW+Q����$x7ƾ/��wa�:�:�Z�A��6���z�H��H����qЫ3�x��C'�F���LX����kg#���|�;�e1��讹r�_�	�>�.d]F΍���"���%��yת�2�Qʷz]v�T3<2k/ۚ�'$yR0ę4�5�E�������3{PM�y^�}#�a��۷|kZ�3����1��aUӽȯ��im�Q�/bX�r�[��,)7�c밼�eY��ହH�nL�2�Xڽ��N����8/�}�u[V�=����O$�x�~<�_��s&��g�������2�]��0�3�e��y+�k���j�d�����`_�Z�x�j�X5��ݝL���R<<{���x�|RC˩j8���5�$������O����������Dߌc�{v���SS��D��^��}�9g76�B}���!�M��K2+��v:X����_w��{�}��H���.3uW7q�2��x��u���d�L�,������ȧꮩU ��q�];��@m{�򦁗��R��{�׷�R�Ni;ѥ�0:B���7@S�ˣ Z��5MV���Qg*��9u]��Z�׷�~��A3^G���2���)�����(���\��Iv��]yg@�+P�SZ��
=�5P�2$�d���gf��k)�
�Z&\������Gt��ӝ�7왊��S��v���
�1R*��`��;Qޛ��ˇ�}9��t�F� �]\-����Ck�wd���U�%Ne���Y^�&��{��&��M�~f*�L,X��k���n���Yۄ~*�:dgg?A)r=x�Jef��K-�.�jJ�]���Zg�bǹ�W�~ƽ��%��Z��FS�y��������1y��N�P�"�;/��%��ӈ
Ť#���Z��g���}�����Y��n��N�)�vxv֎~��.:����u܏Sʽ��ʭ�;�*0 GT�z��nfv�r��<䇖��1�ċs���>�C�첥y���z�r�ċ}eWL�>`*����\�ڕئ�Bڮ���KR�d<߶�XM�<��ʛ~��8�5Fp�r��|3�;��mg��}w�W���4.;*�Mǉav���u�v��<�鯝*C�[śC�/�tۊ��j���ݛB�ۢ�z�G�dw�,�.�cİ����<�k��p[v��|TW�6-W��zƇ�-�K�=/ђCf����f�^��@�>'���Y�}0�t���Vdr5B�0��OD�Y+�����ݡ��u=�s���Q#�ﶝ���O��O�x^�ǻ/����a��*�pr�ͩ�Sq�GK��w�@����C�'��bp<YvE��? <uǸ���槷���w/�R�N`�n֎�v��9�Ң%�򨜇f����[��Vw��Q�Ѫ���۱���ˑ����Y�7bX��=3¡a�7O��<���@��g{gx+��x1y���5q�x��x�����6	���/27Ř��n=B<�+�[����s�/�0(��%�K��Y���$l�\��)��Ô8�=�Ңm�uU�niy�D�ٽ��v ��*�op&<A9���$��V���vV�;$���r����x�Z]�����r��v'?��A!cӄ��x���P�6MTj��#z�3��G���^�*���Ꚍ}@���劯M�Y >܎�kV�x<����j�WP��~ŉ�J���ؑu��Jx�ߋ�Kv�*��O��kJ1�����@�:�c�٠�zh�Q·K��V�����0��q��I<�=��J���,�v:�r��x���R��MB��]f�}����F�2�m��Fl��.�:��MX;��PǠ��h�ӡ ���=�0-�{l�V�v{�9��[��F};����^���Iwv�k���u}:=9��7�@ν�;.6�:<
G�[F�m���S�v��ډ'�{�d<��{.�̼��d�v?]�v�~����c7��5Lg�{8F�ǷA������J�Yk�+���,+�ЦY�
V��q�T|�碭�Sq�x.��a�ucЯdn��r3���CF��s��3��;�=�˕q�r-zK῕�Gy�\<�t|$7ƨE��Y��5�&���K����v*#ҹ�����js��^��}�s|] ���Ws�8��l��ǝ~�yF��2�(M[(��lHY��T67��a�h�gs����z��'�ZD�!��w���l�U g��O#��}�D�Q(v���q���FmB�T�w��N�N�7.X*��o��#�lc��������������n���`���\��`6��a�d;9�lp�ѣJwu9��U�$ɋ.�`�k}��O^�aY�����T��X5�����;t Z�����;f���^���h{4r��U�5�;fr�ͬ5�O/m�հ��6�����u���=\2�,[8��|��h������fEw���h�{=���}1���~��`Vr0��iWD^��"�m�e�6k��g�(�X�(���V4��Ru���d#���$���|b�����l�|B�iF��+���:�#$��v�,���C�<?)y�-Mc�(u5Z>fY��f븅���"���r�@~v�.r"RUw���$���k�+9ML8���P2��*�}�l�"��)R��⳷�Þ{�0�L���Xx�(�9���ṷWWDa��\Ph�$	s���h̞�q�4��{�ӻ�ے�^Ny��W�d��xʃ|#�K)G�F��t����h]�Xo���e��*����d�N�e,��g5j�dF�А�3�9��&�wY�e:�:���k��֜�K%�XX���@��N>�$q��<��U|5��P��@���S���~�14>��҆
 ÃA~g\��->xf]���
��A�7�Bg��/t�gA�N�
����(R#��=���B�@
	�v�PI����ӎ)�4���d֑CN�G� T���^�V�V�;�����!ͬ{��- 2���>�3A���,�u�c�UB�ʄ�ok}�_�r��Zs�]!�l�F��E�X�ރ&�017����P��_�Jn�c�ۦ��R�{-���I$�����2J��h���!^�|�I�����$x�qMJ������/G��Z�Rd�����V�z$�xz�h�틬�n�D^Ӣz��4@��Émf'�b펚���֨j�sF��@�g�+d��'#��2�[��Q<�z%) �|�o��z�=�(Yh���Β�&��	��t�6�/��;�s��)�N:� ���C������V���]��ϩ~Ta���͐�em���;ES#�̧25(>�}�e�@%sX����Dg�;�,��b�鱓�NK�]/��bnf
C�A��n��]��}IG�5^d��tj���1�X���%�(۾�h:0'i�ݴ�J{�7\8�q22�F�B1�G�[Ww+���g<w=4,�Rp��|�ɷ�ݞ~� l�hp�ۖ�L�����L~���UpX��D�7�t
��˴��+����J��y,4;��z\��|����=�1�\bMGp'd��
��o ��Ymp���<��+�\t,���.<�;��s��w��Er�(S��r"�$�����U=dS���	^$v�5w���U����5�x�R��#�p����:�Y�����X��ü�v��4r��*�H���Qήnp�tW�E8�ss�Ċ�-ÜN[���݂s�dU��\l��p����%ibe�&��*�D��p����"t+��<`^9{�Q垷E�ItG9#�WR�S��xv��]�p�bIn:��/#�s��Y9��K����H��-P�GQ˕�Xbi��\��"L�ԥ
���/,\�:�Z�UETe�F�*�"��]YbF��G<�5y�N%ТO9˜��x�{
�=�<i�KB���Q+Tq�TyE�R�;��ȉȃ�B�۽�u�2/G�'5�2�L6�B�y2S�z�q�}��W
ݺ0Y�M�o�W�T��Bx��B�yk�֧�3�.�lw_��S��g�=�P���ee�K1-�aTu�����"�;��M^ח-�Ъ��D�R�[�~�����k��7�@���ߠ�ǍC��R�W����k3Et+^�x��Ox����e��*�Y�	}V��Rl�Y�y���؇�<=�X+��n��Ù�oQK�@臹7K�̀v����<���|��`0�9�xb�Js��&Z�HRx�(�i���xր��+���/�9\&�������mfC�~��o���H��jЮË��55��|x���hvx��T:P�'\��+-��&�V�����ئs���m"�zG��s�
�P��1O��M5Uý�~�*;��.H���A����{�;�Us�Ťe����Ht{F7������r��vo�GD���F�\pR����wU�����L��ǙF���t~˜���?L��7�m5��A�_�??g7L*܁�<B.g��R��<~����5g|*�0���`�<ɽ��捝�粕���+���|̬�?M�Q����+M�e��Ss�]�^�/9h��0��.yn3E-�$�l���{@��8z�M�/W_['z�����@�Sgm���d�Q�C��e�,��~�
��O����c��6riõ�l���I�p�̆�c���a��8��9nZ؂����q��X�;X���Q��M3Ü�C!�cU�[�3�ww�fS����}��M��?�J�}�����y5��炴m�oW����{&�9�֧�}C�di<1)�F�d.n3�Gz�+�pw��O�9�}�������ʐי�]~� ~�eӞ�����;)�#:�m\k���{������#\��മ6��\��3�E9�^��+�]�݇Q>˜����v���#�c�%�~�6�۶<.;��O�8���ʣ��0���MN�n�=���YF�=��/���w�W�Բ@�x�&���zhs�MR�k<�}{&�}}q�V�{'��=(��7��{6w�w�$r7�%������y`_�Z�q<��.F���٩N�r��d&
	X�o�ZW|�z�^������ټ$���C.6�=��N���c�~ݨ~�ك sW7���vrg�o�����f������G{�r*��H�GK
0�Nw�tTw��{�'܎d�oK�p��]�9�[W\jz3v�o�����;����>���@}�#Ѥ禎���n���X"�l��Kq{��^쩡а�����Q�<Q��!q��=���
�����eA�>���k���1WK�a�.��X�NG�E7^5�w��7;sj�㋗�s�V�b�$g�[Isu�h�E\8�n�7s�ؤ��sU�԰�PD�j�V������ux��(5gM4/0%+�&(�S*W.Y���_\�{po=�'������&k�3��Og���
G�>�x�==������Ц8�����f굳�v�h7�э���̘�Gn�ٿ��k�8W��_șr)�����?ooh�>7��|��5W�ӳf��I ��Дr�m�d�_��3(��K��{L Uup��Ef�����(�{dwʩ�������6+����ٟ����z�/}�8o�q� �Swꛁ��v?j�G+��T�mH�����¶3��\s̲7g#��u܏Sʽ����(/��z)[�gj�d{l����p
-q"��c6_z���r����Sq�}z%�j�l�K��.�{R]�m���nUmM����In6�XM�ύ�i\o�}�T�0⛬���zm�I�Z�kn͙�N��]���h\<�u7�X]��s�h?v�S��ޯ[��a׷n�=W�L�#��mODQ��ų#P�dG{����e:���S��<�Jײ�p�%]�}^�����\�}ǆ	�u�ee/�$6o��XO�Y��_�;%}��><�B�O�W%��y��uؤS��G'eJ��|$T�.50o_y���t��<k�T۴���	}o0��3:[�B[��T��0%��%��x��{�|�0ɲ�|�t�J�2*/7v>�8�+��>��}�W:��Ɓ�ZJ�v4�������|�zq�է��3����
3�
���c��]R�H�a��t̋«E�c��z-?o�l����R���=�8ٿn�;��v��*W�.���O�N���r���-o���갼�I���S��v�^DO�,��÷N��r���zt�g��UG���k�@����:*�k�g�zʽz�z�Ɏ�ec����n��Yd_���|���<.2J���:xQY9-����#�b����xq�GˠL�h0:>.�Fɪ����#{3�L�z^OU���
�P,T.3S�@�!l
��ԑ�E������o�'j���;� �t:U�47��ˇ���&k%�ɨʇӤ}ٍ�Tg��8Uz�ۜ�FeT���@���ހ�V9\�G:/g�Ump�|s/�Ç	����y�me��!�'���*7�I�H�z{��ޫ�<g���\���펼�NT�j��f��)�;��&���|�ߠ\����������1�y����MnN]�������po9�k�#�-�?��L�TV�����h���`	�p6�d��u��^��"�[�p~�f�v���+�
>=�!4�.�=�-��ݱ���W)����>���d���)�8��J�5��Y]p�j���������뻅1ݘ�����վ���%��b��9�!o:'/�Z�[��iLyӑ�z9x��d�{R�w�}@v�����Oq���G����q�9}�h1���v�vUmM��	��D1���X�&����Ws��{�W��ekUs�]����`�� �;���{�� �x��V�ө���t�#Ia�e�k>Wb�7gyN+��콟r-��J�{��\�FuH�3L��+8}瞁p���δ����'f�{:�ve뮱���f^�������Fq{7���]*�/�2���~�wC=�8d�]��T��R��	�� ���=���W�c�Ӵ�/^�l��N������,{�sv��&���=���>˺j�d�����+�t4Ol迥ul������z({�Ἧ���
F�,r�v�z�G+z���?"v����h,��?O\iݖ. ��7���$�=◐'kV_ /����<jCq\��n&k)��y�j�^������^~�RE�J}#���?5�ݞg)�}k�� {��t��9u�Q��lQz���f�/'�\���Pu,�Kn��z6��VmMM6@]6WPnn�5�n�P�B���s�YX;s��8*g�"�Ǹ�������`Ut1}vy*��C�t��tmPw�IB�p�xo��]��מ�{�� ���}��+�f������Ĥ� }����$���=y�ˬ�rx��]�u�<ϴr�u~�����=�7�ă2�tt:p$Ӟpd/�}��+��o�?�E�j2PH�L�߾}zj<��ΟP�G�H��ߢ���߽מd��)a&�{5��\�5]�����s�N�0mu��C��O���MZ����ΑќVZ�u>�'��?e�/�Y!��Pz����9�<0�`$i�ޮ�E��TV���Y����n%~zOCܯK�g�N���{a�@��a�ʭ������3]��t(7%��5(�~縭�d�g�U�g;�to��N��#��d���22����h��.s��zq��]E�n��R�v�Dk)ɸ�xc�|����((�ʐ׻��h��U�C�^�;��UX����b�3���F;�N�>�!���_)��[�e�q�}�\�FuH�7�?(~� �)tD����������~��z�$^�gM�ĵ=��n��b�}��.3�O�G_�m1���樽�<�7��Ɏ���n�\K��<�ۤ��~-ʼ���>������0��*{59�s5���w�Zꋌݿ+�۞���u��G3|J���wC�����ԟO�z�k���;�?D+�\9Ǽ}�#�\��-e`�/>[M�E��V����O6��1
����EH�a*��鄰���%RSMj�1�X�.͚]f���KÜu]��z:�	��0�J�'���UM�|K��"χ���.��T�����R�wS�>�����+^WhY�7���Q}nȸ}\n	�����u���v3�4M��>*ghx+��d�ا�u=>��=
pN�w#���޹ĺ�̎�)��.���u��v��Lx�����'Wet��z#�u�r�M�L��f��_�޹�]R/����������)��NI�yi�ծ��]���h_�Ҷw�	c�*j}<Q�������������� Py��&�Ј�9'j��<MV���j���&k�q�է���b���\o��bȡRg��/���n�V�p�Z Ф�H̓�}釽�gf�Y�'2�p��U.D��5�1���l���F3�}���@긽����e䮿�cY8�a@��A�J���5��Hj���"}�/J�=]Sq��9�I���uT��/L����w�p���8Ǵ^R{x{}�ugx��9c*!�)��j�'3�x{a�Z��ܞ�af�܏L[��33U���'�+�gV�Z��]����t�3�$v\k����y��ac��7�(�¯����g�ih�e�I��w�fx�ٛ�B���X:��nk~�~#�:�J@��5nk�<��GehBp�rpLu��G�^�fΥ��Һ�肽������9x>´��uoo[�a���w]���,�%#��V�
����1S7�����w�w����[���{������f~��P�����b��&����ƾ/��t�G`���*��IF�G���91|���O�3},��v�����з�N��,.[V��lW�i�٪��7���*����Vr� ˨Ύ�sp��U�@��ݖ��)�߉a��m�8K7�$uQT/�H�f����#�uV�������%z˕ &Tw��	���2����>&7�,;o�X!�#9��/z��ʘK���)��{<�:|7�nؿ�2�H�ხw��T0�әA"s�+���i=�z�gA��EG�j�+�o�=�*n<���FMׅ�%�B㮢��3ۜw�Opt�Tצ���o#�1�z��~w����%���v�u�9H��=:n!����q+���S>���U:NKz�UH ���0P��՗#{�,�[<37�X�a�$����g���"�y��uI�ի<�ѝ�@������w��7��^&k��z��ኁ`�8�3��Y~�ft��uno��n]P}.l����A����R$����e��ݻd�d��:�K�Y/��=�$�j.���,�f	����7�a5s��?��K<DƢ9jk7ݔ*�x�o{O�}
αp���s�+l�z�MR-h���p�[�CR�����rcK)r{s�J�sO�G��܋5�@���)�a=�t��F;EMr�W�ιԆ%O���*g��R�U�3��n�E�3�M�'�����z�X7�!R*�u�/g����l�/�=�C�]�.�5��xY��.��B�� [�=5�vUp���~���P%^Y����12�"){3=�^Y}�� �{�FO���c#8�� �w��=�0/�w�kݾ��:��M�;�q͵��`7�xݯ<�?]��Dl���6�쿶� �	�p6�d��כ���7�Ǧol��yP���<�-����w��L��������N��G�����e��X&�ƾ5ʽ���觠��NtߘC;6�^���3a�ޫ����?Iu+��]3��os�1[�U�:ԋݲ�z���X>r��P�+��Ĺ��"���0�S�:߮�>��c7�<�{ا;�GD�z{l�;�wb�ҟ��/&_:Ჲ���:��qt�ױ��<���T����,��x����yʼ���e)�8��g>�c��������e􌶮�N :�=Y�ڧ�r�{���ڮ���O� oǜ��mhvOl迗�ó�T�{�D]���W�y�)h�,�eɮ�`�.-�Sn����9�N�i�|N�n��@A�5I6l���Іn���m���oA��%�l^0	�;�� \c�M}'5�o��݅򧽬F�B���a>T�ݛ��Hs�}��}]��zZ��DqWA��n�C��v0���їt0\uv_��|Z�@�<���wk��-秶Qe�OlT�<�P�D�@���r��c����*�&@]�c.e{�=������^u>�u�y^_��a+��k��: +��*����*��q&�~;���3-"Z���+t
Y����\����~do� �����~�-���w�7���DC��ME::&IN|L{�f`��߬�A%����ǻ���5X�&�xu*�<b�A������
���"obpy~!{7=��7�n�&�#����wVd�}�Z���tI����\p��A����{��W\5<�~�={�b:-<3dZ��r�ێ�NW�X��Qɼg���`i�ޮ�
w(�����&�~L���W�ݯ���ex\s̛ݜ�F}:����eG!�J��3�k�����/R�3�O��hj��:7M䛈�Ke��-�C��vr�;���d�Ǘ������h�t�����6��y�N��@u=O���NM�<1;T�ߢ7�T�g�C^�k	^����F�G���Ѩ)�|<�-G6g,��$|n�Kي�\��0��l�y��3Ï'��^S
�'!{|�1�z�����%L����V�l��_k��"�ҡ����1qhf��#psԍ�&i3�e���[���j��Y^^�;x�پ�ݢ��+�����Zd�8CB�pIn%��ƳîL�'=�	��^�Zĳ���s�&�x]��Kr{��i@�؄�unO3QF�مj�
e�[�M��4���7��<��S��)b����|VC����ڮOYT
��W�ܛ�u��̺�(���{o(t�m:`�$Y�/��X���[<f��=&��e�̯5u^���R���S�6��l�Q�/�3�z��Ք��[�BϽ�k��j[�֣�n���g��h�B��O�E2��kY�j�Ay� Jv?�[ˑ���I�N֒on�e��-�`��K;Ϧ�3���LfZ+hT��#�EPKt��a�y|���s��d�&\�^k���b�̜=n��2o`� a#}��O� �c��ɰw4Ӕ� ������2b%�ܲQ�9`��59]3l���'h�e�Vf=)�3@�L�����޽�h�mz�K�c��l�3n�|�S�:z�{I-P�T�:�qm������&w#�o�(�u����I�l��N�g��k���o&�>y�"��=:��j���I�|_S���S=0/��J�{H/�B�ʋ.1ʄUsb�2��&�d\��rK4�F鋬Oy��bl�V!yp� j��|��>6��*IT3M����=�!�)��;����A��p^gn�V��y\�k˶�y�B<9�{�1�� �CYF�;�v+"$-xV�"%��r�E!�Z��
.,m`��}�H�D��'e��W��?Yh-B�f� .�u7�-Z���gHm�i��m׋����r�t��<��W�q�QYQZ������GE�źe=��2f5��h]���� �����ڂ�.����9[G��n�g����2Y4����Z���tK����hۛ_���F�"L�Μq�ˣ��j{A1�x�u�JK�@C��J�4��g�W�=�魅�~�k�5&""�Uu�|�+N�)g�1ܽ�Ο�@<�v��5�yu'��]b�Si:����K���g�c���s��Hn�(RK>DC�����c�(M wb�*�ݬ���b��KF�JhAQ��O�d�<o!,i��`������͇{��N���^Q���-E�.�b׀t�z�}�p6�^����w�T6��>���t�$'JG�k������3���z�Q�F�ƌ����\����v�ݩ�ǵ�.�$W����K����M�邴������ڼj�}݅Ցj>VG+��v��=��g�OL>>�ٝnU�{��Q��Ŵ{���-�	eX�!h�$7{�5��["�C�q�@�������q�2&NB�W˛���E��T���:j��V��F���-N�1*5Y��P��R�ӧ�e_\��5XN3�AG"�r5$����(�nD�:�Xq&�I���UUD�J�#�9���N<��U)V�"�y��|B2�U��hk�s�Tʕ��RZ��+1J�g��(�3P��J�e!�B��K����RL�L+P�Y�)�J�ĕr�.�\�\N+(�B.Z+�\lB�霹nێ8�+��qX��N-D.�I)���B��N����".\)E��:��U�S$>r�%;Ԏ"��->X��SaZY�9�fK
��gũ%t##"T�UW
��'B"*�Y�b<n�ɒ�FZ*�8����`��ҴB��aIҲ�Hr���dr�5@|h|	�L�tX4*��#��α���TP*��r]/��+�ކ�_����o�RѹL拖�@�˃{dA���;}r��wB=� �&��ۖP�E~�u]F.<KL�d��������x�>n�{�K�y�r-O���5�'�j�vjj���oxa��/Wd��sB�KS��a���,W���[9/&��W�(�F'�ns,��ݺ�7��{�����@=U^7��@���M��+�C���F)휾�ʩm=y}i��שu��^�C�Y/���-�x��}TF
������R}<_z�k�������L�wI�#y��V��T�$P]��/�����p�Hl�$��I϶�=��N?�j]�(J������WB�=�C����O�ԎG�� T?S2+���c�D�띸�]���j�˳D@�emV���P��o	�#�92�5�j:�9T��_K3e� ���"����E�TS5�'҇*A��krr*�o��m���}�@mG�ו4<���Z�B���F2}�A���ӴM�P���rGo�=y��r�̓���u��Dnނf����k�W����ꊇ�.&+t/�=b�̯{�>����ݞ���]̒�����F�g�k2a��ݳ�zΉ5Lp�w\=Pn\�u�o*1��y3��jh@�:��˄��[z�g�[-ё����>r�����**B�����}�
��bx���ٹ�b.ŻM冊���3K{��tM�l�.9�r.K;wKI�����V���}����dYU��gs�R�#Uߩ{՘�9�\ʯk��T�����Дr���vO�{.�fQɸ��ӧl��%�p^�C����Y\@�W��L�dS,OOe�S��^�h����`�zh�3~~"`5�Uݞ��
-O�oe@�N�1��g�){g�o��z.#�e��@�n�\��=�{wVJ���w�#ms]�U�b�3��7$v\k�ʚ�G�y��ިO{,�*�*�U���� �Ouf�L�Ϗ��������𝩹��oIo�E���>7�k��v׽Tҙ��i��k-�|���+{No�G�Y�]���hd<o��>����[<�K���é���BU=�w�:�;*��r�.�����â�{�W���`[̧S��F&+����zf�ד�È��LV>�si�|VQr�$6n8���Y��O=7ѝ�*�_��ll<��^��	�c9��1�}IMN��{�º��(˱ %=�-�Ӊ�g[���]�O��ް�>t��'�P7���n�;���7��x������C����x.��~��hR?&��/k��X�ߌ�ci�g'��Hi�:[y���Ǡ�ʾB��;h�},*Q�>��>9���td}����\�����T<����(͠���4:n��]��O�����Eh����"�=���F�"IQ��n{V�&�Y9I+������흌���yx�V���7c߆ɒ����.ztԷ\��U�>;�����]W�u�/ʖ��<�`uw�K�>�����
�����y��2N��hrx��]��3�|tk����M���r6MTk̃�"7�3<L�z^OU�1�+_K�W����v��W~�6�Ю�X�2g�z���7���ߺ�5]�&v��]��5�^U�C�?����7��l�y~���'V��d��Wt��g���zk���x?U��^� �s���}�V���9��KejPN�<��-�@yG&�t9'OTr��9z{�~]U��r��sˣ8)�bl涨l���
�m/G���>�ў9^��|0�98�{��*w�����E��;}Q�}夵����n)�}'�w�u�����?ہ	�ݭ��L��̭������L ~N끲�x᩾3wW��J��䳛��+�[�s�'1��/'��ɖL_�C��q�U�7�wD1�8E�X���	����+��~�:�@�/'�9�a쒆��ͺ>W���?\VC�N���4H��V��|�0g�9�#]��y��ڈ�Z//��۔i���I��e'�viB��-���f��)��$���,��0KK�ueW��.��1�wS�i�.�t]�Uu�^�w�=1�L���V!}AnE}�K�3���ݜ�n�Am��>�$�o���v��G�K��ϗ�<�s��+�^�u.U��\�~�$�VP����}],��Ϫ��	�
�tc�u7�q�}�a��v*=)�[9/&��|=+(��c��ʇ"5r�T}�¶������`c컡��^q>R����_����;Jc^��Q��5��;ڻ¢d�;|�s��u8���7��DȽ%��S�H�r��CD�΋\vQ���k�3f�	�9}N�p���+�=(�/���0���T��v~���V�=�+��\��`\�f�Y�u����p螴��z2�<+��f�s#�XH��2��W���xz&|��w�b׻�Q�/˼�*蚞��h�%�������}����d
�*��q�loN����o���>5T��^�b��&\l��l�&W��TuoTԮ�N�]@uÛ�*#�����C��s���5R�Q�W�^n�\����v�ɯ�dɚ��:�P�u�����D�������?Pzt��4<O1��Y��RG���Jl���;���~�߶���:$�S �u�D:�P�O�:�.�K��nnۺ����b��m5c��n���v૽�|��:s`	�N�V��Q_,�k/���w��g�O���G_�3s�I�]�ROR��ҷ��j����a�7��/Y�!1o����c�|ƺ���p��דs�g]{>�_�ݣ��_x:����3DSDJ9g���NW�X�}9�c<4�m0r,���j��3�w:��h��3;q��ɸ�~z���`����?}톱��k�oUM� gvO���W�foymk�]@ڨ�ړqǲU�3q��Z.ʝ��|=(�L�'���:�=
�Ǣ���#|=JV��Q�r�r��c�����rwOs}ʟN��*;ʤ5�k	A��ǧ�H<wu�L�^~����\���֢�U'>�!��z�R�L�n[����m�(�G�]!�7`�^�'ط{s�n�[��U��`�o�G�_�Ui{��Py�m��wR�Η��VK��<n���G��D{.�a{��M|����Q���ǼWI��[�~69����<z��:��~���s�^�Ѯ�';�tes��p���p��Cf��\�TG���{ũ7<�ٷ���f�]����Q���������:��uh�����)Ra���l�o'�|j��i_~E�]_��Lj���nw;�'��l߷j���7���:�H�ﮤ+%T��s���ႜ�FhCw�� �R#�T�R�t�(d Xw
�A��W|ub-%�ݕ�0ڦ�� ���}�
���b��66��L�<�Q���)�Wm;][Ew`?moz/g�r�a�W���8�>��n؃c���eRH+{\[s�=��Fɓ�J��`.����mz@��Qӄ���_K3�]@;�u!���H��y�ߎ�E�\p����׼)�uw�/h��n�M��{g|%�iP0�x�<B�pQ��,{b����>�	�frT�h��8�)M�5X;3��o{v�>s��~�ᔍL�P��=�V&<�c"��6�����j��3�յa,��\Pצ���(�M��}&�&nQ��gD�,p��F *�jx9�Y]��^����Ҧ]wU��3�q�&�5΄���Qޝ9�~����NB_���.��z�K����A�( ��:>���]����}��q��l��'ɲ��y�Cُ�{�o�j�R�\g@yG&�%���p=�����C�S�=�p����|�,�ٟTק�)�z��*~��;�^1�m�?V�\���h�9gcd��!���y��adv�y����Mڻ�{׌��qɝs����/*�2�S�з�[S~'��i!���	���qJMn���u�lQK�D�[������ovQS��*�ۣ�,���
��y4-�S���,.�Ն�h��&��_������t��:;�HX�w۩��˨C��k���A�1�m^�����u��v<��&��j���+��Xf�y��x�:�ޚDo�V�1_x+m�v�;�GfZ���8���>pY�<c r�7�'��1a?$"iT�mj#����!�˩9܄�GTr�8��3����E���*���{��y��O����v?�Zj-c��H9n�w�b�_z���͍�+����e�Q�Cf����f�5�i,��1Փu�;�F����Γ~0��Y�w��Jn6^�9�g޷l{�쮩~�$����t:�yO*���j݇�/�H�*W�ވ���#{v��ݾS�lʚ�GJ�w�B���oÊ�a�˞"݇�]��T�����0P{�+��^D����rݭ��\K=:y�0:�fQ���	*=Y�@_g{�5�4�@�*S��f�\��<�=l�Nh�=Q�\g��jEl�s���x�;���~�ݞ�;@�(Q��@릠K#��j�^a�י�&k�K��͔D��R�t���E*T�xtF�8+4�MCd�*�wO��P�T�ȧC�\A�C{D̸m��/���Q�z���6���R�dᄧ!]�������k��SF�r���/'<T�U�\x��M{V7�}a���|0�Á��>��jO��q��5�U­�_��/��S7\���h�`|��
����v�9w`w]~��4Un�"ϲ��+{X^���+�\g�s�N�b��X$���{Y>
%��d�D���P�)C�sF�DE�`A��]�W�8����G)q�]L<i8�e��@V�����LU{�ۼ���rlI�j��V�X�����o(^���+o�zW�{�8M�#8�l�,�������J��Z��t4y�M��oR���v���߾�i]�r^�tU�7k=0~�T١�]�<��i�-�{a{�V磗F��mn�n��g�U����7��L_�0S��u\r�����x��؏q:�'���UI��i��z�SB����{Z�����c����ݱh� σ�u\ *<�T.��^��k�G����U<����Ia޺�P��9�e���*��ĩםR)�4�zF�^��'.I���%����\ܬ�7�._O��7F��Q�O�����n:�2���q�G�dK59L�J�}��x��>�1���a�`g�>S��[����u�v�ƽ=��xg������U���F�Ba�C��v���~X��бg���>�R^Ác����t����O�����տ������^�����z�W9�Dİ��DhϺ�/������q�_{%�5
�9���{�%}y>Q͐��|����D���@�G"���~��f������sl/f��#�o�@�����X��n8�!F|��/�.N��Ӽ�vZ�w��;��_4@�צ[��*s_qZ�j�}�V��tJ�k�����)i�m�º�粰n�܃�/v�A�����^����h��mӞF*��(��6Pt��%ֻ�F���޿x��ӈOXiM�<��� +���,��"���Յһ���{�g�¯*nW�^��WF��3^��[>�~�T:�ꚕ���+�������u�b��οb�9[�u����f��8�ʲ�on֙5���j2_M}
���g�>���Up�z��d1=;^��Y�����S�b��qE���;�U�=�N��ok)���8z�Rv��^�����R��S�̸�|垅�����xE�,��+��_Ƕ�a��Ne�s���i�g�;k������h�H˸�68�>U�q�2ovr:��u��79�ݗ~V����u��{�ֻ��̶狋Vm�XP�	P	�t�C=���êo��6Y�y�/ۮ��U��q��������[�n{��s5�7����xe�P��rn!���V��vS��!�ڿQ����Jr�M-����3�0�����weVы�<��.Z�w���rd��+v�&��N��xtu��������A�ﺽL3�w�W��y"�V9�q�Z��i���1b���kd�n�.z�4��U����G�g�0�7!w�L=�9?����oh#K�oswBt��f�kXpڙǡ��i�gw��1�4&�&ؾ��ې��,��k�[��5+!Ś�Oc��o ��'�'�{�<���𶶻��ܿ\�aķ����U������}��7��]��� g�WI��nUǲ�9͑����|����:��o��*͝Ȗ<__z�N䫎�I��\�TG�}�����RQ�N��A�_z��Y[��]tmhNn�ݛL����+辷d��7�$��L�����e�m���Ն�/_����v���$M��s7��j�ݾ3�:% �Ã�]H.�H��C���ݒ0]�|<8_��j��{^�vl�ˠ2�����O�9��/�Q���Ss/�����wz�./�Vߟ�M��s3ܥ�U���t�;f���۹�%��m���_X�����k�<Q�����W��V��ۨ�|�m9�Rԯ�vM���(�ٿ��A�}�x7�k3n|:���#S,N����쌃���9�K7��Ύ�QL�!���� s��G��G#pMTofI�ɇ�ݳ��tI1蘞��C5��}�Ӭ�vwZ�*@w<����>~6w9��Z>�=��胞ˇ��9@�V���9��.yΩӥ 1S���H�X������/�lds�֜����UQ��#G�9�9����q��f
�<�(n�Cn0�Y�𗵜:ڠ{��pt��`�R%w�-޲��fw�\��^��8��PJ:��S�r��6�N�Z��n{QNc�S�Jʵ��4)��ͼ�,��ݻ��NA�rG��K��jG�	Z�o�k�B��-�lf
{O���AÇÔ����d-��,g�M�Yc
C�NaҲ �gv;9�:�i�W�����vbf��ã
�����8����с���t㺙*��˗�}��n�"3�����v�!�,K��v�T����'ۤ��H3�9&��z8[���2w�-�8..�n;�3�>Cu@n�f{��>��Ä���0�X��vlxV0]�y�����͕n�6g~��=����j�^�����p&��/iаt^�b�k��E�{�Of�w=�~���i]�ڜ[��CB���1Y5���]��7/J�d��u�{�oi,�GT�<A����	W�y�x>6�y��^��l��+��ez*k�r�<-��W��Oa�=+H����	�S��������~W�� }��Y�4��>^�7��昹q½��gk��p07���|BbQ�7B��Cr��Ȳ�\��i��w0����K���[/8���<7����+�9����TrV����ne��N��D��eǞ��O5ͬ���v�F��������J�j��Ye$���t��."�]7��^#:%��Ӭ8
���{-���N��g]ڇT2��t�ɲNN�l&m�d��y&uc�x+��6]�<��DWYD��'�����{�� Vj�*Y�LUhIr���ث)9���}�%�������:*&��=�vHn�^6�;�`T��=�vL�m��ve�F�`j8o��̈�p/$`k4ȝ<�;��{VEg6�
T�]ۗ�B���`a�#���e���#>�AO�lY5�o�s~���:�\n,O�@��ף(�����w���Z���X.��d7���zYC�da�  *,L����g���m��t���Vwe�0�>���l�~��{]�~p�ɽ@�1��0�"��}�����{{;F�{�q��[��c��sଝ�Cv�V�,g�U��*��|��fĂ����D�,� ���5a�U���e�=7���dؠ+|=Ո���y����	ƒ�6�F��ْ]7�����	,�*�|�wʎ����3&7�n"f=�KE�#�n�<�i1K�ܱݯ6gNJF�,5�_,�-�v�qrY̮��{O\RY�/7�-���w�sw��B��=���
�[�Wj�t�ޢgf�k b��.�v�]?�߯�
�_��悳-:f�[�3�J6`��t���,�]|�~Ц��a�rɎ���gqh�"�H#�TE\�X�N�J�>p�pjEsQE�%�J�4�˧��E#P���3�Ē���WT�s	M3��I,3��$�PU��<�UDnZx%QZsE���,W. �ۙ�P�E2AEi�YҺU��KZFt�6�\���*Pњ���-(�RF�č
��RC:�)2D3�N楖B*\���e��Y(�D��r�K�+���@]JYTi���ys��EHB�*��<�"�'�r#��Ud�J�-�"uDQ���P��	�Q��_�Nt�3
���xK2�ȹ��qĲ���<$����6"�Y��$
4�Q��E嘙Z��*fo.n(���)J2�2��%
.W=t"�"Pwy�%E��Q�RE&��-������*Q�#��Ej�ȃ$2B��
KCk+9Ei��-Mi!2�%ɩ�%]�1:�kduD�#�JK�np��DU�f� �W9ʂ,ڠI�g<��0���.���b1lDV��ǒR�O�)��v]L� w�s�@���gN��=W�Q���Q���]����-�k!D�H��+F��^�R^���;��7��gM�ˁ�	����E�U�\�OlC��!%\[7قl�vn\zN�]�|x���جdU`�vU����U�b����w �-q"��3����ʟ\�eӑۏ�0�7ܷǦ���S����+��{>yO�B�yU�7'��}���xP�ŭ��w+-Qg��v�4��h=�:�;n�z9T����T��,�G]�*���xK�߼K�]r�����	Υ�-_H;=�د����r�\u*C��z]����2̰j���_w�,��N� 3h(w�f뽷��n�����J��jz6����g��F�(�w�ez���5ު@&ko_^P��(��u{v&�m�=��~�~>H�L6���c]���C��/8���c�=��,�S�*�ǵ~�G�M-�d���Nw��i���(��F���C���6��eM��GK^��ۗ6$H�/�w��ΐ�a�-]Es�LN���z����x<=>t�r�ps�r�����ʪ�0�*�W )��>=�tq�i�d	K�{���p��2������߁c���=��Ww�9R�m� N\�x3|����^m7Q.��T���S�<E��޹�C̱�����_�P��p�����"i���`o9��O�G���
�g%�V�_��F��Q�U��EnT{ݛ>,��xT��seT)>���Oev}�b�7/)Z�[��Ʋ}:CfG��� �w�p%��A껅۰h����3��e�6Wl��^Գ^\�t*���h�fj_H�%U��>�+�~� �GJ�$gx���z!�����~ͽ����L�y2|c�R������'����d49)$��6GW+�󊢹j�p3힪�Ѿ��x;�88t��s���>r}���eS��x��8M9�,�K$��-[z�-x�69��/o�{�힌���dg�`N�Ti�q�՞��6�wt��U���K�
�1bWG��@�n$[�v���붲h��=2;ٓ3"2�*LGi�p�4�U� ����>���ί{�eL?x���9�+��}8���_eVԈc�@��^��/^��o�d���wQ1�CT���{'���Ϸ�A_m
f�t|�u\`#ݕw����FB7���e�C�
��W�f�Mǉa9ٖ�w�qҜ��Λ���`�yEK�2���n|/UQ���gxg��P����X��ޒ���F��^�������/�p*���Ee:� ��^�;��k��Q︊XF��{;��4=���K��YB���H��]�M4f�JF+�F;�A�* �]�1mP۽h��&��mX�v���<�$��Xg_-���T
ۏb���\75�ŏ{��3W�k�S����h2�ӊ�}�R����W��g��\�d�
�_�N����ܯx���ILTN<���6p�7��m�)��p=����͖k�g��KS�D�:�\mS�������R�mhyԍ^�nL�����ud��g�Ǹ����[��p�0y�ႃ�F����2����/E�%t�-�~�(z�\�j���L��N	�n��w��t��;�G�9F\��
uׅLo�[�����tDϱ����`�Y%Hs������*����*����8�wGAghU+�r��=r���Y3��y=���T:ީ�[�	�] rst7�Y��������h�?'JZ�q2z� '-{�_�G��z�u��
N��~u�*��1�A���ULL󺳎��z����y���@W����$wD�r����;����G�f���8X����&Ay����%63�v�e��hq���Tw<3dhϰ��vzr������]��޺f�s�G�{v�|y�ц��^�V�p˙����}��s̛ݜ��>��u���[Q�C8tj��x4����ȩ�3��j������_]��{����wG���NŔAOj�U�T�y��i����� !�S)����}��[֬�sň'p� �n^y<�:��Wh��z8mݚ$(���jz�����m��mT�D�(��@L�I�{%KUc�{���������t���9@;sq
�e׽�4�����}��v������@�L�&���*j}��T�a<P��W��֔y���^�Kp�ތ5��|����~'(���y3�ުv�C�-�rv<만x��*my{�\m��zU�����ڻ@Wz�H���h\G�j{�l7qLX���ꉋ�W�RGmn��S�w���l�M�q�(���tW\�.�{�Wxo����wŹR���z����r=��*�q�yN�d�������Hl�eS�ș�Ձ[�;�dm���ɰ�1����z����z���Ճ\�Eqݛ�Ύ~�ۑ��������d��ɐ�z�}	5]�i�ͣ�.�/�����ҵ@.��)�����w��R:pN�j~�ýu����H��K�TUMT��yC�����e�w(��~w���G2@w>��	SS/�����UX�^T}V�Zw�8�f%)t���Ȕ@�8����F���Tз=����P�OR1��0�T�� ��(*8i�-7�k����L"bY�>���`���8�N�F+��l}�0Ⱥ�1|�٨d�=t�E&e��T�9�^'+P�;�DM��2�����$Ƕ�\{��<�`P�����DF.�����C����'�b�Y�a`�)U,(�4��KF��)�ݫ�F�A�6='����1���������A�7�hy�^ٕ��^gU����u@o:����+�L��g*0�AF�{Ч� >��G����5Q��O�0�;v�ʕ]��{j�y�o�s'V��μUE"g�9��$wO3�q�h�\�J9g��F���E*��wws���}=:�M�� �__DϺE%L���/&���9�I��v�� P>7@���{�"��uH����Ç�K8�l�I����6��ª�z���r}���%n�{�w�2��9_�V7o�n���>���U�"��H�(�pyS\H��<������g�m#�{=Q��W*k���Z�ue`���F<.�Cʭ���_��������¯@=�b�=Cs'�W��K�"�iTf��l����N�����*!��MyT�KL����>�z˼Y�{��l�N{mׅ���1�9�v����}q�"Y�tt��� %�3��׵��x�F�AN0-x���(r�F���]h�N�N��P�P_;�蕔\�d�ٝ2#m
�S������FS냨��=���L9�<�BP����g��rb����g�[�^+܀�[�7ڊ�a��:#�����M����ۖ�}{�]�o�f�'�W�痀��l�v���4d���Z�_��{,��T��/����x�h߬ƻ]iMΗ��xX���Ck�Ǵ�ߑs�.{V�޳9u$���v������[�
�ǹ�n�9��(vL��u-�v|AW[MZ��yi*K�9�F��Gx�R���R��A�.�ʎ�^O�,���(ݭϾ9=`lw>5[>��׊��t2�OD��;�w{�WU \lKsPz���T��{d_������Q"9x��뤲�_}�fpWۆ�ܲS�.�.-���s�j�a��f����b�q��Tm�3�}�����J��K���C��*�wN}�P�]D��;*t�m8���j����O{G��/��n�3Y=�'>��wL\"g���zj;��t;4%�F˦71�"m=�Mg������꭮�e�~p἖:I��o\u�)>r鞙|��U]0��|���z+���$�ς�N�(=����A^!��o�=w��v����I�0�A�J��+�4��^�з���wt���@�n$[�v���붲h^k�5�W��S�k���F���"�Q�҇P��\��Z�ۮ��4��͝@�W��9��4�צ�t�)�� �k۠i,gkjm��/����Xs[���.�927�cɏ��5��=����Wޱ���u�r�AҘ=�֍�)�����r�!��T�3�^Ve��t��V#M
<E�\��i}�4SD^�>����L u�0n�k��oo��y�^N��u�2�誏d����n��f����ɾ�z��y"+�h�3x���0\����CC�٤l噰�F)����Ȃ_�瞫�.S�����e�Ҿ�Xw���P��9�t���G4K���y}~�lz=�2&���nt���t�Y�*�z�<�to�I����Ψ�S�9�Od��+IW�@Wj����:��r�v������PsqU �U썧x��O�nR��p��0�߽wwOٝc�ڬQ���S�w'�uGl��,{�0[��¨�����T�|=>t��r�,�i]@������͝W]���[,{�;(���騾�pE�uq�~��<���Q]���Q�'��(M�;t^��E�J�8�ޝ�b�R:pN��� �=��H�~�n8<�a .ҽc�	���d�)o^��\��=3�f�g
�T�\(�� C�X�}tG���W/ϫV����~�0����v�q�����~b�6�o!�oTԮ�N�]@r�"$����h��������<p��'1�gjʇ/�e�S�`�7+�oi���zL� U�y
�8�y��MaeKK�/�5����R05h�kS��w�k\�k;���a�z�q��H� kN��}J��.	��9�u���n֙9,d����"=D���P��sL��.�n���c���\��~�.H���9�r���|j�'��kAٸ�:$�Sc�m
��WJU�5�����t2@�*Y����MZ��Y3DW"%��q�0����9:���g���:�	��N�ᇡ�� {���RT����^���^��Cc
�n8׶�?O�~���[z;�g�9�[���uNt��\ ʍts]%�zS�c�z#;&�[yS����8r��Pw�#P����ѱt�u�1h�Fw�V�h�K��ޓ�7���$p�<����.&W�٬�Cw_E��;�֎C��\�������<y�yU�b�O&}�Cw�v)O&H��E��4*Yڎ��|��;�����{⚸�wm�+8�.T:�0ϾWx}ާ�9��%��i�����Je�{U�r֭����ٳʣ�:^Y��2��X	�V ~ۦ���+������ {ӹ]���onk�M��6��yN�����s�Pu�Hl��v��C��LW	��!��GcF��<fcK9,�ë��	j�$�pu�t� 5�����z��y���A�h+r:D�ɗKL�{Q�۹@�^뚫0]���-���=�w�<���K��5�u�T����|h��[*W�u�T{BK�#���5����H)��;�vMǊ��Vsu�vo�Ύ~���4{��OI�u$$ugy��b��fN~�O�te��v��h��,ǟgj �r��x�������rU�|�ϳܘ3��5
�WeH�����i�gxD�ݿ���.�����6���*���̭H�QH|�G��{ٕ��s�ȭywU"���5K�lQ�n�M�<�l�K�T*w�;z�0��ނ��Rqj�w.���FHxz._M��\d��<�d���x7������3��|��5Qgُ�wi��I���F�T6B�eއ>�j9�hwq8���]�{��y�ާqR7_���k��-�=��&�2�b��p�L��=3��C�}��_,� �"Q�<�>���.+����g&jSY�:c���S}vB����H�T���3��W������߬�
�	Y�ݙ���J���n2z�J���N����{��S�O���=^�:�nnk��<j���sܶ.!�e��9@�n��ߍd�x��r<��#���	^����FuA�y�yC�Q]����N��7��૴X[�k{Yݔ=ti>�%�b���o|2ͦL]�IvebPR�������cǜ&v�Et��5�f�a�R6��N�v�xp�L촕 ���Q�9;�_��gc��BV���z���V�\��{ۜ����G�s،�u7��M�Ó-O��+���쇔�4�;'�����3�����ko]*�-��c��`��ǊJ�}ݶT��\��G�Y����hS��T̝�������zfcS��S�2p5�ڰ����i��e�������+��7�	r�Ժ���W۷~�~7[W��k���@tB̮��������<�p��<<	|���%O{�ۨ��]�ˁ�k����{���T������>'����cZ�JW�/g�����h�]��]�c��)Wh���i�d���0u����٩�.Ұ�:���߻
�k�$?�<�fd��J���u�C��S7?�'O�_�22:�N�G=�a���e�Q��^�@c�����,F���� ��`�%V�EN�l�~�\MC�TKS�q��o�.F
��Y�h�<B�u�����ھ�B�#2���T���S�'�J׳�t�~�7]�L�^��0�=;���[�D+��φ�ݦ0"%�|��M> .��T;�����}D}l�`Y2��Rٳ���Ц�T�a�P�� V��,���	�,��J�,!�:z��>ܲ�7��ӝ�-����`�>�,��g7���W��zJ�F��v�"�Jq�H)b�7B����.6��&$P�o#�QjPm�C�{6on\��L����n���4��p$�lJr�}K2�#�neٹ�_k�j�5�$��f)� H0�c/<���{7׏�x�8QL��w�]}z��2+S�F��T�!Š�O�.ܽ�/���([0����}нT˫|Z���{%�>�C�c5��BNCW�x�X�����r]�I�x}һfF��a
�&�p���=�����º��>G7^H�/ZcCAw�,aqܢ�N�i� �r�ͤ.��]�a�1Kh��{N><��=�ˏ�Sq�����ds�c�L�-��5ԍ�ƻWK�wϯM�^�6V{2��/:�űא���X���͜eban}��s�O}����t�4u�%��\�.�ԯF�r�������ǔD*_��b��4�vc��Z�����vP��b�Z����:*=���ұe��\���`[�ǣs�ي��Y�0z�.����7��T*�xă ��ﲛ��wbY�%^�8)f��¡��d��ե�K�gJ&�J��G�����/�4/=�k����}:�m�w)��O�zKp�o�q"�w�ٝ���{
d� �u��u��Q[V#��0�$��'�&����;���0��u����Y2���f�ѻ��pA�HY�5��c׷������Y"ɛ�_�#&������z���d���H���]]�/X��^��fS��{�.m]�	*�*v��*�n�e�l�;##).:U��Y�J����%t��|����;��Z��������(R�ٴ�9���2�ns�3Q�r�Wx��4%�v�fR�/�"��R���ݏ�G�0<�Ӻ�3�M�E�2�J�/b�vK�ۮ���;��dr8_&&3�����z�]Ƕ�>A�ؓ��5c{*��ٹ4z1_e�lN�\�Z�CC��Ge��:�N_<���k��}�tQ��{N��pbNJ�,_$���r{���+�^���E֠аd�ڌ����~(KI�_�0���:_��&�q��5Y�P������3�mP=�y�z���0,��YE8g�,{�]�Ag
]'�w��hl�<J���'�F2�N���:r���qgL��<Z��!�Bc��V>�w�";F�*k�-.���B�)A�){�s�"$�<y��#�@ŃOr��֊WS�rz��>��s�牙(!��%^�L�P��s�����IJ�p���ǘ��o��l	:��ԥ����sփ�n�UD�]@ַhe��X|&ӝ�I��T���kw�*$�I�{/��
7�YG0����R�pv�\[�sh2��&U�\�����[�6�
�j��oc�	��ɵ��%�.N#s�3��G.����ʍ�9*��XXY���yiG/UQ�����@�%+RkdJ��ei��Q
f(�8J�!`T�<�!8r���eUuTDG%JL���[*�.EqyK�Y�*e�9ǆⓔV�e�8�<��9�-��e�YDU*��*f*�TȄ���E�J�dQE��/
af;^E���4Õȳ�1=��ý��Ƞ�s�C�8�EY]DY�$��bШ��$���őK�B9��(��в�MC��J�"BN$�p�2�At�:�j�d|�����(�r���f�U�4=Ns���{Ȗ��¢*�����4�M�D��8A��P<dUG'+	[Yْʣ��&I|��I�pE�W2A*Y������nZUr9��UT<q��B���TId�U
�2+"�H�.Y�D#"��&�h%]n	:�!b�*E���ثo]��}���z�k��u�.G�EGheޓY� ��4��|�S;l]��OW@�F�`P�n��뛰B�Ա��`RM�����`;�ڒ��ɬ��&����+�b�UOM�H���s'�>]�Ɖ=��tmRt�7���xB'���;M��:ջ�-Z�0�~):�����R|�	pA����6ҕV���'E5��ę���C,���7��&���e��i0��T��S7�ڱZ�������c��g���Cc���zun�_�l��h�~i[$��U�x�,�՗�e#!{� N끸G�Uƺ���oo����`���}镽w��_�'X�Ǘ
9n	��e�
��tk��� 'm�o��G�yC�z5��������|º�����M�Q��^r�w��[�����4�o��]>�Xw��B��nx_RW��
��V�tU�����O`�F�H�|i������p1�c�~����k��O�ٷ�ѭ�g2�� ӥ�t�����Mo�z
ʷ;���{�P	��#*6��/�)�n<[�~6;�pL�:�ѿd˛ �.\֬�칎�-��엒������2b[�U ��u��_���P/�y��(dmdn��:n��a5%���t��k�o�J�h܅=�޹0w�[�S�@�ۄ���ޙ��5�����W���n��o��U�k�c�}n��󛫞[�ox�q�KԱ��b�z����~�:��r���4�4�O8���4��u�'wdI��k�����T��^΋\vQ�2U��A�>�wf+��o��h�@��yO,/�ij
m{��pR
��>)O�gKZwe�������;m� �=��H��f�\s�̩�ogR�
*�h��vL�~5����ҿDL�3��?MFp<)a�7��>�< U�s�
�\�.�O�f��n�b.���9Q�	���@ޯyx���/'�}2�(��﷪jjO�d�>˗P�2p�dVSZ����M���FM�*(\U�s>���۹D�,d�_d���P��9���moUM���Ozp�lL�z<���,�~�ʋ�/�A��g���5Y�ވ�������$��Z�t�%��s�gk���^��ڀ���4:�v{�/�Y3DTG"%�=���r���ߗ=Gz</�P:��	�	��\�҆�(�i����.r?oߞ������g��@���B~c]#�!��ϙ��WwͻU�\�g_\/}2�M�q:����� �'^�#�V�����ɭQCU��r����ҧ:2�K.�G����E_eV���'+I���\�<<���By�)�=�y���J�V$�8�՘,��l��n�^�~ÉF���ӣqEf��e0��7p1���@,^�{4���9��$���Bg.!CN�|�8 ����T�Zgn��O|�SK(��8S@�EO[����?��U��4�����S�v����Rr|<%lu�_<y规���<��!�λS���p!�9�<�K�ZH�g�>)Te�첥�:�S�l�ʪ�
;��E��sB��-OP[��h����Ʋy{�﶐��ΖO�e��@YE�o�����e�}
� ��<�0��J�\z���tz;��}�$���{+Ü��1>u�9���n���Ќu������������ؽ�{��3[w�՚�xt:Y`_��JO�������7	���m��W��}\nh�Z��*���\�}
��8G�SK^oG�H���i��4�|�f����M����'h'r8=�gv�{{�%���q���Ջ����E�:X�8�e=�����@�r9��2�5�Q�r�L�����o'n���d��֝���|�t���z�S�WT�*�jn#����۠7�u�F}}X3�X��{��f��s��t:+����%��O@��>�.���EN��z:˹�Mw�-�	�*Wy{x��r����EW|�V��B�P�B�hw1u g��3Ds�����F�GwT�q��򍓦�פ�b���vQ��hM�:܊op���c���&���5Rzua5sI�N�~�]���: `\�:�ms��F�:���:U����J%�.:67e+}��ShL�z��E��[�u=�7�������й��H):{��I	�k�#J��2w�~M9�%�rz5�p�ᐮ녢eȧ��z�uP���b���
��7�5�J*�<]����i�����`���jo��+����'�!KӿGg��n��Z��?Zc���k׳����.��y���d/N�{R=}�����7,���d��H������V}R��=�7e���+��ݓ����`h��yW�]���dc7�Gf7ST���y�:n�U!��:}u�#B�;�P�ѽ�*n�jn��ǀ���B1���+�޲Z�/�s�����|H{qHX��T��y�Ҹ���0�yE۟�,�]��e]u�(�qlf����[jWb�������XOM��q��c=���oC����wP�G����"[�8� �^Me�X	>���K�,��e:���S�<�Z+�t����|�|>Uj�{�ןk�\vW}�G#<�`4r"���������n#�F�f5���F���;/H:Ę�'3�����)\���~[ylzVWT�d���9�G]Pˍ�x=�>r���"��P����L֓���N�sߺ/'��- �<�Z8Z�/��gR�|-PS�H�3V��[�!C�|�Ղ��J���"ᛦJ���]��b\<�uZ�tdz?�����^�z��p��u�ً'u&p�N]os���p��AGp������'��c+wO�C@1�X���S��2��yu��eׅ?U:�=�9�0P{�@{#�׃��O�!�u�=}(���ښ�8�s�]q���ڑ�%�=8Z�w��z&)���Ajn#�����`���{&/U�W{<��
��r�R�����$���(��� �]5C�y��ǺP��Tf�}�f�[���љ�&j=/'���c"X��u� .ߥU��>�ڏLn���q=엺���	�9�d���'ި�̢eFKɓYP�UQc�"g��=,�k�a~�T����J���w���_˽4A�n�KNW��x8���#%��p0=������awR����P���	_f��詸�P�ޫ�(��P
p{o�x�{g��q����pW�k��o��Q�t�T��0:yǶ�unv{�.9�M����͈�`z����\���1ZX��-���y�m���� �?_�=�W�u���W*b���{>���L����^���Pww&�}�^tN�G�}t7	ڝ�Ȁ���_��b�5L�{'�9�/;&�k���+��O���mC>�G�!�򣮮"ť9b�������������(s������n���k��MA���L����[��P6a��u�y�*tw�����0q����㎅4�m��xg��
����"]xS��<�V3�&.0�ۋM�z��I%����Q��~Uq�v?\S��R��<O��Xw��/����M��>���&�Dnb�)%x�B�v�����nN���g ���@y�u;�!�>��� �����o(�ܵ���M�{=��4{��Ĺ��@;�����]���w����³�����D�4_��~ ��ͽs{k�Wý&{��q�fx/]E7>�Y���t��O'�`�݂㗦�]^�����7�|�t���'�p^���� v�[���~<���
M>+ /s$U���w���K/�����s��N�g)��T3�&�$tGw���f^`�}�F��Db��{xf��@�G�&=v��}��P?MFp<*!a�7�T� (Ggfd����E#���^z��'�qY�.��qM�������G04<��Ck��?`�=��כ�(>or�Jy֫y����yЙџM�=�]`��2�ɨE�ɚ�c�	n���o��+�.��<jWa�ڕ��tY3�*3`ʚ���w�?P߮��.�9�ÿ�4�^�~��vF��U�=א{�?-�%+�}�5A�Ѿ�<�1��7�V	��V�ƹ���UV� ���Ue	��)�_�Ng�<�i��(�ײ�>��Y{BL}\�y�*3't"뇷�8�ry/�����I�e��ץ�����b���/ި�_�yf{v��K:B��B�P)��5�hu.�،��zfȿ��#�{n;��^��9mߖz0�V��׷o��g}�G&�4��K!roz�.g���T��׽5�;��W:}&��f���*�js��7/r���fR��� g^� 3Yɛ�7�J��êU%c�W���*�8�{u��bݙ��B�,�EN��^�*���8�&xy�� a2��f��a]ǳ��y�8�R[�'<�W)�����*\�C���W�� ��<�U�ʭ�=I϶Hn�X����8*_cC���R�.5x��f��Yr����:�0ϣ�w�Tw�䋈yX懍lOG|F�u9ei�yfV�S�M�Gz�Kd_w^���/&_*���UK�ێ讹�U ��� ���-���=U����PL����MǊ�W�c��&tV3�9ﰱ��wގ�Y.���>|&6����/յUW~|�{�1�e��ǼyI�x��*��)���`������"7�1�-v��g�;$�F����42������g��|W�j��Ss���c�oj���z��$�go�Vc|`93�M�6�������׉�퍶qx�S�t}8�H�#��IF����zr�|Ǻ{����Mس����$�jc�G;���L��{gXaӼMg�{;7��Jڛ��Zңs��\� ��}��W|�IR�_Dgz�Tw���[t:X�0S��۷�_���+�ca��6��{_���վ��ɚ�o��k:x�{���~Y��~h��;�r*���YtSq�];�t׼��{'/�Q�1�86���w��,�����1�ô�\K!q�=���\�@�*)�����:��縲i�C�׆�5x4�{���^8_�He#S,RU=q~�d���[p}s4G9��F�={�O�z���5��n�g�I�ɇ�[�vo��N8g��Z&\�g�z���wO��U���"8=ˋ��~�#�=y�x�����~acLש����y�M�������t�J�=7��Kzhx�x�%~�jz��YDz᪐�nڑ���w���G'�v#e�ʄ���T�o\�E��9�{KuR�����7}LU�a�y�� ��\��-o�z`�U�����#̪�l��⏰K[��U/�xwQ"�Пe��Yr���+�y�	W�rC�~�yf;�ΦT�R[�3ܪz+�{Iok����0m�|l��7϶ʘ]�K�fԢ��=Zb�7�v�����=�]�c��"����ւ�x{���p�[�ҷht�p�z��y�p�"�!����1��Pw�g�#ӽ�`���X��6(�3D�´x��y��\1�L!�-$�����`�+veZ����=w��)��D k�bIv��rh\nUuM��z6�77��b��Lg��:t1����G6��o�E�t�#n*�j����X�1p2�-�S���S��q��W؝p[�H`u7��^ߨ�bo�[X�bM��I¸�]��T��9��% ���=����/ާ�n<a�n=f5��Jw3a&!���O�x����N�\&�E��_}(�q�@7>��nv�ꂸ��x=��(��D>��Ba�l��m^L�[Y��?>������*�ͩ{2����w�\��]J`���.�ʎ�^f�ġe
�27;1l�`}XU�e`�')���zt�͞�{���ʺ��D�5�)G���MGMw��C+��vL��ץ���׎����rXzg�D,4��\l��+��z �w�p/���,�>�^���MT{s"
��q��&|;'�b6��P�+��j_H�%U�Ts�mw��k�uƬ�kGx[�"��X�P���T=�ݲK����{�}#��b	�u�2D&㧬{�J��.zUh�|;�b㗦�5�t�d�p�W��M�r#%�ɚ��}�(��lvlnW�PO�gԽX��^�rV��Q-��� ^X���޵{��FS[]��l�v��1��9�6OJ��X)�f{8z�#<�-�N��X�E�K'n��ݝF&��{��O0��s�!���ǫz<7�g��X�Z󲢼��v�ΰ6��Ϻ��r���\��p��E��q<C�~�I��(����k�h����;�
t�3��x{݊�4��um��=��Ҹ.��ϡ?�E��K�Һ5�̓ u�p!"��C��.0Ux���A��ʵ�g ^.�����ڎʍ� 0��p�d������͘��Sٺ���F(���U
�ū�k�O̚mFw/�1�R�]�3r�[5'��E�L�˸}Hh�B�|�
�g#ٝ�f�h��j<fÕ�W|�碭ᨫ��\��	DoU�\S���*�����^"f��PU6V���N�wa.u}�R)���7���]瞁q+	s�b+.�(����ތ/�V�R=��ej�`�/��&
��s�����������&��^.����;��\���p��b��|�k�4�iُ&{'��S�P�i����
Sq�h���n
Qu�w����ZAqɇxp�NU����+�tz6w����u�Ԯ��7�0a�j��MY�����$ߒY����x\m,�T{��~�f�z��a��^�>>��lcm��lcm��cm�m��cm�m���1��lcm��lcm����1��lcm�퍶1�������1�clc��m���cm�m���1��lm������co�cm�m����������lcm�[lcm�cm�m��b��L����H�� � ���fO� ď���_I���ٵ��+&"z��IL�5���lf�L�aU��lK)V����VKLIk+bm��MH��cQkZ�XS3ITn����N�ʋ4Z�k����q���^�^+ֳw\����in�wwYww��;���jų�!K��֢S�U����ص�mviJ�ٻmwv�QU]�{w�{ރ�},�3f��ggY�4v�E���ٹ�w�n썍M��N�Y�e2��h�gt�֦65���fђgW3�5%�����Twr�����ι�9,m���ݻ�����    ���Y�����y�"����.����m޲;f�n�k������ޫ���FSݛ��@-��v�.�v�n���yU���G��mz�=��X�h�m��oV�   z�^�UU�z��-m�b����EE@�^��F��GE]  :zǣ@ ����  � ϫ�x��ѣ��:�F���O��w}V�l�������,KX�VH��3Ym�  w��c�n��/{���N��m�gum�vڱ���x�z���V�y{�T�h�yv罆��[���[��6���޳��z���aw���ԩ�j�7T57۽���^����m��W@�LG|  ���n��n꯶9��ڌos$�h�Z���7q�v��<��qu[�W���v{��;���t3e\w���j���Us�t����{�s����7sz��Vedek�vЙ�c]ͺ��_  ��}�Өi���z<��jgT���u�v��h����Һ�^���N�d��O*���{���z�n��N��6����޵��B��w;����{�b�l�阴����v۩ml�6Z��  .������;!�Ҏ�]����N������s�M=,7m��N�X��{��:m�۰�L�t�{j��.�[wa��g!�o{����hq7.�ֹSn���#[�%%�٪��U�]��  �π���m�K�w�+�՜ޖk�����w;ݛ���m�v52��:nƑ���:i�9N����R��ݽ5��J�����g���3-�u����X�n���u�ک��]��U���[lǷ\��  ����I����wm�-`;���m誢۽�woP=/Z��o{f�O$�����u]5�gw��A����L�ݽ���n��J۽�w���N��{.��jOek�lҭ�wz�Cl��SovE��_   ��}n�UwU��N�Pj���[��+��oU�޶t��t���yץ[tk�m�����];�)c���ww/y/v��Ww:�z���Z;�����6�j֯k^�ӶMm���L+��ۻd[�   㭅)�[,�f�]5��ۏOZͫ+�q���a�n�zP��ͯos��j�y9�G�r��y�qMW�6Umv띻�n�	�T��l�JT � Oh�JR�  S�<U" �S�A)U=OP��I�Ҫ���  	4�5<U"��G�~����~�����?��?�Ugؗ���ySeOS�Ͼ��߳��o_}��P$�	'�H@�Y@$$?�B��$�	'��$ I@$$9���]������֮ٙ�=�[ .J�^;����J�Vꂒ73g���M�ُ_�Ji�I,&<Rm� �b����3�)�˧!(I��Z(, �.�5:/`),@�5+#��Yf��@k��p馣:H8�y�+N��ClK.���Y�@��*i��W.o3\@�:Vfn I1x��5��kS�h��QњN�f��YQ:,Pe:�Ե�U2-�#�xJӧ��P�[6�&�'�F�M�O�K���Ĺ�B�Q/T[�y��Wi�[2�W�໕<1��fxx�j�v��)�tk"X<��~h�TF��j�q!�%��kn��8�	*�-8́�%`��r9t�S�h)�Q+�������KJ4h"����M�I��-ZxZE�-ط.I��kA���3s�7@��A^��K2��+j�M�j�i�c�E^]��+�z'�ה�����S>�lY�lO(�%�j�H�q�{�6`!X�2��M�zC��
���Y�5z9�R��`[�2�P$)ŭ(��6PN��U��H>�-
I�wpn�k1�m��qTQ�78.�1x)b���U���:vWd6�ti�C�`�t��1�P:��ϭ�g��ݥ@I���	v�3iRan���A"�}�Ch�*���J��^�ƴ�tV!��WF*��%�d@]EZU��Aͺq�f��tڂh KNK��恢���|ꄫ>�>��s�e:�㻈E$�fz``@Viǖ�Be�6~�m �A�����īv��ʲ�e�[-P��i��$�mç��ˣ7q�;�a/'�o,�k8�t�S=��߬SIW�Z�k�]h�^'C7n?R|�&jB�Jr�&	)�F�kw���A�a͖2�x�mta���|�x�b��F�-�85(�{!���W)Z�(�.��{]&U]7YF��29�8�v��֭���8��ebB�͓v���dݚ@ښ��vx���AN��煇�ĝbF����꼪M�ʴѦ��gv1 �X��R�I��F�˱v���Kfn�,T4�͐�"	D<[���Y��O�+m��^O-��ȫ2?m�d�FN^�x�+�e䍼���ۓ*�=e�{Yt��f��v�jf
y�C�CH��î��J{J���	���-�%!��aU���e��h;��zX��%�Y��۔V4����rP�[�&hD����?CT�[3rfU�S	w�K�Z(��Q�Z(\"5{�kVǂ�JZ��Ñ�Jt�
�CS>�KU ����~�di�m?nQ�2Ky�V�n�����*n�1����ɑy�P�M2(��3V�	�=�c�H�1!2{%G��QCW���ʓ*-v�m�U��;ʕp�|�򌣲��h��y�V�:Y��t�����U@��o��#5��c��b�wk���t�o��$KRʈ�A/ep�߸a^����^y��Ҥ��� _I��0��0�/o��*��/k.CW,�#�@M�������g��]37/��Q}�&ܯNV�'���a��Ɗy����w��!Ra�k�%˄�dG�dN?6	0!�b������>�J"D��������|7��k�47H��r�
�2��l�D*^�!�U�~#K���F�u,К�֒.͋hn�d�S��I\�Ā�������'c�����X�R��[���\�P��N�U�4�?q�C�z���V��$�Yh%�3��.�E.ZZ#�ɘ�fX�$��+l��;EI��3r�J��xw�ͽR碪	�Z!����6F+���!�c*I�n��V�wAYJ����n��v���л��0����Eku5�5���kp��3���F�5q�o�n:�D�X%"(�p�����KCUjƄ�-ƞ�ZQ7�>��)����>P�a�"Rɡ�TVk�Zv�{m`�ڹU�F�Ch���D�`��0�S�e���0�@ؒ�N7��5|N�$���}�6��ӛ�q/[�F1pIoQ	�څb;b+���l��87F� ���6*4��ũ�t�Wo69ُ
�MIZP*��~��02|�c5\{�6/�h>n�6��-)�ij�����#O6�����8ىt�%�u{��T�w,������@|��n1��da7n�o嬈�h6��5�]Ӷ,�;#t�Ǫ�}��yv������*5bE�j����e��KMc�	apT�J��3n��z>�v�ͷ)����h^��S-��&_���ET�o�'��Y��e�V��'E��|���|@W#̀�&8hQ隞�6M�+i�17�{�l�B���n^^��n������R˵���'�������j/R�S}hP[{�1���;Z �My�^�qX(���l#����LPE��m],�!�؃�\0 ��H�k�o����=�S��>���IR}�\-��|k"
�~�u+Je2H
��ͫb��zej�C^���$d:l	�Qf���4��u�g)�z�3%hO$ӏ&�0Ta�*ts0�����3C-k�����^,��ҙ�7�.V7�wT�4n��ٮ1�|3%�Xž�N���lp�b��w)V���߇�.+DՊ�k�e�?�XX��[��-�A�d������Vj}��Vb�YI0r�����㣚��)�S�=�3����@���.��S��
��F��t���lR�X(�[��i�V�F�Fk���+%�ҔP��,��7uR�������c�d��q�1:�S`ԁ
���-6V�Ctr�!tT�3m8M�m��)_�w��V��Ǜ��̻OF����[q��мp�x�hئ�p�lJ�"�̳S�84@)��F�]b+C�^ټ��͙(��[4�c���b�-Lt�b���eձf�l�jk�Cu��0�9[�+wYF�k�6�-�(��Շ`�8�`�n��E��&�j�p�M�,lSS)�q0n��\���ʻmk.�ܺ�!�O�j��H��/?�!�4�������T�J�;\X#�5i�hd�e4���kL�֣��nt�m�S;el��d���I�6hd}v1�M)!����&���.<��37V�EzF+���	T &L�޽"�:�H�b�:(��z��V�!3�ӣv��bL=(�^�A�@D[Q)�s#0�6�P�ܵ��[%ǲkDm�A��9&�U�I�-�)���*���.R���� Gh7� ʄ����p�&hB?�-Y|n�f�%��:��35L-�wM�F�*�m'�%�����x�Z��:�|������c�ԛl�1ؚ�n�9�B�ݒ��(!�
cU�r��~�i
�4R�fE�Ix!����Ym�CJ��)�r��[Sw�E��[B�h��*AyVڡ�r��\!�2���0�]��
vg٤�� 8��)brb�w1[���ݚɹ1V��HSQ�N��{�'l4�1��(Cp�N�?�'W��8�*�3s`b�l`���i��!bii��t����o����KG���Y�.�3z�oN�� �V�ft�4V���E��ġ(ߕZ~�C�m���~هQ�*���b>>���� Z��w�2��E��vl�4�&N�gɴ	"��ލDU�7Cʃ��Py��E��hɳbV��ɹ�Y��Q�ja�x�\#�0�ŉ�����ыa~��$��iS[��A+��5N�	N�GK�E	G%������M����x��(��
�(MOuK9��ԁX��MA�H�T�حk-u���+d7�Ak ��r�&���F���5�<�Jf�X��Y6�� ��%���O h�� R伥f:˕��j���+-Ǳl�Y�AV�*�U�V�.�1�ɣA�p��$��f�f߭ L�y�*����Lm�E^��b�1[�J�7)�nn��a4�fʙ�X~ �!�ŕ�.p�e8��Z�u�Q�/&�A^���&3Vk��Q[����sAs�[�������S�d�����ʦ��g�����5k�S̕y5F�Y�e�z�J�XTc�l)w��bXPWG�2��v*8Mal�Z�2��{{eU���<�vܴ��"���S�����0�) �|
:Vk����!�S��
-:�/>#G�����!{B3jz^I�n����'5B�ܺ�c^���aL��B$�Z���)�^Gf<�ɳ
.n]�7Q�#gU��D�z�j.��wR!U�#h)����HS�!F�SH*��Q�Q�Y��Y,�B�Ҏ��B]\/[��Q�o�2�-�%�AV�Ǽ��#+���Y�vU�U��ud�ZƶJ���1��d��[p)A��wY���ҙT�oX�K�,ѐ����L �S'�z[�it ��J�f޽���p	:ɼ�@�0��{f�~�F
Z�#�vR�w-�_�:�F�W
�m����m��Y	JOẓ5�OՐ�J��@�$ F}��6K;M�<�z�$>.jsB{���)L���xdS��Y7Z�{K~ ?l�n���7��?�m��g����i�[&m��E�l��P[+hb��D-`�hY�U&ZV�U�wr�7.��۴�JR4vh�ݫ�SF���Y�'�yxk����C�Y�i��&\َ�"�L��UBm�IKAi�Si�@������X�]˔b@,0R�ZŚ�K���
�<+H1M�͘ )���v�6Ӟ�! �T9l�I�!��eǢ�%��m���f1��$5�_�Kdk��/V��� iH坉[hB��DoEհjkA��UZJ��n��,�[%����"ɘX�GaG�ui 4��	�u��-8�!GiCyn�����70ψx�V8�@!Q�|�۰�e���C�/�/V�0av�^7X����W�VVn�J2�Y�iذC�T'Ddunn���h!yR�̚�C�ȨMcV6��T<:�}3�P��5ߑ�y����X~������D��k'�^���GD��zQ������t����j>Z�
K#` �-Qnމ��F�빥[F=`�X�+�֯���O7	��)�z8�	���4"z��uK*e�"��ƴ\����lt9�Zm��A���q���0�75d9�{�b��	�2��W�V�Bԃnm�8�Ti�#>�	�+r�ʑ��M1�!��7n=4����F���^{o��ė�U���v�� �̑%�t0�D-b�*8����2�|ȟ�7Cc� ���0ދ�kf���-�jT�c{Rƭ2����­k���k�B���J,xN��+��!������Ym!=�_���=�#��	Lh�}tᐫ��
Da�<7'���t��聖���nK#
&�D<����-�>����Ғ�&�&���*��4�	@��JK�Q��Đ��)�}�ǐlKZ�����a]
É�����(ٺJհ��Z0x�b��y^T��%�g|��j�p���*�	�r ��]�"\ll��]�P2��TF�%O@"��+�DLÓȉb'��J��pŨ��J��XATD�z�dKe���:T�E�Ғ|�.��x`4��8�B CorФ�.�t�F�$Z��bK��5�� N�n�qb���"�vʲ��6�VyDk!�7<t\l�K��z���6�.�uC�"�7� R��V�Ә�3eUef8C-�����o�	��R\݊� �̞я��,�v����iړ����P�m��j*�5�mX�I���*�,��K��mb0��u4�mCZ�)Xb�&��~�o��Uu)~���a�rX(�]�r�Ae��`�*�$�!lm&X#��V|]Oz�c��ɒ*%�� �ؽ���VezN��
b�wp<�z�	Æ��c�����E-�!n��
��:���f��^��j�ư�q۹�r����~�V�@L[��ݒ:ۋ*C�V�0���琪�
K�Q���t\ܻt�De�����3}Y�2j�}�fŁ+AO�h���A�Nٞ���<�b�R;Q��)�0��\ӗX���d&�m�%�1Ci#�=b�-(�*�7�bR�KD
3pͬ%��7(���'P��P�r��GsZ��n3�6���vsp�lυ eԌ#mϪ�k.Ѻ�	��]n'�36�*}t*$N���[-R�Te�e��;-o�`*��u��,<N� T�Xhzp3����<8b3O����S��}�d����/�D����[E
j
݃	��*3w�#V�,�*S���8B�e]�3u 72�Xvҧ�j�fC1$bF7��	�p�m�����a4�A��EA��BwX��,JS�-�ͣZUj�xUn�j��!,��u�m�vpa����%��]v>R���)�m7V�śv�!xuSX6�+DTsr ��a�Ɇ��S�Mb[OL��L��]���EL�8nIAY'&����bt��X;K�mHP�œ5�o]�j�-����!=DWsVh׮w�U�5��d���ɉ��c�,ԕ{�R�Q6m�{>_EA\-�K!h�.XFUh��;t���V�YWXh��h�Ԥwu1!6�/r�D�	U)�����`��A�T�Tz7m�k~� ,]z�Ns^,\��-� qh)`�ei���aP�*cI9����
/*�JC�&�Vv�ٗ+M�&�cA�M�w�SǕd�Ą��k&�Ӥ����)��ͻ2�j��b�͔تM�_me#�+����%��^���7F������-+�WŁ����S,�W���VS>:�a3qP\퇫x,�ŗ���/dO�웣+q?���Ɂ�k���[��>��ѝ��޵����zV��M�ݒvH ��
�n������a���7���⯯%�"]�92����B^���(�9>`��;w�"�湿Gd)̙��؂[� ���'���Ms4�s���:����΂��ǧV<T3X�kL����`����M-#(Q����C�ZS�������|*�ʳ�15��%�
�'�>9L�u�A��ס�)�՚��Q�1XR��z�f��������q���jү����l�^��R�1Y�F�n��C�Pe*�\���k�TҭWY.�q����9FU�]��r"eYZ�#�n������u7�,g��DE�ް��nV�Qޘ��ѧӟ*�)���v�����E�×�޷����P�M�w�[މ�,�bY�34� P���%N��2"���=�H̘��:_nO��ؒ�����2��Z�&y���T5%��>��ɵ�W"DSt7t��Ρ�S7��G4���G�(tk6�\�O,�~��(�w�3h��ɝms��U����&����L])z)�7[�ו%u
&�\�x�˸wY���x��aCpq�=�Jȴ�/��b��B`GK�n��kG�qr����`WK��p"�	�ԃ���hv:�yjL��� v<v"���t��L��kO/sW���!�۩����᩺�6��_e>��!21l�j^S�=����@��vWTcj��nVV.�1�4�7���j!����Y;4Wy`�9�d\[6e�2�.|=/u����壥(��|���ȡY������:�i�9a&DB�cW1X1�)�u�Ѽ}�N,�/w�"t<P}��#e��&���׽�.��#mq�����x�+ڻ��K>}�&��]rE,RӰ� �^QD��i���W6��{%��V���"x83��+=���E0
4�;+]0�mR4��.'�v]�s��D3*����(��Ӽ���q��ץ}�.�T�uuX;���4�I�S��&�M�̢V/�ٌ���J+U$tS��H��/h:ïس��&.˩\�3a�%m|kd���0].Ё��'_���t�ORl��g>6� r��1&L[�gR&��lzv��E��dܴa�� ��h�O�[F���l�Ѽ�ln[t]#j���a�!���Y�C3՘��3y	]�-��{�P�q�7YM�"%��fs�h;��I�Z�����N�f���y�ӛ���~!}ˏk��=�wur\8����slˬ�����1��b�T��~�t�Ɓ@{��Fv^s�Nf�\>�F�w-9ٗ�fr�[(���s�Ѯ�K�����,˞i����<�,֔���i�u�X�LZs���ZB��y�y��ifEWHkr(�@�M�Rk
q��׍��յ�v���|}�����{-��5�0�)�-���Y3��x�����uJ��7��ݏy�K�:�-J�!�<�^�˲��Ҿ�N&��q{��͊`'�a;������p�#�@-v�VE�	ʝ[�&]�g:t��4��)�C�G�;u����̛�:x�X=h�3RǭX<���϶�Ir��0�9N`�c�*�=���;����X��o[�p��D��;E�V�;������e�3��\���4�)�9Z�-��)
� �h��}�vl��;�rg�뢃E�t;�<��l/��R,�
���GuԔ�u>x��Cp�X��%]���5%:-.���C^{[2%���d�>=��5K�hm�kNh���n�� ΠY�f���&�*խ�����L��7 g8M�a�C��3Y+2���X->�; ˬ�:�����foЕ��=S�r���1Y`�"S�.F�̵6�_Y`$�W�S@�r��=o�c:�wN~!nw9:7rIU/����L�	��۹vdgAt�;b�$kMp�i�}�@�Շ��(�a�.]ۇV��2��u�����>�B�F9tn!g�� l������G�=��/g=��#�ٷ�aP!K1U��}@�ܭ�K�@�����E�M5��L��p��s�ݿ*Njb�.�J�����h�tVX@�G���۠���:l}yI�M�J;���'̥��"`ǳ�njX7f�f�\JW{��53V�}r�sTNGX������񚆸����ע��GkX�^��2�T�YD�((G{
ݜ�lӕ"����ڷ������Q}¦t֞�Y`�����H'f��ϡu<���	�(H���;���V 3�];E拺�J����o�MUz��*�8W�-�M(-��_B�+n�`Έl�(��Mu�����3����{V;GqK��"�5�dn�<�8��}P��zA(�*$M�ۦ�Wu(�d�Ghy@sJqK�vv��+IX���.���j2��_:���dͮQmǳQ�tb��]�@ԥ]zL��iZ0��(�}n�o�t�8���O�w+�1f1!�nNjh����5<hq��Tۥ�ə�^]#\ ц3��`l�W�	�*�H9��V́R8o�����zL��v��k�#l\g!X�B�R
�n����m>�	�zO+�P܎@&�{#oF�׽����2�C�eM�aSK).�
��@�Qc�B��`���bFӭ%�L� ��@�l<Y�k�MO -zM޴ɓ%"�/����x�T�[&r��=y0�G¹�:�)�Kְ���Y�3D񪽻f��T�⽺P���7�m*�#���nx�y��e�#\D��[��R����\Q��5�������AA�y�9L��6E�c�-	�.�Z��۽ ��tKve��<{�+��-���2�=",^�ᎁw{uK� ͥR|�4a�bJ�L��H�Z��3*C�H�����'�m����U�ח{��-wT�+F�E��K޳�Y�t�p�V��_��܂�Şѻ��8���u�u��<J#B�s�?@�ֶ4��$^���V�p�}�Q������&
C*vWSSeF}o&���W��z%�|���&;�������B������w��Ŭ��$ʺ;�`v��]	H�ÂBZYۓ�zsu�p[�R�R���'4(�~������������ʦ�[pw�ˁoO�;wD��D�3��^�&Od��w�|����B��5����Ư�f�s��f�Q
W����
���{'Q��N�]^E�dp�z!�=�:������xz^*�� ��i�g�j�^����{YN=^M�N�(���zTZ�2F�R�����n1�g��t�G�����[Qc���(_R�s+f;�x�2]�*�՞�T_�o�eܡS��aw�l�&j$���*��[ZJ)������X�"Kw������>�e�u�� �Ԙ�k����Ȟ��*f�^��]�[܂ѓ�\g���8�j��x���W���M��q�Մ�}�a��^�_D�-��A��j �o��Z�#[���20��u�V2�c��ԤK�87f�ۺi�=B�LL�!W��B�Ь��b.��W3p��\��c�Z;e2�j�V	c�U:�P9ѝ\�+v�ҝ��{,�=��TV7������讁���wA�73r��m�&�a�n
9� ��5�P�*ֆ?S�	�	��.X9����zg@+urh��z5��8z�}]|U�\�{�2�B�x��;�ص�p���a��]��gz��ʍ��R�Mu1tf�YJ�--��@�	ю^T�v�_c�S�n_T�}x�5E�^Nh+ԕ]���:ot��)������rj{�iQ�0�DJ�凬���lz��t(�uQ��6:w-���8K��t���oM�֘���>L�)}9������|�ɂ[�X����/�E�E��2�I�&f�.�uypu� Dq`����z�<�I-�f�=�t�e�����l-w��y��V����h1~g��@]*]�tj������ڒa������{k���6H����.�W���	9����vX}��@o���Wܶ�c<���n+0��et�`n��3��1��2:��-��TXk��ڴ�-�1dŒ��^�v.w��f/^����SJ�O,���tt�����8���ξ�y�eɋڡ����'�W�A�g�>Υ�g�ܽpz%&�ݽ�p(>�˸�9r�M��V��j�z��i�F�u�አY�p��&���)��{�Vu��y>�[�B_H�������7���p�r�s�Ö�W_]24�ސ2���Ҡ��lk�J37op�ƣ�k�����r���p\�m�Rf᧪����x��;z��Ӆ�A��-[�!�/lC�,]���I:��=�.�r`�8Ve�V�B!�8��e]���<�ݾ��ﰏ`�!��+��%�L����S<�>�7h�I��Ɂ�7�]<$�l_l���j��[{j-Q�<Pfz���zo�!����J֢u�:�G��}a��6?\�,+��[Z��E�w̬Aci��>�s
�`N+{eV���^+7��y����vM<f{_ݴ��*+Y��u�����1]��82�=�7�\�᭗�w4��:#��� �+�rF�b��]e�v�+J����^q��ʨ��8+LǛ*/�ve�:�u��F۝�_���E��h��1)L啌�������4��#��a��
hB��z��+y�BsIn[�_�fT�uԣ��ܭm����Z�a�_%<�/3�����5�?]�p':���,^02��6�a)�<`�	RK��o9��x�ķ�W�}��a 7,��7x��h�C���xWp;|���[�P+���F�]E�4��=R^�ѝVa��F%	S�kS�.��c�ө�{�����!�l޺Stk~n�W�J�)@[/���,L�8aX�o\��*ʺ1�[$��u~�:\=*�u,s��Se�gk�N�p륁�t�2'^�ް�N��L��n��
�~�rs�e�	�v w��Ӽ��=8���+Тl��ۑ�S�4��8��6�ӗ[�Br����˿Zҟw5�~ԫy,����y=��8i�a�+�~7���� 4�e!s���Ց��<�nP
�\MU7wG.ըo0B�ׂTŀ�U�p|U�^�{�=��qw j�z��T��z�"FŬqb�'{d'KFT1I:E�@V
��jé"���R�*��*J�ua�Jp��b f=���I�j(�R�v--��)[U%GAE�ygE[�"r��|�
��D�s��v��<%w%�N]����5�ցb{}�x�\V��x�8p{`�� �[����\��ٴ��s��6"�[��
ݍ��Vᬽh����:`	C�Q�8�s���GzP���X�th4�B6^�}6v��gn�I�#/C$�vk��A�$���L�^��N|��q�k��ׇ�k8MW�Tp�%�1��S�e,Z0,X��]�Z�XE��m��"1�#\�B��Ҙ
я��_�	�6=�y�� ���n-�B���yU����F<��0j�c��r$%�n�;�
8|��$ ̂.��;�P~��vk���@�nm�\qGʯ$��<EӰq4ylη@Mr�]�e"�-RA�v]��&�(�o�@��f��w�f?j9�Pՠxe-�<u��:�n�Zܔ���Z�R���d�T�P�[��堼Vzo �C�_�!|��wDF��xd�M�u� �tʖ
U.�А`��-��lq�>�et���t�-Z�����#Uս�b�^�0<����oiẀ��,�ζ,q�b<LT�@���0e�V2�����V�FF�\R��$w��; �'�$ǎa{ʞ��)\%���0�¥ �_b����)I��i�����L��g.���HZ��k˹�qq��P�&���E�6j��Kn\��Ġz:���+���j8t
Q�E��(^����s���M���Z�כ!q���t�-&�D�<��Q�!�/��@M��|Z��6��\��Yz�����❋�#�������+Egd���Z-y^���d��J��G���N��O��',��-��9�r��%�i��L�}{��3�@ܽɜ>����4�۩�㖧W=�;�'��t�p�z[��#���.�m �.���J�rKu�u��
���N�U���J��}��ek��\�)���b�i��+A�z�%y��Bz���e�BS+�Y����j}�3�:)*篳�	����ҟ^�����j�M%��ؑ\175�o�%�
o�yTڒ�`;��.��pf�A�g9k���4��Pqֶ�ޏ�� [�ly�Y�]vs�K{E�)q�R�:������R�h9������P1y��^v�j�-\��HqG8k�-�FR綇xjp��2�6+���ܭ��ʤD`d,=le��\�M&�e��>v�`��f�
��Γ�b�Y���H���g:�T�w���H	�����&�W�D���y9���{5a��S�帝��c�,b���Үx䖉����{p*�v�Y�r��vќ�y��dY���]9D�@�1�����8$S�i� ��m�@�g�͋{�����L_}h�6��	%ٕ�OH����2�#rlb�n�iQC�ip����ˆY���t�Jt]�HvOT�J���"�I#J2U��ئ\
)�aT�E%�I�fH�}=.\�ɒܛ�.zIGs�S�[S�D2).L%8��f܀��F�C�k�Q��v`�p�$�����@�{���! ���@�$�׷��5������Gv��=E'ayxt��2��j50s�ݴCX�xC�.C�{�8�L0Q赗�n��ft��aSk^o9���#�,����-y�(��A`���an������|Q�]G��w�Hw�siԬ6b�*c,wgƸW+L5юR�'��7*��6	V0"��t��QS��j9נ��oc R�=�(5�"`b�Y���t�0�]E|c��^B�����.r�m��㋆�4d�%��}����}	��t����T������9L����cM��T��``XO=ue@�ʔ���Ѧ_H36m 9k{�NG[kw�bs/A[����֩&-\�d�mbG��aԂ�:)�=�#&Hq�G��a�+̒yc����g�r��跪��º<6hЋ���{U���硩�\V�y ��#]�h��l=k���3!�M��H}��91֞�c`���ɜp�!��`�v�2�	�k�X}&>�Cu��q�����9[�r�Յ��:����,*kj��K�QG�U�Tp˙�\��S6+6��MINZ�n��<T���]��M�c����j����|���X��c�;�a5L�7b��w���.�5�F��.�������H��������Shêc��2�C[M�b� ���J-S�Z�r��PX�����Ì�5�.y/���l�/S�ř`����V'T��玦�3{xNw�o�*Vʺt�:�,��ͱ��*{w�ۮT��� �<�N]Y �R��6#k�sr��U���M�S�C�w 4��(U���g�[y��m�½]1^��=;��8ͺn�װ�KwFї<4Sj�eJŸ�db�0�ҹ`�����X=�����=������ٸJo�D��P|WM��-*�x�ˑ<Ԗ��3V���{/jq���xm$bԬTC�㌽��Ǧ�y�q;�c�Ag��H�y3��%L7��z��;L2��<�+f��PvoF��đ�?\9>�p�ϕ)�U�n��$_m<wE�r�u��6����KƝ���Hg5���ވ-�w���Kz��h֨6�K
���܅k����k����_	B�6>����	RV�St<J���<�^��M�7�+L�O���A���r�
VOHK��@v7:E��XeZ9ԣ�F\�؍u����B;�!R�7�]Ð�`Ƴ��FY`�ʴ�O�����S���&i��wtNρsTq1E�vvv��R:ҕ#y|Bj���n�8��uɳ{X�ײ!���X��7L�]a#h��qIq͝4*����2�\oW�Id�WZEw�;�j�� ��kI�T*��@�g�����+&]/jv�Lj[:�� �驽Ӳ8C��^�Zu]�84+�y�ɡ{����t�]g:R��iЃ��q6(��M����Ǌ�tFm��Ă|ֆ.���+m�\R,�5�w����u��Zulɨ��N�I�I7��E4]�QjyVwݽ��'�%��w}�}w�a�1Q��V�d,u���`�����Ng84J��d��o�V�6$PF��b�Tފ��+K{(2��v{��)��g(�+L��x�9�ƞᱍR�Ty1��՗!�=U+�ùNۉ��U��I;����X
7/�"�P���dQ�#D�'s�W�GE�49�ѝ*�mɥas.�wfÞ� 7�w1,�R�2Q|tM��'(>ء28�'z��\�nc�F稠V��jJ��	��C#�u&vխ"�!é�0��u����_��q�Yw{W�Z���԰F�W+6�d�ي��}j�
#�=�]��c��h�</l���MqƱ���F]��r`��-b�3��v{]�ښ�y�D�u3�$;ON��j�Z�4��Xy/�1�Gf-:���O��r��xX���9S�'C�ZH�NZe�X�J��R�tÝ]��b�o1�;���{wF�ʘ*�i�!��ti�,=������05wz&��d��$fl�ӏTC')�ù���ӂ��g��IKn��{�[��5�y��W�����~T�7EѶ\��x��z������>9R������U������1J{�WR�p!f��>�1�L�S�����û�Io��9��Sx{�ͩ�8t^��|Ͻ����UcSL1,�[CW3C.|�#7.3�*ݛL���!
��H�5[{o6`�4���%����<�>�Ә��>����<r�K��������Y^ʅ��	�rr�v�|@��]رS�O��q�//���3��O\�Ůd�;72_�<��/�T��K���A�"�����8V�γOn�J��띸Q2�/fA�H����"Z*7��f��U���J��`��E�v{V_v,o'���[�'uBu�ݚ��m-�������@��ny	�֧�/�;�:fw&��滂�P��J��sN�w�<=z˛�t��盢�GR�6"����sɊ,���o&�l��!c�U�
Mf3a�J�Ӕ�h���iw��+����̣����'�F�㔍���@�@E��;���r�e�RƜ�#zn���CN�(əg7��f�"�R�:��j�N�]a�"k�d3��mз\��Ai�����r�)��ޡ�tYL>�8w��WSj��E���ڜ��k\����W\l9Me�ș�$���-e�������������o(�ٕj��&��Kv��V �t�#lh���FpP ��J�b��w���&����#��>�j!8W-�{#%��Y��(:&��@iNdQiZv=I�Ŋ% �D�u���h�n�5u�=����0�ė`���.�� �U��A.�lL��:��C9���gM�H1���E �]7��3L4P°f\���= �����/��W;Z��P�T����emZ��mp�؇�h8��f[�@k6
kcZ���*b�/�nu�+|Af�����å���C�~%b�_�L�Y�	L��R�^��#P�#6�w0m��u����0v��ex]�C�d^�Qى����Պi�d��/ᶖWF�����2g_Y8��Gl��\S��V�╥��,�<w���h��d[�Iѭ*�Ty�w͒��a�5�ݤ$F�3 �/ q]])�U�"��;�wf�Iq7:��*�ݨU�.�/�@姖�VU���խ�^�*<]�tĀ�cU�.�c��gn�է,.�R-�o�OG�1�֣!����(f�l�Bɜ�&�w��a+(�G�$4�
��@z�w��l��9���	��ٞ�)�^TE��u1����Wo_�]��+�{Z߹B�~�XN�P=�����e̾j�N��|ha.��$X��}����:�+h��5"�VSs�C�����y�����q���p��V"I37`�5EN�9�ށy�xVtɖ���hj�t�M!�A�P�_ve7�T�5�Bp�`��6�@BSR�uz+��n�5�^^����cfp$�틮��LK��`دTޣ�L��Dzn!D�&-��)Q,)\ݵY�v�s�t�'RN-55����|S�-�au�!\+V��3��4N���Z�d�赑��F��[!lA���ŃY~DE�<C�ssM�E��6�u �b�Y�b֭��F1IJx����z4�);������cf�{�T޶�����wJY���P�}z�'b�fok���Uf��"c�G�"Jg5\��Q=:u�i=6r�8��Y+�:o���L;�:',�y�^�UԵ��eͼt��h�
w�+h��2�MJ8�dq-�� YT|�6kj�+{yW6&�5t��Q����D4&��'N�k9��c��F���*�D�z�K!�uR&e�F�<�ƾ-�r�a���K�=�Ƭv����%�ueqdހL&�v�)�89�D5�I�pT=+��m��@������UDE�a��XN�!���.�4V�j�EZ��G�8;$ʤ#3�8
]���%�mL}�����<�oU�׋R@�.�@��}���v!*��g�ެ7S��ܾ}�Ŏ�:�kZ��(70Gy�a�wm%X �����P�����u� �g�a�.�53�t%M��ʥ����b����T��UN{%��Ǘ�#Gi�����tR���������DgT��/C���^�A���ua���4.��W1vn���q��s�vGқ���!�5]<�a�🠭'�߶�]+J��{b��������
�˴��T:`�u�{�f����]<���?~=��IX7=���d�\�[Cy�8�K�i)�7(�������TYU�o�W��E fZ� �_l��a�OGU� ��s/n��*Wq����״7�[vS�M���dM�vp�U �e�����mD�P՛�q:i�ve;J�eW���G5��>�4m�!:�bCEX/JGEe�|�n4�p�!������4c^���W=�M�[�5�=�\��P[�,��9|�5c�\���R�U�[���a�
��D[�tRE�^�1�U[0lYѽ��>�Tc���~�/��Ysa��R�G*1��r�FBwj�)����0;�Z֭��s��������ιݩt-�S(1�R�}!zg^���U��)@��QʷLխ��B�����9��<p�v�
�U�⌖.���n]�f���t��Hxx���k���+-Yމp���\i��T�����J*e��BU���]�Ј[�ַ���k��ݕ��Z��Uٱ,p�G�]���	������B��U͌;���V.�cV¡N����Z��Xǳ��Uw-����5�#�Z�e��S�D�e	Rh]1�[���԰'���]���ƻ�"��-��F!9n�؎�-� ��N��A^����w�$�����f���E�w9��|o+��h�2��e�i�h��C�$ρ�~�Y�ʆ �-�J��6*�5loRő=��y��n	�&�.6b"��\��4�V��QPT��GQ����}�$�Ԁ�Fp���F\PX.��S��SI����рV	e�=N�_r�ݜ�]�n��:�"Z1��G������p���2���w�[GO^�r�2]��c���l7{"�{ۭ"�ށ��»szΥf��I��F�N�N���d� G�h��9.�fAI�Nl�V�f�7�:d��Юn�R$r��u<=roJ��
��=��ú��Rpʯܞ�� �F����K�tFtԶwN�f��E��z0�@��pdr������!�e�O3���9:ݭ�]�/+"��֞��9D��[���x4�[��Kx�"]��D�^�^���w�����n�Ս��u��A�'np�L�!h���eG
�ؗB)��(�,��&u�*�3��P�7po��f��r�۶�㓻�t	�a�:��}m:��z�Pf�$�e���	��D��ԝ�Y�F��ҳ��)�8+��*�&�@��3)��BЉ�J����d�ȉSRX�iݮ�D�:��{��$�Y�Z:�n�uK���IX��Q>�Ss�<�g�n^ˠI�[҉�q�΂�y5,P��B$�$��X�R��O6ֹ�X1j1ӂ�h��d�U��9����x0N:�k���������
��U���-��3�(U#f<��O�U�,cSӽ!Ż$�Zw5�5b��bu�����j�m�Jo�f*��u�/{���M}�Ӂ���P(�W[ ��M�TzJ }$��7�;�aBN�ͭ�A��7����� �K�����+�I�6��:���#G�Hv"���9��4H�'�v��LqTi1�ƍ�/u����ث���Rҩ�^�,9�P�yq����l�fv��Ѻ,YT2錀k8-�WA�I��v$=��Ct"d���I�xAX�c��[
�
�[��5��.�Ǝ3���Gr�al6��j���L֗N5�:���*��_�@v�IF��,dE�&�>7ހ�����j̶3bJ�'5τ:�icpw6��a*Z�c<���%.��ʹ++`,᫓\�����KmE e��5:����P|��I+/��hKR\��>�pG5�t��2t���.��ؗu"@hX���?6�-1�N��+Z��z2	������$��v�������ֱ:[���qvv��y�̮K��ǣ��&�x��+{��kqr�t��wÃ�ǋmߢ�|���Q��h�jR`���g+X�I��kY��U��j=0�4$�{�����.�|c�-��z��T�:��t����>���<�g��O�O�p\���6��w� ���@���uQ�n�t��|�r�-���HȐ3j&T�ԙC�{��_��E}ؐ�<z�Pi����Nf���.�df�g�ʃ6&��,1Ҍ�(�YO�+˗{RN#��s��ѠMf�L�Z�7~7>���hQ1�v�lV>	�x�n����;kX;q˃{�����.5���dJ�l��p�����q����*[n���ļo�y����/k�!��-���D%}��槔��'=��_ ��@�t@mK�\-:t��Hlc�Wi�_U�ut��KG������1-ܱ����.�̚t����;sK�B��/@B׻/=���9��t(��} �`*��9OBdE{�Uo̵�.*��g�C�Nw��p�`\zn3H�JA)11�Uز[�LX�}�GǮ�^�u*�N�]a���<t�c��.��2�r�A�SHӕq�W���vHEN����m�����v��Vi�mj�}�3OqAݞ�m�T�Q�꯾�������輪s;{��B�8yc����FdB�J����C�ӊ�=N�.����E˯�V��QN[_<����%e��3����D�7j=�lwr+���
�g�8+c7|#�B��h}���*vu�}���>�4Xiṙ�T�P&����z^��d#��ui�z�����V"H�9&S�3�:��]B��в��c%[�Ԩ�
���9�<�v��&J�˛_���(��ʣ/te��e�w6�������]>:�ζ�}�,�2�ǹA�q����U��<�UA��3��x�/O]sv2�B����S� ;��u�w8�3+QЍ�"����,r�/��oHV���Ţ��F�+��f�VYB��ML�dk��/��
���"<y�.R;Ys	�~�����d�q���,5������z��X��Y 6�=U,�Ʉb��>ç�s>5N
���E����fͧo�\i�ebO/�ɹG�Q>�Ȅ�'i����L����7��s��J�j.�yrK�*�]��[ǂy\t��V��{���ؖ�k5I)��"�x:�u����u]��W�Y@�&�<zcA��t��Ջ��1���Μ$#��?�c}�)D�N9�	,c�V�l�����_iR�8,�������uvnlס����L�p��E<c��p�i���F;��lZ����Vdk4p�����P�nT}�	֝�ݥ�{Fv���n�X/�G.>�X��4��싴hc�*���k돮��\�l�vnvs�����*�5J"(��[Tb**��Em*��	Q��Z`C媩"�"1��Q���V$I�V(1��()iC�
 �c��b���Ȳ"1�����e�1���5�UEDUkX�Q�J"��a��e��TQX%�dTZ�UE�sj�W)P�*�Uc4��������`�("�����`����
��KJ��EX��QJ�T�WM�:K��"�1Ub�"TH�U6Ȋ��)P�0kV1b
�Z��������X*��Q%lcE��QkUcmQ���b�`�1P�"�b�1`�PVf�A��**�b���m���b�X�"���((��#X�TQb1r�J��QU��\2�AQE���(�X�j�U��b�E�(��Db�QF"�+��Z�,�QTAQ��PEbłb��P�
����"#Pd�TAX�b�UAŪ��X����X*"��!Z̠TŪ���Q��֫A?CY�s��`��e��ظX-�b�J�,=��m�d�E[��P�S��}g|��}n����������hȺ��o�}M4d�G1 Id)��w;L?�}2�T������8�U��[��y��d��Rǔ�&_#=��)���WM|e;��W��Ѕ�y�YX�AՕ��7�5oX̶�Wg�۞6��خ����R}eAW2��4�os����֟_�d�����ʣ9}���IƮ8�\�˧:{�W�����x�|v�櫛����ԯ�ɇC����;�O_C��+���E�XR�ׂW^:ū1�y�=�a>�(N��ڒz������˵�VWδ���8��r,=t6���o�߰���v�h{�����|��T��њ�W8��J���X+�j{&m�@�{l���tX��wPX�p_c��|�N'(k&��6/�پǻ�#�[�s��K;�m͌m�}�ʷ�}��]w�e5�o�p �Z�O/�'7�p�ȹt�6����Vs�S��a���B�R�d,�H�2��y>�l�b�.�s�Bt%����sܙS���\��u�E.����w��n#�)S�m��=�K�:�5H�G1�Hz�V�ژG�9����)����3��ɰ�G}^�}O-
=p��f�r��K�ꙗ����J�;�PL�$<:�]y�}/GXɤu�l����ݲ�[X:���S؎��7�bw���Ϧ3���u`�U��W���ǽ�R��o�;J����^�+���J��NK���cg�+�w:��0kki�7��������������'l{.9݃��_�۱(1=$>�N�=1f;]���y
�~���b���g��r�r�^��O�yF�<��'1�U�.�ys�j��xרxs�X�*�2w�k!{C�Y��fvؿR���
.��S⟽V�u���J�<k��8"��;��kɞ��g]z�}��Ƹ��iɽ޹V��&1zhz�5 �`�3q����3��ٖ��y�����+ԃ+���\U��|;��������|��b1������[գ�Ʈ?l*�^a僩b�i�C�}�¶����wpк��$�������x�&���]�.Q�A3�I�d3�]����o�r�z���]�憀���D��<-��Xٞ�NԽ��y����w��:��t�D�J�IN���Ra5|V�[m���É��#�6e�{�t4��Ĭ5��{LT��[�a�����c};�0����ߑCv����:�2�J>b��s@WXA,y��"����x��=Y�~H���8xD=@s���;z��ʻ���I�U��P�+�r\����ۙlf����]8͌f�ΞG#�����m1��Y��fϺ��YJw��k<+Vui=��ӔÃH�"�w;���{�-uF��ٷ�z�Ӟp8���V�3�gz��B�d
{8�q�V1)U��_��3��W���{=����r�����A���}�������v�3�{�S�1L��^�ڭ�V�e�G�2s]~��Z�II\����eI��=�pmmbE��^���/u�c�3�΀y��9�$�W2z�J'ݛ��T��l8�<�	�oq�ژ���_�%�����̬�z�.}��fk�>ؖͅ�9>ў��O����zS�^Hש�����p׫<�w�V3���$�^��+���Z-_m_�R�º��;��s�}�w�Y�+��ژ��8�	S���y���[��ġ:ِu���5����>��=#O��ӥ��՟?�H�)4�]�h��/\y���)ܶ��';�n/zV��rҏn\r�����9Ϻ���<��N9���<=hZ���ǜz��U���]Mn�G��O��=�nJ����~s1H1fv�x��W�����/-qX�q�;��b�be�.y�]{ى�����M�}e�Sr{p����k�F"�!��B6n�[Z߂�r�Ijꦂ��Tκ;-�}����-�ٖ���M;`���yu�\�q���4$t�,�<{7��en�������]��Q̼���ZY�������Uv��bq(x�c}[�����ܘ�i�ےcn����,��lEN��9�,�<��@���_���<�:��'�U�Q[�0�)��'޾�*��{�cǷ�<vp5B׾�aD
5׀�7���������PA^�����vv��Z�S�:n�����ߣ�<C�^��7���_���Ƨ���w�柕��X�*��d*i�.[�r�C�)7�D:����f�;�9�B�č�{�ߴ�vUԒ��n��f:���.��s%J��n/\7�ٷ�^͡�޹��Ƶn{I��;�T�Y���@M�.�x=3�w3���;�t�+��mcl,����Ԙ�]3� ��%?[����ҟ����^���9}���Ekj�v���}����~�ŗ�.T�{���e�<�͋ɛҼ�1G��k�'�u��'r�uH�9>ӞO�� w+[zWA�����Ƴa~��T�e�ns�����#�R���/$rn��a�^
%k�\Zm����~�^��ft��{Q�	����w%%�>ʙ{�������k9����2gy�\�mWzL�I�9�)"%_�b��]�! �`�	�c�X�㷒�yc��뱺e}�Yo'+�{=���̫��37.�h�ǅ��\}��e���	��Z���ؖ���UgU
����{X�����Bts���[����:��������+S|^���L��L�ښ�{Y�[0�|�sR�6qKr�l>���HV�J\z)j��g)*��o�-c���U�t��V��M��}��k{�����GFp�ۢ�{���e]m'.�~�]��g�HwRw�Ӝ��[����.���z�������2��o���u^y��9�dwk �����恝~�������\� ��C�'�<yN��N��1��w�/�}�W���u,���B�͌S�úsV��9I{À����f���Tk=�n����&o��~�5�Y�[���9���ȉλ�u&�Mɹ^���s�_<_�}��{ժ����K��`��v�h�x��ru��(�|����9/3wf�����y�g�z�3΅��u�����{����Yb��|��1���tٿG��=�rl^���z�aO��jí��M��s<{��]��z��3��6c�5��o��7�8/r���=o��L�x�z��BZק]����Ny7ڽ�>.�����x��)p���n�P�{�"E���y
 ���ݪ�}���=a�KsnUŹ����Y��J=#���J՘-���:�Z�*:ҡM9c�u�ˆ�U�V��P;s��̞���,�>�l%����E����-���:SB�q��@�-�4oȹ��ٸ]�0qĸ �\�EՙЬ̐B�m�c��@�u®(W3����W���MK����8C;�>�ծ�b����������#5�or����+B��+��/����L-�j��dե�-s^L[�T���Qʞ�{#;~����W�[7�l��1��:��:ԛ.gk,�ۮ~r�<�s���n2�5�2����"�`,'q�s6����譯xǛ�R����
�w�}׺j�ȕz�F�H�Z���8q��x'wQ��w)G4;�O6��y`��͆��i�U����/~�ot��(�J�U��`̀��˞�V�ۺc~ݐp}|=u���v'�87�f���2�=��FJىWэ�·��gv�Sr`�b���}��v�.Xm�rv�\�^��{z�l��F2��Rkkؙ>�Sk����T7#Y����j^���ϦJ�{mܿ���`��8l���׽�R�m���d(g��ȗ�>eZ����c���)A���Js��e��]w�[Y.���W\Kykr'Z�xԅ��(����DԱ�w{c󤍡��ՁS���ٱ�e^n:}^�5-f��(⧝�T��읋��VgwW�rL��s=N@+=Wn����:��=c[5�9�>|��>������p�O���R3{�y-	��/���(�e�h��;��I�ϻ�Ǭ,�ih����g^����� k��!���� >�;q:�-�xz��{�����:X���{��92w�?;x��c_�R+�S��������x��wpQ]ϵ�����@����So:��#4�}��\���3��]=�:b��Y���ί<��0��V�<��Ì�ʲgV�I}�9��t|����y�F]G�S�OO� \�]>۞���]��vX��jo��:�\�B����J:ǯ�R�.�y�t<1�����M�{X��n�}�yZ���:��2�HU����b�8��1�tj���Y�<'��O�~n�i׍�t�+-m�x�(t[�*"�u!��t�ݺ��+��(�"�����@&x�Y'�T^��d_��B�iʰ��.2��V�\sv[T
8�ty��y�1�F�I���&�ӆ�ë1��依V�����*�"����n�ܓ�Pg�e��5-���$XN8�-�8s8��C�\7'��xoa�I�[�<>s�j#������e{k�\vw&v8�)K=]�P��|fU�ġ���L ���gwn½��(]1�}���~7d;%s�Nd����%�������VN�ܞ���-�U]�~�}u�m`W���ܜn�c�ۓN:��;�;���D���]��k}~w��=�+����l�nWݳlG}������@��~|�)������܊�^�c�Տ+Tr�������ce^�|�޿dm��o�^d�N�q�՟<���g+� ��'�0;�d�6�[[J���:�9:���^�;+��n{��꿤��;P����6�η���69�g�y�I�N#���Y��f��+7���ɠ����T�
���'�xԅ��I�͌>i�]��ܯE��W_��s{<��t�z��3OH�9+qD��7U�=h�')�[nb���´ert}�"�H���a����j�\�I[�'R43cb]>�7�y\�*��b�N0�����r:���=����,Ќ�`=�f�pNs��=���㋴C.�D����D�K-�K��EX���o^Fw�=V��:����V�Wg��d��݁S�O]x]�����2W��f|�������}��c%�gc��͙ޙ���ѳ��=���5�VO �:�F<e����z��fO}W�.�
�JY͝��#}��mVb�>�pQ������up�qq���C~�z:��F���2f�|/��
Ḯ�4���ltBoqUQa롴��[e������ޫi� �Y
Մ����������;�\ʹ����^��M���S�7Gv�L�&��N������,��h��_�wr�;�t�69��6��{����g!%��K�~�]ۇ>ÝvQ�K��m65n��_O�ѽŕ��@����K5T��U�:��z�l&7]y#�Φ��^����[��=N��8O���y�K�דH����1���ǜ��f06��3�YY�����6��m���4�&9rɥ�G���7�T+�	vtd�W:PO)�Z�L/ױ�O�c�E��F%b����ŁU�0�t��z\�{�뫆s�;�<M�d<��"Z��R�=E[o�Q�&e�i�Y4�\���S�u6�e�J�8���@�p��� l��ڣ�]N�5��֜�$,�_{�crD 9�{�~L:��	�o��0=E����P�u�Z��8��wጾ뭨� �Ǻ����iӶ��pݴ�<��(�0CB_�Osq�&�Y}Ow8�����'��/���rT��i�o��!#d�%$k�gt�2CM='�΍�2^��j���^�vs|��#�4��^Oew��s�A�H]_�Cn����f!V�R��ȎT�fT��� ��ɛ�)�OiM�=�3� �+��V�{�7rak��꣱i��Y��7�H��ټ�L�ƥ�0�&�f�};0D�JA�t.�]goHʳ�=0�FZ;ed0*�a�.#��2��=�����,��tJ���31XE���twM΅��.3N��E]�H��0��vwP.c�v!o�:x[��*X���,��n#����Z�]�Ĥ�6M�wux�|{tQ�u��;
w7����$^[pq�������s��Zʑ������5�J��e���;��ۚ�WD&��X�4���l�nx����ݭ��2kљ�S�yq�]�i�(ALm�E�t}GS(�0$�+/o/TSU[]�g"���)�&�E��	��p	�\�,�U�K�o Hn�x�,�l���Sʸ��U�5$�P?!D⣑ ��"i�$�a\��e�~�sH��`�;��� RA�bX_���P�5>d FVa�w�Yt켵�C!@�*�b-ĥ�@�*d�7,}f�EE�h�2��(���J�'x
y��4
�� e�
�u<WTM�nU��e��Aj�C92�6��Ed��Yf�]��[�ʍ���'��k�Í\�&\W�g����5��3'�蝹C��W�EJO+Q*��ݓI��h���Y�L�x��d�hU'����Ue���`�S� �%�#=|+��e1��+�{�}1ɢ�mI��qTަS�&�U��0 �}�.��Z�ݭ�޲�`�J���f� _
���!
 L4�"^�tK������������O(S��[�ӓw��V�譐�m�@7P4oA�NnǊ�*�T&��D���Z�2��b4��"ut��f�AL��	�β�
�Y��b痩2��*2�[g��&+�Kw�HXD]0�wH��R��q��瓍B�}#��|���=)=��]f�:����V��~�bvWM�.�7�H괫82.�%�
n�����5@QCoJTN��|PLђ
�שhn���!�o��w���A��fi��h0���uj��[������e��5�aS��A��r\�X,U@F1AJ�UEE����X��Ub��
�YQ-��TEb��b�Q�2��X*�a���"�*��QE0�*��TH�+�-����X�Qb�#V,�UE�QQ""*��5sJ�A�2�-�,c�UQb(�F"�V�TE*���
L�V"�TTAX�,TQ�J
E
�"1b�$A��H��Tb"a���H���"�1P`��*�����E"��VD�R,Q ��J�-�UTQcZ�X�������X��DUr��F*!A�
�,�QH����
����*(��UH�����IZ #b���UdE�1�1Ũ1V
1UDTL[�
8h,X�"�PAbSQX��G7�c0�He��b��*(��Q �((ƵG��U�EQdX"DE��V�Q��(1R*,V*Ƞ���"��,UDU����"0PͲ�@X��QEc
��"�*��b�Z�7(��r�IQ�S��<�������s��,�	g�`�}�6wS.��e"��7�NX=0.�'s�
Gl����X ,e�t�AfG÷5E�{)��^Y�^/�s��wS��]ՙ8I�9S{��������{O�|�9��mWnA=���ok�F��l(�L�4绪��]QW�Fz���������u�7ΰL���aT(���V�kQ��u��ڼƞ����s�}��;��\�����9,yo�u�,,EO�V[���/�{�ߔ�ɶ�
�\��[��=�#��=iz9�b�۷��v��M\������>/o��w�q��Z~/��U����������Fb�9��}��C ���s�tͻ �Q]�]�}Z0$v��z>�}P�pïq��-<���Sq��H*X�<e��(��*=�Kw�7��v�m=����b�|���aP����z�(L���G0��လ��0�	��MǺV޸����+�����چ�lj��9zwk���+�Rݜ��U���Ru���a�/�/@W8P���֪�c���d�ԫ̱�YF�t�a^�i�C�CzƦ��$�L�����:��B뵇��IV����r����Sݙ�'d�S�U�~����v
z��_�$�
��~�j��1��K��]��K��[��]�3d`{������7g4/+Tp���v g�e��K��C���a�z������}�{3����#�Rd���g���:�g��w}cw���1�O�wXۑ�J9�f�6��F[��k���}�6�sg}(�^����m8�������N�-U܉�y�1��Ź���̜�_����t���y���{�I/`r�Vܛ��x���w����k�����W�����p���X/k]O��y�џJ~��oq���]�����X����ݑ9Q������s޶���^����r�YZf�y��ǰ�]쵷���P��l��7��{���:�{x��s��i�����+G=r�I-���i��}����B0����{Y�-��CCg�XǍJ�����F�+!��̹�/��Ы�܁��cE��;bz��n��|�@�G5�cu<������
 ����dGX�x�S�n�$��vu-�\w��_��Mg�X����#.t��W7/�����u�ʁ�m�����w,.��;���ż���#�&�l�:���	���O��7�N0/��0�	�?'P��	�S��ɶO�P<�|����hq&:�d�0��H����2>�U��WT���>{�޼,���)�N���&��I�|��!�CY�Y��|��3��/��g�0��'�O֙`y�H�����	�uFq9=�W{�G�:��HazcX�'Rh��,>O�'w�@�J���Ğ`m3G����C[�Y�!Ԛ�ؓi�`j=Hy��0�1a�Y'�������;�|����]ӝzI�R�����L�N�aY;�\RO2h��)4����g08Ϳ�͇Y�a�����!�SHy��}�︄~~�}���s�G`ܮ�1��g\��g��|H��>Ch�N���?[!��`+'�1l3�`!P�=��O2h�0_�N�����!��{X���#��E��>�>��%=�O������y�~�7q���'N0��i2��t}�$�O2z�&Y�Xy���g��VO$��{��00�{~J�|����P�?!<��6�!�G�?a����^���y�־���R�q�?0����ɤ�E���6�XG�HN!�	&��y���C^��:��,>�q G�M��@�>D3���
e�ou���7���}>Λ��T>f�C�����|��wX�	�mOo�ɄRL�oy'Q@��d��'l'�L��a6���d?���C���0�=����.������I�B������&6�<���X&�i���$����&I;�'Y=lϩ6��N�k�C�'��	�]��ǿ���w��:�xk�T�z�k��C�fP欟0*g{E!�C���E8���]�u0;߰)'~���1l���d�'m�[HW�������u&��3 �k�z	��m�\�4:�q'�V[�@��Y;�-�<"K+Zck(�*`�Ҡ[�[�6��(Vo/r��p#?kw�9�V�t�~�J&�Q�V�t����SX�W���&p����tT�z};�k�����i���\�YCv�4_{��� [m���-Y_�|��i��Ȯ5�`<��Cϙ!�2�}�u	Y�5�`�����̟$��
��O�?w�dXN�k�N5$�/y���/�}����mO�9�KAP���K��|����e�4}d8��d9O�N���C�8��}y���Cޤ�����d�(N��IěE�G�� ���~���0g��������}'���&��q6�Ěz��7C��I�q��d<�>���	Ě���d<�ć��0���VI�1�`Y8��W��m�=G��jt<�y??�}.��'-'��ִP8ɿ��N�/��N��d��O���N2Cl�!�CI�\�<����l?!�C�Ӹ�N�"��-�y��j�s9���
�+��;i'��u���O�cy�O���y$�_}�i<�y�q3��,�!�>g��B|�r�R@p��m���Z��;��N?�SG��Y��N��9��Qa:�ޱI��&&s��~a������y���}�N�?C44Ͳa��y���a6��a5�����y�ߌk�_{���������ms��:��S=� V�qd�a��������Y�ĕ�&���:��0�o��!�`+?2a�bn��7�';��R<��T��U��W�t�i�M��N&ai��`g��:�̘�4wX��&g��sa<ɩ�w1a�~a=�c8��d�ֱ���G�q/+�}����������~����'�6��M���he!�w�%IS��Oɛ�;hN3(dš�{a�N���I�M�`Xe?2��ߥ{�g��ߨ3�8��P*���@e�7�2CƵ�B{b|��I���d�N��$Ry?�򤕘���N����bT0�2���@�SPQ�Y�{}߃7W��Y]8eG�߿&9L��MYl��^���E�T���ٚ���FX7��PG�T4��i�EJVn@�0�yz�ӭ�/zwv��v�s���P�<Ɣ�#7>�p�aw)��T�9�x�',}���ׁu1R�.�@�����U}P�͝����5��\$�d���<Ρ<�؁�>f�?l�	����!�&��'ɦQd�o���I�_���{I�jv��:�C�^�yױ�������/�8��M�C߬�+>w�T%`|�����!����O��Hm����̘VI��<��Y>@�`z��	�O3Xލ�n,����:}��C:���znÌ>Ŏ����R|函d�!P���f,�`c���He� m?!�'ǵ�h2�u'زi�7�u��������y��������?��s��8���z�*5i�~�&�8�Fm�I�3�:ɤ�!���d<��e�ǽ�����~�a4�߷�g�C(jw8���>I����$�M�xw��~��p��Ο��*,'��O�~���~@�����!�Y����hk��P��2��C�m�a�Xq��~N��"��!�{�!�M�þ?gw��5�?wL�7�ٿ�r�s��i�������>��}�d�N?2u'm!�P��>|��Hu3���8��'�!��d37�u���C,>��'��8�럽�q{�7�m��s��tY2�E�$�'Ȱ�)������Z�u��}�9l'Y�<����`u&�'ۤ:�y3���>���D?�|?�k*vJ/}������Z�M�P�}I��{���uC<�'Rq�v�����5���I:��`�x�u>α'|�`|�`u'�d`C����C�������?o�g���γ���i!�����<��;-	�P�&g����?!���d�,�M{9<�ğ��e�ul4�>���u����4�$�|f��>g��gx�.�v�W<�������o��Hm3�<r��i��2�����8��<�>=�Hy���QE��Mϼb�I2k8��jO['�I��w��u!��>���_~����o������P(�o�U���A������lcq���㡪��Y�%ak��6��E}�R}��Ԃ0�<��kgJ�V�U�o�3M�����EKr��	D�ޑ���[G�\�*=R����{&,��{�Wu�������G���|��́�ﴃ�~`o����g��O�9�i�ʐ�{�u'�0�5�{2d�h��,��2k�M�	�_k8¦�f���l�����w����%����T��t'Yk��l���Jβ�|�m?!�jb���m�:�3��8����9����Œu�<�g��p�C��9�^/ɋb�Y��	q�I��bXT�Ok�!�0�}��!���
�$:�F�6¡�ް�œ	���yI��y��X�0�0�q��>�_�߳�o�0��=���&Y4N�I��I���!�~d�l<��g�c?}�a>���Hu&��O2��N���$�O&�<�	P�����>s����kӜx2ɻd3�i0�<s؀�VLs�ۆ̏,Y�~Bu`~CO��!�C�~C��y��[��4��@�vM��>�A�%�л�	�ѽ��.�u~��a���I0�{�9l�I0�e�� Va��8Ba��?3����,���5�bVi�5���!9�5���;~�rUݽ��~��ӆy��UiO2|��'�:�q��Xw4�u$��&���a�e��I���m��`P�������~He��ql��̟��i�?]����Y����s�����'�O"ɣt��u�֧P�@�q�'XO�s�:�O����`y�RrvɶB����
C��y�ھ�y��k������~�u���a��Y��`u�Cl��IĞ������u���ɽ���<��O�0:���0�a��O����s!�?3(~��޿�W;�������߯y�j�ƾ��BT�x>وM�2{�:�L�VOg:��&��yIğ{�Im�s�'Y;l�C�0�<�v�q��u�<Bu%�w����+C�#�|���=�����id�
]7'�%�D���3���Z��
���R�ͧ�>��j�ڕ�H�����*�b�J����8�������v�n����3�x\�/�����2x����2�������Ϩ-��NټotM.\6�Ǽ�}�W�UTQ�>�����g�ژ�}!��d?�oِ�u�X}�o0�B��}�,��C�q:�L�T�Ł�6����n��@����d�v��4����u��O'����7ݹ�nq��~Ǡa�����'�y���:����H~g�{؇�K�=�E'QBg���N2mR|~� ��>�󤓨cX���'Y������=������c��y�~@���v���:�~�<��>v�By��?'Xi!���ć��0�[�I�g�{1I�P���d��?ZP8������'��s_����k����'�~�0��>��g����b�0<��m>���L�n̇�5�q�Y<���O!Y?o�Y'���,������w��ٽ�����y�Z�M2~�Oo'��|���	���Ӵ'��f��>g�N�O�<�1@�	�s�2�uy��L�u�(N$�7�o�=w�~��u�g|�>~�~���N$�}��[	�ﵓ̝I��&�d�l4�.�fC��١]��C?Y>C����g�0���'�MKa��E!~�����9�>���k�����.p�Щ:ɄS��C��8�N����X|�a=��I_̚�ku�i0�{{�O$5����I�M�L>�� }���
#�c��-o[�����5��C(�L>-�R|�C'{�P8ɋa�R@����I�G�Re�	�ذ?3�m���~�0�~C�>�:�c_`�d<�G�޾�����~޻�����y�=�VdҾ��):��8�$�gX�C3���̘���Ha�nҰ�dyE&�:���3�6����<�~O�3}��ֳ���k����������w�a<o�!�C�>�6�,�G_�H��1?P�l��z�̝�C'y���I��1�T��q�a��ݢ���	���~�7���y�g�%znя/-�`]C���Tr+�#@�4�$�z���0��ݦo���ɷQ��畭R��W���{]���i�Ӵ��a��4�g̊��f�;i��FX:-<}g��ҝ=��1=�b���t��s�# b����w"��.:]��m��}��|O߻���K���e�x��4*�|������ݓ	:�'���O2ys� y3���I0�<�I�C'������v�? �H�֗�8��{�dk�򂽋�L {E'�Ԇ�������>��*l���̘E$���y��P4n��Y=i���&yC�XO�k�G��b�Q��2��/�[��;��q!������I���m�(�*��%N!�C,������>=��d�I��y���1��'Y=l���;i�A�|?�������ӿ�����~sR�����i��{�I��Co��l��ؓ��O�׽�Hm!���b�C�C,��!ԙd��y�I8��}�-�N?��:��`h��}]����[����:����VM$��~�8��d��'�2k��O��!��ċ�̡�Ru	Y���\�����ɔ�"�g��I�������UR�����#=ɷ?Y�$?���u���&�|��t:��M>gC���l���Mr����$<��s!�����<��8��,�E	����>�}�	�=�b~5�s���$ywx6�
���@���cO����a<�ݓ�O�04n��f��|��L�M���:��u2[!���w<� ���R�ś�u�ٚ6^�!:�p�۟���}�d�(OMci:ɻI��0?2k�޵	�ՆS�'S8��lnβCl�|c� u��jr�!<�����i����<��w5���{��M��p�?fa���O֒{��9l����I���蓬��2�d<�A�N!�6��,�i>g�����e�����:�������Ξ�R@�͇}d�Oȳ�:�d����y�������&���~a��'��	��?_��'Xf�f���'�����YZR����T[���u�t�2�y���Ϟf�p��yd�Ʃ�5 ���Y6U�-e']`�k�l�g�]�A����zi��(�[�ۼ&g�%o
�w(�u��c��g=��@�9��{���n�Y>=�`���=m���wF�'��}SIb���By��HH�������u��o��i�'��П����i���5�N��L"̙�y��;�͒q�����'�g8��2gZ�:���3S��Bu��7�w�_���c�:�5��·�T������ǌ'Xy�i�?02~��O�0�ŇU�q2��<�'{�u'�1hk�ć�0�3���y�W��&�N�뿀d|����e>��j;��O�d�=��fC�������$��d��2�ɻ�����uY'�͡�N�<�0��L���d�0w8��O���y�߿=������$e��>�
�CI�����?2o6d?!�dοd���՚C)����<��>I�]��$�q��$���y�ֲ��E�3��L���<�߽��/s)^\���=�c�O2j_`P�?!<�q�C�m�ٲ��'�6{d������4��Y6��O$�/�&�:�9a�~��>7�O�������v[X�}u�CI8�C�[��i6����`a�	6��E	�����~Bym!���`~�~փ(O����dڲLkx'�:�&�4���������s����Y�߷�Bu�l�ń��{a�'��l$���{~d*��f,�`}ևq!�=���d�=�a8�'�?�B���G]_A%yi�Ks߸��ܕ����Ͱ6��d�a>d�?3oRO�����y�׷��y����bM���}��?$5��8�R �u��i�Ѵ�������*�{}d��_�}�*,'2q'���M��>�!k�#�`l����@L�ެ��<�^RK��`�:�}�y�~���R�| ���eu��7$%����9��96$�a���*̺]�~az�4���Ҝ5��fm'<��ɻ�t�N��2����w�/z�� x��wGt�Y��������aV����C\���8����Of_We����(wKo��ݩ ��z]vJ+(5�(e� ֎c��Uj���������ˍt뒊ͣ��e�)�oԨr�3x��C�����Nv��۳��z�h���_҄�'�s���>[��8�M��r��/7}~�c�����=<Ѭ��d�_���yH�g�X�
�v�|��j��ү�,�^�y�fD�Yk��{^��������;���!px�}�b�5��B��A<��4��;�e�D���e��p_��B�6hH*c0_x����/��Q�"Gb�ZW���e?&.��J�݄j��V_Ea{��f��`����1x��˚����n���%^��������U4��Sks�ZqT�W+>cigx켷�-I��$����\.O�*��9���)P�&��~�<���S�D+}�l��{~D�}zd�H��}��>vw�/��Gբ��-�g�C����UF�T	f�1�y0���s�X�	��\ңٛ&3R��$��L�^�s�\�����ʾ\��vkg�؋Z':�gmnx%�f�$�i+�����I�͹z{�Y�I\��+YB��nq
���ѳI�������u�ݺ�Z��.��\&��Kz���P�T+i�����(dWf�5�-�M�L���-�k!���Y�I�8�j�:�U��g�w��QAˌ��|�E���;��x�Z%�:tm=D\��cí�~2;�(D���L/>Ј��\�85!ip�\<���Z+9��̡�S�sz`��eR�!�C�\�/��x����6�$�>vC��V*ʮS8v:pš�`	��&M����E+z� ���32�����Vyx'�tM���H����YN����sڂ�!�w�Ti5��}�o-���<m<]�Tlzzǁ��)��9{l��k����Ӧ�^l���Tt�p��H���K�Y�����{���[�v�ϲ(1��z)�b�<V��`�1�7��� ��ޮ�`�|��lv�W��V݊���aL���K���]J������N��`�Ox�L�8�UΨcIԓ�`�3H���,�鋉������q��W�`�N{��\5w.sr˭��{�s�%�	�C2��Kb�Ru+N�u�K���^|Qřۆ>�7��w�Ĵ�wQ[L
K����E�uT����FJۻ!�IL9P��V�Py"*�Q�ȧ@P��o�él=j�C��%��O)v���ܽe�[�U+	L�9������"��s��
�{�A��Ĵ2��
�t�PAP�u ��_L�2/R�5<mG�Zo��|R�)���#�P�řa�"�\�W@&�6Q�b���E���++%7@�
���Y��mF/�m� ��x=9�/���a�ɠ�&�q↺ps�[Q�ퟦ9�������4�EdZUel���,�Aᬐ���d J* o	2�3lR��������V5�7�����Q�0� ���GJu��X�)��	��
��f�d	h�~��cJuc�@-^%�Y�mT���/K�d��iʁ� �c2�8� Kõ`�>����g���P���տ@M��[@}���+�H(���Y��u̓q�ZM@�DZ*����@�+�C필,؆�D����ㄶ�AR�q�ì��9X���(�:�i��h���;�3:�8	]�|��U��I�!X_e-��=d�&;^��=-����ܮ�`�����c�x��n�=GZW��E
۪��o6v���Y���.���x�(���ю�:�]���7��p��hO���]P����0Vˇ��.dS(S<馨�9S<)�?cc��_�_w��]�����N���m����#x4��^ʻ�78��q*ݛI:��սKV��W!����`0*�X���qK�TA�T��QQb�F(��X�j�UTp�����l�AX�ł�����ETL%AQ�eET�EQ���Tl�Eb�"�TS+�(�*�A��E�EQ�Dm���C�DD\%U\2UE�eEh���"(�3)D�,X�Tt�`��UUV6�Ee�+�C6X
��(�F�Q"* ���p�H�����Q�(�T�QȸB�-���#�UCU����4� �[1�����UZ�"FJ����b2(1XTiUAEȤR8�$�DY�@D�+Y2�1J**��J��b�D�"ŀ�`�.1*Ԣ)�dL%U�� ʅt���+mUE3h��*��X�f�?R��ݽԞ�&*�wݓX��#RG���t����ܺ�U�v�Su�ٷ�sSsi�\�����v�l}�u��(w������}w�I	��{}���Yჽ~0��ٜ�
jc�a���?R;N-pVZ�₮�\��$4���goyU������{��am3�����r�r��;�Wݛ���6WF�̊mu(�j�}��g.�κōh#���r��΢V=�Y���F�o�N�æ�{Ba����S�W=V��g��������h���C��K�k�vh��+��^i����ު���=�C�I+��6�M`�+OIVtyQg��+��4:�F�9K�=� ��~;�3z�V��di�[��fp�:*Xk�����3ხ�gNRg}�����V;�f��m,������ϖ�������e��d8"�$9.����x{:�����%��b�ג��/�d˿��+��r���=^Z�L�>�!>C��~:w<�ƨQ��� �v;%	��Iacִ�[U�1��\2�b�	[Q�w�Y�?�=+��`>���9�0q�Պ��ۨ�+>�1�JØi�+�Q\=���\��ǂ����1��Oaj�Z&�z�/v�d� =Xg�"���%�Z<���j�ې%B�:���G��oRO4�^e�i�xJ�Vp�������͑�r��3���m/��Q�Fc?fp�y����n���99#][z���;+���ۭ������}��5�ǝq���v�Щ�¯ޝ O�AƠ��KI��Y��g��5���6���0<�_z/^}Ix@�Q��c*^�!F���p.�\~�TA��w��:���j�is�r_�z���W%p.$��:�NԢD�ө��%����_{�{�hue�����?��h[�ټ��D��4�ݖ3��Qe
|jm�N�U	5e}�!h���g:��[֬u�zXXw u�����`����<KU����bA���9�Ә��f��f�*��lJF�.`�.��T)�~=Ba��(:G��W~�v@L�� ��O�[�vi��q\��^��G�av���~��ބ8�{H��+�i�	_��3n\���k�j�x���<�o����x؜�3!ӳE3x��;;w��ޗ��{����ZO&C��:Ε|�ۤz��l�%Y��wY�c����^�fy�z�1..��B�����uY�즴@ƈ��Nĥq��:���[B�c7Sݎ{���`�勐ܪ���fЏL�;�ĕ�tGv�l[|Gm_a3�p����jAgmK��>(/=�'�l줖����.�]�kTwo�no�#�>����%ԗ�S?\�D.6#\��GR�i�����O� {�s:��꯾�_��O3mp?�������<54��8F��niAҚ����{�+A��ͼ�x\��e��Y�s�v������;r��O6O�b��֫{���gY-p��U}6GZ��I��~{^'ɉ�Bĩ�����`�0;�6�DWg�9�n@�jn��t�΍�_������Ҭ�R�^P�Y9y-�r��0�޳�#x����n��əϟ{L��5�\�9)�._-��Aq�[��
6*�C�N�2��2�e.�k0gʝ%�Yފv�.��P�+d�`u��
PP�"�rɔV5�b�LV5-�N��}왹�dp�x`6FX�ճ>I���Æ`(_���4]� w��eq�]���ķD���<����r��I����R�V��%p\R'��7��`6Xr�@����U�cu�W�����}O�����`���^/ҫ���
U3�%Y�T5[�DeR�X=��>Z����Tf�y+agL䊵�f����W�v�2��}�5uV�R��r��j���'���An>�.����P�g)�s����u�~�k�
��1/wn0��j1lJUv�)��;|Yǥv��Ϛ��]����T���7���3kA�����Cy(Xv�uG.���s`�+��j�@��>WE�!����}����SE���[d��7��K�߽��׾�Sx[��[���?��h�^o4ؿ��.�$׽�:�zv�GS�sp�L�_���p鐮8c�<�ʱ7�N�y����_`\�o���[YqkH��ߘo����T1+�[\_��u����{U��*�����)�����xf)��ݪK��ˉ`C����w��8�[>�O���\�}���ڭj�Xa]s0��'C؃>���L�e�0{��8�<.O����w[?T7�<��}*��
���5�fm��j�T0�Ch&���%���UAt���2����Nǖ	��j��]��b��͡���S|�EG>������6T\u`V�κIf�|׉~$&���y�=ib+mq�Y�R���@�^��h���X�_�}p��rUw/�%&g��;��o�g��4��,�;�W¹<��1�Sv5P/}r�����
�<���ݱ2�'���J-�K�i��������͌@�f��5��U�3�U��P�+$4���n��
|ϰ�������N�\�>;ޒ�O6f������:򺹩R\]A*�S}Ӏ�دbU��G%�뤞�]v���i�{˝�Ǥ[:>�b�����#���O��z;eU���HI�p�%q=p[:�m�xe`M�S�ie�7���|>��I2A��m��`����b\qG�\��߅Lv]p��|��Bƪd�a{1nA+��L�ܜ�����g���TYhp���&u�z��P�`����̇~���g�N���7i�,�m"��J�и#na(њ�6�m��]�.��P��^��x�AM�=]��&�X�����Dyo+�9BX�g+Z!�)��3�Ja_�G(Ij��joz��VK�˃˕��*0w�Za&�k�ub���X$���a��ud	��	T�z�빃揍Q�bfbɓ+<׾����桊z�<r:x��=�|����x�g�'9�å��E�6�g%��,�A�.����Q/r�.�Kf5�0�sR=�{}�peQ�f����M��Y:F�U�:\C{�����`tҡ���J���jS]303<�����o�G�_�{�|�=�S^�+O��:0E���d2��T/�;�miؼW>����;z=P;g���yE܃���֤��L�R��޻���U�hg���V-9L�lrZ̚9��r�z܌ц�W:˞�x��{�)������LkvN��6������u>�fͤU�{�����7�$`&ﲒ{�rx��N����c)��黮J�-�:�+rb� �7�؁52��?�NѡN�x�; >�}��NrU*�g{�
4p������z����뇄���C����C����UeW��C23-����p�3��4��������PWJKa�)r�����Y�υ׹db���u{}07K���ӝ�_�S��F�~c�x\H\���hR��/\;����/R�[Jr.6Y�^�#�_Y�טg��[�`"%[���(�b|�}���\)}��a�ya�2ܷ0����g9�e�߸�K��
���k�g������䫏� |���SW7������C��g���C�ʫ9}�A��b���f���B��n���;�;W�n[>��uΓ�Ak/y�3F���K�ŗ�ǪE��b�_Q�����S�X}J*J���(mp�c��\<��=<~�<���u-����즘�+�ji"�5������u6q�-���U~�TcZ��R�BĳZw%a�m��|5C�:��KU|�Á��
;��w��Ӏ��m��{d}d�����!�ׄ�_kۺo��Lx�x��c��o�+I>����2T�#���!Yp���^���`�+�@[���S�M3��+�K�inf�V�a"�p���{�����_Y,����P�x���<뺺��jf��Vʸ�{ڹR+�9��H��cjo+��cb%�y�������C:�?Gɴ7â�0����X�]~��3<���Q߶�o>R׹m`���@���G3`ݦz�W��EKF��@��������<�+�>�W��8;�y���}'��o2�K��K��|���i��?,RƠ��_qn� �9�0��;�Mx����^�毁n���tߙ�U]���ͷ^��	�X��ȷǃ$kD���"[��x}�u���G����yu���`̪�^~���=��tV�Jg��"ƺz�}L�����P��*�NHm<yQ��;�mv��u]h�������{�]�xeCz_�����)�:T�~���+��	�yt0�8c�fbFA�_�)J��p|ҁ�2�P{��w�e����^'��KZT�(=�{G�a�q�4\�U�H0��y+��>#�p:	�_W�2�\��J�z�4q[uȬ:����Z���w�=���T<k��,�ˮ(���y�����ILefv���ե���{V�C�J�*PP`�����yK��M��gf&�^�n���+5��v�O9���ԩ�o잀M�D������,�\}əMYy�q�י��q��ћ�yZ�]�~������*�	��<�������������$��5�K�7r͸���rK�7^�؄fuf@�`�,��v6�46���'p��C^�K�]W�{m���u��AJy����Ӽ;Q놀_�;��|>�����6��7�u���
�ȡ���,�p����#�m��
Z����#�V(k�d�x�^>w�:������]�X�S��:��0efĭ s��u0XCO�5��x��֟��,�T���̂���z���{��0����P� n�����jL�2��4Ƿ�C��+��0{�|o�m	L��'�^����?Uz��?���і��Լ(5a�8�kV],.,��?z���c��8Z5�3���'��D��8�t|�+��Q���~3;.��O�đ�L��{���ey���A�o�׆��qy�ꏂ��+)��Ϧ1l��Z�ިbW��=U�1p�1�d<��&넾����o�b��s�=^��P��Q�}���ݢ`|x�o���mL�4&����V���W�����.eؔF�;	�a�ă�����X�zT8�s���ui�nW��^�ΌwDo+��p�����sU����X4:��V%�!��\"�es^��]�7���@g�|�S{=��D^)
�f��F�۰�0�%s7���iւ+�ECk����ya�
��_ZpgE'":��/��hJ�I����P��y��ph���v�-�;��}��|69�nFv�ֿ߳S�Z�j�
~j�.�<fS+�@��A�uB�4�7x@N�3�`�<��{j�µu5[�-w/�w���=~St��יZj	(D��O��`�J�ċ�%�?V��)�ô8��f���	��5�S�����P�S�Vf��c���F��93G�t ��CM,^<�]�g��5F�	Wk��%�h�nz�z�[�N�|���]y$��L&�����/Uz걾:��<
S��2®d�_/"�?Xdl8�^ݟX�+�ĬP(��`1�L�B�u�F�x7���9�xjt�߅J˹<=[ X�[ȃN�¦WS����ȩ�h��ơ�~�J4f�����v�lˇ�Mx�j��.M$�=�@,����T<׈b����V)�i�Zs��6;N+گ��X�D�R�eyw�����G�:⛧�S�V�x ���N42�M�"�2��{2�wO���MN�]a�/
A׍��W�W�{-��x@}���"�i�ϝ<P�L,{�zzs�R)�WX�e�|��X�۞9�"���e�F�^R�j�ѵ�ݿ�K����U��Ly���9�G�w�oEs�+�yz�e�Y�'B�a��l����-�@-	�/e>ݖ�%�I��=�h8�ﾯ���g��{�<-$�9��5��ֺ���v�2����{�@���J�����g�Ј3�!��*f͘
�,-��E����k&&c�O�����,�otX��%���)��}_�bvu���[vO��S�,�u��\����&�)�aa��V�� ��p?���2�s��~���b���r��řr�e	o�C�+��x�+�Ii�x*`:�Ͼ>�(-����׻�z�g�w/�C���������]��e�!ȺeC�uP���z��*���m�d�/n4v��{��_o�Y�>Ɇ�z����D:�|gz�֞�uy��n>V8k�$���Rp:�^��T���y�L&����?	�ژ|-��Z�x}t���y�6*r웵��e�aqBW�z�ʐ�s��i�w�c�_x�%@-�����~a�A�����'7{����B8ѧ�n�����?A�Ц0y�o	�����{1�nʲ�3���ZsŇ�Y�>���a�e@m�Pҷbiٻ���{* �Ugy⾛76A��S��>�P9��@]�4�=wzT�i?��x��Q���	;h3Q>4�M���7�汣ċY��`�N\�$���&%b�Q��:�$9�;��ۗ��	���~��֝�\�+&q�+�����V��P9x�J�s�j�9íм�Ҡ��6�����@�k��QT�m9iInQB��k,z��{�ȡ�n�%�X����X����.�P-�ۜ�i�vƪ��Z�1c]��bG�0Q\��ذQ�N�6��*
�Df�e�Y/=��Vt7I��rХW���B�+5�Pu�ܰ5�A0���ؗ�M�mK?l:Ff��Wr�B� r��D��]f�BT|Q��weʰ«��u���L��^�򝱞���6�q�l�	[����"&sz���,��-���S��ذC>����¤�W�_q��s{r���vqz6=��E�V�eH>=݃5
�j=%\sO����q�z���gQ�bo\��h����:���	Ge���Nw�_v�G2��>^�&$J�:n�N�C/A5�{/h�]l����6�"&�:JrOu�{�j{�+��{{��]s��L���w!�C�DV�Ԗw(���Y��S>����pN����O�F)�xœ��$�+��5gRʆ�����a��I�=y\���Л�zz�DV�;�Wj�ǻE�/�&�	.W(
�%t�ɐQ�ע;����\̲�O4qҧ�w=�i���R���병��Xx�=�)�dh�(o`��^�oH���y�<�$�U�a�ă��S����`��T$q<e�PU>��qHQ�	I��T�<*�#��g��$1�*"|<j��V����L���L�<���{��������\���HHc���^`I/�Uj 5	j=,a+�Q^!�>7$����Y��lƬG���"ƀ�0F�'��L�~<i�ː��1O�9��w5}6)5L�2�����$!7 �xx�]��\~/*ª�<�1�g.!�1�����p;�XcVA���W2:͖!��v[�-@�W�IK�ox,�5<,[C0)ڊ��8�
���ycp�Tf�C��X>eu���Nn�ޫ�y��I����Oj�I�%;����-
���I÷fBe �PdE(D��j��O$���vM壋���f$~g����}OOs� 6���y�l�Pv8�<Z��gSɼ�E��-��U��4��C �[G���e�ǅov�oU.Ь��*�N��U�7�j�̺{�����gVd���ᮕ�F0�X�ƺ�Ꮮ�~�J�0 p�Y���y
��{�Gr�(�Ҝ�
<�;)4&y��+Ҧ�Y�ͰESL�*��"��*�X��lc���mTcA�aXUJ�Tm��ث��DX��(**��"(�Ă�3j��-J���
%AdAAQ%����(�0�"8�ue"�U���U��J����X)�(�m*�EUX��(®�Ȣi(��n0X������QY1K!X��騚���#��(��chV
�F01��c[�*��b�%�Jʢ)��ȣ"�J��5�*1�ڱ`��*�֎R�G6�
��B�EcbR��Պ
�b�\�����J����T�b�1j(��U�l+DU,�X�*��F�Q�V1j��iETQU"���
���-b�ZRČD�R,1��X�����3�|�9��Զ�/��[Z����%g5򙑚�up���b���2=���5`t�n˄
��պh<��,vf�����|ߜN���G�{p�w8�.���#�!� �RN��֥�^�o�}V�N�y�����*��VP������~bĭ M$Q����4.�O�[�&���Jz�%��@�B��F|a;���C �kN���sׅ��g�p��jR���o��LE�כ���ٓp��X�X_xf�%x��jݯ��ȨS�_�Pw����#P�p��[~��ޫ�k�&�~��3��U^����vLߥ߹n��B^����L�W't�d����~�0�g���ɋ��g,������+�K��ܪf�8��0}�j��`���f�	0��7�`��I��jqk_q|ɐ��9�E�
5��.�֫4��v�n{e�j���%bL1Ѻ��	��xA��=�h���Ǟ�4��,��u�f����=3�l�tVm�c���.��r\�g���|O����N]g/�;ǣ���48�	O>�D�^�A`BY� �O�mv�>��W=�n�.�~��5E8�[�4�������?A0}��4.�W�>�g5��BB�#^+s��]��)�k]Oja�A�%b�č�+5�����֤0s;j����g-M_=�[��=&;ݖ�n��ɺ�y�Hq��ס��9��(��1�J൪���}.؝�Z������r'�V�/�(�\2��%O���g5�C����#�Onc��Ŭ�]n�������| ���p9��.M:7U�w���9k�az\<z/`�d� a�ǆ��85s'���_�Ũ�5�=6pVx�C;P:�w�
�
0�a�d��a�C���2X0��o9꼏s�{�,+f���OR����]AC8�[��R\,J){ðBhW*��z[y�$ةfz�"��G�����0��4��u���Ez��D
n��VL�Hxt��n��Oi��y7TyV�}f/
ȡG��w+��b����Y�H���!��/۞&�fn�TV@����ޚn���R��K��ϓ��Je��ac�V�=c�Ē����R�B��޵�"��=��R^
��g��%5���5��
�G��GU�]\U�zw�s�ԣ:^�0�N���P�g�Ԋ�f�����^��t�겧�4#�{de�%�ݰ���]�κt=��]m�����q���U�}�d/A����}:d�)Uvfb�W˪�2L���LᝮƑ�*M����/Z8�7��ذ7�����c����]⣾.�����T>q�f�~�*%�K=�L�^g�A^�MVؖ�`,~����s����y)�~9��`���˫3�*�9�v�  >�ݾ�_E(���j��VsΛ��/E3����C���^�.�\3����ʬ�7�X�>���{Kv�����uq�l�KQ�F����\M�t�k�C|��fo���*�j���kv�t��г
�0��'C؃>����z6�&oҶ'�jF�����$�KY/soG�T�A2.AzT/��FPU�^�0c��j��Ǹ$��C��~�̋b{�l^ί4&�\#f��3��zT����ap0OT��g�ey8c�3�2q߫��E�I����o?�p���b%��d�8��r����7|�ma�OS�K:<M^7І�Y�/��n�o��U�y��~^h{EfД�N���Y���ktv
i��K������\�pʫ�x.�&�<�|�7�?����e�wԲ���ě���}L]��t��Wew��U�y��7�TY�ٱ.�.��N�n�+�E
�.�}�n���C���]�3��;���V"}tj�uf���t�)�cK���rc��i�~%.��N�k-=�pt��m������v�4CҐ�M����#�S/��4��q��јkK
�����˫�#�w���
c]&p2�k�����X�!����Y/��5ݕ�t�uI$�ƈ��_�e��\��M��� l~�#15�Z���&7(._��a��J�����h�"�.zXK�iOOs�s��A��j�p�q�W�P	e���א/"@�]*�Xr�C�C�������&-�����}>��&�����a��~�S��� >0y���R�SŁ%36� *�g��U�*�X�Y�����g��-m�A�g�P�Î���D��Q`�#�������C��y����}бJ�6F%sU��J�\�ʹe�xs=~��r<|I��֣F����41���)���M�N.f�)������B�ȧ�,qό�P�[R��(�Cu�&k�����a���d{�}$�j�M�SY0V�����TY����P$�/=����̱Pw�Xu�앥�qp��/��!Ȼ�y�.։)E,&Y�<Ⱥ���������}A�h�%��4D]��J�x?����	�=j�fT ��z4}Y����[�f�c`��)�>K~R���o�iZ��%���.^��F�Z��<-4�����">8��̱Q#��_��tJ�Ch|<�o=l��Rw�]�]<)���]c.ٲh�_�	qіC�u����" �|�ړ��5�K)t�ɏ�S�Wr�	!􊔼4_����t�x��9�˰rٍo��=�sGU�o����{���k��^�	�*�����9�U�`�.ۄ��ף1�~�Xm���^�j,g��IR,z$�s��^A��L`?&=Q��_�!\��0M�Ū������S��6;I�î�Ѿ|Ǟ{3U�yaꊙ|�+��R�b���x1ؖ���\����e����d1{�=JY7ꚃ=j۵S��M��[a��O.�\�b���s�±{�5n��=8�r���ϩe��8=�p�\�@�"B�:�8U��$�H���������^䙍U\����{IQ�`���w��h,�S�1��qXc�L�R|}��]A���O��{��~��m��n+V=���A��xB�٩\±s�x���fz�G�_�#��o�[������=#=�����[�.�̃o� #�3[��{��y,h;������7�F/]���>��#���X*�e�7�ow�<�9�6��~��C��)�t�+]ezO63kٵ��u�V蚰�{Ҵ�	+�<��V<�+���npw��z�G�Tч��I�����r5{IV�h�,��~��?w8U�+H%_,�>�0�s�(Ί	�sjs���k��0M�V�޹/�B"y�5q�4��������W���ϴ�Q�<4���a�1��rm+(Nww�Ёؠ���i���|�B�'ݝ�{w����b��,�SYF��$i��F6��:���f�^PA�~_}��}�����37O����յ��أ*�-3]h2�cٰ��G�<��e���}������T�{��U;�Yϧ�.ݦ��5^^E<{�.��R�.z�w�1mק��Hӳ�{Z.�k|��*��S3�%�(S~����|s�=��V&��vΐ˵�6�����^�Փ��3�rW�{��k��E�WS�i\���C����i������PۮEs��#cW�g���m��냂qX��<�S�qX/3����X[/�zg��9�.+��M�g/T�g:�5��=��~���C
����+�A�En{*�+z�v�MTn�]1����0,+{�D=�\*W�;��4ӊ�w
6*�Q<����S;�Ķ�DA�״��,����%�ҽʰWA�Z�1�}��=<���ɏ6h6�����zǨ<=�|�7EH�J�xp��Dԡ�7���X�ᏼ=�w�����#u-���B����h_j�ɮ�G	k��}�N�r�B��}����[�8gd����!��}���@�z�{4���ӐY�<�z:.�����
��e�2��oz���p�{ 6���>�N����LZ��������z��?v<Q��q7�k�F���Y��jǥ��mч�T���=�K({|+qB2�:��FJ�^�ڜ��E�b8�R�TJ�XYӓ��ƳH�=\gU�]�s��5�#}��ͭ{��om#�Y؅7� 65cQ`���a�����ö�����:�yl9�N�/�6�)�:��zM�k����g�P��p�ؘ���2�D�ޱ:�����X����2��'�<Vr_�iٞ�ͤ�J}��㣷��b⟆�B�My�g��Arf���'y�N�a��k��t��J��a��䙽��tΛ��YE��j��];ӏs[�*���uqfĞ�89�qY�
�0��'Cߢ����zm�PR�^�}���|�{{zCx�x�[,^�(�������P��y���¡(:<� �ᩍ�]�)���ݼ��&�i�x��[;��\#���!���<�j���f��L�{=|-y=~�⌖X��/EA*ս��Қ�9*��ա��wԠrX�P�=\�B�����H��빐���!��c0��{.\$�YF��8�xeg#�#�nD{t]:w$�]nU���X��֛[W�98�V�R���D�=Mˀ����f�l�,܉�]��/;�(��ݍ�E��h5�m������:���N�����z��t#�	����puV:<N�8�y.5_QΘ�<m[S=��%Qƈ@ϱB��X��[J�זnG��<4,�wax:�X�'���4����C��Q�lE��M���j�1V}��ޡ7�muf�Ճջp�҃4۸�S@�|�^�ɻ�|筲����S����4��H�il|�]���λ\�:m=��{\�ܚY�n�;w1�RcP-?AH�,Ĩ>5+�J4f���o���ne^�Z�x�g��p��옴Kl{5��_���w^�����)J��P�>���@ـ4���-Ǻ_d��4��}�����GX[��Omß{��6��M���j�52T<��*����V�3���Gr�;�P6h�ڲ3��Y�/�����������(b�.��i��t��]�������`��;^�r�_�[C-|&e���Xp#����<�$ia��fmu�2�c�/~=Ylm�LV�hߟ��W�o�v80x��Õ�X�"�{�j^- tX��^��2Rŷ�:�b�|B�5}.��ւ��>�Yv���@篣�zRuP>��q/�v����V;P�<��'V�U�]�9��R;���R�H�l%i�5|����6�WX�k.W y�����Z���,>��������:O6䂳o��=�v�-�v0)�hL뇈�-q�5v�\��*�/����0����p���n��h���x>$S
��t�����ܟ��lȻ�c��Z�%��gi;�N��wC>������*ͳ�|�:5��S/p��3�P�^�P���%�m�׽��,��ҁﾰ�L �_��^z'ُ����u�C��M��S�ݙ�7��V���k8(D#��P�9��y��z��]���>�S��5���|m{��\�C���Kr��EI�W����ن�Qb���MG�<:�uKP��{���4����C5���օP�X�`�ŵ.yx]x�=-�'(���s:;��=��i���Z�~��oYa�ͪ~ϘPP�2�6�a�a�(����3^U#�tC���e���/ԴV��]���ȱy�g=�p��Բ���ϋ���x�G[���{,J����!�D�-4�0*���ՑC�,�l�og�MHQ��ղ���Ll��42��<z�yF#
��:@гW~]|^��fl��g��6���V�cJ+���a�Q��O3ڸ��ðJ���B"ꙴ����j�'Z�p�[���3���4�����l=Ή��k�-�6�_h��k�Y�������8���i��K-����"���a���)f���XyV�*�w�(ck�R�0₃�ؽ��+0��w�Qƅ�;�{oU��[s��h8}�g 4/"��}o�
7��v�ևi���:�Kʁ�Ι� ��[�kN	+H{�0ۮ��_�v���(����]Al���h�|�O�P:�t)�ׂ�����ɫ�f����b��o_ޮ�¼�L��_�G��۞}1�}A�o|�]���8��$���ʱ��k���rٝ+��ڄ�6�EQV,��ͭG`����o�pb�%_Vb�ƕX��,��hv���jݾ7s�;%����amW:�n�~�P�T�x���'���K'��dS�3R凴A�������θ8x><;AzV��Ծ_J�K��{�u�p��^��d�����(N�Ӹ<]��b���Y�8f��f�k��K<�(`SiK��p�%�Xܕ�wG�N{������1�{߭=�ʕ㧌8|3��Ϯ;��r�V$_���Խ���j�E�Q�
1<ӈh�=/�����f��Ʒx�]L�um�&�.W�J���%�@o�k����'<٬2��(}Chv���d*� �w����o�����٠�Bʚ�qu�H� ��;���-�Ӂ���w"Hލ	�"3I=�_���ո�oA6
7�J�t��qC�����ۣ���� ɛ���*��H/��Z9N��h*I�{�L?A�'7�u/�h؂��S�`��C]sn+n����Kta1�I�Gq�`�	��Ź��t���gf�&�	�W`T��y�X�(P��!��$������B��=����&�6<}x#�*�k[��Y�)�a�^O�|��n%���D�C(�1;4���x�z,�a}+�g\r��(��;a�R��E!b���{�l�J�b��1vR�S]�!%��x��ˍ��z����3�9yN�}x�0vG<��ܩ4�X�eW�t1,�t7��{�3�bSժ糰��H��#�NL�����OWUpg�K58]�Ք-�Xb��|�!�lE��ٝ�J\���W��n��5A��#�e�G��(h�z���XX:��C�U�%?>�]^!�T�t(sr����<k�h������.?@Ճ��
@	��S�Ի2�Z;=��44C<��̢e�u��n��O�J��:٤#�>�1v�0�v}.���tZ���:��W&�0D��V��|���Ñ)�$�C����S��ھO*�kH��b��i���G-�c�y$\f�Oz��|�aCI.F��.X����pHN��Σ�!ʜ1�!]�إ(&����-����}��H8Qo��A�vf��Z�����dr��
�v�cl�Z'e�RK}����X����L���,�E;/g�5.n��1�]�x>4xc{�2�NZ�x�Q5-����IV%�v\�P8���������|oJ�*|]\�6��'�+�V.�:Y��JR�6��>�{GD�z0On5�s����ї�Z�mЂVG%\����X~���(��0â�္��Y���55�f�̝R���p�XJM��V>�%��E5ʮo16<T���7Ke7��t9�4��Z�s^o*D
�g+`�,���m3Y����ۭ�i����B��_*���`�(syv���.Ͱ�y�5��ygK��J�Ⱥݞ�1��<.��~��*��Y/[��@��X�@m^��׾�9���5Cץ"���.���Ն�j&Py<xo����=�j���s���+:!Zx=�t�Z�X��^��v!����fw��g��{B�ge-˨v�ݲg|�o�����u
m��u�n���~�}��<ӶΧ�k֫.2G��x��WV�E�]0T8��]���S_
*���.�t�]kq�=��D�x��t��0���!�.�����$��$���\��fkx^�ß�]c��(*��������3�?Z��Q�[Q!iAX�V
,D-%��<��D�&)Z���S-F�,�*�m��UX��،[e
��b�TDX*�űR,Eb�c���*�X��#P���DH�UP��W-Q\Т��+�1��ELk"��E�kb��
hTTPU�+E ��\�+��&���E"���""��e.��1�T���@F,Dqi��[�X��6�Ve���u��A�
�U"�Q�-C�+4�Af1�EUQQQb�PRYY�b��TTXb�T
E�X���ib�Dj@U�X�VύlR�.Gt�|�m^�]!��˵{^�Hr}Ӟ�`C�{-n�`�v��5_l�,41K�
ek:k�<��-���� �����f�G���>ė���^�;��=G�=Ki>��R�
�S���7��_���@��8.��eS%���ւ*�>v����\�,'������Ԫ:���}.��:ߑ���DwѸ� }Uqj.�S~�R�|�l��s���
E���11�H,�ř�&�{Z�2Ht��衦�`��R�r��Go�?ģ���!�w�Y]u�QmM�G�޷o����R�(��TJ�40ץ�tܣ&=|f����e֠�+�܁�mɏ\|��{<����������Ϝ���%i�ǎk�Y�WJw����ˬ�s�w��űMI��uk�u�>�~�(f���e�X؃Jˋ"{��-�c��*�}S3�^�vA���z�o4غ���\j�a�,��~]��~}��Wo�/8i������E�O%d��=]4"ύ��m���D˜6,��1/4,�\_����w�6�ڪ���φԉ��M������a��`.���_����t�8�q/x.���$w����	�H-�R�/ОP���x��Ay9��Gm��л���Xw��2�J���M�6yGЃ�uï�S�j�l	��|(�F�7g����Z&�[Cl�Q$����i�]��J�F4δ�
l��v��kLM=ߪ���}���ަ�7y�f���	��,�ө����ߖW_��k���D�V�������c��g����l̋����z�O;�hj����a`�,�wĜ��]�S�'�7����4ԉU�):W���^�M~�F���l	~���"��ϫ�V%�&��/S�=�~^8�ڿA���ah�TX� ��skQ�������{��Ί�=^ƀ��槙Y<yywG��V��G�Դ�U=M���
�C^����x}t���-k�/���i�a~������\K>��K��(sq��ҮV���@�gt�j*#��nm��d��³�W|
��$���3V)�����~�k��]5�38Q��C�ɢ?s�\�a�0gR�{ꔪ�A����ơ�u"J�ѳ��K��������9ݛ�"p���������˾9�L_���4�y�-�J4f�d�x�z\��h�����ܚ>�Ó�U5{Dˇ�m��n�@�t�;��X�r�5��FFP�4�R�&%�)�`t �3���K��ٝ���FWsz���Y��MޤS{�wM�'>��������O����b��/�О���G��0��nvm:t�.�hPVvJ�U�
�K{�{E��$h|�����ɵd�C��=��cX�8�������9$�bQ���~�8�;������8'ށf^�~�=Vlx�G����8��	��y���ϩ��j�c^��H����
�4����X�[���c}P�p{��W��,��ڛ΋z��ט����8�0vb�W>_���]ْ�{u|�*��i�f�����8���?;f-�kH����<�_���rɇ��r��d>���tO
�3[���=���>ը���%ᮡ٢[0��p�Cܤ��[n�	����,
�fl�{WFv�ٵe������d�pgD�Z53�+G�X��ῧ��1�ǭ?'��J�v�޾P!�X������|X�:�ͳ�R,h�Ml>��u���y�l�=m����9����N�1F�L��i9��]�r���'O&5��p˻hWg|�z�j���t���XV�7x�|���X"��P��;��,R���sꄻ���#]˝��x��t��zz�K��:��҇S�z��*B��c��j��|2V�ٚv�^W��`�fg��LN����f�G�sǆ,H^��)�炑[H��Ι���)��� �J_AF�P[�e����.�g[8+9�� ����K�Ci`���lʝɊH���㖧e �����n���N�0&�t�W��]�S�9��.���ﾯEOxo�8�6
�]=�,F��lbep��Z�y��*�ٴ���wY�����1��nv��l��(^��L�(&���5p�e�WO�̛�u*ۡ˨\�pF��"����0����;���Sܪ �#�����oYixוL�o�2C�p��嶺�7���w�9A���Q=Y�L��)��~��r�[>?��������8tOb$eo���Oᜪ���(X��۬:EPsVQ���^�Wf��(<�pu�G�1�c�-�9����E�e�����=bK�� B�5[�{����tQ�=�ㆎ�R���S��

ם*ّgbT+�����B�|�L��ZӂJ�,=�~W�^��X<�.6 н<�[���Kخ���2� F�ԅ}�u�ޗ�=�w�u����MX�GX��^����ϥR���c��6�4|$b��ZI���XG]�!��s����lT{k���^��M�h�|�r�ʿ7�{2����q=1T��}u��߾�`ј�ll}X�&�}�����~���Xg����[�4������,�ݥNk��_Y7){�-��۩�ml�U�����2�X��{�eg.m�pL���ew4�&���͒bA����7�M����M)���	�3�Xv�p�ٯ���������ك}�f��5��̕NU@a��
�s�Us^Dw�Y�xo�T'�Mh�Qz{^����rJĵ��B����bcC�O�ե=+���R��}�u�;"�^g0j��>����<��^�C~6H����k�����3��/~H��;ܠ|s���i��S�_��.���(s:�C���k���p��Ԣ�����u�6.;��n�V$s�[������+}�Ju������5�ø�:����vj�(��^��6�Z�]6T��2�o9۝Q_�@�t�D�L�ִJﭣ��++ڢ��{��^]WP�'m��a����L�heP����.��~��L>h6[��ߔ���!��+0&/��N�]��z�+�����e��E@6��
�$T�J+*���`��\����V�r���03v�5}Cvү����a�|��}�f���r�W$V4��*�nQ��3MS�T�4��oӺ���@s7�P�Jx�E�Yj�V�|�_uKTmʉ\XYӓ����DZ<�L7~����N��P�~<)�ˏl��Uwk~�����T}�g_M�"���5�¦�����JI�UVkY���'/ڇ{&s��8�emI\:M!Q�0O���f��O��k�a5�h:��lK�}ܤS�ȸ���V�LǪ��sCyS=���W;�3��+�30��T��m���y�X\9���a�aqd^޶v�"��q�~���,X���Ei����r�ܰ�i���@�(Iå��kL��x<��eSfNN�z*���}V��#n��P�mI����f���+�4m���Z�u�pV�b�Pī}C���^u�G��]]���k쇴'ɛ8����At�3L?j>�r�������<�L޾$�0����ײC=���'�֘��tK��D��c����+��a�v4}��Uq�3���� �ɏ%gR�d��v�bء��n���[.���V:g�*�P��~����;���-'�������b\v��Vg`t��p��<����~C�Nc=ᖣDw��GE�4(�}>�U.��0x賁xSV���3�ѭ��I��uƱW�����$[��E���}	ڡ��'۞���>P��rYR�Լ]����+�&��k|���%;<���s�*�Uq�5�x,�P��)�*��U����P��v��r_����4!�=�EyJ9�GZ��������9�lԢ��g#�#����#>�,囚#��P��	���&a�����ʶ�C����Z��7��1�"�=/Fd����@߶;>������r=�.�"Q(����PK@��yn��-:77]�"�����=�bNa���_|�8~�_��XkIW���Z�䰕r��6:隿��x&�9�&m�'R�b	����Z��mKU�ݢ��J�� <k�*o�CJ�E|m��I`�lQJ���{'�x�r,��.���W#~��=O�T<Vz�g�ؼu����:YM�VX�wF�#HtY]�ķ�z�n��۾�f@|�z�/�P�����w���G<�iҜ��kAV������c��1�2x&Ͼ���U��Ub��,t��(�A���7+�^��Lk�q��e���ۯmB�������n�W�We�G|����][�<3�I���׋l�V�W�%<P����W�_���]��g�h#�z��lGF���u�w�^�9�	������pu��룽����Ώ�Ϻ�a�7�k|�L�<Ve�{�\�Ig�
�^Q�;0*��m+�P���a�L���+��fܱ��ƛ��r~�9ʞ�ff3O��T�>���vC9Y��g�j�2�W�{��r�V�7~������w2�2�8�*e�o(B�M�F��A�OQ�J͵޾�0�����(����bU���-	[�J���CWS�j�[��	ܓl��	�3ݷ鉧�4Wr�%\��Lmb��A�.A�M��݈��k�ݨ��O�A+h8���W���������~�KMN�PR����p�������G��&���ů�U�p�"~��K˫//�fz�y-!ސ[él�-�����v����hv-Ժ.L��X�W��O�H4ij��4�-��^�-D�u�Z��L�y/+�4�Boڪ_��:�p�Xt{�/�7��^�8=��Sՠ�+d�8q�Ջ̀v��ubx���Z4�r����6���ح�{4��*frς���-�hXyp�ӳi��8�~B�����NK�5׶�Kw�3W�s�Q�>
h��0�i�3��K��Z���5%�c���O���5+�D�=��z��ʶ�J��b*�ᕗw���\YȐ�ނ�!�S�E��T�rzYu�nz�%ޝFX�u~���tv����Y�^>�Rws�Ș���uzn����y��w׾���6):-�K�.�^��A\�B�Q�xz�������Va�M4{$;7�ކ�s�I�V-���W'δƥ*�(a�<���9�m׶ B��͌Q�B��;F�c�K��ۡ��ɪ'ќ�ct�9ۓ���p��jާ�.�{�c���_4��	�Bg�	������{�OlE�����{��c5v���AY�����1V*�b��l�R�ɠ��އJؼ�|����f���h7����t�����i���;2��K1uq��,/δ��خ}%����(�]q��"���C���V�z�睊Ř�nm E�p�y���0�>�=�w/C�r�k1��X���xo�x��߄��I�l�ڴ�;Sex>3]/�ɐ��:y灵{�I�*s*��@�P��m�G�<͉�>fBϼ7ɥ��<u�j8��'1�ߐ]���P�a����3��Y�P���lI��|%��n��+)����^�ey�����q(�n�%����g��6u�fU�U���1|��{��U>]�������γ �0����3����>���xJy��G�e�^m >t:�{�����߻�>�v��Դw��4r�s�M�^�i�f5F.W.��,�7��_��;W���z.$�o]{�v���>�N��^%�ʷ[����	�X�J��$���Uu��"�U�P�0�:��"�G�ў68:����=��*��C͚}V("��P�&���k4C��IS�w�DRb;��\s��hk�8�*������u�sz���d"��<yt�%�gA�a�*�NIf�mQt���r�\'Sy������ �i��dZ�]����*vs��/ҕ�ɮ����0��"������#�W�'6��E��ܲ]���}L]�XV���.+���P{���*���gF����ra�v���〮[Cl R�
 w����-\6����.5�6ўti{���vD�c�C������TD����|�D�3C_��j�{h�&6�e��~댞��翟ꊗ���~U�C�ۿ�P�j�"���iv����O� �j ã��Jm/�4�ߐO���bw�'�r��Cg�\��^5R����α�X.�V����V��~逵�knz�5��=�-��9{T�d�`�ܴ�)�MˠX����r�f/V�e��T��b2�oQ��f��kf;���u��}\�o�������Vs�B{�q%(9�����ˑ͐,O�hq�=\\ڇy?.,jz��av*Xo��P���.v��9]��#�o{'ue����%�X�=�Dִ����gD��Xa^�ާcAu�bo�$�1�y�[���CE���l���;������G��9|;![
��\0��{]��3Č���^�y̋̉�/����i��cma�	�pϬ�זbw/ky*n��E]Յ�TxЀ���t�[Q�^���bec�A��K9I�\m��dw�&V�1�q`�ۛ�{w3�%=5�h:��/C��0,A|{��.�ڒ��8ІB3���Z��v����;4��܊nc���-'}���+��A��k��SV��ӈ�K�v͵1g�ۮg�עkl>�O��B���;#Hq��mgkX�(<z*f���eq��{�2�K����co�$�����ԗW-�,��&�@�T��Z�V�����N�^����#�S�&'���&vh���CoMp��W1*��5W��r
֎YLCھ�������e�l�/�
;���<��l��x�DJO���[�}h�w
͖8��Ah��1�����e�N.�u���3۵�{���:�3OP���r6�����)���h�e9t�Y'=eGW�\|�bk^��S�r�£�ά�\�FSTe;���c����u{A/9��u�/�h�F�06����et'7K�枹����fۓ��۵4�ѹ�x�ox^�Fb�͔����=e[���kD�Ov��g]Ε|�	�@`�uA�P��N�~��{ӏ[�B6��W�U�ac]�T�:Guh7\�P�eJ�YQl;�8�/\��ú��de�U]^�B{���+����K��jc\���櫕Sa����q;8��e�R5�������a1�OjL�O_L�ta���� wZ�7�4�s!�������Nմ&\b�π��u��(Ѥ0�&�m�f�+�"�o.����#ʳ�rDE��©��$�3c.���DX��v��b�A�n+n�㾒�g}��ξgu�J�]�;6~1�A�N/b���\�I�"���gH�#��M���`�1J��vhnY����b;�.j}��A/�I	�lԻ�s,s��fҰn\��S�`/����6�}�>zI ��j�wV�e_�ՇEY�(�8A�>kV�	Vf��L��h{�q���yS����.t�!es��<��8��v�GY�O��V0�l���@[�c�U�����z�𛸪[Qkܸ���"R�`d��d����'����j��I����'3��g�a`�t5��18~�r>� ]�K��qMG��C� �#޺��z˚�}�;�l˝觕}�z�u��\&*���.\�B{��Y؆��4�6�k��pط�[*��X�*��4�2����74-�Owg���w*o�� ���>��|��g&ώ��9iJº 6�����:�T9�������V�w]�4�6�#D
�1J����P�b���/�٭B�N�,�0��+�l�F׽]*����s���D<��Ʒ���:���p�ܹ9�;j�����6���o1!ݸ'ZCRK`p�%;�im�Q�!F���s(�l���E�,�f:aZ�d�[u�:�ɀ���(��;��vy��NUd���M�Ǜ'kF�H��?��"�>j$�)q�eB��5�J��Tr�fS1����%�E�(�dVQY�eI�`\YmRUB�E���.5b�ˌQH�B�YJť�`�Z�J��U��"�F�+5���k"�����j��Z�V��J�SF1�*Uke�V��b%V-�6�2ڥii-ce-�Zmm��l�c[F��U�kTm�Tm�f�U�V�L!P�]4qKY,J��*���Um*V`[CV\R��֭��QXҕ�رV�5��ZR��%B��aF����[R�ҍ����%)b�V4�L⩆ډj\5�Z�jU�Z�j-�m���-UEZ5�+k�U�V���Z�kT�Jʖ���L�)kDJ�am�h�XR��	��?(�;����S+��q��۷��z���/nk���'�^=н!W�r�}�tg���ǰ�u�3�ֳX��ۻ~��g7Ӹ��I�4��d�-�3۪�+��u\LW����nmvz�SwF1<�����s
���+3�&hd��TP�����0���8Z���^Ϫ��ծP�I�;M��<��\�S��ut�K��+��U�����Cl�^\�>K@*/Gh3���ƅyc���;�W<���th9Y��~U�ʄ n�qJAV'��J�fu�����H:ɿ^z���^2���nWh�A�;���]ʺK��"P��{jt�+��X�U�(Z���	��p��*0w7�W�A}�����c�[j�*R�@x���9�PұP�)��{KEC� ]���o���IT&߾K����-��3�y�{�2��ʶ�q_>�B�q.Q���3��v<�q�6֠b�֋�=Ylv|�/*���t�~����X+�1�|�-b�+r±�1e�{�}M#d�H�[;d�Vz�A׏��0��ˍb�^{nr��0�%���8񃮯�d���oM���V=u�W�ۭ � ����+�Qش����ܫ7r.�Ai�󊈫�f�-�J r�Pk�`�B�r������n��RJ��#�?i��Q��!y+x���^ɓ7Z�fՆoR!�gC�q�����{��Vi�.dK��qP�M�=���P�[�A�@��N�>=Z��9Y=��_'·J���������6,u�9w�_���θłvx��S;`O8�����<W�p���^�N٪��d��{H��1�7<��
��oTJ���Kf[��F�mTr�mgb`�w�b�	�u�^z���5�w��n�C�8��E���W���f�l�s�y���K�+��?.Zn�-?o��@�����*��tVtb��_�n�gg�Luz�y+��<��f�#�c�����ײ0��r���9-E�`���χUC��V�bR,h�Ml>áց��0� ��q7ކz#y\�͏8��]6���J�?�z��\�;��%�+��{2��!ݽ+,�=��K��<�ٍ��ꁡ�W�P�L׹dP�G<E�1��BĹŁ�٥�ԁ p��_�wb��w����΄*�u��%�A�^��-�eb�Bݟ7��
��dP쾝�7Z>3׀�NL�<H��=�-��L�hg&0s3�k�T�����&u�zb�8�rv^�txU�'�d�Vz�h�����o��e�WO�̛�ԫlr�n�b��)�լ�-�ŗ��ʘ\�(����]8*����U�_ekو�:D�:�[.�����__�5��^�m)\_Vf����i򀻭���;r�!��8���(O�`������n���d�h�Π`�VQ�ڇCn����g��f�s+�<����On�}�.���:�*�ț��uA����f���t%���R����(�� ��Zi~��C�0�Y�
�^U�r��h�#�/LXZ��l6�W�w�*�bC@�J��5I8,�P�˅_��j��Y��ye��Yii��eP&�d�=���|t;�ڀz����_Im!o�M��"�9�(�	�U������֝��]�W��HFDu�C/�޸-;��#�պC��ߦ3/�R�\v4À=������'a(Яxf�/�`�f�u�������/n�lv�P?lLo����zcR����#������)�ە8m�X�܋����K �H-�r�3�n�ۭdЫ�k��}�y��S0�l�pIX��//4���z9���mK�+��1L��߄��	<-��V�G^�eX����,W���¬�� uy.�d廘hc<���Y#���H���܂^�p�ϧ��!��}����]ۍR�XU^����U3�8��"[|x}�������W�>�o���C$<�^�$�>�i�ya�`�bcD�+ܫ�P|%|��ﴢ��7\D����ة��sx��4k�%j8:l�u3�&��J2���Y,�w��l���#�R��Lr�(��;���@�[�7.�n���[�;.��̟��]�����2p~m�-V����_p��ť���/�|�=D�
�f��� �K�{�y��V3`2"�WY���Ǭ��}L3^�T������@k��S@��Nu�>��I�&�Cq��D4�g=5�ҍ��jLe��w}���9`�7��W
z����Y+�P춹pi���G��g.z�*B�Tp��Җe�D`�YJ��ś��^}�	��߼�w�]�F�
RmV��khЎ��S�)x
b�LVyM�Q⼲�|��1�7u�&7`�x�s�����ڴ����c�`L?�k ��6� )����X
0�����)�}��h��{,����Z�	�_�x�]�	L���;�ˉ��x+}`��C�������ylr�#�$��x{�]�K�Է"Ƭ��ӑA�0�uKTv(�Eǭ]9�Re䗖�zsy+�zw��	��ﺚ�ޠ�3��z�l�s���S5(*���Ϻ��`�XfMw5�R�mZ�w�ɽ��Wm;�zVTz���^�p!~�pu�P}��Ugp;�q�rI�h�ԯ�S�.�k�zZܼ�l4C=v2b;(�j>�[8�|����W�{o=�{hO��
y�s
â����8�-�����]�e~��HW�ז.��2�M�~��\f��,�7kΘ�s�F���Vw.��uw	0�L����"��*YQr�}U��w����7���s��C2V�n�밽�K�Mt�oU�Ⱶޕpz���X�D�[��O(%�|]Ǘ�w�ҍ2Į2��}��dg)�O:��i�"��h8^��C�.�x�Ou�bG�3e��%�8R�C��/���eΦY�)˭�+��������s���8�%=�R�g]��UqkI���d>�>�R���G�^��v�%/��&w{��+P_yk��K�!��\z뱭�R��^}7�JR{^�4,�i=^��X5A�ʹ�9^�[9`��E����0�ڬZ<#�[�{�F�K��r��y^\�ވ�Uz�ϝߍ�C�1%�ϔ3킹+r��-*/�>�5�ǕüO���FI��;�ih��,Pr���Z>o2*��N�W�LX�J����d������,��_���L�Ɔ����c(�5����4@��.C�������	�z��R�}6f�>������8U�k�ݢ˭u)U� <h)P�iX�a�L�٥���۷��|7&Q�Xkլ�a�n"�)��Պn�6��Sٮ�I_
����E���/dW�]x�܌:9�zWnj�4' ��0�O���+�¾��מ#���ri�#$p�fb�� k���/#�	ld�ii9o/��>���S`ʽ�F���E�/b�~]�z���G�.�@�c�z
F�&ڱiM|��G|�u��U�#,3g���\6�f����.���=�p疑��/>z�>��v&�=^]$�R�ɮ���hD/���u�����%xp_��jn�<6��=Y�{�!.��p�'Z� P˒�,W��V;کd�v�8i�c!��^�Z�\A�C����e��pW*�Ng��׵X�L�x���\�z�+�p:EOve��rxxy4����W%<0J1��`�a+�i�=���������y��[>�}�e�"O��W�I<f�7�P��(q�Z�c]��u͖�75�8C܃�'ݒ�j�NwegEl{m�԰��Ix|5Qg���r����NPw�/ʽ���R�s�w��⼡}/�nWrA^=JII��<���3Չx`u��U"Ǝ��[��w�m���3o��V�!�z�]��c0����U���k����φz��J��<&V���F�=�״F3�V�(U�(3L),%6�iiv���+]�E��ਪnW^)~��Fr�^�w4;b*/�9���,�/t����@�u���BEJ�Yl��Z�]r�)���ME��*d�`�y���T��]��0���`�;�㍣�m�'��Uaz�u����ֻ�W���e�s�}��:�؀�ej������«qx�OWjgk:�u�Y�!'�u[������ٌr�aʇ}�U�
j�`�5�`�{i.,@��+*��h���`��g(�g�c����(�3e��V��6�nO
�\�'ً?���S�v̥��4[PЬV��}�=����a�f �U�����0v�o	�W�#��r���4����06�Օ��]�3�a������i[�
4��qp�!�P���xj[�i���/�d|={�q���kw�M{,��(
�t�����>��Y%n
E�Jt��,�U�j�"��X/vٮ%�ۗ��9}�$~��[��{��W�@r����� 5sB���+������^/R�4��m��e��J�nc{�mX��PuC��.�W���Od򶴬�'a(��Y��SB!uw�"�7��.��֜����o�72�v&��ًk�R�9%i�+�i�f�;��Et������o�vLߥ߹n��P�a� EfӅ`��\.������єG4��Tw;i��2�� ^N�nK8���c��0L�u���l��rꝭ,x;,�jY�Vq,�;#������͡�M��"<�U��/?*��|/�Ts���_ެ�M��`ZhOxo�gR�{Q#������Z+f��A�����r�֬�Q���_���P���#��bA/����n��n�����<}7	[O%@��_�<d�5���=�h�-�{�<>ۏ��C�4����94���f�@��כ���l� �N�����X���\;A}U�b��+�[,~�u/^?T�4j��<�:�땇Z�����CN�ˬ���8�M$@z�c����8$�i�g��;�e )}�Pk	���/��˗Zk���{U�M��"U�X��;}��у�h�	�eH0�AM,�TD�����}p,>���*��f�V��]�T�qZ���C�N�}���9n�T)�(�Tp���|�ˮ(����\53Y�^.#�[��̌=�����X�:|�3(��d�I����g��G����ѻ�s2�}櫼���p"[7﬐���y��`*�P�S$��4��JV����]�H��u_�4k=Yw�ο%�W���h�q�O=2�ʸ��L��~��5��꽼!�71�ݠ� |g^����}632��Iv͵��GA�Y��2p�pdˋU�:T�k1/^���w��]��+�#vt��+p�gXv^��	���w�˯u
�6�y�5I���+,r&xu�Q��U�eT	�~`szw *����On�j�$2']y�f���fh��T�ճ{>���Yi��V�0���Z��mKzd����&4A񺬁��S�3A��.߄�G�X'�X�+}a��j+�^{��Y��U�HN�ukL�g<�u��G�\>�U�B���Ӄ��L���q�ؼ ��}���B����ZS�^���xly�s|��#�|<�W�����y�a}쥰�>�,]ze>���_>6;_���Ѱ\�{֮�+|�;*c��6�����}|jgA�`|=7��]����Zz�u=
��閛ȟ��A�]%��4�l�t�����g�g����º��^ZG�S��r�R�q� ���BX���譾I������p�Ǿ����As%��R�Dz;�S+\�d�=~n�8��Q�4Š���Uު�����(���NPd?��i�������.���>Ω�x�=>�l�� ����l�86��Ö�|~܈5آ��R���bj���F��;���z=���>�����+U۹N�e�c~:/?L����S6��}����6��l8�+��2�`pͣ�`�ȅn���]�E��j�zR
BT]�����kdv�9��A�9�u}]�X����Ow�i��w��Z��W����9��#�AIb%z}L��`�K*WKQq�;A�oZ���ߒ��N��0��c�E��K�\��\�B��L��=�_%�k����v���u4�uLY�߀C�h��%��D;�I3�Q`�ˁd�,� �^x���N����x�n�A�6*�o�U�?*��O
��
�:�mC>��)�4�⡥�2�VU�W�ʻd����"��4<!�oy.��Y��N�a���d:<���������o+N��vz{fvT�uGR�M)�j4o�CJQ�|�2'���G.@�YS7���C ��0vls7}Weu=�T{^�c|xe�WhD'0�>�{BX�<�ʄj��LaX��w��Mj�'��5�@�>�b�P��>��e��9}�bL�k���c�NRR
�5��r��{�O�^�����,�޶|](xM�u�9\W�W����[�u��Z����Y���6�LX"�GMˠx�Q&���S3�������>y��[���:8����B�6�A{[յF�aL=Ro:��1WA�b�,[�{W_P��i���$P�ܼ��`�b�.-�Z>G���m@d�ܓV�����O�mʈM������S�X�f'�{W��3�eOt�_L��r����Vvw�^JJ��Ѽa���׋�w��J�q����MK*����'5p��+`Æ�;\.����q��X��K.+�u��"nu�R��=R>���_&1AҀ�,���O[��8��9r\�|�;~��N�����`���8�F�gv��z�lDQ/70�y�]J�֭���ܳ��Ǚ5�g�t�:��l��\eH���T�c.�$�z�]xiQ5(�9q%X������y���FB����{�����dD��f�ؼSe�%�&�ژ���UF;�.�țrL\���s�����Ģ\�����?uc&v��X�
��Q�������8{(��w��|�]B����]H�-aNW���8��`� o`Pu�v�aWG��CC<_��8*�c�[S�;O��'���e�ߌ��qɍ�o�:J���*��J闛ƵN�&�[�̎��,0�pQ�=��s�1����î��S�vq�N�'9�@*��`���Y�yv�4�%+�X�n3�Rx��.V�m+*����`.r<(6z�]~^sW%��o�X��޴8��g�M�^��[�s�8�$��+��kVgS�Y�ʰj#�Oc;���ױ�L�t���\�uq�˰nw�Ql��iT�ffQ�]C��څ�U���}$�E!P��4b��9�u"�X�fMb��f��<5��j���-�n"[�����^��KѸѕ*��5���$�T��T
Y9LZg1 ]�A�Ь4Ƞ���T&��
�U�`���&��
W&V�aYA��P���f��I�V����..8s�_<���7�W��}%W��%�lx{=m�G8�R�`��I�J�d��ф�"gf(��*���xFGQ�^�#YF���F$_�,_<� 5v�%x�6��i��a��1�M�p�p��AE�<�(�8�U������f�`�������(�� .!	�`we�Ю�הz ��Pj�3�>V��2y熠��N���F�/��=r�Z�mw³���K��,<��-�޼jXˀm���4�ujq��âi�*ƞ�g��p��1n��|��,��`�y����"��(ڣݴ�R�$.��ps��.��1W&��7
�Ԣ�?cZ���5aӥ��N��<2�Up��j�7�J�H+�yCȉ�7c#V�L9�غ*M�2�"��u2�R/{Z���釻L{��S5�_��+޻����#��5�%=�!�$��f'Yw�`o���5p���%���v�r\wF;�n`\�ե}Pmr�p�8��%*#�aEAp�ja���J�-k
�T�m��q�pQ�m�d�Z(�(��&Ym�R�ԢV�����YۋQ9K��-[iV�ŭZV�pإZ�0`��"6��h�kX�k��-����j�h����b.mͮE�Z�� ���p��rd�.��UUf0a�+�\R��S���[+jQ���[E�(*��tцj��[cZ�ڬ�j5[lej��j�p *�J
̦Q����F�[e[Q��A����E��֍�P����
�d�*�ڋЪ�-rԎ-��U\�`�hTX�6ƶ��h*�R���H�7ѣli�cV�
�ŬU3�1ĩ!������+kD�U�X�V�m�
�eZԢT��(���b�Q�B�J+*--�R��ՕAb�G��"�,���mF���#L4\�8��ZҠw��a�q��wL}��2� B��\G�*eH���s����V�Y�����C;pی����D=A.��n�v�����{A�n�I݈L�OjG��u�{^LN���Յ���!���<6���}�ٌ��
��W���`���~�ȧ�,qȵ:��4��r`��/]Bv�z�ν�w��ս YEjl���n�
�}%��ߕ}a����lv ��V�^J۵��s��G�O��O"+�ۣ�E�&3�.����KQd�Pu-�������Ǝ�߽�8�/Wi��a���C(�d8>��T;}v9,�?��_}R��Z:�񄰬��a�t�}W+$٘�X��%�����v�p�����^��k�*�)V� ���6���#^.H{{�+S�O=��z�Y�5�Y�F���+�뢇���Lpt�1�)��P����f��N��d��Ѿ�*X4�K��g����ד�9�\g�E{�,6hq�Ӣ��>6��a�+MvN/��K
��К��+Ơ��m�9*����f��S�!����5�>`f��I��1�y_^e] ._�ɔ�+v!F���rSb�f�uR>�wo�˷���w�����֪��6�_��rW�I"Yu��R��p$w�(l.~L%��ء��ܷVii���{���yQ�Wg�f�%�).�� ������uc˰����+-.V�lG����63��C�%Bd �M���f	�=�%.̱Ng6�~����r�O{�d� i��;?�n���~8`6_���R�(7
쵿B�_N�hX�c\%�׀�,��&Pe��Y��a�^�/M�[C�������D���+��Y�[z��u,y���PU��F}�d�8�V	���ne,�L�S1c�����!�>Smέ��9ܞ���������+�;'ƶl�}.��w�n�a�
��+7��8L���ҩ��J���94aPm;�;�_�ޯ����yH�	���w���ϵi$u�6Uk׻}��4����o����d^���*�gg� ��ϞKG���Ttz]��	��<�G5��>wޗ&w�F�����.�����,��\\�A�D�%�<>۩ur��jSK�-ް5�.��كyu��~��-}�8y֮����D���;�'�ҲR�3u����>v���^�~ʺ�:�;���'־Ç����;������^?�]���5���z��`>�Fh`_R�����;�v�9�.���E�Ô:|:����M7cy�\/�0��ڨ.9�H鈈˳��:c��a����x�9ݽ��x{6�8:^��A�	F����2�s��7vV_u%�Op�M7�!�3����[��&�8΍M��8��Z/������{�5���ą�y���=^u��|'���3U�a�-���~��bQ�y+�A�YbhT�^Qw����9�"���r�����O�C���ѵU<�BK�}n�T3�
z��:��#�E8��3���x���+��̻�eqӞ,=��2`���(? 4t̢�<�Jĸ3,�ag�ς��y\i#�;ݻ<�0^oj��]	R,&`L:�� ���< ��QW�J��;��2��<ӝ*ٺ1�����K��A逸��a��%x]\Rg��9=�F�r�W�������Ԧ�]H�-��Z��臄�^��q'�^{+qB.��AȠ#�ѫ̡t1��2���t��׳�ש�����t��{#_H=|`K���&Q�~*�5R���n�Ϡ������i&Y�/)!��t��{֝��X>�U�B�5�s�&���<\��;�d�	�FySP��`;��ξ��G�ׁ��W�{�Gu�h-�q��]��N_�o\�|G�ӧ�w����V�f�f'�E�_�/��j�`��y��޾tvt�b�W������\�#�|�Ozh��U7�DO�v̽�1̗�/w�-�gK����G��1/QS,,���7�bۮ����YԐ�9��Q	�6i]�8��]۪X:_q��9�:��*�]��89�&Q˃������[۫Z��ra�-�`N��������Uk����~�ۢU����51�R����f��Q-i�>�\_�x9���S��t�����$�\��Yn�<�s�pB��t�:���|�*��I����=*L�w��������VԜcѐ5!�J���_�N���z��`3n�9��.ʙGo��U�E��ŕ|�^gS<����yZ��;��v�U"���g�;��h�>��Tb�#>�Of�ħ�us��[:v��ȣ��&r�5�C^d4GR��K+�T7�W%c._%���q��	6`�&6���[Y��3�^gxq�f��K��T;a��X-�D m��} �X��3�ݑ]����>��$ȹp�Nb^L���wJ�xK+i.���N� :ָ&����Bwd�V�*�S�֯
�{�&-�R�{��i���ҵgZ����)P�^�rVgw2��J�;,�����o˴Jܣջp��̇|��ŏU\�&�/�	���HR�G�����WV=0�h�Bxmx���oH�7M�<��2������#��m^c'��f��[=��I�h�Q�{l9���͎� �kw@U���WN;ך{�#q�y|��;��c+R�mnC��gG�u;s�7���W��K1��xj̅��NS��f�c�K��3�W�G��3��{�USx[��m��o�X�=@��ଔҠ{�;k'F�'�(��|��U���+uf6�j?F�=�����TxX��	6Xe���O���e��FH��DgՑi�_���x
��`�,���l�x,��Z�u�CϽ�Y��#�3��ިw�z���r�^�5�8Ak��u<qGI���G�}�giZ��:�{�@�:�x�����l7�㔹��&��[�'%��.�sy�c�P����k�:���\s�:��m-j�-�o��>u����]S�U��3P�W�����SR����uZ�r�$T	=LW^��Ź��D����:���-�����_��K���ǭI)E,&u-�w�V�g���z�\$7ܓ�̬��|r���A�������X��T::�rV����JP_EעO����3-�wC�V��0o_�3�Ȟ���i�N��Ш������lA�Bx��CA�\œ%S��+��<w��2s���n�e�g��5�L8�mR\2΋]�>o��O\^4r�>v�a]�s�L�r�2��tD� ��j�+(I�N���L��E�c��=�	�ƅG�p���m�:��XG˷��i�7N�I�"�ݭ� ��}��]�)�����y��p���U;��y,�&���գǕ���I�I2W�^+��D�r1��Z�Z��]�7'�Epd�Y�}Xv�S3��7���&I�e����ݓM��ϲW�uo���gC�϶�f�޷��y���j���n%�`p=�3W��X�l8"��|��O*ϱ%�@z��3Pҷbiٻ�
� eӗMp�]9���R*���F�͹�뮃���E�!z
e8S�U��ijP�˅_��j��CF7�UQ�ݱ���ΫE4-����g斛�+��bﺺ��@J��o�M���Nj�(T@�����Y��@[֬u�zE�Xyj6�J�êj��G���*��}2�S�f�OT>0e+�3�W�\T%È)ﮝX^��/"���uȨS�_��u�A��K���]g�z�k;�ɋ��"�/7�A����9�r��m�P֌�u�B���,U����)��4�L�������8�U\7��ϖ:��^YǃTs��8$�pZIv=�/��R�[���m���RS�L���q��ɐ��9�E�!�	���b��Y�J��떫��H��RӾKk`P<�[8��A�x �9Μ1�[8g�xS�ff�*Dl3���`��ˈ�g�ꢠ�.���R�u4�m���X̏�k|�� X'����T*H�Ll��=�p�!0�+��&-r��Cqe�
ʅӥI�^��ܬ��W���zzJ��c���j������jO�wu����=�D��E���5�������}b�4��S��m|��//ڸ+���G��SJgަt��OWy3��ǃ��h/J��Az�ۿ!z;���n��_@EJ��+R�V2<�tVV5�t`8��(�βfz�nb�	�S�[�ދ�v�8N�mq�iq�%|hg
$Pi���o$�3>�\����MGƮO�����^�k��_�7�~:w��`����pG�P�_OR�_��.yW�C1[�>�y\t����L�{=����Ku�}�)�E��Ժ��qN*�\auZ��E��R=T\�;_U�p� �O֧���[U��QbO��2������ӣ��ع���ұ�3:x�d�~ٛ8� @��T��-I4J�!��3c8�m�Ci� ��Q{˂w�h��;��{ϯ�;F�����v�J�bt��bgg���L�E��ܜ�M�+1߯r�oN5풨7�FǨN��V�����V�^����[Yf��!�[bW����L�=wV���|��w��꾮��l��lP�j��)ӷ���	ZV��-J�H�ۡ�pv[;K����{��T�ݥ;��nt'�ט)T����]emG0�Ba8���j+rkz=�ƱP;e�;R���gJ:^����Tg{��o���2���ff���B�N�ur[Ϫ�ϫ��O+��ޝJ�zv6�:�6t�7��K��%lX��goe����,�8k���6<��)Y���]f�YrǪ�I�{7=�ex�z�c+Ze��`Aܩ�Bz냞�G�/���YT�Iz5�ډƕ�z�1L�|��K�^���É�qW��w�z�pw�3���[��apVg�h�g_O<sT��)�?e, |6x[9���$�}�Q+�P�Ƹ��ŜζH�Gg�ɭ�N{��ڭj��
�7KC���A���o����+*��~����Ye9j��{��ʲ�tϺS3W�^z\0�C�_ڹ�V%�%[U����)��X�9�o��{�v���J�z�e(��w�;�/�jx�qB|���R�/��C9AAV<Z����\�=E����gx���e�/b���>r��ofCMj�C��^�Vx;��&�Qu��G��&�]�\v v��5�� ��,S��U��E�*��N�W ��z���Ob*ʿ�7m@H�u?Z3��W%2�L�.TdkAs����Ѭ�dm��t��M#J��6S�[��ʖ�9�kaꕞ�XC}��^w�O�ޘ��}VWn�����չntqEn�'�*�"g��\)9V.���`�ӭ`�v�O�}Nozv�K�Y4��� 6������]��W�UP(�o�\Y$��S�s
ׇh�/�ZX�J*����U���U�:�)��#��f��+W��*� <r�}U6��ے+�a�\<)W+hxC�����f�ȼ5rxSixm���Y��v�͙�-Zl�z��$&Y*�R���� B���.��1=A-����շ|�8�K�ݡ����G??w���V-��3�����Ί�c�Ұb�m`�!9�о?c=��2�rf����:�s����_����4�2މX���c��q�άU��=+b�u���ӆ#���p�mWh늹fZ�(�z�������T0�,��Wݴ��Ξ(sힹ�2;fzmXݿg����{���V��V��,�Cּ"�G=ˠx�΢W��-̯�i�}5�UꆡW��q��=�σ�L�_������W�<���(q��:��J��;���	��]>�f�E=���{�8j�6�MKIVt5E�_����g���G���/����η=��YњP�bzӞ~M[�0���I�
��<�܆:)VkKږ12t�Gn��x��'�oi���>dޣ���>c�Ẋ$z.{���z��zV��rۚ�nq�#�43z��>�y��U���%ow�]��xv������x�%h�K>�p�^����X6I�*�u/�]��݃F�p[�����M�`�,k����w>�3/}��eC�K���� ��n	���-~+d~��� ���g�m�ֱa��vk;<�B��E{���5�^�����F���q��w��#t���6��׾]/	��kw����2x<�3ִK���W�➃�s|aR0}G��A��®P�%�⅌�}^����Ng�]�g��<4�,Qⱍy�P��HM���3��ƣ��-]$)��C�vm3���|���v���p�T!�I��˳1{=rzA������ܔ���c��i_��(�a�	GiA]�[�\|1Cw�9�ǻ��!e�~�k�S ��t)����fp75(���"`<�Xf����)ɛ��O�������<=�X�p!+��"����uE*�0Nܛ�U^��oƫ=J��p�8��P�V�%a��=xX;�T0`u�[�j�a�����}6Y>��v�:K	�L�/`=W+d�m�1V���T%b�����`N����^[]�&�97�ߔ�*�e^�m�t#����;l���B!�=���vi�[0*����/L�~ؑ���|�����8�V*���b��i�(��[��[�zE���L=o�]�x���Y����+c 8��
W�]0ي��Y�;�p6�,��k���@���ܝ�V��n��H�1�ǃ�hx�vsm���6�9���R7�sA����sTX݊�/1+3�=����AJvڂ�:/�N�C��$�Nӻx��<Ϻ�X�?E|W+�X�egd��#�[�s�btw9,P���Y�v�J�%�=�ƸZ�˵;@�ַ��k԰�����:��M�4�d7)��&�@��풯�9W����P#^1���sٻ�����ô�L�Y��n��#���J}"��0�4�@'n���'/��J��T7�j���f��A�a'����#���5�{ ����� �4�9Ky=3�엂*�X�F�s�aΨ���#�]�&J�M-����聠5���f;�l=l�3�ȏ"��M���]�7��g��.��N��_d�k=��'J+ O�;/Q���+BpY��5������+�9�g(�v"�tÈW|ONe�Q�`"����巵ܞ�c$N��~�����|10��ksVV,`:*�7}��kI���3��:�f�ܭW �yA�]q�4�Y�tۅ���&�L��&g&*����A�A%��!��"����cl���0*����i�b������F��5�C�:Ĭ����˂�K��U�.���K1�c4@���PvͣG(K$bb#�Ķ���׊`�ёY,_�!�#���V!�jr�&�ĸ��F�)��U�A�u�c��T2�>���a�m�e��x!/	~HP�MR�n�R2N2C�3
t�G�fY=�S����w�5�Tn�R���5�ʀ�sQ�~�}t���m��*-bQ�\j�+E�(�%��p�Đ��b���k�)��8��<��x�Z)�m3+n���������$�H�NQd����Yم\�x@�Q�Z���h!xՊ;��j��sv�Wǃ6�
C���$�5v{R8-[�T���Z�V\�R��Zně�����|��l�en	_�4z��I�ٸApW�l�D�x7C[�Mh�o-��݂7r|�J+�Ѿt��d>P[h�M[�A=G�\��k>D�6����E�&9�5�N#�O����E�:��jW$��Ą���__Rړ��:ְ3^fhO24T��"]#m�@��Zze��|�;8n��)�©�b���͏!�e��h#8��tu��-�헡d�5��Kɜ��v��-Bx[q�ˠc|;;8�s���Z�h"�K�a�R�lbKR*��(*
��JЭR���b��,�iF���Ŋ�D\6(�������a�5D���*��(6��,�EG�(��\a��ee*-F5�jU4]Z���SZ���p��6�M8Q0�G6p։QEi�
*�%�&��1h��T�#iDeaqj�Ę���
���V!XQ��+��**Q�����Z�B�%`���m&1f+Ij���,�*Tb1U��J�Ԫ�Q��iQ%�q���)mQ�D��iA�ұQ�lb��ZV6��V�l�m.�DDıJ��TQ-l��cYV���jR�V�Z-���DUDeX� �L�p�ڮ)TQ�(�Y�cL1��cJ�D`�ڪ��B����V�%EE"�VL%UV)+Q��AQe�-��+m�E"R��X��D�m.�g�{�,�3��k]��:�#��1�x�����Ge/b��W��RmI�bȄ�2olC}T��ɮ�s^�jm��9�+�Y�t����Z�lo��4Y�s�/��Dc���fg��WY�o���ޙ+=f�%��s�1�ZUk���w�ڮI|W�<%�o ��
ѕ֍
_K]�A��	u���cy�$��X=��r��+u�a�g���Ϟf��A^.1/�Pّ�d�_�kg��?%��1ދ´E��}Σ��څ����v� �gF>L����΅촓�����]^��ͦ����x�:$�ƉE�T�uN(~��-n�{w]�G9�N�v`��^���.gJ��s���_�e�]�:��3R�[���Oe�c�?w"����J4=^��]�QW/��&��ɍd۸gՕ�C��9g�}����ۯeD�Km��lA�|����F���@�2�X��²W�~~t��(Ӛu��]�����߷F��P.�:p	u�q�4[�U��"7��]:�eY�z�FP��J��^��+n��7�i��Ug�+��ۧ�p�b���`�)y���w��]A6՘�i��2�9���\�3W�t�ѵ�]m��}ؽ*M�i���֊���5T�zn��>m�4��k��Ѻu����C��XU�f���l��b\:��eGκ��q��mew��5ىч\�%��&1�Q���5V}�o�9PuBU�℗�5�։^����Zh�a�+)�e�����X*X|P��L�*�T�b�]�c��U�hoC�+r�Y���p����ꔓ�6x@鰬[����Cn��
U�@�/G:4�ʷd�c&�2�A��ah=^E-�W�~5����g�О�U���>�D�<��Oٶ���=k�5Y�L�V4�ZU��a�����s�^����V�^����[vB��Aom�l�M���<r��F�}\��t��Eb�5�F��z����{��G�X'�XHN9�:��@�y��xI�V%�@ϵa�8��j�VVŏ޶vܱ���aN�9^o4�ƺ���zP|T[2	�=x��F:��΀3�	�Ýk��|k���^�����ϼ������NN�n�\�y��b���ӳ<-���@��JǺ��:����o��f�r��f�g5�{S��b�i��{F��?:X�t�`��l�l�I3�(�d�t�(]��|Y��
�f���>{��HR�3�\��,0���Z�S���A�_�w0=�V�$ϢȸJ�{Xw���|R�X%d%��$�9�L�R��=vy�X�^����|�Ncr_�Ǵe,��#f�[�۴m�d���ǻ^]g{;�~�G�īaT�u35��?c��"ͺ�G�]y|"���$I���W!���o��5wN�:��;���Dm�b�a�E���c�tR��zp���}7�|_����\,�`4;-�Ig|�U�����L@4�gb�U����C��煊~ܸ+;��O��⇩��`�:0����9�M�tŉ܏7oҚ0�.���ȃ5����Oj��5hu�3�K>���#�6��s�6oL}����|~x �
���F�gֻ�)���w�`�P�
��h�+��L9s��NoN�h���o�C��זܭ8{:���j0�_�L�(� �uJֶs����y��k��\˂�M�u	�w��nK���F��aݢ���(�L��|�H�Y����4��kl�4����t.~/~���^��®F��ʗ^�y�^��ui�7yy�LV �*�"�y�.��	DMB���Ϊ�^ɗry������J��^7,���o����*�g���p�]l^̯hD*�:�A�|��wh(��V�{034�~f�k��s�V`���o����52W���2���)�,w��R���sl�.�~�M>ZOs�l��e��)Y��F�=N���!�6�ˀ����V*�۔o,���W��TNr�Z�Y�u)�҉S5h~{^r���2R�P9�oqT�=K����u=�8���2{*��_(����cl�8>c��/��z�.�շ���Om�;���u��XB�:��#��f_|�w���t_G�����yiYx"�̳��b�绔��=�R��2�h�F�fJ�C1��O;�u�k�s�N�||9^���2^Ѓ<7M���My�N�g��oI	���,=�v3u�7�9\ո����Mt���TY���!�F�̬�x1���$R��=Tj�+%���BX�C�E܃Ͼ=^=k$���0Tél�o3uߝ�=�ݙ��wk�&e��_�4����6�	M�8~�Y���a~��:�&��7�p�J�9>5���_4���M�l�(o�W&W.|&fI���x�SWhA����	Kܮ%(�OvKL�J�4���g�}I�X+�
T��0k����]z3w�<m�
�;\o��x\��y����]7���� B��:3���B�x貇���uQ�l���#o}n����"^���"��;�g��������mCB��p��G�׍A����r\|1^�~GW�[X����Md�ib�S�����ڽ�خ8��G���%�!#�GXhJ[~�&Ѭ`Ǖ� ���6�^)!����G��)��>�Nfދza�l��_
v��vbb��m��ت�^����f��&v��dڇNx��L�k�Wȗ(֡���CJ��	(�b��p�!�ڽ�K~F+<���U����s�Cׇ}|_.UP�Ȑ��
p��EI[����(T�9f�V��=s�y��h�Q?8}��g���J˷^,uO���)�����֫���b�>`�&y��R����n��#��qUn��Y�:�Y���VX9��`�i��Z�a/&iK'�'W�i���1����u��7�d������S�@���\��1~=C����S@LYOW����a� ���,1�~#7i꼒�^��i�����i��5���#]y~�N-��^�ۭ���$Փ�	���`uܽ�����~��u&;j+�c����T=�sIE]�o�x�ZI��B��,k��y2�9�t�C�4[�z��l�O-���W��~g�~���xA�^�7G���	�jƃ觏q����j竆UD�%�nj�5��\�<�� }�~�2��o�Uܼ˗�>���t
�iO5
��)�q�:��z Ȣ�Mmm��~�[ܫ��HI��G�:��c2a�Ȋ���x��5��>��j��f�vWS���K�։�-�2��O�yNsE��7�Y��E�$���;֪m����YR�ƀi��w�u�9�Oi���oZ׺m^���C&��O���������^#S;\���%/k��D����O��i�'o}#�[�N8B�Q�PhY�d�T�4��iJ��p4�y����L��t��e+���ݳSټ�SoJk��gԱVY�xX��~������BA���/�g��#�%{>͝W�䀡ܟi�gv�{�;/]�N��^U`�_P�� ӊ��w
7P]����&��x&|x�~	�b����j�Z�͍�^3>�y(z/r�(p"t̢��)L���:��o�r��en��e�<|:�~_��!��2�%rҨz�=� ��,��b2��yu����cD����}�̯J���tR��K���pw��z�[��=~�9�8�ͮ���y�s�d���*�:�Xog���2��젔ƸJ��w�=W���K�:f�ӳ�(t�
�C�k�a�����t��ѭY��c��i��.�2�����/]u`E�f��}���*ecV�u��˥���}�2�V���!z��vS����	�k�c�x������+uF�̋4Lݭj��� J�b웗Fb��"̬��܊���i�M\芐VH=���Kqzoc<N��*���K�
ik��7�W]�|$To�$Rjf������0m�"[R�Ѡ`+�OӘ��7��u�O��J�Hpz���?nP9�	41il���uy��N�X�^���=���5{��-B�[�Ah6f�k����碯��_�pV�?�qv���}��3m���jC�ݭ���������vg���0�԰�;��_���)$�}��8m�.']��Ty����T�U7�L�o�9u�+�;0�,Gs��gk�x����E�l��]^`+�|\{'V��>���Ou����05�[��a�h�|Hd����j�v��\^hVx�\�w:l~0�z����MQg:�vS�_Ku���qMYr+;>L��LE��jl���/qE#��:�T�%�_��O_�B��foV�C���:��ik�3�^�|�qm-�9Huq������V8;&�*���v-E��V��q.A]G�t���W���2W�~*}Y��M��&lfu��r_��ZY��L��l�V���
.���9�e9��P�0b�ěwR�b�8��G�����7%�V��F{Mov���L79�"V ��ӭfc��
��Sݲ�׺qM^U�}4٭u�3�M�I�\]x�5c���;���>�~�XMIW��E��r��뭉��|1�Yk�j
��,�uj�lV�R�G��)�8j���R�-f{�Ϲ0�r�ly��C���2�`�s'���W�ߊ�k��Z�EՐ�h�FNb�o*z���jcޮE�2���r��.ۍffo�aN"�]�>���ʆ��0���ÂS�g���g�N��1��y�2���W��@�
C��]5B��D!��\�� �C��;YlL��[���~u�|<\���S[�����e���ں�J�W}��Һ�p��ˆYkD*s�$X{��gO ��J{�#��f�!c�g����uY�;��	8�C�C�ư9^1nk�o����hE��yx^��D�g"�!u������T.��CϪ�^�C���ig]�!WXb+�M3Y�(�C���a����rm;~�T��W\,�5`y�17�7Z�N��r�O��Ŋ��r��3}�z ��gÕ�����8È���MC$�E�����ȷ]��q��|Y���!�VwƱ岹`���J℠F���v	�W���2�A�k�t���ȷ҄�=�a�{�w�>�>��KQg�@a�����ۗ���q���t�ckՍ��*ͳ�*�cGJka���]�z���{�eC�T9"<_��P��ӣ��a�]F����]�`KUt�a���E���YC���CfP��]������/����<C/sm;��E�;���[����,����B�fQ�J�T�p˔�����bG�uf��6|3E�ld���^R�ln�d;[XCʻ�p55v ��zᖔ�y�[��1�Y���ԉv
���
��v
T�.�k��윭^z.�?	v�f���x��y�%;2���5��TtXbT���]yRӐ�i�X�x��2z��
��|����7�~ܞ�y�5Y���j�/�u�[Pл�	V�I�E��6���gԶ�΂w��������ef�|���1h��.�̛�ԫ��*m����b]�qp�!��g��~�u���p��px�.���\|1�w߳*���,�H_o��V�)�QR[󂑿A��C�	ԕ�[]���=Ä���\Y2��z@�H
����P>��Nی��j��a[��9��/̵��Wv!Pk���zY�;���b�=�X>�T0X�f(=�kө��9�c+׊��e�>8��+����=!W�����7�O����r*�gC�2�6e��Ok��x��4<z�ޞ��òV�a�����gь���䞟�L[��^�Xn��������z��n[�<�Z��#����{JuL\Z���9E*�=���j�ׅE_Y�*80)���<�;�|t���N;(.\�K���1o.���<����[I.��j�;�x�����B���.�pz�r��w&D7pG6�&�+��١]^�VC�5��4;e��V5����;�+���S6����3/�����;�����n�nn0�L�.$���ʽ^3]h#�y.3�N(Gy���̍�sL˷�˼�ox��S��Zb��\߆��7W�՘�3�W�Y��j�K��Ը�ꁙU<�3�_nIB�D�5���I�]T���\�9��r�Jy3�h�[�q�;{�^���йq����e�յ����8�uW1A��h�w�V�����ِ謬j�Y��Gs���d�f�X������m��b���BoĈ�h1�)Z �t҃q���E��-���-��̹޴��3/����;) Z�M�e���0h.(H0��+�X�vܘ{+k�b�×���\��Ю!ꥋe�J��c��U��s0�{>ʓn��ڊ�P���k��ͼ��unK����%��s-�B�t����^/3����U�R�X(@k�ҙ�R��Ǆ�~�m���ᙃ�kw�hz�����T��.���6|8]��g"
���L��`x5q�*���z�O�y�Ux��Ef�v��� �tث���*\�w(�yU�`��B���+3��\��0m�cT����d|�F��Uɜ��Ym�`,͉�������*{=��(l��7���i�Onq2���O�Z��P6�3�Ł�mɜ8��2+�+X��D���A(���g�ugwm��d�s�D>�l�'9F�i,WxR]�
t�s@E�j�F�1tr�mZr�:;�3���n*��^Օ��4�����W�J��uK��s��v@��gD͕'>O���J.U�,\��Ů���L��*�5�5Cޱ6"�ׅyq.x�ٶW�`㗋:�,�XP�^W��r��[Ѓiޡ؟me*�x;(`�A��SH�����OM���9r�{���ك�e^��Z��=���Y��S���;��8�4�w*��7�t��� ����r3���6��%+��M���Ԛ�U֍�3��3�æ��3:V,�Ș�1x�6B���9�>���&Wj�If	��J{M	���d���j���(�.Ԋ�u�_)B]��Μյ4�FѲ^8	���._�Y���yu���d2�xݙ�4�Mվ��t�����=��a��n�W+=WBy@�BG�z@�K���aV�w�r�]���D��+���Tϭ�*S>�ɲ���{9y�sq�"������֙u˶d��A��"����ɿn�Yy0�3��<}}m�X��ƭ� -�J�B�l6wK��Ar����n!��JdqM�)�K1%m�m�wI����b����Al�5eR��1awl�O1*%�M`W}<��ʜ��|eb��4�[�ORB�#���f6M�$U����B:�)��Ɣl���ıA</��-L��t�>p�c	pUfAq��*�5����ϟ��Z'�!���p�!C��`�3�0��c�3uu��&�򕙅`u�̔Jb���:"��SH$.`�+�ш7df�ì6����Tе�=�*b��O�:�B��z��"m]JWt!�m
���RsQ[��h|����4D�(A�S�>���JX���"gāC��{}�2|
��R�y�Q��m���s�i�kAƎ�8�p�q�GiZ��9d�\)c�b(���0m����l���/�����}`�ɺ���}�Vyb{��w6����"'�74�(���+*2S�SF�׎B�����5���)]m��r���8�lz�儮�枘s��|j��ӥ�TD��Ϥu��35�aCQM��I^>�c��.J�!_8u��e���J�?#6_M�xS��b�R�fQ�@�F�Ǳ\T�Z�I僳���������C��T-EB�J�jԠ�(*ֱb���p"�2%V ��"��J�#mAQ�V���EEA���$�jĊ+�a����b�����U�(��ER�U-� "V���D�����
��82�*�e�EIJ(��.�j�͒��iQ[mh*�,U��1QVڠ��b!iQUsJ�(�%��Cֈ#"�U�DQ������`��3
��QX0c���\4D��PUFAm�[DPDKB�R�ŵ˅E���[h�1��Z�Ȃ"���X"��-KR�Z��1QUqjV���Up�X�U��,b.-�"�	R�F**�[h�����1DUQTb�-(�qJ*�U1��ʱPUTUX�SITE"���PX+$b��l�"2�ciPTFi�.)Uy���a���o���b#���e8�71f������E7����lұ7�gh��=�m����L�N�����l��|�z��mvg@�0&@���2����· �x�{�ߌ�T=H3�^V�g@3���J,�i����������kqݟP�f��i7�*�O�>��!��N�v}A)�eW��6�]�+s�I7V�����W���`Ʒ�Y��-QqD�"�Ι��aw�GV�	^[�M���:�m,�+D��j��qt��Yަr�X��g
F�UU@��ًz����Kx�����\j�a�*ϋe`kL����3q\ޱ:���S�4c���,����5Y߫����ų�i�_��r]��w�p�pt�θ���Nܑ�3��V6h�����jW��\�^}ִ��?,_���l�H���]�xXv���^Jq��dOM|�'[9�[��a�u��п�S���Ӯ��ª��<%��E�}���57��=�l��Y��r{,��_�}��q�<8J��m�[p�w�%V�xo��{��&��Wﰔj/�!�??g����;�̳5��P�>�A�B�.��1�34�H���LwP������a��a���y����Ưd��41bv�B�%��i\�eV�CB�����+.�v�W2B7I�晰8�r��Ƹ
�V��X��׋_j�ͫ�u´����;6�d�[��С��]Do��QGR�}c.%��[�8u�UŇp�3tC!���[�~8vI¯�~2���:������9���u<�Ъ�]@>�~���:徯K4�P����PO�+<;�9>��z�]s�s~�֠�,4��u�ukZ�>c��2��L�M�������%U��V:|k�p[�:�����{j+�Ww=aS��ސSDh2��V�5�����y`ܗ��g�.���}�P�wʝ�|�u���k�95���~g̪:���OR�ipT8~�s�$Mz�fK��v��A��Ⱥ�:Vעj���@�:�����e��Ƃu���4�T0�u�F\.��n�3������햎����d/=vD���w��i�c^�"�xy�p�ν(�j�\6�\�g����]���p���ɞ�G\`��o�����Αu_EB�9m+=���N4���þ��k���<�ݝI[F�����,k�Y[���p纬��kL$��i���M��YP����Keg����/�9�Nݝm{ᝪ�O���W�p���C=:,�^�փC=P�sΡ�>��o��o^��8���,�;	��y�K4����x;x#�̳�;��X"�GX{�@��:������@.��G5�����g\}��F"n+��J!�O��;q�6g�/��Î=�[�,,�|��N
B���(u�����+8�c�E�G4��"2"��'^���e���s~�l�vy�����z��W`w6�U�t����n6��l~6����S6��Y|�� w75�,�r�$��^͸S^t`���Y�W������;�=��Y�6+�4:�\�eY����<��	�!ɕ܃�W�R�%��竅��[8d�=��y:�K�m�;o��	3���֙�Vx�C�O���=L��vC�tʇi���e{���B��ݯ�,��ҙ�P�0|�[>KGT�9�{2��iu�<)���3��ս�5�`����yu�l�/r�(&P�\�����Bĸ��m�d�7��P�C<�ZK-�Ym�Ao.�^�9���c����T|�\�
�S��5-V�φN��<+E�9G�2��^�5�\�pe�=�0�:�b����(�[PЧP��0�H��/���et���q��ly�{����k,ں|�d���]�]AHn��m����d�5N����K�^��u=K+�3�;�x��e���*� ��t�B�^'��M�5��X��\N�oL�Mx �Ok�伂��[��"Wz��sZ����Cc���Y�傡���Cmi<�6���[W��/�m��0ϊ���l���Ù�������L����z����g"�i�K{f�nʗ�=����ȩ��f����VB5�-��{��jQ#�<O���sL���_��a�y���{tXBU��SHQ�[�������{@��UI|���v�Zvɖ+�8���N}]�-C��^�vjs
��%a��=xX>�B�`B�y�{�Z�|����A�� ���͌J��,U�>\�r����)á'��v=c�FkR�`����N��s�%i罓��⳧a(��\7�K�r�=�Ci=�[m�G������i�dЮ�؟�y���l�c�/���`�w��>y�W�H+ƲpB�M�z$=���;KceQ̩�8��3R� ���}gG���r��=n{��Q��bډ!��kҚ:Ŋ�_t��9=�p�&��,A+"�=�Mh�X�5�P�ya��y:���Z`�SuX"���lI��}��W���n>'Ã��Y����ف+�8�h�W�ض&a�P��*�*�1a����]eh�S�=���ơ���h ��oA�%���j�'�w�/����/BE�_=���D�3�V%�-6�������emCs��Z�I`���2�0	O�r�����udfU�d�	�r+�ݶV�u86uy�V�o��V3�}�mrtFz�<�N�S����׸�'!+�1{���1��(<QL�f��ڗ�5V�Λ�Ֆli&VR�Q�o135�Nx�s�u4�j���z���=nͿ��������oB�(H0��)��Z�ל�tι	����;j��|pn��k��R�OR���ݻ�
�V�r���3�3-U6�sN�h�q�����=S�>v�����]����瞢�C�(@kGOve��`�)��=�]vQ�*�f�	BXW�pTx�+�z��i�χ	U������:�C�s��<�j��S$���*�J��;��+�Z�7��+��krW�\R$�y���2m��Z���^�qM6=L�5��-)����J��9�g�q��9<^7�����*F�,�;]�Ҟ������ 7KA��Zc C��j��Q+,,�ϧR+�5�F��z�ʖg���eǝ2�HzST��3�{)y`ế���0X�V�gU^q��9y,3��=�9P5�U0�v�+�2n��W�	U��Pt��J;���{��x�R�o�{.��I�������t#=�M����q}�Ζ�؉���Fk��{=LĬ}�����X��� �7E�)ڱ��C��ӝ�������0?TgNYW.X[�	���vgn���f��^tN�Њy����y��ٛG7Pp	���` ����<ze�f�m��nY��q�m�f"Һ 2������]b`����ۀ�(���@����t)�EvV%V-���r�#oN�y�9G�ɽRd���z��~���u��S��:�w=��m�>�-���}��o�(\�Iq��M �齁jӹ�i��t/޺�����+ś��8��0��>��ݍ �3�{�����b.�y����ath��q��k�ja�_/	�����|1��c��_"���#�U�<u��Ǫ�C*Y'��krab����3�P������*��.>���qRM�w�}���Ѹ
��@���fe��r�/>��^�*��տ47:\>Zj}C/Zc:�nt��f�/��f�B�{�2�-L�D��p����>�\��fz׵��g�6yf��P����/ k�Y���Ұػ�W$8e��_�V��ZY����ov��|'�M{"ge��\>�����q�,��i0�=�^�G��]Z-U3������G��^���|76�yB��)P�m`�i#	���%�yr�gźѪB����ML�����K2�x:��1P�(bT<�CJ�a(�j�V�A��ΰx��J����λ��	D2O��au�3RJ&˥��!�g��z�kG�4ϼdq ���z��.���wls���X�.�GHSh`��m�I��Mů�[��!^2� d<��|x��؎\���¦�5H+�����ΰ/$���xÔ��������x�tfq�7��0U�N	f�VOmÀ{����<�9�^�hj�Y/�}��}y�>�X6ڱ����U��A���g�V-=̠s�P�o}L���1���V����F��+����t]{��>���_�B���X]!���:�{�@�^ߜG��Q|=�M��-ai�(8�������6��y^���W`�	���uL��L��F���.�7F���ը��o�%�m۾,�l�p9C��+���\�^��G�m�[��L;8�U��^KF?�o�&�[zrvxt�A���r��9x���6�QGP3Z��6�2�@b����9�m3�`�}�!9���E���|S5 �Ȝ?Yv����^Y�}n}���[B��K���o�ե�֨+�%��^���Z���+�N{�wz#Y@��c�>�.��dW�H��:ϊ��K�K���O�J�	�=�
�*�]7��÷CcI�J�tt�iĴ`��pi�m�$�4VV��Ƽ��h5�V^�L\���r7��u%�����=����V�p��&�����tl��;�e�ݞ���5U�=��&	3glR��;q�S� ���˔�`�.O=^�I���*��X�O ��c�҇U�נ�n��!�Ҧ���~��W��m��'y�y��L�|0�R�Z���a�:�e��b��L��������k�N7Y7#ةfu��ιx�k��WU�+����k�V�ˁ�j��bO����7{;��A��[��)A\+�o�Q���X��u�Gp�l�G씩�;h��N�i����<�2���K1#ԡ��
�)���՟E��R>��x�1�5� O����Yޝ�O1U|eWaBH��� ׊�5`���^��}���V.W�뉎�����\�Sg�9��M�/v�z�����3y}��o+�� �Ӄ�D����#^�k�k�N{7��V�A�݊���^��o�@��h3T1uY���iσ��X{�V��A��X����R�ujcx��U��3r�3� ;jB��i��!��Zl7Y	�z��iGjoA��غ�}M�<����[�8��=xo��	<-��V��ƻiX��5֑��ɂ���=U�{���=�OZ�%�!�`R���W�W^�;_Q1��w�A�H�,Ƕ����Q�&ᙼ9����Ub]���\��<1�ZɅ׬��:�i��]�yd��ynX��{+�s-�y��5s��f�$����h�vtA�r΁�s�V]$+�#ڏg�h�
6S><��l�ۉ=�|ɸ��f�;߉.O9���0å>�/w�iJ(i�z��u�Y�J���yR����xK��1����'���C`��2�{
�`�T���Ɗ�0M�Jz�=,8�`��w�+�~W��u�:�;Y�0��x� ����ե�Up��[׷�6^k��vA��_W�3�V����;�;�}�V�8_2��\��]���MX9C����g>*��!��A��u�Zk|�%���9�k��цu�q�[�d��뽛�[�[��n*`�w������yW:8��c�G��G��h�]���>~Lhs����33˽���c�Y\%��6�XW8^����#�,�9{��
�˳��3�כ��f�Ltr��NB�Ke^�he�(/2t&��������Þ]'���k������=�i�y�]����=��ϸ��Cq�¬��x�{L��ᗯ�4B׈�77pL������/�>��!Q4��h�z\�9�>[y7r�����C��*�����=����
���v
���M�i�+��m�1W�!��Kj]��d�`B�����rᮨJ�����Ϋ%4�¼'��V�_"��/��y_h�s�4�j�X�W�bO=�.��,��ܬ��[��<�9�|�m��j<�=��bib���fC�R�s�vR�&o�/}C���6k���;�����c�/;�Us��u�{��\b����c��ݠ}�n�寰��;��7g�S[���5�V	���d���~�1诮Y>���������=���`�ɀk�|�Lۮٱ{���<�W�M��ܣu���ܱ�'I�u^c\K��*�����es��ϥ��_I/�J4^��Xe��q��J�̞�Y��#vp�����{"~���sx���u}w*E'MLVo��0Y}�~c�#׺=�W�E�Z���z�Cn�� ��y쓀if������`�(�{�̟�.�:�W�����R�Mm�ޙ�ocz&�¥���a+w!�i���1�{��c|T��C��2���V�Vvxɋ�p}0,��[�rE�<�a�	Ϗ=�4���攝p��
��([�T�K��ǅr2�2�D��yIs#�R�w�M�n[;�Ql��:j���h��gZ��xo"�J$�e��8NeI�Ճ.��y�^Vkiق�	f﹊�5�D������ݫ�
�h��TD���A����t�7<��0l> �6�<���Ƭ�u�5ث;s����M�#sa"�6ګ��ӻ$�y뷻���ռY�}� Q�51M��q���^N�츨6';�y�����n[�����3._�qUq:2��G��h�]��|�b�YF��)ˀO7����=q�/_w�paU����P��/m�"�'G5��q7_�#�G��	�=r�(M�1@<������Gv>�p; �;�vγs��G\@�S7tv�j���V-�����������8�P<5$\�N�:���O���z�i6 ���+��C[��*�{No��Y9�)6�nݺ!7tҲ=���>�E9���,D�S���7n��"� ��lޜ56j��{W[�)d��$c�=���0�0�ͭu������ ��5�X�Z�{O�^�z�S�[8ƌ����V 䜒�L��w�<�j+�5��w+mգN]����3>4�^�)��&+��l�L���+�L�����F���k�������������^�Q��5w��{㊸*�ݑn��%y�����D�I��-����/qn^ͦ]:��`���-�4EDv��1z��gq�]0o��=�>Yح��{(�*-P>�ѽ9��U�=�0�(9�,�1����Mw�|G&���T��v�\��SߝN�׷C�c�j)Ӄ�|ADd��Cto�[�b�P;�W�c:�J��0�qF���Z˫
��pX�I2�&�����<|̚��.�	��|h�pQ�߽�_�v��h?��i,���I�SB�J�8�cʁoN�p�ԕ
$���p��a�[r`�n��;����&#7G��8��9�6 �>�[J9�j�˃�-V��3��O��겥�/��h�
hpC �	u������D&��a�*=�hN�om���k�su�z��ܽqS��a'� tM��W�G^8��M�n���x���fM����	���M��F-��]r�@X塥�ٸ��n���k86��Y:�����#�!]�X��ִ��5�8v8�����cG͡��~�/5T��a�E�51�*]E�dHt��{,rڻ��^T�y��c/���&��J+87ov]G������y$�7z��w��W`��7�
��{���,Yq�υ���[h��=��|I�������UX��,F,DE��J��b�'�VDqJ�(��1b"���������0�EUU�[+"�EF(�U���#UUTF
""���"#���-�(�c[T������b*��X�DTKJ+�FGQb���AX1UUX�Qb � �J5��"��U�)�T1h��1J�*���P���+b�PX�¢���UX�V(��(�*�F,TV2"�������U����`�`�E�dUF#U#DTQ�"*�T`�*��PF*�l�*"��*�Z�*��QV(��KDV
��Q��UU+Z�ᨱAE�dX������Vi
1�b"�2�H��+"�DQb����QՖ*��Z�DEQTd`���"��+Q��S�X)�E�� |) d/t�V�\���9���|y��n�-L�j�ᵎ��A(ya���+��[o�,���.�ȭ�R=c+KX�d���<��r�����_���;�52��}O.��u�܆�i����Yg�p���K�ӆ��R��kF8���:�U�=�z��fTa�m&-�y�훇^�[�Ϡ� ��F�@��"�k���=x���Z��ϵ�/,�*�L�a�/<$9�Z�E�J�Q�H�L�nl^�]fҨvN99�d�w�둹;��ei��W���S9۝�fF��K�cos�%ɴ�7��+:��Sr`��B�%������륹���������	3��j��������X������-��{�.��.�k�J��rP�Mܱ�_�=9��v�z�wu׵��]�C��\k	�d}�)�A��%ޯKʏ��-����9��}+�ζ�O=�U�WW��s��1���a�ױ��n���M�H7���c{9�� �RZ�������sT�db=�6�9�����C�y�5[n��^A��K{���lpy�r���Ԩ��8T�Xv��*R�,r�ޣ�F@��L�y���/�fS'S�.�F��uwI�k8I�˕���.�]qz�i��t�k�-�њ;�����\�"e-����/g8S�\wFs�^�;��:OC��m�rOtV����L?r\�晔�{��e:V���f������s[���.�<�^6���y�bw�V�}}:g��z���H���liܺ�X'�}-nH�oby��sk���+F����׻نn���
r����,�v��4eu���5�:3����V�Z�����:ew[��u1u�h6�x���W��/�Ey%3�Z4�#����e�~
f�9]�ŷN�1]����7���������S��ǄM��|�U�ek�F�d�$�[{tJwv�׽�d⮱)tj+{�J�X�z�[�̏,n���k�CB󗖐^��' ��]i��.�0zb���xev�M�
���L�1m3�s�܁jS��}-Zxiw�T��	�e\�zb��Lvn|������5�9
h� �U˫>��y�n������v��E纴=<D��-/����ٮ�㮮˳\��Uyh���LU'ud`n��H_N��\����L�ڛ����\
�;D�͚:���<��9K����G6�Žo��<�[Sjm)<�9%l�W�5\��V޻]9+���`�[c�C����j����c9����^�ݯt�^��\4[�+��%�֤�{��<:�����2�;b,�C~��`mz�.��y�5+mþl�!ݯpuJ==ZBќGt�]���2���i��4:��W�%`�s���|W�N����7������g;�@�� ͝��1��c(H+]�ۣ�fC�����~�������L��񸑞���߻>���I���?���+�΀��|qkOӽ�Sy��S}�}����x����>���*�����:%5��әi����tT���s�;��s��$ޮf�����9_(���U拗�/�������>v��_��B��R���gS+����x�n_�M;W�t�܍�9�H.�&�m/'�
���I���P��w9��0�fs�v���@cT�;��q��.^�.�ɂM�d��*�s#�M����cG�zr�M�s�`N�{�R"�bl�?Osg���G��1�2���h�/�o/z�P�מ\����uq�x��-�N�ob��y��}X�V#��1�*�ǯ췶f��y����Y��댝�o��^���U�"K
8ѿ�⯓�����Z1��]):߻ޘϝ�C}}{̨7����q��H�|�T�[Ӿ�A����d�ϔ�����^���{������P�����X<5�!��T��q�߿g�3��?��~ڤr��� ��t�A�i�M��H�������-�2)��C3@*����{>��3c=��ˋ�S���Eׯ��w�s�'�/�#vr�Պ>�j��{�D
�6K�̀�R�&��-��y�6��w�]�l��zvăk���Vz�S���b�o�	I2�!����k2���rϽ��.����՞�Lu;9�4Y�W�%E�u-Zm;�ꤝ��t�]:y7���a���6�hS�Σ�Ėo�pm���,5�&���X�,�U�;�Y�r
��s�>�_W�gi�Ca�x�פb�k��(-��EQ�8
��#�&�2�e.��d�j�*���ԭo���R���+���lO��6�Rی��a4%�;]d)���:�[���÷�+d�q_��8��������`F��w�^/�ΫI�����k+�V�od��s�n�<f��3d�v�9��I�d��n��ok��W��r�u�6�/RK���݁�x��{�ݑ;�$��'K�xj�I3��VO��=�N��3��w�9����ی���J�a����o�ѻ����@/F/��4b��4.�r���0�}���Y�͝���sk�y�Ý���k&�W�u*m�`K�S	�c=3k����1Wﲝ/���J�����;�¦�|�i�Pl�zE�ф�k=n�ܶ���2�������`۞V+2�˸�a�/�o����jh��)ػ�3�=���n���Z�3"��A�@�^`�V���uB�z��r+�[��p(��3̿SJǩ̅�����I�Մ����#�%4��ƅ���p��l��RgD�h��ܯgl���#Ԝ�%9V�ޭ�JF�o�}5%Y���9o��}",2jnխ��Ž&��_m��r	
�������Ğ9kN�]/rb�h�Ԅ��}u'�����<&�^F�j�7{��6&Vay٨Ξ�d�}+˝	�3VQ�n��j��4���v\��y������N7U�U���5�9�|�x�=�+/ҁ�ɛ�cg������O>�x�D���nh�i:>)
Ϩ�^Q].O:���j�&o5���TzP���z��.���V�I�ƦW�5w^%���S}6�����k2+c�n4���.AW�W��QY�q����рJ~������َ����s����:��A���'�,���\��༻|2S�����󯷮X������<�+�7�B�G:�q���ϼ�+>�1_r���bn�ŗr���W#ޖJh���Xg���n�se����6}�Ǘ���M����³٫�$��]E(\���B�x�i���V��Ab�5 u�A�T|��V�f�n�8ifm��{p�h���6Z��`'(uAA��Nga�=���P�N�U�\;&��ʶY���|�ݢ��9�^�\���b�ut��װw����[�X���=..۰�q��O2�t*d�hp�PC��"2���:+�#����|���^�ݙGo�y�ȹd�Ρ.�A�K�ao��zK�;y�Z��]{�����q/�6�a��(=FA��s�o��G��(J5,�x�����]f=��t�V�E�^֍�\neS�UA@{|��z	[�>�����^�$❾�~e�Z��z��gOs�}���w�g�2�N�Sc6`+�]�*#a޺�;��y�g��{}Yk���C�*rGn�v��{�cݸ#�gK΁>�otw/r7�	<v��V};�}X��3]���������=�S�sn�[�Ԅ��C�K�������v�l�f�q|=�,�����!]��b}��ͭڃJ���|��@�����|�,�O��Ӛ���1��;��uR�Wd�m\�}u��H/F�_vxu�C����s��զ����ޢ5���s��v��s_87�!�A�/�"�}��.�sB�_z�����_��{ܫ��@!�����p�P3���HkErT�vX�o�(xM8�]��w.l���=C)�u��y����DȺ7�@x{���Ӻ}T���<8N^z����zn���5�J���AOO[�o��A<]Gd��]�����s�^�$7{�H�]�+�>��|��d��um1����ˋ�3�o����4�g�}���Vܱ�7��hd�z��H�g�u�������ح<-y���{3V�̸}[�.�3��Pw�6�̠�ݏ�W�c�׾�]L��{-����f��Y�ӑW�0j޼s}ù��\ ��B���S�x�|w)��.;k�W��z�4Թ���_/�Y�|k1D��tF�ڥ«�g���j���y����1w�h-���82{7*�z%C�u|d|b;�*֨8/C�#�^�Y��x2]��Ӕ��F~���ޮJ�ne��ŏހ���(�a_o��8ϬڂN/��'��׆;����co$���9ƹ���
�Th���ss'��F�ɀ]�����gv����[���Ε�]�̲��Լ^2�{�}zU�8>.ڤv��j���n���s��b)�gOLx��l!.��C�4d:���S}ig�;��5����QoP�;r�9z�Ž��k�:ah�����96N���M^��@�7A��^C,�82�pO���t:�q���{�2V�58a^R��ֳK�w�=�νW�bX�\.����:�k��mi^�ŕݽ��:�V��+�:��������qe�l^#�BugDu��:P�b?u���T��cX#��{3&��fm{:FMm���	x=
������{����o�Y��zñ�~�J�-̙G����m{��ݹ�8��/�;�`�?s��Xx�J������o��[�㺔�ި�ԫ��ˣ�O��%��'��^*��R�S&S�ǯ2�J����[�hF��>�N�]�N�������:����/�.�#YY>��u�2Hkg���BS��w|�VCV�.U���F�����vG
z��y�{�5�h�*����.V�ǹtgT�)i*��3J꼏q���//uמ�X	ο�@ۋ�⠘�q���)�׭^���Zi�ۢ�=l�7L�5L�9��zv-������u�7R�oqs��-糋}�Z��p�=�r�D ����9u�vK�%땈��Z�����ɳ*P<�۝1�3�s6!s�Qn����
o+Yb��\���[�Npȸ`'-�黇f\}�j��h�
�	���E�~��dN�c;���r�X�ƲM�i���:k.��S<"�}��Xrٮ������ȿV>����c���y K�3�����Xg��nw=��*�L��ݼ��q<�' �_-ͷgv�ܗ��cE��yr���͝:;;�e�`���GJ��/���`�����<���J�fK;���\�u��^�=���ZL��{��+J~�?\@5���~�NP�!��s7�]��_��
Cr��B�͐���a�_vͱ���=Y��>uپ�Yzs<3ov���H�V�r�mպ�G��M�z����ǟ?s��J7ò���A=ӝ��?@���j}���1	�%?=X9�s�.��Jv�U�^}%�j���^ga	�$�W��n�Ԭ��kk�g�5���u��C���IO���$�� IO���$�	!I��IO�H@��B��@�$���$ I?�	!I��B����$�@�$�B����$�$�	'��$ I?�	!I�`IO�H@�p$�	&�IO�����)��=E����8(���1%���U)%H����RU$�RDUJ�%I R���J���R����$��*I"R�)R�B*�E)P��)B�H�UTP%B��	I%H)H$ �3*i��5SlT)(B�*�6��P)B�J*�JU���*Z5R�kc3���JJ
�B�4�UJ��U))HR���E �PD�Ti�JHBm�(��B*%J@H*���ԄH��   q׍��m��hkGAәU�Q���@M�h4�Z�avt;T�)T�hYFj���u��L�hՕ�[U��l�� �)�4� �
J"�  �1TCfW��Ɖ1�QL���¶@ *�*�ABf���M��l(P��3Q4�-�u�l򃜻�
B�
.�*�BKC"��"�Z�p �
(P�
.R�(P��@(3�� P�C@�eٸP���B�
.9��(P�B���(HP	�uV�Tj�������Z�V�j�l�3R���U($J��5JP�  Z�UF�P�02

�YT�h�3#iZ�m��K�j�N暌�QT��1��Y�hi�n۴U�5ݩ:3*�lh:�D� ��FڪP��  z��%K�P�����m�@��*mB�5Z[��6TZ� �S��S�jU�uªqV��Mv��4(���$R$��Q�G�  ���MSB�SJ(UZ#i[Al̬Q�I�l���܉��	CiJV��1TPe
K4QHh�!EJ%*�RQ/  @3�= Z%�4[`�5U���h�e2� � -��A4K��L�4�i���J�HIJQJ��   �Ѧ�6�5YV�`U �LU jcC@5��
+-�mlɲ��0 �hj�T�D�T)*�)� z �W�KF*��,i@�b�M� �PT 
چQEj��h�i�� f�B[�9���BJP�i���T��   �r-�wT]��)�@�!��Hm�5�P6Ա�4�е#R�V��m����w�� �4�
�m �b��Px��T��  ��$�*   *xS4���  O��Tz� h*y�U 0  $�D��J�� OY,�f,�y(�3�1C��L	�
<�	h��k�|�y~O_~�+]�{�0$�	'=�?{���B��@$$?�H@�HB����$�� ��;L�Hg�?�q��_ŧ>�ſ9y�G"��%%n̙ƫ��;�7FMњ��&,ǒ���J7�m��{�v�)�C�����D�pɷ������ ���)�a��Z�X�'�X#w07El�3�)��	�v�����I�c� g5�U���;x�-]I���m`8�(f;zi;:�����@��4m`!YZ����ܬ�B��9�*�xJb+�4��ޥ�.Σ�W�mR��ZE��6-Z�yCiӪ]��<x���r
��^I��F�܊VB���w-��wQ�&�4KݽR��8W�����mf=p�a$ҕe�c �B%kFB9),�N7��9�EU�����fZP�(�ۧES5zc�:h�!Sm�Ij�6nә�Y�uyaMOn!�R��d��+�\hT;yY�+�s.�$X�+�vQr=6�z������cފ$�!��khSA� �4�VVV'˵Ww*ՍK�U1KŏR�Ma*�XeMz�ѻ{�
1Gbې`�[�޼�5��ԥb^
!k��ӳYL��]A*��j[��.�ֆ�wG�o�o�j]�+p��+êVH`Ulh�0��Q�3q�%�M�����ګ;��3�h28K�qd��&*ƨ�t:��A��"��cy/u�kS[+W��x����n���7�� ��\I7*K�Ɩķ$�v e�& D�E�,���2U7Xp��:�D���Q��-6�j��Ϸa�(���w�I����
�C1�0�Ä-T�
/I�����5YV[{y��"���dSu�su�})U�A`X9��Q��7��TE��4�N�˰�9�&Dw�kCx�)�,��(�]LDaQ�	�r���Sr��㰈wo�����c��~J�C5-l�����*�M�P���`w���۫�A!X7VS �
���,+�Z��1�w�	�m�A�B"�e%���tث��Y���%
��lp/6��l��]*�!D���aD2����J�Jٻ5$+K��FìhŨ�ފH�.�"��w���t�z�^�����	�U�c�3U���F�k�Ls���{t/v�y��ld�bdC+�����mMWJby.қ�(�M��8a�~wOP�-՛8bV6��a_׺Xa�7��'c�5��d�"�Ѣn+qTӭS��$]�tUD��FoU�	����j:;G0�vs���,���w��h�Щ6�ٮ�זN+:���-zn���6�^ȌeJm@��2�s,���ڴnj�[yf٘e���o�26r��[��&�����,n��J�5�35��M F��2�(t]�$������rE${��co&X�Q+ċVh�"��{z�V���E�Q��B]Zύ���R��Q܊�x��Q��8d;�Ѐ�è0껕�"�"�x��&-iz��j����5b{cuN�X����9��T�n4cg24�C�v�{�t�r'��ڎ֩C$&�����	`5���ښ��[�ב�n��2�͍�Jka�!+[h�X�9�v�Gxh�@k*lưE�2M�D��GQ[.t��`[��!�5����6�m��WJu���J�&_LOHdڕyVd@
{�%^Fj�a쬦�[�S�Kܨ��:��t�4NV��:�{,�ܳ��lR�U9��4ޅD��ϖG�,��7xu`n���w��)��2�n�h'�lPzwx�+)������yx��)+��mmK��8�@ʱ(�?]:S�%*2��aH3�яP(�CJ�eR������DY/2�f`%�3%��g>`� j�M���C�jjH2��x����jR+�aBr��ދ�N�eC���V�/B��j�ɚ"�J��n�f�q�$��+P�8��D�r�oi��%)ˬcpEi!Mj3J@�tF�LH��	TfQ31�C0ˁ�WjMW��Dӕ��v�Rؓ��J�8�Adv5*UX��-�Uu+la�Z�Z��l:�	YRybי�����)%��V`�
�4�LT��^j�R	9z@��b��W�٩�U��ڣI�:�E&�,�kX��*Ե=ܖ�Ğ�w6��![wst\Z
�B��[d��Ĉ��Zi�Ѵ�ڂ�L��0��d(H��gS/%��&�Ts��
�*W6�4.����1>�ء-�*ކ� n��;Sbtf�Ҁ��I�T���`�3H^���j@�m ]ʳ��,j��{5]�1=Q��^��.6�$����*m2]Z��PI���hd[-��TV	��AQ<�Kw4YͶۥ$fk���{K7%LWcp���JV�M�7h��욬nD6}ɠTv���DF����d;U�	j`��C�4�p+з6Y�j���i�K%ћ6f"/]8�K/$�1��#�1��E�m�țc6
Ϟ̇T����k����&�(��52�nV^�of��i@E��)��`����:���H�4RK5�#0MQ�ڇrIUh^�ɏ,@�i�kn�k����v�J\�.�'T�m]�A �9k3l��`ӉB�d��ɷ���on�8�t̊oG��]��^�M+��N5.<�ܺd��Cv��֍p��: �c��)Ƭʬ��`��Xr=���.�w-���n�v~J�(�m����WT��^֘`X٠��� �N�n�6�ZMNm��.�U6���^Ҽ�l��J5��BU�i;�L߆�3fkEe�l*��dh-4��e�Z^[B�Y��m�p�\��mi�`�s5�A/ T���4�rh�8ƌ��x5,$ذ�@�i���m��6eN�]��"���[�\��z4��Zu��Ǫ�U�(f]��R���Wwj
�//T2C� )��e0��AK7��l�7n�2dᙚNS���&2d���W����T���~ �ʻ�.��[0e�ʜz��[gD�yL�Pi�����c"��r����	��`���WY�n�֪���F��]�u��:E�Ѐ�j�V� %=.�X ��Ut�ɒӨB�uit�X�h��i�:�ɖ$��͚�����؂�vVU��d9�a�E��Y2H�h�JP�Q!+�q���[f۶��(�SbH�e��2�w�t�b�`��Y�B�M֗{�5�S�?XxFܣNV���m��x���͡�m��!�F��]�M
�E[v1T�`6�'��4�@<ڽʙ�F�(I���y��e��BVS"S�0�\U��^F���{*%A�h�J��$n���P���G�Q��Z���1}��N��e���q�8�]eF�R��o�"�tŻ��Նt��=܅`Î�a�̭$��z����-?1��y��պ�� �8!���y���!yf��R�����]�! r��Q��%� %+��ѻ��rb�k~�e}�����A�EVV�i �2�9C0J1���j��w� FJy�)v�Ug��2,�dT�9�]��řl�R����`eYb���ప�̒�*@E���U�n���EtxrfU˙��z�ҹ�	t��p�/ig�n�Y��m�R��J�P��9�;ȅq �!5�* ��*,z�n�Ÿ�Û{�ң[H6��`�� �NIml2��Z�PҙEb�/l�Bmn	�V�KwS�H[��;�ƆFKܤ�,����Q<���F�0=�ٶ>�Gea�c܃%�2�y�z�1y�Ӎ�ϒn�ͻ��h˖.�Z�9Gc
�UEB2-��Uum��K�iP�i�@Hì�����VLwR6�l5n��e��6�*c�,Bf��x���<ӑ���!�����$1![1^\[�-ham[��OnZ0���X��Lr���b�j�\�Z�8i={�����"2VZz�eb�����\3+����:��xh�T1�N������Y�[tkN�A��]8���<ͧ�ef���U,�DlGz�l��>P��r��SQ��� `� s4f}�h	�^8�
��0^�iɲd�aƶ�Dʃ#��j䣨,�*�t�56B��{!�n+ٽ���D����G�A9B��r`�L;������dȅkw�٧��oi�;Ci%/6I��t�R�	q����ř`�YZ�QT�n7CN�U4b�G�4ib�r�1P�k�E��e%�K�]�Zv�sV���.���i��ۧw��斊+1�
$ l�n�ݤ���	8����TY':����0��0^e�WO.m�*^�SUڊ�=�4L�lQ{�.P�B��:�:\�M��^A�n[�lեr@�wZ�̴�V
xN�������W
�dդ!Cv"U��%Y �`��@��8�X�G��hw��:���Ue��K�����F�w�j��m��ku����@��6�tmm�4�a��d���H�k �)c�Լjf�-����h���t�V̀�NԦ������ifn�@=VP��W��<E��n㽕����Co��(e;lJK��Cxݼ��*��6^�Cq��u�	�5��c��ʸ�HF��2��e��&�*�q��
r<�(�Kٯ	��� �NS�i�#�.���ôqH�ո�El�Z�5�g4� ��4���)e����N�ݜ�u ��S{����2����2��{6���i۲	"f��RtT�3U	�/i�Z{!U(æ��jQ�	�v��hKP�
l�Z7\��B-}f\u�>9V��n��&*-Xjڙ�����J*ԕ�a%�!W1a�h�w*
*�$��h��ؒ<�����ͪ!�ɘTe��T�j�Bf:ڳt5�ۈT�HφE^����M$L$e�&�H�k��$�]��\hR��Kv����ؘ2Al����w��z�3��mɷ��S7j�9[����0���1��KV+,�*hGbȂb�B"�ע�ٳ��A��v�+U��6CL0.G�q�Yb���;)`e:懰�S#�%�����HiA��L���e�������dD[�!y����"�Y���[�sZy�ͽ��U93u�4�aӽaّ����FK�K&���r\��0l9t[*H�;��ڽ(�(���@�j�֒�X��Zr�m^�[Y�X���r���YK�8~1ʛ����a��DbǸDa%�2�݄ò�$ԯ�`��wO2�H��q���[E��wZح̗��f:�kl%5 ��Ҽ�1�j�,)`�n���f�!{4jˤ�R�0nk��lݷOh܂��J���Qb.`�u������Q;ӢҨmǄ%k/6��6-�1���vT@"�S��t@���UЕ�d LpԨ(`͋2��ne-���Q����sE�KjAy�����-� ����(j��i�G*�,�4�
(K��;w���w�b�H/�m��U�V��H�㌶���T�Y�
�֐yH7 [Wx��d�gvGQ��f�F�drkS0Y�c��bP�f�p+qd�gEcZڌ��V�����&CL}V��-�p(Y݄��Y�����U���h[,�d&�4bU��J��(�X���Yh�'������ٚ��j��77� e 51r��$��8(��	{h�T�#�yFM�z�mȪ��h�̎�wH�
�i;ݷ�kyDj"���b���ce�Y��r�%����. ��/q��&0��bD\B��w�#�U9w-k���`*WBT�yKtAjR��<��d��)���N�@XH҅c�ly�r	����Sl�N[{��u���T4m[l�H�M��y��4�6�v>5,u<�@����$��Q����r�$b7�o.�js^�m*�e�\�a���r��:%��K˻Z[�v��s[v�JM#!ylǴ+]]c��%[�\y6��-�Ul۬M
��bZ*�-"�\�w��Y�M��՝y�pŚi� �1#`�k	j��=�a�Sb7�X�V��9NrYӭ��ڂ��ܼ��g@e`��k&�۹Sܬ�Cuµ����A�U��aMV��*ͽ��u`+�Z\��ь���6�F*�X���b�@�����l��La���Eb.�J��׋\����P����R�ݣ������̴�($��/��J3s�
(Qo+_l�����Mx^kQ���{7q���� (e�{��]Lж1x�i�)�j���(�j!�u�i��+e��hǹu�K���x�cW&��7fh�bB�m��4h"�3c5��X��#j0Ҩ)�β����#���"k{7�9`͊�B�V�֢�����:��I7YjU���*( ���2�X��9�jԗ�S�"R����l�`6uՊ��x���fn��;aᑐ .:�6ٳb���3bۙ1��#b7����EW�ܷehNZ9/WV�&�hu�֞+�r�M���Yz�fS�v�g%�j�k9Y�ӱg��<T"��I�[,��t`%��ӷy�R�H�p���63vF�����wF}*��71f"� �D���h����([�}7dC4��-�S,Jש�	&��k���5<`��kQ]���lѭ�o�e`����1b{
`ޔ��]�%,�r�TLTC�����҈w
Wp�Y�3m�ܬu�S)n�-�I����6��Yx�,!�G��ۊ5oE_���8+J͠���:�Z���
�.�Ʃde%voFˍ���4V�̏�����,T�zbn�:�T�X�9Y�ͪ�%3i/�+{�,N�T�ZٔL��B��a��z7\"Oe��͔�ʑŗt�T�@��(D�G��0�0��0��;iY1Ro	�Qze�M�Q��*�aP"ٖ6�-UP���Ὂ����ه1�\_�cn'�'��v��u�\�q�8$����Ve�z�n�<>���7]�+�mbi�׷:�ls4��L�FX�'T�Fz�+H�ٶ��04���5*�ܣ|�z*��/V�=�7CX�>��.���ٽq���tu�I9-#Rҥ;_J�q:��ݘ2�>
�;;i]�#���E���0L�b��k%�-���@���s���"�tRTל���.Cqmvl<��&��1��N�=[��`J�բ�)7�Y0�wag ���)w[�����ʇ���*�#�S@�]�d�"��Լ��8��1�97 ����u�l��˲ҤO�Y*�v�n�"� �j4�w$��8�B8ga׸�=������\f�;��kWQ �U�.��
|��
s
qܩON޾WP�-7��kgήZ�ҟU�B������w/�n����f��WC�ѳ�npM4A�}F�/0�ٲ�K�w�΄G�.TYH:��O��mۗ+�'�W%[u"����w��N����6��zM�����;t��*�F7e%G���o�����*<�chWe��4W�:�*̍O9
0�\n�֫b����o��_pS]5�p\����F�;l(�y7�hQ�r�>=��e�� �+�S���׼8[�νI��8�)v�s]�;����c��#��}[u������~^s%qKS^������%tح�������x�#���z��rUdm+�e�2Uv2J͓+% �n)&*�7�u:�������'Pu|�ۖ�^-��`���ۛ�H�Ӧ5*���A����®M��g&U�*�o�������B� ��gg�� ��Vv��Z�%��ux�v�
b�`GV�f\�e9k�Lk'Re�W0�:�2�5mu�t�ݦ\Ns��''���-����E6**���8WHh�v�r���pW- ������\z^��{z.�n��-+:��Z�R�0�*
�]8�����$lv�wΊ��Gw ؏,��Zk����c{|�3��du���%���fF�J5����6���;z��V�<�[t���+0+���ĵ�|�]��[�1�ȥ��>��,w^Kc'O)-��*��]�����	��j��N�%6�Vɔ���̔�V5�c�@mA:�+5s�|�wgf,ۉ;#���[rPr֜��c�*�G.���C��p_��[v����r��G]���3v�p��Q�=ѹ�h�� V^��8&���T��b
�f�����8�л�&�bw�J�ܱ�<%����tA�8KW�
,@r<��̚��ޔ{v�T;{ʧ���:�v���Yv���\PZ}�)X2-�f��ڦ�+���uCI�B��k���P`��T�on��q';���c�6���R�tp�ׇOE��U����Az��:ɳ�\]>n�6�-����S���{Ӷ�v��V^������k�<���.�޹BZ``M�gtQ��\�)�3!(�c�k�gg��>ͺ��+\������QF:���Q�7���V���j}�b�Z�u:��N2�l��Eh,V�i�_ ���c�}�sp��i���AKt
Yƺ�����g^Y��F�׋�NB-�z����}$�C��u9��^��@r�e��P�L.7�u�S��5��Ӣ�<m!��+z�X�U���t纶NS��n�rWN��mZ��-�	��汕5�}z�SP�b����u�u�dޫ��m�J���y�jw�r�If�9u���5��v�ˮᢒ]I����hK4���2���"���z�W=[�B��9��X�T�
�%��:M=��s����V��mҩ7j.����{�tŵ��Ft�aaK�,.VPG���Π���n��R��yAd��x(�Pk%1�L���㣙o$��ع�_S��w��	���j3�XI�����~�9CGg�����Lp�2���g��sc�Z2����J�����"�L�{LVK��꽴v���SSm�3���p�,<�41�6��ʆ�M��y��)!p����\���dm] G�X"��;��Œx���H�\�Zt, ^�i��++*,gt}v�W EI*�c�m��!f#D_-���ALT�̓u]A�m��Ǵ�.��83,࣊�n6;Q�����D�?c�od�VwJ�֊:���c6(nz\�ݚK�q��ttMm�e�P
ȫ�Q�/�8�)Z8��u�Z�s���7�ڏ�u���$�W��k,����%�y�9�Ru��c��Ipm����fS�]ڳz��=�Nj�(ֵl�5�;��B��ݲ�!B%X2d��˽5Y�J�T*���4���U�{�Rk�grH�:��CW�(��v��;):v�]HVf��D��Y��n���b��Gv@B�u w%q��՚��%l$�^B1���F�Pݔ�K�:1�e<;�WA�kt�m�j΍�j��.����
�Wk��C�Sf��ow]�4��a�ʂ�8ʱ1!Z;�H���Y�bQ�>gw=#�9i�Sh⨰�-OyuM�\d$�B2R8�&�l�Ò���%+8��R��aɜ���
V���M��e:��W,����,;\��l_��q��#���'�եE%gz斎EJ�m���u!%�Y�o/����v"��}�����M���}����.'�!(��ٷ�c�������I��
���\�a۬�U�7�mcov�;n<Q��%-�}'׈��-t�ɺӗ�gosw�J@v�gu\J�%i<
2U��r�[�ilGB�g���J�q͇5�w�fs�v�o7��Г1�v���Y�K{W�Fs&e
)[����X����)�5�hޜMȸcKU4Y9N�;l��[Oݥ��@��è`m%sn𧢖[�t3vⓉ��mWW(�0ڥiY�:��*��4�o���jS5��e-[���;-���E�����0;�� �Ɓ���� [i̗R�2���e{A��]�A3��0Am�ӓt�N��eda-�P�������b�o٧9_)�r��ь%�7�o[��~��K��{]i�8'V���q��ȸ)�s�N�i�n�X�4(�{�e���Q��v���+0s���nԋ�-���V������j{Nk���H��P�1v�yӚ��~�F�p9��?�����l���{:�O_\��Of^G�"��bNOR��뎌��<�������yk{��}��]r�
�R�Zw���ɛc�D�[��r�1.�jw��cja�j%L���B὚�n���+C53˕��k9�I!�ׇ
-�˙V����i���n�"MмQu�����cRS�{WWO��E����>���)�s�؄�W[��6�Wo^�<�Vv���3FR�L�r�سWٻκ����Sf�C.�<�m������{V3 �S2g2�[��qq���I�ܻF�Q�5]:#X���F-��U��z%8�l���6J	v��/J���y�k�4�����o<�u�)oGP�r[�ܺ-�AK�tCB��3����1�E!�Nv҉�Sn�Gv��8>�k#n�쭮��h��ة�j6��h�WJ��3=��7x3��+��q�]m)b�^�cy�8�͒ll6�R�;��#N��N��)��Y<�U���=����E��rј��&^nW.��؉�R���F2q7���3u&��vj�x$�l��v���ޑ^�%���Wc��n�c��ݹ�	K��"�KLގ�s:�!�4��"�HKR�JW��+��]�;)c�{;�[{-R�g��l�b��`��GMc׹YJ�^�wRe+v�k1�`,L3A��bf��ǚ��|��v͘���g�j����q7�u�t�p�4K�-�B�R;��(�5icm�qD�*M�`��m���n(L��Ub>���[�pw4]�8��-��Q�!���}�MhA�p���aT�bn)��e$��_g^1��62�ڹ��*`��Vyw�FN�s-h�X8g�����mCA�ʩ9Dq.���M���F�M1:���v�c�4�8�˷�;t��ǔ��+�C'+ �9mv������f��
޷v��7`���ɻ������zrX��e�)g)��jx��hs���97-��s{2&*ʕ�[���+��N;�2�tc:�Dw�0^V7Ip��R��;;J�D��;靭�d]!x��=��]*�l�ӝ5m���]��@'H�����ocΩ)���=�/KoA�C��k�u�F�c���%���b�\gI�nF����$�>�-�v{������2sŐ��L�5o6��s}N�7�S�Kw^ݸ�(�gE�n�*d��wS������s�q��f�K�ox�,�C45C�C��V3n��v����lzkb�]�.�n&:eKޮ�kB�7Ô�:��B��wBk�ްnL�NB�ڼ6��%P���0�Ռ����}���x��{�&���;����l�=2�͏�lh6�,Ԑ¢��0���e��ǎ����\�A�-��}��)y�D.�YheqAS�$�*����)e�+���vZ[��r���lV3����|��ڲQ�%r��z�t�)[v��ڝ�"��.��әi�\�Y�Ylfu�l�@L0kX*����m������3	5�1���]t*'@�a�t���7��{���Ë�����wZ��vF���ɯ` � ��!�G~�]��.�,���GۊXpG3����T7k�d�"���a�D���h�Lykq�
+��%V��׽��ޥ|{"���VIJr��(��w�h+�5{�iV-�@���}��Iɸ��W�Թ���]V��vaq�v`-�G���ՀԬی`J_m��|)�u`J�=Vf8����ȩ�rW�wn��XWnn*m�f�2�ޛ���W|R�)��:E��'YY/h�kmkW�LϪr&�:[$��f�ǉ��U��!��N��.������n@��`Z�Oi�]@B�c�A�]��e�Zv-Ĩ��@Es�&�X2��-EȔSt>���E��q���X�i�5\�S��%˷�e���-V��W���.&Z�cp-�X�Z�M:|
Z�Υ�rNw�m����]�S�J�wt�z酓����v��9cu�([�����+JZ���.,�-��[���� m�ݙ�#�T�Nws���[/SV�]��5�.�Dc{�Z��Cisl�����*"Uj[X�=�㧶�f�=G�����s��	�"�F2�&n�늉�O(l|lD��ټ�P���R�����}h�M.�7@�y��G2�4o�y1;x��:��[�V�ώSW}h���g�V���Wc��qQ�ukl��r����O9��1|�"�q�dp��v��chgt|shs�r�3fjiL)4l��.�-�$Mؐ�*,N�-��d��˶���z�t�eX�1a�1L}L���ӻ��0����6q�f�!����Y�mB�']��Ѽ����%e.�sCV@�)J���_XLھ)9B_s��W���3	^�
�z��y��l*�+g@!O ����m�������wb�KfQ��;h��<.۸x>�ıcX3Q/;;jw
�|�s�U�b���aڲ73(W4SX�c��Щ�W��s�����3&�{�` 	lH�Z�ѤU<���|����:N��!����)p'��'�J<���0�{g7����6 (����+�N]��|��w�%�Ml���I������F���V����A'!�+,�u���V5ޕ�X�b�r^]J��ݘvt��[�פ���V9�����.b�ٮ>r�5:h�r���DMʜ�f��tȫ���W^���Ӏ��N�2	�m�L�c*t�����,�uG� �g�o>:��;ڶ����C���e�w��f_#��5��S�|"�/_o��ɦ��LK���:��]?���W��D{�b�uY�D��w�<��`��b���2��3y�s���.� �T�q�>�;�׽G�:z�kg�]+(雔),�L.؜{ҜAWt�&n�N�����X�0]�;�1Y�V{S4ޖ���
]�42���n;4��r�;!�&;�@B5����8~ޤ<8ӥc�^��c;}�4:�1Hl�˃�ޗ��{{D�Y��;Bq��i���غ����Z�`;(�[ś�c\z��(`��B�`���P,-e�;�t�M�\p-��3�=�Z���z�'�1ꋍ;�۠F�֤\𧋲�a�WX�WJ�c�'�_%0y\rX�M�M��БA�\�ܔ���U3P6+o:�ժY;��cLA�����1�u:�!�3�����ED��;� 󐔻uN�qӕ�1���pΦ4fd�{�K	GB�VS��BQk������Gr�*ew�
�v�lO�o\�����{��u.��6�t\՟�h��6u��]�5�wB����]�]����w;S&�>�0�a�B5�e\�´c%�aHk�F3���J�r+�m���8�V~ݻ�oEC�g;e��RXs�N-�5J�B��ڄp��*&E�r��x˭�9݌�)��q�w(��J���;x����狊p��{���;�&��K��f���x�
\,�n$��u-�+Uq�g�Bd�������r�[ ��@�43���hL�g��͓[�I�Եa�z�w"����:��XY���\�����/�	L���Q��+��؄�S��Zl۠�&��͸�`g�LFom9�������ܧ)�٦�u�.�ٸ	���T�}��;��Jٴz*���7,�ȸ�*uqżOR|7;I����L��e��ɮo3zr���ع��7wݫ�15�R�xxx�x<���=�J�DS�q���tf���a
j�=u8eZ̭<L�N�m��W!�U��V#Y.�
�ܱ�-���&e�:�\;��EH�J�E�u���n+����Ӑ�WV�إ�jr�%c����ǗTj��iu�=�q���+��>�>ȩS&%W]}�7�Hz��V�듊��䩷1�4�K3�d��Ŗ�u�NqQ��m����u���lWzTD�Z�e��=����s��䶠z�2X�jG��o����5W]��1��j��+K��3k�a�ga"5q�5)�vb(���o��wɮ�t� >��»�Q�ܫіۃ+lZ�ԗr�Gi*�t8�YJ�_H��&u�3�Y�v����e���)[i�Fe�{�z��v����;x����y�i�6ķ�Nf-�Ƿ�e/��	�R䠢$`Un�����K��t�/gvf�Fjpy������k+�ҭdK\C(L]چLG�k[���K/���vR��WM{�;�.o0^��vƗ�.C7�I�F���
l̨L�2�����`Ze���$�k��g")i�܉�'Y�$��nҕ�����2�|��DpԹ����c�Gg_g7$yN���{�
teӽ����Av��m<�Wa�����l�9D�I�!��]���R�O8�c�����z��E#�(ӝk�^G��q�V�����!�[��u&�����(����L�kCe���"�o�T�b�푓G'�y-�>�L;�A�����iҮ�o�u�Ĺ��Է���;B%�:�u�Z]o�����Ӕ{X��h˶���j���w^)m�2��;��i��
=��V��+w��7��n]�#B�����uةGZ�w����[7��<,W
�k�W�9v�A #,Juh���fLEfu��̰j*����{4K�sY��]���t��Ģ(	�{�*Y�v�]iWZ�w8����k�A�i�#�#��mJ����37f��������n�t�V��Ȓwxj�SxI�,�7�41�^eu�"m󕽨�B��yѕ@��@�t�7S{jS��G�Z��� 7��J��8]�\�Eޕ��!��H`9ml쭉����V�t��p�C��ڐ�:�0�WX0�>奊Q��U��F����w�*��`U����ui8���9��
��ٻ��ri���p���Va�^��V��[�����G���bTY�+��Xru*䗦���i0���S�Ut��:$�f�
6���}\���f�F��]ٙ)�Ͷ�y9t�)��;�	��h��K����i�vfn�9+�	���J�(�TՠXY7PYGusԆcZ؈��LQG/�֚�э���W,��\s���dڍ#�n]��9�*ХP�1��ј�C�v���n�.+�Y΀V�#u��xˣs7-w�|��x0���:�}X����=���
'[�W�F�y�.�����G.*d���<'3�vp�٢�d8*\���P��rU�w�u��6`�;͗�B!�N�a۠j��q��;;`E�R��o5��v"���l�j�v̖j���K��FS�k��̝{.O��B��@�A�����E��\�uFH�jr���_�7,#ՠ�E쭝����6�g׌HEN��6��C�u��9v�mu���/��^�U��9F[G�^^�N=r)$	qq��k&�:���3�J�}���#�{����ѧ�]��O�{չ�y�(N� %��B��6ٸ( ֧�Wv�>�z��f6�Z�u1�wd�/��]=j]m:ԑ��Y�a���)��냦:��Lf��R�����0av��|{�R�ꌖ�X|n��A�s��Ӵ�7�w7���R&D{-WEN��ӎ���vu��u�u��`���S"���O�Y7%$.�y
��@����Դ B'lώa�z�Eljk�V8��
s���%Ep76�3��:Xuen�D�P�N^A�V
���a�} ��4N�e�e�N��mfQ�����"�^��]����T�b���f�F�VT��0��xSms2����J��уM�u�Z��2�r��j��)S�p�'�/����T�Y�>�:��JML�k�1�{C�����5ȯ��U�m[�p���2QO2W2;U��-.=PZ�R{l(^3@����ufSĒ�Ґ#st}un��^NM��y���w��|4��9ս�nSkz�Ut��i���0���
{����u��k]����&�2$9�Y`�E��Dϵ�+����!�s�c�ӵv9S�2R���Ds���np]�v�xd����r�8�돮8��eD���;��I�s�{/��Y����7b�R�3���\�s���e�楘!��!܁�#k�ɜ�`x+*U��{�1֦��J�G��]���)v�����5��LTv�;'''1��+k;5���^ �)� �ݣ6՚W]�4��	�[�\j��V����%v;�X���C5wG���j��R���4�}`غ�X�K�\��w����s �V�^я�')��bL�;Q�]�-�Ϫhf�ه�-�]�"A�Ĺ`թ!��Z���ky��Ed�Rpfi2��v*�2Z�=��i>k�+�`��B�{e7�j�;�5@ͷLwc� #I�5���ϟ�3��.���Q��A�c���[w;,�:�nY�L���&
����z)�n��L#�;(!��s�1s�M��\of㐮�s���3B�We�����D�C*��f��X�<z�Z�\�ְ�ν���jܧX�ӱeBW;$m�@�ReI��mˣ&R�(j�n�Kx�5���x�Z3/e��-Ā�+l9��c*G�T�\E��!��C;��nAdW6��n:j�ǰ��f��APv�}��iR5��}[ِ�R���b}V�wl����-R4$��-���۬����*mNX�,�6���F��L�Q���{L�5+��R4��%�x�`�Pa�A�s�t%���_[DڱHVmf��m=�6Y��N��ҳm�#�ۦ�K]�i��,m[�ƟCx���VZ��T�W�]�7*�0�VRɢ��Fu�J(c�;��c��$_MR�u��0K����#�����^^��m)��%���/o��nu�)�Cd�7k$�k�Y2�z�c������R�Γ�9�C7�صƕY��gh�)���I0C1�Śy��ͤ	��1��]�(Rz����M12���.t��h�5*��ʟK/�����LR`�Q�q*�{�7���V��M�H�W6�� N�EG�;jV�%���!��\yrd�2��&c-=M��������)TYǲa4-��C,,h��./���3�k۲󑗖�ɷ���;�5մ����� ʹ��XU��ZT�2�r��xLJh[��{�P�4g9�Cр'�*S��䶕��N�Z�;z�����	����R�*�}ۆgh|����GMDOg�5�k�Y�b��u'�<�}��lQ<�XUy����+[�V����J�u��&-���ʕĬ�UoY��o30�������V'<}���Jvgt���Gu_-���ݎ:�tq7�����q�2�����z�$e�,
h�Э����.v��@�ـ�O��+�Fh�^�vj��8$���I�&u�(d���`�2�`o,�$��9'l�e�J=���ap{�̜z�zd̶���P�RG���A��9cQ��5��u2b��^�t��׋SYE�6�b��֍'\M\sp`�u��b��	�Q�Kp3���Rs^��sUrz�.�tDV�Q����Ah
p�3�Z�M; �zWK5������G,�$55�PChv�����J�sp�3t ���&��]�@�5r��:sV�+:-pS	+2�M����[���x�wk{�����f+��v�9ĊKs��V[�C�ڻ��A��3�GP�o���s��,���պ�5�FKYMି�헚��0֛�\�3b�����d�-ZVS��:��nF)�J�X�w�@:��K5��B�]Zt�]B�������u����=�6�s�٣`������vm�"q�k ��P6f���ܷy.�w��bO��E��`{ʶ���g��Mޣ*%�Ela�Ր�Iޕ��R�^�ƀ���b���%�;���dY�(�1d��|�&�_.�n�����smb�R�nS�og2K����e�(��=��Yc���ù5��r�P�
�Q��5��a�9rj�6)ͭ���qG�u;�\�)fp���aR�BB�-Ӂ��ٳoZK~����}/D���pS�MN皖r��
�]�@���j���`���V�Ģ�sx�/�SY��!Njge�:���1H���v�����jJP�"�p�q��xe#\CZ�HX�p#(����3#1�S�@��.���f��wr�J��Ҧ����YR�����w;�@��4�^K�v���u�=JB.��%�y�o/���xc��wA���j0�zz��\>��d�}-Xl1#'�N�ki>�H���<��}�mX�S��$-5�	��̠��U6���į�|YZ̡��U�)wd���S�eU���Wn�8�'q� �}�p]n���1kw�T�-��W(�A�TkI�������6K���(V2;[`�p���;���[�^Jml�o��)9�8U�޼�d��ܓ�+^�j�:�ʾW]�\�n����7&��G���6�xJY+�X���|S�Nm���oL��ƻ���R��PE�Soc�;Z��\嵪�r��8�ǝ�����l �pes�nXY��Q#�˰۩��u�^gҭ-1�4�h��b�o����=:R�q��L�ujv�]���rL��΢��.YfJu����%���;�YS ����L�T �\E�G�+�,�FL��s�}rrZ��S��$.�iX�;��2�n��xP9�/�Q�IB�U�I�^�ܬ��X�N̎�l�:�I�G���]IcFUj����?��f�E��<��Ck�3F���K�������E@%K��*��.|�V>�0*���!
P�f�I�qB���W��ٗ���΁E��C�[���:򝆎���.�f��U��v����d�7��M�P2ƣU�#
a*�:�^��Da�R,�K+���ho�4]�F#�Z�Ȑ��7˛��*a+&�脌�O9X�~����,b��+[��0l32�8����i��%��\x�<�q�]�CI�X4ʺ��3e�-�=sIQ�n���ڽ|�=����5x��L�gZy���c4o��n�f7f^��0<'y��!�W���|���Y����|l
t�;U��:���Q}����39�Y�Mn]-�q��kzp�Q���k���J�}�*m󲌁��4`�9a�噖ۼr�%����0E#/7]�*n�I��o�Ɣ�#��>��YLܟ�kG^Τ���I�+n�6	��1MR� n����tE	Ֆ�GR#3f���Q���
2�lT��w�](��8`�D�Ӳ]��{D�v{-�F�]3nN멮�f��m�X�O%�ު�ʽ\������V��"�� �6\/�#�B�Y�{�n9���
���@,�<���̀�WZCmk������U���ugi��Rnό�n�Js&v'uh�Ջ�������Go"�Ð�r�+�I��z��bf��
��<�Y5���Y�R��ַ��`��������f�9q�۲3��N�
�jU�k�A]�d@N�*ڎZ$_DbP]�Yv�

�b�ُ�핖�d|/eh�@��Z	�7Z�[Qĭ�A�,�N��@e[�1���oY��Zou��Y[�:���k��^��&�_Lۡ��X�`RBX2�k/7q�[���h�9J����@��7x&o0��d͐���YJЙ��
�uj�232邊%���{�-Э�@r��s����:+6�]<���o�=����#�}aC��釵�V����)�*4�����X��ݹɵ@xX
��@hv�MŇGZ�iv��mM��*�a�V��]#��"�g��C���}aIuُ�)�i(*uG4>���^�}��Sn���r��\�6m�K&�z�F�[�IB5>T��<r���� ��XF�T���hnV)]B+퓖mb�]��S�F��+Y���J���s?`��u �_M�#��6�3p��Q�A���fv���5%2��g%��K\5d�ͱ|]� "�m��Q���{���ܧZ®�����'���B����j�g,�Y��ķ�N����u>�i��io[fn��%��U���v�[��N��XX�7]���8�u-�8۩�pK��ʽ�*�妅�k8�|eu�d�V��p.ʽ�+� w-��(�s���z�Fn8��bvs8c�ge
h�}�� ��a��3:�z���Qs{w�|����Udt��U�&�X�K%i�u��h(�e��q�t'!mW_@���2s����]���	�yl9�*���j��(X���lg5l�����OF��}`htH \�l�.���<WE�v/�<�����X�
8�Π�UA���ʚ�X�[�X`t�N�X.Л�oi�v�S;e)��q���~�/�弇nn�}h��28;]�W5R�U�����*�Z6�[aR���1b���_eo�@n��]��
�bɧbe�kV�r��0�k��1�v���rY5��iS�.�jq��[��vy���۝�����E��8��7��;��S��RH8�ׅ�Tw]Fv�hV�]�˄Mc�	���Cj2�4#������(��b���+TՕ�Cy+�sљZ���ٌ!+-�ww���n�>�i����$�	%��f�x�A7	{�RT;��}j(�8� *_NA�+��9|A,@��Λf�[�Nfj�:�D�]g1�}�ޮ�]��ܡ�n!*4UD#F�</��H'�����b�?j|��8���aw���"ܽ�k��jN���:vu�,b9ɪ�3*�וw����lr�Z�w.:j�ٻ�$�!p����G��]of��-�#AU�:ygF��P�'����(+�<�㻚� ��n��h㹽R��ˀ.�A��J�ޭ��]���6�@��5����v���=u��↗��Xm�<&_�r=:���؎�x�z{9�S�۵�1*O;'RJҸ�0^�Kv�h��{gЛ
곹>9+�gv���<���� 1�uۥ�ݽ�pk�SOl�P��	%��Tw��d�i�ە�&b*�j�hlI#�-
�>���WB��NV���Q��˓����i�\7Xx��7e\���xܡ��p�;�������$��¬6�MRAh���Gvsv�s*�}��R�[�LI�Y͎��T#]�a2}�h�F�WX%L˜�.VV���ޝ�Tt$%�C4+�ޱ���F�i۽YV�i�}cR��t7���"F���.*ޔyŧ[݈��&�����}ơx�#އ�e�����7�ϧ1�j���N�up,�Բ;�(>�kL���1hB7��eӎ����V.�M�ZzR��s��Ft���oZ���ᒕfblPܩG`�ޔ�eo۟]f~�����"�1U��T��Ue�-DE�"V�+F+	Z�b�X��E�UR���V*���+
 �(�*+Y(*�J�b#E�j�aPUR"�""(�"����VYmE[j�Q���jP����V(��(��Պ�"�[�1�**�Um*��V ֩iDQbEU�DT,cYD�����F��mR�`�b�QQ�E��ҴDUb ��T,DQ��V"*-IV�e��1�[
�*�D��U�,kZтEU"�kPE-,T�UT��T��Z�b��b
"��1E�UX�D���+*[E��T+V �����h��P�UTDTV��*TVZh�*�"���b����b#mQQ��ZX� ��D���T��%�DZ"ҥKk�c-��(�1m��j1X��T`���DQ`���B@���I!&�	}�9�}�Į_�]��燢]XE�\�z�1pk�����It�Zi��P��Pຽww�t��I�v����2�4������o	V75CL�:��[���i,�-\�US]t3�hu$�a���(*�Q��8� ^Ȝ�܍��eW��qeF�ށ��Υh-Ļ��Q�«M��>���
�)֓�рp�Q��3�®<U�=~�6��2�C��w^kX	���޶��Z0R�1e�T�y��H��b��z�p��|x����n.�*��z̾��[ؕ�D�nl����G'J�U��)�Z���=>���a����,�Þ��R���Ȝ�_.�e�p� ���P��rϰ�(���4�n::���G+Z�Q���Ra��@�Enθ*4ҿS�4K��P u9 'M�������\s/�ϫ/f���Ȧ�C�����i^E+�=T�-�$Ď5��c��1�tЍCy9�%:b�n��qMI�uw�*�4�7r�"���$�*��Q�i�	�=�d%(��Zy+$�ؤ.�S�Ш��p7
j%�,?:~(�/�ѱ�.��b�J�BT:�֡��!o/�!C�.A�c�[���������Px}h�2W��V�RoF	H��KJ����/-����l�`�}JJr೬S��D�=6n�~��O�}���biGО�{���C���ܹ{nwd�鋫:��<�p�bK���L�_���;����,<R���0�r�;W��B"V��CF���Y5ʠN�/�7[�G�+O��ӓ�=����2`��ȖmQ��Uv4��U�sQ"�Op�>a�ty��*y�p$��.L��׶Arr4���Z�J�*��O2U%s�ժ�S�3�{#�g�r�P+G����>g��_xT����wޱD(��F2�2����zf*3Э^�<a�ih���uX�׺�A*�v*�y�տv\�f^=��9��s<�̳ta��t����Ӿ��H� �S�:��G�w�y�w����Nf�4B��⬰�/�-�/��cص̱���F� ��J�E-�����.9�M11+g:N�c]zCR�9T��3�f���F��J4+k���q�f�
�K��Gpp*0����tȳ*B:G!�Zs\�AԽ��PX������Q���\��~�+cM\�\�����������˨Ӯ���g-;㚲����ڊwҤNV�L1�݅�6����ey�g������\Z<�XP���ߟ�%3��t�ҕ-��X��9s2Vy�VYc5�f3{f�Q˃*�I�Cw3�p�[�ֻDQ���o9���,��2oc��a�9��8���<�,=�r��gb��+�˲�sk_b�����8��+����wn���S"�Us�j6�+���a�\9���n2���2���)ר*�l�/,uq�w\*K67���>h���\N@�T��Z�`f�X��wG�x��P��8��<E/���v�8���J�����Qt�Q�	�.�*@&|3��7�����n)up�ѻ��4)�'�=��ͧs1端���!~��x�>�3��d�|"'�^q:�rj�����r�O�Ƥ�2�5y7yqM*�{ZDT�%�C2�W�g�a5������*�R���.�6��h�2�~�;��c��x�TΛ�#a���Rsb�8���6|���6����e����N�nR
��x՟3Ly¬�XU���4�vra��q\�F���n�OK�9�Y��nS���4mX2G�J+Ę�
��*�Ĵ�/��������"�zW$�͔|�'�s����EVy�;1�胧��N�%аE(F�Ez�Ё�]��g(Y�ޣy����U��<��ބi�(F�.��X�<v��0w8Hݘ��_�U�=+�h�����­G*̢�I�`���RE+���	&��k��C,W�D�S����틫���V>���ɻN0�����oWG���̜�w�Ri݋i>9��]5b��k6t�ּ�k��qw՜w���a�^��F>�:x��e.|�'�YM>�:���;%^���b���6����T���-�7IԨ�2	��雱یrv#X�������3���
s�%�<������5�OgϽ�>���U�g��TC�/wf��1���{�s�	]GaL
g�tR>��W�)�֝Q~](���j�Q��eMo�YPN]�\m�O�P ��,�}ԬH��^�9����2"
2ov[�#J�s�w-��XsVR�xҧgb�^V(*�Ϲ�<W�T�+x�h�B��BhK����a���ђ�e�&��ݑ
S��e���F|"���9S�&� -e��q��u�J��u�	�	ݘ�7�OPnrn��nQ
�k�m�bS��.�'�e���vj�hN���ó�y��Td�,�����0X*l��F3Ė󢸃�:��"9��7�n_6�UU�`�a�0jcY�[u+�U���.^*�A��Q�s5e�]���r��s,o@�P�O	GW̗Պ��WCa39i���b}�u�{�	�=ۆ�	�4��ױ��2��{�L_�������-ܺ���1��X�޺�<�^��S�E�Σ���5-��\�Ɛ:�*����b��m�fE�%�����:��O9���WUۡ�0�_˧#r�8���q�o��=��`at�3[L�My�\���:�cKj��T�׃K��'���l��V�<&���=%��ͅ7ϭ�Ը��Ev�p9Ѥ�0�X4�m�]��
.�xΗ*����}M��������;��u���Rh:�{;f9��e{6QI�������݌|�+��gw�dėD����w��z
P���j�iуF�U�=g�{�罓�)�i����m�tGH�qe�=y�Qי�L5��:��-E�.B H�<h����˯jV����'{A��փc���q��<=|l����`��I��h�5�9Ety_�q�Y�%Iv�uv�6�w��l�/%��w�T�-)w���8�2,�)��Cu��T-PG5���Q�ֵ��;�|V�^E����׊�D�)�WB(P��y��|WLsR��r��h�Vxǭ�MŌ�!�X��]���N�Y�f��Pl8�}^�Q�޹"�	#^y1�ܫP�K\s�vƸp��N�זK�-:�h�	Il�ap!�i�>����j��B�3{vBwL՞��?3�:���[ ���wAƬ[�>,7�ؕU��Q����Y��z.j�O�MP���H?I\5���9�p��ޥ����y��rg*1s�ḳ�z,���#Vs���˼�0�]ݎC��S��b�:����q�����xLH�Pخ1��j�@Ћ�{nۤ{�³�gO�Yaf(����`ZʓC��T>�4Cy�]�83y�1m<x�3�Gb�q[A?��*x�5��Ͱ}f#u=	�ǲa8��y�Zy���T.<d�qJf�ث̼1&�LM�8�c��z0Di�Ƭ�绋i����j���t���̔Eu�&�:�7ާ�E���D��ӓ��b9��'37CL�F�*�4X"��6�y���gG��T��Ÿkۏ.L�ן�B*���{�����0rġ����/�E���Լ.b��I}�����/F�<�=��)_���d�ۛ��#�æx�[^��.,+U����|aœ�V��k�Lk�u��&�n���\�&Ʈ�T2��3&�G0���A�񍋇>�4��K���`��	�<ts�]y���[�������J{�;u;��R�:9�(��V��Z��F_/���y��X�¨�[�m�b�|��Y�xk
�Ó��8�Y���֕=���*Lkp������]�fZ��й���N�z�.MK��tT$5\��^�=s�嵓YyC�G��uٳs��gE����c$Մ�,\��z٩Օ��e���òTX.�+i���Z٫�wL-��	B5�a��W��!���U2�,�Dd+����P
t(j��qjy�q��r[7@���*K�/��p(���X��y�u3	ĔAE'�F^)iOy[����������8Ɉ�F��t�f�4�*�i��h�߳U�'�G����/'� �f՞��D؈��[Y�
�x�iG	�N;q��G�V��������q9��zj,�"�}JV�v T[�!##j�e@9fM0����J6�2�z�]qsT�g.y5;ymC��E���gE�f(t�>t����*�#g�Ϯ*"�Z�o
tJ�Ɲm쬌��yuD��ڀ�^�K�KrJ �7VVZ)��3��ù㦋סEl�n�Q=�8,����A��蜚jt����횓�z�N��m7����籾���(�Kfgs����n�Y1S�K�������{��,f��6�]sr:٤,��҆�Żܛ���Ç������idd��uc&��{��� ��C���8�E�DZOȌzTh�Q	��:5��:��ҮV�������m(�q�R�,\d�xn���%q�V0��{
��PO;Wd�+�@�̫�M/���}���)�ˡ���FZ7�~5����y�Ԯ�ϣ܅�f�u/������/�+<�[ ��[ћ���U�n�+��w�:�Lz��sƬ�;�eՌ��_���n���H
�֜�:J��Le$��3Y���i��)KUc6�������!�f'G�K�׍��&^���ѫ����u�"m�<�ɪ��ln �"��R15<5|9AY�J���*4:cC}���鏺!Y��u�PP�#NP���(ӕ�A��Hݘ��kwn��cj.�O0���D�X���F]F�x*a|zVs�yWa�)��39���2�?*�����%x�d���4ѝ�%OH��]t#^���qB(׹����q��J׋eT���w�Je���-D�xS7�]GaeH�D��Q�<�Ν)�֝P�L�#�n�A+�[h$����Y}��w�t2�a��Ҩ*,J߷��xц���o[��-�]�$�s|���+wB+ #�]ei��K/KYO���>�^S
�2��e
u�P�2���ב��S��N�(��Q^y<V�\
*��MC��9�j��f���2Tѹ������r���Fh��{vϘ�|t,5ݨ�JX�Z�wE[�+�V\V�V��|�}N7�,��q+7�X}K�m.2���S��6���Ǯ�W�؝]bձv�*U�Z�o@0(�V��dS!y�7�ٔ��|3�;ko����w}V�2C'�NW��R�U˵�^��G����݂�v[�1#%�iDm����&=Ŗ
5Ӯ�E��$��eϦqn���]�;�z�V&�X��d�<?���` dt��0�ϟSd�\@�%�g�K՗J�� ��qu���6=f|�E�62�i��.�4:�3V:l��(��x{"��{k��4p_�Uo�C�I���>�5.��u�A3����
�{U�s��#�0a�������H]�ET<��zﳝ���%�hV����^F�����x���we����=C���tjQ.+�X(�d3mA���X8�A�4�[����wX��Bأ��AmO���!����MP��t4�uwƶb{�V�����^:��x4��>0yzb�>���Qxht:���6�>ݝ��5�i�|bў.��_U��
�/���bz����aЛ|������jx��lw�E�5+�̏�B�cV�Wvޣ��DQ����1���4#��}Ӕ�YN���V�^���Mxo1W��s�kv�+�u;��)w�nEƤ��[� :!�,VS=�z���i��/y���W]�u��-)k��y���0v�&3�\ϛu�A�C�O�������^���#ό�
�5J�f�բ8���aY����{�M�6�ᣅ��i��(�!�q�(�d⠌�<�\�7��2�F��H�(�����!vFn��v^⫶��/!��Uj$�t���##rt�u\(f�<�ճ�v���׊yo��^����\���s�:B���[�ӗ)�8Y�f��Pmĳ���w��%'���6T�70�k�1C+�
��ȑ�:�]F�WN����Ө��.���x��j�A)��a@؅>�E{�˃1�<O)��a�5Ѥ:����CY�+wx��|��Gr(V1�V��*25�����K3e�a�4�d�ǔ�`1*v��+��9�M���[�`+զ�*=K�+�-��?k_��V}f}E�r��i�%d{r),W�Q��u0�kniE56tCqNf�s�]⚳5Q�y��ӆ�J�\�:X�Ԓsu*��ݪ��4x9�k�Q5�um1_$_��Dg�83�ӗ|@C�Xl��ح9L�W��\ҭ�=�#V`\��؉>A�ty	�O Xqn��u&{=�.t�<��!M^TB��[[S�l����0�I���_3�si�6��/G(���͵����F�o<|VȂKE��6���V��A+�%�{:�y���ʺ�f�t�gV�K�xS�2K]��َв��WB�W5M;�OM�΀t�%[��빝y>����J���X��"��q�[C��ю�ݼ�u弩k؛���lv����ȓ�e��Xi,���@�xMk��*�ފ��,�(]�Zm�b�����c�d�9�"�S���u���C�f�媜9�-j[o�q1�$��u8fU�-�)4PQ�d�
l����=R�k���`Q�|����u�h�Ǫ��tL�/�pWn��H�[~h����=�H��Q��>6�"�N�r��A��nW `�+���Y��+���	��Z��fwvԄTT*e񓺁������@����N��IR�>K�$iY�c���[V�b�Յ*`�)����v�6�a���R��]�.�U�I���3��DQ�u�Ryʀ]�/����s�xߞ�St�g��X��WO�؇6ٝ-JU�0L�>@���_r|���l��c�����O!�{9�Y�#�s[6�mO�٥�9��y�]� �$C���+��ٺ:�L`��
�IO6ŧ�f��%D��e]f
B�ܽ*�=֠�����b������8��8�i�"��9C����/4��V'H��u�$q��kr޹Zgi*�+�M��R���HE�����]]��v\]yVP�s,\t9�)|�[x�[#[)�Ux;���-�y�y��rBhȏ;cel�J�k�HFJ/Nf���cl�!u^�¹��N�K���p�J�bmM��$���f�F�U_M����L�/����BG�oE������J�SZ��G�7@�v�Ɠ�fl�t�dwPm5��8�|��,��me-ţ���g�wwA��G:R�opdbY���L	_]�o�=��O�����Eު�A@��K7�֧����%��C6��u� T���_\�AN�2�\o_ �Mbba�#]8�,=�,�.�>�fc��I5�jȚ]ѽWՍZ��'|�%�f7A�z��w�f^7�H-�aUrX+2�剁ݛ
�t��r�f�!�4yA#�iTy�=��Y�b.���5ʋY87����]���.�s�]�kZ˗h=먭(��f'm�(ֽj�=�Z��]��Ե<���Yn⏭XN�/���V��'�-������ߚꙙВN�β���il����=u�f�L��Ϋ jC}(S.b�!���&:�f܂ڌ�y�<�tp�y4�0qΌ��o\Z@�\{��j��s��l�2a	�rcfe�O�a�޿���3��������"��5��DYJ
UҥlTE ���A�*��eiR�mF��dF�E��
ʫ�*"�`���YYjVYQDEPU��+ADDe�Q�ڵ��#UE��j�R�ZQZ�+DE��iZ
" �"���6�1ZP�mUTE

����eĩF��db��TURҤF�X��\�ii�L�"ɍF(��j��R����J�JV�++*--�er�Z8�)cZ�A��
��r�,q��PAkAF "
���j�Kk�EUX�V.R��b��Sc["�UT�DAUAr�TT"�,LL��DV9j��a�C"���b �h(���F*�(�"+mV"�"#+*1�fZ�5��(�~>����G��Y�F�W�k��43���m	���o#�	�m���QӶ�p�k�(DU� nԝ�e�������Pڮ��u�qG����ٯq\f���8}F�	g,l�U�&F���U��,����͵��@�ý�J>l�+�;������o�W	x��K�ݖ���^���C��g�VM��i���x����f���t�T��0N�"V�\��QX��pf{lw��U�3��q�ʡ�`��C�#��.�U�"ĵCD�86+6�j�{�uq}�t��
�J�k�5c�K=�� �LK��U/jL՚����ٜ��t��L@8S��N��:�(�p�0(�v֚��Xm���qE�øn�,��׽�15֎�I(�s�.�q�'i�6_)3��2t���g�m�;/q喷Aڸ�����Bp�3)|{��*9�8��n��Qh��,�,�}�g�mx.�0��GTX�`��j��Ĭ@��8�26��z�5�i�-w�Ά�J��#���֩�Z�xݷH�E���Qrr�Җ`@ҡ4��,N�d:����
s-M�u�JJ�����x��+����%B.��NҬ�o�jӒ)�;�`v^��m�T�J[�<�V<	��o/!Ȯ�n�<qW"9�.�k0ʏ�=��w�^.R/;�ӕ�����V��i�
ĒoqYmR��6���=���{sLb����{��{��D�1�7h�6�Qy�%�'�n�vT�L�n��'')�Ԑ��b���ft�ܢ}0@�}[���k�����hUqXb wT���*�#w$���L��^��y��a�0�cp�����z��!��!�;���a�2�ډus���Qu��ňn.�Ңa�혁��F���ݍ���c�է����lUF|6P/��Gjo*����-���(?���ݎ�nV��Hz͇��*�A�4��Ƙ�z��r�H�OQ�hÚ4y��{r�:`�B�;e�{lf��^�<WPo�0���\VΕ%���m�@�BJ�I�ӭ�<��8n�A�b�)yԡE�bX�G{3�U�E�zƥ*hV���;"�ίH�aCq�E�E8O8�R#!��9aK5F�^�&Ft�cryw%�BUAT�W9A����Q�4�ǯL/�L�[�]����2bH��9����p~l͐N������%OH�n�����ܽS�F��G��V�!N���5�{�%.3G�^fŜk�� ՗�,�mQgJ;�mnS�{c�ř����,�;~UR[���8�'wm���"�o:���7�E97��P�Y[DU/�*Xk���
G�7��*�h)�;���b��E��2�� ���AItsm��9�ٿ]PP�T�s�+h�,��{%G����:t�fP9�$Y���0������ج��y-�;�ኁ@nY�#�HCϻ]T��}"� �'�%QBѷ{ى�J�p��0�H�˯VV����<�j� U��S0��'�ul�q���j�ԞؽS�<*!D9�AX0:�%���\
*��f*X=`r�0Mp�
�3(Ȱ�k*9w-Ǥ���ֳah1r�S�dxV s�뀮��,v��T<=C����\>a_wtV�cT;E�:5B��L�[ a��>����۰���R��|p2A-׺+����vz�e^�LgJnӿ3��ᬡ���o��>��f
Jo銽��&�~��Э�.��+��T�"h�`���'��q���zM��!dP3�eU�&�L�u��on��X�,��s��D�����	u X���u�>�v�Ih�@֊���ב���hl�=�9��{���T\�b0O�t�9~�d���X4�vE�(���~z6R���g�F�L��J�bZ���*�7t+����b��\Pv�9�;se�¹P�9Һ�ո���T�=KJ�)==�v�m�3�c��쉄��$�]��������o9���˧��Ƭ˖�qE�[�T����G{s9�ꯪ��{�����ۂx��ȀdR�0�`���q�(#��O��X{�MW�`2�<E�'����o0m��\]�^�إŏ���
�C��Yg�=�>���I@ّa�U��s�9�Ne�`5�wW����G���:W�@�R�91����WB�E��Տ����pK��X�����Z�Dixﻪ�§\h���z���e:�b�Z0{ r��pf�����ōf5Nx�⎖3���+�`�
��#�a�
F�O�s�,D:�KP1���JWk\��D���Ʀ,��^⫶�׋/c�M����=�ȡ��m5�:E��6O!���)��T���U�0�
��+%�k�ӻ��3���IL(7�b�,3u��}YY��]|���Y�1S��Xb����#{g\i_�ޚY,k��{�����\!�b��V��S<ß[�"�-̲
�]�U�cn���֜�c)*;�)�t�m�}\8�Bt���G�*5�4���\"�P/Ec�N������͕٦\;޸&a��jR},a���Gͫ]б�A�<_R�t+���񊻂â`��ׅ�jk�n[��|�1�����R�k�P��A�8])�S��p�g+z�}�c�(v���G�/�S��mK��fi8T���*:�,0g�+Tp��g��< �}��Y.Oo+��9&���#>���Ê��}�S��EY��[pW+���@������js�<�.�~�^��Px!8�3yϙv��;=;5fm�Җ�Y���s��t����hu�9�s8b�T��NC,�M�"w�R_��Dg�83H��G�lW��yv����{����j�W�Q\�"M��>C����ŸgFY��ݹ1��+�\T�,����*�}F#M�,FϞ��2��;?@��x^��X�]�n�{x+į;����R�r�>��qaNK��p�U�V�8[�H���"'F�v
�Ӎk
o'z�����-���<�ذ��j���8��`60�J���%ڂV�.�y%��tԗ�O�_�y�IWI�=��Eis�%-�m�����^���役�qh�{�9�E��`�0۟"�7i@G��Ҭk�5c�+����Dd+=(��B�Г�.����Jf�/@LC:��&��1iP�R�ۊp���5��{O�ޏȧtyY��^��;�5X��K��޹H9	�Ž2��Ρ�L��7��it&hۃ��-Ԥn6^����!�Ī�����nXjY��0TU<̊[����a�'�)=��jL��@lx$v�ױ̃�Y����o���I+o3�u�ѻ
V	D��-Z���xf�-H&�b��U��(2?z.r6��r��U�1(��R,��̝:�ʽƦ*������Uo��yP' �+�YD�����B�N�g�#TI�k�hI����%߽E�|��f��f�Xr��c�<��c��������N�K�Wn�:�f�J�h�J�����0���/�)�4"��,�j��U�J�כ��,N�d:�q�x�|!Ԟ�i�'+$7����y�"Jq��y�<j�]�T�L�n��;,�,(�J�Y ��0��nP��Ȼ���
�d���^�ɦ�N(̾1w9.4#��	&祵������j��]���WiS����]f?��U�s��9��C�r<sMYU��Y��J^��Wi�}�VMl$!n�!��^�%n�=*�_N~&�TV.��q=�o28oUN.�\�QVn*�]���!P�R�q�-�:�K��f��Y�4ǜ*�`�����r���X����Ɇ3�X�ݷɪ���<�d��|���a����K"r���ӡ�:�-���ʈ�A��!o]*�!&�}阀�bU(J훴a^�>*���𱫏P�nH@�w��jt���Ʋ�9W݆����+�3{J��'T0�0;s�n�]�?����k�ޙɍ�:�ҹ�W[����{���r���1lU����1�R��_K��z���/�|9J���N��+���g-ߊ-irv�WR�B���T]M�F���7ӎ�h�[���ڨ1�҄pK��v�����G�����lLb����(8xp4���h��Y���g٬u9�T�[�2:76��ư��]�:�N1ҍi}Dl�%Uu d[�n�wB5w/T�
DC�i�LOr��ؘ���e��󰛼��]4W�yxS�cyt*�b~u<��{�&p�����b���(�w\yC�G��t��T-�0�t)�W�uR2)�P���nm������&u���n[��^@����ұK-�d	�J��,�[�h�i~�z��i�;h��`f�z*!�j��0)�{rYyp(��3�`��0M�@@�t�n"�>{�fXn�a�q��3�0`�3�k�e����*Lz�e���5�&uK��ƞ��Wj�>�k4)�d�M��S�<w��S�Nk�#l�@��%�
�O����6�ک"�ۢ�c�v^x��ټ�nTP��G;��خ��9+Ӹو.�
�������_�U
�:�����2�*��[�sg�u��7��������Q�5��\܄r�8���Y��j�zv�N��a���*���^�D)���9�ٽ[ws�[�)* �-��s!������#;�KH����F�^�("9X��\̆`�����]�`7������z�R>j�{�W���᪩]|���6�
n0C����������&+��MA�}i��)o�����.�P=�F�=�u�x�뢪[ȉ�"�A���%�`5��Ԫ؀�=�錦�0���4yQ޹`�D����l"\pW,��`8�.��c�������;��w�n����ĝ6EU�$:a���AǴ��ST.ӡ������H�ͪ{�!��6c��@%�;����Pg���9a�^�g�
ȭ��wO��'��Yuo�K#� s�^k��s�Ҧ�sS`[Po�T�q���c���<S7=��b�CS�4*��ӏv�?��F����댞		��ڰVu��{� �t�6�L��v{��0��J�:���:X�αت��@(B�(�8R6%O�sT=��Ś1yV0D6��v1�F�0�ʽ�P�!���*�R,9u�B(q��z��T�@���t���X����{K��]�G<U�5#]C�]b�V���0#Ʊl����x]��q~>�\w{Qurn�>P-�������gS2�t�F�/CǛ',����]����s����x{���AS����s���訏�����Q�BȜ�_ �����2$�=-Y�=y��KS�F�3P��ÿ�Ҷ��������𧸳ƥ3����MP�g{;&��݋�m3n,���f���H�|6��㔍����v
)�֬p,��o�j�F���L_$���I��EV}��&�?S2��u�*�E[���8�|�m����ɬ��ݨ�����^�JжZ�=6N����	�*x�5���>��b�v�����k���cv"j}*���f��n5����|�F$���N�Y���c�Zڍ�C��v���y��]�l�0(��y3�([W&���:�C�ܔ����-{x���y� ��>S���U��p楼ljz�1*�X�wiՏz�ΐ���G��ʞ@�9�y��-	����(vv@�Ӻ�.�U{E�1t-���b����ùO���6�2V����`,񒦏��,봂�g��z���=������5F���������i�d��w�:�R
n}��ğ:CI���l1��v���iցį�;���Y�w!��1<a�9�`i��WlX{���0�������d�8�P�~��yt��y�g��y}޻3۪��6��������3q�Vt����ݎh�Kub�6�ɷʝZ��
���s��=O"�ٺ���ri��1M��똛�ns��8�Ɨ!����:,��;��
�H[�z%���ꪪ�GB3j�WI8�{��լ��9����(��J��9f�m
��l9�����O%�I��R=O�a���)Y>�4ϙ+�W�;� �0.�yM���C���w�5�? ���A>LI� Aɨ��p�W�˔=۽����i��jt�Cl=aRu:�X,��O�v��ì+��Ì�I�!�a4�0�?�E�{����x�2Vc
���v�����	�C�|L��K#۩l���ee�c�e�3����6��C����A}E�C���"�Z�h��&Өu@��c�N3^0��,���+9�rM (���04�{dğ3�<ͤ��� I3 #�'�O�LA��9��G��ϼ��s�߼�4�̕����4��zɰ�8��|`^S�[�@x��arì9�Af�{�9�'�Cg��i:�N}C��>�*�㿽��C�@���{�& (����;�z~���<��6�g���N���&2�b��h1�VLM����Y+8�Sz��E�2Vq�ϰ�&Щ�4j��x��<a��Xu�皤����O̗��4�A�z�踨|7�Xc��W���#{�������~�?'Y�C��{d�Vb��>�p�,
�u�l�0�N�Xkka�Ì*���w`��g��mE�C^k��&$��q���$	�&���܌�y�p�+����!Ĝ��'O,�:�Y�
�5�Z ��J��:ũ�冓��8sn�\E�C/pE �G����)�=C~�i?3^!~ݛ#�"=�>�u_Ĉ�_����OW���s��~z~d�����ݓu�bO��̞O��|°�2�M� �:�X{��i`,�NY�:�����7��*�/,��$���������q�	 X��o�0q���z}���|z|�I�7��l�Y�)��H~��e8�g��b�Z�bVq:��`���ez͟fL>aY73�;�+%gR<��EVJ���~>��� A��\#s��u�~_	�]� �p< �YUϬ�>��P<6�]��%}d��g����+�{��m��&����8�f���2�ެ�+
,��g�I1
���w[jt��|>>O�=����ۮ܍��U�d�аb�L2��J�5۵R���ƻ�q&fĘ�W�Z훺`�K��J����ʭ�xM�y� lt�zvڢ�x�:F�Zxcg
�B�X�|^�U��8�{N��Y��k��"'-\�R�w#|�)�ݬ�\#���:U ¥��I!��b+>:���s��s���rw|]ͽ��u��+�!sR������Z5�ǘj��n��ڴ�R�v�U�Be9i����%-a�n��/�]7γ:�3��;�T�oSWBA�GrvG��j1��XI}(��؄Ah�YՖ�rnH����{3�*nw�b͇�)vA|��b�rJ�rƪ�
�o�*>	D&<��I��K����	�>���v��6���
�v���^]+�ݔ��R�9o{h�bx�IR��H�(iЈMggN_!ÖJ**{,��>d�]��������mpފ�[��������0�a@p����8J��:��71!LТ�Շ�I[|k�ȱ��H!�f4���*���#5Ç�Ζ�bU`en���ծMv�`X��o&R�.�\��{$ڽ���B >�xo�`��Y-ڕe˩�ԉ��A����Și��V�sb���Wv�����a��/���qS��F�;FU�4x��s��i��&eD�b�W�{�a�J��/)�z1�47N��3�%��\wx�f��h���
�B�h����h���&N�t~��Yuyt������b]q֑�bo)PP�奔B��U�C(�:�K�>�!Q����ڋ�Ʋ�ht4��no0��u#�lYmb��U���Q�{n�R�Z6��9��.�;���u�@�+�z�VS!�aF�9Z�6+��)V�oVD��}aW=u��(�ݡ��1C�a�и���B�#�v^�uc'ky;����	Ŷ�$�R�.�f(��8�.��B&���0̷\��*��ƴT�0ku��y���]��08	��5Q	a�X��Y��)r����6;s,��gr�f&3�d�7x�ty��|o�\�Jc��K3�do\����l&`��̮k;3r��(�t/Q�|6�#�6��C�=}�gJ� r|sC�'8�
��[T��Α�{B&敏��.���峖�𮴦���)�S�	���kU�hY;�`�M�����G�9G�;)6�7�p��
�]Y��N_e+�D�oq���f���.�}f^�M;;/�M��H��7+{��Ü�pq��X6��u�-M_gd��Z�oWt)X�t�ʚ�W'���` 	L���3I�kos!1��5{�/���݆����W�p˺��	�F9p��k�U	*v�)$��O�:w��Tn^��nN�G���&N�b�.��)�I���v}w��x��-MC𠺡+�����m'�.��B��b��6Wu>1<+�@j���e�
̌vf`�gk"��"��3�Y�,�jR�n�`t�����:��+��:���T6��P�Uf61QE+b�h�*���3(P`�h�U�(��UQc+F+Q���QDQ-�DU"���2əfZ*(�#l��QAjŌ[lX���G���-V�*Lh�KU�[Q�1��"j��Db����b8��%J�X�PR�TAZ����F$PUPEEE�X�e�,Y
�T���8�.eb�����r�.e2,B�֢�R�.X��+a��F(!m-�j9B��c2�`���� 5�Uq��iEb�nZ����PA�ZҸ�1s&1J�L�c2�"�U(���W�M!�"��]����kc�G�:�a\_,�����]l��ЬYu��7�,���GQ��6����d�O�r�]���U�:�O�w�{��z�>a�N9�t��_�<G)[>T�E���3&�S����~��hz������7��0��s7���rg̕��s�a�c&��`��-H.'�LN��.'�( �Y� ��M@�\n<�ߖ��@QH/'w�Bé�;C���M?�c1�m
��d���sL��1E6wX��w���oxz��z���'���M���a�<9�:�Y����G���$� O���\�_v���}ϟW�׾�!�(W�N�|`T=Vs��� ��Y'ud�QIϨc6�I�����hĂ��U���$?Z��=M�I��$�;�EĬ�� f���zO���[p�fF�'?~��s���@�T:}g�쬕���bEY�ONk&�*M�S�Xz�?����~�6�dӽP<�
�Y+���[�!�������<M��_Xd� EǄ���|�S�N�����N�4��n��l�+Ϭ�������!��!Xm������t��m ��^2iE���i�zɉ={�hq�9�C���C�*�Y�Kl����Ȉ�Ԧ��w�{6R�����ߦ�V�Y�LE�jAz}��
�3H.3~s$�t��,��N��X��x�&0��1��u��-�
�ղ~9�ڛfvɈƤ�>܏zH�g��/g ��2r1�y��
��ކ��&!�_�g�a�
�i��M�|�Y�O5��2�����5&��+�/,+�C��S\�>�Av{M�}�'�E�2Vi'IϽ�i���������~w�|���<�Xc�1!��7ܓ��q6��b(+<N'��&�u
��y{�~b���
�_w�Vy�+%g��EV�����J��(�a�1��i��H���U@�E^��Ϻ��請z17U[��V~d��K�}�I�d��w!��)���p���L�N!�R�|���� (�8��_����B���Xz�0�k,P6��?y�W��$ H$D�ϟ}��GÚ���W���q�q�t��T>I_�d�Sl=aP�'3�h�3���{܇���Y�?r��B�j�{���*c:�����7H/}�>M (������/��'����m��oʏv��5K�Y�6L=�T6�i��m'du���=��=�;|��,�� ��!��y�pHi���U���qïj��n�^���$�oP�Y��[΃p�Wk�5�<����U9}��j��z���v'����gW�9g\����o��?  ��7��y������>H9d�b�!�����yd�O��q��Y��O&�OP�:�z�o����6s�C��P+:���Xxʪ�t���d�E
�<;d��C��<kn~ם���y�������������R��ٮ�c'졤*.��g�1�7�s�H/�<-1Xq�`z��R����'�Rb(J�&��B���Fo&��I_|3��{�TǠ��}*�6�ӟvv�Q�����T�(��к�i��*M&�s������_����~d��Y�Lf2Wzy��<E �I6>��b)�`\��u�C�Ԟ����<�3� A>gAg^�U;$Ӻ�H�����i�'��k$붰��s���1d��z�������~a_����'�mRW����a�*���~��d���5E ��[�I�ω�<����>���W�oj��|ֿy��
�f���$?ZA|�~а�<@QC��]���c���4�]��;n�^����Y������c�&�I���?w'�=B���}R� 	>| �������3�?U�{��>���<a�S��gyCL<eEY8�����P��}܁��*9�t��i�'���6əC�+mR1'�'�;��Ci��ޡU��c'��z�x��M�ٟs�p��0a����s*�`A "�#�DO�:r�3O�RVf��i���YY.���M$QE�>�I�c%I�7���&�v����h�*m�o5`c>d��ܹ��J�Y���oz��s��\����g�b��`QG�H�	�sE���Xi?��Rl��c4����:�:�
��=��k���Y� ua�>|d���u�a���&o��OP��������~��{��}}���������T:���u���3XVz§��]�7��OCLZ�����Lg�*C�`~k�Xu1E>���a����q��?��A>��x}�=��K_����;'���vLgN�!�RT+3�<�Ci>B���v�|}@�0�v��]S�
��|Ԙ��TU��9��z�P�Y�����0+���ayH~����'�dd%Og.����������?P"���M�~�a߂��u	6���~ܥ��1Փ|d3�<�9fX��� .�S��Hu6�P/��U��f�B]�bf���^+�ʊWn�sf��,;��:l���]N�i��,ie$���UHx*��k�6�պ�*���[����Uy_�$x�G�}�dy� bA}Ny�mYS�ý��TJ���z^��A@�n^kSi�I�+?wx3o�)+'w�Cl��yea��{г��"��N2c>d��p���Ϸ��y���~�3�ܟ��>d�甝�aS�M~�}� ��J�;̓����[�J�É��|sY4���a�h~���!姙�iAf����x�
���f�5�1��w\�]���f��}�}������%E����'>I�|�������l�z����K��z�~�q�����	�h����a��P	��>�r����W���욜���C��Gg"��ću�h���LM�̋�H/�y��f�gTYd���v��7��!Y����O��7/p+��a�<����~a̦�+����%�	>I�̄�x���;7ۣ�5��Y����{�}`W�{�5�V�!ܧ�P1�d̡�Y�4�Y�7>�]���1!��P*����@�(JΧy�Ci�����LI�"En ��B�r�'�!7gk_����J����d��e��s04βT�~�Y�%g+�k̅CI�&�x�'��m��1���R>I�n?2u1 ����&�Xu1<����U>�]7�	�n�To�C����_W}̜AeH,��q�1RV�Ρ�m��l��l8 |��gr�Ǭ��/쒰�q�f��~�x�HT1��9z��0�g�9�0�g��~߯�+߾���7��t���M哧,�|�QC�٬�$�
�3�:��!����d4�Ld��ri �OMXz�H.�5C�6��a���d�݆yJ�RT+���~�ھk��|�۞k��O̞$���CO��a��hc��S��N�2�Va_����J���4��^$��ɤ:�.��w;� ��N�?oY����M��L�� �����2����b��~���[��y{< Ua�H}���Z%c���
%N<dĞ'}��6��J��d�;�o��4�d�4}�hu���<�f�m
�d�ǯ�Y�(�Y��8��S����g:��&��G&��cv�Ao]v�Z��ظ�wSM��x8�\�z�=3���%dt@����.�x*(ű�$e�k�����к�0��O���&0fS����ړ���+��)��5��P���5�;L�,�ݜ�;�L��0�4��-�Ppٷ�� ڪ���x��M7Q2�W�Z�~C�5f�2_iRK?2Wl8��y�|`\���0�<Hj�6Zn��T?[�gX�Y�6�08ְ�]��0�wT���2cB'���������c��zH'�Hd�=5�M$�
�����ӟX��<9��$�{�*~���M��7hx~�"�̕8��Lt�_��:Π��զ�@^"é�5>�H/Q|&��dS��T^w�*Bgr�|,�H��y'�.�Vt�'��i������(��7{��Y1'�W�o�ACn���_�c��u�����|�Xc+���`,񒦏��(i� [��7Ǎ��K���sq�9�3q�~'ⰾY;�n�4ɣ�ޤ����s�x���{���r��*����y����_3�x���E��M3l1'�sA�O̮ذ�ۧ�>��}1���B��uN��Wd��i����b(��%g�79f�m
�d���a�=����Y�x}̆�2\�d�c>d�0�����/��7y���<H{l;���YP_�������\j�������`��^�Èi��jk�8��z¤ߴ�:���O]�(��
�s�q�i>B��Rc�������C�1=Ձ���m�d��5i�hϙ*���_ir�؍^�_*�������<	D�;��OY�ć��w��,4����i��SG�q6ïP���I�b����d����{�I��;�3��1'��s��N�^�@������׍}z����o�|$�I�����:�Xx�^�Vβl�8��|`^S���m����~��Ԃ��?'5d�QHn٤�q'}���}dϬ
�:��$=�o���Z���a����~���'�E�	 A?w�'��|�a�y���6Ɍ�X���h1�VLM���쬕�d��wH��+8�3�%I�*cj��x��<a�è|�5H)���&��/iX>����;�N�/�)������i����i�o �`]���q8��[=��O5g�,�;�b,
�u�zfI�+�o�r��8¡�y��;�ǌ���
,*ʾ�1'�GΫ�W�E������F�m��s՗t��J�=�J���(���w��4���M�~��Rիp�Y���i._��y�%�����y ʸ�a��~w:�c�Ϛ���i&�R=��-wKه���U�ݴ�:�"]�۸���V �&��Gq����]��%�����q�$���>@Dy�O��yf��%gXT�k��Ag��6s0:���9��u����Û�a��3�H�����PSl<z�$P]$��;�����}{��羟}��o���[&2���d����
ϼ�bO_-���W��O'�l>aXxÙO7�L�%a��2i`,���M��Y�[�C�G�\���x�#����r��"2.�,�2f�;����&ڊf����?8���1��d�Y�|����'�)��:��b���Y��}�X(c&�^��I�>aY?ܝݕ���</3IQed�����e��~�Ͻ�Ys>��~�~d�O��:�믩
�i�[ɴ����R��S�J�d��g��1��Wך�!R���MnÉ�i!��7�8����ZγGف�zH|pŰc_NW����jLO�z>Fz�0�
��I�9H)Ǐ�>։���}N�bOY淛C������x�h~I��C�����J�a��a�c&�u��� ���0��� ${�ʖ:UF=������w> �]�á�aPR�﹡a�x�Chbs�M?�c1�����['���i��& (���P�;�ɈkT�$��x���ާ�=aXc#�i����o9��,�ʾCu|"'�ݞ3�U�������}d��i�P갻��!uH,��z���i���ϰ4�c�z�O�H/�]���.!�ֆ�(z�f'��d� ��d_m�u#���{�r�ߗ�I�
Ɍ��{LI��T7�:����Y��i"�,�&���d�6�M����a��̆�������³�J�%���c=d���͢�$x����3z>�n:�6y�_}���l���9�C��j��~�$�,
�q���Ci>B�y�ZN��=Cg�HF�
h���&�Xo��i�zɉ={�4�_���y��$�T�����G�7_d��hȝ��6j����+>d��:^��~���0��7�E� �;́��Aq��'��f���mE��ۏa��z�?�X����6s3�*Cvɳ�d���& .{�y�����3:�
�-֖�
�r�c�&�ψ^	���[ke��U�"�m�N��6��c��;Q[8_f���9�ܠ�q�00���C�ն�β�^��Ԭ�hm��u�u��	�#�SbjڵӀu�CNa��{M5�m�=�&M9�_0��z�tv��ǐ����V)ئ��e����35���9&���(�C���<=��=�x6�ֲ�ߞ~�~I�
�|�b��I�����̆�q�a�6�Z|�Y�Of��C�TU��}�5&��+�<�̅x��b�S�k���H.���>ݓ����ͤ�8}��k�n\�<�{����<·�����Xz�H~�\�L�,�����@�Y�8���$��i��?1IXq�O.���YY+8�kj$QE����L�%I�����π��歸��귏�Vt�f�}�O�?'̟�5I��g+�K�pĂϙ+���C��R�<�p��é�i'��yHe�J�×H
,54wY�6��T3��k�c��Ā0�<+>_��{[�d]n���|o�7٦J���g�1�=d���*��;d��m��*��xs��8�Y�{��{i�3��06��P4�z������`sT���@DY 	�6�����c̩��/�#�JX!�y�
<A>D�:}�9�A�d�bl��4�¤<�<g�ǩ�Ld���g7d��I�'P������7��n�@���+����|��&��P����߿w�*�;3y�+����>I��@�<>���3<�&�����4�c�oT��6�_Ry-1Xq�`z��R����'ǔ��ҳ��;��8�d�3y4�P+�e</����k��}���s��?vM�Yed��s�IR(�ϓe�CL�%I����z��Ǭ
���+'�M<՞�d�c%q����Ҥz�e��é���5a��(���L������m�C�B���ka����|G����(ӕFb�T@��Ɓ��z�#��+��a�V+6*c3�Y�{�Ps�z���Ahg,u*��R#:Pw��29�D��qA�4&0��R,��Xb���^��<I�k�o�q����jÛ>�:	@�9�>\�7#ɓ��������7]f��+�3�t�����K��Y���6-�PY���/n�gM�n� <�\H��͊��]J*�-��JI�ë�}oR��P��{9�a��س�g�k�(�ZI���x70G��yL���W�UW��'�Ú¥Ց������ۖ��l���J�D.��.VgL�'F�������oktj�0q��D
U:m\ᜈ.��>����qJ傏\b��}���@�_��wÊjwC�����O��`��C�:T�8@�_Y���l ����yE��������&�&��W\~��ڨ��)�D����>�S�\�Ɓ@��C�x�V�n:x�SW;ї���v��s�F�7�3Au�5Ў:��l:U� "@�L�HX)1�o�w3�&߰6%��O�K!�^��3�)�1�:�G�%���`�ޱlA�(αv��93�x��Wc���X�J8�y)ӧ�:ovp�T�Q� j:QI;�*Qq�r�`��.q5��%.tl�X����!��qK���e�u�U�$�x�l��e�w�����G'Oj��mGyEDH��W9}p�q7���E4�چ�+�}�(�c�������Q��>Vk�Rak�1���_�s�Wl끚���BK���Mv�yK�ڥ��׸���Y�bk��?eY��7���vQ���u�V�4Tk^�	�
�Xx	����>�l�3���=CݽX��^�͆�Ro{\�4�f��ws��7S�9�3�D�۳3_F�Q��{%J��[8��]!g�{�����ڒs9;y�qM֟��@��:�h�	TR<�ۋ��,��˓�N8��,��;qk�����rU�1ȧ�l��808�6+�(b\��/KYGd��9[$��Or�[닭��T\,8O�Y�%���;�P�9&����a�e_D�f�7b�eOW��R^���(=����7Bȱyv�}S�Xٲ�����ϙhę�x�w&�k���WڝEU�Vn��=wM�(ہB�pŷRt�@��e����wB���;�m����"�(�fxR��c�o��~̞
�f�����X�vUK>�0WW�V�n��p�!K����idQ}M��3��=��Z�Wk�@�W�y����� r,�ĺ�	&"'��q֥�(��U�ݏ��x�
K~�c���s�T|نW�9١�i��ܐ��Ә�X�bЫɻ1�ܬ��-�&7uhc>ث'�ρ�b�v��U��}q]X���ڷ�8!*�M�*F��+�mO����W���qJ�B�v���8b��A������X�]��L��[�
����{��uᐮ��K��{�@��ɍ��Ӷp���f�E`���� ���=���_h. ��Pf3��4�uy\({��(�N|�
r�s�f�{�[�s�3�^)��^@���\#-e��������بV�c�����3�#%�&/�����tZ���Ҹk�5����l���h�ޫ=0�2�2�(���T#��W]XV5b�b�Ez�{M��]n�q�K�� �w�M�e�l�'S9K�,_�
*������s���mpx}���[��͵W�+/�^(�l`B�N��GK�F���q����;�:x7 �8�(���F/D�[�w�����ee��R����h�T.��y����NH�J!P�����@Q~�>B�26�²o�=�kM<��v��у>���pӍ�a�v:�ډp���]��5~�gAN�Gb]ۜ.5����hD���+~���u2"=o+	p���)�p�/�q�n�hؙG�:�G:�sD̡y �=�+<ki)d��`bcƁ��i��-u
��v.��k��ŏ���3�Y��.�Q��Tu?��,�ț��7T�v�^{%�x��<����׬�=�}�1tnOb�U5}B#џ@�VT[S��A��\��Ps��0
��*�'3b�P��қ>�m]s
��T��q�ݝؕa;�	4p�6���-�c�wt�)�1�ݯF�	-"fV���A�W1W����%�V���6�!$���t��B��;ʈ�/�w)�ȩěx����u<Tv���{G�+���[]�*P������xRk�/�lw?z`����,�dH7Jd���P�X)�=D�u؍��yu$��O����0�75�i�:����W/�0��ǃN��/�X��X2�V{s�_������H�v�����Of<4�H%�9�K�����y8Y��*p\�qe\���I^�0�`�86,�bUz�	EH���
�:�7[�
���p�zH���o	�G2:n��1�^�F=���,h���S��)�QF��t
]\B�ȻX�\��7U�w"��L!la��TpU �V�n�\�(�ڒTOP��W��K���g�ֳ�+j0�;��q�(�9s����[����
�^�A�jV��Qj�cd8�vR���p�m��%ǭCQ��ҝN�Q˥�:GX�@��3F�����͸%m��&6�=!n�xC�����O �c"2a�86�
��,��ei��S/ �6@t��y�_f��X�;s��NMp֟y-Su5�YvP��R"�:�m�TV��2�QU�e<5u����/��yOVf�o��.d�kXi|�.����ܸ�n�79���t���]v2�lV����#n��� on-�殫��Zs�kD�o���8H)�=yqԢ�wVed��5�VḦn|���}op,w:�vs$��3�R���M��_PWDJ�V�˭��pĪj�t��ZmNf���pj�s����*� iІ�q�s�5HdQ�gk�m��/r�2��@�T�����J��cO�}�+7��Ō3�ڛ՛I�!}Eg`��esn�gw.�s%Ԋ��M��0us����4Z\L-���Z82�)y՜c�S����쨞s�I��8[��2S�c��4\ږV᭥v\�uG}��'氆��+�ع11���UʾYǨk���D<��Gc%VRS�s��[}���+]�z�r�#�F.�@�Ϙc�:����T� ��0��2��ܻ�Wr�O:Y7S�Wm�]��4�S�eacr�U}y�N�kZ��8Iv���\�������+`>�_+���Cn`��D`�2��9�a��z�;t���?��9���{[���i|��T/�Ռ�2��N�n�\xV�В�;��6m;�o�U����
�ռ9���C�g���:�֞���V����u�݀�^$C����@:�PYG��%�IXF�|]�=]'%oL�j� �m�t�n�k�t����ҝ�
�H6���@"� ���ԗ;T� ��J�w�4�5�d��Kז��f�[�W����l�<�����;_
X5�[��X����VC5d!���!��w�7Y�DV[��u;�;���ɻݼ�,K/'��M�9{vl�Z����.�%L,MX��И����ɓ%����﹡Í"/!�8�<�]u!٫o�_f�R�0��N�v��O����*��<������ά4�V9�Z�ݵ-�!�g��ѪW�����l^	��-�������5�y7�
��hz��Y�\铲>��n�s��u�{D��Ew+�gWU��V5k����Wy��>
�T�'	ɨ�T0������I�Lk'~��A��`n�xw"����Q�G!���#A��H��AKC2\��L�F���j�1`}�t/�ݸhk���tH&�|�n�_j���U����D�stд%q{X���a*�B�f�7��ȶ�VR�]�,#��7,]����\�sᏱΥ϶[�G�;WʧFr�^��U�D����ozRF�xR\%��`�'Jռ:3Ac�ͼJ�̃��SHJm�.������7��k�y���f�����psƉ�kt8^�.r������G ]f�QT8��}��_aT�l��X`θ���j�;��s:�nZ�O�J�>�W���['-����@�Ed0/�lQY`�/���%״����t�B���|�,�+��
�[�U��3n!�\e�\b��\��S�������P�*\��(�f$�X�e�F-���Ī
T,J�J㉌�[�9nY�X6�"����c3+j�X�Z���ԭ�*T���Vª,+kF5P�m�R�#��Vڂ*��ثR�V5*J,�b�25FX�e�LaQU��ʲ�Db��-��K**[T�(5
�jZ�%#KU�����**�e�A%�Z�TE�������j6�f&ch��EF2��P�F�Qb�k����ڂ�lkmJ")YV"��B��ZUU-�+T��YimB�e-)A%@�(Z�e1Fږª Q��"6�h0�����F**EV����� #� �@c��y�ErO;���ݡ:0��R��sIǵ�(������8�����jQ�S����T[�{f�g b��<�  �Y-\�TJ����7���+����̣5�u�竌��+1UZ�`�𬀮��k..��[s���n�u����Fb�i�(3ƙJ��W��絯A__<	��A�*o)qIq�ͪDp"�aA-�Eq�u���^�W�T����!�c�e6�B�SlJ���T]�!����tIa[�j�(>Z@��D��?xߒh������V]�h{������O��l>	�O�)��r���x�����o"�#�^r7����J�g';wQ�����Ǭ�z�	讨+$s���P��.��^�J8�=Q�Q�thܮ|�K�0��oj���w���4F*�s��Ɍ4Pq��AG6�FH�����`�^ThL>����q��} ���J�q�Lq�fp�4�ϭG.Y�T��ਥbt��@�P�hm�
ϫ��os��YaH܊�A��uꢦ�����J����wys��3s#D�o��i���]R���J�7��F�3�yL�X�6JB}X���̺1�3+	$ю���[��͓���J�k�܏���:���\�{b��Y<fm��v��v�ފm��t���>�(��yf5������o6+Xi�S ��9���W^sp��+v�Ψ�]֣��f�e��Y_����{s�8�$j�_:LM�få!��q�<tgui�R��8����Ge�ż�IeaH�.T��'�X��aмR��qK���y���[�L��C1]�|f��ؒǝ*��B(i�Ҝ�j6�>h�U����eY�]fS������v�s+;ę1O����h/�wB�ۖ}9J4&��¿u�(O+E���0j����T��[�J�I�8�ޕ����N�8�U�x�"�X�2�Ý቞䝩���.��3T�g�V�,76]��6hti�Ď5��7��<�΂�<i:V�ZDݽ�յ��"u�A�5Oҏ��[ʓX���%C�9&��8����`�sv-�u�e�f=<tո�5@�u�^���.�l�8��Y�2�8��(�7�`�2�I<�n�Ws���3��Č�q�Jۥ��
bq�M�u;��"}���5X��{{>[zr�N�=If=!t��E�!o����4����f���\�ʨ�{�P��?Z����Qo��+rue�)�V؈:�+*V�&�<t#� �,<��إ4p�-�o��~|�e��n�y|�o��z�M��wՆ��C;һP]���Ix��7G�Yx�ķ�bn��*ͺɕ�pΙ�sQ�|�g�� �{�Ɉɾᢣ��:�4�I�n�L�cB�	\�0�l����1�}��3�:����ƟYc��8��E*�9���N����F:��1�ϛ��Ae���ݹ�Z���A����4t�(��(���9[4z�����Kdm�O����h8e
��a�bȬZ�k��ɝ��ݬ�95(yr��]́�Z�>�c�̤���)�`��0JAT\����/;�ӵ͙����y`�3E��.��bc1O����(R�ү���z.O��s��s�V�^#�%y���\C�3�
�J7~.@E��+��Ջ�(�2���Q���ȭ����"V�/��ty��1ʝAb�AEVF�(ߦ���'�ܹu�~�x�o�� �l��R�<]F�v��rۮ<�� ہe�0�$��x	��DTԹSu�2�[Ne���^.p�z6y��O(ܹ��9#J,��8BҡEß!�k:)�c���薇d�ut?T���0hr�H:U�˽����NY� ur�z��i��<�f��^�ge�C��#.s=���+*U�6�8��(0�͌�0��m�RK�*޺E���;��Q����%^�V����w.rn��-��̽�V��̢�arn�����l�&����,��[�/��,U�څ)ʸ��	wqŹ4ꗗ��ժ~�����y�=K�ZMGe꯼ ����� �^�<t���Q�a�{  ]��b��`�)�%���*yfw�l���n��,Y�% ���(,^i7����X���1S�>.���2��/����Y���~۾�I���`����}`���4}7�4x0����p��\b�t�����0��hR<'��p3���Ԟ����3��ã. ��r~|�����x�P �3�nb��.L/<�t�W D�`��X9��
�"���u��۟&��s�)�Z��fs�M���@�
�<���#[�r���4h֭�6:{-M��OaĮ}�T��s�w�J��y��t:��t�aп�879����J}�MV�j�2�	��{c��X�LZ��h(ܠk��+���R�3˄��D	�^�d!��b�p��7{,D�U��<����(��S��8�F�j��9F��cGE�
�^\���v��t�YĬ�K����2�:l�V�^�A�[l
N�E�T�Vߡ�7e�l؀�O]P����0\2�e�]~Ԕ�Z뫸�+}ļ����*��>�%����3����)r�$u��@q�uh�cݩ���Bɑͷn�҃�ud�Z�9��l+J��5$�FAB�o7����8�� ��mf���]0��!�F��j�QEr8��u��[����
:zM�Y����7q��y��'�㰝H�E�=�k��ӥ;�N�]���q=�0nY�#.A�E��;vޡ2%zc��B8����F���H�^�c�"�~.�YZh,n�kA�������a�}��ht�����)q�B�n�B]/k���W7%��DIV�s3Uu���Gy\�0x��>�Ñ�<���K�{��3����0bFK#k�5ǵ���B�w^ZO;u�+��\���D�AE��C�1�i��:�g�g�ɧ������e3���һ6��8��a�%�6B�&h���lۛD�6yhѻ۸�*v2vcȊj/Y�������d��Rҽ1��$��n�tI�{����`ϗ1M����,��A:ߺ�P�A�k�[��ۭv]u�����E9����VE��^��UK��B���.�w��L��[L�K2L�K3�X= ���@��X'������+�~]B�.Ǚ�b������qS.!{u����Wo����J��r�:v�|�<��a�ۚ�1��I[&�\��ܺ�tpM6�!�}���<���e��]�ӹV9
���3�t��Nwij\�#&�\��u
+z+�V��Lb�X�F�u�u]����8uZ�91�n�쀒�� {��C;�A�Vw������mA��n��,(��
|�Ҡ��Z6{N�Ӵ!N��K���[B�_��f�ڨ烥)�E���v �G�)N���up��ct�70�t�8�aE8�wO��Β���X�}8wY�N����]`+�$�L��9�ɻ�y��3�� WN��݇���t=�XF����m�<Q��x�,.��P��-��o0�}�c�v�i��W}�,r�Z}0���n(���;UǊ,�ѝէ�^fa�U4��������^����8S7�S�`_��X��[���A�)�{��v��f���ws��C��;qO�VtI�N���E ��W^oh_|�-f������X�����#���L�M�e��W��(g��0��g��*�>ugh��@uoJږ��7�٭�����ɹ0Q�)��F�wN���`�ӘJq��ϕO,T�o�E��3�#1���A@9��Sg�f�xti�Ď%�<v���S��]F�Ƒ�J�}:XV�Ә�7�2�uj�o� ��nz_:x��8��)҉n���{N���w���v�=:�[S0�M�P�!\�1�6(�Nc��	�0�)F#�����,\�b�y�QA���qt=ó��Y�1�I���:��ڹ����S+k� ắ�S�'r���=1fw�'��_]I�r�;<b�;rM#����e�����K2RՏ*���P�k��=�j
�/Ђ�~V�x��p�⃙�]��Q���%ж֩��V���p(-9�S8�m�oFR�"�����I�h�D�2���)vѳ|yb�H��Þ�e�`z��:� ��7��(,ǐӒ���࿛ׁ	f�W:C(����3Ǜ��PɩC/�N����H�O X-��V��X�^� �9l*ڜ���Ź�NJ�{���Ū7�=�{�q�6X*����O����Fy@�"�W�M����@go!��M�^6&WbQpý�4,b�0�b���i����f�[�QUvu��� �����D�Zoq-
02��.���WX�r,�4-*�k1��w�y��WI�=�N�[�'�k�+"Rt�7���+�Y��-P�1x��M�7i@G�N�U�	1#
��n�mw������P�*sW��C���B�tz�u~�R_>N=[�B��A��Is:6N!�tU�w[�CF��dQ�Җ%��u=�;@l5��	�A�WXTZVj�aN�͓Γ[t:���;���ӬR���NW��$��R�;�}��/��.X�@�O`��Ȥ��m��p�>l�KY� U�}�%H����_����)N����}�y�L�N�gB��8D:��kM{��_��s
\�c��
<���G��>���J�����E�{��B�*M�9IH��<Y�Q�]����YPy�@��Q5��=�QS<��t`�ã==^.ti:��t��sŚ����0B�j��iP��V`��í�}��H��^�zx*�V�M[��*�3�y~��j/�嚋�:4Z��7rq��D����0_�OJr���5h��e��T�v�CTG8�d�bN���R�)���6'.����`d����c��~�����٫�AO�Ǌ�,xû�Dm�'Gy��C��S1�*.�#��"}��u������.W�X�s�׮�?j�#��X~1_��=������d�齉z� >�2r�rv<�e�h�qqI��S\RƝI({�`��o�ٮƮ޷f�*�u:��=�P���BVO�:�2�QWQC���rj�0taS�6F�Lk��+C���*�Ur���;ع5,$.O��<k����a��Y�nͧJ���"��6<3jt�B��n����=Ʀ����5P�idM�^d~Tѓ}�߂��*�S�	Mh�^gP���	�zyo_R}��n���`��y������� �[��A��njo���N�D�ϲ������y܋�Ծ<
5���]G�Z�jC*��C"x֩.7����J�x����g�>u~���;��9����{g��k���l9�܈�t���l ������{$8��.�z�I�؈�x;�ڝ������������y1U+˜���oG���'*���|Y����"�)B�#���lJt�,*�N+.��.xDmI(���^9�˛|��������qB(ׇ9hg:����a�/���[fT1YF�:qj�s]9��,.����`��*=N9B�ӥ;�N��.�w��	{d`=�hm��O b��]�]�U�Y�ܺ^�W�L��seY/�x0��]�*�`늰xyZ�,u{,QǏbw��Ԙ�qQgvΔh�/!��\j8�t\�_�"�r�ۃ��o����O�h�����ſybͼ�e1Q���]���	�r��gj{[�[/v�XŞ�e�[.᾽����D�0b^͇�e�D�|Y`�].���@>��D�Q��f����d��LNtn�T�m0y1ŗ�+id&9B.yo^�Ã����< $>EF�������v33A����d�I5�y�������N�H�s����!��8�����ϙgU��pU�س����U��W��A�ػ��џ{������*.-�P����g�7L�������<4ר���Ru�x!�̥�+qZJ������F��j�;*�`8}�����j���%��Ny1-Ň3SN��p��)��SG���S�s��:�Tīa����[w��k��&��@�SLj�#��-򗇱��x7���y�b��r����@�S��ȋ�+|2'��y��p���)�.Wk�H�̻���:5V��Wb��=�`�P�:玕��v8�gkÝ��C����c#�j8tRj�ߓ���w\v���סV�e��qɦMa�Q���܈�SX�7�B�W��`7,颁Yg�<;���=�Y�U��{�b��Y����0uEXVe��|����ʂ�"(�~ʝ���E��W�~#n����u�k���J�蓹8��
�'J/��W�t�X+&��1aR0��0ly�UǊ�����kU�e���w8&�ro}I�F#��8��l�O��l��V�B�nc
}�^� x�3+�ި�Db��6KY��i��9�g��YG�����R�7[����`N�{���� ��]&%X�}0˭�r���@ڂ�e�O���zg3V���q��=�Z{�, �YL�.�)�츏Cջ;��M�/Y� �O����W l"9�m��'��׊���4�t	��n��;����^�;n(�q��{j)B�d���GUpB���8��4L�K��hqק_uX�(�6��I>���Ԝ�=G�e
4<�jqǦI�b@j�w*�ŏ���v�i�o�7y�kՃ�e�yq,���mZҁ�U]	U���\睖��c+L�n�-����tE�(�	q�؆���T��`vLF1,�+��֍�s��j�3��V�Wdo�ӕ�WSrj���*eXw2l���d�X��k�O�Ȓ�H4x*�9���@ѭR�pe�I!CͥX�n�Tܨ��
�j��p���r�v��Z�t�� a������ǔ���_bڗ�1���<˥��e�03�iJ�WV�lN�mO�&�A���A�D�gCM��=3�kTRQ�*�����|{�g7¡���n�Ǜ@]�;�ZȷC������X��35҇)��m˷��ʼ�:6����5���Ũ�k�\��-�l74M���{':Z�	�.����W.ȡ�tV쳟|��s��o19�ԽM��{TF����PݸS�]����1:e�aLP��٨r߷5q`;"r7�/$�&�\����tmV�μ�+�cymc�*����0������."$k��
�#��*�Ò��۬y��<�w:P���
t�ɶ�2�+/k47hʁB�7�6Jo1N�d݊Ǜ��m.���W�\��z�kx��i�ca�����T1�[�-
��.�3�CyK��PE�Z��>U9��黙x5�B���E���*�����w��C<6R>�#�U-�U8�B�'�7D	��n�N���n �kylm�AU}�wG7*�d\�9l,l�w7��W�i�v�%\�!����Ƕ�7F(�˩�����4�wvj����Zx���n%G�)�kE^f��UKӄT�I�Y[�I&n�򊎦C@ ���Ǌ# �P�ѫ�hX.ù��n������L�7P�:��s��(�բ��%>��y���NC���ʔ�V�����1%���P�sTlğ"{730#��k����=|�hՒ���^��d�MW��e�5�*fø9Q�O�˙4S`ñY�i
�:�Mp�i&�	ַ2֞-�GuwoG.X���˛�����3�T4m=ʕ�t��N�"j��Γl �Z��9r�K{�Ay܌��u��l�ѧ���)fR���&mw�B['H~��������XD�����{;\�5w��P�x���T(X��ZKliIQDVҔm�X0X(��m��m5a�5RVڥ-��-Kl����cX�0֔F�E�FJ��Km�,�-QQ�Z�mjV��kU�ڴ�m��QVVV�Kh�
�Z�Q
��m�hUI��ĭE-KE�V��
(Q*����*�e�b�kXT�l,�-������X*�F�J���EPPJ�l+-�j4�V0s0ȅ��AQ*�-�ĳ��)J,Z[*�в�Z��KKhҖ�em�j$kF6�"V�l��hƋe+Z��ڍmj�ŕ���m�,���,�؊�(�����2�����&ƘƆؘ��K��i�Ʋ�c��ʊV�b�V�s2cV�kT����ֶڨ����5�m�
�XTdFZ�*B�(�R�i�-�V�V֥�ȣR��(��	�&�I���}��1���.s�z+����޼���0B3	t8b:�g1��3���v�f���"p��p��uA��g22���������%������˽��8���Y
E�.���E�9:S��mGR���ޯ]��Q���ᑻY�c��k�D+�����˔��܏�+��x�5�vګ��	Ts��ڼh9�tQ�Q��ui];һe���8�A(L����^B�{��bVC��oV$Pbua"�����^�Q��[`�0�ӂ��EV�؞<���n|B�n�2yu;�켅7����]�(�ƛ3�0���8��8��wx�(n	�3�q�a�W���W�C!N�������Vf\��->���YV}fRj
�*�!U���ϱA�x�t���w*�K���ژ.���g����)���:�M��� �i+1��%vp�]�3RuE]��|�Wvi�XW:MuE�+�1\�A�y3Z�q����t޼K5b����D��U��b�/kmc������5��4�T���M<��<�t'#M�V��(떄��mF�>����n���|�������T"������s���"B�2����0O�X��%�)v�O��dzh�ԕ���e<O��d�j���A���~�RN{��*��o}n�\�u�B��Ks+��7�1�䠵lKsOv$�S�x4��w�dI�uO]���l]:�̈́�����������^w}���y��P:��ĸ:��u��{�D���7�(񑕐4�}��1S}����di���Nʺ�nT�0ZU�<�{yyW����_�־�������Vm�&=�^ؚN����x�p��UE��ԍ��e�n8Ҁ��]�^��,��wru\����Ҝ����[108����n�.@T!ʺ��b�5b�$t��FFC�Z2��"�Q���U�Zk�[uNb§PX$���D�~�>4n��ڌ��ŧ�
�[ft#,9��XΞ,بӭO��Ӿ:�`:����=Fi�Հ	�ӳ�[:�<��R �N�H�r6S���6��<'$i�}B��~4E�'��r{�1���M����BC�>B�Fո�T�fU�"�f�g'��z��~^vf=�-�r<��0�n�3WԌ�R�Z������u�	k+�sj�85�γsmm2Ei�o�s�[x2��tO���{��t�?y|���$���7Pǣ��/%��kfY$U�.�m�N���j<>�2$X��QӲἊ'֩6xT���h��U�T���YCZ�x�_7}�2�jΧtd��Ӆ��H�i�8�N���\�8tfE&P���,ָɷ|� ])Z��u������c5!�x'[2���o �8��"��
UGT��Sv����5�	>37�v����@e��2;��0hS���OX~	�2E�Xqpܙ*�Wn$.�o�t]U1����DB����v7G%��8���j%з[6������^��4�S���̄z�{\�f���:gM��$l�]�,�g�rB�v�J�\X�ρ
�(���w�v����P�Y�����u��V9�Zk[�w��L�Y8VUQ�����}I+࠰�g,���Θ,�S�tu�,�5��U�P�9��C���q����cX9b���y������D+���񁧨��6�`
�B�m��VI����
�-jm�X軆k�2X]<�Z����FGg��6:(�Z���Vn�l�!FPY�ڸ�W�x�n_@�]\E�R�z�u��6���0	���fÎ�(�`s �ItDr*9d��H��3v >�k�r�N(E�q����a��3~
���ˊuY�].�Mr��,9�L؜f��������Tw��)�֝Q~](׵�{�kٻ���jU��y{�Cߛ�����Y��;�ة��`k�va��m�������|�4� �&�Y	m
7�Q��^�J����d��v�G��o���k�j��G>�G�:m�f��hӒ�*#M�\Eu���_���-���Ic7l@(��)T���S��O/�dEL#F��)Ō��d,�}#"B��vM���]��۴�:h��RU �%�,i[�+F��_�%�Uc�k�C
�f��k}-7\%���G2(�8�2���`��[�Ȁ�
��K�o�a�Z\��=c3v6����12�zh��Ly@�9�v͗u�,�Q��Fb�u ��%+����n��Wp���K����G�ȉ�Xd�;�m��󢸊�z�@b#�0'�w->��Ӎw7&e_/#��Y�6�)W�b�(:�������P3��My1-���43"�Oj������H����u|�z(���;���"�	������OO��7�eȁ\ߔ��u ޱ~������� i�F�jVو�s�2 ���9`��\ 8����{�sN�dv�W��6C1Q��鞰�=`�:x��D)�۝0��wmvbG��-����c��R�&�V�:i��;P�1]�UiV\���� "
�r�k%V�*N��uw_I�Is��C]��o�39't���\�ĵٞA�;&��^�
1���d��}��Ip�̝�:)����܈&z�`�������}!9���7-uʾ}҆��=��c�/�^�z��������\����N���p���:hdPخ���U��
���NV��m��o���z^w�D����wBk猉Uj�*������~�/R��|��6�3��ﮥ�����JO����K�{l��W�͈HW�l�+}N����h�6G(�+��͗/��/°�:\�4���B�dFQ�S�
��ޤe�zT����"(aмR� L�^)�0��w+3a�oW�PF"��	g���Ua�L�e����TO�>3/"0�����s�8jT5�ȿ
�e�]^��n�8� �%P�ۉg�3d�����smwj̄�^g8�O��YR�0%;�c�"�g\�F�WN��%���܂�P�GAX�0ٜ����+y�J��V1R�@�%��,�%�;U�=f�!И�Ķ'��&%��輝���ī��\����B���(�W��ۗ��R���#=�8ܾ�PQ���y�d�#,��`ζ�]��zz'!ى�+��� ������bc�vm(��pIc/%<��f2�k�]G�`R��d�{!]H��==[���:V-���bWBu-!GO�W'����)�E�λ	�5$�[Ϸ�:��3�U뵜��z�{V͎�1]N<59%��^���(+Od���v�ƌ{{0oV�:�-� ��W*�E�5�2�C��H�[��>�X}h�6x�m��т#LN5*�v�;�.�E��w}�$�!����d�*�i���s��E`���M����밂�9ѽ�ϔ�ky*��tܪ�� �j$]=�$�!�:<�����n���0g����rr4��5(�˂�6��;o'��n���-]���C�n.�΋�k��ܝ1���T�(.{s܍�_w��Ԗۿ~'J,�w(9��ϱ.����ؘ��\l߁Kdk�K�1n�<�ol0�;7p�aƜس�q���L:��%H� д�	�c�49��%>g3�>7�e��WWSr�pz���j��u�� ��4�S;b2%�&0(�J��S�ޞCn�}w��&%l�@��N��|�vF��.b�R����p��6T��1��<&�]c�CGk�ǂ�Y��{C�tȳ*G(��ӎG���1aS�,Q[��J4�����a�tE��*x��a�!�13j��B�"�gK6F�w�^�9i�Օ כ�K�Bq��I��*V3��1���Q�rP�����q�oVc=����������>���*^w`|<+����:Ү��y��#:λ�N�u�`Fk���2a}�F��7u\h}%h֜���N��m��܄P�}���WS�VA+F�]\���1vǎ�;6�����8<"�_-�~�F��qw��[��ᴭVJ!h��w}���uZ�i81��θ�T 8�s�0�Ӊ ��̫0kҝz��q�2�(��w8�\^�N�Bu�l���\N@�<&�,�(J�9�N/H�5�F@$Z��\;��E5��������T�ЍTp2W���^x�g}�!��m&��_������#=Z��.�/]�ӻw���vPE�jԣ�R��|��k�΋�p��q�8�q�Y���L��$^s�t[�C�cԚo��c�pv㱸9,f=A����aj2 ;�9R�GcI��;�L�U��m��CO����n�ǃ��'����W\��������L��/;�1r;���K#�'�:�LuY�{���EPy�n`#�g���Z��ra����Mqy�CJ�G;7=��v.]�X}�����f'��BU�P����Iq�/T��w�]o�9�[�����k�;].��(�o����
0��t,�5"3ֶ�	r�*�5��8B�ޭ��L��_ީ(
Y,��.�w�b�zpXSB­Y��eZ�Pށ�7"��1q�����������뾝RC���/B�<�a�<��뻨eu��b
�R��U��ʷ
	U�� �%^*diű�̮\)S��ܼS�Rfv��؟|
Ѝ8ބhחKP-L�ن����|$�#�(*�Ҏv�&����4w�NF��t��#}�J�U�!la�K����@��˦md��#b8�Ο&�f�3�_���;*@8-R7b�F����s�F�9s����S6hl��ڮ�p��M󊺫��<s�i�
F����@�DV�G�nuE��ҝ��:���Q.������a�tp�M��3"��Bz|�0\S��`L{m�xO��|y��[�M����e�J��*��ǁ�u��������C{��Յqx�v\#Ѱ��gv��6�͍m�����g����r�0M�@[�T�U�[����St���3=�_E:��7;3yr�Tk�h0���.�D�K,ht�39�}X#G*�m�Z�ugfq��)c�z�Y_<x1W�uX@���^�@B�C�1��\Q���릵����]^��ւ+@u�H��OL�>1ԩ����%� �Y�d�V:ʡ�2Oi�� �+�Q��a˭e\�������b��  _�{R�S�[T6mʴ�;�Ӊ\�����W�.�v�"0�Sv�.��,b��ad9�t3K�_���������t����VV��A�OI�� �L}
��C��v+�eu����n`��nek����x���us��Y�0s�i���gj3���ŚB�-�Q��{й��uY	�<f{y�]�i-(�V�<&��8'��h�ue|�a{,y	�,�)�]�5<OE+�y@�d3�YeR����
劕�ّ�d��U�K�͸z���Ő�" ���iaB	���;���Fy�b�҃�������!��h�*�w�VY��D�b�	r��}��H>���R����zh��fl97�9���OV�J�M��i�u]`6�[Po$"ڞ5��t-��l�Z݄m��ۻզ��D�z���[��c�6KB}�v��S�&1R0���(��+UǊ�C�K�*��������gog�n��
P8�%ox5�'s�d�pPܕ��TgPF�M=�����7�N�tgs/��y�<F8{�ͨ�~t���E
9:x�vU��@��~`���|,k�����724��b�Yv���	�<@h'��+�x|��`�sg���y��'Z��Z��Zp�Pi5����N�y�s�=�����"�hJ�u�U���V�����]O������pN����qÜ�s��^[���Y>�
3���ss���b����7�٪"��9�S:ګ���`�86Ǫ��ӫ~D
�W��}zh,���;�oś%e[�M�1j��S1S��%1�&��E�E��'�)��U����^��LH�[Ǝ�&R%஝��{�`�Ha��9���jk,#r��u3�ī�:1���)CpL��j��Q���OutX��O����oz�ầ��ꊳ�15.����
��2�8�����εow���Zx�,!⼺�M(�-��}鉣��;�U�L&�3�q7-N3ɮX����1GL����k�Q5Π�z���*#=(��'���9�687�A|l<�/XƄ$k�wL���ȑy�I���ʞ@�zہ&é�<�kM�3��\.�l-x��Yy�z,�޵fzk�2�X��WԼ.b���j�>��j��OG6n���95x�2ڝ\+W���h��'ҩ/a��N��0�b���r�˸IJ4i_vXZq��ݞK�7e�[���C����5����NK��o�T�2J���b}�+粇z����I��9�;�+z�����e;G[}���z9�����qL�Cj�+H_,yL9��X��8^ �Gs�Ҽ�y
�U�VJ]����i��vOfk��k7m9�%n���F�6�<K��{T�gQY}�0J���:_lG����R�N��b9ou�Ү��$����U�V���m��U`�S��)V�=k:(ް0���w\�Sg;�w�ˣdWJ]�m�,<��۠��O�������y�]^�=C���ݙ}(�b嵩��5`�qKy܋����c79���u{&��Թ7��u=�4#�<��<��X���3����>�P[WZ���ҥe���I�4��Z�$��ת̽Y�z]b���{ݣ���V��|�k0�%���B�k�ʰ���9�[ln;�;m2�˷�.�i칹��fp2n4�Oq�����oDVmaqD�aK�^��z��m��5��qd@U���f�W<��q��9�6���o�q�zM��wF��4D	(k�/�ůL��T
�u�7s�sj@a�:7�v�6ʗzvئ�ZP.jؾ�?J��)m�:��"�,χ��^�yI�	�`�:�y)�b�dQl`���D����)}�K��;\��4@�e��o[�j�bP��9L���P%[�+�l�Y�i���P\ɴ�4n��pz�vc�m/'gw:Zq��!��n���Җ�C}�d���c��V$�Z���ݥN��q��<Ct)ܻ�]+�6�痯�c"��T�V���Nl�B��@qŵӒ���T���IA�%|�>7��ճ1
#o9�洇{k��u1�Nb��2\)s��<8Mo��f���r��yY��T<��Q�y��6L�X�q���E�	��a�$m�����0;P[��tprRU÷�I)�å�Z�I�Ц�W34xp.W[�C��qdb��ifM)VyPhѲk�MW���|���&:�k��˘y�݇��sbg(����$�s&/���4�)7ur�>�WJ�]��@��Ѹa�Ft�Ukb��/��pn��+�Q�d��˰���s$���1���������۰(��{ mA֖�o��wz\��j�{ ��8��<�Y��(����B+�@ͫ`����ۉ<�st�a�1�����iV�Qlh��Cs�T���2�������b.�ې�H��C���Z��a<��ջ�09y���z�,��L�V���0���a�Z���Sa�=8˂��.�SW<���]`��*h���	N��v�n�l]��]��S�J��v��8�ȕ�5&̀mk������MiwMi��b��
8�ᒝ.�ޗt������V٭�o�@ǔcӻf��VLq=��&÷�U7Cy;olj{E�L"�[��C��m�p$��_d�������ee�#;*�B��!f;Q\Id�z�Go���_C5wB��g:�6���I�z�K�L�N]�Vsm�����9�8H��N�D������ػ:���[m=�S�B�W����ڴQ�ǋ$���=F�7�������1�����bQ*(��Z���Z�R�왎e
�B������Ul��e��4��E�
�ڊ�U�YQ����e��UQE*V�e�h֖�+���j������kEKm�4Q�Z�4J��T��)Q`��TP�A���hZ�[X�E++)�����%JҖ�[*IF�+E-j1��KKEkieZ��-�UaYZ��m��R��l�-�(YZ����KmeA�(�[U*��cZ)1
�ĪV���U��#h[d�3(�-Q���E�KDaKiJ�h�B�����QQ�Uh���1�*��EYD�T��*�Pm%������E�iYmKV[(�bP��kjJ�em�E���PT�Q��)h��KZU�P*+�Uh�E��J��J�µ���T���[
�mF����j���HIc�|m����$lmKB��[J���(��C^e,�߬�-��QW�w��Lo:�Xe�2�����En���m|l�֫$YC6�bk��s3�>6h`�]8p�A�N,j�\m��Tᴫn�ǲ:�m��j�9,��a�s!B ��n����%�s�����F3gR0p�9���Ъ�X�jƉ�
<Fb����^��E�A�x+�kێ����8��*�\����Z�R5`9L#��L��⓺��OyÄ#o*0mm���H����!P�������u9��z ���Ђ�9yQt�}P��`A���*��
t�No*�p3ިӮ¯q�����YP��8f�Z(�)rɞ�G$���Ɓ��R��~�F��.񕺷�\Z<�X)�^�ۗݳ��ht(���b��֝
�!g&�I�$3*����tҍ�����SP��{Os��Ì����ڥp�T����Y�Bh'פX��{B��W@��f�r�6Gj'=W��������;jI{��Q|c�CtKҤu�˅�L͉��S�w8t�|0��Z��y��Bc[^��J��u����MN�R���{���v"'�N'\l��}ѯ���f�������ͷ\b�E��@���؊ !0�0�j/��Ȁ��{�J�l���d+��qԩ�rq��Z����WW��z�u��(>�|F�x��w}�He	㳏_&w����o$N�q��tUvi_�ݛ�LH��E��k��v�
���Ĥ��ң���c�AV��~�f��cv4�T��E��r2./�#{b �
����<˯{�@��ѤP��5+j2@��FMi��bp�nI΀Uqy���o)bf�/�m7�}��ԡcǖ�O��'�1:W����c�J�c*j�>N��H�ۓя�xO�U���K���)>�b�y�����a�B�����W�9�X.�̽��������(n0(�#F��y�Src[U��n��<V@u�z���A�]����x�E��O�+K����Z�ʻ�T�}1@��"��i"��k^^�bb�eaL<v�b��3n�������((E�qΆG^�{j�5e�,4bf����l�t��"�D������dPxG�|����`�����5"��Gv�p��-�^���@�!�bDX�U�����䲬�=u	�x0��]��<�t4�r��o6��+sB+ #�X���������>�k�>^R�
�&Ʌ]'� !O�{�o�J������� Ŝ6��j7|,Z���9��\��3���p�ƻ���qd���6V�B,�:�����-ɧl�l��4d���t���<����s2"p�v�ݫ����':,w74\���L��&B��5�
��'WD�,�}%�ȏp�TyF�L@u#��ہEQ3��~D�W:���y�	:�{X|+뽸+�0p�:𕳒Ә19(��cJ#l��(��@�w���4�(WSϟZ��(���wy��R��h�d:�.���'i�Z��03�K{˭������ڷ�Q�g��
��fgU�*'7Ī}+��?��=f#Pru=0�������P|�HC� ��]�gI����,��������n"��|����W<�u�A3������v&E�w �|S�֜t�|�������|�_t�f]o���D��֊�K��1����r`�q���ry�ݥ���-J%¨`�8h-��LSͨ3�q�bt�D�6EΙH�s�5�-
98$��0l��AǨl ����i���N��A�b��*g9��"����kW����R���C���ᢺ�@�c`ߤ϶vN�e4<�Ϸ#�r�|��-3S7�`�75�uVL3���4*ʃc$"���@k�]����"1J���1��,e7��n�ٺ������-�R�;4'EG�L`� ��E��c�<A�}��NI)C0l�Cj�]+��+��_S��c���i��)���.���rc�5s�b�)Zu�+�M��|5����#�7U�1	�����9#�n�y�N���Ts#[��Ps<c��hS�`��ZLP��8��3�/C���F?��o�uM�8k���>�<�Y���q�t��8�H����,DH�mm	�����]5����PE��=��qU���@��^%y%��x!㓥Xu\
᧕[���Mw�<��w���@=�}T�8���,��˰W��r�3��*��u^�	��8��Y���!�ʗ�YP�ܘ�s���df��uiK�:<�X>��mE�y�x�J`��֜���0L��(�[�8E�t3,����4J;����i�^"�D�e����`5z�1�ّ6_��-O�T�p&���6%���0��k.M�r�Y�P�uI܈�6��$�Tr��$1�0�#OgD�g��N&4O��^E	��X�p`���=������љ���:yn+Ϫ�ӏ2ю��>ߑLl��J���ތR�^�#8ס�<nq�}w��5�,Zչ�A��J�`��Mu}i���W9u�wArz7`[~f�x@�T���l���d�pѭ�D)�w\�֍�Ī��:[�UC���z�Ӛ�/3t�LO *���K�;.�'�a�4���e��&����;�*���6�e�ԭ��ǀiV�N��wa�z%�,	#��H�vv��&��bD�w�3�ǘ�9wP}3`�cԹb4��\쪎�y���gG��ʞ@�m��n��Yʪ�KE���O��9Y��`�9��ڜ�Z�����~�_R��.�΋������]�d��F7�cq�Qǣ�.�߇;�?����ӥ�W^Z���ч�o˸[W�)�S9��۽|�J��<�F�t�:x�F�h*�Ӳ��d�A5�u�Pnj�V^�����]5^�)��a)N;*GlMr�c X�<E�S;b2Z��c��Ҫ���������J�����luN��}�J���*e�Xz#!A�F�9L��^�m�R���{%�P8S�:�b�;c"(\S�ўQ�*��5�Q�Kذ:���}���mp�]�\��]h�H䒋�>���8�������|�(%��C��ϥ�G�2�Ʒ�@���a^�b�bVi�5bT?Bx��ƨS�1F��l��������<7ٔr�$-��Pi����_Cu�j���W\e/��U�s��k�ۀ�K��m���n��ds��b���]��]F��E�T�˳�tѣ/PaPy�l�l� M3ݫ1j$�)�e�2�[gVT�1�=�8�[�ٲ���ȗdx �j.�3����Z�uX���O}�ӏ;r��7��+���qPy���d��� +>�k�����F�Cv��G1�F�%�;��KtZ�`f�	��^�cf*F��qӘim����-��1!ʸ��+�Qu�<KrKҤs��������v)��ø�1o�It�/^�8h��`āj��MΜ���\�L΋�p�u�>�N��n��w]���%ۜ�I]0��oi�����8**�U�DNKb(p��d�:��q4���s������� ����~Uؽf|�;��]���>ت��]C��Pz����u��j�K���6�����
u��oኬ}��Hw]@�Yt��i�� Gְo��B����P�ݕOJ��X=��ԡcX2��ٟ2]���R$�Mgx8a�n��A�l�RZrv6Ô�t�}ϫ�7v���;&�5�k����N�&�/�<J��g;�-�59SB��Fq���+:�;(n0(��4O8Oض�A�Q�y<t�87\�fI��]Y�P恧��r���#��\5P��0�'J���j:4:�]�L�"s��J�j�{+hu�}/A����«Q�J̓�DN�^^�n��%��{�LJY8N���J�{���P�ñbQ�l�Ǝ4��{��>�wl%�0����3w[�+!fٺ�4���im*������ևZ����r���t.l�����cˁdFԒ�WPܣ�B7P�O(E�9ybЄ)͑�v>3
��m��{SR����/�?�����B�kU(R����[�F�)�*�]��F������S��7#K�H�R;��b/�ԬP���U^Kj管8�i#����w��=��%CP8�X�,������F� H��Vr���91�$#��M��K���KG��,�]>����0\
*��MC��9�l��s:��S�����3���SQM��s���fH�Dm c\{l���l�r�_*�<}C���<k��S�<��ԛ�hW�!�i�J��]j�<�Aګ��'\Q��@���x�Rs<���n�VF;�[�mR+9h����pMюO#c�BJ����]�~�jc� u8ݍ�Rn����pL	1I�kn"ġ�Ҿ���W䫡��������5͗���-I�[i*7`���Si<�qx9�Ns�3ǬFW�<F���=\=��K�q�i�gfmХ�i��YV�ϻC���RQv/U���p=_b�N�udJ�ʘ=8<�b��.��^�8��j5��.�J���%8���З_a�<�ѝL�&<�HC�3���#���:�;�A���u�N�B���Ԓq��o�t���wMʫ�ؙ��ǗG٬5,.���M�c����3X�1P��h��&�v�t�'�m��ӹkK��y�w�PR���l��>r��s���TG�N�R���N�*7Aҹ�ZD��Ԃ�=;�T9$�A��P����y��~�V<+��}�:���!ʹ��H�K�}_o^D�Ǿ�&�1[��m<ЂW��r�RS�qX/���)�
ļ@���\����qA�����o�l#�[��z.��-GF��T�1j�X+ݖ��:5��)����#14��[���c{�+QC�3"�!>5go\�J�!����j����3�]T9s�{����M�4RE���ڷR2a�ZI"���`8�ob�Y8�g<�V�m({��Nu��J�*�v����a�T�ۯN�C0�������n�v�ȯ�!�$I�\����+=i�n.[y]^YZ煪dD�0Q�<�Ř�m]�m��Uz�����Z̽�YQZ�Ѯt��W�J^u.~��{s�~t���c��$�xT�6�����iܔ��'L[�i��k�>����� ���t�v��C�w]'R}gc'�f�!���"�b�y�흟vr
닙Ԃ�z����}��s�v0�~��{U��L�Fu���bY�t3	�V��R2�L������ќ��������<��
A�D���bc\P�^\U��l��T4d�]�&�O'ǦvPECSjh*b}�9

\�xNk�<�<؝{�p�r�����Ê��j�e��"�D��#:����a��ƽ�w%�-#��H��Mｓ���ƻ~6���O����yOm���Z�g� ޼I�USkf"ZJ@</TlVy�۫�ҫ�8����*��#��wc��J%Q�ɫ~-��[�.�X��͸tn��r(E�.�.��|)YwJ��J���v��F���f�k���;��4<���:��T�H����%��9�U��1��9Iu���f�$w,���-S��M>�y��$v���a�D�n�R�`*�C_O�[�)�G����/+�d]<�mIvI�Y�k�W.��m�gN���*�u9t�{"���ɀ�Ro���Me����j�qf�1v%H�ojSB�2���Ӫt�BᲱ�Vi��/y��ƻ�:A't�YL��/�Z��y���ys>�}쩎�J
�sMޫ��w-�Y�����I� ��2�u֤���_Y��7Y:�.�O]��T-�ߨ��:߶���U��=\�]�D\m�Y92���{#Uʁ����:��q���f�'$�ez��v�Z���W�זs�V�*�m
n���U�fa=��<6���R0�I�S�0��wOiP��1ܘ�&B�eD���4�3��|�0�)͝�ef6����K����̧^�*z86`��n.�V���{)�"=�ko�Tdɻ3N?|���=�=�(H�ى�h��p�����Y���_7ݣt���:3T1�5������+V8�\�bG#�Ociٍ�;�y;���"e�ڲ��D� V���*gmM���� j�s���q����-�oŢ�������_R[��gk�ϴ��Xi�R�A���'��B����F���X]y*�,^z��W�N:�Β2��VMn�����E[���R[V�'efnW*��x��>����ȩ�!��HZV�ŭn���3ʡ�Zs^���`V�z�K�{�Z��{-�@�"Gi�SJm����:Q�ɞ��Z;��W�G��ޮo9qv���,���Y�n^]<rҚ��Xu�y|��yn��t�oY��
c,)I`޽��:GV�DBm�X��Q���D�v��Ω��5�����s-\���x7)ѳ0�m���,�U4�D��Kr�$�񅚰��'�N��`���������Ɫ��{@�����H�{��7Cr�����WdI����Ÿ慛D�F���G�V�G�s���t���)~�|e�'}h�o��
1�U����-ٻ�-q�# ��w�t��h���pERw72>�U�Ut��BSO�pl��Pǁ,��ʃ��;{'X���\u�W5*Ŝ��q�a�y��M(�G;ve,�mEe��3ga���ގM�u�{�-���z�-�f�\�J���?X'�ـ_M	h5n$n������e�*�Q�l+�,��i.��x�潩ˮ�Q���2��c�x[h;�;I9$�J�u��r�G����n�m���p+�X��N:|b��n�.x`o:rs|;G\��Nu���A�%}W�y�rDT@�++�Q�d���܊��H�,���Ƥv�ٚ��r����j#X�F�GcȨ 5H��p��hVL��j��y��C�=���R�r��\��5V#*�U��vu��a�9X��.
�[�]��9�5��KH3F[��Z#,;��B�
�9_A�\;�Q;(Uw�pL��Jט�J(�[PEA�����1WE����E&�Qբ��i�'w[�P���p��*`���V"���[��3�S"a�ڈuΌ�Y��V�P���
��L�
ԥ�kO�3fQO`m�wWK,-g"�/Fn�ź,r�&�<�u��T��1��m[��#� k�s�r*�R�Nw*97^5��o����F�5�Y�qYiV��7S��"�z��@�5r�B�k�]e�s%��MY;���<�Tu���[5)�˨~q��{���jų��+�D�r��c&4o���ǫ,�~'32��ݝFQw�M3t���+�R����w׏����h#[wK,E�9sl��ڙ�[��n\33�`'y�D*�$�vRV�/���[1]Cv��u��Gζ��G���b�Gq��t��|x���il�c����7��T�	N�3��z�R��|���$�Db��=�Q��7�库}��܁)�t�]͢ե�w���ًk�FD67�6Y��iq�u���<�ܧ2\}ݲ��ɛ�S��!me3.���׭��G�bȒ�#��hF���U�mE��
ʕ-�(VV[[kYD*E*Q��F���U��DJʕ�ֶ"��V(�[lm)l��1
Rт5V�m�-ZU�Z�J�F� �AKV�[el�e���FҪ�el��kF�ʕX�P��F�D��cKA����*��U��+b�E�+�V�։U��ҌJѭ���-�)U	hժ��kmEZ)TT�*Z����-�Q��iiZ��--b�Q����*V��D�4���*��E�հR���"�TV�iE���4�%���kK-hԵk[*�6֪4khTm[)TF��KmJ�E[-��mKlQ�jʱ�b�m,-jѴEh��j�e�I������@�m�&�����EQb�1PK[m-B�X�Z�E�kmR���Q��Ҋ*�%Q�Z6նV�P�ň��kKl[h��Yb��[,���c+-V��ER��[A+T�me
ڕj�-U��-�J��R�تVQF�iVT�TX(��#h�Ow9I��K��t[|$�s��\^��Ʈ���r���Xwr�n�<R�0�X{/n&E+<R�b��*t�\b�Ğ��M�W�p�
�W>�]n&��=5v�����-�c.��Ѹ�o"O7!pYZUI��mtPw��=�6"*�Qf߉�i�|�0�2E������j^������WlPm̰��`��R�u�y�P�3PSx�V(*ĤF���N�t��Pk4��qz�Cܠ}OT�V%�=^�`� �l+��>��U�Ut�_�r"3�T�Vg,C����;1;Nˠ����82�Z�=`�΅v�WYy�r&�_f�)\%���X�w*�ޜoz��dKl�@t$+#B���!�u�.k��7���J�>������w��q��͜X����}I�hh�Ԕ��'+�ZNj��F`VޓqoܬȆ�l���ryKRi�����I����(���-Zr�=�[��5�c�!����~,�w�=�^�wM�^����1��|ݘ�q�n+�luaeܕ"�DAˬ�{Q�׽7g	R�ڴs�v#�P�N���Z�.n͝H��K����̩����xt���c���hG5F(Ŏ[ƣk�r����*����	�qzU����G(�ȹ�\��r�nЖ��ꚙ�W�y�ot��'ͿBx7[{/�SP4�r�]b;���.�F�����O[�c���8�K^����Nn9l�oұ��|�5U+�CCs0��Dƻ�������V_�j��N�3+���͉�š90���ԡ��ā�ǩ;u\�9��^��
v-?��έ�A]^��ƫ��+�d�s:���9u��q4i��^�]v�zf���ϹI����j��W����E��P��������k�Y{�$��F�5;�����Ub>}:���鏫�T�zj�W��=��z���D��ɋ���A>;�u\�H��d	���k�k��#2o�o(lʗX��ӿ{����gKH� ��Ӿ+��)�
ļm#�b�G<���Y�)��RS��}ʇ>���Q�<�x�
�mN�s�z�,y[�'F��k�IG�|zj�uN���޾ by��8�V�Å{}���N�Y��wl٭J���&,M�x�VoB��9֕��o(;/��__T��
4�]y�ji��sOtv��݉��+o;���9m	�Zĸ����9�l�7Iqt�Z�-���2�ϩ5s��˹P�#���*+��2(rB\M3}�8���~S���Q:��6�׺�����-7x�&��D�k������Q�ÍB�7��\��fnuN���^]m*���L�����q-��a�ř�"&�!V�)��	�p�لŧ�v�����6Y0��gkI��͹s7C�&6i2�s�'-X�q�W`�t(�]��f�g4�w��i�EƎ����e�%��� ��t1�ҁ�8m�\.rN�RV��C���� ߺ8R���87!A\�z)˚b;\s٫l=��M7M���[�o��߾IÒ�ٛj'i��{�	�+a��;�u�m�y�+H�ґ����������S��3�� �*n6F6"@��1#��{V�����%m�=%��ؖݘt.�1�*v.���V2t�ȹyCPV�q6*å礛�\�,��19}�����ӣm���w�揼U]���Yo��lT9��#Ӵ���I7H:�sq>z����΅���]���o��w]���1�q�L'x�m��m����G��Μ�J��.ໍ�֊a�Df�yL�k9�\�4Sc��jK������7j�Y��ҥr*-�v'Ǟ�v96��4��w6�m�ƺ��UI���(�&C�o�=O9K�EG�WP
5\b�����N��{-���9	.�Ƚ�ە���W��;hȹ�k�۾G:�5�dt]�����J�;�[Л�S�	{�����18�z�3�z6�J�j�X4�ص���}k�Wn�<|����֦���w�/v�7Ԃ)o�6��(��}:�Ƶ�:�'_�;�z��".�m�cw�vCl��t4(dj�s�%]S&ul����6GLT�E�M��n�X�>��T��p2���BF|k�ڑ����}���Z���m��%)�W]��Z�rb�2*'����j8ԝ0�0�e���XNL�D��ɥKhN�	|x6`�7�+j��KJ�5g�v�E��
+�=�]`C5g��H���Y�fw-r�8ӻ��J���H�nbn�rMs��M�HB-�zN�/���$�] 8���q�_`��:��<�g��);]M����gv��������Q�^,��-,թ!*�*e�un:��cֲ'�I�0pnGl�0ی.�V+,!}�m�L�SYA˱=\3T1���=�y��	�P�lO�!;&����w��]g��S�Z.n7,���_+:���Xܯ�^\nB�q�}i�m1]@U��vI�������ͼ��VF�n�(fW�i�;N�'J���ȳV�A�����|�ey �S��ں�N��En�.�lC�nnC1����-���(���X��A�AJJ�Y������M��3�lCG0�$�s55����5b�VH�ZD�}:�n���IU.綫�&�l.�J(�>��:�����-�=\�X��X���к6{:��U��8Ӿ%c�!���k1�dEs���s���>
T�s��h�\�����su�훦󵴘���w-k���,��S�
<�<�Z1X�j�������=�@r���W�?%@m<�d���Q�4(:T�?�Gdb���c;ihݻ0���p�(�U��\������|(&,.��X���2wf`����]�o�jϟ]C��(39q�&�#i�ucvԒ�송������8����|x7֢�it���*d����n���c��1Q����!@�O�óہq�ُ��-Of�{�.����ʴݽY"�XA�5�ܪ��K[oD�N��B7W�ٟB���yu��KS�Lu{���&��>�y;Y�$��{�	��D&���5soh���ө�f�K9��������aѳ!0���J�uBg-\��7��md^;{fr��V(;�}i&��m��c�$7�á�Lv��;ɚ�1���.�t���cU���g4Mmʞ�|��Тc]�"x=&���9jCП�&+{7WMԫ8`�����H��b�J�	�Zj��� 7^�}��4g;��Xy�Q��*mu���:�_��E��c�K�lVA�S9vP[n&��1TRS����w�zy,����`�o���qu<�A&�[��'���)����ݨ��)����uc�F᮴P(9Z.�N�[��kvaR�]�մ�s)&���w��m����K��vCW)�j���&`B��6�k��񌓩>��V�u�p��,�hf�=��s�N3���|:
��p}X4vt���x1�Q��i=��ٽ�Kr)���.�lC�jUH�Z�-�j(l��b4/�\��x�9W�	�4��U�[㕮:���bE�T�~H������]��-�������c�t��uy/��_)�������)�
ļ�Rj�|�0U\^��}N�+�s��wo_�7�(Q䨾����z����Z�C��nP�\�i7�˷��Պ�W�����L�17T�.��0�֥�bb�w��3�[\/ue�7@-�ޏl񍜆��u�	]Em�Us��t���XY7�=�}�SK�ղo5�v�h�������r�_ki��
���n�ʸT3	�OF�٦(8u���|�i\+i<x���x5N�&�&:����
��K��h�F:{S9(��W��NS�0�Z�P�=k=��O7J�5����ص�4�X+��`���2��*��x$�������d�Nu������z�_����m����_>u{�F�P���ժQ퀌�)���'�q���D����L�n�&���h!�ۖ
޸����B��|�{*�G���z�ɘw�^��1�Z�[���8R�0}�Y��]X=I�x�8[j�wh�r�Ǉ���|�m��;��[�f��ϸ7!A\�{�S�4��_�<�肮���u3*�+1���5jo�8m8ͤ#Ԅ�e[$�m���F7�(�c�#y�gW���˙�sc*��V1�1 u!�Ңc/F*q�]�鉝ʫo'��`�}bu���W,1��^�ps�1b%L�̂k��V����L:�/r�t�V��V*.�lC�jUH���uB�"�ڱN�A�"!�Y�����N�r�M�߇5���^��Ca\�I���W����	�-vk��r]^I=�:J:��m�}Oy6�i��CEm��yUMnf�Q�:�v�i��ˀU��{U{�6.�����!�Ԅ�S����S}'m�n���TW�`SUB֪��t����m,>y=~��#���%���J��\�=F+���Tj���V�yÏh��d\r�����x��%l�Wm
Kj�f��fJ}�)[��h⚲�͎�p*�$�^��	�\�^�8�W��t������ݘ���z=ޏ�f@3e�����|�eGL�\B!Q�Yˏ!U6��Z��iv*#[e��hW�5P:2U�T�շ�`�e҈�׽�Z��0������j���}I���"�m��\���茺0��Ŭ���>�l�B';�m`J��^��c�ܘ���U�*6��K��U��|�T��P�g=v�j����i{F�l*�!�B����8�'��۵�m��QB'E���f�Q>�Ol���A�vr4��vzit��7zF�"��D�(׷�{s5jlc�8�$m!1����5��Rc*w�:�r�+:Ɍ�]{� �c�lozNT�5��)9�+o�0�j�/܌x+��nbt-Ѕ��<���Y�g,�l�Z����򋘼�:�\���XR�U�}���M<�@�^.�e��w�5�d(�2�)L�K��J�\v�7�����)*Mfkk�٠�H��
�o`z�ɺ�i�X�h���ӫ��;���� �k���q�s0��R��W����M�������u��K�Բ`N$q��R�χ�Q��UnU�w�oWl=ͱ�ö#�y��͝	6���Ub�Ԙ�e����E�Ӻ�-M��j��5NVH�ZD��A7�S��W�5��05ք⴫��̠��VC3�~=�E�+��?.��N�I��Gsuv��;m�'�+����,T��������8��/���[=`ȶ�W��M��9�kyQK�z�j�IP�7�$=�<W�-q�Ѕ������fP�y�����"�K��S�ԳP����-���x�T� ��l�BK��lR��۹1/z�حn�6B�����j�Z&AmU�J{�P���AN,�v�8!���u���vT4�1��oBͳُ���3*�#�/������P��2��u�e:�����ȤJꙬ���7լc����	�:��Z�K̇{�ǭ\H��K�q��ֺ�����K��HhcEYA��C��D��N<�Lթ�zG����X#�+
���!�]��.��=�ʎ0D���t�C����5��kY��j:v`�sF��2�{j;�i	�ׅXRGgBvLÚ嫷�Jxh��ݺ*�4k��)��4�;�������e��j�cT�,;:�M�gs��*�\`StZw���o�:Mv�%w+�c00����\+��M]1��%�h��S��C���q��ρ���<N+ݘy���vR�q]u2����L��=����.���5O&x,�W4޾]E,�n��}��Ӻ��ǖ�7N�J�[P�w0=�P�J96]�x�Ȋ9�a#}-mh͌��T䀤�K�o���`weQ��uy@�3����g�8�K�Y�j�!cz%��Y��L�Cgs�8�xԕ7�:̋/H3G,�2�3�ge�W<���Ѕs����ۤ�ǆ��Vۮ�DfJr��j��k�/��v^��0j�|/D��2�IK�C(�lYݛ,t�Ea���n���ٶ:I���{;��4Y�����o��8���VԺ��BK��%�u��η�h_5
]��7��^L�>�Gq[=OB�r�2+�=t]�ۺ+���p :��wZ15������t����K2R%���3��3K�Fr0n���r��Bǆ�Š��5_u��8�nlɎ�p��^j�K�]}�kT�g�nٲ$�X j�ʗe�f��.��Kock,�e�4N㷠q��BWb��Yڛ���E�5��a���5�1���ݾ�PZB���Z��3]E<#:��P�WJ���w����F#�E��N���idmf�,X[���ݷ&Vl��
��ܗ�>C� ����:+-O6Q�)fB���e��H�ki�-}��8E�3�b�;eu�0;y�_2��vv"@K�����
�k7���z�J̺N+���|�k�ڛ�S8)f���S��Het��E�vc��N�Ĳ��i���Z4 BoR��v�T!�֑:E[������a��F§���.<�ʷR�U��脗j�f��Bd��f�h��h��.[��Ά��F�K�حh=��-=\F�S��b�\Z�s�YN$rΈ#U|t���\U�u��Z�݈n�]�����6�6��>�κD���zC:�Ewƙ�7�n��*��^P�Y�w��/-,O1V\����-I��,q�"|���&t{ݲ�盂�V�4��]��]�Y)�CT��f$7����t�N��z���(�\_
Ÿ��ٝ��<����H�u�tժV�Ys�K��q ��n�5i$fGR�<�N�Ŗ;�/k�շ���R�2+@w+q["�f�p$����{��[4%ꇫ:�v�y�Q�"���"0d�����*O��@�+oU5z��
��p�U��uծ-�5��0�7`,y����t��'���[gπcG�t��-�b��}CaA����AO�%��w��qv�JÖ���qY��b�n��d�)y�����!"K�PC���]�v:���2�8����Vo���MM����7mXQ��ٍ��گ���<���_R�c#��T�m�˫��
ԭq��N���OP�6�� -Vŉ��2��ŊR�c-��m�XQQJ�b�*#IhR�U�V���Q�EZYeU�lJ4�Q�F*Z-[h��l�����(�VԲ��(�Z�D���D�J�eD*R����*V��F(��-l��eE������R�-ml�D�X��D*V�-Z-�¥����m�U�%���bֲ�m+X"���KQKT�m����6�T(�Dmh��,�R�Pmj�DAU�*�h�J����db+�)Z�J�VZB��[bT��ڂ�)h��bUlQQeePYZĴ��c�b�QR�BҊV-DV�V����U�UUQDDEJ�m�
ѭbVԵ�J�kJT���mʅaIkB����D��(��-[H6��6%H�(Ŵ�����KJ%��R-AV	m��E-��eF�T�����A
�X)��j"�bZ���Uj4lmTTB��Z�U�hڪ(���m�s�-�}�����W�:_o&Ұ�|���v�&e���/�T�7��ه��ۈݾ�07�\c4�c�����태�<����
��Cb:>1eyS�f���c]�"z�^�����+�37���5�Xs�mvW������1<�]���<�y��0ӍlNӱ�*��Tj�0v0��[j�,�ȼl^��T�>���ۉ[M�e��B[���MT�B]G�m:"�=��)�T2.@�P���{�\E�+��|�sJ��9��P�h)�ux�A��H��z�j
�1���lMc��)����P䲹v�7�q��*����(둝�L�ãrhA&[����UVΘՙ�K�?���̏A���?�+�c4N�2�tԕ�]���N�^�kH�KGS�kT�{!�oXT˥U�J�,�?=�:�w�N��p�g]E��ۚ���w$;c��m�jM%�fWu䧎�KZ�l��L�Z)h��"1Uk��v�y�n x�ī��
[��"_wA���w,%��v�"^Q���as�U�����.;;�۰1;h�=�S~z�G���hT��ܛa�jr�<y��ŮO^Q�l$H�p6�,)��]���um�=���KV9Ԍ��ɻ�V�r=DLWh���G����s#m��!&P�:�e��N�ƭ���nch��kg"J������}�St��֙K� ��v"p�+��٭]5�q��;Y�#S�P��wA�L>�[C�16�-v%�Z�,�s�b�mk=''	,=R�ވOG	s��j�C<�(:�V�#jo���W��!�u�]S����)�(O�7==�Ǽk�ҵ�l�z��0�n�9��FǼ�m�Y5-�[q#e����28ny$�fz��z���v��3��\��8n��:��W`��Ҋ�!��Z=u�r�[�����:ꇳC�+�5�s�Z����򘠷Z%�O9��v��+�md��t��ent��x53�·��>b:��4SS{^�mw%1lU����! ���JJ�5�~mA�y�;W�6��6��J$f���}z%p#��Dހ��E���6�UK��2���J�E��==4��R�u�}|���w6�uɝr�y��t��;��/Y�j�&�I��,�޳c��6n,����k�p���ZEԂ�zGe��ܙ��&�<w9l	�R�������Pw��q�k�9�IJ�yj��m���񉎮��,��T+���/6��ÅBr�"}i϶{z�����5��C���/.�����'2�XY�9N����D��^jf�+�����O��ж��r����iJL]�S�����R��P�Ʋ�/�O�[Dvfs#��y�i�b���K'u�������l�@A+>!M�c��~�'��41Vm�%߸�5�e(�o1�ֵ^��V�,p$RD*�"�oQO�]������|ݒ���z��J^��[a=�Rd&ggԅ��1F�si!�����α:n.ɺO(��)�.@���l,ʽj�\m��q1(^H-�*�1�+�8-:�:3	��m=�Bx6B���.�/y���|�9�ì�T��Vg�ƺ1�.f��_Y���Ży�^5蹀̮�5mı�RﹰkYX��K�/i�}x�i�FV��q;wF�/1���EH�w������}cwGR|�{�c�����W���o�.�MӘ3:���j1V�"�f�(Ď���}
�z�9@řyں�����cw�܇�ԝd��,n8�zͨ�"��Trb�v����1���"Rs�ĎV*���|C�9�T*�;&ߴI���{�J�G�6���.*���>��KO�y;_��T��o�7�J��4dU�l�zo�jF\��d�k؇O���&��}�de�د��Z�t�@C͠�ƹ�
Uȵ�m��A:*{��]4gtmN+��կR�2��5���Rc.�^�ռ\��*慤D��u��F鼸�(S����&�e��B|��54��aZ;�M������f�7���N����L=��[�K�H�ͥ��P]HP��p�`�#9<��������Š��V��MP�N��K{q���+-�Ǝ����[s3�G�˃�y]}*\J�8�F4�^�˦�n+�zW�~�Ի�LTl���؎�}X��IO/����{�E���۠�Қ���ț��:�7���9�F��^S��/_Qy���'$+F�#[��'ܴ$ �
^m�e.q��Q4����Z��p��a߷�G��l�V G_^2e���9�QWC�<ya1�;Fm�����P���B,�*]��`�=��[J���Y�B�S��q�7d^.��I������p�,�f��Y ���[�����m�v��;����,����7���Cb���X%ۊ�&=k#��bp�Ts�3{���!�s���,5C����s�k�8�"iMNX������M��SC�Q!SS[LH�㙅�7j&5�2mW�W������S��Vo.|4���6��#6�����nf�f�̔i8����N�M�V^d�,fP�ۮ��VNC"�cbu#������6&j�Tw39o%��Ȗ�.J̠Xͥ;�K»�8�������,)ɨ��i|��M���F�/x��	�ɬ]r*ޙ���;C�X�Z���3=�;
u>�䲇.ئ���s�vy�Х=��u���YN@z��c���?MY����)����W|��" �͖%���g�� ��Kg��'Ed�Y'$���I�v���>��M���G�N�q?b���B�����Λ��q>ɽ1���b������t��K%n�Y�G*d;Y��ݹڳ��C���+�D�Z��\�\,�����6�_��PI��/��Z"M�Vk�u�3���9�o�z�tȉ����j�^����R�+�;���P�Wk����fk
M%���ѵ���z��"�v�]4�w*�n��0;�l.F!���a�+�%@Ҟ�Z'��b���Y��Ս�I�؉�zqw�{v����+�uh{��
vN�ެ��.�J�e�o�+:���D��y�l*��E/v�3���9
�i�Q�od�έ�֜D벎&[�`W]�"H-��916�"jv\e$.���'5p���b	���L�ż�T���넹Y�"y�U�W��
����ڦ����A�
|�Uo�U����մ�����u�U>��[��Ɇ�D��+oѯhL��[�"Ӊ�B$cc�Ɂ��4�z7Oo��]��.��q��K�&`5!f)̑jE�2��E%3/�6�/�Nb�u//�z�}x4��3��6>����ta#`wȲ�:�ˤ��=Ki�s7�z{�:�&�+�I.�ý��,��:�Wt9Л_P�d~W�e�? �	�߽�9�l�6哴(�w�����L*�#_HyN&�՘��{�*0E<�;�=�T)��;��gxzt���A꩐5nP��P����.�lC�j [Bh�.�`�Ź4s 6��dl�5�	*���S�5@���Y[E�V&�W%���fOS���r/���^O�j§>IJ�yj�`R�pܡ2qZ�>�l���bCw��O˥';�)�Y��_M�o��x��A���$�`uȊ~��Ti�	J �
�m���f-������w�X
���y��z�MΫ�k^7���p�!���A�R!�s�d^�V��6���wxa�֮;�n�[�;6@��^*"[e���>��q��tҸޅH�ە�Vot�������y׻ue���5SH,p$RD*�'��uc�O�[�3�R}\�Z�L}C����X�Y��J7�PR�����ISk́]�sp�bPz���t[GFI�9\-�������V(�;�ǒ�[+Rn��,��r�������e�D@��_o���/:���N���fs�˕9����TgS���9y����9������1�:�v }P���E �o�f�,M]�!�~Kq�鸟]���7:!4:\��:
ʘ�Sw�]k�tb�"y"�	�qQ9j���÷f�{�0�$�zQfz+���m�h���#9�w�S�'�zC�tc_�j���ϱlq�$��yh�/nR��'+�n���s0��I�Lo7*1]L�ӷ��璽!�#��3HLe������M�U�t|S·C؝um�nP�x���K3;3�9ڝ~�
@����V�r>�ׁSɠ�Lv�1���׫/���.�(FRX��v���k9ZT�rWi�L.�����h���x��^�꾨�����UF뫕*�Z�7��j	�J���I�,�������ʄ����%n������|�:����o/��v/��1D_��rbmkBqΫԓ#6�����h�:�o�����[�̔+�X����H����l�Q
��j�u�Ir�xE^���<ǫt��a>�%����A��6]q�3@MNg0WyL���M����kz�lh�o!�<j�;�I*]j��ZRJL�nu�U��<��BjyO��s �]�lu��E�h�w'�zT^��
�����o���k�P��3�Rn;�#"��3�qm�!ڡfhp॑���U\��:��T�oz�Y��,t^�Lca�W��ĉ^���A����"v�:dbN��՗M�Y��m��n�V]"�qf�\>*��E�0oG?m��U��k�G^��hژZ#�u�hI������J�d!���j��c�i�����5s�M��څ�ڦ��pU����g7W��g��d�+Ov�T:y�wSJ&v�G!�<�f\��s��XkK�����;�bT�n]�k��X��&�"�FKs�e	����\�w��"x{�����&^�ԪfU��ٙ�S�f��B7(_3����&��\iԄ/��;+c�{��n�tم���"�rˎ��z�3]OJ�\�m�l�C�
�I����e�O�e�q=�K�IQ�O3VMK�;�_7�|C��^�`�׈�/��1��u�S�/���]]p4�˘��79�	kZ�~��&f^�E!���5�;()۠�:��*�Eϱ�>��u1��FcgufA��A�Bgr���q4�f/7�v.�u�&ޔ'���Hjqj��=j�[�s�p��!>��V�o�x��H8�.Mt�H�[��ƗC6��{9<�zQ,w���Or�ч���.}���SrW��(���5E��=7Q��h����P���w.���1��k��m�^���poH�lrx�V�o���'Ш\F^�]O��R5쇼w�ɼΧ=U;]uW�c1>|T�M��`����!h�~��m��WoU�N�����'S��yuak��9*��a��,�C�*��U��Z��uMk���V�7�ֈ圳9�y����Mj�Kmu���
�dj�E�B�S�1�T�]Ƹ���ܠ�[:a?%�Bq��U��ZdH���
6��� z(�P����Q�~I�����;���c@��&�N���.=��u�hGm�G�E�rK.�(�X���S%ʴ�:�{,��BǕaϊ)�ԥq�Aq�-��q�����V��Ȫ
�` �����J�!^'l6�R�CkY�Ʒ/s��T�3��<��|�a�.��orKĔs7v�9�Y�)7�,<VR@���M��\Y�/r+�����X��V��k�m6�X��u)��N�[*�;U�ɥ���M�o*:���)�q�DUn�ʇVp�� ��J�E]ӑ �>
�]����E� �V���xr��ȫ4�A,D���4�ݛrwi�vR�ưҝҮ���x�5����i��@��W]�)�2f���:s6�ww^(���6�������S��<AoU�Q��uE���Y��*L���n²=�Ip���m=BT�;Vm���n��ȅ�;M�Y|�K�4��U֜��9���wh[�DwV�����Q�e�
����齤V�}�`7cpm�ւ��bX��	��:�$�SYyKz�oe��rL�rI��<�]*�%���V��$���N�=��N��e�Z�[ó`4sLd �溸:��h�NftST�=�p�9���u��[[��/�3z�GMp* �\y\fj�-�Z-��LV�����S�����:�E	R�4E��8px��t;L��J�p��\W��K��)���zh w��6���	FF������Xz�[W�\�R���G����h��q�I����^��U-��T��*Z��7���r�e�c3��L�U�
*��a[�s��&�J�(J7V����T�����i!������0������|��4�ĮKD����J�|/�*�P�o����h����z-*��d�֒�N��y��#n�
3$��܃u�:��c��N��lr��[ �����M�� ��`8�ۏY���,�؃�+ӹ��t�0����V2�ZfM���qʻĲ4K���9\�tW!��u������n��-Kt��ڠG^]��M���zo\�޺q��nNxƌy7Y!V�l�R^<eڭ$��${���.D�2H�̛�]ͺEj���lK�����f�SoA�+2�4>�V��QV0���ള���J����7S�u�3m�Σ�Q(N/�7��&��t���ϰ�j:��tM�o�����{j��ut�A�׎�H�\տ���cT0��u�KA h��{v��,6�d�R۱HVVGJe���6�������]ц�d1�H�jﷳ[�g�Ȕ݈ú%��]���z�t����^ڏ�EM���Z�(n�%��/�mPQ�����T��B*9�I�۴L���V'@m\v�b��VҢ,KY7�6�!VWc��+v��F�=ʳ+U�� WX��'K��݋�醷#�n��'n��,�v��g#ru�o`�e%�teL�1�s-�X�#���(�)�(x�I���b����R��E�Db�`�h�"�"��Kl��E�c���QVFK[AT-�iUX��A��Q ��ڶ�(-Kmm�h�ĴK*�EU���ŶԨ�R��F�m+A+Z���*���%�`����(�V�����KQJ�jX�V���`��UZ-�R��J�TQ�X,��Z�R�QQ�eAmiTUUdKk���ZR�����J-�cZ�kE�
��j��V��m��"�j��D�1��!64.4�Li�&�60E��1�H�D��,��-eAdcl�J�Bңm*UV
	l
5mcVTm%b� ���ZXԲ%�ZP����J[k[V�Ԩ�DV+iJ��J��Te�e
��TTm�RҨ",�Z1����[j�+m*��ѫ-�Q��F1+(,UD�B��VT�E--��*�)lT�Tb�ib��Z�X�X�E�QB��V�eJ[*Ŷ�T�e��m4����aMOO]{��y�]Jgl9f��sz�H�k2=Zmt�qFgw_LYHSH仧:�B����)-ܦ�zm�p����J��	�/:�*�ݑ��l��^Yn�v�|�rb6�5��M�����#��L~�Zi+�F��O�>=�����le���w^�snl��#�YWܜ�/�G9�����x�eі��l�&�ı�󋄯�ԶK��h	���xfӍ�"�W����h^��r�����ǫ9��Y��"01�nq剝�62pȷyz&�dV@��׺;���CFʦ9<yN%�=:=�,d�"��9�
ժͷW}�ej�z�ܺ7�gZ��$���!T�չ^�5o��9�3+�+�N^E�&�����L�u�z�6}�,�j|���Mn��9��4�o���1FVbAM��Ub�r�E��/&�֬v�;�+����e����+P����B;���H��(9V&��E��=�~�j�!E��#����I�5�� r�L.wi�]#t�4�^iT����2�qgm�r�v�X�W���t�� #��n	,V����������K�%q�V52�nkW|1k`<�T���.:RxQAVN٫�V�Zw��a���[���[{�"f�.ߖr)B���UE�Em-��M�Y��s��DDe�`���5t�1Q=�����k��n�(o�]v�R��lWA���A/5):�c�"�K�u5�����i���-��z	Y�
c���CbUrU�Rt�d۶��u��Wu��n+j��E$B�'���Ӥb]��81]�h0m�1f�mQ�	�W�Wd�=-I�;�hO_�Ab�J�kippe��R��@ˉ��N����(�o�S��;�����������6��8�R�!&ULk�I�\����3U�{X,%oe�=%X��$���*C��D.A�Qb9�t�W�� �;���7�L!�,��y�n��\v��&$pB=���STu؈����:�j��o2c&�HCF�3a��7}�r���穎F�҉�j�зqM72#rC��j\��Zi7(��[Ա���a�<D�]0�k��Ar���Owj�A�H��v�aͮR�D��Z������Ky���Ѹ.�7�g<D���}Aзo]q�Z#h�j�xRL��[S��'S�U�ɡ���Bu�Xy�w+�Ye�nÅ6����Q��^�s�ګ��}qR-����ht�����i=�Q��k�MSi�!��^mzn�mȫzUd@��!��V��3�R=�c���;�端�_^��C��y:�\	XE=�j	��6��e;Q�-�
j�VZ̗˖ڤ�m�]���oX�V�w
I\�	_A�֌��^.k�αԧ��>|���8��+GWNX�N�g�zM�i�1	1���1G���������f�L��9/'ui��Ÿ�x�{9� ^���d_Uo�x^'An������8�ma��'r�B0ql�����_Y�Æ�x��<.hNёS�vu��}MHY��ʷA��Z+i���v��I�C��"�T��P���ȍ��f�w�͍=a��������ڊb��i��Rd!���bp���Wb����S7Vpr�.z�*�O:�n�8<�^������gL 7��sL�w;:���C�ks���O���<4�&m�6�p�f�xu�9ݻ��(ʷݺ�I��V�U�H9�Gk#qjMQ6�g�J�>��.���S��nJ&�Š,�΂�>�h���p.�����VR��^�Uv
|�z8'v�{+�״�����b'���k���W�n"�Gh�����o�*.$��~^m�.x7=j���=.5�O�2�[mOt��	�!�fi�B��Y�b{Ր>f�����B�۰�X3�AUD���a��:��fjܚ9�nFB8��{Փ�bu�F���zNQ0s=^��N�!�>s�A��8Ud\�lH���LAE��a��잫͉m5�0f����(��AN�ӭ����Y��C��i���cLDOm�Ƹt��}ϲ���+٢'T{�3�W�����Z�X��7�v��1W�E���6;=��^�Ko˷h��_�uW��ͫ���\G���A�WʃS�"���uy�T����u%��r�'�Lk�0���WV=hT+���^�A�1�Ek���֩�C��N���LӬ	Z��(�����xa�����3���;-��,�_@tXv뺅5י��rծZc�sL�j�qgv\fa,
�ܶeM=��t�1�Í�s&c
TG��G̀��0{�${wp���a�a%��
�h�`OX2-����i�]�E���>�����<���V�ra;*��X���j/E$"z����>l]�sqm��	�5;�R�[�^{�2ӡj���Dг���!_�ٴ�Ջp1^��V�k�I��ݭ�J�%�aW�2'Խ���;������Gs-�"�	ׄ�^�~mM����v�} �:�&"�!4��c�5��')��v�b%W-0û�����&=o$cW�e:�/�YmZ��הeX�[�kHK�v������s�������s���ȑ���$ֺ��E��sZ_(Bg�f�?W2o���ߙG;'�;HD��6������Q�7��SK�C�Cf=K�q6f��D�7+�u�Fڝ�R�4�^ū`�%���ԡ	�LO'[����׋ݢ�e)طf�ma��ɽ���(٬����ޣr�^e���i�2qScw{1e`Ɗ�_ʨ"�AgO��G92k�F��_v�V�Cpɦ�$W�f>糧.j���{��VϖwW3�u"*'�� 4�8�J�<��v�ׇ�ӵ,V@y�xu�X�I����gh��5'�����uj�����1|2��%1Z�+ݶ�kڶX�m��F�{rL)>�l��;5��}쎑�<��)IU&�l�FVUїәN2��tr�)36��~��G�6�U�
�e��(>�z:�Jb�ي�8]��7��ʣ�[Ҳ�Gr�C頫�B��B�"E���K���NM�p���Bn��\��B�w,&����e��_B�V'�ڮ��Z��U�Uw`L�ڌ))�M�*�>�����ӊS�
�J�I�]IX����3�֗m�V�A�֨^�s���zF7�c�ݱ]	y�*��S�d]�ZBy��η�82\�9꽺���Z�	͐�7a���V�t�n�w�$V��5S4*먎8Y���!Xtb5���Ʋ�iP��6[c�ݓ�b*q�Y�p�3:�6��=�q؝7
�a1�OF��Sf��=;$�̺n�I��ALY�zY�B�i�yؖC�#��b;��9�c=���힔���Q��u;^�Mڽ�K�=tt���:���687#��9��������{,w1�9P+K�e���:Mu��^=�" �co��l���؆���\�������~��NZ�:�u��t����]��e�J>37�K�3�Pn@�����(����_��/-�G�v�{����ɛ��wT�/�B�����$&0���DOQcsiR�V�����3]m�Bi_w[��\m��2.�۔.u�=LH�c�]!��>B)%��Z����;ۺ�Y+��P�붜׮p��E���V��*c�^�"#a�w��
J���!2�k���A���U�"��+^ 򆠡�j6�DZ.�^�	�y�h�W���O�9cv��.�m�E�T�E�i�q+ۄB묒2q���s��u@��૓S�>[j�b���6��\���\�Y�<t�F+Q]����	c
^�Jѝ��yzPS���@�	Ճ��"�׫3�!���
�b-�O��=��H}���Z�����Ե���ċ�ܯ�k���^��׫ٸPDa���Z��_ݠ��{5~:�W�A��)Ɋ��+r��o �8d��sz��ʓa�.ƙKU���s5ݔt$QuwU�W�Zq=��yC�jNgx0bJ�	٪fѓX
�`Ku��+�(�YV��oW&�-�X1��j���l9�ʦ���z9��ӫ3�,�o(	����u'�pw+�pg5S�*���1��[U��Yu���a3��fl�]�������H��hf�Z.nvf5h��K���A�q��:bU�WsӐ��X¼z'ԙ
���v' 3	���ޭu#�_>j� � ��+��c_&"B��Y��+�rT�8�7�Ա{�����{�v��a�o"qZ��%��,5C:X���.^��A�}�ٷ����`Lչ�N�Y�������a���&,u�=���x�U��#����Svz*��W��R�_Q]���ܕ��yZ{T13�E�v�%q��L����|���A_j>^�
�f�ۭ�0���\ͮ�OʰOK�<�,�W�ݠXͥ;�i֌�(�*�$֙ɖ�?om�� K�M;u�m1�Om]�����g�.��IJ0�uҝ�l^�۬ˉ�Ѯݾu5�)�U������s���H�깍���(�mrFꐨ�j/U%E:��;��Kqb�0��"VwWr6����gl��P���}�#��qrJ�����}�^ʞ;�:=��'�O��c���Y�b4V�{3Ƕ��Xxf�;d?7ǰ�k+g�ٝ\��R��ٷn:���NP�7w:RKy����nj�{�d����[�ֹ_��������K푋:h�o'��.��J��[T{���lSX"}I6����­Z�����y��{�n��<��a�Q\��S�/��E���g���T��\S���t٠���H�h����ЅMb�"X��f�9]��Ә�*u�G6�FĹ���l#&*�R��X�{4��2a)7(�~�Ӯ¯q�n�⩀PnA,wD�$�J37��O��w�\7�Ž2���/9B'#Tn��c���	�Q`���8V�
/�� <Ƣ�;�}��.���o˫���;Wt����ܪ�\ע�ptMVf����r�5��R�׼9&�C�v:z򝊰�ꇐ	�Xn�� ��E�&�fN˹z���V]_^�)�WS���Nr��j��u�L��=5<o�.�*����;9<"n�f�EB�*D�;�h��]�,�x�v�%���A*�w.ɗճ��m+�՝��nMlK�,�9�졚��<�IV�71
p�Y��{�:��p��خfV�����8,���*N�3�j��æ��A��^�ɦ�N�@��.�u��x��|�������3Pã��?g�+�~+<r�7]�Ct��|��],�^��z�MXh�q!v+"��#��� x��z�@j. >�8�`s��2�kJ���2�k'y��ra<�t��#=��}X898�G-̑@57;e��(���E��L��|y�S�5J�����;�fU��oL�ŝ��+}��4h֭�7��|���4-�i�sW�V���`۽��������c��J��9�ehu�K����$�ɩÁR��$�+ۼX4w�d��~j���\A��T�b]W�#r"����c�P�p
-���[�\R&��ࢮ9@j��l6��넕CTt�R�˜����ҋ}ʤ��1�E*����WO{/3��n��X���ST�9[�A+n3w��F�Y��Z[�=sR�}�Au�������ܭS�(E�q�s���[�S�D�xS0=�5ЁT_\Lq��7x�N�]��W�<�zr]�, �4���/2q;����jG�r]��e�`�OTCsӕ���mqo[�K`8���46�;�m����*�d����F����n�5Y���|�7�8u�'�_ҭ;�YX*��3^��Z�xF٫�0�`�,&�t�@d�ixU<{Hn�0���]��%*��,VG0�N枳k(s�h�;�0@ˮY�w8r�o9�#�	�T��b󵌢a�G��F�V��$��M�ɻ�����8�v/ ޼zM8gi���Ǘ�a��!U�{��y\�Z�`4 �]b(�e>�,q��	ʸQ���	^�|�A��wuG��{71�2�/M���%��L��fu���`v�p����73f�mtj[%\X ͔seB�"#f��w����+��x%���[���om��b�ʦ��)�,y�ǎڎݠ��A��x�ܒ�M{������k4�턖n2��Ye��.j�rQ9(���i�ȉf��W��R�U�VtT[M�	�H�Ŏ�ʝ�5i�e��(#��H*Σ�,��XݼU�E��,�B٬�_�,���OP1����%˾�zT �Z
�%u۽�D�е��
����:��ÜЩM�g9�wV������E���NN��*��F�'��؜�\ٶ��ۦ���s�m���ʴH�4�ol��6���_���o.�@�u���UK���]��
��1�\Y-S	nrT�@�il�7`�xT�ϮQ�I���*|*m�M�gT��s30�d�z�+e��ɏ�ܕs��R�4�d�]gOW��D�E���+����[.�Z�c����TƗZK�[�xlp�/�4�PV�=���P\*��z[4U��Xg��ʤ�Ҩ�s.�4h���Z�9,k�@����n
\Gs�*���WI��RGZީ5W���:�ܻ[i�܄6�r��"��Q��W��(h &C���O	�ܵ�fGw7��v<���鑪ܮv�ͭH�fqg����e�Y��ZbL��f52Y&d䤮��wv�ꕤ2�^eJ���5�-��v������3s�YWI����2�RZ�*�Dp���u�dȘ��bvS��l��^����� �*x)u�
t���Zv��H��"�tBuoЫZ�EE�L�P�X�q��_²s�{1R@��jm�Pݒ�t��r��k���e��g\�$mU�մ*��J�M0����o��u��x�V)̲(�b��	�pJ���tKv��kjӕ�5�+J�2�����I�֠0ie�IٌK��x�l�*�:YwOχR�Z]w�c�R�Q�.�a���]���\�AJ���� �#�Z�؜�Ma-�շkI<�Z�D�G/�N�]���>���2m�mE�X���*(��6�A��*%�U���-Z*���؋�m�F��Ub"(�#mDTTjQIR�b(������Q�Q�h ֊*���-��Q��
�%)b�V��%h[((�1�EH��EdAV1X"(�[U�(�F�EkTE��Ȃ�[UPUb�ʔ�DQU�+A��EQUA��(��1�Z�Uª�Fڨ���X�+�KB�$QkYD�U
�[UF1E�(�b֢�E�D�V��""$Q+D��"�ԫ�E�TUFT�jU����`���,U���Z�A��������VV�X�P�� �"���Z
��֪��Jі�U",b+dTE���+iEU��
��-��EPQb*���Eb�*�(�X"�*��UDETQ(������(,Kmh"-j�PDV"���+R��� �	:Efn)���j��T'j�+�40�.�8�7B�}�bƷE��Y�xw���:��2�AuG�C�i���h�9�[��B�xŭ��G]m=c��<~:t�wZuE�ҍs�u�� ל3lEs�3��w��sB�9��v�}�6U�����]�*���J�xy�xu�Ҽ��xfy��'}����5� �*YB�'�NV�lI2�DE�6�`+�2Y{�E�P�VJ1�U�\ɉ�����m*S׻%���K��,���vb �^����Ϩ'�q�,iI�Y�q����tg�
,ht�3u ���P��6�>�Z��HE�{ܑpI�9����p{P�B,F|�͛sh��\�H�퍪{+�
�!��z�vY�"�C�={x:�Y�cKJ��xl��4:۱W�G�:	To�
v����|KâQ?-=0g�E;��1���*���n�,�3QeT�O��;�PY��x�뢪U��]#�Z+O�N�N���{������*�-��T���+EK]�N�p?5>
�{0o�Q.(+��V��E����-OZ���+�0m>p��=��z��� �X�P��������]_nL��R�[GА�21Ua�fέ�֑n��1��խ�չ3:��\0n��k#`s��z�-.�I�P�U�l�f3ضp͂'̻�s&���`k���bi}�Fɻ�L�X��Wg&��:��n��Ō�|��co7+;[�V�綧e,��wZ+d�Dz����t7u�j1�b��V�e��q�.�a&TQ�8`DT�MܸU��52�t��P;�(ӍJ}T��j�����>'���|ԡ��\{�n�������r�qَ��$���8���g�5�3�1`.��cv�갺V�4������0w*�b��V�dr���Z�h�G�B�׃y�4�O|ϙ��Z�n��I���z���6zzE�����]��к�)�qU�\_z��]i�e<�LI���d{�\�����rt�u\R���Ȉ����\����+��N�Y�sY��97=�O357ٖS�ӗ)C8��IL(!�>Y���v��,��+�T��I?5W��xE�+c.L�CJu��Ti�.�����w �f�TR<Ñn,�a9�0���}�S89��r�<4w�Hp`q�lW��,LW�O�*25��F8c���M��C�;:E(͙���2:��r�;�P��4D��q,C+�:�w�k�K�z���嫍Af>�NRtsp��(w�7@޼tIe�q5��i�&I��<�����k�\:ac�A����:˚�=��]�z��I���v�e�zi�;�����\T�$g؆:���V��> .��n����������N9�j�v�sx,.�5��r�Ra�sz�E�yÛs6�VB���U��)�r��AN?/���1A�6��s��Y=��	�f�=ȥ��?X�x���Ld㾕�-1bt3�*-9�U#!�\:�K3�8�S3��D����(I�C��:앃%k$�-��)=v�Y��>!<��T�~ƺ�@lMJ~��t�ty��J/ Xv�I���Uïm'#M�x՟=S�W�Ex<����g1,�yG��BQ�,^�p*�:���*5��"��Vo��o�<�r�n�B�U$��0�뷘�YaW�=�ĸ?����bc^���݊�}�''��É���K������[.�����v\�0ZU�;�b}����Jx�I�Ǫ"p�@���:�zBsdK�j����t�_
���j�	�|GR���6/�3aT�]�72-�@�;8�u������Ux��W�ϵp���W3�(Aҩ��0�]�T��x�zx�j6�e����gB�~p�u���C��_��s��,D9�/%R���C.�R�kD�����Z=�.>}W<<��k�-01�K��ʭy#�WKЇIծ9����}��_T2�:o���+4�.�o�V�GnCsRe_,�
�+�r���q��Nr'};��P�(c�}���	)���8q ��rӮ=�*n,ot�2M�Ҍʪ�7��[.k�-����c�~3�Ѧ���Q��,��4�X!^K��iP��ٙE��s|�Rb{���q�j$�p:�h��Ju�����|=s^��?/b��.�DE6+��CeDD�]���e�Z`f�ث�^�{��/���Y8pC��,%8��(��ޏSP��uU��D2��t`�Tw�>f߂)d��`�j�w��z$�Nt�G1�p���D��ģe�Z��g�\�D��ʋ�s�,G�؈�s��9t���!&��y`!C~�̞wW���>��=�jBD�LE�d�w5���1F\�`s��8l���Vʗ
7���W�b5�=��D�1R:o�@��@��,�'�2F57;`�B��Y�N��jMe��,:꜋W"�U�U������c�>Y���S�̋{7%%�Ra�4��?_����Q���@��W�1>��:���ƽ�K������%^:RK)�������'r�in�7⻈��q���nm�	K8��S��*%W��Nd6�!c	o��/J�W�k^�*�/����{��ro�u�M	lb墍���S�)�jR����GlB�0^U�I���+Z��1�N��_w�n�J�4��=}����
�"��T�b]R�nDW�m���7��G]F�I�v�{�]���x�a�-�S�kF#>����cτ���B�$��f�"�o��+������HL���ɜ�r��!p��U�#a�΢���Q�e�7e����%P��kw�nj��yͬ� �n���r�N�C��5��^��ÛS��xg�{	FP6 �c}�ٳ��՝4�vzj��+`��ӞP4�殴���:G^*�����uL�d^�\�_6����T}�*�`���rYV_����ȣF��2���,��ei]�O5Z��{|�*,����E'P
�ʩXV�+x�)��B]G��|rχ�6�<o8y����N������7.�ʜ�5p�
��T�߃��ft�ʜ�A�¯|�� {�<�~>�efs��`��of˺���X(�.���@"�=8mFy�V�j�ob�
En;l���0�~[L�}F����[�<F�����+��(3Nt��*�A�:Ɋo�Q����R�ٙˉ]̜����V�ږ^iD^n�_�"C�2h?j������e{=��ډ�"}0�����*Z�w>N��@��{�&�ft���Rs;�TҌ��.��	X�U�;��yt��wv]��o|��cpn���ҙay�k>����d�]b��<��ʫHAUo���r��ө��Fp-qK9���?��\�n��	�<�U���P^5�-�4�G)�]�XT�]Zc#Zo���;:�b�N��s�3Ǭ��2�@�3�z+V��e|���B�ظ/�a�?z'�P͉W.���*����/6Uy��=K�(`��s�J����DC5՚��u8�]��Z�3=�c���8tPMP�N��n��`} ���ZU�7���^�؁�������!*+�ݤ�
�U�`1���-Ey)�'<�b��W�4[j����ٰu��Y�s$�1�)v,�XU�����6����� QY�C�(�1�<�PS<c���r�k�Fnv�*)vF�\`�O�r�+:�b�1Z0dQ^�򰫏~�x�u��g��pͅv��è%Af���25�R���F��]OW�Iz냍X�_?�tmY�JԵ�k�ǫ����;ƯfdXnh��(P�kJ�{B�+���KW�<���~�v�	^ټ}C�V�V)��	b�6��ճ�A+�z�Z��]�uf�I༇U>����m��
Gt�7�y�eg֩��`��$��;a�\e�W;�'s��#[.�n.�Y�|1����E�ݴ��e�@V�p�R�^r>߲N�+;��o�鲳�Z���V̗/ϫ��Nf�)Lt�}^�Q��^�����p���y[:`�ʋ�\2*(Ƅ�0�"�Ψ*4Һw��K֜�:u9�f�T�^�"�S����NS���E��	b�+�G��c��0���n��K-ψJ�+"������L���	uYcM���'#��ɳX��v�ܓDH��:
+����nT�p�x`Τ�j������|������b�_�e���ϱB��[��{[�8�ddu�]gB9�����_�S
�Z)��;Ҵ���R4�,��gy �g�S�ӳ�P�J�Nv���o�� {�B��S�"�ʈ�J�V�<����<ljՁUX�d�}�BǷ���
���X�{�L5Eiq�8R�5�o�E��X�βë�*��=�������y+Ę��w	�ɜqo��q���q"�<��
�<}��՟
�Exs���/ȅV-qfe��	��|��g�gK��h>.������ؘ�[�D�v*�[ρ��S\fz��/�\Wy;6t�i,�:�N,��N.��G.9W���N��I��
֪�ԍ�VP}�zM���f���ck�:�V���b��	���'fyj�n!#�7���+� ���1�u��o36�}�-ڮī]u�mbD���$̭��u�+�G��۝{�T��k�+�_]��5�f��	Ꮈ׹��+W�2U���t�^���j~-�`����D�\�y:F爢�@TV��jF	��U�+�Kq^��,۬����ϻ�7T�v[>�'+c�+�\���Dd(=(ֹL#��S�`�{V/��s����[Й��y�qJ;�q
�mi�����ŅN��b ���%�>��ddq��u
Mf^(�B���0�S7nu��ŕQ�]�^�>�N�김x��A���L���ݫ�~�bn��aS6KZ�"�N�f8�v���7�h	�il�B���E�;KVc��o^�

�pyV�@9��f7>åTm�e������
r�t��g�K�}m1�ِ-�еH�(O*��^�b'j2G��W6vہdAN����fLj�\��V��,tO��W�@M���R����a��D9�N�`]ѭⅬ�ކ��ܻS��EN�G̹�=�K�{�,@��ǻ<�u�禫K�ʫ��L�g��Y�`𹤁��$�kX���2q��d,��wWj�վ�]��Xm�Cpn�| �,޸�i �&EҦsg'n�ؗoTqv�^�@�:6L$I;O;�uQ�%F�wnb����}R닶I܎�2��.��g�4�f��tɁ�;�z{����f�:8��&���<*U�Cޡ>�!�#˘w5��@w1Fh9;��}Cz|!�u�ɽCx���n��U1���:lu�;(^�����Śq�U{����}`�-*�rw{o�+o� �cƬ�ت;+���	� 1�ڪ�ja��V:���O���ouc]D��/{SU����}�>�f.x�t-�%Y�<5Iq����볤A����<�tX'�� ��f	��u����}�FߥаEyB7"-l���$���q1�&1�V�_s�3ڰ(˄ka��+��U<va�1q�%�6�+DҸ Pjl]9ݝ�	cL�3�r�]\_A��iH�j�S�cU��-�2����t	ڷL�<
)�F�M����W8�q�G�I)Ӡ��3w�#uT�Q���:�_��s7�]PPz٩��V��x�Mu��,9�Lܾ���dP#6
�M9�t��b�N���Q�{^��:\鞑}��������jx�k�]*���^Kj��l�%�<y��eY�/�4��ުژ�#H���R��;kJV+�<m$=쭩�5�vO�P�:C.o{���Ξ{�M��%��9�q�nf��7;�P�L�YV4����K�x:یA(�x�:�fn��ׁ���-���s���q(��<�ms�(R�Y���Hmu*_'�����^%~��L���)*�U���=�p
ٍ�"��n"��
�\=����݊�Ŏ��Gsu�w��QȆr�0N�2P3כQx�=jY�[�a챜�$sg�
} ֵ�b&TtQG<�W�by���l�08`����SN�FN�8mF��\��%��s�\�9U��pbq֙5���L�E��d�6���D���T���y��	�l�|�ܞ�y"�gW=�6:̢ۨ<���_Z�(?�s�zX��⁑�`�\�9s�1uB�8�۰�O��u�Ǩ|���V:��׬�����O�ȴ���O�[�huφ��}�9����O5l��ܭ���9����V�Ѱ�V�s�iך��#���z2탼��{$������0�t�[eױW�E��P�M
z�e
U�$�:aV��vmEݤ��o)�l(��&ΞjqI�i��^n��g�H&.��*˛���١�A�:Zڮ�;�����D�:i�`tY�X�;�3:���]Pw0ϧ��xxI�$�	'�$�	'���$���$��$�	'��$ I?���$��$�	'��IO��$ I?���$��$�	' IKH@�x@�$����$��$�	'��$ I?�	!I��IO�$ I?@�$��1AY&SYDG;E�)ـ`P��3'� bG[�{ٵm����͚�Ue���Z��LZ�m�b��*33jSAFj��Mh�mU��km��!���mf����B�TԪ��h�M��5�f�6�jX��bmg�H%ٍm�6լ�m�j�i�-��jeXڛ�kv���f���٭L7��l�^����[6�l���[YmRi4��Z�6���e�bf�LV�M�3a6�F-)6%jm���U��m�)�[VMT����m6a%XU�F�Xdh��ZJ�V�R��jm�T�(�l�[wqG6�l�Q��g   ]�}���֧V۽��,�Z݊n�v���U�]��7�v��gw] �c���Zu�:탳Zn���ʶ�Fc�n��u�֫����Κ�6[���Bi�-�l5�ihĪ O�  wW�O�5M�����ѥ�WA�n���iջ�{�۸��ӝ[�t6��gWx��Us-��g�����.��v�{�I�]��Q�h���oZ��iN�µ���mM�� ���o�  G�C�m0f��(]�)�>{ޞ��۷wkםHV޶���;�{��j�u�^z֤m|h� tQF�Ѻ(  ��{������th��p�( ���Z����kS�i�)K� � �  @m�Eth �v�( �5}��_I�+�J;d�wkf5�'][E671���-*&�z;���FG6�zq^����ڬѥlӻ�6T�)%�  <�H'��豨���y�^�T�"]zĹ�k��#Rw]�g]k�.��[�GX��gz���V=��M(a��"������U6��	���ڤ���  f�o��6�����כu�V�V�U��U�'����J蜖��n�w+G{]�իZ;ק�vkj�J�����!��,�v�iӺ�[N��kݺ�d�UT��   s��g��C6Ǒ�k�U�t�=���v��=��]���:��V��'v�9� V���=
��#����r����޽���4;rk��T�M����m�kLI!�f��6�I5�  <��ww]�v�}8��l�Z�s�{[�T��j-��ۻ���n�s��vWK7s�-{޻�ѫW3�+v����[wv���ݷZ�����s��C�ܴ�9�4�,�[Ml�L@�5�   �v�o�R�v�w{�ks;<{Ы��h�:^׏R�)�\�9�Kj�v��<� Ҩ9޷����=�p�5����x���l��{qʗ�;�V��b���ڳ���ل�[f�   �x�o[\�eV�����ݝ:����/Ez*]�{Ek]��gI�]WN���v7]4�c%��^�t���ק������y"�MM�=�U�w�|E?�*�� �O�bJR�4  5OdĕTdz@ �JTS@�S�4�کT� �J��R� G�~?O���H��?��
-�����/�J�-�������O��.~�w_�H@�^����	!I�B		�H@��	!I��ID� ^�����q���s���4����u�wkp�H�az1`�x�i��ZL)a���{v�@�[#���T�M+��b����_\8�V�.`�]���2e��(���E[���n�֏^C DQ�صe��.��;����Ș��Lܬ�V\�	�CE��lR����K���!�����	���Ö�7��wP�fh4I�Tt�3W�Uܹ6�m�Ǚk7i��1Ftь���I���Z�f�j���$E�NJ��!��Zx��$��Rz{/	�G �Zdb��0B���S��K`�Z��5u�$GF�n�D�����?l�8��*�'uU�  ��5�U],������d�[�S��t������m�-rG�����71n�dq�cpV7#*-ûU�Ygd)9�;R˥D�V�O1�!�9�yXۣ�÷�	탸����/H�*ډ�Z�͹`E�]�b�|�T�w���-
B؂��D���u��ZHM���:�qLo@� $2-�#�Eu0�	9����-ӵcqVab+�J�s>& ��oj%Zޙ��טs�l�jC������XɃ�Y	�J�[T),`�2����oc$)B�1�Y��[o_m�fL��μ��K�ujʞc��;�MY�W7Nci�_bj��*hX$�n)���v�u�����Xjێ1��wLhR&�];i�l�U �c��+�Z�1��\�c9�1\�UΨ��{�P�6����a�l�F`�X�h񱖊��Hh[�!���qN�{���
!i���n���Y2j��}� "���&9�@$�g(�Y���k�J:����H�8N!bK��Ʋ�kh�!���n�ԎɃ.e�Z`�&*�o.a�Qr�6�b�ymB�ge=уDQ�y+ ���f6f��"t0�⅕�Am ���Ln�V��)R�g#�B�j�b�F���^@쉦�v*�I�k"%�i^�͌;fN�ʇ�2��5�q�԰�@0��s ��;B�b�D��VMY׆�!�1#�����1��і�n�ū�4B���N���LKs2�����iH>�ɨ��3o\,��hq^�h�[0�m[�ՎXe��J�1��	HϢ�٢��R@M���q8E\��HK.Ù�h�!_]��V����N8�r2UiDQB�����'����T=Nz2��[æ��qeb�{r�0p�e����ViVآ)�f�c�'3Jp���94BL��B�w��1`��:N�����q�S*��A�ks�<}��b��ꮌ�r����_�Ɯ����$�ι*��{:af։����^�H�����&M��F*̃v�@A��z�e�At����b�ֽ��ٱ[���x�3g�NQ١��GuC&���ÐL���.��UQ�p�^6e8%\���cp�����su�w7�ːVa�ic�]hЊ�4Mn��2Zn���zu�5��;�Қý��k܄�L�t�Ѧ�:
�"��`j�4�Tq��Ϲ}��q�ū�6E~�%
��JP�8 ��5�G6`��	l
�[M���b�]�l�Ln�-P�����MÚ�#�%��rHe`[��E�j	��&h��؍���E��"#kgrq��h5��Gl�kzH�`�Bđ�v�e5Rg>R;%PEL�y�'(m��Ͷi�]�'	�q[r�748��Ø%f�
���C0V"�:viZ�J" Mj9�/Ŝ,�U=^N�9�x�ڝ[�����̉��|q�kLc~<�z8�=��xG� W	�wi����gT$���	g�M��|2g��tH�%C�wu42���2����k2d��썦����2:P���@b8f�xuϛF�2�`וl��.)�VɆ������j0�� �iX��R�W��m��q��L���Z���)���Mŷvj��a��y��N.�3��3Le�ZN�1��M��M#R�[B�&t�Q��s��js���R��gE����P��9��c&3��*5����ȲG�9��az����A�M�k��Oq4P+u��.�,U�7]�;11-�G@�ç;��h���0m������Q$�& �=�\1\�����m�-ӧE�ޡ�
�c��H�q�3�L�F/�c�����Q�Te� �- -6�8~�4@�|��[��hr��bR2�%ّ[o�i�a1��Pu�s������@à��쿠N��m\�0��9Xu�TC�HĢ�k.�X�G��:�n]��ut�*�ZQ����[I�<D�ިnv(�'
ɭ�f�:e���5��6���xg1R�}ȑ�7�F!��ԫc�d;�����b�(r%��9�v��Q��ެ<��N�D��&���Ⅺ 3�͐�4.��孕#���J���3�EŶ�#�M��Q��EF����K3Ul�u��8;����pڻ�����>K���T�ݘe(�[l�k�J��]��ҋ�uzd�\������iT
ٹ@eZX�
�U�zJ0f����LBc���I��u2�,����i�0V�bU�C]a�U��q����蹸�1�r�VtȲG���݃q�s62�h�^���4� :�U��.\ƫ$�i��%T�Յ<�A݇(9�Jak4[:���[���Ĳ�0����z�֑�c2�\y�%wY�`zSP�U�Jm�ar�դ�(���ͬ֩ˎL�1����HT�A9a3��-AF�dI�aխʽ5sLY���LM�Cb��0f���CW[�P�t8(�7)(ɬQ�	�Q��I�
�	0dړJԮs�M��p��X ��#Y��N�X�ycX�N'������"�j�޲�c���{��� ��E���,�KvPcN�2m�T��K�/CX�srh��kKB��bs��TXj�	X"%!�=ϑ��D�6��*m^Z/jc[�U����vnl���G59U*n��Z ���A)�,GH��C�}(llG���B��@��Uk@[܉��gQ�H��ac�y��xK���jY��*E3&*w%=� ���di�nK9��AۥV�fI�a��;��jU��yV٭�=j<�dYtU`�7T��!��5�:r�<vB�#6�3����T�YM�7���n:,�%&���f����Aˬv��^ȥ��<����AR�ۏ�ɇV�w�`ySp���n���M���z.�$��ږ�D{�WMR
�=(�&��ʛ�
@�sdwF�F;��*�m�6v،X�W�1ᔓ܉R1�6L��'H]��.�	�wll�3�I�OrkI���F�-u�$���{q#�$]���EG�#IM�U�ceM{���k1\�1���l+��:F�|�Q�lgB?9�����݂����X�O\A��nۅn��uw�V�a�!bɚavUj�qA��~<k��qK*�$Y?��Ŵ	���z�o8�B:NYP\�����L��a�A�T%U���DNU�²2�T�C1-X5F�^����ғ&ާ.�To	��V���7C\����"ʩ6���f���s��ɡ��|^r*ra�4�)�N�*>��8pb2T�.��ЭהbC7T����rô&=� r�1�i�	�#�Ie��	tٰ��n^��z���qsH�p��`������X�e���T�z��y�V�SjA���of�[�ݶB��
�����8�5��7��p<�gm�oT8�,��:W�\�Sr�E���iJ���4ɵ�L6�k6�5��A�w���C�jCwZ6))��8s$i�1�5��]j� ��嬕��V�ߣR�f�g���q"��
U���nGct�I��t��-l���J�eAh1be��)��e��cC*)w�gtSvehC�R���N����n�X*C����h�4��e��ѡ�
�M�%�;V���Hi�,��eb?�T���D�e�X�kİ�m�f�FK�YS9�RȒ�u�\t/�1u0�����̔	�\�Tu����_3���lP2r�-r�fL�LVTÐڗT�l�s���7�O�;1��7DI��ۭ�Y���f4HǴ�ȒuTg)4>hꐮ�"�,ek��ǈ�M��V����n-�m�t�p\�"Z�pǪ7 U�,��N�����O4: @EB�3�ʧ(	LA�ggi�v@;j�c��5�hq9�;)��.�0s�'ظ��Ε���R�����o
)�Ǳ�;�0bZ(B���h���ds]�RX�U)�kq`V*�����A9�LU����V���]��dWFBj��
�-h^����r�Owu�[��w��R���mSt���H�b��sBB<=Qwmz�'L�c9g\�p����>ʘ�n�V�zXݻ��ou��on�<��m���ܑ^$r���P��5���c.@��zlI�M"����h!�CrUսJ��c'f��QL�zT0ګ�zJ٨�Ja�=��)		n�'�z��q�[�o�!�Í�ʌR�[I�����ud �&��#�{�w�
�R�I�7c��N&��kl���m�m'L'����*k-n<��M��SSӮ�C��-$[�/ �	��S�cll�ڊ����ÛNl�l^�$i�q-OhAu7$��� <	���r������,����m*T�RPkʂ%�^c�hX�ҧH���2����*�~DRq��LE:*���p�>͝Yr�`��� ,�a�Nc��8h���ڐF���^Coq�ћ�m(�xU4�n\�4��s��C�¥չ9k�]�:����nl�h�Э�V�1�̧�8/6�����цc״�É���P�,bz��A�!���G��c&d�;0�{��q�E����%<nR8拰�^4#!��ʻz�ܓ�*�j�;�S>���j��+4<�Ay�09HHȃf#�weA�"�Un	hT�5�B*f��<EI���V�K-��@k�/����7�4c�l�AP�t��?).���z+6�Y��[\<�F��B���5�pAQ��v%�t��5rf��g,9b��"(X*��rK�IP��<�N+E��B��e�t�>6�-3]�a"Va�tOQ��h��V<b@�D�9��8:�I:��=٨`�^�w>��ĥ�W�X,աrM��^e�1u� ��a�bŷj4(����2Y��Xze�ú"�s2Jh�L�����:�����[I�oI^5u�*�X��`�E�dm* cU��F�̬-��l�&� �:̆�8��J�I\N��J۵	�f�T2=�i.d�dv�h����k�f���*	����eŢm����Cq�c������.��	wT5Yٻ����6�B����`3R��j��N�b�Ts-4�rKTÙ6�;GA4�i�-��ܷ��p�vХ�L�.��:�ô�IA4]m�:�m�C,��p�yB����B�dune]��Հ��6%��54�"����Z �ܻ�@Ҋ����xu���J!P�mdf��-�hֹw5��,��R!&֋z)�j(4���e+��:�q[���̘�7dŊٔ��(6��ԝ�zʸ�5��5�����C�	�*�P�φ���+���(:�.5kw��;��%lxknY;��:4p3jS.n�l��f���"ղ�S�:�*�>�	��RN�u�Ey����Oc��Jݷ(�&]Qɓ3H��t�o�w7K1��!料��Ġ舰��*M�q@�c�\�ZPmU���)c087�T7YԜ
n�u���^%%Z5�����H��rt��xݫ���Q��5��a�i������N؍f�֪U=������ZU(�̷�!tsD��))��,�+�Gr�ʝ�h-�Fѷ	Q-X�-�����QJ����Ő�d���-ֆ�![58M��1Ite��u.^j-ʁKN*d]�ˉ*�-�yZ��ne�a�Ȧ�XMnUú�����t�tc*�8D^���f��[�5e81��^3u-.`�8�x<�,	�>�8�Jt[6���6��2��s8��`ứ��K(�q7"	�F�*�1�LcT\{���I�gL��+z6�U��m���v�Gٮ������2�p�c̐Z�˰%eڣ�7+c2��:�cIPYȘݦ��2�L2u���t'��ŉ���O1�0ܲ�L-8#ܚ�l�BR���v�4���2���<�&��j�
���t��b�V9�AU� �Ӓ��&1;��`��(g1N_tA͡p$�!f2�y�`�-Ū^SdP�[�]Erbxh[���n�6d8 �#\
����Ws��Í�&�U�Y�
=�h�o]�@��4�m�-\�+
K>���s7mi愮�
���4�Y�T�OXK�HB6����5�5`)��(����z���ݼ���icW2��L^F��	d�R�V��,�vK,�έ��Jb�V���$���&�WRY��!���m�3.T9�����J�v�(�O^�R�X$�K�n��2���6eR�B�.�ik�n����X:���*H�֯�����s��z
�ގT2�B�rb��R��5":Z���z՚9X������֞���
BS�V�͢�2���]f����|���D{:h9(8.';��j����^aOk`�z&n!w���#,�9�t�����2�����7�h�9�H��ᚔ\I5Ǜ���J.���3)Dfj����F�M,�P�4�ݤ�l�̽R d/��:gFԗrf�fUv���%�|�:+��{����|v+�.Ie�k����{h�v�[�N�Pd�8*��μ��l�n[HwtmY��r�*���(��yZ���)ٳM�+yB��k.T�y	7J�sZ��������觜�}�r\X}CV�Y�N�;�/5��E���},��oww�񫖊����/���u����軰�F�U�۱���Sy������B��Cu�(�%�nf�=�q���-kOݣ��1��SÈ�{��yu��1;���e��0��݆�>$���,բ:�Z�.�q�mͻ�V�gN�̬�8����C+s���.Y	\^m�]4[�Z}3ëa�6�G���-�b'���h���1�6���r�T�k{�Y��fz�+�O2���J��og���L��c�ǴK�]�8f�Oa�����CDȇ�����O�9�n�������ف%>�E/�Ŝe��u_c��ޞ��7��uri݀ݼզʮ���=��tx���u^����m�Z�}����̳,��c�$�VNӬ���Y����T{��f�JC�l�/vu1T��	ua�.΍��u����s}'��L
e���=B=�&�,u��o$&�E$��c�cFV�c_
&Nx�5��r%�}s������-�b�$܃�������^�/�;�=�
x��#ۭ*�-Kq{���v\=�s1Ѣ���Q��.ߑ+��̻�U����V�+�O�*��-Jj�i�k��el��;´���4�A&��M��l �\�V��@qg��B:\��n̷l���4.wz��z#�&N��_v���O!76��8fo�Y�ϾZ�>[��W�&����U�Pu�.���H�����%u��RO����ل��1�U�I0��{Ed��Q���9��s�aao)_^/�,�;3���7b��V��G���vc6�����Ĺ���/��]�������6;�]�62�a:4�S2�s�x��S��wtA�*c8`ʥY��j��#X�O�yԬ:��o�It��e�6Y��|��~�}E�>9r��z��zX�/�Y.�5m0�����y�y�����X�\u�4Ǣl�u��Gif<�֝�2C�J� ��A���5��y��9�Ӹ�݇�=lI���U���vI�Շxu�����"��o7�Yk�:M!��0��.��,n��=�� �w:|��w�ލ��2����Y�2*O��Żq�ִ�+n�2�t��
��a4�<��V,~p�hf ��.��VADE�0,��1Ո���5)v�qoܤ�|�O8f��]Ng���aT�w�lw�����ܘqI`*,�y�ݭ��-#.��\`%�x�;�:��ª$fweԬ�:�7��m���7D�j=.wgJH��j@/J��Uw�֊v�����q���M��e`�hr��M�ɫMF�5���6x��f���Wj�}-j��š��iu.��磺�_�9���qr��+�y�`���s��m� 9��Uf1+}�%@���cp���jc�[�e ��.���tDo)��`ڌ\˰�m��ww/��;u�wN���Onk���\#���6�X �ɪ�q����澸ۆw6o1l���W4\��vien�V&N[o����^pI׋>*�&q��<��{+Qf�6�q�;M۽�huy�����Z��ݷ�:�2�>�Z;�	0�\V�cB�!g�����А��R�*\����TS��H�݁cFV>�M���q��9�����Z��6;�FS����e9v����4'eР���ɤ9	���2��pp2�l�v���t�s� Ӿ�;z1��b��}!����CsqK���	²��Jh
��ٯ�T���v@D�8����f�=���$7��B}�Za>�]��S�K�ҭ��S��x��|�:�R;�9��@k.K�v^�xض�[w�,�w�]���<�%�ORp�v=�{.h��[q��q|��J�(��Yoz��z�/*n00ǋ����8�����yo��Y|vc}ư����e|��j�{�>Қl���Q�sɸ�ޯ�����u[�l>���>��Y]:[�Z�hN���G9�V'��%|�[�nI�J�(����HQ;��1;뒷!�ƻ���>-�;�k��s:����a����-ݜ��g���<-\�MEs�]����.�G��r�`=�������yI�ù���ʏũ|�a�WR1����(���eΫ��}�g)V�*��tX�\zG	h+�2i8�b�S�4�� ]y�nJ�W7���o�cG�Þp�L���"�.�5�Y|��*F�;_k�����S3A
�5��)nfyK:s������:ףv��J�L�K2E��N��'.��/���\qnJ�Йq\�ۭD������d�N���6����w���ԃɿ`·���b�V�����s �^�h5�q��$��B�pD�ް��U�����p�/�
B��B;0��H��&�d�v5�l�mc���k���V��
��v�$���)�����h�p����na��(7�������}9���p�\�,��w;���[q�Ú2�ws{ګ�SY{Ŝ�.��#5�Y��iyv��5i��0^b�_s�k9
�9�=4�O�<�pXGIsE��{��~ѳ�뾶����>s�Nhi}�Je�4͍rEz�\xp84.�k޾ʗ��e�r�1]|v�[yE�0ΥG���$��!�Վ�y�=@�[�IU�rW����Y��g;h�duj�
�}\�;�0�a�v�X�	Ӓ�ѥ����0fMy��ڃ��a��4"�ܲ�=�.��u��O���x�����߶��am����CǦv��R��!���鮧�ɟ.!� �[R�.t��unk/���vR���,��l�Q�t�jWg^��jsq�,A@������
��Ձ'&��5��v�p�d��"3^���9�ذ�ypＥ�o1�yK�^dcFfA�NG�mb�r,+&�a��⯋{������<<�V�sٕ��Sc�3�Wc'k�|�6��,��4�w_[�@�覰U�=;�5�*�f��B&�N��������CX�S�,pBά��`ͻ�}YK ���[ң�8���$'rCE���D���%k�F}��A˭}�}��$�N���u�(6��nQ@�+�2�z�eC�0��	��bޫ���]�vs�Mo_,��ٜ� k׋�M��t]�7�޻�-Sj�bH �ځ�,4�(�|��ek�j��Eoe�3-��qa����f�CBđ��<���,��B���޾W�n�S�Mff��ZC���*�f�`�3��Q���2�~����_.��E�4f�ݷW��5��x3�S܊���g���}.����4�̬Ҙ����U?���:�O��aH�}�}�t�o	�]h.>�TAq��:��=�wB0���y��Rd�y1k����j=�E����()I)՗�<[P��{�uSY\�����1$`
˛E�#^M��1���+FX�-��T}�"��G��:��=ݼe�����x��rSs���'�J����q>�����9��0�3�q9�:�{���A��v%�Y����0��ԛu��AO{�V���k�������S@9%��GN�5��ܕ1N���D�.aS�%�6�0�~�wO���/�����O�%�Z3�aʴ����QŎDH��4��L�cn\�ӝ��!2�Hە���ݤǩ�����G��R{�V_��4��N�D��7���!�\�tN5��RL��e�Z�K�c��R�<�}U�*F���H��R۝r��s�M*/�!����r��ҥf�	]�֯�[�D�]�qk���>�Ye�E���|ؓ����r��R�� V,���Ř8��A�����1�J�vg:ʈ�d������(�N����<�@��j�s(�*I�׬LPAq9��.������zy�ܓ������l.��s��y�QS�BfzW��8)�������$�ɻ�r1�y�B�M�'�(�^�Ec���b��$�5�7=�
�7�O*��4�:��z�lb%�(r
K(C�J��۵{+��l�Q�
��[$�B�[X�PZt��N��{�׾���}�=2t�
�W^m�c^�����Ukϝ�9�U��I�f�t��\
�%�)�x;6l��{��c>x)
�:R�lր��\�k���;��Gm�_I^�9
74&�3܋�;'>P֨*��X�wW�=b�փ�OK�����w1x�ȝ~x����z�̞�����ۣ�纛���g��9I�51x����4ٲo6�l���b��YY�c��cp�扥Oi�k�K똎!9�.�cq�f��|��A��[yiM�z�5���tᬭp��ۑqGʙmn/�^SN��� ׻�K�B���2�b����h93N����]�L��:g������J�q���Y�-x�e�q���r�;�N&(��2?(�OW��g��5�����)j�`�B}ݱ�+�� �zDt���ꌉ4읕�e��(�;�48f�);���BMԮ�S���؎��B'��O�{dᔞ��'W���z��P&+����{Rov��[���c���<+�U[4�hܺzi�J�VW8�h9�_k���j�gV]s�{���LjY�/77�j"�G��5�]ɣ������,C�2ghҬ�}W(��NZ���m���90̣���(3�kʙ*_a��v0ʺda	���*�V3�፱�W��!;3�Z�7S��29H�'!�٘����AM��Sgf�כU'|��'��ŕv"\���ז�tI�|��v�3�zW�����������T���Gr�;��d����h��v�To4Y�h-o8�ROJ�9���0��m�]cWMg���Tar��eC������;���`��z��53����w�����t�o�gc��X��%ż�CYo	�����]�w�^�4���bdvT*�Lpd�5ۉ�G9uێ�#w-
�gs*}cl��K���Ql���ë�yk���N��}e5H�G
�69��-��K�\6n
U�þ��%S�w���T|�nԺ>�{��Q�W�������w�)��ͯ}0.!�_?cZ�'�Ƌr�N7Ft����nEg�5�Cuj�d���|��G�*�I�PN�4(�z�Y,��Y�#i����9����2��T��9_ۈi����
 %ra�Х�T�b=͕�����]И��Y����E;/�.���6^#�7=]��!���m8l��޸R"*�����juvW�.]����X�����\��_5�����l��.���~����	��`,�\`�L��N�,{*i�iOfצ��׺fe���E�t̈�̜
����N�]��oq�l���B�1�R/Ѝ�E�ܳ-�)8;Uln�ھ�7� ��n�fod�(ʩ��1�:��Z��e٣Iy�S�-B��W.J\x��-��^�@���2?@ ��Y�4~�������6Oq� ��=:U���7:�"�,�Z���H�E�����բ�a���hT��F���U�zR��!���k���M�b
��G}����_w=��-��N��<�
�_�wז���p�s^�qb�o�1B��=ma�t�Hň;pd�h����ͩ1L��F
&
�9�|����䕗�5)��5b(����齪.kʜwIN&��N�D�����h�y���5�pKW\c_L�y=K]'�#_��Ǧ����0���9u�m�A�^k��W�����+%HX̝0��d�ޕp3��P6�g�7B���<��L�?y'(��s�5�bq�.�\����nf��Ѧa�e:�n�cu ����K��x����\�C��fh����S�b�k^*)d�g*T��@��oF8m��z�Ż�����d${�&[�!
�)��G�N*L�����FO�X��&��U�:븎ڔS�ar���gE��M��a��n��"8�挥�C5p;P2����`�WUu�b���|+%gp�����먑���(�o/�v��}��y��)^�:�.%�J�.Z�7Svve��l�W]��9�b4��������8S��vk����}��7�c|�2���G[�6�͊�y/I�s�鼦r1�����l�8Kw�̇<�N��O7�`^hx��x�x;d�(����>���xWZ�0{ŏU�Wq����U�̚�����J�6쾳�I��m#kj��̏N��]�q��O��}������h5���T��*w;�t[Ƥ4��gg)�{�<�]ޣ��I�A�iɷQf����䮝qZ��5�v`}tpB��%c�"�ظ��75jӶ��1��yj�HWY�3�>���}���/L��xomZV*��M�.��3��ȣ�Ѯ�C�h:�rT�*Z֧��S���j���.�70m&v起9��s�J��=�Ȓ�UZ�45�3���䟳����C�4�>��z��Sd�c�2�hbѲ;��Cӳ��OS�6��ɹ�t-�}�u������$LU�%��t���?<����G�\�-)h����:#�%l�D[�OyW'|�\�V�r���Xf����W�9����k��SMY��}�����Z(�/:w	����WM0����v֯4�|k9ͼ�uƂ��V��1���9����G�N�D�:8u\�;�ʾU:��s{�1s�~��5�r�HH@$�	%�9o�N'�/�[�'��i'���1<0'����I�x����W}�:Hx1nq��Ca���P�:'C&���DF<t>�P��9a�[��&��V��`���C��IK�z//)X�f�����>�#)ض�)v��|®-�3މL�N˦��٘���K׺ �ig�	�+�9���\?^K�*��$}�GL	���Lؤ�u�������%H���}����'�>����;��ᓞ	�[����͵���PKYغB�*U��������b��/l��S��sv}������P�ou=��6Х*�XЖ�`�[��Y}�yvXs�γ�-�Np3��8��*�����B�uI�j}7K��o>�X>,��gR�{؅[WӦA���vvv�֊F*.�{ΐ�4$O�-\ �&Q�n!�ޛa�5ޡ��yf��v�����2�sd�wf���zf��=zf�rVŵ�/g���|�k��N;GO6��O��]v�f+$��O���K��j��M�Ӻ����Ř���T�ԼH�A�{�+���� �wt����sz�
��n2Z�x6q�3A�6z�\1{��c��u��
��J�i����6�kN�if
]+�]��3q�fD
}O�Њ�u �\���
�OHU����o���ڳ��Fg0(�Y�9dҀފ� �`�ŭ�!;�#�[�+���A�g��8�&��+��w^o;2R d}Z�$E:g`�M�J{�+�o����d�K|�o�P���䲕M���U�]pKdKR�{f�λkm=�)��Ǖx����?'���W�=ɫU�1Y�m��݌�րp�5��ΝD@�����=�;	Mր�����͵C��45�z���� ��kV�tK9�Mj�y)3���B�M��&��k�\��]��ܽو�#Iԏ2�m}�����K#�����ʷd}�5��W��u�|z���@��עf/z!���;�B[�g
����a��=�y,�یض�E*��ˀS�Q���zv��f�i1�3�E(h��;
�|�ƺkś��[n�೗��b�EF]\(q1�ei�=6����ӣF��ŧ����7�O}�5 ��q�Y������>!}}K�E�d�O�u��29.s�7G+��{��QD�S��W�O�:���-|�N�f�u+p���J)	ϭ�#�\@N��Ƃ-Ɖe�鯃%����IL��c��q� ��]�v�vj�������Y؆�%�+��:w�[Ͻ\�(­�Z����ql�ܻ�Y.b�׼UC�|�bo�<=[&�^��6�ԡ%�l����eG����Ƽ��.a���$�a�z��y�s��eӀR��W!�K�Ϋ�Tʚ{���+��W�1u��������GZni�G1[CM�NI��;�9F��G�<���,^Vu�@�;��fLn��x�j��g�Y�vi�ck2��y��~��l�˕-���b���������/�r�����{Jغt���W(��Ko��&9à�F�l���b�fLd7��I��\j���������Q}z����*|���0�ʞepг�T�nE��t�/]�j�J�F�`F�*q��宻$E#٬[��<c������K4�2nu9KBU�K�d�(:�Y�m�ka��J�T���Zx��- �<��x*��0@��k��}�#M����Ӱ_}g����߹�&gb�l��G�?�U(Y5nR5��;d�9�ŋ��Dc�fnf��=�k�;x��DՌ�i�PM䚙t�� D�����]�֨������t^ڐ[}(�tv�!�r#8��$����U|wV��3:Bpt�]��c,�ck��P�-Ʌ�Ԋ��D���h����D�|3;m9zW.SyD���G�4�'HB@�Ϧ�6Ǽﱟq��u�g�ͷٳ��$<(��U��ƹ��`"?c'��7ӫ;l��q�����Mo�j��m�h�.IvOA"�{���/d̡���H\X�o6&��aKUu"�1F��P���e�y}|������3����w�u�|�R�%X6�\��������v��X�:Џ����(���(�aGF����-����{8��z�K!��X����!1U��%3c�7B���LӺ����/0��h�r�;��>��n�	��4�"zslTJ����[�j`*E\{G�����9�n:3��M���饘8��n>9;��!'����AD�q�ްF�k���y�I������3��/.Q������/@\�qm�ȸ��[HZ�6d�6���Z��D��%%��-%n�h�v�e�n��Xv��in;�u�``v�;*u��Rg$o�s�����kNgwAj��2Po��]w�&<2��OM�$���s@fp`���LtK>�MFBS�y��?��ٙX�;�í�+ރ<' �Ώ^ǳ�'�}�E��7���f�	/�h2N玝_`E(wv��BV+c��i��ʔy��j����o;�W��� ��)۩�k�v�!��Μ� 9��\�pv,���7��N�fe��#�d%|N�^�f0���-�4`���FL2T��!���B�קH�`�ݟt�m�pΪ�[Q�9�b�D�#�.�$<�����j�=in��qѰ���],�^�����-1e�Q��u�v��Y��"8<��[n��`h1q��א�%��2燼�<�`Ŭ���4�W%ó�.:�޵��7;����w=����`~6ۯ������o-��yx�[���w�9#N{�k�|�����*嘔�w�w"i��i�J���\���%�:n
q�&[G�(F\�̶z�9֭������K$�7�FS��Z4��;���/&;��c"��o�����	���Bӫ�Ⴃ2u���j�M��x.�#�ݼ���u%�2���X�'��e�J���B�,��uLֱ��S�w��vu�lQ�ͼ�	Z�.�m�R�	ڄl%+X��+�tP�M/��t2���#	�k{�V\�Xc|�Z%����Yl��1|_H=�/�fr�=M�]�{2+���_��yMuy�G75�=8T;��{��9��K�қ�WAB�&v�� ��l�:����ZL�}l�>���v�K,V鳣����x�0�MH�p�k;�B�D���9xNԶۺ1��#y�!v��^��h�}W\���-��W͂M:��to�7o :�M!��+�X]8HK�'NHt}M�Х0��r�@T��+-��A�d�M�x[!�	�9�oa��]k(rW�p�.gY0���%�L��d��5���h��ݍR�ͩK��]\ ���-j��o��n��໕�Z�Be����)V������'��)��e+�{CG6���w�zgێ�����v���吶H�ȥ3k��tg�EP�bI��G'ò��ڱR����#�qw5{|�������)6�����2i�ޠ��u;"���+�I\��/$������lwr\��d���=�:�d��WqN>�:�|$���gIt]�3�6ﺞ�g���@��'9*^R]�d�-�w|�(��Q��b�V펔�'f�s/^s-<�Ѿ���p�xC����ڵ&	�*�>מ�)�V��,s�ۗ�h���G��^��-l��V���j���ΜV�Pz�����î�]֦����+����{Qv,X�Ѱ�sg��7G�D�����lί6_r�����x��;懒�9%��e��>Cy �k�2M�x1���i�#�65��-��Əd=��]�A{\��	;ƕ�a��vs ��!7�nx�DU����\^�"�E�x��1}�-�'�w�t��1�����
��xd]w'�a ��[xUrܚuwE4��sK�i�P3y2�����m��Q�t�����Y��{�{��Bh�Ns[�+�ՙpհ��<ػ�5�AkA�0
'�[��ܭ��LT���.�NQ����uӬP4�b6膆�����*ܽ�[W�=ku�/	�V�[�xv�8J��v���Fq|�?8 �nօ��HC̖_c.�(�˸����md����UDvs{yM��钍К80��'tΝ�(\R���l�n�΅�ߒ�3}�{����Q�-aoxn�0��b&�ݚwZ͑b}���:S4M�_>�+ �4��>��bvO�+�O�ͫ�"�o5| 0�2IYd�և�������B��Bgv5X��{�њ�9�@l;4����k�Yږ��X���W$�pڃǒ����ҝ!�C(q�{��g�m{��#�Ah�\Qd��$]Ap�Iݳk����իN�˔�����͌�+��3#���j]F����oC�d�SsQX��x��nv�U���oM7��geѻ��MQ��B�|�tK��2����Z�u�+]��"#��Ӏ�b�o��3Mxshb���t�n�-h�-t��Nh��i;9�����Z��l�6������rC.�:=1�ј�̖$U�WY����'��kq��2M������C�e���v�vTC�Ɍ7z�ѽ���wS$���-.<����"�p�yE%c%#6�e�@�������$݄��⿱_���g�Q����`3Q审�gT��e��7�OO�fs��shhu�e65C����>wv
̀!�����R�ͤ��d3���Ab�	����=U���qB��T���E��t���U7W]|����;��S��5ӸU���1��u]��`���!���"5V��Qǈ�▴;��zf�ǯ��-;8�R.������%�d:����b{cX���R��8U9�^w mN_�??�L�=����y�u�*��\�bZ��8�W���t.]5�o����:�d<7�}�%��ƨ�)�Aג�m�OG~�����X��������9pG���A�Wy�b�w
�R-QgR�g ;�5��)��U��͗Ժ��qO�ωΌ�kΠh: �����4�f
��Jd+�&���U+�"r�F�������B�B��wyӹEW�X{,����VL	㾓B�1��`N.��.�]ke$��@�����vWNXs���c�n��l䓥)J�;��r�o7Lz*�l�[� ���{K��)�x]���� �Cq���=	�fȕ�W�t�:Մ�̽G ���{wR����x��N�g��c���c�-��Ʊ�^мq��c宲!��/��]Hq��� .�e����yN�+����[�}��/�ˁm]���u]>ct�Đz�[k��_y\"���KԳu�桹�g�ik�>RV��Zv^WM��*g.��I	��\ z2�D�fp��D-Y��7�ݝ(�%;��*��6
*	3.�m������8�/^�jg���Q�Q"��qf�3-�lW�p�V�}�y'��F32r7uc���N��3w��"���w޷��Jܢ�э�y���~fh��8.cMde �
}�����ޠ:]iƎ�q�rT6n�R��!DE�=�fګR̐�u.�"z`��<�/3��#�5����>�=|�/_�t^U������e�ƹi��f1�{�9�;%5���׊�l���M�s{/�������]�v1=�Z�����Ky�yM���>9ܞ�W�O{�{	Yp�����aø�C�4�Ɩ���D�B���8�ֳ̽�-�'��T�hN�`;�Lk��t��=�FLV+0^ՙz�P!p�����m�#J���jt��)���=l��r<Ѵ���a�uN�D̏3���t��O\ɔ^'
�������;ZDy�WCg��x�y�-��x.�Tf,r�����`�0���X�Za�]+�%����Fhu:�ev���!S��ܓ.9�z戄�m��
}���۽{:ŮT f���K��۩i����)�3��r�# ��5�%��kreXvZi�AJ�T�O�R��c�%�y�zŮ<!��x�:&���pQ�n�S��@�n��F�w5�X	�^��2�o3���e�k�7���OZ6��7�J=�׽L��J��p��v!˺�W�G�<���h�v��ױ��B0v�D�7�)�`Νl�b�N���N#�^S�/�)�����(Lܤ��}�.�ܚ�v���Ӝ)�zK�H�o�֡fC�Wy��]�UN8L�&T<���'@P��U��乘!�X��{��H��_<�}_�4ۘt<3��O�O�1��5:ZY�#j�b�AŐ�ϭ�o/ �d�]������gY������e��À�H�.��YӳN�P�X�m^p\�Kw&c��q��J���2,Z�9Z�&�`a*�FJ���&F7QQn]9"F ;;حĳ�][�+�U�~��n�����W.�$k1��wº��~��n�5�����.-�X]�̬5ڌ�#�ָ��WT��m�e�N�`�S���!6M�uG/�.�͝Z6d'^���I�Dq|ͱ:˩��;��f�b���)�	1��7�+�;���eȹ+t�6h��N��ˬn�o�6�F�+�,�d`Or�W�и�W&�%*s�<]Ӹ���v�i�c��|%u��k�(��m^����R�K��>b���6�w=L�l����o�.?���j���Y�,��j>�����3�4h���=���{x���9v�B�v�J�A��������1b�\#+���~��e�-��5m��x?'�ut�M�ts�dٗ#\��U�{XIVbzr�����7{�&=A��l30F"���������̮c�GLgWS��yku�/	pZN�gr���Q����TL���̻�9�	���ƞ&s��~�2�&��H@�Y2�[����x���c�n��+B�4Ỵ�-�M�.z������۽�;�x�.=m��}���)i�� �[�4�8O,�Qk�+Y�d��36�ТpS7{/����W���10�V��!�-V�F�tQ
���{{t����R�R
�6��X4-����.��뢃v�:!�2�/�`��;�\/秣�E�)���������#ރ�����-���ʊ�|�ً�<�XE�����C"��}\x�x��qҩE#Z��>��p��Y�X�#�*L4���-tpQ�d&��vd�9�rV��ZGU�}�p�WV)N9��S>�7�(�jD�}u��=,>��ӌ<V��2��P���M�@ha��]�b���.jE{ھ����[<�����p��O0�_vo�*��,+��g��A��:���cjv� �j	��FŐ�DmK0S˳��ALPۘ���@l��J���40�h�4�utD�V���ܑ�e1Iִ�?��c��э�]D0�N��]�G�j״��<�[k�X�m��h�%I;��_m��'&i��ud�i5��C:*X���[�D��kl��Q��}`�X� <b=Q�3��ꦡCڻO�d�$PS�
r�@2��ͮ���w��oP�}i7A��G�!�Y��:Ռ��s)�{���pp�ȩ�U�ܮ_;=�{*�����N7�)c�Ů�fJ�&������bo[�t��燢��f7U����<|�x�sؑ����u�Q�����d\�l�%2�*(��|��n�Y�7�a����#
��^i��"ٓ�����}�C�L"-B���Q��AUE�TKe+iV
+R���*��Q+kU�a�EQb*#���+Z�Ub+*-���kR�cH��8q"�Q��Z"*��p)AX�m��*.�L5*V*��DEE�Eb�iFE�B��X�m�Ŭ0�B�b�[E��TX"��EL5b���([b1eK"+�l�Keb��b�2�j2��*�mh���PD�a[ZEQI�Rak�PX��&��#���*�L51J��PF ��)R�[aJYZ���-�iQT�)Z,�l��+Kb�QbԱ�ƵUm�DTAQ�"+(��ң(�b��V��Q���A�Q��V4�DDF*+"�
��cl�EbP���*����A��Ub���1��eB���`��HƵQFڨ��
V�PT���N�tg�×��*ݛ������C��7�9�Oq�g`��p�\�n	\���3`��Y��� ��HВ���ٓ���=FhE��'���;���<(��\�s'%�A)����Cx�lG�f_3�:,����W�/�#�7�{<�-#����CH+���oӛ�};	(e2���C��f� d��WO&�2~�ឥ�ʯ���%}sS�)w)k��x�w�^:��ͱ��4G�f�L�Ǒޜ��^��R�\^�����Cj��JSS�5��J��M����.f����@y�E�X����\py��ô�sʿe���,O7�8������²rF$�oZ�[�>�z.�|!'�a�]g��oH�" Ї��V�o~�^��p�,�̔��)����c*8����(Ǽ�����^қ�"�̿�S�)kü#�W���4�׷��~vl`�3�FKvu�ᣀf��]�2�m���4���8����əa�pOϼ�4�XU���>�}�[t���A�B#u^y�L;��_��.��n�X�piiF}�������ҝ�z��9�i��Ih�>Px�R��Th�dq�;O��Z=*��!��z�lU�	���|��Vm����\^Z�������qEGٍm,��}xkf'�r�#��.̺���!�Eb5�׺�͹5ϊod�B�������[9�w�o�L����:S�Zw��q���4�-��۽�}���SM-���5�X��#��w����Dlۈ.�� ��� i���}QC��s=�C˰-ܲ���($���)����mq%5�x������@1u޼~���mG�WJk�swV���P
�b�W�K0��%���)�`��ؼIN�u3ƺvt�v�[z���/�|�2v��L2�)m������>�ļ��:T�K� �S�BK���5�:�Е��B��ǵ��Cز�*��g�U��Ͻ:l��C*��6x
��^Һ�������|%� h���[� �OLT�^�pE{&�։�+���
��8��+\��NV���t�^��lmd�,�zR̮�+��s��xy�D�v�@����z>�;���WS}�!�Rn;�A���N�%�oƯ^�vr���lUb�ee5���Z�L	�{x�Y��;D�/�E>�*��R߶���v��K��*��lk�L�G��rL�z��"��`�9�N�pmqL�,�����]P�k ˗���zh.�(�+�
�f�yS9#�.���������!�iv�kܵ��B�=�f��Z�^�7� }���k�Y�!�Ke��xK^��G={/��}�G��݁�����i㖆d<�]�JH3����fG�n��cU}�01Ϋ��v�6�ߐ�[Z\5�>���;��WD�蓼CA�'�guh���*�ĹEU�v*����L~�M'n�g��xw*̖�Kw����őT]���	��'�w
����t.g�3��\ �j_
!�]g�p�fV-k��F'�蠥V��c˷j���ڽ��ս�/_����Q���)Џ+�!b��J6�*�0Z�~8Z��`�ǯ���3�z�JʫN�	��ݸsh�po���Y�ۂ�d5�N� i�5�+��{��sR���޻p'�-8 ��tTa-#z�V<ɜ�;�3�6���� ����a�\(�b���i(.�D�!"���D�S7r�����z'y��
��t�	3㎧�k�n��IS�E)wu3�H�VҊ,�4����ca�$=B
D��5��&�h����n�K���
�|s�Y�ݐ(T\��2�'-g����X/�M�m�m{�k�P}e�*U_��~jA��Z괖3픀���.���Y3{�E>�&����x�ߣ�NN<�l'��{ya�ܟk8���;��yg&&+�t���=��,1RKS���p�U�N��U� � ��RE��.`��ޓ�Q{�K���{�%3�b�Z|���Ͱ�{67OK�\Sy�i�6͖��y��̙b�6`���d�c�E�u�t��z���(gj#�/w�	�����)�����J�N�b-�	|��ᴼ�X��W���]�C*�xia�&�!���3c�T��rο�j����e�<��K"�C?.q�e�kp�5`�_�X��7z��6���Wh�LJ��}��t�7�6ehW��ȩ-�|4���X���ʑ4L9JKbo4?s�H+=9ii�5곳�N�g�_�]��s���9_x�Wr��1I��V{m����6�ӽ$מhN��t64��[�н0U���~���*��S��s�3��]��w�O:�~N���#R��:!�G>1�Ǯb�K��|Ώ�7��k�C^L<j��oչ���z��~�����P�X���_|5�b�h�M��OJ�5.�g�<�]v .��iV�9�����R�$|L�ͫ� ��<,�a�(}��y��3�x�Ty����68?e�ۮy�k�B�d
���%���n��P������#+ق��U��1�oi���(��,Nu�W�墷=�������	؝�+Ӻ��ĺu��k}�*A���X�17��%I����we�o׏{ޫ��u�>����y��ȳ��J�;�	
����v��s{`ͣ��$� ���d��o�v�|4~�-�]lz�ȗMPF�8�E�����TTV��H`�ɩE��H�彛�͕�L�{����7�n� ���.��0eSH�T�XFa!�t���D7벯����Z���c�K_M&���Ԧ���Nh��* C)�����c����-�"_��b";��$v5���hnr�Q*ΏCim�T�+�
/�N���`l3ڻ3��v8�'�]�\������Մ�yc�],���o�;g�n\N� ƻ��l�ܺ{�\k��#>��C�sK�5S�d���l���GG�F���S��i��y�8������n�vѿ`_0�]�ܟ5K>jz,�Ɏ�Ità�Oϸ�o=(��Ols>����=����w�67�ݯ�>�c�y�Aަ��91��1�ö.8V��t��15�v��Eڕ�6�˓��T����p����J��K�4)�ຍN+xfNF]�w��q���\%P��T'*���(G7��_��5/���\p}�������
�U���GN)b�̣u.�Z(�,��E�����V����zn���q�{;�1�ݯd���L�In����|h�;�|�˴mi�2��J��m���N��}s�v�&�W[��s��G4�+J?�u�ʙ��*%h�p�<|��[�_,[<3�~/��T �8�����9���k�y[7�}�n���pyV]0Ǒ/n�U�.�����K�@��z̞Z�B<z��Z���j�`˟W;F��æ]�p�&>YE�B�*�S��t�Bdg 7�5{r��V�V`�(cZ���>�D�#^��T�`��(]uܖ�g�����w��K�ԯx�w�b��bX�s,]g�̯Rco��b�#f�q œ ������:89Ww�	�� �[��3�O	�޲�`�_)��Īmq%:��xް�Y9!׷��yy���)�Z�[h|��@k� �#0��BO-�G���P�ҳ+�ZͥV�nf��������'�pL��(�Vۑ�XV�wO�z���� t����=b�qDbz����H.���LP���/�6�Ŕ{}1TW���Q��	��/�|�6�B�N|v���z�� ׶�������l��5����ܛ������]i�7����^]z���RC��b˘aU�}B����g�[�r���rd���3Q(��b��r�Z�^��|��5�=�^=f_6\�ȝ`o��8�|����}m�y��|�����~�w��|<���`��XyN
͊�u����fuj�w;Y��V���c*s|�z��dW|��>�3��g��W
���[M��
�CӦgV�Nop@�������j��ݜ�v��Y�b�i��$A��Ü�.1�&�yz��O��yxw�xr4�����򨮅U��P��+���.����=�O]�y����y�d����-��k�[U냙�=3�)�"/� y��T<��XʯM���2/uK�<�a���M�5���r�t����3��!��	>]� ���m�:\�_���:�F��x�sm���oJo�.�����˨�וw�Z���HՊ��<��]��ڔO]���κ�3��@p���1�d8���0QN��77�38Fnm�[�x�9�1�}὞�B}���>D9�w��e�7�ML�m����b^8�`j
xO�{}`CxjR��Mۇ6��2��F��ԭڽ�����6+�!&�f��v�s������!�@gO�� (@ʮ��"�����JǙ�:�e-�H��=X��W5���[��9�ծ��~Qu
ڝqf�.OV,2#�m��2����ܝx�J��{7���
���;RKߞ��}`<������Zp鏍��W��kX�p�]�c�f�l^"�J[y��e���<e̸9W,�͖�u������u������鵝vJ5��x��t>�� D*(��dN9���ܳ�^>��c���>u���պ���[�����()}�wS>�Um(��YVؙ�'v2��hh�u$I!����)�� ��"f�l0�l��.��+����M����+�놱#�cu8�z��Av'͢O�M}g�oj^:����Bp�Ji�M*Yuچ��sm�{�s�a�u�%{<�L�0��yh��x����]��Κ��u���%z�`�:J��-�����6�)�whQ��vhp��g^op{��oB�ˡ���{�۰��ћ��<��Wzb��ЕP� �g��t���-�^&�Z��;�a22��HG�x�׽��.�b����;�ϻ+��]�8z
_1P�_� @'�
lheoS�v.�ף�U�H��k%��#�vǆ{���g]D�Kyr��9]���t�S{���g��J��Ŵ6/gU��ЁJ
޸���Pxg5�t��kc�;>T�G(G����"�d��'���O��2
����ʃ�V�����6M"���`�9�0�|0v�V�l�����T����3&���.�a��O���Rg[��v����L[w�3[y�KI��DŋM�%q����t�%K���Q�zh�D�M`nv�[�¶�C�\hb�e)�d��W|j�ڧ�)�+�Z�f;��p���qv�k]�S'�]0���h�:y�sk3�`��hҩ��Q�!�1�r麇��i��쪽�<W����-����5��+�m��0xZ4���@�.��̜�B�:�U~��/~5{�}QJ��ə��\o��m#�q��/)T ].�<�e�>?v��F��z�q�e�HZ��G�3�佁�׭��X���T_�����~ĪP�z���@U�.Y�W�G���B��������6j�r��.�6��%ʗAW*�$=}��>�Y�.p�7s�Z�~j��8-7�� �`�y�3�BZ�E��L�" u���.�C#�:�uzuؕc�'�r���N]�W\��� �Z�TT0_�/CY���:��3�o>��z�_�hj="��x��/��E�#>����Pڃ��~�]@�fi�`5�W��槄�,��v���cD=/Z��o,{k��t]�!�vτ�k��rZ��u-6�=^z�EI����Z���գ2%mTmeL_m��5��e���GQ��a
�_.�.�n�u9�v$�3����u��8��nZ�0g��c΅L݆q5�.�e��}���x��5I�{O)\�S�nج��Z-W��w,���7	R�Hq�^Hu�/��s�?^����*��2a61��(���.	������g�Q���#�{n圡���=h;�l`�����ˋý���!���qx�4&����/�h�g��^b�u�G�0�_#ܫQ�姹4�pAzl1���V�=�R�w>�K;���N)�8�������e =�Y�{f�	ڒ��{'�<��2֩��:���)���p���ch�\���_�G ��)�����Ժ���p�J��">>��S4�U�+�i>�ۧ�e˃!B#t� # y%��W����o�,���Ϫ.oo�Z���&,��~����Y�A������쩕4��@Fr�2�7����ޛ���D?�K�����A�wc(k9��.#��*�_���t�.>Ë���1��޳�0��4'�츀B�i:��{�0࿅�h��&6���b�荗r�W���w�Q�\�Q�%���$�o�c@�:o�Ss��Ǯ�$��,��H%m�ت��F�G[���>�:ޮZok+EF�겝�#gUa�/�QF��b�.��2�]]{��3�3��tG�]���s������5��Q�U�n:�)�� 2���9���I�����D�� f����'�v��s7��{D��㨅N���Ƃ����_yuO˝�P[�̭���㝌�h��m�q;�0�SLb���̺�B���m�+�t�Ѯj�A4��+�,���U��Z�Y��{��;|�>�|���_�N�*��q��^Ӌ!�v�Z�6]�5<�y%5���5�%v�=Ͼ	�>ܻ��j\9c:�PuhFb���&em�_nu�-��z].�7k��}e� ���^��o$AF}�w<�
|3n��M�w@�Ϧ��r�G�mіRv2�p�iI֑��.͗SOQ��ݪ\��]�a&�4v$�SV�=σD��#T���iWf���g�g�uo��\�M�<��*����ߞ���9�_��f��Oo����0]����I�,�ǘ3�(9
[�{訩�첮<�k��c8�A��tx��;}΅vh����r�L1�-R�M%���ٹڶ6s���u�۔�j�=�c4�u�Vn+3[��[81���ó�{����0f$$�b-���[H�#&1F�	��+����Հ�5(vea��FdL�^Cm����q˼�&>T�׽ux:�5�-�`fA@_4+�*U�x��Yb�2M��	�4=K(k�)5��;IMx�L%���s�����Ւ���,�Fk��\-ч��C��,�X(�˦�$ T(�{�A�V)]��$�"D�P�-�\q�3K(�!�\����U�4����V��2+��nU�a��ǂ���e��j�,��v�\;��X	6�^��Z�ɳ��C1z���͚��B"�m�\��r=�N5�6�*��wB���2��lS�.;`
/����� �U0��w�5vՇjR8��ۢ���umǮ
�@�C���6����a�ePv.�V
ld��Z�1�EF�ܺ2��9�L�"��X(����&�eJ�yr�T��5V���K��Q]A2�Y	�qPUQF��t�&+��J#1�r��Lbn�D�i@���7U�*�[���3%�#+�qezi�]�fm4HpP�Ʌ��Sʚ�ߞ"k
�����ɪ�-�&UD�f8���,�V�[D{&��dT�V=ϦE7 ͥ�.���[��AQ�n�.+��Y$�[�,3t`V+Ԧś.<��ڑ�T%9V��� �2�0�e�'$�P���hulR,F*,Qc-��ADX��ldJ؊��
��ƴPQYX��ZՊ�eB�
*�EA�Tcm�%jԤQ�
1V*��)U���TUT+J"ʕ�`*�*�5((����2Ш"�U�E��b"�"-j�������Q"�EAc
�Ŷ��ֵ��+l*��5J��UZª�b�Aee�QRڊ�ҍ�T�
"�ŀ��E�����F�V$Pe�T����X�������1���Ь(�b��TQ#AU������A2�
�-*
*"+*�ImQUEKkE�"�� ��+"�mE�Ŷ��[UEQ��H�DQb�Ab�bť�"��"�
��V"�2؊ ��� |��rө�2�������O��׽��K%q
�|�7a��X7�v�&A$���o�����lHU��O�t��dwj�s�;�^Ң���%����W�����t��Ρ+d���ax��Gl ���;�Y�=�{J�qgk�Y��(�|�
��
���W�2�u�޶K7�R��=	��� �uH��œ���LW���xR�a��]{���ڳ���}j:=8W+�^��kgͮ�=p:n}�1A t2��>� �L�z`B�r�8"���:�0�1����ã�����@򯼗�4}^��s>�K�B�ϭ����uy�7[�='=���CE���
�yc��<6���jߍ^�Vٕ�m�͌xxQ�A��'�}ݸ��so�Y�zʕˡyQp|s�x�24��\�WF���˳(؟�7�䎻�/*=�s�l_�X�j3��E���8�.["���V7�V�^��N�W�p����iLO�s�3��>�E����7��5���7��]<-C<@��g�g^��0l��<#*�\}���b���4��Ǆkn���r�uUu���+���xtW��K[V��Jz�_4��g��:���]]yv��`&��j(e�a�Η-���r��v�T&Q�xcP�'{�8v���sQծqNr\×�B��r�^�u���]q�vZ�۔Q��
��)����{��7�`C���D��_J���� #/�u��3�x�Ec:Sx=�U��z��m���l�{������Y�I��t=�|uΦ?�{ҮE�%s��i|qhw;Yt�^f�	�[j��+�Uӻ3(�E��\�=�V+^�B�h^5���a��t�@�/^wVH�m��	��6T ;��EQu�f�ly�S��*����l�۔ܗ@;��g����7�)�{�/*:���(pߌPJ�����+�D�]���݂�w���p�M�6s��E�ݻ�%]yAJ����$Z���%��H;l{t?�y;�Am�86r��n'{��z�pX��<�#��`�:}���9r�y�/�w� ��q���������ϛ��>���M���HC},�G�(sRb��K�����y.��=�d+F���;W�"�;��)[2^~�6���낈��Vg��_K4<<�j�o�#^��M�;������xQ�t�<�X�:��3�Ҋ��/ �|{[��e�Bg��1ו��>O�����F�gh���!{n�fSQ��{�,��j�)Xur�F	�G�)���ýe�e���֖�c%p�{�Z�Ѡl:2�7i%��M@yV�9F��x��6�W���%Yu�
�Z�I�P�d�}n�R��c�+�W��vu���6/��PC�o�`��$K"�Ct���ӑྭ��\b�ysp��̖��V�"�Fߦ�0|�)J��e
d�/���wW�S���\4����K��&��߹S��w�9~a��L�"�h��H���K������\0^��ž9*�|+���'�r���[x��۽5+�)t9F)Bg��ց�㐑b��V�4;n��:*�����݆�Ggr�͓���;s�n��lA��s�߶�f�:���&P�.��mr^��X�w]��m.�<\��� �v�ޗ��T�pHX�}+.	�ك�-*�!x5��%2�}��^��o��	��ȝ{+iٯUg*���H�:�@�����Y}1}/*��ʹm?p��7�S���N<�CR�k85ў+]�^���޻�PP���@]r�')ݑt��u�u��̙y�������53�.���	��A��]�.�PF���$��S���;�Y���47��Y���>�FCv&�֝�F<�b[���g�:␁�Eo� L=�f{-xd�@Ǽ/��7`�雥Fee�l�z�ݭ����X���^�kč.����Ī��b�Yb;T�[�7�-tZh����w\0�Qyge����w��+�ríP�����q���:��R�l�����qg���4Q�ޗ����p�F�0-���ꯑ��>��g��b����[T#VV�z k?|M�����םv��\�����V�̋\��� _�����b#n;��BC:"O:$h�9[3p��8�]P`P�N�(��v�cJr��s��}F�����}�0(2������w�� x$�lސ���K��۵t��Хw���u4��'��3TGg�򇨼�[UYS�u�g�����2�xRhwݞ4f�!-˚or���dqwZ�w���|�.����t��?m@��W�;�j t���o��b�p���.cr�x�׷r�i?7޻��l`�91��˃j��F�k�M�r��_*�$|�ɧA�o+s�� mLۖr�fahA���
|k6�=�9�]�|��#�co�F`�5��s�)�1�Tg�y,�{tc5�n�jHy��=���P��O��
C�X�@� ]}��s@8�)����+�^k�4��S�zN������2���8�tk�Q��^�r�e˃!B#oB3��|ź���dE̬Ǘ����]g��Xb��ǘny����ۯ�J���	oo��}q���0�ٓZ�YoWq*��3q��շq�9���th�Ni��g3{��9����sV��骎�U��YR�
Z3�)�r��+*�T��_諭��R�c���GX@?�S+�f�V�"�]��������U��QTU@�����<wn��zU��(��:����e	�+�bU]�s�^&>]e}2R0	�]�&���=]}���~��
�7��_K[GՍ�5C�r
�w�o"�^���>���[�L��ȳQ^�y'������R�_���[��&Rc}eh�ML��'ͮ$�U_��7r@��q�X�3�rxH��GM���>����F���+�-����c9'�.T;jxP������W��>�uu�T����2�
,�5�vL��n���w�OH�@_��姺F�嶗���+I�yS�o�'t0�ȯ�Zτz�^;���������� d��9�R��`�%�_dx�9�v����yT��yM0ܟ���T���t��mg�RhZ�kX�n��p�5�*E�9F[j�ӂ}<�#3Ԁ���)Ua�ok��<qk=J?A+��;+��5�ޭ� ��]�Ä�{*��}���Zk���;�2ǃ��+��JZJyI3��e^�ڃ�~C	;�=�]0�(U��7����y�:�I��0��ϣ�rawȩ��9c��;N���X�Ny��</v\�/y��<�g2�c���f�h���sw�b��FT�\����*�=�w(�T+3�F��}_}����ɣ��֏�7�&�)��7�u�1����$O�'z)�F�i����_#�y�/�V$>�h�ϟD�n�9�Qp~9��ʣ:�9]:�B"��Ӻ�x�Ǽ�}�m;}�9����G��m��k�5�pK���^I�Z6����nW�[�`Qٻ�P����j{�8, 35��*�D�K�x�l�:͌�o�.�������W�a|5��g_�0���z�O��Nk��&W ��
#5m�87	ff-ixFz�^'����w�VT�{��� �W�R�u��5AS��A�}�|��Ysp���Uz�)��/��9ʶH�k�i�t��yq2�bb���w2����T6�,�e�E_Zb]5^�;P���7����6���G��|!�:z������d*�ώJ	1�n�����uc�3̺�k��޽RV�A��z'�w�'�tn������6*P�n�P_Ң		W��(1���{խ��Ӻ%1ڢ���΄���˯j/�H�Y\L0��9Uuy�Է&�H���6�hj��6���ֵ���=߮=���d�ñ�^$���)GC�sSK4��u��"ѧ��\���9��~s%��������W����H�t�$��x�{��%��s{�\(Ѯ/���m���x/�e�f�o>�Nk�����������B���u�������V���=U�,��`j�K�� ��,$u#m������/x��c6ӖE�MM���3mx�:@l0;?��0���smO<4f��zw�3�D�(\��[Eâ�*���ӓ��2��4<�	���>{}S���]{�~@O���j|�v��r�f�{,G�*�6Ļ��e3K����ރ\��ړN���R�(/r�:WK�t��S_Ho����N<L�l��yF^�'>��u�Dy�M������Q:+.�]��(;'��e_c�T�i�����VWG�X���Q�О\�Ԟ�{���Y:Jv����3�P�F[��7�;��
Bz��1��Kե�kQ��is�C���;�.�����W�ʿxQl���Jx�޲��.��R���W�G��o��b�8ff�u��}��/�����Dc�2eǦb�-eV�N�Fh�L?��F����"����c��<X3~�˳�-8���G3�zй}<�Ǳ��F߽ҍ�������l�&���0��Ի��N���v���o�r�k�;C;�i�{:��pt�qBᦇ��_o��K�%�5�[|9s�gG�ܽA�㠱af�Łv��nd�l.�{�6I�(�U��F�M���ǚn(wK+�r�(��s�ś5г���ܻ9<�r$�g��)���Us4�i��{ θ��*罉�-@_u�N��G�V6�ꯪ��ٕ��^{ѽArG��pV|��³4 :�v�K\�&A�~��"�O+�V���O{˖赡�����sU+(��@W���,&P��R��]r������.vH�7��U��W��<�ë����وL��Aؕ�mPF�#��(N��Գp,�K��J%�H]^U�$.b3� �~
���c{����y�2�� Ƒ��{}Ӵ�Y/{e#ҟA71!��\:���]5B5tV�z k?�!� ,�ߙ�j�����w����H�����S/q���U�eq?	�0�F�w�+������,���fb��U�i���hn�(zz�ר*�C��%�T6 W�挪~q�h|{����7g4�E0���������D@7�ծ]�S|���<�	�����Ƚk��z}u��(�8y7r����|u�B>��-���
@a::<���g�OE��>�Ȟ�����we�n��{2��� 1)��i�o2f82�*Y��W��1c�qcK���P�_b�<�E���ʏs�w�·#gY�Ԗ{�I��_�(񅯎wu����)����q���:/����������k���������<2���>R<K.��M�n|������[2Ȃ�vc�΃��73zI^���=�>�&u���3�MF`ϋ�l`�4����p��\�Dz��G��:B���u��7)%<��w��2��\r�A0]=+C�}Ju�b�^�p����o^u+�wa)�F��^z�ִ��z�t�Z���mE�/A3��F�v�߼�/���tW�	�Y�:=�w��ɃO�3(*��PC��>{�#�y���Xؘ@�8���㪈�:�2�ٖ2���ܪ�˧��ˮU�#g��Τ��;��˲�*�K�-Ph(�|M��7օ{�i��#xZ3�ǆ��k��o�l�k���3�@S�X�J =$�ϧ�լ:_Ļ۬��U�H�G��Q?+�ބ���s����>��G��݀f">2B�$��r�/(%�Ў:1U��:���O����ڋ&b�J���(�p%�L
Q(�V�e~�I��5��C�*�#���^��z�Zo5�xw3ݡܿ�9*�l�`�O%��O:<_�+����-�X�۩�oI��1��ۇ��Ydc]˯>|�ިz�a͌��a4cN��9��I�-뇥�t�r�9z�N&�$�o�{�9��/@1g��>��������ާ��x�cv����
�7��]o(_ƦEu����T��v'9�c\OWo�{�x����6#a6gv ���
���J@W�`	���G���^���z��R=#����֜�;`Y�wkǕ�5����C�F��~���dڽ^^���tOC��H2�Х��@�~�������F���{B��(.����V�8pX=�i_ϓ�4�>gؒ�N�PZ<&vM�6F��o���U����V��e����C��u��'�������t���,��Iܮ��C�t�쎷K�FX�Ъh��wc�ZjC�Qp~8�2��L�t�A�� :ݷ}��3t�������j�(���Amn�|;��Z1�M9�򮮉Csk��͞����,	g��5���V%^�J�W���6_-�xs����=W�-�O���4Vd�:�J��J��٬��8ֲ��.�c�%�|̡p�>���w�'�;-�o���҉o����LW���@1�=�̋>>DH7�
���������C���+�!jXo^k�۬4_�� �H7������P�"����"��٣��U�R{�)Z��15ol��,3"���-���R��!�ôs�;.���� �DK�>�[}]ӇFVR�n����ͦ�̇M�Z����{-������C��6��p���H+�p�*�]1�j9*���'�{�t�/;~p$�����&a�	)�q9f-tX��3s�/�>(!EEq�{L"�[�^.m��D�_j0x���～i]=y}ۜ��z��:n�$��^��h�4@#���jK��}ЗשP�dd�2�����Jz,����ڢ��N�P�vvZ��Kɏ�����J�k_<�p�unK�/�G�o�˳��h�����_q\�A���V�>��h2pf[�z��̓�<���N��f�;#��c%��i[��C�6S�^s���o{��:�p�������\�b���u�t���Rvb�vT���XSא^�ќ��Ҕ� F�r�0@�h�6���)��#�&�m$���mr�'[�u�Ȳ҃.�Ʈ���>Cmw�:�j:���7�I�BP�cQ��:/.A�e�x�jǖ$=��[ڡw*M��6�S�|��a=��|�/s>R땉�������YW{�������R"���[:�3���Jy��Qx��1���-'k^-��2n=�}�@����w<64��}"ض�wZY{�gQr�Ӭ��ke� �0���Qy	�F!^�y3hW��*��7�V@�n��rܨ��fˬgj7��,�}9*��:�nK![�L�q�4��e��D�\�p�|�i<� ��� ��B���t7pk1N
=�i��%;��V��,Yt��i򽭛�D�m
�����gQ�Iѯ��9]����෗-��6�;�*�q�ƃ���p�=��P�$���e[[�ռ�O�5V��{[̱��BZp%R�a{1�
乼/�-��f�mom�fn�úq�G�y���#�jV�������X�gGvX���)P����6l�pWb��ܸTZxd��Om�A]7
ǖ݅�{��x���f����LuZm��2��Z;.^V��w=�k8�!� S����҆J�),,�"p�I���Wޕ�Lc���B���ˮ��P`�Kvi�2G�n6�f5�K�}��h0�����{r��S�g�6^�,�4��s�Y[/S�B=�W	��)*$k����2ak�(k�W��3%AßZ=2��x-�DVf4r���+*-Ǖ�^7�VfJ�=VbD%��;��.�G�?iӀ�&5�_:�^�DT�{�`6��B�w���#ϷNx�^Ȋ��>aboF��G���o^\�P[�7<�'�5_�V�g�+D���m���5h콨��Wz�;ލ�����R���>X�O�=6�z����IR��
͹Y��������v�MϤ�}���%�C��xy��4��͞u-Mfp���`ṓ���Jt�����񧃞u^��X�-Z�Ӝ������F��csR�K�Z����G�$扙F�ȁX2�S_+����G�|4��v#u�F��������L����߷�s�|~�b�UETb�����DQTV1k""DDUKB�QTV�UF�l���1TX��E��*�U(�TUAE���IF*�,Q*�ł ��Ԩ(�P���Q��",X��X"��
*�X-���$YEQ���b" ��A��*�AcQ�l(����b��,QDUEXEDDTU�"����Ub(�*�X�#�,R
�Y�H(��ڈ��UR1X��Q�6�"��,1`���,�"*����1�Qb�`���*�
�+T`�eQ0X��V8�H�Db��H�UQX��8il*���b+�`���0UQ�",���� ��(
*3H�"��E�"�P� �}��F_��h⾷�/d�hv��ksV][�
�8|�&`�q��1a�;�����d�y)fm��B����������rٮ��ϲf��޾�0����k�@�6�b�������`�jZ�13��|0{n�4nr�s/�­g�qt|��B� U* ��eF���V<ʈ���>�����ެM���R�3�6�/bUc+��
�5(N2�P_ҢP��F��N�U���k�;�[#�2����$��.Ai�yї�<�e��fT_x�Ʋ�QE�(�p���z��BW�����L���5�A����Յh>9�,�Y]pP���a�(`K��3�zk`��h�CvS�+��oFz"M �����׶����y���]/ ���^��i���s"�}�KFW�=��\;2^��(\�<�7C�xRک�O'�ǌjBz���U)�~���@�	���9�T�b��Po�񃂏���Uxm�w����s��6%n��uz��xx��~�iO���v��C�����3�X������;L���/b�D���6W�X�j�::�D�僯�ܩ/��B�`�*1R.�OU/�P��wo8q��i��
>� ���}��MP*���6���U�h�`ܛt�rR�Y�Sq�xd�~�3�[J�gWD:�Nl�Kn�X�R�3�J�%������
����[�P#Յ��
�ź0S���:(��J��}t�~�����7��G�}=�ZX���ORXL�A
�n�d�c�,�'�m��5�(u]��x��=]9����y1R�E�ʱ�Rl��	���8�z2�ُ¯�`��:JH�'�����u�
#���̿W(=u�|�k;f(:+o3��޻B�V?32=���1F�4��Ƒ�QơLo���vU���|bb+�b���W��-�e+օ��L�<�|�̙�ڝm��{JW��ZϯixAY��Ww�	��*`�A�<�P�(|���W�'��m����E�:��ص�|.b�l?�G�ܯ *.[~XL���#R���
G�e�ӥ��㯡���H��Q����e8���]��m�0\b�z�:9��_/un�Ǉ=�gj��
�a�kr��5!&�,O@�}�f��Ct:�vA^LO5�`ͨi�����"��W��������o���B5emצ�J���@`e8` �p�����B��x@�����w�v��$DD\k��hn}��.��F�C�%��Q��-�>��%$5�RḴw�n6i�}}Z�.�������o��n�^!M�cu��D�Iu>�	��Ӱ6{�5���?A��2M�j���-��[�����=�Zm_<3�.#O}��Y��ɿc�s��_:����=w��{�k��~y��k�}U�}����c�\��㪮�w�]uQ��7\�d6 W�dz�>�	�d(e��� ��^�jAĬ�%Y�`�U�P�V� ְQ���'�,�wS��?b��<7�R�)�f�e�b'tÃ'���bU{����T�
Ϸ:�Ik��I.�Ծ}sҳܽ8��o���K��SYG�����E��]�6&%,�G�y^������=y�Si��nկOs�q^�|P��.�e	���\�W�唹:y[�+�@ߦm�;">*/���Z'����.�f:^~^\,��9��9p{~5��1�:��l`�4ɳ��@m�FN9O\�#���`��%+���Ԑ}�[ͅC��3���+��t�>`q]:]������l�%H;L�z�L��;}�`V'�NL�y���Ce˃*%u�q9���R�bǀl���a�@�磓��&,��j7Ѽ�g���e�;Q�]�q��(t*��*Z�dgӳ)	g(��e?`w���e���k	�HvS,��/a�R]��k{`��K�4�E��A�q�%�i�C_
ھ�Y��t���8��Pl�xސͦN��Ɔ�T#�-ۢ��[���x_a�7��:����nT�En��1\�Q�{�w}a�Ҧ�N]3w���}�>�Ik�����E�s߾������.�1��]"|=@��t9(��3�W����+>(�b�":�׵����$O�wug7�k�(J�y7O�_�LJP �$Yer�8���Vf��t1̬�uu�>���ܨ�SѺz�Q�h5S,��p�g�̱���.�0��	xt3~o�/ ����O	m�=�2]�^u��:<71BJ���T��WY�iA,�`^���"(�m���ˮ�<�^ ^���yO�cHy���^)�Au��f�Eu\Pj)f��F�1�Ξo��wٓ-A��L>���؄q�����9B�m��k���,�&SV������.�+�i����ۗ�+m8^�Bg�����̑#|��y��
̂��7y�xG헞|��Z���A{��=���>]�j3�f�!�%�+�ڷ�W��[���su��ܖתx<�{ݎ�p��EV/�_2���˨�9�8nrD���觇���V��ez.���ӧ����uYҸ��1 ��U���L����;�Mp~9�8�3�����,��tm+�-��cr�W��x\=s��'��3��[�<۸�>B&&,M���^����VU˞��^JO,�����.�sr������� Ɍ	��3�ݽ^�Av.MД=��2t�t���̼\��aJ�xXɛ}���{ݲ���I�e��wY�U����}��g�0�^&&@���-��gb�{T� {�i���d��6�ߑ�wQkW��Ed�^mѩ;�z�<���ρ��݀:ĩ�3_���r"5��N	u{C��6����g�ö=%(�u����y+��^l�f�O
R��p��{ �
!b���	���V<�-���a	�h�d��()U{fT�9���L"�n�˛��&��yc�)��ރ�u�c3�t��}�h���Օ U1���X]vY�W
��_�F��ExF��0���O���i�ưVi�YF�� i�7_��T )Q �:L�In!x���r�O��_����}� �S�ƭ�^60mx���N�0�|<%�0)Q �kd��W��;����g	gu�!%�g�w�))`�.�y�T^$r���QvW����ɾc�{�k������xn�CVC��g�n69�l0��%�˔�X�}j���˷E�y����S�8;��~«���+��˞��i� ��PT��J�N�O�ݹw��n�l���n%���94�L�)l@�w��ǚÖ��3A�:aLUv��w���j�� ��=G��#}]���+]�W%��5�����Jf;^T�.Q�U��LC<��'�[��
��#�zw�����'��e�2�+�bJ�5�a��j����Ŧ�c��b���X�;�NOvΛ`i�"R��T�/�#m�����Ly7fw�r��,�;��}U�W�|Z�Rt8�R	���vV���f���4���+��6�eC�P��� nX�:�����+��ð�O���h1�]5�T��<��%%l{��5��V��/9�t�MD:2���Ai�4��t�`\��A��3.��2��p�3�j��x?N���M%����-h�}z�J��q�[��_'L+�>�Ii���j��	���sU���(WK~��}3H.�O��E	�e__̛��vY�V"�vǅ.��I��}}9�%m�;�=W�<*X��ʲ�xRl�P�����4������zyƲ�{|Amqs�_:G=Z���w|柰�WH_m�vx8_z��o��m�M�<%?wL�w6�g�*�}U4��R|�5d�	�u���y� q��>I^!��d�=r�y&{�L��i&��*E���M]���L���@�?<�p�Q�I��춱Ͼ�u_k���0��1&ө�CF$��`m��*dä�ì�B��x�!���>I<�S���fP��~8w��<�
��u������4c�4C(M����=�!�H~M�Y�97a椞fyCl�~d4Zy����4b��Þ2~u�}э�_�'������<�!���w�Z��`W�>t�S�߰�"���;]`Q����ՌΙICZn�:ա=ѹ�O⾢���~7����g_�%H|�Y�����g��&��P�gP��d>Ʒ��6��'�k~z�	<�?}a:ɴɿ�5�u40�O١5�g��>�|{��u�~η_��_`)2�Cؠa�N��@��py�=a0��q��q�E�(O�$�1���MLo޺+��$���O�+�ɻ	�O'���G�}�{_e���5�߹���:�$��]Й=g<�OP0�u����?o����2�a8	��:ɒ��	��?Lc�����8�i�_�B?����Z;�N~���C"���j�b�f'���I�5�bCl�!�jC�?'�k�$<�L�؝H~Hh��6ʆ�}�J�a�O��M��>H�g1O��/�f5�?ַ�Y������~�n���]�k;�`�(z���8�ݰ�}a�?3̇��?'�<�(O3{�����M��l5����*��߿fbԇOz_)E�5����E}�����$�&s��M?2Nl5q'�Ł��q�����Ԇ<�?S����,:��y�ƾ�d<ϐ��2����[��Q�unS�����`�m���>��W��l2��|����O�>/��2L2jg��4��e?M{e'1Hk~�����`�Y��|�d2��:ϐ���z���"�[��r�h����8y���޼,�8��vd8ϐߩ�~����I{`i���.>�טM�n�u��m4w�$��	�oI0�u>d*C�����}����x�Xί|���C�C�q���O�0�N��Ì'S��N2|�	�װu���&��I�����d�����N���?D~���_�U@�\�	�������~9�]�HV|�!��Bu2o8�H~@�q�O0?&�B|�&��=��I�i�&!>;�@�N�ɠ�ĝ~���=�U��O�B/l�c��1#Y���&v����ۘ�W0�b�[eL��s~o�9}�Q�f�
��/c�R�� ���z�.�hVa��ׁ�Xu㭋�7o�6e��9�q.j�\�E���ޔ�+�Ԯ嘉�Los�1K<�5��� l4⇬������	5�w��{����M�?���aM0�|���p~`VC�e(O>xì�;�N�����7����&}L�d�a��?h�>d�݀��l���~��'@w��f��s�c����*��E~�߲d3�o!���a�ﱉ6�!��SHJγ��&���S6`m��c�M�W�?2d�͙|�y&}��}�^{�z�����k:�9I=θ���y#�J����?}�E!��'�0�a��s�I�u��~z����M��'tg�'�$<ɶJ�����.��럌}���7�y��y��?0=�q�$�M��w6u9���2���O�*C��Ʒ�!3����6�a��$�y�d4~)&ޤ�����O3�����u�^�g�w���xx0���������*u��� u����"��S�<�a�3��S�������ِ��x�O�2g44�Xa�ɾc|ǻ�wo�[�<����\���}�g�?0��d�g�P�J��:�Rs�LR@Xb{�	*���<�d0�sX�Y�8ɫ�}����<ϒa?l�]�k����[��s�I�L�ְM�VJ���I�N�ya���C<����!����g���<ɟu��d�<�<a0����>�*������5{߱;���P�I6�a�{$6�hǾ��C(|��߰N�VJ���N����i�I�?D+&�Bd��C�a�CS�$:�)׍~}PW�J~^��~9��۝l��v2O��*Vd����>I�y���m�$�0+���<�P��k�!��CP�M}C�?'��H���
�*��k�߬���Ȳ�m�tN�I�C,�{��>d?$5=�{G$���!�6�L�^�3����L�2OsW~I�o���`o�k��
|Ϛ��
�\;_��V�m�}I�_�E�����M?�+�j<� #�\��N\]Q�lm�g���6�
"��,\�Z��ն��FMt���^��s�>E\۞
������*�y��yME�s�g����M��s�;A�s��b��.3P���������������}��q�ݺ�C(u4�a�2f��=d�Ʉ��`��'�O��`~C{>d�&���2L2h�w�5�$��k^����Xi���u7�����������1�:C�C߬�|�,8Ì�Ha���6�y�N;g�}�Bq���~O�2�׉9�w���d����
o��`�����;�?-ǅ�#���?o�~���M�����2��gS�Hu�o�2d��3�u�Ə�̇�<��	�~g}f�a�����<�
�W���}�������~?�V�%���O����	-=�?W�x}Tm*�_T��х����~HVO&�d:�ݡ�C,�a�:�����N������r^�|�M�}{�o�<��|<Ʉ�p���|�RsF>����h�a���PǨm�������	Y��`e	�����H|���q�O06��������{��	�z�'M~"{�w���L<�d��&}�I׬�=�I���y�R�fO�"���ěN��S���!Xu'��ĕ$��$6��u��Ü�1���~�:\}߱��e��h{�!�d��2��y����y$���@Y;�&���8�Y�{��5��s<��CM3�m���� Ex}_�O�s�����FrwB��|�W��>3a��z�j��&�+�5���C3T�'�5�����y�v��'Y3`�!�M���a�ϳ�g�l&�3~[�7����wC�9���}�}lp��'�~MnÌ���jc�C�p�:��p��)00�=d�I����L��9��u8ɫ������U��Pp�T�������n~�����g��CI/u�?=C,�߬'Y4�����N�wa�L�Hh�ya��
�y�`>�0�d}_ O�}(���V{�3EłJ �����m�>�>\X����6��re��̪$��{�X}��s��ЯI���s$C
�R�֯Rr��{�eY͔�N���A:��7�vk����^����/�Lw����]�p3�Nd��,�Iu���o��E_�#���_W�R��wk��}�~�@�0�RB|ϐ�� ~I?�?}���CI?�!�0�'�?��'�m�g�2��g�I_2�؞@Y/�5*C�k����Z_�k��5�_����c����q�2fO{+<�h.0B|�'�o06�h1��I����bN�VJ�����Mg4��g�I^���e�=����
:��ޚL=JW3�pG���u�6O�x�@�̙�!�w�eL0�fN{+Rq�%߽��&S6ɦ~a;��$��f���	�J��	��N�|��q�_�Ƿ���?t=�$��C?&�C����u���rM�<̧�N�`s��+0������:ə{�l%d����4��=�X��UwUY?w�ߜ�߫�آ�g�,{_�Uk�P�3ݡ>`)�o��I�0��d3=L$<�!�:�(O3	�S���6�RC�Y*��>���L2[��Ϗk>9���;�}Ƿ����������)�d�<���T���l�Hy8S�u��(u�C̆5;��f�2h��L�lԻ�4y�AU��h�_xW�1_�˼��]���{����@���G�c�$�&9��&S�]ęI�Oo)0�u��� u���C(����d0�d<�'����O�����r|pы�����Ͻ�s�M!<}�y	+Ě�� ~d�N���&��s��u�e��߹�?0�~`led4��Ѻ��M�C��Y7�����Hm=�~}�������}���Hi�&��n�l'�f��0��h�>�����a��
N��>�'��y�B,ٞbO�/l����i!Y֫�*���U��O�*C��ۆ�c��s�����������Hm?w�Hq:��?3�RO0���a����IǬ��ؓ�'t�5�3~�C���P�k����%�o��N9�>��!�i�C�ˆ���	s�����W3��l�:��<F�\��b�@�m��j��Mw�75�"�x�>�I���C���Ւ�5#�����`.�Z�e,]Գ8رBV�4�K�O���S��*'*k�Q����s������c�ut�lT�ƈ���bYS78�j�|w�ҥE@n�Ð���|��I��ɟXщ1q���˦ʋ��r�b����N����MU���bS+�i�	1�;���]�DD�!uL���_�� �m]$iK������b�	b�&x��*B�dx/��.à��Ūcc!�����}��C�k�%z �#����i���gI��^�`S�VI��c�Ƿ�P��}]���0����<0KZ�zy��cF���Z:\�4��ۃ�pc�>�b����di���0{�A�ơ�F��);T��`/WחI�C{N�<�l�G5�x���1K,�������
�c�mq���^��-~8�����~��.a��&�3��V�H�[�Ǵ�r���J�07�b�)�f:Z0n��Y.��,%�-�诐U���JK��1�\ܾN��!b!�h��Y'P�Y޻�lKL/�v��VbW*s�"�%��]���7���8_B���\lS
�i��\�m^ҷQ6u���Y�Š���n9��":5�ܥ�������UWzr*m�d��]�G�Cv&�ê}1��7���(Tn.S��|���Gw������>�yv-j����H���%DC���n�ۍ8ff�.$��[R����"�����#RU��Y�Nd Rv0D*Qo���!���8�cw��d�b��#����"
�(��|�,�T˫7n�
A�,d�+�xY�X�v$r�t�2ߍ����	�st�p=4D4r$k+34C$��xpjܤ`+� �."Z�4);Ee��� 勒��,�0����6�X̣&f	��Yc�A�N���j����S(;��Q��F�1��̬d����r��S�B���2�>wH��(IV]������������R�Ҷ ��t�La'-��i��U臋 P�6C$��S��tF�?6�!��R�
�yvr]�,��+�����nhW�Õ�����kȩ3��j�`�ʰ�L	,�-)f�h�k2]��ٕK�sl�"i2��Bf�hm3�0\;�pe�V��5X�X�A��2�X�.DCA�G��Qx�˸l3YWG,mB"�k�[4�R�`9�5A�b騈b�����i���O��K@�q�q$�<�(�Ö]+��:-�&���������cN˓�^b,��	u�ݙa+yQ�� ��-�A'yxBX�JI�Qa�O�A��T�M�`7u�YБ�ܺ|�Qm��o[�0 ���(*DEU�?8` ��TX��,UDADT���Q@Ub�)hTQb�"��+�U�,b*�V"(
�Ũ��VDTF-L$��X�PX
ȱAEX��ֵTX�T�H"�ʢ�b���Ȫ*!R�QUD`�")U�a��� �,Tb���aR���(����C+m()"�U0�TUV#�jPX1�"��(
)���(E�DdX**�ADb�DAŖ*)�`�E�E�b0QX0F#* ���5%DD��E-���%dH�E"��+E@X�*�m�XJֲ�"�����W�9t���m�2墶�+���h����:�"���S\��#\�	 ����j�Q�僂������+�����8t��Φ?wM��:�~u�BVe����!���hu��f�>z��z�Ϭ��6�&���$����Of�h��@Ru�'/��0��'',"���}��c_�}p�����M2a�c�<�X����B��8��VM��']f��<ϐ8�̟$����u��3���$�`(i:�nsب'Y������~Q��Oc��&�d=\Ͼ�>��Q���2Bfw?fu�a��bM�����I^��s��E��'�J�!��u�̗�4v���/$�I��5������?{��~�uu�>fP���
É�Gԕ!�y���!�&���!�M�~ğ>a���XO��?&��y�'���6ɗ�CE��
N>C]����z��Ϻs����9�� ,<f���(?{^��+2�_̟�u2d��e	�:��1!�C�ky<�l2~ֱ'��Γ����LϬ2�I�����y���s�����C	1��i����
Hq��S�"�����L�M� Vy2h��e	�䟱���Mc~��Xm�,�	�M$���>����\w�2�yw��sZ~�9�p�3�L0��CN�O�h�^P��l�§��d:����&R7�eC���C,�2���m�N�ف���q������;�gxξޟ���{����N�W��w�8�Y+�3t'c�2�$��,0��u�����C�0�a� VO0�d�:������m�0�~a��
�dѿZ�����ܩ-����6��w>C���
��%�ɿY'�'��@���,'����/(}������~g�N\$:͡��I�'��?���C��g��}?w�������2����{+R~I���]u�e�l���{���Ł��,����<��O��"�<����C9�3hq�n������������xq"|{P�m���:�R{�]��ީ+��gt�`�k��a�]d��r�+�G3uM�S����W.��^b�\�����hY|�h8�2��,,�k(�`��˸��u�����M�ؤ����fZ�����e�����~�~�9���1����4����}���d�>Cx� |ɴ�/��2L2h�w�u��e?�$�Nb���"���s��!�C���<�e�sX��}{��{�w�>n5���a�!�C9��3o̝a�	�h}7�`q����:ɆJ�%큦N2l��ϘO���g����)�J�Y�3߱2��'R�9�Ff��[�8M�o�g��S}c����䆐5�g�i�v���a��0�O����e���d���I�wq���}ܒ~@�ǳ�i:�V�;�T�T���?Tz0��<�G����C����	
Ρ�����'S&�ԇ��z��ɯP�=I�5�y�$��̘x����`w��������Wݾu���2=���>�x����R��>M0�=s�jM���L�gP�5���|�0>��y��<�����'�9�e�$�*U�W߃����ol��U���g��3<g���&�d�Lc�d"�gx�C������1��`~�4������m����y��-2m��
��}L}��T}>��.E)~�f�[�R���n<a>Iߩ��r�z{n (y�H8é�?}�E!�c��!�!���ěgP�Y��2��?&�O��&q̞~H}�w�{���������NsX���c�|d��_��n���I�ӏRO$��e��%y���u'/>։��Y�?}d2����3�|�a��$�y�X��oRi3�����w[��|k$�����2�!�a�N��,4w8���#��Eϳ'�,"���a��&��4��<����̆�:���
��}��������K�:9ߤ�;g�����N��a��ə�x5�u�C�?9d39g�
Nz�F) ,1<S�E{�y2�a�kVC����e	�:�ouy�n��*:��D�� ��s���������Sc����aV��ݛ�{����ۗ^��b�$�|lMͻ����z��)�r�h�}��^�����5\��;,��9m=�Ŏ�ej�\��gc}��T�DVj˦����9Н:E֍�K�w��H@5������c��78��	�=|���&���+�$�d�u��u��+�C��C��x�)0ɯu��Hy�CI3�q1|>�[W��?���P��~�������Q�<�y����!�F=�O0�&_�6~��y��WНdP�}C/�O!���e��4ԇ���!��ffoLo0/��2�߀����}b���A��C	����a�L�`�I�䟦1���|�;�kԛd��$�&�o|n�u���a�I�a��������:0:��95�}�9��s�{	��~C߬�`m�!�`�!�!�o��ǌ���F��̙��g�&5�o$��$��q'��CF��,&�f��O )�b��/�_c���?q߱�z|�B)=�����d0��bC����d�ɴ���<��	�wy�I�����?2}}��a�F{�ɯ�&\��p����vI�;�UBkn���|�<n4�p���>��C	���:�,?}a�u�0�C��a�P�$��7�<���?yJ=��d�{GwVY��Q���Z��t�n���8���UW˺�m���/��y����J���f�����W�g:��鴪䛕S��S�����l%vb����u>0�����+Fp&o\���#�o��M�q�򊽕�/���9Gg��LN]N\��mC�,�W�s�S��A�*��u||G?t�w ���i�Q�?76���N/V$����f�3`�T,7��1�����V��3�]"�����ɱ���N��j�{�0�]�,��1��/Y�_L�J>���{��=��<�qVm�Vs*�ޫu�����W�X����̜��,�y���dZ�e�DVgL:W(X-ܙ�ޞ�����
};L!��&k��T}u/p3^X�MGʜkC����+���e�`+�}��٪�z]H��z+�*�!;�^7�Ȫ��oӍBm�H=Y���g|.���4z�n*�崚��_Uj����]颷�N]:�q���ҧ�;���E;ͥ��\�j������];F������ʭQ� ��Y}.�n�7ef1z{�.�ܢ�:z�CU2�u�eӧ[�^F��^�T�	�g�������b�sO���.�WB��Ƙg�ڱ浻�޶y� ����H�*��']�2�ݺ3�W��1�V�0�s���y9fk���	�[�z�@O@;D�M-,۱�����e��Dv�K^��_X�X�/�:�eˇ�{��ܿ� �z2�6�9g_ � ��2��%;�Fx��v|������'�� S��uS�iaU��!w�Ԝ���1l���L+��^�\�3�_m�_}�Ceu���{l��1ս>^�­iV��t�Y�Fh��9`Ԣ�㚀���@A�:�a���R�a�,��or�ؕ� ��U���Q}��;���~K}�\,a�ȟSH�T��3=��
H��FՆ��#n?=��y�z��O̻�##��lE{�k��yb�����O}�n����ң9��3��{��֏g4ud�swSһO�x��򧝄�=Y�x��g �nW��2SԪ8�Ϋ����������������W<��%Xk8f�ous�1c���;�-<KY~sR|�5���S�5��*��9]�����Xgz
�9���o;8=]b���<7�)r�㯽Gc�G~���]J*�Q�y��U�۫�N�K�r�:�g^��֮�@s�=Gv�������ܙ���A�~���IC�W�%Bz��&:��lf�o-�W������*R���-�K�jK��EJ�Ou�{:iO�_*�<͛�1p��#�P~.ð��@�)��t�D����z��T�NHFv\�Xs~�7n8�l�Mr��ߑ������&���p�|��}{��"=&v�m��Y�C��z��46�r��;�+\�>�)9S���� ұ�9�l������T5Ù^�rpńm�:�c6ŷ0E��wu���kyun�:E,���T]��_ʪ���=���^��jo��eq����}=n����B�S����o���o>Oѓ����^�p,n]���3&W���!�9B��=a)��)�-�Ə�0_����>��Z�V{����}D�
sf}��L�����Z�'f2���%gz��N{v�v�ܐT=<:��.�w�g�ϛ�_UN��c���<�x:u���n-�Zc�~�׸gmC�i=x���y>�~. Z�lvDvf{����r����H���s��##�dUC��חÝ��=���>�uȳzκx��ܔוlw}9��&�eG��gt(<��2{�c��eog���B�/ޏ��>����.7#<�{��G��F�����x�_��U��@��.<E�6�0��^W��\Wם2�=�qڞ~j����\"E�AI���Om����A�w�C��r��[,>Y�Қ�h��{M��v�"^�,立;�[�&���Ĭ�\�3�d��k�R��m%�K��\Yu{�[�`�ӷ3�=r�E΀�ǋ���/��R��my�����r�G��<�d3���\�53��.�^��|�>�y�w7\п����-��d{�/Q|�M]v��ƎwG=PzY��֮�f��V��y|�o�ovwF�w��'��=mѯ�In�U�GX=(j��o ~�ê�X�S�O��ҳ��\��.��Ĥ��Rm��e\Έkq�ζ=������z�g��=������Y�%�K�t���R�zC�!;����LO)�ƺ����<g�Q|�Y���U�5\Dr��fJ�=��	�I��ngW�4[gt�b�=���iy��=�bE��q@��M�U���N�cV��@��n���r��渨O�; ��
�:­t�-�h��e�t�E�|�¹~%������unz�9禨��6�/�{����e+x]M�ѯyxc��|f�#�$V�����=��Y�Y1��vǼ���8������w�]��9�U<�8�R�L��W�r�:+�t�sZ��\��T�����_+���ƛ�Esr��G)���,���������w<�b��/�|AL������0�fv���ho��?y�� � ���!]��n>=72����]�D�GR�Ynu_��׻ʝ^]iW��}[�[>��L�P#r���UW�~�^��z%�G�nb<�����r�s<�ˮqǽ��\�G]
�U��9- �ǲ�LYC�*_\2�q����ܗ�<�xb�5�9OY��u�y��q�q�o��;�ݖ�6�ޫx���7�Jf�����oj���������ޗ2n�q�=S�i�ʓ��+�7����~�N��gc��VT[�:z7��Il��SE7�G1:���S��V;���z�k��	��+�^I��[��_������;MU��)y���5f��@������)��uYZ�g�U^��q���D�EZ�M�T�m�Ǿt��,v�m��G;S͊���6��,J�Y3}�/=�+�A��PoEW�c�b�]P.{b�19��o��˽<����m���ut�K!>U������U�N�}6��۪3�W��k��J�9��oh燺�;:�s,��tN�re�>��O��<��kcÄi_8pqct�z���N��&mbMU��g"e�-dÄ>�(ꭉ�⣐v��_&��s��p�
��ۺ#=�i&��Վ����ĳE��]��܈���磌�E�7O}'�w����^�Ө�l���@9P�镩��^�t�7؎���5��=*��L�㑆g���ت.��%,r0h�T`��C�)�s�x�J�Cw�^o�y����W7����rn���Ǆ��z!Z�u�k�>�&�����],��t�8�][UZf����7�����j�<��7�u\���'|nNC����Y���x�z�}.�3et����{��Fuz���^�Y9��^���)H/�C�uÛT8�+��r�M�Ѯ��
��A��Ad�Ҝ��Z�[�ە9˩辡�}ӈ��n��t;�e$���L��7�G=j'޾�u�3g���=o9�[��~���<�
n�S���wɸz�"oӽ~���ޯ}i3��G��}+���^�����>�B��y��۝�b��BW`��oQ����򌩂v}{�kg�xu�-�)=���$J>�Ʊ��s�����)��{v!}X�7�K�x˱l
o.���u����յ��sN�X[ι�[��`� ��g�/Կo+���h`���Zh�
#�D���p��Y�
w}w�x�*�Ү��0��Ń�y��5���W�UZ�^��M��u��r�sӌ���Nx�W�A����wl�8"���ߏdx�V7�[~��K������t��8Wm��n/f�>ܥ��'u[H�M�����Q=}��oJў��t�A��t�ҏ����� ��F�7	��@�Ǳ_x���Q�!� >�#n��������8���{*zԑ��U[���Q}�D���u�d���ý�/ް�o4�se{�jYvg�6$lg��q�W����0˯Gqg�4x����j�^��.Cl^��5���sp+�����P�{:��Cý�҆�j�+���sN�я=�f,��}�*�(W���>lB�V<
n�;6�'SG6�G��M�ӷV���Pqߓ׋*���~����ˬ?xΧ6t�\�̞���g&��w�κ����|����Vd�\W��{��],|ޥ�qaZi�mg����y�,�v�%��i����ψ����^�e��w��=VOJ,�g>y��C�w�9��&���B��30�/>�ݞY&P9�r�ZU����c�.O7E���Sgی��Ǯ���\�%�.�ܜ�{ze��Qg�k������̏/�b�m;zLvv��؛���_cR���VB#V<u76-���R�#o
��<�5�=d���1;����v�]sm�݁yp~:����FoV|�f��Ր�s�i�eb9|K�թ:Q�۠�=
�8�S�|�<Ɨz^g?��m����v`6�����3��9�K�g1m�̋��'v-s]���W��������jJt�wK;g���,F�]bA�ݎ�k���᮳؝���A�/{�\:]��4�D/\��Y�'������Z���lBTR%6��|���y���'�����w%�ԧ�Xq����&���!�]�D��WŘ1D���f�z�5
<y�f.F��X/�T����Xyq��e��«����J�̻׊a�!=Rw_Z1�{Ҳ�,�.��g�9�01�mޅfĴ�����Qeی���]yH�6�đOMTj�(?y0��_���Oc�[����RO(dCTj1�V)�2)w��r���\���YN|�4�]%�����s~-�E��#Y�fL�W��to6[�һ�T3:���>5���!�ylC6eA�hO��a8z.ѴQ�Y)�Ê���Dx�q�;x�����7����l%*̈́��B�rׁ�3(���ő]�L����[�7M6�m�dC*f<�b����6�Zi���>���M��R�E�x�P�4��`�Q7�y�R<v�Z���.:���I?�N%�l�v"�x��7V�Ka�"Dq(��s+˄jLrY��,�j�w����R7e
-f'-�VA�*��0��	�ct��\�W�a$��5A�ɡ�J֭�R:�ُ*SwJ�#���tS:�/N�;f�>�L9fe6f\�iWm�x�{�&�]X))�-�Ixt�U��k���v�S,�E{Q�bo�슭HF��3a����\f��i��J�$�[�
�,V��-?���rc�oV�4�I�Xण��v%����*�+�YSe[$��|�Nc
�ȃ�h���y��f�`twe�.���ZR<n���hgJ����Zt��$Q\d�M=�6Ƣu*:�6�*�gB�`���M3?��[�m��z��w��1`�PX����eE���,�Ŭ*
 ���Q������(�E�T�#m
�X�|�"�!kUeeJ��"���kU�-�Q�������m%J�������"����(�T��*(��`VV�VF*H�Q�EE#i�((���PKj��UE�)Q�*�TX%J�ZX�+Im*DAd�Z���kE�Kb6�إK�SV�T*B���K[DVز���a�-�J�T*�k
��µ�U���h�ťE�"6��0�PF��TUY�����,c+Z�*�81KB�Ս����j(VJ�U�,Q�q[@�E���(#�U��U��00�
�V1��R�b�0m�-,	b
+�Y�,U٭��=q�>&c���9�\A8�Ȩr�E]CwsOs[G%����0�f`~xv~:������$�)'1f��W����Wy�D��4�φ��z���2�sܧ�\�z���;�A�y2n���>i�l��j̸���V�w���l��+��ʾx,;c�ɫ�����	Uo���{*1p�+�����v���71{o�Eo:�����k#�\�F��}��p�U^����cmqt����}�mJ;6�k�t[�;�2�V���Ҕt�Tu��{^�}0玵��	�_����G���e+���x5��]%�MU�A�({Aߵ�*��G�l��9��;���z���xE�j�8ό�Ҳ�m�u��	}1��H~?Z����yb�.2�;qf.��n*w\�*P�$#w�`����D �Hp��y�S��<�+�Q��G;	�+���z�/��*�(F%���<����x	U[��W���`�i{T�����뾗��U�h��k���<H~s�����uh���cO�=�S{�S��%2�7�&�Eu����B�����{g_���W��yo�*n�w�f�,��eNT+Ud�wsSG^j㖱�[p�.W25$x�H�)�����,�������V��I�(�
��ͷ��着����,���J7��n����J�@9	��D�y��vKaWT{^`
0·����§�nC�\�S�.�n���}-�Ug�lN��^��G�ز�9�Y�wmJ��_t�n�޳�!ϧ���k��uB.=����1�{���_X|�C���ؙ���ό���5ޓ|����,�ۼ���-�a�[�~g8��E�%�|̺]����:w��zI]����n���p����+|���6�+�:��o3��jo2����mj���E���?S�t}�׾��,O��f�7N�vu����[뫸���lW�f¹y����?�,�Ǣ�J�N�ً����1�ʢt�=�U��Vz��5��i,8N�|���t���8Z�)󡣝�պ7�)���]XM�s����f��,�#ʭ�9=�&�]s��˧h�u�GO�Cv6P�����uk<�Z�c�Ϊ��D��F��2��F���|�2�g�,�<���g���ǂ`��S�{;S���+�+�I,��圩c��Gr���ڝ4��'�N���:����wd�!�Y����Oig1�9W���8��խ��ש��y�|�hu�ݰ�_H��g�n�Z6��$���Z�YC���~�����F��h�3��FR�#�o̔�R��U^�������Q+��/��/�[�c�^U_N�(�J��b�0�we������NC��	}0Z�eT͋i���.ꡊ����E�}hRޚ�Gy�����eJ��W�N�|��R���g�7||���U�r�eV�r_wH��P7+���lJ��xz	�ze����{�Ԅ�z��]M�*{9���Χ�L�.��mN����@N��T�OQ;��u�!Ԓd�l�V#�O��7����f�]+��׋�-���.\)Ƴ��׏kw�yi�b%QW�N-[]2v����l�}B���2oό}�3Js��c�/�I���&�kY#�����Px3���AOz�t��J;�;�|;��a�͞#���}��U�u>�rr�=e뵵mq���ʯ�}.^��� r<��I��o��Y�#;Ӯ��=��y\dz�cyTe���,x��ƇG�=�Yoӭ��We����j�ɵWe��]LwԽ��s���<�`��r)#{�P�nQ�2kD�u�H��m�קnWW[������,����Mn���U�J�Ƣޝ����"/'���\��C<ا�哞��2�Y|f�|���}�O'�[����ۧ��[�o�N�ޙv�Kq��̣z�x�����E�v�]��\�?F�m�=���z�^�87Y.R�>�����ʲFE؅'��2U�x|��y�o�zZ}>��O12���Auf6s��'����z٧y��3B�}4*cx�n��ϩ�5A�:�S5�C�R�b7D��]�>�r��F�v׆���=����C�M�su�Z��R�϶�2�S���Q�jt��CYU�s�l�f�"��/'�y!�s��eI��Ѻ}�doX�U^�Mt�L�a�������\��N��=�Mȣ�n&��rMW�f@
�q�D_S�
����J�@M)j����`�&�wJ�yz�X� �M�r]��LN^��+���R��\/e76Ӹ��RD��ϭ�X�[Q��󷯣����s{�tq�#0[|�qnc��3f�O���v.�p�yk���)���'jD��ђTB����)f��X�[�v ����y��Yo]̒��}�1��08���]�2�}_U��7���}m=_�f�.�˵�&{����}A{:��s;C3�����d�y�wxAݨ���ϲL�7V�~��|�ߦҴ����h{��݃J���g,Z�&�7��i���"���/zeE�I���g>��ҫ!��+��X����:�Q�w��3�<�}5����u�FG]�P�_V[Z�Kdmyۀ�}[�,�vL}ݲ�u�ɬ�����#�`�mN�������ǖ���j�S՟T�k8�:��ַwY�nV�~ʎ/.�׷�5��[��x�g'�j:~��J����S�xg�r]S��~���o�����Dx4n:��cwy+�BF���oS�9;�vW��j+�,��Μ�z������r�e�Om��ח�q�WS��o�t`qTƵ��F���/6�4y�Z����3u4yS�Tr��_�v4t��x���^�R�4e����n���ȶ��p���= LC��D6�U��R�pP0y���G�5�G��և
�78d�<��^�}�Y>��q�{�٭�����Ƿ9��M�&�I]��[��L��[C�^����t�%~n-�w�:�_T��}Tv����%���7u��ճ���Z�X���z�dJ����m��"N҄�vg���Cv7�͛��1p��-�X^�$�W*T��-|���C�S�%{.J��DosqU�sy�&WJ��ѣ�� �#�N���7tmVT��UvȂ��@=�zbSw���]�ǟP�)�x�One�@-�y�0�l���S} �օ��A��N���Ⱥ3����,=��*��z��/�p��Ǘ]7V�z���Y��'S}�����+��\����9F��N��7��Û:7[����o��溹t��o�?z�@.>'����v|�4��w�:q���{\����8��{ǩ�n�8{D���r�ݏ6u��k>���x�ױ�˖�w]9���#c�wf�2�(<�����=l�3�����5+���`c<N��@'���ktnK�o4�K|+EIR�Zފ-�95�����i�{ر��h�N�o�<�-Rt*S�oG�VsOi̽�<Θ��;y����!����iX�.2u�;e>뇳������a\���m6P�>�k�_U�=�y�t����������7N�v]'��Ⱥ��D����^��w��>���9ՙX��zM�~��C-��/*�]B�k�r9A�_�'s��.j���h�b})����ڡ�}8�����h�5n[�7�J�3\���7ֶ��>�g��SEɯ��Q��o�vL�<i�0MZE��	.מ�r����8>�����xW�>�)V������}8`��'bxs��*K����P��`�j�hK�7�ֵ�UßmvKeA;WmoS�h�Z݂S���EO��R��A/<n{*�|�o(=����6\����(=Y�����y)s�oB�Bu9�O��^���T������~�.�o���<�zj�w=�O|&K��D�����M��ߓ~^���c2�K��Vpm��<r�
��K���_���	�^�������Qd(��w�V�Ԝ���a����,�[Q���[3��\�YJ��+�A��py�SQU9�35�˵�8PDPX���Zn�>_F������nAt݇��=���aj��x�Y>����������V5��F���͇7��pX��X�_}�{�}#�嶍��
�q�~�����y�*�S��|���\�4��v���ϻ�N�.ѹ��Yy�;������A��x�b���k>�<:����>��m��u��O��m�k>ֶ��Sl��^,�u�Nk\��9����M�q��F�뷕�G��cy񗁗i�k��އ#j����3������~Z���~rߢ���8��[�g�1^P�&>�j��ܞbo]�3�W}2�j����OP�L~__v=�7}��9c��yMٞ��G,����:�k��Oa�x%��^�~��L?%��
��� �E�c7���e甪�+���vP����	���㋂�+����wm�]Op���W����-mo\5/(s�!���qu�W���͛S��<������w�K2|=����1Vy��L	�Xw�����7��>f�ZчȰh��n�)	k��E��n��/V;�p���kz�I�s]�h�S�p�nD6�sn�d��u*V� �ܲ�����q�!�V�18�7���&�ڻU��{��EIxD+�B4�3�{T�Q�۞T��+.�=װ 7�lt�.�^�����fq�Y}��{����:��(�#����	�<�)�V�)�v�o�T�t��Y�ܪ��>�vi����tLU��W��U4'��U�0����:r�KK��ϕ�g�;ޔ����9B*���Q.�w^�����n�|�Bu�(�{�C����X�Ps(^z@
�t|��㍈gV��K��.�ە�zk��^)�~%'�Xt,���yѮO�>�z6���;�o�Y.���T7z�²v_�n��@2�q�So�~�=�v����t;{�c�3�f�����VOWu��7���{����nrϏbOm�Į{-�t��v�ѝo=2�~�g�qnf{��)t|�~�K�ϩH/�T^ug����V��D���_��~��g͇����#ܧ�]T�z�>.��'0���O^7��uNKHC=Z5��A�'z��4�����w���ӞԱIu���۬.�&5OsĐC&e<���Q�X�w0���9����I��ណ��K]�"�h�Rm�v���du�֌�s愫)*YW���ob�-`Jnv[&����̹QԺ{ӏ���Lf,�\cv�T�M�
�&�qZo#\!���7|4^�+�ԻXu2Q��1��zg|$�t{�����S�ǁ�ۓ����L�G�{=�)���5fOv���P�1���LN����zw�L���I^$P"�E�s}M��+��7Ӑ{=gވ��+jq��o�ຍT!��[j�=O�o����ɶ�R>�;Ͻ.;:8�����*�K\��[�̫S��+]�^��'�W���v%�)W)Ny����S���%�t�!�4�1���_:�t�9ao�	��N�=�#����GsH	���X�`�<��xg�_��}��j�����wֵZ�+19tzS�]�����J�'W��<c�^�R����h>�J�j[���c�7>�����D��~�+�5�	��J����̏.V�˭�j?sS�r����{jd���q2̺�ʩ]t�[��>�?SE-�U}�4�)�;�{�3���,��Ά��[�{/�&�Sa��'�fr�_wY���a�o��h����X����������n��z��ǽj�#��wb��{1�2H1����n@tVR��xKd�6���e�`����Տ+մ�y�ge��ՙ���H[��v�r��ԃ�	t�7����j��\[':���c>5}{��N��6DV:��rY�����hp%Aȡ���W8EG��Gvk��'����KN:6��oof���(��^F{�Ot�� ��vw1��� �i	�+.�2̝X��Òݲ�p���z���Oԓ{U]t\h{H��X��m�÷�2F�U�+�sS ���'G^˒�Ot9׺�7�uz�~o4�f3�#���ݖ tg�ܮ=����7������+hLͺ6KR�*�f�R�9�>�Ȝ�1r�v�[%��Uf��%wM3����;|� �+x;;V='�	鲷��X��ϲ�eJ��8�������WI-nPG�4�S:c�`��ŋ�hMv��Ms�i3��|E�;�ٗ��(�&zj	�a%���^��E�td���Y�K���F�P�슇K[�<��ʙ��d�>��a��������[u�1���gc:,��}�,ρH�W�8ep��.u�F��B�f�)���ϳ���j8���?%Y������=Yx���8�K$U�3�����b��>Dyz)��ۋϵ��f��Y�imM�bK�E[Ã����Iؔ�s7�k�s��t`TX��|q8b��hXƫ5����rpp�?8�b ���f�c��,�}f�t%������c'���n��s3SĢ��3�4蘵�sŭ5'�D����k�k�L��[�i��j����rK��%�a�9������Z�9.ِ	bkr��,Ӛc,�ͩ)��^�!��6|�e`�Ѧ�>�eH���T�r�dh�z��I<��f=���N��}�����^l�ŝ�	��tk�m,
IK��sY�R���ESx�\��΋P��ِ���B�+�/=��ikr��e"S�0�;���sSߗ�6n����󕏏�-�L���7/*W�e�*���,l���A��y7�5Ã�6�L)�ʊP�z)&�M�D��R�k�0���Φ4m�Ow�Y	%��R�2�۱;Q�uƦ��_�<8V\�@�#ZߦEBU]x�~Ev]�-��
���S��%�;Kj�;�Y�L�r@s��� ��c;XOu�ٿ?�5k�d{�9]Ϳ��t�Ʈ�=kz���<��z=݆`Շ�y�����mcUcg7���:��^g3Dh��߮�T9���:��y��;����X۱2e���c�_���	�h��w���_wW.V��0��DQn�a^{��ݔ0���/%ɡ��r�2������l�`�����p�u��9��.���e�9c]���e �/*��@ %�7uc�{�s����W�Ӑ����Dl�L�;�ʺ�f�:+�rEw�Y��VO���	��Ӕ��\��V�P��uq��Uo�Mkw��g����!��U���*�&�m�h��ʐ�h�AF�Qb�V�R�V(�X���()Z��&�Qqa��U+
$�n.	iQ[l`�Aj)+*�X�R��eB�m�ZUJ�PF�Z�V�U��T�**�U����E��*�J��0�W��Z�QJ�J�Y����j�P��[kYX�6�q����K0��L[%�cVʴ��dPqe`���E��mXV��E�E
���**�R�Z6�B���V��++�10ʕ�.(aqbԨ�T�E+��Z�#�
4�m����*�*VV6���-fR�[*�J�l����V��XE����`��Q�J\bB�ŕ��D
$Z�F�l6�Ŗ�ذ����`�mX�+��$��M�(��&5΁��`�ގ)�wP���9D(-�e	����ή��̀�*�/Pf����|����I����9�����f�zw��rM����w,�+�a�S��)iۨ�f�wA��_w�GF6�����+d�֗�;w�i��}u���=�Y�'f]^�4��+�9�S}J���λ �����xޠ�3�u�XZ�x�?-7��~~��*�|�}7�M�$�$b�k����������8M��3��5�%��)��=k��:q[���}w���]^��{f�t�u�A�~�����V.��ӽo�k	
�	�ێ�ߚV�Uo>ܪ���S�O�C>��.��8�+r-#Tױ`��߫�B^���M�}5lP?m�&v�wezj/Vh*oL�����#���*�5���'-�����ߦ�;r�:x)�R���ɕ䉽>��z����
�W�V;�����0n�7[��p����z_��vE�r���s,cv��{ʥo,h�u��0k[��c쯆��ӄ;.�⏲�����|�{Y����oU�z���;�j���4f*l������72�Z���^yf�F��Ƚ�؇DK������E�};;�V�W���'&q����.	��$�d�'_y��M��՝R�>��x��U����^�\���ٴ#��~�Y���ͣ\G�u��&*�^��\E]/DN�:��{
�1t�u6���צg Ulj��pi�g����$�v�˳�ȯ5�[���O� 5]�.��n{���8\��r�N<��������{���x�+�	SӖ��>����ם�:�sa���4��*�!�~�D��2��~���^�eN���e\\m�V���>�y[����ޞv�l�=��dK�&�W�yk��^u�ܡ����|���\�U�sF����lV�=˟d�o�rN~�S����r��o>2��V���=g7l��͵�]S�'g��M�O<�~r꟢��ӈ�E�hA��鈭=�f��>�]��Ǧm}m���x�y'6w��9���^�6�y�,����,�p}���;����G{�Il=ǫ��i�4�>�vޝn�;Xg^;E��:</�Y���hb�v����G�<�gc~��*���\�Ӟ���|�{/�}=��1M�MŜ$�ۢ�L��P�nWi}�}�pm
�u �s�/_���K�ΐ��U~^9����W~w�O/�O?G����� V�:k�N7;��y�+���ϥ0�
�7��-|J�1G��%���5�1ێ�o��s[V�[�]���I瑨�8玵�A��D㶭�C���\��0�v�R��S�]y����+����Բ*lfJkЯw�W�������2��|%t�(��J�H��	�@�:o��ۜ��"ͬ~��U�2xM�(sҙZ�{�]�=^A��'*;���^��c���!�~純�����k�����#/ꕑ}@{���`�>����Oq6'�����X� ��i{0j�t~򓅾�LE������ �x�-ݒ���w��5������R%�T�s=<yȯ��3Ǎz-��<�ьҜ�U9v���2��sp�5��Pmޯ$��H`���Q1�AWK�g'��N�P{��5���Û��B��Kg��8%=y�Ag:��to#}��_\u���/Glf����Z�GRws�59g���SB�Q�C�\��!���C�K�J�o>.�R��-�A>�Ó����O|�z\;�z�ͺ�:��~ߍ��`��y��L���jB��|fi�}�q��es�n��|�>�ԣ#W��mM=*{o����� nU��".�9��=������:��L�귱�����̾a9����*���9��/��ֱ��zڭn��/}����@_�<j��K�t���]�W�:�>t���b��X�>ʫ��h�����~p�x�'���};�]S�M��vgR���zv���C6��Jn2cxm�o����M��I8����ƥ�k�{Qx_\�����'o>�����;�u�~�>�����JtzKv�pFz��I]^ީ�yD�1+����gf�W]�����Q[����}=BCH`� ���׼�=�{"	�bߧ��Fk �&�b��MzW� 'O���`�4�T��9�����"\9�/m��(��iD�p�Ċ}���)�IENL��g��#��yz"���a����"��#�ʎ��Ή� �P�*>�Ȗ��81d���� �z$�y ����N��u�tJ�tXOM,�u�C�+�b���KjGޱ:�y������� �%��9�gj*թΓ}w�P����R�l��K���`iŭ|��1zh��Z�Ea+�աf�R��]S#��P��ۛ����T&�*S�\��ݵu�~v�c��Ԫd?xp�U3��9z$Vӗhz��,h��ٝ^|:���K�U�����-�}Ώ�A��}��R<��;�Z[{'F�����<5�	��&�w����G��97���~� ���<�	''u��z�L���/�b.����.WJm�{A�s���:��e�n�w����=Ow���##��?z�������o9�1�R��K�Na�=:h�ƯM�}��E�z}�x7N�v]Q�"WS����)����F�g��$۷�oʫ9��׌�����OE7B�O�����Ϳlg�Mv3����c�g�{��:U�k��ڽ��n��
hp��W&W��7<&H�������A؞
����=�E^����wi�gY!�KW+�Dէ���2��2�k��d�v���iĸ�WW2�y���:��F����%m=ᛙ8k��H�E�I���WX�>[��j���=����͡�Dd� Q�A���I��X޼��O��*��5��޳�/�� ��UΫ��+�O�t�ԭ�����1����{[=/����-��]y���D����>�S��r��}A�}Uk^���myc���;�)Ӄ���(�\��J�(��CY��������W�	�7�,��t���E#�I�k�`SJ���"�*r�^��/}�%}��
�Os�2����˞~cq6�t9&�nd ��quܾ!�dW��f�>��=��*��V��cy����A`z|:I��l߰+ܭ�����hH|6exp�����Ϛ����>�X�殉�y��9�_� w>�_���I���|�����:��Fo+{%�Ph�<�?S��l�͡��,{U~�9��l�R�ۙ�(_�_uv9�T+F���:�ƂrN�T��V7^8�51���P]Y�|m����'�]9����
��w4Sم�}���z%vu#+���.��;�K��Ss��v����t��B�{݇��,6��ͷY//�YZK;Ϲ�ݣ�3��ډ��vt���u懺5�g�R�L�J�hz���N]j�n6�8�����|�{w�e��~��̹���\����PyV�ŀk�s��}�����/�oX���n�Ӟ�qM��퓈���g�"n{y�a�q2����ה<��d�~T��{�_G�Ν.�^������2�r�=��S�{(O3]�(S)pګ�U�{U�;+ѝ�9�����9�V��ns�8�	��\�o;3�}^:���:��K ��-��e=�"�_G;�؞^w�o����+Q}�5WAQ�������φ�~e}���K��P!=���̻�{Cs:���F%Ӕ~[�LF���A��x�`��X���{�i��|�w�����K��/�/�C��yYh��>��_��4f��ߊ�ް6�K�^/���	W:�f�O��DZ��{���x��^��'�������v��=v�g!�߱��
������׆��>��~|��pēK ��9��B�[
���P6�9�$-q�����;-dlo��e�Zf�ӱ�>�G7z�a� �v2��n�:��#�\�[���)u�b����1�C˚-��!���^�a�e+9�bd�k�
�L_uڇ*6s�\=ie�~u�s�wI�֪T����ay�Ká'��R5c�P��:6����xl��k�Ͻۗj�"t<>�g+�R��7��`�hpe����5L�l�-a�s8L�>����g^��P�ks�ך���jz�Q�T�#mS�F����xf�b-�Oحz�FS]�n�;>�V��c�u/��Sy1bd�����O�T^ҕ�n�Ś7���튧=�����8���.��H���B�z�}l&f��S<:+���V�=kW��!(A�`�{i,���N��A��C���3�1�;ǆq��$m{+k��v��L�Y�����?���P:��{2�ڜ����kr�����s}|/Q�'��2�^����F痃�ʑAg��xhk��� x���0.���R��=ʟv	�H�g�w0�[�^�7��I�ji�¾�맟KB�d ?)����,ND��]zgL�����gG�t;I�&)P��MǪ@w��/�E��9�������yץ9M�W7���|�V�xڡ�k񖝿+K;x|u ��f���}j�I2�bxlhE>{q�"��e�Ҭ[��l�k��/m��Z'x×k���)�2�+J��s�vՕ��ɘ)8����P��+��3�����]�����-p��n�t��D�9u��ML4z��'����wu��u��vEa�̖�Vۼ�\�T]L��xR�_��`���ȫٷq�g�z� �^Dko���!���>����|Ou�_t��Wngeо'-Դd�C�ss�%=V�g�CȇY�h[�h2j#�CC���W�Z����
�u���<��՗�f���t�{�Y��>�6x졾���k�7���N4��ֳ5��IAc<t���x� U�	�g²�$a��3�S��ޗ�;�ˠ��هP,ws�l�mʍ�R[�7B�A�LR�P��G�"q�K���ì?	�V����TGyMĜ��^�J���S+�-U���(Q|�ؽ1�p�Ut��n;���A��nJ\���^�ܖ��ʀٕW���5�
�1K-{LK�PX��ج����~-���c��l��� T�A@Ԛ��Ǥm�2]m��2�Y�4�6"D�\?d�sמ�vv:2r�U��
F�ڙ&��<*�=^���r=�~HA{�`?��
1�:U���fc�h������K+[Z�4���w�i�Pɔ�c5�tl�"��ȠR.VR��B��_<!ͮ�o&�������e�[��Z'�=����.�V&��X�#�MX5���^	�l�)�V:�]�
{�Z�l��?tǯ_NF��@�Qw�����:0�)RkYA���B[�xd�z~\f:p�KW��zL��Q�3W�ݕzO������`<]٣�M��#Y�����'�"�k��C����iދ��)�_��s�2�u~��	���<�a.�����2��R�����9��w�vk�y��Wl�G{{<],�m?��Na�r�{�>��j��g5�`����Yc���Y�M46��ÝMz��ΞJ�OB�b��$y��޴/�}=������U��kt��>W �j䛑Ή��.�2��&�� �K��R���ދ�9J��)m���L�o<XD�Sbk��~�`??�wD�L�Z�z�ϫ�:
�� ���#�U���ϔ�SM��k�5�<�u�/�"���KZ7ٵ��;)+�4!��"��QPUʡ$.��J���R�����g�Sk�ubY���"!��3��p���^�<]֎�O�Iŝ��ܬ�B^���m� �c�y|�YjWfk2�O&l�}�����7��^�����ߣ����-���}��^YS���c�n�Ñ���<}��%������$h�����A��ti�t�c3�;�ϲ���68"-�+�$�<�������\�'�zz(�izo��Fs!��w��D�x#.��.������Sj�b�ף��|��h�c��7�l��=�-�3x7'S���G�R�x4��sҴ�k����ǝ��E��3<�Dy����l\��;c�vX�49ط������9�:}kpe��)ӝN����A�m��5�X�ns�$֔;ѩ���Ȱ.��{��kA�E��k9�M�eN�n�Z�Va��i��:!§>V�*�q�����.��s�h&��G�zm
����|I��LEx��Q���m�� �GbIq�؁��k����p���y���Q>#5*��i�G��JVxl³���jǴe�%�I �ę��{]*V�R=B����;]9ь����i��7L��+l�ws�qn�ͳݥ5܄���$�#�\���u�;��BY�^3���;�\E�Ǎ6�>���Ir�{<�y��Muّ&>������;�[9� �M�{Y�6��$���b���ȯ�C��T1>��� 扮��{V9�Z�P�e���h��7�d���s�f�5yb�f�I(��i\'��iQ�ԕ�44j��t�&bRWk�=K��█�S�w�HpA�n�%��P�m"�)L9f�e`�ݢ�d�f@��a%��Y�e<���N�ip@��-�*�.��Z��Or|�B�c�6�H˦a����J�,	*&#�LړNV�RL������mVP͘5��Ph3l/��c(�3vӊH�$������Nl�5Ddˑc�.&T5TO�Jv�ѹ6�%*��(iuu/+�,�q�RP?p���!�����ܻ���6�C�H3n�]�V��Dx�l"�*�5+n�%��dww\�Q�/�����o#-��.��R��P�n�*3)�`o���*V���i���G���˺0���YE�5v�N�Z��Æ�?;n;�w;5���
&�ݱj�mA~D��e��b1T��V�!$�SU��	�+�nXN��wFF̭�*9+8Jh�L_Z�Q��&�İ�6T�z�neȖ@��j)&k5B��Լ�1�m�S/�Xr�]�R���u���5��{����E$
�Rک�+�V# �e���jQ�-Z�cj0D*�Z���j�[eF�*�%IP�jTQ�Z��R��j���PkEV��TFT-�ef�QlTZƴD��dQ�����c0V���J����-��E��\S����YR�V�E+V�YQKKR�P[aUJ%VVKikh�"��ړ	TEX�
8�m�E�(� �R�ڪ[Jƶ6ʔQ�Z����qEkhƶ��֋Q�����FжرPQL[0�Zb� �*QZ���Åp��b�*#KL$�����*V��+m%T0�1-҅R�+Qb+P�Z��DU�Pb��)akDT��UV��,�6��m�����."�bZ[h�(�ʂ#lX"-dJ�TDiJ�VV��X-�F��"�2ڌUe�Ҋ)U����ʃ����0�F�~�(Z��\x�L��*�.��;��";�)k9������J��]����qV7�9��<���y0
w�l��1��W^V��{����޴.۷�ck2Y]m�/�a��E1	���a�,[q�Y�ŃԻU*�m׻IU��}D�8o�BMד}�y \>i||��5�e�{�>�N�6�A����I�$!]�� ��m]p�<��s�
5��5f�В�Ϭ���a�aܳrΩ&�H�N`o�F���d5�3�{�(�,��	�{���^d�п��̜���W1}����~�Yz"a��&�߳��}��2�EO{7���(gz�wTxAw\�5K)���h�����L�4��g_U� ��o��2t({:��&ݨt!�MT�k�0T�c:��36�C�{�.LK����=[o��F��rt;)G��J+�v�+�0�ڬ�(1�k�ul���^�e��~�qee�>~���y
޽�1�/�8m+���;�%K}~xLֈ������p�MT�ݓ���,`�^5b��@1c6n�����B�Co�׎�=U�C\��2�����=�'QZ���k#���T��f �|p=��C��ё�\��=m�{���IS�R��H��aWW!BI;�_%k~���4�z�������`H�v�&.�uт���񑕁�Z�c�W3jL�r¿��Fz�y����^ڎ^N�mm��Q�8v���t7��`��@@�]�;�W����뷆�d�ߙ��6���[�D�XD��d�YL�
�]L�M�a����d�bΩ͙-��r��a���^;���w+�.���FQ0U:e���5B)[��;�a)�ܛJ���g��n����>�鋅�������p�Ǩ��['Z���Ǥ�_D��=U��S�o��jPcUb
t������Ĕ�}�+Z��#�Mj��ܓ3Ԍ����, }EX�H-r�/>�����Z�JF�������ubܕ��Xy�;�7�x�d�ϼV���pP�Ju�)^|��#>p�=q��S�*@��pv��A���m�T��WT�:%W��xR�(
w�(8s�*���e~Q�=0���k
)P��SM�ќ=�yT�`mr|`Xjo+���/�8e7Mh�1����>�)�\�O���=�ߔ^���D�r��`Nڙb���O{_+����5�s�s��6@;1�����6˸��p����/[髥Ｕ7) �XسZ��.j�-s����8�N xp�e2������ʾ�H�Fl��n����Zt�X�Y�f���<i�?"���\]7�}�g��Ӹ���>��T�U\�:fmޛ2��xxpB��V�V3W�U�<�����������Z�λ�OҺ�zs��>�^�*��#�Obw�=ư])n��E�',OF�������Ҳ��i���}ω������������q�9h!`�]V�V�r����U�*\��:A�K~�e#J��D�=Z�3Z4;*���W�C�=��ꗶ���E3Һ�9�ݿn<�]>>�i3c+6>1Qbu߂R�3�=�u�.�S��5�S���u�Qa�������R38��@�c�DJշ,���:<���3��O`�䮥K�g�9��\������L���-{hg�*��eqh��+��BLT�gd��MZKձ�1�V`�|�s`{[>;(yA޺��BdP6j�Ӻ5���*�d�M��Q@��_tkv���@ޔ *���>�v��FQ(s9K��JW��#j�#�y)=�e�9m���4s����
��@��
�PH	BBE],��(��q/^����16 x��'�޳ʣ^��r#u%W���6�\�g*��Qr���9������ ��_]B#k���m(ԀQ;AU��xH���:�b���^͞Y/|��}BV���2k�k��r����=�;�ܙ���Ax뎱9�f*��䤊gnj�Щ�nV�#8f���'����U3�-S&(�B�*�V4Fb��|+8���vJX��o��d����2�M�+ӟV�drϺ�	��f3�vњlO\�+Rv ��>bn�I莎����\�@צ��G�d]-u`O�����Y�/O{2'�i�V�i�s�����^<��[�r���SRm�ѽ��yX�P�_6��D�Kp��m&m�X��bc}�y�>;q�Xo�Uxm�	w/&h�.���抩�c�	�z8;}��r^�3�8w�^��ߗc����=�G��3ġ�\#�S�+oH�{���[(A��/�������!ѕ3V��ePs��,t$�\�k�O<����^��;�C���VD�V''lxz��7+Ub���*���]r\�{�~䤫��^iD���`A<*ikK��e���u�t��߄~��=W[W��ܙ����} �V���ѯk��E@gq���.��&sYUf�*��w�K����i�吴�!�I�F������E"���6՗i[�\�C�_׸y� ."j��g�7쾩�:�{�<��@��'�\镱�Js��gY&-�ͧĻ����t�CсO��,W��N�2�s�ǖ�-��63�v��ھi��?0멓 ��K|����Ui��\-�au���*�L��[V��xw.4�5��'���(�-��GR�(�� :\�ߙ���k��r���w�t�{�t������=�����g$yb�pJ�5k�mg��	(l ���<)���;���/7J����7��x���d�X_W���#YD�%EC�BH~۬�Cte�>�=/�Cs��^����Z�	U����'2
�����0���"�0�uQ ��G0V"�ؑ|b�����Z&�����7���s~ ��r C*�0��]�^��@g؀�Uׇ�W3u7�}w�� ����zE�~��n�:Y%��H�K�o¢���+�P�+��{YOJ��'-:�2���f���!��U�s��;����j>������/�4�]	���,��_dJػ�2�������$P��9����^�����]�<��wf�Ju~��y���n��G{k��CTtAw��T�����9���.D�dh��n�Z�'�k�w�l���G�0�j7�l���s\�x��)	q��־�i�8i�n�V�7�|GF����A��R�B�����^�U/s6���z��;�ٜ�'X˦�ɹ���y�Ӕ�gz���I/��z 5�G�\�A�e]��#͝:���M�i�=B\��!TL��L�}H�q/ab���3*�o�c�__>J����f�ϫ�2~CMX�f�ы>M:>M�n(� �h�H��ł��d���0ۗ،Ϻ�z��VB�����3���4SdB�~�����ϼ��(�N�ˢ�s0|��;ݭ[�*M�}�g_`7�~=<����V=U�=/ᢛ&rk��4-��C����4��^�kjƮ̶��_��*i>�e�3u���e�@@�������<���~�T\�Õ�aC�x_��#�^�.��!�>fPUW��gޛ�G�>�^�s��K=�syپ�Q�t�]tE�C����]�6��mS��.�Z�Ѐ�(w��<jW��[p{b��i��gk4=͟TJ�(�"a�,Z7����Uz#f�����	�=�.J첟�\k�5Gw��h�̣�RI�>��V��t`�S�*�U�d�k�
����{͉���#Ǿ~@r�s0}uqV�k��^�:yh���2�?}\X��^�5{�6���n*��Ζ�t3�V���1�ߠE�{��	�������	�@�{��yl-�5J�����1;���{�+���]˹ؾ�^7�{��)J\e<�V�\3(�oO�9���i�@v���%��vOyU������K��Zsٞ��\���b��V_���D�N�ߜ�g��+f5�kg�/<Oz�I&���.��k�<Y9>�U�ߏ ��e�52.8}-QZ�j�Viя��#���:������}����y������u�Qv�E�Y�ܯ�pK�d���]5V=(��">M���`�6��E�Kկb�m�7Y) �uدC\��N������ٿe������� �30ւ��U���ɔ�����ZRC�z�b��U`'xy޳�(� �S��$~�XX�i�a�3���3�x�24�����q���ho�g��P#!u�n�X��e���۱�k�ۧ�5�d�X7���}F,�v�_E�4�$�Q��鲦^Vt��rf�(O>�c!JC~�z��t{>��!8և�;����vX�'�0�I{^��nyw���]�i�f���Y�po6�-�j� ���?J��'�i������K��u����R� ��+|̡`q�V3�x=�XU�J���lOCֽ+��TZ��0R��)����݋o�i���T���h�����x)�R��=t�y�*�ԝ/�I����֍�9�WA�O�g���^�kì�yu�W��G}�5Ӷ���f�L������l�/���{rn^��Nv��&Md�Ϫo�G��:��Z�v��.M�n�1�M3}K��ֹ������Mz�v�\,S��$8�ve��ab*�.�P�� u����A�����8���ЧAk�C*%Q����R�ZW�{��ؕ�n���tL��1B�X�9C2�sg���z�9��q�P�q�(ֳmPۣ������h��+��@s�* ��U�&P����%cׇ̘Rޞ�ٰ�T�m@�;vW�M��t�#��ۖ.�5(A�4���
���*�Y�QKЎ�iΨ��f�s���8n�_��������]L�H�WM)-`��˱u�B�
ua����0��>�P:�s�F�,�x�'�KyDn;�c,a߫d�9g[�*��a�>�]�f�˽�˓���U�W{M���&��i���[�מ��e.�{S� 'W~0��`;���s���S��-�>�jN���G	�u�ulyp�HY�S*Eg�}�u�իN���c�}-��\P��QA�������,7�*�6�K�����4�#+m��D��A���ɣ���>�/�M�V�縜��뼸zGhvGh�.�0�+3��4ѯ%���K����Q��_;Y@侤yӐ��o���+�"��{+K|�h�ݞ�o�:�V�h WLw�: cw?eڱ�5X���Ưz��+�/L�-��4O�^X:��yY�j�胙��NftYŎ����b��T�����ϗ<є��g���N2��Ո�g[�L���t]C�^��[&L�Ǯ9���\w�D���G8�=C�u��Ŏq"��낶����k5z-�V�bp���u9�=nW��]e�GkC˶+��.F�v�U:{h�e �t�a3�t����h1�7�e��%�/�p*xXw���b�b���F�Q�-�C+�<�\Y�y�>�8��xKap��z��^�S�k������ ���wr�|����>>���B��^�I\ݷ�7X��q���V��=1E�D�U#(h�@��=�dAR�t����K_�M����������ҙ���%�C����^��>P�8�E��.T�
�4��G�]�v��tI��Y�A�QWL�T��<&���U�.��XƑ���jT� �Y�t���8�u�.��C9�сx�ܧ6�5�]v@��� �<�����f��r�ځ��a�z&��	\��M��2����m��,������K	�vn_�m�Tݿ:T/Uc��'��
ew!��r_K��!�{�{mk��:��Whc͙�:S���PfpekQ����CM�Z�e>���١k�tC����ˈ�5�[r�k��縖𲟏�'�۩u	N;ў���D�č�6�*ml��o�(l*��b.-%��dr��[�Bn ;��ؔ�YU=ҟz�1w��l�%Wr��e�/5k�ݻ����]zhSÎAѾU�u�&��3TG*��P���7\��>EtN��ǃ��p��4]و�s���}�����R��������{��U�A��y��֯hSڽ�v�	��7:q�S�Z��>Z����%�є����҇���맭1cj����37T����.M��R��K�P��
Nzы'A�o+r�W�O-�����>x��]ʲ۵pmt���7����J�#v�O�y���0g��+E6x��c����ݡ>;��]��N���[�����΂g��1K�>N��l��s���]���WO����2�m�qZ�>p͈{7����;ͯv+L�v�:<����̎���pu\P�w���"����j}������oW�V�f��,O�i�pOwyj��+��9�#) ~�[�=�>�;J��e'��kfU�J����C�w�(�g��q�cw.�F��J�+�D�����'s�{�XB����5��Y���/���Rޱ{�Q�헲�-G9���wS��!�ÁY��3�.�|%�Z��U��(' �u�q���C�|f�+w�Nz;Uv>����܂��n���y���{'�'��/{<�;,��]�9�WO�FZ�zd� ��UV�f�:��r޼BY)�Łu;��x/f�c
��GU�ؘ�.nOn��N�u���ð����:è{���CD�������M�e�_����|�_(;�kx�6�Zi8e^V���X�نG>̾��%�ز6�787sB�%G��!a�^���u�a?v�.�.������T���:��hz���W�"�#�Ps��zo�w�����E�=��=��/;� �Š�
����w�G��զ�(4+;{�q)�7��b�P�>ɧv��$�W�i��e��1��3J�\����-�r�p9>3B���6vsԱ��
C�r�|ēT�τ��[�{sJJ��j*�o��[$s ��ڣ�'3:�U�u�T���1U���9Z���1q֨G&lJt��ZY۲�o'5���%���%��\���9{�+9�K2s�9��3R���[���;vX{d�^L[�M�U�}���i�¨*�|*G���*�sGi:f/���W����|kY\,w,R���6�R�sr��Z;jnX��Ľ.5R���bp�]����H��h����WV����sr��`��xk2�#��r���h�v���/Q�lP�<�6�k��S�Od�u�epڊ�Nͣ��a�z$�ypq#�^֖�}ï�~1�Kw,�v*��.bZ�-�9��f��p�OIN��	_ ���}���)���!N^��ULR1e�w��:e!��7r�p.*\j��/w;8M�p���R&M,P,��Į'��Ds/.vnG:�Kh�%5U�Z�@hx��;�]��ruou���Gpg��ʵ2�9)&e��2"Or��G3e���Lqe����Ԓ땚4�w���1�z������; �&���f��(���S
�c��w���F����R�J�NUȨ;ױ^�V0�>��WH�Rʨn3R-���w`*�"�ŋ�rl�u�˸��㕫^���!,��ٿz���.>���7�ӎ ��j�����C�Oo̮����,���6�fUFd n�n���r�0�����W2��t}�.�a�YĦ���!ac�l�՘�h���c����մ2���s�gg�8�*��31���g���w�B���6I�n̛j|!��>�u�o:=�?�9�:�.���Z�zd�?X8
�&8����f���,���6^vQ�V��Ğh>�mۼ0]↥�А/d&�����+<�\�bJ%A�K7:W>�gw%�y��qJ3�
��e���|������G��>ŻDؐ��O%�/̣�/в#<X|���$|�h>���d{��3o�Om�e�lo�/�����ՊJҒ*��Ō�sH��}n۫�ί^�)�f��䊬{q��o�z�7����롔~&��
� UE-�ʕeUPc%���QX�DF���TQKJ"(�m��E1d��"�؈�Qj""Q(�J��Ƶ[B�*
KUa-�	iQ1
ű�Klm
�p�qh֠��[E��щ*V[LZ���Ke����k*�A1U���XŋjJ�V��R�J�*,b2�J�AX(�a�ŢV��*V��QDjڡQ�ֱ�m
�)qq0�����[U����(�,R5��m�A��j)YR��*��*����Z�F�7-UQQ��[�X�JZ�%ej��iF�؈5��J�JkA[Z�H�F�maR��50bK�D��"1X��%���)UDE"[0�Q�֥cR�1�X�jUKJ�Lc���-��"UJ5
�%�ab,T�-�U��
�U�*��V�P��Ա�J��)V��kF�±U%�cR��TB��~ Dgw.�7-�喰줜�� sI����W=��{}��m�Z=�Yof�k���fr����ܜ�4�w+���FM�,�3�c�A���xq�����5+��1t3����k�xgܕo� ��<u=Au��5BW�:]�g��D)ҋ�X���D�u��(u�ބ`�f7�:Uוk��C�e`'�ד� 
��K)ݟr�[��b��Θ��Q��o.j�����3����pʜ�2��]������^�:���2��kE���v|nvt��=�s�z	S��AP�������0*��9^�J�9N`���:��FN���a9��@kܧ����Zγ=F��V��i88�}(:�^�]qA�YSE�H�uP�Ӄ�W�mՇ��o��ޠ�̀Ġ�#j�<^�Z9S���`�`o*z`Y�����۝�����2���Z�$�4{�F���<��y�~�6n�!w�)�h�2�L�f�7sg^JQ�%p��٥W�v����xVlِpϴ���1V/~�Wm[V�j���Oe������{OT��j��[/��x?���uS�h�<��ώ�P:^}wB��f�wL�{��0t'Rj�N����Md��dw��M�F��
rr�x*�`|gF�mӰ	��2����%�q$ҵ�wSl<v;z����	����I-w�hf���z������'����'�f���#�M+a��%*��b��veO���Sz�y��\�p�a��K4�l��+M>;���;�(δ�T,��� ��X&F�n?y�E����w��b`K��+Z�cN�	}"��c����h�e8��K~���M�w!YHS}�[֝�K2Mw�G����Ү�3ʶ2b,�g�x����4xm��3*wi�/�]�樽�7��}�xj}�Rp��Ž���ym�87	���V3�Sx=�,'X�=�6�vI/�M���Β�,�sf�؍[fA� 9�����-�U��������L�n;��_���է��x��/�b�s~�	Z����{h��Aǌ{g�0��:f��2��/���:�Hΰ������:aP $t5]�h�E��׵���oV=���]Eh[����I[��m螑�!gE�
��J>7U�R��ɁJ�BBE],����[�,v���>'��U�:��R�>0Wy*����QE�
!�u.ś�ևf�
S�A�wW�U�ۖu�bX:���Id�ϫ�5b�fi4bƫw�xϝ`��B�1�^^�:?�]�����+�,c�eN�UB�u���Ƿ �,.��z��`�y<}��A�u�c��ػW���	_=�#��c�ڬȯ��<9�{]�$������i����Ѕ�]9�@��-�&M�N�y�-�i�vA�������.����I���Cp0�Q�q9�>3��O9.�U٬�;\�Z��]q����p�}�K������v�����l�Cl��7���t��ӷ}^���o%l���U5�K��#�̂}��#ڢ����)�^>Q�ݙk��˛5=���k�/NL-����{�7EGuћ���{$x���-���W�p��,��zg3�����R���E�D=>�Ps���RZ��`ߡp��<�_ö׎�����ʺ^�`�jXY!��9��8}�*]��EB#���sg��c�����y�_�o'��Ƿ��K���*�~�9�&&��]sH/L,f�}�Jǝ��A[�\�<���Q�|F��r����]�cFzmw/LB�T�����-f�Nѐ{P����fHn6;k�!�V���k��Z,U���`�G3�je�\�ڻ�K��N� �v��R^΍�v�B���^�U/�tK�̪U �K��R�|��Y��z��;�X�]ƶ��W!�bx���[�+l-Ł�g��'M��z��Xq@��V�R�ڟm����3�m"�R�^�{F�v�/����L[7w�*�Tܳ��sgm�����3���y�}+),���3k`Ճ�(�Ar�+*�8^kg�v��g�a��`����5R���i��(��e�Q2���@�f�ˌ.�ݚ`�#����b!
�f	��P��y��وL��]�TQ�D�B��-��{C���4�ѕ�\�B�GڡM��,�����ڮ6?����`Ƒ6/��4�<�U�廌�Վ�'=Q!�ipa�W��R��'D�S�������]�&��]��׫�	M-fD�3�M��Ft�6V��y�"ǆ�X+�j��YS%�'6����X@PS�t��T���,ܳԧ-��F�[�.��e��.�����ǜ��_9�޼�Y������V�;�q�ʽ�턮5FM_=�Y�;�a��	�����Ѕے��3��{�"�z�QR)��!�����^|�5K��)��겮�\qn��7C��fV\�~0��þ
�A5��U6�Y�>oȇ��l`�8���%���r5*K�gg��˷�X�z�봘y4�q�u��� )���2ȃ<X��t�>vwQ�oh��v�L��i�����JX��3������&���3a�`\هOu���j�H������c��W��Ɗ�L?�����8݁E3���a1ǹ�ڭ^��	O��s��7�������ϣS�+��/ow�=�\��U��*D���;u�3Q|m���i�f&�ݔ�l{~n�W�yv�}�ǐo��{t[��}���W���s_��矙�^]� _��SWw{��GZ�s�U���݀����aN+��V��Ʒ��*�h�Ji>ߩWB���B�f�h@FF[�ǁŸ'��Q��~�څ����e���]%��ɃLX̠��Լgӆ�M��y���gi�0�}�@w�|c���^���P�Ykh>���L�/��NK{��ȧ��^���[~�l	޺'-P�v.C�b�a�bk�c!�Ltz���[��ձ��׹a���i�{�
v:P ��L���Y�e�o�����a#ĕI��Qf�v������L���_ܑ�t� Ȉ�G���u��.���y.�	���wby�]��y��p���S�����^�P3��&Y�,�L�o � ��9�sK��V�w�XP�1�#��;�H���o(]����>��+�Fp��7^ޤ=�ǳ:���G�4�핯�|��h1��u�|uVs��*�jX���q�k�L]�*����-۫Ӛ\�ɞ��� �3ÚiY}�=���}�ݥ���d9�0R�W7�Ǣ:�k�$v�o_[�> ݐ�E͹ڛt��;Δ�@'�V�ϱ��i�2��R��)�:��;�XpKo�]�4*�M�ܹ�g��ӂ�~��QC����iLݺn�&��j��`yqs��Wic�0�e	�#j�<^�v��=f�S2�[��OL(�圣d�r��q�����>.�X�g�YZ�gϲM,]O7��W�U����}srac<���7�oWYs��9{B��vxA)ye�4gx��#����9�G�o�O��&�9�{�Ð`�.���\�{��|�����<rD���E<��kҗ�h��{ݨF�
g��ܶ7����~(jUgm��.��XjC��\'�|�3�3�3�P�DV��Ru-�����^�׭tX��y`r�ś��ڬ8&}�/Z�:
�Z"��m-�L��f��ϰ��l�	���kEۻ��ϙ5_'�=�j���e�^���_��Z�2������e9S�;/��2������yy.��C���8G�;o�f;�4�Rr�7�G�^���y׽׷���W����My3.*/��84��lF�*˛��&�J��o��b�qޠ۩�|��x��P��������<��Y͔����l�41�#�w^��:����C�i_>EFwkkF��.u���ƟZ�Q����y���`�5�=�y�{u³��-���\���Jt�M����MJ�[f�§f͘�� J��".��vѼ���3��Yѓ�䇹���Q�O���;[Id��{�f�~�?J�5w��	}��k7������g!��x���m_������	*��]$�q%�ߩ�_ �*�c���ok�o�3�#���2�<(3Q^�X-;L��e�{��<�Պ�M�;°���\��&�h��J�r�b�)ޥ���p�(�h�~sRb����}�H���1�~Lg�T�g%���p�����>�2�O�o�`�e���#ak� ���
#*��׳k1�)De����ݙ�ң'{�l`~�`8X��j쪗��r�屚��X1�`�<ބ=���<\�>_�f�`�4����81�tP�Z�����?L�|�q-?HUS���;L��-�5=�ٲ��W�����& /7���X�������f}�t^U����QX��qQ��}JE(��噗��N_��s��o�hH������̛λ,�������:�}Lngӕ�*�t��f�s���G}��ѥZX�%	�BXf'}� �x��z���fr��8��{f�yg)6tY��Ŋ38C�Hc�u�N|�m�ئ�L�7��yOJr�!������s��]��;��	�J��=_��L� ��۵�6`Y�֨����w�e��EY����A1w@ڵ��T�
t�GiC8����|�w�.����qޚ(�3��g�_�����|b���Ѓk(��(�A�t�8��I����}7^�fU�{�\/ͥ�F���3����xNh��xR����G2w���toXz|ߥG����m��
���]c�52�:.���\�P�>}ޒ.�������J���(�W����ö�j���k	t:F:!�{��̲��E��]��/K����;6�#�X�g���͵n��F��-����s��"���C�'����\�S*��$�}\��g�|��1�c���,��~��꧂9�	�B��=}�����DD��,k�\Πj�9�)AW�J�+e� �]��2f�5v�Lb{j�:2�-���0�0��]<-ʩ�$�-c�T��?hr�p�N��g��Z��C^�뇔@*�Uq2ݪ�.Y�S�����{����*�g�u�8��W]�=$~�1l�ɶՕ3$����w~��uƕe�n�Kt�(��ܽ�.�G��ww����y�t�������ם�ݱ`�X枣�=��j}-�녞��9nӷݙR�U)[wО�}7ޜ>j�K���V{�3��$I��U7� 7��N�t;�ؖSU<�)7>����VIC����[GSij�=����"v���i��T�
��R��o����WMI]߼5�f�]��ߋ��K��SD�����.f��YN6<L�xP��W�֘���|}=�����˞�뛓��cr_��0p��,�򯓡ع�n(�iLQ�vD��U�D"��\0{~<��Q�0�6�od��(�er�=�#���T�Z�oN^�I�9v����e`�"I_�*���V��G3��0�E�=�k�;�8h�qDS��a��w�M=�J�;4-��k>��A�mVyWL��&���]QAp��r]i��8�v��݂ǀ~2�b��|�ΰ_����z��^�}{P	e_��{�FM9��BJ��Ijݑ���{X�i���E�,m3�a25�<�:cɨ��|w�����e#�����vcYDخ�kF�>(�j��"tz�<������h)��Y����r���fT��f�=�����5�Ni�������Mc�X�Ҭ�Kq���I��ι����^��`��ܜ�z,�6uZ��-�+��km��L^����L����\��!��r��_-tB��w&�I3�R���z�rU�S���;�M�-!0���/�x�� �&XX��k(�c��wya��~��<��H����Ԧ����nT��i�2�"͸�2">��Ö���	h�-�;����T Y�gW�7�������ĪGFS$�T�mN� A4�jq�`��֢*�z����KŜ|�<��N'VN\�@:��e�e^U
��x�
��-��<f@�y�'�a�٭���u��;���W�uaZ9�����z���w��wg�c��`o�R�PX���(6��F�ߟ���}�j��9�ÁR���jV]��"��T�5c�E�"�3�g�@��̂�|�J4�x�| �� �T_�������;�7�*Y�yRz{6e�~SG���nㆲ����ƹ��'\|��v���;�OY�������m�~}��/�5�W>k6aU�Y.�U;�.�
���<q�pa�i���fޞt�ZXm��J���)s� �\�gs��ڮ���������jĳ�_�:���ȪP��Sp��.TTXϷN�v�E���_��x��|�_7�}�����tk/��\��&5e�Y�Ʋ^�K�	{\N�<��CN����'�`U����[|�N�m*q�i=�rugO\4�KO,?^uv��-����\�ٕ�J�X����,AԽ�F�ywҸM�����4�1^�s�v�ۼ��p�A]�o�7FN����93�$z����<;�Sl�c�6�+r��.����Y��\�w�#X��S���Lڷ�d"��]�����&��o1o.�����eJ!<P��a7`��l�#j	��CrbD����{���������O(�f�%��9]�|>��]&�B�s��ˋ2Dy���.�}2�Ci#*z��j�jyB�&=;D��ZZ�bC��2��ۜc�ʆq�`7Ϸ��Ѿ��>?4s<��;�^��w����(4#��U՜�M�%�g]�u� �|g}��[em>��v�[ԫtX;���<H�_R������_���b���;�:gX�ܻc�s�f*��Jd �_mb�dKg�%`��7����{����
���S�P�ưJ��)��*�as�%���u��x��ѥ�:�����t���K�᳚�Vk3!��J])����F��<�{�
��>�q�۠A���'ú��/�$'mI�,U�����IrL�h�zpf�����f*�@�bY.^�0�'e�h`_#�Nu+GI�S���gK��u���rD��^Of�Q��m �g���	�,�n�X�#�^�ʈ�8�1`��IB�B�Bk��ajʵ��s	C(�cz쒦n´ q"Z&��$"ŅҒ:
����0jX�wY
'LRLd'�̬1�e�ʔ�a;r0D��*��Pڨ%��8��&��]��Ć<n��k%�t�j�jQ�G#��y7D�!-���I����ե�U°����+4Qj����Tv;HȂ.An�\b�1�e��G]
�ףS�ݹK#(��"f!3�P8�Ɖ�l�:M�-e^a��R�T���J' Z��01���WX�F�AM���$�~u���eYR
J��W��r�p�Qe�R�*�!��Jg#�)��p�T�H8�ɲp�8լVp����P��D3S�j�]�* h���xq3WVJ��5@[@h,*��2��X��C�s�-��/)�)�!*�_�E9c �����S���5R���$�k�h-��NV	lU��R���n��F�a�	��.=\�+�u@��úN��`Ӥdϲ".�.�3�A1�]nHZ��i�EK
��]݈��]��D{	.��UŲ��a9��;6�N�ba-(����t�>.�0��T2M�n\2۷SH���[�� ؕ>տ�&�$��H��k<���q��`��[Gbi[V��mF1`֍l�UB�U���6��ҕeh�*Ŭ�Ѷ�kZ�
�IbT�j���TAm���*�DV**�(�Bֵ������A�F�J�

*$[J�6ʥ���DUm�KX�TTX�j#*UX�\Z�L%�+%��Qb�Y��-*X+*Z�T��TL%�XᢋUZ"�PF�k`�جQF�TET��5pՃmV-e������V�EEX���F�1+�%AUT���UEPUDQm�*��QXb�����h�j�`��DZ2�aTB֩�D�֪5��[DEEX�ʕUUkQ���X�iED�%,`�J�cmAk@�X���c
�TiKV�*�-(�U%J�U�*$XbԶ��X")YF%l��b֬H���EAKJ-iD��j�أQem�QV*�%��""� I$P�H?[V3�^�W7E�"��Y(��d�ف���[\o$4�Ӿ����⽣R���ϖu�<�p�cO�u�����Up�ty��p8�.�XnE��d�ʢ`�o�SJ���2�z���Og�Ϗ��;���d��z��ҭ�U�8��Q�	g�"}wg�^K�j�9����J�}��W���zro��J0�4C(�)�*�U7�yv�P1:9�!WAt�C+�TE��1j�����K�.�o	��~9^RൕJ1J^ �^8;�<���:�,�:F:_:�ǘ*�i�KiWa6i�Ctb�0*=L���<�����h�e�m�z��,��}��1�Y�]i�o�];�?J���p��=�<w��7o%yL�+��r���ڢ^;Fz'y纥�3.��i*�yƟLd��U�;M����m|B�]mغ���&��W�D�w7睅?��c6L!���j�E�x��<_�Ω�(��vpI���.,JԜ���&Hk�R��T� Q��@���F��aS�7~�=�R�z ���:�Q�.�U��0�6"l{\2҆祁�T"�D]��M?J�\���z��~�v�p�Uݡ.g����n�W��wgb�r�����?;��U,��˞���R����JjyZ���	�-����s�:��:/,�!~���[�wz���r���3�nx5Kޮc��M����`�ջ�㓴Y��an���P"�;>�C�Ȇ7�X(���{%���9lg��۪	ذY=9��mG�]/3mRw�^:�� ���e�ET4G�h�>��_s�1��Y���C�<5ε���5��z��uNKZƬ=)+.��b�U��P�.ɍh�ַ��Z�k�ap�xS��N[K�J�z��Xi���8�&��o�h ��_2}�vY��Ո���f�>���w7|��F��x��O[yG�*���g>�J>M��կ�@����S�ؤ�,�Wv�r=6�z�K~�4+�Â����G�=�pc�(�=6�����@g\�%1��KrVz>����'v�,|��>Ǔ�\�c�T��g���
#.�E��"#x�'�3i�,��ƕ�nt�Ac�ō������/���N
Ǧ�ԈUn.�@�ߞ]�"��s�w�>ܔ��2�l�(0/"��8��U��z���>�3������]��\�g�`��1f�w�cF��z��7��d��\jȨPO��,�׭of�u*X���^O^�ثM�M����fV������M̖o��I3I4���g�F�����$T7�(��hR)���:ɾ��=F�������x�S�~�.�_b#���M�\�	����wy;=B����0�̶���O�Qξd:l6
��@|S��.U&��<X9�D���1Y��X!�H����7�\�i�=�!�bW$EN �� ����+j�k�N���U��N�x����t��}���J��^,O�[TK�.���	gi�Hf�`g�^ܱ�q��5c�sqv��Ҕ-b�L
��}��]&�U�zL W,��r�_tme���� �Y���6c�9ఓ��Q�Ȅ�z�:�'>���U
0��P߹=�3SZ�/���`~&m����L�Y7$�o�
��)��=�;�=�lxeoS�p_b�8U��C��!��0f�R�}E���u�4��\;+��B�<z�[�(˙�~�w<lo�r�\;H���m�2��C�SΒ��4��`���܋����+=�n�O��r�v��K���O��f���Sy=�)�:�[�#Â%V�x2�O3��3�& �p��%��vP
�t���KQs����_�9�hJ�^����"3c�9؆Rw��9�Q���/�<7��}nE O��a�auA~=KI�tH��=��� ;����99�ȝ��J;"+�檷:gz̛V�E��V��	������U%ԗ��6�n&s}���o�,p��-�zi|�����}0��`S�gp�;#�ٵYsv�Χ7Jtzt�#�u��L�wΦ��C��$J��ڤ��zo���:w�^�.�fQ���wP����Q́l�y���6��>�:��40����V�@a��Z�g�+��Àƞyp�j�p�O�T6����U�9�����3�@8p�/����zf��u������]̡��-}��`��CS��A��Wm	���yS�#)�24�AۣyZ9yP����|5S0	u����sd�1s��v�
��Oά�6%T8�İ3�L�$�A���h)�(�D)ҋ�X�<��R�sC�����d�zKXrD���$����k*�V:m��Az�+i^�go�c[�����!ՉC�N��	���0ۈ/�h|�D����h�-�ċ��^��{Y��u���DtAb}�p%]nS��(j_�Qf�� �TUc}�Wνu����[�s�{&E;���D�x��C��h���+:8Q���^Ș!��N ���kY.N74���)�q�0*�����xF����h@`x|�|Ć8���;t[Oa�ͅ(����^��_A��hϽ��>{)O�d�X��o��g��8^�!a��;B�î���m�l���b
������[�!�f����=�<w�~{���>����(?y���s�\6`�2ԏ8\>G��#ϗyT������υ�*l�N�M=ٞ:.�rs�~-��[.�s~�B�Uc��W|�32����-���z�Nئ��U�4�ۭ�k���T��<���Y�X��w�^�Y��,t/H�M�߮�!w�/N�j����ޮ��Z�P��)s�ڼ��8��|�	t��+��Z3�3�'�5+f�yz����evӕC��r�\��S yU-�ī��U�A�[<u��xm�"D�xA�˾���N������}w�SV���FB΄�'�^^�(��;]�3��]��FZ��y7�w��m�f;p*�<�t~�̨��γC+��|_fX��
��ֆ��h�\��}������i��F�ļ:q��j���]*��XH���+5�˥м/�l}1��m�V=W��hT0k5t��<8�S���@GF 6T@�5��u�[�[���>��ct�\���b���Y���*�â�����֖�����o)��1ڱ���uOC`>@�ž!��T�_e�ږ�qAb<k{2�R])�un��^V���DN����]��44�)�V������K�r��V��]��	�6N�У���"�.�[)n�/��U�42�Z:�0\%���	ٽ0g}�zXI�BsAw|��5������º�����pi/��x����3.��J���׷�8j��j2#�K�ᇩ�+[)!b
D��=H���ݙz�UC����	g`�����.��sT�G��b�rXtg��fE�+�|+FT]�1@�f��#Fߖ�5�ag�-�1z�fdX�'�[[H=� �\���aω�{��c�T;����6�\(���\�<���8��0u����W��(k�DA�]n��{*^�����۱ߜ�}�&��]�x��G��h�v��K)�\�҂滊g�[��:��g�~�j����"v��s��Xw� x5��>J�Ҧջ�PσD����3��6������s^��sϱ&*V驕sp��!�%�;#��Eջ�3x��=�j�P�W~��Sm�y�?,}s�#�߷F;'��l{~�cn�{��>QU��9U�&Ro ���4��/L�#p��!���N(1���+��.�A�b���Ck�>Ds�1� |.�:�r�<��f�ڼ̓���'�(��ʘ��=T݇�Bذ�-N��F΁�_T�o�њ|g*$f�2C/��i����\��lai���ۗZ�fu���ql����3˯�S'J|k��`S��/>�.r2�5|��R갛��_k=���]��8��C��S���_7c&g���G�:G���aDj^�;��c�g�r٭��� ��s��s�;�zZ��5�j�����Ӏ�	� EG�D5-�al�&��r^���W0_�Tu�_j�u3S�^薳M�F5E�(t34�j�m���y+�݇��WOEܙ�0Z�7Y��G���q;�侈z^�u����mҁ�f��s��J��P�Ydo)_rVVK���R$���>�
o�Bl�R�?ap�Ȃ�}'�&7V)��N�~�ٱ��S�c$=�ՏH
��	�Oeb�*�O��˹�)T��I�ԧ���|N�Ur�IW^�r�`d�>�%�U-��9&��nz�r�Y%���.o}�:���s���6��vB}�\�-b�L
=�A}�ǀeC��4�c*,��&'%��������,���oʽ�p�\�ƀ��Ok���K�槥���M��	#N�/�g_���^gF����#�������u!��Չtpx;����`K1Y��%�a����OҦ��,VL�=���}�
��rJ�P8��<RV]^�t����rp�8ƨ
ɕ��*���"���C�r�2��t�ft\���rU�Ϧq�c��w�]r���K7w���v�F�S����1;o2�8>��Vl{��
����T�{ܮyW?K�YD�ϩ5�p˙�j���2Չ����o":����f�^��k����+]��]Ō��fE��{ƸU�N�b��}�A�5Za^������d[̆+�A��6rݾ}�Uw��Le�u���w�ʹ�eQ������2n�L�uWv�vh>1�����j��n��w�,���ǵWc詻�{����\��Ch���"�&���ts8� ��0hZ�ڀJ�(���_������.3I���U[�)od�l��oL��+V3���z�9���f�pA����b����;_0_����<����S��lc���^]��/q�-�S�LV�8��:	�n��}BiC�l.�h>���XW^���3�=� 2�m�2�Tɴ`
�L�{�獚v5dخ�G{��b�lR��7�/��!��R��{���l�ul,�xO��z| ����T�e��,Ʋ��c����>�Ua�q��Q�ÅE�eXϨ]�IV�º�b�#����]��J�[ �.����W~��!B���b����]e �Kz������6��l6t/�%�}�-�����۝L��2�ۙ�P ������\3�գ��I�8��^=��[Ozd�oY'�=g���k��w��8�Vy�<��hH��Μ`"�o y_��78n{l��F	�נ�,`��P����0T��#�S&\�h	o}���4sXo��t;�M�7���Q-�\h���t�lu��ʳ�ߏ��,]l��}���x#��Z�+qx+2m���2����3p���z�Xx���5�AM{���3+�0��Ub{6���b�=w�؇�}��w��,��R�O�M,\�|����8�\�Xإ�LY�	�\�^��k㪾�8el�C�1�*)u��{6�(��Qs�}L�
ʾbT��}<E���Yw�s+)�feE���2[F4��;Ӟ�r��z�+{y�OHOxV��kjfP����j�qmv(/�^�U!��Nw�x.��uA�.=H���zv�;G�C]	l ����Bu�6ꍌl��̧9z�m���I���v��!ئ����Bv_�,�a�8��uS�uY�#�� �o��ϕY���{8���c?Zу@��L��ןy?3R�'���. *���Dg�[n͂\ѵ�M�_���B-�E�&����Ґ0�#,Yu�kɺ�Z�O�=w�rS���������/ݾ�
[3P�%*�-0��˞�#��Ѵir�N���f�{Ӕ �SEf5�}�o^
��a'�<.��{��~�z��sz���WƤa��g��NI��A����`�U�u1�۵C:Y�a}�b��]����Cp�1&�y��ћք�J���Q�7?/�Z��P4vt��9�3���m�]��W.� ��*h�3�!�3�p]/Ɲ]�le�Nш��P �Dk��Z�f�^]r#�X�ó�����4o���.��۱t�0�
�:�{
]쳳ծ����*���Zd�
9��4��n�m-x"��`{�s����U�����O8�{����1��ĳR��2��N�غءI�AC��6�&���|_��S<T:9u�t��ݳ�ۿ̐=U%�\�#����υ@�}`���&���=ra�?� �4Wvix�T�����(��X�gu�<@��J}��7�)~��5��˽�����Eϝg��'pQ����Eg�U_��d=T�,蠣5�V;O�L����=2��Le^y9�{�i�%���W��Na�iFiAs]\n��f[���LH�n5�ǭ��uoK&kd�뗼,��:Ƭ>u��EŜu���I��ze~�e����W�=:�#�)l��v��Sl�tr�Ԥ���
!�Ej,!JS�o&��3���X�M����"g:R�*;�9�r���5��	��`�1U�u�pN8)��a���[Χº=H��;B3��ۏ�V�\�g&mZ{Z^ +�Ͷ/��'�iI���pl��������"r����$:.��9�P̊R!�@��C�h'����T�0���!�S��rG�V�Y{ ��Ӯ����8w%^W�p!T�~��YL��{}9X��ش�g)�O	�AI��yO04����rO����u[R���].zu��ŰX��t/i��JTs ��	��O<�v!d����u׎�?y�mo}�\���?�M�GeOw��b�,�g���kRe�Ztr"��\9�o�M��wŠ�,]g~Ew9Q5t�����{ۢ�5�l!_	-����,N�q?S��+>9X���B!�*�7�+���K�/�l_ܶ�AS �'Z�j���g�;�׃N�bG) ��BwEA�2!��jc�Wvb�iu�.�B�����DG���*����õu���R�m��K�xZ�C �WD3w,�|�x�����]��!`&��&rbmyK:� Ѷ��u�����y���V�G�jo�>�ԇ	-ҙ�^�Μo/+W+<�{R�Y���6LY�ls�d+�{"g��d�bx?ի{_l���|����V�>��0k�Uj��5`�kC�������o1I�b�f̤�t�+�B"�tͺ�0rdbL�
�D	Yx�*P��&1Fd?`�"%�Y�ĘQ6��@�V�5�*����92,�042ػCK�� ��h���,����5̫�[a�C+"��Y.\���w)��ké�&}NCZy0�R2ڬ�3��p���Ѱ�����V��n<yYX�E��*}�Rq��0GvH|qcj�8$�g��e�%#	Qẍ���(��ϙ*ֈ:q`�6�d]9-���E�3m2S��j�%���٠�q��nĀ���PIФ��N���SE��FD� �y��/��7���b��9P7
tdZ�B�%��)ip�v���,��e�`�b��B)��X��
r�P`��2�c TȾJ�t�����N�����v��̀ݹ�wv8.ј�Ԝ�����5�<��鱉R5��H^����j���]�*X�V�4�1J��ae�A%���홋

Ё�aٚF�+�Ȕ���٪8�K�ͱ�A:�ѹ�PV�4��B���ɪ�DDU�-b���TH����TPQ���Z�TR[PE�JŴ�AEWa���T�T��mmQ�V-m� �meb��TAVҪ��F�EV"�UJ6���V6�Ql�UB����-TA�ŘB�VS�ūR6��b1VEQe��cmm��ZUB�m
���m�Z
�mUš�R��e�QDZʨ�R�h�QF�+F���`�JŢTdEm�A�ҔX* ň�QQ�U�"[j�jQDX�VԵJ,TZ�[l��+ieV��T��"�1J��XT��Z��iE�
"�bb�,UPV,AEUX� �+QU�Š��%Ij-���KV++e�EVDEkb[eJ"��*1ej[KiQUT����V������DF������VҨ�(�����+l�a�*�Q+b��եj��[b2"�E�DUm�PQb�6�EQ+U���("��Uc�QbQ��*[T[KZ%�EĴ�UXSD
f�����sx����l�NV��͢-��r>�g��WUZ���2V?�w�x����5/Y<�Y���s`C�}�N�
�k2�K�rm���T]�Ih�.�A6�������n�3��<f}���0m��mW�����R�m��&RX)7�$n!n������Z�z{Z�nw�?�Ϸ�����|}낻>$[�N���7t�`q�H�Yx=äG`�s�_]�(SƐ�i��&<0:�X=׏�ח| ʣF��z)6r�����{p��lC�W�~�XUٙO��Շ�D���װ�����]��]�\�cOՉxjW t>��yc=����.aںpW���Vf�V/�Q�v�X�<�<������U�W�7r�7�D��ݮ���oQ�L�_�X����,�B��d="���ۑ��e��>G�!Ё�%	�� ���ѱ�L/��M\��K�ᗻ�l�j��L�ؚ��c�_�L�݆Yjw��ڱ.*�("([�g,*��M�����K��+FѾV��;)�������LD�N L��v�Ab� .���P�&U��TL�3��7��qg�����t����&����K{��Ȥ�/T2���\����
r�V��sՙ�u�P�t���"r� �=�'8w��9ޚ�{�g����]��Ze\Y�ͧ�	��J��Uө��zּr��w�Ct{ݞ8�uXx��wK�v�o�u�m�6k�)���C ��vk� ��(П���#:H��(m:6�ilj�,�f>`��/ď.-�
{B�-YBCe������D��u���ϕnV�{/��wbn�F3�D�6����g���+���֬QV��^D��A��sZ��W���Y9����^���ɜ3���:ΌF=�J~���u!Z�COO�!ړ,s<zřk&{��:g�+W��,�s���\�b�x��G��*"��ə��,�a�^�4க8��լS
�����ؐ���!cs湙�p����²rF.�ϱP{�U��'�^�OG۞`�8�n,g�|�����s�U�?��s;|���1c8�$;i���=@�}O��WHgb|C�(�=�VaP�V���J���.�/by׳��P\X���v��~�2�,���Bn:˹O;(���-ö'b�;2�τ��]�����Y:����:LE��s֬L=��##A���@UQzf��uڬ�Oa��i��WHM�'�q����j���2�I�Q�D�Bœ�~�v&�^!���0��t�nY�ד�41'����n�h}��@�9���� $c���-�s�'f�l]I��39�2E|�t	��6���� ��p�w�3��v"8kOa��K}�Q����؊��#zv��՗�)�9R5�fo�z{Ճo��j�x�H�g_u�t�\��b��Rn/TsvKmN�e�ot���x`É������RYR���P���p�Kn�Uqz���<l�6�'����{���:�ӄ����>1S&��Q䤵C�>���3[�To"������'������{�"�ǃ��̣�YD�mo�e�y������zC2�;���KS��b�f��c���e���ee�" |�¾�����7T� ˖��T@w���66�t�K��vpZ�G��;�g�D�fѕ]�R�C��|Qe�,�`��.<��=k�H�F�]���vV�$��*�e�X�3�Г�c�M�[5�H�����$������K5�gע�GFUzt�}؆���uGC�u<9�2gt�f�z뽯����	�K�˴����V��Ζ�	є�q�V�9�Á�W�~�\����0��m���<�3�� 9�"��a}��_x�4�yK����r�߇��.�x���E���z�}��#5��o���}H�s*�hAu���\�g��-�x�<g���*@�,�֌A���8a~�=��s%��C�g�p>λŽ`���9�ꑷCƝc#<&�����%�S�+z�f%�BƗB��V��L�X����yt�5���(r�Ҝ�Z��R�_h�Y���*y��W�Ԯ�G�Y�r\g�Ea� <���uC(��|Tw�ܮ�U������r�}s�=��l���J��K��e��ʞ	SKȁ3�&����Z�1zg���F��ȫ�\Ɋ>�3^lX�ih�j���\./:��ϟ�'U�ĸ����k�|�}����@A-˷s�t���wS)�۵C:��"����&Z�nf���W�$+��h?�*�\��nR��ŭW�Z�� �<���x{k�{���1��W�
�pI�)�v\%�
wF��UUüR7^ t�* 4z]����~�ov�+�e"T򦈹va�	X�&r��]8��ͣ��>�l�m��e�J��>Ix]:����B�|pN6U��K^	K�������xV�I#��өm=s����SĆk>��q�X��K�u�YE��8����4�´6_���lsN�+�l�0�b��cz�<ݚ��~ �<��u��BH�t�՜�ׯ������o�O�3/�b.�3�Y�aݧ2o+�Z�*��3�-Iٍ�׋��N��d!��"�o��gl.�s�k���T]��CKS�r��n�_��QxT����h�lE%�X.�h7�<g�Ȭ�kss��R)�;ݽ�R,丟s�[cӮ��L	Mt [5��4��<�F	P�PۻX�a~{�\�d��nOpDՑ�f�'��(��5�+2����
y[�b�|��F�A�������
P�Ւ��w�Nme�����]0��,��%s��mo�PwU�D�W	Д��H���?7C<���uJ��k�i�:6�ۇ�C��2��m%c�R�͞U2t�b���{��nb��6��ߚJ�am�COƥv%���&"wɼч�КF�������u�v� <���m����E��=��x0�(5�1�Qp�t9yEX�j�Y��UI� �\����=�I�w�JV��zpS�n4=��pg���kz`�mR���c(�Y��hA�L��˺�^�ힾ�v��FO|s� ��v�ֶ�=���(,vU<~�(p�u�|=3�-�~���	E��8���^���J��#�׆Y���G|�VЧ=Y��'�L}]���uѻlᆖ�<kCݲ���/���b��l��3zs�C�6T�}�{�Y�Xj���&���e1�|Y�i�;�/gZ\o7��e����kbv+jЃ��ٸ��L�֞7u�1��X���O�n,��Tf�΃����)`��4��B�e;��j@N�{�V������x~�w,�G��Dz���,|���7�EЖ�WS�a�(1
��(�P�p�A|:\�2'��puյ���b��L臦���v�]�n���Ԉ�Uʂ4�C� ��Bh�5 ���U��	ӣ���u�fҩ=�չ��n���z�w���0m�� �� �҂�פ�[T#X���̌�)�.�/'f��T$�5�n��i.,�WÑ/)���q*B~>�nӊ�574sG3f֢����x��H��xB����;��0(O]W���[�.����`�\\�cy{}��sN�X��6�7�v6t�N�����;g�maU���Egy��<F5��E�������a3�o�TG�͑z���~
M���<U��F�U���Y(�.�G&�V��w1'���p��:�:]��~�b�8]�O���OC��\�b�yJ@���2-���fo���80��c�٘`#��Ǹ=�1b��cs�32.��Å^N6a�Mu_UƔ6����Oړ��o�7NG{��6��h@Y%BV�N��8���'Ԩ/E����2�^�m_���x:�hҺu��M�;شs�:h�X��f)�M�W@�ǡ�"�mmE9��%��y�__e�Ֆ篐��I��Z7�gV�����U����x��Y��ӟP>���Z�e� �kj�S���58�����:����er��cw�S��;:��5��Xs��c��%��=U�n�{���u]o<8>3]z���Ί�u����+��s+�yu�U<_�G ͩ��o���^:�]lZkj�ʺe�h ��!��>�k'�8Π�噄���廃*v^�t����}�q���K
갬�Ī���Ӧ'e/W���c�$at|v�'	�Lx��P+�ԖS�=QP�:	�Kn�UgGYC���ux�ed�S�s ����zϫɓ-�Y���t�T�/��-P�׈�9Vk��]v9������TisB���c��_�����X�荛��@S`��UzI���Y�id��D������d?a�-��6$F����*�U]�IW���rFq e�C�k�91���O�,��$�,���1���G�0h�0�t���Y�9묃O�I;�)���V��#��¶�,��O.��K׼e����'kS�Y,�,U+&$�Wm�~����l�Q<w+tuǶ�ح\>�7�1h��ꅡ���3�,J�Oe�w0	J�#ػ�N�f�.=��`fpe�E݃�u��ើ���LGϝxR��O'W1�^^��74�51��BK�n]��X-�'s��}��M*�j�P��Q͇�V������lm.^�\S��a*ɼ�-��>�Ƿ��`t�k�)��.�M0,�Sy[:=y���H��CP:�z�U�����~��w�/q}a�ї)<�B}F���E]2�@Ⱥo]r� �R���j��X����=�Ƭ��Vw'���?P��Z�SM_Sٹ�O�'C�DA��Ub���{�\����pt'˱���x}l�(�OfXC_�w]�M+?��Ck�oaU�r�C�y��+Z*A�O��f���.�W#���|��3�}��cZg<�| ��b� ���)����0x+��7��~��(g�!��ẗ뮮�C�T�@Hr�d	k;�@�B���_3h��x�u��#����0G�]�릠��X����=R�񮩢��x'R\ m� ��_]f����:}m���DM[}g�0�Ͱ<����P�@pK���QUr�<h*��!+o]�l��^�y�W���+�1m@�7�.�Q�W\��Co��K�:q�8�⁗g�z�X� ��v��ɾ�c�n�%��1t��mнܥ�T�y�Q��^���u1�(�}$A�����ķz��ۣh�&��r�Mx�\AO��s���k�D{�u-r�`�Ϥ�(=�쨇 ��z�1X�J�s��ʾ��)�Ԯ���p���
�}�f�ou{�,	Gx�`py�!�,���уa���4��XTÅ#����u�݆��%����w����:���y�[>;Lg��z%+�Lԓ��xE�]9�޾��^�٭�J��Y�e2	cD�HH���Ͱ��BO��:^����	)���^���7�K�jP����k�PSIU��8��CQ����b�b�$.�<U����/���O9y�W�,�Y���B��KL�$љ�b�mt�oFW�$��o!��a`k=�z��+'�B`����t� =3�k��f�L��\�DZ������b�v��.J;Z�#�6�\(�=o9S��9�P�ߵ���w�	�jϸ�eߊ�������q��Σ��9���Ǹ�3���!N]f����e#�wJ�7��'��F�]��X+a��^?O�3�j��M�C���.&���IݱI4�C��x��P�a��!� ׻�v�!��t�̭��\<4���X����DÊK��.UFVE���KB�\an!�r�� �~�J��n�_]{����c�ۚ��򑊯��<�_g����H�f��=+x� ��/{^ӳ�߇�r�����6͑g�o(��!�R��Jo>������k6�p�h��c9Z�U��4�r	.���]�D�i>W���;?��f|j�Z��7OE�9yEYN6�%�� ��.��t�M��FA�y���i����nX�x<��Px-�~��r��Ipb����G��J�̋7��Ւ"�уU������ܺn����R�Gӱp�w{s�>x�ę�������	*�2�w�,[;��]R��W�����{MO,��	�����1�K�*������'a6P��ЖC�>���y���o<X�&wIGQ/\�w��g���J|u5tO�s9H�s r�Y�WP(�<�mE�3�hы�J[���u��o��9�}�h���f�렍*q�B\�to[��V8��sQ�U+�	n{;g��\xi�2�e�U׭�5�`��Ы��MW�n�/�H���ɚ_�z:�.���6��>�w�i>�`o+���� �G��p���7%��y�/Y�Ǚ����AQ��ĬWPE���(s���w�~��	!I�0$�	'��$�	'�@�$���$�$�	'��$ I?���$� IO�@�$����$��H@�xB��$�	'��	!I���$��$�	'��$ I?�	!I��IO�H@��	!I�B������)���;v��%,�0(���1"�� x�T��PP(QH �B�B*B����U*��J�EBUP!R*��@JUTH�JRT��R$=b��U*�	
	IQUH�T�IR	RPT��T6e"E_mI �Q@T�u�R(�JR�@(�*@.��� R(���)D*�)�B)J�M*��	H�T� DQ!HP$�HUR�R�@JPJH��*�RE*ld�
�R  +�T�V�]�����e�[�`QE]]ݭ�r��mt��S��5U]��Vr��B9V*GK��
��"��HBU%A"�QB�A�  ��E6�S�]�kv�smE:�쩝uR.l��5���$��.�4��:�n��4܁�j�CX�d��DRR*�UE'M�  cw�6�K�n�[��J��N*��˅�T:u�,+mv.��u`��Z[�+�e��]˚�M9.ki�N��ڭ��wq��]���kw3��U#�"%EUDU�m� gm�^;-)l겶ݰh�7Ev�� �Cޒ�@�
(t7�[p�Р�B�
;��(P�B�
 ���C��CCB�
9�(P�B�CB�B�]��B�

 î���c{F󊨪*���	H��w� ���ATzv��Zʶ	��Z�Ͳ�tt��]�v���g'�[��۶n�c���]���rY[nZ�5W:��5��m�k*۲�n�ʓ��wn�]]���E
��P�T�  ��%Ur�ݮq�v�4��)�v�EU.p�wP��S����4�]�sr;]:l�s:���nwm�R�������@vSi����v��Fm]��P�E���
�%Wx  ������[��n��m�u9't:-�Tܥ]r�����\���vM]M�ûm�[���t�ݴ�ӹݭ�{�N����l��]�I��t�!)�TE!Wx  s��Z���ʮ�Qmg:�ܬ����쩮�l��[�v�ʠ���U�I�hh9�s�i�uw%k�e���wv�8�iӮ��[�.�3��AJR�)�  ��ݜwnZk9Ww]�:rl�]ӻ�v��vD�t�m���Uɦfq�\�\.��%�;5V�w7e��l]�;��뻜8�Mvm�:s����Rm�T%E�*U��  �zi�JjꫮӬ+��v���wu�eV�b+Wt��vpG)��j�탗j�:�ܥ
�T��Zuj6�O 2�� h2Oh�JJ�L��MOI�M  S�A)I@� �S�&���  $�B&�R� $
X
�D猒B@�ވ3+�W9U�Tv^�+�X:��eA����j�����B��}��$�	&�! ���P$�	'���$��	!H��BJ����������3���s�;Z���`�,�� �0�/� �-�7��n��t���Juw���!��f����8U! {�z*���m�l��Yq��Y6�M�Ɔ,�J�f<�aU�d/h����_��F���u�T���c>p���tݟ��RK�U�`��1KA$^C+落S`��de ��WfYo��T~bk+K_`�ÑU����X�D��s�BP-iմQ���E`�I��WZ��SZ-}p����y^%���*�q�m��]I����R�^c���Q[,��u�Un�*q'��
3j�Z�Ԩ��T{��R�E�QU��
Wi+/m��H�Ƅ:cw�{.�8������� [1�kr�^ 
t�*faL�[f�ূl%t�n�wYY�0P�L�@=�3}�1m`��ͤ�YV�5:r�/E��*���r�)V%�U��� ��k�b���Y�����e�,��@�I���?�n\@���Y*哭�M�{f��M���F���h�
X�(��J��!�$�pk����tQ��b*IYH�ܷ-�
���d	wF���Zh�G�59S!�n�D�~��&�T2�\�ͩ���CZe�!h����tN͍J����zCQEn��Dx�b�śL��Kʘ�2h*��svh���1�GaUunL����%V<�,�*����l����#V,@�\�Z�n��%� *V/��ld9NL�3X�)7z�Ņi�	�E�h��nr9�N��yy�	��,<!�TN&`Nk�����5c2��U:i1�ƫ4���*��]flYkhRl˹�e�ۦ�A��Kb^���KQ�i�a�������KVf$g�^� ,��Eձ� e�E(f��Wh��[˖�i*�1�ٶH���l{�&!�Jg�*E3+w��(�q�$��v����h�h`�ᬡ%!���lٙ���l$�^F��[O'Ɠ�
74^�ˏu�9$�Ci�a����Oi��9��m;!6��ڽ{N��SUz/�ww3^U��@[-��V�j�?���;����S���x(��v⭙{���$�5�lߡ'/U�O3Lxޣ%Iޗ���NU�m eֵ�#�6�L�6�o!�݊�t7M���,E��w�(�奔u�f�Pܢ��.�NS����1�7cq��5XW�t<Z��$��N�6`ebI�H�&+�iD*H�`�U�i6�,���j��(��jh���MFg(ly�ci�'
�2l+�r�"��V��f�r0��[��[�r��"������R�%��%�ei��欣�H�*��
k �F�g�hۉ��������$y��wt�Gp�ѨLZ�"h�F8wqn��FLX�c��e�W�K�V�бeU�K0]� sL�Vq]n�Wm;����*FMgn|�M�SF�)k!)JaNC��\�"�7S��v�g.<w��9-i��*�,%��MB��6�����X-$��;��I8)��^`!@�f�Z��(j�3�-#���#E�bʏ�2�(����@+��-#qֲ<0�\�SZgbD�8wG�cq�=q�4�-'oq��ڔV�/Z��t�4�1$�.�D�^Ru��]ɟ�P���)JIv1�h%O"36��/"�H �cA�ݧ4`�T��l�l�Q61Ӌ�u�0&�q�(Y4]����NG4�
���ͨd�d�tI�-���{.�GZ�g5�z��F�k+h=E"V����0���"�Va��T�%J��M1)�ֆi\F"u;�`:lʙ���n�ͭ���iC�ҷ�]��X�+C��vXՔ��&Q��E�0nV����ɥY{(�̦Fj{�F������4�I�j^��.��P�d����xd�
��mf�2֠�N�e^1��d���Lw��x��t!Ye�M�On�2e)�M�$��mֈ��8C�S����wB;t�+�ݛ��5��j���]-��nbn� ���6}r�H��8*����w�Wy� �m��Lm:�3-�TY������K0�ku
z��Ѵ���n4�Ŕ�vBέ�KʶEOehї��' F�O�ښ2����t2�)�X �3L7b!�F:��M\�\c	��᥹`@�m���͋�P,p��Q�"���m���Ӽm�ɳv���c[Ghm�`)�]�v��`"�hq-��Y-/��n�� �7�K�����g`T��[q�����U�Eѧ��n�1�ϋ�i-sR-�X`�Z����7-�-<���ӵ��l�ղq���hq;4>0n�i^nR�S.^7���B��0�N���3rV�����4�e���m8+Tۚn<��AjJlmf��� und�E�98f<%��+U'�*7T�a��� IC��,F��N(u����Clԕwz�M;C�]�F%ܹ{v���I�x��Pl��C]�5��\9��)�v�v�X2�6�"��o%�m3j������S�S�Xh���^dJ��N�J�Mb�W@5�ӛ�惘7{Kڇ9m�Z��/^Q/�Ү�RY$N��y��e������V]�&��+H�׌=8_oS�Y���@��"���+��ӲdH/�<����a^��0h��F��b�i�d��]`(�{���&� [v�ed��Dn��1Ї5`�c
��.������)1Nӟ1��R;D-�d�lI���w�����/)l��
S-JWzm
����y �kP���9lV��dbD^VMݳ�b0��3@q	�J�)U�%��@�v��CI����2^��oUG�� tӦ]���d��)q�5���VC����`Q˼�b�y�vf�M���m6ͭhf4qB]�Qvw
���0��1Q��oF�[!��Pי�
��
� 2�̳Y��iT�:��]m�iy0V��Q`��#��r��hT[p�̏
$�ݚ�݂�b�KSo2���K��w��a�AX�����Yk(�Z��Mag]��(���j�q��aˍm0�Z��Q��Sie-*��ώ`�xu����"�EG	��C.[��A����Ūihz�"M���5���,[�Z�SC���A+�D*�hnk$n��	�ϲ� �m�6�^���dxh���fєJ�\yJ쑖^���k�9a`V��-�e��(e�{2�Uָ)6�r�n�V��b�r��B.e�Fb�Y e-�R��d�����t��m@�+w�#"yz��Ԗ0Vih�f㗔,�k$3u��Q6H�S�,�Q*�r��+mbsr��l'��h|L��]9���,��oj�Z����b��4h6�/T3iҙ��i����i���ӧ��h�*�a�lG�J��Ao%Zwl^w.��`"�w�=NV�k$�zj'jh3Su۫�ܠ2��,��J�����Z��Ȓ"���˻P���V�u�;L��nS��-����G6��1X�@�١�i�n)����ʀ�U� x�&��.h贲KN�fh�1ݻnV\�{y:a�3E\��d�䶷����7��ff^욲�:VX�M�q�X�Ra���G\c4�Ƀ��ѧfL6�К`0�*��"7�^f@ �AT���(�n0�kב�.�6vT�v	���cr(0b���[���5.!`�6��jb���.�^"N��@��@m���:��A1���ف�h�˫q���p=�Bkp`����oCA��r<��<�k�+H����?=�Υ>Z���-�+d�o!\�r�v�W�[2�2��Ab��Ԉ�i<J���tƉ�� Ix��ɀn��1<�u�Vuk�Ux���Y�:�!�ҶD�7W��:�0�%@���f�~������Զ��kL�e���ĥ2�ض��h��E�P�j��!+(�6��q6�x�ρ����6�*7yn�L�0%�L�����ÙY��/c�R�Z�ח�M�ua�!	f�U�@:v��ٶ��d--�5R�쨄x�i��u-�*ic�hL۸$�b�Ղֆ��2MwY`0��֪�QZ#NK2�)W��X�Dhͭ�Gl�B�Uh���j۩):��)+w#�+��b�S^����c݄l:�Ok���[m���r��Vn��M^
i�*tO$��x����f���'�C��~�%l,�o����g��Ϥ�U��*Hb�R���;x�K*�nXP�t�թF[T�wd��n�/j�s,Ǣ�fo�j;O7���6M��,PxڴrR�/�*ӱK���-��-w�X�2Q�X� CI�6,R�0VTt�T����� �l%�#tm����}xfB錵DF(@��ome^�Y�a&�L�\7�Zu8k�b��
AZr)j�8Yrt��X�K��a,)�Q+,a�;#%,+V���o^RXִx\0�ni�(��R���@��� ���B��a[�ɺ+-�Z^*ص�J�n��㻣KdDV�����Z�uW)�w�@���cim�B�xŪP4��W{�:PU�!9�v��u��k��:�e��QOkuLҾp��[u��F�6Z��8�W��.)NP��qa��M��n9Q��j[ߡck�v鯉�W�+"߃��n�m���B�Ѫn��*�sq��N��t���ΰ�`�σ� �u5�m�^4�m1�[�yG2�T*�*, ��%Ր�ۭ��ڱ`ai4��nT��-��36a%{��[Nn,5�];�gd���t.�Y R�d���~���0��3J��hT+
��J��d�lУ*=R٤� R�0l�c�+j�02ؙ+�
�G�,AF��ҹ�U�X����)�ڰ�ڌ=�#Ƌ��P�.V�^K7mx�`-3bv��9&�ҩY{�S���4��Е=�yN�#$R�Ӂ*�j1O\X�٬���y0�T�h�"GD��IF����hE���S�h���Av�hـ�a�CE&�4� v�)���vY�K�I��V��)FpR�E���*��6�&ॉ^ݭ��귴�HS��X�M`�`�ѵe<jt�Ϧ\5���3��^�XR�f�e�Hd���w\׮JI W�9` �;��åf��M]4�ĳtm�sLm�1چ��#�qZ�����A��8�tl�a�Q�Ͱ���V�#�[�Z�3.K©=rckj�M�#M]�v鷉��
�jȠQ	a�̲њ�Z���1��ݤ%�l��%�MVZ5�\��$n���������y$�&���J�sP������V���ޥ�In'Gv�p��R�F���y�<��ڛ�kFr���^8�h�	$���a֤30�I�s5"�*������s4�IcR��
TD�f�WVV}�TE4���n{�y��/M��R15Z �AT�Q$5]�v)2�o��mZ{��55K�3q�)nAt-�c�*bx�Mֽ�n��C�Q�#]e�*X�F�*����_+n!F'n�J8�W��Z+N�qȲ�PXƁ��a	�^
�ٙ�k����J��tNVKT�IH-�.�4*EL�nf�o$:)K�oh�����ʱZ)�N��i:.!c�j�������i�������Lbc����I�kq����v�\�Wk�UˍJ���Y���e������� R�ع�)d�r�i����r+���T�^�[X��L�R�5-V�ge�uzw~�F;"�� �1�����^
k�,j�eBbM�@�.�	��NEA��f:`[Hvh�TK�y����m��n�]:NJX�ܲ��=5�2�hfͣ�h=��Uԃ"�&�f�"㘗�:Nmj��1�
�����ҏ)Yq�ܽ0K����pD�d,��80cH^]��IMK#4�rj���ʻ�E�z4��4^�1X*��Z&(M�zq��J	C>�i��n���2E[N�ڽ-�H�h=`koCX<�-�,�j`�+je0���bp�����n���M�#.�@�I��W�+ʐ��k�G�[P"���dU�ʚֻU��yT� T2�*��q��#/�B�m�5��殒vDs%mc!ڷ����������@$�W���纜���ρ��iݍe�P V� SF��`��qv�em圛gfJ�-u�-��,�F=�&!QQ� ����Â�"s]��ׅњN�$�m$�t5(��0 IB�U����R�4S�1�/Z� ��d��m�֝�)���Ld.Z�r�Yt��14įU��7� ͻ��F,�����"�%#R��gB�M6��];�������pbv�he$N�\Ոj֥��P�զaо���i�ě�c���ߵ��*���w1����\J-*f
�?dQ�[�����T.<��#��h!c��|�A!h�A�
�s\�,�����D7��hA͘�ZU�D"J���"ʽ�eި��J,U�Î���*�ŭʳ��܂+ٟ�3��&���Y��*�ʵB�9/u<��0�l�m�Kb.��v�tUM^32�hmC�S�,o��3f�5)a�8fP,��.�ڲPl���j���&�u(fO�H��.FZK(��a	]A�ue�ǎ��H �=��#*F)��H�B�R�K\a�RT�T;�AnP65���[�tv�	5d*Y]M&��gE䠩`I�޺M�Ԇ��s[̏J���,��Db�i�	dQ�u`�rCU.��n�$�vN��,�ےnM��lZ��~��S�Z�X�Z�X�-�^J��1�,��)IIM�� �K.d�[�<yb�/D
���7$@ʶ��[���L#��qe'n�$>@Z�wl�NL�
��x̙7tm���~�6�?+U4m��
������[��CV;=�k����GN�ukz�:�wG��bk��iIkt.�+t��C���L�Yo��u7�z��@ lgv�M�E��(Cvmk	sZ�9E�9kJ��H�9���v��;��\+;�:�u%�o��揉qf���/v�n�V�����=]�1��H����u>����
��V�]\��q��Cq묾�fpf��Q٩x��	�Y�qaڜ��p�т^������r���>ZE��5�[�<V�U�v�j���+�ee��D[����9C�"ۥ�u�R��5�R�ث���b�YM��x��C�qi�U�k2��[�j8E:/N�B�-=����.u��Wh���p�^=nˆ��&S��bLB��&�:�^ZZ�Tl[TuM�]�+v�5�iV� ��,��ٚV�+�}r96wSޱ�P+�x#I�\�+�b�+sz����l��}آq��|�Dx�4v��Z��]s�e�cuT���A���i��<�A*�����uw��mM꺎��uղ%�_Q+����2�v�Pl�O���	�a1^�Gb&w�1��Z�7&��YR�]�s�
��eA���Az�u�'u���e�wy�=�@*��w3Q�� �Y���%
Z5Y]2�3�Tu�E�Ƴ{;u]6�i^�pʚi��3��5x�ȷ&p�\ �v�9�}G;NN��L�-�7w�̛e�j�)��1R�t�C�e�t��fT2��7]K�����թh{O�J��:=�7n
rWu�H�S���z5A�<��J��G����q䒆$��ɴ�����ʇ�t���ƚ����l���س�s�e�e=
WLv[��"�wf'u�"��Zm+�"�]i\C.��ի�S��*�������㶗R����Y�T�!Xkp>�˃�	7��f�=�Ϊ@d�v(x���ɐ�]�=��*W537k��C`E̜�b���M�!�Ko��w���.�"��;n�dPw6�F�/�4�
U� �(�P�S)��/-�y��d����(F>L�g6��,�T�{7Co��t�h�7h^���9@�M
���.��>=��51)\.	E*2"�qL�����_M���2����3J�VQ�껹�f���_A��xӮ�O������'Z?H���-�17{:��P�49��I�����b��W�e�)�wDl���c�0J���62��k�����;���U�,P��a��L�j�ҙ8�u���.���ۢ�V�:tF�`o�\Gؕa���R���V��7H7$����������+ԇջ���u��]�`�׍$���-�'L��y̫��v�*�B���]E����n���u��vd�CS�����ܤ��r��n�$��W�L�r�ظ�y�~W�>~nd,.Z����hk�m֪ל�!�AK��tctmf.:��׀+`�q�/U�l�ȭ�f5\@���u
7@n��g;�Z��8���G�7�����{��S�����e̽ήp_@��i�ۦ��K]�]��1U��]K��fM�1v�Kw�,�ɕ���I:�x�#��y�B��% 5ܫC0�:p�~ie8��9y%�i͏�0S��m;�p�S�Q֎k�NҡhgM{#��b^t�����5��f�56�:5�����Tvo-c�k���=�#	8���tNn(E[;wK�X�P'��qܣy�iF�Y\˶ٚb�V[��Y��\��W�5��Y�}>�w�+yMY��Vۋ�q��&{-c� �O��] 4Acz����K<���6�۞���'X^�3W=nҫWi�Mr-�;�'X:]���#�	�M'*tf����B(�~��+�n���9�N���;�����̺�K��=�+ő4�v�֡�Y�ab�pLd��Z/v�c�U�Gl�� ���n���~ػ�r�<�p ��f��������3�0�;���e&时Wa�:�g�SZM�Y@4��=X�ij�z�fWw>koI��归��_12)��h�[)�q�G�8��'�n���]2�c�VZO2�u.�Y����}-k�����̠���ːnwA����]V��h��ev��\	p�F�������I��!����V��rw��㝼s�[aټ�V��,\�Qվ�)#F��f�J�c;�1��qs������d˶��f޻����]M��Zw�zD�R�-�s�R�1CW��r�e��PE�R�Q��A�H�V�M��6���ok�i)knT�p=qa�g!�K���0뉬&g!���&��(7��Ő6�{n���;�V̜6�:+B:��ĭvV�5��]]^�a6q}'V�"u�W��+d�8�r���t)�y�B�;�x�6r��J�B��wZ��d_�5��\M�u
����8y�yR`X���i�׊�Gϓ�,��#���V5�����`Ãq=��$�b���Uv��-t���%��JM���xes #Y����F�Z2��HC�P��95g`M��@�����Y���oE%a_�.�Q��w��5q��WX
 �3���9�Ҩ;�e<��5m	�Jip���.�d�T):�JJ�� �e���\�����Ҝ�� J�<옵�6��O�Iv�� �܍$�U� ���nT�{����{���+�r1�a`Z��4]fֳ���L��[s�F.ܤ��آ3���є�:銲ر}�4�\���RC���a�t3��g�w[K9�\�o]��0��[���(3�BsIWu�w��|�T�Ħ^��3p�8v4��L�\��j'gq�FÛ���Wo�A��@��n�ڜA��l�%�kೄV����-F��-�l{0�@u@q]'M^��-��-T��7jX���ثQη�v�v~��4F�+���69.j�Eg�cN�-����Xk�VZ��2�8�������sw+P,�Kt`=e=d/-nV�|�8�n�s\���җXy�U�U��{k,N�h�B:�2�n]Am5B�1�or���b��.6�e;HR��h$:��o啁�Te��Jk[��;YG�_m,�2�����75kQ�%m.���2%W6;��scw�`��O�:����:o9��U�\�&p+C��d�n>�α��O�89��f��[Da����n�X�W\�"��B�ghM�`@��,�l3���:m<n�a%J�N�mp���4�A�ŵ���'Z�ѧ �K
ո_G�/V��*8�b��Z�'�	���N��2:�Qfh�x(�F^\;I֨#X�^qU����5�	y�s�2�b�Gx��\9�ܥ&��������{b-+`-I��[H�Yɥ����@/��gwL���.�d$� ^0bsM�f���o��U(�q�}���^�k���u��wg�J[g$tE��u/�.�ʛ�.*���mW�N��;!F�{/���	�HdV������.�V]�����w[WF�q�r�v�҈�ݳӤ��{��o���k��eR�t��ƆjV1py۠=�̠�U8=���ఌ����vGksZ��Q��&D�R�������/hu;�b%>�*�{i���Ԯ�= �"K��X��7�b�]�u�r�u�xK�¦�y��P����!�ѡ80�B燝�x��Ų��*f�E;�^���;2��x��h��t����}	f���إ>ә@�\�W�0�i쓇 �%MX�%O���b�v���
k)I��;:Žֲݾʐ�%2q}�K-��WX����v6�y��o>[�
�%A�� �_[�7Vr�D��R���7�.��m����Vn��5���ʧ)2Ǎ1ɯ�V�TP$
~��-�}W��6���� d�ë5`롈��rfv�ڑ�[f��[���KiR���$8��h�����l�1u��4V����-�}
}ǟp߃�,^m��Eb����{�t�ݠ4m�*ۣn5�n��TO7R-H��9(�K�_u�y�B�v7��R����#A�V��[V�K�Ź��t�о{��[��c4�1q_Z��m4^{�ӫn0�}J�����T��������<����ִ�-��x�5���ۺ��=8G�,YHM��D���C�(��a��]��.s\ճ�Z�wy\���E�u�C��K�:�%G�.RZ��gk�� �<���!�\n��J�ʽ�`�8q�I�אU�X:7�1Z�0��8W/�Cڢ�M/l��+!��Bhf�[�M�����sxZ�U� �Sa��S�S�S�̚6uҍ(0C�nJ*l�o<�t�E|p�J����Ω|rI�,T;���Xq��K�������'[�C�M�$��pt���@ɱ�A���vbۼ�-�TzqU�ղk QƁx*nj$V�Ff�{�ʳ�9�����P�Q��H��v�U	��U���qx���;�GcT�<���A�ʕ��G)�
+��2�K�7��Z8�W�h<��a��V*d���J��@뮮�m�:)D�w��W���
n Q��c�.�3���O�Y�<�ߦ��n�k��1���Kz�r��a�@��ܩ{�����.�HM�f�]�E+����x�hU[hN׋f��-ICS�"W�WAk&H����m�8��X/8�ĕ,��`u�T4�O� d�+e7����T����Vt�'$G�� ��y�76���9*8����oGMy�Gl<�Kю�����2e�-�
ᑲﮫ�=X�lj��B�]uv����aT�/��n��UO7q�:����6�M�w���q'�Z6����ҥ+���V3�����/�uw�<x\��H��锩���Y�p��̰��vLud���r���t�p[V��co k�v�Z�������"��y]B��tv�J��|�Pťwa�Od ����vy��JDZ��2�r��N��$�+t^m|�>�5����������5�5q�sZ���8k����'C+����um�]�Kx�_n�Ŗ������O1E;��ņ��"���&�zΈga0oh�QPs��p	���%�6�:s��ws�Z�^w��!0��'�.>�[����~F���^ ��>��+w�~�1��M��t5۠λ��Kq��n�m$����2/���#:u3����g[�S]�'2%y���n��`�n�q�f���g��j�� ���f�b�+{%Z�z����ָa�Z���ZGfq�v�=�/���/k`#0ɫZ�Ѹ��=hj�u�KQ錋����(�7L���ܱ�fu.� ҅M��r��S;c>�����C�������H��iV-�'�>��5��uv�;J���њQ�=��;g�É�/)��gT9�)���v6N}3���:��E-ܴ����}��)R�":X�hvo[�P���`�i��L �d[#��T��j�ՠo����XL�,����Ηq��/.޳�Η�Zt;�kJ�Ɏ�&U�˕��;8]�d�[��!�i<]��� ��:��t��(&�i��\ar��l�u��u։�-fe<\�n']��%��5�ғ�S�g(F2� �a���K]g+	j��an�>��O��wpn5$��u� ;��i�O4��8��������[j��ӷs�ޫ�8���H�܆�ښ��L�+�X��x�e�
ӳGd��:>�mܾW,�b>�ڵ�Y��N[��<� ��d��u&�ٜ,�s����7�]�zNk�)����H�n�Ȳ���p9H���t2R��q��O�<V�˱���Z��b�S%Yx����Q�� e­=.��:��,�A<M� �ɽ�gJ�BMo;
1;س7��["��`�EޞD)L=�r�>���G��X.�39��9�	���&2uu&N�����L�*Y���%�����w6�,��P���a���)e��lM���D�V��
�������`b�O�(�o6�m8�8�.���H�A��.�h�$��;�4�_]�i�^�Mg<�WGȵ�Yqrghi�I��#�)ٻX*J]��|;	���42�̾/@s/ƕv���M���J�(X��u�#���AOu-:���S2�P}�Lji��*Q��Xoiƀ�.���D��@�u�Cf�����<+�=露�e�X��}v�>��p�Vo�>
��ou�3;6����C.���r�V��v�-ҭ��f�L�LJ���
�xf��Y�{KC�V�ngeu][���o��l^Yc5�Vu(����э�/u��e���.e܈�8yX�v���9��]s;#̕���B�v+Bڝ��;��j�۝W\��� w��	�q�5v���&+V�*���{�_P�U�(Khs�[��rq�a���]�/����9��y�'Gc�\e^7H>4vK��\R=@'�|:cͩ2*��4N��~�ɂ���|m�Ui6+��Q0>"���W�-`3�7�f���) ����V�#����B�T�!�(��`s�P�h�@�>�W6h�C�8�ʴ\��\>ن��2:�	��`�Ѕ����XN��S�\������l�����ҏ���7��3=D��;Wi7*u&5�����d����X�7�ѭp����Ht�%��34�:d�Anq�.�ٯSa�Tk�����Q�6f
[��J�\�ܡ���	��\�>�˭v�X��t�vC���]B�ٹ;f�˅:�]ݒ�:{4ͩ�W�pl�^�g�����:�=����Y6Rl��hQ��L��YB��&��D���^	d%����L���h�:���3��`���r�ۍwε�u�:��<ۻ��GtU���J�Y�)J"7�!jQJ���ϡ�ޜ�Φv���s�̚�qG9_N ��7���˹�w�XkT�|��Z�b�t��U��V�dX���~9�7�˯��翏߹����BC�$��Dz""=�n|�����6w�Z2j2�(=��sh�)�t'KG
�b���}Y�Hj��1��F�^�f���s�� �*Ӳ�6�&�7�k�oe�K�[mk�.��82Im�"dΚt�AhBN�ʓﴓˮ�q�q�̮waZ]l���|�R���c��J4� �Z�l�-о��N��w�;R��tތg+e��qU"�ᴱMQV���Vv����Y���7o��VA�Ǹ�gE���Fq'/�^��x�s�f�������N��������Z�\o�����X�W�]��R�B�;�V�g@�%ɠ	��t-k�5ʼ�+.X� �+�l��Φ����>���U���b�i^^p v�k/�QY���'U�b��Z�vT(P�+�EA��}$aAf�u�������+7*�K���bYro�wo8�c4k�ia�j��C$�x��wC��
����,�s�2�Z�,�6G�
C&T:��3Ǧ�[i�컕��'U�7���LGV�z�Wj�[�W�]èY�!�HX��Ǆ2�+�mtWWfRm=�N�e,'�sUF��:�}��3eX����λ�;7�.Y\z9������H���j�,�]�k@�w|Ƚq������B.r�AJ��Rز�v��7�:([��'7P$I���^��e� MEe�����i���ohO�V�Z�KmL��kh����vM"�ve����1�m�X�-]�Fv�'V\���ʽۥ���o�l6F��q<	]����*��GM����}��S�_H�}����`��ݥ��ԭ0]��J�(�s�f�>��u6��zN���ӎ�΄/K-�YG~N��:�2ʘ�QM��H
j^7Չj�؇`8Ѭ�vˣ���Y��ug���]k�-I94��(� �g!Vd�ġ������b�P�{��}��
6�ʥ��p��z3u�{B)뎥�T��wj²�\X�:N�e�����Ǘ�jvLg5RYk۾l���1�I]e�cf5t�dɮM��t��M�Q�%o)Ю��{P�n�����l*`
��J��Y�|r�C�������<N���1���e����g&�[:�ۥ���V];̓*h&Wm3���`N��<ʈ�yw*j����T��k�e#K��P}�����~���;��iU��U7c�B��j�!pO�u�E*XA��}�C(�W��<���:[��L/���r&buW��彳��,Nm�d;�h����77-�@�'i9709���WVL՘�q�f:c��X�$�<�{���-�u��C�-�b�@P�W�
�]�a�J���l��hJڷ�~|�Kż���ĳ1Z��t�WM�L�����x#2���ZW����K�ʹ.��vv�9ݧ{�\ؖ���3n�����V�,<{O��"�3�wkT8tެ�����&���Ť�w��H����e-�����=]��tlg.�A=��o0yC@�g>���(��fTzw3���At6;sR��ZM��YL��j{Z�M���W�>z!��Z�m��1u_b}m�5���r^=2���5��ziՓ�Fu����>��7�5����3$�P:��^:�JB�
>�e7�Y+K5�w�hY�O���V�����򺘓'"�0d�F���.���Xwz�c����Nu�|����t�����Hx�Ãu��	Թe�p��-��s��D�˹�j��iD�dΠ��4� ��vqw-aγ.t�=��Y���SϘ�5��NAh��	���M�����,�y�(�c\���n%ө0�o�&����ɽ޽�Gb3�e��{��w�8;��)+��QD!���zƅ�;�ڵ��U^�*9(^y ��d1��;���[ڡ���&Z%w�A�J��<���;v��Dk���v�-�G[	��p3�U��<OUe�������ˊ�YV��t�;�X�x�����#��mT8��3_%��R��ȻM4�[2��;��Ä��������ad#M���W^ы6�a�]�3tٕ��~�kw=��<�r>�u�O�B�nL[6��������:�:j��ֲ��,c�[u>�*E`�YC����D�k������h�cN�B�� ����84�O(�N�[��u�Av��s�$]����������	Y�v�FXS�3��#��c�]4��h���3$ �vp���w2��f��p���ev@��ہ�(Hܩ%�^S���YF�ŞJVxe�\f�Ǚ|X`�Id:x7��L��wl�8����z�Y��7�dy��9-����	³5EF���Y�����T:��*��n������M�c#��A3]��MyR9Y�n�Q#؍�Om��ݖ(m�bSU�ˍ��Dˤ���ngnf������v ��Ũ��$e�������},�3KBĆv�7����̄�l�/��F������9_$���z�҉=6N���w��]v�TW:��n��`%&ξ'��Е65"�5������A��%�V�&f�"mYį���R�w1{+}�ޡ�*D�39l�+�Go���<L��������7)��t*p86oh��o�
A�]sT�[�������>�д�5Ϩ��h�:�[�u4f�Ṿ�0���1�뙔����5M;0	�<�p���2�<�.�&Y���BI=�C̏_8��������{g$q�n�vSG3���3�����S��׏zz�����ꀕMҢd`���D�.�MǷ��7��_n����S.އ�e�۰E�L�)�(Kf�Iy���B��tr�Q�ޓ��92Y�vtAMJg�8�%9v�޵��%��8j�L0��-����gn�e�e�F��*pl9g���bם�%�P
x4�DY�,Ya>�*gS��1�e�k���"�2���̝{v"��6xu	�)�˔�|59��̷k����c�^�Z���Ұ�}8<�"����t��ew]�տ,GX��e7�.��Es���O�=�g����Չ��5:o ��Y��2r�����gY��GyD��Vٙ�X	1�U�@}˒���4ɼ�*�e�N��r�G�'�]԰S͇->��#�-:I:j�O�쥒1]�/�Y��GH8��ɇT����I��CH���R����ڡK��=Y�4B0n\F�Mr�2 �f���D�VBwy}Nu��M��Pn#ظ�Y1�K��=7f4�R�Ǯ��H֠���˅9��U{\��m��<=��	��S/u�Hx�X��^9G'�Hۭ�.fJȖ�K���ʁ#��Z�쑋�Z��`���d�W;�4�	5��E�蒡�(�6�B�]�Q�H�_%��۳��.%5��;�ũ�!�t�f�4��_E��/��u�T�ڭ�ȮHu+�U��SMc�.龊ZN�p�����y7��K�9��olp������Z�6�f��n�ܳ#]	ֻs%�ґ���h˄��}��9�v�eM��^q�\�F��qjZ:xԫ�v��[}�y��F��r�	о&����p��DǍ�b�;��I5�j��������+���Nv�{�峘��A��M����|���7�j����9F�C=�c��T��:��K����H��Y:ѡWm�{e��nu`��E�w`[�L��"���aKD�T� �2���Z�n�[���MWp�y-�C���
{�gJ�k/oz5��rR�"ˠ��ɫ�����k�2��F�uɌhӱ�6��p�,Ჯ61AT��p,�����5����ɘu�lF�+5���
�Yp�b�a��oe9��t����6}��@n�;��b<9D	�:$�pM#R!��b�u*�'7��RQ܅�Ӷ7u8hf�9@wL�;N˝zh�4-��u#:��r>�͕I��8opݰ�ʙ�m����Y�����K*���RQ��9{�1��h+cJ�|H�M��+D�� ���u�H�vd�2|j�ZM[�V��GQ��������B���|	�?]�3�W��X�Ym����X��J[�DQ�����ǎ�V���,�
p2�	룢N��p�(U�r���b��]Ү,K�v1�2�p��U���^6:��5ܰ}�,��vb�Β�K�J����a݁f��	1��H̡��*T��Q2�W�ۀ�(Dx��ٺ�'���C�b�c��w���07!f�-GR���J
�����+�|�7��]O;H���A�{��^���<ʘ,m&t�fE��FQI���es@X��C:�n0n��-BQ&Q$���+��b2Š5�èu��NQ=ѮXയ��R�=g+Y�����
4�_Y��Z����[u��>��Ӛ8�7��v��	w�F���C��ACRd�U���o (+��(���O6`�i:�1
�4�nf��7Z�n���u3S����xv�g0�:��s��yo<�jn���Ё�-���ov��-j�\�݌��^6����g�)�Ml�;(U�kf<�j�b]�3Ff�޹�op��Xa��_ݣ��>.�Pw���o�jy�i��6��PbrSQ�az��u`@������d�Xm�E��cK8�p�x�S+=���.K�f�I2�m�%���)Э��Qz����VY� ��qk�N �c��6�:G�/C����F�_n��n7j�m@�a���V�7h�v��OEU)PD�ݎN�v/��,p�Q̤xf� �����Irt{�UƮ�a#B�_RT%m�b��ucQrvƝ��Q�l����.e�/pc�3�^mA aԜ�9û2��ú��B˂�Z�M����'�o
�R\㗊�;w.}5k�������l�,��ׂ*T-��E�]-�c2�����R�nk�f� �+h�)R�ݣ]Xٳ�,X�\|���T�&��/��r4a��v��@��>w���n^!�u!۲�Dz[u�Ӎ�ѐ9\�ѽ�Oi�]�����N�[i|~����}���L��+zx><,AM�Cp�d<� \+x�tf��d�˜q�v{3)9ցU�����]�7>��['4�;rs	u�p����U��[4��a���g0�#�q�R��2ڥ�eS���}B��C�	vSW�ƌ�M���;7����v�E(\uӴ��X��V!X9�,V]���R6ӗ�����C��л�z�!�:{}����EA��Js�p���i�7+�52�s����Zka�-$I�l|P�����'��{'��]04��V��ы9��B��"��tpb�zE7�sa=(�}�h����|�O� ���q.������'����:&3m1J�KXoyA�.d��
��VvV�nS`�ĠU�ʖ1h�M�*� �"�\�ݹ�/2[�:�q	d6��`\�oAE"e�4�9�Gn����=��Qm��V#��y��H�kO
�Ѳ]�'wRzwښF�Z�*U��@�Z%5���������P�ҧ�Q��lpF���ثy@�ڶ�eq���T���X�w|�i ��ϵ>��Q��К�u�ib��;x\o��_Y�]�Yx܄��_�C8)�:u	^(�f�5�v���>��[�\�c��t�֑V9�i��%�N��f�o���e1Ֆ�0�N���1DY��,]<�g�T�߭��;\��Ƀ,U-l�!򬮴�W]�����-��-P̖�N���M�k9u��3\陂3��Sqve�(-�.�7�,Ң�dt��\f�ob|3pI�h@&w<���6m��}7�
��,�+���U�l��^����Z�W�k����,Q3S��(
��M�7t7�h�}1��`�ϴ�}Q48�3gnAW�����cH������5��sF�!��:���b�XƓ���)}d����&(5�8�crٕ�ְkK�r�6��[L^S�g�k&G�YT{�<��"' �]��f��w�f�tJ.\�@���Ne[�@��C��:�ɯ�Gu�땷H�\C�R�{3\��35����]����!*;)��@�qr�&t�Kk{���D�����ٵ3��3d�S[0��	Mܼ۫E���rfG�]��j��쎻�����^'�Jj�&��{޽}���M�6�_VrE��Ja,ݙf��^�X�4&����v�ar��t#�\�*�)��\fNID*�^g_�W�����E�;@�]���;��(n]��=��T�s&�
O��'tv5Fw�rI��.&��K�@��tsi�;����M:�s y���ݣ+�{}r^��WP41C�����(��)��7!tS,�)�]�����70��\h��k_"�4��"��:H=7��7�*�eN���xK]��i��X�
�u\���M()�u�:%ʁ�r���;s��k.�l��B�3�2�%���
g�՝���NO���^�Y���MQ�]1���{�+�_8�w�z�hY�̏��%Be㹀R �M��]�/��)��k�� �Y�J���Y�����v�	VG�	���B�����٠�Q]��=6�V�{;k,�Y�WY�+��N�תp�:�����6>Α��%��Y�c��(*|�-R�ʃ�s:��`��mV�B��x�+�#��l��%_uC�h���-Q��-��W�h�J=3)Qȍ�.��K�gP4T.�	;��3K{]
8Jި:�g*T�iՃ�1e;�Σ*m��"�}-.9M��$ ��Vw�N�C��rP�|7����CcY{\ɲ�<1@�ئ 	�ѕ���ӴV��`�ٳ���VDĔ�u7�,����kF�lf�w(`
꺗��Q���
��|�\R�p<G��G���G���ZI�Bi`�����,gIoU�X��4�-6x��A����x)�|��W�rb�����u�GWV2r쪓���kj��9Jڴ�]gq�����br��t�^`���i1���沝�ᝓ~�3V�軚�p���M[qQ`�l8��<��އ6��t�&Ԭ
7i�A���H�ohMIVWS��T���䖑�;K��q͚/��	����$����>��/z�z���(R|��3��'RƢ�W-�l�ʗ���7�׵W(�����%I��#��	,ۉ<ۢ�vn������ghd>6�.��_>\�r=y'3�W�0��0���BX��2#���;^eqV�Z�&�F��4��3�Ws�WIur�%�9t���'S'9_�O��a�|��fԴ%pC����]�wh5f�+�c.�&s��%9�סHڱ��F*�뭁���0E(r�p����g1Fp��l��|��T���K��j�=��5|��sm�OC��""�er�L���wS;(�᫾�B�
��˺R�Hfs(��þxy��+L%��w"Eh*��i(]͓��`|{����<=�#^=t�T'\%>#��@ۺ��Z��qJ��Ǌ�I^d�z����1����Z�Y����
C�v�� ��_�?��T�;gnq�_��wM�2��sꃍ@�哬oV8c��ڊ������G�K_���`i�Xd���V�²R(UR�(*J�A���EP@P��bL`�Im�$X,�i28�UX[H�ڵ��5SZ�	�J�S0���,�VT�)D+-T�*Q�I�q%JZE�$D��YAJ��
Ha����Xc!��PuJ�1B��m��QX�
Y%a����*���%a)R� �["�`���ڂ�`Q�i����$�V�dHi��5CHCL"��!Y"��L`V
iӌQE��
�
����PXc]!P�� �Pդ+$��VE �2�Qd]-�3V�+B""�E i�X*��4�1f5����L*
DB���Z%f�B��4�VE������rgD��8��������ȶz�5�Dd��j���v;�/�Ŋd��o�L����Yۇ����@�.G��[�*V@��귗*�t��٘0���̪R�R�BuJ�s��_K����SIs���<������ʼ8�X����§j�t��oa]齨�����\s�ћ��^<��/e^U�r��)ۍj�a���	��MƸ���=i�&}����~A穧����g��*~��h�Y���{��};{k��5S�ߠ)z�掌�i��\���,E��ڗK�*���\�V�v�x�?{�߻���W�r�:���ރ#w���`���Z���H�G��u�Lr�W�9���⑽P��s�!9뱚�k[Zyʼ�9Oӗ[p�Șx���%U�nc��-�Q�xדe���g��;6�s�X5��v]����*#ew��R�{�3i�'�惧2����yu�]��
8>���mFfR�C����olw����{�{D��eݮZ��6'�gEKkN�h̾+��qL���n�QU�EG�V��/ۈd�*��ύIEv��.��q�kN�=�t�Q�
�$.T�[�A]w����V�h־�:�w�+m�'��t�:O�l�B����N��:���^�����ծߗ�[�X���6m���nv�s�=Cvw:�ĵL�{	�t�p���/Ξ�����O���fF���qz����5k)m�|琹C��<�09��`����re����.]���*�{����� 9�O`�������P]Z�s�v���z��"�h�a���U(�Wj^nK�}�nc�11
�^
թU_k�k�N2��ҵ�����5���ޣ��)y�k�u0r'Uo@�=��r�VkBh*yʟ�� OZn�Ԋ5�eoy��E�.^^m'^��YAT���m���b��T�P喝[�zL��^/6�ʅ�CA��(V���er]%MC���7�ԭҵ�i���ͱ�4�6�K3&q�}QӢz�gr���J���¢3T򕮞kU��u�^ѹ��9�Ȗ���Ck;m��ΫY܈-���]�F0'^����������V^���^��-W����B���Uғ�Y��b%J�p(G^���j�H�~;�T��lm���8�X܉�c�O;)`]WLE� ��te�M0@��
����Di+q�ݳ�N~X�������ì�V�%<���y�n<˚K���C�g;�t'٪C�ٺ����Vڬ�QلO��x������s�w{�tU+��#�=${���pR*��.���e��f�6�ؖv߱Y ڢ�v�b]f\n$��{ƣ�S���m���7r뵊��I�'<{�&xj��>�=���w�my�酃�×�/Jެ��Xt7����yg+��!�b�T/j˭nk:�ĵL�z��>x8F*�"�mq�9.}<��X�z/�#3oE�w�Tƾ�~����S�;p�If�EΫ�}k{��4�����WZ��}@�x��ٌd���G�ޅ�UoVp�"\�N	���oc�W����"��͈�Xj��=��{�gؚ���F�nɊI�͜�]�1�X"9S��r<��ˇO	�Y�r�d�k�g�'���g��:��v����#�N�vm'sx�=`�ls�$�|�����kJ]�{��t��e!K��v�ڭ�|�7/�ۭXkN��r����n��)m,��.V]o����t��K�+!y���y*`�h��e�����>\�|��.Qy�Qm*�}�A��J�q�V"3j���T/3%�!A��O{�i$S
�v�0��j����ؗ]m�Z�z9�� h�EާM*�螧�/+�,�<��~�S�su�ڏ'n��V�Ɣ�Ԯw�7NL3�����]Ŀs�vmo����a�csTƩ;Kǟvx���O6��#�Ty�y'i���:��W+�WO0��b(Tf��rO
q��d8 c��s��;2��r�^I�\;BJF����2��d*�Eb]hu1X[R�Q�E�s��,������東>)Qav���]!}�I�)��Хډ;x�bS�z�9�+��z��cATK�.�/&���^�F�x�������u��'7�y�|W�m'ڱ���U���݌���G��ѹ��'ޓ��ܮ���nFiR�W�8�n��������P�4xzVl��οb=��t;�o�ø�����+�5�O�+���b+�wg�ݩo�`8 c�'i�y��`�4s��8X5���)��4� [.)w=��ە���C;ݽ��kT\�v7R�PR�*[t��9]�jn��^ѱ�6*�T��wY��	�f��\��D΃�>C��멟r�tV�����Q�����Jͯ�*k��x[kkE��L�Uo�j��s����|״ܦ��������gm�2�\��7��J���w�xN���ÉMU�&&:ڲ'֝G;���/�ܳ�]Ww��nv�UVT����d8N,N��u�N��6P�Ҫ�w+��]+�����t���-����'��<'7DX�8+]ks;k7�3�k��ӄF^\JY�)E�J�mk50y����SЪ�vj*f:R�x��]ХY-hͨ
3v�м�yn�2�U�*�s��7��d�!+Y `���u��ٜ��� �����%���j����|����&���!��i*�{s������N����=�|s������jr"�Ot֧�;�M����픕��;���T�|�rN�Մ�9Obk���z��YG�ϐ���E`̸g�r�5�vweN�Y��ZG�U��/��� -=ժ��+����˹q�/��
��OY��֘��H7��u�V�4��'��GIVv-ݜj��Q͝��F�eͦż�92�oJL �6��p�1q�+�Q���R��>��SJ�?v2��[�r�[��w����OYgN�]K���f��_#<�W�Ī���[��n:׼Pt9
�����G������n�9׃��qۺҮ�%}��)���R�J.x7��yً�8{�ױ{�
8=�ѥn���{�8kt;�z�2�}ۖ�wa��o��u�Oy]�ʘu��.9�|eY��H�s�IѨ�X�LO)�)�6��mx71�J�w�:����>�\q��CiTuh�8v,�5{�꿁��� Uz�bf�	S�P�7�*�1{O��_xm�i�0kZ��kBҹ�sR�K��*`�����.i2�!bt�[�y��Ȓ�)5OVĽ���b۸*��C��%�����(\�GC^ˤm�JC�nL�I�-� ���V\G=r��xm��t��7�g�7Qv!�}HM���
c+5عH��w�9�Іu�*2�@�a���X,_;�r� �Y9�b�&��0$_'�p ½�	����J{zteR�O�X�l7��N9Ju�WH��X4�@Nwr���-t��pB���滺 ��O�n�J��m>����rMjwZ8�y�n�;�$�OZ{~�Q���5�������)�mN�l>��+72-�@�'n��;p�F='�͝��ɯm�Pk�������?�{;�N5�D�=;3zuMִ6�+j�u�3�t��l����n#�h��{���duE��K����t�a��I�\+���3��a�F�Uv�L���ߚ���gW,�M�LC�"V"�E뺎JySw��Eu���V{�y�ҏ��3��d���b#mÜd�J�{��x���J�-�W#��.���9�<�ʞ�g���_>5	�>)^��.{������9O�>�ԊΫu1_g?L��'�畾N[�u�{Ʊ��0��W`г}o)�6���v
ҥOM�83c�{���ej���r�F�Y���m�1ѽ��&g�55�n��~���wr�N^����^������]z�pܧ஋�w����1.�B�����e��D�i��ՠ�V�ld�6]lv֮T��`:	�xї�54�Iq������cD�W'kޞ�|8��xəc��\�+���;�:�،�+��v3�܆�l��8�k�
�j�e�u|k�TF�G��q�]�~�da	��v}�+@L7����; 9~'��Q�(^��t��O2��ϩ�V���}�@��ϵ��xK��p���5��V崅���T��.���o�6�a�]Z{W*짚�4V�gn����ꦦ�1h�5��-4p� ��Q���t��BV�볮���<�b��q�y���a��d�
*qū��A�^%W����$UEY��N���<�t�^\��\f�&�V�xA��.8�^ʫ���[/} \)1����/Q�y;+-c5ѭ�N�+U�s
��Fqp�M!رn'���Lt92}�f��������}�W�3ꮾ��sܞ���isW{K:ӈW�b㕌uMx�Wn�:��J�P��x���J�k̒x��-<��-�����ηh�_����2��d*�y�]��:��<���<S���L�͸�u�jĸf�L���1���}ז��Qg�ln��Vfë;�:5�.��Z��V`/u�����|����xH��h�R���'&�|m�E�6yz&L�̇k+�3o�:8�y�<7�x�WLݧz^Eg ��@������4K�s�a�'wd�(+Q�{�9�	�oo5�	��m��U��p�J�@b�R�i�~SdOc6�ؕW�W=��[ε�Ƃ,#���Y��pe)�ju=�����>;�a9�8o�/r�O�1���U��U�H�{
B}�z�k/������=���3J�eW�9�O8hw���L��w�4�nɂq|Y�8����o�J����30P�f׊��9jX�Td�=s�Z�����|���/�uϡ1-�ѱR��ʼ6�+����{Q�-=}�^^I��2��3+���%�#͋��>R%&+t[�ۚY+��i�p�WP���ZՆ��j3ϣ;3�Q�W	ŉюv�j/)�QٯQ���kk+�}��'���.9�-����%��*�z�����ɧ��Uծd-�C\"7�8��-�o�-���qq�kژ3�n�_O^ؖuu���K&w4m�X��Y�ƅ�ݛ��H��M!���׏����_��wK��O�9AVNb� q�D�p��Z*Vj��w���\�cXc��'z�3K�ӹҵ��6�,9���5���-����]�g�;6pK�n,��n��W�7~�ٮ�+j�����k�Y�g���8Z�^�3˸[L�}[n���|Lš�5�/6�#��+��8���w�*!*�k��������o�+o�=/<6ac&��p�3ە��&�0q��)Oٗ#�~��W��;�Nd�U�޵}�<�w�$m�t�=��%`���%W��t�+6��"���N뚘�\��tC[��h���坮����oZΥxm�Zy��t�:l����Ī�ߧ9ҫ��?
�K�7��O���Ťz{����������O�����⻖����p#��>5����X��uX�~���.4����L�N<�^��EE���=nz����}��ԛ�ͧp�:��Ұp�r���x1.җ��_��ʜ�G���²�xy:�(����N�N��z�p��\p��1�c�WK��-u�1��{�uܫx�̝/�v�:�z�,n�����5�S��0���	��y}�v�m�#*r�ΰ��ͫ����1=K5��pH��g{T���*�z��ɤ��n���f�J�v���� �r����T&�Q%��HvX�J�d�����Y����sz�6:
�t���~ж��wS�|6�Δ�'=�8٫Ł �`�	^qN'���Ĩd�Q����б��
˻Q`d�!��ST��c�.
.�$��7i\�.������J�4d���R�Z�[��[0H�K�vݤ˼�l���!�v�(��S�F9olkV��A;y��R��2
]S�e��!�Db���"�1dɻ���:K���ӳ�G��1�l��	r�[�)���4��Ay}�%oX�J���	Z2&;60�Q񣣃}��r�9a��Ew"���v�è��/!�����ژ�����S���Ɋe]^�ՠ����T���OWT�i�h=7V�7�%��u2���e�;pS�ju+��k�b&ŗ\o�%���A�|�S]Sr桂Ίq��%��]R�F��#Q���oTV$�#���:ݬ�{�������H�w��t2�Fг����5� �:�'��Z]Ȟ?c[��[t/1(Y�����	�ٽQw`�*��f��V��t��
����,�>�/�}F��ծ䕧)Z`��RM�V�:�J�[�YW*X/�*Y��v�I	D��S'Mι���F���VU��B҇8=A˘)]&�V�	�@��ǏN{5!iAFԺB�"[�^��]`�a<��@뱒�dV�-c1ed5׎�Gu��]v�9� �U��v���\nV�sz;w�G�m���gY��v'I��wᮨ�cz7��D�� ��S�>xo��÷]X��(B�+Ftw0T�p}6��/V�l�M[=Z�}Q��wM7�ͷhn5J�u�7���ݛ�
[Z��E�����/���^���u;���-���Ye4^ݾI���%'��<�ft퉩��wZ�x;aU�Pv!R�I�w'=���'P�)���4mB]pm���t� 4�(�et������ �E࣡<a@V�On8uɔ���X��SU���z�,�2��4i/q���v�8n��@��p�Fi*i���qۤJ�@��SG5�T�)ͫA�Co�C����®wv�֝���Y�h��B�4+:����s�]�q�����Kn<�E��q��8қ��|;�ӓa맱�X��*���5)ܟlb�D)� R�z�Ŝ�`�����֭��9����y3Z�Er9#� �5��D��EC7yɲf�I�"#"�����,h��
\2Wk)�x�p�̡vp�gU��0A�;e��m{�uk�ށ�P�z3Y�f}u��P΀�����b21\�t�=o-����Cqfd�J{�D@!P�$�@EO*E�l�=d�"��$�LC!��d&���IR
i	PXE"��X �D
�`
E%@�&e(�)X�%E��1�YX\`bT���b�,4�CQHfYT]5 ĕ����Ma\L����L[VB�(Z�h�F*���kk,�*�±E-�l���l�VA�`Q�t¤�%b� P4���2���)+$��1��ʣeH�@\a+1���B,�bJ��!X�����iFH��,"��*�
��Qf�+��)+"�SV�f!X��DQV*ņ��YE`�M$���I��#�Uf�2`��݌$��Ck�t���I��q�ˣ.�ǣ]��[��7��s*6U����tr��Y���-��u��*z�\�T]iIf-I��b���W�ޟ�j�߄�G����0�J���;%�M�X��{:e�ӷ۶
��&cځ.}�7
	M<S[Su�U�,�x�T���tV��c�z۞]/�1צ�]�&���i�w>�kbֱG���Y��:�:�`u�N�B#o.[�9Kb]�ǒ1OQiߦP��z��:�3�Jb���y�VL�1�Pe���܁1���n��c�yԱ��*y���j��hN�C��p�c�g�͚/6��p������%zM�����Pe�z<�<��D5*{�f�zu�"�+�gB����6� �u��ͻ�YV�O�ic5o)Z���f���)h�0-L�i�}
�M���:�"��iй[�o�\�����¯]׹.R�+���tӊU��u�N�wU�z�*CJF�u��2�M���W��_u:�+ޠe�*`�դLzݺw;w-�ĴM"��f�Ғp�1�+]�e��X�����C:D�J���ݺ�f�ޱWOj �@�v��aP[���/��34q�6g����-�Wx�\�ԓ?1�����TE�N�k�wNB�ގ�]R�=m�y���&����0�b�{Y�-g���&�a!6�C���e����[T�f���}�������ŬV�[�VFk�+[V�q�*���Ϋ�7�yT;�*�:Ε5,u0sq%VI.�[2��^�{���"r�,�mEgR-K�:�C�U
ڳ��3Wi�I��DԽ9~���z-Vf��FmAy��+_Kw!V%ί�ع�x�����s�0�K�Ɖ���.�a�|�68��7��3�w��é�=3��V��zS��"]GYA����j�O�nJ��ץ��r�q&���C_��j=�ڌ���8�ӕ�cQx8ez���8T��f�W-�˻}��8�ov�@>��Ϲ�0�ү8��I�#6s��9�F����w,r��b���/,Y�ʩ(d�΅>��+}<��^��Ҭ6(E��[ܫ"&|���C���ҩҵ��{����i/�L5Nv��F��M�c�(*��!f�7j�p18�0�	swoU����gAk,U�c�Hun��=`]�˛%8s8�;���g�l�w�z�Q�ǬK���5���RU��`>����[��^R�/ʻ]�n���	ۊ����a�y��.���~x�{��;�Kͻ�bk�����^r��5��w�G�h���Z==��r�OWw�5\U�w�[�c�k�r�5�y�%b(%�}x���� /LS4t�x�g�q~�2�����]�]n�	�7ZY�
��J*AɕQ=Sy��Z�H�G������弭<����lO�EW���78T�+��-���T�[�[�-yx?.���'���:׼k7wT�Ҙ���3�wN�}}A4cV�Q���Δe�Wyʳ�3jS���z��=cy��u�ߣ�C�f���F��]el�{pS���1,^����5&�ܭ�i�Ϟʜvl�#�y��5f���Y�IX�;-�.��Ŵ���'�=\��s�ݝΦG7Ӯa1-��T״�o��</����8~g��ч3Mn_u�Μ�e+n�Ѵ��쫙t~��z���a�I���q[�< ��z�F�.Z-�ںÍK�<�青���P�SGcE+|�������Q��⾮d���4�b3y�,�ŵ�xe�=����>�\�RA]��>1԰<m�Wt��f������H�b�SD���o�z��V�zR�y�rw����pe{w(��v]�VTj2
PИi�)�՞�bͧՒ��B�)��龮ww"���i��8�/^e.�q�<����:�e�Բa�vrΎ�4�;��W���f�mZ'8�H/W����}vg�X^8�=���RA���N��^ eOZ{���}��ymZ/8����7�����'�d%�u����P�;�ů��/'Kͻt�+ʷWfv0%W}}L����~��F�]��J�z���_Ȍc�k�vޱ750[��pi�[���-F�O�v2�Fk�r�Q���Y�;��;�>I35�eEwv�is��Ud�p�:��H�hRt����\�9�T5�ȹ�K��4o-F�k5He�u���+n%]+�M�0�W�W��Nv�;Ϯ����G���
���s�|͉���3��D*���+�dl���($J���i�k��കP�{�%�˥Xʷ�]ݜ+�	�z�-��V]�ήZKF���I�'��k:�=zq�:.2��}�v�3�M8S�}�r�g�|�l���C���r�����!�3M��%�<avE�[V����F��%�g��J�è�4$�gR�B1;��9�/��������6φS��o��u�� ��q�8���&x���}�{҃���ʘw��g��S��ms���f�<W��+�ݑX�͠�gJ-KrvWB�	gK�hے����W����~��i�=�7�[�C~����T�j���K�G���@s�a������AĐ3�+X�ӷK&ݼ�u�1���7�=���E�nd��̾�w^�f	�a@�I��@o�r*���P��]�
t2������⹢���H�N=��v���q��-�vU�W+ ,�W��!uX��v�(���� y���ҧbq*z���"�/I��M�l�O�.E?}=q�:�FO��S���ۄq�O��x�J�<]z��hv���{0X�H�NUj�Eck%m=P�5�z��s7S��x�xo�p�M��|�q2!��vAR����D%����9P�ͫ\�n��l��վ[�lr��NH���Xe�sہ�퉈��4�;tu+J8���Ev����_}��YnO���PsaO���8�}�����:�>�<��ON����6nJ�u�� �-�R��'ڪi�y\���}������v�6�t��!J���kw���;�/�Ǳ�:��ߡ��YV2"�E뺎J2o���NЬ�]iN̫\�we��v���n��[p�Vڬ�^��&#jG:�XU"���<���s��Sj���;�mA]�{�h��P�s~���i��x�_`�gQ�w��o-���~�L)��:�g�M�t��֭n����Sf�se�ۈ��5O�9��گ$Ѩ��8q�,��!3M�wkt�wp\q�����\���V]ksYԮZ��Q}VX��ts������aO�����JӅ�ؽ�=wet������8F��^�عޯ��$u�9��%�AV��>�|r�T��_�kf�o�]���7�vg�N ��ܴ+8�CrLk7�����=�]�TWY��+Ep��V	���Ft5��'mk��\�xx�-	���i�Xt���\�Z�&�qP�m���] 9g�{�T���:�.>��g�t��8��/(��WO��?}U_|:'VN��;���y��N|�K��"���۪P�����wZ�D��w��B)y�}Ɍ�ƣ���'��ԽE���[F^	�v\�XzzӗڶK���w;�'u�>���C:T㚰�w�&E�Oe�������}}H��J*.8�[t�0�y���	�[ݬ��s�ٔ֬�V�t)XK��6��ݷB����y������[އ��$���mY�k��[竽[|�=����u3��<��:ֱz����V��'�+� ��wX柱�3��+n�R��{�޲�MWB��fN���:]�R���V��u�Ɲ溒�8/v���*yq�:�'�nВ��n:��Z���rp.�Jj�}�ۈ�v"��ZWQ�Lr�I�v��tƔ����\��ή���g��K�TmS8��[cx+�w��>�s�s����1tMQ^K�+&�t�Ӆ���w�b� v(9-���)��ת�q���`H�V�Q�,��a��[`*�݄���ڔ��5�K�ѓ��GgPm�i��-;���K����e!����M�D
��E�D�ⱹ֛�P����ܖ�VK@����謁����e��?1]��|����Nm<�?/r�O��&�a�W�]x�阷����>�8��8�������T�=��]����9hw���F�];�Fs�kr��m+�<��0�p���x7���j�0��P�����]2Q��4��OlP�����S|.zhy�%�/�sU�Uu���~�]|�.��eƼ�/ �y�W0Z�t�ʹϼ&(b���+l��o�����1i\�8�Y5uj��.��g=���!CA�o*Ll����ij�Y�g["z���Ȫxk�V�Uʼbgl�rc��y��ːf�tw5�R���>����f�:�"%���{��_���/2->�C*p�'iڸq�1Y3�f���f�l��>ڴ^v���)!^0��XN.��n�W$
t�:����������ۑ]sL[��2��K/���Y=���{N�{ҙO��� E�m��jk�z��w�(
��ʺ$	*���HZʭ�Y��.Vz<·�:���<�C���X�6�0�)��1G�P��i��(w�ݫ��|]�'�1h���	��9�����Gv��	�֒R0u�|/5�������4	�y�Xɪ���z�X��۸��ʓ�3^Ժ���ľP��s�Tj��泒w���������g5��Z��KM��ko�2��VuC�"V"�ZwQ�O*����l�҂\#���F�����hLF�5B��+n%].4FC�m^%Um�"R�x��_l���&��V*ռkɲ�XSavE�[os��	�8g���(g����@T���ӥe]��s��<�oz�1>5�Ʌ����S��}ƥ��9~��p�ꃳSs�a�Y��0*�O;ʞ�E��ï��q�+(�݌�_a��{=����=EZ�sҏ����21���s��Y(t.5�Uw�y,�=�B�~}�J��hVNz�ۿb������7�-n	(RY)�%ce]�x�m����݂c�Oj�I�Ӌx�7lW�N'�%�4��:d�'(k�Vuv��s����z��ӏyӬnLzxTXsb9p*�3�S@���Q����sH#e+r����{�n��"���gvU�\�e&z�5��/�;��N��5��LNٱ�m��3�+�[7�{�08Ш��Ι�*�������Es�jqN<hP��:9o<TK�"��7ٹT�׮�T=����F��sP�LR��U�T`?,S��J����-`u�,�1˥�^J�;�1�F9/�:R��We����ɫܜ���S��VJ�|/+�nP8l�d��1r�ws�@��{C/e_��q���<�}N��zK�PN�F2-=�3�$.���m�ӈL�^A����;O�ok��x�w7U򝑚�ڄ�N���z��.���N�duz-`��X�[�V�x�[�ž�K�]ʟ5w���8W�a4q�tΩ�w�YQ�t��X�E��M���Z�q�Cy��p���Y���7�#t�:��Z��u��V�G�7o�r��R��5�5uW���弯��V��^�ْ�U�hor2$	=�Y	f�.Z{)�&;�x�Tf����yֽ�Q��)�#�֊��w��0�����K:�ˡZ�QF�Q�ZSN����-��S��H��{a�c�+��7/6z�/�`����K��g-T��nP張��q��~뚧U�g�!��&�x9�7L>X�Mm#>�x��C�xۼ*�W^�)z�'x;C�����ҙaW]�pf����N�i�n�6s��֌v��s3�k�C
 ٙ8g�˱����H�j�C���vB��c犆4c��.� #���0�I��)x"��wׅǘ|dX2Íu������D������Kb�WkEk�/B���n}�檙1I36�J��N��� %=���A����]�^��.;EF�u����:�l��3cw����2i9Y�e��c�������Tw�*v\)��Ǆ!�UK��ugӲ�uq��խ���o_e�ū+��T�'uA\w�����^"��j��
���L�;�=VԵ��q�;hsEZ[4���p��X���9�C�-�	�Վ�qj����ǧuM��#�f�!�cM��Gs����]qd��u5�ы�bz�됼F8��~��ْ��ս�3�8nhUz�݃�)o2�}ʃ��	�U�B���q��ƒ�Vo�e��dڎ���ԛ}��l�/��&����V;�K!��=��b�V���-��),սׅ���݅^��K�wk+��eXI�O�Z��7j�w9�*���D��ʗN�:� ��O��I9�ݎ��:�EXo��ce�*�u%ʍ�1֝h%]j�5H�n�n��Svg"n��9�U^��� ��c�⺳]P���\4�٘_?�n�±�QU��i���Y�]�Z	@a��u�#3��5/�h뵒�1v�B�mf����k�V ���JGd�������+�>k)U�c�bg-5+����i����YG)��JV�!]2�֬�Ǵ�wh�B��hjU��9���[W�:�jM�����k��s����F,�VF��#;z�M�P땻+i�3v�ܙ�6#���Nj�āڰ�V�����8R�����r�<J�W>R��ܱ�#o�K��G��q�}��@f����uG�D�wĔL���G�C��g��θk �k�D_o�|�.��:�����R��,:��h�wUwu[䊲bo*�F�Q|���@vX̝+8�P��Х�_l��Y��i�'z��g�����mE0ܝ֦�"q%E%��t?DÛ��:�f�hvР�5�]����v϶S�:�&�l+z���mE[z�(6�����
'82��co7�W���Y8�$*�M3��$hu�٧�N5�Nuڮۭ#�km�x�1���� *R��}c*�;.-O����3n��J��\�g���͵�k����۶��0$�p�%s��\���Yð��H�j�^uS����s�?ق�Ai�b�'��^�؅�����%�0_^X��yJ�O�Lf��;9[]]�W$Uܷ��\Q.�7�v]T��E��X".$�
�R
##��̳T"2F �,R��*�Q�Y+XTg�1$ӦH�,� �Ү0�
�$�P�TU�*���@r���&���%@X��0��0kT�d�Z�J�m��X�i1�k*VC���Xi���
B�UA`��
��-`�
Ll`�J�`�E��Jъ(*�"�P�YF*����H����L�UE"�"Ɍ*���,Uq��E�L�QDT��"�Z��Ҍ"��,��b���i%�Ĕtц[�4�ƫ!��Dd�X����P*ȥ@�Z�Ī�U ��Y��)Q"�"*0���P�c"��c(Ȩ�H*���XVe�d��jً1��Ll���[���Y�.�N��ͥ}�@�q��|M�ݾ���ZߋW��l�kϝ˽"V�*���y&?ꯪ��Jې����7o���o�ξ�Vz�]�b�dW�;�-�s[Gff2��q6����=/�^��x3���e��v����oQ���ҩ���gb�[غܕԐ��pȩZr�]���S�T=�^jsF���PM��]��F�ӏ��[rSe=�r%T&4Q|o*�v�۶
s]�V�Uùjo���u�p�FJ���\�����My�U�p�t+W���8�}7��W��ϗ�fT�z�8�'F9ڕ���U滽.��ZW�r���6�����2�]��U����4&:T㜛S���z����y�6��~��P��Ҿ�>�D�+>t�����Ow]�	��D^�ො���ߡ�1�O!��3v��^W�Y�����~øiJ���,�[��{�{�1���U���i*p�O���+�Ms�Uֱx�^��Yᒋz��#w.>��RI�^y�,ǩq�8y�e:�`ޣ}��ˡՙ��*�{������z���q�E�AǗC��y��k��Uw�i��F��wuuH���If���of�p�=��@%a�ݮ��,|R�~�{��q���')Ba^ٯ�9�m�5N��{�z����p�:�I��:vu��m��lr�L5��޺�ܩ����w�>=w�4׽S_R�G$�[؛���7N2�R�"^"��\�r�W	�m8罾���=V���V/5
��OǙ�8fۂ��f,���<f��*/T���ͅ��U��ps{�#�Y�^PN�(.��m�3��GҵH�V./����;���|�~�qތj���=ׂOR��]�K�NW)xz+,sߨ�]�y����Z���-��[�v_^���_Wy̩�����	�J��lE���\O^:<خN���߷h��	�t���ߧ'B���lwj��5=��=�����/_�3w�-כ^�*}�K�y�SDVL"�M�Cӷ�UN��c��o{�\-�����u�ؾ��G��*4{U�̜���㗰��f-}Of��j��;Ӻ`��΢}���a}�KQ����f�s��[i�T������S��{w-�z:��x��N]cg
&	$U��u������ʺ�0-�b���=�wj�����!�ܸ(g dv7B�g�ꯪ���Ӥ�<���Z��ڿz&���Tt�,��s8�l��W��FJ�U�)k�hM���������FmB#�/��k��ܻ��߼�4��;�[�WF��D/Gg1���lަ g�}E#Sl��x�,��F���X����������ց���\�����<t<����*�v����6�r����rv/;8Ӎv�)|���=��r�yQ�ᴧ��ZAhݖs:�U�W��X��yJ��onί$�*z�y\��s��sv�����s#���+��FB�P�N����@�L�K���y�k�w]����ö&
F�5B���t��[<D��6��ie<���z�W��&N�O=��˙3WN]����s��G��R.�)u�v���9�=�M��g1m��>�y��Ob|j1��!0��_`�+s�,;��g-�ʖ�R��].46l�/�r�I������)��6ܧ�Dܽ��v��'vnB�ڵ���ڎbTp�A�I���~;�=���S�QE��5��}Y��_M��մ��ӽ�Ig\ݤ&v���rҸ�[��Q�e���������}�ڭ��7��Y���j���l���3μ�t�`�D���j�]�u�.��^�^�̹nEn��A���W�;��qQ�\]d\��6��}���oR���{^��[�ÈK����ٰU��[Oqҭ����{{U���\8��Ay�xLb{VJO�9��̀�W�ɋ�-��V���[iJS�4��	�MQ�^zC�C���o���s�d��\z�jJ/�X�i���b��l(hg�3�k�G:�ڼ���h^�
=�z��|��\���V���1�	��C�<���c7N7�N���j�����w��G�[~�o����W(d�qLt�N���¦c*��7FW'Բ���.'PΑ��ڳ�qY>y;*���5�׵���q�tD�������z�F�x}�7#���q3hwM)ͷ7J¼,?f��+إ����Lut$JU�a�����@PW��`n���#�33����+A�Y:u[Sz��.�C��_nԡ�(���w�엹]h;;}�����{��Fh��'X�g+��"���t�%ϗu�j��s��6�8�[��W��]�fe��;&7�v�PC�9n���=�u˱9jvg���T�'�q
�L&�c3�y]����=�+!� �V�}�O��8�;rU�^��w����R7P�=f��ϰ�v�Y��2�y�r��N�Z��U[S���y��{�6w�"�8�ns�HAW=y����ܽ�%r�/��>]�'��o���s�����1�<�N�nV����j�Ƹ�w�s+n�Q<q��.���T��X��U�Q���{u��Գ�ڗ�F%�,G6ϱvW��P���P����5�'���^\�{)����\���q=��Ԙ��hu+N_�[�7��P���f��u6���S�]ʮKj��������1}C���9��U�]T��S���'I�[������X�o����!���.P�j�ɯӝ��Q}c�#����8��=3j2���Tz�C\'���OT�����t/�ݩhN�=����ﺴ]�����Gc���F�Γ���2��ӎ�C�v>��v���x�d�����w*�5�W�=�ݑᮭrZ��uf +m���dO��ouv�e���Hmc�a���Xn�R�]Et5����F��Oa[����F���b�p�v��Ζ���Q.�\cگj�c[�1�	P�"NcG.�L�M�����{���3aF�������]ʸÏ]�`͋�2����sٯq h8u��c�=&F�y@�y�������>�}�I�=X���-�����5�����mq�g��� ��&mP�g�{�fs��v૱�ŭ��TT�q�Ӯn�1�ۄ��O9U��'�+��\��hX"��"������y�t�z�n.4/'��{���gT$�ڨ%#V3�'O��u��IZ�ur�(S��E=��/�v������Z�.����]�/O��/zH�mW]�����ދ�82 RS���պ���`s��׾�l�Y��K�L\��W�8��]o˲9y{�7m+0Lx��F��E�!��
�ȃ��^<��UL^WS�vG��t�s�^ۘ/�|���c�=�i3S�\�N��,:m{M!���!ow.�Vc�ї傷����V�A�H�'��JW�-� �l�V~�۬���4TL�/9�G�f���m�J�!{���n?�or��ڏ+CYK��n�Ό��ԯe��f�]a�{��r喃Ų��
.�>�x*�2Z�B8�Ë>����q|�R{ϯ6����P��#b����S����by� 1�z��]G�����s+�܇d��=�u<��vÎz*B�.����i��Zj&V�4U}���"q,�LR�������zm,�"eM�B��̣%߳h��3�D�k���9E}s�;*xP���:�xn{�o5�� g��x�^�G=O��G���*�]_(�o�5̸@�+l�Q�;wFW^[s�٢�҂U����=�ɪZ|co�h�i�+���\,xR
��l�.��Z��h�J�!���j:��2KU��z�=��]g/��������n���"��L�k�9l�Sx���.&��R&�\����"A�Ni��w�b�!1N��EF�W��]*qx���z�{>댙¯\�h�������=�Lk�R*И�.qd�x�R��lek[�Z:ϫ W�_[!��>�ppu�݉���l¢�����2[�������Yۨx�����+����z����ۗ�9�N��o���K؄��D�r�>��K�Ù2�R� �I��S �޲y<:�|)���n,�O/	�+�;�b����eG�10����/���z�3��M1:H��m��7�S�m��N�:+|I��X�&h8����\�<Y���X7�}X��ī�X�CG�}�G�����R��h�=��W��W#-ϸV�U4�⽿<��aZ2�X��F�-S��
�[%�3݋���TXA�s��Sȼ�����G�5B�m�%���v�0~�Fr���=�����/`��)��/�b+��.�1Q�ttߓ�%��aO(gx�tP������ݻ%w�����&߾���"�y�%�l[چ/��\�b�`���1hW�g�+�9v������륋u#��z�>������;_�꽨cC��A��_�gN�`��ގ��mb�dĩ;�	p
:*�L1�s��/MG�Ni�.X�B�V"�KG�ޗo�.�5u�y`W=$�uk�t��+���F�M���yW�<&b�O��~��ck��걵'SN2�v��w��#xXq;Hz�%�J��W	����:L������W� 5��R�-^�
u��պ|�?Lg�v��<C�ʇ�ם1�b�D�-�i�6r���v�`|�F퇒���û�F�0K�`��}(1+�b�BQ0���!�����A`�\��G�sw�#v������{�}@�ֻ�R�E���֛[�W`Q85�6ܹN�nm�眵�p�4��,o[՚�2]��v��ѽTo�gL���' �v4���[��5����F��t��O��2ہMM�۳���96�pXǣ_P��z�)U�;�s=���=���G'o���v����[�A^_��]�Wء)?����N+W��k��eN@�0p(l��t^qIWp�Ȕ`�=Z�ݗ8C�����,,p���(��R����V^ڻJ�`�̓�)�����V��Y��꯭2�zV���r��\���5±Z �W��u���7n�Ƚ�zm��,�}~�Нj�G��V���`���P�:Y5��_��!�(=��9����r�58#E��))�gdB��Su#ƑƄ?�-�S��4ϼl�@���G�z��)S׳�������_u�+�*9[�2<��S�%=(���{�����NѨ-����dך����7��[�K�;ˏR�q���|:��B�F3[�IA��!
��5]�.�Ŧ��K�W����C��g�֨�Y|О��\:˫����=x8=e�*X�I��������~�u��.Z���71veT>/W��1�20�_8l��U�C7�1Ӯ�x6����דu�V`�g!]��:���R�v_c�bJ�b�׆�*a<l}�^�X��&�9uWp�j����C��wV���5����=Gcw1�\�`�4I���2�ȏ��O�������l���2���OXd쬔ڔDy�m�}���0J��A�mv�ƌ��S]g��;-s�M�3('g��P
Kwu�W.���G��;���/�\���FQb�׌�M�
!�V�z����*T;U�Q����i:��z8�iT�:�hE��2&a�Qأ\dm5ǁ�a��.�{��QL߮V�U7-�ٓ;�q]�6Y�G�$�>#|��CYr."���?�Q���Y~ �n��ٴ�:�����
~�m�˚'���<��&�i�N�b�J`�"@י�������u+nFfwRC4�������g�G�|nݳ�X��	��*�����is�e�U�N����N�ֽd���#�>�1@���σ�|%x�J�Ą0�g��₽�p��]V�A��鳍��I�ie8}�%����,��z ���ztB�Zp��XW�e�� �^���D�D�m;�[�MN����qJ��l1���H��ARr�x�A����re�*��"Me��5�� 7���h��5��Fl)V���u��T'$`�p���M�����];ٛ�k���ō���8����A	�WLE�JΛ�Pzb�ڨ#��I�j�./$d]��~�cۢ�8�r_f6���2�lx8ѝnh�c�=���S��!G$����Y���I���(cwHݏ�p�Ρ�[%K�j/�Mˮ�^�H��G��P�1TH�&p�&���Z`�Y��:�t�+�ʕ� ���6_f!z)���v^!K�%��Ѷ��گJ�(ht�Wr�I�Y��ZI��/�c]4�B�i򬢆m�/��S�U��t&z:Yu�T����p�� jSx��c{%��jF/��p_G0G�.���4�}�vV������u��4	�6�4f�l22�����N�Z��ҧ�<�!���^m;w��/�:��Ĝ�:���^����m\���Y2E˗4�nk�oszʦ�n��Uى+؆�"ܾ��F�	�	�m�=kшzfr��N�i9�+�+��9���-r&��"�M�;as���Y��~ߨ;��Ij�f�i��s�<覺�����K��n�r���RB:�	dš�	Sѫ�
:�U�.��1Yd�	�{����(����
�=gVCx�-�,�D�Vc�Ը�+{�$w���]�&��r5}�5W P�����mrPf��#C@΂��	���l�b��z�����t�\��t�%=]ʞ��ɗb��;+MCt���N��Gz��ڸ�tz0�/C8�ަ6cL���kZ�O��u�U5u��sd��-R�E�oref�@�O��&���}��7B�
�bǡ;䷖ڽ䬕�˓�R�י��* �Uԩ��Tf�B��On��!��m����U.Fuݶ�_0�������q��T�OIk��I����1Oe!OM��*�I�o-^h�B�,�v�h6�;D�Z��OT��QKh��ɐV����ۍ,)��a֠�n��}R�G�cP����c��Z�G2R�3ZNV#��Mm8��ɥ�D��
��9E��*�.��g����-��jruh
��"�4�q��΀y�2�+7�i��[�G�M�	��b7z�G5��i�D��]W�Hv������J�C�:��t�e�E�/�7���TW%��
�ӗ.���K>v�1�ì���Mѽ�a��)=��^Ts����b�9[�z��ט�cA�N�l��5��&��s8����#�êo�2Pʡ�mԳ�nor���72�['��5dҦ�gh�bP�=ӏ��C+J���;��ɮ�Ա��F���_<^gYN>�Rg��<�am��u`�NXR�u��ϩm�O�a����S[&V�3�&V��z���{<1���3-��l<D�+P����ǈ�T.1�k0G��׎X���K_�����&N�Ug��GP����T��a켼��w)6�����15n!�=u���ogf��!�ź�����Μxe-���ɢWw���k��!�xu1�;�V��� Ua�ЧN��R��e�^)�zdY���N���bIB���ұ��̀#�@ ��uB�r�X��2
(�#�m .��4��-)Y�c�F��b�
р����-`��((�
*TDQb0X�Z��X�q,Y�+iLaU�����u`iQd1��eh����*���̢��@Qk+*���$uf�1!XWFDDH���R�,,"*�@R�"�Ƣ��Q+ �TA@kAeE��Trɤ�b��T*6�V��T\˒"
,X�I���DRi����aP�`(,R,��b�B�E"�X��Q`�VLeEm��҈�ċ
�X�H�"�U�r�:�ER"�b�r�Ȥ���5����,K�Qv�����9�[BU9�) F�U�TҵRE%�K�>��s�c��R=A�6�7�� �A���������Ĳ��-s�������b\o�7��W]��܀c"�O�_L�.�I1���P�ΐ���W��B�F��/��}��'i���τ��Hq�7Kʰ:�$����D���hX�U|�S�����ʆ@�+����f�2�k��7�u��C:aW`#G[����fa;��7��dȱ���s{�Sۮ^_g���/0�=��4gnQ'Wa@C-��x�Xx���������r��;{����QƂ�p5_��!�����t��<#c��s�e�.>XsU�^�	m�|�-z�f.�]�1����B�4T�~]GO��aDwM3 �o�U�%1U�k}r�c����c�l'Խ��>��؃���e�����ǚ�_{aJީ
y�K�<�a�;o��ݻ����b3�k�V)�'�~��h�ꯗ�{�Mk��fش �%��R���x����5�y�<�zWY��m�<"�%pSk�Я=�gP�Sԫ�vw���vޖ`�%���:�U������s2��S�f�cDf%4�h�\,*|(B�L�3m��>��Z}f!{��ٱ�7�Xg`Q8n�21r�� �������h���t��T�S���8Um�W�򵔸Q���e�5+��W{R�����z/
��N@�J3_�k�e�_Y(���������Lr��M=��:~�8v����,���:Dו�-�8N) ��19�ˉ�<2w��,؏�u�w��"���햕�z�E����nn=�[�{>�|jD:{,�F��̿#��}-Q��b�m	�f�����c��Ҫ�9��fѮ��Ϟl���w�-�WI�H�v8�X�,*)�Y�x��ђ�����k��&}Y�弫��S�଩%Xn�T�S֭fh�-\�g�W#.�
�p�i�{~ys$�B�i~�,b²j�YQ}�M�o�Go-��=�A�S�m��^��G�5B�h`��������0I�yū�	��Pm)K� �NN1��f�>�C�aנt�./
D�z�V�Y�CN���׈
�ّy���\
:�ˠ��h�>V�n���_�޹�R��LWT�i˛�
����$Pg�e��˷Z'�X�e.Wg	��v�W�:XrpK*�,�L�����/���mbHw�j�׺���pt^ne�C��0�\�����9���O��ߍ��H�F�3�|��;%X�-���w��MbRk�@6��T��u#��f���U�L�����V�R�Z��k�No������i��v�󫩝XT.�N�h`ce�t�N�NU�[�ۉ��yCWb�jw1��TSZKw�pS�o}�DG�c*�ǔ��n����3Ǯ;��&5�
hb�qC~��.�)q��W�7rBJ'*���j�V�F���f�#C�TǮ$��Q�������:Tziײ�������ޫ��=V���Ve���c����P�R� C�5��[���R�Ov�ݘ�O�1��<�.��/�>(�.êSj���B��q�q1r�D���Ȇ��0��[,��;�*��;�Io-V�������:#mLB�BRgCAֹ�|#�l��b�v�A�RC2DT�w@\���Fi�X~t&�\=�b�w:�/���H}q�XT���)OX{�~q5���Rs/X�t�o�O�z{������������x���9��"��gɇ�����AM$�~��0�1R�r� T�=a�L�y����*}�6�d�+��3N�Rm4��+��Y>eCg��D�Ʋh��������jݺ�|ߞ����Y�Y��Y6�=�I�
�2bs����N��S�<;a�=IXu7?k�L@�)s��O����So'��6��+�8wY- �P�s�9偎${�I2�;�c��T���BR�3��|'+�?{�C�	�͏X�{l~�i��=köO�H/�Ϭ��@�T�ϼ��OYY16}��(i%Cԕ9�d*~q�d�/�a�??3�����I_Y�{������֧��ӆ�6���G� ɏ@�,G��d��I��AH��q���AO�+���'��<��<g�bM��󤇶�Χ�6��+�}���'��s��/wI�*�a'w�R�_����Ե���?r���K�[�"9.�'*��Pl�4a�A�һPR��4���c&<\Elܺt0>�O�΍)|�S#�
��+T\�/k�J�3�*�jͨn�k�͕,�N�7p�����Vԣ��*Rc�zwaM�*�Lo�g�ャ�E]�^��[��/�ٮ`�7���  1���'z�o�� ,�,�?/�LPO̩��d��n�@�;�|ʆ$�_�9�4��*0㜞wD4�Y�����)>C��N��1P7�;�AOS�:x}����^����߷L�ӻ��Z��֯�!y���`i�Ru4��y��i���*p�0��1��P����c%d�ϲi&������|ʓ�<�n{�i�Vw�i��p������z��l|_+���'�]��f����8��t��#�AB������6}�4��l�e��{��������=xͤ;i1�q�A`x{���%a�
��X|� u*x�{a�O�YI���}Ν��\��}��R��'�P����G��!���C�~@��2J�_Y��0+'�d4}�� ~d���}��57̮�yz��h�`��2���=���W��ж��4]g.T�gގ#����=�P��x��̩�C>eNn����q
�_7a�?�a��w%Ed�.��Xi��3s����CԚ���Chu%C�'����}sJg^;����?��B�9H)��&'�<LT���T��'�]0>jA}�I�N����\$�i���M$>�N�����L`|���B�g�������B ���#k�e�#��`폷7������'��6��������%g����i��s�0��c�&��i:�Y=evf�wH(l��	��q'>���'r��R
|���P�����1{���_ݻ;yU�OJ�]� �⾡�*#�>qĬ<aٽ�R|ʁ�T�'���>ea���<���|����'���K��ĝq��Os$S�&����'̝nP8S"<D|=�L�=|��m9�9��-Qݜ������k'�&$�����m�4���T�!�x�N}�'Z���޹���'̬�3�<v�!�1��x{����Rq
���&�+�0��U��8��-�ߒI~�ۊ��~���ӌ6¼q;�1�9���ɈT����'�2���SP��[ڠb~a��C�}�uH)��8wy8�Z�ٞf�2i1��T�4G�C�7F
Cr�����^�3{7�o�}3n4FS�sT=z�J����$��-�A�Y�P� غh>̎�~J�V*azeXڃ�V!k��9ԯ����Yܐ9�����iv`'t���e2��)��ъ~�{�V$���� �ف�pX���G��B��=	Rƕ��C����{�H}���ӹ�Y"ŝjE�;Cl�O�T�����+*Oɨ{��M T4����]��
�f)'���;ϴM VOS�Lm���`���~ihzJ��g�[=�>G��ܽ�$�X��T��'}�z�H)�N{��O�f$?Zr}d�<J��P�����;f�<e@�_{��c2i����gۡ�J���Bǽ������w/��uF����9F��Z���"�3��i�J�Y��2m��M�~nRxZ
���&��Z�AAH��N?'
z�Ԛ~Iǩ�Nv��D<g���3���M�ي��=�#ыs(���.7𥗽���矿g�t+�8��c&�k�M�={��!|;��6�_�g>�tz�E"�g���a�
��OL���Ԝ��`T?$�|~�!�}�*
p��3�<g�X��|�S�=LT�ߟ=/�q���|����ƔqWھ����"D}�����d���4�T6���p�w��䞦���d<f�[�O�5����|ϜdX��vs$��I�8�?w$�'̩�{���P��s���^?s���e�z����$F�!���c�:wXE:�Rjg��6��X?k4���?X�O&��i'����Nr�$���S��i�bCӾ�{����T�����������m3������Y��#ޡ�"#pĈC�z%��/F��?e����Ld�?8�3����
E%~w��X�)�t��_�����r���&��J�����j� ����Rm�i ��w_��ﾉ𫟱�J�m��"���B#�1�D�!�6y�M�>jCg<ցgYY:�Ρ�1?!�1��i�+��I���%@��~���(�Y�C��?0�C����'̨z�=�m����Q5rX���z��e��""�x��}>���7HT9�z�bg��rj�N�T������~a��0>k&�1�*J��w&�j~I��nIYR�k�`Vi�I�<�iw�_ڑ�����q���M��!�����:pY:ʓ�+��y����O̬�=��.��C�ÿ�6������] �Xx�������t��Y>وk�&v���i'm�?[�$�_���	��u����;�0:W��̦���Ֆ����Į��j��i�xU�oJ��yqou���Q)�׫ {ф���jn��s�M���V{�oL�L�w�4髨�9to_�t��Fդ�WT���`�������z=��n���i�i}�2}�= E��~�jO\f2f���CiP|���h%gܯ�+'̬7<��m1�a��>{M2c3(u%��M2z��g�I��M~�Vi�"�d�����76~
W�T��4#��c��d�޺!�J�&�w���H(,��ɧq�4��a�P+�&�SI�� �t�!�|�g5���-����.��<f����C�i��YI�\׿j�o/����q��eu=mS�E��� :�+�0���}H���
��{�M�|ʇSg����L
�Xp�3Hc������H��3�P��T�Ok|�*C�Ho<֍�m�����'_�	���aO,?G��a�S��Ak�5~Ì��R���'Y�;��͝�\dX��P���'��߰�x�&2u�����C���C�i1��q��f������"�쉝1_UocZ����=D N��!�m�ܡ��&!�)3�'2���PRa�u�;�bAMl��u�O�f0��Ձ֡�T��c��WP��q�d�Vj~�B���z��n{��n>�g3����iNo|���y�0��3hbJ��=q��p�h)7|Ï��E>a�,�M>3�N{���RT��I���P]��'��?2�+�&ަ�C�C�R��>׼���u����/��X�E=�ar��̬�{5��<jz��c�y�����Y��q!��'�}ާ�6¢�O.2z�����ٴ�xʇ=��ߘ̬P���큿?_/���щ�&���Z�¦�]�X�<���{�w��4��T�_����['��d�b~a�L���膟̨q+8��YĂ��x{g��OYP7��}�&�P�Rc���E�4~�4�dc�G���ӕ0ግ�}�e��)ٟ�$CxɌ�N�t��{����|���8����a6��aSG�}��L
� p�ђ~ev��)���!��3����Ă���|���5�bA���2c��8�g{���a���No[�}�~���fXj'O��X�����
��+�����x��1��i��>�O9�P�J�0ϾͳL�"��A~f��)�~��I��bzÒ�Ƌ��"�
W�eX���1���� � YY2�-��N���x{�,��:E��OH��������r��Kņmc��ujp9׎��CW��W�֝�K L&cY�,��oU��s=KN-��ܜ��٣��!�O�-!ئ&bnb���{�]Qz����ĿE�Mۉ?%H�I�����N�W�y�p�C��w��������}d�Tu�&緬�֧�4�>�d�+Or��T*$�y�X�� @��� nd��>t�f��"���+��<���2zʜ���<������D�a�;d����g�q���� ��6s�Sj����'��� s����K���E�� G	��tq,��'=�|�I���'�T���Y=eC�a�ٛ`~k"��<��iN����a�*q�&2l�jm&��)�&8��+���h��a�0�ͽ`T�&��'���菥5=��xfME�=�K�*:�z�>����Wi�|�]Y?e����'Y?8������;��f��2��X5&��h.�VO���(*q���sT�3L�3ܡ��I���&�N�L�nU�n}=��P���PXvj�OϬ�,�}ɬL���p�������&�>��oA���&>&���1:�_��/i�s�0Ѕf35�<�F����*�����0������ݟ��+mOPuC8���e�&Шu%x}d��aQG�XLd���S�Y� c'���͡�<���S�y�Rm�m���rAH��4�9�H>{�[�!.���L�˂����XT�Hn���2M&&0ۤ�3���n���eH/�'SL�eC��G,�eC�M���ZȦ���+R,�eM��CI��LC�ܝf�~&�9����g��c��}t����=IXm=>�4x�PR)���8�3��?3�l4�Y]2k�}�AB�&jwP:� �v�>�N嘓A�J��|��il��{��� �G����W�k��g>�]�+Q��A��'N�+4��T�<C�g>ed����w��=I�6���6�tͲTq�'_�Y=�0�I\f&��$�wH(i���I�O����
@>�E�'vL���-������w˽�%@�������Hj�l��Q�1a���C�Ag��;�%f�jx�;�!�N��s=���)6�C��H}q�XT�h�Y8��*�����B����pw�o��U�7�`Pʋ�R�9)z!<6f��E%ZU�7G���w$?��+��p>�}7e%�v�4��Px�Bx�����{�ii�^�:��w_u��ś��]�q���C+fgL���k���H��W6��l7��qv+f��.�����
O�~�{�c�OZx������%C�s�VE"ϓ�;���R
i&�}��z��Z����z�n��w�J��PSy�l�e`o�f����i��W�����'̨~��*�VI
���:��=��{�s>��'����'�T��LNO�<f�|��O��Cĕ�S�~����PR:�u
�������y&�?2�C�e�- �Pѿ���H.����<0{]����=)+��G��z��G��>��'�l���6���?w4��PX��'Ɉ/��Y�4�ԩ�?'�}�N2z�ɉ��s����RT��2?8ͲTg��i'��c?S;~��L抵�z����Ij~�" ��z{ۇ��ܤj~�:�i�O�Ĝ�P��Ԝv�É>@��6�6���R`����I��󤇶�Χ�Ͳ|��Ʀ���Cl�2��w�.��ȫ�t���|��}��ǰD�w5��i�=a��|���'YS�Y�|qnw0��I̿2s�i�T>a�9�tCH)k����)>C��'Xz���r�S����sU\tq��p+8�����P%d�*M�u����~M2z�k���m��*s�Û���C���,ƤY=��4�HT��O�Y>eI�e6y��>IXs�=t��*
�	Z7���g�ݻ�C��L|���N���:��oϲGt���O�Cy`|����H)?['�f<�YI�'�!�����q!�I�}ާ���*�q�P_XT�����O���[�x�J�>U�3�럽{�<G���ry�$�u&���~q�d��v�E'_��Ss��4��RW��0�c'�� �;��I����q���R/�=9�W�Ă�2pﹷԞ;M$;o���=�B�*��8�\����fm}�"��LC����!堳g�ɦN��7|ʟ����*rnì�t�B��ɻ i���3�*(�Y:ˮ��V8�����>f��&�����Chu%j��kkk%	�W��G�ɕ�Y�_PAH�=�!Y������&�z��72�uH)�z×y��H.�{�Hm+'YP�\$�i���M$>�N�ut�j�5<��V,��R����d��dB� ��&:����kf�U��kWQ(�^&n6�we�호��M~��`qh���{����Z%M�pI������R��p`mn���;�x0v��[�>��[Λݘyּ!�H5�l{�wH�0���B�!]n��G�ѹ[{����h�m
�x���d�'YRz��������J�ߩ�+��AONy����z��bu�z����� ���N]�:�NO�b
N�'r��>d����p�^}����f�����ߺ�m!�ߵ����TM��:��/�9��Ru�ĩ�y�Oq��V;��(m%C�<?SL��f�.�p1"��3�s$S�&�k+4�2~����M�Q#I�e�s߳QDT��&�ǽ�1"��O���
~Cg��Ӊ6��`s;��C���wR-Hyh;�N3L�2�o9����6�2|�r��{��B����&�+���8�<����v�<q�i�߿p[���QH�c�cXW�3�ܑf!Ԝ��s�M!RT>Mw�<y��ACf*3�R��(O�<LT3�G)6�O�'��X�3NB���N�j��N�ꏾ��8�>?�~M0��~f��&��M!ܤ����$X��H��i���6�<;a�Jʓ�k߰��i�����*�O���1H��=f>��;�""��@��e*�)�9��d|�b[߻���^�f~��,�!��LAI��=�Y4�Sl���6���֜���Hx�����H%A}N�L�2�u.����d�+7<���؆#�DX.�b�E�
����>�lusZ��{�m?8�0� �P�?3��2)P+5�2m��M�u�I�h(z��̞������y�p�~N$�<>���N=M2u��A�?'۶=���I1T�tg����5i.��s'{��1����;���~C�c&�5�Sl��I�ü�x�h��p/�x�E"�_y���0��$��'��u'�y~��T5?}���9hc>C�~Ձ���3�k��N���Z��Բv�n��#�D=D�!و�F �'u��C0<k'�&�ʆҲz�k����'��������Ó���6���/�2,Y�R>�$��I�8�?w$�'̩3���2�ߏ/w}��]��e�fSh�w�4��=q>@�?Y���c�;��u��g��6��X���B�I���'������>��YĂ�0���<x�N3����5���|y<�����&��~�9���eBwG�:���$4$��Yh|:��۹�ʞ�[Ŵ-�Ҳj,���/>95L��xa��/F���;�5`�VZ)g1I�Ί_*Z�NH��1���|�ާ���5q��9?�P�F���[D��X"���ވ�{�;8)�ڜ�����*���i���>�OY��2|��d����RVn{z�L����p��AH�Y�bȧ��~�A~f��'��L��hu%O��=���HT��>Pf���"j�J�~��;;�t�n�I:~���I8�M!紝� �x���M�>jCg<ցgYY:�����~C�cZ|����Ri7;�Щ*8�}�a�QH�]����¾8���ώ��ϻ�ߚ��~ֽ�~��ߺ2zʆ�s�u|`T>I^�ܞ����
����,�8�ud�1>@��'?o�m �����<`|�n�������w&����Ed|g�#�G��|2��Y��Y��ȋ΅f��)1�gw��E�<j��,�2��
�\�U񓌝eg���T���s��6����Ɏ �Xx������?3N��'&�P����#呱�_u,w3�l�3����s�wĂ���N��B�=�W�n~Z��(+����e�x�?����2���u&:��㹾���ﻂ��%gxg�܁_N�3&�5b�s�D��B�h�=�]|{ð�TԎT�U*kiq�V <��9�38rj��l��<-:�%p2c�te7������{�������g׬}P�cyĪ�;9�P�6��2��edrV��^zֲ�)+�$��ϝσ���7����ŏ�,���t��+�0\2	��,YͰ]���`�+�.��w\�=A�8"���T�}�e<��s�~ͧf�������+M��G�O��eW��2��.�ҷJ�ׯ�A����@�,���h����'V����8T�Pezҭv��+z�	��RG�Cu�v�a��:v0hu�6�̢+r�r\�e!|��J�N^,	���:��c(�Z�LD�*U����J0��tgj�Ӆ՗�"��eiޢAټ���1G��7ڶ�kg;Z��C��0{6» JMn�أ�JKv��Q�z����۸��$�ռ��#��fP��]�+. �.�u��>���g�^���ԛ�m�W%O��e��toh��nL�����e7��=�wHU{�/��"�{��w�ʔ8R�ۦ��=:�D���b^wu�6�"��s��ٰuL�ػt��	������E�|2R��:���;��T�=ەaXVt�O��<(�Y�����6n�S����Kᕃ!�O�f���BaT�w�0-j�<��w�t����u+h"d̜Ƿ�����u�����m�XTk!�*8̷�f�����B�ڥW�)y�A�zr�[G
NV�����k�ĸ )���.]/)]u��[��{��H�wfĝo�]ջ&�Gnv�%�	rv���S*m��KG>��֨�ͣ����&��{Z��Mb�+_ל�����$�ouo�VJ��5�_cJ`�K��z;"�m��-��G�sr��?vu_gS��$�\`�|2^��G{�5X�u�/���jV�Еk3�K	;o��)6��T9�x��lP�]O�V�`{��ᇊڕ���\u$K���f�I*Q뷤=��]��<����gC�x��t��/!�C�\h(l^4��p�W�6Y�q1O��U�p0������Zm�wt�j.�J맕��т�t��7��]|F���d7ڂ��NAP7b��U�h��8W5L�׳���N �l�AT�{k[�_fE�a�ʬt�ņ����6��*�A�E�#�����em�0*R]Y�h�N���]�˺Ǯ�*���X�*��{������w�k� BN��n_eIa��η�uk�m_YՁ2N�|��ȹ����4 ����휹p�*��bgWN���Wx{�p�gq�éOmJ��nrpLƅH�N���B��y�t�J6*GnaMM�DZ}�\ ed]R`���Y��5�k�����y����<K&[/��*$z�I��nK��Z���ٴ�KQ�].��k�?�d+����U���4�6�:�6�:�jj�r��ӆl兑��ӣ�Ķ-6��A�ѽ2���w�R{����5��wU㖬[ؖ]F�Ď7Λv���_Xqh�IM���Vܑ�;��>:r����j�*|w�"���Me>�]M.2�L�؍���4�;�X7��y�H�~�m(ݳ5ϑ�e ��۔n��g'e����o�aMq�[2N�뻢��b�@��q;)�ƀ�nU��{QN�h4sz�(�j͝��Ē�w)7J�$�� z�F'�Eq��UUWv��
��(�E4�U����b�b�1Db��TPX��V�E�",TI��b�kj��Uf%c�+Mۦ��X�*Aa`��U� �J1H�6т�Ab�4[J�,��!�T5e-�,Y���bEPPQQTA�*%�UDQV
�EY�wI�ճ��)�n���U(��n�,�(#�fY�b�e �Qf[��h��E���rન�,b(��8�%DQTݢ�;�LlV2:�PAE�v��(c�QR8��Q�Kh��0*(�����验v� �¥�Xh��  �  @��;��zFq�V�\`tshS}$����m�����*Bh�k�h�wR���]}4[� [����U�ٟ���V�4�s���޷Ƥ^�'eVÎ��[�!��P��Ѕj��z������������m$�^�G�j\s���1������h�}�l�[۶��X<L�5|��1A*�Dt��	t���q�_��|���;=��%%r2���+M�T�;��O���&�b������Ň=ܷ�Y�%�9C�7ܦ8!|�8ߚ�E��)T�_�B�mØ�v�mR�]�SW��Y��_.=��Ud�LS�PW���Gx�~[0Ƴ���;bY� !R�@�Q�ꎙ{'6��G�C����tP��̺5���[����c�	���^E�1��ɷ9=�ל���P@��B�T@>:,���|��n�J�#���2�.�p�}5�L1CO�%�ɫ���X�^�AE��G�	�t�u/���9�y������`�Q�#2��n"��|P6-U�ν����ܯ�/��x�B�|� b�ƞ��9co>l\n�XϜ����Rn�V,jqmcFЩb���ũTǮ$��U*ӣ���t��z�s���̭wn���&��a���ΊƄ5#2��[b4�M��בyЖ�Ucn�c$Ƌ�U�[��r���4,N������upwܠ��75QN�i��܎�&�J8w ���\���8Gn>�?��^�Ļ��g�T�>6��ͅaz��  b�����彴�`Տ��-;����<�'U��C�"�]Z{��bw=C7|gt�f�#�\�>~�q�]b��t	�n��B�(�:���J;`ٺ���M�*1��H��Q"t^]?O�y-�r\b��a�����*�8�=��d�V�n���f��ݲ��R���
�~��(�hu�����\ə����9-����=���J
�l;/ �qŦ�k����@c7f��*���A��Ƹ#=VN��<�L�n����8�ʫ�4F��3�%f��l�#���C�ޒ�X�����Xg �㗼;{sB	�J���_oU
��E�v�b��������tF
�4Ђ���V[5kz0RJ���yS�i�d�<U(��u��T�7�b��,C�wH��.��mG/�n����M�2%����6Ny�Ur��|���[�	�2�������2Ԯ����sgPt���C[=�b�*���)�C�����>������0��<��G�P{S���,�Nt���g]��&��R�{�+�R�҄��g�سz��\�\X�XKg��t�gD��.��q�QP�����u�<��+���r�D���bn�s��3[{|�W[���	c>��ݗ*E�ߣ��]�#���=�,j(}�h.�Ά��<_ܕh�p���~�*S��n�p6�(� �_x����;���ÂՒ·;�ţzH����r�h9��Q��������<�ѹ��ٶꘅ�V�ZE���u�.&gF�O�e�T��r��hVf����I�K��ү��IX��硊�(����sA�����L9�th�����d�����g^�'�F�{V]���9k��w���i)X�JB�B�V�0�IUD�Ui�Y��]��jD�=���C�tVF߅�+�8J��C�ذ�+2tC�TR��'jAi�ƅ�����T����%jj��(�������Ԏ�Kǯ/���k֍�r��S��Χ�)��N��=_FO1%�Z��`�[�B���a�o8���,�w[��u��Ӽ~�a��t9��>k�z���Ŷx[�(��#�qD�ʬ�+/�V�$E���Eb�'�����Ud|�訌��w/0�����&4��Y{e{��tj�u(5/,0-E�U�ʽb��;V��A�9׶/.�ʰ�ZՈ_�J��x%�9�[��c�J[V}\GA>�%�i@v���m�و,s��Z�a������RN��-ެ��gU�⠕>�ˆ��v�c��3�UG�������Ah���f�=Zi�V�3��N����j�QT�y�^��N����i�x�^),<�=f�%W��ux��oi���O,gz�s��2�u�gR֯s._��ū����@1��Β�j�v�W��KO�+L�Y�d3�5�1�ȯ eurs��W�UҰ�cx��0��F��%���:I]�4Nye�խ~�=+����d{U�>�p�ǚ����������6<��®Ó���
1e�Ií릫q�|K~b}�)�����1�5����|�x��N*l,���%�+٩�{�����0Ϫ�ђ���쑱��Q�4x�f����b�4g��=�^�[�W��W[��MbHq�'I��^�p�1��\����C�t�'٧K�*8�����m�����b����/n�/��+��2q&<,��WU��7~i��yH�Cc�FS��Ǟ:o6���G�Y�����(�r���My2kdcg'��|i�#qx�x��;�]�U3�S7A:��ջn��}�,�}�y.�Z�g���g�^Σ�;h�a�-�f�63d�q�o`��!�ݨ��Ώ��)����4�گH��;G)��V��Dw�}`�Ĝ�L���j��%�O8>9H�u���\1��U�ڲ�o;y=]��6J�����C�v6�gkl��:6O�H�")Aa��H:�!�#&���s�4!s=0�̚����jl�u{��|��ꚺ��E�zT"����괡�V��)�h�Ue׉�z��ӈ�� }���;��a���bEz,�.�1�Y15Α4���ֳi@�rne�&�{��d�棡a��T�7���^?�-�S��4T����Dt�Nhu�!*�����Z�hޡ�����7/i��w����	�V�B��1��c��n���V��b疚�;S�-��=Q>�5��5S>U<��bUsZ �v�l���q	Xlx�֢fdRU�ѯ5�^-��q��Z)^77�c�������'��ϸH�S<�_qg�JK�f�V��W�> �}[�V��\}ZƖk����W�=3ʊg��y�S�WUb7r�h}�n�z����R:��5�b�9J�ä���}�����!������в����M�/�ßb�jc�Y�Hp�%����������^Tp����f�T=�K�r����{b�j)��6-w�^���w��Ǭ��2����0Au��%sgU
�}�m�(̙o�� j���:�������F����]�ū��ed���|L}U�ᣘYPuǯ�Ү�c4�Y��aX������_}^����Zڋ|�LQB���a��sl3b�׶�Hۍ�]>�n�͍��غy!S|:L!!�|[�>�,/R�)�X����'����~b�D	�Uy��3ff�kn&�Zcܓ˜j��3��y����x�BĈ�C�S�����K�ѯ;���W�7�_�kMW�T�P&�X1�4Xȓ���4�*���A�C�4RrG�t��\]`�U)�lv'ǭ���}�wZ%��0�wʼ��ʇÔ1P�k�"<ײ��>�<�r�[.��,�\;=�C&������`���"L\�(�$��Ǫp��9�a<�pH�)��궅+ח��|��.�O�|!�q��}��p缪Tb���u�t��\��5��p":�֒u���(E⯔H���_����,����	q��?=,(�:���v����5ĝ|z*=Jg�__b�u��X}A�ݗ@Ņu2(pW��N��>��]'�']U��1�6�X�md���{�z}hup�uQ���:���^�Y���9W^:l�� �����ESk�^�J۠CU�l]��vl��*k�rv�)n��u�h�wg��AMs���d��b�-�z���|d�wL��T��.�����u�!Ɋa��2�ܨ�f����Ԏ���]G��⁐oW����7�'q�K�zW��0�n�Ma�kܪ�Y�2L1IK�嗠�tFxF.��Էm�k]���C0W�+�W�S�q�p��X�P7������_
,t��lX���{��$��N1�� ��=I�����U��ّ�Qr��~�s��p��݇��U�'�-OM�y�A���Pu��G�kg��C*���)�C�������+P0�b���.���Y�=���w��s�P��C��rU�ɕ�v~�>�]vjp��={8�[UkmL���t[:U�dY��5&4N����(G+��&|�\ύY�R+������mTά�cőV���2(s�l�.>����< B嗩Vf^���W���Թ*���B�N�~������;��:E|���2����p���SߟK:��&�f�ir2h?�'�.�Ne��8f��Wxi�^������a�.E}Y崩�Lb���Z��|�E>�*D�V����Y|,+q����C��(A^$.����Wb�6�6Qt8,��0S��b���c�lRڴ���eܮ�-�{�y�K;�Ԕ�x��,.��e��^�;2�CM�~<���L�Yr�np�y(&���Cd�4����I����nWp��+䳞���)Ӱ�T;�[�d�6��G������H_��I�A�?F��Ϛ8L<�&�l�����b��r��z�dF���:��g+����{`>6g޶R`g0�K���2y�~DV�o��=�<c���WJOU���[����܈@q�#�3�>�5��ĝ��!�����D�Ԋ/���q�	eΗ~�я�������6&G��KC��T=�W$+��7�H���9v�]��:���R{xŽ���� p�1��}5P��~6+*�N��Y�Ҳ��]<��+�G�缟{��&'�T�}�ݩU��#F1=f�Up�~tv�5i
��n_��~��!##�����';2��8�+ߡ��sRF�Oy �EΟb�z�T���t&��W/U�+ROz��=�^�=�]r���.����>)T��!㞗1��]�,Zp*5+Fa��
�j5$��"�U��jP�s��xhbc晿7^
��u��2�b&���|#0����Nt��yn}9c���r��a�*��9�^[��0�m�Hb%Oes�uhj�P�j��d�P�t���=��n�a��T����aR����W��m�/9��I���x[=w�ԗ�ϫu��6�˪o^����k�y�ǡ�a�i�:VH���d�l�1���"�/{�F ǂ�:��v�^A����l�
VS�Q�& �ܵ�{ѵd�\�;c����k�5I�Y�4���C^<~G�C��U�3*�0^�����w�z�T������!���S��a�����ԅo��뉟f��r�Ś�B�wRK.6�׭GL]�����j���K<,���g���fe+6Hab���;��W�˟]^��O��uB����(:�5��h�P��Պ|����8����D�}�,B�ZSZ���"���F�O��)�C+���FqI�7�e�zxӋײ��X�̒A�8���Wo��]��:C,\`�.z[�%��$͊�� *B���4�}{|�T-a��s)W�oӂ�	����,����H��,X[��E�չ��t�u]�� p�ӑ-���԰d�6D�({-|�c�g֕�L�{��ML;�9n��Lپu��5�-�
ܡ�Ǧ�r4N�%�g�:4�׭�c�Vphb� x{�d���{s����:�¢�!O�l�s��|}l�顾�S�źʁַrE���N��^0湮�"���B�]�N�Wt�;�VkB�s��:������8��}����c���]��u˹�,lE�w��H��+�����ds�B="�5�c�����w�BN��TtRx��*�'j_��n�e�|3��Y�`�w`��ޏwN��=���M��ڦ8Tj�gq�W��ߡexLsW#.��
�)�Gj��@����Ў�=�n�j+�\�0㱚D߰�u1�cza�/��jx;�4'��{]5^���ҍ�4�ʔ�o(��8ɉGn�\;���+�f���(+��~�xo��1[lN��s�>��xg;��,Ɖ�ű���ҡ�5ƀ��f���~Q<��{]n���=u�뽹S}"�ُ��vV��C�(�^LZ�f�p�����+�����C0��51�1�u��W����o��m�q�La�QMS�
��`�&�K��#��P���`WA��+�7֮{Α�2���#�d�z28k�ί���S�bDt�©�Z�Pط0\��c:�wd����!�O��>6�J�M/�U1���:�EZtG��>C�U�[���Q|�T���Yqo2�v��E�.qc|$0�̨}���D*�z]V"�S�e�=~R���o +��O9�o�߅�rY���_���`�툓��Dq�P<,Wy��m����Y<�}br��@t�:�uƳ*�;v����}�qn!�����¨�ev�!����Ԛ�߶̤W+�7^X�d�o�m��2��/���N�W�v��Lּ���T���#�v�{u���x�m��F�k�C��ͽ����[/Y`>�XѬ��W�W0�	֨(��R�94z�[hŵϨ�Co��,�h���MnZ�l4'4����[�̓Ǘ9����k�n�v��2N��Ѻ
��w�[�G�w�M�h+�R)l^��&�;cO*X	%n1Z��j[_`��س]�)q� � �^���!����
�/�f\�l:oY���rp�՗V�۫qwv�i�H""�+"�9]���Qس�2�;U��rb�rN7uy9ަ9֒�ۢU�S:k��ǲޡ�mt{f'���+_ �v�sz'��#��`��_��p����&��0���xʖ�ӾT�\(>���� a��U��%#��6��[R��dԣ��p`wf'-�>.ӽ8�j"�Џ[��z��s1M����XYHN`�;�I8�`i���]�cm:�y��b���!J���tb��39_Tn����B�f��H�p�Y�K�5��M������	�|�D5��#�u���װ�g:^�y}��w��}]ՔsF���u`q:�+-�uc8mǵ�S���!We:8s�f���D0�VxKs�nb̫�cGe�5�A�-�w���z#O�WwP�H5>)c;�Ϗ4�!�pRj�G]GSYV��(s�s�\�2�G@�m��ɢq]��)�'���Vz���B�B��oI�T�B�<��{���q..�p�}�����VJd��7W&M4�-�&�yc6���r�0܃��MJ�':ħ�u���k~�R�UZ�ѥ8������Y�1��A�e�@����%kμ`D��x�rů����4V)[�0�y��ts�pI�j�h9���u��bw�vP��b}5��5V��=/����m�D.Ū3��d��36�����ky:���;Ĳ�^u�{Z�	��K3�P<�:����!M�ܓ���<�^��[���wS��pSTY�p��|��[|.N;O���D�Mu�G�u`]���;����e#[5㒂�@<��6�����A��ӳ��y��k�^��аr�7]u��X����igc�x��1�K�7�����;�D�^�:�v}�R�wRh&[�Ԭ౺k���i�Ԝ�Ju��z:B��!�7wI�0��;��f�֚b�;��Ǽ�����`�j�@�ej�B�i��.�ƧDR���J����6�)xGd�N�1�X�YAj�.F;];_�oi;{K(ɪ�(++�a��m����p�x8um>�e��a�p:���tqn�u���Y:>���)�K��o�ٻZy�n%�=(s�+� e�V�Lå��	Ep"Aĺ��P�Y���
�Ԕ����t�g$<Eـ �� b@����\t��"��ACVQWiA�1b���6�(�mQr�ED`���� �Q7lLJ����4�U5(�j3�,]�*��ʆ���e�DƑ�
m������(��AQ�V3y���T�Ej[LeQi�b�D��Y3WZ�E��mT���E�� �F��V�i̖1����#��%�XTTkD��Z�Z��݆aA�բ0ƥI����n�����f���#�cTdb�(���+u�r�-[j�6ʪ#,b
�e�*�42�.R��PT���b*�,F*�Gn8�֬P��Z���F��f""�Z�rin�ƛ�U���m**�j:���J�V[-��-�b�lW���*R���TE�U 
1]�q��x��y
�q&!����oQmq#��r�ku�����[O.Z�G��.��:>��L����	u��$�h������������Uy���g[����,�ʴ(e���PU���]�[/*����B/��}H�8�Oedކ��k0����DN���(�/(�g�QU���CA^S=%g
�]r��p6��e������}�yJ&Qa�
����MG::}^f�,X2��NT-?=n�\�}��Y�O��b�f����-�Y(u��[:�š���m��އm�bk�T�Y�ƚ����<y��Ɯ�è�*��hE��P������E���f�����r����H�����6��劥��k�ƺ�q� ��=����2��k�g77S�;�'6�ެ�de��Q*eI5�P!YAQ�|�]��W޽<���W�)W�ϵ�!�^s��8R�;VZ�Ή�Q���	��A�z��3�<�Y'wj�J�����e�������q��N�5�30���Zoѿ���щc,!���ϻ8�+ڵ�Z.1�pt!XXz�xظF0��;VyjG�P�S�3ӝ����G7�[ۋףE���a�#nl�
��)I���I�玃�sׂ����LE�&x��0���,!Jj�+�J�I�FK|� G�S뫀�-e�[I��8�aU���`���щ�nJ\*�a䥓ON��S�U}�������y��uy��[U�-P�"ε�*:3�7�x(@���3F�V�J��gq.�jRWV�����^��]�T;�e,@��+�ș� (s/���#GY,�Xd�/3�Sٗ
��px`���Ю��'���8^@�S�m%(c�a���Y��y8����4VҀbyPH���}��FE�co����\�=���	b:p�ţ�����UQ$�q�'$N���g�T�0댚ٸ�s��l��*���ӓl�i9�K4wd�{�f�.�^��Ѭ�Ry	���P[@M��l�x����W�M��3k2e�N�.�֪Ɗ��bB�|�F�q'\���p�_҉�3�"u�\��p�$����p�p�����f���"2��C�Q�a�5��^�D��ZDW�gy�U�:�÷.�Θ$�L��z] �W����g��e�������ڭ��Ɲ��cY��4{='v��?3�u����OY��U�ź��n�zً>��L��m�&�AY�pgK1�����Z'��ɁbV��P�]��ηNA��r}��X��^3�9�(Gu�[(-T��Q+�jl������w�T6VU�*�8�y���z���!]0J��ɚ���v�5���6�4��Vm���z��WN�Uѩo���wy-<��!�>�B/OgM����HՌn@��*���7�qq�8L�X!���ܽ�í���C�<.�!p\]����l��ѪB=�Ug���պO9��L���N�m)�q)��G�W��=�5qa��~ׂ��<�����`1K�i��yF���c�qx���=H�,�Gؘ����ezظ���l ��9�ݸ���u�t�V���oQ'ŀ�C�������˿Qւ�x�z����{��hE�=�Q;ݛ�z���Į� �V'I�:U��1��\����!_�Q��3��P d���KZ�c����#�Q'����	�ı8�t�(J��o�,�����G��WJ��_5�N���۞�~5>�e�+��"�K���Qu�}ѯc$C��
���J������l��:�kZ����#���T�\|ki�C�p�@pP�N�jd��FMvq�9=0�A7��pk�m+����4�3�Ա���0��E����b5�D��Ao�h:Ad�4�-���S��)�����7^m�C��z�4RN��_A�����-�+Q�ЇZمA���w9��N���w;qj܋hS4�unV�|�[x��1#���4�������i�k�1����%Weq�C�a����S�^��D=�N��H�8��o=N��~�����@yKP�����A�|�i�R��z!v-˗i�2�$>�'4�Pv�v貁�[��/>�f!�T���6���S㓻�\�t诬�c���v"�}s3Cx��ӕg-X�.��S��1��$��Ͷ���&��^�{���rf�#�Y�E�)�͛�s����S��'5�	������u-�Žu�B�%�b7!�d���l�w�8V��w!�B�����E�p��Z�'��uK��&�v^~��O_T��M�)t�	���s7Ǣ��"��]G��s�3x�������?Weg�;��G��3�/s�ǽ���Z|�!҈��wu��K��{�U�C�11�ʇ���Y�Du�8�j���<��e'p�Ah�w�;Tw$	�8�:��)b�jbРF�5��z�-�B͋��{r�Y�yz��mWG�;.�7�X��-����S*cE��W���.K��7�V&8B�����K��yhwE�(,*��C˕*٠�mH�u�vZ�4���V{�����n�ⱦ��6hR޻�o!�!�A�ۃ�1	��.���r����b��k���b���]���R�mRYP�0�}�kQ��%�h�9��.����>u��P�ۅ��QC>�/MD��^�,T-Uc�2N�Ls��P1WSrY�ڋ��[�g�U���bS¯𺏳&?
X&����*P�ߦ��S����uF��잾�ՙd�7&W^5LVG�<G_B�J� ?8I�U��!�K�fT<a�ׄ�wA��S�t��3p���x�vgǼ�m��-J�,|���x�-�lD��A����]	=���y{��!�JGW*�X2І����^^z����.����B.0�0��Y�sVы4WA����YD�;:���aT@��v�Y��TH��^z�v|xc6�Gc��o�r5�&p�>�:�$�2�~=��_b�{��|a��gn������yѕWܔ�C"C�;��-<kE��<�h�u��x��\6��u�D.�5sf
����so�a���v����`Q��~~A�ڝT(d~"ϻX���pމ��Y� 1��v�U_H*_g;*zR6hZ8����B���o��1>X�P:<�G�V�*#�R�R����n�.�E���++�Yٻ����-d�S�Ww������2��<7VK�U��N��(�VZ(��oU%�{Q���23 R��j���]	P�vTg8F�)ɞ�vC�&ҥ�٩�/�Ld/��k��z<�9��J�kj.���P�j�*%#X/�����<r��Q\�9�B��AY�]Q�TUM�ٻ��jJ�X���nbE�{�Pt����x�a�oK�B�y�֑w�i��6=i:�݇��3V�3�c��̭#Öj��dcJ�����<]W�d�������:|�����&�ڝ���*�X�24������*�3��r���;���P�b��4��'{{�>�u˶��>��3!i�[�dU�\"�8h;K����F�Dܾu�����e�wH�>J
���.*�*� .�Wc8i�R���SW;��'����׎m�ދ]7&1�u,C�6*]p�˻CE��wU��4��O=t�Cy��d
��h?E��ܺR���%#|a�j|��B�*5��N��tV$�@��8Om�9ߴ�kB9WW�͚��%�C`b^��G��ت/����%}����p��b�6E �T��o}K-��\����l�4Pr5�A�'�y�
a��#j��O(҆�9�r��q%��/�@�&twW>V�&�
l���u'��ys΂�)��?5�cԝ�ޱvhz�5Q�׬RO7햻�g`S�^b�Mqj�cǻ0�<U%�\�L*�_�HoxP�(r�w�kS�KX�v�胷0e�����\�r�����y3R��Zͤ���Z�y7�6�C��<�da07�$��q��Ģwv�ʻ�!�Y�)ޥ�F��q�mp�}�rz2*�z���q�k�y*y���߻گ�����҃�J�_B��ޓ^�.����r�u�N{\	P�.
7�yU��c9��*��5����M��)�\��~Y��l�hdh�u~ag���}-�3�vj�u�C�6s�ڬ��Gw6'�'�N򐋈egM�(=1n��I�p�@��*���+jv�Otk#�K��Q\߫�k��Jda���c�8�[��->!����bS"�ڨ#|c<x�w�v�CM�}���*���i����^y��]�G����\l7}��������2�!���7���V=��XA���s���#U1�S�
�����`���`n���2FJ��ﻔsb�.[V �~કi��f}���x�R62��3�xz�V���<��+��^����-�hT�A�(;S#��d�x�/>7>b�n��[�i��G{p8�5�
�i�S�#;����3:���Ve�^�Iw�"�Q�WLQ��^�3Ko�[֢�h����ѽ�;�oL�Z�{��:�0Mu��IjWtT�I�,�V�����ōrP�6���-�.�"�jjLٚ����
Tq>x<���m��}F9��� S�nv�s�l�c�_b�G���h����.2q&���p��������cuS�چ�ZL=��M\r��^���^
��!NKSduJ�P��'&�@�:rw(R�
�;���z����Y�4J��ݢ˪�P�4᯹�8(b�+���SG�ߨ�h7)7��}��i�1��3��^fy隹c��`t�8�R�p<���G;���ʤ�O).���٩���y�r���y�8?�����a��|��H2���=3�`�«�o�7%����A�ㄝ664Qcaw��@��*�E�W�߶��qY�y���x�r�Q՛٩m�����sp��8Ⱥ^c2�X�x�|]�k�l�4r�U���J���T�J��q�GS625�'���J|�f��C����M'EY2M���[r��;y	Vr����{�)l��M���c�����P�PA��Y^	���e��X9�Y���K��\�"ĸʬg��v\�0�D�g/�a	�0��s�m���S�H�	+��A@��9��B0�LLD�m�WY���D(W2
�������it`���"�os�K�K'mp��{)�ɇ��$�d���`���q'X�]ʒA]�}κhQ���cio+!h��b�ʾ�d��.-��Za�ح����Q�6�Y��}���XkZ���jޖ�G�:���K�J}p�QY^�Fr�xt�U�R�w��x�.ڥ�&Q���2ڭ]۱��<�7lH!�t®��
��FY�>Ƈ�ϹM�L�c��o^�=��Tb]gb���^W�;�u��E�05BbРB��M!����b�ع9Q�'�-e*t�3uc]y��Fk��Ai�>��b4,�;���&����\�5b@��2�]�[
��YUy��f����0�S�/�銽Ub,4|�ft�ā��GX��p�͛���Mi\rza�+^�����붳��~1��W���,g�U1�c�*���U��{�ֽ�*2k6H�_��);�w^�Qo,qE}��{�F0�a�p�]cM^�[���w^����K�Z���}碻"�`7���6�� �JJa1��5d�;����pC��i�M�x��׃��`u�,���CH���TP�pw��EFg��RLW����%��\��:��>��#�tT�(,re��6s�� o�*�k�:{DDN�#���d����R�Y U��z�8|�Օyk�q�wA~�6���Eju;Wuu>��s˻�u.ޓ@���5��X�s��5��c�J]��
��-кzo;�b]ZėW+�}���%��US��T�}ϻ��㈉x�->���8����J��P��}��k�>8ﮛ](N]IC��f�	�U��S���A��Ƹ^��|݉Zk�j,S*��և;���3}q��;B:��q�m!W�Q����j𘥕LĽk9P�B�2U���AmN*���<�7.Ƶu���IѠq��3�ź��H劥z|�\!0�����b	�O��jve_F?)�F���~v��qv%{Ժ��㒫����v�/�<�c��F�AQ�:���H���n?��پc��(bӛ��)�|��ӄ�J˪CyWR���1V�sڌ&�i�bx��W6���5Cᑍ�Wz��j�0���hzt�W�\����>�Qݧ��;2���{:ѥ���w����'!�Lh�H�w{�r��@�&��B�߾�Mn¡3��ؖ1߱��{�8F�>������.��O��窆�<:I^��Ń�Hw�bT�ٵ�w�^��]�T;�L��R\op��3�i��~�tx�q���Zl�Ώ�eS�î�a���r��F���`��clal7:a���My��&��[ϧ<;�Ǽ���f��,�&.[���g{-�V�Zum�� ޭܜ(1��G6n�V�Ȼv�T%*�{�#}+k`�\�� Ɨ��g�����`M��rwu*[8;b�Fp���7�d[Ƶr�/(&4+҅���h�l�f�]r|�gm��8V�m�]or����]�[0t����N��-����EL�J}s.([�i5Z��u��:�(�g���on#3��,wΎ��f_bm���;8�>� C]̙K�ݽ�ޏh0
�����Kա2��ŧ����9 8ʾ9Y�� :�T�8$���c��mv�7�,�ɜNl�.7�u6e����Ҧb&�1�uX�51���,a5d*�ڷ�٨�80��'m��G����s���pz�Ct�����P-�JsMv���ް�!�tnH��x&����ct�ңu,��6rM��� V���跌꒻�@B�2���T��R��e�pWn��@�������a/#=P�7;{����Hm9X��+ӗx���WOd�+�ᭈ�`�QM�����`����nĈr���s��n^^�L���.�$΁�
�ϒN�j:������O�M��Z<l�Vdkc�S�`(�R�6�/Or����햳0�M�O�u�9m��Ք�5J�,
zA8���p�u6��wwJgs.)[v^��]j�(7RT�1X�Jj6�L8�kX]��H5{Y��<�Y�D�wb���T��dɴV'&뱵���x�Sx�__Y�b�
Ff�f8 �Q�]����&��A��jkV�/0aZfo<m�6��Gp�[}\3Y�F1�n�︁�s\Ô��R̕��ɟ5�u)�CZ��p���.�[n�DK�l�֞��{�k|Z��K���uee"�����{^;�6ֽ����g%͛���ևkgW'G��n�",�GsMs�Vo���cǃ1=����qi�Bl-�fe
a�Y�,�Ty �_MJb�z���pvhm��m��{km�����v#B���{*a��;7��=~R�{�jQ�2s�RYE�wK&Mf�tu�(�Ǒ�4���G��#F�����nm�'�1[�y�����ЮR㩴��h�פq�3dr�P��Y(ܤr�WW5�����k���<��W�P�Dߞ�7Ɋݤe< ��6�%Z: �����3�DE�]��H��>g��T�+ O>=n���ҍ��]�ƓN�ή�L"���H�S븰ܥtwo$	b2�=,���өuۀt����9*ͼOc�qv����N�S��96�]Y�ڵ���iXs~��u�{#8i�1^�,A\�>����:���gm���KZ�3��w�)v�xK����ޕ؜�V��i
��H/p�� �MQ ��q0�f\�MDG[�N�S,�(�QDD���"�4�ĭZ�[�Vj�q�
;h��"�2��M3��r�T��DTLd����r�+c�UE����Q��"���*���QXe�\B���㈢(�[ITU�UJ���Z��T��a�JTjTGm"��9���*��iVDb��UѴ�TD�TPE�k,`����-k�1U�ҋ��Z��h���Ьi�1��R�Q4تn�E5jȊ�Q��1������q��EATF������+
cFKJ���D����QV9KiX�� ��Ҋ�YQTU�Q+(��T*�P��b�DU���+m�*VMe!�
�Uj*ĭ�Fe+��2��+-mH��2�"�*�B�"�VT-�CVY&[F�%h#R���jV
[k��E�`��u��%���g�����ۼ��y��k���M!G�����A����.Vu�ٳKa�+�hS5ۑ�r�#�xъ��{�1ڻ�{ި�y��ܓ��>?c��1�ғP�6F����ē�	~�C��!R͓�̙�Ԝ\���`꼌Rڹ���X��6����&f
�W��`���3j�yyhAˋ�kF��aw�T�A���@6���c�Ʋ�G�ɜUE�c��&��;�(��O�p�x�����r�2!�*��n��fcҩPI������ĨpP�toh���m�}RMf�߳/���B�	�FC_����A�Ca啞TV��)���.k�t!������Ue����v�u����2�O�N�;�"�	u��K؟/Zg��B��� �ر�0��f���9]X�:!��!�G+{KA��\^y�����K�_� ��B��-	^�w�s!���s9��������8#6���Q�H�X�B4����ӗ�U�*���S�����Tlf��m�{-j��&E�\8PRP�r�l2���A�w8
H���*bVNɨƯ;h��W��v#Q����1���R��8!\U����l��wk�hGzWG�������^p�6'�Վ�;˾F7�\d�!���21�,G�~��?D�pѵ78�i�̭N�p���唸.k����^����6;E�mg�¨7��-5�e�9�R�<#���,�=L��bgPi�9�T�Ԃ�g]
����_W�aAL���Hq�'����<���%�RlE��T\sU���qVG��G�X�����d���/�t��C�l®�2v���<��Ԥj�>jy]a�V�SʰxQ�^�ݢ�W
�<��݊t��F( ���T��h������<���r�xk_����._a�r5��}Jz\�CY���Q�A\C��sl�+q4����5�X��}����C嵪e{J^hI'��S�0/f|���������zX��]P��gΟj�=*V�ԩ���av���Y�E����#8���^T���+��"6>2��.��cg1�/j��C͇��źs��?OW��F�j��tp�2��&�t�g	2kt��w��bV���,0-co�0ۡ�{�&W��6Yb���T"�s�a�w��[}�r,���=�<I�>��KO��Z�e�����6�C��a��� ��Qr4-
�)"ۓ���H9�mjZO*7:� ��
���X/9�%���n��/�>G�j����J�fnl�TwFt���x�7�,����Q��>H�cWn �i}Vs�$�P�:fa��V�D�Y&����}ـxQ�~�m��ô�jS�.t�;o[�O�=�#ϩ�ժ��wX;����h�(G,w�nL��4M]pHhz	�R��+/����`�n.���F���@�|��>���8I.b�w�_9Vr�
�g,L/2���ֵ��Һ���F���'x²��fͷ:||i��F�Qٹ9��u�V�u
7 k�ݹg��oz}1�a
�6�眡h�A��Y^6���aI��y�uwf!~���'Z����n ��b�#H���婄&9L0���$N��NRR��ks����V4.'���7��bQۊY`+�����Q��p��\3_���'�e���*Z`�q�Xu�OB��.4�U����(vVUڧp��j@fSݚ���z�����۱�Ǒ(����LR\pޚC��a���oOT+1��bt�o2_WT�܍�������3E1��}��'�4�%���(��i!E�������Un�RKw��.�L1P��3<5�}��Y�%C��Dg�N_O7:]�(�hp��/�ϝ���������u1�&�S�sve@%��ѾH��l>�����r7l��RX�!ˀ�X�GI�f?<�~y}xH�?8��̊��P���%��E�#}	�n����r]�/n�n��RmN�KQ�3���k�Sys��.ӕ؏)�/���a�\��}��]��Y����.�JO�XЙ�Z.D�{7wB�g��}^m��_�%����th����]G����������d�u-��@dca�w*Կ4k��^cW/�pc$Ӛx�oܑ����=��C%=���ں���s��U6Os�Na�9)Z�B��q֪(��H�Q�u	�AY�����	wO���N�p�u�wI)��Ǫ'���IG-��B��!C��:Q.���|#�q���|'�"�PP="��u�U�s��Uy��u��H���;u�^{ft���5K���W�Z���^������ެ�ŋ3�%FϜ���q�&0,����T�ѧQ�3c8���L�,�/���#g��[�y����W�U-���(
߹������2�~�t�.$z��1cܧ�7��L�:Ή���>GF��DkuI��I�8�<HJG�-�5t6{3��mscym��+�3L^�K��*R5�ۉV{�Gnڮ��[�kh��$��yc������「/i�q�}1�z�"��{O�9m�'��GZ��Y/:�)���`�#DŚ9Tz��<v�z��wm�಍����n��-���d�H=S���$���MN��>��(z��ҷ����a��e� uT&���SOzZ�i�|Ký2.�a��[Se(�A��Q�����
��y��[pǩ. V�rTd��G�����N_,����1b'ݎ�Z0��{HW>�"��,^�����*��GV�qV=�����B�Inr�(Q"�a~Ǘp�ٱ*�C����^9�l_��F	5���;�p*�b�b�9k��đ k��g�\�zg�^�+�y`�j��S\�)���*ƣ��7�bjS�{'�v�L�ٷ��\x`���XZK�>x0�?�
�����3�������n�+�6v�S�L
���6�_��ߪc]'f��4FԺ�9�wh;+�����r���`�o�.�;ˤ����a�p���ɘb��s�J�b�	㢱%�sxY��Z��e�Ϗ�1��<�`����+�Ƅ/�eȏ�2gQ}�i	Z��og�2�׻d����ٽ�U��T��q��H9u�~��2{ѪA3�b��ɨPXF��z-�6��f�׳4.��b"r5�Z�J&����^����<��L��"��R+���L����{|���v8t�9&FBck��>�;~WDFS�����q�P��<�_�:\�H�}��!ꠠd���0`亸�Md_f�ӛ�^VͽZ����W��q�N���Z;
kHM�F]�A��\=�W���њK],	�%s{'L��U�'O�rh�_}%�����:o<��t�Hwӱi�/�r�w�Ih�%No����Jz�t��ݓ�j�Q�(B�7g�MM�����^Vj��ի�@�X���Ws�Ȏ�*��`�GA��
�l��d]Q�VE�{
424l��*?gl���[|6��;]�2���I��LC�n�i��Â��{VSl�鸄PzaѰs�#z$d��g'rs��t�˅4�7�V\�\��eI,b>B*-K�P�'O.������.����گS�d�wy��}.пWy��������k�ih5d{���P�p��y����s5f)�y]��;�̼3�|S�C�q�[�X�l�[�O�)����X8Tڼ�>����x��͘����!���/�:j1��&&"}Ŏn4�~͛g��֨�G>x���d^k�秖��e����|�	$&�'�ߙ7�-&�����׆,[஻���Q��1���:����Q��8z�}�B,`���S��.�3Bؑ�&���-�AV8��mѳn쓣 ��ǚ����B�������.��DJ��A�V��m��'QIA+�,�:�Ŷ�X.l�92�2Jky���oT�d� ��I���G���y;��woJ��*mq7�\���ky�#�YN�"��؄��BRϧ���&����������͉Ռ��:��gR���mt��D�����T��������ZLh���;7X�1Om��6B<h}v�*��4᯹��H����
�	�s����z��Ќg�F6�a󪯻fW��7�Yw����C�f�XɁ���Kw3o'��`?h�aW��>�A=2��r���y���b�K�gm�3�y����gJ���η�W���Ƣ'N�E�P�c���H���5�un��ݟt�t�f��{���8��ú��>P��0��G	#��T���NU���DE��P��Ν�n�ZM���kwX*;k����+]V�(����>Y�m΂������[�G1Zɝ�ԅ�̫�huߙ���K�f����/����\cB���n���8�֡��j��Ж~�G��3]�:�jm�&�mL!��f����mj�������7E��5dM�	J�z�u�1(��,���[(LAW<���|<��x�+xL��5pH��9�Ύ��	q<L*���r��AB��s$�.�L%3��q��ƻ��rT�P�L�X+o�DX� {Zђ�<����<����s�z�Ჺ9SO`�9��J��sFg8�W,�Ʈ�Z4ZEZ���mE��5c��[�Hr�Gz�p6��m4If���^R�3j�1��鏷�����r�sv����<�vho�ݕ�p�z�׺��9�s�l&-
.8n4��"A֨n\���}in�=��������2�Wʝ����Xh��s���@�:�Ԩ�'C�u���k��_Y�X#�ׯ��1!�t���Y�*f�#S�����y|eJ��w3;p����<�p�Tj�ڔ���_xxsGڜ�ߝ���C׏�����?���dv۴|z��Doeo�i��\<E�j��w	�M˕'*��v-�B#(�� ��Q����sx�P���8����=7��3dZ:��]^P�͢<����-6I��e�����j!�Ћx���?ry��Т�1*����}(tAZ޲����r��O���#M�VtU�I�1w�I��rGlz�b1i)d��`k�W�>p��:ϡ߉�v,��m	��̴����A�P�q�-�;u�V����ѪY3^R�5�,/G��.��f����c�@���a����4�y<X�C���	u[E�s��|a�RŲfj0UR�(�)"	� ���t�wll\��`�"����v���d�Ǎ�4lbMP���q����1G�}��C/t>�(b��sy��c]^���ŝ/n�	u��K�އ���g�;�L�-�$�\p7�������RV!�&���V7>��C�U���8Mm������Ϸi=���w�)�g�R���a�)�*�3�e�5	ғ��H�B<�jwZ9�x@����Jc8��Ҹ�S3�w������m'2�	#�OD�kpUs�b8��٦\�c��Ż�ޮG$��4׮��[�ה7��B�ŧ6;�����ƙ���S���O&y��:=��ߕL���A
��7�Rh�.5�p5��bZm���ڙ����Z�:Q `�����~��iP�O4+�U_��Ve��hUs����ڭ�I�ԅ� �h�R��}ef��zϨt�~�4�Cؼ��(n8kB�=-�����hP�<���h�X��x'���Z4�Lu�����\=��)BYsx�qk��\���_?xup��\<�ɍiђ�#DLT��9���4\cHf.��`��8ZL��}RAg.�� l�� �/���6��>L�*P�1V)�'���>lq�$1�L %�'�wE��N���Z-.��|��D�9��@]5��i��v���]ͳ4>C6����]���y�R��@I.�Hqa��RJy-V����PκI����B�ƃ��ه�d�ss�[�l��e�[��k]�e<]�5vo{I���q�֚�V�;�D��!z̶E�HL��)�a���qB��n.�Od�s��'q<*Y��
�G�7���8U*�e&20�ĨpP�[o��P/1&��u۷�� 둑^�4/3Զ�J������XAف�����ި��2%6��wa�/�޾���}DIOO������9Z|��gSDz��Xbɽ2�ᐆ����x�o^��s�v�H9��VF��&�񬚩��M9�ďV�� Eں�* �L滖�%E]Yh�������W�U��3�3o���[�l��Ѳ��\@l���[���%^�N�Xy@g�m�g���h%
�YLE�+:oȠ�ã`��`�I��0�e���{U�s���y���O�.�c��ܓQ�h�[�
�B���zx\3���+�60�/�B�Vj�))�z�^�{R�t���yM-���1x��[�+��;J�͆�;-��ݣt�>�fn�X��U�A�Cm�ujR5R��S��𫯫tRc��N����'�,2��ٙ�SNu�ī�`%h�#s;�0��v&�1��po;v��z�
��Z!y�f;�%��CE18t3��ox1+t��e��띺�n�2�.\���
�S��%���U�K�z�%ѥ�Uy��裔p�?�*�\��I�+nhm�=��2��UaWVqA���Ѣy���t3�g�Z�J��c�S;΍��y�ݐ�F���x�V� �ki����v��nG�V�yohbF�lktp!�,�`�+�08YKF�"�mf�v�
F��b����c_[t1bTtu�e$EF�
�*@r��Ԉh�̳%��!j��:�γ#pJ��te�q�2���&�x��q�ų���]�2�A[.X�\����㢵��E�b�ݮۨ��С�������q����̈́LV;�4�eh�n��X��w�/7ru��R�/��)ՒI�.�k)3p�=G����A�G�{Q|���g����/EN��r�C�*I(RH����KV��+���)=�I���=ò�ЮՄ%g፠��M̸GtS�a�c'P��u��0nNbKj;ֈ�
 ZsI�BDy`׊�k�h=�|z�.��T��n)��c)�25M��F"v:q�5�)j�RU��khvcw'�%r���|� �!I��su���ԩA}:��t�Z
r��[�ɴ���[��V
CXW�.n�فg�Qn�N�p��2^̘ ���̘"���}#�ooSV9�#Z6]8hK�����t���a�Q0w��'i�ٓE;�m�z[pu��bI^��gU�;���t���Y(��,ջ�u�R��_WU�Op�鮤/N�ier9�Cz[C M;y�Qf�ؠu��u8Yu}zNʜ�Zx��sR��{u�f�w�uH-G�� ���x%�RgN����ӷ6�J����b:�U�^�;�hE\7�f��ܩEAM�6M\����H�ZsL�#If�wY"w�R�IN����V7��9CN��$�@
��*���I��R�Ix��8�����T�����F�E#K4�'�����vr,�8�M[�Df����2����.�yn�\�L�v��1Bi���%�vNƾH��W���d�a�1,���.��췛���h��+6+�Ʈf/��0M=�#�D�(-=�X�d7rG�L�)�Ã�E�\P��>,)��nfe���ƣ������NȽ&9ɞ�O������up�)l@P���Tٯ3�O��Bb��%�`;��.��#}��-��{�D�up>�N�]z�q�Qځa�"i��I�Յ�����Nh��]�W��>8���c�W0R�#���` g^�5�-%ikc-c7�N��p����q����ʤ��o*mS�3����V�SOLсv%;�z��k�k��g/��������k�;�7Q�$��j�sX�n��u��5�Vgئ��������dÉ�t��tu��v�=��K�����~$�H6�
��3�Ө��QVKJU��c2�
���GV��r�j�F�µ%m����V(��s1q�6��Z�V��
�[@�0.Y�ʤ���3�
�$�TR�Mec&Zk(ZP��s�h�2Ɍ�HbU�ЫhQ
�H�%�Z�e31q���J�Lb*VA�╊TS[j-BVM%Eƣ��j�L�ZU�TaSL��+ir�&:h��YY*V-�X��4��r�dR�G2���0�B��	
�+�+KJ)���V
�A`��[s.�UE1(���b2
eAE����"&ҡ[Je�#l����!����`�B�j"�Z	[+Qeam���L�5�J0�*D`���TU
�\ʬ�+�IZ�m �R��"�mB��11�E���h�VL�R��P�C�{������㎯�Vd�'��Y�Pփ(k�Z] Z������nqmIf����!+� v���^7�k�wLM���r��>�نZz�@A���`4���h��=�6φ|�x<�T=��{2��͵�H���O�9�[1Aۘ�o�5��Z�q��Cg{׻&_\��o���ߪsգ��t!f|��솆�4y�ʦ�a���=:���٦���yY�F-OM�=F�l��ƌзw�JXǇ"�5yS��/�C��"R���f��bE]���@ϟ��} W��YN.���ϰ�Dp]����xu��b��b"�[�+N�FE�o%��މa�W���=|Q���[x�1�Ӓ}���ӆ�8C,_0T��_v߇y��>�I�Z!�)Dף��	d��,oHu��s/meԠ/-��+~,����LM�+H��z����YJ�|�u��.&*7:X�X�]��ἱ��)�Y;�a�^.�8�zp�~=�r��t���>AӖ,u9L�1��Ɖ��o�#z(soe.���7�GYuL�+g�z5�^Mw�}r��U���!��|�ga��`f�5C���\]���SX �n�]�׊tw�g�!��`!�fSuj\�����b�"��F��#x�vN^�`nEO�A-k}f�̬y��Љ�|���k��	T�P�h�bRʞ�v:����ً���n���r*'�D���ޔt*��;т="���z�P��\��'���>�|=���ٶc�tX�YP9n\��d�ToO�C#\�{:�
Y���1^ua�=�$&w7�p�*�y}��F�^�P�*I����&��8�!�vL�%9A=�t��ʋr6��Jxkț�H��~g�egw���Q���y@�I���˹�Kw�j�2����/��+C��P��8V���i�*J%
�\<c0����*pI�Oe���u��搌}�&k�O��v9�4��,^��e\���������#�{�zce?\�gd?K�!��5�6k3+�������jt�=�rz�@���m�l����{9�gڔ�S�X��Q�T�Ի����	�*|�߆J��ΈϚ���F/)`�Ǳþ��٫��U���w��(`�1d�9cn'>��f�+�#�bJ/��)�;E9��v�|Н�8T�!�ï:�E'$q=N����Y�wt�|�/(�1�j�p���(V���+�ag�g*}�b�ª��D:����^�I�xi��L�ߴ�%k�'5b��m{n�y��}���i���YH�Us�����J1C����BLaW(f|d�t��AfV����yv�|��y].�ɝFd5,�,��c������-��ݽ���]����AH�k�>]R����*�3�|y��J
<b\L\�J�hj
�?��]��}����W7�nr�ĺYz.�]�aZcC �n@���4")`ư\6]�����w�NNV����Wp�ώұV5ĝ9�׉ib㏰O�K&Qa��V�WP�r��u޾�v�L^�)b��y�QC��_���e>6,屿��f���3٣s,nX���4*��o%Nvf�ҏ�{�֚��5�F	�����*�Hd߰�#``�������������ߚ���鏃E��u�󞓁�X��o�w��8��Y��z���Ŭ�S�q����S�c�A�;8�^�>#,b�w(F螮(���n@��l&_������Y��{�j�ڌE�䲤�����9��޸Y�R�Ǝ�W�����D d)�Ԏ����f�s<�״ʫ1�	��:"��X�j�pnc��}��N9��g�h;58����zқ��w+�uӲ�'"��q��x͛Q��D1q�P�:���e�v�:a�D����=G0[�C{���V_S�u�:m�\�E(l�����Peb�
�s5�����]�j.�
@�XF�^��9�fVoؔ���t9p"��K����t/X٩h�;��yA���Vgv����Z��T���޷�G9ƏrI�k�Ł_�)�x.���,��˥��>ͼp��kr�/�P����9P�|ס/'�����r;�7J�)v��O�_��ԫ�Շv�lۼ�vK�Rg*V��7�ו�Љi���T#q3'b���A;4X�#DQs�o"���-��*	w�F��\�����Qy$�[(F�3(sY�#!�n|��B��1X#�(�Jc#��YO�;�+���f�F_��)��X�I�BEH��̙�P}2�(h&a�+�h}��Hf��3k���\`���#Q��/˪�@��yU<<O��j3�P��6�8󭮝��P3�(�`f�5x��C�8o,Ux�G&Ą0�gu�qh;{'�W�m�7O1'��"e8}�%�:��ht9Z@���4EM�[��0�7�О�hKL{�Qm��`�Vcus����u�vE��'���5S4/��T��^�G���(4�N����эw�=�u�*�>T_�j����ׂ�L�Ob��7
�U�LY�+����௲�f]�Ȕ�3O�����N;ViԤ���.$��Ȝ͓�f�Q˂G�� ��I0�ͱ}�I�d4��8,��[���;Gr���V�.֋�e���3�W|3�e�=�5W�!��8[�k�!�x�X���+5��i�ݚ+���4�2���Xq��{�9|(�U�Hf�+C�C5e1�ΛE�0>t�Y���:�l�;H_�Z�ʫ�rLb>B))s�!	ⷥ�.3x��	�3˦���4��ܜu�?W�p���s��8�7��c��W���ʓ�/��r���[��E�Z�iS��p�/T�N|Yc�L*� 졽�v���JF�c槑3�v\�w�Fc"�x\��^]X�ݔ[�Ѕ���pc�<�s�R�>,���d�yx�8v/�����=T�m���q&2�Ha^���Mg;c(���byͲt�`�&�:�ݖ2謊�LjT���$8�����wk(��tp���4�X�<()-}ULL�8�s�o��WS&���`fĺ��X�Z������G��#<b��6j}�4OȕF����"���9����>[�z;�[	�����V����I�\�`�8:�E�W��e�5A��cV�Z��e{��.���hZx�����se�N(ÂQ�W�c��'��+�N �,��衵�][9uR�6e��י���մ�3:լ]nk}i��v�Z�wwkX�ΰ��i.Gz��Pj��V^cǦ�$1c�~�a����))�#�Z���{x�FN�ƎHv�����eM��B�����\Ď�w+�{F�x#�m�͠Q�wϑr��*L��G"ޔC48Kȫz�w,UQ�;�w+��_�[��'a���I�N�Je֯e��P�^<W�Rb|�o=�E?d���< 3�H:�\�F/��;�|6x��}���X�UX�w��s�.��uꁗ�¯]���Eۛ�pu��C AǦ� �޷Cf�y����D���c'��hO�k���7<ݍe��^�>Y�[7���1�w5C���pQ������'5�	�n��\C��>'�5|�yWY�<sB-XiJ��y��kYp4,.�W��j�e��
^U]��w���]�HW_*�kb�|-à�8��T�z�v�ژA��A�S�o���ב6%*���׶��R=���Get� ^�/AT�m7A6��^A���(u�;�)��s+\�鸄�%��Us����႟S�4Y̶{��}������.β��[�8VFϖW�n�{^�;�u�E�05&-
�GI�����s�CQ��h�Fcۄ0P�5��E��i���	�Ɗ��e8����k��W�bț�g�jV�X ��.W����k�́.��.��ˮp�e���-|R8�#�����l�J��DRҤӽ�\�G.�B�:m�:q;�Lv;��:�m�W[ˣ`VMi⡔8�_��V�^�]#��wq�L�/R��5bVQ�Uv��t�� �5*peƺb�M��x'y��y�]�{u[��=p��=�����ƛQ�xd���zW��@��VZ�~0�?q`�s@M;�\kJkFi�:J�=rPt����Թ�8�w^�V�!�`�F%���>"�|�N��&�ژ�E�!�fT>�E�C���)ڰ}��ԓ�*f����!�·s�������Tn}�ݸy��ł��,�E@�B�X�+���p����cz.�9%��}�2z��ԏ��i�(y�wĥc$�^��` J�Q����-ߤ�v������ FiDX~t&�^<�'�#�z�,>O�g/�/�m2��IC@��f��V�[����bv����p��z��)��ˬڰ�i�\/qu[��a��=�$�r�ϖ5LS�شM;�����A)�^�<�`�4��&d2k���e�o.q��	�Q�e�n�^��,���59�{c��U��a��uQ��!�)�:��2gu��^�'0K�=�q��*�zs]=���	�������[h"m]�n����Ȑ���<���L�䕉5���2�ݾ��Y9@�.���m�9�`/0���Pv������?I3P���!��9jk�� G�emmDk�Y��)F�,�:WNO����c�vq���|i��/Wr�l���*��$���og~'�R'B1G��{��xF����s�e���g��j��1^�:5��IA�h�b�G��g�؏2<�K�{L�1���"���	����W>�"���c2�"����mtn"��eE��� \�(��0�%a���q�0S�\Я	~\.Q���X�J�`#&A+���.�����ϱ	�P��;�KQ�����}����ҽ�-��xc�ggs�`��ͼ��FR9����Op��fR�Ŕ���O, C,�J�]XqX��6=��.�2�d� j�c�ˈ��3)Z����B70�v91��O*P�#�NV�y�-���܏�}���WU݆�@� ϊZ��C���*�U�}咙�)��ۓ.j^rX��6tF��!��<�7ι:V�I��I��5�">ɜR˼�_%��J{O������K���ׇ��¯/+#���q�=x�/9s� ѭD���=�qB����8nt�4|�u�񓫰�Sp�����=8���4j|F�W+lp�U0�t��/w@��ڄ5)�;kA���W�wD��8�8'�%�O���'�l��jY���|]��zek�9ml���]N�e'�gM�����Y� NO*D�<��5x���_�8o�	���Ʊ�-���}����wRaN�ԝc��8}�(��v�7�Lmp��ӷ���y4�VA�wסL�{�|�Z��KL�3���|�{]�b�Ţ�<�pu���w�f��i�����8v�{�x�SҨ�N�.C��n`	��ۮ F�ڦ�*5ڸ�R������ێw����#��]��D*�jl���h���,R������3q���
J����+:PA႓z�� i� �Y�0s��� �{��&�x9B�eU�w=ےhb>B*Աwΐ�'�<��ӛ-u@�T�:��a�	�na�ٗ���|�-[�$�*�-h����(B�t�֠��V�Ժ�����H��F3Z�xͧ^.�,y	�]�b��e���jR5�%�?*�赜�վ굶�k%�b36X�s���l �MFOuP�Xj�M�/���awh/T&.��uZY�Q��f]���{$0�}��&���#D��ds7�@�X'�\�
��dΏl8���z�wT�GC��� �)j�&$�+�5��wq��＞ν[c5;̎-j:�{H�iے�S]�,{���{�/tNq[�,M�;K�]8��\»8f�dp=a�ᢧa"�?�DQ颯�ÙWI2�w^W�W�
B���3q�ܗM�S�L0�~*��4�գʼt!f|�����A-��S^�=t�!��vR#��Ŗ��=۸�s�� �N$�S�L�J��a�㑙�d�͢5����S��'���0K�a
U��M��V�B�t&�P��ٿ����+ҡ����xлj����b�S���������_0�:AוQ���ɳ��\�f�
d�ğ�|���\��#��u,Pߞ��o��`������J��,DLs�҇�˭^��{k/���b9H������v����01s�Y�C��5Y��i:�t��D3b��8r$~�'4ʉ]�����9���v�>�d�Ls9�{>W�8^�4�:R���-�"�eo_;n�+�r\jC�&�����q�V2}�q�{�UY���y�<�����X�u�<�>>�ܵ��7k����.������'5�	U�n����A�b֢^5���c����3�������k�rd���¸����+�a5r2���	�*�G3����2L+FQ7�]�n��q��cW�������+cx�m�.��7D�`7�w�s!e�L�_(7;yl�9尊X�f`|1���+��P���q�b�n����4U+YiΖ2­t��}D
=>F�Y�șiA�����^�hAxs1�M��!���B�u��g�ʐ�Uۂ�Y��Ś#-ԋ�(>��>��N�$�=F	���Tf��;�M��/0��x��spA�P%[�*��r5�;��:H�ѣ�e%ݼ=��o��dsG#���L��R#(L��IW>��9�<ɳ+Q@�w,��0P��s0e��bçZ{�ܥ�Հ���{b����dM|9��.d��o�GZ�T�h�xAܹ��E-~�SGj��|��E9��o�P���f�Y6i|�VC6�:��
d����]IĤ~l5�\'�Q:z��p�K��xL`��L�Fj��j����zL#.\�FVe>4�Ӗ��͊黺5����t��`�،u���R�hIfvl�����j�̭�/$U�u�	P�YhE�f�3,s����|iKG@�l,Kqv�ب]��-��}��
�avF�����Y�g�<)����x�@��A��NVT��9| fu�����S(;4���^�ٴ�W��L����Ml�.a=����e]w!��K��z��+/@�����o�6��¬2����] 	�_#��X�R�n���������j.��J�eӾ�S$Bq�ֶ�y|�5S#�~Z%��)
e�=�ՙ�m"���y�P�+��(ytc>�gDiw��l�)�9���h�?������[��n�z,�6T���V����{����Ek�x�zT�/T��Wd�Uv��z[���y�2�ں�eH{
�Pć&���ڌ�$M����E�����XKB�����V�J�DS����s%�`k������X�ӕ��,������[��lwE��\�����s7R��)c.Gg&W8��h��U�P��W�2���v�������Bt1��v�1���I�@��r]�����_��Z�A��
���%Or[K�����ר��g{Y]A5��Q����h2�]�I��k��l0��oe鑱d��Zsw1�0t`޺lI2];�>�d(7[۹)!�dY�}�i���H�d��5ґ��[3H)CŁ��j����a��paؑ�>̓��;c[�:�<�c�MT,^��@��`��1���胃 �wh��:��Y���d}[��m���h�gQY�8V��9U��=������*#"ͮ���T���z���;ZQ���g~vH�IQooMa8�3I4�P��7��ee�U��Vq�ir��MSbY@No^����b�Ũ�]ԑ݅�Nܷ���P�Ru�.�g�U{6��e�w�=�ׇ��<�	�;�ߴ��5m��R���;�Ju%)e�_xV�y����ח�u�p���h7�ɹӸ��Y�W�?��@�I��-�-TX,jҲ�$����%EX��\ ������T
�l�m��* 9C2�UTb�@�Xb��2#&0�J��e�
YU��mU�R*�����1`�6�FTU��,*Q
���h:��C"-,����YR�,P\d����X1%ek4�$�j�J��*���E�6�J1t��� ,�*C��B�$rŵ�����*-E�+��j�+�*A�`,+-�I"� ��Q�%eƘ�m����XkT2ڂ�P*֊J�XTX�,�ȈJ�*V
,�UH�)ua�0Ab��
�����T���T��mAb�`�&�L3Ud�V�Le�X���h�j�����yH��E���u��+t���v�M�	e�c�A����P*Y�+-v��<�qJ���᧊��
w�]�_�x{V��NK~<S���R	_fF,t��Q i��1��RԔ�0Ҙ7�~�¼�8�,��ãk#ï�B�<��X��y"*�����ݮ}y���
Ϩ;�9�5��<���f������c��O�Zw�T5L]w3��ii���s�;H&�yax~��g�6�Y]L�,�3�_ίj
cCq^��;m^4�*��x%GR]F\k [<N:��I��S̨�� �%���c��r�9�	��ns��*��{E[Gr�Y����F�Hj��f��v���=Yv�	nI�ז�ce#��[�Ԫc� �Q����MEӥ'r.��hK��۹H�AR�n������e�X�P��h�eC�b����>m�&���s�Fg*��$]-�g[���{����q���@+>F���L�&��4�4'1�l�4rl�����=��q�6nD��;X�˖6����֦!C��(�C\�%s��&�������da��U�'#��չ�jdVV�φs�H�t�2����B8���!�t���2��r�xK�eգZ�BzM3,ǳ�/S��'m�wq��M�e�d�$1q}Λ���_e�
�SB�]�x�r�s��*W;i�ߖc�e^�x���Bl�Z�n	�6��:�K>>���O��ʿ\��g�cx�����3�I�İbW�O��*�{� D���ab#�ش�O9:}�n˫��Gr��cy��p^�Z�c�����^�۝�#�c��-��Y(_c��V�>_N�?%XyP�t�j�О4�u�N�hJ	�wq��y	���"�`�	c��3�e�5	ғ��4"��y�ʻ�٭��z�3����l���8H��R��>wQ��
�n�s�3�E��wHR������5�6����>�Qwfّ,멈Ca�T�P�#r����r޸Y
^��i��;��k�y�٘&���z��ƌ5�6w^(�b�^��d��̊Ja*�i
�}H{"�����;^�N^n,��rN�a��P+�N�5������;���Ei���B�'�	�M���[W�Ҟ��Wݱ.���`�0ъ�c�T,��
�.���3�^�V��*|�9�Q�UT'��Ҕ��]����KU�7"ε��t�}�<�+�XZK��5�ቆX0�]<6�
'u�m2�e-V��e��Ej���`����3z�����s;��,��.&c7ET�[^���*IQ-N>|,G�R�kd�������l�v|�l��4Wf�4���ڵc!��5*b_vN`�X*-J�#�Q�e�����u,ڼCʅ�n�0�J�1�����<)��:yR����)�ޞ�ޕ�1t5�a�Y�&��b�tT��^I%�l�(_14ͣ!�O�(ԒZ�`�@:�����r�{�����݊t'����o�Õr�	^�e��	f�!�!�T���O���`Z�w��ܯl�$�*��9�CkSU��G�WA�ب��f�z�x_���S�/JGʏ�T��W�`(=:�,��$�"4�x�e��ו^0�TY�z��eŃwP��[���7XO�D�B�!�X�����Y&E&6��Ӛ����ËG�R���;��|LҴ�L鯳���d�H>��m-"tvx�MU�������tM'��z)S}�����(z��0y�m�#"hS�j#]*�ES���ێw��s��ql�'y+��] �o�=�. ��V_IeVW.��V�!�{VSl��c4M���6�2U5�٢�Çs���oE���ܪ�ع�[�̈��?p���疍My�&��2�>���1n�˥ȯ"��.�eLնr�3������f�2ۘ~]:Ц�I��Y�:��Mf�Y� -=�1��v�"� ;���a��b�N��y"?\�,Ib�lscz3�Oc퀼������]d�͜���Q���N��z�5]k,�y٬(�o�/�MK���1�]Øb'�R�z�#|r'Ɍ�I+���&�Y����U ���L�*�d��NM]��(4�x��F3Z�x��u��X��
�;(o{U�_����b�\c���=��T�<n��(FW�i
�1�����nt�; q�&&"}Ŏm�{�{��i^ֺ�R�R�Z�x{��1>֨�S�xz�}�暈������� GK�H�Ֆ;�u4��_�m{񠆋���b�3k(��t�o���R��V�<��S��9�NƸ�N�9�U_l<��E�5ű�s'RuO�2<�X|<j��5��ȔY�h��F��1YѼ����7��J��7N_u_tJ��!�okψu�~�p�4E�5���KQ���M�[�k2R�t�s�RƐxDg��:A��%�(ÂQ�V�i�>�z�~�U'��G.��v�7��~��ބh����"c�҇�˭^�^��^�~�K7y..v�J�������bGaXk P�W��$l�J��j"t��"�T6_��_��#/�<}ۙ��n�C'�k�QSF?�j���>ꘘ��R��^�HoV�h�Ն��9��\���ܲe\�����N��)�;R�<�	+�,v�MI���+�r�	U�S�f�gB6�K�:�Iԩ���h_wv[���{��ҧ9Wu�#��;MBE�7r�^{>W�ɜ.�]�؋�7��s}�������k�"����
�#��C��X�]�u�{�YІ���Q=y�y�]�Rfvh�f�$"��s�o��A���ۓ�45�� nUu�A�b�|L�_v��Q�Ve����w��� �M��(Z7��W��tB�����%�ft�@?�v�4����B��)����E����=��)�)�'y�a�Ꜵ����}�g�	_g��i�����A�hn�oT��xN@���[0mNv;�+��-9�Ύ��	q<:1u�53������L}��kO��g��m��C�q}���B��֧y���B}�t�=�-r����5��@!q�q���z�T1q���/�ϳj�}¯j��>�b���:���l#f	�9?�h��R�״�7�#���p��H{5P	�b�O7]�S�|d}�ڛ�k�vZb��:ϝ�Ζ��y�TE�Ɯ��r����Dn�X_j��"�o�����릮�0q��J����/��wy�Mz���-��Y��aOr���w�REٌ���Cw)EBVt����d�b�w]���ڂ�/%9M�Yg�� f��g5�3��
�7; owPeoh�V"�}o�{`1�!�uB{b�>�P|��Ķ{���7�������=e�*X�7��W��&��{_�!�)jt3jj�V������ڱ�:�� ��Z�#B0�fT>�E�C��DC_k.�ILJ������M��oo�-�=$�\�>{%�=u��v�Ʋ�Q����ʄ��+��m�S���&�3���9�4�2���	�d�~��&��DX�1<JW�Q.���]xʠ�[�3-�w�WK���4t��Y�%t��W��R�V9Ļ���FV�lΖ/��\d��ڋ\�ɞ�e��zh;/}#�-7^�GO�8�7�bcy�ˑxgvPE�"l[��V���(���v���p�E�gVJ��:堏�Zy��'�{ެ0�����
nS�F�
�ޛ�pH87�۴����w�Ja����셗��'JN���Ƅu������sǓ�{���Ez��`��2����|��r�q���"�wC�@���}���y��uүXi��;z�|v�j���Mh��qq��3|�[ٲ��{�[lxb�����\��6�E���z9㸛�b�mae���B5 ���X�r�}�Vwy�v���_���d��f�ڻَxs����W���S���ܭ=�r��W=�+���`�{7��j�J4m��\ M����o Ў��pg 5�U�!X�B��9ʃ␛98�y�˶��־����Ô;W��R���!˔Ϻ�c��^�i�-�{�OS��ˣ� Op���b�\�X����JdHҰŻ���n�E{eT�bt9����`��������ǃ�]y�0ьdڮ x�u���}��u�vחd�|�n�=óm�?�!V�����4����yK�S�a,�J�]Xq.��~��eMTZny,Ļ�8��՝�&��ǘ�<o0ʄn&a��q�}O*P�<��X��������9��9�whh�|r��fa�G�$�c�a��|hl.��C�gC�| @#y�u׎Z��j..�u݁A���W���|2���=�	A�^�zݷ�4�=!̕�9{)rؽ�O]� �OB��с�����~Q�-�W�
�h�޳AZ9S�X�j.^�irax]����� �`&-�p0��D�g���(s/m8Ἲ�rwY�=���Y&-�V�-;��XN9S&iO��%�X���Y&E&6��a!�WZB�fŘi�W����\ޅ%l�v@�UPe�~GN���`O;��vt���b��H�J!ޢ,�wӨ�z�V�Ք���.t�&FX�au���z����d��FL$�,�[\'[Fӄ���x��1eFs���r� 6�\���wv��2���W��|pd�ᒹ �t�#ii/<2j�D�2�Є�6;�Z}��k��s��s_���'�+n���1�wƟ�gx+���I�Ϳ{a$���\�`#�ȋ�-�ϗ=f���8�9�����hb(f��!B��ت�ǐ����Z�̹p��-\�)#X7Ϥ2|���W��l�fDM_�VN^L��BT0z�`4��������jg1����0���g3ʱhq���x��5T��3���������wd�w�hC�<"���x�-�g4�N�Yc�dGL*�#'i �e:E��V�:iiY�n�b��ڜ҄e{6���szz�zt�LO�<\�D�ݪ���܌�v�Ţ\��v�Tܠq�������^ʇE,4g��=��7I��j�Λ|�i�i�
�z\��{M4^FJ���Vy�=q3��c=ǅT�5��	�,S��Z=�0N�j���KS�L�	R��6x�ݲ�K�Fx��Ux�x����_��� �.j��8ގxԮVG��ШK�4�����txZ�w�.���X�����&r���Ң�}1V$�j�Nmjۮ����3����)S$g嘨!L��٦��7_vɎsz:��.Z�w���aU0�dH��u�.�;��}^��ۺ��z�U��t��6e�ȩAסS���^?$!׍����w�DY��ލ����6�h�|�9�Y��ϱ�_�J�K���:A�J�E�2l�ʉ�e��:���y^>f8���4�<6Yb�\�E���J��0�-��X��5�2�������Z��8b���+x3j:Z�>>�^&��H�D3b��8]���u�l�8�(�9�~�z��hJ�i��H�Ǚϝ�����ݩᒉ�F��$f���S�Ŏ��Ӳ���ݻmp�YH{x*�����=�����Ǳ���ppy��x\��P�o)�J�*S�9d�����)����=�B�N
�������Id�����ۇ6؜��*���1��ͣ�P�n+��H�}�n�	qf������º��ђ��"�(1��0T��]u���R�r�d�/���u�kbl�U{d��&wK��;�N�̡X)�Yg�I��W�4��U��]������b�Yֳ�)�Oh�>A�����P�Z�	�VQ�Q
q�)�o�ʂw'3�"�S�*��K�cż4˦�'�
O�X�&N� �k1��4���u�|Wgk��1�97�[h���u�H0�2��w5o�G�g���W_*
b�671n]Xʽ�WZ�%�1�����~�� �o����ܵ3]z|��k��g,w�5�zz��M��:s���6/�
��G��l���}=xf�"8� �>�A����X�m�K�j�)"�y�S|v}LCGyNOf��sԨJsV%e��XU��������Ep�4 1��N�k7pS[\*/UX�>}���Ɋ������ӓqNXی�e��c{�f��.���������V�lR�vmV��,dEJ�=rPu��W	�M˕'"�w2,��P��IJ)��5���R�_��7�}(z�.u�F0�ŘC̨x�Q7��DC���޿g����wy"�>>�����p�>�,|��.1�X����5��Q��F.]��7��#���_w�jݽ��=�hY�e�4#�����]3-��1WV}�� ��������#�(lӹMvjAV� ڏ	;N��<���P="Ϻ��yl��+vgK'�}oR��J�g�;.6x3P�����v-5qΎ/��o1�x�g��,}�Nd���et�x���ry����8l�C�w,r���,���Օ79�#o{���Z���q�xVgxz�Ɲj':��Ƴ��wjp�R�'V�.����7��w���c�3 ����7C9�x�u.�������Wt�pS�a4۬e��' �}�ЧmZ�������v���p�d���O�[|e[;!��׍���wY�DP2��CSZ�ֶ���ֱ6[�|�l�+��1���=R��̥v�sg��Fh���|1��}�}��Uc������s�-��r�mq�!̹�.�c��z�(]�Gjnus�ĺ��V1�5fȁs�ڣˇ%��ݳ^�ݛ^�����7᲌�ZyT��<qN��,������U�4��m��˰�d��$�ଌ�]V�m.���[��a)�J�yZ���M�7rk�T���,�E��P��:,�wJgW)H��m�;�ՊK'��wi}�W@��r`n��_�LwRD`%s�}�#@�Gm�b�4���c ���í�Ϻ�D�+Z|�άp�'!��u)�:�	�r�چc����eX;��Vړi��V���.���ۚ�K|n^S�jR}�VM��W��kil/P����)XL gSAǧ1m���j�f�lX�Yu��EG�ޅ�����<��g{�YR�`�`���}�4(5���`�wy��·v�
�ڀI�o{���a>kG̨�K�g����ѭ�gQ�-��=��wB�e�G<�K�13ٵ�Ǌ��s+-�];�=A��J�f�ә�i�j�DͫJӺeb�K9�� �)��es�Rm�v��qJ+;질d���ZsB��6��z>Rp5�g�eJ�B����$􋕅�iC{R�!ҷ��U;7"R��1�8invU�.٫������QQ�U+����Uy�v����
w��s�#{�������Eհ-t��NC�n�G[��-(�<���]w��]ە�7�Rj[K����*t�X�m�O�a���ݴt�w�Z�W��Y�UGMQ�X�%,|��>x�w3r3���m��|�fsm��cc3��@ELX;C[�ܰ}���r��u�+�k<���'0ogT�`��Y4�#���:�Ӊ�w��
]�K� p�o�O���)���:��/�\�Wap���)�K�+_Z-gL�jkf����uuPQ�ڹ�)���龤w^�vY�R��p4� �A��C7V)Kʜ�H��ʉ����Ʀ<�
�h�N�:T�91�	m�K�R���Ks���+��yYƧ|��:� �F3�uH�sN�������h}�7��vR��Oh���H91^M��]e����yGj���Jޘ��Y�PH>Ks^ƥL�K
�W �%��XF��7n��Z,c�B���uu�Dc�BS��C]���`��T�>��a�+���U�s����v���9lR���W����H�H�T%k���+
�B�+*J��R
(���J�T�21*i
�0
��B�ȡXJ��Y���dE ���1��b����)R�`���[CL+`F�RT�LWJ��0P�,�,�*%E��`�m �*(T�"�t�R)i&��X7W1�X�dR�#
�( VKhV
 �s)EE
�haq�ŀ��UdPX��
j�dELeUBc+��H(%A@QKlP����1�EP��Ta*T������`6��[V*��!��DE@RnUX�Z�P�
�c**�+
�a,��"��M51V�D1�C" 
�ʶ�%b��f-��"��*G^�|���ߟ?e�y�p�9���7KДf� x5t��9K�w_fDp䛷D��[�7O4W�l���
�ϖYt<b�S{�k��O*<>�Ө�s��q���,[7%�8�{��p�E�[B�<�]��/;�gV�=i
�L�Vs��c��`�0��R�r��w�ғ��ɉ�<2�<���S�����y3�Ū���8HJ����ܮ�N�6#�3�%,GU�;{�Vwuo���\�
Fl=t������W^��<8�*>fz9Ϧ#��¾�w��� �bba�y���n��8���%�
�R<k[=�-���n�!��&B���-�6����R�����Y�uRh�.5�p.��^g�Ur@h�g�a��q�������i���/���Ki5V��ȋ35�,<_�n�#�^>��(\d�YG�]-#�}����Uq�Ԍ�|�$��벨T՗Lx���y��74����yK7�x, C,�Ga��h��z�sّ�[�T�%t,ž9/Y��,�@ǘ�%���T"��ta�!ls�S�?PD���W�#���N��+&��+��p�/������R�8F	�46Q*���t x�"f�%���|ʷ�>�u�9���"$��׽3���5W2������Ӏ�9�u���� Y+�K��=����2�~�%bu�"�u���jG�#4�kQ�u������ݗ��wn���H�Pс�"�n�&�<����o]�5s�;z�|��*�P��i���g�a�B�v^Z��FJ�j�XxkħO,k��NK�ݽ�w�X-��3��юv��Rx�G�X)���B��e@<!����h�����^E)��Lpĸyg҉��<���2����8o1ݣ���V����I���yj�Hbxi��eD�qu8}ѓ��V�4:��ט�v���ZgW`t�����"-���,^�Gn����H���u�+�xCf�
��֟�r� �.=#�:���n_���%�m�#<cBy΀�]B��}��qY;hG�l�Yꦻ���J��zH���[��a�w�8�f�W_4<e�����CJ���V��Ԕ�ʫ�_K�Pzb���)"�g� �J\��+��n�{2"X�?p��LI��+�u�{��:�$�}�¼�]�b��j�1=͚�g�b�3m٬�Mu�Y��|�>]Y��zG�..#@�p���\l7�5?t�i�Y��,P����Mz0nN��7e�,���B+14�%�=̕������<}CW�qc�5�"�qs�l7A��#f��+���q5��V�[,�T��H�!�6�Md�|6pet�:\���t5�x31�{C�����fbZ�_`���H,EX�գ8.#KI����i�?�������^?5<�
�x�9�X<'�l3�!�W<I�v6��t5�^ٲW*��#,p�|k�߳kl��u�t/�S�HA�}��
���x]<TǞ�q����|7������"K/R�R���1p����F�ҫ�B�|�������_,�L��v⎴Wk@��ss�THB�P����{Jy����q{/�zZ{&͔ԭ|m��+���SX~�5>�������P�.��cςBx�^}u���>�It:���ƒ�yE(��ý��G�}v�*�Ӿ��\ W�4�R�QhG@f6�D�Uv򩐳s2W6V�&\C��Tv��O��'�)�sЍ�X _qDLN�J�L�lk�P����N�v�Z/��"w��מό4�{�[��� �s�	�(��!�#$�J�uAc�k.���L��_��b���z��kċLe����/�ZV}�@X��~=�:�|�x�9!5�-�
��B AǦ�W!1�?����~�X��q���c�8*�
��4[k�Ч�i2��ך<����q���"�ڿ���x�5kZ�촳ayn�&]���}B_SǊ���ȀR���ƽɠ<�WM�T���oz��-ps l����J��S����c���k,[��"���`7�W_nip�ܚ�3����p�+����}�w������gu19�{����J����d�9}ԶRWjM��z}���sl�(R( ����	M\��s�&�W#��Ӆk\>,��Mj* ~o*I��eч���C���oK��M�ĥr<1�RW-sh�	ή�j:�O&%��y`>}Y@�{Le�����wW��(�T���w2S=�"���3����Μ�}���Y,Tl�W_��6����M� �o��y�-�3]g�>�R�Fї�~�V^]�۾��x��Ɣj�0v�q v�o��^��x��2�����1Bn��Rپo��]�`ShМ�'�4�%���WҜՉ�Z�a3�+/��Po�|O�����)�]���]1^�Ubh��LΗ~LP���i�j��^>����������ٽ��{���KDƈ�`݁R��z���}����=�Di0Z���wS2�q�:�_+U&�E�{zm����Q��J:�E�CY���E�UݭZ�1�*�Y���YÔi>��5���u��MwX�WC΃	T�M�z՜���1�:�x�ɀ���;'5xf�H8/�gc0�h�]��è6�����ewd�wN���l]�V�;b��lܣ=oa�~7�k0��1Weu���K ;/4wR��(y�`�w���X�s�C�߅��eW�\c��P	U�E����Jc+$L�{\��^�{7}�W��VkC�PX��d���&>���ǵZ�Y*�Hm�da����C.r���8�4�8ھ�B��:���Q��Xn�����2�op+�lK����<�m�n��W<�����6��K����ΝSu��'moc~^�~�e�0w�/J[Ԧ�%�Ԛ�=���9�^�a��csTƩ��v�)|�εx���W��T�ǖ�'�q�Cf\�v���0���P�f���9SE򇺵?Oh��Z�{��پ�ql��&#m�Nl)����;�^	��P��J��Լp�uq���]����s�eCH�\�-����U�hk6-].4C�inV�w��(Fn�)6�&��k�'���Z��cAT���av����!2Ǵ�S=g��C�[���lf)�T�㪋�ieD+mX�.�^:t�*�P��ΡǁUW@q���{.��'o.�����	׏H��hj���*�9אn�qv�ua5Bov؅2oy���e�w�����9u���[��Ut=�2��K���T�ǹ_N����Y]�>z�v���4k�V�Xj�ݧ<�W;@�ܗi�Y-��P�.j6Q�	����gWy̩�dI|��HF=1,��΄�:\9��c�ׯ����S�{�Vm糩ߤ�}5Cb�䗂��>\��O���`ѱR�����[�3W�=כoU��%+�������:���.[�"y����Ց>���`�]���(��xZ�U��{Y��oU56��h���-4p� �7��\\��S7QZ�eO	v�w�u�Nkq��vi�8Nt���c!CA�\CXDq��G^<�!��o7&^$����c*�daŬdj`�4&;W㏱Y<�p���S�Le&�M����5���Vyx��;��P��[���Y���/Ӯ.H�{�.�͠�mȮ�C����X�-v�!��7+A�~��o.�!���	^�Û�)�N�<��\p��<�mP���$-r8�8�kB�eZ�&���AP�F�Z��d(Qʕz&�C)&u���~�M�T"�݀*�ܳhO{t�t�͎��Ή�=��F{Y��JX驧+��P��͏��9�ʚ�1I��W�'~�c_�c�h�۷WP�J�X��:�".ܙ	�E=瓙���9�J��u���6�:s�U.Ț�|@ m�����6�t���W����r���y���;bJF�5B���l��'�2UR�w5U���|W.=�h�؍��J�-�[�e�Y��)�
�.�QQ)s\msk��mT89�^�yhL�l�N�,��4��9�K�);��!�釜��N��u��=�9�RKxױ�y��C�w����7T{Mׄ���&I.^�vm��;_������}����E��Q�w)���x��I�@Lł�R[o?�w��S���|F�LK�<&*W�t���f`*�4c5�ps7���q�l���:ķ�}ꔻʹϼ&1=�"}i��^��v�r��bņ��j"�	�F5�%�$.t|˔5�}��+��ެ�8�TX����q97r��v�#HY�x���XS=:�W��~o2�'Ȱ�V��z�=M�A:QX�Q��9�w!���|K<��{�-��\��!���ù6&�}ݜ«t���1���M6������em�����v6v�H^u�\�A󼶮�X��3�)<�Yq�jg��f�W#�GC�q� ��P�0���V�!o*�=�m^D��r����q�j�\�3��� 7�T)�˧=&hwRCw�1�o(/�/�N`^l��8�5� 0N�״/��ɚ�z�i����y���mȫ�Ye�x�I���W/=�ߦ;���:�ܛ���j�P�fߓӯ��;g��6�<�#��ݩ+)���v+�;W%!���yʭv���I�*����c�c/��)�{�E�"��rC�Z��E����_�c��r�����p�
�\�Ȭ{ݾ�̫���:�W��s�Z�y��!Wf/��O[S���y�3�\V��=\�{*ˎh��W]����WJ�ȝ�m��[I��=
�>K�ԕ'u��}�5��~�q]�Bͷ���7s^�E��F;b��S����u:<LJ�NS��n�%=U�fu��X�6j<�r�Q��w�3�u��xt� ��$����r%d�P��WΊ��7e�v����ڡ�4��r �+5��G\X4�LL	,Z��W��}w��:���_f��wK�խF�r4�(������<�Wt�S�:Η�>�]�=�]�Z���:p�s�k#uZ��fo$VE/�3�{]��T�k%t"9gK�䗐#a���31w�&�鯅/�3����f�A�6
�ߺ�����%9r%9��:3��3�wL�m:`*��/�KM�W�1TE�^l���͌�L�aF͆3R���s�"n��VPO�n�ᨺ��Ӝۼ���ò�f��/n�p�yN[��ccx8�������r�}Q��U~�$[�Z򚏵.��n뼽|�L�A��&:U�Ն���Wж����ެzLs´���ų���7skz3Sba�[��I�s��n��V��[na���[�λP8����N�e������6���N��1�����O�cl�I*���\�����W7вvX�f��Su�m�N����C7xG�y��]��]/6ѫ����-�D��Cgwi�eIȢ��Wf��OX����y��Y��Rb��8�sX���{��ސ4�����=�ٍ��9���p𝕔���o).ۙ�z��Sfwj���M�����-���8f'.��Rū���+٣�j
�w�uq�0ĬE
�wQ�r�k�3g�Y�l�z���z�\+B`�n���ۅ2��d*�E{!V��=9O^��\�Qټ�ͬI8O:�{y�cb
EW]�Zڈ�t�����0\fc�G��m�����<ި��Q�x�Aw��<av��W�i���*������c�C��󘫹<&mP����kgE�p�����ώ�����f?$s^p,�;Ɔ�b�k��4E�<2��{a9y�7�grk��4�K�&*^����Z���	��^	7��|տ*��*���j�ئ�=�]n'�b���&[͌�Sw�����k�ۋ��4��5��ܶWN�F�=�6:S�R%W���o���Y�t�������t�9�Q�<G=��+�����_o?���Qy@�o��~��$ I?���$��	!I��$�	%�$ I?�B���$ I?�	!I���$��	!I��$�	'�$ I?�B��B���$� �$��	!I���$����$��IO���$�@IO �$��b��L������K� � ���{ϻ �����~�	)%* g�V�Y�ԃL�t*@J�gq`����%���&Í�6֥̒��I��n���`Ik6����k6P����qBr��ضѫ2�M���f�+TM�m l]n�5"%SZ�d'qkRTM�MkmUl]wQ��fmkM-�kNs� ��4i��4     ��JRj�2�b`@�b Њ��
J�Q�     L#C��L� �LL&4��)� ��S@!� ��0 �9�L�����a0CLM0j D�ЌL���T�򞧡<�&�ɩ��}��ҽx�(��H�"I! �?�%HL	�!! �	$��\����?��c���(�l�3�"�!2HH@��'�$�Ip@�E��$@4�����������~�$$ �9�*�R����3:i�������R�o˷�/�*!���?�����^R{���qц���>5ٴ�@R�w��WȠ�݋/.�o�A�L;Z��BKB`&�ne=Xg�DV�p\������ef���ǆ�L�8-�퍧��%X�#�2�7b��WJ]���
_��e���:=�Z��d5����Qp�V��$���	C����ix����uywh-o��hR)� ����±�JT�,��� ����f֛Ä�b`�[V�T�b��P֣�!�wUi��'(�\*�9�����f��*�q2;v�ܐ�)���H�����rV>��V���֡5>U���F՟�,#�����Uxp[yY)_+oq��Y�Ma��M�ͬ�T�#����� �g¶��Íh4_��]�YsJD�N
KbO����kyPVRW�s5-D|S�yV�;u�������U�2�.y�F���m�͐콢����Uj*�x7icd�D���QU���e �)P�v���۠��R��O5�ӑ��Uu2�$�����E��QՎ�U�޶-WKF@�*nV���נP�&̠��f�re�kv4񕚲���;Z�sF��&죈�&��R���]'ɽ���6gWv�i��7j뎐��}A�if�F�U���H7����gL�r�G%���P�һ��h���*�V0b5w��(��ѵ���k����� �y��T��5�����V�)�ҩ]��{����D�`��T)Ղ-=�2��iSI����Bӏ%���X])�	�X���*x��.`���Z�b�^�,�Y�f��j����ۦ��!RS��2����:�h���F�Q�$�0��,�v�6��j���Д��93*Ts@#B�ա��p�SІ[i�֫��CE�j�(�����α���oei��Ƶ�oS��!�/����}D�7��`Б,��[T�*�]�'���ަ���g�                                                     5��)���Q�w���mJ;sG_-�AtF�Ji̋�9���u����w�G�<[��w3�/�P�M�!In��T:�ݷ#;�*�AMKK��������ȑ�.�iN�nN4J���{$��Sq�� ��	]�5I�qb���7��pv!Z�D��{ǟ�0f�.n�5��1��o����eG�ʾ��Q�\���sK�s�Q^:�;p����V�o]p:X��+��6	3U�Y��5W�\�l3Cl��MT���TٜxC/���D�@�D]�ݯ��McH����FK3�����R���BeZX.&����(�nbOXC�	C��jM�ѭ�Q8]`D�3�l4�S��&�����e4���ĻW@�*법ݕaL̕+ed�|8<e���ˬ��V��fE�S�����a]��j�;-�xx��30��Ozq��]��"���Șo
#�Tp u�����{Y[r��d�vj4����`p^�gh��ԝ^>-˛����̵��|���G�7fl��
� =�$5�9����Jv淲�]��b�&R��MR>�9`%m�=�M�[�EIjin_g ������f
��zT 0�S�F�	>i�K̭��3:p�F�q�(R�2��             4`��"˛F	���12���i���vH�	Bʙ���Iyp�+���L�yj4!�R�� ��M��}.���vWE<`�\wv�52_B%���R�Ts@��r*�t8������t�����⨳5ˤSX�2g�0��`�d:��,�әo'l�Y؞���3iW\�щ��4Q�'M�s�&_B_H��!F�N)	��K@� �T�#&'A     �'��/տw�?F������?��y��7�=~ ����$���=����\	! �A�<{���^�|���3w�{7��y�꠵A$��!]j�����r�����z���V�N��XE�ho4�����ɳh�cn� /#w)Wl�!ѓA-���ܶ��r�1�:���td���r½�k����p|��H�,p�z7�j���0�l�hhfJ�V�A{\ T-��n�R��0![uA�,�:9��M�Vk��aQVZ��ݐ'Q�����"�fA���钦���&���Zw��yfOB��CWG��e��u���۲���˽<�/F]p��}.� �Xr�E����R�n!RʜA�73B��*��2�vՊ��5kk�Z��t
��l�*�� Ԯ�.Yg�it��A�IFsXq��t[n�jt�.�� Ih�!em�f(o�Z��V D��Y��7L�Ғ1�lTq�.r��Y�j�v(�P~Ǉqe�Fq�}�曓2�q\o`��q�U���/)���Ⱦ�#�b���jT�-�n���t0�iJ�p�7i�옻�V���~rtO���*޳o�us����%]����6���k�����S�F��i�Ѥ�"��Y����k�j�RS�w�j��n���jE{;6h�Y�<���Q� �ɘovk�8kT�+2����Y����Nl�U'`�!��Ϟ�s���M�L�t;�"����բ
D�*��\���U���̶ʺ;B�r���������S���&��*3���Z5�M��݇d[�kA����������k�z):��ؘ:��Mb�ǩ�-�-�e �wB\!���������G�hA#J_U�� �����͎u��}�,q{cR62��Q�Tj1�rb�U�"�Iq�U���ڏ�ɖ%�|�Z]�V����̕�'D��*�� ��ة"�<CX�X����ۤ��9u7˼!�Q9�OT!! A�� w%�=��x�<R2;;/����   VV��H�F����Dd9
K(Ta�'B�q��8ȗ�9�a��	�pp3	��� (�f�'$�J�/�PJ�H��5n�� �E�4�+����������ë�)%6��8�6���4`�֚QT�����QJ��Z��I��x�nMd��cuBa)��)�YiuCT(\A�j�e���**J������o*�Xi'GƩϋ����z�]��߾����~�k�?�4�s���Ɠ�Ӗ,�i;� m�a��&k�����e8�&��g����IZhXgtKK3,��ˮ��{ɱ���e;E�IǙ뛼��m�n��L�Z��I����wOxۧ�e�>�+�ڳ������K�|��P����{s���lq�4P���U+(�� ��>9ra��b�U-��zu�0�0����ޯ02�v閜N]�l�;gN�u��9��Ftí��6�@�:��v����KB��6۔�3rRq2�3���je�-%���9��,1�FET)�V!!���?�ۙ�օ3�Fkw�`8��N$7���5�M;N�)']�l㗴{��4�4�W��e8��L��֫8)7�X�E�N��4�!L;y�8�N��k3i�
f��e���e�!��dR�b�f�h�]~��uZ�WYo��헖���Nu�u�/e�S�q�@�n��L2q��Kz��l�6��%r�\;NW.m��%!f(����Ci�-&��
�L�ӄ�a�-��Rq03��p��{�0���eL!}V�2�%!������{�Â��*�t�fG�y�E�5m�)7�8�I2��Q�7:�+��t71߲2�d u��,�C�:~�C]��|�+��V2N�R����Yj�1_�ri�d��+@C�PӠ�v�������9`�mn�62�eazz��D6oD3=��8vAm��R��
�t,�3}[��~7Ph��Fs�`{n{U���J;���fz�����֕�fc��%}���?���ۋ�ܲy�F+M->��eҧ��~��OȜ��_���-��'`��q��眲/��k]^� #i��o�3���xT��3�(����Kʚ��&{�c�mgm���N)�j����o~n��I���K�[�.S��e��T����&\s��ǝJ*L?70�)9+{��������y�9ʘs#v���"�U��y��1�ag�*�ȡ�B��yٻ�׬�Gމ���4*���ޣt�{j�o<-`�������'��}I�����m:�E�yu����Οr�wsL�*�fҺa� L��V鎬�b��1�T4�Ssw�E�Yp��wW8� Cy��)�X�:��dc��h�r�ذV,��S*��w���U������   ����Dej5'[��s*s-ǐ�h�[j&��$��<��9��k7dfF2�L���A��4�Va���B��Z|��5qL�"ԁ�*)'��L������Yw�Y���
n���Giv5M4-5Z��x�R�R�]L.�%��8�������u�m����N�[s��}�i̚�~iO�zvvZ9����Y�>�^����t�_¢۽\�?�;�W���bΫx�]ʢA��/�*��[�Gǽ���+{F�'��\q�]ڿ�~�w]�o�P�Wz��������]�8j��ZJ���.U�G//�1_��1V�P7�����W�e<�����f֎7�u�p�~1j#�v�|�h��oy�͸����H:��3ا���7/x��QN-������*�Ō���q�t��y�����0�J���<��փ[�W�<<�G�`�ʴƕ�[�dMi�������1�,�3�xo�E�v,y!�r�֬^V-ÿD�_���#gMx�^ӂ��١�A���Z�4ǈ�tq�~��=*$1����`&q2E�V��ϰ̬<��O�>7��)p�
W-��hP�qE�����c> j���;����rI���#�tz$\[ֻ@�Jd�w����zM)RC�ջL�T���(GKʺ�eyz���R9��v�xʣiAV��H�	᪪1]��m������@Ү��FS]��c1k��������U�9׃kh́�����5o��]x|��]ʑs�~e��q�k0�~�ǭTi~��w#�����RT�IY\41�#Y�pᵭ�3�C>BrҪ	{A'�F��TC���n��G�[T����"��{��^+II�OYD-��ޭ/E﫟?f�Io�����]u��x�\�v{��Tn�O�oȚq�o6 (F�����������4�6��w�cX�����[�e��և��g9���� 7�<d�����~��4��_�̹�YW���nk@�R�]!^�%�F��405�_X�ϸ;f�F��S�M{���L�m<W�J�z����;5+��%v���^Ǖr��^��֎�[�ۨ��   ��.4Т��>i��d,��C���P7+8����}=Π-P���p�;�>�����$@2K�0��FU:�����SN�4e��U�q��?u�{��e�5�|U6��U���K�ʸQMT�����U�-�ն%7e���EQf<�+�s���,A�ULE#-�i4��9sm<�F�m�T�T�hwʌM�3y�L�ḍBU�7�=3k����eyQ7U�Ͼt��(	��s�����Fl���.F�e�p�/�z������KƏb��4�qq~���n/H��F��	��"�����}1�J����Lnҿ9��_<u�{=Yj�ku�ߤ�.��P�����ĿiM�HL������)�d��x��YbIU�I�û��k��]6~0,��Y����vd&��D+������5J���&d[E�Վv��J�=�'Wc�h !w|λK�w֗�iv�mj.)�v�vpX��{}�4���i��6�O%��'�uɓ8�r�D�Ҹwe
�]�*���3qe�E	����d���lD��X��	�0z����ҿ����BOߊ��	O�V[k1�b_��R�[���uAc�Q�۬��P��rF���Π�`5�P'��3���	�y]���z�	���Mȼ�n�y@��2�	��c��ң�Z��پF�z�6��v��q9��xK�M��׷Kƙ�<���#oZ�T�_��X���/�n����^����j��<J�;��ɚ�;�_ܓ�6C29�#��%�o4��G�s��s)n�Ʋ����|���]��Wt<�����o�ݳ��QmzS�8sh�W�����D�,�^'G\�Nl6D�u�؋��U��`����3g��)�o$7�mI�2-k<gj��>�Ә��˦٭o}W��[�!��9�YR=���ř����Q�B�����e���=��W�s������(��p|��X��~��*��⸍�;&vk2+rg�ydn���3~�4��$�����'u��{�gq5cY�ˉ��v�ji��Ý���+Fێ�֍<*aC7��Y{Q4�ݵ��
h��m�\$��(�ԋ���G���5=$7Cd�ؗp  ՘M�C���MVY��ͥ�NK�pĴ��@z�/�!�b!�V�R�	�U�a�$�2���t�������I&�QD\nG'�Uv���T�髡heRSU��qs(��3uTv�n���bW.�TJDb�I�D�	4M�Q&��J¡I�qp|�"�� ��D��������?����|��|+*�����[h�(���&�Տ{���,�����Y���`-9���c��4Ë_�0yM��"���c�_,�3j����_333U���u�ĺ�(./+�L�5�-#Qs���y�<���t�/&/	�7W�3����1r��uN��:~|d�f�޻O�g-�5�3y�-��g騾��Q��f���?���듣Y���d��W0c�nΥ%x�;1QS��u4�O�������56v�C�4�����n�_3{�w��y�e/?	N��Em�_ֿI�yc��[F�;��>tt���yC���v<GT�N8�t=֐0���-�=N�������u�y��]��o�J��Ŏ�fEY���
y��~D^�)��g{�Q�H�������^Cn#�=��p��L�kw�6��Z�����#�y��6fy�R��q���r�J%�<�5���������=�r��G�oNI\109'���i_�����==Ɲ�g:����Ok+t 7��ՙ{z�W_�ڕ*n?�~ڟ��x�F��G*g���6�_���0���k܀&+���\��Vg�P�M�K�O�׷;{����U_UK���5�A���Ibpb��A6ON>�f��c��`n�����aO�;�dln���	Z7ƞ������3��D>�V��b 5}���9�t��ׯ�P��/p+v�(ػS�ā�o������sZ�CN�Ш�^�����W^f�Q�=z#'�3
{"�M)�ȅ�4F�[ݿ�����2�~U����W��aM����Y��\疧���I8��L$�RO깂K`t��!��8$	Lo>_x̐�L I8��U$:a!l���g��@a%���I��CI	��0 i$� �v�CL��$3ʄ�xްI2II$����B�����tu���~��u�j�7��a���cova�4oP��9�qE���0S&����9�%ͺݼw��N9Ka�yjA1*ŽҔ��s�7ë��yx��5�Vb���ua��n��[t@��$�I$�of��ƋBj&��R�
A�a�(���Kz�RZ���޻��rb@f^LrᓤƂ'�xzD�6Uw:��ȔQw&���-�  -��S�T;���CT闈v��U�PFA^��U����QN1R�,������0�.���S)%��c�Lc � R����m���N��j��b�,�V!��l���{�)��$�L��s�o��!�Hq 0���e��	�Z�$��(��L!0�<0��B�HHv���� ��hJHHS$�9X/���w�7�	�t���0�ԴL��9Uٛ�ީ�<ԕadK�ce_<�W�  ��y��r��M����p����s;aN��\3#�<�]Z�f2^�<!����Û�z�01�:��f��$Z��/�����o�k��ia�/�u����[��������J
�+~fC���a�=̵Y��y�r���'bd��v{{tϟ�
�$����H@%���ٕ��ʙ��u����%?<Ǟ��=:�����x7^0yV+��El�k"���c����Ė�ӜU4=̗�#Pj�33U�}�������K��V���P�5%?6̄٧l�æ�&P8��]g�R<J��Ԍ1�-�Z]�w��N �T��z'Pw�.���!#��6e��(�v�"}�Nh�Uߗ�|�c}���dy��P��83W���Q�1�U(�"����pfv��~��c��^Unt˭�� �#�w{_���@�-���:�o�/�V�j���ֲZ}:�Ǘ��D4@�
��j�+C�K���G��$n�Ǫ�����Wa�s���Sg�s�]�!�K7�J�o'�Gl�6���Tkа���Z|��&�Gظk�Ǽ���%��k�{���e6���cTOK���[&X��;{����o͙�k���<��)�L�?ՑQ�o����X���yL�m�Mm%��Dp�&{7|�[[:��;��i�Z�b�_������i���~���a�o�	�qW.g�;�V�/��5�ғ�~>�a�ui:t�(�9������*�g�����o��s^�P�Jk��yhC	�4�/S�'��j<��i�y��
�}��g�Wj��}a}�d��C���e�ܩN�$d�eT��d[�>l�U�,�,@  5p�ç*Cky"���QA��^[�	�b���')u]��-�(I��Mu�drؚ�؀E�{�(䑴Uu$���RSkXnWr��bKM ��*��iM!T��Նq@�q�N��+������IH���ZUj���)HR)5ui�����w�xv������/���2�c}���S�c,������Ǩgq��r��n*�U�^_Oy^�|�U��Ւ�5�s�g�'9�j/J�"�o�Uz�؀qO�����3�V���EA�W|��� 8o|T���	����Q��8���@�M0����ؤcΏ�S^q���C:X�sj��@/�v�e)��姱�B�K0����,]��4=��/x }��^g~΂�l&&e��6�j����YN9�oS�l\Ϣ�'���1�zX�lk�����?}u�'��CsQ�	��pXH�����"���W(aGm\:�k�k�[�r����<��ڭ��0e���՘�N[�ev `���?�<�M7�"[֮5�ֺH�/+����kn��6u���,���>��l�yr�
�����e���ؘ�����qΒ}Ws߾���}���g����_��_�]f);E���tZ�5�檄�ۣ�kE/�q���B���OzW������S��Q�bp9$��ZO����(�q�����,������w�J�WE�r�\�M#Lp8W��{�i�GD��Wn�-z���tSu��bK[�ɸ���ԥ^����(���;+��;F�_�b����f� ���Z:�~(�K�[1␭��ժ���QֆR��d�t6��guH��E~bg:�j#�G�_J�p��~�{�Xݠ[w���	U��]�q��?Ӱ�~�|��W�1�x�f��b��f��g�!�G$�����N3� ��h}�]���JZ}�jh�u��11�J�^�f!��ԭl?4 �x<�k^oҍY����^˰)n�*�m�{�^�A�	�4����t9�����´�c`ђVXkV�Ω�j�ud�[x�h;C-��{(o\UFn���)WJ��&�$   E暪n�k����I�nsʳnr)����;��)���ec$l����Y��L}Ӝ����J���rH�*��v��W-A\�yr�Ÿ%�  ��=�7����鴡	Qv�L�7Tm0�P)�Ǉ�;���ݳf|��{V�N�Xe�E��vJ��.�ng������Z�Ӱ�&���b�5nU��K��Q��eӱ��B�&g��l�w�} �"���쫭C)>FV���.7�?��9�6�D���Rv��KU�[Mc_�l&��lz�;b7�mݢfY��R����%1Q����e�ێUe�jg����7���@h�Ӿ��b�Cۻq,70�Ry��Yx=؅
Z�恸�_�Z�\��Og�ȋ�/�����a��Zv��oJ��0��怜"8�I>�G���x�yȃf�:H^d�����WmN\P��E�\Ѵ�x*��x��~"��'��<�<4�ʖ<C�RxT�+p]gs,j�Ӑ�#�}Uĭ���d��
��)l�,_=��?N��N��M8ó�L����s�g�=�ʯw|���U�᥇��'c�EK�����������:#jMm� �^�|cR�#�+嗹�ߜ������^t�-��j��֊�:q��d0w�p��a~n8�Q?]����Lw�~�Ԝ(��Л별ӹ�V#=��]h�g��Q^��1�dT�~*y�?u�I���:y}����q�����������2�����ܔ�_��� ���p�]א;�F���E{�B��\=��^��{el��;01=�����YC	�����"8�G>�$?��c�S˭#�`�0*���*yO�̘)Uߩϲ��(�����{a��DӬ���vҌce0�{kn-2���d�G��1�m�o���8��U���j�,$\��ێp��B�Vˬ11��{95F�:o��}\�(�IW�Ε�)�=��O�?,�6���@1�v�V�jZ��R��r�~K_4s��i��7�3����:t˔�k�h�@�:�޸f-T���5��Œ�����@�
���q�`�wts�y��˵4��J-��{s]]�  �B�s96T�s��	ȉ�n���NI50%�k�\���M���X������S���N��ԕy��RIe>Ej�e�1�����R��8 �<_%öWu�Z�(v�vR�EM�б�b��)�.�Ub���mviwvy�����\n!_����N�h����b�0#3$��1���OY�E�x�zS� {P��N��NSV<.��N�'�pf�CSځ�;�Q�c��b8�}UUD�D�|o�=�kב��i`X����گV8��or��KR��{	�t=mf,���<�	��7]�TP3{�j������s��)�nU�*��h��ն�����[C ���[B�w[젖�^ɏ�%��h!���A�V�
0�����w�q Ȏ9�Ϫ�����J��Z[�M}���5�C��/�Jibx�谼Ǯ�S�<���1/5i�eT4�&�f���sF��Qxa+}r�VH�,xsi?$�?�~�����ݟW�Ȫ������1�0b��]���۷%i+G�(�dv�vc�����Y��%���]�Y��o�e�81渓q7��_�~s�e}[�41�V{V���
b�k����\�4װ���O"��Ymz}3�n*U7���?#Li��]E�������#�7�ٗ��'Gse�GP���uV�g��I�u��+@\�-�/�+#���%-z%�sֶ�Tr�1��$�{֫�ė�.�9$�7����w{��4rn~�~������^����}�3z���+�\�G��:d܆,�2r�WA��V��c1��V��lʖ�"p��,@P���^_�W�Yh��%Ю���d�ь��&<C�cf��~��4�c�)�E<��Ď��h��L�:�����
��1�on�W�f̾�d�^���i�����{����{��Qֽ��x�m�ta�I�����aW��ǸN���{w�P���&e��(�����6���3�����Q�$����:�ڎ+v�ή&���ܩ�NH�yG��;��HJ���&J�����
�]�f0���U0n�q����.sav?q&j�   FVhꅪ�C�\n,�0*x$���$冯�w-I��}���+�u)�P��17O�M�����ζ̒H�J����ޜ���#9#T`��TƻKS�C;����c�$���/I3uUI�OB;�c�R�pU��������&�H�.�	�f����>��c��絮%��Y������=�|ǀ鴐��СW�/����~���5�U֭T�0d�����{w3��{�ܩ}ϕ�x�hAs��U9�Y����v��ӌ�ں�K�%��]��:�~��9Yiuv����^�O�e��k�+9uX�=;�%�_)�*�[���ެ���;_}�)r�}�^�إq��C��Ζ`y*[^�Va�ttj;{�_��&�}��E���>�K|�*�:̯u�Wj���76H�"8�G����N�ir��6$>�n�Q�+}*x������A���fj:L�4�,`�^�V=f
�J�h������L�.�#O�j	���7����u!�?#b�t���q��~��\wQ�.z�~��ȦM��kk�v��	jē_��-��;N��s��d�n�k�F�����x�}/m|K���_8a��m{Z�z`�צ{S[ds�X�KY��^5%������a�z�1�D���m,��4��I-Y|�P7�-�~*�S������, =�3ti?ml�Gv�������Z	�m���̈́�w!p	
SF�}*h���22����#��m3E�9w?DlG��L���/��#ފ��X��6�/9U���T��ӌ=�<�x��������f֖��{sx�Y��U ������r��?Z�efG�5׈P�t�L��V�p��9W3�����SMv���/=�zs}ͅ�i
O��>�Iy���-�f�g/�[�S��}�����Dן0�`��_z�-��
ggz�=~��j�{T"��U��c��p�>g�⇯W_S�u\����=7Q�y_c�cx�͢�����b�j;�s��:u�L�u�p��(�&G[����g8d\��S�
V]�:�t�)W[�s��SbɇI��g�h   UY[�*"�6��Y��%DN+�Ci�.�n��\��đ����k��]���r'd ���-��6��0�dq���ZAD\쐨$s��n�
N��M&l�L�Ib���A�Im�tQ;L2�X��#��;i���

�����UQ�ˁEUb��ؙ�D���s���6�"
��Z��1*�ҕ�Y.���m6�Sl���u���p�4�79�V�஛^�-]����L�~u[���h5�t�K�6�R�5-���7��K�s�]ƣ�G�}���3̴�g^j2#�t��ďe%ynjYx3|�O0��C�+�B�_�x��Z{�h�/נG��.�}Vh�盨u0�{��{=6�Xs�I��'�_���LGT�b�_��5���ޒ��F���� u���;���@S�Vl��"�x���� �]s32��C{�'��E�$P�}-��>���6Iy����w��˫6�Z��S�h�Ź��\]ub�	�n���e xߎm��՘�aAqF��'�nS���3�*,):gx�+l�0��ˣ�\��v�$�i��1ίV�<I��eÎ�
�y��4�Ht��ӽ��;Nn�
�U��hC.S�����f��Fm6�@��ل��E�풞�<�W}�7�W����5tRz��� �3]���0�w�2���ba�a<=b�ꡚ�X�q�AfS�N�<w{H,�%���i�4�ȥ0�X�]����:N!�N�G}��;L!�T�˶Z���[8�0�M�/�g2`hf�ImwE]�p�*K�L%V]b��{/����v���	2G�����3���i�0�%�;��iHe�g�T���	�2�ni��wWwH]Q��N������\x�RӶ'g��,�0vfO��v��v�K9;Ad�Tu�dzG����/;i�ķ|���U�ۄ��Zq)��myx�)d���&�����D�rI��I��w�,�v�Qi��x��Fxah��xƓ���G;�Ghe0�i�i%�Y�a�p������2i�i�0��]�R�0��m�Q��m:fMԔ�C)��\�����;u��{�'����g{���X��z�#"r֤o���x��S�=Ppo���1����Rw��a�8�10ö��6�нI�)�3I�í���X���3)�u�N<I�R�Ii���N�}T�`e���R<�6j��awX��n�e�m��Z�X�d�6��5�v�L��;�o��A��#��_�F�2����$��a�V��m43I��I�)3�gZ�,%3��s]�zY�G7fX�L���;���e�Vh���4�0)�K�v󕌺���Kfj5i����Pi!uC:�`ᖝ�ӌ�i�C�|������)�UU~�4HH@-���		����D�����.��UFV
����~�����i؝5���7�E��0�C���`~|*y3�L�eI]�~��e����/��>�ә�����Bx��_'���W��}�=�2�S�&���z������.�~�R9,<vfo;��RBB�D����^X�=���nOt���0I� �����aRY�<����h�O��'П�J?����l>��|�Ϸ�|������s��������1Rx�/��d�}��5>�F���גWD��l���
���3��4?O�Ǖ珕ϻQ5W�~���d���/hc��^��#s�~$$ !�r���+>u�J��_�M���<�����)�i!^�_8zL�a�)����D_��T�W�C��C>^$�����>g�d���_Kw�M�^�eI	~�S����Xy��O���z���1G�OV�*�rP7	�
���#^����zI��>���<������~�l��"BB�h�{��?��yf���~�Q��dF}�'�����	������?��ʊjOe��^X��ᐢC�̟SG�� �U��\���?��<�� H2Q2ld����^��:�i*	���3;%�֨�-�T:ٜ���0��u,>>��>�I=��>�BBY���2�|�`{�~�����x;�@#����OBY!�����}��������/������_��y�*��{���Ϭ�}E�ITP������HH@*O�!��y,�ߤ?C�O�/˸z��=Y�O��5�lf��~?<��o��^i3�I��x�3�����_����,���3��y$$ �����o��׿��>�
������'�g��u^�P~P̓��=iBH@?�$�[���@���g��z����T���{��>�A<�o�D��c�Rp`gw��|��jb,'�	���|�yBx����rE8P��'~