BZh91AY&SY.���ߔpy����߰����  a6~}�R    D�   U   ��E"���    @              }�mT�kfm�J�Y���(���j�	 �uN ��Q$��I� 5���:������G}�o\{��}z��T<�ל�ocҚ緽�����/#�>֚=-��<�ޡ׳��;h����|�5��n}���#}�t�A٢�w|���_[k&�/���S��@ql�AZ� }���V� �R����>��{�m o��/����ǽ�>{w,{mۼ�o||��	=ڋ�w��C�:�A��{ʾƹ������Qo���9����}��vW{������>�}���l>��w�ٚ<����*�������}��i��v{�{��S��.��l{�_l��6����oX�o�(oy}�]dA��y�l��#�ζ.Ý��Wp���7m�kֹ��������kAKF�8}����N����l�wz���|��[}ؗ��{��hp�^V��x<z�[��_z 9�J`���t�n�;ޢ\=��=�Y��'�n�^�|/��I}����`�� ��+��m��:��C�;�K{kׇ������yw�:n��ٱ��������k�� �z�k��U�t�E�G}��{�׮�Ǟת7�{׻�}�;�=���      Q@ 
         D P 	T�oT�R�3@b4` LM4���DIJ��h144h144��MFFL4�)HMU#FML���@ �%=@�J�0 �  dh � H@M��1Lj`SĆ��M6�OS�QB�UI�р5=hр4��	�>��ad�I��D�}I�?j{s�Q&�E@�h��?ͨ��!�$��
D�T�����(����(��1�R׷�1��`����������¾40?�?P@�ª(��S�0�I%
�A�n
* `�=����$�I>QLZ�DQ�C���+����~o�=�/�Z2_�_�W��-�E>�����H��WK0~�c����el�ߢ&ەB&;����>��JD�R�8��a��J���ɺ��ܮ�4�Ra���5l���R�-�Nc+��c���,{>r'i�d��nI��-�%�A6��ݲ�~G*�̕�9�:ΗS�$�d��������<;z���%�D��)����F������yL�R��t8Hl�A*�j�~Z����_W��GsBi�rK3\/Q̕��_f$��.J܃��gȏ�9&Ƣp�ʮ���t֣;T�;$L����'N2�6�%l܈�����U]j��ܐr%���U8L���u�~��s$�o�rA�ӽ��#�+fJ���9��k�|��n&���nV$�Ăex/T�~�OT��Va�����%bKbK�%�J��IOu-�IH	C�jIbIy$�R~½��i�y,~)����}Oi�>��M�I�%NI��ѸQ�.���jM�'4��t�
���#�f��N�a�@|�P���k�Њs�	��c2/�!�!�!���%��Ԝ�i���5߰��o�3��[��9��6����i�9G(�E��t�u3g��M�vI��Q�:�0铲}�n��$�#�Y�8�b=4K'���$��,ݖk�6���u.����7���w"N|�D�#l�?#"s��D��gM��\4h��%m�B`���)Խ}���'�(�"6�l��:&�5�(��0j"u�DNo�4:ԭw����C.l�ג��W��el����H��D�G�k+�����_#�(��5rW���|�H�"#ܕ��jV��R�8�R_Ȼ����D�e"o���u�"=�[ �6Q�$�M�Dr%ϧ��R�-Ԥ���#˕���+�粑/�+bi�M��e�H�=���W0~NQ�ޥ|�͔P��m�H��RX�����H��R'�E�Xpo��~{)��N	o%tM9)8j�_WΥ"[�H��WK1�a�KϜ�ҙe����$�W$D�ɷ*�'vʡ��U.J̙�:�л�9&�	�Hk�y8#��N�UӦ���454\����}"98^D��VO�$6H �粒�K�U���UL�#��4�R,�3\/Q̕��J/�d�V����G"?_C�P�؜yU�1�W���$L����'N2������ȍN�'D��T��+��d�G>��Raۈ��Y�N챹�49 �ӽ��'49r�&^D�9	��k�A7�����?(�]H-H&W�ړ�I���ҽ��0���,ʒ�$=	�I{�{R��O�I�����bAy$��<½��R�y,l��2MGQ����9��ܚ���R�N�)g>��esR�$��u�<��㪭��j]�����$I��	C�H�>4�o=Ҽ�M��A1BBy��^J�D�ϻ���Q9%�ѣTU�"]$�&b"�'>�Βl�'0��'M��$M�',�N�',ۄ�Y0I���h�E��*$H��N�bN�
xKѨk�	�1�g~9񿬄i7�D�M��H��>��u'S)&"lu�0���&��M�7���7�R&h�(���^��	̄��L��̒a(�d�gH�D�d�Hu�q9L��'N钎﬜Ý�3�[&C�.�� FO�A;%rO�dԟ]���5[%!hu!�ɢ�(�V�b]�L�'J/����:%&}�D~���Na"B�N"u4&i����kBh�$N|�D��`�L[&0��~N��w����i8=6vģ��9����'G�������0�ݓ�8r�M'G�%	�I�tO�3D���"s�7@�o	G>l�%"wIǐ��ĘlNM�d"$�h��Ú�bU�D�G�\H��$DS��h����}c��6O��"X�3�Q7�>Å0�!8	Bj�"w�d��p�8�8l�|��l��H�\H�JNW��5M�&a����9Ia:X��Ç3��F��$A:�#0�,~Б�DD�4A�J���M�D�L�NɣNA����G�t�)5��>la�8HB�h�H�6t�ț'N�6	�ɖlN��B����7'Q:��'Nh���5ӢRY��Dd;^��=�DX�`�L5SGnY���r%j�Q�sd6#Q�����$�\���M�	��E�J��$D�f�lr|�f�;f��GG���A;�?t�nږJ�Zbelٝ4(p%��O��#hz�)<��xM6�I��v�����zl�C��+�'�B}���K�4x��G�Gv��Q�1�,��h�\�l��UQ�wE�g�O"}�����M��}N��Q�����N?T�t�L��ڜ&D�aD,�tf�#�TG�!ͥ'i�_njk�&����}�5>Gr	fT��Âf56Cra��DG��܋U4YF��RĢq��,K8Y�A�E�D���"J*��ܩGJ�O�n�"hYfTؘ;�,y>Dd�u��*&��6,�8]�L�P�e��#����j&Y-J���f	n�Qb3�r�)$�I�+L��$N�'Mϑ]D���4axlD�Z� ���m�֦�|�؈��Q:jڔA��G�QO*P�ʈ��Sd}eT�vDwʚ�*"vn��7>Dyu4".TD֚�'z���'n���W����D�jQO�9B&�h�B3�;��ɑ)�V�E�۩�\GwQ;�TA�Lj,��TL���57*N���ܲ�f���iBV��ML���YZ�Th���E�R�+Q6�M��Q2%&B��j�|�������D��4h�eQѲN�3U�'�u(~�j'r'E��9Sdފl��h����SF�%�u4�,����})��SBWZ�'m��h�u4J���>u>u>G%u4^M�T�T2P�r�:Wu�������������o�6^�V��^�k�K'd���Wq��9��
*[���\�.y��#'�~�_sR�$�K�'*�r��G��y��2�I����h�>Ə����<�t�\����Z�s�����ǯ$_���=ϊG���u���}�H�"��Y,�4U���j���_���j����RT"`�:C�N�kUNN����}����gG�zO7��(�;�ac�}�S���^��.�CǨ�M����{��+��9�B'�sS}��}
��7��sc��j$�љQԋR�d�S���#��wKZVt��>�:p��+0�q4|NaY��4z=���^'u�r�=���:�NH��VM�٩5P�K�ʩC��UF��&5+'.�&�r��Θl�Z��QĒ�]Mvnj�Ȣ �
�!�aj��>����ZJ8�Gq0�䈝�$��6<��Y\,��M�ܯ�Ȕ[�L��9+�~D�\�M�2",Hw�ԭ	n�"qԤEԮV�${)}et����J�a���4ܤN��J8nO��&�R'E�Xpo��~z�OK�gN����!�Bɘ����4X�U�µ�HG�+i���O��zH�<�#��{���t$�0�r�����Ǵ�u�!*�(EVWg�w�_v�Tx.g�xn��ъ���������edɌ9^5�ђj�N�Iu���)�f��N��8iՐ�%�r<Y%d*Z���U��X�CuD���#���}����y3���'V��L��_��a�#{fN�Y���1����=�M���WFH���)�%��,��(��W�^^����^�h&a�[u�k1�F��l��l�B���X�B�:��R?ld�\Ai�E��=0bgB-�<�x�4j�R���f�M�H�QT�ʵ�{���?�K0��}���{��D8KB�PH�c��Q�i��%��pb$���z�^�uӧ���|���E�X��	V��e:Sl����a/k�zz��i%�Qм��=�4Ô�Y�'YH���JE��t��L�;R��]+����R5x�zi�ϋ$�I��f�F%�a�5���I$�D���ѻ۝�(�l�ѩN�ۧH��zI&���*�U����(�$Û�3ҷƲ���L��ƺ�,�L(Ӳ��vW6�jef8U��ݯp�la������L:]H6�'�^"��[��n��o�М�Qw\�<p,D�MǜG�E�\ZQ�������aӲ��"��*��>8G[N��׏PZOMBN�?}�~7����;�������d�Tg�T�k��T�V���W4I$�w�enVַJ9s	��6���$�����{=�8�p�C��N7�֕#��^�A��m��cV�z�T��)"�u�������7j�_[`��M�'NS4�{U�x�X]'t�m�d��!,����Yڎ-��}��g��rYL�Vg�):w�r��0}����H��s�|�;Q���xϯ��^���Ř�l2����̕�h�x��Y��0�۹����㻌溭$��UC�gs3�u�[fg��g��GI$�p����K_{n�G�_YT����s31�5g/\��ɂfzsl���xr�y��,M��,+��Q�۠ۅ��hb�d�@��Ay�3�Jw���_Yƫ>$�+4Ʋ�eX*�S�d������wΛ�Zj�Ŷef�q�\�PZ+��
�&nf�3Wz�4�Td���7q�8�N�{��'�?}�����|��[ܹ����`��z{�,޼#AG�cÌ��i�I�i�(j8Z��R�^�)�K��݃�aHw�%��?��;�j��{���ڊ4h�OuDne�:h�Ay�r��Y��޵��Q�{�|+u�V��Hc��:�ER��ٖ�cg�ٚ����Y4�C(D����̙\���^
�Q��*ğ��)�
m�� ]�\~�.�wc-��Y"�U�R��Va|yޅ�x��`��Aw��N�W͋����QX!�y�mm�������^�v�v�l�Yk�1�#��&�	�s���ޯ%�HgN��wph�{4��h�va����YLX�ǌ��宊�zoI�{�v6Y�wZ�-�#i���I���G��ra��9�C#s^�n��mt�k�~y�a#���x��¾�����S�u
��r��.����O���K��9QcJ���N���0bx3wپ{���}g�(�h�9D�?�qd'�^!�.c{f�e١��贮f���-�k������m��������e��VŬ>w:a�������r	2eg�p�o���p�N����P=A���ɤ-���K�F����ԁ³wl.��L�h<������8�F+Y��K�Z2�5�0�tF�wp!J�����}?	�;��7����2����Ϳ�vR7e��������i1�����p `(؈�٩i��t���$��sZ�-�+!�Iλ�?�3ru��a}�YZ���2�Geyܖ4��l��5�ba6Xp6g�m�n�����嶖�C�|���j�>�*��i��i�l�l�y���zp���s���p4��c0W�ò�?]3�z?z�d��6Ɔ<A�/;��۷�>�L��e�M4��aS'uKNm�Ì����٧&�dٔ����(�o�:V�5��{sF�G1��(�5m��h��<pcT!���H���%�I�.HI�t�{�"w���׷Q~ϱ�׌���y�JX�-��9�f]w-[��S��7�ߏ�ݽ��[��Uah�6�a)̤�3.3�����ڟw�ڔQ�m1���	�q5��H�R&�͸WK�s�N)Y��c�vi͝ޜ�=�m_����w�e�p�̧S'�z�;{�k"/SJL�f;Ǎ���T-�˾8{s;���cM�޼$�j�aS*�&dT׬Fmy4�j��:]�s�w�����n�>}��kݣOb�����:��ݥRy�*+Ec��I��$���Jc�����+�嗷�/�������,{6�Ly]ah���1c�1fei�Q�m����n�ӇN@��d�Ic���}��C��=�[����V�{�{���,�.c���"h<����8F�&ǌ����BYHw��v��Yc��E\ǝbO��d;�7�����|"���4���̯�v��ܑ��]���<7y��	�r3����5OYA}��s��?x����c��l��!�\k]*�2��{b:�[���=�a�}��`XV]�s��|g�����g���~8�&�?B�2���S?/Fi2�i�e7�N�jI1>�����M=9��Y��)��&{��ر�m����s�q6���(�'�tP���]}&f<d+7)n?c}��F��-�e����M�+lj�oY�}��Y+e�~��;<W���������wq������W ç	Ǩ��g0���ċ-��Ү�0��oJ�mcS}gkt�?c�.-����V����Y��8�,���O����/��]�Ӟ���Jh���UFY���.~�aו��딤)W�'�:��X�[�.4�dE*����X��ɑY0wWN���9��ݭ�QÙ�ѫJO��^����r�F�/]!��el%���ר���Kf���M=%C寸2E��􋤭%Sa0�p��w�L}�ǌ�頻�IW�V�"p\fe�.d�cBd��C���M!"t�3֝+���"�ߣ��z��ҩ�=p�]t�u�e�^�����;5����1���c�=;/E�˙�>���u"��>x�/�ak_�;�Qٽ�>����Y��-U�MO�z�L��n�����`�gj�~��fk9SXH�j�MY����U�V��/٘T*�a��9b�
(,��Z��D���0/�.�iv#XP��h�4$~蠇C�zd��Ǎ�Sd���p�y�+wj�Zl��y���w�~냫$9)�l�Y��B(�fXϩU׆�8�F�k�������i��骤�-uX6��$a�
}zsu��fnv�ۗ��jw�'��G{D���QE�~�]�B*<�/Gq��/�|��'Z����9�aϴ�O�X��P|��V2���ُs���KōSr�V<�2�V��0��['I{;���|����������~c����r�z}״�F�6$��J���}��.�5[\xG��QLd��%J�dd��]�ğ���d�p�r�i�a�kbfDk��.���F�F�>�Z�I�͋4���>��n3M��E-�S�)��ٳȝ%�ޜ�������I�ǧ|��iO�F�-��if��[�m7r�W)�=��a�;.�������eS��y�$j��K�����Ӟ��ڛ��SgH��v$;	�@�h����c�O5�>ٯ3r�-�[�Һ�d]�e��LGP.�V��9͡����?�����Q���O�Zą�O/��BG�,�4k츛q���~�>���z}��v}�.���m�����[�0I�E.[�/�:]�s���IiKޚ&^C��p�4���t�,�c#Ս�3?��Nt��uu����e�"��AD�L������;u�%�n�4{c5.�M��w��>�/jʯ,,��0�����I�k>X{�Ow��Jx��\�-$�K�Ć���w۫�t�{���u����ΐ��lwXL�4����w�u�R�u�W+dk��
�w�L^�N3��u�wv���1�L4U�`�����t����u�[��B�SZ��Gxm��sv�S�d�N��·jȠ�ŉvw�G:9���V�MmuW�s9�<)B�l0A��	^���3,��5�4�Y6��3�����p�-�L���Ưtl�Y}����OH��&�#�=���mbm.�L˦��w����?L�=�~�K����m3#���$���g� lb���N�	�=�9���$wP1�R�H"d���u��9��^i@�"�`$��=[�0�IlB�<\�[!He7�8ؙ�2�,�S�����"]v�Z�W6��2+v�r:H�.WZ�Uc�-���mb���Z�N	���bBD"[�=�N��K��@�vb�o6j�#��SSV��i9�z�ii�촔/3)4*l��뼆ɖ�p�ds׊= ���cj���,�;s�3wf��I93R�-���\d�%���{n*"�r��9X�.I(& �J8���|�UL�0��_v�fZ	iDR5�)���H��í�3u����Y��I8T�V���}.�� /�~�W�<�4m�=@v2���������Ƨ"D�*t�a�ӌ`8L|���$�����#�_J%��-8����0�����&�`(��A(�ҁ�o3�Ç�SI�Kt�s{$���YwX�k�<-/"\��M��6��E^#�#0l"szA���N���G ��zQEH�ؗ��݋dL��':,���t�JH��-S��Y�g(G��n��m�5�[1� ��C⪺Df("/Q`��s���K��~n���f܃��i����=���"�Kk%��-�mj�]�n_�[�ac/����a�S.0K!(x���>���� �F*������Ւ�B��e�kK>�'�b�g�i���UR��!��d�J6�$�)�I�1!��u�E�Q��"=���E3p���!��p�1�#���pF����hDړ��ڱʯ)I� �zZ��p���%oa���Mr3_�eupd
$ �|���نOlu��c2�_2�(���J�����Ϩ��u�3��U����?�<��U��?��9O��G�`�>��� �FO��	�U~���Z�.#�7���=ZW��եUx����mUҫ�WJ��]*�U]��U^+j��Z��^����]�J��b��,UU�UUq���ZU]��ZUW��U��Uⶪ�Uڴ��V*��U]��V�W����Uⶭr�]�ΐ�|rY�$$ �KR�eDR�-��E�����$�E*�	"�(��"2*Z�����D�dZK@���	 ����� ��r��z��������J��U\b��V�Uⶪ�եUW���Uz��j��Ux��WZUv�j��[U^+J��UUUz���Uڴ��QUU�*��ۥv�UҴ��QU^+j��]+J��U]�s���k��s*& e"�H�5������[RKd�V�T�T��P���`%@���V��M�$��Y(��b��ȩQI�P�>�}>�$���o����U�Uz�UW*��*Ҫ�UUTUUTUUU����UWUv��UW��եUx�������j��[U^,UU�UW�ګ�WjҪ�EUW��եWJ�եҫ�Uz���Uڴ��QZ�U��Ā��PFj ȭBI��$a!w
 ���ߠT7!��{9��=�yWj�U]��Uҫ�[U^+J��b��+J��it��]*�U�U�*���UUEUUEUW��եUx���ح�ڪ�b���Ux����t�*��UUTUW�ګ�WkUqW�[mUҫ��uJ��'�Ep1s08�08��	PP�*"(��4EBFA� �Su-��$����Gq��(�J�
��*$n��XH��S�����H��h��F@_|ϟ�?b�(BG�?���������]�q��iG�?�l���Y����"`�6%�!@� � �	��Л8pN�!� ���l��B"lD艂&	ӧᲄ6 ��AĲı �"lD���tL �tD�:&	�0DDç��P��b"&	�"A�6"pDق"tM��N�d�,�Gb""$8P�Ԉ��DL	b`�:&�6!�%�BP�FA���CA�K4"YbpN�:l�l���)i��0�q?[����y����vn'����ø��$e��1bAE�g�tSR<h�#��Bk2�b������$�d���a��Ю��ٛ8Ͱl����#�fm�BF���rL��������.`��i�=a1C)�d��n!�`����ڽ�ʛ�����s�.�L�I�X���;�����#��,�"g��m�H�nb(mI0"��TK�-@���}#	V�_���(
"�>�2��Oc�����_z1�&Ε{Z�&�����u�X�+Ii��1�|�T0�0�Pe:ՠ�� ����I-V�Q�64�����t.�RV}}I�Y�u�}�L��l��������-��"_��.���15*��s.�B!V��I��UƠ�����3qn��eԄ��Bc}}�qԉQ�\0�
C�����+E�b&�~�/�|`("�D��my���ZA�M�٩~�~?*>_���\B6�\R��# �~�Xk)_o��RZ����=j��d�U�BM�4+�ae�Z����8�蒬,.Ql}�m,���z�|uV2�J�j]��l*�˷<���by�i�������h�R[�FÍe��%���qX#�Գz:�O��GzX�깹2�4a��~�_w�m鱶q6ȉ$���r<�K2#��F��M�m�y7�F����V�Xҗ\im�4n�f��c-�X��ɡ4�:��m�k-ݍ��*8[LF�n�w�}䯝�8Y��7lBV�Z�P�vo���E�f+4&�ڕت6��oiMZ�XL٩h�͞R�[ZkuїW�ƺm6v�fV�A�����K�O��t�Ì�,����Ө��1�Ş�r��am�[�6f�6�la?,�����,ɽ�#�q;:�Č���^��-�6��x�73˶p�~��ʐb����Kl2�\�d��de���Z����UM՚��h��2��9���U\b���}�}��~Es33�*���W^��{����fg�UUq�����務���UUq��� ��}�L4ab(��%��<'G$M%?ڿ�92��(O�A�dєˍSU�fctclZL8!s-3e����j������HK�+5�CV�9�5]k����R{R�^͊M6੗d94��dCZGPm
������ke�ʕ�]R��� ���v]lq./8։���Mu�2`%��t�Ǥ��r99�U]�2.�d䬥R1j�ZŝcZ�5�Q֔���~?żXa���B��>���F�mc)GXu���xѤ�a,q�$8�1��pV�!I�I:h�i9'��B{�'�Na�����r���BEIRQ\C�Lϵ�~,M9mh�;�R1ኊ$�2Kp@L�jE�f�aL!s���8Q<�9��9lө�K?c�lm�ƕ�z��?<pDLF	GD�iܽ�B\�I!ģ�z6h㢝,\���\���x�F�2q�yz�d1�+ub�FfSi*e5�!%�,,t�i)�/RH���r8�J�Rd�ˢw�9/޷1��[�����n���z��,%��W��bi�g�L<à�.\!�ͬ�d���S���ü7QD��䐒
���p�.�|�,�h�4Y��������&�<��л��A��i|V�j�XR�US����p��8{�ud�u��$���D��7��m�������6�5�Ã�}�#l�l�8�٧y�M��}��$�����<C'�:ߞ��Rن�b�)>[u�,�`����TH��$���Ѕts�|�s�p4��d�#X,a٦���g{C�	��u�.����t��1%��)4�K��$��q��,�9$�o�4ae�CF�6X�0�8"&�xzC����_$Q�����{ľ4h�	=�0`��_DH[������ύ�ڷ/����ܹ�a�HK
)�C��Iƍ�t�l�p�T��NGN:��G3��ִ�uݙlm�����v��e�;���"�!������<��D�}��R2��Sl2=t�\p�&]?*2p�c�r�\�fa����D�4`�tL3f9>*�[�{��|�eIeiO|���rZ����!�P���o!��[���|�[�ť��^�>�U$�`z�A���H�!��E���YBZ��hL�f-4ɫ�����5oh���e�5�� 	�����)p��Y�5���5.n	ku�����挄<�p��Ms��0rgGe���z-V+�s�觽y��ǤRg�3:�MK˂�)��Y�R�$�!)��'<�8C}���h}Ȩ���u��B�aHw��������匢f��{2��\$�?>w�3�0�!�<oVL�	#�*Ul�M�gEѢı4"'D�0ND�+e�nK�I �o�:;z8��G�������z�J�'$чm�dt��:��$����3�:
�$�H��<�f�l�ra�Bd8>X/�m �g����2ؤr
�H�Rf=SܙpէhԨ[�����N\��A�T�O��ھ�i�n�Ç���a�!�E�,�GO	�0L��0�K�yX�A��$�Fs9ᇁ��v�(pr���\�a<>��Ǿ�I�4�"����g�e�	�gY�9��N�{<c}��kl���a �]�:�1��X��:�>���������>�ÿ�K���!0b��72u���s��yo�$����fD�1�esN�v���ʤ]jY�U��D5��mvXiSv�A�G\ֻ5�ݩzU w��^@�¸ߏp�.��*@F���`�!��M�C�+	�����lç(�f�4(��%���"`�'�a5'd�*��$���$�g����I/$�W	�nS;rq{b��\�p����]��ܭII[����hٴД%к\����)$npN/|�ԧH�9��%� �s;<�^"nC��0���ҩ'�iM��t�;��&�!!�Ւ�n�����lI!0�.p�c�7�BBbx0��r��\��޷MYô��0d�gEѢ�pч����&	����+�*�ԇ��g��m�E�Y��FlB��,��]bm6I�(�|�{M\i�=�p�Y��w��{�|=s�Ŋ����-V�3Yl fؙ\�UIwLKfXZ���l��u���i�ȱiM���UT����!�:�uZ��0��-�l;Y�i �KV�$Dd�FjP�8cG�J ��J?�!N��踽�8~�L%.Ha�	��v���k���+m���p����D��A�y�G/M^△#e��w��;ó����I$!��i#c��ԑ�wI��*��
gj�C�|�c���#�<Ӗ<�f��˕ݹT�!@{:d�kI:J��t��B�\�1㞵GO,�CF�0���'D�0ND��I�I��ⓗ���9,�I�Y��T���Fq6h�.�\���07�H[P��o����)Ik�oe��5Tړ����1]l0���?9a���	��I�4f����v8vC�g3�p���艣x�d�Ԣ7��$	�j�d�d��������2��
�6X�j�Ӷ5��5n/ˊ��1��;�W�RW�>�"}�����~�W�|��ڕ���M8����(�0G�L��ҲCk�母1��qq��1�\_��mj�U�b������lk�j�_��><���:�����b�|)�R�Ū»cUr�X�V�ұx�q��51zZ��1�,�-���q^1���z�|�5��S4��<%"O<Q�'�I���e�<���qZ����X������,�ƚb�1��vƘ�V/o��k�Z��x��m=\^����n�b���_.1���b�q~a�{\...6��q�L\\|�+�;m��wn=o�q��mLt��M8�&�â|%�ŏч	����|(����"���'ê���ƌW׫��_Wך��_��'��(�F~���^��(��Q�^�\�w'�q����^����\E��/������[ӌo��^\OC��*>�̿}:��/\�=#7&n���2;z?���n�KsZ�m�X�������)��|[[��ff~���������7��Fd�����b��"���Z׵�+333�Ŋ������ֵ�fef�3=����U�U�|8Qg
���ٲΖt��ǎ�<'�����p��.����7��BHss�R��ކ����Q��U�4C���0��i(�D��J^�P q�I%���ժ�7(>Tna��H=��i�䠺[$�.>b�~��,�B��˓^�/M=�f�5�Z��[]$������s>��ǃ�6�M=m��J�y�4�8�4OD��pOpLs����V5�#n�Gk��cl�q]E�����<V���c��i������5�Fڋ#�EYS꜔�>��8�WK�V��r,<��s���z@��
!K�0p��.޻qҝt��6���??1�ׯ:>�>�S�m�Z. �	 ���`H�OQ���OF;l��EҀ�l$\@<C�SL�`�z!�E䅇{�m5�ٌ�ڸ�X���j�xv�C����x�X�b�w6�,�oϖ�*�Ҝ � ı�d�
2A͹%0�]}b�: �^��3��.���C��G�r�2��`����ԧ��#R?>�Z:Xu�-|X,�r�
 ="釅��&�]#R��h�Q[�Z]F�=Y��x����uonG��Ȩ�֛����Y+�Og���c���v��)�e�,�h����0L��(�;Նe_�J��Y�YP�D��;�"ћ#)bP~��PM��	�<P�F)&,L\��fQ��QK���c&�x�"V�M�)�����O����X\7m5��v:b~zli�ךCe�ݣѿ�$$�� �x�^���JVЉG\�8K��r�%v��xk���n��l[�&�񲖢����+�b|!��RE:���v��H���:����T%�����Q$��Hy���~U��,Tma�䯎�[Xa�~ϱ;�΄>�L�sE?��F�E$$�U,\ݎ+��Gp=b���9�b�a�7��H����
��j&��cRXƤn�'�)��t!������f���U$.ҕ��^Rl����D��9q�Oe��[4UI��w-j'�UT�l�94y�[��}:m� l4l�͖ag�'���`�����oD��kG���BHI	 E2Rz����"��ERUv�u%U�d3�����H�`�A�')@6�;4UJ��KD��Z�^��B\���A-<{��� ��X*ؼ��`H�0f~!<_F��˳�#|ؓ�cgAI5e��0���ܝ TŮd~���Ɗ�G5-j+�SF�%}G\�UHJ�a������-ۆH����J�>o���T�p8'1&\�b>���i呉GeM��Hm����Ʀ��M9�t!�~�R:�X�z!rat�����j�$O87��4@��e�rX6x݌i��t�0�ޢ�9"u$ĭk�J�1G{i�ç�ͺS���ٲ�t�l��"`��:A0��8�ݻ�ۯ]i݄��@�a��)�ڽ�Y�W����c�'��Ez򦽍V��f�2�}��s2���Kme� �g�o�p��� i���d��5�Y	 �t���R��\cW2�a�݀��I!-����X��M��_�~y:V㵓�m:S��S�:"�!�ak�a*�nK�H=Epp>u<�G��Fv%ɸ4˛�:�5��&�Rޕ'��:2_)�L+q���u����l��J�5#8������ɒ��A<J.�ve5���IR�M˸,e�\��!xE4Q
�C�r@�0��ؚ>�Ѳ6Y��<l��8"&�������V;$��D��H<���@��y�
'�*��I
��I!,S�h�Da �b��1!�	=���� �#��r�E8������KH��=�qSQF� �	�8'�b0�Y��C��(�	E����ITn�ǲ�V�1F�y����A`\���d6�=��!O���J!&\)�������CD8㛐�{���}��Rrf[�~-u�-v����-	g����ȥ٨�N{$�]2Bɠ�i���(<�r�(�,h�a�\�,��lO�D�8t�`X���_�M��ue�˳H:��dH���d�66	N�X��#F�K
�IiBT����i�-%,�!�f�;i��g����7��sf�[0�\Pc���6�U��8{.���`l�w]",�0)�--�AH1�{Ib��OOM葴���L�����WY�)%Gӷ�TʏP��GN��iV-{����WG0:&��&��0i�>{�ً�rȵB�{+�#IH��nn�ֵ�y����E�KPy��#C���ݵt}��ddٯA$!4|?a�ۊgB%B�i��cl4���0���x�Ժ������U�߾�ݵ�r72i���8���f� !G�^6���(}��g8q*T�����^l�d���`Ȯ��5D!��)�	E��hu �b�l���s�J=��B��HUJ�y0���d�駎�O:WN�z���O�����"p�Ú���=����k[����誢��� ��u<�h�UR|i,�)�礘S���:���l�*�bi��F˦��͘��(�%J��_��!��������٘�1ilvZ�
i3��<p��m4e1�N���`�xA�
�(:�]n�m3�꿐���˷R��y7v]��b$���)!J5�7mM��ށci�Ӌ!��<�I�ǜ5*TA&���m7Ƈ�Id�:�H⧧l_�#���}����>8Y���ٲ�'�g��D�:;���`�6BHI	!�LN`�+b�Iw.%�K�M�胛��]1j!��=&�R���:Ѥ�Vn<!z���I�$3���q��}%ފK94� ��P!�e/Ctj�ڻwwM�>4��2ߩ����:>������Q�=ɞ�1��Id�^F��r`gmF��t�\�"u�onhs<��,V�cVK%��.�O]<&i��9���_�Z�p�R�S�Iq�1t�ߓo4�ûv����t�ͽ~t�����"'N��I9�:]�ϵ�TO��I	!$2	�'�λ]��kcI�[l��S�9ɴ��q���/�fD?1+e�}�����yD�(r�u�6��SK�s/]��*���{=��i�gİ�#��Ԭ�_1���kRXxA�_Y�B��M�.�6 ��{P%T�=��ݲ����a�Atۛ0�]�I����>;'����:_X��8���s�OV��հ��)�grfUQGC`� CIg�!&��f��<L���+d�n�k����_ϵk����1�N��j�[\Z�VKn;][ݷ�
Ūū<Wj�V�V�l~i����⛞8X�✓fJ�����N����O������}>9Xk��\m����5���n/ˋ��cƧlk�t�8�-]�d����O~�(�O�~�I?��Ǝ1�,�q��cLWx�1}\W�i�~Y�c����4�4O	G���O�'�aҴx�L\\m���Ӷ�X����<kK������q�b�\_k-�/�i��-��cƘ�����lk�i}v�\\^n�c���b��{]��-\\c[cX����	�O	G����8%aҾ�¶l����b�].8�V�K��W�|*�
���|R����b�ƻV,�z��Wֽ{��N�	��>�,�Ƅ�������RǤ3y>#'�fO���MJ��Sv:���`J��o�$��5h�H��E�	 �i���7]��T-�u�f>e��[ �&�P���f&ָ�hXM��0��B��Ԍ?{��1��H3�(�5i�m���fՀ�Ō�����,��N&cdv! �e;"�O����������3T{H�rf!���B$Z#�b�P��a-F$��16gP���&��U�qA1��*8�j����AǬOZ*�/Z�o�~|Ojϗ�}�ڀZÈ��N��Z���Yg6M�m�)!\	$�e�X�ːVmVVJ!����:Ce-`���bh�  Yy0��"_G�����R�e�9.uk�,���%��\�C-$���p����x?29H)��ۏ#��f���dbq�A�bɆ�ѻbD��kľݙA52��qcl�������髐��0�,�b�F�R[%��#* �0�:�GO�o{k�ipٚ�7[*Pզ�l�M<�����o|�]Ŗ-E�s��ǥ ̠�A�rA5�EҰ�BdI7UZ�e
Ȍ��"!��=��,� 4�;s	F�,��IQ����S��tt1�Q�UaB�*�Y�'E!g8V��TǱ�p��k�i�N��%-zj�/t~Ͽ�/;�]������g�=�yWV����k3+33<�=�W��yz����Z׵��y���{��{�����ﵭ{Y�����qZ���{��V�}��Y�6Cf�:Y���8"&�ӢC
�H@�>ְf�Me�tevz9v�.�:��M��!ۮ�]��mk����.ls�e��mً��Sd.Ήe���L������(6bᆻ�&���vsv�d���6����T�-.��j3V�{��U�b��K�י5B3[av����P�%�	�Ѵ�V��m4ڶ�&���d!�����.%�4�oGJйK]��q�O�""$���>�������g�sl"����{�Ij���4c<er���A!�af�rk�Qy��ש|��4A�a��;����$4k\nBw�!%���%�n\�Eݢe�a.;!�q���n�9��sm�����SoI.���ܚ�x۫,�Hr%7�$+%�n���g����'�������d�$$��Q:]�����`0A�g��]�W:m�P��5�G�j�ݿ�y��3-+%�����|
B�v��$��/�z�@�QĒ�R�=$��:��q�Rśz�ʵ}��wǏ͸���JٲΖ&<~8"&�ӢC}�^vz��8b�2�`�~��EQF����E�m�u�r�/��
I��p4q8�,�����v�rx�Jh�l�y8��!���<�J���d���Lp�܇��X��d�g�COrzhx:_04L�y��n{��������/z��-΋�]1\�O4�"7�V�~ItB��U�4�����0�&�70L=!r�m �`S�Ś����-����.��	��������r>�;�+<S\t��6����؞8"&�ӢC��*���]���Nlzc�12	��3�=��9<�<X��%�!�ܺ[%�:L�H:#�6f�HHE�+Od��|Rl���w	�$�/ �O�	�G�p��̌-������Hݵućb}��Hy�s�7�7U5(h�a�S�����aɹEBG��J9��`���֔�Զ�W�KM�4����j�b `�Q��J�kI0��q4��GD,D3DM
�$<D�dߣ&qhUS�nC��zo��N�у	k�M:vx�cd�4l�͖ag���㇄L�DO���Kǌc�&A3�?sy�c�ɇD�q�&
s�8t����L ���?#��ٻ6�Uɬ�&�Vp��X�9�QH��C9������M7n�)��/�L{$������� He�r�|8YP� Տ>8�w�2lɤ��N`���l�Dg��SČ����:)4Bj�t��I�FBͯ���UzIӆ>%;D0[���NT,�l�f�:X������4x�~ϖN��A!h5
8���}�ǘqAH6�� ��Ͻ�q���	����3Pg!����`H�Y���8َ1#=v�}�*r�=1�
"G��ĕJ�20A�L!	B4���tc���pɉ��h��c�12	�é�4�&�����~�H�xm���y��������uE��n��Z7�7Z�,Ys��~z\�Y��L�/5�sn�&�X���G�&��$8�8v�.��a'[��%i8�$��#�k|���8!NcA���]�n;+%�-ww,�e,�(�;�������L�7�.��.��$&�8�'���m��! \��gE�lI!w���OYߐ�]�Czղ�3;2�J|��J�մe��JԌH:�)aG*7s�:��H�����:��L���J���^�Z����>)�ӧM�S:m�N�co_:~c�>D��!���ε|�J�oYsL��!<��1�c ���y����].%٧��ɦ4��H"`�� �$	wq�4�᫔�l�m��& 臠D���̐��Q������1	��`xD+�͹̢�c	6��9l ��xh��wp��=�Q@��}�g���.L�����9�0&�@��5Sp��*T�0�,X��-��lQ2μK�z�
i�n����c)���o
��j���K�q.�d�A�h�.�1��}5�#6�/�?6����N<q�d��㇄L�D���h�������1���fvu2��I!F\�@,D.�L]ʑçEvj�d����xS{�!tǛ Q���g��tϺ�ϓ)�.nb}�l*�>�շZa˘�R^���r�A�J�$��a�a��\4�ݟ���|�~��:Q�SGk0�a�{RI!9�G�5RJ�^��c�9�>:΃�>��+Ƶ�Mt���.��:��l�g�c�8�K��
��X�HFLO�:7��|�rNy�4y�9$$��v��cN�_F �ƀ��6�mccԤ�t�`xY��j��)%��7��+�����s%�t�g���Ǆ�:tHa9Ky�V�,�֥rNt�1�c!Ƈdh�Tܔl���It�1ڭ�{���d�<W�����5�l�t�����|�wͶ��|�Mw܋��V��!s=4�	��}d�mO5I��'��[i�&iU!�a�3;M�{�q�;i�U�=t����Wg��}��:�i\v�>yznM���G��j��l�e|Xj�:����t{�N�J����m��t�M%�a�:n�ɝ�uZ����4�Qқ�8�+��Ѹ�֤�z���zm�q�f��0��㇏	�"t���sh�u���zL#e�&D����#�a��8�(�zS0S	�md6* ������X�6Չ�宛��'Y:WY;�n�%���pGw6�w���ya��#���F^>�|�δ��K�L�v�W:��݊˄��:Wk��zIq��b֣�v�JX@6W/�\�ԅ���7:��t���2�6칲)F�\邒6ٲS������8��m2�!��y);�'	S���d�|��B�t��L<c`��ʕ%IF�$�T*��e�
N-&��6�Q���fI��d��RC�$l\!č�	ri�ۦ��UI��,L�we&���+���W��oo{�'y��=MGFBs��|��l����C]�$�`�<,^9H'Mؤ�s/��:]4w���Z���!�&,9!�Bh���g��D��!��ď�u�c�u����%"e���F�&��.�)\i3ę����a�i;U�,�:�n�R��{�%Qa!�6�O��TRJ�HC4�2S�RX�A6kD,���I!��mk[I��sm���h��`���O�ߡ���m��6[�>�iaAͅ%�Э��L��'RM��i0x��2�y:STjd�v��t{�V*�Vnq�I�8�$�i�v�@%%�	�/[7=������#����q4�ߚ8D㦍�h҈<��z����'����H��<%�p�\+����sVV-�X���p�~NpOV��?x��\�N`�F	r6Q��:Tc].7���Ʊq�O�7���ۚ_ć���<[��2x���ʝ�8N��g����gK��nj�W��V-Vb�Ū�b���^,��cLWJ�i�]�X�+�b�cOU���|��~cU1�ˋ��J'�$?<P�+�O	xN���1q�m�m�c����qX��=kK�ƚ�f��+5��׬z�+���|�cF+4�M:\Wk�\k�ix����x�X������5�㦴��i�cX�cX��X��5�>cL|��>k�ǚ����v�4��v�j�ڝ���.[�\QW��*�Ɠ"���!��f+�5ڱg���z�����5��|:{㄃��a�DЮD�Ɂ#�ع�9�D>A��3=jG���*xZr3J�8�0=�es>u�W��D��@�x��"k4�"�ȲD��M��!-H��E���F�^)h�x�wHg��r!U@��Ixn";�xZ' 9������yRB�@=��b����ZTg<����&b��� D8w�2��a�p�zJ����g�~�y����i_{��x������k32�3=�+J��g�{޾�ֽ����f{�U�U���{�w~�ffk3=�ڪ�c�{w�ݶ�xm�qǎ<q�1����_��������V���St�^1�c%@(�I���m�F���Α�:@:D�
!�3���B+
��Q8y���
|����x̒f�ęi4�� ѳx��rF1����!�����)e<���W�X�6����0EE�*��?'�{�Iw���,��bi��N��$����6.��^��$7�d�
6�J0�-����JLK�6V��=��*�A������'���=�a���z��T��'���TI1���8�Q���uI���#�h��Gm��6�q\q㏜c�O�vx�"'N�!�Hϋ�.����zc�120,D�G��6B��`���E����J�Q�w�(�-�z������g����ݵn�.-3�LK�ù,q:R-��`����Hq��5j9y	ڕR6�(vC}aI�I�J.�J�#kH0��II���/��N\=�}*����8��-�pzH�T�����#�훯R�����F�'�)��<X�%p�s�ٷ"�6�pۊ�|��6x�p��0DN�l$8򦾭T#��a�^��0�JD"TQ�d?�b> N���-�FT�M���J��%��0+fX��	FАB%��p3�+m���ё��g�Yqpk@fn��%{MI�g��_	<!aO
�b�̻瓶�E3���1�XKC���Z,޺o<ԋ|$���{ϼO#+m�d���W4�7��8nT�N��V��n@�t��2�tv:$I��OR�8zz��O`�$��!���it�d����ӿ���ɇۜ8~T���6SE'�������R֫x�4��v��r���a��NN�2d�NV�%�@��2qâ��뺒`��	�v���ãߒ�6٩n���y���]/�[��~iw�������:��ӧ&�s'����n��]G�8��>*�U&���ٮ��t��A��i�ۊ�z۷ϝ�c�1�X��F��{mGuH���A@mPL���l��ҡP*�\��5-�a����f�
�Z���z�NX�9mI���r�Zj�3�uX1��R8dߞ�$%QUKDM�6���pP:L%�%N�;��ZZƖ��N� ��b��Mh��4w�%U\8�B�����?�uIF�W�m��6
�eJ�@��
ؑ�}d㴣R1�#
I+!)a�"���X���F�+�N����ļÂRl�m���jBQ��ضX+F�-�k�"��[+*�mKԈĶ���Е5����R�-F%E���.H֬[(���*��S�*�0�Ncb�̫F�P��і�md�TYHC�).i�n''䬷"8R[��,qQ�X�ex�65��T@`�ÊUH���1���2�2ڗ35�$����ݴ�0��c!Ih�4T�Yy�$��(rG%æ�>N'yٝ�zzuN�����[��YA�^쌒+���7����~<�.�}���2}i`�:?p=����8�%Ny���p�y��ݹ�h��H���{V��#m1��N'f�W6�g�����<x��'N��z�U!	�|���L�v�$�17�<Ͼ줴RK��(lSDrq:>0�mı�cP�v�;nq�֜n<z�ꧫ��#��[4e)�Sč��L���X�U���Hy��g�~�Rg7��Ձ+kaL�= uǸ�\(���p�:�0�
BJpkIc�t]��t���E�Kl+fݔ0��{׭z���Ia!#�Ѹn\.s|3p�)�MҎwӴT��C�R���t˵��:d��������OM��:m�����ǏxD��!��;��ݴqFKHS��$���fC�!��;M�At�d��K4\
̎l%�}�1�{�R�~�v%в�J/���l�Wwv�.��Ğ�{ϏSdnA�Ԡ鶓�6fIR����K�%�%h���M�c�#��a0�0�9��&�$
JC���r�ӂ��硝ڭh�6�{$M�aƓ���0n^4um��d�IUP��C-�t>�
�2u1Csm&�)�[��c'���|�ӣ�m8ӏ�|Y��p�~:x���:$0�$�k�*�S�9�v�^�ۦ��T�%������f�b�D�P���z�i�u�;�tk*o
TB���:UIbW�R:�6�]&�֡m�/�8��B$enƣ4"�tȏﾘ�V+���6��4���z__]SR��mp]�w��X'��m�ikm�/�Xng�a�����'�X��t��RSb4���N.L�m��URQ�M�,��o>Ou��e��ɞh�[N%��\��0x0�C�z��%�RZ:���m�}����}��<�8�U�Iw�"��e���q�4DٴՓYRQ#j*̱���!4�.��Ҽ�-��R��e�F�����.Qs�ŉ���ǎ�<xO�:$0�ed�Ij����$$��2.�;BG5I��Ci��&#*��]��LKA���K����o��v_���*�V�?I�z�U���~�n2�:�xk�˝�&*���eܝ�4�+*\���M�p�^N����0m �3��
��`�����]��,-?&�:Vm-kqepa��ﮟS�f�,K�8K�Hen�ɼ�ܵ�UW7$,kjX�K݁�u(����n'�I�'4xِ�X�b��.p�	�����Ǆ��ӢCs�Mݵ�2s!ƻ��	!$$��pO�៏������]#0�SNSuΤw8Q�� ���Y9�	f�p��_���S����_%Ș&a`�!CGQ��qJ���{��`{�<F�q�����T�8���ܭ�zUT*U��g �.[�XZ��WsEȉ�[ǉ~�*<���8ort�F�$&��X:�섅�T��ch��t���w�^����n6ӏ\|������<'�N�����,�{�����*���l��q�iV������Oz_�v��s��s��}��Ov�۶M��L�[AV��g���e�,T��[M��a�d��2���eUI!U��ӽ��<��0�.t��ḡ���N�aF��ݧ�\��]2Q�8�L���=l��w�I"]M�gką�:<؆S���<W��W��i4D����=Rx���[��ƻWK�°�
�mb�a�S�k�J�*�j��O�ڿ)�\~jq��K�]?4�x��\_[k��.7����qq�X�_Zq�*��L��㶱q{x�ۋ���[�Zg���ƻW�°�+][1j��Z���V+,�G$�]�x�N<J<C$�(���?��x� �!�(��}�+�I�x�x���x�Bx�	^��/����.�x�m��㦱~W�Z��ƚ�[cLV:k�
�Қ'�,p�W<S�:<Qs�'����W�M6�Z��1�����V.=cx��:kK�5����b��m��X�����|c^1����/��ӄ4��?��>)��g�~O��t*�>&*�7m�����X��m1[cS���Y�{���|}	��G㳛��_������(���@��&)HC�� �z
�3~]K4Jm��^Y�ASXJ���;�����P�Zj�2}�c���ڝIi��
��&�@�P�������W%��\��,��f��������z���޲�]>�t�жe1���+5�|�WL(I!ebWJ"a��J���fc���D	��|�/%%xډ��]:u��<<�;��k!9v\�J#�B04�ح�o����uF�oI,�y�m��b�I��6L:W����E��	���<��AVq��l����	���!ۅ����MH`m2$ �YT�ݑa��0.ZiF>,b��"bY�8֍z���Y�
��i`�ճ���/�a��ЈgIIk�%F߯O{z�r�/{���8�d���o���e��.!�YLjѧzT0�*�M�^2���e%Q�!	���sN&�����EX?+�aJ�I<fG!d2S�M����M��4̈́�.�:�
��e����j���OS�L�6���2�X��\K@�-8�^̳:Uզؼ�Ն�5�r�b7{2������h�3ks����t�i�]u��Bl4��a�L��!�x�K��Ke�d9PJHɇH��i�I1풔+T�o*�%�t3��s�������fg��U�U��}�kZ��33Y��mV�W����{y�������j�Ŋ�Ƶ�k333y���]*�X��l�e�B�Q��<m�;c1�|�Ϟ<<��z�����\X:$c�[���5���ܒ�)%�m��[4��
Ym�0���6�]v�/.��a ����Y]ZDR���q���9Q40�3D�%��H�m]�o8���*2�+$�N����vN�[�m]{:;4�urZK,-�Lhj�4ʱvB��I,M6��c[%{ڶRٖ�h��o�_�V+��SO C��Gh�4��]��۰M+��ֱ���(���y�	��@t�r��9��<�䪕UUU����8ɨ��ٹɛt�����M�I���16���J��ч��|�w*�V�%��t�����m���'�I���g���(�7(��K��m���r:X�h�����=n:5ۚ��Em$�E
!�ZB[�X�$����#6M��k/+-vsN�O��\��i<j<㓏��>�wV7��8xm��q�c��o���>c4+[�5]�h�����Z7�FY�j���p�O���ώ�ON�7���V�bHe����I����	֎���Ƕ�j��uޮ����%X���ʦ�խ��a<h�JS�6mI!�΍<t@�S�]:"y�����a�c�/߅,��H^f�`��l��(��u����ە�N+1s�3t���rl�J�-*�I+Cc߰�6�K�c�͝�����DL`��KVK�Ka�]��ĮHB�n��D(ۦ�q��z��1��<c����@�aw�ƒ(!���I�h�Jn�.Yƒ�u�,9/�S�I/D�Q���0tm����L�N$;��04=4��x�R��<��m��J;����۴���>��z|�F����K��p�#�%��.<q�$*��m�9w��mm�	�28q��K�X6-�0�&�I��`�LJ�UJ�(��˵0l�����X���r=c��6�����o��<x�<'N�L��OotUQUEU}�rY�H4�!��)��y+�|�x��t.?�S�f��Cb�vl�J��]��(X�p�{2g��e�s#�u�|��5D�I�.�w��M�L&��%/A�V�-%';,m�͜_���ө$$z�7<��d��ty���Q��4�0`�G'7=��X���t����w���!
<��$$��?;8m�q�����o������F���K�2QC�$��/F(U�Q1b�
��I��4s��5����!����1!������!륖�GLHP`��Ut�K�':abj��4b<&���\���Cř/ioi��˰�i�%b����E$�;]x��y��LV+�g��+�υ��k��lm��uCK�u�.-�k�[d��?������?\�.;:��IE�MJ%QE1�l��[��zx�Mi�i/����6��.67��rҋQEؐ�h�d�ܥn�8X,��T�Ԗ.::iZ5v����fJ�a��L��9U$*��a�]���m6X4D�..:(��U�d";�o�K-f!YA��̙�y�n&�b� �T0`)�0y9�<�;K`�|'�h��G�l�aP�^�m�Q���Ώ��8����ۂ~:x��<xN����*�uE��h�	!$̇y2vvi�s���*pnf,Rt�4�4u�q��y��r�zL��&��c�=ZJ)��7��,Y�șM��Xnm2�u�zIU�ǟ4���%�Ʃ�Mbl�P�s���~�/{k�6�g�i��(�l��f��u�wk��N���`�{���:qG'�B��t��C�Ӻ�^�B��.����4�6���=+�l�Bݩ(�Y�����M��;Hl�zm�qǮ>q��|��c�1���'�-oӦi(*v.?��X�j��6nB�kS&��2�Csdk&��2�^ap�e;�UŦ�~�*$&�q�)��(�K6-0�p������Y���E�NF��@DMl��o/�k���;��1>����}���S�e�U)��t���L�t�N�i�̃�������#?-:�0�^�׏�{�{V�˂�J�I�Z�Љ�;&m�fmc�-�.�L�b���ągT�w/�̦�}�I6w��bm��0��Kt��Ys�UN�06(���؇ϟ���~^�?i�?;vzm�qǮ<q��c��1����-�V[���!$$�A��t�*ֲ��t�=�It��:����MZ�b�z���4Z�!�\YCs��섒ʂ�H,��6�~ì�~�<�$�~Ïd�a�v��:���־#'d��h�K��0]4l�1$L�S��.;.vXɷ���BN�'Z8).A��X:$CLN=��[��K���4�}�Ia�LF�oB.u"u�R1�Wk���J)����E��n+�:qیc�o�c�1���h���9�0����s1��0��1�m��~�f\A�-o"��6N5a$"mEk�n]�p�"��&�[x���+c1s;b�'�^bQ��
rC"s������z�f�%"�\���[���)�YIf��}/���	C���4B[kz�ޅ�����1X�VsO|�π��m��#T5p�pfԬaM,�շ�D�ȘU���(�J
�iEd����l��<�,����IM ����M�5��&3 O6l�:7��%Z�G���0�F'r�����f�t�a��{��8{˓�!⸗���j)2fBI5��7�L�y<x�d!g-���l���A�߽�,�5+f��a�cp���f�2������B�S�:�J[�����#�id���drZHN���񍬯1ϲ���
(�C^�q�ϟ�<c�1����<W}�'��D�N����C!�	s�?��ۤ�r��{�'L���sӍT�EUQ)�wBS}%���)j7vt���E��� �!P�I�ȧ`�m'F���aM?9ٹ����Cp�1%�i�-�x.7#E���i�zY(�19y3�Г�q"��I5��Ob�<eݚ黭��;����.6�0\h���y��1$%��c�HH�׭N�WmG,V(�m/柘H_k�%:~4'C�ǌ:'��E �!���M+cclq�1��ھ>||%���:X�$B"pJDL6&�6YB � ��EvDЖ&�M��8'D�0�`�&	�`�0M	�N�=x��Ϙ�8�8�=c�q�"CBX��:"&��ؚBh�,�|��"X���'��I��"&��:pN	�f�К,K�x��x<a�!����P�%��6$��8lN��,A=�����v~��ks~�TIʟ�����P��[�p�,8f�����!-ћ���{�ޯI�	���t�zF����Ij�*��IKT�++2>��>���t���`X�'}����͞��5�wٛ�}�WJ�եֽ�z�337��iUҫ�iu�k^�����{�Ut��Z]k�ׯ3339����Uv�.����,��4t٣���Ǐ�c�1�Ǐ������Kw�Y���Մ��C&!��a�=�҉���$r��`��(4� Y�>$d��3��W��K`�JN�rB�,��txC��3�,3����=,+�[�y��N�,Ք`O��+h�ɧT��^�ۥ!a牶��	DH;4�Q��at���B/g��{�l�Lh���5�,;����^��M�I��mıh�L%18)g��u&�;
g���vC�S��p3Ӳ!�V��J��6�4�8�����<a���������+�|s��BHd<.]4al��jUQ*Su�) \6�u<鷌64�,MJi��K�����}��*Oϖs�Nd#'9�����jLt���p�|}�+��w��0�Jz$ι���Әu�(���E4��Da��N6m,RC����L$#pD�m(��aԢ�x�dƤf��O���'�D�x:!¸؉&��Mk!�ۥ4pᇇ#��ėyb�M�ӏm\i�m�x��?<v�v|||z||zvvvw4��9>�U�"��1��%�Lj�>WIeǒ�U�m���U����2�5+�w˵'��6�޻u��>i<O�#�k���b��طSd���͌m]0$#Sl�iLbi�/ɾ1X�Vs7��5R��R�	���h�J�S4i��͵�RX�n���k�G8�����p�d?	�N���]a��m�+�=��C�vx�M4[��b�K�d�0��M�*Uݑ8����O&�5'%+��ێ��R�q�Gf�R���v�)z�2T
*HY�V%�&�x�`������u��R�&h�RR���^Q��%@�����a�����6C5M�e�����R�?d<<�ܘy���4t�;W&�ZUZ��yE��M��8ڸӎ�t�Ǐ_�;~t���x�:t��UW�PO�TUQUAEfHIc,a�ԇ��˵�yrPh��������0��y���
xX}T���<&u�H=�v!O��<o[�z9G��n���ErATE��vi��E�S$���H�\�3�e�Jl��«�F�z3Ą�Z+I!�O6�\��iƵ*V��H��^�g�R����!4�w����ђ�����/{B�v�G�n��=ky��]��4�v���4��G��!��^��Ѩ�Vp�:�L�~}����ȪU:}�w�m����k��Ln4��$�=������(�y,Q�����Ɯvۧ�>c���c�1��gg|PDPM��!$$�� �ޖ�1��#��R_m�*J��d�/Lo�y�{&
�\-����7Kl/:�ϰ��m�p�#h��&buϾ�ώZNSS�-vK�WRL4̷�|����YE��Ѝ3���)0�"D6e(��}���)rv���]˒�t�"K�ZlU̀�Ko���'�	ÒB�[7oׅ�Mi�@�[rً;$��k��)�~F��+����t��Ύ6�4��;q�����c�1���ٳgo[�3��	!$$��|,g��"u�I��`!gf���o���/�@a��5�r��z<�4�ŉ:�F�
[M�sp�Ǹ~�祗���{2d2q�F���u�����
d.9@i8�p�I$0�!7M�n�u�	����u�sQ��u���(0GgJ4g���s;;Zp
oY��9��9�I"#������<4�Q(:h���8����t�8q�q�6�㏘Ǐ�1��x|>41�����	Z�0����E���!�֤�2�L��.W�aָ]a�#Dvɇ������0g&(MA7�D+�,�N�2.�ZV�.4,�	gl��g�aq����(��'��+���_����L�[\3]�mց�i5֝kZ�j�K�f��cF�rU�K)-!	rga�3�=�=�d�o�%˘ljHfBCgw�ǸF�9�^&:6/|:�X���K%�0��R�b�Ar�����>!�ith�J�M�8�D!E�(��Y��,�ѐ�v޵�C�҃����g� ����
g�_����l��b[K�K3��X+��,�h�L'�%���,Bɲ4̤4�M.zS�d<8Q4��)��1��<c��|���m�~ozUQUEU=�m�b��
3�5�%Q�I�LpCF͞ۄ0r7l\�8R�$<t�l��T&��d��<rb�A�|�d�&w�X����D��_B�Dp�`��
|B'M6r��@�͘�?��N'Q�<Ð:���J�66C���ؽUHmzB��(zC&��~>Øp����B�e(�������!�by2�gIK�IAlHHKx94��S���?8q�q����ϟ�?<x�1����:Ƿmi���ֵX�_N�$���ì���{���g�Ş7I(!f�6i�1nq��UsyԓtQ*]4���`�n&�n������P�����R��c*�1uw2�G��"�YJD�k��F�8M<;%0M�.G����v&K���}UR��Ƀ,N"�I�����}$�t^s�NQyz�䢞�P���d���H�J0�t��i2],�2�8�(��}	�<��8L�]�Oe�p��,�fZ|��j�N>m�z���<c�������>�Y'�[	!$$�3#��;$,i5ڕ�ֶu�	m�F�9&L����p�g�
vzx},�[-���i��^ ��/��[VT���N��j3��X�D=$�[�m�a��$����
�U�j�,D�]&�࿵�Xu2Yr����3)���=m%���ࣅ%'��5��}�Qd�r��:e�
19c�t��I$�e��I<�8ĶMJ%Ut�q���N���l�K���$Q%�X��4~�
���g	�6YB � �'���x�ǋ<Y�^&�4x�""X���'J ���&��`��4l��A,A�8&��4"lD��:&	��:'DL�Ή�e�DM���E�DHQ�Ə6x�㧏�^Ȕ&�КE�,��bhDD�0L4P"A4&	�""tؘpNhM%�BP�%M���M��P�P�X�"hؐN�:p�Ӈ�	�������L�Q��")��	I�%�ñ$���"	w�c0�䬯��F�L�2��ƛ8��d=�4�'U�ܥ�-��D��iUc�L���@W"F80����R0�.y�<I��(F�ް���=�|�4]�y|�p���m��0�{�����!eX��]�Z]Yp/&�7y�u��kB�l����[l�V1/{xp�]�6��:����̳]�­�\q4]�W��jV������|=U�AI�-�D�d5�d\a��w��uu1$n�]����E)erI$��R�G�m���p�5����d�$3�"MKi��2�p,P'xCZ�!�Y2kbĉ��.-�M4b=j�-��oL��=7mA���x EadL�d+���^���@�uG�=�F&�@�Rw)?5���}/f��u�mV�0��+v�Y��vK�{�Ӯ����³B"��Z��@\�]Q����/�_�b�!���Fΰ[���/\k(�ii��;��ö�LeO��O�2.d�B����y����}W�[~�K�P,�>r��4�Z;Y��f������j���F��f��ל�ŗ�B	=�Wm�
��(�5�؊8^��!����	)8������2U��[�޷!d�>ܭVu����>�Uڮ��֯��fffg3޵Uڮ�mֵ�z�333��Z��WJ����kՙ����z�Wj�U�[8h���!��<m�1�����c�����K�&+-���չ�c~힎<��Y��Zg�:if��[�i.����Kmq���Fݵf��]|/��6�j�Xzİp7�R��-���Ҵ���o��-B�]�Z�u	h�ٌ��Ґ�l5�7�ns�ifz�͡�ms�;���FX� ����V+#.|��J�!E�n�cM5��g�vHi����,1��cY�L����9��}��=9��W���r]<Y.葐Τ�4]<�4y���)׉"Qf�l��D"7�xX�&a*����c)d�����olf���i���<����	��Ge�jY<]՟�v�q�F��*�6�X�:8�4X��G��u�R��[���ůV&-�H��"��Dt�`h&hX!���֣&w��gs�'Ù�٨�g�՝�t�G�ծJ���8q�q���ۏ���1��1���ӳ����I	!$u�ϳpOq��)�0��8{>�R�7�j�3ݷK��@��^;i:��������Τ=8�|g?��d}�wIû�~聓	���Ô���T��p��ܘ�1���!�;�0�(���,a��H;�ˋS�GK
v8u��f޽�M�d:������2�)˺8`�X�s���d�N2���S�u���/Rr���d����Ev�O�m\i�Ϳ;q��x�lz�>c;x̕�.�1��Z�Z�Zѥ�M��%X棜�쯴������Rp�G�����Hl�v��,�a�ݒ�����)��8?_g�խm��X��l�}7g"FQ"W$݆�wn���y���>�'��h�bM�K�����7t�M�G8�i���m��>cO�i8�5��z�C�;�G	rdI�Nb�Z}v�ZZ��]d��m%&R�u�R�z���ބ�$e�J+)I�J�X�t��Lp�j�N:m�ۏ��:~8x�Ǆ��8t��{�f��z���VBHI	\�\çi8��٫�M%̑;��H�G��4ܻM���l3�7u��ZT*S�I듉b�ݭK4��H�N8�R=8���LH0���,�x���gD��n��1\d��#���p���ٹ$�tPp�&�H�3z�v֒Z��Dv�.0��B���a���RD,@�l�;�U���4�q�l��/#�ރ���<p�j�N;m�n޿?<c�=<xO�K��Iz$��7��ղNV_�=�L@��J�{)\�ת]�R��}�a壦�g޷�OZMx�U&������r�	��d�99��� �Ēl0A.���1�m���bS-��pQ4���`�xiL��fD�\K�'����de��i~䵌�V��:̲^Ym���r���mm�ie[>�����p�14Yv�9��z\8'��C��%3�aIt����L�!!!0a"u��k'���i,@�Z^0ry�d�k�73ڒU�h�.�N���BSt�)L��\�Нc�����Ol6���eM���U�&�R�3ٓ���pY3Ԓޒ@���JI�`ܺR��A=�fz��|����*%���˯#5Y1��m��ϝ�\w)��`�)	���I�Ɠm�i��޴�Í��8�ͻ|���o��O��N�뾳�)K#�����J*�����G�3EM6A�Y4�]���F�4�a|Z��7�Y(�K�(�6�)i�{Y�QkQcA�臧�1Č�t�|zu���.2�ĮD�Ju!M�N�ps\3M���mI�f��\;���y�\�t}�' ����.B�^g��݈6�K1��i���<�B��-�m��V����S����?ap��B��G��e8�2�a���F&�tC�RhՒƹ(4VL�{��L�F�)pSI֔M8Qsr�q�6�o�_�1�^1�����>��~������V+���4gܼR�:��7���C��m��KdԨ�(���G]bI�ވ:=�9x�>@|6?1o!�V�%�ҏa4d�0�i
H�6D	Ȋfm�t���f٧Ǉ�{r�pA4ɝ�Q��I�Ha߇��qr*X:D�N������Y��k�G���ش�����X���k$�ʅh�i-��p.6aV��'Y�tS��䧌Csv]v����˖���Z5a1�[d��,���Z��]�GO��b�}z��m�P���6��m�YD�m�؆N�#��[B��{�|�2�̚1�Z)
�������#Fk\�.�:���vtiYfc�VY���u�5�%����������v%Έ�ռᤃe��U�tFi��).Fhs���YudkGv�Z]�����2&���M-�`�VƘ�HMw�X���Wq�52=Xm6��ᴸd��\�i�o�KH��3̘n�i�	o�InYq)EU:�2�1t�s���ĵ�����E.8ڸӎ�cn�??<~c׌c�1�ǯ4Y���M��dwd����QD���Z�����v���&�MTݑil.�p�Ӝ�C#��[beC52 t�d�pNl�0S"ƹ�����J�T0505(�N��P�G �^��I	!$	�M��UE2ɼl�a(0e�"e����cK�&�;}V������ݲƀ�m�p>��Զ4�H�۹Ya_ry�]��F�<>����]lzh�+:�UF�)��Қ6X0�MT��SP��Ӊ��,
v`�X�IgO���4��ݭUj��z2/ny��>�2���@���i{�K�2�3wL8B>J�i2���̧����.E�6t�gGWq�o�x���c�lc�0xh�?��W
%W]��@ʖ!�:�$jbjF�{��b�Ie!�k�	�g���{Mf�R��˕9%��w����*��֖���"���k)��˗K4��4�[@�7Eaft�Z�s]4�GM�~7�I	!$q4�"ڱ�����[�y���C����y�򐶅7V�TI	�Q�Φ�ypkoM00Z`��M&n��)�!�3̺
_|G��EU��
N���<X�i(!���-I$�dl�p�!��I=�BIwmRh�&I
<�;�9R��I䱳��WL&݁���,������r���cy^p�$�쿳=��$ �`k�$��*��<K��2�:�z\�`�Ę~�^v���\���8Q4��������c1��=gM�~많 ��o�7\,��wa$$��!��$�Itɂ�ƚ��Nb]!��C�In�J���O�p�Rͧj2h�ci��t�Q���r�cb�f��II			yQ$!�S��N�Q�s��\�)��?1�]�X8s{���K�pa�}���Ԭ��7m�[{5���J3 P�K?Y�s�B���������m�In��	�~;��3U�z}ܸt��Q�I.b]�S�!c�˞6h�����6&�(AA>>>aXScclc��H"&�DD�:P�$BtD�b`���blM�� � ���4["X�"lD��d����0L�0A8"Q�:l����'D��$(K4x���<'���NblMp�""X���� �"lDC�a�"'M���F��l�%	BP�A���: � �%	�Dѱ��6p������d	�(L�7�0�8��ظ?^]�L�dC��\;s5�_R "by0�I1�bz��b Z�`��%@șU�=�s��&W9הJ��ԵP�j����֩��TS���w�̎a�`0/R�!ӕ�Ayj�I�-C��[�J�^8� s��-�GQ\Ĵw ��jt�7��8��"q
�L��9���&a�j�h&�v<������nw<�L��:α5�_��^�9�����<�m뙙�z�Wj�U�F��z�333;�R��V�mֵ~������J��[Uu�k^������z*��mU��W$�h�+Rt���:x��ǌ8x�<'L�UYUd�u{�HI	!��d�{U���ED��9Cd-�ɖ�E���,��$���#�DQ����.o�@ۄ7������!� }7?|�+�Y�s����5_{�'�zѶOk5���K.m-j���l��7<�u�<�=�%:c`�=Is$$L8CX�����KL�w������p����J��<��=Y�j�^x�T]�3>�׉D�V�9��7�&��%��t���ƹoM�m�������zvxy�BV6F���HI	(,�7/Y�J��2�Oy4\=lI�|�mtv�+����mu4�1ܖ�2)��T����Ӯ������_']�5!Q��m���0��n�)4lO;rh�I$�i˽&]wE��i6�N����W-!V�-{{��x)-��bD9�T�Z��U�Z�J6�j�M��Ϧba2��`]6��N�zז�q�q�[�lm��1���G�������{Dxbu� t'N3r1T[Ff�e����zY�o�+J�����.Â@�Q�0ij'h�-����M	����V�ZL�E��k�Ms���V��Kv�(��bM�ea
H_TA$@U�<�)�����
�p�
9k"�n6A1ї��+|�2����"��|'��e+v�lJ/%��lD���D�M�&sR��I�Iı��0QI���fI�0�(�SƋ��q�Z� K9�v�Nl�0�G���Ԥ�h�e���=�ִ$�2�k��E:���:�����|s�8=�8���H�qH�@�}����Mvv�F��$
$�dԋ<f��I��P[^�y���rt�Q���}��'CE��Z���Y�0N��x��<xN��2}U]!D�(�%EM�}���@�9�p�vw�)N�CvL%��
��ɴ�$�^�(=�O6Om! LL�ǽ
(�QD�
|��֌���b�����b#�B�:z͉r] ��2!xl��
�5�&*��?��b�j��ZӤ�m�P��A���Hs�I0�ٖ���]��6�R��������ɤVR?���0;r�t�K�ap���&3 K�N٥ͻRT+5'�)���k�.�&	�3ü������D�t4�i5})�g�����x��<xN�g�����~��Z�o�TUQUAI�t�<m��MyN�1@�p�\&{���D��o�!���&��&
L��I���k���x�����#Y9�]��e7��Ur�!P���ç2�H9��b�j�)�Z�D�Í���.�g�m�͜<�5�Z�xj��}wnPl�O��VH1V9���g���|�G����3������R�����73��|�-���ƹo����_�?0t|0|<>��t�0��$l���l���@����v�䓲�[t��'�`���t�l���Q�;9�?t�(��ܦ�6���:ڋ�4n�c1F��%_�Sש��%&^7hɟB�TT��%�R{E�Px�K��d��M'�q��I�/S�tعFIe�mmcf{�ʕj��Q��f!�,��M0�*9���
!RL��V�p�;ѹ��q:\��n~>qp��욼(�M^�af`�?0���x�3�NMj�j��I�C"��4UB�4�HEHx Bq�q��+���h��=h�B�F�㐮�� ��4уʗ\(U�8�Ӓ��]}b5�Q��{�4�Ю��!nͷ,X^ ��R,-�����)C�nȳu���?c��b�Y�>6¶�WY[mpVb��ѲR����m7\ViQc���Vz��?`��a���u,�UT�*N]0.��X�\�ar�̆�q:� M�n��{#M�''�6L�!��a0��x�%����p��I#�I�l�HZL���ɳ	ĳ�-�8��k��fH�	'+���XV_�fHüғ=��`tx�������y�`��f�̛�!r�&K,tL?<x�ǎ���t�HL��U�rғ��I	!$8u��xs�s�']i'w��a7��`ċ1|ċ��;L�t�,��NzI*ҋ�p6Kh&���-Uf{��fZv�K1��Hz�UT���u�i`��6��F!%re��,�fsױD�j�ZZ��^s.6�#U�n�)-�v��yra�癟0�y�I��x�l�y�J������N�v�o&���ғG�$��b9��w�Y��U�t.������ƹoM�m���<c�t�çN6[�4[�UQUEUbd�ٲJ��0auٜ�]H�8a:�P�ۣ����{f����i�&�P�i8ܷS1�2kWM�V�q�U2HN7��b�I�푶,��N���q�Ѿ�$���I��C�p�
�������k"P����p��z�c}��>�ٹ�49�Ƈ;�_jW!���jr�W�x�CEh�bh�����x�������'|�=��E�D��z��Ρ$$���8��y�2���8��N�W%��]L��7H�X���`��9wD0Є6Fk!u���Å��^pWr�$��Ӿx�Ot��I��p�*�F��x�����La�I	�I�O��L�O�'K�N�P�Tf�2�rp�[�UA���$��%���r5T����r]����%:���O���Ǫ�ӷ=~z��1�a�6&�(AAOb�i�sx��ӌqX|�_b"&	 ��:%""t؛e�`AAL�,�BX���pN��Câ&	�`�DL5	�:p����&%�%���"'����:p�I�Ƌ8Y"%��4t�H"&�D��&	B"a�6a�h�,J��2|���`�4A(D�@�f�J:p�ÇL�f�(��jB��j����'�!d$��ډ�7F�WJaIj��f�H&@E���!�Y��S��f-2�B�(�LS9m���1AI4�AU�$�n���ǝ���>Ծ8��������p�4��@-,�Q�׏!��ԡ�:�"h�%I����VSn���%��qu
kI�I�R��Z)�Ӳ��0�CW` ��3Ccl�5���wל����/%Z�>B!$�mx�.#ӕ$mx�6��}�e����@�/�Y H����Km���X�[2*h�M�6��/
W�@J��t��;Sl_�؞a��s}k�϶�P���T��
d��[|3fZ3	.�!vY]nt��Þ^t��ËZU�zTJ�������g�9��%ϣb�t�ME�ÖHl`�X�0(m���cL#�_���
K_bړ҉l�`�Ag��W��`�>b5��(AdM\p(��������Z���{%�-�&�u�F�R�V�q�04�Qfպ�{_J�-a �������Pv�98M]ub�[B��n�$+}Wkg�<�%�F�mυ���� :6�j�ak��B�U�ĊPH\��p���Mq%�a*��FUS��9����7��.�KE�h��Z���%�Ǳ0M`�Oj�%fB�q	��kE}tC�^�묟�ٙ��?EUx���ֵ�zffff{=Uⶪ�Z֟�����EU^�*�����ffffg��UW�J����t�A��h�gK:h���t��8'�	��lٯz�.�.�5(S���ԋ�)���m3u�Ʋ͛6�$�E�<��JLYaHo�>=|��"K\k��[͑�[��c�:��b�=�g�Ĺ�a�v�ةu�̸K�����8"]F��Ys��;A�ŕuг�*h�ujcCͣ�=M+��W�4�t�A����q����I�䄐�@����=S�B����/7(�c�ꭎv�lݓM�dR1��S�էxL��\��._���L��M�tjk5{�2�&%�v��q1FP��:��4c���V�)aM�2�b�wn�=
��)��R�`�BBRu��L88�������R�i���i5j�5͛Y�n���Y��g�|rG���]���5'$�N-͔`��Wm�o�1�<c���1ӆ��û�L��U		�$JM!A�.Rv�ģ�%aۄ�i4<3n�NS�.nGG��zS�� r6/9j��x�X�F����4�N<��RL<7?e�i�� {�K6E����KYo�3��@�J)t�2�)�RB�ތ,�$�2����I��I3�M�x]���Ӷ�i\q�m��>c��c�>8z||zvx>u��Md%��QC�o���4��J���4�xppp�?<n�᧬4�<�Ӄi�t���
2���A����5���9u�h2~ַWXWn��TC����:Ϗpqܮ2IF�SZ4�Ʉ�sn��
�Ģ$c���g7*�U�7�%����:=����g�9��}���e��6rtrr=v�~�gJ��n�4�8��Κ<~�x�Ǆ�2I˫R֕ؗ�EP�y�y���C�u�Z��-��VڵɌN㧹�Aˇ�a�x��F1���F��U��vY5Z������J�vWs���G�%)�'��p�C��ʅQQ��|p"i:��Ѷ�M&u	$aP$�Ѽ�����i7d�3KI��`�³��0].zrx�y$�I{�pl8�d���m:X���D4h���4t�'�x�Ǎ���t³�1��5rH�6�FT��1���k�]+-DK?�}|}�g�4�-�[ ��	"U�Ԇ0v�*BTBl8�je��z�xR&��e)����ʩ0ߐ}�2�dԮ���g㈢��RC ɑ2JFG��ED�[�Cf���a.jJcK��y�v�S��AQ�~\�?���"���K2���F�:q�d~{����s�BX��(���/pt��x��H�bLZUW��A�HMHe���:�x�wǇ�7�R{i��>)�^�߭b�v�C1h��k5��ˮ�$����B�]c�1���צJlP�Ѡ�cX��*:	&�x�m�8Ҹ�n�v�����1�X�O�<'L7��j�(�����Zvm����;?+��-d�ҫ�c���,]餰Rs1�[)��{R�u�{�ӡY9�zn떯�!!	$��S�='M�L�]�-;j�bU�Rյ��Ri�
�Ѱe!�k�kI���0�4�u���L�<�����id��Z�Zֱj�|�^Kb�m��6��+�6���>~c�<x�Ǎ���t��Uy�r�/Xn
(��	�x|i�
ȶYe�i8og�p�x}�)�sp�g�'ֲխ*�5EUi4Cid�u2�L%Υѓ{���Q�[�˜�&%z���Hi�U��fi3�����y���uV�1k^M4�v^67�F��T�&78裠g�t�(�#*�ӕ���O���-]����t���B��H�I���q8�&č���!�d�)�s��]J+5�f�=n�p�W9Hu�O��20���zh�׆)���;�F�#㶯�r�vr~�l|۳�+�6��4"'�x�Ǎ���t��VsN�ػHk�(��;E���B��Y0���I&��,�d=�0�o)�=�����Mu�#$UK0��$(�]�PԚ9ƃ�Ie�{M���a8�䖒e#���|ڣ��a$�K�L�NI2&Ç4�6��zIL�RL$�hÁ�����D����<ba=�S�ӄ$�v��I1祇�gOΟ�|q�q����=c�1�4'�	�������7W=wr�B8̏1q�0&o'�K��%��/kx�$�G1��}�?I�lP�l��ˋ~z�d��b�pV���*E�h����6����:�."SSq7X�n��"1K�~A �Hqr9$���t�j��jL�e�q]˭�f+`]+*S1��\�{�fr����zi�����et�`���I&�F�i��!q�=w):4隻�&P�[sa�y�W�wn�(��9�u����}��u��t��4��DF0x�,�(%lf{�|v.;�z��Q�������e����&{�g�?���J㍻m�1�Ǭc�����%��իV�8��#�zU�B%�^�N2I�|�M=,B���A�?۞EI##�;ν��X�iU�l�^I���CIm&����0���~��5����]�9\��R0!��d=f�u�	�#]u��Z����-!{�]��\�����t_��R��U�:`�ף��o%W��!V���uUT��p˔���FJ4x�f�=|����|�Lt�L0��������LUb��1�8�N,���"&�DL�"%���&"`�8&��e%�AD�D�,��%�b&�N	�N���0L�0DDä�Ζ"YB&�:P�"Q�B"pD�H��bhN���ŝ!��ܞ<&�p�H"&�D��&	B"a�6a�h�,J��2|���"B �"Y���t�Ӈ��'
�fV����d���y�~>/��O�����g;���7�*#�ZkI�pwT!\�������
Kvu�����g�y��f�=��sZ���4��o{��c~�gs33����ZUu�kO�����yUz���Z֟�����*��iUֵ�>3333=�UUq���p�g[p�J㍼m��lc��>||zvx9>��mdI,��E!�6�87��U�O��F���h�4C�K?$R1�j�������&y�|(��!�N@"��(�b�~���CqǗM6��&�\k>g�9���zn~G�C��L�����&X��ӳ��i�>�􎡑s��a<�>2��,kl�\�y8\c����'K�N�d�ܒb�g��t��p�^����Ҕ�ƕ�~m�>c��1�����h����R��'�X�3�I$�?w�8(��#/U*��ś[��f����"Q������']ǓF	ĺͰh�--�]��DQ�u3�$�lPx|gR`�b���7�U��`=��c�E�g�E�D�8?��:�(S�ȑٳX�%B�΃��D넁�9��E�<��J���׬>��dw>y�w7��q�n6��J㍻m㏘��c�1���ǭw<̨���1J	�L퐮J�S��*#7L�eP�ȡ,��[��C A"F4Se\6�)ڤ+���IQ�3����Kq
)�V)�!��abD|p��:��b}2�z�ԃ�9Ji	�K-��w�UPz7��ۍ���l+tBu���6���:37ZLMu:��mc[�MV�n��A�C�w�����Y.�
�l�ƚ�Pe8�6C|0x�{Õ*щ���	�nd�\�r^�k�,l���;�:�s��.y��߼����k����x�����S�~�1rv�߬�w6���J�"���d%`�f��~͙+�h�ɣЖ.���4l���Dq����??;~c���폞=jY݌�#�qUP���L�y�g�_��8�qI&`I�;������iv}��rg��Xv��.������J�{��jU�ԃ1[2%����"jə&f͒�lT�۳�jͰ@�Jc�4�IFdE�s��L�dOR��?�q4�n�=�D*�Аۧ)�����燸p>��M��$�m����IK�T��#/E��a9�:�v�:�M�9�N�e������(�$�'%�A�:rq<dh�$f;D�	$��8C�;m��Wm�o�x��ߟ1���	���7F]ˮ�I$��7��$䖸N7�����I����6�p}��Ifɬ�tg�rRl�5�D?��������5e����l�U�	H��;��GI¼v�'�#�{���4BC.S~7$4j٢��zZ���d��%��>�l냧��;��d��S�zL�������E��^�{<z�ro�o���'q�N1�n�4�8Y�����p�0��<l�{�9�UK��84S�4:�0��'y��,�>�ъ#�?v�k��ե�-�퍶ۺ�7Wy��=�O0N�����7��EUd�-���+�����S���k$�d���n�ܒ#	EJ�5US	�4s�Y��2��,=$��E�5�l���w60\�cAr�h�gKF���	�g�´ucJ4<%	^Z�w#�d��kx,6&QER݁R�£Q��MI�b�qR-e��K�
B��<-�!v>��'�� ��� ��K4�26��6j�}|����N�۲Vm�C��U9xHǦ6:� � �"�T"p���S���E)X�ݲ+�q�"��V,�$�F�<��Ō�\<�:��^G��SG����ٸu�gg^#�d��6�i2G)I��i8����������a�� ���wۊ,:5��t7wj�7n���~��g0�><���:!��H���"Y*\�Z�b�Ĕǹ���:�6���w��uu��Σ�>tۣ�+�6�gM8xN���x�gƪI$��%��Ri������f�%�Z��\a<;=�z�EN�*�s
~�e�a5rA��bm2d��z�B�$sH���8/3�C��O�)�IuWvBY�֤���w�?a��)/.[��4Fq�K��:�Mm/�M2�ۢ�H��tw���UX��z���c��Ԇ���.g9\yl�=���+���vq�q��tП��	��x�d�;*�?96dE��UU9��/cx�g�u�'	��n�OO����̞đ$.S	t�q4�,x�`쐝�����ם�a�CZ:�RZT�wMѵ�Q���9�gd�C�}(�q$��vJ�Lvh��t��������m��N]�p�����?24��}֚֍,���U{c��h�4Y����?<'DO	�GáBε�����I$�9����;;��d��:�z�%d� ��IQ�Y�ads�$I�v�@���q(̑g�!&&�4�[�U7s$���;,�L8cs��E�I�7Պ����l��w8�ղ���ߗ^4�����&_�~��2�i�p�1�c	U��:�b�\���~x/���RA��I>�# I$���P�?����?�Oޛ.���f��s��X�Q�t���B�E�_�1�ƥNx������U$���ZH�UUR�*��(UU,U�U�j*�J������UJ�b��V)UT,UR��T�T�J���U
�UT�J��b���*�Ub��U,R��K%UR�U*�R��HҖ*�Ub�URX�UU�U)V*K)T��T��K�T�X��)U,�R�
R�J�����,R,�,�UR�YF�M*YJSm&�(U,�T��*X�T�JP�R���P��R�U*UK)U)TYJ�e,T��P�K(UU,R�X�tM�E)b�JX�T��*X�R�
T�J��
T�J�ʉe�U"ʒ�*��eJ�YEQe�5R�QT�*U,�U*R��R�b�*�X�J�)UU,T)R�J�YR�YP��T�E��,�Tj�r��J�e"�K*R�b��B�,�U*R���H�R�,�UR�T�YP�E�UB�URE��E�Q-�,�TKDYI,TKX���RRRX������RRRTRT���)*)*)(��)*JK��RJ�J����h�)*RYIR��K
K,m;)0G0G3��dR��%JK
K"��J��RR�XRXRQIe%JK),),�����)JK),�JRX��IE%�K
J�w��IE%�%JK"��%�J��RR�U#E%JJ��)*RXRYIR��J7��F�IIIIIRRRRTRY�IIQIQa���RTRT)*)*JJ�K$���)*oCt��%)*RRRP��RP����
K$Xj�i
T(�E���E
*J*P�JB�EB�E"�EB�$QP��F���UK(҆���Y"��EH��EB�$Qd��H�P�bT�J�*X��%J*QRĩEKJ�J��1H1`�`�`�)"T�*J�%J��*T�EJ�`�H�$�!$�QR��,T���%J*Y*J�T��dT�T��T�*T�R��T��D�R		$�$��**YRĩ,T��b�EJ��**QR�H��R��*T�R�J�,�EJ,5cJ�G&�T��EJ�(�EJ*TT���H�*QR�JJ�%K*QR��**E�R��,�QRȩEJ*QR�H�*QRʕ(�bT����T��T�*QR��**Y)*QR��QR�*QR��**Y**QR��QR���R��,T��EK"�"��T��,*J�
�,��EH�T�*TT�T�R��EJ���,T��,���(�,��)*QR���Q�j��X0X0BX1B$T�T�T�EH�T��P�R*P�d*X��
�%KR**,�R�R�T�R�J�K"�%"��%*������R��
T����R����JRR)b��������IJ��������
RRĥE(R%))QJ�E�R��E*JTRȥIJJRR��d����*)bR�R��JT�))R�����R�))IK�Tj�TR��IK$�%*)QK$��R��RR�J��)R�R�(R�H�KKR�)RR�K*�R�H�KJ��
X���R��R�R(R�R�K$R�R�JE*�E(R*��E,E)���R��IK"�JJY%*Rȥ%,�KJ�EE))QJ����B�)RR�R))JXR�RRȦ扢��%,JE��E))aJ�Y)`�E,�RQ�I��)QK
TR��R���Q,�R�X�E,Rĥ�TR,���E,��)E,R��)QH�JY)IK"�����)QJ�E��R�)b����)QK%,)R��E,R��)QJ���R(����J�Y���h��QK"�R�*)QJJQJ�RR(��X���)QJ)E*)d�QJ)QJ�QJ�YK"����Ij��5%(��K%(�����J)JY)E,��K��)cq�E�TX��T��(�Mi�b�EQe�TX��TX�U*��*��YJ���J�Qe�T,R��E��4��b����UIe*�mh^h�(�X�QTX�R*��U)T���U*�U*�b�J��J��K��X��U���T�UJ�*ʒ��X�UU�UIT�J�U�UT*�UR��*���UUX�B�A;� Q�d�sa0�hL�� x��3B��H
��������+���������ӿ��_bp���������~C���>���޿��;������~#u�g�!�ϞP�%�?��~z`�>���rB|�~�>E;�?BO����l��(>g.��((�
��O��x���������ڢ�����UE ?� DI@���2?p��s���}�C���A��"P�ŗ�A?�n��~����>D?�?�U �}���s���!�H��A�4������_�P8G�_�hV��b~D؟��8���̚?��)�k��tm����@�H+��O�˄�0�̄�?���Ĥ����@� ��!R�"�� ��@֓PRĆ�$$�H��R�)U iH��I��ܚ(d<Q�%X)�_��儸���?Y�8'��$���54"EQ�T@�U��%�Zh@���QT� ]����O�}���o����?�Z>�~���2�``|��C���?����������aC@'�,��H��&��&��.~��~p6A���9�?����
����s�́�C����q�D��C�!�~�X|¾H����~�G�~��ʨ��� @g������>��8p�����}����ՊD @!�U ���p�B$W�	��?��~�D�����x���`����X�M$(���J(��5�$H�l���q`��̖��))��N��r ~l�a��{���#A)(bzR�(�Q���L��4�� ؍�\�:���%�'I��pO�@
G@���!�Q��g�~��O�H�*������
��4�ߗ�)�i��>��������-�|�������$�'����Z�~���h�~���������O�A�w����G�wQU ��+���,�7��`�����J?�U �?y������� p>�~p�'�>a�>�|_�M���a>� �H0�Hg㟸p`�B((B�>�6
?9ߊH������;�`�p~|��?A�τ���7s�paU ���}B�����j��O���?�P���!��C�G�ݧ��m ?|	
5��Vl��ƙ�|'�"�
?�S��0�F������'��QG�A��t.�o�K���f����\�`�O��0�I�Bn))&?�?��_���"�(Hk�� 