BZh91AY&SYp�	�ܾ_�`q���#� ����bH}�           �A�D�4AIM)"�&����4E�@ P
$U�H�*"�D-`�E�
)TH*B�T�l�JG�U]�)B�&��V̨�l1	J�U
P���	v�֕*��U6dE(�Md���AB�P�)� *^��� �A{2��� �("*.�j!@�4 l	HR(�QUR!���U�����-��4j��TB]�
9�i����yD  1�`վ �:�
'`ƕ���lV�� ;���GTi`�ڕ�Ve5�N�r�F�4iY��f�jT��ȍb)5��t�   w�>J����n�J�����)T�Ի��v� ���n�P(:êT�);��R��(;��JP��΂��M�Z��4�T+wCT�����E�T�v��Đ  c�`k�Ji����EGc�@)O^�Ҕ���焕J�,z��T�'<��Ru�<��^������T��Κ]4�T]b ���'XUU{�  �x:}����:�AXu��
P+�ǪU.�UoK: ]�wE�=
 *�n��,��^��%;z�z��=J�[קMJ�Q�*���TRU-��+��  ��9��R��^��w�z�JR�R��:�JJ�l����
Ol�ov�$��okmh6��T�C�z�4�cAS(�iT	wJUIr�QUJ��> ���@*�>��<�Ts�Qփ@��w
kAS j���êR�v��tqN�R��;��UpmM`�j�%*���TB��A!)�|�  ��0}��� �� �M� �m 	�  ;�8 �1@ �kw �\s��1EU#m��� �� �|
ŀ@��pb��0 4� i t��� ��F h�  ]�� 	�J�%)]�$��MK�) ��^���� VV  �;�ti� �p��s0 (�� 
�w 7
 �J�:�6�D�����  π ,X ��� �N (�`:
#@�;���Q�@�W   ��4>          ����@�  CM O�bJR���&Li����)*����     5<"e5J���42d2bCLFJ~�%I�Q��     !I#O�"D�M�a'��M��4ɴ�D�o�����_����?�
 ���7�׽���o��f��]�rd��CUC���� ��=�`�����*}����z!W�G��#��~s�#�?O�a��T���� ��eU_=�"�
�k����HC�y Q���~���eq��1��\eq��WLdq����\dq��Se1��Gq��e1��G`q��f\e1��Gdq��Sdq���`q��e1��`q��q	�ddq��aq��Gdq�`&\e1��`q��SLe&�SL`q��Se1��Sdq���L`q��S`q��SLf`1��aq��dq��&G\dq��`q��C&W\eq��Ge1��GI���W\aq��\`q���\eq�1�1�1��W\dq��q��Weq�1��\eq��&S\baq��\dq��d&WC\aq�� �G&C`q��Gaq��fS\dq��G\`q��	�dq��Gdq��W\e���W\aq��G\`q�	��GLdq��`q��Lb`q��\`q��e1��`&S`q��\`q��l`fdq��aq��WD�dq��Saq��Y�\e1��S\aq��	��Gq�dq��W\dq��G`q���Gaq��`q��a�dq��dq��`�Laq�1��\`aL`1��\eq��Weq�a1��G\aq�1��@��aq��Weq��`�`q��deq��S`q��Geq��Gaq�e�Gdq��`q��G`�`q��1��Gaq��I�eeq��Wdq��G``q��`q��&L`q��Sa1��e�I��Le1��GLdq��SqI��S\a1��SLe1�Ƙdq��SL`q��e1�e�e1��\dq��WI��Gaq��W&C\`eq��@�WCBde``aq��G1���dq��W\aq��\e�q��G\eq��\aq��1��WC\eq�1��W&S\aq��Wdq��@�l`q�� �G\aq�1���\eq��Wdaq���Gdaq��\e1���aq�1�1�1��f ����P�U�pfQ`&T\eE�DaD1�Wq�Wq�Aq�fL`E� \`�\aE� \`E�`U�Q\`�L`�Tq�q�Tq�Tq�Tq�Gq�Faq�@� CEq�Wq� �Q1���`q��G\e1��WCLa�\dq��`q��W`e�	�dq��aq��q��\aq��G\eq��L`�\eq��dq��G���Gdq�� �W\eq�Ƙ\aq��\`eq������\��d����2���2ƅ�}��<ͽ�A��^3e'{e�o/�u�6�U�Ⳍe�3�m��9HfSr̀�T���q`��hU�щ��0�;�.��J��"t���*�cEû�L#��p�Z6Ɖ�����N�j�BT��1nhi��9uhS��[e;���$��˪	��7X��e��6�Yn��Gx�i��K^S��4��8,Z�Р�z�EUU�)e�A5Y�`�a��D��ɹ����WFttB�X�,�NՋ�k��v�����Ēd

��QbA��.ef�����ҟ+(�u��I̶ܪ��-�z��Fl5��-�y2��5�&�*9�<\�!��:�3t;5�ePy��(��ln�)�*�eX�3f+�u�8���&SUM�n��q^���7��*b&R��p]1��]�uL�+]\��*H�vJ̼�^,�O�$I�aK����v��n��SD-�c0j����J��n�yr�Sl�,���m�g��*�Q���S�,^Ùy�3;lY6��+4�^�H0e�U�x)��\)[�1��L�to���q�Fkq���Yg
�B�����b;XE��Ƞ�+!�`L�u�>���Z���ܣm������5(�fz"�Ŷj�ۼɃ�'޳R9�\c�R�Iu��e����M�M�J70ћm7
˥�YW���[�q)�ݣ��Sb�Yƅ��|u>��0R=�U�V2��b8ۘ�4tQ������%e��e�n�Gc�Uc+�Z*�v�N��B�'7P4�����rѢFn�D���j��p'��	��2�<�/�Sn���
G[F�I���'J�oE<.�0[mLih%f���\�����r��M�Zmc��EX��"<�z�n2�fE��w0����bQ�e�\�QV"ɴ�78m����.���vH�ɸ��[�q�!L���p%�,�dh�W:�Z�;�r��:Ği��</��ļ�ޣK��v<M�-IKs(���6ժ!���@�VuYbգ�V!�*i��M:��~��X(e��P�ѕJ˥�`�.�5�ǳw�k$�ʺ�R���j���ʛ�k㰌[	�wnd�u��UwpI@�ۦ��,��Q��Z7�o#��L��S\��1Ul�On����t���){�J���K��-NêX��SLs0��lT��7�#l�'�XU�Ҥ����E�ů&�$�-�فǶ�۹TLZ6e��*����,mfF򰔱�#]H-kM�b��h���i�d�F%�mX�i�ǻL�0�"Uz�Y�ѻq��S�i*(�hVR��V$Ӹ�7�PѺg���Q-G��he ��b��0�5%e��Mԭ e�owC��I|����w����mWQ��ӎ�LF�ھƋ�d��$̨5�r�C��x�,�m�"��<�Ek�m��%�:5���E��`F�6ݭV�[*��J�����N�7��0�,�
��jm-�ݼ��Fc��������[��c���������A�̵!�3h�>��YDYt,^���m��v��͓y�3Ak X�%��QݛB@�IR���Į���n��w*k�PJ{-����I-z�mJ�Q�����f�F���Ү*�����i5����]kǶ!9�S��ȩ���Or�3v�2�kZ�t�f;U��h������^,��p-6ń�Bh��`�	:�Z�j������0��x'�1'yX���y4��+ tP���l)A�5sj�t�XTOpk��0Hj[r�<6U��^�n�n���B]�{8�ʫ�c3T�P�U,:G��S��T�NR����1�u�D]�Wt�)���v��,7S�ل31�W�7���$�
WT9m;�U��i"��V���T�3��n՚�k�Ѣ<I �t�����I��V槺�KCY�7k*�*�x���0�L�j�6ukS1���V^{UQ
�,QYz�`'61o��c���D��*��.ܵ���2�����7^�����Q��[�`�j�.��b1��Z�&�y��Pz���u�S�����w����KsV�ɖ%e�J�gn(��S��1����۫���y.�ee���Qn��؉M�r�\a�t,ܼ�eK�6��6�
�1���۵.��$e��#D*��v���p��G�;��u�ːu��u����
(�y���NfԆ�f�E�����A*�6����5Vɕ�{��m��e�'XwY����(ۡ30ѽI�Ȟi�D˔��-�cۂC,�ZuG��p;�IL�`ݚZ��&�6+r��w�j�*�(����@q�e�	77  !$��)�eڎ��{oS9� W�!7w
OMd�W b[$�O3�oZ��#CE��y����*ɷw�e�[j[?O�Q��Դ�l�Z16Uá�D���&��0�����/.��n[�����t�h�ܔ�)a�1� n�n]�)��M �ݦ�B��lY�/ce�j���8��-��E�,QM��[�qP��r�<6��{R��a20�r�i���^�&���m��)���i<xŋҨ��I�CY���������nް����Lh�kp���
e`���j�&*7q��ƛ��mZ*����*�4/im�������nf����Tr�bOu���e�+L��J��6Q7S��lЬP�Vo5��y��@Mi�+��f^V���A�"�K �"NV��m`ǫ	[{E��ܠ7,I�h��}-�tQ�I����u����%Hq�D�lCtfm]n��Yt�U��h��u�lf]�k~Wt.�[GL���dK$�R�!HӔ�u�+Z��ڪH�����k�=�1�!���@���7������h�k(���9�ͨ\�!v�+z�c�I)�z� �ӵ��0Cmi�ʼ�e��(��b�+���RJ*�Z�faơE
��H����0�hl�h�=���ͅҤ��dl9[.5P�&�$��>�e\٤X���)Y	�W0]e5cS���gx���`��MY�匩�mZ���h�e��V�E���S�bMavv�bX�������*�Y8έm�r�-2��;�Yy�lVACbĂ�$M�Y�iM�[K);˚Q�v��2��n��"h���f��Eo0�h�X���IGb�� ʙ�II�y��щ��b=���Y#Q4����z2H�\��:��x��w��oM�i�M��YYI}*�M�ݿ��dn�u�I(kʲ�݁m���̺p��,�I��2�ҽ�R:��f t�(���N�Z��^c���T�V�Vտ��M�J�d ����R]*�S $˼ӸJ��S�ͪe�]�q�@Fs����YL�㚪&mo
�z��Om��\UYv��-�V�L��Ԣ�.;OS��ˬP��nP�G������cr;�ffj�DۍmG�0\j��Kb� f��u�"�2�`�W�C1Ճ�f7{0��0Z��XIA������n���ˁ޺4%����N��J�%�*�e�[ER��-�N�W�!�B��^;�	�&���k�� �Xkf`��y�ֽe,�q�wf����!�^˕uR�b6�޽EAL�e ,�u`��ȹJYZ�c�M-(@�*)j��S�D�M���0�ٺ�D$ܠ����n7�s4��ٙ�*��b�T#WV��+(C!٢Z/l�����Z���a�M����pm�A�Be���ё.ڂdǹ�;�$��n��%�,�;/<2��.��[Ʒ6�ܱ,��@���wJE�" �Cr�^SSݲ���	�q��-ѸD"lR��]y�pս.8�ɛW��J�n��vl�̤e϶�"��-�ёі�u���hf�`�sز��v݌1�}*ʺ�3;A��gm��SnQ$b��1�ۢ^���i/\0�`��E�F�yy�%�R��DKOmn�<����ƽ���D����Nm�W�wϵ�d� !��1���b�2�uj;���;���G�kN�2���j��G ��)�ɶ{����)埃��Y���(��d���B`�V���[��N�XyvMD�Ӕ^�э�Fű���]�^6[�k��n��v�b�P�pwW�Kfa5ya�W,&"[��$�9�����1ؗ,�E�ct���N�[�V��,l�b%tKTŷ���Ve[�ۮ����bf���	
����,=��yo���˩��6�(���#yn��bR������.�f��:��׌��f%-�ЖކSѦ8�2�U�D;nn�q�t^f�lW�f�� o^�/A�扴�N?���\��N��nД�O�c�LO2mX���h�՗	�wX@G[����*�jj:YZ%���ѱZ���-��g�M)�V���(�mԺ4c�9��ӕ-���E$mb���&L̅���&��:/hM�oBxI!�m�31ɐVT׷R�]Y�ڭQS{M��ݓUlNK�0�b�Nz�d:Y/�`|�<��ټxy�Վ�oi[GdU�i���DdۙbL�:�V��2����ʖO��h��J�/t��j�5]�.�OF�Dy(B�q,¬8v�-ǶCL]�;x�=D�rR�[�6d͕��8���&f�%f�d��P��xD�l�X7V�V�Wgau~�Q���e��!9r�G�[��v���v<D�Ca�NS�H�`�UV�G]�Rٚ�F3��������n#ͻ�zeQ��$�b�L���zj�#B�ͪ�@v�\b�P�������JC]��v+-��11]yqL��E�4,u�1+ZA�@��:{*���fO8.me��i�,�e^e�+X�ƴ�K��^��I�CНLˎɎ�/��vM��i���p٪U�Tw5�d,��F�Ś�KTQZ�X,�۲�v5�V��	��&��L(�b���;wcǖ̼D�JKݎ�o2�n+A*�riJ���Ǵ	�f8
�+����7�;'�c�TI�8[�\wtc��E�Bt��Vݜae?Y�#�����Аd���jN��3`ܻ��d��ʗ��m25�w2���e�ݳ2V�6���,XWDݼKC̈;g�.le9��Vl�UK�YW��������kV(yۤ.ć����v�Q�m�uA�#bS)4/y6���qenE �U� �'N���b�e1V�I�ب��W����I)S�#�����Ĝb���P�l$�B�*�*��n�f�V1z�L�2)P�ܸ��-Yw{V�v[��XU��NH���V��[�Rf+���/KҎ�C8�8�V��gcj��<�o�`�zE��*H�104A-#���y�My�����x�]�z5G6ɘ��_��R�SI�\���QO1Z*�����`8,�2U"�R�P)�&A����Zp]��X-b[�����&��Kz)l!����j�Fs��*-xU�����u�֋�5m#-1W���wN�,	�R%;i�c%���7,�w,�:�y�ū��f��D�ʪL��R�/tt�n����t���"��%=�����cű��h�f�j!v�r��U�̕�����ov�TvN��7
�'5<(�^r!mQr��R�g��c�Q�@l�=R���
����#�Kn�v�-���N�	R­)���di���6� ٻyt���:yy#I�hF��C/AR.������T%-��qP�YM�t��a�s5,ZZŨ�k��勐Zwuw�6"��;��f�]쳯)�d�zk�b��VM{���MZ�&k�
�V�h��R��j�4!Q9w(�A�OeHn����M���_�US�&h�OB6�d��l���	%��E1��Ԙ���6�e+5��-�u��t�գ\�p�P=��d�	�e$�/n�ǀ�ŭ��Mh�%5�nؠ�D��Vb�&F��wٛA<u�,^xӌ�L,��{1C������P�w  �]��0��JŪ5x.ռ٤�e�[њcc#�-�I-;���+1Veid���Ex�K⒑]�d�"qs]ʫ�>Ԣ����q].I5�[<�EY"�-�����9�24�!'�L���F�hǱ]�i%�M[���>�d��n��ZB:�$x�6�$�ƭ+�������R�Y9<�5N(��i\R#��JV&c�P$�i#�س��R�MX�g��,"��U��0�R"��6p��Ã�D�dڨvI�ҴR�-tN�p�l��Y����J3��9�I���Qt5�t�\�%����"�v�Iꨯ�d�I��k[�㗆��M�J��LT�<v��,���M�L�:J�,�ȆY��%�I'�<��al�'iVp�Iy�{��aa7�Y6l��!=9��W�.P���{0Y4=a|w�\��x���(*�Vᓁ������xA,��3vC9e���i�9ǁԏ*U��WI$�V�V��T�R)�4�փ\�.%jڶ���

mn��HGd3���y&�3L�	"���5uZ�Db8����SHj� ��M�.���E����R*df���D��ⴞ(��0�(��=�&��a0�J�vEȆB�s.�(V��	%�Eu���b3���o�Ei�2č2�2� ��ٽ;�ɿ��݇~-��k�h��v{�������V��ġ�v�qD�0k�f3�����:��I�;e�o�X��JR�Xյز'�Ů�;yU���W�D�������t8�d���a�g�2���u.�>>��w4�zi�AMR��EiD�N*�_"�㹼�BQ��-DB�[;g�w���{�����Є�9���3�0�3���Ne�z]f����ѓ|1aD�b+�DĪ�4�J�_f���V
�&�P��ԩ��MX�V��2��ebg!�V���"K(��ĄAY�Aq]"�Z�]��s�"֭��Su{ĢExQ!l�,�,�A(m��E��h�]�&�d�L�#HE#�8�)��i&���GM��k+�}�֥�����w���}�?��}��z��|���Y�$�ï�<{��ޭ|:jQ>�R%:���L��%�m�Թv��2�k�m���g��gi'AK�z8�U�ҍ(�)\�����}|�{T%�Q�+*��7ӧ=��|H�vk��;z���q��':�x��2����>X��=ZY��w�풳l<R�������:ʮ�+���U6֪�#�r�.�X-�����-�\�t�\�b�D8����t�oLV�.k.��`�Q�2�vœV�?tZ�aܜp�uBl}.�iRu��/�:����P�w��4`sr�,� sN��3�?�I7���S�V�|
��Ú���^��y�gT�������]�\�+���:Lsfb�9>.ӛ����έ樅k"�:�����S��;�@s+�h�	ֈW����J�1f֢�'ƍW\��:��9`!��v%ՌH�*7���^^s?���|��y^��h���+6����J��)ң"V��qD�,u���+wN,0��w���;�j<�ˮ�\�ݥ����;��Ɋlq�V&.����:��G�Xڕ`�,����ж�Xb0Gî�+�V��r_ە5�7��J�w���y�)��p��te�v/0�p��[zU���Wh�5���7Cfi��{�ɒ���h;�=�o���b��3�;/1Kn�CH�k��5�!,��~B�S��5���`��{���y\9���20���&��^f�
`ު���=Dj`��a�u*ˑ&-0q�*-���32�&<����$��:�gFp:�V�*�,�-s�yj;��s��(L�^�"y��8�}#��wG!��I^k��u�1zA�����!�\�U5ݤ��۫|��e�)®�@���mSUe�Mk0d��>�awd"$�H��Ҏ��Y��޲��[y�XDʋ�S�çom���c�;fl�r�x�ám��ws�V��#��E�k�+�F�VVԾo���:����mgh���z/FeaS%Q�E ��g�^���g�3�X��}�-��V\r:Ͳ��êa������+|��ͽ:UÒ6^-�2��ۮ��ޕ� ?S�Lݛ:�R��.fL�+�,c����� �yj���"2 +/�f�Sk�κq��ۘ��pU5����Hߺea�v#S��8eu�#���N����8tG�2z.��'d��b�Q�\,sݐ��6)��
�k3�`!Jp3�m)]!�W1W�7�9��As��<��jH��:�H��3x��H��w������A�v�֑��ϐ[.#.Q)ĉ��K�;݂�U�ӡݫ�:fN�ם{OP�\�VwHH���)�.������Ht*(�	���4kk�o�P�o���MvqQ|�Ӹt.�P�z�5u���Nj� [*��u°��\*��(So_�y�@��m$qL�_-P��^n�L�b�ʇ�����fy��g^P��2RYRh�<'z�E�L��bԈ��B����y��4��u��O&[��L$�II/�����{��c���ĥ���mm%s����C�}9�lʧ}���	c0:����Pb��ػ!�[1�D�f�qa�2���ܶ�Uq�L�K��Ѡ����
w7M-�Q�V��8>[����]���&�MUԖ�m,׶�u�&��k�yki�N�X����K���Ԫc%�L1e����]Ư���4U�S�9��t��7F�a��D��w		
��[x��r�ٷS{�0d��;��޿t%]:ڭ�
"�?wc�^�R�݊`_����μv��z�}0��a��@V-��lNN���5�b���pj�׺'���ʝD���ks�.BVf㉴��䣠mvv�[�n�'%��d�B�ۤ���=K�����o����,e�R�惁��Q��[��H��.����Y��tv�ȯI�1���j�[�&�cf���	����ÌSq["7�%2�d�]��<��F�\��n*����[��Y�	U�j���EX���<(v땨-W�f! ���P;H��l�a��9JI�s:��9��5׋Շ��l�pUZ��/Z����:ﰴW��>Xڬ�+�rh�o⇕v!��,}[W~�� �#I�Ys^�wA�ԕ��b�G��0^S%7�{�Y:()s�}6�M����26�7�
�V���]Y5�483v�]e��NI�U�B|[k:��qC4�nM'X�Z!I��{�xewB�=y �4r�5�]}�Q��!^뛮l�+��`Q���Π�Ò�=l��D���H%t�-��C��j��֧�}�j����{�W�f�7/����2�%x&Ǐ���3wKJ�};��wG�L F{��4m%e��������O�QK�����klW�̘.º����)3�;/:bx���U�5O��v7���)59�	����|�F9��^l۶%�;�����r���Z��v���d	�k%��f���5��X�:Mz�6V��w`��7�Agf��;=;F2ԡ��r���.ĝv�.�w}2.I��ۈM��rf���*N.�t�D�]��S}�/z:����OUҌ��p��Dea)nm�N��bY�����A0,ԡ
�۫+�î�1n��0���ށ}{��=�9�1m[�:v_*�
�vK�q6�޾k���r@'��GX�pm��r���;q�:���� ���E�*�&c�SSQl	��X��.d.���{pM�Z9櫔xG0��mh��@�O�k*��/N8TP2��]n�e����<��G5�Aԫ*�T�Ӛ	��w�|�����)�ME�ՃN2��q��J��e���}z6��"6s[ӎ��*�9�GZ}q���eᭀVf}ʪ�m���W�jӐ-@պ��V=f��/����b���u�RSy����Y���sط�y��n�Q7���W��%\�*���[��N�.�L̤vj�3�7©�eӱC%��Jȹ�|��}�!�3��׃������o7V�'��+���vu���S�G��7�V6�ۖb�]Mnc���M][F�����c���m�er�+m���wEZ�v
�v�1��cT�2qU�+�et��k_c뱚�E�"����k"«��롷(�\�.��G(N�hq��ՙe�l�%0�vpc�Fņ�;N�fZ��gv��h���ae����1#�;�]�\7-�:�a�kN���CH����o����v�U)w�]tW0�C�N�jpޗ������ka���ͦE���;�;+��n���S�We:m<��O���ٕv*�н�v[X�;�w��Sd{��ڮ0A���Z����;�5={#섑��R�!�t<���=h�!n�jY��v�;)2��<o7���ٛ���R$��3�e��'��gt�5^Ӿ�����#�C����#<��
]Y��Ww'��YJ��HZ+z��m�ÎWJ���[�o���	j�#4nQ9Wk�G��(=,3խ3@�=���C�UڛjMɶ��L���q3B�zEI��������%,0��_
;}�Tt妯�6�a��%_�s���R���DC�wl;)AI^� F^�Jm��n���̆�z�B�e��t�f�Xo.�r]ui����j��^����gz�9є��1k�2k��kBIFj]UjR��Fؼ6�kǸv���d,�ML{���5&Z�h�ð�2�E���iڑKK_Uֺo�n_
��6�ɝHVMj�=cp�p*-��P���X�YPk~��umX�v-�E�i^[���u��7�\��8����c µ�5SQ	�_w���ݾN�^��Wk�K��ohF�[ag����Ei�ԯq�85�f����r���=���r�
Q� �c��xG-�.��#ݷ�O�0��xt�WS;#���\.����I�9�-"Wi��v
⣶^�Rn�L OD�b�0W����RwZ��Ux�c_4��7�tQ`��{{����ӆұK��!b��iअ��{�v��t�cE��}��{8乬W@d�\�N']"u!i�kj$ ڹv'S�;]ԉ
\ˤ���Y|{P�lGע�����>����n���^:�u����fI�{�H�Y������B�
z�&X��{]J��5��&H_`U�;&�Md���,��юgS��������92T�RU�ꮢ/U�f��*U�P���Ĵ��L�{�&.��͵ة��1 ��RS����6γBQdj]��ѻ��5�n�ע`�bXd3ǲk��#(E��\���ӽ�[�Gmm2&a�7`�9�a�p�&PY��v��ض�ؚ��xg2��\XC���֥o���&_N��"}@f�Oa�k��z�	��u�%́����::�Ci\yu���7d��Opf��v�ZMU�z;o���t�ބ(�Q�w��`���9��L�l���\'�W�Qޤ}�!�V����S��w�˝>�Y0��+t��;	�);;�ܥ������4�J���{�e�wL&���<�Ȋ�B+[��Q�Ƈ�W!r��9��EME���a{�\F8���IS2�08W&j�x`��m脌j6�y35�M�/�&��٧R��\}X�k���h�3��ܪF���v� TV��f��:9�Ok���r�z͹pgR��DF��U��w�ۥ����=P;�cz�]ތ��u��մff*�"cO�J��OϦX�Tl�>*�qئ�֌��Wz�����]��ٍ�8�O(��c��:4�yW쫕�Z�]l�Ng �Dܓ�=M����ov��[@�Z	N^p��\��Z9�9z�v�v�+ŝ�,��m�9n�����c��Ηyf��;�z|$r�Q̒�im�JقS7T�?��K����n��9I��I��m��e!�v�����f]�Y5h�v�J�荌�۹p�ٮ��yQ�ۺ�5�zPD+W��h�6#�\:Ծ{{��t�1e،GuE��m�+(sej�[����$9��5�MR��d2.�fq�靥9����4I}�v;���Uɨ�w��w��,�,X3>��z��v%�,؂��e�|�3����k`��i\u�S��h����z[�1���{\E�o_mG��unGOb�
η�)�z.__��{ykzZok X�lr׷��F�Ǖ�Zeǔ����y�kHر��gz�s,��L�$wE������ɼ�)�MӼy�C��P����Ƥ������3e���,�1��Ґ.�yp���KT�j��#��J���3�t�k����B�![���T�����o7���wn#���C{w~,�S��"�U��V�䵆&%�d\�J�ۃswx��;�]s�p[�/��Jn��L�g7����ܗ��X��@^���"��K�S3�e�/trv��hv���7+�-�{��b�Ze`� Y�m��2.�|��u�f��<Q*�gz4�[�Wl_+��$���;stl�Z�ɭ�h?{ْ��.Z�:�
�A�J늝3q�OM��s�Ƅ�����8��mԬ9�ua�Q�҃�~�f�����)U�R^ؒswv+��H�\�+u��G
w��9�]C%p`ѮI�[��.ng��z��KMT��P�R���ІAp,�l���R��9�e��ҹ����8�dX��З{���RV���o
V��&o�L��F����n�p7��Q*֙��+�9�}�����,�%��M{�K�U�mP���6�uP+jq!���s����U���Yh�S���s��ࣅ�t�͛].7�t{� �q"�$e��sxW},b�|�,��ؿ+<���=i�_\���V"���Jn.�Y𶵪|y�y|�/���N���m�6�ڴ�R��vl��pm��j��Cg�i�w�J��7�M��g_5ܥ���7���2
�;
�b*��Β�Wz�RZg`��P��ʇ\�����qB����}l��3qw1[��Z�U���ϵn"�`����)�30�r���l�]�~�}ԋ�䶪U�4"ڼ�K[]{A>AQ�Ө�z��{Ƅb晗1`�9���G]�X��l;'iwtSq�kO�S���M��N��3T���gsOY퓫�h9V�\���]ndƜ9����I5�7�'_��0��7�w�����|�m���} u�@�o�r�p_;�u#�[����\}���wϮ���O0>�����<w�r��s�D���*o��b��r/�D۩j�.�$P%�4�@w
�:�৘̉����'r>|�������O�'������#� ��~���{����OR&�Br�)5��^�|�w������UQ��?���*�(n��o���'����|��"?�?���!�c�}���_�����?����������ׂ��X&n��t1J��ݷ��H����������%�V�~����O+b|w.}}�w��
xA���O��4�z��Y��b�.�M���0�+%�R��:����V��"���j˦��P[��b`u^��͑Tk'���Η���0Y�T�&���V�ej*���\.��[ӫ�ɾX�RUk��-��3t��ݷ��Cqg>��g;����oU�̹�rs� ��¢ۤ�7��i�DJͫ�#�U��F<3���0;U�%��⮃*��`��/��$��UUM3��t�|��+e4Z]}���z9A[���W�5f���٘Ũι��AlMQ��@f3X����!x�җk(W���-t�G�\S�lh4�Ŷ^����`��E�d�M�*g�@e�6u-�ToC�Zs�E�y4a���Z�w�@���뵜��7�%�q逎p� +}w9�X}o�U����=
h�WU+)K�-�:1�xPN���W�\��[yl{F(f�c�˖�)�^�{�b�|�E/]ԪӔŊ��.��:*�CsgS���rM�-�/f��8��@�Ξ���>Lw�V�,˸f��Cεu�wd:�wN�=-@Mj��;3,�dc�Ru��d��>t�Md<�ы����!S�X���,T�������=~oo�����]}::뮺뮺룮�뮺뮺�:뮺뮾�u�u�]u�_N��뮺뮾�g]u�]u�_N�u�]|:�u�]zu�]x뮺믗]g]u�]u�Ӯ���뮺����]u�]u�]u�]u�]}:κ뮺���]x뮺��]u�_.�κ뮺믧G]{u�u�_N���뮺�ۮ�뮺뮺��:뮺믗]u㮺��]u�]|��:뮺�n��뮺뮾�g]u�]|:뮽:�>^<u�_�뮺�u�]zu�]u�î��Ӯ��Ӯ�믇]u׎�뮺�u�^�����~X��1@�`�S�}|��<|C�u��*�x�)�\sJ�fYxu!򮹭��+�V;٘h�c������&un.�eu-�'��ܽ�+����:�P���1qGh�v���(u̷Q�v\��Vɗ��!X�r���%�:�"�=�PM�]��Ar���UU�|9�W]�o��Ur���8�P���\k�<�ݑ܉Q�i//vu��|f�7����o%�+�	�Mxx�Wk5v<���\���*lp {Y��]���*їV�+��.܅�U�uFD��Y�9β×v�9U�h����� Y�ݦ겷��a80���Q��Ǔ#�2�KY�V�$������w�Kq���uۻˮ�V%�9�D�"�Y����0*N�:�ܘ��>}C1�cJ�K�q���:��w�jj)N�
֩{�z^�8eIS��]��ʏ5�:����(.�9����R���D�4~�,��E`��-��Q`�=%���Fg՝��կ�T̆>�w�d��h B��&���]}�-����jU��Z#c��w>TxËR����-���}S$ү�K��g������/k�c�8��v@����kPUc;zjg.p��D�%EZzq��x`��q5��K�v�m%�Ws
���c����h�v�.\s������7T���s������{}��_��N�뮺�u�]zu�u�]|�뮽:뮺믗]u㮺뮾u�^�u�]zu�]u�뮺��]u�_.�κ뮺믧G]u�]u׷]q�]u�]|��u�]u�ˮ���]u�_��C���N�뮾u�^:뮺����]u�]u��\u�]u�_.���]u�]|:뮽:뮼u�]u�ˮ�㮺뮺�뮸뮺뮽�:뮺뮽��㮺뮺�u�^:뮺�뮺���Y�]u�]u��뮸㎺룮�뮺뮺�:뮺뮾�u�]u�]u��]u�]u�Ӭ�����{�ޛ~�ś+SR,X�Q��)N�6�N3UAy�N�B�e�yz,5J��K�=4�T� ��W��7;ݙ#Tٗ�{[էT6��4M���iF�R��������&Dh�v8.�*�k����]*��2�@7*�ٺ�ġ�k���id�{� $� ��Tw/h��zS���gt���^�ѽC+�8�U�;*�<k,WS�h}��ޙ��6�1��+��i̱9ȕ]N���k,!ww_U�:Yn)�Qg/v��l
�m�j���!2r�]�>C���6wd=&����F��LC�U��\���ﾰ�����n['�U�^=0*���eUc8�����egu�/36l�w�KZ����5k����� M�5u}��9fƞ̗�
���Ax�s7��K�ǘf��tY���R�Dc�w=�*����P^>�U�8t�
��:�<��[��o%A*�x#��/t;�cp^^?z���i��6�������|��_ka-j�p��	�n���-vE���j��:����{��R]=�2Uғ3Ue�"� ̗]�i2��22q`'M�ggr��&L�U1�Кkz��e�o�� ۗk�������7.�_T��]rT]�E���p�@���X������:ܮ�R]x"��3��!VE�U;2��֕��u���W�͘�����01�);��Ǐ/�V�����M[BS]�b��k[ٽ��v�2��߻�8��|mU4)����K��ξ��u��J��ˁ3s#� Ӄp�#Ϛv��޺�����Oy���F@�c�l�rVa��=֥��q�r:ɺ��5%����V(X�c�)d��xB��!�swcmѮ:�T
�C:�=jϣwYs4�_�) V��%E���&��f��^Y]�.�8��Ш�N@�v�t�o�;�tsJ���p>��M�"�	�\o����:d�m�i'J�M��PsgnY��qE�#��m�ku-%�'r-�7{����Y�w�w�n��6_�UxԽ�4i��G]".�
A�9f�y�u巶)[��k�����x��ʮ���,M��Iˍ�s&J\������y���=V��D6���L4�ޫ�9�=�� �>�]��4
g�u����Y�
�w`�Fk�O�̛��w9��ՙ٘�7�Րڵ��[�*L���ҨWN��
���l��Y]��^+��.oh3���7O�)�6��c{dj�R�щ0ww�Xs^|:wU����޽�|�(�Ă�tb}S(@aEdimֺ5d������%�O�
uш��uuY��@�3��wC�fp��7�r�%�-��n���9�t@uVQR�A������ت�.oXFR���C�L�8S{UWؑlzq��ܖ�.x.��^Ӻ!�w��c!��;t���ų1�*����+l����+���j�VΙUBI��o!�l���iU�w{ݹ�4�l4��u��w�Sڭ4/�*�)�J�#pb)����ҳo.-	�|�H�nrs��֛>[��c�O,��Њ�>�ޙ��1ܔ/T�����.֪��=s�����Y��S�J���J�Q2)��~l�AZ�j��Uolj��R�${�m7�X��iڰp60ڼ�j2S3	�rAni��j��}�بp
T/L��튷����9�3�p����]����<�oV��%��.�{�F�2�/E{c�cf�D�USd�uO:�UY�lU�R^*A�з�x�b������*��9:��]���Κ3ʊ�tpi=�7^v�)�8��\�����9n�3�ud��%tM����)�*4�_J�N��
�W=�;��'QƩ�'[hA�7�n@�e\L��u��hhn|uG��)Y&�`�ަF�f^��&�Q�t�ֺ��RWYY�*X<}�{�uv�bq����js��*�@z�	��^s�D�M�P�[�]2�.�o�5�6�̣��y+P
�o6����GsJ�eZ�#Z��^IpC:{z�ƶ�ƍ�n㵘��|��U�Eʢ�$�5%
���g[
���OVLx��}bn�m�wB��Ē̪�,"�Wrw�*/�\a�ˊ���qg'wU�L=#��ⵝVsC��\�gK2rW���̧N�4'˗
E�Y��=y���kgX9-�De��K�X��F�P �k���C4e�[��LR"-5��u�/�dH�P��o;�+-}T��u�O��u���ڐV'H�ɕ�lx%�؆�j�LB� ����:��0V���y����q���ڎ����������yl5W������B�F�1�U�-T�Ho=�R�R���U�:EFi���*z�)�۲������3e!K���c�����ƺ��wҜ�W�^�#@�"V�*�d#]�jG��H�����NuS�<���%����ݼ�,��
�v�3n��	��V�`�i�|U�"X�:�� ��Ӑ.�Շ/jJ���M�]bJW�(�F�*-X����h�J��D�{���y:v���َ��@tu��E��1bc歵W����RY���;kT��,��r�(&�F�ե��h��b�$�L�B^fe�8K�Z��f�������`�Ƭ�*��7x6�lF1ݏjr۴O}j��ۮCy�p�Y�˱�"7�d�u =2�8�4s�4P@hWY��\���5zK��U��`��mtm��j�DK�)g5ی��NЋ[��9j����&eA���)�༒�4���!G���|/�<%�E�7�[pY'{DV�GQ��E�7�=WN�3�������Tiw+q�i��\�GR�s�0t�z�p�����^)}ps������e��*sB�Xw�yb
{�闏�F+�y������)���b��V<H��)���/����D��3p5��1�����=u:jBԔELo>�l�����H��r�׭W"��0q�-u����Fa�.!�%,��JFu��ޕ�(���������41pն���n`���)�}�&�A,\�Ȳ����Q.�1"���.ID�����9n\n�i^�,r睗9��m����G��n��շ57[�ًsB� �߇�J��] �7ǓYV1�Ӆˣռ�|��ͫVʢ��3j`�o]"��Wa�T��W�G�'l�!��nSf\Ժg[�����2��J��ES��$8kMjy 껭���r��kDgu:c�a�.���S�Cm�A˚�X+F�Js�s:p�w}��U��dXk#<�,V�k��������&]��	,�#Zw+�G  �坻���Y��d{��F��f��fT*���D����/���vN5�j�Q�c��덌ޚ65�>�ll,(����7Y���Q�3q	2���Y�
�	�]��=o0ԫ��}�n��quɜc���t��p����=��8�{�Xkl��ݶ�A���1��l˼�湰���s`j�(�7�1��Bˤv��>t����N�4�MP�ͷrL����*+1�z`��tm��/p@�FS	��k��#8��]4�)L|j��7�qm'�]36
������yBv���yw
$b���V��R�Ȫ���5��*�F�3�zzYG�md�-��G*���lF����7�^�ދ�R��vV�>��|Ƭ�GH��<y��W ��:�{��K�[R*��3��
��\����[�gV֪}b˃�	E���)��o�.��9�u�w�qU��A��˨!�K�]�m.9XpH����;�!���</`LԛM-��v�BB���c�U�o���ŌY&�*��F�t��m�XɗYk$=׭���+{.P}v�:�j�'@�����.Vۢ=λ��)����Z�1Q��ޒ�ؠ�uv�k�;�{����1��9JJ��q�Y�f}}0�g�:��^D�uJ�6�C@��J��� h@zʑ]�CL�~�k�!8�s�8-=�K��p�x�n�]��	n����c6����ن�i2gt�\�a��P�i^*>���T�PVVv�d�ݝW<���. �Ωt�o{wb�5(+�S/;���h �i]���R�LhfW,[�Yy��K���D\���R�qS,�~�fQ��`�K.1}C�[,��"K:⇥��V�3&��o�3�ZSr�-��=��!<h5t��Ʈ�����WM����e�ֲ����T��Ҋ�]�ǡTiё̽���G��Lus^_f�ݧ��S0����R�e�)�7���:F�������;S�Qʙ��Uh.k�1۝J������pnɉ*�Y`��o����ï�L��	��H'����	un�M�i=#��\�h�V�g�v,��Sܣf�/醋UhX�Iv��9J̋yn�h�ĵ��Ļ�Q��^��i�DU�U�]c2�5�U�I����������u�jV���o�X7a�C�'e�@�|��m�f�%�w��Z3�S�n��
N��bc��:�=x��Mʼ�BN��2��y7���t=���q��f*}�^(`�9&����ԓcȻ6���f�.��x�rN��5��cy��ײ��ˊ�Aj^SI���ط%y�q8�]���e���Nj}�����X�����L�"�
��O�Oc؆��]+pYǕ�r���}b*�����Ӻ�]Y)}U�R���kv�E��c�)o6+#�6K�N�^u�M�L眃�Wl���#CY~�5����\���=��N��He'��Cr�>��kbdL�G_����k7S�0=!e��J���Z@^�z��]f��y2��1J����ӝvA�M�ڜ�ye�J�ػ��Ac&�Y:����ǆ3��]2��put�87J���S�!���t��������fHjK��ښ)����w�3X7pPXZc9]kIN�9�v�����.���ng�W�O+,Eq\�{�� �dm�ҏ�s�nP������q��V��0�rgV,�t��5͐w	N&�B
/��u�� TTp���$�캶L���
�6��U���n�cv��$�.�N��6���]K�7	����SUU`�;��9��N����Xc���|�n	u�#v3��U*#t5s^Iq<{(�З]Zl>Ŵ��Ɣ��'� *�Z/��_�}����ؿj���?��2����F�,BJR��%T#$ �)10�$��A��Ap�q�F���MLIC*2]RA�<�2�>DɎB�E'�TPJ0SQ��qB�cE��M��9"�M��	�Ɍ"!P���E4X.N8&QTEBi�T�rR.����JA��lDKMЧE4�ZL�RQ4c�O6d@�e��(�p�
���Eq&�$�F�	�m������� ��<s���*���E@�j�%#a ,D.S&>*B6bi��m¡""�m"�
5R�%D���B#���	࿨��`��g^��>�{�D�meEI��w;��&��ٔ���諐�ł�S��En�^�Qœ1���yv������yI����=��T'.��[�/�J}Z�����d�ݠ$9�+��v�f�b����ecS�ߠ�	Ā1Y��+ct؍�ؕګ��v�|��5��U�(��v:����[E����s�(���B�)T�^��ћn-�VȶmVfaqSM`��w�ˆR��^��og.b.�D�et�[�ټ�tl|��(U����f=$�Mf�sk���T�D
jfS�1<0�M�tO<{�.�\41�wi�Q���%o%j�٪�H-�뀫"ӓ��D徝٣��ݒ���b�n�����緲�t���\-u�U[s'74U��Z�gK�y�ܘ����)6o���0eӶ��Ύݍ�y��n�+[�Um���I���t2��ηX�n�a�*��v���ǫA��J�gz�ʠ{'�r�/6��+c)>#��WE`;׌�Y����<�B���&L�8��]�*�����Dəιw'�Ff�+!�#�o�)k�9Yg����r멊���\3�gj�`� ��CGw:�t��t`R�V{*��ښ��V��mh��r�RB��q Ɂ5�� x�$I'."B�%x�B�J��㐦HQ6J���M����8NDҐ4Em�#P��m4�pB�g��(2_d92
<q�!%�$q�\��fB�Q���9
D�j)��D�b'd �F�,��@�b2�8a9aN���Ke�>j@iG�mBa���2&�12h��p0��Am"�8"�%�PA��Xl�#�\|Fcf%
G�s��}z���g��|�v������a��AԐ�
�I
4LM2R����F*�*�&�8Ze	n2���Ȇ(�i�Ah��	�de�J�E�.B$�,4H�Í8���\1��0���$4�@�b�!%�Lh�ēb'q�� [l� h���ƈ-�
A��q�ƛ�� �p��BCp���1�!/�$��B���C⏅�q��Ci����8c"�.*�Da��GȯmO�RT���$:"�&�r4�	�0I��۴�+i������ӛc24�gYѝ�6���s&g��=�{}�룮�뮺�ۮ�뮺�����ӯ��ȥ��$�BڜEmh��)ˎ��1��0s3<��8d��3�.��뮺:뮺뮺�u�u�]zzzzzu�=�sa��Y�aV]����u{E=ڴ�M��r��ѕ;h
,���Y��n�]z�kR3K�{�dIF���we���5��Z�)�m�k<�&j�֘��{���l�dl�mn]��c ��r��%�[}��;�{{ޝlݐ�{�xF��^�B�=�s�m���Mk9-�y��[�l7n͖,���n8��m���q#k�w�<�mv�4e6�������mإ6ѻ�w�h
S��}��)),�tI�rL����T�a����[�^X��۲���Ӝ�å�����G��/%�-������/�[��S��k�������y��gx�|)
H� "@�༦\,&A8J\!���ȉ��J���("
Rp��ED����9,D���T�����k�oU/�eӺ[�n^�0�,Џk�_U	sh����+^�Y[7$�7�R�2PŮl�=];�6��ΠR�!�3� ���A�#D��� �D�l(�p�ˑ�l$���iDҌ�&b,(�)��O���&5ƀfBI��$��p������%��b��.���WC]+��`�+��$�+p�̲��	�MU�Y}�v�D��.���3�9��:��3n�5��~���N�3�����e�ҝ<��ĩ���h_��R�HʨE{.�"ND�m>�e�V��jԧ2����B"��o��|E,��~BIv1J��L��c�jT�7���F�r�[��[8�O�U�B��#l�݄������T�P�p���-�yR82tL�љ��H9u[0F�l)e���a�ŉp�L٭��l�}[��)E���m�L�a���A\жD-�<��(h��Pqk�e������x^6v$��O����U�0�B+�1jD7�ΓL���8�aϣ-���$���u^���2(���,Zʓ@v.ǷoU�<xig�fP`_�,�fG�J��$�ķfPU^�7u�F�Q������N�ט;��& q��U	�X�n���&�9�����'�x�5>�*�_\kB��Ɇ��.��,.v�0�}�Q��Ѳ�����$���o2���M5V�[o#H��E����9�எ,���άw*��k^�˹rA������:ᕃS�hf�W=��oD�tu�ﺹ4�i���ok�a�͚8I@e����F�o6Y��Y P�H�gq��ъ��ΨӗE-l��E�pI��Xs�ԅ�0�ע�&��d��������펛����n��{ڟK���9�訋v�BA���)���^�1�)<���y1-T��*�I2
�$j-²��Vz%��1�**�\��Z������g�`�zX���BqJ��my�f�jh��xy{��v��)i'���� ��W�ʹ����W�j�W�o�=p;�xD��jttWL� #y�{3�)�������u]�>�}�p���hf=P�9QN+W�NnE1)U
����b�m2�j��{+�'+H�P�"�Q,km	F�f+U��}9�<%Al�����R��/�5����Z���2w"+�{��(�l�{=�%+�G��3���*��`A��{3��&��4TQ}�;v�N$llI*�Tp��R�^��خV9��bt����8�Qv)ܕ}�j��k�B��4����\ڗ�>q>�����P��m���]=�/5����S���"����W�SY��������������[�I�v�'��;^�-}]{��j 7�� a��Ăw֊�������4��/	;f4��i�lA���P���KF�e�;�ąx�-�k�ҧw���ߵ��o8
#��}N]
��5�Ŀ۷7j�����o�~�K����yͨ���l>���
�8b�e|H=N�0����ޙ[� ��ғ��;�z�گzfz�y�(7�|��^�E{�Jʓ�ִ�YH�v�����(���x�fq*��u���@m%�-�G��� ��
�7�5�ʟ^��>6K@8(϶���Ml�m�V�k�������PF�Q52��3#u)����E�˫�w͆ŚR�Po5�61@žh�`�!�j�k�ED	L	DϪ��\(��
]e�Y���j�u�6�@�g�h%^z�jv�H�o�lVeө
�摒��ʫ��r���;��>�l4Qͭ�����f=m�خ���l83q��fI�x*\�	��^^�#��P^�ͫQ�5Sd�y,��B g\�(*[�>H��vD8�t�ᦳ��w微�4��z��,�}7[��D�)#l�hR���|>�q;�"滹���g^�%"q��#H5�%)�e_�Q�&�p�S�Z�|?'Y����Җe>�S���l��I0�A6-���+����k�a*�EK���.=�N��k[�ܧ�nh�'vP�u}sE���#<��ʒ�%��G#_B�ZE�S�	N^ZeO�A]9["+�m���o�l'Ue��P�g�ݝz-�
�{�ҳI&�[;!�͐�B��l�{`
1���5������wc5o��{u���H�Z�ve��c� X�͟���R��K,�q��G6*o��2�S�_ג�/�Fd0�[4^a^˖��K4�~2��W���H�X��5���N�lo����Zri6���K���hɏ8[�TxI��;���P�$��J!��T���)�vic+&s�r<�խ3mma�f��"��,rA�c��εs�K�g$bLEW[}�H]F�%����e1��f<�^��1��wk�p�_�b����31�B���{��S7��;7wr�.��������E��GiN�;�q��S�w]󤁾ق�mU`�-�+2��X��nX׮�����l��P�d���	�Z�X�c��Y�d�ZQ:I+�Bjn�`d3���*�/0 �>�0$f���5oX�0�2_Q;tW�h�KA�Y~y����(ILMJ���^��N���ŊNJs$��|� �Bu�VBט�`�i�W����L�6�ς]"��n��}��]fnu��^���d�@��ˏR��*��YVM%�ھǸ�l�t��Id���ϩ
nW�z%4���O��n��m��FH3R��
�f�f�灨
*����,�I0�%��6��S
��KV�:���n�m1�4��Q�wf�Ƒf��N��N6SС~��1�����01I��yPg�.�|�ֺ[0���V���g,6����l��G4�8
��H�(l-���4d�5�Avä��ܶ�m�=�����wY�t%.5Q��Y^ϩf��5���W��|�n�>f��W��]��D�+jp�R��%���*v��4��:���'J�V��I�O`��q�@J>���fd�5J`w#�X$�w�5�� �|�7��]��9��W���ˍ�������2�>ʇ��dy��k��ؼ59y�-�p��M�v�Yt���+�	f �`i���i4�/uiɉ����X*S�7�z�l�&IGi"jkʄ^�+!��V���!�,�>�����0�S��!W�YՌ0i�;�GĜ��i��Ŋ������4`,B-�\*�05=�쌖� ���m�$��.��_Tu�>��
 ���W�o'�l��>M��ߞ�U&��M��s�s�b�j���|�y��R��ݕ�-<�v�S����b2U!��ͺocK��w�e�r�O�r��J�U�(mf׮[�=;Wzw��.J�)j�9�')�NSp�(�-�w'J�c�O��9OQS��؈U@�y�VҲ.0���i^�v\l��2�Бk�c�AJ���x!��nF�p�3ud���8�jX��L��7��I�&�2$����� �>�.9��^H��y���x��G���١�u�I����2��g��{7j��3y^N�X�u�:��>����c�VO>k=���Y�2R���uZiV��ޝF�&�����}5W�6K�Y��ff�)O�R�j��)��	Ӛ�!,�<�N�{�V�y:��
p�RZ�JD�}�ۧ[�pi˶ԃx�N=n��Y�S�א��J�e���KCU�R;$ِٽ�M�C#&��X��,Z�骝�bj�Z�Hs����=N�e���	���[�e�l��6lL³�[������_����s�[�[1Q�f0m��i@վX#r�*�4&-�pߧ���Uު�8��ש?-��L̰�U�*3j��}���a�M���9skص����g)��/�D9�
7j�B�R��8۪ufDV�̇xL̸ٓ����-ǚ��Fd�T�R�BzrX��S��������6�P�r����~ iൟ?o��l�:�#p�އྺ$P{�wMjX��j�O���D�Wt��Y��$��"x�]�ehj��b4������\7�R7]��v���T��ޞ}9m�z�m�vqȆh�$0���1V�f�^�c.	*�>�^VG����{�����uT�wt�,�cuZ��E�[�џn��A���8p�8"׽��5���١�_��-C����#w���'@I�f�܉VR�ּ$D��!���lS��
�T����mi �\�j���H��(-�#*�H�d�MA&����,�j�"6��n��NzP��t�I����vϮ%�7�f
�� �J�͒Z�f���W
�"X�Y�'��ہY)J>ߟ�W�߻.޸�8������=Z_5!���/j=�(�6"h1��$T��T�WT�F�h�{{�H铱�渕��ӏ�ᡲ��$��J�e\��|����dCϺ>��z�ה7J[]P���I�6�W����s���屬5'#]i8��{��Z-���a�ҙ�+mv YE�7����XBP8.��i]���n3�z;�'=I����o�,k�ŏ�G,aQo	貇
^���%l[Ζ�(M`�Oim�	`o��d��x�γ�0�뗤���n� :���]��cP�{X�.��J���l��^�C�3x���e�.���0,,����[�r��`�ˬx^X"�C�4L�LV�!gK�'��*	"�=���7�����0�r�e�z5p�K�no��}+��TJ'��T���{��fY���/1,��o"�L�cx	UD���tW���n@�&F��i'V�cŊ��@��M�ګE��m��I��m�u��!�
�n@��z����=�^A�X�����A�ȸJJ�*tk�Cl6ƄF�g���d��>T��u�nc��+U%Zs<�ױ:�h��e�a�0Yg� �=4�	�5�m�v��0�^ܲ�ω#Icbs_d0�zKѢQʖj�+b���yx���q�V#%R��4��L�7N��ڞ#��F�av�����Æ�a=ڇؙ�~F�(�4�$i���TK��lF��1yR�Vsh�p��d�WY�P:��2�F�%0*�����dp��h��@��ψ���(��]:ϫE6�fd��/��c���v��(fu�q���-�Sc��ݩV�c*��{���*Dgtz�;9��dr݌?]�D��]��x�Qk�8]��:�w���x��R�݃��V?�8��}j��n�>��م�"����"$+&�I�ZIݵg7�-�ڦ>ۼ�c4��&�q|���8�I��1MOWr=w^�Q��	�v�e/2�il����1�-U�^�@6���!�i�cV�d�Z�c�Ӥ�f�JRFH6��P�L�4}���x���ϯ�sGQ�HCn=l)�/gbI����/)�zgq�_T��f0��Փ���o�}�H�]����g�ןz�B[��ͅ3��F)n����a�P�4���͘�S�#6w@Ki)�7[[f
y�"�.�ܨ�XJ�T��6��2�o�O!r��G���f�T��M�)ӗW+�c$�Aڏ6�m�`l�"�Guu7��"�ex���g��ݳ���>w�7�l���z���*���^�n��'�����{|m�"�NY̝����=����N%�}u<v55;����E�rL���8VQ[��:긨� �i��H ��8<='��#�ͮw�)��6-K�9�0t«�,�n��Ѳ]׾/D#,ݗ7s��J��ٙ�|(:�(�j���[ʎ�S��h��#��d�$l6ť�L���w��pa��I�g(���F�l�we�t��b��]�l�En��`�PhCW+f�s�&��`}[�'b���H�7tc��7o�� �q�.v�0��Pc�t�31^��� r���b�C2�_�gL#)��6I7�T��r�ҙݶ�L��7#X�<!�{Ν�-�Q�i�r���V�E��=ǵ�в]����q5kr�;:�__[�Ws̒��e��}��tw��k/C��r	�R��vX�(I�I{��޶E���[����n�NLM�u:��"��K5����GLy���l�0�^���҅�I'j6�M
/tT�}��)��
a�嗵Y��_�{����*��҂k�p�Dh�#xH�zH/���9�UK�GZ�hmQ42��ԒK�3h:̗��ld�K�!�\��cK�ɕ� ne�͙��j�m�Mƃ�ˎ�r��F�x�p�w�6H�}ӑӾ��]w�
7�S���c�ntl����X�78�̟- X���P�OcHi,�W�Ui���l=Z��J
�Hu�8��#��NQ�XT�;�@�Hm�\�K����V�>��y/�+�����ق��9/�����̾vF䧘��
ˣ2��-�N�2�:�R���Y�["�0�r�;��(��T�����.:�n�;�0����l�����Z��D��]���M7��ü:V����W�N��.[��]�_%��;n�|�!��*�lέ��6.��1�Ϧ��I]��ܮ�wui�z$�X���(p~M�0��8����P<������U�ԋyN���*j+uMn�F�ݑ�T�R��B|CY��4z��ЧDbs; �1��GUd����C�6���4�����uauI���{���Wݒ�C:ȅ���oTΖK,�.��ӲF;܏z/���MH��1�dHs�L�Ǵ�ti���:�A)�--�t �|�v7�V�o��2ħ�/��Ԫ'�X�7{�&���k�-b��J��:���b��Aj�T��;#hU�{q��C��w�}�S9��yO,�;x��6��O��D�f�{��eM8�2�����ܦ�,swQ���.�_:t'A�X�T�ѕRc��ު���wB��$0o;V%qׅ�@=�^ꋁ5�g��+�_��d`0o8
-���ɦ�+c���
��S���nc���:����Ď�c�D��^����=�����[ko���}/<��{�Ҵs��Vc�>�[�]��e�mk]��j�מ�{��T�r��ywO����1�39�s�&G2!+,���==>/o�����뮺뮺���u�]x�������ps͇�
��̘��֬��n^��3��ﳺ�l(6�d󜌖�%�&.q.� �Xl�ݷU�yG���{���m�f�v+���u������ۧ�������}��}��]u�]u�]u�^<x��ا}�]����]q^5��u�����z�Ͷ�f���5�ڶ�����_U,lۛ�~��{'�rߍ�F�to=����{��|�5B��]�������kl��MϽݤ���k��s�����N���z޶쵮����>���w���ܴ�v�z���'����}��o����^�ΛH�����^���ONw�mϝ�m��7�N7mW�����{P����}�p�i����gڳմ��זq����|��o�^�}�='�a���pv��j�D�������H�jI#�{g��<�m%9�y�k&��z�mv@#4IH[�A�gxYf�����c�X`��ׅ�ޱ�f�Y^b���Kl�8�{[�/l��%�
lr�u�޲'�{�vvGXmd�"��~6�_�e�G�"���)*�R�[m�����k�$C�;��eXYYܗ!NQY�q����8�#������mf	�k`�-�q�����B�v���MK%W��0��2�UhLrG��)�x,��&���D�c:����."M��zQʼ������<����Ub+��o^k8j��<���c�O�d�l�n���gAJ��>�q�7MoS*oG�77���{�h#����~�QU�+�����[�����
�;���_>d�/��՚����7�7�qv�D��>7��^����,>�|<��_/�C�VҢ��z�^��u.�a�z�̼J}ɾFkp��߾d��U�o ��g���N�?�t?�N����o��ϼ��Y�[)T�%�/��k��h�=5��;�O<'�Fq�c��j�?�Z%xy��a�;���#j�{��ֆ��V�U9����c��D���ǆ���)��{�Ut|j/l����o,O���q{��+lJY�c:�W}�^���t�1��8�>����)��r�kk�� �\?W�</�#zL]q]g+/"��x�pY��;�_�$É�W��lu˯�dWP���%�.��Пg���v��C��F?��w�~��`���އ��=%���<������\���F���[s5�7V�c�7�����`y��9���t/�Mz%�i�g3��CHk�旼����U�u��A��Wvܷ�)�<]�/�4�k���r�8��kb�s�(��H�ME�ư�v�og
�Z�eEi���]��ʯ���K�D����e�k�v�J���t��Ղ��"��d�k`n6�C�<|�q����eZs$�����e/��y���g�}1.���B��|w��&/5��s�����˽�C�u�\�� ��A[�t1����
��W���_yՉ滕��(�������Y�2�2EȞo�^5�^��}Tδ��o�C��"�BP�g�O��Pƭ��H�w�yƖv�M���v��$Y�����)��[��඼����5y=�p�Z��ˋ��;�J��֎��;E���xx��������`	O^J�HJ�e���Y��Ng,��O|=��/l���/�pvޔ��YΙ�&s���ϼ� ���������o�/�:M���Q�3��p5r���^m�d ���d5n��:\wN��9Nm��u���Q�+���}5� �5�{�xM����Eyn�G��>��v�����z��ٮ���f�ɶ��&�lk��7����"��{;k�(8�������?y�m�;Ʋ�5�/��u�ϼ9�����O�b�k1t���=�����gp*�7����>��|z��a��~��׌�]<�;��NwA2dV֭"��R�RюHe�����wb��T2�a(ȟDe�e��N�L�؛/Z�[<8 ��p�����W��ś2k�).r69����f=s�o��P����&�T���N���)b�Q�;�mY�W����^^�|�G%�*lz�{�c�'p��u�`�{o�h�+{}&2�j������d����1�nq���9�p-�O?_r�����тXJ�M,廣	��XG~@Q{'O V_<���?��X@!��	�����n�����N<'�r�v���[y7��^�^����\B�;��6,k�>������@�[�a���`gC=�D�
��<MD�~�ʝs�ɠn�4^��_����e=Ԏ��L��O1o�>tg�nP���<=������6K	��4�e�s�tG��o�<��i�]V��ϛ����Z�گgN��`�2�%�#`v rO8�	u&��0[��T�O-�Z]�6�"�GU����S9��Ύ�!���>�a�@�;X��o�S{��#�P#<^��'��u�4��[�i�Y�3U�(yg�!��a��y����&�[��L;7\�>�Ú�o�	�ū^��O�o��b#��wf�!脞HM�03^����N��X����>�I\{o�0q��.��t^k��zO����|��?_5�+�1D��ρ�]�F������	������ǰk�q¤��Ѡ�>�]�9n�f�U��Ұ:ԊL�<Ѹ���q=�*:�V��^�Ҿ�:f�[�n�8��%�nw;Fa�7��*T�����n��=\+o��}��ؕ&���1L��$�8moF�����=~8����\�J�������/
��*��~�#�vp�����f~	�K��N3���"�<V��҇��k��S�0Z���Ts��<����c}�{�N[����mA�ݚ���zU6�i%i`Θp!�q1w4^��!V�E6���</��P�Roc�����<����6�����C�1L�-�X�L��AyOm�C'ۤG5_��n�YY��fAݥY�����:~��5eFR?���0R����f|�j�c�=>�N�j����ܕ��+z�2o��T�����#ƹ�����]���KT_�[ۼxHwknnN\���EA���1W��ʭ�fks�V��ZOƽ�ff��D�t�/�� [wwIn�/B�N)��1�q�B���oͅ;�6�-�UK�吳uX���n�J�C������=M����3�AB�MN���zl��s�Z�Ǯ���x{|1���G1�L��<!��R_��W9�>?Be^�=j��(����=�(�t��;���70�F���uB`�֑�ʼ.�S�^v���ob����Ee����5(+��uޞFm�ߖV��+$4gm��	�/1��Y1�٦�r��s���=z��zikW��q���.�ʭ����qr�q��1�Sǜ�F�'B7�,�6����=G��Kc��;�IbJy8e�x.��ja푹r�&�6�bw=$m�����?��*iZORxz5��M�/��G�"��<#Xl���^ŵ��$�M#�n�{]���������ܼ�'���Cc���q~,~�bj�-��P��}	���?������h����y�^/W�`�i/\<r�.ǎ���ӯIAi��Iz���[-}���IZt9��@��)���M�Q��:΃Օ���5�R��>���!f�7����ԅ �
�-�� k��1a[M���i�i_a<=�ٝ��&y=��.�d�6@s�l�n�'����;J}�a�P�C�A\���f�P��g��h�И	�LSЗ�zV2}wFD^쀘*�(����n�3�ͥ��aA��>�)��^1��@B�7�i�C�l0�ߗ���8�ќ��/a�Y�>�ۙܜ�5o]gjr��,���L�z����N���,?'{Et[j��-$-W��c(�wۙnUWe�vs�b�jd�}�^�S�+�|g1��zǄ�n��:��L2���V��N7"dc�ɧS9�xx��z�,���nos_r�n��ty��A�Ư�~y���B�6������7o�n y��K�c1�bj`���^�ok'���<=�U���2g:��{SV���aB9�-c�Fv_Y��-^��֎�Nۻ��Kw�M)�i��3kӝr�U.b����ɪX����ܗ�ʻ��-m�n�4�蛫-���_�������9�U��=m�!�����0���Ә��vO��˽������J����Ke���n#K;�Nd�Cǽ�����c��`��}vkB��������d�y����lY���my�t��)���Q����������|�.�l�p!>�D07 �K�J/��zgK7)ƺoz�1���&��i�����ޗd<�zi��{�1Q ��R��M�Y�*�����óaI�ǂ�y4[�����07Up��>M&:���~c !�Q����L^����W�,�wsƎ!����pg������c�<�^�B�����m��AC����f�����\>��2���~�}߷Îd����N��!��2+�Ʒ��|e�NǥyL�ڟG�_��dlo�?m̦z����{��`��j�=	s�s��b\NdM���<�$�%����T���1q/�jSCĴ��g��_ßv�ш��&U��|	6����P|y5j�	xN���m�3j��{l���ZO$��;pE��h��K3�8"Lx ��o?yPj��}c��k��:y��{`.���nKE�F�2����״~�����\$�� J.����в�Q�����e:8��:�JU:p�i��vwD�N��V>�W���|N��d���"H��f��;\�P�a=Ěeu.a,�0������=�@�Ge��q㧻j&_�^�ܲ��e>�Lu�A��L�z����cUn��L�@*�O@A���G��^]�-3ϫ���ă��=ŷ'�zn=$\�-"n�֭�;ۆOkSձ�����w\�p{�R}y6�ޢ���%V>a��~�y��r�ei���x�+5p����xt��9�}�\��(#����-���Οm��r��0�7}�Tͽ�����1����-�7C�8���M;Հ:�L\qz�� ��+��tz����&ԎN3��g���䷬��_~I���`U�t����>���|�H��E��<�ͯ̓�:����#��Ǵ��
���Ӝ<��W�3zcW����h�l���zn-�<0;��}\��9�c	��n��y�n�ևީ��V������%�rJ���;ݼ0���F4�~�4&</>���N�JU��J#�m�{���Co���~�ܟ�1� ���_i�D��Ҳ�����A��>
�h��<�7�p��BCw�����%�Ռ�@�W:�x��xõ� w?s�K�z�����nC�xi�����%5D�N������)�xh������iu&�ɘ2��5S�Sc��{K�����U�fıִ�
�,�Λ��\q�Om���/�J���~��ܕ�mWS�;D�j�޹�8^���,���M"�Q�ݏKGuu�6J�F�f��;Yu��y2'A��h�O838��5d��,ⲝ����4��������G�{���w�<=m���������ʦ2�Y���f��H���I�\��P���{=�/f�K�Ñ-�N�ΠG�p��=(�"O��T�<@����ħ3Z�g;`G|h�ʪ��������y�@��[5�'����A�Wz��@���z�.�Z�D��R6+Ǻ��i�წĵY���x�F�3�K���|�h�e^0-�<��zn^����C�<�y/lc�v�к�v���<q�xfvS;zs qz� �┻O��'I���'����;%vܙ���=��r����e�h��{�9r� rx��A�#͢�m�����k��ӊ�4l�L�K��h�0h�� ��O@��w�#���|�=����fgނ���uz��wt)����q���M���y����6>;��_L\lP��h��4ûA~�=��6}{�"y��ͩ�ՑFD{��i�Un<U���%nP��]�ګLѫL���ٞB�����s�co�Y��VM�&��z;}X�T����~s�����x���B� �VW��'!Ŵ{��z2�D�����O��{/I�K�ކ���̵Y���6w�L5yM�]^ ]mk�Z�8�nt�ۻ�t�سF�e�oN�@�O<�H#�(	�$Q7�����D�&������0]�ćWe%G�ׅh�
\�P���7�.A��Ӛ:1�+&�'߼����{ށ��z=�<��}����_��Uz{�O?c(��{�.��_�{���
��z�+���sA���UOPc���#�k��vo��l��r>x�����*�O��1M�׽�iBo[&�;��+B��0C������x�7O�Lp>�`6�k�P�BU��q'�t����2oW�r���Ң�їg�噶�|9�g��av�2Ǧ5�i���홚�Pmg��·���]J^�dk�r:0�MVf{�v����xĳ�����C����Fx�c��m���Dn�����򇅹Z���zw�{r�"ϐ�~���t3O�"�F�A_2GN�ߗCD^0��gRۘ^�om�t��4���ɡ���m)��Е���_m�OU��|��X_��+^9K'���wҾ��s���2uv�&�2�����2���c�wOW�ECǠH�Ǉs���TQ:�;[����,�;C�p��i�_u�� �[i݄�
4R�d�)��W��C�m���\Mp��u���S����a�����s��{8�thCz��&
�u��p���-X�؋:�N��B�����އjdm^��r�S��f�W:�ޣ0VF8��U�����ki>�8_�̯��c yD!�T�ߤ�e�`��O�l�8Z^���if��jptz�o5al�3-c�b95S{Yd���^�Ajlȫ{��z����@�z=� 2��<�3�$�z�j�~�]M�P�E;�3����ވ��JTX�=��46�o�]�G�a�fu���.�m����<�����>53�	w�-���w������%V��n8�A�9ӫu\�L=�H�׻72�<��-�׻z`&�L̽�]�����%�^�P��U�s��xyG�B~�>��+-o0G8��[��w)����~`:�X`����iw|H����V{��ū��[���s�u	���� �-r�9��è�~ow8����N�Ϸ �0�E}��R^�Ӿ�y��o��<$~~`��T�6���4�$�Wk����������0zلT-&��V�[��H�}ϵ�]aP ��Es���_�#�ra��_� A�z}��]�`爌�qT�ub'��^5ͅ7{94��f���z]Ǉ��j4Ϗ0�&�m27��������f����Ȯ<O��L��(%��݌�xw�c�;���4��"KЇ� ���eq�5�a�N�nuM�\=�"�a�2�&�]�+�Wa>�nx���>����u�lA�A_dc� 2%�:�uL0̑�m����2�vMyNΑ�C\p*��{��m��i#֥\j�񌢱�3\�[J>|��n�h�h^�F�`������ZI���
�=���b�5X��N�ɒ���n^,���Em��T���.�[ǅC4���������ze����Fu�R��T�1,�省g���e=n�>��3N^G��r�u�83�@�3v�N���G��M�Vx��ԝ#%���>;�0�32�Fe��\A<�-c��J��ve���^��*�.)"._wP�{��R9��X	=[Y�y�nWwH)�H��;H�ɬN��5��9e�FL�5�nG�fv����⭙C�n�o&�7}w����
G���]+��$6n����x�O��t�D=��b��@�ѯ�~W��W�mBa���}[����U:BM��x��q�OpIf����p
��p��)��%7�Ƅh�3���/�sY��Ƿ�TuKz���ח�=�-��-欩�Y�:y��E�h���1H�t#�w3$m��C�nК��z�[L�qZK�k6ɭz���՜��{D��p�iNi\fZu/��r��Y��7��]�fB���۩4l�UUθ%���o-�b�쬣���L_]��MSӬ�㼷����Duˎ�e���D��ϭ����	x���՛��s�Ds���]H�%�b	�.2v��W���u��n�9}�}͵gM{��$���4v�Vݰ���z�(}HP��c�=���l�!m땽G޺ӷ1uo3y�š�����v�D�J^dg���N! ���{�p>^;�|�t��w���iJԊ�&�xy�2NS&�<��BҒ��k77hs�EFw�en����s.e�T�l�܇�7����<
�h�w'kM����ʹ�z{�#i�D'3K��4Y�����,�g�h���m9�z���к�
ʋ����Sxս*���9�ף��n��@np�˶�
W�Ǒ���@�p僦[u�*#��^·��0+�(�5�]Al�_����hPYu�"Ns����t���ھu�b١���NU���NW(���j5��7ԗ�:��S��n�L�����jCz�+I�_TOZ��N�2;2i�g.��s����oa8�\[�w�)e��)f]�6��w*#���
��芾��" lqZ39ЊwA�qF^t��*��3��W3Y��7!����,	\;)�ͦ������	��!%T̠���GJ�Ӳj�J4]͜x�y�5w4v�]wѫ�d�d��՘T�R�cf��*�cJ�#�n#�$������E*��K�z_�]�$��2�1�v�w=9���$��q��m�f�R�w9`83i*����gk�&�����+�|�
�hv�bat�.%w�q��l�LKG�u.���L�P����ɜd" �Q\��N�N���8r�hBI�j
:;~=�ʂy�BT��FQxgx�����u��}����}��n�����]u�Ǐ}��TE�EL�=�9%ָ�@�V{�Ғ����A;m/�;v�wO�����{u�}��o�����}��u�^<x�������5r��Ș�2�2�#��3	�]�S�6����Z��KkP�̿<�I({��p�������mY��ΜI��U�8w��nm�Sn��䈧NG	�C��Y� Xږ�g(�va����G��n^Ok�`m�u��+m'Q�[�m�Ns,�(�@����:9�h�ͬq#�nŕ���k2T[7d��\C�6�');lJp$��76��J:�88�m�6�����=�H�:9
J;.�-y�pS�n����L�Zel��N�wNߋX�y��q(�gH۲�ΔB�i � %�i"7N��Ƈ8�w�SF�MGD��@[`�F�?5@��)2Ѧ�P6	#�H�䁲"E�HA�0��E5��	U�P�j��v��ܥ�t��M��z9:�9����Η��������Qޡ��Z�x�^�vꕼh��6�1􂊄'HP�Ƙ|q��p~T�D�HB`h2��e�����e��m�j6��F$�,�Sh#(3E�#FY�WM2j�q\a����|����||`  �s���m��M�s���E��>�rMpsc�!�wI����E���/���M���\h�}�B/�e�
Taz�~�x-����f���tδ��ۏNЇm�8�[�\훖�t����6�n�&a<���tǞ���܀8'���)�Fo���ݐ��済|��Δ�4�.�Vbe>x?c��q���1���^��Ȑw/	����+u��-v)*����2nѮ�X`�S¡���I���/�ސ#��UƯ���^G�9�FH5vu�rr���ၑ:(0�Z���44�R�)��e�d�`0'#��N0�����⩣��V28��a����_��"��z�a|_�s�׽�_e�jU���RN��'F���Ү����N�1��I�����ѫ�-ύc
��w�/�Ku�X�v���'�1P��r:]�C�zN��<X3v���x�ϯ�/li��ק�#��iG7_O�
�=I��ޞGEo��W�����;��0᫲I{�~�v�}�GFʞO������4>e�4��=�Q<�����T�����^o�>�g�����&�B�_O: ���/ '�������~�y]�;DzJ2���:1�훰M��,�}�W��}]b�.͓�-�n]Nil�ĞQ�8���f9\�
�W9 ��6
}ɨݺ�67z�����\p��J�J�A�Jq��^�;�pb�z��Q�+~wwl�����u�c�x�}��wa���&�u�'�LW�dEt@�J�9�/^w�xh�O�#�=�F��7��L���\�m�$u��*n�4u�7&��3M�Am�`�z�Sש��x5���MP��f�|�Mv<m�FcaE��9�5�J%��l��p�"yd�	����PYs����2>��<;�܇�k&�96��U+yU]�n�<Xo ���"2�y����NI[��u�+0�n�u���7��D�1�v,��&r���m��lO�7��ŗ���Թ���֣�o����w)�=��w=��Ռ36$��c8�SG8y'M��ۚ�j����Ah|'�H�|/�H���Y�fӹ�@�j,}w2��L�p��8�������W��� ����>�{ߠ ������CM���d�ʗN�Fu��W��h�L5Q��	��%�^�P!h�`ΞF������%���y�M8iubV8y�ˁl\��`��qL��	}=5z��nԬU��U�@��֕�>��w�xYy�B������?��"���E�N�/��.�׆��BNB�F���B#m���m�[�"��ǴN�{�L[���hc3p�Z�}��b�.�zK
�!�[l�\�1r�!�"�|���a�Yd1A�ieQ� �p�$�dH�Ͻ�yœj`�y*�w����U�X���ޞdZ|ԡ2.Q��{d���u|��է~��|����χ������e�]ġ��c%����ň�8?'��������M��:��u���챻A�q�3W3���I�߼/�'H���Y@c��4!e�c���P��}ύ�Y#���~�N;�\�%ۺq�7x{1�1A)����f��zigj������X�D��7 r�aO����[ڮ���ئc�!7%�X���x�{�Vq��Us��(g������y��ӎ�-�l�gdu�bЙ��#=;�,U�F=,��ݞe4���i���cv{��0d��`{����8�:���m�egj�+�p��q��9<2���)9*A1I����O'�cݜ����ܷOb��^������;�E��13km�z`ٳ"z�r�Pe�(��Ż�2Pk�6��ƶNN`<����-a��N�A��@��c�p��X���z���nt�6y�]W/�3��9lˁ�G3d��<�F�C3��N)_� ��N�e�;��u񠽛�k����4�I���[ӳ�R�s��o��\[�<_��z�]q�UM����0z���� ` Ž�@�������٪�T�WW1Fv�Y˺��9*[,Wk�a�1�yc�iW~W��Q��5�)^R.���{W�g$��$NWo+t��v�)�i��.$�:W��nU����c��]|��ѹ�5O�s���'u�'m�j��_R|���x��<DU:�w�>�����<Y�)���eAI��^7��ZU譈�Q���ϋ�(
<����CGPYG{�h��+�^���e׻�ݏB]��}p��q��`�zZF�f`�!jS�DE2j6#�v<"��gj-��7	'��Qwfa.C[���7�~���*�n(xK�݄�
E�))S���:֔�]]R��g�4�b���T:�O���υ�����N�`�x���>]�W�n�a�;/�[sq[(���Ő��]ċȲ�T��uB���<<�
��}|�q�ȧ�#q�c��j�3r�)�]p��2:�82�wM��tyc����|jg�]���݆�J.:��!������_�����Q�b&�Cz��\��ri��� pnj��Ms�T[�c�M<'�[�Ü]V�Q��?y�]7����4���@�p$��U����L5(���Fw �ۮs�U�Iv��P/l��4sZ�Q��U;���xsM%��1����8C,r|4Q��/��2��n�y��v���7�w\�[^�z����.�n;��{��E�t�|\cς�z	ƴJ�L#�;5�7k��|u s.K� ����]ѯ(�F=lH��9�f-텹{J��)GIe�v��^���Fs��̾�8Ǧ��f;S�委�]F����n�S|�I6�����J��lt�ړ�|-�f�����q4�^�N?��ܽ����ga|7�x�u�*�.���ǌ��)�����U�Vw6�?�ͭ�nN�C�GƝ'Gw�5.6�לfE�k;!��_m}�=QƊj�g�ʲ<h���Z��ƹ9����9�������[\��<��d��,ܫ���#�����x`;j7����O���h�#4�I�2-�p�֐!�.$3�k��|!!"����o�s���5���Ȫ���^h,����w9.}�ԃ�|���҈�!�>��9M�@��Ϸ��t��g�����}C&W�߉���d���uǤy<����l㸛��`4n�T��.qh���<_V�H3g�x|�"z��.Ň�~����H��k�H��R��j� �
T?����lgE�;��z�[}a#T�>�\�i�M���<3s��1�d���a9�a^ ���֔**;�'<Z�'f�C�:n��|j��12���"�G�Roֶ���ud�ǀr�4�3R�o�����_/�'�О	:j�VU�r�����@�?���ߗ�wUH~�5#ň����l��^ʡvO=wG���D~=5�ѪZy϶t��ď@+���~�UN��mH���3̦�/t����U�MǦEE5��{2n���HkȦ�,YyMU�{���u��S�^�-�+�S�qn'C�=Y,���ysT��\nud�ǳ�s^��M�m��+;f�J���Q� k��*��r��0��h�\��:B���jX��jt�SNw��O~피ǧ EZ���86��*h2T�3;�z�z��M����G�>�l�<Lx����{�eR���v`�~!�y��zaB.��[�@c��1Þ��7or�g�( ㆆ���֤���"xyS�:�`�y�����g�Z鰺���L��W�pHΝgu�Bow����p��vF�}�0�T�4U���c��.��y���x��|ŭ�sky6��:��D�GE�`�4I��X�n���C�GOs��FΑu�g����N�F���}5��'VT�Tr���=4N����rZ�\݌�swy������Yz�o'2���L�D�mE}۫��	�C�+5/�Ty�yn.s�3�H�Fg�b�Q���XSz�X�:+svs�/l����fx��[�y�Ư��R����,�9<���{�*��a<��%o?>v�r�ƛ��p_�}�݃�s���|���*|�rJqv�0��%���u�:����n�����9��g���hW<��sl��4>~�1�[z#�<LIN(�x���C)�T�Oe��<<u�:m����j��}�k^��P�S� aw�4O�T���p���o�W���h,8eU�|��Zz�Là>3���Z|9veBK�������'7c!���7�2芗k�.� \���|��ɾ�N�cW<hV3�&�*om�wI�/\�����w�ǘ��٧Fh������ޟ7�� ��z= {��������.����~�/��3BTH`&S�gS퀜�0���b!�M����8�:�/I���o6�&f���vi�j��x��z	C2�aP�E�)�>�˼
�c�b܌�+�G��cn��EE�vC0�w>�h��#��CT#�>)K��X�`/^/��+]��)}�)��ܤ���	�8eǅ�H�@/���R�2����5k��.�(�&�c6�<�9��f|�^|8D�!�_l}k*�=!���˂w+�`D�|3x�=�0�rn~���}�Q]~�	��z�X�x���Π���{�xE�><G�g8H�@c���X��qP	�.�z�9�����hNU���ԭѪ��hAm�o�7�(�y�1_�ƣm�S�;��pP���Kd������&gm��P�oHnfSPr��I��~>�Ù���"�W0c�^R�Rp.%�}����Ӓ��)�zή9����3Յ��q�:�Y�+�L�s�yؖ��]�\¼�,���s�a�ɑ����жN�Cņ�px�O5���K�c!d�Y^�<LZ~a�0��זV���7N�����S�QC?W$5Wq2�'��YZ8���w��_ʓ���3�{�K̕WT=�f�E�A\>�]Zˍ>�,K˙��������mPݪ��b���O-�m2+f�/��J�n=Z�^s�>�wn�w�y�~^3�� 1�<x{��w����i��l׶�;�>D��B�"m	�Ͳ,�4�9])2���-O
�ڕ��]��t�)�Ӱ��<�/W0���k!x��@��a�O���#9�>����g/W��l�K0�{��-lCy�㻆w���=,�h�	z�i����/�O�>x<7ü��8_���[9(fY�a��@�L�`㪎p�a�����Ç<^�t$�Oc�#�3U#+b��U.�W�Q�؂r��"Yӏ����9�Ģer׀�
>��C+Urg��F���^|�H��Pgc#`3e�VsP;�o��>#Ó�	A{Τ|{��"y���e��'�Oн�C2wA�����i�]w1i�iE�g��,��+�.���2a�K��%H����=�!3=��+���{���Jj�؟8�W�q׭���\;p��H}3r�-xh�p�n�o�7sܽ��^O��O�"��-��uݢ����<r=��@��[&=$믕j��g��b���E����A<�ޘ��hf�)�#_8�y��ՆO��V�@^��~�.��8����}1e�VW��I>XB��@?��L�}���~�z���f��y�N�����L�F>���idZ��w�t�k��|=^4�V���(���5�nJ�
��ة�]�nR&Q"��:
Z��,�Р�fھ�i�%�ld��AV�K��[w�vw�"|���	��� p�R��n��y����N晳���mǳM�a�P_^����ua�t�AƘ��ցM>׍{��v�|��	Mw�g�sP���� c
F3���зf���0���J;����]�1����o1 ���H��֧�A8�� ��#�H�~��5W���M�d�[qۇ�n�=����m�@���c��Q�C���v�k�8��]D���H����s�\Sn���է��M�H��ê1���q��G|z�C�췭���������"_r�i&wb?�2�k�J�*M�Z�O�*y��}!�>5��Ӎh9H/����b�b"h�&��(j.YK��E�b�`�0g���-4;"�<n;z����V����9��gOCI�v%��^��-4o�su=��%��gwֶ�_� ml�<˘�sB���Sg%a�����w��_�ZusX7;I��3����CX�@UR3\
wv֞
�/�%�Y'N�ƈwu!�0�C�y�mu���� �B�(��q~6�e��W�#�T�i]9l�P_�����{��_L�n.{(4vs/���
�Bki����.�� Z�����?����(����������u�|`�e<o�$��e��c�v
6M�K����|�.��63J7��y� N��ul��Ml�o�#�7�bѽ��M�K��ʿd*�3'��搼}��3W�hTVn�%�Ei�sd9�=�~��x�< �oG��{� eT�q�[��έi�׍s����W.J6<�&�kZ���,���I�i�a�����E]m�p���;0	�v`��}6�^׶s>�����J�e���Wu{�=߭��W�p� �����ݞN�������6�s��p!��'/�mG��{1i8;Xps��}��UŴ
Q��`��}�\�wO�^E1����A����QG3��8�[����Z�!��i�O�9��Tw>5�8s�8���U����F���OSL)�IsUQ�H�;}&}�����O�!T�OQ�v|`v��>F�V�L&B�{Z��-iܣ����|����D0~�x@�*�W��熾���X�ԯH��8t�6�;�\&��ۊ�&��%Sy�Ɵ��[����oW����ߣ'HΪ/������<����8W���	N��o�ϲ9i���}EM��r��n�7@-�ldW>���^�1e����� ��]�s{96�Tebޮ|{�Lx�>��	n��P�7*Jt�[��1���94����z��%��2:!{��cKm<�������Ɯ#���F#2��Ւm
���X$����P��C�t
<kl�n���aЃ�ƙ�����.��L�ܕdDfgV�W�e
dyVKڳ��r�i��T&��Du�h\�z���NvI��]l�8�XJ�fM�fvJ\t��]��y�Dlo+���Du��2�(M�ki��y�;<pv�KSכ� ��t�ywhU�׫��&��s5}���]�w���o%Im���S/5�U����{��Hw�]:�&�V_)m���󩕩�:bwAq�b>�}Q���M2�52�nE�T��)Kx�^�B�:�]%�@�e�6�bl��9{�u���)L��-�}oT�5bY.f�5G���idȫ�N4�(Z8v�y�ٰf��cP�L�!{�z,%�#�X��v��U�5h�-��+SAd������1���D��7��wS���ƭ
���y\�se^8�r{S)ޙ۪�%�!�u*	H��CpT���N�=%�O&WK��y�K�l��,l��_v��;��s@\*�/�U��V_Szz�[��Ƕ(`xIB���+g�hr��2�S�U��U�F�}ӟ"D��C	��os��z��cϵ��YE¸ECF��P·]��+`���0Y���}�#|u�r�Z�fiՕkO&��4�|$O6����FQ�鴠�ZR��^��h�i��I�0��ʽ�\H���@��J�u��{=�tud
*>�*6�
�u3QQ�%��Y���ΌN8�iU>,~���j�g/u�_�6o�,�j���o,e�S��W�wt�/��5l���b������gn���wU���+��M��Z���f�T�]at����7�S��b�#Zb���H���� ����e��3_Z�JSuU��=��eZ7� �����%cf����1Nk3��y_N�LY��BlK�Dޜq����q��upn��EB�LY�vZ�&И�*�K�*t�I����Bwd�
��&�Z|u�c�b���=����J�v˾ ��hgQބ#]�8�p椦�{��c��R<`��l�Y�ҍT����mf앛'\q���.7�Ύa�h�w�Y��8��Y���kc�;�N��q��O0��E�\�BG�p嬨eG�v~��$�bvө,�DGQ�Q2�*�WgE��&�g]nwtn����wtT�鴩�f�=Rhb�J�a�5�hs�θÐ>siS6����;��TV�:��4�n�k˰��]Qfݜ<XQ�{wD�#)�s���fv	u.R�_]*9����yc�M�����\&��i���΋�qUݶr�6���mQ��s�p�9՜���Њ�g7~�#ʮ�N�+7c.4;4p|�T�]JYůo�,u���<g�?{�
(�f��Y�Y����H���G�Ufnzg�>u��u��뮺����}��o����Ǐ}�;��IEBE�du�gH�����ߝ��rQPQ� �HGv��s�{��w�����|��:뮺�n����}��<x���{��Ya	4T���շ6�H�;r�'c�rӜEP�w�BHH�^۠$␤�npD�C����K���jRڐ��n��h���B��'m�m��vQͪΑ�㨢Y�[YǛ��=�8q�@�%Ŷ�˳�(�(��J3NI��N"��("�֊K��q�l�rQwZ�j�t���b�6��mXeXE���C�\!M�MZ�۸�����&�gig	6ЛnF��m��G9kV�q.�P���D�"ppe�tә�z�O���%�u�Q!�R�oq�k8�
	�BH�t��}a���=�*�܊���/IŌ��Gy����s�5�� !δ�;X%ے��ᬶ�k=�oy�O�Y��A1�<x���3J~2�9��!���� �Zp,6��r��8W0�9(����7s�wo�2�WP��MOet��j�bs��V;��G�:m��[Kצ���=۲�������݆u��Qr�ut��5wo�Vo?~d~�9D���G�������|�[{�B�ٖ���;��[n��t�ˮ�~��{k�UzK
�-���٬��=��/��at��4O��	Q��m4e�v,�`�݌1�iә�r��1)�I�3��w�f
<����{�v���Mn��8��7���m�M�@���;2�ДEC��W���B��,������gw���s�O��_�N����S��ȶ��}@��Q��IS�P��#�v�,z�ϳ��I5�1����F��%s�v��߼� *��ݯ�3���z]r87�����cZ聵[��ۄ���ǸRέ>x]�5B�-<�^�
�s�m��~������7S��7ᓭ�5Wm_Xe��AW�J�^h�i�o	Ɋ��yg��=c�4��Ay��W�w�<H��[L��y�@e��@��w��u�P�; 3-��w�:�}Ĕ��O>��x�9�`IWn�t�S����[/>��	��6L1�$X.#�w�F>��,鮊����,$J��Q�O��_���KnD�k�71��� �^oo�{���z=�����Ӽ�\���tAj�� �P�T|�_>
��m�O��oV��Ol�
u�+����8��f|����)s��ԓy����>��k�Khr����;�K�ǽ>=�����B�=��M�J�Hg0�Q���F�Ӟ[kbu�K�{`��
��G'��8e4��'��us/EŸV7������,�Q�Ί}o��-�0�v��Q��rT<���_�T�~��)�=C::J�i�M�����9�9@ܟw��d�=�|n,�c�,hLxs���JY�)1�ꦮ�J�B�y�[���5�w���W��W��/q����.o�M=�e|�\�O7�h��/G��q��B�)�~�>��P�9�˝cOƗx�.����6	 ����T�ӱ�uV��/8�CV�Ȗ�3^6���J�O~=	=�ߺ�@[�`Tl/�Cd0gB�d%@��I��a�$,�TC5�g`���(�U�hig�|�jT=T��F�X/A��d��V�]�]-���$`�'A���5w�q�K|�r;|��/�����hx�H�5C�н<����?��jQ9�؍�l����g:Tw�w��{u+chb꜖k�2��4!�4vt�.�������vq46��?�
��IL����n�.�V̩�<7ͨ�9RT���gu���Z���s�3foW4d���d�+	�.����D�<q��/�������;�N�J�����&g\u�M*�k,��0�T�M�2^7�}�E���:�	)/�O�! s��V"������ʶ�v�n�	<l��QJ槝��ٓն[��}��!>�N�P�^ǖt;O^��/�\��z��~�`|��j�sm��OS��܏N���'z�!CT�qmΚ����-3]P�,=0χ��~_Y��c��Χ�u�������1'dp� pn�]XÚ�v�͋��c�;{���x[5_%G�q�yj���׈�?ȿ0����J��<�h�����_�g�0�{�v�����VhL�6�����3hN"XE�xf���M��N)(��{�@��{�R���F+܇�U��s*ΌRo��7�E�s�=���?���@�A����4A�7
~�n�:������m(�� �ݨn�8t�]ⶹ���xz�DǠ'�>��5���rT8�齃�w���*��Ƙ��xp�Զ]��3��k���uk�yN'm>�a�@� ��'�߼&c�\ނ��3P�5�O���0Ҳ ��R��=��Ai�riK���PJ��|�%�o:��waߙ�f�i�&��[�>��^d\�V��V-ad���F/���]���
�?��ľ[F��:I*:�a�.�Q8�P����(�K���r�V��J�j!w]΍��dN[�a̺�x�r1��k>o+xF�u�|z���[�y:���|��/on<Tg��xa����Z���]پ������*%��*��䀲G7K�\�������Rxw�k� ��~������'{_��Y�8׎���}��8yL�i���!��2y�=��Fsm\44���xon^���s��A>Dо!���>^��	p5�}jEu bK�����{H����͊�-�u���y5vbM��`�Z�A��΢
>'�N h}�|l�"�fJN��TD�KUd��՗Kn����>��m|h}8�438�l-(����^i1��swY�_j.韻��6��ڣ��[���(�%ɤ%���9��t�����x-�����1[�i���s� 
6.��� ����?���*Xݔ�txpc��>��y��l�gQ���@��g��5o!��n��X���(_&�|�r��?({��4;���^M�'o{�+u�i���www���q��^��`�Q�UJ|vǶ����Hޞ����p�qʩߠ��i�+������y�%�*\[cX%ty�\��;9z��[�C�hen�Tl8��}3z��Ϧ��,�
������=}�Y9���>g��YTX�����z���T;I��.�r^�˯^��3A.������[S�U�t��f.T�@g1�,�/��!�3�V����]r�*d����E��Iћd?{������{���?���������IO�q�ɽ��A^O���gv��+�'<Ǐ��[^�s�P�|@r�9�h֓���Bn�\)�~�R9GOs�}�o��� �7�C�G?s��q���Dd�CL*�܍��T]������H�eW7`e~��݀5H�z�Sy��Y�C�-���a��4�Q�ȵ���C�:��HA<0vW�jr`��QL'�c�s�Ny�DIs�Jewc�c�i��p�"���`����Li@�@�s
�rQyjY��{��-M��\�*���l�ކø����4ƻ7�v�t��caxhO�*A�rJqv�0̆0��w(�;�Z��ptH+:X��b�|t�@����z`ct�1U�������W�\:��G�7���{�&om]�������Г�_T}��������#�W�U�(,�RQ���T�����c`���heu (v����-�P6��k�*�RhQ퐚��a�N�fq�@r���93}����c�G�}�ˌ��9hm��x��|��C��Д�")�
gN�G��V �+�:���1�ln�jV��v�:�j��{�`�Sf��{WEyڀ�u�Uw�,6�Sr4��e�����8p]<8(�&��iȴ�	���+̌��(�seQ���i���2���BQ��+\�{u_7�G��OŦ�zߦ����=:��Bx�ǀ 3x{�y���>�q;����T���D<��!�Ml��qL��	}� �(v���y��^fb�~��;[�᫽����'>�Bo�@P��Q�j���S=�i>BW��.^����$�t�a;:�9��tq����6�=C�\	g�,Bas���.i=ˈ2+}B�"t,G�u��K�+ks)Һܮ�~Ѓ&�]���� �����P�E?���y�fAvy�NI�ۙ�����U��k��pE	Mm�F7_)�g�P�c1�ޭᦞ�h[^c�[�Gv3szo��| �����ٝj}� &�%������GwP��l�={^�������3�+{j���d���ӑ��Ssȳ�G���u�e��`q�Kz����+���̮Ჷ�z�'p
[�9�=m��@�ށr=0�[L8p�9�'�9T�~�|�s��cv��s�Ӻz�w��}+ڼ�����M�G��Dsm	c� ���_X��<Г���×�*����{u�%�='�����V9M�Z��%������Ǧ=i��b�>���~i_b?���ч=�r����`�;��nU���m�-��+'�u�m���[Ҋ����ٷEn^R��~����ng�m�y=���u���K@xy�A���R���+^�J)1�jK������8�v�)U�h 9�~pp���.0Rx�ǁJ�.��{����߿F%���֫�L�c$��	^�� b�c%RS&�6;�	B��C�%)�=>�R������~�K߻`Y��I1�axH+����+�������}���8������P��*�Ez@���	=����@UR3^�nlٚ �r���Xj>|�Z� C����D������׳�4��3ʹ@�c�|��ѳtJ@̵s�n{��5�v��3oz�Fz��"�8Z��,�����t����T�~��p���5�d6ȿT�^��/��l�}ΰ���J�G؀i1എ���6|��t��`�Ns (�̠_��� G^�c�rt_�?ų�6�U;o�A���a��Agn�C�g=K�zڒ	�5{�	u��M�:���q0�$İ��V�.��ȴ增��Ö�C�dWg&շw[U>	��ٻ�kN�U=��K�9�S�G���Ê��^(�ܺ)����e��9�uY^�"NAw:Y����z{��n�V�I�>j��}Q��O ,���s��>�Nk�#<���k��r�0�c����E�<�N�:J�xO�ס�4t�������q���Q-����4ݛ_�{�z�ى⊬�nF�9�Y����)��9~�gs���l�V�۸/�&^���M����
�ۛZh�"���h�*�5��g.Bus�#�$�6��<"�;݇N��{VΕUY�1��GY2��c3R��S-\#����Ώ�C��ˏI��"	H!C�7ڌ+޳�����E�<�{w�xH�Ο����z�}#E{fV�?G7tgK�\ 62�����7�n�@�=�>��f�{� ޠ���&>g�����D��s���Z�W�Fo�Z�{;��N;j�w>�L�����O0M~���x�a#���G0�SmY�);�+t��Huޘ�&�ƥ��-��� �sã���hv%��s1l���3!n�va�j����&=/��=�}�n�
����K$st��\��L��x׊�e�vi�\��6�W��c�&D��u��SM&��3���O<����~N���r�y�Τ	�
�>�:H3�aB�@#�˟:�X{�z��4�̡�a��ݮ�U�����y��f���Ͻ�:}zI/z��7���BBLXlnO��}j{ͯf.97}}gti�J�o�W�7~�o
�怵�IAi�_�XH<L���E�.x��߭oyR�14���^�љxl�ٙ��e�
��IC ɒvk�08"��׶s�!��D*�W.�w�m��3`�#��^���Z�c��vl�Txk]on��c/+��"���j�ӡ�۝����o2�jl�0�-��[����`�̮�����+� q��`�!*v�3˯��T�xt26�N�i��=j������㼧y�ne7�,~�~s98���D P�P�O�{�}�ǟ}�o�>��IH�q�a�?�Pj������H6hM�#�.�!�ǔ�&֠9��xV��fJ�w�co5i��7��u�L![��W-�JtX��O|�/������<�!���[�5�P�N�}3�������,���"Uc�����Wj��폶�c��(oGs���s���ր������}��G=���U秝<\t׫'��]D� ���~�?-a���ۆSO�h��m�UAm�e����iO�co�zCtt���1��\<�S�?M��H�~�^_s*_�R����3�u���ɩ�zu�|Q<�~�T:���oszv`�$S�����}�1�ΐ�,��w+��!�A�M�7��D�=\݁�n�c"�}�H�)`��Sߝ��O�ɸ�y�ssڷ_���OS>�O��}���6N٨iܩ<�<�txG����M*�`0���WC��cw�im3x���	/'�Fx!��(ؙ� 煩h�s
9>�z�9[���2\_=��Ɗ�][	�
�=�.چ���q�U��1��r�x�Uȧ��>�sk{[����L���,����|k�1�cM�q� �M�H�vU���KM�.^L��}4�[�>���j��}��{t0��e�@K�	|�Ǝ���쪘D�m�!q��������\.�h�xZ5�e�!��h�=�>��<����H� ���W�{|����a�o�U`u��B{mi �;�P ����"������.1}��4"^��Uo���4sa��D�q\��{��<�X#Q��b��ƌDy���3��x_�^�⍔A+�v~�ӸUO���f���i��M��3���՗ɲ$sD���Tم��D��0<!��kZ'u`�M���d���s���3-z	@��E2�j���2�ݲ�ڪ��76�����J%шx�`{�A��@�ׇ=}���
]�j�P�e���Ii|U��i$�v��ӯ�ʀ��àO!�o�L�Pݫ/�m�}��^���MYsk�{_sv��$`�J��.6׍oyS���XHc�{�'ܯ���r;i���̿l��⃼�jím����~�2�
�R�}+6i��\�C���ŵ�t�x�}xc3�W{�IO��VH�07H�l���n��p�_>=}�_k�Ur�ZfJ�9�)@�߽�f�=�ӧ�maxFzA5��n�խ`<�)�%��;�0��B�F�c���(�xs�ć�����k��$��t�j�P�}9X��`:�D/xU��#�*��C�O<9�I����IM�hk��ͳc4F���d�-�-��շ�⺃f`��vT���⛈�s	�]C�D�I���`�:�uR�խ�R��@M���Q��^��b��{��yF���.%' ���&�%�VL.�����	�Zx&�ztzڻ�Fڼ�kT���5�.,��L�`���/�2�%�v�'ԗc�؂�[*[鉱��(�kB'�`�bT�j�KcrК��J��Dcq��n�&ӫ��j�+7��d�G�,���`�P�b����iQ����\	K�Pm4�&����B�B���lu�=q�Χͪ*G��n��/���5D�*�)�n����l�c2u�<����jKL��s ���X蔱��qA�X&�����f��\"�e����_�uTG�-E�b��}��F�X��d:t�.V�8��O����k����f�e�lۧ(��S͖rv�JOuK6�8�H_9ԯ*>���Д,q�k7�3U���W�Ŗa��X��%�+%�R�*�>����+�eC�h]XOC����M����P�[v/m���ARP�ŔE5u��ya i�X�{�Tv%\�o'�[߲�<�����:u�֎}Ԥn8�j9��Վ�T/;��
����~��DY�/�amh�2ʓ]�MRT(ITH����Q�ۊM��QQ�t��X(�$}��j�='X���nZN�o{��zc7n��':�R��a�c�ukh������e�mz�ٲ��k���YS��N����|�5�L�W��}���y"���xc��-2�	�I��&t{[Թ�)��[{>j��m7���ۆ>��Ƹj��Y�w�WE��j�Ă�K��!WnGB*s��|�
�i����[r#�f�Ӄ��e44Q,�ܰ��b�onv�˱=�[�8h�p�F���7M�+)��޻�T���.���6�M������R�ia�Nj8�׍\����[~�B4�k�r����{]�j�[c5�ot�m�s�h�=�����08��L�w]㖪S42t�>#�R2��e��i�T����6��g0�2�?su�v���Tya���p]�=6�ʑnՃ|������2��;"n�M[u��E'��Us�YJ��2�c�bt"L9nL�|Ζy��Ա��_ٛ5νt�%I�}��bѓ��]Vs\�j�Q��ͬ�.��KlO��*`:�����M�K��ΝC�E�+n�<��A�l���Y��Cw��ErT�x̟r��<�V^u䇮r�yr
�}��V᜝>�"I�6K(��*�����[z&����9֖S��j�OJ2�vA��C�?]���ΈvAd�"�������zQ�y�AE�Bm���ǏOO�]u�î�㮺뮺��뮿/�������$((���)��v�36�B����r�cJEDɓ�zg�OO�����|:뮼u�]u�ˮ�����zzz}�=��eFXfdeT�]��$E�-��ι�m[Z���@�;�r@a�Y͒N��#�r�X�$I!=����%8㎜�@s�����Q"����ى��{۞ҽӻs����/�n܏k>���K�|��-(��(̮V�P�۳�D\�wtY�a�М�v�$N��gZ�HDGq�m�%~�Q�]��lVG"$8Rf�qI�6�63l��n�aI$�Z�����DR\wyږsY�D� ��8\GNH��p�u�~�}��88��+�������|����%l�#���%$�!E��ZP�ē
C0�#�'�j���׊�g/��l*���ê�"dMm`���%9���/�j뷹LËy��靍.��7�b�)^'9	�pB-�e�[e��PC��e� p����P##l�#nF	�a�Ȝ��51�!)`�Q2�i�ԑF�p(dr�d�y�ts��̎p������*SE���UiQ�P�w�~Ӿ�)�j��;��@�ӽDTZ���Ř%��m�~��~�X��/_��s�`!'zI��~�Q-��^[��\�! V�|����Zp�qa�>��Wq��cP��k����~�݃�{>o$�'�kvW���]�O���Nc���n�n��@�P��S�@r�K��S��^���ٳ"Wu�Ss�^ՙ�^�9�^��g��^���	�3��q-F0�������<7;��e7��6��յ��6������o�ɦ)�4�]B�%ԥ�ݑ��C��/]�O�Ӿ㇮|\>mn9|�K�����h`��8|�T&�4��ȖRdְ%Gk�C�uN8U#(l[���09z��k���j���F����M�OmAZ��@d����m)���o�������!�*ֱ3����5P(��	^a>x?|��ߐ��v�3]��'����#x��(O�]�<����Z��f������&ۀk��RU��zC/|�z_ɞ�{G`=���D�sa�r�݃�VV�Sn��\�q���F|�Z��魮�S�a�Zm�~+o�~���ܩ+��I5b��f t��/�҅)�$�F�;#++&���y._J;�IT=����?%�a����}�����e�Ue�J�{DRjJ����1��vJ���{k*���Q��ݹ����u�A�j���G�i�X��U�O�ۏ�<q� P�0 ��#Yk��2}ُ��=��"�g�H��!v���ǣ��Qz���yg�顩�Wm[ۻ}�u`�Ü��ۘ�k�KP��Bˠܺ)�d��P���{j�<$��ƞ�;*v���^�0�q��D5Ǥ�������G5#�_D���S���fk�=*�7ێ4�2���D�<5���|l{T�X��X���A8Iờ�͛H�1��i���Mu���'�A�Ơ^���[��
s�qp��� h��Z��,ވ����6u����m���άwH�[����l��aȸ~/���Q~fi�"a�n���V��]*����--A���;�8��0��G� tގe��Ewt��Q���^��k����P�96p \K�5Zt��}0Cl�p#�v��n9`�����g���8���sL$�sz#7���D��u�Q���y�h����#L�*\9Y�P���S^Y#���t�>;�Η�A��0��W���;��M��>΁��y��:b�'�;>��*7�l�ZɎ�v<��Ao)y+M��/sv��SV�Fv�ů�7�|7�('W���;{k;���,��W/�JZ6�,3���]�9���=U��0{�|��M����$��n�yM�	5ȍ�w�&w�;a� ��B�'A�1�i�NQ8ӳ�6	.��;��<;����'�xL�Q �"I3�gAu��p�3;3��&A�b��v�H�xBjK�|���E�����}Bݘ��q���[DdT;BO���-[e?{y��1��g5e�A�91�p�SC�Ҏ�'��v�gb��e��Ȼ�1�si��E����S@[IQdƝ6'��#)���
S
v���G�Xw{����zq�Ldhd��9jg̈́�'���Z|�38"��׳�`C���h Ҥ�����#�������?uSTn�c�ly�e^;):��d�_;�g.�ǈ�ǭ�$�3���j7`�vC[���ķ�)�b���
�zƇu�g�D�������(7v�y���>y�a�a{�9Q��Ƞ����Ͷ��=��X���~��1�v��+	�8�=�J�����&�*P����:C�X&�ó���m�]�C6�OnF"��U9�Z�������9������^~�}���" �/T�T-t���#�z���ݽn��5Ѫ�IS�Q��{��X��[��:oD���w*�(�3�&��{[:yu��T�����I_�y�.�ҟ�aG���F��{�.mh�ӭu�	�qF��Z�X��+�|������}��K�׹����R�����.ᙦ�i��޲�+��ӫ���w[.�޾�s�қ��s���DVJ�v�"�7��c����|���'�xA#Iy�f\r\^ym���/��DO��ڸ�!�0Ȓe/_3�e����Es�7��\�;��d��\Ӆ�ni��u���fpy�k��#5Ah3콌���t�n��\s23��ڣ:���n����̣��k����q u0�<��!��K��I�r���^Y�_s�O�N�L;n���'1���t�z�����3�uXH��!x�lx�>^�>��׺F��4�e⢳0�V�]8�JS�f��_}��'��ӆ���I�@��N�	�k��=E{h���L+O�yW~�p����J�bJqA#<^��	=��A`�<:i-Ѭ���S8����qS�wٞ��+c �./t�0��'W.
�`ZF�yu������P(еQ�,�`&���I��'fk��N�f�1A����_X���VI��^�ֈ���ʂP̵��@��࡞�m8N�u��U������/�Ǟ�0�P|�O�|���ϽlS�l~k�xJ���==:+�i���޾�v����Ơ^-ᮽ�	_��
�C����EV�еfpsz}� >w�.麻\1Cߗt��&��T0S����!3S���l��@5��ы�[[�v��z��_W`��W
)c<S+mwt܃��t6����s�MU��$�],�(>w�k���qɜ�ԕ�\�wA����i�ei�Z/F�{�x�z|��	��	)-JA�ߝ��oXl'�������ov��tckv�7�|�����v��.��W#�U污�CR�֩��VXzC�Hg�@��|�{s�{a�{۱�o�T��{ٷ[�@H��{���T��6-���U�,��5����i�,��w��rل�n�ȧ�on�Po6�MV��n�|�W=�,�A�{i��in7�\>��B�İ��vМ�ń5p�Ty��ӭA��� �'�{>��Ra�~���}��7���\U��QU�/쫞���YE��'|B��5f��c�VAF}�ve'X(�M�M�=�L�	������ˁF��9�.)�����[�0Ƹ}��dt��}⌌Q�m�N^5Tf��B;��t�ë�y��bYPXhu}����T_�����O��k���uR���gc��d�8�L�%�[�|~|�my�4���;�)8_5�=l�g�v���Ss���������У*ccN��a+�Z����k�o�� ��8�|�U�Am}����bi�$�W��y��23�c�ڼ�=��?�,$���9BOt�:�*���:�T/:7�gMzkoh���8�;�8��j��yJs�WE��;���U��7���� 2Ȭ[FB���6�d&x����&��x�jz��7�plz
������:ku�#���ۇʽ�Q�]�4gN�f���p�	���'�P�@�A)҆o ����i�KI]LN����X�}�_|�F׌�S���Փ�2��疥�yJ|gI���f,飌	��U����~�>`��PP`~�@���D|��M���� ؟}�:o����<����G���e{��`tt��h���������Pz�o���c[:��v�J���Q���̖�\�)K�l��y�'"Y�p�H��X�W��v����7��������u�4�=�A�MHA}w�R�0uB�����!���f�w{G&��B��ތ�0�~s�zm��]��L$nC��g9�ؑ�i�b�s7��ñ�q�N�ŵ���"�Ҟ�%�>q���]�g�sW��y��PW��n�v/V��������%����~��%��@��v�����$'���3�O�hn]vl����?��M��q��|��=�eyAJ҃�+�O�.�~!��&K>3�\�dÑ��̜�f���~�7s�u��;�g����ڙ���p�F<�i�"�n�wJ��ktUe�h�;�!��+��d�⮰SѸUi׈\�..,> ��e�#�(-o^�Zݫ���ti��b��}�*����9B����jT���@UV�9k�����kq�7rM��3�ޗG#�l�yz�]���OO�P�8𑂁�) I)�hZ	
_^����߾{��f,����cXt��%U���9�Xc"��u&���bz|�<l[n�Kn��-[�b�,���Ʀ�6���ژirt�	=s�[��F%�i���j��/^29��� n�4o�a����qp�ϯRb[hnu
����
Y#�����6s��:m�ܶ��	���M0R��D{�c`!n��~;�a��c��N�k�es���Q���۰FR���9��kH�����=Q�j��I��|j��<x�a��\�o���n_�ࡍi�G����.ǎn׿r3�3�%���6�#��4�@���y!{3���R��g[Fe$s���w�%s�a9�`S<��O{P�G�|US�6/��#XX���{��Vr�Qѵ�Ϸ01��c����1)�v�jP���S9�:�[�FEn�N�Æ��9���S�KW?nG�]ѡ7e'\�i�.ѫC�
��S�kwv:N�mO���2����0k���>�X}k�؜&�3�~C._P�~x����+�6֏ρ��=�/c���r�Z��j��ô�����*��j�˥�������p]�������>�W�l��o6���|�<Ugz
|1�呴{p�������룲���x����nA����'��K3���gQ������x��@�����N���v��C|x�i��c�P-��ꤘ>`��`{���z�����]r���g���u��_[���=��C���:�|�З5�`����	��g/�ǱތSoEV޼�/�'
8;Ku�{�\���`���B���&��Ư�>��[�<m�K�S�F��zk1{�1��� m�mj��s$��Q<�c�P��t�8���a;�ml}�A�&N�i�T��4��D9��X��n�O7�7O��bcg=��5l�榇h�=��i����G[�
�-�.��������+/c=����%�}��kB\���e�6���r;�#u�F�$�C�z���`	���|���~cm����*�u�tہ0y5:c"X��ז�z�K�t&U�=L�<�A�[}g�C(�t��ߕE1�`�8�����.3ekbR�lp����.�.�a��W��;���.�`�����r�ped�h\B��Z�Ĭ?H=5��C��y���{�k��ea�V�1��if�?|[ngן=��������f&7n���匀��3-)�K~�kS���7�P��`ͶJ��䩰mQ���tn�آ��f7��u�.�P���5�r&:�]��]��XW{$�3s�E&[۽����y����<����5� #���.~���=�ox30k�z�X�QuB4Dv>�>7)T�ur��pU�9m朎k��	�h�v���c#��.����ٹ�@�18�8�A*�l�r��'V�۪��׾�T�@J�ax/���o:*�u]���6�>{�l�s
&%=�^�ܙ��(�����I��b��C S9y����Ϡ�����dPt���Gn�&߉hۥ�)�ml�<N�
@?Pi��O��*&v�X%�MW<~B��&qk�i~��c���S���9,����.5<5z�7��\�p�{5��g��+���Ö�z��L �tEhׄ�+z�V��c��z�M�`S]��B��zqzǽ=�-���;���#Ȑrk�Y���ܬ�:y�p�`��|~jb��}^&sU��Wʅs��ym�U���^v�W���Uz�	��>��0��H����q�����ӭO�Jd�9���L9���8kvM�nN�7c8m�j�d�'��?:�I�$0Mry������4w�߫��w?L;2�mj������4lږ�������{��(/���q]Ǫ� ��#�.��ep������n{�L��0v�[��������|C�/7.�i!���4�q��D�ފ�ARQ-Fʼ/�$�퍐H$H���$�{�ߤ��yvǦ����yU��yygD˩uc�c\�:�����ڗ�9����{z�͘��IM�����T��_����������wI]k�N����R~a<�T�~�QM�7U�[��p����8��Ht#��z�&9�r�;���\=�D��P�N)2�=s�=ЙW�r��q-`>���:�\���n��õ8����:n��}�1�5�p����K�K��n��K��`!=��۟<@���ًi�K�{�;|a����G|�߬H!�u��bz9>�:z��~����nln�y�pr�{\'�-���;�.  �<����D�ԭt~���2�<���>��<�v�=�T��Z��2�k@֐��� ���/|��-���v	py>`��r��.��Śjn�9��x���po	�G�^"m�XX!�5��8:a��p��]�r]O+|����F��Z߭�>d1�,�`��Ͼ)�)*v)��o��v�tFĳ�p�]+-Z��Û�pgY��k,~��z̏UJ����vg�r�f�)	s�����3J��w�U]���w}�^���4:0���[�[b>=Td�߽���WM���W!���!���F�ެSQ,�T�ys��.0z�Z2exﺀ�k�n��s��.�!��IMo�V���Ys �k�� ��`�MM�Ř%�d�ևќ)���@wR5ݍU]��w>�˘9�Y��PU0�x���[�Jծ*ef:��vJ�1�w�1YR+u�S��˕F��3�]nlk��]fa��1�W���L��)c΁t�Sy[�c�ie�k�	��@:�T���!�jo�N�U�riƓ�6vb��;��>����l��*%u3N�-�{��yR���p��M�.��T��C�VwL�V��h3z:����}��v&�R�f���;*e�i�ŭ	#����F�UE�#D��^:j�ɒ�%��f��.k9��Jq�_j�����H�rxw.4��/w:��o#�ya�:�j<�V:�]+r�e ;�+�b䈣�PX$�5�*�s��w>�����6�v���뷌t��O)b=������5h��^�5�@�lط]��1�I�]��j��x�kVF<�b�U<[�&uJ`�zp���Ɏ���*!T�_�&�VlS�&
��̷�7�OU�1�@ia��^�T�zU����ywL��)��X$�7S��5���T*�wQ������Ȟw`,8�S��=�J|�a��A�7)��B�O-vj���ٸ�2���*�N�D+�i%]?�E����$7q���śޥ&l��r�+��0EsF1�;kP�gA!�
U��ϑTw�%�a�!ϣ�����Б�e*�Bx��,(~�>��!�<�����<�ڨ��/r�ss/V�Ru���7MѺ��띱�b7��z�Eٶ	ie���P.*0!a��H�S(��I��7O=�x����-s�9̈m�m�[���p�^J�t])�H��&%]6��JK̎@x+�MԶhM��|vP�B�yҦ�۠�(�����sv�y�Ur�Jz��ib���W!9-�y�Rh�;��W�-f�zQ�go;�n���U;�Y8oBl\�#Q�Jn˷ùR�ON�ZB���iVWiݎ�e�Ԅ兎�re�]І�s�i�m�!F�����B�R��:���a8C��-��k	3L����opt�qsA�N�F�<͇;y'˯�l3Ka�Pj��v`�h��8	ŝ���ʵ@h��G�m��%�1Ы���}��w��h;;�mv�����h|4<�Pڝ�v�/x�&Çr�����|����Z�O�鴺��Tv��3�YE�|��'gj�L`8�Vb{S.�.��,�4`����<ڊ>��jV�wy���>o���o2Ly2��,�{�`��ݟM��4�u8�>秵�W1wF�zJO�P㘢�ǻ]�J⎗ÉFL9�ڮpQ���������������"���'���4'����]�J9D��XXpweF�mm����v������_O����]u㮺뮾]u�u���zz}�=�@PQrdTz�h���<&�\"����QYS^Ǐ�_��u��]uק]u�_�뎺���zz}�{{.H��De�u�=��f:�
�n7W����I��m[�	Kk8;mrgr_kq�v6Ȣ"�Z���]fM����}������9������t8	�ͨ-á�㎈�Ģ�f�Y++E�ed5��Nmm[۷�8<��j���vj^������맞��y�=�ݖ\۳��w%&vv]�	'v�3u�hI�c�lw���lj�����#�mYŕ�d�M�.�w��^�%glI2������BJ�`�)}�u���*���}K��|_{�����a�(RY�#5�]���{��,�D�j�G��bv�dءU�YK���Nc���R���u��<x��D�"���&h�.M�;9ٞ����l�vE;Ň�a�;��+��*�Ϝo!<�h��^����۷νiΥ�L{��j3�+�f=[է�V���V"�l}�{�zq߫	|��V"��gf�&����w��-�������W(V=ŇNr���:�u����Ls��wH��\�F�^I[����������Q<��[��\���r����1�?�ۈ,'r�:q���3um�8t:���Y<8�Muw;'�]�dWP���y(��#�-n�>WNF�	�2��X�����~���mˁ	�o�ط'�%��=�7HM9��4dsF?d�<�h�����9]�;6����G��P��y�����	���R��n��J��=��t�c�%��'���#�&��+�&G��3� �ԏ���H&�P�X$��7<x��a��ƕ'�+�'���v�<��uϣ�U#+��#�8A��ς�P4~^�TX{Ly-�`����'{6P�ocF���Ѭ����R�����b �tssC��qZ��]}���:%����J��_$���'	vj�e�e��9n��&u�v���������e.��W�%�m9�4G�D]��d�3i,%9;��Cm�s%s3�����74�fo�
���W�3$n��{�ɼ�1���� �oW��8�L�8� ��~<���{�CRxf/�ޯ�E	܂�����%�9�MJ�!���?_;�Jy}��cۼGS;w�l�L�:���c�콡@����dҔ3Sx��[�=���S����۴C�2��)�H�S�n[ <4 ��c��*j��}�ʩ�>������d.x�������Ik�$�9�.��V�i�&�G����[���\zi媺p�2�3uJ�K���F���7Y(5���ɶ����K���a{������+F��Q��^Onv;��F5>5����!��ͳ�H��*/��{�1S��#��t/2lV��c��#w�7:~���o����nu�%|�WGJa-�#��@�{)����藨h��I�qm<r:�v7�c�g�`��#nkc�s$�D��r��Г�|�a`��-Ȝ�F�4v�V�op���9�8�C��O�|l� �����(����z����ɉ��ؒKi�p����PJ�3�N,�:<>zc^��͸��0���'�!5j�nN��8{L.'�l{&V\��&����W*o�\>n����z����6��8mj��5:����(�M�Ӵ}{17u�\��]٤S\�u��圻����4�q�{"����D�*X�V�d�f���[�C��G��{����{��R�`�]͐/��C�N��;���j���ȦXk7�A��U;͖��V;V�&k�ϛ�cN$�5���^��x?�75���/�fԉ6�6���׫��5�հ�iĮzk�]�_�3�К�T0�xw��]Q!����Ǎ�9_Y�Ƽg8;Oۛ�7��sޕ#�B��Iað�n��l�(A��I�hP>���M��/�k�&뷰�l;�.;<��= ���EQ(����/c��	=���,$-��-U�yu�h5s��i��IӬ���8!f�ol�}���e�.m�6�t�S��{�P'R�[
<%���\S��r<�gwx[c@W|2@^y��R����L�o�o�Y���g�9A�Gf3X���[~<��8�E7Q�l��.��� �꘮|a^��n��f�̵��@ތM�yI������@;~�*�}A|P�=6��)��@v�hP'��8��yY�~���ꨳt���vdK�w��]�/��~U��
�}\2�Z�ڃ)r�,9�w=�����#����Ֆ�;S�*k^ĸ���M��S_�[�C+Q�c�DG��Ȧ�_?y:�ɗ~��2���,��\1Hi;���u�J/4ә�x3LCf��*>c|�z�S�Ru^�-=�� �Pj�`�M���A ��T���+�8[y�����5]InV��\%W���ؐ�q'N1/ebH���w��e�M`;�'��|������7���W�8��� &���v��Z|n�_�+����/��b��O,���A�jr���M��٣{6߶�s�繁k�<5ٜ�!���� �}���������.�j^��2�(�f���BΡv#g1�^��Ȭ�z1ރk�?'�q��Y���>x����a�T>�ll�ݕz���-�����Ů�

�?,"�1q����n�]Jr��D���S�a���\���9?s����N��k�`5�ޛ��_�=:�	BP��gsw[��+�
�F�dOP9JH8��ג��-���=�O��������ďu/�n>��gهu���o1�[ZDp��	�O����JE/j�R���5�@�����yE�9��l��t��]�Y��x�)�{���֟CTĶuzdKv��a���/}Г�?n2��ՙ1y��rv6�!�ٙCb�p������-�N4qx�'���{��f7Rۧ�rd:ۃ�ue���S��I�϶��Go%`���;�uơ�ʀ�q�,pO��͕����T�z�h8�r+�{]�Uv~����q[���[)�^m�;�u,~�l�(�r�y-{�e�q���(@��w���d�nȵ��rs�]� <�i�uk7mI˒��+�<}H�L5����s��ئ��mB.�oa��=Ԇ~��>^q�������{V]�tG_~�.��!��(�X�Kig�x��x�b��v�cü �`����M�P���7gc3z�'��G2W��*�;I�)�g|Q�j�-���qប��hR�Ϲ�I��^�C���n��/V�ld����	��U!
���^=�e-��zg���=�d�{1����<{cKO�qi�?��
zl��,�ˢ�sKѼ�B5�9z�i�f�~ݜOC���)&,!e�^�@��A�d}��g�Ʋ8E^�`�y���H�q�M��zi?%�~����U��r�(xy��"�j��c[V�fѹNj3o{�p��f.Bq�(��{�i�纅P�8���?<�{w��s:qPS,(k]����j t0�pu��w;'�~#�[�M���jc$O�E���_v��C�G"�n30�ϊr$]ΰ5�qF\Q�U����u�H��wRc�f��zq���j���������C����Cӕ������gE�nN��������!�驉f���ں:��C�n���pDF�:4Nl���P=JC�ޚ���U�s�7���32�%uwV5^?C>��x�}���W�x\��o�Ϻ�s�/Jzigw�uoIO9�IV�̕,;z�Kwt9�������$a�G@uN�]g������������ս\�vm����Ji��i��p�� C��]�q|�ƁΡTrQy�-`�4�-�S���֛��w3�c<�����r=�Bxw����vA�[��T~;��j�A�3���Qr�Wo���h���cFTW��ݷ'ʯ�8��Pv��������a�T��d���[ek�M�<0��6"Nooc]�ȣ�(�a�^5�^�3ꠦu��������1�V�����bU�e�1n�;[�m�� ;k��̌��\��s4hR����.y�<�ţ��Q�kγ:���~�hp���|M���M�kxfF��|&��wINǪ� ��ܬ�F0��h�gx�v��f�?����:c��*Q�/���.�h=�I��k��gq��-�<�ZӜn�dG�ņ�w��S�&����Y�>�Xw^q3�����"ǔTy��}+�&�@��ɋ�N�c�=�a�w)7�m�+�j����`X^�]� �w�mF+��s<xiȶ�n���"�n��X�L�A��u���â��~T1�J����sf3�1od��"�`�^9�rv�⋳^=x�+S����	�tk�cf߰ ��O>���K��Y��h+�zb9�z]�[_;}��d�ʑ( ��\��g-{�-�<̦�W7�3�pV�-��9k:��~�/{�yy���d�w�
�⇳u��]��qMZ��+����K9ml�uvJ�6�����3�de��٦�0�!C�>�X���ȯ�a2�|�WGJa,��� �d:٭�a��*R��D����"9� ��u�^m�6�Z���y�vO��d'P����E���6²�OR�,����B�Kc롡�u�&��F��`<�|�iGa�cL��ބ�n�����(<x͗���i2 �X�|�m�ymF>��ϲ�3:(��Tk�22�l93�Y٩T ��QL���	�@�Fh�;�ׇzh��� �!��71~��E]L�Csg��p���N��
��X���s�	�=>�aC��m5�H��,��慔6�ͺ����#"�S_(N��9'�Z])��a��]S�5=��1.�A�}V6:*�Q_Kk������ <y�Ku���f�Eqx)Ƅ��{�t$��:����γ�e87G�I�t��֭ɩ�{)_����J��L�����V*K��4�wP6�����N�K�WN��8��7f�	����u�3􌀔0|���@x�����v�N�N�JU��{��^��x�v."�sQK�Lgb�Z����5��r�#j�c�Ξ�x�UtZR4�F����mo;'>��Ĺ�S����J�<����śE'�q���ajy�9���)2fR�;1���z�M1�����^^^��jp�՗�@b~a�u�4�"�jW�K��>`]�N5<��t���U��+}�5:�MWi�a:���s�W�1��� ��sx^�v�"-�O�i��@f}1<���x�B��Y��os�Դ�����]�F�qق��L�>=�o�����7o�Fb��^Y��@ؙ��R�t���.x`{�.��*.��TX��7�C"-]^JV8z͜ahÆcU�;�sh�M,�\�g���X�K�!=��wVO�t��FG7_)��2�-;��U2�����:rk�cݯG{53�/G�p`�f|�7���\�2�0��%4S�2�����w)X�n!�����h?{�.��ު����Z�L@��~O�}��b��CY臎���}ZNw�֦W<����i����3��k���9�.+�w1�^� ("#�c1
�NNAV��f�n���=�d7�p%C��4��_*�O�ץ��T��!J�MN��ޙV;�Qz]Q���}��׹�G1��_H�^9]$Re��/Ns���L��C��[���}�Y�,���\����1��2L�~�;����pZ�c�ޙS%�v]�_{xc�sh�hu4ٓtm���d�=L3£���y�T�����Xk����k2�ytuR\$����5���c�gs�h:�=��.�ñ�پ����?���i&�[ݥ���f�SeW����`�����|֑� ��B�.��Q��H�	ze�4UO�є�Uϳ�ޛ��gة_@y��ZD�5�0��mG}R}� �Gw}=�1��A�����E�5��C�^��F/�;�1��P��[�^*���R^YGeCu̡u���yl��O[u��\1����=^|���y�%�3��q���`<!�}���n6"_[c�w��9D��Q�p��\���z[K8��7�+�C�4����,i����v�Mef��tq��������!�U�v�~N�pcȥn�C�?���B�nUb�}���H��f��C�i	��1OR�oJ�Ey��ȋ��O*��j��cv:!tte����0pm�'��o>זx��--(o��|��ޟJ{jk�n������I]E�S��z�8r%ƙ�,:L>?����sϔ�e~�(,.����~�1q��`�z�����K��i��nHE��Ξ�W�<�;��
�z��O�\�^b�,8E��ڰx��Dn�!V�τ!G.�@e�+�"��2%�w��;m�|���Ц|-9f��2ﺤg_�ݮ��q�;J�BJ���>��_>YǕӷeRȇI��ﰝ��s���i8"�맷����\����ǪDf	Ҳj�߫��|j���y� {��Je.8�t'�i59��	D�s��SM�=�+���a{g�{w�$(�&��MaQtp�tc��00�W@"v������{u�����ܥ53xK $���΄7]��Vu��E��x/2I�;����I������':�*�O��2�Q��q����|��u��]C���$�IBq�p����K��w��~@�c�<<��7���N��j�	�m��M�nOA(�riw������{��sJ	�Ɓ�bXn�}�-y���F��P��}����9y~�O��g����;(�<��q@M����|wæU�C�ڀG�~�b��B�@��Q�͘d��v�Dt)��ƻ���a��W�~�J��DŻ��`�1a8K�k.�]f���ˮ�k�e�\�M�����,2�^5��F=$)�b�O�B�F�OW��2��|�̷;����ji���b�ؾ��d���ә�3��N�Nm�B��ُʲ�sw��+��D�%�&`��>� ��V؍���o�����T(�'f�'C�*xR-��Oi<����o%�
���Ǔ�|�.�� GI�ݖ�"�@��(2�Scn�eҁ��moro.�5 �a-\�כ}�T/8Du��繯���S�\����u���mQ�6�C���h��*��M�z�uu�a�z�1;#�c����C��Z��TZ���,��5�\s�d]�.oB͔��j�&��79>��ƞ0ow{�M����؝N iWmچ�sd{��a���1-�b\zg�����{���kI���V���z��xv��@�+w��u��T\�n����Z7H<&�#��Yc�HA���hڴ�e.J�!�p�>8>�is����]�Y�=�sv�ے嵦�]�c����:� !]��5-gn�ff�9��u˽%jLc�1�6Z�x9�#׃��h��˹�$�ҫs[��!�/(�g*�����"n"z_$c�S�ʷ���|/�N�X
3��(��dc���j�]NcpeY�	z�>5�)�I٣zuP�B�.pԧt�(�1lE�r�'����Ǯ�ڴr�	���$��Jl��\J���8b�5�k��r�n]��A�e��B;l1�tSL��0N�.sշ��Tՙ�a�5:�(d癎eÁ�ޝ�U�;J��δI���*�݁7�4��y��t]wpl��W!鷟Y9G[�Q�d�-ch��*�
BGLU&и��$�V�!�)��}�% Ύ�
�	}�jRn�IgV�(����G#�m�^쭍��;�o��]Ie��t�K�
�愖9�.")�v'��emE��\��RU�1�	yț��9|Q=Dh�@��E+��oA}K���s�a#1Q5%��
�nXPi�Tm�ˮNl����S1S�´�,�Xql���V�S�f�ǯ3+t߫��:SCs�j���'Z�R��,X�xNfMsW�4%aN^e&{��Ve�tƶe�F�{us�.=|���ܧ
W��/�"z�|uT{��I�{R��#�]�uT&A]
��l�]�\wkyv �.ic�G-�/4K_��m=ٞ��`b(K�#��7�`��-����8�s�!Y��q�{m�;Ϲ��yv�h�Aȫw���W ՚�X89w�W%&�=�J�s�Gr۝�By`r,���p��=y ���#��;;l�Eن�u�OΦ�A:����3��X�%!�,��L+�m�ř�i�';�-
�:�#� ��	�y�_���&�6�^]��ʻV2`����/iR�l���\ϲ�U�KwSI3��Ѧ�:A&��[�$��k��t`�/y�r���ued��<]�Mo��*r=��C�\���ݗJ������ � ��H��ۚĻkEqd��"ɵ�Eï=:�|:�u��뮺�Ӯ�믇]u�]zz}�=>��☯-Z�:;�;BA���ќ��[��3?O�G^Z��������|��o���뮽:뮺�u�]x�������|�w�SDMw.���:̎���J[ZFY�mҤ���:Ӧ����-3�m��o+s�������ok����{ۑ����Qҝ���H�RlݧEne_���>�z{�ͭ�6��l�gYE�ߎ����Y֜lsq�Z"⒂�섛b-�����8�mo����e�ee�7(�R�Ȕ�Y�w�6�+0�,��mض�;f���$���fq^����ٖg[^��ֳ�!��۴��������$������('-�-&ؒm��t����V'f$��'2�u� ���,}vxxy��""(R@�`8с7	��m�0�@�|	"2ف�1UJ��7`w�2ֱ݋����
�\��U�v����.=���AA�S,�\��Ι��F�>��e���X��-�2�lc`��E!P�3q��8�a�-8���ar%Q�J8�E"@"l����.qr3C8RJ������D�a�8Zg��P��� 0@Ҽ�>q�����~jE��3lȸ�ۺ.5������vD�ۏ6�!���(��x�E��j3�$~�S�++X�]	3\�Lq��o����o��=��f�n�XS�3�3�N�b~ �y)v�����?�����x;!�nϾW-�B�<�WddNa�2qSuljq��x!��w_	�B*���k
@�`��9�a�
g�w}�5lL�z	����]^�d�E.��ܱ�t�꽉��X��Pخ����M�/�#C�6vQ�p٣��ԤWT#^��b�޶g���YRָ�E&m�Y�t+���y�mv�7��>e�r�o�[��D�^<��MsD�GN�+Ϸ�[�9����v��಄@@;��m\3�ʳY�����pҧ����u9�P~�0���C�]���������ٚ����JF&���M������_�r�\����V�&74�</aO�����bU�uw>Z��t6�e�fQ��*���͖������Gr]n����Mt�ZPۮ�,,��7�:����}=8z����^��*y�hb���ڼ�Xx�ډ)�<�T�h[�B[Wn�M���Nps�W���&_�E(,v��w�OR5�)s*�cgNk��o}�������1Y��V-�q���K�z����n�����z��>,��,4�C�f�����.�qM��
�w��&����I��K�81/U��|�;i$!���~=g@�q���ON�Ƃs9��q�\]�5�Q�����7@�t>y1њU��yЩ�4�^;�#{�7�ls,����Z��c�Rs�L�V�v����V��S�������f[,�sr��s��FgI)4����9����[5M4�iwZMV;�|���DMOP��@��wEK�iu�<�h��Ǔ^�o^���a�7��WG�)��\ɨsf�*�"|��jBJ�*V��qk��{��vO�4�a� �������GWt����fF8��m=�qi�� ����s*%��gA\{�n|��uא��՛��a����M���o��޾JP���M�%eec��A��⬚�q��cŀ�w���C�^dF�N��YRlʼ�����#����up ^�VP=w��d>�Fv݈l6H
��5�k���z��O)�$�z#k�W��<�8��j�u�uV���#I��^�!�gz���G��'���T��;r6U�0E�Iy�{yI2"����Q��	"{��2�O�@8G�M�V��y�-빋�©���=��񻞣��6�l.�d�!6�n�mvgI����,Z�F8��;6aH7�mla5��;��ǜ��'��D^�S���mn�t�[f Po��f����_4d.鄌���\�z�F]��n�\����ग़\�o��S?��i�a�i����ߗ�%V�Ԏ�w�E�{߲sC�X��I���Wn��yE����m	�Ǆ*i�vfS��vt����ܒ�r�ON�E���ރ^��x�<{�O���.�f�v=^;Ć�|+�.�	��aś�3#K'p�4k�5�[6P�f���&�:H���Ϋz#�z�[��/�����E��{ow�L����c����|�l��Џ��7�]�Uh�)s�$�2�{��q�Q�[$r>4�wf���3�wD��� ������
�\3mY��H�b���O���W�˽��(C�N�Q�ň��]�ED�gM�榌��p����$dQ���.F������?�H��Wq5�븏g�,��������U[
�/9��:w=SLD<�Ý�S^"M6y�2R�uL�p�U��bf������t骓w�<
m��yQ$�"0}��\����f�H��6Y�,�H>��x��Wb�V�
��e�@
6�t�rI�w
2��#�u��n�%ԍ����)��ne�g	,x*<�r[4.����S��B۹޷��a��F�gK��ڭR�ΝX){)���Y�7K.�La*.������KDc�|8�Qכ���<ϐ�q#���!@���/�&{���.��{{&Am��x���ոv��21��p�v��lӬ�{d���I�}k��o�w	9��@��d���k�̶p�ަCT��كE��Ok$0͓���q�7S�m�+��;��8��[_f�G�ϟ��rS����e4���
�E���Ŧ�I	�	�tʦ�ʮ���x8��2�0���Ӵ'���2$0ve�s�Q�����:�C�Y�͉]a�]<6�"ۦv�IJ�ޗ�VY��I����&�a)z��:T����g������f�����iL�=��9�{SxLU'�ѻ�#ڎ"Vj��R{L �� <n����G�z��K�wt)�*�����0t3c��MK*�ۜtS��}t`��a������&�d��}�h	�O�1U���Nz��+�㪪I��������TS-���:;7F=���d���:�s}�����`����h��>Qs��87H����-/����Z�4�l�q�sݼf���`:C:#��u��>�W�*�������ާ՗r�跎�#2��(�R�	�Rj�Sդ�[2j�b��,�Xo}�r�RGj��Oup�#]t��-��P��Z�|׼eu��wV-�����}]�W���������s�V���(��r�5v��~&��{��r�#'�"6<k֕f�nT�\ah�Mv��Ϳt��$�ɟkdK�M2�::ߺ�=G��Wd���g�:���;�{Ir�Y�}�ڛF��X�������
Mz���O���}�{�@7Cf�KH�(|'pk�g:�s�}z��U�fΒ�4l�S�3�dݓ����4<�H�.�\�����dᗰSA8%�+�:�Vq직��{�!��������N"Ym�=�������E�@�t:t����5�*s��gv�+=��w]�7A���rkEK���	�?q�B�휧Gnٱ�B��yvX�έ�.��˒�����R��3�l�d�j�d �����Z�����mc�饚��Z�zX
/���Q�`����wW��)O�:p�mi�܅"k�VJ�;��.ÛS�<#�U O��O����f7#	�W�w9"M�;m<���,.�	�_������ob[m��5��A~�Y�W|g�ie�{��!���J�=��n3xs��3�a�uԞ���g���\�&,���ue��^0����PeF��0q����vOD��ƨ���x�A�������&z|Sn%~8$Ϋu���8�i�v���}+r�+خy;�2��t�3'��䐕��`�ח3e�z�{uo�{����%b-'���*K�Oq���U���&�S��4h��IR�y�N�a�um�� ����iW]_Q�m/��E1띖��`{�v�)��;��M:�H��J}�lWN�͑�خU��O�[̊���Lq;^�>>q�������ӈdkD3��� ���G]ۋ�^kR�z��G�oo��j�g��*3�4�H�v���/���&����ϣ�}���Jk�m�;,�g2Oh�:L�&̾�{�4���EP�����Ι�GJ6D
��2�y��gZġ95�n榝Hl��EۥhY�	N�I=��,�����a*	����۹�����@�����Xn�Ms[2;S0w�Ť���+=$�.����e$�6g��e�Q��Z�n�_,��R6*Ϟ�_Eyi�/y�2�^c*�ۛ���Q�o�$>�[��GK���l|�8��c��ml=�{��B�Fn;9�V�:�,�h�D{��0֠0[�c��	���{���%���ȧ�
iu�廗F�jW�|����0�L��:�G3+b��=\Y��сuѸ2��aw��)^fĸ�Oc��=��a�w�����l3=U"�rDR2�ߎ0iQ�1�s~�}��8�'��I'�iD���;=�pu����;�h���ց�n�^��m�S��ҭ�:��[�/e>�6��1pO��IM�����?��u�|���on�~�wq�Jd����Wl���
�`��ޛ�jC*�E¾�kN����nN�,'��З{�{(K|� X��}ߦ��M���e�>�	�sd@7��=��,c4�� �:$��J�>ud���u���mp��<���� ��8��1�w�h)�j,�FK>��Y���ͱ��)�r�:faE��y�U�Wt^wRha���\gޝ�z�`��������᪹T3T���]e�=�NU��?�R@ϒ���cO�o�]w��e����[��)4+�nB)^�NA���X�󢂻�1���q�H�\K���T_S��:kf�i�}�Gp)(䑄��ʮ��%ηS>�n����Ӯ4��D/l�-�3�]��}��]ʃI.����q.�0jQ��j--nY�F�f�s�킼���
۸}Qx�sa-����[��V�9r�M�&V�������Ơ�;��:�@��=|����r��t�v*�"|�����!��wv�����y�L����k�����'\@n�z������f4�f-%�moaX�]�t|�t[��܂�<�3������c�l�dVvE(�5"���JV_x���Ɋ�y�R��;����3���r|2�T,���a<[��yj�T9b�{o�\:�ڒ[��{����KZnj ���N���շ�Շ�7l_�;<�� k~�^CNDq�窌U�68�=*��H
͓q���ӝ�=Đ���\i��lx�#ک��X�m�aw����X�j��ߡq��Lyu��4��Ud�5z=�P�qޘ�2�zy�}�Z��8��خ����jL8��I*�l��fj/vVC�7�-�-�����`߬<�W���f�}�j����p6����ҿ�[�+_N��f��+vii%e�����a���47N���wP���v{����mō��(�^��׹��۷�. �n��]v�b����)��]-�4	����d��(�y:zW!������
uH07�
�q������l�}J�{n�j����|(��tU��}����\�F�[m�j����.���5K=�u0S�Ax@$|
��ho*v����`�T{5�}q�
~��Q�%ϯE����͵ԆPV����9͓z��q�����k����͏&�t�ɚ��STt�z�#��H�"]v�?`2�8g��DdH��m�$��6]�>�u���x#K���cJ7�Dt>�ʙ�ը�r��fa�g:��bzǠ�veǲ4+�Jk��_Aj:Y�:�Ƥ��z���幒f�= S8C�{�\��δv��� �^}>�`��ȹǩ��*꽃[PO{R%U�����s2E�0���H>��Pz2�/'qu��ru���}��~g�� �6��T�2�|Ǧ;��B�Q�©��Ku<N���ݞ,B�tt�׃r��3�[ot�&��FL�y����L���ۑ{g �7�`WF϶�U���+���HZ������3�P���'��f�|���oP��7��Ǩv�ӻ{ӝ��v��ӻ�L�/p��~��6�����9�jzL(�l��!Q������-���[i�ц�;Y���T�Si��c5FE�k�b�p;��0��P�;��Y'w���+Z�|�&r��.�ֱ�z��Q;�˨b� �+m��E&l<��a�87}]�:UZ��I6��:*�}x�;煊dm�U�'r�4T+����t��H_Ue':���!l9��p_j������0�˔��=�E+�`Sg]+���[�//B"�ﲆ@����=f�����^?�5C�fA.�⩊�\5�suu\9Z�����X͚Z���n�˩)���'L6����v��!/��}�ɀ��c�b�K�,�͓�<��\w��q
{�q9o�1��.�9����R˙b��i3'^��5���V�zy�s�M���/�R�չ53��h�V�c�gP���ri��U��v�:�G%h���W����Ɓ���šOܘ���iS����u��U�3Ht��(�Q]7�2�RA�ف]�G��͕g��;q2X�-��ˉ���ƝtѾZ,��ۡ|�����Z�^�Zf{95� ����tI���ay���zWD�A9a������7޹�O���ӓ4�%�m�(�öf�9��1Ǉ��4�\����U;�];M��ĳh�m��c�1-3N�h�aJ�%n֛��n�U�뗶)9��H"�R*��^�Z)���`*
��,{��%�m��Y��:5�m�`U�>m�ZWv	]����&��?75��׼I����҃fnԹ��s�g���z�i��x�f_k�G5���L�]�[�fDa�8P��gR�J1X��4����Z�0�t�nh��ΦP�CoL�k��jr��1�y�N�7'Nn��U���GKk� �W�c��F�*�ö��}�Zs�q�I���sq���W�v���:�W�e���i��9U7]��%�ކ�\���c�F+�r�vÂ�j��sS��{
���}���r�et�����/3|��]9F�� `�\�0챙�Y�A�e�ta�����f����s��FQ�F+��"�^	]D����`QU�i��E7 �r�HgV.��;�������2�I�l�D�4=������-IG���:*��|��]n��w�j�KN�U�+8��6�tu�k��gz9e�|�BK ��s�x�1��Vu�\��#�5�)�}]�nܽ� ��,�i���%��HAx��89��v�\���1�i��/�'�V�"��C:�Y�-�����7(��=�Ã+��&�Vܝ�7WKNOmo_�]ׄ�������mn\��4]��o�u#������'�t�ba�:
���3 �Y�a��A�k�D���[/��t_k��Rn�դ��O��(�|?v���"��O0"���ӏ��/o������]u�_��N��zzz}�>���v�v�ۿ{j����ݓ����9n�H��P�/�}��wO�]u���q�]u�_��N��zzz}�>���vffY��1U�5(D�/~���g������q6��;�	(����ﶢ���;n�r-��z������붓���"^�{̄u���8(,Ӷ������8$D�:9�m���Y":D����qeؓ��H��k�w�ڷ���Gm�׷��4���Z��������l�������m�P��Y��Ӟh�׆-��K����ID A'�e���h�vSY��d��vw��u�srH5�1OHڛ�]uݗӸФkVa���2�t�&��F���?�7����b|�7Ƹ�܈fp��V_�ܮ�ު
��g᥆s�O<�����nEke��۬*�NPF2I�#�y)�n�0ga�#E�x�e�}�/�[�$fV$P�4�]�= �Y)g��6U�N��U�#j9�l֚��O<mw����O��R%��9�I�%��^\��g}��xD��E�Zo1�7C�~���SRj��`�jG��y���l�E�N�Z_LnN�p%���oG�Ώ=ܧcs7ܳ���|bB��n�z^�o3;�>}'�y�����GQ�, � �;a���_��{*tKքٙ}.f���V��k���<��G+�~��mn�U���,�v�7e4rws7\��)�J�w�p�*|�(�*H�?wKeV�7@�g�l`M�̤��W�����S{�"6�I3��̣����RP��ٖ�~7�z(����]��#�b���v�Їy��At���SF� "��#޽$��h�&�,���,�<�>!�Q�x�r��G����U���8/�XD��U�S�%vE��ӕ��j
�[�X���Y�;&<�z�Ge�uD}�ƾ??��TZ�V�/X��4G����'��*���Oa��|���X�L$[N^Rnk�5?�N�,���2�ƹ�ڟl�&�8�n�fb�'�_)��\F����y�>��t�̵���#c��й�Ɖι���L��"��oZ�0����`B�ĥݠ����7�>�N;L����*鬏z�8��h�����⸶����tz��V���/��Khn�0��żZV�F��t�FzF���Ŕ	S��L���}V~��_|���G�䊙(��	c{p6�}ϛj��TS,d�g��я��XR�q��fn�&M�P���������d r�ρ=��>N�M��ث;s�֒M2�a]:�7#!�t3�(���E\��ϩ��i���w3�땰���w���ht�b��W��X1C��{)��}]�Ͼ��B�'(�9���-��@���S:`�[7 �/jg\e;�8�3����i��z�<��j�󲥇G3�T��L��R�������n�f��l֍�l�����x��z����K���#g�+�6��jpC�W[��~�����������__[pg����B�jƤ}�''ݎ�쉽��8n�?���c1���#k"0a��4v|��IWwr�ћ}7MѲ�ՎLQL]�C��b�ӑ�m���^�x�"����#�q.��
�=ח{ե�^	yGun������@z�؁IGq�S��0-�Z�٭��;*�Nj6Oc�{S@R9�H�f��`�����$�T�3��2����ݟ�9��30���-/>� �zH���L��h󗞙�]���\3hx�-�c�ӹ���@2���!,Rُ�^��\C�`��M5��m+��&n����zr��x��ʹ+��-��v9=Ct��z=�-�{�G�%"yv������2P��&�j�<q������^�3�[]vm^`���P�̪2��s�γ�>SD��~���$�z��z�u�T��m��f/�31׍�}�My{����("6�Gk�a�}꤉��*܍��uճ��X���/(�ʴ�E�_�R�ۇ����X�p�<�;nNob���ت��f�Hl͙ u�u�w�6�$�@��;�����/AyL��(e�W[�A]�ѹk��o!�1.c�;bҦ&�"�y���&8�6I�G{=�q������,�]N���s;��
Y�3���BdR��>��/��L�Yh��Q}�N��-�1�+��I�A�w��σ�u��Ճ��.6��߲�]Nۊ�A�d�$dm1�C8�c0�~Ȫ��"�M*�%��y��en��/o=����r�����������Ĉvu�4��Y��ĳ��;���W TХݴ/H]����L[k�o[��T��üH edwV�sh�)ꧪ,����u?��ۧ�H������e���G[����R-�w��n=>�3��+�����R/W�*�i&�"��3�Mşs�]���æ�=�Nur��hSoMauY��:�]��o�����E��m�c��5��9P�s$��nq�~ՙ-�uȄ;3�12�����R9�="3N�'�����O䥫�{Mv�w�2螮�g1���舧��E�8��I.��(��o�p�7
�x6�~G@=kje^�j�?^;�V�Y4�vl^ ӱf����Z߳��wN�E�`5�P��]�\Ûu'b���e��M?e]ɗ�����h��N%	�8;�����z=U��GQ�ٸ�7>��:A���<�qC9vrm�d�a���e�=񐱝M������q�7�
tn�l��UG�W]���d-OՖkLΞ����3/�[��#��m(4yC�7.��7�px�vO��i�W�����	,����G���-���ly���..w���.U�C!���xӴ�飮4�����b��G�l�L`o�h,�4Ì�qԢ���Q��on�|�ś]}�����R1�N�:���O�HL�G({Wphv\`s�[T�^��c�)��LzU�e'X$ϴn��ɦxB���)�Z�M�Z�J��gh`ǻ���|&}��;�.�Gh���{c�\��en�D��;�F�}x ��_L����H��ԏJ�36���Z�0�g��-�TC��F���f?_��	���g{�v{�lϴ�5�5��L ����g>5"@ŝUO��.�ד�u;Ә�Uc�ŗ�i��h[�Ƽ-y�%/�M5FY��_)1�.����̼�^Z����B��H�m*���U�����b��n�f�,��^8����d2�l�imz��*26�y}q.�l������w�Y��D��2�s�
�Uf8��3�r����>��fy(�g:�d�:g0jc�o;'w3z0Y�=��׆Cj	�H�?wKeV�i�&������망&%-89z���QB=�Uz���6Guvʐ�W�sg�b*F��7\ݔ��c���
�9�Б�6������/!���=B��( #���Hm��׺w��� ;�^ncO�5����1��0�瀭l@�Lx�NDy6l�k1�1�8�<�yL wŘ9���c����K��TGUmqׇ�Y�͛����W���+�!_��l�4�K��.���D_V�M�E曏D�[z�\{�{���A�����`�yhH�����c�8N�t�H��96��&75����I(hCj��6��Z;o:0�6�z�ԏ�}��Z��̔�N�!L�Ļ)M*��<4�;%^��ը]b�kboY�E����nRg+pŅr{t�e��ww}G�ƞZ��ڹ�U��Ŧ�$���p��S���̰��A=Z4oNi�P{���qqqs+��vK7��#//�|�;����
�z3`�*�B��%���9VCB��@[W����װ@��c�|��\��K�v������e��e�w^Hkf ��(x�U�b���b[L >ܼ�M�x��U�yw���h���N���A�Q�9�盅���9L��u
3�uy���7']xR]!.q|(�h����S�p,�Û�U��t�=ݳA�cU���vc���w)�t�]�ʽ������,��)K]�]�Oe�������z%^���W�G�:k���@B9��s&�\���cp�y��3��;�̆�0Du�m�P�;���uwN��<����S
���x4U��E�7;7��[�y�M�9Ef����ܫ�a.�?GwZo���M�3��Y�����qW�A���TulyG�+n��ϐSY�'5��V�=G62�" �ڜ�"�פ�J��h]���t�v���;�-]qB�Pu�ϴ'��P���M}r�Z��ؒ]WEݶ�q?YȄ���N�:0�G���m]��%��F�vTk��4W[�v���Q��#�ҵuX��bU���s�vU����V!�4��1�I�2U���j<�[��dt4?|}~q�����f�:i^����\�W�N������{g��"�G�%��� b�����Vv�Gp�˟F���͵�&�t��\;z3���P���4�c�8�n�aa�T^w����}�erz�cͪ{�u��TW�__��e�:`�L8z�YF��bv�
�
��8$
�q�J ��ƭ���m������l&^
y̭�I<2�C+�0ўbK��^����v�1��Qde�����:gN]_p�[v��iI�� 𷦒=v|�Bw3[��ɮ�p�����LD|��	R.ot.�W�!�� �,v�8#�=�"�A���%��n��k%F��u��0��]WO��5���uL��ރ^��-�܏�3�#����D�Q�/H]��;����p	��f�T�D����c��c�u&�۞�����Vt)�{�S'q���פܭ)�g��DgJ�=`;˭]o*#�F[���c{��aH�m�,���r4�2,Bi�6�������>*s�[��	���]Jӳq��;��jd���{]�M��t��c��G"�a������yq���fEw���<�?��5�y5�h4Ş�[}P*%�s���a�!@w=\���S�캅=�g�Ε��e�J� ���I�xL�'�ow]��(������.͞TkI�A�.����Gws�IU>_N�O�dN3�Gwf;5�}؉���Q�����3�gu�Zǻ���OrR�[>j�R3;-�64��d����dY�G]ٝ�6N��t)�/ro�}��e���9��FNML���q.���oJӂ�.�,tW�dB4�lm�8�+�Wq�&"�⚫2Xʜ�@������r�}���<��hD.�F�	z�%������Vp躵���ٛ��W�ϖ��a�.^U�[ӝ;1�W��'�Nw	���hb�,�I*��#[ �y��Ad,����L���'�'u��I"窀� ,q�'3����F���=u3�+��$��:[����gT��fq]��8r96
=���!��ȳ�<iM	R�׹Ye꜓O���3St곑�pw�R��Z?I�Cn���E�װ�����({7�躔�h�w�=ޭ}uj_+B[BԺy�H������6�s{�|����������:��\"s����xS�TL�2$$���:��u�k-���J'm�"_լ�39���J�c��l�s�BJM��iTC��mhk�~;�K)��!�/R/��@\�3�\u���V���_jW�lJ똵���p��I�ӧoB����x�M�z��q�{�t=ܪ�0&[!E���p�٩�;��������@ϩR�7~z���կCH�g�T;X�/9R�~ۆ0��Տ9[�6w9.�S�#�ʏm�\۩��pb�=�A�e��<χ��M_M��݃�Y��G�΍��~)#�B;�����F�u��-�s:gt��-�,r������������*RK����9]��Gr��*u#¨x���\�^��g@8��:.����]�SQ��/#^3N颽�L���@K�|(^�|�"�)7����C���~Jiө�>��]-p��3\��1k�E�96<��';æ��q�4*�+.�S��6�[.�|}/�p�t�Λ�\�mط&�^�#�&�p��c�*�B����*�
�tK���yj+�u��Fk7D��NԔUk�gS5�S8L�p���_;;�XŶ���|ح�~���nk�G�LӰ�Fnf�(u�X��^��+�/��^�} ؐWL�,(	bbb���
KpU�⭚S�*�	m���|�%YʆIt)ss�+.�y����M
��WR1�����7�Vm�)P�G�����c��#��]���Pm8G&��s]���n�u��-L�{�Q�̸�e�	RӮ����;V��ɇs:�|��{	x�L:+� ܩd��PBV%�CB� ۭ\��΅�<�f�w�2�ܽp4��!`��ie.�4�{�V:�z�;-������5tQF�k3��1}.������&BY���]!7{Ԙ�%J�O���fU<�u�ݵѩ��et�0[}�.�YQÌp{b�B�7�S��g3L{�Y��oz�l�B��mk��Օ4Q�O`ɬf����L{i��&�b��ջ�aHd�M��t�D��{k!����u��sq��۹��p��wE�D�J�Ѭ����w�(\U-uN��5�E3v���C����R
#*Vwtv���+7&^':���.Ty۔��RTen;�y���Б ��H�^�����}��I�������9-œ�y�&$A��H�"}�/�f/b }H�����bIS:�N�嶥�Ⱦ�۔��n!����3D3Ps���^J����z�Hw�Ń1ށY��[�gRэ��ܻ�m��zܳ��b���\x�/6�QV��/��� ���w�b�/3xガ���
�v��5�(m��uj`���:�;vm9KL�}s+6_f7{N"̨̀.N��V��wq�i��G�CI�s'n����!J�t�ۤʲ$��#�	�e��]v�����%32��s;�γWSm��`����/��J���;o;��Z����%�Ξ��Z�/Rf�d�������%n���Z����9��,����9%)uD�\�{N�|Ҡ)�=zn���/�ܒ�^�����
�A������#�1�Wz���y{ֆvX�W�	�ջ���<#F���w�j��)��jN����Ty&Zj���k^)�����e$��c�C�B��2ub�x�m)vx`t����]���Vv�L��ӓ!n���un�\�����k�o�*��]�4IC:�ϰMU�Ї�^¥>�T�/*՞�*e���+5�[��J ���x�MTa��\꜒#�\�l��3xy�СS:]����D�ڻ��4�u�GT���}D�|K*d��֯~>��k�v�lGr�L�>��ǧ����=�Î�뮺���]x뮺���������;��9�X����m���;m��՘���x��}>�Oo�ێ�뮺���]x뮺������������23,+m��m�f�?^��sy��S��m3W�g��n�o-��K,��pm��o/2ܨ�ݭk[k�W���x$(̛E���-�{V�H��ݓ��mE��z\D%{[�,��m��^�w��{[�2�#��'Y�"ok��bF�_T��+y�I:N��[������$��N'̒�{[�ӂs�j�N�6p���ݙ���+4�1���e��m�c��o�	���ai��,�i�	
!�(�l�=���sr,�.;�goM6��s�V��U�G��=R;3aI�����n�Aw`7�E��sF��2�$�CY!4e2HƄ0��qq������(�(m�"��nBY�HY��1�܈$M�#f3�6Yp�8��9�!�0dE$N5 *D�Â(H�-0�I1�;�������u�k�LaM<h7���[��s�T9�vz^�YZ��P��]�QX�dSk�ɑ���>�M��ԻS�1�[c�F<ñ�ٙ�v�7+f�P�l���;L��|/OU\�}׊%-�W��!o��љ�� �KJ����=Uʹg74�x�z��Q����{��=Nfo'�7�5�i�Gh;����i��FTy�ޘ}�j�v;5��<J�H�4y��/���~�s~����50�$�A�3����z;�>{u8�=I�o�Kl,qu�
���S-3WXMM"O]	�ʏ3�;?� `J�j��}����BF�_th��y*t�ӷ%b��J%�خ�b�c�{��
0�˟�*�ʖD;*{��ͩ�w���|z�*Bu�M媟C9���^B��?5�ɖͫ�;�����T�SZ�C�+�ܵ�k�[�l�l��hb%��;Y���}�%�a�T;M[�xu�Ít)�F���fk8Ó8�c����v�8v�h��m����mC��kV�TI@44�o�m�2�[VM��T�k�+�/ϥ�3_;5����ɻ���\��Kѷ�T��<�$��aSy�]��ԧO-sخ�oKx�N�fهss����N��^o7���r�袉/�=�©��Ft��l@�H	��=�K]&���c�Շ%�����:�V���齖��WkO���`�ˊ`�ys�q�-ea�W ��^�Ԩww_����� ��������묢�2����杷^�%+QCa`H� �̈��p~ar=v���M=7O�ƌ���'"�t�z�A�|�= o�UǇn��� ��X�M��O�:�q�n��8-׃�]" �����΍���Z��&Gt��8�O;�NO���֚�N���ˏ0��-��p�dli�'��C�Z�Có�\U�Wg'⎹�a�]:
�{P�2����!��~p�H����lj� ���Y�ǲ�T7��̨��¨��m��8g,�ً��O���P;)[T�<�� t��"��5$��n��e�+eY��]������6��η؃����I�V}�-�٨���.�5�x����h���X+n��b�~�%�~>���j{k�^ ,�������=\.W��Sc�g	��$6WU֙%H�VoBpq��w!��%*!	I�2wX.v��yt�/���;|;o:����$���|̮���
ԁ�����n�&�g��.�����I�]�W��3���n�\��b{o��K�K!�3:nvZk�`��͙ͅ��"��6�.j�����
���w��o�{��Uů�w'J����A�M��U���[y����
L��MDó��rRz6����>����������î=b1��rћ�:)��<���}o���m�8W�#*���i暸#έ��pT��=�'n�6_ogN�zG	�#y$|Gwv�rxJ�>_nS�^̐޻f͎�:��5z��.�'�܅�w=+�S����{�*�ef�ӪμȪ=Y3g;��0�����^�����6��q����my�6��9ɵu��K��)�ӗ��M.�\y����(ݾS��W]�
��]1�����C���7m�H��h�,Z4pZ��ɟH>�;a�ܥ$�s$���Rt�F�w��Jʐ¯a��8WX����3:���5��b���4N8��D7J�V���2�v��Ptnm��������ۗb{��p��O�>}x%f�:m�˺X�l��;%���vat�)^��:�f���|�u	6�ķ"����=;��x�>[f���Ps������T��'��}g.�Ʀ�����{���> 6�p���AhCH� �/�����2��{�c���; �JC-\�E�Bd�i�㤉>u���f�b�8�䉅��Y>I�	55�b!�n�Y[�d�޷Ψg��p����R�|���wMVODpaar�d�Y��~��ǩ5t�'��Ʃ��⇇�@<;�
�pP��Sj���U�O�+7�����f�˫�Kr�5Q�替o{X�=�g�<;��t��5k�Í�]�ړ4�ᓧ�9���� ��N�myK�:��zb�^��͸�����j��xsV�.WM���U㫺����r��Ҕ����o�৻�v+(���]�>^qO����{�������E^u"�<��1��#�K��_NkF}�u��G`-^�HuIR��+�B��]��eŨ��{ׁ���=vU4�ԉʾ��y�A�r��<��\5%M�ە7[�Pf`�M�����:�A�3�p���_����۹߿_��I�&NN!�s��ZI�KK$��u��M��_���ϼ��m��j
Q�T����m����\�g4LD��'q���B�P��T�g��2���ܐ�!e�^>#�����ލ��H{�25��P�d�У�z<m<n��ɻ�i��wr���s�
A���6d76ߧ�n8p#��;f�u-�0�w�ۊcl��z���]z�mB�[���H���29L���y�;!��8���wJ���7vr�ά��*X������J:�� ����|eS>�p�M�&��Y��_e����V���q|�Ѿ�k�Mx�ƻ����379]�m�Z�"^⛳w�߬Wz�@q��.�*#�u�*v�F�G�����dgu�ݚ���Pm�j���9��6ӎ���|��s:n�z�C�t��\�5�X��:����Y����J4w?�C�O}��{|"�n�XH1P̡j�Tm~��r	��w�'I�8D�J���d�El��Ǚ<|h�x^����V�بr�<s�+ۂ�&3���@P�g�B�Z�����42���,e��K�s{w&i��ȸ:��e�v��'K�h�{f�0�y�Udb����ԣ���R@)4���S��g��S7�9��<�LՍ7�0�nQ��=�nfT�37�r�'ڋ@t���rZ�]С+#��=9�9���� �w����}U���Z�JU�]�[6�.�n�5B]�f����G=����=���̛J|*�o!�^G�W:�����Í�w��h���y����C&������1ǳ��[)(�d�y�1ު��m�ƞ4qi���B�t��_�k�[X���S����$�q�Ev�;��OuzڦXf�v�m4�4]J�wuS������C��r:�\ƀ6�4]��v����l�G)��c���#Ƽ�b�6c��G�ۤ^2v�s�NUi�g�2=hI�ѓ��y�*��q�n؛��Ro0`���=�m�Wo�)x�f{7�m����P�"j�^s(+靾�6����x��E��3���z��hm0_��ʳ�Ì��Ujk�0�GlSs�έ�l	y��mY�#-vZr�q�8�C��ۀ����l��h�5#�H#B	� �AF��[��^L��Lgn���ͩd�Uu5���F�O`Snt�X���l}��6h��,��y����Kp�Vľ[l<7��~���;��c�jg:��ޛ��$��3��m#�V��Μ'��f�dy��3H��r�܁jz|`�K��k�L<4�>�N����w�GU)� �f�m�f��Ƽ��x�;XK�H����
�q>F�f�+û@��G�e��JA���>������#2�%;<!��yy�g��a�;�l�F���A�D�� pA�bq�;��`�Α,ܐe�i���C�)��=x^���JW!��>.9}��q��Dڸ��ZI��|��D!\�i`�����/@!!up��-%�b����M�I2���Sy�g��P��UIp-�q����ɻ0��D�9w��*#�f�՛���o�o��f�n*%��h�q"yܯO\$fOV]��ί'���t۠�f�)N�N�s$�<M3��w\G|�Cܜ�O��o:����"��^U�cWIZ�SO��~6�T7����ۖBU�jv��¥�[G-���n1�'ylUT͡���s���`o���p�utґα�chT՗�hU��q�3z����!��/�S�w��<�oY�d��E��!
��6q�l���qt�@>_N����)D̬���p_��lZFٽ�\�d�����H��]&;���x���a꩙�A�K�n@~�0��~���p{<�*�{���L�Ȟ���k�[�0�b&L��;���M�8�q�R�6F�*�q `>�t3��SX�Oy��'1��µ
:�n6Ck�ò{@5�D 
�ي~���j/VTn�h��ٞ'������,�#��8f�5�.U7.uk���o\V1�V������m$Mu�F��]����4���q�[Mb�)^��$\/8��͗5�g��sU�@"ޝ�x07R64��_L��n�����ô��G������W^&T�=��+g�h��7��u�骯Oȼ�����-@x�UR��e�4�cީ�ѕe�IdbA�����l����2At�|W����g;��.ʡ����U;wh��D�XO-�A�.�������ǁ>�ْ*}o�X̓w�;��N&p�b��l�K�ڐ�N�B���^��V�c�i��딦t�W��z�k���_8�������yfр�gl�Npa�2z2���a3Ac�2�>7�B��+���������4��𿟟�s�虃w�ʺ�-\���-Җ��9{���V�FP���O�o���kw�Lp�=ܧ��<��2���݅U�r�������%I'i�ǲ�Lө,�)0�Wq��٢����X ��ov�s������W������<8x�H�~k�ɹ���v�0jn����+B�l�6��#�*���J�uf�)�/�w*s�F�e< 2�D�8�`��Y D��l�vQ1����wE����[P$^-�l��飛��9�kwW�p�|���7˗����-��ڥ�k6"ݘ��7���<c�&̲m���C��۾�Rng��{ۂ�+/�|%S��xm�=��o�D���|�ߤh��~��;��uy�������C��7�,���4+ΉKf}����^B@B��f����K���ejP�2c�K��;Z`�3#�e]v]+���%n�`6��"k9���2�3m!�Q��Õɓ���i�DL�T&�f"��o������]K����`�kc2n\*ď�ÛY2Ss�l~�y����F�:�>s�z�F�Q��|m�q��k���z���|�*�̩y��D�������q�#遼�@܊�u1X�_;(T�D�hSL�K��^�[��ټ��]���;����}5!�}�"\
Mq�Z�ʔ�d!�C^
��=r�8-l��; �>4�+��Z���WS7��S6�ng&�5KH�[����$��^��#*A�}�����m�����'\��y��&�(�]��?Vb�~���\g�n���6��c4��0Z������AG,GB�*�b�C�%]�ܵ�6����D���ܫ�:I4�{%��:�Z�(�*��:��\+�Ҩ�wWO2&6�j��y�7��8`!�&\�ӯz������ۉsud�Ú}BȄcݜ�^��4 T�8{-x�U�И�J�w���d�P�z�q̟�髯<�C�}	{#�=Z��~~b�L�3F�f6�ռ�����&�P�c&U�Nod�͢��2�I,k� ܱzFH�O=�x��{P4�^�̉��<P��Qx,�i}�����B�J_*sr�T�Z4;9v�����sV�G��}meH��	�Z�(��ifi��.��S���q+��d֮vR�k�u������:ݼ����ׯz�Ń�6���2�F�뷖���\C�NW>[fXy���Oz��KjX�bL����9Hk��@�����y2�g�b�r�ʸ�T;�o���@�}#�۩/��Ǒ���F�B�4�8��-0�YF�X�D��u�&�L��3�����ث �7���>�囁YYj�8�A�m��Z�냗9��,�B��x�Y1�
���ޱ��iq�i���z���1m��0j�TYy���5u�S�6.��]3d���M9ʘ�F<5Z	]��9|�YoU�惸�C��Pn�O1*��V�YÜ�ڵ8�2�.���^�s%�˨W�3����F��Fi���A�+a�kgS�ऌ��;�g:�7��Y�o��%m	}8v'SdR�qKoS�'r��n�wd/�f݃�s���f ����r�jh��ќS�Ir��<��Ӡ��&K���yG�+34k��L�:M�+;@�K�ֹ�!VtNX́�(RH��M6�:�-�߁�s���x�:0ˊ�?�oNS��� �H)���dG�� ��՞�g۸~f�Oh��J�޾M�o���;L�֝b�B&�S�Rޛ�(.�AW9행��{j��7k�s�:YNd7Oo�]�p��Im���M*wb��5��'s92���p]��m���3�:򶮟7m>ṥ'��F�y٧�m��[�^8��;u>�쇹��92�XSh����Pp�}x���cݸ�N�bӺ>�����}�`�/P�N��ךt�w��Л{����dc�	U�Pu�dG7�e%Ȏ��ҫXo�j�.W�oL�w��݁��HN8Q��b�]�i��m�5V�o�E�ԯyJ4���6�� Wy�)�����ݖ�.SF��w^ˈ]b�P��f���|��R=����SSf��nNCf�>���:qGٜ���hKt΅Y�ܜ�"�Gm���)��t�PlR]��Sp���F�)BV�*���6�%�!U�L�#�̕ף,2^��bd�l�e�ά*��O�����K���kLYX����R�u��c���$����L�P��uio�ΓgLػvf��K>XE�3�ޫ�o��OWE�`с���Ŗ)��s=Y�m�	2L�;��A�������pL��閾Y�Wy��]�gm��{���{nN�mߧϾ����J_{^�5�iI{w�e��浔��x����}:�}>��]u�]|��u�]zzzzzu����;-u�y�w铗�ٛ���d��{v���~.v�w���O�����g]u�]u׷]q�]uק����_>H��	����ʩ�8��$u��6���ex[~v�Zۧhi�2��[�y^^�ŷ#��d�Vu�G^ێ��%����#���Zui��QG6�l�m��ޱБ�Q׶C3�����,�^��{��mgZnu�U�k�г����N+H�����mc�yy�3]�%5`�n��l��z޾ؕ�ݑ�Y�ڙ�n���k�ٸ�ku�޷'�۲]���Y6Js��I�c5�6����:M�E����ycd�6v���awξ�߷��_�Z�Z��UvnI0a��٪�WN�(ξǒ�Y�.p�a�?��w��>3���5�P�{45����_�ί�؟v�����̖��V���ݞ�����~���\��6�D��B��\��!brawk*�l�	)Z�6c�CE�;�6�co5�oXw�����#U��B��x��ޔ�� ��ؾ-�OYĞ-���q�k��N3_��z�M#z�Bك�ѵ��8]�}d�GJ�����X)y�ʝ�dlޞ�������0�@��#:D)���U�{�׼��w\Ȫ�Jq,ݭ�(et*��V�g��V�4��wL�+�czE�w/\�I�n�v?v�"j���{F��0u�I�9�M�OmZ��x�M).�Q�l��_g��2��FғA�{a�CD_c�4�J��������3����0a�㮉 ���焙�b��7���+L�I��:#�*���rץ>��W�Ӌ�N}^%L��F�ٓ���r��dO�E��ĝ�"P�j�Х2�g5=��d�Ů�Y�G]mi��{|V,N�����>���*��3[�Y��Vԇ	V����(e�/q��h�}�t�����N�ݦ`��̖��7m'm�i��ӌ/�o7�'�g�t��կO�B�w�U��?��ڽ#<�]GU'��0�9G�4��G	�wBբ=Y[>޷�B¯G��t�L�hȺ!ۺ��U�κ�iS꺀�K�@w>��.�S�K�����nD��bg�����	P�l�M�m����N��x����"��tzuO�e6�&��%��i�%=44�Y��Mvov�`T�De�KgrV�;�w.d��|�ܧ��j$F]rL����'���SfDm�ݟOr�k�� �o�rL�7V޳J�Rv3A'3�ּ][�n��\^<��v_=�'���B��Ұ�I9�ԷO.�ǌ0J
�p����}s��M�8g������eξ�2�׸�'H�S�Ͻ�=斍ƨ�ò{K��Vk�T�i�J�
�sb��5U"�Wa=5ջ*��N[C7۫�8h�#�5���lS�J��,N�ZiuT���U�ۤ.�J_c���;�F�� ���L�96pngv���9�$$�D�a��R�mÔY�:�pT�����/S�,��z�����3v�1����!y 짻M��޻��V�<�(~���ϱv_���px��ɑ����N�:n�81�[��m�U�0.J��� 8x���l�����H���Q�#Z�߭̍>`l>����O�o���7x�8ǜm@�*w;�y<x�P�H�ԗ&�X�2R鍢��`�hRP�t@{���H�tk��~�Z)����k�̿l^�Wf��$܈�/�̍�����?R�o�T1�ٙ,�l<Ol�}8�Q���yy�ey.� � v
��.f�8�XOy�=wLMIj��ƅ�LRٻF��ʜ��Y�AT���Y]{�a�P&�9�*2��s��V�̀��Skz�^�3����;����r���Χe���^�궣\�ѫ�7aϺv�b���
�����G�m!m�Mc{_rv'T�]v#EjӦڃ;D;y���·\��J:Ѝ���$_�[˵�Q�P�Q|�dޛ99���e��4�rɎ袆�]����c��9.ɺW��'x1���F�|6��;�F)�7��]�Ǿ1^u�:���e�ӱT*�{ǥ�Dh�� �v<�7�m�ZՖ0k�Ӂ[vv�����G�{ukh{�CW����o�4.���Kh�=ru�SW��:�Xuqs�������n�7��7��HZT��f�Y�91���l�]?O�L��cB�Ǣ�=u�g�34U�v�
2WX��]lg�v��6e�d58������V�r��_+p�-�LD~����p����k���)y�(oX:�$�;t:���_b�����o�AG�fim�!q�sV��%�w��0`��}���m3꛼y�[q�[��t�󾋤_@q>:��X��|' '��;3I��-gl�l��wTs0oj.{xh�8)S��i�[��8�U�y�ׁ�wNV�ֱ��Xp����,p���{P��j`u��~v�oV��i����{3UN�a���M~,N�:(ϼh3�v~�P�֕��c�7<E�g�7���Zڻ�\�|��ڔ���,tJ��u>CX ��8>�/{
�:�=�,���g������q�-�ԧ���Hí5/�e�\��"g$vw�~Ny���zV{�!��w����@�:�\^[T�K�0u�f�
��v�Qᚡ�9A����+�yǓ����I'H^#q���*��;��<����|��DmIX�)s����m�/Euxިv �d��?��M�'�W,G��N_Ϗ����&���0�d}�4j�&9֊���t����wW���%{[[ݻ�KV���j-�w'J�c,�6;$`]w22}i^`�u��ѯ��6�ض֪�-(�Ŧv����K���:�9��c���#*,_H|�y��+*�,�Y���^�����C�OTr�n��y����c8����S	n��N�����W}��H�\'g7��v���]R] .��^sm���u���a"[`u�ko駚��T��*,�~&Wu��A���z�^K��w�x�P흭���$���i���3�:�2���7��J���7�=|Z0�8.n��L��H��wFr�nyP͍� w͙\�'2����w�-�F%F<8ո�e��z:��#��6^w��H~)�9��v�M>�kF���7i̛�ó�WG�VH�g�!�������p�6�����E�7�82	y|8M0[�tn3T��
k��
�wn�E�o�r��e^���Vf{-����=�:��mI+w�7AN�}D+�3l'����!t+c�m�=WXGI}is���d��fjn0n��g7_Y�}���6J�Q͋��7���jFd�ol����}���8qɱ��N�e^j��NI����}�E2��El���ϥ5��B���w=�	��~�*�*/ݧ�ly�]���$�%��Zy���õl��h�4i�	�X���q}4W,^�ϷR���0b�E�bGKV��o��Ge�-�F��)5W-����䵹���^ԴD5=T��D��=�����zߤg��X�:�]Ez'ׅG`r���]u��m�;���{���D�����e�����B7O�L�:��*�4̲���WR{,kU�f�U�ɫ��Q�@r� SO�f��j�u��w�T�<Z�_w�;��C�,���[(��s:�%v�}ч���WuQ�o1u|��y���&�����-I��:(��^RLO {�����w��e�=^V���G��O��W�]u$�6tI(�ާ�-OqGൖ�>ن��u���T%� �%��l�@��� �I%�n��ϯwq�w��G�2�έ:5�.��J�״��nn�k�.�U�}���[�n:��f.��l	��^o7�]՗=Ƶ�����6k����ٸd萙hW1Yy��7e�A�FaƷ�j���O�z@�~Yr�5/}������{�>�����{�����wg&�FL��8i����8ϣ�R��YO8�E��ƴ�t�:�{����O���c���5x�a��H�����Ϲt���:z�֬�o��D�eg��J=^�'��wU醜��4!�����o+ζ�,�ӄ�VC�3�z�j��8/eH *B;�I]c�ǖ�١4��:Z���{l����c��(v0;A��J�nwNg{�vde�}ݟ��W������ۢxs`F�2�@]++��L��ќ�������SN{�I�gӗw�D���Z�}=�P�Z���B*�V�y�<�o�w�YM���ZFqO��I�	>//>T�G28V5w^��y���Q�ŕ�o/;���^Eo#҆��V�I�x�g	��鋿?����_L�6���3�4�Ӿ�+�I��U�t&v`-ә�.n[�� �ךN}v�W�M�X3xяhy�Ё�wg�>�c�6z�`���J9]lg*b[f�<��]�	t�k��ս�����he�_QF)z���!��������ݓϤ��K_�����2�+�W��R�����R=sN�zX𭨗�z:MeY�'1�����ҭ����GQ����S�#��g[��`]�鳺S;���OKg�U�u�7.�u�����A/%�6�*'��U�1�̆�[�Mr�:�j�m1�4�Ǩ�3�E��� ��9���ہrL��dw�}AB4�RIqx�M4�#\*��r�!:g����.vیIZL�k��r�]lg���l�&�^qò��UV[���޺��}l.���͘����kbA5��;��=ǜ�)����˨�����+t��������Ȃv}�ʨ�D��Q!-�W��=vݾ�ˤ�ۺU�;��k?����̍yDoh����~$���T�����rocM%mNO����������c��������]�~�O`��%, ��=�}Ⱥ`�^�:���k}�㤱]i�:9U��Γ�n3�Mw=�]�U�5����{��@Wp6��l�D�cW`0�ۻu� ��p>�s����t궞e��ήю5�#y�S�]��|>OV���잵9�2�Ϗ�zN��I�ۅ�h9�9@s�0:�'I�3�W���W�V�79�,o	�E4����>U���̲��xv;��.w�}�>�Lz�o�2�h���^^�d6D�Pɷ���A�'N�X6����E\�ߪ���w�:�5k5*�sp�F��cog͜$�X0l��Yƍ����K"}rj���ǘU����Yov����a[׻�3IpK�p̳>�m�i���({��KE^���vD
�7�,�#�3m 
V�;y@�};��9�sN��8uO�A��{:�&���m�+b��jp���$.�����GG)[U^��~�^;���J��hk9Ud�\��wf�<Ļ�Lwz�6��n�TJ�����.n�~�\vDs=;=bW�\w���2�'8��x&WpǊ��*R<R���D^U4��>�fX����U6r��Xt�.N_v�վ��,�Zռ(*�ݍ[��5ڈ՞؂�+��r�R`fm�[MRf�ʔ�Z�g.P�V���֫�02U�ĺ�}D��hޗ�I��T�����n�N�N1X������흂�6v����B;>�3=o׷�zzR�<;Ok���`1��E���:؉�<���ZƝ�Gl�l�����mS�7�k��t��{S�14bs�ʎfwu�v�����v�o��k��ޓ�*i#̃�}K�.sp�ڙ��$�+>%T�)�ݦ|�!�,)�{g<&���3�Ng�c��2.7��^��-2T�����}�a��3ׂa�ޘ���v�"�?_c���Q��]�_eQ[A�B6�F��[�Pu6ge��7i߳��N�wp��|	���7������z�Ru������c�ʘ�$O�6A?[����o���7u��R��Įh�Yi�wI�n��z��)�S���J�KNhV���٣�tXO�J�򨫚� ����4�����S�9x�) R�7�tM��N���HJ<�S���?���~bG�" *��DD{���I��A�(����.��yΐP���D�!XeX`VVV@��P!�a	 �U�U� !�a�a�`VV�a�aV �@!�a�dXeXB !�a�aVV �� !�BU�!�a�aVV �!�BU� !�a�a�eX`VV@�$XaX`V � !�eXaX`�aX`X`V@��U� !�aV@�!�a�a�a�dX`V�a�eXeXeXd �U�U�E����^p�P!�a�a�eXeXaV �!VV �U�U�!�a�a�`°�2+�� C ʰʰ���C(� ʰʰʰ�2�0�!"�(�2�2+� C*� ��+�C °ʰȰ�2�0J0ʰ�2�0,2�2�2���@0+� C °�0+H� @Ȫ1T d@HhdUQBAP�� dEBP��bUy��*�@2"�!�CC"(C	
!*�CC(f#�0��2C
�C(!��(�CC*C C CC
 @Ȉ�09� 40	0J� @ʰ2� @ʼ�U��`eU��`aX ��`dU����<e�eXV  eXVU��`� ʰʰ���2�0�0,2��1��x�<�o�UAE�ReDd���=��>����������<G�������p�������2s�]?��/��Gӿ�}/Ђ *���?����(���$W��X�p��} v~��e�)����T?j ���i��#��Hs�<���?��@�"z��?�? �l+�2��#)("" 4 R*�
(P
�(I"(D��$��,��)" @B $�  B2�H\$@	A� !BP �H@U! U� !V �I$ � !B �ID�  @P� $e�P$�iV A@��`�_���T�b(�� �% �P
"_�}��_���~����P���? ����_���Ý���$}�u�������S� U�g���������'�T U�A Jy�����aР����hB�����~���.���'����� ϟ	�|�$�r}�t�8� *�'�?A�ϴ����� �
�}�����θ����{�0?G������?`@���8~��s�$WOQ�����A ~�:���hy
L^������?f�}�ݠ��i��I��� U�jf{{>�������K��o��"(�p������AE�����>��!����PVI��E���)��` �������f���ʪ�z�B��%��[aAR�j��I!B�%KlDI(�jk*U)ER�D)�	A*��RTUP����mP�VV�[-���6�-���}j�)j�lRl֚�Z�mUV6�)m�V����Bٚՙ�T���&Z�ԅkm����F���&,�Vʬ^�],�j[Ul
c�d�mV��E�66��l�m����"�+%f�Z���j�F�m��0�2�KQ�e�2��Z��%mU���k*ٷn)R:�#ln�  ��V�C�]>�x{wWV�V�er�sNۻ��k��u�ܫ]ڷp�w��'��M�޵�:�oy�[���w]�9�q�e���q��{[�.�u�{�ݫݫ�WR���5���VKcMVYj�`U��  m��"DHR���!�C��2'�*�H�����U""�
(��y��U{�kev�.�WZ�U4���붛m:��{���n�Q�3.i��U��]�۝C��ʶ���Mn<�5���l�6�Z�Mf���   �x|��5oKvk�׭C�t��2���ݷE�yޠz���l�+)����h&+]��k�n�a�w�^�ݺܬ�]�U{�v�u�v��s���hFU��t�kF�zTڱ�P�@ƛe�Z��  ��z���V�z.� �k]��ծڂ��ov�#j�͞�����^����7��P����3����U=O;���tۮ���bޭ�ޮ�l[Vh+Zȋm��խ�   =�{uvs��xX�V���<�V�ӏF�Vk�;��m��p�ܓշwY����m��	R��t�˃�q���=u��s���<l�ԭ�FE��"�m�M>   �}]B���{ݶ�il�{z��s^���5�u5UUTs^�V�b��;��Z���ewtU����j�j�W�z�<���8�֥�Sf��VʦCB��   �@��\  ���� �=� (��.zP �L A�V�AoG  ��<��  v&��YdIl*
�+3_   ]x  �  �훟@ �� =���  p� �)�Ҁ � �m;
( �\�@�3fm���+-
dU�_   <  �Ӏ ��Ph�qW � ���hQ�;8p  5�n �چ  ������p� 8��ZړTƙ�U6��|   �ﮟ@ 6p
 ]�P 3�  �8�tn��  z�ڵ  :���J��n��{���t �"�����J�� E=�	)*� h�A�{&����CMꌘLO��SQ����@5JE@� �)PLUP hh3S�?g�~���?_��������K�#߼����4F���3n=V��)+�P#�=�����{�ן?/���1�m��  m�������l�q�co�61�m�  ���?�_���?���ٸ�����մ6�0�M�6���%+U5�էA��)��o�e���r��7�����F*.����q� a=N�li�Q�f�Mb��I�i�iZћJ2j���lL��Rgřj�X���W�.M�i���^����6��Ν��*��I��0��I�v�ڧ[�]���,6QSjlm-��\�o[��Q�Lm���a��X���v�h�Ѣ�˹�fi���+���f^!"G�� @(�d���S�0�2+N��[��t(1n�j�W!o6�`D�&}#6�"J8�((�li�B��"@�p�<�����K�bGc	�q�j�?�k%chV��^PN���<�w�<&f��1�M�"ElHdr�lY[w�9O��ۚ��KNR�xQہ������OE!��̺�OUe����EV�7n�ɭlj�`��8d]Ĳ)OqSƈ�=D���V�{�0��$#IZꕢ�oe�Z�k@RJ��4ĭ�$<����j+{J��4ഠq,ݛpZ��B(l��f�fLKd+tŢ�Y{�I2�Q�)`�@0% �*&'n"v��CmLj�GFeI�c5��«��XY���!�a�6���A���/�d����wB�JGq��< t�h��vn�-C-h� �`��4㑰e���yHZYJ�u%�d���]��L��-�rل黢����d׀m<�O&���2���
ܛ��8�l��#ڡ�I�����{CRS)��Jҷ����i�#�A*��8.(v�fa�D>�%�	����n�8��qf�L^S�!r9V2�*�pT��c2�ܚC�!����#$�낅�M����]N�����>B�c�#�uڗx-���ŷ�R���n�V��3Mn�+J<����|ʥ4�!�i�JTd����0�E���a�b���iq�a����"����:*U��yw�����Rn�Z6�V��I��X͌(}wi�ug��B%F+�FU���V�o�Vkߣ{���K+]*�C%>��%f����#��#�%��)k��7P6��ٴ;d���J/]@�ʷ,`x蕳5�Z��\%j��oXȷq)����!L�*K%��v�zK�t_��N�w ���6��#��"�LotV᳥���#����w����`Z���)��V�ٷmP�.ъ�v���.f9��dl\�e�H ��r��N+wr�2��֣����nӴ�v�Te�Wr:-Z�IA�AWz���p*RӇ0SX��,e:_
M�Yf�"�D�n��8,�E�����'�t�"��c�'�A.3��z�w[L�d��̷�-�d���@Um+K3m���#��B��{��g.�W�L����vm٠ރyvnn(R��Xۭ=�f����e��/R!Vd�*ܹ�Ķ���M�9��5v�#�=p�{ZTEV]d	��ee��~jя&�N�x$ڶ�Ō�f �*勏c H�I�ʐ9���eH2�`�Me%��"���Csc��X0�ue�-+�'a�7�&�{o6Vf�&�Z��+�q�-N���m��t�5�J_Bݐ�6�7W�^�]J(L���bݼ���Y�j�m\X[����Ϙض%��#L͹�2��:n;�Z�	���Z�O/^=���1����aZ��*��N�*5����,�I1�ZV���S(�C
8�Hmee�/ʛ�'P6��+n -�1e\��⧊�c,5MdٷC]�L�,(�N�-��weZ׭��.kkdt0j��L8Tѕ5�g�N�T�T���/X6,�u�)�Z��W,^���iɨ�t�u2�En��ƴY����9��9[5ԕ�$�j��h��.��%�1�9M �̕B ӷvSc# :�\�vi����ڊ+YfR�X�i,@�V��Z�����C���aD2��!�@�5b��n�í�@�(I���D'>ݐFՅ��֬�2rK�#�<��u����@��N�Vm�Ԋ�X�:�ƨ�U��:C(3D�Ċ��58 H�������C�e4(^1���l��%eτ�[�m[�V��,�m
�n3�Zر��<�Q�n��\$�n�=T�CJ�.�]�����r�F��VUe� 7nV4�aa��nj�tv��E]�v� ��w-��]�2�փ�W�N�����Z5֢u����QqeF$K�G0vt���v����˴f9S2b�m�42/������e-)��i<w��,+؞Xx�OvO���u��+M2B	�X��a	��ν�{ ͧ�\Ut�1[M[.e�*�é��
X�vK*�af���+x,�]BЍ�V�`ֹ���ѱy�b�gر�m(����:b|��d�si���:���x]���@cl��2�&m��r]E�7#��,��WoI/][�2������%6sL�n)���i5�����)�DCJ��=�BQ`k0�r�R���,-�sA��T��)V���V�ZѐQb�|bz1MD����
e����&��ۥub�Y[V��3nʇEa����nh #�k��Uq�bN��Iv6,�{��Z����
���4աO���# 8��X��oԚ��֜£�Q��a�V�y�m�`�6��`�3 �a
�a%��w�-@һ������;�5�Yv�Xf�i\��K-r�0#kQ'e̩hӻ�k�0,�
T��f�P\ɢ<��TBG{�+C�3RN�3�1U(�^|�Ě;�z��E���Ŕ �t�5Z�ܣ'c*�� $�fU��� .f$%�pYnC���#��R8!w��&d4֊�1+��Sb��56�]�v!u��[G�Z�"��Q��GΖ�t�Y4-�}Ec��^�.�Yu%x��g)Q/[�@��(��ЗP.e\j�S�խ���N��C�2e��j���Y1h*��kd���p���`�d�K��R�rŬ��Z�q��7q���ҷ��mr�82��-��x��N�B�bw���Bn�U
֕)�c��W�DkvZh������$H���j/ u�
HRTj�aw��cY��8�E�1��]ǧ ��!jP�1�1��ӛ�H�I��{[�2�ȼL�X�a�)|���r���6v��e'Z���l�%Pr����"�*���q��\j�V��hu:=ԝ,q�e3�@Z�u����6�ҕd��ґF,�X��a�/��e�Ri��6�=�w1ar�u�BS�39J�Y��P�]�z���Ev���Ģ�na�m6�'ѓ���A��ی�	ѭZ�,9�v�����]Ń��==`��S��iZ�ҭŪJ�����sJ.�E�w^#-d2X�.�=2ZLV5i��ҧ�Qƈ����E����Հ�P��L�{X��l��,��.�94i+e倞& ���}�����@)ZR�[��؞}c4"n�F����ծK����m�.�%���/�)gDܼ�m�l�jt0�2[�Lm���*	��K&����A5��.2�3*i�X�I��Y�wI"��bK��-���qkt�p2��S8��q�6��V�ܢ"��Ļ��Q�U�m�4ub���b���;{'��M��!���/�ә�n�(��t-|��jә ��&�$��[���҆��	�=�H�p!z��M꛳�ْ�[5G�p5A}�S�ޫeZA�&Jj�%���P��F��?���j�
m��q;����v�*�T>$,�Q`�7�sjM�d��f'���I�HBV�}���ɡ
����<6=圧�N�iЂ:��MV���ʹ��+2��l]�+AT�f����BsR�qF.��u`����	�[��f�E:�[9��8.���A��=OV��
\*� YWyWyFI�F�?�E�PY�T�n��P�%�J;rGY�ä�!W�n��.9�f���vU֬�N�);Z��X[5M�z���⛔i��Z�2W�9��v;k�'$����ӻ#6ݽ��{�l�bT�Z��פf�Ҭ�N�/i�b�nb�)�>:$��a�:�w������U( 2�c�oa!����b$��)X��S�����B��{K5��jy.U�%�.�U�SYbV7�Ei�>˔��	�
��H˵����nhKs��2˗������v�B/�J�\k��5M��趥d���.b�m2jskl�F�FD�q*Ò����IV��:�޴��04Ѳ��ˉH�Ȯ�q3�aշP���>�H�m��e��n �<U��Qf�����X�n� f㼡���ц�L��(��dP���gt	�������{DQ��p���&+z��snr�aۗ� ��z[D�.nAz�N���ؖ�����^�>�e�fF�0��06rJ��6Jb ��Ѵ���a��p��1m��OÖSlkP����#�]]�V2`��qLA�jV��7���Qs�/�u02虊<���Y�G�i�$㩚�槨5r���ʹ�F�Y,�`:a+�͢�.���'�+v�J�r�O2ƫ�i���A-���"Q!R�7hee��0��U��Y��^]��ͷtqGH�@��܌3{M+r�H��"�P�)m�%9X駋��d�n4��,����]���n�0���i�"��*d��Z��p(��򬖣զΡm�2ƿ���%�+Hm�w�鷬-���Y,�S�DZd�NԎ��M�Y@�7��åV�F���~XѦWע�{r]�ю���'�*�9-�;l����V;ۦD��//-�<�h���J*��)���g�I]m��ݺ�â/��yV�X��,�9[������l"D4�-[z�m���n���jY,ƌ��{���iJ�Gr�ݻ�Su5ǨG��ʥcr]���ASL�J2��9����̉�IU�t��:�CX���M��U�SU���S�FfKE�´hjCet�b��6"2|���ИK4��h���Ƀiy�Y��NI�/C7#��Vm�I��כX�j鶝k����-ԚFǒV^V�%� �u��
�SM,�O^������SNQy�"�l�^�q��:�*a�)�jy�h�N&9��ÙN�^�ҵ0�vt��Eə���0��ƒ,Y���'jdߛ�e��%�I6�[s6�%{rS���l�k�����r�S.�5�k�&6��w�R ����
�dB��I+�t�2/*�b��QG���`A	�Re#6�L�l��<B�݉I�%�/"������dt��A�4-�^j�$o"�ӂ�l5w*�ikH�f���kMV��]IS�SXI���Z�i��%�Gn��h�4��1�$V�b��%m
©]��{v�d���BDӨUJ�Akh�fe4l�8�i�,챍9f�Kvk ;�v�1�QJ�v�\ְl��Ol�ՙ1GM��8q\�����M�U;dV���m��^�7,ɻ�fK��1�B�۫��m��RY������9z�YY��6E4a/#�f���	p�*e-h���V�Ы{�Ĩ�r�K9�
����X�����m�5f�u���Ր(��d�e+
f���f�km8�:�Z�#�fn��i�)l˶�"�V��)w�p�ӓPv�{Df�ky�C�i�+4��r�饷V-k0��X�
��T�۷+ࡓ+2ޠ���۳'()��j(�Z8��z%��6)��i�ӓnl�tk-bm}���vmդ2��QdܤJD�#U�T\6�l�������hū啩��%��(�9�j��1:̭�q���v��J�[E��i���6�ݣb��V�ib�F&4�Ԗ�1���`��N���]��4-��6���+B���1�:���[.ʨ6¢�G�itn�8ްtT�Q$�ehݫ5��,;��j��KHt�$�J�[�kt�nl�m��8�V͢qI�e-�a2(4+�P��&�In
t@�6��̒����n�zd�ov-����Zwi^TU`h�s�N�ږh�����LwXS���pYR���'��.�ى؀���%�wZ�֘5]��y�Mjo*h�,@�ᒘ׬,��@�7 ���*�c&��-�ȕ)�RȬ�Y7
4Y*�[��5���Q�[,݋�E�dP�1� �k��r���
;u�Yf��>���ǣv��.h�� ��W�*d� j������V��7>��K;M1����3 �R��A���^�ċ��u��bjѣ��SNM8ܻ�X�Qزn^����.k/n�6|�W������y�����t����L��Г���?U/]^��f;��4Җ�E�&fUųb�S�EX�䂈�@�;��j�3o�VisDiPMj�4MZ�3kl���A�XÅ��y��U��3bc2h�f�iH�ˉ�76֚��;U�Ì���9S&�6�8���^�H6i�k5���@QՍ�y��
�1�:l�
�d/0����X�1Xi"+u&�CU�{$I�M�K��Y01��*7�.�oklś��^eb��mL�Q����,2�"��Yɱ�����v�<W��'�%6<�TRefՍ��� ~n�"��X�0�&�V&�YP��w�_kPݩP�x����;�)I�V^n������^[�H� FjL��(���V��60^b�2�����ż�n܎�'d�<ښY3we��SVt�qi4{:מ"�.j����RAv���T���ѕ�p��넡n��yO5���4*���u��^F�1i��d���x4��͹Rk�:1�����iϮ�f��f�� /K��z�T����t��*3D+mS�[M�T.M���{O�F�F���y���G���[R	�s-'z�;R!Rn;Z���Rp�����`��c�E~��a8ܻ�%FwĂ�7
�V=Hfj}�t�y5;N�Ӽr��$\�Vr�qt��U�c�o+�.��Q9��wW14�q�WJHڱ�o� )���Y	���_b�D�M���Y;�ꘅ�V���1'Ww�l��%-��c��ml���s0����XU�=�0%h�jw��,y�����N�a�ݷ�v���7�}��q��3-�jN���z��׍�?��/�~�Q�\����sy���4�K��*%݉�}mtt+f�}��գ��{9xs�û�C��kۙ��cupr �.�h7����$শ�e�ot���a���]�HZ�}3�{��[q�f���Ҟ��@Y����E)>ۣ%�o�vN��v�����Z],�F_!���Ί�ؕ
Л�G^�q�a�_]��G��E��rg��E�\
�r;.��M��}ڸ���zfB-�q�Fƅ.Vr�N�ON��{Ip¸d#�:���awnNa*���J�ԪI�-p��k(�P�va��?�R��Ϟ����t�Z���
��E�"]�H��¯6�s�<����)�f�[rVV�[��\wLs�����3(�=ȃZ̰���q��A7m��f��[���t8��7A㈉*�]��96��Q+����=4��;%r�J|�f��N�Up]�o�g%h�8�Ђ���<�/t7���ȏ6�N�ԭ�M��F�#���vʍ�M�f�ŋ�R䕹�\�<[��R:�y�Y��Y7A�3.������V�R&!N����7).ץ���\r)[{v��5�|e�E�fb�nx{�F�qR'��z��-ز��]-�[�n{`�z�kÜ�W!��/����(�[[�׉�o��Z�	���Z���L�)u�S�T9@=�؎��Rb'y�T��`�K&�JR���9��_���Nƻ��m��Ÿ�U�i�9���Q��Џw��E��ML����R��Ӯ$�l�T{�t���l�w�^C2ʳ�#��tB��@w��=u�MOC�X�����ڦH^�%��[9W�O��ĺ�̮̆��I������<��=�=-���R�bx7��y.�������+E�(+}gh��W�x,�7'-���y�-
l��W��,�V���ܽ��&^FO{�H��}D�/ݼ!`����(�-wQ��S��}���?^���Nvrх��ݭ�*��H�Ƒ�P3��}{`$�y>Mb�Zh����G1τv��.����>t�l�c��b�<�59��L����	��"���;HO&��{����or��3i��_nt;B�EV]丫�o�Jn��U��*��9MF���� jG��)V�]l�EmG���v��=�bN���pru�U�il5�a:};:v�0ѭA���4nR�-�EUk�����Ab���[\V�Rޗ���{r}os��C���Qբ�^O����-���1i��qq�/b��x�m.�����]v�G�<�r��HN�����:��tY%`�XN�v=.�/�IhӰ-ڗi��,����kv�m�e-�HUԽ��z���S�N�{��؏��U�O.�[K�D� ov]�J�"�h�¸V��o#�ר�>y]�-1�#����Jt��jo�Ʀ5�e���9,�G�V��������v���}76N\��%6�T__p
ckN1���P�3;4��ٮ���%��R�a��u��Ȍ�j�F��oh�0[��x��'e���M�o0�����n�g�U�&�5�c^��(�u")b8~7ڀ85h�Hl[W�v8倬��uǅ���!~���p�R/h��Td��hK�6���%�K�̱�˥Sw7�R��ٍ(��WO�݉��բ[\��u*$��5YX �4�"�i�=�w���1,�G�ٻ�J�Ӎ�	�^�ӌ��Ԛr�����,Zk���o޺]|t����fj��-��$��ϱ��{D��^Jw	 ]V2��*�T��m����xO(Z��Ӄ^�.�2���c�c�j���rrr1ZU ͓�֩��\�����yzcY��ʬ�R�X���ê���[VI����b�v�˽�m}�g���k!��7�7�Ө��#����:����\a�Q����Z��8yΠ�r�;r�%ts��tKjj�Fv�S���Z�Y��Yj[��{r�G~�+���jc��>��EY�;��s�@�������	�ޣ:|+���KH���h#yb��z/�w�
N/LT���N�52;�H�[�[����D�.�{+cQ�t^�#����1gi+>^�VUYr[#��ˈ��A�?��)�G��J�}���;�c��v��ހ�x,<P(.b)�g�ra���oۖ�Ucȶ�jɝ�����ۖ/Zz�Χ�>56��R#�X۷�V��ڇ �[��l.Qμ�#78oK�_,]��gq�p��K�T \L̰H61rp��ֲ���fƍ	/kx���:��s����97��E�v���gB�{1�`���`����ȭ}�+}�͵r�Os*�]<�cy(tGt�`�uX�t���^ӒB=�7��Fw<"q/PNG�X/)z&��Ҧ�����:�j�M^T���}�P�r�\���o��U~�ޠ�D�/c�i�D7���ޖH;�P��}�e�Gᾧ���s�S6�4�����Mu'��V{;�H�Vu�l("`�k4��7�py:j��K���)��u�X\����c�m����ٺ���%��a���g��O��W){2�˾�F7�ҵ�=jqϝ釘���B���Ϯ�+�:���5�P�j�}�څ1()�&���0\���Śí'v=�rn��ɫ���[��W]�	]��ԃ �:�^�sӶ�^�����
嘸�W��&������p�Y��R��
� ttL+փV��3N�W��N7�F�Y;�p�4���Nί���dýNk��+ݬ����\mZ�c�����k�0����A]�\�8ro֊�g1��RR��us|�4Ш�A����0�-���9&�f3�MՈ��aO~	�"�']�7�p:���J*ry��枡�+Z�9"__h��{�\����+�ѣ�Q��Cy����v� ,�{�#={��v�ĝ�Ȫt��?,A�Hgj�o���w�h����V^�=�<�P�|2��v�'k��8��S�|0^�a�{���t�k]Չ�]�F��ڵ��4.��ғ�-2c���l�!��j�d�����7\�l����Z�H�4���o]A����I�T��M0����K��g�b���aj]s�x�-���z�19
}ztҰ^���гy�:m�;]�I�V�����SyF<�j�\���7V+��v��
Y+j=��;�G �����;���ל����vÖ$�W$�c��w�2�ynV,�g5��@ȭ�<d�J�񻜚��^P��l��bTݡ'mk����k!�_W�c�6���(�+*��f|��i��,c+�9|t�n4u��uwH��
�Z�2c81�t5D�"˽�=�v1J;:람�ok����]��IҨ�+��VUi��*sbݾf�@ �L�v'5���%�ޣ�["��\��d��19��yf��q��nD{M����9���ᜅ�vڰ��x�U�"���v	2K}�f:\gJ���0���,A��달��K=h0��`��*|�8yEg4�&�N�9fcX���/����/��h��
��ڰ9�q�z�,dĜ:u�,���_��� �h���M;�K� �w����E�FrΓjٱ��r���m��Q��;�`Keqw(i7;:��O^>c�J��+g÷����Ǚ:��W_4B���q�y��C�sJ�M[�wYU;^n'ۂ�YKl0�l�m�نd`3�S�7k-�ͷ�|����NtN�Ae�@���&S`:���d�3���l�z4{H����c�}�"���e���-R9
�q�@=;D�t�|9X9h��\�F�^�������͆���yqzY�n���5�I>Rz�}��4����W��q3XI�<��J�'��ąe���w,��쑍���;ە�,� �_	��6����<�3D����L�L3�`#� �'z��G+_��K�^��y���B���uش>g�!���٪���tƽ!��WM�F���ZLїZm��#��L�[�+z� ��mL���G�{����X�l�꾲m�6N,��+���ʫ���T�]ys���l����q�m�6�@�%��b܈�\ڼ��4`s�����[=�"���3���Ӫ�XU؝=Or�E.�n��wj��"G��i���jh���-ˑ�umƆ�yռX��jKE��*pz�S�_�͏Ka�3�-���uƪ=�����C�k��2��R��d^Fx2a�80���L;�I\�EA��zJ}�72��Zή���q+F��:���)��c��d��\s�.3�:�Ֆ:⽂����z,x�i�H�x�m[�.̴�;z�b�]����a!a����6&h�b��X�q^�0VZ:�@Ӏ���5�\��5���ͣ��Ee�"j��Q&ijR�V(p���ܽP=�;_/hU��	ݪ��K�q��O~��Z������]����d:�v�&�A�w�=�[��`�^�ݩf�Z�%;订v���L]o]��;��	)Y��"�WSՆ��Pʚ7�m05=}׼�/����͏x�ڟ;s�Cb	%�+X�7�V��ۢ��<���tR7��P}o�K1�l�ҕa0z5lJ=F}��<�OT��:=��\j��	���l͓:��MӞ�(=� Yd̹��r��P�U�p#:�ើ���q�sՎ;3P�l{�lgU��*�nJ�V�dW���NĶ�vˡ�dI�Fw�}ӵ Z���<W.��R�e� D9�k����_]��,Mp�\�쓙�1R۷��h/_���;D4kE71��/���ݕ��b�oCu�u.z6�g[Q��sf�,W=쎷�7�y���۟1`�^�VOK�����q��=I�g��u�����=:1�,�R�❼��h��oo���0¯7��2zv>��վ������3Y�-�C����y���k�Sע."� ��N��\w��GyZ�/��j�uf�;XZ�
���Q,�gT����M������`�
�d�b�.���d�+��JQ-�-:�F��P$+=��-�B1h��z����U�H�l�.`�MN�t󻬹R�Q���K�y����o�5iL�F;F^e{I����bhWLeV��]�O�Rsq���l8�x����p5o�7Rn@��cBѽAݑ��P����	���L�)֌�p��s�s�n��0��0��9�S�_mukIf�y��ZN�AP��=�&H�7��r�%��i˵u�L{��F���)e6��g��kS�t��ג���.L��6�Xf�a��c�ʻ�I肵��sV���*��t���a�}���ĳ���_=���y��*��t�'-{�.tQ4=�-.vIc�#�Parmq����-���v�"�mH�s&��V�/�m��#�����>��>�}�]�r�ÍX�]u����F�Y64̵���!��8�-40F�l����v(d|Z5k/4�K����}�w.M�ٹ�3����vxd
����9g#٩�.��m���{w�H:�n����gZ��uvL�b.ThhP�NiOjv���l���(UʜA6�.�azNV��5gg���a�즗>5-��i��V^e�d�&k�휷��k��<J���&��t��ud�Z���I�� ��os�S���/g
���c3w~d.[��YW�re�B�M��{�/��,�-�i���n�P�d+�R�*���s�!������&��|���XKD�,9��f�	q�.��zY:ܵ�(5��KF7�mCH\���lr,s�n�x�7�h}�2�k�@v'�1<����Mw�q�hӘ9����瓉�$Jfj]���$�9�J]�z���ps�N>� n�t]X���b���l⻖�=!E�Q0��{�P��m��n���¸��ݧ^�v�dNj�&�ӏk0"�{4XC�T��y�eW;�1��Gqr�Q��[��h7��t�Ic�x�6�2n�AeI��JH�+sd���	�#�C�]��@���{����Oh�k�pd��� �k]��kO��_b���!�s�.�2�����X����8YfN�.�e]�xZ�h۽68����=��/{����S�s3d����� �wd����8q�"Ŭ}h��^�(謎�n�_<�!�$QTWl#�Ob1Õ�����:�$�����R��vf�b������;����_C�4�s�\�P
]�۔&d�U���[�P�7k�c�ft�'N�}K{��(0^�쌺�A��=����"JZL[�B�6=�����7��5�$�	�]�c����N����../I%�W�X4�w�Ł�[���4��h�\�9m2�.j��ft���'���s'�n���X����Jիr���e�s�S
�nB�O�g�Dn�'<t�Rs�Lޏ޹�u�h|�q��]3nf��F?]�<[�9�q[c�n��ޖ��O����|�t��?UiƩ^�Q+5���"��|���5��˲���Y�/.�w�V
B�Uttr�ۤ�DS�_�>3�goy�W7h�r��r���Z�l�љ;�@�嵼���X<c͝C�4JTVv��1%R������۽
w��0.Yݯ��O��}o�hS���[��i�ɉGq�������n�E�����
u��S�콊hY(Ce'����vz�|ڠ��2�K[�mA���ts�u��v���,ۓxN��DZW�N��\���m�1��{���mv�0   �����������'iJ��'��Nɾ�a�wn���K���I�I�.�IԬ����3S�=q��,י>����r�g=��Vz�"6#$����n�{q��rT�,W<�+�bqA���Y5ܽ���9̙�$<�0�:��y3:\��>wqJ��g_E�&)FJ�e��g%�8��NU�/��\�W�T�񄲰%x�%��z��W�.vpC��qTƣ����)!���[ƞ�L]�Nb�����U��X�=W��;��_q�*�e@��S��q�e5�s�3n�D7y�>�9YiIU�}��rreJ'2Aݯ5�m�O��k^�==�	��jqGI�W-_G�3�d8�C�Yx����%���'�5ҙ64ʼ��u1N��a;����uOk]OG\D��x7��^��
X���U:X���޹H���SW���o��}�X��l{�; ��+�`9ǯ�K��n ��Uʔ�p��>Չ>6zRs1�����UKt�]#�O�^Rսu�Ԥc�B��>�����+=z#�.9-*W�����q�n�ū�Bj�-�o�����;mi|�yˮ�t��HN�ާe��":lHjW"��N��k����@�7�������X��u���1�[��n<�|��}j��Nh�X&d���/�o9���<a�v�,3B[�RJZxQ1j
op�����kT��2K��N�m�m���+�y��]`z1��2�Q=������g��)�4�*����$@ܑ�nu���X�e%��u7�-�}k^�Е�b+^���ѵ�,Y �؋Y5r�j���
R7.w|�^'y3�����ֲ�W��w;���y ��a�J�qU��B��W7�\�����q��Y���q`+ٶ�P��v��z	P��W9�^�i�����O�T��O����T]�S�F.3�8���kRE+O�W�-W���t�z����+�R`3mk�VB��N
-�f���ul�}9s�xK*˷���p{��E���B��om��|��T�"�:]���:R՟qzT��N���b,� Rܽ�F�3@ָǩ` u<%�jj�t�woFฦ�_*����v�})�0O�9Ɖ���p����c&<PQ��K�&��^�����M�Z�A.9�v�L�e���M�D^FE��ћP�$��c�N[���j�ev���:�'nLj�܍4��J��@���K��43|�<�ڎ(kbԉ�&W[�z�t��Ø��L�a�*���E}F���/p
a��>�4�S4O�I��%��P��ȝ��d�B�ܝ���QB�vn�eZAL[�5:1��[��/�Ֆ�^�!e�;Y�O\�-;Pe��NL�Vv^�cDg(&X'n���������-Ǻ��	�w��,�^}x����$ͤ�#�虎XT�n�+Ε {���4���]m̠w�(��Y�X�M�߰{Շ�`�0��wjs�OS퍚غ_ ���1�[��\S=��a�b�	�Z�p�t,^̨�����8�WOa�x�U���\���G�1��£��f����vNu����h�T�d=ҤB�Oc�]����1�׎T�dQ��Cz�����=K���B��r?K��C��i��\4�Wnd����Gs�[��A"ux&Y�*e+D�)���:���0cȾ�dLi�����#z��EW����}�+� ����f�Þ��f�{Ǵx�h!�����N�U�A�8`6sT�����cV��7@p�ܼ1l��,��g>*��tx1�!������c����t`�E��xS�QTϖ݅�Ӳ6�탇9b�v�4^�9���Z���ڗ�����zr��l>߬�6V�&K��ۚ�x���\�|��-�wx�|]i��Vu-9ij��Uumr}[��]�a�w���`]ԔX�$74T�FEM��n�m����T�f�[�|S��IuC;e*�t��$�_9,��}�R�Ӿʱf{T���{Q|,G��'7�D��4�i��J���1�B�	��Ʈ�������C۬t)��L#�t��K�u=ȅ�GcA���0W��2�jt�1P\��_?DgLb��2�H>�b�{}�f.�e���^3������u#WR�Z�7wq]�D���.�\fg�HY�y*n�֢�R�F3�(M�C�ʱ��J�VܻȄ!KF��98��2�:}������t���S�]�z�����A���	`@m��Ëq��Z��tr�/�n�������������h��&�ĳ7��C8���)�Sl�lΫ�􅷻cq��^���p�SZ��O������wUq����Tp�C����I�L�5�m��wz����k��E�ڕvl�5��$kP-:�Ww(} B��ǆ�:n֪�q����
y��5k�7Bt1�/N�XEn˽Ӧ��J��Ǹ�W()�`�ܓx'�*� qm���v��ߞoT�T�O�2.�&�m����mG1��YZ<x�N`6����:2�׆�ےn�v���t���I,f�rٺ�a��B�v#8�;���+);��N���A+�V� �KJ�iH���=�&��ߠ��wd�8h2\ZN+��o�Akp��f�󧎗	0J'"�ɐ��e�ͨ�)v%�v��K�>,�=�f����!Q�G���Vw���A���#�u��H�k�g�-[XWfd|U�hm�K����B��y�N6:��uP[����T!��̓E��:�̚�(d�KZs~�;�#���xƅ�H1V뷱�C�Y����	g�7���ޮ$����篁��`�E+�5)%�
�+��4f�����C7�"g�R��]��m��m5��B�ۢ$�j]���"��vp�)?��������Yz���9�Z�e-��Pm����Y����D�{aY�QW]���$UKƵm"D��}�6�C�D�r�G-��9����:Eu^�\Eo@�՚��,��4ǻV��go{�GY�w[�N��%=�\�[���_{n�_e85ns��r�e2�B1*��o������{n�fg,b!�A�:-d��0�=��<�'i�N����<[O3���e�Z:Lqj�Zp�{k]�.�75Ū�ԑu��-�@I��z�f��"i��Q*L�9�ek���x=;��q������Xp|+L����ui��Ҳ�gx8�^�������4Il8�0 �#�։� �Y��9]{���m�02(nƥía��ݥ�t�]�� F�����c�P�7R�;'�X�d
͡ٸ_W�0�Gn5�w��ţ�/��s��j�82��M.���񸷝�&����>�D}3��w���r�U��}%�w��8{�.�mM�,�P��9|#ɼ��7�cC�'\w\�c�@�E�9Y��ӽ�ˎ�� �%}��}V�/n�yU���'���+rO�FrJgNZ��+���'.�������cյJ��wA���(p��\����Į�K���&��?2"����wBOGFnu�7�K\���7�]�"�"jZ\�����@�������%�s�� ��%5��K�x��y�lVko5Y��!h;���|E���Z��ڻ�1,8;�5Z��E�^��8�x�l2����F.��nbK����(�-P֠���K�ͫ��'uKg�s�=ޏ���=��*"�h*���r�K��Ýi3��M�K�6�V,��X� �k�7!����*6�&�u��cq��J�ӗb,
t��K~w.�<��� ��?%�=*x�A�C��g#���7)8��EҮw1ftFd��;�Ľ�Z�n���}p��w�ExpAԥ�̍0�xo��,�d:d8���[������t[=�u���;ܴ`�*4;��ax�J�ܝn���nc����}�hChҡ�V�v{tܘ,���{%;2�P��/�kSz���7I-���]D��[�� r��<%�r�k���ﭷ:�s:吏�B�� n�;�#��R΢�4�{e�Q�T�5u�#{�)mn��L�o�*�f�nl�ԗ�(��,��*@��@�\m�D�]f_EW|�s��5i���z!����������Cْ�ٲ7��U��s�`p7���8�[�Z��t5��y0V�q�Ka{/b� �(7���+	�r�b�5�e���j�6m]�e��N���mŲ�˭C17G�:�eY����z8�E�uí��#FV���F���{ne��G�F�U�M�<��ZA^���j�P���|�'Vד2|�F��e�g���&LG��]���6��c�O�r���Y��kx�]=]	�:��#\�R�k�Y�m�ݍӫtz��WL�f�m�X�`\#�zs�6�	l\= ($-��x�� �ؙ��}[�{qo^�5X��%hΑ"�t�I�)|�����P]�|)o-��/w���Hg�M�:��Q�U0
��a�x��Oaʁd���pE���EL�;z6�D:'3���G�T�'��Zl��7�e��k]݅.�a�.ct�U�/��8X���伕o= e*�m���QM�H�i�Ln��5��Eœ�wY�Ӂr�{�T)����&
o"ߨz�P��n���n����h4pq3�,-�/���=k�w &�`��b��3Pl��J�R��Y�m�7��l�9�����i]\ݏit
���Xm�љ���mPnŘqހyV /u��b�QnApB/�����k��)���ح�I��滈����>�z�a痓�y.dБ���ҕ�����j\�k)��A�v(P|R&9�|s�ֵ6�����\�W��k�	�k���],__K���<�|����ءn�:���{wye�Z�.2�kķm��D�^ёƾ僙�r`�9�Ja��q��u������x���G�wH����D6s;9>r#�XN�x�JXr�6\z�ض��iD�-��!B�жF=�7��o��q����U�ȹ.�S��,�GG{�Q��vf�[��HX�qș��� u��U��mjC/���7���n �C���i�
�]��ݧ���W�S`���M�FF �㥔���blEZ�Q�g�5�R��3�J�T�Cl�{��������p�6�Gt(���X�}���t�mBp���3@�d>A2�f��gd;N��OK�A�R���۔Nkrk}w0N	"��f�0��<�hZ4oQ��AU{��Ҷ���z�wqf_m0��8醓��R��iKS�hot'��ٚ�)|���j��fS���q���쥣^=�8��Gj�p-��e��.��6�r,N:G�\jflٺ=�]�=N�Kj]��c`�j�)Q���[��g[w���܎lDm	��X5]GH{��T]K�S1�� ��՝���8/z'זT����;�]V\�qe�tV#C	Fє�}U�b�!g�zQv��.�o_�=�k红��k�gz٭s�bڃ����u}
̩w�>S����Mr5ܦ�n���6��ǻH�O��.7S��z3��~��]��i�X5!�}�t�g�	�E��qcifb;�Q�o�+� -�C�HWq�]C$���J�[���kZ| �5D�snM���P���`nkՂ�-X�.#	�3����n�經R���֞�N���TR(��ES2�m;Mp��u���S<���tӷ�U�)ndUx&!�K4+p��ΐ�X��n��È��U۾�����R,�t�.u:b�l=��H*�eꮻg�����oy)Z(?m:K���ρZ;�>AR�6]ը�Sü.1x'����p7����5��WZ�A��琥�l1��ȡ؂���UIf��cLU�{J���ӭ���[P��r������.�S�i-�1,��际p��'��*�)nVn�� ��b%Ʀr'��d�MϪ������y�6�_$�/gA;����/.�IA"�K�.<�SM�>�w��CR7N'-�i��p�bX8o��OK0�����j��2��롮7{&���њ��Yf��c�{�G��u=��@�KU�W�hLT)�5֮�n���-���ܛ�y�/����p.�	�8Qk�c�b����W�Cxp����w=nS�+����݁/���{�2De��5�[ګ;�D@ �j�-hjW;���j��nV�ݦ�"I��\�'9y�q������;��l*�qG9�澥yzG*����!V{��%*D�'j��}�i��A�(X7j�do3s:*Q�1d�dU��Ȏ�J����mY�ҘTmo���Wwe0:�y��"���*�tu��vf��w��X.��T�nh~7���W�.��N�Ԟ���a��V��^��kbU*l��9V� G:`ЬmJ�h��zC#�yr�������)u�����WAnm���s_[P�O�ng`㮥�\����t�3���&Y�ҫ�<��dp�}&���y��[��`�vS�l��-b�zll���o�B�۵�,�g_py�&�O�Ǣ���öo3��vEB�ר�$B�#*���l��6fp�w�솲��v�
��F���	��C�ytn�K�Ŷ}�V)���ץH=gr�E�a��GhՐ(h��~Xn2�[�ٿr秬&��S�Σ�r�Ɗ���f���"�&W[��t�:�T�uZ�z������E�M��yn�i�*XU˒E�]����� ��I+��_S�ZoM��&d���f�{�ݡ��Z������Bn<�IKᾙ�x{�بi1_r	at-�!��j|��.�)����k6��N?���1%��EAL���;v'Iu7��$�{S��-�-N��m*ۮR�� �I��΃�uFE���!}��g��(|�Z�쬻B��e0ů���m"���������yn�(���}kPs��fo���@�y���BQ��J��.��_DK���;�@��WTf԰ڇ����N��;"�+��>��^9��Qy�RSo���R���峕1�A0C�=l��װ�M�m�q�32Q�D��z�Bu�N�:e0�vF�����
�BP��;�.�D�f�7��j��U;<*���R�a��4�l�'��[�Ԛn)sUl.�^����Y�\�/����N7�X�@G��˵�հ��}��Y�/�[����s~�Q]����ι��B�F�W���Η�.��ł�v��P����p��W��CEJ��/M��ws��x��k�5�Ⱦ䊊��w]��s�C��2up�ͦ��˻}/��Q�ꌂM{ԁ�l.mX�����uu9��?t���^	������u�y�9�њƋ�M�C=��O�o;�]��i��㮾&�Ӻ�t �f�_==�J=4�ΞT+/�ؘ����{�M����|���8�RB�泌Ry��<y/RJB�1돓i�}3�i&��s׊�O�!4�K_�f��Ê�|v]�ɈP
Lȃ��2k]�v�[�>��դ[�hڃ��9����s/5E�9�Ӯ�y9=�n��Jl�6M�[O>V�(Xۆ��<͸�n`���r��{F��ܭ趃:�K�����*0��ja��&�K����}/#���U2tFT�
�W�RD�|	���yXU�L���\�Q4�"P��<򊤬�ErªI)PP؜"�P��Ñ$���i�*(�A*�$�]9�Wp����NXX�BL""+E��p(�D�"�.U�����ɔri�hE˘�А�$���"I4�r�\��t�!D�BxNwE�+@��9tV!{�UDE�E!G��l�P��U"dG3�%Ht2.9���!n��̨��	�NQ�EIXd'HLP����yA��D��P��\�)B�����v�R��t:q'7E�3�*��\�w�F#�#j�Νʙ�4R��'2��N��&�0��
��W,�2��H����TL����֭���de�A�/��.L\�
ZɱV���̍�R'%dn�@i$���ۊ�N3l�i������cof�e%Uv�G�h�]T�=��F�D�����n��___R_E\��ؒ�SW���]�^�ͻ�i~} ���ؤ+�=2�zWbg�{qDrz;�-���1�kv�����95���$�T�FO��7OedEPA��U��_k^~)��p�gR4�����ڍo�^E��u��
�d$�\,t�/eV�*��+����-XΡ:M���@��^�6���N�?9r����`W׉Xf�́>�smX�ss��ʸ�#�'�)Z��M7,uo���G����
|����U�XYY66���Q����.Uw�������+�g>
oy�+�=XǩZ]%zL%dt���)��^�����Lޝn&\24�F�����ke��p���S�7�*�F��O�w"����H�p��3��Y��oN���8F�-������[�HÇJ��/V��:LW�i`
���O�C�<3M6x1�J�Ug�r�#}m,��r�IԖX�b�=�B˛e��(�Ȁ�i�j�1
�Ε��ySy�@1�Ç�;��m�灝��p�b���׫9g��iA~�V�������u�}�m�BgtL���I�=5�� oV���ޝ����$�$|��{�O��[��x�g����#��r�Y��<���}DV�[q�f7`�=>3t�y^��f��_��Ї���;H�O�����uBb���
�R���&�ϵ�i{8����B�1����\D
�8G.��������B۠�P��d�&-�w&+����i0��"p�O�Mau^0;7$�y��䳐a�g��b��;��)y�=������r�4Eta�; W�ӣtV�����B��
{�o�dޥyip�hg�}c���[ѧ4(�n��Q�N W�#+�@[rΟ�;��,sh���Q^+k�}ے{� "�8攪ܓ��R.V�D��-j�1xS _#��nuZ>��j_��{N���lv)��]�s$u��K�`ŷ0o���4PuA��],b^t�]Է�ԣ�ͩ}�K�^�,V����}fM��_o��j��ΐ�z\\mBb{2#��z��Ըs*��	�؇*��3�r8�]VoK�D������	���;�9��ZU��l��C|�=S��ZX�N����d�:u�����G�����M��>�ã�IA�7z�*o1������0M�/��j��n�w�!�j,�)��{H�ˌҙʅ���Ǉ�5���ײ�V��N�Rk�vuX�m����SH��B��oJ��!�k�B`���mZ,u��Ύ��t�+{u�@V}��tY��q3�ee�y"�uꜶY����%�A�Z���F��D=C&w��T�u�yX/��c[�d�72{�`u>g�Fe7C����Zd�C\t%��	�{���R�c��f�+4
�k�x^���e3��ޣ���5: �q[$�C)�y��B��璜��ٸ�IΚ���GK4&c�E�D��q�>���v��G>���M��{��L��V��c�1�n:6I�|��bI�=3:5�Wf��f� ���-���L�V�+y�S/H�΃ݛغtJ��\�U�����0��=q��5��JW>��r��8%��Ʒ��ݽ�ڪ�i��!aq퀍�NW���q^�I<@�!wH2��^WA��?Jo	�ۿ���-Ko���"�,��,�n���3���=���B�jJٸ$05�B�������؝�¦�n����֔:|5�>V�!�Դ�Z�&CsmA�s!��#�2$���5�]����۞���>�/�r�6�T�͔]yv��7��k��n�H���l�����ŷ�Y2��m`6�!�+�����a��j�:M�P�T�ɋ��e����Ͼ�����o"�\�p�8S����?rnc*��!Z�3����X+Dc�P��M-�R��9�r(��_GI�0Z��Ϣt��&��^�R��;WWq4~3y����8�1�=V��m+5����u����.5+����', ����UW���/ϧ;�U~X��҃#���vc<+ً�U����_y�6�d�����L���+���=�6�}���&��T^�2GW���,�+�'��Y�^ɦ��ƻ��}ҽӨ`�.t0�e����`���A���6i���V:S�𡿉��r:c��9&o�v6�-�ջA��Z'�&m���Oпj���E
vy`A�U_���6yk6�uūР�@b^A}3���ݓ���:�7;ˬ)h^Pn�P���>۩Y{�����-�S��A�>y�YQ���H��-m�/l�ϻ#Y���w�_��i�#[E]j�����u�{f�ԐH����F��T�
�ePA{�߇���=~t���e���=�5ђ�������u� \�%����tܬLC;��.���/~3���}�n�y����V����b�{<v�su�CR]ȓ��ZLx�>���F��L��'}Y>kJ�����XJ�ؠ�t꺻�"5�[��h�r�	��ڗ�C�'�Y�;<�� �a�����Oz���Qދ/4���{�yOV��	����K�rʽ�}IP�}�FTv�K6i0�=yfS��b���cH�2�ːf�s������X��Ӱq^%��ؐt�.�ai��"����������)���@b΁k+Ǝ�D+�ك���:$N�!�3�oF�]6�����W��a�nB�uU�ĥ͞=@
�=��q}Պ6��wn��|0�em�I�CM`q�c�w�q�a7Ԛ��6��t�Cٕ!n%�.��-qUj�����̐���HD,=
}+��q����<k���n5'��'k�b��<j�v�Epz-�AG��v>ty�FUiC��;n�.׌ʦk�ӫufz���[Lռ̲=P2�̲��cK�^\i8���86���CK��=R�(����һ�C��XK��{�rٕ�}-���?}�	aP��
�m�F7j��VDU`*��H}����D]g�� �/W�:|��F�:ʺ��ho���i�C3��sp�S��+��k����󔊙�3�y��k�#bҺrx��}a��9�����W�m��|_�ef!�g�>���7#�_Oa�N��
!��3Q6��Q��&=�ե�k�`���U]��A�C�:�����~��ޫ�Yz��Y��j'�
V�=x�'���2����z<�F�E7�}�Nǭ��X��Ze�5��^�����+8h��Ј�m��*��+���N9}����-�p���H�Cf������VPsr�����	�<,Y�zj]�m������{!_@���Z��-+�ڵ�m����j�w���;̭����^���յ�g�>g.#��0���>D=W�G���e���pʯ�Oi�_���-���X�7��hPs��_�n��t\!�V�����2�neˠ&���{�GG�N�9ջ�L�@{\վ���`!��}A�Jm���8
6��@-z}�&��f��,f�\T�$o�J�4�<.�i�b�
�zۀ�z1T��D�MM+��̛��ǃ	�j0�I<��'<W�p���q�����U�n��yg��OEn�*W��`R"t��=ѩ0��`vH�	�#y�q���Z�VE=1�[O^։S<�͍<����j����J���������c=�2�Ǚ���Z�=�A�e�T��s��q%��Rx:�`�"��wl�V�b�Q����gG���N�T�^�dW�-6$�f�������A�S&�n	��Q-iL>�.6,*�D�4u[���+�k�p:7�R���*�"�R\�����e�Z	k±s����hzOsF��+A���i���\�W���ԫ�K����A$\��5��y�N����lu�,��Z�{6�Ed�:;�i�]$�|���4��vN�%l����X���j�4�1�!F��s��+���)�Z�NS�X�)�	ҽF��|��#�g�L1w>;�yNފ�6�~5���6�%n�m��o�?�sN7Q"�z�y S��$_�&_���Q�1 t��XHW`�@�XK:�n�;]f�gb�go����-v�k֟��"���7�u�=���U�(�Sخ!|<�ΩEV;�vPU���z�.�~P��Q)������ܧw�ʖ�b���]M���e�F�B`��Yec����������|�޺�|�T�ܭA�K��i�u^g�Ƒ�܎:t�-7W

���^c��z����`���hy=P��tϕ���#`��k�����P�5�Y�� �{�(ZgF��7x秠y��H���B�4��Jnw\��Ѕc1������g)5p��R����#J)�]��o�OW���]+�	7�@���U���o�w^%s�<-�-�!�b����Ϯ5`�Y�TQP�ܭ��5\����z���]�Ik�v�S>�>�yB(t�!Ӣ��B���mz��j0��ި�"��R��4�z�p��Nnܭ�h�p���s%�k��66"���L�&�cÛ��v�̢�.��E�̹�PW�c��N��������.��e<� �Vn�$��ϴuq�wVW�+���V)Yk
���ƪ#��z��(MCuE͢ D`��@��Ţai�ɨJa]YKc\a~Ƴ�U�R���3�>�8�]�B6z8):<<5ڰ�(��u�<|4�6s
ژ��Z�e�k�'
L��wm>W��!�Դ�CSd�smA���R#����Vʚ��Ϧ�լ�V=J*�����ӳ�������i�w�j�p��P��Z&(n�ܭۣA�J�Ʌ<�Gz�3�mXdV�{JǇ��C�����ouT���q9�$���7��,v�7)e/�4��C�'hd�l,��y]�L�d�|,:���n��A	��9`�\���O�n_B��%�rb�{��)��:���Fb�Qz�6����
�=�>���ͨU��\&�b��S�����"��l����J�6�tv����u�-6Eu���_+��>`�Uaok���<.�Z����?G�0J�;5���۷����?^7��s����ًD��rd���>�-s��7����/(7Y�W�ñ�����Js�(2Vk7a���ڜ�Q�ǘp���U߉�w���E�?NKM�Q���*�T��M�3��1��.;E���A�C<���c�=�[�M�2]s[;�t��Z�q���zDWX�w�.V�&|��
������*NԬ<��[0�¥��Q�s�`��Q^�+�1N�rvP���:�3��"��5��S��ȴ�9�oH�ᳬ���kH�S�g<wS)y�<a'�'����ɓǬ�՗�W���gݩ�6�#�"�C�����}U犣�t���.S�R[>P<��*R2K��YT~�ȼ�w��S�¹g�m��`�L���~`��޸����La%Z���:Pa#�Ǌt���Q��{�w���Q�N_:W-����j��Z�~�\�����<�!N���� 3�U\�z���UE��H,+@��+zp�[A����V�"i�)�SLE͞.�B�}b�e����y��M�� ��`��5.7^+���t�:���o�5i
䥷C�q�f�`p7um7�)��^�jz��DwJI�0y�=���������x}��@=O�ɯxa�2	��K��",	�L}PUS�i��ώۦ�^3>f�-?��
��|$�W���e�Z���&3�A9`a~�f���1��]Ey�8�����*�؜�Vǫvw�^<��&_�ǋ��{5�n6��h��ua.����*��Dc��Oa�1���J��A��'-�%�.��i�.Y�N�{7]ly�`�������Fm��(�=���2>��P��]]A	�	�E�A\[y���+�pń-�����y�ty�^yz�W��XQD]{9�b�3���P6�#����RQ�
Ќ\6���� =�Ï��l|
�x�z�=�0i��h����+؅|��V�e��#%Kp,�U��-��n��Q���3�A�#�Jߪ�+F�-�H��J�#�����C����s�=P=�U�aF���%cXv�Qh�l���v�
eq�#~�\�頉K_;�
k.)�y
�>��47���+v���ol\n'��
��Zς�����I��%��dd�+�rv)�St޾�|by�3�����-[^�~���r����t�qek��5�?u�I�3�\�yJpKZ���oW��Ѯ*d�a��'+�jW�?����;�#Q��i`
�څ;[�����ŋ$���B��<`������&�+g$}A�ƙ~����d���D��X��N��f,�w81Z�'�|�qf���`}R�^��d;�����j�U���'�0�eÂ@� ��ױ6W�s����r������H��ױ\q��ʽ�Uͻ�	�}=�䌫U=S���% ;~^m܃κ�9��I�� �Q���:����}��vБ�G�C�F�C��dw'-��B�~Į�n�Y��˹�/�\��ہ�r��/�0�m>��^��j�R�mk���CͲ�ռ<�w|�ƛ2�y8면��X�7n9�=1G@ov��xu�zt���[\c��ӳӨ�����󭶷���՚QA���Nj��q�O�m��c�X�jfz+#�3�y�poy��l��F���ڰ�IN�meX��ۮ��wbO��໵*���8���xӹ3���*��N��3�c�7�V	�h��+/\�s�ڗ��:�Wr$��e��(�{RPD䮙1��F���t�
�y�i˳�G�3B{F����L��޷�*%N�9K��1x�a��#���1�$2�+�;e�ٴ�G}�
����2,��=�r���QS�z����>X�;���:_��Y�"�f*���El�2�[i��o2�|�J˂I6=��7|�[�Wm�J=��f��"�V�8�q@��f
\���r�$B��'EmaOV�=z�V��Y�c�wo}P��W�i��<F�w�q�)0��n<���`�e���.>Ug�%��\4���dwk۠[z��s�Ujx��ۣ{C�1>��?q��ѹ��n}�s۔@��S���a�-��a�{��p���ed{a�G.���l�#�ʻKY��or<*"^]��F�֍֜�%攟��l�,�aw_v���s�W�=���.�\�������t�tg Fi뚆,�^̺Twa�$iik����B�ϻ��Sm0����̅[�c�Ŵ'WU�,�Jכ9%2p�/ �ˣ;O]�-�A�QZ%�Y�\��I�m2����iڥ�7�Y��N4vZȖ���������X��*G�YۛnL�Ƕp�����эӓy��ŸW��4��ې�hBsT�����}0�L�l��Jdx���+.��� ���,�B�HV+���==֛c�;Ou	Ի ړ�XwW�.C�3����>;���6*8-��6���Ǖ��˞��}�|��[�/q^km��Kgs�%���ǃ��.<��`�k�~��zk��wR�DXj�0��0�|�֧��:�2��v�اG�9�����b�^9Vh�q���Q�
�O���[�}�Di�oW�"	�{��cVY���fo�����C�98�����(Rw�^ Ήd�M!��d�c����!�D�:5%�BmB��n)�o3~��{��J�<�f��Q��m�-�w.g��{�]H���R�C�y��%��0y]L@F�ئ+���NR*�xW+���x��8�L��),J���Nn�'Z��nAz"��G\z�@.��ICW! bSs����/�/ޝ�E��W|<),*/ЧW��{.�;�z�	c�ٜ���Ǔ�G �
N:��1F��iuJr�D$�%�]UŐs��9�e�SHѹ;��\���P��,���f�-;����t�*�L�T�$�h��%t�,�U�8U$f&�B"Zds�nI6��	�$a��F���{�	eE�Q\�Q6��KJ�"�AuK�	�E�眼�5#L(��%�X��PQ��W4а�EBl��k.h$�`�(K�#D�BY&�f�+(+J�DҰ�!#Ow9�E&�I�\���<��g� �D�(�dQ�I7!���M-0��YQ�"��(I�+wnʜ�JIj,��MNt����A��9�)C	Gt��U	���n	�9�ަH������Y�N]r}1Y�қ.s46S;:����B&�3���Q��H���U���Ft�����z�?B��'�|,������U?���P����l�w��h��$����t}�m��'!�r���7�C���?���޼.��@�Es�}�l��y#K]W�e]|��Ι�̓�G>�"	#���#�A>ݹ;��߼����j����O���]�=<v��$;�r�L���9������yO���&��w���AG�璒<	'��yS5��;]S�
~=�]����@�< ;&�dA�������'�|v�ߓ{�w�i;����{�SzBI߿A���1;��x���zM���L>�۝�v��9�8�|>&F�D�� ޴��|��]��d�V��A��0�@� �5x>��A��>�#��|(} Q�'�����7�99��ϭ��m�<��I�����o(�Bw��v�ՂM:~qD#��'��$����@��;dH�<zj{��7��G���y{�*��^�A'��|�� *^�b�����0|;�=dQ���?�Y��"�/��x�E��s����x�l�w��=|� Y Q��G�I�b��P�7�w��v��F_�~�? 8���@|����z?8����� '��}v��I${� ���"	 o�xAdp��R"��G��������x�}��ԗ������ �H�����o��f,��%V����_#��<�7���dIdA��nw����y(��
�ㅟn=�ɇ�y�	��|v�<�RvyB�+������*����	dA�y��<����c���Mo����d{�2@�I�y}��#xa�O�'��G��"�G�!�����s��?�n��aw�=��;����U�w���Гy<A�#~B��z�� B>�""rx���c�ݓ4�*�_s�q���0�@���#Կli���eɯw�o��������� �"������������"�{�}�z�B�A�=��į'̏a����iG�>��#�$�I���L؝����C�v���>��}�A 2�3�x�l�wžq�	'ogϟ�o.��ۿ@s�~�ޓ
��k�~�>!&q�������]�o����ݼ<���\�����O=mɾ�>��5������neWq%P��Z[�c��K{�,�7�ـ�l�k��H�3ݟ.�~�4�Mm�]������ڵ	������Z���a�"���j!��#c�ݫ�̎m�ܔ'���l�J۴��Xv���ɷ�V��b`�j���Lt��;ԟ9�GwM�u9�߷'z�N����<[|'���<��o��I�N��xp}d�=g���0�'��O�9>�����`�}O�9>#��E��H}`C�#gÈ|��hG��>>�}�돶3$�K$�1����̾����#�#�!�^�gÈ�>D �A�����zf<#�x�O {�-Ǽ� ?<�C#�G�����$}�#�}�2q�Y������9�\�v��}'�<	t@@D{H�M�F�99���u� $�q��??��I��x~�'��������ۑ��}�@Br����Y�������{��򯪭&zn����J�_\�D�y�y3{HV��<��0~��ӿ'���ϳ�p{O.9�S�z�PP��]�	���t���Sy@�C�[�;��n�m����������
1=]+ύlu{d�u��5��I��y�c�E����|4}�
 !>�"/��$z�}D41;ü����ͷ?����9ӵ[Oԟ�p2���S�A������y���|\������z��O��| ����{�,�@�?H�|��/F '������G�}�XG�ސ9'|O_�v<��I�'��<'�n{�b|��yv�����]mΝ�p�u.-jd��o���~����#H}P}D`������9ɯw��s�!�܇��dD�O���O����ȃ�2>�#|BM�	=~�<z��N~������'y������v�	w�	�<���N�L�p�On�q��� AR��oi�ޝ�&��ǁ��xv�5�|B��a�P��Ag�#���B墳c����<��ra~}��?'���@�� �0����#�����K��o���]J�^�b>��4G��{����ŷ|����<&|C�n���L>w���o*�nӽ,}O	�����XP>��v������aM�	��ޢ*P�G�����^��H�=��}Tv|�N�'3m������q�>�K�F�%	�����݋�S��o�����NL.�����oiɅ<��7�ۏhs�G��	2�O���@�}��T-T�Ͻ �G�>���W� ��$��O�e�U�F�M��6f6���+�`��)	Zή꙰�+F� �S;��mJ<��K��m���WR�?U׷fJ�bŬ^)�vI٠�4wy�-��vq(��+!�r 2��Ɂ6���ԭ�|U�7���:3ϴ���M,sO�S:ϩ�:���:ܳ�N��=H�G��
!y�� ���.��'�����~��<;˴�����<���W�I�''!���]�1;��'���0���ͽ�˿8�Nv�)z	>@D{	0�f��i���~}t]�6go���1q�<���Y |B>13��g�m�"��"~^_���P���|O�=��zv�~�Ǵ�;s�{q��x@��[{w-`�~wǐg� N!�����?
��p����k�W������'8?y�ߜ~Nq��NO� I�����G,����\Ϩ���z$����޿[w�|>��zOI�S�z?�v<���@�C�=;r����>�"H��a�쪑��;d\ng����䟎���7�~�x};yN��}�K���@��}���^�=��
�yyM���h�>�]��| �}���|D�O��"����#H�x��c�QMe瘰�r�o�|{�>�4�Hs�j���~���u�Rw�J;ſ���O��?;x�N�w�}C�N�^�ֽ�xw�i?&��ֹ�<	�>�4�g����D�`��zH�#� �Ϣf����eC��Y����4���C�iP��D�H�������>'8���+�	7���S���q�����N�y�<'��8��6���K����xM�	����O��}��G���UCM�?t+>������aOC��N�����(��m��Œ|#�i�b\xY�|�DG�o8�}Nv���rs�w����aWe��|C��w;��7 0$��#�kބ��̉���ΰjk��ˮ�߀D�I#�=����=�#��@|}�$�O���(�������z���g� aI��}z�	6���l^t�V���>x��|v�	/A��=K�k�&<��?�����{s?
(�W  ��&G�>���/ծG�G�>�/�.| �#�D��<+�&��>!���x�$��<����d$#�>�_@k���@�$���#�	g����a�e({�鏽Y}�u͍������#�"8��Hq�D��7��v��9����M�?�H��鏫L}G(��w����܅��UMI��$u����۷EDk���허dB5��r4��hv����ś��%��xG(�*�j�qaVa�Q˞���[�S��M��_c�^�h��o[�v��P����0�C��o��fe��9�rX�M�����v�g����u :�;�2frfP��oN98�0D����_dI�O@f��q���t�:�ķҚ`$+���4�Q������,��Њ�=RE����X\)�؄M�#si49k^��D�mACj�9F�x��: ;�o:���EnY��
�Az�-�#�rT�Ķ��&����T��T3�"r���B�|�G�d�{�$�x86���]W��t�ؗ�B>�1Q#�V�=��{b�G�Ǆ�]F�ٮ��PM��+�ع�g�ׅhF.q.�K�Y⋢��ݟw��o����a�p�E�^���_18�؆gn��7ʵYL�$�\���y��kEh�P�c%	�k�-+܎'kXf����o9Ƭ=͹	�ڪ�J���i-�f x�l���v��N�|�uf���A���t)��L���n�I�窷�lϛ��Y�N�8"���|T���q۔1�Z|h�����������<@{�I)��LB�uZ<3�e�_<L���� �kpѓ~^�^��O�������&�kE��hR�=��!�
J]O��'g0i����w`�]���4U[���{Z�=,��J�Hų�u�;�(Sɵ���8]Ox�������>���v+3��YmD۽�p����h�����-|�tjtu�b��+�.]�Ѽ}�3����0q���KJ�p�]��C��=,���i��X*V�`�Ò:�ɏ3�͓7|�?=�n�CRPh�BA��;L��,�>�������)�ca\�j���bu��j����Wd��\@))����Gtyg�8�f��uܳϡb��^�B�\m�P��n�C�=��<����G�'\�H#�3呯bl�@�s�����>gF�^kO���ܪ5M��n�Lݠ�P���7 �>�/�	�J��#�+r�.Sݺ�_���v���E^�q��@�탒
�e'��@C�b(D<gځ=�BD�8�}T+����[�Y6�{�q��~�5��9)��Ja�Q��Q0�S)to�)غ�-��V���>�<�/*!r��a�1md�;k=���w�Q�\ҕ�m�:�g�H�a��q�����K�Vxzs(b�}�z�ǅ��T��Sb�=+�ں��a�iH���Rr'�Eű&3Tb/q�b)J����O@5��+�+�W�ؼ(�ֶ�-�̛�t����l{�w:Ń��,�Bd����%ۣ=yѽ*�/�em��˪����C[�OpcP���K^�������x�B��Oer�ƕX���]SgD����*k������=��hh�Q�Y��>ۡ4i{�U-u�v�%�v9}��*���]��}�qq��oj����vk�U�.��[��1��d^!NM*�R�j���N���SB1������9iT�f�W!~y��m`�w"d+�:�38�ȼEK��q��ǳ+�s��k�w�ˣS�e��Z�Q��V�frT�ډ%���}���Ǖ�m�j�j4�`ĝ��Ng�u��1���u�W�k�-�
[Qw��}�I�g�^�G�l��=v���Z:4�ʥ>@ha\v�o�`����=>��q,���3e��V��uM�B`X�o�q���4�=�]Gpϴ<.x���-cG$��Ý���>��KE����0��ᤞ�+ _�<%4��Ih�_ǹ;���k7z8Ķ8N�3������UZr���ҭO��A�\��ռ�����0.���o�랹���&l��6Յ�Y�y��r�q�/Vcr�r����r�Ć�S��I<`aA%P߫g��amy�x��֚�^Ek��n׫��riY� �&ʠ9�Gh:�)����c԰T^\��h�k3��Z���qf�ݸ�j��u/L4d�J_Ӂ���ҍ�p_��l�(׋�^����k�B�[��+=咖d�6+�ht+���ѩ�ι����Ue`��[Aa�o���:c��M��6z����crDS?�U_}�Oς��>�Fi�p�aR[m�hc��is1D�smAV,9�޼�bf���#�=�y";�p5�� ��N�����!YZjLV���.b<�S�����)�:���^�f�:�#��]���U�.^��Q��=>�� =���}��Ϯ��]�`r^�-hex��u��?�x�cv���Η�ٌ�d��V˓v���l�I��a�)�u��Ij\\cq$H|n`��Z�f�b� �Y+�x"�Y4�T>uԯo�^����(�԰�$�h<�fu�����Pz����k՞�o3ؖ�:��Ӛ|1ZZ}L��;URw��\���t�6���U�c��ȚC�M^�n�>��PϷ5�~9'N��P�?"nO��H{0��ݏG���е�x�^5.�� �j��3�7�T7w�(=��E�W�Tb�A#���j��ΠL��֘�]�����j)g���d���_�lz_'PoncR�/v��4&!�O +�v68vs� ���72v�o[T>�_�ݡ������u��eL���qvU��]��_9@�N�灏'垙q(������*J�đ� �+:�Nh�2�k�.�@�=�h$w�9����M[��b���>L�TyMQ�)lq�+��U������d��ۇ'8�� q��<^�u^x���:zҰ8o �>��A]�;�'�����b�k>N�t�%�#�>���J���L���g��|6����aP�����: X	�܀l��d�r>��h��P��U��q�#8D��^��z`���㖍U:�W���"-c�Z�'/lW�������Np#�iGb�q��M�e^.�u�*����-��*�e>[-���[�4�6&##fV�#A'$��B��0ǯ�P������[Eڋ�;(�zމQ=�n��Oי^�:Q�>FV�GtI�T�"��I���_niւ��T�~�)�J��>=��D�%���d�DQ1��O�L�ZQz�m�k��2��^�������r��������}5
�o�(Ϲ�'�Q&�86��Hiu��R[Oc���J��(;^�	��h��R���׋�%���\!\�ۙ7A쬈�A��%R;�:q�YUi#7�ו �O�Q*�=T�%�LO���L�1F�z��*����'��߇��z�c�0����.ڳ��[��x[졋�r��5ҀBjEIx�/��&m�ө�O���n���RL�O�%f��\���Җn���NٴE��ci�+��=�Xhި��9���o���V���U�x�P�DQR�ޏ�>��.-^�_���<la5?|kF��r7��R�d��q�xס�K����:�Z�zjgVm��yЄnw�G�ef xU�[C+��A֜Ņ���f���Mw Ɖr+��]Ol�[{�sn�~�|��{1o���{������ܣി� =���Co=O��dZC7M��^��8�	��[��r��s:l��^�<�;~�Ԗ�H�Ek���BL���g�=}��d�����[S�2�Y�-*8C.�j����[Uڌ����Z%�'��Zҩ�xo���$��׽;���Ѥ4SGF�p�g|�3�jK/�cUi��dh��������9^�J4�8Z�!K	�ѥH+��W� kT�O����>�;H�5'
aݏ>�=��oM��W	z��X�W*��ސi0P�Iůbs��"��8OmxݤQԛ�u]��O67+���-4��;�P��-Pc����-O"���^]өP	.��fP� YV��/b�.��%*�/d�ｋg���K��':v"�:A=�% ��4�mߨs~����>s����&�g2w�j��=s��|��]�J�&,�2if�#�,�]��망�ϝlu�H�?^	��L�o{5�+��G//svE�@MP-�v��P�\'���j�^JH�.s�ۼr�@k����/��-z��!���B�YG�U�}U�q��ٽx�>1�06��u�!�>��Jv\�e"I��eTtӈ
#�nqħ�L�+ͽE��c�}�w�N�咫ź�{��;˚R�6�w�����ݟOj�R��_��&|�<��=�����\>��Ӱ�}��]��[��u�:�B���K�`���b:�T�p�)$��YEiQ�$� o��s,Lx*1��V�/
,u��-��I���h׶�q6����,s��|��U�d�Ja�������t-}��n�t�j����`���~������0��{��J�,�)�/\[�#[��sS���ex�Chy���yu*Oc��N
�.D�;����Jba�'=�lzUT0-L1粟�.�O-�|ּx �U��`�Z9n���s�R��2����˪�:����I��:�XW��q�fPn��Μ���un����>N�Ξ���D��v�'��ݘ�R��n*��)���3����aGw�s�-��aoH>�\(�Q_�p�
��Z�$}��+j��}�9h�U��ڧչ`�Ck��mp� y/���B�����^��
P|�_G4o���Û+��_��r��ӫm�2���1}r��Q�0>ԍ�e��֢�E��p����b=ٗ�9�!Cqw	7�Rg/&�Ղ�Þ�q�ʐ���K�#�ǎ�=[]��,r�qR۶��$�h꺉WM���w'}��-�z1�q;�'��=I&c��J���>���ySkݞP���^oI�5��L�����EK�7�(��mWy��*�ܣ�p���>���2s���ە6gsn���rto6N�9`u��q�[j�q�f�i|����(mLv�5+�z���ʣ'�p��7�q��N��L�h�N��E��[���X�LQ��8�]��w�gKG�����j� ��tH�5=6����t%kV��wQXt���'U�N��rh���g��|�n����m;��#G�T���j��d���!��s��x�|��QZa�!%����k��CW6q0}kR�粷�L�a曰3CGY��=�r؇,u�w��2�c�4Mo*+��h�ݞ̆XuG�_P��gZ����gSۖ��p$&�I��ă�q�����G���u�S��M�o�#E��S���l40�P�؆L2��岍[Dq�wt{*��8�w��mt���]FMBPx�ڑ��;�J�Xsx2-w;e<)ij�����{8��ES[M����FV��E9H���]���y��5�t+�^��(Ahf�� l7����0,��u�a�#ʳ{aW�:�pmح�<�j\�!��ŝ1]��N#��:v*�n��o+QJn� <7��;��6�wfE$�i-�˷����E?���O6��1a�EmM��\AK�a\�j�\�[�v�����F�t��b�H��iu��=��[�1e�ޞE:��->��學�m ���jʍ��澘jCn�Z[�J���]�ӭ���G���1ZM�3���>wz��\j������'%��]n��wn��A�� �k2/��پ����ˠ����~T����\G��hE!qg=�]#�p����;���Ð�>��z���I��z+F��
ٻOXO&e����뼓[��N�
�2��F�d:*���[��t8A�~ܞ�8��0u��V�i���y)a�P��U���*V_TY ��5��B@�*J߸�4��A8�\_%��A���낆nm.W�͸����Sܯ7=N��f��o0����[��;�[�����y�����2Xx-��q�s����rU�E���B��Σ��M���\kz�W�v��t#��/�=�W��p�7r#4�y�,r���%��v	�}��a������1��@׋�!��z߫�y�w��N����KC7�!�;qp��o�9�B�8�)��k��(�U��f0ۖ��g��%�H�jJ�HHG|�,Y/.�(Ԧ��(ͯ�����t�k����Yx�n�k�  �@ A��T|N���i�*��Z*I&���r%3mP��A*��r�Eu)J*H�g��e,6e%VW#�-B��a��B�Q�V��&s$ʒMS���<��f�r̔Q6ҋA"�J����:E�WaU���9�)���e�٢�*e��tĢ�ȧf���T�'T.RID+�9T�$�<�8Z���2���\B֘p�R�I"��b��[H*�є\�d�l�g�Y��2J�$���+�L���\��3:t���E�Z��U�.��	$�URj�!.(J�Yhl�Z�tS4Ģ+�����������TFAjˆ���J�)D*9�Y��aR�4�*�TTIH����(��v�C�Vm1j� E�[�p��R�AIXX���DB��
*$G0�r/"+X������ߕ��[�K$A�ھ�6�}8-�Ȣ�5C�x�E�C8;:�������H~�jJ7�(K�Ĉ�W���~���� |����\�{쀍�X��6�ۇ��GI(҄�)�Ѯ��	�&�l$Q���V2��B>e�ơ�w�}E��j�3`�@Qr�@f-X�n��r�%T����t*���!�g�i����1�G9S�܄�q�ne8�D��9W����L�K�b��v�<j}`�z�ݛ��N;�8�!�8ɲ�ɻ#m�X���J	��~�.[����B���!������3w➩7��ݴ�XN���]mM�qy�p\ɽ��iYC��rDnφ8�x!t8m�v{���:|{KF�ow��i�s���#�ͭ
!S�QqZ���_{����_k!�K�ՉK���Tk����0X�8=�&���)�KR���"�؉�]r�Q��܃#a���;hh}��H��^fFzL�\���"�:pĪ,g9�/����%�E�H�>70F��T^����d��%�^Rz$�%��h��W�H>Qg�X�x��cbU1[������=p������5<W8^f�;�hF�Ld�+�\�ʭ׳��/�sܸ�l���k7md�髍z�����_v%�}qӮ�f��'(�.�ܫ7n1]D�����Cĥok;w5uJYJ����j��r0��=Ѥ��^l�Yu>nu�v��q�NN!�o�f3��}��V����ߖ�?��kV�Gp�eVj�5�U��T�o��{hc��΅n��n��x���'�D�ʚ*_�`A��ko��Ҍ؏������ǣ�[�CW=��c$�g9]����wB�tvtT�WucB��µzH�+��*1q�.$��xCV�o�U[�Wyx:������t���K~���[���Z�}s��Fhݨ��51U	�$q��9��{y�E�v��YӬ�Vlc������B:�OIr��R[!@��9FgT)�묶��~�����3����?g�<V�C*ܒ�U��;a�םb�K����O�����kf�u�����Й�Py���E�����a�����ӭR�ys۫6b�m�����!��:�b	�/�kH�;
�8[�-��W�ح�G_�j���W��LΣ�e|���:���������z�}��|8ea]#��x�*��7{��v�G\�M!Z��u�)ӡ#�\-I�1���P{����>��qy�D��L����z�4�v�ɜ�80�+�bʜ&�qeq5k�㝒�{GF����39)�8���GaYtOJ\�/	%N�.��ܫY�Q��p�~�Ut�ՌwW\cJ1�d�&��q�`ed6�<*]c�P1ujH���y��J2U� ��m���4��_J2-k��nu'`�d�DQ0ܳ��\*V_�"-��Λ��fs
��=�PH����4��g]q��\o�(���O��Y��0�CK�������1�秣<��"���E0&����6�]�H%U�09��Z���a1/s��8�$����=3��R��w޵�1ج��9��bxmQe��ey�+�Z�ޛLRr�cf�vG�����%����<�^:M[5�Z�Қ��&^��Lk�ǥ�x}9b�2��+he��eC�iN<�>�ܘݼ�5>-X�h	U�
�������Y��E���W��]1�S��f�J*�v�~s"��q�ź�e���s�!��ύݻ�~�\Ձ� �Dfdʾ����� )н *�s���9du3��[�K�ʃ�*5%����=���CJ��O�^�Zn�q$kR`�R;&Y���-*e�·4(9�g:*t�̈^l!�cG:b�gn���)+J�e�� �����	w��>�jK>�^F��@L��
���WX��{vnc���~u�uٽYbZ5���+B��w��V�]9�S����8��L�����"��Oq�N�o�O�p�\K�1�S8�k�5vͽ齻�u��=W]���u�4�{ظ�-�`70s}:ĝ�F�c�!��">��٫���[aO���3�r|�G�`�iRS�Bb�^���<.�i��UUL'�Hw�����׳��[]��#\�C�U)���Q��$�Z�'
� 
�8`�DgX�(<O��:��ާ�n���|�����Jې�h�<�!���A}>0N�u"F3P
�E��]�i;�b��t	����j�9C��œ��؊�xϵ}ݱX���r��ة���Z1:�>e9[�2�c�v����Ҟnt�`���Ł-ݰnU[��U&ֵ�4�Pi ��B������-�9�=y��yw�g��=�.�Z2ʳj�f�~޽�]!HV[��+�
c	ym����l�z�Hݫ�׼�
�y��8pUa��hf�S�����X%@��m�˄��D��@jWd
�p�Y����a���48v�+�k*��7�%C|�6�.�f/t'깊ZZW���>*��MW������&�mvX^\���;���ѱ�����������(R��_����(�S��W!��~�?�����Me[5�8�]Z�F��O�*�Ҭβ�������9v�b�ʹ�����8�Z�V�9r��˛2hyw ���R�]�y���Y��dn��yئ��+�@�]����٭7vp]�q/��XV�y�ZH���Ә���㌚߼ ���uoc��Z�����Bm.��}���L�O �<��<�"���<�x(�p@+N�x���O���Y�󱩅!З3�� �J�`�<I�n�֚�U�z�i��ǍD�<^N�w1���[�8v�FǪZ>4��KF��T��'L�+��׍􃫊i���9�1�zR� �|jv�_����۽c�;:�x������Ep���	o-�rb����􊦑u�^4'^_��M���.�W�<�[�l.�����3�R\V��\9%�|�KbW�rP�y����Խ�v$5Rǅ�%�d3�,h>4ݻ�K88Wϻ����ݷh&6��5�k$���VRzs�����)�}+D�o�sބoW<��ϓ��'�̧Ȓx���+&���x(}�P�or��p=�Q��'ϡ�r��>V�&ʮn���#Q�(�95����9��J�B[��$ _-"}�3v
z��:Gv��ZC<�SK�J�qB�!:$��Ӈ��W$��7�
耎���&���~<vА�xlsE�����z�)�!k�G2C�^⎡�׹L�a��A__[��[��m�o�OB�V���t�[ƺ��"����d�\o}�rQ��\4�B[�^{���ң���Lo펦G]ǏM%%�@g,�����Tq��Zm�7v��V;��7�t���� �����m�C��WV._��55)׼͐{�������i��ub.^�\J�KnU@ê\*�ЯUN���:�,��q'��G��znAهpJ�g�e�����=9� �/(��W�,V�V= L����u���Sʘ��A��%�'KA��N-������xp�*9�ٕުվ`�t�P�TU� ;9	:y2�f���`��T��S��|�w�d�*Hy�?�L�����BS�Wloh5�5�x�V����M�f��ߴ��P	i,'�2�;m��߭7)/���(͉O������F�b�:�/c�z���q�K�{�#��i��Lv 5tn�ep��V���:\����3����nc ��opˍim�T �d�\D5�o �t��(�K}���F�_t&u���yV��}�KwsP��z��D�~�K;g9՛��չ��ê��B:�OZV�)�%�x=|NT�}v�Obo�_�Sy�g{D4�ʾ(��it�H��x��&�W��/��9�su�X�{7)�f&ǉ�T�����żK����`W�;��տ_ڮ�E6"�'d�۳Ϲd�p��.�NSkL�fVQ麁���oAS*�Js&:����Ф�A}$��<p�����������s�I�'��˛�yNr���9.a���ո��Ӗ�u�����v��S����{�xx*r3���q�n��XL���A#QFt�}�\H(휄�Z}a���f��0�b0�P}�M�N	��oTYDO�#�Ϣ	�� �(kZE;z��`9t�U�v �<�J�{�sW���}ݮ��V]�7�~���<	#4NG�ב&9k\vF�s�.��g�W�{U�<��.�Kw�x�I
䥷^�:�C���u��X\�L�^!'Fk{��hݶ�/���浯O7:��\2q�"I�ܳ���,�-�Sˍ2*��/+��TBj���[>f�Zun�R�����8��_Q�p����5�pm�ъ�h�h�ؽ�Z��\��9�VF�!f�QY���9%��"ۈ5�.��:91�!��=t�ip���g�Ry�Z���h���
�{Ջ���)unz���_�I{Ǎ����2�ʬ2����k�P�c�5~??�b�����*�������k�9}Ӵ�����j�ĵݞ�[�Qʸ�U�@���=\vj&�reV�,$�a��{7��cӟ��m+W�SK�40{"*�W_j-I�kRa�I� sox�����T��;�Q�i�ΊY�4R�������=�6���"�;�s�ւXU}V��woZ���t�����q���]�!-\�oat���NPt[�;�I��xxx ��v�S�֬i?umiF��|�s"���>�Z�4�{�Q�M%Ɍ��ۺ���aRJ�n�zޮ<�v�����^���H��Ln��q2ᑮ1ٵ�s?o�3�4@W��&5�Ou�νw����?BW�k;&Y�Ja�:��(t���^�5�F�*�[s�C�o{�wm�3����X�]=1H�BgyP<c�Oc����O��T�D�o���i'	�i�h�1a�ٽ+�gf�JH"`�4�6JbI�fWgþ�οZ�h�݊b!�+#c��.|L�e�7�b�^�\�܆C�0��pD�ђ���*�]N����/�h�gu��/��z�յ�-��J��Aj�*yzCpS�D��p��ԣ�7;<5S\���F��꼧���^�}\o�.u�~ha����%9t#= �i�;H*�f���G'�9Y��Ï���U	Z�e�c��������Jv��b�n���1��"�{hݬ]uT@e��/W���a��T.�#u��퐌�G4�W�rN��}���q�JjHE��}��������}5��|!P���Lׁ]�+�pc炉��)��B�|�3��;�dr\Gf_�_T�д��漢�Jj٭�y��T��	�\�$��J�o-�Z��]d������˰�q�6TH���/Qߠ�d�_�DG���EO'%��ە�㢠
���]�S���m���;U�ú�����$`�-i�폺�޻���}����^��Os8Q.���Wd���
���V8M���G�틤�7�b��o^Qņ�'�Ň�I�.�3^n��}W1KKJ��{g���:�0=`����LZ��u֬o�:��S#���V����rb�~����9iUL`7b�������T��D�n���8�gб��$���f�C6~�Z���{.�T��g�5�����9��$*i�rYl	sٞCF=�~�n�R�z�\p;Eq'uƴ�:�3��H̼�\�Ȏ�e�Y鴽뎠�����h�<	`�������^(_:�α���}��M�3o{gB���ǫ�^�j��!5�[��AR��6���rb���TK��˭���Awov�Σ�zxݸ�o�<кs����G-It�Lx���	�{�buV��yl7�a�~���L3f����*����Rn\�z�W*��ހ�`=�Ɉ���񬎷�^�U��M�#�潳���R�b��u��f����wW1����]��X�㦟:�۵��/U;�XJ�'��*��1�I�n�Gu{�67�
�#*VB��gq\v9ذx�r��Ր�*6��W����y���feYՠ�u���W��U|����`����z}u��_d�9������CtF#o&�rP��K�gfO�ׅ:�*���,� ��}�N��P�v��Gf�{����qC�n2l��7Hǒ��(�_��+��:��ˬ�`~�酻�(�O�.�͂�o��C��m���4C	����D��8��<��'=X]��������Gmbb�\��E7�+�3Q��B)��K5����i��J���b�����4&*=������]PK�tB�c���Zˮ۴Zo�DKy��Z*u�����Z�_/8sI�~<0�Y���	�{�~�xzS�߫3f�<Q��^�KՊy�^�>2{Z�W�}��+�X����W�}W`�2�[s��9�r�=V�߰�nyZ�=�8<���O�e�l~��M�fe���Y;��q~�m�B[BL���qnOZ����zx�잣�g��"�ؙ5��L��SM%��N�l�WE��(3���ƽ9}���v��.���?N��c��/��Ř�*�\�1�	8��6�ho�GPЗg���K/5�{�����rՙ�-
�y�іN�J�R�ɗ�������ͭP[˨�¤�P'۬2��Jֈ:싡EЧX����˾]-�fmZ����-��(�MV8[OT�u�����L���;7���b҇b�"mk,h�8�s��ғ�ݝ�c��+U'j���~ӏu���]J��L��q�~�6C6%�^>��f�Ò����L������5�a����|q����q^Ys��.��M4G��e�e��;�fW��dǳBķ)����ˑZ�����ᆸEvж��W�+%I�D�{gi)�p�/n��⁝4j'-��o�5q'�H���ӷ�������fV�w[(�uE�I#y���pbU�4�g="�hb���}��Q�����rU�`�cr�� ��t{ϨI��l��*��53�4��`��V��F���n�gz����Hr�B�t���}�R+��1�]-ڵ	շw��F�u�4��N�6u��m�/�}Y.�jr��A���"���5:��t�W
g���&�:@\��!j&�.�8B�,�Y@׷��E�Ѕ���s`�6���/{���%���i]�[)��kr9����-k��sS��Mw�r
�&��۽�ѰƧo>di��pX���N(�#,��7φ�*f����j^�V��4����;Es�2)���Z����i���ԭ|�^ztYôgBH� X���.��4�bV����ƙ��OC�s;&��2s/��b]�PT�ֺk&�.S�n�m�������s'����a啺�+L�L�g¯B�R��
�Ӝ-�[�z����ί��:�.�h�m�4�ה	1�9�.d��氕@O.1]�^r�b�%�G�g)v��[A+��J����}u��,���.WZYj����i�=�9���I���c�Pn��:X7V)�0sr-�U�m3i39��F�d�Sͫ�w���{{�)Nhcv���;xH�YL��/5+*�����$u���4�#fZg'�\͉o�����L�������x�}=�E��l%y����Kᕓ��hV�8�-إ�*
�-��6�@V�]�����T4�{[�s�=���:��Y}�Ņ��K��ȸ�-����=��=�I�쬜��� ��طK�Z�2���PJ�T[�U��rji�[8���q�R��T��	�����2����g��v�k�MWH��c0�A൙�܆��@��
ٛ��d��7�,�6z05���<� }��=�3�f��*�G�>Z���ˋ��Ma���%t�!6�ʸ�͒�9Z��3&�8�> �N���������3�ʬ�m����
sl����{:�-�yAk�q���iF�r/iI��d&Q��99�+aF�QL���(Y',�:�,@I2R�Q&�dqn��$JB��Rf��Rr:Y�)��e��ŤQ�V�3���$%[5�H�g�:�ȩ2��Q"2(EZ4���6*'�$�'! �
�u�r+�TZ���3�J$Y����¯%�T�s����UQ���+D����H*J��E�T3��.G+�tڡhbȪ�r&���W�Av�O2�LI,˹��(DĄ��'!ԫ�9	�UVIPPA�k���*��Q�hr��sr�C��wQ��9����V�3�+�*�I�p����S��"�;�Af�*/f"��P�CCHI�$�QX��r�܊����9�9B�D���Г
$Ψ�$
N��4�U&�UQ�G�Ă<��EA"�h���;˲��L�3��o4��ŝ�1fQ��N�[[���e�t�шr�i���Z���2�w���{�eb$Wz�� ����?y��NW"��O{��ҙ����$�M�9�s�/-=]���9��
�`��\�8d䔞�+�������힄q��#��f�[0�4ca���疞,��S���'���[�z�=�<���n%}�].��7��U�d{=毹��]Ru�I�w�RTV'�z�8~ط���O%��/˸��gy�An}����򯒯��r��R�֖5�z=��qI�̵���Bl�y�s���k�M��Ն0��Fkٰ���e!x���|r��/�I��~��3M�N�.�Ӿ��O������зO�U{�+^;�Dۄ�7���D��}^-�t�2۰\�k���{F���:=��C�����Ԧ�{�;>�Z��M�v�;F�[�(�f����޿{�S�o^���pk�4���ϳ��'ay15	��p���p7[�(*��|�K�Ԏ�r�_r��4�r��j���{�+#7����+[��w��E
�����W<0ұ	��d��耓@�� \2�E���U��;���Y���އ"I//�G��#Hl�v[)��ꛣ�j4fy���9eh=�"�Tl�ve������L������.��z��/a�*=<�J]������\,2�Um�6�l�yj�Cƫ�2�JK��l�)�է���=�g4EEg[������v�z���W=�x���֖����a�߫9Zߪ>��ye��HZ��k�Ot6��y�{���="~k�H<l�T8ק*Èt�Q�1�ମG��W;��Ȥ��=ޣ��諼��3� �M�}�]sՓ���y��>�w��&�k�m���:{ث}��퉚�.�>bV�� �Len^-�s�[-H8�N�J�T�_P8ٗ���s���ǰ��u�����}��Bd��:};j�I���w��?x�K�#�'��V{kOonq�.յ��T��K@C"�n��Ҩ�����:S	ա���~��l�kw�{ ;�rܷ�K�gr��{���)�)�1��"��G�=V��7��P���B��oopg�nf���LE�[�z�󭮾Y�r�;���^��M ������`bM�Rj�
n��i��u��WgC%�n�̀� �|�Z�4��\�+m�����*�mm)�����6�t����]���F�ݸG�q��vϊ�.��|��K'j�f��ov��E�o���u^/#�����y&�xT&��B!V�����
ս��:-��X���>��7��H�Nc}�RZ�oCP���n+�O�Nn}uzٗ/%�\�u�_�P�&ս�?e�ۋ�f3�7�T�{��ktS�a��	R�w;���kӬ�{��5{�V��Dw��2�޲��1��i[��y仰w��ś���������h���5� ���g�߫9y����M��}ײ�u�Y�6���ף����盌��j���7�K����J0�X����u�
�u�'�Z��&r�S��}3��/5�iEir6Yt�;��/�.��v?D�a�VC��=R/O�=F�<�;ŷ�Ύ��mX�*��*y�&��V����:.Dp{ ��|#ۯ[6!����\M,��>�i�Ie�r,A��j�~D���a'WrR<#!�o
�n������\5�-�]���5�ez���iȮ��[��Obw]}CcN�ƶ�+C�k���i��:-܉�wؠAeV�������14Ս���@؜Av���
���v��|����T���>b7&�9g}�mK�P���Vf{&.�bF�f���ˈ���ε�{M�.�`j�;��NV⫗:��t�w�f{u��x_W����.���+=#���'B�Ӆ}7}�Q{ b׫�5���n�쾒�>�1ڭ����~��Ǻ���=��q���g������;&5�+u{�l{j��K�UD�l�̍�������2E5�������N�,��	�*��ɏb^����k���'#w�����hv\��O���z`����+}�RZ�5��8�m�O'j��
�Lz�k�(�f�H[P2��rV��m��T孜نtS�ۑ~M_���h�&�pا��Cf��kp�d�ʥ�X�o6�p����}:��3=��7ˍT�ѵ����c7��>��Gf���Rl�$��g����sf���@&ͼ���&�s]�)�ջ�5�A17���h�P� N�*������4��~��SL���w< ��V{]<���#4�+jv�:�������3S���FLf
;OL*8=G�0l�4w��f�=�ӎg��_}����^�]\��§�\��(��7��#=\=U��|�)��^�Ԫ(;u3�l����{{$����r�79�S��cy�8�\,�|Ϳ _���#����u���-.�8�'�[V�O_�r�$j���K����O{�l��퐾S|��+Khq���Ëk:�6�w�����u���GS[���%�Ӛ�7x��÷cv�q�|<&���&��f6l��:u���{F�@�z�_��|�^h]Z�Z��hZ#՛%I3�k�y4�cZj���%�U%+�cw~p߮<�ۇI婽W�z�����i���u�y�rm�IJ��/U�RTV'퇡����D[Օ5�T�Yj�]��M�U�F��i���c"�n��ҩ:��Ix���Ʒ&,Ug��W��Ku�����#����������*���=2�k����a��wa����ճ�J��ڴ�w](�R����������⥭G��v4�k#�'Z(�<Y��R�
�W�(�ם)(ă�3fm�-z=����zT�0]*�tF���]S��Jd~#o҄��2��G%P�+�aN�8�NĞn+�����y���i��>[��6<��L�Ro�~�ד�J��64�n�f�Խ���D��B�|����@��-��G�Z5� �K��
�Հ=����>�~����ga�����q-�S3�h�Ő �J�o����-OZ�,��勊�ߕ�Tk�^LM}	�Ɓ�t)݈�yHYQ�U���H����=�-�����*���{]��o6��>�����˺r�Bz�b������U���:�$9YJ{VR��#��~���.�Ɵ�x��IG�x�?/=�����imL�K���+W��o$�h�^E�%{��#��fw�����=O/���ߊ�V(m�,_�"eη7�X���p��6��i�������󽆪yM��&m�v���ٴ=�gf��g&�kk�!����m���w���?w�}緓�}t�(��+�2?$�[t��߰��,V3XC�Apݭ��^��^%S5��	B�#r�a*�BRZ�jN����T��.Ĕ�y$u����T|�s���^0��(34�z�{�ʟ{�r�������E��־RPL��-�'0l��c"J$_%�7���W����z�j�am�@0���R^�J�T�P8ٗ���Ϟ���[+��H���s�]f�Y/��}��	�v<� ^���Q2�_ԥX߷Y��CO�F�(����׻ {����ye[w�P�X;�<_t��uA%U��m�鮎}����^͢�����5����P����~���9�P�N�F�J��:�;��f��䱊~�XiJݴ|�<������t�Cp\����L���Nnd�uoF�k�k����jۅ�~5�^IX&�(�g��(��Bkcۮ}bې��p٩Y�By����k�އ�wJ�߲i�W�d��CN=�f3�a�H�rT�X�z<]7���t�/�������]rX��0��fך���Z�2�@9PjG;�6�.{K����Ym�/�v��aOp��ͅ��.|�F1��v��뻠��#C�<u�\���c��d���f���*/&�y�#<��u��˖C�ܩvW�V�t�
��?�:��;S�� ov�!���kgsn��i�[�:���3C� O5�V���Nvtg�`^wm�NQ���ޢ=�f�tTf�E�*��x��a�_6oE���6��z�ݎ��8��\e�%�Z�f��ч��]?zT���YQ�n���dV����13���~?zg����(.酼�'��~����=�����K�r�R�/O�=G���WyIO���qzz�N/2sG<�C�����*�9�g�o����s��@�[9����|�0�;�,q=�gyzlL�{�o�1���MX}�=�*ǋ�T�	F�V�c^#��K|=�-ؠ�=��^R�����I��Jޘ��J�S��x�ʡ+��l/ݐ2�E8W���W��O��|��ޡ��O�@�r��§Z���um+��ݽ��h����JVW�S��A��8yoE�7M�a7�2��ѫ�ܳ��Ω�z8��'�P�k������e}:�u=�6=����r�1i$2�{+�/�h��2��}�0��`b{6O���jZVϱ�:=x<I�;o�͗}-p��}�s"�)N⥌�����jv*�G�g�j�kk!�秭�%�dt���J���������3F�=�<��m���+,��
�Xn��6b1AE��:�Zs'gw�*��d����y	�f���	r԰�3��� ��9tؘ�m����sO�˃������:�$Gc���=�e+�y6�"�б�"=���p�������������Q��t�mJ1ة���{����J=�x<���I�a��B�fF����)윥SN�mC�3��\W�s�׫,P���L��������ô�z&�vژ���x����֭N������i�՛�{R�W��o��{�-���A�SIˉ��[x;ԝ����.���9YJ{5k���w����w�P��4�Ǎ���ў�=d��Z]�s�/|�k�Xt�/V?[����^�������n:�g.���l��O�̠�+KOJ��f�a��<�|e�Vd�Ss���J��������r��ϼ����C���r�>��C�����H�x����VJ�����'|������k�*��㳀d^��s"��Xt+��V:����x߈x�Te�\]M��x��#s ���:0s�P�n�����XYG�-}�K�۱�Pq1�,<����W5瓸[��J�'��x?m���=-,ܕ�E�x���N��!��e�T[�=�ha����-H3��1��}��D]]{��j��;��/NƼ����n�<�\y���˅7���#fi%f��Sȹo�ɶ;Ip��z�B�B{�)Q������\<KRwƳN�&ruF���n�F��6B�T��7D�in	�?orU��{����`�X4��y�j��i��mZqݞj��o`C�kد��"pKX�m�`�}y�/��P^v[{��6�4u�np#:�*�Ӟ�4U>Lw�����.?U�ʞ��54�z�~B���횂��k�/G�*g\�g�^������Nژ�ЫV�����h�7L]����իÒ�=�r<��l��g��7-Z��.-x�UN�\�ם�R�֊nY��q8�_�ۓպh?c���2�A�s�ԇ/c\����=��$������e�gD�z$�f�U5(=�݋}-~���ڻ��wsf����{��=uf��%��w0�]qnμ����v!a��88��p.�Α;R/.�X{�F���.�m���[��&��r��.���]e� �쎴y{��8�3�ۻ���ݫT�M��F�W=�3D-�2_eu	�V�ԁ�%;Y[���n�::"R'n��|e5ʱ�@�h���w@�.�����m0s\U"�p��EM��A�hY�3��9X�1�N�7vN���OD]W���r��upXÕ��e�G��k(��߭b�{'QjTj�Ivu��{qU��ˣ�N���Io*�W�{�&=�a!�(9苢�I�{JpW�����7���َ��gs�Y�)a�Lv�Y������u%�D��il�[�x9F���s��)�B�����ԑ鄚��.����U�v��v��yHI�D�)��ƺM-*�Ⱥ����R�K��5�ϲ�ծ�i��skХ,�7[�{V�k�뛱]N���=��r`#j�sZE5��	3Ҟ�U�<۲��:�a�}��#']�qcwG^7�X���tR&:�����ly�������FICf����&�G��t[��7V���ݒ��뗻k���
������zPh��^j�q�ۗ+@���kWc�Iӫj�1r͖�i��tC��ቻ�z����L�_m#�fm�\W�1V���-5%�(P���fP�f6��)LOm��r�%q�xz�e��;���Z�F,�MOdSf̄�Nw�F��l+QT�Tv��0wU�L|�����,+o1�����[�R[�yi��[�RB�v>q8�]�w�u9˞j�4���jӶ�ozc�n�Vj�*
^S]��vK�YN��kOs��!8����M�/w��=�㉹ �q�>#�H_��!ef)�N��Q�Ck���ϟT���b�n^w;4F7�>e�o���zF��:, ��e���puwt VM�*b�G��N'-ܔڝ�%3�����*�G6㏣�Vɕn�W��3���Zo\�z{<b����N���s�IGS�t4;hU���t�﫳z��	q�mt�$eݔ�|�@�:	c��f6��hW��[�N�ݫ��5f��e���h:�GVYS�T��v�8��ye�Ľ�vj�w7h��"����8�eu�3qC�F�f�m�ǃb�c�p0t�u
�2@/� �~^���ӓqi==�z:�ўiLe��7�	�lXGP��,�ւ��a�JDe�Q�z�;ͭ/1�>��4��e�_�{�it�i�d��G3c�P�m�1�$w��Q[HD�D�N���V%8�n�m��t[�,盽�x��p�ft�'��.�(��wgI�9���g�-t���*]E���1=���2����1v�in;���킮ꦡ1���
��jB���c+�/f� �|Wl�2�4��&ϛ�)J�m-�=�]w��Q�����[���[��c�u�o[ֲ
���R�u�2)�>է��P����/�n<V��7�	��B,�sC�ߴ��U'YD
�+SD��Q�W4�.'H���I� �UEp��+�s�*���jR)�"���<�p��)�+Q5n�wC��;2�B9E
�*��*��:IRK.h�:�%T�)9�W* �*��$�"�Ԃu(�-.���N]5#�9��Uȕ�t�����s�'J�"4,���h�B(���X��j¥�����!�T+2�\�9Q)�9���\�"g#$�DJ
t%�NJ"V\L9F ����P\�U�Va���a�R�g9QȤ��Ή��,��UAT�*"�I#$�� �r(�I
""�QPA��d�TQb�wNX��%F��BF�Fg(���PGH�\*�ȹF�h*UUVb�QQS3L��Ȣ-hQȋ[H9UEUA���C�9R�Q�I6Qu�Tr�i$DPZ4��Qdf\�(�A�TTUeE�H�AkAR��<�:T?�{��c5� b@��� ��ڈ��i	d���_>���}kM_Iϭ
*�{{^��?��*����gؗ���x6��)���Q̿��;*��'��v��(#O֖���K���͝�V���kb*��\�}��VV�<Gg����~�n?5�y�&�\n�0����d��$��z�d�?�uE���zz����諼�5<����E��S��v�b�RMm�N�]��Y�D�{C�6��O�t��o��k�ۋh�ROr���Vw#��,.t��"�԰�l8x�l����������^�oy��l=��Ts�oJGu�%���q}G�����+�C2mIy�o�Rn��o�ӽ��o��zwLx��*�;�G�ל&�Z�����ך��{_��7-�*.|;�����C����qr�s������}d������ogI�}y�������-��!0 �r��빦׷|/�HT��,��Q���clzw�� �U��v��^={�J����כ�.�0���a<&bY�d n	�pTu���Y܄�!\csp��t�ս�����_i��+�QN�{���O��	�)���a�u���Xf��-��^��`hG,����	ݾY��M�	zd���� xV�}k)��8G��#3�F��J�zϷ�%���8�R�۪
1+�� �o���)��TǊ�k�!ld��K˕������L��bx��w�%���T7[�L���zh>��<e샕����H��^y�Ⱥ�z)��N^�f����ط�з땼��Ǻ`���a����7��W����YU�O�<��O�ˌ��d��j���	8'�j�?='(��`�2�{V>	����?zb�K��y�M�G��2>�o�yӚ;�ZZˋۇ����VE��C�z�x��-1^���r{���:��ɾ轵�Pg���P���-ίM��6�ua��X��}�5�?3���ӑݻ,G7����<�[^�;�����=7:�#�+���=�l��L�mI�؟��nnO\��U���΁�^��+%t�9B}Oi�Rݫ��f��g,�l��Sl�������e��;��`s����9U�m��ww���i��91vw����Բ��^�줵o{T=��8gz彧-CX?!���8o���\b�y�m�qbR���Rk�r�"]&�h���������x�����9}3��)j�7w��׮��i��^�x|B��t=7���	b����ڎÁ^Uu���񯔧�^Q�-����(����[�qM�p�q��� ,�#��mLvH�x�tv�{���l���~|�,NH��ˑׯ�e�ez�xy�}�FB_by(,��b�-"��VwWBbg�t�y��x�W��9�Z�ʇT�<�=C���C}���=r����s94�J^���&�4K^Ư�އa�
�f�|�4y5cQ�rav8˚�6Adlf���U�mN>^�R���s����S�����b�r�����=ܸ�;6�q\��I�'��<�P��>8�^Y�o��R�_/8sI��h������tIjQܑ�OI��}�E�g%��^e�՛�Ok+�^^[�~�CFTNBaa�~'�V�'Ow-״j�Ok�wΔ��]b�^�|��C��[�;r`�G��[Ƽ5��DE����(�x�ة��$"ӽ��E^{׮j�B��3�a��|��$ت��L͕�Kў�`N>1S����4koL�]]�|��p��/xO��Ww��0A�5�ڦ:����u���\�S�gh,@��]��o?�}�D|mֻpe�{uQ��eN�����l��u���-.�Ëk'�[Q��۸���4����=��9)@n�l'Y��_�϶�kӕa�ײ�� ����\o�w��X�f؍��!k�)s�����d<�&m��q�����W�Z�s��g����ۆ�F�kq~�Ϩ:������ē�&��������g�.�����;�ƥ�n�<�y���yRj������F�1���[U�(y�d��TD���/U�TV'퇡��A/{[J.���mm�V�X�YV���U��T��7D�U'S���m)z/31`��N^��3��wע�_��K����_j�1�Q#5���Tr�a�[^XV=�LK��t>�j���4ټ�>]��~���ީu)�/5r���y����<�������w��q�۱>N��.����c��\NY���\��Ǭ����S+f�k��y_v.+�Tsվ�ż�N��y�y]I2y/Z��Hn��O�v�53 �]�RVu(�ɜwn�n���ۘk�b�שF�|��Z���L�&�wK�%�28K�K���
"Y�4�8���`[Ш�������azrɏH;���)/.s��nhU�Y�އq�lc�T.#:+����soY�
�&Ӯ#��ƨ�-�W����=}+{�}}��z�5�{Ȇ�p�Ջ�s��>�0�f�y�}@{')ϣn�:�_U�ɮ����Fm��r����v�};�W�%����jg�5�&�f��|%��U�G$.~�.hyՑΟg+uSz�y�.{�v�WY*�d�t\G#�*���{��#5�c����`�~�~�nS�[^eyZG�+��=���\ޯf�]�O}{��Èz\uk՟E��zz�x��yHjyOfj�������x�Jȓ���Vt�FȎE���|#w������u{O�MP�Z�n���8Kʖ,;u�l�[ ⯤��Q�����d2232Uv=�D�����z+g��mtz�9F���;����߲�@��0���T���Y@�<���}eX�>U��T)�k��no���Zb@)��՛� �H:��f����Z�$cۺv���mz	�H�i{���3Q���Q���xC���q���0�?����֠�_!w��.1]^bs}3�{��O�.Gj�����f��=-y�~���*ۼ>	h}�������lce��<yKj�p�$���iJ~��Ƶ��;�rr�T_{x�b��l�F�;^��\���������
�~g*"]"I�3�h �5UkoX����з����������ck�s���T�����>�����g�إ������"7H��B{5�޸	�o�*���~�-�/�t�cG�̅t����hˆ��7,��ju�& ]�ڋ���ݎ�o��>�{��I*�5��4�bj�g�K�%*�O��XȨ�ݮ}[�m:g�͘}�ԥj��Sza������6���=6�3�z�pE��sG6��.�&�a��/-ȣ/�V�<d�>~�.��,�����f@�ܛ�E����ʝ�^�;�/|�x�N�K�[��*v���Cy㧰�%��g!^fM�{�1�u�:���5p3�1o	 �<��ֳd�bg�7��Kr���@<6 ���gZ�x�Ү�R��j�ݝ4)��{r@o��n�]�T���0��͉'�mkH9c��j���ˎ��j;�j�^4pc�xk��Fd��Œo-�Y�h����#Q�u���}�V�ׇ�E\�^Us�cj�N��������]s{�eq>�ٳ����r�U�Pg���5n�bڬ���]Sn�.�=[I�Xz��\��4��:t�{bf��􇝋bN�� ���'���``T�7pa�G)��##S�r�Ƕ'|�r�x�k�*��X\���cՔn��+������k�T�Jd����c����\7~{^�y��qa_ֹ������ejS�7xp}�n�Rw]�^4�?\4���XR$h��&4U�[6�أx�Q��p�#� ����k�#��kܗ����~�P�z�s�f�'ޚan:F���_j���b{6o�] ��2��:��5�r����[G�.����͜q,.��6l�F#�bDv;A�ec�N�MKQ�|�Rj�*�zՆ�;��l�Kv�D,֐��U��v}�͢r4d�s4��!��cQ�
�-Y�bNY�Z�W���C�%��̊��)Y��q
�/��i���4����O��^K�C�V�\��F�t��1gl��+w����ػe��a�l\Y8gs�Űk��u�ƭZ��G�����w[2��o9\}�������R�2�-�*���5��b&*3�wӸ5=1OZ8$H�r��}��ӺT��O61׹E;���NΒ�׻������;oy��Y�nr�|p���=���x{]V�q���c����c�tǼͩ���x����N�Q���	��bZƼ���	�'N�N�C<�6���;��y�ϭp����?yTD���xzhFmJ�.z�W3ꇚ�"���O잢;��W{\5O�my���ih�~��(��@��n�����]^��R��-z�ys����7{ <�[SGt��L�/E
ʺؤ����V9�dF���ہ��Z���j�kۂ�}7;ja-Ƽ����/�k=��Β�˶
ޑ	��8oO�#�cs�[�x[�)�̕k<�]7Mx߼�=������].�Pt/ӵ��>ޟ>AV��Ԑ�ܸ�_{�G���6�3�K�/:����S��E���K׌:�w���#Sr ��:����+���4�����,�OyY��%����G#�����׷@�]N��lQ[U���������m�yb�މ+�����������z�����&�~�;�=���b���ހ
�//�ۂw��S;��5���)�Q{x׳h�)��o�=�~g�.���l:���1�%(�{YU����5�zv�V�ǵ���p�l�y��V�ʗL�!V��ՐR~RӬX���_k���Q:���o�*�SI��ý	+�]��ؖ��0gIyܟ�u����;���w}��������Ὥ6���lc���&�Iǭ�ۙ^�����U�U#ZB�xG5���K�~=:`��v�4�[��ڰ�'�ot�X�W���o�;�M�g�Y��^��rJ��߮��z��v����~y��-�Ӷ�qr�S��]7�K���I_�S�WsI�R��u�*ej��L�iw���{������/֕��jz�:���~q���UI9���Ej>�Z�<~�Vgy��g�~F}�PPyP��{��/�N$��zB+�v�H'���7m�U�)�X8�=4�[���o�h�������W
Z
%gt��*�ߵ�k�I��y�6𝜇MS�|��XH7֞��_g�r�D$k�s��w�"�̺u���S�V���3r���'�9�ҟ���r�q��oKw'�u@똨�;>7�o��׬WC����	Н��-�Q���'�5Uf:�Kz�/f�Gۣ��ז�]^��^�K�N~��;�w�+oY��o/M�(��v-��v�9���>��V(T^��i�Kpz���m=�]�k�ͥ��w�Ы���'�Yw^���sӵ��לn��������^��p�<M?iV����r.+.��V���B=��m5�k7� ���]���F�k�Y�ޫ���E�7{P�ʪ�u��οU0�#�G�wlP=���ΐ��z5�G{���R��Z�}�M�
AޱY�lJ��`����{���d����&����Ib�)Q3;n(��{7�X���\J�=#`�ψ�y�LsH�{"w�C.�K5a�zxx��~]��.#sW�
��S5�-�Sg�k={�RX�f?[��ò��ʬE}Ԃ�U�:�d�W`@&�l����j�4�ӷ�=z�������wq�Il�'l���n��E��q��jX�a��Z�l�iZ�-���8�:*�~��I�:��	Eb����t_+�i!���觲�0A.y˹ry��2-n�uV=�n0q^�4N�/C���nL�ٓT����<�3�2�,]��Aέ�Q����8��l��kDhcW*�@��W�EW-'k�Mw͌Ќ�.���1����!A�7N빹W/h�g^��yȬ1ķ0G��,&Y�Jw��e�<���p=�c���J-0o7z޹�w9v����"0��4d*�Y�
%�&� z����� ���@=�gM���b\t�}z�]�^��B^W_L�:�fо'���ysUՎV��w�L�v��1u��(�@w{N\���_wA�4s%��NeJ��%c-��\z8�H�6M���o�ۊ��gE�ߖ�O�Q�p��y��u�.�y�yX�s:D �&��c6&ҩQ7x��W	���y���䰭)���6#f�A[�.��n�&Ѹ��MͫsG]I��F-�g"O\z��s�*�5)��M�.n�
]ws���F�]+3Y@�mK9��N6���}G�iUгt�u�YM��^Zq�ۜM'��$����Gp1{s��mn���̮� "�e�����y�R�-e΂����G�{gD���_Vy�x���u�os�Ǟ�܌�aV�����<�;�{,kZ2�hM��,|5��-Ӏ�oK�Vt��'�4�ӝ+oV�y�����a���1r)��o�{������3v���LƳx����y�硯���L���7�a��S`�j}y����'��W*���,��ag
�"��h>��;)��t6��h�{���ӆ�����4Q������ѯԭ�x�ou]�R.�� �U��o��Y(p�m>�7+W&c<����::
�J�ko�8ܽ�eIU��'r�8�j���\�E���Y�9�qA��ɪ�g�l�DA�q��)�r�qTF�;�M:[��)�3J�Zp��5`��J�;��n;�6�M��]W�XZ�^�3sk,�l���<3X�F�^�~~����C�u��G�e��E�X�{tmBal�vXU�+!w��$09E��|�daU�J����Ι9O�24�d�ԁ��e|��>{���-s�}��0J\��8�
��͚Ɏ�^�t��;@lu�W��:�_M������M]�ٸ�B��l+�X2�кG[|)+���HS]��=�G�E��ɉ���j�����g-��������T��
���ۍ|9�����W*��ӫ�w,=]t�|e-\��ǩS�q�t��ӈ��ڶ��ܩ�E�j`չ�G���0�3+hY�O{;eǽ���Kݣ'W8c��p����g.�ݝz����X.�'�}���B�����|�9ȧ�+�Hʪ"��Aʊ
L��b!PFt�H�*����M2DBga+,9rM0�R��jAUU�kL�E�D�2�ʲˉh����4D���iuB�5�TD�AȲ�E(�E�Qm�,$T��t�J����Z���7J�3,�DF�
�%B#����t."���� ��D�9EG(�".�.r��B%��L�9ER� ��s$:dQR�����UU܌$��EF�U�
���Z�L�Nb$������VJl����e�%K�S.Q�*��G'A$Ȫ��bI�B�	�"$®Qr(̹QȽ�QG*�9Q���G!K*.ES,6AQʂ��.vZ� ��i�p�(���s�Pe�E
!s�,����U��'� �
"�\եu����YM�q�0������ݶ�޴*PZ6F3	��>tO%m�
�ј�(�B2�^`W�voE��|��[�]4�7�ק'�^ʑ��Ķ�>2-��Z�2��^׀^Zt�����_���9�E�ċ�nM:�r�u��
�qr��c���!�o;1�za��t�Ylr+���u������<��Éw.2�q�1[~Wl$3��=8yQ�9;5������g+Z�ڱ�9Y����N��_�c�vbc���^Jg�ؘ��F���b���qʿ.߰�ܞ��k�>������B[�*�*7goQ���ѷ�c��ОS�H|l�8�7��b�ίNs"^��pa��T��Y;��~�ӡ��ɟyvן1��hqϬ>�u��^���FK�E��7�=�ɸ�Ϟ��{�ղ}�Н'n`��Q$,�1��{{Ե���ОϢ7]	��y�}t�����Q��f '
�� ��V��Z���@Ɉ9-D%�;���R����\yי�7�s�EX*z��ut
��Z{o�����Q�߁��9stjʦDV/��C�Rw)V󥸖�M��gv�o�[���Շ�|�MI���[�w����-s3�r������SֺsA>�S%iw��C�|��F�_Qd�������ٮy|��rw�ب:_j�*�+�8٥+v�/.��d�ѷ�ǟ�
�_���o����=��`�s����(A�\��؇ f��mS�Jj��$ǬbleC�sC��f_O�����ťѬ��qn�O.C���T�:KZ��އ�LT&퍡��_Op�<�t��uٺ׹9X���aMtH����=#{eN�2�b��Y�{�j��FRYR������G&2���-�|�Ѹ��5*5���ς��P��k�m�;���x�f��@�{�j���%����啫OI�L��f5aԅY�������E�z�rڜ���ϱ����LS��u����	T_�H:�ٲ���ۋ�E��/w�y솿�5�_�k�ZZ?L�K�.~uQR�������t�u�n؁7��tk<�ۮp����zC|�-�q�;��1?m?[�ɓj��]�w	f�����l����oz˫x<�W����e۞��.��F�5~��e����F�_�Hߜm\��g�*��:	G��LNk�@<��ywS��S������>��ŵ,Y�wr�)C�!N��z)oRq����G=��ŉ>���bɵ�Rm���[��k���^�����>bb�cO��K
�D{0�G�̘�َ��p���6�[����u�bv��12<�����N��%���;=�����zGdwnw��wl���M�o�U��O.ޫ�6-QϽ�)揷�ϐ}����܃��g5-���ۡ,���oV\m�a�K��:%�_���C���({vQ�'S�`瓊oƣeo��X��m?3�I\C6<�﷑�>�W���W�έI�pQ^V�H0j���y���p��5y��Y�ͿrԮ��qoe\�u�{�8����"�Ԧ���������M+e�p��Ā�r�F]TR��j��8G�����@ǎjVzj<��hU�Y��z�X�+ �U>�	Sy݇�NgS3��ԍE샓�ͬ�,�\��o˳��Q�~�9pV"KwD��J�zjy�
ay+�r�T�b������>|��*�Z���W2u�˽���P� 1�Bܛ+I�d�K�!{�����gxɛ��bcxʥ�gn3�*t��Y���OiznRcq�-u���Y��z߄�ܽJ���-�&�q�^z=�t�����t��������AV�n/��6�޿eM^s���v¼��zl�U��N�T.����+���}�p��Y'٫O3���S�<�CW��O���[u("؝�9�.����u�����Vbꕫ������?��H��摘j⥸6��M������9��ե�r��Ëk;�7�]Qt�'�������s��O�����Cۘ��;]����b7�5n�A���תR��|�'SO@�iM��I/��j�W�2����,;u�h[
��(v�Z�MN��v�{=�Ƕ%x$�4���yjoj*�l��7Q�����-j�y�Ik7����q��R�,o�C^����iޅ��Vz{I�!C3�N�.�l���;��{\��q�K=���>��~M��Uσr�P�PQs*H�J��̴*C6ϸ�QR�"ά\U=��y�Bb����7��Gdc��n����B�1L�߭�-���'qi*�d��B[�����cyQeG�(��cl[�U��(���Y��}�;��j�)|'�c�%Rc�1G� <��������sy���g�X}�ױ��=Z�H�������(g��N#�X�ʅ�%7�\�gA���`�z�P=�6������1���KG�g9���/Ww���ߧ�ď8��N��F/{���<��)&Ѵz��/X1�/=\����/ĺe�*�et����L��*v^h���ǗzԢ�yŔ�_mT�j�s1-���P���y�5��/mM<q ��c���Rj{��LG�|�ir�����J��É�6N��zlOwmZlgG�Vff(���޷=��߳����|]V�<d��c%ܸ���ɚ�kNACI�;9�>������鶗mVM��V�w�V�"g+s�����>�ų����x��V��5��A_d����Wd���+;ë��q���mC�;�׳��WyHjyM�2�5��߇���{���";�+o�]{T{򗶼�xogj/���T�ES=�]��ƙHՇn�.�K������e��������%Ñ綽M�����7K��
�m]�l�ގ�m+�"�V^t��jk	� ���{;b�`!�����ˏ+�t3��z����ڷ����%��6A�7^�{{7å�7\�mg4wg�q�����5�u9���Onz�߭gm o��&�G>{Aμ=;�����N��jJ�i�����8|��yc�\������p1�x��m<Ŕ!Ag�P'hjW�klק���AUIJ�N�KƾR���XW����b˜��g�)�X�м�yV�n����=/��/����!���{�]B�ۦ��Ol�-�������+;`����.�IR��;�Kl�
=�ߟJ�Νޮ�w_���3�	��uNB!i4F�k�3d&��3�	a5.'5��n�o�*����v�����,��;����Z9w�G�X����sg�ͥގ_Nx:�s.�l[�r�1ibs��cǫ��[y~�:��KH�-��H�Y�X����jwi^p����hj�޹X�^�6�MF"�PUh�ͻjhw��)�T����veI���7.ʧ.�o�����}-�xͮW/4�Z먴�gd]��
�dX�Yl�����!��}�T�+��E���,5�]��7�G�T���x-s����o�����>�le{�j��գ�Y�/&�f�=�'���xϓa�T7�R�/��s���CCƫ<5U	�b������-$�>�kt��b�*|�+�8�~*s���u���p������BQ���q%s�Sm^�99�l܎�#�}��]�.v�^W���̠�ܭ.�Ǩ��ěk�-��)�k��E�s�؏m��Z��O��̦�n���{��ȉ�3������fz���W �,�B�����Ϣ)��ޡ����ޞ�-}]#�^�C6w1�1l���$�*5d,���ܩt�����IF��I-�Z��on'���X����������Oz��o���X05z|B���<��nކ���o{):n��Y��� � ���Q���;�0x��(������l�8t/����M���W>�=��x;���6o&c��.�T��s�dR�����h�*��n�>��ۻLS�H��r
+<�^ n�]G��<Gx�����;%)պ�QNˮՖ�k�d̛�ېJk����K���l�|LVn˚4�Nȫ���϶�Ջ����}��aص��4=I�M�����\5�=��ў�p�l�z����ed���K^��N�b�ֳ�i������"@��ul����L���4��qV�I��lx&���Pߨvp�~����k;.&����ӽ�9L[�B����t��SMڎ��K�����������K��o��Y���}
�"��p]EqC�t�淝*]�1<��^�!��5��>����X�b���_s՗��W���{oޚ��5�yt2�A�n}P�x�1���C�ϣ��l�1������2a͏v^y8�O%�ߜ�7VUz3�/ٹ���ڬ��j���{���T�n(�x�R�.5<v�^�c�(�Yje��ˇ
���qʫ��Xqmgz��ꋥ�뇸g����<�J�uc�����[�!�Mſ9Ua��d�ίM����R���<j-A��
����%�ag��.�ɮ��w�����x4p��%Z�B�Tt䰹�����P��ࠕ�y��޽��{��ϋ�4���.F!�ι�vpBW1�o��f��{�ېEN�3�{�w�����m�F�M�#2�{��r�����*��U��IO�v��u��y<^;��l�V�����.2<ݭ>��חR�Kt"۹;#"�YX�b�������t�Z����u��`uЪ��βTy�'=/w�X9�D�j�J+�����ypU�x|<G>���H���m=��V�� �H�ןR^4�?\5�k�y��|w�!�*���M��x��X�Q��{\,�����|��1�vt���ο�}{Fle��S;������H�<���r;Ϡ�}՟_/usu��
�]�YBq�"r�e<W���Y�9�C���=����{�79�� ��o��-�x|�v�u�z'���4����nآ����˩�og,�A�������a�U'q��.w�T��f%�1��B���c��z�O^7�o���N��}Ȫ��/���W�\�l8�l,֪�O\���kY��ĠZ*C�D��
��J��7�Ҟ����9�oȦ�s���<��<��g���}q<�Ӧ6��͓�<�+)�/2ۇ1�3s�Δ7-�W�BlK�ۅ
�)�
<f�u�fn:]X�W��U�!/
/��9��mL��h.�C�yi�g8�����X��}��4gu��Я~G/o-�$�3K�^��&�`w��'4������L}�#_�����ۇ�r�{ҵk���U�y�&v���5��y	�v�\���[^�A�Ҿ�W�ۇ��=�8ni��^܏6�l��u�:�Կ=�jI�'�A�V���?5���������z$���gW�jתm���==Dt�aS�_��T<Xvhn��+�_��?*�G��'��'�>߰z	^��g��]Y{{�{g��d�n�Zq�{s[}j:�-�ݥ�t�=�
ސ!n���OGp��^�@</(oYQI�v^Ȥ����8���-���~�w�
����v��w��)ڽn��x,�mwf�͢j���"���ܷC��ޏ,�V_���r���L��}ֽ�����\B��������>���-��؄y�WԳ0J#��L�i�?��'v^ɇO�n08�kE�lT+�{��w�����=���h���+N\{�j��p�}I0篔�v&�~�`��GW��d��ծ�:���i�,ݻ��6ŌK䕾q��)C��]֥n�w����λ:\n�r�̙�����|�m��"��oE@wMEf�`9�\��i*�(>G�DK%c}z��v8D>ѡ�;v�Ws��F3٣;,�1��CU�q�GH�-�\�;32ܡ}WٍSnވ�]��Q>/x=�}fm��=�=���ͤ�,�rru�{ͷB>�i���ˡ��]�e(��9�Gv��ٛ |/�v�"�A��ڸ\�����j�VXOZ�W{����j�=R6�~��n��7����̡(CԷJ	BU�Luɲ:.�4��]@�[i��ٙ|�K��'L#�icG���xP��u+2��
��C����@&U���]�.���� ۴���ޫ���fiw�-.l��bw]�O��aw|&�0_k���%��D��q�-�4�ź��.�T2m��b$�38�ʽ��H�����b���b��)k��Nq��8���-Ľ^E8]��b4h��O�$Uv���;�:�T���m�cN�̹gU�ߺ�wN;����bok��c�}���Ѳ/~G��N}6��j�05
%�W["�)����`͓�2B�j�U��+�]]������x6��e����ME	`�i�	Ǝ�r��7`�B`��w��v3ki<ɖ�����7T�[��8��َ��7
.7�e�'b�eh��n)Ƣ�=8f�}n]bA	���m���S���,[�4d�o���HAk�V��	�h�n�fT��r�D:�2K7��;}�4��{2C5�{9λc���u�r��	L�K&��M����ѧ��O�;�r��{��z�L��ۼ����3�A�5l�0�q\�����יK+v��ұz5�-��r�p(ӽ�Y�a��6�yu�0�Z�����{�SN��;�@��+�vL{����;�+���!̙���j���) �9$09Wu7j7+H��"����t��g ~}v��}�=9z����Y�ٹ�{����>��f5��!���eJ��u��\�vI��u`]�>��[ԅn����y[Wʯi(�LX�e��O&@A�%�K9Dtg�������6����2�@�g���T�[*�3R����t����+z�����:Z+�����M�;,�����F{�-$o)m4��v�"��܇
W �{f u"n������J���|C���#��bU��x:�t���u��g�Tdᮖ�N�򫭗��d<��� X(����/x��Or�=�<�J�'.�#o{�k��n8$�Pm�=�(��"{Svci�w�����M�ĥ]���\Y^a۶0%�!{���ݻ^(�1��������}�_F���=��1�_f 5���_2.
G�R#�K.Q�y�w- �����ep4���"R�rr(��Gݣ�UQR���s����tN]�lS,S0���9�	�Dh'8Ar4Ģ��\�	�H�iIG4"��Q�G��T
�$ˑEZ�QY% ��
��G�"�9G�<��'�"�,�I�Tu"��%B�� Y�I4�Q<D��]n�D�U2���〳Թ�ª��VTT�r��",5�UQ̢tM�u'�φ�U���r�D��힚���ݖ���J���K��9JQ�%r"�CX����4�("�1�*�ǊU'���� ��L�³��G��Gt��P�=���Ur�̣�Q=�S����yx��:I�ɑ�n.�^��t�U�C.���)X��$�9��IQHT\�WE2e2�=�'"�X�y�\���EJo~={�� �����EX��E��r��(X��k���6E�Fm�/�+E��2.�|ͧm���w5�rJ疖��o|�OZ�[{���^�4ZJ�%�g<)62�S�*B���uЊ,�T��'��nu/�����o��}�T%�\�8t�hj�r�n��ZbqD�	�����J�T���tn(��W�K_-VC�����'���wp���c+>��ɜ�gG���XG�c��6���ۘ�����/�VL?[�|=�n�J�{�+�}�^73��v�4�G���2�W:�̨����;���t^ӡ��>�ɚmA����5����{n�gF�UX{��:M�]p���ΎL���(���Q���p�z��T���k���j�G<&�G�#W���/�5���>�ڮ�������_�0����ø�;#���ۍ?�R���U�oDT�.+g�Ų�ؼ���\��
%��>�������eΝ�
���뇒�RW��)t��<��7�9���|��\�]�u\�^G]xn�V�wf��+�c����~�u�Onx�,����g�v��uR7�9���C���@:���ߓW^�|_�=R��Q�-��@C�r�9w�e��'5�K����1�^��SF�b�C�����ՐBv7|"��:��x9s*�]����m��a'���%\��+�x__'�i5�J5��Ϙ!�b����c�nO�ۻ].���S�R�����=����|o�n���K��q���*(���h�UA�r���{2öoч��M��u4D�$�;g�T�^z#:��G[����4ωwP$���~�ʡ��2���)E�u���fnFz��Ր3��E��;���O���x�ǹ\=��q�F��Y�������{^O{��{I�����xb��W9���\:v�7�mD��θ����f���<T�[5,^lw|3���q�p�|d���q�jk�Q]z8{�vǾ�Ͷ7;�i7�:Vμp�����C��}��E螉SE�D����[F����R��_��=�ԉ�Lg�7G����T�o��d�2|v�'��t���� ׵�n(�9W���&�jq��*|j�-��גz1m0_�W 7��x
��_q.��b���7f�{8+>�|r���#�a�7�TL�w}�gR����ˍ�B�w&��&���{�3T=�O��6:T���p6|9I=S�/<��~���*g�U¯악m]Gj�0��WI�����t2�3f�O�f�X���7³�bt�b啯@��+��͵�����Ǚ��N8�T�o�G2X���">�d{q�H_�V�p@�{{[����2��yp���/�yGG8v�{ۼŽk¾W�踨@<� �N�b<��<��;;e�:�9Bw�~�f��97�KB|=Z6�^]8N^JW�~y*��z1���v�q�ﳮ(Txl���m�����}��pf�9�׫��S�-m�Gל����]x�:����̙//��-��e�o����vߪG����(��}�	��T%?����d�ƨ��/��s�>��;�qj����3��g��R�.�B���^���\��;P��Q�.#f�^����>����l﷽|�(��9>�ǫ";����j�w�����d��RIU2¡3��E����Ov`�ݮ�屮�����#�^���ި(�������G[����7�9Xe�DZ�
�p���FnkFVVg�=���|�b⧩���}惛�{��܇S��<v�|�;C����<{��G�,��+g��(�㧙D��3�L�"������m��/��y�s+9Qªb�|��}��ImF�מW="h�B�WE�e�[��l	�� 4�*�L=5��q.Z�Lo>��QS�����P��>��Hi7�gT����؞�ӱ�9�uG�r/� �V1}�'���쌣;�;Z�7(��r�I���>nA�wi�;SWJ*#��E�ܺ�˶�f�W�m�9�Ċ�^8of��ӤD�2��r��Uϳ��!�y�>������X�Y�7
ԵI��v�[�u���u,.��Ny���Ph�#�$��u䗔n��K=��w��>���=�:v�}נ\GU_����©-M��}HWwK*�{B�T{�޵��;��=�٥�S+4Lv�j�M���<G�y3^�o��J$��;f��7<$Nv_��Nj;�F��^5�d�ޒ{U&&����3�3Q诹Q� ��/�����j>���y���侈0���T����]=��%��[w�Ʈ����O>�w�>T��U2cy,5ɛ�y]ǛP8�V@ɇ�'0Þ��Ϩ���o���eZ����pP%{�b�Xw��j�3=�Vl�23c���=�'+�|9�0�累��'�gk�$Q��v=�J�!��Ƿ�tN�,'��\7��Up؟蝟�~Z�5]���y�ߍj�c�4��=fWQW�=��G<%���zDn%qř\@Q���}���i����2Z�����e��I��s^q�KVoY~�9E�!)���W��p).��r����7��x�\v��D]TqB��L��];��-K�Vt��K��H�S�ʿ�M^� X�W
P����;k������^���Xjk��\u�J]p}ؾ���g�d��B�.K�mn=2��0��R������Q7ς�h��̀�K���P�:T�sE�}��7��%����5V�Jy٥"S��7/2>�����3X뗩�ZP�\��h���'�B�Oz�#�*��4j�b�e#UO�Ԇ��������e���z�g�rU��2����y<]��MPrI�P4_t�^�����[yq/jV��`hu�&m䕍�3�Inw:@�+ܨ��������'�L-&r�~��@����n����r<�}\��n;H����;��W�r2zi���x�8!Q2��0�q�\�4Z�����Ƽ'�p>͞��֎�:�lǺsm��3�M�냷�wƁs%���@��|zo�j^���<D�@�=74=];�<P�l�pھzr��q�%��5�/�D�YL�"z�추dQ�D�ӳY&�̐����qZɫ�2X��j���܄��=[ �v�4��}�Mh��&=p9�t������ED���慨9W�-�koΫ���3iڕ��'�m�
�_��2/#�ˁ_s�Lʸ��pr|�uf������0�[]�������}ñ������XTc���T��롷ΎL�����G��F�����[�;1������(rI]�{C�T��m(:���l�~�r&�R��	jzԗ*F�|�2��X��G�Fs:�G�$�hY�H
�h���p;�}��w��-���n�յʴ[-T��"ܺ8�,�{it1���(��t��ќ���1}�D���ρ\/���s��`�ƾ���~��5�c�7�[�ݵ\)~�Y���3��3���_*�j�z�ǣǫj��j���`��'�pe9D学E�/GDK�ހ_W���C7�c��1�S����<�����^�Cv�������	h�>3�>� r��S�c�+�\��K�Cgƹz{c�W�;p_XVy�����J[a���v��WU#t��U��c���%t�5��RT/l�E�����hp^���C��HJ.Q%��L9��.eG�e�]�:�X�V��.޿g��w��:G�g\>S�\7��h?F��.�r�%T΁#�C�Lͽ���*կ�~/k�ʘ���E��j+����/O�;d�ۏr�{�=^�ލ3��n	�yp
<g��l�n���s���L]L���n�M�v�7�m���+���g��
���Q�x��i"��[�~^�y���p@J�2�́PvW)�@,o�V�
:���Ͷ7�w	��P�5ћ��Y�}���y�l�V^\IfJ9��ʠH$���t^��@�j�o�b�>v����n�^���d�QW�p���ӓU��WW����A��*�z0�J��6�q��f0�����ᢡ[��+������I
x��Sƃp��Ǽ;����ցщĉ�[Z�7��R������ս�:��Pbk�в��J|)wY컮����#+qI��u.�}�I}������Հ\D���%���|��� ׵�n(�9WP��l�[��w�M�u^�{i�ﻺ�=����|�x�%���Z�<��;6+�{X)��Q'����P��+Ŏ��!����S����|M��P�f�z��G�u�����
�G��n�ml�v�z�͏fj�v�8�	Y(V�����o�ں�Lc螒�'��uH�}ʎ�d.�A���g*�e�-$9�l��X6�^Np���P�˿=	Wo�������k�.�[k��d�9�����|���qD���9��z�MӜ-m�E�+��u׀��;}[�{���j�+-��흒��������.!8�7p��.��]t�v�φ��� �,ѽ̐��HbG�{������H���ᜧ>��H/.�B��u�W�l�)/Yek��O�|_]�ũ�~�um�dNs���; 6G��1P�R�Ց޸|_R����A�9�P�I+fXQ�>��&�O{�O�^�z{��s�9��<Z��P*Qe���|W���v�ב�W�����}��ƽ׭MƁb�3�̣�wwB!V��ّa�����A���>�J����l�.�1�B�	dD_sOk�c�n�	Q�VȚI�Ӻ�]�FneGĹ�=�ˤXHjԊt��X��afA:���$"5!}tyX!T��{2�Qn�ar��bه�*^�Ti����q�`��J�2�y9�������`�!��{��|�;M����.v������5�:|at#�Q�Q'��:��"�KfIAv�~�!�����̬��|�!sң�)���yŜ��'
��Z}G�� 'Pf6���qU�ʉb��U��LďA���޾[#}���������o��F�u�}�G��9 aߋu����N���Ʀ=gs)!������T;��m�'�{����m�^�}U|j��Ū���ā�	� f㝌�޻ȣ>�O�
�����jh�w�6�����O���P�x
�����2�n޿EN�(ԡy���zx�]�b�ru�S���%���!��Ra���4{�@�bb�v��m�iΙ�"����)D�7.r�@}^1���������䱕n��F���p�uJν���!3g��k��sZˉ��|2�Tl�]' =��A��9��)��ll��Ee]0�P� �U(�nt,J��e7!�*�Vϣ�hm�����<O���neC�����xO�����)=�~Y�6�oLP7u�N� Z"���.h���k��Z�p=�ݻ��ӠF�Q�)L�Z[;%�ݝ���n����Ʈ#Q�Z�)�ʲw=N�u08[אoR���
@��l���E�����,�s�V&�h���\Ռ%Z�r�j]e��QZ���רV��U�S=T�Bu�x��X���.;�Y'=�_�/ƏNT�GJ{L䙜��l�u��ڏQ�%�9=�5qމsK�u՜V|�.Sz_�zg��p��LC��۫�7\���cΐ��2�I�83���a��w�K�q��t�N����^F��F{U˗e�G+�k�Ǣω| �cb�y�!�dr�� �X�_
�>��Wh꜇��f�ǐj��y�����Ŧ��I@�iPeSJG>����:�Ì�mv��}�w��� w�WF�!��c����A�NQf�Iuc`LU⌶n�P\|��>��鋨�SW�T��^ͮ�S��zI�;������De�u��i�� ';'@��	����Tx�h����wZ��z��f�+S��t�"���wI»:�{b��������p��]�o؅C8L���۝j8�z�W�
NP�@/MDymhnz�0�sm��3�K�9�w|h)��Rԟ�������-c+��GT���@����9�9�x*Y�C���cǹY��=>�^nCu]�SvF�,"��嫹��ʚ�=ǵ,sLn�����,V&�]u�!��L%W�9J�T�b`#Z���ZPh#d�DU@[��������wc�kz��H�ۜ�c;HFU��)�:�X�4�e�te�vM擛�c����Po�d�F�Tn������eĖe��2G+�;f*^�Q����W,uB�d1i��u"�M����^��3��@��/�d�1{�7��z�W��}&��ۘ�����~c��$��1w�<Q�~���u�������ݝ@u_ϯ�����\
��zfU�6����;��¾^�Owy�^�'�R�X�?TƖQ�]�&}���v]p����Co�����Q�����o�p]�7<�E�׷�~Y���}��.*w	�q��Qy{p�*k�ǡ���=�<+W����?��>!Fs��;���Ú�!L�fun�Hr.WD�C']O���,�dB�`U�/G�u�Q�����jwN�)2>���37���_�F?}��s����	�:��,(�Ma�� r����X�%|��~���{�W����m��\��/���9�+���甅���G�|JWa�����H�S���C�X}3�����ϣ[c�Cݦ��E�1���hp^��C��HJ.Q%>2���n������'=9}�ב�ȿL��5�x�Ǽ�)�s��Z�gĻr�'�%�w�w�~��ـ�ly+��{�!�囇}Dz�����n�W.���Z�h3���W)�C������ܼ^�K�[�C�'f�c�2�`�<��BU�b����m�=w:G1���ay��W��ޘ�hhvM����]L4����MB�A�v�WA�ӷƳ�T��A�]��1}��0��Z�i�:��
}bf8-u�f�,�eܳ|��[��TT�E����_C�ü3t���J�@;x�bV�F����IfoԵ�!k$�|6�.��j��>��e_Jj�]��s��{ۊ�dH�]_�d�;*�L{Kk���XH<r0�մ���_��d�v�+c�VfYl�����D�T�d�=��*���x�4�e^MYo��y{q;��Z��m+������.��O/��Q��9��1>�D�Qw
	�٪���7�<�>).ΓE���\���Y6��}K)
�yϰ�3�Պӕ���$;HκOR��lh��|ok�I�Z�mkވ!��:c�9����^�=D�;�h��+oT��6�㶥�L�dt�1�N���,f��77�`�C2;[�4����� tw��a�m¶�b���\=�i�i\;�))m؁�K��h�R;��;$|4s�CSOs4�/pw�8���v�[�x����$�5>�4g�f��B����H��wj���N�<���{��\�Gܴ��S��*`��9!o7���i�!j6�P�&���V����3u}�»��^sk���8z��]f��z�8�+8��4�@]Nz_q�JM�,eز���I[$�S�ZY[�H4�s}�{��pF��]^B��2�.$8���=���vޮbz��Z&m�O�Eg��VnP�}˻�e|G�zd�m�Sϼ��^��>Y{�������H��+;j��=��[�79TV���qM�+j[5W-8�o'��+'yɍ�Ym�o؋�!,gk	��]�=��(WS�"K�v���⾸R��m^�L��sA7g5Um,Q{7�H!ׂ���aι���GU�/\�����X��b���{g2X�će7j����c���7EN\���v1+�T�H�C��uέCdVلWU�Ǽ	�̼|Y+nK�܍�Y�	Nl�W�\�ѤwS�����Ǳ�v�H���q[�I]JQ��\�T.�,���I����2�G`�#����Ö��v����qK�	`]��2�*����UrZE;t���u�#E�B�_����'=�=��jxם���u^����3m�N���u���Wу�mw�)�r�@��ۡG��%�H���o'�Aw�pڰ6�b�_���y��<��X�W9��Kj�7���9SU&9Yef�X�W�z��=�}1n��S
�j.{Yen`�$������,�X���.V��]�Ȓ�3��꽍,��s��QF����˸"b�F���鯨v�co-1ǡ��E���G����Ϯ�_��PQ[�uh��s�A���aQEI,�t�bG�W#�M�A��*���%J�w/+�i����P3Mͺ$ENKL��EȊ��j�t���3eu&�ZGn�NTT�rD�#�W��Tss(��-#��(�G��jR��ʊ9\�Fj��dus�t�w���ݹ�䉮h{/Gq�*�BL�"NZ&Ug��:U9��VaW*�j�N��(�T�p�;�Zby��E$;�^�RHBt��e^��9R�q�v�p�B��.�9�C�ETr
8\u/t\�S�����T�](��Y�3�
��.r)2HJ�G	*�6Er������=�
;�:���2���*Ԣ�e�&��W�Ěp��J�D�#Wf�ך�������ܫ�a���|���D�5L�w��
�#�en��G�3�t��ZG�2�-x�%�n�%5Y����$�L~�T��E��V*�=��X^�tG�\=������Y�����B���7�={����������ۘ�S餧�[�h`o:���|w���'T�	J�J>��c1lnulOM��G�Q�p@\�A�\��^]z8z:�����cm��L'���+&�(UR���O-ۃ�믮&��m�� h�+�h�Qz{ �Z�|Ct��w�z'��]^/�����F��%��Ӂ�C�篽K��FIh�ƽ��q^��=�D��/h*톯R��"�D��|���>�@��W 3�׀��_\�L�|�O)�;6/�ۙY��_�����׈�
�3�o��yqބ�ܛ�y/��p���&E�*8E}μ:\�g׹w�f��r��}��R�ว�¯없�߮���zc��+���9�R=N�F��$fv��O2�F'�zc���qS�p]9�r�2P�ʫd%]��}����i�_z͍�W+�r��զ����O��,�4�9��,�Na�q^��qNp[L�y����[+;��[�;j�'ƒl�u�镙VS��;���t��n^�J[�ᘢiBL9`��R���~�9�ԫi�� ҏ��Vj�y)�3|�}3h��q^��>��S��Mq�NK�{2v2�s�.����u�Ce��vw��C.��$X_,�[J�� ���`�>�ޟG)��NF����H�>'���0�z��|J��O�Oz/��3ٱ{;������.%�.#�C�ᜧe ��-��������uW;{��B�z�{�^T;l�QP9��Q� (I��Ց���:���瘿�]l�=jI*6w`�%���õr^�ߵ��.�3��}S<�.)H]/L�j�@��Qe��>��u:��漎�td�5��{�=\�k^2�Z�W�t��T��T�s�sA�����:��Gm;����u�ձ�E��g��6oL.Ӕx�2�.�� �H�=-�%�m��t��{@�	��T20Y�j��kͱ]�>͓��HN����rx�2 'Fc`In��;+��0��>�8���aA]x��k�z>����w#���n;:�l�S��Tzm�9 i��@J��m�˕o`�kzoc��o@��if���o���g4����o��z�U_.d���x��#]��̫��g�w� ��t�_�:��@=ơf��pھ�>�D�����M����$mn�g�H!��ܡv���P��:�-���X�/'T>G���:�ݏ���b�k=s|A��U�=ѽ�
J�Z%!'��!cB��f��5�^�\zVb}7��A����⺢p�K��˞�DT�ǅ�\�j�t�ٕ�˞�8�u�U�4Cm��.��E+���?�F��
�:���Xj�^ޒ���Ŧ����z�ǯ�\�����Z��p��]�Z&}����(>�m�0�+ˏ�N&<���
5u܇
�S�������x^�9���{��@N�G?Ea�C*F�� d��9����C��ﶘ����X,���Ֆ3��z}��8�d���ߣ�hm��zG��>�Ñ��P�\�����ޛza[�����xM��F�*e���'\7���W
�go�w\�O��8����I�n�jy��{�T��YT���%9.,�qމ3�@�T븬�}�	yu�7�>ɝ�c��DyYb�$���׼s�(�/�L�W=G�9����w.���t�^�}q�<2�1w���	�|'_������������gK3��!��2hr�����z�W���9�ˑ/z�s%B�.�ζsjt<
oLtw=��AV�f9T��H��S�:u!����e�;���R'5r�\�$%����#��1�W��H?F�������;f�-�L;W퉨~ۯ�-Ʈ�2��J!r�����U�Zț0��]�排C{B>��ǐ	^�])l��*�A�����������WW�S��&��Aǯ[�Z�s�zʛ�>Y�L��c,YL*�^�JJB[�����s���Ł�˧�f����a����P��=����ݗ*w�}�O9�Fu�}�H��]��F��.��9#@���@Fߗ]���97[�-'�p��M�FGa��]q7��Y>Ⱞ�8WgT�lWU�7����w�׭���غ���پy<|H��@/��^�-��Sf8�)#��;���;��97�����:���z�N�&N�$�� g|
jh\S�����d;m_<{��5	a~��mw�짪M-Ŗ�'<&.o{�&��5�mL���������Qk&��9j���n�A�Ǖ5r�)���R7�#���%�ܡ���.�{����29�1�{Y��_��ɛwn��p����QЙW���Ԟy�U��Oz��-���v���0{H��ݳ�X	�]2\t;ʇf����F��򮣱.�����I�ˮ��롷ΎL��l�(�WD�����곱�v�_�`\2tm�W��\T���5y{p���������>��\���c�]����XA]/�@�`�/��Q�Ve�}>�a��S�8.)O�e��y����]p���C�eH�׷�Һ�O���F�x��c��ܕ��c<BP�/k��`�{a�쏊oC��5�
�Y����Z�Q�M<������^LӔ9Y����­�C��e=V^�dL��̚u��Ve�z��xMR����	;@���	K�V`Њ���P����t�4��/�����>B���Tj�ĳ)@w>1�&k�q8��9h�`TB�hk{����pzDS����֯�tuK�^u׆��we!q�k۔}gĤ;>�3������ 5����µ�=ݭ�nW�z��:�u.��c���C���Z�w=�
�$�CҠʨps�d�sWv���^Q�#`6z�pq�=egH�����}���z�~�3�]Ô	*S67��m\���xn��K@p��wS+�.�R�L�+ʻ�r����l�;q�WGM��*��]�N]�>�O�7�=h΁!���1T�}>�-��7�����[G9I·���ܘ絞G=�͛o<�s�nr�L.G�Y��� �@���M@cv<��p��L)Ld�z��ll��^�e-T*�v�ZMǻ�����sE�D@j�H&
��7^��0�n����~�ۇ�J�%~�"�y��=�ԉ�@��ɸ��X�_z$����FIh����2��
��z\�n���{c�J��ڄ�-B��W�o��H�ë��M��޾�]_L�$�E��г}��\.�l\z���"�������juDq�c�-A<�R��\8���aދ*����xd9[����u��%F��vm�xy�x�fC�:�]���t}��O]ͦZ[lY�
m��f�L�l42�*��c9n,=\���-8�a��)c����>�*�u��q���ѻ�p��n�M����}�s"�r��*��ET״��]o��sf�mvK��r�X��wR�ฮ��W�K�_-�\?}���Ǳ�WI��'�N���쫷�Z�)es�n����za��X�Oa�,�>̔:�.��U��yӥm�����_b��	��k{�
���rϣO�fc�D	�0�+��e��)�7#Df@WI)�j�o%�=���v��>�����)��N�O�e��~�,'2U^���u�N���q�k+Q�1��#��~ȭ[��,�ݢ;�]K��ᜧ>}���.�C��IK��\���
ǎ+>,��U~�f���gVUq��=#q%�V1���ǫ;���Z������\Gk����檺�~�׺.��<�x���g��t?T�S�Nv�q~��P*Qe���|W���vׇ�9qSs�߰=��O*���}��xe}jH(�h�u*����N}�������`�܇SS���W4+�9����;k}�Y�=w�.��;�i�,��/`΁ �H���^�M.��{ׁq�&��7�<wa1���
�eg2���Eu]�N�Y_N�Qn�ݢ�\n+^��O����ʹ���;p�Ս�(sߎ��i)�b��=�V7���`�c��!H�5��}��5�37*ou��Ys�+B7µ�5�X�|4'���qM����J�_1����ޡ�vJ��]P��W+�My�P4�^[��8_@+}Ϥ��Y�v�ty��>���MyC��Gs��4�Ι�]v��GuQ�@�#���i�A����N嚈�ؓ�����Y�����ϣ�sOq����m�^�q�WƮ]Q,��W��������?V���T��f�qS�pg�|jh�w��7���O�q=�f�PwJ.��O+���y�2)�:v�$�9��V*zw���V����z�i��1���4nŏR� vGL���{}ܰs���b�N���zJ�s��;��������䱕n���^�1�5��q�}�X���
��O;k�����Ī�d���a�WVa�/o8��4���c'ݨ���x!�/_���U=>�P�7�V:�}�Cn9�=#���r�Ñ��P���f%e�U�P���T���#���N�񼭦6%U<'����g�b��`��VI�)�p�v|��\���F���v#��u�7E�Q�9.,�qޓ;��N��}�Ժ��=O{k�^�t]����y�7��o$E������V�Bʠ�O����h���:�Y(^�Z+1�g�nGM�R�)0�u&÷ឹ^=Լ�(='T�bc|9T�mr���W��ĉ���E�0>Y5�|dG�TbAy7��gU3.����v�x��&�����.���ȗ��	h�k��r9M��`+�%ָ��K���m�y�Ǽ�5�	e�p]t+����*QQgĤ �bI�2�GXɡ��1� ��M3B�^�4�7�D#Oº!:�+�t�o��#��珬�A��k�*���e#2x';�;<�++n|�W���x��z�;�b���h�g=�m�p���%ܠ�zK(i%��C�C�#M�|��=X�osK�����3����eĹu�;���gP��ʈˎ���>%��@	��>�;�9�G�]�X�jwX�|7��)|d��WuCr�"����>;�vu�ˊ�g����{�W�m`t&�C�U2��P+�u��P�Y8u�ُGNm�s��3�.���#�T��BX+��[��ؙ��S0_�j����dq�l���!ZJ�a������C{�22���y*��+�Y�O�+�����u��K��7�)��;f*^�Q�-d�9>�^�{�m�0��E�5~\B���\>u���O��E�������L��2�ۧK���8�U�;z�^�u�?n�,׾��7cp#g���,dV��$-�~K{+u�@}�����R�8s��e%�@~\�8�����}wP@m�����QO}=ѻvG��[��_��!z*�R�yE���ۆѕjhw-t�7&�9��.ǩ�L�`n�,��s&N�+�c��D����8W�PW������e��u�W�6���ڠ�fR�w�G�5O���xn�´�K�_^_���>�}@t��ˮ��qΎL���Yiɻ�wSS/9�Hr�9::�N��Su/	Áq��ۇ�S]�=�}�}�U�}�zn��Gz���i\�gȏ�ؼ1�_���k3��ۜO��ȥ?��[L�W�]�Ц���W�g���۴�]4�543}���eΖ<O����ȱ>3�Y��z��AG���a�z��~��FN�~�#�u�@�Us�}Sc0�vR�nQ�Y�)ό�C��{�?>�2&qV�]^��FpǦC�|�[���c�����h_��nB��(��Z>�Χ�Οu;�^���]�F_�=����0�zzʌ�{=�u��>��\7�:���%�����6����<�ww|��p��wTt���}Sԙ�E��k�����'���OQ�Wf7�uR���G�lt���p��t��@�sJ};�`�.��ߛ޶��Ⱦ9�,U������(ݮ3��I�W�J
+��Q�bM)dyY�� �����8=���X�}vu���ѽ�7X�G�z�k�i������z��ح��Y
�E����{,�ܡi	�`�<t��#�1\��-V\��F��Ҵj�f���,�TO���a��>����:������k�@,myu���v7�Ш�$�[[#=���;C{�p��냦������4Y�D@j�H&
��7E���۾�1�&Ӯ������w��b�;c�J'�����Vs�މ��U�7�-$���D�}7����n�
>���dj>�ʄ�|�
�i��6���\ �bl���7��f=n���*&m���!��f���)�96*R�qR��8�n�\?|���<��Ѹ}�n��^��QEw�U��6���Gz'�љ^.}�qg���+�y\*�2^�u>��zc�c讒#yws���լ��l���X9@����ˇ�p͛�Ĩ�e`w=��9�r�2P�ʫq�U/"����w{kx��P�*���wus���KѝqC�������\�Us9���g������U�=�l;w�N��@�v��{��w���ޟr���om`�T�g�p��3Ə*�����d�C�����>J����G���W )cVEĮ��9���)��hv��)\��2��:F��Y^�9O�}�	עEY��|��л.-7�O]m4l�f�@�F�s1���L$�/o��]gi����Y�Ý�f�tqS$����W��V��9{�3�u�D'�A$&D�:�(��|3\�&%��ۧ
qɮ��n�D_ep뚚	���2���T��ɽ2�ӹ��˽��OeN�F)���Wv��t�����\	�)��7��,�ٝݖa <�γCt��o]pB�R܀�>���1�?4��9��_U�����6ì�T�@���F�n����MC՘\=ww-�xFP���B}��Q��Se��.-�|���H�Y����5��g8jډ����47�GFgWM7#�v�]IT��1����/����]Ջ2gI1ǽV�]Bk>�t8<�L����c�t�$���ȏoS�4�l��k�*�e^ʉs�o��,�)[���"E�\��/4tz&�o��:�ɮ��#��i�����f�]H&U�8�Ế�Kj��f$ޑ�C��_n�H#ӷnGk%����c�T&p��y�Yc��!���8�vv��z:�[ObT2��fD���\��	���x
�P�6d�f�v�73/X^JF'��UNh���+=y������_C�]�r��%7u�st
P��-�Xv��'���8vEjԩ������gIjMǕ�ccB��{����t�L��=���*��T����3��s&�Q��9Rp�)b�]lK�yg
�$�v��tXv_Z��_g0�s�r}�/	���E��\���w�sqQڸ�{t��n� �������Ӎ��,]���RĠ����@m����|9��rk2���r�X�^���-$�!��l���Q�l�1�������G�!l�֣�Q�w�����䇪��{�-����o%]Y��eh�mR�@�ѧ�N�����sn2���jeKL�V��Y�Q3t�����
�zz���V��(r뛒�xD.9���y�����x}�J�mF�w)����5�fĲpr^�s^d�ٸs��t��'o��e
J��� ��I�o4�<�N��g��@��-7�&m(��:ef�}�´��2�c�y&a�vv��=�T���M�+[t׈T�W%�+Gn�*�dΣ�-��p쥋�f7f���:�Pz�l��o.h���ovi�/wd�Ɠ�3R�Z7*�*|sZ�6��o/8��:�UcîsK9\��/a�a`N���R8:Y����k�Y�il�dJ��d�ŵ S�3������
h�3���{�}s�T,��ޅ*��oL��lml��`*N��绵��R����ok�!��eVo���j�`W����J�.kq)�3��x�O.{܆s���p��7i�J-^�׶U&c�9|;p!;�M�٘"�\T��o=�Ys���&WqjAQi��2T��%�t�DK�:���u����M\0`�� ̢���G
�NR��05	̃QK%)l�,��Ap�I��Ü�wp�9]�"�WP��WuB�U�9DRa�I\�sSH��Gt�tCD ����LJ9UEʨ�@r��G"+�9�-(I/P����;9QU�@���p�D�dU��H��\����+Rp�f(,�E�9E4K�E7VTr���a¨�Dg(��q�T˄C�<D�T\��"s
9ʨ��(�젢�D�ENM�Eܶ��r9��ԝӑT'H�Ȧ�
�(��IE
�-
R��*�H)�e\���A��IHr��K�r�3���T�҂�(��s�t4�Ԋ'H�4L�#�e�$$�L��Uʢ��Ԫ*"9TEB�L��0� �8Ut�TY���Ƞ��]������/�Y3�^��F���q=�÷P�d͆/a��r+Z�}{V�7}[��C���rw#�i��ѥ���Ӿŝ(�2�:⺩�*#prz��:�t��gz��~��W���y�6}�zH�m�g^�[�'âܒx��:�L򘸧!9zg�P7��,�+�����NR�]�;aN���~��^h����7���3��jH(��X��	��˷4����=��zk-E�Yq���v@���]v�|�;C���4�XD��t	"EA�l��2���8�*��q��ۭ��;��^��9����C�edoP¯��Bp�w_\w���<X�1�'��w���13ut���sԷ�g�z���1���On&��^A�O#�ӣ	�Ωq]v��uQ�d�E%���F3FtNz�9F��Q���P(g_�L=+4L=o������x����^�}U|jb��9�>}����vuI�5���䔧�d7HUԽ83��4�ECmWIP�y�ǧ�OvAUn�O�J��[�n�:װ�D��%G-V*%��uҰ�㑻�C��ܘ��geC~��*�Q���̯{*��^*kd����J���9\	�-exg����d��N����4/%	W���G&;Ѻ�9���[D�CP�1���TWZ�ioi��)��+�M��m��tR����C2հ�:׳��l)/�~��vG������G;��j�c�i|�=��
�:}i���{�t�O���)�ya�/�U{���)Q�^зʎ�����_gPꛈ}<��V�2�Tl�*�L=��a�WVa����V ��ʭ�.�lvaW�m!����[����}#��ʱճ�df��zG��l�9_����O�;��D���,�U��+����=Ƣ����J�xO�:�}��V�#;}��Ւqug�-:=�_�K�n������Q�_��7��J4}.B�w�4���]Y�gϲ�/�6�C�3�4�LK��������/�#�%%�l%���u�r����W��p�\`��/��k���5���t+W��x�_ݯnQ�����= �c�3��S�ʱ�C�+�٥�]LUv��Z���@�J�+����G]!��1��nx��$���r5U1qS)ړ
}��,�^{a~��?h���C����Vv��s��Gm��;O���~ӔY�Q%���ⷊ�u�1�+�Uԣ�}�Fq���A�ﭼ���N����s�Π;MǹQ�Uð%�/���3"����q��77�ޞ�8������FC�q[�q6��G�g8�9�t�*��둌^��}y���X�3��wPE��
V�F�^ͥIz�=�xyu�h�zCeϵt�lw�������]6l�G�ډi�}x#��N.��tsNqc�B�.��L�g1Fo�|vSش_=�b�:K���onq2�,�k�ޑRq"i��v.�싞�C�(��0��U�ue�+��B�V�aq�#� l70 k�B�/O�Ά�u�c�ӛm�_:	�U���ފ����L��n����4.]Qf�IA|
�4%������d?�.��b�6^��~ZG�F�;��>=>�_��Q����>O�3�#�>a�K��3>g݉�������=��7�����.����B�w"���q=���g1Q`gp������6��Dm�Oq�_,��(��q�y���9W�Bח�ɺ�6��}|��3C܇�G:�̪z�R<i�/p_y��?�,V���z<��A�6�(וw~&X���7�\+{�F'Éّ�9����W�}����AX���\2�^��5���J��0�D���S¬��sh_f{˭X�B��+�7��>�g�����8����S���[L
��^��:�4V�@Ʈ�|���,��-�3�};n*~/����x042���?p������ r��aU�q><eO�9��zy �kA/�z��Ҝu׆�����kڎV+K��j|�d9������W�iv~G���{̯�I�7���'n��Vtl�1.,]Imo�)�'����Ȅ痭�s��#���$�m�@=�o4����%��:m�1�`�F�S���p��b����H�����k�d�*6��N�K�z�Y��6��띻5�1�fqP��ЏﷰV2�0�K.鬾�9�:���h_sې�r�(��ў�����������G�3���7E@\^̰�:z�gH�ٝP�e�[����?�.G8X����.Q�d�:	/�g@��ʣ�*e���*z�>�4B�}����z}�'��nQ�˫`�8��|�4Y����Ұʀ�3�B(������}m�	�t�[��9]앧���R?�ύ���p'vu���u�0��Q�p��� l�er��,oc���
�Vm(�@�y�ٽb�:}lz:sm�Ȏ�ZO��������4Y�D�H& ��������Zo���zoc��oD	�u���->vǣ���86�� ����Mĺ�����Z;���>t�3=yݎG�X�:!�ңqq��ʎ�P�
�i��7��=�\ ����x
����>^�}Qf�P�}�so�[���铮n͊����*{�Q�/F�e��&����%�4nu���gu{�^ZR^ ��s�W�����Q�χ\EJÂ��p��xV��<�]w�/Æ���`K�x)�U����t#�K�{\�G���,��6�䚁7��K��d���o�Yt"Blԍ�[�X��}CL4���l4�Qt�5v��;��=8�4�c=����c�oOu�o��[w 30�ح\�<�kA���7Y�,N糤������}���^/{��rz7%@��wC.9Q�6oO�������Oa�q�	�(v5�+l���pҌIe��:#�=�z#;�oOi�5����Q��������}=�{ܞ�� v򼬍����� {v�ؕN�Bu����49)ȍ��˛k�c�2����q��Z��֥�~پ��*��:�V2��cVEĮ��y�p�S��)��h_k���hdJ�G�ً5k���=���vz�B�������r7'�+�
�'K�W]C��֮7X9�
�,~Go2�~G|��c��� �g_	��yL]9	��ٮ/�z�S�,�>�y����Ϣ�]�yC���ΦsiT<�s^F��+��IT� r,z��U6�w��&<�o����H2cbLr_r[�a�H:c=�G���q��.��;�i�,�(���,��g�O�}h˹>=�^�Զ���_w�H�O�<�g\oP¯���7�u��{O���1�+���S��z��緳7^�K	�8�}�ׄ�i�{Q;���s���}�Hi7�gT���&��=9N�qFt�����~&1E9���5�K���;� 6y7*kJ��6.�G�J�kN(e���}���~��Y����u�l6;sfb2\)���1�q��P�m��m�]&>׈
P.ۖ{:>
'b�\�KHO_e84Tk�a���zf����|�]�Y�B��V~���zif��m��}�L��;X��]o�\�S���6�^���M�'G:����H҅Iz|=�����]%|�yǖ,� �g1�3��p4ɾ�^��^�E˺�6�Hj�Ղ��]+\d�5��C�Ә�:��q]��K��ƕ�u٣o��oz!��E}ʏ��?WI^�s��;��^S��W�o:(�J��}�S;�w��^����}w"��P�ǀ��]�7�e@��%F{�0��:q=8^�;���Gf�8�o�6��Q�����%U�}����[>�q��������W�ɛ^X*���CQɌ�������5���T��;�u�x�9Up����]��ȧ~�ep����=�r_l�8r��������0��t�\
���;��<�8�%�6�_���q�&z�CW�o���L���$�˙c�&t+��8.)��#h�p<���v�sٻs�Xޯ�D��+��3{��׷(�,�������,I<�S��\�і�X�1��V�k�lfj�����p;ą/�$"ƛ��ʻ�FoV�R����X ��$i�Lm"�#�{�s�t>��h��������r�7�NN�EWA�f��\��X��(�<G�2b���	�{l���_YT&�܀m������ONK�����z�R����}�Hv���1Gs۞>��$���r �c��1b�[Y�)e������wC���Gh�g=�Gm��c��%��z=%�4����T�{�w�׵� W�Q���P\}���n��G9<�}�i�r�3���U�]|��-�ɼ���N��� �H�.u@��ِCÕ����ED9�����p��\p���}&��F$uf{fs�\�kL�UBY�����a��_J�zj<��7=M��Uz���z��Z�y{%c�*|��L�p���]�̖qT�Չ`.SC��x�
o6&�㻩�j�#��oڕ�Y�6�1�=���q/�ƣ�*;��q.k���d�������!2�ӧ�<h���S�J�'f����Z��UR7��q=���gz���=p+�~��##����ŵ
�����=Y�}�<>����yQ�k彗�ɺ�7:�꿟_��2/9��.�y���{YYS~���d̾��pr|6�f��{O����U�<���O���g߲?���{�"��X��- ��-6_�wƳ���O���ݳ�.2������oGG9��kJ��������v�f����Ywj��]Os�ή�J�b��J��9J@��ކ�%�ފī��fbt��V�B�z�ݭ�F��3����]���q�:��1�������
5��X����W��xN¸�^^�?D����D�$iO@���W�v�⪨�������p��o�����|O�2p;��Q�qJ�i��g���]i��r�W����6����x��Ou�>���w�b�}�:|��fa���,\W����S��Q}���y���=�7���W��E�+�z��ҜG]xn�}ݔ��k۔}gĥpf��0Q�~;=�v_�^��m��eW����-�
X�wMWK��CU֎��{r�fV���t�R��mn��I���5�����dtν�a�oWx�Ǽ�3�)��n�lҠ΂�����W]ar3�v���S:�j��-�g�=I�fAϡb��Ȟ/	�D�Ӯ}}��m:����,�����^�ލ3��n	��'���ȩ��}�`��W�ݟ���S��է7�����h�ܤ�Wvu���]�������fl�_��j)�YNj�ԱS��un�x>�;������Ͷ7�w	_{��鸮���̖r� h�}�R'ܹ�Q�y]�7`�Z]����ta^��d�����WS��Vϸ� 䗛��tq-K�V�͌��]�|���e>ԑ`dϹ]!��k�kJ��a76�*��Y2����G��6û��Ѩ���sW]4h�:����c�vj�zD��sV9닙J�]�G��	�T�|G��Oxt�d�Ϻ����Is=3^�ד�R1?a����[�L��Hٴ���xzk��kB�����}ԁ�� gz!��,���i]N^�<wwˆD��zv�%S�$}�|u@��x�kߎ3��sw�\?%T���_G�9mA���>�#�۾�/tq�NO�ϹׇK�|nx+>u�ü��ײ�y��Q�?pYz�lJ��bqɥs;��+���tS�}��'o��e�*8f���U|=0�d�{�Oa�qNp���ȗ^u�>�n�[���?��~=�������;f���u�꺖r4�̿�W�߯��R�wȷ�$�(u��}��,w�\ ���c�*��>�:���r�������e��C�'1�>�_���v�C_��5훥�}ш�uq^��ty�'��
�\B�U�9N>�Aze���-����{�:�e�库� !��\�s��ze3�<Y�b���w�3>��Be\ǻ�L��z2򻞍�'���_7�B�뭒�"ID��·u3�b✄��.3�؃�Og��/@�O'��9fDBv�=s��e�ks�ot2�:Fs���j��Ÿ���Y������E�Z��9P�B#�M�C{��)���|^��nJ�/iC�vnAG�i�����=3ףeg���g�� ��{O>���wV'W�+��K¼�RH�ƍ�����[���u�o�2ϢԐU�&�X��U!qU<����Mg��2W.>!]�Y��OD=^���u1��x�|�;}׸�h��X�Kt2]�X�ϊv�{ٱ7��c�s��v��OTΎ�}~6>��{\���U�R���㽧�x� '�޳=T8�4m����@_Pa�_yv�M�k�y�W#��Hi=�23~��b|�������Uz�P�F�� nj	g�ΠT��N��ᾶϾ���s�k��m�ȸ��ٶ+����z��?XUxh��P�U'� �@}HU�KӃ >;�EC����~�Q��n�����_����Y�O�+�k�Wu{�����2CV6�w���Xj�%���53�j�؟jWi����Wra��4Wt��3Q��G�
���+��9A�1薲�lN��z�{ʜ�����F�e�ۿ=�܋y�:���'5w���܆T<JφL=�ttۘ��Eř�W�q��ޞ�0����XV�6��W��cЕWi�>��n9��1W�ٷ��ɬ�+╈�(�=VW�K*��FpdiTU�ʙ���Nʷ	�떙ϥ];�{z:39]�5[Wڙ��J��:�+��G�l��ދ}�V4Nӛ�N�e�L�t<4j�s�����6�\мˣ󮾜J��)���J���k Aέk�8-[�I�P(�nJޓ���0#'0f�q.�̥ƥms��\�\r���8sF�(�j�땔��+6Y	���Ì2@`�ͣ��Z�����:�~f(�㽻� Vuʼz��YK(m	��}��P�W�v���	���K��]'���w����[�
[��?V����~�Ap��e��v/X���gn�vv��=KH���8:� ��U1,��K$��z��7�7�[*�E'3u�WS�-�+��eW����%�ٸ�X�ð7jpm�x����V���o��]�`�U�uN�ba��*���7�'�΍�-U�+��}�C����mI�)F��,���	Q���2ۘ\�7��c�8'f�;Y�ѴY���8��x��B*낏e��x�&�iC���㎬�; ��Ҩ�G=��Vf�c/F��w�V�ͧf�,��嗽ւ�%�O�҇�xxJ�0��FVٔ�k��$^i�˰�|x������w���*��ɚ.�9f���d��T�.g#;)Ni\F�-=ʝ��dW���E%��;؛�o�G�ک^I��6u��Gp�{os����^��k�t�05�`Dk
���-Wi�g]�R ۀ�ܭ��E�7G�&�.�>�X^j�z��_6)-�k�.e��t]�)���i�*$�n�����o���"W��i��V�9�k�z���Vec�^�2��:�q5�i���L��#���-Њ��lhx8P���m�si7p���袱>{�����`cx;�Q<�v�R�l��\��l-k�ꗃ]B��
����a+�8MZz�8�I��l|4[V�Ӣ^��3�wɪo5����%�+/AͥQ#�<2��׫9�j	����7B7}�����!.�.5���4�?��t��s�c�ٳ� ;l5���6渃�Es�_[L>/]�B�;�<1v.��)��ol²W';�DW�OM�2f0��%��:Qv ��e�R�[��*��\P=��u�|���ک^S�{���%ܱU���'�E�n�
�w�l�N��c��{��X��.Ҟ�N�%M앝�F�t��-�G5,ee��ζu�����n�'Hmwn��2as]*�Iz�����^�%�S.2����CG�;��ud��x�`٬�8��i^����qPޖ[j���s{r�U?u�k�-��s�]�ھp�yWqeq�EX���t7}��oUw�t�:i�[Ò>պ%�:�_De���:s���B�I��S��t�[�)og-��8QU�3�R"�c�:�Ŕ1�܌]��9��ٝ����1\6o)^$�����&��m��K����y{�yx�""TUUr�ʊ��?����r�nIA�J*"��"���8�UES(9�"9DE"��("�Q��r+��I�S�*�I�TUG"����PTY�r"L"�9�8'NQ�,��DU2�#�	����U�#!C��sS9���.��&gK
*�u�!�\��!�Vq�H�%@�R��4U*���skhp�STU5
��jY�3@��(������eG.r��/5��9��Q�J�(��&���P���$�)ʕ.�"T["ԦA2�13d���YiD�9���iZ�u'0��H�(�* �+"�
8G,�1*K�Ҋ�I�L:�D��Pp�V��Z�r̮s��⻉�(9T%��,.S* �8�P\9�5�*�&.�X�`���*	���J�[��uKks�#�E�e	�������B��wr�_�Yx{^A�i�p�T��מ���U�*�=�J��f)ID���\n �Hظ|�ޔ�,T1?�d첺!�L7?��g�j%��&�<�<O^Z�՞���S���XA?��χ�߱fA�߀���@���;��=��Bk_-�{�������\��o.5'^EvϲgC�>7�x[	h���pG�?r|e
~�[q�nX�������Iԙ^w����a}���DY�)Y�=@Ζ$�G��c3��љt��t�Ց�2���/W R�=|+ϩ�^��C��^F/��<}eUA��n�H��r�>�5�}�^�>ƴWX�|n�xs���Í���>��;o�}lv�K� �r�>�h��=�0�ط7=$����Q�F[72�����mӾ��ry��H��d�:��i�2�/��v�kư�أ��#>'n�MD��:[2xr���n;H��qZO%<#ܭTvaX���h�^����wض�e�]V���<\ �ِ6`7P(}(T��N�v:
����pV���3��;g�s�w	}�:���q�7
���H0
�4.���o��O�q?���ڝ��=�NB-U��^]z�Lp�Yu��˝�F�����]1��`Ӊ��Mr ���y(g;�m�k�����U�x1K;{���l�ev�y2oh�ʠ+w^,aX�S �`k���7��8_�^u՞����b/j�S�/�gy��ت�%�J:�W�B���1�ܬ�����ƣ�*;��Y���!��l��;��Y�w}����X��=E<���AR�dp�M]�M���<sp������̋񳋬�n�.�t5s���b==PR��Ϩ�r�a���������y�U�>�Oy�����e<�s�����'��Ù�������[�c�
0r����X^>�:N�;0����T�&�8z��U�x+z�o����l�(�NW��_�/	Áq߯/nw���{����yVm�IㆵP��c�����ڮ����5_�ؿax�����w㸴1t��9���Y�Gkʋ@s��GҺ�/���>������eΟ3��Y�~��O"�~�iڎU������A�2�t��;@��\���>����t�;���׷(вR�#�5�D��[^Uj{س�QfWU#t�W*���
X�wMWK��C�K���~��KΏ�����y�����=�,�ƢKD0�Fy��&^̰��7��}�8�{:���;L�So$|�MT�V�e�n���+l�j�5B��!�i^i�uY|נ>9��~�5��/�>��{����]܄�wp�4�,�B���]�;�ӑ�.���iֽxoY]��rO�-f�gP��i�k�9��>�q�@����]~����t�}�|����E��>=��kס��3�y�	(�`r�w2����&i�+�'_?lw�M���=��6)~U'����ϰp��~�^�u{�h>���΁!J���/�^���z�_�-��zb�~Qw'?�ͦ<9���r9I¯��'.+�ه������ �@�|o�"��z��f��.��t@:y;�ç�0�6���G��������4Y�D��b�D���\��v��j8;㾥F��)��,�!��O���z�=�3���� ߧ���F=�76�)o�ǚs��L�q�[7�cVӣ!��fT>4�
�&����{����:$����j�s#��n�;徼�][��S%���`���R������n�\4�T�cs���{�{}�`��4z7��ƨ{����åϾ7<�����e<�y/}��n�lN�oW�Uf��*;����L{���7�d�	��|��:8���_�+���8�zhW�՚��g�xMY���~%/.>��=�x���$?���,�O��SޢQ�#]����ǻ�K�(��t�ln�O1E^՗���0*U��uh����z�n ��$LΛz,��v��@qZӛ$�Vs�q�Z�ݎ�%�w�a��˄�D�A�i�q��b�hL�fS��r�ϵ�b]��
9:��{x���a�ytVTs��0����2�쌦 ��m�T��:�v����49)���_v�.F:�^b^CA`S���!�J@³ǕGO�p�Q�%\� ��Y���x{�T>�A�v��M�9�閽�t;S���l�<K��v�\WU#qE��o���tNW�,�������eϢ��+��t+W��y�/���C�jI(��L�wS<�/�r����Bzfˍo�pv�|���9����^�w�������i�}���΁?ȱqR�.�ۜ��h~��א;|��ht�w��rLgl�8�T<���c�r�7�(��΁���tIVk"ϯǣj�MNV�r�>$w�ӌ�T���o�$[�׃��k�Y�C
��Bp�u��{O����Ov������%��� {�c I]@W��eW�L=5��m�ۦ����r;�wRM�vuH��>���ΟD��/y�E�<�QR���F�����^~MB���l��sOq�ϱisԶ�|o.�v(�-{^�`�-��.:���˪%�U%��$��
���{�_��*��͸��FQ�N�ک(�ܡ,����G�.��oG�X�1�x��w�&�ѓv�
�J����ap��y�Óadv������+����	�ô@#��\`�6i�/�犉j6B�q[w�Y�َ�~�`�N#�Ӿ�	B��l8�ͯ'sM@�^꣞P�/$Fv��βY��q=�k�TwW��q.뤢HkFՊ�;Ƅ�^5�{���ɚ��: fp��.�Qڏ<TF��w&}F�����r��s�t��s�N��+0p�;�_�x����M�'�s�tVK�W��W�n�8z5u܋��Pꛇ��N�.�V�C*�%'��P�Ǉ�7�KS���AP����_���M���,��_wn��7�8��eX���t��@�4z:�gȷ^����Cä����ʇu��n��p�a|o+i��UO	�u�x�}�յ��v�iL������;>���k��a����Ӂ�W���Q\J6r\
�g+�>qo�P~�ù�7)���c9i���S�u��ߦq��U�Z=dټK���-*��8.)��3�rql����׈ڛ��h���R}k�}.�+���7�w^3�*Q�d�,z��1>yuC4/��ڱ�w��^��C��DR��Xɠ׆;�+可��#���C����1q���\Q�N�]�Z��O\�̱X��}�9(uL�7E��C@����v��s�c�� �����x�vy��u� �hW+�eb�a\��gs��($�ɏL�7�YyY�֢g=͸kU��n����f�]��;1
6n(I��v�)љ�O�%X�h#��Z�>�7�Wr���E��eҨ�v1�}�>�{��gzP^�N��Dti�b�����d��7���ǳ��Ә�gk�h�$�owT����I0	�^��T�3�+��'���~�'��3��E��{�QX�=�^��,�WB�Z�g�� �bN�1L	�ґ�2��뉷N�����˹C�n��F�m�V��j��_g\���gO��"�&@ـ�@�w���V��N
�RV�܋p3��{7�_:w�Ǣ:sm�Gt���o]�̖P����١�=�U	μY/#�z�p0��DvB]|�A�Vx� �����@���\M˚�7
d��������tҞ4�V8�n��GA��F���&��{��dEF��p��'����3��ǀ��\��*����^��[�W\��#x���J��q'���=P�����M�ɷ�ê����i��&WZy�5Ȝ�GǖW1��\
ޯ�M��u՘n����0��u!.��}��yy���*w-��K��f�'�%	�u#�r��7{<
#�7�Վ_��xװ�8;�X�NqD���w5�1Ǻ;f����=�<+T~�z*?~��b��x�f_m�w���x�?���j?'�w7�޳J�+��'�Vk1.��R}NC����t�s��B�/ױ].�y��e��"��b��T�x�獒���4���jK�{a��%����n�`8ȋ1�T�Y�!��q�����z��P��P��m�O�r�jf�g_G�r�<�� �g]��8����]u����M�u�0�}�"�	X��Q�����n����LX���>8;�ɤn"�	X�`R�hq+�z��:�W���we!��\}���C�{���Wm[��W@1�j�FK�ӑJ@j�TpV1����5�}Ls�#5�f�Fl�;b}אuz�;[ۑ޹D�k�<�|fa�{O��������ޮ�q�9�"�[��d�ͷ��)�y[����>%�C�	*�t	�r�w2�TL�j4��0�Ƕ��nᎨ�s[��z!),�}�x�WGM���pm��3�O�J�ncTמ�Sw���Ҋ�^{a5�{Y���\<6޶�G)8U�TWu�0���x��	ј�v�V�O��s7>���2@����w�-�V���u���KI�w\7]u��ά[��v��n�5�^�y��G�@�	�v��a�,��|�3�{��d���=$`�:jkg	�QY�_'s�{�ڔ�5	n�	��?J�Jz��2�Of��ڮ���R������W��y���O��J�k G�`��K�M�L4��p��H��|^�
f��8�~D>�2��޵&z� ���:�F+�浽�	��7*�2v\/��&�{����j�ֵ�p��̲:��I��5��WX���]I�P���y��'wЋ�t�ޥ�r�(&�|���#^�]���^s�U+�:F%.��9T׿fV��z�گGm(������}K�'۪V�Av��ju�F�}���M��ׇJ����j���aw��=�����'����;�T��G.������~}�m��	��r��EDi�U�{c+K�����k�u^Jk<���8:(�9y:^]�1�J�}��8�vMq����;��Y���:4D��s����3Ou{�7��1�^��qNp��bkݶǥS��	�oO�Mӝ鱘�=Q�d��3m��Fm9�d݃Y�ʼ�F�ϙ����c������]K��ᜥ��#�ӊu>�g���ۉGh�����k/��'mωC.e�ѝ�W�B�����\�����ӽ˒��/v{v�+K�ya�wQ�_���w���;\�Y��aT@���yL]9�E����Ҧ�l�[���W|1T
��Y|}��|W��������7�i�}jH*�3�`)��R.�����n	YG;â�w�i��z�xz#�u1����o����]xC�rQ�GI+���6���01��%�-���n��h+�{]c��e�N����E��W�g���$�]Z9�qIH�F6$oMj�XS/�Co�{7�o�a��R���<�K�juOuq��c�enp2`a���Ie����k���&.!mr�G^{�3����骍U���C�ኗ+���툶��E�����9�wѝC���Bp���}q�w��۝μv/����ki�;�D�c LtAr��E�=5��q.Z�9���:��i������k�G�p�T���K<�Vޅ��|��� q�F��t��<��ӫ6��}m��݉�}�������T:�yN�p��7�k�dK�%�U%� ��_T�<3��<�(t7���;Hf�oq������[��OA���k�W���1e�t�Io�j�DK��@w�&�c�
���ݵ�c���FN�[��w���	��;�����Gu+����@1ɐuǟ�^�o{U&���b�a\]�CP�>��_�};�9w:�T���6�]q^7�T�q���p�ʜl�H�%���pF�>��=���m!����q���TF>��n;*�V��o@����x��[c��Y��X�*eC���¤��x�7����*���qO	�/��.��yr�+�a3�BULRT����ׁ�ʴ��C�;�[���${G��Z����tN���엡��v�jN��^��%��b���5AR�E�c�x��W�8f�+1�x��9�{v*;S����
ݡS��o,�|xV�����h�J�NZ��䱤!�����2���jr�5�{�텣�|j���Ǝ>��I���zj����F�}cu,�����(!�=՜S�սw�W�W�h��GD�!�h��_��߯�VuX�5��m�
ױ��A��+��%Ը�_K�����w^�^�ӿX@HFu���ߧ'VЏ�K��KS���B;���7�t�U��z;�*>���|_T��ޘw=����:��Ώ_o�v���}��F�3���R28'���0���������a�C�c���7�j���K���]atB9GM�(�0d	���\Q�*T�\i���]�s��t�Ix����L[u�*���玣-w��{L��9 '5'@�`P�H��d.3����h�|3c4c�9�����۳�V�vuH���.O��pB.�d��@��tL��<n�K��-��{��\;�:�lǺsm�wN�/������r�7�T	Jn_B��(��l%�f�}Y+�z ��}�C�I�=�Y��=>�n;�=���K3�c�[­@ ���S8��ؔ6��Of�Z=iy^��[����i;.9�$���{�������c�6��c���1�m�c���M�co�c�6���1���cm��c�����co�61�m���6�1�cm�c�6��lc��c����co�61�m����cm��c��ٱ�cm���e5��js�]�M� ?�s2}p$��<*���R�$��J��l�I� ���P�HR�BAR"J��5���������J��)R*"��EUDDP�	P��RUJ*�
@U��
� �(�R�EI(Eu�T�*�D��)R�5! *�S�UB�����	R�JD	�
	J�$T�DU@�Q*���*
UA!�UD�%JR���2��J�B"I �5�keFض)p  YN4�[�� P6(�*��u. )�n�r�N��nK��ٶ9���5�t �t�Z��T�E4R�UJB�B�RAD�^  ��z-T�֝:P�'V�y�QEQ@wJ�) (��(�袊(��(�qIQE�c�QEQE�wP�@�����QEQE��PTRR�R*�*��E{x  ׏B�4�]m4v�5��w8]�n��n�uEw8�5�CLcf�dΌ��:�F�uv�s1ѡ�W`�@�[u�ZT�J�QER�)*DQ<   sޙA��K:\��t��v]]��n̹]v��AZ��ۺ�ۻN����R.���]!]۵ݡ�r۪�m��W�wVs6��5�4�E�r���R��RU"�h�
P�   �K<��Q��:�+I�,�-N����k�[�����-��i�mwZf��Rvպ�r�k;�V۵�C5��Q.�u�G�Ѫ�n����ݫ'lgD��J���RU%<   ݞ�m.�ܲ0۲�aws5����F���ԧ[�h��+�*�f��v�jH��\�˭��]֭�Z�k�pڻZ뺌�5ҩVk�v�˥n�]&$��(�"�k
�T ^   	�悺ݻj����ۭZ�팹ѻ;��sP�-�m+s��[�%�]�봧j��Z�ڻ�8vݻv��U[�%�b�C]�7n�j�]�ᥳ���P���5QIT)B��<   �uP�^U��6��Zt���+��.�7:�ܔ�'C)n���\�Wjd�8qv��ݲ��uu+��Ml�u:�V[ca�۷V��]K�WWT]��1JT���A$�J�R��  �{iMV٭�ʝݕv�v�Zb�뻶�j]p]JW+���R��֮��\�+un�MۭʻgY�,�uwSN��Mc�����wt�v�Eٹ��!*�;(A�  M���[+���γ]�n�Wv�L�4ݖ�Y�5��Y��܍�V�e�vۭ��m���mUܣ2��͙v���U��l�띬Q֕D�[Zso 5= ʒ� 2 S����  �LHɐ  E?�SM�ɐ�T��	�S@�	4�LeTSQ������Z��d�F4T'��j*04W#E����i���7���$��2B��B!!�$�	'�!$ I?�	!H�B!!�������6k���i��x���\FjF3-Q0����Eu���d�1��D#Ome����QK'���!&�̻۴b�L�k2H�oh��r^���V�Y�U�.lYq֙f�6�5kV�f�$ؓ���q��$�Ӵh�Q����P��o����i�ɘ�~[��&X3f�DY���Ǭ�E\t!�5�y�1�-�*����F�MԪ���rc���f���w�e�R�\Rh�(a�2�Y��q��ξ�P-�8#�� t�wz�Sb�Ö`�HS�W��Wy���SXy@$��j�w��A*�Y���M��Yh����ܠ��m2���0��� ƒ�^mKD���;k8;�&�2�@��]h��VŲ>8H�7���'�D283w2���a�e%��U��8t�*�'Y@U��T��=�EL�M6[`'���j��9�'M%{vwV�Ŧ���h����5t���VfHT�6�zؕd(.m�e����3�A!+����1�ʱ��led��G�͸��M�r�ՕIAu-�iȰ<7G)�d[�t��
��*�Y�lM(fE��
mTvE��]�I�{��/a�V]1Kb�մ�J��B��fm��ص��!����ڔ��Om��բJQ�Z�S8̼�19I���Ĝ�Z�AZ;t�5���=���b#w3�HRh�R�E`6�F����" �l��ڔ�ۥ3s�ʸeb�-�䫸�if�Żf*mV�bT���Y�4����Ҕm:��{�&"�ku��_���ˊ�lY,h8�a0t��mʷx��@�0)7!ÅYX����**wQJ˗dZلGh�[YYu���3yU�����Z���24�	4�n�tR��o4�'�6! @��R��v�%!U42�K2nU��^J��4�Vn���SKMж�^��B�Yn��,c�f� �����t%*&�]F�f$��r���S�2�㰋�{�I�зC2��e�%�U3K*�)ֽ��u�ݍ؆T����C/+UǸ,��K���e�ZR k^��q�#W
�+9�+.�+Bq|�髰��Ju�nf�z�G�4�fHl����+A��ib��f
km�{�c~��9�жV�����z+/B�>U��&�5��f������r�x�e^�z����N��nɴ�f&���Ca�-<�z�&-�����6�;B����-TDd#e;��4�H�r���W�[y�I�;6�n�,*B&Q�Y�-dy�[sM	X$��j�֊��Y�SYT��`�ׂ6�6E��n+�rie��q2d{��T�������&�0�n�k;R���b�8vAGm���t�b�ĩT)�4�é+��R��e+���0���BV�ojځlX���Hiț]z�#�]`���k�l��o3 �'6&�<1����kɬ� QQ�c��	xۭ���x0�+1uhR��5KU6�omL����%���+U�J����{���H�U��L�)��l2ފ�X%�;&RAAP�&m��l h
�ϟ�Dyv��ʃ~{�M-�Y3"8{��a[��ab���"��_���8]#1�0�L��,
��I%ށ���+N����{�I��Tϴ�suU�N�%�bd�ݑ�R	W	%��Q���
)fR	�/`�C;p5��C��.ܴytB�n#�\�t�Ս��u�+d�^"������"�U��c]8i�F�k����œd�Yxw/����v�<�"7��� �Xȗ��C^�*fԭ�,;T��rX�oi
�]^\e�٢^3[�%7]6i<�&]1qY��K�[����Rh�4b�Х�n�. �����؆Qv	��f�D�C%�͚hZ�M0㙭��+��拶b�f-MiuZ�ʏ3YB�YW���6����<��9%U��i�Q��8������R��p u��U���x��J;Y��je�a����e�46=m�V�bDe�w@r�kZ���I��%E����`��B���SaV0fT���F�%��b��
��w���1P��]�Dݠ�, �.�Zwz�p�]�n��˻����9�`���GA����[��2ѥ�+��B�+v��F��#�vk	�L
�2�f��
�xT�SS&�Y\��'6��u��+į�k15�$�ѣ)��y+$�P<٥Ed�����MXݬ��YR���h��1i0J5��t�PU� b�7/#�Q��,3Q�D���oe�l��92 ��߱�.ùN�e���Dk�tK�/�e�:7P"��rb��7(fK�]-�l��T�Aa#/n��{�
�ٶ��-�ČⲎa�����t��hw�J�3�g��9h7J��u�]���)�p�`2�pLzw�0!�c+Tu�c�%�.�Yz�\�m$��t���Yf�e	� ]��MPA�����gb,�XQ/>cVT���F��B�˒�$W���n�;Z��l�an���m�#��ՠ�ƱL�X6a��ǎIp�1��ې��Vd?*k�&|n�G�Zҽ�Cx�,UfP;�Q*U��]'���i�)���V�$���	���yc7R�藛f�G�Ψ̐���4: �q"&eKsv���k��{n��(��L�����;ijC�D��P0⻩,�u1`��ZIn���p	�E�yyXL�EKL��t0�V÷��l��i�2�4]+9��ܕt���	KEj�G�X�$��%B�eMp�rM<Nḝ�BYwuw�HīUz��� ��V�$#C�cpQ2@�1�]k��@TC�,��Y�{��I;F���o�Qd"�&.�d%�&�!8B����ϋV���O���R��v� m,��h��D����n&E���8M��{Fe��5)Ld�Y���KTc�%C�f;2�� �ط��5{�޶X��xe=M:�h�Oqe����'մ��ӭ�lQ˽����ثNGb�����%zܽ��&�����ueHfc�!���S[�4QN�폴$�Y(J_&�d*[�6e;�KXQ��,���6éW���ݩCJQϴ=��f��i���t�4I"�YB"6]K6�o\�umX�����F]�L�m�u��^�[�.�:��9&L�Op��
�E�SnL��y)2��p�d�ؕt%�8-�ۏb�@h�U�n]�mK�m8���\c(�i�;�nK�P
U��WSFR��.�����y%�ʻ��.j"�[��(\�!4%b��Z��.�[{�b��A�!�D��{F�ֳ�k`ݣ�[mS*�MŒ����ELZr�K���6�"n|[�0�$�f�I1P���9�B�P���3B���IE���ũǙۉ����k.�U�����GnWB��S`���P
Mխ����M�p[9�FJ���zDi�˪�n�[[�^.�kS/-])G�/N�n��ƪh��d�g)@�R܄l�I�+nL���6iѪ�͆�B�3QՏ�����Yx�����d�Ow.^!�j'���黨YD���v�6�̢\B��f�J^�~W%K�J�X�2k��1�;�EZ��g^ɗ0��,���e�0�a�N���.e#)���S�غȲ^�B���w�&M��"ݧt�n��6�xr��[)Kq��"��V��(L���N��M���6mʗz�N�t�ѫX�s4�q]�9����PlŒ����F��z�m���cг ���H���T{I9�(̛��
.c��M^B�)r��v\����h*��DF�QX�+1�2]�	`��"��O@�*m��yY�J��p��ʌ
�G�CjS�sDmͳ�~�5OnL��t���']dmm�ۺzŘّPD<*����#P55�Ȕ�<KZ����� `;Q���څ����(</rL�C��(JX�.�5#�Y�B�HemK�M&�<%����5��'G���(�+��q]���J8��U�T�	��3jRKN��kH���K%dv%7m#6�Vd�"��5��i,QU�_L�@�t���Z[YuvZ�p�

`R�۷�k6�S4�#�Ⴒ��n�x�������SMfmc�)5�gmeg]���U�I0��D+ЂC�Vhͣ��u�$u%�:u�n�٣f���EbZ�ҏ�ҨܘŸ!�����a�jb�'a�6�amG��\�TFL�e�>cv�4�Jo3չ�$EЏR{fTEЃ�(���R��S��R���R�5mR�4�"婣 �BH�<ۺ7\e#/*4�U�*7%�sJ�72��w��S�yB䷨�·���L]�l���1
�#���o�@�@���%,����yT��N����)R:���i�kv�"�Z�Z���"yW������1��	^f��� �M/��c��fnY%Zol���-؂w��;��r�ǐ�o
��*�*�N|*�#Q�RL�YwFA�:N#��d��^]3��u݊PVm�V�m�5���ddK��̑�t�)k�Y&؈���� v*ۗI�&e�Ɍ�͆pdT��[D!{n���e�46���ygU{["n�ڠ�%��i�RPٺ�2t�	�r�t�j��Xa���r�6�Z�ǚ�F%�����9vU�B� ZL*����8輡��Pv��B C�PQ3�M���n��e��%�ū6$#˛tҺ�vbǗ�YQnJ�H��zX����D�)�:TU�m��t]���@nm�؅���KnV谪����t�޷��Yr��Xh�����qVl�Q�j�ű^hJ���;��r�wd�/x1�� �S�"�M��t��G�Y��:&ks5�b����k��ץ����Z�����V�ŧ S�.�t�`��81�ܡ�ŰS��{s5ݽW;M�ǜ;5
��V�֦k�aͣuu��[��a��-:���0��b�l���O	����K����v0���I(�nq"����"���)��ux�����R���ZZb�XK��!�^R��r�
l��MMùo1^
ܺ�f*c-�Q�M��ܫz&1���u6�#���v�R&������QL����2E/7ZPG$v�1�ϭmқ�F)ٶ!UB�R�`bw��tT4ܻ��Y�-� m��3��Q�Vc��­.�Zja��l9+/���]��#���^wA(n�F�]�*���b�f��ȥ;ʼ9�ԣ�t�սgWz�VL���� �q6/)l�K[h�BN��3Y��j�̦wYʂ�s �ܱ7S�b�A��AP�%f9���z� 6�YW�ʚէIÐ�.�F�퉊n�Ń72�`���<!��A�p]��Qc.���� n�-PU��S��A*�����2n�B�du��[w1ҫ�e�hc�v�IBJ��]d��#�4��k�z�ٷ��*�p�UDwqZ&2�h�ZP�5��:(S�bn����(1Z�dYyf��gڥ���d{O>ݨ�'� Ȁ�]\�d�Ә������巐�uq�3F`N����F���ݬ��cTl�u�'����weZ��Bܽ�*��f����_�*�iN^[Vt�)�4
[ ���4�v�5��Yj��x��0VX�t�n�1R�BN�+Bu2������R^�Z6�ˑ'�ˎ��L�L=���r(��=����jɥ"����u4Bk*7�je�0U����▰$L��I,MZ�.��PVH0���=�{V>���Ű��7m��H�U�E���S�#�0m��a5�A����^�HEY�ݪj<��wy�ZGX{2���%��+���3�Q[1f�ǅI���P���Ȃ�Ȕ̓/�a��04��UG���dL�,ʇr頢���Q�p��.�߆�B�Pb�y6�흒�X�<c]�����DH&�Z]nޛH�jc��]o9]1V_i��EH-`����Ph�֩V�p&\�`7�c����Й/27"4�,�Ҭ�R]�c�o1n�5h�CwV�Q���#�#.�knZ�0ݦ�B�i4��p�畛C)95 n�ʗs@��mnֲa��M:�Za��L�a
5���
3(TxƧO�3r%z�I�
�\�ޑ���j:�� �V�R�2�V�S5�D�ª;54�j��M&�Z�^ާ�NɆ�x�M�G6�Jc�`i��Ш��c�H�@�L�{ ����y��`O��)O�e�V�\q��^7�.�W*·FG����2��	Y2B��� �ڔ�՗[$�k+0�$�y�����A�h�l�!b�	�B���,�yJ���Ѯ�J�ͺq|�e��Wk���A*F��i�H�1��&�Y&^�Zx ���C�A; V�yV�L����Q*���n�z�X���݆�����ڬ��D�q?�#�&��f&�L4r�oX����b�׉�nb�rU���sucAm� /JJ�^fIvA�B ��'n��a�)�XVjdHݺ�)VCH��X��dzQƨZȖ�vZ����%�R��5I5q�L�g5On�=CM6j����]e���Vm�e���)(�gƦ����܎�{��8��B9KEމ���oV8�!!5ŗ�tҽ̥z��ѦO���v�kZ��lBӰ�YOTQ�j�.�Z9j����
�B^T��w!�8e�>�AU�XZ
��썺L�ӻ�T
5�Xգ2^�����B.PBj�D���)Z�|�S+�s�On����Bn�e�#��GA�KI�t���ۑ<������aD�0�I�vk�x�Sb��M�^<��{���JMz/ �'"���m�q���xP[i�3���B0�{YnF��$����	%���sM1�nlC/����ݬ4ͷ,��]B�b-owL-��c�%.�/��FԜƸ�#�`�X�^�U�b|1s_*zY�_c���F���٦c�cn����a�Sl���V� k��憮\D���d���EѢ�_fv!P�2�--�պ}�L�� ]bÊn�T�P��Iͻ�Rԑcy��;/���հJc0V�颜�-]��<�{��R7���TB>yO(#hP�(���5yyPrn���hE9�}����AA��t|����)Ei�du%����oK��{l6�^�{�e�˝Z���G���q:ۭ)�oa�Ǜ���N�+T��_�P����/�f�e_H���|�I!k���Iׄ`�;����5��r��P�[+oon�u׷����ɀe;IN�/jY����uM�qe�أи���z�9\�G`m+��<�v 9y{ӗ]���S�����vM �y�	��U_1�oBg�*=�վ�����Y�D���Y��m����P����;*���蠪g7���̤����Y�I�ܻ�1�.(%�9\�͎��mf�l��=�K���R�d*�����	QA�S��:%`X%���Nz�6�2p.r�C2�.��{b�s�X!�+p�ᵚ�z\�ݗH��#��%S; �r|�d��r���m]n֨�t�w����9��7D�-��j}:���7V�z�V[@L��wK��s5�ӣ��W�2�Nl/�'\�i��&m�]Z�f>o6�	��|�I�b���p�SE	���&�`���6��h�Ꝅ�y��%!�
]ݫ
���t+c9����C���F�Z�0�Ŷ�8
��Pv�e����Y�0u�XF�X4d ǯ��U��2�>���VjK�fi��]��)]]J����K��a�!X��lz���!�N�쭴�U�g=�)S�m.[|m�oy�Դ����N�Xk��34�r���U-Z�4}�E�u�T8)"M@K�:���A�y�֬"�KB�(�u��k���$u�}y�Y��i<��ݲc�d���xV�i�Z�kiV���ͱ;q%�,y�;��E�
���Xu��u$2Y�ưn������J�o��qڧ�}W�a���w�泈�9�۬��v7�Ul�΅e%ܜ�ݽx�N�)��Z���b�(���.2\;0@l�W���n���J�R\�D�֪:D�����4��n���*kU�AB�W�n�P/rT�*7tlv��q�G0V�D���ͤ��g�w8�����٫�GKd�̓��I��_ڹ�0�g����Q^���j��ӉfL��9,k��Y8�@!��"�6k��Y'9)����v&s{��l�R���[�}\��@ϩէt 1�+cۭ�$4�k��x��p�Q
vhU���)ڕ�ݡ�Lc\n��(w����|�ޥ[��d����‎csN�i�U��N�K������F`��^b3oJ4w��Ý�c��ボ�9�>�b8�a�wn�����䷍�}�ؾ=p-`te��!u#���+�Z��4$��q%�D���� Sf�/:�R]rP�E�,��SF�;�r*ӅV1B:Ҭ�k*9^WfI�95�y<���_+�m�z�佝�e����&��٣��2�����]Q�Д�Y��Ќ�:�U��H^t�\�o^�Ҵ)�+�&��	�p��5-�-áq
��1nE�b�1�ms�sL���\�
��b� e7W�n�W0\{�w{3��Y����>�傻A�\/���"�~u���ħ��k���8�D&�V���L>�������Ԟ�U��Mz>���vn�۳j=�uu�b���їEպ�!ᷛݜpZ{��鞎^C+�l�F�d�F������q|�X��ĝ��J���9���n�������D&��^r=Y��\NԮN�\	w9�^f�5�[X��VjG3��X�L�%�7+.���k���B:�3p��lM�;�34b��S5�m1���,�(P�yAf�Kn-�J�ye�M&(_$�Z����{sWP�N��i�ڎ����]�T�zhv����T��b��h9�ж��(�7��es4��w3��e����<6(�(�1��;	�G.�<s����a,Y�9���	�[=+ ٹu��;Ҳ��{Y��Z�����֩R���pڡ���B�:��Zt��6^�NX���׼=� �mK8�a��?��ᕣ X*U�)��7����:J[y�f}yyFi����V-sVH�vkZ/e�md���p�l�^��J֢/S��CKs�lWQ�$dRg�.����*�CJ�� ��+�#���h�͆��z�|gP��et�����{����mͮ�0�/J�\U�t<S�+)��^�r�i�5s��a�z��`ҙ%ɶ��ͅ��ey钣7��<�q��p��f^a�-#����Z]p钇N���K/F�2U�d��)�#��`��{�v�u�-�OR骶kUإ�iܶ���#[oOU����"&,���'	�n�W�K;�v��ve٥���l�	kǵ�F�U���m+��3��"S�3���i:�;s_i#5wQ��A�y�U��ӌ[Qpգ��c�ܐ�-���^ٻξ/NԔ��MM�J��,V�o�fB�1r��t�a����9[�k�q�=`�#�$^G��u%r��e�OV5���r����!��s�ㄪ�f�Y�f�[���\�8��d�3��d��Er�W��]����T0+Ia�U���ʾ��ق��qe���D�Z%J�<���A%흴'���H)�Tqs���#&����Ѵzf�{�z#���q����#�ԑpv�&)�1�X��
�u/o�
I�|�N8���f��bޥ�Q���(����y0�":���%���X7A����\6F}O�H����1�ۮ۫������j�M8;M8����ݧ���p)D��ue�K�1$p�dh�����C�Τ	�;5;ds���
�諵">n�J�Z�k5��H�GóK[��W��X���+[N�)e�І4�qR�s��Ջ�4d\�㉨�[}���.�%�h-�X\@��Z�)��/��ެ4�W4-<��λ����gTf8����*iP��&K;��Uk�a�+��W@-c����LvL'M�M�����0�I�Z7�����[���lk�ʆ�Kb[�Wtw�p*���[U�"�Rͽ��b:�A��ao]�����*�Y[�(�����u��v7�)�LwRw-�W��ڵC$[4m�G��i2��ce��ݗvv����d��ȶ��n|5N�Fog�RǙ��P�+'IQc����p�>Us�A�$/D"V�`g��I�4���y�W����e?�L���Uk��n6���8�����s,�w7.�dGRj��a��=�n�mIRk)q5�ikc2��)XV��M��T��+�Ʒg��=��h�35��|�w���5'tv�/����;qM�e�ov�Ļ5*5��Ç�u�ʯ��\�7�4���'��7ܙ�g�/�3�{���՗�W�+9����n�G��I���8�kh���*�E*٧�{NV�P��}5��(�J���O3��.�7��r9�s��K��ض��d�-���h*�>k�(���sV��a�"ˀJ���ap�sj
Q��־�wT[�9��^���&�eZ�{j���٪�[�f���Sy�j�Tl����*c�za�����v�Đ�z�1^J�7C�b��6i����an;��%���o��xI��Lx)���|���8L��B�A�mX�W�U���r3�+.�P��&#�W��bނ�%_>��r��ӳ30��Ĝ���F��w�w:�s8skpv��I:��jL֦��L-���ͩݕ:���x�^0�V�v2�<��;��.i�~�bJ�5%`ޓw����!��U�W!oh��Pv�����o�}�`N�սәn^͝��Y�I�$������I!5Ի�@^�ֱ�.ot�44�h��ol��s���5���'z���y㙃�85�%2`��%��]��,����sN���%݄�n�����Hx�	�])�.櫳��`u�oa��1y���w�
���U��Y�$G홶:U%�f��e��L׷"��yw��SJ��%Lo��I&��r[kf|E�J�c]�W]mP��l�3\���[����<�r�R�qh._gnf]MO|�|��9)���l;X��ǲ�����_9O�)�U̼/e]��Z�	�=�K[�h=���LqH�wS��P��t�Ս$�3�й-�9���Kw��X�P�<�D�1�k�Gnbl��P+�mƯ��9e�8m���������bk�kҹ��k%9�T��w`m�R-���3�O���S6�Yy�16�?g������S�>��s�I�9&���em��n�M����S������mrd��;e��-8HͶT�y��@����N�J�1�B{#�+�c���)J�+�q
���G+*�(�^�q`[����52���۸���/ gt*Bv�:d��Y� �-і`Q�<�#���z�C�{��h$cP\�����޵�Oq}�ڂ���z�x�=p�wRrc4\U+�n�/^\������2�<5{�+Zˈ�c.wtkN�� �AXe�V��o�p�޳/�<s����H���T�b��8ج$WV��u��8V��nf1s������}�%HuJ��z]�h��We��R����rt���V���OEW$�;��������η��T���vkD�Y��'G1V�M��+wZwN�]���y������
��/	��:Ŝ��I����wS��e><��v�T�k;ė��M�����۽YV`���9q��5�n��\�P�Μ����v�Vt�P��_��=+���k�R汉ޣ�>�Z�7o�	+;gu�ar��]7�`\ei�@co���f�^A����]dS�\M��m�RԷ sO
�fJT�1
�Wvn���M�s�*(;}z���OP�wWT5�!E��wi�D M�=����Hһ"#�۶B��l�L�����&�,�L��z6Kۍ��]Z�}}F�Tۢ8�]�lY0��գ�T���,C�cᘃ(����9.i�N���>����TV&�̳a;��������*멺���Umv�\n*���D�(jGV�<�T���C�i�XT7^+�N17��Nn��v� y9s\��̦_e��H����J���kW1�T�Vbwm"au��z�Z9�W�L�2�>w�s���F��֜������<GI%����r�1M0U��,���M�x^������,R��c���5\8�Ӊ�í��D,�ͣ�ל"�Z�{���N�d�̫"�j�,LF��>q�و��b:�H��k����+!`�´˭ϡ��G�d�T3Cm�ھP�i����/�m�E4:������U%uz�1B�����ǅay}���u�Q�VEb��[�AS�G+u�u�]�k�/2���u"�miͧo�Ax慜�;Q�Z]�3fn4z�T�\��EVB������lf���gp�Q|ήǯ�V�{qwsJ�'g���eu�ԃ��nh�|����I���-RT�wW2�8�p��t�soS]�X�(��;��}1�|�\m��]�$�/*�J�����/K�6�u&҉�}\��G� ��(s%͞����!ܫzhV�(�嵹�;(L�ww%HH�����c����x�%�rw.8�uXr�s��'�����w-�Z���W�X�;Z{�����o�fs�9���%�O;�U��%YCb�	�L���#�J��DV%*c�1ʲ2Wy�����0����P�y|�gk/�7&u���D��	Xxe9y�xs$<Q���"�	Z�r��c�&�zË�\GZ��Y��na��o�b(�����X���N�ֲBj����;�Ɲ��$��^!�h�_)��s+&֮�3�'�J�]\�R��WG�[�h=�z�0ђ��O��H޳[�:�P��h�a��otIݐLՌ<X2���{���E���Ֆ.��pTH�s���aU�D���6ٳ-��nS'aװbh:��e��o�qQ�a
{�'|m��)h6��\�i�ⵝ�c��-4��d�,��Ջ�ܙs���D����������[c�����s���s�'K�4g��QrL����S��=0�Rf���*��؛�U7X�4�;ْmSX��Z��EN��դo9���w2�X�59�l85�͉.�-$!��_�Z�K�.������Z�7A����ά��Ek�л}J�ޝx��Z]�V�񉖈\�k�MY��GT)���L�Av^��8�f*�CbɎ,��eK{`���oT����9t@x�wB��K.fM1��Ιqe���ۮPkS��R}�fd�o5E֠NU��G��X��U|�>tk����*��b��`'u��4�wT�ݷ�������`My�J#��Z=4I�����qcr��O�7�Z�S叫���^�㡺\Շ�ǵ,�)�l������5Xv�HX��Z��V^-����$;y�qm󛢐��U��X�`4�G��9��51Fs�{�)v�&hr[ղ��V��d�r�t��X�ީ�A�b��˜�.�뤮X���K_ol��f�#m�%��WtBn�(�u^GH�W�l��`����]�-���P��ۥ��@�aΥ���/��Ya�E����8���9�v���Z�܂m_i�0��5�@�F:��N]�D3
�@`t�SM��/��Oc��ᣨ�\��d�6�7г��R����VK]Ӛ����2
�7�9�3��6�y䯲�W:�d'��>��i畘�Ҍ��:�5�c}��Y��E�;��bXV��9�u9��>�9�>t�tr���k�T�Jn���:����N��_< �s�=�u�����		䄐�$��y�?u���%S�;��
++#��ud�V��lS^^4�d����N�R�F�c�Z�ם@��	uά��P33���Z���(�*�U�1)e�Ы٭Dwfa/^�]1]�dR������ǡ�dU��e�T!5hwS[go�Bx]�� 8�Ԋ�q�Yn�4Vb�iV��쉩�����f\ړ���Mش|�e�{J��X٘D�,oТx��]e��WP(��s�nTOK.�^�7�R��r��'��́��z�����)[V�­B���sq�o,}�b͍7v�P���Qg�m�a-p�z�L��{�i��aݮu�Z8��"{��sZ��p:a�v�=�"]��� �#��Wp�m �۶$SE�bw-�6`�������,Q���-F�X�h�;v[؜2P`Y�F��F�suګ��r��	C��f�J���HiK7H6��>3��[�"t����F�7�n
�+^��[i�k��5n1V̗��E����ux� xJ=l���I{5�DHjVx*(N����v���8FI�����4��X�����\m�*b�� �aRnM{�w7t{.�}q��jp��]w\3�]�]�7C���ekeJk�����od���_٠1QP����	�z��g��u��0-��Y�:^n���`��M|�[�r�^��n��N��{x���:��.tf$5e��g!@�)\s����.�\������8����X����*ʖx�l�Yj>T;M[+���j͗�[|(i\ų*���������_[����fldo3�g4§gj �fI�i�=ܪөu��J�%0%ZH`5��x1E���f�]�d�t���a�>mOY2�YVӖ�՘ͨ`黗PnP����=���Ýؖ��6�l���b��	˷Q�T{{b�{1�Ks�.;{13��Z������W'o'˶I�<dP��t�
�YF��:a;�VkY�*"���oPH��,�/�(��
꽠�'5�K:��r�qV݌�|�������[�2bԝ�{���ӵ)���0o'}2:)��a��֭)����4��3�.;���18Q�M�SDV��[ܡV3J*]�3�+��e�yJT6i"loF�H-��oP���bs6h�u���RT�ɭ��΄h���dZ��[�XTU�:���F �m�R���ʁbj���K�8�J�f��ոDe�R9ׁ[�=�xLS']m��1T��ۧ�uoC������a�-6h��/��;�h;Lϋ�(4KKhFt���`�Z��v�0�7�d*��N�d�s7C-l3��d�;=O{��e}|�xv����D`v��)B�[j�i��� �.�p�z��d�[8��c����:�HZ}+&WX���M�8�Ci�mҾ����n�uu	͗+rӈ���X���4����+��v	)Z�kU['�hl=s��|zܻD�wC�E��t�S*�P�*`a�Z�G����X$��c���1I�q35�m"~��\�lͅq�z7QyW��f��%
U�v�3�.��CI��;t��]���Q7��;3U��g@氱�%�r"-�4^�b����Q:l���i��iէ�v,�L`�9*u*3��;�"�r�0��:��N��.o5�jM�H$��;���W�A�C�q���G0�j&��R�n���N��#2P�(Xƫ���Q&��U�\ן&k-�m�rd��]v:�s�̋��5ܧ��A���6�rT6%��j{m5��������{���+_
wA6���.Ĭ-��9�C�� �mg�����]�:=\���ҵr�\�ʽ� ��6�h�(7�Ι�i2��P���Q꿺���6H�X�����Cw�{���#F�Շ6��,dȸ(�\ޓ�j�Z2���n��;���t�b5Żʚc�(�����X��٬h��>��&�Vk*i�p/��u�Ry�!��񾱠T�MEܑr�Pʱ-�����\xK� zt����r��t��%�\�2���9և���:�����4��օ#��|�R=�Tu��6�*Ȱ�����q��ժ��w�u��8�r�9����H3X-���/U�b;wԺueEvDW�����鉀Lۧ������;��v��+ݭ��̘(.��9xҫ
�F��3%h�����TK7%�Z���ZV�\�d��%-k��ZN�:ݽ���pЄyX���L�u�._4��٣Oa��`�aԄu��/Ufml��M�hO@��X���]�VfY�5乼�!O�I&W-��9C��<�zO�҇�s��;�%H
*��Ci�@^�*�X��t���,+�ks���\�b��r���d=׫X�6��n�E

��S/��0�[�)�d��B��83�^��
�dX��W�n[Z�4�毞f7w�p� �e4��ur��x8�{n-A'b��,���1S0]�Y�T'�r�ԝ�7��"���iU��y�)�)tl�:�`�.�☷��ja��=e)9��u�n�^u���ń��쩱OK��]1��t�(Ѝ��-�Hj����.v�y��'�Ŏ���=�R�TT�|����5x2:VT�nI�W ���9eȭ:b[ݺ`>�N^T[t�̶#���r���P��z���3k� �E=o��<pKݒ<J��-Kh�@�U��)�{I�nrx�*�u���}n�bse9�2g�*��ʻ�W�Ø�b�4)-jS�/�h}8�Đξ�%�p��o��0g! /�q��PA��X%#}[IVT�;�#ħ�
<;"B�P�Ƌ�.q�����6��r����+UC�,e�F�+��l��Z�K���4�Ŧ�8�1xn>���v�SY�˰��A�f�
z�t�ܺm�;�mRʬɣ%�WҖ��NǬ��4��#ܔ5���.�g;���k�
s�/aIr��M�Z�Ct��&=��oVVNӵ�t t��ՐuCXf�.�nZ3`g:5e�{r]n+.��*�2u�.�.n��G��nm�5tO[�)t�^�U7[X;i�c'vG�U��/�[7���c��o���lvl��T��lɢ���+�����%@Er��7Phwή��E�@���i�{O���!����Nc�:���h�p�K+C�(��l���왅-�����[����Y(]\�v�o�wu�0�;��v'RX����w�ׄ�Sv��)������յ0M�L��5V�8�^n� g5�٬�t.�E�YnN�����ur�s�'�PLv/&*��_T�����q:�D���:����s��%r��v�����J��Y��w�Iٌ�Pĩ���YC:7T:�4��k!�z���[`;OrYL���;k�;�J����x�1:�-W���_,ԁ�.��
�����J7�
]w�V�:�ܼ�a똫k��/�z�=<�9�T��j��P������� ]Xu�!��E�#��肽,]�}8uJ͸n\��r��t|�Ԭ˭ԻM6F5�C�uyE�:��X�\X��G2e��
�Wln8p�x��>7S�����7nN�
k]��[��@���v�{s8��hR;�IY �n���n�9G�wm&����;=����p�
�3�2CZuV�jb
Π�G�Z���/Qi`�t�D�C#{yj�K{Q�U +8վ�(�FY�P����(���,�_in��!���not��
u]>��pa��u9]twuq\\�l^��ݪ�\g.�v�f˔�˷w^K��[_;j�6���pc�(�]�%T��y�8!�X31k��<�*���G�}�+C��o�]����n嗢(�����t���2Da�ܳWe��ݮ��5:qR�%�ݼ����N�S>��(r�Լ����"|���r#&���4n�o�!R.z�*QqY�y���}Hvloujy�����DUvV��+��X�]�TIZ��\;���]���'B�	OL��]�#���qN�F��uiE�t:1AiZ���_v�XF��������
q��uM!P�W���]\�AÖ�v�7pq��h�q�y7�re���V]�*���r|4�4���V������܈_XF�#V՗/�|�\��ݧ\f�׉�rL�%k��,�ӭ���I��6��}W�ԑ�җ���W+k5�{u�l�$)Ʃ�<��ۺ���%[�
r|(�%6��-dEK�:cđ����XxSv���,�6��!�����F�U�@�s��.X�$ذ�Y�rܵβr9	w�l�U��0N�e�n��J�;@�9�(�ûV����x���H&�wdb�LM�u�x�V�%�!H�3�;�5M��fZqf>8X�V��vk�*�u'�hd"H�l�X����V�1�'�w)(�u�x�RYyb&gFF;c(F����/k�^�R�X��&K���Ңo9J��rçN�9w�wn�gbi�c�1�*ДӶ�9m�:U��f(����D5Ո�KD`na��mn;���<��G]�_,�w�c�¨��|�b@JU���#�#2��ӷ���c
�-n�C���@o��ti���SS��ݫü��[����2�-��Խhs��������Ow��Z��䫧�h��j�٩�:fmt�_��#�I�`��M�����k�闵a;9�n��TʈE�F�N�Eݚ�;w>�G�.Hq�{�U���SG豥��;]�P�3�LU�nn�2�m!WL�]f�p�ȗÌ����1��,јh]����4պ�7�s¾�k��Z 뉹�JCsLW|�>&�9D���$n�bÈ��M���3GHᾮ۰څܥv+j�K��G�X;v�w,깰��cM�5�x�4ʦ�ofM�;)f��%��f��;�
C����8{k�� ��g$6�S���GWb����s�AV=�}V8��X֜���$��a�2
��fZ2؛����s���]�`q����u�x�'o]�C�B�ޮ�b������Vrz"�IR�SfY��f�BE�[W���2�$F7�qrZ�S��={�-�+f7�侒��gT
��}ptf�f�Mq쌣�d��ܫ�#=i�ˬ�����-��5� �KO���vL�g����Q�r�8%�N��Y��It�F	����lJ��C(��j3�Zs��t�X;;+�8�%H+N��G���m��&����k0�?0�	oRx.�
OͣPR�F���y]�[O1>9�#�3�����O3*=|v����U�Pۡ���1ݫ���mno:C��4;
�Vt��Ae�0`}���ss��O]�t���*R��r�%�%�\º�47��[30�������i@�}�(X_f���u���mokrn����J�a�w^��m26
�Ŋ���"rnvS�n�#�jv*uE����NL�����m2�ě����'��hEËl�d��HM-����oS�7i�����E>2�+��̬��lW±m��
щ��U#ʜ�pn]݌e�q+�I�x��=�����i[&YI�oE�𾝥AX���7wR��׫��.=޷>�ZBܠĲ(�pwe����,1Z���yAv�wY�
���!E�:��̜��-���ec8�`��g!��me�U�B<wV��чt��z��ˆrm�\�S8����.�+G�(��Ad)�(����� ���Ta;p�8�i%�쌮����]b��ڮ��̧@�1L�W�j�Ax:����W)�W)��f�=m�G�\�w9�.�qҮ��W]�gi�B�ͫ�kp���(�K+�	��B��w�Al.���ˮ�W����D&��YN�/:�KM�E�c�����ɝ�
��"�l�u��'th��crl�����W�B�3#�F�hn<4qԳ㴁�HQF!]��=�*�spn�֥�1���-�[�M�t�ɴ�M�jX���i�n�'��%��u�n���nVc�7�n�Ö�_R
���@ss�)n�E�<|�8���i:��ʺ]�l�D:����b^ō܆��Ed4eAΜ�t#�}ų�P �tĜ��<�ZY�gw}ܩ�P+ucDŲ�:����Y�d�] ��%��'�rO�ۗZ�r�b/�Oo��z����J�'8�K��N��t�օz��x6h�kj� ��Lʾ��,����q0rTʕ{��,-��ʃ�i�f�;��q/�P�Z�_QA��)vKq)b�{�^Z��z�F��Żb�g��X%=���twS8�`���j���0d�;X�fGR��ĺ�O��l�U-j۹{�Ү��LP��,?�v6�[�P˲B5jV�ʀo�Zm�;������U�䒚�p��1���)&w�Ţ�̷�O���$U�bPGDp���{�hُp0���/�9Nw��;B�"���k��t\�ٸh,=S�2�)_^J�	Ӣ�qa]�oIz���>v�t�H�z\�C\f͒���Z�6-k[⩳���bp���+;!�Ψ��q�mI�����p;U˸���t؜w]9V��l�jh�ܻ�n9+F����b(Vm�:�˵E���F�Ѯ�a�Y���ql��]4ӤЩ���2{t�O��ׅ�GSWx���l�d֜K1����SN�޴�7�n��I�y�@-5�{������%h�iI�k��([y�Ō���K��3��w�æ��v'V:�+V���q�R��=S� �`'�`�uD��z��ws��B��%�����׉%�Z[jݞT�=��4z����8��ɋ��H�e�l[)��c�aX���ck�^��uܫ��NWb�{Hd����
7���dp�I��)es��zc�Օ�6ֺ�/[ߠY8��	����xx{�=r�a_;�-y
��˽�y�q<��KuƆ13��W-�]P+�?ͦ#��ST"ڜ������+s�T��p��9W7"�OdI�dMp]Щ��'�;�T��oϞ�@�3��tR;�oTD_VK�F�t>�R��sP ��]�OC�lK���p��oҒ-�I�ߚ�̒�f�r�r+w[�'ͣ1S���R��ڸhu�f�4/2S�f�FD�l����gP��A1�XC��!k�d�]HW���t+"UU�X�i��4_j'_sm�M;�/���+;��|yW���կ��s�zm�����	#X�����.Nw�o�C��Sl��oj�\d���b������!Ӷj;וo;�M���;�f��k��[,���q��@����Й4v���?b�ƥr=��:���f^3��Е�
d��\CU���kP��[�P3�=�CR�s5&s�#�N�[:P�o�'P	�֜�|����l�:���v��=ە����U����J���A��;�MN���P�U��[${��۫m��
o*��N�N��vf��%��/���]�t��`�U�LIv�f�qof�
;����L�>��ut��J���;���:wRc 0bt/�v̻0�&f�s��6ü5($����.�47���e�"��ٷ���ln�Ջe�p�Zm3W!w[mu��w"��<��^O`�|6[QAYm��-J1�E"���G-�8�m�QUEV(�DX �Kce#kQE��b"���UrьE��V����X��aY[l��1e�DQ�KTE�(�X*"�-�R�ZTF[P�F�QH�iYRW(�Yr���"�� �TIP��)IU[hґ��B�F*�+4F,�T�1"	
�+Kj�Z��1W��(��JeJ�U��*
���+neT\*�j6�#il�Z�Th-E�F�QdR�E�Q�e����*R��fF� (��j#hڃ+PT�X����6ت��B����*���"1r��mF��*��m���[K���-h�����G!K�:��E���C��{�E>B�U.�3�˂����`�A���y�U�	�gjW�GV!�yX��_6.��/Rv�ɻx����x�:fvW_ܴ���G�Ѩ�P3`.��5�g1������_�4w�w���o*J��t�d�QJd�:Jy�sڝS����9U���[A½l�
m�5O]�ۧeN�Sn��N���U��0���*��2Z�#����
���n���O�Nw.�YI�	L�]`<_�[l��ʛ���y�x�W�A��v�,��2o�}�r��a���7�O��M�kEf��%M�\3%Z7h�',�rR%u��G�:7^]{˴�n���2ͪ/*�k�t���k'e���w/s��I��+*�{S���isj7t�o�ݘ{��B�Dշy��ww�{}[`�ld��Sk�Z����2t�0b�k���%����z�t."��OÔ�N�/�g�'@)t�t8��{�pm<�/= � D^�w���68VQ���4���eF-7E9wP�R�Wo'�������9��u���Td)�J��;���%4"�;�Fۮ7Ru�	�]t�k@ݡ[��
�w)v��kB��u50�4���}�����%�z���y�g�^Td�u��"u3W�"������M&�^��Y��D��.�<��l7����=�������E�k)�c��SQ�[�.������n���+�/(vu�+|Y�>=��Q��e�������V���V�X�f���������ڜtu�9��6E�%W��X1>��v9+��tڹ����;"c����B%��R����2���=\Un^O;!j�;ػ޵s=�v��N|��b�h�394�b�k��e������}l��$f�v!S��S�4l#~��.fΌÈ^,jh:�VN�����+��gj�3ױ�,\�y+��xMղ��4{f�;�~+	uîD-��� Ue���\Vg@�[�rs�b3�����b3ܚ��=��新�+*��;tr9yI��.�Ԭ��5��ά����ê�ښ���Π+X����{��|��<���V²Nػ�]j��}���]J�PF����t?u�����ޚ��v�xt�ނ��N�ޤ�9sR(���#ue6��=u����g�W)����q�r�O��f��%}�)�I�=�cݳ�9Y/Sf��f̕�9:�e��ꨆ�ɦ9�d��w��׵1��k�3�d�)��XɗM�w����R���C�MM�x������&����'7[\��^����Y�Չ/WryO���� 	օ_jge0��U�;{i�m��wNr��S`��69e��n;{�hY�-|=Ϋ}�}�8$�2�2L�9�Ɩ�07n�r����xҾ�<[�=}��^W"ftm?&���%p���oCw���O]�|�Y�5���=�%uȳ0���x��7�]�n�k������'�5�4���������D�14�zMk����دV1�ss]*���<�f�j�,�����>���Ku�^S������g�I��y��J|}Of0z{;�gE�N����ju�oi�lf��B3~�M�+�o�r;9[��Z%d�E2f�w|^Gl���	#@p֦���Zw��g������!3������rr
�+܀�9�T<Ђ����pt�:Z뤯��2-L�wS8[ב)T���K���b�V͊N�HX�#��V����X+�(;�뜮�ݕ����O7#y������+,�h�KyP�:*��GL��5�+n�&����7�ڠ�޵s�Uz�B�r��(6z������`�%��u0��BQ��6�ͩr���:�v���Bt� �Xk�N��I����ؕ{܏*�*���D5y~�.���y�� ec�A�Zr��1؍ڸ}9��)@���P��`/$�.iH��������m�'P��g��^~b�ʳ�4�ܟ�K�һ�/(�{t�!�};���={�yj�e��/6�ޤh<ow���n֩����\�����[�1���c��;5�ʇJ�������㷻aU����u3��JO6<y~���/3�+�	|"8��/��k-�[����ګ+#!�^dô��X�\���<d�	���}me����%��"�ln�[[���FC�8T�F`qԕ}8.w ��r�'���Ug=MΠ%�5Һ��H���O��q�� N�ut|�	��Ʈ���:+l9$ۧ��#\�����º���^tR��ө�R�Dr�K>�̋���AH����!�,ض�:d�n�o%w�7U����@�Ɩ�Ԯa{�}�7`�7�u5��w~w��y�`��c4-�����G�Şk#�z�z��n|'w��r�uAy4Fq/p�%s���7����sa����e��DO#�J�#�
�m����d��rx���IRX�VL��G����#ڰ�7��#m�]��椋s�_jSP�޼�Y��'5���:�u����o(C���vM�+���ޘ-Ğ�z�0�^�n)a�9��V��R��3��{9J����}SY��g�・l�Z=Ec��}���۾�}�ԣ%�~��f�9n_t]AwMY���\�����-�J����h�t^=��\���[��Xw����z�,�y �Y����9��j�؟�<D��$#�K�;-�t��ɣv���ڢ�S8��=�n�;�(T�KL�t�gvYF	vz0{�����U�V�E�*,�,�&=p��#�q�p.��]Xs��4g	wױS��wd����$ѷK7yH��!^mp���v�=VR];X��Ty�w�r�_pw�Ϙ���mn���e�U��J�y�v�mUn��չ��1�8�f�²�P��m�hמb��}���{I����nl�O5�4c�]�k��'5�����TJ��ɭ�����ݛ�L�̋ؽTݕ\7�gK~O,,�ja�b'Z�����:R��C챭��K[款�L^-��SFߗ���#]	B=:��|4���S�uT�Ҍ��3��_t��y�ٶ�1)�Ν���|w~=���;��L���;WßS{��k�1�֤�,��Q�̠ok+СVe:�ָ-��O��s3�S�Ɋ�{�����ȡ�<7�I�u��w�6�����</��rY�'�&[U=�}T݇�]<5��ǉV>���SZC�(��!>�*@�̣��`��^)��5[.�M��cI�ϣn�8h�g��V1�ݍB �*뾵݆�@�=��S�K_8�'�,�|fT�o"�7rڜ��*F�GV����ҩ�'WW]�%�S��`'4��ou��ۡ�V�n>`�����T�@I��x0r�7�tʳմ�R\�bV�R��@����ƃ��:��U�+��293zkҶ@�T��3V;���gn
��S��x��v�E_<�8($�ć�Y3�Gn�k���u�����h�U뎾�-�f���9x�R�g�kg�aY/�uȅ��<ٛ���U��+/;'/m�)s:�ރ=�D�M
���x����6�e)��J�^�27+����bW=W�R�i觘��]W/@ݬ-^�{�-�M=�ӊ���ұ���U��!��C��n�1��i�v��3�t)Y���V���:�;s^��u��Ô���P�ƅ�ʺ]f�n�u3}Kq q��.�{w<�wl7�[[�l腆i�
ڙ�㯲E�*-d43Ӝ�s�N��p�-��s����-����^uG��"�7��Y�ݷ������֗�6j�t�v5��'�{xؔ��yz�ӧ<~�6��O��W���|�A�W^2��c*�������
�}m�a���S�v��	ӧQ�p���QX�n�s�/�#fL���PYb.�kX����O�KU���,�������8ݒF ��z���'�]�����e����w=Y�wP�=\��j�b
@���
+�n�=��/l�^BW�9��qt)�\X6t?}B!*\���O;Xr=�-�f&Wd���C�
�v��n�,���`:nn2*q�_���S���)��%ٚ�з�+f7q+㗖�&�5����vѽb����ݗ@c�99z�s�*u��׷N�t��^X���C�j�ud���2�V͊N�4y�#�㐷��m���ۑ@�Ku�ܛ�ʑN�-x!�V\������A�$�����Miq�\i:�u��Sqص�&6����U�ʚ��=a��&S+	cO�]�	ݍ����H�<�X�W8���z�A��漝 �Vt4p��F����ɓvt��]��Nu�ب�e��/>��.�k�[�X�]�I3E)dJ��o�h�����_L/`����z\��;^�Wk��yN����H�݉a�F)��̅P��PQ2s9$CظV�Fwo�k&<�<3�"'�Y����w(�tw��I-�A��ū�4ˬ�Q֦{u���k	��	yb��:
z���c���`=.�|u�8�E[�D�gFR��kut�*�lM�i`<��a��٩ܳζ��z����uc�O�m?U�<�^�v�v#=��Zm�,|Px��+�Ͻ��>��gǐ�q��ѝq\�^|R�]�K��x��ʇJ��Mm�����7����bӣH��]^���-�G\�g4��B �hU�H�O��v����o:{���2ś��U<�r��ᄌa��eeFNЈ�BP�L�	Ao�>v9Җ��^n���k�ϨV������Oj�Dj�s���&�Xt��'��m]Q�`�(�mC�ݍamc����P��>����*>�.��}�t�^��V(�S5����[��t7�CU�X��{�x�i�Sn�:K�X�MMn����GS���f�7[7�O������x���Syg^l>���T�Ǻ���E��'5���+ΰ
u�u����(�+���;`.N^E<xu+I�Ar7�8؋(�i�e>��#��n�G�od��м����*�s.���㌎wԧX�rqb�Y�7+6,�T���b#��근�O��f�T�Y��v�i�r�YbI�-��SeG��tRa��T��U'NgjW�=��x��dY���V��{x{)�������e������>�v��;��q?l�+�3�z��:%t��U�dU�=�̓��tĕ�S���`����X)#��vu��r�y7s���ζ������v�L<�W��|�B�x��G%���Y��|;ȕumȪ�ůj�Z�K��U��HX��kY�>���6���jC��"-��w3�oM�ޮz��z��j���mkE���>櫲f�*5�&8%��8&�.�$�\���ή�ا{��sA��`oČ���v���1^=����d��,3HN�2�&hbN��u�m�cw���=���*�^j�n�������#]J����5;Aؗ�����u��5}�,���ڊ�c���q%0�ʇ*�F��<�2��^K��;6!����*��ɉ$Z���i��i6���YA�Y^��ŀʦ�ۗ\f|򬬩r���ZҺ[�s���,_Qь3��$b��:�M��5gMt��+l����W�V����V�u�8�o<�*49�A/�7{����(L��T�FL�Ҍ��Y�]�6�Ⱦ���+W������R����Q����r/�s��j�4�=��+�t���e��,�(H(O�Z�ڸ٬��WÙ�4���]�p��N�K���V��/q�Qd�p�%Y����}��H����r�n#0�e�BD�y�����J���%��.��Eg�YrWb���tXw�XQk)i:�ڔ��[rn7�{����x���3e-pj�9+z�|�:�X�ʋ7Wv$�ܤ�UFi��)J9�É[��&h��������݌j�P��r�����
�ǒ��|!u��W ���i�Ee֡2L�p�|�D�_b�YN��n���<�A�)�^;��>;�f��+-���t}�}ܴvr�5]�³h�ػ�WyO%˵+]a�k.ŸG�nhz(Ӌ2F�wv�<��;w���1��7J�n���r�D�*�
t�VaAnn<�¡�q�
�I��@�m�X�ɛN�ϝ�u��m}�¿��Ը�����Y�w݂K�}3^�dB�5�i�֮��iĻ9�Ӛ��L�����[����a��t��X;�9w_�5��Y�NV�᪳�&)���;_Y!��c�2n�ַ��B�L�Χ&���8	I�Ӽ�%5�j���9_E�&��s�zu�J�Z*[6U�}�z����|�<��p!��pSVj��CD�R�NU��
�R���2ޥ*R`�������r�\���ٻ ���#ǝx�mַ{�lՐYL]7��ˬ��D���w�P��BM����+8���|�M}�V&k[������G)>Ȼiߒ;�7�N֕iNB��r����0���R��c:��R�gc�,���Sj����NW{؝t�1�Z��W[X!��sg�*:Ƿ;�wo^ةz�y���[(J��u���2��.n^)|ॼ��zyd�"p\ȻdF6�E.�]���R����FЙ����|WY]6�#/:ѥ��s��2����VNG����.��RLW}���
�fC���q3�mS3�%e+�<��Q�5i�4�Ebĥ�*�Ts]�W7���s���Oi(�������E�.�\f��s��z��"f�V+��7X�J��Vd��*�UtGC�-��o(��J�+yOJ�]JRU���6���v=�y`��g��q`][PMƓ�����Ҡ9dj���W�k+s�N�[2GgB\/�e!��.�;w;y�)�|�U��j�NF�W]����;�4t_F5JXҩ�YڝkF<��[���ct�^+���J��(��Q2���[k���Ieȝnf|4> ���LQ�ŋZZ5�(���5���,F��V*�
��Kj+[k��j��Ԣ33U��lZ�Ue����h�j�h�ETbȥeJ��V\l*�(�Ȫ�Z
��&&D���Tr���"ʭF؃�r˖�Z�+FڱIR��*��PPQeeiR��¤�Z%Db"�!Qr��-Am�+�ڂ��+m�)Z�[j����-+k-���\��m��[l�E�,�FVشD�Q�
������-���R�Xҵ����0LTXcECh�[V[YJ6��+U�m���Z�E��[iR�-b�U�J4�m��[
�E
�ʫ[U��#+F�m�YYQ)lAF�R�\�S�/�bŊ5ظ�m���{;{����5ζu	RVn���Q�N���m,!a���u�r���Yu��A�o�;����c*��1U�!N��kKo/؃�Ob���b�;:Ԕ���f�*�<�ΥF[�yi�nQ�X$�XhSވoz�ڪ��c�9wq+/�]��y��$|tCs�P}Q������K�d�j�^̷7�U�=NQ�[ݲ��a����,�|x��B|+���é�`����i�(�沑P�in��Ld�+]!7D�3ĭ酛�eW�Վ0���w1]�V��'.�*{-�8)�����u���J�Yqn1����\�QEk��F����B�l�ͧ���d��y�\u_;l�n�c_7�)���_�P��3��"y4)���h��J}�N��^�z�y�[���k3��'�qҿvK�g=4;��o�h�A���R"�u�{:��'*ټ�����VVKV3e
ʷCSKZ=�zR�yMv@��J� ���cq��'��	{W4��v� Y<���l�1S�M�$�8-��(��M�#�-nZ���'[�_;�L��׶��]={���hEŎ�>��*A�fWbt��s����J1�l��/Q/%[�Ig.<��݉��g*/zL��ܼk�m���Me�:/(�8)���^42y_�H�1�'"�*���K�3��}�ͪ�����i죫Ad�����t�K��a��)ŵ˭���Pr���}�o����9o�+���F���2�����z~{�h_�ZN��h�}�vm��,��������I�����6����y�.�()���5z14��
+�ͽxx�ʽ������x��i���+y����W5�4��76	@9���7��&��C���<�y}�y=�;�H�s<$�P9Mt�]x�]�����5�xj�DV�ַ�o+��]�gtQ�:�V]c�$r<dB�#�
�]�ӽ�7��k�՝I�o5T�ոY>o]�SU�t�8���"y�2!oMJ�xn�S�ɽ���&�v�Un���No=�m_���u��.C
I�p��:�����-@jS3�ӣ$k��q�\n)Y�ն��p�c��i\�̱J��)�Ule���*h���/�����R��j��bwF��,��M��BwCt�"+��5y�G�l�5Ԗ���˜3����xF�5�u]�K�{��L��7{�G��oc�ԗR�c���_�)�ζvv�C�V՗(W�=��{A�SM�
�뤊��M����e�/Ԫm�{rjyO��W�۪�P{[�	��Xf*���j�ܩ��6�k�	L,��f�}�m������;Z�'�S�An�{�4�So<�v>k/�U�׫Z�opK���ڡ��'Y��S��j��(8��ۆ�a�t�̘��[j���F�H�3�ؓu�:�����o��߫Fs�̖�5�ލܽԯ��C*�N�ִ^I�޽�%���z���ݙ���0c|��]�.��&?c�Vj��|�vK�[O���}���ګ�dn'�I�.�[�b7�:x���c/�Gj�+�gDֹ��>ٞ���+�u�P=��d���L��H�G'�`��gC9�k��X����6�Չ[�.�<x�a�ZC�=I�V�OP�c�2O����O�X��:���~��}���k#+�v��_�i�ŀ��Q�������l�/��E�e�{�h�����i�}B���Z�5+\��-q��b��`�+�:ّ�@�|��bSw*--+�]Q�gt*n9܏Γ�j3bJ���`����RF��1rW`����)�e�/2#��^L��T?}������7�aԟ<a=�XN'��y��%I=g��IX|�{N�Y>Aa����z�����>a�m�{��ߡO���Rwz>���+���yl{��^`x��N�!��2������&2o]�<~d��I��O�L�Oy�D�'Pߝޤ�(O��VO�XyhI�<��.%��F��mv���������6t���O�[����Y߰8�Ğ?0�9�<`u��<I�OP5�'SL�0�|o�	�6�}���:��}��1 �=��Ȫ���"/髿�B;#�G��w(I�OSf�OY�t:�I��7a�J��k�rq�=~a��a�����2u�l<@�9ܓ��OPY�]���#ׂܛ�jHuy�;�τo��y!���ڒ�I4v�%I�+&�����|�٫	�S_�x��7C�+�!�=���6{�?$�I��^a�N>@��l�X��}��te��>� Y���x��kz6�:��^y�*T�G��+'߬
����u��N0>M�|a8��AzɈy���I�Xf~���$�����Ws��3��	�a���#�9��>A`o��T8��7�a
��M��d�a��d���;��E������'�?>'�P�`u4n��~I��#l����2���Fg}؏��G����q�c*�u�T���'X��ĜI�*��!Rxɩ�h�	�M��$��I���)?>04[�:�a��LjK�:��X�wg�7��}�>�|��&�q'�Ɍ�A}<�	<C�n}�Ad���u��M��<IĞ������zɾ��_$�@���%0�O�{z����޿o�;�k�)=|`v�z�|�3|���Bkt�d�����4��g��O�q��'Sl��~9�d�T&���Ĝd��O�`z��!�:}s�qKYE�ˈh@��������ns"�MaXq�Q���#YM!��|�n609/B��v�����P#d^��֝㲤m5s�e4�q���e�|�Uu1Έ�*�c7�]�gkǋБ�:b���l�+H-���ZV�"�f�ڽ�ή��F}g����$N8�|�?XO�̛M�gY'�Y�:��O&��i��,��d��uߛ��$�e�M2O����u���'>����$%�=�s�a��X��a��@�ò|{Ԟ���4I�g��z�M�񟲄�4���Y�I�*kt8��5��q�ъG�d{��#\�G�>�\�b�#:�(�_I|���Y�y�d#�3�'�ì�I��'wd��<~���IY<`nr�̬�a��!�i����2OP�bAd��2u+9��.�������y���)=I�*t�̐��a��ï�'X~�d�N>0��:d�x����I����oRT�Hl-YY=a�2��d�T���8���g�
�[z��?V�}����ޣ���ޥ`h��I�N�C�y̐Y8�|�_XLI��ru'�O�ޙ$��ɳ���+$�7�oRT�Hn��+'�,7�����|��:{y������{��	�'����ެ>M2O��Y>v�x_�8��N�C�{�'Xh�s��75�:���$����'l�����Y'����z�w[uϻq}p�D���@$Q�� �|�áh$�'�م$�'SF�>M0�f̡�'_̆��d�O��3�C���s���O4��}�u�d��Q6D��&�~����;��yϽ��I�<����5���䬚�z��l��q������q�݇�<|d7}Ì���3�C����x�f����~��~}�#Ȁ3�yi��{�`N��K�`,��xw��%J�h��aY>Jɬ�q'��j�5a8��h�aְ�C[��%|d?s^����?wn���*���{�l�}��|8�ӿ�a�O�x���T1��=��HuY;��XN�y���I=��0����6e����wTެ'>f�W~��ߝA�JQy髡��V�1�2����9��{B��1��q�q'Z��Oeq��2��ǖ@��6T�4{&�ۘ��dޏ滙���AVe�p�N�m
�ٴ��R.���OZ���QTO��� *����ɩ>ް��.�ȝ6�oP˜�j��|G�}�!�}aԕ�&�o���$Ĭ5��q�Y'?=ɤ�AHn�B��'�,��p�I�MNw���N���5%J�u��<O���й"g+(��w�}�}�~����&���T'P:��o���>C��u�Hzy�u�bV�{�Y&?rΤ�
Cӽ�T8��V���<ICﲽg��}�#l���
�.)^/�J�\��I���E'�2ì$����P�d3T�:ɴ�a�}`x�2u��u��
�}�PY&&�y�Y>J�l}���{����>������~H���f�_�����HT�d���ԓ9�%v�|��)6�`v��$���q��t�4�ԜI�'�c'k	6�Xp��> �� E�_l|g�'�go�5�����VC~P���O}���'��;��nI�O7I�'S�E&��4ϲ�2O���:Ì&���i'P6~�x@��̀uo-��f��8����,���#ȇC����I<C�߰�'�;�d�'��<9� z��O_�;�=@�t��ɦN��d<g��M�d�%MM�qG����:��Ffb��_!U�淟Y�=A@��2OP�'R�����I�7�a�m���fd�����P:��ԞN��:��'�5�$���8��I<f������5�*+��oiee���{V|��RN��!�'R�6~���'�g�`N$��w�$���:�����L��ORw�N�O��淩+}���V�&��ӵ�|��4�>�q�2����>M̦$���7�Aa>u�2|�����E�Y8����d���4o�;�u��fI�ē��L�d{O���;;���|�I�� {�+$�t���Jì��C��>Aa��!�'SfSO�q1�O�Ì�%`|~���d��{ܐY:�F��8W�X����y�.���R���ue5��4��"�5[kk��[G��G�-�}�(��-��N�@v�"���}}}j#`�*0�Ṡ���G�'cNs�F���c��t�Vf��s��A{��OB��5�w�=�
��^u2"~��\��+���ND���W��{�|��p*���#�x����Č�{�|ɿ{�P����y��J�����B��&�`|���M�d�$�m��'P�'��_�8�ğ>!�=�l�8�O���:�6����i�|>��ȓo\�:�d��O��'��'9��a:��wz���5>��VO��k(`��".D{�D{�*��D{�g�;�.��v��w1%_ ϼΑ�T{��d{ w;�<I>���&�~@��rN&�=I��`N��M��z$��|ԕ	���J��VMe�=d�Ӿ�ϳ��w�1Ј���YkV|=�>�#���{����J��k�ru�Ԟ�!�s�:�9�{��8�����:ͤ�����:���3��,'Rn�z%ea9�|�g���������f��Ǽ��䕓Ԭ���'Y>t�����z����I�<�C�+�&�l��a1�Cg����Y'?G�i��)��!P�'�,�{�:���]�����A]�M��Uq��4���=�������rE���������oVC�SG�|I8��X���a���ēP������M�m��)���}�./���]�T� ���dA�}�
��O��4�:��y�_�I݇�"���Ya��?>'�Y2j���m�~���4�����	�u����|~�%EE�oOs�%��z�\�>� �7�d�'=J���0�a�&���z�1�g߲K��8��I��Ì���>P�N0����'Xq&�뾜�~�[�lr��E�>Dy	��O���~è,'���ru'Y�̞$��Ԭ?w����o�~�̓L����N'��|d�y2Ì'��r�{�QF;�s^U}�fSU�z��g�χ���d��g��u']��$��n{�:�d���=�Ԝed6w�:��O_Rxs���7����'�ǿ����u/��yb��N<gk��4�������ePwX@y��x4�Z���ݖ��c
��8�s�KN���V�����֯ ��u1�o�k\�;�8?����W����E�s�wu%׽L�p��pK�u������\�B�5�:�ǧ	IY�3�=y'������=��_k��d1<d�?���$��6��a5�d�'���q��S�XO�q���É�I�?���N{a?w�:��O�Q��'���#�~�ޣ���ne�F}��`m'�d�����=grΰ�!SF�:��f���'PP6~� ��'����a��u��q�y�u��X{�Q~봾�K��}��R	>��,�߾��q��O_�[�T�H,>J���|e��I�o.2OP�oVAa>vÉ:���?}�Rq��Ss�2Ad�������=��'nl����>���﹇�:���@�Oό���I���w_�%aԆ��Y>A`�>CԜek$�'ڰ�i�|�I�+��aދL[���cf�f>|�e�>��{3�Y�vo�|��c&���ԟ<a?{�XN'���J�z��9�IX|�)�+'�,<���z�ԣ$��|>����O��ر�=f�9�ָ|#��?5�̞��v���N�u�'���:������75���O�4���4�����V�o��RT'��+'��)����X�UOq���g�G��̈&�x�!�Y'�v�w�!����N$����s x���p��Oz����u6��'��'��M����:���\��j��tֿz��>#�G�ʓY@�'��&����[�ֲN&�a�J��h�ܜ@�O_�y���'�'�,�&�~@��rN��=Af���T���vq���|��w��~�@d{�O��,��7;�ڒ�I4^$�>ed�:��'Ο5a8��k��|�St:��2=���=�6��'��Uu)gՔ�~Su����a�D��O�i��l�0'P��}��m�u���5%J�j{x��}���Rq��N�q	������N0��Azɤ<�8������h����p�jrD^a�O�ӹ�nT9oC�n���9[~w�^��%�&6	;#mf:�f�Fs���6ǲ	�nP�^�+E��Y7/v�T������휖ֹEA����vu+v�C�ձ�q�n�*ӆd=Iu7Z���*&��{�Bڽjq���?�}�I|+`a�I���m��,��
�<Af��!Rxɮw���N���2J�d��Ȳ}��)8��Oω��	�R��߼���k�[�y5{iW�Ady��#�H�'ߞ�̓Pןa�IS_s�q������<eC��*O̜￴m��'۲Wl��CܑI���o�鿡��fڹ���o��H�}�Ͻ��4n�3�M��Oǖ��N ��}��!�7��u�bs�u��ON�'�8��T?�@���M����$���Gw�oW_����=�|�+���=�)?<`j[����I�'����'Xu'��'�i��.��~C�o�d�m�z��=ì�J���<I�O}��{���yi�L>?S��y�{�o�_q�ل��������ɴٖq�x����ԜBm�d�&�?!�N��y�ȏ2��2,������S�~9���;O���qv�a������}�}�����z���>�$�����=q&�xʄ�1���Y�I�*kt8��3^�u�� �{<����CϾ��֚w�_Po��r�?�#��|6�q|=��>�8���	��ì�I��'wd��<~���IY<`q�Y1��+!�1��R�O�|j�Y&���5�����}�����p8��VOy�Ru'YSs�d�d�O��_�N��̝I����@�'����ܓ�'S}��%IԂ�A���af<�
>�#�1:N�g��k�ټ�_��t�x�m1�|�(|�Ԭ~���'<���d����:��bOO���>x�~��I?>2y��+$��׽y���q�;_E��V��x=�!Y>Aa�`m�q72��u'f�>M2O��Y>v�y�8��(y�rAd����$�ɳ]é=(�i��}#�dY��R����;�+`�J�b`�i���f4ј
�yJ��}�B��O��Q�.��i���ۃ2��9�}�on��&)ƻKY�,:][JEMM�Gq^�s��tv�䬰9���u�\"�&0ӽ��󥻼���n콜�98Fd�
o���Y�xb���V�a��xA���ە#�@$l�
���Ğ��7�$�'F�>M0�f򇬝2�8�ğ���9�<@�v���&�<?k�gt{��.���|�<�8~�1�2q����$�m�p�hI�7�h�	����䬚�P8�ԟ2�':�n�検f��=I�� �N0:�����X�)��x7-?����vO�����T�>���@�w�'Y�OXi�o��m�y��I�7��ԕ+	����䬚�z����V�����k	�3����3�-�w�;k�&�J��dz>��[���<z��a�I��0�'�<@�;܅CL� ���C�O{���o$�RO^0��;@�e����wT��yv�1y]|�\,{�>��y�|z��q��>I_Rm���g̓��{�a�I��ܚI���܅C�OY���'�4��M��I���RT�'_�8���9���/~FR���<O��H�N2u'���5B|��m�|d�'P����d����$Ĭ5��q�c��2u'R�r2x����T�#�e6ok�"OnOnW}f�	��>��^��I����?�52ì������!��:ɤ�a����4��6y�u��
���I���u�䬆�W�uL\���Ǫ�O��y���D*O5�?{�&2o��%0�O��|`xZd�z���l8�m<Ld�N$����d���M���G��纺ت�����Ob��k�w}���wW�j�g�[R�=aS�;=N 4m�i��n'���p��n]e�M���q^��y����|o��=_E���ML]}�q��{ҳHj�ѷPL��.^�T-���Z�޾��t�LcƧS�b�aM|�dL��kF�����c_g)jJ݉��f�������a�[�,���x�h΅����41�`9�V�x�dtuD']�K:���ɻ�On:l��$K�&����p!M���\2V�v�Z��Y�f�R�s����P�B�z7���|Gs;�J�PG�:iw
�G+\�L]/��Ԡnu�N[�i�u��K���V;��g��3�I�8��2�*����W*]_Ҿ�����]lڴ�̇9e��q��{���\3�����R��
�fnVc��o)2R�9__:�h'S0,Г�U®Pc]��E��^�>d7��k�U�J:�3���E
*���o��Ww��a[s���v��)�a��hT�j^Քo�M�{����q�4ns�0J31q��O�ʘ�e��8K�.�J�W�7C]��X�sFDs�w��ؘIj���M�HH�]���W6o���1޷׼y�}h�
��
�����p��6ѫ�j��TRb��es�T��U�Fu�|�d���/'L�1�ɗ��;D�(5Ԭ�*Q�]�iF�%����V��;��Ukrk����u�R���n�̼��e����k�Q�6�ʱ�6���C�=��A*��b��)K�D8ia���h��U��D(�+Ù*�8��:��r���f�[�lt�6o1�Z&ƴu�{�C�w�Z�AT��GnǸfQ��{]�}(JK;�\q���A�ٷY��!�oc�Ń���H(d��x���λ�٨M��U�ޑ�֏�e�}�FR��
��^�]�⠁��Vlclާ�֕k�4�U]��Ͳ�Kr�#�0�S��t�v���kޮ��U�v��d���4����;B�S,���N���������kلv3��A�j9DP�Z
�of�ҀOgY�v����k�e�zT�T�>��B�R��viKq���ʦlJ]��Tuu�fe֭�ʙM�:"�P�n��El�6�,��m,Ǌ9yz���b�����J�L�3�Fb����C=��q� E��̹�)�K���vV�ǜ���� ��^�p���պ��5��]���&Zz$���1;M�0�t��NGt�S��3-^�hW,�7��Uu>2��X��V�P��ِ(�c$�'�Y�k*��'Vg��2��Hng:9
H��{pkd�ZtDt7�)���^9
�դ�;=c�vp0�;+E��2	���n���OE�gW};ҋ�@��������I
�w�ì�DN��)�iR����c�Zn�|�ⱬl�r�K��9��7-)��s�]Gy�!ؔfnrH�����Ι�Ē��QD��[���;1��mp�隳�\��Ω:��ɜSJ��u�2��u�y�>��Xt�85��P�Y]Μ��9�Idƥ�;@iz�7mg4��R�z��"�3E���T�X([KRֲ"�(�[VZҡQJ*Al�Tl�֪,�jְ֨��0m��)[[+в��J�dD�`��E�Kl�J�J�6��lm�T(ڕ`�Q*�9�
�i+[j5�c�čE�J�[`���+h�D*U�����Z��i�c�m+j��-d��\��)FQ��U��ԪT�Z�R�QJR�V(��e�h��Ŭ*����-�Z�
�R�5�֕�E���%E#l�FV�J���JY,�����L�L��DX�KE"�ڬF[am֦7,��m�-D���&&-J����FV����j�m�)Kڱ-�Z�J5�Z��[*Z(#E�PZ���iV��֠�[iKUZ��--�,DYQh5(��kb*Ɩ�TQ�_��n��j�	���e�W�t�kQ��۝8ZZ�'z�Y��d=}}�fFxB�g��/��F�\�N#{@�ڗ�������]]cޤ?=�/�3ci:R���}����t�;ʯ+�#90���޾��մ��,R'[7�#޴�)|ў�f�,��NKHM�j���	��6V����O�q�|���O]�����tn�S��p�ݾ�W���vΰ��<$�B#�z\�\o�y�8r�Mf�5=Z��/�`3p�u,����<���>=��ޠW��v2�q��z��v�5L��z�P��*[W7Oiv5�8@����%����l�Ԟ^���N�ϲ����B�Z��SU�t�S�
��$g�,��U �@�쵘�V��Z��nE����$f��U4�r��n�X&BF��)�9y�l��������-SB^��ugj��@r���7͞�x�ݷ���μ���q=�����])�LWJ��`]�y�w��*��6�!P��z��u��b�����=�b��uuɒ���V�*v��S�|8�ˎpm�]7�!l�Ɉ��j���ʆ��}c�"���aLK��|��G�Έ��']���1�MkγF�ŔxS�}�Ǎ>��cs���8��e�W��w&W��x{��bj�K��c��Xh$r}ޏҺ���ب�ˋ�%�ҫ-y�L{�`ВF�Ξ��m�����!��ݬ:���{�mW���N��Ҫ19�ъ�@u��ۯ�6��k��.��е�O3�ߛݧ��Yy
�^TЭ�][#��2Z���:�ӣ������c��js���A�{��v����V��4D������m@arc����N��WϽ���h]��޹�t��a]���<��j���*�q�.u�|<1&��T��U��f�Ӗ���.�?n���;}�YU�ǲ�d���v
Lϯ�Gc�r�����^��m�v�8|�Y��qE�;�ļ"5C���+Z5�����֞��թZ�}ifpN�lP��X���gkب�g��,�hr&3sz��=ܰRc�Q�X$�^5�}��g]X���}f<��>C;�R!�;d>�iP��H� Л�ɻ�}�y(�I���1�/1-g�|+(���-��ja
�r� �7M jn�����`�)�s�x�[�4M�y��v�e�t�*���<��bќ�W�7����m!�e.��"]�\J�u=�Z`��lڜ��x{�����qw��G/���Z�%��4�^u7[7O�=�Lm���f\�>z�::}�dPǍ ��C��<;J�y=3S���W�A#%�Q�m.����f��[�����N�d���e���n�v���=���`\�����3����0���]Z�t��I7*�6kg���'ڈ�~�Pe�漝!A��W1��6�\�^#Q�7S]L���y)�����+7��s�C~���Op��?�	�?J��	ɟB�5�k;eTB�����#����`gd}�D����i��a�;��u�˴ۖ�⃕��W���=���[̈́;�V�S����� �Ȓr���S���H���=����{�/wq��4��x^H8er�r����9���U�J�.[a�}�����mmlV\d��Ȥ N���}@{�^R�4c5�X�z�b&�O�Q�f}�t#M�e�V��$���
��bɢ��t���kwi"�]�*�������l����VΌ�Z�b��S�S��u%nR��|��[}F7�
eΛ�g.Mw�F+!D�j`�
����3h��/��� �MV�:�Z07޾�N];��}����v�l*���Y�Z=���õ��ى]W�i���{�o�f�lo�-_�vm��q%�:2��T!{H���ۙEo�v���ֹs/����^ �R{��b��n����i����-��;�p	�r����zfl�sy)7�����Y}�/�gq`�̣�b�'��%k��WJ���{�GOEi�f�av&e�A�~�ղ��1w,V�st���:�dO�2'0�z��i,�o�l`ٗͩ��e�b:-���f�'E�Xݓ>�xȄ�u�z�Y�d�0r��\Nc}Ǆ|#��>����3��z\�����&�$8�9N�om�)�R����:�٫pxo6��B�g�6o N�8���2���
v���f[=�<Fu��r^��pgõ�ɡM���wE5�.�����Ww�,H�G�}k������,
��n��(�,t��#��y][Q��ߟ���#o+9��f��	�>Ft��S�}o��!5�]��r�bV6�ݭS�i�t�U�)S	t�Y+3����C��>�_7��R'Z[��W�������f�{T0J����z5㥶gjھ5k��Q_����T$5�YX�MťUͶ�&Z�5e���6���b�Y�^�y%S�e*�kFl���A4�#�+3Y��,�U���#A�v�{��\���Զ�XO��s�\�<���ur��R�\XЬ�]o94i�{��'�O��Ҟ+ꙐR���ɓ�w<MfbR��9�_ke��K�}��m��y�j��/+d�܀�v�B�T�r4��q�Ȧ"u3W�#i>
_;P�_���򅲟�n:/1�JgP�
��r�ˡ���.7��ш)���Ʒv]�z�����ݼx�Շ�7E���A�Uʄ����Oc��{��7O�s���0��f���[ٞL��G���U��G�5:�_e�ff�k�S4K�o;��R�`��j�o�w��st��%e�3�� BމGi��ɰn��t����������������ۯSkr����Q8���Uy$����
ّ�X�q�1�K��٬ 6ı	�m�C��(!aK���}�
�z+8^u&:̛y��S�6��7Y�gFz����6�ʰjo��}/m�o�U|< ���[�ctw��~� ��8��Z�2����S�	�"�v�Wn\�z�m�RZ�(����~�ٶT�����Tҡ������~��pN)΍���r�N�ha�3��M.�N��o9�:��r���B��˼����K:2�!x���vV�p�!nM	�7X����� K�]�LU}�켞~2r@n^�u�pXh�HN���n�uϡu�ʉ�Hmښ���Ԟ���،�Wn5�ec�M��a���c:ͮ�
w�n�M��������/g�5Z�1N,�B���s^Z�yq���zl�Z�,7�+��;fA5�}.��1��ଖ/2�V�[~Zѡ2M��׻��Jj=�����N�Fr�����{ͅ0�rS��b�м}�>�������]ʠa1Z�.yhJ�1j��ݰ��i��Eˡ����:د_�bO�w{�H�g��#�N�l���V�hz�bV�/�EL�����o���d[�:�9DFb�K�e��!{R�
T"�>,:�,�䳕������a��"���1$k�:���8IS{`����o;Lr��j�y��)6mw;�r*�-N%޽�b�
����������jJ�w}��/�R��o��YC�^FJ�"5ׄ��I�!'(�{R��=oi���)�o��|�Y��$�t<x�ڨDj�$0�u�;�n:�o�\-2=z���>��o��amc����0a�X���۷���rf]�^����`�y��վQB^uͷժ����ӬOV�
,'y�3���+Hu�	��@�>�*���go��,�nr\EZN��f$)��\�7{��ex�����s(�<���c
�>�j��҇W����\����5}{Ӂ�O���o��}���URƿ~�3S.eo>Q=�Ҵ�bUU�o]��Ym�����ea:�QX瀕Ԛ��2�=�����n�rW?pٚ���9Nx&��\�P��=e��.H��ڗ��q���e�Vv�c���-�VZ��Y�� dM��=�w�4&6k��wAgZ8浛;3x���O8�=25�љ/w;lժJ�}���a�P�N֖���w���;f�6��Ы��E��%l�׼�_L������"1�����p�5ֵǝݥK���nV�*q�^.[�ި㝱��z�I�Է.z3s������ZM��gJ���-^\ҟV:V3%
����X��kaLT���0��d����ɇ���6����׶���o6JY����e��d�v�y��ukQ��'�"t��nKG��r�}YZ��$,�"�)����ZՖg�2m�Km�}��{<�S�q|�!y�"�Z5�f067�)^kyKF�H�Iה�v:e����OfJ��ЬY����mc^��wFڊx��4kփ�o�-_c�l7#��'z�K�紫��f���@����z��=^���5v�B�دs|�����m`oz��]�x.n3<xP=��L�pzb��S�z����ca�Kd��}���uZ��c�$r<$�drY/��n	ܦ�)��hʼ�v����t�k�k&�5sb�U7a�0r<J�� '"��C)���A�DS����F�c���K�T��}{ʊg;i���]�5�u��u�K��(��1�˳t�
竕���3}$B�H�Z�p)�<�Vҽs��G���^P���b��S|���gA�����R=���P�S�fq�W,�[[��n>�Ғ�(�=�s�}�=�	���f�15Ig�s�]����!cvO3�=z|d��Tk���f���YS�Zrs^+�O����5��$��F�:����]�j�(��nf�c����u������y�e�=��9� j�}�j�F�I��s	T�[y~�r*���1�{5�����T�1<�{����I}!�����Hj�k�f֌��w����}��9����7���79)�u`؇�x�k�rq��Q����R�)O�%�P
}OgVܬ|�6��F{�������֋����T��c�4p�l/a�����VD�׳{;�ޕLwN
��������>)�{�;[{�y7�ߎƻ�K�g����{
~��g��u�]��6�P��e���t�'<���J7�@��K�O�S��hih�����L����)|�CY��n���U�]��J����ح!�tVU7
���K�O�Y�K2��8���>nS�1�"��R�cB◿]���j���ҟ^G0si�ǽ���N�s)pw����ιsg"�XO��.��א�������p�� �<��f|�;�]��]K>������y�m�"�}ܲ��CN�B�^��^�:����AA��׶�H���؎��éZxƼ=M��o�K��J�ǅL�t�a���j}��VZcXsOz*[��	�ծ�V:#�ᇵ�WJy#�R$Jy�O�����/d����ٞծ�o�W��s/e*-�<�<��:�c��*!v�*����&��ϫ^j��^��5[&�J]ŇV(*�6}�]�Q��9Ɣ.���g�K��G9�~��T&��ꇽ0�YK��3���u+�e�uK�w5䬛�>�DbY��A�䜹��e����F�@;SB�T�b�)�C^�q�����+~}tS�^�GoѶD6��'ַ�^��o����i+=�[����H���+�����6|ׁr��s�jZfF��6Ӥxm⺦xM�k�}<���]�׽�9�>�/bs)��ue���@�p�F�����םrEE`�7c�fw�Y��᭘S����kf3�p����H|�,osW|�z8�l�ꀟ�
�e	��q]�'M!t�����G��s��,_&�}G[�Gu)c-̠�����ӭ�#sz�(m��E@��7���Ǝܖ.�G�9�;q�zU�f��ɗ@NX�s�h4�؝I�49W=�]��0�b�)ks�X���un�Ԩ)�����fBM����wʹ���KdL��i�����y81����X�d]�F�����ټ�&�u&�4&
���QF�S��r�wwwY-6t��޻�9�\�;S�f��sR,�w�A����7{���p����m!���M����V�����æ�U�'m��|�tZ�k���]%W�nm7���Ւ6��[�K���je	Z�\��<�Kv�%N_=�Gn[�k)��Ƿ�A�>�n�TZ ���7�:�w�3�N4Wk}oV5��t:4Aب9g8���h�ԑ)	,����4�uo^����x�p���F����H�$205�s�@��Y�c��˙9���8y���b}�_@,M��93:J�NVK��0����Z8�u��"Ts)��I��Yʵ%P�	v�<�n��nEr�v���rnҎ�C�1)����Z�\�Ԕ���i��澚a�Mhw�n֦���4��\���'lh�g������!��*�Z�tY�dv"�M�E�N�wUغi�;�6%3�ؗL�Vg\��;��.l&�Fdy[G;:��m	Q�Zb���)�Fh�ў5��̘*vlr�LsWW�ڣ{�e��ңW�IO��C�����(�N*J��X%��Ų*{ݔ�n)�a���L�YɧR}�Վ�`��YBaU���Y�b�7ڶ���M�؇	�4�֑��i�TzּIgh�Q�[)4�X�T�Z�;��}�:Λ�կ�el����q/� �oPJ3O��uF����B0���D��H�>�}�����IoX|�k�U�����<��pr×c��3EK]��A�W���S��;�Mt��f�*C,[MV�;<(�W�X��D\�T�]rݬ+��c�[��uԷ�2Шi�y_-7)�SxX�/kx;o*�xfԛ����յ}�u9X)�s.���6���P�nU���*�,6Iι�S�d�3���s�Y˝�k�Àf)ϐ�,�Զ�����1��j�+{�f-�Ӓ!C2E�x�kz��۩;>X,q=�ڍp��2n�Q�n:M��H|2��Ϥ�v�Q��1c���}��	�L��P��&����Z:f�X��*.��¢;�U��4��k���d�u��©�S)`��϶�����iqa��f����� ��*�k�ךQ�{Ht���d�ڔ�Bn�D8�]"p�gJ���˙�aN�A9�:Dr���6��8�2w�0x�u��h�z�o��uF�弰�N�ھ�-��w`ǣN��Z9����5d�$��̎���sjI��ʉ�G�h B����Ѩ�V�Zд��.%�*#��5���VRՔĘe�*��QAb�V�(�mmaP���,�U��**�De���4j�Zѵmhђ�R+FU
ڬ,R�U��"Q�m�J(��lTYme��UDch�̸ �˖�J6����V�D���R��lEE1
Ѷ(����b��edX���D�T��Y*Ti[e�j��*�#DJ�h��UB�(�KKD��˘��iQ�UF�X�+Km�jU"�i���m�1jR%F�TUEHѕA����PQ�X��"�U��"�J��Qb��k
�bZQUQ����+*�Z�X�T��QcFѤE����K*(�����*��0G�X�e�Q�*��H��
#LKh5�@JԴ��̱Q��h��m�E%B�V�Vڶ�֠�(�h�imeV�J#"�m���J��U!U�B�ѨR"����i+��AĪ�[[J���b�X�P��̸��j�F���73:��Y��nƠ��ۘ���,��w;�Vt�YS�ˮu����+���s�X%�19BvW3ĕP��;�5��{�xx%H[m���S��sƯj�{0��t��P�Z�D\��.K>3V��͞�o�\ݨ��^�����i�5SZ.V6\|&�eZ�"66�Ҩ���s��%�+sx�o&���d^��|e��{�����q�FD����$�t�N"��"�S�;%>�f�eWm��`��<ާ�:�Y��a�Ub�Kz�$<�[�"�U.]*z^���K�"����qˡ�ꕑ��)���27�;~�ڇs8���Ym�dT	��.jr�b!n.x��1�K�3��iC�eC�P��>ͱ�1q�f�
aA���b�]͢�����_d\�K��;6;�!\�,�/��8{5�qmuI���$"(c�Cn�n�S����楤�f��͘3�qx4t@U���`_�>�T:�.�'��,�uo�	�u�2�<�uAJuD����돞��:n]�X���_�Wr%B�D:��^�T�:�hC�8t��cj�7��V�<����ԭX��%�V��u��֢P�l�˞���)���^��D9jb�퓋����t�����Xy9�u%�}�\q����*����t��^��z�u'?���r��{D��ԧx���+��ӽ�[��j:o���wf���r�D8aЇG�g�[x xw'w��]���Sb�oh���w6M��{���ᕘ˹ݓ�N|�q�N+`�:go�� ����'�}�\�봻��(1S���B1wܞ��|�t(bܣ&�M�����>��:,:㻳 ����4��hL�{��K}㭆�Q��E0:�¼���bb(��4�����:\V�>��H�:�$s1j�O��;���A�W����z�3���7����@�z1�XVyjX'��r�&���ԚǝZ�V��g�yxY��\�1�;^��Y\F��=�^s� )�V%>9���Lŋ��Ir�˶�i�(�oQL����9��O�r�1ՍAˬ?l�"���*n���͡����=��*z��U�\�Qiu�V�������R���5�uۊ�X��{��gb"z8UN�~uN�NyC+U�68F��[Ӻ���7���Զ��v"f��W"�v�v�ǽH`~}#A�}%C�D';�pt�[�Y�ǖ϶�h�6�Y������������NXѾI.9�4ꄗ}D��g���N�/�?j��j�P��)�Uc��{5{]*�v��i��`k�JE�8�x%����__g=���72�Tx|�6�hPa}����n��E˗.S')�ܹΫb�9c�D�������3-9�u��{{t�Π��YNij��2�by3��en�@B��..�6Y���������GPh�1�FD,�Q'�bx��:��L�hbF(%R{bJ)ˢ��Or�Qw�$�'9�k>�M��1�%2<_�(��]�"��C�5�`S��`Bt����%�C����N�g(L��4gϺL�z��[.�썠G���S
�>��x�R�X��-�[�5�鮵�f�M�Z|�+�=m�Ȭ�H��C�%�vd��0I���@��L����������=yx���V>���<��[��eȫ�������7.�1��	U=f#����ڪ��s��/:�B�d2�֍�sѳC`#�,J�c�����X$�5w��p�����P.'�{��No'��GY�.Z)�F�B��͜�3��e�e� o����XX�e�v�.[�[�y�Ё�P���!2�^>�(��@߈��yu�1��ltS޲hT�<vT��ʏ� � �2�4�9M�X����
�	܊��w~h��P�>��hK�r�*s{Ȳ��j��Ra�C�;�{����{V7��c���(�ͫp0yu�E��#N94!(d�R�0�7	��$^�F!���F�oSG�x�e=���^��)�y[�(kj!����nԱ9j�9�5�<�Ɨ:�%Ԯb!j��[G���3��0J��1���n�ø'U��[yj×���X�kU����_W��
�����oS�Hq�8چ/.�(��iZ�D<�㺀t8񦧌�yR]���7���Ʀ�M5.Jݻjq�k%ڨ��H��lw��r�n輓�dpH]r�_"���B�=գ�{}=DXI�ʯ��iNQ5�DfV�Ix돬u*��r�)F��ޫ�uU�+����p/Sլ}�2����t��M�)D^*�[AP �egb���/e�*���!�xNlQ|��4��D)�BbF���DR� ��sͲ�����9��`�;>�cǌS���
��t�G�
4�,.5����<�H��n68�ꆆb��۸�����:�ܔY{���h[�re�޹�̣��.
7��@'0���썵<ŵ<�b���Z�F�t����8�����yt�c@��;U'��"���ۄ��<5�@(M<%�7�z�TUc|J����6_E�P�|hF�̦�5eua|��q*�'�)K���.�N�ޚ�K'b�d�����$q.�pv]�GJ��	A��NJ�eg��gG]�f�tLLӡ}Y�7`'��c;��үC��v+]��ƥ�Bo*F�FZ�@P��yY��ר�+=Ʊڣa�YR^S�X�ɧt��Cy��6�2Wa���UNU��rI���W��NЭ���f-�k�e<���pup�MВ>Rj�躉�@��o�U}����^�Z7��n3���B�A�S+8-%�Z<�~e��hcN��C�r-����U�����r@#�jdU{�{Q�Br��X^�X�»��Z�6�5��ː�m�Y�_�t�ͮ}���_�b��r&lƼ�{�掵-2ͅ�:�=�^�G�ep�s4�R(ڛp�
������������%��(ז�@�y�[WM{^uɳdY\���u��wuݮeE��f8���U�.��fmkP�V���cll�%M��e��T=4�7s�;;B�+;��\���i].V=*�>b|D�X=�'���uDm��р��u��VZ|�-s.�a�Ƚ-���5nςU�<)�8�}4P7��N"��"�>):���VW:�jѶ5P[��O�]�;�;�_X�RƁ���#Elp+Qw��7k
�jT=紌Ӱ��U:���.��VF��]�� �p���3����~�W�Ij��\J�\䮩W�����ƌVJ4>�lyK�Q�X�f޻�/������%*�^�k�z8���j*�`�7�^�}S��~=Q���!�=����.��p�7�g+����4��F��.Ƚ���%�2���ch��u:6(��B	��l�5.yϒ�=�/��QND�������v�̛��;�"R��ϐ�yS����5�ƶ'q��U7�����߀ {�W��¦�3l|&eu2B�|c��f�.-��(���D�e����!s�v�(�\�K��d,��#��<7��G����D�a�w�y�{};j�{��U�;-�Z��`#��#o�@��%���\|��U�tTGy������A����smuKZ��)V6t��wưZ�q~j�%Ϻ����B�z�J����^�6�������o5T�z��
��eKZpȞ�a��.�񸬒(t��#5s�ǹgKG(zٱ�d^5��Q^�T$��6�pS+#�ٚ:/��;N�쳂��E�ט�O=z�\Օ�ٷؤɵR�P˯e펱�\Uz�ؔ���F��`�z2t���d�igM��*����m�;�vh��R���YJ�t��Oя��_&��W�e˥�A;������_\�z�ڀ�.�/���Nס�x�8���!��Ohç��s<+u��KݒC�]�������ʌ�P7�T�ōOɂ2���ͦ|6�+Ƥ�:���Q�+�{sQ�3�뽉�Azi�t���r��hL�}��[DO��D`�@v�&S�d.�����qv�5Yhg�=��Q~1��]rE����Q᪔�����;��<��8c�&� ,��Ek��/*N�����vf�S�tr�詪_x{��r�שz����2p��+�a��݌�_<X8�tHh�Qp�lh���3����^b|2����Y��1����T�4�VŇ����H���A2��]�>|{}�{)��y�33�R9�	+d0h_Ip��%�W���:����w�e����vv�QM�c�G����o0�;�>3���t�M_I)�R\Qo�;
-�Ġ��-�u�-�D�7{ �~�s(x�'I�2����)��Ғ�/��B�u�ٽ��ۻ��l+����N'ڼO��3{� ���oac��S#ŀ�K�'��Ou*���Y	�#'ʙ����u���>D0'��o�w�&5�eTW��A����QDp$���D�Uu��4���u֤%��t�bj�vC���\��'�2�[t�+-�7p�	g�' �0I������ڴ�n�fp<��򝆇_V�к8w�zG�Aھ��Z�_�6KH��M�Q�;�}���w�E~\�VF�di���[O�x�W^�c�60ܔ��%	�W�R@]��|t�{�����m/���sy^p<�K=�Bμ��U�~zMk��,�d���冰b��ͳW%�s��D�;@��r��^�#�N��'4��:����FVeu.��k��ެ!�e��mQ��r���;F\U�vFu�H��y�着��.R<���:�?���$M.��'�G*�.\lٿf���,���� U��uݗv�O�ܢ�`��f�dR�.��
ڈ�'Q�-yh����I�qp�<�U��}=S�����x��].NH�_�ӄq^$�$o�c���Z�·�P��o®��g��Z�m��Ay�8��|�|�����E�g�l�ߧ�"�kڱ4m�B5\����'*��*D%�^���5\)��uPF�6��]P^�O����X��,y�b��[��)����F�mt��b�P���624�(eP��v7!8Q���d�Ff���gVԶ�]�^!0V���-�����=^��`��Z:u*��C��y���M$�r؝bL\+��_=z\�p�e�1�O�����
�W�F�xT�X!��n�1v�Q����A?tJ{#5�[ӀY�Uw
�j���EVz|ߨhN\L��b��l��]��#p�΢S�CK6����l��ϺkG�iO���qi�P�0�����QT�m�d웂��gg��k]6c6�xl��2lYޖ�|O9<��9Ψڮ��4�����5�;�������{r��������e�W�Oq�F�ګ�C���%����7���ok�{�qmWYm��옷R�.yj��dM�N�~��� ��j�v��Wҫb+���5�,з��ا#{'fQ���f���ۖM�o�~��^���I������5�*>�`.�y{V�Zaw;�FܨEՇ,m��,4��v�^����ˍ�QX�/���T��)Q�I�U΍g�3�óVR�c>��u[��5b�4SMq����z^v�>��k��I��ґ�N�q�߄ϕ����>>r���<8&�`��]�Y�ӷ��ـ���m5�ה �'��O8-%���S~����U��u+:����S}7��vg4���K���~l��6�3��Ѕd�w�{"
��ڤY���Lw7Ѹ�lNn�R|���o�ͱIͿD��c^B��OR9�-3�hNGn��dr�lt��r���y}&ߑ��3���8ޜf��dE�!B(-v���j�顯:�Ô�M]�'���.��X��V4�Ó���ofY}흨`��:Ew1Cl-v�/�v��C��'�껮��o09g���0�����be�G��m5�c���0�'~ZdF��c�N�&]�ة��=3+�@���=W�#!�;NUЗ"�À>��_n��������	{���]�݆:��̻e%�]7qS� }zVۏ+�t��靌F��9ڝ 2�2��O"Յ���ٙ]janm!Qu\z����J�������F8�y0k[���-��=���jݟF
șn:�h�lf�qh�r��t���cYg,�]vw���=t��^K��wX'�О��O�<�K�]B�E&m�/3Z�S��BYq�}�T��.�z�ls�g�;̂́�;s;P�}*��^ͮu6����o��C�����F�Q���3aK�Q���6��"�y�d���M�l�"�_g2�����U����uDs^��覬�F's�rl(g�X�$"*�^gR՝y��i@�я��_�L�8�"u�UEX#��I��,�v�X�/(�[�t��W��^�uڼ��kb$M.�/��壥*\<����U������0�+�i�+e{�O��0�^�=[�wŹ^k���������'KںĉG�\��Q5P�f���i.;���.�R�k�C���
�q�q[��;T�'����#�\R39�jY�_l��K��'�t����ʭ�Y�=�a��!����Hi���_��ه>^���yZr�n�Κ�"%)Gn�r
J��\i��3��S/5ᬹf�������
�:]��Y�ǎ�S}�]\�ՠ.֨*�3 ��n^ԼAū�9 �д=uyò�ݷښ��3�f��6��d������D�6n�fҾ�k��� ꕖ̱wJVtŲk�^
U{���փU
��9%%���z[	����Tu����魢2������Z�7z�J�����3��Z���L�;51;U�����w�;̙�a��"t��z�+=�M9�nD^V��q ^�JVI�ވ�ľ��)(}�fո�����������Ջ8��8�v�Vsi��N�D�Z��q�.Y�m����̀0��v1�Sv*�V�z#V9������J��X�!y������+�%k��Y�T�X��0�����b y��\&�_v��i%�ל78���of��2,Zz��#@���t���L��,d�� ���w�����Y�m�*p���g�]/��$����w#%��I9�ZqAx�7.��f����N��R�EJj�e��Uj���si�G�{�ѽA��Xz�I'�b���P hĥ*'7&ok���������Ÿs��Հ�;P=�L�3y��&��4z^�BP��1��2��#�ɮ�^K����'8���.��6��ɹr���B#�d�놏�鲺�8�Q_m��x"br܋�����A��Jyr��uY��謷�G�t��-um�ޥ����Nm�a���Nƨt��;3��!�op�w�s�T�o�u�Eؐ�p�f��$/(t� �W+��[|hL�o�'�I�i���ެ0Z e�j�\�-�e���#���K�S%d���L9����K�����u���Z8��-e�c{n �g�ނS��!��O:o��(]�Q��	�9�ΰ�:Q��um�{%L/R][v�u��g7mw`#[��s��Μ�,�AR�_<���Vd���������5�U��ߌ�����P��A�iF����U������6��(+����JD]p,uc�C���Wi�k��S����Ky�]Y˲�L�)�qQ0ܗ�/^��3���ǽƔ��u�O1�ãs��z��m�ژ�1v[�|����yǇ��ʼ�>�{0��q�ι�2;hb�et����*8�tY)S�Zu���]�g�:� J��NMk�k���e��:9�9�gy2g{-���Ҝ�4�'yc�Ob�w.Q��d�u�;֟.y{|{޿��W�ȾVs%ME��)Â,�}�.WC�q��5��	C�	���W���.�b�ۈ; c.ٓa�b�m_P�o�o$WG9�G�u���\�����jw^nr4��ܸ&�����kw�*�W$FWb�}���N�om ���m;�&�WeY�@P���ٗK�]�?q�ו���Ŵe�'JşeC������en�/0#�N��őSXސ��!h�&���k�ox9*ʕ��V�b�4b�����ōQ��TʩF�mR��J5�m(����QE����L��J5U*6Zʵ��QE*���QE,E��FTV �--Q���F��-eiq�2��Ŗ
�Qq(�����)mTY���TX��m���YE)Z-��-������aUh�F$AD��(��"�������j�2����!m*�2�QVC,��`��1F0X�Ŋ�V(��UV�X�P��+����eJԢ�(V�Z�l�*����jV

�il�*T�q.Z���ADX�mT[J���%lf[qUb(�F�"Č�X��.e�[
1��b���& �UA���l�%e��l����8ܖ���Q0A3&&68�UUb�TU�Z5�k*�""((�*6�V�"V�6�X��S-UZZؑ"��jA�m*Ҷ���f`\��aRҋZ��,��e˂#�V\ma�(�T�QV�VPX��Q`(�TTX��LT���Zɍfe�Ĩ�c�F�"*")�LeV1U �T���q�q�3%�TS)E�cE\���v:@�_I���wo��o�����v镮�wp����ڄ[�3o��4��b�d7Ӄ���s�S�������s�Y���;#��/�n��������ؘ��RȚN�~���` ��8/J���4j�����l���T8l7��&K����Q�H���5�%ˆ'��Z�r��[������p�m���Fϧڀ�.�/�ʤ���x^b|D�UcÛ����o!B�|��X7���\I�Zc�����k
>�S9G�P1|P�g�>x5+�d�k~�R_o�\/ �帄�*t���Z77X�]��}cO�o&%���ƢT,k���$���ɞz��
!��h>�]N���\i�(el[���KzwV���_'gU{�~U�L׊8�ƫ{ݻŘN�NJ5lԡꭖT8�%�R�v��Kc2��<�}�;��*���Vbɳθtq���۪��XU�[���p_Q>�W��N��C���s��XMZ嘴�&�(��t�ba-KqX)�X�\}n6}U5k���,b�Q���{�����<`�q`ڱ.��ky�xhu���.#�'�Ґ�U��d�&a�+Y軬.㖯::���U��$l^��֩�맡������/L��G��'��'�-�}6��6��!=ɷk*��D]�՛$�9
Z��VQ�4�h�D��P'�8�ڮ�I}}��'�)	������]��YJ�Ԡr�%x6*�����V,�R�ݔb��_k�U{|d�7�4��*���A��w ����	9.Y���7$��'k����[\��ʙբi��ٌ��<��n�R�0��Y,w�U�&"��n겺6�V`G�		EFDb����}�(�X2��c�zּ��Η�����e���͏��7Ƕ��H�N���Z�ኧ��qi���qr���U6��F	y�S��X�V�o+;^��M�q�U��؏��"��Ȱ'墓K��,X�|q1/�'~����f{gKvVa�W-��t�Ev�t�
IZ��bg���P߂�&*W�o�Pj�����$qv�S�V�՗Ξ�ݓ�l���%�aZ�6�o*�X����V�u�7p��x\ܰ��Bᓶn�{}��XԵ�ZSy�Q~�t"W���g��K���HM�n�V�x���pWv��x^\KrwM!w���N�7H߲6���@)��Ak�ov���C��ƍǁ=�%���8�mu�o��U�Rw*z��i�c����(�x���-;�]v��I���J��[0�Ut�PfiΙ5��tch�}%�6�-�Te����_�����\��ֲ��t>:��>"�SY�gn޼t;�u�x�٘��y]:Vw���a�����P��+5�C��N|��98���u"�	ocN�m�8��^>����<��%�����|b,e3L����N��`.s=^��`���ڹ:��}R��d������q@ê7!����y0A\)Yh�}���.��z�ĉ}Kވ�V�^8��:�^��s�a;d1���`%���B͔Yg)U�(L9��1J���x㘪߯�˔��.��LS�j����%зCK*R+X��=2����#\k�%�x̤��wO��<������P�WT��q��/s]��o�ɺr7�p&e��.
65٢E���R�{&�I�id{�tx0��R�}��W���yi����QBTc]^]��.N��޾z�:s����䒇��P^!�C��2�(z�m.X�s�Y`���c,u��G:�����;K�l��
�PVۀh'0T���ٵ���:�'C����T�?yP7����;�e��f�>o���mʄ5bY���`o�rO�^�1�n�d��4�qb�o��&�+�<� V˿yі��}r��.C^�b�dB{@��q��м������R���;j������63�MV�L�|\�<z>�XP֎.�I�sp�n�{r�T�F�ݧ;�y.����<����^i�.D����6�L����ޢ7K%M�9H�%�Xo�Yޭ�NJsR�r=t�;�Z�r���r����k(��=�z.�G��[�6�?ה�"���v܉�1����O4u�-3�B3�{Z�_�=��&�F�����:�5�@7Ń��͌jV;��+] x��v/�\"ٸ68��vT3����|�/%n�6E�9F�0R+6p
�F��S/=��Q�v�#;BA�����k����y�'�,tٌfZ�|*��uK��[\2b|D�X=�'�����`+r��we,������mLj�F��v�OtX.�t߷'f��!¡ߛ������vuݚ��%�K&w>�_��]v�n��]�Ό{P�69���W�"�jTǠ6�f��L*��	��&)��X���Y����%6�.��}�R�a��R����evy�Y�FQ� ��ޫ�Ţ���R����d��9���$qe�WAP�-�(��P�z1�����Q��jg�!�|����Gp6#��<C�xoI-D���J�x�c=�K���چyAݾ�T.�<�s��t0B�7l��uQ���B�aqr!^�TU�����'���Ƿ�&�3vE������*�SצB�nQc\p��zB�p�9;���/��\OY
���M�2�P�v��_*Wry%����ӹ[�u�%����poB�P���}K���jȶ�4��Z��B챛�w��9r\��U�`�����Fwpd/�<=�/�4
i`*ت��+k�C�o���%��J#�*8��(��Q����j���#�祼���Jv�~�烥o+.��wŹ^k�V��gC\����r�/*Tm�o���#5Eח���>�r���4�vvꖴ��D�q÷R�'�0[����Fa��8�r�y���^q��'��5��Z�z1E��\C����>��:/�;)�a}��yش��'��hi �eY���ڛJ����Oq��o=��7W�g�⋲�mm������q��l�@Tz�[����fֵ���&7�0�����Gn�L���%��Tr���څ��M�dm��Fϥj��?;(p�k��T����}w���$>n�c�F�6/6ɚ{H�+���Q�j{���7�Q���f��8�O�	*ʴ����ج�n��J�$�eX�f��Z�7��+��mO.U��o������X�uҷrӕ!�D�ڦ�F8b���Q�T2��dbwZwc=�**���l�[줹��XOhc�1�+������b�|��*�ĕ�R�}�����u�6��H>��_w���kכ�$;w_N�8��9��n�Ċ�;��̣�s�8���\�3�)ZxWf�]lZ,�#�/+I���R�T��T���  �Ⅾ�1�:��&UB��v"�lH�]!B�J�(�₧w���>�w�����e]�`�h��p�H�ڳx[����Κq~��.�M�A�BM�'�*��P��$:Ayw�H�r�.���o	gz1�!םP,�'	�3���tv?6:|���ꯩWdL�g��BV�zS��Y �y�s�7���+5_�0��%2<XJ%���T��'��S��MZ�T��\��J�v���37̘�m�a���7�C��h���#@>#����+���y���t�`ѩ�ʄl	�y!:gV�i��fQ�m�Ȭ�H݁��hcÀRb_w�p�9D�n�(q�@�X<�!Cy_=�_=�`.�}�=#�ej��U��zճg�.��o�$;��{�듃|���R5��.I�U�O�<vِ��f�8��[��
�{��m��{;�T=�D�ժ뙗�|<|����Fً�E'Ip�X����c>���`Y8�U�3j����<�`�̔7�H��K�˱0�ZJ�J-7�߈f�׏�o� �g_r-�����R�ܛ��=ۆ��*��C��C"ir�uA�ȵY�)�ۋ�[�B���m���Ab9梵^9CᔱE���N���2v�ZAA�'��+V�AL�V+4U��PW]�S�9a:ܛ]A�UȐ���ѹ��c��sx�wꪪ����L}��d�G֕I���4�5�fQ%��r]0���C���^�s_*i�?��5Ҝ��0El	�n2�Q�3��-j��q�lE�5PD�w�$�a��x��`cFc{�R�b����9�u1�F�F�!yt1���#Myk�x����F4�fb�z���r�@��2��G6��P�W/*�<1icc���۴�x�8箦��4<S�ȁ�,�9V޽g��u����IX�e.X�s�Za%�>�5%ժ�CW���uʬH'�O`2�nC�:w��!8�+j_�k����H��M�d����l淲��x�A��K[#5�[�^~�!�R�V¹h����Foܴj=�u�2w�h�urO8T3u�-z�,�}H�bV���_��Ac()�;���K�/H�lS�f��"�7͎��>K����d���޺;��qZ��{p�����gZ�}1��D�م��x�G��P�]�z���4�o�I�S�E�t�'��{^��H�6ޓIa,�ZH�t�x����v�Nn�r�T*�kc��V
���z�;ehy.�L�Jc]ԸBo7�r�8v�����n��-���LmK��������7Ӫ�P42	�9ǚy"cpʆ�����着l���X��`r��v�65]@4���yD���!P��&�t���D��p�!��L�&fZ���ixu�Cϗ��:�A[{p�
��s�U����d�T�.���Xn�]�[<��5>��3o��|f�;�P�h6�A�(L���H<ഗK��9M�h7�`�	V�A��,PkoZ������x�J�W�sJ	bC^�o�(C�F���ı»Y��x��SR�bO6��d*b��k/k��X/%�Lv܉�5�X�׵)�G7�-3
o��
�O�yM��C�u��82���>ͬkƛ��ϹkA��5E��(Myk����v**V�޾D��og�%�=�ɳdY�Q�2�k w^.��f����i�6`gի�Y�����1}ʳ#'�J[�	T;���1+-b=>�U-��X�����b|D�X=��h��G¶,��;:����Q&�x�6G������7�[J�^# ܋݄�Vnn;���~������,�Eڧvw���c�ճ*��^`�*x���9S��':���+��g��L��A�'s�:���RI;|�	+h��i�R�>̻���lbn��oi+.�%gT���߬4�kg8�;j\sFp�ս]�M8����O:��� ��������W1��&y눮����qE�s���+��>�]3�AK���n~�7�WZ��N��H�D	ͦp�T-���*���.��VF��{Xw��.�j''K�X���5��ʨW1!@�\D��*Zۂ���R�k�ʝ���ŭ�	͜=B$4z�!���<'��Wa�Ϋ�S>�j���N���xn�Qx�Yz�U�]��~������:�(h�
/E���dM5�vw��׊+�i�0M�����p�j��Wr��d)��$,uP���<U�����ėC/[`�Zy��i��iW"0�B�yeV�`C�8t��w����W�V�#]rO�^��Vk������yo^ҟ��B7�j߷��{��Ϗ�Zӟ�o�;b]�(�qd��h�-�%=�q5��C���q��.��s����2��p8)��ى82��tI5s��H�
�=�g";�8g�t�G��R������%u�>Oj�ґ/yxR�7�/78��<3yv�}~p�B�W�� c>�|7��}5PWf�u&Ku��f��R�yTE{plP��|ιYW�5G�����b.�;bz�F�0�MbF������@��,wWf:����s�C�9��;��D�>�s7 �]B���]w�V��w���x�8vHR��80e!���:�^U4��p�m���ŗ�#��:2���zk2>S���B?{��Q�Dds컣ad�C���g���Ɏϙ�}�X�����qz�q��7η�ɚ[L�(7���5r�쫔�|6���r����A�骾�]�Ɵ�:��R�♱��=�;e��~�#|�Sfx��T��P(����EX[)5�xk�}~���ֲ��mD����dc�+�u�_U+�(�����ޝ�(ԦL,�)�mW�c��œh���g�սU�T�8���';�s��؝��/�t�����rМ�" ��m�g��E��`|e$�z��3��d��JF1Aq���L��o�����=�V��k�g�5A"J�bĵ-Ģ������ϒ�H���D{�*��Ms�FP�9%׭��%��B�'���	9������|$���__ʘ���Z]wێzQ�tz��+�.�f���;4l9;٦�(|�yPz���Q��=�FB;Λ{���̅q�H��WJ���w	�:���O�>Y�rۥ�Y�t��;�Y~񑽀�{�]�w�D�n�7n��`#��m3{(�������yF�'6XKC��RP�'��\�,�M��Ui���%\�N�a2j��N�\w��J��j2�p՗1�r�rS�g��v�����P��Օ��0����Ӱ5��b=*P{�Uio\'joVn� ��&VA��e�kp�`�~=��ĔN�Mo.w=�r�8�2�{pqS(Y��v.E���53��aУ�ь ]ӡ7fU����ц	L�)e8.b��W\��{8<�GR�1��K��P^�Vd��!���]�%@N=�V���:D)���YPK(�s�J��;��+_g�y`\�+z�BN��D&7+C��DP`�θg��o�嵴�$��W1{R��|^�-h�k��*��f�K�[�U�h�r&y`m�#�ړܑ�(�+���t��oa	���Qɪ�_Z=�l�O-V��tG�ym�� ]V|�%CMYԭ�w�8h��sB�0�J��DT�6�2����L���l�t]�k���l�a�����no��$ٴ�%�h��H��D���Ql^�*��K(��������o{�]�+bܒ8�[.0�˼�l���7)"BT'��]Y�E�&�o�\j ˺7ou�1Er�$j�fa�y��Y,pTgbέƇuq͡��rӆM�y%�
	Q,��YgWK�Yb�����1��D굪���U�wg;�gS٬�]���Z{
|1��ݖ�<;�&�*�-��K���]�s���|GVt�c(/wTނ7�R����3��bS�����RZ�ژ+��'�;:��{)�����srS�ѣ��q��5���(c|�CMڎ�w_�M�ɹVEwFg�r,�nVwkn��9-���)�\�r�L��[�e��e���f�6Hi2C���]f{3li������O`��3=��8w�̷)��ͳiTH��
HHF�p�}�L\�s�����l�}9ˍ7�Ѳ4�,���ؔ�V��Ń��A��.� ��]&�=��VN��EZ�-��s��rÅ�����2پ��I��;j���X�E�&u��)K���w��m
̢^�q]$��t;*kl���e
g���M	�[��9ǱwZhs�+��Ϋ�L"^򶴂�O.���ceJ��������ɴk�,�Zڙ�<�5�1��*"P���4�7WJQ�X��{���$����bE���˶�k_A�\謞z��N��W���^������^H't���ki����э�WZ]�_CP���M
��9U�0���M��1hU�Wd��pe�G�)D��Ih�L��.�0�����jJ7ݕw��d(Fy}��eέx.>X�9V�5%�;V����0����5��L䃟[�Be-�ڝ�NU�^C���_te�-E]\�}6F�t�6';e>��BvF�]e�+�1}z��jt�|f
���S���_WK��7w��~ߧ�1�b
���,QV
(������QE�(�P�DˎȱUPPW+V"*�-(��$P���rՌ����c(����D��*��J*�fR�\)W0�b�Z,DQb+"��"�Q**��((�S,�ZV*���@�Q*f7(V��U�"21$X�"��-�bAQD\j*%aX�PUYATcTU������U`)Z��m�ʱU�eLj#A�+Ke`��
��TU�R�1Z�aq,b�Q"�)�E"�
�cQ\s(8�UU2�UAE�h�UUH�cP��E�����TV-lVe������1�b��1Y1,EU�QFe%�Z",AUQT����ĭVR�m��eL©",blV8�F
*�U\j����J"X�eTER"�j��b���(��UUUX�P�*���DDURڪ��.3(,V�b�mob)Vk����X�L�]��3ZX����J�(Z1�>�vs��k\2P�6[3{.M����@�Et��{�J���<���]�5�����L��x�	��!Pջ��L��u�+Pv��z־;��K�^f����(�;b��]��<�:"�Q1�w �h+���!�(J�ad�h�,�����λ~��]�3:�X=�W����|��1yh��ᮋ9��(<���v��5��>��<��U5���.�T��H��%,^�؛����7ཉ�s�7*�[�'t�]
�/3o�\%(�;0�oT��w+&iHj	�6eh5H��}�b�8V�Ǩ�\6QJ��מغ�!��Z5p��g��`�>pX��Z7jW<�2^آ%M���]ܓ �+O�dh�SJ�eU��!P����1uk��%ٖ.:HW����g�q�iE�d�]�=>�/��&x�d��BY�]V�o�L��1pՈfL�9�/�f(�(.��J'�>���"��Xϩ�g/�Wh=1r�]N`'��"Z��t�_���Z;9�Ʋ����c�r�)F�7��� �/O�q��u�*���6��+˷�2e����Y5�Wz����7
�tY-�-�ݸ�S�����VH�4��g�e��N�#�3�v*k��ne�,y%g�9�з�>��[IE(,m�[�RV���1-4����v�\�'Q��J'j:]�y��8�7�������]@�'�[|���F9d({A0�Z�5�[�g1Uæ��UaЭG���_� 3�gg9ry��[B�>o�w�y�P�͖Lw������X��9�{PU��8���)g(;5;���Eep,DYB �������'�/��Ʌ��]r��N̣۷��X�m�t��`�Aø���#�����5���g�Wq�\,xf�v؃���q�756G��չ$)b�¸��f��@4��L��,H�D�
�y5��eoK7Д�=I�����A����	�<�KQ���	=N]Ú����
��s�U�����	S�y�9P�<�q����x�ً�����s�B5���T!�bX>���ഗK��9��Һ���L������y��7�d��+�U��a�+`���:�!����kJ�rJ62�G*�{����yz��dV�X���L�x$5�J�2t���]�foo��%�lX�Y�?��m����+g���^E�V�3eKGw�����>�a�+9� ��m�b2Wu������/M2�w�-%!��n�e$;^H�Dݜ[�#y����s�L�Skl���������nJ�]�u;��]6�{���n=an��Mo���n<�e�c1��Z��v�̻)���.k�j�6��m�O�UQ�=�;��5�lq����:�!>�A�P��<=x��qps��G�4j�#�]�L����U�cE05��>eqdχ�c>�Sp=.�CU�//�c.��٥�3%����yr�}���ob7G�ˬ*�uDj�h�O[��w��}ZlnV҆�.!��1zإ8J�3uf�����k!��h�63e��n�v�ݝϺ1�B���j���%�w��:��b7��*�"��^��qr@@��t��3�����E�
��3�]6�W�v��v���b��z���Pt<�0,5�Z�]*C�(q�>��B[pQE�3�]r��<M���U��L�q(��ߗzD�p����:�G�X��.b�\b��=��%��d]����m�
�������k2Yco=v�Z���x�V(/��6U�du��t�yg�J�+6�s��7n3T�NZ��b�,t�N�2��$�C��Dp;
x��E�qK\�Ī��lij7yx߸����Ha}�F:�ze�ެ:p\�|^}q�Ո�2P �rWCW��i��d�9�E��.n��F�H�vmgc�ofE_Dt�w�}�fƋ^�z�ʍ���9L˅D�S��E<:�{�ޥ��^�yR��G�{e�1���ɸ��t���Tv%!��}Qd����uˇj��]|Վ͓��S�{�Z�㗓�j��3fo[�U��{��f����Ҳ�ʡr��������>n�p�-iρ�=F�qöK�|uɺ7��]m���3�)�$_��Խ���br�+�nR���b��U�;�����:2=��!�'f�g{L�Lm]�D�3qQޘg]L�{r�±��U�l�I1ިEdGy����'���/~���Լ�A���ⶡ�e,R��@���S\=8;1c>6�{����/����6�!��"���a7U�G��r1+�>�Ç���&8N�/����������H�n��k=��87�0��vL��I�Zc�����V�Ο�S;o����x*:Q��9�R��YC�Q]Ɇ�6$��n���K4t�j��=�������<X8�IȠW"�����Ļ�=CI�H�����L���uR�F8b�ˮ*��\i������#S�U,�T����`敪�������}U�KP�L\(>��k��J��N8N푰����2[j�f���f��|��F��,�{I`|g�$�z?0=^ :����\�5�Q�*ʭ��'�#&N�پ�(Rk��f�g��W��Vr��R��� >�Fv�ns�������k�o5;��;Gs2�7u�7��*]��c3�'ob�G#}�;�.�3�{����(/���kL�z�<�	�Nj�5�j��oOr.�7]��3�3�U}��O���<��Po�:�ڰl㼲(Db6L�-�)y1��V��͎���R�4=�Σ�s��]u
��	LZ}�lC/���v�`饏\�D/�\K�Nk������P��.W��L\�'��_�:df{]����ɺo�i��UF��=��w ����(L<��ʢ�4��F��-���P��桺꘭z8wڣ��ӽ�F��qK���ת:��ŕ�[][@��!�z _
�s(��x������q/u� �MEoX�OжdUT4��Υ��y�~,ϪXp�2�G�\�}2��#�-�
��F�������&�s{����Y9x1�T0�S-�'+;
cI1ґ�W�J�)/�E(����vw"P3���nR}�ʅ:g���'�}f7�dH�G�R�ǦI^�����:�^�4;�U�6HC�ý3s;9���Z*G�^k@��@�!�&�2�4����hVvTdx�����9Ә���S��¨�#a�T���ˍҚE�07�l�G���J��h��ۗM�N3wz��[���+|��|��q�v��}�Z����k�)�R��ѩ3O/�>��gj�ώn�Ϳ��5�a�H�y�̸�;xb�ַ+nf.��kT�8e�!"��/�-�;ghK�F���z歵����r�{�ݹ
�� ��uR�NV�7f�g��ͦ�̙N���Ǎ�ּ/-���)��K](��7^c���ly{/���V:�Z��ܴ ��mi�K�<a�{P1i��O�.��:XB�s���ՋbB��:g�����LZ_چ�R�V�`W�J_�4T��`go)�_��u�s�OM��`V����s���v÷:w��/M��*��m� =*�;�z��ы�y�A�����S��,�
_XxK[#5�[�g1]_@B8��~�r��ܮ
�D��t�U�H�f��f��ܡV��T��Z������<�	�Q�޾xD�X�r��� ^JW�_�lA��l�h�GG8�N�+��(�Q{��h|�M���읎�B�.\&���ΆI�+v�:f�,�D����Š�0����:e�f<�����.1��E^ѭ\C��jz�C�e������<�Deq�����kTB�*պ{�%�5pd��\�g���;���4���;�.�`'� �	�^�<U]S=[h˝	FrI��f��r
�g5J�vWK�0n�; Ps	.��muY�s���d %��Q�H��=8�~�;��_r��V�K�����oB���+z���ѵ9駡鄩�y8��8�
��N`��ȷ�h��e� 7�p�r=��$��-�{Ǩg���yM��^������kA�*�a�<�$3|k�F�-��WTʯf�8�,�ݾkts�7������xө|��=p�%A:2��9�x:�!�]���V˸<���B����)u��i�m����������]�DȔ�	���9�Nm�[7��N�����œ���b+ʳ�'k�<}��^,+4��S'~��*��LJ��]��vb�׹&���R��Yч��b�1��
��ڄ8
.�w�r�z����;P���6�ote���[j�l�y���T��Ψ�Á�oc쵈��U-�K��J��k��1�ҦJՏN��'yiA~S��66��Ѳ6���<P�6K�Z&Wr�a�V��j0V�^7�P�o<�������>�L^�0�"X댟y˳�:1�`=t��@y,�c����V�9z��uJ�~~��w�'z�.h0��&(@D	�L��^��2��)t0�R���]'�Pz�q�}Z�+���/SԈ����䱟kEZ�U���ĩ�q���>��|�2u�K/izWb�X���]���+]mAP�u^4�)�ee�j��t]��3w�6���\��X�6�T�U=���j[�8����v΋��1�8ī����n���X������%�wX=�:](k\c���gZ�ו'eJ�;��D����~��v>x��ջ$?���=��p཈g����0xo�Ih�i
�T�h/᣼}�Npv�����'+�D>��m���u��x�����kW|�|^=��1~lp����3�Z�����)�5��ꈃ�)d�t���˞�9p���5�!e_�4i�v�<�u�O��껳��V�=�<�1��D�Um�Ha���=hxyʳ����q���"�D�@�1D��ye�c�O.HL�)_�]
���u��-[��ؽw�����"EX�|�eT���a/g^��'@���+$�����G���iw�pu<�Y�t��Sƥu�".z"��y�&�<�Z-�뜐xY��8V���j3�]ǵڭ�^�'�'���v�T�]/���M��]�-D(���:k�.��d���P�p�n5��L�9�Lmq�z��&5'��3�F'��Īb5�"��;�z�J��e��E��yYGЁ����^FM�1���t����n{sU�&�[Zg۴���>}�ɦ=�C����v5�P�7*2W%�م���:����oY��1�N���Av���]�~���Z���`bR�fa�;����pc}C���.Ԝ�3�*�	�UuX��i���(m��0!�x��o��ԃ�|��s5'�a���.�t�'>��L�<��7Wb6��k�읝V�Z�_]��߇�u�r���t�|l�4�q@��n3bJSe.�h鰵��m��ʩ�o�΃\�8�}��ɡq#��#��N)��Cb�"'�P<�V^A�3;K�>ɳ.[�J�E=�r�,�����g�[�Ú������3��5}%C��N.+�YY�[=1�㷶\r��qcg�l2�9�����;IF�,��Ih��������q�Rj��Q�ږ�0��0�).(��'��b��ITX����T�U�O���>�m%ۯ3juf>��4�_D��h�$���ߡ��E��Ӄ��=JdB҉p1Z���t�^��V��7�ّ�bαR��.VE��Fg�1���F�rw�M�P��6cG�%V�/;V%p�D��!���펿H�νu��C��	�:��>��fQ�m���k-�Ξ��ޮ�q�N0�����'9�d����B�纬|������}q��򠔏�)������*i�^��ΞJ^��%@H[�t��
�_¸b���E���h.�s}�b:9�N���t:��<�a�3z�ҙ�.�)�F�\�su���w�oL����m�n�6�I˖���s���G[�!G�m�6���!��z�r��U���F���]׷�7i� �G����,��g!��^�]�5����5��[{+���ubzRk�����8mLi'ґ�V*W���*r�\ȷ֔=퍑�_���x�����R\9x��1�`IH��F�z7^����+���������zf�g����Pi��8cO6:+�Q3�Hj	�6eh50r��U�(��k�����$�*��P-蕑��U2(=����5-tZV�@Q�=�֍�dܛW�w�$9����tR��SreY�1�����0��� �[7�Z�2+�-=��q<a�y'�7�������A#��b�\+��R�w�W~:��P���7�H��7z=Z!I�kxZՖP�+����P�(���Y�F�Y����>J�C,�`R���5�n���{y��ߵ:��K늾�V(t�0[�������/O����S�^�*�ӽ�K\�����=va�N5�� �!-�X�L�
_Xx��;��<����o{R<~��`G�!�{)�dVcE��B,���07�X<zԨ��%��薭��ͅ/��%oM{��A:��d�,Ts��v���tr�����)���ɢ�IX9X�,�;:����t�W�X4���YZ1�n!uω���&���i7����&7Kl=�y�c�����Ver��%wWT�ܛק_��	I�\���B��W$6vW�*�{�l9�WmI�k���J*�B���0�6]�\j��)��dX��ÝV�ǒ�m��v�*�+��[
�����յ��mC9��I�]�B+��tS�	nW]Qsm8kt�y�����u�/��"�X=�LKW��lܧ{��+N,�}������*bYie�Z��,�#�j�
bK;d0�f��O;��[4��L.K��ƺ,p�\���C3+1ɬ�d���S! PpX 9o��� P�l��+s�]#��ܭ����ʖ�J�7*aNZʽ��|s��[��.E�|LAE�R�X(��sy��:�h�׀S�����֫k9�.DFu>\.���9��;qM�&�\��U�eN�
�VJ��U ��O0hm��;�(L�Q�9j�&7��ݵ���&�_���ݶ���ټ-;೻&80B�[J�ef�N��v�r�cݗ�oS�;̔�\ߚ{��sq��us#ڕci�:t�߹N��:(TY�<��[��-__N8�7g0����W|X�T�e�j����똵z+v�t�a���9[mK놓�c:��,ˊ%vK�0�����Ծ\I<�.�d�����u�aĝI�Ub)�ֹ囬+ ˳�
����	��Eio�n!�WƉ�u֋�P�m4�'�8�b���wv�6E]��|�{
�I�ec�GHff���g.fȞ�v����.�ahѝ��u��R���[t�u���3.�!Ư.��vnR�(omH{v��h�)ҳ���p�Q���Y���f����NaQ��upY[G�Y����;���{ۘ�Vғi�S5�܂ė�۾�Xz����QB�rQw��\;���9n�v9�(Z7qY��Lڻ.%�����>�S�\6��$�r$Ef��}�G����s������ky�|F�/�9Z���N���F:S�[�^_v��Om�Go��phu^��B�>Ti�׹�C�ǝR�D��	�,ޱ���*S�_V���FM���Ε�v���Ӓ�Fܬ�ԡ�0Ƿ��k3\���hq�.N*�wtGsx7��髼���f1�ei�����)���0҉:z��z��	�ǡ���Z�i�y[]�k�v-��˖-�م�x��^'^�	�3z�m��bH�k.���}f����gt���_k<�F������(˙�(�
7���2��m#�v��Z�a�6	��`�EQ73���h��&$ۥ��7��6P������B9�D�s���jV�:�T�"��i��e�^v�Ր�\�75��x��SX��jYDQ<�W=wX�����.��n����+��F�u�jlK�@��JO^�!����̬�t˺�o�4��w��IT�,X�h�A,P�Q��J���mmUBڋ[*6�E�4h�V ���DQTTb�QX(�E"(�V�b�R+jёU"*��eT�UA�%��0U �)��+E�(/�U�ST��(�E�V1EUX"���ʌej�"�V����V�kb��j[i��b���(#2�QG)D*EA�*���ud�b,bDTkX�1U*�+"���[(�K(T\�paD\J���Z�E�Da[�EAAF1TjX("� �"֊*
�&��Q1T��X����kDŊ�fb��ɂ�R�*�b���*"WPV�PU�2UDUL�cZ�b�X�kH�D�)V
+��Ub(��Q5�`�)QE�fXUU��b�0h��--����"�*�EPV$Q[j"������E�U2�(�1A���b�\c��Ϗn����Fl�G{˰�n��s{M�6�J��K}C4
O6��#'K}؆<�	'��s���w�$5�}����VLN���z���#	�\%�F#������WDW�E�k�Y�[�rT�D�L�E�Rw�V�v7T�wg�s˂��2Jpa2�Ѩ;�]����_q�n[�g�;�*�w�[��[�7��7JY6)�ۋ,4�뺀S�Q&Y�"\d%�T�k��0=�k1cFw3���K��<^��qF���n]��t��\�����
��U>��U9�'�J����9��-��P~>r�m�we3��!�h7NYȐ©����E���o\I�������ލv�6gE�.�\2����l��6�w�%�ϲd�r�L��+�6+G�)��v$}�^��ayz�1a�z�.�Q�P������V��}\�wEѼ�}�����,xJ�!�=Cm4xm�g�;�yjֆl��M��đu�Wl���`6�[\d#�~j���}REEwQ����X�]�p̹�{�꙽س�-��f�8��|���Qc2g�̱��njݞX�����3�X����Z����u4&Vwjΰ����CԺ�{��+��b�*��r�ӄ�ȉL\��ۢE�`I�S�Ӆ��u�PyPp�g;Օ���HEh�ќ�Nɽ����VMΤt��I�yu�x]��n�'�_;��PuwVӗ"��6��k�t��׌��l{�m=�=�\����h���}ѡ��E����{����e���^�W<�2TyDl
��M󊾚(��E��E�uG7��-�a��_��7��܏���{���;�O�e�3/�ެ���R�&(@B��8��(�����*���yK���7��*zR��vg�u	�����)��� �Q�sBXϢ*�S�]J�p�75<{�w���:U��m�X/�6�ȶ��}�1p:�L؅0���8�&g���;&��ڈ�2k��5�;�}ry��Z;ѝC��j�5��tdn��r��#��^=�^1�2.����o��8�G\�[��ΗV�`����m��y���c%��^K��d
f@|U���}�k��rC�'�i`]��]����
w��#z[��C@�Rt�Y
��*�'{��{�kA?T5t�W]
���J��-LoG��/]�+����q����]��;�����vP��H	� ���_�����'�kŋ��oJto���>��\yV{`�	��O1��r�jMS�ק��%��I\�,z;�8+;=2���$���t+�h���5��P�Εo\�E��&�8x�w�Vgu�Q��r��ɨ��]k�t,������눕���$[��fVeӾ��}}sfꫥkV�C�f���;N�쳂��Q�au6B=C/l+�NÛ���w��dU�\�WNY��ؤ���"�]�l70�BrN�f�Ld>�E���J-�s��h8�SU��������Er9ѓ��S^���� h78�IU^�,�ދw�+(�~�d_.@��������Rc�|�l</��O��dats�el�H��j7c�<V$H�&�:������a#0������jq0FR�f�>����P������5t��iGNV�f!3���1�JՍ/ݝ�Sw.�����WU l1��\WL��%��rd�*�ĝ��U�n�R��l��mT�sCUS;P�e���lH��𾒡�u���Qj2���YD��c+n��Kc�a��2��}L�9���V���48ɷ�ʩ�V�B��u槕����b�
���L(t�0k��g�2:�\TF�nE˚(��d��k\�ħ/
~�E\�q��7��Z}�lC/�������!'4C7���F� �Ω��ٙn���]�h2�f �T����[�������ȩA[ܭ=6H2��C>AӚ���ݼ4t�ش*��r.{֪6�9�>�H���}�f+�ӎ,���
��9�^+B�OU�U�*���o+GLVUl\����;�޵H�gr�u��Q�bYS
a�+"��鑙��t-��-�6Y�"P7X�u����i@ꃬv��>�8VC�	9P��o���.�ul:��O�e=w��ؖAF:��{��&�\�)h�XɃ �H|+���w��.�e�Y�����P)>�R��;p�{���jȱ�SRuKZߜ,�a�#))rN��u&G{�ב_W����|ۍ^��bP����k������Nb�r�:��1��JG�X�\Et&��Ʒ$/�㥮o�������aw����'>���2����k��d'uA�+j"<��ǐ�u[7Dtf�c���ҥ��D3X�i����d��<�r�{��|򞎫���%��V��y&�\��P��p��W�X԰�-)�8
,l����ԍ�J3�dᖳӟxt1ĵdW�kڱ�Y^ږ�8��� ��c��k^�[� ���7%R4��=��&�'b-d��R0�{��\�������p�\��s�v�l(�44�����M�����G�:���
W`;K�@�i�lԬ+�J�Y���!X�v��A�G�Le�1� ��WCfamvض�(�9����$��8/{I��_G�6��:�.:���-Će-�F;��Zv�uZ&J�w+�Ka��>U�촳��81uC�9uC4Bp�)�{���L�*��X�i��m]�����u�d��/׻+��^E9��g0=�}E� xeOc�U��(t�0��v� ���.`�
�J�t�ԫ15��o���v�-W\T^�#�<*D�#�?�S�L�kdg��[Ӏ���#{��+ؖ�;qA<VrhE���#Թ6U@x�J���K/pvK�t4���"GVb�Qv��y���#�T������Q�����<�Dw�q��^|��6Y0��n�*���dtX]с�{'fQ���f���0��;�]���H��jy6��wv�橞��P��ҍo�ɗ���cn��7=��'��K�x�G�0ˀ��lS�����(GE?@}�^��/zvT�����r��FÕ-]Kz�2�=)%bo���Z�|J������Ƽ�c�����Lk�ß�oV
�8|%T9��P�p�P|�gulN"�5=���F�Ub$ׯ�q/�::�7����Y��:��%؅pʿ4��l��#K=
��{^LE�AY���*f)C��xM�� G)`e���n�c��)\��eE\:��WZ�U�!^�H�YQ��2����kG��yr�����u��_u�x�H܇x�n;�����"��g �v�ӛAu��EWu��ͨ�n#(��.��&���JF:�!�y�+�����+�?�NZ�a��}�l����r{Ŏ����^s[�/_�ym�j�����X�N�-3�hNGn���i�9�ţDo��=���_��y:��^�Rl�fb��s֎��Έd2�t���"�g\���q*���J���[Wu�ުGXs�Q�h�b��t����J�y�2��ջ<*�]Ψ�/3��U�T����X}δ�{N#c+L��3�Q�k�(\�/�K[�����x���,�U�v��kU�C�3³>0Tr&/��y�����e�˳�х��{�����#���Xʞ����0i��<Z)kA��C����
�8�	EE�h"���e��C�'�T�j;2wIW�]�E��=������2%G �>�Uh���U����+�q�>$���ޣ��XSӻ�&��iy�����F{X�f޼�Q�Xi��0�8�30{~˱SbT����+�Q����|��q���j�����C<�����f��z�r�)
��t��pڬC����n��9�2S6���rLf��ݲ��It�n )B�^/:-���
�<�{�ׯ�]����㺭<6s����i)y*y6Pj�uK+rJ��0	���7�F�������P��,4��`I�K5;������d.�{�`�)�ʢ�L�p)O$3��}b(K�ޝ���V�$*�w ⣚���$�r��$TAQ	�G�e�ʈt.x�4)���E��l��n�`�J�e�Ċ&�;j?=^A �`�*x�',��h���ᰖ]9���G�P�x�wc-r۳����i�L��(.��Ⱥ@8J�
[�t�>îSu�]�\3}e��s�V4�pa���C�����0��C 1�jϤ4΋Pî;�0���p����<�7>�딫�5m紂���ܤ�Q�
u�N��P�,����Ĕ��_�'K�چ���K��f��\b����1�Hv��[Ǹ�v+��j�m�Z�r�����wZ����y�ر�H��c�6˗��t��Nr�m}y
gK��߷i��ha�wK&���I�1�J�=]���.�c��.��]���>�k��߂�,j~O�2�qc6h�cn���K4t�֮�;����V[������Y��Ǭ%�����7���O��6Ƞc-��/S&���4fܿM�,Wd4�'��صp^�IW��[���h"����!�s@>�ƞn��U�����w�4Q�b[L���mJK�GQ4�r�U���Eݛ��w����g�*����VNd}W#�a���!o�/��n�⡽��'��ةg䭾�'f�{�G��>�sc�n-��]2������UkRǦY؋bWH@�sy��ɚ�ҩw=�Iu�v6�#�S�v�C���(�<�d����J7��ē�ϸ�Ku<�.��x�t_<Y�
Iog�5}$�b�).(�Hv����!�e��*�6#r��7{�;�.�&SY�y�1(��UEX-D�$,�PJ�Z}�K/���b{zyᐕ��n,C��Ү�]��9�:D�"2!J�혞.aL#��d\'L��D�1����}R[X�9�1v>}�yy2�{�2��m'����{T���uB6'��\'L��u��.�.w#|�J��CS��ڢ��Yn���Ʌ��H���С蘾4<��w�f-๲�w=7��sD�Q炥�ej�W�k�~�lةa�e#C�:K�.���p�t�	�N��Y��ś�[�B09���N�����vLa�=)5��br����%�#֖��P�ɷ-��ǳo�U{���W��=�QmY��%�}�7�lIH��s�]�K�P����'��%t��`��|�>�§8���E$9^��͵\i�D�.a�p��L�b���l����%VX	�6�\��EX�m\k�jg�.��k�B��f�L��E��1Js���kP���N:Q/�u�`XS��Ǜ|�tna��)� :w�gkۅ=�3q�˻r�$��Ώ#�}p'wW(���f��ʉ�R�i�(�A�R���׃�����Gl���yaDu�·�P��nA��|��k��_ٯ�֖uw�,�$�sۻ�mw],�G�E�ڮ�"��^׵cb+�XN��x�EN!������ɛ��q���y�p���,��C��7��Xɯ��}�X4?rЃ�miʤ�a/��f^e�v��5z��x�#�̍�9v7��S%C��{9��
b���L��n�z{4��Y�o�_���ORS��5�L���#K$�����SA"�0ȻV	���;xm˭��+{�E��sy���#9#ԺW?���W�F��	n"�:dW����D��0k���t�;	������y�Gƴ�C�O��bF���*"�!,��vK�t4��;��6<O�uٜ�(b�n��:<���Z�#\k�iq$Gy7~�]^�E����&��{z����~�j�ߩH�����z��td��:
�x�G��GT��a�@v���>݂ۼ7<+"iSӤ�FՐ���i!��o��xL�ڏ�hz�5X�E��X�������M�gh�����T�����o܃��"ީeE�Z�F�.Y�ji��$����;�p����wk�EZ7��Jt�΃N\#z�=��!^k��jwo\DB��>�t�V�\��sb���J̳�]�I�(��g�u�3e�N�un%���O�>Y��~ɨ�����S�o�y�le�wM�r�!А�<�(��V�����om/H�|���>oF�T&����{Ӟ����]S;��u���%����
8k���h�b�b 0ў�����������Cr���z�ל@Q��zur2<��gܡZ1q�tΩ�!����u���2�,e�3c#��BcɅӢ�v�P�.jq�G�f��3���5�J�2u���a��tסmY��5��W�Emiî�C䙻�;}�㯐}�1('@�{c�=��ذ��Ӯ���6E�]&�(�/6��.�qWk�_�Ɵoe��hDU�C9a�6Ƕ_����\�5ibvu�+-b=Q�sR�$���U���-\6�[��ӈ�V����t�#=�8��_rٕ܄��q��6�3~�^g<:�3+Ը�.!��Mȟ��ρ��k�������u�u�k~�My#�#Re�`�e����4k[|���u�c�@���_e�U�ty��5>w�!&�rVU��&��Mw^gZ�=8�КְfY`Y�S�����_V�렔�q�jD���t��O�ݢ��҈]����,�݆�Ɲ����e�ǻ0�Z�eb�>�G�[ףs��=�d1�CM�����:nK�/�H_
����37��	��ج9�Ǻ�̕+VB��u5���K;�+&)��{����j$���u��u����syliԭ�YTƼ�����wHW16(��lv~�f
�n��G��rթk�&^�GU��ua��7��>y�jqFX��uIR� ��h��;��.g]����8�r���w`\I��"�H+@u�83u��@�����NAU�HM3R+�ʸ��v=]5��z����v��DLk�O�yW����e���]�����뒳�\�B<L��Y�
B&sB*E���h[�Uh�0k"��r����Bf�3N��s�6�t%;MŢ��0�9�:��W[L�{���=W�n�Nru��"���ȝ�,��}pf ��*I�-����Llɲd�IK ��R�+.r��%���-cGs$���+'wA��u�׈�B��9��VSO��$f�Y��Uxr���S]ղ���B�uga�Z���y$x¬���r�L���:_S�5[,�X�m&���X=�%�WbZ,=������V^�4�IqN�=��I�۾�]�Y���?��f���{�����������_h5�iA[�� H��nN����C����t6�#8�]��oh�-����
��6��M����ib��SW�0����-��j�o8��r�e+��S�C�XM�N�s��]ʻa�	��[2�^F��r�I�ER�`!��nN��-d�����J8�t����A�	�����D��R��:�9J�=�(�cY���+zҮ�|n�h]�ki��8 �#���4�{�b���WyP`��l�`E�2�u{�Zz�ۙ�![Ժ�,�]�ðWs�}�A6�g[�p��Λ��yWYYܾWջ��,]��61W}!�5��ǥΰ�vbP�U��VCq��uϨ^FN��v���&ŀ�vgw״�wJ�a�"�U��Ӣ�Ap�&M��y��[\�,y�׭�=OD����iHwE�k���泙z��|.!�4*��m:̕t.rj�Mf�qv۾�9 ��[�y��[H�<d��Y���]�f೐�ɡ|t���h2`J������ҟGVF�(w�˚�0Gh,<Y�f����\���S�m���|o\�ٗϚ�go��c�!�c����Y���K�0��L؜�X�dg]�Wge`�sm�]b�لS����aPqu2�w-��tиz�e��6�lo������(�dl�:l��#�d��9v��gmgNv�29>��p����[o��������Ib����V���Փ���XT�%�e&Z�ib�T�AT���ܵMh�Z�X�رCM2����#s3"��6ؖ��m�b#��U�L�U1iTT\lB�2U�PYV��q(��(�j�TU�DQc1�
�����*�Dr�)X ����b[(+ ���R��-�(��r�X��"
(�m�������:m�X�EI`����+�
�Fڢ��e�����b�m�m3)�EjEX*�U,bȈ)-�cPF"�AAd[kmTEE��T*b�b�SF(""����²�U,�L�,r�j�1Q�,]&8���ɑDX"*�����#���-�(���Tb�b�1�� �AAUL�V��fIbb
) �,Eb#D� ��Z�Qc5�MTT_�\��\
�}SS��Z����΋�����G�:�|�ua|�˥����\���ٴ�7c,��.�RY)���D�-�}��_评���A�a�eYxj�H�! N�`�p�T_��.�-���땻⛖$��a��/���]���r�뫸(�FQ��ڇbbGBP��xx�M�Ѐ׮�PE.B��s�(��<_�>�l)u�0{X�f�E6e�S
G�X3ŭ���B�:��kฉ~�Zb����f�.*�뒋<���Z�#�]�EØ(-Mg1��P7�_z�^�*66rC������|�t��з�ا]�v�C��(k�B�[;�E�jWZy���� ���@Ѕ<U�"Qu����B9R��S����ӂۻ�[<��T3�*�dn=�YOW���`�� �3����L-��"P���sQ��7��۪=%��b��{e*�1�JM��׹�)��7�b3���¥�>6"�H�җ��5s���&3��y(��x���鞝��y��/j�	���V!�t_�vSlË�p���<3�Jg��S�o+6�k6��&���*�>�
n�U����N��^naF�N��^qu�Y1���$�)��t��������{ӑkp���W�מ�}~w"kU��m���F1v9OE먪z��8\諵R���� ���Q�N�n�{L>���y�cy�7��^o\�;{��i�tН{���عѼ�m�q�7�iBf>��-�}w�Iz"���]v6��_��u�N���i���@��"5����컣��#n�qg:�9S<u��}]�d<g�|_���q%��p�n�(66F]�ɕ��#[�Zb�U5��{�9@�(Yj��n5���jjP�Ƨ��JE���c���00�/~��7(ߓ����%�Q}�͂�v�݌)��Ń�_D��I�WTcU����ddPM/ڕ$N-W.;b֬�Ty�V�i���z鑸�l��y�6��]�>'����u���Vx��z�xU+�k)�R\8�	D';�s�.��,����5Vo
�(�RXө��n8��ݽՏ�9��_(�e5�Ě���ьP\p-􆋕��ģ��u@���ʑ%�
������BY9�����c�%�$1�HY��I�~�_)5���q���?�����g��2���%��ڤ␩Uؗ+"�'L��tK�{|d�PΘP�!��uu�{���.�m~�.�f4z��v��|GI{T�B�y��xJZ�f������lGkw
��!iЕ:�c�XaˮLں[/~�ݕ�"xp��W6D�����z���S���<r�B�͕�i�bZ��<��ܣ�k�Ž�ٵR�=�{�'�Ѵ����wNޮV�����m��|)�n��`���Pїt�i��ц�V1\�3��ٻ����d6>�9�K��g#�t��;�Y�fI�I�9��⯌�nk���j�ԍncj�,�!u3�a֑�2��`t�Zׂ�p�Q��~2�F��%��
�eg�m�����r�g]`�fG?\�l��9�+���7��*0X����v6�4��Bk�c�}���A%U�w�T"��ؙ�-E�����I1��*�]R����2/��z�g$߽7�j�:~�'���#�_��g
T˸�_�Ǚ��@��@��{�je\Q�^��/n��`՘��tN���8��p���z�ͪ�h{A�_,jZ贬lQ|f��ڽK&zWtxJ�Q��h�9��{������Xڨ���F�tO�zj�
�A�b��Ku�G-��U�A����c��X���r0����Y-����x�<0�k�]5�t�W�ז����e�Uh8t�.dj�������Bbdp�-�s�ئ-:F��Om�������9��Ϩ�)Y^)�~d��Do'K$�T�W�V ������:�PE�?m`�W��=G�t�IU���7ms��l}��$!y��/EQP`�h��֩X�&l-ҹ�-����D�+h��e?�^�����׵�{�}|��K�/��]\ɱ]�U��*U�rE7�u���n�%�Sˀn�ʹo��ǹ�ѣ)Sf��"<�z2�'��j]�}E[�Z$m������Y-8��Cq�Ծ��D��:ĵꙎ�]>���bE^)`�Gv��B�b8��^#��X<xZ�X���=��o�Qs�L��[B��]�V�3�����kfR=iX\k�%�y���uC�UtF�c�j��Fq�)c�ܻe����d�V�\��#{'<��z�;�p�Vz�����Z9�l�I�7�S����'�U�#e8[�,з���9d\�;p��g�������BL��U��C�k2Q��#�\d25��t���a�S�3c=n]��~�RՊ���9�=�����}"�m>�l�bK�=�y��O��\��:��NJ�e2�s��4s�5Kg�n�����P�9��ƹ&+��;��e^� �S�Uy�z	�Cױ��֮��KM\�L���3�ꨏz�u鴶�G��K��\��*͊r�<��|���}euY�l���9{R�ѓ�KL��Z~�=����٪��w�s�~�Y]hުpSq�*awwn�g5IHh�,� �R���͡th{֕:�����WvZ��Woq0���X�tu7�F���cz�a]vè����a�]q���O�^����bj��Rwd��S����ð��Ⱦ�O����'a�
�x�N������8�v'2o1��}�����f�S�K]�l��v/�\4�:�"�Γq��T�_u-�!���_�1���qhu1�fmkP��tm�e�+mo�%�j��g[7k��e*W�� ���p��?�+*��0�"�Y�J�:#o�i�޷}ъe�l툁�ˑ��؝9����R�,nN�3~��*�"1Sr'}L�fעW��e�˳�8��ŉU�o����b�y��e�����aߥ�w�>���O�*��9���o�+�c�++d�K�E`�v�c�9t0�R�5 ���y�Y�FQ����=�u�P�ڒ[:�7�5�����Ip��n5���R�`��6��"�Xi�@�<�h�ᗤ�؋�5:�JŇ�":
��>�bȌOݮ�򇼯킇�c%�7<��mz�]m�����Z������L��#�'��з��:�S��1�)/wN�u����t��m�`���_�Wz.TC��#z9R��Uie�6<�v�ײ�Ě����+���8���^&'n-���#Qӯ�V]WS�B���]e�v8�,��^h�}�7�,�-n�G'Q	ǚk�wNO_2�˨T��3l���C#7�wq�س�Wq����w�8Z��sޔ�@�bvwG�\����3Fn�|3s��&�Ԋ\2_?Z��F"��k�Gڻ~�^=j%�R����y�\c,�������vN{N.k>��6p튗d�؊�s�`9V|��̮�Ø�S8Dv��vk�T�;j����ª���3��Pì}ݘO��:��N���SĈ����7����;D\�)��5mv��sv3U���RȚ�whnaF�	�:h8��U�\1w�K	#y�faV�]�w5`U�P��r5���,u��|3|�;Y�Lz1�\��Z��X�҅�ae�j߹��yn�0fR��Nj1|�)�yN���҃cdau�왥��#���t���~ő܃�Lŋ���!ߧ.ڽk(o����8�O��FR�^m3�m�*r���<;��jz�X6t�c_+�ov��`�<z�X�q�vtPv2N)�����ǈ����Y-�᪾�'����=��*�S�Ӟ
[�L�U��+��L��'Wo��d��rY�N�Gs���X��``.�J��N;ʝ�9��lc�Y��<�}�Y�7��kcw������{̪�U�}�nmޝ�; InՀ.:pwQNq�',λ�=:�9.��M���Z6����7a/������,�2��un��C�w_Ө%݆�Mg����@n�ނ��jN��S/R|�����3�I̶i�u���㟯�����y�b�6O$Ț}I.)�S��������-�j-��%����#:�$nj��`��p7AQ6OY��1��V�J~l�-DB�ъIT->�%��EbR�s
�=�����,%����f�C'h:'p�"�t��g�^]f��� ������&3�WB`�Q��a��w9�oe4�cG�l�@�|G_%�R�Uo:�Y�t����Rc�˳��7���M��*���̣���dVz�#w��^L,�;ԉ4;�!C�z��V�Sw�-c���j�O�-��Tέ�:��(;Wҽk^_�6*XpٖR=�U�f�⚎w��{1m�!L0C.}h���֑�+�{%�a��>�R��F'+�Çc*�F�K���;֒�"#��\�Rt���,X��E�	��4K���o�ؒ��Ǚ�6*�u~銬Wy�J!C�v ^�D"�W�����w<˼�@�ހ 8)j�zGݎ�w��rۣN=0. >�NW�ʱ]so�N�W��g6e����IX�D �Y�=�d��X��I���YW0��,W$�ӳ�^��vtۉQO ��T����W]ej�6O���A�wG��<v4���2U�ÿ�(+���)3/v�.����v<�]9[��J�[��n��n��F�Ww��[�dԺ����j��7�z�7�X>������\0�����w�$߻Ut#]�x%�y�5�:J.�sS��\��\޷z����j�e��☍+\������COO9Y2^���ͳ���cYVyY-�F�Ƿmͣ��%��`���ɑ�:]P�	x���\{Ťf�9N��J)��;��a.�K��+�Jb�&���+L$���u*���d]��U���W�#f�2�y@{�v}ח��B����.��xҜA�b��,c�B����bztr��ؓ5W��J�b�5HcxKސ�9���!da�D,���e��mJ���K/w��n�L�]i<;�}�,'^mx�}H��j��񔑇~�p$����
uC��65v��k��Z���ܵ$l�0AS�r��FT�p=��H���\D"���!9`�me�<�9*ur���~�#�N��=	B�C�K.�z�ە��卵c���������9O{Ԝ�Xs7�Ǒ���G�4<
�!�y5��eoN�S�l)���ܻ�&�˸�������t�2����k�w�	S{خ�3<"��,���kJ�U��K��m�ؤ"���L|�'6��t�\��.Η��������f���H�KN����-5ˏ����F�0v㼾m�4���N�s��[��^����#g�f�Ǯ�\c�e:�q��"8�K�G4�7-P��l�P�e2�T����s+�q�S�S�ʰU��!�B�`�$�It�h�7��S	VhcN_4=G,���$���}���GF�u� m	�^�b������K�
�N��k��Y�����X-�Jn�<��O�dd���LM�6c^�{R��2tʉ,�Pn�t�ɯL#ٳx�ep��\n��(�'���MZ�_2��}I̦N�o1B(-v���\4g]ȳ�\���N~�v��,8��ٵ����p�YJ�}ZC�1�������.Kէ4W���B5�y��圁c�=Wk��F�[O��ǧ�q�s�%�#cm�*�����>�s�n���j+���\�:������-�jݟG�l/���?��3�sW�^�~0��]���zw9er��cU�,=t��Z�w�K�l	|���Z�k�91C���,{��"��fz�oK��u#4�<��PuO��K���5Kc��;��dO��֥ͪ�T8��Ӯ',���mބ0���N�i�֓������Ye��ޝ��:ؾ����),܅�#ޞV8�9���_35Z��⬊��Вi7J�Ypl1�BZ���ɐu�N�9�]E�gfڏg#����W�nR�;'j�n�'��7��Vu2���k���7p�Sp��.r�%uJ�:���u��@(}�R�`�'ٺ��E:�L����4We�8��rI����2B�2��x�N��K���yxl<C�%�6��t�;�N��C6۾J#�3�F�(���L�!��w��֘t�.w�U���[kK�)���X��s�vIX��#��S�@�]B�h\�O)WҫK˥j��~�6�xԦe*�b�Η|���z�+��q`�X�D����������P�qׯ�6!̡w�^�����3F�|����^��0ʖ���D��mK�|lEd�])qLR���l{�	us;����-H������0��ʱ��|j`>oڲCL�0�ل�#��u���J�p��^M�A	�y�\�[~��sw��LE{��&�wh�(�a6��g� �R���]dc����mf7�@T�6�p�2X�Ō�f�(���NB[�Q�sr�LvҶ�ۙv�=COR廃j���6���~į
3Y.�viA��0��vL��|���E�B������M�:o�gf(��b�֬��(G&�Ԍ�p�ܻt���[1��Aʻʴzۋ0k���b)s�2N�w8�a�T�ޛ*=I�"���]6t���uX��/; j���cT�뎇�1�Z��j�Z3�5 �y�\�9�kGdpv�%Y!*�3+SltC�ovq-m��R�V��l�3��
�4����1�W����8���ʄ��g�8V��*ܥL�|7�e�C��ɓDG�K����3j�幨ݗpb�W��ǳi�QJ3N�x#���ݎ�N���e�:��p�q�#i@f���<���v�r��뼣O�U+�Xunm��ԃ�n�@�z1l{8.2�FU�v�r�j�՞y�T.ZW(��u2|�=7(��%�Q���⃚��X5��p��]3�WR*�WHɄ-��ԓ�����;�\�θ"��{h�����Է���q��ۂ-!�L�G.:����Ü�A�
��,�G�S/��}x�t�[���\�����`Z�ɹ�eE��1��jҺ�D�	�p�k�U��'x��8at9X��4�]�TΗ�ct���ha�%�Y���
���Ą�9��0�ׇ�QC�~�fU��,6T;O�p#���p��+#[�]��Y%�0�IR�{׬t�]���q��q�\�[��w�l��	��k��V�K�J`v�)7�ܾn���G/[��D6���uJ�
��|��k�����k�':0�o%kz�g.���Q�;.�u�1�Z�����ʻ:���Z�LA�ò'.}/��������+e�6L���j���q
,�y�K��/�}����7"��Ѐ���nK��rU��K�}[0r�U�4t�o]Hh ��=}+�So��5tл9;�x�
�^7���;�)�}��d�2n=�>q`tK������zcJ����ǯ�=�,W����ī��n��*v���
z3���D��ӯ
S/9�Z�N�J�eqw���y�}�s�;z��voK�`��ai��Ɂ����Q]6�[��Mj��od�S���؃��,���b��(��X��t�b�t�Z�S̫�W�]�y�i�=K�'�c&���κ/;��ܫ�)�zy���"�W�V�����$������V��������n�է3��RY�-���܃*S���zbg��u�:����VU�8q���OQ�%y�����_�֎�|��N�	[m�v�2�fM����l��\x�/6|:�W ��bG��Հ��2]�M�׸:�+)6�k'dQ6mu�I���L��vz����j��iHz�l��C4Л\���-]|�%&k�ت<䇥jǪ/�7��%Ѧ��
j�uY�N�%���.�AXE�Z/�����8��R��AW��5n� �9�,�)�8�������Vn��Y�Mv����,G���|Α�S7�E�͸뻧
f�&����ľ��{���޾�|؇��Dc��aPUQZ�b �Q`�HZQ�U��b ��Ŵ�V.R�D�*���ˉ�Q���F
��S2� �&�Pb�b+A��b$Q2�Y��X��"�̵�e��Ŷ����,WV��f��EU2�F��V�PUEB,*(T�QZ��"9F��Tm����A5(��)Z[*���GYLVZ��،JڕE���2Պ��-�#Rګ�E��""F��EUuGX�:�UF"e�R�B�DF���5bԪ�4�����Uf������e��M4PC�J�AE�h,Ai(��"�Q�mau��Kh����Er�EDAQPfZ�[X�ň5QLJ1U}|n��}�/���D�v�(�c��+�G&���P�ߠP.�V�Fȡ#4E�7l�0�]�~G�sl�Q�����ou�쾑t�]�*��~ֲ0Wu�vyv��5���f���My`#)H�f�>�YǊ����X�2�e���'M/R�)��l��r�P/��+ȍ��~�g7+��y��Z���&ݭ������������uR�ӁC+b���#p;�-��lI��K��y���8��͉f54�D0�H���ˋ�BqJ��=VBp�=n�e��7����XGE�d�K%ƹAK��댚��BM�����-�aC���ģ�
�UF�7�U�ɫ*�C�t�u@���rY���8��+���bE������֥;GD8����Bb�`��Q���ic���D,$N�_%��`R�=JR��.Q�N�̃}ӫI^�q��<���6'�4�pEkʃ���QDJ !�F��V`ޢ2�ru��^���R��`B�e�:���]��m�Ȫr�t;B�%��k�G��λ�����y��y]�kc�W\K�����{<3�`?J���Zח��԰ῌ���@�o����Q���m.�V�7�}	ް%�j��_o5{u�v����:N¬��5K�N��+��Yަ�kL;���+l��G�Y���:i�V����Z�=�㐛����:�Ҕ���/�K��S,�i����l�a1𮐑�ӞoZ��Ds5���x�I�J��F��lБQ��Y��9+������)�$bj�����
�ٕ��Ȏ��dD�W��q�J�.�5��	����*�]R�T���z"������^���f���}���!�
��s�"\)��bǙuy��H�.�e��o���|' f�-�(��A��hp،5�im����yt߅1G��{$��Dgof���="�2�аq�=@���bÌ+b-��'�=f�`�7�Oo���=3N-���{���c:�#yP�_P�S���J"��#��:_F�:^T��g��+�woF�u�y�d-���f��S�4�2d#�����x�/_�g���k ��1Ď�I�������U��ں��1q�}R#�G�mh�U����.��dv�Cs�.m.Ё����s�ǾF�gǖ�\�"�xT�^���<y��I{�1W�;��q`� ��,���V�Y�ߺ]�5(�UaТ9"��>o�`�|Mٙj��!�-��Xx���K��5��5����:No�W��)�>�;�PSyd�N]f]�s`�[״aQ��v)�n���/��ڑ���A�������P��E���}WQ��t��`'����vP�9,��v��[w�#�{�[A�}u����@�s�J���`s󡥛R���!f��ø���	<B���-���ܲ/R��Mc\P�*�"�e�k�Y����od�L�=��/�*�����FT`�^HK��ܓA|hև�e��>��K��p�f�*����v6�+2���z�p��ə�� ޜq񡌞>�xN;���V���l�k�vmg�ՆytW���RУ�y�z���k֛�z���T{YS{��#�ϗ���Ixk����a��zpJ����Z�\��:���]xa�<�a��P�bz�H?�ƹ&�h�߆���P���җj}���%eW'mĪ�dӍ����M(ٕ�o�B`F��^�Xz�R�Q�~0g�&�����{�yCi��X쁏�w�)9����ߤ5�]8cTa�j~�=�[�@�ͼ�MtI<Y}�`:����ߖ�Z�c60K��aw��<y�[WM�RvB�`�ġP�T^6��4�i䛎�{;�+2�kZ������(h�G�X��˒<q��y*��PL�c׋���t�X�w�-�C�j1]�B�+)VbN�_�T�<���[�Jyݼ������sՄ��{����aލ=�(tU{×8�퀺X��p��*���c <���r�=[�y����n��L����]���p5a�Pg�����VO�@;t�Vyo����V>ŦDlm�.����V�%�y�	=����:�,҅�Vb�	+���嬥�� �E������<�7��Būd�����=Yg(�]vw������$n�y�M�|���KZz������)�=�7;OA���yjt9	eō���T�6:]6j��;�wPw�4a�L�C�����[U���w�/��!0���S�*:/��AC�fԺF�1>���b(睇�ѝH���M;����4����Ih�����Z<:�C���؄�(g�X�$
�̄c*:"f�җ���j��!�N��1u9���a�y�mh0����dC����)��ιr�I����Z��i�E}q�W%��W��u���,��~���Ey"1ʨ�m�N�&�6�A�:㚜"����yq�Ո�� ��T�܉����3[���i�x�&���rT��W��Ug��K�Ӟ-�lK�seݒ���H�sb�0솪��0�ܓ*��oR7Q�9�o��}j�浽x	���[����:�
G�SZ�g�l�yJ��o�}˭���U�B���,��N=�L�e�Dt�6u��MI�1u;X̛��֎U�Y�9�p�f�O�9��'��c�u�0��[���|��D/��Y9����y�ՒgE���X��Ck�Z7-j�&���̋���o���ϑ��i
ƣr��v3e�I�ިC�o�ܔ�h�##�\�׬�MS���K�2͏�GO��C4|v�R�4]���qC�oGI?��0���
�
=YC����6?uN����}����\�t&i����
Q�2%�`a{���X���oH�OOdv�5�Đ��?iY=Zv>b�{��>�7��/�0TG�z�׍�c~��\5�،�.���,�+Z�<����Xkz����ښ�t66�#��g&�mjՋk�(��8-�2�OX�q�QO23 WZwc��c��h	z�ѝ�L{��r�vu�=v�V��𮐁�}(��D';�p�Kc2�:�}|O��ʶ���F��1L���3i5�i�H�Q0>�Ib��HŌR�o�>�Kc#����<R��R�z��]^�ň+޻��JҾ��f'��tz娃C��,b�Py��?y���e\����q>��'FFǥ໒w%l�;�K-sO�h�]��*�i�՚~U{��Y�ͶB�H��� �8�����j��Hs�]('o�J��K4�gu�*ue�%:�B����jI�M�o���g��W�I�m\��;;�!E+�ܢ��a�y��b��X:ic�)�	��Kqy��:�ؗ(�v���Z��y�P�]��UY	�tK�[��&[�xY�Ƽ�=z���T��Cƍ8c�e�2oz�1��|�+�m@��`���ǧ{1��~�ܮO����������L�A	˺�ʽv�kΙ��=>B����׮j�ҙվ�ZE ����r�6�Z�l߄����o{hK�K���mW�UiK�w.(5�)�C��Y�{%�`�7��q`ث���W��X�o�	��?���?�$��#C?��O�`B��N6l�lÎ,�����,�4��Y�t�*X"�y�`4��N��&"�z��'�p�ˑp�<�j�m^�V�ىd�sT�l�w�bk�BPKf%��h	1ر�J������T9��"�����2w;�{�ή��p��΢���X�jW<�����8��j6��P�X~^�>{w��a�z��a�ݪ�D�+��1�LF�z!c�G��Á�V���u".��|_r��k-m��-Z�x�!�Q�a	},�x����rn��vk�nd�ܡ��:>=�{i��;Q��4�.M���5�ط���˚���ew\�&6��C�o��>gu�w#%�w=ܕ�������.qT2��#�Z�3�������a׳�����'�̌�nY�{T��di1����cqz/$�Grɂ��vC�Jע��;�Ǩ9����n�ݠ����]Nt�z��%� ?��>��R�ޕ/�o�G�������\}A��^Q�����@V�t��iZ.���H��B[��N���LĂ���+^�*�v�y:�s0�H^�+zp��꫸P68��_��}J�Ko��Y,m-<=���w�$�,S��Oب�I��ʇԎ1�Pt�=)i_ˍp-.#�)���+���<���7�L����\
J��߉Yҋ��d�Bڨ)�޹���z���F��b��z�]����_t��֣
�	C$X�-��5o-0��w��E�)2���I�0�w�q-�1�PaA�sԼ��C�V(/_>4<�CfS�vl���v�q�i��������8�`I��/��wR�0TE	s�X��hU��B�)x��~˿!�j����r��+NX���ەj0ǹ�M_��i.�-s��5�k Us�=b���!)&Ufy}�!wJ��Y���Nt�9Bþo�.�S���ٝcq�}Ϟ���J]*��kΨ��W��z�g^.�m8��g0�����#΋�WoF���4e��
m�����w*t���j�\қ�\9�y8���e���=C�z�sC��}fS�$5�F�u�dCa{	a�m#ڣ4�Y
OYS��y�3�fm_^R7��U�����⍂�-�X���KL�~FЁ��k�{��:����:�;�*ɓ���Z�90�t	��(Erv������̣M�TKYJ��Bvd�DQT��e�ٚ��<�6���H}�0���EVz���M����\��e�4x��6f�G�R�E�ǥǡ�O�Y���A�I�Bo��{��֪��"��\�z�v3��g��V	��	V~K�¡_7�.bg��ġ�>��m+��,�W��b5=��犷N���-���ݔ�F���wk+���|z��`�~��w?;[�!���lg	EŁ�u�T�6:]-�Y�S=��2�єwr�(�pC�����zfR�ҕ��
a�S�=����ʇ(�1>�n�F��\.���:W9^�P���xN$�<�i
�Iv�Ə�/��;����e|E�si�P&��(-���=�덽��ċ���]K�7:�����F���k6��C�T{��
��+qAWWW{�:�p�f������Q�K��i�9�⡼�/� �F���+$ۗ}/�n�r�{��u�Kc9��x"ޤblUЪT�j33V�_B ̣C,���)��Q�Qk֪��2:�Tr��wŐ�{8k7�bA�˸lj0�YY"kb$e��/W%����X%p��s�Y�a9��=�3�t����3k�1F~��p������WY��
��E�Y����=�����w�޹����TE���U�⪬�.�N�QC�K�|n+$��K��[��c��G�ݮ=٭��@����<k��KS����S�v7ڲCL谡�e6!���ֳC%��{���G�xWB����Qܭ���IW���o/
w���y9Q��%ً�u��v�G�2<`��S=}D�D:�gθ����őC{��O��am{=ޭ��*�P��vg,�u�"���죑��n��YeB����x8_د�`_7y�+����QYB�]�Lu�u���כd� ��]��uڰg=t�#nіY��t�fS&��/kAQ�L�u���r�]m�c����֮��Cv3����,�Ʌק!|�{zRu)'�s��6��v_\ʯ%+1�DR�H^j`˸�qC#l�#�PS�VX�^Jv,�Û[S��u GV�':�o@[k2�6���I��F�Y3&<<a�K�$%}�s��:WC���S'��}}�iE��wo�%K}ٕ���ݭGz��v�_z��)�8�uP��c-��ut(e23֝����ۉ]�R+�O$2{�oQ�NA������a��$O�� o�%�)uL��t�e������ss(K;G���j�
G����ῤ���«K�3E�M ��&�	H��Y��H|��LQ�&���/�[�WV�>r��¼|*��%��.LiG���s��H��]Nĸ���F��Z��ܲ�D���_�/��{z�t�ǯ�L�XH��[�ȭ=�.��uD�	Rz%V�j�ic��#0j�][��&�M��;�tV��=~�v���p9�Xf)�=RKu����4g�U������镜�O�>Y�rۥ�X-�7~�p�c�D��(Sy;\Y)pĲ���2T.�KQzD3��{KU������=(;]����ȳ�κk�9�9�8Y�@׸�J���t�x�v}lБQ���qx�+��������2�������,aBy�yPc5����6����H�jWLUx��1c\^8��x���ļ;�vh���>1�@2�oq�8�u>-��'��m��(8븥f��GW�]>	W.�a�ާm��>n��0�v�y�F���j�Y����#�eh`uj�V�U����Ʒ��}��ä�'VՄ��i^V���1L���]����]��h���8���F��w	i�K7����W]�Lป���|7���U�Q�	W�̙P��m��^�f�ڐ�]\�����o6Ern�j�K��k"	ۀoK�}J�Yu�����j�AF�$b��9n^�7M��⋢�Q����ɰ�+Ayl�M
ә����ъ_�;t�)=�/o&�w$��1S/��eta����)��Y�S��S����4���" T�xS��S��)݅��%N��W���[�wLq<�b�`I�v��|���|5�:����g	��;wn���7jR:*o	����D��ͣy�����o�W^un%٭D��՛6��I}3i:劜��B�7Yx�Y��\y�֥�;�Lm�ҿw:V���I�A�ћ2�Ah:=�N��1@�CZ��n믊��+�W<G{k�U�uym\h14�Z���B�V���ڈ��^�U�γ��K\���i��v�-.T�7��{���}{�bD���.�Ym�,j�rj�\��84�/t�X�"ĝGj8s)�َ�S�[�,�|��m�����	�mX�u�HK�[vC�w&f �;sJߓ�f얯%.�i���Ѭ]��gG�ٺն�A}����-�=��Z���3t����wŴ�B�w�h��͢6bB��rg4+Hq�Op�>���k#�0� :�w#�����Jv�MҒփh�����E��v:��F���ݙ�2��<�|�ɷ׋Z�9-k��0��ot���Nܷ�8��X�J�Ѵ��������z�a�սR�d*�H1m{Fu��@���P=+r���`�3��I��o,��|D �y��0�^q��	)Ú,��wU��]����#��&`��/Oz款�۶sY�{;4��5ݪ;@��j<F��+7����A�y�ɷ[L��q� %�c�tlu��a;�;�w]��h���,�.:�r�{5�������v�@��G�j��ո����+H�#S���d��.�{��4xj�sju^����ם�\���b<���qu�3*�Z.�t'%����tc��Uԭ
Y��]��J>���i�6��/	��\�N�O�*8`N����&f^!�y�.�>�+�p5@�Jh̳�x ;5�0�L7���hK����e�o���^����m
w(��ೱ�^m<9�N���3�Iɺ�f�w���ĺOs�̹f4�g�NFe�eJ�+�݈�7�������6�,�;B��s)�I�� �7B�	� 5�A��r�ͥ����u)�H&����\}~/�e��iU���<��46��QE@B��U�)Z�e��S-�Rթ�b���Ya����PF1S
و`1DAc,DX�e���YlV"����(+P�QJ�b����Qb���*̵�
��,F(�%�b�H��2X���R�U���X5*�*"����,�`�%"��#TF*��D1Eb�UULj,����TF*���EQ���lU���1X��a\�VEEbE�*9s%V1U��Q��UQQ�6�4U
�dV"�h�3)1�2"�*��e(�FH�(��ZEdkDUJ����kE��Zշ�*��D������ZJ��mˑ�Q��ls,Ϯ~ۻ�k�G��Cv��{;Cg8�;�s�pǨ��h���+��P6�5����;+mc)��C�x�]y����]ۃs{0�6o�U��S`4����<mD	�z˥�	�Vˑpjg�
�^���،��v�I�|�MyHj	�ٔIi#y��i4=�+�1^�s~W�㧺�f'ǧ�m���5h��;�
�����bÌ+b-��1�Г�nDˋ�[K�Q׸b�.�l'~��95y�5��<�(P���,�#M-t�/�=�F<^�W
�)仜t���d�l�����ߦF8�[�ofX;�!
�Ukڝ��{ǉ�U�]i��Bc�75�s0�9�ύ��XX�1:�*���)�a��'K$�T�[�CNj�GGLԼN�X4�z�=���0<uǰ+��`���j/V���|�Bܿ�K��+�t{(��؇�T������(��Fk��!���vxԣ�U�B��H��-͵��+����)b��H/˧b(g	e�Zr0�ж��ٲ��b�O�O��\�Ҳ�L�T�L�di$a����%��a���jڨ4���	�G��p�����.���n����͑\9/���=2	��W�^Ǘ �,$��j!�Y6��3������\�=m�ќ�\��x�Q��$t�٩��H��p텻�NA�q��@�\y�<V�$�s;�T��qܕ�R�ք�\��i�^���zӖgp�2��������c�
R���ܦ/r��޺5������4s[�6)'s�6.��N>��D�:3A������1Q�J��\��z�:�o��X�]�a($����9Ƨ<Z�OW4(�*2Kz�2��"8���t�/E@s8M�%.�O#��
��K5�y�����YA�-�;�DkA��B�B����c|k�u��W�Xp�aၼ�-Ǳ��߸�=\huMz�T�UC+�sJ�̭�a�gi�Q�^�Xz��3�GQ���c�����=�y6�[����x?�c�c�nzR/vH��c^�{U��N���a�Y�/�쩝ؕ��<�t���+&���ʰ�����f�h1�';�ޗ�l���8ʞ�bS�:=�*�,�wQk0����t)�p��֠65N�C���{��ʈ�؉��Wi<w~�W���R�J��3����5N4�\�z�ѓ�U��M��a�zSs���,ݞ��#Oq�ު݌N{L���-b>��Q�P��4N�鞉���凨)���!�%-��~���q�Ŵa!_��ev�������8�F�)��@e�vK�P|Eg�?tż�I<E�O��j{y¢Z{��NKKf�u)���Or����@x=ɘ���#L�a�Mu�.������Q�T��U��W��+Q�X[-���.�;���Y��t��� O0i�;��ɍ�X��'���8�+{<�|�Sǥ�Dzoi�c4K*/h"�ʩ�lt�[WȾ��	=��V�0w]���u7�<�:gJbeT+�ĄE	bD������Ѡv�Q}���H��'׃s��:�i\�a^n������e��4�Q
	G|y%��搭iv�Z<:�q��؁��ojibU��ըU��y�@�_Q����tX�0W�<�ft-U~�p+�ʓv1`�b��y �7/ȁOԟ���ɞ�V���Ll�E��_ڹ-����D���O;n*�"��<�Cg3U��'�U�~�Z]�|��m_�u�W�# ��*�b�K%���w*-�ʔ��[���B(�D�Xr��'�~��#xgl):
�8�׷�<�pQ]�*R�����Y
�nR����|�!�|�j�!�t\2ξ��k�M��}κz�(:����8�k>��c�hm[�yQJ���%^�,��uH����k{b���9�mX�-�w�
���#�@��r��)��Fq��p�BI����6;�v*���'S��WH{�n��	�s{���]H��3�/ZOz�e�
�1������E�O"��4\�F(M-�u��F�t��sk�%�C�a�i�=˳Lzp�{5���G��[#�Pª2�h��L�,O��D�^V�&n���y�ء/بp4�r"���C�m���� X���"c�v��>�7\2fFϟF�f�|�!3������
��Zc�45�X�YQ���7���b�^n�q���2�����#��Z��{4~6�
�t�F��֮ܑ�����Y��ؠ����d�f��e������mt�y;bN�ȸ��z{��XtyC��G���;�yތ|�ۓXYU~�U� X�̿'f�Y��UC�1pP����\\���v�t�[cVEc���ԳԈ���Oy�,M�Y�T��>GG��O�SP�ʾ^	[�g6^�cӎ��u<��eS�^0�$���f+�L�+����<����\�g	p��i��FQ}�m�,�R/��<��I��N�>��bt�Iߖ4A'{�^L���	]X�<k�ʙ��D����M�o�i��.[.�썠~��/�m�M��+��vt޼H�R����w�����k�]^�fU���w+�k�>~5���e��������꼉ʚ��x
�禈T����C'N���		�'nkȳ�����F>�{�d��od�/;.N�������ҙJ�]{\N�s]�]��da���7���L�(^1o��1X^���O���̣���dV[�n��k����v4����p�x��,�/�P8)o禇;�5Z�8w�V�҃��y��:�}����st5��z�����`z��K�b��u&������qz��
Z��C:u���3U�.���3���15(�C�Ki'ґ��Z):K�:,X�Qx�%�2��i�Us+uT�\?\a��T����i�£lA줔<ZQi��W��C�˴p��ۑVf܎׽^0��y�����"�t6ek�L��X옸
�Od$�ޗwt٫y�f�+v�½�4��h�ť=��Q~��jV'�##�(�]�K��'�.zx�4� �I,�[5nz��#�
/�c���;宔F����{w�~V�@��-5��)�*8��GQͫ��T;��,^���!
�UQz���P+���t�M�fꢺ*�(�ky��)�h��a�f����)r�_����O�J���6�Wv)�{zuԴ����kB����7j�dk�i97D�8f�m�ZI2��bVgpi�,�����s_�=�:��y�W��x�:ܼ���lN	�+L�ԇ���t�ڶI��-Z�q�Ǎ\Vfik�j�����]5b�����Ŏ���Ù�w]rr��Z��dͧ�j�L��K��{�^^�i��2���\�f�:v���8[�K���e��%��E�t�P���Z����:���#Ƅ�}����YA�u�{a�o%�7�VпO��|]�D��C�Li����K�G5�[��%��q��]={K�+�=����K#I#5@�c�ҫ�(�Y{�]��z�뒜W8�h�p��˵�y'�m�ޏ����,z� ~�#�0xhth֎Q�kZ��0��c}ѥ�����*I���yR�}Uu��qz������]�g���8�A�yD���!���"�f0��}�1o���K�vr~�A���>޿i�6��bLI����|��\}P�{6�{s*���u�t���>�'�6V)~���Y�C��e� �e���t5䘩\|�������)��b�yS�Ȅj����RU�W���Ӓz��덲!����NŉuꖹFG^0���0�u_��F���͌D��~�I�;�Dׁ͘r��};;p�f�*S���qn�f�
°��c8Y4���]�:g�=0�s[�>+7%G�Żl҉�[�*;�$�����s��(���?��z1iهn߱ky�V���[���7�+���[����y�����1um�۹���U��J]��G8��1T	G��$p��ݚڛ4j����ht�{)�Kǳk�]��Y��h<��%��Aoz\Ք����c�S�7�9����nF ����!�G�Ӌ����3���
�̍3U:7�g��cEM�~J���.K��3��:��B� ^Tԩ����p�c-c�qx����������¯����F����4')E���ӷ0�daP��:�WE�ɫ�yz�WuZ��:͖��J/�;���Y=t���i�����6�S��u���lG}ܵ�k�n�5���t���(�����T�ΗC�ۧ��S=��:�zT�"�.��W,r���	�'�EV�t��/�q�.��ǌ�x>>��+��a{�}W��6M���i��Q��w�K��C<�?�ѧ3<\��&WK�qj
�.�1RB\��������p�J��E~��Ot��>Du0xo�'���c�%[3is��4�ޏ������^� )���e��9p���+����wp��׫��B�e����F��㹡J6�@:�y�+߻3g;�3*�����Ӷ��Kk���C�n�͸�i��ڔ9G]��+s�X欭<�Tב8�ԗ6��P�}�/im�/�,�^n�[����:#u5�y���3����NñtM�v�=�|��N���ŏ���ri�o�Y<)�z��R�ҏ�Յ�'���s^+F20A�5�I�#f_lh�m���ոVB~�(������U����^�����KZpȞ��B�	wd��ٻY5�⧡����Hx�LR�\�9d*��KV����TC|U]������sAF�N�������N�܀p��ᢲ<3�e3�_�2WL�7y���P�,����BNr{�x�׎?`O�Υ�);���i)�,
�\�˃����9|��������l�V�v���Us�{���T,IK���Z����=��KD�'^��o׃��2b�d���s�׳��⇃٧Q�s�f���$7r�Ƶ1�^םbmeFC(�3��j�pip��/c]�}R�/h���LucP{5x�kU������Xb�F�jxh�g�G7}{��Bz�Ո_)>Z���R��@�#!^u�_���iE��J#Wn��J��-�=A1����ml�����d��0�SԩS�]A�5g�G�`y˸D@�=v���~=}\�T=����/{�U���Ų��wrwa�x��f�cln��#tQ~�����z*�p{�7�'�F&�j��_NG))��mu���rE���϶�����}��.Fv�PW]��klr��e��:�����߬����vH
��wX��qg��g�aU��3�.��!bu3W�#�WpTm+�U��įyVz�us-]���ͼ�4U;�B_�}Pb�$A`�	G=D��9v�5��3��I밡�1��c����<{ݫK|31-N�֪�tgW+�O�r�F�7�=���-�f���g�FF0mon�Se-�dm>�%�W�����P��K��u�|�lSj���vnF��sq<��g����� G����5�(k8���]�5�ن �K��R��8���T�M���r���V�v@�}�:�,]�0N�#�,��eOcNpCv�:�TL�Q�V�<�n)�7&<��Xy3ӧ������B|����z�e�+	|:�䘹�w�^N�qA�v��Oj�X��f��kr����+�N���o@�Mn.p�=2��IR,���٧KidQ8����t��;#�,ڒ����$]ħ[���Vm��;�ǈt����t�Ԣ�q�QD^}�p��̜�z�������E�հ�ZO����]�ܺ�L��L"��N�5H�@�\�{˗S��s�7�"�6e�n�M1{��.��=�zky ,|���t-м=����z����a��KC�\���Y-_�%�{�ƭh�J�DZ�u'���yt�k��O�KkQ�T�Y���s�2P�ƅeZs��V��u<���Ճj���F�7���k��m��S�F�P��E75҅�uٜ̎t�V�>�ot��?9u���z�㥙�V֙�p�}s��ފȸ�n72�l�k^��3A'#��:�R�������=��ƨ���sJ���L�b�r�7��?J"�2/�F�[�O��C�x�ͽx�܋˼w���冺^f�H=��~�1�c��_��G����p�Ps�t���N��-�����ۛ~�Pރvμ��lhw�Gd>�<��x�O�L#�����b
:Z�t������ػ]GDD��O�k��y��H@��	!I����$��	!IHIO�H@�hB���IO�BH@��	!I�D$�	'�@�$����$�	!IHIO�I HN��I!�`IO�H@�XB��@�$����$��$�	'�$�	'�����)������\��8(���1%�|�@� �z�JH� J��  � �@ h I 
 Ҁ(*� ( P( V�[aR�i f�T��J	)5��mF=��`#M���֪��4(IR	R�ƪ*�dݵJJ��ƣ-��)-�*BB[JT�;��EB��kh�U%M��XV��l��V�H��ʐ�kID�B��R*��IE�;%,m�DJ�RjQ
��UIv��J��Y�   ��%Mh���)*�˹ݭ�b�M�*�"��R�ʦT��k5(k0��UpH;r�����h�UA��#R��S�A%D��   O[hR��33l�LR5+[a�&)�
R��ɫm(�i�jSZ%�[e�-�MV���S@h�mfR�(+oM\(�ܔ�6f���ZiJҵ%�n   .�
(P�B�:��
B� P�����B�CB��z�� 
B��;�
(P�AEr���
 �B�
�(P�B�TA٦����v5J�0�D����u�le��SfZh���   q�����R���-�,Ԕ5�T�X����Ҧ��J7]8iB�������l��4Ԩ;u*�����X�lԕ�JRm�T�0k$+�  ��I�B��J�)R�f�TD�mݤU(v���H�CkL�X��)gG8�PU��ҫ�CCc��T��
(im���k4�f%[@J��JO   燠	5��Z�MIf�����Ф˹�V�T7g:��P6�ʕIUvư�Jҭ�֜��*��ʌ5�m�SZ�U���]�cV�D��[ZUx  '��,[*�jT�U��ҥI�m��
N��u��IRgk�����-Q��XZ5  �����[V��Z�RJ���-�Y(� � Ś
�hV���@�V@6���*eU� 7���M�`P1ݸ 
CW[a��M�(�Z-��ʣ�  n�� wW (t�Li� L� l����0 :.���4�,V�Lm5w9 �9d��iYi�T(�  ���&րc�W�WU�
0�b��& �AF����S*�2-��Z�$��M��S�*P)�IRP�OѓU �  ���)P  �	�0ѓL�H���H  b~?����?~`����?F��Ks�-��n�vwNQ����
��ސ���{�������$���BC�`IO�$ I?�	!H�B!!���ǿ�C����~����Q�[���:�i��mS)�v�vc���ɞ�ySG�X��-|kF�x��j�೷zս�Xq��~f�.�I�h"Z�����*�	�%Zu&V�tԬ��Cb�s74gƶ�ݴ�V�-�d�G2,��N<��jùYJ�����[b}!�-!��.�¨5�vy�pi4���*2�f��ely���2ؚ�p�R��6^3V.a���!�3oQǒeK��+4�d�����$e��Bu�CJf
T2��k~�f���:p毵c�y2�k$�ᆳ&���.�I� �hn㠕me���0[�ٶ�g�h��P��q,��H�ir٢\��KT����Q ����+Tǖ��tv9%�R��v��Y0#�)�z���0S�j�X:��,`43���]��{oOv���81�������i^�6�6����Q���أ����{@jX�ŪK(5�D�c盆�*�U\T���托�=�3U�/!q'f���"ղ�-�Ң-�*�P�Զ�k	U�W[b��oQ[�e�]�E�8��&�F��I<�EZ�ϖ��#Wg1ش�DTJUilQ͂hm���"քߗ�R�`�k�5��{Cc������NZ��(���ś�r��6̷f��<2�iGi��Z6�x�e��D{���B�{�a4$�M��j^�ٶH�(Zݣ�\�I�L�mER�5�U�@ȧͷwq�[��Ӷ��3of!cNFf��5B�ٻ]eh�I)S@j�����
#lMa��� Y�g,����.R[m�X���;/ܬ��ʌ7`���n�7��]՛�S[�L�.VIo�U=8��t!��E;̫���3-������g� �B��\A5��A���"r�z�+a�+*h��l඄7�AK�'����k��:7E��"Ф���,n�[z�h�-��@��X�N7��P;͂��t����/A�Rf�6�̪b�eC�+&:��2+Х�f�Z�̦n�VlYV��ƞb���9r��I
�2fEy�^ZWdMSD�.���6�b�.���d�Z5f��gz���J'I����-��.�)��.S[+N*E�@2�(���押�%��ˢǘ�`-")ɨ������ó��m�.�,V�����|)Ȓ�a��7��5"�ó��Jl�õ��B�w��-��.ZՊQ��n+�*��Y�3q�������D�BL�rPn��e��M�oT��ۼ�M �r)v=���X�$ �b��4��th��{w�
���Y����?���:4����tjv����ffk�Z8�U'̻�y�n�s5�'	�l�"%�[5-��0K��O5���&nr蚺�i���T|��Uؖ��޷���-��գ���q������j�a3sa7���b��&ۥ3n�z^���YQ�@��b$0��q:�k5�Xھ�z�R�T�.�t�B��k��`���l��*�S)��v|�@��z�?�0�"f�Ɔ4���3+3�ޭmb�5͂�w,�I�ř�NH$����.� 33C��Lh��VVd���F���Ќ��-�n�ZZ�Zn��T��f�u�F�Y2�\w)��N	��k4�%kZ�]6�fkCsZ���R,���wSM��ݺʆD�_&�K	&U�ym��sM0�� HV�f���;�yQXxhL���*���AY��l�[�.��n�J*�e�B�E�8h�;F�0��Q=�;�;��'V M�\2�D�n�G�(�Zh��&\��{/t��+���U��[E��DB�2H2J-�ݻ��)��R63a��n�ѹzJۨcѕ�meZO$H��J�gw>�2ɭl3/׺�&����iÒ	x��
�/ᮯ6	�������W�ϲ�B�Ȍh��ST��0��� 6c�yX�[Z�-3N3���+a��R�X&!1�}�jTfn��w��Pu�{vn�����c�Y�K�7BV0��ښd�t��`m�L�7�!Zȹ���$u7ve4�����fV���h�5�t-Ƿ(4��+��a�u+�[�"5�m�=t+�a`vo���t ���ԕ�f�*�R���1[l��6#�M���]�ǘ�Ξ�uc��2����ϬاW��j׽mrZ4�x��6��Kw(悬e���[y���ڻ�0ZWK[$uw��-���|j��o��E�6��d�DĨ�iJ���V���Eَ��Ȥs&ܻ��`�����	��9 JÈڽ�F�gXq
x6�4���Mb�J��2�'P˔�FK"� ��3v���L���oP��`5�l.���%� a,4��7�jaks4ؖ����E�f�:Ҙ�TH�m5��b�[1Ym�8(�k-�5�F��-.'���[施<`�t{;��a�tH���y(;��0�B�� B�U]�I�Ŷ��,�ǛQAy���rn�b�0(`X�B���ՔU�6�g�@ü �,[�c��}��� ��u.�7���7��%��n����a��fiE��/q�X TŶ�~Bc�z�Ñ��,*��2��N����Ve�����n���n,��L\Ɠ�P�8��]�J�����i�.�9u�=��:Y����K��иr��C�K�xE�Kچ�2㸩�fӋ1୔��h��,ӻK�7i͗X�#{��gn����m��u��ZlH�-P�o5l����-�h%5�&��y���7d=5*Qv��ԓl�,�����%[�&K�w�ʂ�^ѻ$6�@�z�4�L�&n�T�h+4��0j��摗I�C݌�ysAY{wl#���`��WYD�X�;N	Gr��܌D����Qк�oo5*��34o*k��I�[����Z��f�wzt�j���S@�|��F������2��Lص�u��7P�=@Q���4*�hT�!96l*�؂
���2���9h��9m�b	�ޤi�  ������$��gq�8��z���n�M�^抓ۑB��EL3vʤ�LW]�J�\�C��n�vW��9S.(H��.n���(A%��%��0����hlyp �f���6��gp1Ł�sj;���Y��Y-�UC�mc��]\��]E�y�,#7]���&V�2��=;��74�<��`�-S*��ɏa�fl�.�a�و�̩Xe�rbĬ�6Rٻ� uqN(����[�{��)��)��Z�;�eѱW)��U��\�0<ߪ,U��6��
軋7L��F�'m�;��.�b �����ݡ���0��b����^��1P�SB����u#��ꔙ�A�d�ݼջL�ML�Yz�FM��6���ȫJ����D-�����]-,�ǯU�t[v̂�e��%���@m�B�ټS۵A��sV�t�%��D1�o5̧D�nD+��;���Z��)���zr�6uⵕm=L��[[��C;�Ώ�� ��#�]-�,�P�Գ�x�Rjʘ�w���IŘ)^�͘�"��w��JQ�7d���Z.�&���s0l�Ú�e��QVA���F�Ub�pU��f-뱇�nZsJY-�C�"n�M�i����c%i¶+��*ϲ�n��;�bK�lB�S�j57w)�(�WHÐ�jh&#*S�6~�]Ӈh��}�<.ŕ,�F��35�-m])y�Ġ�3L�e���"�6/�i�v��ꭏp�CpL�N���Ie2�P�a�'�+4:�'�od���EL�m�uޑfڼ��;X�)VU�� 2���4���1Y{H��hQ�(�Y�:w�̴2Dw�Pj�R��Y��M�����]��f���R�pG�t���b/�A|6ڼ H�㒎7"WͫSnXk#��2=�w��-P���Qb�Pݱ.X�P䉹�v��r��
2�Aܦ�#u�(T��ӎ�1m��g&���6	[��j�<�1D�B��Ն/\� ���J��_�of3z���}��G.����sM^VX��гWw��բ�]���1]�`��Ր�p5��e2­e֚�`. f������ �2�S�1�^21�,�+�:���!5qj��74<�-٭�j�����p"v�Zl+��A$�E�[�[��R���p��B�[z��K��U-me�j-muu6��4d`fnU��Y,d'�jiw`e֕�^M{����ի̕om�;�`jYQ�d�O&V�{4�c2�,�E���&��w3��
:����+Ӗ�֣��A��u�5�Tz�������yw�a=q,�hC�[7�Yw@��¾��$�^a�l��Jf[y��������7�^k1kn<f�jct	Y$F�	B��#����ues\IoK"�nTx z�u�0ް��2�W�u �(^	YH�����*�Th��w]�}��.<�r��y���v�Ų�8n�.�	qų���L�͠�1Z��V�!4�UC�ʗtn]^�ӳ��C�C�jM�u��gwRr!���P��
�e�X�.F-R�*�J�0V�%)���{z�a(6j2���S6jY�$ܼu�r�J�Ӆ	`��Z��ө�nZx�Fv�U�r��#��G�zb �L_ayF0��E�⭑m
N�a
�v�kZk3�(����w��ç���69��u�����v��� ;l���!���/��[��4�!�����h5�%��sP�Nj�q�!��֛ԩ�+&�\˫�I��4���b�7ҥ�W��n�5���{���׬�`���,,�T�S+�[���k�*��ƪ����7&)�n�ren�R���*i3M�T��72�
���m�m�#s�1شfn6pI@)�Q��q1�ѩ�$����&%��t˳b�d�m��.1���bq7)�/Yd�rf�d��t��������˫�߮�0[[[�����8�t�V��50P֊L,� ٶ[��h˱�Tܬ-fSr����F\#2�p��|wG�麒{ɗ��wX�Fm���,�ƶ�z̠�]L��(�%Gj�VEi��G(�=vCkV=�:AXsqi��e8��fP�]nm<��V-m(0��d[��D�2(��hܻ����(�J]�k����.�������4�9��cj��	a��y4�P4� �:�b���]�׉&U�bQ��*b��:MnU���|kf�����emړfr�ۊ@6�v�P!ʔ)m�RUiJU��%#U� �!I�j�A���.����%:ӏ^��8��naI5������eeh���F��n�*���e��V[��!ݖd6� .�;�m�� �A��S#��(ۋw7)�(� �кvk�&-��5�)V����^*�X��E8�Ĳ,Wb�a�ӤT�.e�k:������"���-�8/YĆ��u-gF�f�Yc�uo+J545RQ�c ��Ya�7~��Ĭ�)Xiڼ�j����l�Y�QיFʽזE�w��nd�V�C$����(�XsR�`h���⫀�B3XwY�v-6�:ڊ�їw�y�mD�i9V(��e%�V>���u5�'P�⽛����kB$���Ȭ^e.푙���YL+�F<z6�hK.<1��᥵�g����4�Sr�n����U�bj���-���tŮ��p9o��c��V37.�5͚ὃ	:�b@n�K�w�%�cJٓ�H2�ݷ��r"7]��̪UنiW��v�
4YlL���"Yr�g"{����he
��у0m��V+���&�ʻ+t��X�Q%����F�V7u�8���^VP˶h�@M�)��*�ɽ�X
�{���#�ؗN�7M�����S1�+���ֱK*�^-R̳���6X�P�1I6c�B���S5Y�ݪgl�MͫJ/mb��FfEwWs���-�ˬqR��.���nU��`U� *�8Uf!>���[f�����UǬlrT�-��yh� �c"߳h�պ�=��Y�j*��+�#Wj�7�A�wa��6fI�j�ڳ���qj�0	s>;\�r�˦2��d�o+^H����)��6��ԠՃ(-�إ�`$��1�w	�ڼ۰���h�l�A���� �Eb�#��6�a$��jɽ�X�]��k���h�����l:�-��v����zT����CfYYH;�b�%�{�Z�U�@ۡy�k!�XR�E��M�k� ��ip�]t�����-8�yicZk�^�x�W�"�ո�lkH)�YH�cz��r��Y-�WD��Yʎ�Ubg�Z-0�W"L�ܑ�[�
�o�ˢ�n��-Em�	�t�i"�e蛦��xb5f�JD�l���$������u���V��Wst��_Zx��	�1[K��T*ʬ�Z�Y��Fc`��q(���vv�fʽߕ��uOwMͻֱ�"W�c�N}�5��H��ޖ�2�Z��t��)#���B��֊�-Ji�'c ��"���teE����Zfʊmڭw6Ve��E'&�Ň#�r�@��NB-n��In�a���f�m)ͻr�E���D���:�&K����l�!�
�s"��nC�LbR�,�K�y�s�`7W���މM�9J����h������@CP�3aC0�{e���Y)��(�#&��������Y�$0լ�b����M	���l�EE���p����2+(ՅS�bͩc[2��9�Y�܏,��N��7f�/�e[,S�4�Ul4HE���ǆ?��Yz�,	�@AX�9l`��kJLv�����ڃ+XG-�8K`�m�4f%�d�t۸��YP`�����=��ҷ�o����W�"�Ǜ����L��$�Pƍ���*�^����c���Iϒ���v�2���md\�p��<ǽ/w��1{�h:Uej���~ª�o��6����h6����]>�([�b��q'��tz�s�Sn��M����]t/;�l=�գhdLzy�Ed���Εv�CYżr���Ǹ�4(؛e�냡�;t��\6p�,q��q�Ә��d���gL�޸����W�_BUv��gE%فµ+�F+O�0	Q!�\w�ӎ�=�fi�=j�l]u��~B4�����ae��C
�DMQT��&�]�#���}����l��ڔyr�*�8�%���EJ�9h�
�kB;��oik4ǽ8����M�����H�'�q����N��P.���M��h,�MdzFI��;.�ġ�!c/NG�E�|)��ۼ����q�)a��
�p�R�+TY]N���IZat��R�yi�_��[���ë;�Q2���WP%B�fƪ��5�	_r�(�|ƍ5��f*@�k�'3�Q��(UTB?�,X��Lv�5IЧ�Bq�&�ݞ�t'B��}&�Q5vb<�s��-9HF�]p?;�6�]gb茬 ]�4�J�r��)N`�K*� Vͼ[��X�T��N��ɠ8��<7۱����fӓ>�pQΨ��]\��P��O`dLZ��}�^��ȯi���X����,ӱ��&�PV�u��L�����#��X�s��F.���6^���yzd�İO-�F%�9g5��[{E�gM�t���2m8ܙ��x؆����<�KU��\:�Pi(�\����2�i�.U#�.��m�t;�a���*�2�]�*<��� �t��#�z�S�'-�6Um�}�̕��v�U�KaZ�\ZA7Z��q>��ȸ6:WHQ��&�é��lvu)w"R�FN{w5���y	Ȕ��&�6�n�:����VԴˀ^l�W5P�΄��ؗ'�K#F�m���cDN�Bы���+z�u�8JQ��l�s����U���;��3u�,*|�3�(b7�h$���w����_?h��Β�aζg��z�0ӎ��j�D_+0Lo0۠� /v5���kr�>��_Q�ĭ�ibɁt��Mʳ�'P�	������٫�ܻF��u��֍fw>����+GQO��S�b�ƺm�ɵM5.����腒�lf�aj��Y�6��m������L
��\�V:������+0A�����QCwc�0+ICX�����r���,���+��˗����V���(�<\{efl�[����JU;��M���:h�̧K��J<�&҂O������ù����*�hnv�j�)I�t̼����Re��ٌ�=$�+��N�"l�Y+i����C������M����L���<
eq�5�fɒY�ȱ���|Q��[o�&�{�0��ؐ�b�@��J�]	�S��I�޺��V���5Y/�Ņf�6X��ȫ�z��Zt��b�P��l&j`����d��h�M�{
��HV�<�i���&�ň�6-�e��к��,k�u����ݧ�Ś_�4��^���£�ej��2��9������q���v(�,uh��J<�1�woY1��(좛�ru��
�b���(��L{���yо�[�5���nq�$GxR��2�۵���q�$�TOA�]��P,�Mp�f];T��gG7j��Ͱ"7�@p���k3�Lj�b%���3\@=�`�g�[�|��ɜ����
�z�l�$�y@1��C�f ��I��WՌfb2�'���R�3C���u�fӸ�ó^c�u��;P���Ԇ��1r˥|äaT��4i��!N��<W �㶡̕cN��Ns�ﺇ8p�7!:�#[�˷�*��QZZ1T`'d���ւ�}}{Y��Vk7�Թ�u]�9��EJe���f,�����eiX��������X����>�Kt��w�I%��3%-����ՓR��BU�tޮ��+o�
��hZK��\V����f�H��k���B�]�.���8L�(�7Ru�s� ��]�bQ�#wJUt���/��B�����E���<��)tG+�e%}7%�o]���O�y�X�<7F�Zs8\��.�W4��/39e���D�w}��� �Pչ�ھ��yw4���8��9k�P)f|Ʈ�"c�Fo>+����Xk;����*�n�2��פ�+dfЅ��at�F�<�]�l�Y�y�T3rb<]#v/ Գ1Қ�n�R ���B��@S�u3��Z�g3xv��+�+q�k7S8��[R���/�Q=d��� �٬t���l���eA�8CN����˨̺�g��_L��zې{RC=۬�C��� Ք���3��p�
��R�_>���Kp�.�#�:�%S�:ɩ����C�-I�!�	J����.-R���_4�7��ñ��s��h�\�;�W՜t�ۦcG�K/�I��i��������a��Z�ɷʞ�&"�m���ZxW�eۈ�L�)'rꕂ�Yu���v��3y<�f��NCK>e��:���-�����Us��V�n�ZX�8�:���"4��v�	�Rh4��jM��3�"�`r���&�;��������0��'����
��*� ���P؂Z	��d(1aWջ͢!Ʌ���y�n^Zh�n�R�z�6c8��Y��Y��hv&���@���z�p"����tpYS�#����6�山����8��K#����b�=5�qQ
�&�Mo�gCR1�zH�IJ&����)`oN^:x̯��5��8����"�-gմ^���nef-�*�Х	�����f�V�**�c]s�8+�N�e&�-��H�p�|k�h�Ge�2PK\Y������>�;'$�cd�vr9����+v��l3��У����r�V+�;tqs6c/�E��Sq4�C���e�'n���������bZ����Tw���w��wxJnsT�ڊ���7:�Ղ(j�n+_u��bк�1j��Z�\��+r���Ԗ�
YW�	Aeb�@�n/.g*�w.]*���8�e[���1���r��D��y���Bj7��.�Y[z��/���Qز�e9r���s�奼)W=�6cY*`g6�g�ΤNn�5���3����0���I��c�8+��IG0�m�g�|,�R�X4cz3\/��[��6���s��x*:����c�;���y�A]Ω�3'L3D���^�Q�e�ӧ����ݥ6�]�J6�Z`A!�Ou�cK��y.��g�.�^��L��I��0���[�C(.�ݥQ��*Ɏ�5�H���mM9�k���9x�)w=����ä6%-T���%
��b����u�%Df-\��R�e{38������R;rU��s��^<�k�YV6)��,��d�����r�̳�lsuj�MڃTz�v��K���ĲDՂ��F�K�<�7�vPI�f�eDfk ��W/fVQ�S��.ەvB�xz�:E��5`�@��%Z��AW�i��6}��e�2�!Z�ϰ��ʹ��Cm���w���[KhҿiC�Q6��� � x�qۆ���n+a�.��tV�][�\�1Ҷ�7�sz8�]|'.�AM�;A�fؗ�㦂]�6>L��݉��09��|
��P>��1d�K*ػA�1�d�A��S�IN����ao�WZ:�jWݍ�M�R��z_�qݗ��JtKn�r��Y[f�J������ګ&�tBok2�7Q����+]R��v��m��2e��v���ׂ�]N²��k!��y�H�]@���}3�ݫZ���ݦ�kUմfk�F�s�/��b����\��f���Ԗ+37��Y�6�w6�ͺS�ȗn���x���Vw�Y� ��\�Q�0NC�1-u�bɉ<�CF&��n��	��w(�r�Y;}�\�X�i5Is���;s*ڼ{%kYXhf\�iI��?^��2V��/k#s�rb�g].�c5�,{)��s��C\��;ԟπP�T��\��ٯ��^��d#��U�$�a"��rGLqwP|jZQ�i������l|'wU�(�\�̻Bs�;��P�+�]כr����mc`���E��UŐ��n>���G����q[bu���rp���n
Ja��B�9	��r�=�V�S/��iqsuf�V��s	��g��Cy�g�]+�\
�7m`�@�o��;n^��:R�83���a��e�4l�wg5\�M������=Q�>�[����-�.���Y���=^�B���MZ�Gμ@��$�n��WWB�ɚ�?"�0`/�a�-ų��d=;<�M���k(Z�Au*�-�qx/�HE�[�5�:�	j5	���|ZVo�x�59��ʁ�Y��+��ۃH�CJsr�������+li5�v��0&H�+z)�����\��W/�
`2�h�s���ch�[��J�Ү��t���h�,�Yz��;(�<lf!+�;�ƊK�/��@W&����b�+P?a�79��J�7JJD�O�idn�%�w��*��T���6P��Y-�1��Y{��5��O��ok�1)2�������Wa;��Hf�Д�[RJ���5�sC]z� ��A��<��(ә� ��"b�s\�����NJ�mJٙ��i	^���Gfs���W؟[n�`��vwm��F9�X�c�x��3��FP�e�>Sy��,ܝ
�Dm:� �p�/h[Q�WK�:L��݃�k'�v�d�𙽢��*K�f����v�Y�m!�;Pf�Lel�ư�_0��t�wۗdm�����g��S�q܃5>�Y�-
.�����;F�l�i�B4T�r�ZX|[ �S7����8q;#�����[�k�D=�̹-��'F&pl���o�f�Ԝ�LY��[7��з�9��j����"p�����dr�"���l9���*Vc�F�H�%�l��'\�{YY�
R�' �����"���>��p-��r,��1ū�o-����3 _T��Lx��b]�>˛.䥚�*�&Х;��H���k�h����m���7����v�.wÎ���2&Ɗ'J|�?N͜釽��|Y��/4<��JE�ȝ���'\!gWdl�E[sc���Χ��M�ϲ�F�;�'��ڑ��Uu�ŬD��-�CMn�;���!},�<7}��ň*t��"I/ƞއzɼo_^��5N�4�]{��81ܚīx��+4��!0�.��熛��;�T�^ڻ�eذք3A�MY�a���c�6���*Y�
��	����
��jL)��+6�T��hW
���Ӧ���p�ݩ-�]��N�Wf���&���a-6N-k��ʴ/)�+�B�ܔlk}�(��8r��� ��Fb�-v�����OI��$�����_22��:d��A�5��,;����p�vn͠^�xjVM;���Ć�,�w}y�%v�Z��8��k~eo'x��n{����v(�<v,ނ&4�)3��&��f)����wO��7]S���:L��DU��*_%V �V}����	f�Z��\��!W7���2�!e�z�pIZ���sikV�3����p��I��@Y��".���Ղ<�˒P�
�٭>��m�6
�<M�zc���Jt�H�fWV�*��!ÜQ�0��
���E�i��E(m�&)��"k��m��Vل�j���CtCi���*�>޹����SXaj�{Y5��8�
�'q��,��K�[m����T wW2�/��\�n�`���]̽�X���L���ޥ^��J�3G�V�s|�A��@�����G�)G��Yq�gT����ȹ��aA݁M߲���G�!uk���$=艷>���&�`ں��rAB^�}$Nk��'Y�r�>5!� `�J�d��+��3�N��ֻ�����3���d��O�=�jܔ��&
W;˙��j�X�*�̍F>ױ"+h�9���6�s�#��>x�'��2̘�E�(T���U*�
�S%b@fX6�.8�5�:��v&��˧�eu�6��w�}n��G�hٶ;4ߧ�8RV�T�x ����cU=79��qRl�V/��V�����p�{ubR�S����C�9i�k��8������U�N���f��Q��CW[NM̝����Wj���'-`�p�NN��T�a5�0���0�k5��욗e��O�G�]\����Y!V�vk�C%u���%��P���F�� w��̄�\�+F���1/.k��5>7c�h9���yѣ͗b�c�K�;K��nA��Eb����E��p�:pM�.�Nc+3�s]6�'Aj�R��&,
��d��t�R��홻�G� �xO�,^��&�d��t6�u�ÃW�s6oS���Q�v��P�[�>�^<,��_c�9��N�t�;�ݝE�,
��
�J�m6��V�d�mh�G,p�VY�̊�.�	�
o�_e]�Z�+c����~�d��x�v�[[o*@y;55rY�R����`C�vJ� ��V�f�"f]�h3��zX�
u�{rgA��N�j��Rk�-�_CVj^�u���4�wq�&p�N���ۙ��\���dr�4n2��	u#XgW:���1�α�Dj�3�B�i�I#ڬ�+���F6C"�a���g�٤VRvc��%�q�ԏ,.����3|"�Ue��dNoTŐgP���,u��M���[mҼ�gL2��Z���[%<��
�zzgR��cv��ڧ��N���c2�i-�wy\�v-�%2k�}����=���{���k�8�=�~�z�e�Wfh 4���۸�`��E)�U�ۯmed&���.�G0�h�����v�0��'I'Q���*�TU:�v�d��{w�j��H���;�DN;b��2���*ʙO�1�q�`E�[��z�Y��f�s)��s��� t�r|p^Y��n�0'����(q���ip���ld�!&`U�5�݊�� j��W��Y�
�mm�((�u�.��c����0z�"yyP��I�Hbc��A�X)ѹ��^�8AiLt�8k@}��nYP��[����Ŭ��7*�:�b�mf;m�������sPxL����.��`C�5I^�ל�gN����;����;n����ˡ����X�p�asƅ��M��m��i
����6p��L�oM1T��f�WmK��r.�fm�q�Z3��i����T�U�}Z�oS�<{dc���*�)�qh�z��R�txgrG�1gA2�8e]�{yл�zh��1�R�j�R�6M�g��28{�3.Q�ԚI�h�r��=y{��7!b�t�;4��"z4U(C���vkZ�FP�i��_-$f=z+0%�s6�r��+V<6He���$z��bu7�]`��%Y+�-c[yA��b��}1u�������Q�Y�r���S<ʔ�M���R����j5���]
���5��^e��f�F�X��њ��fd*�ɦ�fC��f��O(��>�3������Y���L�7�Jp�̤�Zq�	-�M_G\����3�^V����5SÕm��6���#Q�m؝-]Szv��k�zT�5b�&]��(��b�v�k"�۾����NϕOLDz�ʐ^Գ�h�>J��Ze�z�i��p[m
[3�'��t�B�]i���+��5Im���<Lh��,%ݫu6�����u���u�����8�`��کc�,�q+�Y�P\��i���]��Ef�]b��)��ҷ��k��m6*�-�q@_[�5K���tNv��m���b����P�]�$��sf}I�9�v1���_D[[7i��ݛ�#Q5��h0b�-�ⶆHk�ցy|�P��ޥB�&��������67�/��]ucU��B�c[��*m�@l07"��qm$���e����:��Ǣ��9M)��n犻Ws=�SQեؤ>��񠐒�(�}�H����q�n�����\���Әn�}�y4@0�{�b�t\붅A*��x����w���m���Ue�Ğ��K��f��H�_P���y���&���q]�^�0>�L]�=ۼY�]"���|3r�t�41�(�v��Y����%Cs7�IܵRU����fӵ8�в��CFrO�3(���s��1I�I]���ࣗ�;�ۥݢ<d��4�MZ�zXɲ�N����	�����n���˾T�.��9n���Qk\��C/ǵ���i0��w��n$�+�!v�n%
�oZ�5]9˖Xj�y�gx.�����f�0q�wרU�)�������6h�:;>�
��o5�n�]�SE����v)�vSw+TJ	�W����aMe�w�Q$��b;l���S��(� ��b�5ӓIeN��5B�L�fTw,�P��茝���g��˭Z��.��� &ڡ����۸�"���G�V�C
��
Ƒmš^�`aݛ��݄mp�t]*�$�ؽ΢P��m��9��a�	���sL�I�Z����ej�K]!R��=֫v�J���|���eu�D��e��9������t�b�&%=�6me�ٕ2p����Z�;2�0��J�t�����4<�`MZt�Ê�"���~��'�h����*-�\�A��")�>1�Wu�K�����.��osX%VQ^���v��;�m(ICu���Q�_ni"󖰷E9��a��X31��.����Ѻ�][iTrd�9ڦ_]'j�u��>�ܩռ���1���驽X�U��}�]^�L�ڇ>X@��I]�P�Nˮ���	����[k �8��V�ܐ�(�
�8�\;|B%��s�����λE��/��x ZR���k��"^����* ą��p��o)�'�v��5��Vt�ڝ�C#�گu��˳�7a�di��$��do'm�pI���uĥ����
0:�y�5���Ի��8j���Da4	�����26�-����ҖN�g� u��sј�S`*���J��Z��xv�Fr�˹M��Av�/z9�v7��fP�E-��6ٗK4:�u��lնˊ>���v��[�!FW%��J�Wnں�I���(�l�V[��ڽ����<C2�F�EyZG�3v�ZN�d�}y�_�Ct������4��`��U�B�+zN�g �eLwݻʃ����V�}V�B���8Mִ��OMv�wL_(:�{����k�n���`x����ַx���ݵ׭�b\\�W8d��L�����cs2[1y��cf¬D�K<�]�\�=d�	A��-�붜�԰o��H����4�ږ�ԕ-�u�6�j�|���ɇr���I'lV$��r���P�82��h}5F�zɭ�!��d&=U���`���/[�ΑR���lc]�.�#��@o��Ż��T�i�vZͷ�PP��� )yf��S�F�q�z�<��y�-���ID��f��К5�X-eҮ�db�Esw��TiԺ���8^:g`��9u�kjƓ���<�����x)�7+u���,��^�+sW�0�������l�M�A)me<ʐ����v�)�>T��Lp4�^6W%�� @Y�ɮ�̻vࣼkMc.el�4� us�w�a@�]��j}c#}S\��K����i�悆�} ���@����]��=1�ƴ6�Y��p\L\-�UV�����-A\���4���D_(֕��/.8^sˌe7v�Uu��`Uc锏���������)�C��kC:�<Wb�q\�;q���!��=�~�X	�R�	x�����>w��
YLrx��9f2�^�y fiέy�u��d)
��e�H��}�^k�H;kճ�{�9Q�圩��tC����1�X�YyO��v���
�qf���D"�#і��6^�5[\�
�(��^5wu��g�`�ʵ��Ǖ*]\Xt�uƌ���ɦ�f�MVc�X���3�֜ fgT�(��Esyf� }Υ�.�1��Ԕ�%�� թ(Ѵ�����I�%�*�)�Z/l�.�.�լ{VTr�e����Sv��ϟmF2�ט�,�e�>�k*�*\\�.�@ܶ��j6/SP����QP�ܹZ�P�u�w����0ou;�3'Zz]=�.v�����}ǲ����S/`Y����ږ�)`ԠAnvp�otX麵Q����r�K����О]�EZ´�\3��qTA����k�����Ƴ3{P��c�0���-�ۥ�y�.�T4 ��6�fY��)�@���m��飀b�:�ge75]v��u�MB��M�ǥ*+��+��lUL��B��Ͼ�f����ݜ�K��dTj�n���絀tJ��f�&^�e�A1G���|f?���RG�с���ق��Q=��Z�N���=n;�ic�f�����&��Z��t�}����DBpu�mU�0t�Wז��1�4��t�R@�
#��0)B���V�M*��K-�MX�q͵wpS�O	ߏ������j���,5�{�U�zG��Ctw���w�=!�ݸC��]j����:p�z�ne�1pw�A�:�n���9q���i���mcA���PǬ�"½*�V}�v�)��[��P{�>ۺOh;��n��V�b����3Xp�X,���`V��mċ�aP�*���na�5�h�L*Q�w�V�řv�Yf�v��r�
��qg>�i�@�qf|��]K��u�1X� ���t����Pۑ�em���Fݘ����ۺ����*��rO����Je�e(�U��讦�h����[�NG��L�Ԁ���O�Y�ĩ��I��@�i���c��:ǅ*Z��W�\wW�XUNɼw��$mc�[���(�l)��qfI�����ikMEJ�������K6QХ�͆���V��$|�t��U'x�J�b�� M��0�U�Co�މ�t�ev�����jr|I�2�e�&;��zs��] �W ��P�5�_^����y*&�v�-���|������fV����+Uu;EđvK*T<"#�n�5e�v�6�2�w)V���f}�j�:���tRv�خ�qx�\����򅁪�#A�Lu���Y��1������l�l�����f�\+���'�dQ��3�҅y�w�x���VAR�����˛]ָ�r�x�E���Q���\!a`F�jV��$VVh4!�Ll��}_*��ч�[zt��b��Z�dn5��zչ�E|�E����_Y���S��K�&PW]�B��tӕzt�4�����Ԩ�\���Б�=2`�{�(l"7n5�m��T{�e�0��1��I��U�����w�G��"O%�`u�O���p��оvaQ�,����l�ٍɏr���	�-�<mˇC�e;t��xZ,���))x�eЪ�.�hا��s�:� y4Pⶱ��zp�]D�%3.����f�LX��΢�rD*��*[����	�+o�C��0�
�9������Z��/4J�F@L�.����3�A��L������J��/;Ų���J��B�u��
�(��+��]�z�7�=�e)´�Ò+�i5{��,�'�Y+��h�D�G��:��ڎmEʰ-q�\j����幹��4$��MQ��r��44u�TYj�W��s4�khD&�^*P�[�n>7C]���B���-Y�|em�ë/���6�Rv�C�Թ,WO��w{Ϸ\]ktUΰe.�J�sJ�=���ծ�c�7 �2¡��L�Q�Ȼ��]2���q%�4���N�e^�JMҶ���̺�f���f�5�����uGʹ���K��v�)�4aD�a'*�\7�Y�j��#p���9|�

TN�\�ְ^H��̋ԋ�.D���.q����<;4�S��"��0�qF��-��iub��L�jV�B�J�wa4�9;��X�q`�ut*����l�L�\�@��b�^<
��
��5q�V��vVh�)-�6MD�PD�F�����	y��Xピ�^��M�Օ �[��!�9���[WS]���beI��͎P�i��{�1wT����ζ%���i�����ŵ-���!jY��Թ0��}1��u5;�k�)�������.���Z�V�Z�f�o":k!��#!��AX�4�.�m�J�P�3x�҃�l[u��m"����)z��_-�cA�/`&��5th;��<�b�^�s��@`5.?7��!�3��
T�m�� �l�pt�+��dʸ���g8�Q�&"◎Ħ��@ب��5��o�/8i+ʼ�&�!xHP��C��X��>}�PIi��@��|��#Me(0+��r��zP���;{W�����kF�f��d5f���;닺SY��� ������x >	�V&w'��d�+8ۨ��(�/�˧�$pEV�]{���r�t�4�v��Y�1W;��wd"�JƑ�9�M]��wN�w���W�M'[�+=°���w�ը�{xn�6�f�є�R������X�}C�K�eP�&����v�}�Z��EY7�}u|�L���υ��C��;z�D�f�6�A�t������W�R�qU��r[� Jk8�9���Y뼼��f�l�� E� ��f�o$r�#�|�q�ȃ��t1�V0w��[_]j���5��@Q�������X�ͬ�ahe�%%�&ej�ˌn�OS����B�l%�l<{ջ6�%��/�M]Ƙv��cz;��{�oV��w��X�B�"�gM���{m��ST���y�kb�4��>���W����+�M��r���Jj�t�/6򥤬��Ҏ�7��Рۘ�$uS;�+�F���*H��]p^[�E�#�-�X��+�v�T"a����dڦ�n�1�U�j��u���t@��8@���`4�7�6�����g{��ll�ILV�L�`�k��5��l��^L�.�G_
n���9�*�[�M����#�Ը��P�6���A�5�[�򒠯y镶Şf�CM�1;wǐ�fŴ#�7��Z2�G"�=�XB�H\�$��-Ԭ�U�m!ӯ.\s6s3*)���B�UٻB�5�[���;��쭼B	����_[��iҵ7�*+�������X�u�f��k(�`�YT�f�ڽlb�/�;�!��s�����PV2_\i�+n��,b#!;�ޓj�乆g��M1�Ӈ��qe��n�޷�� ��y�q˸��]g�w��b�f�M')���OVS�;h7�H7\vÀƔ�T))�0�Z4��=�چw��qUoa��n!}���7�+ֽi�R���%�&.�ޠ)s{BP�j�ٴأ�B��VWU�@倧'�:��%d�F�d�:��_k<o��Ox�X�t�Ie-�q�v��C�`7���:��8�)�kb����^IK���7�:oʎ����� �����N�뛡��@���ib�Y���K�Y+��d*���EJ��
�r��mi=�+��ڬ�B8ή#��e^ُ)�Ǵ(�b�>d��#����嫵��re
g.��:��:���L1Q��q���nj�6T�8&�J�>a�3s���p\�c�്ۗO�M�9� u�.�ˊ��{�o��{��{ޱ�z��!<Xa��Q�D�M�ԫ�`�����gEfPU�rvG�5�u��$ƻ�"`��N��̛Kn���b�q��I�-v�4қ��=5��'K�p�l�n>!Y��*Y�\f�ؔ6fTP���%�C+`� ��J�C�]�v�<'��J&�a�i��, ��U��3v�;��S7��3Q�Ѷ�s+�ǅ�D��J�Ԋ�*ba�vne^ֆ�S�1Ӯ��`��2�r�d"�&��d�v� ����.�#���4o�Kq���~܄�*��
��_63��$*���5O�kf�U�3s�^����g �VZ�Ww��t�E ;��Iu2��:r%�^ǒ�XxNSJﶮ�6E�M:Zeer1rŔ5�\w��VP9i֑ƈu��}�:4�@h�M(����sO���)�enԹt-,��.�kU�q]X�]�1k��`�t�1����F��Z��4Y�΂[[*�:�p�소Kܼw[���e��V�����-�'\wX��0̆d�14쮶;p;U�蹒rr5I�.��Gh%��|�GxSjfX}�t���-��<5��Jt��w)
6�座k�<�Vi'���o�>ȐvqZS&_m��C��J��bC[D�꼫Qe/��[V�����ÖL���m�_g�U�����:A�:	�s�l��С�$A4@KYF,��j[
5-�)e���Z5�T�kXƲ����j(�([ZV�mJ���)hUDcmQ�ZV�R֢[[k)Dj��l��#JZU��bډD�����!mk�J�A�"�����(ĩY[*ڥ��aYe�"ZUQ���lQ�-�5��+�Rҫ�U�V�U[mJ��"*�ZX��"��Km�k*����Ub�ѕ�6��EQ�X���6�UR�m�l���Z5������1�ؖ�j%,-*�YZ�U��E���X�E��A�Kխ�Rڊ֣F�T����6U�ōZX�l�b�QF-j�kX(�Ĉ��mV�cJ��F�¢
*0d�m�,-�TBڰQb#lR�5��U-�Tej��EE*�Z���meTP`���l������A���A`���h���e�`����iA�bŖ��UPTEb�R[b)XVQ���ւ�U�( ����e�������������}0�IŨ�/lV�p�hb[�o���P��s��Xv� r��8�oS{���:밋k��E�Z�mP��:p�F8��T0}֯��q�&�C8���#-f�	J!��{X����Vx..����$���>pX�t@�9�W�Q��Iu�ƶk0g<�i��v����˹���j\	�ӂ�<���J�*El�X���AAΊ�nD`Q���-'K�Xط��E���d8G���;f�M_Շ�G�0�2���$4���ޟ��M��K�{ӧ������H����8����˅r�ĺ�2Zf��^�04����`�G2}h�S�˒I��QR�x�6�ǈ͎!E������w0O�,G��ň��5�
�t6V]��`��TK�:��S�m߰R�Gp��7�PE��ƣnG)�pl����lB��õy��q��FM�]+;����.fA#������}�Wh�X�e���m	�U����5u,먋��]tO9қ�����-�Y��l'c*H��`�s�9 ������ꛝ��
\�8&n�pˇ�b��p�m�EBa�>��M�͓�h������E&m�Qu8d��������*��u�B�-�a��3�o�?��n'f�0V��*�#%c���*MAU.Cg��R��_h���2����0���y}�[ )��3�������'<���] 33��#[sy:V�1YN�m��U���]Zj=��7; P8�W`�Qt�ORSR��E���y.�ǌN�锭��Ez�ꔬk�T�j~5���0�N��Jjؑ�4F챕E��6|]�Br����^}~�1S�˱�0�oV7oy��va�QBn�B�됣��,�X&b����;q�:�N	U�K���ׯg1�e�s{b��.��Q|���ȡ+|��~�5<e�Wg� �{��{ ^��+�ʶ-�>�����!Gl�a��>C�A�: D ��D��j,b�:*�>};cq�Pym���F%��B�5�Ι�@�{*��qu!@��AVJ�H.H�^�<uI��9�mL�M�*j7k�dT0s��r�����;ʺ��v�����:5\"�Ha�Y�ӊYJ��A�ke2Ƣ���#i��'e�B�(V��`S;��L�&�ŅN���
�Y�"^�c�m�R����\��~�����x"�j�v+d���q�)�[�tN���!��6�Y$��s��������U�ª-^
�p�b8��j����t���xr*'��%lEd֜��wE����wr��mCzV4�6�-�ݬ��9�M.����X�9A��
'�M;*pV�]�9I��gr�{�-�М�bPsi��ru)��yd��Z��f�sSd�c��8��T:����N�nuĔU�q�\[g'��{�e�ݫ�"%�� ԟ4+�\+\�*NHV*�2���v��y��
�E1;O�K��D��";��1kǷ�s�f�"!#��9GEa*ϼP�YWq��T���sw�o��QҹeGl�����L���S�_b;�����Է��;������
���R�}\�<��`q-N�F�B�yȭ�
A�1aG3��.76�e��Spy�ˉ��ib��^����b��] a��u�o�e���oÿYb���2l�=,g,�3�i��Eqt�K=�և.����u�z��x;��s�
t��{:�JP��s���P�IOt�04��Q�8E9�R*��[�z2��\6k���pg�)��u	2���ײH�x���r��qB��#¸V�T�Ǯ��%��S+��)�<���ӥɄ���3E`���������`5�TW�P�nO�@ٞCH���x�6�&J���\��j�1�E�3��X�X�)B�JduVyp�r����| �w�򨾈��}P�˔��C#H�'�ɚ2!�S�z(�xM�^4����,�y��,=����J��y{ƫ"miA�[����iʁN��ǐMy��>U��:����mo>�����i yq"��'{}�Gk�V��f�эQ9|��1����v�O��3�-����圈�$����c�\��g���M������Q�veG{G!�����y(���^P^�x76���J7�d�t'�3U�R��>հ���;Nw�!)��CT�N���xd��4F���89
7����)y^�j���>γQA�Q�=�gEk��&\<u�!A/s,�[�n"�D�D�O;�Tk\�}�20E�W4#J�(W@�&c'�!�0��ƸV�.6����r�^�{n��˦7�V҂搐ȇ[�!�n�ʥ�\��.�ztU�0���Ε��<��jNYm5Ko��c��Μ�T=����Ce�EE�-Ezhs��Н�(��#F�[�%j������2���U�X3�ۜ�.7C�o�V��6�^�X� ���*`"���O��{r���3�.v'gT�5��ي�Ō,��(!7������J�㣲N�j�J%`�X�aSK�����E�P�H��M��b����6�K�+��;�7]
�WVl���Y�Ϣ�37�觅4}��U�����Z�}Q^-���AO`�n	�v�j��¬TW��h��T�S|�\�c���d���}�s,�J��G/�׽u:(gP����s�{-N+�:֎)���
3V�J���}���]�>w����7�\x>�0�*1�c�����:��J=�\,��8���3s�﹞��OT�]��ӌ�O<��φ�%��T
�b>�\P��r�t��*�m����`�[��`M�~q�Y�ã�\�g���CO�Ⲻ�]��Z~W�^e;{�O��q�i��IR�X���j[L�	L��s�V���K����eD��u�ƟI��Ԅ����K�(4��|���T�1�L�����3�N�����o1�ug��rK�{����ʇ��cΒ��̨��;Ps��}(�XnmNǻ��C���(l��ն��a��g	�mmʙA@B�|~5��$������b��q�A��\���<7��~�%ir��͍���zH�*���ԟ?O9"�6T�]'±w���V��7k�%�.����Qf;%l��R�aJ�q�ɛ�j��h��Q�	}��Bˁ/eߟ�����]������p���/�;�>�
�ŉd�iъ�^p()��na� �羝*��.]�1��\�Q�7#6
/UI�؝���� ���4G����_ ��ʶ�Y�e*%�H*f���X,R9X��R7��#�W_p��u5YB�<t��B�ҫ�C[�@&m�Wp��e��Qa�
��]F��Y��z�r'�It/:�2�W��[���u���?rZfC�����m(�R�0��3Y�QY�6�'�t�l��h�#[��Ռ�/8AZ���U0!�%I	�tȗ3��4��$��q��M䘸���+��xHq���݂}�B�����&ǹV��{%9Y���r�哹K]y:>A��iQ�%�c*H1��X䊜�U�C����v��wOX����b{o'c<�HLp�aN�� ���7��Ƀu��]V�]V�b���>G�q�1B7 q�m��v��� c��mt����7�ltg��ښy[�
���*��[t_]�x�6h�����r[�!Ԩ�\��.���ڢ��S^d' �y�606��X��J^'vZ����iʮ�Tc�k�½G)��U�8 ��/��E�N� ������ј�Ύ%��l
,fڊ��^��0��G��W�P;5<e�We ~=��yRe�+B��|�Qb��y�;d+
ht�u("��Bd!�"O����Xj^m�������/4'w̏y�K�jf;�3�U~Ӌ�
@��
��`���~&��y�_�hQF5d��v����5�lw':y(�wf�5t���+�V�;I��r���Vw�x5�ng#Rf���Tp�x4��j̗bfB��2�n���Xiu㼅4�W[�{�˭a2���dO0����6	�O:�OF���׊rl��&*���W0�Va����w�VWf��M�\z,��&��yWYA�\���^Up�����19�3]�c,I�;s;t�*�:�e��t�]S=
]eϒd����U��gsPg�{y.^��
c�>�|�C��PB�r���p/Us��B��O��c�pB�
5&m�N�ޚ�����#�:D���(���玕׌����Uꩂ��tf^.�����hO��a?F��*ۂI�b��k�*NHW꫌�!�����qy/��+5���79�|�F��0�3�a��m��JZ(g�9L�_]ǃ�ؽ�V�fw���aq�y{�m�N�oԾt�b����>ړ梮�\L�g�V�"�`�M7�y��'���LZ=Pu�8�CY�[��N�9��}��Ɏ�O��+��8�'���Q��n����*�Yj��$Z>�t����		� ��G�L�͝^ȭח���n�q+0j�{�*)L���$VW\�5�U�$��-הn�.Z�E��)��bXi��KV��d)�bH6�����gq5N��ܭ)Щ|�Cp�wÍ�J|�����2�=�̾b�c�}����<�+%cgjJ�t��Kޮ��z��uxyi��{j��Ҭ�4����lZ�r,Ȳ���^!O�;&ޚ�vp����ؤ�d��
�Q�c��o�)�8/��H�=�!:����
��}ތ���vZY���v�k��=P��q�z�]�
���Ⱥµ*Y�ȡ*��>�ђט7o�����y��^ĘP�21��X)�����]�U�'�W�=��2�/�b��'�g.<�uB_aP�EO�U�E�b�-t�E��=.UeJs1�4�.N��㺠d�g=���vDx�r)�z�lM�NG�S�,W��'aA�fTX��*o���{iZD��w<��0��܊{B��*:+��}���Z ���������X.������Q�<���Ԭ�1��,�3x��쀽�=S�X���>���:'\��p�Н��9��+��U�9��	�uj�֑ �T�hE��"J�*f2qX$C��ʉ� �7$���ܜwז��v2�2�-<�Tu�=����	�bi	�u�醝�
q%
�xúX-�@���tI�{�۝!���vk(�!@�x۹�Be� L�W����Bve����Aɽ�fr�oN�e��f��6�ob�O�S'P\/Ot�Z�kmv-rxR6��G��h�m^1�X����l�J?:������k�� ���遲��XB��v1�R��(]�2�=p6V�m��S�i�����'F�d��Ԯ�[,�$fW��!���[���1����h[2�@�>K��X���,��[^�!��,�#cv�=u����2��ՎX�6Z�q�V@�3װ�m��M����]��c�F
P�H���}�\le!C7ۥǗmd&wa�fqմ�~K��{���3{S�P��e��U���T�x\K�2���^5*z��Űj�;jWV����{��W�i򾅾�s��3�������-̓�a3�uS�Mڻ��.x���,G+$u�m��l����음�$UJ�eEa�UFϲ\
�s�WC��Q����g�R��'7�\�T�j[�'a¿S*1� ����������K���>���ѷ
�(aN==
(�(�9α�������	�nU��4
SJ���S��oN�=�q�t����0�PQ�<ʋ�����W����ˑ�wU��>�|�x��������U�B��z���>8,��2�k�7<�>~偞�ǵebH]�ۮN˂@]�s�V��Uy[��l�m�Ѽ�;�t]�y����Gw�ЦM���>4���[���s�փ}��5��ZȞ\P��rY;u,�V���:.:q�X�U�5�r��/}�R�VX�c�������ug�ɩT�umr���?^��7ہ秠�R�H�:u$��$T�ʃR+��"/��ib�w]k8��y��*�0�݊Q�s�WLp��;�<�h����G�0�.R�$6[�����̞�
��YI6�k�=�;��bs��Ω�\�pw����p�\_�����f��%鬳0��t�ŷ�s���5ﭭ��{k4�7��tp�L���`���8�=�A�#M��oU\�w����=�h�|�n���������؟�wDEz�dJ����݈�V�\󅼈�2���wG��V�$�uԪ���޶����<1�pot�����-�W�; �Ϙ�� ���HLz�_���n�޺�x���X����
+�h��nD7%�ۼĖL�g]��~TpS}�n ���o͓�G&O��E3nB���uqz��`�2�hˌS�E�B��ck�a_f�}C#c�5�ښ <;�6���8[���[�����ޖLV����_�r\���b�T\�u�h2�8��m��� ��8�:���ab��H��6����JSSqh��Xi�["�r-*݆����ݻ)$�r��+�z��S^p��CN�t=HX��	�%��]F��L��Vo52O��=��w��X�$����x����g�o��ѭ��P�B��}��V���ee��LE�M�2��/��WKa�j"��5��kCTdt��+A��:'PdF�G�`�bS���,Uγ����պ���"�e�w�$��T�kh�΋��ٕ��N,obU�֓w�����5��wn�a$����[��i���Nx�v0���3��M��g*��W)Q2WI؋2���6�V8L��_D�Q4-_\.�TV��,L��b�Mr�Fj�O����kj�,��D_D�q�0i0ho4��"3 �M�}�A�u�9�YĝRef�;�ϟR��5�2W*JT���}�q.�]61�`�)�� ۜQ�l\ɿ!�_4�n*Sejc>Jȱ#n��[Z���eìsR���Ҳ���ݥF�7n�¦3�f����б>��aG�t*h]т�b|�T�+�jt��8�M�=��Ej!D����U��'��$�|�f��U�h]�z��Z���z9����o,Q<���T��6���<k�Uʼ�4�.WJ
�iʶ2��{Ho� �i�׈GdJ��k�=��Po7��82��,Xl�ww8խ�b�Z�X�B4�V#u[)E2��B� �J!��J��m������Kw<y �:��cR����P�0��udO���y�]��VwD����k*��!�sVN�劃�P2^'�6�VΧa�Ӓ�N��1r�me�+7;vAI
)f5\ SΫuf�e뾣#�,��;j�vD�	ќ�L����z�����cS���TY�&��t�)�%�KJPgo�w��:뫸�0�3�}��bM�� 2�����1^�RSMpt@�jrܣ�M*�x��:��KO�%���e�[�w^Z@�V�ŝ��*�|��㒣f�/�
��j�`����RN�g�oZ�If��f^cڶ�e�c�&�O����67��vM��O�'�X�M�e�1�\6�֞Ä�J��@���R)}��9�`R:P[�7��,Jt3ܸr�W��xQ1�flT��u-Z�sJ��yױ!�͈�T��:�z��f*I�(��z���ǱR�q��7K�֢�V�\�ѻXb�L���SRT�^�O0�ծXhb��I}�Y���W��[�5U��5~ P��y1�zoM]>z�� W��7��f�-$��ո�,��ӡ�
��s�K+�y�b���%&�Jwi�F��
���0�e6����m�T]�\�@fj�a���mn��sC�1���&tźM��m�pZ�z��*#��fˑ��G@�ݣY�(ӄ#0os�x�h��w�/Y)%c�&����}�^}�_S�v���XZ(X"�����-�TD���2ґDD[B�Z*Ŋ�QF�UYm�-B���U���m�bZUk*V�DE�@DTX�PUDҊȊ*�U�#m�ZQeJE����X������A��R(���XQ�F**�U���6�V"1U��ƥ-� ��TJՊ�QDjTX��(�"��T�[b�J6�b��DQX��U#P��APTX�E��#-�E�1�-b֨�iQX�EQD�"��,T��PQ+-�ҫ%eQ��Q�AJ�0X��(ւ���*�V+m�-������QD�Qem�[������E�P�b�A�iUF1 �� ���"*#Z"0m�eVX"��"�(�F,A�QX���"�Ċ���"�j��QdX� ������Z���*��`�U��h��A�EFb+`��"���"(�
6�DPEb"�1AUQD*T�DE ���P���Z�^�$,ˣe����
�Ef���ڸ��#B��sZ�2�v	�L�̐����L��x�N���:�\��W��[;���_yt:�5��O�H��j�~pL$(}{�um2��6���,R��0tޢ�)5�|yp��=p ��x�|�����]n����La�%��+�63�N}6��g(����͂�� _��l�aM�C��)UR���:.���+7s/ws���Ғ!E0.�	�P�KS1�c=�V�R/�G@��
��`���\�d;@��qX����.yT���No����]]�}��̫t:���v��*�F}j�Z�%G}���`�ql��4��Ϋ�nt[���]L�O�&N�Brb����y�/pR���+��ǝ48��׏x�V���j�r9�W6�k&,���������b/g���"xeter4���痆�5E+b!����� u����U��
���!\-:"��A��+Є�'$+���ϫf���m�=Ԑ�8�_{Ӻs~]B�缨�_�Ȅ|>�v�ɰј5$q
�0L��s����VT�u��{&��$E����w��M�t��+�݇�Λ]p�.��wwyT�3fM(�+,2[v���lη�}/�%��E8� �r7R*�f�=r���i��[�6�!+���rK��	E\�1�x�f�U�U�U��K�����ܵ��_GР�2�'<��0�8�zk�L�jKQWS� �_T�~�q��B�yyNbl1�н���Kh����r���Tsc���-�	�[Ŝ,�z�Z��g���	��1�(�2�˂+ko���ma�@�U��o�x�����Sb-��/�T�^�����pVx���U2��)REe;���
��:-ϔf�Fܼ�*-�u�{���d�V��I1Py
��+|��J�p_Qp�iz�K�Ƽ+���m)���5�LC�'��f�A�s�C�.�\��]
�Zh�cLJ���2�U�Q(�s�19/d�O 髁ѨO�}jz�[/"GFҫU]P�m	�����3]�+E�r:�?W2$�e@"���3�m�\]o�&�yS����fQ#���V��*�Y{�;Pw��}��mDyF@�7�]J$��܋ɵ=Ǌ��e2!ζeE�|��}�b��6�t�Ʊ�mp9��
�TtTi}��@�Z ���\��5!�?*�W#s���D�QĮ1�z���2��s��<��{���_��f��/+0���^�9K6'(ᵆ�ZO�`�S��r���®V�XU	�4�s۔`�y�S%n�e��ܱm�6ˎr��"d��k
��	͡�U��u�ҁ���R������݁�p��Y�E�g.]�9��xf�#qB²�j�1n���r�x�{*3�u�zͮE�I>ӕ���r��ݧr�}~��X���ЋD�+�T�d�H�W�` o>��������I��\��}Az��3��qq(H{�=0CL�M�K��K�]"�表G֭!����\�S�$�<����ߓ�k�����5�\�)�6X�0``j+�C�N���o�yε�=�%���
:Z� �l������Vg]�9ˍ��q哢	��Uz��ې��_uN[;IrVo �z�EAhK�mJK�;?-���T��U똽,g�-HyY�mG#Dƫ��u�X�]�@�5�KN�T���fE,�9��6��.<��ˈ{�T���P�m�z�"��ջޝ��PE�R�5�~P�X�.%����C(�̕����Oe�2��gc���p�v��u�!�8��=���>������
\�˶�Q�d�8m�p��Ᾰσ��b^I�g͜��S�]���H���ʼ5�Rh��uEzn+�^�!KK��Ż�G%����ĕ�q�)+�R��]C�1���!V�#׹u�����\�ڹ'0׻=Dx��{<ϧ4z���{�*E]̳/2�]��:�3l�o,�4����;l��w\�j�cF�����^Wsj;���ꭷ�}'�.�,�����
��VT��*�҇�`"ݧaºeF9�P؝rH9Զ⛌ȟ�O��e��xp5�k�IA�1p.\(Pl���:�/ x�w�#�sz��P�7�o�c���X�%i�+��*���'��F�
<yҍ�;Pp[9��t���1�uuh�9ֵ�6���#cɋ{b`�J�B.*������x�*..gaE���d����nZT�n�I���#�)7l�u�>���mR�4'����ǼZ#L�iq�X�A^�!L�����A������AEՁN:���ؙ�/%�ǈF)D�;	�����G�i=�sW/p�������$�Ω�T�pw����p�\\�pT���I��u��g�N-g�Zw�0���X=�U_GI޻:�u�E�vO\�n��(�2�uP��9ï��\��>��t�x>h�
���-����}j���ۑ~�S��\kw�1J/���y>�����^�f�U��M7�W�#!� �dP�G"��ptU%qGӖX��q�=Ld�]�6]d#���X�u�Ί��C]J;H!4)�-��
��k�=�]L%oh�j�XP+�g��K�V��]o_���������9%6S/{�fxy�7��>v�7S˺ �5z��`�Yk��V�_I��r�:{mv�/���쓫�������	���:=~m���^��f�I��d���VR��8)�X<�]��SE�e���;:�^Z��>�jw�0��ܣ�#����y�ף�]WU��[I�$?"��D�R�?S�x)߰-�%�����A[=�}�|F�Fk��4��AW�-.��',�u7�"�GB�ցT���S�����JxmQr��v	ȇ�FF�T�d�]�g%�f��=Yޓ3B�Wu���gR>KS�m�B��e�&b��b�j��2�Un���^��G�Zu�r]t
�	ڊ�c��$N9�4a)��n��r���cW3����b�d�@����yRU&� _��l�aM�!���^�Ey�D�K1�f)�F�m>GUڻ�.�:*�y��b�+��c��]V���ԋ
G@^��!X!,��,բ�1d��&�!�,WW��g��άR*,ǡ�ϻ�L�2������v�����E�:�|;<�s�wu�@����P�.O�",)��W���P.���WL�O�2pα��Z�,VC���Z�zB^��Nj6Zu��:e�FjՊ��E�i#��^a�gay3rj�Z|e���^��n�7z�ȱO���}\g�±7��k쥶u��+`�w�'V�dz,�Jݔ���b�Wd��wf���^]�&��}�ˏ���NIv	VM���{����Wdq��w�V�� T���C���AwU�ȱ�8�������{����P�8���l��⡺'DXנB�r&�Տ���`�5^/\^yxw�@����F�3�|��f��3��G@a�;��DU�� ԟ6+�HV�"��2c ?���9�".��z�s1#�}U&��P��$�S�ϲ�4nM�fI�8
���R�U�x�R�W��fOK���ͫ�!A��P���q�c���@6>ڒ�Uԑ�*`�;v��{L�R��u=�p&
���nv3ѦU�����曨i�&/&:A+��qV���]y*)o/��-��i��[qc��n�fB/}��X'T��;�[bڭaV]�s���)网�r[���+4��D*��`�Sb����[X�#��[�A��ߏ�M�^�[s�g�G�ܖ��pu�"^u�����>��dp���H{��7��a���.>�CX���e���+��>OϏZ�^=��T�p]� ���H�����z�B2aܻd�(�n[��h�r�p������f�<��8p��6Shm�%�5�+Q~��$,sЭ��vE@W�6:f�$a��,5�����g�:fr��9+�ض��&��Q�&z���֤Z�Z����/�y��!]�ʜ0v-�æ0���Sy�Z�5�R��)��`t��`5p:/څy��K��LD���VWD��k7K�Ֆ�^=K9R���(D��9h����3�Uc�~�)B�eL�s�T��ڗ3�8"hEt�����y�����A�G�#��J�IŹ�jz���Y��(<�I���<�x?U��_Q�I�#��T�����W*:*:��������aF�����a��O��)�)Ɗw�����Ε �x���t%h4��o+�*�|vH��ME��C�`�?u�N	��{֯�9A�<�ON?>*:ې��}~����SɡPdIB�Dd��M_�ڵ�5�vߌZD��c�	:��Fſn��B��U�W0�{e�ġ!�:���i����8��s�Ώb�r�b�As2��D+�#���N�_�C�)C�n�	L���D���|��ӊ��y���[������[��G��'�a���̯M�P(�]�9�\n�K�HYN���x��e�8�}�����way��@b�E]q|Ş>ưk��u�����0� ���,Hkk5��sno.�OK�aCb�^���f�P��*�p�+Q��}p�k� ڠ�-��M��Y͞=q/x{�r�z��%��.Z�!�+*f�1����tWwm`	���n��;��jQ�X����U.f����9�oW*:N��x���ڲ�g�9آ�_���n�]b/
F�k��qJ���aq����t���F]��"���k����j=��N���l��5~��\j���ʭ*�`��t�x\��P�x�g:*��ޕ�v����L)�ta�Cݨ��G#S�}G3�%NF�L����������1Q̶��M�@rutQ�0�dר�:��9ҧ%�음�U+<5��fe�HX�۵�K�T��\��>�T�j�bR��\�ȥ=cP"��;�eF95��b��]Ozh��`ؒ�����}CE5N=R��O��-�9�-�@	\�]�t&V=�%_.\�E��_��=�/�#LQʇ��cΒ�>G�Q�[*	�E�j'�V5G�ct�[��WN�	��G��퉃�\����/��
pBUB�=,�������:�w1M��[��a�n��U�8w���>'ہ秠�j�	Bt�H~�rjceEQ��#����Jw�i���"�B��@Ί�ns�W�q��<���&oD��>ڨ���<����H��+UJ�ȳp�>��ѳ�DtD�N�j�\�&u{�5�s��RWb�s��0�琡64l��6�L��e���P���_���Xf.3d�����۸cX�:�T	J�[ �����F�D�w"F�V�n�=�;�IPt�jx������*h�J����?UFKٳ0��k��Ss`gT�*oTS��	߉�
���'&�C���
ĸ��{�.�w>a{澀tFˌ��!a�s^�dQ����d(�U&_g���{�Y�NKU�5B䕈��`�WJt��x\.�h�|�ntՌxˊ���U!�*��:����AkN3r�l���*O��ẗ́��M�Q�U��M>�P`���K�wHuB�ӭ���s�mjY���P_�7�ls����5�ױx7�M��d��LG������@�=:�����M�a�*����@�
lv�x#����M�ia�z<%�Z��;}je	�a��Ƨ���,��U�Q1�9�Jz�L@9����)r�͋�5�ښ�U`�3T�wp�����KU�:��m"�r744�\!	N�ӗÙ�v�NF�<cP�u<�}��q�I��\�
g��	���׃�Z��h��uVj�,��DD�pKڮۻn��-�Y����_������*�vK���z��A�3ǭ�%��~U��},��6ǐ�Ψ.����<F��|(V�55=�Xs�a��9]<���v@�;����l�����C��n���;Ī�e8-a���Gu�,Z�Q�8¡��M	���ލ薥��l%Z.��*vL�lNX&�Y5��R= 8���?�<v��f�VI���g�TD$}u�7y�;d+SC�HC�A�: W�B�>��3wJܼeJ���,v�豋�(��ߓ�\�3}��U[t��B��4/HNal��f6��)s����2�~n�-E�O��uY�<is�r���gfU�sPE�n���8�S���&7�Ϊ�� (uU.:�h��L��U��u^�s��@��]�+�w'�-l	��;k"Ie-��%��\c�v�T@T}�1�48���.񫭃���ػƦ���z�wh��d��r�rB�^���MV�7^�R����A�r��EA�.{U�*��s(���"�)��0zl'A@!�;��u�4]W�K�-�t��Rұ�hف�#�Df�n��kz|���x��x�DS[��|��C�tnj�3��q	V��W��W��l�k�eZU�#��|�:`_,��;�q��=J���
��Ɉ�i�N������|��x���w,:�²}���m���ͤ��sh
/�M&&���4������T.���v�t��j�L{*G��=OX�'��bC-���ěJ�;�&'��q���
�|�{<�a��b䯷�I��qRVo��"�S����������3��'���
����e�c��<�R��դ��*s�&Wk��l�݃���ua����{��X��E��ۏ����1�4���K�3nI�3D)E�Rˊ�ט%��9�614[�[$R��� �e,��7fX�c�,��mgv��BL����b��:�{i��*D��ܦ-�{
���-^}�WS�C*f�nD���#@Ü��$�1նP�pW,.G.ۡ)�G���a{�9-귎��ܛ��u:L�Xz��e��ڪl�b�X��"u��!pj��2:�ܯ5�c�����V̂�eU�h��g�ܜ�]�'�9E�oR�`U�PY�Y��gG�������}�hl�I9�̘$�=�����;:���Ȣ@����Ǉ%��V���#�">I�2j3/2��yf,�i*Fn��:�i�6k���Y��E亍b�V�����"2����j�M�Mk�i.�S0�N!����R�w%�6(��ǣh�&z7��9@i�#����C;.��5g+��ڽs��v'ԭ���aU�|�k̋k	�vwd��X8s�F�a�t���Y�6�Ų$�n��lt�8��쨞w3��K�9cG����w�!-�s1���Qax��Ǜ���n�<�p�̶:�nQ<��"�ֺj�#�ĵmL\r��|�0;y�K^���5z�@���"=6���0hvh��[g00�h(�~FӾ��O�ܮ�g
Re[�D]4�����q�d�w�D
�Np(e�ݙ�O	�1m�:�+�W�I� Wϰ��(3wXP�s����,4�����\�&���gE��/��bgl�9)��gðu��?�6��:��Yo��֞�Uf�r��+�PҫujѼvT�y���LZzہs��ZQ[�hö/���lz�۔kD���pm��rBnJ�i>i���o):���+XP�Mز
�)D~�:�u�yz�a�i2��y�öȣ�49̬���k&�k����Oi��jT�� �uYb,��xp*<.�uҽe����"������핐|��2��D�{����ʤR�֠�|�B�˴�	AӸ7]��,�o�9$�����H��zx�9]l�*�G��"���l�ZWV�hI�V��6��4l���������B�N	�-��s�	,��/#t�Ҵ���wڮFkh�I�:��#]�`n�U8սX�0�(�]���5T���i�C*<����߮��܁��3PLչQX4�p�w�n���E8i��S��P��H��AQ��f̜�?JW�k�Rě��ds*-�x�vNuc�%��Cu^�*Y;*���y�ܬ�ݻ`N�⻩��.�R�a��l�F���p*Q�Rx�7=�S�IZΪGt��[
M�N+�����~}�Ϋ7	�-[}��"+}]bv�ڽ�TZ�F�ѯ�Nh1�����5i5M���Y~��},M�6\P��(
� �O� >�(�����+Tm�AUFҪ(#m��E����UPY1�(�*
( �1DPX����UUcD5�V"(��ATD�PE�1�KeA�iEEE��"���ň�EUX(��F"���X�������F+Q����*�+m"�Q���Ȗ�(�Fңm��EP@QX*,Qb*��X����"���QPV(
��*1TdX�ZUE�(-J� �Qb�UAPcUb���b�V"FX���+@��dDF(�*(�T

��X�jڕDDUjX�FE`�
�QX�ADJ�EQFEF*��Qb�"$��ơPTb�Ȉ�V")�VҩmE���"��ȣhTUEU1EPT+Qb�UF�b��QF(��eЪ����DH�$X��VQV5�T���@Pv��A�w�_m�_G��wmf�p��XB�'Ž]�*����)E��L�6RC3�{2N����3d����� x
ַ�m�b|�{�����|�H
)�?��E�u����k
����75g�2y�i����~d��6wz���l�h�qYR�o�rN�a�B���g�8��Y�v�.���Ϋߗֶrkq��<��`BAzy�m�a�z��1��v��Y���p6��*a��MO1E=E%q�!��gY<����0�³l8���Ag̕6y�&�Rr ��[é��t۞���\���,��Y����HV3����gSI�3��'�~B����I���i>O{�����u�)�@�*����,��z�"�L*w�O&��� Lx\xK����%9�{8g����w_��׿y�6��������J�8���&�^2u<?w�@�=C�Og|�q��!X[�C��8���5���O�I���9��|ɧ��~B���dD��T [a�V�f���y�����ϻ����I\d���:o0�0�d�噻8��Xq~���RZ~�Y1E:Ϗ{���q��i�O�v�ia�
�ɮSL�p׼c�=銀;Z֧�M}�JF��p��������IٔD�+*A��Vwa�B�a��M�c7�p6�0��6y�i6�0�������5�Xb)�j�8�3�٧��L@^�~� (��p ���n�.77|�z��g�y�����g̚�r��VaY�j}TuH,�'2�%UI�*|�E&3�0�Xg)
���������l>LC�k�&&�z�C������<!Ͻ0�����n��۾�:���s�q1� ~J��!�y�&!���iaS9a�{�i:�a�6��Y>q�T��"��d����V@Q~dѝ§*M����I�����r����H��
�ꚼg�0�ӿ/u��ϒ~q'�{�ti ��O�{���H<���6�a��1'y�Sh%f��7t���S��E&?�qCz��g��Շ�٤
�!�r��ޘ D�	��J��6A���_���-}�ɷh�~��'>s�Nw��
����_�˄q��M��C�(������+*��0�ir�J�|�0Xu6�Y��QCL��E&�PĬ��'�q��s���u�ׇ߾�QF���}�H%6Q�[�w�#��v�kt7�c}��PIՖ1U����dʩcEp��Dp��>�M�L���t��[�N�K8�:��*k�%�q��}ԟ�w&t뒸���'�_SCR9H��b�`�y`7.v�6Ԧ�ɜ_��� ��f�X�E�~�3�c ~�2x bT5�a4��d�O%�*(|��z��?s���'�����aY�y���r�Y���I�%UI�]�掠m'�ӌ�|�a���D�~]�f�%��7�c�#��P+4���8�E�j�Ĭ=f!����H:�y�,�u� i���m'P���LOIy����
��g��CĘ�a��;�|����`ҁ�]�Tc��}Z�F)����W����;��z�"1�}�Si�
���ud���B����t�����nɌ�'�{�1��ɮ�0^!R����M��l1����6��VuY�w%@Q`y�]�磷[��پg�������RW�C������&�a��T%d�?s%՘�P��0����@��z�'��s�n�L=a_̛��h� ��%|=�I��H)�s�rM�8��9���=�9��]W�3W����1��u>
"=��Uq�1 ��6�!�z¢���	��?0��|>�O�Cf��V�T�~����La�Y���J��ٴ��Y�M�}�vB��³���D��>��p�}�ɾ9�����#�#����Ӊ*�N'�~�i���q�9���)
��y�3����1'���Y�Ɉi
���
x�L��(��i �B�b�N0�O&����B��>���ӵҪ~ڽ��6�.��#�Ǌ��� �O�Vw��(�q�3߹��<J����}�S��@Qz�w��x��*Ow�<�|��ﻆ�z���q1����$�Ѻ)������^o[��������"��q
��Z�@�c�a���L@�Vq��a4��ɣvbu����y�oD��'5ON�'XmԬ<��ݝd��hS�O\O��a8���M9���i�9}��׼#�V��Tx8�1��H,����QH/r���'U��H��;�w�`i�a���f��1�aQO�f ����3��1Ci����OgXT'�}��SN`��G�J��
ǽQ�N��P���3ý�x��Vc�Q��B���vj���Y���i:����sI�I��w+0��+��gl:Φ!�i1�0�be��}-1�s
��k/΍�֏<޼�r]7�\����p۾I�f���o��H6��Tb��_*���!=��^TB��f�����]ʳob4�k��`�N��Y�qŶ�uȠ'+R��@g#`����h���^�R�����D��X�_n��  �{q'qy��~��H)�����x���1 ��톘�i������m'�+7��2m ��9��P1'����N8���4���Y6kX,�%H.��^��.�Ǣ�	̱Fcc��*#���؟W8���y@ϼ��r=�mq������ݤu'\zs2��>O{a��VO�{�]�x��]��y�@�T%M���������:f����!&������t���������~�a����|�!5�2d��@��O̜t�o�I�'�l����N3����<d7��$�Xz}��@""=�}�dh���[�yJ��~��Vx�3l�ְ��g�16k�Ci�/2E�aP7��C�J�:ɞ�wD4�W�O���T�!Y�o]���p�a�=�;����� ��u����P˿8��ׇ��z�ߺw�{�J�����l\a����j�g��gSɺ2��b��I6�e�&��uHx{����Y��O?s	SI:�g�S�w!�Aa�o;�Ny@*��'�7����y�����j���Ǐ��ɧ���:�h%t�YEq��zr��Oɉ�
�Ն��vOYyCٺM0�;��}N��4�����O�7��$��*�I�@�*<>�>�"wO�Ӿ��ٹw����J��w��S���<�T�)+�~�P�A՚a��p�Xq�@�+��g+1���O\N!��i'�T����v��4¿��d�r�$m�G�Ԥ?�8�����r��xΟ��I�c'=�(��Nw6�r��S�������0�s�3�~C�<9f�
i���w�!�bA՟"�gV�g�P�%z�a�鴂������*=�_i�Χ����n,�[�I����o_a
�o���6��r�����~d��J�{a�4�@�w�m�������Ýɶ3��f��� ������
���=E����2=��Q1U�ت_f���~���]O�1�Z|æ��Rq
��}�6�Xo�d4��~Og�`���,�q��Xii^�;a�Y����~���OSl�{��OP��M��w��z�2�{LI�*u���y��c��M~E1\��wٴ�n _3Sc5��Z��qD� �d�EݟfN�^��U������xw+���ykn�9���E���E�rdj���77
�m}��S�OhC����2�����^�Ng���{f���R���@�]���}��W�n����f���O�� �H�]$�TR���N8�!Sɪ{@�c߻�b�P<�1�T�Og�kD�)+����|�H;����{a��@���6��l�����/�S�����{��F%��{�D�`}�C���!��]yHV���鬛�4�Sz��4퓹E5I��qߙ�I�!�:�8�Vq����L�:�3���ɴR
m�g������~���<���y����ă�����"��+=�rM�ĕ�q���P�kt�]�bOP�Ȳk;�*��a�m��O5C�%N���3�B��6yCl�ayC�Ϻ~��l�|��9{x�~��IXc?&0�:��m ��'�;惨TR
l��P��C�����C_Y+i>g�;��J�HWs�?Y4���E�'��bO�������ɽs6������������V����p"<�ޘ��*�'�?[1&��Y>O��[HVaܦ�{��T�Ag���p:��Ԩ�x^��'�/�s5��LfÔ~����5b��ʒ�+���=��}F�Lg2{�*����I^����H9f���ya�'�����C�f�y�f�S��8��⁤�B��;��HV'��O̞j�`~;��:�_5�S�����3�o�E�n�m���o�v��Y���'}�Շ�B��:��Y�ufv�H)Y�����8� y=�{a��4¾o�'ɴ>I^��<��E�g;������U�2o5C�c����b������}p�M���g�4�P���&��J�a���O����J�\a���t0�>La�����Ͱ���H|�E!�~֏~f!����w$�,��<M>�@@�p&�2�l�?}z�n���o�|z��Y1E�~�����b^��1��]QCg<�]��
��×Md����4ZE�N�'{��J��dמ��)
��B�Z'��Ă��`yE��@�J��}�9��&����v��|��a�q���vo�H<�x��w�}퇈J�{���l��*O�"�R���+XuH9|��'����Cz���C�g̨(
)�OM�ͧ*M!S�s��so��֍g}�:����p(-���;;��f��ds.��x���nE.9n��U� Ϟ�nQ��;�n.T/s*�:���_a��e��.����Sr��J��k|�	� �f=�A�EԐW8��G������HN�~����+��JV��z�.G���TǄÏ{SL�O�ɦc%v�ܧ���D�}��H=�{a�V��a�4�Af��3���H���(��~C�bM�n���8��������̤��c������& ���z��z����NޠbM��d�8��w zsX��+4è�7;�L�J�f�ܛUI�:��ܚI�x�0���
�l�c7�p����ͧ�}=�ר9�Y��u�g8�,o}��� J���bO�c���X��y�Xmԩ</���g��m�N���ܰ���m���Xq�1�d�g���J�6�Ý͠(��4�t�𰫁�Y]}�2����� �z�5���Vk)
�i��:���LHoY��O�$�*,�jɉ�'\a��g����l;�@����I��qRVl��CH��)�����?!Q�3sB� �����v�}����G���l+��䞦��i�;���cȸ�@�?!��aY?grB��g�2y�i����~d��6y��R
z���N+*A���}�;�
�3�̟�!1���j�9t}+m/�@�q䝜���E �9��8����b��%���E�w�p6��*a��MO1E4{E&:x��l5OP�:��w$�ݚa��f�q<���A�(��O�~vkc�V�ĊÙ�X�DB��*|���Ci<g�0�=>��<gS=�8Φ�7��P�<C��ý��x��bO�ӻ�H?Y+StSl4��T6}Ef�děE@��1�0>�}����E�NFf�y�]���߽���1'�6��N�2N�a�=����J�8���&�^2u<��G*OP�S���5�B����Rz�L@�S�O�$�T~��i>dӌݢ��H?�?y�%󗗇߶j��$m�޵�+���D��� 81P 0VqRW��b)8������1��ٛ���Շ��� x�!���U�S��?;O�*O�Mw&ӌ���G�H��r{U����NZ����ק�}�d��+�t厨��&��$�YR�Ձ��8�Vl�2M�c6y���*,��i6�0������d{a��y>�,4�Ĩq�~�M�Ld�Ѯ����|�}�r7��V�*��h�Z[K�a[�x��eLN�V�F�o:���G2�0��!ݬ�W�n���qI���f9�q ٗ���1J�ڞn;�JoEE����u��q�lZ��wp��lE�+i�Wt���'�Iʬ�={��� �I�8}�߾��%x������m��5��{32��+1*9H,�'2�%UI�*|�2Ȥ�:�k�r��1�<���:��_���LC�*,�|�4�0��C����>�\��}�}+��Ky|���>���vя8��W��2!�{�&!�(b,4¦r���&�u
�Hnv��d��aSf���%E�La�
/̞w
�@�6����'�^R����k���f#gܡ�v��8��`T}����q'�u�1 ��N8�1�
�~�����x���bO'�é��J���3h
)5L0���Re��N�É�bJ��>���;D:%��RcU+Ͻ��L "@�v���
�g�ʆ��'\�ӝ�l:½d����.Y�J�6�C�(��;��=VT�sv��,4�W���Si��r�g�*)<殎xh��5�=�o~w����&���7v�m�bk������p�x�d�O/�QC�����D�+:��}����6ì+<O3Y8�R:�w�i?$��1��GP6��i��R_}:٭&�hoL�y����<%�=�E4ì�1a�c6��b���j�Ĭ=f!��a�6�ud�,Y��@��=��I�+=���	Qa�;����i1
�I��ɾQd���<:��#k��ķtm���r�+�%E�<��4���vʚN T�N#�OY{HW�P��I�:��M�1����M����H)����� ����i��!Ϲ��mĬ�"=U�8}ۢd`ӧܨ�^.O� ��;��I�)+�����0yg�Mj�ϱ�T�d��亳*��0����@�٫=CI�'\퇻��XW�&�}�?2W���N�AM>{ﾵ�'������/��<�#��}���>�����m�a�Ă�~�l�g�*(y�p�M��M������ �a�6k�QeaP?%M~����La�Vb(z��x�L�OP���A�\E�����R��7k+������XqR=gO߰6�IURu<�߰�~@�<g\y�a��
�'y�3����1'��`,���4�w<�i ��4�M�(��i �CfX�f�8�����s�N[����v;�!a�sa�(d�g(�zg�w�O8V��L'�SL'wnN#�}b���I�Έ�o'B��m���>��������%%|��O����J� �0���D��8Ej�Gk���a�'b��Sta�܈�įP;we��� ����]ڸ���}�'�>B�߬��7�E��T�o��I������d�?3﹆�<J����ߵ8ɴ��w��x��*Nw�n�������z����:|ǔTT��Gٽ@��d�?~���5��)����C�L�V�_�LaϬ1<7I�iiY��s	�Mn�N"��0�n���>d��{��6��VՇ5gY*?U���dT���X�gC�!����'�8�2i�l��M��
���<��>a��i����Ak�	8��)ԇrÏǙ��q�{q�gP�q�E<���gb|�ܱ s�����}�Dݶ�����3���w��J��2c=3�"�������x��Vcϰ�a�
���� ��bu%UI��`i>@�1���a���w<��q.<>�}��&���9&z|^�	�b��]&3�����E ��q7�s�>LC���rb��1��M$�
����3&�XV�_���V{�,3�,�q�ڰ�%z��B#�=�@�5Aiό�����}�������&���g��Փ�.�7�a�e'��ӝ�:��>s2���S���r>0\B�o�ɮ�<La��yt�ԨJ�v��Xg��T�=0������tI�?LV��w�������v|�~��N���: x��e��Y�J�~��H�>q4���'�T���n�y܁�0�s�{����^SB�( ��:��S�A�,��x�|��Ȏ>Q�9=�A��xϻʠ�t�t3�yy�LމN�⥸�kr�q>�s�uԴy�4�������ft��)����fF(Z�-k^1ѓ��Wl5�J���l6��X5���ʃGB�j�:���{6����g6_e��v<��C��'Z��30vN��C���W.wh�'�N���i�"����%g&��Nt9��TEѣuM�.`��R�Qǂm���d�q���5��(���~�"��n�M'!k���t�q*z��8Li�����lI����x���۝ݾU;;�>��Ce��"kX ������5�e�Ռy�������by̮V�yU����ʦЕ:@�N�dؕ����dddd7�Hen��p
j����l#"�/�MV~\vA�7M�7�ʶz�f������7�O��@u����<���p��q�ە���T��P�QB���s�@�
lv�x#��rm��3}��u���R�nQ�wc'���})1H��P]#�׼xm�B��ck�~Wٱ��#\��=�hF��ܧ:2�Cjh��ؒ���Tt�"�IeV��(Ho�I������=R�:�6Z�km)��D+�2h����8��#��V�BlT�87!GEJ�N|���囚�;ܢ���ؙ�����'n y�j{ʫ�O&TTu��P�8�j#*\d��:��>zy��q�{ܫC�5!��� /}��맼�WP��5.\K��r����Z�<}�R�d!�|D�J�^,=`��Ҙ�	KS1�뮫[�R����������?`'����M	��h �i��h�%��ٷ��¶� u}�	WP3ݛPN�yd���[�J��;�${+��"�
vf�T�� �Љ�x��T�X�o����} ��(hb��[w�g��Yy�"�Pٔ��Vv�� {�f���R�%p�w�6'>�AriW��S�6�Tw����w�)��G ��1ª2^��5��g=��Tnyx!U�e$0�/��l��U��{-΁n��"�Ou�x����ɻ��g�9�뮍�7Bx��԰�.� *��<chqW����4�Ж���/r7;yx���'½�]E�Q�{e�tN���*TC�<2�0
5����A�֏<�;����!�V�EC�EE���.�L�9�� �@�~��DU���Bu�끓��崵K�*hȷ꫅��Rs���""X��c��>���y;+�����ҳ�wZ�%����e()��P�Ywy��x�Nw`�LW����zy��3�T��p��G{��QvG����l-�b��sp�^%����(A��y�\TB�=z����;�?d���Xǆ���}44/j|շ�_���T�Y�A�"֊�[}ʝW0�J��W0��x�ܼӴ</M'~z�!g�YEB�b��cZ��~�~���&�E�H{Ლ��2�h(���Th@p���_
� Ua��b����z�C��n�+��J���8��n�h3Ժ؆nb�Ԕ[8�m���j��U���	��y�G��(sԺ!��n� T+�f]א9�)F𞜈��P.��!W�����{��/�-b{��Ѷ5R��Ar+��yװ0��k�3�ENE���&��Uً�O�>��Ht_2v;�G��Ҁ�f���v��\X�ΜS�UwM@��Et���6��e�(��qO��
���]㈡���2���.yL�*���K�<}j�Y.h�7F�w�G�b�26�1�q<'ۂ}�ЦP�)"&�(}EO�6�/s�'R�9�Y ��ܫ��Bk���|s�ϑ�|H�T�TQ����J(�~�7
�,�Y�Z{�U'�sBq��ڗ��`u�����e0e�<��!\`t���/����]�0���!��ɾ㯷��7�Zr`%&t5M�:�
�]��&n(XV@��:���-��f]�S�i#�Q�W>��ѝ�Z	�
+����͑�-K���"tIՈs7}i�gv,t� �U�~����H�7��ߣ�tcU�;��&\]�4��}�=1���xou��f�%�v�m9J��]E��V�¾~���8S�~P����7s@deu�L�쇆����(O+�q+h�d3*KYt%��n�I	�w-�	�+uI��w˲�@һ6�y��+n�����"t$?Pʇ��v�WK�,>6Z��yT9�qT G-ԛk1���18U��8��f݋pw:�mz�k��]�}�I��,0���%зXr�ptf�g[劉I���f�N�S���V(�d|t�ua�}�d�����,ǽR���c�+��}����1��@�����J^�ʵ���e��#�x:!�M]	T��e&�(buc^�&�����.��m	2'�ha��HAY��1r�J����،Tź��iG�J�ZC$o4��q�Hp�Uq���%.���ا+�F�BK���ݕ���V]��C�,|_G�'z%���cV;isD�TK&i���Q��ećkG#N���^Z�;/��u�뢮�v�-3e����d0#���@�����g
�Sۤ�l��̦��;�A����,�=n�=�A��T��./)]kR��tp�tU�<K�Er�q�y�a��FN����6!ׁLw���4��`j,S�f۱|*^��VN�mg;�7GZ<�p�� Hx]�w�I��n����V;R%�-�����R��z>w%�c`������u�a�w�R�t����S�I��T�_iZ,JO�qΉ��{-��uu{���ܩ��d-VwT��R�@7��wϾx��J:vE���=;�n��vX�����y8@O�|��V�M�0Bp4{tէ��
^�Z����u%it;6���ý�%��ȅ!���/��^�Kt�Jl��pt��9M�_bܥd���R��ι�p��b�����d@6������e"�1o^YY��y3��T����l�]"`G;��W&���u�1�Ԡ��2�2V��u���A���Y_��X�0�8y�k�*w�mR*α�Ne�E�m���d }f�+������L�f��a��9@�H'�-\�U�=M:�]r]�7�n��t]o}��;�)QB\������q�$�|ʚ�0�� ��Xf��4Kw�\g5��[F���e����ս ���G0�����q��7f�d;o�8�/��w���D�4�<���5�Cٔi��@sy++:�V�*��#%�ǒ�]���8?a��^6&S�e��D�I�y[!幚�R9*�>w:��w۔0�Sśe�6qa
��m��Ѭqn�nvP�����Ż$\X��̻���謣�����E�&�g}6j�S�9��:ˡ@Ă,�X�����ĂG��33ά���7GzY6鑕��e$:�v�v<4!�u��c�c:�4����s���_`�[F��vC"�L��2��d�ݱ{��@#r�b9>�]"��ʍ�:���}z�9m��lKc��8,P���u��v�q
�7�
Q�r�Vf�u�n00�Q���+W35ݨچ������ �RZV҈��j**������*6R*���,���
,b��Uk*Ȉ�V�"�cm�����X����J��6�U��*E�F��U�H��*#Z(�0UE"
"�T(����Q�DE`�[j-((#�����V(�*�",PE���#e��(���b"²��
�V�0Q`�#Ub��*X��*(�E`�T`�֢(��DAPEcl�[����J�*Ȩ��D���`�KKmPEUP����R"ȌX�*Q��1E+���ZT�UE�Pm(������X#1DQ��(�"*(�$b��"�D5,EkcDEEPQX"��(����UX�Z�X��(�EX�#UTEm��PQA"���ŋ�*�*UT-��Ŋ#
��X���Db�J�h,DD��AA� �4R"��E?P |*��
y���sl<����3�0mh�ʲ�Zr9�w#u5���cX�m��9!�嗛z�V���^�R��n��vo� ���f��=�Dt�މ �����+a��:���2�%�P+3�ۘY�-��8���ojd4��i�I(A�����f�Ez���E.#�,��|�c1Xؤ�S��R>����[.��C'��0#DU�Xn�O�����|�e
p"6+�'\�R2
y$\��^֮賯w��0�W�.62����ң��NŹ��*/�[���&��к��r6�W�
Cޏ�����Æ���^I�8a��{��p,v��l��O�����IS6.;%1(Tfw>hK�{�
e�����PبR�ߏQ�c&�@��y$T۫��(�cb]�v��n���|��><=S����8���~���B��;*Cx_�i�.�z��B�b3qf��B���aC�L��0�dVh�pWK�[F�)/���t| �j����6�z0��)Ø0tX��`{j�G��?@�!���C�Eq�4q�lN��_,.*�G�b;?<v�峟J8����S��8���n��<�����îE�����8	��v��I�7r�:����`Le�i{15?�L�����k��A#��O��hX�fe]2����g�{4y4WV�@��WL�xS+P�ֱ�0����Ie��v'ņp�������x��S/dbF�n����N�}�}U��f鉮�gW;�w����.a: yʽ�8O�����y	z�o�{:�U��4�����k��=����f��#L�iqk#p�(#:+a��΂��������9����t�w�U�$<�,�8���4��x�2!Uz�n�b���g")ýcׯ�S:��Fa�ޜ��WN+74p�&򙺓�¿��#Lb�6�*�Γ�v>X��k�-c��o=�Er���ԙ����`����qb'X����c�m#[�"�x"��wWgi����tޮ��EC��t\�S0J���Ա�UO+����*�}d�o�T
�m�z���T��>�t�ˀ`z��7���v�ܫaǯͳP^�^��	��t�Ɛ����8�{"�]���HH�J��������i	P�bc�	��@}Ad�7��ܪq@mj��ѝ:n���n�%�Z�u[I��jG��Eԡ3�!
���
��%��.1���T��IjQ}�26�SE�ؙE���T�j~5#����G��!�=�9�
�;_��2
��koy��h�?ZC��KՄ�y��K��R�l��WXa���X����i�@vþ/`�81K7��-+���☺>'�E�|�8;F��p<�̙��I��� f��뮓H.�"5rw:��.��i��_x{��:���d�ܺ�s�>>*�	�"^u��m�>�EPg �4�t�G);�z��Pv���:�=�L1t�c��R�z��. w�}=3�'y��=��/���=]�b�H$g��۾�NE���R砇W@��S�]iWg� ��}u�� _��l��GL�`;�\�`�]7�R�q�ɇBt@�28E.DI�w�Lu�(�����>��u�}�k�ʧ����høV�;RHp+�!!8!-��U�=Z��mȨEq�g<-߹�ҩ�;��������Tΰ�;���L�	�'N* �YU*�=&�"�jac�M��I��9d��C����e3��X�w'֙8d'55\|� @�}�1�����B��O\7��Vdv£�rB��O��c�pE���`4W�X�4�`��ʐ��Niͤug{�v!}�Gq0���?���ئ�	�P�A�=:"�� ԐدD�T����mn�O���S8�����`�s�٧'���x�DS[��S>�v!Ѳ���͑5�)^2���§�}�_Z�y�%ؙ�:����rO�ZEjs���n�;�9���W}w�������ksu��]�n�6Z�MD�wb�(�*<4��fM�"8��I�b��&�6�W�%��Q̣���5��H����k[��.$议5����x���O7ݓS��b(8V��3W)�x�@�Uq��fQ��.78���y�7���e}�*Ϲ�d�g�ڋ�
�{��}G|H�,V����0���#cL�g*پ��):;_9�yw�;��o�A�1aν9�Ɛ6�e���U���>�}��4raj��N�D�4j뙚���K��ݗ򪝺PU|0QN<	�~���\=P
vo��%5�EOd����#n^xw� �Bq����k�}�����G��|�Eފ���0���¿b=�i�W��^N���c�U8����J��j�w���v�MˇEOfZ�=�W*� 1Q*Y���c���=��O.�X��>oZ���G����lKY-r[�9]JgbXB��'� mL��	�e@"���3����D���iw5q/����5�i��\.�/>G�gʤ yGd�s*TM�|[�6��ݘ�x�s��)#**������lʋ��*oؕ0e�?�8�h`��}�l��[{h6b����eQ�*��x���X!0f�EW����c�'��mM�~#g#V�:	3�tҥ=P�
�lɬe`�(�ٵ���Fe�	:��Wה��K��_j���	t&�w`�v%�8��R��E!�2�]iT��t�
�<=�{�*��tƢ�g�2�8�x�9�r��r5Jsp9�>��613qB²�j6=(�T6����wE��h�W怢U8�ˌ�rד.:0W
}~����O&�fx�-+�w�Z�_"^҂�Č9�Bǁ�{��p�]l��2��i	5�x9�O2�ӣ�<���]�:,�&���u)w���E_Ȍ*���;T�Y����!�S�S�������+ӴZْ��� ���49�qw�+a�x�sd�/�~u#իw4ʍt�/��xq�v���!�\zB��f�U�
b
�ԻC�V,^_n+s��(����ogf,�J�Lf�oV9ce�Ud�:;$�"�E84N�'���}x��g����CXz��c����.<�ݧb��eCE���:E��n�Ԭa����@QE�Xj������R��_����jT=�tv<+�W���O���{��B2]M�F��:X�|�zNK��4�]{��R�ߏQ�y5��#�"�r��l�Ju��;�����.��49�o)���t}�� ۈ�qt��G�<1٨�j���G�@d�@|4��ٓBv:��q�(��W:C`�c��CrS�1c�yU��g6��;�J�o8��WR}3Ԥ��]����ehɼ�'Z���]��uc:� ���m��n2u^��l|'(<���uO/k*(��5Q�����@�(��Sc$�P+f/^lAYk��.�/!��'f߃�E���8R�E��t6+lr�}b�:*�U�/����	��{}�(�Ş17�у
WNu�^@#��G_�d[����x��+ʣ�A��S�F������K�ӳ��;�J��9��}���s�G��saNǸ�}ba�fi�"⢴��5�lN�1�D�t;�q��<���Ap���;
Π�j�GG96-����p<����gI�u7y��JV#�rwp�C݊#���F�4������������AE�ӎ�s�#����)S��v�D�k��G?6oD��Q��P`9)h�!��7L�U�����7U����bc(����M��엻��/#u����p�\XtN-:1\y�Q*0QÐ�ơ�_2*����Q�G;}%u��`v�#��������se����Mk>����
4T��L�v�d@n�Cצzr��}Q켽�<x֚}�§��%JhV���MʏTֻ��b��uZ�"���&f-H��X詍�h`+)R���m
.;'�S6�X�wP9�j�Ve1G%����HZ^�4H��ި%���"�(G�_��t���Á���Y��^�����LGg�|�įj#t�h��h�[��c����F��J�3aM��� < �}�,g��j��v�F#N{ۦЛ�[=a�j{}{�3}$���I�4�om��};�`̵1�V)"� ~��※G�2�捠a=�F&GG]ƪf���b��0�{z�`�&��$�m�%�Z�{I�_~5�8�{ǆ�R�g
��/�ro��������N���u��V�V����.R���5��Պ���46��*jF/t�N�w2��3�X�3�5��r>.��NA�l6���>�Ex��>�i������f��j⻱r\��H��jC��Yp�f)K�`�v���X�W@��'j*��:x(N����{y��Wp��L0��q0m�Qp��f�Od��.N>�:�w�.v�WT�8�\����n�5jR�*phN��2�I$_;Qc��j^ggރ�B\��[�t��ڒ�:��͔��x�]�3���WEԋr:/��P�[���E�T��7��Ɛ�9�f��q�ULuVncB�o.��f2��u�\�������$0�.�}'��~�]^����(�����<s����k^�+
d����Ȝ픴e�-ԨI���w|w�->(uۨ׸BBn�+M{�۫�v��q���fۍW���2_�q<�L�v�َ�Ǽ�VU�HV�峡�YG0�b�9[!���wZ#��G!�ݍ�sy��o�����w1(A��%��l�/�@��]�)u�>�'�梆���a����$�K֍lܐ�ޭ�Y��FR���p/Us��B��}���+��{��H�<h��|~�gn�K=��T��F1 t�QqPoqc�#���S�r�!ߡ��a� Լ�j�d-2V�6z��/�ʳ����W�a����<v��~��
�E1$7S	:�Æk��=�v�Z�r�٦3L��!8�NQ�XJ�������<�Ǽsܸ�1�t��'����ֺ������}oE;�G����J�{��o/�wM��o��V`�v߼tr��XYy3o��9�g�+�`i��jA����u���dk��>�n$4#-
�w6W�r�sy9�n�g�� fb(CBuH.���x�U�Έq{"���ET\��M)��� �ʚ�KyF���y��Ay:7���6��ۗ��E��:Kν�����c>��T9W|�I��+����.MH�j��0�t]K��f������ (	R�pk��l�Nf�	y.���q��~>�Uw��2[f��8ꖪ5[%�0`|\#"v\ن�K7�:h�\Pv�Y�ri3/E-������T��G��)�3d�Ghm؂�Ո��]L��!zݽ��H��K�n\�Խ�EjՃc�TVT��V��{���4�ƒ�(W�W"�´��E	@��2���'I��5
�\�\�ۏcW��ʾ��xa�0��$p��K�J_j?e
���)��8y����d��*7�����*���]
Ʋ�C��*y�|����ύK���ix��V�E%|x���WZ�7!�ڞ�eU쳉�Pk���/=��i8y�'^B���%�d�ŹM=���3�z��|��o�!E�{�:.BSq`���u�������
��(��<����4��n\�S�ߍD	9J<al�9�Z��L�x�E����y�P�vk'o����aT=O��E�\)0�n����v�
���G�ު�~��{C�ǹ�$����!�n��B�IB�ą�EgԈª���:�N�_�BO?\���BS{˴��N3:��~�d^��Ce�H����Mp\]�+a��S�u�0��>4}s��b����q��)�u����0�8�\��e��^���R��K���b�OQ��Wz���V��򻫷�Yy�$.j�vc׃��*��E�������*�f:��93�^�p��i]Yl��a�d�b57�}�$������\v���p�R�si����[��tl�]YՎ7%��kD���j*�w��"�;D�;�&�� T��.N�r��"�������9�1�nX��R,GY�:;$�;�O��@h��!���l_���vʾ��R�FA��92�24,����r��ݒ��>.2α�$p��;=(zZ��R�B�dzT߫+��W�0�E�\"���ug�ｼ]��˙3��LF�YM�)����3�%NF�L���AE��o�ɉ�����X]>�S���rXs��;�r����X�p����Α�fo�	�G\H����R��V��eH]�o'dL�4�f�s�H����m2%�eF9�.��m�lWGA����U�����e��M�~�[{ �좜�:�/ x㾙a2-��g`���QҠ����v��,RY�<t���e9�uT:=^)���s�G���zD�ӹ�8��s�'�����Զ*7���8!��A�%n���}r��ۜѮ�7�x��四�FX�� �5�pQ���g�a a���X���(�譆�9�Qu�R7=�Jj�VH��	r���h��w:	-n7v�+�� ���ZD_e,Hʵ�@.$�x�nK�A�N���Y�3M1p��sA���rv=��w�9��і�t�_'��\�
	��t���@l9w`ʾz'�gD�N!|�Y��˦v�oY��zu��'�A<zq�s7oLqY���b�8�R9���M�y݉�RJ�Y�s��e8i�[U���-s=��`ȡuc,�h��� �!>j ���=_W j2]�̮�*�s���ƨ	�d���R�����r��N�3^֍8���ڻ4�2�ŋ;he
7sO'Mn�&ɭ�/*�+*	��r�y@��y^ڹN\������N�
��'��s]���+�$/�l�Z�*K��ǣ-k�|���������q��T�:���af�8;Ƃ܇N�z)H٨>����9�U���ykݏ��굫Y�q��&�	��7V���U6"w���dv�W��=��
Z�g+Dp'/�;�cC���P �K)"nMJë��U�������v��[)��N�0��h���<`��mm񋨅�v�:����e	��v>O{\�\b�#���Y��������&�����t}x���|�۾��������]�ҹ+�|k�4 9	��va	ve�W�U�`�,�b�uI���f��uY�t�.|�R�'�ʎ����p^����]h=Añ��J��SY�R����w7'�$�v�-:˒�3�:k�us�F�X��m
Y�]�A$Ns�(@.�{��f�]�\�@�3i�%}R�e!|���X�=t�y��s�"�=S@TS���Űs��aM���uv�V� �{QK�i*�<ǌ�Rw�ND�Z3si:���c0
�ܤ�ks[.��)nFk[3�Heݴ����:��0�4�^չ�s�e�ud��c�D�[���$!\:�fa����1H��Ho�!� E_XoxD��y���R�0L܎��*�2lX>��k��Gj l��|u�i�}�>˭m`�z��Ë�tC�'�/�B#DD*$����>�t���N�Q�{0m]=�Z ��+4��C$��k+/QFx����P���ᘶ�=Ef�WqKt�՞.��1�ˍ�֮@PU.�&���o.��u-o�Z�)L�܀�+��V�f��X�!w>���wСؒ#��9�m�}/�s]B�R����8V�@���ʱBs@�0��Y���8�E�͆�\��Y�|�Ph�꒧���C�11���lP����-���+W[N�\ĹB��vQw��-��	�d�ԥ�u�\9�#mE��/4nK�5mlT|�]7�1ү9nk鮴�6�nZ��#xTo���S�Ym�v�Xf3+fıcٺ�J�V�{lZ$:|���
���i�'�6��y���.F���ڰb�o���,� ��=EX�`���G�a��`�Q�E�UQTX-�Uf5EV(��3db�(�Z2Ҡ��b�1�T\j"����9J�,�h,F
����*,X����X�
��A@F(#Q���1��DR"�Qq�(�#-���J�Ȩ��1�%E��V1QPb+L�EU�(�Ub+m��H�����lQE�Qf[s
���DH�����UB�b��*�iQPE"����L�T�"�(��Q��
�[dR�DEQ����Db��U�#PF�DTV(�c[�eI1XȨ�+m*�T�Tb.Z,ImD�Qf2c�*̦8�P��TX�TEq��b�%h����"���QĪ����30`����ƱJ0QL�E*(fc�s-�����S��r�U�QU�Y�E0�Q���F��*5-33̴TQFe�TAAd�EƲ(*�mTDQ[**5V�4f����(�X{_!.OO,�����Ey̵|�m]<81�Ƿ�������P�u)i}Iv���^�=���{�Nokw�w��<n7�#z^:�(��KDi>�@B���ꌦ�%�g/xF5����j�%i�S�[إ؝��p�\_��͆����8�F�'�Ƈ�U{^�g�wrW�����Η�]���ö"ϻ*z�t�{D8��P��A�d(�7
S�]�B�#F;���YT,Ͱj�EEA��`ߵr/�LdJ��L�u{&�G�ba>fu���n�S�u��dk�Cb�	_��E�r/���m	�U����٨!���^\@�l��ۙ��֤�Vm��>J��BF
PՏ����j���� ��t�4҇nKU��!f_=��׉,
��o��l�)U��23B���.�e���VԡJv���Rwi��\�����P�ç ��͋o�h�5���c�\�ct�g�S�G Ky\\1L��V��+�-f
`N��oj�����v	ȇ�FF���X_��A���ӌ�U�B���V��I,�S�������EB�3�����:�N�;*z�Cz�8��{t��y\���O�k�NLJO����Y{8x�QÓT�j�lB9%���əu�V�RD^�{`����Ej��䐆Ӕ��]Ve��5��%�m�i��K�ǲ��Uү6<iY�	nߓ/�ݫ�#����<5���]:E����D�r��p���'��0�Ǣ`�T\��X٫SТ"��>�:�n�c�gб����S�:�O�Ux��W(*;B�4�SH�"�ڋ�,#��|�l&)B8���u��ޛ��.㯗%3�/*�5N-�k�*��R�]7OŨ�
�=�ǳ���e�L�6��q�;���<��c�����zL�D��x�p��2T+�I�Ȱٳ���M�`��\�Yj�"��zuIS�2�_����i[5<PU�.}�}�0���9D�,7Dڭ���z�슗�Ybs�z����<�r��e���pE���B�De/�w.3
//��s^��wcɠ�.@S�t�T�\X1U_�T�r��� CkV�:t���Ą�����o���R�u�*�xj]%c����߳��x�bKu0�\��]�n��L��ޏ���W���R�
�%Y��3��ⱃ��O11�u����2�X��Ӝ�tpn�LW����L�Qw�Z/��D>��$f+i�Y����S*��WC_M5/wl�^��S���,n\XCseLN���B裘:�e���N�u�RɎ¢f\��
�2�J��-RVvok����:��De{	8���r)�v��.��,Y, ��ط���������z��V�ӇWV��7�����ɐ�u��U_V�rsțY�OOG��;�����Rm�� �w��V�25�|�qek�[��)�mj2���-i�t8@��,B@N�ߝڏ'H�HprEY�}�T�=��wN�s���إ�[Yr���W�GA��6ƣn^w�=:��``���Te���4���r��y@�z���E�"������1��|*ui_Gz�F9�;E�3�R�����ɽE�Rg���K��W<�T+�jT�ǯ昔#�L��~.yL�W[�S�Βo�Jnt��m��]�z���TP�jR�hO�@��E$Dۥf;�lvu�Bܬ2yJ[��)eܣ-�b��J���d0��-NL�K�&c�iz���#�8ȯ�C��P�9>��T�/>�sƯ�7�®�W��'���&�s�o"����0:Tn�����]D�MRh��
���t(ءӰ����r`%&t5M�� +��3�ъ�s�ݧf�WR�U��ҶH1j��5$�����'��p��܅���LD�\�skw�)h�����V���'uGŠ�+?"�W�m:ܽ1�흕���P��t9�p��P��>O���u��C�kc���"er�8����#V!�a՚
�w
ˉH�9�ٻ[T��p�&T[(�*M�����6߳�{��7Xfr�{�ޖyp:�����?z�ʡ~�)p���f<^��L��3�,�n�A��}��),����T�c�c�$��ߊ�HB���I���ɠ["��*hN����;�Qkw�t�rFˍ�Q�~N�	L����4��z�]��.�-r�g4�08-Y�n�HvV���鼡�)�Ns������;ƥB�E.#�;WD,9ٛϕj;.y�Y�+0��#0�#zm��j}Ԫ�o���'���o!������Y��2"�9}�\l^�t���v-�&ʋj��LX�S-1�c!�YJ'/�s�7����Rt]�J��������l�X�H)��n���]��,T�d����c]��]��]��X�=n�W��u*�P�G�7O��
�|̡�VXM5�swru�K��nR�W�QqG\�o�"�V{YQDXDt�l��9A��Y�i�O���	Gǖm�������)O^�E�	�p�ҋs��lV߹Z�"�tpj��w�Sãc�J^�SG^n�m+��Ρ,�\��{bfx�`ö�U�uY�f�f����w8���e2p���AN�3!�Q�<4�맷��e
h��x���a+8���ҽ]�ھ6����n��a��f�i��,_q��Vk\ؽN~W�W�ur�N񰦘��z�$ʎ��Qny͹} V�w�#��\��v�}J�Yx���efn W+��2a��N٣��(�xeE��c�=l�Ҏ����v>"c2=US���xı��/x���5���|~0�	-�|Ĳ�����Q�!��(��%�=��T����{���˹r�N�>N���ǼZ#L\Z��@�8-�T�'��qW7�u��}�{*��lA�L��<�]�R�<
����Ԑ���>��zܷ�fF�xN��tzv��q}�N�L�W.,:'���}�J��`�j7O^=/e�l�o�EK]�Q��q�B��Re�fb��#�C�5�h�qj.ެRw�!n(��7�*K��aԌs���9��A�FޣnE��l�R|�Lߓ��-�j��0M�-�vd귎�I�H�eepC	����*��;��ڜ�����N̹t�dޮo^t+ =��e�|��-�s::b=X'��H�q�h��Sr�<�����\����n�$�)q���\&zı��"�J�t���fvye��0Gp	f�+���Ss^�k�v�X��5��&[Zc��Y��]`�8���	`�Q\�f���^����6ss�f��E��]�.��Nwu3�ɍ��i���[�}��q�VOA�6�G��D�]e�W��9Y?���n�B�����G�x#�Yt��&,KſycIB�]2)U�U<�[�\{4{ܫ���E?��Ar��z����\��Ū��m����"�:0/�4:1OmQ�^s>.�	�"^u��m���392��Zy��r���VZ�6����,NQ�`�՚���� }վ��������1p�%�~�be�<�}�;gK����ʍ��M1)ҏ��ʠ�S�`.� ��puȶ�[޳x�[�'���r��
;d+ht��J$F�&BM"$��ڋńtU�|�ma�Z�ik��u4f^-�/#X��dc=�V�R/�G@^��!X!*�NeO�ORt�T�em��ok�n�%�Ȩt�������>eW#�F痂f��_$0�-��]��w�k�'�3��cWhh�P-I�J]�P.�}
����6�<XT�u���M��f�xpbzN\��g֋�48�>]]j�7ƪ�!`��lS�%���]/1�mkK3y�`0�oK�uxM	7/2'X�s4�w&B�u+|���#����Svn$ ��w�v4�k�c��Z<[$���s�f,��|v:�t�X<��ЖȀy�+0!yg����=tY� ܩqS��k���d�\Ș�ѣo8m�I.S�9\�~MV]�~z�^y�_9Ű��<��:@��R��x�և|;�r˱����z)
�&��uW��x�&��x�LHT��+��ړێ{��4��}q���D쫪���� ieJZ)Q*ϼs�pR��<ࡥ}k����V��exg�pt����}J���x��@6g�RG1WR}�*`�µ�;�p,Tە-�d�me>x�5_%��3d|KS���2���"�l �ьV��w��o�#^���66E#�W[/��vN2��	��ٮ�W��\�3㰂���G�L�͝�8��G���o�`Eu�i�,dYѝOު�+���Y�kC��GA�^Q���k��E��)�>��{���I7�Xƒ��~}�+��<$�"�T7d�W��FT�"|��F9|���*�u�����2{�RJ���9�.g�j']S(V9� хA�?D��7�甙�dYQ�����˛�:�WG,�=�}��B�el����Q]D�)}���+O��dTo:��J���J7Gaf����m���!6e+ǣp#�o�g+[^���8y3���Sz���F.�p8T�H���piu#��v	�@�om6Oόzi�,�\ľyY)�Si���zl��-���մ�o��ɕ�q�
X�;�R0T�n���dyA�j�qhw��R�e�U+���E�3����)B�eL��E��/>G�gʢ��������վ�1X���J�v�)�jz�W��'aA�[2��>9Sx��8����p\�d�� ���*<+Β����c��7���܄��ˡ�m:�
�}w�l��P��:0_~��q�
����d>D[�f�����ʃ��^ˇ���5׳�a~̰�t�����gS��3��� ۥ�B/��'�W@���UB�ʉ�9M��:AM=���M�&{zԽݾ]1�:�~�B"lz`��7SfR�.R�H�:*�Da_?yҞ1\��#l�մ�u-��jkr�/dt	���`��/ � �b�49�qv�l84x�c��%]�����^~�IT:fu�s���0	q�YZ"�򓆵LF�c��u�Օ'(�~��h�_�}J3��us��5��1Xؼ,���B������\qU�1�d���|UΫzgov�
����i��FE'T�T��윆s��ct��ӱnSuѻ�/R�vs}衏�r=u��i�X��^��Oũu��e���������l��WR�Պ�C�b�[������Y�v-%�j�J'�9ڽ�7��+&#��𕾩m]����]��ҝ\�W�Б���5x��ܧѢ͵��!����k�{&�Ӓr}2�R|������YN-`'�g���
{9���ZNMf�>�km)^�+�މ�GN��.8�N�ֺ�@��-̓�adO�=]�(��w3�:[y��"Ԑw�l�J�t�����U+^u���}U�l}���h�l�d~��₹��ٱ�T��J{P�_�8WL��8%�ح�V�M����o��[YS��(Op��1U���N$�p�AQnps�r�* ��}29:�xKg`��:a�B)�ʍ�V9��'�
\���ч2z�2����9l�ҋ�����U�i����7�\�����+�(��?r��M��G�N�u�W*:9�up�41_,M\N��U��n�ʘx<4�((�uS�ȿ|{��#LT��Tz��ʽ�{Kn�^�� �v�E�앲:1N:�7�Lމ��G�0�/�KDt���dC�^���X�Yo2z�ձK���1N7�N�`�؝��K�r�âp��7f��PB��{��l�K�9.��Ս�v]5qU�|��B�Ec�ق�`��ڙr
�S�=�Od����43k���w��2�~Y&��2�:�*�\��)�݉���k�]y�����$���f�[M.A��Pl�)�б�uڑԦRj�Է�bR������7P���I;�q�E��c�B�J�`�7 f�!F������[,@���k���g'�SL��V�9��`T��w�W��T(��r/�Ll�RBh2�B�B/c0�o�bؽo��Ibr=S^�s2	��A���n��v�E����'��8�fP%s�)Nʹ��m���2�E�]�{5��^����U������2P�G��T��[+�(bz�:��Bc�K�{�㱲:�PY&��0l4rg���4Q�S6�(��2�b�7%LL�+�+�L|<��De��u]'#�>] �_fŷ�ltf�SD<;|�\iPU��}����֣n�-��S�46!	OmQr�s>.�d' �^u����� ��f�imt.�B����)�j1��`�(�����nB��e�&b��b�|���U���<�Ͳ�PF�OŔ%�ڊ�c��"q�E	X��C�*�٩�4q��۽G�!���)�!���h����7�aM�(u("����	<�Bņ�#����af6�����ar<�f��l&��0����'�z31��i�P#\�y|�NdŻXv�h�n�fPc������\#1�ɻ�y�G�i�5��2�
��a!��� ���4����`��=��nu��ɖ�s�p�T��c���ZѴ�r-t$ۼβ��XA��|T�
��
�vA.�]۩|5�90k�ZT$4;-+ɝ���j�U�EV�(^�������\��c.����x*�a�R��bGMl�ƷIYO6Y��ܬm,]x�@vb��˙=)
*u���:e�3�<9���vvR5-nv���C��`��RhZg��2k�`��1xu9�ڠ��m#�Ez��-���6o@
֞�-�ZL���r�f�Mt�O�ރ,��v�/��C��=�B	oh�ƛx+��ٺ��!;�P�J�0Y\\�W0�e�I��[��n^�5��AR��4���Ua[n�d	k�p�Y�_Cv/Z��e�+��,����"�\W�Zy!0e��#���u;�Ӊ������dY��o��T�	UV�h[��k���Wr�N����
�4��������-8 Vڥ�sSˊ�Z��6�3��Z;U-�
-"4֌�BPV�(��әYW���5�	,%̈́QHE�BƐs6ƌ�\Q��L�3+#	�����ۦ���rE�{ե��3��gc��x���Y�eɓ�9���j�$v*�$��m:v4d�S3k��]�<�4�Qs��+V�E�^yc$��n�|�K��^���72��u����_{/n
���}���o���ur6�kV�;���j�$�&��S%����v������[�w������:V�J@��d��B��rJ�72oS�V�I	5M�p�Ɣ�7���0�IM={H���1R���O.�	�-�B&�8�ɶc��D��)�xҹ6�\Cahd��ԫ�����p�u�J�1(gV*��]�P�s]sx���Ox�e����u�v9h+��Ԍr"�������$Y��,�]�ҭ�� �����ߖc�]���l�(�����ܜ��ᡆmC�2��зS!bQ1�\�mL�ǻ��]4P���=�I��j�Ϣ�n�a�	���C��c����U�hmv��:�|�4,Ƞ�����ne+0WG�/N�	=�x��&���-5Tqh�"�=kEšs7�H� Tyw�N��;3�8o,��-�w4�;ܢ���&�X���c8ܐ]2���n��/���ʊց&��I�w9۾���癉���F�-�C�֌dSw�+�����OE�S�$r�6�\�ԫi��m>��e!�ЪwXa�j���;��E��v��������V�TƁ��SyW���g�g1)�[�{Nv��yL�>�'�CYW�w<<�ҭαX����8=ےk{��F���PN�,n<����O������T�hTU̳Ls)UZփ��j�f	R�1r����%\�V5�5Q&0�1�UQ֢�EX�Pb,bĈ�Te�s2)�.e��-J*�p�����[@b��s1�UETJ\�5*�"��,b.[���k�Tp�TEUQ��X֣�����F��L���ej0�EJ�R2���PADA��*̠V0UQUX�
�X�jUU-UkEV�U�DE���kB�E�E�[-�� ŋ[U��F�c0[JV���Pb��(�"�*���T(�m���-��֢V�TR5���`�mX�"�ee�AahՋZʩim�m+Q�Z*�*�l�"�J�YR��R�e�aY-�U)J���-�U��aR��V�V�Q%m�dR,�*V*��-��Am�V�,F
-h�ԨڴT*X�#Kb�R�J�dm��J$�V�ԣZ�b�XXTYf��믾4U��@�U
9̪�Z�u�:�к�h�}2��)ms�I(��v�'0Nu�1�OD:�	��Q��b�.��fE���-�佷?���jf8�g���t��E�#�W��*�B�BV �>�^�#�J����R���4e��)W�p[�q	��V%�\�i�6�8�5\"��#3sZ9��ۓ�A�=�b����o���[��@��]�)u�>���6!91@���E��뽼g6�s\Ҥ��a���RύC���r8j�7T��B���\t�pE^�FOU�[:�j���>��D)C�Q���$v�T]�./�1U^��.l�(���;v�Y��y���dg�+!��E?7�蠅k���*�2�������/%�1Uب�ٜ	U��Fm��w/��G������쫯FCG���)h�J��g]�b�զ�z@t���jy���t�Q���a�8����@7�&}�$su'\T�>�Z����ǋɼ�o��y>��@FLZ=]#��(R�pܯ �,��{hŌXEE9��Do���r���|}7���Y�ԥe��ح���>�@�3�
5H����y:F�w���E>�Hd�D��
��U�.���a
�{&��r���3�kn,��v�I������߅�Mp��-�E���t�@.�ŕ�<�7�;q��2�o<&Ѽ�[B�V
�n�<�,�9\р]vp��qӉsQ�[([�Fc��k{0�oZ*P�|�x���&��O{�[X�#���Fh�m���T[���>�� 2���粚��5�}5�Ϻk 𒤊�P�\�"�ՍxT�~���Ų�a����n��/ggk��=P��4�p_vd�]O.EЮ��,��i�A��L�����uV�o�(����W���W��u�1y�>ω5E	�vR�W��Z�x� ����8�3�RE�,v ڢ����X�X�(V5�2��9�L�>�G�ʠ�gc똅wՏ���ѓ݀|��Ɨ�^\�<jÇE./�GR���0:�/MX.�����(�fK=L��u'15��څC��TtW4��F�A{��,T��Oʶ�ydk����a��͉�y%��X�f�U��R���/�]4x�����p�rӧ�	�K�R��U[��j���c�&1�U��_"0A��ЋW�(WE"F�M��Uf<^��-9�xX��ߴ߶tq����:�25����P���lz`���ߊ�HW95'gb�`���&=~Q_W��$z{�5�+ru=�}:�Ξ9MU��W�,���	.�:K���X���n�l��#��cE⺸^x E��_����y8F-d��X�t[�y6
WY��<f��l4�rY*����`�p6)�v��wu��^6"g2N�x�l�B]t#ԝ���7��XW�83�>R�����e��$T\9���8.-	�q�c.�w�!=�=�pԳ��^��P��=ˍ�.=!eh�3`r��W�1́c1ٷ-�r�^�k`�+�D:Őʛ�ј�l^}Df���,ce��� v��4��[��)�8�|�Ԓ�leK���'T�*FAV	�g�0���B�fS�-��.]�u\�".��O+v�ˮ|��fwr}~�����
,e�
�Z*��X�.c ���^5*��~69��ݬ��i��l���2�b��}{�8�kG�|��P!X��m�b_���|�fK��G��j�z��\�T���m��l��ĺ���WT��TQ�i?rY�:��n�O<�̓gz��8`�����No$�P,l�Sڅ���p��Q�r]���D�iع���=R��m�䮴m$[�S�P���"T(Pl����9x�:�u�E��/}�`�ߒȓ�S���N�;о�C��Bp)�4a�Tz��T|��g>�q�a�Д�NfQ�{�hHշ�3�mep��&��禂�r�亷W�ium�m/-��$���F�����Jz_��^�置ׂNP��o��U�1c��Cf�)y�������^f�%�9	��@D��('�^��y��Z	�p���ok�{Ej�>�|�x�-���x!��8!+$"YQq��FuA�����}���Y�{Uvq��N�iIb��u�ہ�E\���P$A	ө>~�� i�)\],���?G,Bu����ί�VA�����:
.��C�f�Rf��]a���@�e���'��&�mx���8���K�=Q�۵}��@.��|�)��'~&\+�j��4��T��Ԭ��û6ڦi쌛�GK��P���dQ���6
/ڪL��'s�b=���M���Ɉ7n%����GoO�-Eň T�nmX�U�~_8���~5u�>l�S.�j6��_Q;{Y:�o"3���^��[,�M�Ԫ0`����+�r/��;�P�E�v8��u��}����:w9b��0��A���ش���2�LG�㜩�X�����Vz�gk�L�g]��j��
lv�i������7��Ƀa��$CN�0*f܅�̓� �Y���,2�h���R��P����{] �Wٱm�����xv%P�zk�A~���4���əQ^��)��ytaK�ZMb�A��x��K�^х;�o�x���=̘�^
�޹'od�OWy�y!	�vQ�Et��6��t��]���][�-���^��Ь��7�fMLK�1�C��Ĝ]Z���t�b��^�o��+}sCL�1	M��E��g��!9Kα���TRQ8f�ɢ٪x�F����n�:z��t�Q#��U������ʢb�����q�uF��Qo�ʗ6�]!k����G���u��F�x�(J��,Y𮽺��l����]d����: �
���^
�����u("��Bd!�"o�P;M�����9�z�n���)q
)�>JoɊP�����n\��G@��
����IJ&�J͗�U��-T���Nlc�r*,ǡ�ϻ�gfUˎ��6��iӊ"@�B#I
��]Cs3�u:�Y7S[.�"�t�꽖�P/}
������6!91CU��Xi­x1��ض�}Z��Yg����Av<�ȿj�7�W9
�f^�q�eΡ����HO�-y>�
#�Ka�4hdu� 9:TTxˋ1UX�S���I���ڹM\K{�ъ�|�Tԁ
��DRQB�t6+�A
�$T���
���Ϩ����.�^T��ne�3�[Wv&mE��X|��|{��p��S����G'X��@ka��YS�)'���iE����]�TNU���A��{~T�TΝ�M7���O���m�˝o�	K�����^����qE�'.�l��c���;�VCP�[��B���*��S]8á\$��a��X�vU���h�� ��KE"U�x�8)�f����۷2������
�f�7N&)힀l&}�'��� k��${�o�
Kpe�>M4�{���\�f�b���t�Y)��F�Bܯ BElڐ{hŌX}'�Ϧ��VD)5����p�_����!���Z��!�m��:�R�a�v�,�Al�ЙW�5��8��
Z+t�����4�Z���!g�YEB�e;����V2H�>�^Q��Fܼ���=�6"�)࢕s�5���t�8*�W�]E��"��/��i	�;*�=X��s�q�;���'4�XewC����q�p;E���N)�����Zu�$\+U*Y��M1(:G���}e�Y~�ݽ.9���k(����>�1�B|�6�{>^sO��5ED�)}����+OZ��|x#j��x�����:�K���}EO�U�E�b�+�T�/k���z���tOuL�\�v�ot��a_+���@}
0�0�����p�q^�<��u�*,|r��&o�0�]��}�bJ�>����<��0�����|��H��xP<�b�� %0����E1�6�d$2�dY���c����bc���G�v��S6�ƚ�1��T{�Z$��m��
wӇ)��q3���fq�$��Ӫ�{�<��P
�9mi����EB+k�߇�4��J����/�U��D����!)��CTՎ��i�Tx�uZ틗��w@��xf�$n(X
�ѪpTźV�� �(��=��:��aLΞ����9�)j��N���!�"�_�:#n/iT.X��.�r[t<UY��t��/
/[7���q�z�a��x&\]�!��=0CL�M�)Ĕ+��a�n�[duׄ��JO5ݐ%��ݼE\�sY�z1HP&sw0HL���$T\9��׹�q}&���wC��ʊ���׾�&5,�l��J�S��1�\zVV��<��.�#�l����K�Vo �z�E(Fb�|����V6/>�3B����>�O7@�꾾/iU�����Gd�	��4�DhU�wĊ��V=���4b��6�_��a��=.5s޸|�J�H�%-�*,5n���ƯJ���u*�c��|�x\K�o���ڝ~硭�����Jn��x.7
��|�#��>Wдs9�T���6��%eu�],��kt}6.��ZD��*G)	����i_�bKr-i�������p�����Uܻ��4���bƔ��Hs���,�����(v��bT�|7��U�E�AZ/��a���f����g�rSSLY� �4PN�8�ډ�b.�r�����\:�`���p�E|��o�k���{$�γ��@��.!�뜍䊩X5�}uq{7
2y�콝0-�,��j�)D\�S~�.T���
�NÅu�޵�����@�T���}�#��lu<�iTiA�1p.��Z��=�Y�x�����%�H䕉k!�J�\��5�s<_�TC���z�<�*��<ʋ�c������у��m��#�^�G���&��sO!����$J�(�tA��y�n��}���ӝs��Đ�5�X�z:�}�	�8i�����~���Di��<O{ȥz����H�R�cQW|5��pq�l79΂��㡑O/#�&oD��q��P���f:���Wt��8\�
��dC~?+��C}����|�O_͗
�ź'���1Nh��^��U���\�9�`�V�x�y��t�Q�`͆B��L��'s��b<�vFq.[g����5��"_�� �8<�Z<5�e�c3����N�;񫮈��x���s»2��h�%�6�̧M��B��lȳ�%=���P�zS�$�}i�����|���R�����£�#�:�@�kl�lps�u�D��N�*����*)[�(��e��X,�j�b�%)Wvb�-�WӂgnnlyczS{��/'EE�\�����^� �����i����싵W�8=�^VF9�)澚�+���r6<�l����/ L�I6݌�=1�+�*rWC!����f����]Z��X�-fo�U5;�m9��7<�>��M�g6L�r����Ӣ����ZOZ�^���S�`Z+�Kgs���B���R=y��њ�mM<��m��y������Չ��;��@����u9\H�p�.�6��x9�~d' �y�6'�+5oaΔV�Rtc�fh[���2�}Mx?��(�#���W!GA��T,1J]�`�b�⩺ˮ�4�Z�^j��ZV��E�X���	�	ڊ�c��#�0��aA�AE�N{��B�S[s��O>~��A;����S���&��p�B���L�:�P�H������m�ʽ����[�ꖮ�C[�(��>�ĨHKS1�뮫[�R,)��HVK���vY�u٧ӥ�WY�._Oϡ�7 ��ekL�ʱ.:���7BS��P�9�����h���ӑ�]n�D���#�^Ċ��I��G�̩mZ�[u��C��9��2g�ps�5.6��Ҽ������C3s��v�q��	�[�e�4c	;6��u�;[G�Z��H�.��V��fvk|<����)�����A�k��ήuFǾ̶:�.H����] �U�:-ҁuL�.�w'֙8e�B�u�����#J�k��U��|+���SC���AwC˽"ƨ�p5O9�Y
�xf���A��X�5�W�C�N��zJ�r&�zj�u���矅��V(�e��z�-u�s]�[�|��쬑�𠘇�DU�5��+\�VHY꫌����ط�����ӭ�3:7ø����E1%��E3�~�F�4f
/��(�%Y����v��rj��w����N@}�r,B���(�s����T�����Q�Qh�o�!�kUƯ��nld��W��6(�}g�c����(n�l�i�i��.�c��9o(8��1�Ѝn3uIWoW���1�*��V�ڬ�E��@��v�,uH-���G�����M:�M�I�k�{dt�L[;B����7YNϑЧV\�~_A���xU��;��s脶Һ����e�^����k����:GPP�4��t�%��}H!ta�����Ga�e�v����p`�%�\4"���ջ�N�Y��V�D��.!����]Χ���@��*J�q�Y��Bv'��7x,R�8�,<�a�cgőw���=U,t:��{�����ueE���_g`A�ҧ}���i|��Ũi��9<�a���5d�Ց�՚���ʅ��i讖�T�lf���:b��u�M�[�9�{BSGi"���v�����˽��G���hF�j��^e*��׸[<��]s����Yͼ(C��'6]wd%&0#�T�p%w�<�2j�q�=	��xs���M��;�4ҟ
{+x����e�|�9�9���ʻ�b�ݓ��Y�~\z���|��Y#��Iu�r�KX���81t4sL`']�n�§��U:r��Z���<�I6�d�p���.�KƩR�Յ��]4^`g��e%̚Ů<��ѽ�"	������3jC��o�w�zc�ԛO�؏sX�<U�g	�\7U��b�R*�^���O��#���8�8������|�5&6�[�7
�������nVi�4s<sqZ���٬g�T�2��m�VV��L��	�m�)�G]��*�kz��?*8k;m�weX�ӽ^	�oc��c<�&�Qd����\������|�]�<���h�xJeQ=`�@���ïNbGB�[��L����C��F�#����mw.��B�\w�Z\#/�.���A;�s�]�$4Ȭ}aq���� 5�t�}5����so;�����傒�5)J/=�����,��w$��q�׳1(�ېR���K�X���_>g9p�2�Xwl�/�[��Xάح�r�$��ޒ�`PR}�^gt8�Y�s��8�a�z�TIr���[#'p�F���������k��X��VLTL-�2wb����@�h�k9��AP�����;K)cꆕ���1������ܦ������ئ�9VQ�:�ܗVZ�:���r�Et���GAcM�;F�F�N�R��a�#L�xEZ��Qip4�ah��R�	P1Bj��]�=�-Q��Wl�%��t�8��jh�A�*P�ñ�Zm�y΄Ι󬫘.�	ǓN���FI���Y��fb��-P�R�j;-��h2<*����4�w|-v�酭^Ի�q�oIܝ���+W�8��\ژ8f����ə����2��B�Һ*Ī^��+n�寥�l������"��Ћ�����db�nIP�t5�;�p��A1��:�������Wh��� ^~��Be�eR�����t*M��żb�-�1��k�O�5��'��"��fpI�e>�'wף�bXN��|`�	����H��0[L Q���l�`u>�o_(Z2^��d��"i�u�>���쳽ܗ`d��Y.2ed�����c�d�k�2G�J��Qh0WQ�S;�����S>���>�(;�N�9���I�1��Ke��#�E�U�E�*iZ�QKKmF
����,��DEKV��6�ʋ#����m�*�ѶFģZ(1�K+Ak�F��(�+"����-�R��YE����ŨV�m�1��Z4F"��V�+Pm+-��KcT[E�(�J�lF6ĥ�Q�����Te��kK�AEKj�ڡD�lmX�+lF���j5(�UkR��UQUUb�[cm����U��[H��im���TR���ʊ�mm-UU)llTUF�E+ic���F�)Tm*�6�5+VZ��1�[J��DZ��mkkD�Tm��"�KjڈŖ­�kV����(U+F��Z�Z�Z5�m�B�b2���¦'[�I\�i��Y�Y�u��
7��kVw���T��de[j\�>��ͦ.�@��WPNrS45P�F��؁/p�㹼\�9���+���8i������q�{�qB�yr?p��T�Ǯ��%<�F`�2�Y�ݓ�ⷜ�>�_�JT���E��F>�
],��35Eu�]J_oQaV��dagH����'�� )4�J��h��*xΩ�!b�-t�C��=(L�K=�h%qOOb����or�������(DH�4������ư8xW8�O��'yi0C�c����X�̒��Ƈ���9d��)�.���~B�
Q�Q��܏��Z ?S�Ǽ������{@	��x����s�H=+�5Е��K���T����~SZ�<PU{L���;;�|���t�=8�
+�������=�a\2%	�38��T�f7F\*�V�>���u,��{��B��K�fu�\]�� 3�=0ӣS�
q%
�8��V;cxF��R6�[j.fab�|�t�Z�
f��>R���o�(C���p������&�JX���.���Ppi��P�;Y��d(}�v�����q�+DY���e�J�ٻ�
�=��Vة�:���2��&��Yڰ(��vc8��&o��El��Y�4U(�h�È1�wKԵ�d��K��h���&��	c����	���ӑ�遯9ɑ�3#�r�ݯ��S���`��Fܭ��^5������>b�a���Ddo���̠�n�c�Q�����Zx�:��عM�ѥ�@�TvI�E֊p"6+�'\�*FAV	�g0�ر�7\���9<`���5�$����ӱ}9��*,����E��[�u%�W��qg���w���"��]�	��[Wk/L>4�m�eÁ}���e^��>F_:���_[���L���=���>~�3ѿ9��]���oƐϳ��CC$�Λup(��t;'c�����eE����y���5��ӷ:�Wp}rB�RϮi)ȧ*�JzƠE�NÅ.�[�FƘ�B_u򍢃{��?}�p�Æ��iW?���C�� v�ns���
�<2�z]�\���sxu��)�o�H����-Ez4QҠМ�U(dU�̨���j	�K��ȍ�CQ�[��WN�r���{���sO��`�O�`��,�����2���^�?G�ϥ��4���Y��9%�Gp	��y��9"Ԩ#S�R��i�͸�OTa����5r��]`�z!
v��ܸyr��o	���vSi�, �IW�֝S�f]�sYf�Z�����A�nJX7�t���E	�
��t�)��K�Htd$��r����tƎ�]��ky�}�J `eYY��b��������)=�Z��T�AP�9�[�9
!N:�7���"�|4|�
�������Ӿ*�ffys^��l?$0�7�"W���/x�r"�7Z��_`N�L�W.-�8"�CU��9���R���y�澂�W���X&��5|ȣ��q��f�!E�2���s<�嬸�ק����\��~�b'�����,X�*F��������A�}r���ۑB�1���cu�ܾ[04zc��Jz��+����+}d�o�T
���7�ws�U�� ��ko"q_Jh�	�ζz�l����/f�I��d���P�X�c R,���%���c�ߩl���ꋷ��:y[~}��C��>��M�͓��g*O��nQf�n3V���*�(��2}	OA�L@>��`mt�}�����w-�R���^#<���}$t=���Ԭc� �SZ��Z8*;*�xA	O{j��νM2�R"�0�C-<q�qI����˂�{���G�5��jr���Vj���2�����K�����JwX�v%;��x|�J�՗�[���jc�s�'��{w��&�[�,N�5uh1B,ڏ�H&������m�g� -��M�!����^
b�Ҳ���&'��GQ�k�deq>Y�S4���mmV�C���U�4�/X�} BέS���OZ������G<z�bSKD�P�'��ڭ*�s}�EX=%����	Q\�}u�� X�����L�:�P�*d!���1g�*[�Z�\UՉ~�W�c�VQ���(P��w��U[t��E�)z���Z�ޗ��nYO�U�gk�`�_�I�^�ժw�ՎB
r��*�s�zL�r;T{�@ʫ
u�//pwWgU\TЦb�F�h��)2.�
�t�����wЮ�ܟ��y�G4yX^��,p�I-k>�§���'�}�1�8��c˼j�	����̝K��eb�z�K�![,V<��D��נB�r&���r��EA��..�,6�����$���~���� ��B���PS��Q=�Z�jHlW���MI�
�U�F
}p��^<�P�>�[��Gd߱��P��$�S�}���j�*�k���-.����&�/���c�5o�wBWi�騸�r. ��0���0�t"%c= �L�jy�5=��Ǻ07M�x����&���:7�DV-�:v��mGC��%�8R�1d��u�	�#�%��RU��n������_g
:�CvN��ZӔ�ǒG�J����v�l�|�h�
p��0��tK�b�i�ܽ�3U�c8�l9�&ԍ��hsz���k`�3մ�/�wf�_�mI�p0�-���(A��y�a�i��9�����-}s�&�k:t�H/Uf?���dk�4�:Z���t7W��;��9�Ѕ�uH.2�f�V�V9���ɭƒ]w��l��(�;����iI��r��*�H�"�yF�����we�TQ]�9O:�ar������9:Kν�����`g��5�xIRjECvOA��H܇t�q�Q�Y��N���z��=q��n��qB�yr.�W
��^��R�y�w�Cfrm�����S�Fkzo�Jt�$���j�F>�)y�>�GQ_��r�{R��b�*��Tҹ�|����S,A�dI�T��*xΩ�#X��zʙ=��R�Df�x��<�S��m/X���� @}]��9�^*�P���7
�����<o-k�m�����r�3��������]?�(A������| lr���;Nz"�ɖ�"�q��=�gO!�9r3e��da���L�P�+ /F����s@S���^S�Z/'bǚ�I��w�*h�,�t�9�Y�&Z�m^v��q8*�ޗ+rO*˽#0���'�[m-U���|�Q��y��jd�z�yl҅�*fZ�x暮�o����j\t�z�����>jF�����6[��^����<���8s���)lWT���lR�x�p�֋��������T��,y�r�
 a��k K��;�s�g�������!S��+���G��	�b��u����7Se
q'��<+�=܀��$��oP�$,0W�DaTy�G��4sK�S��T=���(G���n��h���{rN��۔>�+�~B�Muk�3�9���Y
�v��<��p��.��(.$�!���3W4d/�+հ")}�a��Y�즰k�V6/�Y�����fn��v��;s��<┋�*�㣲M�v2��8#\�H�*��g0��o�D�*Bj�m5�u��B�1�Ty_iط8eCE����/f�ۡu%��	�)�YN-c�+�eL��&߻�?c3��{�>���ԡ�}���G#|�+�\��OJ��4�X�Q��2��yxi&�EދԾ��TadO���~� ����\�h;�vL�/ڵ�+�L����z�j���s>��A�r�%A�s�8�].�-�NÄ����|*��4|M�W�*m�g>���W� �iF��N�6玡�ȷfu��<����T���Kei������L�]bG�71.�K�{�WLNOzG���Sk����cUƻs�rޜ�>V9���ap����Kg6��t���"G�..Y�N�&��&��+���/].ԫUs�K��< ���~[�;�W�S�M��&t�[����_����\���P�J�AG�eFg�=��ֲ/w,�J���?�-��ӎV?�nz{�c�7N暊�����	������x��b��� �jiC�����χOsN�d�-R�"	ө ?OB���m=��R�rT�ɆH��N�
C���n_:
.�S��/�jf�E���N���mήOrR��{�>��4��#4W�r��uL����_`N�>���L��d4�Ȯ��{��8��(tp�ɤ��+���aW�
��3��U��i�s���!y:g�ʎ��
Q��:�nL+�3^�CD�I�Y\�^ɼ ��/P{���Rha	��j*hs��1E��Q��hxgX��)��y�WgWU�s��m�==��gh�b��Wq��㊎���'x�6od*��JnP�Գ*(�T=��n�{�krm�5!���X��N��R�$l�\A�����Q�����iu����/�u�u���遬�^��N���V]�wU�ל~i�Cy2�M��d�"E��ޝ9�h�yt{R�EZ�u�r	�7I����s��y�Ziqy����Y
9�C��wΜ�hƈ~#���;~��<��P���w8����
��qh�����[��]�ƹoU1��C��-�7)s�Z�T޵L5���*�����d�z�Z+����A���U9N5����.�SF����D�J�]==��r�����i�yڔvΧ
�"ޚ��J��Go��w���VS�i��/�P,��!5��!�Ұ����,`=� I���Ok�`����ﯗI�o�Ʉ�֣���[y.���srk{g�*㞽\���q��9̪�+�Z>���ek��qOa1��-302ɝ��^u�*m%�,v)�w�@İUuz]Tnu�m�Һ��p�۰�jV�kU�n�E�c\����(�FA�CUH��mb���1����#���.��)����5ي5���r|9��$營cОEV��t��(8���4g ���;C��u���-�5��*�Ks�r�Kd�{�����8(��[��������䀬܃N��1Bn�N�r��(�D�u��O'r�֤����F]��]N=Cz,ǥM�p�w�f�:���ܐӀ�����"��qLWd�VY�4�SI�>[7�՚}���	��4Ht� C�Z���q_u?g���@z���p���0d�٠Qt}�֯�Sn|-�urZ���;�_wZY�@������}NQ~������oR��oVS��,ۢ9�ՍOW"�\y�%`�s�Τj����x��y�fR; $���ɫDli]����w���/��w5�qCF��H�txn��32meE�U�N��nƮ�+m%�,�>L��g*���P��X�S���eW��r�ˉ5�eY���9���sZyX�EߙTy٭����Qrڒ��P�ն2N�oz��T���)q�Mr�ջe2!�g.��O�����3+�	r�2��Բ+�]9�+Һ�gt�Sj�W�B|�5o��ȝ�;m62c�-v�����}G���f����@����ߥz��`9�jssk�t���ќμ�[f��P��Xiu���\]�Kg�e^F�]z7��M��^%RnU�/הڄ��/x:��t���-��)�8zf�TE����P
Υ�u��I��u�6��jeꊸi�)%݃�ۤJ���.�:���(H��E��Z�ZƱK�����t�|�&�;�>��c��E ��S�J(tt�Ճ��^�=7b^���Ƚ��}�t~k�=2DgP���}&I�p�V;e��E{7"qű�7p��~��_��|��}WEL�5KڪE�Ek3�;Ί{2v<���cQWx����ߩ�"__XL�6��(�ᝳ�F��0�iv��ʤ�й�(t��H�F�z���&������{��LO8�,�C�E�͝[ҕ��&�ء�R��³].����N*��p��7""��c|5��PH�|�ᮄ��UߋR]*����L^է4��6X�ڤ�d�|��p�J����\-d�7b�*��ŷS5v��C��f�>��x1��,�=��i���g���^�N�^����%eg���4N}�geI� �������Cns�{w�'D=];���tc�G�f�C�D�o��q=���tx�Mu�I���R�j�6�S,Cp�A�zPͩ5�A�t�G�i Pߊĵ͗�VnU�w�txڲ4�q�F9Cċ�v[�D��?��m	ܻ���j�o��W�z�|�Wx%<\��G��h$��v����3���f<j؜�yeO��&.���t(0���j�7���+o�ǗhR�+�6�g8�+jڪ�J��-k=tBQ��vM�%a=0X�{X�a�rt�u�+��o��<ӿ���"��˺1�x�O��y09=���s4�ȏv�X�r�؂�M=�,7t� �%j�Jz���օ�p�cF�Dq"f+k�xC��0��ףJ�);�ܬ�	�y��N��n�}�PsZ_br�i���\��:��6q�-�������T{gv��}�:�R�;:;vx�!�0,�y
O���n-lJ4�W^6I2���W��wG�����jM���S�a_���08�!M9z��4v�@����bUj�lln��ۉdm�ZE��m샦V\5_[��b[N.\B��I�c�j���T�2�lq��w]�B��C2�ܘظ�}�S��n�ƛ���+��sSjY{�DL=��PQϯ���Q ��͘r��J$�n���P���B8�t/.��Nu*��"n��t��v�����X5��|��!�ϞQ�*�T��{7�R�	�ɞ#>�a�wx<���`L\��^!)sfFM�"k9�ᝐ��xa��d4�nS�ihٷqFW��v�H�X���F���v]f�|,�)O(�g�f�U;*��QYY�V=����j۸�R�d\ҹ�i�7r}R㬈�4[	��ꔯ���\�N��C��k��k{�Φ�Z*�S�X��}2�\/��hs5� 7a�\xy\��bǤ�A�,�3�%H��O���a��i�\9UJ�,�jT�͊��xx#u8�4psd�K���ޙ�,5w�E�j�k���j.0�w����mu��t���
q�ˢ�u6d���ͽ:2�	�k��bd/J��.�2�
�]�gC w5u���Q�!���o��:	��it8&��(*���Z��x�0��6��>�&ՓOXռC6�VJgIc=5}�q�m�����@�-Ze�W+z��tH]�e�N��q�>]k�K��̥i�I����]%^w����l)�AK������b%�[lԺ�r�T�(�Ǥ�c��7e������d$T�e1M�CzƎ̔H*�����i��g��-�7�o\��Us�
9�0ŷ��:\7M�k��ew���6�N�-�Ρ�Y�+��
v/G�Y=���_<��&9�t���:�����j+g=sw�D��w�t.T(X�poI�;/d�]=W�wt.����٥6�6����'+3��=Ϩ�����ڪ�X�.�k�rT{�}x*�U��[T�*YJ��,��mk[Z���m�m���%UjT�5� �PV�-���Qe�[Tm�QKmmKZ�KZ5� ���J�m���ҋQJ�صcjZ2�--*+mkKU�j*ڶ�m�(6��%��+cEh�[m,[`��m��bR��	R֕��6�h�6ѢؖT�
��Uk,�J�mEV(�5�P[��մ�A����+J�Vڢ�-���[j��$��e
�Q+F�DmD�+UKElJ������(�����U�B��m���Fգ�l���Tl���ѭ[B���Q���KZ�DJR���h,�JZږ�Ej�h��De���R�Jե���:ټ��1epC��C�u>'/6��2:2�'T�jfFͻ�T��0��$\�5�҉�PL̆aӴ슱.����V�b9k3vU�3�)�M���ʣ�w4+,�U.g6�sv�;�����R��39.��h��ޭ��h���чr5�I�=��=F�����[)�c��;��_�Oj��F��sO!�xv��f���#/�:���Z�Y�/��k��@��⣦Gnkؒ��9�2��RKGGfV?rRGn	�-
WEҹN���3y�G�a;u��wz
#Gհ�V����ꑃa�:��8�V&�S�Wj�}��}�����;�8��ٗjD�wX�AgV��{A����&�i`N�/��u��+�Ղ��z���>������������=��a� ���L��ץ"����sJ�(vw�]%�3*tecZ�#I����mF�5פc�#f���9ѥX��	�]3?mr9���OMw�^�DR�F���Z����_9�u<��tF���fp���|�=B+�.�)��H���\����'^y�q�c/�=3s�wfD��5ؕ<Bh�r3�F�Å�c��Y�0��a�ݽ�;K�C��}�������c�v���h�����&�:�9;V��l2�M��d��xC�+p�s���7u���h3�v�'|'ulTV\���x�D8��vW�V]^s�Ko���o_�E0�-	��:�j&ps���*m�*qבmB��3bJ�v�����]Z3#{�����L��W��U��]-����;���xZ~���R'���F��}������:�qy�׼C���>���;#�<�b��YYT[�(Y���nqJ�6ca�dj�1�λW+�x�*�͊���"-7u����-}��* `ĺc��%=�m�+�g��q��/6����=�����L��~mb^�Ŭ�wŅ5�cQi��C�Ŋ{���8�(5����b·s�7�>��{�^[����d��)���&��>�J:5���s��7�3q[}�� �-�Úm�R��w���e�*��gBv:�K�E���]6C[`��_u*��Eۓl&I{���%�0nn@���\˙�����8蛹�ط�-]��Ĺ)WR �qҕ�mK[Y-�(iǧrq�;y�Ԅ�	�B@��@����V��a"5��|wͼ��H���NR<1�,�H��60*�t'�(�G�����J}�=��Ne:˲�Y�	�u�	̄��/wL�����*��L��.�78���y��9C�je ��L�CYRHl/79��t�i�
�!��[DP�8�����v�7cپ��}뙼��?F��nH�p+҃������A���OV�R7�<��+n_�WQ�:�	�C���1��⇐׶��U9������sh��JJSG
��V���p�B�r�W�Go��ޜ��=Fzr��Ķ��bk���X�F��c��-���t�u=˰ϖs6S�N/	���ʩHU�������.�̔7;ۍ4V�hCgq��5�x����=��W5�q^Ѯ�9�ͺ��Bո*��A��XdnI��B�#)	�0򯹴Z��W{��w:���t�d�ww�u"���X$�)��9��w����F��ں�7�+��˴��v �N�Ή��������G����h�k�a?<���t��y����D��qCў�8�s&d�N�Y;�kHL���{TmġWbU�3�m�d���[�w���%�ש�S�ڋ�2���f�rw��QG	[����� �q+�t't3�c�y#��O6�u�+�|���>�/�`n�j�#3g�hu��p�S�b��;�Rj�W@��$%�e�|�cw2]י4xv$�e�q��0l4,	BE>�zy�궯��l�=��Do�l����䠰��[���OB
����:���΀:{hq��A�__g�nO%�L=�|9�[ڜiA�~K� UuzZ=�������K���΢�,n���s�/R{k��S�KڨH���c�Q��^\��'�_u����ѭ�H��ľ���-=�Q��"hJ�Xe��k�i�ˑ�$+9�q�3�J�5C=i�=ؗ���D�L������:*��m�̢�DpR	�3`E����iSNU���
Y`�[H�j
�86�lɣ���=^�"�M��N`��&�L�̠����э���wTv�-�,)cL[W�_��n���ʾh�$�^�t�6�އ*v6��:����Д���OԂ�q7}!anh�G5�cTS�N(�9Yp��m����$Bb2�
���"GT&���ԗJ�8���S�q�r�9;�q�w�t0�$k�tG#�B��*�Q�ފ��wc�xލom=�2q_�~	j��o���6�ڣ�憸�����f#8�����I�cq��ŗ=y��aX���7ϩ^�9T@j©O=)y�שYg�c����p#�WTv�t�������f��{]�Y���8B��v�����C`�1[-�J1��r�RM�]&�����>���ˇ6�|���%*��W���u9HF�ap2��&��
�orҬ^�6�,��H}���̬�jh�6Ĵ*WEx���d�'�gF[J�-�f�Vy���j�G&��%��7��0m	Um���,��Μv��+�g�''PZ98S��[���	��J�Vlmя%�_b�}�Nvo��ܡG�M�Ɓ����	�����!���:⺋�)�A�M�ۙxxq]7b�
�\���RG����>��uK��W;��a����xOWM�b*P\U�|=ش����� o�8�}rCl˵"W���6?G���]��hyn�=C�l}��~w:�_q	�{�[�HϪt��ꅢƾ�R�$��������U���Cվ���sJ���}//���r9�	0�89/�S�{�,��ǲ0⼆��nW��o:6�'[Gni�Z�y��L��N��6�Ww�W�R�bPW��?+��	�"E͈{��j)@�خ�N�͠�;^EMp�Æ��G�	0o[/H������I]��8�3i'ÔS��TC
utZ���\1Z=�zwgI�o�QV�������w��~m���)�W4`�����=�L�!���X�E�]�Rx%�k8n������x���ZV����ju+s,�28�+�N��3�Q�>T���C=�U���*JjoM�}�;P*z�^��X�k�8R'����0�\�7)��bk�qj�i�PT:���*s�(i��O�����
�;�Ԭ�%6�0)��0�-�ǃ�ls�d;\�c:o�I��a=��QLr�U�*+f1@49\���Xz�ɘ�-{�g))��i��,���<g�^Ә���ҵb��۱YH��h��q�][{/�)��vߞ��&���}|�b�9CE*��D�\7��kK����0���_��-�O��|�dC�ģ�u8t7+�-�q��&=Oz��ݫw����Mȥ�|�5{%v�O�>���;�i_��)���>�ܭ��O�Ƃ�h5<'�TQM|�u���H�Q����[{�49��5vs+�i.�����R���E u���}T��y>�q��_OIO^5��Du�g.J5�w&�2SsOܫ�1#U�%�F�{m�ڬ:�zRb�C�K�VkY:yn�U����3�E�d�CV"�46|qΨ��q��f�S|���l-w����e��$`i��Z�9���NɁ�okOuT_p�;nJ��Č�O�Uΐa���E4{xQU��f,�?V�8�31֞`)��%�]�ݞ���/�=%S˱)5�iִ�7�z:�F��;K����J��F>�:�<��ȸ��ܣ�tѵ��YYe���H��l>�\!ڨ�k���4f�m�Ųs.IR�t:�-��������6�����8]f���S- ��W�#n]��*/C:���*��I`��:��'uyv�J���奋�q�W�������}Ns�g��[9D6֨���&.ں�Wk.[��C1�R�̞!��2�9-Z�!i�8�gG;���5��&��'�5�p�\�5H݁��[����M�β1���v��֐�Y��ڢ-ġWV)W�]�9�@�go�jU�ː6�.�}�@�ߵ�ݨ��eRy٭���=�A���:I��/���v$�.�\�7O�ԩ����ɮVڷl�a���u�^�yA<cӭ�]�����|)<����������6��\��ryV(%�,�
.Ν��F7ޗ��ҦjZ(S��^�uz���3������KV��r���!��~r�Z��)C旑�*}�[ڒ���g��p�5�v�Yti�%:��:M�7}6�v����h^�̽x+��1��8��=�Nmem對'i=�;8gL��|��ͳ(��i�V��/��̗���]5�����U���ip��oy�SMN�k���ncZjg,Ŭ����RES��]VH�ءoL��PnX~KʮXʛ�u<��)N�J��U�q��/�R�ue�Oms�mTk����ݞ$c�Kz�R�vP�_���B׹ѭ�H�|ȗ��g��\#]�TW4P�r/����q��U�z�h�L��:&��������a�z̑H(�!�.�C���8Q�k*�E=���s��.��ov��Qx�F5h#�,l�o|#}[[�����&��Zm�Jk���Us���{��Bq<�]O����%U�q�x�Q��M�Y�7f-�7���Cw��~m�{]f�L�Q��s�"�cy�v�n5���=�mb�<��^��f4��.�|_���Q\m(Y��Q)j	մcF��Ui��<��p�ᜑs�U٠7�z.쒣�a6�m��9�,��פQQ�fW�߳���O�+�i��ݧY:֫���s�iƯ-ʌ��n��|��fv��]��x��;p��^�	�mp~�^W �1�L@��� Y���<����N�.	�o�3�C]t�ky��gh����Dr/ln��R_ftW�t8S��n�U9@��94��Ӑ�)z�B���u�*�P��z�Z��JU��Ex���%�r�>����ye��R��r��� &��֬Bݭ�sS@�ڑ�BZ�.6U�N���@��yt�'�h��:�#}z�gGջ�Q;�z���ՙ\�x���s���_?�j������>��$6̵���Y�U�4[���]�|�7����w)��Dg[�Ws��'�������n;�zm%�!��=� _q�ږ�z����i]Y|�&yr�&Ԡ�g\M��os|p�[ ��(��BF:��m��W.����ޓ�ZI��{����H����j�i�zUz��JeJ
�w�Ɏ���ODO�����Y���������Sh3�SQS^|p�Bk-H�B�w��}�2GVf�~��N�%Uj������W��+��s+xI��Ii�D���`�e2�G:��5��}cWh��ح�řܪ��P�d�yG��9;�M�Xu��ǫ���J�=<ֻ��c#��R[���Ͼ����R}4�#{T��M
�r�5�E4G�TU.Co��s+oa�f�0]�t*�^
_=�+r�@�17U�=e��F<��M�n�۳(����L����C$]�����q��g���z��3lճAg3
�+!V�sZ�e�=D��HPm'��
��{k,���{Ƶ�mH�W#Y�9S�k\�؅���������1���������f���\"�2�� �:b�(LJ�G.�u�8k+V˭?6�֌LrU�uv�2x��1Qخ} 8Rl��짷��W>�|(�b�2޽̓Ew5��F��&��ʅ��ҀY�(�<D�:li��|Ìy�'Wd���}\1U��n�Zj����9f�ި�\9ke7Z�k��b��޲��4�o�u�5 �ә�̺�f�n�?�(� �S.o�n�rëȶ�7�峹46�(�M�֣\8�d湗eg\� 3ZE`}�B�Bw"���P��޾�8q�A�f!7D�ZW-O�*P�1�2��;*0�8NTS0θ�R!���Ы��
qd�!/'�8����A��C'ڗ|ť�j	6���+v	 ی;�[���m�]9�w�ň-��X�A��*��\c��՗T��V�yz%��:�3����)s����I������T��uq44�E.}Ƨv�:{7�u��`%�1 �pvY:_�bSm������O	�gsU\<Pķ-rp_W\ �O>LR�t�����t,�uG��QMu��˟&m]�D�WX(��,���=����g�iY��3%�gF�P��ʝH�8tꬵ��Ķq`�5�ς��)F����1��3]�bʛW(+P�λ�D�;�S�s�M�xԚ⽸n�	�våʢ���! ��c���g.7@N�K��7�N0��i��ٴ��t�}�ͫ�)H��j:!\]9���4oM�>��;��bwH�֪Ӕm�H��}4y/Q������[I�e��,�
�{�!�3f��ج:��v�E�k�un_2�sU�Sb��u�u�w�WN9�c���:�[��[㵗	f7W��	��mޞ��꡹�¹����
DN�hes��+�b;Q�
�+0�J���;0B��#+y���86�:�OO#�^*\��9C�|Me#g*�eY�Ջvi56��2��+��4��Ut��bAu� x�v�Of˂�Y�3!};�q�W����VZW).efW6�2���b�cPS8v��.��j��pf�`'����s1!)�l�HVt�^.�LF����)��5�/4��"�����r�}������߿}�l-�T�[J�6��kj��m��[h�[[EF��Um�#Z��څ���-��mP���ckE�­�Ym-��(��J�����6�X�Ѣ�UQcVڶ�Z��*��[ZV�մ��j��֨��+T�m���U��(�ml�mQ*Ee+J0UmU���YP�U�m)mV+jڋD-�jکFUk-,	ZTD�DF-KF4��,A�c*�����m�m��QcҰ�*Z��Tb�R��h�$F"ZQ�-�-Z�bŬ(������JکAF��F��"�Z$�������U��EQmK�B�ڔ��2�b�JB��-�ZZ��mm��R���Ԣ"[e[`�*�m��V��F��b�X�+(��B�Q��`� �OJ�Z�K�y|��>0aP�ښ�tOY�u���������j�I�z�	���ڹ��X���'@�ȸ�N8TW��y��cE���	sޝc���TC
ut|�T�8�{���s&!�9�Yҍ!�/\��F��o�*�a{����{�b��,9��T�7�У$�}Q�</��]��(غoln�nb<���yM�EI֌����Z,b��>N潡�h�����ż�B��ulF�8�$�ƾ�+m)\��!2�pw�D<ؠ���N2�%�w��Wr���}����6;�+y�ڋt�w����OX{�@r�R���s��f9���Ij[�mdJoZ�l�D<�J;gS�dv�P�Y��3V۴����t��b����5cd���q�V%�w���\�Q\6g��C_$a�T�R����ZG��u^�j�0�֣�젟���V'�������rU��E ���]�J(�w�uw���<\߫`8��^ɭhw��5��cb*څ.jJ��h��`�$���&i�^��/2�/��bc�6�D�h��mt;��y��Ӧw_�^�� �:;�7�:���&rD3ԝs���MUoi'4Ud�V;�.۪&����Ѭ�<�ݖ0�����Ώ�u��]siT���Y#"����1ڶ"ι�%=�������I��Ƙ/Q	�+�Q�̂T�T�jF��̳h�f�R鱪���j1-]Ǚh�}}m�Zp!_ux���ܞw}��J-�t:Js^8�ގ*�C<����pKN���,%=��/n�$
���mMf;2JS@�TFk�c�S��PM}�x��4V�V���79r˗y5�(k���~�ʻS@UgS|9ia8հymy��$�!ӯ�dts�'+Eq�	�n�^U��t�l���s�*n��S\5�x7���֟����v���憸��h�S�T�ú4h]w]���S�ݬ��B��H;�]�7�Ϝ�ʭ��W�r�<�0�H^����/�f��Q��.�b����酷��~�E�ejz�{ϯg��D�I�R������B�����f�+:�,]����;�3oծm�,�K�e@�9�/�Aa�x󧇯�*�{Ւ�����Į��71\r)�/�X$F�n��̂u��!�nl�.���4�Km2��O�/��W)�w�v҄'�t����΍ui�҃�v]H���P�95ɴ[�Nvn��}N"os�bT�֖����;hH�S����3�C��Į�����*c�a�Jz����򞸂s���T)�KB�%tP-+�N��Щ97��l:�[s˶��Q��ɢ�<��S�Hr�ʜO�� ��
ʾ���]ѩ�-MҶ�.�U����c��ٗ~���9Wu��!(��y�3�x��]���#�k��]άܞ���(�FAM�R�Sb���l�L-���L��S���@΍n��+�|�K��L��+�od���:O�9!�c��u#��q�΍+T:�	����k��tFۧ�-�fC[r<��U�-�2��j��Rc��³a�^����QM:]�w6�F*�A�DX�*k\"GT&�����cs{5��f�6�"c3����X-a�:�b�w��v�4��A.}�����W��~��U��ތKs�a�2�dީ�|f�O��S-A���u�.���:v[������e��X�7ʒ�.�w9:���
�])�&�N�f4yI��L��N��{��\9���SCTEWT'1�gŗU'/�;������v�Q������ni��6;T@�s^�Z&T��o5ds�q�-9Zzqh��o4n���i�{]e����9�p����X�����@�)P��&���9�-Υ�صW����ֳzS.�8(�������}թ	Q��
�F�hø��[v��e���guR�kq)\�fvn6���A��
u9H֏�W_`sj�ʹ<ܢ������)�i�yذB��������	��2#��P���V���Ō]$�l��5����&��>�V�R��v�k���;r	�T�X�!=��r��}%�/���~	�����>�!�e��fS7hf�W�uC�9�r�P=����+�Ղ��{�MP�r6o�wc.,P=��MA��$����S��`p�'1���qs�M�Ykzz�U2 ���/fYa��wZoH;@v���!4;�R�n��Sag�nRK1�\f��,Tч��:�c��w���Uۜ�p+�k�g�D]�FX�$����74�ʄ�Jg�Kd�;Q׭�?Ih�
�R��黒X97z<�}ʮ�֙�Q��cYC�D=}��.�!/k�á�/�(\��.��ϔ�r�ݹ�4�P�W�gT�gX��bMC�U�K2�%5�m��\F���ڢ�XM(=�b)��|p�w����f�&��n�]eU�ujҜ�Ҩ�;w�QL�PMv残QSZ6�NZ�[V��U;f�Dc���եuyv�-�G0�c��/͹����X�:��B͛���jeЗ"��A��U��9�Id��t���@��u_��9��nw�s�1��r�y�}������xh{Z5М®�����HeP�g�FI����ΕV��h���v7]x��ڧ�U�
U8˱YIbf#v[K��Z|�c���=M��4�{ƣ�n��;5����VX�J铔tf�������6�yݛeiͅ�B˩�������vQ��ㇻr�/*���n]�O/��c�U��@��z�=O�N��,A�]ݾI�U�"tt+0��F4Mʚ������������Wq<�(�5��N �B:f��鿓jԩr��$�l����v�fv,S�=i���ڹ�穤{_h���'#��(N�3ܥ5�l�څ>�+�:��js�[QuEl����f�{.(p큃o�����⺵��0��b	�܇�4�bv��.J��;��c��!�q�t%(�l��]W��ؼ���'J��a���'�ۧ缈���&�2����*��L�5Wv4f��]kt󳨢Na�Lx�������9F�2%�]"ڞU���P�o���(�	}�O�o���sJ��__7V6ӁBPqi�b�.G#��4�u3L.X��$+:N7���X��j��ae��W~P��3k������ulEfK�X~-� p�>�v��S�n*��X�q��^�Όj�#��rCqS\�����ǕyB�Mʬ�n�L�Gm�u��=9;�Vgm�)z�e ���y���S3<i�7�.��P��c��
�=�e�@>.�5�c�9#�߆��y�����j� ��.Nr$CZQ�`��$b:��*�m�㾐��|#��c����N����I��wLǱ���:��;��}�c��ڱ�`T�"��1P���.�Ӭ�v\���Ym%�6��u0��#V0@䴅����v���j���9�r�? �-���s>��U>ń]p�g0��K������j�����v"�m�V�|�}�|-17g�VU���L-�j-��EߙZSս�ϯg�*�nZ�n��z'��(a�t���nzV��h;�'����OR���9��};���yz�����NR�Q���=�]�=���B��;�.�n$>�N�n;'7ܔے0m	h	�ߤ�����%D���i�v�r�Oy��{�<q�q	�v��S�AU�#�T��M�F��<w!��z�������j�U���&���}r۩|!9���qd]l^V۱W|�u<�����LοJ�@��s��Y]ί���V�i58Z 5�!�N!B�j�����X-N�ZT$1��d�������4*��#��v3z�s�N�w�#�T��B	��A��u ����ާڦ��*|y��A-r¦�X���ںH��|6�8(�w]�m��d@��Ag{�S
q��Q���T�+��>_s�G����8�������sJ���D����8�x�[���y%���3(!��cr:�"c9ѥj�ZV�W8O#��roU�'1r�s���:�I	3'ԃ�j�5��Ps�NRř������J���Wbȝ�Q,6�>�b5����)�k���œ�q�ǥE���&�"��a��υ��#��&sTEWF`ۘ�8{����QV��U��X@�]��6,6��u��gj��s����5&�
�EOE��K;�g�*Ds8�]�7M����v��Ԭ�\U���>F9r����˖*��qZV
T&�V+*�o��Crs���B���nEV�iw1}�{Yʮy��e�Br��b��Vʑ ���˦�.��L��/�N���S��C���6��{�D��G�_��[sfٴ���Zí�B�[LU�3D�\�+�zk\��"%v����<�Ӕ�2N����(
�p��^ΗmU�3fd���|���6�{;#�T�ѣ�)��-�e$�f�kL�*n������r�� K2�>�#m�R�~ʶ�}k�L*��].:����X٤���d&��<�Av���S@�BF>����!���y.{����v�s�����-�)���ŵn�>�W�=���D��yz
޸�K4]zxJ�����]��=�g��(4U���@~��X��&���0�$j�	J(�������_��y��.�ļ['sm����ˣ[�tm3!7:�ʤbF����Gj>νo�]c�G��j��Mr˺gY}a3�iԍFR�	Ԏ�������S�<�v.��S|��Oݰ��k�kh�/��sVNJ8gg��;:(ۑVx�	N�Z�]E�	~���GR�QO�Uΐg��E��GC�˟qC���M��"��v�x�Ȧp2�����
��S��{}ʮg�Ԗ��̩JX=�XVXE�������Ŷ�:**��;_[���۔��r��8�5kw���=QWZ���h�'��� �v͍��}y�>���!�9������K�7j3٘��ӏ9���kvZ���,�t�g'��T�=���d�!�0q�A�/�*C���e��Kʚ�s�+�/�n*u�Op�Bs
���a��{�H v����{��)[|����:��=�ה���PKx���y^���a��g=���Ƒ����:��S|k�kt�7��j�y�H�*�8�ގ,���2���I���W̛�ߋa�G�ک���;7<������ѹ�#�;��'������T���릕��w�[��dC�ģ�t���ާzio-Jb{^�-��FoU1S���&�d��@�|�ՋV@7����/{D��o���!vҷ=�mzF�<$4��i⺵�t�F�Ɠ�Ž�7v���yݽ��>�a��v�/+C�*�%�y�!��׼�n�$�UY���<���6�J���*1)��wq�<�[��[����U�q��c�ΚF��r����i�Ȫ{T��4@]7���q��a���|����sk�����4����g�w�5mXC=��m.�T�ћ{dd�{�u�mݎ��ۡ�aսvоZ,��~A��N��g��Ό��n�@78��n���� "�����}���Q�^��zR�X1�P)R�NG�$��;_of�YΩ��K�1\�,�ݚ�1J+�D=7�+����� T�[Ͻ��JK�+ˏ�)��嗛�Av���HzQky]��[S�֣.�Yo`wz�T��?�!���5^W��W��x�q�#�S�*1��*� w!7[2՘u�9a��;����u2�Hc���wz�.v�o[�F����ߠ��kT�h�i�-�@���ٻ��d���fG�&1�n=��N��4��Kso�Z7��� 3IVGA�2�޴[㯩���X�Q�[\4�%������m�6I���O��`9J-��o��*�ŕ�zGT#�H�gGW��>�	�B}7j�n��WtRV`��Jf�#�xowݹڎwsT�6�����٘E�tܔ-��}�{_� �	��_ÇZ:��Z�Dd�b�e�;�a$��A�yr�b�>ݩq�p� ��g���W�$�'��9��*�sw5�-��D.�@B��ĩ�,��NLMWS�.�D�ʋ��P�j���R�Ƶ`��Q3�+/kC�2���'-u
���b�:ӫG���lI�a�D��	��mh��p<�_*Z�F^�^(�񡻦%��,��lk�?��s��lT(I�n}sh�X���a�&fX�r�2)]f���z��oٗ6�_B\��f��=�SC�1���ł%v`������4�OG�̼��	�z��a2/$N�5��w�����'f�#l�E�Ǹ����Oe^�kki��pU�u�*  ��%�Wm�+�fǺDK�b�p�/`8X���05ɚӆ�3�l�Ƒ)��^gvt����u�s{0��x'f��F�l,�N'�\�Wne�	�`M�d#r��L��	����e[�5x-)s8g`"�;��⾆6P��:��-�vk�8hH��^v�^ZWXr���F�՘B�����z�31�R\��}6m�-��u�Zյn��8v�).f�](9,X�`�جھ�\�l�8Q������䔑�D��<�+4_=z iAg"��B�&Ӱ�4��cv��	���\��kYG5cXsFo~:�<2d��2	]�����ͻN@K�r3;admݳ��u��O;��c�x�غ��*�3#]�Or�.��V�����2����Hi���ŬB��z5aD���[C'^$��BF%���ݰ�9[*���!�����|��t��3���ǬZ#ol	�i^<s��s����^�O7�Bͭݗu�+oC����t�U�)xH�vm=�^��� ��2eaWCt]�ѐNm�WVܫ���3�C�opجB�gP�j��:��}��$��8���=1�S&X����:�I4y*��[����sd�*n�;��2�4h|@�hP��کi*��im��EE�Z�+lZ�m��*V�jVU-R���kB�X���U�KZ��e�F(����E�T�FZ��iD�������-�����+%ՠ�Z�b������%J�e�Q+�"ţ�kT�V�Zѭ��m����Z��
��-��Jѕ�%����V5jڢ�ը�VҶ5R%6���m-+YKKFֵ���б-(�U+B��V�(�V��-AQZ[*#V�RR�m)Q��*�hб�m�
�*[e��V֩UDb�E-�ԥTZ����X�J��X�lmR)KImm����PkJ�ET�Ղ��em�*Ԫ���h(���V�(ʩZ�*Ѳ���b�Z-mh��QUZ�R�6�-���Z��z'fGG�2S��T������f�k��J�NV�5�C�T�Y.E�� �e�*C'A�w�ej5[w�]KnP�27�S&�tkw�+XD���l� Zp#Ḻs�Ѻ��I�R�h�!��H�f��98ލ��P�Zh�A��ܔ��;j��lwj�K�fH�R��Y��d��ʭ[٩��y溜[�V�2.����y�Y,Ee�]��+|_����5�YU��Y*�_*��r���xXN%f��9��f��T8b��n�W�e�ȁ�vz�MYI���3f���fR��@�Z|����v����6�k3d4�k��H�f��o���Jp�Uw�n�Ø�W��-7���f��{Tm�ՙ��îa��m��m�ѲŊ�G�VU S��ޢ��������͗��|lU�bQ��ެ{�U߸S�NSv+�.v����m�c���2&36�Z�2{�RK_<���X��Dv�/ZL9�'��k.f�q�f^OZs��],Y�h���.��u4�	)�>tHe��_tӑ���(u��^9���R'��ֶ|�׳*�,Λfe�2r���Y012tW2	E��v������ozLBn�#�Rg��V��=�K�W'Y���2��
jY4�-��nc{!�9l��	��	k�=���B�]��V��BpU.Eˀ�\s�u�oyΫVS�S]����c����%5=
�*�J�=Ұ�q��ک�`����r�:��|WWo��i{q���.�8�3=R�j���t�o��4&}T�Jd��Y��p+�Ղ��{��|r�W����u��f��ۊJ�.ސ��K��H�����"�3�[摪z�n �_6�q>��X�,�m���#
Ւ1����os�JU��Q��5}ۅ^wd���Q���Q#�ջ�V$�̚A� ����WA�:�oK͝N�7��8������X��ӊm�X��k�O�Q;�td.Ή�Y�o�N�j�����*��8�~��n3����.��}w���Q����s���R���Oq��o�]�P;��m�==�:ʬwf/=��ݝ�#`ǫ(��w���i-�*�@yV�6D�[�w�kw�j!xI��<Z
�vw�5K'+�(Lz9`� ]����a���;�VmHEl �$,4(�y2��3����e-��ѕ�~U�5c�P����f`&你�Das���o:ֵ�y9�f�k0�X�1�gL�`�s���]�-���yi�y��}�]�7��]��9ّj8'�s��{_,�X�{TCw+/*��*ri�2�����rw&-������uD5���`q�!=[ٮ���ƄV
T')��F3���ⷕ��4�]��⑞��)(jg�
�䩯2������)�G A��N��!��1����7p��$m�l�6��N��!4�<�X.����SDv��F�v�tnU.=�+�]'T�	n(��S\6J������AnW`��]��{��cGl-J��6�� $����[Ue��a0�~Q�9c.Õ����s46�_Kn�N:5yHF�ԥ���}0�I��X��=�y�lO79��V�Ѵ��r���H�u	l���͜4+��^��3a���++7�0_#�y|�]h�̂0�X$cF�TN�b���Ue }Z�N�M�/�W֎#XFS���� &���fmO �����A)G#<�}����yH,�-N�fmO��ܣJ��G�ރj�8�K�Zh[_z�T[_�����u��W-���M��4��Ԉ����v��S9�F�<�8"��M�X..�:���]�\qF�cW;XD�K�v�4�i��՝.W��g(ʪћf�{�vĐ\ˬt:ANN7�z8���Zh�A�;����1���޼�J�E�$�U�ZS@�Ts����!�TCd�y��R��ŉ�Fkv]�w%�lN���&ۓy�v��*��-����q}CĊ*M��e�3�=�r=N���]�J^�	o�'����Ӥ���ɽ��9���a�h>mj��;������h{^Ѯ�0���gx-�Njx]F(ۧ{���v���1�3���\=����pk��/6+�����i�ɑV$K׼�o�]|멑s�[uSk�a����&��0C�-Ɋ�>�^�}�J�s4����)k+��\�"饱)��n�L�v+.ن$�R�;���i��-�/7��ܑ��P��c�&��d���CN�A�Ӭ�PW�1u�w]>�l�Y���\�\�m=荧0��5yb)Ǽ�_G<.��t�1K���#�r�#�F{��u��|VTU~e�����n���=��S��<�ս&v������b��o�9��v�9O�ηm�v�v�-��'��X�wwC����T��Ԯ�Y[g�פ	�G|� b��6:�{4v��ny-��r#Z���p^K�����C闲�(���We�m���\U��=��W��K^GZ�'�����W���5�^�����\)_o��KRPy�_��>���Z煥ue�)�+|r�:����Gu�|w3��Ao����`�!j�����y�2���8#2�%�׎m��O����á��BFg�;��j�[�4z�����:��Kۋh6�	�5���L��yu5���2Anh*��]�Oyu�����gV��wo�n�dN�����j*k�2��kqث�j]�MRuѢ9$�,��}u���|��a���.�#�F�f�DU�R���Zb�+�������DxNpc{>IiOa���Q�sZ�6�D.y泝Hm��]ײ�o��!�3T#�BСz�B�u7il�2�)�o����8j���4')��������D޹�/�rY�5��r�o��W�݇L*H� w8W&�6�zۥ��&wq���]���c��g^�r��S�u�"h)���9�'a�w�����O	TR�{��a���3�c�
�t����pk���Ť�Iu�|�v��Z�!J3�`��-�H-���}��K'��uL�F��YM�)��㕯�z+���r������Ws�
�,�a^W��}|�*I�袆n%'_Gг�s�R�M�R1ק);�;��ǀ��3�Պ�pm��w�bs^�Y�i���۞��J8��6���E=� �k��W���j(��X�z�K���}�5nܽ�jz+�r�Q;�`Ίm�>���X��wL��/�����U"��4�=�8��ٖ)�v�4�V:Mb�ei�_����*���v�=�o��]ά��{�������o��LorK:��� ���<-#U�8�������sJ����2o�'W$P�ż� ����6�� #
+�j����q:�{
� Z�33��6���x���MR���o�P�(��4{t�߬�%֞�ow��V��4jwtf��{�D�2蜳��ݬ�������i�t�������7[�$y[�t��y�,Ûz�fmT��uɍ���]�7�i�� P�����v�=�y����"Z�~�V$�̚A� ����RY��z_V���]wZޝ�Ǌv5E>N'@ma؊�Mp��SU.�M��>�]v�ͺ�@ZSGK����(�9��|.�#�B�6u���뮔�s�ͧn�TF<hNbWW�v��e��(�l[nh==��Ogn�E�f�{�eA�EU1�sC�EP����~�uv������\��z�Y��|�YJ6c��˼axo��j�W+0JٶU�YU���2�j�(�;q����Um �h����{HoV�k��!���0R���f���+ؤX��guK��Y8��5���.�)�;7<JU��Ex�������n�̧c����EVg{�:mQ��.i;��YM2!�b�!wWXMOXj�tx�f�wf�f�HR�u��9�b;��I]&���ƠY�8�5l�1C���3�w�)�
y�-�qԼ+h�1VY3z�G/�ل9]k�oUBr#2�7IZW�oGG�n)�Uu�u��ɲc�^�3'A N�ݬ�	�*�r�6�o'�N$=ى{J�VOo�S:����޹���:�-t��>�yʣo�sk�*V%71n[ܘS�2t�O��H���BZQ@�D��T��Ʉ���M]]P��to������P~��K_뇂�CS*F����}�����3����ᵶ�l���g7���G�z�H�)�~�1)��Kf�͙�`K-M��-Y�Q%��瀴����//����̂�j�#]]
U��Ug�Ui���]A��l�\�tiv5s�MWK�v��
�:�Cr(�ݽL����y!`zN7�Ij�}i�C��b7���O;!���2u�,u/ҟeK�e�nh�TFs�c�S7
��"�m�����#�5tBqS�"lp�SV݊��v��*ј[�/::���1�s��=SKOa�&v�Pf��U{�:���X}��5.g�a�/��W���@������`�Z�����W384=�h~���e��/� D�q���e�2x�o����7��V�;�^��ף�Ss��ٷ3T.��7NR�N�jI$bӢ�� @jF�k��#��/��5�(ǚ���t�K������Q�sx���g��f�`�qּ�%9K�����Cz�����t�>9)�b:��H.��G��o'a��!�ؓ]�Gظ���d��t~��e5������Y:
�(�5r󸨷8 �Bq��٭�ʦ;7&�;��.��y@l� 1'���Pݓ�aX�G��Ӏ��5���]��8�\O9��L+�Z�{.ro��!g��;�
�u
�Z�,�릘��_���>
yI�X�,�)��&�5qsKs�>�;6�<�[,@��T�v%+�@O�@�\"�H�6ʀ�%	�����5�R��F[��"��P�ҙU�\.,GБ�ύH@��4�z���v�]'��ut�/lz=�
? |%�p;,�Ns�*-�]M���e�Q\`-r�Ak#�3GS��j��JV)�����Ct9h��{=sŊ��)�V�i�@V��߱3q@��g/h��fl���� �X���*b�u�j O�R�{*�tV�x.:�rO��n��8��)I� u�X0C��Db:.R�H��:ۡ��/�/x��\��G�����6e��.����%s��kN�M�x���DU~��v$B���4Nt���Z7m���L��YK�9Qb4-K��c�f��=Ozk�14��Jқo�T�y�[&/����(��H� �T�H����
" ���-g>In����=[�t�<T�Q�Z>!Ԟv��K������"��DaO�t�҅J��;���d�qE\���2���w1A:C%�EE�/��49�qv���x���JЄWw�1��̭���j�Z�/٤t
#�s�t�cՔ|>�v�f��Z�(1["�����^��7���Ef��>r����&3���Ϩ���YXH��`F���~�Gd�d]Ftf�ެfҦ�����q�5�����c��x�:����#p��)��^[���3/���*��W+:t�⇪�Z/j�c�?(N���豒�����8�3I��=��9Bܤ1��wk�)<e��6�p��X��-͞�
�Mz�e�ҝ�v�k���S�Y(w+�O��9�(��u]�GH��.�Q�:Hi�Q�R��Z:�M�R��[ͭ�}��}/��p6�����ʌs��lN�*'���/j��eE�ݞ��x(�;���y���*�<4puo��>�K�UZ���kݟ�ѿ����o��{�hB���IO� IO��$ I,	!I�`IO�BH@��	!I�`IO�$�	'�@�$��BH@�BB��$�	%�$ I<�$�	'�!$ I?�	!I��IO�BH@�RB�� IO`IL����)��`!V�-��8(���1%}|���%�"D�!$��UH���*EQ"R!J�@�H"*(J%H���UB�
�DU(R�TQ*�U ��UT*��P��)*�N��Q)%kkV�I�_Z�%"�UJ���TUH�)��T��R�R�*�E*��&i��H�JB�TP�(�)RJJ�QE*���Q�$P�����I"T�
��H��
�P�Q"��$�T���d�U*�2�  t;Z[�)6���l���� d`ڨ [h�J�6hHX(�U4�P�b�E*��-iM�li�&U*�@j�)P(*J%Z��]�  ���S�l���U�QZa+ )B�h�U[5J&���ۀ5�3hij�F�CI���DHV�EQAUT������   ���ZP��b�
�JҘ i@SZ�e$��XCM(�a�T4�b��СC���$(P�C��p�CCB�
 ��K�P�B�$(Pq)UP
���PT��Sx  ���(P�CCB�
��
(P��А�'p�B�
(hh[��P�I�
��h5M)��hТ���*�3h

��e �׷]QU*�*����("�EEx  ��(ѡ��hh���ڙP����B��,� �PF`4 J*�U�"��$RR/mRR�]��  �P�4b�P�"٬�EP�U�hX �%@�PU��
�iKV� 3%T^��� DRR�  �EU����4�f���KE�2�AD=2���f(
�Y��M�
Ʀkll���7R��E�ʪ�%�JR�$O   ;����*P�m���b4� �`�*���ʬ ȫԍ�4ؓ*���A�CF�ضM�H
���eB���R�IR$�%TB��   ���4M�4Rʽڑ�
V�5@����0i�����-��[ �@�f��Ѣ�¡�()�V�0�U(Qb��%A���D���  r�(��M+f4���m��)SU6��h���@���*���L��F�Vɘ[�`�lȵ�O@2��   ��a%*(  ==D   �~%*�� �� �Oޡ6UU1 &�H�2�T��d)E6�%I�D
g�� ��1�{�{T������`ݣq%κ�g�c�b3�x{��zOkԿ��$ I7!���@�$���$ I?�	!H�B!!�9�?q�(���!i��񂥕�B��d fP1�;���	GJ�)@[�F�ʂ�v��
�?b0������@6���N�	K��wl����!�;T�D�P��E����@B,�إd�bPl0^]b�D�pdR����5���[�A^',9��6$�UƓV�r�xa���X˰�RE��E���L�?������Е����uVbu�L�`i�&�Ӄc��:�����07L�%֋0�5nDS%g�0�YYf6䣎����hj�<N���j���YD��mV�Czl�BngI��+>�ǎnD)�W0�0��1�U^�V�<�1S���"�<�'{��(��]g\��Sa�c"9L�Ur�֭5.��Q)"��ф�����������/��� ����:nd�Lk/V�QZwG��7���5��	��������J��E��oj	�+nP�u2�(��q��hͿ�����B��XA!��L�h��E�$��GF���ijѧ^Lǔ�y3KR��<�UkmP0�m
�P^��-m�`�\DKn'��c�4��;����亽̖T+b�f�c�wt]�V-��[�y�-2����YYK*�g���
�3�cMfP�q-,���%YǗ��ԝ�Ӻ�A5қ`�Z԰MN!Б�7Y�g���C[*�TC1��BZ��0�x]��I�!�#�e��&,�T��tV�l;�-�e5���D�nҺ6� '��X_ԯ�lQ2l&'d\ʊefӶJw���AU��p����`��7R\� e�����Si��#ݼ�*)���)w���a�Bl���P)�.�2a9����o�!����# /9I��+�̒:��+��Õ��T�[g0諡�i`U�{�Vc2�iAKyZA<���d{���IԋSԡ��7��ECl]��ݹ�>�Nm�ytV�n��e�����Xd���b�ҥXב#y��n��^QV.q^E\nj	I1�����7uB�;QJ�&�b`�c���Q8��q^B݌St�.b ���  ��̲sj�G))M[����S�jGuH#N��le]�ֱ�u� �5�և1���^ۤ��amI�lI���t*��l��y�&k	BV�Ԡܼqݢu6�HΝ��pjR��Yvr�L�pm=4�ɕ�����	ť=w,��:ȥb1C0�7H:�¥n�Yg0=��9�"�.���ƍ:_6�c`�pc���̫e�4hq�Ͷ�b�5OQ��[�uax�Ő�֣P$1H@J�.�+o�Bb��!�̻�T*�+j���QV�;�<l%R�.
n�ɷl�V���6�̤��.�ƥ�
�M��7��[�n�&R�4�)Qn\�5��@�~�(�j�8�%�1��"b�X�h�^'-*���s��BX�[*V��CVmVMs	IПL��uB5� A�AV�:�n�@1(�Jմ,���Z쟁53Y^j���	Y�f<ۢ�
G�/H;e�,��Y�p��7���N�<��g���B
�*-�1GJl9������ثh�ymcՍ3�h�(m�y�/�x�#(�-�aV�c�Y���T��5��f0p�c/@�fc�Y�V� *�#Z�vӥF�6�S��|6*�w��F#^ԋl��ѓ����OF�@/���M��ʰ1;ܷ ��y�hF������(�6�ZՌݡ>�ẖ&��,K^��Krd�st�����]\f�*����֣Q���h�k��+%��,h�9���
{�I%c<�!���J�.��9L�D:k".0�ϣ8*!I^&j߯E F�â��!�BD�DcfӼvv'�)P)�D�zR5��kHz5�
��x���6��gZ����|����Z&͉-�U[bl:�h��Y*bQ�ʗ� �(���T�Z*�bL@1R��ot�����W��bw�b����ZѺA7X�:�ə�����.��t���O\����oHi�X"�
��A��NVʺʑTG��p^�WfMPܖ����[d�B-+]��xe<F�n�2�ܫz�L��)�f*�)ړs^1AV��b��̡�a'^�e®T:cg/U���Yن��N���ƴ�P�Ӱ�ΉX��.���YËGv��cAm��mk���օ�e6�7��8����+�l�M�/�'f�5�T���$����r���Iͨ�[�Ie7�z@�
�"2�B�콍��4�3I+7��7	��Ǻ��OkU^��b�w��t�7���^����-b����ʎ��93Ҵ���ڹt��Y.����%hYDZ�KjV�VH��5�:��Ē��m�X�d�j�Zٙ���ŷ�]�� 0\�Rf��J�T�6�a�S3�wZ�Y��Z�K�r�fܢ�̇v.����X�;����4y���k2���q���+#�w��n�šP���J��`���]z�T�յ���vQ��+��T��tokm�1=1c��)b��@�� �iK[zX��k6k2,���@]�r�T���bki���u�LWքy]1��fКV��ʆ��ɪ��	�ӛ�
wۤnȚ�dh^�|�A *W1f����(+Kw1�SM�`�qlxV�1
*�n�j�o>�y�e7�Uʍjx�c����dH-(<�8��@����Xѱ��4$��u6���Z�2��Z'�B�:���.��u�������{�>@�s3A�a�,���[���s$n����Цeb�\�:�VP%���BMP�5�@�y��j%�IC��n� ����n������ �k��!XE���NJ
�����M86�A��F��kv�ve\��S���F�q������D��������+7-[�c2��e-Mn�a:���5l#[֯r\hk��u��\V��Y�Y����C"��GGb�֪x���0�^�R��Q�ke��!%�c�,�yzW�"Π�Z���W4Լ��Dͻ��N�n���&}"�֊���.�mM�5��*_B�R�
Ƨ�!�H̻��F�ISJ����`Exn�4�0ӈ�B�'Q��90V9��;"ma�{�F@{���f�-��a$�U�ܥ����,&��c���!IT� �[�wa�ʕ/A���0�7��YO7�e��[Ji�#��z�t�����5n=l�ʻJ��Uӵ�Im��ځ���V������F����2��Mq��b�iB�[�H,���P1���iP��)m���t퍅��揵Q	�hau
+	Fΰ�e�֕��ұ�|ң.㔄Am����X�;$�$k �!���^�	n�m��o��WXJ�����eb&vV��i�IHqPZ�oF*E��#������Q�5{��W2Ƥk2enDSb��Ln�6F�^��H�˦K��;���'3>C�c`����Cu�H%L:�r�r�*i�SC'H�e�kou0��&-�ZQCGMn���dج;��z�}��![�v)�W��:�7'Lݢ*�lc��Ԇ˚죢[�4�
x�����a(%P�u�f+�*.پ+���Dr7��Y7�I+`�uou�]F��#8�:�Ubt2����ux���7wSk5W�nV��-��n�8`�©cutb	B�ض�� ��&M�����A�Vo.�^�B�0��c��g�|*��nF�	�[Tu�屹qƺ����StY�X�l��oc�Ӕ�'
���XњeB�o3Dm�V�]��u(�0t�q�kr�������N'Z������ӭ����#aL�wz� V]8t���j�*f+�Am����`AөI}�ie����#D��][����J�)bfͨ��6S��R�ZX[/M޽�trT Ҩ�k5�ߞǔE������ԧVu�%ecf�2AT�Y�x�!h�
���㳯�/m^'6'�]Е��7f�n�d@-�iP�dD �`D�VKU���`#V�xl��L�����9a��rˬ�Ԁ:R�\.�*j,��Ln<�t��PFf��6�mK,Z��E�.�Mؕ���X94�ީQ�Œ(Jܷt7qVm���� ����� `�t<���7��K.�6��Jd�6��Y2��/`��RG*L��;7�(´��#��v%\uv̴�7��4��+D��6��K��b�9�����4�N{�.񜻭&ĺv�ղ�ץ���ژ�5Nc&!,M�C7	I��[��n��Dh�����nM��(\Y��^m7���k��;Z*C!+3b�K+N*d��Ð�y��7������fĮ2#��Jûݷ*�݆����wloJ��9`?�$(MF\�i'R5�L�JD�+���sQyF�7GMf팥��ʰ�{I��ff*V�E1��X�ީI�Xv)"�WY`S`���B7�d歊�[��w�V9P�"�a��JV~F�Y�P"�KxB�nf�3lQ�7�^�S�c2�[sFJZb%;qxR�L*�dв���T5�<���Guo�`fQ��3�d���.RBm!V�*Z��*fB�8*fЙ�i�f
"4{�Y�J�9n�g�TٶDb�v������2=˥d�n�b��1Dش0�vf"v�����fͬ��P
WbX��ʆ�M���T�ޫ�"���2��׭`�f	0fܥ�j�L�B�xtJڽ6	$�]ݪ�X7 ��S��L�ED�H훔VX;���c���#;�CoCu1�
[4�����@�w��-CY4Rt�q�k]�a/~���=�5��KZ���1�(k�I�K �l�.��VMږG�`��Op*�HKa����j̲t� *R �ܹu�B�V�а4��18���LU��Pٙ&m� �B��F�Y5y�5v�7�
��#�	�{[�6^bwW�<�n��-�&�5����uJ!��l�7P9�d2R�UmY��@D��YPjݼ�E�u�#�w�V������4�=DC�3\��Xq��$R�2�:�	r���j:[ܡ5&�����P��h��))�Te�:�b��Ê�Q�K4��Y�rӬ�����86^�?5S[�Rʘ]�Y��8"�K �K�M�@��w��ʹhfۨ�
p&��aV� ��z^�r�>�T��[�D.�8�kZ�j��J*S�6c8�1{%��=.��l����Ռ������q)���(U��)���{��T]�y�PNcwF�w��2��DT���A-enlB���\�Rv�,l=X��gC�7[�h2ḫc���e�Y���СBR�X��A�����Q^n���*���n쁘u���
��bC3N�h���@^ �M	�nE�K��R���X� ����f-;@���m���+9(%������i�r��h��&`��V��l)�����D��&0�k%�VZ���[۴V�cq
�ҙv�LJټ�e h96H�d�����&�mZ�46�[x6��3R��_³[�V�Є�U���2RZ�f�ĕ��V����1C���#��2���IM�k�)�WNVN��*�y{�̢20��dbDӁضE�"�^h�Ȩ�I�g�h���d<x�*i���\N�kQU��ں�%E��)_�3*�J[XVe�n�Qp��l;KsK�F�C48�� ����6:vF�l��f���h���A�% ;`�w��V� �+S��K�����6��B�[q���Q�6���չ5T.�Q�Q�3��a9ZT�g7�T�x����5��N����4�1�Isof�r집�ye��ύ�_Qh�عX�b4�+�Ō��`�&�۸L��̫d$��*֒�hw�:qK��,���6�a7z��N���j�-K]�hZTZ%4ZŦ��r�m�T��}�R��*�\ڒ�Qq�%�HV`W�UQ;6�h�U\M0�v� �I�YĶS�W3T$R�t���ۣ���#[�Y�*F��bCd84HሥooD�t� EV�����.�3��יO�b���N��RX�V���=�R����(Xc!zӣN�AIV����c����c����j�.���q� �R��++��*̬�gU���b���|�ָ*]�wf^�*Sn�T�)]�z�J{��mՓ�DC����8U�*C�Gڀ�fЏ�M�9�-1V����)�j�u����f)���
���LւB���^�.U��/k����!����{B��6�R�I��)�1Z�6�l(N�rԷ�nn�޷�eȭ3v4P��隈]�V�	Q�XͭNK��ˀ���LMʰ��d{�Z���va�0���V`lR��9>crln�a,�4vM���R[�ՑVqfU��i��Iso��nT$S�/!x!��df:ypi�(�+f���]��ŋ�Ł���d�F�B&ڳK%%�YC���j����Gv��[;��V
{�䠱űi�j�vݱc4�W� ���[�H��ʬr����1�W�h4h���MZ���#;C7iQGr4���6k�$%uz�L^",��	���X��J9�i�mT3X?BU�;�(c ��W�r��͟Z՜ȶ���[6�^Z�pm h'Z��CKS4aL�u�U��Y�e��Z��k&	q	Ql$(vT�n:�B�t�3J�D�ɮ�\٥f���ۘ�x[����,=�)��c��+��k4Jsn��ȱ����b�{�S�������Q�����"�j�2L7Y�����,X����G�O�Z��7��-Y�*p��P���. k/,l�u����*K0 *t{��ʉn�k��]�ݳ;���H�9����4z���Y�.X̙g�Y���
���&��;d�en�a՗�z�3��!���;M�$����
�K�s�}2�{"b��v��w�ߎ���5�'��!p^�qyK v��q�)�H�89@IH�ejX�姴�*]�1��9|s�r:�GK=DI���^��s^���}Ӧ����sN�-�|]�c���V�+���[�S+^K�W�OQ\�R�`F�=�f��.��k"�X\;�@ސ�j���}�r2���`#	`�ɏ��tY�u���lk����ë�7��U:4���bޖF%��n�|޵Y��mD�H�$���CI|�ڗ������9LYf���i�pn�� �L8���7V��� �A�7񚉁���bI��*3�@%����f���J�[ST�L2 ��d����L�q�*�L�"��3yk����`��eI�i���gR�}"��H�dv9M�5�6 {EÁe�Yt�̧@H�-��ޮO~�Z�foo����z5N�Gp�����\���D9���K$]�6��sA���ɇҴn��P�e��5��ٷlc-YxX��klʛ��BkO(u3$ӉCΎ�}]�J��>ٽ
�9(�/6W.����L{�;5d�t� ���W.�kc]H������+U>�l�p%ʹg7�đ�]'������/z�I�x������3J�;�	R(��+.�۳|�"G6���U��Z�^�]��Sz���VQ��gV����-�v���B����Ѥ��elTଗ�C��*�Jޙrn&��l!K���սm�d���\O9�ޥ�3:.��X;p�t�ľ�Zg��ԯ�<���ϻ�{�s~j���u9�֩��}�"Gb�R�*k�2�^L���jD3	��z����K���-�]).�O����ok5��Ӻ�	ׯ�����5�|�o���*.�s+g���]��B1�ѝ �Hfm�.�����N.��I�̆ucx
�8��7mu�Q���{�/R!g��N^�VVjOVť�Wc�>������;�Z��{$ym�=�ʕ��;[λ]�e���cG�l���0�Hp�B��2kU��u�]��b�ٮ(s)�5�;č�n�W^�c�:�^�x����NL(����Y#���d���Зn�y�����n�ŝ��Z7]8�+�¯Ci�6�;G2l�0k�䮕�U�C��6N"����0N�����n�A���/�]Ww��ᬬ�6.��͎Z�l�Ӄ�V�:�,iR�x��M@�ô��q�Zj�,�|#׳jv�1AVc�;r����av��f좐�zIV˕y����_y�L��ۏ�^��n��TT!�M��-cp2-v�ӷa��[�J�wA#��(Z �!�ԥ4v���s�sqf# ���BWx��}g��u��ևhDH���o:���t\�R�HkX���ʶ���6V؏(7�0����yJ��wU�f�6�V���,�N�hQev���GR�.��ɻ1�S
�@�u�0�˵J#�������"�&=����v��O�u�/Օ�q���h��Λ|��ѳD��������aA���k�R\'=��{�V�巓NdX��{,1{i�SI%�Kr�|�s�=��`�jf]vWm��
�z�D��л��s�v���h������t� Z����;�S�b��cMwvo<�W���W�u�V��J�˰��n�V�cU�������A��ts�X�r�Y�/*ه~*R�;�r������m�Wc��So�(l���o�!�H���r6����j::�V�B�=�;�S�o�y��ܗWFQ�͙א[j�e��u�`�Mv*�8��Y�76|�9.��ƨ�?6wn��B���Z�ܡ���U.�#sf١ϳ2�+L�=v�v�"�7�3����k�������G.oǇ'.U:�%pv�������s���r�9�7&�( ����T32���:q�_+5���<��E�ݵ܎��x�6�Qul�rW��j���q���Ջ�Dv��օ7�g]��Cac�f	�`�okZ+�陙96�w���y9��6Q�qrhf���'l�o��Js�0nY�㢌���\+�d��X��z�H�HwԴ�)B�뮂�p)���C���K;:\R�QU4�3!)�nͫ�����YX���T��������}ݍ�7a�}�*t�Ov�gb���xі�![iwr��,@��7v��3�A��U�o$�C:6ԎCAC���i�,����E\%݊IQ��l�8(^
���K��OF�R�4.32��B�~�0��u�o8e��>ӵnŭ�\]�3����+O@ߖT݁��J+4�� �ܶk��J�i�{4�VՄ���#]n�zә��=y�^p.T�i�`m���9f�d�\�A��&\�V���e�-�z�_$��a�EJ��m1�_�I�&:P�S�`�rj�"��v���WY}g2�gR��[V��&��w��.#������t��O�Úz�d�Hm���r�����Ǫ��O�m��@őQ�_.s��=t����+���׵4pAgHz��GR�]�w������#�n�逎�X'�3���BO����o�v[W�_&/�ⵓ*fN?sS��x&��0���XM*ӽj��j�id�
��Z�Z�9���m��8�Yt�׬�.N�f��0c��x�=V	DX��je�:�@�(-��(\�����ڷ���I/e��x.�Ѷon�PZm��Oe�kH������~vX�Z���)�펣�u���<��C���ȳ�I�V������7�J^�/h\7����0XBźpl��aѪ�R��d�B����#�\.�Ё���m��>6�͝���g�J�L�tSަf���k�{���/T�vm��\�3��B]Ș2N��,mŴaڔ�4^z_m��p�j��jmH�HxL\����9S�e��V�[]\kgd�@���$Z2#-MU�{C}���Q�C�\1�Z�jB�lV�
̺�g���� �1�ݬ�k����ܶ�+�;��:��!ɀ�c��dO�KK;����bl���*e:�u:Z��mH��i���0U�2��w#�,���f����H��*���GkG)�0�C���j����hrek��:�;�_fǫǩ<��sH�J{�p:���Ԧ�0Zl�"�L�/���Nb�וֹ�т��F1
�H�.����J�ލ����dQ�#[��H\Z�����]���������<�*��u3�(�d�kH�ݿM^��x�����i�
�Nv�Hq���;�����7�U��$��_Kcv��<*Պ���k���C����M���\�9kZrc�c���Wu��w��H��
FP兘)s	!I��b�tO:3{��V���헛c|r#'qB�����xe���r�Ƙ�;����զo;���)[B���Oiu�+��T�7�I^�,]�<��l!o�XH�{�}m��8 �La�o�2jb��2��;��k�s����t5���/oy��۰*��m:KV�#]K����1:X�-�[�Wh��p��ؾ:^r�j�N4��y#㹹�_^	�Y�U�$�=����E��)r�qk��ҫP�Ϻ��F-��5&��t�-�Y�wD�8�+��:`�Evm�LV�N��fuI��늃o��^Ӽ\��H�o���@lu�2Q���y,J}�w�øo[H5���J�,�ťҶ��)^t8�\���K��]b3pV�t�f��|�Rt=�-�S/erS9�
4��Z#ot�%(�/�z��N��:�p�Gj���1.�a��$Dʖ�uŹX_22b<�΀��cp��^_.�6��J��0�3pD;����\Х̎��e���-�0!v����A�;w�BNL�4��a7\��XaU9.]b�v��f]sٌ�G+p�n0Ud��A!r���8t�ͥ�M We��Nf��kO�k8�MKP��r9\�K����{0�y(���ʕR�*J�5��}b��2:4+�t�.	�P��.�J�z#�/ �t���gaC;k�]�T���*R�o�w���B��Ԃ�,�$P�2���R3KU�=�pɀԂ'�v��[��:�$#)�('�q�f�I��V���>r�77�_B+�ۦ�� �N�<VJ��%��N�A��U�VFc��z�.�vL��R�ak���vP�`=�%k��������� ���7K+��4M�H,���:@G]�%���ܲ�Z�%�@Wk��ek�N=��ZO
�h�B��u����u�:��������z�C@�쭽6��ľ�kW-��sVâ��EWt�3��x����i"�l�(�I��ց�+����H�{΅gJ[�HU���as�m����Q[D�|�]�������Қ@�K���M���|G6r�ZP�|�������e����脕�C�y)E`�v*T�Mc��7޽ұ,��T�>�ݫU�l*�n�|U+.����3����-EY����+���A"�
M][9�L����Z1؝rk<m�)�;�:����HKv&]��
�飔P<��^��nlHvQ��m{u�լ�X�h�a�%����j\��w��u�cE�\e�j��buu���"�����+{n�u��n�x�\���:��jB}Mu)/m,��"�wHc�l�0�F�N<�c��!�)6xEy)&��қ�.u�#)mh�M��5wR���gH��ه��/�����xw_ί��Ʋ�h����/�][�B=S�1��1�u�,�ǰJ�9�[��M���n������s��V����N*g*�.�Ù�����t.�9����n����j���^��U���H�>�0
a��G.��&ή��AS�!��'�z@΍M���狅�u�����`0�j�I���	k���e�,�V�]f�]��,�-��{»�27����4[FVl�5��ߵ(�;;����wY�vA�sT�%�"��ǭ��#�Η�]]���3�'�3��(K����i\�-X��lϘ��J����8�M�.h��oG��X������JP�:ޠ���t�.�\\]&:b���z��ӗ�ς"+����Kz�8��mD�<zL�;o4#�G.�QU��r���R�ԍ�B��Q�s���ܣ5���z������]�:{c�@e�rႚ�������7;W$r���识Է�F����v�*�G�=���Aĺ��(��=158������ّ��\k
�8֜6�h��io�R�]y(hy�5���azyk=����A�y.�c�.��55�C�H����2-f�;��iN��T�v�[%l����m��;GUM��dh��e
h�0��33�h�oE�εJN�p/.��!D�W�hq]��Q��)[e5�ة
'N����ۃ��`e�����1��f`��N��hU0�o�W.*�b�&��T�\�n��SJe��e��\�EQ�܌W����D�޿7}�oe�zN��1*�X.�L�&n��Ĥ�2Nܚ�\�/s�q��X�  �e���cZ�mk�Cܸ$oo@��ғU�O��S �L���� �[+1��qy�U�������Z3*w!��B�XԼo:J���#��k Z� 7h��5�E���'y׆�uC)<���,ͥ���3��
U�T��;'5�r��H���]�t�6������s`s�X��Ί�s�Z`N�>'\Њ=��M��5ڟnp�Z��HN��K���tY�9�ś�Ǯ�0vK��l������U�K�%+��e5k���U�;�| 3��B�őm��A]:��͘�Y�r_E�{Ǒ�˧Yz����!Km��M��7;�<�r�M���2�Tw�]���UH����&�Y}���/���ǰ�g�k�^[۳�����ս.O�r@F!��.}����ou����[�6Q���la��ZU�{Mv�G�q<w�ͥ�Di��F^��٠}Er���u�W�|���qe�ǀ�����j�b3�J��}��v��V�<��̢at��M�[r��V�%K=����6��ߍ��0FjY����ٖ�u:ʱY�1R����q&�gM]��)�Y�v ����<��p�:�8���q�}�[��@9�xw9��:7ŝ�-�4�[���
�3#�7Q���V��)��yN�����N��.NЛ9oa�Wn���;��r��_��ǎ>/�������řS,Šs6�#Lx�v�c��R{%��t3��jYg1lY����� ��ԩ�5�*��l�ţ#����gj��uu�p�w��"����^]p���lA��S������t��ғ�DC���<�����u-e��&1r�IM#�-��M<}Xb����9��R%�7�#��(V�nI��M��z�s�9��L�WX�w�
�p��$`����øԐ�R�JW��H�fa<�9�4J�2��d�^�ҍvP�ʍ]�;G0K�v�ԋN�(m��E�b̬9ZЄWY;��!W.ub,�N�5��ó0N�vLR�%����j�rS�jnoX��+n�YyF�`�١o6�;�_tlqmmz��$]P_,�{1}�!ܒ�^�+j�R��jKm�!��յ�|��N'�iIGw��u>8��v��oq�.�2��/3]b���<\�j"h���g��9'�˻9Y��4>�ٙϳ���j���"�,&R�!��ia1�'S/o���c�8�|k/���i\��s7���L�]��&�g$�N���[��}����=��<���=�|�������&����,��eV�2H��V��GNPT�*J
���S�`W�ؓ���B(�q(�l�j�=lX�ʳ�g�����jRƎ�+����չ����K�|(g7�M���n��
���(�P��i��j����^5�����"ՅεSC]��:7�W�6�<�ϟYe�}h���I],.]t����m!B��s	�Y��p�Dav�ڼa�l�I���b��oG���gӬ�6�n��Eb�ܩ����b���+�C��9W+#8��וЫ���<�:;ԛ�F�2���ޚc2��g�x��l��$�u|/���V��E�����ޮڋ���dgڨ�[�b���xk�ID%��}�d�O�^�f�u�{k�cQ�|v����ۣ���\d:�n-��5}맙YGjX�hj�]K��MV��OoT�IV��5��س��G!�
n.�\:u��n}"��:� o2.ێ��Zh���k�WB^����Vm�|�-��؟mi�"�C�e�����'v��V�k{[���Hp6�C�۫�U�$ol��2�c�M@/"�2�:�u.$+ǹBj�fIJ�n���W��P�L�����#V).��NƦ�Tɧ)��Q�=�E���j�����p PMf���T�J�u���a�G M���v��F��9��L�Qd�#�:��c2���(�um\%����3�J=��@i�Ǣ��dF��w��_IƇ+{�+2�.[
COw6�R�Fw>��3:�s/(Cɮ��<���˰�{4k���p��W6E]l�����|`Y9u u	u2����(�Ԗ�,�k�/�	�ݽ��f�kv�xK=HY)���-�y��J��G��b�"`i��.�����Գym�uk&.���r %L�Vڍ黼7H*z����o�*�����c0�N��pK��f��-5�q����~��z������੆�}��b�qZ:����ܨsa����<oD[ԕoBw�Ce��́����R�n��E`�P��4�L��/�}��<0���lt�����m�*�xki�`�@��r��.�4<�p3��u/e8��$
��B�b�2=�{p�2�-Z�����na�)ؑNJs[R�tv0��&���us]�Ӧi�e�ko�Ai˫�.��MYqp��|u�e�8��U���M���u�������n��ވ�V��������Nv�&b9�V#t���M�o�&�a(�9[�wh�v&mHePnR����� z� �ݥ��\���}N��ݪ{B�:9ٮ;�,م3o�@m��E#PwT�J�p��5���/��v�]N��+���P���逌AU�+�cqː�$��P��]A��;I+�e�g�o[��29Lܽ�#4(4uvV�\{n���_f^��Xvwb1�;����L��լpe����+X2X�֦��D"�ѻtnY]��rJ:7քr�P�{�b�gZ�:��y���A�:�z��"� ��w�,�4c�v��Wu'�����Y2�'X/6��9���r]^�o���ی�켘K���q@�
��8�B�;�I��4%A�V�fY�Q��x��${S�t}ʚ��x��'�j���[��� ��������G2N����C��R#f�$8�i�t�=��ظ�)B�s٪�vU����SC#�U�H������a=���yv�o����A��[�k �I�Oy��W�tks�
�\�&�
Їu��[[�(�)�"�T��ݝ�V���-0��?Z���.��%���[���a�����Ѓ ��S�D?.W�����[U��],��5f��ҕ��pm��5�}do �;�Jp	�G�g ����s��%i�>;W�'R�d'��L��ʝ��f�*���Ie�u��c���S����T<:��v�����o�3��/��4�b��3t�岺l��.r�E�+��ܜm��J��[��&��Z�-��X�� �(������U�-�֛�#���5n��k�c|2�FI�=�e�p��B������Y�XU+uz�#�J�|)�N�>*�)I�y)3�K�	��Gғ=xu[�e�\�K�N9C�7��5L4#Gh�Jv��:3�U�u`��4�՟o>�2��J�!����#���4�f]�,
�,��XZGj�G�eo.��+��t�=�M/�z�"S�B6J�^�7{pv�wQ{AcV��t:0�S��a�G��_�$�Y
R�Hw1"F��V�-'��*�5F1�	Wk��n��W[t��;݄�{f�w���4蝕)�C6�d�=�5�O.'v�1���1|*�򸨝-wJӫ%�F,��<� Y�EOa�i�u#��ĀJu�S��-��:�Csk�<%>����A�۾����ri�*I��
�����I���Y��B��ԶL����й3�1Շċq:�}C�ɓ�z�Ug�쳥dzs��w��g'ب9����Ҧ���ʊ�!
���u\о�+����h��C4vզ�ZupW���k�5k������V�v���p|R$��Sw�3����ݩ��5
Fq��;凕������&Y�;%1��ٕfg�e�7�#\J�n�a��(J��xS��1�Y,Ĕ��$wtp�����u�U����{�=����E!pe������ţ�t�'�yzܹ۽z&ŋcB����'b|m�U�{Nj8wWt`�N��`y���Xr�fIO�I�p:�J{M��#չ\/�iT�M��`6�\.�撳Q&`�� B�6��a9Z�3�8�qp:cF�*��Z��id�{��SYw�V��
\�����$���N�=Kr���Ro�b�Gm�'�ś2r�3j��.>�.�V)6�GWtfN�L9��rܥwR�O)�dM��e��ѯ�:�(s,Sݽ�M��Q9R�g5)xX*�q�i+�(Qnuncy�
O���Σb.�ѐ0f��6��+��4���hm\��ȷ�wfT��E�"iqS�Zܺ��(D6�=V%K[����y���*J�X�qRЪe��9N�����U�:�n$�,3�*�6d��n�a�o������pI�H`�nv��|�#	�a�n��	!�9������D�HվتӬ���jV½�Θ����j��wJܵNRΛ�E�L[��StJ"�#'+s�$%^���}��"�C+����4����Xv�CB�<�i�:���Vi�o�L��JF��(�f�p��\7�u�\R.^�Q��@����ʜ� �Wf[;;�at�!��Gk4.X%X�2^]˥���f�]VzG��9wp�rLV��"�f�&v������{f5�1�\W��0��*el�ˈ
T�܎SŚ6Z�5
�vư�d��7�Q�H����jH_AQ^��Qg>|������q<irތ���.��5>$��c9�}���t�|�1pxq7�U�
�VpZ��U�A�)��wf���,�絷S��j��<��7R�`���� ���$�s���?[�����1d�,(�w�bzq9c�Q��o�W=�x�h�gm\�z+�v��wĂ{�-�vj#����i��'|C����Mr������-��ʍ�������i2nhM��V��uI�pG�)�o���5�!k��܆�Λ75L���T�m���՗Äe�djܡ�3�J���ȵ��2�S3���*��_^R�{|2��/:wAN>��e�6��eαx���X��\aH���S�_5�6�Ȗ�ˎt��0� h�/��ǩ��%�RV�)�D��F	�mr�)��[Ώ5ӻtԚ�ړ0+��$��5iS�k�9�4��m���`d��<�Q�m��j��q;�yӫU�æ�����̻N>?�J���`��JM�;�ٳ5d+�b��^�S%y��y� S��:���o��Gk�>Њ�<���ش�z���v�m��:ʵ`n�F�s�9-�����~�iT ��W�#V06� 2����p>�1^u;�+�'�eb���ŀm$�pAMU�QĀPi"�L��SK/�JW�˩׻	�d��]��\����� �΁��V�V:W`ǎ)�h���@�	�$U�)�ݝ[��0��n۪�Uݿ�;<�73;���Zo��]=�h�ڑ�,��䶬�1Tע-h�ʽ�Ef�=��K�X<��)�%H0�ƕe��a�bUa�'{�� ]e��l+���o%m��9a;�ޝ��&Ɓ�Fᣑ�]I�˥S�4�
G�Їt���wP��+�:B��f��ٶ��Ց*�ojX�e�ѝ��]��6�؋ 7�A�������c���1&.P�xr&���˵����[碘e�$=ǔ^�6��v@�.+c��f١s&����f.[�i�qsV⌜��O��;1D������b�t���I�Kh화���Y2V��@�>�X'l�G��nT:kE��fKAoX��<+����+�vǷ]��[0�|�$���4t'�t�O�w!KU�Mp�X3-���x?���a5xiŚ]�	��A�Xk2S���i��!�ݒ�t@*���=�9���Y���u��{\2�5e���qXY*s�4���&V�LM\�i�c{J�٭�/r�P���t�z��zK��aG#F�G�bɄ��<�L#Y��Ѯ���Pot�l����j��.t��M����ֺ�����Ȭ;����]0��N=[�K�Nf����Z�u�:���-�E��̔�
޼wl�J2�Zӿ�"��ݝ+��޲��+����aΦ�l�9ʓ�r��yG�mXzi<���9�����������-�g�B��o�MY�Z���Ń;5�#�.n�8�H�V�͸�z^��7��-�"���+
��o���R�4�dF0�ќ��N�I�i��Ӡ(Ջӟ1��F�0{9�5�E �As�SS3�k�60�a˥�1N:��.��ˁ��LI�s�7��E��{)��ؠή��[�v���5K�bεu�'au�(6�m�K�9Y<�������G�ʴU��V�/�i���('p�ܱ��NV��2dq�qG��s�]Ӌ���V�a1�+����+M]My���j�:���ج-���7�(�7{zl���Nu�3�E4��n��u;-GC2�]���v����!�I����á	}&�*�t�QZ�hŷ�����=�e?�Djp5�W`�&v�r���%�F�C)��SV>5�Z�l	�f%�GGSi��[�$�Na��y5&::"Y�iѤ���Z����V�3�t�G*=�ģXM#R�q;v�u����tu�+_[L�wG�6k+{�Y�Z&j��_KZ1D{�mn�Jѳ95Մp�)��Kx^�v��: ��}ˊ�	��<EEӮ{j/mu��| Z{{R=�]��\H��[%$oM�\
�ʽeFV�[����Ŏ�p�ɼ5
ʌ���<�􎼤�w^��w��k���.wT���ȵ�Vneة������Y��}Þ�\s��LF�nI0�Z��շʝC�����~
_T���;��Sw�ūJD�U�-���n��������tܺL��W�x���3��yPRQ�
�V=)v��ɼ�*�K%e��4z�xc����ei$�jˡݛ�+'�]��oD�6��s�r�m5�u�V�͸\�!��z㈍��b)Ƒ��Q�m6o�"8�58���𶃻4��05�&��P�{�F����λx`�/*���9���2�i=�q�Ge�x9�ޑ �ә����A�p]��lv,5�*�"s�kQ�4��Ь}�e4>6�Q�Ű��J=4�MJ�#�HR #{�Aj���\�u�0�|��n�����3ksUwְ.���W�i�IL{&����!�b�d��=��Ν�x���V�������H�Rs}ɂ����`���W��Y�`�����SQa�J��g7�=�#_,"*y%��]J2���*9�F�z�ػY0`���Զ)n�dջ�[!u�~Y�*�Q�L�v�"���7�v�W;�����s��L��9�Z;F�������p�⺨YӯnG�tb�va�2���i	V��vѾ7����!�*"J�S�tM\�9@P"_ed�d��>亡sm]^�XȦL����zW,n°%��X���5��ˢ��Ԃ��u���I�����x��ȨIȒ�֨���I�fU���G��mz���7���D�TMY�W�ҵ��m��Fc�).���CN��$�=y̱K/r�1�E�p6.���Q]�h���ު�)e4�ZQ���H̭�G��׀��n5����ھ���96p_'�M��%B]]c�J2˻�Pe`�j���A��-0���PU4��.w���z��w^(�*.3������1����\��"oo�o'��f��oʆ�sk]����V�d8�ɫ������L�gI&�1St>!�:�į��-T3�w,��g,�yu2����v��ONm�7q�(I���H yЫ�:R�$��/1р�������.���S��<ə�4*��t�m_)�F��j�lY�|�sڳv�-'����,�(ZRUњ�ſE%�@��LC0��I�4A����f^;���v��wQ�x=n�VЈ��������"��N�\+ks��`��^>�h%�,�pf��%`�{�\�e�X��Yc�!kA]ʅ-Om� ��s���u�r'����cx��1�����VeH��5�zӝUb�%	׫Mp㏢� "[��ӯ��ڞ�5.͘\�싦!�y�RZ�2�kX}�����Wv.ü}f�X��zN3ǩ�'�����$ٽ tv�h�.Ķ�͵K�}fDV����W,1\���{�����D\�T��n��e�핺9�7WNV0�M������������{Ke�tV���t�j5�+�j+��<���^ج
:��,|���gj�e@���mZ:�s�����8�Ӊ��!�}����;��u�F�XG:�я9ڼQ�Sx*ڋ�$9O5�Zƚ
X�q�/v]�Q�o���ء�n2�P³��H9��Ҵj��G��ֈ��+\Ku%[�}��S�2ʋb��E:;�QL�f;�kw�YZ����l*wA�(�z^V�/�ăϹ]q�@�	��ʋ���<�X3��t�1,Ѐ�ܹP��d�zfJܽYv�<��@	��(�M>w+��/��z���r,�^��Z��d���=.��[1D8��b��c
0r�:^X{ax�.�xf,,p�E��Ȏ���I�ܯ�����2\��M��x��=Kk�m��|�n��,��0�F�����}ӓ�k�<�c9���`�ېvH{5%u%v��x�/��"�'��og[?vY��QlNb�b�X�C4��e<W��ގ�)f*�����{GǖUMΟ�ʭG[,EE��g
����u��#���7���xێ�#Ȅ�fuNҨ�i�5�H��t7=O�T����g9`�h������բ��'՚��ͷʝD.��K;_i�Ů�3����wA)�xJ]��eL@���@D��$U%���"*����Z�TUb¡Q`�
�ajւ�QE���b�PUF(1h*��-±EQ`�R
T���e�+*�R��b,A��hV-B��UX��b�AdU��2�A�mB�ԣKLLDETH,1(�k`��E����mYU(�-�j�j�UE���Tkd��R�k�V6ʶ��ȱb$��V��6��lV�eb单V,A���m�-@�JP��m�T��(V������R�&%LX�U��1�����P���Q�ъAX�X��*�F\3
�iV�H*���PR
�[-��)X*��ZŘ�qm`\�rգkZ�� �e/�}|d��-�u��(�0n[�<�x-�.�c}���>�����Vi[<UE����^U��Kc�ʺRs�����UȘ�q�Y�/�n�w�"_Rk��V �+MXwYu�}*�	���hWx��p@��.SOǢ���{�1A:e��4Bӎ8娣b��&+ǔZ:|��%�n��V7�u���^༹~A�}B��ԡK5��!Ҫ���0O����	v���'���e%Gn;c3�S>J���O�qeqS�{�uC�}F����GDp����G�Ж������OU�Yb��0�����b�n����9u�dc��٢��٬DԮ�ժ�Vb�+����nH)_�A�[@�=!�DqT.E��N�FB��g��'��䯶������t��3�|a�!Ru�nlD�ⶄ��.����}xd(�(U�-��{|��Frt�.	 ��6�~�V;�O��0<�~����.S]��ey
V�o ��Ϫd$z�<\�VZr[�q�e�A4hm��0�se�t��e%��7��`0�Mhr*���g�	�܌�㘧���|�)�`��Do{�b�������l>� oX�uLo&�Qyp/����M�"�Zb���u
�
f,�fw^el����P�K�� $#;]�q��H�R��s��0�]s7��R��Q����asK�ǣ��;r��:��>T�����&�B\T��O](I!ٺWI� I�Y�����	�V�<'پ�E�w�\�yE6�5�AIbr���֮�+D��lL�E�f@�	RG�D^eq[R�ٟ�u��n��kn���FD^&�HG����>�w���\V�����(;DT#�E��=o�-NRz�+��{�x.��;Q~�3��g��P�B��T��,=���Z:SV��j��|8\8���픻z{V�4=T4Ucٚnzi@g<]B;m�o��tV�Z��V#a���dw�=Ǡ��[ ���>���<W9ԩ�0��
Q�w���	[������nߦ�e���y%����PHU�T��+��XШ7��F��p�%�E�U�x8��:�E8��W��x�F1ˈ��p9����Ixw\hh�4��6*��Gxq�mxmuc�g��ɾ�__�w���/ m}]��Іk�Ǘq���^����P�C�p+[�й�Q���7b6(<T$�4ҋL��;�B u���h��S�@���7뻿a^���-r��e>bg8��YB�)x��u�����}��{4��K3�X��$�};�NjŰ��cBMu�Hq0���o:>�{�����e_=�]ʺ�̘���d\�묱1w]_q����U�����1-�iG�p1��Q����q*�O@��'2oVul�'�et��u�b���u�y��_�۱6+�-FaE6$��$@��^�%�%��J��X=^���d����ق듴Vx�C7��mE�ݻ�u5�:(I�`���=�niS��se-���x"#r�*�mAU�5Ĕ��C^q H����0:��YK�r��]�?:��:s��BL���@�d#]�WQc�4�2A�
�^m򓇳����Imp'�<g,V�����	�G}1�2$���"��Cuݑ;,Ѽ)����$�e��L4Փ���r"z�u�����^�էpT�#{#�Fy\c��tY=�"�����eY�TFd?b�g�3��>MV����� ��-b��xL%yME����oq��9��#׻AtĬ����=�i����߇��C�m��F�m�q�5N�����E/%��OV�� �V
_d��#�R�:/�ky�Nk�3��եQ�R��;�ڷ�n����T��p�S�"��%�J'FO(&�H��Kp��o:�.k:Y$?{`{��2B�Ы�ՖۧL���^6�d��xf����	�KM����c����;�w�7�P�#8~���M��fv�v���ˣϮj�Ƹun�J.5�oq�"+�'f��h�pV��؎�����).啧���j��n� �+���u�i�z�s�����{̊7�.��Z��mX�Z��ꀱ��#p����Q�U<�ap������e���e@�q���%��%��2���P&���8M*�H��t�\��D*��d��$���Z*��O�2�\�E��sS�ٹ,�;^����!��^}0C���>�q�}1�<0J]��뛼�o����8ѭFm��}w�\mz�a�ҕ���#\i��a�rȇ=T�'�e�%z����y4V�� �`�=&7 ��t�(H��Sg�!u>�8�+�2N����s��r���Y;o;W�*�@a�
��Nn!��TH��:��B}u�Tv�!'<a�..���In�JG�sF	�W�J��O��r���5�;_��5Z-�;]t�b��{��:RS봽:Ja��Yn �r�<ќ:\�d�^s�>��v<uMw�0P!K���#=د���;fD�4G0���,v��[��9�&���6�8`��� �z��Pt�k2j�,f�MV�JӾ�ˀ\vn;�����㽳xu:�L�S�)�^�<���U�Ji���p�tN�ә�D4���ܕ׼��Y8�yU�[Xr����;r�\�y�Ըw7�:��u��3���i<ƺ��R c��r�>Xw�hW����2�jw@�~�x���oi�2���վ�W��W�

��*����5ȫ��*��i7'�bwP�=��z�xm��R.��\QS2,�@z��.q�X̔.�e��Y�I��Sz�/TѦP��_:!�*�ן�7�S;�E����|&��������-N�NC�rh�Yݛq}����]�~p����`:�F�.�B�c
�������9�*v�lRy+�v�FE+���Q�3Dg5���%[Q�j�ʃ�	a-ѯi��n�e%m� ������r�u�vL1�h(�b�T�q��6C��oBp�(�NY�
�=`��G��Q!���a�����?	�o��zo���3�B�ki���H΋f6#�����y�<��'��{��4
�U4��SK��M����Vusѷ]���}B}!��Jb�7�n9�i��'.6��������Ip�LGd�7r���B��	��]�"LUŕ�w�[Ң�W_,4Y�R��5>�nH)�,tP�^Q��j��ϵ�n�sO��/|ѻ���Y�S�JȐK8��{)5^]��xWuӮ�3�?�p�^L�g�yq��[�.$+8a�s��5�;wϵ�U�R����b�ӓ�n�W"+pQ=�<ٸŷ���ձ��.��n�dρՋ����{S�1Fm�#�c���t�����������+:��j�F2	
��z��'���53˥�IM%9���vU|Y2)�t5�p�!�P�uy:�q�S�K��3J�g� ���7��Y3���sO��J��sF�"1�s�}���3�C���ѡ��2F\����U%��a�q$�m6�t�s[U�8�ѽ��=�`fK;c]iw�\Q[sr��҇G}�٠�)���n�'�X�=U��Y�"��
�̉.���9^ɫ�oy�����"mϔl�h�B�u�8�K-X%j9B[u�2�Ga���RE��qYC�Pڐ����҉�c���_$���9�;�趫���^�W91����X)���l��3��*�;���a-�U�V��_��G\`n���k��j�{��Q�d\��G#h���8��:�W��p�kv�	�~��F���z�'��pP��m��x�tV�z���Q�0��m��2�N����]qO�;Ṕ]$����|��s�=J�s�[�"�J7�8dN@{=D��g�>�U�e���F���q��ُ/sy��ܚ��*t��Q�L5��$�^�k��������Ʀ�ɭ�ᅚ�yC�7����*����׵���ׄǵ%\Kr�N�U�x_V�K3������ծm���u�v�4]��L���܉��t������
RJVԑ7����i8��n*Z�[��9/2���r�K����8X<t�4�����p':B��g��<hb�F���H�j#�$�me�"2�!9�-��8�7Q������D+��J�85Q��L�5�Z#�Z�wWK�T,����]â�P�n��F��"K8eB�fv!��B� pY ׌o9�eL�m`���h�>X���{r��p��U�F�;���c�Bx:WdZ�$lI-�'� �V2kf�j�}bz�ތ���+�͘.�'h��q���m۱�bq��:(I�C���׈��ckt郜̒�ƑHysN/6`�#\I��tCf �h�ʸ�+\�C�u8҆�t�-�ζ�E���
�I�^��t�x�b�_��+���i��Q��˽[d3��S+V���[t	���,�4x�}��=4p]�8W�U��f��i���+�7x�:��q6C	�%��(��'� V�ȉ���#�C��x2�j��zG�|w۬ԁє�u�YY3�q�r�n�u�/{��S�I��Tj�(^룬���Q*{�)bƣ���O�u͕�;�ZsB�7ԈdRݵ��,=m�7�ҷ5!�Er�#���E��YdLѳ�y=�G������J�����m����7��E��l�lԌ�م��͹�e�j	]�v(��bgʀ�-X:�{r�f	ث���<X�����`l���LJ�:)�8�sN�uf�Z��m9ٍ	>鍹�e����嵛��B`�
�I@�Ϟ�'eb���K�K�ʯ�K��(�^�󎜻���T��*��9�~8p�@싻3;]:�!A/��H�kx���U�5>\��������=�y���k���:�(�[Tu�T �(�诊�\���g�W;Hx9���y�V��r�ޤ��Z��`�JF�[^�{����G���E�\*��i�l��>e���������%4y?9�`�@�oh��°�ЇJ����i��~�Q��^<L�Ak�u�ɥ�V��qȥ��$:��ӗz�)[9��3��`���U����>��)�R�5U1;-�DbYܪ���$�,Ǟ�	���t�h���N�t4מK"kκ�@1j�SW)�zz9����g!�`����I�D@#�}6}��>����s�� ������U��tsL�5v��W9���p��*8M:����7�vX�eV�H���C އ��9�n�E#�c��),�[L]^�����{.�N.up��%���U��'�6�k�������(}���K�.���^Q6�3�����y]��1��\w3!�|�s�[�*��mD�i�>Ҷ����"��D���b�1�GUO9{qosK+.�r3�0�4��~k+Zaw+��5��~SU���R�ӎ�8�؈O!��V�ɡ,'�u��q�r�<ќ;��# �:��C�p.ǃ%���#v��z����-�.��"���뺎�`����Q45�F��g s����Ӱ�����w�N��D����*����n��2���O���T�.o�U�=6���Tػ~�wvx��F�.<»-�¢���E��t*�o�C�9�sE��n��Vp]<��T�b�Z(�<٣V��=��b��sq�1��!��^��>����Og�+��|���{� ���yl?k}zs^����#�@<FB�gb��@���;Z�ݏ�l+�Y���Ii�%�uL�����g�x�_Ӟ�V.|�DW��ԑx���05k[�EW=��a��1�C%��P	S-�	sd;)V�`NZ�2�1����y>�ʅ��b�m��O���.�(ܥ����[�u�}�q���#��Wd^#$��H��0q1e�zg��p$�H�wvxkKS7��=yY�q`�S����gk�Jnk n��0m��PauJl8�Vv.��q�X#���w�֯��s��^��sx�6�5��u;���i�*d�k�[�A����u(R�`�!Ҡ�#:,�тOU�rd)G*w{���z�@���X>�T�qc�3�s>�yŝAN�ມ�}�P�|��;�sk��{�oD��QJ�H^#	5R�������ݹ�=��5͜��ͧ�g!I=[�pq��6gjY�'>�� �~����l��VP����7]0��u�����Sl��C���T3��Æ�n�ѿ:�p�A!W��Csb �dM�g�K;5�����q����H��`[�u�je�C�8��,��uX� S�K��3J�3�:��䏻`u�Y�;����s�vi��oL#�hI��N!�y̰i4hm��0��j�h=�NC���<��N��ۙj�D�
7r}bzVE�J;z�KJUE[>s� Ҋbh�9�2f�n.�z����.���)�I}�E>/c2,T+>�<-�p𙾓E�o����!�.E]9�
��{�Q���M&�؛�[	t��t٦�W��]	�V�|]cU�U}y2�NYZ�� �+�,�kNn�N�Ƕ��ۭ�
��+�{z�������LpQ"��%�I�٥n`k!C��3�"�ZC�`��}���n-��$wTb	���8jXTs�ٻdc6���1Z;������,;yj�sA�
����j��Ns�WS6�з��N�*�zҴ6��5�ۅ-]/�v��Ј��o���ʼ�ׇZ�� ���t���*6�ub���Į�׽�a)Q���ݼ�;7N�?��n�u �:^���i;�jf��-��!�|�7����Jֱ�;�q���5��o*����'J��ri8K2_
�}{�	nV�PqYK�	_ǪA)gm�@w�pݝ�������[j�sά�d����{D;�ͮU0������.��;t\=BIF�L��n�Q�3���C٧i
�)�<��殑�n:儻�ӗ�Y*u��E���D���˱Ա�[=r�3O�zU'�{z�3����6,���x�W9ޮ����맂w`�:�G.K`v���8������b��(��&@�s�n��|GW�T��iT���\X�|:>s=T�uc�ghu�O��z�o]u=}�x�mbrI67A�1���	�i�(/OY�6��t+�Q �閠;WL��=B���j�]�1d��v�VL��]>�꼍�x� �u(����be':�SA;Gr�Wt.�z)��A)��{xDCn�u�=� ��5Q�w��s��Gd�K��G�u�kdN�w@y��]-�8� q��j���8D}]a�<iU�v�_=Ы�gQkK�J���m�{E�U���.�ݏ�U���o�,lU�����֮�)G��wGf�"�٠9E�ɼxI��1�%0�|fԨu兓�k�f\{I�k���t�a�L���v��w��Zf�8��:�VX޲��b�c��ۙL%FW!����n�peAe�S6��B�w��"�o5�]rI޺�\�ʶ�����=r���޹Z��]��,�ȝ�C7��pI+�3��f���ݔ���VV���ǛS��#|6V��s%f<컰0�[�M+��GMgv�u�˹W!*�a�*l������M}]�����Newu�y]XwH;�Y#YƜ��:�6�Ь|�.��s�"��N�a��⼡bj<B��:v� �l�J��*%ݮ��:��ВW;.���ɖ���jX���
��1�`�yHQ����	�i��/=L�����Y1�d1&T%������c�t�\K����Y�)q�]��Ϻ�ekjd�xv��/gLA"-.�e��t3]��t��oo:๡`���n�x�i\E1w��Ԗ*���)�ST��Xt��xc����bĈ#"r�We�;�{����k
G7�����=G��]'<�N!�]��Ue���W�3���Z�=[�JxW�ŊnO�ޛ%-�0ʊSʨ�ZV0����~��F���|,mٙcj�
��"�P���*�4[�p(ZADU��m�����­�mb���Zũ��#T�)[VՅEj�m��PF�*��U��TU-���T�Җ�j�,T�X��h�T,�Im��ł��������J�iZR�mF�X��
��j���J�D**U�Z-kK
���h�mZ�-B�j�"J��A��ŵ���*�Qe`��!P��b��YRTb�)U���6؋i��*ڔ�TQؖ�-�ڐm(��m��EҢԭ�Q��ȋ"�H�ڥ�+h�E��j��(���(ֲ�-�QVڪ�j�Q�EE��RŖZ���Z�V[e���XT�E-Z-k�F"��[b2��J(������V(��6�UYZ*D�(��Hh��{k���]�t;��P����E��|�}��Ver.�$���n�v�#*�+�����r�z��W���{�Qc���~H����Q+����[U�	������m9�
+���9N��O ��=���3/GDg�+�MH��48��u�7T���,ۋ;����0GM��}o�J�c�H�=�;��K�'R��dp2^���w�#�TW��Goͻlc��[�S�
\Y��!u��y�i�^�(Q�0��$�����`�q\�L�m�56C �ѯ��\�g&�f�[ka"&���\�P="��fHf�e�_�)%+ڒ,�e�4�Vy�n���^�Wu�v���[�o��e:���H�@7."(#��Π�TMp$�;�44:�TŚ����s2���Jk8�čᬐ�S�>�(��m���B��H��z/�Ex)E��PȪ��{�P�'V��a���r���)n;�5b6(<T$��T&c"�D�z �+(L1��E�v�q�1�������q)�b�"����H{��v,c�JR��AR�� �u^� =�L�ɳ�,I�w}UĆ̀NloF��+6`���!��mCt�k��p̸���(s$�E��q�NP"��fǭ<����"��K͝���p[\�;I+����Q����[������d������LD��8 �+`�V1�{u�C��GǓΤ����R����7y݁�ceMgm�F� "t����C3^!}bL=1������9�@�~���sƯ.�Lq}�R�E�ͨ*��5Ě	:�Ȫ�W���)�B�;����~����>��;�F���b(V�����A���QdvP�G��ԘI��l]��MA�i%��%�L�N�>����k��*lu��H�2��^uq�Y]=�f�R�UC��'/yC�9Z{vB�$�R�$ĆՓZ��[�x9��p��5�/�NГw��Nn�2�5�����$�X�݌����:alXΖ�9fz�gɪ�"ƺ.hC�N���j�"�*;;�o�Ջ9�-�Z��G�+���b�E8��i���՛-F�	5�<���qk͚ĵ�ܺ͘L�~3�:6kb\8��6Q3�4�2�H�OU.s���1A�S}#���г����l���YgTȻ�fvX�TEJ�_X�D����)�lc;*��p����ܻ�-F�N��9GJ7�����ADWED㮌�i�3�)}y/��%:F�ws�ھ�ф�'�Es���]~F�Z�N<5�<�uAp�T&���+t�<��P��κ۵w�#q�,��joL�sa��|�]TlmZ��nZ�H�\�}�+V#3'
.��`��`����]�:Ox�<�ۛ� *[�E�-���]�fZ2��c�s�U�t ͶF�x�su�L�ܹ�;�`�"��ֺ=���ٽ}��6��f��s�\h<�.'c8/�B�7�!�Ұ��];�b�� v�K�Bz!8�.]�W�[zr�i���1�ѣ�%+g0s��tc�$;�I�S�LtAQ��\�*�	>s�6M��x���4y(��Q��u��JV�$�9�n����dM��{�Zh8!E7��%��tu�����+ ���D;"��C�}qNW8s��/+ie���:���<u������P,)�R����׌��}��zV�;B�����y���gFm.��tF�N���qZ]��y:�Ȱ�s�Mi�܀Cr�k�s�E� ��+�ft-f�Hv�
!�0�T�n��',�^�i�1�μ�k�����Ǻ�Z#�H[�!�+��<�O�v�Y̋#��뻨��(Q~p"G5D־��6!�0BX�a����#��F6�f�Z1>b�F�9��(��VEoH{�X�Q�)D�r�5�\'�u�!FE>>�T�o'����#��u;�ȩ���G�][����+�ubn���'+m�v��|cCeяU]��;e���I1q��EF%ӥ�^9��Vu$�2I���"�|E��f���`��Ou*�/�W���w|$[u�u_F�s�����y}��{�V����k��\��J+/���|�G�5z����[��%1�Kv���y�m_,��Zr�{��J�x��a�yC��B��sq�1��"�3r�+ F�z�ree�9�I�W�}���>���ק5�](�Fh.x�$�Da���B�ޱ+.ļ�8�gWBE�g�W(�J�e��Ɩ߭t�F+U�TX�8r��BB�zC�.n9�E�2,QC"�+9P42Q�%L��|
U���n��&#obu�n�9���V$���L�fgN�L���� �="�ػ:�)f�4�d&���H΅*yV��!�]{ȮZ�B&Ͼ���$?��3O�iw��}>o�G�Y�j
����Nl����+�z^���!��Ȱ��GE�
V"B� �4�pA
�7r������r)T$r\�6+cR�8��lѳ;R��>�-�+ �����	�j3����7���t���}$a��o\`�;��8p�n�ѷ]v�7��:�6� j��Fe�od��
TJ��7��k[�W6��$i�0����臁����䧎}�f��ʙ*��ܼ��I;�ق���+]]�����!t��w�b�:	o'��,l\���fnM}�L��j��H�}��:��J�:�&�.����x����WC�)��f�:��v��՚1�Q��M��Y�C].��	o,֨=3�ܥK��X��9���1�=s%��p�8Cz`���kzS�q�e�A4hm��0�B1�ss�C�B�^,���q���4O�!�r�ּ�fU��<�zw>��[>s�僮0�3-�]�*ދ��q��� �;�/�Ȣ$��Ⱥ������Zp��4h0%뮼�W�
�*'�IF͒%�:�	��G(N�u��O��+X7f�.U�2�t&�V����T�_F=��o+(Ic��݆ܓ�=����s�;�s��ߎ�,�EX���+�zCa��h����_�-�W�4�8nea�5ns*E�s�v
�|�[��ENq���C����ѧ�X�O���.�PT;�?L�t�>5်�v�۱�-��U���'�xNI��;v�w25����0WG�є�Z���7����ț�M��-��O�Qk�j�嫖��\7�ȝ��L@P+�\2�^� ;�WP�����Q'�CTں�y[W؊݉wPYS�+j���:t�5���@P8�gPWQ!fYK.��t��vq�
w�Ku	���QN!vS��8�黫9��\Q�J��w�h�ϲtr�|}A�x���!��7K�b�;��uй-[�s�7�����<	 ��K��B2���4�2;�4�?�Nپ��M���8�]�

Zz���륖��R�g��ݳ�.�(؇�l��=�=]҆T��2��gp~	n��♳1I�{; Y`UN_P����j�l<R$�4�3�c�I
��:¸�]F�T�U���f�w�1۳$�}=�p�R��
�!�pnwb�;v&åvB6I�sx�w-�(f���s+p��s�2H�F�	��d��^L�����C6ͨ�ݻ+.�d�L:�N�5|���aΊh8�+2NɄD#�吋�f�^��JNz!����D9U��|"{��d�4����1Vۨ�SSY�:hB�k�	�_��YC)��sr��ެ|27[�*8��%��C�};�(O��<ԥ���@��ve3½--=��M���	w]�v�
�`��T��;U���Q&'ͫ&��9��@��7�L�xY��41�*u���6��R,�8WE�H]0�/:X!��T�؆��	��"ƺ.i�t��ވ����ךd���@J�Q�R�Dm��"��W�4�tS�q�\Ӂ`cue\V�!�vX�:5�r$IFGSv�fqh�E��%#�Ë@d��WWG���B�^a솺J��G�؉�6�Js{g-�6f���yj�V)���̳�!���md����A�T�ޓ+��h�'���)�[�
�A�Ʋ�!/5��/)���q{���ޝ;�|+/�� ��#Hqg#iK��e9#H��/T���\�I��o�7��u-�'m���<g`#d-;"�����ꈡ*I}���d�N��fy�����p@b\�	�ѽ�8x߱.�=��A
"�*'h+���~��4-��&�1���L�>Ί�%��&�5PD%!.���n��B=0�[�f(D	7��Q���톰�����[�����`���Wʡ@�hC�Ҡ���z�p�I�́g��@������q �!��{"�*er�z�)[9�C;�� ��X����^�i�����^ts�n6 ��	Z�O>0��8�}�f�He� �;j����/�Q��+�\*�K��JՑ.]W@KDʏ��7� j��0�F�ڃ�U�~ӣ*�c�t��m�c��{��c���[�Ω�k��*-����D�i�``�;�廀�A�
{�uO��VF�m�xⴻh��I�E���J֘]��ck�x9F��Fz�Pmӥ�O����)c�4%5��++OB!���YO^l&�J�0�ȷ��zi�@3�3���f8+ �Su>N��x�9t9ol�S�̥������v�@;]����Oʼe�CQ��[{�M+Z��N���zᡙC����Q�}3�5�(�T�"��߻v���A��k�5��\�d�^s]5�qι��J�z���X������ӳ	F�0�㪨��(Qa�`�jI�}Q�a�'*Ѷ�owJ�듆k.��;^�S�r���Ҏ��{�<��?V�A^��/�2n�;��n2W�W^5��-������g2 ��Fʛ1�(��ҊUT0�:�Z�B]�P�mT��[0&�_��.o��Å��r�Έ���#�v8�7Ĉ8	�moL�5�\�a�w�P��L�l0%U{^7~}�Xom�܎;�\�lDq�^1��6��\Cu����W����ddq&w�s��T�%đ{�g�����L�*,ߗw;n��NX�����4��*3�ʁ�D3䩖�%͐��z19j(�,лj�����Y��� i�2�ᾦ�����PQ7Ξ�P������V�Ha�T�H��q�v��Ю�LlGE��qhDq2	�xJiw��|��g���k��@���Q���ĉ����2� ���su~4�GØ��Q�:��s��cLN��ڇ�^>>�jS'��˻�����RQ�~g��[s��j�^D�e�'je�:*�\P�ݚ
.��A\a��`=�V���JVU��ò#v�f�j�?xxz��B����F��8�(��"ޝ��RAJ�HBA����(��⍊� �	�.&�[=נ��o�oNp
�dc�x��<�J6�C�pAK�D���Hfy��ӝ��[�z.�\x;L*F��W�!N�3��Æ�ݻ�n��1�HT�Csq��ȷ���f�xzlZ�y,�[qZ�!Pޠ�C膜P�Qh'U�d�����u��/Zkt�{9�>RΙ������S��;2D�ҜC�s,��״�m��l�^�43��iƜϤ���.�ê�,�"L{anO�T����ζ_�ߍwo�~�{�*��>S%۬/V���X��W�W ߂� ���4=��T�!�7fS=g�a�vS<(Ϋ�ꠠsk;��\n/l���Dз^QA����؛�[*�`Y@�d
T��`�q�&fMfY�76��0��#y~�{tJ�~�>����YzqT��}��ú����{�������ĳ�"�1��>�`[A_T�F��u�7T��>�f�]Ԍ�:gc��f��nx�{��rCh?��+�.��e��;�n'��^��1�H��l��u�	�Vj@��PxE�H��_���t�x���CtߤO��X��'�9�Ζx���H���ӕ�N�(��	R�mJ��4����l�8V�CQ�]u*�wBڑ�?  �ok������j��ճ������;X�3�����.��݌;�G#�����xz�p����LX��SP+Jk��R�GP>s|��s�=�J�s�xa�[g[���s�;y�v_*!��k�nY�>\�c�M��������ƅ*�w��7�3��3�t.�����~�����_W�*��H�^n\D��Π�THF�e�������Z�p��嚌z��0�!֪n"<�=�G	Gۓ���i=-}]��П��^��qi�T�I�qY��홸|ʳZ#kC]���f��whj�lS�BMyƚQi�؇x�B5��$ڲ�wU-���O�:�����N8�4)U�F�9�݋�;v&�} ����ҍwz\�/_�����p a���@w�@Q�4��8#��]KDo��R.G���څ��c\C���U�(Իo�)�΀Ý$הI����:
"x�˚pt3j
��5ėB����r��w(��Vm�r0	�C/����y<��5�0:=��#�e�!`��C����ι�oB��h\�.݂�:8���v�w��ZNĔW|�,��E����X�bt���ln�x�yW�$c���~�Lﰖ�`����f'��S��ꋱ�}���^qђ�[���}" ��E��By��`�\j��Z�;���=��O��O�PKs�P�Ȅ�˻��}�u&wO�;��
����ԏw�I�w��Ԍ���=@�+Vڬ�+�hঢ���U��*r�
4����9��ue�l��|IZ���k�����a����*��_L�P&��X�J��=N�-ɪv;4#�J�됏�b��YU�lO��e��.�{�����=WJ�Jܛx[�63����;�0](x��BE��r}$k}J�B���H�����C~H)ρq��K4r���f�8e�d�ĕ�\{/����Ӗ��诹�c���ޔH���8�1��E�ሁ��v�;�-G�g��@��I�hv�Y�]��X&��{_.u�T�8��Ҝ��<�.0��'ԙ�����@��AL�&i o*�f���۳\�iU����~��{&IO�֗��:��
��.*��1�s���f�� {{ݸ��{�@mt��ҙM��ޫS�o`y˸�uc�/�
Zv|���:t�J%��{�9���ʺ˺�mQY�7����o�	JͰ7�����X
j�*�=	�����4�2^�s�{��x����l��[��D�)��0��;�NB�W,���%�w���5N����Ȇ�tyݫ�~
���[*�v9=�{Fw.
��qޞ�b�	I��J��wkx���?���p��7��O�,��u���9ݡ35�/+��i�SW���mI�Lt�|7�_i�]������SUb���[w�=�֨�u�kMv�5���FjN�;|�8��'���z�����꽸�%d���-�x9p��%���d"����s�U���Xw9�At@�
)r���[х�x)���<H�xn:�;+����[��pB�
\9����1��K	��+6�ި�;]������I��%�8:]���V�S7����'3+������u���7+�[wg;��VL�`ċ}SW3������ʙ!{������whkqv��l����Y<&�a#�&7]N��t���N�S��wc;��;����ɂ:jwP-�7�r�k:k�|���9f!n�ȂIo���9w�](J�Hi��\O��g=�.[m��̧�R�ƻ\��0ʝ�,���ʸb4�M�ݗG�u+1��=�%��V�%A{��aގ{�C{�vmok�*�t�S�oQ{R���f���K�`_tW���ML����y��CS�{|Ҏ�s���p
�W���ަ�Ƕ)�h��I���ꕔ��۷���3���]>*�n*�V^KK�L�&�-s8�9����|����o�4V#t�I�E��Wtc�nݔ�[5j��TUPkkRQ�-���h1�YF
�"��X�Eh�AKB�mDJ����h�`�V��*)X�j����(��U�"Q�T���-
���Y��YmKjZ�+j2����
,e�"��ڐ�B���Z�-�V �b��E�b�UX������Ƞ��j��-EkV�-ZVR�*�UUEZZ,e1�`�TkV"[m��ieaiV,b���%b�b**���+�҈�Ҥ��j�D"��ŋl�QV,F4�Qdb��R��#mR�+%���A�X��*�1F��T�*+(ĭ���+Pb��Z��"*��#m���""��
��1TE�V��҈�*�([EUb��ڶ6����TmEAUR5�Ŋ�-("�j֒	 �I ��3$�`EZ(f���/q㋡�gem��εQ����w\���/.wT�e$ە����2VR�����+꯾+t�;I��X���'�u�\D�tɮt	�|r��u�j.Pu�z uH�2׷׽Vo��~���ؘ�mT��CX�6AR�<���bCjɭr@�s��l�nk��E�k�S}ٌ���kչF�^����
���:X!��:�f�5�MVr�.P�)���/1��|�F��-Y����T���<�����0tS�q�\Ӂn'A8�͚�ڵ�]�RTX�xi	^��rP��7Gv%¸��Ѳ���4��ٗ�Cކ���yZ��G��M�D,����,����Î4�@�dp�B# j�:�(	RK��R%�\c�����j�����l�%��.�b\�����F��lco�Έ�8S���])��=Y���]c�����2�U���Z����r�"��[^�-�(��	[�f(^u�`��n�T�v��ĩ<m��?V�./���eĨ�̚�0�Jmq^m+j����:c��Y[+��U�\���:x�E?L�2`27"b;���=	S7��3���Hw�b��	�t�ӃC��g�ٳ�ۂ75ۃ�̬r��ݑ��ĭ���yߌ���G9�ک����4!>	=�}b�h�!�u4�����8�ro9�\�NՏ�ď:��@º��R��¦Q/�=ؔ�ښh̎���e����G+��Iu��?{���K�[/�[�Kc�: �xd��Eh
��"���t>�8�V-٣F�v�u3�HEȅ�6)��zxia�DM]v�b|*\^9 �F	�A'a� vT��S8F�1 ��O7l��}ær4��)8{胧)��|�-��8*T[���AP⨜/���I��v7����Zk2�VD��E�q��+K�2E��n�+��k5�r=|9v���=xn��{c�a���n���*�n�Th<S�4�I��".s�9�Ov�١ن5�/w����ҽ�6�<v���쵔�iu�߉�~�:���8#��N�i���{���Ĕ-]9Р�6`����;^�w#z��	Z�t�k�^b�G��h�'^��
:#+�F[��{k'bT"5c��4ǡ����gڷ�ؖ�u�K��.U�F�$�ؑE(T�sE͌oU�ѭ��B׋�h��
�]V�L��P/ʮ����Kg۹}���o!�Q�UW��w�ѭ͞�<ۣ��D`q�Y�!/ ���c#^��)��Y�R�P�Y��z��܄�][���r�5�bJXB���������J�mX���=V(eՠՈ��QH�c'LM�&�RT�D;�.��uu�u��ڊݣG\�����f�{ՏsJhu��ڌ4I��]s)\l�)�V>�x}9�W�i�TX:�mK$��u�2z�pC�#,4�=c����L��s���=j���R�O]��aL̲ �q�0{��)�r�w%�%,�
\�%9�~YX#��N�<�����4!�+\/��*���5۪|�T(^�GJ5��"��n�Ƿ+ŉ�n��[����ٍ�6��8��f����})���\A�Vwn<���$pMY��C�}B{!����GE��R���Ip�h��(�6b�q�������l��������ui�hߌ�J6s�q^�$�$��A5{�uYxOK���,s��X�wo�B�u��0S��p0���u�l�BN}���b���S�[�������t�Y����)aW?�]{LS/��q#T_��#x'U��&�P�n�qwb�*5\�&����s��.c���³\����������
�2�M�f�}:�l�\w��ei��L��v�̭m��(R;-}.^�.��u��T�(�H��D��C�i���dʜ�� oQ��6�t3�3��c�˪1Iz�`�A=����8S������������c�-mn,6lt�"�KC�3��U�t�eK�.�c��Nf-�LۯE��}ֆul��|�K�S�d��J�����{������'> xxL]s�I��'�1�jX4ڊ\՜4%r�Do�CہS{�l��	XxZ�f�_��uf+A��lQi���&��F����:9��ʿ��1��*C���w5�t�F:ۺs\��O�n��{�2����_f�t}�HO��������8=��Έ��V�����F��!��И]��<��uMl�g\g��e>�G��9�!�AʾR�%��r�4ʃ�`�e�u9Q�*@}22[6]j���P��ګck_p��)p��Ծ���nvaY��0V�5�tO� +]���oJ���;�Ă	���r.뢷׾�i��.�R����^��|��r�����)}JIKf��-��e���Qϸ�Ly�ѤfԄ����+
U�:t�4ܲK�ʶ��޺�ʮ��q?-,e��W7{�[���_�0���ک[��BGnm���W��$p.:�y��sX��w�_�;F>�똠�W[���BWP�czS���V#b��P�AƚFWx,'ԫ�&�{�(h�4�smq�O��E����)qyVۂ*�%N�h��mP�:z'}]D]:��Z��\�#K�r�Xj_���\��W�Z�f�=���x��]]xnu.��vz�J���u��o�CT_D��TZ�-V�+5KE$�셃��� =n��7�7�$O�G�e^1�M�PO.��9�()U�F�9�݋�ؑҶ K�֛�o�.�Syh��	1�A1$�fIB�"5F�#�*�`�4��Ď!��*�o^i]O���v���nݎs�9�BM`�fI�0�� �˚.�ͨ*�gIh(uz�g7�8FD��8��$	ѡ��ָ�)�o4Ѯ�����H4{��#;*@�&+9ɾLv�,ea���\D�n�<����,�Z�nTن��2^x�pf�>�c(V ��j�9���>!W�]�fnպ�Ⱦ�D��Q&4y�dֹ�B���u [M���v:ʆ!�0�t���,���쫠�GL=�����T�ߡ�'����UZ�F4��c���j�Z��|�V�~;mp����[�
������N9��[�~r�²_=쪝��N��j3`IN2c�FmPX+�P<+�����Y���_����W(jWˣrU�~�T�K"��5����;Q��V���s$d�%��}�:i�6�7��}������/oRX���Op���ٚqH$�Դ`���`	5ܵr��g/P�X���G�b��_㍇n|V�j���x������ye�.�emBکȻ������&v��*T����Ae	��jNvL� e�{�{�ʫX'Sy��pN¸'�R9@�R�<uVr�s��%�G��"@(��1����kn���0]�:��GVL�5��D�r�"����;���u���^!�%�ՠ�'qd��u^��R�я�Ѽ;����3F��B�+dC���&Z�#Q�n㠙��.��ˑ3�5�,�GT�>08��)*g��z��T�l�s��t`}0G@��ޠ�)~6�[:���ͭ�۰x�E ��)X��d��4c�⏹F��Ě����[�+~Tn9e���S��FmF��#%�5�]v�g��R�C�'�YףeR vM����y7��IJnļ�I>��u���s��NPݳ�g
pT����Cy�qUD�!�p[� �1�W�kynD�BںȀ�;aI:�V�bD4��
gOLI������U�Īé����<�UƯ�#�eHdg��
�۷ux�h',�@sF��s�m��"8�ɋ��y���P�w�/�kѰ��ˏ]��W�W���o��1�U��À��z�M^�]�r5*8Xfimew�v6�@�WAw�9n���s��н@ʝ�a'������wd���d�����uzX���S�^��z���u��v&��o>N ��p�:�k��q������2�,f�P���t�=����w2�����~��ﾪeW4��|�;I���7�G#��}�k��s�r��Δv��Y�G�U�K�Z`k�)�Q�3*sn&��o�U�%g��~�4v����>x�oR-���,�"{[�ι��X�Y�h��T0ߒ���k�.lcx0��&�mOm{~�B�HW:ӺǚhV3պ�-}�g�S�Wd6:����vg�ҽ���n�㼪9�8�F�s�a����T���#r(n�'���b4ʊ��{�m�"L��\��,�E��g����{��w����CͤR���6w]�Ps�B"]B�+"�W��C%�RT�q��6Cpjr�N�q���z^=P�f�b����ڽŉ���@���-���%w�1"�Iǎ��,������}�x�_<?}�x���:����~��Z�H��K��]_x �>����>O8���Z�?0�1��=�8��1�ϐ��h��!��Z z��O����L@�_7���y��7f��
E��4�H)|��]0>���>��l�7���xA��z�dS�Y?2���l�I��:_>�c����~�0Yԩ��V��c>LC��0�k"�'2�$��n ���*k,:�3��cKc�A$��q���<���=�(� ��ěB�g5׌���R,�/�ɉ�O\g����m��l��h�������I���g���$FLz��g���+#l�x�P>q}w�u�h��"��ӽJ���W�F-�Ѹ��z�I�Og|Y坤�98�杹K"}�(�_�t@�NX�#�N#�\B���A�w�]�h��P[k�>f`z��2����o|IH�)�Ε���·2�:73s/y9K��]���KqJ�T/l~�� �W�Ñy��k����a���dު���Vu=a�TRm*Az�o�����c�s!��|��������+?2]���βx�����Ry������$�>�Y������~���wGܒ�<=AH�$����X��^3V���i��P��O�Hu��k���T�yO�T�Ag��M�gX|���5�OX|�3�?���Èbv�
�@�+y�e����]�y����rٷ��3�ޒ s�(�z����	�1"��M �Y�5i�״�f�oT���Y?2�N��I�u�=O��=�ܞ�`�IX�h�����'�$<~���m���>��{���E*�;������ú֥A�IP*}�d�2���b}�M&�i
�*r[&���x����
G����u�����HJ�|8�����A��)����#���������~����t��1��>�M$FN�LCs��i�dm�gy�bm ���y�I��bAk�5�~j
b���OhJΧȳI��z��1�$��ǽ%�i����Ƭ�tV��.�7�ycj�&{>�dDA��
��1�^�N2ow�g�>��6����<��R)Ę�;�k�Aed���y�/�� �g�w	���M!�6������-�?!�1 ���{�b�I�GD݌���[��>����������c1�����Ax��3~��E�Y��)�O���zs�?��*J��d��M��"���m"�w쇉�R�g�wh3,���{��~�썗�H��-�����z�����<x��;�C�Lz��f��|É�1��T��J����z���<>�f�yIP<�kF2u���ɟ��@m6��W�ߵ�)6�I�Ͼo���p�3��b�}����x��Y� }� z�4���>d�%|g���i��Rs�x2m1��wH)��ɉ��gCE����Ě�xu�'�����Z�AN�S����~�*駑Z��Vޡ�8����z���Vx��;�x�O�P<��4�$�l=C?y���4�'��H�x��3r��Y�& sɼ4βo/�
���J�U���b
E:��)��Ă>"�Ž;����L�?��C�xn�ܛ{�cqK׺pQ�����N��wIN�	CQYWե�݅͠�W����L�Z*�M�����̠S#�*�Ne�+ʜ9�9X�װJz^n�˵���c���)^r�P6U8�O���Y�m$^MӺ�lL4��V.��e�1�{�	����P�%��y�
#������8�M!����m���,��!���:�b�0�15�<a�1����4�_|�Zi4�"�Ļ5��'_�1�nÉ�*H-Ǆ|�W�5EC?^|�VkΟ��=�
��}�=�`b
E��|¦�HVi�R(Ne�9�M>�*O����O��?�+Z�g�Xo��i�a����Ă�ȥ�3�|����B���2���3�:�R��"�IXt5f�L�2��Xm4��R|�}�����B�Ϭ���O ����i�6g>�3�J�ĭ��'���C���CO̘��'���AH��޿^,%����H��=�?9����]|,�#i�e��i�?8��P�Of��Hq:��x�H%f湇�6�O���솞3�1����Si�~I�|�&�(JΝ�u%��>����J8#�M�S|�O�G�}����si*+%W�d"�&KC��i��1����L7q�
�É�i?'Rc�����f���?g2i��X��=L��h����6l��C茩ϧ��˫��� �a��ĩ���aS2c��$SHT��l�I*2�^~�1����Xq3�B����|��I埙�'�yN�G�>'p���l���s9$�N0,6�>J�;�L�é�9���m ��|wzѴ=N���u�R,��+79�%d�Vs�(bJ���-1�VE&!]�_�̞:Caّ�@�#�N���"T]A������/}�f2T�X��z��Ss���~d�Ǭ�w0�AH�����M�~d��u����Ă���I��N�0��i��AN'�� i*�m�OXi�J�s�߰u��k\������~��~|g�1�� �g�6~��YR(%w��|ɿ,�&!��Ĭ�&e�N��$�+'��-`T�~�J�� ����������3�0��d�25x��4��s���W\0~I_����ϙP������q
Ŝa�t�Ax��1�i�x�$��}��<O�Ry��q6°��i<5ܨJ�I\��y�$�T6�Z"�� ��ߎ��]�n�(�8~�u}�08�)|�r�S
��'v�oy�+�:^�˗�c�(���$f)ۜ��U�Zv.���x��b�n��FE�;mӴ[���mk$�� ������(;Y\9Mޜ�:�����;�������/mK�JCW���Џ�Wh9Nv�!����C.�=���j����s]s����13V�l��P=Ne?e�����ǌ��OP�䞛�H,<k�����1�0�c6~���m �B�f&!��� y�1�E������E�{��>�%������َ��>YK�zP*T���|JȤ�w�ͤ�����H�T��~-��L��Y6j�4�d�c��wI8�2bc�� �FN��I�C���kvN>�'����a}_e�]71I.K�� Q�=� �s�&:@�)��{���P�g���"�I_g;�4��$��xK�>Ci�~OCO��;5t�.���I8�βf_����I�*S�D�q�Xz��e����j�L���}l��PRw�֏q��AL��&�2{�i�m��^0�?s�x��+��z{���*C��yy�V~B�g�OSI��i�i����ɼ���dYG�+b�F�K{'����bw�~�}��+
�~gyCh�B��~�{�T*o�a���lA�5�L��v���ɶx�P?'s�$���S��08ϟm
���9��k���T�Ͱ�0����[�gמo���u������ ��wa��?'PĞn�?$YPyCg�iIY:��yO�d�J���4�VE&z�i��O���"�ĩ�s����|��\ϙQ���,�z2��ϤR���/��֕����G�zH�*p� Df����Ăϓ{��Y8����c�8�����,t����q:�@�T�<�&ى��M>�6�\gRc����� �g�ߙ��y���ޕ|�t&�ymo��Y��}���>�,�'Mw*�3/��i'�T�P����,ݱN���I{ɦM?2}�i���c��!�W������O�M ���z����k�����v3mƊij��4�H|O�?�È� �a�����3�c��٧|�&%H��쒦�V8��e&�>J�b���Vyn �_�`b(�Y�&{a�g���;��{�~��{�������{��~Mr��+��	��q'�W��s�&�Xz���ju*Af�l�����Ă��i'P�<�&5"ʃ�v��
����n3����R�̡�x��A	?k|����sp0��o�#J�Ȗ(+��]r˃��������z��:�y��7�5���;inN�Q�P�W�Xvr�����B�uE��=xv���ާ��u3�+�
�e!B`<��l�*Fq���/� ��w~;�!E4Y����_I�k��6�i5aS`.PCVӝ�/;k4�B[�;^h�b��*�I	,�Eg/7%���g��}������u��Yʇ+�b�L�9��G�C{�o%�6=꼾&�u�4e�c犖I���˭��L�/��ӗ\���L�7]�WgVE�y�AkQ�[����}es��%o3-�����,ΥfƱ��Ҡ��KOj��3}��{�˺�.��d�gJ:�|A�|x��F�Jv��5��j]Z���Z�ε��*����+�;l�ގ`#j����갔�PR��;-a&3f�J���u.�`�}t��0��T�Ֆ�w�(`�ϒ}��Aޛ��m7h��J�8k�6rl}'C����ۇ�N��D X%�ȔU�T��J�P�w�����C�mV�Ψe�h�V��P�nm�2�sǍ����`��]|/e���V5k��NW����l��T�U�E�ly���YB�'��}�X�g@ L�����&IO����;l����s�n���feً��yN�<R`�����?H�ĵ^�@��[K8;�u�"��Y\ ���-��%���6RCs�F<B��{Tl��}}Y�s�JB�ď�����M7f��!����jC�f�-h}Y�r�=&qn�[ٝ}d��}k36�m����_[:b�رs;v^��O7�I�2�<�oi2���3�w̙��}Yuͮ���c�ӗ"�s�WW�
�ist_&{�ͺo�� ;����'Ԍ���ۈkJ=.� e�����*v���^oT�l]�H�?��}佻d������@��U�L�$����|��]K��)�G�R�<�s~a\%��̻'[{�`��p�[��Y��m���m;��eՉ*`��+_^��߆����k8$��Q��%�g$�f_���φ��/�!���5���0icz@�Tں����nfA�<(R��蛀mD��)P����^�ˎ�ىh_k�L(y�0�O����.�����s���Y�������;6�F��=c��3iV
yA��V�ͥ>�׭k�}���ΡO:u5��4N�H�V\a��ͮ/jh��s!a�8�mt:��	T^��+K����\�e��ђ�"}����O&V�zy�5�q����3�0�f���r� ͬ�����Ty\�u���	<CY#��
����oX:��`�_vU��(P�[��̤ص��˯�k��c����*��{�nn�|yR�i��L�{݄e��Q6a�-{F�Y�t�s ��p�A�ܹԠMa�еi���_7^y�ϱh%�UTPE�AX�B��F	j�UJ«Z�F�E����D�TZ�UV���T�m��+
�2�Q�Q-(�mJ�TE�
0X�[Q%�EPU��cYUڠ��AAEkT���m�*�"���J�Ɩ�1jڈ��-�1�Q+F��j-U�[*+mQ����"5�TQh�DDb��m�"��"�[kT*"5j+U���k*�J��ilFZ�R�Ub�ڕU-
��b�mTUF �X�V����
�TZ��-��(��E�*��DX���4AJ�P��*�[l�ڋ+QE�AA@m���������1+V�0�X�JŌE��QQ�EU"0DX���b�Qm�KJ�V*��)K(�KUbőPQEA�V�kUUV("��V��iE��#Z"���eVڂ���*�����۾2�Σ�����wZ;.���97n����q1�w��&ڮt�m�0fGu|�eY`}x�>��Kه��}��=��qp��ǿ���g��ꁆ
E�h����'�3�J��5���~d�c�=32'�W�&�{��*
G��5'穉�Nk��wd��Ğw�|@�w��i���8�^}~�y��c�̍>Y���"�� �(ϓ�I��Ă�Ϙo˷�C�pϰ�&=eH�����m�2\��~�s&�=Jβy���0*O�T��w�6�X�Xbx��� _x_)�@��c�&�����?>��A��j����1��M�g��m$��y�Ag̨~Cs��m ��V.�S�*i �g���6ͳhbOo�����Xns���aXT���&�=D:ߍ�e8�;�Z�q�I�H��y�h)��6w[�)c�}b�Y�J��l�{�'�����M$�:�OP�����X~k?%fҤq�����<f��sO�u6�/�h�'\u]�V{�{�_xt�� {>�vM�T��9ߵ6��d�
�gr���q+"���!������C�h)Me�i=d��?2_��&�̝L~O�Y4��W�6{f�o�
��	�6�����Hd��A���Y�YW����$��dwd��y?w$��I�;�l*Aj��5�
~B�bW�{�z�f&�b/p<LH.3�n٧��csW3�LzʑO5I��<d�������y�s_.���}���������`T��|9�dڿ��}�i"�I��L?O{��6�^�k��������o2'��I]����6��eC��ɤ��!S�j��?&#��oig+'鷛�Y�������;7I�z�&%g�T���7����:�>���i6��~��m��_{d�;�<AH��>L���3�Jϧ��?'�Y6����`T��#�A��u�C����{��m��cNk�(c:� ��yC�Vg��4�xȥC��=�� �H��伤�*�d�6ϻd�O��m6��W�Y/s	�*A|};�jO��)	�t����~�S�"�;c�"8�}��w�p��]2u2�01'�W��l4�~`T٪2u�1v�8��'�Ɏ�X��!�>�$��,�PS�Ty9��R����!E\�y�bv��KG�Z���̈�C����gw!�Q�#E;�3�y\Ƴu�� ��:*X��8V]l���6\.�}\r�o��;:e�`t�����E�v;ż�ehz%��|7�>�X�792��Ǖ�r}/	��SK��G`W�'�����r�sؽǯo���Ax���tM�����;ܚz�$�l�<7�h�f�.Se�d��Y�y-��~`T�O&��%W�w�1"�Iǎ��,�J��^S��Ă� f�-����|�f�p֨����$YCԕ�I��
��2����'��A�dY���q���c=C��p=a�bbWya�%aQeO�1�oI4�3L�1���'�����Q�e��B��[�;v��;�)c�0��
ͲWg���잲�����&�c:�M�>�c�����~��,�T���p�=M��|�����M5�J��f$��"$�v�� �"���E�-ע>u����3l���wvi4���*�m
�tg���'���?_������S���6��_Y6w�4x��Rm
�u��i��Ý�$FLz��XϤ
>���y�p'�r*�<G��g�������t�Z���a��H-f���
z�d٪� |��OXy�x�R��S�6���1��̆�Y�Lzʇ��`�~J�̗�ާY6��A�}j�����#�vrl+���=���B����Y*�2vw�6��LI��O�,ed��Դ;�6�]0٪~a��4�X~��M`T|ʞ'�*bAg~�LY��2s�ɧ�>C����M��'�� IJ�'ytЬ��=�Kӷ�>����R(%a���i<}d�g�4�I^n�Ύ��CR/9O�4��g�S����a�i��,��_��I�u�<��!�S����>�>b���K+�|��o����~�;�~a���S�����T7��ECi�'�ֵ*�J�Swz��+;�&'ڤ�i&��R��l�B�z���'�H)��8�N�~2}�ݟz����ѿ�W����3����=�J�>�*M��;�~d�1���&�#']&!���4β6ɾ���Aq��6�?PĂ�Ӛ�?51
�_w'��%gS��l�Ҥq���H}�ל��%T~�7�
���.���{�����6}����O����>J���q��/�
�}gP�VJ��ry���S�1���_�+%w>�5%��$L���6��I�8���Ag������/��hRל��>9�q�N��nm���}\k�NE5k��᳞�1s��Y�ծ���[���)Ky�|nsX�gwŚ����}I�;��t�o��t�XйǙ��[3Y���E��eogn����#��x�[M>�I�Ps�j*��=�x7��I�m�� 2$�G�!�,���c-����1�����m �0���6�H�q+>La���La���M�RW��=�6�HT������"͜�5S�i
�3^��!�XT�ٙ�%^nv��+v��0� �����ٚz��4θ����
��q���Y1��0�cg�5T��J�yN��m �C���m�����c'YY�l����M���E��*6���f����q?x�� A������ɷH(y�a�R��=q��a�&�1+��Z���'5C̚L~@�wH)��ɉ��gCV�>�$k���Ğ�$9�oٹ=B�o������]��� �$F� ��0�L@�Vz��u?%@���4�$�l=C7�!��i&<O�q"��Vx��zɈ�o3�����a�1+%W�z~��
E:����q8̃�v�Cm+��c��G�>�=+�'��I�پ�zé���p�|`T<�&!��$8s����4����|�4��bn�!������Zi4�"�Ļ5��'_�1�;�,嵧%�%oo�{��$#�r���4��(t���R/�S�*k��f��5�P8��&���ߘ'��涓�+�O��+Z�g�Xo��i�a��������ȥ��07e��u��K���d"�O��f�RVY��'���,6�@ĩ>B���dRm
͇�d�k�'�H)��� bT�&�s�c>d�J��ϵ'���C�R������'��J��_<���񫌶��{X�~� "2|��ˤ�ϙMe��Si�6�Βw�1��َ�8�
u�7�m4��Vl�0���<J��~�i�:��|���$�Lw����E����j���[��E-�����qK��Y�&$��0��zəx�����T*VJ�6��|�hq�� ���f>�}�i�ọ`W�O�I���I�����q�C�>Ld�9�L������HI}'��E�����ֵw��~a�Ϲ��Ci���4'�R(��EaXTǌ����%{�<-&�T*
d���Aa�.3�L����d�'�C��{O���G��=�������s�SJc �,g���~�#����~���y��_L�C}���]��y6�0xX[�;��ES~ޥ{>�3��|;�L7dpML�RG�K�.{B��۝ԳP��� ��f��o7}��l`�7x���s�>�G4m�ja��ٚl�ů�Ω�Si�҇�� <;f�:��O�w�%� AF��kP:�:�<;�L�É�<�|��x�_�?޴mS�bA�;�z�f��J̆͜��c+9�<�4�R����)1
������H��E�L�?a��y��z�H�,����1��~z}�_Y8��Ss���~d�Ǭ��&�ɩ�y��H,���;��O^�$�7�z�����<��v��q<������޷��ue���8��U�������|4�(�>�J��c�����~Cg�m��P:���a�&��l���f����I;�4��T����ޖ�*AMO{��_ω�<�w!��N�dBO?~���r�!�·|#���$>���6��8j�|��^o!>a��m�|���d�M����̋'$�8���D��~�� g^A���#��ޯ|b?f�+WM�<L8�}��Q��	LՁ�w6�̕�̥a�1��X}5zϝ��
��L���g�|�+>a��}?Sl�6�^!~��~A$����>��z	�����3o���ls��[�_{�C>�>���_��I���FV�tO��������G�&�'��{AUY�}9��٪��^��Gc��7�k�p���~-FlIN2c4�tn��RP<2�/��j�|�+K�K�z���=�ٞޑ2���e��o8��}S�e!Q�b#`q�r�b]�6xrY�e��:�+���PO(ㄩn:�9nx��c��j����V��4�ZNn��#ȅ_U�W>eg�g�;"9|���0DhJ�EuJ�+�Lh��ηH�n1�^u��ʐjzw�Y��)A�%d("b7���h�'2��Q�]s�<m��E�쵭�����smY�t���D%�N�ٺ�ڭW�v�K�n�o��۾�fHw>V�%Un���%����	��Ru���)}+:+���8-�a�.�*ck%��G����¢�%.%Fd篕B�["'V�t��wf-;�����O�7���,e.	<N�>�R��M���.,�JV�����I���&�#�(���ﺅhO��>�؂9�R�D�2-�^1�q^>��މvVT�{��Rgf𔲴�Ǣ1Ɲ��4�YN��@��T���H!׌���}[�T$��J�a�t�v��B��7���A/��\'t�7vϬ9�pX�Q����ϭQ�����ZH����7U\�X�����Ȁ�;a���0לV�\�8�PdH|!"6�F5��[�-E{�y�yY,k�����E�U®��
�n��_��
p�4$]lN���ez����˖��Ȉ�+��X�C����ǃ.���VY���g�f
zXܥV��z��w$�gP9P��0CjI���2�8`�u!�����r,�)�"��l�[ ���l�l+�T�S��K�Cډ���j�7�j&(_��6� /������H��X�h����[���Lܑ��b��4\o�L��t9a��X�D�n��N��*�04�7\�C�]GԭC3��ߧ'�)�˭M��C5��
0-D[)w ����R|t�h�<~������3�wn"���zV���>���z����`����_cz8J��X����q%��,�ɣZ:v�u	/�� ����S�Y��i�MA��K����.�5�L��]3��,m���ul�V�^Be_{�͵�k���w޷��t''aۈE����)m��Y�9.�1}�\L�X�y˖R�a�Ӳ��w@ƪ���C���B�%���Yӷ-U�3��wT�=:�]�c��v)�!O9��~��q��v幺*&�����t��_�E9zR}�v޵�OPm��7ʽ0�)�;�W����q2�jw/-�U�����~�.@W�4�Szp�^J���#�R��NP:~�6vW��[��g{�pǺ���s^s��=���`����}�d�����+p�\���BG-�])/tu�i�e7Nr/�k�T�([�g�j��^��X�`���n�|�|'?ez2����xz_�e�ʔAi=�]Ҟ���
���d���7.��])ru(u��a�Pj�\2���X���
����g�8�[飵n./l�>�~NnCu��r��.Ig8��K��YwK�o����[{GX���q�[g"wb�M������K9Ӎ��� ڭ�)=]������	�+Q��t�%`��[#��'�f�꯮��l+�ݸ�Df.}ã%��v�h�plp���0���չ�%<�N��>�x#f�c�j_�1W�uM�כbZPg���{��w��w`O(	P�M���������4�o:��kj�(��Ѹ�f7�(]�/�UXu뮇��Ҋ	8v�ī9Y�#W|;��x��ˉ�D-����c�6��|9��zsM�Оg1ު3��t�h��� ��P{Y���_rʍ���v�����R��jp!����iu
<�:)���=��VK��tl*b��-m�}��]��|N�|<"Ω+���Wf��#S�r�E�^	��E�mەn�R�M�䮂�{f؝Ӟ޺F��9L_z��/�k�_W9��T,K�.�����M�rF�߼�q#7K=5�RU�SQ<�.�WT�:��m����	��Wr=b�{-M�h�/��U�Z��颟г��.>(�:�����lX]t�Z-9WY��"���U!�EwT��*�6f6�[3�Vg�BU#t~��  58��x�V���w�2���2�Dv���w��sChQg�g<���[�ބ�$N�~��� �҃ɪ��B�g'���Z�.�2LUK�:;5��Kr�4p���g��#�׭ۥ+�e1�.���a��cZIFmn���q��S��*o��dLjڑ۹��e�.�s�gk8.�kVb~
n1W��3^�^<{6�0w|���������&����xr],m����ݺ�'ŧsF�'8ͩ�4:f�ׁeni��)���;��!m�[�v���k�35�؞h���m�BXwt�z9�>൩�S�,C��l�-̹v��ɵ��;s]*��5[���*�*�\Q��]r7܏��SXby�Vwf�_�Y��riP�^͵ԔUϐ>d��-�wv�No.�W�����Ʌo�J���u�8<���x�M��/lvN�r�B�S��B9ȡ�+b�3��^�u�B�l�^ S�����`�K7�k�����U���ڽ=�2�nF�ZY7��+K��0��r�	KD<���řn�)�-�|��v�8�!�Ӳr�y�́3�!��  "�o�J�N��;w�]K��z���x[Y�i�e���Ss�u,Ed3����=৽��ۣ��
�V�б�v�����N����i��o:�P��'��c!9��@b/������mۚ�}�׉t�rx�G<�̨ƧSKR�ۥ����auzPK�_!7Ȩ���!w,�m��
�ʕ\���O{�Ϋ~|�U�n��|o��i_�:E�U|��\��;aS�lSt�u\��}�ޝ=V�(����	��b��e�\(ΡOc.K�FW$�[��h'���N�OH�V	;�P���^�HMU#q������G%�6�c	���sA�R��C�o���_nmi��Q�����eHyV^>}�ֶ�q�M��g��	�j���W���Y��Hmh�9���wbD'�$'5eH]�h�n1�:9�c�\|�����K��[��쾫�hv�y,��ĄO��^����7|�BH�ըE�����d����nw�F�\��W��r�֍�����S�X�"����Ϙ��+�����5�����7r��x̊�v�٢��|�﷬���哻�e����_���fcW�ܭ[6���sNf��k���W:��r�ƞox,c�~������%���{+3����x�:jY������yo�&��5X^q�<��qw��A�&�i_5��o���C�#�|��fK<1LZ5z���*!���핶3�qV�EБ�^E���vxf\�{ilM(��mi�Q�m��Y�+/��<��q^��k6��=�쩺�x�܃�}'y�T�u8�Xq��B�}�Dt�xݾ����=Y�u��j�$�}��|����$lN�X�����1�N��p��Y������ܼ�=k�ޜ�]�q]�>��_��Ω7�Y�:�]�RNm�َ_����i(�3	ws�N�vm�K���7AU��X$��Ý]ʴ��ϓ���G��)̀��M'`��N��%�p�Vg
�T��f��E��vç�ڴ8��GT��,6*䷕5����QmgL��_��;�Lc�ĝ5�	B���<3&�2=���V70fC����&\x��P�uԗ=u���Պ��֭P�k�wcw"Ā���旪}V�h��5	e���z�<���._�W�]��%@e��/������ԻL!ɐ����E��g_��յ��{E���T�u���Mq�n�Y/7�A�Xq*��֤wj��KuTt��r�x"�1|6��̃(����t�Dh�g:��7|*!Y���oV���X֞m@�b�u�/GZ���Y<Z���;�x� ��.�͊�j�nn�PÍ�Ϯ'��ɱXL�7\]VEJ#s/��օ�ɬ���F��ڇl�.5c.�׸�OT糊W�|;jas2|���\5�9������������+�8)��Z��)%��Ĕ���u��:�e�5p��.���t)�AV)�\p*����b�ζ嗛B*�c�K�������U�rΟt�J�#���u�nku�V�U�Whad��&Y,3�u<=�1���3E�T]Y��z�NU�|hJ2f�3�6�&�E2�=1�<ʳ-�-벷~,$��0=�Z����*�߻��]�*gu'j�oT�MV�EF����\7Nʒ�8'3-l�I􎯭|;s�j��5�5�	@_wpX��Bs8�����b��N$'o ���I�K�f����Q/yi�M�o^�����+��U��<�o�mGP-VB�3��yc ܻY���.Bw���2���4�x|1�ӿ��P��	�����vT�h/A��kك��;�ޢ��{������7��uc�|�M��!es�[em1igm��{ ~�]gm7{ǡ�}N]��Ji�b�+���U�.��:��֖gVG/,��k2�W9Ÿu��1�t�K�>�u�˗�V(���E�L'��e�:�=P�!mZ�;�D�U��v�$󑳤亵f.6�J�}��p=aI�Ջ��B�3)�W�iR����i��謔&����pq��`[U�l���nV��e�WT�Q���*IC1��9�t�q����Pl#Զ�s;k����y�>�����b�EƸ`�y��Z,N[b:N�j���e�۬��<*���b)N���0&8���#�,�TX�a�[�}b��2Njí�Gs�;�l�f��:�E� z��� �x��5ү�/)MwL�y.nG�s`;V��ۊ�4��5`�d�2>c��3�G��8�	��x{���"\;נ��d���ph��c�|4���4)�{�z����"��7�<D���l�iXX�`eq�R:�O+�tEE�@w��Ì�i܆�ں^֨#K*ēO���Ջ�Y|D���N�-��J�������}}��+�o��³��n8�ϻ�vnҁ���l��ӃR�q>��dN.8�Yj�vm����F׷���ʊF[QTV�QT�[J�*�ԭTJ�ADbm`�EZƕ��ZXČUF*[Ub���ŭ� ���R�iE"#--B�Q+(�*""0�U�ڕQ�Db�kJA�UF)Z����������ke�F�Kh�+H�Ң*�l����"1R"+���m(��0QTcl�1F1�
$APF�X�-*�EAF��1U�X�DDQADbĶ�`�X����"1m��XV�"*��������V"2"��[e֥F*++�U[KQTQ���F�TEF"���`�DT�,PX�Q��eUb,V1`�*���%j�T���� ��	mQE�EDD��V"�B�J�*6�I+b����$D�Ŋ(�R 0�D�`��U�
  �물wN���TC֦T&��^v�/z��yh�f�to���E�|�Eu7��ԫS%YR�M]8�唺����{��`����]���X�d��>R�F;��&mw���۹��H��m_u��֓R��mz�Ա�'�*�nf廞L��4�iQ�V �����i���3��8"���� pX(N��=��mL�����������C�	U�o.����3b�Pݑ�VĈ�C��ok�Mo-�7;.F,�C�4���0c�'G)9ƍ�;�0���lO����{��%?s�c<�d��d�� >�5�͗n��rps�=Q��3C��g�����q($��^������4;r��|lg<1#���ʄM�V%���wn2�����̾Hg9���a�z�(�ПsG!��|��i�9�sM�U7�8c�9eQ̘�Yr���#'W~��R�w��}
�hg9���f�UKq��+�d6��q��sM���9C�oW����ˈ�Yy����7�8�f�U{����k�9(���V��[F�5j˰l9��s9��|�ܲ�aܛ�;����U3�$h��^f�ú��[�ƙ�-	�.9.:X�o�q��V�俶vIm������KN>�=�q�4,�S[�6*89�����݁}���LNcRk���"��K�z��籴\lg-s�����]E%�U5��[z���,)��
Ry�t��}��t�Y
����K��]a���-׉p�1m���:rm�|�ŉM�r����&�d}�!�o���_YN�W��ɹ�>���=����*�(]��Kyi��=��9��>���|����"sԵ���a�b��t篇fv�����b�'�Q��ss��ynj�:z��*�o���	�Nf*.w����
�%�Xȝ�����N��4Ը�zgK�~H�����,�v��v0F���������3X/�	�׭ӊz�6!k~n��+"@�Z]�-j�����h�����՜�˺���v� �=��q�Q�ʈ������]{�8;}w�v�����iSۮR|[(1��'8ͅ8�ve�[�uP,ͩzL��j�:g��驮��֕f�nH�	,ό��c�Q�8(�nJ[Ȗ��b��ż��+WS��X��%G.��1�Y�|�^e����4�Û}XB���ӷ\�ɠm7k9[Z<K�	��)L�
�gL�U��"��� <C�<�|kt�W|����yee��x���k�34����{g��9�sZ)j�u�p辿��/%[�e��2mV뭰;Ps0�BC'����V���LJ|r(xbG;j��{�bU��3���Y����#�*M�۵��T�ls�:�R���,��	^��%���<Ě�%#[��]9�mtT��{/��=p��۽
ܜ��_���������)8(M��i9�.��zdl�V=+^y�}c[�1��Ue-Xt�I��iff�b~0���a��B=|����.Sn�sWA�gT�V���U�E&��$^�lr��PX��מ�}^���|�r*I!3�u���n���[�o�2��WJ���\$�*�)=֝GF��;��Z�V���T��H��a��4���]�:z�%p�o��ҩ���Ȼ���}����dJ����w��ta4��b� �o�0�%������k�S�*�szb�J�F��=)�k�g�����^��>��;r(�-�{9�������"*�Y���4����Q���gvu��ި�*�qQ��jɹ�x?W�}UV�21([��n>�/�{�M�}�^O��ӥ�!.���P'ΜC5ؕ��a�����n�t5v��y�'�O)ˎ���V���v����<�S�:�J���'�$ݯHY"���}�ֶ��q�y���,�z�z�(�NM�ل�ƈ�1��`�
ؐ#���No
���h$���|�潞AF����{9���3	X3�Z��VZ���ّ3�&��Ɓ��9E�INea�%4r��8(s�4:jX`j���򽖱��|h9�y]��d����ښ����e�5���OJn���ڷŧ��z�g1�ޡے2iPޕ��Ê�(�Б�^E����G�;��1xSb�f��sz�m�%Y��'��=�+/��<��qO�mnԺq*�kc�%�g�*�.�b���H���z�tΣб�Kd �jTmڊ��u����I�ءʮ��w|�D���)�a4�������!eZ��a �B�Rq�ދdD.�*&>�z�����	���엙�A���=C��#�����Z��,=5��S��Yp�\KH�Q�aGF	�x	��iM>z���d��-��2��Q���A�b|��>{l^�T��zwՖ�[�/<�k��յ=�]�d����n��i���^/�-l�O^hvݮ펑��C	��T���7����/�=t�Gv3<y��}�v^�or��۷�@_"��+��L.��OSl�B8X��w,me/N�����/r�����j�	Gbky�9�v��M��z�v3��7�%�/�r��Tۙgyn�	��|�^n���Ř������v�Ϣ�7����5�}�S��JGKݳ٭]t��l��e����-������9��#b���8-��_
��Qs��$��9/�p��a�eیT������L�V�[�P����!��@~F?Tžj�9�ͪ�޿VsG)989۝3�m7I�1[�刀o&ńt[����QnITp,V��a&LLp�	-�6.�Q��(��;�%a�{t�$�<`�ۄR��u����-���gAԺ�r���ĵ!�71�N"^�xx�
�\�>��=�w
�-�.P�����5��19g`L���U}1yZ�:���S�F���W/o�J��b[cZPdkょ<1:]A��&,U=�v�y!ٺTZ~.��X�ku]Įη��4硆�]���<�7X4��Zuw)�]6T7�a�vxfg�[�����'U�?m���j~�cU�S.�t#ϜZ���{�z�������hLO3��zޫq=�U��ov��I#����'~���>K�a�_K;jp!��5a�K�����ni+bZw�zH~�>��뎔�z-�6�1���q����qx� ��8B7�����O�dʣ:��8�)�~r��)g&�s�(*�t�Ͳ���dU�m�n��*s����҂U����U��TRĪr��󄷴="��cf�7��]X��W	7΄�U0���!��*$~��o^)�ɤ���5mt�������k�W���%�Bc�Kl��i���%�#���7\	�:�Ü�n�;!�݂�U-�{"�sk8�GZ8Mܮ,)�\�T�7w�#v�n!���1ٸs���ǖ�S ���ᮭ�SUwf�f�{-�*XV�nU�[����\8�sꌓ��qG4F��t��C?x3�jk�Mr���H���9�;I3���r8,w�zG-u��׷�{.�_�r�s���^����8�=N�`�M��� ����D�ܹyQ/���ɧ#v���}���fַOo�g���DBC�+�]��ۻ�}Ko�G0{�Dn]m��V�딟�1<���Nq����P����˦#���fg��ɹ��`~7��X=�)Z��d�=���ؓ\�^�����D^�<��[\K�@5�j����˕n�Z�6�\䅴�VfH���&y��l���SC_�vc��Vwd{�~�g+9�����W��R��h����wo�w�r‷�Bj�/����јU=�׍V�kDE��{yr����E1� ^ꮙY�/Z��7T��'���b�ri��yt_5'ojX��S�z�����qҵ�w���g��1��d�c���kgp{إ��wj��z}�.{�*u����Kӷ+6&Ы%+wd^�xς�X
G�*E`%m�,+�sB���s�M�K�JՑs�TR��t�;R�j:ٗ[*�n$�r�:��l�KnhQ�Y]�֙��ʍ�(���i�� y�<��<�ٽ(*��7B\�(>�b��7�8�M��_C��O�9Y˖V��4�v�5AU�����d9��|��|�-�la��9O8��ƻ�c���kz֮�b�� ����ޙi]G@��o&����9*9w�`&�ٰ��m'`����U��@�{~�����i'�� ������a���_{�/�-ex�M'���K����8h���:=�v��ӄ�=m���eo�O�N�r6��=�Ou�q��OD4剾�Q���i��w�̎�w��ڑ�5g�Ϻ�^�/����'Z��a�G�T�^�/���lF򒗵��"9n_�'xV�sA'��koLV$�U���[����tr�s�ڜs]3	X3���>��Y��ܥ�w5SGgA�m���ͳ)���9Z����L>�.�;
�ؽ'���8vV�+��E	˧b(�YP�Uwz8��)S����]O�Byc���6S������FWJ墇� W-v>V�Ա����̮���G
�2��o�)�����Duc�SXyGg:��X�xx�WlJ�m�ٙ�&�ޙ�_ �li	���{^�O��tR�v�ܻȖ�Ҳ�X����riV����Ê�JC}�^E�������q�=�<�Ю�(�
r!����NFN�镝���<v�FÑ31�9Z�y��ؽU-���q�t�u7;^�g�b ��jf>"g?w���$nο,}��u*�w6������*𜝄n!�^S]Iգ�`����<V�F§ZE͵٫ؗNإ���]эT&P���*�{��b��<��c^	���I�`CV��-�M����ρU��WB,uS��Ga��{��	�}'��֣�_��>M&_pZt�y�K�H\I������]�W.3�<�N̊�M�R�G��ɏ���A�R(����qv�K��:u����X$��c���T {s���&p����m򄙔��]E[��޴��WVW��ό1���^\�M*"��H���cR��Nw�,؉�jV�O3�r�,�2�}�q�&���p'Y��m)�ê>
������?.�%�ޖ`t��=��Ws�9I	{��ӹཻ����L�ޝ��6��av����ݵ-qqٯ��T)����":�� �u���mL���&�S��+)1��b��wpO_0�19s�z��!'0��
ؐ#���������u9�O��UZ��՘���یT���v��3	_�앰����27�i���J�t�g��Iܛ�9ܙl����NN
��t�>ʌ��Z��.�3�y�=�'��5Y�j>[I��鞴�a�=����Ҟ��֚�SJ�5������%��W�4�y��kj�(rKت��'����R�A�g"��@�=^9�
�X�g(g9��]�~�_�0��_t���IlȻ�
�t�݋���Eڊ��f�a/�%<��@�~z�ߗl7����hv-x���ݻ��y�q�9T��h�����&��O����ꊁn�s�BJO:[m���NʸZU��������
ͷ��9�G�^��S�ѭ�NZx��GѢ�̾��t���(����J�ޥ�,�īw��B��u+�#��.!��\x^꭬��{��]�	�uc�/�՞�%]��ݽ��m%���	b��CM��v������Y�H�n��ysf�픩vmg>b���õ��"m�=�n�kq�������g3)։����M�@��is�
m�tVK���K>Z7_X���ʈ�S_r�%!C�W��6qٶ�C)�Փ2�6�Y�Q��������ds����^om��Nʓ�iN�'U^���`�bx��s�o2���rR�MgC�5�ґ��#qI�8>�P�l�))��]|0����bv�Y�ۜ�/���m^�N�J�g� ٭�{Z�@f��:��S�i�!ۖ�,��m��G��ز�D��V��M֬�qh̵��"޳� r p��)��_vu�C2���+����8�E�m�p_u��WM:�9t2��Z��V>U�r���\��h�6�6cr�Y���\��/�'�WY�f�o`(:8��ұ�'����qe��f�o��ֈ�{z�b��k������B�ڋ\7�OCx.��c����f�ǈ�Z����q�gD�4������M���*�ح��%��)MK
3f�x�yj-_n��9֧wR��4��v�qS�
��m7�3GXRc��T�QIϬ�ɍWam��̬z�թ��%�v�$��`n�l,�ۓ;(MX�ٷ�6`	x8ֆ��f��v��GWǘu�&�Ew�WF��aC�#?������ʷgVx#��8��b��m[�޴��������P�|6\%�8�Dm��;�'��mdE9�q�/�
���zu
v@���U��v�7��<÷,������>�%�m�X�2���A{A6�u��JX�1�����|�.U�J��A�f�QmJ��%��"&Z����yd���o��Sùv�;��\�83Q�%�F-Ʉs��UV�*lWD�(k�|+-����X�\4�L�Ք.��T2���o�M�FC;s1C|t���H'�2�>83��\ n�$�m���d�דy��Ʋ�v�k����b�k�2r��e�{oo��\�%Y��JL�����(t��<ڱv�0�R���*�H�"�q���غR{�h�/7���0�Z��Dp�E+��3hY��h�fևz.8z��&�X=��]�ݝo�D���^�`�Q�&�Omf�t�,\�yM��:�Mr��އ\�9('ۭ�K8sO�o��Z����`
Wfoe� Z�����ոB�e�+�X5��'��C��&���gKvEr�+��*�>{�n�
����9��h�pJ��*n��	���]���:i
]{30�E�5]n�DI�Z���Fу�l@j	��R{5��=�j[�9�ˍ�֯���ּ�I=�Yie�DU�jV1-*���U��UETV#T+
��TRڊ�T�[bʕU�1ETF*��(�A�R��1E�P�1c�eTX,b*�dPA�*EDE��*���QU�B#F*�DD`��Kl`��X����"����*((2,[Z[J)b���TE�UT�dEU� *��T��E�E�E�UQ�����QDDDcb+U�
DAb"(µбDZت�1UD�*��"EdX�b���T�!YX֪EUATX�( �Z���
�[U�`��%kmH�DUUU�T���DEZEb(��2*��؈�*QdEE�UKlPUFFҖذUb�EUQ�
��*b�����V,"(���EEDE-((ZR
�" �x�	$��A �r��תk ��^e�k���ٕ�_Z�l8Nk����R��f�]�Gg��Gc9�ˁJ���%�؄�r�=���y�CS�:����eН�2T��$_.q	���a+�M�뎝f(����a���k3r�5]@��auJ	VGH�uWȨ��T.��_Jo	+=�^oێ{ю��珏��-����X7ʄ�U�0Һ���\:�:�ׯ�+�b�	𦩭�6�OU����N��k�Tp��Py9��{�N��⣪�����{�te?so�w�u��L�}o�T��I�p�2]7&k��q����6��6;u��^���[��;�Q�y�7Dta��uu7��b)Z���\�1�Rȫ.C�܋�پm��s8��09f�J���2��������~(v�t�{4��漓���9����s$��W�t��g��;�������W�; �ɡ)�R�Ǌ����2�K�͈w�&����-UӮ�;5�����~��P�H��|������� ,����@uhL2-m�{sj_�=���^�ddzf�:UӼ)6��t��&�Ͱ:u����T�/A�B���u��7;�l*�}o��i�w�#WZ�o<�my|k��"�m�Z[�Vu�&f+/��M�qgW�2�55�����h[@�hH��"���m��=̅FȊv��R�R��[r��7����Y^핷��9�9qV�Jj�5���jUZ@��r�x���E��l�ֵWL��wS���ݵyS�=��3�ʥ�8�Q�9U�m�ڽ�E0>�7;By��@��F��z6�k��ٕ��̘�gA'x���_��5n=�| ^����6�gNTtk���v��d[|�^%Ӷ)%W���MQ��+$��t�T�=&���������/�����T�J��T�uL��*h��9��u'ʡ��cndR��l--���Aaô�%o�;Y#��#����t4Z��bb�]Wΰj[�奻�O��8uY�3v�Fq5�����]]m����ojSں�w�wb�N�;�4�GR��D���-�4���-㡍!4_s�A2�(���e/����}�u�K�b��ud2�j��9�����ԩFQ�f�Z�	W��ʔ3'�����&��o����cN:쏫2Qu}݇�Qo.	v���%�FY��ջ�L�������#z�ƻ9����7.�3�t	��N�����;*�>�kZA��]�]RT<T�(Ԗ�Ss6!kt[�: 8b7��N����YH����*��!�%��y��^	����6��0���k��"럫^�s}�s��r�ۧ�Lr��5�i69�NNv�zK�3ՙ���2�Mq<*:R�����cn�+p�S|Î�m���|ls���X�\H�����[��W���r�8��n'�3�>��ug�=���)|��I]=�q=�bQ۞���=��:g�c�'��/g�f��~�T�ۺ�uKV��,4�j[7��Ʊw��:[�:�����K5���WA����0�{�I���~:|�#^��zj��;k�X�W�][���Ι�4���RH~�}�
Rx!�W�[V�g/��^���(w���[��x�
�ؒ��]�ne�Ty⮇/���.ܼ�c Q�
��]3nWMp5�P\o �.�v��T
�w�;Kp �	\�Z�I�wx3z�c����&TN	��Ȓ�kgd��G�Bm-]��۰*\9.��X��d��;ue<�H۩�IՉ�W�B9�g$|&��^	6���Ml�)A�z�`�*o�V�˛[rVv�u��t'[��|���=R�N�Y��=�p��g'k��:{ϫ���4���p_9��U{8ve�Ҥ+iV9�������S{�yn����o��n�U�M��n��'9-�I�^{��;�a�-<��q��ӝ�i�:�� ���U�Z�#cjm��ɶ��\�>�1����<�ӗ-�e�5_!����#��J�$���r��m��]�ͭ�P	�;
09��a+|��M/�_�=���\}	��!3dt��nc��L�X����s�*�����S�CՔ{����;��yn�z9]���o����cr�Po/DUDE˭���t�A��%:��v�C��T�QUD���Mί/?k���ɣ|��m1�wL�uCϨ2��oܙ����ؽ�]�ɓX P��M�D�yK/);f�\-��z�&���bv[޼ŏ�m�\�N���^
"ė��7#��6f ��B=Y�Ð�rP�E�\�t�szjb��6KM��d��<�a)���ף,�ս���Ą��P׆:����>��,J���FJS"r�m�:�k���iq�D�hj���觉5w����9��;�t�e�sR�Ɵk=�=�Y�s��R���Z�7/��ws��2�Zn�sy��q|8�6�~��ݑ=��{��@��|�;n��o��5ӷK!wV^7.����J��<����0�20���=|��.qbSm­ig5{k4:1r\��[l����jmA`�ubОՐ�_9�EE$�@�u[U7�����{�o�?�[ݎ�&��p�|�����u7Ξ��==/kQv�]c��<�#bm"���V_k��OZ	tp�o��҃��6zL�xo�^u��p�f]���|o��H	�+L�t��gM�J�m���׽�{�}�}|{wOcz�g[�:ps�
���������.��� �=�r}��Hţ��<r��ƙ*ǳw�ol�*�r�Z��O7�}��һ0�����7�=׷'{��{�O+Q�x�ۓ��M�d���r�ۃ����79Ս�K}�[K\E�:v��bu^�)�r�I\�f�;:`;��\)���ė�S�k�ݡ!d�Vys��[���눷8[�UU3��k�K�W!�ry߈��&;-'��H��4���o����hЬ��\u��Im���s��8�L�W�`�s����V5=�R,����g�V%rIF�~i�M��mЎ��l��N�O{j��9v�ɞ;�5��垖ryd��R����k�9��^]�խ*}�̙x�<�p)8'�hd5Nbֺ�����}�H]W����cv������kSz���w�Vr������+,wS���k6���# ,�,�]k勷+6:���>���JGk8E�������}��<���[���ǝ���������O
��toP�%�|/x^�Y��n���&_����o(3}�N��1.��V��� ƪ��Z��ރG`��FnP�(�o���w��*�'2"�ء�V��he9�j	St-K.x���wxp����@ќ֞�s_.���F������[���L�6�vu-��-4�3xʻ����.�Vg:х��M���B��d�7}�d|��vD�h���n�p��Wy[���3�g�����3���`?'�4�|���M�t���Z(��B�/2��)��σi;+�����i��݇b��1�#�kzn�\m�LjWU�s���������}N����yD��!���(`hG�ڏ<���>J��v�����#n���yg��z�}��n]�C7�缺�Nb��
ߖ�6X���Ge_c�Iׯ��tRv��H.���J�zs��6�:��j0B���N�9	՞3�c�L^��W�33;,��[ã��vZ��FPNq�
1�t�%`�ϊ�4�\@=;�ٌ�ըl�e��ɗ�٠��|r�NN
�<sC���5\X�oj�]vl}��˹����멯_ ⇛b@i	��6+���F�P�ViIkn7���Z`���ǥZ��̉�f��3�qV�E6���j(7����oZ���E�W��+�x�N�=�����Ã\,y795��/��VvE}nN�O�uԔh�w$U�-.-7)}}%s���qWZ�RW��f�M�=%*ξn�3�����]��N�����\��.K�,�j����>�n���1 �U8 �ޞ��kWU��a��Ʌn�m�3�8�fy��ܧ�R�w'�y\.[�Q����&�jls9 �=@�*x�'�*�P���S	�L�G..
z�d�C]$��T��Հ&���uo2r�i��}u㜨NNД
p�Z�����M	Z��צ�q�&wyP���s=�	�W�tcOj�4��W%.n)n޹��#��	�Lגm؆����ɾ������81<کS}y����T���1�[쎑|�|�r�pM'`��=Ю;��cѰ��[̾Z�G6L���u�7O��ݥ*%��D�(��bk�B��{]+VrÇX���X�_u`s��ڍX%�v�y���n���שn��9�V{��*:X$�#{
���Q��E��ˮ���N[wU��]��A�r��`��o��ds�UG6���ޡ��&��p�-�j�tlZ�Y�I�F�`z{�r�DT%�������=B��p��O"��hoQ��5hl>��sH���r^���9�mf�S��δ�AFSjX����L�0rރv&�r���U�� �����%�9��]�S���b�@�.Fk]aC��8�M�W��v`sAL�Se:�8��z�y���?�#r�m�Y�71�re�����s���b'huI�}]L+��nf5Y����u���wt��7-�P���ݼ�Z7�RS��gy���P��ژ{�r��+��~�u�m��2uiN�`�}Y<%����r�-4'_�׆:���[��g+��K�IL�K�9��x�N�u�U�c~��	!��9�)�M]�k���љ��{�n�R�ݭ�[�\ѽ���}�L�ړ=�r�޻�mnՀ��QzmD-SQY��g.۝�ˆn'��ɫ�w�<����^��>��^狟���`�����H���,JnO�8�	�\��6�9WP dڔ�پjy�哽m�����!�]ȟc����Ϧ��.���]<_���Gp�����.�w�ieԫ�Z,q�s�k�Sr�#K��"7��o"���u\�p	Z2�����N���+=9q����l%�\���k�8 D;���5���9k�ܮ*U�Q[�F���4]t4��"�n�m]��-�Oi��v<�UJ�t�����X[�ɸ:
�_,��O�u����]O\u�Z�쉧�k.Ot��q{�r�s���]��OP����E��[��H\�K�`�0MW��[��(�>Ζ7����%�D���g�<!*�wm�6.w���(uN���^�ime?=<r�=��7�V�Î��B ��W/�j���V��_2:�y�H욳ҹ�XQ��q���=�,���;.iɚ�}���ʵ�������
ؘkr�'>�*}��h�&L�H���T���-������'Ω�4:f:����愧�J��۹٬\1�x�a����2._6̦��G_<sB:��j@�����ε�.8ͥ��N]4�l��W5�T;s^m>m	��(k��v����s7l�*j�+E��٬MvP��2iV����zܨ�7�SW�c^����mJ��Dj:F^�����R�&1� �*��6P�b�n�K����\{'\��oc�]�1k��Q
�X�� >|��Y����@��27O+y�·"��ە}oS{Iӑ9�����f�r<SG�#y5�n��Ǵ���v��S�p�Wc�.���1�m�3vg^c%�PoEl1�Ǜ�9�{��i�qɽs�/��:��sc6Z��I��queM�o��&�U�=��s]�<6`%�յ����V���\�7�ҭ�8rG�(a�Y�c���`��ř��ۼ�-TJ�[׭n�)"Րo���\6;F��7�1�!��Q�HS��W*�7bLTS�vհ�dB$X�$�n�!�:�^Y��3@�oI�x�T쁧we5cwǚ�i6�^woSsB-�7V�b1���m�-��̮<j�tZ��q��em#�7��GP	v�\s�]K�Iӧ,ճ�i=dp���Qf���on��t�J�B����Wկ���\~br��P��ޛx"ʷ&<="��������tmL�䭀��1�N��TW����D9x�P]�	���Η��PUp���7���k2щr�-���P��>��gus�������c�����X�E���?h+�@��q��y뮘[o
įF�
�-���{���{��,�z���U�i�7�mڬB�.�W�������cF�u��:6�V��5�$ipv�(n��:`��j<N��YYۃ4�fYRʆ�N�Pp�-��n9�Gn��K�f1�N���֣osu
>y��=Ԉ����2$/Vmu.�%a[�)ݥ\�+�p�A�y������p�Ŧ���{�Q��ꎁ�n���
9>|%��� ��}�1�w
����{�BJ�wSh.����`u��v���+)�����em�c7�bz��v�U�c�]��h]Z�$�]Yf���v�,\3��-(���1�=K��үi͗`�<3���;xEHV.��I����Ov<���n��9�Ys*RڼVs��ӻ>o�]=p�ok�CS�Č�h���n�_[��\�j4!9E0�oq$���H�Z�]FR�clv���P_G��%sm0�`6�Rg7��:�v�#b�׷�
��a�rF�*�.o.T3�Y�p����Gy��grpc���J� �u��ݘB�((�9�ft����f��l��H���#b�
���˥�K3;a�����X�:��+)�2c�Qv�3*/�]�%��Ky-wN;ű� ���ijw�����,k-WYyƎ�Hc�\�O8�V>ٖ�8*}�=Y���Y���hWjw�����|�-k���5��=��/�{�a}�	ܡ�:�&@�y��N�(����>�6$���Ry�5|J��^Qk9��՝R���zՌ��P5qvm3��%����%�)�U4�Y�5��n�vŕ-듳o���|��Z�!�d����|�lDJ�1�����V*�[DD�D�*1eh��PX*��Z5�E�����,X���m�mB��X�*"
#R��,� �TbȊ�����ň �X������m�R1UF*��E�ڶ��E��X�#QB��
��Z��$��b¤�V�U`**,�c�TQ-�
61��V����XV�P[j���%d��"������hUJ�*���YX�Z؊(��ڍB�(�KF
�m
��,��hX�Ab��eHQV(�b��AV*1���b�FEF"*1VV"�*�E-�R*1[B�Tm�TA��edX�$ ������U��Qb²�`Ȋ
��ԋ
��lE@PT��dU�A�DeE`� �Ũځ��$HĒ %f���_of�\On�����3T�'u^&���l�c�8�@���u�e=&�K࡝p�<踫�+���3�K�#]�G����Y���W�ee���=pշS¢X%���\�Mj�U,>��/��򡸶�z�Ҕ�S}pr���1����wfRW�d�[�s��i�XǱ���d�7��`���(|\����^�DEKj��p��i[�����l�T����ۃ�uK�tU�݉)������@BV)i��I1:�K55���#����8To8X�c�g2���E-b������+K�2�iaõ�(^n)	p;�T��i(���W�����v`��_sg���L}�5p9���x>���ㄹf����j4@=�\�ym]G���k닛��@}f��8j�[3�K3�0�r�XoD;~Z��(�@Hkk׊s�'��u�NO�G�Gd����_{����q�ѱ[�ݑ���Bh��kԭW+u�v��t�	S�4Ow;�v�j���3zKJӝV�2�
�
K:�+P㾀��Sl�8r�ڽۙ�i.M��)�D1�-�E*�j�ˮ�\����ds���>M�˼�owJO�Z�t�}�Q|��(��^�:��;��+fD6t��e@f5��޹*���� ����n-P	�e'8ѷ;�0���+\�\
������P��gCk�����;v���4bG>9A98(s�5�_S٬���V��\'wy�̞��G:%���1��A�6���'_�8�o-���͇�t)K�̓�>g��*�nU&�߳�q@[�tu�`�׮{-�/��A��5�:�vz�d�V���#'y��z�� ���$��kK������a��eO3h�=G1E��3ւ̈��Wj�>��}eKS+J�����]׭��ף��[����<��t7�Kmq��in]	�X�Z�:Re�����t�:�]��-����w.7)co��n�:;�_!7ɔ�j����L'����4U.
��]���;k���`��]R����/�U�)̀�Ki=�R$��}&]n�%l�Q������V��u��jȻ IaJ��&�׽��u{��Q��-���@�1�D�ή&\��HU��y_M=�Bd�s��\80v�:�У��]7�%Y�N�fu�Y�^i2^�#6�c�h��G��9Q��BʍbgG%��kU�����l����.E�O��v�����"�WN���g�,4�'IoQ������OU�%@G7��s���\U⫵R����E�9���l��.6V��~J�
�_?�`����]4<����t�W��_WJ[wz�5��ڌ�-�p�j7r�3��p�U��C7�����*}��X)�vZno�v���T�ˉR��Z���;Æd0!��v�i��s@w&]�c�6�z�R�q9C�9�J��kWN ��4�5~3�<V�BwB�ec�C��{�+z*
b2p�,�[�8^�[�X7>60sȞu���U�}���ޞb��{�{!��9�,��M4-�>m|n5ٍ��fz<��6��D<�y1�z��s���s���^_��������"��s�����gEt�U��w����D�m��,뷗X>MS���k��<���v��A�n	��3��,q:�	ŵ��q��IS�^i�wV����6khKȉR'y4��9�R���3t��ӏ1ʖ���o:�o2$]�s磹[\�D���X��Q�L��ǰ��ql�[i�aR��gZs�r��-jΙU�/[p����W��1
���|�"����Oo7M�>�&�jR��ZӰ�lt�m���ŕ�t���_qw���i�̇F�Lb�K��������8Jm���jT�D�ӯwN�b}YҹZm���J���臱ûr�8䈕q;�7\���E��m�P�ܬ���w&����7ʦ:DC�F��B�pQ�Oy���<ս7VUz���>o�ߋ�oN�;�p�|v��6,��fn�U~���C�`2&��o'��ۭ����g����C֌e�PIks�uw[I�s�opHOj����=��y��q@9�.M��q%ȨMt-�o��X/$[R;&���}֣[�b��EEׇ ��Ub
5%���9��lCPW{[��O�xT�k�ܠ�s�E��U�X&���7(�WS���e��Z�ԻO�>o���>��yZ��H��V�oi-0�FP�Օ�_;�7��f7��mr̸�k�g�-3k�}10.Pߴʾ�leȚ�hP綶P���G�l����W�f�:�Fw^�f�RR�o:�cڙ��/q���%��y���j2��eE���1���x�;�Q�^�e�	+66z ����fySZ�3A�'�3��
���/���RE�*�fUE9�U��$��X�̡�{Cw��s^m��|s]��v��[=+�`ŉ߽ی��1#Y�mR��*��/o��n7�y5yf�
��
������U��We��y����^}���+;��@k�Usm昉�I6�,YJX<ڛ�{^/���1S��������w]�.�{���>>苫n����_�=��r¨��;��a�/�7�pZ���^���!��X�۰殃QC�����}}�j��~�]_o7d�.{�X��r)�EF�۸i�K55��7.ڼ�mJ���h�vv�v&&u��GM���<�֖�O�Wm��f��!�h L�L�)X�������0�[����3�$(U��� �\�È�"<�t�7�uVǪ�S��0JV4�î͖K�VxBGiV�|��h�:��<l�g���w�:��k"�(�9��ʚ��jf�u�2f yd	|M���_e�uǻ���L���:�;���h�m�sp{��p���Rݰ��w�:��$���u�6��[���t˻�4:WޞU���[��qsm��f�k32&�SbЮoV����Þ�i�^��$l�$�8n��6�<u��-yn�r��s����Zm��Ӡ㱣b�E�#��	���S�*�T���D_5����r}ݪ���v���18����@s��~�AO�{ԻA+޳��d�S���g#�jk�ɚ	�<������E�����LWn�\�������2�mڠ7]M_ �l4��z�i��kX�[��j��(0a�	�>�b��9����5?y:�=^ =[�cp<�n���m1>Ma��ux�=G2a[���9Y�FN�7\;-e���iqؚ`6�;�ŵ[��mM��8��wΩE�|%U'�޹���^xTwZ�)3�����[yj%q�%�}�m�ݕ��<���oE;����t�v��S�7�]�([�J��sDbuJ7��T��m��T��8Z���Y:��D����!Jjwӗ �++�=gz#��Bt/GD7�`���-ѮrKH��՘�j��Vv.���^׺gz�t�x����y��<֝�����9��5�Ѕ �ͤ�ƺ�oN�բ:Re��k��/t�j���qu.޽ٍ�>2C�$w' �ڝ�R�ud��B}|�ŏJm�5l%�3�2��]vr���{zw�:�|WP1ΦP����|���x=n��u��uV��n�շҙOU�:z�l�p��^�J�0ұQ�k�h���W�;���j�ncSI��#bo�>�e�7�p������%���+�>������Ы�b:���j���w@TB��'<�MtXQ�P�D�:�SqmZ]:��$U��c�aw�]��VK��Jo��WtC�������n��a&&`��m��)�s��'�8�7e�QB��	�����\y��q��Q�nݎ�:��"N���,鷺�G�Z9cw�s�*5\�%����'d� �����"�f
��J�N�!�k"�0�����<�K�GJb����f=�b����w]���5�Z{�Ճw$Tl�޵�ƧO�8V<��e�(�q R�B�g����䳖%�w���	E���;<�ݙ�ǹհ�γ�ݯc�)݅��+�t��[�fw�lN^@�U���j� �Z��v�M
��W�<�F����g4Ѯ�
�H:G�n+�տ
��w\e߲��-��v��֠�&���QڦM7B�_�ls�u6�l�Xk���ƜȒ�z���<#�����ChV>[�^��K��$Ķ��� �qq��-Fz:xץ�iڄ���pa;�t撮�$�X�݊�U�W��a�^t�g��y�$.�;eg���@a���'�r����F��,	�[=R�Dn�oh+�[���sN�uf�Z��P���{�>iS����w�{h#x�ҁ���N��2�`�X���]-o��>�~��S�s�L����]�����~nx�Ŗp�@싱�;i�
	}�H�������N��9��ޮ�"_v���Q�S�:�(�[Tv�D�DWExD�`TK�P�
�d��ڡ�ŚU�\;u>��d�����!.���n��;0��L�P2��@TOt$�����Թ{ݮ4#�B^��0�O-�+ͥa�j��L鎱(�I�T���~����21���I׌ȲI����5���_�rH��1.Z\���l͵�g�n��6�]i���=�{�N-+��EV�m?t����:�xbY��� ��"���N��8!�6J
2댧�+�l�r��H���f�uY��+���_tVs��mо��.�d�����VH��u)ˋ=R����t��p��R}T�y��A=�7q�EQ�g�;�����*v�Q^>�V�t�h����w��~>�]\�ث~I6�}�g1]%�q+��� :���:Tkm҃���G )��a�ebw��.--]�x�UH��3��N
���Cy� �'L�[@�:�Ȁ������brs]â0�N����|у���PdZ��S~�2��E��ڑ�;�	l�g����0����0(���!P[�ux�h',�\ѭ6s�k�y�GW���vl�rܺ"s��%>�l>R����[��vZ�W��������Ϋ��^5����y�g�|,ZE��Yf�]5	6;7Jщ�^�s�p
s�;:Q�ګ"��;X�Qn+�Tqӊm�@ V��c��2��h�^�z:»,L,�E�Sf3%�j��aUP�~�����'��lO��qd��Ӗ�7�z�0�ʈ��D?�]��N7�U3�$aD���d���efʹ���{�*��(��Gsm0�o,�i�;�
@֞��΍��ە�m�f�-�>;F���
Q}ʦ�X�c�Q;^�����"3����rg�#�n��p�k���}+h���U�m71]��b�ř��6�K����{S���z�Ԝ{���p��{{w��z�^�������4�5�#����@�98�y
���19�gWB$�ܫ�`�T�8��uϧj�o���.2�+(%��Is�W��rʛ�e-�{�s��"�3����D3	K-�8�)V�`NZ�6)�2a*yW9��]���/�w�.KIX�PKF�צJl�="�ػΥ
Y��!m+(�����a�љoC\�����^$�N����4��i}������,j
��.�qǡ���Z�coi���WWD��:�N�tX[0
F`a$�w[�/�֍���k�f��E���m%�[Ө;^x��6��F�s�qBܐR��z&�4Hfⷣy=�����sq[��t��[���)��g��7n�ߝu�8d�Ź��x-�$����B��lƄ���ͱrH�7�C�7�.���CfE���N�b��]E���K��z�����N?�0��nH�k=�\�u��NgxF9�ѡ��2F ��+g;_M�MӴ���c���|x���2�4���o1^�}�d�:o����3Z�=5<ڗ��%�SnO��6�bׄ���i$�zr����`һ0$0���z�kI>�i�rǓ1�E�s7�W�$Z8���Q��RT�]�֨{���1m�o O�'��ۺєT��ӑe{ݕk<��5�t��W|A7Z�l<��jD��O#��f�:zP����� �_�u�	Czs ��Wӻe/6.�F���ü�H:uI�2*��;k{��k"k5��)2˾w�;���y]���Ľ��u���m점8Kb!p����V6�y.
��2�,�+�=�5�*#6ض�S;�������a\�{33*�!Dɫ��W8 �c�:pz����u��*��&��t�8i
�T�S�3�ܬtV�mk��ɶ���u��ofY�[�j%jl�3z��[��m ���U���ѱ]R�w-�Gh��;��nU����N	;f�ו�����Ұ��N�{F!f�t�������S���6�U9]w�h�(w)�W���P���6��Y�%gkk��֚4Fn�eX��֘|Z�
Hw ��G(?���3��Lڡ��H�/���Imb�7i�r����xp���ZCO�m�"u�\�[��FdHN�rf�����x��D�1&'R��X����:W6��<Ps��t�)�r���RR��7m!Vn)ƕ.��ނ�.Uq������9�1�؋��3��b������Mq)ɗ��}�i�GF ����Ev�Қ�DV��G+�lժ��l�d�s�S4��Ÿ]cʎ\=b�1`�U˥&�Bh̤���RuH�ٮ���YƘ�Cjnh7�o�1��|������X��8�V��fU�*,�(ݰ���e�ur',��i��i��m����qm����f��V�+r�l>g�kFa���4�%d�Ä%��&h�=Il���Y��������7s|ͥ��j��Đx9Iֹ��4�<<�IDa�]x�^.''�]�;9���U��F��gS+Jˤ���1ˤT�,��w�|�8T˾�(r�ݣ�U�GZ���-\+:Pb�QS���Ng=Et߻c�����nn����o!�g_l�Y���n�-7�#��,;%v���vu�:��.yzC�!��a�� N��t�>���^�ˇ�(Rκv���lu��|�F�q��G�u�B�nH�*y�׶:�uL v��5�S��ug�>c(o-zo_�ˉ���n×˦���B�s��M�Sk�\)T4��wv�2=c,L:}�'�E��$3��R��xˢ��	s�f�*���𑘦�@"7i����5��j�=�Ϧ�� �f�F�m��q�He���HT{�ܣǮ����S�w[K�Q���>n�e�Ó\�[A�N�G�X�s7O!3���9C[����X�*"�B�iEX("��*,U���b�J��(�F("�,
�DUD��DU%�,H�$V*�E��E"��[ʨ�������ADdkTF~�����+����b��H��"�VL�E""�*TEATQQDQQ�6VTQ`�*�9q!��Q9m�(,�iU#iU�����
(��ʂ��rъȢ��B*�VE�b+�+���(*�*!mp���EcR6��"
��G)X��A��UR,PQE`�%�b"� ���EX�V"�Uc���A�ʂ�l`�X�S�
�#Xe(��cl�bVUEU��*�,�E��
�X*+dDlX,lT�S"2)��"�*����b���j�Ŗ�E��J#X(Tb1��&YPDV5��-ZbD�̪A���ER�AQ���JR��͵���m��>��C������y;As+��j4��ǆ>x;&e�cxn�t
GP���|�ú����;�_T�*w^���g����m��P��;r}b\��̔vƺ��*Wml��72���d���.�oE�a����ds���@��wU�(l#�울F���Σ�:1Ae]Z��I.��D4��(&�\��c�lL�0,��a![����\@Z�����`��<�l�x�YBK蓙	)'Z�t}�j�I���������8�S�EX:��h�D6}�g��h��%��Qok�M���u�y��V�FiKʑmN��+Q	2���3���s���[��6ja�汞�Un�B���/<�S�^C̣�۱�-���p�Z����ټƱ-̍b=�j�\z|�3�>@V�_yM����"lR���X|���!�ۄ��-��p��dNŊr� (��fHA���|��1�J�����]Ƶ��QѳšIc[�C��ZVx�\QçH�^n\DW�����j$#S2�U0x��:��+8b��w:�t���(���"�f�]Q�����z!^O�U�U��k��ywi�S����!%�YY�D2�j����Wj�(�^dຠ`=R�fN�x�h�7lfc,�v}�n�F-Fv�"8�u0��H��#����I�t�����auvֺ�]�A��=�4`�$%��Y���`�媟H��^-��x��$��d.�p��poKqݭX��	5�iE�gb�HU����]��N���N�(�ڌ��_�v�ߪ	��`c�"��:C��7;�~�nĹUDj�$;b�=��m�̭ã	�fI�7 LG8�,B�f���)5.�gه��x�Ե�O��l�f�r��n�-�Ű��$�q&
B	�}�Sa�E�mA]\IГ��q9�e�\�����N �f�ZsZ�FyVۨ��4k��G���`��Uo¸	59�p�l��Z�*�\D�,�j�O����ֺ���5��4&4�E�"��P�l�]7���HvN
�fn[�Dh�TK��$ĆՓC\��+\�D��XZ������Q+���j���<�R,�8WF�]~����?����6�L�����.^�ܩ�6�ڡX�2�Nx2��]�b_��p�n#2 �[�
�T���q�5ĸ	�4�6��o�֦�t\j�%��vc ��7>y��/�x�X)b^}��n���0c~�B�e9�Q���W�ʔ��|��l�Ӭ�|u�릇i�;qG֜��X�x��5�.��yv�1�q<�9�8}tqB
��B��]3>c�n~V���gb��X{6�u��h�4�@�ط�ɯ~�;����	��f�{�#�ˮx�8�I����t��;!h;"�����TD(%��"dd�j�뻆1gt�p�.����(NUY�QҎ7�GxZ��Å=/�+t�W���+�h�̓���Qr��������ŒM��"J�W�Ȕ����f9z�31FQM�R��I�fo��p��ܝ}�$Ǵj਌QYѾS
���iXy��q�Θ��1�>t�ż�c���z]]��%�D��{"�er�z�+g0s��tc��P�O��#9��l-P�,�q�7�I}q<L�[s�ܣj�a�J�D�q�n��B,3�0�S�=�_>��"�;��R��9 �	<
�'l�(H��Sg� >���t�̣��^�f��Jc�����}��ߓ�g��8
,L����� ���t-���<���Ƒ����ݙR�*T��Έ�nƐ۞0ٜ)D�6XN�2-J�5�����ƺ���u����9�2�lj�2�K�Q��Eၯ�n�,�N �r�5��~.b29����<:�K	��w2�V�ʘ�]�[�fe����FzrY��r����!/����5��=u�3�'X9ާ�\�x����-`�F���Q��S�9���Qd�͜�=C����V���(5�m��;�-f_u�Vn�wܷ�´o4ж��w)��}וN��'n�[,'�׫s�;-e+܋!W�]�E��P.���sTMkꍁ�(���<�X����\��,[��P��S�pS�q�:Q�UdW��=��ĺ�9�ro{�輞��O:�^5��/ϝ�0l5�u;<g2(L,�Eʛ�U�cz8NmՋ���^�R��&��7rۚ.o��Å�4j�:q�k�
�5Μog|Hug��/=uy�鷊���xﮡEU.�S>��yl=o�N{�G�B;�ih�#�C3�]��������V&�h228�#y�8�*��\D�z���%;Q��j�ʋ�)È�`��!�ܡ��d?LqDh=�C"�Vr�rƄ����Q�U������WSP���r��{�� }B(6�:SHV�+��
#P�v.�u(R�`�!�a������>ts���=遁����]�4�D�i}����8o�U�9��V��(+��!&/�����(�`�E��"�ӵ� �b$!&dr�Xih���w�%Y��w*���
��0p��ԫݡ+[�g1��5��|�xq�� �����r�:� \�YKK�w&�i�@���kg/{m��U<�KQ{�~v��9Ќ�OvV�\e�T�
�1ծ��sqa����ok@ڙD7�x ��zl�X���"͊S)i��-7�	.��;�+���7Pv��[4o�v�N}([�
W�z&�#�3�.6I���"ƮT���c����j�����}ўS9��8p�v]v��$*N����"gF�gd] ���cBY�=BX����$q�xd*�E���9�g���h�QJ��Y��ih�m�';�폔��y�e�pn@����\�"GnГCzS�q�e�^M��oz���3�g�w���t���eT0UIf�c�r}r��X̔w\�}�\Q[s�A��YYbȌ��[ս�8�!������ds���<dQ��3"�C7��Pɫ�[��L�����ҹ�7�Xm�"-ϔhm`&���6:ؙW���s `�!�yTE�حp�C�������-QG��Xu��>����=����w�;��o�'��xËt�{Um��#uF�ΰ��`O�����bB:L3��g��E�)yR�1����ۗZ\�wk�����5pS�:5l즪�K��PT;^y�)jj9����F�pu9�ʸ���S�"�з{Q7G��.��I�֥������-��^}�G�����a�gܞ��4V�uh����ָp����Y�//u�J�
����|ij����\�ޘFc��������߄⯷}*K�(urQ+B
J�r{z"p';S�T4ӝ��(��G�/�t
���΅�
����SzP�BlR���0a�H�٭gq��o��Q�q�=ǅ+>�ˑ.�*�>	
��^�)�%+ڒ,�=�1xfC��n�.K+[6���=[�oC���(�t�[�I�ʶ��޺�L���^ʖe=�n�d��ng�Q�Ug*a��:�M�G��:8m�������w2�h#5�B��Ov��/7�Иǽ}иǪ�b/0K�Q�)�v���A�&��M(����v1�$�jC�,��٫�]��	��@ь{6*	O���AJ���S�=��s��݉�J�������Fw>؆�B��L\?cJvd�<�1�\e�]�0Urv����3a�ډDR�"��mf��k���s��@�9�BJ0`��2N����ʜ.�j
�t�q&a��M���c|�egTG# r�"�sZ���Ϲ��t�P���:@��F
���,��Π��m�Fm]�}{Ii�]G\D�tɮt	�|r��9ֺ��l{��{��B�t��t����kO�A��r�VK���z�-���M	L��aA�Z�7���9���v���qne���Z�7_��CsFM�u�l5Y�%���J�����`2�h����z��5�ٰ8Ec�hHwM�AǺh){!���Hd�o��;y)��j����>=�P�쎮̠�������D��%�I��d�� �qq��-Dz���w��S����m��ţLT��]�����zP�	�	���$ϓU�D��S�w�*{!�{��Vc}@��T��a�W�m�Na��젬uM-��\k��iǥTlfD�t���^5�O�)Ĩ��n��a�ٍ���e�V
�I@�>'v�f�T��r�����J�HEg��~��?-,W:�J'nS�b���[�d-��k���)1���v��XNB��iҼ;�QҎ7�Gz�"J"�	�]2��w� �x��fn{f9B���8m���ʠ���%~���lB[|p(G��n�����{]�	�qq�}g�{��}���*~(,?�v�՟M�
�[B&��U�XzgLt�����O.17՛�k���� �#��U3��=qg�R�s:�F>�"]�X���h_\ۼJ�fe-���)�R�Ă��ǹ�x��mu��*E�;UN��j�6�mU��9\�F�%#�q#Z��O.�2d��^[�e�]��vCr�[�u��|�gVVM}gO<��ĳ:K/1�0���&{( LKm��\���=�Q�'��s{���p�����E��c�6��K�1Vҷ�'��e��1{'>�xi~NYA�]�	�p��!�	�z��.��t��Uk˽Qb�����7).��9T\��AӔwl�Ù����2��	��*Q8:{e�T)��.<,e>��B;aA'\a�+K��4��n�}�4e)&O-R�M�YgyԾ�	�}uՆ�HÕ�CH��d:�wQg�q8d��5�x E��߽��gg��`72x'�F7���*l��Zw<*yF�rF"�[���Gl�]E��dO��&t��Q�co6p���j龅�8�'���g�w�|��t�n
u���j}��~d���rQ2��Z�z�u�z���v%�dO�X"Ug��~�4v�����G�][E��h fi�ܫ�y=��"|Ґ���9?�uՉ�YA�*"��D1Wb������V��]�0��-����rK
o!
��D)�c����^�ק^mQ���h:Et���[1�7+��G�k4҇Q`뽡�
$��u�2US,㙫�k��|{����w�j�nWynJ��u�!Ǐ:��sCƻ4ɋHC�c�Ki-M�N��ˎ�:E���Et� ���s8�b���JZ���	�&����Z��`!CqV���2�{�0�7�\��%�����]g[��q4�9[�lE�b�Fwe̘I��������sD��6�Ī���ط�m�����dA�`�EdS��Td��	S-�:�!�)Vt9P�^]Y��k���{���X����C�>	h�i
�ѯw/�ܾv/:T)f��i�̍M��®ŧu�vM[]��Y�{�t�yx�Q:�f���cK�����|xo���/Ϫ*�4�k�3Xqt�}B}!������ـR��	%�Q��x��	O5C�.�O4:f���������<����x��"6e	ϡ�rAJ�A�B��l'�}��oLpK�$Q~�wle!Оw��3�で����1�HT�z�V#���l�'Wk�d���x�z���́Z2��\��u�0�}��Qe�4������=�\v��M>3��3���}>�_Y�ƻN�ܔ���0D��hIބ� �X1����(�w�p>�|�����H�i���.�����L=�����Ϯ���x=;�B�(�*��h�ŉ�YG}��6���ܘ-���j�`S�A�S%��"��^����z�1ּ���H��׋�AY�J���-���\���M����l�%�Q;���_]������ד����[7 ����"�L�t��ͤ�d�pwm�S\un�/�e���cyT�]��wr䉮�+E�ֺR�.KU��p�:&J<��XX�C����`E����ز��9��"+���)�����S|�����٫\��yiy�;8����>�۠��}���j�=(u�[�`s����-��}u��ш��Q�n���l�����90�-U���nU/0m셝SA=0θ��X=�(�)yR���ruu��5n�Y۳q�8�Ppl2��*:�H��22[$m;�'��s��#�$��u�72���H�s��Lv������#�)�@��k�菑#�'�o��@G�D�Ϋf����f��DO<K���K��X|�gG',�ؕ
b+�<�	
��^Ҹ�ݵ�
3+2o��x)GK�y�	��0F���!������9�H�Mˈ��p9��HD�m��uv�pc-��r��;�:q������"��0]]Q�}��y�V2|����Qק�˳R�<�Y}�C=9�`TO@F꧌.�G���Ոد���q��&c"H���r�gt�+�+8ő�I"_����jSu�鱎p��]�Ta#��ذ1۱9����0�׃ƍ�G3r(�M�`�.r���L(�R��L��3��
�*�7�6��GY ��:�6W0usY�W5�Ü�˶z�֡E>2'H�,N���Ft�6��B�$D�I��Vo�S����$3v��.�fMy��VS��,#C�A)�;��mG��P
��i�[��yj�1���u�ܙ�:aͰ�+&����a֘a�%ҽy����BW�N'��ƀ��v�a�R����4��Ǘ�#��m9+*�T��0:IM�����`���|�4v�=�(ձ����ѥY�;cQ����e_N��mpe`Yc4��!ԛUy�ٖ#�g��sz,�.(�	�R���&�
�+�S��pw���#}�%i��w="��C5*��sL��Y0ۆ��= ˚9ɪ�Me�#� 4��v�r}9[�����N��eJ�)aFQ����S���wᢤ+Um�v�v�u�ML��e�g�D)�g��6��8���%M���[îV������'U=��n1���ꀝ�	�l�ǥV�ۤ�m-��|WQ����T�k��m����6vvU�	Yx���b�}��vN�;{P�d��[}g��J�+�q� �w�L
pVv-�X/�Xn�U�Р��'d�ݬ���[KnL�{��*EC  ��l�)�,��2��\�O�N�!��Xe����J�\��r�W+\_o[i�G!�&���p�f]�1X�H�q�Lv�iM��Ю�:����Nw���:*��]��p��%DiX�C�Z���J}h�[�V�e�{��+\o;.�p��ڶ�C������A��єݳz.��҂�[��k_5[�EIU�Ъ�b�v^��Ϲz��.��%�x#[����Vk�˰�'#���j�83�бؗ ݁;�+KK��W�z&�_'�z�Ⱦ9��2�P��ѵ�Z��v��X[�����w*nX��u���*�7Zկi�0���r�b��i�S
�yη�Z�*�@�iZ�j�+f
eI� d�NW��O���,��.�����|	��3:?oU�w,V��V�u(:p�n��!9H/w\(����OJ��:�<=X���6mwl%[$�����RM�wc�n�+���#�D�hn���ӵCyY�Õ�b�������Y2ʦ�^�'X��Q���-6C��>���ťƳ�e��yҳ,�Z�p���G��[Ԃ�'_J�RK� �{�2�%�m��v
��+�H+zy����1��r$Qp�w�c��ֲYo��b��w��}�0�����oS��/��|޼`�[��"�w��}m�+U���OP�u����T;��-el�o%������d�!P_�P��n!������,å}E֊�����}�}����ڕQ�ӹ�02�ξiv�W�;������WJlV��V�+WJ������I��w��}��\�w���d��(����h�.f�̔`�UFV��EG"���UG)S1-DG�E�J5,�fac�̕DS)��X�B�
�H&S9�(���
��6�PQ\�PA"�K�X���`���k
5���s&cDd�(��C"�Vڭ��.XT-��TUQQ�T���ܥRڪ��cU"(b���)�J�!Q`�
��e�*�l�9B� ���عJ
"(-��Ea�*EPQF,dEj�,ƶʭ�QFDUEc&R�Eƈ,SV1TA�*�1U�������Ɔ%T�e�QUJ�TQ"&%�G�X����Ŋ��#&5[V()"���c9J1ƙK#"��1I1��TV�FJ�T�
���fZ�\����
��*A11đkDPPR"��1�PU�m�[�lY2�H�1�kPģ�[k��}�qt49n[�ΏiB8����O�:�U��.��z�	`+qV��7�v�-*V��$�^	ʇuj#�T�3+*4DE��I.�SYh���a&:)1$� ����5�bEf���)x#�g��5o{���"y�]�=��*�Mk��tP�J$�J��vL" ������`�v�����C��]2�t����@�h��Nk\�*�u����(`g���_�(��mf>�>S�öH�yXB5��WQ~���7L��@�N�9`��Z�nTن�\l����kTr��-�|)�(�ě#^]�~3pn��;T��,�LHmY:���."u]�=��y��.C�t�6��E�/�N�"��C#�Pʺ
�鏶,gO��oW�l9D��R�U�=L�͆�mjڵ�Cj�����㓆�%N8�G"6��oh+SK`q��k�h�6j���sH�s�d�qn�什����b���`O��F�X+��a��/� �V���'g��aJ�:wˣrUȅ2��Ek���<g`#d!�*�F@�TD(%�T��F\�r]��/;�o:�*	ce�\�r�bT�<�^p�V7�G�*"��
zYX�W��_�]8fdѽ(�̏Y���t���vW��9r�齘��1��a���C��<�R|�K����B��V�\�r-���A�����	�u�\��;u,ӈ�̀�t�G�/y�^iI��r�V� 2;�Ž����[rT:!jo��l1Q����<k�ʉ��PDRT�!u�����zaS�f;�s(�Rh��'wJٷU�1Ktc�to� ��Y���T(~[BRiXa��񸷂������t�e���L�bYf":#����CJET�s��Ş�gq��S�^����u����5#������D�ͭ�۰s�u��ܞ� _�C��t>�8�y�z��0�+c�Mʦ9$�f�i�����")�]��R���H!тzA��M�DW�B�.u�Q{;B��61���j�Y�9\��AӍ�3�����Q~nn!� ��������Ut��a��Pnr =��DRN�����sF�n�*rW榴��I{��o�f��eC�$[Ok�sO?�q��r��2+�̅C�n�,�N ����5��s�x^4N�Pȍ�Cu��S��~�^;
�vl�b�x׼pJ�Uaق��zFen.��ez$z�!��ښ�7Uu��q���-i+�A<l���}�;^�s�r���r���j�a�J��Ư�$GVE�Vo�W޷�@��g.e�eYTgE�뻘��Z�	YKø��*��nnT�V[��[5��*Z��
i[ֺ��U��4˧��@:��V��eЉ>W(h.�>,]���o7P�~���S#��gR�� �fT4��M�(��P�^LL.�GQ���G��T�r�ܷ�ȍ0�,�<�fE���fQ��2,��.s�招��a�3׉�7Έ�=��b��sq�9o�T�I~��w��{.j��}Zla�5��rUW��w�ѭ�aǛTuGb6�cH�4�����|��EiI��"\i�Q��_��
$��q�J�e�s4F_5��]��1xXq���o����6w]�Q�b�K�]��u����:� �%,�	����z)l_N�2�2=�[;*���Q�r̘�T����T�k�`4��"M�w��P��傭;Jc
V
�KQW-�̹�Wb8N�x��6��|��4��'����r�:zR�p�.!�ip�Xl�����(�G^	�E��j:/�fJ�B�	3�r�^J�y�AMe����=�g���'К��x�C���px��6gjQ������R�z2�4D��C�@�sVㆢ��{Aˑ^߲��������ΆYl�v]v�7�FCvɧ�f�����Owv��B�����JQ�8p_L�[F"_6��<�JY����B�I�%��7Gz�5��)���w��ک�k�]P�%T��{6���\��ylra̼�������H��q�W8����n,'+�"���T�\�{�}��	R{hM	��^\�8ȼ2oP}�R�!��9�dVF��n\5�}���z�d����y+}�T늘]t�N/z`����T�w���ܱV�8�y�d�K��ϟe^��45�d�:��:fd��I���|s��":ӧ�w�*�)���受��R���GTyL0��h4��W5q��8D�u%�"���3"J�g�c�d%hm��G�I��W�|���D��>Q��׹��&�ζ&U�GQ����F��U����ii����E���3�Ή���~��"�������d�^���g*rOy�X�â�����n/���{tER4va����ec�mK��SK3�+�qy�NsU�,��&Pţ�V�� >�(�['iި���ƀ1��?=I�x��Z���V�9�Cx,����V�י� +]Z��oJ�����u���u���ZJ,©��Js��aJ7��NY�b����T���!�̾���������B�#)l�;"�Av�!WB*���Ĵ5,�\�Yh�b�]%O'z�b�8�N�(�|�Ӕ�B���1,�ϧ�Zƍ��i|������B��wy���е����-s �V�2���\��,7���`$L����4�7"|�Y��C��o�'��n*Z�^�qGӤq�ܸ��T��#:����.rs87����3e�L;�E�{$X�*�.�(��L��=�'�.�F`�wSy�N�r��oB��2F��p����k�&j���J8_�� �p>=�dՇ}��8�u}	�U��Dc�GW�����cy̒yt���JUwFB�u�������4mq.8�iv'�ꑼ���ķN�l�
7͉%�2H�BB���*4:��u;ǯ��)����^9��J3�DR����u5�:(I�yD�)XI�Qh�˚p~S�932�6Ky��6Ñ�h4�yā>�����
��B�����V�=��r����"1�X�^�DH��:�p�/���8��'��2y�'��9(M��5(�<�Ѽ5'��L]�5����t]��<+���n����zA[��t��I�mY5�A�D�����w�9S�;"}�s��Á��Z�s��L�:c9�"��Y⽕t�L}�c:~3�g��6���s�I=W	� R�*úK�]��ҹ^���bX���,���|��C���*�����B�H;cH�zm{z��'y�:���;���@p*�Hs�=5Ϝ8Z��;������ӓa�w Gf�D\� Y�3u9{},�
�Y&����x!2�dGb��ؔ�$��aԃ;A;@��r�G�&�Q�{t֟a�Ե��i���u�1I�K�*.�4�[�Vl�s!;��C����T�|�N̔M�{��Mr�l�5�o��C
f�H�J�\�C�e��y�Ns�v6BӲ.��g`uӪ"ݡ�[����x;d�{�ZMs
���KPM{��p!Cp�t��t�c��-P��D�E��Z�!���t�^n�x�������2��3�+�̖j�Q5���J�W�Ȕ���
�(YGnzF�R]��W�j��36@�'�kev��/�q��\]��g�.�Cý&�&pj���fֲ�8�;��s;��Ft�\��D*��>08�!�"��2Ob ���>��{k� %��`���=�=]ӐC=�W�����C���D�2��h�8�}�6�������3�ys#V�k7ۺ5v� _�N���,��uڀ����C���YЍ�D�>�%�����-����:��ϱt��=�9\�p޷vϬ9�p,)�R����Cxd�U��Q����B�Ќ�iT8� 3/�ݭ��1
K��@�*c�_�K����i畭]Y��\����5�1��$�ge[�Z��`��R�\�w�܎�^j�k�ُ:�RV��f0{v����69�r���\T���/�4,O4�m�8�܆u�i��C�S�&X�cȅ��>�u�P��dRN����ۚ0p�N��*}�_���
�]Z䤃o��`x��,s�n�}MV�wp��5ٹ�3g�q��I�sF��·��꘎��x���"�9��\u�͚���pT�orF"�T7]�E��P.��܈
�l)�ʫe����ӢS錃�C8`�u!���H�;��)N8���n�b��^�	���� ��-������,{ډ�(��P����]���vm��Qr��㱘�yֺxLT�W��z%3{K�/kv0rJ���]�W�yQsc���,٣V9Ѓ�_P�����˘�YX�0Ŧ�z�I�/#��\��o���`���w��c[�Ӛ���g��ڧO��&ͽA����w�37Y��ڌ3�U��@�D�ι�*��q���e���ӷl7�k��Ľ�=w�w9��X\|yX�A-����謊qYʁ��C1A*e���x*�t��k��7q��!2�c���Q^��/���-����r���S}*������6o�����JL���i��Y�;��/��/S���1����.oe��2���Z�O�h�/zL���ث!a����C���d�%d:�wq����5�VV$M�Z�U��^v�V1M������|���Ja�"�c��dA���u=��u�`�W��R�H�9Vi���:g��I�t
Oiw�盫�C��ù�=0�=C� l�"��.�p��q	�G=;Q�al�)_�B�	$!F&wE��m(Zu�GqR�`��F�g�:5���a���{��� �ԣa9�8�[�
Yk�Iݜ�{so}�L�P�&*����-��s���3��0��ݻ�a�]���Y<w:�n�tt5в6	�}���zA{Bjg�K�$q�xd-���K臞qCT�^�qu筼.du�MpT�}纠^�D��K|g�k�ʕѦ�%8ވ#GnГ��Fwd�m>ƛլ'ONQk�)�ʈ�~s,ё� �'\�u32Q��5����η|�*����<���kM4�(��9���Ҋ\���	���inPT�*�v},�f�̹Ơ�Bl������3Fߪkif�,��㚝"��F��k�;by�D��`Y�%1�MJ�N�iLmިp.��������+jB5�%�_���]I�p���k/n(N[q6s2�p9S3Q�}x�=o��#mq����:���;b����*��8�w�5!���G/7.��ٔ2���Pe'&i5�\��@���z��Y|;f�X7ǭb�-\Pdo&��A+�wɸkqTޱlr2�m�u3�I�{�e+U݋gI�2�M�޷���F,a��;��_u=��R*�:���g��eR藂1�U���)��T�Xi]�Sy`8g�{Y-*��vSU^�^�@ϊ�#iި���ə��5�{Z��|�l)�YU�n���+��0S���j�a�|���
���}�s}�����e��վ펞�gH��8%���:99dNŊR���W�ə}
�����q.��&��I.G�_#I�`CqBZ�XJt�0�Z��
�Ѣ#%��혭Ҹ$�����A���44?��0桶�V�#�]Q�}�����B!��Q5�S�9�y��mF�u�t"�Kqu�33�L���w���yv�Xl����s�!G^r[��f���DsrI!L�
T;�v��]7�s�R�]т�b}䕕:�[KR�����}	~���X{a$X��L�BIJ�2H�Gdx����X./��3�4ym^�Q��OzJ�;��"a�ڋ۱���k\�$���@������L$9�a۵k���ME�r�Z��-T�L\.?�<�赒��|Ս_wf:��W�f�U�e����7|2�'K"Gd�Ѽ)	V"C6�
/�-b��%��ތ9�k�U���uZ˖{;vʗX%���P��kn����T�l�j!��e+��f��,�\���5D���CAā#�418�p#��m�XU50�bN�683�^�8�⫮��9qf��y\C5��t"�&�tɮt	��_�n{_�<d����fs��<XS��t�X��| h�3�tW;���k��= ��$�@K(��Փ��]�Gջ����s��l����e��#��>�9�j�����q�J?���^��+���ݴo(�jd�FU��p�oeB�=����".�΁��*VR�~;5����b���@���#���j��ԒGc��0�r����Vl�v��s�~>�F�X+��@��|�N���{d;S�p"�+]����dHٞޑ2���e��y�Ns�v,��*;"�����g	괐c�&�=x��Q�XMf��ܓ��W9<��P9��R�<����Ⴥ���͜���W�^��/d��#R.Lb�*!VL�k�ʉ�g*�"�T�B��6!-�:hOY�����_�L-���Lk�f+�Q���V����7P�.σ��<iv*>2����K�����p�V��b�Z�h���f� x<TG�t�A��[i��9b�E�tA)��s�ni���<n��!L�5𮬹��V�J����z�:9�	� �Ș��1Vժ�v��k�TQ��V����Z���+�K�{�;���]�MݷZ2����0'ڶ�݌	I�8��ri�+�a"��Y���1=��.gU*���w���m�ԗ���zC��Bp���eA�|llj�1!8�Vl��q�g{Rc7���x�o���G��].���umj�ٖ��[�:+�k�#PPb�gW:�����ͻ,��k��y���GŜ޼�tض�E�l�H׋#������y|�����W^N��"�{r�+�F�Tȳ�;dc�wIԭ�t�r}D1u�!����vns��ˍ�j�Վ�K�5��&��UֱDrN5�rl�b
�G`�o��`x����Z�� �ή���ʮ�6�mGc��K�uAqK{;����\Jx�Se`��t#� jJ9����԰T�_,��*���[S�	�O������LSr1�k�D�}1���A�Y��r�����l�tE����vn��Wy1���v��ҏ+&�<���<��m�5��!Y��3y�X����  ��n�mamL��[q��w�pO�˧&�ʹf�׉L��>���͸S=��F7e� Zϯz�J��+����q�k2L�Ԧb�i%�(w^ 4b��
Lvr�)j"<èi趢���3��W]`��J��d�����0�x�:꼾��P�@�3��ն륅�E���ZEX6l+�q�-th]�P��p�,�H�\�m��&W	ٙQP9YVXF�ٵƛ"'S6�N��-l�ʥz'+�%���R����ţ�ݸK���Lt�`�X��7,ή����R��R=� �)Ǥ�2^�ڇ~(�j��ϓa�2s�2_%N��/sE"%����3WC��,�$Jv[F�hU7���ĳy���]��oS��ݺ�I_gN��\PY�R��J��>�,V�*smh�g'$]_ub����p�ܛj��e^9�3�`���:K��1��7t�f$K{t�vTܸ��ҭ�Z(s���Q��yd7�ܴ��;;(Zux��:R��x��G����2�m(Z;d���Z�n.��3�u��Qa� ��
���.}U��};;5A�S^2U�w�F�QDo����n�(P//�m�2+��� U�|V7��Z xW:�sk��&��4�Q��.g6���h�]�ZZ�쎑���Q�yk~.��U �V�_X�:SyA���g����/��5:&o
�2�{
/k�G:)9fY�F=��`瓣�Sc��ۓ��͝v7��7E�,0��o;k�Q��Y�����ٰ1о���Ӷ��J��jƎn *�;[�R]e�r�o!�d&y�g!R�%�7-�F�r�g�l�S�F�ⲅ�Z9QV���Y��(�}}U�fg�,JB�&$��z" A�>��MZ�L���H,�T(#R(*�UTEdbG(ElR*���Ua�ȱEE@DƢ"Ȋ�I�3�m& `*,D�ŶEEEDq���T�m�J��`�V*��*����%�f`c�
�X�bEE��U����1��-b��"* .$�*��*"0m�����Tb1b,�"�Y�
�DDDA"�"���������A��`(�R#�TTX���H�"�Z��-��F*�RҪ�mb�X��,�&[
�X�b*DQEb�B�PF1X��
�@QUAUB((

"��DQb1kEV*��b��y��J���ݧ��_R�'h��:@��s��+rbu���{u��m�ʉj�+�/E�*���֯Fs�������)��}k���;��;�b�� v��&A����3��=qg�	J��%M߲7n�4�mj��Gvn`���i�ۇ�G<2JV"x� ��4{�Q�(�u{���QY��{K-��o
���"5Ɲ�7CM�dC��P��R���:�zL,�TV���s5�a����"�M�9��8�S��'�n�8�p4)�R����Cc�������?y���������,lQ��^�
�#�BNx�N+Kq&�N�2Gl�=�[�.�����W��y�y_ı�v��h�q�
w૞�H�;Ď��VL3�٨��2�p�����`��dj�掿����K���k�pO��XY���;���I5I�St��i��z�ʆ�0D���}1�K6`��t`;^�w�|��oW~�"��L��<���[�ʳC�#vj�-�tKr�3�j�65�D��p#��dP!�OzB���͵�YW�Ni��7F�W��\Q���a�wH|�\Ir�7���͚5`s�F:��tEs�8M^�����h�eN�(��=�o���\�E��C���9SPs��	./b�Yհ���v���Zr��Lpfk潫Y�H�����ܻFU���>lu��_[�\en���e*Z�\(�v�����tk9�t[�Ȍ3���늟�n>�2Vq����g��c�\^��5��nUW��^{���z��lEZ�1#\�n�ǝ�6v!�E��ugb�/�h g!g�ι�*��\D�z9p����xܮ�ʳ���ӭ�ܷZeE9fg��0E��ȧ��@��D3�վ���LOS@�<K����SG0Z���娣t�0Q�3<U�S$q�S�E�F[�w���'�Sb@�;�^A:K葏�҅,�F�������-�؎����I��4���&���/���_3�|����[^��yE���=�uC��8��}A�~zv��������k�_��s�u9��ڗw��~��l�E1�۞��{�:���[4lڔl'>��,�=��w6V��AT�hq_�A�U�ң��U���ֿM�|��3��ӆ��txT�`�"���7ڕ꺴��c ���z��'���4&yt���#��
��>��/�%B{�}��X�S��Y���X�A]������8,��Dyr ϶|T늿
�ѧn��_ND�gsf�LmDR��H���zx�g{+M�m3C;�.��g�8�+,)6�.��ƿZ� �l�����s����w�<\�b�F��ݙ�w"�ÕaYPZ�݋��kl�[����ԝ)V`疠x����0�ӵ	M|��F��Yt��T
����<�X4F��s$a5ΰ��URY�&=��'С�:U�ѓӽ�z�;f��v�� %J⍭�9��`�iC��}��9X�o�C�t1F�ݴ<�%��M*��iYQ�
���ca���f���S�DW�ה6�����r&T�5���cL��v�����T�"�!�FVP�0Ή/"���=�wG�BڿpvS��dX�8�5r���2�ځ7\p"͊�R��:�m� b�PW�4�L3�(����Jw�-�q�o{.;�0�4-�eH��鍁ڈ�gGuSV�Ϛ�������v/Tw3�i�;<r�e���صp��8��#�۱�-���S�
�`Y�caeK�,�oe�D����~�SǼ���=��hB+���Tۜ����oE�,�غR�"�R/�A�����9"Í��*��L��h��f�>��_l�.9Ǩ_#I�c��P����\Q�t�[�s\���2�rxbi�J���P�Ό�$�w_ѡ��*bif�#��:8E���j��M3X�W}�qըȘ�+�>���M��X��rH�l��v):�r��s�M�F���Q�#��|P%�����=+�mi��.���u��^XF�X�EWr���%Vf�Yb-�収Q��Tz:���o�Yar�Vv}q�9x�P�H���Q���EX���Iq�ˑ+�9���"Go�@p�uD�ت�5�]B��Jqݠ5b69�V�n�U�5-��W_`�ÆiE��;�c�I��
��o9�O.��9�()U�9U��D��;(ri(��7a�;�x�ؗ*��
0�
)�$�fIB�F��bBŽYV�����˪�Q�6���a��^s6��v�s��p9ΊQ�-2NɄD�P�p5�wSu�g�K�L�͘/�b�($�yā>ѡ�sZ�F*�u
a#]��;��+Oucu�K=�����G��A��nQ��n߅p������ħ�L��} k���4VC��壷�<Ը���ͥ��,H}L�W���n�M�U����RK�%�I��3�u3SMg�Բ���A�<��D�����`����x1b����.�uҏ�aC�{�m���C��wҢ[i-��E�uL�j	К�"/���.;�'(�0����T��j�)2ǔV;/f��:S�խ=�R�q�\Ӂo]Y��n��i��m�k�r��\ҁ��`aݾ%�sw�/s��-Y�rQ����:��d���|��i�4��k)m����'K{.��
G�-.��y�{F��~^�E�kG�/s�;�ç�1��"��Aj�G�Z�g\��>p��:��n�|6�n)���uX�lr��LU�V��/�,n��h��'���S�`s짓w�Ώ8_kw�k�3�e!Q�x�m��rr�:�}�ląybv�'FO(&�)�X��nJ��y�:Q�����Kw)"�M�}���ܤ�)�es����>g�W;HxM�^��"�T��ȸ95� @j�7:u8Ior�՘[�za]�f`B X7�TN����7
��σo3Ɛཾ��\��EP��[Աu@������!�'��' �W��6��n�c���3{E��p��6Ӡ�tc�$;�V�LtA%+<L�	��O���&
�j�d.��s������^�n�GDF�Ӹ�5�rȊ�P3��qx�$��"��u��5�n0o}fz	q��T�"Ϟ>��� S������g��8�8*T=C��
�t�۲��6�llFp�z��@�/`H!=YGl2($�<qZ]������i���38�������ϞZCgM��2��E�����r�]E{��v��E�x�B�ܦc*!�<���	��ºh��bo��x�)��@�l_f���.n���E�{|��\+�����N]����3�׽t��>���݊��q�7����nM���t��Y��V|��g��C���x��I�Jr��#�£��(�e۝�m����P�&�u�9���q�b�	[Zw*S�;p,�Ȳǝ!�͏9R����>�qWP�NP.����Q:�c �p���>�v�>�;��=Jq�&�P+g��t�V���;g���ګ"��!l�S���y� �[FŪ~z0V�~"��ą���ׯ�#z8�l�g6+Ե@nU��'6����C�85�8݋<<�f��"v۷�/e��Μ��i��{�������a�w�� ��Io\���y��=�7פ����%X{�Vo8�[���r#�"��G�0��
����D�ι�)�Y7˕9J��wO4��b�Օ$[��ؕmF�ZeE�
p�3�A�<@�Fq�ʁ*v��9��C`gMu7��J.��E(��l�e'zo���%?/�����搭`4���4Χ��ۚ�T,׽"�?k�x�K5��!�a犑��lGE�."	<M�Ќf�/�m;+�&"���dvC�L�����>�yśqUǳ�uC�7��R}A�a�ڎ�[0
R�����tSLP��$�Y��X���:���.{3u�W(ks��1A����]b5�S�z�M���w�K��[��[���u��5϶soKy��79-��k�8Q�\�r�f�G�V�%m������ ��O�].̨��ĎmN�����W
n�b���Y�����b�Oe����g��y{���3�(��wL��茜����Zw�qj+L�{$�БV߲����M�8ޟ
�xw��mm���(֖�V�n��8c ��'^��{<V:N����
�,��^�ZX�7�`U�qj����s��9�guX�FI.����$#�c��R�4��q�M��c\}��/Pͫ�O����Iz帇�X4�46Ù#	�u��_UT�}�k>P]it�����PΩ��G�K;cz���T�(���ܰi�"��8hO�X�7�!���k���B�n������u��&���<&��N����jtH��^QM�׽��K��=��{���^4����j
�f�媺�Лv�|_��pzP��[�`��wG�rWVo�xL8�v�UOq��>o�s!w�`�c�A�(��F��6�yo�,����\��-)5�Z$=�p�{]@��WmT�,=����F��j��lu	^�m��K�o�YI�`��xu�\6������[t�G7�սL�8+4����Kã���e����ʧw}�=K	�r�:�p�Rh��8�䚰��ܦ���V��=��+�ň
z�<aC���s�����Ŭ��㭸�fwc�5�T��c��yN�oWR�r>fm���'�U���3���u�B͸��B��³̓*]G���BSR��.fҽʂG>�d���|�OR���XE��z-9dK���o��T�:u�{N�I��P�1J��[ق3���/���9�	j�a)ҊN�Ǡc<Ԯ�������b�ވ�nGq�[Q!�2�Yu'�{�7�z�ol�EtqF{�r�p���o��[����=�<��Ϣ��	F��Tn�xԮ�f��)�q��:fV��-�b�-]�B2)Q�*L��;�D����A�s$�[+��u��o0��k�ޒX)�c����w�۱6�]�~Q��QM�%�2H�@��5�����5�f���˄[]����&�N�X��3~s6��v�s��Ʒ�)��wQ=.)��zг����*CпU�'6
�5=�S)�e�N�!�y�C-9�p#<�m�r��4�?j˖s��<���h��H4w�/�d,��B=�5Q�-�d�:�8��ӖU��(-��d4WP�
��}�{��ϱ3{ȭ�u5�T��6�S�f���T�����1t6�CS�'N�^B� ^���i� &Κ�B'�;g�+���;9%d\����p�6����IS/��9�j�61�|��T[y��1�󶮉.p���ڬs���皔��>��=4p]��
���f���􂧻U��/�#�Ӌ�g����~;&����+\�D��]aj0GO}:sEH�0��5!/5U}��nD�u�t&��&��@�~�U��)��"ƺ-?���������\,�)`;���8��[��&���A��ݧi��sc���5�8\���n��`';1���gHJjQ��6f�[��2m%���OFD'Ᲊ��4��̽R3��K��(�C[�:s�\�!�o�^a̹�ɖ�z����ѨD(�uQ.I}~�D�<���#��-���^p�kD��~�(���3��g�����[��ra�p�B*2Y�/�^�UBRf���P������ݍ׺��|���p��xj='��,.J��\�[�2�{�#8j��ɋ��ksި
��=~\�E�@���C�m+ -V����Q��@L�3���ґ1�pH�[����wt��{+�{zst�����Z}v�<�c��%+<L�`�û�X�9N��Ƃ[��jW��I��ɍg
���8��*[)�l�jё�3-�8Y�,��E���j\iV!�T������ᘶ���*c��Ή�|W	gj�n��!�:Ma�p\]����� H���l�쩴��Tq4�L��7�6�;M��	V�}"�!��0M3U������~����w�nYN��@�'¥ŌrAD)˸��!՘���o��̒P5�K�H�T��J�}p)��b�n��8�py��q�̼{0�B��3p���s�d"4��OJ"�@N��"=��Г�0��ix��o�ݒ�ol�e�hq�*�0x��C��3���:���8"(�x��j�Gʐ����T3*��vF������=%��7Q�҉4F�ߋD����ɝ�v<t�x��e�+F�b���e�k7�����t{�e�,8<�C_Tl�p���>õ��r0�ެ�ȔiK{�yI�Ӎ�ӂ�X��Uv���~f_��xP��J�D�c"�3GD�/:�n.V951�ܡ��Q�X��fJ/��qF�U7��!������l6h�t)���g+'q�c�ܺ�?t �2�*7�3�HY�^��+[{��sg�ޟz	UQﳵJ��"|�h�<�o�;7�׍���r���`�1����m8n��y��{��	!I��$�	'��$�	'�`IKH@�xB��$ I?���$��$�	%��$�	'���$���$ I?�	!I�B���$��B����$����$��$�	'��$ I?�	!I� IO�$�	'��PVI��n�Q��w��X���y�d�������}
(@	�
((���J@(�
P	�(� P)J�*�� %
J ��ݝP(��P�!J��%%UTR�"Q
")$�*��*)	*(��%UR%TBT�"UT����{�)
T��D�(UP��R��B%()	 ��*���D R"�J$"�R������B������HU   ��km%��%��ֵ�J�4deTl���	V`[Dْ�0 ,�R��Y�bR�ȉ U�  ws �� ؓ
�m�UUJ�j��%RULa�Ѷ͔%lm�kl�(�b�!�
 $UQ� A�40����%+`)����&��ʦ�(�0[`�TcZ��Z����l�A�*�R�*�l�T�QC� rJ�	�hPLfV��
(��QJ(8�
(���pB�
 �B�u[�( (P�Сn�� �B�(�A�;� B�w6b�R�% � :�j��Ъ�+[l5`���U3l�#-�իZZ�,k4EF�j�&մf���f+@�5��[[CZ%��Km��F�I�ShUE$�B�T�\  jv��kU��L��Zʚ���3ke��Kj-UR���m2���d�h�m��)C5�m[F�&�&�-��*m�V�X��PJ�*$U"m�   6�Z[J�5�kI�V�E*��IVmkeU��5�Z��cl�(m�����[Mjd�M�h
�J��)Zچͱ��B(��@�U@   'S
U�S&�U6M�i�!��MV͢iUk1���Z5�h�-[U5�UI@�L�55���J�T5kV�J%T��")T �\   �UڭeR������R`�Zֱ��[,XQ��Z���#V�LMPMTDֶ��ll֪�Vj�X%b��5�m6�DPmP�D8   ��J���`Z�͛B�ڦ��`ʡ�����U���L�2���نi�Z��K[Y�Tаj����m.�*�D51�ʔ�� ��COhaJR��M� i��4�U?Pؠ��      O��J�� i���M�iO	����& =OA�	4�T�L'�i����&��C@ee�fbP�o��&V�IBJ�i+J_J11:U]�U:�J ��]�?j��EG�p2�@PMb�����ADTf�K����#�D�����"M BB%C�$�@��Ԓ�i
�l
*5�nʽ�R�A�����j"� Y]��I2��I������s��*��BL�4*�,�a�0�3LQaأ��А�s*�4.\�
K@�1r!]D՜U��c6�}�Yb�,�se ���8na��)F���0Z���� B��W��j+Z�'{h���G���˻��2��e�ӧ��$M��T� �*�0�ҽ6̻8���-��5��e*Vj��b��u
XHzӔ̀*�
����d����y���@�4�bV��wN�x6S��ĩ
j[�BVVn��"��M�7��q���R�\�f�{q��;Ve(�gm�l�72��Tڴ�yt�E*�ik/&�9&��S��	Z��;��j�n�v��9wtsm�4[�!W��-sE'TV n�]�>N�W�3
�N��C)��u�� Әkd ����ᮣ�b�A�$w[5a�껣u6�Z�ef�@�+(��[V�f	GjУ#�Ӧ�+�[f�����6Gn]�7KLJ(���Ip�Z'	����\j�QQi���s�ʻf�k���H:6���W�7i5�muhe:�ܻPW���ӥ�����j�u�h9���sCs��VO�0m��Ukh9t����c$fc��`Yz��VP�R�]X`a�%J�S3u:��3d�"�[��� ��L�i�2��yr�VmK
�aY�ꜻ2h�Z�jզ�)@���ol����ئ����t�!f�L��J�3%�sN�4� r} �t�m��F�K&�ۤ!�E��ԥ�5��&���Lm1d���*�j��){ZA}��nօ��+��9��4V��-5eo:y��K�<g�v���Xy^f�@�Z�U���JV����f]f��gCߊX1�֠�+$�h�O�m��n1̔��r�x��R��Cl;[G1ڀcPM�L+e��ڒ�WkD���y�m�`=�N]cv���uc�D$���`[f�>��8j�3����<CU�qM
-����Հ�P&���>XDT�^2���%4�YUN����7�\���Bf��X?nIE�5|�̫9�(�h��� �؃���ũ{���xu��)Q�:�K��"���(�A�����.�G6�sl��*	.ˣnLQ��S���*��*�(� hȰ�wWH0����7�/(����$ƶ0L�n�K6�7�� vj���`5ݱ�>u��> ^[包O5S��s.�S]�+������"ۄm��sp:�u��ܹ��H�Ω�m�I�b��f�M.�iG4%hV�a���ɷ��v�m�J�b�z�]�4�[J�[[ՙM�HY�&Ô�V��jcA�Y��d̲�وenY�βq,��?��n尝�t2��%�²�іū���J�Z�6�QHv��hj��62��fJB1J���%�e��#. Bx��E���cݴŬ#3�OU�K�) ��j���WCvZ�"4Q,K�(�KݔpF�˷G���Q�i��6�%�0�۱@|�]��xnP�;:ޑ1^�v���kڃ�|���w�9�.�=X�6)�Z��8�i��Ӡ���m�Zpi�Y�dz����-���b�*�T̢�+���XH^ϭ$�jnhڙ�4�0�k�AJ�&�i��6��G�б���;V�r�Rgq�6�`�`� X�B�d�Y���q�VD�����sh���|�Ou��GB�Y�|mh �jU�F�͂+&�I˚��W_j
�������N�j��w��kn0�Ԕ�ѧvU���kͩ�X�S[Z��豩@��+kwִ���ч2EU��lwvF��(����,୽@���Ցr�(l��8m�r�U�Xz�^nk,RGe�,aF���F"��ۄ���W��^�v�꼬�t��38b�`����w�J�g����n%ݐk��_glլ:j٨Pٗ�r��5kk�,���OΒ��G��Ye�+6���t)`XOR��i�ъ��sӃ�{ɲ��:9s�A��6�AZ�d�t�^ғiÛ� n���dQ���J��|Ef�kS�uD��UjT��qQwjf�ת��k\�	��Xyy�]�x�d��`cp'�1�=���GS��[3B�ܽ��p��9� �3wy���N���I���gF��ŗ�r��� 2+SU�[�S�t���  K�J�Tʵ��Y������x��_���B�wi+*;vB��jހ�VY�W��#����Z�MDTt�2�,�VL�aFF��
*���5�|�+Z��l�;ê���ލua��
Dv�lb��=�f��I�eL�̬E�D6��0�L�����["��jN����:kd4M�u2�ob�"�71�-<�BÓ
XF݂�
n�\���2LLaj��5�4�ǏƬ[�ǌ\sT�����7/L3Qź靡6#��ޙ/�Lҏ6M�*+�e"�5o^$
���]��+-�C(=[�T�U���=�0曼u	f��B�s���w�Gf0�1m��ž�f��M,��k��fV]j߮��3A .�F� �%n��7��*U�+#�ڃ���)�w��R��Br��d,��+�3fփ�̵��S0SZ�Z�*�����9xL�LHP.�Z>��Kw�������[�!�T�-��kA�K7-ܺ��!�e�nZ��[t�$V�*᡹�RRd�E�ʇsE��+��	���e�-X.�m��-Z��ո�z�u��_Z�X��\9��ϷYu�z��{�oM�K�n�E5�9�������6MѪ�fXS���u�2SH֜�sף�7X����Q[��E���R���H�.�ϯn���팺�+u��2
�b��QQ�.�RY��X3° �A��l�"�P5v�a��Ḛ;�]�*�OŅ;*�x�Y��Q�r���n�[�yR�i�Mr�dv#�Vf��������cH��_b�[�I�^��g|>��Xi���2�-ݶ�&f�3k(RyX&�U$���ࡸ�(�2�3EI����WIكY���Hц2F���ޤU�^�
��bQ:�M�r�Z�m����l�*@�ou1�V�-a�x7om�
�̢r��fYg]X(���n�hK��2e\�.t�'(>#�S��Y��v�B�,	�R�*Ouwc�`W�ea�j���Vv5Ƕ�0��W*vF�stݣE:5����I��I��ЮЅnf*�:i�W�.�ٵ����+͂�LX ��,�
���x�Y��`�Z�֒�Zi��G9�^�$F�����&�̈́�1�V�q�,%�m7F-��
#:�-��h���VN���&�
��36�Z@Y[�ͬ�A+cs~6��C6Q&����f��v��E�8�(*@�1\)\x�˥�|+r�nm+�l��M���M��Q9��f,X��G{kM,�=���w��)�[���G�6(́Z6��Ġ����tk-	p��4��
@*�]V��K���i6� �{�'l�Wsa
Gt�<@�1cv�͉+���i�b��հj5 ^]-��L��`V+�d�B�ܼ��6ҹ�q����m\�v�+SRѳsX��5{[b�Γ%�-�A���q��W7+	�Y�02�*f�eY{��.��r�@V@B 0^�J��+i�5t0�[&����ڣ�V+���$��mo>o��:~̏t�&mab:ڕ�\R�}�ߚW���.�а��r�cN�b�i���}�wj`h��B��QB9���ȡ�/,T�6�[�ݡ�fa�Z^��i��Y(t�1[�F�<���U�t�nAIw���e�kN7!qؚ���ͥN#�{2mL�	b�̾��|q*	-�4j�_Q.��s��ݙ�%�<�)��_\�> �lW�:�6塒�.��2[-b����i�x��d=g^5u�[��7�=�ko o�)�Z[�e�h�Bb��V-,ш�Շ����⭧��C/M["����KH�6�̀eH۽�g6���U����%.���H�l�r�L�M�m�Y84��֑Gp�Q��ib+��c4we��*43ql�[1K�V
�F��	T)+NT�T�2=S�9�_&4��Bc�Ѝ�h����@@��9����/F����*ʳhY�R! ��e��!k��[�B�"�J:�g��dZr��VU_tǆ���j���R�[�W|��6*��f��c�2@UEf�n�T
5˞��4>�Υ�ݬ�;(���[��^ػ�̴���8^ڼ����C���\��ˮw�c�f�Tȱcwo�j�B,�▅��*�8#�ݵT4;�e��lU�����K77ڗ�Z���!��"v�0�������T�*N�v����
�ی#0�0�A��ƍ�p[�(V��H�rM�VR��%�LDB��e��n� ���J�^�1���t=
x�;jf(�%�+wu^ٸL��S"� �j�]��mJ�׺q��yG3.'[�1�cВ* w٧S�:F�d5��v�M�j�&�ò�%[�*fDBwSF^0�,�8��z��	���Ŋ��I�&bծ�c�R��݂_�IT�<����˃fAC3.��'�k�mâ�PY���:3���/n��TFv&�j@�C�75Ga*�ʶ��u�,��o/f�t͈^���j�L��`�lJ�]��KcUӇ.�>*V ԠP��#x���RWtc5�lY���)IY*��O7��1R6૎K�"��wY�/w*q���l��Q��5��;G(iz͗o]�gp�Cm��D����vVv�<�>ܥ�Yl��A�J��8f�ũn�dn�O�M�%*mm�J�˺��sj)�;{��KB�0��t-�a^cۛX6��0���Yʺ�^;Ŧ���vJ�ݘsve1�����Үݔ�wi!����p�84��6��:��@������
��a�D��fi�-�@J�#{sV�ͥA�5y�30P�	�N�)Rc�� ���Wz���S��b�Ik�ʲ]��N%yVSSf4�ɺT��(���2�A��ۨ�HJ�.�64�t��(a鈥j.�A+�ٱ�@yqi�R�r�Y@e]7��i[ty=!X8�L4RIU����M�KN�]�W�Y2�f4�ww4�m(�u��Xnf"�q�Pe$�Ce��h��C4䷤)��c2�h�:��	k&�Z��ZN+�;��k%��Ё
zD`�Lx�R�EU%R�p��]9j��r��wF��$���AaZ��T�m��B�>�n���.OH��z�̡��@�w�u��N`YX ��ko>l���#ud��Ҕ#���w��M����d�8բ�W�8�`�*�`1�Zn�/xo;�oa}wX��QW��$oj³������Rx��M�ֹ#v��N���}��{�c]�3Y��.��巡�B�3�J�}m|ź�TNY���-l���KY+4X�U=0 t�Q[�5t��v�a5��⽒��]-kV+͌�O�K3N�[���R,W�ڤ��{[�R����C+ZM��	�o7n��%hku�2����h�>�aJ9 V(<͡S0F�$M�t����$5�-ckj�s~�i��ۡQX�ܰ�.�fD��fU�+Zx���;O ��g�F�Ã]_7��9�D�+	|)*�W�{ՙz��>5hJH�-sl��v@F��`yv^V���\t�^��� �Ы��%D/Y��]X�Ly`��;�dv�8�=�Ѕ���n�v7lh��̬�K7�R��bO��ʰ��v$R(��P��1�nY6�,b�:ۻ_X$lQT9<�3E�+E埞*ٍ��J��!su�ާB�fZV�7I*�c4��h�c.�f@f�.��ȓF��O,��v�V�mX6E��az�
�/uA����a&nK���h�>8kl>)�|�p����j�^�.��^
��ݥ��Zzp`}gK���n��@0I�nYRۧ6�ڊȬ)�7tECFm̓4�ه~:����J`�A�����C:ַ���j�7F+e1 ���-f�3ۏx��Z,��S��h�ȭb:���ܚ�7�U�to%T��A[� fk¨*E��^b4֋��ݛ�f��|u�yk-<Z,�V�T�m^T�O0�f�D]
F[�AZ���
Mk�'l�sz��T �.�o@��z��i#�mĩ�kZ�9�e[�Ԃ(�!߇�6�K�� �z(�4"&�ݹ� �z��̨�s0i�7�����U�--;�o'Z�ם�[�rg����������	��ו;'�{�UE��qh���K�S1H�Rj�P���E�wݸ�C�[ŵҳ���{0�M�-D��0�CI"m̏��e\�"z���_<�����os���t��t�XΕ�.Ǐf���Ըr{0eZ�˃�P2홯���-ʿ�)�#���k'�e�M�prثb/����f��ѓ,r4��}�tb���>°���oh����fIu��'zHq2�}�c�Б\���y��8�sv��s:����{��_v�3D�f���n���am�O,ƪ�(�m��m��[�fޓ����k[�{p�9�G��Ssz�����=�����]�qep�[F��͖کP�v��Q����S�y9\�q�����jѓ5�|F��|�1m-в1Lb�-)h`M<o%�>2�ĲZ��-ʄ�u���b��w���9	V��@Wt<�٢#�����8�L�Ԭؖ������+�4�.s��"!H��XT�k�jΗy�)|x��-��X������e�
o�띛�������p�6v|���Σ�/
,N�h2s��@*�QU�0�9a�Y@�<��e�(н�p�=�����?�
:�h�n��z�G}���"�6�]�uΝX�(*V�3�K�R�Mr�M�f��v﫵]�/�i�!Zs�������S������=C�T��Is�Yt�e��}Ԛ�sq��V�|@U�̺Ŷ��� ���c�\7�^��ħթ�,gX=�AX� -=Oc�WnH�}�/��lE_VFs=7IG9����(R�&��H,���|���KۘL�˛��"�m��J��ֺXz�e����R�u�����7u���+v��tN�{�sp陝KkX���P�n�������toV9����sYwӕ+dНS~6]�sCfT�ͽ���5,�W�4��k��K3�HTQ�F�)�$ ��N36�|gX�Q�L���Q,Θ.���!d)�\���q���f!����ڲnҷn)y�F�����&����'X6K�%J�>�o^�5pEح�5�{��8L�:�۫7P$��kN�Y�L��N!w[	�sXhں�+uV�3xH���B����N:U]q�E���b]dע���<�5�޸�ζ�{�3	w��`��nP�(���5�v�m����Mϑ�4��tM��w��`�	�,k��Y�QY��֪�dЇ�,6��5�a|�.���Jæ��&��Z�OS
��fز76����NK-Z5t:^-+��hX�y-���X���X�)�1�a����[�,_|V���J�ݢ0A�8�T�l���Н�=�o�j�:���g�ǈ'��r���A]K��u�:0\�p-�r,�3�մ�0헤
�����J�a�zY�ʹ�w�b#q�Ԟ����W2��s��p�u� �a�L_}�e<�v�Ϧ��]A+H�g[�%�;WACJa�4V����o����x�]���Q��P�����v��+E��y�F]�f���l�"�6�jr�'N�[���E[f�Z��M��ޔ�m���R�-z�'=��N?w��ޠ�M���n��5�ӆ������4֛�Ȕ�@0p���x�$!�={2o<�|�br�ޘ�ڷY��r��D_K�hԜ.I� ���+D����� 0%&�0)n��-nU�+U�*���
K.t�E�Y����2�G{�����["���>���{�mսV��˒
���
���t�F����
n�$E�u���F��Z�WZsL�]'Q[����md�:t�lgdgk/�rh,QM�[\�z�;zp������J�o���<8��g����A�/�m$Y9lwv�.Jb#��>U&�N��2^f,���Fcޝ���S.�E͡Q�X�����(v6tP��nwVf��՗�64�Bӌ���Q�xDŕ���26Zi;{]�ۙ|�s/j9����F\�s�E�9ܫ��� (��#ki�y���B[P[�ǫԧ72LB�z	VԵ֭��T��*rq�u���r��ٷ���k\���R�������V^��{��/#��<�?�0L����@ �w�,�C��mi3��i�1�*�VGzN\��������$�\��ՃN����i�Ю6�>3��-!��CFT�`>[O�M�W�S�c�/-�paqr��GWQ�s^*Y�o�{�IT��[;:�u��"�n�MVzY�J�%.�@�� �z�ϻr�G;�FrDW�g��ɀZp��xy��Y�.��MĞF(�wkt:��7��譬*�����0IZ��|Qv/�%���OJZ	w�9��4DF��e��
w���x��IC;C��K�S�B<�'��{��"M��lu��[l6:�.e���ޮ�@��{!�gbB�H��n� ���غ$�!��w%�0�̴������Ó0�ܝݜ�v��&�K殡��ooe$��.-(��mr�[��e�.�����l��GnȬ���,�ռ�Qw���t1�p�>/, 7�ꂻ���$rP�`:��-#���-2�b\���N�����y����M rO���e�IQݗ1�-<�.��1�(�9+F�Nd�&ȁ`��)]���Spi
��50o3$��ܵs��+w�,�R�n��B�]�r�2M�ZYG�a�y�����Z��\u����Ѳ��B���.��Pōa�óm��j\��(�ob��7bm�.�F��t���N�i�s������0�9)��E!�fj���T��O>�_�c��X��d��,a�AL����w��wf��qÈjۤ	�Wu�Րl7���K�ʎ�\���;VÊj��d!�m��lS
ދw�l
k3�d}*�:^��aү�Y�q��3:��Z�hf��q��n͎���Rpo�J�dX���Y�����,^�;gt�K�<��Ch
�y��������Y�Ŗ�;�mq�zSv��(�!3{�s
��oD�Ks� ��w��7VI�By4r�R����彆�0U����H!/'������јU�c6��L�3��>���L����w��aC���qL)�m���upwr�q���]Y$��H%1��b���k57V˰���O,/��ʱ��u���J�H>��f\��eq�P�HZ�������6��{`�2ļ�on�-��t�@f��"�ѣ$bl1��3B���
{���[���e�۝(�}ka���R:�V4ά{�s%�ev��]�0/�ƍ�W�u'��Ϸ�R�[fY;�hݽ�ip!h�|[������&�-�̼se��	�t���hέs���d��nҾ�l=�V�q�\\qh�����0���%y
- 6��¬��:<W��k[�����|I� ��+7�Bz.�8�ϓ���H(��n������fl �]K�7��j�;	$)eVU���e�WG��"�6�6�62����v�A��௫]\�j�)8P8֛���V��:�\�ȝ�z���k�v�!�y ���z�M� c�َ�5Z�G�6{�l59u%��T�r�cv�-a��J�ɜ��iξg)� o#��w̥]"� �&M{YE�Т����u�u�O+�`vr�ԭ��@�N����M�\+喬7Nr�dV٦ᇨ�{8���s'7]R�7��wYm<�u���'%�>�7�Ҟ�ٻ�9�z�KQW"��#�v͜͞�]�Fʺ�����{ey�Ux6q���9�F�sw�32K�{^�%r�*�gF���*����9����B�(e�0S'^�:+�ۺu1k.�H�8
�;���Nx2��$�w���g�3�dT��!�.���}e��En�A��tO,
!gKzj��/�Z�#k(A���>�5�a�ӥ�C���]u!Z�(v��$��37u�L��.�@���.͕45�f�A�T��JR���\?p&�ҳ��*xR����t�/n-��\��`�)�i���� �(�h��Y]�7���G;*��,WYJwׄ�w��ą��N�.l�8F$7�c܀�69]�B}.��2� X��w���>ŔI�)�����a-�,�z�
��s8�h�w�I�h}�{�Qb=5�r���+{���o7�ku返��Ean�]z�`�ՒB�i����"�H5�D���۶�L�c���Mj�X�Or
��N�тh*�u9+.t�RPBL	��]Ru�"}(�%uNsU<�HѱГ��Jm탁�A�[D�]I�T��1�2�x1��!]h;��Y�|��D�ǻ��{̶HVr�J]�N.��q�R���Nx�� ����{/���u8.g�j��b<��U�9��4��c�8Q]āL�;����Qt��F���u,$@Ǝ9%^M%�Ƭ���.8��Վ\x!�uGB�}���j����$�
��wl��ʆ�ֶ+n[j�/�)�q��GC�������އ����a��5*�М�)+��j�j󼣬�\%�0ǩ���6oI|���6�*s�l��c�L�b��J��&'�~�I͢a���7���S��ɫ85�u[k��K�]��a�j�Pܷq�������2�ڴx���RS�J&Mz�/��,�`^d�ZF���#�E�ʇcY{���I+��VK�d��>]�^:�ƝM�ŤK��B�Q���Xq����һ�K� �)����ef��ǦB�su�X��4��M���`޷5��'����Z�*`�kWM=R�	4K�1����(��Eޢ��{����>��'J�r������e2j���),vM��%I��^��o&��zWm!��w����ޫ50�h�9����镖�v	�h5���똾�����Y�o"��XA��`+@�ꔄ�ed�G@��3���|�3���1�iY"�i�MY&�v%"��_e�X7�p���],0�E�"_(M�V-�"�j:R�^���)V,�W���Dޠ�t��[Qv^���p��
�J������}�P�:L8��)����}���]*�_�l���C:�i�ƒ�-�����Ǉ�Q��-��=X����ȷ|h�7&�:��Ϯ�U�k];����ɒ]�<Ju��Z�
c���lJl�����Tz��-��B&&X�:�Y��]��]����h�Ug�eA(=����k+.�⭉U3�T�\��py�Í��6N9�nl��#�ͤ���ڭ��<Qn�A������YU����+n�S�)�(� ���s�m�N�7��7���)7�<��k��Nw�5�퉓&c�lp�{ʓ�-���ba��q*,�\J2�|�ïu6�غ�-�,�0WE[�I:�ɌN"YY�E˛m�v~P໣o.v^��֏E{��7N'ټt.�)���x�����&ٕ����k�� ��+
��S;7���篯�6P�����x�U��׀'A����g[�9)L��|-�{0�ItN��5��{KN�Q)�[�0�% q�V�����I��)�����n�����Y�Iq��u0X*�CS�Au�$�����8�.K�u�#�"'�6�R�����4�/z�9[�-� �Y�(W_wV�ewW]����Yz�Ot�}�]�]L�x/����;)����N�Vl�<�R�ܷ,�HY
��u�5E�e��%Ǐ�s4�	��y�d��[�̝N�r�㻾�!��51�y���́�̱{)9FAy��u����'��9 ��oZ͊�E�>��6�Vܪ���*��7Qb��%�Y*w2�F��&c��-��"�>��J:��&yTp�ST��ю��b�/	Yxcgj<��۹�U�CVJ�V��y�m�\Ʌ¶i��*U�h(���c�+U�/z�[�v��,�+���7t�X��Jؼ!m�]��6�,�]��Iʄ�r�R^�\Ca絻}ܹ����Z�tRqD�doW^&�U��7D~]Y�2�����+qtv�b�1�T�n�%p���m�R�uo�u^�#�Dˡ�x�uH�h�ʟ���0B�VkY�]swSgW`A����Ѷ���=K:�s�d���$��=Å�����o�{�qT'��0єbV�<�%pw�	��}��VF�.2�8� �F�J����l+vՁ������m�ku8�e�\�"eJ�.Vsva�;�[�6Ѿ����u�Ts��n�;�G��e�څ�g) }.Is���_���� >�e^��+�llU��tՂ�#]M�|�[�;u�\�I�2z���q�d�y���pT�2�Q[;gmQd�K���ce����/�
���\�]T��}v�5��8\Lp"CU.��rZ�(]�ٚL���L$<��m�"Qu�@�۝�_e���*�r�1��.K!��bj�#�v�"��P�t�I�Y��fd���=l�Vx���S��=���������[h'�P��]���q�����3+ �e���� ��r��GT��@,��U�-�0����LW"@�Lu���);��Bz�#w�څ��3/w�NJi\'kh��/uh!��u�r�J���ٶz��dJ�a{Q�k:��ֽh�v3Y�5��`E�%saU�.�K�J!��q͑�1�̈́��cl���fJ45u*��ס�vZ��D�̓�S �}��جe�'�:�iڸˋ->�sEpf@�V�kv]�M!������͗K�*�RWr�X���cz �HU��K�]��:����N�ɚѷl���[MZ��ݻԺ-��hn�tqTu����A�`��m�ӣd �Ԛ��&��yYP`��eWl6�S��y��G	�vJ	X�fV�]���S\�V(ݎ)䴪���G�5�ΐ�E�3��ө
X+C�ǂ��=̷�jc��-�����ڰ�U5l��[ތ�/B.WoS}�c9*[ǲ�A[3'An̸��.G�A��}��&Q�� ú�7A�(�P˸r��$�s�܆G�*�Qd�S$����e�(�ep@�Uk���mq굌V��2�+�F�Ϝ�����Gc̲Z*a���9��{aZ�0�A��`��8X�&�����W�p�̨[,���A�W������JQ[��F��=�N}N��V��'Ɨ8���Yr%n�ܺ��u��8��.����M��c����ϡuR���G.;�b1���K;+zu�m
Br	��+F�cA���i:5	�����w�R��%w�&0>*X�Q]K�Lֳ�B�M��I
���ɵ��9V-�+%e��u��X7��.ɤ��͇f�6�ӴN_o,s(���uf7Ԅo���Ԡ�z�xCI)�VK1�#9�Hky��u���Ǉ縳)C\q���X�t.��f�,;�`��-L��W�Q���\�6�ނ�fw;�T������9-[{+��bEs'>F��+����mSN�H�#E�te����U2���v��-���3�u?���o�,�ĕ7)ͬ��G(v�T����@�zӗt���4蓋_N���e9o�m�Ёn���\A�3X3t�SBU�Em��h��椭خ�GdmP��x�c	V[:�;�]�b63)�����/)�M[
�#��W�y�-c6���Ӵ�}�*i��F���Q�Ӏ,$>錧@�c&��{ĥBw8�uc�pQPg� �o�:��I���t��
}`�2�������7�Ao��e<=!u�ծ�B�X�ڎG���oj�GSU�'������^T��gP������.��uk�J�ͺ
�!!cy�Akp�`�����T��M�� ]�����.H%���ۇT7�	H�՛�SV>RuA"��0�@�ZG���۫�o�$�F����<�w��'�y��s���Kxv�Ī��Yo�	nW�
ǅ't�c�*��w����H�3�풒81���b�(�4)UC��;0��>*j}3G$�}�rp�3��)V�n��9.T�G�Ü�P��5��K7���&���\s6�sD�t���U��A$� ��*(e\Xi�&�D��KtT�H��3ӬZ=����g_#D���]c3<7��
�Z]D�̜��`�k��gk��t�[ծ����F[�r�j�\��)up\O1v���Yu�Sm��*��q�-&�5tf�����ڜfTg\��(���b*�ޚ��fꂙ玮�5�ma5ݪ��e)[{.�]�z�Q��	�����)PB!���m�[�n��Y�zsPm�����A�JAvȵ��f�&�]h�*Ν��Eݰ���H�D��}/���h|PO@���n�9h��8��@�E�G�2�T�a�^�kz��)�Q��κk�0�訰d6������\�jU�8�W-VL=��i��p+a�'����5�(���y��?��+�5�.fA5fZ�Q��2ު��ݑ��v8c8ť�i��Bu)�9b�m�������O�Ηf��yә\�;�h�Y�]9Y㊐x��!�@]l+�Q���:��+2�ڙ�k�M�nת(+��sV.�m�[Z-��.s��l���7�Yԅ�ÂH�B=�km
�3�']�f�Z����j�[3e
|鹗}y�7�h( �s���Z�=��;M�c�L��Нn:Ż- mҝ��\��'V�s{�0h�Y��E���M%�+n �^S�@b]��̵�Πn[Ń�G�w|�t�iL��h��a���e.j�DS�Y�����e��-/9�t�� L��M<@t�����4�F%{(��.</9���hJ=Ԫ=������ћH�9`q��ͦ���4����os4|`�3��Ki�Yc�������B�$���e���/�=�
����rR��3h��ʥ1�'vʶ^��H��m*zw5�o7go�4"���f�{���cguP�>K� �7�*}5eB�^9"�7��\腥
�y�k_e�Ϛ����-"��&�B��S�>[��&E���k;�B��1p��;�x)[�;i�COu��tK�E�OS�T��ά����{���\�<�����qm�q��\���yyBJT�#�ޖ�j�w��:�hp�n��:̈��-�-͢$�}��q�J!Ձr�l���
�W+q�8�(��u�Y��H�VX��
�v�M�������)I����ZOgK�1I��W4*��

@,=�|zi�]���fZ�P+Un�������≼�bX����OWe��\tk��V�r�B�V(q���K�}�p3M�/m��j$�PW��_Lcc�f�����f�ގ+w�Gl��*Y"����`�ϟI�����u���"p���f��c��&�LI��_e)�` �DE3iV��5��"9ׇ
	n�C���!4�՗QY
��:�yh̤"�/l�}�0l)����E��[]z�����3�z�/�Y�E%۹�&�u(1:�+��H+)3bX��2�i=�q}�0�$�&<�<���.B]�h:k!E��g�����z���G��Lrs���֗]�٦�c��{8��-�"#)uJN����2o>���̈́a��d�+Tj�#Yۑ��R��d��޷��_ �!�f<��pk��Lr�Ӫ����:��@�4*��T̮YF�@��;�K����(�F
OV��i��Uf��،t����X��L�*ҡLJ[���=�of��79ԆI��w�T����L��:��7XM]�ŎZUˋMXa�ky\�������i��\*h`�}\t
xݼ�q�#���T���V�&�f�=�к�r��+�u��%D�^��{c#S�v<�)�יV�@v�Yia7���s��t+�W:ood��_-�.�I��P�k\�;Vl�ڼxc�0	S.n,,�.*�8��+�y$x���0�Rɤ� H8��Y���di�͵������VrnZ�!�Ӏ��x� ��*�B��!�\�az��w�s�Аt��b݄,H���n�\M�]v��|���|�d�;�6I\���m�l𥒳�fmᔁ�e��@�7Y��_(�)iя+B���S��5 �P��h�e�9�!�w�v*׉Vj\�7���"�ܽ��Zh٧�[���A|�<�	}1
���Ϻ�de�-�	=j�}�}��M���Y��Gب���,�J�ų��#2dg;v;��[��q��"�f�K\4�ޤ��\�;��ZGo�7xT�Q�N�p��F���)��)oٻ�t���t�q̂D�A%MCF��3Y"�)q�k����g%���w�H�Z�z��8����c���&(&�b���ޫ�<)	]ʠ���"�.6�!�\�1��f�R�7��6���r����U��m�!�44>Cv������6�.�dX��I)�F,G\n�TۭH.]���+o�έ�ͫ�s-󵣸����ɴ�f��:��b5��]e��/�8��=������Y.��UK7�0=²���WJ¶-�ҭU�ab�8s��˴*b�V��Y኱�3j��h ��<���>i��c�6�iY�����!k�9�:�l�ğ`a���_�h��^Q!�g�E��\���[����Y@�t�����pM���
/���W$��d�F�ltMeᛵc��e�-��/�t�E,�+r��ބ������Z����h�4��|L"�M��$�L�<*4p�/s��)���ģs;-�W��ε�599�%�&5���to��GS��J�K�������;� �\�װm��$�vH#�àe��{�Z{�!Y5w2�v�@9��n�ra����ħXft�W�h�gp��T������x�$E�
8Ve�v�����⡊���k-8���D���tsaA9�7���w��(
[��0uXm�a�U��s��ْ��2�������n� l0f��5c���R���5��v���3#y��;|23KM�'PT��Ku�̇��p%B-Z���,e�L�����������|+O$t;�=JEn`�yA;:�n���XJ�.���N�A�,�^�4sl?����ዳB�R]�h��+Xf��I��4�W��tT����ڧ�똉�s�Ł��]�c�#"�풞9g�CC���W�iV�M=�#2�Jfn}���;��:�-[)M����+S�{*�	�6�V^b��tB�V�0���w\�&1!�|MX6ӣ)��o���	�v��8�"���-R���ˀ��8[i�*�s&�W2`��&<o���7Pe��+���Z���kV�``��tT��� �3nD�.�[j�C�\�U�57�=��Un�5�;�l�s]��+�Ҍ��0n��\&e6%n�ܫ��$;�wf�W}��h��[1�s�fɥ�v�ғ���yX��P��Uv��7ec��[kvkwsT7]���&&��	�v�k�Q�����\��}6���c�`��h�T���9��tz�e�)υKY�,[��wrf�������(Y��n��S��o���#����γ�c5dQɆ;����h��>�5:�4�E1�Kh�˘�+���M�*��`����Ki�&>:�l}�.���E(u|�M�X�+���4	�-�:�QC.��c������U_f&��6�8�`b���x�9�D%��95���Γ�1��ܢր�n�+�38�G��}η�e��Yo����b;��k1
�{��Q��uor�p�xs��K]]5�7��I9[� �2��c��2���S�����u]�n����l��ma���Ư�ĵ�m|�v��s���r�w0;
Cz`T��p��}���GaR�>�R��j�3w8��A'��rH��)�-�8���]�I�]m�.�+��[��-p(ؤ8��K�F���l�D�[n��E�=0��[������VR˥�A���F�>Aʚ��<W��p囘���b�2��k�Ȥ�������\	-[�
@�ϐɜ�t�[��K<f-���ư�4#jf%B����p��L�EwŪ(��"j�rXo�>�sXo:���a��Uب���]�؃��櫖��Wϴ=-6�ͩ��5��ۘ�]]��U�cM���;ك36�;�Γ���]�,N&�T��.�Z�	|�:�x%&�#��­�W:�uh��k�-	�y��0�5�;{��tq��F��S�vnԫ�:'Z7BfM�Ce��V���\s~|�'Y��/sR��^�4�u$�RBh�*v>�lZj-���c��6*��a ���`�$"w�������	�+:n"�i�G��_�lU�#��2�x'Y��V���J�q]�P������\�J{�7�V>8�1>����_db���	����tc�0�A�T7_7�i|w+��l���.se�j����t#dwl�Ĵ�¹	+�	1�q���]��m�K��qЧg Ū�K���ׄ%��gGŵ��-8_t��U�]�ŕk��s�g�-�mu�r��v/� ΅�@<g3�+4�����@(��l�Q���M�om���ݿ�;yk�x#z*�ْ�6�=��9u'�8�t�L��M�;W�3N���_�߀�����/���2Cw���� �������z��ir��$��pNm�߭L�fYտ;L7���Ng���I���ww���z�G��W�k;�|^k���4�6'Vk�\F�hs�I�I*�]s�2�sj�N�S���tA�1���_
?�C�]DN�
�ە8�n�{������)�Wqm�Z,
ݶe	4�5�\f�����kG:���wI��=�.��S8FK�~�E��g��q�([�2�ȫ%Y��s
n�ʤ�]|(Zo�ټ�Ҷ.��}Α�癒�:{�h��Bܖ���ZX[cF��bb�ܗ�7�89�������@���<�>�%�e��:j��/r*��<g �=��� �����˺EW9Y��\@�����f��(]vQ�A�'l��)�	�Z>g��-PΖ����F�w>�c(�Y��H�m9:͛l��V�+;+4�Գr�5�]n����IV��{]4 ���C�"C���_n죏o�r������q��ҽ�dN�GP�%b�����ʱ��S�����̜�Jh�wǨ�F�a�O�7�ln�!&a��]�E��ՆtM�W���%0��r�r��vqQM���q��,m��:����soI�#�>���J��4\��"܀��:f���f�K���U�n�\f8,e�V(�"�2�D�E�T4��"�X��.��\j������b#2���H��d��E������"����mb�ëN�+AW��Y�[���,h�b�����r�h����N%J�jɥ�2�j��l�Eq�����,�����T�[5IEj�(��1"�&�*�LB�TYF�,r�.e�6�
��ԱEMfdEb�(*�UʵQGnQ��UQ
�N��QUX�+�Ĵ��`�t�(���5r`�0պ�4�%DA�+AUU�����V���E-��5,U�E[qJֲԱcF6�(�Q��uj���Q��b"KKED��#�M2����X1�aQ��ET���.Y�EUF0F0D���a��1r�m�Z��%�fS5CH��b*��F��TU"�I��.Q��
���nQ��O?�?��w���3o}�w-��V2�Y�& ��ஓ�2��M�����d9Mu�ӧ|0�WJ-ɸ�2BY�U�&�M�o����]8�3>�(�2���)_���vtbͪ��q��>�$�2`��>�rU/g]|�p
�w��]e�Sj��wΚ=I1�:��N�9�*Dc�|�3�����n������g'2y��zeu��'��Z�'/k�	�ȾH��n5���}j�N'�c�K�Xq<�	�"Wb�)f���i��2i���RA�[~���"fW��Q�{�J��f��ߗ_���ϯ'�ؖ��<�Չr{������MN�:�h1j��,��C��LC��
�#��Gj��sQ���ѩ�vլd�^��;���.a�mt�/�Q��#��J'^F�3η"�����2:2�c=���n3�>�nz4J�T�ߵY3ܕ�Wͣ˚���ɀy ;:e����X_;oh� A���/�{"�}3���M���Z�6��d�xN`�+yV�*��fVZ�F���9�l�ҕ���q����P��������cؙ�q�ד�of�$�3��Top���]'��{��r�k>sE�8�"_P�(��q�����QQ�f����^�>�6�M¦n��/Λ�=����3��N�<�wB��9N��7Uö�.��'eڜ��#�W3�mb;r����;(=�a��9𒺼�8�5^�q��#R3�����39[6�dE��g'�mu�uG����n1=�}]����c�E������I�����Bx�o[�{�gpڛ�N=Kdbv�2��7fZym��ƽ�"�O?��-r�z��x �k(#	~��u�˾ܒ�</9=f��h���q"��<�O��b-J��8����?)��t#�:a^�Նv^
�1@μY}�v��-
���||.�sՐ�A�[kH��ɥ�R����w�LD�tD�b-Yy��n��m��{��3��Ͷ��!��_	�_=�1���G#�x;��_��)(���$yр��P�*nE�1�5�>x��uZΰ��9�)
�����F�Д��zS��'gVn��_p�T=ir9���z�L��n;�3��E�<�+�i6�Iq��b>��Xɞ�J��<���=�QϬ.g�l��4ޝ��˷-�3VQcw��]�~aR���6���{j=/��h���i,��ByCp�!9^Ӝ��"�]+���!���h&<�7��#7���wo�뾹W@hN��.8'�\��r����kj\�h�\��E*����������	�]�n-��j>���!w��Z�6>�Z�Y�%��B>!�%rT���R�W��,���f��kΙ��_v��ϲ3z���'�sa�Zhi!��=�x�z�{�����޳y��;[�8K��7�v/�b���݋P�\�C��j��3�G,�-d^A��1j#�6�^��-X>�P�9�v]+l�k%]&e�P,?q����9�=G�����<"��Qu�*��7z��m�'l���cG*NY0$%�7�h��ϯ���l�5+���3&ٹ:M-sz�C7�A �dsa��|l������l��Kʝ����o����\ ����WEz�A��5�{ރ��>�>+h�5�+�Ns��䧧y�Rc�t�|�Q\��6&z��J�o1���DoW��m5l���b��\[��=�kΓԢ�3Q>��AO^󓇍&Y~�^�E#5Z�%�Jr��z�;��J(�t�t��R�O.�|��1���r���<�M֟��~d��e<�}I�aGh��,eN����p�^=y��w��Ro+J�M��8��Ni���?���@���}�z�3ɕS�{���ʇ�eS�w͈��������,z݊�h;��lJ�o��%�<Bm���Xl;���N�4�dܽtrv/ ������Nϕd���r�*̘�}���K�C5Q�� t:����!r����B�� ��\ɣA�"_���|+�glAV�w��*��-:Q<��% ������qQ�m�ۻͦGu�y)[���!b�_b����ؘ�X�8�����ј�Iz��$93��8>�Q���.6�[!��]=w�b�߾(tل�����%ߔ��/U������釽������No�}�`)�[	�]I�<�oX�;+��&�/Y������8���:��F�Ǯ+�1#)����5X�d�y8|н�b1�}e�;���lJ�¬��,�����Ym�Ů�{�C9�Mf^�X�[���MfF;����Su�,h�%k�x�3���[�O�)���c^%=Jqߨ��k�	�_8,�^3����0�z����ڼ�K��>�ז�ΛZH��X�׼y��:�O��ʰ<�������y���u����*��=-f1i7���K���;�;��Z�狡ov �lyA7l%(-�kN�]mMڨ'��N�
��)S�"�ZC�B�?cDeZg2VE*,rM��`u�wP)1}OM�v��2��N�q��'�C���k��:���=ʯn��r��zԆ�*�y�ڥx��Ű,t�B)��Y�.6�}���򼲔_'|1ux���69j}�10ϲq��Z��q���TdmS�ZLv����9�����D�97[��׻��r�<bX��C�N�����҈:�Ɯ3ηt��lE���qI����#ޠ��=Z��>���l��b�~3���n�Tof^kQ���h����"�#1A�z<����\Τ|����9z����a3�w^���hܴ�D�
rb��:̭�f�W۬.��U�\�;J�s��YSَ���~����s�kh�V-e����DM�:b��vs��_H�H>�㚌�B,jhS���u�G�C����"�]q���3��63S��v��t�2�<i�\z�ӽ}8�p5qx=�PO(����#����G8tJ&��S�����&Z���&�{۾Sm����ڄ/Q�y��~�G}/NHtb(1m��_qׇ�[�����jG=@fή��u�	�{�s!��fl�K���X������])� �+u5Nd��Im�0�sZ�(���yS���J�旋͜��t�v�xyܛ6iQT��E��G��+J��X@Y��7�k�/��Wb����p<;y�j�3�	�`��#�g��bv[��>��R�Zt��b��QZ�kY����,BڜB��W��]s竇�W-ym����UH�ĵ+�O�jQq�Z�
��8����E��/����ff���
��չK�򉴅kΉ|ʿCS��W�6��(G>�����E��o l4�yGy�i�f��)��$;��ϧA���O�^ӛ�އ۾'�S����T*�qP��~s�\(�v�}}oڑޕ~#��Bk6vK<�c��U�o$L��'���ϵ�we�֩u�c�Ӊ�X �U�i�j�|z2���#D�ΊC�f�+��!q������Uf�6��Ֆ߳՛�1lWy���i�����P�j+��)T�F�|@Mq$�ԟ s;	��m�Ib���6�]����s��:I��'V�6���Ļ|�xd�����F����Ò�;$�7�����.8����������}~΄8����B)Q�/{�H�y`��v!�gP���FoU;R��pn� .lEЇ�ν_4#�h1؜�t��8��Zʸ�j�L�q���e�W��P�{�V�9AZ�qa�n/�egd��Ʈ/w����~�c<�1��*��{�R���0u��P��
�y��vϹbp�;�i�{�{wc���zY*f�> Ξ_���^�S��59-���ú��L��{��OFw�9��{�buu�����i�\����y+Z�N����U�1�1�:С:��ӭ��|P�e�̯QG�*��Oy\�m�̓Vi��������j`귱Oc1y�S��Z[݈<��+ɻv!GW����T�	�Sn��Y#���� �����M8K��N���#n�<Ғ)�G��7����R}���mHj%d�Բ;��]�2�	��.�x3�ۗ�3ve	7����1�D0�Β"�\[�N���O�E)�܎�;��0oD�3Z�=]�>iPG���]a�Hv�&���(X47Uj8�Ҩ��Y�u�}�bt;5KS�w�|�PYr"�Z���ìjKj1j|�R55ޜ�D��AǄBw��ku�H�J=�v�����z�����)GD.�k��u��ī�h���>�sJw��/*�\��ʚ�t�L�{�q�C�*t�iq��=Nj/Gs{n��=`���K(�v�&(k�r3�Y��Z�b�VV�X�4z���.�����;$sɳ�GY����WNGX�2����	q�s݆�QW�Br�-cq`5���瓔��>���#i,I�U HX\���v5ԯ͌�o8�v�y�{'dn�����1ϖy��U���-~�s���<���md\-�ה�x��Of+��	m���o�T��ʃ���X�&-靽[�_��l巘i�=[�r����ټ���=�Y�)��-���0�7g)��TKMqc��[z�X���%2��`����|G<{sDIᕇ#��Y2\��"y0�t��Ï6���w�E�I1p!���� �Gq5b������y['��j,n���x��kIY[\(N�l�ӽ�5mc��ҝ�b��z�;~���Ϫᘺ���=�Z��_{�4�ys����u{�.��؃Ϳk�	�w	J����t�02�Fi<M�scM?C#�*l|�X�����c�����	�5u�b}d���E��W6'ћ6��}�zH��v1:5Z�혎�S}��m5=7���hz�j��J�q���_���y�t1�;�{�^?�).�'����g�����gu	Ք�8Q���GG��<y`��<��lf���_��������I�M��4^y����<��t�eV���*H�A�]
�䳮F��3! Gr�5IE�n��^�����ǁ��LM��j*�n�Ӈ��(fMJb�i�K3f���G撴L�b�X�H�#	�V�a�V�Wd+��V�D�U�l3���1�ChG6g*�'`�T�Fsn}���[�ك�-R�b'���/F�u�Ű�>{��V+��s^
=X�$I���h0I�F� gm9�梛C�uڱ
��v�ξ��Ú:�7��)��id*���k�ع7�s�4�W[�ȶ��aOP���;�')^��T,�r�6KpF�mn�\'���xi4Z�u䍈�m%�v%e��*$8f=�1Q�.�g&[��kf=�p�X4�^awS"��o��K�W�Ytg��nU���j�����ëۇ=d7}�\�t?m!�\��Fs�Ի92,����eꧨ�:¡���|q��:u\�u��K���U�o��si.���HΑM��\���+MpGi����P�YZ8� f��W4K�_bX"MiM�ņpI�Y}�}�ep���	���c��R�4����L8����|z�8x��(�Q�J����N���tW;*��R�lJ]虠w��+5�Y6q#��WO!���4Q톓<�z�36���kGmkV8u�rI!��MIg:�<�;B��x8mm�o\
-ܶ��������9�K����bu�]��ʗ�^�f&�[IF�3GD{�vb��ږ�Mˏ���3�!�MA7f��R̈呡}��?�7����8r�h���gY��Ern�XG��l��d_0/g�ldW�:����$ �xjޡ�2�=�e�������t0R�wSγb�ɻ�l�1X'-e��K�z�j;�R��dG�ݏ��u
�[��.�3�ݓ9��5�$��ټ!%v�� ���>`r�X�1y��>Ir� j��"���<�ta
T)>�|m*�XZ���� ��ku����Wp���͏����Cfb�����ucXQ�.�\#��I|���;��T�eL�AJ���:WZ�h��N[�/V�X����(�+D2��Juf��N	y{W���܃�S�J��T��Xe�X�*��;��EN��E��˗f@�#DSdū��+pގg�@�[*|���ɲ�������r��NN�i��M�/�sҕd�V�VJ��C�#���k���aǹ��$s�ځ̶ݤ�^��YD�����B�6�ʘr�T+a�d[��ǯ�5�,��l�؜i�,S�	�;���(켡&�~��8�ͳt�vq�c��Q��:�Xow�\�rA�nf��2�y�)��)�4��9*C��ݑ�Zؐ��Գ���a�&�̚��G9G.�l�Z{�����3��_�z�9kgu�܆P��/�oFadr�"$Ų��(VVnZ�X+�J��"�R��\ƙi[�F1\�1U#VVVЩ�AJ�C0���څ�P��4l�ƪ媣YF"�M04���c]9�e�j\�GVJ��b��b�R�.5���TuI`�R�4�V,���h��T4�]5b(�����+EU��j��kA[j�0ӫ���Ҷ:��T�q��sG��3.e��V��̭LLb*�hjㅴX�m+��˓2�Y�U�2���6�b�ӆ�p2մ�iT�-�mF�WZ�n&���U��̵�TKi���֪�2�3q%V+�2�KK��*�,S��&�X����
�".���X�J)�l�ba�]5b�Z�F��ո�)������F*�j��\b���D� g�Z��?)MV1w��ϫ�k���Z����N3H�A���m��A]�gbV�]k�Q96�*E�dǯ�q�����z,��7��q�h�Q���+�);/����w���	
�ٶp�ftŻ��Հs�~\0�>V���M���3����劲r����/L}���>V�x�g�2�O+��*��f�G6x�ܘ�yC�{�k���%�2����>�\�D���P�}Sy��kܬ+�P
���HN�o^�Z�B��v_j{d)�}
<t/��+\^/�ߡs���9^��T�x��{�Է����5���,S�z�{A�<�{�J�;-�Վޙ]z�{��;(�:9������K��S�;�E�>z��A�gi�*��E����5)�<S��v#���`P�\r�"�Y���leb;���mq��15�-3{(���Ħ��O!��_Q�o�A��>�y��xu�)�7�>ǨͲ�]���K�N�s�����~��3�iq�Q�a��1�J�UEX���ݾ4�rVw�U"��t�s����2=�t�\.�'p]������W��I٧�d��2��T��8S{�޽-<��p���׽�pO;����­��ʳly���ui�)�<�81y*����\r��8>W�S:+�,�k^[�]oa�ќ�ycՐ���Qj���������"7�Tb�U�Dg�nd����_g�A��Y0�(]�E��v��S<�s�>K<�Ǐb�/<�g��Zܠ��o���B�CY1�G�I���ꦬ���Ψ^�x}+l�u	g&��Q��C�/o-$;.h�ܜ�t��<�p�X��!q3j��>�ˊ�����φ�x�`��)G����W����'���w�x�̪ᶘ5�Z���GIۜb���J���g{'KRn�9<��cǾ�VX��IΊY�w�������E��<L���3�^�{tJ���e�b�L�+&
�M[�N��{E��p醎Y<�i93;涍c���b)�[�<�~�x�r���"{UJ}&��8UȝO��x	}!-Q�)�n1Ah��ٸC�{�A��W	�(k��4�)�kΐ�����`�J�h��?oWcvf�5�Ls�W�Ӊ<��8�"{o,r�]~�Ĉ��Z:�_$e���՛|U���+�!�^b��<���K#�l��:�-ץ�x󊂋�[ȘTNW��=X���,|�-�y���&�؅B;k�c)R��r����^O@\�����P9���ް�.���UXMO}��߯9B��J��㪹��fi�'^����ؗn��+΁̭�\�{���W6%ߝu��|v�u	��������m�E���v��S̝͆'H���:6WTaDV��ػ�n����=x��]+yOS�;.SM�B*L�>q��§Nv��ڌ1����Mi��{��kjjc��a1�buME�n�p�_a�� ו�~���.��١=:��Ȅ�I�n:,�u[�F]^%Pkp���L�Ջ�9�����O��������E��0���b�'��j�.�]�ɀE� ����je[�#���Ȏ�ń$�|���	�x��9�7�7ug�w(��2�+c�.���y6}���/]ϳs:�o}%�xKؠ����+��%+k�j2���G3�WFĢ�/s1&�w���m���8�h�����mM�m!5�]u��b�(#
�9q������/(v?GDL^�o3��۹u|�=�ح0���=�Oq^��;G�f�\�O��f:��b7N���-��v|�'���׉�*��ݫ���}�aby�T�Z��|���GÖ�����yO!m�7FOh�T�pD�I���?J�������.����z�v����c!��+ӆ=#*J��_��֚�s��MS�}�S��H`�%��W-p�����-���>���zO����tsS��T�r[�>�N0df���B�V�!v���Ȇ�ȹ^hDU��mj�Zk]�I,hH����e����V.�r5g�Q�o[��;l_7_��x��i����.���"� TMe�>nuԳ�ͻ��W,�*L�iP��S-�l�(���Ns�T���v1�޹ズs�u��}+�>�8��S�;A͚�I.JLB�՞S��N���[�VS�+�ъ�\�E��\QJ��.�*�����p�śbN����Z��+����:��4
���MiU���q�8�����Dh��>�Z|��jra=�����Wn��(��q���Z;Y3��L�#v!teve7���ź�=���H�+�휛!���ڱ龡(�`�}hM��Bt��g���Y�b���ke�}�o���=Bc��4�ϜO_��]�.��j�;Ũ��H�}8�p5qyu~�;#F�����q�W�������.o���aY�J��9ރ�Z<J~�t�Z�z_���^�as�����<���޿���gQ����jn��ʖv�MA�7�;PKb�W(.���0\�C��ԅ+�v*���bmoL�/����#s�p���/�[[.���,�=J�C���o���yR�K}h�.G�bs�B�`}g����
����8��ҡ�������ik�y��R|�ۦ�U�3�V�>#���Y��u̎z���@W��j�D�O��k���ߖ��ߡ)���`U)����G����K�vi�<�,Ku'*�S�~^�_��ՠܡ�B��B{���\F��)!}��s\뉻�cv}W�y��7���� ���V�c!n�L��o��!!hO}q����~����DEgծ��N�XF�
�ԔL��#�hV������؝����&菭�E�,�`�=��,�-�rr�a��!A����+�.2�c#U�ʲ'bV�ҥ�H*O���)z�i�����=��cM	�}N�Y3X�ه-��vF.�B;d��q�����5��em�z����'�	ͻ z�?0l�N���8���6���$����[0u�-�ſEY�1xK���̑fe��,Z����������ZH�k�20p���˝��W�5�:<�zV �tZ��-��[�i�u+��qe��q7��9��8�v��$��ݜ��+c����.�vd�y8u����M�˺�L%	k����`�W�OW�2���X�5{���'��{��4Ķ?f��^n�[��*�����)�jQJ�owYةީΓ}]�<�r�S21�r%�wm2w���j��yo�Fwe����z{S�m�oQ���t:�N���]j oWoe�qM�����a�ݬ�ԛ/#��<U���?�#S��SN�>r�*kd��w������y���%>cf�����8߭<:��l�+�/u*;���]@��Kz��~}A7~�n�՛���y��)\7�M�G���x�����]a�K�k����]j�>���כ�#5Ʀ��t�������B�8�vj4�;��艨uǳ�⍋[S;R��[�KgPA��f�)*��\�k�s��� ������]�',PS�ans.��b8TL����^��0y(sŬl���c�[�kr�ckvP�n�VDv.��}Q�yi���Y26l0XL�nP=�R�-z?}�r(u��3�2���xa;�G5�ulJ56W�B�n۝��%���Q״#ʳ�k�W�U��́��\|cq���S����T��z�C�#
�9���㐖ꆏY�J-㑂Un�@���d�
rb��dJ���oB����cnU���G���qDM�2�+c�є��䄋̹�3ov�xޤ�in_\b�7�l��Z��)>�������7)����̣Ş���=Ke�N�^�}q�=7����[^�q�:�b>���-2��[D���7�
����]W�˽׏��5�bͿ>=$M�\�}�#.s����l���y��_�������au����IZec�U^�����oH�ז�ΛQ��'/����T���c1��k�mzĦ��	��*e�b!�,5�b��ʱ+z���âB-��� ������ �y\<�f0��'��:opUɉg=�.C��U�ޡ|���@�����Q�-�I���ђ�7ze9�t~��6��|�v��cy���\V�X�o�@��S�~��:}T:#�K����sF�P���o^ �lk��pn�z76���o��mJ/��Y����q@F�����Q�C��R��q����|�m!U�gD�l���xCᑶ+�ڸ�wc�Cク[���Nar��#�)�M�ޛ�����S�K��ͱ�!��"^Lff�w9F���M[��$}KUؕb��YO�w�<�2�׻�ٳ}\�lGkc$��<}���ݤ�%�J"��󎋛Q�*`n>�7�:�����ϩ����ʀ&�n(3&ݺ�E�b�,���V���_�b��t��;�d��u���L����@����%���x���γ�.NB:�驾�e�9��оŌdA�O'�N�����؜�-������$�����f���7�Q��:;Zp}}WXҡ)�Dv�k��t����Re�E`�{�:��N�:��Yvv�
�[�j#f[)Z-Akb�4��4q�C&L�I*CJ���u.������[m��͡���'E�;��;�:�^���No��qG`x�4�x�ڷ|�[�;T1�ۋ�{��N�ɦ�//��L��w33��:�V��\��ik��æ��Ԣ���9�{1��k%o;�Ew57�ٶ�m�ê�kkӵ��>�\��W�g'��(��K]B�wE��r��S�J�k&1�$A�Fq�{π��G%X���	 �$�)���Z��睾�Y��'��Bq
�P;�s�y��ɩN�ݮ��oQ���/t;�֙n݁	J]��Bqb9t}a[ٷϯn�2���۽N��7�m�c������~��.:+�w��)M���kL�}W�>�y�\��y�l>�wSC�N���*z�C��0�������t�]dC��O{6�/�'+sZ������Ki�����R+���9sa�w�R�쌺�+[�q��rΗZLhu�!����0{2��f��������2�8�=!e���8$S2fr1h�����9l�,W%�}ux�F�X�E[�����VE�dy��Ӏ`��;%�wX��8Ʒ�d�bV9���721^Yʵ�w)oT�
�;��f�K,Ӈ��[Y���y�5pt�µ�������98[���DHr����'S��y�n��p�<��ӷV�\��(��rd^Ͷ���[��8YV��j1.a�N������,74�gK�ϸ�qjoF�T��"k&��R\]���w.�zx��NN�-����*�����S�����F����&\�L���&�4t������uvo��K�l�|���6�A���1t3�l#�6�s���u�9KcJ�&�����
쁔ռ� �WLpWŚϱnޱ�R�=]�B19��7��<�سǄݎ�ҏn4�)���]e�Ӵن�~R���u=1�to�;tp<���gC۬kr
@-ҕ�����ㇵ�:��;��m�<[���@o�.=9�cqp��1��k,SSh�hi��(:���i�j�I�v��{b"��f]����72���K��K��6��H7�d�A���/\�1�IKr�v"Rt�Y���Jᣣ��Mؽ2�?��7������"�*�HS7�NΠw���C8�8/2�[�.�+{�ţ"�J�c����J�����֩�g���O�J�u�W5j$�X�ce%���h���6M\O/*\7&mH�m:�B��.� W*ңľնMJ�N�g;7��{V49��{�|a���mX{J�!�P}C���kn�i�Ҧ�&��oFO�զ��,�.R�p  �&f���Jut�S� %�P��7]V���G-5y\l�2�;b"	ũR7g��>�u+c0����2��� �h˭��	��)��ٶve˽D��: ���{Z�)_>c�
����ݨ:��]�\���K)�t����4i,3+d��+<��U�;{�ǅ�N@vr�Δ%�ںI��4�,w�*��h�t�}\Im���H�]/Bf�ƌ�h�>��DyլJ��ᙑ�ɛ�;M	LV�P����<�W́\vb�y>Gƺ�崄5>�Ӽ�WWv[˹)[����V��M�I �8� ���̙�fl�M���CzjP+��H��*�H��]ٴ�c|F�m:O ;*��N�MG��P.B��1�X�7v��"�lӂL�c�ք�D�÷��.�0���KB�F�ڣ��%+#'lv y�͔��L��2U����O�#G�(\)V)iV��<s-X��b[AQb�2�4j6��Vj٫\���A-�eZ4�QL��.UE*]YQ��ш���4��WkW"�9f���TTƎR��F�i�)D2�T�p�K3)�EQ��b����AJ�Tim����q,���H�.�QTm%eZQV[FڑE����U���j�J*"�-�����b �J ��D�,�U�1+P��PTˬ�-KV�L�TQN��-�kTX���Q���
�M%e��ӈ���[&2�1c"1��X�h��3Z��Q���J!��3%��QEڪ
 ��%JlEQ\�b���������}���Ѹ��K�A�]�7����3�s�����K�������
�j#kin9J@8��8�����)l�~���B�����T�Y;�1;۟��}�M�|j.���1�?H�ǘ�f���-ބ>���Z�(XΫ�����6ݦ��js��w\����+���\���@N��p�ֲe�ʌ�Ii��q>R����)FRv]�ɡ�G��':�����5D}Б�N�"E��� �8��.��w���=C�hF�@s������w�kl��.����5�ŵ��g�͕��pl��WA'�J��\{>v�ԛe�ԣ�op7ݺ:$KuR텹z�e#Ժ�����b�xf�#�j�;��j�~��{8M6}И�OuO}9-�E�z���Q�U�R�he�WZ��u`�i�x����/1a	&�;�	��Uu����hX�N6�Rڒ0�Ь������Ⱥx�b)���l a�n����A+~�ܱ+�Kn0mY�t�TC}҇���>�Q�
Z���l�Gg����"[&�Ӫb6���g1�/[�s9��%����0��7�;��StK��5�&Cl����툪Q׽�6�v�T\:ex��{�~fվx[�ѷ.m�]���>7<��-�����K{��o�e�Z2C8.�e���1����P����)�7ˬ>�E�'9�%� ��[�kjz��(�q��]��������GԵ=̮�r:��@ջ{h8�^��,���yU�@�Po,تA�����'7���g5K[��nb�EF�Do#8(��Yٵ��1_)�s��]���kK}�0j؝��]Cz�	,2�EI���8���;<���ҳ��9��n��v��H�L�jrb���yՌ(�Y3=��w`��bׄ�n�c>�"�H��]C�����3�E4��	�ٷ|!Y��"q���Sf�Zȡ�����וS�y�W�g#F�dy���y#R8q�g��	b$�7A�νNI]3�Zeɋ*�s7y)p�^+r��z��&,�ј���F���Z/9vc��Kt���僨άJ�p	�=Ǡt���-t[y}%����y�O2#0̵�Go�W����E��� ��T\������1��|��������Pf�%�3[R����œ�,���N,�j��}(Nu	��5 =��n���f��/aN�=��PZ�E�[S{�W�����Iu�Zs�s�=q�_������|�j�\�㷧Һ�<��Q��{�i�om.Ť�O)�ǚY\�P�wI���ym�q��i�܊I�\o+��f3(J�Bw�据�x��[�1�УnL��;��U���K"m�??Y�M^�9�cj�B��;�o��C7��t5��$;D�5<����T=��7=*�}����%R��5�)��󅈽�iA�߼tVNao��}f�g���bڂݞc4�Z���MydS�msS�(���b��8V���帞��D�ow���]�ƹԪ��mg���'fp;Gݱ5�#K�y��>F^��9/n�J=Mu���[ٝ*E��B��/���2�e�7��k̄qdJ�Z��I����G��nc�S��	j�}�UW�/�Hs�x?P�LvIp��>5鉽�N�DP�ĝ����tvr`eobj�RQW��,ﶱ���Џ*�@���+[��n����b-�Ǌ�~�ɍc�	z2��;�gZɚ��<�{n;�X�:K���Vh]�����Ҹُ����5Fh�ka>���:�\��ݘM]���Z�Q�BX�5��+��l�zau�Ƀo����N��f.�g����#[�E�o3�cMy����;�y0t��x-�[Җ��UC�6��u�R�
���|��uR�x`�3�{�n�e�E����,A,�eNScd�\�ϵ�!g'��yp�F�'����$z�&5j��b�'�g�*����W3�P��P��9�g˫���I�M��ZD���Vk|H��}H��y���`M����ֳ�
>�8F�l��o36rV��Z���������yx��r�[�K�m/p�<W�Zr���3��z|;}�c���R��/0PRM�9�o��m�Ý^�eP]��n�yL��0�n�W���/^Z�,��P�7�5���������L���1���q}��ym�2ݻ��K�F@Jp9t���0:�N�&'��^��{��c���tV��.�Fi����]���]$�'a�;���y��[��>��B]o���!�,U�wR���)��`B�^���U�]{r�f秳��W�}���
6��r��n�Kf�Xf��F��r��
�'*�3��WCC|���&o�/w�4Ze����8����t�u�z���+�25^h-	�x���1�� xo=Ȧ
oHTQ
no��5V�>y�o��uI�ŬamR�˪�̼��R�a1�FPN�Qs�X�o��Q�Խ-�}������S�'QȺh��}Iٓ�'�#H���<M���0�7T�ܾ/��Bd���J�	�W( 5��Wn�I����!ȫ�s����x
>�j�NdQ���ծ��	����=�צ��������%t��u�1�`Zڗ�������G�Q�org1-�3/d�q�vaOW��%��Yo��X�'(𷹵s�����K��c?���館��{�!ߝؾ�6!|�.=Vs>�s��gp_t���v=�Kl���0�^��͐ٝU}�F<���Ci���	Z�9��^xrB�i��O0+�M^h׽F�j>���`^����߶�u�����NZ�'�U��V���7��W^>&6GZ��ZuU�q|c��K��gj�/��C{8�<��6�E����n22��@��2+�:.�]�Wa��-W�{�����b� ���o_��z�PMۊ�qWS��$��Z��~+��>���T���w�k�<1u��'�m��u�|D#{�a�������sa|�l�mxOv�q��=����zʽ���m�[�C5f[����Bˑ]nv��� K���q��hF7�^-/.0����e1��'��J�J#O+��4e|{P��g��Z��[1߆���^	|8I*!e�9R��W:�`9΃ΧԌ�K����rmͧK5�ĥYIt�P�j���s���cG�0.���n���M\��vC�fvA>��}������'۪_v�:���uB�I��s���Mn�U���~�<]��\��˅V�!�S��H�%�Q�&b���}���S7&���JUG*t��.6��:�>�=[��)ey2]�Ɍe]�1�C���$�"m��·V��21D��%En[����ggsw�:��k]=W�c����lf��t�nu�W�g�)sB���QN�^$�M��ѕ�{&� �rګ��0�:�@�{4�0#i�fSG̢���k|y^>�;�KW�9b�Ceu��]�z�\����s�Q^���ؽ\cz�w����i*����Y�̄���3w�TgMOI'N��W����dr�ե��ޟJ��OgqŊ�:oP����lT�Ɨ��F�#�g��5<8�so	��b�]^�����պ�f.�VM�\���u]|�f�<y����n���9K'\� !�+q�P��1m6rP�h�v�v^�t�ӎV��ѐ>"��/:�m���l�*KR���X��m�ߨ����3�[��8J���ʽ\XڙٕBCҮ���3+2�[c_�][_vd�SΕ��.�������5u=�N$�{�ݔӷb�D.�#��olN����j�H)(sS�봐���x�c�X}���=�c"�{��J-~OM�~Y�5����]G5�Z�w�6�O�WӤGvY�M{N�۝�G�
G�r�O��O:��KUܫ�s�H�S�O���r�W�鴗����k>
����8����T�z%�/u]õ�^��]ϡΜb�ɹ{��,��E���9�B=�
TBB!`�v���� ���<[�y�m���ǧ�z|�ߕN�UNE��M�QZ�iO��͠��	�FPN˰�&��u�'Mzo�Yj�9�*��p"��7W����)��Zp�-w����;�����}�7��z���7��P9|S��"�hot�wӊ�����Om~+��/Rۡq7���fA�w��5e�w�i�$��ׅ,4��]�Ⱥ��(��L.�n�vM8�w:�ea��,��q˽��U����R�����H)�*��y�ɏ��r��8��9Y��7DR�>�e�֍[��u�߽� �m)��JY���a�����;���eOsTצ�*0��|��L�Ҙ�l�8��k9ʽʬ�k
�Oi\`Ua����a���=E���x�Q��ګ���ҷ�O����"�z�E��{��|3v���u}�`v�+������򁕟P��M�ζ(�����'9!O�+���,6��n��SA.�	N3�,;����I�ִ��E��眔��!�Zh����[���+rvm�m)�1�7�M�}q��U�X~^~�pw����v�ܵ��ҡ%Ond��*�>���b�m�˨Og�ʶ_�i�%�.�,Z�w�ԧ�׳<a�)^���}��b��'{��v퓻;V�.:�n�}�m����oB�ʇZ�o��>��ċ�4�V�7���|!]Gw#��7����r�tRX�ff7�H������Jvt��%�O`����Y��c4�=>ś��P=T][�1"TC��>��G;%mq���y.u�KB�A�h���ߞ�2P���+��ZjKnي?��U}UT���tS֮>UN�qH�����h����jt�JV���Z���=���{�e
"e%�e'eߔ��՞��	�D"/.Ӧ���c3�(J�����Q-M�@�N�N̞y9�"%u�Ģ.�6��""Bڂ���vn��^�'+���j�����4�_v��k:���Ϳk�͸w^�U&�_�V�sh��Pԣ�`�To7cె�1�^���}�ۚ��Y�!�+w0MtG�FN�#��qxJ����5p�y�Rw�%=8���Y�H�N��S}��'�/zZ����º�����i��"{o/������_3*�4�ubn��6�r7N������x6��(�:������O	{}���N��-t�S��ob�� ~�n\w�kk�A� ܣ~����1�g�	Y�.v�8P�t�h�������@[a�kw"�3���-N̴���0#�1C*��k�9gf�It������d1k��hF����Uҥq�̗�V��㋒���AU%[�~yN��r�4��e!2�=�uur�4�6▏r�L=��\��S~ᵍj����-�|���\�C��2���Z.:�h�� �wRZ�JjQn���|�0�n�4N�TxH��؋�NL��󂡘M"�㾢u*!��5`$r��pV�Tz
��=�%_:a6���d�r�&��2b�|9�˼�7ϳ��jY��;��E�|�2vl�����K�B�q֊7�Red�zz����y.�e�V#�.�Ν�ci�:���7��f�R\�.Z޸��p��?#P���Zǽ���$�y�LV������%��mf��faVNG&^��%�������6������.�N4ON3��<�V� ��GG1lm���Z:�c�x4��,�k��؊�2�e̲�1ܔG�;T��lK�#q�8\o/����\�%67�{˻�����Np�
��n���VdSs2� �#g�S�R�Ce�{g[�,<�WYj�v�o��^@hL[�[ȭ�{|����eb�V��.V�;�8�C��J����#���)���&��+��ɴ^K����pf�FM5��G�+��+*C�+/2�Ø�WCj�#�AH�6٠�*ѷ[���� l�����`X��L���&���>4uK��f�TCb��M�d>˜��x�~<l�zeuc�Dju�Yh0�Zk�[�]s(�jiH���OŽ�9f��.m������X�H���V`�F,���.�o>?]p��\{>dvs��]9q�v�t����*ިh��'3,��r­JZభpX�mdw���L}W֯�ٴ��r�_��;!}rP-Ce��=��X�I�٭j�]�ې.�0)�4��d"̹}�ҹ���v�;�통gXU�v��������Ք��.zѮ�l8��[Pt��N\Ǥ�]P
q����*]ʆ���a�cI�T�����@c���s�f��X�p��Y�)�}¡�=WZ�����[�RĞX���t�r��������vit���Rٜ[�|�Z��:5���n�m`�[U2���9y�p���Mbuh��%�v,V���_^:�[sQ�:SoV[��}ܣmv�3+��TR�ynl���ے�t�Z�yn�m�Μ\o���F�����\�I1��H�ŗstǜn8%##B��bSim����fiW��yS�R�hA�!�S{�13�O(f�uX���������b��>Vڔ�ݫ��ZhZ-����e�\p�.7L��2�kM5K�W1�����V#�Tu��j�--kX�)�r�6��%F%J*�n�k"��\�*��5.DM%Abj�ED���[[Z�b���ZZ��s.6��[rܹ�岴PQ(�Z�ٔ���Q-(*�\LĥfeMe1�W-*ȷ3���amD�(�b�b��ҊD�%a��%�Q���)Qa3.
[*m�b�]e1���j(*�JQTR
��kY����s1A%DU\lPY�q+2�@Z�d�q�c�0`�a(�XkҲTX:�TUTQƈi�J�&�m��[F�s1�Q���ne�X
�	
Ȇ}>�" 4�~�{�;�!WR;;��#2������ũ�:Z˦�x�+�KM�ؠ�#�N�����_q�{���r\Z���(��t*�vЋS�>�k�߱u��'�D�
���4�QV��t;uV��8\i����N���N7."�T�nr�b8�b��w�S�Yr(u��3�2�������Ў��qO��^�xN�#�j�:]̤j����}gfm�<���sz@�����ڷ��K���D$��Rf(>q�v��]��4�E,��I����#ƺ��=;�eQ��yT��[!���2EQ���M�5�����܌p��x�2(� �@���3^��A��-͘�����O:�{�gP��%��(-u]�-dgȬ�v���C��Cok.�C��gg9����1d��+a��h�59��j���4�k�K�R�m���{'m�/'��7�t-��{W�4�`܅��e���:�z��d������,�t]su��������i��o��Mv��:g	N�:{a�6"��ɮ2��<�
����u� ���V��Gl�m:DNݘQ��frT���t��2e�]��L��������d�NI^�^�#%V�����_7���<�>��ު
���{7�u.�3tv'�+��*�j���oaq���qʔ��E�u\�������'S"�"W3�Q�cw͎�p�n�2+^�kQ�☞V�Z��2fT�*w�_5޵�9��9�=�۰�1�]�h1��E�t<�^&��JQ��#=�������x�F�������w��ί6��69s�eRMOW�m�9}U��^4��o��k�z���g#������M�
��!_N�w�֥���e������b��%vp��@n6@�������$TT��_^A!^���5JT#oK���O6���oqW�K�ۙ9j�ަ���l�W�(�"_TaS��)�U���4Of
�� ś]��<}F�-��ڄˁ=��v1����K�u��5��LW���KZ���q�	qA-�z�S�����Ώ��t�.��fX���|��>G^��W%*-Ou��������c#��]�X��G�u�{���sD�nb������>tJ�)Ɋ|:�nF"��qе�8-C�꼱4�*�{��}TB�}ˣ+��v�&��u�:jo�K-	���<TUf\�L�5��q��@�؜{�ʫ�}u��1�;f�bY�0(r�Y�JH���������{���^��Dt�W��h�f�7(�}lG["w�$���\��aԢ���9�˼�=�g�޼�ԑ�\���W+`�"k��r����\�ε�/�/bxN��Q��M̝�uq��^XOz���8�=
�.O�q��Ə.��u��5'�5�ڲ�=X���BX�o��1�S�Bqu���G;�:���.�O��;+�o[ZD�l%)j�t�M�xWwU3��^OC���wۥb>��_�����MZ�� 험�(�+�Y[g���fQr�S�w�&R!wN�G�u�����i�<j��B�n�4-�o�3Yǫ����[������YTcɽK�VT�7�_~���b���F��^9���R�4�� ����*�+z�0�^�O.�U��<=�
֑Ɯ9�5�G(�k�.g�f�8�����}Ma�L�>W�׶c��A�kbV���Y��g�����/��2���H�~����;����T?g_=��#D��\uz��}��Oi��UH���o�*�+�`z��_՛O4hZo��:���~H/3�:���Sn��TWg��|��d�flڃ����=C�-m�,�}.�,�i"�*�=�aǀ��xlP*=�!�'�Xc!�'��+6ɴ{�*N�پd�:d�gsy����h��,��Eǆ�}���ۚ�Y�V�.Pm}�:=�ݷ�I����t��u�N�v�`u����;@��uް6ɴN��`M��*uϲ�톷�;N�La�������:�o���rz��Nw�%d�&�d��N�3�q��;��B|���`Ci���RL5��&�Lx������=�z`U����������߾r�{�l;�|d��&���L|a:���
���E���y|�M�/V���!�hc'���1�v�ӌ8���>�t����h!���Tz`y���d�9�!�'�>��>������:a:������"æC�<O3Y	�B�VC�NR���foU׺�ٗ~%���[���5Z7����M�F�]��*o�t,�����z��NmD�����;��/)m�M	�9Գ�:�z[4�2�DQ�8�IZo3oY�nm�z����jMU���AZ��N��WBo(�7�4�X��=�{�V�˴�u�c��������$����̜Bo�2m��l�7�Hz������I�'���>t�}��a�m��I�I�5���Оw��������y߯�:��=������m��'z�w��z�i��O��I��C����'6�|�q���I<d����HO^�I=M2g�W_w�;9�f�^u��{��Z��p�M�Y
ϐ�'�Y<;�|��6Ύ��&�l>|d�'G�$��!���XI���A�x�,S�q�� ��}���Sz{jZ���{����4���'�&��$�L�I�I�)��|ʓ���8ɿ)�<��d��:������6���C5ע @��G���/�eRS���3�ވ����v�q�������'�����x���$�T�V�Ì�0:;�m��N=��a6��4Y��I�9ǉ�}���N���C5?��������O�wϰ
�s���CI��hc'�,�Z�L/y+$���}�z����e�i8��ղm��OS_a�s﷮�7��ώ���>� �)�y@]xt��C��v�>Jé�d!������`k��C=Jì�>I�MK�J��W��tT{�X��*-qo�Y<��=�{�ۤ���t��2����k�a8�_o�N���	�+L� �OS����&0�}Cl+'̨T���z~����Z�֔fr�U��������q�kVM��lwa��x�;�Hm��4{E4�m&�~�2�7�I6�u�äht�:dĬ�5�s�.�8h�}w�7�Z�}��
ɦE��'���gI':5��ē��'W�������זChL�Qf$>@��%Co���ϼ�C�.U��y��e��\dژ�%,\X��s��=-"#�k���w[��vW��
�+�1_{z7X�k��c{�=r��)P�vHw@���]��'Be�BMP��fa��r����^�V��N;���fs]�� {�
[Ǚ|z�=��{�ߝT6$Ĭ�����R|���,2zɢ��� k9�u�$�i��;g�Y�IR��!N�!��`�w����sX��y�:�����=�2m+9�������@����&=�����a���ɷP���2���h�xi$��eՓ�bv�$�y�CO���G���ī�������|�/�= )*'��L풉�o�'��8ɷ���LB��|{̞}|H(i�p�3��M>�H)�w�V���4�S)18�~��b��RKہ�t�0
&��� 8�'+>۩O�7����
��aêm�H)�<f�I�
��}�!�N&$�u�0�= �^0����T=C�SOo��HW�w��>{ꐨw�{�t�I���* �L=G]� ��*�~������ l &��3���v�C�=La�tyLt�P8��3LĂ���Cl��!�:ߘzd�+�<&�æ�I���0�OYY��0��I�TI{�RqWq���{��3�> ǁ�:*G���!�J��^��d$52�Y�I�T�:�I�vN'f�� ��M�:�����Aa��:I��c'{̊|ɷq��j�Y�OW��k�w�[�9����퇌������$��=�7�L�ʟ'i1����ֳ��Mn����V|�d���2|ʛdۏ��1'�T�}���ACl���_��[�����a��~��k"���:H/I;}M'>�N _l:5���md�7�Ψm:C��xCi
ʇ�Ă��9a��
٫�aS��1��� �]�l�ɷ� (�}�*��w�s㷩�P$�32�Ğ��B��o"�L�O_�C��0�H)���4v� �;.��m�q���p�!�6�à�pIS7���1��z�>a�t��PG����<�T�Ɨ�O_���Ĭ_S��4���>N�t�=d��ez�o�:O�@�<��(V!��;��!�+�o4���<���'̩QIRq�����AC����y�g��7^��o�r�cz3]k�*c�b���M�yn�ON��,���+�[��6c��Ʒ���#�U��]�ְ+ӲL#Xf޹�V�ո$�f�.w�<��zLݴ�\��ξU�n_L�P��xÊe��f8L7�>��I:�޻�������>f8�S�,�t��l��'>q���i��@Q�X>�遶�[��4�T�s��:d��6�C����Xk�<öN�AIP�ߙ���J$��{�~�u���y�ε�}�o����VT�N]�*M�S^�9�I����M�:d���'O���)��|����8��yz���@���Ǥ���~�Iq�� (4��?|�+�W��"w8|¦ �Rrw�O�i�M�0�˦��_,
ɶT;5�O bM��f��Ls�������O_�O&��S�k�)Ǥ��a�>�N�yǲ*<�%l��ٳ'#w����������3��ô��î}���3��*q�3�1z5@�O�Ym�J��R>Ь풲|��tÌ*g�z��hi��i��v}O��ǽ?5k~���_Ωsxv�+�������d�UI�T�o���B�a�7��Oi���d��M3H=sz��I��c;Փ��8ì�;C�ځ��0P��06ײ�<J��LyjN��>]������8��=0i4�=��O���4Ι/()+��`�8�D:7�L�ʞ0�|�Ǵ���<�f��Myt�S�QI�2m����1 �$�SI6�}��϶��z��Ͼ�9}��4�Ł�Y�Or�i����mH)*gt�'R��L��h(T;�̇�a�8���x�1�,4y����c*}�v�N��1=�
f$�Ϭ��r���=��ڵ6~�֢����0=��dAH)�;�x�{H)�y݆�xΜ@����AC�8��l8�Ԃ�=��i3�:>���f!���`�=k'��A�0��J�ơ|��_����|���{zy��|: ��z`{嵱�c
�n��n�|�a�8����4��T:5a맦d����UI�=�Xi���;�OIZ�v�l�=�xi�Ƥ��3uG;޷�s��د�vw�ݪzw��p2=��	T2 b�I߿a�P��@�w���IP�J�e'l�'l��f�4��+&'�3L���t����%�(��������\ &�;迳������-�p>��`�Z0��e��0qS��IJxX�j�(��L�Tٛ�p��m�J��e|e+$�9���\��-��4��(�v�j���O�Qٕ��qNy;[#��6�Θ�IRU����w� ��ΐ}����������.��}��&;d��xs̓I��7��Ă���g0��|��{�y����̤��AI����M��1��8�h(W��a�8��{þ���O��9ǝy�|���,����d�:���W����sht�$��X^�*IY�kx|�� �����i� �Ϝ�H���8ì�󤂇�u�0��Z�DF5\	�0���ַ��s>���z���vLO�q�����X08�N'{�b���6נ�Y��>d�w��,�0���N�q
��;k���C�*w��6��Xt��M��G�s9��9�w�����ʕ���sR|�� ������O��$�
��Rm���t�Sl�8�;���:`q�w�`i>v�v{̋������tɌ��2�[�4x���B��������s���{�us�rk1����`q��'R�OYSW�'�& V�M�}���LCi+�'y=��_�A�S���C���u�O�b���b�x)� T|o*�� e�&~�y޽� �iy�!�&�Ru��M�L1>Agv�ma�/��1����H�0+&�̊���:��m
ϒx��T!���N�t=~� ���.�[���Z�b�|����}���m��;9�'�I�>��� �����*T>f3�X�a�1�*��Y<:�M1q%`o��I=B��J��l�8�B��CN�Qz����h�O�/}N�i
�i�.'h��4d��Yѭ�d��P�>æt���w����&���^�d�K�&َ3�Y1��Rjg��:H)�M{tÎ����S���Lb�A�-������@<* �ua�%C�w�,�ed�5��T�&$�:�쒺gL�t�z�,���Ѿ�t$M��oZ;dǤ�
�yg�i��.�|j��J퓜��޺l�/�s�IT��#��d(
|�ɜ�����8�!塤�<t��R
��VO�P��LLf�bm�oy:`cXz�Y̩�t�jw�a���
��|�g���3ns��{;OX�]�W�=�8j+��!���ρ�IE&(]��ǟ:K_u[�1w���L�q���e2��V���Ú���m6#'+2à{Gu('�7���ʱ�J'6,�eE �x�r;�G������5-\٢������1���4��+=I㝚�D4��+:�����'gT1<a�q�g���I��y@ۤ���ΰ8�0�R?P�J���s�� �0񘜮Ɗ�]�g1�g�z�@ ��O�<f1|IY:���LB��F�6���:��$����פ�Cht���ü!����z�ىP*N�:���M�q�{Ͻ߻3�4`�����yn����z�������`VmC�ϰ�����Ϸ�׶}C��@QC����� t��y��&�Y3�1<N�bO��w���Y�$��*�x��8qO�/���ۣ6�߼�}��!ؐY:xyM'l����z>�D��l����s$�I]��z÷�
P�i�'�I���w�e'�1C�a�R�'Z���`tj�c�Q逃�B��"�U޾.�g��z��l1>g<���k���i8�$���AH�`Vzo���I^>��ߙ�|�g�;�3�~��WϳR|�T�λ�I����$�� 0=����~���w{�D˘��^MY��L8��;<��R��:�$��ӹ���HcmN��3L_Vs�zI�+6��;��'Xz��5�y@�'�Vxo�|�Ӥ
��o|��s�<��q���A`zצE*Ad���a>eJ�Y����&Ҹ�����7��g~u�$�>���:H)����oL8��2wy��E��9��Ơz�<�!ϭ[ۻv������{c���ǇޥCbt�N�bO_Y�Ι/Y��I��gZ�I� ��S�i6��*)>B�7���偈m%~gGt8��� yL��{�@1�+K��_Q���������o��Ob��d\Hwhp����;`q��vbLB�m�0��g�1:�04���:��'bv�
E��|;�6�!�J���H�� LyG�\=v~���%}4&����&#�N�<�*C�׸t�R|�T����
|�i�;��M& T�9��;{`t�f��C�i1��Z��m*�+1 ��=�y:C��1����d�eb������:�n�÷�.�+|���QZ��uc�&���d;�<�6�yR��R��*I��ѽ᧩�����R�ٜ��2 $C=�{W#���2,J�p�uv\�^��'"g^��{ol��+�5l^*%��o��%� *�Y5��R��]��=�xy^n&y<�_�x���+=O��2m�����)�I�.����'+>��x����� �|�o�:T�ʕ�����VOR��sT���>�N�=�]$]��ڜ��y��>�I�bAN�w�|��o�b�a�H
(v��̳L���(q%d�+=�����N�c����k1�n�ꂒ�>k�öL4u���c'�&!�=u�k�k�v�]s�|��I1
�d�~�]$=I^��$ۏI��1�&>&�:<�h������ڐ���SHcma���HVM�7�R
m�0ε����mg}#��w}����<�滼>a�i1&0�ف�PR.�:��ɶT>I^�����B���p�={HT>O;��q&?j����AObq�׶'*��q���bU� T�
���q��-js>ի��|� �z�9�a�:f$��<gHi1d�=��Leb����'�Vxg�&�>eaֹ��w�m<;��z��'+߶m&���LH):��z��}�ֹ�8>��z�4ʕ���b�&Ҹ�{@�1'�C��a�;{H,��0�1혐��kEd�|��'sVM�@QC��<�Vځ�]�8��m�����i<N�c5��o�2��8�^oo���x���t5�%@�/N��J$���<gI�N8��7��&!S�:��<���P����O��
z]��;}M!�Rbq�I��k"��R�_yr�ͼ���aKx)����G�Q0>� THV'�Ă�3�y�t�AB�=oA�Cl4�LI�甝�AH�ON}}}��55�Y���L�T����[������X�GA�'b��M��E梦HX�����lXOƚ<m�©��g)�Ju;[���R�\lh�B�;C�u���@�$r$c���r�� �޼y��u�]s�betY��LC�E�,�_��qTXލ�T��p�rc4���١��-�2;�q�c>���)�#�p-�7w���Wl�N�\X������lm��i�9M���N���WNWE77ttTyJ�%.e��s��	[BI9�.P�#N�2	gwnLR(6u�-˺�u<��]�e�t��wA8�=��4�+�*�α����O��a
��h��*xGt�e�e�t��7���͵ۛ��`�iM��}�H�ʻi��-P�Wd�/��w�BH7!䠥�����N�N�l3�U��Ŝ;�n��6P���O��]ݤ_*�2���:�m6>5+(bй6p^O��੄�:�gz)2�e.9ni�ڽ��N��eu
r���3��W���n�:������VX�;R
�0Ѵ��eb,��qE�<Ww;�7�����<���#�U��u3Y�_N�t&�:Y�A����f�@G&���Ru�}��	YĒ�����CV�WEU�6�{tf*s����i�Of>h�"栜5��U���,WKF�q�ZyŷK7zXW ��U#Q1u��K��|�6�Cb�h��3����=���0�鬛S0d�C��C�4
�xw�� �xoP���ѡ���5:N������e�V厸��k��w�>b���FWQ=����Y��q�,.�}:>�Vm���o�a�������L��Co����Ӌм��,��ƑJĮ�4^]]���H����+�2�J���V��`Ɲֻ������gCX���C��cY���wJ�oI@Cة����Tч���4��T ֏C�lSh��'m#�-q�p�Cf�彲/j].pG��k��AF�(���U�6���镲]ԃU*��:Q�fr9G�XH;9��y��A|�&.Y��8���k�z]�bvΕ�톊o7����,�g^ڵl���VeGt��rd/-V�ø��'��[�_c���_fu'F��gq=]/:���&p����8y���-�m^Bww/,�6̏�V�ڙ�j��\���9��=1^��=Y�iu��v�0�E���ˉKem$q��Z��X&�A�	p�ܙ�ʼ��'������O:`������ܛwY��4Ǖ(+�ޏn�Ʌ�O\�&�\���_��k.;�;��%�csox:Dx�	�Y��� 3��0��/.����"��Tq�xp�[�-��"S�-ر�����t�`V�q@��i�FA����q)�c���m՗t/N�&��E[�Y��gXgr����#�<W��оC�me�˄�K)KZ�[qۑc�Nq�(jJK�Z;�����s��Dవ�Mwcc"��rGNlc0n]�%`�>VJϳ2�VV"
�q���²�E"��Z�F8�LY��8[i���̭��$X�`�ڲ�KB�"�Q-��*L����ؕ*[ET@XԂ�e\��Z��*,�(��C��[���kB�e�8����L�$�QVUJȣ���4R�XT��l1�"�d+jQR��)X,V�3T�`�`���Z�J�DJܸ�%q"�X-Ɠ+E��Z�%q����E�@ƥZҰ3(
>�MaJ��+KbȢ�%E�+X#*��V�6�!�7Z[c�s��U���+Z��1�8�8©i*��ܷ(�Z[q�r�S�#�)�~B�$R�(�%X��\���[!�_Gҡ=)��[(��v��>��!A��މ&��נ��n_�P*�V*�ŋ�����x;'{�=u��{�櫓}�ֆߑ�f�#�9j�P�Jo�k�ߥl��LI��{81��v���=u�C���(�XQ���t`��9R���~��ϥ����kv��p���;�&j�g��!Oz��>�T��	�.�R�G���=Y�[֥m���G��S,c�/�N:�aF�L��1�Ͻ������Z�����5������r��~�����̂'��lL���N=W����w]
��
+�,Ќp�Bth���O�gsK�HUA�	=��.�T\��L���
eԴ����Dt�|������{|߹���}G���2ر/���Q^��U����6�=��C��^U�7tۅ�����r��w%�v!;h�CG��_��C%��ƣ�aھX�����]և�S�����m�u�n.�']�$M{��=�>��G�
vxqQPɷ�2����qx$��,i����mv�-��A����j��OE����{t�W�2�"��V�-�.�Ѭ9�8
W�3�\]z���t	I��)F�+�\o��^�X�q]Sl Ԉ�*��>�k;�/o���A��$b�Hk��.�t��:���v�(��}ȢMm�(��w�xI�^�a��0���gl-����b\���lt}J:���o�(C�����c���B)U�@C�[VNZya-�~�������Įu��|:����/ez�g�8=B�rs'ܫ�����8�����q\Z�]���!}�Ax^��pt�1��nve��xe� >�5�vh������n�:j�+<�Qs���2Ŕ�o�h�u���ФlH��T��9�;����R�꧊,��,{��R���W��4։|���ph�P�����V�{M���j�v�s�\
�(y7��}.8Υٞ�����.8ɞ��i��;�VS֭�2p@���b�t�J�~
��]���A�q�T��Ł)����4�&=͕�zۯU��͆�*�1��%��B�6����S�OFp|f29�,������a��"Ł��P�Ϯ[4��$#��h�jw��>~�WwZGU�6VF|�=���gK�����v�<8?��
��F�z0�m��K����6�;6�������P n΢�����٠س>"�"���`�+���y�j��4�	�4��n����Z�T�Mϱ���~C&=�_D3�A�S�z��iu���"u1Fͨ�0��H�b�2v�y�d�Q�b�7}�� =֓�׍�����:�g��]+ۑP�@�H�;�/#����^�7x���כ}��螮�Ýr�:��E?��o(�����1�TLz���km�f�i`��p��(��mA��5j��J'�
�L�ٮڨl���u����ĕ{�V|Eu�]E�ҩ��N��@�
���*��K�̢��=�]��5mⲸL9���(�f|�x?�L���|	*��,�#�C�Byb��m�;F�4O����j�u3(|��7�Ù��`��r�ԴB����x̺�{��\V��X�����]Y�.�;���ν��8A��V���d���^�<ۉ�Q�u{(*�3f��7J�W��_��U;��5(A��,o��{�[�_�V����~�}��w�=�u<�^T��������n�	�V���ak�1杫���ZvT�5�[ǄX�P�r��Q�EƆ�p�;.6%u�\�K>Z(+4���G�f�\@�[y!g}~ڻ�	��H�xGR#� ��1;�X�bR5�]��TwSx�~�jL����=��]��e ��N��RY\�h��r��_<z{���z��/]o
����S��a��>��c��K�}��>��g�m6�����:(@����Ѱ�I<�X�C��HZ����^,�x���)�<�,�mcS����η�6.f�pa������i�&�h�Z��E��v]��}=��"c�|�%v��2�=ڈ{"��+ ��[��S@\P5���y�.����ƞ\l���J)!'���j�cc�gaYer��G.��D/_H��/#�%�
������C%$`�z;Zd���P�Ӎ��Ј��<ϳ���[�a��T@g��H�^RNٿ<O���e��{
�1��E��W���vg[�e.r���~r�N}��Y\m*+�Oݙ��z�%�#l��yI��#%CوPc�J
y�:�K�A��%ō5�p�c��H�Է�8Yi�<>���mp�yo�������T��P�>�
���y�=����|�ҽ�7EN���X.�c�mhk�Y먳��9}`��W\�$��o��fA�k���]S���\ ,�g�'l�?;68%���t�"m���v��IDD6�rI�K����t1
A)3��VJ(��YW��ꌢ�s��g�[�w��@�n���Q6{
��E���oaR��]Y�n�|-�r��)fV�B�
Fg^�:U�i����������f�ti��hu�����=F��Г=F�Oٵ�'k�mJ�5t���FcHם�����(9=2���zF�U��s��5u|��Cc�GC3�b梏P�c����9S�/0��Y�YΚ�սf0sOu�Z�&&i^�eD�������A�df�S*��av�V�9E�7��ur�3�^G/�R�٦U�5������5H�ו���![ǕP�*�@vUV6�@ؠ�e��{�d��gUl��%���hl�X�%a`uyDK��m�w*nW�c�T��m��y��P[(V��:��,w�T����R�u#9�OP�XP�]J���K�s^w������p�ߦ4'Pve��{ݕ��$eb��Dڢ��ozs[��=���tH��b�rg��#��|f)�7jGDv�I��W�Y6&��[p�;�Q#�(��
x�	������TX+K�oB����R7�K'�C�ʿQ�r�l��}�B�u�j�A�43��RҲ]����kk<�ݎ�G�}kS�")vfgk�#˵��'����{yp�L6���?n���^��R$
��N'J�X��F�8��ǋ��};���T7�YW��u�KטQR��Ŏ�;�>Y:<�����eb��� ���m���^�{:���$E�hi�p���,^G�E���[H��ͥ�/C_O|ܢ�
~'_Y�g��^���&�h�:K���,pt0X{��N���j.⎳<�X���3	�2�_�]��m�i׺�Y������5=>֔��_��cC�^��cLm	U�
�$K��r_�VVP��T��y+�MY0�k��Z*ƪ�ˣ�
�f�(�R���	^68x��B*�X"/|�sp��g=ǼͭU���T仉P��O����j�9�@�.f�*�.y�Qqu��g�Ea�M�@ҹeb�Yܽ�貨z��� 8P�nUD�+�N�{�n��!��nsu)+ v�p�{����<WԽ��mN��	F(.RoC����^X<+�]�)Jx��ޤQ�ct��U�h_�:W��r��Bi�LS�2����%�p{V]�c:y栧r�ec:�+������&�h���p�O�.���-Uc�K�3����P2�l8Zv8��1�@�g Z�c�C���%�*�5�]dz�[��T�	�j[������;�TۡzQ�q�q�ۧ�q�2�Yw�o
�y�P]�&4�_+u,*�v#�ǻG>^X�8�D�SY������Rԓl��9���W_�cx?�w�J�j��=����7n:e���׽3�Ȭ(�=��V��=P�R�`	yAO#�62\,�a������Sz�;QW�;�pYk=�fn���]��@x����!�HGW��7�X��k�<c9w���HyԢ�Od����R���������h�V<�^Kd'����"/(a��Sܷ.{V�"�jt2��N�.}�B���R�L�R��]	�Wd:|5���ܳ�8T���|=Ƹ!Թh���[��4��|LGA�l3��8�k�o�r�����4,�����И�r
4�|��Uɘ'n�'oq0dͤ�����E���6?�-�+��5������[�K��gޤx�f^s�5{���^��t8=�%D*�F��^d�џ/L�)��)g����Z��Ħ�d�G����W�>ܔl���"u���=H��D��x�;b���*.̎hB皬�O�k�}ƶ�uT6����Qq����W�c����$�7n���E��*
y~'I�7�[م?y���ψ͇1����.`";ְ���S�x�7x�-�:M]�A=T�5N=��r��a��}U�R��K�X��jh3��>&�
�2R�����������Ep�{�iC{�VQ{���t��Fm��fϭ���`���V��Gqzk/�����/ǹ+��&�%�D�=���2���;�й���=���n{�m[�̦�|�lGrmﺉه"��QC�*Y��,p��#��FT^��p���`��:��Uw]���z�>�͍�ثCt`_i�	��r�uA��+���BtgN�9l���I�+ׯz�l],*.VgT���=KC^_#���TkG�ԫ<5�_�K��qbD�hGg�Fj��*�{"���>O�<.�"9�v�n����]_h�y<zǽ�f�r[���(R��:��3�`p7����x��'.�S*#"G1�5ֹE�~�����u�p;K�������~^���
��t@g��gt���m�0�jX�*��H��lßϊ�/;Bz.9CB��(_�V_��>�$�[܃����o�[>��QOeXm/VPǂ�ΗЭ&�]�di	W^�a�~��p��H�U�Y��u�>Q��ofE�	{W��r�@`������k�yrV�:C��i0n�dB��0夣��b����V&�����H���IxmcU�o��gM����2��Y��K��\���;���Y)؞Q�]q��_��hf쨳�v8˞�#%��p��;v�'����׿�P��nT��[����!�S����Ԉ��Y����a�3ޠ��a?c��;�E�,�3*]�E��uTxw�J�g<A9���f� 3=n�d����k��Ph��p�债��
����3��#^v
�����Q��w*�ｳ�%��w�*�*[<%B�~B݆X���T�K�>m�Fh�s��-�FZx'B{�;o�н���ZӃXJ���Qɠ�]H�T�PX����3k����y��@��r��U�ɭz8Ÿī�V�nV|S��7<҂|���w-����oa�&��r�q�>"V�b�����F��b���Z�)ã��mC�:�����\�䕻,S�,�ڽt��!ƚ]aE��`n��U��r�g�m\��&�yW� �^����& ^3d��cV��e�*�]s��0T���[�Ϋe�VEp]��[5�h:x}���M�m�-Z��Q��*���x�j���TZ1��Y���\3�&�%�M��):mt�A����[��\g�磌�<PI�{RĮ�|�vK�:�ʿL���B��g:�aR�Q�H3���8�����r(�s)�����L߱S��*8�B�93�C�u>3��C����%���q��\#4�zd*�����y�iq�9�E��.��ʠ�B������-�����ܺ�n�v�cSC��@S��j_��*f8�:K�)��[���v�U������24�+�ʅ�
�/#��9�m({�a�ܝ��'�ך�l��4Y�ʹq��{7N�;52@��3�$SZ C�`�|'�� �;��{��˰x��/#��^h��H��_���3 ��Y�y��B�u�qw<អK�=���=:<,hS��V�b(m��>�E���=|V+U���0��$���O�"�"����z:�N��(p��vQB/�r9����Z�w��Q@�^�Vg�������?�~��Q[,Z��lC'ک�̀?X����oJ9q�nP3�T^ቍ�j�Von.��xԫ��;���Q�yK׬ �w\#yڮ
�<-��P5f���N����z\�k�����;�"%�Qt��`{Tŋ)��Rr�|�(!��9Q2k���;�ׅ�fd��?��5���_LL�Q��:sd�KxU���K-V���C*�Z���tƄ�@co^��u�_:�z��ۢ���gR9�u*�lDsifa,�7)����^V:[�Ñ�P����3�]c�!�����v�E�]s��p�0�ݼ��6�5z��:�ؾ��C\�l���yC3H\��pӒ���C ��8%�*���  ��m�s�Tx�Y>��ơ;�w�Ȳ�R5�M30Ng���b.l���%����W@Y��.v��&��V��98�`�\�-��ۮ,��B����]�̩sfr^a��gT�9C�Kj>�9Q(7t /�s�Ha�����Ma��SgknBr��Nu�2��|���gǦ�*��!�ӏ���n��L7X���`T;sft��	
��ƪ"�mX�b�j�N�/Qxk!IaV����x�̱��=�@��H�B�J%��Z{ae7ady�fcI�"��.���K+m_�����;76n�2�I�tu�:���+Q�CWIh���S�vJ����K��c]	�+�b�NVR2����r��Yo@���Oy&�񻕕9q�֗��C�c��J��X��s�O]jՖ��X��Z^;׀ea�M�����/�7���0.Ԓ̗%4�d�P�ـ_F���bK]���룴$�kw�E�^ǰ�1�>6�U�K�vCY�d-f��h�::�OG�.�l�R��ۤ]�F��;a׿AϫR,1��:��:o���1�W@rhMe���=�Γ�L�m��}rjU��;Z��[�^]X�BI	�ѐ����rrX�;P��Jo��u##F�n�.t\�e
�Z-WC37󗣨�C�n$�p`����,Z�r
R�i�-�G6u������֗�'fbg3d�w�f��V7�R��;��޲쑎���r��[Ӡ�cN0�O��{����U��gE���� k��՝��:��Y�A .�����֊�]W����.���7ِ�G���1�Ir݄d��=g$����$G�^�F�o���W�'Z�G���0�zq}�O�eo7��U�tm���.��71]6�L�ܱ�+Zw����	X�&���}a�����x��{n�ulGU�ٰ�Q�{�r>�LW}��ɽ3�AG4�Y�$�ˎ�V4�J�b�Y˄�$����al.<���I�k���;���5�����P�+�>�
�`��ʦfd�"6�IZ+�!X��RV6�0���h�L��dR�CeT�,1Y�T`�"��J�`�X��*�9���YRĴ*�U\��Њ�5Z� ډQ���Ũ�
[J�lJ�B��J���U���$W
Tm,B)m�q��UB�DKH����er��+r�Re���Rڥ@U�V���ʹAcE��˙X�+md��$���Զ�qrŪ�DUeFڅTQ��L-T�,�%-����L\�q��q�rو�Vԩ����er¥V��.F���`Qne@��LaU����̥jT1&e�-K[m"�C�3���p��r�E��[E1�d�*�,\QPr��-ʩ�����]������~�ι�_��g���휤겫�N�3m��L��9�jJ�J�<��T;"�rg
�Ye����+G��U��D!���S_?��V�S�;�h?��ȼ��/L�j�p�0حs2��m?]�x�xvoO%�%ΝG���������2���<�Qu:�'�(.&�5����D��;n�}�����{�R&2����Δ���ƺ�b\o
w�Q�����0�d2�[#��M�쉋�B:P��@�ҡ����h���_�mdd��)�OU���&�2(Lr�5kG��@䫠�m@�1߽S)\�6���%�����P�;cZ�[����4W�
T,����Gy�7��I�ń�r�ׁ�w]9YY��D����7��CNˎ�q0�
;O�V�"Q���]����s1Si��6���b8�Ν���S��PyUQk�0:�.]����b����ۜ�"���+�q���:�q{�*��`���z*��ۑPN@i$v�6��u��=����9D?|֎xh�
�o���Uʸ0x�:�>�v��7��k0Q�9dӳ,K��by��$:8�G�^Kӥ���z�yu��ۈ� -�"��2�-�hؖ�l�	�
�E�n�Y\[������*D����Tr�mfم��T���i��}dm[-)��wi��2���ɱT�p8Ɍ��� udso�*&>č�t��r#&�:�w�
.��ʍ蚄5PQ�"|��^-��}�4�9�z�Ìp��"�U�t6?��e���ҩ��N�����@��f<r��k��8f9�E�ȰҢgR#d+�Y8tg��%Jf��Y�38�B��(�����\��#�t�4q�v�6_z�B�Au��F0xh����K�f�,�(;�c1�9����`�P]DR5�&ڭr�pB��C튾��__܂�κ�rY����憫�)+��D�Wc���F������ �z����B���|q�i�ii��p�� �����y�R��i���º�fv���PW�C�gcy7{U���k�r$$�����L���@u� X�e�
a#��FT^�6���a�ݺ�Z]�u�
v��z?F:�hn��h������ҭ��z�ڙ�CǊ�s;WBG7^���<�g��v�b�VB����
�3º:�������9�Z�1me�y"�����z�i{x%æ�Aû�oe@W>��'�s!���I�ty`d�
�5e	z�����8�y}-7]Ҍ��r��{r���פ5ի7u�7O��QeIç����i$5-����U_Wj\2#&{�[��¢x`�y#����[��L#萺L୉�s w{���a-�f���u�K\*Z���`��P�>��a�LPx��_��R����(��p˕~���}����r�<��.�6/%C>��*��n3�𨛗�&"�܅x2�6�R4hıSzY��K��]*c����x;5����z�p7�x������Zv�3��k]A�|:�R��֒O��������i���.��U�.E��X�F�y��Β[�	P7$���
���K�t�n>�[����g�>Vf�7���̓Eٽ���Q�0�U\�\�a�����D��Ԉ��U���<F���˔�ۣy�e���D?:�W ��[�# �Sǻ����`2;&}���ۯg�D���[�c�vo��V7�Ei� 5t���Ɵk��I�VW��t�3�@���%.^'�.|U`UB���r*+ǨZ�b6*s/.���=��#~�`���,��v�wu��&�]B��+��Q�pN�!����j��xZ�+�d��J��|v�Ւe'tR&Bq��wī�0w�9)K�p��~l�˂j:�C�;xG�����f���G�^1�BF�����J;��ev��g]5�������ݝ!A�%G�ʸ�$6����F��z5~��įx^�����6n>�#�Y�z�����c_#���c�H���,�6S~V�?y�w�S������%��*C6����G�>u�i�N�d�Г �q�|w=o��B�����]y���O�u�%aFv07@�)��|{����k�fL�_�=��}^D]��WL���1
{Ճ�{a�A�J�E�D�7i�g+Ƃ��&_��^����WL�*p2�q���PG&y~�p>��zn_xk��?�`�z�.�����`U߭�?�4���x�
�r�@����<:���͸��@`��5A��C�Ѷ-��iuҢ�b�xp��K׽R�M]}�5�h�}f�u��{���V��a\>B�p;.�`[3�!jVh�n�[���9S<:�>E\��/&Y������s=3�/-�X�6�k��a�x�\2u�cck6��Qk��:�����YY��%4�0õn�R�2���d�w4��m^=kȱT�<��gd�%��-a�إ{�N6��\J���2wq��W�X3�$�%n�Z�d�x���	�����UV����}����`V�W��}��V�)Vb"���ᒹ�+��驐Z���}9C�nMZ/����si�>=��K>���8�J.�Ckz)G�]S|�]Ú�����7ԷBAZ��U���1p��u�Y����2�(��!C�
��ͨ�%5��ɾ"�z��e�g:��hxl���u��u�M��1�
�� ��t&�Y��ap�<yU����C���?u�/,/�)j��&+���*��3�T�qG��N�Q��h���s4������n�h��U���Ю�P\�ގ��w�O٣o�B;:�y]@�{Ș���[B�<����}!4��֘�|e��_*�I��_m]A��w�=�s�����;C:T44��@W*�m��nl���a�-c9?@�o�1��~�.h��q�(@5*ɹ�*��T5#aGm#�,b�6L^����O��O]��S;:;�
uǅ!`	w�����+äU�z{��VX��͊X�G��.GJ�.�����L��EevP��C^�����z��ZS{�]�C֪7v��Z�`vm�Tp%��c70fӫdIͻf<���5�k(L�J�묩�=�zm�����[!��Y��g�h]�-��+c
<��������;��o`�?�tS���b�7eDB��D��"E+Ϫ���3����r�bP�����륋˖ԫ�CoB��>�&}���J�p.����U�vR��S�ϕ�p�J�s�Ut"��Ɩ)죞:���9�_AWlq�=ި��מ��}~�PA�ϕ�֋Ǝ!\-�/q�Z�Z)�l���5��K_�hBZ�����iwkG��m��x��hY�6+¸;!Y�1�ƸULO?#N��c�YJ0�uN�f��Z�>5|1U#�J�x�ɪ�O�_+���sC�F�Lo&�=�CD�G�c����Q�Ԉ�
�NK�'ҙ��|	'�0ܬ΋=�ysfop����Έ
�=��'%;&�!䌍bf64L���A���9�Z�r}�D�9�����j
_f []�����U�d�+{"�<l}xG�2���!�T��H�i�}�'jŷ�ίeQŒz�}Z�(JOO�c��Bf�y}u���K�V[\�䙙���8���IX�Q$�`h��o�0F[U.��S��T�$��s𤋜9~"�8��*�zz���8��W����qk&�Wu��VS<w#=۽��Ж��  'n�;�[;�����h\\�������S�N��&ia������D�T���qʽ��V3;`uy@�|T=Vv5��x�����ͧ�3Ws�/��W�*9��P*��"�B��C��FT^�Mef��x��iSe����ߧg�_}�n`�g�ثCt�� *;���{p�8���QUl���vr��^͍b�{+�<0O�+%����.:;KC^UJ���e�Ϥ�^ep��/۽K]h��c'���m���-걊�ȱ�VBn���L�r����J�C}�����0���f

:�ð�S�AǷ����ً	өB�˝j�Mk�#]!��V�ؗ
��Z0X��5xx7����z�<>ԋ�fh������X���u�|���8�r�k���0�}{biE�m���d�X�'j6���Wk/�kr�
�j���洙Ip�2:�����j���O
�^�˧�_U���c8ntnH�O��<�J�QaU�K���C�|4k������u�o��h�3�(�9���ب�U|�&�
�F�]��$�T�����,�꫰�o-�tV�yk��I��)@�cn�vS��9�0�||@�\�@��q�&�D;o��󎖬-X��Ęae�'Ȩ��R���Te�F���9�_5� =�q�\�b|f=Suq��g���R��y}c>�l׸D��Q"��5�_Z:칯��33ώ�n�	��6~�Ի��bTxߧ�w��������=����x;�_A�R��p�;W�lIk�V�Pks83u�`�'B }������y�W��z���6YU�-�A|�T�����ĺ�����O
�p<^,�	���1�Y[�!�Vx�h[R�쿏�dg�`�����;��/5�ڋ���gcb��63ֵ�֖�5�8�@~V;Τz���X�%}������ٴ�l)��}<���%����Ce�#a�,���z�R��vAyN��=�:�"㿽�ߺr��B���ڿk�=U��q��XQr��
Ͻ�����vK:"��l�b���o�����p�mS�!:�����+<���h��+�D�	��zpǼph����/��P�=&��T߭p�Q`�z��o�n�Ӹ���\��������<���;V�s5�|���lؤ�����˸�#���𝽁:k8���k�,�0�ܰR�8���Wu����qN�����6�}`�g�sF���|{:�,�&��a������c\�2;����-)�~>�x��Y�TX�w�ǭѱH��X���x��.=@�
�3�0ҽW|�Y@Ǿ̷���������>�UDhm����ʈ�L�p�igf�;a{9׃�{Y=�f�u���AS�di��z�d��SA�
a�r�\7���s)�l-����G"�\S��½)��icG��Z��Q�/a�$����? �!\0Vz��6]��}5pZP�X�]K�oe����%��*w�h�*����y���VH�E���Գ��+G
�h���!uLd�	c�0���'$gv�:H�%��æ����4*VTG��p��z:���P��1h��|�����O��h��]��y�%M���E{���zڳ+=H���q�*2���3jE�BB仉�L��]�X�j��m�6����ҵk�صF˯tDL��0������M���٘3|;�Ǟ΂��!ʭ��':*�����5����#�:��2ņ�ew.�i³Ůä����~�N�AD}�$ޕ{�ډ�o�����m�.�x���\C���o�gU�K�NC�v���_[<$�����v��j~�T!l@V���7���ܐuu����B�FHL6b�}U�Ww�EH=�7�Ûo�+wF��Nn��Y費�����-�HM#C֘�el���'���g�� �ܱ7^�T�czX�Υƒ��K���!�ۖq��%桧N��7�"@1�]X����&z�XP�0����)W�%CR6v�=�e���&n�����E	�ݞO�G��\8U�,��={Z�^�NTc'����O��G��܄vm(ams�O@���AM�ɗĨ�H�f.z�e
�5��m�&=����1��Һ��<����S���y��NUOzt)إF���_�	�.z)]o�;�����*�2��ҧS�.�fW���4#mP��1P��{~�����c���� �nµ���SX,S<&�^R���\k�mև�w5Pw2���m�K���,W���b5�ZU���<�f��X�J5�a�1�[갯<�Pt�^�o���~�@�rf�/S5�Sz:��F\��j�*�<@���a�Y�(�ۅì�M��e��^=�����)p�x��k��|0���h'#pTy�9���i�Oi�p�"�|�e2.�[K9ʴ����e��D���kN<6J.��7����ú�$8���1�Wa�s���4GTL�-t��N�i)M�[��0����|�]"�k't�<��nc�&v�v���/���+��Ô���M)řM,���GC{��K��JT��WN4�\f�ۻ��mi���^^�[x/��t�f�aE@�Ԓvnn�8h]<�UsI����t����l��ѽ(�7 ��	琇6��S:Kw�C�s
���n�3���%yW�z�9�2�Cz�F�2ɬ�i�Vq}[eأY����#-fx�ڊ\k!Ȩ1l�enq��"���{4ڨ��wc�Mi��M<�]��We�t�3����9�n��[f�8Լ�fn�W8��#k[�p:]��S.�ܴl�v�����b�d�S�e=�[�1�]�7|%�L;��s颟 �$��P8C�����F��1H�]�.�u�oA�.�ťH�O{u��A��Ҳn���zŜ�DK�eu��Gt�p1��eD�ˮ��g�]6�u��iڗ:�N�K�8h��ݝHN+*6�c�pm�
��$:��rL�3�G���V���i�h�r���LWycw�ɂ�R�=(<(C�0�����C�<���f@Y�;:%��K f�G�X+{h8�A+Pv��Ϝ V⬨��z��}n+����a�f��ۃ���̔9��#X.�W�F�yx�r��JO4���B�2�nZyXz�/�e'y�~��f�]�[�+�z�x���V�,	qh��&�7�X�h�w�F_6���ա��|�@~��q���]��s�]f����X&�o�Z�7Kj��R��i�겳q��ޔ�
V�v:%��9�b�������*�e��Ծ��\{w�yk�[�����WE/5`�d�[j���O&G�X"��)�����Y��֋�(��ZU4*�u�t����p���Ԁǖ�q&3�t���X5>�yst��gSx���t�8a���˖)ݷc&,����vjb�'X�������1�w�MM7�z��	�U^�į��)�k�\��U|���'�?��"k窲��f�\b)%]�y�"k_	�ܺ�=���)V��!F2�-%�oV+< eע
��B4*.�t/u�9@wC����8_R�F�18Q�ΐH�|�m����B�j��H��)�F�d�r	'c"q�i9�\�\nd��z]��`�w�ʥ���98'��ҦVϰ���cEf ��s.�e�aFeU+1���e�.%E1�ۅ4��˙12�cr�lmS�ʕ��\L���!R��V�B��.8���˃�UC"�b������R�\s(�Z��)P�A�+�\f$m+\[`��Aakm�ne2�1�JR�d�+PiE�Cb�Q��f\@�a�a�֭�s3Ʋ1 ��j�5�f9hW�P�1��R�s2�V
(�J���,r�q�eL̰��S+hֈ��R�8[je̪eZ�����\���q�"6��`�-����ђ��ffn���Q���2��e�V)��LAC��T�ڢUe`����J"�LAT��V���+Rѵ2�eZʈ*եVȎ5�F.XV���-�72ʹ�FZ�TQ[jZ�i*%�b���!R��a��*TJ��!Z�Z�U���؆Z��@#"���3%f5��bX�U#���y�j���]|���C9-o����b���i��x,[��v\�����C`��!jT��b��:�O~�ԛZ�����v�T�21�χDU�z���š�L�!s���򺝙���{��I�dT������������m
�5}��FD��"�çM��-{�D������o���S;�G|�ߏ��u��N�&w�����{o�J�6K}�E��K��*�.V����d;��$����:��\�s\K�Y�u&.{o���mn�U�hٯ| ��ɿHV[�g�41����}.�s�~_[���`y�vE+�Sܭ�a<���e�`�E�g�P�\=��Z��n�(�Gx��e�^����Æe�Gz�<��?v�4���_���wt�z����D�Af��^\���U�{�����Y���+�ɗJ�_�aFuJ����@�@bX�w��'%�^�F�3R�`�vU��-���W����&�|��q�yQB�I�T%mؒt�����!U::����@�=�(ں��
/�~���$ez�FV���[p"��uDm%�9�.1=�r��÷�R�4��w,^U��Ue��vd��%��X[j��!b;�J�^1s���F�!�VH�T�I ���C�����%f���*��WZ��R�R}�S��^v��&�1(X�3V~ <=�C����qF���\��?='Ғ�ǖ�8{D��P|V�q���D��)�c	+�=ܶޱ�x��=���g��G�.Z�s��8|��(��Y�W���lR�O�;�׫�Ap���M޷}p���1��Ip�2:�)���:m;<=�{�v$��A\�G�J6�1�Ӄ��w*�y��u�4O��� �����Ȱj�^W�{ف���p�=��^��N��h�Qc�������d;
p���詁plX����s:�39�*̡��:�!�H;�^�`���2���Z-��B�.�aND��¸7'�I�w�jFJ95gԼ����h�P�v�`/��p�~X[�ƌƆ����؋w���=K����b���@k�| �tJ��UOUE~e���.d^	UHm>*j�3R�:����l���_�O���Z�ܴ-�`�H���^C���Oկ��7�1�t�!���j�}���W��^��Ÿ�5`ڵ��ټּ{V¶��Y���D�$�w�yX�s��ߍu��wv:jg�Q<TI:\����ir�r�;XC[��^[esY��Y]˰�p�N�ܥ�`�l���ե���VJ��5c}��Y�k����ujx�8f�ۊ$�=��,��_��+tf�l����U@{%"|}��J��^Jxψ��y�*�Q�-��b�SO�!kF0�K+Ӧ�j�{����w��D*!<p�}��xW�o�T���A��Ӡ2�`��t���9�1*��N�9�yt=��Bpw�FVy<4�� ����ċ��zL�łeo��{��	�Y���+�9�3=tz�K|Ե��Η����EɈ�����P�؃�2$n x��"e�\�.�}�Ǹ�WՉ>�:�r��r�0wHqm��Uu�@p���MH}Z2�#�iu��.=1h���D�k+\g=g�iHPiv>�.�������oy��U�����{g'/$4ƶ�~�V�v0"�:�
�]�}ȫ����ا`��{� �~��lփ�za^��7��6�֋�:%�~X���h�K1\���94���<��/"��kR&�6#�F5�lԳ�P�^�����۶�K�(ŏw�݃���y��c�W~�3W`k���¯3J�Um*���EJ�tt�*�v��bPC�ŏ��\�� T�V�V�w�ϊ��ʳ b�9�A���36�Fvq���K]���/�c�ރ"/�Yv�W�P�T�jw��Ş�G�Xr���ֈ�]�m�K���\2��:+	�e����F���v�ݫW��zp�ϯ�
#}�=DÛ@��q�#/ҹ��e�Z!lp��YV�s�l-�b
z�)�.{̍��s�1��CXf3pE8�;�y/О�~���GM�6���u���d$1��N�J���o���5���R��˩rZ����sT��-^����bآzu�u��d��r&3e�����x���wQ΅L�4x�ccC�B��_��g�/�j\��4���� ���(y6E��pr�Da��������a:��TF�d�P�+
�#�ĺ�x�����*��Ic�S�U�g���n�� �on\�*/v�\ᇹ�O�
B��N���eY��]��X1��+s5R���iQm��fz���^�E����'��t`�`V�\�bub��b�^��kx�˹���}�4��(����B�A�P��b�xL�X�,չc��a�֯:�����ɔoX��}o�.ks�IyG��/����L�𭹕x�"T�S_[�o��m7+�f��Q����8�G2��*���gYgob�@��]��J`�wV��i@�S� n�E�"���}��E��ˎ�h�u6B��.:�tU(eo_��Z�	w]2���y�ʵ��*m�_;GniI��ɕw����"��^4G��X�C���TW�.�
T:�Vj�{p+'��6�Ur��Ǳ���m(*f`t`�$+K�Q>���W��zQ�b�[�ep���A4��M{��!f��{�`�^n���P�{�n+GØ���e���ҩ��[���HTx.v�B+av��;�ꏄg�}�Q��Ԉ�(�c�;ڬ�.�ӌ�,������W=���	3E˨xh�.����޹׸WZ�f������/3�Rr�Fw��e�g��\ƺ����D�8��K�F���Vs��	��˛>�{O[����	tHG(Cc�(�g5X���6���ao�������E�)����������^�S}����.�z�6���N�1��И�]��Y4=6�y�L�w�Y}a�{ӽT򣜡0[(p�K<���\=iV�f���������W��:(J>�];�"�32�m_�8O
at�W˵+��m�ͫA��O�͏�Z��8�� �=wwo?����Yx�����C���<�e93{��bA]jWӮ���*Rt�s{kt�nd��E L��Z�%���7n��)"�Fy�8ؿR콌	���"=�Т d'�j����p���ʕ�SO�kHW�E���+�������s7��04���U����b휙�x:�c�p�[�8�ok���*'���Ƚb�M��J�0�.����+惘�����T�H�^��t<��p������ʼ>���j!�A�M�T>z�/\X�>��x�J��*]���k�%�P:<�`�g������Ξ
��ȍ����3|\͸��o�Q M���,�_*^Z�t���a��`<W�`�0�Z}�o<e��m߾�D�Ր�sph�|:�R��i1.X�p��/�L�~o�+�V��M��}���"3�'H��4����N�Z;�h�^>hd�h�fizq��ݬ���{�t��Y�u�.+ER�;�\�~�l$�}�p�]o��:��4�����zT��|yTj�}qf	��*�|bU��c�M��;%<����V��u��W$f��>P�Av5��R�_Jy��6�o(�<*Ǳ[Oy�p��β���ƟKr9#�IjP8T�5��i�	�%���};�I��cXM�T�v�gp<JZ�>@���L\ά}au+��.MD��s�y:��8�p���}�qUt(�r���*؝����P�X[����Z�Wq9�x�l�x\�&Y��-Z�����k��-����Q:b2��rk.�},�nuL����-����t�^��1m���3��'HPEe(01�e(�"sk.�3�{��{�����\\�p7<����F�zx�����@��񯭈h��^o��w��3��CJX���H��9W*�y-�>"W]�b|EGb��26{�ȣZ��[X��R��4��R������C�[!����=U��q��(�.�td�q�Ge�X�G}�������X�p���)�ڥ����W΄+0<��,�yk;=��x��^�<8�D����C���*p2�q[D�tv�u%Y�k������r�h���k1��}*��ր�b¬t��4��tOi�8�xC���V.Y�c��+Hp��B^T�W�4:�!�
Ѫ��4?����<�]zǎ�7Gi;�;���WL��#r뀡J���W)�e��9Pd�Ȑ�)��z�3y�=Eڧ�g,���@A�%��Q5^Kp�4�l�/U�t��E%������g�W}	S��0�ن�E9�0i�Q�������=��b5�ϝ�P�[�C�)iY9K�+#��g�sE��2_ݞ�d�b��͜�!D1�E��ţ�U���+ʽo>��<]=��;�'f�G��&����]��z4�q(��ǃ,V�f�#���
����=���۳�����^��iy��?��}��ZܖtW��r����1��������l'u:�ބc�ݵ1��]�Q9WC|9���#��F�p>j�];W���s\�}�ʉ��N���jl8��
.)�`V:����S��+�:@��BN��s��&���\G��Ф=~���J���;gf]�:,�y�,�Aj��%���JXfr*0N@�몋�m�bT)�WA���s���do�ʵ��]/wjZ�=�ޓs�D븅@�LQ;�P��8�:�����׳�<�W�j�)�<B��"c*���I��]�<3�h��l0����#�=BU���X�
zxW?�p����c�}P��du����n�!��˴��(��o(z�fˣ��D�%�V��9�5m㈌]��������z�x8rZ;�7��u�	t47&��16t�ݮ�Y�q�0^��x�O�X�i�z7%t�8�o?�?"�k�x���\����U�)�N�o�HvJ���z�8'Qҡ̲xH�x[E�hG`�0��S�^��ؗ��4)��HX�]���O#�"�:sV��C�m���c��#�mm8��r���+�m��c �7��=2�a�b@ؚ��$_
�~��*�z�k�'faˤ�r�Cg�^9�������*��#��1P|�*���ʌ�*�sgSP�:�*���������)Gd�U(d-�����p���o��	pœ_�R�ڻz�,[j�Y�4�#�/�ax7����@0����(��ꠠ�:��/7]�B4���[�o��NX�~����ցiWO�?#�}7��{p��{���'u�˟ {#g�2&�7AƐ"�:�#=�֣��luO�[.W]E�k��vk��uB�N��{��%�z)
!F�ʖ4�Ƒ.,ˋ
�Lbf8���g����`Ik�}���Q��r��%D���B���"�C��~On!^���Q"�~�>wttl����m�Kᕆ�;�YnV���&�4ՙ��ŮT�z�H)�Y���*٢��64��"a�b8�P5�GI�f�[�ڑ��<�����e�+�� G�N��s�ԫ;�P�Z{��m�Q�6�T�S|c�|�.-�����z�j��¶\5����)Vr���ܳ���ÅXU~�) .yWU�/1
+��F�%�����,Uѵ�Ҋ�ۨ�14��^UV�H�Bw�y�6�=����5�H�P ��{T����g���� ����4��^7��
�ҫ���$��Z��2�|�z����Ƚ��v����ݖ̭�ʎr�Q0[��
K<����p���0�{�Yx��z��[R�:E��h�Q~��]�0w�͍�V���/�� m;q>%��S�!o�1jX��������+Q{65��re�D���R��;�%��O�k�����.��ʫA�����d��-�������<��X��yn/�Mds�]�=ۼ�k�	�q!���.T�zU{�U��=AG���ʃ�r��:��'d�)�Ԧ��]���MpF­o��Ғ�Z0J"_�QB_�$���K�_I���Ά�	f��v=���v����n+�+ϥ�T��������� ?cz�e}��O\OGݔ�2�VV��ܹ�p��8�7�
r&�ު��6͞��6Lӷ�C��d�-ܼI��ݹ�zA�:��Pu��_w[�J.�^m�9D=�Z��ӷA�e��]�$�A�4X����[�ݍ\��jѹ%�R8���.^��Xe伨E��F���n��j�W�N�gV�y��<���ܶ`�,&>ޙh��˜O��s�:�p��w+�̾)>8mX�e1{�����;2�4�,'W����s49!Iㆯ�+!�pP����g����ɏb�U'�eI܈ǔ9P��N�M�K#Ӥ^�O�]�E�m������ڵ/��1�G�E���)�f�t��v����əg/k��m�[KP)}X����9�9ڂZl� Y)K��+��lޑ�_VS��5�{���jZbȆ��l��O�2�⌝�dmr�D<-K�����	;9�#m���R����S�o#����]8M8��h�鉖��|n� ��e�p�]u`�br�6-���2� #SZ��h7wQ���=����5
O�-��lV�g��h(oLw�M�o����}!"��I]֣��A
�ۆ�w
F��ϸ�֡W���X�
�9��]٩F��4�fi��e�>���խ
���ɨ��"�(h⣊�m�V��Y��r���ORLR�0
��ET2�ٺ�"m��xV*g%]̛h�GMw�;FwRٲ�q��͜�դm�N�m;ov֡�S0��KK�n�G��K뺚Ax�/��u������I��S��J'���B��f�h��n�6ʁ��O��+;M��[B*����t�{f��vN��dP����G/�_Y�(�á�pѳF�m}�*[�������i�Ju��(ij�;�Ct����gE��N�ɺ��i=1�`n��>�Q]��s+VJ�r-ӥ�-�ki�r���dY��LrT�.�B٧݉}��O^�P%�]����V�L*QN���������gGPg�X��7^���V�L�GYw�뚭��һih�˖N]ڼ��5c�z[i�d���a�t��+X��㻿��C���5�1����pk
��bE6�<qIS\T���=c�mq�����._̗�׻Y1d��{m<�F��t�	˺��U�d�Pu/��y�"R�a��r���$�x�W&%�< \u�Nޫ�b�3>�f+�I��baFuGK2��	>�{�n��`��ٶ�6z�o]�Q��Wv��&;M�WnDֽ}�tȝ�ʒ�u:��e��k�y��c锃��ˬ��n�X��+v��4)0��)0�ǽl���Q����UH'�`Ƈq�5����=���|DR`)Ե��7x٧�h,)X0=iɆf��s5}�so�)t�EZ�B�*�TX
#�a�b�1�q��R�HV,�10b���*� �Y�l*�����[��\31�EUb���eEZ� \�YR���!����K[R嘖ؠ��j*�h�Z�1���81jW�h�\E3,�1��1���V6�"4���-�R�!naV*��Ҩ̡�嘙pɉ�f��ȉ\LJ���\�pJ�8�[q�)2ܵs�Z*���LF�̈�*�ڶ�rظ�kmRڥ��Kq��1L���r�01�.�m*�\�iTIU�J)���iX�)kmL0��`�*�2��l�b�Df5&YCƫ��
���R(1��G�,dr�+���-�D��B�iLa�K�#mq�%kU�
����6�\h���Ƞ�nZ���-�Z�5�DF-�\q���QXT��0��D��c���6�����Q�,�ֈ�F�-�Ua�b"�����\mV�#L��km��VI+�^�&ve��Ic��a�j��]&i�#B:Ԙ�X�#yY�M׻e	0����x�SJE�i��ö[<���\��������Ր�3є:�R�g5�ϒ����+���T!�^�OTɽ��ه���� x1yN���PI��VjeÏto�\t+�)�n�)|/sV�1H��u����VG�]nˊ�T��T�b�g��2���FE!��$z�f$�"M(��pd0mV�K�Y먳��D?Bk���F��x���%/S'�<u�dד����>�ځ;f._FlpT��ڸo�����nK�;N��[b��<��~��>�G�ϔ,�w�ڱg���b�=l�ʖ.2�����z��.K*��K�J��,�Ɣ.�nWL�,�����W�Q�4�k*si���ΐ���T#�]>�����z�S�'��WcQS$,E��Vv6�(�^Z�q�q�j��o.�UA.Z���9�26!����P9����K&�R9K���B�n3��~LXo��˾x���ٍ�bn�
4��]J<E�BSxk�ܭ���{W���V!Ƴ�3�9�1���L�|
�\������'�:�*�/U���(T��e��M���+���1�6���a�n�6�sܺ,ɛpp�C`A�f�c���^�<Gn�hkw���E�]|��i����йo6C�ƚ�2Mǽ(ߨ3�F�y:���Յ"��9��^D���S�V&al�	pL��Y�D�A�a%��U����,�/���i��ϱS��*8)��Ν��w����
n�s��S�5���� ԍ��2$n�I�O��9e=�s�Z^�c����5�w9�]g4��
�[xzc"!E<�PVq����Sq)�!$Լo��̔v��x�.R��W�VE��;>�T�m8:�Y�4[��IG��1�X����O]����P��c�=��Ϲr✼�f��B����9gMevk�'+���!:O��`�Z�e�,G���x�e�@]K�iu�t%�{�Y����n�wGm#�52����`T��'#��g�X������^iy�s39z9<lGb�1����La	��<
kU����z���3n�5�넧j�{�r_�:_��^��+#��сA(E�lp��E_�D�}mY�Q0�îuO_B���%�[�]���]<��wAn��I�������f���y/�l��������W��I��=b�k���S�R�]}@̬�)eL�͐Ã�_W[9O�S�ԥ��t��/�mI݉S��Cj�K�]�c��<goQ-�P5{ʟ����+�W�K�����:�`��Pa���r�q�{�/��]��p�yp8P���zۮ�u��%WE^þ9�G��77�y�.�6�NV�RŬ5�1��%���j��йUE��ѝ)�l�hd:�2O�'�/�;�ڲ�+��׎F/��������O�<+��Gٚ��)�����EZ��?%7��o�D]�$�U��q�O��q�(@5*�甫�Q��`����ɻZ�_R�áУeW@шS��ێ�T���%UB�� .�tS�Ua ��/3���İ2B���I��NG)Z�t�>3&��`�q0�J�����{n,�ξJv��w���,l�[��4��ڋ���R�$;���s!��弼��}7=施h��88:8��h���J��ɕ�O��S�����JXck�H���wS�<R�ۡ���"�t�apoʈ�M`�Lp�>+���^���0R��Sn̰f_)W�a���7�e�L��2�ZX��2��aܺ�Yp���7R�l;>^�-G���A��n�%�4�\��* w_���y*�|ĹR��Jp�JN�|�U�T��ۓ�Xf��B�3�%J���V��3́�� k&�|LF�J�<~G�,�0W��-vg�l���:�*T6�7!FhD���W&c[��>�luMl�\*�`������y��M&x%�~�Qو��J�d`�h�]rTE,�"6B�e�鞮���N�=w��;�+G�t��1A���|�[���9|D��O.�.HȰo���r�w��}�.uC��h�[������S>�@+kx��g���*�`�白^�b�S�^);ӞE+=K˱��P��3k�Q\;q`bi���*�X���V1��M����<�3�����~W�T��gJAe-��4?���@��0v�Ά]�Ϛ���k�|\=Vv7�����;�@�T'UX7f�@�t�uTƶ"�+�z3\�]$(�d���2����mS�ʌ�K���M�����V>V�_(�ʷ^�Q���7p����r�U�a>q�h,T�q	��	��+%���_�|����� Z+^{6�$��*5v̫P7���,��]�Ta�JtVh��"4}H�OT^��h��+�ElOUȺ�x�d�u��2*�=��Z�䬮�vj���n�T�-�6�i4�륽F�J��pH��lD�3$����&+�ǕX%�����VB�/�H[�~�!�bnU����"󱤭�{[R�����5�]���^%�_h��G�����8v*|�<�E�)�/0^Wn�i�Z^��c:�)�1a:u(E���2$u���ҩ/
�����Nw~�9�|^$�p���1[���Dؗ�&"/����Gt�輵�1�k��S�z�c]՞RV�v��U�4�ԅ
�FP]o��sph���l䴒xf����g���6�ފ�?{C6���.��T��Hv�].��qiu����Y%=��o�K6?J���ð��Jz�O�]l8�2���\��{#\�!�[S���1g�w��=Q^�����9^��bC֠υveK���[�"x�s�O�����$ �Ş�}cA�L�'�� �Y��\2�`/�kr#t�3S��������S�j�3�]�A���ۅW
����Kh�ݷ�E�x�8��O��oY��l���ZiR8E�5�QE��W]�g����9u1u���V�i��Khc@Qgp����<5f�	[�.Q��`i
ؑ[��'I��h.��N�����F��I��8�5˳��/3j/=U{	K����_����W�Q�4�M��ɟ^��8xD��E�J�k�+WC�@��Ϣ�\�@$3}t��j��ҋ��YUҐ�Ҫ�;�n;<���
�}~;�Z���y�N3>?d#����u�ZM�؞{�U�76�6]WU��z���C8/Z��j��ã��:<:�r�Ojƺ��E�9�ڷ��7<'\�8��(��7@�t���P�lU�n��=Oe8�=Y\����g.u7���1��u&觽X9״�n�;�*U*.e)3��BU9�g�����LP�I�X�VFV'����?*�6�)G)�5���A�5�:�]
��zM6�S�m��HX�'��#.e���*=@�V����Ы"!E<�P|��G��`�j�(WJ�..<|�M�b��C*z�=X��^ߤ����������Dr4;BV
6P�s.���y��ZK�|V���P�]R�]li�P�O���C r+�vL�'�gnZ���~�o%f)�7Ej�OӍ;76������' �ʗ�VaјM��t]5�a��R�)�\xa�����&�>��s��a�@r./��-V�j��Ѓҏ]s�Ε�65���Yq�)�Y]V;89׻��3�S�N�ؠ9�nA�Ǐegޮ��%����5�Q,ht,xV�����z4D�C����#F�s��I��ީ��=��d�9+�D���rl�}��r:hӇExW�T�a#�~YC3�t��f�"=�;A��>�D[�\���b4�ԏE� �Z��g�Nn��o�t���b2=.�z�(E�!C��`bup&~;�r�`����s�$
߃�{�_���9�i���\�ra��ЦO��r�?>
ŗ��>���`-�I@d�߂�a�š�LU��Q!�{α�
f���y�imk��.�ȴyv��U�G��*�P\�ނ��a�9#c��E��R���be�iL�^r�~�ݒ�p�?zpY�|b�V����(E�%C>�z������]Rw�mZz�:����EÊ���s 犈���tg�쫡r�M�˸����Ÿg��O<$iT2:��^!N3[.5��u!W�E!`UX�?+����,Y�>�a��5m�V��޴�J��r���UX��@l�(��p^p�F�.V�nc�E��u�q���!��M��p�]q a����h�f�:�󹕯n.LժV#�y��~=�fʹn5�u��ҋ�(lkn<��ю��1�-Q����)��o$t,�!t�zA�*�c�m��)��2":���h���j�:Z=Cx��>]�Y᾵���n��^ȴ����}+K���٨Bt�wp�X��G~��l-V
�^tx`�������J�:	LUT`j�Mֻܵ���L�Y��qP�@a$m��:/��1��q��Ҍ�Ů�1{M*��3�#����Ԩ(x��~�r�|��$V��m�Jx��?��M���l���k�^k �SưE�3�4��U��Ȑ������2�� v\V>Ft�xd7��ϖ�[O�q5��o�!DhY������G��*"�z�2�����q�<����{��ʑ�'�>,h$�
=[B�V9Z�C��y<>�y�][��n�������Dpd��"��կE�%CPR��h�q��Mo��k�r�#��A���k"{�(*�㢬���W�T�z�����T+�Ǥ4��j�WԮ����	~ܹV��L`v����{��*�Ȕ))դv�yP� vzh�����k5�q�{��`)����W�+�fs�jė��˫���^F�N��vǊ��:84M��L��tVF�����ʙ���R�n�:��{>#f�浜5H]�z�4J���_V��b~��ɣ�r�2���}.���~S�Zs�mZ�Y��P+gF_�;�e�|�R^�;uc$8��$s��c�pR��#�m���V~�{���R��I�xqM������QQкH��9W�'��-T�qϯy�
U����X6�y��k���b��U��ž$V�qc�.{~=!oU⨇�:�P[S|q室��%��{�hL�s~�Q�����|�}J`����"S��G�աUs�{l!��������1A��:�"�GB6bդ�>ã���D����go�H�맙0�u��vR�¢lK�u, �l�Xa;����K�Q��\�����\����FX���&�8�h8pD-�s)u�y��P�5Kg5���`��^:*-C���)<�QZ*-�����а�HK�.���<+���Ju��'xVҙ�2��~��/�]��9��56_��xWr41���>����k�~��l�ʻg���t������P+/qłNԗ �*�M#D��T7���o`b�HC �\6ʾ���k���-�3�P����'n��]��Q��#Ńc^8����<<e%Y��CR>��7�+#�E�8��W#X��S.��x`�6�C^R�3��o��J�/!�޵:\^��Vl!���8]{�O�@Y��혏�A��ׇ�j���Nd����w��(U���� +�����21�z�]�j�O��6Y^�1nz%���*��n�,��P�.���s�2S���lm�9�Q�*�Cxg6�g׬�JU��y���������r�E�WL�S����lXO�ו�L�E7'��\h�.��zPNe�u���5��A
���)�r'��\���X���1�x��<�ם�8���|��e�j\��h���G��U�9���M��G�X�7���^1K����;�����XP��g���~�i����	����o���6�<�����)U!)JH��Nd3���UMs۸t#u�:��H�\�n���rl���	���n�vՄj�\��X�ؼ@h�{Cq,���f��k��A]����N�ÿq'r'�08N�R�u��\%,�W�NU���hX&��X�!X�D@T���Rd������.�jA{Gj�ie=�Z��:}*݀-��5�����Q��m�i�Mu

`r耾鹄V�iC���n�33a�J��0���F��H;��m��.m�)���ݽ��v���)��U���k֑�����v��y�mbAU��m�m�8�d�F����S��*�����.�b��� ���6�J�e����z�j��nF*ն����e#M��.�3SU�$ⳓ�ݷ�L��s>g�Kng2Et��6�Z4�R��aO��]��K���f'���'���k�s�jPPZ�$� 9x��qAS��t��{��/
�� H�o��^5��q6&V7���4�P����T�����b��:�wH[h,�B��A��F��zˮ��W_�(��|�jw_e��j�g���C}�#˽*XbT�O)����9t�jsxS[N(�:��ۧ��:�Z�N�'ˤc��]�1Sݾ��qvR�`�ٷP6�k��k�y���{	9764�Q]��zֶV�\�t�>Uz�	4GT��Lh��̉[E����8��� oe��<ށ�:��S���VB$4�S���[�D{y9�]�
�Weqy4Q:��ku�s����[pV�1��k�e�S�E��Gp;��_׷�S0q����a��@���3�`�8�)���� r��n,Kvev�wWp&�QV�;3Ф��ja�틫���C��M�ťd��	��-�)�Xr�M&��|*�0#⯤w����n�Lh-���+rtJ������w(l�xm��	�q���C+��%[��w�'�T���v�r�x��&I��S	R{���r��[��3&�0t ,���G���ۋe�'tl�F��K�f���_5���GxÎ�oK��a
��h1��ӏ�U�'ϵ�m��(�Ko�!�<9���Ѻr���NJ�D�������j�cuj�\x�؝�����ރ:�>*�<�����4���_9�Jؘ���R����F@��ٴj���J��
N���1<�tT�т��f�5b�d[���M��_-:�
�Y��}�%�I�6�����ǹt�"�9Y@�.*��p1�i�wt&��>Nf�-˦�ԭ�bn+15:WWC�(�I|c!d��*keI�������ץ�bf�����t�q�V0�+��A|0f�R��.	E1m2������Z�,YZ��F"�+KkR�"���U�A�i(*�6�h6�(��*�eb�.9�Eb�DU
���ګq�FF*���5��*"��X����iEe�R�fZ�e\�qj�Z-��QS-AU\�Er˅l�(U+C-ķ)��$EU-�1�q�mJ���P�ڊ����c(����ʂ"�m2ʎR�-�TYR崶T*�5�+N�b5��i���Ukm��`Ԫܸc[em��++L�D2�f[�̸&*\�q��[lP�TE�11*ۃr���Ȍʹ��嬹�-(řh��
�%�֮[q�1��)�!V*,�DI\pG---ʪT��.5djb�Kh��2ҹj���e2�W3r�
���˘䪅�c���b���Z�F\Ƌ�aQ���(�+*��0Sz��o���{�[��y�v���7�7b���)���dO���b�C�ȝL��fMn�JL�ُ;�.��>]t�v+[��L�#�q�FѸ��.8K�ť.����^Y$�#��p�J��^WFd8�7��S����}��e��յ�Cޤ�y�p[��Lv��g�޵>'��u��Gm��9Y��a���U���������8����pK������V��Y^t�R2)�&	ܘgJ�+.v�fhO�z�Ə��G h��ׁ��M]n�y�6�����i���wG���nd��rWp�^�BG��Q���4���8�o&���g+����SOC����)T�˸x�Ԏbe�?du��H�@UͿR�7<�wB�u�jB�A�@���(s���
:�D:�[Vfz�D���l����	z,(�(Mⰰ]a�r-HBGB��5X��y�dP�[����U�v�ܤn�yY��7�h��.�V��+4]T\+��J�3J�8{0�fT֕9]3�����>��+K]S�D�V��vJX�&�M�]��'P��A�Ck��&��<��/2�);��CE�S��X88��.�����n\�[}���^��f��}���:"3�
(����e�Z`�[畿��u�m
�P\�ނ����
Y��2c:Ԍ�����=G�B���b3�<�Y^���͗��j+T��_�U(5:������oT���T��^6�l���+������q�Wn`�Q�㈻��3����Z�;F⶗���KW ��<��HDu������B�f�n�u�J����)֝�:S�G;۹�m #��� ���L�
��Bޑ�F���c��Bnˎ�׉�>���r�s\h�|<������$*:�L��}j�����aX(��m�B����i�2�4y�ǬJ�PC�n.GjZ�����Z�҇f)GF��P�[��nj<��<�|��*D�W���w��<�r�Ô-��t���5�V<)���1j�����w5k[�ڄ�Ր�t�#�`�&!_��i����ցiWJx��{�L�	u�ߊ�wC������m�!���K��a)
/B$ʮLƷU��.�����י����d�X�d�ډ��{S�_��\������M�	W�*퇎�x�;�%�ei���B,=F!!ıN)�cyVG�;@�S�0^�ekU�L&�K��Nm�oʕu���r�5�`S��	j�>�R�&�L��{�S=���X��tj�[���R��2��q~UB`M�4Ѹ�	P2cg.��:d(<qh>v�BO,�������	T0V�/�Q��ۅ%*Y�VLp��=ţԮ�� ��Lt2���V�E�3�j
� Z=�z��m�L��W�ЮU��yE���qv!�S�墙�����u�!ic�̡��]�F��}.�-�J�^U��vaJq��f����1��v3�����h�:uL�y~�}��spM|��#)mL�.}���f�f}�4l�;'�o�5Qޫ��˭;�9�,]pX���1謤!����	��Q�}���K��ˌ���{	�TmW&��YȚWu���⧰+�X�ܷwt��냂,Ͻk���S|�\����%@grx5�&���T���3�4FX�G��kG���%�~]��1Q<E�E}�᯲
'�!�n$�؃�ud�[��Ba��c�ux�GW�)�5p�ڮ)�v��8�9�����`�v��vz���:�>�GTɵA�*r̛)�Ѳt޻�;��R�T�a.J�Q�z%u{��Du)���]��듣\z7���{+t�k:���2��Wv����#r��c�Q�b������t�U�n#�L��ܺ�LôH^N�JbdtT�P�x��C�Q��<�ε�ɽ���w��܍��@��.)m8�����R�&"1���l*
��B�����Aԕ�B@H����g����V�a���=����j��kI8�0����a�Ho�7���ȅ��Y���Wg���HK�.���<+��ҝB
�J����J�wȕ��.8� �0o�wrݐ{e�
�P}���YIR�G�UڱW|�E������2����٫�6�.��P?�
���|]�fǄ�A��lx����*hi搎���3	��uN��yw��`����b?5�B^U��Y�ݡ�j�ڽ׬�&�� .�Ng�ё���(���ժ�& 8l�*�Nˮ����cN�aOlA��0&�ʘ���9����Fh�s����MAo��ٿ3[��%e�;y{��R�6�R�ٕZ�w5�!S23U)�)��u���<#c@���5�N���#��x�*]���ˎ��^{x�o�2��1��ZK�H���ܸ�Y�,њЊ�(Ƽ���u�de@�.�H�fgL�̭�Cjnh��ؑ�ƴGk��G��
\4fHk�[��m�<��%C�W)�{�ŗ�ʹ�PbU��6� u�Ǽ>p9���^�D�px�(�|y�zly�{�U櫓~�t���#a��j\�q�.v9͌5��Ҡ%*�AVq��a�Ӵ�uy��u.���;�a�U�[����f��#��g*c���^)w�Ba֩V&aGA�<���{H�
�HP����̊�JA�i�ZĴַ�/���;|L)�.��y�S���#��Ѹ����vO*�q�/��yv��*�?W�fA��똅��(���g�-�=
�2"��������
�-i�T�UG���ʘ�>}��5��>'�(����Gm�� 7s��R��w{q��fCϐ]��
�x�ڋ:��ר��W�z\[�j�6�+�+�z�b#�6���`5���u�4?��
�ׁ���`�J��㛟{�^X����9i�5b�.�����U����#�o�/��v�5!â�_�
���;7�q`�H��yR�NIY�n�h�H5�����h]��͖#���I�p
�u�܀8���(C]E�L���K��v��<�T&�!ܑ��.O$;9uĶ]�o9�%�Lͻ�<�A\<��Jׅ�8=м>}ȋ}�z��F���WV*}��,�ΦK^4�a���M���B�D�t
YB,9
��� �\	�9ᬑ�3��'�͵5H����\e�y��2nE� B$d�)��ܹ�}�oB�b�*㫜w��igR�Dؐ�舗�,3����J�b�&�d(鑐Nzܷ�ԧr�&��o{�郦�w�X��HW1Ar�zMGd8d�����瞋�ֻqw%7c_V�E����e{SWc7��z|z^(8v|��-xJ�t�K�įh��h��TkK�T�9NKj�6$Ì�h����3���z.�y��u���N�mn��Q������7+�_���P��9\\�)�n7n:dT(�=Ơ.�v2'����M����DdOu���^�M� �ʆ�߆!N��1����dSk�s�����[q"8F�8�2+Р�Py��~�|�J������y��K�z�tn����ⵝ��m:�
�NЍpzV�K��t˭��J�>+8v��J�+�>��JKͧG�{Gh uv
;ޝ��u�5\�Z\�I{v�Ը^A\��1Ńٓ�ρi��ݙR�ea���՝�9yѽ�C��R��}���O���Z��F�zȊQѷ���� L�Ҷ�hW^u��ʏ��v�ʹ�츨:�TF��"�N��Y<�gp���Y}���s9m���d���r�ιW�Z)����[�ѧ7��b5�|m��U磪LYp���}7b5�hqU<�W���g��aZ��
$Uɘ#[5ң���ҩrI	�{����,3=2�� P�1ѻ2��Di��q����
�6���z��E�Ez�R#���`g�].}>f��W�xUY�>�(`�{�ox��]sg��<
��=��Z"�ԢF�'�D���6|9�j
� x�T�c����[;����,v֩s!@������dXg�T�<tUѵ����v�*V�	��v�}3�G���\_����u���{>8�4а֙� �����׸���ήM9b�r�\�ʚ��Rϝ�>{��P��Oi��C}}Bw���j��v���g�<{m-�]�][��׳����;��+_��J���1)�3G��'ו��GO��}p�&r�ؤ�
�C��{��tC�L����?J2]���hoǐ���}��E�\�,�.[��֗d�߄�����'Res�u	{�e�Z�,t��$r�����;��;ޣAg������KT�7֫C`�aa�;�üzcx=�u�9�����&}��/R=������Րp��c�|١AB�j�=�YAc�B���oy������t�;�o)'��3xe{��E�]dyn2U	�bB�"pP�OW�tu}�����<\b�e���g�O����Y[+�s�]V��)��:�.o)o������y;�e/G�֡�P�Ӎ���DH͕�.,7�DÏv��wx�ۈp��OƷؼ/�Y�c��b�|�N��+�l�ώ5жC�!!8w�����
�����@���zn�.}i����b��W�L����D�
���:�T���8RM;v��צ<�)WM��K�ށ�w���)����N��g��)*�d�ͺ�r+}��i(�{q���l�N6�>�1\,a�Z���|�2���,�u��-k�A݋��-�#�^jb#Uį�Y�tm�(��gP#����H?� �#�
ve����!i�6>�#4]of��t�P�E�����������.A�%�7�XJ�е�MN6�v�Q�ֻ9� ���W]�v�=�v������x�r�~h����p��m�$!������,fЊ��ʕ X}�9��c1�ή��� �?L�g��rw�?_�m�8��h��n0o��TQ��2�R�p'��-����t�_Ԣܴs���8q�/J' Nx��4��+	���׸��22�2�\�eZ��֜K����-�&����yl�/���,Z?5�x��{���Z�ʯ�|%��sld�h�c�j���ޯG���{]!�����jj\Աx|���7S��xh���f�g�1����`%^z�<�8�K����r�QF�aBJ�3(�٭�w�ڌ�NOWw�����R�Q���.�u�>��w
�H*R�:+���K�Q������	u)�s�,�X1ţ��4��V�07�1���X��RϘ��l�xx����s\��N�ss+���n�+]�=
��	�^�9T%C�ekv�f�엮o3n�n¹ELI��*��a�ܶR{��ޱvڠ�䓷e�׶��Y`S��2%,I��>�֕F��X�
9�� 0�{V�E�S���Z���3p��]���W�Z8�W����Ks��ɓ�Է����`bF����ʘ� �!X5�*�}׷$(dv�P���C���hV�K)���^�~β:�u�"(����Z>T �	yy����V�?K*�7��n�k�]�g��fr/ԩd���䉺8�$��4:�cµ�^͌�q^}�3�����0�h�J�^�ɺ��mN���)ig#�o=[~:���kf�-�J=CEp�l%uo�4Mи|��ލ�g������?kx����m9{�}��6��d�������1h�>��\<w�l"�Ŋ0�ڋ��6�y��:�K�L3�\e~���>7C�Q���u�W�㥁�HA�E�}~��q�p���C�����E��^��X�Y�t����w��o �G;�x=n�#`�N��tߡ�P#� r�PA��Q=�0xP�]볙%��S����Z�ҞV��)���%���ڊ�77^�:�E��?}-ʑ��Wv�7Sκc�X��mG��Z.L��X+k��"���7z�`�z�����V2ދ�ۢl'N��{�L�Ci�^��6;S*
8��FQ&�VY<��oP��:E���K�����a]�-ӣ"p�j��B�O�Ֆ�h�T���oT8�����������>|C��rcmnf+�J"���6��'3��A�
�ov�9�V�c��r;�۔�Kx�m�s�#�u���-)ϯ]QgVFN��#��˽��V종�/l��>9cA��s��\
r�9��<D�%JI��]Z�4���� -��c�oʲcW��w5��j���ũM��+d;2�[�mi0z[��kE!u�*��L	�bU�oq���{����k�t�'}�{R|�=Y��m<�T�3e�r��)a��v�A�l�;J�K�M����;b�3���`7�������AXҨ���^ջ�/9���;u<\i�Bދ�R�&������ʘtcTq������*c��>��+&I�m!`�6�o��&ɢ�۬��Dmn�R�#F��������f�>P��0m�S�$�D⫱'FtF�+;R�f��F��9>�%Q����u�:#Һ�"�a�p!D��*��dX�kvT꛻�3g��Y�,��4�Q^��g��ʳ��-�[ڥ�r�0�¹h�̝��d�Jͬ�S�(�9���w��d��#��f�w��HBu��!�)60��0s��9]|KL�}R��Wud�J�� !��o����T4~Q����x���al=��0K{ٛL�Xc��0D�_muԂ��hV��Nu�˽�Z2��-�Μ�0��衊��7���η+Txr�q���WKU��ԍ�\YH�V���{�Y�Roq��I��7�&V`�ǯ����cS�-�#����oY�ԛ�3�	M���'��ts�-U�)�˦~��1�C:x���߱d�MSTl�wܲqw�*�'*U٢��Wd���*�����<�D*��F�ɣ{��7m.|��(uem��/�*l��c��	8�n&�\�Y'T#�v�,��pwKځK{7u�w��K��zqLet��!����=F��XE�A�g0ܧ9���X�q�'�@�ҝ~�]u$�u�5B�cm',jt]�q������#v��� ��bFU�ů1�$M�}A:�iYv�w/�K��uѳ����Ӵ-���u
}�ɹ�� �#,��Ը4p��֎�,<�*IB�޼��EMy�����0�r�І�nG@�jCf�H��KԚ�M{([�Ĳ�B<�.}���[
N�e� ]B����m�7�Y�m��	r�-�%��*��Q�YZ��b�1r�1´J�FV�l--i�*$��F1rܷ����e��b���.Z�D+��[B���h�a\�ۅ�r�J&P��X�q���Tm�*
��؉��n�.�Dc\��UQSV�h)Z��4��c�Q�Y��ә�UP���b�*�.4b(��E,�*.-�m4��&:sUJj�H��j�mEDR���m
F�UQT�s1Z�EE����-�F`�3��)UT(�V(ۉUUq�!��X�U�jbK�b��ҮX���mTX����V�R
�((�.�q�EP�[meb+]8�.�eci�X�J(�E��AdƘ��1�kY�P���QDEj�[f0�V�DD�*�H(��)�k[���`��]4�"]eQkE�N�TQ"�aSYnPFEV9lUU�P�Q�a�l3E�AT�(�+Z�^x�;�����s��b��(u�����5oXR��ˤκ�Rw5^�J�2���^r��b�0ou�ք���g1�+wI���T��B�b�s 犈�q�/&m雵��N��_r�{g��e�*:f㜮�C>��Χ�͕ꁅ
�������L�;{�Z�P�C�J��
*� �\�L�Hp����}oH<�oM��h��
y`t�/2��d�L��lY4�te
��x���i��}a�SͰ��*2'�g�󼪉+5e��j�2b��>�kР�w�#�(Ш�Z5�����ڼ��&�/!
R�)��'8�B~��J�:OLߓ��١
�Ld�R;��
�����D{ڝ�֛�}��{���/��r�5�����+�T�|������ȍ뻀�-��甪)h,�� �".h�P�E�b�y���\'%UùB��**����]\��ލ��L����5��m���UָU�#B�1=S��_�u��
l����Mys��,�Q���W�G��.})��)VxU�54"�{�D�&���"9�O9�U�Kp�U�����c��"�)��F�t��q�9��b?m���N��2�yq*jM�����K~Y�=����=$�����7DbxK5>���;�]*�u6�[a��Cٴ�b��͙�xea��}�b���u�溁����p����o���'��gò���UAYw5ZQl������Z�g��<|Mp�2�2R���SÇ�E:6�5÷kiL-�a����WS��UV�w;.���G_U����B�֙�����%UJ�]Ju�r�[�T(!Nl�ć�L�^׺{����_G_�9�C\h�{�L-Y\�13���7�G�sK�(}��W�(�8�\��q��8�������G=�y���=V���Z>�X���: T0{��ۍ��-��o�Mf�k�v>�"�k��/'�8eQ�|�q�0��וR��|L#��"�G	��H�6L���lGg=����<��]d��q�U	� .���*Tux�GW�>*�6�`���:��b�GP5��"�P��ܺ�Ϫb�+�<=�U�ҹ@�R��Q]{�d�gщ!!�<�����%�hQB^�ž��z��ګ�� *�氀_���
�Í�5Tt0c���kΥA�#�����T�g�U�W8�b�o����+%R'B"�V�P��S����f9Y���P��grz����,el�M���-fX���}���T��[����S��u�\��Z-���1�
Ґ�P\C�&
Zq���>ӣ�~Y^�]D&��C�nf۰b�,C�)f�3�W�V1T�%���5�U��K|_�a�ug��ω(`t��P0��+�����I��V�Y
�>��Jt���_�|>������|;V+}��~#�=�奏�)�S���C�|7*\���
I��]T��;ІmV�K�Y��צN�g��~��֩[k��&%��J�
 �i�Nl.��#�r}8�0�� NٕH�����=�Q��8�r�(\t0z�����d���� C�)��3u�>L�e:^�"�7�X����⛽>����%�мr�b)s8�8��cu���N?eA����8����ܿ2t�����[R�U-O\O�<�`j*d�����XϷ
nߤs|�,��;J�5�D�Ƈ@`�h�>6� u�cޔ��*����n:6	<qW3�.)/4��6G9xn�k�^���{]!�����j}�pt�x|���$a�+�/�Դ&��2,v����-�݅)U��w9��6̰/�:$�Aα�z�����g::(���+]tou�����xX����JΖ�8����ih�a)��A�a�K_����N6dכ��wc����<�7^z���H��䮑��n��=C�)U
D�u��r�5�����=�>\*\c�9@\�{]*�m`n��٠�*�B�����Zhĵs=>]�����	��"]v�]���8
&yNb:4�1�7�%�Q���:�F޷s\jEDQ�2��g�A*:��WK�����y���oB�\�We����)=��D/I�=��x�5Dh]��)���D��!u�ηٸəe�]�+yf���u�}���n$��.��Uh��y�`ǋ��S�}��X�梻]�nv|��!��W"�.�+����H��h�t�H�D���,z�����#�6�W�>bs�lA�KHp�W�Q�n���J��h��6�}<���ݖF�M�5)	�[;@��Vuo���x}�H�޹�DٌT�O��N��l�DT����q�:%�����!G��@�YEp9��0L�c�nwa(��}��v%�J_*e��!36�2�v7)d^YȘ��P;}9������K�y��5�t�̸�F�Vf��//���S�Bb�՜���%�;���:��ҝA5B�z�wrt�'ǝ� ���>���gQ�m���z�ɯ6]�w�-��.wuJ��Jۨ��N,u
���/�uEm�S���Az��zo��
Źٗ[�E��`a�t�1N�ج��8?.�P#�fqE�s��í����{�ؔ=5S�*�^��+�1As�އH��=�܎#fk��Z�w7L���C�){MH"/�<�+�|���\oO�����������W��7B7�=Wy=�= �l�9NM����L8���MS񙴁;�9$x��=z���Q�]w |�W���l��֙Y�=�ێ��8dm֭�[��t����y���@�Ȉ��X�G�ld�,a���-�&*jzn�qֆi�T�6J���c ��[���ѤD��^�s7�y���o���nY�jv�i,��#��L;�-��]8�(S�1PS�S��Ѝ���X+]��]]�X�~���f�i�[���޿J�N�z����Cܺ�D���Ot�ȡ:0��5�ն�P�b��<V��dVm�I{��r�!3t�zw�[�jl{�z=����R�et�쐊4n����b}���r��٫�t���Jr�$�a�y�8��^fμWsju"ˉmc��%�>�1�a�37��U�
��˭��d��^g*���Z(j@v��i�7��C�!ΞU�@X���N��xQ�<H�:UH sV��pPeA�a_�B$��Q(k9��8SY\a��g���X�Q�nT^&�0ZPGF�ԩB8��R�Gw	T޽}��o��͉���+:���c(��ץϻA>���`����ޅw �M����C�����NI�yw�r`�*cC'��)[�l�v5x]��0:���յ����>���#\��U�\�P21�"����e�ge�@"r�A\W=�$�ԫ"�A�"{����Y�<(^�s0Vanq���꽟U�h_�Zg]H��:o{f��!V=H�:�heMy��ҧ�}~J��o�{M��6���x��N�*��P�us7"q�a�P�9_dc�c\P�u�uyݓy�疝�p9����Zf�,��4*�x�w�b_xf�:�0���{Q_F�G�Rt��q�v5��[˙�Dt�O�w[H�=������k/�{�mŌA����:��D ��ݾ��*]İfk��C&a�Ķ�S��)�:���9����� �Jvb�$�)lج���n>c��W��a��W��^���+E��#N-�)��s��H�jT	�KD:u�ko9J���[���!oU�U�E�u�Bo/�hL�sj�F,Ю<�9��M=��r��s��N;2���[�>T{{il�+�CN�J:i�"'t's���ob��S��@�HC���m�<b�Ͻ�|��}��� 3�V.Q��8k2g��.i�}Dޖp/���<^�����Z<�xx:�������/8AZ6���vo��k\��T�sZLK������/��8m?���M0��ˆA~��=M�%���_.�T�"��A�F�u_��� xh�q�Xpn�׎'g�>�#�ދ�g������fT�xJ^���f��H�i�ߨp��6�C��,�_�e�U��A5�7/�pX��N��i�+�/�r}�����	�2���g�{��$Ȑ\��Ǳ���z���_!2�(a� �
s8ј�5�!3���$��%�&��t�,W35:n��IQғ����CS+oΣ��k΢]��Tk;q�L�x�<�M䶝��me���M=�;�]�V�sX0��b���JΛ�����)x���$I���rI�8����h��e�7}%����ˑ�3ZԅHd�����xW�A��Qb�T�VX�\�̐�8�{��W5��z�����(�-�#1g��0b�%WB�B����j�LŘ�ј�k�sW	�;��3�����4:P0X�~��`�+�_80������U��������$��r�? |s�G�nyee�f�|8vV:�VӏNn�r�:#.S$-�n�oat�4�Ҡ,��7^z��+���FrtGH�.c�H���mQ��§c�H�^���g��0��ЗyMϲ4�5��\
��oo8��Lc*{����|v�Kż�+X�8�\f�S{X�&��mO�<��6��>!s+6E^q�z�Y����舢�+�s\������
���6ǜ�*��q��ؘ�=e[�{�����W�y[؈��J���U_[̞�	�f��=�ЈJ��,����$���v`�����[d\�H9,ͫ�o���JԹ:̬�h]5��*�d2Wz��l}�ʙ��ͭ���L��\y�LD9W�ɉ[/�GF�ȭ����53���	�*L�rnЛ���z����2P�u +-Շ���ӵ;,�E�0zcǯD.�tR�4*(�����[
���[�m3���bJ�b�:m��T-d��rz�a R��춢�@���gaI��++e��B$J�>�t���ݨ��t�!�q*2*�HP��[�}4�s�E�����ZU~{�	�}f�T5�Ν77V-7�_�3����!�A��6W_����h�ۗY��(�j�uY��M-۾�JX�����~�N���J[�����L�p�ȷܐ��L�ӓ��u��:��imOB���]-B�߻�˙шߟzb�E�uN�iкս=m�m4��v��"r�d�K��꼮x�1�օzu8<���{�~&W������Y��ڀ���`�؃Qz��o�&���݊�y� ��W���HL�4�o3B^��}K��x�t(^�&�#��;V�-Zb]{ѱ���Pf]X=`�K�Hw6@�޼�I��=v��L����#2��;sI䂊v����j��7�f�|'�����Lo|^�B�~�f-���oe��Ű��buz;j,e	��`����#p[ev�Y���ky�Z�}�MO{xE��v�ǉ��l��]�-I�j�7�r�m�"�yܻ�O����`��\����'9k+�)�TB��{p�9^ߥ]o���z��G����Qոk���%R�Y�&3�s���*ɉ�ߤ��SqyP�X�^}]"n����������I1H'�k�f�Z.��u5��qud0yK�o��T_oL=�v�>���In���1�V
�}tbf��M��GY��⩶�	츏o���p�-��+K�ۉP8��/��f���G\v���������~��ڟ�J�TU������|\VM�������_0(fW��L��/�h�]�=h��ˌ���aBHD;B�pd�~���Y&���_��i�!	!?f��l��4Gu�7����'m���SkJSUDLք��$��~��<�_�����?n	6t�K
��AQ��7���l��H+X�"���'< "*?!�,BIj7��WBk�k�
/J̃�4���6}��Â���h��� r����" ��;9�v�p�dS�0�X�}�� L%-�`+Ө{1~�daW	��.�$BHG�?0׹V������?��I	�a�Ҭ'��^�/����tx��L3Ң�Q��k�%�_��h'��,ӫ"�nx7�q��_��C��	S�q�����6ȋ�K�0�ؽ�܃<���3�$ڲAX����ݩ�	���;/ӂ�Wջ��,4� 	���`�_a~�Р[2;��� �m�w��QODQ ��\r%�A��I�(i���!$'s���Tc�2`��_�zO��!		!�Փ�� ���ga����D�Ա?c܁�q�$�3[��V�<f��ba�Y�V`2k DTj����\����������q�=��R�G�~-�I��7!��g+�r�4���-OǼ�Q�dU�B�G�� DTv/*���,&}��ȻE�='�?PL��u��������Bc8�-�@@n�e�W����z��$V�pi)�[B����m[N8�O	l��%�ec(3�D�� 3J�),q( H;�&xR��ϐ:t���۠�ͳ8�"��uGA	XU}a�d����,��:�,�뮉�"��J�ԻAY���"�(H4�Ԁ