BZh91AY&SY�d�$�*߀@q���"� ����bIh           {�F���Й�@hdhM�h�D@�+m��ɐ �h�R@ ��kKlQl֔ h� � �;��d5��SXЫcE�#kZ������i��e�[eM�Qchj[l6f�%fld�����fUm-&�L�P�TL��ٕ�� m٬�f��S� ۱e�cRѳe�2�m2�ed�j2�e��le���F�P�R�h��kc�f�X�֛m���lf�B��63Yj��   �� ��e�im�n�*�kc6vN΀\�v���6���Qsga�����:�4A�WY�5K���+]��r�zÅ�jlڲ����b֯>H�� ��2PJ��ܕ�i@Y�*��Q��a@�wUP���

[�m\h4nոtR��o�Ҕt5�=����m&�-fմdM��Rk(�X<|�  q�ý����@jQ��@
(�;��]��QnO{�@� �ݽ{�:h<�m�7���
����
P{��JF�=�z�Ph=ݛ�= ����D�����ű���Lϒ@ �|JUv�i�t���@�ҽk� R�����Ҩ	������t;'�=Px�p�d3{{ހ
{x��7����v��tz �Tt֍5�[RѳR�ٴ>|�  <�}݀(�i��� ��{=G�G�]�p[�����R{��=P Q��vh�j9j ���]y馊�.�:T�]KZ[J��Ѻn���i� �}� B}�h=P/��`@��.( :�  :.���n�K���+oD������
(��wJ�5�\�֙f�ɢ���%��|�$ (s���| =���@�7��:Nݪ(y�ݠ�����= ����$��J�@p�{�= ���x {�L�U�ѣ4�SD����)�� �Wn���c�x�����{ATꇵ� V�S��뛀:9��4
Qt�� ���m��mR �����پ�* 1�`�|�Q�������5CGt�ht��wm�C�F뛍�;Wr� ��pU ��� �(֫�L�iJ�kJ�6Zm��ڲ�})P�{��R��U� �u�@5F�8  �\��M���Z� 50V����(:|       �  ��RU(d � A����*j�ɦ�2d �M4�&&�T��JT� @    �*jT�d     S�)(�*&L�210& CjI)��S����OI��f��zj~?����/���{�$!��	�FZ~[�ffg��۹3�.�w#��Y��mK*_|  AV ���T@~�@W�?#`���?Y��� �B/� X�d�I�6� *���CЉ�3
!�8@A?��~����>���XŬR�J�+���+�R�J�#
�+�R�J�+�R�J�+���H�+�R�Z�k�R�J�k#���k�R��k�F�+� �R�J�+�B�
�+�c��J�+��
�+�B�
�1+�B�
�+ �B�J�+��J�+1J�+��J�+��J�+���
�+���k��#�J�+�R�J�+��ưZ�+�F��k��c + +�V��k�c���k��J�#
�k��J�+��J�1�k�V��k�R�J�0
�k��J�+�F��+�# �R�J�+�R��k�R�J�k�B1���k��J�k���k��J��+��J�+�R�
�+��JŬc�R�J�+��J�+�B2�J�+�F��J�k�#�J�+��
�+��°J�k��
�+�R�#��k��
�+�R�°J�k��J�+�R�Jưc�R�J�+�B�J�+Z�`��VX`��VX��X%b���)Xb5�VXF)Xb���
V VX1�X�b5�VXb5��`�X�b���X%`5���V	Xb��V	X%`��V	Y�b���X�`��V!X%`��Q�V!X%`��V	X%b��V!X�c�`��V	X�b�V	X�b�X��V	Xb���	X�`��VX��b��V	X`���#X�ab��V	X�b�V	X%b�X��V!X�aXb�V-b�V	XVb�V	X`��V!X�`5���F)X�b�V	X%`��V	X�kD�B�J�+�R��+�Z���
�+�B�J�+�R�#��+�R��k��c�F���k���R�Z�k���+ �J�+�R��k��J��J�k���k�R��k�#��J�+�R�J�++���k���+�R���#���k��Z�k��
�R��+��J�+��c��k�F�Z�J�k�H�k kZ�Q�Z��PZ��DZ�Q� 
�1Qk �
��DB�Ek�kF�@#k� k�@kR�U+�U+�+R�U+�E+#Z�D�J��J�T�J��J�T�J��PB� �PJ�A�J�T�J�T�P�A�@����UJ�T�+1
�E���Z��J�+�R��1J�k�R��+���k��+ +���k���k ��k��J�+��J�k�k�F��k�F��B�Z��B0�k��Z�k��Z�#�Z�
�k���k�R��+��+0J�+���
�
�#��}�Ǯ��p?���?������~��]����4Zn��^bS%X�����N�KN�w]���y��pҝ��ˏU�]aV�M�ͤu=�.�^�f���s;["������˗5�kn��ɫݏL	�\"VL�,�=ue&��DƄhM�!%ӽTs&غ�X�QFU�%�'en�KiY�i�Xs]��o���[ڳ4�Kl�ѲɌI������(�gu��;���@�u�u&�j��U����*ڍݭǎ�ص�Iҷ3c��=�;��rV�G�^�t�H�Y�F��%öF�YxM��1\/~�5Ǔ�f�r�,�ڭ�Q�CH:#	Ӻ��m];OGk7e<g����=!v��!vKon�)Gض��h������YJ]9f�f�M7�ꛫ��U��u�cl�n�4��a���ȝ��^�ܲ�m��5]��s]3�h��wGf j���(�s.�I�ЊYUj�,Hke����܉j�-x�)>��	��H�#rV4m�h���q;���.�����/Rol�y!W��4��;W��2�!��6�u�͎��L�{�Yw��$����f5{����J��*�e༇|6�H�Y�#^]����BIK���6���B�!�E&<��{V��7�u,�Lk2jܽR��Zjҋ�k����pVv�H�E[T`�6��ɪX;��-�r�ՙEɶ0���[hm@���a۬i$��*�7*�*��!���H*��]���Cm��-�N
i8���k�l���ģz�po����;�//y�]�n��e����5���u�Y�tU�j�SL��trtŠ��-�y�ˮ��7�y�GZ#<WxާM�`$3Xђ�43p^x���qc�]tɧ}��֥��E��[�{�l�x�*����:Y����5#����R˥�<�Ͳq�g�sa�稾�5^-�n��)BO�7n4��
�ys6��mH�:�N�S��Z����+B�������Lm(��lhJɹyY��)�1ãa�u���ټslܧ��C��˹�[�2+�-�R���!ң[J�1-v��dUf]kܓ+%k�Y.2I/s(�)�5���2�����G�{k���c��L�iQB�A��ڭ�y[�Q(^�ٱ�p]#*��HwTŢ��HXr)�
{Dckr�Ȩ!�q�nV�6�(�s�-�w�ޒ�=)	R=*R�fкP��o,ޭ�����VV�������ij�S�P9���5o&0�giqOV�\��5�����xk.���%OI��m2����Ir��nȺ���
Z�ˈDY6�J9v�4hֺ���MU��ل�Ua�-K�N��8��DK,�u�A���΍2�7qm��!��0�2;�!n��a4�E��+*��̏oc8R�Eƥb2���z��h�C"SCw���	�ȋ���0՗�ʨ�8�En�{�+h���f0��˭�Cb����V[T�� ����wZ*�'q��8R�V�UbD�ګl�=�f�U�4Kڂ�ʺw.�u��R��N��Z���:C:�N	=�wi�� 6RT�Qj����O-9�/,�wvyi��j�}����dn��'KN5��f��u�-nuղ����g�兜�,�$�M���+�õf�SHJͨf8)��R�o%u/6��Z���ow%�s31�Se���4�N�Q`ɖi���n^ �m�n`W%���5�aN��ti�ֱ���H��Î��2������slެ(�f��A���:-8�n�O
d��'vF]�ʠV�����T�V�Q�\�������1��Ⱥ�;k��<"��!�������+C�p*��OF7�F�����UP5���F��������҂�	���=t�� �-(�Z�vߵ,�U��;mf�N�6r���w�N��r5�*<e���y�_uuӱ�u�u��4�.J�P�eu��r�_j��uV6���^+���/#�ZF�nط+rGCni�4���-��Uv*�����S�i�O�\�>O-�>�79mb���n�c�V���_6��V�VN%�kr��{\�z�O�z�/(�Ѹ]d�	j��]!���B-��RDFsk0��8uF��:e*祬�`�36Y˻8�^�`�Ile;���9�<��LV�UJb�$EK�����N�X��Kͪe).�ѫ2��ȥv������o�A�7H=K3�������i�K7^t�!�v��Wv�
���4���˙�,�b)�{��DH;�,�Qju�hlB�b�Zj���k6�*��c*mf5�f���J��{�Z����}��s��/]/
Z�w$��+k����Hm��s$r�^e؍_�����GF-��&�OFM&$F	��Hڷfk�2�V0!^�٭Z�0�g@U,L��c)�+ ỡ�-���8̗Ҹ
,l˭Ŕ5XuT��O�e9BG&�Z0�-8�Pʳ�
`��)�6aW1Vbj�v�����Ўb��ɫLע�2��ǚ
'I����U��xʧ���;�q��-Z�%!��G)٫I����n��uS�j�����wo2�j�.��Q��(K3U�渒5:+t[.����;�RV:"���m�gH�[��,9�У�-�`��F����s�+E�T�;�SU)8���V2w4:ڡKڥd �t������,�Oj���u�<�����w!�f�aN�'ucK0��2bFf������Uډb�#H3Vj�`-�WW� u-U��v�Y)��Dr�mceU7�ja��Bzo^]�1Z3i��I+`�YMh<8f�v/e;����"��R-h�V��nVFVmU^m�0�Z��Ѵ��lO�n��Z�T�Z�i*�U�V�5[���r���ŰRA*ɻ*��uT��{įendX#H�
3m�!8\�sX���w���sv�r����Q���`ޛ�ԯW5��Ô�	�[G�pumе.�X��[t�:LX&�����T�ܱ�;�˒[w�����vުD����m.Z���a���_Ԯ�sn9��Ӻ����	#1-����ܱ�F�(���N%[���G80�t�ÔA5lŸ&ZZ���j�l۲\2m���X�U˙���V%���t��vo5�!��*�Զ�
�bs.�ՙ^8���c�#[q4�{�Ҍ�����h4ʘ�f�6�[��ۯ,��}��޽Ç���%Iu�j�����kvzhL^�7��oj�6R�w�,��]cܫo2[2�&e�h����Yr͉i1t�����ˑ�(�Y�)�1��U��v���h*&�X)���1!ylKE�K6�-�3eÒ�.���4��V��#TF��{yLf����y7�>y��dj{իzɑ�y**�i��iRU�.�oi޺mY�#�n�N�5���<�a�Y��oXC�r��<8����;�Ol����V�o�;�]+�N��ǁ%<;Q'NUnx�Eb-T�A�4��'��l��(��4�US�æV�v���o	%Ѓ|�:�sS�{�F]�h�-3�C[��V	���ʼ�kc!��ɕ�!�ܕ�ƴ^ݘEU�auiXnF*i֌ʭݕV��-,T%*Ueټ�aa�(2��$���p���4��Ҏ �ּ���W�.�qYxl�:�!R[�jV{u�6�udx�
n�nӴ�Tʶ���֗[+n�V�Q-U�7�I�Wsi��[���
R[�ܵ�dn�h�jdr��b�
�n+���v�OZ�ɤ�{O^5q�w�̣����Z�5Sy^�J$u	wkS����r!K�X�KF���oi��b�Cw���=N�h���4�n�a���K��d�YxZ��2=͛T�x�fS:��r�m��J��Y�v�M��5[i���P��dCpin�J�Ebb��6�Ę��.�ӔS�K6d�5R)����7=QR$1u^�x��}+TNU��+�Xj�i+֖�`��6�^�^���2�V��X�3ܸ1����Zt�3����Q�̻��i�e\���J��$XԨf3vbV��G*�ܹ��\���4�N�n�n�߈dIe�jц�*)̍��1J<)�`�W�]���&��c�[S�պ-�Zj��7��U+[��ఱ]�kw��4J���i<덭}���^��W�r)C*R�)����y����qӛK.�5�/E�OR-�^3{M-ˣ�%��-C�ӱP��9�Uv�ƈ���mV���Me"�e�n�;��BP�6����@�֋�Ԇ�B����D4�.����jnl�&།l�t���+�aeD�t���i�.X)�n�+N�w~4i)xM��A�+�V��*۬�l�i�T,��*Z����͢�SI&���T*�w+qhĤ�nC����n̬b��FU��k<�JQQb�a�q�i<J�S9\Z\P��_.�OaEЪ�[�%���}i��{�E63P7u|�g��dl��b�:xL;dd5�'2��R�wW���pĮ#0�͕u�i���<[���5��2�W�7�Z�e��b����Q(�-���ۣ���h���H���X�NY��ni��[�-�[��	�:^�Ml�krƽT(�V7vL�Y�pl�r��.&��2���a��2Q(,#-R��CN�y&F������XA��d�M�,�n�թS�kwBŏi�����Bj�Ʃ��'E�(pѕ�ߪ*���F�-Igv�3�D�[���m��"��Na�l����x��y���;GkY�S��B[8C�p��dS�UB��ǎ����b�ŋ�Yy�.�d{쵗5�n����f�{TK�x��{n�!�dS6�⭀�7���6�����ŻW��إe����h�rK5�^�7q�l뽮��U�_��ݺ�m�V��y��e���O;�Մ��t�[[�����*m+=��Z&k#
tY��X%����	u������,�;���F��m�q�&Ԛ�i���Lt
��[�VYR�h����!�U�x�L��b-��W�.�:����y���+T��F��{Uf:�V�~�[Ԇ����O�=���<g^U왧�mᒊ���%dKI.�T�ݦ ��37L`5�8���4�GF�эS��T����]jխ���N*�Sn�꒡���,myV`�͚��V-�B����pW�����Ye�sE�I�[`���P�F鹺a5.�Sz�JL���F�֊�ز�<���}�4��\0�W�vr�mU�6�RV캵3u)���3�уv���x�`�ɕ�BTt�ywn�(S��W�2�q����E:Ş;�S"�r��!��I^ݛ���̈́�!&��[4ͅ�/m^�k�6��Z�]t<�vi��[�U�;���f���C������l�uj]��f��R�uɢ���o0�k��Z� �z��o%U��u_���^X͛gJ^yt�^�5�V�S�i؝N���U�60�a,�>{�O��K�Y���M��[B��q)�y��iԫŀ�5�f]9n��F��CY,����}C��wX˰�4[����w��r]K�Ѕi��YA����j%���.�T�V�Ŗ�=e�������w7t�jĴ0�cؖ����0Z�!�rm��c1Q��&N�(+�GUYEP�Սep����G�%�a�X۫����mQ�8�b[���9��-¯�5�v-%	zm#O5L��5 ��EF季������T>woaWu���¾�a��+�vZ�:s++S:���b�ZS$��e�+X�%�~�H�n�Zgv�ՙ�V��WB�iN��HRN��K��Q�-n؄E �#�Pg����i�[z��0y��i�[\h�/|�P���l5^J��
�T�N�A�km3�[�ͮJҪ��R�KX{�ނ�n��T��l<��V)�ꎩ[�S̴]���{WF��Yui@����r]S��Z�|���~綱h|��{B��Gl���,��E�up��&=���P���6�e�x�9&Wq�F���J�(������S���<����F�E��M�URݸ�t�n\h��Db�T�n�1�4�.���n����r���T���l��w� M�@��:���gQw����GɕE����*�m�4�ɺw�͌L{�*j��[OT�3Ay�i{��;R���.+�-^�ń<]�KR��_��UU0P4uj�U�NT����Rv�zS�����J&�b�u'w�t�V;5��=ɥ�NT��<���Z�I!����kDI$�)4�#j�m_值I+����R�n�	1S_�_,��(�"յڝ-h�-U �&�\�WfTZ��*�n���Wk;MGJ$�$�j|��K�w�"ĿR�u#h��e+�V�O2��������5���b6�~�n�j�"�s�V)ʩ`5K$�]V�j֪*��bJ*���Er�7�Uݒ�)[V�Ě��2mlKĵ\[(��ky��z*;�x(�7rz���z^/ȵk�J,�)0M+ĭTSUD��U�n*���''J���]�%\����4�%�⸸h�IlX���:p���=QV�ƦR#U[1g]c:/�����In��E��Gփz�*�;J#���k_EhȲu&	�E�rDԭSWj����A�X�b�WD��K�1Ѽ�J�v�ҵ�_�x��ű���]����km&�/Թ���Ē�W�}[�~iR����ح+�Q@N���ژ�埗�[k�ZL��(*dؓQ;��G��u/�%�mo"��U�ayIg�R�M�ʉ�m% �,�x�����I�p^�@�K��RF)��O���j��X�Z�R��4ZMd�x��A@�E���#�o��*q^�J�T�M�R�[��g��k��w/�w�N�9V̷�D�IlTC�IM|ݳuJ�i8�
�s��x����-�WZ�j���&�%�m"*��Q@V�
�A軔5t������N�\`��]i��7ky�j�Z8�Ҵ�D�WI$ڔ�W��5@TW��;��R��_2ÑKT�`��k�lQ�kuZ�JZ_���-IĚ�r��3/����G����H��YIE�����]����J��YH�.jҽ�Ӌ�yI%mjW��7mRj�t�����h�mn'�D�����j��k�v��g��'%\�Q�-�bۭ��Ц�N/|��֘������KW��� �z~^��%0r�7�v�wwwwI$�I$��I��E�'���n�m-=gRkZ�tB�,��OiQݝ2�AܞX��uuM��\� ���3_-ޱ\�Bu�lOu�\9榑as����B��.yMW�DnT�"�#����m>$�`�S���0a׉�8ঙZCʝq�a�0�����{o��}!��;�<u�����U���B󣠷�&qąpQ�tB� ���/�7g����_���FhݝG�lbF�d強9���l��.b��� �)�3l�eM�d-eM�B��E%׻3>Ve�[2P�^�r�j�^�ōZG9F;p����Z��m���������'gM�ʎ�ʉ��gn�yЦ�X[*Qn�����R���ǔs!ϧM4h]�ڂ
7p��hT��ж@�/��w!C'��i�M���5�:�e��s�pj��P�Q�1Nuk:q��[�]"�^d�t�v&2�ff������'\j*��J�(a��Y���{�)���PW<�U��Á�[���j�ͳA	�z8��֣c����Rk.maVVK\�m2���ġ}ʟe�Sn�gbY9�=��F��mx�f�z�f�4��t^��h*��{�ץ��ݻ�3��2lq�{����D���gwl�n�N����"T;�t��󮏳.+3g&ns��j�Q�,S[y�ڇL+�v��j`�ÛVeE2��vܩ`�9�>��D9yu̩�x�.P/g��h��p�TD�w�F����9�-���N*�LV��m�tؾĮ�C&��޲!Lb8I�n9+OWT\��%�k�6Ї6��r"lJXRl#E��'ooU�8z�,��C�\�ٺr���1B֦o��g1m�N���T6��q��ה֎����"�UY4�]B�Vb�]�9Į���L�^a�挂��E��: Fۻ;ݳ�Yi���;�g
.��Vn���N+
��E,�L�Z�^ܛ����Rs�DW6�U��D�v�7.��6��1���{��c�߾w�/͌6�Vr��C�.���h����KT�0ɮ��K��� �\��j[M�k�M&�CEtѸF61�T�v-�~��z��p�Cr'�����,$�54�5o�$L���m���\��s�4a��E;3s&L�I��V�c��3Vٗu���/RK��J�{��/B����m�k�]*�>�+�׭/�M�=�R�L=��1��c���������[���L2j�ڴp+"�`�2⭌wSX�@y��̃���0����w6U2��OS��vkZe7�o'Y4�=NL%T��'�^��*��H��7��ƭA�V�n�J�h���iY�O舑B�Ψm8�h*�]aϔE�C2�45BGCrۺb��nB�ch�ڮ�u�EX�4h�����f�k���
'!/J�Σ�U]bl}�-*e�2�Hڱ%�cĬA����KTq垦"J��^�!.��I����Ԓ����o4e�5oYZםN�Ğ��۔�ٜ�9����9,�-#�w^U�[�����N�c[eW_*�Շ+P�I�����[-k��s�yolى�NS�9V1�C��`�Q�L���gz@޺Yz�ݷ�l���D���R��zоZ�#~x5m�ܼJ�4���ت�b���԰�|��W�9��o[DÈD�*<�##<�2�C����ƙLlb�U]���nm)��~�WM<&m\,'��+�����G�b�
���[�q;,ߛ}��QO�a�+%D��ȹ<�k��H9��#i���T�fUJ�j�]��j���`��v͇u�f�Y؃�	:p�$�YDÆ�Pu�݉#CtnM��.�tM��mAM��z=K��DpU��/�we�w����]l�'F��kuc�W[;*��ٝ[9TB̸�Zb�&����Qi�T��T2
۾����I�1L<�Il��j���JjsY��qb����;W(V��#]R����X�~t�z��;u��{���$�.��6����ށ�Nӗ��p�r��Ȯ��BO���ĳ>���BG:mR'7y�{f�8��q{zH��%fEYU4��LOl��WkyWc4-��,������Y������9'���fʾ��L��}������>�y�� A,)����X�F2݈`i}����i����8tzp�|��t8��U�Zo7���ʣC���i4n؃�Wkx��bG��d�>y�CJ<�A�"j�����+��	06�j�ӷ]&ʽ�7�ХL��wٙɪ�+5��0�UFʘb=��v����i�����RB,v˷7t壗n��$�v���H4��i糟V����$���X��V$׈$r�s�[��UGM�����hڻ�V���1�I�Q�UP�wT�ڸ��fc�v;�V�����'!�
"mw[jTQ�ӷ�p�8�����\���c5��.9O^�mZ|[�f���Z5��a�Dژ�ws����?p�{ET�Ȇ��u/�Ӯ���w^k���C�uxX6�;]
��A�8��KN�-J!n���^c�=a��*�u�C�s�fv�AF	|�(s32�]�R�h[
=��-��ňy5ې,k�x�x��j�Ȍ����J�mih�}�hR ��z���z�-3�$6gX�X���m)78��>H9�Gt�<ⳔuR8R��bN_]	��]k�l�r�Zdd:���X7j�-['̨�¦��m���
��:��թ���d�����.p�;!��/ xE��k�o��U���铇!�8bcO�Caip��{Ֆ�cO��pvQ�]^��Q�R�1�����Q�Աx�=�\E*U�MB��N���=���l�u�;����цbx�jE��4��[�]���b�7ELׁ�Qꭼ: 媏���U�\r°�����H����[y �6n*���u��IN��{B��݄#�i79���p���Z��#�m�|#��>5,�ɕcO%��xb�G��7��\��g�Wa�uk�E��0���EݩXWJ�oe豋2�)x�h[��n�ʚ�ַũV�ef[��5j���	���.]�妞l��5�Wfn<#���N�M<�"��Z!LZ��۝�8��Ӈ4�:1��7�㘍k�4WU\��������8{ɳOJx]<�����>�\y�q�a�z��ʬV��q���N���q�k���et�\ݕ���m�s�Z�yx������2�Fi�Ү�p�m;x��mkvEݥ2�:Pw:���(��{-K�,���)ug.�����`mI�Y	�-f3�3!�����6U�/W�O�+[���h�T���; 6{{
�齁഍e�/L��n��!�"Ӓ���Ivs�fS2�U�6�>�;���f�h�}���ۄp��Ŏ�cpms�#V�ue�z��%Hf<��nQN�SD�=O5AF��.*s3�73��+FV����o;2�3Ja�u+�������[�2�!,��װ����Nd�ܹ�ANʆceQ}A�ƔSrп���Ls��3i�V/(aHU��7S�jӶfiƷ�ɧ4]	�,ySa��`�W%�ub��xӸNkɱt}W,�Ϡ�Q�7�#u���uj��,"Fq�X��@Mgk�[������T����e��E�v�;�/���''���7��X�1�L��Tr��H�w��i���wJʼTq�[�l���WB�_JC�B�+�Q�4�N���4)�%�j��;�-]IW���y�mt��\�񸔻�6�Kp���o��u�H��ʩ�w��߹�.�6��K��Gh��YoТ��L�g��bt��g�I�Q��f[�b�E��T0��ݗvtl�Y��<�d��������Z�����|v����c}$V�޵]yq�tf<�%p�]d�	i�nm�7�M��k��J�X��{��E<4��*��:��ŽvNM���N��h��[��Çn�|"��w��RO)�{N��{p����\`�խ�������\�i*rR��ӸȎ�U�Jc����ʵ�_Y��{٪k�t��(��m4y�'fD�b�p��|ICquq�Y�1��!��|�.��u�-I��R��3�50�)C9t�m%��.Z�
z���E&9���-Cg�U������+f��7Oʏh�ayG�i;N.��gjϒ����4m��/t�,5�\s�C�Ƈ
v�6���$�O�"�$�j5z��yc�:Z��ۯ�ů9)�V�܀��ɲ����>S6C����IR}�4w����������!lf���!4�8o�[�v��W�8TI�5.��Gn��*�-М�ն�l:l�c��U^z��'.k�b}�}�_w!�5�5��[$��m�!Ppr�jagUV�[5� �2��R��ͦ�e�+>��Vv�T���^:j��7�"�KV|�M��J�!�bV���=@�T�U���Q+%��˳o�"�Α������=�qen�]���=/��OY�x�7]�^�֊@����̻��=>�:ձ�����U�ah+&���{b�!�| W�N�-��^��i#�"Ǚ�U`���&�r�ͥ�-9Qk+���S��ۼǨ��)Y*� V��H���;��M���f�SԲ����ؕ��z(PR�Š���Ї7��r�SS1\�?U��c�/9&	6RN��sM�Zn'ϑ��q���F��˽{im7��.d�
�|�*�A�n�'*̅��Q���n�0@���ᤪ�:ج���{tYW��T��+��Y����9���Oq��7�������}1Gҡ����C&"�rJ�a��-���lA��X���${��P�v�u�N���<e�Haʱ�[q�{g)K�F"uL�s�"�N
�2��۹-��p�u�_ubY��"�Uq�,��m=��E������1�\�dc�ì��Dr��ۺOh��8��DɆ���<�-4��B���'�X�/3�.��Me�P�9a�G����3Ft��Y�Bq�Z�V�,4�Nk��uˆQ��ƪ�L�NtK*�v05�=7'P�م��M��d�Y��'o�um�Wlt������+��f��Y�p��3h�e&�!�W��6��T!\��yW��k��bX��pj�k#�|n�vB��z9��_',�}E�I�F��&�P�C]�:�M�{lŝg�׳���Tx�[0�f���9c��$��N���@Գ��md����.�c3m8w^�V'W���\Uh��WtR�K$�:N�`嬤�^�ʫِ�۶�I�N�Y��a�D���5-ҵ�HO����sqj�v�P���f��{F���@�l����p%SgVK��n�eٷ����_5AUq���(��x+Z{r���.����N��-[짍��J���^ғJ��C�ޣw��ˊU�-K[�T�u��m�]�DkS�75S�'�gx'D�́F�tͺ����f�AEM��ź�	�U2���t��Ì���y�p�5��Z�+���&Q������:�����O�gV��씜[b���ez._C���'O����k]�������U�xuf��)�������q��'����6M��<� �%�捹j��{pŇ��i�Ab�����Zζv�]��k�E�h�Yp�c�֭c	��Z����{y"k�����aUG,ur�"��a��]*��9a2�ձ�p��1mu����K�D����̱hjU�uv^�6��r�H����Y�y;7k�y��܊��m�t����pQ��y]�"���n�ӗ��y�a���F��7^��N�pf���YH�'hr��V�MK��_b��*,�+��Y���y���%Z��q�s-��Dm����p�s�Q�Ž�I��	R�dF�;�����L�N��+'$��98k��T�_v�5�%�3%�WpM��$M����u����yQ��tB�]�}{�9��֑H���]�K��O�N��0��L�f��rTű�:��wi�U
��i�NAó0��>��dwj����IF�V�fq�fB�\��ʼI�#IrogI�I;&�M��4��}gSr9$��$�I$�I$�I$�33333:]�u��y,��N@ܱz��w�K�T�Z�:�<���)�Yb>K�.騧p�u���B�3ɚ��)�~��"=Cyz��RG�j��Do:�Hd�؏Sɢ+�!� �H�+�l�y���T	���4!"dC�)�@}���uδ/&���P�󪯑����S�%�E=�@�s˸��7:���E�Uy�!� �%���,�@n4G��9�<Ȧ���ɐ^C�T�e=߾�M��O��͜ {.� 0�����������&���7G��'p��Q��a���EP��lg���O�����������|?�����ַ���/��;�St��\K%�Q6�[j�$Rޗ~�lrc�ۏ-�޾.�2z�<��4�eEm=�Ӡ̓�v����p�Ƀ����JeV˰�túLA�£�,u��nR�՚�waٙA��ۉT��K=/K�m�'uj����P:��lre>��J��b63��to&;�Q�b� �V[
&���pK�=姌��E'XVk�_]����i��E+۱���u
2Ŋg�T=3���9(m�OZ��c�ʉ���ׯ5,��\3i�h�j�v������㵱��d@�Cn�a��v�(`�m���0��U,�LU����a0+�PT���Ի<f#4bnA[]�6�Й�|~�	�1f�=aM��z��MEl�-_��rr����Ŕoە��7��=N5�nd��j%)niZ ̉�v��8�-�pu��7�A���,�K��n�y&јY�	o&��2w�}Ji]&&������j�nл��W��^�bb��ڟ4�w`-�z�(�0�6J��T;ۯ����x��O����;��k�q�V����\�Pd�t�]5�Tz#̡��'y�AU,Dn�{��l�ժ�{L�]h�4RyE�{.�{:<�z���~M#R���D�5����XTf�'s��%�vi�#������}�?����8�q�qǎ8�8�8��8�8�8�8�8��8�N8��qƸ�8㏎8�\q�q��q�zq�v�8�N8��q�8�8�ێ1�q�qノ8�8��5�qӎ8�=��q�q�q�8�8�q�8�8�q�q�q�q�q�pq�q�|qƸ�8��qǧq�8�8��1�q�q�1�qǷ����on:q�q�q�q�q�q�q�q�q�8�8�<pq�q�q�s���{���w��e=�ng/{�"t�'��,�<Ɋ�?���b��hw\�D�i;�Q��T��q{�;hӡ�l]0Vc�+�ڳpg�;�+6/��8/�X���-��tFu�Ǹ��k���5
�����R&��5^����x�!��Ofvu�-��^:�e�H�ˣ��){�s6�� l؎��
�0>"?�/�ު�E�Fy�BN+7U�	��Ϸ���y�f&I̒^���T���}Qw\@qa�Q|�$Y�iq�h=p��I�L�bFn*ʹK�J-�X�gi׹���}�a^Ū������G9���3�e�O#�lCrŅ:�ê\.����9#Gi�U���S�q���╗�e����wW
X�_������
��@��ʵ��v}�[G\�m:��g<v��=Ҳ�wKv��x�f��֥Y�6ꦲ�^��-jQfЫ�t����GF���R�N�v��h�mp�aQp�-e�����ٕ�S*�ǰ>�Q����_�����f��kW7{\���<��X�t���3��}N��axz�[;2��B���:���%�
s��_;R����������y3�B��	��K��{�:��jq)i�G3\�(߆�ڏ�N{3�Y8tT���[ɂ�gDs�r�{��+hT�/+N��D���<��}��+���Ƿ�=�q�N8�8�ێ8��q�n8�=8�8�ӎ8�q�zq�v�5�q�|pq�q�|qƸ�8�8��8�8�8ノ8�8�88�8�>8�\q�q��qێ8�q�{pq�q�|qƸ�8�>8�\q�qǷqӎ8�8��:q�qǧq�n8�8��8��q�n8�=88�8�8��8�8�n8�q�q��qӎ8��q�������c�8�8��q���8��8�N8��q�q��qێ8��q�zq�qǧqǿ9�ȳ�>�=�k���ɱ��¢��E`�[����[�$��a݇y�k���`۾�v@35eD�[}��j�RZͫ�m;��E<
kz����n��~�n�M��[��SY������We\ܤ1�4�#s�Q�ڸ�乩�.�,����Nv�k'o��|�T�єC��)K�s��s�T�t�!�߂inҵ*e���-=�H���n�yx%��������ާ�X��Y8ݲ�����1����J��Q`��t�U��k�[��:uF�ܓ+pY��j���uP��Yif*����]7شNGK�{�M[�CJ���R3+���b�3���F7���Y��g]p���ђ��-^<ӱ�4 k��@��4���ەq�{qTo�c��>V��������#T��vwZ��v,)6.�|Vm�Ͱ��/T��������)c�Q���k��3��!4GG-ue{�=�H���;�fax��9�v�y�0<�Y�݆��:U[s��H3�ml�6b�8o
�"�� M>�uy��Cr����$�DV&�VYj�r4��g������bWS���4��C�K��U�o8Ⱥu���]msW�,��5uÅ>��C!���q�$\�ˠ�Y�Iv��nu�(VgL!7S��FuS�N�kS�!�c�a|r�R��uVv0��UЛޠ޾�Ƃ���r�R㖨 �
�������̅�b���)������1����0���7�r���b�SSᔶ��-Y�����fh8�u�X{sv�Q��㋊�������z����c͚�n�c-�n�d#/��a���r,6�����Uv-�W������v%d�OZ�ݭk��J��[�%k-.�S��<h�Y.B2m��T��Ҹ)��Q�~�_�%������ݖ�0��v��#DT�m!W��-u��M�X��V±�Ӄw���Z:�:Y���[v9�N�]�*9x�YΊ,Z���4-'*!Yc�"n�r�*�����l��a�%U�m[����:��sm5T����m�U���73u���v�Po'ƞs�����Ԩ��׈���[2�̀YKֹ��.��Y�|*e��P�Wzta��H�Mb�nq�
�c������Z;W4�nՀ�P����7��ɺY��Z���_�U��Si@p��},`),ނ;n�Y8��Y���Q�c�:F���9jUݱ��`˭3e�m�ꔐ;\��ͥ)/opɳKqPl3� �Նg-�2_h�í��ʻ�CKB��m�<��D;��ؖ[	x��lL�3���`��UYf5e�:t\�DA�v&��pe���O"�'��M&0��=o��.����m�@�R��b������b()5cQ�3�5˖cf�����MP�fmcSE.\a�0*����e�I1�ud����(F�ŕ�����B�8���VSHl�>�p��JӡnL�1���µ�5�jh�F\S�r+#|�nP���O��ڴ_,s3���>���8)N�v�+$�f\�Ţ��Ѣgvd{�7�A��j�F@z�C�k��Ӻm��8S�9�w��:���u��GY]mQ)ˁ�5��٘+fKW��/S�ݼ6oK�Y�L�YV��^��%��T�v�y��O��������'���u�i��,:�;�-�H\Mo4��+{$�VGnOt��̡n[�,EW�/RS�������LѲY��8}9AH�=������\6R�e>ܳ6�O�|&^A"m�a*RAvJ��{���7J��Eϳ/����Ug�q�0TےS�:��r��(�t���١���}��N8ӵ��}�⏇��Y*�r�Hi)��M_�!I�n��!d�D�ڝ�L�D��]�U����b쵺����ӓG.p�5}�Z�6�(������/0�H�>���
e�u���N��tzP�C��k*u� к�{�-��⁻N�����rrq�TR�*�`�q_"��s�d��yؙ�B��ծ֮�cZv����Rþ��^M�4X�ZU�S�/$Ǻ�#�Z��_a��3�G3œo�=n��=M]���[P����D�;�+h�c9Q�OM!uխ抢��l���[�R"#��vn��%Ox�4u+�).��:.9�"])��d��Ϗe��Y����60�__Va
]a���-�l��"������Գ�^m �;:59�ci
6��*LS�i���:��P��6�>�8�,��N��޿�-���ŗ@�UOkn�T@c��ܜi5r��h�����������5�uCx��Q��[u�Lӝ�|r5+����Z%�W�ɳ�b1�+���Ź�����Y{k�ݚ9Ь¶�[H��*�٦h�V�tOi��@��J�wC�L�z���>;L��f]PR�ȴa������B�]�z�
���̬����e����È��޷�ݵ������#BŚ_
g�.�"ё�U/�B�M6�sܻ8^orRY�V]2��7*�{�j�#0Cpmd��R���[=��oGt��3z�<���uy��{g`ԷbSv�]�T\�M
(����W�6�.�aYo�������ko��gDǷ�:�4n��ʎf��R��i�L�37��i�iVr�ˍ����eb�yT�;ؤ�V�ʝD�C�8fh����ZѬ-�]G��õ���V���O:$��*���I�k&���7E\o3�]Is�T�gN���ûu����nV�kJ�wn�)ݤ0i�+z욭Efų�V�]KU@�9�T0�L;��ں�U�4�G�5e.�q��T�����oVܽƪ=�Q����qg4M���;�ܶ7��"�q����ͭ�fU�5�I�Zν\�����VPP��B�\]K�7;&���l�!�q�0qX*��Y�I3l�n���N��6���s_w�A��]:�+
l�՜&�c�b|*�6���6���I�N�MU��vb��m�SL�qˌ�]Yj�>������az��}cnu�Jк�gR��/�,��[�+V���3^mmU��bεw%r<v���xt���M�Z�F��!Uj]���[�:5��2�޹�}-"�(D�[�ivp�����U�s���:c6z/��z�{3�yO�>�c�z��'VoX�EI�umU�=�V�dOz0񷷙͜�Bm<��x��l2E�E��tp ��7e�iV;��Φ�G.�l��o9\B\������f�>]2]�]�r�؈,���\u�
k����wvV�I�%̹�j2��b����ua��O�8qpc$�X��z�W��z�2���Gha.>�=J�λY:�n��D^�Jk{fr�gk\vVq�O4��!�=o|b�x�}\*�}��j�v�v`�80һ�:c�&�2�'1��	oۤ��6��߷��١6վ}ɻ�R�aن�)�)����q������s+�o�ϕ�*�"AW�m�K��b��Mɔ�J���!v�b]��7@ͣ�-g[���)
�d�]����[��(����\Nŕ������0�"�=��x�\/2L��޷�c�<v��"�%f^@aa؂��C����Yt����9V��4�\*K8k�>����Y�p0�w�~�݋:���c��5��4��1�#/#4O���LUUص�B�w�o-�n�}�,N�-=g:��<r�"0�U�/�]Wn�H�a�M1�*��%]���Lv��e�K)'.��	VQ?j7˗��
����*�Ac:a���;kjt���{�QB���:HZ�[��]�I�����M��,��٦�I�i�����6�8v�`v��T�a9r^;s^��♗ه |G����؟�:V�Y�Țz�DW^	��^1���.��0lG.��*�9��fڇh���9�]S*��Ɨ��Ɩ��l[n�a����\4$��*��%�V�sj���gr`sq���;5!=�39S,��}�*�zb@��CZ1F��? �^N[-�ER�F�%ރ��<��_.��������՘XY;�	Ty��8�	�Q�E�߮��mZ��>��{A E'��N�a�f)ihԠf3�U�Xέ����M����S�A��En=��*���*>�9����K�+������u��<gE����0ڄr���Z�:�Q7�,���*��<ՓS�SW�(�A�+�Y\;���!-��Zʱ���.XJ�n-U�mL���K���[�v���W�E����Z�鼡����*�;�bm��ϊ5&�2�<ՙleR���,bX�=yƕ��1^�|��5C��w]E�dƳrw`���6�Y"\�>�MVR�jv�"M=FYo�fo��J�l��u�Мf��G�Ž|v4�+; �`�ҾD�
5GNJ䞯���Fo-
�$j���"mU��jW�,�Gt���<I�q�U���R�n�Rr����S�9���Jc��s�N�Eu��&}�ϡ�w R��e��V��U�̢a�[+Osa	2�tWy�&����Gwh�H[�r�i;K���u�IJ�N�,�����-si���Sw���C9U�Ƌ����VIs����e�߀2{��;>�.�FAc&��8|�o�/��Gm�8�u�
О�E��4w���(du|3(�KN�y'�P8��>d�q�Q�6s���7�]�mM�-�R��K��L3��i�{,���[���E�|>Țve%�_uVp5�Z�\�j;��꾉�
I��v]Wk���Lוi%��Ҕ���C'�>�J�IY|Pb�BKܽ��u&��I겺k0�젝D˽�n���KpT�٫E�������.�N��Vp.|�f�TD�p7�엃WuIy�,X����Y�4��{�FZF���|!��&������]!�3��DJk۽'V�[�c,IX�l�QٮZp�&쓐M�]HT�:��tg`�T���&��uդ��y��ѐ�{���i���<s��v�}!��{�Kh��[�x�*��}��!�%F����:x�[�Fa�Zpd��? ��Q�O;���5OJ�� �.u���뇅��(_!AƞL��Ü�4MȮn��fa��t<ˬA��`g�9�i�.��&=�u5T���'K��R�iW�+��+��D�b
2���mN5o�:".���-Kz&'��%)WZ��D�Ҷf@�b�J���.��?���P _���_�������~�8�<?���/��J�3b�%H�e���1h�i'IQ ���U(�@d&HX�G�V�5-)pE��bB�XP�J�m�BiE0�!a��l���
,#IF�H9�tjJN��iz�f�f*L�(C�R�@�h�ԍ�ZF����R(h(
�@�H��(8� ���MƈHW��'�9�b�D1T���g'�BC��ALQ$�F�5H�S�Ym�������'���H|Rm&�M'�"%G�[F��=e�ہ�e(ϣ8���fX/O݃p��b��+vQu2n�Y3{{�vU�� �;K*��m�(�Rl�ydF�^;�eWlCE����y�엓�W�ۗG�%W�J�%g�NK˺8��C8�U�	��;��ƻr�����Bx)��}B�P�јt̕6�W-�K��x�������F9��7��������;o������u�v���3�W{��P:X�Ta��[�3�kv�'"L���5W6�Zp��������\�:��j
Kr�UR�$y���G�x�<T�=q=�l�yA�f�޲�A����V/��R���T2�Չ!��f.��Ancq�Q:ɢ�<(�Z��Ons�J낹gq��net��D�k^�C[�IwJ���ʨ�km��U�
�̦3Ye9׊a�ۻ"�T���˹{Y��:��)y��^S5N���\��&0�+�¯s�k98�g��p/���;;�����K�1D30����*�����J���oBD�X�Y�NlY��OK��wX�r�kEV����-v��W�xZP�xc&܄�J�7e��9HlS�̻��Hu�K7/駷rht�<��fި��F�ԒB�G�I�fW�� ��㈈��^Q��`� �0��f�P&�-�8K)$�2El"����&���ȑp��p8#*�s�$�EFd�	�N@Qo"�*�Q"�ix�E4S�Id����Jm1�I�fH�9$"�@�e�h$�a�0�F�$���x�\*
pBI �%�,�"�6�n1faq[d�$�$��`��i��&�A0PbF�(��$�d3$rH��3-&RM���. �A�<�1�	$�gɴnB�a�f��1�䐠�H8�i4d&
%�SȂML�[�y��EB�I�ID��4J�l��	����M9#Q4�.7�R���I�j?������RH	7p@�0C"E�"�&)ȑ%1"LH�09��`)�QJ@��&c1)�$��ă��q'!E��pS�9���!l8#'�8�p�B���B�U!�9
Q&c�n@�*L����甌�ƽ<W�M�!=���G��F�yE��m���m��g&_;�����χ��tj�k�����8��5�q�|pq�q۷nݸ����:�y��&j3���.�|�<O�_m	Vڶ��ՖQ۝^�>><x�ێ8�q�q���8��۷n<|9�Kyt�$��Ci���m\���/<�.��v�z�?������k���ڜ�ۧ��ŧv�3Dghg[N��^�������ŗ�n�ά�#0*-��.'�Q�Z���S�{�#��ƻ����ʴ��; ��}�:����m�~+���!~o{t��j�8��Zy��S�N�vJ��^q�]f�o?yw_;���;������m��e�ۢ�����j#��_��4��RG\IG���;u������ߏ�����q}�[޽��j�֞�l���.jV�[�y��	Y�Ӭ��W�C�f ��D�k���t�Fժ��y����ཿ~��C;_+���m�no0�s���b��7\vK;WfRڛ����{km�l������̇/k��{u��}����Z��N�g��<n�����y�&i�kj�[i=�ֵ$-�d YE����A}v�)!	⍆�&6q�m̂&�)��)&�f M b@�7d���Q�|*���	�Y"�n���K��֒-��4��U���˱y(��hO-���Q��*e�;��8�4ѹ�e�
��\�20��@[cN�B�Qm"�rXe�≈[A�14�a�I���&�I�R6����)-7 q��-�E&e|Xj�JDȑ�L�OP�;��c�G�^�w��]�kԳ5Ţ5dѷ^$�A,Iv]ܻN��H[���9|�>QdRM9��v���3�1��:5��uyӒ=w7{�HyPyO����{�s���H��ot��[m�5�'���7���W��y}�/l_��M�|䜹7�n�Й�jn��:�������V*{��=����/�������o��Ls�d�$o����'���5�� :��k�k���إ^�o�Ǉ���Q�i�I=�3���w����<�����-ੂV�s��)	����9luI�Ot�/�a�ۍ���ۻ{5�\��/'�>̚qL��vOL��ϕywg�K:���O)�.����8�?w{@�*�$���D93�~�E{�@c2G��1�MӾ��3�0�6����:�b\�c7���.«���Ͻao Y�r_ۼ�Y����ש��k�)�ݚ��1(1�Oj̶ib���[�ݗ��=��v�a���D+oL��n��P�Xrey��ri앃%��Z"�+vQ����5�e'��p]�K�et{�^�ت���=5Y�z�4"��\`]/�w���~?�ގ�SfL�~V���@����h���q}cڂ��~�>���D�ۏ��"z���g��SW���d�YO��Q^�*L�Z���S6��ݼj��|⺡Sc�^_�\_�<1 ���s#��v�v��<W��g����Ϸ�"�������Ò�Þ��<�WU���Lи�֊��� -���]�1d��{���qF�Oc^�ַs+Zm������xL3I;֬��}6L�y�������&4<I�����s��#�dl��$U�L��g�ӷ7z��<ؤ�����o�K���v����g�r�I�=�B��#�09_؍X�Ǯ<�����C�H�xܯ[������C��c����d{�����%�Ƴ�X\�=E�E
�=�j����ag�zK�ٞ�T>��g�ʾ�C��ݞo�.���3y9�)��:l���;a{����Z+R�]1fY�E�_\�JX2$Cl��c�]n�Dsߏ�P�P)}C���s&ڭ�ϿŊ��KՃ$c�eS��챈T��Nŝ���wc�'C�{Q��ż]�O��.�o{���||4of��9{ＰM�K��|)��@ y�1�'H8Ns�����|eU����̺~�B-�}w����x�w�h��-�QІqK��=k��/�}�q�:�}V��|�q~�����s�޽m�ˇ�GO�'��海c�:�_؀��a���@W-i�^�[�Uv*�Ҷ��FbưP��E.��_�y�ޞ%�������R)�A��w�T~����!H-#����V��B����ṇ#��^lAB��<8u��}�ːLJȆ���yW���{|�����Ao��:�_{���K>�~�����3�vN��8Z�J?Gt7w��z��0p���V��>���H@LM�6��v�'���;�9�R�p���Wv1�[=�aO�֯fԘ��f�`�Խ��]Z���T���]{qH�b���vŮw9m�*�l�"vx�1�e��ܪ����^�[�f�`[����]0'���w��'�v�I�Gf��!gQv�"n�w~��-Pq�~����+����E�)	����t���}�c=:��n��~�Ւ'D��(�c.��^�yߤ��o+�N����_�(��;x����{��7��sٝ�F�]�H�oш��zāy�-�[���.8���T���3��|���=ès��>-�����n�Nh�́��n<i�L�y����cA�����l��l�m_�-V����{���~î���~����oK�����u&6���VY����;�4��n�; g��ο�l���V��T�s������6	&w�-�c�0�88�K,�3���x4Z*I���~�=���G��w��Y5c5}�A��'���жo�$�F���Nx�?7��{ݣ����m���Z����������`��Xo��g�{�ԶVɊJ���0`XnS�9+�-"϶/Z��mך>Zm+c��טF�D#�VwH6��N���@�".�\���[β,��&�ڼ��[�>dX?Q�׶�(��fu��Y���ɻ�!����3ܫ��k�me��J��VS���:Vǝ�&M���n�7RN�oV�ޮW���i����_[���ެ��$д��{BsG`�$I~З��3���g彵��3�����H��=�_�N���G�y�}�yό�0�mLYW�/�;�����e��>B�Mq���ɓ={ݾ�=M|��[J��Yo~�C�f}�/}�0� Z���ۇ���ϻ�S^���[�ͫ�8��������+�vor��h��އɀ'���@����Q� ���^Z����p��6��Qyk=���Ӆy���=~#����~��C��=9��H��Z�-UvU7�s�{�o�
���������AeyRg��<1�ټ7T|�QI��O}s���LP�9U�V'�����3\�������a�z���[I�4m)vI�s�{��yv R�j�ʽ��/���h���mS��]����.r1_^�O�x�{��&ȓ������K�d4��ûΝe����h1�~�En�WxX�]��`����N��<��ԣ��\Y���v��\�Q6�y��'L)���Ǡ�f�+���x�,4�܃�%���X���]j�$�7hIt�DJ�#��IT)s&���Z�18��s�+&}>?�=[�L[��|L�捳��'w��H:_d}���c�b5�[�ѥ�Aן{�3��'.�(I�ܽ��y�sP�{�z��_�MTZ�+�K���@�P��PK�}���$����ޓO��U�����OlX�� �H�Ϸ��u�%	�)|v�������v���/&k�&��U���M�.y��y�|Ȧ�W���Z�!��4kys2��ſR�ӫg����u�ď0�W��@�Eo��M������+3V�8銮wf��97�,7MOp���CŴW7�����������E=N&��3�O�un�g��=�8V��TqN�7^�G5�=�7�^�W�i���Q>���_[����D�4�M�.��[�w{�k�!��	���T49[dl�j�;��[g7���y�.um��t�rS��e��6Y�Х����3�&rl`��|���ʶ�n�ȫAك%@�ĉ�ĥ�Z6׎5ّ�#�I*/)���*#n�Dt�E��b��,��s>�x3T���]�i��:�-UP�n�Y7����xڥ�t��>� ����w�gF��F����6)���������ؼ��Z�O'x�$��>���x�ho0o3`ޓ$��r5X�k�������
Le�k�����C$�q��߬�$�6Ս�s?:&����k�^��M�nx_��y��^��$�/�%�`��]���5F5����n�z��$]�����P> c�������~�|��W�}�-9l��a�ݧ�}�߳��+�Nu�3ꥮ��W��&}0����	�\��P?lSVo��7vWU������/�s1�Fc�����߻�̝��ZWj~N9��x��Н�K��@�@�����W#���~''-jz��]
�k�#2�[#'��ky]�/�/�~�� ������[�ˋ�ļ������'���:��H"c`3$�s�~�E�w���j���=� ��ܹJ�vL�/R���̡LؽTS��5�pF�S�P�|���o_���8�yOJ�V^|(�����ic.u�t��n'��]��1f����M��V���1N�^�-�$>���P����B�p�a+xw�������rG0����?O�=]ݓ���l ��B$����$<[�fb��L��*�b�x(k��/�g��M���l�=�.rW:Ow�w�����^��\Yj��l�$z���/D-]��Z����~{���={�ra�^�>ߪL�վ/k��J�z�%�\#�W{��ei�n�&���g��ỽ}�� ���v�z��Q���s�X�{�=u9�s����M/�������~�}�=	[�����{���e��J9�8�J�y]Nx���+:=�N�y�Q<Xǉ���s�)��|���MɊ\�G��c������47�4݂M�~pK�l��4����N[~���
����u���8�����E���N�q}�R�Z��K�'ɇ��敏�"��e��Q��({���3-��ai��APpT���Vt9ޛԯ���o<NU(�����^w���u�'�b��+^zo_&	ԩcZt1^�u|.����&���U�3QE(ˆ��R�{AH��C�_���e3���	�;%��9�e��N[F;�3���� '���Ψ�d��|}��L���tM������X���c���7*�i��y��m��jw��Yړ�G���$�]�e���H�͊`�N�>rox�I�ӟ�E���]"BO{<��{5~��� 	ߏ�=���e��g���� }��x��ّېH�����P�;��{�g��I��޺*�W�����V�˗���8ǫ��~4m4K%y�^���hfU`��ߞ�X�h,��w�2.�3�Lطh�����lcb��<�|��%<�S�#�|�{^��驪o�yUb�g�������<޼��"��y�ސg�J��Vm�T��/3�~�iO{5+��w�'>�\�=6���gW��ߧ���j�<^m���z�*���vO4�8�M����x�N��xf?{ɾ�~����Ǯ�
��b��8�k_/k�
�W��,1&]�:���oh5�Om���V������B�QPs��j�V�pZ�R8�z#�TMH��`?�b��j�f(�5�6JOT�։�ڣRW������X���꾧.�dó��aY])]F�Oac��Q��z8l�oKGi�.o8�;3!��Bɨ��O���nXΙ�Q�i�;P"��~���y�13=.�z[�XW��eK��b���k�ۛ� �M-|��8�������`����/�B�Uqf��do����v�����~����&A$����NguHrq�����݃�Y���;c�w�4߫�ɓ��&̝U s�<=Yz��U�8}���oˆO���!�`����&�k�}&����e�IV*שּׂ~ʽ�&���T
�5�`]7��{r}�^�y��ϙ,a��3~U��GS{� n��,�ua0ó�;a�˹k�ѺNP'��^M�t���L�Z˄De��è}����Fy����;�D�咜9�[g�8�C������#ׂ�̈́������`�X��xya�5[�xX�c-�\��o|�<:w���/�zy�gg����ڊ }����N����.�{>�ӹ���Z�����Au���#��6z:Qb��u-�2��{Ԋ�̣�5�:�5/ 葆ݮ�g��o:³f����9��5����bh�P��|�_s8���t�18Y抛J��Fu��]���bP���+��%k}�K(�[�js$o��{�+����b5�F�����GA�+��xırvXyWD�E�%Kj�w3�p]GFO*�z�41,'6��ȽR^v���:�N ]�ɈՌ�	��:5-�L�8Q#5��)`�Z0��6�Z"v��fJ�Akb�\�2B���3���E�%"�ֳ���B�sY�����d��4��s���匹Ո�9՜�9�.���O.�1qܙJ�6Y��Ky���:tT����NG�]�b�|EqL�*�*�[���3E�d�R���v�L1P%��V�nB�-+qw���3�.�*w+�K���n���I>��B%ro`�"�j��^�s�UP@U��"�(����nBīZsҥ���'i�/^46�;�xpFBӋҶ��n��,��;�aWlt�-��J8�u�ۭrɮTB����n�B��.a.���{wV�gb�����G,�q�]�h��,�>x��R���K������q��"���B�d,ۖR[2��%ZOdz^t����k#Yt��9r���NMf�%eY�;-��'���sk,y�T�Ȁ�"�K�M-Z�/�	�/MX�W��ƫ��c��0�\\Yc��闯�v�q�Y�������d�Qy�"�����y+=%��Q��rά�r����.V�U!u�cr�%���p�Aڦ��P��펇�vtD��5��#��5v((�;7�.��S7�p+��J<?2��C�՜د�*�d�mX*.��6�"c57R�f��0U���� ���ˡ����VQZ2J������i��=¦ow)���N�"�HkY������2����-5^.N���Z:��yx���}��C+���/5;u��X��϶�H*��N���=֡�W7�հ_݅��'e�Ԙ��1�؜�cwETSF�/S�f��b�uA��n��l��^�Պ����ӊ㽗����]�V
jj41<`�;Yݐ�z��'ޝJ��an��v�oQv"�*�`������o��n7z�n��n��y�V5Z��I��wO��7�g,έ�i�Υe�b� �N�k�R��c�:R��܏Zt�쮝�g7.*��oU��.�K{xgnu�7��w�S��rJ������]���u'{�\ƽ�M�F=�k
���'�#rKi�#*I#�$�M�F��94�Xi������ l��Xn��T���ƛ��k�i"HoF���}�Sd,�zޤ��e��u{����kO���w���ӫpq��D�7S���ӧǷ��^�qƸ�8������>���t���Ǎyɱ
����[m7��{�S�S��{���ښAG?�޽��z�{�=ݖ�:��-s�=��Y�Ǩ����ַZ�O�O>��8�:q�qǷc�>��;v����ÒI$���U�����ɠ��9Gc�j�Rs!z�z�޵���ݬ�r{n<�v�����㾧Y~z�����O��oZο��ݹ�=�A�����m�u��4Y�4��ڐ����ݟn�<������n������xwӳ��מ���߽�:�5�yN��w�#����JH����K��󼲾]��kN��t�����z��艛�����ѡ~�9���J<�����}{W�9yu��I�Oռ�"�B�u�<�+�^�?��� {gmnG6�Ύ����~�w������~kN�9�[�^�����;������޺�۬�[l��g�'?Z��0���n9=�AN8�3-.'JP}���w���OͿ�8:�h��(�
S�D��d�q�~,�q%�~?� �I��W�'�ח���X6o��ٕEN��I��2f)qYER�������7ҙ�X���f�Wd͝�z�|ޯ8������Vk����X�ϡ���Ad�����V�F��@I�	"�&��8�d{���y��,���\���u2��2�����Pp����M^�L'�/V���>qw]^��$�s�H!r��׮�_������J�?H �a�DA&e���[���=���H 5���
c�Ɩ��@��ӓ�T�Kͽ4Z�P��e@��	��,����F�z�����X���b���RO��`��`xǤE�=q��D��S��y���nHe�;m�w����y��j�LK�Y��M𚉷�$gA�zi��f��v]�������`�N�]W)��j�A�C�v%�thNxd_�22�%*AGc�W=���{o;H.('����YY�J�f����xam��� ���	}~��=��Jr�	`�&�~�d\:� ����/m�켷������!�M�g�&�R*5��nOC�Ou*�|�|�)����*,9���N��ȹV"#q��]�z7m6��+�^��}�3���и���cn�/5�]��M�jL�~ZH,n�r�����V��C���53L�{��]��=�*�_�/�?r����B�t.x����= Ň�fF_;�lMپ"q��-�9p`!��{�k�(oV�O��{�s��j��]{�¼�e��tG���/�-Z%M��q���*��������ܙ*q�.
���Y�F�]��g�����8Z]:<��A��si�z����ǟ�����dv������g?�{��
�J�0	D?�l/�Aq�{��@��A� T�D���*�;[���Z���-���q@����MG���e=W���p1L$��y�_��w)�2ӥ���{7�ؿ������8
W}�?��(�a:��o�������5�K}���d�*��0S����]���J�>r��v����|�6ddnO�8���
� ��}��j�E�&[E??G���t������#�͉�HM�VL����aq^�/^&�I0]ćn���Ζ�����tF��VV����X�kܛ@}����6؜�����Њ��`	�����t���=�+gfi7�3�;}�~kOÞqz<	X>bO��՟�,�잪��������Jѽ�G�	B�Q�d�|B�ޛ�l���x��t�ӼXP"��p$Cݽ0WW�1���Íc�,��C�y~3m��l��|��%�$k��c���T9oP��h(u�12�]T]$���F�>�@^���?'xO#c�l�c���G��=���Z2%B�>�*?��鿁ϙL�������5a�ɻR��ى�[8��Tt�Y�2[I'\��/�oi�18v�j�5�y�g��6�y5�@�0BA$	�8j�Y�ޭx���vE��\�ӓ�v�Y���ܛ!�k'I;v��*�!uֈ����9ӎ��n%V�����///o������u�:�6���\Z���>{�.U����P��Va��7��r����^YE�����# oGB����m�8V�ml}��r^�ħ-�K�J�)8�cV�U,�)l���q��H���	�����`խ�������C,���`zΩ��&�L���Zq�Aw�8����4���u�<�^�u��EP��,��v��W�7�{�b�>;��3��u]H#��/@�y�N�t����̙v���{OV��~����� S,u���	��K��&h��\��P^+a�0���r#�<�T���f�͝���G�����+�.��o�YQ��( ����@>M/��(�_�����jvR6�����C���^��u^��{#��~k�J�a^Y�̩T�/l��Ӽ{0l5��]�v{e	��۝gp����P`���]�n�2)WD��� ���������P[��F�>�z�jj�}v6f���C���(}!�z��3��i��]٘v)��`���J�ߋ�ֽ���:�܃	��;3=��\���C�\-
���X(���<?%�g�?�i�>��v
��y�_���Ԧ�6�%I�[���E��o>s�;6�`E��3[qL��^]���'�/L��r�ѯw�[1����;aS�Ғu��<<\W�$x�.d�Oo��oqh���Rf9�^��jv! R<�x�8�K�H��PB^�	*Q0���ɹ����*�� ʹ�sQv�S���	7j}1�U����/��>������3*�q�#��ɚgy�l�O@��A�r2�'D[H׊xn�����d!\A��P�����;�x��g�Or��-�]�'��t�M�U�B��O�6��87�g�3j�̕Wz썟�R���<>[��L&�H�~
�xG�+�D�R�mS
�t��HZ���f������a^�(��jXw�]=Ô�� �0��#�Y4È�-lZ2|��%5�dC"-�P}bd��yJ���=]ڇ�������T-U�e+(����f�m M��x��Z��u��-��MڬṦ��I~/�a��	�T.�g3}�l�逷{�`�1�:��p�ɰ_@#��ͷq�F7N]��'���`�B�,g�O��%�E�<�H�%8o?E���������	�vp�=ClL&��r��
�/;KL�f���8�> �	s�]���E�xr�E��L�oP����7�k۽6��y��좦Uf�֢=���Bl���F�F��wqOK�Dŧ�I�J����k ��?i�[:�����94{a��c;{Ck;>��4�ؕ�"�ˁK#YM�w=��EPt:�Ɯ�a�%�km�:v�Z�#�����&�Yx�K���bΚ��4v�i�VW<�v���a/�w(Y����+ik���
ּ�}9i�
�ӎHi���C�u�/���/l��^t%&�mWl��u�|t�d�^�g�y��=Kdf'���zaP%��K|���<Y��.#'������g>�'��}��ܥk�w��0���Y�oX#��UJ�x~���]�����ss����qp&��; ͖�,��"g����e�=��s���x�xǇ+x���z1���4��"G8��@fp8�ޖ�A7BC��A� 0���Η\O�{��ի�lr���.5>�<[
`+�@�[��Ah��],u]U��%��$1���gu�H�^8wg�s�zj���\mT2Cd_U���n�/@� ��gb��-��^��r-��+���{)u�����c$KN��O���ܢ��ލ��]�H�v@-^cee(R]Â6R�kwg�M�&�p��<��Q}��ہ�<��t���{�NlLG=4�$�u�Y��5�����,�����U��k�����B�ٜ�{��AM��!d���Eǥ=�=�>�c��"r�m�)����S1. Pа������z	�Fc��n�f� `\؉ar"���:��10ٍg��Cǟ���jt�$'�KY�BF)���#�-�lm�<�ۼ	
�w$e<I.�����+��@��Q"~���߶�Wh!Pk�y��_�1��p«~�Y����vD�Vy�Q�.X�UTV����L�u�Ө�>�	���cߏLF\��ųT��j|��A"��7ai�9�$8:�I]3Q�P���<����������t���\����H����y۝2U��)9J�$d�2��(���0M�����]b��({P�5�4�����X)���zH��V��M�t	E4�jB�^�mCcim�j|�ռ���x�?R�.~O�d>�����j�|��9{�]�ۑ̥�zO�ca��#hw�m�g���Թ���@�S��p�<]���Lh�Ѝ2ڟ&w/~�Q�Te�Y|ǵ:���o`Cݞxǖ�X��1����;;�=���!�6X:�vM�&D�x�6��~��L�����C��ܣ(����pB�$�Z��x�O�j���b ��i�[�}�>��r�'f���q��x����޶^�mH�]�6��X����2םx�c�GP�l�`ۈ�tҜd��zwN��r!�"���[��2��ԋR2w%7���4"�g�m9`7	�6o;�,���S	�ɔ�>(�5
M���C��p���B�tIz& f,��g�P`T��u��G��Q�EÊ��n���e}[>G�B8-q�|��7~���c��-�38���m�3�zTGMܳ�H�6�	�t�!9QкLӮ7*��n#Wl�����y����5{��>��
X��8"\��m�vhZj�����*P��h�_Y\~�Y#�\�6r�#��X�Fʍ!n`4�1����q�����y///;���W�C���}�����9��ea�n��T����os$��R�Z�6�~��矗�%v��֋Q^���~����m� =Ų/sp'�Ǆ�;<Y2r�_J$�C���z4��zގ���co�{�Jn�<PΜk�Ο�	w�<"ä� ��[�P�u9�����ջ\G���ޘ(��)��N��οJ	�8�K:m���q"�*��k�g�rH�h��[�Yy���pH?�9�@{�3���Hi�h���_�+|�ҙ\�B��=J�(9���Z�HB%��}��?��%ש���oB�"�	��m�8@��Rmky�Ľ�1)�FB{86��1P���=����7��B��;8�T:q�C�lY'��3����7z���Gt�Lm�lLqd�vq�C���h1�E���
\�[!��,�3~�~xVy|}�mÞ�;+�w0vi;fWY����x�s�^�s���@Ⱥ��Z^��vo׷zhA�ǐ!�2�T]��'D�iW��ޡ��-�(�M՚L*�I疠\��XJԩ�HO��>;0�L��Xm�+��<CcB�'�>�N�jG7��8���^N.3��U��`Z�X �kL����G�au����3����qM7�}��b��@�㫐��Gv=�S�Y�X���u������z��������WuZV���ދ�fa֭����HR�A�RKn��;�����m;y]���ո�j,��9���G*.}���//!1<쟻�q���,�C��7����YV)��:^|�	�\�_�����G0����#��f#]�z�b����mz|@@�3����=�� ��M���-�8�i~܉�g&<"<��۝6x|�f��"j�x/f�������9����X<h���e�C�$�n5��!�E��Y�Juu�7�{�G0V�y���1�%����4:���yw����\�b��7��k
��U�����\��G1�r�=ۉ��ov�Afz3T|+L�H:��N� uc>$����G����묺�.�:�u���pn�EF��З�zk`)��Jw����\���r4<�}n�@3��n�hh�c��YuY�ڐ�63���C��Ob\GT	jħ�c�tʭ]II���F�"3��}������*>�j���O�ŗc��k��=�Y��	����R���'����w{���oµ=ۃ�]��U�hٌ�`�c&46;�Pj��'yW!���\���=ĈY���RX&�	}B��fb��+�FҸ��_~YB=�_�jU�֧��cVO0�p͙��kةa���aZҼ���8�%��z�%F��TyZ���v�`��m�lۺ��إUQ�7s,�	��P�2�|��[�slcb�{t%�٦Z��L'd�2��VvKo;��Ը�!��k	_�L�빿8����w�����1�k~���9�+�;��L�v}��ƽ#�'X�%�{uz@fTJ�
�|ᮢ���q ���]e?-�}̵�ٺP�ka<�K�Ϋ��}'={�,�ag�Qt9�-�C�{� �]K��6?�����]|�����"5�?�6ྑ;�~Ȥ�,݆z^��O̓�Xߊ�P�b�a�h>��,ε�zXS)؟4`�1�x����}q�������n�]F^���SY�)L�s3�F<�C:��s9���!����g�7��]��8>"������W4�}��B�
�n�0�l.�z�o�.�z������=��s�1���ǄU#+b�>����GO����:�1��}���*��B��Գ�w���7�NE�K������5���{$O��3�N�f} �E�!RI����7B�7;��{[[)З;^�����z��Ή��������!�#��M�8�]5gm�M�]�{K��@{.^�z_+�LG�fz���4��/D�GN�H/������^6*�i�%�Cn�����hx�6^р%��ZH�_
���fZ��dWu�"�d�4
��."aMT���=�,���z
�gDy����Y���eҿyS���/��d�h�����D�_+�8���oc���@��鸡�x\hMz��B��j�i�8J�!��{�i����ZH�F��O����w"}<�<��/$�^u�O��k]jk:B�*.::..98�#�����ݞ�o�w!�/��
ȴ��6����a�C(���ǣ�E=01$�`�l:y���S��'/�{9_o��=lP5�$�͋OmL�H�x���� �؋�.���mYM����\�vg'��γ�G�_���cC�b�OK�+�03z�Ui�Uh��>M�ʰ��b�Tg@�А�,�����<_�#]{�g�P���c�y0�LK"��FR�T������Ο=��O��e���܍��x�p��S��,^��"�W;s�M��ħ6�L��*Ml��!�c��z�wԗn�!��0弁@N-���"}����`�nOC�wJ����b�7H�Yɥ�1�S�ٳݺ��5����gB}�?,"�~~a~��|�-��V�����/sa��<M9赓i�=�O>��8��(6�tz�����]�=�*�� ��/+��a��l�,��b����T�^�u@��t	��a�t��0	*���c�H���ǆ�޾��?d.9�vu�P��}����� �{�]8r��ڑ��/n�1�3����ŏxxx k�i�{�"i�]��c��>W"������j`�s]ے(;��E5�*�Q:�t��ѵH7b�Ū�\�E`u�[P틩�<�
��[yټl^�N��wr��>�����PE�Ue�w�	#��ww�"-�}��Y(�D�I�z�c2b	�]��2�q�+4���"�u;�������6֛m,Κ\�8�0�tN���p�]��w�]�V��G���UK;+���Ge
�6�1��8#�o3%s�2.˃7���<_j�w&�KL���uT��N�r����f�M_Y�[�����Xs�[�7H�*6B��P�ܖb�bV�*�aJ�l�h���*�f�ͫ%�*&�6�hmb������"��;
-AYo{�+/x;���ͤ��cf�V�tO] ߭*S\�.�T�2�BB/��s%M�r�G���5���$S�ǡb���O��Ok�[��,5�Z���Y��2U���m�e�ہ�] u�r�W���\��mo$ZwwCT�X��� ��z�ɚ�k]�-��.g<�\EC�	,�=�3���T��:R���h������/��=n��k휞Ig^��	ܛ��.��P��g���N7�CNa�E�Kv�a쐡|�+�,Kk�N�,������㴷��]�9;I�d݋ʗ�%vD�,3:�45�U��Q����Ph�y.���q +&V��=�g�t�WS���5G[����l��v6�w]V̕c�c��DK恩He7Ua�@:�8��'2�Z�u�w�C��H�D�KL�V]�=ѻ/����g�}튪ɹ�������jF�H��v�0��	�2��hŖ��j��JK=�c+/X�Ӵ��{�Ve���n��Veb5{n���o��]��A�/�9a�J�7�zۮ7�e�����Ym�ժ#�űqk��+1ہ>7�u�[�ާWeG���n@��Mj���̵�������6�G,nV�!��4��b�̛���Rɫ���u#�K6r��X�ϵ�Q�So&����̛9S��˶�zڮ�z�v?7��)��X�Dn��%�w� �G�ȡ[�ݼv����M�(��7���\yq�26t��ջ��뒵D��C�ON��t�pf���B��1��o/�*����m��l�n�y�(=;[�-/�\�돆�����U�{l]�}Q&��%���AQ�;R���YƯNX�su]��fU��4Gn��tr:�v�ɬ$��r��+���9�"�='J+�ӕ��dD,�T�2v�Q):G�sm�d��f[Z�lj��(�Y��7xl��GW��!�w+�~��@����0)��aw�_P~�.ꊮ��c9�
ֵm�T޼��X��;��ݑ\�q�����:���"�>JH�8�fH�I%t�K�����o�����:���\�"q���S��{�wo$D�����q�;�BI1ӷ��__]��:q�qǷq�8���������I$!)�$��[N�{�n�d�vq9w�u��2���X1��x��Ƿ���n8�;q�q��k�;}zv����]��v���,��(�Rr��JGG*3>�NO�Nr>�����PI_�܃�nH�:��S�$�壢Gp��}�{^��'I!�|ߛ�s����� ����ۢ�~>��ﵢ�����?5nQ�^ۈ�|Û����w>֑������[����'G��۞��V�8��N�9%�:)�a�s�K_n�y���^G�f�>���Zů����u��ZNZ�Y�k�dS��܉��R�@��֜)=�t��h�A'��I ���V���/��#(�"�=���a&g�b'h�B
QJ"zFl2��}u}4�|[�����5�`M���\n<�utF��i��Y�u��[P��r��%�ǆ*�����;���!(�>D��BBbj@�,���2d���@�	3�!d��ed)0�(��m�1��lD["L-��Z��}�>Z_=�}����}�Ik��SG�S�8��c�@(��B*X-�������w��*��;t�4F����͢x��v�����St�L�ܘ�D�_������P�8�msƲ�%xϩDk"�u��Hwm�"�b��j�S�,'��3D<y��ɀ������1fFnBN;�~�aD��:L�;�)�X�{���|���v��k��B�ø���:`�5���Lګ$��^A���������Ż�ܝȣ����~D閫�a?/�5Y_����X����D�OB�ӛ�l�T��z�oj) M���5��>��}�]<�7�z���^�z^�e�I��O8�t�38��L������ȾF-��n =(�_Z��C���tSE(�qW�� ��W(5$d4��V/;O���y~`%޽`�|f���C�%��{���?[����ۛ�T$�ם'�j<%�y#X�@�c����3���S���;��d��=��̐�6b�?���; |`���=4��[�zѡS��儶^�f�JU:�˿�v��^��?�����}<��}D�L^��l���/�sil&%��JsqU<�P3Z�g3z�WC�};��=��T�e�{�@@�_/�B5���������Ψf�߃3o�u���	�͘�0&�v��=r%]��ݍI՗թ7��6�$m��}��qUG�w,��4����-F@�*Y{ˋx����^ڣur�^ag�&ѵ�A;1���N]U*�[bX:�pʽ��2]K��.w���������<����{�x4������7�*��D;	�_��Rz�Dׅ9�/~w�xa n@A8��?p �~B�+`XC��6�9o6� 4��ʞ/~&)�u��iZ^F���W=p�����jތ[����ۻ�|=�.-�	Iz A����2�}"Mz��
�ؽH��ۜ/`% :��	���q��]����j]*���<X�����K�sBL��.(�<�,�ss*�u�$��xl�Q��Z�\��Ւ=���p����5�����?�4yR�D�N���������M��������������C��X��.%��ۺ��"|����@��n0��`�@�[C���sg�/k�=�����4���`=@{Mi=���P+��	{��o���uk�2'��R�$�U��e���������O@�^�1�DSqL��4;�@�����|s�Y�b 0xy���X���,Մ*Zo>�BBn�����?r�?1~!�&]y�p�i�ަ�:�m����6�v-���x�pQ`s��\e��>�Ƕ�|hpu���	z�W>P�k�zޟY���]����4~S�o���k1����jn�5hZ�2�2�%�XMQ��HfeE��6;n�M3Շ�1�k�}�"U~�3O/�f&�̚��JU2�P�O=ۈ�}P5>��
U�+h^m�J�<4�-��I�l���o:�\�g}���>�C�X��+�:t������a��i���ݥ��N��!�|���_���APQy��Y��{������u��8ɲ�������=�h*�d|�Mm���e�2�#�5�[����M@WݦGL:]q���]�>2ç��^������Y�W�8��|E����z����ҰTd���YJ2��;��qؖA�Ai�1%�ɔ�	�BJ�؍�ǭ�F4'�o��g��ɔ��9ҪC����k�Z�=�;h����CZ�L�齎[�,�������~�gYg�us
��_8���!=�_F����̅z��਋a�1^��˜1���]0�0����d��sx�[�S��{�M
�]�{����ǜO�!X_�s�����zo��z�T���!a�WS�`�Z��%��^�"���Zg����i�Z� ����B�p�>ZD<T&9���q�%Q���[�]y���3V��FdHgj��!��8��n0����t~"0�>�u���^�ˁ7p�E����1����&1���^J�-�� @5R2�E���97��鳋����3V��Bח�6��)�Iu�h�+�0r�\���9��[~�K��
u-�kX؎���{A�#K��o�c�*l�<�l�a��K*VDk�8Mf�-�DI�c<����wI)��7��F�S�vM�ޗ�ƦECa�-jx���8�wed��}������|t �:EA9ι�����^||mg��xb��;�mx��dϧ^��c���V
=H�Z9�o����n��733q�!�]��Bc����`��	<{����=���by}>?g�-�W���6{f�y�ր��\����ԇ����=�A��#�q>�3e᱒��}6�ǥ�v %��ϚA�q4�p��4f�?V�=lѷ����6�S��� K<y�4���ɒxi��r}w]>cvK
�Ʃ*���j�#�L
�K��^����p!��B�.,��|�v����|��G~���%1MЫj/Gv�$�,�k�M�LF�>��'Ʀu�"����[vP������\��WLn<J[ǥM�p��XL�#���Z�B��Q)�$g��z�o�^z��	���d�<���;ˬ�΍����6��"/���=�给��Y1,�ߊ��P�����l��qo��_Wg��A�R�/�.�0X@^�1�΢@z|�ܞ����Yp	*MmS�1��n��~��y��*[\:�x�D>�<�İS�=~�ԥ' �PX������c/iմ5+��z��t��4#b#���ܴ�y/P��ݪ��应�n��M���w w0���B��H��dB���:eG�=WZ��Z�<�<��GkPe�WB7Bu	��T�?����3W;��r�� ��S�X��P+�:t��o���ާ���H��S���A]]��nU�4�.*nk"�>�x"��հMZc���~^w��c����?��hG�6[^/�u�]��!�����.U����m�^��,d\0j�,�<�L$��-��k�#�O�|}0��e�sMa9��KN�Cٌ�=smǲD�Os����Q~(%�6�8[jiߚXa��:X:�O�;bS��9y�y�ƹ���~B`K�\�~t�z�Ϡ�H�طp/�8�h�c��ץ��ͽ�({��<;��lFGޠ��z�'ߏRgNe�����q\�~�~�����龢_���A��;n:�3L��D{X{;J
6F�`$E�1�{�f��>ܔ�ì�=�D�a}�]���n�a����o����=�<����i�.���(O��
߮`&J�Hf�7e�:�>w/7dé���s܇��y׬�w��RG���OC�ʀ�e~�K��0[����m9���Yu�r��,�=���^��^���*<����׹��\�g	oHA�z�g6GE��"�]kk�_f�n�HC���7�����?�^�ME\��䌆�ٶM��[:y�t��k�ӷ20Fg�F񷖷3?y���o��T]Dw��;ʸ���;���s���������|riI-E���2��4�������B�7cs���7n�X䮺��3`ڮ��<p��J�Q��\W���"�]���N4U>�9�6x���z��'^}"���t5�:P@ˌ��[�x�q�C�8v�����V�SO<�c^t ��Cy���c=_�x���~���l�#�O�o���'�}D�����_�S@8��g��,v�zx2�<z+FD�����_8���ww������m���� (��g��&a,��ǃ>Ba'�pD
�M���3��=0LĽ�B�W�zK�}M� ����:@��L,8މ�{d�$����:�.9����U0��*X=Kc/{��)�,�Pm�):Dȿp}3��ZdA��x`������v��oh��(νCżp�qk�f�O'�g��en��i[0�h��>X��w��ۦ��"j��]����b�3�`�X��r�lȞ���tvH�X�B/�(,u)v��a���&ُMZR{yL7��ٗ�0r�"#�[SԼ�T$�#������@���U�����8Om�ԏa��C����SӸ�p���@B��C�ǨG�����>���I�Z�����ָLL
ݔ�W����V���S� _�+OJ�!x�00��U�pT���x8���ϯ���=��n^RBѢ��mmV��ô����=/.�e=O#hZ���x5�*���WQU�۷��Luyd�vfnN����B�ĭ����A�Ż�1�ٵE���8YǓ��F��5����6���zwG��[3�7�݂����1��k�:t�*f{�9������<��<�C��'�ρ49�����`*M����B��W�yk�o�^�G�ꥵQ�Cř����{I�(�J�&�=`@:"��`�k˼ ��]X����,���P�uݢ\�QQl��a��)�Fd����ǡ؀t@�5צ�	c�����LC{�F�_N��`̼�bOx`y�~5ߕEV�ի,]�� ���~\K���F��2�pk\��;ۧ��C�r�,��t��V#Y��r��DU��.#��"�#�^ם2��FЦ�/c'&�Vq�0�nW�q��G��� �����dj�׭�O�������G:kd��`o�'a� ����x�#V	�Z4)=�G+���.�)��0R����f��o��~�K#�]#R�V�+;�r,=a�=≮Am&%>x�UM���%B�6s��_�
�l�w�1���hz�f��S:�x�w���^��	zos
�ק��T��p!�9]�%)��
{���j\��TĹ���]E��-ƻ�xs(}Ǡ,�]繽 QtÔ�.��)�-���.694e����ˇ������=�qs�20��xJ�r�Zzp�bH�%w!eV�Q�ƫ���Y������oֽ�*9�*K�����ʖ�_j�W�q=j]���%^Ӥu/Zqfa[\΋�b��o��<��u�ܝogҀ�>1ۤ���x =�OW�TY+��k�|�]��P�d6Ä۾��	5}I�ð�K�1i������b�+/[+�8�^��|C�>5������?��̅����������Goy+�ۭ���T<t�Q]��z��2��� L������4��3�n9��H�s����;��M5G�=��[��G��7=��z<�k��y�U%T5Sᕱl6}�3�K���RNF��z2x���$=������·�(��ޑ�� j|^ī�Γ��.�;=�Tl	�ϒ�U�ݽTG���tDV�ͅ�]����3^\~&#G<{H,MR/�N��F��1ߍ~�ٞf�g��{�TP�Qg��xw�hr�7'�5�)��/�����׻� 8V��/D�][�k�r�p��-����/�\(�����b����z*���6����}�j��ޯs��l��yqV��ù�y�B���ˊ���/��-$(�SY��/3�0�'���m�+Vo���wzB��PJo|�0�yk�ދ��{g]]���[@.B�y8[�{UU�l����uI�pn����m�����U�*C[���L��^���6���gn�c��b�u*�Fj��D[�&G�q�����a���	��8Gc:+so�mAL別��}�1G���s]�=�u�sW���O�vǧH#]1ӡ�ʏV�Ж�1�X�5�ݻ}�u,z�!�N�RD�&)[��`��c#�y��	�s�DBj�҃&�Y���VU�įG/���Z�3�8=�����������l<0�r��<��znT�P��q@�����#4��+�~���
���YR=�z3���x��G8�r�� h�['^�@	�v/=���V��U��jI%?чƽ_�~ϕ	�EÞq���͂�	���
}`�rz�0+ĜV'9|�tU�Ysvwg8���[�5Ȯ��&ȸ_C�y�l[/3�b�~�Cg\.�[�JQ*�]��$�����G0^��Z~Y�Pq��������g�~�$��x���=�C���/-�c//��F%yڮ�c�Y�פı�{Լ���[����	����]�1�pރ�5��X�q%�y�"�q��rz�*��怘��S��ݮc��	�>P,FW���Z�\��������1�+����Z�t��FhX?�A�� pr�a�:/����"��Ö������������8�$�4���wV�/_�!ݱl0c�4�1gml/ޗd��ˑ� ܔ�u���j`�u��
K��a���:3lp);bYkv��B��������0u��'5%Z�l/�u��d�ә�qV��~� UӁή����5º�Yo)�W~߼�s��ߺ�1��kk+-���r�5Hr��I�O�$�7�DM��R�'���ǷJ�]:k�@ ��[�Vs�C7�iO����#\g4G3���
ߡ�d�[�g^K"����}����΋��	�o���`j��{g�I�e��)��(>��RV㑶5��y�\f�3:vxz@Ǯ�ծ"��)w��P$2,W� m
�ُ`s�8ht�g	-8�X���m-mY���m��t^-�QL'���1b
�A�0@��dޟP�ΞѺ�j;WRk3kUO�C�.h|בv��쐍��r~Om�:OV,��[;z£8�]�/9�Q*z��v�2�p�LT>P��hLoK
~^�_?����R�@~?�8
OUQB����<'�N���Ǯ-���y�v��
��I��_�M�&晙.L<ʜ)��x�i�s��H������a�vFڢ��/L!x����8v4�l���ى����u��^����|~�I�0a�E'I�K��|��{��3 @@�0Wk�����suj���U�-�!��cN�;jJp-(�E�c���A�?t�T�� ��<."����-��֥���Ljn**<�������UF�רY�9G[���R�vim�ELȐ�cz
���24m�
]�'��w]j����g��q��Ƭu�ȸ�u���V��m���%N���mqm���ٕ$���k+���w)]q��T�^�Ox��IB��1��Ae�gG��j/޷Ho��R�����|�s���S�����Z�=�mg[[]|�m֣�����mf�ѵ;��(��r-_sF���t:�u�a1k��l=`��F��4:m��X��z7�����αT�B��D���u�9�٥n6�!���Y�x�`��Fv��ݲ�sS{Z�tPNо(�V�*8�ʺ5l�䁙�j�d�u���u����7ae!��e���ݳ�u�\�n�p�(�J�J�h��Ϊ�;ѯmV���ouB�����8��j�S���-�c�����]!u֭u�9}\��e���^G�X��oW;�3	��P�.�.�^�����;sLٲm1%�=��lk�s���&7D�gFYsi��Urt�:�e%��3������Z��M���"���뫳�HDwTA�}�0�0aկV�8�em�/VZ<2st�����O���+�ۣn������]���I�j�~���ct�a����]����	��$�{FYl˲�N�H*)UnZ�%%�鼬Ԝ�JzʖԙE�"�4r�vUr,LSً�A��X��j�mn�U]*�u�����X�67�>�`L�Z�0V��(��j�P�d�}	�X�L�"���L���e#��	��v���75��UO�oNz�:��^$މܸm�R7OC�&�j�;��6������dp����\���%��q���"�:*���=��p(�ak�;e+ڶ���ٗ��KYA���un99���2I1�5\e!In-��$`۳w"���&��WL�«n��YJr���#ƛ�Tv��-�]��tz�'۝���q�5s۹'Vk��\��N˛t�mµ�Y��0v�G��p������)����������e��w�_[V�l�qd#j��̷�R9��&�-3o�m����w&�F����V��ASm�:��������^�Wb�g��RF��Y�xN7E��:p����\���X��v��io��pq�K.���8$C\�$2�sRQEtr�E'>7UaT��4��zv��w�\�Ę��W1���K�v����R��/E���(ݮn]خz�{4��]a6���[�ˋ�w0g�^��\���B����`����O��4�F�����*�Tf�S��kyE'���s�QRG����$���!�[}��yX��Q$�~ �C��+$)��Շ���P�f�Yӽ��<}q�ێ8��q�zq�t�ק�o��>I$!�XZ����U�Y�H�s��''_ݹK�� ��;w�}ߝ����N8�;q�q��qӎݾ�;}t��B��@�D�!$$��=������{���I��8Y��� t�tp�5��kDN���1���p'pq�I����8�t�D!C�q�rp�s�ND�8�G�H{n���H��Z]���c�����r�v�@�}��(�tI<�X�t�@��+���?6���ޭ�T��"��Y�����q�QD�:�'��qr��k�A$��d�~�H;��."Aƚ?�):/�v�؊Bq��Rtw$q_�Z���"�vQ:��q��Ҝ�D\A�@?n��^<����]?	e���;�=t�3a�d�dS
A�pJ`���vw�Y��x�*D�d�R	�Uj�*'���:t�B(�_9�>|���Y�.&dL��f�p��)�]77��	���&C�O<�ʄ_�Pb���S���\��
�r�N�5��p�����"m�/%�*@P4vJqv��1aK:y����k�*�9��a7�X�R�xB���1*��A_~$==^!q|��Clȥ^~�.5O�X�;4ۻ[[ݛ��w]{r{e5�����s�:��+������k�D���%�&���4��ְ�\{k��?Mk�0'k���<���3���y��h04B`cnL�; �DT�ͮ��9�hL ͥ�vk�m��^�0�u���	<"���ŕ�j�5R��A�}�� <:�}�����
�^�d|�U�!Eg�}��v�ϻ���0iL����k�%��wc4d�ii���޾7�ؖ��P��I�w�	�o��������M�\��r{��=�n�g_Wwn��h��Jkx�������5|�N��>>���D]��.#�}!��)ݱj�1��z���'M�8��O�%����|�^��"q�_��觟g�����4��ߧ�)��#�?τ�u^�f�Ms!v)KS>=w�{�:h��]"�����g���3G�s�O�S}�5�v�*Y�N0H��||��w3w����z&��ð�hé��v��p�����į�dwV�˪ǯ`��u�����;/^�a�8�:t�H ��<�޳�m������_���eV�
Or��,~�b�Ui�J�/��B��w�2~:�cC./�������E�� Ժ5�ϼ%0	�Nl%%�j��}���p-���+J�b�}�<N}M��&��`��ʟ9�>{|�"�5�ާ/��;�Ru��K"�@�uaJ���~z��U��YՊ���{��3�E�!�)Q�1�C"c<�Fvz����/�,i�E�7E2�dy4Y})Q��=x/[؇[�?0>6��CoSG��t�0���S��y�ߩ�e�sɕ9���z�C�k���;�F���^݄Ɨ/SC�̘C_l��d�!�	��"�~a��x��/�n�tf���y��ؼ#NK������ܫ���ƽ�i>�����#��?���,�ђ����źt��_lo.l�*�1�F�݅�ekߒ��-m�k��*FVŰ��#�7�gA��_j���e:�k~i���EtMϪF�<j|&=��c����X�Pxn_St�[=�����\4́��N�|l/_eո��^~�sR��BA	����
�~T�_�<�ٙ��AM����*�7��Vr���VK�e�]���a]��O\�l�LV�s*�~g^�����ZU:�̼�Z�N�Ӱ���b��n�p)�m�p��t��3�����GE�]˽�,�����ii9���VǓ7y�;�^�:��k��>�8�H	y�y�  ���;R�uW��\9�z�I�Z��5l��la{~�ۺ�e^wLYТ�K�>����:R\E����Se�K�%Y!��[xCN��������|�WW?5Vu;I����?�*k���!O��/��0��L��h�!y�##r���ɖmN�ogwe��e0��H#Ls��z�>�)r��#^Y�9hjC��<���}���Csl[ؽWP�������צ-q��
�`�.���l�z���x]]�`ql��@����̬\ڶo�3�v\]���lU]{yMWЃ&6�	OI������o�������W��bf0�GP�fl@���W��y�nU����2�I�W)W�M��{�dd�b��������Y_()ZNc�_/�H2���́�j�u�y�&I��a������yS��"��J�޾�@��&�[\vI�p-�������}<#\�S����� ���q�b��������u�|�b��E*J�xsP+�u=���x�����������7K/�
�E��j�z���t��i���4枓�yP9�iy^=4�=� ��5��t����<��V2��e����)��-�so�'�2Q�����V��M�K��e�����X�|͢G7JnA�v�A%g�ԡ�|�����~}o��k�w1A����g�4g�����A�lEdc�W7��(;$��D����W{�x ?����P#�Mt(�"�u�=�=�5b�.>�����{�*�%s�x��_�x�x����=|g`H]�M�0Чj�-��M�)��wd�#\�T�E7W�wQk�M��8��<\
��}5R1��WGuyvTn2���پ����� ��Pna>A�8��x�;6g�ȭL-�y��<k-{'�z��q+C�:V�k�+�gW���קPs�O{ֈ8/��4?W�(1l�}"�ۓ�㮮��@�E�ƨ���ٱ�X�"��\���8���H:��h\Q�0�M�k��>?}4h!���W��:�mx���%9.�X�faM_�k�i��ұ�A�0[���5����{no�zqX��׮��_����Sᕺޔ��*<�^<���Ҟ��6�hl�k��b_,�y��]{�$9{D[~�N4'���S�D�%�^�-@��#�z�m��Va%�;�:w��r�=;����=�������#T$�n��ը�M���#�z������gW�|����4+�r��@��|��aϐ���3����XN-�,����T��3�)y��R���Y��#�s���Ŏ<je��8Q��k�hkD�5�G�Q���y����E<�U�n�F�վ�-���5o޸껨3KZ��Լ�wq�ǻ�ise����J���[ь���U�6��p�[���6������?O/?�:t�H��*]y�3;�=��o��5�_�g�/g��7������f���T�~[��|.'�q�+_l�kU_njǍ]���������&��F��R������l�L׺q��t�P�i���!E��a���b1lCM�=�i2��b��n�I�$M
�|��v��s t��v��خ��V�?f����ף�8@��n!��x�Ϸ.y=�b�'X�y��i����,��z����^�dnI���vln)�/�!�=K�����}I�P��-^9r��PX���d__�����=|;1;	��p��5�k� �`1�Dn/S��O�$�2I�`�E���fCo���y�y�U�R;�-0�m�#�$�
���!�~_�#~��@fl7B��z�#��7 �/k23V�q8�k���2���˞��z g�����9�f�p�hsS��̽�r��*�V^
�M���׽p�y��߇�����	��4��Z|^�9���A��{R��H[)�ڕ��ݼ	`��^��2ב`;5Ƕ�&�^��h;	�:"�^��^%���ζ�y2nf��q��n+z�}}d��r�&��F��Ֆة�f*��3�9K�Q���Gh�.����hYյ���y�uVˬ��.����;@�������oq�W��6r��n/�L�ns�-��s�9�ɿ��������5Ҡ%����Z�1�p�[��C�wh�訶F�Y���>d��r�CO.٪�jY��&t��<�2�)ᮀ���T��	=	z�����s�X侘���<�3k���܇zk�7o�]1p�5B��>!�� ������(�T=���Qx���5��A�Y�]d���[Q��<�Y�b˱��`h>Qmu�#��n�/Z���6fǗ�p��g�&M���O܍�1��=��[I��y��ޠ��;�˼�֢S��W�i�S�O�Ib^���P��w9��L���s�R�����Ş\�G:/�&���t�*x����ꔝ��9��W�T�h0��ټ�e��#�>���]��A9��� ��=�{���EL-�R.�st����Uʚ�z��7ʋ�f���c��p���Mn�ϲ�6ﳤKxׯ�;�xB)F�;�n�������Zt��%��P�Ʉ1���L63׸F�x.�A��V�������`��|l7�b1�4��F�e�_�o��JPۭ��xe�0Ҝc|��fV��{�ؿX�����'j�9>{���o�;6E�ꈖ�B�r������LS��`'qL�|�~k�sY�s\�wy�����Jt鮄| ���菼k��G����f5��j�썫\��H:T��'9�݃Y�f�5�+�UzdkJ�C�}l�E1ק~�^R�/լӰn�uG&b���1�We^��P���BdK����?y($�{W��&�F�Ű��Z��[��Ղ��nn��=��;s�H�f�y�*�T6��x��Lz1����#,_6�IQ\�5%i~�a����p����ӟ�z#� �	����P~$ɿ��mV��}�/{�����ԥ^���X?PHަ��0/�!��^��|d�+�/�CJ�
$.bوǽ����٧yՑ��N�_E���P����0�-(dv�I��Qr�c�LĦ�b��u�gR�}B;c�q�����ŗ�`�o-���A
|֧���c7�m��}6r�y������.�R0�h`�[��±xa�*o|�5�%��3�b�����I~׵�w9�ҵ_Wf��������K��?(��O�������G�)���A�ZxN�E� �>d-�Ӱ�>e��Oa��%^<^.́qq�,*�@�y +�:��	�d]#�zXomȞǨbX�K8���6��z!��jL����Iw50�G��ݝ��9��=������}b6q����V��� ���ݣp��봮.��B!���3:�����A{����|9����{f�4���񉓾;皙|��u������] �N��A�3x\fow%]�=n��?����_
�Ak~c�'���x��4O^ïA�&I�����Z!�b6#��G-/��cIG�&�~���r�}��ŵJD��)�X-jQm�>+Y�Y��v�D�D�DJyp�U�'�:��Xn��Z���32Oi��<���`��&ةxZW8�X��w7�olr��\9u[>5[��ߪ,�N؂���nx���a=����T-���S�=̕�uo{��gi��ĽI�m�^�]�����]'�k:�e��ýgW0YZ�����D}��ڑ��t�j����z}����'gO'�W>N��l�:����}�4�b�1�F�A���":aغ/��fE*�0�g�X�RړDS��uW�w��mD[$�o���ca�8��r|�_Y'�.��>�#=��}5Sgj�1�J��W��;�X/" &w��\��W�+	52�.(�� �M���:���C���ؾ���:��I�=���^�0�X�f�ou��=����vD�ǂ"�p��^~�^~��W���e[�K\]a���SՍ�l)H��a�v���Z8Xͳ�}�y� �r0�*��}8X�Y�Z��Q��Wً�l�a������{:¤�&�d�8a�V��m)��bN1��+{���om�ac�*��K��{��O�8�k�#�Mt�����<$��g��q��r��EF��Me��.�E�E��@A���i�}kO��e�7w6��:�N��̂g�#@{�lOsq�oO��ԡ���qW(5$d1�����Ri����LO�H�~yON� Xb��=����)�T$��μ���~����ej�<�p���~檿\�2㦾�`������$9�Y����iֶ���R
�q�(��Y��G[��;o/�[���νx})���B�),�'?vo�Nu�jR��������'��2�����>���N�u܅�L�sPuĻ��F������6q���BΜ�C�5E>�l>�RÝ�o{�˅�*t���n�
S�qM�^fOA"k�����I��;��;�'ic �{�Ʋ�9�5遣�m�2�V�z�n��{��|���!5.ב��ƳE���l������J�g���	H�8�z���.��̉��L'���]B煼)>�R�uogV)l^Y��$�L8�}���h�����m�%�:�2:Gd�q�}����U���Y��cc/�f�C7ص�qWz�{�z+�s�On��~�1i�%LbM�a�\�������:�=�EC��������| OԺ���'����Yy7O$p��.�e@�us��y �r�ID��x��r]�8�HUeU���u5�� }�]5Єt鮄RD���I,�}�����)�_��XI{mn�*j��W��2�E>vz�~Xi��t��i���'����{}�:�8�ҵ�%���Q���j���|�~ ����-�s^{�e}/�.�N_�޺���ݙ��e���c��{����hsH���Hg7��r�v�w
�[�Ň��zЅ�l!�.��Ľ�5�٢ù���f:�L:3�l^\�ᥡ���NZ��<��à˼ ��D_�~YhT"��`�	
��Sr�]��?t`�,�-1�oE��`�i׊xeC 3:
�e��	=�Ƕ��]فL5Y�b�;��}o�s������]; �	�M�ۦ���}hg�b9�<�
�ɢ����E@��3��ev!m�)��z46+öa���^��&� �s[��b����H�o׋*��:9	.���������Ǘ�3*�
O~���(�ǏP��xjkgb���dC��s�+1����Ny�8���x��Z�Y��-���JK�	*q�����`����d6�£$[c[`��z��7��<��4.j�o��*��u��b(8�.�*��v�H���̧m;��?'�3o#�4WX9*sO6\(�&��*omfEą���[هp��R���)jER�+BZ��q��UJӍ\b�>�I�3�t�R�ׯ,w�@u�m�j|�b�W�0O�)�r)�p�|x+y44W�"�Y�Qf��f�<hn�.�|�P7���yw�]D[��uKk����Nq�b�V�+�%ڡǼ��x;y>�B�{l�_c��4e��f��t31�b&6U��n,ziG]�� ١Y�X�RAm
�|Қw�I�V̈���#d�GZ�w�l)����1c�X]�}��GvQѕ�V��Ʒ$�N�J�n���܌m�՝բ�l�	do��jU8�h�����TMi�=�O=I��׽`�ՂH]Eޯ�+�%WUԊ��(C��T��4N��W��b���5�e��Y�\�ndiU�.����Ku��gp\ڧ��G�l�^�]<7�7����|5�k=2
�W�?�;�]�*j�[�6x6&ׯ+Y�LU�(K�WUqD��9�u.}����Pݒ�u��g.�5��4�U]�MQ=���B���y�ۺ+39��T�k3��y��#2f���zs���e�"���T7I\�e�)+���-G��+��*��j���A��+������;x��f�hVL�j�]b��'�^�K�#�����i�I�ŉ�OD�xk:�:�/����Ǔ1͋�w�����:��hw�4V���J\v��g�_l���ɺ[t�ف<y�R�[��r���fQ�*Ă\��q�.LǪ���go6֎i������ꤗ��99�#ÎPk��y7�%y�X�0����Ղ��������;�Qb�;kp�nu��z�7�Whe�S`;�7H��\L���a�V�h����[w����*���i��|���4���8[�Uꪫ�,6�rdY����j��e��il^bǛ�"��}�L�.��ؚ�kB�US��h�̧X��&4�Nzz�:�(aS*�q��n(�f}�
�p�A�����5�7
��Ʃ�N�Yj&4-Z:�k9��."x�p��:M�N�	��W1ҧ���ont�Nʀ�l���ý��*�kt�R�,��X� j��%�������HR�n��J�Wz9bv�Lj��/W˜�[MͻUw٘�(�[�ŕ
��{�9��5��Z�͋]k�8��8j��
}������UJ�HΦ5k�t�ǋl�TZ�[��7�N�¦�T�8��¬e3h�ή��nt��"5a��Gg4֨e�q�ɽ��_1}K��p]Xr���i�{��F�Ŭ�y�H��H�I&A��ʫ����;���i�dGG�e��ۻ}���C��	׷bBI!P�D�=;z{|q�N8�8��8��q�nݻ~��Z��Ȉ RRw�g���_���f�t\t��\��w���׏���q�q��qێ8�ݻv���׏����Bda$�X�5�)����B�z�:���,H$�����N����_�E�� ���d����J{h_�8���䟚��U8������)����bs�3�T�{Z���~,�AOv����B۵�s��3�!���)H �ۛv�E/��		%�rNQ,ߍ#�$�L�f�dy�?7X��Nq)��7��:
N������W�G�噠�_��D�ZĒf�QIȤ��I�:Nq��qC�����$���"9#�+˴��tTH��?��ｈo�爗T��aM@�����L�C<�-2D���	�|LD�|�(8v��˞���1�Ǉ��X�41�6����\e��q�U\幅#��k�WT�pj�ouC��(�uD���f�h2��Jy���A��d ф�D�k͒}$��l6�mI (��|"�b	��
 �m�R.@�RH�P��1�<�%��#��R�� ՉiK�I,5�Y� ��鮔�#�?���{��s�d�ztld��}rϒ��������z��}�sI��{C!�ۇ~�����Jaz��Tc����3��I� �%�u�,�^��"�%����*���R��� ���ʒ�ϡ���L�a�0�O��3}%�}�]0�h�9O-,��4r�{::	ǵ���Gp9j}� Pw��.<�<��`&�m	αE����cv�1gw{kǡ����.�z?7%�.��@'ݮm��`鱧��5�;t°��*���w���o�a
�LU��]�F^�F��}C�W��8��E*q��ZGU��
��uNʺ�9��k�I�1,�@�K��7k�gX�?s�:�W����dgX��Sq"i��GS好�CHd9J�.3��r��
?�=��������z��ƣ���n	2#1e=%���]�X���vŰ��E�=���K�	�}o���mv�żW����97���g8��uo?7k$?��O���M~�~��kü���qq*l���%Y!�	A��׬�U��}�u�2�s��x�v��-�;P�C"Y����vL��B�iNɛ���wfDc��V���ۗ8:�?v�d#��^���{����;��6M�GM�ǫJ5m{���/��4���Dz۾�|xsp�������Y���n{{2��]Æ˔���c���)ɗG��x{��7�5����K�צ���] H#w�Y�y�+]�9G9��g��m݄���28�%P}K���}����Q���=<B��U٭��4i?E�0���R2�eEM�MA#��ѽO�}o�a��'���՝�����d���C�.��4dzdŰ]B�ڈ��cKJ�����Fq��L�^�3�os:�t-��9�[�!�.�D����V@S�ZͮApK�.|���U&:�v�m��{
����C��񹩜�SۼH0!<Ba0��q����)S�e���ί��6ӧ1)�M�˒UOmo����uC�������#\'��'5N_*�/�sN����<L�x�a�nq�'ܯ�'b�A�E$����cz/�獋a(�Fʦ��K=�}���w{�AK0C)�dzC���i܎j�L��`e#�Fr����L'��;��.K�����8�8"�3���۵�xl�^�]��$&2���X�n��.�g�k�W�ݟS�|)�ga i����A/BZ\BgT$W�un�5���ׯyU��N%��yW��,�fYՏ��w6lx�4��ڪ��lݺ�OZ�8��jՍcR'�v$'�x���UK5*Y;��@����i���}k�R������%,y���t:r�=�k�SrwV��� �	=%$�-)J��p.������~�?5�tȐ�B'|癘{�����kj��,�５����i�½���&��}������
�C��6��'{:p��a���g{9�t0����g[�i��$w>'���F�ܾ��?,�I��!�AJ�k/x��b�J.��4¼��t��-�友�a�@׆}��^��)j�f�'3*����Y�`C�nۀ��õ�$��{�O�z�_�-�@:f�}�%ߧ(4_H��Ϋ�+'������x~.�-EΌ��h̺���%�p�h��HI�sd<DT,V�������W�{��MN���(��P�DZ�g���H)�@���~[�W���"��I�mz&���g_uu�ӑLW@�~y�w�(��<�{������6�8�/���*�rZ�w�AH�~�^�?Q��{��W@��0�\3g�P.lD�<s�Ol���6r|Y�3avs�Ɔ�{=�ѿP�ޥE�5gd�T?�{��0�)��ހ�Ƚ8����{/������ݣ��s� V�=�}k̋ۘ��ZF��GԝžŰ��к1��5���m��(x�5�
�<�\�y�k���"W.O�A�"�!i|^�"�Sv�Uɘ�坭�6^`0�����i�J�Nv#]#����(&��M��ˡ����*u���۹j�vL(�GHĚH8Ɇ�s�7���r7�?{�������� ����&aۗgScaq��A��M�i��u
�i2��1W����&�x�8_���=N'U'=���,���L�wխKމ����0vX/�;OeI/d�2.�8Lq�b�uN����_��9���:��?a!�3��~��E��G~ ·�K4�;]��Jk_g4�3{y�c�����Jxw3�����`�DW�&�{���U9#��Ηژ���&qvv�8��.�ΞeJ�a���0r�^s ��(v������������Գ�!�uM�ڭ���-��Q�2K���t���*�����{w�pÃ��a�Q� �w��o��9��2�JD^=z����sf�T:��ֹ.#7����H/A��צ����N��/Q�@��xe��$_�/��8E���d����;�K�0�עg�3#���1�����̄{^����l���.����f�O�F�VE �=0��6��K.�`�mg��S�?�~�o\�e�+���'D[O��ײ3�`Je�Ӥ�/V�k�[�^�����J���>��>Ǩ�u�}�s��j�^s�o�A���՜ʢ/N�$�$�p���U(��o�kNI��SǙϱ���"BȂ�w�=]0#���L����;�1[`��#bP�6���U��V�n]���y�oz�^�k��N��$�$%��ך�ݽ��x��&-X��.����umԊRW���wQᙒH��*?ۏ�.���w�<jy�_����P�,>"t�L]�.�O�"y�]���r�{���ֆȦ�-l�k�A�7@��=�� ��zq��K< cw˝�V(����w���C�-�[�v�z�P��zd���hR{�r��ǡoV}ͷ@����Sn��d�!�Aip���b�!�µN�>׈�ļ'�	I`��%B׽ᗝ��2������;���2�r�\T��5���[C�����+z���.p1�nn�i��T�����[piq��@�d�aO�|����p��`\��cH���WHY��L>��զ��īuL̓����Z<����'\�:j<ʼ(�L�]���
<�6ؘ	��^�vUB�EM��{��������OE�I�=/Dŧ洠��ҡ��k��>h�y�c~
��u���w_v����]��8"q��<c������ZMc32�o�tklח�;���q�bT7M���f�� ����UR����[�\z|�a��%��dK)vy��*�Fń`��uN3ʪFr�NO�_gUj��R��Y��^:b�v�j�&�7���v�T ��@�6�����<y�T:s����"5]�ȹr����޸E��(�;i�ḧ́Gp۹�-�a�0F�N�����.K�[��o*��'��"u�)���9�Y������%�x��:t�DdI^5�"��V��z��>p�5� ����}t�!٪�EtS����<j|�gӯP[���Y�g��ޞE���	����@��l/�}��߾�3ӊ�X[-�m��E�N�G7vG�4�ow@�p���~$nP�?v�G����&��.!�t\LR�O���ğ2YֿE`K����gR��^q-@�rC����k�3�\?����dm<H@���Ah�)GZ�+�]wY�Ӈ��Z˩{��V^O�)H���O�Ei�w/b�׹��q�&C��	��x`��L����[s.���?�>S�G�%B���e^*m�d��}͜N�:,�'\��Zw��3�t����u��cN<������j=���WlŨ�O
�3��<�Z4d(�㦻�zU�@^��v/���W�@A@�.���Pܪ֯>��x����W7��z�8�K�*i��T).�g���?0������>"^����m�6妬����M�˨w7�S�}c���X��JS[\vH�ȸu@ty��	HlI����w^sdds��EWF��=n_l@�Y����'$"4�.�����૟�Z5��^�Qk,�y�v�]^����Vy\Z����M����[�����V�ˤ�3�)DLo})��#pwO�"���9�<���;��������莝54��滼�N]���a}8�$É��4��LU�H�^J�j�g�G�}{0�����*óe4MqsK����&�^����V���s+�E������@�P3�%�.��k�m�ݕ��N�ތ�!�5���G8~��|��/�����5�z�Q���v�/�y��u�������C�H-��Yb��ܣ_�~l=_4�Iՙ8�wO��)p�E�>m���ܖ7�w�sꄑߦu����8!���>�ȇb�z_[$-��_�$��2�3N��,�[α�Dǧ�η��h4v{W��@���?~W�O�����z�u��MnQ�
@�N:�~�aD��:L�o��נ����k�<X�gh���ޚR�[��ÐA�%=Äڻ0�������Q>=�Y"��jWj>H�MKS�ޫ۽��Qm����h�,���p�֜�G�]�P��%��.a��O�9C��D�X���̩���m�+�3/`�ĿB���-z~��y�:/����{�ɖ��g��S��P�%�rZ�M�Cj�u۵�G�ű٪�$��B���������yd�u�kk^�*i�JR�_N2m���?=�ӯZ�Zē���Wغ뛻QY��� T���(5T*Ɩ�;:~��smwr��N�]WIq�̆�!�>��yy�??/0�0fo0��n�E*��\�zd4�ͷW1e|�*J��*����TEo��P�%�̸sM�Eɢڈ���8;�����Xa�����5�J����&�*�k�
ϬD��𥦥���z����vd���@�3' ����&5�F�+�E�5�8�:���TE�w��ok�X���^mf���B��]n87�V�6��������F��B��]���7"��6�k�~�ٍ�y]k+˛�-.���A��k_�={7�U��L��`&(tSR}#�)�8��ٗ:�}��Ю]D0���7 B�S�L9�ϠK+�.���dI�b�Q�T������:���c�1���#���=;�׏;��ړ�e�n�3>f�ԘS����2�O\����;ٽ��<��r��Jԩ��('�p��X���ǼQ�l|w�E?/�����_;
͚�+w��ևl��*,)gO2��"~Vt�ʹ��
�����c�fዝܨ9w���F+iB`s�Q��<\б�(%픿0;Q������7���~eHiC!�q�v�vU�ll��!꥕�s���ONЙ}��X�'�s�����-X�%S�t]����"]�:�r�W2)O�ṉ�X��r�6�IQ�bSSq%.]�T�u.;����.��&��)�;w:�ə:�a��'^S�����:t�P G�f!��s�:?��w�򅉲�G4�G�O�ja��vW8�ǃ&I	-�f�Y|{��'^j�$1(p��j�U����h1M>����̮�b�&�V%C��Mk�&�29��,��`�))���S��O������/�����]q�����ك�Ra^&%=a��ǧ�)���Te����6"�сl�����qCCᬺ���V���c@�E7h�H=���۾���;��P�u}�I&]��D[O�z&�X���f|1���.'ѐ�Խ[�R�5�����Yj<��og8��dD�$ɗP�:8�5��r�r5曍�M]1p���ň�2Np��ЮXC�J;�����R�捨�z6ށ׬�L~�������1��^�;��N�͟��K��W���:�Q� C�Ǟ{nY�n�)��ʗH��Q�Fc���ιv�밲���Z��}ghC�iN%�a�
|C@�S�A�-@�Pp*��4,-v̨�R��۴�}1!�삢����t�Gѐ�A�4'��z�pƽ>�I�Ɍ�J�''��w_Gc���)�%�|E.w�PO�u>ZB��o�0� �CFB�J(>�ј�!�m�8c�S�t��|徳�����6�;*9��V]-V�f۶2>�c/�Vv�s�q����ߚD�W��ڲ,������D��99Ǟ찲��
�d9w�p篰F���
��9R�֣L�Au�ba�]U�cP����q��G`�����ͽ�?��30+7���Z]ع��J+\���Qu��)�- P��O��8nvkd-������c͈�{�w�ox�b�R%U�q=�z^��O�a(,it�~j�k>��F�k��~��	?��� ��xfxE����cH񎼬
�a�"��d�2��5��J�s�qͥ����v�A��+v8���:"1���ϥ��W<Pبzg|�ʣ����+]&��� +���\�G`eb<��ۋ��+�ql6F�`�s�!��ͮ��;6[�<���Ck�5>(��~�}�9tk+wV������=�\�:�����a1�|�Zp�3'��3]�*�?C7�z��ǥݝ�`����^g��6��w��{D��PI�r%��
(��H�<��WY�qZ���7��׻���;	9!��q4�?��^��鮡�=I�F��8���ߔ��-�8j�B�sԽ[�J����e��1��ߴ�4�.�/�w��m��OR=������ξ��U��"�ZF������	�G<��@��J��J�T�����|]����WT�`w��#���`w;��&���Z�D�x�{��D9��q;ׁ����
��Ie��s&t�uwZS����:�Y���1]V���G��f5��,�M��7] �/o"y�4k'=��qv�]��9h;�b��٤²��Q�u��u��6$[����*��ܳ5��+ȇj�u�^WZ�V�H8�u�Z�T�]E��VW$bS��j�>�9R�� ����ф��n�K��a�.��-�̓:�pЏ��"�VP�eZˤlև1�yػGZK3s�]p��y>��]�t�Q6�ܨl9���/��1]4E�̺�]F�TG;�[ًy6�Z����p�O��M2��w���Ÿ���T�9N��Z�hA�g昧���Q��kJ��W4U��c
5pG��[w�%���:�̬n�i;i�[P$4�>�=r�b�[u�l��qr�N,¾�nv0�L=����<e��0@���DS�7��f��f�׌S\��U�El6�ֵ�gY��w�̲g�������\L�V�N�L�h��[☣��=�v�ֻ2gc�������Y�mp퀄�`a�-*�v���In�KMf�X�A�:4��q�z訯{:79��[q����x.����f����@�=�,:ŭ����]n��͐^ʘe�yte��j�9u,��p�Sc�l�L:Qp���b�iۏ�Q<�N��G`�Wm�d�?]'��~�S�Q�ĥ�U5�Z;J�/R ~��*�x�0��{�iye��g�{+��]W��ie���>��>6b�F�O�ђ�6	���x�ed��Qva�e��h���ʚ_H�h��;ڷq��ٴ��(�.�E��2�3�p��6���/�77ݨ8�Q��WTY�u�Yf��dF.�H��Oj6���� ��7M4���bm��
��0�L��X�MwݱC�{�l�{�͙��6�D=�P�xh��QRX�Ϯ��m�QŪ��ds�m��)�n�S*�$�n8-�k�(Fb��WKgV���4����J�Ց8&%%E)C|�����vK�[]f���'D�9NT��7�(�4Ǐ���ê�������u���'a4�٢��[uz�P7�L\���'Scz�y�_c��N�Y���wc��nW��yS��FR]�) �Vi������c���a��RU'>j��]�X���=\�4*em��K�.t�AA���B$i��_^��9XQX�1Q��rޙ������:���}�l�}׵�X���qg>ymgST�����N�$;���\=�l��i
��O{x�*ؕ��eDU���'k9�;Rj��+���e����&R���	�Z������ѽ�'j�������NjGBNi����Q8S���G.93����2[�ܲ�{��aIBŁHJ��#�=]��Qe��\�p�qNߛ�Q�;q�>��q�{q�8�8�۷n�_X��$��$�G�]2r�|םgs���../+D	I�<�T�IedX��������\q�qǷqӎ8�ݻv����;���"HBE�$c�
p�ӯ;��>_:��";�L㓼��y��YOͤ|�ydQ�%n��(

�i�c������+:��J>V\TQ�!'^YHDY�u�Pei׶�̳9�r@��tDS7���y�vO>z\���)I�٭qK��|�8f������D�9p���-:*m�o�ג_�_����9 ��I.��#����˂E����:.�vqG	�%fp�wjTY���m�vr<� Ok! Y��?�TG|Џ��ɡ�ֻ2�$�9'��_Y����{��]ꔦR����m�-��3���aջ��oh�h���U�*T�U�[��7�ouC��U[���~�8���� `���W3�����<�'�?Ai=�`�H�Oܖ/<��j���HJk�`&�jjٺ,�UV�fZ�h���t��X����1�ޫ����ft��a�o��K��
}r�YА�Ğ�Ί��M��ą��K"��FR�T��}k'ѭ��;���qu0����9����ٔ����0 L���]�,��9�Nl%"�PIRkk���싇\�♟Zb�ڡ�L�Z�����a�ʟ!A�	�܃3��$��LU�H�����Η�d<y�n�N����7;���N�2=|#[�c�l��Cy4��.�o̍�,����2��!iy	GKXJ2��^�w=a:��4O���Þ���(�5X�����]��Rrc/1��i�{Pb��(�V)�F���4��(�>�6R ��S_��}^���f/k��rի8�������ٽ�'� 2<�+`��\�����#�?�}a ��y�b�K�c��%1�MW���Qn�;}�7���g��u���_��9m�M���_y`p[���F���Yu����Z;�ݮ�m���j-!u���Cl���Y��N�]U**=f��71C��ї՚�d2����I�T��]����lT7z�<�f܊NZ�s�T�2�w*sn͈��-�K3��g[Y��n�]��x����͎�5Ԑ"�X��u������9<��m��xorp��7�=�킜�հ� ;<���nX�=�q�z%�t����¦�a�����c;h�	���ss �5�~gǑۆ�X��'fL����k�^Î�j͇��9��K�Z��9�@����g�؇����G�]�P��%���6�ay��+�绺:˲�Ʋ�0T��ۀ�����o��߀Y2=3�jNK��[�ϵ�19�x��m��!��)7�l��g/���`���;�S�p	�.���fhW��g�F�i����t��^�@�S�U6Ͼ1��n@��463��\�%���Z"Y�V/����t�sx�f��7~���?�cC�heo}���2%B�a,@=��^����3��<��Ţ,!(c���u�ބ@]�O�5xL��q�+e6� �	�{���������k�Z�h��fj��Z���E��kzS$�v!���[�H��Х2�0a�E'�`��5= �w��wel�9��c������� ���ܟ�L9탲�ާmɎO6��m�[٫E]J���m7-�-��]�"	�{���_}}�N׸����M���ս��ݼ'V�n�4�%�������6N��7�V7O������2ζ��V��e�0��V�}Be�W�\i�Η�y��܆u�9��xxO���j鎝45�5
.�m�O�7[y��ݜ��.�f4sC�D�F�i׵Ϯ�н[�u��x~�Pm�+�'���@%g���_�_���3��D|A��P�r*z�cS�/y����-b�ǖ��(�����J���<;�4�{f7=!�CƧp�y��[P��@w55g���.�(	R�I..�*�
gO2�
�X������4�|m*҂����c�k�+�����X�	�L�lȣO���x���iA/mj����_ݏMC����Xw�ȕ���n-����0By���)�μ��C��6���%C���k^�0'hC����ڗ�bm�&�VoWl��
z�#�!��
�rϦr߰Nz]�|fl�RXw��K�\�@J�Ȥ{���6��tE2���cB~hw��B�߬�����Υ�Aߢg'��T���r�y0��0i�e�N������@dge�����9����D�]�����^�s��e%�/��fGS�W�a'��B����d]�n��{זx�����CkN�+�{4..���xf�>�E4JE��y�1�9@��>�摁嫯t��{W��_��V��J��6u�+:9;#p�|/[�9G��c+m�&��q���h��0�u�0��<2�m4����� @�0�_S�N�	je"ib7���9��:��KnB�ж�dS*�ZL�z쮉Zķ{��KD�������A���OW������{��xfh���ҝVq���h���>��A�E�W�� ���0�f���fyʭ�ģ������Q�9�yܽ;տ�~�_Ui��@;(���]�ń5�@&B��Z�Z�H��LJr��g�-J*Vl�˙�=��u�54�cg�2)3��{gO4��y��A|�0y��|k��l���z��oB�{��sμ�)�JS׭p�Q	θx�����
t[�C�0����W�LwZ�Iw�QE�Ԣ�pL�-4:�r����υ�4�PB��s��i�Y�o�w{�4��ƶr�]Ď�=.K�~gJ9��~e垁M=0W��]�!���]V�b���3�t7�|���(F���}�&9���2(�=.�Y�i*�K s@ث�U��7ٵg�c�k�^�f��>4�
���_�y��u��X�1�P��r��iA/t�L�!��W��f`;gzv-�1w�1l6zC�|�<x.��靀f�y�=�n�֗�|�����&5o_#o��u�~m�=r'��;t���l��:/�����%�>e�l���'B�{�X�p�P�ta�<�8)iv�8�*A�[��8ʹi�R�w6�vT�@��1�wݶF��yz�&[���T�� �\k�;V%J�u��DiݱZj;ҫ�:�Н�;T���4�]��E;���)�1j��٘�x|+���������<��7�7�x̲M����	g���N>�Cgp��H��xE1j�;c;�������n��	59�Z���Z�u/�z�Ce��k�K�$@3��j�z��yDu��g�8���Z�+����YQ�0�ļ4�ɸ�^m̳B({�S	&�Zg�ċز�=�.�-�0rwQ���:��'�}�^C�5��9�1��OM��W��!�x8�6ކQ����=�������A�c1�ޙ�`K����=a�yq���oDy��"Sng9��⸜��U�A�:�75oz�Ф�����ޭ�zݙֳ9�l3=>b]K���n4:�]��Z7��z̲u���� �R�T�����ȧ�xO��Q��4뇄���������v.Y'�1)̈́�S*I��5��\�Ǩu���n�z�fE:Wj���AS�h���Ͼ����=#����L�Eל�b�@��Qa�K�{�0�g\��O�5�~�t�j�Ѭ/����m��ۗȭR�"ߙ�LZ~Y�R9��њ�_G�Cr��_u^WYs&����$�­=�33v�;��eqĖ��랼3�nZK���4��},YQ��0�}�����7do
0�Mz�V�f�z�%��a��ѕ��^�����n�GqsC���FuE���v�������]�Kv`\p�u��{|��<I�����0fff�`�޼'	岺�m�y��fm�O�h�������������^T�'Ӈb���_��(�l
�ܱ��y�߇�k<���^����xǵ��dF��U�=���}��C�7��,����՝�8���{�qK:x�*���n��3���<��<�vN���:0�7��q���n�������dUщ,7���>���1��}���z��nϡ�h`݃�7B�,��F����,jelq��K�|��#rRq���C��	�G�:�Z����+T��ۋsZ_/�СG��&��粠��c^�{����L8%}'x���X~Ȕ�~���װ�k��L����`�9����{lN�ly��ЊvR}sh<A�]JgZ�{����42��v�'־~h���!��(E����E�md��\ST�hs�Q�����]���Y*�|���{6ʺ���{�Xt�}v��0ڑ!bg+��+1�r��j�/���7z��#6Ͼ/��qGT��k�
�?C2d.3ߓ����3��s5�+�[�K���ˬr�S_K��I�.v�m�v�^�U{��ͻ4�l�`��g���|��'C�\^��ӽz.�;9�}3x%��m=�m��ptFkF�g.����8'��o#}����o��x\�w�w��
.�::o �_cR�Ōz�ɼ��u��WH~w���j�Դ]�H=4�鑶�Lzm�C�<��k[c[� �o`v�cBѡS�t�ל3W�d�o��r�&�ѳ>��5�qs9��Ѳ.������_a1/a�Jsi
�JN-���Bt�ٔNU!�9��9�S�5�* N7�H{b�8�!�e5�ozD��ޥt�<�b��v��d⺛Po��j]Z*��vk��3 A1�I�����q�սNِ�M��E]��.���q'�֘��u�c4��_�W*�@�&���/��&~n��j��ca���*�JOO0��ٙ������PX�\�H�q�����M�y�Ȏw�x�+oj�/睿AUr�y qqd�,
ΞeV�����������Y�Cu��)Zv�w�+c��1�n�0�Y�J����'�k�J	{k
����6ʗ��	sF��}�;4����R��`�8?���4����]G0M�q*e�k^Ɂ:`ꇳ�uC.�!�E6d���A�ߟ����n��Gބ���f.h��.��ߏ��?����͵���H���:S��Tk�%}�գ,��X��5*�߭�wh��n�'����r$RlZ��54�qq��]����oB������G�[c\�m�hV��b9_q�h�L��?,.��\�1�*�x1P��ok(����W���f��`���}＼�$GN��"�I�y�=��{�3�+��0���Lw��zi��-����.������^��=�y{dX������0�ћ����Y���>�5=P7�=��L<���x���p�ae����n	R��h���Jt�*.��k�U��z�1<5^�K'��B��<�@:n鋇��,�wɪ�k�i������ݣ��p{.$E��<z�}^jE��"���1V��
JV?��l����W�ʞ{���p�t7��-�s��q�^�*�O����HL��ѡI�N��cO8�s�q��+�X�ߟް�̥�ؙ�
v`�0۸&����Q�����"K*�"LcQ�ʱeu�O8�/��XrL�B6s��<�{w��ڂt_*`$���ۙe�Fr���/{��yR��� eȽ��d������/�Pw0�����0-�0Ʒc�9��T��]ݗ}�~P�������]0�w�H��1�l��пu�'\�p���L�LX�[��Y�j�fީ��	��=���+pݻ��z^��O�5��.���h�=�X��'ntZ�ˡ�Y�:WU%��'5,��K��M��k(qa3Qu��F��n�+�jq���nb���6Fj�>�auո�P�[՗(�
�#�U^3O�C�ݪv�cګz�N�W�����@>�?/0�����# ���D�E w�|����o��
s�;��s!~8W඼�I�y����/��vJ�/Adk����܅���!�/(�=}�(K/Sӽ����pp�_�	�lT&D��ݮ�r���N�ti~�)����?W���p!UH��dlX �~��.��:�(�������H=�����8��p�!o_��cӮK��9�3�k�j�� �E����_�,f���ʵ׽g���|r�@fQ��-�r`��=��wW�htx��4n��9LRQ���L^a=���<�DԬxlm\2Cgd�k݄^�"�e�����?:�:T<,�⁉S{}'L�g_cF����w��v����݂���W"�i�w��݈��%�;WHvT]n0�ǖ�yg�顫A��-9��G<��F$����e��XɁh�� �6ꯑ�̭x�d3��|��1������1�2/b.=2�����y�k��+��9S�	��౵{��'�Q)�Z3�(�ǫz���u�v��P�4�$D_�O�,�w/v�77U����ݎ仲��;)�h����e��d�����U;>�ޔ��ͅ!}�x���l���$���R��l$� I#��b���
��kz�zE��o~�R4��+[=��V�4�gQ��N�so��s]��� ��̙z���H�4�هj���OmtGN��	A�BA� 5L�a�]s���ρ��j��qD��]���er�
������Ϋ��n��R�@�U6m)��W.)za0�J	���2O��Jr�	e�*Mmb�31$�H ��X��m}g�հ���B�=���"m~���gA�}�5*k������M���T��t�/7H�q%�1�,�c:e���1h[.|�g� �0�X���@�ô#�v�����De�?~TL^yG#�Ɛq���@������ⷠm��`?KE����i�s���Z�~��-P���̈́=A��j��oo#�*̉�uOa(�z�,g^���,q���ݓq���;ݾ�
�4�k��V+=���z����h|�-K�Jp�����<��2���~H��RZ�?m\7;_�)۫���ej�0��?K�G)W��S��|��g�Ο�r^��d�އ��jU����f:E�>5K��.�="�FO�%'e�i�x �\���nZy]��C?dm�V��������L`|Qc����_��#����Y���_I�b�y�.x!���\�/(��Aܲ	��d��3+6�h�;�y����9ceU��K.�����\ܘ��&��zn�&�pkFv��TQv+ܱ�v���M��[?[ �n���"U�<���΃�k�l%9K�R�y���G�Ib�гMԹO1��Q��e�����t��yR3*hH��M䳵^�\6�vG�&��75�V��Q���cev�b�W�:��#O��0�8�ͮs.-.�nͬ�®7"�ӵ���]v~ŧ�va����U�v�N�OkZ��T��{Ѩw����]�Ȝ���Y&�Z���U�N1]�uV7ڂ��G�$Aݳn�ѣ�Ҩ�}���x����Σ��+�[[�9��V3��#���2
��A��wUQ���Nɜ�D�:�oa�o:��\�!q��K�J��#{�ś�����5#��kqKQ�ȍea�ñ_�Vq�6�r�3��%�T�Y�&�&���wb<
�V��ދ�T��f�j��r)��ݺ#7.ĩ2Vۭq���GY̔b{�)���{
��eu�;���ᎌ{��]��P���fukd�5�FQ�<�Xp�>ǩ��5��ۃ�Iu�{#���c�ȖM�,H�p��Zn�6w�sl���m�E��O3)n��Я!F���1�f��\�޷x�PT��X+2�)!ީ�Y��y��X@�ǏⰬ����KҴ!�0b��`�wj�&���6�m_��ޔDr�SjUFE��H�A�;!�Yij¤J;�;D:�w�8c�cXٺ(7�R���J�!�R���۾�sy+\�{Ej���3:=�1�%*�|Do7<�7[h��R�{Q��gUN�"W5�\����i��®U�2!�Z�]��/7i�R�aZB���Ɲ�MNuʙy,_�e����f�X�YAVB�l��`z4�ì�ܡ�c]h�e�U�6�v��NQ��i����nTl�\�ㄆh:��od�r����λ\e8w��o�VpP��o(?�q'˫d��Ѭ�V3��Shv"I�ՌȆ�wi�gFK�Ki�i[YS3p�����Ӌ{��z�*�jWX��}K$˜UE' ��}�iV/ܯ��fP[$v/� �vV>�VfK�NlC3�ja���9ɻܛʹ��Z�ɻ�+zY�17�x����@���zV�olSb'*uvy��}�ػE�M-3�����k��6�p�1V�5Ou��|�m��c�	��+���Ī�����|������=y&�C<]B�L縃f����Y�v	1��2UCu�,���b-�iݚ�$D�ǈc��j�e �GZ�?v��/z��0���e�++�j��rt�\ݛ�7�nt�d���<��5���Oc����,`Ujܲ+���~z�2�vE�|��V�GG6��8�)+˷�[������ǎ1�q�q���8�nݻq�<NC�e���d!$yi��?�ݓn���yהm�����_�;C��;x����q�q�q�8�;v�۷G���,��ul	%"j_wN�N�/쬊(����s�i�u��Z	�g'�j΋�=n$��$�ߏ�.)#���=��GVVyZw��W��ƾy{c���h��M��[vI�U�%f�q���o���iO_�U�k!j�GvMj�ms��k �K�vE�Y٩vn�]gY��_��"/ͮs��.���<��],������:��(��[$Jj6!���F�\u�\}����8 ���N�(��3�=�+;�"}����K�Q��vDu����?7�>o������R�I�¼���^&"A�DI�5�&�bAe����򫤌����j���� y�y��R��kou��Oe<����w4/��}R�^����˺�a$���0��aLY)#$j$�2"�l�jy��)q�A�Ɏ@��2"�@|��(I$"3f$�-)a�i��P��q�.JP׏�x�����M@�	0�.��ܙOn��矔�[�t�TqR��x�Z'y�q��d�?Y��>�Z���U��X�o�ba'��֜�G����"�!ǙZ���U�Övj�t/�pi$˴�ִ��O`3h�����{�d^��J�Y��k'O�����#s���C\+%^��B�4�"h%�ю�S���T��㻴zjS��.�IWBƠh�Iu�'�&➰�_-��37���)�;݅,@�b�-_��k��hU�O
\�J�l��ۆ���q��k�ݖ�[���X�m�~�%xW�Y-���0�����k{���7Rp�ݞ���[t�̑e*r��p�ލ�H�E�`��y�3z�9�ѫ�߉��[!��ϳ��\��0�>P�yi�u]feݴ�݌Xz.}������5}@�#[�pZ_d������ucŬ�%�c֬�����\�\گv.�7H�]���J���o�7Wm��<w��և�����d+��q.сγ\����<�nq[��+1=%Y��Gn��}4�x�f���Ȭ�]6FG)��N.�ˤ���-�J�_��^���ߟ�?Wn�3S��9e\�8h�m^Z�S����d�_k��k���z'{�ڽ��\I9���<y��.%
����uI;��B�zj��*;��
�L��:��X���#4^Utu�\�=И Fl ��;�p��ڧ�e1��|��t����Nu�Fs% {6s3��XV9��{����h@�q�b��<W?v��<zݤ�NլY�甛�&s���Vb�Ф��2��Y�.�LL_8*D�i��L3���wmƜ���F5"I/�=��������<*=��	Wo�έ�t��V����F��2�7qH�H�İ=�����"����pc]ݽ݈�i�,�p����ҿfV.��jSʈ�=^O^��R��K��3�F.���Sm�;�F���NP��L�bSg9��h���\��a���=���Jg������gB����wz��L��
�ݫɐZ7���'�|�]�я8�6��jiԊ�>7K&��L+"+V�ٳ��s0n�o��va�2�F.������Z�'el�ӧ$����*�^�Y݌v�+,�\8SY��15gL��Y��Yj24�x"���D�Q��*��v�G��PJ�y��c��]���%�P�'��_�y��#�3s��{��7&��<�r�y���؎�5�d�!��x
��ro|~���ޕT�h/��Q=�	*�>�϶�@�g��H��L�dk���[^�4�ަ���X݄�RR�0�yl������u��7���X�mve�����N� jQ���7g��ia�	K;tw_�y##��1J�4���}����DWm�ɣî<vs��kU��9�خC[LmH��V{v)��b�>~�ֽ�Oà;��F�F8{/��R�N���,�
?-�"�Ŷ���>4ی����,�{K�
3�u%���������ݻ[�2M/@5Y>ڽ���G��e�d���tK��Gwfn����ܣ	�Tt����B/N�V��Q��V4�����
��u}7�w$��\$H��м��h�Y�]vi���]l�]u�����]^�r�N߆�#�u�;�� ƞh�kZ%�K���|�{1	u�N���lT��ͱ���ハߞ(����bI��?�~ꢹ;8m����\��=��1ʹ����ۗA���r:��:��,����A�tƜ���b���V,w��jo���}���}�I������MGR���7ϟ6u_F<��܊�1�B*�м���>�����������N4��ίǷ�ͫ,��@!�6#��hI>��4�d�m	��}u�3Wz��>���"��ի{z�fڐ7'��@g�s�#�	Ps�ꥇ)����UI�;wwv�=ؗ��+��
iA�OZ=w��Ϩ �@�x,��kk�P������`Oƈ����y#*���s�a�&�B��P�sW-��q�&;w�p�-�_���};>b���o�a)�I#M�f���Ň�m���t�=�\AO��?��j���}[���29ۛ�[�������뭥�YΖ�fFk
�C�Z����'S?��S��(n\z���.c�I����?F�
��~���r�}��dǳ��^Yv����;��o�U�PM��ɦ��v�l.ϝ�|������Uf�c]!-�ͦ��� Tã��*C����G��D�o��e�7k]
�O[؃�]o6�B�eUG�r�KNT'`��x�l���U����}ԝ:�H��ݝuo	�i��"�/�0t�܇�H���n��:���b��� ��<�ϟ���`�o0��!ٌ
7�_��*��{e̝ہ�{���=X��Y�����ks���w�� N^�?�����V�6B��#$����t|�w�����S׹�i7���= �d�ށ�;CZ��YZ��38����p��z��F�m��ϲh�c�	�[����W��sw6���1�EPe�&q��:����38��5[�g�;��vo��ob���!8������y�w��4����M�f6a�U�v�Ɯ��4O/$�.bw{جx�=h�`���h�B�i�$�F���`	�^�����R�y.YJC����V8z���g��syʟ1�w���m��7�}�O>��n-%uz��*U�4��.)�GgQ�ѕ��ݛ�[�3q��PBn��:�;P`�ƅf��:���]`��M�9u7k�ѭ�g�>���U7���ϡ(��pyŒ9m��쑧�V=��9��?X|n��U�
��5sx�z����;��
M��v]���������Y���Yu��}�h���/P��w.L厫W�)�'�8i��(={�5�����M{뺷�����ض��������Ӧ�$$VH$���Mw�y�����o�������};5 n[���١��\��y��2�j������~~��̦��?~��e$N�{���v�F。�r�}�4m>���OmmF��9���ϡ?���@��7�Ԥ-/�����4����%{'������wMb����+������a�7(�K���I�q��5Hh�=[Yћ�y �L:;����w���L-�Yܦ����Y���m����˚�j���L����q��v+0���ڲ�<Rח��qMU�6���q[��"����ͼ�M���hL�#y�*p�{�{q.g�q*�x���0N�wU������d�4��ν;�ª�.�*v*�'n�Y_X���wJ�H9>%��7^������Y>�ۍ�i]bWg��(�;X1�wM0���"x�����:)�b�����:.�?Ϋ�ˣk���u���j�M�W�.�W)��N���b����90�$���6�a���sŇ�r��T���pF�ܔy5ay�d�s��n|�d9FM|���]����/�r9ER<�'��7���v̩P�����|��?�I2:t�QH0$W^M��9���3fHI']��]�R����Mi29Q�M7��.�Χ��\q�[��<�K8�[w&�?*a8��������if��벯����I���=�~�ۄCLi����
ҟ[_	�-C����`3���{zyw/_$�h.�m̑R}p�^ǐoBٶ=~VB�Ó�Y��r����3y�{l�� H���	�����Jۮ�Yw����G5���Ol�����Dn׸^��}% ]d�Jm��u�=i���=Z�e��jZ����8-~�b�{���{�Fc�깾+�6��������^j�~'{�b���o?���ӷ��;t�Y؞�Z�#>8��M���N����+\�V��p���Y�~��^���%z���L{3 ��ޑ�٘�i6�A�{��7��ۈ�"a�O'b����*�k�{�����e%�����TΑ��_���qA��B�.=+�;�j���h��J,%�I
�J"���{ϥ�]g������1���Zc��4=e峕8gc����뉬���+��qX���6�Ml~5=����������<���k��H������\u���U���ۻ� �p����{eH���t�}�ʝ-��vO��"�5���~�/ޞfB)��U�*���Q����g�,Xد:���ȗ�����qt��--��O���21�Nv��n� 7kr��w���)@ѥ���_������i�iv���ˡ5�;��ǹ�JC�^��l2Uǟ�U諓^�w\��Kcrj�Y���5O?v��j�en{]���W�c[�|�Wߩ��U���^\t����gs�ϫ��e$����}t��P7a��em�׻��c����z{vά\_� ����=�>��2G��
@I��s��k3�����=�!�u����i�
���FS�v�}��=,[1{�ޝ���Gs[���F��:/�G��7�r#���J�IQ|�0aGMܹo�����	�������B����jа�c/������h�!����1�kT5�;���˞b���u%t�u%ڎ݋��}kf���Vֲ�GT����<����j��ʦ9�#���T�7���s�:��}{k��Ӧ���H�Ͼ'�~�z徎'�
�ϻk6�(�V�7�Ŕ�L��ia��������t�>s�zoy���@%��>�jl��=��}�ս�ڹy/-Tu�<�.��Bَ�18�v����E�mb5��^Gj�Nlyg>Ol���o��.��O�?I�7���;�j��{3�p�:lH�H� �t��9�z�k�,�l�]E���O
9�pڏ]��ڌF��&|����)[{w��� �d�:��<�Qm�h̨}�*�l��!�~��wJL�i��>��{���mcv��z�4��{8q\���A>k��a5e�6����4H;9���*����t�M�ɠ�=�ϣ���;:���㮊�[�zo1ꩠ���X��Ix�fX���ߗ��'�[�!����
��Xᒜ05��m��W����F���͞�˱P�8�>��Bf2_S*�
�h����[X���Ax����ܣH�:�J�P�rmu�WC{;���/�]-�
��u��}� Fb��7�w]������QJX
;s�d;�0὆!{*wf����2Ÿ�b�H2�bN�#5�<��s��g�̒���z�խh�)$��uw�qm.���)M?���]z����i�.��Z��Cf�s��u2���]�Å؜/U*�^�ZJ�� dQR�$q�R��sz�V��{OT�縁���������H�[f����[��H����n�ޮݞ�Cڳ�g��i� �7"�\'!^o0f�7�����j�Buӳ�R��s����RC�]����ĢE���<x���U��ʊ̧�8��k��L��6Ǽ��ҥ"@�6��G�9��K��WTu���]sDs8m��1��*��hے���#R���v&���u��4�M.Zt'�Ђ`Q���j�a�t�%�t�С���t��Xz�Y��z���a�u��̺�=צs�˒���*к�܍�����+��w_d�)�qI����\�-���&~1�زG��7�����U�]9\��j��t8�v[5���{4c%eP��۫fgc���)�B��B#�p��+D�ݷ]��g�:��4��/}w���CA�՘+0���c�(8�
8�+F�����ot�{c�Ǎ�
�'ͫ���43�(>в��u�>�k� �
4�B�uo5wd<7��7[i0��A}�]e�8L^,�j���xk�t�
w�8�|
�bܺ\�]�6���[Smn�oG<[��P�]\�Md��u �Y	ކŔ4��xx-z.��\j�]p�]��^�g�r�ʛx"v޲t�U�]Yk;H����Ry:�9���y�lL�ڢ��d6s�e�׼�+Ԫͅt���Q�l�����n4��c��î5�V��qk4;X�Rx�V�?l�i�Q.�Q�-�vR嵰*�YAn��-G�f�e�F��t���z�[���WGv�v�2�u�ȫ�MT���R��ٰ��[u�JeVA�pێ���k�|� �ф�7t�3�
�Y�F/f��q�X�ӉX�
4_�g�d�v�6�a��;z<��Gl;wU��M�n�kS�7�g�/c<�)5���A�é-��c�e;�ǧ
-�����Dk:�_3]��j1Yɓ���՘�pݥ-4Ų0'k)i���Lv�%G�=�:��=�7B�ɹ�QuE�`+��s�P��;�'�{�iY��AT\6I�EwJ�a�A;���:�y��]rUu`��=�ѱgC$"K�P.áWyR�xMnl\^@{��8��^s��I�<��j�U�i���Y%>r���|��{u#��ڋ���q�YU7�c�F����C��[�m��{��gv1�.���;;4�!���2�.�"��$j�f���՜���#��\�[��K����]���7���^���UA��-���n+{1��;E����6��oQ�z�$6�ka��R̹!�E�m3�n��9�f�R�Lq.���K0��o�q��aS�ݭ[ӻ�*�fRiS}�TA��]UO-@DA���4�K���ba᱓3�M�Oz�%��-��*����k������+�9B��Ir�{b�,$v��u
4��-C}�"�_*��#��vn%9���Z2�.�Ҕ�M+�J(��\0��^���
�Z�<��]S�n=���S�Q��MO����f�"X�i.�<r�v��
O2��U��I���*Y᳎�RɗOw�U���;�uu��7���f�Vv]�;���N0̦X��5%Q���{d�i!ed
l1��=5�q2�h>ut��kTxFI�{���t��[��v�Җ)1�u\)���Fa�:�,�z������nHs[y�4��r�9P���'s�k[�F��$qG$��Υ&��:�����w�����9��j�H�� �	���I
��F:t�������8�8���8�nݻq�x��99���M����6%--� �?;v�����q����q�qǎ1�q�nݻv����du�!�<���#�����:

"���/���۳N�ւ_kE܋�7ov����۲6��Y?uY_���W���/~��sn�����Q^g��8�^��D�Y��5�:���dS�Vt���転��xE�����w�G^���2��϶�Y�]�IOk����^�gO�w�DG>�n�w|����+N�{\uEG|.���n����='�x�D�����m��h�cRN|�òp_]X���j٥u�MZ�w��i�v1U�{[�����}`�z<���5Vf�W"���s87��N~���Oy�[?�oK�P*��Jpc�\��e$������_�Ц)_���<�����e�p�*�˼�ZӺkz�s���ny�oJ&$i��a��������z�P�ֱ�j��g���;Y��h�qwM��Kx�<KG�
�y~3Ӹ����彝y'N=;�(A�Ѻթ��S�3*���<9Q�<��.{�h6�=n�usL��E:�k	�����(ؗ12�>��&8�a��et����Wѝ�՝m7��\ө,�"�� G����`�>��
�X���'$�ӝ�������L���ۺ�s+����ɟ[��^չ�-����㥣r�9����=��H�)��w#i�	�fQ"G\v�SL�L��:�w�t�D�A1\���	.a[$�Wy�=|.�\5o�lZe]h7���=v
2m]^8��W�yպ�J��;��\��o�I��f>���aAu\^n+{pöF����g!x�n�+ܪ�
*�&�5�M�mʳ� ��vMP�]:���{NT6�����K\�2����������e����<���{�f`��9��ѵ��ȏ?|_�_�����4��imҖv�X�U��q��w�u� &���p�,�ղ/�ϫ�@��;��)r�=�/-&y��j�+�7Z9�ѼA�^�9Oeg��^���s�т�CY��Gv���fc[35�Fs�Uq9�����'=���O���i
ه{�����7�q��?f0�SH�os�')n��u��{�䵇�����U~^�w��u{>�0#�Ĺu/�ۚ�0��і���)3�����u�gh��I��3�!�[c	V�z�xg3�|nG��H��7�r��n\&A8����Ց�vw�9�j{�1.����k�ť X���s��&IC;:���u�p&Z��k�q"lR��u#!��������O=M�y)N�N����b.Y�����[���hW��[Jz)�FK?�t��8tu�!�qmA���l�"b�/^fQ�Ѻ��1s9��,�p��Ez�螴�{�̙�jx�v���ǁ��t!㞽ت�{ɩ&U�Ǔ&���=��J�4�^w
3	���*��Gf�@�m�}�ɫ��n��cZ�=7���;k�N��$����2to�����)7��ے��+�+Őm�l��Ez�n��ٮ��ƾUጔ�[خ[,l���1v7ȩ����'4f�S�ݻ}�e{9���v�� ��I�{�ɺ�3�+n!\�l6�c6���hg>�Ȏ�=����m@���y#*�;Uydlf��GY�M[mnf�t.r����6�ʔ���r��rF���*Q�vl��}��kn���j��ꗋ�>J���B1L�5>��(�T��@��nk���23��:9��##=����lǏ��L޸G�F@��Ow��Y�#;牯M�3�2�*\��Yϝ�+��]�f	{������;$u�UV�]�w���A�[рm���2����h�-���x\�nh���%�ɾ���S��U�`��Iv�������M���������y&[�mT�f���V�����q^���أ+_N��մOuQ�iQ�L�ԉY�N�!�L�bG�;ھhG���:��*e����*zw����ݭ��_��.;M����+�6����V�����Ҥ�E�؜q�eE�l(��)�����Ƭww'C:�?_D��O)g:�DS;u;]*�׆q�mރ��߼��|�����o3�GuaU�5��۾����0&\�U��(��[��&��n=`Gqʳݜ�/&���6�O��*gU�#S�24ýk�jg�nz�𬈽ݸ]}���v��|@����>h�L���=������L���/���=�ͽ;~Hfw��rGԊ�Y�u��:=;�X��;�Y��[{4h	�N�s5OE-���B@t).=K?
�w]t����ڴkzm�x�짪�B-t��ԕׯW��(�If�i��!n��{���n���aS���5�;_�QR8.�d6�9Y�q<�><�;�=��/�}��8�F��x:o�m`����)�Ӌ8��Wf����U�9��}��v�9�R�y,�<{p��]ّ"�.�����!q�1����ӽ\<�6���o���w�?��"�7JH����w����3|kIE��������醦���#:���=���מ��v�Җ�cɔ��pmΩJ8(������7.nwȒW������u��K��H���L��k�Eʴ�w��vه&��-w0��p���z⦪�\n��-����}H��F���I$#;�9�ϟ<�>k%���S��}F��6�и�6��֝zE��k�\��Z���]�ʳ�%���7�Q��Z���ݤČ�F�ӅY��'v(�CxCy��e�sms�i��i��a���TBR �O^��\&;��kD���Q�෯z� HVG��M��P͆��d���O��2���}����|�ӓ[�y8������ߌ��Y��s#��~�oW��j*r귻�{#ɖ4w6="_������h��D�i21���ρtf�����Tcz�M�o���)�V��2H9 ��[�^�;r������f���֖G�����'Y���wh��d]�����Ŀ��%��=������� �*5:f~ٝђ�U�[�j�ɜ�Z3�UQU=uug���N�K;A�9�:N^��VZ�^��8�x�����?LM�W���n�w�.g|��u�P��-��b�*@xڟ�x�UJ���%9{�wm�I�r��w^6]]'����:��v}�Q�b�hw˜�>;���m+������� x�����Y���K�cQ��	�Ζ��Ի����V鳽����o��y��|��n�bWΖun��V։��i���][���:��������E^�ݼ}�Y;o[d�>��>��\��*�#rv�D���p��&�FN�/qgb�������E�@/��!�����O$�-�ۺ����n�wٷ�E�Ⱥ�'t�[�(v���/���3�)+�F��3�IM�����wy3�k�f����;�Y���c�V(�-���ZY�V����]����饶�<AW�:��ݣ�[w��>v�k^jp��q�n�ퟩN�ŋs����9��G�^`j�Hxq]#�?#�����7�X~w*`��;�i)�M�\��a9��t|,�D�Ή'vMǗQ�m���6=� -�:!3��X���7��͛�;�ԉ��*�3ߟ�������r?�i-��y��q<�@7]گ�wq��OG��0~����Y�-k�xa�cYE7�ユ��S�9/ �*4my�P�����?4gl�����߯�j/^_����5��Z��@��@�cwp��j�V�������Y8��[z��1�h����IôZr믤�����{9�G3M�����<�8�0}£P�)���[���[���F��I'T���9E3(�Mc� �}"�-v �Gy�0wFG�ۚ�i����?�ބ��*����U	�����T,[��瑺�1b�8�ݺ�������+)��R��Ng!���nI<�v�B� 2`��Gvwv]�+y/$! j��S�~���X��Z(�
�wS�og#�+I=��dqv>�2+PS�'֝#myK�=t�=��xs	�2��P�q*z�6���lP��f�Ƥ׏ ��'���g����ᕨz����:��X ���
�E{T����p�@m�Ue�*�.�=7����w�6��=Y�}���?��jD#��ZwA����2�{i	.�ݙ6G%ט#ʬ��6���y֛�r�~
%�����2G��K�lb=�z7(�4d�'�Q8Fc��pV�-��z9�}nE�I��S���<�]l9��[�c�yx�����\�� ��ɫUWj�AG.��])}Y}f��9~i�j�,��ӕ������a�����)�3�j�B2juF]#�����E��Θ�6������8�Vr��}y�[qN�������������b���YS�{�<4m��kƽKH;��;���w_����iiy�ܛL����۠������6����@���jƂ��-��$2%��;'���;�¹a���0�[w��$�w����w�-��u�kDd�-�7lO�ŀ�f�P���b6�S��;͵�	&�sa�P��T��m7�Ӽf�o|��f゘~�k�'�'��j|�^�$N�yl�n�7������K�/d@����� �K�S����+�G$�j�@U޶�E^��{w�Gn�9���I����z�dd3����цG���i8���y�39��{�K�����
|��;ۉ�烣ۨ0]a���S�� �vM���qe.�!pJ���Ee*��ѹ��3t�+r����z��:�\x����
�PRT��-��gnRN��J�������ce�>��+�I��v��}O�B\�`@����2D��{g����d#ѝ�k� �D�M��iH{6�F�5��N�F�ݎS
�U^�^��A��V9��ث�me8�e�8;��ge�<��y��OW�yy{�h���R�x�\�Ϣc>�:��s7HT���d,L�Yk�����m�Ξ�U�=B9x�W�fOM<�P���4�ra*3�x��Z��S�Twu�Ʈ����B)y�5^|��uٙ"�%i�5��V����<�G(w�pf��!���1\P�Z&|�`�Z*{�pn���R��w>��=s<x�`�y�ۥ
}[�;n'��4}h�m�+k�6���Qո�����=��GB����=�l֣T;A�GB]ӷ�!�S�h��3��zz�^�����}Mp��x�սP���=2r��~��W��SR����M?�\=ҽtT����l��!����y�&`�jL��.Ս��\�v��.�n�u�gc�I7��<ʓj``eJ�sl?��O�M����Σ|�¸��vrw���'{{I^W��y×}^�l��k\;ި��e�����d]�^m�P�Ĕ<*2��=q={f���Q�^�z��!�+�M��RV���$��d����5z��i�"ʍ��zoTΧR��hVd��{�9��W�S�9����h2A*��c�y���_�y��|��u}ˎ2�~x�ub�>Q�`ɏL|:�.;��r]�O&s772��rj�_i���
>�f��֞mm��w޷ݞ���q-�[�F�U&4�M����K��`�##g�8�b��ILMOP�z���zL��\.��H�I'�T�<���-WT��/�����g�칀�_���y˓�gA�9$�}��rh�=myF�\�6�T+���r��}|�_5�1=]~ֳ�e{���޴�Z2�B7'n筅\��0���0���k�v��S>�������~g���o�Wv�@�=�䈄�1�z�3��������9��r�97\DV���$�1��nɒIO9ܝ�bwY������v�i�^� �-���H���>�l�x8����Wފk���=6!_��CY�x ����#��o�`ɐnq6�e���p!�w(^�v����M�x���(�ڏa�7�'�ppw���#m��s�Vƚ���N���
�P뼃$DpO:�	U�;�k������"�k�<ŗ�:���ų0'��F����kB�m����K������BY5Q�����d�Я��L��uƪ�2>��ٸ{L1�R�]��z雪��پ%=ZmjX{R�ջ�_lUgjn��1=��Hcc	��H��o�,.��r��|�=����[-|�f]�����҂��sZ�٠�*ɧXm�wg��~N�Pm�ڰ����pj�s�*j�+�N٠�Q:�/j��J�Rc�S"��d����[>���	��8k'N�zw�6�>{YOrŷmT�ٹ�^t��ȴ�t>�.��n��)���=�u|�kZ��6��N�s
������#�5s��}7���^�v��-qĲ�J�LW��y˼=�S�p��U��֪6+q���es�fk�S`�Q�Ҳ�M���M� +�O'[����Y��ۦz��v�-}���޽v+��OZ%r[E��7������ڜ�}AY�.���Ӧ��n�uD�"k��,�0L}P���%�H�F�ר��] �>\qg=-���x��'_3}��rÕg�(5��
��-s�*Y<��r�08�R�
�3�F�_5�8�O-��V{��?5�I"�Z��c�Ӌ�P���[T�d�;���N��4�:���+h�,]'�bx��^3����(4����V#=<�o���J̲r�v�Ն�s/��d{G0��z.6��[�iν �,�˒��ŶX���M0��)4�����Gr���ep�o:},͹M</r^�Vٌ�#j�.��Ņ7qԾ7r�zb�=F��s�;m���D�1�L�]q�ɥfJ�naI��.J�Ct�[��ty8^)H�Ս��]W��Έ�v2M!*�4�ձ:��ĵt�T��J�/�&�H�[�Ҡ��9l=����������3��v �9��s�ht���i��_@�h/+l�ۈ�I^�uj��E�=���iAui`�oj����'ye0�n�������G&�n���;�Z�9aQ���xa��f�*���[�u�^��%��[-ɄA&mK����Op����xT�7I���V}���c��b�x�a�S9*j�VFj[��T�zZ�qU.�'M/#�
p���ײ��%9�G�����UXa�ά��\�'4��4��}X֛A⦮Ⱥ��pS�z�db�p�v*o'lX�A�w?�h����UC����&P�J�F��oe(���9O��P��%_sR��un	v�$�C#�uM|AbW7XB���l1'r�ي)6jrI�wI'-�H�NI&��u)&,(6$t���H��}�{|����˫ܿ�t���E�gP�,W���OoOo�����q�q�q�v�۷n>�y�،���c�D��,�l�P<���>5����������q�q�q�v�۷n>����H�!I�~����{ug󬸻�@���:�"i]IF��t������">qYq������u����.�����u�W��-��,��,�,�w�wdwntuegj�,�8��N�����w����~4K��g	�|�U󬳢#��]��Y_H�U�a�e��j����ם~�+,��¯�ue��"⎨��i�~lI��#��8�㨻���׿��{��B-(�d�Q����4D(Ph�(�q�	r4�ڊC>)�:��O�ͳV���Ɓgn�I�TU�[٣��]�	a�W*�ߦ��E�Vk.���Vq4	�l����(�)�>�iAI�׼|�H�d-D
,��
R9A�ِ6�l��m&S�6S1��3�$�A��!��E�I��EF�%����POC�!u�mֿ$��yϗ��_>�$�~Rm=��.�AR4x�M��2��bIm�y�[���V�vm�Ν��r%r~Ќ�����,��3@��&%�>�W'#di�קw��ש�.*���bB��N��	���p� 0��:9��}�9�:�.�o�n]���:3Uw%�䜚�=W��w�!��d6_�w_n.@�
�;T�ˊ2�>��|W>��j�� u;+�]��~�U�;��d[̜"���xRg#��]�˅v(��Z;^�2;�fs=��k����LѻmޮΞJlUώ��ƻ?����E�I�E�6/n��*������"�����@�U���	-:+u��2�wWC�J�U���U�Nk��ʼ��C�k��%�����Y'o�Q�z�ƃ�[���O�ŀ���S�}ɽ��إמ��6�s�V���i*H�Nm���:�aOUl�-7�K*�N�;�!��<�ٔs�j�I
�ǻ�+�8OZ�م��^��E��O�u%��2�̆�V\��"Y�{�hz!Z��*�rΨ'ղ�]ʚ�Y���3�K��:u�U�vK���k���gw���F�r�5��0�U»���-,̶ҝ1Ҩ��q�a,�]�5�ez��>o?��j��u#��i��F�5��к�N��l#�x�F��4��K����ꣴx�v����Q�n�U��I�;{��{oO���TKv#Y���.+��"��y���Q]1!���DM*4$ު���H���J���9����7�w�v�-�'�u��9��b�<i�L�����h�ۯ �� !l�yL����'u��� �D�6Z8��M.V�ag>v��rL��*`6�S'���t�n�#|:��[��T��g�mj�kc��<?"���;�R�+�2 ��ow��9"��ހ.���z����?�����
W��Ɠ	�O������o^g*��5L��`F��a��"6⌭}8��mZ�ZѬ�?�:��Xb�՞;���Z��@�k/�A�'������ڵ�����A�D���d�=v����"ߥ"o�= �A��N�g��vu].7 V�a�k����1*��I��בϟ`��q�2�}(h�w�H�9�]��,KY��t�'���:G�PB	3Nfw@���^�W4G\�n=������kazn�1�X�ۋ"�]bM�*T��}����۵{�/<��o|�7�����W>?3�Nc�p���)��w
� x�X#��U���g�L���U+��CN��!�KEi�j���2
#O7,���8����r�2������j��y���H�^�2U �
v�Ɓ�93����sD��?��Oo���FM���U&��}t�R��C�����t�<�{7��L�ߜ��i��̋�u jg�vםAw�#�q�{5R����pg7=��@��9�b��(<��GftK��8C|Z�N��D�}���6�7��{�n�[�9�$��$��S�n�ݙ-$�����WV�w�A:"w�v6rEXn^���;~[~s�4ה��ϑ{��� )���킕|[�}%�؛@JB���(e�*4�g�6ǮN�j�!�8$+�� ��N���֣U�z�('��zjΚ�l�9�;���ZI�}i<{:�?
�+�8��vqz��8Nl�(%|��:�열�RR\�.7\)�3i5���Y9�>�o���n�-���4m�uYx���[+5��k[j��=�ㇺ�
���W��<�o|"&�5�%�Y����>�[,������}[����zs���Hf�GnOI��ٽ�ؕ��4n�&׏�=6���!��s���OLv�Y����t�������Ƭ�����*k� �z{��D�WA���y�������o>.�T�L�ck�͌.��0��j~������^�q4��܋���b��lgrͽ5����	����O��$]�I����`���*�;bm��<v��Ǆa�!e�Iȿ[#X1��Ӻ�/Ȑ�;D3wlś���wvs�bH
oؾ�X���৥�{W�%z⎍a�3��!v�nH�f�EԸXy�6+:�rν�5��{�e���*���w?��?+���]u��.�^Ktc�=������j��>�F@'���3���>n�4��!2	�w��y��Z����.k4�����M��@P�)U�*��{�V®��c3;��o-����9�wv�mw���/Ðr�k�M_�׾-S6�o��N�߫'�V�����W&(ܖu��� `8�W5�4�l�[�0P}*:�nPO��츯5��Q4����-f&��'������2��H�[�-��Ypz|�����';�,[i�]��G���I+KfɍI�o2�!c>�BS5�,#��h^!�Pt����[4�0������`u�Z�i�)#3��y*�{ʛn�Ĵ��b�{�2������ѹ��Kx�f$.�t����{�%~c�ד������x�nO_�P9��O�æܜ��Q�e�c���hL���-�'ɓ��2�R�dI>S��_��Y7��r�	��#�슗ٍ�Q������z'���a"W7�r0}�`��#����ge���,�k&�OU���~~�"��U�+ݍ�;�E��h��4?BD>]?���5���d$��x8��;Ҟ}�����V�D��T��7)m�0���ɋ�8��|����S���w]��γ ��t;��z:5��E�����S��Lt{p���+<<��#�;���K0F_p�Wb�G�rҾn� 3U ���!��ս�8n�$�WaT!���u��8F���]���6��^G5~L���٤װ�W'��	Y��t7���"u2��݉>g"멑C�Ǭ/WymOM;)��J�Z4���T9n� [ŪpU!���(39"��p�gi��)�"����F��j7�r[�����;���c���Q�Az|����o=Nݮ����O��K�"��#�Q��~������WK�IC��Nr2Q�N�1�P9�U8��O���G������z�f����~=���#��R��5�0��0�����)�_�q��mʹ�)�~�X#o2���5�Vą�4wC�̎�f�ǵ���
Pd֎OQ4#�<�#v�����i��~"*��B�3�,QP�[�^�&ґ��TІ���]��8�7g�����phU���sN���,.��<-�tr/��I��+8�B!�Ƶ�9D�4�UO��.�ix�>y&o8U0ĳx���ۍ��Gy��`�;̽��J�,�E�A.<M����+JQ0�O,�����G���Y���΂irU��vʞ�)�&����ɳ�ǅ|F���L�G��	�26ᙃ������ce,ڸj�WO+$0S����r�TL�-]��51�seG�
l*��Ʊ���7itӁ�-����B9o,1G�NA�]X,vk��ŝ�!ȪS��� r����v�yI^��G>�ά�z+X$2M�NT�Z��ct^e��tжj�����<�o}3����6��aQ?4����;�<x����I��h�OUث���g��Q��=7��@���Ľ9PX�g�!��z�$_n�FT�Ν�.�"�f���g��uf�wf�SFvGm`���c|��[�����l�`�E6���#���{s<�iY ������"�������p�W5=Y۫4h��0w��dB��0a�7�}�8�$v��{h7c��)J�ư^g�o{��(��p���N�¬��=�s��P��<��mU��p���TJ������c�k
�`���{�כ�OH����qX�H�uWa��O�o�z���#Y\t���4��UWX�="��RK�0q���0����NtQ��l��Q/��\����8%�=Զ�����C��tM�+��P�#�M��yU�藠&��<��|���g�U��I.����mGڭg"$K�(Q7�����DԮ�m���ǖ��[47m+{�D��9ٻP���=uo��*y7TЗ[M��t ���$gt��&M��ʍø�C���1L�J0�Zw[nAA��m����>�7�MnwwV�U��Iܐ��"��\S�i��l�.�ݫl�"���X�]_N��r�|�x@��݂��C�RI�����,������a�	z��W�&��mх*��v��6(���?ߦo*Y����l���{�v������e��<�p]@D�C��>�E�]���]�]\�r`}wѨz~��+c�}}'K�Pە���Zַ�/�UA�7�v�7�%�ۚ׺���9��t@���7��U�G7���adf�vp����1V�zr��V��n`���X����[`A�wZ�F��i�%y����Z)�l��Zv�;��q[@�];�s����W�=;@v��I���6�(�����tM�|=�y�!�p��/jx��YH��g������������QsX��K���Yg�4�E��E�9;��lh׻��78̀�j~�K�wD�/��l�Ug.��fcu��#Y��JKM���]3q�9ǯ�w������Ra�Yz���g
l�&m|0�:�Z�$Ce�͵����Vū��v,�h���ܶ�o6���d�t/V�Sc�b�q5Uv������<�o܃�G�p3�v����W@�6 �zw{V,fb���[�쭩��p|���>N*5��E��������O�jz��c����ނ�q��Vwv[���Kz��<��{����#�� �=ܞ[X�ꩦ�6�utwU����^��Q�-�z�o,��9�jB�(�ek{b�V����!���=Yۀ���I�P�Ҷ��i�Vgc�%�D��͇�gH�T]�&��@�G�A��и�H�J���ڋ�ge/֪�9����f���P����!*�q{�s�%~c�c{D�|�l�흥�|�w�����?_L+��P��?�J8��60w0,^#q�`�����Q��<E�Ago/:ɺUz,'�l�.�&+a��.�:�kvws����� ��&st�����3�>�_{$��z�/���3�e�!�L��j5�73ܺ$�	ݯW������n_��+�؉� Ļ�l�����vq��3�j*Ai�c�z�Y{�.RbѰ�9��j��H�̫E��F�b�~�k�S���	�ٷR�s%;����C�h�y�L���>�e�5N;ռ�����WT�b�|�Fe�� 2�V��_���W��&���7�a޶���}"#:b����g$MJ��{���l���|e��z&�,ݪ^O��_�7'q�L��]
ȩ�Q��ثw��LzC���r���'G,�R���&ud�I�����2���g�f�-�*�O6�8�vj�+F��l�];�}#ͬ!� M��<5�X]�����ݩ��&����9�^l����o"4�O�݂μ�k���`��8|�ʻ�<������T��f:�h���j�VT�_*[S���u�ɿ�䃥P5}�Hj��J:=T���!h�I$��v���t���=6:��^M�m�6��j���`�� ���x���<�yR>��'E�za�~�O?g�EcK�zG:�J_��eľ߅�B:�� �@�Y-�q؃��~<���q���H�w�.���w#U��U�/ER�ц+4�E?a&�!�*�t��eғ��kԎ+V�bYZ$���z�D�_0�ZԹGd*�%p�\U� t�ձ����^�4ZEvA��U)C�sFU)��;Vj!��:�r3�����M��*�ђ^:5J�7HfGv��7�]���������FIўj���)��A��8x���n�yα+a�iPշ�d&a��a�א�"����֖srٚ^V�IE�6zfVv�>�Fq6Wo�N1V[�b�'s�����kǍH&J���Ξ��A
GI�X7�i���T+�ޥ>U)�Eظ����,����V\�����Y�aCy���X	u����DR��|�C����f���-�gcK���	���×2sV�[�*�k�b���,�5HM|�-쑋���4teS�lv.�����N��c��+�.�h�f;�4��X�[�xۼ�i�R�����֖�d��7�Eg)|��2����#����Q���������/��]�t/p��| =��&x�ݤ= ���1����t���R�����ya��wl�i,[x0�"��=�*eAj}Y�Νk�ᬶ��㏤u��1��=J�,����u�\-u�n�Tǜ��wۼ!�=��Z�S�y���|u���B�G'��^����FS�0���N���؄��ChN�Y7:U��{�a��A��\Ujb�Aw��s�V!	T�N^[��	3	�m��W��Ȋ$�+�Fu<�3�$�fY��vj�T5�P��g"��(��ۛTC�I�e�E��֯�z�9{���jlܙ�
�Gc��v�ʭ�Ќ�Rr+S��I���s%�6�]t�21ג�ލ[���[�� �sr�v]T�d�m����u����׫%w^+8gTEF�W(��
�o�Rk.֭�';6]%�&�>�鷛���ug[5�Cg0�/5�Ԓ���k2�Q�Y��l��)�����cc���9���*M�f�Fm�I��������jo^V	[.��������nUJ�����h�����F"��{�U���U��'�`ʜ����%�;�/�<yv\ٖr�CU֝�ӸĤ�f�f���*ø�Vm���1e>:��ئo���ܝ��+�����8�.-Ե@ջ�t�L�`�rw¦�h�5y��E���ɬ������R��-򂸓]�*fΨ��o4���S)��ܙ� �"����!��GU�׺st�z��
��Y"śi[���:�yю�s_+������0��ۮ��q.��KSΆ�-Mj[��U2��v^�7>T꺣=jSW,ކ�Y%^��{��-m�W�N4�3%gNٗ��.����9���D���Z��[�r]��Ut�ʬ��(Ļ�ⓦ�$�#JI:7$�G$�G$ʏ-*5�>��]����)��s�PԱ��l y7;����o�΋�YY�n���������Ǐ����q�q�x��8�nݻq�������$��uvgV]E�Y^[��/s�]��=�x�����q�qǎ8�;v�۷^��9^o��7�k����m��*����.��7j:�Q��Bu��BD��u^�]gVq�;<(��w��|�/.�YrU�s7q�������Tq^�":��
��uy~{{o������w�8=�;�K�&��uh���=Bһ��ըY|��6����xwYݧQ���-Sμ;��q�_3�mtu�ݕ��u�FE�����y������Z6�~k�:/����,�*;m[b�Q�b���ƴi֙gi��!B(AG�,q���K�~���S����-Q�-��g���\��gv���ڃ���1s��5�]�Þ;�&�M:�;)��ܼ�~�>�����_wg���x�@q��0ڏ~s����	T�Jx��N�K�����60����r﷘Y�j3���;��C��t˨�[1�n���ƛ;\�y�Ji߇{���j�=�d�Ab�m�9�M�]t�K���G��������� �5�v��Q](%���k̖���Zg�C�V�U��=����11�3�2cf��~���xHMϿ~�����m���M�鬓t��d�3�=�6@Cz����d��Uv�a�kUounF��~�V?G�/]zM��G���lР������	ͪ�w�g]f��/��\}�`m�����T	I�;F}��.�9�8�":�R��e����z8�r�׾������y���@w����t;*�L�k��i�
4iwo7����.�wI���{O1]e:�v^�y�����2C��}��=���[�n�+��h���Tl�]��yw��VxZ�2�P�W:Ϟ��C%(��kC�D�:�+�7Hq�ߗ.�Y���;Vk�Dݴ���E��n5[5�C���ު}���7�l�U�����������-\�����h���a<!F����U�ҡ��_fw!�q\��^G��J���e������W�
]�tz��9Mw�z�k��Q����j;�ͼ��g��&�2(�Im�*%̌,���w���ټ�-��2rZ(�ƻ���G���JkzL8fj��+�{2�m暂�\�9�J�ѝ]��D�^������Cڴ�c	j+�䚯>ZܧCm������W�f��5�"�7"1[�oG��$o��mҧ���`��s��ѻ� 8b����̖x��[q��}���+��F�U�ٷ<���4n�UU��8�uăg��V �Y��$����i �.�E٭F�r�F�V^��0殬���5�D�=���
7�z�A�b�; ?v�D�J�I�FiY�{k�t��'���*s:�T��dW���;��CB>}��g���������R;}���״��CQ�*u����7)�LO�u����S����v���@�nҾ���  ���-}�k�+�mw`��P++�>S�j9����Y�	e�����it��4BSWL=g"N_Mԫ�}�����[�#EW}d�P�9�ѥ�W!�G7xQ�$R觜�h���=������*C�=�	�ʹ#]&�``o��z��Ё�xz��sp�M�@���L�����\n%�_�(�f'N���TDE9�+��}����������H���$�]�5]!��N���y��ٽ��Mvt��P�xV:�-�Фh���qV���C��n�~z5b�9��2��w�5���G�������|�1@���Sږ��R鄵�ܛ��:���笯G����y5�#�o��i/�H�u�\�u�Dgq���^��>�ɉ��u{�Ϩђz�o;݆��3X�	�Ve��4-_���Y�9 :��H��# o^pU�R���(J(}���Y�yY86��T��˪����s8��dŰz��
H�\�[x�q<�2�X���뚬D�n�zc�*���)�@W�J+��[Ǻ[q`�[���W�:%��z�ᗙ�L:�p'�5��tƝDs��9Ԑ�B��ܼ��K�q��͂Vl��O�#a�:�=9"�;��0[P�b�ŕ��ci���2�M��3Q�.��nW�G�ex�]'X�F��0����a��������[%}�v~����@?S�����g�=L�#��5����f�1�y�/��*wv2��;\�3��+����T��_0��b����K����E�����ckG0LW��"��u���Z��K��1�^|f�7����y�*;Q�-[�-ϞA�v�l����� \zX+�gMog����3���C�dnFi�Qǻ�|����S��1����w_�R[Ig���M-�"6 7%�񘬾����W�n�H�0�� |Z q��eخ�;$k��ݎ�v�s��Z���9��Y������@���a���W�_s��q��AJ��z�9�ݺmԮ���^���Pgl4@�=��³|���C÷���y�F��=��F���{�O�O7X��b��>����҅�)�*��v���M�soo��T���YU'=��!t�Q��myr���us�<V��o��ܤ��e?�z���螲^�D8�lmm�;p�����ɠ_�dA�(��K
y��꣥'�3g@ae��w�V��Lu��lI��S}:�A̛ñdDɋ���[�����K�t]h\�&�GZ�ӫ��F�t��BV��>?��3�M�9��12 O�Cx]��T_��]���� q��#��.Y���I�Nq�����Gs�B�����`�ɫ�B�ys|�{n��Az�OoNNVm��&�P� ��-�+[ꄽ;B��ڋI뺝�n���Y�R0���Z��
��S��Pζl�KD.��UG5����be��\ww6w�z�1�I$�����m�N�=����"ߜb�凷7���1<�oy��I\O�o�k���l�f8S��꺯���f�J��xZ�#zc���쾶��J�J�+e�sǀ�6�n�ɋ{�ݾ�<��xW6���k!ޕٟ�1���/�<"w�x�7�;s�<,���ڨ�y�����[<�3ŵ�Y�ú�.��<gu�{}m��-}��}�Wռs{{���	��h��{)���F���>���oF!�6;E�N?[����d�6�+M����;ns���f(T��N����p���L<��6��a����e�s	bϳw;�(�8U�䱗bL�^��Ş�/���_�aV��X�J�7AZ��Ngb����ҟC'oM���}>���Vp��꽻��yu��;\{����9�/E<������~ǲrq��6wj?���n/��{}[͐z����{g���n_����W����N*]�ܠ���b�k��'�s��<�y���^����R�����]�E��^�hh���qHy�j���F�x�(�~�8q��XK����Ƚ���c+,�E��,% O�Q��F�sG�v�������H��[���ך4��c���u���VI�V�GK?��	5�]�x�>�OZ��f`�][��wj��������խ #q�u>�� +�b�UZ9$�<l�9�v�GG֯/͚v�Ir�Zwǳ'��f�ͽ�uKLvi�f�G������ț�"Sx�rMP|���V�M*�B�ai��t�^�n-��ŷ��a�位�^��@�=���䊰�^�ݬ�c"E��
�w�䵣WQD���tUQ����.'�n%!���S�г��׆�����l^oa����		.�I�9@]
 �@�D��0�lK�:����x�SD[��76F��(��}zSF�_mve������f��2���5S�ʏl����y���n�y0������ٻ��R,�{5k�����Y��p(� Js�����U?Ӹ�&b!t�#b�)�ѷ<��D�&8�l���鍺�ڎ����췱�4��p]0���/iɫ��8o#7v�;Е�5仧�K�Pϸ�m��}[�Ww6k�����w�;|`�d׫�Ǐ*���4��7���`C�׹�4����ʇ`����"���3�&�	��~� ��'�Q�o����5��^��=�=>>!3�������7�?}�h��#���Z��Y����)���TcC8�z�_P�T
����=z��	g���u����'��ح̍�@�Τ������֕j�lo_�x�/L/7R4G�㢣^_�_2�l�0��I��lj������^�>�Wn.�^ks��Ҭ��ɦ���S�ܫ�D����Bg�����j�񻿨�(K�ǨWZ�l>��L���=������걲�ɓ���2zN��"<����
��ysJ�e��*9-�+*P��u�=���rs��7/���:(�u�2��K��?|~����LJ~~��0�ϵ:�0vO�W�ѣ$���Y�\Ӝ��CC�m�S���39^Ð<|ov���RV�.�#i٭���,3\�[f֮��p�OQF[:pɹL+"+VϥƸ�_�zQ7��x;�;#x�L��gV�_w���������@�^Fb�\Dz���cGe����\�oF��EqRXh������pj��Ck&f�qj�TžY�O�����}�\Q՞��7J�,�w_!�h��	��e�T��ӻ����3�F���qlgb@�t�^r{�^5=�F��Sp�Im�U_nFv@ra]�1Y�Twl��j��#T�Y}N�]&y��YK�Dz�Z����Lc]�Ƙ5O��yQ!p|Ξ`t��'zH���̬q4�[�׽��f�鋙�P�F�Ar8�O�`!�T���?�~��e��H������&�GE^;���f��4p)�?Y]�7Tv~N�VSe�+%���;~ĳ�����f��l��l�\JbO���j7.��*�[��e;�X���ƒ��G\u7���7���D�����z����N��?C�w���9@������ͣ�HF����[��;2����s�ߥv�e�:	d��O����0g ��>9�Rӻ��$�4h�Z�Z�= X��yu��k��Ɔ㩁ً�U��ܭ�*����_��{�	�u�Њ�5mU<���H�DH<��5o��٦�<�ޜ�6�?��U�,���KhɆv��9���r�����J�-��]Į�3�~~�E+�5<����z
�p#�&U�V�Q
���{@Ӫ�'zwF�[=�j�{2ni��AU��,���v�j��[t�ѽS�;��i�vT	��$eW����N��� �Ns׍&�4M�>�v+�8v�m��3�*t�+���F����PI,��vGe:��m㲫"3]_%����
��A�'5�qh �\��q�6�|O.�p��)�5Wn�dUz����M����&Fm���xw<ZP�9s(n�ͨ�'v���]T����8iv�ܶ�p�{oy�R�&�jN����=oq�w�tw��
�mod�v����	G���8��ej��8ͱ��}͹�Y��/7�ߪ�S�#��S�wW�öb}�m��&���4M �[-w���F�~'Omw]m�WJ�P)�d�����g�Ѳ+T���W���Mn�^a;ϫqS^��뻌�[܅��YQ��R εSkb�Q|"�7ON#���$�O���M�J
���u���Ia0�Q���#�sτ�V�>�z؂6L�jږ�=���wx�h
O�}@���1�`/Ϗ����w�e}�Ey�M��2�mb:�]�#E�7-0���0�Ώ�Y���Z���ι�p��1�\�|��!�`��<�7gͦ��<�4�v3��c{��^���k�ƌ�x*^k�r�S��]�w�эS�9�l����c�V�gE��B�xB���F�וAc�=&a��EJ�����ݥ;�}��"Oo���uמ�}�5��=�W�������~+����( 
����z�����(*��� hu���D�RH!1VP �X0@�`� ��P�`�X0 �`�B  ��`� �U�1 �0@�0P�! 1 �1V �  �BP �X!`� �U�`�@ �X0VAE�`�  �X0 �1VU� �0 �`�1@�1V@ �@@ �  �X1VU�0 �!`�U�`�BU�0 �1 �@� 0@�1V�0@�0 ﮇ[���+*���A��b��A��A�*��� A�t�Z1VD �X1 ��`� A��A��b� `�*��(`� A��`�`*��� A��`� `!b� A��+(b�
���b�*���A+*���`�b�"b"�(bb,(A��`�(`�"��!��T������	�+X�"�
 @b  @` @b���A� "��d(������
j5 0Q@ ��  0@BP �1 B �P �0@B 0Z�:DX2`1U���0 �V�X2 `�0�$0���b!�$
��@b!��A��
�ZЁ�n�`��� @b�*�`����5V  �X1VU�1V�`�_�;���p)����*�,b���������_��?���s�O�!����_��_���������%�����w�O���}��@ q�������@Qz8� U���?�@��I�E�����?rڀ *���~���?�Ӥ�~ܞ���������t��xEDQFU"� �$��� $�� �2
 B UR]UE]T��UN��b�DZ�D �E@ �� �D ��@	  � �@�E   ) "� �� �0@ �T � `U�P !`$U�0 �V(�#`� ��U�AYҪS��:�J�J���8Ez?hBQ�����O�DDdAI @$ �Q~�������w�	���`�����( 
�?}���o��o��o�~�$? 7�ЇG�q:>�� p>�?D��:���( *�@ ���������f�P^�����"� ��@*~֔?�k����<v(�_�I��;,~;
@�B ����O���_ǭ� 
��vb~�������?�7��?P>�'��p0�o�A W~e!����@ U���������Wӯ�4~@JO��������'�B �I܁���J��`}�@��Ë񩞯�E��l
O[@Ql���������?�1AY&SY殛HY�pP��3'� bB^|���1[9�T��)!l[%P�PJ*�ѷWeTQ%$�nEu�(U"D�JM�mR&�U��a�v�$�vb�-��Ռ�K�4��wwv��ק�m����:�����v��i�����WNm�V���m�qݮ�;���;����ַw+n]�h�Fv�]\�t�n�E���w:�mk����4�����s;a���.s��vvۧUݕ�S��s�g-�ݛ��k���WsL�Wn�����Nn�;kSv][����u���ַbݜ�㝻�\m�n�wvΛR-�m�L�u��ݮ;q����M�]���  �}m�}�d���ڴ�����=�F��L�k��]�h�۳���릵���ފzh�Wz�k�n��	����۔wuƺ���{��ö���ݽ�n�:t�F��նvۮ:�'-��*��[�  ���H�#l�q���ˎ��$H�v��i�
7�5�y5�*�ؑ"����҃T۷_w��Pgv�V��u���JӮҮ�Cv�9�S�av�Zwp�ct�ib��nV����*��^�ղ���V��n��ѝ�]Λ�_   l�����ul��s�`����;t;�-�{{ t=tݑ��v������T׶�9����:^�7Kחn㠫v���J�'{g5�C�;w��ӝ��ً�:�:��-n���վ  �Ϗ�(���N�V�ռ��^��^7{Ƥ���k��==hk���ֆ�U�p�ڇN���\�	ں��n���uڜ[kGM;ݶ�5ҹ�b]�ӻ���nW\��|   ���ﶁ^���V��������´4�;�]�w���ۺ {���[�� ^�{q����xأ[uһzn����th��uծ+vӮ���k�6���   ���Hu�����^�U��]^�V���=kӈ/v�8�T�sv(ݺ:�Fw@ su�J�*��
�����v��l�7J��ps*i��3kT�]�   ��z@=�  ޺��h@��c� �g��  y��  n緅 =�w��� n�� � ��<z  {�m�:��-����ʼ[;e��  �|� ��� Ok��Z �^� B����  �On  �S�� t0 -�  ޳� /v�=�qn�\�;n�n�ۮ�5�վ  x��(zo�� � q��^� �  ;3��� 
;;{�  yۼ�=  9�0 tmz� �;�=ʷ�Z��v]�6W��s����  ��� ��\� �;��i���:  =��o@��G�  �׀( x�w ��Xh �� ���"��JT�� ѐE? �)*��h�B)�14��@  S����M@F���'��D��  OT�D�UP  6S�����_�?���?����?YC��ϼ���bdx�K��3���IM�A�����}��cu~���ֵ��Z���_��Zֶ��[Zֶ�����m�����߿�����������M,���#��x{r�-n�ܰ�N�$��t�8���i}��}�D�%�AK��-�۸�ay)' ��֍�� E��ĥ	���d3ǎ�gN�x��'{�TV*!͡��EQ[$��Ӗ^�"I���Zd2!+2��-Q1����k7�N�[��-�twBӻ*Z��Yݱ2�B��N�V����@;���V�d�b�f�
�4#BbH_����jd ZN��݉96��p��J�\2�� ~"�Q�)HE�Ӱ�係��;Zi+�
9�(]
2�SCe1�-��@�Ԥ����-ɐ^��
�P�d�V�V�/n��,�Lm�gY�:,1��9���K`�N������+M�p������)��Hj��]'[>�Z>
�ص�H����������G��!������)t�jz@�uY	M��P���*C�z�#e-֕+͌��ŵ@\�(<v���֧�q�[�(��P��F�	1��ɠ����|����Ř��
��oL*Z�fbt����mLeLQ�J�^�[�e<ٮ���XŴf]`j��oFL ��0e4��B���H�u��2ۼˡϖ�'Y��R���3�ib{�e��5������#rj�I�F�CO�A��L��v� ��{[#�jڳu��H��o�)�A�Պ�R�+u�O>!o;F[����S����m*3(���� ,�ƴ�Ҍ�)�C���Q����d%��d���tV,e[pP��� �۔d�4��ͦA�H4휧@^���t�v^e� 4qc�����EůR/jb�F2�D��if,����ہ2�RF�c��"텂���#SC16Me�M�ŏ*l�]�����1a�67�{MG6�#&n�aS�b�)m�QM Zq$FV�1�5�`�
���]YZ$L���Ϯ��P�͠��Mh�7��̇Aɶ�e�U�BX�	�1�&u�X��aR�=�g�R��;�A�Q7���^���^���:Y"Z��`��L��e�Z�)�A��<�i��a��1;7���qU�K	Yl�
1ٴm�v��D雒۷��&�e�N`3PSl��1�溣���ywn��Q-�^�@���d,!jN%@�y���u�����യP#���E�Tn�h��@��x5h�sh3TM\��EC�-ttjv]�0]��ժ�Ȏ�W��Y�qZ�t��k$
�a�4` 9��M���n�x��co�ҩq;�d�]� *�	�B9,-B�MR��ẽC�p�+D��c;`]1������1;����=	kztI��c�wb�n��XV��B��W��h5s,����Ҍŕiȕ-��2e�����Խ��1J\�K��̤怅�Ƴ���ެ!���K,n��8�A6iرV��A�,n^��nA����ٖ�@�%ۧ-m�giT�35��+]�&��5$�2��R��OE��(ri��V�
���/J��LP��^��]aS8/x�OեV N�gRZj�ǖŘ�,ͽj�/�e���(|��麎X�@6��0&��5�x����@aČ�M,�uF J�Y4ix�}�o�,+��ӯp�@������j��0�ͤ����`���e�Z)��m��Q+��9�~gB+"#z)L���x�X�ډ��cQ"'I8���υ�Kq���e&�K4F-��x҂mһ��W /Z%��R�ДҤ���1JTKo�֝�̛CNPQe��KCTX��ZکF*]8/(S+V�̓%H)d��z*���'[{J��(�k	DIt�Xq����`:j�\ѳ��E��Vnν8c2��b�e&�ʺ�%�EK���ZKx���3J��@�vs`�CP�iL��T2ŧ�a[Aə	݄�3lE;�u]7{%���۲d�w��@�-_�5���]�sEݑMn-�T�mXXZ�"�y�,.-��C�����^��77u<� c�nj��;Y�q��iՊ=|<�͓�NaƏ)�P����F�)fN[���k;j%�������V@:��W��W�ީPȔr=�kkX�.��@�(��� S��4>��C��Ձn�E�E�� �dl7J�f�Vi��Fh%[ƱԤ�o����f��L�GC-b���m]wvp�7�AG�X�IU��ɱ䀽CcSSq��kܼ��(7YH��{�P��T�$(��j��ctH�Q9(�`�	Č1���~A L@��i�	KW&�N�㶝&I
[�i4�R��)��uUe̡ ��D^��˨�)������̎Ԁ�Y 
h�[�݉��p�WX�a�F�E]�!�ovB�d�q0(�-�)��S sj�u��^JаjJ��pG`/��+s,�43�} p�4I	��2��N�Hi�5�����}�t�Y�w��U�	u�c�m���y���YZ��oٔ�v��&�A^��M[����2)"Q���r�n����*lYu��Zk.�kw/tf�7Q�QՕy�E+���A.�bu�� 0,E  �9�9o�5��xϡ�Gs���������Y6�M,��Z��,h׸�2�`ء����������}�Uc׋E�f�4-Z)�v B�]�Q-ro��Wƕe����l�N󚤙�K���-���ȵ���n�����Q��J��{�Ո�)7�{)�u�F��h�	��B��4h��2�XfI�֙��#�-�t��m!JVK@�56�%V@6�ssVk�l[
�C����q�I���^閂���M�Ź�����Wb��$�6��nLTkNө����-i�����f�-e��T�U,��n�>�tq	�Dk7Wh�)�X��u#H��Z�1EIS�6��t(lz�Pp��H]��m�6c��%J�E�ػ7��م\zRV!�����h�e�����P�6B�ۖ�2�
�om�!����m���k%�ڸ6�)��'�-��/]+�I���d�ČVL�o*�f�j�#p�t*�� ��[�InRDlZ�(t��{�5����B�(n+�Hǹa�f��^��V�fZi�������5��xZ��eat��їE�@����=I�EY��&����x�1PY`cIZ^�B�2���e��(GyA�Ճ�
�o#l2͍t�K��K[hv�ۅ�nU��&�/Yi�5�'�AT36��i�E� A1�p����}���Ú�~3*�H��ѵ��ڙ��b��3*:�cfఝ���Z�JϞ874�n�xdN���<$*y��Ƅ0�N�iS��k+��ޮt@
�W`��J��`c~��e=6N1J�)Xw[�L@Ӷ��)�D|����\Fjtn�b+i���;�Uc��
�,�N��A�Rl�'6�v�"�-�G,P+����*�M�j�z��L���$��R���� ˩�s%�Sݡ��m7��;��2p�{��C�"���=;�qj�/FRy�f����V��Ss����!��#���ѭ�q)z�ލ��Q8�������X�RbdP�n�ݡI�w,�R���Ӓ���3�,���e�4
��S�6�u{�CVŵ���h[Cb�tż_]�b������L��A�د��$�wO�]%���[����a�6���mީ���xf�p(�
��-�QIE�eS5�򱷺km�n	RƤ�K��#y�`�(ƛ�ӂ�a[�Kh($ 6�]�{����B�Zͺ��A]8�ء�ݼ��F@�mm��
rX�WZ��z�!FB��//S�	.<��mn7X��z�� �:7B�0��^DMǣE���H�����m R�Ul�2��0���ڤFi�֞%��j�M��M���ڹ��5� �v��qgm�PJ���
-J��(Fzʨum�2���4�������i� �)4,Ipҡn<d^mm��:���>ޭ!^����/J�7G\�.�Ԋ�|�@��8��-j�����	1��E�hJ&��h��C*Q����� ض�2�Cou �Ք������LY����ͧgE�
�,�h���I�)b��M�D���$օ�E*V��{��
DUn$c�ŕ�Yb���v�ha���z�PWB���
f�C��9�Z�����ư8mX��ot'2,����Pp�8�t3�P��;J���S�7p^\@��譆�ܷ[c��n�ce��-�		����TR�P�吥[ZrFE7���(�Y���p��m�Ӵ�Z���%�h��P�i�N���i��82�jFd*bܹ�ՁX8�gu�bS�h2�!U&勛�A0+)�R�bF��:�n�r
Z1S���"�/�Tܠ��`��PV7v�B���-�4�������oA��m�q#�]V��zKBd۷���Vh*��sSS=ڗ���c�>���'I��
:6���Lj�͇�O�+t�4T�c{��ǳ3JC�~҆<jg��F����~�M
b����Z�ln�i�$�,V�q�&S�0Ƽ��v��I�A�i*��Yn��*�Z�'b���`���ͻ[5nh�)�v��I	zU[!(72�܊;Y��!P��B�b�3IAB�)Q�͏u����t��x�E��uu76�$����u��?�-������h����x��
�č�M�#i��L�&��oHҨ�jquϘ��c8�P���o�Ո7f�=vl3j�j��'�,�{.D; E�x���DN�ɸTKv�E�Q,x��KV��kbE��
��YJ��U��X/j[G,]M� zBf�.c�	�GiʚN�-�hՓ+S�@������+
���>_R��3]�*��ݺuw���g!ݵX/f�U�94A)�T�4�gX��hb$#�w�mR�[�0�E�^
��k*�MB��W��-���VM�B�ʽ����W�5,����G�U���,pT�G*¨����C^�TӼ`I6M5�/V�10�c���
��+�=�G�*��f�ڔ#S.ۀ�)B~Gn��XC���+ח�y8�d��"� $3I�6u4*����Һܡ�l�YOIMR���J
�%=�y��i�5gj��+Hg(�	}��"��� �V%bۗAE�T�6(�,ҙ�ych����0I����ݸ	�G�w)�U���=��=�����DOqg,q�I�G�cXn��/m�.�	��)�yY�J����f�s�X^�˨���W�eB��.��&���Q�f�P�*�z�c?B�kb��̙l�b����ӫ�����'��щ��,I�# l��Cc6�������8���b:֊V��2iUqn.�<����o��&M��O�L�3n�T�[-�#9�������Z�N��eb�X�өH�V�+��7V`���m��`-{�y]���Zt�Z�f�*�h�c�5H�d
E��M٭��w�iY���6�)A�;W���93K"�*�Z�سSM�:��P�D%�ҍ�V&��f�VF�0$;%n�4\�@�v��t2���vCU%�4�in�stP���d,;:�nbDQ+)6�����0��#qenFk1��s,E��B��ݙ�������W��>�����i$��J7hR���+HO6TJ��J�]l��.ܵ�"�JZ�۲5#��nh��Q��>m��%2jc4�ۊ��V��/v�1�)A������\Wt�+̧*��g2�<�� �+Q���gҶ�Gd�hT�,���hT��"E)�)n�V^%�T
U�KZЕ�[Of�Ӣ�fDa�Z�4�M! ��x��S�.���j¦!��>�#��$� �.{2�ض��P����S�Aj�t�M�dZ��Mk��F��-��[{21�H�֐WA��*]ԱQ��G/-�Co�Ân�M,�� 7/���xS�<m��$C�7s%��2΍m��m�KF��YR�g+FTDڌZ3K��Աpr�&͙�j��)��ۂ85jv�c(<�(ff�A���2��ջ��_� wXl���sXE�R���L'J�'j�hW���)Eƅ^B�)�n@++%�a۶M�͔�bQl��iYf�ߊZw[��I�r��Z^ImH�싒��MJ�*�dn��s�W��+2woD:*���&�0$3���&(��`YذwL@��ѭ��I�l���GUay� =	���c~�ýѢ���;Ԓ1�Iђ���"f��|N����_��#�G�5���[F^E�k �ꥣY	X* d]�.щf(	FC�Yd醯��\Nh�Q�Z[�H#Q2��[�l@��P���mLۨC��ۤ�43��6r� 1�Y�(�B��´��Yf�a(-�X�E��@A��	�$��e��wi�Z)h��:�¶�G���W��HȸvE�sYSV1Iˈ���yL��X��.g/sc��v[#i#W�;�0�2�$�b�AZ2�Ua5Ql�1GQ�Ǯ\�r�ϥ -�h���T��=0����3_w� >�Ht��fm��:�ue�*�e�0�R��30��!a{F��ɿϦ8V�3��J�gC�w&�(^Ҡ�Z����,�P�s`�D®��ᤙYG*��R��H�/��ڀhT�s/>�J��n���Y�`�n5���W�.31���t�3t�$q��ٚ6j�9Z�m�(&�ʇV��]��ԧiY�Y��z줱Z̳"�KF+ڸ
ò�Q+1#svV�-IAK�l�v��̈́I2�s1S:ñMB�[i�
Va`�4�o�P��*șz�Ŕ�(f��n񝆶�kDĪݬ�(՗u�0H�{j(�+��jk� �����9,'�7��I��ڈ�u�^B��T���σ����}�a��]ts�`s��Ǯ�E^HudB�pq^\�A��30�ueɼ���撗 իw�6��x�[����T[.��ι���6[o�H9��*s���R]�{n����][����Plz3Ԛ��]��:FM��S(�2����:V.J3]Wx7d��u#[Y���v�).P�O�X��8k����㻺\ƚ]�nBGIZ�x�(>f�����ñ�7��ci�w�X�2�[f�F♺[��j�4v���v�˸hf�]j����H���rSW1���*�Ƀ��q���܃pr���\��:���|�t��o����eh��:��ޛ����jt��u�p��8z��v��I�b����;{�lQ��۩�Ө"%�]�0v�`�:)%�R�����f7պk6�*�lK��ki���w(�;����
��3��v)�@�V�S����7�t��`J=��&�֧b�x���lY��9�wK6�B|wh�=�i�
G31��צ�%:�?M��+I��u����n@��e�u�!}�^c��>ݻ�a���o07t�pA�t��.l�������H�ԁ�����î�]yw�U��66`B�F��g��88�J��*�\�JQ�٭Wa��lԹ�D����.��1��O:�pW����zx���R`�5�N��K�OT.������Їb��h�Gb�)�<���o)����ʗ0V��A��+���4�!���1C$��7x���^�"L~Ó�yUsQ_�7��1�-99�uz���r�-�`mrr̾�#&P�-�;�Y�Go���V���Bh���˝_t+z�x�g]+����d[y�=X3��ё<��"�b3z��ىj
Ѯ��Mu� ��޹�,�f���u��AW���do�o�Ѫ*<�i;�e[E�֜���HE��}��k5Ӱ�o�M��L�F�u�7�R�'u&�FV[;B��c�[kBAvm�����ޒ����6�V*&;����U�U��#���k��[�i��C8Fgh�J�sx;;|��"�w��ެC�)���q}E\�x2vvىv��h����]Z޷3 ;�a�q�ʮܗ��MM���Q�.�����2�M�W���kL�w�1��/�Z�3��Sd�ʙ��P�B��,�>p�5���Te
�R��TS���T�q<����3��+y�Uu��\�I�7	�"J����8�}4���*��^g���c��Io���|�ܳ��o���߮�����8Ȗl�j]r��4�"�v���c���N��3�U��9�-�1?��m�@�X��.�N��.�uޛ'5��vv�7��..��rqQ������]ԩ�̣�f	�Z�Y�y3O��M����ࠖC��[�9
�i��`{�$��9�>&Ņ�r�4(���&W.���K�k�ժF�il�O��X���w�;C"���w'��U�$�I��@+%�	Lob�Z���Dk����VE����������&b����hٻ���E�Cw(�+:���Tg�r��M�V�h����7N]\a�[�Y:�9=�T��y=��0ﮉ����'Mt�su�.��������1�a����K���c�(�y�[�\<0cs~�Z���-+�Ԝc�I�j��p���İ�<�Nżr��nv����YG2����4Z����n{o�]����֥�Y*F�xd����ʽ��`�}䥴��'t(r��.#:e�lR�2ت�N���_EG��8���Jޖ	��b�)STlo٢��Ovr7(*�Ĵ�+FT&�c�9�W#�-㶔S%�X�Oa��U�]r��r�ٔ����]��Z���(�໐O�7��[�j��мD������]��f�Q�=���G��y�Gm��7�GV;wΗRR:5;�`����ݠ������ڢ���W'#@ՙL�S�&��{(�R�u<Ͳ������X���yןx�Н����G���٘�n5�L]�˦�xA`n���]M�҈���r�N�xhaJ��]J���`�H/M<a��C,�j���>�̱r�[�X��V+A�k�Ӄv,��7�H*p;mg�:8�%���{��ν{ҋb�.��)��+���⭵�z�!+d��(�����K�{���Q[N�x[n�!�G=;\;eAVӫ�K�ȏf;%�;{)�,C��AcCh#{�\w��5�v�L6hp�;��
[�]-�b
Gc�?nȝi[+6��V`=j�Wx�Xj;����۬��cf��wg �#�+r����<�i,w����_N�[��*��,n0�l!����(I7�q	�+`��2�7
�)�G�zѕ��6�ǯ;�`��2N���\�[tE�Q\���W
�\Hry��d�v-�0-v��yQAE�����ǂ�p]�KAʶ�DY;��v�2�]���J���Z^�]������AZ���)(P[u�.�k�K�f��)u^X�Y�HJ��U����P�8���4T�O)�RX� �36�7n�nn�������w�v҂�.�aU��gUs��9@��O.��Pz��r�pq��#X���u����^�osPz�9����k�".�1�D\�x�Z��!��jw�F�
���<�S��O!���4XZe �RՅ�g�p])@y>(£ܐ2w�&��x���f��vT���]��`n#�v��Lx�.aB�%2`ͫu��E�]����G��j�Mţ[Yc��绦D�vo[�n��_'Rhvn+�:m���0�e�1N���5y��v�՜�Z��ʮe,�
�iER!�~-՚:Mm����}3�>�3lMι��2<���u��h�'�ԥ�(����M��X��z��>�,+���Q�LUް�se�j��,��(��}L�B�٫�	뷣*�%
����b3m�&��SK8c.�� ���Ea!�^�b�4����>���@���w[ܓ�B��br�]�a�\A�]�[�
����z���̐Mu��:C�ö1��`���xu]_�ү�G�qB��^M28�T_�Ŗ:�NVz�1��X����mB8�>�"�u����o8�m춊շF��b��I�Q����h�D��Kݮ���H�/5}�d��pq�S�D��"~��'�y-���>�{���W�Gz���ΰp�!�/H=V��﷢�čS�%eՉ��x:�Ɋr��n���#��eE��D��}�*:\�Li�k���$�]]L�����b�4Њ�W�G)RFLQ��ƌu�"��n�1�#����N�;S5�x���<�D��E}2�|p�JPp$j-q�{���c�+=����>�th�Y�����o%`	�w�s5��&g,�8�R�Qr�	L���bi{1=�[�N����gU�thh�嚱Ү%FK� 'B^�NR��-�;Ʉh����n�mQ���k��G��옦��r��n$�'Ǔ��W����۾z�H�4�]�ñ��ϴ���/f�s�!�$C���=�;Ҭ���3@���ާ�F
�/Uqī��1ܐp���{�E�hD��5��^�1
�sj4�&^�r�����.�4*�GL�N�{x�Ih���YoUl����̥Q�n�|����+�f�Ft8�3�/����:;K|)��t�* Hc���Ӽ&��Ymn�{P���
�x�k�5#��'^Ia���rΔ/�nL�8w5pߍ��{ѢyA���ɵ���uȨ�}��@� S4���w6Me*z�\�F=wInd��՝Zp����n'�,ϓ�mv���³���͒=4���t�)�R�b� �B����4Q�:[Y��.�lg�휊�����c�J���8Fk�Q�=�{��g�C�W,�--��-V�i���/�����o�y�}�W��O�s��8bяnC΄���Qpڴ� ��f����7�i��!&�;z�mh'(����p�2�{{^��)I'F���p޸�9�Q��m�t��ܾp��v�4�L�Y����w��|�y�V�k��<�=�3��t��K:�g���t�Xq��,bǳ�	Ǚ�_+��0�3�۾�懷۠x���BY�ڵ_�`��-v��S%^�&��!<q�6����^T��b�B��+���������n̩9�[J�7|!��Z6��cW�#�f׸���n�Ӄ�H�\5ʽ��̈h�a}�.b	���Y�۶r>W ����j��y
�r�C�4cFJD��S����6�d�\��pt�qp[�#.��ڨ�`t���s���}�4u�P�n��'��2�oRg2�ڈ��*�
T�71����p�ɺ	��(cU2Z�ǚ�)�2v)�.���%>�Z�싱�SVK��-ی��7���u�	 cG�u޳:P=�!�lc�Aq�[J��_n�8�V�ic�:�8A&q�
)0�>�34�U$uY�M�v��6�4Oi3y�c��7V�kfr�{k3�ӧ��.�|�]i���/����V���0�my�ĳc)���va��LǛ��$n�
v�
5/�E��`��dѕo+�X�/p�hYNod��r�4ᄭ��w�JmC^>w!]����y�7�z���^���:�>p�5�srg.�B�i���L�W�ݻ:�ӌ�Q�c~�������Z�L0����$�IA&3�G���xF������@:
�W���6򲑼$z�E�Z�>�~��j�ӯ���7���c�J��S%ބ�>�n�����<�;n.�<�p���O(	8I��[/L	�����ou�6���$��y�A�;�;+�f�9uaK�w:Hc���̃3:�ݸ.�X���q��❚⥽T���d{xXt�ëqfG�HuG�����R7]��	�����V��
��o��K#�MO��5z�F�W�G,�/w�kGiG_s|���T�m{&נ�v�r���IS�
wLՌ޺.����6$S�&�+�u���o!��3f��uRd�h�6"I�%���+b��&�!�#@�u�QXP�ϲn���%��9�Yo���;�և\t:�l�o:b�x��4bE�7U7�n�S�*;~�
7����b��Q/����w>a%8+37^���)\t��]�z3��![�&��3��zb2¡�q��D����Gz,Wlˎ
z�A~௧h������!L��k;% )R���Vjb]��6�E��bb�˼�2�r��U�Â[4��Ջ���B獓�{/9D���q�ӁM�2�c��R�^sdŽ�i�Z���B�����{�j��r���]����������`�w�ͬ��Vj8�Ҷ�ߩ�WN������&6wK� Du.�'�8��i^���T>@SO�u��8�N�L��j;�CWv�����J������x�:r͗�c��o���i�X0|�Ǳ̳Fϑ�M�ո�L�e������neq[��h�"�i�|�7%v@��.]6�����aJ����9e亹y�(�Tu�����P:��.���7@�*5m�/�ff�7&�[ʂ�t�v�ÑTy2p���ykT���v+�Dҟwmf���Gc�~��M���21�E��{ L��Z��m�
=�8�u�k�e	����)N�Pm>��V�ӻ+����2\�
p�M�H
�B�B���]�C7��(QF�k"�w��+Jy�0��s�nmػ���I-��\���a�����gwns�ע�t�Y	&�@T��q�g��`V�8D*�b:/8��M�������x�����_oJ4�iG�1��]HyNmZ~7�&oQ.��pt� ЎG�)�����_����9t��o�S�{�}�} ��A����4��f�U��aqɇn�Y�N�wi,��57�m�ً��y��o&�5໙��s�s�}Q�o����|���J���N�`!s�-9�U�3���Ѳ��5f��֧F�dP�V���R�g6�ة9x�̩��e��^1O�:/4���������|b=�8��㬺4<s�_jr�4�j6f��{�#E�a��uh\Y]N�����˫�}2��Np]��皗02�7
�Eejҵ\�L�.�����<Y2u)Gb��+�%u��[�[x���H�\�R���A��!�Dנ��v�����>�[E��z,���R�}vt�A��%*�݉R�\���櫵�������l�K4)��G<�s���a#b�P����iN�%��Z2�.r&�_ʞ�\<�ṽx������;DZ�V\&�����Yy��L���u��x(��i��]���	=��z�U�RJ\��Y Qw$��:w�7��Pb�C�f���{�^ZH:�M�ĳ�aI*V�l��燳�U0�-�3S\�O*D�3�K�vQ��o��w$�+[q^�r��q�r��ٷ�z�d���@�1�z\�%K�8qh�[��읦^�V4���2�����i�7/T���.g_���9�lެR�N賁���p����p&�c�ðšVɹ�c���l�v�u+��4�V�q���4(��Yѽ��G;O��9iI�㋺�퐶y��v��s���]e�7i
ĳv
t�R
(��R�܊����F;B��*����U�Sd7`5{� ^�)61}����	�z��Ж��,8�1x��I��C�b޵Ym�A�Y��9*�������0�D��eV+w����:��A�3�Ps\�T�$�]�g���SN��})ѕ�z>�>��b^��H�^sk��c��}q��m�)K��ҵ��Uf'B���T�]W6��r�
����1�n�r=�"6�p�tNNlnI��j�f�Ǵ ��o�j���/n�w2'�2��̒�58f,�sr'"T� ���$��I=�S��W���UUDDG�}�>�>�����ј`᪓S����W@h�\��Ϥ���2��F��Miƈ	*Y�8�w�*�"���V���mýM�E؃s�r�P7�'\Ӣ+�v���_L�5�!�a|2����N�����'ZE�5{���4�K�U��Y�9]ä�y�l�t{�:�������oEBE�N����*��4��i�m�����IuNo�U{�g�1j�gX�sI�)]��Ih��F��-"��.\q����H-��.�oX�ȅ2,żöZG_)� $��y����+A�3w;��4�;�*T�uKń9]�i�w��-'�fo[��JYi��y�0��f#���8C�w<�A=�����͛uBMW�/e�w"o��XK��)�ē�j��U2�E8��i�}&4���R��dє��wG��t1��(�^��k����ff)w�q�7Pl�G�/:>NfD���Q�J��P�eGS���+&8!Ԁ�����\�\��sZ�0�V�뾚F>'9ͷٳ�>�;��ٰBs����2�U�J�YP`����w��e[QXl��m�f�����3R��5�5�.+fngh����&�����V��ְ!�;�m����9�N�v�V�z�'�ժ�R�C��mqًX�c�z�ʷ�i)I�ͤ��E�
����K��V�AY�r�ȉ�V��,Ǆc��ne��i��t �Yg�Lzk�j̵(�`!��=Qf��
S`�+0�����y��^���^�Ǹ�����铺��];ݙa�Oq�i��Y�9�|*<����N�@q�l�W[�.�{`W[�ɷ�\�<7�&�˵�'2ؚ�35�sꀖ�]jr���"bv��O��ǯ] +;��Ŧu���$��`mū܂9��%�	֪�����r�s��b1�O-@�ޫu��[1C���_cv]Zv&E�G�� ���'q[�eH���t%UEj���䕑c�[V1��Ы�1�=4��4�9k�>!��j��sQ��h��Y)VY�֣��n������,b]/ֽJ�f3�ylSq���B{3O?�B�ʆ؜*@Aˍ�%o���{�)��\98sʲv�φ]��dƏ"�@�]���am���̉k�r��1D/_4]�	W�z�Q]s���+�}B���sx�x)�Y^����n�$M���R+>�rJH9d��ve4�XD;(������C\��H-F��N12twia1����WS��e
#�9�F��]�sl�!0PѮ�I6S�4��.�:����΍֗�Ƹ�]�V�X���7��Q-��n�;.%y�j��i^=�țy����`̮$�b9���b�8��R���g�Q�%��Qm,��n�V�г��Y�e��wh�P&�^m��jl-f��V8ޕ�%m�6�x"ޮj�=V�T�2q�����&�Si����ƯJ<C�3��{:�trq��ibaU���i���y�R`�k�0f�����8�sn^��^X���\O�+�M��NXy�Va�5�Jr]%![h5�E�ׂ�@.��.9IΖQ�1�q�Y)fFrs�\����3j:-6Y��g;�I(suRʾ>�;�2o2��D��(V�Ks�9�bk�kp���/:w�y�]���嚊<g5���՝���ڼ/0�>.Z"0An���]#$��V����b\���s�*ԕ��Y3�� [��l]ڳ���99�U)sc��rj�/f(�;J��Y)�#�G�t�v���=�5�ogK���5�Y�p��NO��5���h	��T�8�����#�w�h��o.�n�nt��eĐ�j#6��yI�9.Z'2ʉk���:�C��C'��P�Cv��4�$�� ��U��!�:f�i��lN',-�acÌf�Vx i�b�TC�]'�]R�EuKIVc*�ac,i̽
�q�fIX�^�$[�f�'�fF�K�"T�B
de$�o=��#�ZRwJv؈�`�A�7w�%e;� ����
\ѕxC�Wh,6���ZΡ*"�3nd�����h��1k�T�$J�����dr���f�qv|�`Y]5sLW������,OG>�B�-d�{�Ĭ���B<�{qXѓ�>��vU,�����)����p��]����C[X�GgX����J�b4r�N�6����i������k���`��1����ئ���xmYw�����ҹ�a��E��2�8��; �d��/]���p+۵2�c���Т�E)M���z�sknCw�x5��>�`oQ��� �=}��wD��\9�.1mw.�\qR��ܙ�4�O��"�o1�o��7���%���aK��zv��w�>�ò���!�0*�݊�����p�T%���kU��Ι��Y�x�Zg����9���Yx��o�7��*c����5��3NOY>pu$�RkX�n�,뭲K9U5u�rq��v�*Z΂�t��Ty���qWV!#oj�W�L(�#fu^!wV�Wu9��`,�r��-p�%�+��_@��{�����N�$d�ϲ�=�xg-�l��5kr.qZ�9wD�@�թ�f%�R����!���y��>�p^8�n�j+�������B�a��^�qZ��[t�r�MV%!�Jrbl3z��5�M�MD(�O�����=f�8B������XMr�F0险s�[}��]n=�˺}q�7���j�Gt!hfu��vS�Y:݌U�
a�h��_Lt�V.�8n����y������'sFM*;M�Ei�l��c1u1p��Z��ls �4�޵e�ٹ3G�V%F�#���s0j���7�A��a�{��%T̴�?O9��dncN,gѩ^�em}p�˾�W�,E��]M��]�'wu!�7��r�.���e]�[*5�/C����ۤ$9Z�6�ɘmr5�i���D*�#�k�m�)F`RZ����e;Hu5Ѡ1t�͚����9�#�N��;
���$X�v9򆢔��],����(�������C�g%��4�&�(n���l>:�Y�VU(7�Y����zo�3��68��HT(����eZ��br�+\��¬���11yȷ�X�a�6�lm��ǚ�S�5�9�`@��'����jm�����)2+@1b��L���U�.�ռ��A\fM��7�{�8�ݰ��<�����j�@��Τ�z��6�іxQx���#/�p���Aq-�*H�c؈����L�#�%�9)>��&']+Meȗ�9B�<,ٽ��8��:q�xg���%a��S���w+�X<���9p����9Ɩ�5@ɩ�XX3.�S�N�X��C�>���*�멒�+_91��T[�(e*1"S��]�l�SX)RS_gL�fw9M����t.��+��	�B�m��w_S�5�h%���pI�aV^nsn�4��W�L�氭6��k��wN�u�k`͸<��l9oK���n�[�-���;6��}�M��s�"Ͼ~egr��V)��6�Χ�^UCz�����f	Pw'�]�"���0��C�x�i���������;�z���y����&<��)��޸�����S���=<��\�s1Em�;�5����-vB���5�E�f�����34����ޣJ�iᶥ�iM�Y̶�]��_ �Fk=��@�҂�J;�uqDR'�q�$��+YC`K�hM��æ	E�4ѷg���}n�ǨC��:k@b!P?Kb���w��S�10:.���i5`�4�j�Pm%3aF��X��w{N8���&�;�I���tɐ@}(J��G�|}�9r�^����ޜ���] ���prTծ����
d�l್��E��;�4J�믝�^��8P���'-����N�^^E}7�V�r��=J���2�;���l��)�]��Z�wH9�x���Gu�U&u�:�dy�Լ�����.͘���IG�\-�WdD�(G�6T��7���:^����)_���{9�8� ŧ��ӕxWg��ɧ��Vq׷..�1����t[�8���#�!4�]^�D����M�f�jW�2���.���|��2�{�e���v�B�T��ٝ��)�<�Vd�w��=�#��ʵ�شE�a8�Y���Lu7�����bk�O����G��ݥ�	m,����vyk�I:4=ޠ�	8� ��yʾ����v��|�sT�V�X�nk(�jr��)��Ս7J�8�
_V�h_jk���oجk̊�w׻�7\�Yk��?XԪ蛮�Pt��^�X���/�Z����Ϋ�I9�Tk�|&J�0����S�=
�j&�������oWW>v��9�0Q�����Ee!.�����A��Ny#q�p�����I�`Z�{w��1��&�F!ԫx%�d
c��>مGj����V2w�,���cך$�["��ټ�MǼ��-p�VV�dh2��ph˛�h�H)��e��4=$ԕ�hr��ȳځ�3g
j�1RE IUݳ34.2�X,�g���v�����6�=���d�q���kT�˜D2{uL�\3(ЛV�&G)�tl�����*
*ЬI��ʜ��HVp�Q��\O^K�5*��U���]R)CmL{��*;9Lܻ����yZ�^��w�&
 �~�&�힦�#Y�-�;f\W���VHɻ3@�+6Ĵ���dk<�ɪ�����ȴ\�#}��toza��x5���Ո8��i���X����d)�L����2v�4���65�i���n-Ӡ�`���}UTF,�������E���,ju�tĠ�yie�%�mJSa�d��B	Ν׀����9Xׂ�����2��ݒ�ՙ�8���Ѭ��y*��=�lr�� 2k7��zsq�W�a�V���"�Bp㩌��ٷ|��5��;g���o#�qKz���'dz.t�(�q�	,���sYZ����Vq��S]�~;NI#J�������2�ӂ����.,$��b�ӡ:���7\#`+�m���/Mm)l�\w�˝7*d�tmu��<��{lِ�+"��#��M���Ң�� S�>�/^����KMi`Ry+V�x��L[��/�z�t�돬�o	��ꘪ�{�>y�$xfV�ں�~>R��������Q�4:���\V,�E� =��9.u��X���!�F�!�)�x$v��S��^�_`��B�#j�:M�F��qK6�Y���8��V)�:�Ŋw�����I���3'���Q�lSo۲�.Ng+�������(g� f6��C�'��r���&KЬ��t�7������>�`=���G��mO{g2
	�Ej[�M�E�S���1*:��� �B�Жtb���}���k��CD7Mt=b>fgj��PF�in��n�mPv���S}׸�%��^��-���rmɯ��x2+YRxo%�ϭn�:�'#2hn�^���v��������F��L�;G˧< A__d��͂Q�K�u�E7��L��*󶨓ȟ�{|ϭ���ܢ�5SH�d[���l&�j���Ր:��BScm�E"tL�D�V7>�0��-9|��z�j�
�J@��,�rȨ�C��Ҹ��mb"�%����*H����W�Z�r�fp����+��!�ԫ5.Ne�ﷲ��®��NQ�7�Q��!Eղ@�7�Z��f@����7��Q�iQ"�+[/����SZ��ѭD�[�	��q��r�Pt#��o��W��$������s��,{Ja֭}����hs�{�����	���nHj7���b���r�r��I<
�~�Z4-D/��a����P�e��*l
���:xǢw{F����3e9:V{�oq@��S��VW_
�E��oU-ÅdD�*�f|hEb6o)�2��}�DR[qB���VPS�WaLVSg��~0�e�X�m��r�[��b}�B�_F� 1�k���9 ��8ǈV÷�w���oimm�г�z�>�lҤiz0�C���H��Ymz�mv�����k�	�d�y9�
ͻ퓋o-n��U�,�Ӻ]&�kg+mW6iN�)��ʛ�;3���#���yn�"Jl��D�ݚ��=�<8$�&�Ƙ��X�|��`�������|���;�L��u -�b	��V[q�x7D3*	�c� }������`"-˩�)��sB��:�Kͣ�j�P����J�h��[A�zmF��b�ݽ2V��s��w�����˧Pn:�!�4z�E����9���;�,�&yc����%�1�\197r�EAN���.���f�l���}�R3eb��rU&�FUڌ��PQ<]Z�m���4)9ۂj���l��i����&�t���ƅl�i�"���Ev�ެ�Nt�um�qZ�G�ܦvC���%��Z��e�)9���k}Xl�����N��qDw#/i5��d�C���1S��o�=��|�b��^λ�I��i�#�@�)E�|�=�w�S�E�o�͌�+P�똏'[�(�|VY@;�rd��M΍5'��H���=0�Jb���	P�Mc�z:N'�濸'�t��چ)�MZ�omv��e�Bf�on�A�4�?���v��S��zp��A6�o���2������d�o>����ۏ6���M[Qz�A{ngh<��˃U���i<��d[�XA�˫Eˉ���^���h"�i���z��8>�͚CZ��I�k�+&����k����C";�٘����}�
�:�&Z��V)���T��O1�|������4��Ey��=#�]7{+>p�� ��������\�&f�Vi�ޢ�+����Ss��R&�6��4oLݧ�)��A<Դ��h�CwL|���z�\!�7�Y��N�{5V�ע�'3�Mw��\u����N5]��SZM�r?�}wp�� ,�$G�����}_W�}����ǋP*�d�RiqL M*��{I�ad3`�&�4�{R	r�d��JgY�c��1��+�]�[�cT$��r[�뜊c-=ԶdOiQͻ��\6����(�,�3�vscݯ��tW�]=�똳Wz�'M��4KQ��j��:3Ͼ��j?_�[tujd�U��zV�}�R.�[��I#Lwy�ks���ջ.�ǯF�f�׋5���*ᑥ�㒥mvf��H%��:� ��%nQs�3gZXʽ�պ3�ھQ	�	�GS;(Ͱ������]0���1�-s"��eݹ��ٟi��mZ�6����7��
���*f�)ܩܱ�XU�S1�jP�n��y�_sdg/�-n���)�o�9ܾb`gmV@-�jIG;�G��c 8��K���*M��n��op&�Q"�K0�9�����@FѸfڷ����/C���B���@�#qJ\x7C��֞�Ź�;)��
2){���C����b�/�oSY��
.YS�� *�R���D��%:�����0"����&�;�_��2����9��ӣO�<��h��B��t�¡H3Ve���Nˑ7O�D��*�:��b��A�(ә�tF�i�9͖R�2-���5h8�4B=ւp�whc���&S�m��.V�-;�f+�`!�?�=z�ҹ���,+*m1�kiE�U�I;R�� ,s&���&n%�|Eo��1�X�=u��;,l�F��ۗ�ѫƸ�l1�ɐ6�PL�3��d5$J$�*��cK��h�]�]CW5�u�؂#��n�$��d�A���w2&�B�"����u�ѸfTGs����)(���4�2��u�Qd�wn��M2���GKF�7+�͸b-�ڈ�2Q�9u���<]`����.nn�׋��nV�X���� ����+��v�"6�n�]�,���7�j*)%&��<tn[��x׉㱫�]1q��A$�>E����y���t�oc�
��{2��u0�����`#"�S��=ٌ�b+;x�`)8��(t:���Fht�w\
��{$�q�����{u2�r���!��/4=#��Od"��ֺ�z�Ѭ�ʷ��g��<�;�o���2�yT���_qXb>�h|pTTG2�����'�+Aܳ�����5�Z��lf�I�#��q��t�IZNS	�KA�.�U�}Q*��������J��b�1+#j4O��X�7��F道�DK7��˦��]K�˞';e�z�C�+�c9�sC{Uk0���v6wH	������}ҳ1a��E
���!�4``Ob�\�O dK�c���4�{\R�
OQq�_c�r� m���8Lt�"pTuG���@z_�]xS���s�Oj��*2llfA�y�e��oCX+�E,���&��v\�'�IH�~�&��D��S
9���l��^��|�bwX����ڐ�������4���-|=u��/�cx�*`�z�(���uwj�y�S;H�RYb�c�:>.q��gD�p�LA:q�N�Q�����,ā�0� g�!��{{W�1�i�U�SU�3��e뭗���/��|�XT��vDJ��.�����I�u.����I���3xȂ��Q�+�Գ��Ӗp�|#��*>z�AS	v�[ԅt�&^
7\��\|�s8z��Ҩq���A�����v�܊3~<>۩�*h�e�� 9�G)�*�o��-=]���x� ƀ$춦�B&;h�R���q�7>n���z�'�����M��z�e4�X0t�3_�@��F�\&�m�RMZ�f1���J�^	Tz�[���~��S�-c�˧��������6�C���S4:���^&�j�KV4��l�:�zl(�q�P�"�ϓ�`�B��S��>���}~�e��i��m\6:�O+�.�5��L�NS&Kn@֙�ڎ��	��yş^ꆋm����ޭ�k^���W����S�iu������^9���pkwCn9��"���*amRbϔh&�Wsٻ�4*��u��oƝaA�Aާ�jtW��;m�P��G��<j��]��lȻ�7����Y�1��L=5�+*��P���8�^�Y<��=�(O������� ���W�h�vh��T`�g�R��xUj�}3��1su�)�g��~t��0�L㑮�
�g�d���C��6��H��,*�ϯ�p�'�X��\j�5�V����8��8�w�Wi�C����}6�y\,���gQD�������}�䠩b�;[&7Օ�S[u@f�vU�Ƿv��,���d��D�����6���e��t��@+O��`��5�:U��W$�}�t(:b�����@u.(�;��A�͆��ƫY��0֓��KG_�/ESP�6S���M�;�3��;0¸��`2��nS+)����S�"Y�$�2�y��l���0F�{<ٺ��d=h��J�"c�>oC�3�gk���삫Q�Zj��o�v��1��8�� d� ���qS0�L�yh�p�X�pЖ�=%��s��<0D����5�D�l'v��G0c`� �G��U�هڨ�q�|{C��=I� f��OWNM��_˦�d1)�˔� !1�K��@�:��g"o~�s�S2���i�OI�G������6�G\;v):�T���4z  ��<`��=��/����ɭ�%�Ǻ����1	>��&4B�2VC5�T'X�uU8�#_�:�T��_o������ǩ�������oQ��Rb�N�9�ք��'C�]癁*o����hU����{�b��۰�T.L���Kvt{�cd�8��|
6˴)�̻�%N!L���9��Wny��AZ����^��/8��&�	��[��΋b�9h�#O!�Ю�u*&�g&hSlӻ�f�@�v�|Ķ骙����sS�N�ܹ�ղ+��ӵ�<�Pa�u��]Ȱ�f�� v���E��!���k�~�T��T�_���V���C��caQu�_V��f�(u���]/�:��܁@��ڳ��'�2rVی�Q��� �|l��+����������[�L�\%r~�0Ga�Sj��.1�1=��vh�쨑���*��8�u��(O��^�'�K��K���vp1����s ų����z�x�
��������#v��F��n��0{�v=,# _E�}�_���2�.���^��)}�ͼ�]+�3��#Jv���7;+���Yb름T����&��� ��̱�2��ph�0�!�<Ҧfr�������A�G�z��_DJ�kua�0�����N�)�L7էvݍ���[�Qq�L<e$����We#$���K��S<�g������[��M�0�tB�oz���^����IH�9OI�'�`�|<;��e��e&ө��ח6���#XUGO�y��3Z�5�
��R@�u$#�k���rz�4:rX�KX<���+b���taV��M���s�̡�KY<�jĮ��Q*�m�e��w�Z7d�Wz�ȏb��r����lx6j�u�|�F�
�(�'�᭧$�������P4}_y����������*�@�J`,*����u�-v�wc��B��*��!Ӷ�g���Ӑ�ƈ���u�S45UT�j�B��ʌ>�{=�ݏ`�J
Zc�(C,:�:t|�'h!�Z��1�_6�诜۸�Eq��Ha�ڵ��7d��q�d'��5vP������OH�j��nx���4:�����,�X��thQ޷ϕ��z���Z���xbuX�n��	�4l�����I� ���	Ufk�V���?�O������	�P���i��M��ѽ1�W�4ߖŊ����j��}=��K�]:�Nkt�qX6��q���ݘb8Yہ�P��e�8w��i��Q7��ɴ�8M��Y�����;����q����%f�m�X�9��Lec�nnE��kT��L퍵�qY��}��j����ֲ.f��	:�s\���Z�`�3e&����J����.�����SG�*��,��s�<���1��y����V�d��=�كU+�dKE7q�]�; ��ޑ��\�5��,X��v����0Q,�[6�ֺ������삚�Q1P�d����h3�'�̹p2�ޞ�ޭWP���ON�6Tl''CwN�Ή�NM��PN�^�]O@��.�G�K��#8z��޾�f���L�b~�����Q�~ S��@U�����kΩ9���ˊl�|vxE���4n7��5�C��'OD�����|~P9ɖ8�:�]ou�M��h�\#�e�w	�-K�+o��t����	1�Z���������ܼ���/�c�]��/F�B-gZe�Yxc!��p�F�}gD�iII: ��z�O��|v���h��N+{�0�f7�_MD)A��5��;�Rt��~����p7*Ymc���{�ħ
�7<T�h��)�<���硋T��B���w=w�_}K)��ju��e�]?8{0t�"T$��4:�0��n B������b�hV��-\��t�n��%f� �U�"�Ȑ�Gq 
���\s ���	�ȸ{3׈-�/7dޙ�%��k�lN�F0	�;�������"����[LU�_�XX�s2��zֱlX�yl�Tn!_W>�"�JS&M���9���h�t�`/���8�����cyƷ2�^��+���Ac��=|S��<̍�7�V�[��f�7��
�^�Yc/B�<���ǻ=��c����ȓ���,��$�6��c�ɩ��V�զ&�G�朼tp�,ܻ�!T^5�{��+���dyJ�T�^I�.}R�v�şt�E����΅�_<���������/���;s�q�i�j8���	�e:K��J��-	���	g��0vUâ��ϫ�O`eo��+[���tf-��I	��E������vk�MW�c��{n�]�`6�>r{-ɒ'��Am�n��	Vs/��=��Oƽ�Ѷ�h��W0~���Z��e�pT�K�O����r�^rY�����%R @ƥ~��V���j���"�p`;j�9�3MD|N�EW����N&���u�#q,�o+2n`k '��s,����7m��*1��<2�i����t�W�m˗��2L����P:8�	t3�_ECǼo��2���z
ơ9B%���}eOiGbLbt��{+�퍀D`q*�]T�R�ȅ�t���:c3�0���p�>*���9(�W�;t�gk7D����%T� w2�aO{h�p�X�m	hŽ����K;)�p���j�5��AF[�R����p5��>]ǳ�o����;�}uwn��i[�[B�%����6Zu�Ȟ�Q��V�l��]�$��C��S�>/t���={{ׯ�����7e�G�x��-ۼ!q���S�rLt�%�[���tF'!}�&���L�ӆ�{���b��0�ͥ3��'�Sˣ���̙��d�i-媴e]�mQ��ق2��&���7���d�@�(�d����q�63�4V��Nn����{3n���5�7���B]z݊O�"x?�G��$
!��W]�)��\��	[�^��vx��Q4T�[G�p�/�3����	�3A��HϺd�ŬX*�α��]�nt�Jq_��X�&�����&ьԘ����|�b5�1q����j8֊�.��5�������?*�v�TKڌ�f�!����/�J�E��s5˻�`��U� ��Ѻ�;��o��M�u��2�צ��~t��
+ً��/�f�=����=0n=��JMqp2��"��ɊsՍ
z|Lu@��7Gv�NK�",E��<�ޖ2�:
3�0�\�ks�+���Ae���!��uLO{�x:��FZ���qȃ��]eV�^�*8�[Z�n:����K���ojw�/�e�g�!����]o^�p�N��e7�Ӣ@��[{9��z�<GZ;�&^����A�\����,Fm�{�/\�P���8Y������Skwk3�����b�e�j|�J���M��7��ő0�GH́�W�a�����k�r<3���駫�E�I�}��7��$Y��g5񙏤�s�{0M�ڊW4�b���E�s�\뾽��u�8����ӱܥA��"�`�|���`��+E��Xx[��5�q���ǦP޺��y�"YL�\}3<��������~kw���u�7��f���?zEG�I|w�R%�!�[��L1�]s�!��K0���Y<^�+�	ix���_g3��¡d�Ճ���7!�|/�/�`<�̡̬�sn���Rl�.��k�!��HvK���@��*��9MDI� p��0���.����H�@�N�����Eô�*̣�o�\r!��P�ֆ_޷|{��)�u4��H)�����c�ho�%&t<HP��^F�}+C�t�l�8�ƈ�x�'m��4��7W�7����k�fp�O�b�B���W�:>U	;ArՖs�F2i�q�W	�붧�R���-(���q��7�4���_���N�9�d!h�?Wͺ�X홙W�0n���m�;l�_$�@w�E`
���r��n�W����F��x������{�Vb��ԾI.��V�p�������������uJ�~|j͇=;�Bc��ۚlʷK#WJ�l�٘+��j}����;`�&�gL�9É���5)d͈`1���2���+5�Y���Ү�����:̩�a��=픲�F�Q�γo��Λ�l��͔
�ܘ��eF��GK����dΨ�As���
J��e*(.*�g(ެ�ؠ�&�e�Wzr5:ɸ����3|�$�ׅ@,�T1}�,��y�w=�<��Ӗ�n�ǴNJ?H+�R�N+Y�2��ڍ�I�`�7����{vJ��!J׾���|q����M=b�Z�c"]V�'Z�F��������i�/����S���ve�# fQ�c�����7JX"0 3�_.y��2%�c=��)��cr���N�|��S������X���{���&-7��%
x|-���i�"�b :�yæ�|���8ئ��Bƙ�ɧ��B:�]pѸ�_Սm�2�BL-��*?��C�P�| û���ƽ������],����\�ˆ�1r�1�����WQ��<	=Q3�X�ʆ����.�h�Nի���M@�1N�ͳ�c��D��!��m\18�Ϡl�R$�z�L�+�5(Go'����V�b��g���iT�u���(1���i���C8�i�1�f��FS��s�,J�/`��A�``	�����s����u�p�3�q��H����W_�h�%��"Rf%����|r݉���=�/*{�R���Ɛ�Twy.����ȅ���*!�9q�-Pz�` 2�7���O��೮}����V.bq����ն_R���a�[������؞�EԢv�Yv%d�Z����ݪI��!ѧ�?��1�x|�ȥ%�i�i#\55�
]MӂE[���m������TQY�������6=�F�c��%|�[�1��*�7����`C��}EJt� ��*���iƼ��Qʘ�g��_�̈9r��ۑ�`���xW�;����j:�)a]�&�W�5t��X:�DV��s�J��indw��sl�;�_>�T�kSnn�hE����"�et7i�u愫�r���lBo(��ekIJ��}��n�vdt��,�[��:�mN��q����y���3zs(�m�(k�|�LNRH�����,M���5�o��i�s��r��b��ݱ�9�|V��[�V��CZĶ��;����F�Ӥ�R \9M4C-�-�^YQm�3���<��S�A�:;���@ꚑq�+�5�ӝF�ׄ;�l�����o&Xj�jZ�wt�m�XK�L̦:��i�Ƹ[b��L_/�ӝy*b��}pţtw�|����ٯ���D��U����iYFxu�cäTغ���ˬY���";��-���S0����i7���A�p�f�Փn�:}�j3���jJ�/�ڼ�2�K�0�������Q�_P�YՁ+��owy=vٍ�YK/M����7n�3{��V'�Ut[Нv�kϦGR�z�9�S\0�س׊��Q�r�X���2��(��r�vfNC��\{��n��q��o���Z;q�x'GM�=#�F�u�|kC�%3���ٲ��z�(��5�� 9)��c厍��vD������K5*x6�3���:�ʒ��U�h�w�5T�n�>Y�+c+{^ogk�K�$e�G��ذ�Q���r�A����n�i����9�ds��p��U����ϕ���̾��θ�:Pńf�"��4�:�Zr誎^Q��%�fj7z�W���s��x7���£�e�@��6�਎Z�;��%��%��>���m`y�*bͮ1N
pD܍�6uj��[�SPA�~�F��ComS��vĸ�����)Z�]ƌ۳v�|��)�ʕL�A�����k��x��{V�iü��5ۘ�e@�+Z�i��ކW|�Sjvϝu�����̩]�0�Ĭ@���j�	I^"�s���e�����w�(3`�e��������I32�s=k�{�����ߛ"۸!Zv��[�/*�y�t]�p���kv�ҹ��.�%�b���)&��w�Gs79/����|*7=q��'�����n���>`Uɯ3Q��U�J��q�� e�DJ��'�s�m�R1���]����"2�nŎs�G��+�ɺW(�r��,�^;�r�l[��\�Nr�x�����6�y�;�a�k�9Û������wR[r�l�m�y��Ƌ%�W��.K�Y�F�;��Es�\71�L�k�9ʐӺ�9��N]Ewu��<n��Fܤ��.A��v�W(��sE����^*�^e�ol����^(ӻ9���v���n�F9s\1���Gu�˻�]�o-����܎��\���Ĺ\���n��q��n[;��9s\:`�K���˃�4q�wv�;�r��C���sx��;�<M���H��.k�8I;�*$(��lS�n[���79�w�y��7����8/���$��W�\�ΖV.�Щ�1&r�X[���~���.�4:ƅ��I��}����o���R�M�{�q��r�����_�xW��}V)S?S`�KA��y�H��x�����v�����u�zU˛���ξ|��u^/�p�ͻ�[��:�->u�m��=�|DD1E�߫���|DF]ihQ�y:�Z�WY�H��F�ѣ�D�#�O�F�W?x����կM�ۻ��]_���h���=y���s��^���U�[��W�~v�;�sy�����k�okſ=�x���#�M� ���{�hv*�����+Ι/�"#�}�G�]G�!>�G�[����w�����ү����y���y�E�U˛������ֹ�W��~ok�o�oKO����6��׍��׃Q�Ȓ�p������l˨����Իw���B1��"0DX��~���>�����",G� Bjb(G�"�#��_:�U��鷏ϟ|����5������-�W�r���z����sz���~-�z��!#d�����2r{�y��k�ݍ.����#�E�����>�z��������o��7ſ^5�����^֍��>���oKţ�~���b+��^7��|������?�����~*����g~V>0��f���+4_��]�y������k��D`��#�LX��@�>����߭�W�����o׍�ۗ��[���m�x+����o���n���羵����y]����>�>����'G�#=1LU^W�w�3����{YH�3�ͫG��>�!��#�����a�V���_�Š���k�^->u�x���x��.o���o�|�{{U�s}m�����߶����w���޳���e�Z�x?H�`�?Ϣ�2k��0C��"#��1C�|@}(��~����^ƣ{�����W⽭߽o������x��ߕ痥�|W�x��������u��K~���]������I"�>�>�#��<���R�R�N�I.�|�Dp�"=N�>�� ����}?�>|�V�����A��k�����5��������om����^-��<[�]�ߗ���-��םzo���A�V��+Gգ�*��S��z�_�����_u�����>�"�!#�=?DW���1�UG�DAG�$��/������y��������+�^-?��������nm�~�����ͽ�o���~yW���}� �?}">b ����嚏]�pro�U�ߺ\�5՟ϴ�������E�m.��%R���{�{�,}hw8Uب�=��ش�����+iL���oÞ���#"������8���7�l��#�����,c��ͩY��]z��p��yv�ùNAg!�<�U�GX*Ƭ��Ig���}|���1^�o����~{���������?|��W�-��Oߞ��ӻW��n_Z�|[����j�Ƽ_�����~-�ߗ�<��k�^5{���_:�c������|���9�^��ټ=!���}�I������ݼU+םx�����z�毋��~~yW�������_?;\�-�����u���h���C�b#�Vg��(dʹ"��{q�}�}���#�<vb4DH��\�:�u�W���{�v�����k��y}6�W����^�����{�w�zW����[|����߭�W��=w�}n}�����?A^?|��#�����X}�s\��}b>��	��C���>�>��^=�>y_��~-��w���^����TE/�������;����r�{�v�ޛ���ϝ���{^֏�}�W돸D`��Y�㟶{�I��<6�^�Z\����1��}O�"�!��%�Z��ץ^.~��^}���V�-����?E�,��G�>�鈻?}C�(DF3>-��n|\�wj5��<��ίkN��
�>���LW���v�A��1���y��G��"��"<��}�#�#=^�{|k�m��כ����>�������_��[w�~_~����K��~_<׿ε�z^�u�zm�ϝk����[���<?}#�>��>�jO��D��1ӎ�*]���w������-XGЊF).\���|W�x�}���\�Z7�{�����o�|^5}�[�\��r��U��[�^?���zU���_~}�{_���U�w��ub>�C�>�k����&�1��}���ϻ��^-�;��o��~6�^�����m��ޛs�v�v߭�{��[�}xG�_]�~�G��w����#�K>y|k��k���W��ז����/��3�����W�GT�߳/{���O���[�\�}���[�}��y����ޗ��+�v����W�Oz����m�o��ߞ�_��������������~�{Z-�\���筿箵���>����/H�����W�m��{Χ#{1~����$�����zZ5~����4������oM�Ƽ_�����Ѿ/�7z��-��Z/w�������k��kϝ\��x�'�d��~��Ɉ���a ~!�p����Q;��#��x�QIp�e������:�]���\Z���*ק[�K�&�_P�����kks�V�ֿC)�?ih߰V�s֐��*_��7RX�D<�!3��sffg��� +��*u��M����dIu����mg:��"��D�͇?���������W�Ϳ�z��}���ۗս?�O��7��7��S��mzk������^+��ww��k�꿛���_����|~o}�[�}k��m�g� }"��D�V�M�����k�nG��|c�#�e1��"!�#�ߪj��!���*��>}�{W-���ߟ�}[ڽ���뿗ֿW��m��Ͼ_����s~��u�W��v߭��y�����οTV������2#��n�;]{���|^5}��7־/����|��Cb+�����_�O���<�zo�ռU˾z�6��߿{o?�����{Z�����5����W��.��ߝ~��o�n��<��V
���X�bO�q��k�����4���*�W?�]��z�|o?z^~����1���O�0�P�Ȟ����|I��}u��h*��������z�Zw^|�7��׋��{����h߫�����~���_@���>�����s9���� }���zk�^7�ퟝ\����~v�*����w^z��m⯋�����׾�{�و�G�1(��vb(}c��ΰGѹ�=���׭����_Z�k��-�o���}^�ݝ��e[Y��G+���W���\���]����Ţ��}�������^5����k��=yش���W��痧�oj�.o��Mz__ͼk�|^+���m����������n�߽���}�W���>6ח�1����鵳�(�y/�"6�X���|���AG�G�Ӏ5���|�~+��Z��wk��x���|��5�������y�}_��i����zo��x��{���}���|���^�/fȭ����ы��,�DCB>� �y���ُ�DH����󯭼�������^._[�?7����oj�.7ﯾW�~E��O��������j��w���ݷ����U��ۻ�0��!G� ����>Bo�<���k��=���D��=sUAxCD�v�7��h���y��x���^*��Ϟ^���>5��?w��V�y���޾�����K���/��W���x������z�j �� ��}��G��ry��e��w}}����}���ܿ���o��ѹo{���߽x�Ƹ~n�|_��~��}|b�����g��ϴ�1��㨝�wl��	��������wu�P�z��X`ko(+Χ+hnb�H�ÚT�s����ɣ�cAZ��hwaQŗ��)�0uZ���w(Pǵb�����jr�gl��"ubhlTr<�볦�ףF��� �6�Z�Ƕ��Cs���r.޳����#�����48� G@`5�BQ�-�q���I�c�����J�������ws-;�i}^�w\ӌ�D��
J���2����oQ!�����:&���z�S�mZ:Y8�@sϨ���>�So��B���1�]�uL׆'X�El�sᘻ��}˦�+�\�Sr���23`��b9�9*����Ϣ��J�$�pj*{&�Ӝ��׺�{��j����S��w�5:ɸ���̋��Cfn���~7(t���Z�	�}��=37�;��cգ��~�W��}�g>�uLJ�ڍ���fė�^7��p���+��?|)��x�#�����N;iQ�d1��}$�Y�sC{�:���q��e��-��
4gL6o��@f:*�B��<+��c��L�Z���$ߎsN�'��������/�G�����^�r��Ŧ�����B�|���^ U�jz�-���b�&��w�9gh$�.S[��b:����ݞ�&}jah��Q���'M	�Z`�`�����픛�0Ba�3}�K���H��E/o8/��e*PC	�*0x���32�����4b�U݊��\��fVM�S稙�&�l����Ǣb�D�!���=\��#�vU�o\�ݭ8����+��"eY\�Ҷ'F�k����[I��4���N��[�@�+fPLr�M��ˆ�Ʈ���L]��Nq���fLt��S`�R'y�鷣��ܼ�id�F���EDI���F$��v�Ϛ��Ӑ4C_6����e�����s����|q�D��F���1u3ͫU��)A�k���Rt���~�=f�õ���==8��*xwe��(��|m�t@�V��(AJ�{��2=�~�_��.W\�)�L~j�y`cx��]�ޭ&lt��\��yQ�u�P�?�@�P�)c�Q5�4�*���S��9�9�8s���f4a4ۭͻ�ߌ�e3@Fr� ��xwe%^���Hf�pv�k��S]���l�>�*s���p/>f�0E�uLUX�b��ϊ���-�6�w�+^���df3�^���	�yu�L�<��9�5�q������8����^��*W�׻&��ǻz��Z�����;��T�U�w��W�~d�\���>G�րd�QYݗ����(�W��Z�۠�uF�����/�Q���S��S�:F{u;����n����]u5K��
�}�Bz7�G�T+X�o���7{N$�}L��;��8W<ۼ�z���ٰ�����s�a_|sgRK��]G�~fm����83H�e��Q{�ȩ����c3d�1�fɧ��T�5*ޓiEl`8���
��.����ځ��ta���б�Ǐ���U�]��z뻶��ɬ��rl�r��4 �ǧ��Mnf��b�C�~8���<�N��������u���r�1D�)6�uP��(1��>ok�\s��q�+h���ö�����|%F�{-u��<���.�.�C�Prz\��y�T;��V_ݶ��j����<a;{sZ"��j�Ovg��9KE��PK�m��q��u�U�`2��nS*Z����c�*bPgt
���{��o �L��A�*�B�:J8.����+�1]c|�>�ht�3���)����gjwG[z�[���ֳ��p��P8���qS0�RJ	����C\׆���������步���ه�RQۇ1��N���eõC�r�ҡfL(��3.�A��L�P��
v�n����铙�+�.�>;�����`��sA	��͢ Um�Ƭ�S�K�Iڽ#�Ata"��u�p��GΈh㝬�w#�&)gܩ�ƏE�hݝ��Z�#�2���g��*^Z�I�{���̇
ɬ�;��Xq�D�#�mp���XOpZ�Aֽ<r�5ՉeNZ���G�9���{z���14hǔ�Ȩ����I͖f��6�szÈ��Qp���ӗ����R<gevk�����(�C+��x)�ٱ͘�`W�â�$�(dǠf�
��h㙎_�g)��5:�hL�#x�Ll�[y���f${�H���5ʼ?������B���Rb�N�9f#\�8u"�2��N�nκ5�0�P�w*��~�����ĩxj�!��k����+�Ĩި��9�Y���U���ș��x ���b�vP~�KT�tV�����w�����R��x�\��3{�� W��.1�͖(9ٶ�s��������k�g����沽h�=�G�l퉌�f����d���b�1�1<�'s-t�p������m��a~M��R׏����GAU�_������2K�cwu��q��7�1�WB��M4�^o�'8�є:~󤭜��=��ok��Fy�K���ׅf��s�~R��
G���V�5�+L7��Q�b;�� �C)�(�z,�{�W W�g�bp���\ڼ�r���u���8�1�b�[u�,��?t+��t��7��s�lp�q:o3�Ђ�ŘsS���{��3@��Fr�u���>�i��[�����a� ʊB79d��\��
y�Y�������Ǜyk��cI:`�iYjt�3��-������ca)h��;e���L�ځ��v�{	�T���g�j�.Z��wZ�,��u��S�J������C-� �")�ύ�++��E$�����|aUH���.�ڥR'-����Ob����~�z��|K1��C�=�C��{;9%\) w&�XVAc@����;}�_l�v>�@���C��ʢ�G��a��C�"9���Ep��w�R|���1�yyf���3�p�4߾HBGA�S�
�]�T�=;l��/N71��:�ހ����m��u)(��4Ϊ�M�( G@`s١(��:�t|�t��rՖR�8mja��W�ޕ����������
m];�i�����&�:<�g������� ]t�M�[������׻���Bp���q/!�`sȊ"0	�:c���2�e�T#4~·HDW���j�	��=z}�8��g-sW�%˦�.�����������0&9�9*ώ��W���OV������Y�:$"�#���4�	�F�Ӛ� ��a`���m/`Wz+L#2!Ik$]�G#cR��qg�R�]J�t�i�oj���zc��Tk�bVmF�̊UIٱL���nW�KxR%ɍ0y3�q��'���Q�U�ر3�f�ST��u���S�K}<8�VR��~2���'RU�*�&wd���>w�Z�(L�rkv�QZI�5 �.��}�R�x��2��L�jJ!�NVvYe(9���®�YXP�/���֦�V4�\X�P�b��c�Nu8��*p��c�K�����Y,���坨��ђ�Nh�q)�KBc뫴��+��A��+�z�� O��F�c�m��Z����IP��+�}S��g~~X���{���g/���ʺc���,3ש�h�j�&�/'h�ny����b:�%�����v�-BL/�{�1}�Ubo��bՕ��wbK��P��咾!���&`�,o}+o��U�ck�}S��|w�4ߕ�Š=�S#��F�!Ga�{&z��ӃD1���8��]]��1�������]sc�L�9@@]�ʭ�S�����ʩpxp߽�B���2�n���^8�{�z~^��z+���^7]D	��+����P<)T�=]s��/2s��;ܓ�-�Ӂ�i:eZ>������,�B"U@�0R�&������ر=���Euf̘C��[��0�`�[n��X�*�Ȑ�q� S���:��mEpW|����!�w �9L��n�R�$(Y�/:�Zr�`���׮�Wq���\��
���j�ڪa���V隙��Ư����bB>�3�튺�o�ǜ�v ��壛w��ڮ`�ʄi�vl��ZU�C�RT��:̹Uw]��9f��[�s���Y�=�*S���)�5��.�:�*�u?���d��Q�㚧�������Yj��K�]�W��.�*�ɓp��9�3Z����S�K:��;�}�^�^ޠ�%�nX�,L��?\�X+
��WP�ri`�T��xxz�8��My�$�I��f�����$�# t��{	�C�c+��R���Pd+�_l>���hЧ�2۬╥Xw{C������(W�ɣ��O���j�b��@~��a���<6�y].�ݯ�sp�����j��̘�.���9�7B����Mn�h���_�>b�}��F��fE�|�kݓ�EV�L0��3�UP�1og�oL�U=�[��Eo�����z�fy�ĮCz�3��r���|m����% H�u̳�N�a\�3n�B���<2�|n��,�-�[�r�(�:a������U�>@@�8��]�A�\������ϩ���A�3p�9���N���>�b���qc��#�
��(ส��rMW��L}oC�1�E����T����Q��R�53)�\��֎�)��	ʑ���R��W��*gAk.�8�ee�{7�^�+8�8���q^m�N�"7�LWa�RȤ�уl_S�.�l^�Vr��)�%�/��yI�;@��lW8�Ae�wv {��ڥ���bO��6ӎ�~E�o��(�v厎�u�7�y6He��k;&�Gq�(�qAq�F:ݷyWf�6��Ř�����䈃ctVLd)��3�򁞒ѝ�4�k�b�nWݧ�j�[`YqJmM��U��][Ë�҆9�wQ>��$��>0B�c���d%�$��+��p5О��"sv��k*'X.*A�!q�X��oɀ]�S�Wb�����N�ۗ*�V�)�7v��ܥ����p��w9fTi�/��8�-bT�c縫2�-Q=)�9Ak�%��畵��������f�PS�+r��z�RVԴg�s(D葖@;K8%�E#���3���#K!>ϝ�}���5�uzl�X��D
>�X�q�Z��Ǖ�,����qS���',�U��]�B�=���mD�=
J˜n���u���}��}���'�w �J���Q��WEflx-��s�N��ywt�Qx�ͯu�"��Iw��>�j;v�cl��Φ�v���e��� ��H[�ۄa�4f32��.�;w7uv��5(8�Z�؈�Z#��vxc��pyu\�1�t�8��4�����Gws~� ��)��):%m2�㗴G��E9z����a��Y��9��RR��cR'^"m~��R�dA}���٣1Y"ܢn�RY|퐵�l:�v�L���۷�g��oB�|�b�����z��t�Ζ�@�<��YY�=�s��t���˻�u�C��K`��u������J�J,ʹo�[w����U�x&EE����#��_=y��5�ע�������{{��c���'^�Ρ�X�$ Ï�5�r]�i|���X4#��[8<k=͓�ɁBŘe���/��љ�;D�,�7J�m��W>R���4���x��i�Wc[�X�Ĺ�]B��v�pou�u���F4���WjM�X�wX��켘6�"������0���eL<	��O���eg�,�����S�e�놸�'�W0���B�m+�8	z���	�]"*���2���L���ZA�\�u��D#�Ft�];�����.tA�D��εA�݉���@�(�XV1wU�\�����g�k�K��s"���	�Wo)A�M�I(�Ȇ��qM�f�f��Xh�JE��X5���s�w1a�=:��-^B%GY1�(��`Ư��4ѭ���J���u4^�t�۽��-�dR�kl�Òtڊ��m}{���a�0�㸨��@���m��)��y�j��JX�K���v�
rܥs�DM�yF<|��v(���(�r:�Jb�uή�*�r�-lq�zk����ø�!��O�T�d=��k���]y���DΉ쿾�
� ���;��b(��I��b���(�+��A)�ns`�鋥�����˛Ǎx��ܮ�s���t��ͮG��x7GwU�:t��㗋7wh�sp�\��ws]4㻗I\��3���s��Q�S�����Ar.�E�<��;��s����M%�\�v�7�Ǟy��79ӻ��v�	�w��҃t�s����H�͋��fm2wncFs\Ys�����n��K�r�w4ș��$�\�+��x�9����M)r��-�&��p��w\�\��˦g�ڔ0QE�6�ssNH��x��ѣ/<��'+��$��9�h��\黮��+��n]"��^h+��;����s]u���5�n묖�sx~/�����y��e�3�xz�\��]�o5��fe�p
��
�^^ܮy�X��7�%��z)-�5wL9��v�P}����j\�&��k�*;Z��7 �{~��@�M*��%�vvhc^oAT�Q�ܺ����848LKF-�v�sN�Îɔx}���Q�J���"�ˡ�\�v\����"��
yTS�J���w��E�/\�Bi<���B U!~ۯv�����{RN`��
w�V	��ou}Х�E��*�`6۹n��M|�$���
��9�3%�6��)H CJR^�3>��¤��,��'3���ց��=�s�bz^Ό�����^$�Y�f�\���P�1�3ٲBEq�0�tY)�+F��U�o6�u����DMz�]ew!d����}A/�l�]��Z��
�y7��Y�R������`9�@h������3�
�P*9�.��hZ����=�
򊒍֏G��v=�Y�tP|j���br�ą92�mد#�^P:<Δ���-�_���ݚ��<���Q�Q�N����;�C�P��!��uLOg߽٢��*$e��8b�vw޳}��Rrs�eU
�P��-���(�W kiB+�Fv�����nq��-o6 D���(˴��V�sK_ �S�.�o_}gk�ܹC*9��rՆ�m�r����=;P���
�4�j�2%Yֶ�IN�7R��/6Iy�u��6J�.��.��\����)ٯ諭���g(�w��ݧ�W�_]���N�]1��J��@Ϥ���u_oF��6ڋJӃެk5E$��d�9t�t9}Β�p[�=�up�����`�2��o�
��3�5b�F��4׫yhPث#�+��i�?&+.X���t�Pz�v�=i"ۺ�7����EdS�d��	���B �-*�!u2��ԤM�H�-��?;�4^�WWX�wJܺ(PO����L1�e�)�ωW<} �(�#Ğ������ץ�����{��������8U?-R��>��k�!��HvD�������� Sa�p�v�����]���<>��̂�gV-���(�Ja���"7�;����U��K��kv��r��s�cdH�qD����1����L�c�>t� ��Ӎ��q�7�83]�ąf������N��~���b�k����{S�1p���򤝠��7��K�vb�K�\��h�4��M&��6�*�M:72BWx�#C�tV�����Aʶ�
T��msE>�/:��f��h�n��mn��el��󦬏��߂�`�����׽ĸ�\�7�ih��N�߹��f��Q�s:�a�B�����ީ7Y����e���5�k�c�
z��.tE�ƅ�]ʗj�g2� ��Jޭ����W�W�|�H��&p�h��7\K`�5�"0	N���G"8�.�)�C�oϧ��m�ݎ>��/j8Go]1˦��W��K@�����b9�9*����$����oCv=��m��c�T����GY�v.�s�� U��͇�r��<���d��N�V�Q��C��[��/I�q�������;����8�g\���^�d�����!v���k��S�a}œ!�8�N3�}*p���@T^���D��R��`�*u�u��7�k^��U�m�#�y��*͌F ���0����
���7JX"0 "އ5Zj�2��R?t���);���������n{\�/G�i�b�h
c���~�{T����b��f|�L3�ʹ�����uˮ5����UW<I�RR0v�_a���7���<��91���;�ڦ@�L��;��1KT�d��	���f3���Y��[o!�	8�g@���S#�TIc�B
3�]�9�Ǐ��
��G�L�j�r�;�,Nj�Ə:Z$V�WL4i�`�B�`���~Ʊ�ü5�'�6�q�F牭�����Gty��9oiK��� Lo���dd���M�5+6�2WL.�V瓖��mq;���tb��x���z���ɔ�m�O�u��_}��_=���k=�A��@��,�H#I�&O@��/ꙎeR��aJ`���G�h���M��u��ӓ�8;�쯒�b�ʖo�@� ����Y
=��P�E��X��%e%��p<������q7��O�U)���,�" 5P$*�n	��Q�¥Ճx���k��y��e�n A6��k����ф�ͺ�/�X�*�Ȑ�Gq��oE�uZ�}�Sr/q���7��~Bb;4T+��5ۮ�5��.�S�`ڪ�St�*���Yƫ��m�$_�����6�����h�iZ{����TP��L�܁�3Z�gDغ�n_5��v+��/�Zc��Q�:,{�9�]+Mw^\,����㟙)D���,��G;��T�s�oh�W��Z�2M}� �0���Pa��(�1�F�2�Q���m�ީ�jDd�o)�JѨ�p㚠��0�ۆ�+O;ʫ;Y;Q's+��|h!��KH7
�4V(��w^�ȼu�p�T�7]����{Ё|���]�Ѷ���n��Wat}��|��vS=jy��@�F��gfj�t��WG�t�ʫUt���2c�a7�ѡ�A�rCw{/����W��ʍ�Fb��c�S��1l2^��B���K�i�����Tn����OlL4AK��6���f�[���If�15��b��v�T�de�h~���>���%�r���C�Z'� Lpc�u�����e1��C{\"��p�y[F-'��caņ�:}���We��P�)Ui�1�A�p:� �s̲���+/�f�w)�mh+����V���|\$�����$� !PN��S/�.)H*L1�1T
��.�e3�r�b��ګÔ���Uw��f��"Y�$ߌ���.g���T�S�&�+���c퉴�e�ŋ`VE.�O��{bژv�5q�9g��\;�$��>�����J�~�)/��!W�P{Ǫ-j)9��H`q
���Ĵb���Yۇ1����<�Mk���r��h/��0�݉���io>�ϟH�g��}/�ǵQUǕK]�O��$g�`��4��e���	}�NH��ƹ�-��L}���P���F���R�#��tCG�`7���݊K��ґn������ǳ�Y�N�]Iޛ�� �<"�J��d@/�D�aT%���s1��3��imVt�QL��+�,o�m�c�X�m��$GK�k��*�A��0Ӫ��.��G]��Z��O�(���X�_��oS� ��#Q���|��N]�c� +3.��I������{�V�=�H��r�u�޳��/Jܚ��l� �Gjl�.��q���K�Q�oE�"�9A�9�=�9�z�+5csƍ$\�}������}�v�ؗ4��tӇ�f#]�Q���a�c�=��0v�5�����,Bw��B)�z�C�ܧ��l��r��a��e��
5�T
��Y���+�c�Y�lR4���'���o��������YC�M��#!	
rR2!��2�F�Ola�) b���&Vk�nzfl��DS�v��6�Z�݋�	9�uLOg�vh~������[,#�5Oվ�B݆*�h����t/����.�����%Ms dIc��ت��n��H��7�C��V�t���_�9ip�C���%l��z+���u��}G�s0�/ab�����V��B����W-���j��l��+E7���O�oԹ2���u�X`���aW��Y���������ee:��A��1_w�mÖh
���B���[K��kL]>�DSwk���o˓���<=�w�	�2�{H>�_=%\�� �(�Ğ�3������u���x���⌴n�x$b���U=8�K1�d����g�^+��ӱ��rC�1�g�,���s��(G8ij��Cg��+��%|�`��ԛ�B�ó��/�=�;va�cE���gU8��N��m��G0�oM�(�V��WiY�I[vsOV`]}+ �&�I�i��^�RR�u*n*v#cJ�}�UW�V���d�B@rF�8s5Fx�qbۊ�(��Ja���"7��3����7�s~P㒮�\xX�@"�v�����xE�!i��ZC�m��6^�Mb�L.��b����ȧu�a��$�#�K�u* @�ژϟ*�ˠxG�H}2�Ϯ�w�c�-�spW{�Kr�9 �d�ͻ�)ͻ��U4��t�	A�c"$�rj"���q��N{���݅"�k��y��sĵ�2��D`	�d)�tx_�0:��tn1*�ꦞg��Al#.��y�묭�׭��*e�nX^|���.0���P��K�7u���;+~�,��r�p�E�ѿ��	��lB��w�>��&� F�2. �_�wp�s�n7}�!(d�8�"F��/�����Mv��D�x��$T���qZ�&/,,ˢ�c���Sbi(����mnc��ɋߌ1�'��q��"T�9q���ֲ�.b�Lf��^O����:���5Z�F��ys��rqdLT	�B�N�ʝ�bcn~(\m��MV.n�M�G4CR�]��X��Ј>��k�i����Wzv������SALk&X}�$��w����Uh0߬�ް����8�j�2�����[���7�i!��RzM����s��>o�E�I���Akq'���{r�����B���������t�y-nz���V����@ϥ�c=��|�~�a�G�&r�h�%
fv�*ʏ5��O|4D}���B� ���sI�1r농ƺ��ƶ�u$���m����b��wޝ�P����!�
#Kj�X9�&�!���&b׹�L��p+wYe}վ�{Z��5�`$��Z�����B
h�N7Hģ5]�9�9�1���1��xq�Iw���Τ���Fw�ZԖA��/�}ܪ�Sǟ/��`�SS;)N�����{�A��Na�q�2ʅUx	 i��P��OF7�Ev'�6��ift�Z()J�l�<7!��&�븞6*������"�ߌ���gr�T��޻�nykwȈ�6�L7P��)&��s�����m� ���3"B`ǜ!D.߂%��۶�*�E�u�n"�3��~B{4T$�<ۮ��ֆ�c ���=}�֤�kn^��_4n�MTÀDg��+���_�Xv���7�c�(���&M�n��ƃ��4����:S}<��k{=#Vj����]k:r��W�t���������9�3�._�8��Ģ�l����1*l�,�X�W��(t=�8jl N��W��_�4��]�#�E-�}��������˚��H��^�涮�eN����O_�W�TG�zߓ.Һ�F�@�~�%*���(���a.S�K��;�]�Gn�gz�RVƱZ�8U���š�ߤ��zݩ������8� �m�Tk�_�G��R���^n�RP�)C9P����Ud���.���)��q�qZo�m���L}��r���,�6w3�Q=�{��.M�X�w�8xejܦ6��|��}=���t U����y4m����\�R'l���ni@̑�Z��}��W
��O\	� ����J���PcNCzeҞ�-?3�Vni���㛹�L���y)����>oJ^�h���@�<�*)��+�/�f�I���*�k���V��TǾ�G���^#:�|.��ȟEQ���^�΄<����8q�����VVl��z�:�u����xR�8�1�^�
��Q���4ئ}����2�'�U��`������gi�p�)�~��)$�3�L@/�L!E��܋��^�ך��M�P�V����BZ0��s��p8S�P�#��F>�d+ )�ٯu��4�nߚ��T�{�L�Q��+0(�Y�&���m(��5�����	se���m�f�(�J����h�>�D�����_�'x�BZ�l	ma����:��k��]�K^���*��v����[y:�W6,�OHy���\�^�4�~��ꪪ�=�|f��B�*[=�u_h����Tp��>;�����`�fB��K��������׭'�d 0z���YB��.���Q{��R�#�gD4s�;X��	�m�o�Y���x���7�wu$�.4I������@�9�B�����5��%���s1��N��&fQ�U���],MŤ����<��4�;xk��*bE;V�GoQ&���d"��C�F����7:$�|���Ɉ��#Q�Q	�Ȯx�\@=ѵpV�\���-�bg�˪�i�V[�ƻ�i�vm�Tjӆ[q��1����xؕ����S����A��k�*��C��5UlxY^U'��}�f��3��s��0ֱ�E���`��4�{{���S�b��:s�E�����o��w���Hy��/���cL�z��HUܦ�fW����F�d�]�&���=��U�/j��e�n��*��y)���j�v��r�Nb�:�6��d}/>�^O��Z�I/�9��+˾�k�x9-ݻ��bN��_`[��x�eպ�ӭ�^d��[wa��$�OOL��;pX|�%\k��C}|����{(��C}��3�MOt�^�Ȑ=D� 12<�(UM�Mx����k�k��b�+uo������6�XJ]ܡ��u��=�(��J�w;������m����y�b�'	��մ�#��PN�+�d��kU��7l6nX�tfԫ�Jf�6�-�e�ٶ�J5�\w��Y������ �?H �#�O~>�'Px��@��0��jp"�t����յf���Lx�S�iP3uSY���r���(�8+��� �M⏀�Q]���f�ϭ��OJ�X�B^��kA����{�aỺ�0\��[�Ϸ�D(�vX�o�G�ܬ#���Ww��E�.�5������.��
s���|�1���g�(U�<Iu���9h����R��n0��V��ŜJt˃1<�`�r'����J��P����tΈ��TX �-T��w*�dD�UU�`�Ti_Y�-
�j�u�s�Kc�n�c��K��XE �_(��a���xp�;q��=���{�Zݬ�ub���g�W>"�;��.g �I�^�-��;��4��-�c M�+6nݻ���Aa��isl�D��"�gk�){d2�x�*�m|ڳR;�}�4"���])�6�U��*����y[��!7"�,���h�w�UAR�ܸԌ!Y�-�՚�� k̆p��θIi����@�`���Q����f�	�+{ �4��>�ͯ�D�E���h���Zg��N���wU]���]>��E݇r�\�c�bDy�9CVD��0�;ӧkͼ�ǁ1z��\2��;�hMY����d��kzn�
m�k��tyf4���=S;u��e�(5���Їs-�[�������&}6��zm
ⶰ��_��y��v3��SS�Β��
�nB�ϺD�9���2F�}�V
EV:2����Ly�.���+{��j7{
��8�g�$���4s��n�ܴ�އ���O�fd�⸂�p�^��i�سy�����ޚ&d��!��2C�v�����L
��ȸ�������Z��0k�����.�����׏:Ќ�%&i�e�<�^�g�{׽M�vA�"y�,�W3�����²�h�Γr��OZ�xJfD�_y�pj�'f}.?/�eq%	�2�w5'Y9}ۅ�� �|m��t���L�(���1G,�T<kz����"Q���L�"&��b�u��%\�ڦ0�ۧ'E�pT�Ƒ�V�\v�uKe��R���ej/���e2�x�L�ٽG��:�}��5(.-���(�Xq��Ӳ`��&G&X϶��]z��`���.�ߥ������,N7vhR5u�}���ExD+]�ǩt(�Ԫ@:�)�#j�J�IR��G�"@��u�^;�C��5�IS����r�cx�y�]�]�\�<F�;��t��t���9�b�wk��k�5!�%�<�fd�L���
b6ww�t�����D����6Ln�;��w1Gv���m�NW��U��;f�5x�%	d�;G4����aD]ιr�nsi7#s�!1���v�R�"Jw] �p	5yv�s���8o8�ܼox�Fe]݀żr.k�\�Q�;�4\$$c;�w��u��֏<��"J1������8N�Ѯ%���cF�]1�WwR�H�+�y�	9����ݓ����s�h�3�M�㻫��s�6#��;�����F(y�^ut�Rm�ɂ����A% A
�q�%w�}n�Zގ��ۼ<�� ��{=v�4��&����K	^�����o?v�^$e6q05�t�z	�� }��s�ڽ<���
T"m�_�����z+w��f�Sj�o>�Q��ډ^_r<�yG���da8�x����(�Ϭ���5��\�9 ����Y�ݨZ�9��J5����}r�����p7
�\0�3�{
ns���@���8=�X=9rㇵ=�|ۇ��<�^7���ؽ�U�ol��f�[�TU�b����=�R�M)]�	k]��gv�&����C���Z�P�2�Vl+/Wܦ Ɛ�H�}6�}��_�uj�'�L�~�K���c.�v�oڇT��U�ﶇ=���,.ا�}=a�����%y�$K��6��b�{m�B�s\B��Wh��u/?FY�쵸���~#����M1�y����ˍv�Bt�4��2��OL��޴��ゞI�s�cɈ�x���_ZL�����q���zwjI��;��~{��l����@c�v+޴�~O��9@�j\u��,�Dλ�=�LL���ܾ�[(�m��ȻȨ�c�3G>�Tǳ{�m��oҖe��{e7��V�#��*wS4f��������Q�s�4(�3h
�kd��B�F�ĹX2qPBz���������6��^�-C1~�>�W�����4��ڵqζ��k�n�Ti�]8��e����Wϼ��sjס����y��ퟜ�xyɞӻo}X`���Y��{�#�|��G��|���V'���L����'��ev�2ʪ쿞U��v��4�%�w_ǧ�Zo]뗽�o����\>Y79N��:�n.�w%{��tNp5����T\�৏���yݍl��V9��,���~%��n{�r����]�1GP�˛�v�\K����X�OF���ެ�]{�������QJ��_I|Trߖ�W���|�7��}q����h�"}��9����7}d�Uy��F]���q{�e�W*j��᫐n.�h��9NR֪���kum����*�\���lW�!�J�:������v���/$Z�������:�q�����]B�ˢ��	*�~w�_X����S�X��ty~�jܖ=N׳��P�XX�nԙG#X!^"�KJ`�OW��7p榔,�]T�(�'��Ȳ���罞���\���4��Zͥn	���DUK���GZ1�Ц�,�����t2�q�F��v?ӯ<�H�?  � =��{����}S�Ww#��!��OڇT�2^��������
4�=k8��o5gx8�v�Gf�I4�������snj�W9�n�4�����g%�P/�fl���e����BK��m�nׯҸ:\Ec!�[]�Or�=�3�Մ����G��R^���}�Q�'��}��Ϥ�d�X�%�b\�	�ss��,��ӆr&!(��V�Sꁷ0Wf�m_vիs�Y�����o�Zk����⛁��9��D��t�[P3DK̩X�e:�l�:����o���FV��6�m�p͹G5��usY�d��ј�Oؐ�j�zc�r7����r��b��s��I���xET���w�ƾ���Ʋ1��xk�f�{z�w ����c9�r�S���T�)�����y�b�b6qr��}+˺�9���",���v3�^����mD������]��h�.n�;0����: ��� s���j����`�SD���
������B�5�v+������� ����I��//�V�{�/H�
z]	�/����=iH�3�u�gV�ݱ��,k�S���$q�>��}�Gm�������� �bgk��X���{]c[=qV;����uTI}Q*W�%�b�tQ!�2�q�͡5i��o	9R�]q/�YY�	��<Lo���u�z���^G�I���r�Ra5v�7�����m=�+9\³���EQp�J�{����69of��O/�Y�����/&F#[Q����S�"�SŜo"�#SK�RW�*�s�mmJڎ�����Gn63�3���)6a(|���"y�-�v絛��֑�Cg��K�d�7��W�]��na�/	�����BT*L��)�S%���>����}=�%�Jvj����d�>�t�gl\7L�2棈]Qh-rW\�b}��h:4Ċ����y.�d[���&�l8�ЎD��\Ls�=p�Ճ���XB�c����>�n�s�]�_vOoc��J�E��6�Z�\ds�_��Og�YS�M��$ubB�7p���.� z��0�eq)����H�Ҭ(��^װة�),�ܧ��z�Ӓ�����%B��7�ł&�nu��FM����e'C�.�L����Y���`���{�t������3�c��l�J±������*�{��k4V_��Ǜ����*�s���ᚋt��7;�,�ȶ+�����;_u�q��fi�y�eg9���\��	8�q垸�1B0���"��8_��{/g/��E�f,��ʉ���Q5���S�,/+K�B�z���|�r/����'����m��~�D��D�}C]U��s�ѭI��ժ�w
�7{a�[MdK����N����6�L�[��G��i>���۪bS{Ȯp6Z��߻79M5r���Yɬ����C�o�G�Ư�4�y��`�rRU�-��[�z�z�\����V7
�[Z�G3���C��r�5��<�$�V�T�B����kn>z�噊��sj�{��k��fO�rv��Ϥ��͝yR��z;aWN��z<ӯS�s�2\-�
����}�`Ƙ��O�{�X�U3��L�&�	�T�u��S�2�v� ,�a���ź�XW{m�Z.u�e��c��`fǒ6�k�<�W���R�P��uzQi3��E�9S��i-Z��1u+挥�rD��îq�]�ҫ��f	�7K|�&:�7��tcT��ԣ��W�U}�U>\��g'��<��wj{���;N��)���]?
D?+Ϯ/r��}t�∯I����i0�4�0��f���˚�T^��Q�Ӱ��$��ni�����[�Q�{x*�̶�4ˍv�D�v�)�=5IǓQj���v7�1�����S��ɯ�Sɨœ��Tm&6�]�3��M��3/3Z�\����e��퀶�f���9�ȟ��WOW�A��\8���9�U���r��5_F���T@�����٧=�Y\�Bw�G�������ԝ�P�S�棕�z�ǵI�N\F����:��?g;k�M��gy�E��Y�n�}�8�jJ˗��z�\����Q��5\�C�}~�CJ�f������Epؽ���A��.
x����X֩n��G_���v�[�ҽ;p��}�E�.P��#yss����3Z�3��8vx��J4��L�k#U��q.{�{�
��C�u��u�
^]8hs&z̀�t��3�u�I��kܷ��@K*,r�`2Mǃ��d��d����r�l�i��=x�md"ԫt;�U�.u����Sn�j2��g��+��1Sٻ}L~������jxסq���� 䮁��*9j�j5��Cym��7���=��us��
ާ1���W��"��G�:FF��s<��}�O��`J�{b5ɷ�@�����9Ecwp��!���Hi��dd��BL�Q:�Os��� ��>����<�[]�n6�_jG~J0+�F�|@f�M�,}��V����)]���opt<gjR��亅�H7h�(���N��^��p'�WÒ�[�١T$�b���
���|�����c���F���6u�x�W��y�!.������Щ.f����l=���=�c��7�w��v5Q�!��7���֏o����Yط|9Ό�o�HKP�ר��V�@��ظ�y{"���~�Wѧ�w�>G�� �|:lwV�rW6r�Gr�Q�3M�\�+\a��ث�n��o]28�ao���!�)�E��|;�Z��Mu* ��9��z�h YN�%�uuP�8��??������{��p��5l��K~�/���`+l{D[�]YE,w�t��HuiU�(�V�����ڮɬd�ߞ>�I����������Kӗ�~U���Zfs��������3��[�y_Z�>�v�dYF�,`Z��Y��z\K�Q=�*1��տA�Xx���Ǘ�����]4o+U���)�|�\��Ss���1D�c�<�৏�!��MU�����Qؑ��T�4�*�m��ca��3�^���.��������Ē2��9���r��=^���v�t�H�=k�y�����ь^��ؼ[U��ok���0�7�ޛM>��ޗT{#��ڽnJ����*eo�LٮY���3���w/�����n����~�Zg9�q�*Ң�(������{�7�.I�Z�E;փ[p�=y�Ӗ�H�0�w����=�G��Xn;1/�y^K��=��xs�x�\,G_A��:��S<�Mt��Iڅ�)�	E@��an�n�����j�NQ���JY��:�qD��S�'���{:�����wGq�홁KFX��S0�������IR�����5��kx�.p��⾁��B�/$�h�oVX��g.���,�����2��x����veJ���k��
q��+�'&�l.i�}�G�De4��=E����a�U��u\����V��5���;4.��]��t�S�V%�bhٜO�w�����5
e�G��mL������y���t��H����H����}F�I0�q��ȟ����v��=^�oN�4�ȑi�|�������c�c���Zp�|ۍw�Tk��tu:����}�ɮ	eok�n�Ve}/�ѫ&��_s���ᚋt���Μ��2�U*k�]��R��>����&�TJ����'V������v�"�H�-v^6+kZ���s�e�No��2����u���9�YT_���3;2�9G)��5Ƹ������׽Q��v�`�5k���PNA�́�nn�-�v�(��,��.�5�������W?��e��a��{�ٽ�b���.���p1Gb��E4����Vu|���ݾىl��>�u��mr�o�����y|bVZV��Ρ���g$����+����If���(,��K��6*�M\5(<�v2,�\�$����S��v���k�f�%��`T�_,Q��Q%F�v6v
�j��c�8�`ֳB}��P�����N�7u�����N�W�UW�^������Y�.S��kv�7j���낳��7���zs3m5vA6� ��~ʤ�Q%򿕪������5�����Gm1Z�v�*�o�T�1<��Sh.3'�]D6.�zL�;ʫ�<5�х%�{��/�҃�^z.�$�te�?�hgW�ʇT�����mG�'����D�nX���ݳ��i��gT��
Rv�k܆�E<gjS��2xϺ}��{r���Μ�V�9��MS��c�7١�M+e�v�0��ߜۚS.j8�ү�7Sy���k�*��\D�d�cS��r�y���̸օ�Bv�j�%<����ܚ��np�b)z��V����[��Y?n�W�Q�I�_6�]���]��9}�nu��5��FD�%jU���W�dl�s���ɥv�c@m�-�}b�ݥ��k+����K{�6����q����k�f*���Q+Vsq:��O�XY2����W뙶����٭+�R�Ka�Q�츸6bX|�͵�ڨ��j �j�Ј��a�z�.�q�m��(�vX�7��t��M挔�Fѝ�V�ň��ڧx`��/��n�<l����ظ�Y���"�֋�U �b�,�K�]���&s�7b�}`ZFn�c�׏^�G��b�EU:fņ��E��{�핃7'NW�N��dS<���g�O(�]kمyr��<G���Rќt'ܺ�!��V��C��^}��������Zx A+���n�@]G*�
]ˎxpBnr6�z��N��I��Gц���|�,Y��AJݏ�{��(8gr�]�{s�u����]��M��u)7ީj���*Qs��w�u0�i�W{��.�rr�i�pz���#N���ʴZ�Q�+Wd�Y�����R�/f�D�W`ud�a�,�|;qep�u&{.�1���j%�C-N�~�X�����\��S�!��5x�v�b���J��C���5�:��S��x�¸� ������rv��R�̫�+��vv��t�#!���I�7M:���K�IL!*Ŏ�A���o|M�-��b��;���(K"���[s�6anU����8��k_�a�
`���-wa�ܗ���ouD_nk���:�f���:tuZ��غ!�
:�/�,h��'�>D<��VJ��VNm%�V���YH�i�ݧb����:���we��o{8eiܮ|�Iѽ�!"5���|: ��H��m��6��|(B&mZ��(^�{;h�Z�X�`{��ކ&˭th`̵\�4HeK�-룪��e.p�Q��܃Q���]J:�k�eǝ��0�Bd�i�\/{t�)��ݓ�]7��&m����B��@�
��͝Q=�.�dK�'V:*<
�o���a�c�*	�xq����˔����K�ʾ2��hHIJ��n# ��GU����I,������B����h��}=e�Vz�p*��K�:Q����[ٖz������ܱְ���`M��\]]9��[���i+iڡ{�7b�wb{�Q[9�*��'@�)vǔ/d�MSCnmi�K���
�E$/VD�_� �Y:j�t�n4(hw#�k��5�r*X�"��hq_,�ɣr\��fn$(��<:k�[�e��fėn˄6��!K�ѽ�v�^c�����o`�?
���|F��2��^!/�U����T�Ai����%7�!�<7��$�%iq�9�3��|��Y��#]Rf&7���"��h��fq�\(���e���n���г+�B���n��]��V�X�J>m�7�9�8�ap�;T��R�
���Yqv�:y*�(G[��3b�`�tX��J�D���F�C72�Yh��+����"V�Šb���jf:	�ڍu��y�B�%��3��×{5�T�)�B�>��R�Юdm�s����M܏���a��p�s�;�q�1E�p�s]ݻ.\�(��c@���XED�Q"JP��A˶dF�#w;t&i0��Q%�2f336M��9����LWwL+���湐�c�����H�+�4ɘ2�˻�5�ۉWv�']�$A��W4D�]��IwWe\����FR���˝WdRQ�d�cnu;�nWwt�����Cwt3%9ۻ�II��wFdwwN�@�˥���c�6$ӻ�A�CD��l�Uˀ�H	�r�H�P �71\���D�fFPd�λ�n��s�`	�p���hЎ]jL!N�"Qb�!$@�D"P�N]��e˩2`�����x��������w��9�A����4��w�P�27���u\��f_h�@����b���}����4^%�(#������>ڦ	�[�r(I�F��{���?i=���3*遘�m�/�M1���ך���Np��gr��I��^oF�ʌw��s��P�}R]'l"q�.��[<�W�ʨ��ъ:֎<��N޷y�9�cY=�'NOS�nz�3�0Hf��|�R������(�}*F8��cyss�;O���ȹ��(��l��z�>�c��uTI}R��-��kb��򞍑�YI��Y����y���Z����������?�����_�k���^� *_�5=O�7�&A�7e�k�m=�+��̌`l]H�,�\����]����J�O/浮��9����/a}�N�({��z��2��F��B��9-�{�ضk�+��Gk{��3�:�)�����L1O��׏[�|��P�]��l�f�I4��s[ϙ�����P�L�o����ڮ
°^�P�!4Z�̈V[e��Q�c���ɹ�|!�bkL�3�z�掮�Jo=wav��8�o��1��Y¥��S;�Hk�!{f�e+y�K��7wY���@�kN�W�E=��z�ʍ��Yr��#��X�ג҉��B�9Q�T@�!>��[�a9��
��j|�h���~�E��K�4p[g"R�+�6��F��Z侹�Y�On��W��V�Sr�gk��q�xMƻ����*�>ɵg��z��F���x�:�Yرv���&�}���½=�ޯU�z�L�3�������]���:���`|�MK[0?y�jVv�[W*�������nv��M���8��1���v���R�����m�D�_bu��~=+O�\�׏s��iJ*�<Ed3����RΊ������3������AS�v��<O'�ٞ�S�@s�4�ҹ*�o��$����p��3lϏw�!�b�ы�5�\R������b�����;������oUc[=uc��*�U%�J�Ÿ�tNnƸ��Z��fR��'���}/�YYɬ���t�}?�*�x���k�>i'sF�K:���5_\%�L��1�W���tE-�m]�|�
��[����2�֧<a�q��u*W\%�u���k.*���!.B�^�k^l�v��1���9v�^k��I�ed�¯�
�:��Q6�|�J��K�OU���%UE1�����<�e�����ZM��r�ku�=�����m=�+9X�*����+/7����.����}%򿕬�S��h5�����y���i�����^_)Q��K��Pߚ����+z^JR������Ό��ɮv�[�	P�2��d֩.�}�Li��ڟN���%7��6�W���,�&�Ŝ�x�ˬl�
���2�>S%WH]_��N}q{�y����kϣ��~��M�vE����L�
�g"a�e�#�]P6���=W��u��&��\#��\�5��G.�I&1�9�qq<��@}U~����O���%��z��T׎�*5���6�Z�\dfR���c�t�����X^��?[P�ls�ڭYY4�#���؜3V��\̫/v,Iޙ���x}�L�{e���^f��������L��h)7k�S�7����}M.؝�6Ȥ�CVR�L�՚�ǋ����%g{s&�nX4�׬�S[4�f�)���p�;僐���#�a#��s��@KT�"�)2vu��3s� �²`�P��g����f�Tb�����U�C�}�}�W6����s�Eך�z����C���^���O�1TM�T��Wj�*p����*���S��.�����{��o^��us�`U�D���ܦ��Z�o����/U���q���Y.�[��kg��wQW�L
��$F�t=
��nw�rw�6�5o=[�����SM\K��Vu&�x�Ҹ+�Z�v4��C����J����\r��������o.���ꩭ73\M�ի�]T���\O�~|�JU%�V�ij{q�Z���B�f�Usש�t���+��.3'�YTh6.��ʲ�M�:[�����V:vԴ��s_��\�^�<g*RV��6�ϧ�R�u[��Y�}=���fdަ�i(g5�{��3���:����1y
9V���;�!��\������ݷ�f���p���b����9�S.n";�qe��0:�����b�;WI�=1�:������j��m�����^+�^v�9,l�cke�p}�(v5��6RO1tj�kG6�a�x��ȁ�=Ve���N7E����Cw]�ƶ-)Y���f�c4�I}'CY�E�\b˩+���3�c��G�U���� %���MD�ɬNc���\�6�6c�r2� z����Q7As_q���rJw=�,��x�9*5�������<�j�]�9�ˉ��EÅM���6�켕�����l~m�C�t)����o��#V�����qfu��ſK�+���ws<��3
�ȵ뎖3�z�c?)GV%ʼĹ��h��ko�����qι��u���9|2�1D�k�ҰZO]뗽��1�ͫ}���ٱ4^�Sx�CJ�T-����D��#�p�Ϝ\��{ɿ'�ʹ^�/K;ՆG���	�Z����v:\�]^�g�1�J�gOzr����*av��K%��)�׍d�}\I] �!�D��_B-F8̹���-���z��T�i.-=�+:�[�*�����<��]���n���T�W@pt��r&^��.yCz{Ur��n��$Go%B��w#�5�m*�:w�;��>���>G�V�7̏s��[�9Yzj9�7��I��Ղ.�yIY�wPnZM��)L]���o�lyV��qݢ<��CM��x�*a%���]�'��T������x���x.3#]F�600e��:���fk��B�\IƭZɥ)��Z�d>��Rt�m���U
�3UM�:�#T��W�*	؟����-�ǲ��B��o�S�v�R�u�f��.��QΦ��RK�u���#O���,j���Вi/��o���ka�vg�T*f��B�/��o�4��j%ne�Nc�BK�v5��Z��X�B�moZ:q��Ȕ튅6清�jJ�5�&�Ń��)�{�q[}�e��"�ݪ�&�)�ƅ�o��O_����cm}G�cg��.j
���|zl[9�i�To&���l�R�W���Ae?_/V�/c�3���u��ڍn��'iļʉ�{z�~��W���8f�ǆ�{4��x���	+'�:��Ƨ��Ӭ\Mk�Q6��^�����g�`��z׏���>�0&�P��j[�ȫˬv�Z���7��Mf\��:�����M{�_A�ֱ�rC��(Mw�YX����ХZ��X�pɉ_#�g����J���x�b9B;=�� ˍN4���0R�W�S]�e,���&���e�܇3�W�Cޗ2����f-w�������!�a&,��������p��>8����j��G��;'��w�h�`>��sqJ}�Ⱦ����?'���c�^Ş�k:�[ꕡ[~̩y��p���Ի���w.���uħ�pު��늱�PU���/�eC�l���;_l��C"����gD�؋sp�}r��W��Kq\՗|t�Q���L�^^w,����U��%j�+���=���X�
�Wp)U�UX�ef;|���8	A�?}_D�u'��+Y5���h5�C�y�3#h쎙k]Vgj7�D�+��9;%�Q%f�s�)]��#��75=���4��'�c�y�큞'�{�}��.�"$�������R�:;/�>2�����c�zO'�s�gp6�l:�5
d���ls�+]�P�|�̶^���纖f���p�5l��a1p�C�~�dG�PX|�ӫ��B�j;��v�TtLdKne�i��-?{"w;{���g��[������O�	J΁���7�U��9s�Շq%|�PUزux�B�`�Z����<�Z�VZ��R�Lem��c���
z��4�.�T��Q���[�8�
:k�U}�������&�������.��a���=[O��[��)�g�M�TV��U�ˉ瓊�#����Zp�n1���v�A��o�S�k���X;P+v�����
ǘ�nin������ZAqU�ч]+��N%�q����V���[|qy����粋;��~p��aB������Ѯ)�Q���=��O��-xf:?���լj~��_����6�y{�ڥ�p1�ݮ�p���n,v��:��3n��Y&wu<�*�cw�|��{�UMq:'�p��>qpSMW���5��CS��yS�v�[~ry�����}2��ϥ�ꁒ��b��\��SM�{⳹���p�����EhP.�� �] �/�Tr����[�z�z�75'��Ӿέeu^U�tބ�V�89������0�(y̫2�M�o���*�!�Zpsz1�T���A�3�"]N��`X�X�X�֪�::��-&��[�p��E�9��[9�i��}�l	�/loӗQ�ն�c'�Cۗ˖.��y�FN�H��Pa�:�!�0�.u셓�ڌk��z ��=�u*37��J1��>˭��b��aK��[P����wp��!��;���I��ƈ�gE�'�WڒY�39.������gS�r��%a�u�������f	��I�]+�b��*��u�'��9�q��OڇT�VG|��u<��,�*�Ĳ��k�=sS�e�]=�M$����)��Nm�8s
�e(�y�}��7dԸ�3~��=+rq=�૗3Q��q�*�nP�9�nH��^��+�䥚�S�>,��g��jK�7�&u;�Gyp}k2�v��]���-�F��g*5�D�*�S��yٕ+�ز�I��9R���U.�l���*ۈ�ᚶ�m79Z�b�v6:�۱���:���ie�n��欉�n7�VU��K����{NjyF��P_LUr.a�S{+^f_g*=.%��X�ͽC�����\����Q��5~ �:�ڕ�H�R���vh�]V����)	��Dh�7w���v+b�@��X��ݒ��	����,/��(Z����B��	n���T;}�٘�O����_6#5����lN�wkpw1�J�jm��Ka�r���빼���ރ�#��M��m������==Hw���y�e���Jk�K�{ׯ|0?Y���}�ʨ���E܃�R��C��dF���Jk#�#����y4��6��_{����܈���P�3)�Q_�U�&׃������5�a���O�"Z|��٫��"��G�?��W���[��FCԙMvb�ű{��˚����ըz��m8�T.O�v8f!�<�LvV^&�l?�5Q'��k&�R�5�j��Χ�r���nL�nC����J��>�s�|�u{��Xn;�>�bLo�{�he{<v�v51Z�.`Y�}7��Ԝ^�؎����%cW�[١$��|�kkbCn��^ެ��N5�����C��׫�e����Dj�R"y�U�ݴ'��!:��,�g\e�.�0ofp����;�G!:as�-P6��9�%�c���hm��j�f=�'(�����&��#g���������~mh����(���u�z��D�b��+ѷ�A�ճ��;w#oT�%�ᩥoY��0�e��t7&���ʇn�`X[Z��Ν�����,
{��.0Ղ�$�{aZ`<���\A�E�=<���y*Nr����/H�H����@�ij����c�
咽�ϑ �m���{h���o�l5���L�tb;��l��OE��%���~5h��,�H����1_h2���3��к�面����!���r�0g��c١n��+��徹��Ő��Kw��-\p�~R{����Mt�{|�V6R9	�Yr�sĳ�!6�^[�򵝶��E�m���HM���dQ�������4�N{�q�[�pѵJ�s(V�62��vX���]*}g���ѹ-ҫI��ɚ�kax
���M��*�pmZ0x�= �V�##�gU�\��Z�i,���*�3��<J��]\v��3�����Xj̳G�%:���];���M*��S�妗�1�i��!�q���ٖ����֜Zݍ���DsÇy�N���'KD��6�l6�僆L�`
�zFoD�2���w���=���yȨD��aS�r�k���t�[��F�Y�{�"��Tv���{oq]��9���F��S�b�w�U�Ҟ�pd�����o:����9�L�?q�/mδl�}W}/;���;���y!��69%�v�]��eo���Ќ�@B9��4�=x앢e���)��ǺPt3_%fpK�+�����+q������w%��"{��Z�Y��I��ku�N.!��xs(D�I��zE;�ٸ&TJѵ>TP�Q>K)a坔�>Jn���	_,g��)*P��o�dזV�R	���aI��S��$�|$!��Rw�.��V!�c���u}w&ر�Ҧuj�.�ˤ��j	�!��P�i�S��i�]��	��"��&捡�[�U�KKt{&.�Tm>8�Q��yəG_n��u�서J�C.�B�8�	"������T*���ҹ�<�m�ù7�d�r��2�#(Ԥ-�_m�cuVW5QU����m�����
�y���g#�ݩ��+9��V�i�V;��{ۧ�ڬUn��)���/�@��2�7�@�a��օ�j/m8��4*?NC]f�}f��8�މe^��pj���̄�A�f���ѓ�1����k�iq( ��3���9M�KR}٪��1�	Kh�� �\CS�w��v���7!.�����cl��u]MvfA9
�"p���m:V���!(���h�[T$��+��*��jt=�W|�2MX�c�܍Y���w<`��3�Β|��iXS���wkr�J`mΝ���}�Iz���j%�A�*<We˛ۖ��DRǒ8jr�i((�җ���Pc�cF�$�I �2b�I�ВBi@�dӺ����I�$6$�wt��0��$��r�ȳb�l�QwvC3hI�E$���L��2���E"��,LЩDFM�Σة9���I�)BA�i�]�l�&�8 #1�Ĳ�d��0 02"4��R����a�fL�wBP &!,�0ȝ�M21LA��۴��SBR$��A� ����wI�3F.Z黝٘H"4li1Q]�& �4fd��1 T���	6"�I�r-;�\�9�	&�1�d�c2�j�	�P�P�(���ߞ�}����޸U���Ҁ�Օ��3Rq)��坴�%���7�X���S�NF�]U�+IX�����P��_oP��Ǵ�l�F�Q��|�`��B9�.&9۞�}�mSձ�[�4�51�OF^Ώ8�i^U��.�xO{�6�9�V�ȟ��"�,��<�o5	,��p7D�ʈ��n5ed��//�"��#���ƊU�t�[�]��w)h���f3o�V��沵Y�X-'�#��m�@���!�7��Pw���7W7��3(����X�d��o�*?O*���,K�S���=��v�C��}�Ol4��j���J��.r�C�ɚ}�s�Z��a1�j���8����)��7�������PU���J�n�on��o>��c��!u���c���m>��Ϯ
ΨMl�����v_� �r��}y����Y���B�JƷoCv�,K������g�4gg��{'��C�\�Ӫs�)TI�v�d���cz���ʉ�ķq���6�<9yY��ˊs��q��� S�*Z�I����r�|(��yz�?A��TWq���*N{��N���Y�0Ih�=�4����9����"_	�×�u�N�1q�����f�l1�JӆY�1S�v�K��s��N�N�v(���}˱�����z�;�i��}�N���O��B͖�|�wg�e�-W�$�]�}��e�.���S�'%��Ti�%XS���;���e?>U���fuI�p�'3��C;��gi�9rG�TC����Z�`�[��nMٷ̌�s�%�\2�;gV�D�l���וL��*��-Z��\�_�jyd�{�}˨��&1�9	�C���*�V�O]�k#3�{�׫���g�M}�&;^;�J�Zp�6�^IZfh5V��Q��qq�@���Z���5����煕ʪOW��h��u���zl�z�.R:�͎q��5����V���9�.{��w}(�`���ܮ�k���i�׌�����NoW�et�|qcxMhu��o�5����N��׺z��\T�)��6��Z������PU�4H��⽆����Wv��ݓ+\�{�x���T�o,tk钬�7ʡ�^v����'4���5���r�(�Q����Y02��M#�DF���S��b4�!�]ΦE���ͽR�k���v��o-aэp���t�V���3sr��8W��Ui�v9��m���K�S��CO݋�|y�|�����O+���kz�w�ܟ-��zLREѕӉS���]_@�}cOb��)�u���H��sċ52��$�^kw�m�ힸ������Q%�}*9-)tn��o4��}Y�2z�z�e��=V����g(�)h�`�*��D���\��75²�5�5�]��%&��&ۇ��D<�^7qp��!���Hi_Fe���N6��+�}tݼ��+��ֻ!�ί�3��(v^���&6��PJ"����9��b��u:Kf���Z��J��{��h�x��C�s_)��fZ��6�^v��`�&#�Z��w�t�hT�J���8�|�����$8��.���iD�KS.j�F�sq+rk���9s4���ylm����<��6D=fX}^�+As��>��mL�%;��Ln�]�:}��U�j�9NˌEztX��c�1h��[ 7ἭT?c��3�E���W �x&��)��Ѓ�L�u���5�=5\��4U�PV���gϯF*3f��%�Е��
�k'��b!�}h�	-m���1ym��VvF_`�ke/�ꪪg�9�w�=\'��|��v��F�Ȟv�\
}P6�OfT�r|�`K3�(���]�:6�e^kS���5m��nr�5���:b���!�ཷ�B���}�=V���S�eZ�/:18�x垼s)�ʿ��y�nf�x��M�-ow��܂T��ؖ���2�A�m�ҰZO]�k���k����eўr���m�[��Xd��ʾ���Lu@�ظQ��,�����S�2��u��ԡӊ��=�Ĳ{���e�_��\�:�SC�^�r��~K�i�R����旧M��S�1��U�<�N1c���
�˼۸�rd�*h�M����+Է�U��v|�-Q�����Kr���X����7C�SP���������Ci��X�m���P��^͈���z�򅫯��z��"K�q
�M)O-�k��Χ�r�:o O\p�|*�Zr�{�N\�9��޷�7}��Cl֣:^�J�zՍ�a2U�E^��fi��~�2��=8#cAN�w�QH�I�9�mnZF9���#@[����3�Ǿu���D�iSEoax]��j��,��s���n�:�-�su�3��4�1�j[ڥ�Z,���V|=꿂~wQ'�Wm��k�����<l}Y�=j�5B�ˇU����|�l%�X��[1١$�`��wf�zyVP�����X���ا6��U�P���]��ރ�hD�	�S$��Ԉ^���o�b�M����M�����6�^��z�~�*�;x��$�>�,�'����r�5	&
n1�9��c����.�M��&��<�]=a ����Lvի��F�ӆk�m�ڈ�9Z�"cl�1�mG��G]�z���5_��<��[̼= ��z�
���,T�ϓ�zf3���4�)�yUk�����{�gy��ߌ]��'���e�^�د��{��_?k=���i?�,����%������y~�X�������IE�ocy�|�������E\��Y�T��~ޙ�)�H� m��{;4�W� U5g�q���ӏTx��:�TT���Qi�w��2�74'B��]�\Β)R��fA.n�p��y�z�&����-@���3su�������|e����\�#@%i���ޖK��+Z�T��~����)ˠ���S(s�����=������46&JK� �x��[�]ٽ�<��N����/�b���[�������P��pˮ�� ���r89�u}%u}2�*)w�[���x6�ډ�v���m��Z�w�����d�*0�v|�JU���\���֎���a�\%�é���@�Ⱥ��}ғ�4�T��6(%�B��nLC|��:-�/92T3�ð�Up}5�-Ϲpg������b����l��zc*�|����W� �䛖����a�q������v#ϨR�ʓ�{�OV��Z�jnI׽.o�.��Щ.i���q���Cv�%ʹrsp��o�:v�j�4��'��ޚ��8�f����i$øeƻ�]2Q��X̓9��g�Y�^潆��ީ+s."Sɨœ���%Fӆ^�����o~���{=�+�N��t�Ű僔^?��V��t�������p�㙨3i�wN����|r�|3#ц�zn{����e�e�i�1�Se9�zp���Մ{ӵ�\���`o�wңb���:�W��^��r��}ԣ�*>V1�\��]��S����J����S���Ĭ�v��f���o<�,�����we�&�w+F���B6�l��[��_�fq~��k�'u��F�ML��]�.#�����e�$�]��Y�{/~~�9k�0{�f*�FϦ�����:Ǌq������Wݪ&+0�8�6��v����6hT� �`���q�+7N%Q78\.ю&;
���4�}.�n�P���w=����	u<����~UD��P��d���&;79�U�yF�gUd�Җջ=M�kR�1�kg�����`U_TJ�T�R�ݜ�V&vDT����{�䌪$�\���+9F�Z�����D��|��4���ָ[j*�7��vԢᦕ�����Cڇ���/��R�����.�ˢYzhe��'�r�-��b�\�iR�Em�c�p�g<f��%�_j�w����F���m]�q�\�ZG��d�*�r���
�ZVLܼ�k�u��My;#��N�q�TU[�fӹr���g�Pc�ʈ���o��M6.�;�3fn_Kh�H����{� X�]���Ұ�}}��ob׎\��z3�܉���Q�<��w5�f�+P�V;ޗ����^e���z���xι�7��J	T�:t݃z�vG�	^��N�#��W�\^�Gf�I4��e�v�0'�Ƿ�,wK&q����76���Mq�Z䭹����&|���H��8� bC��B�|ʍw�3��1����q�ԕ������دeq���8rSo۝;� ��Iqm0[q�����ʸ�6�Of)U+Q��P>����������ٓ�V���[q��5������j��:E��d&�n����ǫL�?������Y���8�q�Y��)�J���h�.��-���jӵ�����?g����{{Dł�z����r�.X�kZGm��)���x�s�Ȋ�9��k;����^�~~��
��O�k�(�nw��O_�g�T�v&3֨���.�GC=Sŭ��eU��5�<$��i�0�"�\h��ysgu,���s��ٷ��Z����>b��ciuʹ�ԀwmAj����i`�2c�M:2*k��XT�2o^�v��$5�&y\��Q�3�6����ukq�hġ��9Zߘ�QQ�u�@�s��y��d�>]��S�:�����f���nŗ0�YV]����b���p�[�Q�N�m>>�Bj�D�ͪ������{��K[�}��켼�Y9�o9�J�ʚ����կ��{_6��m�(��+[�[}�����p���P�u'��+Y5�<���u�n8��C�{3��I?On���<;���E}'��ۡ���\oa�4!p겹$�-;�� w�xz�egʩ�'%����Q!cW�[١uc�x8�iJ�op{�q4s��C;��{m�)���.��	��D�� ĳz��a��w]<�2��AR|�Co��gh\g��
m�}�.��V2�q����w�/��Ý.Wd�F,����QI0y7и�qq<��uGU4P�Kq�u�����l���Ccj�����7:��z�y�k�s�qZXT�Q9^t�ݎ���bz��>��� %[�j���M�c���⍺Z�:\�A�o��Q2R�x�jOVL��V�,V�>C(��ե��Ǽ�6��\B3��]�[q8�UpEW�����gC�u12��	�"�w)ҝ�`S-�������C�ϭ�k<٬���ZY] �]��1��?�(�T�d�Q[�=���&�5��o�7��^����O��������3��O{$�����ZPsZ�\���=��;�ˈ��U���X�Փ�/�J;���;:�弫����%<�৏���y���V�����2��&=���I�l]g��zW�::��~�|�����m�ުƶz���E��d���bi.S�5p8�/K��2_\Q؋r�-+V����˙�:��CJ�7r{���~�p(=� �=����p�R������\C����Z{22ᗮ��v���V�89���p:��)���D��Os�k&���$��ʳ�#z����²*��am|�WН7zp*_r������,��4J���7���K3�NK�);�q��c9�7�<�y=g��r�I[�R$�xڀ'\�2�ȡC�A�k���ZkYep]J��2m(p��r�2�*����hd�3�Tq��Zޫ��:�y����Nb��!ozfd��Y��NV�ves+�#����2��O�>#��('}�]�}�v���0YJ��ۺ��u�� �|%kV�!gU�u�c�|��U�k�֡(L�*��^��lP���{�٢�z¤�*����~�w9#���P��8�A��vey���3�3#d͔b6�i�����=׼�S�7����Ѱ�l����q��S���ټn�V�X+�Ԡ�Bᓃ���wr^:�҄���n����lG7:T�/C2�|U�Ľk�5V8J�_%J��	���}5b�
���z�(@�WY�r�& �s�-�e�+z�Y���;'����u���|�uAn�y`�;9�M�AJ�|$8����^��G@��BP�+���5\��?�������2�,�˘n1�%:.�A۬1��ZfM�V�f�Z��I��ڭ�:�72�ƻ��K;��T�|�6��>N@r�{�;�V�޴���b���9�VnE8^�IS��;9%���=���4.��S;���6�g7WfT�%��EY����Ք>������(��n J�e��/M@��M%��y[��a�mV�8�q���z��-U�Jݘp�e�N6�:�o/��hQW���k�T�����#t)�;;�~Ԕ�7"�ʼ�hMU�y޺]+��j�q�]����fK�`�]@"V:]��PPu�����%�wa@	}O�A��(�T�����'j�M<���$Z(Gt_e���f����,Y'��y�m;���7w�E,	=�Z��U�h�,]&�a������Xh�$PÝ��e�t�L���]�D�Ś�Q0�@^:��-���pb:�� n�3��M|���UB�c��u�۱�1f��𡁴�κy�n��w�7��8�m�oy:����-������d�5����1�q���j��Ȱ�Z{9.�SY���	��e�
�H�&�>�#O2�>��l��	R�M�e��[��h��9�kϨS�������q��W�ή���]ބM��wv*�V��E��'E�j�{2�/.5�	>�(R݇P��U���6!���Ԓ�w�[׬�y
(��ij�ݴ���a!{q�8
��er��>,k�r�va�+ȯ�t��8�d�Eβ���B#�at6�qJ�(���1e-x�_*`�w��/�9y�\�fLf�b�⽮L��k�x[2L��{	��Uo�h���⫸����m`�,|�VR�� ���������v���e��pcr�C�s[_ �v|WGWv����P���Yż�<��b-�K�WO�f����:^X�Q	vj&��3���oea�>8jV�y|����	�V��Ŏ�������Q�"��i�:.j~�G/;I�>����$(H�L)�1@́Ntbs�%�d����`4��Ή��΅�)J@� I�2lM��c(����(1F���Y�")� �.�Hbh��"F&�iL�P!C�$���2̊�dQ�%��`�2�.��F��A@��Q$��c���H�M����LFE2c(���bP&�c"�a����л��d�Lb\�]�E	Dh\� %%0 �����(����ˤ���Nu4EI���Ɉ���h��23:���2"QT�1r�J�"�h ��E�э�	�(#3�����(&m)L�H�������y?e{U��౵���?+��t��;{<.qw������LD�y�Ѣ���}ԕ��V_$+�N�3/�e'/.Z[o���?�5?,�w
ZL^������ҙ*��.��ͬmj��X�V��p'�ju,���B�K��_p�0�����)�b���6)nVU�e���.��1"6XR�5��f��}ڝ����Y�]ȿ�u�}�|��]�uoޙ���vuQ�D��de������#n`���!��{�zj{o�"urx�*��J��㻺f���=��O���}�df��n�ٙP(=#���[����<�mR\*n�{i�J��8��U���P�q�������/Hɚޟ�A��Q�C����^�?>�`�����{<P�ڵ�N�SOLg��+�s��W��߫p��㓟�g�J����=�2k<��x�2�9Q��Qb��R�����|�<�뀥����23q��Í�m����1TU��-���H>'W���}W���t�+������"�y{ d�������<��{De���<˟=��G��{_]3�g	H��za�z����Ս��k��M^��$��,���ɲK�n��.�u��
���]i��V�����=��̠�����B�t[�e>���3��/�'�|��Omh3�U��U]Qp� |�[����NV���u�|�z�wĉ�K�ʳ'%�/�YK�m���P�g�^z)_��ȟm�p���*(����ʨwF|��3o��u�LN����o���}�|�%���~S��^��;%�C�	*���&�C���nc�"�a��t���3�-�^���dКz�������I��j�|=9��:tK7	ў{��Sw�s=�f��|�������L�9v�t:v������w�):U�}q;q��a�������J�ddN�Z��gwc�B<g�� � W�Jjk :�o����Θ~������q7����~���9ׇI�[��ZQ5^���jt�" 5B@�?��7E����ioYw�����"}`:�\��eu��Q�l��[7NF��r��u�"��W�n�Z6H�}^�t_���~+��y��:��F��>�bH��>�>�������ր�u�w�U����L�)���ة}Z*��~;D�Vw�g=Z'/3�mvÛ;�*7м���c��d�����C5Co��"����|n|���g�w=(���mw���ܥ|�����5HU�5�.���r���~�������z�m�ޡ�l�q�+8l�1�߉��yӭ��}f��׫�*%���W���h^�8+��͘D&Z�Z�^=�,���v-ټ�c���%U�=��·�0��n�'fJ�s��x��[f��Gl*�f���[q��ފU���0Sǡ�!��O%n��L<`Plh�<N���RR�K�^�����_��t�I��C��x�U���~��9���o�(9�`F���,O��;@����i
��3����fcʄ���Y^�t�A��`	���lg�*��9׻��)��}Xv��2yD��}����ʡ��'v��<4|��Ui����m0B֬�F��ɓ�'s*{���+��q��>~��z.����sX���U���k���TC��gt���נ���{�VGovn�u�>��}�z����P�y�y\wg�����o�u)J%�Bg����w,�ovwg���ǫd{���-@�T�Y~>�L�����"�F���4�E� ���jf��z��evh3��T��2Zs��h:}�����1�u�P��]o�z���hM�~�3�s����f�$����fIA{�<�B�?^����+~�{�aݕ��	��UsO��T+�&��{}p���>6Ȁ�A����J�U�a�[�Mb9�)��N��Y���*�,�Dy�M�}R:�wlU��T�m���A#��[���a���W�m��g��fφ�wLc�~t�4\Y��7�1爕}�+.��\)�~y�MN�1k���"��닎J'���Iԕf@�+5�TW�.U�z.�F���!"���C;�q	����e�RV�یB�e�<�ӷ���]\ꛧ�� J]���
6@GU>i�'r�#�W�i��������ǧ�A���|�oƶUIb�Ijn	��P�����f��묯{w�9O����j!o
�pڿI����'�=3�'��h�~$k��Q���f˕w�:��9位-��h�K�i�u����ϴ�wz�v������6�>��ϡ���� <=�0�6�խ���~1�b{-������ciu�3���^?P�����n]��P�w�y��׍z6Ͼ���
r�Uf=�'tø�V鸢������t��U^���mk!W�L����+^���(�頧g�?M��{7(ft�����n}�C�p�^5~����7�[%��r�w;��T������	Y���p���ulL�4}:�eV��@H>�kq��w{�֒��=>�QR�y.ix���[��ێX�x�9���xKk3���8�<�ߣ;2۝矸g���X��	M���ua/Z��2���7ޭFѾ}t�|+���~��T�ܥjP��|g�P3���#qNC*�l��u t-g��Y�?�^�<����H��7��� 3A��֜������{���If�����m���i�]i�����r�=��Ŵ��܍%��%���w�5�!p���kE�9�9������SZ�l��N�3I��gm��e��ۡvT(�騮��X�qld�L���n��5��0��Ǒ�*�������O�yty��������U^�f��ԧ]gr��Y~}|���ϸ�nD�Fc�O�ʡ��e�u2���x������&=��W��Rp�}���9��Q��S#;��dq�%�9 '$p��ٲ��c���Ͻݽ����G޷늸t�#�C����'/o�F����~��nE�� w��=#,�v�q�c={���:tW��[���[f<s�̿L��q�z�z�w~4.UK8qY�^ŗO=]��\���	H/�к�����]���m��c=>V|s�;�^G�F�qX�#[���vJJ&��y�רڙ#�Q��uz��kf�#e�.TC�&��\6������g�ɹkl��ɯh~������'��7�2<��ϥ�n��+��鯗{o�og���E�y�3�3i/.��}�y�����8��}�ہKՆe\a��>�ô^�q)��Ч}3������gж��s����P�y�	����/Hɚޟ�}'�F�W{Ϊ�i��/��3�'*;��c{æ�p���µ��yf��%k�V��*Y�cؒ��M�z�Zӗ��ߨ�UwK�c�+���K��i�Cr9qYd�=�������f�S:U�j�=7\ ȝ�Qr�\��*ť�:\]\�����M���.��y�hT�'h�>��o��l�v�~:��x�>��Wx����V~�}��ߧ<kN3����Edň+%�/е+/{᳁��9GE�t�v�S�|�<2%��@�~���zhodk��5�lw�*/U�5ݫ�f�I
��q�#��٘yBZ,_ՓZn���,Z�.W��DK�?Kq�;�|�`s����,�J�z�Y�{���o���d��aᯌ�C��R7����]��<�sEI��綨V�o4oI�v�z�L7��C�dK�B����Yr�(�Ih��E�2�ɥ�\]�/ۧ�}]N��M.t�a�r��=�|}�����NW�x,�^�"N�wP$��g���P���+�C��6�_������rZ?��К����yI�|s�'ǯ�j�}�վ>�ӢY�p@Nǹم�3~�۱غ���eP
��.�}�NC�Z*�Ӵ47����IҮ=����]�0�۵4���w�w���Q`�x�`�����zW��|K}|<3��lgޝ�����q;T#�����Mힾ��*.&���۸��SS�h�T$W���|}�&[�C�R����]��y�-�H��e`�ק�mV�����"���ƭk3��n�l�O%��lN�k͓y,�$TeP����o��;@��Қ�T�D�e�w�z��3o�z�8;�\�x܇�ЕhM�l�Һ��J�+����:�u���u�Z<�����D�?z���g�*�Uz��%�pH9�z���+&���r+���n�g.��$8���O��ԁ�G�x��f�
~��7��T���G�ˀ۬�;g�y�xW���H�ӻ���:;���ܕT��R�L�{��3T6�CH����s������]�?�K.���i�q]��Z^]yp���F�EzNx��z�m�z���^��9��ǝ����C��{	��󱵡_�+N��N�����/n�1�}�
5����o��ez�u�~���uE>FrY�F{/.���s:�U��ⲽ���:�� Mg��ȕN���o��C���u�9��c�.Z2��k����Z8Ne����G]t�(xM�b� ����s�b��t�O*���#��6FO��|�}�!{��:�+.p�4�g>�=P�+�H���=�h��3��^nx{`Z>=>�j�*9:^>���p�VDW��vDy�1~s������&XW��2��û�����Ve�<�0�3ޘ��!�|gŨ�Qh��}��y�y�yau���\i�:ٌ�����b���0�mHwz��㢺�tv�շdQ��{��3�6�r��j�\��y��h~\x���N�-rez<j��8�#6�Q�!��j��Ndk)'�]�]أ�"����sb�.�)�q3�]��p��n�Ĥ�k�n�gf��%�#cE���lH��z� ��S�B�|��ɠ��}��ўC��������;�w{��}�ދ`��[}����5֌?@ݩ�Q'�g��"EKfIA{����V�>�2�u���ugW+�O�=���������ɟn�@�-��~<�B���j�n���
Q�ܭ~�x��Ӵ��~�8�o�F�����U>�d�5�2[��/O�׺)$r�.���.�N�#�d�k߽m��L�x�zz�{ՠtz�<i�̖5T���$�}/�����_g^��I\�B�9�F�L���^����'�=3�'��5�?M�����F��6˿8b�a�����!�|=V*vy��Zj�e����Wra��2_����3Q��c9��
˧0��>���W�=r�EEK�Oa��|��K>�]����gܽw"����Ne�K��o�ok��K�ќ�� 9�nEi�8ځ],�a���0���n������4^��u�}�'T���JѮ�B������������ܡ�|Np8<��ݨwY^F�'I���{�|�{�g*'s��gq�:k�\zP���0w�~�����Hx+U�@��^��E��g���<����scm+� UσV�k{M�⚤PJ���\�ՙ�6�Q�ٌ9i�5�-�s7	��$^ #j���05�_u�Z��i������ĕ���@ӛmvrչ�>�Z�2}T��n�;�#�U�+#}٢��+h�)�t����P}:�yT�v�W{Wj��g�|�f�ʁKZ��fW��q�����r�[Ʊ϶��C�:w��)k�����@�wg��ia���	�Ԫ:'�5#���P^��>�t�YO����|�s�.xQ�s��ǪH�R>���\c* ��u3�e���C� k����������9V���Y�����BX+����ſ>���(���#�U1u2�������a��y;��\C��N�=T\�K����.RGjt��VO�;E�e]|f:��rfIAx�g�&�;ytA��Z�R�ٙ��t�i��>s����������~ϸΒ��9�<��&�r��ڄ]����v!^�>��#��;N��N�8�w�q����W�\����V�?L���"������鷛��Y�<xWT
�S�+ ƾ[����6aǧz�����o�������hi���g��*�̮�}<}�$r� t�>jh\E9�Ȁ|B޲�ڿ3�O���L�uw�lVֻ�N�1v'����j�LoiF#��[m3c�s�G������J�&��?����o���G��m[N2�l�ܫ�0{V�P�
��Rq#'8Z� ׸k��f���͕:����ne1.˨����syR9æ�s*W[R�Zr����SB�s�]nʊ�F��X��/��d5�[,z�+!�M]ț� ��5Q�9~{�95���N0Pب���^���FG���9�wF_�^W����0���^��3^Ww-�8�y'W&�3ޠ=>�x>`���z6�R�a�P(>;g��n�(v�5�$G�}���7�G���p����괭~�=&��]xOg�����z�����k��K����N���n�7�>�~��hۊ�i:n4����뇑*k�c!�Ew�F���V}�~�����kp��o�P���dM]��;]�k���'{᳣�rN���>'WK��q����@ϥ����23F�;�U}C���ZY�R1�?nm�9:N�0�>�/�ɭ2�]i�_-v�yz�\=�;����zL��ŷNl����W��~�A}�}t�Y�R�3A��s�v)�_�j�����}�v��v�g<��rR�MS�z�hx,����ڠ�\�J5%�FUC�3�d������ݽy���@�/�X~���s�'�۞��9�^��;%��%t� ���w���s��^ň��0:���#m��a�3��^�&�����.�5�}�\�C��8��s�.�Y���r�/cH�t��`9���|ë�y#Zƙ����m�4h\����]j�K�����R��:���(���뜏y<!v�>�	mB����w�e�ԥ��U�ֵZ���i�]��S2]v0=mР��,�d�]͝�讅:⠵�I1ު��P��<Y�C�n���6X/�X޿�	B-�O��ޫX�Q�-�f�őD�l�*���
|~�E
����_�5�R�S�Hs��.e��o34����k<3|{#p$5/P��Z �n��+����*���d���oL�����$���cLΖ`��# D�h�#%evK�*@ܨ�:0�n�P��.W���k�a�˨fI���ސ�.Ju���2E�4I����^���3Uc�$g
Ĭ1w�]�JP,V�u#æ���*Nw����lԈ�m��D,�X�]�W�u��j;Ri�i��=Gs�ln�B�̦��_�8���2�es.�UJٲ���J�:I|������Pˀ�@����-jv= _�a�p�_�2,�*�!w�YD�n���]_n�.�b�"�I�1[sǸ�:��{N8��#f5��\�<B�l�����h=�b�]Ki`Z�c��O�Ww.�pϊ�0�Euv��+h������&�ھ����l{�JۂI��o �6^�[�܉��*�����p0���1��])jgf�)�$h�qS��&!zD�Y0��ق_3�+O��=r�Y�`�a��{\~}h�{�߶�4�kWmp�����Sۂ��}���ѣq�gܱS.R���0v��7�l&S��M�ur=�k�c�A�h= i���i�ރI �vn��	ci�e�C���j��Ž�,��Vn�R��i���ͯ�5��-���3�v�1�3sZ!�z�<�Bs�*af�u���5�-^[!;(y�#�z���ư���Ύ�=�_	��a����,��gWZ�J̹6��bSK޹�qR�l<��d"�;����v&�-�]�C U�w��`E��=[}2�e��V�ʒ�q7[����}vol�&��0�ekKy*l�ko��4���{���N�.����v��+1T�in�B�Ի]��i�4U��,tӱj<��53������;#3����d�q�yZ�(v1¸��s�K����egkn���[�,{��K��cK�\k�-Yi��h�WpƊ�=�WJ��#+p�ֺ�-�f%�M��d�y�̥��,ǭA��Œt3��0T�'& ט�/�L����շ7PhB�Ϳ��+��]Q��֐�͵�,��
���NK���C}0u2 z#��[�k�MYІ]�7N��ĪT{�nTK�%湕�q�<�1pNR���)�O��$;-��!k�58�o����:㴟	;���	��?G�"I��2�@�˩D�+�4F��%���2L�F��h�R)	 ���Q���hj$k��L�L� A�wwq0d��Hd�"ə$��0I6	0 ���(�����M�2"`��H͑0`F&X�͒ŉ
wu7+���s32�D��q	$��D
d��cwp�"D&BfE�$D\���D�(��IIaэ�	BdȦ�.$���#H�b`ȈL ��fB'.�ђ�P��Ĉ���A�y����B��)���C ��<��Aڦ��r�lw6�a<綝<���+�H�YJ�����eo*��3E x��}9��T��ޘ����<�KU��#�O���'�T{U��>���@��,��*��xȸ|fj]��B<�D�#���/L]L��ǎ�U�v��o�m�_���6��]�w*��ݨ�5�F��Op@N��� �@�Ҽ��:���xz|�����n��˘�>"%�{��o������+���Ek��e�� p���]F�>�R���kș��ނ��9��Hٜly�R'����W�\S��T��%�q�c�}^�t_���lI�6߱l�nǢl���*��I���Hdx׀�k@~��.f�S
��Ɓ1��
&�%\�zw���~B��9G�^�����{>M�ɸ�/���� o���CH�^��;W��\Q�z�ܵ��[�;�8=%���W��+Kð����ܽw�3_��&����޺�/5���s{�ք�b}}�!>g�O{�0����}�Eӝ'n6P�^��c#�{�3_�/O����
���<��	��}�g}��]S;|N���*�a�e{��9�v��b��l$@!�r��yS,Kޛ���P@ڳ-óVQ�ձ�kp���)V$�n�/(ߟ�5��t� �Y�5
�t�U/n��z���jJ�~�G��?!q M�k���u3�5��u뮭��c`�O�w��f��x뀫3�ӕ�|�}t��vj�8}��Jk�`6���|�Nv�ijK&t���|�d{zWyV��f��s�������T;���qE��^�}�u@�13��js��� Z��z��.|3�*=�!{��:�+"�	Cne�=P�^�O����ȟn�ݺ��V�Z��G@\F�ъ@�'K�ձ�~+"��;�ϱ��:�(R$����Y��i?���y������	����t��9	����\w�C�,��ޗ�Σܾ.��2p��N:}��{(՟}jH>�<�
E��T���s�<�����FyS����W�bM���N�^k:�Z�X��0�;jY�Q%��_��H����q2��<y���~�7}*�ɵƯ3�\p[�)�8y��>�~�\{mO�� &t�-���^*������)��4�z��v���gL��W�t�xdG�k���ԇ~�T��U1Z�U>�d�4H�?�����3��V������Y�Ǽ^��C~��zgx��}=Z��z���~.�ʹ|9�F=�3e���n�{�׫֫��Ýh����tn�io
�6��}��O���;�|����g�&o9���0����%AS�w�12�]GA�ٴ��7w��HK�n��d����Ɍ����M�p��XVk�P㆝g3�}=f���f�v_3܋\���'����qk��Ly[]n��J�!�W�3qF����PǕ�,t��Xܜ��յ,�[jw��I��2F�t�,���zV�������CMUI�m�̛����������W��v��'s��z&=졄
o)QX.c���b���N}��e���]�c���_>�tMaP�S^�Zb�}R�<�q8w�P+�Ī�l��;��z�M�z}�Lh�R�eW���4��V�%Ug�	L�>�z���Fz�zzr=�ֽ��3:|N�@8=J��;?C�rPH^>�_�F��_����|j���ȕT����ür;�^���{j�ߙ�7����܂�j�	�=���޳�3�}^�f�D�4������ �>g�����!z���9F��Prg��׽>�C<t�D���EK�����;,c]���k�D�L����J^md�[�'s����M�!^�1����G",�)_�g�*�,I>Gb��U�١�5�KY��W��Z����V��t�l�Y�Euxya�j1qϮ�r,�J�1�hʦ.�R3'�>ytm`[���f��B�2�=�*4�~�܈�Q�z���/i�$��X1�*�qF[/�h�o%�yCst
�����z�<�+�9���^�άf	a�����
���b�uՋz����]��j��r��Vn�f�.̛\�<����mD{O��Ӯ05�����|�V.�m��8��6�в�ר]���%�=ٞ8���y���H��ud�v.��/�;���S�����g����j�p�w���:K����8�Ī��Z������eM=�J������Q��7��qV��G>s;��'J�o�F�z�٫~��yzy7w<DP=k7{<R��z&@逺�P)�P��[����z�1�zw���ޙ�&��\OtF[>�v=�.�{w�ZQ>�4=ꪝ6�Hjā�
��x�P���pڿ<|�������C�^ٹ�7����j�:N11�=�x�*��רڙ!��OY����7E����=K���R�|}�>Ž�)���F�D�y{����ϙ��)�2�W��~�q��#�c%�n���v�n�~^�[�����tz*ϻV��5%}������}�����p)z�̫�l>7g��J���~U]�ӊ��+2�︭5{yq섽w�5�����]xOg�t9z�]�w�wRB�Ɨ��~��_�������8���뇒���3���9�����n�5O����}���I
�a�}����-����NQ�t���}{���{ g��{�;��멽��.���7V��3��8�uI
�Ë8�[���U#�?P�����9��2��ݾ�lw�RK�W�My�Y�����vvP�چNۖ�8��yF����H�q"���֫t��K�;�u)�ä�8��
e��r�c���0��n33���*�1;�ߞ��_�n3��;��yB|�Y5��)�Q���Z�;�V�u\6�o���_���Rn^�W���{����hY)w�aᯠ�T9��;���S��<��H����K3)�a� /P�R���"�LyO�_K�B����Y(��D��|eT?]B{�M�x���wb�}v�_L���{��c�u���^R}�d��r�%G����W��{�g���=UGI>�ğJe��KU��"<���9����P�zs��(;<�s��}�u��5�lzDѸ r��x	
P4nb�S���Z*�;CC{�|_�Rt��[��߸�zf}���4�ڝ�N�S��1��O��8 'Pd�[ +�k�c���xgޯ;aF&�;v{ƻ�M�����S�/�����}Q:}U�p�jY�D@j���/OQ�/��>P����W�=����̟C��w���"}�3���{ޮ�Y슷U^��FIh� }^�^~�N������[Y��9�|t�z#j;ƾ\�C���O��@��XZ�z��ê�T�$�Ng���//���<47ؔᵆ�3yI��"�R��0K�y���KM�旡���`^nҮ $��u�����k<���R�����V<t�	�wuwq�src��Fb�7�8sp�&�"�</���>�^�uU��Oc3�]��g�c��S�gR�I��߱��{a��T7	��8��2T{ޠ;�L���P�2\���q��R�r٬]�{~�U��σ�6�R��{^���ח9z�g���9��]��ӌ�㢪��>���o�/��l�2�Q�<�և'�pm9�v�P�^��c>�^�W�.���������1�>�fVo�(W�חL�q�;�f<��{��7�9�we�1������6d�h�N=�]�fw�=�^���^�NGzh{����Z7וC�s8�<4|��Ui9�ū�a� J��={��Ws��i+�� *�d�x�.�7�}����S�{�8Js/3q��T�x�Vfr�J�g��U�qG�$l�
ƺ�:^>���p�T�Tn��c�]E
�[�z�#��s��^+R��'}���t)'�c��!9��^/z�W�h��r#ޗ��������P���J�w½v}�{eq�rԐUD�$"��R���'.̇O}~=C���B��(�y�ϱr��>6o���au�1��RͲ�,�H�_Kf�P^Ǐ4PV�y�=Q�t�E������R~�`y�L�/ݲ�Z'{����Ų):b����|ul�	�ү.�3b.͍�m��ݺz<�rī{H:���z�<QA-����Gf�.�%��5+�v���-+sB�yv�!!��K�1��+h��<��z��O��Uv���8�y��̭�*:U�i	�q��`��`@O��t	-���^*�I]�)�1G&�������T���W�5�g�v��o�Hq7��H�]�o�S�d���"�T���t�������o����1�5xT;���s�;��>;8G���.=U�5n������F�|*\M��Ž��@x�  �;�
��qѸ�[¡�6��}��O��L��C5�L�S�ד8�*��=��)��G�ez���<�����
+Ҵ����]ޢ�j�L6�FO���f���|'�P឵�j�Y�M� U�1��n����.c���=�[X6��M^�K��0�������u}��3{�.��s�<��)���|��ñލ�>%F�}���};�b�����3+�/#ʯw{}��cж��d/U>:�#�o�A��fF�!{7(fGO�ڀpy;��wA̯k�ܟ%�t�2;I����7����J�zNCu��9ު𕑾��o�[GQ�p�	�jF�й��^�Q�+>�>;8�YU���̔o�ˁ_-���@���+}�吽|�G݇b�tp~� ��kۀol�S�:Ƶ �勮�<;�5xÀɋ�I����I�Ț���:܁[�F9}�1pq;3k:��Ĵ9�3�!����-4t��q�Ѿ*�e��e\b��G.9b�� Oɸd���-��7W85*y;x��;�t��A��e��謢����%��R��r<�i`(�P;�]��.�+ӮQ�Sv],Q傫ѷ���1q�}t�E�%+�� �c"�|��NC*��,� ��$���Xq;�R��K�{�oI9���l����Q֣�����Tf<�T��S)�*��:�^�o���f7�wKܺ������u����q�{H<���f�e]A���a�#��U׳�wb��$�h��ۊ�N��<���g��#�oڪF�?]�{#��.܀�<�Y�s/�^�P�nq���:}�qFB�q�T;�t�"���{�t����o�i���>|�h�Jז�<="x����P(~�+"|j�py�m��N����d}ؒ��*�N	���0����ŏy������@j�g���f�1��d+�%l1���t mGR�=�_�^:}��O�����~��&}EB�!�=F2"_W��Qkf�e�*s1KAS6��(�w-����0-UR<����<g�w����.�/]z�FG���Q_O���Q��ϧ����b�n��EK��A
����ӞV_l���^z�#�H8,�Y)��J� .�.Ȏ.�]0�5w}�U�S����I�y�ud��Eݬ�Χ:#�R��r������+��)��!�U(%��;z��A��k��&[�u���b�.}����|���+�55%������i�fhoz2�o�Նe@���V��j����	L�4�Z��^ђ�0��i�����{yp��w�>���n3�^���t:�z���*i��[�d֗N�j=��;V��>���V6tu�exl�i8p/�چ��5�1��+�s}U�+�L�C>���g��9+���~��5�<�'�h����J����W
]/d
�p�8]�_gl�h����fFn:�c�V�3��٘yP'ȱu�Zo�r�l��O�;,E8�*�\��4�JMd��y�^�z�o������r��0�ឨw^�G��=+��Pn�����3�Z��/T'+ޚq~�<��hx"����Ae�$�RZ'�M�=w>�¹ ���R������d(��,(�K���I���G���L�χ/���t엷���k��U.�%�>Eo!�	;��#�0�鎩�&q�К�����O����|z�ڮD���Vb����J%�/�gD�ߠ��FxE@>nb�S��s��Ӵ4c}�h��t��xVh7]�>
�&�R�=`��/hmj��&;��R����ï�Fc�<J����z�	�מu��7�kPc�� �25����r�Z��NU�m>��v�\�s2��anV�C�������9V�LdT��w�ap�H���n�R9,�|�\Nۻ�q�����0@����yM`,uB�_���1���隝������:��zuZ�=��=Q:}���[��f�D@j�H'�]F�>׀ƅ=�|]J9�Ow��G�ϣ�b߼����>��&���p��dU���M�$�n �:y:��?LK)�e﫵%s�T}��F�&W!0����O��@���^ w������U������¨���׫�� �G���6*w�E]K��:���p�7w'~&J�{�y�����U��-)|������{絃ԧ>�r���NqR��{^l�5��ˇ��Za}��^�3�)�����l���L#��� �{n�ߝ3g�%E�|�ևu>Ӣ��;q���/n�0��!%w0�;���.��Q�+���A9��[��uL��|N�1�'tø��q�P=�t?ߟ�C:�d�L��k�� |�p���w��7^�NGzh{���p(�f�Ϝ�;�ó�||��f�����vg���[��_�>���*�� R֬����^ ���t�{k���/|먬��P��"���
/=���]�ր�~�A���z�G8�*�/zr�T�4�b:u����ch=��d��]W��2�g��&�ѦZŻ(K���xv�iCw�SP��H�;+��޼���o�熵f-dt�z�����2�f�o�ci��"n��y�9�y�+wo`�,1�P�f&nu%oH�l��C�_M�e
�&��S�V�wG���¶a�<���K��()ox�R����nҦ���E���<��<^aBDٹP�])*wZ�xRnؙ����� �3R�J�ɖ)]���C&���x)^�&��~j���v���ޜ�mq�}���)ɰ���1h��]vT+A�Q���(J������DR`��QD�Iۘ� ��E��p�l�1�6�)�����t��b�����߹>m�ua0H���IL����h�΢���V�-����a.1��m��a5��5��~����|i�Qx�2�Jm�pr��}7*g�j���Y���YkMx���{��f'Z��0�DL��Kq������'Zg�X[���n�ڥ��bV��:��R��f��q�st��-F�:������.�S�^�R�>}I��=f�R��/vKx]Wp��{�;Z�"vM�U�0%���n��.7g��Z*�z�V;��"YG�kA̛�����j�Sq���r;��#�4�a�O�rH�-�F��ɩ�-�FGE��	�}Cz��o5��%k/֧c�*lMN�0��F�k�*@��w[�nƃ����dV1�nn�a��B&1D�&FĻC���p��u��<��Վ���$��T�Q 9���Mk9v����w�[׵i�\�X7�4��Lx���^�{Y�%�i�0�<:J���Y�w+]�J�
U[[��X.�2ҳ�^��ۍ������b����t=��P􉶥Z0��`�u�uq^?7Ef�n���"�0c��c������twY�����ԷZ�z�̈́Q���������=��Ç��K��W��7�}1}�J�Qp��tg6�nf���v	�̓zA��a�G����M������֊�ϲ��o�8Gwftsг�c���{(ݐ݃]$4��#�ݾ�H�{�ꌛ����Ӳ�'DԸ]�s������w�Z��#&�����o5�3+%�L�,{�8E�Θryx'�Ϯ���X�w�7=s{�<�ХZvkX�9�A��]�7��[E�,��]Zt�#5cT�/E�x�fJpN��Ht�G}�4oL�k1]�����NG"::���x���O����1/$ץ�B�/Wӳ�S�g�2e�tq�{5,�q��2b���ׂ����݄=�4�l{ō�%e�K>3en�\Sh.�Lٯm*x��&)��	�o��!w	:�i]���b�j�]��6�c�QswB6��u�
�xr�CN�M{�s33�:8�ꝧ���_I��� ���%FdBY&"�A�t�r�$�je&,&(
l��
!1
D��#1�1��$L(d�9\�h�Lhs��3D�F�IƂd���;�Ldis���(13fQID�!��2���I1D�`�#	4����ɣ(����0�E	�%����id�dę�cd幒��"1!FL�fC{nTl��(AM���4�ܮ;��KH��F&�v+�^.W8��ɢwvD,c)d)9r���DFLd�x��SL�x�$ئ���;��� I
��$?�b��d�e��o]��	L{��+/QV�,M�O>��D�T�Lӵ4��i��-B�s��l�@ƛ���X�$?�C?��\n��4F�@\5��/Vǲ������H�z?[� ���`�y�ջd��P�6��$�T�
�<=Tϔ��9	�����@{%��ޗ�rtD�t�Փ;O1��K��[�V2q�G�W�ȵ$Fx	��,]J�.�|��ɠ��{<4+y�ދ9�Uݙ�������:��{��|c�;jY�e]|g���"��[72����z=�b����0��Z�v�ϴP�F?uy��'/m!:o���>6Ȁ�A��� N��T[N�_����>����@�����}����5�g�v��o�Hq7��H��ݱV�U>�d�5���շ�
������^���'f�L��&[¡�~��}��>�ߣ�ՠ߽��/�Y�[9����/[��M�s���?V4g+�@���>�C�s���B��m_���ȟ��>�Q-��l����:�cU��eb$[��F��X�Y�^���e�����Wrc߫c}�k��=4�X��^2^�[��C���+ \Ǖ����ތ�>�ZX�TU�<�V�{uU�G����fyy`��æ4��oD,ܜ��G��hm�u|�苡�v�RF�)�r7�sZ�;%��6�X5��en�x3�\��]'T���t:i�h��n�E�/w�x��[9.��LC�Vm]�q�.�BEO,��"�<�}u�ެ�,�3���rW6^���܋�z��oޟ yz�p���ځQ��U�}qwL9����C�����Vn��;�ǟ�*����Ԫ��_�x����������Z�nP���;P#S���p�`]����s9t�z.\�Q����O�ok����T����ür#�U�+}����+h�;<,�{Ɓ��'л_O�8W�wGG��p���%�K�K|�=�.ix��/վ+}��5C����m��\�!~�2q��q�{g5���;i~���5�����VvX
5��/Z�鋽����<�m(]��g=�?\od{����]#B�K�2�T@3ŋ��#t�2�l�������B6��^��|�l@I��)�_�:�!�]j1qϮ�s�(��Ǒ��ʦ.�R>οn���@ї��[��1�_����C��~���O�w=�G���c�r^�>�,�(�����v�%y�~��Y�}b�Vg7�~� �d�	CǷp�ߴ�y����Q�{UH�~���Dq�%�* /=�Iyv־�\��$��*��v"����޸��N�8�w�q����^��-�׶V�UY���J�.�6�����P�M�f�7y������������齌wN;�?38����3jt�;:a-���i������(���]r�."J�25�.��;��&���{�� �D��bh�$�-�nn�x��q�H�[�tY� ��wz�X�{4'Ofu��Nq(m�W�a���fg}D"�&@��7P s��]�/�ޞϩ#�N����;q�e���[Λ��>����+z�w��١n�����IX�:�N{�r _B޲N^=���xrس̓�3�y�+>>'<K����+ͧ��$�t
Y���n��jk���+��S���^ݏH�v�#���6���#�|{!���~�����7��#�\])���|�=����/���#�4�4��������������4�346��F�
^�3+�،C����;+�AS���p�Q��q�/M^�\<�/]����^z��{#޺}�|Gx�Ꙩ�>�o5vbHO�̯zxjO����ӓ�/Iӡx�^�\<�T״�C~��U�ڙg�q˺�"��|*Z��h����G�9�֖?���i��*r���S�������,����&ab	џ>溶�o�z|�Q�顽����/��m�gIݸ3(O�b�kM�N@��>�j�>~�:UH$V]����.v��/d�u��{�z�o{e�}t�% a�Pg���'#�fݚ^��]sxe�������N�mJ�fsQ��7O�y��V�wpËÕ���&r0f�1ī�e:�h�{pF��֧��l��i8��1����b68ɤ>&�a������绬Fn�M�?�_}�==��֎�Ur��L=�2.�x0����7'�w���@��,����{�[�c�+և�/)���Ba��Kz�[�'��94���o]���/��p/�Xk�ޯa���{���yׂ/)�ͦf����>����Ҡ=2k
��BU�[���Rg!�КZ��9R|_�I����3W� 3����n��[�W�;[����Â`�J���I)�y�p���{��=G�9�v�.82����N�~�\N߮�q��p �" ���o��%���$`�y�.Y�R}�ǝ7~��z�;ޞ�W�����~��u5,�" 5B@�0W����ɛDñ��ы�3>1�&�Wv���|t��L{�������J'��tx���\�z��:��M�2KF�	W�|�>>7[��k�*�<��m�<����f�r�M_��ޔ��5�{�����,�Y#�.rW�U]���̟MTǲd���zlT��E]O�v��zk��m���ܛ��&��P�|�y�e�Պ�ez/��Su�Ӝ7>
�c���h�T}���[��z&���ߒ��g���uo�r�m����6�����K�Ս�R줎X�;��0�w(IQ��EH��,Xͻ"	�Y��N��-��,�7-e���d�˴�-а���S��u���DX��(��C���|v<�W֐�:,�.V�΂p��ym��3f�".��U~� �~�q�f���5�kC��<z�+~W�ߞ�2�_����
�W5ug�!���Fo�Azs}5�+7�)�����wnǕ@��ⲽ�gkί|F>.��٫����A�GW�Y�hd�w��u�����oN����m�܈s���+l.��ͩW����Vu�z�T��H�ci��D��T�������/u�q�u�Ttq��9d5��=��ya<;g�v��N����y����r�'K����{����a~QxH����w�����;G��I%TL�('�ȩ�)�������w�=���2��N�|Щۺ�f�c��Y�Ew\5�Z���q�s�RAUx	�"�ԪB���Cɠ�*����z��)���� ��Ô3��>=~��au�1��,�̢K��<����rb�u��c�L�n������tݱ~C�ۼ=�~�}^elyQҮ#�HN����q��>7�"`�@F_�ev�[G�;(���*�=�R����_-}qW��;^G�=�C�����uǮ튷����؍[�U`ng�+���݋�Ux�N�ŀ��tS=Z:�`������U��9
�����֖,���Ռ��&�]C���<��\�V�{%Z��s���ޔ��͗�P�Ϭ*C5k��{��\�RAg]&�˘����Me苴vqT�S�E���f]��H̃�� qf�����L>+xL>��m���;��;���n#��������ݫ���gv���O��)���ЪKSd���~�*K�6>����^����'ĺ��m��9sw;��yeM9�s�5�TCu��m����D{�&2�yOŅ�����\��o�\�Dz���NZ��7Z'�&=��+2o�����z�+�^��c˄��koFS�i�����8
��3z���wC᝕V0z�܌~���������F�
��*��>�;��c���n����8����-�(`轼�2!*�q��3~�v}�M��ܡ�|Nmﻙz:���g/t=Jϐ�>=�Ⲽ�����/Ưo���UOIϛ����UxJȍ�f�<�j�<�V���B��E�΃�ng�j ��M�^%9.-��D���~��� 8���ߧvof��l�N;=�\�u�Y�A��t�>�����΋��yM�������Q�qj�bR���mY�}�`z'��Y�\od{�����}t�%.�,e<X��g��S��Q)�[*�mվ��RT�~c�u����ư�ז�Z�Ł�p���Tڋ��Z]�%�����9N�1@�]�g�iƎ[ݽ�S�;5smC%�+�
:�Aev���u��=2�Ͷ�X��V�V��]��{Җ��=���/=�o��p��C ۝����Գ2�ſ@~������S�Y�C��F.�]x�IU��5U0uކ�a[�v�{�������;�5�������u�c�r^� vԳq�KvHY��Nz�����Ѱ=UB��>�|<���[�~ӟG��9�u�7�U#m���Ƣ�h�ѓ�t�ug_w��[�kђ NH�#�`G�e�M�_�qW�is;��{�t��Ӄ9�ʉ�vz�;t�*>�^��W���uB|\ �$��@�y�P��\:��`� ��������#�/ץ��O�~������h[��f��RCV$��^SBY��|��@�ϑ���
��j�fO��G��<2=>V|s�;�_��@~�TS�S^��!��=f����u=V�ʗ{�;w�����}�����dx&��wͺ�>���f�@��ˁK�~�h��'γ:g��jr�fj��Z]�s����NEgj�j=��w��2uro�O�^O�21�z6�c��$��	L�N�Y5�c��ߤ��Ǚl-�U�o�/O����o.%�9����z��{���~�h�"��:+�d�S/����*��tƅ��>�\�v�Y�Ex�Q�%�9Z�j���0�����0�m��i��5�r�zO�eB��1$0�}ǩѧ��8�]�+#,���OL�.Coj�ju�KH8�X�V�'P�ZH�z3'�+y�c�\S-�����Cfn�r�F�䰣N�7>��zN��=�������?�V��E�'?W-dfn^����ӽ�8<���bV}�����~��,~99�3�(ӡ�T�J��.�~���x��c6�y�s�o��R��@>�g�������Q�ۮ,a9�fT	�,_ՓZ{��}�������_s��k��_=V���@ȉu��{�z�o{e�}t�%.��<>���D�Դb�+39{%z2T�>��+TX5��'Kޚ��1�W���и~}t�q~�tƸg5y�+yq'O���k�.��>Gb��&nU0�z���O���{��Ϝ�u=ގ�&����o�ܻ�;��*�a���wP$���<�T�s>��<�P�_�r<���'3�L��;^�ݽU����6�j���gçD�n	ўB���$��=��Z+�_�v"l�y�f�ԝ�8z����):UǷ����a�mO��8 '_����^ST/a�&�|ϲf�w}��#�'��w��z�������K��o�'�Ǯ�qV�jY�D�H3�Q\e��������ҊՔ���h�|@�\�~�%�'Z��U�(~x��db	�^��R+�e��f�������k:Q�&�o����^���8�t���Bq>y�j�Ȟ����p)y��g-�\$�>��Kt�j��:p���=&��.N����{��wZR$��q{��z�����������G�ԉ�}�:<Mǽ��.=Y슸uU�}��X���M�Ub��CĖω ǻ�Q���Q�ƣ��M_��ޔ��5�{!��+;�/�ԛfI��+�ID߬C��T�)M��R��U�R�v�Ɨ�����<�������2p�l�yp(X���[=�7�r�[����!9��s��p:pz�i�qOk¯e�]yp�<�T�_�
����Zk�{�<�✛�=>�z�޺ޑ�h�q�*�L5ckC��86��:Z�Q�]�����������-���<��F�H�K��׌��\P�~��g>���*�aޚl��;Y�e#��ի����)@��x5���"U;�r�w�#�4=�v;ʴ\o�n�����eIt�&W���~�C�4-̯~���Q^%FπZ�.W�x���=ң�����=�Cؿz����W���noOp�T��ր�%���7
C�k�F3�
�T��S	��D�f��}]�ks�傫ѷ�����q�]E�ԒU}2¨<�ϔ�Ӑ��3���TB7���y�?�R�v�������rL��M�ʵC�rx�,��h�7�2�y ��"]�t������rϩ�-ͤ+Vv��]Q�M�k4ɓ��?zgq����RR%����"nʸ>Anm^F���#W0$���{���w��f{oTא�sc�����M����VW�ǖZ���*ԐU|g��ȱq�J�/誟'+v��Du���||:=y�w<ܹ�^�?c3�z��t�_{��݅��ǣ�e��Q%ўAH����{n)�{���݈_���*gG�Cǚ([��ё���V�yQҽ������ǲmO��"u�ʻ;
�m�w�ڹ
J����	�ǧ�.�L>4��qW��1�ב���&����uǮ튑��:^Go{.���L��� SD�3ΠW��>y�|j�w��9�����h8����Ys�g�����	P����X�\:���p�O�6H!����|tn@/Ƣ�w���Ջ��>�b��l���8}�d�<k@���/�X�3|�ꉌ��?.���]����7߻`e�M�s�oe��l���URc���d�@�&j6+�� TB�W���sW{T���}q�gިu5��]�{!{�ע���V<7�N�E�?P�����/\N����q~'�U�c�W�
��+������1~��[����}�Lh���6����3�������\/f����Vb��V�����R����	'%o7DI;ɱ��C[oz*�(0�r�7��R�XN���S�[�Gq��k��2f���7��ho!��������<����;1]F��^�!O�n�-��zb��/�
ܢv#���f�Fk$�N��t��E<o��iIM�"��y�4�[�Ц�;�65 <�;�;!*��H��4f4t�s!.���9y�V6^[��}��|�$,j�&u�U���f[�X�`��_o'3[�H�CՎeCj�`̴�$�?��.��D�֖Gti��̫�ZY��tvØ`)ܛ.֢��s㢛E-Ж܏u��]�4�N��S�z�G���n��\�&�҃GřV�9w��l�u:���Κ�2$��ҳM��3<�sU�yue]��%R�!w�;L:�ͤ�l��A��T��ؕ\�IdQ4���~�zd�F��z����gd���Dؗ×Ixt�e�J�	��ri�*����}4�l���̽��<W�T�K:0�sU�kKz]ZK�`]�͐
�X���Y�w�4`#¬�(V��1�ٵ;wKv6rn�f�V[�Ι�vH��a������⑛���n��Ea��
�>o�q�N����y�uyE 6t���մ��<X2sl!Xຉ��o:����aa��c���j����`�Mi���.skp�M���g k�(���α�\G��A��L����3x@E�0�����i�(�]�W	Һ�Dↄ�j8h�5l�f��v�3��sL�.��[�z�͛w�ٳ �ib�2�ϔx�v+������۬W���w����񥦥 �ݑ����(�ER��֢F>۬����l+��W�፺�R�zݸ�{��N����|�����z0�OC:���1߅"��:�0�z}=�
\b)���>����v�Ĩ"VK�y��e���7�����=���]����e,��E�9���F:���G��m���f�\�a���w��D��:��FiDz�������i�2�$� �O3y\"��xa|����Z�]e�6\��a�æ�٩6����8t�f`����ۉٳ[��tNQ�5R�qQj�âX7LC�*:;MZ�_��"ѽ�L�;����R�E3��b�`��4z�aے�b3B�q�!������d�Aq��60V���$
�Mɚ��][P	jΜ���vm>\�9�؏yr/uf�g�y8�^O>.ߥ�$rd��ҕ�T�mgto)u��(���(mWv�,$#�b��q��W<�'p�����I�m��n����p��������{ٽ,sJ�sQ{r�ih��K�3���(2��6Og����!�v�L9DzS@���|���� ��3t����6��s4���u��R�)��]��%��� 
D��&��bō0��6�
KI��S˹�#$D�$	F�A�A�ł(��"4Qc���*5�s�� �k���s��鷊�D�HF�6�D�@lP�H��l�Dh ,Q���5�Hđ`���(c�a�3[,����S)�b6��D��
HɊ#'.�w1ň#d���c&(M1�F�i4RC1�x�Q	Ex�35�6&�1��WK�r)LX�Dd��hlDE㑙\���I(��%�tWwY4b��E���������x�g�V�@����
�ü����ȕ�Buǝw�.p�%��F�|kgo �Y1�,�W�A0�M�đ�����O��ҖS�����Ȕv������
�xKs����W��x��^3�ǹ�Ӆ��h��+h�C�N��`�t;�ʮ7��Q��ˁK|�=�旈�}��?\,��glی[+�g}�m�,��s�����GN��xc��m~gB�S�e����́�E*=鼮sϸW�y�m���+)��{ޭfo�]#B�H-|�b�gȜ��1}n��u^bŕd5� v"��{��VW�,.�~{U⾲�*�Ǒ���hm�.szϲ��S��p�L�fJ��'��z�g�O�w�${W�l{�y(5;jYqPˉ����ý��D�2���ѕ�$��y�ۊ�N��<���g���j�1:�����;wx�%M��:O�� ^���Hn�G�gh�zn:�늷N�,��ZG������ݷ�m��GNO��[�#<�Ư��>7E��!����
���pm=%��4nN:�������>L�9���=3�O���UW�32��U$5b@�yM��=�^6���X6:y��Z��b�L��dݕ���/B��WA[�^����3Z!M�]\�S���lk�;����������U8c`�VW�v�9�e*�Z=]z��+�n�ܣ��:xs��ξ��(Զ�Qbf �v\���ӻ�j�T)o|mMXy�8QT��EJήQ)7�~�������^?O�������5�~�\S�>���Hj������]GK���]�K'<�Ƚɯ}(:\��M]ȿ�u�}��>��F �P;�^����>���Naݯn�sAd�����T��;W����MB�m�d&���F?P��z�c3C`�]��#Sy�ʯ��\_�z����@�n;�Ј���K��jj���\u�@���4+�Eԙ�9>L�j+}�w������>���+:��exmԽ'M��x�׷�弳���"��XN�\��^ُB��r7�^�?~��~�9�Zs�g����@����J�v���fO�Js�={���O���D>o!�}K�"_�|r#ޚ�������m�gI���"ǍE��I��YI���B��� >��@R�hr���3�^~�>�����B��>�G"��U\�>����f��I�[��X|g�T���d���5��������1�>�<9K�BO�O��}�s;[�m��(^��,��_IhѕQ�����.f�U0�>���|}���Q��gY#��wY�U��aJX
��%O<�ە�ºP��dd�e�P�i׹*���r�G�	mm .�:q�B�?fRYƺ�^�wnn�^>��t�'�.D-��9��ʱ{EέZ�}N�����rב��P��;D�-w>F�p�y�K8^��\C_J��}0֭	h��s)��N���@���,yT;��[����&s�Bk�����	L<�s�=$�w�g���O�g��Ig�=���V�� t�\ �<��`y����S�܏c�s
M{����f����ٙ���:v�����m�_�����a���S�p��� t���4z�⒛�\�f���)�dף�||���W���zw�ö=�\M�}q<o�]��MK6���+�9}蛾k�r���J���QL��0�|���-�;c�҉��&���\���
�Ű���E���k+|�C�#���`��U:��=�����W!P�U�*=�R��^ w�i����:o׸k_�j�^��p*f��<�O��42_V���_�ѿ��5�w���Bn�H�C'�^��;T��{K�&O�ܨ�}�T6��4�^��9��\���V�Ok¯e鹼�yB�!��4
ꌟu�%sg}��Ϸފ���O�������a�;|J��L5ckC���iє<F{�=qf�='�9D�U~D��v��[� �3ϣ5������Y�חL�q�;�c�ئx5C	�"+����� j�te��I��Y�йet�UW�.�`��X*1>�)�[��.�6��,An�#OP��Q4v�&�U;�ł�]3v�H6�gm��*�Y��M�ss�E�@�x�ś�k{�r�J�3�-Ԧ�gc��,�2�k#j�}�'��>�b���e2X���ldJ�zs������)߻ʴo�*�v�̂�;�G6�����q�椿О��7K��_]��G�%X�`
��YzW�R��|�����N�g��2}�ϣ1q��T���;Ez�	Co�a���B��R7\"4�聮���:^>���,��][�u��\u³�����=��.7κ�jI*�XUg����Bs��kŦ)�I��B�V���͂�z9Q���?K�Y^wY֣p�Wf� �3�H>E�*P�^�2%N^���ٞؿwl�2{���FG��1��>=q�;�vAu�1��RͲ�.���V��v��������a#�\����Po!��-������<���W�'M�_�=���Ǫ�\�*m����>�/����lAJ���2���K}�p�C�y���&���|���s{|�wT�yDא��3���8�������a񨅼*��l�zgx��'��e�X/�����Sku��^����3l��:��Ū��� t�~�*K�6~5]�:�/#���J���O36~�9@R���z�+;�o��M��uŃ4�b�ߵ&w��Y�v״�{f{tb�ޝH�s���]�Q퀱d] r(�wio={ ��P�r��j�f�kc�a�r�=us��f	�q������ �]RtJVD�m��Eg��n��c�۞�6�r@���d���>9��>bp���.ez���Hj�uX�s�4.+Ҵ���C�W7��i���ݦ�c�gqI�^Wra��2T?O�w�!�����C�^���yA�1�Q��|�˷���N<���|s�y�?�����=3q�O�=q���ѵ�|J�U9�{�-��6j�Wz9,��.��aʜ�!�{�4T^�[�W��k���U�ONG�49����دS�b{s�ݘ�w��zQ;@��6wj=VW�IxNǾ���2UW��s��8@�Y���q�� PJ��6���׻x=�V�܅00�A|d�t9ɞ;Ex�Ke���W�gc����ߜ`��\�.5��x��:�V��Q˽Y�V�Y�A�N&�����k�:.����m�5�=��!��7y��H��y�ּ`g��2��~������Tg��qȳ��Y�2����ǹה��;����ٽ�g�Et�U��	`�p�����O��z����Q����B�{wa,�ж"{;�����]��>2�����qE��]��G�O�w"=��z����w�wi~Z~ĿM��5������[2\:h]�׈út]%13��;%mՉ/���L����pdk��W<*�H���V޵��H�j"�д4U�7d:�Bx�����m�6����=�?��1J�k;Xy++�^c�eVq�&s��Pu,�Zu�;� {�aD�����WFR7�L��r:�����<���g��#�O���W���M�d��2�}	`��W���x:vKd ����Cґ�2����n���� ��U��F])���z�G���9:W��#=SL���D�ۂu2Cs���6
�O��Rc
�B�;�|�:��E�;~1��޿�ޞ�}�TN���ƅê�f��� t�+�4/��pV���IV���G�����vm��u�ÏO���Lz�`W��늸u5�(�	���K6�o=ؕr���7�[5����dEG.�ȶ�x�dxπ�g��h�PR+���	uUN���̓���#��쨩�V��>�ʼ�zj;���D&���c�Mǽ~��ef�|(QUi{�u��^�~��p)��*��4�{^��qE��/-��y	z���&da��MN/h��'��`��]�Hɚ��x�91ч߫���K�tޕ�5q��킶�L���5ug��Jii���Ew�o��%d~�|=�׍Yߡ�gng�U���Qo��v.�{jrS����1o�3u�.;���΃���!�/�����{��3ݶN=~W�_�����%��靆mS��<�ILS �t�6�t�rd��Q*�U�X->��aZ]��58�=ZZ�$ �'m�i�l�b��N�0l���đ7g/5f��]>�qt�=z�C.�p/��{��M�u�0�ٷB�'2���4���f&oz��^_�߫�W����.L��#�W��D������i�{��ڤ|�mA�X9z׼{eֵ��ԣ�Ox�5r��J��Ґ�Q�����M8�SY^�#�F�x<F=�����*�c��]t\�J5'���ug�d(�|����ý^��O�������<s"�س�������i\��?yڳ�r�%T�S*e��W#�&�������l��r�sc���}�S%�=���+��Ӟ>P:tK6�	ў`)@��s�B ��r��-�>�_�[�lh�����):U�jT?]� {j|\ �3c���o���������u�-���Ե��rա�9�_�l{Ը����x�z�W��2�Ǹ���\Oou��Ը�@o�@B`��/�>�����~tÏL����tx���\��@R���z�|�MW���:��H�/� ^�W���n6a����m_��ޔ��i�}����if��V����N�y�Sbp�Y9K�t�
��� �U��aˠY��1�9c3ʚ�gT<���%��Dt u�\dLS���Sέ�ed����:��|��J��9j��[(�#�=9�س0���/w��S6V粓 �A�S���ṏv[+d:�ˑ�md�z4V{ƴ
�o-�q�=S
d�B�mxU�R�v�Ɨ���P�e�ೲ�zj^{����2n�@w��j6��0��z�z���p:p�le/W�tDoiˉ�z�ڷ���B�ˍ��;���7���������dTq�*��>�Z�����j���j��#c�Gx���u�xϹW�#5����zi��z�G?^]3�G���i��I;*���Z��Fg�N᎜��Q�qmC��c"U;�q��zs�4<�o��mP\�޺]l��"f��M!W~���Iݸ3�P\é��7�Q^'�m |���/J�φ>�-� D�Bs�g=��k?S���/�G���-F_�XO���EG]t�6R>�����u�5P�ᳱ�y��\��Vtw�������\wg������A}d"�e�Bg���򘸧!���6D��]���k�[�^v_�?Tl�_��z_�ȯT{��8�/J�L� ��1�<�o҆W�#Une���X�hz�wޜ�MC�_��W�������;�vAu��ܩGad��V|z0��v�?N�a&��;�q�7m�;��V�^�Y�f��ձN��-���,p�u�W�$Nezvp���]�m{�Q�M�+��Yq���w:��������Bj�⩎�d	Y"�=�=��945gj:��i\����ov�I7zސ�ۋZ��M�t#n��9]|}�@�1�O�o��O>x�E�t�z2<���{���l�8y��q�t8�E�9��ݷk���g�=�@�Pf6�:��W�˘|V��+�5�d9��3j�~5�&��/����g��kO��3�������T�X #��2R� �<�0��-�p߭�7f�pF�Gz=$�J�]y�G������A���q����ƭ�T�-T����@��QR��l㔓:����������6d�Ez#�����'�=3�%�N��Y��+�n!L����_K�񠹨�;�,ϧ����Vv1�>���ʈ����Ŷ�d[��y����@K�^���;�JQG<j7|G���ֻ�{�ǥ�oD�xk�c;]Xc���?����oޟ��qZo�P%�y�Oע���h���c�گ����0׾�J��!���R/j�;�>������g�ǧ���bf�ϱ)��x/��ۑw
|J�p4F�����/	�q�x��RL��!��=q��Qz�/6}ڧ��>�:�%o��?\�j`a���2}:�VUq�+Ċ�l�@��Tf3����|��ct��a"��n���|���3��
�>,8j��y$w��j1�0�R�!Z��.�}v.��ףl�4K��Ց�LJ���aw_+�:������d�֎d��:����DV4��ſ�eҮH# 6�.�'rF+}�SL0}��^�G+�^��NmO��͙����*}GE��D�J�e{G��6�{7�S���*��I;^02]&VQ��[~��ѧ��	η^q���6��=}+*�,��ig��(�3�q�|6hyF��9k��O�/�:�!�֣���T:��W^�Y�]v$�Ky"Nz�q���bI�;|�}ty�������uG�����#);[��"��Y���z�&�a�nԲ�$�1�&��]B�T�/���i�i�9>s�����]ɷO�.�b�g�e�D>ꍸoo�������9���L�H�!x�{�yFzs�lڻ�RH�/G��\w��:W��#:#�V���������7P w�/ZhS�u�l�~����n�f��x�{=^��g�z�3�������q=���fYH��	�����p/s77U{s|��_)�謔��1��f�
�w�Ǐ���q�Tl
~�\Ué�
��ե{���TfŚ�a��I�~g�<;�5y���4��tEBJ�/!�`u���}�}G�����kZ����Z��Z��V���[kZ���kZ���m�k[o����m�����m���ֵ����ֵ����ֵ����ֵ���kZ��嵭km�ֵ���mkZ���ֵ���kZ����ֵ���[Zֶ��mkZ��mkZ�~�Zֶ������)��֠K7�,�0(���1$���%T]+m�U�Z����(kI$f�ڛU�-�M��4[&��l+h��-�ͫ먎���5�X�����Zѕ��j��kX�[[$Z�#k%��ѫ]ڇѮ�UEKVd�V�ۧwU�#�)u�Y�ܱ�l^��ʮ�ww[6�إ��J{���Ȫ������kѯ[����1T
�[�n�	&�77z}���ڶ�-���6jhʶ���vs�2��u�i�rC���v�v� n�;fM�ܓwu�I9ҡ�յ�jZ�I���i�v8Z*��Vڔ]�q��V׷u��U��A^  ����;O�y��{�m��Wu/w���W\L��[w{z�U^E����*��1���m�ztA�����{P�w^؅V�Z�r�kM����  �_�b���v@ֶ��W
	t��<q�EQEQ��tQEQ@Q��QEQ�C���@P�Ow�(��(��;�iǢ�(�����Ͼ(��(�h�^��s�ܻ�6�m�wwM)�jt���   wQ�ee�:R��/^0�.��հ�����z�����W���z�k�Y^�ް7���n����*�M)d��;r.4�i���kR�mZ�M�   ��e�҉N��u4:5[�{ާ�SZ�{�v�i�U{���-����zݭ��cӗ�h�R�y��:X:Z;��k Ocp�UR��ճ���ܛ4SZ�Dl�[��U�   ����[�������Z�#iѦ�ۮ��ov�r�niܶk��1˹ۭ��*��K���R�����U�V��hs���a%��pGn�LJw�����meu�nV�۱B�   >���[�n�����t����v����
W8����;��z��^ͻ&�;�i�um�l��j�J��۷�z����\��wi���lp�)wmn�:��oj+[n���-ۺV���]��   ws�]�[u�.�R�u�ڮ�n�v��������Ҵ��{x4�����v���������w��Ks)�»�����M��j�v�;�޼:��Zt����MJ�M���[Z�ū����� �}R���|z�M�J����Ht�gCg���(Pt����r�]���ӵzw{Qmە��-�s�M:۬�w����ֹ5�Ǜ��gC]�+p9�]۝�E��T�b�6�ڽ���u۴u�  Ϯڝ�J����m{��5�����Cn���VnT�����\{���Y�c��ݺvz�T�����y�:t�S9�h�;�wG�魣
�Խ��.훇%V�uݹ����v�  �}�����	��{%�ӻ�:��n�ӧ]N�������\�=z���6Moz�҂��of��;f�VݦgZR�u=�=Q�m8qJ�� ��T��� "�0IJR   j��y4��mL� )� �*   ��&�U   I���b�&A�<S��~�����~��k����z��zOQ�:�}���}��|s>ߧ��`IN�	!Id! ����IO�$ I?�	!H�B!!�^Y�?����d����ny�O�3��	�Z�ªL���)$��*^�ܳ���v���)3F��o2;�j
��^۬͸�^N�:��0�m2���#�k0LG0��Sd�dO�grUZ��)f�;M�'m�gi@����#���+5S@�Ƅhm1ص�<��Bҽ��k@p܆h��q�)��wDk�8���p�Y��ĝȓK2fMb�����:+u]^@VCCa��Hm$�«5�xěop��R�F�8N�@Љ��-�-q�߶8�e������]�̒\dl*���[�h������P�HV�4iۀ�<K�R� ���o��K��}>c�>���U��!���Y�MKt2EQC5i�Mi/�G�Ņ���M�^�aˑ���ǻw�7зf,�̷X�R�M3p��qS�S4�f�꣕�Y�;��D�*y�aN��nLz�,F��|V����dg1�(ڃ�H˧E�cC�Ow������)�NhY�����v���e����[��y}ϵ�r) 6��ds=d^'uW�՞���mz�2D���Fʎ8��;�w�iw��ܺ��c�|?�е1ۜ3T�p��T�n'��	�#��\����#��MCBZ�ީLa�!��n�87g�L)��6�w�e��2�0]�z�opz��]��J�N��l! mֺf؛�'�oji�dƦ(�Z��\e1mf��j�whL�Pr����c�I��`���CL>4���&�X{E�Q+Q��9�N�А���Hz�G�xų�8\h�5L�F8��f^Rդ��Z���ބ	�K�t�*�Bt|��a�a���l�[M��cCH�g��)�X5���G�+dҮ
�I�:5��Xz�K���P����RD�EV�cM&�F��\�<�G�,�aHo� J�Ʀ�9e�P;P=_f�8�!�c.�$�n]�Q�fʺ���1���#365�`2�:��2��:,���Q����v-�a���zqVȂSV�GE>��uzi*{'����%�r	z���>���t�ȉ��7�a�V��ٹlm�P�H���y�ƭ��G���A�(��{le6�.�FF��{�/��j,"�E���)6�r��iLA��kS���oU^�3�|j�/j���rx2�l�DQ�VP�������j�v�<g.5���nͬ.��6�cV4����iVT˺)&����xV�^:v�jiq���HT����X�yh���p��W�,d��Y�8&��b�j�;���&�ɹ�rD�����
Af<o]j��( ��!"%�QՀʤ�k2]�v��I-$�n�utZAhb�'u���;3~x+
�\{��j��Ѷ�RìFR� X%�{I��>P��u���cC����]�,OR�bkD�zƖH.Q��~N�-DEn8�,��{t��X�Н�[M���Eǥʺ�,�>�3^�VӘ) �z2�Ym�2�4\/M�d�aj*����4�IN�=�2Uj�7z�F¨� ����u]#l��b���v�#ш)yv�A���ň*��+n��E��U�ڋ*��AjJf��V�[|>S7��.�ܫ$Q��AȲ�4r�ƞ<"�(T�̢��&�qȩa���V�ȋ�^`����"� ���p�ڵ
��LZ��IO� ��w��=���T�+��܈�:F�Pt�B���ųLB�$0�:��6�����ǡ���(/a;�~�h�
~j���
[%��گ�4���nB_�<�(y�LbH���O)��cXF��P�6D�N]H"���vbxb[6��(�wj��wa��K�^�1�IѠʼ�ި�ʂ�k�{CE�ۧ�k�b;�&��MYw}�S����6e��v���[� "5�����q�<޲7|=����[n�B,����\#j�eAz�k�ya��2��§2Cx(�яr�[�œa-�!�U푴(!-�U\t��@�2,��Hs$v�*�FIS`��ܘ�qӁ�n�5�[8�6
�ڔ!;���rR@b�[7��-m5����&�HwP��7ch��׸*(���I�~413z��LQ�чsF�b��K,���#�u�,�6�l5�fj��ku��bh�e_�%/6�l]��ؚ�6�4��N�`0�z�iV1%��^#��x⫕�6�j:��7ҳC��]Rg�԰���ҟ����n�-��6L
g�F��!��PcW$u�4�z��tz��}�!B/2І�֦��m�
��[.&�݉e5S-إD@i�I��4,�2��h,ۭ�L3��ta�i���с D�hpK����[u�_��h��P��m�,[��Z�ýt�YbS��U�n�Y�`-�ldrv������M}s��5���-+��W
��z2�>IU�Q`�2;��ԋ>t<�L[�A�^�5X�OR�@�sPf�$è�F��0��r�<z��ٶ��]+d�@!$��q�:��᱔�\�0}�Ս��Y�SJ�o6�.%6��
�{�M��S��7	Y�	�i�w6	�}�s�X�Uy��Z����!� )Qf�)�Z���{n	Y��w�v�ZX�� �*Ay��[��.ai�P����Wu	�Cr�fY��j��ۧ�%mM���������w�1e1m
��+����7M���ze���,�ٜ�i:ӌ=e�]��;�N�Ś�1�p�Ӌi**RfVz�n�VhͥMCykƲdTU��J:v_I<�)t |�T{K�~7����L���S8ֽ;0H6�h*���YS6��ͤ�C��Ǎ"ӻ�3m<��if�o�2I�[;p[����L�qF&1w<�:#��uj33n0ګ��R�A���t���+I�)�wtYm̉b�[zN�L�z�����]�!7ِ��,$P���f�Se�ZN�P+�Ѓ�9tf�-Jΐzy�CV/�۬��ΠN��?��
�-�Uh6 |��a�,���,7j�k��,�(+�f�,��vZ����BʔH�F�V��^��&:of�� 5m쳅�u�KLnb��1�u�yl��[��C�h3x�a�`Xр�4�妥�Ƙi_�U���,u.��wx���;�yt��F��=�q+y�{6	� ��^��[�7k,.0pXm,z��8�h��.`��$��ب���41m�	YpM���d�Ǔ1Ь�,�/$47W�z0�yL�Lr�M�-��7u?@��h��>��|�t�M�:ڴ.��,�ӏ��[�䛭\�n�$���%��r�[ub���&c�ܲo3i�oT�3l�ܐ���O̶�c�l|�\���YJk&��SiQ�1u%��+ȥ�n��]��I���KلV��������]�7{Bc�8�D�Mk0)v��д9�f�|3E�>��ܾ��������C&5�Y��7N�*�	3��\���0�D�&�ʰ���wP��)�S�(������j[��	�<�v��h��9�Zo�|���J�Zcv6��Ӱ��nV�t�]!y��^�#͢�_�4iOB׮����`��S��XY2�iҭ��ݫ<A�觰�a��/!�4ڼ�n�bi+��:,Py4��N��V�yD[���Z&:6�TVUŃ�&�d O�ҕ�=l��YLl�l�-���`*{L+$������e�̳*ݩt�V�iD[�����ê$?�&%,�t�V��������+r*6�+l�t�A�dFr,W�f�,�q�5��x���|����^5���W.���
���Qm��-��E#��2=������-x��v��j�^!�]h�36+�Y4��c�z�>���wi�4=B6��р1�t*EZa$A�73i+�'m��E��!��v#�"�-B�8CA�`�hf�g$�%d��%g�����ҫ|.���F8@×��<���+������L�7�|N�VY}B�Iww�-na�s1`^�iڿ��Y����.�XA^h��1�fzmu�95���~��lYZ��ɺ�+��i�-m	�cV�Ab�����^��հ���d��efĝ���Ѷ��X�n����[ͻy��Ӗ�5P�l|�8Vʌ`ۤ��.F �]�Q
ּ�M�^�L����cQ��<J�%v�ν�l��%#���Af��6a�'��j�mEė���V�qo�OjF�hA��*Ʋ��#L�H*$��d2Wl�ו!�u�p�U�x�A옾�ێƑGk~�)���G�����3i,/Zݕ�� �f�nMT$ҬY�9	�g��r4A��Z��V��l�.�4[#r��a����6��+ �f�ָ�(�V��GOu����#6+�7&gp��ʎ����Z��+Q�X6�'�MxՋ�⍧VRe�
��Y�٦/n�=�;J�x�Dܺ'-�CH&P�[�J^������q�3�"G�D�3W�� �m�Gm�F���vF�cx"�e`i��˽�(���X�6k2��r�Rf[��f������P5aJ��e
Up�Ԯ�L�����Sld�ՅF��ɉ�E�|�}wX!����Qb�W�f�-.�(�Ùp}��5�f=`�Wݹ�����p7��.�$;<�l�.��D�jɓT37w#�� :�n�h:V�ҋ���NX�6љ���m��-e��,JSw��*B�S5r'MS�1�;�Y�v�]����fP���NV[5��3�x�x�m��������5Md�+!�6c��.���-ۡ"4�)�4�eZܴ����3&�cUݻm%cy�WQ��u�A�ч���|��n�H!�%��3YR�������,l<h�&chn)����7�Z���b�Ѕ{Q#[2�DF��l��7y#����(�|��-�Ԓ�\�x��H/���8�p*�r��Ammp�W}Lc5��"E��'���<�MwY<sA�MSa3�F�b���^&��KN�I|Y��O���)������T&1�Z��t�ضG��O��z�Uh�ɫ>���,4l�9���N��J��&<�c���}X*�H=�+�ni<��C��^a�$MlIRt��l���lS��Dc������ߑ�[_hul��j�Mt��[��ZN9�L�M�A����D���7b�,�c��e��F5/Ef�Xb�4!n�J,��@�x�Z��v��QA1�>�*�ѩm���7Jl\ì�!J�4*H 3B�i���~�_7���Bۈ�B}�pTQKT�f]''�Xb��Q���^9�Qw@D�է����� "��H'E��{��B��Y{mn6�W�fݒ��c*�A�t(Z �I�gA�3`�ě�t�����`K)f�~�u)�����`"#�Q�j��G5ׯG�W��Rx���ˑ�bj�,Q�<	�A��Ɵ����әK2͟�cHaK�x���6��K���[�IQ}����X�\����p<�H��h@�F/�5oi"+R:���ͱ7��E&��:�
��չ���t�nͫe��Z�0������1��n�iД(T�,�*�]VSOrZ���rA���A�Щ��OK��wP�;!�<��>��%��EZ�
ܛJ�*�qfU�ᬢ7Iѧm2l�,�
�m3���i�A'�*Ε�!��"��35�e1��ޭp0��p�76�,�q���8��s�h)�B��x���.�2�SPg�Tn��a���ɱ<W�|N�h���R�n�+�xE��Um�YedVL{vd%��@�]:6����\5��`JY%���ݶ(cǊ����ue\��&n�����$��!Se�"����m��H8��g!F� ���n��y��m�Ð`�MSJy)#[fniٕ@�t��"���� 4"IV�CqSC+#0z��'Z�c�н���+q�q���0�b�-���FU�y&g���R�����ń�^I�D��mY�z��5�u7. ������دX!(tc�Z&`�XТֆ%^�*9�ҫY�k�^�Z����H���.�4*M;i@hPYK`g��얞�A�mh���'�uh�ouAɺ��`h8��X�F��[a� �gҎ�AhM�*!q�C��D{Aț��d�H֢�3+hM�ZXAjg4擮3$�7Y]�!O.�h2�Q	���.��џX�� I�S-匆P��z����E����@����V��X��̥!oXģ�wt�µ`yZ�)))N�q��`uv�6�P.Rێ�M֮`Q�z6�v�Ӕ�;�Gaeoګ'�=´U�1h@� �o4�͓X�o����Ǫ�����@S�2�����p�mԠ[V�9�R����S^/��k����Z-�K
8�q�6M)M�kX�#�"����]��5X������+(��x=��Bcڱ��rk9Vժ�NΌYxq@p���^2L�#�2��Z[�/2�ѡB�mYN�����!
���Q��1c9��_=���9w�e'�«�&;85e��eQt�ɤ���~�Vf0���l�j��@���F�.-xE]`sA'E�O2���a�"U�G/M�[��A���h @-��`1�Qs!�B�F����(�^'�������Օ�h]�.�C���5s2Ί��qVݳ���["n�͔��@�'y 2ېZŏꖅ��P��$��Cg(P���.ʱx�l��X��nPP��Ys6�x�kBݬ�v��%��6
�-��e߲�6 $ؙ�М#�DY3 ���#m��ò"��ufj=��@D��vڭ"s��ں�d���J�+4��r�bQ��l�5���Ǔ�]�u��;>>�^�]V�wmpS�+�]��Ύ](u�Z�+xQ��ōZ� �9+3�w�U�6Kl7��9���j���u3v2�\�0;c��|C��705`��Y�~:t.dx�����כ� �֡	�5���ާ�3];˄�㖏	��u>�WD�VސO�VȌ��q����ᓯ[���oi�}�j�_Y�/$Y�˗z����,��o��7}����ȵP�1�U1
2p�����5]��vlZo �ط<��ޫ��"���,����B�j�y^i��X�cBo&�7H����aǋ-�L�A��Y�ݨ i�T�ݦಯ%����\��kʐ�z����JĬ�I�c�M�b5k̣�x�D�3b�E�ƹ��0�@rU(�	Zy7͢{>I�F�!\oa��bFe"���T�G��E��;�0*�l,ȳ��B�TӂSt�,�lx�p�u�/����xU[UT(����L�c>
h#�z������+�=�|C�/?K�Qj���N��뱇) r�5�17Sz[k�w}���d8���Z��~�!�/(�^��g�q`w&�lZ&��^TΚgep����1��=�h�C�:Ʊ�bD�D��WKKJ�9�C2��9ZߤyP�f���w�54޽��{�ءYr�}Ԫ<�A��[˚����y�0�\J`,ZS���J^ͧg���:ؕ>S��j��H�S�ː{l�]�.;m	͘\L�cKB�Iτ�.��(�9�V�vY�Mv8�5_Lsg{���$I���8��E��9�]�v�-�,���W�Y��vr��٭������]���o�\������dr"Q���N�-��Gc���w؅b��왱�C��4��AfX۩i�awOu�#XW8piL�36
2��!�
��&��PN�r2�Q�:���&��y饢N�>��َd��d	��.��񮲀�v-���o{%�A}�����8_�*�nQ�2]�ș��^wr�$�Y4f&�A�f�^�x���U�z����g��w�cJ���R�n�7�ڐ9\�\Bi^�d�u?w��}�"���V��1!��m�-.��يď��?��whq���.�CCk�d��������sx��ws��{��d�s�	��0����8`�
�Qj+@����!8����:���v�	�e��f9���O
	� �kL�VDz{r�s��R��i�L�3����:��1ҹ���r��<V�ɴ]�����������<2��s��E�]�"۷MZ���hm��fwW�-���	��i�|@ު\zJh�*�C Ū�x:�mͅ�u�i[y:��Ӯ����D��-u�~L�{L��z�Б
�^"���Ü�s]O�q�>@��}�>�Yً%���O%���;��"�_a��{ˈ��o����V�(���v[N��r�x�]]tf;����3�����l�wg`���ԊG�!��5n��e�⨹�_}yd^���*�E��=�\aڻ"�E
�]EV�*�/xp-�����N3��9Op��iWk*N\�z�7$b���-Z�}2+�t������(5ݙivnG�nC{�S���A�J���c
'�Dw|�q�1c�/Q���`�y��f{��Ȗ���E�E�s�-QzUXu�s���2ե����Bv��t�8%rz��x�C��++��ѕ���xn��X]��_ϕ�γ��6^́�k�l��W�by
52TLD:��W�z�=c��a=�pZ��54tW2�y�p�\��"��VvohjH����um���s�c�o"GU�Z��C�v�qR9>φ���@fWE��D�֮N�M�y��n�N�2�c}6Tm:dC�e<�(�=y�XZ
�s
=OOMկ	�.#n�N:��E<V,o	�0��cMf�y��A�n��,q��:�`�o��6�6�9���!�tq�2���d�e���C�ܵ�c|1^r[c�z-��e����6���C1������pqǒ�SiK|rI7N��I�z���������+y%K�A��Ɗ��Au:<�/d��`m���Q�36�}�Z��8�H�]O���MNn�a`EQ��ۭa�m�|�Zk]t���9�Ӟ��l�B�5~��2�t�x���[�\y:T��0�����]��b�gN�W�����5�[�V�we6V'�tY�]<3�cS����2��$�p�L��J��N�c�D�==�qz�5t��v��:�M@Vک�a������q��Cz^kY���IF1[u�I?@VZ�{�%�ʑ�Ak�bc:}���{��`b�ڷ�A(��Ld罣�v��*���s�X�;P��<���y�띀r�;�gp�^�[��
zi��6��^+�gΫʕ��-�O���^����Q��T���%�7��#���%��&��7����v�²��\�~��{c��i�]nx	�ݍ�������ƥ�O�z�:n_�~E	T�kL��S�0x\U7�+��N�p�gP����w9���^fk�+�qd�?\���Fs�aj.���
t��L`oiC*q^�v����<��yB
K5sr��ޖ�-�&����3�|���J�}gA1쾸�o1f�H��|r�:�n�Ē��O��:E|v����A;۾�Dd��:	Q�z���N�"����EM���Yԙ���䖼�T&��((�����N�4�ܾ�/Vܮ�ԭWi�%�\�]������4e�<�3ה��V�����vю�%S��QsL�vv��;�V�'b�iAv��K�����0d���D�q��9��h���X�AaS����\� �າwG��7�4�J�`�j�so�h+�5t�ҽ��]�2���IS��R�b�m'i[�p�ѧef�kE�;q6j���H���tn	�Y�cb�co[L:E6�/�����F�T��ၶ���~���1��CqS�3���M��]eb�A���.�*���<��tI�0��)����#��F�v�=���³_H��?�V'�L���gS�'v��e�wc{Ӗj�{�%\�s��ś�NOiWQJ�;$��zN���7y�y�� |���:;�rl�
8uؖT�x�έ���k.�[����g�x�����λ+I�ι����hXFZ��{U�:��$�]n���ۨ�|F�}�"%ӓ�ք�� �>�9��^$�bJ���w��T�э�y�ՉE;��kt�6FT�Cj��~e��%��G�k�%M����<Ȩ����r��N��a�ZX\;�3ފ��@�>����8�bx�I�ʚ�CV�=6�n*{5y�Г5�����F�鹝�@,��p�K)��]�}�S��0���=�:�Zޣ��S����e#nK��cQB��j���o/�7���u���>x7��Ex�r5���Ю]1���Gևu�2�Lr�Ra�
r�w0��;Пhn�2�,���,�ChK0����嘪�������rF���:u2H{�AX�f�t-�:��3q6)�β듼�ӜW��l|�GS����Jt��m��}��	�Mn��Q�&�뙩d>8 5ʇ0��j^9&�la�¢{����f�V��Ù��/�H�:٨�(n�/W�Sl��Cr�MuR���g�]�����sZK�	L�T
+����J��M��fHV������Ro����\I�WV�&p�;�!Xَ�j����ۘR�F�����)�w��sşX�{�NQ��E8���XSx��/���LX]�!p�z�X�g�-�������P2^1ՙlVd�,Q+�;mVnN9κX��d�[	ݫ��/f�#v�w۝�};�fAQ����3���;�w�����:�i��Ȼ�̗�:TG3�jS0>Wˤ�Ӷ!}�3T�X�6�Н*+���쎵M�	JoP�y�ٲ薣ݘHIc2��Q=R��$��V)���QvU�����K��!Ylł�����r���Q}������*̎��N�e������tT��{��ݙ�_37�	�ȟ+��s��{�'��:���1��{�Hi�Ԋ��D�*�[�1J	����;y����6髻+����v�`{����}���9B�F�#��l��g�
�� �N+sa�N�N�7��D�߻��:Q�jG��h�Vږ�Q�}�Pt�/*Q"f�84�/��88����G����ZЙ|����"z�v�D��X9Ub�7��l�"񖅒�M���Ӕ�]��,*naC6���ˡ��bڻX֩�R�ņ��Nkh�56�������ݹ���u�V�� t�g�4��E[ݖd�\0�Z�����m�neL��z=�݄��ֳ�ڎXܕ-� �|��Z&i��2K˰q���Ə	v�.j�
��nQ!;V��;� ���;*RsiK��p�so:��вOY���l���;MP����&f�}`M��^ê0�]�����oE�\�Ҏ���*�C��a�������,T�)isٽ����J��!��q��s�MW����Q�[n��[�t�ЮB��^��I>��C�{���f6jv�ݱ�����*ۅ�s޾u��� h<���uu� �'�E�/�2�.�sG�^u�!���ϰޢ�m�I������Ά<�u�1��:�=��-�o�R\�=�|Ύ�wS�opQ��wH��۝��b�X��`���!�.�x��N7�I��b��e�]6�v�.V��k�ʢT"�ry�q�i��N��;�.<��v�7�ی*!tR�d�vT��ꥭ�CP��؋�Vfܘd޻�Lem��o,r�l��ue<QЋs�G��)�x��>p�X��t/�
�y���;��h4����om���n��ỡ)PA�>+n��IN��Eg��،V���c^i�6�d��u�MJ� j��3O����v�:�.�ܣ{oU9p���[��b��A뒜֎j:4z���,$�vU� O��Ie��x�w^^��w��%�"m���^u��fs�'����h;����*҉���&�q��-���8�K��r�>�G��'_i^�5�!V+���`�Y>�H��*AB��D;��Ak'�	����C�����.yJ3��������B�,��s��֨��7�F�me�zʉ
ŁjG���k�Ό��l�Z�F��vuƎ!t%j��%��R��.�5�R:�^Qݚ�`0K�����V:�g�q�K�6���JfV���y�#�㼩1o˭�/�t�H]]�0���NLњ�Η�s�Cy���@Q������K�闘�	���0��*4e��5���7g��X5e�z��b%\��X�+C^j;�u�j^��Zskg�g�Q'�2���r��|]���)v���e�#]�Rwx"ŕ�'Qp;j�qH�u�my���I]xbu��g��ʏs���K��t.�yu})�w�����Ve�켧n7��?MKԗ�g�u�X9��:�m��]��ۉ^W*<��0-�����2�%[�K�����t��{��.�lي��`���!܆�����1���������:���m챯8=T	��B���cB�x�,�x���`1��;x����C2�!�f��W�6:b�]��8d�dw�Ba���"�2!Ұ����r��٩�@d����k�fp�U�)�z^+��&G��k��� Ʀ�t,$���v!<��&p��ԙM�l ��2�q�}(S���x:��2�8�I)Ǫ��h�$���bʐ��ʍ���jY�-#�K�
mV��z�h�H	�� ɚj�*� WV�
���yր�tG��u5�6�ӂ���`�L����u��Wk���WE=J�jٍ7�sfvib�N�.nX��u�k<_M)�3����W�M+��c���qv.�7G�m��*���;4`�Z@��� ��.�Z6/���r4��R��yt-+��ӭE���6��Pmb�Hm*[@���y]�;<k- Rh��G�7�qk���Rǵ�����9k&�=)|�ٜ����b=�9*�o#���&�6*m�[S�k)r
���4�, �)޶U��l���ɮf?n��ؼ�AM2�=�s��Rb�١���[��u���x�6V3��j���ܕ��i,��������>q0�mtZ���S˜D��X��iA���"�]8Ѕ�5:�+��E�l(f݂�͑x�H�J�f�XÚ�q��]�;�>�=YH�]���	"[����yù|i�rt\�`�dbX��wi�z��sX{�k31(h�ST�u�y�Ê��!�ikX��F�h��̴2��]���XJn�GNc�k6��ފ��}��|AȀNo`�5�m�rSb���҉ѾӸ0��a��)I�W�M�#�Vk�I�e<Zz"U+W9Y�&��F�9|¤C�ڽ Ku�����_�y�"�G49���<]��%��=���!��bx%��z��Y�)�JE}��*8z�����u�Y��Ko�������h�+s}7d�#�v�(��*&�#��u����8��� �sLS�E�Y���f^�2���N��Qgv��;.�7:�TF��{�ߜ
�ƙƽ�t홳��̛�zv;�7)1���Tp�*Ǿbo(�����p���BZھ���y\m��f�ռ�o��.�e�՛h_'�r�J�iNG|7qc��j���46g
�30s��O&�{�s}Nq�k�OI3f�%��>�bJh:mU���6]<z�������U�����bV[�6e4��b�)��}p�Lc��{�L�MA~�a{rGn�ףdV7۱�7�|��<��|> >�}����$�����mO����_{�|g�����^��X�6�8�?�姑����T��������2B�v�5��oA���67di�
:�q�7le�t����=�e����;�C�pY�OLJ����]�JI�gvדq�Tcx�f�U:�\U���!,� #��n�u�y���]�A.�ګ�gN[���_/)֥ʢ�/Gq�����Lai����nݖ�FVW��B��E�7
9�鸙+ ��Fa��AYڄ�\��QaqN�L���}����]2c5;�s[%��}ˊ��IwPC�S�8�1(!E�p��5��vi+�
ip�7m�맑�8�'�t[���l�{
c&R=�0�8�n�6�M�]�j���s��b�k�Ո2TX%9I󈻧��"���u�%�W`��-���q��ի�O�����:�e�H�a���0�J&^���ޔ7��/V;%�R랰z8���s-c5��oBU���̤1���=��W���{`�WR�yd+__V���.��y�t�8�(Wc<@=�1�_T�t.��_��9)�$����:&MF����f/;��,N���=�:u�q=�0oʿ�'d�Nrk�yt�^��xU|3�Jr,L�E���	��r����U|z�J�TI̻櫏V#�-b��i�^jtR�6�+ 9xtK�݇��E؈���I��W���IJ�Jͧ�ǽm�͢
	��d�h��Σ��s���<�Uy��Dր��ip��܊��>����X��o�c݌čib��d4��t���]���Z�P�l�O1�h�PK�M�.n����k%u�M�zGyzژ�b,5u����ry6�#@UK��6�4�V(z.�֘��fS�ǆڣ�R^ᓘ�(LY��<�mmYnڳ�8���Wd�r/t����Sw���`�8*}�[�2,���������cg_
�r�Wk%���m�ە.�i�֞�#�ws"+95u���=2�f�u��xwS-�i�Ѫ��/b�2�@]%�ȋ롳v�2o�}V3������K3T�^޺�pwF`��+7��1{��vi�g�щ������+��!*= �C)Lb˪�*��!kb,�C-�x��8��`̜҅צ�S1vr[��A�fq,�^޹�^�u&��#μ�kq�򤐭	������ ��0�1cX�9� ��;�専-�-�Ck-j���4E��n̬��wa�=<!A&�wv��%B�t�y�[�q����c�����c��0k��:=��NO��A�qM�{�"M�ݼi̒�Py��kH2�K���n��5�C�7�uj��{1���w�U�:t�Mb�f��gs�������G�fX���^��9Q���,���@��d��!-ՠ��6��^C=��^�AyDn
�QE�Tzv�UTos����E�w�S�=��.K9�������
�Ц���kk%'H蠫پ��2�b(<�����OcK�q�Dj��:�ʎ=<=%o��}�,�T1�I������}Qq뤁��A��R05�wL��n�o�,s�>�6��y��-�Ӏ�9v%1�m�����x��{om�9����'z��u��9+]j��g���{���G�C��ۆ���f�K�2����sԚ[�Z{�n~��J;'�C������A��z���� e+�[�F&em���< ��15/L����.��[㱊P3�}B��[h ���V�/������ ��]�^��P�Y�{q�ݫ�%|�ɽ���&moU�O�=V���Ssq�1�]m��<�5�U��Zt(�H3�:ؘ�#��b2F��U5d���ŤO�Wt�tF~9X��֎bC���̭����'�N�T(@��3��י�j�Z�ܽ#&!���Z���|k��:Ջ
�������[�X���<z_��I�B= �f?�u1�'s�es��i�$�s	�5*�*l���j�>8�[[���+K�g��1��!w��f<.�)A�L�c�V����������U�WC!��$1e�8v,[t�eŚ�0��&5���q��n�3\,H��hF`��G�Ã�LV�/h���|�0�ӥ��k�(���A±���9��Kq�j[���t�l�y���yi��=�F�_�0�����3h������b*Թ�$)���F,��O
�Y*ʈ袛.�>��$݈�|ғo��0s ������A�7,pW�gK�Y��,oY�{�_g��c�H����z7備��C�$Ҡϫ+XnI����0#�gi�v�l;v�������S�`|��*ͣ�Rg!]�D@�
�P�9����T�T���/f)y�O�B��5#<Ζx�н7{7yܽ���+3q���{�R�§w����Ԧ5���vnE�_����n��:�ppdh�;m*Q��[R����MM�޷ Ð��%�B믝�J����-nb5+6#F���h^��)PD��y=�|���+�
��-�����G}r�V���М�q��b�ی��aN��Ճ�c4q���j\^�e�PG�D�Y�����zy턋Z��6������WΉ�M_;ᯨќ�\3u��j�<*k��٩fByT���ӀT�k-�Z�ƒ�M�I`D)�,1RQ�k�U:ˢ�)S��[6����x�˖Gu�v�l�hQ���I��ji�ﹰv�ͼ�����5��೸f����ֱ���{,u�:�;��D`�e���:S�t`���yJ�ҥ�=���	�0\����������Y͐Zj��Whi�hf�,�G!̓;>��P�B�:�2�1N��V\��U��)SX��B7)
G�>� Ր�V"2�<7�:��og=h��&,K�iW���ֵi��v�ɸe��;�Q�����V��u�G����������	������-�ւǙ�ml��E8z�dpd|9�T�]8�w�;Z:'	�}���pko++9a�+�A7Ӯb��2���52�b�Zq:6��C��Ӭ�Q]���7\�r�b�vm ��[�-���Z5�!�+&"�U��/-��L��N�pU�4�����h��ٖkT���~Y���b�/V��d��恣�k=�οuodǆ���n60����������>�=�=�E
��u�:�ΰyVN;�������&2�)b)��c�s^MJ�����yo4�o�.��T�����(t��8wL�b��y�os.�g	wWD��I�P�6�k���.�*�W8Vgb����#��
�ؑ)�ٷ��<���c�j�]R��|��MCCg�(ԬR����ʠu�ΰ.��j�1�EK�����Y��u�K����򪧄��O�L�b���`J�v;{X��}ڜ�F�-�ޚ;���4�	�tq�v��Ҕ��5�����W�NƸ�������BN]׍��,�ȇ;��v���<�,�{�ޥ�Mg�/��g�|���ʃ��0T�V6�!�l����-l�����TN��V�����zv�X7Jv ��\LL�L�5.MG����l7Rľ��[�o��"vk�]̰ ��n�ٵ��.��K�Zj��zuD�$�Du�1o.��%7sU��2
��w�\�2z�1����>xugB�Ec2���
�*X��}��g^>�1CX�9Z��Z�5�y�J��\����x��$�7{��#�j����4m��ǂ�j�R��dKj%V���H��^^mC�'N�����4Gt�V۽I5���MH�.�!E���ښ���br���hQ����ܐek��[�t�X-m=������=�v�mس�(jT��:w46��%ԡ��p;wC&��x���9eiV`�H
n����}�]x�$�)�`�zo[���GK%c�Y��x�����L� �a3�TtT7gt\��V��e�b����/2A>h�VZ���3"���r�(�{����Oi<��I��oi)��|��˽8�F���v`ΥE�&��Xm��&F�hK�HɼLD��޽��ذt٘3(�V�������j���s���笜�*�b�Y+��']�ޛ��5sT,�EH.�o�G���3��f���?�y�!��sBkqg������2���e�zD�EѢ{`(����ɼ��r�/���/G�t:E^��9D,Q��9�g�u��I#v��*#���T�);K`�b�?!��ŧ����lV�v��i���C��p��	L�#e��ucN�1�2�K1R��kY�0ڼ6K@��ͱ���t���M6��Je�}HՋ�u �#��cv��3*,�5r� ���]�me,��Ei�α�s�=�:����zct��9v�t�z�����I���<N{�"�5��V��z�x+�ط.������f�M��ԫG�(l��g(c���EY>�3L�F�֪:����fv�5��­s��v���4upK9`�e��'W)�����BȠ�2����]=�!�T$�fj���lպ�@#��}dt��9[c�tu����9Zw��Y����xe��`��Iݽ��
�ÆfE��#��륰�P�n��w#�Q�m�̛
"�$���eer�kۄ8�EvL��f�a;�"�\���K�u�*�o�a\w��u�|�,7��:��,���ټo}�٬}2��.�ǉ͵/,s��&nǫ�A/J�=�+�3�>�v�UM��i-l�˓;D�� &uuLK>��O4h8��s3.�:���p�JUәjr�CR;N̓s^�9S%ײl�=�Wmfw�4��<÷�Wae%m�6�-��,�|��f�*ʬU�@֥�C���	
nj�蒗{N�u:t}�Y���8��il�w!�}n�@��M�W�������m�,�`��k5�3v3�!	�o�-O�P�i�{�M�ϛ���xia�O8gu��+���;�ك9��w�\�ǭ8Z��*�\MP����V#��
�D&M]n�1e2h��%ƚ`%��FxhW��H_)��m�S�[=&�Aa�&��l�������vQ���}k��*hq�id�"i��:����~6��"添��=1H�Tgop5��(A)����gf9
���3�t$�p0۳��R���"j�����%�� ��տlŰ��|M��M�S�*�hhc�Y8��w\��^Һ����R��3�<!?��{ǭ棝؝�ʁqH5a���;���5��j��<����2p[z��u�;�{�#�[F��	#ykK ��wf�PP�e悲z�=�;ú����Y	\��X��m}�!0�]�S��tr�^h9J�q�_k;ǭ\6����\�
��Rc��k�i�K��l'��-n�a�Y��9�[�x����>�����Wd6]5m���¤`�;6����ll����r�7�u�[08,ym���fm��:��TWdY��l�VqQ=,��&>��x�<���93i���ŕ�5�J]��Ͼ��;��"&;�L����I(<W%<�E`�P ]��D�Һ�a�X�����wp�Ju��\:(��8΋����f^Wr+ �����4���Z̻9�$wf�w��̜x��ˁ;�<P��MwX�Fַ��es����P�烢��4������֬�%g��Km�>��I��M¬�$�6�Ȯ��p�y�|M.�X�d	�vŇ�*Vn��*�\�s;l`�5�=����]�B/�r61���_G�m��A2��褲�WsL�3����gO}��"���Ev�yu�ܒ���Ȉ�B�@NX��+�ֲ��a�v܇�|Λm�B��m�[.<�y2��[��\	��m�J�@+�WIWy8�_�έ҇Q����m�(�y�ی��aua��\�{�c��b{&
2)�+�6l������e��Sd54�@���3��R��|P=2�rɪA��^T:��fbn�wTb�<�=�v�PV﷞�ଦ��a���]$o� ����]M%�#��!�8�aZmӭ��5����OkM��Yki��xނ�C�l�M�����M���ƗηNu�u��TX��eg_�	I�,��屌����MÓ���WU��H�G���=�1Ս�teJ�m��,v��*���m���Pq>9fH��͵�Y95]�*M�u�F#݊U�c��ɵb�˄Y�]�����b�Xt�Q.@ʓ�{������ϥ˕�f4�ܫ���q�#1���{�O��n�]Z̆��U�5D+��ߋ���bV��I���6�HR�mnp���m<U5[��Ric!��%*�=���T.kg-8��i�X�~���睜��yA�sVei��l�.غxʛJB����e��:�x�V���w5c�Y�$��72*�玖��C,iX�\q+yd��a�tNR�=���r������/#ce�r�
��Rl�F�u(_.�[:�ZD�9V�]tVB�;��qV�m��b*���Э�f7�v��Gv�N����mPv%�ȴTԀ9�-�sV�hμ��f,.�fYtk,q�ioj�b�,Af2-3��u�
��u���,>�R�D��r�h>�{�dΰ�f�����hN���U�;�h�
�; L.��X��N�c8_fK����id�reL�ڮ��&+;�=�{فJ ����}���0{�Feo
�֓-)��U��10�S�=y���*M�nA����8.�y{%�q�@֛�x!��Ѿ/��W�r��
"�r:|���t�N�[���o[������{���+��ٳ��ID�ޘ����g�V���R}���9����ý;���6c5���7}|n@������K��5�vh5q@�E���)�<yJ�t��K%6�c��F�U�ʼ�^�b>�-�L]?����9��͵Mx�ő�b�(�f���#vjq%��P�����U�r��n��-�dLqa�i�w�����h�{����9���x^�c�v�G��e�ȋ��j���iIX���@���Iļ���cw(�Z�[[�fL23)s�M��ݍ��g��`�A,���VB1��٤z�6V��PB`�s��ܨps;	���:�����QRK�;}�d�6��uMؠ�O�{q����zH�B�����a�<jn��Z-nr���%�:��8rϮ�m�ЏD��Οg�f�++:����A��AfR���c4���U��Żeb{Lt�GC��Ƹ�L��z^-�p�LWC��m�oxu�D��m�y �2�nwg$ɭJ}�7�Y��7�gEy��n��oM��ˈ��.=�#���'�}��u���*�'��-�]�ͪT65x�:v;(`�a���)�,BD����P`mkCo^E�Z�x���ɰ{3N��6��g���T��5�� �\X��=�qU�)H���]�_P��@�R�d}���Nޡ;i�g�2�%�Kr�Wm׳�m��C�  �X�m��E�ڥ�b[,VѭTKU��U��U��Z�jڌJ��ʖ��
�Z�֭�F�\2��L-kE+B�ֶ�R�m��[m-��h�P`ڪZV��FԵ�FV��m�ijk,R���Rܲ₶Q��ڹ�32�iE�J4˙Ҕm-IZ���mZ�m+��T�Z4[Q,��Uh�Օ��*V��*�W
�Z�
+1�e��PF�eVV�ʊU�fUAh�ڍ�2S"PV����imjQl�dm����q�R։YKe��.\�R�j2��h�j5���TKaZ�U�E��-�Rc��)ZV�V��ڕ�j���8����E)Z�mj�Ң+rej�6����4e�d��J�ѥ����h%�Ȫ��ڋhڭ--�R�G�R�@D����u��w�*Yn�k{�j�_����-��/&u.��w����ND���z�g�p�Dn�:��ܱ�;�yՍwa��|��Fv-���}ݵ��޾]V��'��,��z��*�z�6
�Gؽ�6�K�|k7��q��K{^.�)�P�C�z�3��؞�Njs9��͗��>�c&7Pk��B2�89�e�9��4^'�E�H�ms[�Z:��j��}s�����}��u�bp�2���udC�U��w���V��!���	P�t(�o{j�G��k���r�Y��0�<v��V�ӹ��	��SQ�-W�/'Ý��iV9��[� ��������~mn����5���7kE����w,Z�輐����ƅ*Ħ����`�����NZ�.u���Ш�ow";6W>ۍ�.��5�.��g�������+ީZ��	��3���[f���LIM�D�<�3r�^_gr��貟��1JN��S	ʍ]m��E:��f�T���x;�hX�G�}����1t0=Ji����dI����~��m������c�ϼ���&g��-�e�.���8�!<�U��>�Ì�'h!>�B�zxok{��8���i�j`y�wWa��B�_QRj�xx
�Zo~�y��X�'ZK��з�����P}:���	
����>we��ш�>��S[�m�8y��uh:7(�U�K��+���5��j�9/nt�w��^���9�O��m�v��e�Ŋ/z�r�:b�߈\���UΝ�٥�ҁx�4�X�5���S���6�]�"5������.ΉSWyd��o)���UAj�Yا]7�*ݷut���u��IͶ��&��9�����T�[S#+z�75�ϫs*4���w�Ym*긤�����[��M��ګ��TC;�Mœ5Ҟ��([>�Ս}Ќ��v�������o(a��m*�1ݘ�z��T��9�]7X��گf �Y�*�ì{��W8�.��ض�S��]s���ڬ�d7��:��̑����E�Z�p%&�8X6-���l�H�O�9��L�h�9WX��^r��S_^�����_C�݋N8F�8�.u1�^���7݈3u)y$�_�����s��i��6oP������`�,�Ь�����wu;��ݦ�����t*'؇P�n�Q��LT#����}-g�4H���`�f��6�p~���-��[�������;&��������y��V*�&�+q������uD*鬖�J���t��TbhW�ݭ܆���;Ify��O|��n2���ٰLN��g+߇�h*���t�o�>��$�B-�J�ۻ���uPzk�$VM'�wo�f�mi�~9������u:����ep�#����V�53�7��X�喚kr��5i}�׋�>�'S���b*���{�]��*)�ˌp��������p"��j��=��1v�o���>5�/�4΅o]�O��8yׯStxp�bg���w�O7��k�V�WV�{z�5�{�^T��#��U����;3;1�����{�Ǩ�p�5��԰�冤y�]Ρ�)�t��.��`a��^�D�W�"�}��.ǥ�NiMv�ٕ��&{�U]���IF��ww��gS̯VCh��9�	�C���gW2�̯�q�ܯȵ�e0֬z��}����gk<U,����+w��F�ցK�d��&��xfdF�m.��-��eI�H�h� \ꌚ'{��ۮ� ����,��'V�Z�M���&-���r�q�5G' �ۼ����X��vC��	+zjV�[
k�,M��\�7{���Ě�j���ۮ��lAu�*u5�Sz�T�ÕO� �p�M7�r=}����3u䭫fTTBp�y�]S�~�ǦƯ�x�
p�)�0��lsX��n�1�1�٨n�'�2a��V�̡TYwCoV6��MF���x^L�W�.�u��m5	��D�BS9 �Ӟy��շ-:�'?�jZ���'k�.�S���o�1Q�/���ҷ-�\T����>v~�lz��*Q@Vr�����S� �̼[=]�f�;w���}9Z��k3�
-�ې�6���.���,M���vj��t�fvj�2r,hT�:<��s[�>����*��Z'�dye�	����\����hp�'FG`HR�� ���o1��N������n�~�x��#��T�-Vt��޹YwJ�Ne]�V��Dέ���p���*�����6߄>1
Jch��^m�h})�cs��N��Y�2otZ���o2�V�Aya�{Iq���k�mY�ц�C�<Pͣu�ѳVwlA��Qh�'m{�[�1��4������$��@O�㇝Km�&��U1S��%j�\9��ãj���أ/ӻ�s=@v=���p{������g�t͗|'v=�v�,�ŏ�C���/��8��DíR؂���KS���U�8M��X����Tj���r�x��ސ��Y�OxsI5�y�O]�zy�dB�u��t�k��W���X�D�|Y���z󽥺���p�S�������S��w)��]m���[ڂ�tc�}�Z��F�N��������N�u>�FV�'���ym�s�MpU��+�p:��c��k�����9���y�P�(F
��S���n�9Y��<
�}�=C^_g�u��*���<~K|>o�i�F��(�K2�u�nj�4�?j���h�42|��k�_:ʖ�o���;�����y�y-'#�ϵIjL�}]�ц��m�cO�٧��#�r���Mu����|�gj�g!G�N 1^�-�dI����q�㘙�3�q�w"�ѯ^��ul"c��S}�8`�ޤ�֏jSѳ�c7w,�/�V�����{�k�h�T��Y{�H���y�����h��i�4R6zPJ���kz(���w��4{E%#�~�������l�9T.u��ϛ^��F~e稫��9�F&�_k�����	�5\\e�qS��*�������Y�gW��~�}�k�6q8=�i��֣�&;е0����Qy��^�c|�
U���<��ɻ����5��,%�u�����k�|7c�­�ں��K6i��/,�m�d<��r��TN����+��4��7R��+n�+�����*��CO��5��:�Q�����	8��������w�$�h�K��w2��I�y�s���=�mU{]��c��t����Fk�+�wLE)᮳�Y�
u����wWO���e�v�oOu)�f��"C�z��s\�neDiO;<�z����iWV�ua@��L�FV�����ӛ�[t����kr��4wYC~7�5f��7y���"��L�-YҶ� 3����ƪ#�v����*e�,��.���p�+�S�p���v����M�q}R�L�����S�!���9�R<z���:�����B�����pƣ�1Ub,9����5Պ�Y�[>�۳ݒ����ע�l�����ONX��z�����:��	�6� �rWe�+cfD���R�E(N������g8Z��**��^lcu. �=��%m������Yk`ޭŉ]*����b��<u[�	�p%&����������X�[ysy͛Z��Y�܋�s�"s��Gd���z+y���Ш��h�45�l�M����)�^����^����S��iQ���s��bhW�|y����Z�&�S��;�K��,�輠�e55����9�O:��A,�.59�r^$b�t]��Ѯ-��&���ͪ+(:�t^&*���L�sq/�r�K��_����_�MnD;{���u��|3��R`9&c{���������hT,N����&��,��W��Q�o<T���P9�5Xǐ{7��v|�-��+M�چ�	�C�a���fժp��F/x�[߬�y&����M��u)��}����:U�:�p���Љ�H<���H�/0�����yq<w�6e�Euz���%�����vo+@ջ����ԙ��Ƃ�ݜ������^�~�~Z�[�q>X��㱩�cXphfҲ%��Wf���K�p�-��K���{{��w�:��fCp���\EQ�'�z{���%�3���/z�r��U�׸�ّ���R�L#fj�T<��%[���Mӈ�꣝�Q��O�ob��f^�3�6�U���H���m��:�'N@���'��Z���x
�<+��>�c�[Ӓ�m��;31����uVt�׼����)������n�.[��u��`ҵ��T�t��[�\������veNk�Cj�1P���Q��-��z���x��{w��K^lM\l�ݒ�M��uQ�	�se�Q��-�ɫ�cie�'p��w�R]��-�n�;�\��**���������42t��4f��^e�
Vs�&]Y�ghF^���
�Uw�U����q���Tk�����d9������F��vR=zҮ���cn�n��PJ��R>�ؽS��������U�U�^]e��ك� <�M��C&qj�r��s�u�
ә(�%L�r���w3��+�y��tkܻå�I#n�x�:�l��:b\��J��}};���wA1̧�GSRu�����7�&�Eg�՜�(Ҙ���pצ�k����B�C�w���H���g��qLW�c?S/<\ל��I򬌪�Z_��%����U:Ʃ��N�Os4���}��P�z��v�}��}�+��{Ӄ��v������yq���O2�Z��17��oel�mc�|���{ ��4�����X�$�߂|�i���Ծ�̨&w�$T��;����ڨ�E��+�bo9�f�$
�o�l�����z���p�rg��?u��K.�����-��<�w�fҬ	6z��}3w��y�s��*��������ه�{��p�@�v|isƘ[G��w�������w(���T7�;�긧�P�è�b9�N�$b��;+6Mj��&�B��aLV��O;�M�Z.��]�oC�^x�Q��]�-31�he����H//<�yJG�x����ϝ`�o7o<��2^�cV�� �y{����6�j� ��m�Z�3�P��T��n�H�˷�Ű�����}�]<�[b�(
��Q���؈ey��'�棳V�q��^�zŗ�����{��4�WSk<]���{c�֌��'�c)Y�9�jn�'o����8�J U���k�G|�W���C_rͫ��Y��3=�j��sV��oب�Q��ӵb�tu�ՙ���-^d�&��<�M��dRѬ�S|��'���=Nܺ��%��Q}��W8���a�'�0�6g�i���B5�\�h7K����v2Ū���yR��ak������6�n�&�����Ոr���hS����k;r8c��.bũ��Y��"����+�u�FD^79ʢ*�I�z�g�� Ng�+:;}�b�O�f�֚��l�b)D�Q���:��_nQ����X��\�s���v�nXʅ�pa@k�Q:���	S��Y����n�D��7V5��뀚ˌp��m�4e�(Y�s�<U��,�Լ�$�ؽ�3�kױ�2�H��2�bԛ�αm��i{H4(`�8I��k�N�����gr��빋��h��e�c��p��d5)'��}� �$A=��E�z�>غ_vOvn��.�f��*�C3�娯m�X��;I�<��i5$)�Or�j崖Y���w����g3��cK7�!ͬ.9w^v0yu��eT�ŎVs%^��T��r�vط��:���Cc��;LY�f���M�q3�,IIc|�ݤ�վY-���{��kG����d�p��J�r�]��W��$u�'��[%Ј�6���Q�\}��ُ]�Cٝ���y��-?,�W�*�u�ڍ�(5إ���t;�Z�Ϝ�v1m<����uچ,��a�3=�L�:gv@����K����u-[�YIJ�]6�����8�$-����ѐ��=9�RT�i�K^��kW�2�����d8�fB��P��5,3M��.�L� ��1<3b�֎tk_tΧ����p�e�X;�[��ڵ�3x��bj�X��
��¤k�6Y���4m�}���������xg';���m�ˉo2�ζ�
Úx�!]Qʊ	��c�t9&�K�2�ta�d��z����6&p�UN�Y)Rљg�T<e<Y������g�z�ݴ<d�G}9z��(�2���)����C�/��L*�����wzQ����z��d��jY�A�=r����x���ݧ��new8miucx�;�޾�|lnj���s|Ep����t������]��.'ʲݑ}� *uEHm�݂G��\�u�]�v�ޜ�7�V�tɊ,�����r��hkt��:� �Ҽ���݇�e6z]�'_4sI��55}wx��mX`w)��)�at�%	��9��ն��4�q��[V�\���$�$�0������o�ZE6#�j��̮O���o��R���E1�~v�hB;Eo�tx5�$Z/�]�F�>���if�|�v�f�U!$�J!/�;�z�R��I��z睞-�Ⱅ��/l��!� J�;3Lb�o�oR��ɋ�)�^�v�͟72�X�N3�X��u�q����v]ԽRd�^`���XݱSRN���a뾈���ӭ�B�.cF���+����ܹ.��T�ȹ%q8p��oY}ya���g�R�b"��M��u{:��6��4Ne2k-��as]
�l���J:�&�l9��.��{�7 �CeC����Ġ�Sh��(�$�W{�eu8�0�y���Бk�����S�9t���-C�S�7<�WO@�2\����(Ck
d'Rܯ�z��񲔶2*��G�*��ˁ՚�4�,�� �)��T� ��˦7x���WJ����������w�xZ\��`��������=TW��k]���fC�\�[���HZ��M[F�DRؔ+eQ�V�5U�J��KJ��iEJ���D(�VѪ+k�V"����Vŵ�����\L��(��,h[h�ت+J[`�Pj5+hTb�eLUZ5�kKmEm֪Z�V������i�JV��J�X��UڨєBХ��F�hֲ�V�)���Z�[TD��6��mb4�*֬XD��Z�ij-Z-�lA@Pqh72��Jң��R��k-�)eUX�R��j*!��%m���PlKE�Z�ж�Zصb[(�
��R�EEQKJ"�9�(ը�։KaYm�-�\e�)h�Qb*V�im-�J�lA��U+YU�F�"-+
ѭ�
"1���ѩj%�h�j�YKmebUm�֢�[lQ-�ʨ-h�,���kTh�
�Xָ�p�D®4nfiR"�ie��5�&2��%�̵�aV�bZ�r�#Q\��U�,mKXȫ*�Jb@� �%Y*�ó7�v.۸�
X�ˢ�.�/jl�qǆO����Ӯ�8ϯ
פ�kOve����⵭pYיǥ�J�CO�����D{C�V�k���z����Ƶ!hc��ͱ�f��.�:��ŭ�T秨�|w��9�{�J��^Cj�]���B�@�)hH5����G"�����([�w��E��>�7�)�u]O�,�����.�<���o�!��A��)��޶e}{�^Ҟr9�9�)+���K����֗c��6�)b_vA�f����M��e�Mq��oa\{f�u�♜3�S7Ϝ�m�Au��'Pۢ��]�X��Ta�*�'�ţֳi���Ԉ�h��lʊN�62[�w��՞+o.��-C����4mV�5'�^�b3]Sl	�s�>I��Bp�T42[���H��0�B�0)94�.�����e���';�d��z7��M�`�47��y�tɨ�|�:y��)�X^tU{|P��Sު��\�*147�U�|��j�vb�S�ެ�O.�.�LM�Z(m^J��Mbg�:�!��ݯu�U�	�Y��x-wԋ	�2�y��]\|���=�h&�<.,�=ٰgSܙy����#( ӹX/��V�ǣ�GDJ�J����~���[nIYW5�_�����.�����MO�%Ez񨨜侭=%z�m;�����>)�Ӻ����B�<V�W�+
�����}��_K�;l	���w���Vk�ΔsWͦ�<��$'��/�l��֎ �)wpKṙݨV��+���;���p�zyJh*��r K��GR�]��Y����ԸLv�օ*޸O��p����^�G2�w[yk[�1�6'Ú�I���Fi�N�s=]��ľ��m�,:�i���J�H(�p�è�B9�����xg���7��įz� N[��ڶ�3��W/�X��"��BV9��
k�P�e��{_���ƽ�O��K�{�B���t�"�U����]��,wa��_)����hf���l�;\��c5o+��!ps���yM�p̽��t�9� -CF���E�ઈ׻X���ߠ�b�yԡ�̑nȝ�.��U�b�:�2�w��(^ڄ�ve�+�����<ͳ�=�ϼ��ޮB:A�Z�(�E�db�����E��y\��٧��r��\��1�L��175q���QfL��v����WMJ�ܷ�e�KSu������T�y�QI�بm�T�7��)�]��Z��Nu��5�n}u���Vbs�-ʄ�H���^Nt%s{�*Z�\���SD3����B�V�V�k|)�Ѽ�D<�3Q/���WGen�];���ބ�<����j���`'ysJ����+Ԡb�lF����M�s��5�eFsB�Z�m��>���+z/(,u(�54��S�ŵ[z�� f�ml8��K�e�j��z5�1��/<�Kk�Y�!@f^5��h7���Wz�ڧ
�����یi�t�Ղ֚�.�
�_\=�o�����
3p-��2�����M��-V��ѽ�2�&oD����+�p�¡ðaY�u�J������y`I>��5�c����$9{�O9w�N�߷��<�~��N ��i!��f��$�MO,?��q�Xu&�Xo�>���|8{繁:��or�r2d)�߻B�^
��˞�+��g���e���J�iƫ}W�Mu�����Kp�*s�U�<��XVT0�{gd��픖��WG�����s����*�*)�u\���aU�f�|ME�!۱�b���ˡH����ا��,\���M; ���
��7�6��xɩ�aԛx�~>�,'l�=��	RO���5䕆�KN�Y6��Hm�:��d�a�xh�!=� ��wq�9�Sn�Q���?{d:}�d�'P����C��oO7�`�d��I���M��5>��	XN��|�*
�t��h,<�"�p�����+��$3q���3�����i���h|�I���s���y��N$��y�@���5�᷉=I������M��Bm�I����,��k��{�D�W�ُ\��D�go�)��I�*N��6�����u��i��u=5a�J��}��@�O]���0���	�ܹ:ɦ ~�rN��6���#��ퟪ@_|���&z�霾]���B�=C��~�J�$���J�l��I�O�6��	����Z�m���ԕ����q����4��&��0���"'~��w~ e�uu����o�D�OY��0'�|ɠ���L��?^~�J�$��ĕ��e'>d���	���>��a����֯%JȜM����H���2���>7�!������N �7��z�Λ�Rz���'X{9�$��I��M��<�N2m'���yBq���>��N$�ec����?��F��ߔ��#��G���$��x{�:��*y9�:�����8��T?w�B����kO?�d���9��I����m�?>����֙Mgl�E�Ϸ��_Dh��{��1��I�$�=�=O8���I����xu�T��0�'�5�����>eC�y�>d��S����O=�%t�q�~���7EM���)՝�o���0z a4�3����Bi=f2u�R~d�d����$���7���I�?��q*S�r~I�O�����2m�8���[��Ƈ���I�nVS���],F�G����eu}�Pܼ7�L�{Xn�|��oS�7�C����Yjߝ���u���;j�g��T�{Ml��RJuC��]��D� m>�������n���X33��4`x�m�a�֎��T;���l�q�'r������;��N8�m?0�v��zg'�Y�����]��'Y5���d��=��I�5����$��r�d��	�?.9Kp,���Z�E8��P�����2̟$���{�'�O���ĚI�?e	�x��іq�zʞ��I�}��N �jo�%IĝeMs�	ĝaë�G/�'��Κ��s~K~�"ǣ�=�'XO��d�O�2{��'P>I����䕓��+&0���d=O8��c$�����I�}��N�`]�G�c����+;�{�]8���<D}�HVN0�)�i'Xn�:���'�ޙ�=v��w�'XN����$�:��h|���PіP񓉣)��� t��a�����ws���{�C��d�V�{��6��h~��!Y8��~ï�'�5;̝I��'�d���&����+$�;�2J���B�|����Oi%]���4���Ͻ�E�{D}bG��I��Ld�jdۦC{�2q������
��N�ϝ��2s�u'��~I����'L��w����l���?w�ǪE������ֻK�G��>b �{D-�>I�jaI6���La8�r�̝2�`q��=v���|���so=d�'���u�d��O��{��/+3�q;J�$W��X��л* {����	PP�n�!Y6���q'�6�p��d�i�ڒq����'�����0:��h{�0��&����}�Z�ڿ�Y�9�����x|ɴ�@�o�M�L�a��НC�O�w^�8��{��*Vi��iY=�|ɿ)�,'>O�:��{�����}���~ff��s���{��ۋ��c�������P��O�?�AC�O�Y����'��^�u&�?y%J�y��
���FY8��'|����d�;������l�;u�}t�^j�4[	G�T�M�=Wk1�<���D�t�vq�|s��b�Cq�k�H��E7Ӗ;�&^Ҍ`�j^f�Z*e0���N��*�)5��9b�ˮ�:ǈ$f+]�u����H	ךw�5J޾�5u�u��g����ͥ���o�f�:�j�W�������9%z�L5=�:�*Voxu�Y'?v��'R킇=Ag{HT��p�y4�u'����T�']n�d���埂�?�~��_t���n~����G�p���M�|�5f�Y?2qǶ��&���gY%J��{�8��+�9��8�����8��V;�!Rz�����L'���%.���������ǔ]���?{�H�M=�I�����Ě}LBu����d�'p݁�<d���a>B��t�$���a�N%d4s��q���[\��h}�����K;���'f��2jo�I_�&�SvE'����Y&���톘q��z��ԜI�{d�8���~C�4sxu����f��k�r/�ʝR�Im}=�Y���:���Nr����M����I�&����ē��vE'�Ԛf����ԩ�:Ì'����'P?2z�Y8"�[�W�MP?���$�O�>�{D{�w;���I����Y8����p�'Y6������O�|��}��}�'�2i����!�>d�k,�$�*xjÈ"=�{���e��QK>�|��"(G�D �?!�M�g|�m'PћÌ�	���:����{�@�N?$�w�I��>s_�$���P�VOz�d?2�����j�]�ٺ�������
qorz�'�Vw�8��a���q+[�	Xq��Y�hN$�3�;�$���'_�&�zd$��Oӽ�:�=y�d���}SM�Z{g����-)�q�U�Yrm'��!��J�$�3�P�	��Xq�iX�	Xu���~}���xs�N�d�a����ē���H��{B�Tq
ԽN`�	�
�OZߝ%d�'N�^IXm�ա�T�Aa�6�̜J���N'���ēma�M�`z���d���y!Y:�����Ę}�5�>u��_�/�xu�/1~iPu�#��IO�P��ne�Ax� ����>d6w�C�X-V���'g���.L�<��yn s���Wײ����/�4�]���]:H���܆> =>=��rԻ0�^_�aI8^�h!���ńTOj���Qw���ڭ�C�=����>�|�2h����d�MO{�$�(M��T�AH�6���J2O�q9�g�'���M��7�@�M���y���n���l��S�5��~���z!G���1x��Y:�d�M?k�	�4ɩ�~���{�$�(O��+&Ҳx@��6�d�I��V�I�}�up�����޳�=�9����B�~~Ht�2q�Ԟ�C�y�>I9���M0�㿲N&�6�O��0'P�&��$�;��IPP�Mޤ��J��0��o��<�Q�^��̌�^���{�=��|}O��<��ԕ���}�N0:��hzs�?$�$��ۇ��a��{��4�h,�<��2^����I�ׄ��&wm>�����3��w��IY>J�R~d�����l��g�}I6��:��2x���p�	Y�4s�?0�$�����N �9�$��N�u�;�}��5���VV��1f|�ο�ǽ��eG���s[�M��<�N |���זCl���i�$��`~N�i���8�VT<=�N��	����L�AHy���������k3��{տk�}����C<J�gw����O���L��?s�IY'u��d��̰�i?>���!�C'�<zɦI�}`z�2u��^���P�z��xg��7׷.������4��@�{������ܟ�q��?N�V2y߿y�$�S�K��8�t�OϬ-�I��?�4��&���N��O��z���5���~�����{�ԜA{>�z��4}�:��z��'Rq���}��'>J��{�|��&����d�2{�O\I8��R~}d�k,8�zΧxg��_y��������5�z��	Ӕ��2q�_����Au�I������i�z�ygRq������N�m�'5@���t}�R�p�F{�c�$G����Z}W�ud�kSEgZ�0.���f�x�����T����VC�z��٫�[�9x�%��*l���X��Y�8�m`E���m�U6��t�B��7D��S=f�2P�cZ���9;�ٙB������ޘ���xk�n���4����������c'�-k{�B0{�#�46�|ʞ��0�kx2u�_���N�My�Bm�k7�L��?No'Y9�����'Y6����q��O\��Ϭ�_ʧ�;>�ݪĹr?z=c�#��La����2|�Ͱ�B����
I�ϰ:���!Rq��SP��	�a�9�]�N��y�Y;���X��TTa'탓{����h��G���}��'$��<���C�a���a��!�<I�je�I��k� ��|Շu���l*N2q*}�rB�q����oz+�㜧*���k>�=�X�c�;a;=�(I�O����8�q��d��R�iY6��Hm�q��q�|�^Xu<d�te�m���+��*L�v)�w�έ�p��{�`�����y;��0�2s��M�a9��	��&�{��T��j{�y%a�CAi�+&�X)��'R��l8����t(�<�l:��h�������{�ma�Nj�v}�d�'_P���`uw�6��Gu�z��'{a6�2l���%a:���גT'����D�����pO�3�]?|md�-\�}��'�FI�3��q��i��;�����I��� |����x�ԛ@���N��6�I��rl�N�s��F�6���f>���W-��4�%ABt��J��T�@�O�8���q��y�k$�y��W�C��q�>v��y��O�M����M0��ߧ��E�y�=2@��p��Nf�kW�'�i%���6�f���*T�ɻԕ&�Y<�N�|ɷ�^XN |����&�zj�RW�C��q����4�����d}�+��M��ќ�\��ɶ@���P��s�'P����<d�a���IR��}x��o���)8��'_yBq����>��a���_�����Y�I�;�~ߖ1k)�x�j$�n�O|��ϰԾ�=���l2plmj�R��CuK���O[�h��w-��<F����"^u]U����O8E�y/w���y�U��F���#Ί9�����������z�lB���ՖEP���ǻ�@> �պ������IR��O���u���)�'Xs�2|����R~d�;��d�a���J�d���E��2���I�DdQ����@�kI���eb�����E~���_~I����=O>CG�g%eC�w�PY%O�ì�A`k�����>eC��*O̝�Xx�xɽ��(��y�O�{�Di�2:�ݝt�m��y�T$����P�'������&�u'����.�����}�:��*y?s�q*]�O�8��T?�B8{�=��e!��ߗoP5&����Me3�{�\�7��WO���)??0<�����>CĜB{�z�:é?{d�8����$�����u4�=g�y�Y� ��\g���c��k��R�X;�{��}���`z��'M��>a>`~>����i���M&��2OR�ɪI�'��C�N �~d��u���	����E�{�<����X}���?e߽���ӌ�>���0�'Y9�'���>d�'��}��O��XO�I������񓩬����T�j�Y&y�Y8��ֶc�G��|<D.��nP���ME��3��ϼ�Bz��3�z�a6���d��	�w�q��>x��Y:��O^y���~`s�6���P�����OL�2O�G�.�C {��Kv��������e���}���g��`~�%I��eN�ܐ��a��a�i'X~/2u'XO��L�Ğ�d���a:���^IRu!�C�VO�z�`ud�_�y{w�k3V��>��~���r��$�Ɍ6��6�e�u+�~�*N�s���HVN0���	�M�N�����2I�����!G������!���_{gCck4e׿{����!Y=Aa�`u�6��c	��Mya��m�e�m��jo08��N�Cӻ�
����;I<d���O���'���	8�d~��^���7�fg-%��Jo�ۧ�,�ꆲ26!]����H�Gc����59��J>ur�Rbǌ��x��T�İ���y�Q+�L�Y��#̽{w�d眆����g�ɱozVM�ۆ�+pu.Q���g|��1�#j֢39
�YU�J{�G���u��[\��?�{�cߡ��	�ݝB�m���ğ$�(�m'�La8���:�d5���'z�e!�Xo�ͼd��L����������n}C�=���{�2}�`,��~氕	�vq
ɴ��e�>I�h��q���6ԓ��V$�����a�Rz�3_����79_dNe�Y�ګz8z<�1�ޡ�wI�x��=�0'P�&���I�4��$�XO7N���J��P8��M�MXN2|�~��XN!����]�������/�ml��C�A�4{����=�k���0�$�c'z���(c'�,��rC�|ɣ�k�XN��y��*T�ϯVO���Y8��'|���m]���BǽG�7�;�}��z������&���$��4�^��d�+���$��'�8����r
d���!R~I�{�ɤ��k$�XN��V��\��qy3���/�ϣ�{�(DGޓ�c'�??&!8��}Y��O̜C���:ɤ>���T�?n�Ad��9��8���s�2|����T�����cv��~x����}��������9%t�m��I��a��i���P�d0�Y4��6���d��:�|�a����IS��0�'��~S@*��}f�ܒ��,z({� �G�jHT�2xo��jI�&�d��N���0>�8�4�5톘q�𚧩�'Rq'��'�x��y���/�}o�kd)��L�|Uv^o+��jLU�[����MN�=�lu���T�u<�M�=+�ʄ���f�C�y�yդ�w�q�+�ۆ�vt�ӛUVvy ³V\��=k&lĆe����ٛ�v,hc�Ki6a�����T�}9{tѝ��+-�Щ׮�GT�J/E�ipMhCs�uG�`�����E�8� M"��}��ST��ƏNAzS�4ʁ�0̏[���o}L��;Z\؆wr���^s��k�3h���(\|�v�t�b��r�B5�V�f�ֳԫ�%�;�������B���q5�.V��'��M�{y�Ҷ�ڏ1���bd��vm#��v5e��u�j��HQႎV����!��c�R,���rb����svS�Q�p�ş68�Eꁮu�ƱjPK���Rn{���ԥd�ۼ�*�*�~�<9�(�n��T�	����8���V%��{�;6U��S�g�(I��z��W��Z �׫'�1��*v;��>�������int���
�S�|(�06����C��8���f�eoZb��]N�*|��u���QyE�0�U�X��s�r�o����m�q ��E9~�]�������\�˙�hl:Ey��X��zF˓�r����V�8.<1J\:h�_�f��Z�I)�¸,sʄ��-�!荋�B�ھ[��Eq.��O��ϴs�sQo Pj"{!���Y{s�8�S{�ɀ�nV� �=0����`�)��N�%[�P����X��͓����j!���;�Ͷ�8����}ޞ�I>\�K]���ց�'���h��:�K^�Yy+4�da�j�a��E��@��
����jG���ZwƸ+�s��͹;������M �Evʃ1��cxT8V5O�P�@�S��y;D�t��t��\ܾ:%q,pOQ>���+�H�m��,K��Jr[s�e>�$��K/�!���}{�Y45�9+q�n��@{H}�{�I�fL.��L�["����N5y�p�ʒ�7�3v�|z�m�3���`� hW�yf��s iR��Ǡ,{�A02t&��e��8	s7++��k���u(u���C����[`�N��{�5��+��P�q%1�Ǹ ׻fx��*�Ta�iS�ԁT���	��i�����ϻ�;UëѺ�M-s&H%�Sf�[W��i�\�b�e㆗sn�kk2&�\[��ԩ�<�w`�z׉AX�xP"=~Z�K$T�q�	1^K���;$P�[�M�Ϡ�tZk�CI��1^�o��H��4
m�0�:oa�+�2�<���Λ;@���W�IY�}�{'^��Y|_=�� ���lp��f��;ۭ��W�!����-�F�Y.��Ñv�H��&)�ˇ����KYr`Y�M�#"�h���K�\l��!� �U� ����@�ܿ��5D�-UCs�K�Y�7��3�i�\;��F�������&�7�V���8�*�B���l�I�������;1���a!��׃��6���O�����wCm�q��[�q�-�䲯iC�xNZ�}�f* "�\3�=Q'd�l����џ@�81�)X�j��AK(��IZ���U��
�TTKmm��+kUU�b2��[m��Yڪ�B��J�X�Tb��X� �ZʭRҠ����V#[�,�*T��%����(�ij��
ե[L��d(�Ա��jX�X�"�D�QE��QaZ#X�TƸ�[Q���%�X*��"��j[mij[e�X���ȢƥVZX�1EU"���V�ch֕*	s�"6��1��j�b"��*���[��Ⲩ��V�#Z��b��P��+U�F���-V"���QU
��[P����iQ�Z��UQm��mm(QDDU�EV��R��m\E��U�cF�5)e(���Z��Km���DDmKV�բV�Ҡ�s�E��+`ʕU
���+UeK+m�#�8ֵ*�eJ �Ř�f%�F�mFUb���j�6�ĦV�[J�*�jTV%�q�*��[�E2�j�
�S2�8Ѩթ��6[-��KmR��bŖ�KaA+,j҉Qkh#�q�R�Yl����>�T6��S�*�n�ѐ�6&cΓX�i��*:�Տ�����VoG���2�`1�8�!Ĕ�ʃ��O�������ӭ<���W�LQW��Ns�ʕ�kO�;{��W���j�F���E�vx�;����^��ϵ��G`HT,N����&���ζ����t���v_o4����ez
�PN��p��-
U�v�V]�Ys�męOd���x��'Y��(�����vf}ؓ�|U��W-�a�[6���{�ed�������uc��D��#�z�UA}p�\�SS��r�6�_!{�m>u9K�궞�T���8��9��d�6��Y�򬧋yU�k�V����vR�z�N�z����7b'���\Gr�^bL��b��zV�?Q���%���{��I�{pۮ�������l�Qh�윭)Ȭ���i���-S���;-����y+j�Q^N�L���:�ޕO����No���C`�kb��i��������x�*��.>LA�`�̙}��0�uul���}�B�|r�W�f'x��;��z�?]� m&��AI�X�)���Vu���Ƀ.v]��w��`F�F�޾O52�Na^|z� o�����	��mN[���,aL��[����>X293�}�#���Ѷ���ڹ�ޏѮ�Hd�7t�X�^��ׇ{+wË[�<��C929o�-a?t�P~��&����hhf�����j��y!;ˉ��y6�U���n�Z��jjm5��]��7�ebhT<�����C�騌�)�KaT����>k�rK33�=X���n:"r��7��ж��y^ku���](cK1dU�^�W����Vr�	�t��Lw�9Q�Wk�ۈz��#t,}�9r��J�Ϲ�.
M��P�;�=҃��G`HR��
|�ѹ.�� �F���mo)��I�t�:XT8v+!-��w8���]�`�Z���7��$sC���O��W�^%p�ïxp�ڀՑ.y���o#��55Ëo���WݏjĜ�}�#��÷�e�<:'õ�=� ܑ���]���og�ū�����u眦��+�o��Xu��0���Q�J߱�I^k˱���:��^�r��?b�}4�$꣖ON�[������dWa�a�.�l�⵳u��[웙�9���P�oU��s���6_��\/����8��J�!�����M����3>а��;>K���e�h�$��[��M{��UU}_{9Է�SS#=ٿ�5�O�^TqK;!N�o�u���S��l��	���ŧ���ˍgk�(>,Қ��&��/O�vn��=��]{��/��]�^|W��y��������hl,�
k�7����/y���}p熁U���W�m���2�89��.��`LF��^+\��u��n�r]j��;���Lbq���o6i�QQ	�ئ�7R�X�]su��� ��RD�p�5σ7|�[�~�=�w��ן#Q���~hd����
U�鋗�b�Buv��}4��_P�K��Aa����&�B����ݕ���#(��˹�gKV/kb�`=u��{�**r�D.u���R���7��F�l���SsI�Mv�����쾯<j�P���`j��x�U��e����6�a����kϽ�Ux��0�#X����c���S�����Iu㍂��ԋ�+x����\��]��{:T~�7��EXF*R��^ᛐ si�T7�Ej����6���1�ٚ0w_i�K�8�1��W�XOM�c	$�xGT�]��b�����9�;�%��y+�(��CJ�z����{������y����>U:v9���Վ�����³1��^�j0�u ��R��zrU���!P�9i�����θm��4xh�0�ћ����&{5��5�}^�=Ep��bк![ٯCO��ڌv4����e�u?^�k�Q�(͗�N]:g�dG�c������=�3mLuê���=V�9ȥ�	�zǺȧ�ox��c�3�N��ݒ�W֥^��A�ʵOo]Ծ�n��;<�	��� �s��+s!15�DLܔ��;gc:�u�u�8S���ƕu\RuE�*��	�1�-��[v{�rk��:淆'��ĸZ��ƌ��em���͇5��5��Р�ԁ��٩x���l�KW8錛��|�QI�د62[�{�;��:
ǲ:�v�� WFӈ+o.[���W��X��L$�W�����`g%�^���{�@x>=����5����� *𼴌T$����)+������˃�x�����!ZV׳�Wj�)�2�ٝ�s]��i��]"h��bw��Wѵ ���;�QL�H�k�	^\SQ�����s���� U}�K��.�r�?SDh��:Ag�Q���dGd��z+��j�����2��kfw7[����贆�C�ٯu�]���W'k�*�u$�v�t�xHξ����������H)�|y�U�8*��h��(�3��w�ܨa״^�<A~='������9Q�W~���>܅{����i�g6��*J��"	�b��&��5�����W����G�(歾]���Sx]d�V�b����s4���KQ��'Sa ��0�>����:,��a���kD뵍�W�!��yJ���숥�c�5��+z���QÂ�◹h+�Z.�RYʩ�p�5���txp��^'�z\�\2;z�ܢ��h�w7�]�Ī������<�%��lc��C�Gk��\Q8�,���s%Ykcf����<�b�u�Ӧ�)�T%a�:3�^�8��ޘ�a��髬j��k$b�RP+��S�ME���2,�s�̎3��V��sX���Y�z�Y�!���5>p��c^}^�H�g9��V�R]1d��3:<l[}�;Cu75����Vs�݋4.�x_#v�%��Yz�b6�[{V�<�J�:�s�2w�c�z=�~�y��O~�2�=
}Mg��N�Z�r!ڮ���]Bn�I�ͻ���'g����r��{1l9�;��b�jٗ���or�Y.��x��nw:F-�*cX��+6"�:����A�%m_��9R�[�
�39i@ۤ�%pf��2��X��<V�ק���U���9F�.i�	爎EٝE�	����룮J�r�㡮v%�r�n�9�n���|���و{{=B�t^L�;��P�8�n�t����fu��̕��Z�Ш�<��͏C4"���i��mj5fA<��X�-�x�X\g����P��_�{���Ԯ)��8�@���fI<��sZ~v����)�}��g��W����G�h!���ex,���ʹ�d��/=`M5�+�(�\�����fε;t����#zB�[W��J^K;������
�i��HT|�y�}֣z��K��ǃ����wt]TC{�G�4��֡Q����w[ꉕ/Y✗������x3����p����uG�w�V�M�άu%mMT�c��V3f/R��*.�w�{���M;����7�\�,����*���8v(}��1�GV�ֈ*�mY{Y����=�)��;�	��:���9�����ձ�Un���62�gwr��e11���|��l�BO��Վ����>��ߍ�uQ��U[m��~���C��)<�}μ�ӬWW���U�yC.�Uh��m�{�u�����A�fU�������gg�ۮ�'9c��
1qK���N�.������|���&о2�O�n���%f�{MxJG�\�����Z7����KAu
��'��<��{E\��{0yO,�r�x��7C�k���ۄ�v)��̼
��j�'K����\����~��ށ�
Ϯ��M���EBp�)�����6|%CG�m��r�W�~�h?VǴ+-�fK��`Lg(�QPݭ���6�eE�z,{�9��~Z�zd��^�y݉�TI�˗F���]}�Yd�5����c}J�<�Z��]y�m��� .�&I�VG���Nǵ�1���v�2�մ�3��(iN�!�8����n<������:���(<��<`4����f�b�ݗ�{��G�ݣۋVA��φ��/"++̕ێ�y����n֌l�Hwu�-S\�vf�d��}]���U����Pr�.u����ܞ����`��0��T�|���8+ܣ,����,)�})�{�]`���V&���tz��:='�����׋l�&>a�F�o�,�Q��sz;w:+�f�c'!� �Z��߇5��z��ݸUcbʟF��-d���� ��3�
�	��4���\c��~m���s<fd������WV��;<��^�=^+��v��hR���O���S�k/9����ժÝ�g��%�S�.y5'{��L��5%o����[t���{�krz�w]�av=�C��7� ������i�__����s�4�	??��{��y|���w��p�aMv��̶���;<p>^��9�mL��{]�M.��&Q����ž����d~�Z�ӯ\)0�����U��(��}IAWYnP��9�0A��a��v��S5nR��i(f�j�s@��GS;4����獸E��t�@||��E�Dcq_���ٙ"꧱�'7���ĭv"��I[l�g�N�%�,Қ�?k8�\��P3/W;4���c27V;SO�[~N'b����<
���/��L���K��6���]>��^�6�1��`�(N�y���F�*qى%�uN m����`���O:����u����Rj6W�������q*f�#����}C^]X��t�����xq�-��?;��?TL����g��7y�(5sݭ�����	�jZ���kݩ\���譱�y�3�t���P�������ku��j�k/謐�Wd&E@�Ok�W
�w�;�~���޴y��M
x�nG����y�Zi�����=��_ڱr�ckj�nN�S��LTNr�ʕ�汴�C��V��3��m*ٹ��\���s���&)��LW`H,O�
|�7c�ݠp�$���sP�Qȶq���	3��d�B��؜N�8�q�ƅ���qD^j��;S$a3_-W�j�	�48�ۻ�	WRXe�H��^�K^K����Vd۠�S	�=�����eE�T�+�l[���<����cf����(Y�8p,�#���V����EA��YP����T��']K���;X�*�ZK�����k뾥2���5�4�=�{�y�����g�,x��N]u;Q���w}�'U[I�b����7���a˽���7��]��)��{�9�EN|6�s��k'�v�w׏>=�֔�3˹מ9V_v^_mؓ_�ȧ7�q�(���k�K2�Gk�C���k:T�
�7�<�U��qJ]��qP�]t����$u��s���Z��$�bVu3ן]�w�LEO�����e0��cz�@Ԛ�/'"q�m�ǹږt��r��cZ$��g��_˖�9�~e��f�4�Ѡ�,�F%L;�uu�aZ�J�e=|���(+Hp���D00��BGa����uW1�X���vz��z��ns�	�Z���P*�ZM��#j!͊Z"�:��Q%͜��i1χ+�9y�����~�0�����i�s�K��vp9�:�t�t����#�G�ר����"��y��y@�!e���~ޱ3 ��r��D�����o̽�2���!FR�b�Z���]h-�z��mƆz�)�8����N�mX#����<����۪��Y��͌*!]��m����s��g�ny����V�m���tX��Њ�n���x������X�P"h�\v�����k�5��%������2�\��`������e��������V=W�K63E�UF�'���ר��c?+�SM��j��=��jU%�����ݼ��`�Ļw4�l�k7y����yM^$����n����w�j\���΂��<+'���eB+m�"ʅϵ|�a=�Sf��,���s�n�d���o]֬�xyjb uN^x�71}��ŵ��}7x�(�wX1��-L���߈��t�u+gb�iL�hZ'n��@ps��@��W�����\b{/{+��3����x���~��Yܧ1~'��1�ه���:�K�I�ʅ쌝�86���=&W4�Ga��a
�4�i����������UŹ��Y'�Tk�HzMI0�Z��G�˶>��V�E�Uڸ���N���2Q�~ a��m
����Gs�Hf��>�̄�]+r���7��8@�c��gw#���gD��cm�f���#(�/�dkrGј�4����{��������,��5w�>�ɮ��V���,����D�z�w,�s��9X�8��Z�fV���1���K]Dʵ,�o]h~�,��֭�%vXQ�c�TJ���v�a�	!�֧t5bm;�=����Gkw�޺��.k�{��-�;͞®5V�U��~��1�Ν�0J�b���]ӗ"����Z�p\�����vt�/���|K�.}M۬ipWrY�6w'��;i]�O(	�o�K��AI/2��ދ����IV��Vr�V۸�i�(���N=;������H�AoEh�!�=��W����޳��д��ֱ��Qf<lظ�V��Jȁ�N�-m�i����T��[�w��k/�h(��<�����r$�Tn� �t=���Wڢ�ݮނv^e2��k������\tH(��f|���˦l8κ\�0wvA\�+�ND׾�{d+�L�i�uù��jW�O��j�r��%�Y�b�99��g�A�V�OY*��wgXG*p�u�� �B��X�]���~�]%X��H
>iM�{z���swt�F�Y�l���=ocA�xҘ��"��kT���]��y��{t��~� ��12���k�5V[���p�h�,=����F� �a��̶�:�W�wSxr[��0 ]�Y��&v��u�V���-Щ���}NNS�?q{�`�)�QՖ���jƊ�Ie�R�ZpV��ynd+]�i�⻡Й�b�a�#B�y� t�P<�>���a�0`�gF_?szu��Wm�km-�Z"���T�@\��K�fX���(,`���ic*��Db6�kJ��V�X[YP�iF����.QU"�[R�r�Ŭe���h�Lʫh�\�ո��J�ң(¢�\��Jѭ�DET���J�l�ʎf��!Z���T(��*
֪5�qE���DUlm��J���[(���UF)Zcr�+��2�#[kFڵ���L�A\�kQ-lV�E���h�Z�GL����hX�(�
��b��V5���"��5-V�����c+Z��eQ�Z�ң-�*QU�kF"��F���ت6���+�����2ƕX�ة����XVŭ��A�*1Ve��G-DQR3)UAR�[J�*�������#[cbX�����ب�U�-*���#��Tj��-�(*�ʅ��B�U�r��
��F"�ܴ�`�"-j֩[PW)f[W)*傢AF
**���TKZ�[FV�Ѫ�5
��meH�}��	�,^��i�Ml�G�T�65+}b�s\�#���t��q�ژ9ĝj��[����b��0� +�ʆ~�DDz#��ҙ{{��Ȏ��qhs��Ō���X)���\���|��d�<v>�P��{N]י(�$�֕�RS1�5=8T��{4����u���2"�4\cN��	'�{N4��o���˚y��ֽ�f�d��VR���Lu	x��Ϟ>�����'�������^]�K�Dᆒ��u����xi�Uyh��@�����|�H#���oK�q55��'�c�7ǀ�1a�Rҵ�1ݐ�0�/�	Cngh�d{ꂃ��ʈ��a��ͥo��l�jJ<o��b�},\��q>��v�	�
bʒ���3�e%u��}�zs7Z+�c���e�j8�e���Yx���Z��B�Cw�15��4aԋ�w�˛������\\Y�d�3EP�1]*���f8:���*�֣�q��.���H˽��r�_>�(��� m��ԦfP�z�]e2<lR��v�gl�W.���/_5��g`C��nkV}�ء�Gh�X ��4����P�����j��_��
�g]ZD��=�����:7���z�{ݻ�O^ĸ8���Y(?1�h�x�h�ݝuu��`棏W_��XB���i���YZ���n��گX�Q�S7�Ws�i.�;�;����s&vK�k83�2�0�o^���oU���r�K����ǹ�K5k�Z���Vxb,W~�Lm��&儑A�&U�]��]�Տi�bF����e��\�9��p�R��6�v#T��F�a�q.��`�+��.��j ��Ƶ7�j���e��}�p�\+��c�$�)bCwj�!��tF��X��p�37�����.�7Oy,�"C�cl����y;E��tI�N*y����GIƤ���݌�g������t˲��g�⌄&ˢ�F��"Ό�y��^�f�
v���}ѦoH��_���~K�^�,_��P\�
�4�D�-�V��c��|��⎀o��3=�h���vF;��;�G[Z�8gg�x���ΰ��*z�P{gO�h)7��t���#eC�:����vp`L�7U;���C��O1,�3��X��[�7�}ռ��S�_�����OxP��@lo�qF��ɚ�N��V�Ƭ��c�~Ub�_�I��w�Ϭ����MV6ծ��c���],�HH[%�e��5x�P�\x���l���`*�cy����҆S���Ŏ�-�%wh�����U�%/ɹ5g�^x�Kmz-�֗[��]��5\gC�ȷz2��'"5�GP�4����ϔ����)�_
2@�>�r��W��mL�V3�S},�M.�!�Uم	l�ث�^�������t��M#H�����0
T̮�3EWD�҄ŠM�d�<���0y��t,�Nr$�&�
7,�K��DC�.I�a'��R�f�j�Y�.��}$9Z�MV]Yi���]��eM�-%�3K
�F��:�ݘ^G@����kjp� γ�|������C����9����3{zp�z��c!㧆�g\8z�<t{�l�r�&��!	��.N%��ܥ7ά�Ky]��핇J�3���Wfb��5*�^Z�,\D��b��D�9<M�FA��;[Ӕ��Jƹ�Ќ��5űP�.x�Ƅ-�Un㐙�	�K���}ׂ��fFR�ׄ`y�;���ۛ��\&�/�JdRP�+>2�W-�8촕��q�9]�ru4�sv�py����˪Ė�V���uQ�,�K��5.xf�z��9R�x`tku����{,�b��=����;�5İBRFSyW}�p��;g}*X͙b'J=�(��|7\���{#5��Y�Nh�^��VsVE�ei6�緷:��."�@B�ڶc=��F�h.��݋����+��R������e�g���ҁ����� ;�v�Z���^����K����T�<_&ƳD;�9��n GGn��S���Vy��˦�Tç��n9��tv�L\h�%^����v�B���1e����(Ͻ�G�b�]o��1SqÆI��+*1�.NQ=�yHwo�F��𑕓!��W6�)���簩�<����R�a.;eٕp�9Q����)a�K��d��ڭތz�yb�3Y�hӁr��+�.�V:�`/���{�J���K'���Up�t��	��{ڹ1-T/�R�>��U��(�7R�V�3���N$_��'6���؁{_�w�-���Y+#�]K�pW��=*�D3�D�
��kȪp8U�D�;��f�O�7��'���w�X��)�!���+���0�$x�L��I�-"U�BU�AY��E�j��z�gR���i̦�/�mx�g�yO�T3�b0�'%@�Â�nnL�D�ǩQB����ĤV;�9Uw,E��;��~K1~�t`	�iu��h�lS����*�jI3� t�҃#�+�S�:�E@����<�f(_�K��62Y\�i�ܜ�D|�s���S2�X팘MO�B:Tܱ͚�:�tB;�`�+�zOG�
!�	�$=L)w�]�/i���B��W��]�7�-��ܳVjY֝=i�^���M��0ĸ�&���b�</.�kTW��=@�d3�d�]Z ɓ#�0d������}kY�S:�1�pݕ���ޏG�[��5o�]C���N��Νz|:2M<ഖ�h��k�S	f��X�����y����v�����Ε��}�j��98Th�}�TG,��p�=�o����?
d%������qnn�6D,[PKζ̋f��^N%i-I�f�"8�4^W�B���"��v�ѭ�Ԟ/� /cC��)�s�(�'n�3a6Ց��g]����{W��9� �`��NE\�a�l�q���1:D����9�v�fw�ߦ���q����ɸ�"򤳁�]!W�H������������:4���:��"� m�.iN�Z-d��WӢ��;%��<"��*�5}4͔ɸ����{��$X�ZV�Uev�]��n�����k�a�ݐ�<4��^���BB0
޾v�{n�_QJ�u��x8�c�*_:
u.1�-+^S��0�,�(m��rf8G�T9�<�*��;����1�Yf�m��x'����ȍq>νy� �ı�T�D���R�^���(�^�C��d�N��̒�1x���W��A��Ub�;�W8�
�0�u��
ޛ�.
���P<*=��yv��Y��.�bZ�\�\|v&MQ�'�EH�������OX�K��_���ʌ�<������(�u.�������+�*����k�*�����UFU��j��Yx��Bgx��q0�Tc�Q����2��TqS���|֔x�H�p����Z�
�f:�qR�Oz���E\;��ػ�F��N�ײ�e�oH��\���37�j$�13P�*%�2�-J�����v�C :<=���{ݗ��6��g]���Vo��x��bx��aةp���sQ­b/wqj��i��u�u�I��tts,W~��:��tr�H|�+jw�]��� ���笵���]�ֺ9�-��3���!��c������pXck���08���]1���˵?'Иb;��.nI�϶뀴��퉈�=�����q
�7v�Zr�n��^�W��jp�%y�A:�׏9,6d��),O�g.��W{x���{��&�S������ǘ��7���p�<g�ܡÞ��,��������>_K�����C����w��s�vT��YJgo7��hԬ�%=���qW�p�~PsHf8gՅ�����U�c��86�F���,n�ܿ^՜��wZ�z�:�.��ͮD����:��Ŝ�1Ro^����z�+=i�jH��o��un��l<ϼ�`Lm�T(��RA��=��үg)c�ȟ_]-!zIW5����{z��}WQo8֠j���W�ׁ�3;*{�)�Zs�Dz=炞l���9˱�Ɔ�jȸǕ��~kVD��^X{�
xv��<�)���'������z�PX�[=��b��3��|�z����<ĳ�m�=�h�W[��5���w��K�E�/�����R����)����t*�x*���$!����� ג1t�}�&b����|��],Q�$$��,�����-9�%G![�Zv�:�m+X#������w�T�W&x)s!l�D�Z&��������ƫ�^�\���;��+���Y��l���"y&	/˟32�QB���~R�ǭPR�[ش,���[C/;��5�5hP�o�h����of E�a	M]�(9yn�7}�Nq���:�w_0;8�t�c[3���]�p���yn��.�c� g) 	�o?�k[^e���Ғ���,�L(>g^��TƦgD%�V��Y��Z�,\��bðH]���R��٢6u�%*Β�&P�'�nD[
�x�׆�1��*�a�T<vuZ3��4� �������$����v�\0��7�n�ۧ:�2v���l��y�}�rE	]�y�M}��W\�FH_�5��T��#�ziʮ�ue/�?86VSQ�{coi0ݑv��r�dw��1EG�����WXtF1�%)��Ώ���N��#�_U}��S�-f.�q�j�g&I{�FٕK�E"xm�,s����Uc�a13� �p���Y�[��~y}��� D���'F�]��(����x^̡F����DL���/1N�%��ٖ�b6�࡬�P�J SRF7sQY��8at���,f�U1�.!F����=���)�S�3�^�p����ZM�DD����}�*{;�lQm�9��G�����n鎹��c$�:ʌf�p0Tbt���yHwo�F�槄�����A�+��йŝ���-L���	VpWQ�[��`��q�X�|[Z'���tGϭߦ{}�D�Mik'�X�bՀ��z��/ѓ��byU�Ȁ�=5��A��pD�/ ��h�ri�W�W���B8H�/"]p6T���Al�i��ʅ2*ܙr�j���f��<�c\�+��2�]�bΉ�D�k�p4(��َwz�y�G5K+����;!�ʍYO��q/T�=��tHb��XH�G��'e���j�7gr��5gpڭS>���R�!�.�N֪y7����t����j�n����ؔt/P�����n��s�T8���1�輽o3��3��ۧ;�udO�'H���LU���X�Z��y{/�^����� ��q�f�����D�dנb(=�}d1P��tcz盉A\s�!�b���kA^��n���W�d��|{����`W[��U"������9�pvW�����LM�6e�*�u���0):Mzg���hK�!��iq�tĺf���zrJ����<�ګ���6��Qs�
�e�	�%�
�X��ɀ�*t�f������F��MpRߔ�@���|��i�QqX���i!u���r����ja�,�Ƥ��.�I��t�v�u�t�N:l1��"���a��2!��	����^���]R^���q�O8]�����T��Y����m����J�n�6�͊\",��:�gF�u��cnz�u�����ttO��[<2Lf9�'�yEA����3a7�j��O���w<�b��˽e��X��mYE�R,�
�v"�P�E�S#gh����q��&���<J�e5�`�qR���uϒ�Á��6�m���"�g�\�w�HW�{4����;6���Zܺl�:���mm�����j뽰���`ؑ	H[�tC�Og����^��L��n������gK�0Ұ9�m�]�-���.��pL'���U���;�ݾ�q�y�16�nq7�p.�v����8N�c���#���S��)����Č�_W�U|��� "^�2���'��������4��>Ίl�+��������w�y���+�[ ���}�������	ꦺ]�7W��F���kI&2
��S
nNb���%9�i-���_1�9�1,#~�:�O�S��x����X�^w�Ca�wV�#'������`���?=�������KS�G=�'����A͉A�Q���So5s���0X�nfx;��S+��	���Ie�we�g'�Boz��?~u�yC=R�ԮX��Bc[����W�C��HP��1 �:�;kyz��9�q����'u�et�{�N+�vP�%�T�;�v��j$��)���Cآ]��G�{�R�Ґ�XM,��(��j�X�$W�w���+7�u��@��'��J��
��q[ǳ�ît':{+j���8\ju��7z9��a��%Je�,���(>�ʱK�;��,v�:�J�Aym󽉢��J�rt�w:�)t�1؍R�N&�E�a��wv���Ͼ镵3絔 ��5:�Rk3�\���Gxq��T�V���1�\ɂ�9`��~/Odg9�iC7��	�	�3��y��t�|���0-��μg�X��n�b=�kGj��^��ϧZ��!Bd����Q�T�W1�OpCה��̲��f��tR��cBy2��L�Nؼ�;W��� }�<���X�X�[ɰ��Ը3	�*ڨ���uZ���l5gn/d�0��L��^o(�qvɸ<+��m��y�Q��v���SP����/��!x�IP^�bN�E���d�N����I�{� ��ZLkˠ�t�k*l�;N�\E�9�^����wI�t�<%Y:�߹]�����ޢU?���w;q�(*X/��<�DwK�h��Lu�mg:{���6b�Lu�Rν˘)T�qc�E�����݂T���$�\��twׇy0�� ��{��E'kn�
�
`��I��y��ž� =`؝��L���V����`��d����^e��w#��\b�,�][���s{�2�����J��<9T��5���L��ӺB��m��9N�d�I60�թy�̺|i�[���v^(9Nᙍk[��jn�>�7£w�I�|;��,f��&оv�&������iܰzphӸ��3/���֫�U��Yn��;l��4Z�H�N{�����TrO bի�k���W��v�#�v�7�f�w!tvB���/q����G0�w��8X5�4�9�PUk[<6:�۲��,!���j���f�m-��j�H��^if6x��>����=���p�o9MN"�=Ոm��+*p��G�}h��qZ�Y����f�̷����\|O�+���+��otKE���ƵJ��/���g�19��:�[ûO�Buٵ����B��c�� ��WC��k�|�ƒ;��y��M�%[����X�nW�O��*�}�WP9er0Wsܻ���X: ����W�H���J�"����r&�ͣ���k����ԑ{�cܹ���Z�7z攕��5]]�}�H�ܹ�-�}Yc��oF 6�M/(�-[4 8p�L�/b�f=��M0��6�X���'8�>��Q^W��ѷǞ�b��?��ul�0S���i��g�ɱ�Z�	~�V�C$�u&?��[��k�.��Və��4���u@�݁�&�\s_YEd<P���Y��h)���a8��r��z,j�T`�7�'��A~��r��J&�VkR���ћ��^�;���J�[p��5KV��mX�l�<o�X��Z�m�ufH�J��U�������+��䲳s�]���Pu+��K���p@�Yy/��E@VV�2%ɩP�dʒ�u��PZ��{���z_6���ܭ/$8J��\�1ѨF9�]��]*�9���߻�_<�x���R��J�QrوP�(J���Ԡ�J�JcYZ1X�+%E�Q�QV�����m��Eb��(Զ�EJTʕF[V*�DR�D(Ve((��iTUJ�UD�l"���VQX�Ah���
��T���PUQUb(�F	T�ʉ��[j����*��*U�����UE�U1D��T�"+R���E���kPDceV�F+UFҊ�J�U���IR��"�R#"5�X�Dej��b�,�h�-�DF�+ZEUKh��,D�cF)Z����+c"�Q#T#��"�(��**���-ZZ�Z�F1V(��("
�����EEE����������1DU��VT���1�"�(�"����Ŷ��1����F(��bDTAJ�E`�Ab
)��*�Q%J1�(�E�Tb��TF(����TV1E�*TE����ر�""��F*�������u���o܁�S:=0�m���H"���>@�B�s���ٸ�a36�3�)y�����������7�������S|�V�m�,f���,vV�+!��f;�Mz9K[�P6��E��#m7�x�r��v��Zj)ܢ:/�n,�
�P��k���d�׋���$�w
�u��Z��q���+69.?Z�}^�p�ۑ�֍�J��ty},����(f��"Ό�L��� �"������� � BU=��5;��W�&�
���8h�rd����UJyԅ�3����1G�N�u�f�MQ�Ц�T���ܹT�QL��-]�=���O/EZSkܕmת0:��ҙ�++��D�+83�2��=T�n{��F��x�M�\�nM������{�i�~��e�`g
-��_������]�Л��"A�Y-�h��TZ�͍��yO=w۾�#,{��"�JK�)%��?0WK W�$����Y�_w:Zq�c���[;�K�	V��(6��e�%P1r8NY�Ɏ���ҟ�>K�Hv]fM�e�>+��{a������9/j�5���j���a��VD6�6��ȝ��3�/.��^�:�J��.o�}�/Y��`_-&MG$nS��c�n|��R�ݾvM��w�=N>�}��S̥�sx㊀I���f�� Ц�g���b],�K�W��f�$���z__tٙ��.�̜o-����56�H/�w��J+�Ս�a�^�{��b���u3{�"���O6�P�V�f�)+^Qz��!<J������U�>7Bu��q�$���~�{^�tƭ�5���o�e�x��r�D�<=�6M�)J�'�4����s��o�9��!����:��f�[!0bl�R���Z�,\K��"M˧7Yl;�g�����E"�-K���%/����E��`�~3����-�	�A�����F}��O~O�RQ9��	f��$��ȍ�>^Z)?��qx�fs$�e��` S�ۺ�����@|��	g˸xQ%�PV�s�7"�
T˸�X��i�H�����q<���=�Az��4x4@�N% $^y���5ŕ�V�������뮙�gbڏuӽ�׮����r�_�P�kz�+ؚ�%C�L�s"��1u[b�t�/��u.��>�5�8��e�ۻz��e
,c�qՕ��F'H��yHwk��¡��#7�wkqS�Qy(�n/�7XT�MH�7q2��V���ڧ�Qӕ����R�&��c�����L�}����7Av�cw6�Z���,�Ø�<_&�}t�l�1���V�~s_Z<�_Z���Ο�Hu��s��u�dW��W������W�ޜ�<��c*WNw�u���Mt���p�P:%�U��$�wJ���0�����S*μ�ڷ�G�=�nu7�b���S�Ei�5*%c!������" po�o9Hi�];��WK��]ZXA2���\;!^^�!�I�.��Qr�O��2B�_$	��yC{���}�U���t���-�Ƹ/:Pa��UvQ���c�+$�k�U8*B���u*���f�Ps	~����CO*40�AF���s��
���<ж��tWE�e(�o�.��'ٙ�JTgfc_�]"cA�>�yʨs���n%q�,�/]� m+VLJ=�*�2���X��Œfy:ATK��q�)�;K�9]w,E�����ţi�nU.yU=5�ɩR��сP��J길�0�f������W���tț�~AײJ*�w;�ޓvݡf����P}��@�HĴWS2�P'�L�j�u��Q���B�*�!�}�t��Ʃ��ã�.���L<
���_˖�8߆��0�>�3�9��oFm���;����j\ktB�6V�8S��P��u�p0���~W�(��w#���YuK��Iu�d��ɔ6�kx�BW��P�����Y��Va��:k��F�����ْ՛�a�jmX��3%	�j;)���2�P�bw��k�뵵����V����X�ƛ��o}���k����W�s�o.X�il�V��J��	"�s�~�ﾪ�.����ΌB�\.0���f;�j3��"٠�Rq+IjH�hHaB"�<��Eb՛�2��ܫ֖��.$���(�5J���;h^�X԰k�±�����Y�LGN�sf�4�=Αfw�s�(���Ѿn���U8�9��z��XϨNՂ�}J/q;D⹖��l�۠��ɼ�f޴�ha���;H�Z׹�YTPѽ��U��H��������V�{�x�2(�]y��W۩�*��&^4�qڞY��5X̵��K:)���-{��ja@�7s��)�۷�mn�k1��S��T-1oU5Ӱ�X��y����Mj�^�-J5�A��L[��CSU��gxx��\t�b�V�z�K��N��~�Դ�r��y�1q	CxW�Pn�2{�/i9�:Or��nm+��[PgL�d�Q�-���X	���׮5� �h݊w��n��Ϊ̾֗�%�@��{�Ҍ�4'.��t�_z<��rq0����Qnc]~�!�����	����)���AC�*�ߪ��-Թ�\F��|wa�W�>��r�Z��In����P��R�ń�6���fS��K��Vu��$���ճ�����2m�y�S�5�C���S���D��;�K�[�-���OZ�z���M��z�`zOV�$�Q[{�P�n��j������Mm�G�j�(�3�U}��sӢ��8��ˑ{���H��f m���R�#�(�^��'��5b�h�ΌW�����)������!��y�t��r�G_ޡ��|i�b�������yD������O�g\y�����;`�F]��X�"�N���C|̀"}�zH0b��2�J�횗�s��v�T8��k���Z���7g ᪚�ӅX�,1�.���V�o.A}�6�u�bG�/KG�9.Vʵ����D��J�Ԗ�q�:��k|Ж�˼�y�'Yz�ưJ;l����P/����pw[V��/�Ή5�T[�@��ˬ{��c�\�mΚ�U��M>ǘ��m�Į�l�}���/���T�zeq�>�Z�k�^۴�Oo��2��S E'u��S�n�qW�p�p���s*4�/;�1�,3��ҷ����&��26'%�����VF;��;�K�:zx3��v�>��� �aP�%�n���{��b�{v��ܸ;��2���+M��LF���c��8��,�`̬�K
��<����fX��	-��Yܒu�v5�b��ך�D�	Z��b�(<9y���r��Nۙ�-�y����
9yM�y̔�KU,�\U�au������c�o�+�ĩ�5����8%��؋��}�x�'��16Z^�?����B�{�J,گ&jS�c<y�Ӟe5Q��:xS7�����rW��p6U�����K�)%�ҟ�O�	��b>.����m��!�do�M9���9�,�q,j,1��E��'p�K�
�L�W�~lq>�GX5Ђ0��М�ob*��w��/1���^	C�������ʈ���6��Ȧf�u-C�br�Fꥐ��u5oK���b3"Q���6rg9�><e)��E�]�F�`�SK�Ùf�L�o��g�f2.�:�(]�R�[k���c:xo-�p]��b@1G����ٝq�I�%3����&7��ؾ���K�����V���֭�9��|�44�zf��r�g� f�ԚWUt��o��ڳ��8���f�4OAx��q��m��y5��ƕ�Xmd�� ]�I>H�qyh��K��Ŏqx�}�̒�eg7N��?%k��<[���=��=V{�l
nNo.���Ib�����j��˸�V-2�N�ہS�NP�=��i���giИ�ͧ��w$�� Wl���:u�FB��T/;��L)*ð�[Srs*�o)���u0�\#v����r;��90���F/+w	-p�*�r�sX�0j��S�9����mYa��y]��B�F���.�Xsٺ܁h���������J T5$cw��;�+�b9+{}i��&p�愫��U����7Ӂw^��2��x�����B�vV�mQ/on(_`ʄyi����uq�����k+�L3'}W��6��a�*'&-��.
�N�7�)�����]�X�"�vq>r:yIw�˯^�5�B��i�.K�^���
QS���;�̅,"Bw˰�d����ww+�N/m`�r���-x��.ZE���F�'C W�'��`���k���RZ���>�� 0�Z]�Ѽ�/��g�y�.��	��;�p� �
�WϨc��n�Vq/�!S뇐ewm�Ρ��v^b�hL��C�/�T7��s�Ɵkت�!7rF����"_�D��Y�Thb�}hd{\K�9ݶ����<l&i��n��s��\������OT#y"#U�Bz��C�C�|�r��c{'<�J
�YJ�/��^
̃-�v��Z\�� o�0P�FfXN����iH���\xw��9�\F	�ZwgR^�*�)<���7Iu䒝�RTIx�Ӿv)�c���<�uv�j�����1���^עȩ����Y�h����t��gf����y�֯Ҧ?,�|�Ÿ�X�$�w(��A	����[fH�r�-ĳ{���b�L	1�,r�<���>W8T��:)b���Û�h�J%u\\X((El�s�Y�N�R�����N_��c[�ۅr��t�v�ъ���.�akyfy4Gז�ixnU���i6�Z��y����+�ԍ�ĥ��ac5Lv�)�xS>t���ђi����G�o�G+��#�{ֲjj�vg��8p\���y��w��	�D��V�na���T+�|z ��im�[��U�<�T���9Rq�y���H��?,W@%�Y���ّl�P�������sb�Ý�R������FjG^<氂b�)�Rt,z�g�|W�S�2�~�9�+�P�l!��A�޷S4.�R�|���0:����T�P�����t������<���.�����8���3O�SOX�ao��0s9��y�+�z(E����5R�k��J��?�'�KX=�73�s �s��;6��Mz�e�u4cN�J�s�nΝ�;%���(!r*�5�\��ʗ�^sMN�ݵ���������A�Jwc2�Zb��k�a��ȼR�f�f�-�W��yV�m��!����R�.�s�89 �3�,��b)�Jq`_�u��z����}��I�
��3
/2�f2�(f8C��+o��>`���ɛ��{�x4\n::I��o�"�����tԏp˚0��6�/��iH�6�7.��U��d�	�n��??��sĬ������`�{������=:u*�0�Q�J��S��0�_5���mb�l��SH��VU�Ÿ�J�"�aC�P~�Y��F9���G=�'�ؚ�����9֒V��pn�n��*�*��˪!ت��	���}%����C4���T	�3m6���-8�b+���Wg��rB�C��G��Nlt��a���{��M]Y]��r��ײ�2܏��nV�h�%�ޢD�vb��ŦO�T=���fA�y]�mÈ�<6����v�`�p�����Jͳp!�:�'��ORV��ɫ�[֫3P�*�_:��N�,['N�:��5X;��g�y�+��S�6�݀��`��ʰ��;�ݒT��p��N�]�j�����u-W�}a�GY�?��S����ǎ�y�3ٌ>vU�[�����`m�!�#������:���a��u�R,A����ܴ*�u:�}���yf����.b0�)�|8l7��&K��=rO̝=٬�"���Jy�:�o�⇶��{vqQL�ئS���mCڑ���е��pmެ�;���f�:ëO�W��D�p���K��gEb�}7���.���h2R�WS��2ȼ��N4;#4ͱ-!���tl���ۍ�R�G���_�{���QPj�p4��I���d,���H���^\M'Ւ����y�Fnv���[�����C,`��v�,�N�h-��b����8XP/N�1��q�he��ô�S���o>��Y�������6�w��^B��S���.U.�^|����������᷽������cU���n��ܸ1��٘)����ei�z����Ѻgn��Y'ڱ�������۾�;c�t��ˤ����%��(P�B��\�����fq/�y�y���n�nMf���#���Cڥ��j,䤰>1%������ m��l�in��Uv��X�v���%�&)�]KNk�CQa�j!�@f��w��Y�)S3 ��3*�$q<���zczm��k��-lH���/ ����ןi�0uYm.I�K��J�����Q��T拶���q��T�7�����!���C��Y�4���k�#�]ف�Cž}w�^�b�篧��{�
غTP<]�R�Z�z��Y�2:xo-�e���p�죱�ĕ5B(��ɬm=�`�����G��Q��cԆ���QȜ�h�.���h�s�I���m��G6.�Ѽ�Vqr�h�	,��L���ٚs<`�� ߶��t�a��ZA]�v���yPѬظ��c/ivbm�`�zt3:�f����в��ś��$��(Mי�7{�ZC���:�k)f���8+�:!}]��b"-�۶��!�#���T6��g����v�r��k���<��"��M�|:Ք*�<V�wd�=�K9��ǯWR�QA6�sMI�7u�i�ʁ�R��U8!� ۻШ���C2��N^sַ �[�Q[N�b7s
��q��9�P#v� K�z�7���V�v�k��2�۔�/��Jp`��WW>�	�x*3�:�S���c4:���c�$��L������f��\�Q��X׊�v*m���TK��@ ��P_j&5����r�V(0Gw���n�yaT�5Z󎷌�����'��u�_#���V�:����3E�$pV��!��@c�r�Qe��	���{���ţ��Qӹ���S�9�J�o3h�ݪ�$)�b�;��wHc]��v��B�+g)��݅��f�;\��\sT{�I,�*,�&�)|�
�Ҷc��S���C��jܦh�Kɍ�Im������ym��pc�z������p�k+_.�����<�9N��S�Rf��m�8�Wgi� M�3*�R��z�"�F��B?�2A����z{��-��CU�C7"���n��i��	���(y���z��Z�J]`�v��K���|s�<��qoX�P�L�T��zk/9��u�a�7��6��}�0�#-�֞c#��rn��ٻ閻�!�]`�ݕ����k�����]n��m4���x@�]���ͭ]�gt��fV��h���S�p����}��NӦJS�z�K�j�j��0oU+x5v����j��#�T0��7r�g$.�E��44D=�f�W�(hNzQ�\C�k�ÚR�G��d샆��ݍq�gA�V^����KO^�9�`��[��Uu���m7.�a��d\k[�d�p&9NT�eI�S��=�����o.nf>�7��S}e;b�j�ȝnM�1�cuE��ڽ.�S��Fd����p{ly�Sprx)�<f]�zEn^ީ�޿;�����2�leN(�&Ž���{���-�d��۫���n'���;��˛Y���T:�(�n��ef;�FwT��о�She��b�΀op���ch)�g�E/u��̫���[��*��(�ǁ]L=�
֣��"���g=B��D��k'ǽ�@Xi�2;[Q|�.��n�b�z.T�Z+����`:���nGD�	��N��8��JU���v$�`��s�ww,u�Kg+��^�=��	�18��Wv�������]�K^�3��`�R�V1�����T�(���*"��V" ŉUUQ�F�AEc�ZU�����
��*�mUb"�*-�hQV(*�ZJ1X�F*#F�Z�#�*(�Ȃ��(�F1U`"�F1AQb��"�+[QbȬ`�DEb�Um�1Q���*��AEb����F �`�UETT-� ��b#[QU��V"�*Ԩ��X�H�U"*�1T�+Q��b�#b�A�R(�*+i`1E���+�����UU���EQkEEb(��TTUQ�UDDQQAUEF""� �TF
�QT�,U�"��"��b��,�"��[X� �E��X���ADX�b#TTb(�DTX,DV�*"EB�EE��"���+A�-(��AFDQb��EEQA�
"��ʹ��!R��&T΁�ӷ���"u�r�������e��5�"<����4]k�b�=pČj�}��2�����Y�];٩� ~���<Ƭ��D_	�;�Y�|vr�"O�*僥LO8�㲫�]b�V���X��%>L)�4���Y�}�lK�khi�q�B�w	�z���᱓N�IX��:�.#Kþ��5���=����E�eyh��K��ŎE�PV��F�\���/7S9�I��p�R�~N@���6q����eX�PV�s�6eו�T�����*R�*��;F�lE�%� �F�D Rq(Pԑ��U�1Y]+�f����8x���	����w�P��|��]���V5���KE��5.���ۛ��d6&��<���u���m5d܌��1dM[1W�P���*.+*1��\�N�7��6�'6�}r����+W��{c�E���%�	s�����BU���[������s�뢖lh�9��<ėZNv.�ӱ���������蕌�R��@->��� h��E}�o_]��T���\(N^L�8���W���B+����gº�X�)LG�%�0��j���{=h�sЙ-Wk*Ҝ��s�[�эs;�&d�H;����S�P�K	��n����1+MZ ������F���q���1e%�����Bݗ�r������9��t;�Y�DS�������7gu�96��O��f`����z1.ݐ�_1�ZH�5�l����T���R��dk�z�c3��0���
�%vƂ\�&�q\����c-�([,�Z%����o&41�>�2=�%��=���$1�S�8��s����r�͹l�L!���_���5)��1�YS�WB����KpP�{�.+b����IR�#C��P��E�$��t�����`uR)�Kk���s,;C+mQ��O�s�pkRW�D]8�p��s�L^��2Q;,r7還O��k��O�fg���I��*��K;�X�����U������Y.�P�r�ܻ��p�Y��!�炫�U1��d��nc�����Uoo1��JzqVS<�SrvS� 9���
��OQ��5�#Ь>���h���zj�SOf��b��)�¶f��8��[�chW]���M�źөΌ77ސ����$��m'8�L���K,Dݪ�W���"�
pV����H���U �0�Vw;�,8�"�*�H���;6r(��v��Ӵcu�a;�*bv�j-�=q����'�"���j�����ר���έ�
x�Ԯ�W�;<�ve>��3��i�!����ռl��AH���N��t2�j7�Ea�1�u+c�΋�-�б��=nG�d|8�I�o]���-]�_m���h�mB����%ԫ#�q�Y|s��$#�t�^� ng��s��4m~ ��o�ӄX\EȀPy��r�^�0�gh��
�<c>�]@�AO�����q�a�=^ɘ������B,�ֽ�9TP�����eÚ�"��{A\�g�u;�hm�D?S�
�U��M�;\v-����to�iq��ȳ��5H%z����x�9��/�h(��*��w��̆������ג�vy�dh�|j��s���e���j���=1��0�A�T�\Gh��N�J�Ō�N��>��;�7ulvh^<���[su՝��2F�gr�m<��E�\(;
J��(��6�B�c�u���9v�Kh�_
.�U�\��[y��+C�)J#�T�RD?
��dN]��:\� i�i^���;����m]���`�!��cs�14y#>0�$=n��A�*����^꣊�u3z�d�c�y��;-�[壐��z��وD�6�b
�;묨=��M�^-�m˚���B0Vʥ��!Upwy1��yn�����A��Ho{k�-B�*�A����DZ�MU��v�[.���)�w3��#EkQU�i�A�xcxr�#Mf*��wΡ^�b�P$�uM�<x�2^Ҝ�Î���'Gj�7.c4>�ܮu&�7ӻ����lL��y�/IЗt�v��߄���F�lR��,�H�6��u���«�K}'Mw:��5X;��g�C,W>���z@8m¯-h� ��Q����IRһ�ST�b5�*Υ�����|�Ȯ�^�p�,e˙sp$l���=�T�y�g
�r�Ɓ�$�GY�(k����TF^�+����7]�%"���E�]��T��M]L���s�>r踆�Ա~+(�y�X�@C����Q{xl�Fmm[�vj�y���Is�,+X��ӫ"Ժ%���ٖpE���m�y}��}}sא�1��7>i�z�-)�6x7�\@�an�{0TBwKA�jw������c|���=�`;��*�u)9��P#$�7�4Nͅ�����VF;��<�Mb���`��t��k��E���5��ԋ�%.u��^���%
�Sv�q���''�l�#S�E����-��Ώ�����i�^��Q.:��Aۡ��%mW�5��b�[�1�3Y)u��]�&��֞�p����*�x'6&tR73<�+��+ݒB@�<�N\�K=��8.��{frK`\�w��2��=jM~����'T��5���%�kZ�����{�w2�Sz�R��`��U�F^�]uꇨ�w(t< 1���;=Cڑl��s�8V�]���lŽ����9�FҦ�������u�,;������3i�G����NV�������@d'l习�<Ӫ	o����p]%O*q\)���B�$w����=�z{�c�s�7�~�a����B\��OWg�DҸH�}��s�z�R�Ÿ�TP�K��Ժb3Q�m�j�,ћ�£���wfN^T;���u��=v�9�x%5<�Uu�P<]�\����p�C|�,c�O���t�N֗ky��^��Xu�n�qD���l�R$�"d!9{�,c�ՁԾ;7�dL�_����249^�Z�VWjku*9n��q.☸��'��t��
�X����u�N��DgYo�ڴCL�W{�
vg��:0�C��X����r�I(vA��tD��QeɓۗN��n�$��k�$�e�l�(����g<�]��+3=f�����L.��\�?%���܆6�D8�i\����׷]j7��B7�ĠCRFSyW~��8a\�g˨�t�Z[�\�C:e��V�S7�9E�cΗ ���"ò��j����j5���L��=Y��lŗV��[Ww8�2�i���'{��[�r^�$={e�O���`�8��뽡�� ������5��ro�8&/:GN���(>w�gh��:����+�w�CQe|�����ǇMw��ى�QP�W�Z�On�h��>1W�P���Qu���.NQ0��j�����V�7���-����}ܴ ��=5�'�p�]T��}C*�
�t�T��C��O��:�� nx�%I����j��;kk�c�*4ƚ�~���n'��0=^�a�k��c�7�j6�n�z� D���<��Br�&V����vD+��~�N.K�K����]�On��a5}��zh<$����`�"�}p���c5ĽS1��/�<(x��K:�7��ۉS���ȡ�>0c������M�e�=B\�e��i��e�ǻ4
Y�=,�N�8�ܓRGO����"ZD8����KiX>���^�/��8�;N-�H�d�`jS9Z�AEؾۢz�P��Ex8T �2�t���~XT�j�[\B�aqؗ���G�RO���u�Ggw#|w��:'R�_�Uqq`�����rvn�`8��v#Oŵ�â�v���ۂ��qǒ��	e��w
��0$"�WS2긺GU��U�5O5�nܮ2fC�|��̗��ʓC2��m	��3���ngi_.�eJv+��嫠8��7V2��|%^�ό���%�I'תP�<���Xl�(<Η|���Ҥ�87X���@�-��꾾|� ����u'�v�غ8��jx�*=���8�)���1��ã�%?/
T��:2M<ജj�	*g$&^L��5��o�]�~��9թ��
�j���l0�2�	Į"��Q.�G�1�P"R�[�Fd�7h��R�-ӎ|߇����%���J%��xȸf�����O��VN15�=�5���X�c��vji�᷊��n���sNъ�uM�(�3�\h�����u�[4kRZ>:9�� �e����<6c~�Ō���9��'��Je;s�b1lL[�s�M��g������2G��Ki�V=.>
ߎQ�nl���������dz�`�)��q��.1�k�Ź�6t���|%���)�3�=��]����ܘ�_�g�#�lFl�M���)݌ƪ����{�[�x�N�27Ӷ�k£F(�Q����B���^�*t �U>,�,w��-*p�Q8�׏-U	ܾĖ.����ABP��L�ϩPd_�`(y'䢋~���`�}nIn��K���yy$�X��B����{Qn���"�j��/�=d^�W��>Ĳb��t����̛TdNjZ�}ֺٙ&���!?�i����=5v"�=�b�6�Eܹ���EiH ^��0p�:�Ћ	��fVNVx�
,��;���o�j\�*��\�r۲�8�g^��sbX�R�Fʅ��UL�$C�Q�m	˵+�����%W��\�:�j����po
��a��=3X���ʅ��AC�۷��Gz-���dC�:�����S[:�pu9dU���;�Y�GY\׉ʱ3�%]�K�����9�ݚ��Ц�IU,F
�T���Upw�<����t��P!�:��oz���5�P�q;Z���Iq%qFE���_I�]ν��n�r����:tƷ5z&s��vd��=|�� E�Re_ԻS���F�i�o:���7��_ ؊�4g.�}=ضxˑ��%:v��a�্�`�$a޺�QC��{p��:\�Lc%��ř�6��V)���p-9�_��4C��0����(l:�IA�eX]��#�J�:K�r���8p�㚢N�b�P*�GI�5'�몡�$�|@�;O��,))��Vs#d5�����U��5�Yс�: �S ED't�jsL�_Jy���r`�(��r�7���x������d1���{ӫn�;��xR�]f�'=���gMJo�1H�ug����V�q��ޝP���\���e�.� q���1RG�b��j��u;�ũ	��s���yC�{fm����B�MT��������A���r�;R�Å�s+��>�[;�٠��
���Vj�{�Y��)���m��pٲnj�I��%�.K:yF��,"Լ��Xb�o[��_��ӷ����س9MN�[�]����d
U��)�]�X�>��z%l���K��/%�R�2��E���<>�d��XO�hP��j�njkUv��zs̠Ƭyl{TЫ�j,�K�*�Z=)���� M�O�˭J�:������%E�~	�Ӛ�P�q�!Ӫ��A:N�sAx-�; /[�̈�@y�9-w=[���4L<7�BX�♇�0��'��=�EB��#�<�4��wkhB�w�w��)^��`TqęC�*].%��"�����
�����F�^Q�`4y鑾+�����qǫP#�#A��jfrۮ���K�j]1�a�p�7�2�y㧆�l���$�ĺ�\�[b���6M�)k�!�hP��c4%��5s���X+��w1�"�7���ީ���N�qq���b�˸�/��$O:M$���C�3��e5�39 W��
	��ˬ}���Nv�-Uc}�4�{m�������C���l��z���{S�ӫiH堬bOh�"I�vh(�+y��,��9���T%uIUs��aa�_8��L|6u���;6�It���q���R)�0����K}K�j�֧#ګ�m��b�v��/\,f�4_��Gbẇ��.☿tI�H�s�^Z):K���u�i�[�߄��v	~�:\��rI�e�l�(����8j˸yಉ,Z�����rP���=��w%��j��X+̻���e�u��7��j
)8� �����+";����QP��*y��ÆL[�]-\/-�
T�S�#��်�~���N���5$�9BR\&ߘ�����9uꌣB�EhT56���g�/f�e?�7\%U�g�|�������'����X���.]��on��ʇw��,��Lѷiej�D�a.���ĽC*�
�,z�d���s3!�����V��IM��k��1�v��ȇ:4h�3/fpm���tx]��{ezQ�	{�Ћ���WXC�S���򫅁:zr��Ӟ�=�;+�+.���ԗ�e%N���U�ǫ���Q��[$-�T=�"�
}p���c5ĽS1��
�
0�)��q�Y����f�1�<GR�PבT�p�R�Z9����F�.
}h^z�����4����V�:�X����E��B*�/d��GFW
��y�J���:
'jŧXLޫ��ec5"�����aAU�Q�Gy�yuU�pU}���NZ�r�p�k���:ȱ)�{�9��@����`�]Ʈ��B1��\l7��/I���##��r&w7+J�����b���鍔ϟKs��C�Z�[=��Zb�NnJ��ۺ�(P�st��o%E�xv�=錛��]ds����[X�`��C�	�����s�����ƅ>�؆��|�����G���ut��lhH-��*Vu����e����6-�2�M瞗G�b;xqβ��𱄼��c�^��r���f�L�(�]���LTm<Y[uc3m4��ѕ>=WPô�#� ��̠sp垸�^�|��Zl��y*��)h�8{`었>�d��w­y��a�'�<!�_r����F����7��l��6�|ouV�y�������]c�I�&l�ր�s-�m�c��8�pY�I)��w3wO:e�W%F��R�˒���go�7ʔy8��q[�!�`�e\�o.��!<��ˣt:���)��f����qp�͆#uZ�L�^��c��/F��W�2ü�b�mh͂��u�m���'�����y��KEJˠ��'�� �����C��ۻՍW)���W�W�����8;2&�e]�X���jm��d�yK�;a�M�'j�x�r�4Vq�7�f����E��"��'f�:�(�g��wt0!�:��E(.�)��fb�Z��_>�W�&����:C�X s�H5��fW���{m�p�\�a�}�
��(=B�v���Ѿ�9�=� �]���kU�ۊ*������Gj[�(bi��ˤO���!"5��%#��}�7uG�&P�瓸L���r`��n���.꿟W[��V�K Sŀ.�\��X=.��+8��4�|4��RO'[�F��z�65�jE�)��7͹W�f�NU�ʇ8b�5����w(�5�Ȃ�� es4!Re������K�)���b�J��*�1]ܭZ�I�'m�+�3W5�����9���¶�j[���v�q�le�T(�.�=9��{Κ��⡗�kQ���i�0k�;y�u��:{�8��7j�vv�]׽�����pY!_Z����/B�v��;�%��:;�?���ju�����嘵���yr����S�
�I;��q�]�ԫ��h�L��l�w�dv�O2g.Qŉ��.[�9u�Ȑ�����͢�G��9v�GMﰙ���&,�F!8!��믣y�%�ں|qȭ��K*�^�LN�H-���V_0��Wk�dT�t+�kTģcj��dŔN�;=bB�6��ӣ 6�<�����@T�d�TyF���%�l|��4������m�2��򮉾�8�3[Ƕ�x����]�;Jg8m��rOi޷@�q���w�8w�$�H�7���g�y�ȰU��b*�"�F)1�(��1QQ@EE�DPUUV*�h��(�PX�*�1X�AUE"��ETV"�#b��EV"(1F1b,Ub#�DF
#�b,Q�Ĉ��+�QQQEU�؈"�"*�Tb��Q*#D�EATEbEAb�E��b�Qb(*",`��EE#cdX�*����,F
1Q�T\j��1UQ
�b��F"�cR�b��T�V����b�QD�aPb�QQ���""�(�R�j#eiD�Db(,AE�J��ȌU�X������b"�DA���j"��UUb�UU��,TF+���ƪ"���.%UV(�EDV
����*"��bŊ�1EPĬdF*��"�e�U
�F ��c���(*�*�Q/^���O,�2�w��طL7�
��^��=>Y������]��n���+��L�t�oQ�������嚭u��e�t��o��H���[@֑+��>�m+ �({}��c��Yz4]{V=9[r�w5Z���¾~�aϷ��7:�Fʅ� ̿��%������w�%���B���JG�8�p�WB�\�R�6������wFN���.,���Cg/2�~�uWfA�{�� ��mT=��K�t�՚�Q���7.�\y����5.x*V3v���M���2e��s"�9��K'�t�*�ac5Lvx���	e��QP��$�,I�br����Ӆl9���Ľ<]SQ�zP��js�Ѡ�?34���W�1�b��5B�q��w9�E�	�6&1O��(��]��e�1q�Vb�'s��!�
n	� [������eZ]���u��0�C�:-h�θ����D��bx�Pofp�b (�a�������iEAz���6��dX�m�b*z�6����uN.���PV�j�Z�s��S�:T�E9��/��=�k�W�f+��c�B-�{��j���+x�/��h2/mOf�-�'�.����-i�[��D�DBy���{|^�c{�^7�ԝ+OU��{�ܜ�"�a��z&Fq��OXX����n\ӝV��**cuS�n�7e�t��ά�
����A�a���щ(�yIt�4CՇ�)� S���i��O��\9�/�]��?����W��.1�k�Ź�0��N�cj�DdͶ%M����-��DaqTѨ����d���;��L,0��k��cv+읫ً���}�F���^-�2���4�0V��8��1gզ�R��8S������ү�Y�ڂ���+#��1ݞ��b����Y8GJ��2T[�������m>lf���{�z�s�͙����s\O��^bc��D�7������rH��L�b�\|Ue�|FYGhJ��I�F�V\'%�x��\�E��1��c}.�L.�`�T/�PP��X�'C3�P���iw+���&aٍ*S��c��<�W�N��3
�{]%���@�`��]m9���v*�k��q1(*�d�����ҩa�3��<��ȷJ����VF���6�ѹ'�w��5䮗j�(T.�K%���:k�׷��n�r��̱\G���f)�����z���;v�l�ԙW�.�� ������j��XF<ʗ~�<��h�uM��r���ǽ/��n���{�7�x_pF�V�t�+�`� �W*t���X�e�=|w�vZ�ڽ����~j�}��x+%=�4G�̈́��}��<�ګJ�-c�M��;��r.\��ƭ�ܱ�[]z`S�t��em�BE���h��FlNNX�ӅYc���vf>OF�!Ⰿ�Hpܹ��}k����3s:'����"������ə��Z֎���׀�>�1���r�����ݹ�[�r�w���a����-=�r�V�������:Ny�<i�]�VM����)��=ķ&f��Rb��,dF�� h��7��j1S E't���x�X�)�=������qK�5�Ŋ���@�Մ�3����O�V`���|X�/�Љ���f�Zz+-�6��y�ӹ�v�ܢ�j��+�-��O�ΰ��'��	���?�����6hԋ���O��x����.<��!���US�K0��c����[�բ��~�"*%k��o���y�«���٤�����"A�X�����Pv���X���O��	:%��C��5�� �H�����>	�ӑ�%G"bC���N�ȗ4�u����t�4�NNb�eN�t�����4ОX&�2{�c�s�0o
z�ϴؙ�dq�]��c�{��o�*�3n���}} ��;�՝�Y��^JKY��Q �]{he����"�m�����z����oWk�z�3�LӇi���2x�U������
�������7��xB��Q��v�ӄ��_A=��L�p|=��\�t��<���7C���V��s<�B��"��!�;.�Y�7ŅE��з��9�Oh�5��R��Muف��J��&&9W����������oz���V;��*޴�:�ͿZ�,: 3��&�r�'�u�!Br�f����V:Tƫ�	�Pc^�뎬����'DsFb���]˩��	Kҟ����'I��S�c�!��Bb���������[5�D���*m�&&c��Q�na������$��#lʥ墐(ך�Y��9�=�~�|��0k��(%Vg�%��XW�(	��+���P�]�����^k��+V�z4�awr��=�e�Ȫb'�k.P�N��{yX�)8� �����QJ�v����<�y�$�z�!�+��+Z��z�`z�<��S.��ƃ^ާ ��Ր
i��$��E����se2}�k"�:c`�����d�y5l�^�B�h����r2���pk�Oo7�ځ��TɼyHwl:�+ܴ ��=+P�R%�	u<���B�������Ԣ�V�'7V2Z޻f�����Qs���Ƞ��!Z9;�F��Ty��U�3^��n�:�v��a�/ù3D�.Q�C�z�`���̜D��Z�o�pū+��}�k����\�È�c-�8�Q�ᾃ'���YU�6T���ap����}�=����r�cѷ�����)+�r�ev+��QWx���wN�/'B T��w<��`N���0�Zq����\B'�E�0�r&s���mY�8vp�p&+�2E��-�~{LE���-��k�z�<cv�=���s��-V�l�~ǮH�j6D�,R��*��^Z%����o&41�>�6qL��"g�$d�s�η�7r���=�.��L��dK	�}v
�ɡ�����]�Ee�*��V��[����N
��Yk� jrQ
ƍh�u�K�l�=�w����c�{��]������UC��u.�h�X)��t`T'%Q2�#~����Y܃E�J;�6{�9�nS�T�י��6p�pW9�9���	e��K��W�	��ѩM�Y�>�4�{�OX�qT¯d�
jx�y�ʲ�Y�1��'A_Wz�*�i��3���sͷ3J$Æ��X��j�ꌛ҅����h�Vx�*�%�OQӞV�6=Wl��.d8�d�p�BN�ӹ������^A�n ݪ��#7'�˗>��T��Yt��F;��aF�g�Ж��%!������R�d ��c��f����٘��\oi8A��\5�O�/&��7[uy	��ͻǯ�Lb�����Q���[Kl�{N9M��us�Uf+�s��!!���9P�sk.�7��,�o
�K$�v�V<s�!��ۋEnu��Pδ	�^����M�8�A74���ns�,��T����3a-Q6g]"¨�r�b��\wf�n�nr���y5v;���N���qQ���&��3��Ã_f�'�k�F�[K���rU��ؒ����,OVG��OH��{�O����t#.1S@��cN�g4��:$ٛڧQ�IF+ŏ�RPh芯#��3|d(��7[H;�N�f5P����Mt�����\�G��O�r���R�rګ��[hX]A���\�zj�� �U>,5%i�s�ڣ��M�kyL`|�=+|���w�C	Cngh�q
P�T�(��e�y�y/6�{�P�ݴ�f�s��40�g��N��q>��v�ΰSIDW�9����Du��ԣ����W'��d��MF���55F�)��G�p�N,�!���K��˒��Dzg92�X�'��=��a�5j�Ci>	Dxy��	�y��<��Nn���qXyڡ=�j]�Vb'����jIo�ޫ���X�T�1�0�.��G�Uڼw�ºƣ�֦�sy��b�{AkH���4�V���Hs���*{W���u!"$f2��ʂǽ�_��*J��v!����\K����(C��\���h{���.޷�KKA���0x=��%���^����GU ��y/��4K����|#���d�����}Q7��AiX�54/@����KS}_y�w�E]��O��{���L�U���գ�/N�vL;�	"��L�{S���F�{MCyԵX��{=0;3���Z����ٍBeiq	�������y�x�)�Ѱa0�]h���0��~�,y���M׽��Rڜڸ$�%,An�@��#�ܑ�`;�b�[6}j�C��}U���54���d����!�~Z�;?7�3VR����X�v��1We�绶j���G۝%�@#����Z����կ�A	���e��٤E�o; �*`�'t���x���
�]�M����-��pŒ̬O-��i�%��d(����3"��&���
e�l>8�v]ji)��E�)��d���;����u�,B([���#�}N������zm2��-Ea�%k�ԵW�y?
2�D�[�<�\(����&#����U��}^���(���v��l×=�[���lm�w|�"�S�v���'��u9
��j�1�OGh�e�e;6h<��zݻ
�=������}�����N�#�7:��·"��R�bwZ7O<�|jƥ���qԳ��@E�"f��J��{]�]+�O%(�^�jS�`s��y�Տ-�m��x'6&tR73<��*sn�l)5�i�.Y�����$r��e��@N������Ӫ��f<ư�u�o�9�ˬ�bp�fl>��t��L�WN�+�h�P�L,7�B���/P�(o����6&#�Jƨ�95I�}�ǲMDi�Lf��fRt�\��*P�~}D7�\(t+|�F��Y��4����-��A
�������	3Wz�/-ڇ)�yd��;7�g�un�:t���7Ȃ��I�8�7�xo"-�p]��{
�I L@�7�VV�{��f�Ï
8|���-��#t$��W�f+�*�^Z�,\K��'����t��
�~�6��ո�&��3&�ky]���K����9���j�E�"��sOz%�SԒy�4�i��ɔ;/�����<�w[�����z坛��P9�����96Crp�ywr��c����'.a[Tw'g���1Mc\ԱV�u�VL|�U�t1�Z���[��\�i�����Xj�.v9:=i���VoDY�}��Y�l�i�]���(i@K�u���m��fY�[�X�Y3Ff�2o`��Z�-|��e�¶ڑt]�30��?%9���f�u�Դn���_@<=�]�\ r�����o�E#Fyt�.̽�H!�+�JְV�}i��)|�S�#�>���\�(�i9�ۺ*{7y������J��{y)�[b�t�P�O�x]�ꓞ51*�Xή�A��s���ԭ��5�'��3<`���}q,�z�oGX�͎���Z��⒒ᄹ���O�-/`:�����ªx-!��Xq`�ك��q/��~����^X0<5��JJ�B*�Z�{�gj �,֦���[-q���g�\(N^�&V�ntoB(����/f�,�Q�<i�7��C8����e@k�u9#�Mw%���XS��K{1��%��vX�f�M�����B�o�yD(a���J]*�w��y*%kD���מThc7�,e-����]&��Uvq/T����CxO@�A,�i⿯���R�W��P��KG�ź�޲&N��B�;��84ۺ�7�s�Ġ�#�Y^�y9(�h�u�A���En)k����{�t�civ���Q��f(���ov��9}�^f��m�j��fx�� G�/��c_���Z�9�#(�Fi��۞�ք�h$z��nS��rW�V�����ե��˶Ik���=����.�2�Mv�����c�iWim��xV,��8��X�y��\;�"��N�l�X)��wF'%S,r=�bK�U=�wR�&W���M�Xp��?GL���UO����q�y.�P�]�qP�!����D�n!c�)�ݝ)�:�
�̼|]�P!�T�8*4���M�	3T�d�,�vk����+��VC*^lr�0;��?k�ס.���ɽ(`��;��v��
ٚDװ�e)�����ܓգ�CN�;�8�S	���?+�Ɨ���U����=��t�HK���܂�z���2'��j��^P1�>�!�:�6�G��+g���=-�hɞ*Mi@cZ��ԥ0��F���X^�|�Y��|��Ȳ,��r�
6Up�s$�5#��X�8yT�i�..�[�*3�J{8���v="�ǹ�7*�|ҋs�n6�-Kb�lsˤ*/f���~���ڙ{��/v���0�	��89z���ݧĔ��ɪ��-��ed�Þ�l�_M��)�q[H2�P�j��'�G�s����!ͅx1~��(�A�����Ϧg���3�:e��oXF�ꋀ���Y��y�+7p-�6R����ի)�d�@�^޲�T��,�%[��k��n��9��o-��m^���!�Z7�v�ewn�k�V�U�@l`2��.���Ⱦ
�+��S{��F���h��iu�=ޙ��ї��P�/�իZ����-�F����%�j:��j
ݬXzem���r;Yt;������L����Ⱦd��o�Ѥ�F����4�'D�Θ��a�:6zn2��9�9�&�#F���m��p�^@�j�-�yE�w1�x	}d�q���6�1�%�����1:^vt���Yף:�]F��ò*��:��䓢N��
:�K���y+��WO�|��m�B�.'wR{d�b]��Ԗ�ޝ�������]LU.�衆5WAa�{/
�Z�2�j�&q�(e����q=e�|�t��0k0$�L8��:��:ϣlY��P��g(��_-�M��!��s���.��=�/H��:���o�uw����.�]�<��@Ȕ	���ڲ�ۅ�@�'�Y����>��lw+ �t�;�-tծ�ޙ[�������P@���֎���2���N�t�f|�Q	��'m�Z�4�=��pJj[���FtD��J_z)�j���gȒ^�R��˦�]���7�:�!�*�������u��ۆ4kfݢ �`�u�"��]�����ӳ3���X��1�ݼi=k��1��ؤ�R��bF�꣖ҭ�zZ������4{lO�bb��k���9c���|�)lq�1+pK��k��Zf,����\�CG��{���;�ޮ�vڹMýCv��M�-�t�����Y�VoxJ�����BF=�r�4�i�|�4�dʁ�]�ϱ�޷����k�)�ࡁ����tp#�W�'o�����@��Ԍ��OZ	>Z[լu�Q�e;fV�/��G>�e��2��������N�iaW3�<��Z��*(U��>ӻ�v�[#��w�2K桎��ɠ�{Յ�|Ec��� >�53��g
��E���V��#�76�:��2g�����J�;;M��o�E�)gI����u��|��)oC��so{���8���>���=\�vt�w&���d  ��ZI�(��,Y���^.i'i¦((e8�����>�[�o0�t����J4$S�v{���D�����W<\(a"�R�_��LW�h:>Ʉ4����-�#e���r�̻ˌ��N� b�wM�=����}y;�5��(uΝ�y�����T�C&M�"���A۾�w6dc�癀��?xki�9L�I: ��}�v�݇�?A{iިݠ�bD��J�g���bU�k���o6֮x[".ѡ꺩w�E��i70U� (1D dU��***#�U��XUUE�X�+m�c����ȱ��c�EADAAX�Ī�4QTb�
�X����TD`��
"�*+H�E��(�%�Ŋ�,EbUX�1DE`��#-�2�QH�26�A`ň�����b*,PFDEX�(��Q"
�iP�k����AF�*#DQ��@Qb�P1�TYmU������aX1DTe���@D[k�-Ke"�F����Dk`��R��*��j*1��cڡw�]���~��T%]�.�jؽ��v����@<�I�=˻��_L�w{;�G�M��xY�݇�n��.���Ψ��m^�Z���Y�j~��c��F�\f��I�1QHj�U�|ҡ�V�y��5],�d�U�sUչ�,�GC��F�Դ�r�����G�(j�U��*��(;P�5-m�F̹���V��s'��B�},\�����wh �`�,�(�>Z*�����=C�U�Y�}�2	���	��,�<]t,&y�q0�Tc�Q������0�����t�֥�f!zL��~����I��1���Y~w]�w�
�{\�����n��;�u�����6`?GN���0PtQ-\��*�S:s����{z�5UFuF�Y���m�ĕ+�/�n v=,EƚWJjx(T/%�q��m����Vf����]16o^��4.E�
�/�N�ۉw`!~�6 �d�9�/OT�.7��޷'N��!�PU�E�$���Yl#�!��kӅYca��:������GY!u;E|�V؇�m�H^��Y��sw��pI���4�ځi�G���4PwRŕ�p��@T�ky�';s��3;
����q�o�0�p�s �l��P�ۏ�;����u�|��r���Gf$q<ҡӽD[FU��:��-n���S�{��8� rko5��p��Y,gG��G܅}2��~�b�dKS�y]�P�<���d�t���Φ�p��`�%����S�k�{xF��b��kS��Q؀��ȵ/ғV9�2��X%>���Xtɶ��Pz}y~�VE�(����t~�L����[�NVީ�e��r���r����,�5Չ��Z��'�9W���O��|X���h@p�c.�R�Iml��c0���GJ�_]h������/��ΰ���R��}B�c..kl��fU�ӕ�_�����9����S��n�y:;���-,gҒ��\�*�'��^�2[�?^f�!��),�~U��Jwla�KN2��w�����Į�Y��X��(n���Fe=\¬= ?V� TvI	��z|a�N�����5e�u�*��c�qwo5s���� �{�%�F�h�Xml���dUØ|��?V�5Nkg��a����r����?�!�K�`�OWe*fR����Y��̇�C�<��C)T𵔎À+2&�cmV�W`����^Qz���@B:������W=%���7
]1��ʺ��uhneD�Y	�D������ȓ�oO&1-����en��a��8c-nm�O����SE�n���`��س��|4��v���R��WLs�+���� 1.�[㪸�@�R���ԫ��4�P�4uuָ ��r�G���t��N��)��z��N_Ӻ]�q<7�n��.�W��+���!�a
��f��
�˞�
No����������S���3�����L�u����>�ұ�T!ҖFf_������c�����l;��^�s��X�C5Q��܊;�C�q.☸.�ѳڟes9eRޅSi��a����e0*,����TI�e���(	��)�8noo��*݌��}ױ�O�I�]G��^Z//��Reܔ2F�u�yP`���.ʵ�I�m���X�i�� ����ʸ�ּ�0���z]��q3��C�.� �������q�I�����;�jy--C�7���#G6�(szjي���448�\���R�bk
�S��������&��!��0h�jt �[Cҵ�%%�	�39���t���yVvU(�D(�ʎf�<��2����j��;kk�g���ZcMKa���ɪl)�ũh�x_��A��@LWJd\d�`
���'�\,�	�ӌ�ei�x�%�4S�`�(�׶5x�o��oTٴv2n�v�:�d�їr��Ɠ��5��O	y��f��A�X.h�~�+��#�B�(��?"�\(;�)�VP�O�`����[s;)މ�D��ث;CƝ`4�v������h�ԫ��8�ר''N�o�^��$r��L����S�:&��K �"�O�D-����^J�&�4Pt���L��Cf���)�T7���V�KD��Y���3��&��&v�.�bE�Z�%��=��v��a3LY�"V/��Ϫ[J�D�Lu�͞��j���oN�o��S�WB��od�q(.wD!Ѯ� �(��8*���酄L��?����f3���}�IH�+ø�O9]w,E�Ӹ�X$�;�H�J%׌�᧘�f�wNf��K+�s�RPc^Mt�zwʧ��\�8�.�P�].�����=��ޑV�<Ӧq#Ir烩�;c& S<N<��YL,f���,:=��{o�b$j�n���Z�t��aV1��4�<�x��K�6���U��Df*!ߔ�a 8ʔ"�㺙���	� ?k�|E��6��b�U�P���k�{N9M��\��>�b��4L��}r��O7\^t������¦���#k���.a�s�%͜�21�P�^f�=��<�u��<5-�h͋�WG؁:�%-�k�.�-�-�ڻh���Oy>�tb�W���ɁP�T���t���ʱ�@�[ӝ7t�=+_'[h�1땗};-��kD�zy�Op&�6����c�(�9|��Qgn�3�<K�c���ot��{ȯn��&��*'N3a6Ց���lb*z�7ݫ������c���z��f{�!�8�9�����}C�ث�R�|�og�p=:+ϳ��a���ys=�r<*�$p�����!��B�a6��e�*h�cN��E9�'�2z��s��wW���qm&p��P�*M��頠\f�d�V��S�:��m#Z�-*�(}�1y3���Օ���]���^`��Ư5z��������σ�P�u��$�j�o�U����k�X�:���i[)��Wd1��r�mv
T*
eN�1�u���&�55Y.-IG��;l�*},YN����y�!��1~*J"� ��:0�)'�b݁����{�n��HW:��*�Br�^�.V;��rq`�F:���Zȉ3��Ҳ��k_)��� �.$=�.��*��-Թ�[ʥ�yNT�"Nֳ�]��ؑ����r�o\�(��� m��Ԧf
XQ.���6K�OD�g�u8�Y���N�Ò玲 �cz��s�x�U+�\7Qb��y��ۼYp'@$�_Bl:��7ĺ������iT"�0��p�1�.+e���ʕ6�wL�7-gk0�^׫�`W��F��^�E������2�1��l{u�ȣ2��ۉMs�c(6*�<��p1ϻ�u�9�%�,�{�EƚW�)��ʗu��sQ��|��
G���_z�J�ok�[� z����]:cn"]�0�儐�&W�v�uB5��P�m���M�{�#v\�Vml��`��g*�-�ȃ�]ƽ8U�1q�:�0��SM�f�#�ԯnWp�\��{����~�e��&	�z�J���%rW�we���z-�#D:�c
�8[R��9V��.�c����)2��:�2Y����>���p������Y���ܘ������6���"��[�:}����}.&8*v��1> `��΀+ъ�Mj:`��2a0-�)�M�����x�y,W~ܣ��PsM5����t*������T����Ð�j�r�D��l��֮ё��Nȿcʆ�T����˕K_E0W��]�=���Ep��u|nm�C���W\���{�8z�����vp`L�/T���n��x�kҘ����J�/'=6����k�U�h�~{'�(pn����Q`���]09�aL�Ƭ��Ƕ����]&�����lV�YP�����T�Oy+�0�J�(e@B:���MM��4�iň�<֎�"Ⴆ�]'�m��G�S/�$ǃJ<����U�A]���v�N���Z�k���՞�fU�r6� �̦dW��e��nl���eLhϬ�E�Fo8�X=;�+�?n�4�	��`
���f������\J�D2�7j�dKꀷc2��f�[��:��n$�ԩ����ĺ$g��E��~�s�!5Yx�|��J\�Cײ�	4���8��0|���&x+��TP,�;�.���}D3�n�\��7`]]����T��/��RV���of E�aJj�A̧J���b|����k�QS�Q���,�IÚ���7�2�<t��E�B� 1X�l�R$��C�С9p�ϙ����˾{��Tgl�/���!�p�l�V������.☿`�<��;�ze6��kF��`5��tj^��Ks�^�X�ys�f�4!��c�Y�F��r(�70����c*���^�8)kR)w.�^I�ݨ��)r�I��tX�΢��b����C�a[5Jd�|7$5+=�0�s��`�6���������E���^_��˸�TG>�� ��z i�����<��
��8�m�$��D[�zܧ+m�5Ҷ�Yk����K���a��g�ﵗ/l�xF�Gt��
z���R���k��A�gV��ñ'X�M���pg�4[��"C��mcw�^��D$K��k=���~��aQ>�Iq]w	�_:x8��u��N�H2_4���j�]�Ta�{}��0��؎��B�[�\���Yq��[[Y�oD������"��ZM�TDKɒ���-�MB�:'�ߊ~5�r��3{�dk��{ũ\=\q�������0V'H�w(n���h���#b2�>"ފ��.9��wcN{yZ��T{������8]zË)�`����%y����z���N��+��*���;���q�ޤ�t2�,�����"Z���NO~����@�I�!3�Lc짇)�K��=��X�WK� ���F3��砹P�S�9�]�gm�烆t�I��.��o���ޕY0�D�S��7m^b�P��C�/�J��}w��y*%sMp�j�^l:M����}�23��X4C9�;�w�O�m�1u�x�f�6�"XYu;S>���EZ���]*f�����Ki��,'��I��r���E�@ΓӁ�Y�3�i[�����DJ���U"����}�s,��#.S���wX~��f��ެ��@fT��J�z�gJ�Z�
�\XȡlЖדQ�,-�RtgA\�8��vb�ӗgwN�`��Y4�#v5a����엜��׆4]-�Í̕���uj��:Lw��y�Gph>Sa�	fH�� a̫d�f	tנF�p#v������35��h��yi��[��u�s�=�=̢��yr�{<g��𢈮��@Y���$4�%���R��vY�I���[LvI�lo����e0���9��hSZ�ۨu���d���`���-P���r�B��M+������ja�,�Ɵ�|��y��=C���gq��g��_"pN8:�t�دz �Ҷ��#��ϛ����?	�|E�n�=��٧�9+7Z�"�}pMg[fE�3A@��V�mQP���������)���n5u��:��Z��v�n��'w�T�N�f�Z�0o�g]���OTr[���T]u�mi�XY�4xl^�0�gh��tEF󊌸��og�a��*��!���G%��^�lz��r;T����ü�B�{4�����u���UB2�SA	R@�{�k֐w~�w.l�+k2.+4Ϩu��2�#�,�8U����ꦦ��L�������&�US��Ku=�v5�zb��S];%��Wq�a��9�-�-JX�
����`�R�9�&��*�t��7d�9��\Y�*_5��N��x����)��w�C℡�;E�C#�'�hw��ˬK�n�JU���u�E��?�O��u�=u���GnA׎�e�Ý���B��]�{����]�r�I�x�iu��ֽ����t¶o;��ą��d���PG��vZ�����v'���z�u.�-܉d�!�����[9�4{JA�L!:�˻�I�S��w����ɝ�����T�`'<����ט��ST�C�5�z�ne���L���r����W2��ʶ��ڽΗ+��Y����!�Tk�Y.V9���Z�Ӽ���TMr�F+��((z��vbA��ʤ�X�y�,�u=�s	{��xR�_r�*�2N�����zf m��Ԧz*\<��|��EXz������yK��_Rk|L��Ryg���E	�U8G,w��x>4ҺSS�B�w��q��:a�@�:���
��n�u�u�K�V~�e����]:cK�(�h�${��봂m��!7V���/�\�;g����}a���p�MS����mC��d���#���-֬��݌�-ONW-1��c�*�f��מ�{����b�v�Zr��԰�
���}�*B�ޥ�8hۅ E���g/�,:�]��Y;E��tI��`�u
�w��<�����M�Ac�\���n\�l&��<~s�;^������F��+1ض5f=��T�X�=:��Siε�+�;QT���EW��̺�-������f�z` 
V1��B�ӛ�"���U�ѵ��1���R��W�\]/ HR�jS:֛�7J~�`�|[����D�&�Δ��Ȳ��K[F�b�C��3U��]	�8��;q�m��蒥c��}:u��y��Q�a�f�Ι`��ŕ�}v �8���PK���H�M��j�$�-<���j�M+�h�I��6�0]�T#��e�鹰}���E�nP٬����ث��q0��I��/��_=�N1�rUy|���Wv�H�t*r��v��t�xgK���i�*��Aݛ�����7L]�.~5O~*��_:Q�t�m��:�$`te<<)�G2�:���Y�8�jr�'	��[+���Ն���N�����WӨֺ畵{���	_y���c�Z�zGؒv��]{3��"�;9��|��A�ku�4�EC�^̭�;�M׶f�v���q<V�������s���Y��S3�Bpwa�)��]"�,�w���|.��3����Y�ŭ}��Qp���Z�V.c��w��]do�Kݤ��:��.�y�����ly~��$Z�����Ǚ�;���^`Ă���|�����4�U/�Van�Nn3��S6� B.ew���q����ώ�P�к��@,K�{� i/���p�3�H:�h޿YT��U!���Q2��3ǳ.,��f&/UZ���5g�W���{&�����uYw�=v�gX��	�	ޖ��2�y��1���]�:<%��v�J�-�_H�����)9�$�"U�)�خ�|�c�^'�{Tk�J�g}2�G9w\-r�8����2�dVA�z�6G�'V�R�d��&nS�̫Y��>tjɎ��`03��j�M�S��:�&���̫�Z�4��F7.���]�ô���T��Թ��gʙÏv��/��0������x�d����`��&=8�����0�A>J�c�٨S���r��>9��=A����l�;�5+�_iE���53Mg�'<(�����Bxy���wZ�C��;y�%|�[�y�a"鴂5��j���ya֜����ٖf���U-�,ZݬI�k�s��k)VV;�O|]=g|�f!z�@<�Y��>�`�N�"�^8��94����ِ�c�9��PKgi��
�o�;cޗ�D���Dw��3�)]Aa1�i��[����Z)�RM�O]f�	���y0�8���D��I�y���	�&��2�sb!:�����,u<ǵ�u��x�Hz�W���h�m�z�Q����;�3N�8��E|�(�6�A���TF���s�`�b�l
�nr��SXu�_�Z��k���PLr&2��蹜�#�<!KD�n=�T]�Sڱ�&M���G�ث��Xo{��3<���E+���kiaJд�YX��B�eB��E��TE���
�F,Q��"֢�Qe��EAFEF�ciDQmb��EUS��6���c ֊��A-�Tm(�m,[F�b+%j���Ѫ�)TQ+X�jR�l�1�J%H�(�J�A���*�eJ[UQQFڈ*�-�e�DA+X�VT��-��(�5��������b�Q�EkAKmJ�X9j��2�bmV�UF-�Q��UQ1UR�"+YF��l�Q��lV�[b��*�Zc*aAT�Uƅ��W-���\��+U�
1b��[Vֶ�Z���b�ZVl[h��Y+�F1m�6֖��*Ŵ��YE-�F"��2�8ҥDE�[iAK���TZ��G�|�۽�sx���$����a,����W�遍}%��K>��y����� ��.h=��$n��,�Qru��0���_wl��a�y3gèL8|��x��W���JAc�s4O �Yf�)˱�i�9�"��F��7::��,���w
F)��Q����=���u�URF��7����g�rt-���g@L�P�S�
�F�/y�f��٪�O=�N\Xf"�,}��[�R��(U��ꇖ/���S�C:ZrA��X��U����FN]���~���lM>��M�E���&��,�HH�����t�낆q�<~Sni�//�5��8s00����1������\��`U�gb#���W�����:׋f��ɌK�8T�^i�0�#����i-��*��]u�.%�����X�r�a�16���X�\��9�B����C���#�5ݘf�����(k�2��/7S���;���������.:U0��o�ݎx�Ἃt��va�ǂ���$"ޥL�����b�_b[~q��(����]��U1�\���+��Vz�֭�=���=���������*�*ʖ�
�[Q��Vo(:��;����������"1��y|�c&4��,ֲ�1���mq�_!ҹ�l�ܙ�{>�D��ӳ�Q[�� ~V��Rwg$��S5b|&��δXt�l+B���=4	�<=�x���",�����$����cg��D�95�sʱ�,�j�E�46�zTu�V�ʌ멘��Ĺ����7Ļ��Ď��]�T;i�����17�åx��9�98�S��כ�痽�n�0>�N
�o]�<���|'Q�/��%%̹
���g<�)X����O�ow�� ���(�.Z��d��H��w����x�T�7�M�R�f�k5t��b�N�os1�5�9�:U�w�����=�jX:Z"�����`ʊ�/&�	�����L�J3Ǔ������r���f�P�!K�Qp0Tbt��yHvy�`�P�tH���	����F��+�U3����n-kd�q4<Ռ��ͻ�|t��X�����%pD�R���[\)4,��1%+6����f��֖�%c!:p��J�����kOW�19V ���ʱ��Љg+�$��R��	�l�}3٧b�J�r��Z`�u܆	����w�s4�疕��%]��IgME��z���a���g��4<l��T=��M�Ha�QL�F.�\-yj��v�/�9�@���Q���<����+�̚��x��0�מ��]�/NN��7Ƕ���Lm�x�X���ʗ�ӧ�ߎd۰	�)��N��>�ػ@.u�gB=P�͊�ՎB�k�BU9��b�Pw7���Z���W#t.RB���<L�p���u������4���dKDB��뎞�ǳ�AЬoU��k��"j2�܇�C�T��s�9Ġ���:	9(���ڍt;�vVq[vf��5���`�Eɉ.v���qZtw+�7��|���d=�/r��!z�����n��k�iypK��((ElІ����n�OT��:{T���
�s���:�i���{}��q��n*�r�0$"v\�W,u�g��I�ZP{Ҧ��1���g�Fw�҃������F[�}JMB9u�:e�����V*S=y�~�`�Iy�wa�Lx�~WY�7dYq��;�U�2p����8��]��T���;'���A��d�̶����o��J��}3n��TِĎ��aqINlPb�a�rC[N65�Q�il����8JA�;b�⽎��?���3�LIہl�CM�dh}s"��u�.����p���5dA�Q��t,ٚ16���v��k�DTo8��N�6��=���3C�D�p�=wZ����S��{Z��J��p�WefKp
�����7����Bʽ�-��b%�A8-����t]#��;Z�b��&��T#����>��% ��єIl���/v[�o(�
�Z���R!î��?���ۖWL��:�]{�����r���n�F'�h�tj�i�+�q�s����'&�p�P��
�����eV�$��hq��i�nw��<��~ܝ����|P�3ꦍE����-�ж�sS"���x�*�����^݌Jaa��WG]�{�w�4�cW��KmR���^пp���޽��k|r���*��3��L1g�E��o�i[�yLwc��"��V��r��ucz�~���<Bay%��G���PO��)��'׶�bc����r2�gd;�ֹ�Q��aŕT�g�TC���*�hq�X�QX���98�xP����&������ֱ�j�Ƹ}vx�HQ��P�HA��٘*���;��/��f��C�!V�E��#^ƣ��9��g��^>~ۺ>HИt��έ��8�y�Z*��a��㕥`��qN�jx��]��pM�K�K�8�b��`{�CR�O���[/������jA��kh��}�N`,S�gd)���˳��'L��T̀"c���.�&��pd��'���5K���=�����h����f⥴6�uMgiif� 	�����ҍ��A�t'&�j��������U��̇�^e>� ����h�m�Q9Y��U�:\'m�p^�;oSpho���1�jt��$W�uz�Ax�H�h�\i�lgR��W�#�f;�\q8��6���
đY"�V[�ypW���]gl鐍������_�?.]V��`IX�������9�\7Dh��饛L%���빠."7ڀ���kG�T�,J�~>�����±�b�ns��/�~&�����E��.9e���p��H$��Ș���:2��߆��zP��z�4����F� � C����>���rl��i�.}8erZ!�k/dwu]l�E���b��`�<�`��MY�t�s���Y���P�H�9��Ʀ��$518��ޞ�8:��1�,_�O']k����/���^�Ӎ�p�u�L�D;euvbK&����׭���tÁ]��7�U��Jwhdt������6�=�yK2E��W�u*_��q��ԭn
�6�,��MEt�Gd��7e�e�~	���I:U�']�%OϺ(6��e��U�p��~�48���S�VZ$lB�0���G|���Oq�ȱժ��`گ��V�xM�m��`C�n�r���]K=J!�y��m�YG	')`莫V
Z��+�I܉��);|���cŪo
C)��/K��^�չ#����Qe�ι��ؐo �s4k.�]�O\�x@�t��9'r{��YO�c�:�Lr�� l�;�tvԺ(\D�Ag���X{�������֍���:!מm�j�,ѰH�k�#���#A�0h�z�P��/o#�Z=u�Y�g���^�T�7�����7�2�C�O�[�,:0��
��H�f��]vg�o9�Z�����Ɖ�p���^��}*�հ�Cf&�5*�^Z�,_��S��0@��]nEn���H0�#��K¹+�/����LX���w념�Thl���u��ﶖ�Y��t\&�,�z2K��#C>Z)4�c��cagf���f9���+μkU���\����@��IN��YD�geΌ��
L�<�{������{��uŝ���:�8���+�ĠG�ۖ�������Y=������Ema��2̝w������r�[��k� ��M_���5DD����~�Q�U����\�F3�m,ə�$�vS�^��P����͢�`���p�)f0`؇ӢG.{�Ø��9�R��5!&�Y��X��Ô-{3_�d��0��ez���)q5h�S� �Ux&m#�>�U�L����9-��Ź3��1�쨿eY��I��an��T�A�\���AÔ6���=�U�2�ntE��SIE;�v����/���_U9x9����8+����
���3�����Ӫ8=���{M]��%�>����b��jx�D�����Mt�E��`
���W<��Ԇ�4Û��i�c��z�!9M^�_��f� ��P�v� �zV&5܄i��|��Y��b۱�V�w��p]�x���˼�ǎ�	��`L��F c�(.i��t���K550��%p��u��41pS�C\�+��+.�Q�=���f˃Cwm�'�3��"������8��YS�R)��윈n%~�B�Lwnw8O:�;a����V/#�qf�Ae��
�un'��1�X~y��:>���6�uZ�4�>�����%J3KwH�J+	qqe����ަ�y���i��G�歱Y�G�o2hv�7�1�4ǟ&t�]=����S1..�&1u�xި{]T���Ǜ���6ҬS�l��XT\��)��O�&�VpZK\�yϛ�ֵ�Y�kk=췍U������t��'�яΨ_P�}p3��� b�Kv�f�^�p��:Vg1�lK'C��۹��Q
�ٗd)��7̟�>1	�;/�ư��Ч��u��k3g��l1V�*L�n�Z�H���ہ'�Nަ%���J+C�fv_G�/)l�w  b�JH�
l0�2�'��buu�qL&Ł�n+��u��!����GrVv�q�8��e��}�O�f��l�P���H���/ȋ0�24��/�R�n�6��rcof��[Z5m�n��ly�aI���Xa�����#WK�Q�s.-������c�Z۠|6�&j�ߟ���XϨNՂ�k��NQ*�^n���4��֑[�l�p�u�{������8ӥ�ǭ�Sf��Cd\V��24C�J�ʊ��e���j�H�|�0b���i��x߃Νgd��}3�Y���E����[�8W�Y][��E���W)݌����z���y1���`�|j��I�1EL
M���{�7oհ�ҭ7�T�鳲�ۢx#~�2��6:���<�S����C2\Lhث�|�7��n�Y[�z�b��FJ�)4�=�xٜ��N������y� 6��{S�+g)uS�z��;�.J5�̒x=��S)���1l�QOs�"rְ}�s�K�sJ�t��I�i$o��ʏ��-�+2�fR,�g� Bn�yi#�ݪ(zizKmp�ipf�g5���M����л�8�x��d�,��wk���ʅ��8Է���!Y�@�_��!�ň��z������
N��
�ٱ����щ7�lܔE���f:�WJ��X�j#v�WXF7��u��V��m�nw�0�ֹ�f�����V�JT�y�\<��PV���E���r<��k���ޯl�^s����i_�t��3b{@��p�H휊��k7�&�� ��`��o+6N҃�u��Sw��.��e��t�.�6�Ls�����l�n\�{�R�W-62\UC�Q�K�rt�s��5\����|�����u²}����o�����E����J�O��Qܭ��|�g�w�xS�y��*��q�:��jy5�~�o�u��F���GJ�0�p�n5��L�,O�,�S�Y���<68��#�E�nt�N���,i)�[˺
ɲ�:@�>*}WsC�v�����v���H�_���j���풻������^���݋�K0����W1V�Ŕtkx	�ğn`y���V�py��Q��"��F���G4x�x+ƻmv�gg4���έ��;"��)�P��@�u�o�
�[��fU������n����(�P��'���9#'�5t쮔k����˛�|� �^�_mp���p��8���r�I��b�縷yv�m�2&e>@��&Xɜ�3p�R#O9\Lp�k�\�}S#Ou%}�ܚ�}X�E&�����b��u��;83�2��,E�+���զ�3(�@�em�d�c�}�&�qq2Ɠ^�]0�W�%T�3�)ݡ�<�ia8u�i˚�*A��N�/u���=\��'ݨ��,��ty�0WK TvI	~[,S/�:�boyL�o�v%c��&����
�q��+	Y7fR��ʤV�G�\��`U�i�ʋU*���.�|��#���!�=»]>�'U�ĒtK|�R�/.��!�O�2w���6�wd��n،�]D:��|(*|�$k^Qq����G@[+G���7�����{��ES�]E�/
.XI����fX�x�ἷHXta�v$;%�K�F1o�]�쒫ȓ�>�
ޔ'�m���qļ�ECs��ԫ=y�����ix{�W=Z��[����O�4�UB+"��lP���<Y�u9~��P��]V�9O>K�`3���+�]¤���O�FIu�Dht|�Rt�X�}�E�������铠���1d�	���-:�Й�f0C�l^���s2P0��˩�zA:��x6�0�:��-P�1���ř��Ey.��qX��E��G�#�����R�A�Џu�ѯF��m�!���KC�+Y��3��ݨ��E���X���6�z�3U=�&��˥/U����E6�0��X���:�yx�}l�r^�L�(��4�́�:�-�9v%���ATǼ��T�k�|�M�R�шm��A���ge;�mmj,�NVH�{�Xo����dR�7�%g�����]Х�b&������]�����1Y�����S�RkA��bRcn���w#_0�_�d���z�u;�>T=��`�c�.�S��e��2�p@t�^x�Loh���*�����	�HfC}O��N������z��ĦM+8������S���ka��
����h��;����h�����um��$�#2�ۑ�RoL�*]�j%�L9��j���̼$>�Ĺ�}*�vm �4��5��خL��X�ĺMmb���k�N�ۭ|֊9���Z�2�
��>�wV��_�q黆v���h�E��r6J��π�`��{��i�<�ٚ'��.�)�nbF�ۮ�XG%9.y�_"T{X'U���B��rl�v�k8�V}�N�]񨞽;���D��]7�>q f�i�K��M�h+�=�8��5�P�����d��E괿�-0�Amd���cH�)C�V���v;�_<��W�h\�������^�\)�s���iu�45�{�j���B^��e�в	tk�}:����+K�z�稚T��omb<�[l>����3���}WP�f(d3/�S�{3�}�;Sc��B�{�$l�=m��Ԟ[f���L�1�XD��<�眃:Q9��}ii�����f�^و�E^,I��x�����Cg|�������N_����x��7i��������ǩ����DtS�sM�����W"�-[צ�k�i��6���� ��mc�HS��ܜ��͜���D���ʆ�3�t*~�A�yu:�+�Kdq<jU9M�JO�Q�c].w\���q�n�Q/#F�P3ɂ�۠�1��0�T�Nӷ�1NVEM�ܩN�Vƀ�
6�<�#�;�N��?q����&�bsӵ<r�h���;�yђ+1�RTV=,��ɯbP��i�h9��_���f���YJ�`�/p/��������*�.��g!z\�:����:e,u�W�m~�(\;;�u���I�w,���L�<�ʞ������Z�d�����}�ӹ� ��]���%��n��L4 ��%Y��X�쫏�x�U���
T޺7B�.��g�����~˚]�An�j48g-}y䒤��S괡R�k^��j������C�`%{��虽r���h�й�.��]��`�[٪6�������]fI��)F�ERZڭR�kldh�b�0�	R��U�j[J�DT-���ХTm+�\pjZ��R�b[F�J(��-�jZ�V������D[�1qT���"�+-����R�Q��4e��Z�-)*���ch�JZ-�X��ҭ��ʋUJ�(�l���*.R�[q3-�#���(�+��-cJ�k,Q)���`��KkEX�R�J���kch�nR`�i�0b5�P1m
��Kc�*�������[+j�Vڍ���%J�Ҕ��Q�cq̭���+4(�n)J��V�Kl��--����e�+V�m-��h��R���R��e)E��c�`�5im-�E[Z��cFZڭKe��J�(7-k�}��ko�`Rg��k���hB�7GLʹn֑��v��!�WVE�(��2&�}�N�K8������[�e�}�Ek؟2��{���q�p.�#`T78��{:�'èt8��dK�/�r.2�V�WXmBY�ݎ��֤G��;�Q�H�p�I��R>���x0<��Fŵ)���t.'��S4g��[p�5���膌N�F���0�oS�Ebj�ò��r"���%1�EB�wn���Rm�?MƖ�;  ��0�j��(�vTc7�"�`���p�)�1�A�+sjrs:�sȍ��{�f�5�B�Z��*�/���{2�X�
:r�
\��3�XD��v��}��ۧpv�4���������������lc9T�`.��'��"U� :f�.^o�c��몪{�#�v8o;�^�ei�x�d+���H�/=*���O�it[`e459o��I���;�}�hEAO�-��Dk��rn��(Ɲ
�?��W�5����ܝ�7{��+ pk���
�����Ŕ��ȍq/T�=�A�!�<'�b�k2뙮���4�����#_�����U��@�,=�}d1^x�ED71���n%q�,�5z�r�j��1��_^u,��߆��7�U���֮:��weQ��ͪ��Wɕۆ�XJ)�;<��<��ި���Ş��}FQ�-�կh�W5ƥM.���s��z8P����������,]jݴ����䤩X4�뤄4�}��"��"�����z�nL6
��f{��
][��6�V�[\o׽��櫯��:Vq㥯f{��T��g���@��QXK��>��lЖg�?�*��z�:���a����yۯJ�H�vOY��u	��'$"o��f`\]�eu�x�V�8����,�����>��_�<u�~\z��1��*+�]b�	�J<mS��lE��S�����Wv(4`:��$>Sa����'
��v�u�p)�ر�i�(J�ܽ�|�o�cmzq�y�����b��g�n��޶̋�h(��V�jH�hHb�Ub�sq���r.�ƖM?ri�5��gÜ���u���*�D�Q	;p/��CM(̕�+%�"��Z�va��*DH�
��,��m�
�=�6���5�X�Okws����s�x{eE��^�g-ξ5N4�+�\zLO�U������[kn;����i��HT���/��v�nw�;�����X���-��
w��y�K�1m,�h��o�K'�����8v�5���T0��	�h׭�F7PҤ"z�OkQ�J�Q�Bf-]���ޙqAܧ�R8���1���ν�S�2�4�A�C�P�Nї�/3NS��D��*v:���u��U�F瀃�i���gn������n�ޮCj�@�+����*�o��-0�o������5�J����[�e�V���=r�7��o�@H�GVu�8���A�J��<�,_��ZV��;��Rˬ_�w���mَ�D�N.ӷ��>�A��_C�hܤ�Om/�g:�gJ�'׹6��W7}4*VZ�_h����G�'��ϒZ=)�+_�v���^
�Q叮�܋�]��7ݎ��3m6��v�N�l{L��.�`��|�A�Z�
�3f+�*���^'o�e� ���^<N���Y~��w��GY��43�:NPgV�O�R��Qp�i�2�D���W����,������3��s���v��t��7F:�'�NmnE���д�����)m�ř�:;�������e��������.�/���ۏ3M�= ������*RҸR�����V=CyԵXo��̳��i^N&�E�����TMn
ak�������<z�!���<3�!Yq��_�Ysw��	)#b�P;�RM��9m�Z���Wti{�s�%}c�%췗���4�^M��]H�[�G��� 9{�(w��uד�;�������o�y#{Kh�h�W��ޛJ�.�e.�-=���\b���SȮ���a�B��]�)���bU�P��c�0<�9D2��w4�"��d�ӺFuڈ�X���=l�M@Sp�n5��D���^�Y��3#h���|}i�<}�Ҋ��T8��&�:k��]и�Fϥj���"c���taj�@Y쁻�������nEb0���T�� �U=��5<)���_�Q�Ũ9���
��]�p$m�r5o�λt�.J�d}�c�����-��ah�����3	tT�t�-�;���@���..��\ �����x;�^>r�����xB��ñ����;�tV�C�O9�ƽ)�%��%�	sԩ|�WPm�<���N���KLfG9���y���ރ�Z�E`�[S����^�d�8%�<E�k��+ݒB@�-��(�k��Žs������Or�G�g���z�b�xR�J�D�7d�CH:=�ι��$8�S�Թ��#9�mW����/CR��9C �
�u��M�ʈ���[�2�ii2:e�hx�N;�ӱZx�s/�0�K����Cw����V�f��6���وf�x6�]�x��T7�A	lf�"R[�8�5b�����=fWYR�e�f7����׃���B�r	n��|q�׺X於�ۨ�g�:L�tDO{���mtZ���x��7R���b��,�L�>o�Y-3�gs���<t��y��3X�%������G��T�7�.�X�p�7�2�C�O�[�,:0�3��{vY�y���6�j{�Hܤ�$C�(q�zh<��-u/��Vȿ��_��Y��8��\�ޑ�oUՂÝ�| �-�:K�.���p�<&p�c�qV;��9���O5�Yst�Nbmi��'U���g��/� �-%a���|�R%�,k��qAZ�nFc��m�u��-	�������r��K��yಉ,(
�˞WT�Ne$-���Z��vo��jUe�g2F�$1(��ĠD�n桯,���ռ�����fB�\\��&��mX~�w�U��W�v}��J�Prs�`�MK �h���,�N;dj}��Y���%d܌�'��ɫf+�{U\f!�F���g�Պ]�ه�4:�{"%�+��e����N��R�m⽿"�ܙgf�cYr��ˁ��D(����o˝�me�k*����Ř�W�I~���qۛl�����P�u�*��J-+Fu�L����Rf�B�`�TVu)���U��@0��DN�<��#�A�D�c{�g��6'��R,N2_9��^��44����R� JU���wHf��v,I�=��>�(�s��-���m[����|��z�w�\��6�*���9aoX�^���N�j-^-�v����^��g�v��i��Ӟx�g�����6H�/bUp6T4��f&����e9os��@�K��b}P�)of5�z�(!���0���c�����EM*�^�m�#��w0�e�U(T[�MB�,3ol�M�p`'Ԃ��Ns�a��CX��H���V<��3/��+M�	B�F�w.�R�1h��������A��/��PRn�rv�\�l��<IR�#Cj�!~.J"�(Y���	���g�:�j���}�����P��Dpծ�F�����N#�óq�1~�t`RrQ ��ߦ
>�
�k��PY��޵9���ט�]fh��ڜ�%يNz�w��	�%��c]� ������^R�R�cp�KOj��ׄ�^��� ���Ӗ"����m�b��D�K�
�`��N�m���q�O�x�*,�ʝ�$4h1͙�td'\E��Q.�CU�Q'9�U�m>T���j��$gip�깏�U�)):Q/6{�:�D'���:FW���:��������2�K�7�V��.��l�{�]�a6k��o�@(h��K&
���Ø�����6i��w)IN_#�.�|d�ч��Z�G�ږ�b�WA�s���2t'[]wP�;��AL2�_3����L�4�����q����t3�w�؂��Uji�<6� ����r4��n��MG��T�8pn�N2�ҁ�m�J�H��Y;���1Lv}�Cl�WN.g��XϨO�k��h����_�La���z���;2q�p�P�8��1��{T��R�����e�[1<`7I��]Z������u�_*�x��b�;�;�#
�pn��.9����P�*W �N�*��@�Vwn5�$�v�4�!V��T/a���-ꦺu���O.4mi�ÓN䶸\nމ��8��uٜ�e�zcI�.uS�q�%oӡR��c ��ڗ���c�3a�*[���=;Y�S�跘�4Pd1\(P;$��QOZ<xθ��i�'�˱{�[u�g4����bg�`�%ؙB�����dGT�K��ʿg,��jϜ�in'�V���=�䭫��jE���=�ln��#�4�_$�=R��*������F��yGz�u#z�d��0��{�j�[��JS��$;�f m��Ԧ{(To�A�}��Sp��b�`��;�{o�B[����V�9�LCF3�.B�ų]���	�)B�Q�P��v�ɰӼ�3/�(��m銺5	tyѕ�su�:���`y�vh{'Ҳh����k���:�»����ι9-��S�>֞����y�G�"�l�X{UW~s���}�t��2�y�~t(R�x-'��dr]���r���~Ũ(_}��q�1��k��nMގ�F]��Ʃ���v��46���6��\��H�G�K�v#W�5��JZ�7�4䪾A�U5N
�Q�ʲ;:6�ou�u�a�\�`����xVB��j3�]̕�׎�3=(��b^nK�Ff��L�orù���g��#�wRŕ�Iw�X�6�g�x:��U�z������VWx�Us��i����EA�J�@�NB:M��:i���q֍�O��]R���I����h�U5Yk�^��Vx7�\cQ�w���5���X��<i�u�Z�8X�PsL��n���r���%�37��C�^�*���٠��[X�@����/Tn��膱dP̛��T���w�XQ�O��R.u��u�J��}B
��T�������	�My�#z(�ؓn(�˓ܻ��w1,�0�U���[�t|([Bg"���q_��d�Jgx�F��:��;U1���ī�r!3+��	�·�J�~Uꚋ��fQ3��ۋ��7�Il�1�üq���	��bi=ȕ0.G4^�WG{��!OѯOH�رs0�wnMZ��\.�C�Ȏ��ٚ�urt��[�Ĕ�H�}�j�t^��g����\�b�� ��u�N*$�J&kZ����z�o1½�m�2G����R�[��p~�2%�E(���]���a��~�a[�p�~�;^�u���{�ݰ�M��:�[���w9UGN�-Ğt>a���{��n��v:�m��^��O\�_'u
��挌���S�t�Q�.���t�U���^բ�"�y��x�*j�v�.Gx7dPL�C�l�����~��&�k��=�WW6m��&묾��jX�;���&k�T��<-�Pݝ�4���h��4����n��������oh��
@������v(�o������==y��-?F�y+j�QP�-��އ2�+�u�/ >���R�:CǏ��8T��3:�u����n�'�2[�v&�!Iu���`�n8l�g��Eׅ���76��w�����y�UY�,��y�l2��YGt|3��1ilp�u��4ɖ��O)N�}vWmK0��˦!��@��^]��+B�f�yO�n���D���3�fb�n%���׉�!�G��N�'s����}q.J��^c���Ŧ��������U��W��9�d�vw+����l5xeed�q�*+ݸ��^�h)��(����mSZd��8�T�����Q�yTV:�U�Fz�NZ��Rk"KەU{���q�1m=Υ���o���c�Vr���m	�[�9��'��W���A�^�uk��|���~�W��곞_gK}����L�ˮ�E&����� ���U�rYq���v�mU�P8D����K�M334?N���a��ގ��G`HW�)>w>W�p�5�P ���"sr��nZԗ���:�=�p�v&�!�r�j|�����ݳ2_D�ֶ�QT�u�X�u:$v��U�v<�ԝ�o�>�4��\smMD0S�I���L�Q������tn~��{�<��=����$��H@��H@����$�$�	'��$ I?�	!I�$�	'��	!H�$ I?���$��	!I��IN@�$���$�@�$����$�$�	'��$ I?�	!I� IO���$���$���
�2�̃�ΰ"V�����9�>�&��OPR�_cm��l�J�TU*��)U�54�&�٥
�$Y5JJ���!J4�
�V�ѡT��il֚ThҖ�kM��Œ���4de�m��'
����%:Ժ�+j��F�T�l���i[Y�,�J��Lm����B���1�d�����4�l��j�5jګf+`���6K
TK1��bj�	��V��L�UR��[Uf�Y[3[F�(��ڦ���5�j![2F�mfԛ��B٭���� r��kJ����%!�rS�֥��U��U����W���0��wn�����"�]���4ЕU�sN���N�)R(9]�ZbR٥,��H�Z�x g{m@R��n9mU*hk4뺠+jj���lP�VwJ�J�.�n���,`5J��ֻmV��S��mYmYj���H<4<vԲ)��a�Y��l�kd�  �p�C��� #�8:(P�  �[�B�(P�B�[�(hhP���uz{���С�hEz��CCC@ н����@=�����(B��w@��ҷj� u@�6�Z�h6ʤ64��  �ޭ���'GZhj:�+]:�i�gU�Z;+�֚Ҭ�� �4��8Y�����i��6��u)l�����*�igET�-��Jɥ5hh�   ܼ�)��euδP�uN��j��T�mݶ��Q�BS�- �wv��v2�Ύ���kWjwlh	U,��jR��lj�tS��6fLE-�  -׀:U;bn[����n��+��m��w@�U�0��R�A�UՊm]n[�����:��h��X��B@7)��(J�n�@�`�TMa-��  0�� h{Ur��MQF�b�V�V�ڠ�@L���.qw!N����������9�*����E�[��wu�[E5��-b��Y����  mz��0(�l+�4� �n t�l�4�u�([�sP(�p� u�� :��E��ղ��LV��o  7<��(:�.����P���݃@)X ���
�� ��C��A[� �u�TL������kjԇ� 	� �K� � � 4�8)RU6� ��N��L �pB��wp6Ԡ&n��Ц�� �<�3*��L@��)�4Ĕ�@  O�T�j 2 �~%*$  &(�L� 
I�ƪ�� ��ЮDd�D�(�IL��̬�VCQG����خ!�^-�br؉�C���}���>���?�ED�T@QO�Q�ED�b* �* (��zz|���&�Y���^�2<�f^�84�n^�Qp�$�Vi
���f���F�������^�b����+��7�\j�pi�t-Ƌ�*����*r����!i�f<c�B�\]Y#/dvE-ݽ�Tޡ-@qQQ��[61K4%��6u��Vl�R��&�)m����,��QʉG��vj��375ŧ((tH���[/E��M�468ɿ�!��W
�i�w��^۵��]� ���;u���73	��aV�^j�����m�b�B7&Pܬ��fI*�t�
�f�ՊܷP�J�D�Pf����5j	sN��ҁ��3r��kp�R�7A����O�ZYH�C1F����׬LZ���ة!��s�yX�2���̒�l�lC��q�R�JJjskǪ�[{�hy�ȥ�Pܼ�aD��Z����;H��v���T��	������e�k����SY�C�Bf�fi۫T�R�^�v1"��!L8�ʔ� �$F �������Yx,$ˏ�����s���z���@��Kx��P�BFBj	Q,v��^ڠƍLQ$�+��.�U�����N�߸&tB�=�=�c�eս��d)��CwqCe�^�SQ��Z�f��FZ{X�Ek1�*�Hj�$<Rdѭ4�#b�M��ج�V�`��0ظ�D"�Pf풴m���]؜����Rzi(sf,�6�$�/%-��:ݫ�>�B��^l��Z���4Q&��(Q��\V2m]VAwf7w��&�0�`F�f�Qk\������{�o��'�CW|������_;�atLT�Z))��
1�v	��l+���mn����i�CRý�+(k
��3,d�ڤni7�����q�;.�YCAƃ�x�Ż����_iR�-���6� �nX��>S;Skh+;�	0�=(t�t����U[�u����q`����k�5�j��X�C�`!���sjQ�rjŨ*�l:���S�S5�ħ_1��苣��{�6��5�\��0��_��K)��`�m�����b�hPIh#m۬����x3Y˃p�S\&��Ƭ����*U���0����6�o�#�&	xТI�鎁��-��c���Z�&yl97U!{���	3u�W����V���E�
��S��e��r���Ca�M��W��T�P���a*-�v\l��a��!Ei���ɽ!����<�p�t3�tB��Áf�����X�F��m�gZ�Ut�z���Jy&�NK��}X�&v����̷�Rܻ����g�t��;��kU�E�/+D��T(�`Y*�p���V�d���v�3q�$�VܚmIL<��s��W�^RT7�H�d��RL�j�*g ����4AL6D�XS�y��ׅ��*���+(����h�hp���� V��3���aY�J`p�I!i,7%���L�V���Zw��͢1����撕b�D�ܶe�̣bEM@��rr�x��f7�&��S��i�JL�R�K
@�ə�m�D'�*S�\t6�Z����q�:wsXN]��S��賗���1����e[����xu�y5lu3o�ϕհ���X�{�h�����f2��^T����<�a[��~ٱI�O ����9�u/hf�Q���գ��,^�O7(�.2��Ȗ*l�,�n�ڠ���#q���ˋ��+r�aU� ��$A�2�p��#pU�O��F�2��76w솎̎�Ҁv��e�l�p�*#�$��7�`��Գ,�ڷ�w�=��Ь!kqM�M�nD�;�6E5 ���e@��͍�JMz�Ylf&��@�h�Z���N�[�],�R�ap��,�&& ��HV��8yB�_A7*�FB�L�c$b�ܺ.�J����`HAX��4�c&���G*�EV���":��	�,�F�7$y0�-%��8��_��"�R�v4�V���P��Xi=�m�4�&]��q1`��j@f��cd��*�7]L�n�-�4���ҟZB�Ќ��Ǒ�z,6����c�a��^��.�4�RR���tj�R�Ay��V��Q�Q=��GL�ֺ�u�����[f�Q�AS�[���$zsT��0]k_��$��K$KSs���|�H	�"73+ZN��m���B�����S�L*���8д�z�ơF��5ݵL�<�
F@�ê��%���%Ǜ[Z.���fnN�/3������zڶ!�-�Gj�7�T<�ZT��cM:�z��p[�)S��1�0f�3N&K�
�X��#?H�8�� º�Y�B�hv��Uh5�Uv*a3k0�&{��|5�Aei�eKǓ�ǪB��e�#��ZS����Ŷ8��L{0B�l�2_�H��激�@6�y2b��V�U ��g5���#݌g�$F$��6Ž���x������vaȆ�|�r�]��3z!��H��e�Vwm'�ˠ�:~�BJυ2ޚ��̕��Uێ]�Njl�qn�0��֛5&��.Ĳ��Id+�ehu+�0�`H8��f��z��a3��n���ݪ��R��E�N�QzAC����7�M�M��`�]~��)���P��.��B^f3������F�d�ܠ�ҺG_�kb%�Q�.�l<ڼ�6b��VeV�{�MSq�[[�bj�PA���P������vs��̨�l$�����Qs��&S`�u���xl4ڹ�U���,1C
��ݺl�Hb�vl3fJј�T�NRh���Xm��գu��R���-hd`QӍ)���E��J�����uj�+7�N�ͧi���ZtuH%�����t��`���"I����٘�l^m,y��^�1I�Ԕ���7�lC	��kI%�Y��7W��*G�ִm�i���N%{�Ǆ)�f�
zsh!Bm'����d=��Mlkhӣ�(�k#�kF�c�,#������#w���;�MA��*.z�aC�)��b�\�;��In�af���ZVr��66�ݪ�PL�#F��oi�
:��b��S�+l��ʐX�ނ�X��% 3v+y�Lh������-��J�BmC�0�	G��6�밃y�@�J�M�
��޳6��ܫ�	��W"&�j 2AK`���Y��ۼ��i�šM���T���d�i0�*V9 �RD�jf/��L:��5*�:!"
�W�� ����������&-��X���+&^�(V���f�-���k�f���NS� �,���v���˦1e���3o]'�uR�%��0�ݤ�n�-�	�U��X�(��,P
�K��n��a8kEjG�����6���$1()�d\��9D�%µ֭����n��<�a[�f�xP[��V�Փ�D���H��RR�Qf`di�4�-fFoN*��	p��kr�&�l%�/n����8%�� �a���A�گ[�Yi�uܻ���KvP�#�30�wCZ�&*�%ջ�05f�խ����dU)|���1��|o.���/�%*a�p�BR�0�����52��^*q�����i��{&,���@/��Y�rc�$�����_%����Ғ���*����Asu���G+����ҩx�V"��ڬ�=R�|j���Q����nnjv����mC�h&aT.���)h.�ە*Kɒ��{�+�&�t7-��n��xC�C'M�mZX&�I�YM+�s+~��a��qV4�\�x�n MV�1`2%=��3,�KJ4]*A
b�LwbT��N�N��a���җ�&�@KJ�e�g6Ɖ@CMJ�V�;҉zV6��*�*^^��5��9�]�x ���eUݍxTu��=��B��R:�m�Y6�J�;�+/F�[h#w�j�qб�),L��N�O+(τKw6k��%#��qd� ����ܠ�����gkh�zt��%[�e�ba���Uhk�QZJ��b��hAX��]�V��BSp�I�C	1){v�7*ܲ�7����R���4��p+U�l`L��[u�&+)kb�7i⛄���H�k�v^J�u)�ӵ�R"�J2F�[�y��Ԟ�3n���kR�Kq-b{X$�&���&�/Y�m�N�����N-b-U"���9��r�p��1���s�k��
�'ܭ�A�{� ������p\f�@��؎��i�Z�8���bڨ�p]��x6�ɗUj�'k4dV�/-ˬ�o�c�ӣ4��f�X�ǖ���Q�Lʹ-�,�oE�[q�b�Z�Ѻ�VfT���K8�#��N����9U�����K5f[wX�w�fǑ1B�j���*�Br=@PU&�QƱ`{������O*Sǯr��[������z`�&�۫�mEȞj^(Jܨ�tb2�n���Y��p�sD�y�nӂ�^���Y�rCFM�~ٹ�(;U�(U�n��K�I���)�JQ�`1S[x��+(-In5�?MYI�X�,�*[�${OfY���0kd��H�G�gE�U�:Ѹ�D��S������.�┫i�:�0�f�(�˦�EC{N'�ud�`��X2�c8�ãKU�͊�FkE���~��!Lb��kL܈1������6�D9Z����$8�Z��W��ͷ��MV;�{�:���#�^� v�6�Q�q���,��է�����m�}"��w��+"�P�b��
b*�3䪱l�+Aa��)�%j�ٱR�!��V7�^V�XЏ	[ud�p(m^�V=X�Y�9�L�Ǚw#����S/�U��l��wMB��*�(5+wn�����*��ի q$Ŧd�)��:f9��%�<��,��g(,*���9�]8J��ۦJ{#�&��w!��i,����ɭ�ʵN^��I7J�'8���T0(I��Ճ�,�3mJ�v�sPr�Ie��{b�ʗzk�Lt�aXp�B��%&�(�Ϭ<�*Ui�W�hBi��T�xS�%R�8�T�=x� ڀ��6l�PX@���b�c0����Kb�6S6�
�H-YRk�àl����hQE��0��Df�� ����ç�Nѭܰ��R�T˿��;�uZ�kVX��CP�i��V¬w{Tt���LL��ŝ�k0Ɛ��oYY�j���jQ�	��%k�H�bv)��xgLg���f��\G#˱񲬫;Y��n�Y���-�a=�"�=���SeǑ�xz��=ں���l�n&ڐ
YP�Ȇ��:��7X���Î��<"�\.�n�B� �W�UǙb��
���x�%
Ʃ�W�镐Ps\�"�o^�����$�ۥx:Ӥ�w��R;Im�#D^����f���`�-me��l�Znh�.��h܃%B�j���%2k�u�1ѡ���Y��©�hԩ.]�;��4Ty��r�3���m����"YGfm�jD�v����o(#�رEl������G1�ǚ�l�J؁B�o6�ض��15�ص2F&�cw[�l�:�D�Yo1MǶ���^����f%�w�1y��0�1�I�[d7�F�7��T�� á�pj�����f%�1��]���6k(t�a8��vk��t�O�y4�x��T�2� kq��\C	U��&��E���Cb�����ܶ!&��݋�-�[�3eMV4D��2�wt�Yl"uUn(�P�uMJ�k�k�����u$�n��',o�m���U�(0��R�6at���� &ٕ��T�ņ"���k�{S22��l&I�E�����bՄ��*�0z��*���"�c�����V��n���ӄ*Gc��چ��e������tE�"��|]���)�ʱU��q���O�"�s}#�D^@����W��ۛʣGa�81�S��[��r�ʑ�c*�����Gn�"k��Tf o��k�����dPY[���ܔ�%�IZf�9��v��dK�ȐCR���^^ͨ�c�6&#5o���Z�]��#-�M<�Ѳ�uYh��V��%S)���y�0��0��,*g�C�Ѩ�ՈлyMk�Hz��sصm����7��,4¼sv�(f�%�IZ����G��C�Ng4�t��5�=��će�-�^��a'g뚕�j�
Sd���Yec{�t��"�����(��QYj�G2.�¦]�����b�ph)c$-�Q��٣h�(�4�F�i�Խ6sZ9�b�Ձ	��:m�J�DO ����*�5�,Zb��[Gu�Kf-Ѭ^���T�F�FX�ܲ�Z�zp�GK�;j��B�3y��^�УX�-�US&��Pg;��u���'u~1�C����~u?s5Z�r�r�[��2=�0�MH.��j�%t�̡�alZ��-���DsKf�Xpe=/r���{xɑM/4�Eփ�p���F0�.��5j��M+Ud�B(P,F�;�f���IZ��x��ϱ�v�a{J����`�R��:�O��^���9<$�:"YŮF�)l8ݷr^�)]3���0�Fm^��SR^mQՅ��pnkL]U81����A�VU��n�n"���Yх���:���r�ݔj��t�u=4���Q�ͅܖ[�+k.�6`:�Z��3� ��al��zy�}<!�YA-^��>O7�|t,����ư뺘�ʰn�4Ҧ�(�b��e��n�㲚e�1ܗ@k�sr����`���������n��9ω�8�P��5�k����|��1�0�hDk��5[Z������A�����WJ�7��a\����O�ui�X��л�C&*|Ȏ�ܛӖR�$s�vJ���O�qMeó��n\�� :8'�gc�U��	���0�|��p��Z(<%�w&y�}i��R��p���p���%'�� ��<���h�~��l����C��w�q��0i��H�U9>9���,�.�dSfaԎ,���N�qn������5hk�N�Aq)�p�p�b֦�W˧�E�m��x��n��@;Zк:��ʃN�NZ�N�R̚4.\GoTLR|��)�J)jXy�V�T��(��ou8/��r��Q��sp�8�Q���ᠫ)��Qbav�j��Ujƌ�o�뙻T	$����K?m=�F2�X�.`5����,ȽW��k�_m�s&*�E�����Dɗ�6�۳��;V�HLSE�[B��yŁ��Yr��Mb�%S�=0�{o�\�n������t�4�V��'��5u�;��kU�*�F�˺���ۡ��Hb؞�ʒ��iX�<��\N�%��O-� \���s��ڜ�Y�_�o����y��9��3}gL�w�_M�
Ĩ��ÛO���:��A���!p��y��Fn�R�Fb��x�Zz ��ᾲ.f����Z��ʖi�uҁ����!�L
��7v�hk4L7D��ii��ݎ��L�j��w�K�*������.��3�C+���y]�W��9뾥�xn.�C�X�T��h���\l�(�3��P��oY�k�T�NL�:�������`��;�3��|8:`���Ev�M���罒����k祄V���}7jq�X�B���&Xj�>GR��̔�m^��HK��_ML���*���$�e�k���:/v�η.��j�"����m ��gQO�<��X�{��#b�Q擛��"�Ch�l;�1<�Fl��v1��P���7n�j�yHH5y�)��/gA���1\57��l�4f�i����&h���fV�b�ܛ�+h$�e_-��F
&���0�+���\CA5h��l��k^ӫ�K`�����Dt1�؞Xdjl�*</Z����49�z�A�GOVc�Wq!	�����P��)�R2���Yܤ�ՠ������b��N�qcfM��bh�T��=�i�Z1��2���/��N=��+����E����u�5u�fo6_�]9x{3x$�����B�;zD�m��nu����\':���#k΀;'DwQR�řg;A�Jq��/�f�b��g0`yx^��SD�2\�*˴�;��kw&Z=��;�;,'XMbu j�u
�b�� �+� ���ᧂ�P�/�4����۹m@��9a�'H��)@����X�BC�xFf7�{o]>�K��ܰ�o�y`N�A��Q�+sb�r�R����P���5C]\p���oRt9��א�l�շV��W��o�ګ�ɴ�K�AKs�:/N�f��d����Z4d����Ń�7��r��+�,�o�(�K!#w���4.�o:#4	��U��g7��I-��84�+���[o%�$e���c�TX�t�pg�[e�N{]�G��=Y����S�P���5�*m��pab���˺����
�Z�����`������j��y��]���;P��o�☜��a�2�n�Po�l�MG�tch��:^
Z��+~�6�p�1�&Aj	ĥb�u;���6��01ڐ���}nzV辤��Z�J�§h���:���մQ����:�Бg{�exf����:s򒜻��_f��P�Q:Y�RD��7���v��s��h����+dmj�<��g�Rz�^o�]z�:�(2�)g����Q&��� W�ݞ�;V.��Y���(.P:�٭���^���>�og����z�k
��B��-Ya.��R�w>B�yte���[�m�>trX'^�nG��8��w�b�r�A�[ۜ=��ͱ���˳o3�f�ȝ�qBrQh�����p�e�'�L���^ �v="�����E�4I{n9�+���;O|7��8A�m�:�#}��f}�b����Tb��;��kS���c�=r�'��;Wn���ы��dQ�G�c_� ����<�P�\ �->�>��+��nΙ�oC���CM�{�[e�|%5
)�z�r��̎�a��G���M�"O��29g���h�I뗰���,wIVd�U��,�2�psvy��J���K��؛'5�}��s���3��u\m��>����~U��u����R������@���ݚ��t���}4������l��f�q���^��y��ۛ-��[i�-Su��$���Yp�l)�1�",��ڗFg�����{|��Cf$�)�c�3�3d|mM�9c��'G��Py�����fØ��n^���[��)
a6Bٔ��U�n?5Ƞ�|$Y���׷f��&a�x�а�l�|bʁq���\�l<zc�j��(~�ΰ�ա�r��r;��n٣���5ǯvu�
�`�O���Y�W�6�Ѡ�ϮcQ���f̲�9-�XpmКk�Ʃ�)��'��PukX!�[*���E��R����I�{\H^�-��Y�s�:ty"�=\ gw��[u�>���{/L
�z�Wn��S11�e"�@�L��6�c��`8kM�{�d#j&\���Cl���1E�����핣wM;]�Y����K2�q=^ٹ�D� ���1�]�A����b��+��᥂�A�J�.���qT�
�7�:`ی�z�rX�Y���_�-����]�e�-��ACw�E�Һu1a�c�y�u��9pS���C��<6d��H�qT����DFY�	Y3�GT�����T��aB��ԥ̭vB"��f���2f��7U��ͩ�]@1�/��}<��l�!�$˚�Mz�1��e�s���]���#Rv�>R�q�)���9��5Rb��.�Қ�sy�g�����W|,��Ӆ��{�5'�����<�{��d�rd{3 ���z�xgcO�ײޫU� (#s��&�c�ԅ����s��:W�/�v�G��`�5�$�.zǺ]�Oj�ԁ�0/-���d����Е���^��G@o�r%��<H5�U9ʕ���.�N��;6IҶuT���f����c������Y���s�J`��'kBd�w
W��ʉt�c-�N�,X�H�.����ְ�jX߄fW�M�k�`�{[X�AKa�Όt!���Z	*@3O,c��Y9�vk �ˊ^Cx	sT���:��&�c33ѭ���%J��UУ�dEu֍q��v���'TY��[�+��y{0x��'�1Z=8[�\�e=xO>�M�hsY�9��i|��x��ű�9��sܓ3�J�s�þ��\ 3��-��.�箦M5v�ͭz����x*��NdX�ג�����I���y��$�`�#�Ou���D�)���̵S �T�p���i�:���oټ�SÆdb=dN�v���,^oU���W^]�<K�^&�M�ytKѫ�y�c�Y��f���.����tM-72��UC�����2��
r����R�P�_�J�IoT���`Ձ���*�@�2BI�
ì]�R޻�CY\�6�ܮ��$�m/���30/�����ˆ�������������i�.j�"��8lG��"J�9��V])!�]�nZ\D	݇���W�M�����	&�W�>�lv���grf�B����������U�y�2�����`D����ɛx�٨`�V�t��ǎ��M}�q-R�!��ryq��y�5�a$wN�*���xXp�{{�u)�m�R���"��1* ������R��RD�ޜ�rӭ���{uUrA	)�sZS}�=ˡ2�r�:��w�R/0;仂��m5���M���4D�>ȑ͊}�����]^�Z�:v�>"�zʡ�^�t*�z��&��t�H^2��=��޺�3�����.-������B�qa��o��kW�;�X�=W24��`���#�o*8��^�f�^�=*C4v�OŔ)�/l�<�D>b�ZݚƙGqU�����4F�S�y[�n[~ں\�?atc=7�fbtz����.6}��������
��a}���2������o(,F�1�|�^�F�9� �+cOs��7"M��+j��Nqo[���`��,K��:v�)�s��<�v��9WOS݇F��'/RE��ϵ���Kk1�htT�Զ�0oi�b^ܖ��,�l���
�eƵ�Wu'\��j���[X�a�l�Celp:�Y��z�>��6���C��5���poV*�o9�/F�I���_G�p�g��L�=��	�xD�f�ݹ{�t�ԅ�[{tc�^v$뀅iV��f��X7(��ꭨn�A��ײ�r�ۚ��˜/;�n����$s�Y�::�c��b�+u�{n��08�����L!	���>�ף���{�-`"[樳�BԮ���gb��\I���/��F)�[���F]��;��ٵ>S�j�?5U.`�Ci�yM
��.��y˞S�Y�.h f	S%[�u7�����)�綉����=��$~L��C���ٛ5��8U"�mf%��������94�f$��/o��D���3w�c�F[��M�֡�es]4�vk4vH�>|�3f�g6��g�[�4w�.So�u�}�.�X�k&�.L�4����*}�*�'WJ�۔ĝ`��A�c����Q����Wx��-_�gs�^1jniG3h|���~꒜�n����&k��.���v7����_���/bǹ���ٚ ���=e�x���t�\��������\M'��O��ؖ6A� -YF�ǎ�73܌�6�}��::��:t�)X5D��$�q�ϸ&h�b[I���R�*S�v���YÆh���O-��+�ޚ�2�S�C����gp�8j����U)�ր��綏q%Zz�	K�}��^�n�+P+��=׹���f,�>#���-����f�3�[�إkq���6rɮ�#�X�i��w\ͱK�n|�=�
�����'�r���U)��c\�RT��:�T*���D����NLM��p��{{g�s�|Q�;�-�b�[��г@��(/$�������go�)v�;�E�>W��%��лN:�Šo��8�<�{*[�>�N�"*N�t}���r�m���}�Wq�k��9�$�SS ��A�d᷎�3rx��*�ZW��?L����f���/I�����MM92���:�;V�b����uejwK;��Ҙ��Y���q�����0�י���Tx3k��y�C��q��w�G��c<�E��n�3�l������8h\�<A��y���m�b���ssʥ�g:1f�ʦ�0���x�!�{C�ެMr�GL#U�Y,wfw1�	�8m����b����e�(sg���f� 7h+z��\VZ�x�[}LN���}&�lI�)����U�k-�i��ܧe�Hl�;�wZ��2�1]�xwX��S�]Z0$���E��C �E̫d=��E���KtzRh�pe�#���"3�c�5�v�H��`����]�c�-�՞ᛆ[���r�Է�>fVą�6V��|{��ssGùe �>�yJ��{G�̛Mᷚ�E�b�x�b�͖:A��r����ٛү9�%��X��l!��#ɬ���r���2A�uݘ['͉� ��v��gGz$��	3a�ﻨZ�9ʑF�rL}����&�/���=}�t|YYV�/�v�v0�Q��޷bW��ۡ�ll�-�V7�sn:v��� �%��e]�j̾�K�bZ�7�vMm)0��{��� ���5�];U�wD�fb�ԥ�F�Ӈ^7�ZQ�R�˾�F�DE�&6>�l4
����Y�3ﰑ}�Ne`���k���<��i��l�G�k����R�c^c��k�$<xV,[X<���6�h�<=��mA����o�����zs��B�Lmn
�A�:��Lٛ��nQO*Dk�S��}CI0�M�QӲ+�{}�x�Hw�l>Ի�oQL~�Og�t�F�}�������N@�F����rTWݱ+�WTs{i���`�]�E�Bj�2�v�Y�3���&yObg�򖅹�)ӧ�a��z�J��' +E�H�e���`����(^�֗�����z��Mb��Kyd<�xW*��Xi�x.��)��J5����֔A��k�Q��{9�Ǒ�����ωA�\7�� �s/��޹1���fdNQ�#D��s�ٜ9O:�c2�=�#�9霽�� �==�3�8;�4��|��ε������O��3��o@�MG!�.ڗ�˘��tr���o��V��&wW�����d"U�e���2��-�B��S�~sܵk'u���F�ú:�E�f��{B��I�\�� �ʩ|�U��v*U]������]}`n�"�8�;݂c�o���tg�Z����6�!���4u���^���_NٌQ��vb����o�����)�n]�%��	�\�M��	��gn�a����̚��o0Xق�/Ϸj���x�͎��	xR园^>�(G��elU�ԧrHnl���񾢓c���;�Ҧ����a�����ͳ�΅z��p�u�%v��v��4L�7vm�1�{QD{BZ�X��*��.�X��Ds��}6�[�7W�����|l{r�n�4.�w�p��
{�k&E!�ڇh�cݺ���xmy}j�_o`��k�iC8�]�����_}�}U_}_}_����������T��DxB鵄���U&�I�F�Cm��t_�u��U�"(k�C�X�)t�vTT�E�VZg�:��`�/��5�����|1v혅ϭ'��FG�Q�v�}�-�k�+�����k�7�ݾÙ���?p3�GL��w�t�X�K+�%v�6'm's��S���DVd�n���B�k9���%�	-��^-�����u��^M�\���Q�/����~S��N�^@���n��}���S���%���#|F
X��Ud�$}8�4>X�P�2#�'D��9̤� M_w������^s6�]�ǻVp^��%޵%�������W��6��f��jQXLP����wnQ��E���j��%߁��yRa��&.��-����Ccz�+EN��_{�e�p�8d;�]���rz�:���z���6=��IW��黵�<������5+�*JP~+u�C�}��l39��Q��=�y��w|N���+c]y�:;�r�����^��G̥YH�QL�����*(�aw�g�F���1PV�^cLq������kjE���ą
WS�l;��k�j�	(�@�H|o�z��5�����mm�;V:Ki��s�mȜP|'R9[v0���p�vi��S����5���|�E���zI��� -�~�=���D��Q��^��AL�6�Bs��<C%���#�yp��YbS���of�"w=	�l���C�qs�b��3Y7v+�O:�ƨ�+�8�}�E��Ekq����$�����<�n�L"��u�a��=Y�U%�U�o(.��{��rd��n�>*�4(�n�-X���=�%�jݬ>�Y��&fm�-3��u�:K���4=@��B�����S�}���З��h�d��坵b'��sVe���CfJa5���NR��*7M�|y6#�O!�y��Q~���z�	S*�.�����D�
�%�z���<����8��9���}=�73d7*�ʭ�����̹#��C}K(*>)'gh,R����}i�ꏴ����^{_�ʁcH�m-�\���/��ac�kȮ�^�2�����b���-Z�kk% ���>��-���C��h^��9E�ݺ���$r�ޚ]�9Ֆ�R:�WS����W+W,��V��Ċǳ�����rSR�f�Z���X��uҵr3.m�(���ZuFSQ[v��1)�q��ѶH��[�o<�)��w����ܙ��Sˉf�xxd��>�цm��������f`��Eڥ��36��z�����Z��Nkl����C�	���?,UQ�)�%��&�
ɳ�ii����v��19{���,�g�W[^	��l>@�<���l�ub)��5������u�<�8���ި���Í��ڑkh>D+���B��'�A���<�Z2w�r�� ����AԹ�}(78���x�VC�c9���9�� dP�z�8��5�:������GlU���Qor�P�]J�-�������r�B�d�V#ދ}I�:zI{��
�KF�x�����p��p+Z+t���}�)��}zy{g�;��P۰�>J>��{N�oa/�e��B�9@�QG�5l���;G~���Uud�T.8y=4��Yq�#����p��U[g��lI��j������c�G�w�T��N���m��l�ct���h�/�N��;aokPBm,2D+�)Lǯ{[e��V�(3������O8Vk�r[���$t��P���=1���%�¡ۯ|���q�\�J�$��!Ե�{i�LQ��'!ڋYe$!�}�Z+AC�I�
Ǯ����^ƨ��0��]�W5,/�3}�C89i���N`؃ ����'vm�f۽�Z�p������_:�o'+]���Rc�O7j��_e96\g�޽J�Z6�k�9q5:�ޅ+&�v�gd�r���C��sPt(�[�f⸓��F!#�^�X�κC��x�����hmJ�<c�:�hV��0p*�s�ySu�@z�H�����c#l�ʚ7���cL��3:��K���)T��Z��L�2SenK����Z�iq�4�Ovu7�^�'`�730��/F1�܄� 2�Xj[oh��z;.*B݁�V�
�1Kn�֪Z����kEN8v�[���/E����sU�-H������ ���+U5ԕ%�7����� ��QV�6���r�Ğﻮ��7G]8�T<���֣����6'`Z}ތ�eń���XL�+7Z�iR�vu(�-V$�rk�3��V�ж��`�3��K.\�m�d��^`|��b�,�蚴h�7Ga������u]lÄ3lԮ�4A�(t��2r����.��}��x����v�Pŕ'Xۭ�+o$8+�s$B+M�|�FN�#�ui���;U���^��R���:=5�B�x��5���Uq^r�xm��1l����������('0��ց�Ȼ�`���l82�f���w�f�J�Cq��9�l:t���Y0�9}�b����y4���j1�VֳjFU�m,�ҡ �}�t	�м�Ns�y��3*
X��������2�\R�?h���Q�X�2ͮ��>��(��[��/��;j�m]ꭦns ���=�j�+}�)P��
�8�Kԕ�g.�z�b�|r���L������#e�p�R��D �D<uC�Q��a�"h�wn�e`�+/tNM�����k�c�O�a�b�+�uY�1&^էï(ѐ�ݸO]����'�9���:n�'
�0F.���W>��%�����b��5�,Va��Z	ܝ�T�u桫����e���jC�o�+gL�j�gE�t!�G٨
x*P%����E�#[��.��4�;�,K.��.��S���!;�[բ�oK�,��Y};���5I5�:����'ʝֺ�:�ow�|����Q�����y��g.�,b��y|�Z���r��K���K��gR�(��l#Nv���O'��Ui���-��;,~���z������7�4k~{����L"U��c� TȺ���C w0dpZ�!VP��b�n�J�,k�kf�+2��*��WP��ƭb�RnT�i�������)��ks�Z�0��7Ӯ��1�U]�����3:ϕ]�[J�ۣ-[�
���78�8��w��S��.�!�M3#����d\r0�0.�T�kJ�%�VnWS~���W�!��q��5w\ ;�˙x~:��ʼ9R�7&_U��;�Υ��P�}�1��V:��<��
��`��!�	�ou�6�cG��OA�)w1�R7%)��T�,����P4jjRxtN��G�v�[Ԩ��3h`���)���B�_3mޫ[Czo�kKkr���I�ʔ��vA���[:�=<:zt� uӹ�:�3Αm6H�}�ɅYZ��m�gM](l�29��#���v�F��j��)����t�����Աۺ�ʣ\h=��g\��lO�(�|L�����n{����0[�� �	ob�x�{|�Zߦ��5zrNDq�����;��<j�����:i�*�u%��+�40�q����_��B�鱈�+D��s���nf���r�6K(i�q4�T�+v������Z/p��#�W�Y&�I4���45r+�j6]:���'mA�߫�5b�P�g%�.g��#Զ�㛭'پ@�4��m��� Ժ�]!��mDռ�(��DU����>��+�a÷wxA��*�9/T�ޮf{d�����u�t@_{���/�F=y ��fi�TT�M콧=X�28:	I���֭��Mne�/�RT��i��/d��4 /���6$ʓ)������w�t��H�sG�!-������pX��˕Ў�yȫk�9s�-9��'�H�ws���k��,�Eѡ��l���xM3�/|�(@b����)j��-T�5��n�u�4�.�*�ط��E-+������kf��7Q�Tq�b��
�3l:E�F6���s;����R�l��o�c?)�9���U����<U,�wa�h/���7�n�S�;ݎ۟;f�^mLX�F��[�vbv9�2c�\D<�q�ZlV̪w�#��6~�Ӓ����3�O�����y8�����Y���&�;w\�#�Vo��+7g���t7,�aы�S�I��K�,i�X�f;H���	��M8�l>��'��	�6� �Z�ڻ��m�U���5*e�TZ;�N�]Z�Ŧ��8A��9�rȅ>�;`��XWS�vR�zmhN%W�t���(p��:8ɼ���;�S�[y�67��)/��wi�rmBLz�ئ�����فy��*��/�Y�\p��f�����/��A��XX}3*���ۇ�#<2|��
aލ��E8��`�`�EÒ%L�kxF`kw�xg%�`�s��qA憅0gS����k�HȲ%�w6R�0�E���IxhQPx�J�r�Ŵ��>�d��Z�8��|�����6�?�"B��:Uٹͱ�Pl�[/zYT~K��`<�W�����ƍ�>ٲjE��vXk�qcÊ���2P��*viv�3Pc�*���G�P� �g�ă�W�RhX\�M�r���
��Aٮ�\P؃D@ź�v6U��ڙ��T2�y��C�+�Y��΍s`;Г՝r��!�
;E\s�x��㗆z>8��|���x,
)Þ�0�M
��8�K�1�ѽ��J�N�,�]1�=���m�~5�E*�.�+U+_���\�U_ej=o�]
�`�KR�S��eo���D�ً:ɗ�.�lE\㮱ա�Ïz[�1�4e��)���9H8b���DQ6�a=�lR�m�d���t_g��ZW|_<�h9��1�����X7�Gg�D9�.���}�9�Bs�ލ6�v��G1aÖk�,"�b2�^���Rc����N`�U�^�OwV!�Z�4kD�XzM�	�;Mb��Ͷ�PWۘ�j�]Wx:�w�Ō���룪'5T�����3~R+�Џ��I$-�����!e`��C	UJ鎔hw#��������o!�A*�m�[j�]yVhåif�¦���U�ӹ4��]��h�j*%�J���pQ��یQ�
3 �՝z�COJ��:r��n@w��m�x���G���t����!�A����ƚk�@���ܸDE�v�rY��8f�
�6�tElk�v�SA�J��@�9�J��(��(�R�8CP$q$c[Uwٳz�����|�VC[Xmbx� 5�\C&٠;��,V��$[���h]3xDW��羍	�+��W̺���� Q����v4o�J�����auv��f��LC1&t�V<ژ3�}���hǋ)`���^b�J-|]먢Fy�T��y�����s�y�]y�;V�ܷ�C��H|a�/g��b�^�LuO���2yd�Lu��&�{Y�L[��s�9��}��~�>���u�Ȋ�71�յ�n���8Ĭ�q����4���%�h�yx��s�`����ӁqE<�2Ag(�
].��f{��� �/gCg^\�l�87[A��/c�i�>�����z�Y��2����]���է���5	Ҵ�ۖPN0]*6�;~�LB�_]���+v��kL{R�)�u.Kw*�oP��E��`R�����~/]��#��\}Zz�w7���=��;q#=Æ�T��=����q5�݊S�٠��	N��&��a;����6�{߉������ �.	AX����ʲ�5���y�2{O�.~3ѡ�B�Ry�fZ���GK�[��IB��ś<���s+u�"�J!I-�V`V%�xw��(l��:�^��Y}܄b��AQk���wڒq�;���{ٴ�Q��x��0�r�Jl�w}F����R'���#��<�Zw+~���[s9\yY XVL8quK������iZ��[��[V�:�9k\����X�ml��F.w}��v�r��f�u��_+�OM#{�z��tx��8#����Ç�ݦ��:�J�K;2�[�5��2�<X<�d C��4[�q�j�s	�]Y�R�u�L����Z0�S*WL��s6�7�H&_S��C�N���7�[��4�2>ʽ�)7��EQY���/'�h*
��/1������tƲ�VX�{���j��*�et��f,�iڑ�gE�9ܛD�B)�����㍖6Jzpiv)F^�os�@A�o��vJ���#T&m���L�lD!Kzĸ�YJ�-VF�v��GV���T�!�1g�������V]�W;���4�C��D:�9�T�<���nc���9�v�Cow�4���@k����Z7�X���*p9!��e�B�f���k8,��\E:�Rcv�dZH�ݴ`�tn�U��2��k0[ގ����L��RS���+c �;b���K�=sq�[+�ʭ&9������nlx7�n�<�Q>�o���Իqٷ�v�Ht�u�g�b�Q�5�;q���G����$��RWU]S���M���ts���OJ��#WL;��A?��ZO]K�;�%.�0�"�ʮ�kNs�x
��Ǐ:2T`d#&�0][�5��U�fR|��N75@D���;^J]X�x�J��=ܘr�u��ND�|J�a;ڱwe�e��C}ԑ�FðsؽhTm>�1�Dq������&Sǝ���Y+l�8�7!3_o�iK���?;����	5wt���TEz�w�'`;���g���|>ﾱ�9��S���n��n��V��}{�!�k�sT}ZQ��;0�o��f�V��L^��J]ժ��2*�n\��*M����ԣ����H.�n\��W3� �B���7�s��=�O2�^����s�%����Z�K|N�t��X�����n6���o���N���f��n�&���5_[N�kI�N���uo��FV�ջ|�=��(�tw^���ʪ:���I��lrw�w��AJϳj�(�;MT�v��Œ^�e+{_8}5XWp��#����5x�Ӿ�Sۑ�*�n��:�j̫P\��������ʋ7*�pD��ѹF��!Oô:��CUֱS컲���iǋ��7�K�'��^S���Q��K��i�̀.JTzu�P�zuH]ȗl���I�D	붾߻r���37.l�F,�����2\d)��kH�����y5Ȼu�S��r��m�޽}�Fw���t������q5�����9m:��+:W81Єi�FV��U�>mS��d���`�m�b*�.X"�A�����B����0��T�;��u�Q����4�B4�Z[��ζo
�М��w�������D��-�]��Vd+�X쬫�3������0�XFV�ޣ2Y���r�ӻFwVƎd�؅�i&-��
�cj�V!�-^�hY�G��,�ǳ:�4IWj�N�u�h�7�JҔ4���)\��r��B���*�h�Ȥ��2D��������*R����Ji��2�+ )��Ƞ�2V�h)��$��*�B�2L����i��h(����0�''$�F�*��e�r�2L�����2W h�1�+ 2��)�"D�"i(�L hF��ʆ����!�2L���# �+&�@�22C���rhhi"���(2i)(������
2(���)l��J((k L��%�"Z�")2rr��ו�g�|�u�C�ީAW#%oo�#u��]�婥��Z7�D,�7+�X�\|B����=��'A5X::U��{W�u������������g��Mu:�>��w��ܦV^�D�:hX�z�bN����E���5~���M>|a��ӥ�i�c#���Ⱥ�����v��A�^�pyy�>�Kl!��)He���(8�ƃ��G�q���EJ���<�yWONo�c�`����go��������\����*�#�sO˻^��u�7�b9P5Ѯ�˼��tegH�=�!��`���
����v�Z������W�b�F�N�N����<�9
��7DBV}�ڹ�*��8�?A� )�Ͻ����e;��Z�����u��؎W��R�,�x>Y,cf�@�/D�-7�׮û�=Ś��n^{��5�A�Xc͞y�_z��k�茥�)�m�T��Ȯ����9ԽH�X���YXf㘤�`�¾���Z�A;�[�c_,&x5T����u�{K�'�<��jvR>�;�:��t��D2�iW��A��|}��yGF_�K%�*y�p�vf�롞;|�:uN�d�Ye=��uG��{�ت��7���Ţ�-���݂�ޓ�7v;�������/Vpj���V�ђ]�V�̤�jb��=ok3��j�/l�{@���`;ʾ����K��̎J+��[�p(��|D0i�
b}�r]^�fx�[�޺,��,&��{;=���0�Gwd�4:	dr�����̹�F�S�,+�x6�g�s��R�7���R��]�X��Kz;:�Yb�6�Ra�R���軙�!��+�*{���z��<��*�/s:(pnCNJ�ʺ�~6/ڶ�����k�q�w��SVr�L��R$2���T����Gjɷ^�m�2Yv�[��C@�Q��hgLu�v\e:}�X$eV����>�f���H��ʏ�q�}�i���z�R��Ջ���Ë��B��b�7\7}�E�E�>��|!�ickT=��z�6��G5,V:�ɑ䳾Z���ˊ�lc�GA�C��snK�n�LLΩ�-��KU�w)Q������ʡNp��Gss_K���Q�sK�ʇ��Ê����a��<���J�1U��|)8ue����N�>��hP�5ԁDz���jtk=���W&sY�R�HC�Q�&~3��ʬ�����&Yv>���|�:��=ԯ��s�۠@׹e���jWy�-��N�F�9���Aa�,w����� ;Î\Dg|w�.+��&�"��Y�\�:�"��:�����I[�y2��dr������U�<��S��^��m����t}a���R�/ⴧk;T��2*�py�k��w<~^�E<���m�o-�Gp�Jxo�1��$���N���+!���h��d�k���gg�M�p{+��W���欨<.K�#��\?xގ���<�f*"�j����u�S��lyM,�����%�{^��\���m=���.ҫ�4v5��]jknW�ࣛ�&5�~>�Q�=�ϳ�;'|~G���垘�:�`ƦJ�"y�{�JΰP�[Wp��z�Hk�5�N�����;�0�%k��V_Qcן�r��y{u�L��S]՟%�&6�r>a*�+���_�>� j�
r�}�i���]^7(>g�6'Y/]���b�������O��Y�מ�P�Ԡ#H�ÿ.�U1H�̅g��Zp�W^E�>����o�S��W@��6���ܺ�낇|�oJ�����ߧ>}�#T;)Y���oF�a���1���\1	�k>�0GE�ϧ&l/��Վ�r.W<.Ε�!܉����ѱ��!�YV*����˼q�7.�y��ҳ�����*{Y���Vd�p䳸{Ѻ�ٻ;��OU|Ʒ���<��\�H�S��o7x>�}��F�x�U��ucĩ�ӃK��u�.�SN1�<����h��M�d�d��zl��s��Ʌ���+U��F��t�JUbΰk||�`쇨bg6����n�����
��jU�,�/�C�;��v[�ux|\F��ּx�u��Cv�]冏r�T}��;�n�̝"�W�/Z��6d�_p��t`�<�g(7Ϫ2B���6�v��q���v��!Spe��jn��^�7�(Ǳ}�F�����B���B���M����;���*����7����+��c���:qˣ��R�,�bx�?3{�J����H�XE�m1=�Y0OES��X:,-�H�=��eg���~�5;ʥ!c�;�wF�C����0�f|�ڔ���N�T4�C���A�_s<r��~�!(ۙ%�7�*}�s�i�β1��/�4GڗQ"m�r{T�*�e���j���~:y)o��Q��֝�K>��3�z�[����n�ܮ>���΃�pR��S�2�[����W�>�[Y.Hz�:J_��C���n��5�v�c�}n�������R.��,;�6��	����j�T��=���V:]�d-I��)w;�*k��޾��:w.ͨ�&�V�W(Sw�grЉI�C7j��cT�gtG��<$��]}zWw�����]{6t�.���1|�]������W�r�y��Z"�}�\��g���6gd�J�2�t��#%Ȼ5��D�jNkk��]cշq�7%�ˊ���~���fr��X;0IGrJ�
9��>r/P�jV\#����u����W�$i�^�	�̼;#�=����)���[�'�����P����1����%�F��iա{[N�6���4���~�ۯ���йR�!��/��>�_._zg]�ϜC%�ȶϺ�z���g���5�\6�A�����ya��c�p�C��7Ӎ}���ƬW��W��^�c��cl-W|���r��仨��(��e�墨�!�_\�$T<a�����=�P�4�l�}Rzj�`$���+���	�}Kl,eбHHeڟ_KF�m� �=w�Bí���~�~�^��Fg���١��%aϢQ���p�:�/k�X.�|xz6q{ʀ�����͙Q��Ss�{�t�z^	��)x5ѕ��&|�!��K'��e,G�A�m�J�,y	��G-�����c�o���8�g�m�j���u�ͫ��2�8`��*�`A�?nm�Y��n��P�7��lIm��i��]��+S=ݧ¥��suj�B��F�4����d��~��<Hƻ|�������t��2闌l���Zz�F�YG	�=]>���9�<���$�b�\��k��_*kL�G��󳙽w��sVw��6�qHӬ���;\�߾����k�:7 �Oemu	C�W���H��jF��� ����|��]���O�I!&�8�fϼ��n����?G�9��/��`�>a���p�Wp�gT��+�/�&�vga`�]���a_��dN��|]WO���{�g�v].�V��n�u������i���пK��:K4S08A5,:�7�gf2�7���߻vw1G��QԵG�z;K�8����mYϻ��6y�i�\§G'���*��Ҥ����'��h��������Ydj*
n�l˝�K�%���k�4�?Nϫ���d?61u�x�qmS�T�e/��nXuԾ���.���)_w�=1���L9���خG9C�ؗX}S��5�A�Z�<3��J5�8�ԇyu8�n����w�ĪO�y�~��/�%�|w��ƥ8k� a` ����hZΘ��Ԕ	�wS�ޤ"Z��Uں+_�un��rWy.R6;�c���C$~,�K48�u�
�:�i�,#�i9�e��=JU(R�UZ�+Q������ľ�JJ�}yB���{w2��Ԣ����nag3��Q�y�.8�3ٵ���:M�F�c�	묃Y�{g8������L�VD:G�"u�s,��#�ԛ�ˮ~{˙M;�u�X|��Q}��M�c���ma�W@u?^�O�Y�{�w�����O7u�w�['�p��̨];Nm�z'���%�8D�o�q-W��*!&��{Me�盐�J,o���P
�e����x�̨zX�ÖP�ǥ��<���J���������
�Α�������WX���)G�g���:5��WW
��k7J\�}+�y�*W�X���T����xR���@~���.��ѳ��s�(��^"��#�o*1L�>�ޛ���\��_x����+}	�Op,I���^򸬇Xת=���K����7u4�n��&��UIm������ޘ�����F�Ӂ�&��Q��D"�h�n�/=��~+s|�{��p
��Xl�\�p��v*��*�? h��_Q�����u�sscr>�ύu��Oc&��g��"
_g�1O�^�
b�+�$O7ojVu���H�8֧)n¯�{�ZW��/������[�Gi<��Ԁ�~u�ʗ7OR�>
�B�Ͳ[�x�Alp#��
M���e�w {D���EPS�W��^��b]�J�r��O�KΛ8���Ɋ�OD٠��݁�v�Oi!�w�(���,\�}:���]������R{%ĻFc�T�%1�V�j%\���a�I3�M�oU�i�-���f�3�7hH�u���>��;0
r��ϽBM0�]:�������;�e�Β�c�G�!��}z��UC�@n�����b
���x�����S�Y���ZY�G��mm���O��
�(ul�����b�4��\ޕ8?����ρ}W��:�W�U�µ�9��X���>~*_e��g��}O'&lM���E���uY��+�������3Ú�}������w><v�!��W����3�qzL���Y�ּ����pvG���Q��pj���N������k\x������Ք��b�l�p��R�0@}b�/s6L�y���YHb��k�u�Y���x��
�n�����=.��!eW����ez|׳�Џ
���P��S��Hھ��Ɋ\Q��劃�*Ѣ�{�'Z�MGپg�.�U�W�H�fYb�_K=_�
W�0e[|����Ѵ��>stx<�^��R�i���}u7��0H�ەUu�:��p�5_px|M,jb&Wv�2oA�oI���x��<��}SF��|����>��w���%a��h���TUh�C>0�q;d���2^Q�H�iP66�S�x��5Hn�=�'L������H2�M
��]��)Y��9��Y�������'\qN]��^��Mo�+�������]��_�Օ��3°�}�棔�*���u���uя{�}4DGˊ�V��7�P�^Q|P� �oZ�v3��he�f��75����{=isC. ��[Dh��.��"U������z�=l����Y�"��	�܎�=�� ���N����u��4��˴��/��X����H��Ȱ�2�<CϤ]���-d��9f���?Hb�I������ӿ}[]vB���DP�/O��+�xӪs�{γ>�K�O�DI�`1�X.�{^m�����ա��Ț��W2/���^x�ov�v��}��2�w��-�����a���%<��l�\#h�x���Y���*'~�S���:��L�}^�`�C�e}R���t�bjK��}.x[��/�3��g�!��[�����^�f��J߶��S���\c
�-���C��|�����g�Ƚ����	-vf����Ў_�,yWz��/���iHe��2������=͇��8Ѡ���=�7qOhJ�W\n�b��n&0�x�����=��:칦�Q�0�v��k�bIH�Y�
~���kP�i����b��%�C;�>�)�]N���۩{�%T�n]���Ww��xVL�;�r�s�Z�����	�z�z5����ǹǽ�h{�μk�r�09�cִ�B
�� }����.h��Z�̄j�����R�E���t�S�`�I~u�"QE��w�qg^���,V�i�knK���iֲ�롰�g9�g6Uz���˗���'z��-�&|���*Y8��Rϑ�WҐAwV]z�Z�j��g{�wz���˞;q�N���j���u���ޓ*�(+�@������n�e���{��	�lՕ��8��]B:7/�Ś��L���}��8EK[����7�t,���r7*�f���u�P���z�BMq`ٳ�W�}e�U���OW��+�a��/�F��s�7��}�����c\�Ju��9���
����]ר�=R��k�ɱ(����}��+�d*�_o���!ղ����/2�����	�L�r	.fͱC�s4�Y��}r�o�}��A}�!�y��&_g��#ki�#����ڵ�+kmWVn4�ý���+�=��"*X�~��e������>�*\�k�0ʒ�O4=Z�N���OP�5��Փǧ:e��i��C3Z�rY���U�����0�ܩyԍB��2_E�-�*��olbԵ��tV&��o�;[��bq�]��\I�x2"c�ᆷc�88�r��V��wͼsl*$F��`����o7�8Zܒ�$���즸U�.��L�Ӡ�[Q֮��t�v���=���k4m\�.�.����ݗ��׬�p`T�մ/o����e��=m�`،�=ʹJp<!2���b��J#Um]�-R����b��%�xH�\f%FA[&�ܷ�|�`�����t��k���[G��K�\3X�I���S���֊$<�WE���և^
�;�I.�5\)i�P�J�y�����a_f9%��=j�wB�2�_���s�}S>�fn\����������3]!P�f|;��i/ɺR��@uk���͛jڲST�#�蝧��u��x�.͇N(���J�{reBU�&SB�dR�h��Pq'�k��X!���5a���S�H�τ�2lf�M��þv�:Y01��#�>��L�l����#�V5Ⱥqv}�ѮP� װ�@�IP(�}�ǧ�A���P̚%|�:���<�L{������y2)��P�Iᴗ;��gMQ�z�;&�6ݳz��U��Cx��Yu��X)d��^�������e:��P$���90�W��x�8̹��h� ��U�Eٝ����tst�����v�z;[����'�}P�ָ���˔��A���w�}��Vo��}[��$�pط�V��B� ]�Z��޽�,�-��rX}cU�J+�� rva�&/�����(�y�9�	�<9��PPv�:�TO:J�a�YH���+��c ��X#rg��9WEt��w�{���Q�a��mO>P[�/1��ұ���ymgU�HZ�]/C��n`-�ܮ�ts��6nk��ۗ�2s�����q����ivr�Y�;<ϰ��	4v��3��/��G�,N�H�:��;Y�\���J�>�n�]��ЎU{9�veۯ�\�)�4�`��+ ���Y��rۘ6E�K�!�ęe[弓��$eV��"�ko��&���nr����]����Ҳ��;h�(���)Mc{^��d5���@6���������	��a�u��vu	wj�}��=bT�
���e�ﺅK�^��������+�Y�0�i�W`�W�3%]��1�Q|z��=$ 6�f��]Oi����n�P�)�|;f̃�zQC�>5fJ�sC�ZqZT�b����0�-����M�/7����Gf���d;I�����*�{��٭u���q)1�T�Z��ƞl���6��{=�_EJZd�
r���=7RM��7���޳��O8��={�Ǐ�*��m�;A�@�mECr��Q�6��<��,�3k��J��O��y��8���O[�n�C����7�Y��<�3~�ߵ�Nf	YP�QK�%.Jd e��eY&C���M49	��d	AEAY��d�䑘�4�NY99!��FE�PRd&KMJU5A�BfVPR$IY�a�8T4@eHdU)��䔭1M%fbNf6e.E9dd%)���,F@eFHd	���JVda�����99�NY9��9Y�d�fa.�P�.f9%d4�N���d�A3J4&K�d%YMV`��d4Ӓe@RP�R�KAM�fdNHVHك�JDd&FNH�S�Y�ݓ�]^�؇�NO��ZG֚p��S}�3�Nt�YV�яe>��W7v�U���s3v�ܜ'�I�r9�L�t}�mt��{x���y�����8*kO��]s��ld�J��n3�xw{�n�����l;�~�oX��3���p���Ҍ���)��8떹r�v�E�BY{���f����Ht�e�q↥��	w@���q��]H�^�n�oj�v3}�R�//����.���}5w���V1���$g��Э�����wy��}Pl]�6�XT^���L���M���5��E�ʵ`u1ޞ�u�{������N���h�`��;ֽr\x��LΩ�%�`�ĵ^|�R�:��sop��l�u�3
���Y��y���ߍUC��>����c��\/�P�'��P�y]��r���<���PH~�nUKxzi�8ŝ���8� ����眑r�:����{���|�6|2��ބ&u���M��E����׬<'+ԪK����6x	�/������׫}R�>�frTX��/���T�g-{@{�bpXE��/y_�Y ɺ�1fu7i��K��<�������������Us�	����@�t�w�..�yk�B�1����P�zE?o\ZEf.���߁��xe������Z���q	Y��Ŝ"�TaYOMS��n��;v�&��ꕸ}���_:y+<��"��֚~�-����JXY�;�z���.��@�8��ht�8���v^ Z{^pW? w}�	Y��o��\���f�6t.��7^��C�bV���}^���K�Yԫ6N��;�e�wMY�x����>��1������������_!"y�~>�i��(�/އf%��ʈ?ޚW#�-?)��^�����C�}���sZ�s��R�x�uӯO���݇p{�֡�{��o��3C�LyـhS�!y�,��]4и�G"�\���_�y�N�^�f���G�^vc2��Vr<�#}�}�e���k���c���S$v���ٗ}�@��շ%�������k�׎��O�
^,����Y��*�y��	6��䧹w�.��b�>�-�P]��_��KպsO�'xƵ[�W���w�v'������c�o���:�r�^�),g��g�`L��R �u��TZ��3Pk����=�A�/
��5q�^�h��ܧIW�X;�1���n�B7�] ��+P�{�� -p�2< ��p��ռ��X�\8xC:N�-u�»T��1`ʼb�J�y(>eڮ-o��p̴(�N�f�=��a!7��ǎ=Jޕ���M�rμF��2<>ͫ7�ky�m�ϪU�1l�ֵ�j�i�U:\�ܬ��ЬW&Ŕ�&�!�z�|n�ϑ��]}�.3�����ta��.�Ɵf��]gN�t���eJHE��`q�sօoɏ@��0��}R��qD��u���ًҼ<�E���w6��O5����	��e�K=_]"�y�`ʴ=-[{@��v��U��>|����q!K(�+����S�̪R=s����������ʩz�Ryo�����u�>+���~�C�?Z�:ݹ�[~*�b1�
F��g5�)R�+�8YNz=�����Z6����/_�;9�P����g�b���%��Q�{�s�:�9ks.��߽d0���>�������/�(г:��}���W8A�3'���ⱌ�XT����ų�㲄��S���Y�V�g��Jp�.|�|�v�k�I�,	�M+��/���)��\M���w��*�	���"���Ny����ӿ|p�L@��41ł-�yiXbs_��u��y���}��*�k�	g�ENϽh.fHr�1�X.�{^m���NN�`ht���6���8�`̞�g��]�L]�p�%��j�t�gen	��۽��$pZ�f�-�HKV�Ev�ݚ����G%t�ǧ,���
�p�k�=������<:Ռ����7�,��J�'\�M����|U�_b�w4�ʦ�����Zr�J$�N������Y���[���n��]�kd�0Jw�K�p�����$��>��]`�x��OgUl��+������9.?P\����Ɵ/�C�s����zg]��hͽ�zDz���צ15b�e�����:���+��p�!��}8����\jy�����E���o<�TT('��xgTc����ˎڳ8jU���ÿ
oAr��u��]�:p�z	�ܾ[�������:��d]]'{wԶ�;t,V�e��펵��
^���P��j�#z�x{0t��SE�Io�ЇXaS�^�W8V�^�����]Z�0v�E3�#�X�x��79�vS��+�g�/���ϻMPN���[�L�(C�ʖN~��YH�N�%ܬ���KT�ݟ���w�>+�զ���Ay�+�"�Y�s�&U$₾�_l�S�\G|^燅_: ��F�|Qk�:7/�ř[]BP��+��<5,"��m=E;���p8�ۢcU�u�P�i�m�ЇF���}e��{���Y4��M�Pz�ׄ���[ʰ��{U/WT(�U��CU��P�W_q`c����θw�]�� N��.����;@�#�;�s&�3iZ��u���30gE��]��)�����P��Ǉ
�(��W
��}n��Y��C
݌W�O��䈛���:�>b������}$WHzcͥ�Y�%w�[CA�W��F����|e��#t�κ7ݺdW��{�4�PK��YS�!ղ�����j�}��ctY���#�/)Y�7�Wb��>��O��5�d��1(!�!�y��'�����C�����0a�.�rpM:wm�]J��jiB�� o�U��LS�ҥ·�2���{�m��m���}����v��y���z�.3�qX��i񔃮�1D��]�w3`C&�����v�uM�/=৵�����]K�xI���4�kL�\��<�����.���e��b��g�])?+��"�;C���L�+�㸇qCR��_Xa!��wAe׃0o���g�}G6m�v�ʛ<���&��x$���wu�&��82�X�c�?�6/79m3j�n�ve�}3WC��ލ�?QQ7xi������g�!�o��vY���"�	��W]���W��֭�s|�>&��v|��@Ȇ`�z����ܗ�x��fuHN����"z��N[��AE��>�:�"��nj�oD�&M��$<�^�Υ��@W�ik��f��MB�#XL�-^��~��=��?zI��OwZ�&�Vu�Ի\��;/����8v�#T���篳�y��o�F%��o�c�m�N�X�����n��1�8������[�T��
�*�>=,8�j��:�P�-h�\�\ݙ'��J��90�?�<O�Z)����	�Ѥ3�J��\��L)��ԛ͇*�7�j.��A�w��X2��#HH�X;.������z��/�v�\=�/ 2(w���bv��޹�FA�U��T�ez���_F(��;@�vr����Τg�z�e]	2/VS�,!�*���U@�K�>������F���G��ʺz������k��p������TB3��K��R{��r+�����]��1>ˏ�&�bŜ���������W�F���-+NyE���,��)ֻ0�J ��m���{62W����7�\����`�e���.��s���ևR�~u�5��,m󰶗�^�-sίG�\�(e�}����Ýk���r��N����0%ԩ筮��py1~Nd�h���kc�yAO���`َ�,�e;�u�[=֨H�-#H�w�#���!��Z�-ƚ���9��8���Y,��l^;���.!r��&y�?geI�F�W?w�H8ߝ{*=;V�V��_����[Eht5n���tjo�����e�`�o��Hn��X:�����v�=��]
�R�}�Ƭ��]�;3ƹ���k�,����O�����Sݜ���Y��^:~'�<*�V�q��h|��L�����z�)�����
PR �B�ȝx�}���X�#����ͅ��Վ�r.W��υ��s��lv�����<���d]Z�R_�L��z�m�gM��7��jǽ������9=�1\���FUˡ����7��X^<`Շ�f߫��=ʏ���i3X��Td��V�	!�·�&	�Wg�0oӠw�9@7���d�k��*m�y6��ZJJ2}�_�ˡ���OS�`��I�>�q��hV&"�zC�#j��|�[���3�7t�K�p�7Qò�_�Jg���e��R��,E,�|it��LV��صȅ;=]��������Դ�X.����y߃��N��U%"cnz�z��ȗ�0`�|ϑ!��`9J@e:��e�
������@Q@��s$��U@� c���5����9������PR��]�Z��*��{Dvr��������r\n�{KT;;h���#�2�8��5�jפ��g��
�<���E�f�ݢ���B'nK�be.۬8Cx������NI玼���$j�e�m���d��g��sU'�V3C^�gʥG��Ӷב�],ռ�"��q��˜��H.�'M��o������<�y�C�)��NԘ=�-A��8X���1J�m��#�v��),��ח��+�F�ʯ�%��}�E��䇩��3��j��Z+�LY�r�oƺ���x�����>��b~�٭���J����ߨgݭ}!�ղsΧ�t^v���������++���}[-�Z�j����6Qxo�����V�wg���	"�1�X.�����r�=b�P�.ǒ��oH��f�H������Wr�jyq�>]���:�����ͤ���
�*�s�u�˙ӊ��L`c`o���G����jK�C�r�|x#�p�����f�nǤ�3�!�h�G��k��_���UDHu�]���Lu����ï��m:�߬�����W�l�%�W�g���e��jUҟ_��w�M�Ar��BVxY��{n�}5�eꃙ-c#���Ⱥ�$�𞾥��]%˹�l��:τԼD����t�'N�4�򏪙�h;R_��D:����� ��(~X~��⫶����d��wR������9�F��͍˯�=�J)iQ���tdy�bK�՞xxS�%�}�CC�}�yX���m�K�tG޵�a�v�+�')�Z���:Vvh.u:m�IVR�e�o0�rT�[�8��E݇����?�}���|��ڝ�λ�&��+�y���/}u@�z������_B�T�p+X���g�<\R���r���m�|s�Ϙ��V|}SQ�g: Vj���u�ͫ��2�-�q��n���Ve���ׅ}��]��u��W?a∺]�ѹ��x�+w���;�@���@�zp��ۮ{`����jF�r׭k ?Nʻ	p!�U�W�m��w��U�A͠�ɓJ�݋N*^☹�g�+�r+�=1���I]��A����jȝ��X�^Q%�E�*V�s���>����X�!a�v�ʞ�����}z�-�z��2�;"sbz�ѺF��5%>��w]x.�8��\P�}Q�/X�z���MV��Թj�����C�H#�9��V���U|;��+�����b<s����k,��LSw�^�.{��0ʒħ��y�o�g��\d:��jFӤ�;>��+�#��5��}Hq�*zq�J��4��{��NPrpU)�q����1�C�����\Q�5�A�-i��iF��4�ZS#���G�N�&2�2A��Ψǡ\}�D�V㥵�U��</fu�/9��hV^��z�׶e|P��!P�Ƀ�]�=,Bv�m�1nf>���ܗ��y��Q�؄�[������y��d=vW[�g=͉�5x�T��C�]���σ��O5�Ѝ��S9-�B*�������Pʕ�a�:�1��"�P?]�)���S=���+�����-�]Ro��E��_t�㻮@M]�q�+�v:�X|__^�Uէ��7v�¸Wz���������aQ|z�Q}�E�ܱ��n6�����;�����ϷW�u����Z}G5Gނ��L��i͹/g�����"[��kev��t�����*ɘ_��-Ң�:S�#�?_�A��[�U���!]�eA��aތ��3�g�ݺ�t}��z��ܯ��k��A��� ��.iM:@�L�Y�U�x���h�Mp垤��������!�B`��t#h	��`��XxNW������S�é,䆋��c.��B���zߙFN���}�,�Z�:*�n1V�;C�B��9��o���̶@��Wڃ��\�!�ع4�wޏd���n`d��]@W���RnL�s ����'�nN��aG�sI�RjL��3q������kpW�����4P�����<��ۧ�
8����oM�'���2N�1���y��c�>Z�q�O�]Gr�ԛ�Z�	~�;���15�2��4��O�N����(J>�6}����A���Y�}��>���]���lZ���<��%W1W3N����T9��k�~zw��&���esy�~rwY��ӇW�Ʋ�;=��m'u^<m-�U����M�i�5F�G�W��uh��N�%F����n.q*�7QŉuM��ùX�u�ʚ�9��7e�9�kG=�L��gPwA������=)�aP9�2v�)�u��P[=]�ƎGl�ё��<�cw=kI{�j�������׼��n�ǋ�_
��M\p�?�ü��Y3{ml�J�'LD�	|;|�WO���3R�N�	ܱ��]P�<0���,���LY��mR��a(e�ƶ�s|�G��{n��7ҥ�����HM�m#�Y�e#`��|1Qf��0u&��s�m1��lV.�#�g��A��W�N�;�zҡM�^���d�I�'�d��=j�\*̼"�+�m���=��uqZ�4�}��]l�-�������/�m'����H��\ ��CX�blP+ã�Mݞ�.���|d~7T��u�M�Po�@Z��Wpg_�˅FF��Q�+ֆd9%]cn{���B����c.�\��&@~ݠsfQ��=�B����n��)T^f�����Zڄ����KX�Ør�լ�F����H5����m��a���ˀ�w��­UcN�P[x�齑����nr�����/S�vK|o�����[f��"��.���:��3�ws��i?KU藙���;�b��U�d&�+��=���4�LG0�������_K�/���$��-а����s�$���	;Ha쬓�b<j::�������C����{;���W����b���{tuc��	 ���a�hp�����Ιc,�8�dZ��ađ�E��j��c@�>j�_b�\іǄ���
�p%��$,��u�zR ���̪A��tU;(�0Y�t��4������6�ۀ�۰����e��Z[F�]�N�xcT���6����}�����`����r�c�aY�ʀR�[�9}v�s5��yd���N̞/l=�3�a�'�:�8h�z;�x�i&ޒ���2K:q*b,g:@lk2V���ٽ��������Pd�G��D����C����HS�����c�|���.S,ėjQ_Un�vF+r}�D���7i�r������E�g2Kړ�&��m1� �ҍ�b���3s���|��Z�`N� L��-�Y=�m�z箿=��2q�fTJ�j�5��^d�=3\�h���L���yCr��W��'���	V��a�:�9#�Yq<s��͒�(��s(R��)+�Տ�<�rX�n�8{�d�:W=G�����x7���J�6	UY����{�5���pgM�����ޖ>`Iľ���Q78�����]:��|�"�P��P��s%e/�8L�����9g|�Wn���*��p_`���ϣ���mĺh�y:�I�L�>��M@U��-$FC���d�e!QdM4�AHPdde�&BP��CCY%!fEPfbBRd9C��C�I�R�Hf`SNC�Y�CM%
PeY9P8E S4�FA�JS�%(P�0Q��M4�-f`%f`D�T+@S@QMRd��-VFS U	ҦJ@P�9P�QABS	KEfbP�R�P��fAICHP�f`R3YPұENf�1FIUA�eFFEP�-�AT1R�MeDIIAT�ED��R��Y�dU	NfALMS���TUSMRRR91D�%D�MPQ��15CSIP�Y�EFfT�D%KT��T~ M;`U����	���A]����]��9�n���`�V� ��ٸc�<2��K�rdj�p�:����̮Kz=��������v�W��̋#�=_��4;�����>�[�@d>A��/���dm�$��^�é:�'�r�_�����;���S���v����O�������j��#L=Y���?j/��\��磡�!���a+���ϒwA���o�5�zs��pFA�>�dn]@QGo�(uu}�5���]�_�ԞI��>��k}	O��o�hz���~^�Y�z�4$�m��#��D}��:���9�`�'s���y��y��f����;��2(}�QܞΠ�{��%�.Mu�(ܝ@~��~�A��غ�gXj):�#���y�}����a�SGr_��ۜ�f�}u7v�L��쟤�9��W��S��kOPW%�w�;��!�5���I��&I٭~�=���j�u>��wo9НG����0�`�K���"�~_@o=[;9]���:�}�|���������-K�BQ�q޴=\��5/g��x�^u����]@w	�a��ڥ��9;9���!��sN��}���4�ɗ���W��D~�Wξ��������}�����~�;�����7�P�~����~��K�����<�2w�4�F�)�����2)=���s���`�_��Hu��j(�k$���>��{�w�Ժ��y���r����>�Gڿs7���߶o������;��޾�qִ�'$���Z�)�^��d9U�d{oX�=O-I�u����L�S߸u''��J�?h�O��=�"������O'Pr7��:�/�r;��������������;����j{�������>�s�x���y��)7&G_bs1�A�jZ�)|�'�d|u�F�%ȧ���'PW��0��!������ϰL���G�9����;��~�Ѽ����o�}xs��?x��d}���!�K�W9���2��`n7'{��?}�F�;��ԝ}�@QBQ��
^I��}`�1�/:��;7�P	����\���s�;ϯ���i��-��U�uo<��в<@�?o� By/-s ��4nNI�%��:�.�&O�����=�
�`�����S�~���`�ku]}�'#�Jux}�S�=�5?��~���\�xD��w�%�Ƴ_��G��}��0ul��?I��h$�GX�K8Np91���˳ �26�QK���u<:1!P%��ʎ��������Ȑ�@�g��̦g��{�=��w�M�P�&X+�뢘�Y����v.��K�ݔ��
�&��1�q4��?�UU}Iu��y�����yBY��MG�{�>I��������9.���Z���r���oC�2y.��y��9&Oq޺��Z�)��uÕP�o�trp�;�=���I�0L�W�����_������"3�7:���_�"����!�!��dj�Ȯu�j2OӨ:w��A�K�^��=G$�W��5�yO�u�ֆ�N������'p�&�g9�aK�9'�֭�e�\�{�v,�o�w������We�_�� �@����F�������_'=�2�u��=�����7��������:��K�gRW�d%�~|����bj���@n2yS�δ�R���p�����va�tw���GH�?A��=�w���K� :���s�7X�\����%�j>������:����1?o�?I�����;���r�����%[{����9����#e�:v6ߪ�}Y[�/��|)���~��9��$�5	]��ѹ�O�dPw���s䚍���}��K�&����rL��2:|W��u&��QA��}'k�w�2y.�߷͉�y|����~����n~���W��w��8�E�	O�����r�����q�C����`rN��2�y��ܞϱ�|}ւ���5Pe�٨J7&�Q��
;��K��cM=G�j^���u ���^���;5���<�|��\��5�����{��(��L����:��2N~ޓ�aK�R{?��Ѹ�.K�{查���s�O�q�!��{�}�/��`{����kq�j��i�aը7dP�w����ֻ�����Wv}�����ϳ��k�+�2C����Rs����x<��7<�f�(��oG"�/d�����>��X~�4�M�~��������޹�E���?}�C���ݯ���\��}r���~��{?u���\]I�jO���)�Nu�VK氡+/�!�� �������z�u?I�jC�٩��O�dQ��O�j=��>��.�9�;�y&@}k۾�=��u�sGy����޺���r�{.���I�Py]^Oo��w�d�M��u��=�-��'�u�S�δ�G!ʨs�G���sY'�g�&[{��������y��I���U�k��_������n�5���߀�{��,ї䅤�f<���t�����Bu��i�m"t�/��2�7g����݃����oh�h��:vޝ�Ga�M�ɲ��lg1o��+��<�1-{")�+ w���G:T���<y�΁��|�z}��o����Y�9	G�n?��k�=�A�K�;9�&��jN�u���|�'�`~>֝�Rd�}֌� �?A�����R�jO|7��q�%ְ��r�w��'�y�=9�s���g5��߹���{����xw�A�?I�`��}�w	O!嫳>�y�(�7�4�]�]A���4���ԝs����F@j27̪BRh�Q�(r�O���Kx�.�z��߾u����s^[޺�=:�w#䔿����i>���g���/�V����'�<��I�{��~��*N���B"Ȓ~�O���$�٬L����]�Օ��}�w�s���e�]hJ:�I��^h>�p�x���'QO�d�j!ˑ�u��:�>�.��oKC�<��ރ��&I����7=��Z�	�����~�@�����^�I.{���\(:���}����3�CgYԙ>F��~�GP9'Ѩ?����ɳ?i�G �'g�ut�4�>�Qߟhr:��d���sI�%&���5 �{�~�g�盺��o~�|MI��)wjxs�9&�;��'Zy.@~>�VK�j>��gX����N}���Rd��G~��n��������~��K�rW�d����@
!���AW�֧_� 2!��u�پ��k���p����P�%>�-EZ��eP�X�'<��'�d�/�13���:��y/�Q�������.�s[�	�u&[��/`�>�G�;��~M�����?
��'����j^y�=F@a��u	f	�a��i����'Q�;~擩�|�S�;��(�u'=ތ�Pj�b�QO�d�9���?C�#�uBP0����vT>����f�|��y���d����hL�w��n{��k�����#��]�sI�7��7��;����L�/�ǩ7>F�����k�JI�j/p��J5?��A�rK��v_��O~̽��_��_|����q�~� � ���t�����ZN��`����Z)7&}�/֯|��'P����qO��;<惫�|�GR����?��X�����@nO�kXs����X��QH��]��A��׃�M�3p��Ҁ�ss�i�4W�|���?p�b�X�ym�հ"�iҷ��O�����q��qǚ�ݓhYn��U��w������S�K8c>�&�����<v����i:m��(oG�k�u���Uvm��  1oq:�_G�*�cP���Z��ȡ30ܾڒ��#�z�5� �jM�9�j����O�@Q���Д}9}k`�K�~�w���؞I�s�By��}�4=��`��V�}�����?}����4;��25߱���2O �Ւ��BQ���^���aA�r?@aם�OP��&r�����O�Q�k���y���1�(J:�Og_�5w����Hz3�����d 2>y���;�|�'���}��r�}<�pPd�ë-�j�e��)w�4&A��5=I�Z��>ˑ�r�e�dy������L� �����~��Q�&�'��Y7�?���:z�I�py���%=��v}��A�BQ�9���z���I�bk�\�z�'��p�C�2�x^��E=Q�����ރ�7&}�.�ί���� к�VoPoW�0���i���ﺊ{� ��E~����N��OP�5��~~�V`�&�����#�J}�����{��[�r<���+�8k����5����'PFI��h3��GȀ��E��~
��ۭ�7;��J<��{��7	k��/;��L�����p��;�����QG%����5@u�d}�O�k�=���N�e��:�����n]�
=>ր�� @�/�߫�K*~���ɗ��Y��\���Ø�b}Pd�Oc�{Д�}�S����(J2zw�q�A���G_�9&��ɗf�����r�o�|�{������h7yu�~�k+�?}N1�F�벳�O�*��S���������N���u>K��2����`9�Z�֤�L���u&��ԛ:�F�)�N��GP{E	�|룹<�A���9�K�ع4���Pк~�_�%������ǆ:�}̟H;������
+�>�nMǛ�5|֎A�nL�
��5�>� 5o���r)�\�+���G��x=C�{�^�����L��.kC�r5	G����h���A?�M�~7��9��9W����>�v������%���o���N�9?�u��n|�rϹ���(�Ptk�d��P���p���Od�6�����c���
�9.�k�<@���@�_����^�̮���T��ww��4�z�b��PAr�UX9UGf#�^�ϐ�"d�7���za����\#C�L�,�1����]�m��;JwSLu�ܲUMA��Fp����R垓/t�����%�<���F�����t�9|�������Ҕ�;���|�>�2ܤ���}�R�}��Թn^kÜ�(�ٮh>��%�Nf'�bwPd�O=�p��z�[�:i:���~��A�v����~��~���g�u��~��w?n���Q�w\3�����Cջ��w�c��^��!��j�$��NE�7�4S��rw�i�T?����Zz�s�ԛ���n�L�s�jwϴSt�W�C�u{��4������u�{>��A�@sXj:�������x��b���}�䛀�fsA���u]��Iԙ��߾�y��L�~5�'-I�2_���W��S�?��� A:~�ȗ�ߤ�'�T����S���?Aֱ8����$�l��#��M�Z��>Z��ȧR�n^Z��޵�	~�6w��������5��d�P����N�����:�? 3��g�����gr�Go�?&����&�ˇ�iF�:�z�sC�
(�:9��j!���h�|�4�Fα�N�%��:���5>K����7�BQ�}�h~��K�?�b�x�U������O=WHG��M�ˤ/��WY�Jz���|���&E	[y�n~��� �0sx�I�����u�2I��Ցܺ�����P���Pl:��O%�\��:��2z������?q��G�a]��~3?�|��ГC�O>�I�{�Z�������;�F���O#�Jv럺Oc�<�"��`j7'��7G�ފ�&�7���ѐo�(5;�P��E'Rds����>ם���.}�}�}~׿�����۞C�2N��p��i~�'$�;`n:��"����Zz������7����9�>�4�N��d��_�Ou��}��k�O��j�E��t'Q캵;�+�2�����u������wսWϷ�_�"�ù| a�J�ߪ�.E	G������O`Լ����X�A�{��;���0���R�E����q�C��c�}/���{���q�#�類��v/<�\�^�^����ܹjs�(J9N��T�%�tu�{�NT;��'ѸJu;;�s�������s���`�_�>�~�䚊;}���� ��~���2 $�xuǾ�*�5y6C
��TW��Q�i�p�~�:Z[Ƶ�7Mx%W���,�Kn���.MKv��[��J��Q�F�>����!v�k��Ep���O6���+;&B�8r:ō�+:PA�:U3k�W �3�&�G��)Exgc9�뽝*tj�|>������W�-��(}u�� hA��e޹��kZL��2uO�E�	O��}֌�*���m��hz�Z����u�	�jv���rry������`ȧ����;�������5g�_�_s��zy���s\З��{��#�5�eÞi>�s�x���05�I��؞�5�p��Pr�aK�>�#Pї�r)�=��
+�z�4d}���t�N}�d���ȏ�1lAo������_��ZYC��w���Z��ι�P�y/֯O����B_`w�t�r~�&������w;�;���%|aC��>�Plz��c�^u��v��22>��wG.�v~�w�������Ȁ(��sK��$�����<����~��7'$˒��yw�2~�-�:��xP�{����N@}��s�X��2�h��n�[>��L���Meڂ�'�}���}�����~(]?I������Y�����֞I����ur9.��=֨���}����:�'���t~9��9&Oq޺��Z�)��uÕP�l���G�~���{}{}�e���ν��?~5�$�ØQԜ�F�7����j Ȯ��5'��;�A�K�]������j�~y���2}���}��I��q���� �:�9�;�*������|/۱�����/�s�����F_�ȧ�����{�4n9���au���0L����x>G#S�x����j߰�P�j^��I_A��Y��]���15��y��2yS�7��sεf�o�s.uq�(�9��u�]����`�?��X�g&@n2^���u���
:�Z2_֣���c������O���O�e俿}�p���.���XP�us�y�4o����ٟu������������A�x'5�ʞs:�I�j��:�`���"���4=F��5�wo���%��6sz��� <���0���r]I��u��w�v����K����������zZ��;�/?�??~�szO"�	O�ߞh7�*��v��q�C�����4�`�g��s��Og��>�;���A�;�BQ�5:���(��/�5�4�?~�3�����.�9����si�}{+����;w��5n��q��n�l,�)�w�Dm���p]b1nd�*�8��weǍ1�|a�iV�f�OH������I�V�����w���C4���.>J������
�񵕇�}��}���__y�N��*5�d��/�oz�N���|�@n`�;?oI�0��Ԟ���n�˒�]����������'#��!��=�>��ϰ=���O����5~�k�~�>e�=l*��U��·w�E	GP{5�+�2C�e��jO9���cPFOן����^�x�>����;���Kx�/�a�1�@w'�\�sx�\��kEK��0��/�s�o�*�w�����Dܻ��>��ԟI���x_a�J}�a�Y/�����:!�� ���9�O����>�H}�5;�A��L�;<ր���MG�ߟj�p�x�����{�����]_��s��W�"���c�{���r�=�S���P~�.���i;��2u&���Bd�ɖ��ȵ�S��/Q�r��}��=��u;u�d�I�`�wS�u''��'�o~�?2?g�;ux�z/��?a�Q���k"��r}��������ÿ�����rMI�:���>A��0?}�;���$�Xg�����aI��R�jOz��Q�%��Z)�\����a2�0{�?$�	*f�ǧ����뮿@d��{����9����nO�sX>���9��)�<�v}��5%�Þi>����%�1�0Ƥ���n�����ʡ��I���P��W�W��z�����L��3�s���/1�^:�}'$��'�b��?K�o�4�r_mF��XP�G���*���o���m����J��0�~V.�Z�R�9�������>��\���~�/T!���I~����:�V���vP�'�T~sf>�R������O�<=8�ʄG�b���߼�n2Dᯯ={{��hX�~�l�:�"�!K�^9R�~�Vۯ��~F���+5e|��\g��?���W��{��z�m��Ej��
��Wkp��a�U�6]7��14s*�Sk���q~#
5f�T��/������Y;%�u��ό#�oրM�������5|�tw���l��ԇs��H�9�b����A��7���� >s���y�NF���eRA�|��*���*p�4k�(���#�s���g\�9g<Pc���3�г�v l�"���0�ۖ�kY �vU�K���W�G�x�1k"4r��=�%螝9����9Py┰j�/>l��}�Ȯ�ޘ�ix8��,��6��|suz�X�fu�1=�'W=��{An�tFc_!��{�0���ʞ�D:�X~���R�Um�[�r��Y�+��Fb^�.��	V�ƃW���L��z���="s�+�Ը�?NC���h�=�Sl��C}N��G �g19�(5dt��E���2��}�0�3��	+�޿p|v->2����v�t��gԮ����ʽ����T��uI����<ܧ�ַG9VA��}���)_w�=�]Ӿ��~���3��h+�ڎ�)�FWʚ���c�ʏ{d��B6��vǭ;�ȪRף�;�=CJ���v���N���MX�_���{���P��AF=B�4�{�԰&��nt�u�k��F8eb���/|�{;���W�<#�s����/���;��tǈ�c���l�Ϲ��1���'I}θ��0��(ߺ�N%
 �ƍ�+oq 7�~Aw}�L��;��_���}���9��;dV��c��K�Z��I���[Ԛ����wQ�ө�e5�6B/���}����զ�)�T]��x+��H'h���]��>�Ǫ'�>�"�m�QFJ�!͛�q��59��/>pʵ����5�t�"���D0;�;Nm�{<]M{ia�9z��B�8-��հ��c�z*���,O��8�̑��掬o�P�zX�x߹b����{���.�J�����1��Х�����n�X��.�Q�v`M
;'�OVg��<�F���`�ɝwte�:\a	+�
Z:� ?Q`�	�s%��J�WY~ק{���2݇>'*R��Bҝ��S������U�/�S��k:*�n�'���8�ݛ���*nN��
�P@evr�Y���9Z*Rv�R_�z����./i묻շ����>�k�+����Z���t��ѓ�<�f*!�b�[��n�7�f�ϻ�d7MUq-��|?a����L�pп�p~���Drc8�V,��E�O���S���Jb��}���;�hS�㰡���"y����Z���+9�_?�'�|�����Ι/�&�� �A����*�j{Q-=s'�,��&�j��E	!14i]�gx.�z25�M�oʞ^AdA�x 뮂�Er���I���Z�쒷�F��nࣨC��y{�TAM�4rd۬��+#n��5���A-�S-V�X����o;ko%�?�|� �w�svܯX��&��n}��\�ru��I�*(UӮ�l/�Ѭ
��@��WSW��5��M���!՚O�Ӟ�����j�rS���T}�נ(;$�}�U�=4��T��S�y��1�=b۾���K�2��ϥ��9]Y��~��5�p��\����Y�[��͙��h�g*��~�/�
p�XhZȝ�'�Пb�u��p�ҞcY���� .ހ�6 �.�߾�+�u�d��j�u�]�uy����W����wzC-*�}w쵬Ojo/دT0JQ�6�>�ו�zB���jUˡ��~"��D��)�YT��ov�ɝ���fs)*ꁿvI{YM�Q�5�8}A����oaT�d׮Ѻ�/��sw�xmg��3w����N������K��˞��*z���$"���8��_�6Т�"�ZSu�''�-�9s�����]׮n�u����/�����W�E+2�"�z�5�XH��z����kH�Vu�Bpu�m�7^�!�BvwL�w��5;�T�U!ܛ�+�{�Nc!�'@�:��Rm�q'�1��٦3�Nc�9�����D�z-���o)p�ԭ�L����,�F��)�N�s�nb�	�����Ȳ]�K�4j��֧eD��ȷ�c�%���v��7��� U�wB$�ng*��.g�(`��N�s��xT�[��x+є��j�����	GD��V2�˺��oQ�㧡C���	Fݶ� ��@�)�N�����[�<w8sE�
�y����"��A����tk�dU�1f]$��@��J1���t/�ee���;$�8�&1g52h�w����$
� ��� �n���y�����	Nб\����e���xZ�Jpښ�C��iM�og�K�v�+��;�~m�-��s]s�_*�/6�L�:	��<��z���_r�rn�	�Ҵ?�<��L�orfo8	u1�h�d���9=��S�-�=��nT��/b1쵛�����aO��T��up�9[���oʵ�<�	�M��/q�����X�yR��Q��u2����jwWY��_wP��tbڼ4�t��p�L>�#H���D��I宇�l�0��L[����}�ƅ�q��ힹ'I9p��]qO"Y���"Ż�H�t�_��WG�+Av�7ܴ�R��9)����/C�`#�����{� '��j�D6N�|�=b|;�=�-��΍�!5�����z]���Vo�S롗)��r#$B�(���ۡ���|����Lɼ@��qv��
3�ğit�������¹�;hl	�N���oGe����ʺc6r�m ��`�L�������؞+wf�sZW�{���ER)��7���~��=�(׳G1*���O���jeCO8O�$��7��˞���&Vy��A�=�mbp��K�y��器xj�Yi�\W��K� _wtta�s.m�[�Wf���p�I��f����Ѐ�ry[��n����j���_f�!��s��l>��O��X�R�޵�킮*���˺�`a�j={-֤��<��:� ���}���O��+n�F��k �V=ɛ�Gy<����ӦvY`�|XZ�s4�*���^y�b�VQuS����Nx�;$�<[\�eo�����!�6��Z/��*$�⼘ƻAS�$^f]ݷBL̘
eNw���y;^��:�UCC�m�m�/)�O��h�Зc� ��T�u�̙P�sԂ���[��f�퇖�=�#�І��S�P�Kc���xQg����[��ʷF��U����i������u;�쳻�@vgg�bJ�b����W�EDV܂�������p��9���>��;8V�i���]�鞬���伣�]X�|��bu̫�pfS�tH�%`�I�i��xI�b<(;�?wQ���Y;���Y��17��^(�K�[4�zO���B��J(��j` ��������F�i
�&�� �i
����
*��b
*�i2 ��������"������

ZR��b�B�&���((2��J����"�f�"�Z
�*��P��(��h���&I������J�����fj�����������"*��))���h����)j���� �2
�a�`��X�d���)(�X� *�a
Z�(��j����)ff
*&��Ș�a� �,�JF�(�) ��Ji*�iZ*���� ���(i"��$�*f"�(**
*��&� ����(��������"���B�����"e����(�������,&"
(i�h���&�hh&"���(�����(b(!���;����lFŔ�q��(�V	Ŭ�±ڴ�:���ʴ=�.�j�4w1�r?
�q՝x�wr����"�Bfqw����������7�ʷ����wF�AH�cƫ��� sfy\W�v�LOA�=�$�ZS�:�:�zV���o<��\'Ё
��[�\x�	���;w��8��ƕ�w�fT�ڭ��)�~/3�Ђ���py��i��Ͻ
�K �Bߟ���o�@hY��S�j�T��VO\c=�hף嵵�y@���R�}�ԥ�D�:d����3�Ҟ#.�c����Ϊ�q�6r}�;�z�����=[�`w�沥�}0ǛY����ߺ/;N�M��s8�	��V[�j��M�u.��<�ȶ��5��i����3�"��ȥk�>�3
�|}�L�k�{׵>��������dv�[�8�˰
O�U���a��G�{ボ���~=��Jy�����;�z��A�� c���ҩx���'I�r��r[���V�^���\�d��:�v8�Kϡ�h�k�w]n�E�;꺇����h�5g���7˫���u��"��k��$�޿�Mx!!�o��x���a�R��_yn�A/j;��hGzoa�K�=�52|h�HT1{*�U��_�8L�������+h��Ŧ[7o��������d
��P��v�8h�>�q��}�rQm�D�t��T���
>�)��V_q�D�緦y�R�,h8/����ݤxw{�k�� |ջof�1�8Wi ���VUVӭ�"u�����"�쓷�x_R� �|BAӶ�⪥otΞ����͵��t��֏��t��jK��C�8"Q����y"M:�ް���q�r�G{_#ui�����ܖj�>������]���Ǭ����yW�����^�Y��̍���)x+ϺE��?�G�����=q�&+}�p�m��5{c\�֫/�ey�C��o�&U$₾BXB��#8'J�P�t@67�����0�%�yYz�������ޙ0,�Y,7uBq
�#��Ûk ddNʻ	p!ԪޯK�Vtx�d-��[�%��39z�zb���j�/>l��|�7]�6��Y֖9��ё�W�T��ź���p����Z�A;�[�d_,&K�i
�w��VT�u-�=�n�Ss*]ؐ����y�֩@��ڃ�h9(�Y�����G���8�zD�Sd�i�$W3a�׵�s4����4��Ӟ��O�:939���!A�#�&0�=}W� �w��'=ٙ�˥"`c�<#�,R��j�Om���+���ez�S�8�]r�����Mu��HX�c��e���h�趒YN��/%�����͹L��T��P��q�����j�!d�5[_d���z-ʍ�{��;JWR@v��=�ݬ���ФG<�M��  ��a��{���W߀�|�ʒ���^q�I�NϨ�J�K��@)��o�T��3�b�^1s��:^YPE�+���s>�ɟ	2P�|���Lut�q�ؿK�;��{OJMI�]����x@um],�u,�%��8�ȪRף�;>rg�g�+��uc��g��=�'��{h~ʟlP7cEHȿgLu�v��z�_w���^f#�@$ۡ�m'm���V�Պ�bP#��ؿ
l�e�g�!r�y�},*��.���>�2)ْ�Oe}Ph{�/�2A����O�5�^HeZ��d���x��@mp�Q��;����^�i�����֥��-n���y^|�R�a:�@z���?��&*%�	v{�'p�H��z>]�u��r�>|zXq���vW���&_w��'�*�sL1gnmU��P�I�ޞñ�ӱmXڕ�W
���2�B���ॽ��ެ������Z$��k�Qs���)ρ9^�N_�iR�v�����uSG�>���O '�8˭vJh����c�'��z{�}׉n�٪;��K����٣|�A�8_o]�2�b)��f���b�p��э[s6� �e4y��t;�tM�	v �
I>������uʝ�Hf��,�y3yS�'rr>��m�7����x�[���l�xy��|>�}��=�3��z���ނ�Z`$�o�4E�U���9	V�����v����z�e�!h��F?�
R~�Z�!���j~�t���2��f*!�R�.T���c<
~0���¸7x}&������H��
��J�L ь�SA���[r�:w򽤲/�@�w2���߭���v#�.p=`-!��p��ky�>�G��ǀ�B�x�/�姂�ߔ�G(̻��T�n��΂Z���yy��=ܥd�}I��=ٴ=��f�b��]e8�t�@t�)oQ�}S����۟`ԘR�Lk�}�e�A�w���zׂ>������ 7A�%�y�+�p��SS۹�(B7�j8|k�n�����#M�ޚӧ3O��gk]R�>|�nrQ{_O��֘r�h0~�xP�񉊶ȿd]tb��hO�xQ�dw�<�`OP��]�lcn��Ԡ�q���Վ��ȹ\��)���|���ϐ~M��_������}��~��>@����x�x䶼��;�n����E���Z�C]n��^�h��d�_::��i��3���n+ۣ�;;�h��S�q%����CJϸfxWM�3vB�X���������+=wȩ�-H�L�R����Fv����X���Mu�t�-���T�*�
�Ԑ��2{2�(߮�7Kw;8��W�
�f$�
��1�:�^h��}��������{ �z��Cյ�=1�߫)�����>��%��=�)�4^�Qs��gn���S&���R��}�˺;n��Sm��e�|�=T�ë�n!���Z��V��f�d����At��6�k��G�5-�ʵ}�vtG���R�>�ŉU���$�m�f�bj��ԑ�W�*ؾ�����׬�+�!;(n�^w��m���*��M��M�zv�n��������
V1n�s/�|Ba!�T|k��|����[g�J�Iߟ��/�Xo9����0��#I��ݻ���g;3o�m�S�{�2o7�n�L��V�M����(�gZw�0z��D0��}U�F��e{[��#t��*�Lmy��u��}QyJ������W�;V�K������B�3>��I<g��[�ZS5�����}j��u��%���<��Úʔ3���ƽRo.�Kov�y]޼�$��ϓў�t���R�/��c�#�������+�a�nE�o�U�n�6sB��:l_v���t8�KV��"��r*�I '5Δ
�A9;�va��G�S�!ُ����[ì�%�_]{*�PV��v��z��×ӝ�yā�����������ĺ�(����6d��g^��k�������a}�߾�����\��V{��Z�b�{�{_��_CA��me���Kt'�21d�{z����*�iN*o��!��%<1:�~�F����PZt�Լ~<���Z���FM�w�ݮ�j�eA�w��\���zg]���/!�h�;_S��u��}�����캞���T��>g+�$u|�;Z���g�Ƚ���߿`���ܾ��BC2��*���W)~�~�l57ޏ=����	lT�	��u��]�:]�N��2:�Z�2.��$���}c���|w1Y�1���͐&J�b���hw��Ѻ�t��֏��t�Aڒ���C�9�e����f���=4�t��t�g�����.+�<=g��<�V?�6��_n <�4�մ+�&�ܙ{� ���O���?\����R��ҁ�m���/S�F��B	��Sy��������gs�j���j�k6�t���qA_)a
Lg�χ�W4x�2�G{F{-�2���s�{�����])��ti����d������*Z0�ۖ�k~d���!5�<��紅O�^���cԙY`�}�}!�d�
���ʳiǘPח��|5�]�����f��3R�7yN�ĥޜ��sC�ü���56�Y�p��+u�pcH���(�Ћ����8�[;��;F��K��_{썡��������o��'��W�Y]S�%��2�LR�{V1x>�_`Et��ǛK�,�H��	+�?{S�!�f����f������7�
a�Y��ﰙ/}����x;ueOH�]q�໛X.G���]��C=�S�����)��!��y(�C�Xc\�z���'��Q����{{Y�����>�N��	9���q�<v�C+V39���Y)1�O���L���N�՝*�*묻��|�RX��Cտ8Ӥ�'gԮ�����_)���\Ga���v3p���!
=��\�����0I��B���}l��&:���<k�޵��1�fs��}ד�U@��U�K�,9oi�}�ȪR��t�c�=C*Wm�5K6ukl�#Ec��]��@z(v�mC:c�|�R��ӯ�ˎ�󆑞����ٞٗmy�F	�V0	c�?�6/7� ��Y��w���aV�uE#����6I�=��=�ϣ\nK�����"�C*Ձ�������W]�B����){c�����p��w[�gs%G�G8ck:�z>׫	:��^�)b�.R8E������z�У�X�CYH����UCe�xW�r��|8\Ik�Q^����G�i��֞��B"ч/u�\^��u�]d�фP�����Z�߯{�}�����ܨ�i�y���eX&gTό[��|�^W��*!�ui���K~�]���*<c��粎M�i���C��	ÖPϟ�� ��~R��R�X���:�b�p���.gK�=+;��Q���Lu8,i�F�z)X+�rg]�}!�Bg��xR΀����uŠ�Hߏ���}C��){W�T��Jv��O\�"��k�TR/�S�0��c')�|�x����C�pxC�'K�W����f��� �p����Q��/`�"����s;y��7q���m{|5=��'�yO��TE5^P
\EϪOya�ߡ��������� ��*}��Oo)��*���G~�}DN
�V�۔�Ӹϕ�-����A;�,�׸{�_Ӑ�EUt�xޠ���1��H�nފ��`���ՠ�e�|,�[7g���T/CR���w��|q��׭��C��k%���%�Rp��vm|�ε�}����X3�~ft��Ö}�(A��zY�Z���e}޾�������@P>[�{��ϥ�Z�)�_"n�����z��/k%��u���_(&]���[In���mN�0m^�,��ĳie���
�A�f��g�Vi���9��^~���k�*����]S"��q���]�#�!X�#$��X�6���S��̨Y�*�g�������5��^�#��B7����c;�T�#3��y-8_��9C� ��a��=GWiu�<��;�ӱu���,�d�Z`��_�4���[B�ȝ��}��"���΁k���^�W�V �FT�93a4�c�r.W=w]V_�w"~�/,|���m:����
������v���k�П<9�3�`t���Xּ��E��Z�hCC�� ���-鰡�v��׎�����/�� *N��'.
�n�B5ۗ�	ٞW�b�@���E���=���]���H�� �Wʦۮ�{.7��tVS�/�\CE$-r�h�x�c�=����rШ���I�~��t���yP�����E�DU�^��{hּ*�Y]kn�.g��Igk�NB��`ʴ=-[{C׬�"!;(n�^w�U�A0O<^���v�=��ls*���\�wF�A��dF���ڔ���fޏx�mч�/ޚF.MG�ٜA�g�d���eA�
��T7�dt`v��z��1��\{Sg�����u��S8Pמ|m���rs�U�g<�;��5r��[�X��m���?$�Fj�2d�ܽ��]��j�� �a�Mv3��G�IC>�C���Wu�v̕�<��a���ɗg-������l���nօQb�@�w���������> �l��G��ܭy�z�yE�Y� ��r\�Zw�0z��D0��W��<v��d�Ro	�{�^3(Ig��9s���<~��2�|��׿T��d�+`ˁ�=j?o�2۹��f��hb\"�z�����_?)Vy��5�(gݭ}0�j�̆Q��k���U�Gc���NC��/��41��E��*\=_ZB�wo¼��n�]n:�[G��
���רBڕR�����j߾��Z���	���V���Wr^�Z`�IX��<�y�U�Z�>v���!��%<1:�u�,�ޚWPztσ��~?SFe�C����XY7�L��W��1D�����w�u���8�K�[Fx;_S��u���J��u��1��u�x���P?P5	#k��� ��1�xd^�mx~��K�Oo��5�HfY�m/$�n!&�	A�v�QG�?{���� ��ƍ%����ֱ����d]]�v�Jn�ڪ�#������k��9��b��w���h���!j�}P>c�p<>��q�~�����!]�ݹ�;��3>`��0�X���]�륲2�JD�&��&�n<6jq��'1��^~��m�F[c��3�S�t?wO�k�b��vB�fjݓ���,dX�r0t�v?YV�@�gm�n�������Qn|�!�v�؃>�!.^yKk%���j�G���I�{�|+��Q���
3�&��p��-/��zv��m�/+jZT+�DI1���d��˫��Ƴ��]�*yπ�V���O�K��0���ܠ'=GK�j(:��7i����V������i�y��̶b�;�����Л�Q��mi7�
��Y�de�F��k�K]�ƶ	�^���ݤډ#�9^ ��6���\SwC1zoN�y��I�I���e'��2+ُ̕�&-��t�'^�������"ٱ�֔*�7�>E�����Wjtx���I�]K4��&����m�GD^�����#�[�.�w:evSv�םoz?��j�R�ܼY��� �F<��ԅ�{�M��Þ��왝ϙ��,>=�F���H�>PM/�摹���j�t�wL[J�MZ���m���#Y	W�XKhsDɄ���p��^���jo�S3�1?=������;�n{;�|*ր��t�.��rH������b�͍{d��0oG�,���B�m�3$����V�[�vixGz� �܂@Owy�G�t6D��'���
FU�re,Ĭ����9d���NZY�AtC�p�3��6s�ǃ$�9u��G�%������6��b����iK�Ƿo�zZ���b�]��:Ζ���ա��;����a�Y��Ӎ�f��^r=�O���7�8\'h�lٶ�kЅ�g
��=�+Sy�xu�B����ݺ�d�zDJ�����B���e������ភvzK�(I�J�����̓�,ӣo��S��N�QVf��2 dU���}H:�m�n������R��Z7\%!:��(���ʝ�C�Z��4�j�R�`��v�����z�賖X�"���m\�"oN;ʷ��#A���T��б�n����O���$��s�7�B<]ѧ�Ĺ3���T}�+7:�7]����t���,,����z%�J2Oa�`0�t����j�ͽ�[AJۃ6lM_�����w���e|�ɷ�n��vS�0��Ӛp�hpU�<�����{�"G_){U����Aw
pQ\F�ڼ�םԤJ¬�*ۄ��Զ(pm���*�t��#�)�tW�=���w��_|k9�|�sf�%5��<���x���X�Z+m�n!XG�����(wcʒp-�& o��.�&�^�4�C�#1��'��F�
C�g �͖��<䳎�h��U;�=�GX��\�h�I7�����s���d�N�4���\�Y��ەǗ�-�Awm��R�;"kbH±t	6o���b���$���*(��	��hih�$&�Yhj���(J
)
(���"
i�(�)��*��UEU9�M4�TTD�TT�DU�DEUD�%UYc!AI��QUL���CT�$ID1DEL�4�IQ�1%QUSe�UEREAL�@Q$D�4�	E!Q��P�4Ĕ�T��IQ4UKQTAL�#ET�TUMPEDPE!e�IEUSUE1!Ed��IME4S%SUCEP!MD�EV`dS@P�RSIUAACKIE3faDKAUADPT@L��TT4UUU1�5D�PRDQUV`SQ,EIEa�Q9�M%U5QUR�ELA4�%5H |{������hy���fwp�6��!�6\�m<�[�+�)�a�� �̽U(��*`ѽ���"f΁����}_}�ղ���zu{=F���W�;Ҵ/��������$m{ˢ<�c�*��=��M��|{����U�tegH�<.S���!K�_HU.��9\g�\��,M�^Q������g��=z,��ݢ � �m\�I�I}ޞ������G=�����w�Wah��i��~q>T��T�Q�3�`X�d��6j��r0|o\9���߯�G<��]��^涚ޫ����B͝�I��WK5������\�g��Et��ǛHDǜ�gg�^c���rҒ`�}y�����PNǪV�5��g�O(�W����W���s��ey^�}�c����/2��҃E1��?��!ƾ\P��M5���9�ɥ�V`͆�o����VC�;o���M�֟��Y��Ɍ�b|�� ���{"����Y�&�U���^�/j�����yT��0ʒ���ӌ�.`NϨ��+�.�Z�!����Ϸ�l�`�`���C,J�X�t���0I�����%|;%�Ox��B���62�=����tUz�ɴ�2V�g�~1ĝ��%�%�$�,W���Q�j��^1�ս����{�/�$�`��\ic�[2�wy*��O®�ՌLf+�aY�ˆC���|��tU�ɤŏe��Z���SL���˘N;K����z�X&V����4����9Lc}����ٳ\<����:Ya�cm;�uTe�GHs�e}��/�"<W�c�T��n�ow�����`��b���k:c��GR,�6�pzݹT�w�v�$_�޹�w��V3�c���X>���n�����[>�2��G_����us�mSS�y�AŦ�Ge�X��/$2�}`u26��G5/y�������Uո��T=ֽmܞ.�,�fuK�}8N+n�* �][���}�nA��Y�Æd�P���V���`v��,��Y�a��<���%xB����ꥋ�*	��9g?-�+���T(�]��v�F��E+p�L�t��a��a	��h�9��C�V�K
�7}�z��F����y�����0�/�'�Xܞ�<FN�E�<3��|�/&�W�md�W�dj�Q�! ��]��/����WK4|g!*�>򰜫��������f��֫��.��bt��ހ�84f��Y�Y��FyX��Yܧ�muz���ѥ]� �l0F^5�ko����$��ܻw]�ٰ_Y��v�� ���a�vz��t��5X���pԵH�;���yŶ�o�s�=�z�)[{��m�����LtN�Ma�D'�Q%Et��u��`N�����=\���� ~��/w�ż�����Uo���t�U��75}p2��O���G.V��q�ӧ]3���;l�߼1f�BMz>_yaP��ޘ�?}z�)��1��	���R��'�ՠ�e�pצ�eiSI�l�9�|7�Å� ��x=huc��{@|�\�.���)��^�孵�v$/�}=g��ժ�F�U�P�]!��lp��O@��Ճ��6��f�u�~S��e-8�Gz���@cs�d��Ap�(Grļ�1��m|#��G��Y���c�P�{�%e�&����cN�K����S���C�Ş��b��_�6�b�е�:W���Q�YO�}u��j�}y���c#����̈́&��w�E���uY�5_:�,c�/�֬��frK��WO��(z�<9�3�`t�:m�Mk���
��e^�hu����8�T�\|����]]���u$)��Y��^�YM�V|����	ٞW�=�)
>��X��/L��� �O�����{��j���m��A�s��*z1��_m�
�C��+y�R���p��ء�C��P�R"cݱ{�����Y;�j�UaLZh�,Z;ev��:��_^�y���R��z���"f�9�g�.��Q��'�u7�#��1g�dx�+�L�n��u��t��&;�_}�������+���B��b���j����1K�,K~�}�u�GԶ�0V-�B�,҈D]_oz%6�y<y�z�4��+���k�KF����׬�+�!;>[Jv������3�ˮ�N�_ƟH��Ș۞�z�A+��'�W�ٞV"�KXNlA�0v���0i��m�2���	@������YP{�@���7��j81J���u.��}�0�ha\�MC� <���sޘ6��(�+��R�9.v:��P��V�]�M�YY��|�.(zf�K<R�B��Ϡ��8m�b�fO�v���$=[[�Rř�th�E��d�Υ7|�*L�w����L\��q�a/�"���sYR�v��N��-a���xo�;�N�;*>o=��;Z��C~����3�i�����'�i�vo����P��}ѯP�"����;�{���P�5#k�Hp:Fxw=tX��9d�y�Ӂ%x=u�Q��5�2H���1:�~�F��玭`:tϘ���� �|�u��͝`����\��&�7v�f!o�����Xys��'S]yi�j]�l�)پ�}˅iXm���jy�Ll��>*8����V&��Ѻ���ʮcZ��Gح]�7��]3�˨�i�2V�8H�^��YW���|U�[}$%N^GT~^����������7��]_~���ʕԾ�����\v�nư�/1m�כ^�#U���*):����묳�\�U4!����:��ޘ�9��`~��K�Oo�_Mx����]]�s�3���gs,�i����ÿ
o H._\�h��a���+�ӾR��N�
Vw{tXZ��ÜǗ�p|�[a�бH}#�^���.1��@�q�p<>�?}Hm�.��B��2��]{ش2�5�= �ug/zV����д�4;;���+>,/z�|oܲ^�T>�l�]�f�'x5ѕ��&|��O�+!K�-��3@���#��v��]�z�g�!�r�E��/)͗^���+"��tB%v�j�H����E^l"�Ꮂ��)�P�l�����������}��/5(�����cf�@�/~���P�:�&>w��V�qvWu��5�/h�$�_�͝�Y��F���s�޼�_G"���o^���ӝ��]�m��z��4��^XՑ:�|X]>�߼�g�(������0X�̒�P�0��}��Ղ4�'e#�H��^�������*ĀW�����*(��z�|�Ob}j�*��w���n�\�緪]��z��Uo���{���f�@M�a��J�LV_A�{eZv�q��6�Q��u�g@gN���Ne��kz����������黸�ߜC�l!��x��=����	��%^C��(��%���^�==�	�@������ ��i�
b}�8����fx�^�V��dx*X��ZN�]��:EH���Y�߀�G!}LTw�^�.{��K�%�=�6�i�~��?i_�߆xV�Ci��r�L��[���j��R�XuԾ�����s��L�%|�{�����VA�N��LHy~�V�]H<�ax��p����ey�4Gyv���EC���/u�F�ԙ�`�.��9�m+kv��,��_1�����B�1J6���1�=�K>M}:�]���F���T���z\�����G�V+�P���c��{�H'���z��Y��ɥ��9b�&�7}�E�D���E��B;,�6Q�C*Ձ���׭��W\�0�N�һ��<�;\�6T=AM9�%�.�,3�a�v���^W��*!|�N�We�u����;��:�-�<#��#R�iu�P�����0k=,?|& ���)]
Z+����唺�;�z�תWg�b���,�1L����bZu'~�dˠ�w��WFR�7eP|r;��[�֖ת߬e�ڞ�T�kL�0q���{���{<�H�|�{��[�a�A��
십�*~���
��ǣ�ٞZZ��0ߧ�����t��ӑQ��������(�We��-N�,�R��W&u�ї�B�,!/u^;��"���Z��m�W�e���Xx	��	/�-)�ϻT��2*��y�����};�u՞zܤI��������(o�1���'�ZN���+!�5�ʔ��{������;��7{i;�jʃ�代��8��M��6��Q�C�(�b�+��/fp���=��rf�=�q��
���{mT���mv!��s�끗=����#��/�䲡۶����8��ts����|~Gr���z&)��aLLu��D�v�T��O-�kE3ϥry��������ӿ�r��ys�#��}�C�d?:���s�n�5�f{�E���:_&��/�o�J_����#���V��$�W޶������͉�Kly�5���{�f��t�x�$����T"��B4� ��}�"��@�̫=ׂZp�zx=��I�ǟw��ِ�¿Pڑ��^o;���c�K9�d�Z`������Qsk|C�]K�pdգ��Z̢����Z�&P@�S��V��=��ި�uon�sj!c"d:�ތ�^%=��3p�w�%�љN����ͅ���>;i�{΂�e��V���^�|�'7V���WR_u�x�p���Q}�Y�ܠ2�$��P�q5��?��3����m����ᰭ����Xq�t�NL؛}I��r��.����|볎{�T�L�s��_.|�{�V�ȣ��W����͹��L���Y5�+��E�*��y)�sO�[kW�~Q=�ﺃ�V+�m���t��i�ozc�7j��k�Ps��ph�/y������c��=Dr[f����O�ݠn��ϾF�Z�u���ۮ�{.t.�2u�m{.����]���hh�'��@_0��H$m_P�*<Q�o���^)����E�/d�]-��=3E�_G��,X�Y�����X�U�yF�,"�6�����D��E�w�wmv��]���c��jn9�IH�۞��^���Ȍ)Y��H�e��o��v^�κٯ��9s��+��
��_��G���W=��R�����ŢP���{1[6���=;�~����V�y�����<C�x�<Q��.�ӥ�,�^ӱ1��vJv�ލ{wԠ���l�9O�g�Ig�]�6�0�g��o�w����d�C.����n�ӾeK�4	8�
���u;��{wX�,;�Ŧ�&^�j��'_(dZV��� 90�GP�Y���;F�(	ܯ�oF��񻺡��XI��NwqG/�i�Bã��Z:mm������KE<�Џm�T�2Uӱ��~��i�n7f�a×�����d�Љ_�)��/�&���I�3�zr����뤻m�H��mߞy��.�g�vmd�����y�v6��B���(xܗ������.�� ����5��n���AM��E��V}p�����t]`{g�R8��lp::u�s&�!u8�/U����o�����u���.�X!N�����eԱ�>��^��իެ������!~��&W�-��ʔ�MI~�}.y�z.��!��b�31�{�#5�������4�j�xm�O��+�u���y�[^��^S���W�v���3���i�
��v���O`���+��O�l%���n1�R�1�|���L���2c�۶7��+���xO}�-���]��˵��[�8�ƃ�>w�U�8�^k���6��c�CC�Km�H��轞�p�h7���������g���)�7R�D�[A���7����P���j�������>J�?\����äYKx��#����w/eS#N��`��%��G=5�=����7�͸�Yɰ+��w�P�ݎ��,����ޏh�3B�٤r����	ڨׅ�x�ā��*7����%
}Rś���n�E��׶&=N�At��u{c�"W5�]h`�u���U�vs��$�]�u�8���m3�p#N�6��*��ۢ �]ٹ�*��
�KU�� ��_��tTk:OOnmr�u��
hM9���)F�v<,���8�K_H��n��Kº�z�gr��U9��Z��l����C_�͟z���.����2��X��l��|�jn"�;�yu����O+1�YXe��Z��ޡmC��ذ������bϋ���߼�Q�ű�w;.�ʿ8�Qm��m��6��z/m�=Β����*�k�,��=U�Х������2�G`�/�{��{���:��6���ڽ�CM&C�z��v�o�����.~�u��e��*
n���s��˔݈.{�myƝ'�;>�ʠ��w;����tj���#)W�o�VPuտb�����`C&I�����w#�xJ����ίtU��;����F
�h+�< ��`�1�
C��b���%�a�G=�:����^��>f�ג��>;�w5.��,0�t
}[��]����p?h:��Qޣ �8M����I��ݛ[V�!��5<ym>�s�/A��w�仝=F:����z]�i��i��6��ʘ�$!F��i#m�A��<��s{���C�Z���^�	I�{���3�_e�(�$g(oČd�g��=/�B�ᘧi�s{|��vT�v�g��Yf����w�`�t�ӵ��3Z��7#�a�P��4�Ker��bs����L�Ϸ.�uJEc5�$�t/B�	��A5n�rf.��s�/eޚ<3�_zu�S�<��%7�g�D��S0g{O�xE9
E��_d|y%�)t}ǂP�{�7���
i]���5]F�1RV�
�b��W�(Ufȷ�'h�U�i縨X�#�N�b�.X��v����ݙn��^ac���jCB���BؤD3��fn��L������XdS����8��y|Ӣw)�}�W�op�hCϪ˞=��;�7���E;�����h�nUN�!Vt5�cw�d�m<�D�9�" ѷe�!殺�f�뻉�g��bLߤC�FQ��距�ҹ_.ǂ����]ST��R��J�;�T�ܠ(����f_Qm(?h�s�{��o7���V��dw���sPJH�z{�*Ӕ�v�S�{���ܭ� A9	{�q��wFi�&�^�ks���wq�ղ�,Y��q\2��K�O/�N���捾w�w��d��n)��ʈΎP��5��ZR��_S��M�Jmd\�.�}�#>1$ml��b�7
��l��zm�c|��w�]~�d�s�bQ���^|C���V+oC.���o��'�L
����5�Cm�Oc��G+-�:7ؤ����5���G3kո�R�f�-.x�n�n�4ڡY��Y���{��a�����9��U����bS����1d�';ݫ|��]Mo5皀��FOI�q���C=�4���^/UL�z:.�;�gI%E�wT׼���ڻ̫2���Q*�m�eQ��bBu�`���4��G�]	/o�����v�6w-*S�S/l�F�Ao��=��c��lÉ�-D�xhP�+�X����9���v(�j��qM릶�y���7�|$-�	u�?Q��|T�;���C�L傟���+'��u�p۠�΂v&2��ը�w����N�≕u3F,�@h�A�/sq'Xļ#&�C0�wi�htoNM���h���ә#�՗��4�Κ=���u^RM�ʂ�\jA@��&�	�E�9���d��/��=(w���oh�1������Ef���{��>\Ԅ�R��o�.z��Y����)�����\�g����ۀ��,�t��������	�d�{fV��(���5�ǵ1�Kn��|&��L��(,�NS�n�S��.�
BϘμ�#�4�t욇s��
�)��i,��0\�W��tA��/[�.4&�6�c^ƫJ=ŋ���Y�MI���{w�l��w2,�\-���nڻ�����$H4�U%R�QHP�%PSEQM�	E5TQU@E��8JQ�M�RQKMD�MUQH��FF�D�14UP��+AM5DCEE!ES�5ESTЕB�D4ELŖ�RI!LTSUVfCTRD�%TDIKALEE1AM@SDEU4&fT�eE%%,�EE1T�5T��$EP0HaU	TS��%!�AD�%E1c�L�E�SVX�AY9AMP�1E1QAD�QEED�DY�SCE,QT4fbP5�d�UDMdcP�LADP�UP1SUK�ESDJT@SHMTQHP�4Ņ� �o^l�����X�h�5x���}�f+��*����G�L��F6��A�]}.S��7�r�4T�Ϲ���J����V׋_Tg�M�(�n���Wy��+�v:����7� �����/���U˞^�{u��5���aV�uE��!"�o>�vY�l�.K�t�Bk���z�4N-���筓��!��B� ;Nm�{��t1`S:���p�W��*!|	����yq���sNw,�sq��_l��5�Fx���T=,c��(k��9�A����%K'¢�ļ��k��N�j9�u��~�ĹU�+�m�,��_L�Y�~�4�vs�f�K�!��ŔA��|�.�GY�G��Z)H&��0��k�k� ]0�/��9J�rzטw����8GW�2q����*��!��H��L[��o�1�=��8,"�t��qY調z��� Qv�姌vj�w�^uc�f��ެ�=r]��������C�8m?^&V?Xu�j�1Oy�I[����k�r�.T���x��f[����J�~@ь�^�pW[9�.��s��|��[��|�����������1N��0����<ݽ�Y��k��x�ϕ�����ީ�w.�B��a4$H*��c��㳎�s:K.�)2'��Lݫ��2�݆fj��
�������������-��h��7/��Gԍ�ofeR�/^;��+��yιP�Y�z����B�$�iv�u��e]ڹ�r1}�'���l��yDmvC���d����%�!Z��=e1��Ʃl�#��t�����C�;0hS�}�L=_Z馾��A�_�[�?vT��kx4zUl�~N�kӺx�W�9[��,K��#;�2��`������XuT5�_M' �r�Vl臧c��۞c�K.�Jϸ?����������[xP}��Z��y��\mu��R�/�Y���:.�NL؛}I�}r.W*����C�\�t�f�{��?uW�[�,��ա�Ic{�����u:�o�Mk���*/Y�fp��Ġv9L#�s�h;�@����Ӥ:��n��9aSv��F�r��zr��;���=�̬y��k)��,�7��#$!-���\`�e�8�OC[�7{ks3eR�S��FY[�����oؠ58z�i��}A!R��n����S�|������-;�����.�_x	��e�U�|M�**�p~*p{�ńXh�ǳ���F��Xv���{�l$V+���m�[d�;h=�!��N�9J�/�tmuu�Ou3�|�r�7�9��	J�cSb�:/^�	��Ӓ�t.�w�d��v9�>\�7:9�1=ҁ���o�(lM����8j��-*������|�)er��~�57�T�&6����@~����jP��ݶ�Mlݾ���s��M{�����ʈJv�I~�ʃ�,c<+��sQ�b��%�IZ���e+���C��o+w�z`���{�1]ג�p��Zw�1^%ֳ����續�w��/ZM��5�V��E쳂���W��G��Q�4�����2�|%���f���S��nA2��@;�����B�3=lRS�1g�ʝ���O�sޚh\|9m�P��(���ͼ�#�aN_L�k�����y�v6��P���X=�f�sU��{��}V����3����x�!��^��E*����oʹչ�ռD��ܟ*U�������}��g(f�C,�y�R���f��L`����e��m�x���W^��Z�vhw�8����E�z�0G L��_UԧN�R_�C�s̀�-��[�ܯִwP��}kr
�V�o/
�m�Mw����>�Y��c������?.��߽1�xd^�m~������ư���C����[�Dѥv3j[�zj��y�}}���+�a�Y0��D�ƪS�Z_[[Y��'��_��M7�YU��t�YH^t��Z�W�����}��|�Of���^\*ݷ#�w�V�T��SN�X3|*�v�j�7e:��{�,��}Ҁ�u/�{���Y������ÿ
o�0�K�����*+Em�S����==t�[�ӎwxO}�-����C.�����m�_`���;"�g�OJ�xeJ;��/v��t�PkjK�Ba��E��w�Y��W��|�,V��=&���~z_��Q�t{��v��9��׹)�/��w�]Y��L�/�S���
^
��e,�����͒��ss�r��syT��[�yЃᚲ�CtDf�j�xI�I|₾_	a
��<վ`��R|q�����b�0tՕ��U��[��W��R�g&���%���T _8�K�_��ި�1��9�z3MǮ�O �m�Ї6l����Yb�������Ռ_;]̂22�q���<�m*�H����iyŝi`s���_���!��,����J��5����`ו�{|�-�W�i�pv�ʞ�D:��ٯ���C=Β����%^C��Ҍ���9E���}̳��ژ���:ǤN}�g;��6y�i�\ ��C�fdf�Y��R�5w�N�Ӂ��oYS.l�:7��uj��s�k�	
Y�Rec@]K37�k�~����ð(�����4�V�u�7���O���V����l��{.">� o�O�S��r^��[�wS�%��וn�k���֌̝�޲��C�K��!�F��b���*\��S�,+��^4�:����w,p�8�C�]ҫ�Tf��Bv�:S�ꔲî��(�?wE�́�&J�ҢY<e-6=�@x���x{�2]d��oX����W�3��}4�>�1�R���ϥMP�;"�xz���{��d��;K�=_J�X}�:펷V+���F���o^G/��kUKdZ!:�y��6�#���$�ˎ�}5w�Ϝ2�X��u���$y@� �4�xJݴwۄ�ɽϪk]��O��X���ɟr-6�VkC�X��r������{��(Vd�x7��w��R�=�P]�6��x��)�S[���q^��R��nֱ� 9��R��ԃ�/d�/�����^2�>{�+�l�(k=,8�j�Eے�?f�P;�x�f3p�딮��_!��|�z.iM;h!2qfU�x��vs����⬈�x�z��E��"�>B3�	���� ������H�C����y|��9O�Iov��Ys�{���o+5���e�ڨ��,-����OZ8���٘/%�;,T���P��m�j���x}dԗO��3H�g뢱+�n�ġu�fm�n��XgV�1�&��=���B���K[F��[���@�gxwW�YO:[u)�J�;��m�!E�R����T�ez�CTM��bpXE��{ɚ?Zs�9+��{$�5���v�J��������YP{�K�w�C����jo����"�hy��שl����Ooo�o�K������a=�g(x����v*<f����=��7݅(��GCNgR����R���:w!�W����C<��1�u���)�����^;4fp;�ڏǋx�uߪՃډ�����fZ�e�v��չ�r�����vq�- ?��>Z׭
�w����<��_g:�(s�a�,`SR!�v��b���&R�:#w�!��˟d�W�e�
�����P>.{�_{�R��#aߖ�p�1��Q����7�.�>\Q�N�=�_������`�=Ω�OnxU��,�'��`��_�5�ف�Út����펺�T>�-dR��2�ߵ�K#��������^�C�0� .X�U���ܧ;��W�<���f���j��Ճ�A���/�L�>xsng���;�n�k^V�¹4_����YE�~'\>YG�,+~�6�E�vf��[I�;HY]%[[qXI�kZ��ŻS�W ,̪�Lf�J�6fr��i��e��ir��r*�׃�ɼȧ���勒'`�I��?H�}�m��s8��m��q΢8�/|1M*d/���i���xz�{�����+#]�$y��4VwP�e�cӮ7�^��G��saT���Y���������yy<�����+Um��/Yk_t���^߬��>��4R�m�XL�n���$*Y�uu�G��kҠ��˺-��}���y����}���,X�Y����+���l_K�mm�	M�����}���׮?4X2�i��ۿ�MϜʤ����.����aJ���窮ʝ�D���y��w�0��Q	��}j�v�I~oVT�c<+��j5���n,�M����A:��>F֘����WAgnz|������)�������P�\�+����RP��[���7�g��fu%�Aw%m`�aφ��q��Z�q��{9����K|x�=��e��,� �nR+�ɇoƹ���=�a�C��޵�w۵^�?K>B���:v���m`oW����r�p�L@���8�-�y��K\5i���cكvr��pp��J�tm���ڂZӴ3Z�h��I3�X.���Ųq�m񕢸���f����x9QV��u:��#z��-WQ�ly����ɰ�_+�s�]��7�d�S�q.��ĥP<�(�v���.ӊ���}1��o>��˟�3�8T��2�9A����oi�y_1�z��eBP;�8��"�I���^
�Aˋ,�y��Kt3l}��I�S����m+�m�ǥ_����\�W��}�*Ƌ����z��:u������\�d��e��x�?eA��X�	K'O+�H]s�-�=𖾣�f��X�
۷S��!tN��D���[D�W��v{�43�z�J,w�S���^R\VgS�|~�@�6=0�K�\нY�E�ؕ&���v	L�௯�|������Xь�)!�k������uႲo��^�U����z�o�Kv���HMjK��u�>�uE�����
����`��i�*vp��vo۾��G������򺗎�#���i�	�}����	3�S��ϡK°t��g�����V��*�O}����8�XS�F��@Έ3VW�tDk�77��T�qA_jN�V�u}���nxxU� A��Y_mJ�c}o>�yz)F�v<	�R��H�v'�R=^�[�T�;�٥֛�so���^D�1௻���}36����Kjs��eK����R����i�I�q��p�W�nf�ˋ��u�-o[;bս��w�f�S렋������!��Y��N��J� Q9���3(�r��!�)nt�u�mwm���}]�:�n��·6�|�ȝ�v���W�L	}�9�z����s�K�;*�+�����-B��ϪW���]!�6��m���� �?7aߔ�"r|N�s����n�;c9}>��^�HUo�ʜ=�4��c�;�P��iM�`L�F.T WY���Г��8W_���7�	g����<z�y�}���C���l#Zpz��ݲ*�z���g{'��A(E����~���#U�b���*\�~1�*K
���o]����J��oA~��U-�9�Q�W�\��������!�ua���.�}�!�6��bɧ	�W|N�=d�w���H{�N(�?�W�#��o�y�0R����֍(,�Z�e<}�*�,eH�[���y�C�ɞ���v�x쎻@1��"�P7a���c��X>���';(�v�s�NW�ԧɯ�[��6.;��&��8ᕊ�c���C�:����Ŭ�>w�z���M���aV'˪/}=�t�M���i���ls�t�N�7v�^��Lg�eṕ�I
 P��S܏2�������@X^�BIX�{�bm<i�;Tv���1�ڢ�dG�CI�/\��}>�^��,R";K�ym�v9R��i�������[���#��&kz��H��:-4�=��b����UW���'���s���o|�	��]�"���D0;��snK�<]X�uL�ž��ļ�lSC'-���Rü�\oԨ���5�8�~�]#:�o�W��|�h�߳�xW/���@�`�EZ'<�7�E�&z�J���&]����E=)�Gt <��F��E++�rg��yذ&��?M���N|z�����!I\|)tq�����(��W��6`>��&��uP�F��3��bv���Ȫ0[�U6E��`�W�gET����E�˒�0���<Oo��B��I��*�<g*S�,/��T���eA�ʪ��|��M���S<Z2���0��=�7<s��ܑ�P�5\��
��Xp���[��Ӳ�.ҫ��4^9��=�_��cT�>���g�Ǖ��Xd��>�Lp"�1�~�v1:����VP7E����d��t��������Nf���	���\�;I�޴:�_ν���q�^��s���'w��t�r��T�/P��ε��i��
r�}�i���<z�����p�ޝ�*eZ��TwQ㱻�`5��s�3w���&���Vݓ+ڰ�^SV�I�UL����&�ylK@;8n�E9�ғ5�<i{���W��k��b.��}�]�r�c�	��d<_i��:�ٻ�u�3��.�u��:��U2��ioϰ�a��s�qh[�wiڬ�-C�U��(�ӧ���F���N�;@Hv�=�E6n�p��2������b��^.����>y�aǤK-5�ʕy��Y��%8�M��ވp�5�8�v�#�n�U���v�k�-�˴f�`��Q��e�ۢ�c=���\"������OAgL�,7j�\�p)�o��y��gM�*�� �����̙���1Z�\i�WNt�m��T��賜pX��|N���Nθ�ch�"��g�[s�xU��i����4�J۸8%nкp<,sh�2qU�xi����pB��E�<��GY�guc���d���Ĭ��^^�߈L��]ćyG㎒H��=�7k6^Ro4L!^t�To���t�erY8K5�Z�r�ޥt���ju�-�R5�q48&���XU�*�n��ʁl�@�(�
:&��[�v;OL�Es�Z�$f�Sjh�V�p��v�a���w���Y�V����/k둳T���"��4oi�&�c3{v�pk�{$vU^��6�MU(hg#!ܡ�X7%���]�]ڵ9Wnw*�$�֡��i��;��=K��	Wf����5h���[��x�R��Q��ު'WD��]�;��W�M���V&�	��MYj��r:���@u��u�2�s��͐�ڲ�������n\�9U�����ly�1zRo���fPV�G}wڮen�Opk�[��m��mʱ�_��ۥXb,���\�啛}�Fڬ��9��7�0�ma���*�	x��v����6�����)�����-mg>X��<�:xkњ����z���Ӵ��N.k��,f� �&k#A��R�U�ɉz�vy�ޣ������D�ג���s<,�h�J�K��w���u^d��y\x� y�G���c�v�X�m��������n�/MIo$�1[W`J�����Q��ZL�cB�J*pMwX�鸔�ZX��8�����%-�'Z��+-]<CNM��?
fP8�u�����&;�W\�4b�^ݑ���j6V�I]wT�cUٷ;��.be{�v����OP�Ras+�"�k���㒲K���gVnTL�ZkR���^��J�#��{-YZ����i8�ߪ���[�J;hh�1c�A�JĂ�|ܽ]�$W����-E��J(��<9$AsDr�`�"�ͮ�>{�;.8Z���V�w��f]oe��#:�ˎ���B�B
f��핔99�9 ]݈
%�o�J�{hӅo���u�w�^{��5A��A�1ITT�T�AK�PĔ�$QAA5A5ERPPS5SQ4��SYaAKESUE5AKUQEMST�I$TRUFYILAQ)HD�SL�TSUE$T�QUU!MTU$D�PQASUATPTQQE%�DDSYaLD�$T�U1TQEQP�ME5LTTQTT�Q5EEPEE0D�5DSU3Q98��MVY2SDUD��UQ4�UT�U$UD�D�T��:뻿=�F,Y���1��Z�1Uʂ��[q4+�.־96�!���a���\�� qΙ�T8%u�fe�u�u8C����pϽ6���x#�>�@�_-���=J�caߖ��=[���D��}����U�=�`��_T�R��~�N�N�~��c�K.��0~��V�=c3����g��LSg?�P�Z��3P���і]�g��GE��ɛ	����r�\�/���X�0�ϭ�Q^��[��@���>*V�y}s���K^��4��kH�ޮ
�5���,ؘ�{���1\l�Fd�*�4)����~���t���i��D���n�`�c��{W�E��$��ᄑ���Prvg���b�Ch����7^��5B׋��M�W!�X{�6Nc����.W秩�0VS�/�C�h�랴+S_P"Š�h�� ���!38���V��I]�����K��L�^]L��VU�bo��WƐ"�y�`ʶ/��J~��S��w{Y}�n��7R�	�
BvW�J�_]O8���1S ���PC�?[���r����=�0{do��S�W-�k6�{��* �ۙ%�7�*@�1����
Z���{-w7��eR?Z�� �TܮP�c��lV���_f�K�F�6>�b���W*��޶����tp���N/NԚ�f
?v�A�m��IT\�]���Jw-������J��E���캪�/�D�F�˥�E�ځlr���7�<���������w��0����C�mq���z㳐]�X<����1[�q�� ���.W5u�L�0OṞ>�[{C<��K:`�Q}U���P4,Ρ%�K�ㆅ�c��mv���=�W��u}_sgԝ�$N�t�V���V�}hD��1q|�?����O����`�����U�;�YI_`Uk�\��v���mg�s�O~��;𭮻(�%eu�:V���5�����6\J���~![݂���|��3�"��es�w#�އ�]8+��lg��-�yű�6R�?^�������-�Z��f�.���L���'[.��9%�4o�^n���sC.{}^*Pzt��9e|~�z�\�N�ؚ����\�d�-�w6^&2ތ}�f$/��+U���v��u���`��K��!����:��鎱�v~��������L��
jqYJ�M�$�����׀Ґ̳=�*�}��}�����;�9/�ƒ��-w^�=k�F�����j�ut�����wxO�-����C.���Z7[n��)
�܄t�]N�w����I��P����tK�15Mjy�g�J�9_Eqw�������ҡ�A��0:�R�tέ��=�&�'�ͽ�r��^x1�=�%.�u�v�;����;x����솑�!������_Js�����j<Łr���5ݼ'>�4��C�;Aڒ�ЇXs�T��+�8����{_"�uc6c#���[ֲI���t�����t�某��z;MPN����ث�߉�z�_�f���9b.bj�yfh�=�Fz?�����9rϬF|�o�+ᚲ���\5�W;�eR�N&��r�[�,�1~�-���}%�*���3F���������~�,�[]BP��`�?w�f�c�M�{y����	�jF�r׭k 3���\t~��I�O��U��Qc~�>�ꗽ��C/�b�g�+��Ȯ��<�^,�I�0��~[aߔ��"u�W��)���+��ïT}��	���HT�!��u<$C�l5�f�����5+r������8�QRc�u�|� �ް�>7�hSwԾ�`"^���}�H�S���{`Ӧ��kN�۾�t0�!��*��kJ����/X�ҝ��Pj�{E�b�����s����%�����{\�K�Xqn�ql���'t�;�>:#1Y�D~0<s�����z�b����V�X3�ϫ��҃Ǜu�K���b�^�_Wk;�x�>�_6|����M����s	������)Յ�������V���S%;�}����^�t��4����ʱ���9>�tڴ��+�������\�܋�wo�|�ty���R�1{��Æ�i��T�w�-��{>�#0��-�<'���^C���n������͎�#j
g%�J�2�u���z��㶇oܘԸj�0��Hp��f�nםs�W����ac�.�&���&��x$����w]4�#�8eb��;A�A�B��$t���'��p��	-?QQk��>�`O�T^��!"�nXj�h~k�*u.]�T�����xWYD8����x���AT="Ûr^�<]X�uL1o��uo�f��7=�+&a~W%�TB�D��f�:?Wޖ�5�s��eC��>��g��|���\��I�{$0�C=pEے��Z+>�������sLq�;A�2qfg����-��t��n]��4+O��;Ϥ!Ж�e��K:��^`���	��.Ǝ���4�2�˿��K[�e��Up\�!�*h�W�gâ�F�`�~��V�>�x�^���Oz�[��5� ����R����T�ߊ�*UT�N���mtח#)^U�~��o��6`�*���3���h�s�i�w�2<�]�2�M��u����J�T2An OQuk��^n'n��3���CU\A�z�B����2�.}���6�-�dKz��؁�sgF+�Z�;�Sz�1*��e�>���{�0ǹ�{h�5�u��MW���.
�K��ڦ+}0��[�v�@�y�v��v�w�kyҠ���ѻF��+����"��aP���밧���5���7i�ޯͿ��e�a�~�����9�_;	�ߩz��:��4����ecs7�Ƽw����	���HEOt�0�S|��4A��NQ�ϼޖ{�<]�-��MSEƘ��_���u7�����gR��z��[=֨d����(o�[��k���g��n�G:��W 7�!Y�y�Z��u��՚��!����/��ZY���/���"�,�H��bzނ�b���ȿdN�e޻��},GV�ɛM=X���*���[��խ�oيܻ�VG|C!���r�e�˫Y�K^�z��6�H��)�_T�b(��W}��W����ו��!}^S�O2�ai�����ƀ���/1R����byU�}(���1ש�tv�w$>���ٞW��YH`M ��wm������}�m�a^��,np�pr~�7�����6���/R�d�g^�|zNҴw��s��h+\�kJR(Dٵi�o*<�G��w��4���I�2ۡ���(^�R�K��Ԋ^��pboW]�ʹreY��ɛ�C�x�/3������IN�x��s:m׸_��R����t�m}�;�`3�����y����6��<��[^ݿm[��N~�ZQby����OZ���zE+2�$���ׄqa�	�*�����t�}��v�	��6��7^��@��)e��W���Ʀ����"b�}w]^����ۓ�oy��p�L��xg����9�<�+�.�Ɂ=�R��7�*B��#�v뉫���l�9:J/�q�㚈b��wC��[����8����{H����uZ��Qצ�}�xžE�OL�t��W�	�E߈�󘤭�s���"��*hQ�BK>��N��Φs\dԆ�Nw��;�Ζ=#]_L�md�}$N�(��m��iFF]�)��/�$|_a[YV�r��ݼ��;WV#n}����ܾy�/�k>s���~yK�����^�q�J�<�τ�6��PPF�W]��+wk�(Ϝ��ȥg����ўWػ�i�����׆x9*�j������~!��e�e��2���_\﵄2`��1��k�Ƚzp��<��G�K��]�~ƘU2�.�F���7�!P�^�lA��Ss6[�$�ha~}-֣/�����o�����ȿ9n�\ʽz]"��� ���zp���Jv�w56����N��K�ǳ!��Ҝ�-����2a�*�ޔ.�Ȼ%s�����}ni⁳���;�ޜV�N���σ~?ZU�ǌ��ӷ�S��E��:�W���5oLHg��+��Q]����8����������eV���LX����+?}�����$����^JC2��v�Q��^�Ȩ�>����[�ڃ@r;ϠO�:��Ri�`�]]-d��쓰L��Xˡb��w�O��>v&��%�'�{�t��Ӿ�lk�Ϫ��v��t!�GT轞���,�^���^��"Ը{�t�����8>:����:�^? �M�}�.?Hb�^u����^<�T�f�c�W\�Ħ����S��=_O����C���ژۻ�
���6}�DC�0_����ϱ��<FIg��\{��M�"��������a} �F<�>=ߣO3���wٙx�������ɞU�Y���2�e��S�8;�%z����Y�p�xzl�&d��5�k�|p��oԻ�������]Y7쎋�<�>J����B��sυ6ٶB�x�Vo�1%�ط+\)�����Hka���Z��9�g2�*r���*s�/CF��M=�}�T�.�esn�[��7a�h�L��1X�n��V�78��7�?B���\��ޯ5�s�4�#ʪ�:�|^��Y�;�����S�Ry[�5�T-Câu]�o�-���S%�!���J�K��`s������&�^�i�c2�S̗�n�x>
����_OA�N��X�;*�����a��2�wb�"��l����l�|zB��_���{��#}C&��޿%��������{P	/WO��{��[>��(���~�*v����c�P��n��߸0���d%��1�Z�TR�"�xk��$����{�ɦg���z���W^��Ok~�����n��s�k{��Ƚ��N��m	��F�:�2�����>�ށ[H�6u�s"ǛD��v�I���"��۹�o�=�n�<�����g>8^2D��X�lz;��M�G���L�~k>�ىn*�8���uх3�'��r��Cd���y���y������٢C�M���xqk�;zo�\���;.�3��n�߷���TA�]��}�_t����]P�r�2l,rf�TKp��["]�u��R�X�ts�}%�Z�A���{|O����ä��ؕ�����%���.�%_��N���费�5!�; ��!bJ��t7����g�x�ݬ�x��{9�����jاtb�8!1�Y��.��`�t%s:]��Ϥovz@,�xx��T,�����^�x��n�����29�w�m�8;�uQ#��+1�9c�\�3Ņ��oM�)Z���w�)\x/xtt�<cݻ!̣4V��%y��0����b9rL��::�̒o{9�o9=��8��ŭ�d_�x|T���z�`��u[��ݐvy�;Y�褞���3�`�ύR�^�x��b��-�Đ+�{�r��Kel�����L����p7�{�D;in5�;v�K�v/de������+�P��m��c�����3��x���!L��W�F
�W:&��^l�2w)�[*�����[U��ハ]|S�������bf��O۟����{��V�p�/�Ə�%x�o��e��������}xsΑ�Orv�8�&�}/g/�N�Rk���%���9"�.����=�L�� ڽ�W��]E�Q��8@����)��CG��=�u����E�x�Y�wi��}���wi�%�ö<"a����7j�;2DI���1m֍������ȯ�4^K�D���͢z�#���=Jwko�=_���(<�� SZ����9x���1���z? wK]F�0��Jet*�kc�ҧj�6L̋���Z~�B�����p�l�]tX��sw�p�8B�v�O5�]�F���Vw����k@�%و.�s��p��%���=��',�&��<|�D�O]�����Oo1�:�7=�l]σ�.4;�-aQ�Q3�d�3�=���^����ŌO��Ċ�J��c�W�����ޓ{1b���.��,̺3�����V�:z1�B=�p�����������kF^�Qj�N6ߌ��c�^����<��\���X�K�BN3b��ۜ���𧌫f/����I�����p]CG���=�!`�N���jC���t��J�f�5��O1Q�	n�=I��޹X�Y$<d�9��B;u��`�Ք/#"[��w���i�C�n�:�}�j��c�l��G]�i�0���>t��e�S�c�[��e��.��-q���ӢZ���W�dֳ9- Wl"T�^#�G�c�����{��E�����ؘ��0���i�Rk�v�3=�c33�#�s����?#�7o��`����k�5Ҽ����O2�g�ئ<��k{�y�T�/8��ѱi^^]ɸF���o�u��%B,z�79%��:�^؝��{��v��W��V5�8�Z2�E�:۳A�)��H'4�C�ǚoh�9Ov�nu9:W�Wo1�1]v�ˮ�-ۋ�Z��a���\6����gL��BGB�4�m8��ڻdsQ�9�v+6ӊЈx�����Yr�_sH囘�Ǳ�CwGU�O:�O�x0w��nK�fs*�T�f�|O�Ґ��M�� �<���n>�s�p����q�`Z�V�ɣ���=��W�9J����4��=0K�4=������+��Ĩ�2���fv�aX-*��]�8�.S�;��R�ދ�1�"���˼�q =� ]�4���i�JK��e5��aZ3�`ۻ���4�c�C,'�F�L�z����jؙnN��<D�K�������ti-<Q(�uŌ���,+�!uom8������atK��S=�d���-9$T� ��l�ՠ��i��
�	��7���� ��3F�M��Yńe_V�4�Q|{�޽}�2�+�v��J�ܭ����U���EO�Y�-��[�]��Ш�6K�M0eG��,!b*�W������e;HC��"T��^�I�.�h������B�u��w��d9���u�z��e���qC]YG�vz�;���\Ev���l�-��i^9�u��80���r��lj��n3n�쨫&�&]]��M�+���MQ�uķ:�n������L���������{��z��5��g������7�L�|Z=��W�\+���W8���&!��]W�mS�Y�Vb�����,y2v/u6_��+D��5c�q}2���=�Û^�w,�VÆ�d�����ѡ��8�\gH�Ӈ�]o�ܬNݐ��O[=�jU�U�w*�j�9��wW\��簪u'e��c��h�Y�WÂ�{�Daݛ��|j�G5�*TF��-+��g�|Ιn�b���:�C�!wf�A�P]1gF3�u1�Nގgpr�/@ �}֟��ُ|Ɲ/��nW^!
���թ9���ۑ*p�Tty<���VȞ=Vɚz����C%]`+mĹ��	w�޺&�s���as��ESQQEQU3U5JA4�DEQD��QI1%DUTEAT̕QEALSfdREMME3U��SSQDEPREE1TPQ1EQEU1AD�DD�%EE�SS5EEQDTUEI4ADEE4MTQQSS5e�DD�TPRFfU�QUT1AR@EDTRL�UQQ,�SDDL�4�ACE4�TAUu�5QUMT�k2i��e�1U4QE$S,DD�4j\�(&A��DMAETQ2Tk0��*H��ߙ��uן��֘�p��� ��غQ͕�swV����q?qct�oI�����T��v����汣u���q��֜�Z��D��S�����;uLN_lOs�E�ƭ}�V|�;��x��ߔ����Ou��Q¤��������_k��{fqB{k���ng�eYw]�\�f0Y���m����u}^-�/�H�����<}V뷪9�X�S{{I�7Dd��oŅ{�G���}G�t�2,��N)��ﮗGU �9[���T�;�C�����0m��has1=�WH��*��Юt��0�n�|�ɒ�Mu��ǆ�Q����}�ޕ�ͯl��s��t�ro�ֱ<��$mo�\�ׅ	"��y�ݵ ȥ��K��~�}�t��������O��grk_z=���
IY����O�����^�����.D�5��nɀto}3����Ŭ��=՗��}{��=oȈ`�:5��y�co㜕Ih��>��H��n.�tzGS�ۮuU��3X6~�F��#��5�z߇wtɿ�!�8���o���.�0���v��$^�������vu=���O���~�{�ԏ�K0��F�T����&�n�{:ɽI+��:7���O�]Nx�����(��h[j":�����Hf֑^��]�:�y)L�}�=�[W���D/���rnx�M{wo<��*���q��Z~��Æ��c����c�Kzmq�C�;^q�?I��`pMF<����1�$p�"�G�m�"űo4̾��3j	���j���C��rQ�O�ZP�zU�E=��3�,/��G�rߪs���}}x��&����k�ޡ�Ny�Ӛ���M���<�[R����'����*������/��7��H$��kX��j��My�N�Ҋ�X/}�9����a���m�V�&�\���ص�qT�n��:�	�^:"�el{�����gjU0{=�Zޔp��;>آ���Ov�
}ǰH,���|O���7�����$�m���>ϵ��|�?L�T�/�����zsw���=y6��1���
�~c{q-2�o��1B ��ؗ7(����~]i��|B��0�[+ n�ݫa<z���ʁ�،�R���(k�~ZC�����~���__i�+�-'wܲ�����#�U:�>�t@zy�x��Vk��:���7}Wn$Aa%
Nr���'��������ד����\��؜�fl|�K�W����d����'޿���.��u�5�{',=���_I��0h�jc׼�Oa��\��}���w}�	��ݾRH���}z��<����5쎭�{>׸����-�3�B���1	} >�u�����1V�׮��=V����I�c�҇��>��LJ��/��D/�g#�^ПVg�t�Ϝ��q�=��d�(X�_x�q�L6zm%g7f�R�����S�Zn��ɕ�1�`�ߤc�U��.�v_���Z�zc^}fϺ`9��c*P�)1�(0�}����"�V�ɗ�垷���׆H��������rfv��x֬�P�N�lǅ�q�߫����m/0?q����S���$O�}��Z:�}u x�Q)�v�i�����^��1֦Fg�gs�r�d��j���od�i:�T�gd�(�4��X��P�.
�;�V��e=6�%m�ȶrˏ��>�z���?j�3��o��;Z���s	�y�zN���އ[K������p�ě}�����˕+���p��?}�b���D�}�8������_�y��7�s�
�{`��ݸ�����r�kS>�'����=7����ݳ�_gnz��o��~'ܔ�I=Fkw�3�42vԏ&����N��]^�{�5�b1�f���<c},H~��o�~W�����o��A�o.?K�S�*�۷�L�=��ev�>�+�m��س;�z<�^G�G]���a�<�b"	쭸�H�I睟T�f}G����|L6�B7j+�nY���g�Fj��Sd�=�=ȡѢ�\��ϟ�D�Ԟ�ڥ&�uz�;�o��t(��3滢3g7�>��W��#e���cы����}��}3��6v}��
m����o!���`-?M"�˧FI�]�/'���x>���@���~^�}�5<�.Ϥi_�sk�#���!�e��7P]���m�"*���J�A�뤷�f]��Q�s�d����)gd"ޮ��^^P�}��~|��{��RCG�HG7m��KeΨ"m/�v��x_��S���]o�S����?>}�Yn��u��FbDo�|�X�[�^����U�0:?h�Y�Ԗ�_��'��zAg�~�q��Z���^��	yr���l;���*;!D��Rf1�P�,��&دOf���~H,G�/���b��Z��3~��x�e��f\����<^��֒`���r�_�8���,�¬xzy����������_�bɮ���y3�ތ<�v�$���=���,/A��_����Z=6A�����d2D�sԏ�{�5���H��f{�3F�����H��J�e7U� X`:E���m�����ހ�䓽X�]�vNs��C���ǧ�z�z���~����U���zD񧮷�b<2�i�z0vs�)�n*�炞���C��n�q�-��y��JPy��3}*]<�+Q�cQ����u�ǐL�����
T�p�z^�<%&0v�ie��]���,/r6{.�/ض�����V��'��/�\�m�UVn��yG�kX�5�3��Ǵ�����
$ܜ@'��\q	ȪBc�Q�k,�viV�]1���,,�Zê뇯�V�2�c8ܗ���[Ԗ���ٌ~[hw?�6b�+���Q���!�����}���#k:��ׅI�C���Zsx���xL~�޻s��)��S�'�	��I�MzPڰ��'Z�gz���w]��S����_D�k]�&��ɝ��������د�,cXr������X�9*�!�5<��\F�T�[�z#v���Dmg�;�gä�p�cE�N�k�<��
u�^��g��rJ�z�<�oK��ϣ�����Q�`78?p�E�cώ{�^�鞸�~g��/7����Ed}�98!�F<�p�����'�{(Ks��j*�䖜�l���gy}�B��w���O�����뛘�7z��ų�p�����a)���xv��6�}�Nu�x�і3��Z���w;��g�e����x���T�[�û}�Ƚu�2YH���W�a���#��ܗ[�y��=������meIp�op^��d����kw;���Z�I`T�Fʒl�d�Շ���_b|e�a,s�PO��L����O���gmuԻr�틷��|�]���7y!�^*uw�۝)�	zq9;J�����䚞uq�>��wpzf����g��d��C/Ta�U6��B=D��f�ɰx����d���6��O'l�N�m�?�ݔ=P;Rne����ۜ���v���R8�Ov��N� ��^_����{���c�{��v	yfM_q��j}�ޏ��}^k'}�Y���ق�,r?y�^��t�4߄�E��w�jw	)���!7���'�Ⲙ�/%r�e�G�N��რ��_u�ƻ�9b{-I�o�3
���y{�]���f_=�^q0I(Ϲ��y�	�.��}�� �*�F݌~��Q}պ��2�\�o��^)�"-�<���|F��T�rǞ�<lg��k|��3�<޾��Ɛ���p�.���%�)��v�+]�=�9z���,}�)xvm���^�xH��$��|:?G^�U����À[��4��s�R��Y�c=R�u��S��~���Kp�%U_,�ٓ�>���-�(2:!1A�5]v�ܿP+X5.��uO�:W�}y]�)�7��2q�
�����G]�J��q%kה�������Өj��u�ιz�b���!yC���1 ��HǦ},���p��� ���]�W��z��z����Ϻ`9��P���L��(L�Qt'b������������D��̎�I�2!�,t�����o�������H����O]�yFh�ѳ��%y
��j]$�K�{��R�*��t���	���$z�Ow�3�Bx1x��Y蘚���i���sͪú�����ί<����"�Ow�����&�*��OɈ��=�~Ǘ5�h�bѓ�/��N���y�%������w_=�E��\����M��мipa^�"�GtWr��&^L~]���o�ʋ�p��c�D1�lxi���G�^G��5p�g{�����c���G��T�f}D�L"ۢ�<�G�yЬ��~��T�l���+ǾZx�o�`��9�����^-ǘp�-L{e����罪�r_�k�o3ጲ5)U�$�����W����>�	���	��������3���]w�71Y���A��p�݀��i�v
�=FT��V�6'`�d���I)��o3}�'�B=�'�F��+D��ͯ�=^^�Ը�%n����cٲ�j�����)���4�c4m��bR�|ew;�6��_x>PakK��h�:6��!�v8�'�E�.��)����1��a���w C���������Qv|$j[�3Uc1n�5��R��a���`q�@�(��W��������������u@�dg���D�N�����l�!�Y��B���e��;�+�Dz�xg�J�.�� �o�Z�W�X�uV�c�zM9�Ժ�V!�9ټ���0��Ͻ��p`r=����e�¬M	s�m˧9��qo�ߺ�~̞_a~^�a�n��I��C�g*ܝ�
G<���zi3���d�G
�w/�͡����_�'��|����v\�V���<(�N5�+�����V��/oϮ��*��z�`n/rW0ڐfo���C/�ꞹ��w�]��!���v侪G�;��W�ܗHz��
l���0�ܙ�Ś��ݚ��E��:��.�8��-Od�:�9��/:��ȿ3�mW����o>qÚF'[ U�}m�:
΂��wãe�ޢ��zW����}��Nᇯ�i9u]e�U�e�����i��a��Ӻ����q�}^�$�Żw��Nv�A�i����'L�T����p�?X��ɋ��n�������luӽ�T���~k�ݒ6��ιMxW�Eq�~�~���f]Q��������~���'�<]�v��_t.grkBkҾ}��;��f�)X�gQ�]��B��;vL����
�깗d@++D}����Α�S�HE�E�g��X�9�
�.ѩ�Ƿo��VJ����J��N�����}��x<:K�%g���=ba]�q�-�޳�5�gun�4��5MuszB�D�,���pt~ќU�/��S݇]4u$$���9�VY�l�Kt��1�1�DvǄ���)ν�v�������K�범�{	�b�r�{V��g�����{Z���":	u=�r��Tt�q���H�!�OW���8�(]�`����ltB�!���&��np�m����<ل��F#|���=�,���e��-��ːV�Ǽ�TW�E8�+6;�	���1V��	z�=�����v*�[O���9`�zF���&�'N�n�q���b޺JU��m�n$�,w|�$r��t��2b���ը��%�o1u�W�n���|q��އ�$�d��hӍ�&Uk{3c0�U�4CO넆r�5������}��Zڶ�r-�5GA��U��r���'L;z ���$3�������Su�xm��\�a�d��;�A6Y��epx{�9؍�uCJ��f ��}�a��7�������t�9��u������7���]�/u- ll}�	;r|��3i��T�cR�cD��d9h��;[�ʃ�S]�aGo/a3;�����N��s� �.bn�w�Z<���17�4Ŗ@UӨ�+�#�2�[6�uc��^�(�f��x��`c���r��+��M�5�`H��4��WIt9z�����̞S^�c�'I�T,�������7�Sf�钊K�V��1�s���u�єT�\E��v���ٲ�a�-��q��cv��y�|4?��Q�Qt;�	t��[��-���X�/M�^ٹ5i	�Ǩ�ӕ+�b]�58t�ľpK����Ӝ͝�$5g�����܉Q�3�Lܝ%�Ps����"ۏ-���O���v �@�^׽��b�.�/��@�S_Zm�@F�aC�	��	�v2T�it��!��2�k�|; C~���������N6Ws2��=���E���os��{[��>�!�t������3��q�:�M��f�m�==s�U�.�3ܵg6�k�Z����M���6��z�ت��\^��Gmt�N�GVJ�/�O$zw�����ǫw*mb��6+�&�gkβ5ŵ���\E`�v�w���m��C,�;�P[�^X�+k�-)���@�n����Ct �+��Zqu^N���K�[�)�Y��^�5z(�� ���Yq9Ã�w��{@&"^�@(e�{p�i�W����l�Fm���7>��S��/���X�_k�z����w��/8�L�A
_Uᛜ{~;�pVp=ѯLUo5; ��/���m��;_M:���tOq�- ��{����4x�q���K��<�]5,���<4��&�ưk��Ǭ����g�Ҷ��d�ӫ�>�۸��Ò+�Fl�������]�`��lw˰��fX�,��l��k��������蒶O���@��4�DS���jP}�i������I$��?�Q!T{KBD15AQEe�ELQ�2�"J��"j`�����&��*,�C���b���&��&��Y�54RRQ44�T9T���ՅST�AT�%U�!�"���Jb�����h2 ��a�
H�b(h�b�*�Zb
*a��
�
��
(
���((�!�f�����*������!����")*���j�L����+,��i(
B�����)& ij����'# ���30bhZH����
ȥ
N�;�n�� Oz��υ�-e�Y�h�J\2��c�}�!
K/�6e]���ܣj�=O�@8�Kӻ�-J��i#h+�{����ͯ�O;+�+�ٓ��F=%^}�1�7�U�=H��F���=�Y���ٓ�+�7�%D�s��C;�b��ٚ�iPhw6
$:����~�~_a�su0��� ���0�ç�Nw���#v�<`��Js(�F�������1[��z�h ��`v��ϗ�+��/}��׼y��z�������
�<�v}K/��6��-U}~�d�Un��VA��n}��ρ�!Sݺ�ӽ7���ȿ8���j�x�Y!~����U}�kG�nvǓqT�k��S�;g;�-n��v{&��߇v@L[j�zV������ˏ�*v��`����̶�#�xIc��6�C��,�<��[v���Wrc���3y׭��O�̗�C���0�n�]'y>E�C��`�ҧa:R���{:�*�GhY�>�R�~��f�vUv)&P4vڊ�b��s���˜��BovY� ���6�5�zo;��c[9��Rۭ3�+g��%�YZ)�X�����_;��,ʅ�u�Ƀ������z;<�}~�����n�k������y��DO��m��HWk-��^�WSּ&��&�k�l�q�Fl�����⟢! [!���cѢ7*��T8[zr�;yQɼ����7F��Lj_ghqh~�6�z�(�+�;I��-9g0�O�������,�H�p���ud�(X�_x:D~g�h�̼-��;��A}�ψ������[����dc�G�����!܁�]}5z�Ϥ�Acaw�׽��Bπ�R`o����W�nY֥&�����GЏmХ|�����G�����g�=�����O]�3^��~r
�'��6�y���|Lj��Ztl7�'��ed�����-�5�G���yA��� ��n��I�b{���	�^#����'�m�/�cӛ���\
NX`z���Z��$׽�ǲoU%]=Q�<Ȉ.����͙d�����qˤ�i���u%e[�7)��z/W�\����y�o=��x���7����8Nթ�];���w�iS��?;Ok��U�u!��њ�36]��6�\�n��;X�F�v�
�cx �_@<�Ei��N�u����N�-e�Lw/Y�<�qT�n�u�K�aX'����G5��ý���E�cox��!o6�������f1�v���\���w^{/�݂�i��st~C�ҧ�u`�x}ݣ���9�m�m�x����^y��^�G��}\��&T�c��c��&Su�'p�'qW�d%��ǻo�����S�9H��=�Bk��&s�DO��o��,������.}1�t�~�~i}Q�ۓ�|�,
w'7�'/1�a}$Po��s��/��go��ϟP���xߢU5�Ѳtm��}�p�c�s	�YKw�n�^��D����_���`/4�zD;F����5�U����-}u���g���ρREvį1���v���E���{9�A��2]�d����zoNUy��K�E-#`6D��ᬋ;��K����Q��Ŵ^w����\�k���-��~rB�S��s�:��ϱh���h��;��*�%7{�Į�^4�T�b@��k��:��B����i�'��+*��mkꌦ8,��RM�S�x0e���畺z͙g)����ҷ�yP�3���f5&67�-}�x�`޺�+y���{{M�k����t�i������ ��=����WL�8Q�ॏf��F���'�'W=��V���y�2n���۪`�r؞����5}���xo;w[R���yɄzh��Juqj���(���^��n��\}n/,�H�@Om���,ݿz�v�K�F��va�n;8҈�>�/��P�~~���y�ޢ������b�>�}o�mS^X�k��p�u�WU��l
/�pOw�
}ǰH��lzr\=D�+�^F�ŻY/����g�">�u1���k
z:�q��*v�����y�gs��T��
�ߏ����Ç���R5߲5�3�`��C:���¾�+�=�J�=>�!��<O��s���}�~%�u�v��'�|�m����XoJ�@֛�XZPp.�T:$r��UQ{5�}���ï���!"��M��-���퐌�7~�O՚��Jb�n.�]c�{qW>v��۶$Sm3�t�3�];����vm]wPA׀r� ���X�.t|'[����������0|� ��?X�h� \�v����5����7��Z�
�+= ��A��>:�1��=#�y�6I��ܙ]�$�^��o�;�� ���4�~����,��G������x��RCygV���\�HN]�m>�;>���ID_l����ŕ�7Ϯ�;؟e?9�97kK>�1�`A�$c&�g�t�5L�Uw�E�������kE ��9�x�?d,�yI�7�9(�D�h���I�Ylԁ�ӗ�} V~�(������<c�\�Ѻ�@o��Nn�(���^�h��~��%�n�E�v<�}�����|HRyaaD�2F�dw��4mc���}A��'����mk����3�W��z���hUy�l��Z�f<������ja�+򍪮�̞rᢥ��a��V��h�1x3&dxijﭸ��=۴���0�N�x��MJ�6U4�+�ë�n��O':�C�3�{�>j�c�U���ddޏ�\���mձ��0�UgA%���Q{�E���Wr�h�.Z�/|D��w��5��v{�?�������scQ��=���;&��RK�Y�Y�B�Oo{��&p�Po�'��e_r��V����=y����3~�<.�l�5�_i.}�+�o�xi���ҍ�����GM�OF~W>�^vUߞ6�Ԡ�T�f|���lx>�0�n�ˤ�'ʷ�:8-����2���{nkG_�/ �(Ϲ�c͢x�j�_5{w��U�r��MyУ�y�zcx���9�x>��P~���l��������S5k�>l��vr�����x�Ɣ=�p�k��~�%Xy���3ޫZi�����~�;^vB�wO���g�bJ�u�w�]y{ss������Ѽ@��<z�RYɕ�ݘ�g8-�����]��Z������{^��F"Ll6w�x��j}ڤ���;�� T����Vy$1c��[�tx��/�S�uq�us����D>$�7��~��4m�}��-�Op�
Q��-{������O�Z����{�z�&<��}����W��q��fm'������N�]s����-GiOm��m}��s�<u�z�����a}DeWJ������Y[���J��:�g���7b�O���0���=��i1���Ztl�x��x���aɗ�1d���o�}�{ц�uL�r؞���P��#��n��R���.�['T�=*w��2v�`{��;Z��ST�������1^�����=n�Vp}*��8��_�<��k�?&;���$y0�zFk�Y������m2x�I��ݝ�r��Q�
^ς΢7'��w�gE�myA1���K56vt�S�<��2�i����;|,xi"�Q
7.h��ݚ��:�ْ��c�G#܎:=ޝ\�y�1���,x>@��zMz�Qk��K&�+�v?d��NY��!5�AȌ��Q�}���]w$%��}]�J�ٞ�"T���˃��)����/lس�A��X߈z�¼R7�Z��ӱ&V�E*�|w�H�t�>���Fe~廷�NX�n��:���N�)=k,�F�C�X-�r-f���\9�Z���>H�cރ#�l�>��������7�X������W��J�>��=ѻ���r{�/����L�ɇpx{)�Wy~:;W4�d�?c�:o�*��ݣd�Ѽ1t���k-��~�z�l�cÂ���cY�ǤDu�搯H�h��]E����wۃ7��^���@�L�>G��bQcY�ϼ�����4������������zGt4��}�@\bJ"��ٜC��g|�{q��]o\�r�膳�.1�pH�[�6�����hk��#]Q<<�y�ez���Qks�ж�߶�3��E�X��H09(�蟎8���.�p�n̦����;<�( �7�'��fL�77S�T�&�������>�~��&0�;��c�Lx\�/x|H
NXX����o�2]u������T�#���������fa�w��VR��=�Ŝt<�*M�λ�˖�jS{���|d�y���e�ޢ��7�����x�c��XD������d꼒�gX<A<&��_X��[p���A���Yt�L5�%���	�ʳ\��mp����RL99���F�#7(��p]^	)d��r.�0�R�-9��IY"����>؛o^Y.(�Ĝ77��V;��G���W�]\�>���F�R��#8��T�6�E��m���;�z�RrdyE��
y�t����in��'{�����#�w��׋Í��_ͺ?.�}߲5�)��Jm��\����I�?w����s���2���nW}1�6���`]�|;�9`O�S�����wPc���C��W���
�Յ$��?mx�r$v�nl��Z��Yra�#���1������JhqiO�����,z4G/33i�S��&h���u�tZ{�<z�1��_�_y;o����/X	�靻��ݪ������݌�vm���9L�Ft��ĔE���S�4�|z��L�ٛ�;ò��_,\�����47����/��c�g�Os�iJJ�Wd���=��砢|=�Y�xs���D��)07��_w�W�o��X��OTDQWU�]���{�(%�h.Cy���q�����S<�oc��X��u.��b��+��;֐$����`I������0������=룅���A�}�I����5tƩc}ʻ���-�����ou8�ȩ���N�]�2��rN�瞭2~��Ћ��Ð����77S��ul���s��s���7w�	��ȼL�Lh�F��_��&{�n����U����>}@o�L/����E�������u�f�E70w��/�U%��*�:��spkRv�1�Sݻ�3�`��P^�wի�.�%����gKz;�֌��,��a���.lj\�*z>U}&N{&�}蓬�D�N�W��HE�o L^���}�+S��XQF�ݢT�J�����ؓ^+�n�%�1�C���7F7���g�^G�9�+�Z#���_���]{ ����|*M3>w�_��c����m�t���Y�X3_�����پ�Q{#8���ښ���r�h�s6<�'�G�1����₦ͪ�W�\�ʝ�T����`Sc��i�ߢ!����]�ܞy�[;g-^�>�XE�)y�^9��q\��<c�l5�9ç=��*��Q���3B�b���/&�:�9���|����*s%��̎���<�yբ���˧+u�c&�5����a��hl��uaX�wPJ�K��lZ/Z����Ыe�<�,ދ�u��!y��C�Y�l[�.�.,��i���N�e<A�o2yuDh��I�A����j9Sk@�/�&��,��G'�*/�s0�`�Ls;)�	?/&�˭��B�V�ܠ��ƭL��͉5p��gn��fx"b����O	T9�Aٿ�V*�6��!���캡�����Ō�ӣ����Un	%��<=�A2�.�'���5�8;�z\Ʒ�g�Fަ9}�`���_7����ͬ:G�oc����z�B�`�s*Þb�;����('$#B�5�I.�D�Ӿ��2���Bgs:�N��B���[�cC����U�Y
�TÂ�m	������r��J���o��7�ci՛���Jy�پp	�.��14�!�����Q�
���b����{R.�����-�(�˥]�z���/�n$�y�(wk�!��~Ό
x{k�| �����g��-����ɑ'��u��u/�\�嬱a�Ui�P�☼s/y#��2��No��y���C���Y2w���y#T�&k��lX+RX��)�3��!��:`�l��ed�����.��u�p k5���ܴ%�֣S&M��Ԗ� ���[�.B���<i�����}BtvWt`�L��X}��6wgw/J���wo�b�/�̆_6Ÿ9��Ge8��l�I��39Ӿ�wc�:ʨ�BhU�nM�%��*�U�@��|w���n��U_n�z����K�z���]-f�O%m�� ��c����0��-wB���'}8�#�:�>�7L�
��IO6����h 㫊��B'T���v%�$���<&�
��B�&��O�r+٥�Ι|�ܑ���׶2�׽AGiv/wuu�{�;�P��e^̞��u�J�g�F|�׵�+!�؄��SN>:����9���.#��o�X�8.A\?����2�,\�x�;��;�gYuj�e\n%�Y���]E��z����Ϯ�c
�ӽe����y���#VQ���9��=o���&9$�ʶKq[5J8kz��R��'\�����!�{2��.U�
����λ�E˽��8p_v���,��®��*���.�5v���c`�z��~��CXssD�b�y)�{���vct��݅��2��:X|�t����������9\���H�]W-�x��R�{��8,ǲI�aZ��=��F��}�fb��XYt �*�K��"�H_s�sw|:,7��OV��_E�I�`��}od��_W�a��;��qeOe�캲�|��%�>�]��4{}�3n� ������N�b�����VU�RD�5TM+��d!�R�SMRU%4U9��QCIAM#AMddR4�d%TT%P�Œ���ДP�TQTUTY	YRfdE4P3�Ĕ��T�Q+AME4��4�NK�L-3�IC�KT4�����Hd���9%AI�dTQ fc���f5D@�.I�fdH�(�f4d9P9!�KHR�D�&B�BY�DT�19!��R!�J-"Q�UB�1CFMQCANFFf5H�-�E�&IEP�%=���Ef/13k9��`�V�윜N^���n��t��|�*rӭ����ziTP(��V�\��X��ר��wJV������hm~KZ�5�ѲgF��cK�{�����c���ܾ����t��!ꁇ�ǽȇk�פ߻�'���4�b
�(�E�q�P�Bw���z�$h���E�y�����Ϸf<�;�'O��~+�Uev��= ��烬���ٌD��E��Þ9��Q3o*eS�:x�����i~xx@$��Z��Z²
'���Ik���z�r�n�{m����0�odsz���9洕Q�+N��o@dB��w�[��Ќ��3�{ч��;�'l/�ѳ8�=����ur�w��gg�q��3=��)�XXz�ɾ�'�)�k�������f彣�c�r s8^�<x�2���z�<<�R����C��m�M�Ϋ�I��I��y��5���Y�C�D����+I���w����
h��8�7ch�Wh�@-��(ߘpZwFu�W^��z�����x�9{���O
���Vva�:��&�l��pZ����ݐw��l�wm�3�y�:�����ŚJ�8Px���:F��ǫ���x���x�O��,қUǠ�&���Q��S��7\�"ǆ�c���"������&�Nv�O��x��t�}���8�`�4���Qs���������j�k�;΂��9�NX�',6�{}5��Es �Ig���Ozb�������OTg+��ۓ�]����8��������l��)X�8���y���r���h�0to]��䬯.��m�a>l{3��	�/���=%�������h��{�{ՉEn�|Z�]��JOL����O���ch��	P1����,��m�Ꞵ�ã������5���?8�Rв3��h�z3�y|V-�h��<�R�&��}n���m<w���Rc`��p_��h58�/�>��-�X�m�ã_���OC�/:v sٓ0��&;����G�~8��\N�\/4�f
�Y��ކLD���Ū�wx׈{u0�}�~�w]:�v�d\\W3Z��������r��wH�'S��p�?l���t#�a�N�X:��m�@��ܻ�nA�ؔ}S�yP�/�M���\��M-�x��3[]3e�=�y�����6�Ly���<ȿyL��?,2nn�v�$��ӡ*��:u�k��z�B�<`��K������Y��'�ĩ9,y{�t0�[�&�{G;��8��L�}>3�M{��Is�D0�~���Y{�|3;\���0M��Ґ�3;#j\��O=�8�sz� �xoŊ��h�����[��ꯝoA�ǃl��l
/�q}Sݯq����ƪ�1Bv�g�\�����0rQR5�Ǖ��k
z:�<�S���f���+Y�Ǵo1F������m�]������Jo;�;�{�[��*<�[��p�{�/���~��E�Ev��݅V�_�q^�^���VIX7]�{�}q}7����bIZ'�͏6�'���g�o�/yU�+��f�-�k�pL�/���!æ5���|G�}�0!C��mЀ�7��G���w���B��b�ܚ�GN���@�B8x�JZ&�Y�mz�ޮ�x��C�c������0�Z��;1Q6���H6V��u��P��4�&�g~+���n��J���u.��ѣ����c�ޅ��ny�xE��] �]��{�N��T��1��}�ϥ�����u�.0�0���ym{TK���|�tNY^�wO5ѝ#=q�(�϶ja��+���P8�C�*A_��9�2K?��اt`pM��B����%q��9�����Xߥ&@��`9��c�+��0_�s�E�U����e�U������7����<�V�#��7[�G6��F\�h_L���H����C�v���&3iמS���${~Œx;�K٦}7R��4��YG��T�ں��P��O��mS�ĩ��x�s7��xZ��/K���'���@�Ƶ&v�3�@_�mW{fM�9s��v܍��ݷ#�[�_���|���m�3�%���(�w�f�A�]�t�YsS�S����:#�;M�>@�+^|��}�j}�XR=T����Dp�1��n���t��۳.�w=Փ����vh��K4�Z� �wE<*S�0s��t�n�������.���o�o����Ź�Q���nы
��t�����os��u�{s���q�i��"�=�f�ہ���;8Z���賧�%�Ty��7�7X�k��&��8"��vb���Z���*I����1'��}O���L"۪��m���6���;GgL؋[	B=������r��}���bWط6�����}5���Tmܝ<&7�؃��r�~��o����6�oC��\����F�/D�5��Fɝ�<=�p�gnr�|rPyx�OL��W��ĸ:���ǽy��p���u`4.���5�bfz��IY��/|
DP,J,l Y��>�+;��z���ۭZ�8u$�/9٢�c����zd��f1*���9���I��Uf��v���$��I��(1�x�e�8|5�d>xy�d���,�T����{��O����x��L>oW��8<֒��?N�X�䟵pZ��ۋ)f���;YY��lҒ�^)u讗e"���+2%�Y�Z��H�tq���Ơ�	�!tzL�hvY���n�Z
-�;|�Y]<2�٧��9�������ō5��/K�C��7h>�x��B���<u��b��o'Pzp�i�p���D��F���KyΨ':�m��.����<��x;uLN�_��3�'��.���8�������;��Z��!I�aa�>R`�jdSd]��������ܗ��l��7����.�rx=}G,	�v�����v:T	bA^�'{]�� -�Sݻ��/ ��~C���7�½��gy�����m���l�������(���\~�NӸ9�!�Q�W�5����+�Y[�*8����{�1�ّ���zuw|y�3��1�aF���w�Oz9~~;g��oh�#C���Jr��o�MxT�\ίr��o)O�n�����ʂ}�����l��÷',;�ϔ�@I�{�iU�\�J�HJ�Y���^LÆ��9'�����/�*��Fɳ�J#'e�}�O��U���c�6}���y<C���5���#��搯H!�߃����zmW�~��Cc�B7�#B����d^���������.�w��PP������P����#��Y�d���W67�-3����
˲��Y[8j"${�9���G^<�t=S�77������h@n�\-9��N���XA�mǘ��{��q�3�	��o�Y�*8�ؔǟ>��!�<���)�^�r��H��<�FvH	q���,��"pi�
�BW���^G��y��S�!��P��#b�����5↰o�){ol���uo#1�U)g���Z��c��"�g��$J�{����Dv�=��@����`�,�|=+0�>��=�MϷS>�j�V��'��Ϋ�ڠ~�^�����ƫ���Ȟ |����
�YJ��{tخ����(go�_o�������T��ax��Y�&��=Bu����Z�f4;F[qƦ"<�}󍗟M�!�8k���V�s�-�M�����fT��Ͳ��E#���~��{���7��iw��ι���g��Íxs���\cK��C��'I�w~pkJ�����)��IÎ���*,υ�Yb��=�}2{=���/B�Z��L�/o���["���*�����;eQA��=K*��۲/f����k"�.�Z��l��M�2���θƜ��Cs�=�
�蓵�gm3R'��})���o����F�<4�b������4b���)�7{�����cF9��o�EYF	��}'�s��v�wr������˂��9���dH�n�T~�xϗH�sm�7��mXBIF}·������[+}U��5Rk�gK�k͓�LoL�/���H��D1�����kT�=~#I�۫�Nl���R�����1�cHB�0K>t�)�Sar�*��kϝ�Rw�n��o�{ֻ!zE�9<���#H\b/���ث2;r�1�촺i�4�W+�����әC� s�d�@Z�C�d�t`A�+�m��N͛�jV��\�ѹ>�|T`�b�8y�9&���"eg���{L�{��f��ӡ�S�蟎��+�*�/ZYʳ}��c��gr�<K\���lZNG��0�{8���4��yDN�O�${��gt�ߒDٔ�n'��Hw��l\�^�������w9����wB)����΂񨺥e���uh*tO���	8y]��4����{�p�ȇ͖&�b"��.싦���(��ő��E�5�3�!��mz-�"rV��1Y̹f�0V*Wt�B.��y�iGݸ�T���ٿl��<����}~�	�	㯐q<ݽ�Y�
�j�f���z�Ng�澒�<|7�Ç�߂;I��:���η5��<ru��9c�{�hyÝk�`��s
�eg��������}� "�-m���Ng�u*x=mug�FPy�~s>َ�/�(ԫ��׋;�,{��>ըoa�n�]�@F����m��Q��'���w�X:r�U�Ks_u�P�����v��R7^=oӵz�(i�ι�*���/��h�#hZ"t%��*�o���u��;z���.���}O>���6������GJ��D��w���HUVz���穴�����9��2����3�qzL�gM��5�+��E���Z��[�=�8�iz^EF.���#�t=>'�o��/���X;�1���n���x���vg��ز�Wd_	�z��Ι�#�߭ n��`F�X^2�B�ۥ�ˎS���(�>��.Z�ۣ63՚9H��HP>����c��B�/���{@H�(Է�*����3�R� 9C��ل[ש��.�:�fx�\VG^�%�D�P5�VAjĕ9뷉L�4�ҝ�n��mjv����͹����՞���}������r�l�Q�l�z�7j[�{se]��o��T�e�5/6w���ME�7����-�ѻZ����s�4�v^ot� dV�1ЯKZ~f��Ң|��|�S_4m?��k�eOObsz��%N�zp�,�w��kj�����(M��dF���ڕg��5���m��s`��}������!(��dw��eA�3°�s9��1J�>�X.���:큳q/m�R|��9�L�B{����+t���u����4��m����em��<�{ಌ�� w�V���Y���z�hY�RY���8m�#�<e|��'Y.Hz�L��j���.��aak�nR�/���@�v��<��,�X���R.���þ��T��k_O�:��a��-��u��VvT�Χ���VJ�V�8�E��*��������\�.=�f���Fרa�J˄v�׃m5o�ruh`hr���Z��WOÊ�<���Im�@_��n�KIz��ܡ�}���a��	OLߕ�����qPPzt�����U�o))��n��w��<�@�ˏ0
|�=L����i>ޫύ���_�TA_�Q�ED��D�aWB* ��Q�
�+�B* ��Q�D��W�TA_�"�
�"�
���+ڂ�
�1W������ED�H* ��Q���+�ED���e5�K~PfEE� ?�s2}p$��<�H�E*�(U*�H�P"���"BT*��I!"	��$�T�P�"@"!EQU
�R�URP�U(R
�
�"�ETTJ�@�A�tB*��ֈ�* ��ѭ���J�U
���XCc)%	���II%R�X��R%P"�:�P����D�R��R�IkJ�Q*N����BU��EB�����!T�u�B(�IJ�*�̔�HIG^  �����v��8k�(���[�̦��
H�ݹΖSwl���wT7Zf����Z�wP�t�[���2�܂�VۥsV��VZ���R�
��(6e)%�   �y���:t��K��-ָ᫥hj����p�kv�����ݍ9	��GC�Cuեn��G[���9m�]�Ȯ�VuN�km��ú��n�֪��HDUkI*ETW�  1�ڗ�m���]�Zkk���V��۬jݷK�ڙ\�8��͌�u;��]�V���.gM�{!@�L:
(P�B����(P�B�@z;�
(P�B��R@��P�B�U=�  1�(P
 �
 �B�
1��
(P (f�
;aJ=�zC�º֝��n����T��Uvٵ�kf����@ꨪ�,7m�Ӌ���
J)"Du��  n�EU�i�U���v� .��`�ֺwC,����Ԡ\�sBڵX�n����r��5l�v�-�Ҩ�(�)�%$�]<   ]�]t
ږ:�GL鶶�wg3ڋb��5�j�73����heUmr��*�����m��6UR��-�$T�EJ�  gU�e��B���k�����vѧ:�u)N8eS�����#`�u��9�:̖�uv���jni�N�B����F*�%T� �<  <��zݭ�j5�U��5�U\:�p5���-kv��M��m�����t-�����pշV��m��wVn���V���˴�e۪�ڳ����R�J%R��K�  ��][��[��.���m�5���r�A���1Y�J�YsU�s]�3uۻ�f�K�U��]�m�7u��[m��+�ݙ�6��5�+w�
�@J R�L��  ���r��N�Gv-b]�m�ºն�wsu:��͔�M�v��P�\�]�l�cZ\�][V�m1��*��ڊ���յ�f�gS�\M�v�x���T��h  Oh�JR�  ��xP=@ �J� ��� j��M�R��   �I6U%dFčDE��N00�-�� ��1E$�P	U��}�S�?���~v���r�?���$��%�XB�r�HH�	!I�HB��@�$�� ׇ��T�_�?gu-����SW�8
�n�1�͸�,�(2bV�4i�T�E���4��2-O��b��M	�T�ۤ�nV�_+�,�$��ܑ�2��lO(�ȕܖ�6�=g5/Mn�Y#lCW́�k/_�D1���l�N�����,]@%�r�Bt&CKۡi݊�B�4XBU�Ym�&B��,T�b;�y{.٢��_�bG&0� ����E����G�4��!z#:�[�������Q�G�k��%jC%�QY1g�P��D�ͻ�5>ݦ��Ϧֺ�H����b+6*ި��>�t��]K��^�)�X���Z�gC��x�DQAhǮ��5���,{��1�B����od�L9��-d'L*�hdI[����a-(MMlu�A�/	��U�u����
�d��kUG&�W���{�Kq��f��&%A�%�J��w�o�u=�N�+[�����e��4ւ�[�Զ�������K7�ct�DYɍb��t�)�3	ʍAn��>T�]�j��t���ۋBoM�]@$wQ��a5�0��lS�� IM,��b�b�OJ��iM��[N��1�eh֘Ķ�sn��Tv&UtG�mLƬ�����`ܚ� r��NӲ�Rv%��C��)��L�nʕ�]̫��o4BrQ��1jkG�e�[%�nL��-� ȍ-$�7	�k1лW���YF���C[t/���-���1�4*�K��F�,�p��ۆ�K��@� �G2�Ľi�S/#h]5Kvd��kXT"^�v(*acW��� �m=�P��jآ�ea��c���"
���@��Pbƶ�e
u��4���+�]�b�RԏRݫ�����8��4���k���dP�[��<��q��Vg%��%�wJ)�*�^m�$��ʹX�J��l,ܗ1-#�A2����J6N��C�`�1˭D��g.lIn��M�iȕ��44lm{L�x���M`Bڸ����MS+m�֣�p�"� ̎<��ƛ������4B7���	��f��Emփ6IZ[\k��ݳ���5Չ8�X�3(��B�R�$�5���Q5Kk^���)��pD��3/r���;�j��0��8^��=�n�ph���of�QP��[Y!���U�5
�!����eboA�*-�z֝nl2����K"�fhu5(j��tt� �3�ǗV���Ҩ�{1f�̫��7(C�b2�3/*;��,�5^������*�]��M�Yb]�V���IGHu��QZX�1��h�"ৈ�U��,�Ֆ���7TC`�0�h����Pu���V��	h�#w������6c�Ќ�j��;VA{e�5���Cnl������v��";�$�H3Hڰ�n�%��iʉf˶�4[�h�B{.���A�n(��K)�W���u�d;	��u���"ڼ݆Ւ�mXwQ��u��:�B��n	2Q�ٵ�a�YEїK(#,+���M}r�`זȕ0SuwN�0\ї�r=CY�B�eL5�ěup�Y��X֗��`\0-f�Aˍ��u�Z(}(n����J������\�F�'�=;,m�����Էq����n8�ͼ���t�&�R�N]ح9�KA���@VbZN�!���4d@+ki�cl]97[�+�J:W��L���;�R^J�B��ݢ���p�T���,���d�"��p��ˍ�r񌵕-���^\�9��A���*Ouk�Yvl8㳮�\��w�ر���!,����R�lZ��+4���
�#u�H���p�G�-�����WGq݆ii̲Yt#���D����V����ܽ+r+W��N��a���NMC�d�.�4*�mf�$T�e���Nm�kn��3-ٗ�n�T�aZ&=Ks �m&�ڒ�t�3yR��)1z-G��IZv�&񋥻,f*�K��Yuj֑N]]\w�LBn��e�'��ݠ�o\d�\�VHk(�2u[��U����`�r�-��j1�A�zKԴc�U�PY2REUݜvn�
V��-1Z��w�U�:5�Sw{5X{����B�p�&�٭"SF��w��Ă7-j��S~Q7E�����7J��2Y�``�[�S���l���U^@�*�ęZG��Z�ܔ��$�y��%��e��m+��X���j�����;��
�R\R��`S�AM�{�]e�dj�ô��"�XB����.�nʔ���̩�YCFn9 P�R6u��!�%L,�D�n]^E�uw��+i�PdH���kdh��wR�c��Q�u�Iyv��B�ӭ�-�
�_���Ò�S4��{����E�
e�ľvvSQk#�����܌��@�
��5Q�l�ɷW�i�檇/E�@k�ڣ��<�xT�P-�)lBf�{S^��k�)I�Yr����[��Z��%����G��@���=�2��1Ñ\K
VZX�(*"�4F�
�@SE�AO�)P�Ȩ��>�m�y��P,���_l*ڼ���i���x�]�M���X1�!lt��ml�&��I={��������1��E��J��-��H�v�Hth��x�����b�@R�tr����%e���_]Р4�$���m30<[����4ZC*��ۑ`w�7S)�g@w*�l���ɹ%7dH��$�Tjєc7Ke��h��
�*N��7%jKmj�HH�q��ni,J�
�ZLU��hS���j���H��v u�e���%l�0�@��#�d���S����r��k�����-�a�N�c`fVSnֺ��Ӻh}���2��X˥ou�Q@�nU��Ҧ ���g*W��:�� 0�Ye԰L�m�v�l�N�Gfae�-/��^(r_��zN�)]Jm��%H�m9��ƃZk+�Ygn3V�SW� �n�;�EԓL�XP���kȡ�vZ5�0�Y՚��;H�(�@�g1�е"",7�G6�i]�,(7e�ۚ4%��W���+��&-��6��H2��!U���-ch<ׂ�BS����呎��Գ��nCS&,�n�j(*��TtDyi4j��W�-�6�c9���N{�B��:UAup����rmnn��M^[!�eF��6�Yp]n*�1e�)�M,H�c��05��VWx�Ҷ�p-�BUG.C��!Y���p��iw��_
��
��[5��[�ȕ�A�b̈E'�vefe�R��7EF7h�Q��
h�����y��*amR����0@p�+QZ�XN�qh�s����˫HZ�WD��B��J��$dko6���Z�Z@��YP���fj���
?n��ԁ��b5y�큚��9Y0�B��se,b�`՛��l�W��ri2Yle�0i��m�#�ܱ+�S[t�ח��.�v^cYY���0h�� Y9���2۹�X�e4\�R�Q@��ec�cT5d[n,����V���N��IT�2b�v�*�Y0H컘�U>�t�m��qT�fS����xH�e�R�*�������E:�3d��t	
�ܕ�E0ܩk!�-a�%Zt��ucI�N�'c:^)��t�XhND��/d�8��Dڼ�V1��U�Uј���^4�hiEw�V��8��j($�@l�[�"�Җ��A��Q�"
�W[�n]��uf!��kmv���h�X�ӽ������/!F��&�N!,���!�z����G/\7��U�P2���c ��
{�7u6�4U�w
��+b���GZժ����^��c
��n��u�j&i�b�}�	�oS��\�v��	Yw��7v:�61L�e*�p�0��x]�(��B�����\�*��l�fC@;%�q�JpR�.Y2^�zЎ�5����@L �)�n���팢����P4p[�+](WٚlU�N���
ܴ4�q���g���j�Ei����/)eC�q^`x�"]�5
n�@Fj�F�%h�N��Ҥ�{n�D;��SMtr��m�LM̀,��j�zpV�KYSh&�6T7 �-��4��Cf�j4Ua3mz�ɢ�2�MZԱ[�7��Q�B�0��D��(}d�bEWi�0���L ��#���V��bd�v��jJ�Qe�:�&nA�i'R���[�̥�U���m �,��f�4΁>���'
�+UE�*UhvH�������w�ʇ�#�{�b�p�&��m�pѺT�5�5��T�l��)57PkI��Z���(��&�,�/Hf�&�-f�pAr \�ok�1`�9���Lc�֜V-'�E
���D�E)Rʢ򵗗���봸�ٴ�=YYX��nil[h:�ܼ���J�$�MFh��g��qb�f}2�����!R"���B��e��5�n��P������MM�0�6h�j:n��V��5 n6tl�v���%K���5��]n���MВ�*֖5�F��Q�ݭw�f�۫��E�ø��0�ql� b?�jQ���n�"2�µ��G2`T��B��.����C�$n�ǆ�Ӗ������͎��Ʉx5�ޖ�d �ܶ�0Ɲ��P�V���$7����1SLȐ���-4=�.�:]�Ɣm�.������Gd)�
i;�1cJ�Y��{t�锒sl�J�A��ܤ�'>m��K�M]��Q��6l�d���[[cD��8�Y"xF���#& *�D���w�=ːͅ�	{bV4��4��+-�{$$�Պ� �AB���d��G0�pU픑�SZ�e��D�x>��-MHi��T�{��]����&��H�9+t��n��U��7�Pq�C0�Hs4��&��pkJ����U�Q�/m�eKB*����u)U���Y�l�%@h����ӥۣt�m�ā����h�����6ѼU��Q�ImlqT.��X��O^֗���f���-?	�n�|ս*ݼ��F;ׁ����h޽Vĕ�q�ZܷP����ۺȑ����x�Vغ�qZ��%�x��-�r�J�&Џ*cQV��]lqfb���2��U�C�W��.�P�j����[��g;��fmXX&�K-n-����ue��1(&Z�r�2@�iT���t�;q=�m��`ݺ�yhPW[:�N��i����C���U�Z������!1Z��C&���n��K�YvP�a�w��̬{z���� ��H8��$��َ������}s�˻=�Q��n�J��ͻ�t(���7^M-�Zww-�K���f[���B*��ma����`;�@kݤ�I��n�0Tu��C���z����Kؤ��x�
s*�f��jMB�Q�"& ���j��4MlYmP�Z�c-#����n�l�tX؊ѥ�*� ���jm����(P#	��f��ИJ���2�fFC)�Gg@�mL�l�ۙFR�cI3��R���J�aӷ�#�,�{���,!�M�A97VE�0�ȕ'�uz�#�"7��QfЬ`?�'K��t6�5+I� �Z��ˤ�"(��$6t�.9�)�o2�3b�&!KY��՝7j)r],Y4�����)TP�u�5d����R[��ō�N]]��pL
CE��q�&k ݔ���6,">��X���2B֗b�qy ��*����͡J-�,垾��9ҜØ�;P�x�U�:�1����䩤����e��d�ek?x��R��vm�˛�W�.�e�l]I�ExDe��2�6\xr�Z�n�QnQ�f]!VX��q0�O b�[:7dP�G/[u��ʥfe0
8v�h�iϋvkYt�[������F�6^�v�t�\��' Q!��2�aZ��N��3x5J���OR0k͖��D'�ب���b<��E��5�v!�!GkUe�wZmەb��QRRwx�ee��� eҳlA�����]Z���bv4��NMki9[�,�Y��cÆ�XDvN:y��ly��XUz[���L�F��yp�JX�)��.�*�b�n)P��M#v��l
]6�bʷFn�����j?��Uթ*dA�CL�$L�U� �"�ϴDLZ��+m8)�T飉7r�TGbX�����,�-��B�,�x�뭑*�k�R�f,*��:�e�RbUg.�T�ͬ���V*�v&�۽��ӈ�UR*�QY��Eŕ�7/�ڱKQ�X�[X.�cjXPU
˃��=�����T6A�m@%Ժ��]&�6:�hQT�X�Q��F�.��̇J�������Rӛt[K.�K� ��A���۬���Yw.��U��F��� �vIփ�V�9dj�J�������Fnf$�� $�ZVh��Tq��7o*��Vh�!$�l	�Um^����hK� t���N�:���
��ѡ4�{�D�٫wz��d���,�BV�e�t�^ ��Y�ҥi����VdI2%�,��HoS&�U!.��f(�3��)XW�!HIe�$�;��N���*cp]�6�D�d*Q�����g*å�3B!��+�Z���i,!ദ�?c;�B`O���+�V��(Ғ:�i"Q�`�gi�&�9S:2-Y��$�q
�I[2\d�Eeg�յ�*%Jܺ��<ܹ(��ePSԱ:)3���mD�E'�IlR4�D���7�y�"�CVj���m�Y��۲�T1]f���������R�SCf;L���ݢ#6�2A��Y@��V"���I;ۏB�u	Z��rc����*��V�f�{��ܥ��d2uu� �Nh+1%�J�ɗ�f!*S����W���D묳22�+[o"��$�6*fi�Ȝt�K�I�{�V3��2��
p6�vaEbMo����ޥ��B(�ä��]]�gI˟-�1��)N���}�����m1{xG9�;��b�_�����'�K�`�oK�k�ugH]�_T����\��nwupI�wu�Y����vqh��U��}����Wh*/��`]\^\�����7x��u2��n�u�&\Ifl��x�F��m��d�F���%)����u�ye$*��F��a��e�Lv\.��삺� M��p;9��k�����t�;���˥{��J�e5����M�M�x�8�����չ��"��ƈ`���������31A�S�(ws�֩�{GYk嗘�s�%r���g�Âö�!;�{�l��8�'�`�/c����|4m7�;�Wz	���\��"�rv�j�	so.�q��nd�!���D+{���u���S�c���q�%�#�yŌҺ�eU�a�;�ۿJ��ӯF1/�[�i���8(��k���9`��}$<�r"���9���]W��n賙9P�䂐a�t�[O�v�I�N��Vr��gE�Bw[�iZ&���Ǐ(�N�sC�9�������2�ӓ=�w��c$8MvWwfh�Th�t����fWa���b܈г�&8ѮozƁ0���9��~Mn�W]z��Kgl�KY�f�C��b�g>���㥣]�<Y��.M���Z�)]7ݯ;i��MIe���ܫ���)�m��{6.����b����{N�����h�o��JƩvl-�8㨷N�B��?+��ۦ���y��0uG{�Q_hL)xs�u/v�����ܨ�����u��|,��]YnPˣ':���f���.��CX���ICs��ԍ&s��!³�D*�N7�RvoG4T�w
�8vWR@NQ�-]�&�t�Q��h́��,�:&vN0�u�dЭ�c���wUu2���D�a��LY�'����յyC�u#G{�9�i�Qeв�eD��A��ɒ�fu�l]XP��U��Ek�&|e=w�U�RǦ��Lu#�ϊr�sP4�o��C����`d=2�Me���RLxh�b�5U���)Gs�֐Iį{qR��I���TZ�T{�p�31[�7�Ú"�O&EM�g\ဍ�2Vb���2�P��u�f��ˇ��+`cbO��2n�7��6L�1�y��J���rK�^5M�m�2n�H�<Ux0]>�2J�ӵQ��
��6^C��Cs�6&,��5	3|�i>k0� ����6ouE��;��F�+:+�<u]��D�wj7��K�NѸ$d�xN�PG���n�{IQg ͑��s6��ڨet��zWZ�����FƮM�H�b�����D왝=l;�2p�-�A�{m�̮����'VsC�l�|35m��c�AS�x��֩%t�I/�Kl�S��+�s�x��S�R#9m)�v��,�	!���a�#7wݦ�_.��:Xs(R�ӑᆓ�C��n�j��L9j5cE�0S%.���<Wل�\ЫNHy���_:�̳��[{N��)2��ټ�@�q*u��:jT�h�2��쵌%������h��i��!�uc�q�r���͕�w�Ż1�l��CGi�#`�;�	7-�dX[o�9[ܩw�*b��!:۰��)p�O(TQu�
���MSZ��
j�>i_YP$)��Uѓ^AlZ�,b��v������-� kq[�[W�ZQ�:�;'*{rT�KxKA>�uw�h���Ɨ ��� ˹�e�Bv=P=��6r۫�9���}�ܙ�s_i��+���e�K�sgam�(ԩ:��ԣ�^��ͭ���'���p���<��vc���=8��{vu��}��oe�3�(|ѤLOue�l�A��UXׅs���rJ܁W �����]�u��y�W�[ä�k\z�E��v�Œ��j��˨-���+��P��e�#��㴌���ۭi�΃�l��ff���M3r��n�RGBK���]\�i�`R�l�cm��x+������+qԜ�ɞ�bV+��u��v�j'�@L��)*�/;�Rʱ�p��U�(����s8o���c�vWi�i<��-�'*j�H�٨��t�F�hx��t
��l��U�`T�Ds_s/�XСy�5b*gY�f���&��j���Nb�@����I]_8��(�8�+�[:�����'B�����C�@8�
��X��V���Q�l(�|���Lx�����4t��x�-ʕ���,�i����n<l�V�ܺ�{FQR���t̷�OU�wKz���-�8�т�+�۬ް��c7L(�U�mf%%2�50�tᖥ����c���9�]�<�:�en�`
k5�F[Τ�Ӧ`����{�+Z������#����A�\�t��6;�ǎ��EK�[J����"�%���[��>r����Fn����z����z����a�Ʋ������n8�n�J)+ַ?�����7e۫{�WS��=!����^�����Y�W��Y�ܐ�)��T7]B���n,��a/�wPR��C`u�:�ɯ(��:s티�]��ft�σ9'WX4�U�w.�d�����4H�c]�.V�$Nw.�����D���+1wvD�gn�/A�BL������%+�Hxu�>�@R�)�Yq��{��2&f.��p`��xtwSx\�8�<�yJsb�Q]a����8�+�Uą�;u��WǦ�#���K�%ǫ�\�xaU�lX��=�� ]	�j�����o���� '9I1���l� �>�Fu�$����o\��$�A�,����o��J�3^浡����H�4,Oa ���LS���'��[��&:��q2��:��Rm5O8v�,�}N�.�٨�Vsxɫ��>WӦ}��0f@1\�u�uIL*u`
G"�1ÁVfwhg��O3k�mt(��%�#֪�r�Lgs˫�AY�`���b��<b�j!��,J�sE�#�M6��w9�:�6�˸��	[�c r�C%�ۈ Е2��2�7t�g�X�n�jM��I��|�^��)W����e�B����ƀX �1q��z;,��ݑҠ���˹Q�B�������}��c4�N�T�Mm��ծ��}��-����m�{k����&�Z�{�r���ӖWu��޾�L���*��~g���s]D�\�.]r|e���R�w�}&q��y�j=�իP�vN��՛��]+]Yg(;}4��L��U{9DoW5^�N�Z���6@�c5yOS���Y�[N�|d������J9Ҝ<z�3s��G�Q]��.D�db{u(�]��A	����1Ar�ݗS���d���մ���+����-u�w��E���[Ԉ�hU���Gb�{��.�	��a�[���WA�k�`ӳ,[�du;����p�Ց�t���]ee77�N3z�]�n���zv�
��cx����}���%u�6�hU�ݞ [��CCāpՈ0�/nL:&�)�w�\�e��X�Fv�(i
^ f14-=+��9o@���)Q�-ErW�f��M��q��u��J�7�wкJ)]V
���AΉ0k����K!;��ձ����(�D����g�g�w͎�|�1��M"gg3]+��U�:8���d=*!�u;�<w���f�sg�eK&����+��׻ejB��HR��@�<	\�eC�P��J���d��6���/2���=lw��]F�5��?aj������09����Q���hN�6�}%J�{�3 �;K[@w\�cK�te��z��{J�6Mыu�q(l-9=Q��Y7.���*���ˢ͚;v��n����@׷$;��Z��p͌P5�9w,��S7nn�sqj�N��x��An��}��+Λ��g������̤�]��@�R��Q�.1��m�`�g�.9�Li�i+n�郰�<��'Vں��L�6�b;p�@�;F����K�E�A��f����!A�ےvt�5�6�]����Sڰ�6�5n��,�����Sh��c2��
���q(�	�Y�=�SXhRG�t) ۘ:�mN��V��T�ˁ��6��c�v�#���A�pG���EV�ԝ�zޠ0}7I�pW��/�)��+3K<b�h���4�2�CHJ��V�*��;Q�#��g)�W[�(�Z����l�rA�����j[��`c��E>����D%G��g6V��j\=��nN���+�h��>b��l^��uu*���"U���&�x�)�`��Ng݄ôա͉:� 2�vf_Z:ᕙ{s�a�i.�7�_�k-O]��<G��N�_c�=��d�}K��6]�w塡38�)h�M��ܧ5��v��-r�J�.��w�tB��y��!G����WlW��\��z�6tK<b
����+���g����n���:�㳙�:�ːg+})<xIQj
��T���V���t%
F�Q�&VNx���W�t��{�r>��C��w���-�!v�co1�����^Y�3`��|��T�K�)��]\퉹�,�c����l�o��ō<tR��/b蘎f���o�\j�N��H�}���&L��,��&�R�b�Cdy8k�s1A�N�Ѽ��o��c�먻�2�;-��pך+����T9Vl�#ɤT��;�I���y�]�5(�bl�I�.���'��ѐ%�G��'���Au�&6R��K�N[��T)�p���sd��}inS���-���*�[9�)uvv�[ѯ##a�n�n=]�Ya�;�n[L2�0���]�]�\뫠9K6�
n_[�Ta���wou���2빕4YsW|	�Z�:���g-Z/�eZ��>�����n*�=��/��vF;����*�N{u�#k���C&hce_vCgK3[����;u�#�.Yw+�(�t�t�b���<%j6��\@�\���Dq*/�Ҏ��j���F��Z�����7Z��/`A�ŕl�gl�\�%��wGwH�Y�Y�u�wTN��,�;�J�mu�$�L�A��9��wo-�E�r7z��hḶ��F�S��ޱ�s���8լ:��	����U�7"�݌=*opM?�#μo�����ZW��k|�@S�/W6�|�c������#�&+p��T�^����I.be�*�g_h5szx�{]$�VhEϝ�<��)���c��t�j Ie8n�I%}[��������JªN�ѿ4�z�ث�;�����h�O[<�c���� ��ҩ��\����O�X��ȥ�:CC�,5܈���n��7���5�:M	�o�X��m������zZ���^��%7\9ǥ��/Wp��t�,��ŒJ��Dn�Ec uX}h�����u�eu��G%
���ArJ�k�]��j�ų�F��썊pD���,����aψ�6ռ�|5��e�εF$�U�"E�C�J+�[����X1p��N�P}_��r���g\���"%ѵ�R�jR��vWj�_Vn�D4ƻ�R�p�Y�x2��.!R}c�%̳lG"�y�L��
���٦�-W�nA�z�(b�h�cn�.�˂hnӫƤ�b�-5�V���5�
�!њ�����r�;��SքA��V�:�7e�ݼ��F��#d]MZ�B���K2�:�1���wi��g���fZ�I���|��M*�������v�g �њB4��v/ �2p���L�Y(�+&b܇��yp�ݦTnl��m�#j�mr�j>���N����qx� I�Ow�1�S�Eҭ�{9�\E�u�QJ]�5k��i�T���¤w]�/ #h�Ct�r���B�>bh���{4���s�Y\i��m�D���ĮE�K^j;@o<�Ο;PȆ�y)Y[�5�W2iF��OsR�����/ho�ul����$J#�	X��@'����B�r����)��%�m^�+���{����k��b�i�ô�)�z��S�,�FV��� ���}�����9�f�.{�<iۻ�f���])��sX�_L�j�9μ��إ�$�;r�U��<���,�WN�I��TI�v�T����sp�+�}��b%h�c�
��g`���gc`B�9�cŵ�t�:� g����/4���@ayͲz�4����Ŕi^Aw��ӇPǽǖ>�C�O�
�S�tn�4,�Y�x^Kq���+��<�1QY�_vd"�-���[�n��r�;��JeJvXf��O8̕��Y#����OF9;��y���t�r�h4G%ޓ;�ĺ�f=��]e%*�ft3�^�i-8)��ls�r�hu���!⧕2�$K��0Wa�d�Ɂ���1ճ�a�4;M��#�u�$k�[�����|r�֥���%R%�'�K.����U�)"�x��vQ�E*�s-�p>
�ɌgZ����e�l�$���^�*��c0>3�v�jY���O�PT6�\���;e�H.�mwhj��SX��[�P��ۡ��K���a��O vm��+�����ܩ�`�b�gAҙt����V�%��윞�;8���0d[+�ŬJ���InYY������)����iݳ�O�V�)�=y�WZjoR�hvX���w�F�Y\J�i�s��#�ͺ'gn���%�ّ�8��	��[���A��7�i�=�k(s���C��Ž�qT8�YWA�ݑ��YpN�;Cw���T��dm^W_clt�X�5t�j9���y��=ʍ��#e�4�uN��[r��z�U��WzY��|7M8g=�M3��wEn�N��Es��2���;y�-�p�t��r;^7i9�vW7C�F�.��/J._>��w�.�]1�}8x���5����x�ht���ϵRZWl`����sc�E>U��G��P&�]�m^��W/�� {����=��x���\�G����ˊ�9�썪�5����L�ƧŷIk�T;��7�s�+Y�b�*�%5�7W%t��Y��C�1$�x��g�"an��r��
B[�Bk;g��>��q�^;Go:��R&��i6Nij�J�s����[���CO����P>�k���=X$�;��E���ջ:�F�v0���U�l��OQ��(!�T���H�"�q/,�ܫ4�{3xZ�}�o�JV�:Gv�u��n�U
�}�F�i����4����q����b�
c���bsSZ��/f��6����� �Ğ�$�Y�F�b]�m*Kr�ô_<���4!�IQ5w��h�NLzۆ��ʂEX,���؈sE"[g3)܋q���Nb�)�*�]���9�7CY۝L^����.�+>�#���'�,����W�Dz�,�׽�n$� �v��V��42 �K��	�v�R��4�D�{�yS�:�+o��H�vw��hV�ќ���7Ro�<��p݈f�bmfl��N[\���̍ܺ!W��ꅱ�։����{/*�����:S�E��J�7��^.+%�	�	7�-f�t�����7�+�Z�V�u�zI�Y �9t�t�V�]7e���2�6;�L�H����/�]}2!؜�]âbvM"P�7�w�gt�%d�Z�Q�ʒ��70&	-�42�:��W�h��YG�O���d[��5]h̶6�t�q::,p ��Fr�L��uD�S��-[Me����ve:��먪A)����]"�>޲��6Z���p�;*��,R�R���ڡd��8���J�;��e�to���^Y�#�Ňc��S�$η��t���x���K��ΏѰF���J�������|��%]$I�(��UceWF/)E�ӧ��PbCzWM��cq�,�Z�N�pAW����|����MI"{ip�y��"�mv�0ʝ3h�����'GH��dZy�����k-n���'!h�u�Ѭ�{\�A�Ԏ��]W�L���m�� et���#��}i@�9��7��{_��f���i����&(��Vd��T��Vb��w�ս�����a֖�yN��6�l[>l�oQ��/���H�]��x�^���Е�BC���j=+*�F�WFl��wp �����ҷ�E�̔4{oK�-5v&�7W�b���9w���>oq��լ�6��ʀ��o(��҆i�Hm�d��m��$r��Y�$�[�Ԏ�i��i'�
�B�\t�����㾣�)j�+�B�H'�����9��=�]dT��t釩����Roe���7h_�ڗ)��i:�'��Qkf_1�)�ԯ��x�A
���Zہ�٦�>φ��:Q�z3Ep�w�G �`ۜR#�_�w/�,aY��0�蜧��Z�*��H�X��̡��0�μ�,��#�u��N&��
�ٸn,�U�]�rY��֦e0ƚu��j�o]18�#i�r�D��m�x��\���8��Wu%Ԃ���R�ۡ+�Ù }Z��fP�Y���A���ɑծc�1�r��Ӏv�]� gs��k3�����s/l*��O�ёʃ����$_,\9WSU��&S�����#U��,v4��E7\��k���7�0�"^YT���i��p|�2�f�ԾAr�����P/W%zT}�4vp�(���<9ԗe'U��\��\�w�*+Bt�Z�`��WBX[w���Upv��VT�(TDi앆.l`$�ԝjKj���"�N�-�Ú��n�+�%׍@���j���� ����7��y����Bۦ�M�7NIu�V�B���N��F%b�����Υ�����6�p�(<�xV��9��	��OM�!����w9���������*1(���'�Cs��>ep0��q�q���]|'yʛүY�_4�q�|��v�`���Q�i�mY��u�����Ңb	`�%��,m!]׫@�l��GV�JJ���[oně3�K�j]�N"��"���1�ru.�̤��T��@�5tE�;�f˵� �j���+Z�W���u���r��B5:��'�xQ髖�kk� �.��e!���i�f�D�;(7��f��!�P.y�2�Ͼ=2N���y�.����+��e�2ص��!/�Jv��Q̥�O8xХ�Xk��U����Y�^��}�����8r��j�rGm��p�[.=-�{#8
}R�%r�)��PS�Ѹ���<c#�-B�E[�t��=����C���j(f�]]NoY��eaΓ�T�U�����k]�7���b�3�;��(��5�졶�̝�����{.��:��w�hE�a�[]LR�a�:��ڎ5��,וz���:]h7�l�0	������Pl�s9�\�0f��`�!nb��=۳ָ.�ݫ3ݴyeۼ�=�'�!3�qCe��m�Ԏ�����u�#C���=�Խyf�E�YdEc�[a�����W�4�׎�B�p7�a�Z�J�{S��dn���z�4�Ѷr����.���t.q�7��K�C�5�u]ɓzD:`[1�-��&�dG�V�����fNb�K�ݷWEԔ_�ᮣ\C�T|.��nV!��br�*K���n2oDUJ��A<v:�"T,��&ԋ�����V��gc" ���gEH�[&��'qH��>���9CA���T���1��G̦� �3t�8��:`���r���]L�d�dY��_i�ݐV�N�eJ�����)��m��w��� Ѕ�t�P	�WK83�}�4P6�XN���hKQ��nm�H��EWQu�i'ʠ���+�[w��79I2�1�U�c(�3h]�����`��|��H�pH�9���Wg6�+�q��5զ�J�]ʣ���� :�6%�[��Sx^�v��T���4	mLT9�Uĝݩ�m!v@8��)����Kw6�,������u#�ݓ�*�77r'��0���`N�"�#�+#]�׮��5Md=��I)̠�V�i7;.'`��8�֍p�a��o��r:7�V�m��a�xp^5A�z(��V�%�9ݲ�w=�0k�t]���)i���r��&s�� k'n�S�/��(Ӂ�X]����YYq�82�˄n�=�|����b���X묅I#���\S�2�<.�+�3k�]^4�7�!|���l�&��x�k��
��f0�u�kٮ��7�O�٦�2�#�Uə[Xڔ��V�b*#����W���m,���	�j�G��\q(l'���a}Znq�]�����2]��]9��l"�Œ�T��6*�D�����*���hi.�G�"b�w����/ όz)�t��Nϖ�Q�|7N�3O۸�����V1Zܼ��l��
]n��Y�G%][Vur�g�0Â�Ԣ2<��N{�,N����K�m�N��AG������{��'���%L�iA�õ�b].L�01�J��<T%�Q�ٔ��Ge�P�k6�����&(���چ�;��M��]�5�zS'3�Щ\�uZ���9�ب,9�>�()���p��eY��[x�I�&EM&��­��f	�t��-gQ3����lF+b{$<�pu���{Onu����E�m�Ż��g��hMN�n�{zJ4�]�`�i'�ٽ�eGsm�e����*v�ǈ^
|�r`ڽ_<g��J0V�X/���,���"�R�c;��%�f>��j��������m-�)SAh����&e6��ΰ����^�����@�z�z�Gj@�`�'K�ܑ���ˍ%ݕ'ۈ�.�/�И>k�rY��)LC������o�wr�N�
;q��2�Q��{8��s���k�Smp�s��HS�Z�Q�<QU�n����%�%Om8iМ;����1U��e<�4���E ���ͽg�8��׹���՗wBR�>��s�w����G���;lV5�N�/��R�w+#�b70�6!�p�I
�O�ݚ�M� :2ʃZ6��Yx�n-QgFf]�k��s�c�	�v�d�9��Ӷge֧�M��u�7ϟ��
���P�;��̹E�l�C�S#F���z
Yvv�=:�(&�M��j��ĕ^U�r}�]�&u�*�G� ��P�vb���u%&i�tnpx6T��h�3Qh�t#x{D�V?�ac;��4�ـ�X�0��ee6���Gj־z4��Ecoq����:V��6�#Ln�z1v����gu��,��因�\Y�s��3�E2��)Zl`ɶۑ�ɧo艵,�bX2�Ά�,����u�ꏁ���M)�"���;K�3�m��;1S�8���x��)�p������*�ڒ�r
�$k��e�Հ�;��Rv�{���e[�6�ї�T��ڙ�WOE�`�ᓴ�X58ۨ�@��[�m��#�*r��7D�D�O�	����¬���tŅҨ���/�^��Ǐ.�3�Ԗ�D̺Tq3*��P���h�o��I����
}�	u�R�^����i����K!z
��F-'x@��*�����fR|�[s�s���X)�y���x�Q�7����9�Իz����U�TW�^A����qP�RQ��*>�-֚ytT8v�Ջ���v"!�鲁\00,��̲�e�N�(�whv��Ό2�5����]:wFnH�Z�����PS��ûټ�/r�S�ɽv��=1Vʌ��8����k
����nbB]H��∩�E���V�N��--��]��ZVk��lhq�R�o+��L����DB�D�9�.���悌M�"�YV��ym
�Dǝ�'n��&�;A��߰&���IS9T����2��@9[�|�AZ�;�-��L\WG �dL��'sCbS���YZ�M�uvZM�"Rٴ����;v>!�*э%� X� �\��y�,�������z7���y&���.r2Ͷ�iQ����S��B��C2^[\��#�9ө����ݬ�\8�Ԭ�>Z؇I�a�z�˪���VP�د�7�r��RA�Q|*��a�4�u����J�K3��7SN^ �PuL�j��iU��q
F�*uu�[��d��]Y���`���O'v��l��� ��T�e���-�۲�bX/Ve��k��6\��n`Э�}�(-�F�1��4�i���h�8!���0u�%-�J� I�պ�HA�ħ���t�%T01��'`j�7Y)l��]�S�]�Klm�.�y}���@K�f�>�����
�6*�Dߊw!����mIW]���\Ь%�{��t���tO,,�|�Q��e�N��|�KHK�9�f�Sw-�}�u�v=�<���S�*y��8o�ܳM�C��Ru�D��9;%�e�h���D�r�]r�+�����+��v�e*�Vݲl�)V��3y��ѹ��Z3��;2�W^�h�h�c����9\ͅOU]�WO)w"�3�*�o���<����s����H�3�� �ǃ� ��Y�p0��M�`O7_v-�Z�ȕ��3G%x��#9H>걹2�1ǭ؆���)�}i����qZ7h�q������M�O���,Ȋ�*;��������z�d�������x�
���y�u86J��f�)���h$�`�>��;�r�ץd��V�Cn���t��:�s�(s�[�Jjw4�bB���:�Y�T*�]�7>WRCp��H�:r��L{����"����L��V��^RPN	�&<e^��n�;�Ok#ѸRƌd��u%_s7o:���ڤ��Z������"*������,ZY�h���eh�`P��w89��(���XV�Ϋ�ƈ
��G���՞&�0M�u�4X��C����D:I�H� ��$_���M��>�n�`�Աܘ���a��<�Al��켌0(��Qʺ��¢��NaЋ�@���n;U)ǌ����ܵ]��t�{���-��/2170m�3u']G.%I� ��qWe
�'dW�W��W`xB��jד7��P7�R\��щ�ͩx�s��ȷ`����b���`Z�h�����̾�+���o��2ܶަ�����Mm_tn��#(��j��O�ej�
��m�]L+/�c>LΡ�Aإ�n�m0���1m��f��d�!Zf���2�խ��'�ZR�loFŊ��W�o7i���2М�Օ�k�v���`+��Ā\�:U�2�c#r���^+����{·���5Qݐ]��u�N��捭�N9���F��9D�}���*e�x�������iX�-�x�@��9�V_�]JnpQ_\7��v�O���ɢ�}�ˣy�_0�6�#u���,\>�>�Y>�
�>�x.S8������U�����z<vv��p,��Ťu�+�m�Fgq�%����/7�A�÷cy� D����B�(ڰ�أ|�6�w�m-��{;r���o`0
�z������ �<�
�x�ާ��v��]��%o�ϝE�I����ʍ!R�=�B�P���g�s[���za&�4tLl��E��,�&Ajf��j�D�l����c�۱9׃Iw��{��`:�hG��+!k�Pv�*1���w5q�9<�hn�����"�J��5U��
}�d�6���
;͊�/%ӈ܌�κ[���(A��e����!v;e���ٙVMvcBְ�V�FU�a��v���m���� �lL�ژ��ҹ��z'd=yB�+NN��9O�#G0��
O����U�=�I9]��jڹ�/��r�Y��;!V4k�k&W<����i��]m]w[�� ��|z���!=�۲��GY©��X,1hî��������؛HX��6���!**٨�뷦�'f�72���3WrT�=y�r�?����<�� ��h�8v�7Sv����/�6u8��n=�]��Ꝗ��"J��ڴ^�hk�A���ֱfA|�����&�T*�[+��x~����~��b����/J��v�����r;e����-Vi�%���c'�v�5�������JSt\��Brm����ȉu�]:q&��z-�U�Kb��#b�������]6�'�JU��A�ovV� ��V$M�tOh�5nn��MC�ׄ5�\�&�,�i��!��$)�_ �Nn�τ�[�t�b�'Y�{����-��44*�$�e���˦n0�>R��#���c���yך�Ai�Y��6�˃@s�h.�2�mP�Oǎ�jK6*ޮ���5g����6�ڷ����i��X�Z�������2@+�@_u���:wSz�$z�"���Jf�
9�3&>o90h�7:�7}��C��#Nr嵵e�*7\V]�sĭb��tm�%WZo��$�iLk��PT��f�-QS���5�1����L�|��j�h�ՕÎB�9�9�a]ȩ�2J�%n����l+����{}��s]m�3v�뺳{�@�)�F���3��/�<��҉�jTV�.N#����i�Y��ËS�%���o%U�{��[�6�V���a����S��e=��l�c��9v�X�];�5�-D������g�n��~�yVZ,Y�J!��J� ���T�A ��(�[I���
�J5�ĸP#l�-,��l*�A�a�d��%AH�-q��T��%T�*���H���U����b�((����Abֲ\� b\��*T2�
��0Ea[Q���EU`���)+�5�b,Y�PR�8�
�U�)AE�ڵ��R��I���Kl#�(�l
Ȗ����
[EQ�D1!k\��aiJ��R�lQamT�X�-+J�EE#mR�%˙J"���5-��Uj�QT[h(
(.8�"�ƪ��X��ĥiUkm(ֶىc+QTP�T��>�I$�l�޻�Yێ3:*�u��Չ�|uR����}[u�nq�y4�vr��.�Zq�KF�V��r�N���h]�gs'+n}-ߖ��ƣ��4qX�hL�V>��	�ٵ/z�,��1�N��Uj��eiU��8U��r��[%NTpL�QA�=���˪#����Ϋ����;w�~{�Y[S��ި�Cpz�e��Nj��ϵ�Թg�TI	q0=� �ݶ<X����f�s��Z��[�>i}�)������s���c�7����=0%�V��Q��h�ӽ��`��* ����̱H��_�Q�(����x�8�z��pԘFY�xTj;��iJ�5��U�M�~�l�n���
!�zg�Нo(c�3R%�D#I���L��pcὝ�F�F|��$;_�Jĉ���X����7(�ƾ*�J�͊�x��2qr%AgrSA�5�2��Iw�hOl�K>�G���+���k���E�s%��u�q�v�]ġK�Nl�6*,�72�D�b,6Ս�)&:�).�F�����K��6���w9�;^ti��k��.�<�V�Y~_JN&�T������I\�{g_�����k���g�����k�P]F5!��]����g��	������U*�Ee�:��"JV ps2U���FKO��1�ɝ�7��@�/n�ν��B���RN��{Mn��I:s��ܫ���U�81.�t�	�T��
����������,�U�m�_�He��}�y*0y����[����s�%Л�T�o���r̕�f��".̑��=�+�̡�v�(]���tr����dN��ﶦ���.�Q�{�=�[�^}�d�u�.0��N�U���6�y�c�
`�*m5�K��S�|y��64ϵQ��˸^α���ݪ-+S^�9�����]�t䄓-����ڹ�y��`�m���~��SB"��g�L�����7Uְ��A+{\���t	��ܗ��Wk�D������\_J���3��,���SI{'u5����"J=���uo��x]U{�}r�o���]��ӊ�-�%�f2�K:�2�+/iU��uyJz����ȳ3k�VP�l-����}����*a��6�J��P��og��G�oB��~��fZ�����g��b��3]C˸�W�6�:]���s(��j�ʬ��zp�M�d�9`�6Ga<��	y)�e�Hv�������ΰ\�r��T�r��Y��-�P������^��G��m ̄�۾DV^k�kM�[��s�l�yƱhb�0M��Y�1δB4r��Y(n�y��`ċ����'u�f8g,�̍=<�_.�}.�n�vZ�)��&�'K��Uo �f����p)Εmno	7�u����V���Y[����mNʭ���N��lɂ�ꝘF����$L�h�>ȼ���5*�==Ϋ^e��5>j`M��R.�sze"R�,d��d@�e�E����VU���;}5��vJ��!��ܫe���]��=��SA��X�U� ��Nk4�VdY�߽ǻ'D}T�2kҨ<mOX�R�n|���6���yk92�i:q��onpÖ^�Yu�T��BG����\�+y�%)r����D��vP�^ʸ�ς���zAS }}�h�c�k��������p ��?j�{LEnx��tuhk��e�UX��2皥�׫uk�;싖�-�����2������@D3�P�^$�#�!`�%�y*#]V�~:��$���΁,kSƁ=g��|1:�ّ�����# e�F=Ȩ�����X�V�ĭK,��4vc�n�L�r=�#��\��r]�z�:���S]�}+�pǟN��c|��I���1t�í�}UJ���5"�P��U�JuDh�D��d�msD�:t�RW^,ݣ�v:��|<rS_E��N�3�7�QN��sɰ}s+ +T�谶;�dC��gi-�iP\��Gyo93C�u�p������7�-Rc�Z��[$�;vj�+w�|�+�O;�މe6vZ+C��v��M�X��}����>U|)�M$ns�GZ�ԺC�8�]Ӿ��7��FW��z�s�Hx9��u{̊,z��]My�yՊv��\�u/i�c��㠶�I��n�d
 � �嶮&�⦰d���~�Բ/V����>7�K��6X1_�7�B�H�
ҹ2�I��k�DF�2R���?L�޳Ŋ����r�x�y�pL�]D
��T�w��䈼��o>U��j^��uz��u���V�+�Eg�kג��n�e���:��	�nԂd]9A�q�7�|wf��^e()��1#vb0I�E�C����S�O��O��r�(߆��/yI�������X#�JM4U�^(�u?!@�=�^����wy�>��{	��%�җ�Ν���b`�su�R�)�-L�d��ڼ5Z.�,2,l4����sֺ��ڴ�֡�"FÕ	1�X}�؎���_�j�����s��R)�� {��嘉|�^��~��
��s��!�8`��7d��F!�:�OO����ٗ��;�	���9Ё���Q�p�ɽ�z�d�HBi��m��� �^����@�i3�e%�2�*�˴���"L͇"�.��}��/����Y.��R�j�r���PV��fGD�%��4�i�rԹZ��f�\����Ս��K^�L�;8��~�{Z�� X�3#8�n噵7�Z�X6�{m�ip �;B���&��=����Ex.���:*/(�|=�h�۫�t����+F�5u�i#]���E���6�΀�^:��\�q�1��!՞T^��5��o�m��/il���~��g�|��v�$9qP�`=�*�4�K�v�k������jd���;���'':����t�ݨq�uW��>ׁ��c��ѫ̗[X+�m��\��
�u�$ݺ����Pgu�{\D*��pȥ+"3��'%NTreB�W��2_�e�ޫ��ģ
{�X.���HM��B=�,^��i�7�����x&�����,�3�^$�v�co~Y�+۩���+��1v\`��Ӏ]W���P�a��;1a��I���H��Ǌ͏)u훜��ᘱA��<�Pb�U`|��ih�b��ܿ�m�×�02���U�ժOv�Ȩu.������Q�
��_��Cb����.����cC���ui����#��5uϧp=�o&6l���2żT��^�Y.m�jݫ;��,ΰ�[�&�UӢ�'KzQ��m����b7Y�;��զu���G���ul�N|U.����v�e��]$�yi=B	�U3k��ޙwѐ���S�t=�k���T��!7�v�^�>9g=	�����%�d�H��+W>��e8�)���3$8
�u�gyE�X}8�NJi�5�2��r]�Z��2�(�۫ϞU�?�6W��@z�zpGg1>S�H��z��(�)P��bC	�锳��a�Y9��x��N�-�/y!��I.�*VI���[���q��鈿4��ߚ�"X��ߖ����8����P�t_��+o���t�Y�x[���3}&����
N��ߕRWҺzl��'�o`�}�w%[UO�8G���N�Հ��n�����7����*�ՊU�;��V]f�e�e�Gk�'׳��vLe߹�q���Â�EN��C��OR��%�kEI�oQ�ܱフ}�w��0��kv�d�⼰*�܃]=u�=[��W71maר���L^��
�s<֎���;�{>	��#4gB�3+H�˱R	�yx�so�����N�ܸ�}Q�myg+���B�Ԓ��zF5�yH�T'k~�n�p#�#3skK��2��g�`DZ��ǭ��̻��m�f,���a��%��*}w����ޟLz��o���
WƠ����y�����&�ֺ�nj
jWt�tM�GV�.ӷ��A����u(mt�/+8�!ح��A�m�>�$�SXr���(�IT̸t3�z*��b��,�D��DY��͸�T2M�ڵ\���g\9��+�<��L�����iܕW�t8z��-Pf���[߲��t,�Σ�CT�5��{9^=�\������v-�1v�=�+�<��7aP�igXB&׀�Mrx�����-.̗K)+��*I*�l̎�6g���H+�M�I!��{`�^�X
͒�L�mꃷ\���]�&���9�w�;�*�3�N�����0�k	)�
&L4H�'��Z��T���crhV��&�kp'��ԋ��2�C���qy̘<���pSE�e��FT~�T:W6��(�z^��m�G?|�B4DܦC3�}h��z*<�rQ�*�=�mKxۆ�r>y�ڑE�O>d�AJ��I5I�
��`'�n��p,!퍸C7�ז��1*�y�7Z�-��ݝ����tG˷����E���Ţ�"^凫�A���FC}�6���0s��U�w;�K�1�Y2�K���s�,B���U���Z�`�j��ur!�a�n�CS�݃�v��yţ�ɵc��D�ީ�9��w'q7Wtq�k�^��
̵dJ*��]H����m�y�oTZ��ʝ�}���m�)t��#�k0���n�F�/9v� �.�W+J���S㵢��s��Y����G�rǱu'��`�rz���>�GzB��D���TF��Y�f�5�=^<~�^�$��2p���uh����u�u�[������"�<���5�.���a�⑾n)@39f�����@��Tʡ�wk�q��y�ރ�b�c�����;�_>~~�V��iϨf��S�#��3�m���'��7u"�9nj�����mMR/O<6k����P�}�����)�tV:��+�e3�+���^��w��K >~ow#����1t α#]3�:��!���M�R�i�(ΐ�\�t�͹JH�y�4jI듳9�_6M*^N����"�U�r�V#;�6
һ)�RN���k�P������`�>��Զfu�4�%�=��Xz����By?J$W�;�VIّz#�� �[K705�z+�����&|T�l��~�{%aй�e�r-;�,x��N�7jA����ݠ�\�j��<��JkO��P�`���8�S�Q�����z\��S��S���uy\���۴6w���:il]R늞L���u�Sb�p�ݭ��v�5F���,4��yڻ��c�#���q+.k�%���du����|�v��Y���qNE��oI���*P����ۼ�x�G�<�i���I/h*9�����*]a㮾�2�Y��wGL�&Er�V�a�{'o-�7�9,R��JĤߍ�>(������]�
�#���j��VW�0Rsp��=+6��d>�/>������B1:Ȕ�j`�+%�c��9MV�uq�
��F���5=�����Ӣ�{K�2t��Fĕ	7W�V#�GEau�b��d]#f�iZ��e��4�m�Jf�9�a�dz{�2��0e�0�Dn���u��҆�EG�'z�jc9����͋�t�9��;n�OoR�f� Y���ނ�Ս^7c
6\x/�U�iĝ�_t��5��GXWe��|*.P�o��cz8NmՉY���W��1��p[����޸�|{G@+v�-�b ۝t��Wf���7Č��*��|%koT˔oT�3E������Q���`��S:m��;�(����^����OΕ����;�3�y"�5s�h���DC�o�Uݸq�uW �4w�VjJ�ؕ<�;��q�ȭ�Ÿ`륧ޓw���uY�S��`�P�U�d[.���u�)�-2���h�-zuP����%��4���1(n��q0�����z�[mZ�@wQ�;]=�4�����^֮�7��{b�Na�ᝈ�i[�P����;�u8�G'�:A��O����>�ov������gJnt8i��hh8���z�u`�e܊���JA�����̺�C���PΘ3��������C<����\�^�e�SH촷V����]RH�d�mi��,U�Lu�E�<þ=�F&.<F����1_el^n��~~�X�Qg���*�4�jSk.��4h����=Z��d�~T���n��=[j ��b���I�Q�ץ�(��@���`��Cb����la"g�=P]3�w&���Nu����5��6ɔs�S�!ߒ�Hv$����$O����T���(�{:f���+	`�46�,>X�NJ	C���؋�&R�T~o}��"�q�t�/ϝN�M����x�� =S��Q�=I̵�J�ؑ��)Hi1�I�F�}Z��-u�e�$�}�S�fQ������Jfy+Y7�y��t�[JlI����"�s�B�d�>��*��hN�E��B���qh��C�ɝ�V��K��\@�����3oAH�U�|���f�y��*:ڪ�M��V�)К���-[S�஻����OCq]��C�@�y���À�A)�WE�
��}���b�Pˍ���\dJ6w�
 uH;]t��E��,���˭�D��+���ӵ�Lwp.�y4�:��0<�k�֋ �miޠ�3�c�d���B���\.�'��y��y�6}���H�mq�k�Z��Ψ;�h�N��jC/���Ӵv>l.�9�v%%�d����� <k�`a���V�&��䳕
"/�t3^�ず��2�eE��ZS�y�A�a���=�Ӛ�;i�.J�7'�'tهc�Ȧ�z�q©���i��"���;����S0*�J�vQ���79���\5.mq�8�
��c|5n�h�_sv	�Vb6(��*s�%q5v�����O�kN���e���]@��u��1�ׅXr���9g.^b�u�� �gcYM�\��5��`�-X÷��k�
t���m�|��{׎JkF��
@L�������ll�ST���4�에^�ᦷ�yO��ЊV2�jm���#Q�6�g%t���P�,qT�E<��V�;P�c�n*�y�QG���2�3��z������j�}'	4ӥՖ��	�Z7����v�7%
���A;pzɼ!������0�>b��Wj*�xT{���Ky��6��ނ�Wz�z�k��tS��Q�8D+p<���A;[�s�� �rJ&Х4��s���-��=g�Yx��E@��+�u<�]kLe���xӬ�N���{s@ze�yWv��gL[n(sh�:̺�v�U銉�,QM�$�r���NME{.�����E9��Y�]�^��!u��n�X[N���Yյ��w'H�k�T�}��<�{v�ucz���L�I�ڑ�Om��5*���έ�
 ��[��ݔ�,����T;\�ķ�uS�0_p�dw�S��K���P����3�X��9NM]���!�{���'��!����X�-�e�vR��k�sa@��^0.��*�n�i{a�����̦,`��
�m���6�W�H�a�c�o/s�@[�Qp5�4G(��L���m��[c�p9��f!|���-"v��[�o��R�s�f�`���g"DQvU�
n��;1��:8������Fɤ4`\�1�W���H��ڽ4
�|LÇ����r�45�5��vW�XZE�fQ�EgSDAX')��Z��tq���λ�|��N�9��"�]қCY��꾼�+�(7z+��]Y�ㆨC�0j��W]��:��t�h�th���ɪū�OP�~[=�P�O4X�e���8�q���S���RE�N��µE����a=k������˶O\� 
�r'��U8�q�IóF��uSw�9��F����	JgZ�Jpr9����Ӣ��&�V�ȕH�F�[Qq���� z]c�:����SPk���ӂM��_A��WL�)�]R6�������ˉ;�sv�˰P���P��ic�V֎[�R�b-.faq3J�YTE*W�2Ҳ�ie�%���-F�-�V�+F��m��kX1X8U-��K�F���h��db��F�
�KKm�5KQQEJ�R�T.Y�T��U���b��,e�-`�(�J�mm�1R�PT�30��%UAXҊV�ֶ�DYm��Kem��FV��U��Xƭ�[X��D�)m����Ң%�UEU�X�TB���0�j-ER�V�f��T��(ֈ�)hڢUJ%cj�-JR�q��h�DJŊ�-����-�+KU��UkZ�ʍ,UF��[ZTB�("�%[*��h[K��n\#�ֶ�"ՠ+�e+Q�"�U���m�,J�R�l�Q��V(VA�kZ%�-\J�PE\J·.*b�����l��mm�DP��T*��%�J�m�"�J��VZe�12�m�f\�6��Q
Ս��ʶ�Z��Ң��Q�JQ����ֈ�ѱR?I@���RO�G�l��v:�d��3�!�|\k"ә�w�w۱�ʘyf�87���b�YU�]J|jؑ(%�:x̜�Zf��W�j�),���y�B�}�eǪ���ͭ�����ɶ�#
��`#�&޾�s��c[w������3Ԩ3*,�-r��u�6��P��g������,���&�s]�oowD��O��جL3�MxxT�]Z���B��7�c�f���f1��?Ovi��$���y��`�&j"G�m}(g<�}(W�$�R��k���!���a�����=|��ܦ��(ga�"���*h���1t_g3N+0���I��	�)ĩ̏�uo����ψ�8�J�t8�A�A����uƆ��H-3�S�C<�W�d���m�̡>�Q.�|��m���W�x6��T8Y��M��4!+r�'�=�lj�4Jx]�����S�W<g����V�H+�L�e�Hv���/������涚��.��O*Z&7X5֑i��Z�i�~r���S�dq�J�Ă�����t�I�|I؄Jyx��V3i�sz��C�VE�9=+.����}�~������;�aJ��0�r>�;;F�Z�:��*r�u{r�|����b��N���yh����ܤ�#��>���Q��3���_�-E�K6��ê�PT'AW�<�}�E	�!�\
uw�q�����\�k`s��]��N��B:����fw9ø�uZ�=�@b�����Dvj�E�N�e� 1�e_v��
�Yt�_N�o}W�ޚ'��u+hU���H4w��m����Y���D��&�T��K��9�蚋��3mD_��1�,����]Rjʜ+�̥㺰ZdK��l�Op�����~�?!��vG��.��*�xM��!~YXޘ��ǅG~>���7�.-ݵ�̓���c$����OT�.���e�y+�5#�!gӬ%�	T�c}2�9�� G8�e߳}���R���l��8ͅ�uh��n���!2�#��dTVD+��n�/���K��)�W�P<2�����.}j�R�K�ʵ%����r\&܍6���w}��҅�Q�2�d6E�Tdv�dX�D�϶�46��o��nU���+��I�w��KH^{���t
���p����"�d_"�A�S�Z`���;yj��ٜ�ͳ��ܦ�lC�i��7��xv|�>�ㅵԞM�R�i��ri��Q��)]���������/����\M���>We�Ы�3h4#i��q�6˷F{Z�S�tkU^�����^�7u�r.��Cuub�]C§DJ�қ}ֻ5а.�t�[X̤Q[��˾g�9]�z��(ގ�]u�]��}it�To����6��h���4+]��=ZD�+J�� �Y��y��7/|P�%�Xm��\�#�BJ.��Z1a����wGK�-�@�[��X��:�30C������O1D���I�����kmY����ĜkN��X�^���;ǅ�^���;�s(�JC|EҜ�"#�➢l/S"�;lV����ˎ��轸�;�]��W4v��-^qΆ��S���)Yϓ�i���)4�/j����9��|(���si;�yƵ5�^:epu��VQ�Iv!�d�\���Vz�}p���U�J�}�ݒ��f6�Z�(R �`f�h�˜���bĕ	7�m^�QZ������1ve<1��-��g�=Τ�F}u��c ;CbƬ#���k;������nw]j9�V�Ʀ@��;��^V�_�;{�ʇ�7��k{���G�n�̯1G��jy[W�4�*�;$��o,>���o�fQǕT�a���ST#)����2�wŜwv4纄�L����gwk�v��Y7V�ڇu�A'&�;�H����wz��w*��
�
��4.ޝ�����I��� �C	@&nR�����\̹�6�s�!9#�[8d�ظAҞg>.��ꕑK����4ZgR�5:'��.���յ�I��F�V\��s��	�z�7R%�nG`�C�(�#uw�~Y��#z�42��	'�qwf�'����p�7w⓿>�Ud?2NT�̛s]c&z�&(͋�!�I37���6rK�)�.N!��b"�u�UN'Up{�;���x�tV��p%��,ƥ钦%/�ގ�V/�:��mXޖ��D*��2-�]a����IS�jRŻ���)^ުw��l�7��0]QQ�����Z֥S��^Q^M,T�ޗZor�TM��W��7����g�$�>&|Vi�D�i}�������������8�&<�#æ�<S��]���)�����A�(p����R�Yu\Y�VE�������y�lM{�P"�ͻg�a��3�W�+�D�@��`��.��#��T�4�3|��LWn4�'[��t�2e�ِ�d��%�~�.�_=�,vcmIM�����kܫ��<g٦�_���Z��fXֳ�-7��{���2�
T~ln(���6���P@-G���h��{��=�ԧ��3+�Z1�l�2��u,��;77Í���`�(�h�_I�.j��K<fgN��4ұҺ��n�o��sē���B��r�N�4�k��t&`{�ʔ�Ԋ곲�)�~���s
ϖ{��.�;ޱGܜJ'���j��R��Z��leL����.=�r�ͱ8�<*�L���r�Hݥ��k��n��:�刮�"���O
�]�tK��L�����ќ�4�-Ղ��y3���>��I�^�o�^K���鍰){�o�O��M����;�U<#�u���ӡ5� -[S�{�	��'!	C۲'އ��3�gy�q�����a�g����;Im�+�5az�E��3��\�gjU�X]�����j]>��+�L��Õ}�P��3鵻T2J�^MuQ2�������r�s,iRE$��s��m:@w/}���X=s<��մ!ج����� ���^Y�;+�;4���{o�7�ل�PG@�=�t. V���oJGo�-����//(*4����mJ����e��k�!y`yM%`��"IN]��%���Da达f��B�nˈ].�ʏ�\�u��tީ����w�inJ�+ ����<�A�U{�=^�v�q�Y��>5���W��y��AP�EnTT�X+K�:����9��}.�h�;reLn��pH:^fq�R׫{��^)�JWm���[��ͳ/��ث6;W���8��ϯ�,eڐ&t{{lnhjЂ�̮�W�g&'�h=���t�&��u�0�a�څ�0u�J��Q���;�+�<�m|�C�9�|e6�c�۫�8�8��>�A
7��w�;h٧3�t�u?�;��y[X$�l�I���X�{�x�	um�;��*�aOҰZ'�Vl�"�wܵ:�'���{�>ٓe/l��W <|��ՉiH��y�v^��G�K�h���PK�x�=�x���1��P�!��dN\��-��L�wS����矫�!�XF�RF0���S!��ܨC36�}�P�To��J֟9�����Wu͒�,��Sc0���-�䤚����Q�/�(���XC�p�Wo���7}���咻�ڤ�mag���r�7�~����ҩ5eG���8.�g�z�;��6[L��Of>��ЮP� ����e��%W�<&r
М��tw�5����f�D̂����[���N曻9��4�ڤW��Xg���ި�z��q&�w�,�)ʂa☚�
��o:VWY���	�b&;($��=hi�P>{\~���R����}V�2��'���K�#&lOr��9c���[�`�8�iEx.hk�c�Z�`�և5n➉�\�Y��j䈻��S$g<��[�a	x=Ȝ>֩6v�rf0�WJH�uY�9c�}�L������Q]Y���rl�a s�R�V�$����^P�s��t뫡[�w"��G���<+/Խ�k�mb7��P<1��;*�pkJ�K�ʯ[}���P���9�9�m��GGs���5�x�,��1�.�^C�˲.�;ڈ��S��=�{5��t�V�)���C)y�%�g�r��>~}�{^�$P,��*����1��\�F#��+��p�e��[�I�=С�8�E�J�߹XK�ϙk���mz��6�H&@Ü��Wo���}^�c� ���Ѽ���P��t��k�bq����`�+�,�������'�+��wk�D�P�(;�,]S�Z1a��ߺX��o�K���JW��x�orj�$���Y5�:=y�"�D�+��
�F������׷��˖�������wh�p~���}_,)�8n�+^a�֊�8��OW�=D�&F�A���ޕ9q�)8f�u�s������AUѳ�O��C�b�x-5�V%&�h�/W'�6�	���+�!��J�$w�L��=��ru�G�d�(�.�#u��uYMք��}Pٷ/�BU�A��T���A��87Ebˀ��p�#���M)��<.��v��sR�� �tq���:�Kq9���tuu��_.omK����x��w;=w5��.)c��IN��q�:�L����g���[�ܽ��B�[m�S*�ek�����͌G39�J �.��>̱��{ٖ�2$lIP�`F��Ϣ���;�+]�m�X�uy�wk9w�a�ɷ�)�����p�^e�4�;��4�"�u֢�����C�ܝ�F���Q�������[ؼ"�����ߜ��X�s��)�����1r��Z����{��yl��}�T�6B��OT)r�ܫ|<�'�۫
�ǒz�i#[v��V�!���Up�Z63��6��*��] �Uٮ8��;�C���o���}X�	�*{�o�6s3��ݷ~/S�58���Iʃ��̛s]c�u��w�{Ї&LU��HK�ϩ%G�>�jd���/��wpâUY�ѝ�yf���1*pJ��Э
���s�.̤��D�d���#�o�6����ci�
���h�XDƺ���yQ:�g�./D��Soj�N����QP���(]$G�u�#�t�������W�(�����89�ۏeRk���Vr8�M��1.$�΋�m`����}�Txha�^ּ����C���>(���'��)�@�p�=��Um�n�Zt�Žv���{Go���Yu��@i�>��[��q��n�{��2�ɸ��f�Z��
WI.w-��D[�R�,��qy��L��ع1�&���7J<Z8�wm��{ڱ����周��}����{ϧvݝ_�E��X�lK�}��-�҆�iJme�qf�@f�-��{������Ĥ0��?F�fN�,�X��9K֙��|���Ao>TMzQ��8����j�k������*{�!V}���yI}˓���aӦÙ2��w���+D������7zף��u�t���ި��
XU��9`N�%4cZ�-6$�ش'��z�-U<���Y��]�V���ʩ��qp�DW{�(��S�E�:b,6���u樎��dY=�[E��=S]�"y"8g5���җ/Y�k�Lva�J��5�S˴��1Q��owc�v�7���>���hG�����T=���zτ���x>O�����
�]U]���(�=Q�{~Ui�#kpV��T�$p���P�t&�!�[w��R�|j�x�����s�y�5 ˠc�U=�N�;��eǪ��z�h�֮d���x��,�b}c�޿)Q\x�N���P��
��C�<��r���.�s�Y��*���W��JQ�r�4+�>s$=� <���i�K�&&��th�fw9N2wG��]z'�u3g̪k�|'j�b�v/��(��d�A,s����Z�X�Y���ܕc���9gM=.�z�{����KTd�2���f��r�.�>�Ү�K��m�����\W�{����+���ѳQGR�˭���r�50k����K�]J�Ϣ���7�cGv�䑍�yAm�"u��Q=�a�l��PG@�=�:%S�k�_J�x�/�
wRJK����:��r������qj�Z�*���4��C;�!����>�D��Dh��}���<�WN�Y��r���.2']\_4�ş�q廊���p6��<�RP�8���DFҡN��|�z�(y�.,{D�7��i���J�d:=y'�m|(mf�/�����]���s�}e���2�P��{�������;��y[X$�}��$5�=��R�ߤ�̀GmQ��D�Ճeiwܴ'ZD���{�6d�X*vag;T���ճ��Ƕ�A�Q>���!�
	y����5#�%����Bb����T2)��r����v�Y��A]$[�h�P)��ەb ��R/�ب�g�W���i �*�f�Uf�d�1����$��Am=�I5I�U	�����`�����C��n@<��F���G���)λ�%_"��!.���Mh�p�UM��\�Z��&MT�Ūd7g��3Or��M=
 ��{��A�r�a�_s��L�����YzV�1s,4�����I���4�nJ}Zл[�K�Ve*����0[�����:���q�í��1��WM+���k�871Mv�e�օF��t\��7�[cR>tGp\���N�mYDW���>"�<����U�+ZF�)�,�kUNt2�� -ne�e�ѧ(�F9ǆ�(�M�a�Q�@�Urh��^�T��m�����VO�×X���e����+��'hmb �C�R��l���Wʜ��2��f��r]`��	&ܩ���3�oF�p+�X:i�Φ��j�B�ۛ�g]-�޻�nCXe4N�Ы�엏#L�(�kv�ٽ�H�.(�W�+���q��w�@=��,M�냧(鹅
��ox����wq&m$I�K�h�T5"v���l�`Ⳗ2�M�e�h�G�� �Zڎf����o'h3h=Zlo;B�o+�������q���ïRj�(�[����V��p�[��C{u.T].��g��M\�B�y��eL�y�6��E9�]h`[��!ڂ����V�j���d!u_s��� ��2���6��C�w1���V�J2R�|.��V*奼>�t�\��OeZ�7�	c����������g��-�}�=��"I����Kdlq�;많����}�E��]��M|��/��bA��q:�p:	P1R�/&�Һ-�rY�.Ton����''�8��-THL��q��}��pU�`�;2�"�SA�k���I���	a����H�nY��HSקq��y|�l��{���:1�.�b2�bH# �8���\��Y3T�i;�:DW[�K��]*�4t�I���W���[@�{�זk��3i��:���+ljоR������
�ܸuܬ��b3��k�]��u� �<zU��9Vԃ4�x�ٸz����sH"n��j�VH$"i )}2Dl�YدӨ�X	ѭ���l�E� ��w����2�;ۍޞ�K�f��R�8+�ǴJJ�&�̠���%��C(`2��{Q�K1�mv�}��Z�f��}�0m�7�q�E=W��܉�%U�B���4(cI�H���k��,�ܳ��q}�b�xjZ�1�K+%LU�2%�Y+o����V�c��L�$Yut%���j�[\HT�\�i'�Ɗ��zn�`
�ơU�;���F�I��Ν���e��՘9��
u7s�}�V[���
x���РPg5"����e��9�%wa�Tw�pGE���pn�:��P�4�^��狢;�	B������Gt�L�]�xKY�g�r��0^���Ⱥ�ū�3�[�w�2�*J�ޤt�+w��j]ig;A��#���]�,���>~k+Qj�b�b}jȸ�i�QQ�e�*%�m�AKK�Q�5J*5mFƫQ�[�\)YV�(�3C�U�meE�Db��T�fXֹUb5+m%���*��KlJ�+Q��K�Fҥ�d���jR�)U���FKj��R�̦b-�J2���Q�Ɔ&d����J6�L�1���j4m�����j�-Z��J�b�Qk+)e�j���W��1E����V
�[Z�DZX�Q--�*QfS+jV����+F[lj��eb�R�Uj��f2���h�ʢ�q�1Tm[TR�U��V���Ɩ�
���эYT�Z�m���[J�Z��[kh�EJ�2�qAZZ�صkjZ�[ذ@�lTX�V��ҍ�5*��m��cFV�Դ����hV"������k33إ�mmZ�h����b�
��[���ߋ�ĝ�S.�����s��kvZ�Sw��7V&릁���W�H���w	��C$�����G���ﾧYӕz�s������v���1*���Lt�F{��~KW(����!��3{�z�����������h�"���n�w��/%�ITxMΠ��iU�zg
<4�Ҭ���bSgZ�{�=~���RF�����.�<��P}=w�Ҹ�@H�H\]U�����%U��l���,��k�<^nz���,�[dh��\�_U��;�ʹ$uP쩎uo���S˸�C.	�Q��2rW��W>sJ�>^'gظj�VL��q�ԯ
qлe^R�Y����_���5�yKw��%p�u�o(�y�T�$*� =�����v8�pM{���7V�36��0;��Vw�r�� ~}�y�G�d_+
�a媜����7�y�����`��*���vM��-��o�v|�]��KkԞM�R�i�7̋V;T�,�>��Hmږ�ɵ�5cT6lg;M
�@���6'~#�ZWpʫϺ *�(W<s�knyu� 6���Ju]Ҭ���Ó��{��Q��vRt��x�\�eݸc][�̮x��ގ�f�vF��Bu��������W���α L�+���=VG"o�X[�ً|X��٥�J�������b��m�DV��>{]��3fN�nj���Z�Ӽ��R�sKg%�o[n�����s����XvT��Ͼ�<��ۉ�(ե?Pf`X�*!,�a�ŏ��Bģ��F�&���]��]F%��79s(�3d��)�Ɔ��ul��
'����^�Bv�V�P�7��|��{ܟu����o\S�4����bx-5�IX��r��P��Փ9�@>y�܍���
}=�(X͙z���<�9�⦙zf	VQ�c�.�#��K��p	Y�z�TB��ۢ�eIR^���Ko��.�;cr�{	}�fZ��č�%BLmVEEj�j�����ՉrWh������T1�ك��91�hl^�@W�^e�4�;���q��ȗ�ڰY\N>|�4f�҈�;,>�}W�WjӶ�b����ߞ�pW���Y��x�"�z�{)[�:c�Uy\�\�(��,E�.�[����B0S�+v���,���q��<7����ܢ?i�����Y��O=p��]���;�X�dn�����Oz�gm�d�<�p���/-D?]gI�w|�B���皜|�cl�T:��%ѻ�u�_D����L��n�#��BT�.d�Íc3�ˡ�3K5��/pӦW>=�<�-.�����Ok��d{�ژ�$�ε,�|��|0����{�����Z�:�Ki�Cs+�y�GxdD���KR楒NOo:�R`��+Z����xx�F�
�S�����,F�6��7��::��8���h�f���1*k:jj.^q��5Ε+���g��*��X"ܬW�}��"c��"�5zq�z]}x\}�kPA�j�����PѰA�,_�	V������PQ�s��N����k�Ct���'�����zt��[��e\rJ�#�/��xJiwT��}�Wǆ�:�W[YQ�ʧF���60�n���2z:�:�#���g���*QCI4>R�Q���4�F<�V�a�u��Ex�������Y>��<)z�./�]��-�N�6"�ƶ��nMa��[����ݛc����k<��t�2e;2d�䯌u@�pR�Wc�'j�'w�>%�T(�ƳM`wX��'S��JB�]�C�Xѝf��w�pu�|��ǺM#�P��|؇,	��v1�'9��0+��Q`�'2�D�b�)����L%�=����Z�ߪ{vL�TÃ��L���OgrTi�va�\��^}��.[$����+X�ד�c�)2�<�K��!�6*�/v�jU�=YR��N#����`�GHv�E�'8�9Lf���w�g8��n�>�Nf�.�*����
�s]6��nB����ɤN�Sb���}u�����Z]�_����<]�u]������~�`���	����;~9[u�_�He��Lu����Tn�����x����ٝ;�������׻��S��%Бk�n�5ʽe��*-ǋbfTZ�ŏZq����l����w����/�}�q�}^�7ۊ)�����.;�2?<��N���t;A�I�[�W������Ta�Zoï���WiV9sb�l-93�<wݚ��۽��a䄫8;�ճ������!�ꗭp�hC}�ԝJR�E��qO���W_�dc_yc��C�p�}My�� +]�����Ύ�*R�m#/dC����һ��SJ�S��u>��Ͻ��G踒�*�>	
��^� ;�VuU���c���Z��y�f����X-���_˭,��4�6$����p6��:(2k�\�gO.��o:���ߪ40:�T��6*�@���qg%w�@�&���7j�%�V���^m��<�I�Rs�\Ӑ��tX��20����q��S���c5�Ѳ���ɛa�:Q��t�j���,�͔�t@����]�[Ԃhw+��5��L��͘R�����i��p��G��l�읊��(Z��)f���{X�
K8�.��[�!0�znl�9�2��./�B�7�N�������K�� =�«��*b"��dA� �.b9u`�`\�}ө֑<�[�%���]�#vC���h�e��w�������+S��l"D!�����,.�H����ߌ��CՋ&��>ѓ��s��㱏S�c�
�ʴ#`�H�>�S!#�*�ͤ[Y�������k�;����?*3��q'�P�|�f	*�[OrR�uiC=��h������tOo&��ٞ����Ͳ7�e��}ז�r�%V��n;�@zx��;��υ:£���U{xVұГ��]��G���:]sP�o�nX�dM�g]�U�;�����Ta�^�h�KLE��c5�7ٝ��l�(�q�Qߏ�롄i�5tV�Xx����(�mS7>�Ğ^::&މz��fj�<緣��6XK*$�kM�u�{Eҍ�8h	�l,�FF�[�s�v��©��z$e�ڛ-K;6̇�-��E٤2��XNOt�PX+�%��3�TA@���p�'v*iS�8�j�l��`��TD8�k=�1��ę�#Hv�f��z��	�g�Y틨�e0����QX1o�5j����Y�C����8����%����<%O����!��+����F��gk(�Xfq�E6;��T��Ç7��҅L�+X|��-�J^��y�^S�_R�D�j��+)`�V$��N����� 
�J��l�2�>����_���F+���C�64N�؆�[�)|8S���]9]����/rg�¡����e�4\�d��B���xv|�:��;�ŵ�O&�)*x(NZ{������l�����-�q6�5�;��v��]���	�D��M�P��W'��Ǳ�l/k��K��08����U�+rr:�Ic���Î��� _�H��KHܞ����=�>�LƽԈ삉oq4G1uON���rr٬�@5���oo[(��NF��b�*p&Y�RL���eD��
z�>L���k�w���Y��(�k/\�h�o��#S2�W����}%bRh�j�^(�5�O�7�6e�nt�NL*2$>��Hu��d_9|Tߌ�3>�e7%؆���1�ͱݜ��.i�}sY]�5u�o.�;�B�a��޻��x�����I����"���-�^cݥ�^좲��z�ɿC��7�͘:.���0���~�̵��0e��p�2�D�.��܄�Z�Eپgj�����;hp�mxp��O��x[�A[e�{D���ڥ5D혻��+��a qbonY�0�!k `�j��6�����>��5%�u���`;د.�G9�i���7ǭl��5
F��(!��3�.ۋ�]��VL�׭)�L2�.������4s�s[��:�c��0),���]����k��:�Up
���S�]�Y7�g)��M�'Aj�\	��(���T�6B��U�z�N��Ͷb����9�Nd�W��[Y��2����9�A�\;�2�ld4M�^ Ո�a�X���eQ�ڻ��Mn�os��#��
��>��;\��iߟJ|�c'*�PfM�����ET.��k���l�d��R��";��2M{��Z���*��t{�=��Z��]f�^ۦ:sx�7���Ϩ�p%�] �Y�z�-�@��D+�C"`;���V���.���Jg��eR�Gʅ��W���,�8-}DE:��3�dY�����)�i�A|��Y<*�p�=1�Q�K��Շ��L����K���#�=0�aV�6,���g�>L`|{��Xz�3�����11+�Xb�XTԶbx�ɈK�$��X�٤4��~�0�
E�0˛��?wە��3�'x���	r<&=��LfϽ�=e}N��I���q&�3�~`T�~��,�T���pXz�a��1y��Y�q8��i �H��i*J���L�,��Y�~�}�{��]�<���{�{*m'�WԨi�&����<d��"��!���'��=�r@�_̞w�m�����I�ǌ
���Dd�w��i���N<k��8�3��o5϶]=�L�P-��s�L=�i�lx���M���M�s�tA�x�ei�X����t�]};;(}��P2%#���Ԭ��/���Ȝ�-�s�7���m��L�t����Q�N
H��5PO���˰�*X��!2�w�_}�}�&�O5s�{��j���,>q8�d��b�Y�����x)<J�^;�������cL�CO��&=eA�*�Y�%�w�βx����]�Ry����9@L	�zb!ǽ�*�^���U���~�����R��OL�1���3V����At���O�Hu��]5�PY�*h�SI�w�ɶ,��<�̚z��1�Ρ�^�D�C��z1"��V��s�1�m�z��n斊4�2��z��q��%{�<��HT��S�d�
E���?R�a�i���OY_��4���x��q�PS_~����J����q�Sc:�����K+����9�w����> T�����{��A}I�sZ���%@���z��VwVLL��I���z�
LB�~�Lx�d��
G�k �i:����rM q+����:�0*N��~��V�}���՛�r\�\�T�������}��I����;��:��&����Aqg��^$��1 ���d�����a����m���,�Ri*A�Ԙ���1�������Q;{�ki�.�Ø~+�V� *
�0��5�<d��|>�d�����}��m+%WL7;��R)Ěw��^�VJ���3�m �g��	��&�Hq��]�*>Om�=C��'��5\("����7�v�R� ��6������c<{�H/Xu��6�H�q+6}�a�O���{�2hT�����>�ěB��]o�j�R,�{���y�B�L�(i�UO��>_[ꓕ�`j��Yk7����I�mư��>�*Md<t�g䬛���La���j��"�3�u?!���>�f�yIP>��d�+=�9�I��B�'{��"�`	����<5������;��~#c��t��O{��?%Ld����a�&�4���Z�O�
��M�i��i��n�"2u�17��F�Զq���\I��ï�?r�$=�oZ�"���051'ﾯ��w{�5D�yo���%@�+>N�������*?S3Ԙ釨g�=�?��1�-H�m+6��~d�~7���M���_7a�4����=I�)��O�F������*��}��Y��fVũ9��*�JD\���ݺ�L�;�D[o:��cMӷQ������v�l�X�%��ù$05�j�&nf�!whbl]�2�kka�Q{�d�}��W`�&k��+"���QSv�㕲�dĘ����*Ȝ̵\/u*ߵ���tlc�\bW��=� KĲ������{z�H.�7@�����9�a4���,�ϵ*��bC�̝B�f0�1>9���1f"�H.�|��M&��P8�z�i���̘�0�b	����ֺv����4}�3���|̟��O��(t�1��R.�a�
��!Y����q9�M�jm��Rq���$�
�S����`��7;܆����x��_��������mf���UY�}��-���>RV�Ld���~������
���i�I�+7��&�����߰4�R�6g>�3�J�į�u����=`T=�����̘��'��D==��\z��2�i_T����wi���t�_Si�7-�I��1�L� q��T& |�����6�O����<gRc�����Ă�~I����SiJ����z�|�ިϮ"W�P���l���b ��2f_�<��J�J�U��~N��_]�TW�'ݦ��q�
�É�i<iԚ}`Ts9��>C��OL�M3�+u���y� Tz�Y6��~{�U���[��b�L;���x�%H�y;�h�+
�����"�B��{g��I*0�����F\g�L�HT��Y1���<g��'�ݧ]�P����s��1�Q��߸�y��,6�6�;3�L�y�<��x�_̞��mS�bA��,�RV~/2Ld�Vs�yhi�I�4ZcĬ�LB���_�Y<t�j �"?V&��z���V⭭�����8�f2T=�k�N&:`T����~d�Ǭ�^�4��5�}�M�x���'�S�r�㴝�aٮd4�AN'�� i*�̜O�6�M%e�m�������5��}|������H/Y���2�P8���a�&��l��ևR����I>�rm'P�Y7�oK�
��M~����$T��m���SL�C\ɨ��@p؜�?|����c�ǟ^�$��
��\g�T8���<7a���8�g�a���c妙��^'��u�ҤR~>��l+
�v����RW9ߵi*w�h��X��u��'���ό����2�J[Y0�n4~�i�k�}<��5A#4�)ʅ�g��K�����
�n%�A��KG_t��G�O�Mze���P^����g%�꼤8��"�wB7uhR�5%�0`��Y��؆�]�����=���% ��H�i��+ڒ�=��xoj�,�N�_����`=��g���ܥa�1��X}��q�O�W�Owf�Xx�=K��!���S�i�x�H/�Y��u=C?}�=H������d�i�����s����/���-�����`L|�A�Ԭ�Lg��6�\q��N���H�bT�7l=t�Y+&�x�}d�c��I�+�&&>����R#�&�8��o&�d��1 ����p�ɺ9_^�e]��b�yl�Q�:��6��S���h%@��
�S��M%w�O�bL3ù��m �g�塧�*E�殙�%ݟ�1<�'L�&e���M$�+�����
EW�'�oŔw��"��L=�]����I=��l�z��i���!_�'�~�P�%0/��A�~eC���fH��+q�-?&����L�?!��VCI��5�I����â�~�(�G��xLxJ~}g�i�T+��<큉*>�1"��~��M3�:��'��M��J��<3�]I�+���?`q�>$��N{��
�R�i��EDب�r���g��Ƒ߼.=�:��
���bNɺ��eA��M i+'Y]�O�d�J��߰�q+"�7�4H/2x���"�ĩ��}�=|g̕���N&?�z�T8gTS�_&K�ߔڭ(����I�+���_�"3���S>M��f��~L@�n���$�(c�:@�߷�T�I�>É�bq�"�O��ͤ��1�;�C�����=e*�*u|�~Eu�=���"���Lg��,�N�P8��əx��I>B�f�C��PY��)Ԝx� ��d��O�M3�yd��~Cf���I_Y=��m�e@P�Q��������nG�^�˻o��*�:oߵ���w���C��i�?!��R.�;�)��N<|�I���Y�f<�`bJ͖�
E��&墑g�8���~X.=��L{�ﻢcVSߪ�I+�����J���˄��q'�+�=9ܓh,?5��̝J�Y�?k��x��q1 ����H���uC�{��R,�=��C*VO�k9�*T�(~CO L{� G���p��z�a���ӄ�k��T���݇�v�e�ÕNb���m��4'*�t1>ǚN�:h\�+tdI=z;1�Ŵ9M��E ���3��_+�{�d��2ƭ3"�
�ݙ��]�-���g����(c�Y`%p5��'3��(��V��$W7�v�e��N�=��Cy�U:�p���6���*���1yDf�3zJ&�ޛl:ÍZ��� DR���x��}%?��/� #m>%6kՅRn�U	L�,�w\��Zq���j�w3���I�2�a|�`1�� ��|p�ai|�W�U���Ů+���Tв�J�]�f�rk�Cg��<8�­aЃUE�T.���M朓�B����̢�� M5�( ���+C4�u���j�X�u!7t��{чz!b��m�0�8�r�]��8��@��H,w���g8��n�教�f�/�f<O�&��JoL>և�a����|Vu�eƞ�P���b[ �#��b	��J�XN��N-8`���0ͺ�]>d�uv�0H)�gM=�Зr�1vm��۽X��;��Q�����wt:�0��:���r����c��x��<G��`ց�	��Y:CV+��i^b5pj�Z��aat���P���x{dg{�&M�MɽևN�'eCɳ�P[ta}���T�a7�^R�o�;����qE���吪��SiJ��J��tE]�zFP�WoY�IC�L;M��y)��7V2*�m�L�r�fb�����_A�|w$�ʗqH{D]VP��QT����5��A�YVލ��0`<�r��g.�Z��=�C�O�u*�����S�.�[�ڐQͽ5�x�RT�s��(!���ʮ�-ǕҢQ�9IQ+[Kk0��tMA�!��v�aI��r'��t�p�%3���cd��\�#�9�2�<'n�F��E��8��|+�s�p���쭸�:�s�&������i]bt��[��Y|�eJ�`<��a�*���`j�ެ�C$�8RX��0���o�[}�� H��s�C��wM�ʂ�`�{ը��f�ܳ��� �w�z�&�:t)��Å�б�/���`�լaĬ왤
K�v��d����8�n�!m:e�V����/iK�vF�0MH=���.�Z)�RE���.�� �J���A�
ٱcD�+����u�T7A.��y�����Lڹ,�N�=�k�x�͉V�� +�))���fg/�igҶ���s���wL�\���4]��7o�申�Z���!.V�ӑ���{.ď��<�a�S�B>8����DJR��j�.���wab� "�'L׭!�\���2ܺ�M	%؞LW�qɭ.���z�cy�	{B]4&.�&�����[�z�*rP��)�o�V�Pk��F��źr�5]f��i���Ŧ�Y��EN"�>��M��W���w-�w�l��:�t	�$�H63�`�����[�bV����)A"����ږ��1q*�T�X�!FKV�e*�ZTm��Z��B�f+�-�V�l-kV�*�-,F�mjڅ���X�,Vѭ�F����-+b�F�T�����)YD�����*�Q�DKm��*�c\�ZF֥ERԵ�[V�"T�mF����A#R�آ��QTb*��m�1 ��D[RZm�i[eH��m����[ih6�6�ERУP��V�B�A��DX��Z��[V�-��¥-%T��c[�mŶ�R�DI�UE*��EF*��ґmik*6�
%�F+T�ZF��P��TZ$X"*�Ke*��(�b,Z61H[B�V���m�j�iDh�ҫmF��
���Ubň�0m��b",�B�б3����qv��.�d��8�d�9�:{�Ұ/�)���w��ZC�{����i֭Ij�p�wr��`u����*?��xx|��.x�?�����5"��]�z8������s	�6���Ǩ~��Rz�}d����Ǭ
���;��ǩ���5#�&<LI�;�> c�;�zZi!0 qP�{�����8,��ܯ�����*%C��|�g�1&�J�^��?yv��Ă�ٟa�&=eH���`u6ϙ.Y�=ܛ@�+:��u�X��<B���z�j��P_!��.���qp ��`D�տU���U�2u��}<f�+��򚴅t����q>M�ĕ�7CH,��P�t�Ag�_}�XT�Ax�Ͽa��6�$���^0����ý� u+
¦�y�c&�=J����y�P���k~��_������J�,I^�>ɴ�ܰ7�ށH���g�x[&3l���q?j������i'�~B���Aa�Y�Vm*Ag���u<a�6�����ǽ& �@g;o﬽7���E����������_,�=����m�d�ϲi��Ɉ�wX��
�VE5�`x����{h~v��d�S�O\g��ټ���N�?'̘��W�>�O�Fǀ� �D/�t�*�������}�ޜ?<LH/���#�'�3�d�|@�7�w�H-@��s^ ��TJ�߲OSl�i�!�CiR���1�c�\x�Rc�T�x\�8�����VƏ�O@��n��v���|�������Y��0*O��sz6ɵ}`Vy?}�H�|��{�CL�%zɿ���R����?'��I]���I�VT?&��&�4�Mڳ��$�����_���ַ����������?!�6�P�4��0����2�|��a��a��& u*x}�6�oܰ1��7�Ch)�l��wR,�&xw����%g�������i�����`T���$���o��u����;��{����ޞ�0*��P�q*Ag�fP�����1&���u>g��i�E�4�9IP*T4~�'Y�}�&2{���i:�z����kD� ��>�5'���w���y���z�yX�soK-�y@�=늏tx}Ɔ@��2q3ə��z�}O-��O�
��5CN�& n�gd��1��] u�==�ܡ����Y8���s6�Ԭ�u�'q���<0ް�F�+n ����R��&4}���ͫ���}���¢C/��4�BAfd�]����[1���|R�+ʖ���q��u�˙|Z�Y���<�+g)\���
���GM׮��H�9w�D��r�Ă*�Q��xݘ{xBľ���<��5E������@��1�ƾ�����ُY�&:eIþk@u+1��6[�M x��'��֯�
���i4�U��]��H�Rq�y-�f2W��S��Ă�������n�֚�ܷi�8�������@8ʆ�;�ĂΡ�3Z�=a�c�\k�c>C�� ���&%k
��V<f'�̘�ĺ��1�,g�٤4��~��~ɗ�M����Z��2�w� DDyǄ܉��%~�ȧ5d���:~�$�J�8�g����0*�����J�_{����gɈ{�Lk"�'L�I�E5-�i*J������]�<�۽׻�<��u�aY�9�i����W�i�&���g_̞� �X���18���>��Ch+��~w�<z��4�|5��&�0+<�sI��LI�;��VF�8�����z�S_i�s%�ݣ��k��0 ���T�s���a�S��٪� u+8��y����}N�����I��i��$Ǭ�{{�@�+=d��|��'�J�5ߵ'�^�*N{����~�E?�h�gm��%��cޘ�Q�|~��)�??:|�Y+�5hs�6�]0�1����a��M`T|ʚ�SI�~��1gX|��yf=a�f3�v�z �������:������6�Z�LTD 	��Y'��L@�w�B��5`g��HT��S�l�AH��5-8��HVi��i���OY_;�@�N3�!��|��`T�߲~v�f��5�ͯ�Aݜ����է�������OY�o��Ci�'�wZ���%@��k$�Փ>��i&!^�N�I�*��̞�AH�5�q4�d��{�8��������/�z�}5�����8:<��|]d(��1��s�M$FN�LC���u��O��5��������&~�����S�=��Oh��O��٤�H:�~I��=C��?}����UeF���;��t�@�B�LlxL :
�x��6Ɉ%{��:���g��d�J�U�����S�4��y�R+%w�sRg�� �g��a6�a��i2�+�Ag�����y_��u%u1�ḛ��c��}�U�����5�ҝs2�jҩ	WK���dFٮ��t���`s��u�B�����ۀynj�qTg����(�"�Km�v���}@ٝ���oi��_�֕��ܬS�Rfq�4��t�vl:��-� ���=���Ϛ�� \ �T
_�u���<-����1��]�f��!����I%f���i:�Ɍ<�d�m
��v�ߩ��B��]};�ہ�
E�;�j��Ԃc���
n�N��;M��ׇ��R_���O�q���8�Xz�>�*Md<t�g䬛5f3�8���᪤��T�)�����<�xi�A�%@��5��u���d�g;�2@��Á#N|��.�7�UE|��q��I�'}����M:AC�ϰ�䩌��|���hJ��%��4���9��ɤ��ۺAH��~LM�h�26�����Ă�MO�ï��r@��FLUT����{G5q��u� z�
z�N��	��Jϓ�w����@���~I��~C=9�i��I���H�x��3e����& s��gY7��|݇�VJ��ߴ� DD�����٫��V�{�u�ǎ�*N�_Y;�i �|�ް�u4���tM��*<9�jT=C�ć��֧P�Y�?&'7@ǌ1f'�x�����M&��P8�eׅǅ��{�����c�����#oz�~����k��m
���ç�6�HT4O)�y`b
E��u�Mr�����T'2ɹ�����I�{�涓�����0Xz�>J�g{��:�bn�&��"���������˯;���?����O� �M!Y�=��?��I�O̬���M�i*O���y���B�~}�i�̞�AO=�H*q�fs�c>d�J�5����=`T=��4�d�ǉ=9�{��y��s��������"2c�ܺH,񑴬<x�H.!�h~t����O&��Hq:��o �i���0���<J����COԘ����>�$��Lvw��H�bV_����<�瑩�}ȣ_{���=��R"G�{�S� ��3i*+%W��

E>L->�H,�nُ�O�M04ְ+�'ɤ���I��Aw�Ì�!�c'�9�L�
ŝa�0���n�����{��q�E�x(Q�
�}�o� �]0�]�A�x�"���y���*c�Lvw�"�B��{g��I*0�����Yq��q3�!S�ud���P�`T�6o���W�f*U;�^ˏ�FʼРn��z�<��R��s�T��_��V���-̝1��F�P�r�P0t\�4qF�-۴�RZ���XKΙQX�#G2F	a�sNmK�ޠ6��RJ���(픥�g�`R��7(m���r������{�	,Q;|�51��1��?{������%O��xé�<�|��x�_̞��mS�bA�;�R,���r�!��Leg9g���*T��J�+"��퀿>�x����T�s[�7︔+�� `t�틏S%@����2q1��Ϲ��6�ɉ�X����~�M$m��?=LH.9�'��wT1���CN�1�>�jB��D�,�+p��9)iܣ��Vz�r��Px( \	�}�z�ǾI��<3�
�_�����*R�����M�f�1>�%gY3.�l�rm'P�Y7�oK�
�S�a+㴂ʞ��!��'uM20�~~i��}]�n��;��π� 9�{� zꇬ�!�&�q�V�d��$�==�'m$���2,�t���/�)��ވ =��K����/�azl�˾��E�X��9�L���5`w�x�P8��|e�����Ǭ㤟���?�L�g�v{�1�0�c=M3i�������S�1���4�$G� ��>�������r���W��P:�����9�׿s��.�~�n�A�����l]*ߧ��2pױ�j��ȱCt�Ï����SWrh���/���]�8�vP�����]+�`���/�˞�M�n�}"��g��㩓�f��]��](q���zh|nL�
F�W�432*���1S|�f#��L�:�f
�O�m�hmtD�C���Se�~�ܹϡˋ�����sÛ=�9�F�+�9j�������`g;&��v�W��x�3�:��2�S>�s|�B�_���
UǶܚkMgL����dO9�b�$A�#T�c��s�xb|G�g��;�_n�xxܵQ@�s�:��*7��Y�Y�j߰�8�uY6:��ku��K̾� }K�����V�
�opT��;p�+�W�v:���d��G/���=�ҫkm�kW\����j�L�@� ��w,�q6�5�:s��f�*����.w't��^�yK�6
һ>�)'b����E#t).�Vl�
o!��?,|�]mǞl�ᱻ,�*�v
��f9�Pf`c��*�h��l�D5뾙���x'9ä]��Mr��.������z�X��Ɔ�<.����"O�բEUG��Ѫ���S����$u��]>�%�z'CN�w�R�!�'��R+K�����W�x�I8�s���y�^��a	2� ���(E��_4zfJ��]�G)Iz��Ot�^�i���z�j`�+%�t;_���h���\)�n(+��s�:��n�DfsF>͂���sc�������������@�����k�pO��Xv`�y�����Rdg�`;ю����\��w,F�Snɝ�X��(��,N����R�V�|��n�p�u���$OO���{�w�a�L�X�s���7���E4�iG'm�+a��kuX��B���[a�w���#���$y�ϭy���&�t�,�D�7��i���SU�/ǖ�za�X�OL�	��|�����*D�y��c�xyWrќ�,���9q26�iCWs�oJ���S7/B��o;k�w
0�5��[�˪�eQ%b��l�O���<<=��Ҷ�c`��O}�f��wcc��k�w��p��]���}b.�F�Ľ�C�����;w�%�T��N�A�bF2慠镳�s#ϧL���;E.X�.��}ͽ�y/tG3F���j��|�U6�֫��V��8wp�/p<ߏ��I�����+��N����Ss���bxϻ�⢧�]�d������?mZ�6Hix�E�Y\�R�J7�\����P���I<��k�9VaRi<
{{P���.���
M�n`�S ��Y��k�Ŋ��`]�zy]��۸7���%���lz����yV���*�ݙ�y$��!b��˹�;��:^��lK6���l�"����}Z�w�^��lA�^����o�j��d�v��>N�ݎ�5*0S\�r�%��+b7\7�H�f9l>��T;���C'��wR:���7��m^Y�)�˿�V�2�S*M����I��J��Њ��/�+CS�;!�r�B�����kS{C���gNk=�r�{�g�jj^{��J��d�;a�軳h��J�����5L��]��l�*�����2�+�n�R��=j���Yk8��s�Uk�X؞�KQ��	�'za^�]]�GM����۴RS��?f��T|�D�l{�����۸>�6��p�h	
%�W��j/���V���v�*ÐTm���G�Gfw�5��YY�&uk�k��T���,$�;V�vpqbU�6�[�P��V'j]Xv��~9T&��ēq���烌F��ҞkK�T��f�[��Wa��6w��,�:�+s�Mȵp�j֮���O>K��U=�VK�⠫vލ������'��$�V��jv�ǹ�髨Q�iyN�H���Q�l�[Wro^�s{�V�yoV���<��u+���M�6��w�[i��rJvH����+m�V�Oo`m�3� �s�����]����u�f'雌�yX�66z��߳�)�IXUܳ�{{ �4��	�Y}�7�����Ϛ-.��w&(s3|��g]���Y��1s�2���H��-�bQ�=f�U|����=e:��F�	�9N9K/k�����h.;-�w�\���^w\�&B��`Sl����ov�m^�G��%Z��&��ĭUz��+�����r������vJ�-*��]�T$��ޓ��^�/�����0�ŋd3���φO��q���`��	�߷�'Jv�3�qr�[]s�𵋰ڋe�:2�O���"�Q�K��ד!}'d��-���ڻT��%��oJ�0�3�8%_��w�͉(���3�W�3E*-g#��u�.�y�xӧ������t[�G�~Qkѥ}Yޜ.�z���jL�y���c��Dr}6)�YI[�+]F:b�^sj6�ݡ�Ӫ��{�d��	��o1�$�p�N)6���h:�v�Ԡ�d�m>�m�H������A��;�)c�Ŷ�+�.�%15��v���uW��n�n5��xm�r�ٚK�Ծ��Y{Άի=Lާ��2���.�H��]��;L�&{���NP�WX;��N�xwX��F���<Y�3��X� �X�K���ո�MT�y(˔ѳ���r��:#k�,׽٩��#���ǘq����bIu���xn�B&�����1����y9N�vf�^G�o��>�dv���D4y�s�]�ݷ�zo���� 咯�O����*�s��z���2���&[����X�o+�\��/Vu�fy���P��k�,�ǄH�b�i����{�����'l+��v)�O�U��ґ���i��~�$g ys�
�x^��܊2A�L�m�����]�`.��_p��oL��+9���j{�>��@櫕I�쵯Wy��wK��������.�s-i�oT�݊�[9����pmaIAňd12Y�8��7t���V��Rq�꽎�+ǥ����K ���}�a���X�v?%bxL- �-��K;sN��	u��4��w�d��nlK6��K���,��b�E�[���}W���Ǫ�);�ڼ�)�p����l'op	u�>/zGQ�f]#���#��w}폽E�H�f�<̄��yquc��y�׻A����z��ܔ�<�ɧ�j���F>�8(V �#i޽֑�[>U��ռ���`dۥ�x�3E'��
gw[�%_}�������
��nu
O�S� 9���
S6�絆0_,����(����G��+p�7qf��2'�a	u�Կx  ����ӹ�2����S�OT5�(Є]X��`n-�p�q7V'Vt*�뚼k1E�-ec���/���q�bm��>i���yj��>�;6���R��Mzws���7��	�-!��pX}�-[� ��w,f�frV.�&b�I����}��մ�s1�*��n��(F�VNԪ{՚e�WwE���}�e�槕��#o[�m}T��|�K��-4MV4`�7O9]M�x�vQ��G�G&��q3�v���5e�ꢰuR/SƳϞf�OGb��f��D�K�G��`ߔ��D�&Pg�	�B���So���.�񭚮'Jxo��V"��6�2�J�R��Hw_���'x�"u�R�--��2�w7�ջ�8q$e�8���r�T�X�i]�	0��[o�I@�������t��{/N71���cO\��ap_��������J�V�����R_!�p��6�*[q�P��Us;�-6�������pa�Rr⫏��{�y�t.�Vt�,C�l*�t��ԧ����lKܭ��{���8#���������C���&N�n4͋ gx}����P�c����!]��$��Y�6F��Ζ.�6�.�|���z�%]�,uY/,�GM�
���=+�CJ�u�6�r1�^]t��6L6�|G2n�GLrĳc3��9�j��b�#��w,�Y�D�H��X�cN���6��v��21�G@���<�&�J�8�I�t�8��u��Y{.����)���ӝRf�|^��g	�_jB����~���|2��Ɛ��b��M'RU�G�!��+�73�F�鹍1v6l@����m���V�z���5�����뀥b������<.�l�X�B�Q�Dh�A�M�87��{�PuɁ�V���[��;kt������-+�����Ա�D±�[��M��U�d9��EF%fIWW8�ʹ���D���О�J�e�k]㎎D8��j����Y������ó-��@��ij.K.�ԭO@���%W@֜�m�-ܝK�Ms���{1��#�t�B8��Bl�J��Y�MٝK"�u\B��x;�#k��Kr8��z�U�t�ʉQ�bo�mp�ץ�ުd���Z�yw9@�V�m�U:8ѣx��Q�x�q�:�O���^��p�:(�$�{$)�pp:q �'x�K�-hU��庵��Ƌ�C5�0�y1L��;l�;�:�0ۼ�*.�b�C~��z�H��Vn�Žݪ�9fd9N���m�;�,w�y3��/O
Ֆ1��7%
�Y�Q@:oj�D<ʵ�.k��AR�J7�ۮ�\3$K֥^7N��z��\[}/�e��B'k{��TAֻh��s�~���4�*�\��[k� �]�zY}�rl���7]]���c3:i��.��{�F�1�����be���<��5=���.�v�͕x�!f�M��{aCH�a��\�ׂ}{�A�e1[-��HKYc.T��d��kbl��젦���N�p��#F���HT�)��P	E�n�M��fV�����*��c(_>���q��y�Or���l��-H9:��A�qg�rݺ�s�͍"p�������f��Vat�Hh"V�����)��V�yE�y@�!�B�ivs)�[zG.�Q���j��,����{�V��o7�6�u�uɡ��8*;w��Wt/�f�;A��O��j4���K�y����8V�7��w�tQVw�b�F{T{f�	<������b��<�-i%1��m��uã�k��=E�F�M_^�$5��s��7@Ѹ�1�����+hs\l
�F�����]����CK�m���KX��컁>������
� ���u���lK|,H�B�2[Qhն���b���U��+m��TJ*",F"��TP`��h��Je�H��( �
%E�Ԩ��A�m*2[EX�X��-iZ���PBңJ�T���R�Q(T��4�F���%X����U�T�����*�+mc`#U��Tj6�֬����TX�"��Db��Qb���ƅR��bZYmX�*�TR%���m�V�DA`���E��elEUX�VUJ�+Kh[j�"��+H�ڪ�h�b���
�F,��T-�R�E���TV���[am�UQ�,UUm*��Z�"6أi%��,b��*�@PD�F*�X��h6��Qb,Q[K
ZhT�
�ڠ�*�V�Ab"�DUV-���1UTDF*��"T�,PD`��"Dz L�)��f*�h,9��Es����W��7�sNt��\��b�F�6sp��"����j�� �Rٵ}j��'�Wb�֞�,�
�����}Y��۸7��Z�o�汱׏�ג<K�Gk�������ȟ¡�b���swr"t�վs~�mH+�{r[x�`��;|Zκ^/r�H�X���D�f�<��а���_cɝ�_YX�:������}��0bK1���r.�<3aP�/��U�C⮞f���j��w�,�؉��[�^�zx�OjEGU��,���o�������ۯs�0d#����X�b��/��x4���~�@{����T�>W��V;���j�6)�1E���L��Y~�����Fp�r_q2I��xk�s��[^V��Xua�Ц�䩢e��iZ��:���<m�Y5bv#v�'ʸ���EX��89|;���z������(嚴o���Y2�E��r��8�잴�����/ެ���.�`�M��9G��tN�xLX#^�Yc�
x���z#J�q�]X��X_\X�|A�g%�\s��y�5
���3������Q�} �On��uo��g�<�.K:��%ϖ��V���c�1�1j�ds2�_2�����j�v�D�;*V.Շ�J�<=�U-���%����Mc/-���y�����7��YF�H>�Dq���\v�gr����EM�ªi�uk�&��e*��,D�b�rқ��:p�	��KK�v�l�~�|��� �c�=���'(���h?_ r���,�K����+�;��3���e��mw>k���=}\�׳�̫�S���D�� 994R���տg������:x���A��e"��~�6���G��}ۂw��ʡђ�zJ[�C��Q���W�sն5���i66?%�G�����F����\��9Wx����m�[��Й7��ܳo��ߛ�0�jJ"7%��0D�]-g��;k#�.��0K�Tȥd�^N�x��SrZ�˼����e���O,<j�4®%����a�C]8���X��7�{��������$"mҨ�͡�Nν���/s�,�awM�#kw��`�Y�d�a�[�0�.}�f��n����_���w&뜑���@���u�mٚ�;�yD��.�����%CH�]Z��Ș]�֝]k=��DD����<=�V�d��*.�F��v�
���5��u����+��,�%�eL~�}��-��:�c;\ܫ�� �K;�K��k���.Q}K�2�By�j�}���~��x����f��5��j_nʸ��{4�i���poZ��[��d��H)�i����d�茠�g�����)dj����Y�5]���]�}�2�OZ��_&^[�&�f�=87��&/�A%�l�sRj߫;�'��]2��x�y�;��'̈́����%�,�]�f�ܶ��Om�u�H>�Bs�<��y[o^�/��}z�4zi�5z�4_y��n2h/��b���xg�(�]ow;
�<�3�ow�����Z�������2E���J6�urʩ��n]��o��(;XG?&���l϶=`cd��9Ɓ�����~Q~�Z�9�kB�
�?3�P離�G-�{��Z��;Ψzfb"�\`x�<W�O���D���-�>�1���>�(���|��\�Iُ�����U�/2�"�����Mv�!�A�-�1C��p�ôS�\�lt����k� �Ϊί��{���t+g�f�V�˓����վ����l;����0��+,�M��.�z�)o'{���"�w�ډ���NL�kz%����.E���ݹ٥um4y��!2dv��)�d--��S��%�=yyBY�W\��J��\R���v*�/�H����XN��
�W��<���F��q7W�6��7�[�i��.�#�x?Jڝ����ay�os�ʳR�P��r�A���?byf�8O���'R�q�V�����~�ϩ��n-�� �Mė4"M�7o�o.�3�����I�'�!O�pX}�4���.$-'��ʶ��z�߽��3�L�=J,ڷg��,:OmU�Р�ݜ���s�Ⱦ�5uL��7g�x��^I������W�[���zS�z��h���M�cVaN�k��v��u���]�����cP�c.�U�+_'�XF��1��i���X��/���V�ѥ�o�*�:VwEk����囱|�,�\7&�Ar���V�]]\��2�]ڙ�^�,oy�1��;-�2��F��ج�],���>A�}��|:�l�{�"Q�\�1uN�
�gL���IQ�X�.�������G�':o�s�yG�÷Dr>hؤ^�#��P<���8��lt�QsYt�梎gf���k{L3�_o���ۃ�uH�g��l�r����)4/2Ϯw{��[�O+$�)�g��I�0	�����.�\���8������s�1��g8N���4�y���cOI	��2��z��s=���t���b��ԥD������x��W����no�ew��W��E<�T�8.��yn�1��8����"��c��5̣I1�Du�^J�t�Z(ANG"}���$Gai��9m�nE�+����͕�����s�M�7�:}�.~�buf������"��U��q��1��̖>r�\������xk�Q����Nr���I�z��b���
�&��y�y�l5�{��t_��7����K|�ؐ�e�2�U\��� �QL(� ٸ:��*]h����dś5Y�J6J������:�a�0�G,؄m2��ښ���*�d��p ��vp�е,]f����
�F�`CCo��wRwBP,�2�/n�3�Y��EI�3Qި[�[D���  �r��K;�Λ�����z�wu�j�&�4���ڭ�r ��&S�����1���v:��wsԱ�n�#δ���T��51�i9:&�ԍ�˖d�c̛s��w}/ʸ��t6��w�����3���ِ{iԫ����k�M1����9�2����7U�Q�\�oڄ�H7&.Ț��y9��j�M���qI��yowg[�ҧ�,�VeA��v������Y�zu.���Q^�%�U$�:�؛:kϘf��������G���$퓱�ͶKuu�
`�J������+m�t�ǄS��
q�	y|���8=����?D�~�=t�V�Vs���K���k��ԙ�N�:���7��nf�h�
9�ԛ��F��c�ќ;wx6Fܪ�NWu`�٩�h�K��e�f��ؼ�zxO�h_w?���oQ�ɉ�W�2�Ƞݿ�#��S:�tg-�7����9����^�`��F�yDR�N9��U.j8��1�'�Χ�莊��[$��b���|6�K�V|���v+��v�x��9��+��1d�Fn�uvv���Qg�6���ʸ�J�{� �N���2o�w��kֹ�3H�6?%�:ah�<�P�BAƜ�}�7{H��+�f�J~�ւ���'92ͼS�U�����C������eV�%�ح��Vv}�;�8�3#�3�VL��Ӣ�[�N�f�+�Է��kӛ�7zaW��a��Ͷ�\DLu�c�L�9�&�2�%)�bMCy�P�Պooqm�z���uc�8�M�{TC����l��Ve_fg��M�4o�Mjӳ; >�Q�s���yo�7�Xwt2���p���x��݋���&����%�L�o��=9�����=˃);�������ˆ����
a�uoxPmn�y�F8�ᙡ<�O�El�t��8=�}0��_U=����}M`e凼MV�sӕ�d��i�d��f�F�gO�i�wGX�$b1^�XU"ӷ̭�D=�.�x�%��&k�[���*��w0
�A�Y�a��z�)�d��,'�x}O����ۇvga��a��ŝي�mNc��R
��w�������U�3�]1�&�{Yę��n[�]��we�<���f�.�ta6����,lƗnU�\v�P�ˮ�D9B�z��^ė�ڲ��ilWއ�~+�������`kg1�}���k�[��S۪�Tx��e�z���(��>{Ju���3�ќ�X�,�/�:B�����u>}�Z�2��{{5#)ۈ7��9`�s=�~�6���'T��~Bb��qe��ְ�&��=�=�lv%�	C�2���ES�1nߊg�����9�{S�f�v�X�����[�ca���	�@�R֠���uZ�y���`B.�F�X=Ďź�d�;s�O������J�k�췼w�^T��:*7������vz���oOml�ԙ��䵹��ƕ�#pG[W��C3S���!i�H{��pn��U��JԳ��s�
�q����T%�(Є]K��Y����t����Y��X��|3d5a�+����`ߣحu��iy�w)�|W�Vm�?I�����N[(bg�b�A%H��-��ֆ.l�8�AޟlJ���+o�6��k��]3���f´��#��V�[�����]'��zz�O��,����=���\�]Gk{�����n�ѡ��V�
iyvr��ZU������Q��&]��tyG����ewV./���?eb⪈�AՀ�M!����@g����Z�5�XG����gs������ڵ`�3��ëmRh�ݜ}�:&⳪8$su��6��G��k��)�m�N��+�V�[��`My�j��?{�E�Q�Zn3no��|����׼ ;V�����?_U�T��ۊ{�0cr'�wM�_,9��/�No�F��܉�th�����#9	�k�Ot�oaImɽ~U��7�ob(�ś
��� �/�R�6im���6g�ٴV�%V�aK���O&|�od��`!4w����-�O���Y�s���z��g�{9ց��:�6N705�٬i��HLx�����*�g9�׬�m`�_O:ݙ��JTK7��]�m���ؖ]��Ok�.{���FE�����-+<�]Ȏ;� �'@���N�a�Xk1B%��]�]M{}�4�פli�+SVb��!l�*���/{"��^���`y�қ��om#��ԯ9X6����-Nؖ��p��j�QC�����{�̾����7�Z��Y7�wSIX���W�� =�n�=�I�K���ꪫ2v�$/�����u��z!���H��-�Ohr9�΄����9�]�nwz`bo�S��(s >ݱ�⿂�����FNr�R�^X}�o3�5T�)"��X��P�y��8�3#��E��^�u��cnwJ�Y��81��X�1�pav�7�&������� �N[u:-�ss����zF��Sr�µ���Z��Rø�ƽ}�U؃�H.�Y��j[�p��h�5��st�ٖ3r�A��w,g +kj��Zx����Ux2��w$��������N�vE��j]a���ݡ+�,���@mߧ����D�>܉�ڮ��V�X8��J��{,6��2r�Z���k�WC�5�-'�T�g���{`�Za]ފv�Ɂ˽�{<�̼��vwf
��˅eO*6�FNR�L����Qc0c�F(�+:�'��v �;�2��y�Y�=/y��NLL�ʛ&�+;sد����rȤjXV'�z�7mUJ4h���/[}[���w��]����*�P��q��TV��-�iw]EС� Q�ۣ�D4]�W�Z,��ܔj�T*�x*�P[-�
x�׀ҫtK��Vw6�އ����Mk�F�f\�]jfܽ��X��������r\��	W��`JJ���Հ�4�ʲr�׺+9q�V>�<5u�{o)l'��ݮ�23\��5�4�5�.�	����&m�l��|����f4/n��HW;]v^ �M�{��(�Jb�<��}Y�V�멬j��TԽ�m6yخ�k]Zg��f\�!�(Y��T�˭��Ï�C��A!�&q!�`�^m���v����;�	�{�f,�we�l��4�iq��d�U�V�¶�h�u�0�)n*$�l���s1h�5��9SW�60�2�1
��y4&�YhK���]9��Ӯ��܇_j��GOd���뙴��3��\Ժ�M�
�ɬ�X�
G�m�&�y5;�ֺ�1��D�[��R ʹ�:9@�i� ��ee-4UW2��;�����'-����P��f8)���os�y9٤��G�Ye�<���b�����f�]�(\���C+�J�Ls�(��%�:b�Ovq�����O�:#M��Uu��s�K���d��:�X. ���*�%&����
��4;Q᥮�X��2��w\�2iyO<��n�p�IO�_���ϰU�d��,�X£sv�9�-�u�l�9�@���'�.>�Sɳ�@��J����L+8tZ���G�Vef�-dȢi�{���Kږ,vt�+]m�F)�Z�W*
�j��	N�Zb�i����r�����!��9�����U�+E)��Yǰf4��Y����F�o�r����6g?[��#�r�㉕T(�z�ӵsp���v)��&/fS��®!��cv"b*��x�]"�<��YU�Lk.U�ܮ�\��R�8pĜ�1�W� Ɖ2��Qd�u��t�<�]�,�Jp�B����u@���VS�1���ҟ<Z�ҋ�;X�����+��&�c1�1i	i�㣦0��)X�$:�'����Eej��Um���SL�����`���w8`��K�Fn�}�OJ�����й�κ}�Yj��J�~�pg=��n�?�;�S*,�-,�� �5�ut�����;F*��-eDV�;B��-]���� ��v�]܊9�V�I��e��G��M��r�oP���ī5�-'�R��:�s˳+G]q[vӗt�Cٔ�W�]����;��m�mpJ�M��N���W\;K���0���R�h�͂��0:!���C����o���U+OZ��\E����X��Z���?���2#!'�;����8/�f\ٝw8����˝��C9��,P��6r���l*� �� *ŅeF
��PATU5,DV$Pb���֭b�2"kY�����V��hƉEb�d��Zʨ��V(TEUŋ*�E��""��"�#-�X��*�PF("�*V�*��-���EEF"E��(�PU�5�j��Ȳ�U+�

��īj���E
+E�*�U-���(,*UKh����T��h�X
*1Ub*��,�TF-��V�l���X�bȪ��kZYV(�EUdU�+TV,Q����AJ����cZ�X��
�"%�V-����F�D�(�iAkX���cm�cYB�PEUb+Q�J����UUQe�*��Qm+�
���m
�Z[hV(��Ĭ�++
���[d�P�,�V���("T�V)`��)VڣKh��*TF��B���Q� ���TG�|@�@�93�P�j��Ἲ�y����Ip�],�k������!v�Ŏ�t�c)�^>�2��ӽ��G1c�*sB�H��{���g��nrd�/¶����m*�B�r�*�nz�A������a��k
�T��IL@����N�L7���.��e�ۿ�w:���Vj�h���]H��Yk^���q�9��&�R���1�����8�i��2�ҹ�m�b��q��kx��p�4!������>�x�ݳ�ӯ7�gicO>���|�ĳkca߱�+���-�uV&�5�������Yw-�`����si58%7���;]�<��%XޗK�+'�R�);�5���>��C^������.���9z�k�S)v���gyv�+�b���abw�{�u~��l4f�eVkB�1�D��'p�eW����=P�E�v����*��mI76.��;k�*Ԛ����w����}���)q�ֹ�*��A�gs~]<�u��N� 㛀�w�Xy�:M76��X_vNUnxVTO>�[���,(��[w6)"���KzW\s�`��t
�i����O���A��R=��k�p��r5�QŐ��΄��o:՗�s�!v�w]uo�f�=�l!1�S�Ğ�tn-iU(����<W�G�s��W�PuoP��|f�홠�5�L>ܚY�q�kFu����Z�C�W������uO��#�[��r�=@�b�I*�M-��{�O+�nF���]2�O[��7��;�H6`�H'�
�kk���#sN;hM��PH�ɇ�̭m<k |Ν�S���̖�Z�o�EF1�c�`��)U	A�8a�y��Tۭ���37׎d_Y��V�����`�'@B�V���)��^����j�d/��:r9-�}��-�}��;qe!S�uM$g\T��je��Md��~�Vj�I�
{o؆A�҈V'��΍�9��һ��*ܽ�7�<�X�V�z�K�R'���tߛ�z�A��j/��q�Nn�7ܔ.�Gi�`e��I��KyL�rͫ31�㈸~�t��d��?s�Rћ������)���H���v�h��»����WP�6(݄ƣ�fU�=���t��ۼ���YX�,�uP�ذ�����e������JC.�pܛ�+�Z��Eµ������U��B�}�=��\m�ڱ=������X(z7�����*��{��>�g3R��o��[�w>;3��˒̙����Ok���l*<Y�;x�1Q���c�Uf�ſF���,y���3�	`�5���p��Fp����L��)ֽ[��ܐP��X����=��	�!绯}��Fd�i]̣m]�rsy�̡�:�&]X�J���P���w��Q��˭7=�ۼz	3�<ࡳ}Y�3N$3K{Ë�=�I�|YS�����QX�����^���L����ry�b9�[G�e�ϞiצG	�J�!�f���]�Ϲ�U���������8��M�Vj���;�bi��R7��ͬ�e5l���vw0l9�#y]6)�²���W��S��;��ؕy9�s5�q��2�W6��P�O{ӕИձ��E�#	r7�ƎK�ګ*�ֽF;�����]��z2�s�	݊"㷐;3���~{��G�(b쬊x�z����&:|�������;��Id+�E��$;�S�s�U��p]�-�Գ-��NJP�r���uf���z`�ī��3�w���x�j�L�2���(׳�����&ەmAlͅj"�#��MT�$�|�[�h��7n�����hΗc9�+���of���Լ�N/es��� 7=R�b���c��TH��v}�%�^���3�6�uN0��WROچü^J��	��`T�y��Nst�kF�77���I������k�v1�+:D-��m�*w�P�P�z&�ɽD󍵖�n&�bt�f�X!Xl7p:alВ�`���ԅ��r�>*H�VR��l�Β��/��ܼ�+&�+N�x�9�⋨�έ�ͷ��v\��xՍ0w]i���6)��npkX�&%�f��Fj��$�]�o�*J;by�Z�ת�w]_ku~M�6�,�!䕛���`�s{;�k���C}p��K;�K�̚Z]o(:�=t!x)v�x9�\�Xn���C24s낅�v�D�B����
�z�9[��2�+�X��+���A���T�[�O�_�*F��N��%+{�p���܎�;;�ι��vN��y@���\k{7r�0gV357��$mN��<��rp��5}F���VS���@O^�i`��k8�ߩOb�kM��$y�h��Fue����?���y��>9�6���ą^�g+�	���ܞ����N����1*�oê���^�M`e�������
L������=�����w93n����1^4���O N�g�l�2��6^#�Č	�����qB�,
��LN��g1^��c�$J�>޵Vwf��\�w]��+�J~�PD�¡3�+�u�������Myk�iVL}Һ��S{>ק�HM�P9���u��L��o��-ڞ��:b8���}��Ǆ*��y�k��lu�	\�B��#|*�qG������wМ����3��6i��v1�+�z6�}��,�y�U��w��/'�#w�YQ�N�L�&�ۛ��w������j�Ii�˝����lݜ�++#~�%kk�M�X���x��ojW�J�\�YU�k�ƅ��*����9��|��;Y�{�\ |����go>���H�+J�l�i��R�s:5@�w;��Z#�"K2��i�}�n�Y���˳R�ݘh�^�.�mC&�vм��S����'oaͺV�s�FU�e�wS�Β�}1��!����N�aQ���l�NG�үhIx�w��Ӄq^�}8�:�й���k�n�[��-�h3�ݰ@��x�o�7<������P,Ƌ���z��z��e����ql���ܾ�0%a��E>�G���a�y4%4�Ѐ��Cm��JWƱ�r���ܯ3�r�o�.b����[�]]��fΕ@>�V�-d�9�QU+��w_d���Y**�~���5�2�uR���|��;z���Tr��6&�"�Փ��.<�اᲧ,F�u�MA���V�E�x�i��WX|K3fo]o������[�	V'�=2�r����,���f�m�U��U��n����킻{(����>�ٵa�A�%��aL�T�a�<�-d{����:n��K����] r.ƥfs5y2���F��LN݆>�;��v@�z6��br�;B��V���2�.�ˉ\�o�Ⱥiw{)�[؞��ػ�>�e���뮳}G5�9+s�v��9YjY}]\�MbIn��ܦ�
���9��:NÁ�e`EB���T�"�v��$�U���%�!qu��k��BʎU�>	��Om�C ��}�ᵎ�B����ֻ̧VvfnMh�bW9�H��.w�"pj���-�<��!��,JQ.{�M�<���Vվw\���I��N����skk1��<��{r¹�i&�=c���`���A�~�U�/�!ik����7��'v��������6ȅ����h��=�~��iv"x�`;F�R�vsmy=�6B���W�Jم�VQl/����^v])Q�;����z_�-,f¯"n�8{� �,�)h�"�˄�4J���A�r��,�S'/�_}�72�}�Y.��PunAQ�_N��G�t����vJ7W~�d�k6.؎�g3,g[Cj�Kg%_�m���GO7M�������ULlon��ڤ�Yx��}��c���R���x2��\i�MO���mzU`�kc�qA�}X����{�EK�;�88J\��j���mc�C��Lt�`W�n��y5qf=}��8��n�>4��F���.�UBc�;���OBu׌:����y�y���Z�u�z�n=uViƪ[㝽�v,�ҹ����Ou�%�TZ���7:}\�	�q�zOPwk\�b�;<�ܛ�6��ЛV������h��=�#yX�FP}V����H[Ϋ��O[�(:�<�}2�@:�؛/VN�c�Gf_�N5�c���q7Vs��]d��'��b���rm��s�{�O+v��}1�9ś�kN<�w���}�P��/u��ޮ��y̹O�� �O��R���jU)ͩ�Y�-l3w�&o���L�c뱼;w7����U�W%�e�Sǰ�k��^��i��n�������K�*�}�����t�e��:�9ۺ���\�ĳi��o���:ao���QW�}#���N�<յǑ�R�����Ov�v��yr	8�E������o)�0��^���w��{�>��̢���p �J�v���E��3*q�_s�U����Nw;���|��qi6mF��y��F�u-ҟki(��@�S�'w�av]��	j��,`n(:�S�w;_ZL�H{wavR��m��|�� r�䬙�x"��ǲ�Ĝ��qw����� ������w]_���A_G�$X�_��]n��e�nR9s0��Q��yc1m�z���uc�J� ny��c'/�˩�+�cF�,[	T>DK;���YYV��]������#�]mV��^�uy��HS�o�z�Q7��gZ��]q�=�;E�ݮ��kZ]��������y����6��o��W�
缞��9^�I�G���y���!#w�N�S/S�����5�����T��.䉖�Փ�7K}��9<��j1�L��M:��M�el�]=Ⱥ9J��y%�LE؂���lW��9
<��m�t��i�̰�{o���F4���vCV; ��xR��s-�$��0�o����N��5�6�Vy�;��pF�յ��y�D�Z�t�:V���k�8�R4#�?���yb<������%�a7݉z	.w=�V4S�ծ����8A�:�>�n�{wQ[�ۘ���P�Ag:����Ŭ"�\�n9�ړ��X�>�Y��w]���YVgo�&P��qyڞ�m�*hYo��E��熰�>�s��X��� ��Oq��lhb�ᵄ�7ݲ��b�\�?O%�y��,m[�6����c�V]�6o�t�IV�Խν�|���G��r;;��6;s�;��1WL�я/(�ӥ2���1�B7C��#�}���;N��l(u���+�{��<mX��T5������:̈́x�<�C+��f�'dFq��y���l�f��k!�y��x��*�9�7�ƴ��ܘ�vߩ�Z�V�mZ{S6CV�#j�<t\{��gg��Anb�xu;9|�[��KT&y���Bx�폶�j�ɡ4��o_l���A;wQ�*�Ωh��}zJ���*�oR��j�S9�,;iU��Skv_d�P��A��܋�!�{dҸCo�TV,�B
�{4)e�Ӝ6� N�gXsN�5�{���Ž+�gQ�_H��i�t���}}��Pf�Fs�1���98��co�;���s��F�j�֦���Z�Yy}}v�6�s{����3l7B�
d`�nu�ޜ�I���;�[2*�������NG]��yk�k���˝�Lɚ�T�LKh�w6��_U���{/���(�ƭb�c��TD���S�VsY���)�B��d���d��"�i��[.���f�x��z�Eucj'�a��|O2oI��ԋ{�]��"�H̏��ɦc������(��Z{�֒9d��eB+����Uh�ʕ��[�����@bH�(�܁�����Y}��6Z�I��E����E�c�Q���LW�������_��$)�i'[k�d�e���PÝۼl��o�i�֟�)p�աַj�!\�,+�w�K��֎Z\�N6�U���ɚ\��m�f��٫��n��^*gR�M,���(KX����˺8��p]ӵ;��-Grǝn��D����zL��v=Hn�ӛ��0�˽�nM �������<���qҲ�gE
w��u�� �u�\(�rL�h��\ �تA��G�^W�0���b��Q���Spv��Yptl�uf�%�Bh+Jk/�AI�!�h���U���[Z���:c�6���)�f�*MR=�|+E�J�B
�ӵ���,6�]$4�fֺ��̗��LC}�ދr��k�m�s���k
�wV*��jD�8��W�j�\����IK����eT���}	����[��0���Z�v^k2�@T˰KU�_#��.�^�8�[#�[��/���d���b�0�e=44!�Q�Z�����u��*�m&%������;�c@:f̢u�Y;2�����P�pE��M��䋜7ML�9N�oR�hQM�%�X� ���u]��1���ZK���GHq�W�Mö��3�m�yN�)�ɨ��љj���6R�����E�6�4W7#8��b��W�kD�}�1�L���Tcr��KB��T�q#)]㏑}�*	ۼ"=�z�#G��£G���R��y�w�^K�� +;9f����.���/9A+kv :v<45�+��A�Ҧ{e�L �ҥY�se�o5d�)��=�z��2ph޾� ee+�}������V�]�����{t�EV�u��2��zs N�i:�xV��.�2�i��Pv�;���f'LI��� Va���uh��bY��+��;���8��������?L���--'Cԋ�I3SF)��oi쌮��Pܤ��ة[�T1��	�
��s��B�(�:-�T��ά��]$9C��܃J����w.�L90)s��Y���@7���o�n�*48��A��r�ݎ��^��/��wy�����v�a�Et]~�Mh�G� ZQ�K[H����(�YYY+EV*��FJ�k-��VQmڪ(*,�X�[m���(�5�,R-h�+کP��XĶ�Ub���֪�(��i@���4j�X�*��V�-���Z²5��(��,�UQEV�ʔdQ���+�VʤEQR#U*��`ҋ*ҔJ ��ȱE#�T-),b�5�TUT�
2��PUkVKj�[
"�T�Kmm�R�V,%aV2��b��QU
"�Q,B�YPDjTU�-��,b��TB%mdFT��"1Ac��*U���*ȥE�FҢ"���QF[U-�X �b��`�(,� ���E
�2�X��Tm���+i*T**�������Ȋֈ(�m��X(�(�����V �Uj�T�UR5��UR�b�A����"�D(������b��҂>� ��Ɋ���toFV�v�$�s)֋島���f��n0�daK�';�'��;Bi����tWq/�jQ��r6|J���Gs��>���Fީʱ�Kp��o���^LJ�/OTZ��~}Ϛ=�yZ��mvU�<���'��,��]b���KJ����3�~�̓ԟ�?sV��+��xD�(� Ό�>�޾���²�qY<�ܛ/k��W��9ol��XB��D�u/����@�9�ʙ�yI$h�[�Ʉ���9���d��˄�����<���'y���O.��z�+�|��e3������J�bP7�,��'�P��V�L�AT���q}��z_�̋����x�Nj������[�S�Z�d�)�X.�r�$H���>v+���"q#�n�z�*�{rsdp��i%K��h�cӮ�x5�]�� Ȏ�Q��F�j�G�+Vo�������e���ȨNC�����3�0���K2a���ٶ�;l��.�w3/ʷ</Q豙�����3=�P���"f2���siɗ��l�:}��#��v ]B��/��"B�ʉ��3o s�;&읉[.4��}���Jz��p�s9�^�JkI����5#�aB��q�%���Ȑ�T�Y*LKd�[��,s�f1�J�J���Qoz�.�ΆD���pe�ͧ�7���E�0�w�u~��G�$K��#�u�U� ��Ӕa��oy-b�{��ݻ�b�d���Aզ�4�y�t�7�Ӷ�!y�R�K�ݤ�e�܆��G����+kj�Kg=ŇV�U�S�ճ״�k���_Z]����|�K�;9c:Vӛ3<����G}��]����>P�>S;,-��5X��L����6+�P�ep��i]b�Ī{�f��J�c*���L�	�l���vw h����S�{��������ٌ�7ǄH�'�K+=�I=�v&͇�gqf�X��ݍ5E4��r�b��D�9����[��(g'ɷ�:X�)��m�y���{b�dݪ���&~���t�X����Ηy̹X6:���C��x+R�8wy=6�'��
�j��⻳�:S\���57�Owu$����!�ؖ&�gn�O��[��Hd.I͠8a��p�;�^�v�&����2DX�� ń{6�U\�JR/g\t�<��m��~��ֺ	7Q.��@L���8,f�}R���<��[����PD���S�0����5J��k����}&�t�ia}9��0����p#;�R�L�_��ܾ�K	-�+id�Lm�si �ü~J�#�B�B�r.u�E?r���[*�=<P�g^7�o�=�ݴ��3L�X![a�:��;-�\͎F��S��g%�<��|/#�ķ�	�0퐝��z2pٻՍ���m,�u>څo���Fj^光�u��ᆃt��Y8�Z��Տx$���eA�;؞�K=hB;r�e��z�wu�kuN�u�"�&�.�"{���4[[�}����]ϗO;�|)k�^ر���~U�w,�E=(:z���y�NK����I~G8ڗ�L}�l��-◺uq�w[^?S���3_U��Pmn�>���m+r��'�@����¤� �z�5����7B�d��$8�˽���=�;E�Bc� l�s��\�s;���K����76i�U�z����{ې1}λ��t�Y�-���潫c�/��ݾH�x{*!rV���X�*<���ұ���3d..�}iJTy������^�M`e��ݢ1�bmQ������z��n|R74�cՔn����#��VuRi�=���~m��y�;wS\�<�X�
��w���p}~�#9
<�ʦھ�\���Wl�sZZ�g���&�w��v�S,߫�u�3��#s/z�x�@�NG:�����������!4_
9�Ժ���}��:�钯Sƌ���=q��s�1x�R�z��	B�̲]*Y[������:��ꮩe���h��[�ٵ���c�@��*6w#���svu��v��w��N�l�d�&Y��b�D�;B]�2���������{�셵�y[�������sF�5՚;�n����j6l�bU	d"���r�yK���,w�Y��uް/PǦ�9I󜫁��ְ�fGv�)p��P.���܃��Z��f�ף����C��Td���*�;r�?z�9vm�"3׃	�\��x���l�P�u�vY�}����*_A�6L[MwV@Q�7"YҲ�jġ[�vN��u�S�����6��]|����O"��z��=����q�ם�/^](N6:�f�4�o-w�ug���b�SE��`G�Z�3���幔&�G�rѕ/�_s���÷��d��ڃ�M	����9o�e�|�X�w����SN��^6�q����U�߷�mZ�z��qa��D'¼��['���^���t�d��%�G�FeI�pR��׌��U-�z�7��r�#=�|���[uZ�>]ǟs&�0l9����7[u���f�e���"���;Z����χ�>_s�{��r�V�pD�^X�pQ������US�u��*��w���ۚ����FN,
�
�AZ*_H3װjFR��n�����[B���BՎrH���g�z�EB�I�����-��+�l�1R��H�s��<,�s���x���1�8OM���KyP�N&K,^5����#L��=.�<�-�\�2�W��!��ů&1:�n���i������s��:^�yՊ��3rN�4-(�(Qs��R���N+�t�b�����RU�h:!���w�x4g2t�-|.���kZ}˅����Y�<�;���W�s�"pj��H':.FiASN�\�4��6(Z�t�Gh�]����#u$�K��Bgmu߮v�ur�oX��f�OD����:�z7����]u�nxߏ�W$�=�Nu���M�Bv�ǀB�
�n�v��׋5L�J�ְn�75>%���6�e_9�a��9k,I[0���]E�5ỻ���I�u�~��f{<p�T�~������d�|�䥢�{7~B3r�3���\J��qv�T���<�-f<d��;Pt���S����J�ᖟ\�nJضf�d.��Y��R�p�6�u�,:�S26����6�J�|ki�c'p#}ע/�,�q�9��Ҟŏ�u�qx.�/j�j�QLiC�2����j���pg�Ѻ����8�{6k��[�m(x����Ķ�K��u�M��ug+H*.�n�s5�<qd�Ӌ4*YB��8"�@⺆$z�Q�7*��|��O
�9
gj�˛��:��E1�]t�r��{Wmm򾆋�Ge�w��EL:����.]�7�\���pPJ��;����u��x��:Y��f���eka:k<�����{D�o+��<�X���UF����M�c]�P�c0e�GU$�՛ּ�%^B�&hhDC��wd�\�m1��N��LwXڔ3����:�?�<��]�zB�8��Qb�����i��ɯ�����b���~��3���e���L��f��A��4��9κ��S{`��2`�sE��KK�P��yb7%�[���N��Յ"lfc�]����6:� ��^���&攇=��G���j�Q�V�k\e��s惁.���ޛB��������H���m�|��5�eSU�kr�'�-��ZE��ju�O'��r�J��F|�Jj��Q2h��]�[�um��y��D#�g����X�R.�nc/A�8�qJȱ̘<���Z�\���޹]�r&��G$�t �>��d#@;r� ̿�֋��=r�(�2���y����5�p��L8�O<;�j�PkDφ����7�+�)gh�%�q�K3hځ:I���j�z��f�+��ihi� lþ��^�\Q�M�x�N̛��`e��4,�\֎;;����a���Qض"2gL��~_s��y�wS/��G����&R�+,���N�[��&1AC�y`?gf�\le�������
�uo¸=�q����O�>��ʫԙRME�����1���+���O�r����D�p]�8W��AVͷ����X�z)�Q�ɺ5�̹A�W�xL����iWCXc\���{��''CmS�����)��;��<���Xy����9ƾ3U�_]:�ΰ�Uʠ�*�k3���.��v�<�N�u��^��2p����F}��^}V�c.�09�&EE�H�Q���������K��|�\��W��a^>'6� �V
X���^��|���hh_K�z�9'�����e�<��y`�i�U$���T�اK��\Z� 1·D6ua�1�
�q�Z�68�wo����ڛ^,����{C����/�^��Z���v6��{�w{�mxJ����mݙ]��6jޓo������p:��:[^��T)xd
9v��!��ǯ5{Isg6d�j5�m!/Ns�Ю�]���	�D��f�ZWg��O4��O� ���v]+lbGU[۪��
�ˏ����n&I}*�ݕsh��8Z����s��p�Zll��1I�����]OO�g��q��2Ԃb�evuNvvC�]�����v������S[��@�нѝZ�K���_a)�K&NwN���OeX���n,=b��w@�b徔H���+��:�30#)�ua�z��OX�k`
��{��+�k�/M�o(3:��Н�1Ӂ!��W�	��f�>~~�6�{EW(6QK(��
z��4�X�#��Y����p�o����� ħj�Y��z�<����cЦԇ+��	+�M�%�WS�a2� �hl5�#|=Q{].��6�5�/2�/L�VQ�bK���%V]VSu��5����U��3�^�Oni��9߲t�o��O�Ma�ٖ�=%BLmT^(!׹��ο������>s��.��ƿk��>��߃�E7�_�~̵��`�Xa����7;����D�Ȥ���fi�)�'��D����� �U��=��PMU�����X�s���7H��е��^v��<�f`Q0ƽ��:񂎰��G�|*|�@n[���7���mՉ����[�'A�����D]���2���	w��phTt�\�o�wċ>��=R��Z�g��I|�K���{j)��E� u�!7����p'�]�4��i��K�,�Z�}w��/}�Y��v�=�s�������^�Z̆���R}�nDC���[ �9j�+K���G"rΫ<509��#LQ��ic��7EP�*uȤ`7{́��pk�0V��ۡ�Ǟ���<�S���weGl�3&Ú��\C��yX���]FJ�:�]L17W�5�/``�kI5ϯ����vUY�=�|y���+%�h�y��a�eYo��[����g��
��Z�U�{����D*��2-�K�"c]{�D�9Q�� �v�p/Wy4c�۷۪���GTGDn�G�gL�o[N������X���1�ہ�$�qL�=g�y��<oO%�}��H�\H9����%�O���g�ßy�|{@�؎�+s@v��9�;zf���j]^�����(4�AJmg�UŜ�dW�{����xhu]�L�/��j��i@�^sn��y}I� �|�Ȉ-��{@��]	�G-�
]�c���M��&}{����ܡ��6�L��T��w䰒�+D��ʏ�7A��ֲH�ʽNe8�i����bu9)�Xְha�%��^Q2�(���=����ʸ�9��%���4\���c�s��C��o�N%�P���JCI@P0�>#������fn�ǃD��a�� �ُ&�K�Me�� �D첻o2���͜i��H�A��I][�Rs������j�o[�+��I95�Xƕ/E�����J
�AB��q��(���7��k�F����0�gU�	��r!-}���Ld��+#䊢�V@�wlfK���SX���C�[7���; �:�����J�C�w6RY�V,c��Rsh�Rmsg7k�S�K_mN�qgPJ���Ɉ>��dCM�X/� �e����u�y�Y� @��z*H�
�����-�a��˞�TX%9�ve�Ir�ى���j�����n��5�uBѝ��]����T�Ǹ3��
S�/�!$���Q��y��`���G)a1V�F^v'�ܫA��B�rԝ}m�0�a��g\u|2��j�]V���5�ԧ�m[�.!�G��Z��7���i��U�$ujǟ#���kr�R�h,�\[���A�T����n)��<�ګ���	��պ�������͡ 0Wv���n�b���O���s�A���{�"l>�ʚ��������{~�^��t2�k ግR
�W��]-lb]�3�{`׈re���F���<�3�z6��f�#w7�[L�m�9�K9V6Ji�\Pv��WG�*cd�{!WS�x`7����X����V������z ���7��լYY[+N���ۖ�oj̉f<%q+��"VE�e땦��U�.b[eM��|]�J�gm���QR�[[������gqh�}�(�����`�A��Ԓ�i�u���S���z��S������euj3mS�ʵ�x�F�X����c�%[�'-]l�7+P��c7��b*�tjY�Khk0� �{^�����Ѽ��`��"�9o� ËBt�k��ۻ�<8 qi�������]�K�2���F1��>�.�SYeA҈l�:��uKk>�hjY�r�Jn�2���
��
�TwBĖ��P���*�F�$u̡�-�L���n��fZ�Fͮ<8���<m�:�̗��Q�K@�L>ܡRb����������ۙY�I�|�b��� Y����/b����*�l�d��	����X�[��7y:邰33����
^�j˜'� dqov�]@¾ŕ��Х����B��6f{�[�d���]�h�89�K�!�@V���1�Z�����z:-fb��kW��(�����D�A�� ��3+�����v�TR��b �A�{�,��F�)���B�f5۪8���d�F�wo"2Kxo�.v�`̖���Xse���7k����ۉ��u�s�9P�,�
�SS���iK�>��[��F���1ge@.�����*�Ht&��Χ��tw0�݇6p}�+��멼����-N�N�ӥ�pcJ�ݙS$8[�{ze���q)Y�V�� ��aR�F�VEDF[AAF�TUA@X[b�TH��d���F(��b�**�� �YX(%������EQT
�6����Qc��V)R�
�E�EB���¡kB��őaZ�
�
�`��h�E�j���V0E�iYFVb֌"!!m�T��F��؊6��*�+")i(��#hV,�PX�X"²EU�ԣ-�҄QImUX
�@R"��*Ƞ��-�
�QU�V�(E�)R���H�,�E`�	XV
Aj��T"Œ�`#)J���UX�PX�լ� �,+ ���T��Q��TD��h�TX�i*Q��R,�b��B�P�У	RB�"DH)�u�{���i��g��|�@P�#��W|�i�VR��XT�k8H��A��`�W�v�|��f۰��S����G|�qFb㫧gs�2��]w0�
�2�׳�����(9����%k&�<�y�ߓ�"j���̛��ok2��oZ�S�2����k��ќ����C�X�Hf��Nx�iRj�ݴ�j��/��뻈�ߕ_%�"�ҝ�Q��S���:�+u�MX�c���B3�N���^������5���Al�G�a�6��sz���q=�X)���~�Яp�i�������1�g���N#a�Mt�8.S�g��4Tڡ"ҵ5꣓ܳ��y��\����o���q�r�A�u^}|���N���Hq�nv&�lc4�ѓ&���i�3{�ݓds��}V(��Urt�.>�ھ����q}(V<��k�{�PQ��@��.�%��p�^���<���]����.�[�[�]���~�f�W2�f�Z&n{�Z�{����z���lN�Y�GJ� ��t�a�A��-�e��hu�;��g;b�{=��k0f�{C>�D��>\Yϥw������o����Y��e6��V��Y��l-�
������C�e�\�Ƞj����yGz5�x�˳�f�\�wj-]�V]<���y��6�5s��Bt���j�ƨ��-�x�y_m�E�ĕXC��ur᪅ث�}b]������� ��Q�
�Ʈ� �_c��}ٷ2�A0�}h�E�#�jj��\�a�=�"����^Ga3�ڐ-Jw�,�C v��o�f﯑��f6L�Ә̫��~�������c�g-�'ZD���{�̘+*va^"SDo����e�3f[ٳ��Y.��� n�a/E�`O��"��sze"R��>4ς�<]��l�+�ϞN"����ǩ#'�����b��Z=?�;� �7o3���ѪF���}���U���%,�ZA�*�����Q��'�!�T!�\���߶`��e�Ζ��>��;�XY�9p���?z`��׹璋��KCH�3�g�z���"Ĩ{�����=]�+ �^���#y�2�Xd�N<&�PX�唫��h]\s�Uf�qx$jK7rݔ���Wq��d�e�����O�?�q�����x�"�j��X�ʑO���Q�4�i�����d���5��{EӍ�9�@Hͅ�4�A����#.�-��,s�4jzet�\R(�ƅ6W��E�+B�«�SQ.��{@�3,��wk�t<}�W\�q��m*�Etm�a�#T˶�t0��z��ͺ�q�����]�C{�K�]˫:�V퉭]�;�Ԣ���JY�zeǨ�[�=ޭ�S+����WVi���vM���:�g8X��o�ٴ�O�_TM��녆-x�iB����;����=�83
��n\����WLv<)]s��H�Z���\����3�[����ߔ#��ld�ls�h�X�|�'���Kg�pp��lCo���
zYX��T�Z`��N�wU�]����6߫�ř�w������vk��y�nq���ۅ+��9�3[�R!+�Z�V��O�ʍr�S5�:s�Эt\K�9V`k�=ԡD̪,"k������v"`(a��.���6{�Sy�K�-�zQ"�w`�:�.PK��]c7�B�oz�ѽy�"��p�'J�F����~�y/I��XKb�����^���fh���p�n�י�4�.�؈"O�➢mz�[mA���?iЖǢ��< �ys�7ێ�{wVϊv�<�~���bx-5�JĤߍ��Q��~C, ����\�-o*��o��H9�OS"��⦙zfJ��]�F�%V}]VSu�Y���n�-�#�o}��6��3,B7����-a�"FE	>���
+������I�����3t��Lr��;/�H�<;[蝕�z�@��9��1�q� ��$�k�aV8`ܵ���9��9�o�a�hJ�C@���<��4Ԯgwuvw�4��wV��A��5��^�Xʽ�SL|ŉI�e;���*ɀ�雦<ivU��n��FJw���>��~�Oz����ouaޗv�SZ��ݓs��Q���,t{�������Q�A���"
��/�u�{���^B�����OV5d���u6�T��n����yl�`�ؒ5��
:»/�zυ,n7����X/C����^rwge�g�
��y�V�����YX�.:�G�~�~Yk�F�2j>IŒ!��[6�Z,�W9UH���<�S������ڙ�^�qp��|W�P�U��+L�7^�A��}�lp452O��9�wnk�� ��[S���J��[wǴX;zYskp�����76�=�ƫky�>�i�
�9�2-�Xkӎ��{��Pݭ�8��C�L/{�ӟ���.��|j�x.��6)�|Ons���jU8�5�K��󡻆7g���Y��y��� ޣ�E"�#�q4��4��i}������}Y��F���43�1�tq\oW���뭮�b��mr���-��|P�I��@K�hۦ�q�Wt�o��YS��ø9��q
��O�
���Z�� �Du���7��m�0��d0����@̕ �ዀ혨P(�>z!ڻ����Pn.��9^%��,��׼���4�y�aTgE����r��A,oo{�h�Ij�{����N)jT�n��_W9ݲI���Rg�<��'|���8��5*N�Q^J ����I���6�Uu[v	��]�T�bE\~� �w�=�Tz\l3�M�2e:��%���I+'��Lt��5��)l�u\�-Q�f���'"����Д��]�Z��2�a�n��:�Y���'��;(��Ϧ_c�N�v��	N`���e�;�p`K�"�ڛ}��ͨ���`�{n8���2fu锲��,�"�����N��n҃��0ҥsq���q�H����aK�q��M	|�(ȈY"a��g��dP3�ug֞�sɝ�V�	��w&�0�w�]��fJ<�OT@�����z	����G~���#���.�	� ,��2ش̉�j�7ִ�J3E)yt_�j�W�_eǪ���[hṶ� �xd��C�u��Hz���Z�
�����u(�K��ht��*0�-N���B�Sڡ�щ2N��`BWq�]WS6wy�_�����u��.���j`�/�*��k@�hC�Ee����`�'����7�K�)��S�8I�!��[�U.ʏO_`�-&%��9(̰+,;:�Yz��a*�Ɏ'�Uˎ�:�J�����74�댼v�b����;}�׫�L�DJt���c�����`�M�<��]���6���������WB��w;�8��>�p�=_5�l�X�8�{D���$u�}(g<���P�yrJ;���݈f7����2��z����B}�q%�U6���%�2� ;�4)}�}��1ď3�v/g��O#�x��w�A-�1�ZY~CH�IQ%�p6��Q!D̸H��P�K�����ɔhߋ0fг�FeoQ.�|���J�d;�K	�k��eV�_��"B����цr�-�^�����>���\%6�:^�PL������_��l�m`�W����$:��0v���b�����v�0��TI�����/���-N�����]�!���S�WAr}�b5��>�.$]�&AD��$`!��^k�h��+�E�sb!�B�u�uk����}��o���v��5M����xh�P)��ݷYf^��v:�����)>Ԣ���=ϰ��HU{��m^�k�z?#��2k������H�01]6��}I��U*>����7��ťQ˄�A���p;��υ:£�o��'J,�)ͭU�yO�B����V.2�g�����v"��'7���ھ��`����j�vs%K��S���=ޛ�4�Us3sR��Cv�<�w(��Z�(�c3]��J���I}�9���S}7���đl�쌮Geo�z�-�]����%-d��_q��wCqCX�_�3�:&[�Xd�AǄ�AZ'VҮϢ�1�U�i���-�������#�\Ս���~���q���}��B��nN��qG�u^ݛ&��%��xb�+ձv�K@2�Q���9�{�1�)�4���F��a�2t�K���e�v0�Ys�W:J�>^'eV.}V�a>�A��c�,�8�/�gm?B���>w���X\j�s�J'n|�أ�nU�Ǚ��Av�F(�c����I�fЍ�H��-�ߔkŜ���{C��,��j�a�S�m�y�sw����z�&������:lg;&�ޖ�\�7λ>g>�s�mm'2�Jd�����nˠf_5������w�5��QEs\1SV5Cf󝦅g�����4*�br'�kb���[v����Q0I��(�k�/�Vo�:���nR����r��D���+�p3�P�c���G�4�FIϞop�ϲ�Zz��Ļ_���W����^K�y�e����L�#��N�V��JuyNW;����V����O�6Ug+�Z�Z�p)P�
\Tv���q��̈́��V��.�j��3���+�]ϰ��r��r��$������Nk!J����y5�EJ���Pӵ�Y̍J�������.|�J>��s(�9��N�=���<.�͔H����OQ'ɑ�B�߰�������c��5'�J%�/z�S�;a��~��dCx-5"��f�h�lWS� ���̬�ٝ�;�(^A��aO&G9\T`��0W�@���§ǔ�R��r�Xӕ)�&��x����5k�����u�R68�	c���C��T$��zp9������͞��B�u}ݩѲ�\�~����V-�c��Z���\�3�3��!�8pꈋ�����i�kg'>{����Q;,>�����էm����A���zC��X�s��Ȍγ1%�Y�N=c����iX�C����
:�+����R�(�|<����R��n�����7Dx���:��ڮ���]�ݪ��� �]���y9r�QǳGܗE���2�C��)1�u��U^��皜|����*;@�d��.��%�+�ձ[�+Q�M��MR�Z���p�Ot��~ww1*#]Os_��U�]�����pQқ�,�T2b�R�үºmo���Sۦ�w��{�+k �M����h�pȯ��i���6ի�$F��c=w��U��Gu6��.�K�Ku��\����Pu^�5��-���Է��F���)�膸3;�S�xoX; �-��ǝ3M]ޔx��ſES�u ��#�of���v�D+Ý�"����u�,�啯��I��][o���j���*�u���qt�v�����:`�z�u�(�d�P_g7U��S����Cg�kb8�.��H��q4Vrg.������_7��<7����9�{�5��3�v{�����:�#6��� ����CI5�R�Yu\Y�-~^C�����쾴D�o��bz�J'fG����/Zg���J ��P<���`�s;]�	[�5y�QN�(dH��r��,u��Z�r�A�N�s&Q�S�!&�!�^���M���'7�r-�s}�3�tD�_�U���Sr�hf���',	���e�hJBΉ.�*3;�����Z��1�{�t�GԊ_J�T9g��4�L`;I��0+��Q~�9�;.��T��q���;��s��jËԆ�t��Z��H=��<}]�+<�zw>��~�K�X�vnq�4}�����aX�W�%��-��dU_�H�G!�,u�~���N=��s>�'8���,�����I�!�:JȁDo���߶ѽ��V<huv	B�n����~Y9�f��4���CP�l;��y��>�J�1Z{֮Y�,�n�=i�N5�ɸ��0w��J���CrZqq�uV��ԗ]���n=�c�u�R]�WN�ݙѣ˝�
����ÏA7�mn
����&��+u�M�*ґ1�������N�nS��h8������{��q귽�mm�͟�%�*�M:
�c�����~q��D���6)>Kr������3��}'S�p����5��-�1Xbq�᛻���a��ţҩ�gcU^�����/�/T�5�:"��d�]gWh��2���{�֠hbBz�;ct�.>�D����3�./�
�z���4�����w�%4��=�WG���>����i+.�pH�v��,蔰�w��μ�z:�R��S�3L_5{�PȮ[�f�����0�<$���]�ް��z�������}5�s2Þ����U0���کW�?�i��y�q�,Q�Y���H��C��S��s67�f��>�˼e2�k��mh=��4���s�lcV&,C3jp6(̼�H���Nl�̸��o�H؀�����ҳ�D��϶V�i��[�u�O-r��^>5��ַ)��=:�!��qf�y��L� �ԠU{t��Ք�]������yH����v�_w4�12�`�����[��tY;�v0��ut/n�����܉�M:ηz*6������t)�0��]HWl4W�H�ob ��5{�be�$/��E y�����Lj_0R�[76F��������㓀��G*�[eX�XPw1�����A���L�v�8��;F	���zڎ��!��i��jtK�7� 1޵qw��.ZO�4yt��IĄ�L��,^-�X���oD��,a�[��'Q�rڼ%��< ���N͐殒� �(_R�[Ƭ�Q+yN��#�0tI�'%����;}+kk�+���
�I\�E��9�(���ɝ��_����<⡈W��o��%=C�| �b�"5�F?��WW����:+����92P�q�QwV1י�E}��Gl��l\�Zb���&�Q�i��wL'G)e#Ӫf@�_nt�����#�V/]����w���M�H-�	J
o�<��n���� ٕϬ���5��Q	Įe�A|A`u�3�p��e 9vEݒ�󗵲N���l=7��u܄W�S"*����IL]��6�g+_;�V2�i�&��2Q��ܳq������P�c�.k_u%����l@1��6e�	Z�/]��y���k��Gh<d�<�ʲi��rv��4�Ei�l��\ϖ�ť��+8��+��vVTR=��l닭�X���w<���]n�4�h ��;�+��,�<���a_u�j���.�;����lM���><���{���i��G��.8�J%�ͥ��šb��B�'Ѝ�&�ٴ\ki�a��;H��6i�0��cHef���y�/��H(�9ש�(Wq�cͱ�#�v�y��E1N�3Hqu����z�ҽƴ�
���s�ܻʺ����Р���3dt+��2��k@���1a�f�\��a��Ec�,wBv��t�N��]ݕ��z������IӺ���5��E�ok�>;�������I#EG^�acyv[����*tօ-`NFqyR�<��.I�,�W.�P[�-�Iu�x�����Sb�ݽ�.�U=��n�}y�Z�w���R�Ѿ1�Ӹ�@��[g�5R�퀡�v썘�5V�,���8[4��ԑ)<
����.�M�b�X2�v>��Ȼ�b�͋;D:�@h�ح
�H�	b��8�F��������{nE�����VN
҅f��֮���ZѴ��n�<��i_>��k����n��a�z�z�K-�A��y �)�U�js곚A�2����3,�����q�vV	�KY銷�ƗD5�,��s:����v���WCkA�,D��q���U���X���s�L{]�}i=�����ʒ܍>���S�X&T�:oC6;uN(�oXAE���+AE�REX(�E��mȨ�6��ATEd
������ ��XT����Eq�KJ��ň,�q��P�+0Aih)��̢%q�dTQ��3
�����"���V�DDe@�"e�� �E�0QE�Z0�[C2�fe���&0���2�EX���m�Ҡ�((\��UYZ�-�-�����T�AE+�c�1XZ\eq�ШVd�d�V�*���)�F�R���"�ڲ�"�
���«2�������\d*`��@�µ�q���Z&[
��ʈ�aGE
��r�)�b���"�E%eF�,YP�����1V���IGDB"#wYL�JkE�[�m)*��:��k��@s���M�^�2�L�+�;n����;U�d�ʜ-�=p��&�}ũzZ<��<κ���.��&L4H@��PK�z-�c}H���r:�Y�oj/�9���|�w%��S������dC��a�E�'�
d�V�N�k���#���✛�OQ�ߤkP~To4�@T|�f	*�[N瑟R�ɮ�����H:G�o�R��V�|���^��(�K{E��ys�."Ua˄�v��<w��ҩ5eG������|������rK�;=#��1Q�6�V|k��L�0w��/%�ITx��0ӯj�V���_�pI�0�[Y��N�9�+��w��C�z�-���~���{�| 8f��&";b���#�u$��|����	eX�A��֛��<!7�b�5=��kO�Ս~[�6�:�sV���җ9Т�z�?i�\%�4�����uҸ
�|�N�\"���^�����9���ݜ6O5w6sh0=w}μa�}:o�J���8jl%��y!G�Ū ���=JW �6��=�ɓ>��D�t:!��H��o4���Y���[b W�@��F�YU�Bo��j�d�̫�r��p�-�3����n�MƎ�txHL-�x�b�ze$i�R�:z5��ap���a~��9&�d@�����4�
���!&���r*k��G�{%uwk�ճ�\�gNr�[�V�}�9�ԮQ�	bi	 ��ۄR}�X���;g#)B��G�z���CC���w�Ȣ�y�t�[>��cѠ��ĮR����\�b�s�JW|��x��Ū�,���ڲ�����v������H]i�]������x�C�UM��oJ�*)&��4�IwJ�Ň���w@�b徔`Ur��jؠ�&�����ÄS����Q�DX�(��*�A~G
���~�q�;�t�ù����ɳV���w����Ň`�X�uWSٍs��,(� $��k�ȿ�!۽�j�J��zPLe�{��g3�<���{]�4��+�{��Zk>��)4@�O�7~ۜD�y8pC��t�+�׋�!,!:��ԇX]�ȱ�_�3�YG�v!�d�\���a��}�u���v�~�S��p� �hܱ�P}�whx���J��ڬ>QZ���	̽���^����Z��#��bM���Ȗhƛ������0W<�H��qu3��R�g`�/�8�s��g]��)+�����{"
�ob�u���Q̯1U7�n��n�hZU�-�����ٶ �a 4���Uu𨲝�r�O$G{J^�w]�&�<�{S}��v��l3�޲���e>r�X���7k��,Z����W#�Xw�8���ꝷR�jk��҈�$�9�Jhb���j�[W���<�-�v�����>P����\	�n�w��uH_�a��Z)=NR����P���@�j��Z[�20ͻ��J�l�/'��"=۳q�"��t�vk����$� ��(&�'���fb�b��ˌw|�UW��~|��ޘ��ŝK}qq	�r#9�'Y�i)<���W�2�\�+�� � �s���8�Uph�U�;�l�!:g2y����~���V�N��U�X��`��V5\[΁��"|�_���7^ZN�Aq�������cyw�2�EX.���.�#����h���N������\�؞l%���s��n}�ޘ$(g,h�^NJ�#a.����]�4��F���Y�r�m��0۔���l-��Q��wo'��_����)r�tAo(4�JSks�����#��E\��{_gzo���"�s�������K'��G�/Zg��Y�U��F[������z��+���Cb��=�la�_r��r�A�N��̙EN���K	!��G�1e*�}w�%�k`�[\�>_	��*M�[���� �9�o3؃�8�N�7����y��v�u1�[��ҷ�>õ�p퇵A)�A��f�9hsy��P�úPwY����CP)b���͑-��,n:��{k6���㇗>�_�[�w�9��k�}!��s�]� ��U�tꛔH�Y���u�ȵ9(�2Ƶ�ZkfX���ܛ������{n!��Ly������t��v���0�lTY�Ne̊���S{5����D���h0f�cq:CI��L���hÄQ�~Y���"Y�����Ҍ��s��'I;2��Y���R�*T��W�%��t����_庨�P�mG��ؖ�C*�/�l��"�U���t>�H�m��ǀ����;�U<H�`��2���ru��yy}�y�ؿ(�Klm���7AE��=�΢A�\z������j�gb�cRRoeU+�L�Ѭ��>]^"�(xإ[�W���
T��F�P��a�5�����g����gc��z��2�kB�ţ�5l����r���@� �z�y����$!���s�<r83��e˞Oƕ��!+��zP5t
����Z�}�7����~��k����1R�gr��
�.;�$�B�ǔ�A�}���Jr�n���[]%�Nr���6�q����+�B2:�.��ۛ̔��V@t�dچ��@�c������:����+��!}9!�3���nI�N�&�cj�9N�|K�Vf�9(�<�AM��=����\4��e6�o+��\	��ru��9�ӏ=}.��h�>߱��dR���ӿ|FǤ��V��2��uc�nɧ1�lot��Ԓ�{Thh_�0���ګ�i�:8����tz
�O6�޶�*4�LZe߽'y��A@ew,�Mr�,��9�#�3`cV&,C3jH��0c����~�7��]6Y$�hFm�`�t�$���V�`&�ju�O-��[��9�ۼ��p�ks�E0(���QX�Q2`4H@��R^k�o��H�71� ^sR�ӧ3n�3��^m"��mcY�&mJ��hSE�o��"�D��d#�m�!�s��>m��R�T�>�~E̡�Q��_%@{ݥԟ{���u�#&Mt�P��=���ctq緷��	}s��q���`<�~!��yk �J�.q�G�O�c��K��:���.��o�U��9әGJ:{��!��r�՟X��	y�8��v���"h&�"����:n�o1��zU>�ޖ�ݥ[��j��b��}t2��9>��'Ꟍ��@�����%��SƐɎdl�r�9���{]�*a�xw�J:i1�$�7�O��	{1�6�,�NP�3�tk��|%bi*�����}ɝ�L�û7aڎ���.��y>�
|�l����m��;W��`m���ʧR������}Suf�ntR��/��U�蘟%DmY�x�ߚ�d���P>{]0g!^x4-��Z�gH��[P��Y]��UnF2�!�F슂�2q�:W�\ҁᏗ��<h�<�^�"�o��Q{�TuX�
��:0�!�}z0]{V�q�Ն��,5����۽�����q�u�y��O��&��D�:��Se��ڣ^,����{^�'�t��"Ӈ�5�ws��#��78-p!��o9�67���v���X�e��1�É�Ǌ��9ӎX� W��C��ʍ4�x���T6lg;M
ϵ�1Xq��}���Z��s7=�}|��
s�e���UĂ8��{�'�Q��wZS�^�� H�fGƷ��s�c����D�邱�̋G�$E���o U���?#�D5�}��4b����ګD������~��&
t4��P�u=�����[N��Kf"��w=R�w�[���Ĉ�
���ӭ��?_E<PӶ�d?�!��Zk$�JM �-ʳ�Ǿ�7�r�����|o��BF�hRϳ�������1�I޻sU�sjn7̲�v o)ogkF�Sh�m��ܯD�n2�Z�*UgB��-�(�]F�}B�u�#�V+�&�j���IA>�r�(��:H7j�+;W�R����ܳ$G;ji[��ݺ�<��絅�u8�G��{T!�r��%a�QF�uA� N�Ufa<�iҢ���ffw�FD[�C�U�or�"��A�{ٖ�.$nJ��ڬ���Ո�Ԧ�6�o�E�Sk�\��q�1@�c���x��e����γ=&��y�~��5�'�<c�7x��z;Ub}��M��֣���EG�'i��_)]�N�U�{z�Up�!U�c]ʧ*����ǘ��B����m_�o�%{m�i׌u�vZ=g¥.P�2zqy{{���;�LC��}ͺ�<z��ZUü��۸�Ո�a�X���B��AHeM*�\�<����-lH��	�<��w|Ӫ��s��k>�v�����C���R�����B����O'>�~�"�<F��^Wi�;�8Y1��r���ÍuW �4w�l;q]�!�_�=�������ҹ@�i�5\E�Br��ܽ���t������vs�f��ij͞��eީН>��r����A-)�+CF�ܾno�M+�4�^X=#��AE���.���붹�+;��-�Se�0P�ǘ{���$e�W��ȏ�B�խJ��l�y�816�	�$l��29�\5̃b�8KU���f=���î�}W��ۯ����Y���sM� ��!��D�J�u�Tr�rݬRhŰk�n��o,��\�IQ$l%��Yɜ��%53�}]�M�ɎO�1��'�5���� |%����\x���B0lk�}��-��Pb�(i&�{=��N���Wos�8�AuP������ϼ{S���N���(��>���Ec%[[J��tj��%�Z%w>�1�B:$B�N����t��:�P�:o�2e�َ0ݱ�)��ιu���M-�JV�\@������S�@��T�%����@V�,*w�9g����e�i+8}�$�}�5o6�����4���M�],��� ؾ��ƻN	���}����T�]��K�]^R��zV��%��`��������3孑�(R��Z�.^�*��&1��
D�:�E7��tk�}�q������*q�a\}��	x�:#�Fm�L}�7i�,��ѯ[�Ol(�t��	�=�����Q�����.w*�ߕXq�&�kpVG~��I�:���˽�j����ͽ�hAYBj�;��lsW���ʌ՞�d���g�&�}#��V>T.�q��=�tG<[%��ge�O���j�K��`��;�e�tmv�b����w�n����z -#��ye�w��3l��/�C��;��ZΫ�cz���M�Scth��뤔朖Ƿ�o�l�s��I����'��^Ԗ�ҷ�$���4��� ��7J4�|�Y=a�*ߕd[�p���a���a�6jkx�Z�GCޭڡ�V�}�Z-)�geSU^�c�]2&���L:�xF�d��3��je��=CN�<} r`ӂz��yk��O
r�XzS^gD|��Z��/��uȄ�c�9�:�G��Z�q��S��m��۽���;�$�B���6]����.\6�=�z�׻9��u勇�U�)}����Eb[�f�����0�2&����g��WrB�;���/gy��@�RK��hh�4���6�K��У��8�KfV�b1Lt�tM��$�g}FN���tXž2�\k�6�5��F�绝�ٷ�&�m���*�����ԛSX�%�Ht@�`��{�`�O>��ZE��ju�O*�>�����y�h�]��Kx�Q�����p�v"Q�Kxv�Iqְ��j/n�Zs7��,w�_.����f����|�dY�0{~�W��M�]$[� xQV�X��Kq�-{�s�L��[T�Ԧub}�y��ǍeJA�W�B��撄/TH�'	��A�͕�X��E�VV.b[�oU���pU�G��pTg58ut춤�|�]]���R��2��vS�ݩ��ڶwR�kZBEڒ��fXG��PT������G$�G�wf�ġHlʘ��
������t�v�R}�'�4OG�w�ɓ](0K1���tet������`��n�v�ۄC��v�����c�������9�T�8e�4+r�Ť�U�g��F&OP~4p]��<+�㮳���zA[�D˔8���	|e�41�ܱ(v=�+�,�*C�jh������t_��0v�d�<�j�-��~3��k��z#!��O����I��w�u���wj���BYQ �i��t�b���K�=@,���2q�X�i�[8m��ܚ�!���/���w��z	�Q�љ9�=b�I��V^�k{<��Kl�M��3�������]TK����s�!�CO����bp�+�b�%�ֵ����軎g��߲=����!4N���&��艾t:!�;��-���g>Ӳ�k���v���3��N=��5�l�#i@�ؙj�ʌ?mQ���vM�;D+�6�_��ζ�U 쁫�	�^}���y�����r��]�-\M��b���GFr�R+5X�;��p�a�ʾ�]D�
0��o67V�k`��gJ��m��� �iũ�vؼ�y��En�{)h��(M�A�;x��������jޑu�w��<8�>u7^��kv &��K�M�Ӫ����t��4[�����T�0v�%l!<B^�t�j �]�C� NZǝ��za�q�I�A��juP����\=.T�m��@�ҥW'sUf4ȂWQ��vvXװJig]����,�Kut`�\tw�P,�jܖ�1�Ê��j�X ��+����*p�>���'W�g2b����wA�N0$�=����� 2R�qs�G�HD���F���V^V�jf1K�SR�:
�k�]���֔�˜��h՜R�ÂM4#�@��
N����_SrT�����cHs����Z����T>[g[W�Ԯ�*:c>wsS�G �if�N��9�,�#��:�������K�WO��ff����Ҫ�m^t�Y���y�U�I�$�m��EI�*���������7t��Υ��l��Kv��h}��I+7-p՜�rd<���k���C�yRWNt�Y�
f\��kJ��;��9�^g2�7�8e��R]���z�wPCkter)g*K���ag,h���j�)N*P���ʜ�+�;��XV�b8��{㶤��إ��I����GC[|s"2��u��{��
���L�xV�
�q}����#�V�zc�q���nU�gvv%K�R�L�>}�����Z���}h�j�|[7|�ڰ.YxSm��;��J�*`�;�H䮙�`OY�O�������#f�]q쵷���˦�-�[t8dy��!�,=v�R�����B��G;v`����.��[0N\�EYؓ��	�Q.�Cy{E�������볁jY�]���68Ld��o�,�˶��+�L],�ۊ9�S��j}��f�{N\g�a�|Y�ӯj���}0Z=e��}v��f�9�{.&ѝ*`�f�}�����π��>��)�0�-u���R��u��;�\�H���/��E�֖��0��:!SDJ-�f��:/A�]Ê���*��<�ސۑ�V,֮}��iѴ��'>�jC�7XS�j�9�;���Sy�:� ���jd�p%���e,�;!�W`� �%�Vx��!nY��{:#Hˌ���I;�;oUۡ�6��U
s�pZ����{m�䬱ӛ)L���cM�)6K�]a��T����е.��)�{n�+�� �v�.��i㝮����zN�W,5!!a�G��nT�{c��H$ ����[2�t/2����L1����ko���X{y�[�z�em�U���A�#�t��aڧ�yݎ�����]=�v�j̌ح9y�c�L���;,Z'4c�z�4���� ҙ�;�rt_u�ee&���om��˥+� ,sg.A(啶��q�l��6W�_
m�>�Ȣ�*cb0�P��*%�q��b0TVT���1�����2؈�E�+Y�(�A)�+&[1��H���Z���6�r���$D2�XV(���T����R�m�b(�(*��ɖ���!�[B\��k��X�QV[jUEX��,F�XW-����Qm*�1��#h���AQ��*��!Z���Z�8�ŎZ0X�*�A��5���������[-lm��TƢ
����UJ�R�m*e��)X�QU"�Lʠ��PkKj���SVT�̹E1��s-��q�e�ڵ**ԕY(ՙj"��2�B��*
�F������De�6ʪ��1�:���{u��8��P\,J�A{jFN�����D��|�u��ށ�v�-*]�y^F�dt�� �+����gA�0��c3jQ��+�9�~]��V��JLʿUq4P�(�����Z1a���š�������7�cvY���Qo��J>H� �[+��S�6W�׺�Q%O����`�)\��WPĞ8�A:���'`��n��R7ɑt�5�x����Z��7�ەS�J��֝�P�L�x�v�z4J7�Y�a<�~�+"ؤ׾��)=y������s�����
D�FT����$��H;���qQ�zf�YG�.� r�k���F�ֵ9á�s=�6��TK�k�r���n���W=̑�4w�����R��W���VdY$�Og�k�8{
��/���_��g����eкNLg��ؽ������r�5DEL���V�zz/b�n�KSnɹ�u��0�4G�'i��JWjӢ�l]�u3�:hX�t��9v{9��U�/dn�c��d�cVc@�7�J8'm�!��A��u+e��M�ӓ5�N��b@�����ЍWC�ݍ��t��+[�2��[{����rZ��~�D=��5���MC�t�,W�m�.�VE��-n��N��i��Pf,d�Ø�0�X�w�b��R�΅-��;�t�T�7���9u�mr�O%��Ԫ¸Pc��Z���!�hU�;c�n��Sٕ�E��k��5szھዓ	v�����o��К�����0�ST<:��J��k���N>g>&��Zi��y�
�۹����:�A��s丈|W��L���&��K�UCJ���3�]{����)��(w�ޥ�^�4��:Ӹj����`�r�W����dB��9�}x����y���w�s�iY k�yo�T�G&T(� ���R�ȑZ-�r�
#u�#�g�pkp��$�iƛ�T���B}�
hoNtu.Y%D����h����m^M���:*�=ӻgv��y�9�\��O՟0�����W�.<E�'X�f���`��xM���,���՘�;��Qĥ�1�����(f�O�m�Þ�ߵ�!�RnTbu�r+f�D���m�i�ZN�Wk�
��K�`�=B���`�C�]3�hN��;�N��̙E�Wy��ӵĔ7;s�矩��H�u���=^�lU�r�zT@衛���pzU>�x�1�J%�9ñt�]�%��������U�y=�e$Q�����Et�%r���?S�.�u�8b�_*9�x�/V��\2�j��y��;g���e�P�ϫ��>ז 90wQ}�j�mؠ��ԡ�J�b+ya�}KK�.��rX��}I}Vc�A�2Y��F��/�n������ֆ��k��N�G.7D��wX�ֹ�����/�����]y�kS�3jD�ߔ��Ս0��_���2��G��J��k��в�[���rWM^~�׳U�'���v�x��JÕ�ڰ�>��z�5�yh��B��F�oX8�<��=9�j�KOW��9��C��38��H����Մֈ��JwcVj�j����i+�����t
q(ȿR��9�&v��9����MC����9���[��A��[��$���G3Ϳs2m�tR��F��,�m�_0W�:��T�ܨ����_�jn�EsÖ�9��2�eP���<u!0b�ѫgcU^���PC��Y��E�T�I~��gg
ے���!�4Y�&8'��W�ũ0E����w=� u��Tv$�L����|��`6g�P�.I[.^��5�yg�Tp΋�.�*�($+�vP>�in���ѿ��/�ݽ���A��G)��9E�7��L���~,��GTIuV]�l�M�%�w����EbI���E�T-�ˣ�ƺs�졜�m>\YϥvO������W�;����]��K��(5Kr6�M ���6|x=�)�e�hX�f,{Zi=�XSzL��~	ל[{�h&$`�A�"$���M���8/ĹVj��%C�W���t1���Sb�tw��u�t(Nn����p��:�w��sq��q[��
=;��z�A���j�AgXVe6�Z��9{��L��x7��Vǃ!^Rw�l�����=a�~]ԧ}��$;@r/l+�*�<��l�"�n��et�\�n\�Ś�gv�~=D�X�Vz�f@�)�
&L��!�
K�z-��#,ow�"��Fh��^4s��&�ㅾP�!��dN\��J��j�,#e�#�|��D1���՚N�儵{����Z�b����z����c��Ji�G��`�����䥀S�H?f�.�6�I�>��y'oF�h���QE������f����\Y�W9p���?zx��f�a��EN78�>��۵�RFv�X�>������^wu�,�^g�+s�~U�eg��L�ݫu��נ�t��Ob
Џ�iWcW�5����*;��d�<�����S����ߴ�.1��Uɖ^�20�t_I��ڽ��N��TH#���Қغ�8���_�7�wx�'mZ֋�dcud��!ۮs��܌���=Ȩ�7Fd�s�+`X+��a�L��ؐ�3��� U��ɕp��R����w;o,s]\ۖ�Xc4�{R-���o0^�5�t.��ֶ���W�:!N;I�Lj�a��b��ָs�v��m����B`�C*�v\W�ѱ�u$����<.u�/=���k诮�\4�ӻ��rR��g.}JF!������y���]/C���>{�c|��I�R6�43*�L:�Ehk��=�)���
���Q=���&��承���u"�%�ۈ{���?=�w���p���rb�Y�����YȮ��-S��;�j�7���v�\�7λ>g%�ds�aG���Tx��e��p�MK���Lߢ�xgH{j��Z��[���P��t���C��7\��oJ�ݷB6X����fb��ϩ�RN�W@��P"7B���.x`=WhrG�zi�種*ߜ����Q"��;�VIّo�$E�Kx���9�߬}<<�a�Yh�O&���a�9��NE�{�,x��*���C����"��D�\�h��Kk�*��IyS}��LR�A���S�ŧ�觊v�̇�R�!��Zj�}W}{hJ�w(q72��!M2bb�]L��a//R�yB9�⠕��*�8k����L-lt뙞��}LW���-VTu�+=e��x.���a����{��5r��Y�'ۙ��H'^�MU;�LjeWr܊��z��e*YR�H����-�q¥`�����dkU-�ˉ]n�
����*�:��ӗ҉\q�j�̠i��[�FJ�.���vw]�9�sԳ3{�-pђ��*��6��խ%���pU�ޚ�uqs|���to%�M�蛻�'��a�g�M��!��?�c���x��j�?��]'��d�>7�u�S/�]R�r���C��CNɝ�X���4�*<�8z��ڴ�ػ{,�qFB������}�,��uW�����-`��j�7c
:'m�!qa��G�u%��ő�˞{ѫ氈+k
�ۅ���>�ƟrҜ�.W���J��Õ�t_ ����{ۣG5)�P���w�fj��ʈ��e�UW)����y�3�VDҥ�Gk�d�s���wG`P�/Xj��8���L���0t�Nt��~ww!�^�ާLQ���5Y�Jxo:zYߥvs�r��<eV.U�SF���+��W���tq�r�r~�v�<�z�{���Pg_�u�L���"�TX�P��X{WI�i�uF7�z����\��'h��T�Ӌ��C�i`���K�}%D�'�³�'R��ܗ�G��Y��]����g�/�g����Ã�;��tbb��X��B3�mr���-��s�'����=����h����7��L��y�u�����EE�z�B!���K�.�r���xïfܮ�뺸�z�g��֙�w�F�����Y\�K��[�N�i]��;i���J�Ӝ�\ō^-2�֮���%���4w�
��%;���O7�P�M)�e�CVE��h��ޒ��Gp��K֙��P>�|j,*�{o�#�w��m|�T*S��!���в�t��'[�0�Ґ&���h'a�陝}}��۾����a$K�K��X�<�V
�}Sr�h�A�=a��jLs�,�L��j��j|�7o����h:B��w�j{d�H��a}���<\k���e����긻�-�(eJ�s�稉��أ�N%�J���1�{TG�[#�
@�����7�}�M�F�'+z^�88z�,J�M�kΦԨ�Յq�W�%��-�:�g�<�A1�1�̩���b�l��*6���g�.�x>�H��:q�'ѵ�)�\�U�D�{/zwr�)�W0n�?�z�Մ<Klm�����f�*3V}�OM����ٗy�1�Q���nR�W�>�>�I�^��`O��-�t�Ô;�|�Y:�χ]Xf���c�eS���%�Q��;�J9��2�eP��ę�����./���`�r�L��W�ӵ!��W%'~�0d�b�s���ŧ�"�۬J�u빉�ܙ�m���8\
�<7�kcD�'��7p���%��two6��o8�vB�MR���vl���R�&��QK��8���	������u��&�U��lyv����� ��̜��\BYg��&9=Oʼ���"͂���ԵǅƦ�e�e���Q*��>3�^З���.I[.^��5�yg�J�/,yM%b�1'IXQm���'oZ]�P.��~�c�=tEb辱�͸�~Pȥ:fpiߋ;���8�|������,�;]9�ξemL˅@��N�=sA��S-�]7��lgQ��||����'Waж��g��e���(`�Fe������[@MT`��2�\k�6�:]���s;�I��I��w�n�d.�H�WN���S}�����
�S�$��Umu��)L����`�� &��Ϛ7]�W����-�rk`3:�9�
��dx5����(�0�!|C�(�ע��K*1��u�9�v(wt��ƶ�"�C���mG2`���{Ц��.�-�}�wF3�V��%����>��B?s�d3�����uEF��䦃(
k��cueșYn�aނ6�/�՞$��v���T|l�b����4m�����<<J}��=ʈ���G�2�x|sW�9���F=����Q
�B�^�[ю�D�I֤�V�5�٧\�&y4ej�g�RzOY����0�������y���0��?H{�p��J�X��,n2�D�//Och�.��:��-��ӱ��̟.�vf�g%ڲ��e�`�Yցёt��>g�y�Wu��P�?�3�
����Z�~���׊+�W1��;�I*g�곕i׵Z+ex��gV���#L;���j�:��u�E��{��Wlq�|���H@�3����]ڽ�8:&'���6�ص��v��d�r�X�ՙ}�U�{��шW�7�il��Qr�긆=/���Q�j[�Vq���ͣ�*nL]��'{��1y.����8�@���Tʡ�wk�q���zo��a�\)]t����-7q{!:�|[}�j��5\��\�"��3�m�Ck�&��C���IN���kś�o���c�]v��+���v�@�p/��ѱ0Z��>�����y�ɽ�h�c���!�8;��7@΅�{&-�߾Y�e��I�ۅ+�� Q�Aص]�-\M��5z���� �bI=��O.wM�x��g�P8�	�����+J��)'b���~�ҡwU��3��O;��Z,�d�~�9Ѻ���\�
dئ��>�!��u=H�V���+����޶�u̪^k�Dad��7�R���&�.�S���:K�B�޶�o�3R4}�D�ϟAj�%N<Y{B=[�r=��]!�{v99�� zM��*�᝭�2��-ӯ�j:���S�?/��+������kH�ܤ�X���k<dddEӵ_�EWA?Q�W�'����Kb���c��J�+=���<.�͔A��;A]ٹ!���6�ӑ* S�I��h��j��o��\K��;a���.�Ȼt����E�.�JV�X2���K��@�_%���@�<�A��.����{�d&s�K5����Wָ�ZU���yj`�+�X�C��9�U���\)��*�vޛ9���ĠA��M�e�$zZ���qv'��j��:�J�Ȕhƛ����o`7}j|j��r��`c��9�9Ƙ�s��#vM��G��B<�;A���dA_��$��Z�|��.��s��)�PMU��z�20qb��3jo�- cv0��Nۢ,Ed.�7/���5���y��g¢��Uo��7�Fx+��2�>��l�!�n��lUu�r�}��ͽ���6�B]�ߖQ�t�teO(pu��Z�����S�N�qF8<̹�%;�z�7Pc@��:+U
˦v�:�[AC�<��~����$�hB�����$��	!I`IO�H@�rB���$�	'��$ I?����$��	!I��B����$��$ I,	!I�$ I?�	!I� IO�H@����$ I?�	!I�p$�	'�B��LPVI��EF4 
_���X���y�d���	��J��+� � �lyN������b��k˰QM��R�	��Pª���4AT�"�F4���    ��2T��h�4�i�b0�2 a���J�SF �     �O�%)SA��  4d   �?
U@ 4   h  T���?Q��=A� d h   � �L)���MM2��Sjh1��Ld�ow^�/u͆�`����h� �t ��G�D������O�J� �@��aP?Q`����+ :�D0=����7	���=�:( ��B��k��S��z��W<��

(����3ǙιU�sJ&�QsYzCi������{�m���r	��X�U��&�h����(&	�3�CxѬhX��%����˭��zxv/�p��`��u���.�VF�\S�ʝ�z����x�T�R�nM�w���ͪH�鴾=����n���m֥����7�#||]^f9Kc��4�\�[��|���6��z),m�ukmrw$� ���E}��m�T1Y�E�Q7����b�jp�r��;/=�`�G#,&�1b�;J�2��yn��Y�?7��b�,�xPh���X�sN:=A�!G���s���|�g��u�e��<|��YO$�S��yİ��
�i�c�k�b�(�����{�պX<�0{�Շ����3��>����D-�6�K�o/-W�Z�y�G��}�~S���a�o3��GE��@�B��{�����������l|�	|�"����L�$��S��l�t3]E�@�nEƵ�;/�o)��F�m�6e�l��.��^��cE�ٛ��J֟ЛSn3۽c����]�Tv�2*s))�b��һVOP�nLo!�.o�}r�btUK��{�Y|�nl�粦)��Ҵ�*9v�%15v�E�v��g�3 -�yA��/n��1-Ur1�MS��Bzd��giX�gԶ�E��u�nY�.�Nm+��S��mgtcn��������L�u1]��goZ��˛]��a�}q�{����c�l�Y�T�] �"]�c�/�;��Z�#C�0����X��U�u]L)��vQ�˕[U��>�����XX��t:��L}|Cw֤S�/�v�:�[0�Y���kN�'c��D�SS�<sd6�N}>����"k�'�Az6Hm�i�AW�u�(zS�lXP�Ə.��z-X5�Y���>��q��u�M�&�TdӨ����W;&Lh�wv&X�q���N	��!�K�z�R�9v0sUu��T4�ԜP�����h��g�V�b�L��#�[ip
A�kB(�k�i�B�l�٦/�ERd��EƧ�P�嵎]�rL!�yGX��y�R^�K�L{�r�.=XѬ1bCD7�r*�t��O���>8y<�#B&�;�
|)�'h�hFȱ�.�Q���D���5�\ֻ��JY���.%Q�- ��)�����!��Vy�%8���	�	a%��X,��.��	���;.����YIQIF���.��z�:*"�+���{���YEb�*�j�*��8 �d� o�{�^��?�0cF+�"�~g��h��X�թY�d�nM�\ed�����|���{��i��lH�" \-�[jY���}@�س�?Bn�I��v�p�0�q�Ϝ3j�\q�Y�?�`�p͡7�(�fM���\l[��u
M;�4V�'.6�Xގ|�.ͭ��|��T�:�
�O�b�y썞������n֞2ef�u���bի�Z������ۆ��őC���wY	.ᗮg�5�}����:�QQϋb��G_+=S9y�bnDn��l��>ZS��س+n��.�Iw�{�w���Պ�,E��F$3�����".x��t�/>��j�5�B{nJ4��O�O�%mi�}�K\(z%QU���H�SER��O���Sx.�t�b�.�������N�W�؞�̝��uX�S��p�4�67��z8ԙ��0p��Nķ�#�l����6e�@���FQ��;%�������xy���W�D|���	�D�y�|��A���_P�t�jߡV�Ȑ�93K�nWz�Yb�¾��έm�5cs�/�WSݻw�M8�ٮ�b�j�|!���қe2�ūa?]tJU^�H>�sc��A����,�jԙ���=�7��D'���R�5g\�3Ӊ�i�gw�����?|�_/~�������=��w��ɩ������P��3�].GKB���B�͘CiY�z&��Ne�h%6RQ�# �aY��:�8�}7��P|S'D��9�	YS{[v�h$�vR����rAj2vuʶ�m#x�33p�3�f]�1�ٶgUa�~ﯢX̬\����S5a~'�rpz���{���k�/6��6.\(�nj[��o�;S�x�wQ��r���]*㌾f͜jt��m{��o��{��d���˪c~;0�O�!Vf�N5.��Af���B͵sI�Nb/5
�z�����F���F���1��h�-���X�* ���]����x0mo��Ԋ�[�8�]�^{�9w��j����w.�Ȅ�ǎj�`�)��V���b����M�}�<���k�}'�i�r��f��+e;��l�y�yRaർ�RG�-���t�^^�2mm��m��o�C���v�W0��S��-�$4���GC�
�H���׏�vkuo ��1�ْ:uq*/u�.�4�d^M�q{j���Eql�;�E9�}aƪ3�ߢŤ�<Q�D(��aַ&ZW�]	�/�҂Պ�zGaTd���;=�����̦�ue�@OC l��VfV�g*n�F���ޡXp��x%�����l:��Y���-qoKd̜�fнF.e��⥗01�F'
�Y���\��3�[��~u ��v��v8x�)ѥ��N5��d�������tv��R\�6�ϐ�� !�؊!�Q��o$@*�*(�� ��3wW-�.�����{
+/5�35��<t���xڸQhI+w\����	hE�^7�)x�j�KmtLB׬��"5�ΰ4�7��!Pδ�Pt��7�gM/���Mvŕ�¢o��.��� 7�%�B��[*,��)�ٶ�]!�M6�h��"�	�L��	O�hI@�-۸+5k���g:�@u֔�W}5��]�GX@u�!!Q�P�D�;�-Mj@$HH�i��h�7 �o���O�©����s���|h@Y��*gzBE��;���Yj�9���D��	P-!�Y$D�+$Ņ�%nk�M�*|��E�E�f���M4e�e����"^�����7�ka`��}���_9mkn��u��f�w 4m���O.�.��u9,�R���[9ۗ���[+o/T��Qqď�y������[�v�\΍d7�?"�Ժ�=��x w8'"	����Xq��"��;+��HfEM�ѡ4o���a�&�=v�dm�Nۋ�̙��iw��w�nP��\�Dp�yZ�ϓY���b�m�-8��!�)y=�T�W:��B涡]��}�9�W��q}o�U�g8A{�h�G�\����-�^�d��'��**�3/5e�4C���P���)�o{��u�h^�"�fPq#������=�u����=Q1P>[����Q�/����v�*�^��=�/�]�O:ƃ���t$s�T3K���F��n�.�:\/�ϱ��w!����s���/t��D���=��c:�oV�6��vP�����Ұ�.�6� �LJ��6�!��7+hl�K�r?������;��w���0xm��D.(�Y�{7{]>f��2a༧U'Q�{�|�tb�SE�=,ҙB��1�]���;/�&�C-��ĭ�����ř�)E��eE�L��=d��!���a�4�%�z�2�sV�x��P����S�ڋ[�is��p��ֱ��O<D#���7��= �*T�C����5K�Cp{�]��Y��A�v�v�L2�Uv{���Ͼ�)eI�A�azcP�~�7	F�Z��I��;j�i�\<<�h�,�{<��U�鬥5/J{X� �M�s*q�4Yi��ż�Z����-�����N6��;P19^_Cɗ�!m��f{W꣉�3!q�%�jF���zI��+��Ft��];�D��p`����1N��|��!���}F�,e ���娄&��}�����5�Qή���h���(�{g>O;V���q�rU��L�@徹+�%8�5�8�֕M�>1Դ��6�[���ج��;Wo9���ݡba�i0]��3������k|���2��z�<b�D�R����=m�jx�;���/t'�����߽��x��x�:I�$�
PB�!��{�;�'t��~CC�]����K'>��W'Sݤ�������\9f�Hf��`� `c���g,z�E�bT��9�&_6I��A*^L�kQ�폑:�5p���B�đ�a#�OZ�H���+殧g/�(&AK����r���]�yچ�FN��������!�#��HNS$J�̌�ɲ��.� u�p\*0B��f<�36�s85=��Q�q;38xF6�R���7/6�]	���s6��Q���[Ve��j]8i�cv޼����'�F/x�)h�m�ط��3m�X��,}�y�T��r�:�'�F������8܂��o<�';�ƽiMx/fIyܗf�g'	�,Vq-pw>fG�J�Egw��9=~�v~��������ҁ��ʎO��
��ȺrZ�v{!�Z׼��t��|}z=�!YYe�d�	�Ta�O+���'9!3ى��k�3G��mf�h�{����e���	#X)�z�&j'����x��#���N�D�Ry�*	�'�9KQH�1���V���s���h��|1��LJB�����!��|`�9���]׸X��i)��ì�s �^>GS9�V�m��*�q��͢�J��p�o���̱�L��_<�zX�B����M�Qf����VG#lZ���s�Z2+�m��D��h�.#;sd`4g7I���!@�UV�x�B�N��c�^,x"jj�f�`��!'�� |険��&���p��R(��Ę�Q5,q���L�@�ʃg[�W,�mA0�2�T���Ϝm��Qr`f��"�����X�޳�=7��s5L���rߖn�^A�bs��{�%n�6d㝐;��5(�i�q���\CCs�e}�W�2/w{�zl�(�RY�� �(/̅��*�`�5c�\J֊�w�r������*/!�����2�� bE%�o���!؁�1c�J�����A�2�<@� ��e���g�H�f�AN�/3�x����80 <x09F�� W�ɯ�H뙞�K`s�p�kw���KaB5���S��cO@e�8�7gDp�s�ۚ�sW� '��5|H:yNǁ�g]��96�!�� ��C	���LX�+xw����|�{�p�3l�#�xֹtD���;�����H}�C^�B�)�{��
��҉HjF���Ni$�EM�f\���'c����Z%�0gL{	j!�3�%ҘɆN��fA��\碪oq	��E��@'�8JV��b���J�e)����Va�&�g����#:����"�`x�`=���fJ6�-�u��d�ɷ5I��pocU��YT'7)�ňlח�t�Y�_5�*����L��S�ѷuCz� 3�`���Ux�0�}�6�u��{��~�����B.�۩��1��~3�GE��� ��ftS��Gbz���k�<���B}ھ�D/y��E;�V���j���R~\��36����yuQUd�^�)�'5�����;q�X�|�V�j�Δ�7�v���+%��!�P��9k��Fs0�ݵ�w�A�U>F_��X��_�y������|�o���ޠ<I4ᝯ��g���{ըF=~��������C�۝W���z�ڷݾlk�X�N\�cثvU�{V�E�B�V�)�PSf��`|=p̃HHI,�B -�_5 �ܴ��}a&C�V�
X��-����X�k�F�������Ҩ�P��;�W�Р�:p�n�
Zރ�z" �yI'��GҾ[g�x}��z��p�>�g)�uܖ;�x�t���H���,gnd:���p�æ4/���/�]����{{߈%@�~ae@���Y���p���I���C�[�7��'g�x��P���@���},�|	 06�ȀX��@�f������W�+6��{W��X��o����q����^��R�5��%��r��g=�d�@�DM�^I�E���!V�=0h&�����z� ^.G0J�3�/Q�[�����	g���
lr>wW��1��
<�#�i����( ��:�8/K�s���wsT`�}Ӗ%:�A�}���'xv=��]��C�;��ç��3������@�N����{F@���㮡����$=yXB�Q�N���?�,:�>y�
^�}�y\na����F �3��.\�6�B3p,ؐ:~f��h
��.)ph@���0�66Xc*��eCl�l�����U'���_ZO��� ��ß����o���?`�Η�@�~���?\@�����|��l#���</L���ۤ�C�����=����)o˯��~?�� ��_��FO!�=B /j���	�c����ۣ��G��r�բ�� �!�{�@��u�w8��p��}�m����~F�e�`�1���� ��,ߵ:z��[�v�Ma�F��`���@������p
r`d�� /��|��ǳ� �G�A����ڽgp�2����c�R�AƖ��W��! �ć�(m�۠����H�
ս�