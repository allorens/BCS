BZh91AY&SYrH%6�_�py����߰����aT���   kEP�      �    ֥� ���m���QA�h
;[1�kFIJ�����A�    h�z�X0
`p     �   (   �   ��n��v�g{��[֜6�=v�=��]^�Wo^�S;m�����R��� ��-��S���'����}R��{����o��{>�ws�����G�����}�N�����ã�wt��ۻ�;J:� V��x |�#�  ���*7��ٔ�j^�m}���(�������lPm�t���	i�|o{ݞ��9���zz���{� ��y��#��=:k��oA���)���Y�r��g;�yOf��I��$k�������ܷ���=�  �W{����R[.���;��K޳Ow1���:g;���u%��]�����y�q��n�v:��e�Ugw2k�mەc�G�ם�Q��C��%;��O@c�� ����nn橺[v;wk�;s����%�gEs�W9z�k��Z��ݏ N��ww�ӝݣN�ݬ��z�^:Ε���M�^ǂ��;w+Gsu���bS՘!�  vS�/=�)Ͷ�uqݷt�y9�-��6^�v�m���.S׺����{m�;��Ԛj`�/^���kf�.���x�Wm飷\�s���                  �*T�)T             J��4g��*�1	�d4�20CC �J� F	�d���	��12`JmD&R�Q��&L@0 	��� ��H���MM��L�OL�5@�@�M�Q�D�	�� BmM�6I䆘�24zOA��L5J�FC �1 � &F`?3��_�W�R�!wpb2�a���apY�������"���8ӏ��� T�Q �*�z�QP���(%����[�p�����6����Bl?|��a��Q��~��U]��TE@�N���_�B
*��'"ˠA{�G���?���O���O�l���Hݏ���7�9ӎ�5Wd��D:��L�(Fl�a;RY=�N	'Q�Q���s>�$��ü8_C����"o9&p�}ӿ_�dnT=��ȏ6J��=㇑5�Y��eL<t���^JN${nsnw�����=��Uӥ�����[��F�&>�H"%��bX�ʲbA)�H�S�c�I�͕��2�py<��䓤�G�D�����ty�_#�(��M���+�G���G�͕��T���D�r��x�W�N;*���8`�����a҈?"[�H�Ģ��h5)��M<�����Ҿ~rR'3��%���k)<__W��D㒑=��*�5�i�̕����p��D��H�ܭ8<�}�5)��D��D^Jӥ�{��~Y^0�rWD�ґ-e'��+���H�rR'���~�Y�K�;'��ßx;'H��벰M7̪;�;R��[��7�ژr����ܪ/�}�ݪOc0Þex�U2Yr#R�z#��6&u��}��C��	P~rV'�T�8S*�7�e�nJE�&�+�.)�Z^�d��+g(��n#��v%`��IcS��>��5�0{�I�ϧ�w��G$�u�~�ԒA�Ӳ#S�dGf	�eW��+�d�Mߦ�T�I��Ld����l��G$��3=<��+vg2&CC�I��t�2f5��xt�)��+%J��\���Wʷ���Y����v8ol]j=/S��;����X�G;��I8iYR�ܕO%';&�rW2c�����Ul�%�pjo&vfGc��;%��.N5)��e`�oez竒�Ht�=��=7�]�7ޯݛ9���Mڲ6^��;����󲒸��6U��S�URv�Z��Mü�·:qI�Y�Ipl�ĻIi�������'M"{D�����H���8Y���t�ӪM:mt�ea\*$H�����0|T#�r�h�t���G����'A%�m'��o�?x~߰ϱ&'��IvZF�����%|�;��1L���;ӥ]��܂_�����54wd���Na�F�&$1�bz�=�%��Np�2{�&��2l'��%��vFt3פ�vG�f�rrbF�tBд<�!�g����B�]�ZJ�D�Џ��0JM�D���/N%��ɩ�<��bm�W��(�B`�I�q��&��i�������a0�R��<8t����G$�D�f~���N�+�	ԡ��g�<> ��D�['�d���=䈘��w��)/�$����i5&�:�>FB"Nx��DLML%�\H��aN�J9"z�")��	�D��D�����>L��p���DN�M<W�!<�I=��"p���Γ�Ll�#4�8p�"x�"'S�}ώ"'�ӥ�p8�0sġ�&Q=���(~D��I�jQӃp�$C�DD�Y�Ɩ��_&�L0zC>��}�O�O�%����:$�~Ϭ�Yސ�%�"D�I����I�ޓ�ЗZ�� ��o�O��+ސ�D����|N�{Ri�9&����_Ş���Dw*'�tNtH�+ӧ}<9����dʞO^��<M1�S!�.&����cSN�a�=�D�2��0��c�����9�����GҎ��!�!�g�r&���:�K��ʈ�J�Y<{��4�=F{�U��W�4vx~�����'v�n�[��5)&	�p�(���c��F����[Q��N��N�g�����Oóx�����dNy�ӝ�=�#��#���ƻQ􏲢=ji��bt�QD�N���(�v7UD�$���TOtGg�=��x�"#�DE�'�g�,ϐGj�x�C�3��f�9���Q��DY�ʟ#ʨ����x��gȋʉ��">ډBq��*P�&��"x�AU�$&r�%�JѩdO� �	���`�L�(FiѲD��'�I�J�D}ʈ��N�(LƧH,�<q�J����j��W�A�DG����R�f�D��:A��4HT��to��DK�*p�9>D}ʈ��KZ�'y��ϓ�3�(Fv�#ͨ�|jQ$��*".T��=mN�}>A�6N����s*"���O������ݜ�`�O��.�jNr����rQ�!_2|x�GҏP�cS�Л�6�{�B�M�,rtv&�4�aX{�d3*<����ڈ��Ʀ�ȇ���d؅3�$&C�'��(�`��<7�|zl�d��x>�}>A���>�S>�r���ߑ�c�����i�xk*#SDi�Ʀ2{�O'�;��'��S�~M,��I9�j|�|��/��!l7��8g�fS��un3�$�{�㑽L�/X�V��5ۣ�k_z5��ַ�Gw�9�K�䰲5ʍ�G0��9�I�;&�N$7�+�G�R�Q��_T��+a.�g�W��Hi����v{�MK:O[S���b�śܩS�*v�9I\K�WSZV���3|U��R�:_�%ܻ���|�u��;��}���c�W3&[Pس�d窧$�	7��T�#��Ol����#Q�r;�)��Sѩڝ�K��5�ϝ�*�zN���G�Q��}z��s�'�\��IGi�~�桑���&�Jȕ��RY�8��z=�;ڎN���z5;S�e�Od�y�kRɭC	$= vNUH7U0{u>{ʝ��꥙ݩ�(�K�F��ɥ>�aꈘ�R"'���,n�Y� ��!��1�������]8<��d���,����{�&=��~�ty�_#�(��M���+�~D�)�D��l����X���DE��*�$rR'q��~��l����aD~�<[�H�D������H�nR'��ȋ�Zty�_%�H��J�>�'Ra|e}_7*����4�aF�M:<�_?,��8?"u���I�9�7�"q�H�~���Ze�	ܔ!݉��bq��KvRx�2������%"{YXp��}89>v&S+��>��!r#r	n�xL�*��jV������0�K�G��Ļ����L쮉��a�����,jY�*�z%P�û:��>���t�A*�JJ"�}��!	�D{,KrR,�7Y^��."&�ӻ;�Rl���}=��~ϼtj'�>��5�W���D�ʪL�a�C_��$�;"5<vH#��2�̬8{d>G~�9UI�rV��s�8�?'��Ϡ샟Lɞ�2<�[�9�2���~/��OA=�l�eJ�R�*W%"s��em�<���K=�W����J��U=�N��k�]�~��{�c���������S�V�S��Jvleg.Ul�%���ggz��_4��*�KR�V��Q		2%����,S�����N��0�G�E����|S��L!�J�*���W�E_��9�o�8�b#ps���Z{��N&i���:V�ߴ���<���+�e�w2������/�D���t��?��O�����O����gsjX~
X��J�2����;(刜nl��\�'�qg_�.�?��Ns�#x���'$Lpd�n�z�v�ߢ-{4ח��ήo���g}��vq�=xzIW>���!����//{���R�*6��E�}n�#|�|ú�^]�9=5|����{~Ծj�޹3Vq`E��<窭����4톶>/��.l���.�k�����}�{9��Y�E\h���Oӳ��K�G0Er��:���}�
�u򤭗vy%�?>,�AoU��]�l���N�L[娂�x~�6�n�>q��$���������x⍌f�ėN��ζd�J�w�g���$d�����~�]�}>UsË*%\�ȗ�e_l�h�ö���������sGǄKx�V�|���.���q4�Jn�曬��]��9{�����U�}�}�n�{G�Z�}=��ί��?0켿���_~]��8���U���ԕ����7�{\ִ�VJ�;��g���������v��i�m�țz{n�Y��k���z�w�سQ��?_��_׷��~��Ǉ}g鴨|$~{���˦��G�K��i���U��秛��u}0��[�o��/%���${���_9!�F�\��<�������>���ӷ`��ˊ��>�t��׺]Y�5����xz���\ʌo�W��.���x����{˜J�Ϲ��;�����g�:{�_�}|�G�$\��ݣ��g�qwé'��>����{����~�o凒�>����g7���|�1וDq{bw|�{="B��YO�R5�WV���Q��������sg���5�$eJ��\�ΕT}9\�MjI��u��fS^�.����%��'��JH�I5;�������!*�&��ł\Mj��ލ5�Y�A��SU%��E�������j-�z��bc�*�I$����L�t�w~�۫Wzj��������5��\N�$�}�SM~Mj�qD�B��U}��ė��$������/��I|��f��իT^/^/�|�(�TMyuj�:{�s̫����m\2�Ýi�s�k��/ɞj�+��q���yge���>}є<�[�,�c�,:��^r�����WB�A�
�x;OM��r��ʁ	O������)q�5�s�)�I�v�}�����3m����Y�!�5���gôBu3�jK� ®W��I���Pf2wY˾au���MƴPmI��r�
h��s�h��h��S@��4XmZs�7�~Xo9Vc�g
NG\(5�yf�|V�e.=�WF�H��Xq�����>q�@��>�a����"�3�e{��c��]A��<����C�:����~���Fk�������Ǎ}��B�S9�-�Vt� �;�2A�<5g(�X���*��H$%�NL��l�ȼ�'fTgy��_9M5��Q�Yu�7��f}�6�Y�?�0���F���5��׳ƍ��U�`l����<������Z�w0�7+!S�8
����,8���@m���nF�םM}+p��'�i�%$=ߋ���l�J�gx�*Č�el�}:*��Q���x{�������3��VToY��C$}<^i�����4����yj΢|�#���;ך�Q�οC�x�5���%)�����k팕p�Ȩ���*#g<��Z�ו��<��k5��s�,���Y��X�������R��uf%V#Y�^3�|�{���Փ�ee���k5�"�Q�Of��lϽ��icK7�M�?,�?4���~�p?,܇\�f���x����9N^���Ƹ��qaհ��F�^��yug��<�.$���˫=v��g���y���>��qg��[�>����^�r(��Y��6�*�S	���w�տ\X��(%���<�{�`���z�V�I�v{�O��)�ig��Z3ߞuj�~g,��#V%�t��g���Y՞YՁ�I�nقlgvg��Ǟχ��7�f�����6��.,��s���sz������fo�|��d�i�� K'd����s�|��ϼo9�=m����ǹs
��A�X���Mi#�����#|gM�q��Y��|}�n�g���M��z4��&J�������G|���!:����if�h���n�jk:�9��u���0�ѝ߽O��w�M~�w�k<�Ig7`��Gҳ�yDE����&�\�Fs���ʒ�x�Īȳ	��j&�ci�qLIj���R�(����ı=���i{�}v�,I�K�}�t�Jl��Ұ��ŉbn�H\t���SQ�)��s5>�=��FS2W!��\�ԩ>�#+��&��q�G�Vf�߫����?D.?I��.�u%�r�oJ��yg4xyV%�v313�\���:�-��-���U�u:kp��2���z���]h5	ts��;�,��j��S}*�Q;����ҵej9��F�b;�\dj:�cQ���J���1���1��n3eVGVugP(�׍`�o���`��.�(�w��n9���&�cT�<�%d���N�w�v��&�Ԭ���vV�0�NѧC�+�*J�e�̭���4�j�s����<��E��]�Y�^\5�1#�]�mȋX�'VDk�|����Sr���������aj��M�D�f�j����d7ޗݿP�Q�Uvn���X���]�|�BZBN��{l��\�%zS4�J�/�v��&y��N�+�]�~k!��CУ@<p�g>��r��yX�2#��C6�}�o^U�X���Z�皋�C)�I�jtd�ʹ[���ax�P�����#ZM7ֻ͙�;���o����5�-�æ��Q��gV{��Gԑ=�x�3�J�V?h�#��I�<h?a��~�����o+r�O͎�!�X�I!��w?���ͥpb������;�C�=P��}��3��*�⛸=��N��s�rv%��@Km6P�a=G�H�!9�v��$#�~6�|���o�/Me]��q_"����?\��C{�T_�e&��9�� �fsf���l���A�>M׶_ged�J�h��n�i&r�hԦPd-MuS�;LՎ&sE�����Љ�d��G�,hꇺ�%u%��6|o���y2�/�:]�D��+!<ԕ�W��{F���/�сj>O[[��R�j�h��S;Q>D�\2�;j��mkR�ƿCD���^��|����8�ǇVr��'��q��%c��X���GTך�u�YQ>g��8t��
�����zr�U2&6���I�l�wi��v*=hO=�7��>����gS�����r�Y�Ó��{#ع序!��ε�Ԭj�]fo�����'�C�O������?G��O��~�����K���~���!^�J��X�׷6��'x����J�ۼ��&��;��l�vǷ�˫�w�F��>�����#��q{�ϸ+�Zs�}�7��b����{��f��rsxu{v�����^���9�Y��L��E�����[/�W�Q]�-��ͳbH|�-�~5��V�;��s�ᯯS�z续�}���Gk5gT6�S���g���o�����[�r�ڮ�qts�|�/y{˵��ݑ��i}q�WcD���q���z���뽔p��{[�{�O4�7I/B�K�ޤ�|���g�ț�W9��𝧧;l����)�s3�;�f]���7��s�䜹�7��NݮEkd���M��{����u�rjK�λ9���j���]ȫ9�D��:��Ayg�\�����?I�U�g�ӼʙF�w����ޒ�
^����U��W�9�t��{xsy�y��==^��QSL�=�I2zڻ��v�eQ°k8p�/}ߘ��~�|�uw�ȝ�>]�Ow�V<sn�ޭ^�2��z��{����n�~WڝԼ}��l��6w�t�|��5�o�n����W��m��~�S�X�~�ͽ7��<�W�98Q��Ԕ����ts����(�MT�����?_���%�C ��v���۽�!���a.�rƲ�6�J�D�1*�Ri��Y��CElˮ'\�&�Ci2��(����O��8���A*�rTؿĴ��c�f��n:�J��Eq¤�ur2+�<��*+�*��D�,��]a�H�uF6�&��x՘�Z@����d��*��T괨7�X����+$.��^��m2�6���-PQ���֧j�QQEc��q���RV�c��!��[
�!E �<d���jZ�F��Ǒ��:��M��v[*I�U��^�5�5��_c�,ČmrBH?'�lȥ��tnF��K�ړGVj"�m��R\ʎ��2�uE>PXj��L�:���Kh�w��S<��W�%�r4)��	 �Ě�5��))��l��ʬ����D��q��,�qm�F���x���������B��,��gt5Mms<�b䁩#�۶�+b,���]Q�k@���D���e�dPHA���*�J0����[��*F�2�yDq^<K"��v��dY#^�]lF��8������"�#��	 �A$�\�u�U��D",dI��5R�0�e�$�b%nڹ���[�+���*�֐Ղj�D���Bl��%T�ė�h��$&�YP�RXH1w�~�c�|�u�am�%2��׮I2ڣh�Ւ9l��<�(������Ge�F
(��&Z�phHB�"K"J�#Ĭ>��Ө�f���qĥ���MTӹ%U �*1*�y���1��uƃ�*}�E���Q$f8�-�ubA���5��3%qTs��c.,�^TeZ��Y9��.4j��T��/�SS0�c�!14�afc��\���y�b?m���+�Xfu�0�u��fa�E�~��.W���L�$�;�a��`YԄ���#�����^h����,��A�1�B�nD*Ǻ��Q;�C�d�S�s7v��bɘ��8�b��\M�]D�}�3��v�v�������1Y�F@w ~���`\C0�y $C0G0q55�733ķ��W�C������(����z�?��۱�1�[���V�/w�����~��|�v{%6�����������1"������3�����uU]b��-*���U\ZUmU��U]EUUV�U�^*��*��*��Ҫ�VեUqUZQU�TUUu����UW�U�V�U�UUu��������=U^�ڪ�-*���UWX���K����y��1I�N@�*2,�̬����6i6�l��L�iXV�M��Jr
4@�dQrv�9�{������*��*��*��*�UmZUW�UqUz�j��[U��b�����-*�U|�*��Uub����UUUUqiU�W�Ҫ��UWV*��{���UWX������UuUUW��t� $E$T�QH��CH���,�,nFZ�+51&��[im���Ak���|��U򴪮*�U|��U��UuiU�W���[UUťU\ZU^�گW�UV*�UmU�W��U_*�U|��U򴪮,UU�V�m^*���U�W��W��{�UUb���J��W�Ҫ��UWp��O��'�Bi>��jVQkY��Y�ܵ6�	>���B{��߽���U|�[Uz��U�U꭫J��*��Ҫ��UUTUUTUUťU꭪�U|�������J��^*��x��U�U꭪���U]b��W���X�U�����X������U^�ڪ�V�[Uz��U���6����7&g-����z�������0�m�f�cu*��n&�Y��q6r�,�յ²��2�rr��V��F��[����������w��u���v��Cف�����O�~��d���~����!ӧN�<"&��AN��<xL4D�0�,�A �$�
,N�<'��D�MD�0M4�����DD�0�$���D�&��d�tL:'D�ç �DN���'�8 ��"x舆��`�ı,�'�(J �#'H �	��$DK:&"hx���x�Rt��B"0D�Dât��ACD�@�Ht��So�iH]9��8���]���

N�!���nZ���QJ �8�U����J�9QAEU ��IEq�b��-������M�d!��R�n���V��"5�B����B���e���adcC*��1��bn�!�,s(ƅAc�}�#q=܃���������$RU2UXVGGGP�YQ�E!RI	��+��:���q��hX��2,�b�f&ư푭�Dl��bD*u�L�ɔn�,i
[��G�Աh���tc���T!�e��,m2��N[X4XX�XӍ�q��d��Z�m�[$*��mX��r�ދ%�h`�Ur��chX��h�����!�H�ƞ���[�0de�NV�H�d��4T�r
�eB��Ƣv�����T��I
Ŗ��,�Hm�2��"�+��E�`�x���0�Re��E,��"�b��U�G1��Q��J��8�Q1�	I�R:A3*��T��*�u,V2��ʤ)��d�2FFD��J'A��Ҏ��x�7q�dcR��F'�J�5��:�v���<U����HZ��"L�n�FJ���V�$��H�	��tJ�A�V�U�#]��
���*Lv+����!"Dq�D������.5��-�X�rL���B�R��FW�2&Qb"
AC(�d�y��气�pdb)��R�� �\���Q�����)�2��
�J��Q1�t���
 ����
�2�!Lu�
�Wq�;G�"�	jm�FWP���HT�!h�Q��J��*R)Q؄!�ǒ�ȊZ�[dYiJ��DVT'���۶	5q�7��QQ��,�7�H�l���xZ��5�V1�ME��H��e)0`�lN�(!�ǒ2��2Bұ�ah2�QQ'T�vH\���U�$	j���uq�.$&4��(&�S��x�p�I��2�'!H���[f��w$��x�Z1H\���c�P�c˒�aKd�B:�E)`�ˍ�౐lR��FD2QA`��V�HC49G��*MWm�:$&�AR��21�*##H#�㖥
��qH\�c+n))!X�E�YT�c(��6A2!̘�bV�l���D�y	f"+#��T$�c��Q[�2�	�]���beR�<O&Q�c!H�b	FYNYJ�	�
�0CjR�8*,.3�q��i��%q1MƩq!#"2��+q�JD,,F&UZ�6!�SJ��F�((�"����F!º(Y%v�V8�Q�P��RbR,d#©r	�I��؁��e,5����b&N�
��@�Q!8嵦!�TBex�@�B����#�&��Q���!A�*�TP�BTb��X���K �R���DD�1C# 4Q�I�#�C�c���*r����H�7m&A��J�W|�#����H��bTI��:��:7J¤�IY!c�+�u�&8��Iք4"�IE���[6��EYI%D{n���nLl����ڊ�"r�d��$L�*M1
9]�$�6��n�ۍ;̔�4�b�/0n�I*f\clJ���%bJ��b��:��*�UH�%��n��6�v4��T�S%W!����D��	�q8V�ڈHV�ݩF��e���HE~D+��n4�o-PHi��-��H�l�<v;\v;�[$��j7��\N��S��J�rJ�Nښ�u!�Q+*L��c+E��q�G%�QRԡ,�JVZ4�R1�J�d�-��.����BF���i�J�&9b�*+u8�MV�'U��q	�*�ʬ�TH)
�u5Z!
ǉA�*��c&5bd#��W5�F�9�T�X؜�i�N!E���»��6�p�+r�A�6�H�)k�dj�$�q$FӪJ�5mWE��d�I:DY"v�b+OV�M�G �e���b�F䉹S��eRZ܂m��+��
�Q8(ԈlI�և����%ie�����]����)UU��r�P�*�a1!<U�m�UibI�BW�Q��G�	$vGl��Q��V�X�u�+V4Ec��dc�	����B+�
ՉQ��v��v<r��H���,��Kq�T"�F䕎E�7Gl�*5rHLVʡ[V�Yd�*!�&�I2������kbc$���6KaEk�\C]rU6��K"�jF�v��m�����i�b�$Q�p�ʺ��9
�UrW*^�O�����*��*�wv���>�[UyZUWU��� ||�����*�����ۿ���mU��iU\X���ֵ�ت�E`�����[K~�"h�'��4�8ѝ�BH�4rA�<������SE5�	Im�b��Ȑ�P���I�����Wku!��.$퉥)+*X�i�c,��uXF�-X�P���[QiE!R`��d!J�C.J5�u�E
�U�X2e�8O
��H�c�': C�k"d�GU�B YJLR�p�(ŪBj�I�BcC��� ��9r�6�Z���%��(�V,���R�F�UE�Ab2�h��L����D�U!���I��J�	LV�Ri�)2&�Q�,�t�h�d�� EX+ �*��mU�GSn���B���Z�����i�b��'�m�"DE�*\n�$GETLm�I�)-I�I*rGYPܣ�q��J₲����MX�ȔE��4&�l�B��hm�P��)	%R��J.׵�Y`�d�[rK*��%�[M�!Q:u$�S�7���$���|�:vF��T"g�#�s`��*s�㽜r�Ht`�ӄ���w�(t�k'z�[+i�k�w�G:{��.>sƳS䕏��<�a	�Zן�d�F��nQ����O�L2:�4���K=UT�
�i���98V�G���n�l�t�/8*��gj�Ѫ�l'���s\+>����M4$�����r�$�����>W�0���-�${�����Á�t��F�����o]�r��HI��t��E5��~2=�x:6d$u�a։��ļMZ{J����2�8�_�y�����D�4O%i<p�m�J��K�LorI$)�[���8���B$��{�w3��-)Gce��!��W����V1	>�[WU�v��:0�J~9p(����vݑ���H��8T���e��I���jM%4kխ�{�盞Gt��e�P!�81�jp�!J~2Μ#����4iu��y�r0�D��L�vq�q�M+��O*�am��l�M�"h�'��4�8Y!��u�@��.�X� `K�q8��Ȅ�V`��T���He<$�����`�#%��h~$�[�JaUf�m�㼸 Χ�:��̔[�a�ѣ�M}g>�����m���c����I!����-������Rϩ��W�rRL�lp����%�����c]�zֱ��JC#��Jq��Hƕ�=B+��F���F�g�f|��·�b!��p��OǄD�4O%i<pݽJ�r�J�p��I$�f�&i��$����y_j�xGȬĤVi�eŌ�Lr�j�?	�8[j8[k�iI���{�L�~g&~5<M���!��m06p�`v�0���6HD6�c>{UUN)���Fdٷ<��<^���3��_!�CGNl��2�ޥWG��u�dr���i���նa��ˌ�˭:�ͼ�μ��ç�<xGN��u���e�#F�i�Ø+�-aor��Dk��h��E��q
�U�o�4\�BmÉbMH�v�i%��i(�E\K��I$���&�]�];�|q�-�G�s�>�7~4����6��^Awgs�;�M�:�z����+e���g������ӧ�
:i]ӗ�i���;�����~��;�t��&[�oZ�i8}��{�'f���W��:���^��Z�r��d�{�p`ލ��GCj|h�s�ð��Df�\�!O��2�QCa�08bfn����d�Yq�3���4Έ���}!
�;$e�s��
/$pI	[�&��D��d��c�wL�x��� ���AO�&%��曑z���(:���c��L5'�C��f��PJ�
���,Θ����4�����,T<|"p��,�~�"h�&$4�l��UJ�J��0�,�nH��I$2�ǤN3&���3�
�QKW��n��\%U�M���/Źѥ#�6}�:���s����MbM>w�N7
���%S�J�	�~9�Mg�Y�<��Z0�÷]뻺�A�����#���CrBI-��5�����Kݭ�CG6Y��V��<�μ�Νum�Je�2dY+fD$�yS֒I#��%B�ǐ�:b���d~!ё�ւ��W����=ġ�Lc$$�ㅼ!�)��0�s*�N X�F��>��dz�ٌ��e!DQ+�ݴ�J�FB�ЏD-� Ӎ(h4�,�C��{&9m2C���r�N�:[�D�n�ђyK��$a
��г��Ġ�T��Ѵ�E�>G�e�/4��m�u扂hi�0��E&sn��]s�T���wM�$�H߱,S=�4f�J��K�Ҥ<h�O�l;��W�n�uL���4��|	w�:\�g�.IX���%@�	Z9^l�C�|�#��<�v���r�j/9�>O�ε�$+��7��%��C��O�nn�F� �7�0=\�~bd��ѝ���۪!�˞:}�d
C�<X�'�D�4LCM!���]�;ź�;jd���k!��"2!����[�7��yɖ�Xp�ڂ�g$�X9L�:�j8�����ԒI��]�����D�7���gd=:l��vO\M��V���ӧ��=IK�9������4�Q�w�g,��ѩ�Z!r	yOa˽*�_��n!��}=��g�I�(?�y�k���ﴩ#�zQD���]۪� �H`roX)���p4��|&F�?B���k&qr���:���=6t�_���v�c����F+��qX<�ju�&��:}��fM�8X7~��Qe���f���y��Ι�8;m�_��tXz�Q^�q1��ĕ�$�kaq����S>��"�1�1�!�	��J�:m)KÇ��=�3��aI2�����]fO��$���F���ӂY�~<"&��`�<#�}������m7Hh�Ʀ�PڒI!�2c���)���b�E�3��d)����棊(�!~3L�L�}b�E�a*�:,�QʭY.�V9�A�I�|G'�I'�;P�YS��+u���r(�nw=X���W�Ṟ�&!�xI,�������>�5o�����a���h��p�5 �O�hߏ�<�#�0��#������M#	��?1l�����ql�Zylm�Kb-�E�ů�g�cI�W�-<���n�M����fKb/DZE�H�H�d[la.J�h�a-M%[LV��R��Z>[Jݦ*Ӊ�ql:�G�ao0��v�n���[�-<��-�O-�'S�|��b��l����ť�����a��[ZD�Kei�ZZ\�bөV��'x�ܞ�<tk��2L ��-<�̘�ش�������a,�<>?�?���N��~gG�,��bx��O��l����A��<8OČ%�K������d̟�D��Rފ'�OGމ跢�-������V��㘓�X����8�6�N��<0�'�g�g����%�ǒ���|�$���>L�lE�TxR�T��	�I��ÏB�QdYI�|F�eO}�z��P��G����Z�H����N�{��~���8���m��I���}t�ܜ�wό��W�c�pR�I"��=ƣ�|ka�5��]s��m95{#:J�Ž�!����Rd�'����V�����|͞�0�p�i��GR�C̢���s������<_�U�fx����M}�����z�����~\���w]�9+�E�y7�Z9�����Qs������a��{��i�UU�w?{�~����{���������w�|�Ew�������{���]��]޳��{���w~�W���~��s�����ww����Ux��X��v��i4�]iխ��yםyǝ:��u��ͅ�oQQZʅ`W�;��������9,dJ C-����ᱱ��*�r�� �`��}�%���l1`��+Ln�D�"|�r��AȦ���(��bMp�	�M���T�ӆaw�+6W ~���:h�!�%�/ŖC�R�X6ݖ'S&H��ń�P�d�S����$�d� Q��@�
�J2�6���[�4<!KA l�y�X`�V�������ti#�-'Xf�	OP: ��ϻ��e���n�ي8�	T�=QI)�!��Uh���<ˬ�4��6�:㭺��Vî2����cY˕�Z��**+B@,ʰ¡�;)�Z�J)v<(��`��J��<�=�hO����������Q�֔�\᝝����E�3��2󎛪vEns���{3�:&gL�鉣�6�j*�x��Z�Xe�);�T�x:��BAp�
²`u#�"e����PMB.�L4�*����+zwU�e��'���L2$�rSP�8�	1����9�P(���*F��P�)�m�?X��nM)�/�IK[|�HC}3��R(i��E}��� d����0"�T�V�X�ꢛJ3��R�ӈ�̼˭<��xDMD�44��F�s����i#��6�*���6G7k8�NH�\��YE�4�B�;�:��Pi؛�#zԵ�X�+JZۤbS:�b���$s٫�������s�}/ݜ�Y�2�����&B��z�*�aF����:c5�λ�*�CיX{3%r�2�&}1�'M�8p�߸zW��e}3���=9+Ǫ��}w��=���g5:�����8N7�Ϋ|�����9��}'�mq��lkS���[pZ1�r�x�� ӱՏJ����$� <$��xL�1��q�����Vd�q���Px0\&a�)�����@�N<CF�"Awd���� �DI�2����r��0��9RHD7Y��8a�G�
 �ye�8qՌ���<�Va"i��+(��LNn�	�#D6й ;<CHY�[���c�H�y~�GfJ��A�Ev(�
 46�����쁌r�ŨI����W���VU�J���M��oF��ѻ#�:i�1��h���5�l��"�J���G�u�Z~[�o<�:�ǃǄ~<tfB���9&�R�n��**+B@��
�BŗM�-��#���q�����#UW0��dI�}�����00��&!0F|n�'#?�ݹ	\Ƥ�w͏ʜ^�
"����!��5\�Ѳ.���5e&�% �!7;M���m#�/�M�֯=�v��SՉ����R���~�:�U�%������p�X��K29�,a~2���y�E�]*�4Y�U�C�>0�FI��7���`8an(���!
�p�3��	����r@�A(��Lw�`�lb�'0�&.�� :�RQ�:J���T}A�e:FeW8�e6|�8�/̺��~m�&���hi�0�C�����������[����y�TTV��у�z%dh�2`���N����tB��N@�����E��F��i�Ȏ8 XA�����٬���IN;-�C�6��\2>T�W5�8�`�b	�{	NL�t���N8(J� b�y���1:�(����R�bj:(/��j�4Z�,{��5��^#&������PeW��J�I�դ $,�d?�[�5�}����2b_�*��	^+iW(>��)��$���Z"P�$L]/����QY�1�l�aF�S畅o&�l�9��x-aM�4F����A��n�n�8n�ѡ�����0>#qa�d�|�l�\B�Q���FL�h�-�e�5����p��2�/�ϟ��m�u珎����ugDbO[�dƤ�n��#w�,w����	
��?r��wĝ�)j�#��`���i�a�T�1N#H���4eqws4A�D���Qb���b���&Ic�g ����(�a���
!���j4�mQ������`�"L+Q�4�Q��l]4fB�� �9��X(��t�,B���	�C�\��&2�W��|�"�J|!,grn�˻����'6���QL�?+-1|���f��d�i�R@�	8`��å�0�4'�hh&�&`4f�ي�ֆ6���>�wUr��8��+��Ȅv��0�05Qh<��YEJ��+L�0�6���/:�o��4DLCM!���;U�F���}<s�:)�����y����A7�i���e�ZƷm~����C$���Y靈�m���()[e���3I�|�**+B@���<�����Η^?)|2������9��~a�<Ow[9R��۳U��9ż��>D6���oy�~�b�Gߠ4�����v��1wy�^c�{]��{�}���G7I)˳�8�(L5GGO��B����0���)�.�$�4�lnS���[�$�xҵ�Hɹ̢v�g��`�-�e�h���4i�!G���l�`'�:�j$�̥�:죭r8#�$�� �*l��C�)f�>\����P�� �6�h#_1V�A�i�ޟ��)�Fa�q �|�i�%!��L�l2C$d16zBHP9 �E�0j�*!d?U�M�;~N� b��o�vT�^��B�f馊7+�ak��������Cr��J�|1M�0A3z8m��*�t�|e��<�F�#�̭��_-���yמy�hi�0�a�6r��v�ޗfJ�7��r����H���(oc����MYD섖X���_|>A�i?S�J}?>VZW�Ds1������h��6�������"��L�p��&H#�4��i������@��!m�������zC�S:�ۓ�}!�?P����0���OFځ��Cf�.��,i����-d�[���M]hyn����ܵ����)�sDcfCd�dhK:���#y��Ն\�Ym������l����g���*m\�>`�J�a���|�<�BS�:S�Hu��3!C'L�˫|����yמyǝ:�8���tX�nE��\�˗�1��7���� �dW�LG��P�-�A����@���8�&k���Q��l�Q�Ң��Oq���v�k�Zx��#�A�)g���t:䤚%
���rN���Ҙ@��$�|�7i��}��_c2>���\8kz���i���oe��Z)��p��B=�#��4eJsC�N�C�0>w����J \e8&��l(�`�nK��� A��0��&Pڐ��\�bba���>|��p�$3FÇ��!$�1в��ݒ;3A��@�f̛F�e�][�6��u�q�N�#���慠�OjDN�m�|B8X8Z�'4h�Y�c�0A��6���UN4>а��Tr�|t�Ep���VUl�>x��� ��kkI�j@�?�?�\Jȕ�;�������4�I$�vm��l�4>G��&?%1����'���xlK WX�Ppr�]��e	� aP0Į
>�`�G�(6@�ջ�pU�#��zd>m�:{RG�m���d�,�Da�"��YP�R�(�m�A���nj	�B)�)	�O����r��>���`p��p�b�SeR�p3Q�Uݽ�"i�Ϸ��"� �%2���M�+D�(t����'��xJ���k�h�&�C��]��-�d�<|>'��Ʈ#�C�il�2�ZmlY-��KKy�V�Ƙ�>L��K"�I.��H�dZFش���F��i�����Z4��Z`��|�-�Qi�:�V�y���Zu-��KO-�G�Ǔ�1����b�[-%�ť�����c���Z2��5h��LZZ-�:�O-��mlU��5%��m-:�M���ZE��[+f��Ӌb�ǒ�c	dZ�Zeճi�ص�i���-��D���<lL<5����xp�-�l�b��	i$����Dm"�Q�!�Q<G�|M�|l�Į���'d��c��~����~O-�f��b��^e���ش��Zq�--l>q���ҾL��K'�W�V��O
^���XF�T��|Bɜ��N׹���^{�p�^$�S�7_N�|�����{ɣ��'���w����_ܫ�s��sa�>�n��r4lj���6{_M�jsw��z�=:q�<M'�t�uw�&sy�s��rww�pb�Cy�B&�p���?#��Xq�_��N�ƴ����� \�~�qg���y�^r��s���~�����+^�5Qjb��n���i��:�����ԟ6�v�sK�4���,ĩ֕Ę�����6.p�
����F-��9��'͏�o��qV	�m�Sf:B4S��"^�'��w��T~�x����<�s����rw�T�￝˺*r�m�d?p©c���~�3�N����v�y9ᴸ�|Ś����ױ�����g߹k�q\����s~���'�=o���|��v>���HI�}>p�� �!H�#YR�(�e�V' �U$����-��6LV�+��&j�ƣ-��݊�b��M�ښ��6�b�	N"A�6�܌r4�6*[UM6�M:;�v���v�j��_�r�����}\������:��U򴿻ۿ��n��~�^*���������ww}�����U|�/����v���w��UmU��{ڿ���eRa�u�Yu��[g�DD�44�~0�;'Z+���+��HZJ�)jV��1��cu	�,(�+S��;RNԔn,�i+ZiH�
��<���D�*Q���ˌQْ�1�s�qD�d�!4�j�1��J'�t��Z�����B,������D�E�F�"�ڊ��!a���]Cc#=$*(�QLB%lT�er�k�Q�"���	!+ ��K!DR8�Zr��N�G$e�-�$�,V�JISEK8�9���y,���ub���$��(��2��2�d!bH�%��p���al�.:"�L@� �hM�4+!%M�c}?�*&k��1Ek��2�,J�2F�B�I[���F����H��Q�F�,MD;}K�J^1��ܪԄ�!1�[��R�+�QDJGcw(84D�i�$#h����CI�U.*K*v�T�q��+�݊�mn�IJ�HQ�!lp�y"v��!a�JX�%�%N}���1�`$�w��؏秹Hp�?s��_'gNp,᣹ɇN�ٓ-j�;�2��0�^ռ��h�S]+��*�[�}�����qnd��o>�F�u�w����l��}��|������s�h�)Jl�����E�Y.���^���d%X�;,���9h�n
=���UQ:h����ܹ&�k��E�*����47��gÌ! #�'2��>�@��2A����0���QQ>�����{�K-��n�>A�C�X=���!�����d�̓C�cA���e�+�
��-?>s������&���E6��-�C�<���%��1�@�kx���&����T�d�rU��)�����	��Z�V-���~9�8���6mvm���#������1����$&S�2�����r���� H�T��V�p��ĭ	7�ID���>|��i�^y���g�DD�44�x�}�jI�*=���c�0
�M~,�ŶӃ����m�1�Ƹ�P奮i_�3QZTj*>u��>t�	��B��A�$) �
���tB�:+՘T��P��II��#(6A����c f,!�Tz�-�p@ ��P�I��a�VR�U��PwECꄒ���M����4C��(�	C��Pm���]�J9C�ko�8x�f,�3Ю�L�0��`{˯���l�C�vS
і@��q�k|M���*�C$<i��qocia�$����Q�d衈9.v�]�T&��Y��:���h��u�[Keoϖ���M��Ha���v���|�(`�J�.�ZS)��$��Q�c�H5��Շ�GH8SEj���hs�d�
�CD@��m�(�G$l�i�# �ÄB�G����l��&��zݻ�[��I���%%�)q�3���A�Z��n�nZr:��k\i�}Id9ʷM�w��a5L<6����#Qq��.�9��N"[=n�kqd�P�d����09�� x{�Ύ�}&6;�cNe�Q��0�s�%Y��(��te��:Q���C@�2)�����3����|f��):���S^$A�~G,L�iz��l�an�(�L���ӌ���~mkyמyǝ:�6x���ew�^&.Mzv1�c@ z�<���l��Fu�Fa��ӗ���I��k�6�wp�r�N�:i��f5��4A���$�/���C`�!e��\B��F,��x��<�8C QAf<�ܤF �b�5{��TChD6�ƒ�JJGq
r0�8�C�~i�A����F� �h:n9�5�q������B�Q
0�'X��-��|�n�w��B[CeO���$$(.F�)�<Aѹ&�L��#	\b̙C�fJL��٬(�r��/J�L�EVL��˧ S���@�D6�S��#!���2��`�\9ba��6�4�N������ַ�y�y���8~3����zs-֊!(�*�m�Xo�)��7������b�b/M���N��
�cIk�'�#�*����e��:Թ�dc�0(�����>��K��������ǸM�����f1�9��xۺ��{�Åot�U]�9��8i	�I�a�΍s���w�{g�׺y��M�۾�K����wy=w���GH���l��{�3�T���EKƍ6k�y��A��')�o��!�`���Ǚ �����Ɏ�eD���n�F��H�6Wⵁ��>��UJ���ϋ8�4��|M�o�rw�Ҹ�$S|C��S_"Ճ���MT�R�8�Xh������F=4��I�٧����,��X	y���t��R����A���> P�^PY��c-R�p�/��i�~aQ�ei��n����PY=��4�4O}MN9̜p�2Yc�`A{uZ$"��ȣv١���lk�I=5�O��K�e���v�rCᢘ@���#(,�2R�D=���ӜI�r�J��4J�F�<��:����ַ�y�><<#��{���)#���u4�U*T
 �������_n�L#7�C#��MA�v�zP�5L�&��\�8`��
+1�?�A���,��qQ4�R�㺙zpK�G�G=6[�lc�KK�C��%q���ME,�K(ccP(;ad
܈H�N�к�Zj��M�8tmq���$��4�e;+.��iɡ����i"�!��-i14�1�2��ϣ��'��9F9Ye���1#!���v���E���O$8�G�G����	�`�@l`�$��hq+�|����U9QO�1X�wZ�gA�� [���@��h69�6�wD���M0M�����_F���4�N���������^"`�i?�n�fO�Rr���r���L���]�c�@1�y�D�qi��و�t�Y��R��dH@���A��ˡ8B��������)ǍӫB��v\,��E0�rA�{�}	��������N�4P����bQ|''Y2Vht�?��?�Mnd�^�
,��%�WF�6S�-A6�B���T
�J�%a����d��f���
������,04A0�F �%c0�lh-�@X�2�#3�A�ͩ�n5�څ�Dh#4�£ ����k�Ӽ��N��d�;��n�<��g��}��3B�TV��H��;+Q�Y5Ph��q�y�^|��ַ�y�yӮ��2�ߞ��EEUQ��1�-c%�s&F1�c W�(�B��C�?(jA�#�&��o�x�3�$�4����Yݭ�4��,k�"�i�Cj� ��)j��#e�#�a�f��Od�P��*:!����p��XU���3H#���*�Ɛ���l��i�解��a�p��$0<�a�hÂ8`X��!��CuE��-IU�9�^*����d4m��t��ҙ�ٖ�4�$�I����@���و2Ɔ�� ���D�@d#y>�M�924@�x��7Qب��jɚg��#Q�O"�q�Zy��~mkyמyǝ:�8�|���{�k�aĤ�����mpj@�Nn���9�7+�����w��8ҐP�Ց����Y,�!��=�1��<_ەϧ����~��;��,ӽ�el�_rt�p_i�>g���1�������ig��>�m�bߪYOo��������ӓ�5��7j�=dޤ�{}μs՛���k��,�*�W�q���/���`�C�:�L>;���Q+@���K��8b��!0��a�!�C�b8,o#�Ad,\߾�\�B�HT�Ji��F������81_�R�������9|�X�*���pt��4E���4�l�283$G��i����H@��w��2�A����@ȉ�0���p�n�'N��n7�8���q�r�lX���`�4fM���Ѻ/�Z����m�����܌k�ӓN<�W]��45���!C�5�䰢	�L��	�G�5�-���q]~~$j�+�3�u8�:�m6ӫ|��ַ�y�yӮ��/3\���A!�r)�u�.�ǆ�.&1QZ��C�ϳg
�_�p��"�~6S*�:�<sTq���~K�O��%��w�����r�g��[0>�lk��J���2@���a�C&\���@����^J��$'ORT����(q�WyL�� hh��A@ă��Yw�=Uь&��cQ�(;ǃ
��h�cz2a��:���-�G��MkE9&���� Xs�,tl��l|���`��M�٪�w��~�P��ؚ>666$j�C
|t�'�2x�$�>#��y��ť��k̶--�-�%�g	iů+f��kb�obey��io0��[FI��Ix�K�"-",�i�"�b�KF�H���-��|��Zah��-KGVè��U���m��Ŧ�i��-<�[�[̺�M-�p��[[Km�E�������ih�Z-���|�0�KE��R�[�m-*�r[|�䴴�m2�$�e-/cKcKb�iin��O%�c	e�ih�ص�[6��KK�Ƌ��C�xvO��a>%�G	��0�,kŲS��Ēxj������Z�-0��J��m-?#�u?%\���ZZG�~g��-�#��g�~^'���?$~c��&Vͥ��Ţ�b�KKy���kcM��:^5xrO�<)o��I�o	���t�*qz.'��=~�<f�������&��=�����������|�f����m̥��nV��l�F�ּ�tt���.0��Ѱܭ��*압]'N�;e��j{����Xi���p�..V1Aw����<�~>/#���w~�/{�Y�T��ת�]��o�߽��/��:�\��#�/�"ӕ�ܝ/QP���I�o��I/2�����_��"��'�u��x_x�n��[:=�l)�9;�K�Y���??-U�W�����f���w��UmU���������o��UmU��ݿ�����o��UmU��ݿ���:î�ӭ:�k[k[μ��<�>>!��e����$�Ou�̄0��j�J�6-)�pl�L;��P��8":r%\��k==��c��ُ�8
 Q�'�X{�).��	���lq�6� C'|FC�$$8X�~h|t�c^��f]8@��7��'0S�rd��m��X浹��K)ݮI�Ʋtra��	c���D�s�w��Pr:�ݍ�
J dQ�����|�zI0|���Е��Z8˧`��h��ы�,�仍���:����s2�9�;ωRU9{xX@����#���wt�\YGN`���G嶵�מyǝ:�8�<����9���Rے\�5h���	������ɦ_��r�ƈC)n�aXJ��HYw�I$�0a�ƽNM-�ԓ�i�f�{4!�2fS4�8��>�4?��K����C��L�lw��P�Nt<��t��70ۆ�Ə��$�#&��CĄ!M����z6�w��!��LpSԁ�m?¥��Y�<d�e����~���.�O��}U\r�����L��ɮ��_0~��8A���`� Bę��	m����#��7<��|e��2f��)��O��[kZ�y�yӮ��7[ex𳂤v�)ů6�]C�h��n�!�'_S�f�n�[\d�ڬl�/l�d}◉�:8�W"�U%�UK)]�C�w�m���������s�I*8��Ex���w��t�t�7�0���4$+�
g�s�\��Ù�Y<l��q2��_y~3�=������$�5����5V��{�>oo=��s����w母����u�OrY9�sђ�O+�u���y�c1g��$lk�l0B�3�q�����9�Ӄ�4?'Ñ4B���7D杸)������1�DLm���'Gn���oL"HW3�:a�z>n�n�ӀY��ҵZ8�͝���j�D�G��HI&�>[�� `����K`�]E�������*h9�P�]�>r�����B�ٔO���/$?����w	 K��7��܌������5�hQA��=z���e=tSЧ���0ѦYa�Z~e��m������q�N��-�50�RI����U�j**+BA�VH� �8�$�sRn�0t�����h�j�_�)�Уd=�&�"��2�B��×��п��[� l����&��8V�8lv����*��x{���GQ�2r��:<�����1��F��"�aex����:T�!$�o0��/F�C����獝�ό���I�?l)�!��0��J�:~c��3���ΖQ�F���m��ŭo-o8�]G��s�^]����**+BC[��nY�1$g:krՂ륝L2��0i˷������F���aD:�2�8'҂��i(2C·X0;㳵ڰ�����ɐ��n����#QcI6��1^�W��QZ0�zDB;f�HSLY�g������:�� xl�'��j)�-�&B�eqe:��ɦ��B{�OL}Z?��-�8p�麔q�ݦ���w�[���c��ܮ�h����gu �(�ˌw<I������Q��y�V�o�qk[�[�<��Q��9�,�7b��m�\$%9�}�TTV���i��@���Յ���?V�$4l��`lp,��O��E$�EK7&BFp�]p���=�k����Ż�LL=7R�\�6!�1�;r;tl����ي2EvU�>�8@�:~��ӹ���wu
��9���(i�ـ�XB84LI���A�y�`���
<5�Uܖ�%�
�HC�Ӊ��+�؄V�h��,:���Z�8���ַ����]Gϛ|��:b�I8jY���#�Cyx��&q+�M'7�b�Ǝ>@J5""�H���1̴Ʋ� �/h���	<���r��w�l����{��爛�c�G��_�aF�^���8^�%��u�G���WN��G�m�������Jo��p�}-���.zoK;�mߠɣ�I!�l���fp��;��#?ACN�m���IR����)Ɖ<9Ln5�kt!҆���4���3���>2�Cg�A�,I�L=�Y���5[�h|1��X,!�0��;kAd>�8�7���VGkN�1��0�jI[ �����������|"��k���rT�j��ޙ�34�N��!��!��rl4yξ�So�$�ف���N��N<����ַ���񡦐��v��ۢB�(k��W,���m�,.f�����А����.i�73���ҥ��#���z0��|q"~��[���)FZ6���n�L���<�3ٓE�L!��8lӒ��Gx��g����AS��l0g�ϰ�i���_M�\��Z&�7�T_�B������w�w}�/I:C�T��H|��%(��ٛ�
���q��L��Yd0�6��<ӯϟ�~qk[�Z�?��4G�>�wz��o�e����^����**+BC����U�0�5\��1�h��3�-2�g�H��%�2;���t��wI�I�����x���6i����Q�,���e�F�!�[�(�l�ZA�U�{;��
e�Npã��d0C	�NM9!y)���=�{�O��m�Cmz>xp`@�:���F~�xʪ&yÑ��K6��l�~�eQU\zm��?9p!���c��������[d��<��i�4����8�Z��ַ8�6����U1��Y��&��Hi�D����!�������~5�6�r���	��v|g��a�?���&1D�9������c�3�w��ϑ�W�Ź=��9b��ݓz:4":�rZ��*9^�1=W�l�>�jq	^y��V�rL��ٴq��s-��9ĭ
�7\[�՟���Ѕ�d:��v67�6ѐ�y���]�m2�m��(ӈ~��b��7{�+��<��Jh�`��$��D��!�>!���q�~'����u�%�KKay�žb���^d���i-x��a}����>FS���O���	�I�I�=i�&��4����L-"�m��Zq-[Vè��-�+�an<ͦQi�ԫO-�%��ż�S��Y-lZf�[�,�Z�Zu8��-a�����i�ZZU��R���ml���il>KMƄLO���_�����<xN��O%�cb-�KKԘ���䙴�<ţ�b�a�1-�����ӂY�x��4�1!�|>$����]q�u'�'j���^Z|��BөiV��\O$q�%�����'��Ҽz��0x�O���^4W��x����⟏�O�}�+R[Gɔ�U�Id]I�J�/
O4𷢓��q����TOQ����Y|��������i�M��5���IZ�ݧC�{�q��qX�J)ؚiϷ�x���\'/�~�T=��w�ߑ-"��VK=��/'.+���sG�BЮY�~xp��_l=��=�>��M���a�K��s�Z��45)����ߺC��ϻr]�˻�o�m��5�{���Tb�l9�w�ފ�G�gx{~�G¨&�b�F�]E��.}�K�]�{����3�<O9��j��X�>g�4sF�DRd 疟/gM�ܣ�w��?���Ҿ���J7޳d�7!��f��{�X):���Mr�ﹴ�'�y��}7�a�m���s�����׿f��g����m9�㝨�٥�e��ίٞ+��	k_Dy	W��n�Z�X�v�+��UJ�PQ�H�ubi<�KkZ�G�%UuZ��㎩_n�4mier�+cIđJ�e��B���*��Q%i��65Y�F�kSa���(�Q�&:�]n���n����Ӈ+�^�S9˝���|U��׎/[Uz��������������U꭪�w���n������U꭪�w���www���W���������@�Hif��N��n-ŭo-kqÎ#o>�<��T,"��V(�1��K-�m �b�B��ibĉz�D��Z�Kk�(���*i��v�5̐��֭�:�d���" �lQ�C�$�x��IlV��CLU��9aG%�UWb"*��(���,b �;SQ"B%mD�1VB��S�(�[�
��5q�d�����QE�&A�I�j`��cQX�Dd*q���э�
R�mF%b��"B�!:4Q�,�8&1ZD*���ІZK��W)k	����5I���G�d�jԄܢ ��<�-4�)�B�$"�RH��Z�+��H����7Z�WTh��455��ێ	���ɍl�,VTƊ�V�2����i-�$�b�X�Hl��$�oKn�]��D�i;m�bh���Q�����*cfD���V�I�E�m4��FT��l�qD,N5����M���rA�Ȣ��Wy����x1��ײ��~[`��wu����޳ܕ����<����)����{7�Ɯ�k��Dkg9�A�g�?s�Γ��az���ro�������f������o����M�)���֎����܉~3�Ag�2�����O�(�T���I���C$rBg������r��X��Cw;�A�_�~��P�F�>�|T(�*�Ύ����V��$[ߞ0�sV�4�<�;��ȗ!p?CU���$U]�ºe!�<V�AgwQ�2�A�������1&n�E�GG�����d�J<lxSg��@�
�2`���� Q�q��y��_<��Z�Z��!�����]���/kRc^���b�\QͼEEEhHYP�oz����h,�9u	�&�v$����~JG�i�1$+d�3���3��#���v�=Yq�}�DN����'j#KI��G�jM7R�T���2��?�=b �c�E'^��6I�nջ�g��̕/�~1�fq_T0�����=�M��u�3YV@���d琅a�ܐ���j_��[�Wu�ɇȶ�i�u��qk[�Z�p�����}�#_}$�٦�|[W�Cw��m�������ǘ�LDQI&Tg%��ܟ��I��c�Q�:�u��>:�LӀ�_�t�*8{	��ͅ���C+I��}���,7i��K��3j#�_�n�N�3�2���a���z:g��C��O�m�n��r�p6A��\]��m<4V�����Ԥ�l�,���d��%Dv�N�3�C���@$��y����A�*t���e>ui�ik|��Z��ַ!���=)���\�r�TTV���(�����l��4H����p�0��li{G�����m�3��XpF�Jg�!q�cMX��]���$y�}d����Ñ�v9x(xC���=����zO���
!���[0??<Ƈ�,�T�+b~<�ӆ�,��*�o�Z/$��]���T��y80�φݼc�W��0!&�=�����$р�AY�l��q�23��֭veM�i�i��m�����?8���gN�N���xy��;"j��Һ}]ӌ�歳�&is�9ɛ�)4o7��l�7��	"U����P%�伉-�`�K8��!��{Q�e��O��x���ח���+~��:��w���;g,���ϸ^0�{�E
��|};Q�V�f���9�t���t����a�߻��G2�{�9�ǯD�,x��m�=������l�<HW��\�_z/�'�߫�]����iq��IEf|�~ P������v��Ð��Yx��9O��u���_I�_�y�@�z�a�I�۾4m��N���o����jz],�#��{����3W5|}����@x
��h�u��~�m�l�0Eb�8��2��>qH�#�s'�lӸ�4��̉�vI�JpN���L����X�A�µ�O����%��/QM%F�wH�Z49r`󋄑XWʾ>"|�4������~qk[�Z�p�����n�g9�o�z���iR:�H�zEEEhHl�(J�Z�a�p��;����u��'������ΑTQ�R��:O8l�SА<�yՇü��d3���i�]d>���n�@������b?�����6��^J���!�L٬kYxp��a�N
�A�v������ɢ���
���&�6b���p!�X�\�eS�[�6|�>|��N�����ַ������:|o�S___a�d��w�\T�~�**+BC��F�+	�A��V��>섛08V�	���f���C��B�͓ۄ�l���S\�˥�):S��XQo�×����|��[�-�TN�tX��]�4:p87��uv9�#����/#�M(��������>!�������+g6Ig���2���
�p�8S% ��EW�V���1�1*�5���-�dt�h��_<ӏ��m�ŭo-o8����I�9�!\h(�K^��6���
L�ܚ�:-($�m��^tY������/�S�Q���'�S�k<��,�%��R"������ٓ'��#!�D!�"�=�4p��~;�{���������6j�oOD�Au�Ą����J����t7�h�92�~u�f�y�쇜ɰ0�f3�1���g�\�Ǘ�*�돜��r�����`���̾u���q�������F�y��b��xļ�V��(�^%*��|Dcb8^B�Q�E����UMJ7�G�G!��\�ѥ�q��<N���kclm��N���ydr��a����-/�=�-�{q�=|{F	����x��Y���� ��Q��gL����7�CO���z4$"ce�N_/)�>��Y���8|lE�e�_G��=��/u��_+����x�4|W����R�Y]�Q�v�uΙ{:V��tw.�����R�
n<g㇅�4G����O�\��4�rO~Q�Z����x�Ee1$��{=Ђ(�CNOB�6�{C���C^��h*�Ҩ'�vؘ�-�^���4��Op!��e����C'3���փ$<7��ӓN��p!Dw��h�O?��� ��ߜl��e�SQ8�{+ݑ�B�Kl��Ӆɞ�(B��8C�Ã���|�<���2f*�ۊ�h��e��~y��Z�Z�q��5�m�H����*�f�TDu���BJ"q�Z7��}ꊊ�А�e�¹t�!��ۃ�����/�_d�?��Z7w_�v���U�>��\�!c�RގP��d0����GՌ�j�I���_/��>Cч*uJYH� �����[\��:��/<|Q�d�B7����v�vpbdO<����V�$4B9��o�ǃƌ�n8`�æ�?��?�`~�"&�pA�b"xD�:&	���e�� �x�8s�%��,D��<&	�h�&��h&��h�"h�a����$N���'H"pN�����,�:"X�ĳ� �%"X���&D�"X��4O"i�ŉΒ���X�#'�&�C���"X�MƇ�8"&�"~4��~Z-kiky������ն�o�ag�x��Ǐ�Y�l�����Ŀ�}����������g[�q2n���|�L����h��:K�	���;y�Ħ���y�}S]ܿ=G9�>�w�g���y�d�z=˯g�}W&gYCU�F_$_RG��*4l�����o�/洒>݇�{�vs�g<�x����y�}�{Φ�fx���-}���'vv�ޝ�I�ن�9���;�g�W{/s�wk�U�{�w�w����޿�5�J��[Un��w�n�����Ԫ���ww�M�������U�Un���黻����R��W��ֵ�]��GQ�u�δ�qn8����qa����"I=���0А�z�U�J�~��Mgb����&3�s���+�?�����>!ڇ^�t���M$8���r�|
c��ŗ8i�G��L��"����������`x��t>0C�C�Y��8ܙ3�d��;C��pf�$pF�Fp�l�s��ǏN�l�x�2�:Ce����ꬍ]ٓo]���mӷR,���3YV���������,#�?2��~~~qm�����qa�ّ�W1��Nk9�9C���&�H�����clmА���dR@1��0�-��2B�e:x<�����k��^܆Ho���A��DCZ?�^��W )R����Օi���B�#��I	����æC��d,lv=E���htp}�F/�ܩ\+�] �䄔f��e4��ic�M��KM�
!9��z2	�Tp7�lk
}���0��#��:]�x!��E:����ې��GMlуg���n-kyky�Gm�K�3�ӤK������ȩb-CYrl�$��x��j���NKc|\�5k8[GnF��NR��Q�&�R$Q�1�=8���Аֳ�xp�ߓ[����J5��j'�HC�`����ٳ�~�{�l�֓�2��a;�yw�`����,��0o�x��.�1+���|�~���Y������S����k��3���pM���c9���u9ƙ*Q�06���	����>�A�2c������u���~�9Q�ׇ��rP|B���9���o~�eG���\��7�.ۺ�W�y���\g̸��#�kw��ضe�8퓙�9+N�R�ΐ��s2���s��R!��i!�]�_�Hq&Dەt:8O��c�eUg�����BI���at�mXJ���؏��|��iŭ���Z����8�0ۛnZ�-�0%0�1(� �;ߑQQZ(��'M������fP9�!�h�tɨ�2���J��9������ڭ�YD.��H���[���>���t>�ia��5V���H��#��CƦn��$����k�����-���ayi�!��K.I.u�c�ǯ冞������q�U�퐈J��BT��F�C ;�����#�&���N�ym*맛E���.�ӯ?8�ۋZ�Z�q��L�N{5�b5>QcE���!��G,"��HF�S{��͢���&sww��F��
�q��d�z���^<:Ӝ�h6��A�0{c���Uy��Xt�t8���<�,?s�ce����ϝ)l��m�ϱo�?g��LGPC?�>8%7o
���j�M�J[ve)u���PST����C�J�C���,J�[*�ѐ����p�!�>���m�YI�Mꌼ>���u�/ʹ�����qk[�[�8p����Ϭ���*R�I	Qo�q�0���XO�!�LGc�զ���<t5	q$G��J�~��4�՗^�i\Ě��M����Z0�%����q��x�p����z]7vg�}�S(\Fpa����ӕu��"w}ݷ��q�;ξ2�����
o̱����7�a�di�߇��s��t��,�a�]��ע�<�VϚV�0��̵�f`l������p�Gś2ێ�������󮸎0�?{w����)F�����I�I�-6�j+���6A��4�Aw�r����~/�H�g�N�`�`V1J[]Vc3/7��x���Л3|�>�ܼ��-Ԏ�b��ާ�>C�mKDçN��/�46w�������Y!���ϫ�>��ҡ��2�\G"J6�i}�y���>o������Ĺ]�ؾ���1�F�⸋Y
�����`rm˿�1���d�A�=��4j�f2�\�!cN���e:|<�<P���0�4�0-�'ђ�*�:>�w��٩���0�	M>&�(�e2p9��2lx�r�<���N$�:4�U6Q�hˠ��{�wbv�\p�p�t��*��ƛ:P��Ĭ|,
N�V畚���m��OߒYm"�u�-�ۋyŸ�����u�q���w&"MV� ��S�,���cm(�@lm���0!�9���J�<�m��0	�LCC�4�|u�$!��dg�4d>��ɑ�i�A�k����A� [c|:U�!�')����O�&S<c
{�ɷ�߲/ơ�J�@��4�F&�����(~��&<��~aO�����ܻ(ýIA�)�$'�E92��~ l����`4�}=wW��M�/zH�����fHh�'Ş,���q�ŭռ��뮣�6ƾ�^n�z�bH,ո7������#��6|{���R�WWs��b��g��.����4g'Bp9x|`�N�y��t�������4I��Z>>���3�(�Hۖs�s�Q������2f��n�c.��A$�k2XD����ɀӡˣ!hx�>PH�Q9U�fܻ> ���׉�(��Q		*�!40�����9�L,��~e�N��8q�i���l���~qkuo-o:���x�/���S�{uC��Y��6X,ͶآqŚs�����П{-DEb��rM��;D�[r���CZ��2�v��ft ���yPY���3+�[���;�Gm����8t���M�>�`�L��)�c�� k2�2��6m������<<�۠��0��3�Ć����i���$�I_d(����G��kg�)���%Ym�/ Y�8��ɡ���W�U�����}im���2��<"pDDM
D�"X��4DD��:'N	�!b �tJ(A,N	b'DO	�0LLMD�	�h��i�a҄H"%����ab	��,L4�b"Y����%���'!:""i�a�H"%���DD���ı8'�(�L� �AD��	�0DL4:pDˮ��μ�-�Z��ֶ��<��-|M��XYe�Yg�>Y�am�f��}�5��u�{����Kg5���^t��4�5�9���9+klO�5���m�󖜴�^�߽~߯&؇%Ik���t�3��|-�\w�|�޻9o�S�׾~��S^��>�nVI[mӻ*�՟+z����X[G���D90���:�Z�����y��s���������.�"�ޛ#6_
{��EÃzA�;l/��}�Ϝ��;;�ʕy~ẽ�}��3�.�<\�J]9�}i�8ڽ8�����-��n�B�p���D'm��m���<so��6�϶|3x\L��É���о��wo=��C�UO/���z�����N��uM��^���K;*m#ܑٚl�-�6�}=���T���N�'���O��NY�z_[︗;������RU#������+e� �c�E���&�9Tb�+*��ȓIvH�LiM�Hk{\\��UA��j9ZȾf��q��;HJ�R%+��WRR�I1HJ����Q�ʘ�n)���&q�w�s���6�y�C��~��{1iU_+�V�����������UqiU���񻻻��EU\ZUn���n������UW�[����ua�Yu�\un-ŭźx�����g/ƞc��cd�d��n[(�����!V�RV(ҥM%M"U���o�mؚ�J��LbHNF4�nL�6W7��,]��`�!"��]��BD�)�.6�"��n�",�,h���%iB:��j!�*�1�D)	B�e:�Q�D8<d�B��![�X��F:	�$�%"��Ց!R�C��)Ud,�i"������en�PEDZ+wR��1��m�L$��,rV�2	RX���B��!TB��"W&V8+����B��Ek��1�R�+�M�F쵻d�D�E"q	�]U6�A�D��4�i:�QLmF���X�MĞ[jr��I$�Z�^�j!�D����X�[v"Z�*C�Z�[���-�JYiHYf+��v¤6��8%����1���Z�,�)0��**+Bp,��]�X)�F����ש��M�w����/���&7�h��}(U��9���|y2�M�%������}���+/����FQ�o�~��پ��l#�r�8I%Xɞɞ���_�
��ֲ����l(�ђ��p)��&�Û�h��X����x�G���vw���5t�wo9w�9��		�)�	���L�,�6�饴��'gfi����I��dv�)�`���{s�+�JMt��װp�IR�[)��F��1	�R���M�ua�������h<thx^�!F�����5��:m�y��e�]qo�?/�[�yky�]Gm3�^}�|���Ϊ�G�z>���Z8�;�u��QZT���˕�����&��	���·���؄+�QR�κvl�A�P\� �<�,{��0�(�3�Dj@��ԟB��A����I]�$�0=�ȝ{��%�͘o��� %�~�G$3�.\�o��L�3�\ܓ!��#c,4J�_I#$���&�faф�#԰�'�Wo8�0�XWK��J��k6C�~8ˬ���q�n�ż��㮣�6s�|�aR?}�TTV��9%,Ucv������l���t�p�ҳ^n����3�[�_Cq!z��$�����{����1t�Sǧ���קꑵ�������#y\������ n|hx�φ!r��[���)۰�@pɇ�g�fKL8y���fԘ		㺆l���Ěz'�0���M�49��Q���2�-�康��󎺎0�2O��,k~�ǯa�y�MBZ���G�H���	�+�����f}:j���l!gh�&�h�2�� ��:�{%�Z5a
�G���^��tYei���.��b*^|����C�����A���Y
�h�7v��++�l65\�>}������I������U����}��qfKfF��6�!��n�h�6���w�B3��=!�O�T��S^+A��l�����a�f���ia�Y~eǝy�庵���󎺎��=���￱�}��Ӆ��WKDi��7iw��u��1��Ehb"ꭶ(��7��-�ȄBV�,���lV;"uOn|��?��QQZ����9��mk_������r>(��?i�ĺ=�=��:��_�Sb����<*N����|a�䮙�(o3��wp';��u#�áxJDw�ym�>_OQxChO:�%>�/g�9�6QG/����[��4q�P��x��4;����$��t���7xn�UK9���`��9�*'��t�ķoL��=�C��똗:t�a�D����A��ɠ�6dx4tl�^:�� �S��M.�p�i�u��nͲX�L����F���.?���6�ke�]yո�������|t���Q�X�DĆ�Q�2�Ҋ��ЖU���~��N�6=�!��������0��A�nxl��	�W��#��ށ���{a��!�A��,7	CK��.��3f�0��&2x��r�3�:x>�!����6��~46}��A�>o?�O$8�(~�$�iy8Ap�$�jݛ�܆�(̙��r�����w*�0I��I������8;$:EJ� �uM�4j�h�����l��^q�n�n<��㮣�6޹O}>2�Z������{gQQQZ��5#yZ?NI#)9CI�f����&��h�cS�3������Ǚ�+����㰆��㿲M>zg<��:4- �"���V[m�Dd���a���Qf�.�t��2�&���#0x�~�UF0u�e�������J�O���c��O��z�*I�3�̇���'�����Uw��O	&��}�?Od��A��Z���_��4�?0�l�ˋu�ŭխ�V��u�u��&~�f$��y�����%��,=�6{�/
2x0֎�q���Y=E,�N�z�8`|{ߤ{)�˺���[{�Yx0\��gXhe�=r|S�m�z0,�A�K��0{��M.�:,x�ll�8��U�2�&�Nt�ĎJQb����Ki���?B������2f3
3V�(��<�4o�>i����c�e_��Gq�\e��V���Z�uky�Ǆxg�����ǵ=�ާ�h����=��=��<\9:z�ܞ��;�<�Ӹ��Ve�Ǒ؂7S����"���'|��{]�Lk��2|Gѻ��}o�J�����o-���L��N��:�}�k��Gǩxp�͟tCx��dY�f>������k��2x�s=��Y޾~��>vy�W};\d]�s�|p�o:x��9e,�<jx����(0liϻ�)�Udl08ܙ��ae:��5��Y3&C����J%VƋ���2tn�vJ���\>���;�p>l�A��c��Y��M��cu�I�j�Ngw>H^Ԙz���:?��7��K�UE��G�y�<����l��@��!Dq�J��Hs��
�<ï2�.�ո��V��Z�p����r�eR��ܿF e0�4ks}�QQZ
�a�tv��[䞯�M�]�J�������zj�*�m��٧.��"O�Um�^q��ΔDHI!����8[��2h�p�����.7�8p�p�א��d����5�,���h��ߏ�-�.�7Z�@C=��M02l�F�Oh�-dt@�*"8��I&��&J:�$�d�;���Ww�ۢǆ�>ᐛw�:l���,�tK?A,DDM
D�"X��4DDâtN�(A �xA�'�C�'DL̘&	�h�&��h�4MƘ&(D�"X���&J����DҎ���<%�bX�pND�"X��4I�
D�"X��4Md��,�'P��	�2|�!�A(D�<'��:C�%�i�&��~-h����m�n���8���>el���mYe�,�E��u���g�?M�����N��ms-���ˆ��s=����-����Q���]�:a;<���Q>r�����穾/��p�ݮ�p9^��s�W���'���w+�/�r��^��z�Ӧw�#��pu'd�}��䯭��t�λ�=};���kG�u���<�F�s���g7_݄b�{$���ym����D�Y�É=�YP�(�3�Yۿd�|���~��𪫋J��ݿ�����ߑUU�*�wv�7www~EUWX������www~EUWX���kZ�����u:˭:�qkuk:|x�Ӈ��>�e��~ޑQQ\'߹�Q)cB�m�U.p����h�t;q�NO���Ð��6;c_�rS��tl˓g�$�AAӃÁ�K!^��dho�>����+A�bs�x��N��4��wm6~�h��X��$���H��s����ɱ�Ē����9��`��_�,Y�sET���0^�`��~]��5�IMK܁N��3\$�����˵�����&ٗj�#��O�q��y������[�:�:���n1,<��5 ��x#GP�b2J�E$	�Hg{��������8S���:���Lw(xo��|�|��4��7�����
=զ�Y�c�]���4BB�ͺl8;lˠƃgL�Udv:0k�rp(J0�,��{	$�'G����6d��e?�͆�O�EH�.���|A��D��c���4`hzx��G���a���ѧ��Ӧ���8�2�N��~[�[�uo8��<>�|lJ���5d.�Lx����v'4�ƨ�"Ǥco��OjQ�E[�!
�)b�JQ�PϷ�TTV��ϡ�}���z�������]%�w���^z���/��e�;��r��>�7X���t��:VM&v���kS��1l����'9�����ݽ'9�y�2/jZ�G�N.y��֝>|�!�g�ɠ4<xP|�;�|�O��_����d��$������Tze;��s>�g��4�>���t�5���ٛU�ey�����q��\-XM0���ta��P$�aC�9	53����~D����W�
��,�����b�Z�89���ƻ_W��iroo�帬U���v�[��¯��q���#�-8��~~[�?-լOƟ��M!�a<ti��W$�J�����6K�B�M\h������=;+w,i�'��'�`xp�O�d.�¦��p�ª�U��}xɎ��÷�·��B[���I!'�!�!Ɗs���@���̖��L�e��i&���HF���f��!)8~��l������8|X`�D���\�æ��l(v嚆�獵����x��ȹ��ȯUau��ac��.���ͼ�����󎺎����32a%e&[NkH�������l�*d34�ʵ�ʶ�\�0�v�$I6Rrv��D���tI GZ>�U��=0t,|���M�U݇}�T�_;��B7Qf��X8JL�MI%Sp�|X�8�џ�r1���95�H��C�ݽ�o=*l�t^��|���A�_�_��H8㓠���&x�Td��y���ݎCF�d���[O-m������󎺎�Ǐ�����%�*Ɏ�EEEh����V��x���a��ÃM���ɐ�q��0�ؼU�WY���ۖY��R%\5�����x����t�W�WMVώ>�Zt�Ȅ�׾W7舓�1A�N�N܅�㏝�v��[��Plo5(�⑨��%�ˆ��?5���?�Rx>�333�x~a�����$$'����Ð���׳��
(���>e��~m�庵��󎺎�^���s#V�b��2L�$��FU*�ޮE�E�2�SǙU��ml\�CX�8� "�z��(D�li�+j,J�J�$�\���#��_�QQZ&���ʜ��O�|�܌�F��NpL;�g;�osfI2!t�I��Q��<N���'Dy,�~�m�y�[���-;���gϿ]溏�>�����x�����%�.�w����co=%��)���,�aO��s�>��x�8i�	>�C �A��V�U�Y
�/s����,i8���P�Ic��A�t��ϲ'�CC����f1�>�9c���òdې�r�p�j%+�*x���i�����>�9�Řl�GH�}WR�S��Ly�qc��/4��6������[��xJ�*�D}l%�R�u�j��*�84<��`r�����v��#P�y$-�xv�Q d����!�11�n���A���N��f2��ca|�O�mŌ���y�w�ݔT�Z�0@Ğ,�F�4���%x�nb����l���Y�2A���a;{|H�$4z����!cF3Ã[t0���:ˍ-���������[Ξ<#�评\�^�F�d�	#x���������l��i"���ƴ�hّ�����h���8:�#׃��u��CsfF�v�ц�
��@�t��s��L�2a���%�R�9	����l0��:9����P}τ�C?s�V|c:kl�V?���#&�I6=���}$d�=���$!���vYr���?6?(�\j�߾
v�p�2�C̢��[-����ykukyn:p�����2[��6k<�v��nk��**+F��vN�HsD��?`4t)5�;��z9á��Tܺ�1LLQ$��D"���	E��w�`��a�`,y��[4?'�)�I�w_i;��f�+]̞�%a����a�d9F�hi=����D.�H�TRA�зdaa�w�d������x��ÚI:3����D���|t91���m����67ß�ZD���Ő��	D(D興�x�H"%���&���:'D�B�AJ0�8pD�8"tD�`�Y�h�`��h�&	��D�	�J�K
��p���:"`�:DN	�,K�,�B�DG�"xD(O �D�<"h�'��A,���Q:YL� �$0(0�K0�4H&�!B"t�D]y�<������kqn���6���>e��Z,��,�.�#���7:)y#e��J�,>�w����;>��do��9�]w��l�)�Y{�tpҿ�=Zs���}|Ҧ�������q�y�m�;�}��s��V>ٓ���͝�����v�����N��4���ʹ8vR{�r���W�}�_z{��h�U��:K%��r�������6-��I�g=̺l�eg�*/����Wy;s�Q9�{�v��:ʪ��ϡ�W�2]nΎ��ZvsO����i�s;E�}���Φ�8j��n!�,\:�%��}�������_0��������p^I��;�w?n�=�k��n�֠��}��7.�М��t�]sH�W�>�3�����M�n�f�tӞem|�n�י�sf����\����7��<�D�]��z%Uq�TU�%P��J:����Z�\����N$�m̮�)vi$ګKݷ�4L����HѕX�MQ���Z%�r�u��bnc�7��(FӍ�pEci��=y�;��{w���T]C{��?��������*���V����7www��ª���wwo훻�����UUQU����������𪪨������M!��4ᥝum�kukym��uq��Ŵ���;��� �J�C�N��H��'B�P�Gq��"4:�E���CD�ʘ�v��Rțx�D��"E�ѹ�IiE��D�J��4B
�,D�h�-��Y2R\�_��Ś�BZB��P�#$"C���)
<TN��pB��("��P�I��K^H5!$��ˑ��:�&GF��d��%d�kSm�,�+j�,�6V�[kb �" ��	�$���+��!D�

XP�X�!1Q�f �!J�!1R��(�*��� �L� �QL�dQ�6+Hc+ˈN¦Qь�o!��.&��A�E!F�ē�#��`�F��c*x��:�r(:4�EnF5c�Ƥ%N$ڰhKv9�%
'crGciƝU���*L�Yh�"u�2U"�&�-�,N�v�J��8+[Q��ac�Gj-Ɔ�j���
��Zr4TJ�*�WJ�V��h�I�J�X��QQZ=�{7���O㷻/�O�[��Q\�����|���p�ϸW7��h��<��ǜ>)zKy�s7�|{�,�M�=�tA��.��ĥ|�+�u�����;-�g�R��󛗼�)o�Õ߭��X�i�\7����:OM/zq��z?����zC��pi'!�집��*�����>vd=����H|4=���x~���-тN�<O<<������ht?�|߉�Xᥲ�G����˘��v<�F!�CC��>83�k�aUGG�o�Ph>sð����������*�����Y�mJ��u�6�~��=���<��DV_a_V�2��2�+i��Z�����[�:�:�,;���Q���S(�����`�;F�7�F0���*�&���:Ñۗ���;z.n$	#��G�c^��!.�l6�q�$����\�ׂ��a$2�#&Ɔ�f|N�# �`�ƙe��j R�6��"E�H'$�\}u&&�7�	�$$��?||rn��g�BJ�]������χL��秕�|�=�xy]>eq�̼ӏ�m�kukym��uq�^I[���(��m�"���!!!,<e��T!Up�h�d��í���B}ɪ�?[���}P�K��j���%B.~3����MȾK+%A�2y�e�N�w߉'vBN���'%�zUl8��XGl���3��a�f��A�Gh���I��xY�J�enEgi3r�:n։8�l��,�f�-o6�������󎺎��J��ܱ���je��̥�,_�gs�/�й�9������R�h��"t݉�6�E��!�@m�;^6��	!r�߂�Z���7A����O7�2TÏ���^s�6O�9��EC�Y�?�,i�����*Ux�{Vk��#���~߽^�c�ԭ���ǭg�P&N���(��S�F�>4���ai&x¹�~��e�e�]eƜym�kukym��uq�{�w8[]cR�å�iW4��E�W�5�9��@�b'x��С�u�ݢ�ݪ�gP�7Zθ��D%yf��CE�F,�ք9�z���ߊ{=��㿱�C���O�-��s:�.���}�7��6^������8y��t���|s_?r�QY���Ns�7�]ü���,҈rp���2��f���4o��>����-�w��#E�^zm>�i���X���o;x�M�y���e6p���1�8x<�:䤩8>��.�C���NXd0��t�Y����a���9\��t_~I11����f��!!!4�ZG����h��p��>��UNHh�ao��3�0�����ա;\��ϟ�yf뿇����i�r�{�.uu�w�4���}7�K��c�<~(048��h�6ˬ�ӏ�Ϳ-n�o-��㮣�Hi�}�v7���T�˩.!��!!"D��g���e����#�	:>�8����	�N���`p��y�ē�N����ev�cA�˶'F�ڪ�O���C.M�al���A�|S�OD�;U��]���_��\�N<�SJ��7�	+�>�34Ő ��J�24�}����ҕ\0i�[���㐏a�9�l�BBH����|��[�mo-խ�[�:�:�-���3�̹����>���f�ă���j�sTJB�e��N�dm�
�A�z�m6����g'����}�)�S����*�]8������I�'�����y�Xa��f넩:'�=2?^<v�a���T�#!������f�t�y�]�ֲ<{I:�M��c��dpL1����b���R�|��.<4����g#�!�[iտ6������-�uq�����h���lx���:686�#n��!	����^�o�2�X�Y:VKSLi�Q,|y�8��o98��ä�+�QM׽].�$���G+u��2����PX4��8.��[IU�C��č<4tz������"rp��!�a�dIN��I�)�mG!��C�-����ѷ��G[e�\i�^mo-խ�Y��Ǆx��V�j��)�9��|p鼜=h�ͧZ���Ts�!�:r���T1�!����&�V' �%o)GDk��!*R,��۫g�B�R/������$���uin��_5���T'�26�Q��ϵ)3/7�}��uG�ә�b�G��<Q�4a;��	��/�x�W���L�sh���ɷ^�x[[���f��N��Z��Vv]�H�/�R߉ �m�n�}bPˇ�Պ���3�UT+�����~j�<fwv�����|8fx=�{?�����!a�ޜ�L�h�������l�@`25f�]�6B��h8;p�0nF�)�S�-�ˋJ����Ɉ�u��٢�m�����A�p ��$2���ۓ��"�e�.4�����<���V|t��:B��|(�5R�nuՉ�K�H�%!�E����|�����S%�x·�]������>r��͜|�ܸi��I/f~��q�4���C
a���>r�w����%���Q
�Fkh�W��C�4�c���1�0<yd�<������F�����B�s4��4��<�ӮrT��ϞCF6�ݭ�i�_4��?~Dy��"h�G�DJ�&�"h�tN�Ӆ � ��D0��8Ȗ'N��̉�0MD�4MD�4D�!�	�J�KD�"p���h�"&tL:'D����"A�"&�G�A�7�"nȚ&	�:%�g8�BP�A:FN�AH`Px��D�MA<��^yכa��<�ֵ�������y��>y�,<x���qe���g��,��S�v6/�;m��_�\Nqn���~���?r�o�H?;���G*�_�޷{�{IZ[k齟��)�0��;����S�l��M`��L�����p������-^Ϻi��� �>��m�x�:w�;ť�Ϝe��}���$��y|���3���P����������K��{�ۻF��r��<^.4s�������Y�Unwނ�H�|��K_Ю��&�c_-6��{����g6�}5�Fv�;���y�o���"�3��rz�w�S���u���Uu[��n�����߿EU]EV���۵�������UWQU����۵�������UWQU����ƚCM8i�K4�����-尷�u�u�_s�"J4Ve}>-�lJ�'���P�{�/��كΕ(<'5-���O��!�ɴh ��G���mt�(��Y���̢�t��4�ڊ��Ng���.�������>P>z`���W��Ր��OC����_����=eT
�u���\�]��H�1^�1�����q�uo6��y張�󎺎����N^Y�`�B�q$��ݒI A�d�'��u�+�!��y��#��r���x����u�<!��R��66B$2?�������T��@ΉC�̛xp6�6<<S�П>���6F������7\;�o�D�~/�5��=^!I��cci��͆Tlq��R�ę�xc��0|�Z����M#��m�yo6��y張�ӎ�#�H/S��R�v��k�� Qa[��x�s��9/!*���#�h��(��^h-���JT&�Ă��jG6GIr�U��X���2L�)��o�I$���m�^ԗ>��n���4��[c�Yi߹�
��
s�ӵ�>����<u��Vs�:\ӾШY//wz򞧻4�W��/nʝ{�WN�I�%����Y�4����]�+�r�$ڰ�ņ�;�����˙elyf��I�^����X�Ow��z8ϡ�3C�?Oy22
'?��M_9d����p;5� �2pvtc��hR<�#4&i�vMW
�HV��|�W�|�rfWL��?�7�8C������)�CO���^-�N�����덆�٢̖p��_�[�<��Z�i�]G\e�F�,H
,ϒ�-%t�b��T�ӕ$�@��gc���0ֈ�Bq���}R�=x`փ����B\2�1$���~i�N�I��̆s!�Qt�d��8�BG����71�3�Bi��a�n�u<�-�l�9��p���Y#vH��`œA�^z:ɠ��#:l�:~6On�%@�+�����0�WV֯��[#h�L��m8��kyǞ[�[�8�<t�-9=h���:�I$~��n�,bL3���yʏZВ��z�2�S4r�붛ht<l�^�j��26�~Ç�j��t� ����!�8�/��3������]Owf[�Ι�����$&d��}����v�L���hpx��h�D�6߃�ƈ� �OO]7iwH����G��Z+g��
�U�Q�����uo6��<����<xG���8� (��O�X�o\�I�6�)هL]��t��.ƍq}�BG�~Q��0k#�ǕS8~ק�Hc����B3�v�.�!�����U;{ϙ�
Ld���T��*�C�z'C%��>,$'�G�ωU�>>&%T��_Zmِ���L����c$�I��%M�U��h;ͮʔ"v�MC�P�9!��ZG�[+iǖ��q�����<tGN����'	��X��!(�|��qD�r�܃�9H��xE��7sc@�g4Z�U�%CP�UZ�6o�$�H�����M���nϋq��i���n�@��仈ե�!���qw���9}�[��	��gs��ܙ��֘>�z���I�7N�9�9���s�{�������s����-���Y��N?Nf�N��5>*H4���Ơ�	%��%=Tl���4Y��pv��6�(��������)�U#�����6ezCE�O�a�RC	��;ӳ��`�lK*�p��A`1�=ԣ@�$ِ��Q�};�oL'�O�(x6{A!Y�&�~·#M��y����ߞq�yn��]ӄ�&�jL�:$CjI$�?6큇�v��ɰ�BB위Mt�V���7��6˻�4{����f<ݙ
��vೣ�ݦ�u�0�[��d�懇�殊�X��uJ�,�H�d!-�Q��=�C�=5�0�;~6^�P��$�>8>��z>z[gφ\�>dD�>4Z.I	��e��-��O:�ߞq�yn�g�����?,ɯ�5��"ǈ�K�4��*�Q! ��ir�ԒI��/��F�mu���30´ꏤ�g�g�60lá�93�]���Q4a�m.�:,���_,[��>����OR]m�p����o�p���%/-��k�],�K6sox]U�%J��
z?�ϷR���'�Fߟ�i��s���l<s<n��K)%�jW�a��p�N��vG����������+i�V��{�yז��u�q�G�>�b�����c�RI$#��L�x�c��|WK(�h�+�}�Vv��q��0G�=�:n3&�����g=���
3�|����K���G������ \��2��k��nJ2�w�Z��f^{c��b0���]�M�'��=�rJ����ɂ�N�ڛ˙�6�=�_.SJY_%UJUlm�q?�����sէ�?/O�vNSMQQ@P`C!���ش��m�E4E �L�y��t�؈�����"$DMD���M4������D�i4H�I&��M�D�Җ�$��ih�Ih��i��KI�K"h-$���i4��������n���KI,�K"d�i���M,�E1h�&���Zi�%��&�K%�HI-"m4��$�%��,��I%��3���Y$�mi$$�ZD�I��I$�%�I��m4�4�K$�H��]q���i%��I��mi$��I�I�M�$�D��BD�I���d��H�H�I6�D�"[H�H�H�BBI	$$I�HM���HHKi4��$$��&�BD��Npq	$$HH�$�h��L�H��BB�P�$$�K%��H�M��ZI4���bmd�Ii$�4Zb��"H���%�i$�m!,�M��I-,I���I6���%���I��M�4�i4M-��,���I���I��ZY&�Z-�����D��Zm%��-$��mi%��4�M,�M��K$��4���<��,���$ZZD�E��K"h�mbZZ"Y&�M���$��H�M�-"$����kZjkC���&�Ц-4�M-6�i��&��&�ii&�M4M4�M����i��֚i��MM4M-��M4�4�&�h�&���M��4�D���ZD�Ţ�Z-1i���LZi��KKKI��4�Z"Z-M�MDI6�"&�%��DM4�q���FѬ�ё��LF��#L�m�#Y��h�4km�X#Lѣh�mFq��6ѣh�m24�F�dkam���ӛ�n�I���a̍�f���F�h�4�4f�lh��F����F��kn��Y�5��X��4h�X#}�6p�؍F��CF�5�F�F�F��b5�k4b5�F�F�h�26�F�#X#[4h��25�t�8ka٣F#h���h�hѬ��ƍ6h�5�#i��F�F���4klѣmF�m6ѵ��M�4b4ƍ1�F�dh�k6F�Ѵřf���[�M� ж���M�	���Ё�M�-� [;Yɨi��6��B̄��Y��!16M�[i�ɦ&�k	�&����bl��̚bkm��&�i�ɡ����&�i��&�s8��D�MZn8�d&�Bi���i�kMm4�e�I��M4�4�I�4�$֚&�i4&�Bi4�,M&�h�i��hM&��M4Mi��i��I�6D�M&�Zi4���iué�I��&�h�i��M&�MM4M4�hM	��&ɦ���Md�4&�Bi6M4Ml�M	�4Mbi4&Ț4�4&�Bi4�hMd&�BhM&��4&�M6[M4��Y4&���&�Л!4�DКɬ�DКd�I�4M	��M&�l�֚&��M&�i4�Yc���,��Y4�Y4�I��M4m4kLZkF��i�5����h�h�De�4Y"D"�h����DD�E��$Z-4H�,�B�H�M"�4YE�4H�Y�Y"E�Ț$5�ZH�mD�D�D�E�����yp�hH�---FYE�4YE�4YFH�Z(��h�DH�E�"К",��D�E�б4H�,�h��hkDD�E�"DдdD��Z5hM�(Z4Кé��hM�&�ѴК"Bhi�M	�D��DBh�B��F�Bh�hM	��4Z&����dMhi�4&��M4&�hZ6�kF�n�puhZ4дmh֍h� �4B���h�!h��ֈ��h��ж�h�Zh�"��#kB#Z""6�h�k7!��l�DF�jѢ-�CZ-У-�BЈZmiii4Qh"-�� �D֖��"��i�i�4M��"&x �n�����5�b��@ҚhN��W��`֍��S`�I6�OK|]C5�?�_�5������6�R{�����O�VK����������0 *�߷��?�p38?��֝G�������'��[�/ſ��{|�6o9?������s��;o����x��i��?h��O����>������L�M�����V���6��8��~����o���������w7�so)_a���������'�e�ߓ�?w�(����?����ڦ��lw{�l龞�����l���&-��I�������I���E���ݭs����+�����$�?>�'C�v�yҨ}W��~7����ן	��_��-�8� ��҃��c1����SfocM�r�[Q�[�cy��:Zf��@C��k����v�쁶<g��|M�ޏ�����P�6͔6vl�F�5	3$6�P@T������'� T?�b��N?<7�� ���� �q��pR{���J��D����?�$� �?��/����������n>N��}c��������+�?�����?��G������S "~�	��0?�$��H}���?:������?�������m����5����տ_��g��i޻zt?���~C��UP���(6���~�!m�������E������M�����9O���_��l�b6`O�_�P�
:r��$�=�0���%-�DTB� 1-?�G��?�Ж0:q(�����Ji���b��P�<����q0[�����~y�>��?�;A (��w~���>����Ҁ����ʟ��g�&����=b�?��C�?����~?_��2鿳��u�3|�����ߌ��6�����~c|�m�;��oᾦ���=��ݷ������7�7>��c�u�}�}�jը�Z�jը��(����
+�իQZ�j�
�EQ�ejQX��L�+)YYF��L�Յ5b����QJڊmEb�AF�PV+�b�X�V�b�X�V+�V+��b�X�V+���X�V+��b�X�R�X�V+��b�[S)MJ5mL���Q�(ԥ
V��J�VQYE2��)B�)L����څ+)�QL��E2��eaJ�+jVQ[R��2���)B�����[R���emJ���J�VjQ�(VVVVVVSR������+++eee++j�Օ�YYYYEeemMB���հ�YYJڅmYZ����e5ej�Պڲ���MJՕ�)�+VըVj�Z�mB�e+QZ�mZ�
�����Z�2��V�[VV�+(V��(VՔ++++VV���YYYZ����ej��Օ���++VV��YZ��ejڲ�յe�VQZ�mZ��[V��VVV���Y[Q[V��VVV��Vիj�+V��)�SV��mZ���2�b�++�YMZ��S+VԣV)���V+��b�F��V+��m��e1X�ի��b�[(��V)�SVV++�e�V+56ղ�����¶��V���j�J���eb��J+Q[V+j�E6�B�b���[+e2�+Sel�YX������Յb�Ej�B��VP��S)A[P���jիV�Z�V��++)[VQF���V�EjՔڅj�)��V�Ԣ�ڊ52�(���mZ��J�AMX���P����j55mM��
�b��V(++5m[V+�
�b�V(Պ
�l�V+��eb�����b�E
�b�X�V+��X�V+j�b�X�VS+R�5mMYMZ��Z��j(V�5
�R���)����jյ(�EemEmZ������)���)�j(ԭB�Z�+(V���թ�j+SP��QB�P��������Ejje(�El�55b�YYYYYYYYZ�����[VVՕ�e5
ڲ��b���յjjڲ������B��څejښ�������QE5��V�VVj�Q�e
(P���l�B�
²��5
�P�L�SV�52�mML���+)�mZ�ڙX�)������V�b�AX�Vjj�b����+��b��X�P��X��V+�Պ�+��b�[Vղ��V+�ڊ�b�X�VՕ��b�X�V+��R�+m[S(�����j�+)�Z�e+Q[R��e(R�e
S(������YEmJe�+(QY��e�VԬ���ej�J�e++j�VR����)B�)YYJ��5�����eeee+j����j�Ք+++++++)B����eeee
�Օ��ڔթ��J+R���ڕ���55jjjR�X��L�5++R�Ԧ�MYZ���5b���|?G�|�����y����lw�=����g��g�}��<��g���ȻI9A�E0�ݪx��0Qw�"�0���7_����_����V��9�)�|������L�
�O�ҿ��fII@~������Rڸ�������?���^������#_��̅i����Y�ڧ��_��?���1��́��3��G)�>6
��OІ�������=jm��g�w�d����|��t����ѭ����_���"�(H9$� 