BZh91AY&SY��i�B߀`q���'� ����bL��           <�  
     �P  (  �   
  P@   �@  t Z	S@aja����$�R���$
l��jRU5�((�*���Ԩ��	�P��h P�%$*"	E[4F��4m���UJ��eD��i��b)IP,

%J`��RR�(i�D*�� �
�TE�T*T����%I�*�c�8��
��!]��@ rkٖ�8r֎�vj�����2�*�k2��ֻ�����n���Ji�F�l�M	U�%�ƦNF�5��\5���l�� KA����� 8��!�'_7��ۂJ�.zn�iJ�R����IR�g���Z�)%/x=��n�%;�o\x*����^�R�$JG΄�c-NwR�)UM��$���lւ�RB>=)J �Gw��ԪQR��=�)B(<�x�RT�T������f�H�i�ＥC�T��:UJR��N��T����ϯ�H������ןR�*J�>7�}�%R�.��JyV�5���T>z(�� �8�t��%W�*����{�J�IHx>���U)J8��^��T�>������U^�=��ġR����zP�S����J�
B�>��ET�Pxy";i�J��U)UYi$��R� ׭=��DT�yO��T�j��G��I%JC�,�U ��h�)�/M�O{�R��I�:�J��\�ה%J�\S���ے�UR�+^�UU
���(Z���J 1��(����p��L���P*RR�J��	����&t�ROf����J�+m*�^碔EI]껪�AI���М�r��`mTJH}J�{Ŗ�  wtp �&/� j��g5�Sn�p6��t{�@
.R�z=�T
�:8 ���= *��J�S�Y�*$���T�<�̨P�;���84�Q��H.�\ت;�� k��}x�*������h[k:�Z5R"��HP�ւ}�H��3���	�N Q]]]���{�E�Xi@��:v�8AGu�tn�� �� �Q��T���a�jJ��ԥ( π�6ҷlu��:��(ۚ��])�����놅 ���t*V�Wu@��P*��p�(<|  $*�
 S eJ�  �    '�F*JR� !�фɀM2b E?%)U=F� ��  � j���%��bb  �   ��%!4�  �     $�f��M1&��jzj4hML��~߿���I5��W�4��ގG�m��"�����uktW���r�7������w��W��
�
��Έ *Ј���p����� 
������������������ҧ��@X�RI$�� �*����PE�����_�`��'�~�`�m%�t��%�m�lKb[��Ħ�-�l`��6���`��6��%�-�lKb[�[غ`�ؖŶ�-�Ŷ�t���m�lbFŶl[b���4��4ŶlKb���l[b�-�[�4�6��LKb[���%�-�����Ķ%�-�lKb[M��Ķ%�-�lb[ؖ�`F%�-�lK`��6���`�ؖĶ�-�lKa[����m�lKb[��b[L`��6Ķ%�-�l�b[ؖĶ�-�lKe�#�Ŷlض��&�l`�ؖı�lKb[M�4Ķ�-�l`��6�I6���-�lKb[��Ķ%�-�l[`���bF�-�lK`��6�-���Kb[�6Ķ%�-�lK`�M%�-���-�l[`��i-�lM0m�l`�ؖƘ��:b[ضĶ-�#-�[��-�lb[`F[�����-�lb[ؖ���Ķ�-�lm�l`�b[al`�l`[�Ķ�-�l�Ilb[�Ķ�-�lK`�-�`�ؖ��%�-�lK`[�LclM0-��-�lb[����lK`[�����%�-��-���[b[ ���銍�A�"6�R���؈逍�A�6�Fب�Kblt�V� �� �
�A�6� � ����(�`�lm���T�
6�R1`l-���� 6�Fت� [`l@m����+*[`#lm���6�Rآ��` [`#lU-���A�(��F�*[`#lT-�`�lm����"6���K`�lQ#�6�F� �`�lm���6�Zb��*�b#lTm����(6�F�(S؀�0�6�F�
[blU-��R�+�[b�l@m��A�(6�؀�`�LV� ��@�� �F�*� �*�)�lK` i�lm�l b�lB1���Q-�-�U� �)�lm���� ���؈�X��*����-��� -�-�Kb
�[b�[[b�lQm�1m����[b [� � [b�lE�"�[`� �� -�lm�l�F�
�Fؠ� �
�E�*�`[
b�؅�`�-�L�-�4Ŷ%�m�[���m�lKb��6Ķ6�0�b� �lإ��!l`i�l`[�č����%�-�lb[���:e�)�lb[ؖ���-��m�2���ؖ�ؖ��%�-�lb[M�-��%�-�lKb[��L-�L`�����m���Jb[�Ķ%�-�lb[0��m�[ؖŶ%�m��l[`��6Ķ�-���[b�ؖĶ�-�l�$b[ؖ���-�lm��K`[�6Ķ�m�[c6���m�l[b�L-�Lb��6Ŷ-�-���Ŧ:clZb��%��[b[ؖŶ%�m����6�N��*;��L.���o����t�?��E͏D�k�ܡ�f撷�s{ބ�%��\]�w4��x���Z[z�Za�8qV���k�����A�oƛ�9���e�!�3�s~\]��Dp�M7i:�bs�{
�ں�h��%���V/aK�\�u��m�Bi@F�nl�.�a��Z/Jkw5�0ng9�F�齯�3�hOoC���6�瘝�?�����g�x/9;N�U,d��ZU�5ئ��H��q:J�j��q�su^i{^�%�W"�T�ۃ�3&�͂<h�������8��
5��t�]�n�d��8d�J��;�]����ٳr�ww D�4fn)�!�ˀ!�=�_i���d�Y�;nP�+��%�'�ۗ�S��29hK� ]�׫���/Il)p�^Y_��e�ݮ�9��Ps�`�F��cỏ7D�fs����^��T��ƒ���@Nۈ��\�s��V��j�]I�;�9���"p��N����h�8q�N��-�Mގ]��M�g%��P�7VdOxN��;(W9�}����ٍ�rq�{y�v4���Θ�S'd)��e��l��؀\��Zg!�wFh��n�i6q��]º��*}�\�$�n�+೪r�d��5Q�8�an&�k7�w�v�,�Y�	�кT�3���H�ǆ)�0����[��͵���u>��.���ˠ3=G��{X�i.YÓH�#��^-�^�֊�'��W\I�]���� ���m�kɑ��x�!G����7n�x;������w0�,�$kn�:����d&����ߗC�gf�pG>�jUgJv���C9��8�.؞���7�i�`-�P��pk������4l]�L>ՠ`Z�-�Cy��KCLCt_��ķ$��Ќ��霩&����������G�� 3���,�8,\&���e�S��[���_bn���Z��q<l����i2~��dJ�o��q`q�C�|_�w\��sGh윌�"�&��<В�i�1����̺q����b��O~N��F��7���68xs���f�i�r�o@���.�!:32d�+y�tN7#=�õܠ�T��X�ޭh�Z�v�b�t�k�J�%�����fW$�s�z��\>D�%高rh�E�h�6��޶�׍^Cv ����s�1l(r���{ij1ڥc.>
Y���ڇAJ�ǻ���%�/ja��lB��B�=�vND��A8��۽rf���`��p��:c�>���rN�Uʦ�c9*xoU!��M��jͼ8��7�*���Ѭb�Wyr��{[7�h�$�vf��v\-���;%VC&�����>ȳ���v���bl��sp����2@D����L�3f���=e��
��
��6��%a���!�;{{r�眲p�yG3,o��`�	x#���m ��b���6S7+V)�He��5��i�\���]�i����y���.Vu<;V ���D��!����S(%�{���6[ת��MM�Y�<�3�1:cDt(��{2��z��:���_&F��Rˢviy�_W��涇Nܻ�nN�FoӉ�5�j\\����.���bu׏�/o@�$���6�D<HC�.v\a/�	�.�7E���q;תŭG��Np]u�Y1�c����k�>l-^͇\�{@8��>�W�fvŨX���i���A��܄Iwy)��"��ڦM�\t�S�v�n�:�^z��u�syOdJM��L��+[-���w��<Ǹk�+p�����ŭ��FM�v3Xc\p��@L\�";cG 
#�bΚ{�r= G��'P�$��}�۹���9���6���szvNԋ$I�t΃9�����yf^S�݆�vL�U��kn��� ��&۳;��v��"��#��׸oBx�L,�/�z�2���c����^I��gj6hi��L�5����h}���ّqנ`vn�f�)�m�Wv�U�溋j��;s[�y�[Z��{��]���J{iu�{W`[v���!Z,jA�I �u1�3p�p�˽4#{�����3G<�4<ٍ&������i�h�:p��*=�w����E�8��	N@Vu�
=t�+��Wk��P�Khgq�4L�W]"f(Tȥ���0���\���E.y\��ɻ�
��<�bk&���'2Z�[�чB������)A��R"�Zkie�[�hǫ�+�Oj6/ ol�.ü��ah�F7�%k��+�4���\Ù��9"ئ��Y�V�ѩi��Y�:]�*��mᔇ�2{V�!}�Z|K�f<,�wr蛹�j�{�ᛛzᔥǞ-�%ѷ-$ފc|�s���R���m��7EL��2o��l�6��3r���Ud޹ܔ�ro|�׼7nۀ��0A�ͦ��IV"�`�M�[�������s,Mo��A���5n�P7���)�ˋ�ެ��&l��|��Cjb��\rf�M�KJ{o!�)�#��=ǁ|y����ո�<�Τ*G.�1	 �s�^�~����]v�U���qFt�x�^.v�o�q��/�^�}LJ��@�|�Xp��;.�VgH�����uq��sڤ��J�]ءX��*�B��%2�LL��ƉoA�5�oE
2	܈�ۛ�7�Zb�}a�Ce�՚V59�'ˁ�q�#Z�Y��t^�S�J�r�p������	Ǥ{�3nN�[���r�wR��_'a�B
3�FS��zom�ɗ��=�S����ǋ�����Έ.��@6ڙ�K:���9Dn�4R��X�F��ׇm����o�a}�ۇ�Ou*f
��g�n���GU���$t.N�h��QĞ��o"s/m�,���Y�n�"&�}R��a�yv���Ie�X�nb\q���O24���a}��ǳ�kg��h��ŗ��8�n���@����4.�&n�N��u��.�,�g�s\ȫ�t���ݛ�m3��&']��������t��.߱���#��v�ךy�Wk�a���w��­77�4���k�(�ܻ�ǀ�����6����Йy`�/�T��拆L��Da)탦�]�@������`�3qh��q^ߥg��m�rp��1�*N��Ōwq�@���#��x���z�G����C=�v�_h���mq��Ӛ/�Vڷ�/�8�&������}���ӂT�<1�׸'n�i��{�.�un۱�9��d��]���\f�,�7EW�ˇ�����8��=J7M��qs��}�v�et�l���(6ńe˜/Y	i\����v��[<����\�[�`�o�{��@���6>7��4nnWB�Kc�:��pm�yݪ�ϻc5.���ex-�ހ-W�-t�&ś��2<�II�@�ۅ�&ج��Һ�`ܖӻ���h���!�Ps�����YK�.�r�u���zJ�]@J>&�R��xn	�9	o̞�y�lU�#]%���;����U���f�,�zu;�cۏx77F��F?�r*l�o]�"�L�����-!����L"ʎ�;�����Ï �(�9�;̌��K�q�C�X���2�
L1N%��GV���E�+�8=1��&�'�/I��ld �ƫ���*l��c��lЋF�ؙxo(�pC˴���X�u�fvw`޻w1���ͺ���Ê���?.:�V��΂�g���8���<���&��H՝~[�h��s�
}�\��$�؎�q'�vp0�`T8��8���KR��Ɛ����_d<{�k���CFj���C�;&�]�]�GbBҔ�\7��xŰ������&,R����k d��� �`{���r�Ȕ� ���}*0G����9�Ǔ�`䵚�9�x>�RwHzk�IW����Hub�	x��@t�03�&�Qu������2گJ6-Q�v.��e)���A��l/�" ^}�l�4��x�lU�熎�{�g@�6wyn�Scwz��'U�\�JB���[���#-�Cb���鶗E$aKw,0Ly��<(e��������I���al��%Ͷ����;��]u�����V#d�l���z����0����=f? ����z� �r���X��w��q`��a3N<K�� ����()�� <�(���Z�������S 2;�8�gU�w{����]{G%8½�+:.+�#��-v,��\m�>	Ԉ��Հ�cO
���< (V��Ӈ����NN�bӣsq>ʒ���'pTu�pvqW�(S9,��W�3ڴ� �tS�.�������\�n.��cV����M}'���y��涣%+�8{9"�M�����I�A�L`�8��I~z�DKضda��'��3Z��m��h4�qr��4���"7�w�	��:�Y1��P�`7��C�c��.��ģ�zgd@`�D���{ غ�ƛ��؇K��n!�����Q�q�D.�A�y�\wG.�O�	�"���ڱ���*w,En��i�IG�G"x`Ѽ�T�Q�ڡ���� ��99}��i�-y�rB�)ww�V����-��8�Q9�&ݎ�C�oj�	�si�@�l�Ŝ8�r�Gd�gr��������,��u2
�#ۆa8k={���;.[���9xK�6;z& ��p�����'Mɱ:�Ȏ��۪$���f2S���z�Yf����wQ`%���%[�f�:�����ї$)����4��+w8�hd��� 3���زi�.�M��\�(�3�ҷ�Aȳ��vI�Wڴ,�����N=���ۤ!�q�ܯ;�7퓫�<��S��.B�R�±���,�*ǻ�W���y�$�ck5Nƻ/1M�̦� �v`�,���h��P�`l�[�I��,֊��駚��1��C��2Y��M �3�\���(�E�<��sD:^�aO]��\[Nn�8]��q��NTo�{�����[�Etikǿ<Z+������kUK���Df��@��0v>G��`SJa6����ݨ9{9��؃�����/��T#v9����vj��-3���.y7oN�N����ه��q�LT���2с�
��[�9aZ{�G�vƨ����]ۯq�7�9���zX���ŗzv� =�W���>u�:7���m���S�,:de|����Zy��GGܘ�D�d�g1�X˝��*�W�퉸��v�����wnM�w������V9�-K�Q/p�8�z���!*��osYx&��qc�������hUaI;�h��5��ۨ'��0>�!�,���;�۷u��f�
�FR�qX�"���I�� ^�td3J�C�R2�����m�I�pՄwu�-|�G����븈ޅ�ۥ��}�&�a�U^�����)�@"�1Lo�A�vġ�v�Vo J�b��n��w�Q8#��auYe�Ht�ە��tHGlS��9j��V���4;:�P�N�;r����[����R����K��"�7�]� y�:V6�p��D:s@:��Ç���p��`��:xv;'![��/��g]L&(y��l�K���~�۹��9׳�eӍjY��cҎN�e��;�ܛQ�9�˕@�{�鷜g"<s�����1卐',/Pʞ���rz0�����O��P�42�8��G���+D������<��jb�Rm4t�8��.�ѭT[���K�oy�X��:������������,NP!"�.l�I��&��j�Ш�g���wt9��ph�����8�3I�����oH�%i��ǎq� G�:އ��J!�����$e�{Սfw.K�=�)6��OJg���3I����I����J�<g�x�I���J=J���\/IE����F�"�m��:�B���n:Qt���:^v׾;f��=���h�����z��|1�"�s��^�k�����OF�S=8�-���I�q5x�Y0�#Q���K5L/�������7Ǚ0��{�v�_�׳�E���Wh�
��+N��R���a.�ƞ};K�S:ue��/;��1���Zy�~�NH����_)f��yw�{g�x����5��w�a��>�՞%��l�ԍZ.���RQ�VS�a���M=ƌ(�6�x��ЯzOq���sb�&���'�s���Ǎ�HY��1o�P/�J�#���4� �{f[M��`��v�r�0�!\����k,fw+�z�ku=��"Hsݹ"W��F����a35s�g�WΜ+H\'#x����m�ǧ���	��t�����_�L�sѡ`�_L�9n�Ǹ����=f����^F�]��)\�"�U,b�)�3��{5kS�/��G�pW<N�'��� ���U(�M�q8�'�b|�/��z���|O��
��3��$����_��Q!Rwtvh�d�P���w�x�l�)���V�w�qk���Y�촚����r�L��=+�zvt�ʒ��>��O���x�>���x�ݳe�|hˀ#8�'�IW�Nd�ų�
L%�ͤ�O+ʵ;�z�}�􊧇�s�I^X��݆�ln҈�U�%������[�I�Fq�oۂ켢�8�4�Œ��'���l���/`4̖��>0v��x�3�RQ[/�r�}��W.5&�b��Z��q]�p�Դ+���4ve�Y�yBcVzYlV
ؔ1�faHV��p�Y���ƹ��ۖ�8��]�����0iޑӾ�٨�4`��O�A��D�qK:й�r�&��co]j{'�����;�3p.&HdY�X��Y	������??;|~���_�����I ����~����v�Q��gkot-y���a/��.�zޭ�|Of�|�.�WG1O�`��:TΖ��b127�\y5��v�9��%��;"�!��V�ݐ6����Qx;���VQ���&&�|�5HP��,�ӌֽ�VṚ�n@k��ή瑫���*ʜ'A㸼��6M�R��4���̗�ۄ!������|4�.��}���^����Lse�_q�ш���=��2I�n���N��ŀ}��	㻎A�Yc�}�k�_T=�M�J�=�3�i�3�l�x�7a�Ť�ܧZ�����邿,M�T��ݳ%x��;a�\�9�.I"����2�����u�cfʛ6���8S��	t �s�����Ǵ�42vP�]٥�^��3�'�於�Hg��7��uGh�+�'c�����mm�۽�GV������ӑ���o��ѝ��[=/Vv�j��ÉTs�ۜUtgH�@��7F_'[�������Y/3i��qE�v��X��m��a��C0��iJQ#�{}ްb�n���l9����<(���|�ۇ%���{���S�����t��ٓ����;d�|dΝ�9�ej��X[��њ�t�氧7���.�.���·+���UL��G�=>�	�9=8��I��N�Nyl�C����t]')�J�鳰�io��;wCu�/yhE���i���f�m2��o���	�],�݋KN�-�7�]��*f�y�a~�G���a�[R��vw*v��VM{H��YU�3,������^�E�^oC�������,&z�b}����9�5xv�sd�}��78iд�}�m+{{7z;D 	��x�Y���ڰ��w;�>����Ǣ�BM2�.��Gz��l���0o��)^�.oQԍܮ�~���o.���j
���[P_S4�0�34C?�nca������/p,1��$_X�ņ��Ujq|�C��5�Qe:y�r91����g"��)K�̲)�p�.�2�]�A���e!i���q���e������Х����͜24i�l�+%�[�۝�6;@*G��l@
������Q֯;�ln��y�5j3��ۋ.�K�7ϳ̭q�.sy٨�f/I�\+{(�&�8S�PNW�lPd�����e�6']��_��6��XW�na�)%�SfnYpZ���ѻ�N�YX�%ǥjG��w%[ٶ�7o��g���Ǘ/ne뼡���p6���9�ڨŞ*��]�v/c@Verc	Gί=ɣ�b�V\Oއ���F�O-�����rŞ~���I�"�Ა�P7����;��/q�9�­�f5:u*>(�#��'6u�3�Z��l<U��ӹ�8��͍5�nt��l,RGk^n���$��˽]�3���2�y}m�j �b�97�1��n��;Q{d���ߞC��ݵ�jR�O���#;G{�j��V⸏I(z�t�iPL��Ǘ�h�QƞY�,u�/��@3r�C���M$���T��z0�+훬��gU%�Lc��%Ѽ��m����h^s�������.Q�ɭd����zͮpkSW~y[d�B�H�b�:z
��x�fu����Enn�&����%x�'H��X���:ZX4kn�v�u��)e<F���®N�"Vo��v+d.f\�2	Ք���v��3m�/��I�t�)�{�S�0�WM��m� �����;���Ս�;"�.��;R��5p�5����&�릳,���/	ʙ�w�/�J_��:�{��{'�;��]O\���:.	��� +Ҳ�gK��!�!x3��n��$�h�@Q��7�
諾�I�hV�N�ޏ���"�_�y����:��np٣Ѹ3����)��p�ڕ3�U�\���̩4ٞ�@������j����t�Y��j�������ʚy�	��gT.��֭�3m����,��Ǿe��3X^r���ɷ����t�����ǋB&J5��rJ��u*ҺӓV(�a���<{�O�����w�n�����.�s�P��z�k���,}s��U3d�������2ˍ�d�{��6�՞$����7��{-�������M�$Q�_n	�w*R��}�T�Skf� ���LH���>����g`95��ەr�`s͆�-��l��Yg�	v�b҅���7{'�x�G���e�4��J��� ��4�<|
�{ؕ��QC`��N�1;ۛ`�*�s_�k��ə�:}�v.��;�P��Yh�zww��n�,YL���N�.�)��Pţ����O3��cq�Yβ�S��� $��!^T��L�H���@�[���\��bA<�wF�����x�';d�̹{�K�ܞ�h��&��[}�V���ݷn��w�2�B1�V��*�1�����s���Lv{W�pS�u�a�ѓ���7����*�v��ب������w�ת���ܘsH��E�J��3~H�U��l[�b�tm�'&I�Y�.��$�p]�10V���J��v ��7�eb���b8����Z#�_V��|�RbfP�a�'ͫǸ���#Fm�#\7�4$��g�9�D۷�Z�|�qi��\�&(�;a����������k�U�۵PWLʝ��en��0p{���:�{���l�=���e"��{��N���֕6.��,�;��[wjK�X{D*TR��r�k�o���A�Z��{�����i��}�N�n�v?hK�xzX&L��j��'D��Rdzݥ��R.�T�-\�]���2�q�ج�joS�y���z�N��/$v;�_	�W�wݔWe]O�^ʍi�<N�2}��|�=��H�ί6@��/z�x�ה7�<��vl��d�k1t������q��7ő�w&<׊���<ʃ}��Fr��mv�e,���y��bW.Q���[��wX&Ω.�S���SFY�q&�m�Խ��5r�CO�'+�R�Rw��;2R�&�id8�u�Y�lu[�4��+��F(	Ǌ݆�o)���d� ����k�P��������e��2��:L��������XgU�w;�����ju`�aFZ�,\�u�wN$��ZjL�۽���nm;�PM�.RF�,�"eV�����{�%���KuL�;~{�P=��:p��|�
��	�o{�2���L�yJ�t�VP�u�����PknPx&�wLӂ�iN��+�n����I �%^Lon0!�̜���40h��#�t��/�	�N�(9M��Fd�ն24l��sE�);T�!�$��0��{Z������{%X�-�z�mt�NcW���nm8�F�h=�k3Y̛qQ
�����h�|WQzM�^�68Th�z�F���ܭV�n�sy�n�g���s�6�v�R�%z1'\����`�cђb�0&q�N3,þj���-yO�,��yܺ8�3���f�^�3q�ڷ�༞q���rz���p��s���غnX8�=�p��M���LL�أ��=Ƌ�{>
޴�����NJ�uL�i��<oݝ�&:�wK�ܷ�^Y�hcl�4�u�o*B��
��\��.2���䨝��G/�{e�Q���e��h[�9D;<��\���6+��=*��{��Os���r�"����+U����q���{R�2f�d4k�}�$����qy&�V��Q/���ޣ���h�{����22���w�:�>/�k���_g���>�En�:8g����'��{�w�� ���ޡ��ܙ�uszҼ[%���"Au&I�����C׽ŭ���<se`���%��;�(�<R���T�F0�Y��{Q��M]<�l����tb���7���f�#�S)�c�Q���5-�ݠ!��ѹ[�(�K��Ֆa�]���{Hf/�rҝ�;��x&1|���NRJ�V�k*{���6l�n�e[�˻��W1�;�J����E�̥B���hR����Ⱦz���������]�:A��:?@�,#�Qm�z���\�0=j��p�N����n-¯{L�;�e�ONdۈ�$������_�����G�7����gm����A�{���\�Jљo��X��;N��%+]^�x�fFqH3�n� �v\�d��ܗv��j�ؼu$�{�aeC�vs�Q������#]Ĵ]�|�����1"���d8$\��/�zI�xi5����35��Y]Y��!K7Ga��;��A�C�
��Z���ļ��~ãt�cdQ���g���tk�Y�O�2���:����;d��C��,�K�01}�Y&���1j��s6jr[6�:3�Y���RifY�XөH"$r��9bT#PQ�Z[8��9��VL͙�}�7��γ�q����63fB�{���8��q��1z8�zv��YC�ٛ�齇=�wT��J�>�t��q[�+o���z:�>;��l�6�=���\Ա7�ָ��H��
nh����&�JAs2��vI�]O�� ���޽��{]@pa1�`q�ū�wc��BUӫ _Lv�*�}')�|�ׇf���=��l����Z��}�
l��cO�朤�dY�a�\��$֎Z"֞�ک�vNxsN.�P�����h�3v�ك�I/l��U|��H^�֜�^�6��O^0����+.���V/�p��P��R�����J)��t��\͖��9OG"ei��^k�(v�4aO-��z9wd��p�b��r�ip�l�a�=Z��<"h�;ΰ�V*�������� I:4$�M�ǰ��<vp�V��N��=gSe�B�m_�����#���� �3�`�ffǳ%!W��2��{�V��\�Q�b$���y�A���8����ƅf-}Km�]9,Ҷ���t�T;���5Y�;<H̳��+w��f��6��zqڵ�M�=�.;�7R�`mJ�]�L��R�4��p>�g0�zO���f�@kC����#P竢~){� �8���kfv;س�6����;sv_+� .��V�[��l ���^Q�[X&�DՋ�oS=̱6QƄUq�d��k��=��\r�U�[u���&�z��i�(>�Sf�m�륬��o�+]���˝̪i ���"���+����j@IՎ�"e�>�gvP�hx��٦o�Өey���iJ���vb���۽��,ɚ�����r���d���]�)V佤������,��N�Ӭd����6Wb�i��ޏ�Y}���W5M�A�#Jnݱg ��)r\����L��V���Ơ�4�7�Q��8�C�K{�O_"��T�MR��<y�a� ��ٮҀ�3�H��i��?�g	=3E�������](�<��ɳ3�Z#
�W�M��}���q���o�[,�7��'�O�=��v盤��������z�}���sxx����M֞��8��'��6c�Hezh�ee�ق�*���ҍ�)� ���wk�����P���;�S܅\�뱜Ӝ����݉�fP���3�g�[^e����F����S��nz�S� ���ϕ4�OO}�}�{L|vw���Ʝ-������#Xs�����a:`�{"���3d=��E�_�$�J�5�０�����`ɂ�θ]� uu�bŔT�.�,ҧ�b���˯*۬{ӄ�lbS�٬sPOA4��<���^�����Jo*�U#T)cC:��v�Y-�8C�
��Ig-�r�^��FJo�L����T+��� �m�����)�Ao��pL띏����9���Hf9��>��"�7�&`׼��F[��7k�w����O{m�ý��u2��h:b�XBz١��dg�F��R\��r�]n����C̙�:�͹���CF�������F�m\�˝������}I�9��4����~�����%�CT�rv�]�*�Ckf.�`м+���������&�cc%*�Lr���F���FzXG�s=�
I8G�Y��^-hb� ��38f6s�ϴ�IG��:|�n鞣����}�fg��f}y��3��[2���1 m۰d��&H /*��pC��ϳ�E{����1c�|��u�&��#-�#�?d�l� ���BML�n��(2+���ײUl��&a�>X>�4�q�1�f�x��130��T^��z3t�U�9Q��#�-y�> a8}��Gٗ(��SQ)QlX��~�$3�BG�L'�0��ŏ�� ��d}�pџ8Q�27	��p�~�%��}�г9jx31�v]��MRD����Ġ�����M�X��1��ί_֒1���|k<1���Q�����043��0�' ����n����h�ύ��9�����]R5�i����M�zk�TP�7M�2 ���)!$���\c)�L�8�+�Ĝz34b����}�a�ぐ ��|������U���\#A	��oU��h�uY|��:3? E�{�MPH�$7�<��T]Ө�MS�h�꧇��������,E>��}z	����?����������W�_���������t�J{r�G�6B�9�e�\�d=�c�\��O��zS�Ld�w=&����{kw��n�Ѹ^B�J��Y<}�$�,
滞^�\No.z����.L܀�o���{�qq�Of�p��F��{m�̴�m{����Y�-�Y.v����M�M (����޸�DjL�9klu�κwA�.����Bg �jf��[�]c�\0<�d>/q��7����s����h����
G���O�站{5Z=ճ#ᨼ�$��
���3F����c@��l�Z<��x����n:BƴWîu��ڣ�iA�N�>�B�9�H�*�:p^O��t��e��.=o6|<^*�p��k���Q�r����1f�V]��=�!�eO�ù��v���m��aY��jE�;욾۔����j���[˃���p�H�X��KO.�Κu��פ�]^w������=�ے=���v�+
 �u�1�T��G�H>�h�ac��v��ݗ�8�;o3��b�t���R�œ��t��rۯA�~~��-w��׷��1"�Vejs��
���UT#�gtfZT�2-�Ǉ>�G�RW�֩��Eh�u~�����t���8�8�8ێ8㏎8�q�qǎ8�8�<q�8�8��8��q�q��q�q��q�q�|q�������\q�N8�8��8��q�q�q�q�q��8�8�N>�㎜qێ6�8��8㍸�8��q�q�q�3�謞ٯ&�;�ޒ�9i��;m���0v=��]����ɱ[\qf@;��b�Z"���O|���uᵲ��Z=]�L�{��`���b+N����_�G�,���э��@֕���XjE���L
��E��`�)Y��Ruٸ��B)�����-J�=��5���gfMX{%�U!N�c���Eӏ�}���ĆL~�K�y�J�p9���� �ō�Ĳ<�^=�ﲢ���$��]�_ �c˸�g̉����gl[���Y�R"[ڏnvs%}��+{)fb�qsg�E�^G|ߟ��&��z*.�Df���YǕ�[8Mዖ�4Y]7��) �*�-<Ֆ������L���#�+fCP�E�q�&{Y��%��ӣ���/��2gG�|F}����{�	�3Bt�`��hꍍR[�oaJ���+hР�E�����{�7���7b���x��[��\���'!e��;�
<Ċ�)�J�F����5���K�`����[�cY���>\b�e�Vu���$���V����m�����^�5u�ջ��ͮKk-v-����,���F��X��A�-�;��7<^0�̑��޾������H>��2�\��J�z����ӵ���z{���88�8㏮8�q�N8�8��4�8�;pq�q�q�q�q�n8ӎ8�8�i�q�}}____\q�8�q�q�8�q�q�n8ӎ8�q�}pq�q�v�8�8�;qƜq�q��q�q�======�������9��aN��˛�;�G"^\�N�y�r�Xؾwp��Vb[�,���&/��NY7Å{k妆���;h:t��m�yuD�J�W|�]w0�Tv��\�=�u]Q^a��O���mN�]�-�L�W�G��ޙ�wX��1����F^�ܫ䎒^���;wf�:���C�(��W8b8� oh0i�C7s%d�(��ww\}�0k��ɝ�3C���)�,��Xw۔O�xzk�'�4Z��f=�kcb-ɏב����4�/�	��g.K0��K�Z����h�N��������{�1����Y�ew8�d%�N�W|����:�m�5�W&7�33���h�RT�Hi���΁Z;o|͹l�}j�']��}&��/��V�&����/E;t}H��Ņ�$X0�'sN#��-�ïco*v좫jv�ĭM픁є���yI�6�7Jc�84
�b� �>:b���K�z�ߏ^Ƥ�u�r�;���e�%>��Id���6��+�J�v�v���P��Tv4Ux�����ЕZ��,�野 \�����l)��a�d8u������ȷ �>tzZֳ�Ս ��e���>=���Ü�{a�QO�;2Fp�z��q���6ճxG`�un�9���+|�R�{���y�;}x�c�8�8<qƜq�q��q�q�q�q��i�q�v�q�q�x��8�8�8�8�����O���8��q�8�8�q�q�x�q�q��q�q�q�qۃ�8�8�88�8�;qƜq�q��q�h�ׁ�d�{���3����=��&j]�3bdq,Ӽ��ԍ+-ڲ�������Af���۹��ܚ}������8����VU�ߦԞw1^t:�雍�k}ǒBܻ�h۲ɽ|m����|���d#ϊv	��b��eJ�xW+N�Rz��]�Օ'�]uZ���u]���o��)��b�v�QJ�(�e��9�S���J��6�vX����S�=f��I$��`g]��*1nc[^pO���^{�,q�f�{��3i��^�do��^��]��1q�ub�Cľ�P�h�ͫS��n܌�;(��~�M�'z�$̎��jxB�̰�nYĵq���=O1,R�7��F���Gy��=���Hl��~��E�[ڛ �TP�WF��������R}� �WE+:H�e��=\<w���rK�/��u�m�A%��
b�y�
�h�"�/��u��K;��7z�H�W]ǚ�@�����gގk�g�Y�)�y�� 3�2�f{��&����Z����-L�u\5�v�쉰�����H�}_w��jܼ���ˆ�$��6��:��v2o�39㭻]sb�]5�Ù�һ�t��p�l�:�,}�_G-�nI�?�KǨ�;J�$w��W#�ќ��gەt���7���6��$#����5�9���{o�ݼx��8�q�}pq�q�q�q�q�\t㍸�;m�q��q�N8�8��4�8�;q�q�q۷�����\q�q�8�8��8ӎ8�8���q�qێ4�8�n8�>8�q�q�8�q�q�88�8�;qƜJOp��w5���钬���f�Iګ[�-Y�%����x �r�X���P� �dA�a-7�g5����=��7ޙ�-4x��x�� �����wT��f��̣p�n�g�Ly�}|V�\Yh��kg���O&�=9yl/����Qm*ά$qj34�C���~��n<�C��_H�8P�v�Bñ��x2������.G���c=;6t�n
R�N��M����ι��ұbM��3���8)reE��,����N��p��8RP~I�c��/,o�=X������|�u (fU2�#���	�Y����/��UCn�^��L�3~�5t`�Ҽ�ȗy��j/oh-����Π))���Oܘ�������2�ؖ7��\�U{#ܨ�#�g�Պ��wY���c���۟(J=}_����&���G�0g����*z�����o��o��K3�v�5�lzb���2�M���<Z�g���S�x�glK��
ۡ�v<HGE/5�c���v �Ͼȵ��`5M�}ވ�7�u>�dZ}NzW䟦��`��Y�s,�xL���9��H�z��v�L<�^	B�Ž?(���%�囓���ٷ��Z�\�q�JY�n��a
FF3��R\fww�2��(ތ݇r� k�n����='l>�w��:|��Ad��S�� �h{�͡[�T��/�_a�BОkq�w�Ӝ_mb� Żfs�c''w-��z����7Ddf�r����ձ�J�+��5u��Μ|�;a{0���l��;>�)9�W6r,���{����O8�T0ŧ0�Q����U�oMK��k}����I9}���Pn1�|SG�f�������7���v�sjW�Z��#�e�2��o����;۳Иs��/5��&�I��{^l�����>0�v�mQ���kbś.P�\�z8��V
��i{=KMU^����Y����*�ɹ[\H���!�zfsՏ{_�Þ��}^H�����2b�|Z��=��=�H[��.5�m� �f���w!�q?���71Q:%��4���|r6W�-'�8�y\][y��D��X �ŗ�������R{풻��q>�;4�Cd���(G���wӨD��Ȉ���7{��� ��9��o	�m��j�T�i��N�3�ͭ*J嗘�c���ۡ鸻FK>�
"i����H@|��#�٣O��lc/�NnC*}�v��������f�/��NcB#�ՄpX�J��j�n;��/v_?[��n��Yr���ͩ[�D�e��{Wd�+�6��2
������l����ԝ��B���N^W�]��S�(��H��Q�.1�[P��a=�������d�݆�T�b��0���xx�FL�&�l*jp6��-;����uY����qM�ל��=��w&��f	��M��ڒ����2`k����k^:&nȨ@������$ǢX���G����}s�.೗�U�n	��S@�m��co;�q,Q��Ƿ����Xs��+M�~O.]�V���]��x牓���,�]᥆��4{��
��"�ĩ�ۢ��qi��J7��S��S6��Vͭ�goT/+R"�u�ixv7G5��nN��$V��!��Q�Q^W��x�w-��c�{e�; ����>F���ku�]�ˎ�l���Cx-_��Tk�����vl��ⶒ٘f�7�b]��}�l�8[)���B��˚���kM��-\<�n玛�r��޼T�v���ۉ�m��e�廏vuM&aCK&��+�G?�x����wQ§e��b�	�^X�Üݑvs>�=��ě�r����H^�6�K��\���f�b�f�N�K���KSR M���^�3��r���w\���&�S�)�\�ğ[l�f'��\`L�z�M���6uk�Ҭ���C�oE��=������^�ܻ��*�ϳpc˜j�����8�Qhubj3i��bn�^��7=���ܺ�-\}���\�0�yg��	�m��ʪ������\�c(�<!,�޲kw����R���[u��d��͜��I3��ab�����Hm��.!;�a|.�.����M�e,}6�˛2��-��Uqxs�cJ|�/=�I��w�z}Q7���"���v�A�H�,�/I ڼ^g>lINo<���ˊ8p[.��r�mJ�9� ������ɔ�Hc��|9Aņ6*4lPF�s���3���X2��{g��?g���U���o�fL�g�6oTT�y8����.Yq��f���Jq\�ii���=ׇ�A��y���׈�<]l�X����3�Kh��]�y�9ΰ+v�JL=�kj=t�zͪbۻ�lL�U����	�2P�kn��F�疛��0-���C9^���~�IEv�!0���������u������Ǒ�ޗP�Ew{��{��W�8���eu|��.�׮{�\ؼA6#Q�o���Ӡ�Ob��ge����V�D�A[4����H�����	[�:h�y3{��EH�ɰ˽&=���9�b:u�vo���{r\��ݼJ�;�����4��ܭ�Im����B9�.��o9T�5=�G3�����'2g��I���}5H�m���YkB��DH�pV�i	dzf�����j7��ʹ�pÄa�'��˞�i���/�_����G��V��C;N�f4�0%�z�)�ޗ#W�WIbf�+��yI��v���70z�0]��SD-���n��HӢv[uw���7]'X�h�ym�6Un/���(�.��~��$֋���Ԗ���s+ւ���w��7�2�-6cc�C@̝Vp�xv�l��Y�Y�y9P��Zq�P���mA��ܺ�@�<
*����@��wo7A/�<V)C�()�*cn�V��Z���C��q=g97�n�r9��n�M91r>�Yt�^���w"�p>��M�YN��'�����_�&��S�=��c	��=����_��G:x��7��9�3�X)�=��h��S�C�<�c3&���wn��^�ݹ]]K=2w�̥�
��b�j�����(Į#p�j�G��:V6�WoWu)$4��F��{R����t�'56��6�nv��a��ζo#N�㆕sdܮU��Xs��m�(8�P��sʗ=>ꏮ۷.ݡ�n�V�,VA�Ë1d4�'���yj�fk:\|�9�b�y\Omqg�ja	�l��S��e�k����֓��V875	�DBb��]���q8���/e���UJ۩0��1�����:P��3�v{9�K�t�r��.��c��z!��������٩��"���z�5g%a�p;{�z6�QS�e	ǝG�\ۥ�dX\���J��6v��p���k��N7�BCaՙ۝*\��x�͔��2*�*���	#��U�(94��w��Srj�|m����䷦��\�k3jʓr�q1�&�t9+:�twY(���4��Z7º^��@��6n<Fi��Ԝu<2.�ϥ<W���op3�\~���^Gnʝ^�pi�pZ���>�`jٯq�W�PG�-���_g5��5�y�|�W ޝ�UJ$��;�f��*$d���Bm���+�N6e����K�QҲ���)�p�`ʼ�c���z�>����gzi܋���-Cr��=s����f3x�eZQ�]��۠����7���JVb�{\���I�50C���*�အ���>י�g,u�J�fN�cj�=�759ۘ��/4�;^u�}�8k�`t�x�V��G1q�������`4��Q�@���-����A	�M�sT��Uh������TY�=����jj���1%�3����^�]�W��c����<aH�/<��f�O�lb��V�S=���d�ؾ1����%[���KW���Y{[2s��`4�&�_R��ێ�"�H'%9�r�^W)�I*�,����O�ɀ�r�=湞�y�oZ�-/��/�5�?����
��@�����W����/�C������*>~7Z������^3�7�62Hk�l��-1�6��M�	"P85�(a-�xX�?�cx�ǋ
ÌC��+�`2nA�Ԩ�[h�j��E�
�$8'ěh1�5d��G�l\���$�m"�D��	�!�2!��|~����ДE����1Q!M�E��+��"Ck��K�8���x0i�������HV<�&��,HM��  ?mx�n��$Y5�?$������yIv��ֳ-��"�93�S	i
q���Xw����	WaA_^�B�5P�km{!�Ѿ��Y�������9>���p�÷�Hmr�q
J�
��cc:G!��o�潸���,�\CT� �O�/ uئd�k�LN�r�R��|p����-:V�3��x��r}aP���R�/s6�A�����u�^�9�MW$��o��/�;k��#��-eV m;���CK�IZ�+q�r��mkǥ� �3�������A;:�:��+:P���ّB�e��A]�W4�9�z���Sɚ^b�r[��ur���4J�_uv�v%�-����,f�k:;MZ1^Z�\w-�d�
�8zǕ�ex����'���4�L���g��9����Ec�U�Q|�;�}��~��\=}�|P��#�|b���n��F��t&�м$(�q c�sp1��r�����Y�FK��љ���'�0�S���
�'
���J�a�7����x�70�d�z���,yw�6��촥�"�s)�ʹ�f���u����h��������;�=)�P�5�I7M��&����@�J�s�ouo�yFhm�ncx�`�-4J���-���������a�
l�-��G�@JSp�$$[%�a?�M�"N�&	�`��p�M��8�Xo
 �,���!!@�*h�&�P�-�0a���@���"	L2ж�� � �W|�ف"�q1�aɲ A��Ğ�!�r�lAa8xNp�(K%��ą�W�q��0��)b&���0Z�.AN> JZH�ZA��A�P��I�!��i5�dB�C��0L$12����9�b8ǀ��Ʊ��Ěŀ��)��lcI��^(�Ma �Gƃe�Kl����/	(��&
M�-��څ��R��C����5�:�o O
a��<`�~2��*����G�i5	UU�K�Ou���?����^�o�QI BJ$��Ӧ�;}z�۷n����s~~��KKӤ�:�����^^��v�v.��7n��=tB%�&7:wu�c�q��nݻv���1�$�C��r�Y;�n�.����tRBgwdY#�����$�Q$d]B�4�;q۷nݻv�����rQD(�
j�EB�;�\�6�ys�{��u�=�r��N��\r�Γ��;�W9yoK˻����+����ׯ]�v�۷n�zǣ����s�ƻ�滻\���ޚ������;���v9��p��4�m�ܒw[;u����Wgy�Ͷw�{(�^��X�Dr��㻹��ݫ�o<ֻ��*�o7�K�����F�� +s��h#�]{m����]�M����t��ٱ{���w�{{缽��Ww:m���a/;^{۞���9#������B�����Gnt�����:�����{����ӮN���or�y���ؗ];�˺�\���s�뼟%��׫�x�&���ۮ���d�����J�Q#т�?6~�dH2$�-!i��}|�$�gtt{�����F#B��]�p��/=䯎���<�E��H0�d���:���Γ��{~���u/�dO����t����R^u}7�u?5~��W������l��)��8Bh��pchi��}
Q�""�W����$������x�x�p��{N5֬�g��;��)�<���+Ckd9��%.�9Nͭ�2���l剰�M�[Z��J�CP�'�('�[�iD@a2ᧈcX�g�,#@��~E"�,���b��	C�" �@�͖@߾��J�ȪA�Ƽ	�;�ʹ;�~8x��Y�2�Vf�o�ә����2����<�!Gڅ�L��ye�}Muݡ����]��{Zm�xA��&A��}�[SN��3w���=�� �@�9�@о��K��-���{��R�)�Ƌ�mw޳sW�D��$�����臿t���'j�nh���ܩ��@����$�Fb��h�\fs��O����Kk>�<���\>��R�p왯>��E�|���&�{	��~��i�ֺ�fs�C.�%������f{�x��h�����A�{�k�0�q��� ��F<WsB.���:�"x%֮�ھ�U�s�gտ)s�����؟��Wճ�6��a�H"
�۴���j�"��{v\��S��J��uMi���k��Ō����h\�؏�C��;Y�Vq�J0D[�J��_�T�{X��#q��жɢ�\�qsz�`2��`��#M�'�(���dmL�[��>� ��_Gjf7�^n�S�w�d�F+�nɝ��{D���k�{Ӊ�:��]͸��I�{t�����{􆷭�ת��s�7�"����]�x�-����TY��Eg����wfN��ѱ(m��=9�y�\�U"���tӴ�o	pNWq�}��Sӣt�>�B�����o�q�����(P��s���YG��x���v�h��a�f��?a�/�M�h����ͼ���s�.���z;8�؎37��]s�go��m�A'��6�Z��kg:��=rf�nNf�2ς�7������;��{â��=�H��U_�����ʮ7��2��Gl�jSw���<�;?E�Q��6dݵ{�O�9�7B��DEef�p�k'���k�������U.�VM�N礚�<�cK��O�^w�}��;��j0eJ�6N��-�4w֥]݃*{��q�/�s���7�xּ�:��
l�������6������'2�?b�k{Sc��S��ؒ��Un'C�zy���xi�Ι�]�N��:��3&^!�Zc�.\-!՜ԝ+ڱS����ڊr�W�qbM��6��.ty��}�Ì�u�q�'9�`^���l̐X����T���������^�gq���?^��L�w��;��Y;"����/���[;ڻ�K��E�42D%W�V�VԈ����Emc�A8����ED\|��f��Iy!��k/0�˻e�cG��֎qZ.��ҿ�<��C�����֫�q�����W�7M�6Lϼ�[��y�z���=�_f8�����|>Z���7A��uo��Qd���{��@�ø�Arzx�٦���{��*�e�t
�N!]!���i� �8���u,O*�}�������<��qY�����xyH~���A	O��)�o����շ��ͥ*�E	������^ڮ��3���Meζ<�8�V���5������^]H�c��2�@�L=T����%��1�-0�Όs=뼸�����3���>�%k����l�8L��Ix���&7�z�b2ݕ�s��������R�(��7�ܜ^�U�g{����VG[��T"�u���SU֢�?������Du�2�-�&[���iU��V�7ji��{�NYu���6:K�b���;�o��q���W�&ߤP �Ў���t
7C0p�y6��n����Egl	���&�<2�I\5I]l���S������΅0k���N���&��Qs.���4����ē�.�s=��OP����/�،�I�9�����o��=�4����`�4�%���7R�ܧ��j~[شeJ� Л��͹���jժjH�p�s�)ͼ���g��h�[���J��љ�uek��׬#���ztL�&8=:�٫��ѱ٩�7��Ѧm=p��ʟ��2���T7c�4`��1��f��{���9�~��/o�xJ�B��m�C����cq�ZD�FvC��7�vH3��.w~���duh�>��:�{��y
돐ۉ��v�v��o��Gl{�:�32娎��k�2����rz�!��Wz�͙���kN�!F���2
<˖�\K̔�{y��"r�e1JJJ�����M/l}��#�qSy*e%��T1�˭�ǁҡ]�Oq����s�b�"�z8KX�R�� y�_e���Q�UwTг�fѽnRjd�:D�S+f3]�-�s�g�WWS�%:^���O��Kk�]�95�Һ Wp�/�;�;�^�V<�b�WE���9�s8�y�A��.8Ϧ�v�4�ݣ�O�����C���hK�"�7�H�rk�9��ŵ��M-���ssc��q�'N�5=��Pʑ�p���e�H0��/>���3�)�����!8q��]`�Tˑ�r�����&�'���Z{~��s���I�$@�f�5d�X͐j��M�&6��V	�f͗��=X�N��۳7>&Fp����rx���}�5m>���8w4sG�*K�\�w0�y����ڀ��4T�Z�۪Uv�m񃓼�7-#G,6뎭<g�����}uc�:��7��|ׇ�g�ݔ�z,�O�$Ϸ$c�p���=>���;g�0�0,�N�{���Aƛߊ���u��N�rԯ�/��]h�jS�F�V��4$%��wkJ���C}�oa�`������5ؾ�w���W�@�T��JyҬ�3��rD#�.*�qʆ�uc%%��{{%�v����7�om����m̈�'{qP�ULfr�oc����Z�~��V�����o춂��|X9nP�ڙ!+���u�`7��j!Z����fFoKߔ�>l��*�G�1�Hw�E�GU��@�`�@����`7�]�^w\}:{�+�c���C�3���ܽn5wBX�ts��4��q�]G�g�>������ē|xi�s����#d5@���c
�p�;]Lm?�|glb3�I�]S��f�=3�L��痣���m�`T;J��Ny���W�t{���'r�,b�J��sNnn�%�
@�g�/�q�\��9��u;��ӫϪ����>�(���zƎ�p�����G���g!�x�LUV��q�]Sb�����}��;|�}$�������ݲr�Nf�uY�'u�Dt#Z��MnȮ��:i��9�8�f�-�9�K�������z���YZ���j�b�(OMm�g+�W&	�CB���Po�u`hz�z�/n�Q�x��#$��������p�Oh[��8 �@������Ts�Spn�
��^�ᬶr.��n��z���B8���ˍfM@������ǇL�w�C�c�����g���Nf���������,��V �랈�G��:�O�1�[0�b["�s[i��������0뾆�=C]�N�v��`W/*W@ͲAߤ+���F?Vf��6y��ȸ�����g5�oo�I��{0�ͻ�����}Θ��A؜�/'U�m���x��[��E��W�GLq�c^���D��oz3��molʈ�ݟW�/�Ƴ?[���N.|�wZ��x��}.#M'5��=��oj�M�'��ܰ�5+����f»�ɱZ��M����=6(��3���s�ޔ�h�hol;��4v1���:t�=s��.�.~�k�̙�"��[t��x\��'��2g�,U^Y��/$ߞ�D���}�O��<p-�<�a����qna?0s#��67�Նj��M�:�!��3MJ�*���n'Qb�ֽ�ǯ1�`�ڢ�g1�(v^���b�"�aWu�u���c�e�d<�]��ܺ�rWK��e'ḧmtMMw9d�N��U��7�:��Ϩ\��}��=x��Ù��[�ؙ]qb�_���������d�f���pz�O8��"&3)�}�?r4Ʌ�j��7yAg^�b��,�~lp�9U=�-�G�wX��w��_}�r2}ba��"Y[����Ot9��<��*���;�)�����z%ŧ=�B��MVn~��>_��>�3W��Oc{,�E	p��"GBn��S�*M�Q��ǻ�ft��f� �{rP�=4L��3�=�r�<5�s��%���j��*�hO|�TX���vd�}ӽ��}��T�S]�|,���ˇ��B�u�b�5��bsDVmzsd��-�ћ�/eHzJ��>���B�Pݼ�P��U���=b�?�4ͼ�X�F���q6s!WnK���p��de�h� &:�b��,���v�)��"�yI�i�[.=�y�ч�2�w'+��Y�ozi@�b�ƻ�i�g!/�`=�,걹�&���k9�ݝ[F1{��Z~�י��5���{�Um�#�E�:���l�nN�r�u��Cܬ-��'1�M9qv��2��I^����p�Ouxc��;��;���i94ąuqԐ��Z��
�Eos޼K��FE�g�!dD���oon)��dZ�*�A_C�73Oʫ:�ӯެd]/	\��Y�X�x����ۿ� �w�f�A���>�Ӕ8�Uz���'�M���pi��3/ᓞ/�����nQf��z#<}��G���=��>��9m���N$��kER[���Q�\.��Z��]�����{���w�O�����f{0�������rѦ-�+Z}1Vw��B���I$���7g��;��Y��k��9�}����_�e1�_c���4M̘0Ü���Ξ~3�~���j�Ŋ�;�������r���ۈ�9�8��,�N�����8A;�N�X���ȧm$�N֜�[�>���?D35݆�n�k��(WP��g������$��54gs�d��-&�S�4��S#�����w�gزa�xQ� �a�C�tH�g3u�ev������d�S_�TV��a;������j��r��1I�z��{Sl�!NJw��М���u0eݷ�VdŶ(9z���S[�oor5^Ҩ��1*$��s�N�Ġ~��ۿ��K�]������ܣݳf�6��}��i��7��{6*��&�vF�]�]��m����τk�g�ƚ2x��mt����dy���6�=C�{��ñ0w5��i�����q��b������Z
��P�Z�(�f��9���Aح������ב�Gk�����?/�Á�^��1$����ʖf�@T�tX������Q=z�ofGVn��\;zN�\wN^��@�&� m����23�����C|n�"���=��xؐ]�Ζ&����=���l�n��+=��s�#�?>gnK0s���3�����O����癠�*�8l�� ���[*��.Rr6kb�>�L--�TY���]�S>����^��|��v���̻S�b�96D���1߰e8&�����ZT�}�1��������;�[3%B�c�b����d�v��Ή�5�(�ޚ#{��	9����~3���h
!q��;
���F�����ceo2�]�y�+5�Վ:2#AT;z{�i�����sB�օ����5v�I���S�	l�u��㸃 �1��{;rR���]!�����f�%�:�����fFp�
�R������چ���MeK5��ÛF�J0�
�����z8vUI�C�ٺkr�[{ �5MI����c�+�{�އ��°�Pvܾ�aNa��;������Z�_.�ȻrK��kc��.�O�V�-�5�IȝW�%�vv��O�v�˛�\�C�k"��4��;P���Ԭ�� ���K�Y�:�9���� �q*�!f�AdR0P��^r'Wm��.N�E�gt����Ԛ,o�:�e���BV��m��33��!���<�^+^����|(g=9
�䔠͌uI��j����}�o��U�
��>6d�����X�p<M��<6 I����z�f)6ʤ���H�.u�s�J�����Vy9lH��olg۞7_h�<�'5X,�N���ޱ'�N��ځG��qܫݜL�Qu�	�9;h+9��=m���<�꼗�MXu՘>Ѕ0�&���/��d��Z �R	�٥=u7Ma�>�mc�f�����Z�i���T�*g2�^�����u��p6�%@ɫ�N�p��Gđy��B��bK�3��UϭZ)�)7����Q3�:8�yaڶjـi��U[������P:N�Luv�9�%g�F�ɝ���quAy&7d���W�x�F�Ӏ��½��v���y*HV�Xc}���˛3�9�:�p�����:��}���0��
�ԭ��3���͊��U�t���}M+T.F��F̴�����"��ט�8��Ņ�������U�Ԃ厳l�ܧP��ܮ�܍�bʆ�wg�}2۳��z�]k܎8�P�~�a��,՞�Gxj���:/=8+F{�_�D�ed��*���`�Gg��m�uk������wr�ZmU��ӧY`��P�L�8\��3��9���nF��\{��z���v�� �2�DUމ�X#���H��s݉�G7{�b��g7��������*��z�$O�H!�/)��	r��CH�![��{;�#c�Z#WѴ� q��5�[�j���BjOjܻ�V�VZo[J�Vli���,�g-,�	���ܙ�/)��\�or-�i����39nvzg��;�0B8���D���塶l�2�V���+��c��ub�)��/(3=���y�kn��9�WF�,ȃ9W5���-g��AC<�D �I]\Aݷ2g.ez�2i��USG�	�$�#n=~=~;v�۷o^<z�{��UFHE$�]�K��ѐ��!��1st#��0�7n�z�ݻv�۷n8��{ړ#��'% �]�s��i��˫��YB�^��ߞ��}sQ���v���׏�v�۷�~�����W�]��dC�;s���R��}��G�ؒ@�
�w*H�N޻z�׏<v����w������:WF��q�۩.⸘���#14�/wdwWH�����e����u��W_n� wvBI������wk��r�<���p#�UԻ�t�wn�������r��ɧ9��n^�{����ً�]���빎����\�v:����=�w~=#ݸ�c����K�����Rs�����I'8�9���7+����(Ĺw�u�pr��Q-��� _2(R�C�¼��� �j&�;�{��Pwnܨܧv@��Ȝ������Wun��]��h�2�i�f�Oh�t�T��y�d�t�1�b�u^s0�y���~���@q�[�
٣�f/�:��: ��g�	C��孛pP]�������n(x����i����Kս#���Y��-���#=�{=� \:����xOc�e�Q���F������Íbd	PVe�'�X4�ˏ�������@Z��!�{��`Z��JY�i�fX���G����|�B�ӑ�l�� �a"��7�5��y��Ky5�'E���!59�Z�]?i�Mh�@�'� �g1=Ux�>_�V������f�>Y��}aI�|M�+�Ǹ\a�-sN"0F����>�� 7�=��'u�� *��G�4}c��~�YJΙ-���IG����\X��٥�nQ�@�O8^��/``�Q��1tȾ����e@�T
4���f�ۑ#�.7�s����A�&��3��r��CH
���:�`�^��'z=E�|!1W�"��a�y쾢����i��K���a�=
��!��5�����@�(�sЌ}X��P�KE���Û�H�=��Í��p�qx� ��i�$�ߚx<7�	�����9	i�� F� ��Y�z�r�L��}�Yַ̖��*&4X�!��m��8ޗgyj�Y�S��.�ӵ%N=Z�6%����d�[Q����Y$k���Ә�~�t~�}ׅ�|Q��s~��4ɰ.�e^v��BL)�y׈7St_x./�뜯��
h:n�ܓs��~1�H�#�5���k��2�kۏ�@OÕ���b�[�\�X�M� F��1�-����_:�M�؎��d�������%�g��R�>���Ӯ�f��k�Q�&<��7�^j��`�yaw4bt���x���R+e\i�d���V���]9�)}d4r0(`D��}Y
꥝�N]u����}��'�4�j�G���b+ �@�ğ��A?����t�崸�*����C�g�W���k÷#�x}��0Arb������~�L�W�|</�Э�K���s���!fδ���ua�V�{�?���I��qMi�ƶ�C�/#�w;��7�l�3:�fԿH^��p`���(2���mi圢�� `��?DR�GܨF�p=T.-�Of�)��[11e1;0e{���� ;c[�Ɋ� �Ԍ�3zE�[*�Δ}�OȱC�t���uJ{%M��}�UW\fT��?���eSj~N�v�	�� K�]Ϡ�[�\<Û�(�uQ�i��Z�x������O�m���`1�4��� ��J�+�H�=.��:�f���JkA^�^�f��:��i��^}@<:4aKͯ�[�% s���}�ء�P�ن�r�[cE�`9;��k��"�Ɗ�~�`��Us�q}b)�[�2	�bV�V�|��;7)��e��``*��'}:6�2����kqW{��^J	�a|�`�^���� �o�;��L$�'b7r����J��Q��*�I
v�}'���+�0?<���z<vUxe��/ [��j~lf�M��� Juew����T�>ejf�zz�2�7�c�x��
� ��c���[Ar�L8uW�����eRc���Y.}n��r��T�9���l5w =��^���C�k�R�2#���1��O��������g] �Ȩ%��ך�y�;
������Kkx�^n�[4xn���O�⠔��_���S� <w_/6Of��
�����s�:�W���I��@����P\n�3����@<��B�dI �}�F�wj���!��o�&��:�t�p3͇��k��5��p�ʈ�-2�J�v���/��L�����]���
���9���{a�`~�s8��{*	{`.U�O0���X\l�n5�O])�����G�� #����!������ '���ʾmT�h�ȼ��ui�[�:_]s�!̴�4��;th[3/xq����9H�Q��^�@��}A��
YJ�=��&�=��4�����S�y�ɼ�FɪC��שpއe�q��tM?X���I� �|"p�딵@Y�>�f���Ez�£1�9(vsF8
�]��.Yu֬])0�6
zs�q�=�j�ݖ�Z��]���U�������
��J�s*ݻ䡱�v��#����:�P|�Q��G#���VF.�k��U��n�)]uU~�c�#;}��ɞ�tS�$�|�=����<?� ��A��5⟼ޖz 3:<&P�.d<��v%�o��G�gz �^��zj����7��p%�v8�	e9�u�n��L\<�,�Ρ�I8ZlY��x{ь�A��q E��{���5"��>չ�T�> �����W@w#��Td��W��}�*����څ���L8�r��nO���7��ͽ5��/f�
N�c��ӱlR�{c�]��vmς��[f�5�*(����E��I������5���d! sB��.e)�x땜�+�{��i��������W�8�֑��� J��b_��\���=�5�pmf�f9Pw��s������D�| �"��<��7y�Ş	׵E1�
4�Ac�BUT3���@����]�x��F_L�g`ʝ��sH`9]+͵�K����]0�9P�]7�tE1:�,��{� �&}���O���c&n�l�=�pw�|k�ݞa}>j�=JP��ր��^Z}���=k��"�_U���d�}��	�~"��C���+�X�ǕT�i5 ����00�������ɦ�N�p�j'~�۬4�f_���ḹ�ل�1f6�wstHݵ��/2��bU`]�k8H{��b d?��yt	���w~�غ[X*c�%��,���\�{��{�H��V���.��o2�'�߾�o�f��>0#��G�$��3,�ݠ< F�d<U7�&c�~�y؉��dt F��/b���~l3�<���k��6��	�li�K�A�l+��٪��jb1 �$e���AZ5�<���^1�@t�u���񛗞��[ѽ��ę^ f�xr��|�3�������|rxx��IP;y�J�Om57!��5M��ZS��w���-^�h�ڧ=~���xS�Nz3�Q��#4��#vG�n'w�J�Di��t�<�X��0����i�{� ������.=�l既~���!���[��F��3ݿ=���P��F5�К�9��vԤ=����b�)�g�&�d^��[�{/#�W]Bk6@,$#r��@�q���M �=;�峾���k5Qg�,�TAx�̀��� bs~��.��N2��*' �F?v>֖�㕦��킺�8�� 7U�G�/r@
o"�M���Ǐ@����'o�D���|��9Y���v���&�DfR{\Ď�.��pD����;�
�Iz+�E�з�x/B��,xy���I�\�ǹ��3�*���C��Yri�D;�X��=���X�>,*����Ư�@��߆>�ċ��[G�|�Z�ٓ%�cN_�
���O_i��ϰ�W���^GH�2�ѧ1�hN�w�ݒ��8Rt�������p��7z�Б�#s:�t:�,�V��]1(@�\ln��GV�]X9����;8�s��y.���4���ܜ�ȳ���*{��Ɗi��h���|�;�k���\��/�!���	�l����Y��~u~�>ģ)��Fǭ��Eí�gky�����	�� �R*<9�ж|&�l�kx)��w7�RN|�&+���U���xt��44%�Y�v����<s�vG�j�,j����#�k�v@��|�<ќZW�+5>Y���Vv���-鱧aB��I^��k�m��Cxb;ޫ#����g��yᆸj��z����4{~ꋺ���_��%�}^�]S𭁇������yZ_)(�DG���5㼾�F/k�9}�OL����/  -��VRk���k��;|�lm����u�܄:W!��q��5l�aeoh[,ՙ���2�0gר�^���1kk�H����بv���3�@�r��������:Is���{���p�Ŕ8	�=z]����R2oe'��gC�Y�7�[�ޣ {f3{�5/ǘ�U����݊HC�7��~dAEXZ@G��H��!�>�q�6�mt�'5�)�4�#/)�*'�ݖ������ଈ��?���l�-�>n�A���_8}�+˲�ߋu3��>k<��P�p􈙥숪Vq�U�R�a�.=�]������-"u�&q���KʫM����5]CN0�����Q����IB!Q]��N�p<5i������.P�{��S=�>͍��3{sN�
�cٽΪ5�a>��n(�e�ޞB���n��}��߯�#T��I	���3��w��x_�}�.w�S�ͫ!=e+�G|��đ8����$��Yk���c�k�F���}8�(��J�O�ܠ�G�g��iӝGj�n�O�`�| �,���/V�pd�?��d�0��l�tgo&�zw�`ǃ{�BO�ܫ�6S���i�K��5Á,���B�cΓ�v8'+ K�]Ϧ:��E�M˛�g��v�D�Q�Q���ǐ��[���K���Q�>T@�Vo�-�$ :�^��xQ�U�)����,!h���0�߰��N��Ҷ�+JcC�>y�
��E���S�Ʒ�M��k)Ղ��d����g4�԰ۨ���8�6��-����$~b���r���8B�l���4csԆq�뜛��y2�x{yĵ7�6���I5�^~��f�ᅋ��~��^?x숏�p� B�3����=Xܣ����v5=�d�2oXt	�z���au��\�W����٭���$sRt �*�Mx��9��5,sGB��v,W�<�NеI�*����ܦ�kJ�%��5�)��:�Pc�W�f���ԍ��gW���>�@G/��<~��c�%O�M���qTZ<�k��7�T��h�-%��M!�����̵{炠����֪�,l���j�k{&���&{���[9}�$�ʝ���1�Η���B��[2�n�si��{��	V�8�R|�u�@�����۪�9�^�{��Z��K��{��x�7���%(ue���������ꭦ�F���9S��;��o��z�@~HRf��_a��
>�]}!lkz9O���_XW��u[}VSq���V8>�I{"|Ġ<1��oʡٕ��O7�i��T3�`sX���*�P��r�i��. Y@@����8� ��	����^�
Q+Z'���k���k�K���棭3Ԁ�ñ�Jj;\Ӎ�<"�сl��<�`R[㠁��ʉ���	M�FTk����>�����Y,­颯$�!���i�f~��3ׄ0���z���dW�K�ޚ����`�\!�֤SJA�&��疭�%�&�HB��H����j1p��\jqY�ٳ[���A��gҽ�HhY�C�*'� -����=��fjރ��]��/z�PCC����NH>ۿ)�����kH�����%1���i�����[%cgϹ�S]�2)�k�~M0"o��/������@enЮ�z��xi4Q��ǐ��SC��p,O��Wt1鎕^�ν�Ti��E2��5γ�&PT��7�C^�מk=4c&E��Y9}�vu�'脙�L�5��r����X�ok��S빦U�af55[�7�������t�����xTa%�g�]{�C(2��S�,����464�ۺ
QɼeG+tڜ;1�޷O$OV��@M=R�����N������M4T�4�4дdFEa9��f����8h�`F��q�:�u�X��5E1r�&^c_�Ϸ���7�!�b�u\P��vEU���x�x��4���L��})�|�����T��>�m��F�����;���,��.g�Ū9�\@� Ŕ���t#�X��}�Э�]I�_�}�㾜Yؒ����b�jd�s��c/��k(\�G�}�I|����d-6`=|��釦N��E�X7A]J��� �뽻���ś��f���bK��x��	N�	�xF��h/b֙�X��^�d���E��vf�M�@x�.�B/r�)@�L��tFF0AB���#��P���d2rׂ~5�t��3"��_�%'|\���Ʒ�Ζj÷v���g�h�H>���'t�5f��3O����g����Y���?[4��_��ؙ㾽pe5�o�:rt��)#�en��ޚq��qGw������}!]%񀣢�WЀ��H�ح�!��}�w����f�`��<͍s���e�ۆH@x��9�!�L����l\�!�$�/V�p�U�P��,�-����5�\T6؂�,.��Z�c"��fT/,�v���I�t"��ʎ�c��w��llFJG1ڹ�,�!_[Fz���Ҋ�ǯaλJ�Z����;4o�t��ّ옪�ۉ��'__m����f�s=�y~y��=�<�}m�hj)"ƚ)��
h@j�2(V����s�z����o>ǖv�Ai����WJ��j�*O���KÍ,o�j���7L��^U�[m��ב~Sj���)1A
.��g���(y��6��!�	z����>�և�}�pހ����t�Ū�Izt��(�S�)��L����<�ŇU��P���HT��lf�g��=� ��M��k�	Ɨ�I�IM2�J4*�v>o�����$�d��dǔ�W\��������T�0�+ !>	Q	�{%���ƁF�[\m�$��S�͵��I�� {yG�<-�����4��@k���z>���@ޥI>��hS�Mݖ.Ou��E��y�2�]�����1�!��!�9�嵨z�z����z��̠��l�{H{��s�- �<����DF��)"Ǉ�k��3�OS9}p�-�4b��nSN�O@�:;^+�&泹����v��<~�3��G�s�؇���Ue�p��&'�ʠST��k��)8�]<^n�� @T��طq��t��C�PB������|���{	 e�w[�u�+��g)ٹ��R>#6l��~��b��ݴɧ۠δa:�mg)nm��g��`�MW�}���!�)�Z��n���6)S2uvJΓHx�-�[���,���&g]��4n�;�N�I��{,��T�zۯ�"'�`~h�y�<��W�8S#w���s6i`uM�2kp%����)��fu؂'�A�E�нy�� ���:wNtٗ���.>7˺+޽�SE\�s�⌜]ts�UbEq�t!o��.�<���$����q6 �02���햯�{B,�l���c6�*[;sf�δ�gdӑ�̲$h[ɻ=����/^KC��KK���Wf�MEݽ�0˖C͑��9�t�b-wf����M��[D��⫍g*��"	w�f+y�k��*�w�v<�x�lɯ�m]�H3�!G��a=�,���+�w<���ѩ
�.v�':�L�ԇG:ܹ�^��{�ӟT=�%�q�p�4]A��D֗��J���YT�͍�c��.�4j�	�ٵΖ���הۤ�J�NX�f�.�����2�E}�x9�r�G0��ټ��,�����D���%��q�т��Wa�Pyx��a���y��u�X�ta�/W@
�k���kG�-�I��2��2�J��ař�����:�_8	�1�
�r^��P�1�2���ӆ����*�u���l(��m5��p�縃�2�v8H�]opv�/u����G�{��� /20��.��]1����;PF�-��"n:�u[;��؁����ս���,�"5 \�����BS��~�i�N�X��cڏg�\C4g}�B� dqJY��5�h��'d�7j�M���$��S�������`��V��{Se�e��l�0�m�t&ooJ�/.�^� ��^���&lz8@fq�]��{��f|�{C��U�5�������6��[��F��W<k��.ɪ�����[q�3����}�t;�k9�ܔ4QQtTf������f-�D/��^ �vVÛ� %�g6�枷�k8����m+�cb��۲\>F����ӣ�ٹ&ES1!'.�r����5�5��{�^��X�N�f��])��*X�]��Ɵ<��f��k�`���i(W+�IV���ͳ�ҐKj5ۜ�n���ڎ�F��sz-FJL���E/��>fy�� h����ٷ�x����ɜ��jI�|�^�-�5�� �&vmv�\�z-S���aN�������tvdѠ'�7����d`�^B�ӊV%����9�f1D/j�}.6D]��t�l����y�UY�Jm���q��`�M�����0��1˾�k���E�@v��$��˺3��'\��`�.�6��-۳7_8����(#>���3}�dfe�J�����?�H��HL���7��q�~뫌G��77n�[�7��׏<x�۷��,��I��L?{�a�(Д���7o���w��o^<x��Ǐ^�:�H@���J�)0�%�wD?�e��#���˻��焰��;���Iliӏ�8��׏<x��ׯ��A�%3������.nC��wt���RBLiӎ8�޼x��Ǐ�x�H_��Q&a�4(O�vB
{�bC7w|\&6!*�]1,��L,"$%4u��1���$	ɏ��}����ሠ���r�PbH{��g777&�3���,��b�ow)B�$�BD�L;}z�/��q# _]ך�&c�tDf!ݹ& {���;Q!�7:A)�G��"I	���<v8@�D 7�v�P�A�8�:�)'����r����� ��vm�M�P8���V#-�`��	�[���`�̗�9e��%ә1���U���Grܹ���M9GV���l޼ƥ+�_0��{y���е����o�ALP�M8�L q0�l�e�>I���ǈ� @�X$0L����bxKa��x0�Ii���CE�X>m/����U�U���dF?j)hZ���v�m�Y�vڻR֨���x �< E0=}T�0�f����m��\��0(��Jw�$:�M^}\�MY�ax�s�O�q�mP����������Ѳ:�sr ��Y���dz��~A�!��5�92|�� de�$㹏M0�(��fʢ�M��Ͻ��ۗo�՟b��`be?�>(��$(�o�&d��$6=�����>�/Ֆ�ۛ22:�!]�����TwP��:����*U�x�K�Պza��)��5��q��Cr��m�n�昃79�6���N����!��cG�r�^Z\�א	��Bl�k{�d_F!�Q��T��ci��췖[q��{rdԖH5$g|�C2,�~��4_��R�9���j��n'��gD�N]�co����2[��'�'ƿv������x��g/�� ���&�l+�;BƘ�*�u1'P�;����BO�>�G~�k%���ί_�fH�aUs
kvLنT���A|��c����;Z�#=��l�j �E=��|D���,�������;�R~^�8��O�Oճ�h.�1d��~�a���y����yن���}����gFi�}p��� vܛ�wp�3�ԧ����։1�Į�����2�/��\�i�7 = ���a�E׻3�)`�K+���|d+�S��'�5��ttݖo*n��W�a��[3R�`n�� \���C㲰���c������gl�]��RDlW����������
����*�
 H�y�y�>y��X��td�7H��#���ٮ��Сv���ym��5\�^c9�c�ϹK�gOy	nY��?���m=��S"���0�H�#f�PHO䤿(��~Ƿ��Ҳ�S�9S�ᕆ�u.�&̉5f�
��K��CY�\矛��P�SøymZ��Vt.�<������y�d�~0�=���6�ؗ��&G_G�⨰�Z��3~�Z�5��6v����Y�J^�(XZ} ��45��Bϧ������ⳋ�V��������ة�۶��/a����{}ک��b���sۿH��	�41� @|O>�fW"��&�z�xt�㊇Z��]��*�uW{]��9]�<��F��q��A]�#0���)]-�d��O"0d8������|Nz��|k��-��ϻ�c�9=#X����t���z����,�-սj���G����B�����p;T�1��v�1�Xtc��ȶ	�n�%��AP}9�3��hg��Hw��`:{�0���2ji��3������w�?�t�s��cY-jW��W2���j@�#�626���[��]l9pg�ĭ��.P4��?UU�_cW`���X�׶wm�'�<�>�n��ؾn�"�.i�P�&͞�;Uq�it��b�췶��� ��T�t^�kX7j��v�nl�;qTC��������ޥ�L�J�=�,�G��h��i�Z������ �,���H�\�����=�_;�I$޵��PS������!�'���&���"ڼ7#�2�t����U	�H�i���l����H��]?c�N81%�
Lg�O:ld��>qZǁ��`�4��X(�-f\����f�]��[�/T҉RQp���u�)���pc�Η�ıty:�g)e�Gcqc/>xE��ėW�e0MAIT.�f���^���[����W�*�q_T�*�P�{���m,�"�}����ıZ ������p��uG!`*�~S��ZZ�5�I�F��bū���R�*~^�`�TV�J�\�L/ܪQu��LkP��NX��?K�g5U�d?]g�κz�
^	ibǟ�Õ&پ�&�S��/��=q�K'洠�t�FO���N�����޵�����A�5W��������tc��釤a��`qTa⦃�y5V�\��A��o+(�b 4���U���R:�� r��8W�}aß��ֿTĶ*"Yw���s�CD��^ig�O{��^H�k�S���J���.q�_�<5ු4p/_�vzGW5�f�-˺���\7����b>��m�!���*������@��:?������ݶ^�~Ϫr���tL#��V���Ar�!Ѯ��ʔF��pC+m7J��JwZ���t�t�}@��͗�vRmvS�6d	"`�o�s�97~�5�̯	�r*B
��hA*%7nڮmhش7n��ͦ���ڬkm����m�Î-%�-��v��E��#�6F���>�]�NvT�"uP(�c�(k�������{F��?���.��L�s����P��~�n���'��WI:�Jtx��A���>3z�0����^\t=��+�*��=6�	q�|��l��_��,!�\��- �'��x�e>vl�X3�:Ϭb��ܵV�o�}��z)鏚L��N�o����D�͒�[��ifMի��twl����B�9�+Ȳ��6������<<�CN������T��Y���<�:�se;�C+�Q���%�J�t~㖨�@����X���?��/e�S1ܒv���nGP��s��B�d�Ʈ��i�5Z�/Et��V��z������ǚ�$�D���떄�-Do=�@�&��t�4ĲO`$�w�F�R����t��	&��Mڽe�+_�a�V�g���<E��AȭgP�ľ�D�E@�%t��R��v{�Ô��'.�B�/}0M�zm�q��τ�|���O�g�č�T��LW1q�U>�{#��E�N�2�5ۧv�9o:�� ҥ�]6ow�P#+��7!�&�R����6��N�v)}u��+Y�b���2�;1�-�M�#�]hS&V��,��)�Z�NX��ˌù]����"�};We+���iЧS�\��y����jn���
&���E2)�����i����������m�j���mZ�Vɇ��`��g%�Ji�3�y�K�uvZ�Y��A))3Q�2Ee�Bd�J�=>#�~��,TD�y���A�������/�ϪhO}Ej�Q=��l��Sk��Q������8�"7_�l]��T��=0�B|ױvG=�]����x��0c�ڭ��Ț1���La�%�%�V�c�Cqj�!����W�U�zW	x�?EN��L�O�:�H���wQk�1�E�.�/&��L�el[��c�l��Ę<���m��3�*��C�~/R��"Ԋ�h��_�[����0k`q-� 
���B�ӥ�>F��� ��}\�B ���~�p�� *�^��O�fbX-�W[	�y�'�gn�T�߰�Z�XdT)���E�
y��\Ԅ�X��ב���A|-�2gfk�G����B�kG�3z	"ÝS���|�fD
z@����5��Y�.�m��B�s�F0�-��ڡ5}%:Nm���%�_<�����k��"����[�mO�Zqm���v���	���E7z|rU8���ɫ�d�����/"��	 /+�:i�w��>���r���T��ж�'E^�n�;(^�8ȼ�㽨�����l+G
�v�0��R�-�Ծ�C�~C�Z��#3��ax��Z�ګ�AK�[�& ���\�l�k^v�*�9\0�fHcyZm�'�	sycw-�W_�UW��S��J���ƚTJi�Q�� F� �L�ϛ��w�|1������zaQp׮m�ˡ'ƾ�A:��A]Z�@�[��׬��;Z2Ԟp�}�w��V�b�Pq�~0OT|9Q���-mWZ�t � �H��B�F�1X3����w�S.���ذn2i퓿�����
�!��)�lҷ㺈��n��N暺h�,w�su}^��)��R�$^[����?X�� ���	�n�y���jBe����,�Gbzv��c��@�	�/��u
k�RUI���v`0���*�Ɔ��雗�b:WX�(s�[�l��v�ڔ^��7����˾��ܤm{�yHHD�ْ�z�87�{�bY��>�O�-ڤt�>�b;=}I�P�熳P��PX��P�S�B���<sfD��=������h�����0���#��"�	����ʵ��c2�X>^�1t���K:7|�6a/hW���|HzBC��45���`Rn�.7�J�ǋ�-��UZ�/�����fAG��cj���2�^x/d{ĉ�(���O�_F2�l�_��_d�DI¯��߰J��� ]�gd#�h�Nyx^���}2�u�l�v�[��Z�Uu��9;M�p�]�=�A=כ����R�	�zᬠ�#���p���nB;���֞gqY��{���1m��oN9z�kn�[��q�k?���h>�Ji�Z�$i�@�,i�m�mUZ���U-�����x�V�O�F�y����c�"�zp��$�� ���>�����#q�&��c�M�����4��x�($�mƑ�\r��C;j�s�x�c]���C� `%w�X�D!������;�/�׈P�穒2i�qW�>�8��f>�"�Y�N�:�+�R�	U���C���0A�	g���>z^����*�s�V�O����F���#-笼�>���)��£�maeH��~B� ��P�_Ѓ�b�=������enқ:z�r��Q���g���Ό2�{lfZ�?�9D���~a���VL{<�KrH�曶�_G�]�ݽX��P������zi���S�l�{k�`���	�Z��9V5h5����.������M���*S��Yn>�w��A�)7����ob����7=&%��|K��Z�C���J}6e ����y�>�>�r�K�~���m��,�v�����ш@��E��~J�=AO�$��ޟML9L,t�<S��~n��R.��l�0)�����)B�����f�j.;Yb��Ok%<������ZT���g���s*l�5Su'�Y���B��E!ga�7�k6'}�y�����v_d
t���o�eJr.�>ç
ͣo�=��9f��S�Lu��ܙ��&�3g�[>�j$�~�F� ����"���*(�jn�[nm�Z��M�l��H��) �(� ������o�J�@�%'��������<�7U���h���l����1�����\vbu���p��qS^�t>�0�GXY���B�C����H�Y��ӣ3�	���xU����Dt�5��
�D:���Q`���9����v���!��0l���Ķ&���*�7����+ѹI�q2��r^�ȥ�����Dd�XDwŃ[t|�քWJ3ż��ʴc�\Z��'Ԣy��=#'鋍��0o@�-w-9�e@� �����N���-�9ku���t	i�#Л<�B<��&��⸎hj��o���V�{h�nc��	�!�(T^_hXl��_�̲��t�x-��\�BϽ5bAQ�����;�]�@.%1ün�z��0EV�]��E�}ܵ����X���'�/V�r=�u�$I/���v�<�nk� 7�A�ry�Oc�O`�E7������x�"KH#�/O�')���O��kډ�m�d�v5z3�U2�ݡؽ3�S�$rC�E���ƅ^��hb��Ov�ȝ�l,2F({��/3��dŬ�>T2K��&�qt�c7܌-޳ܰs�#�9�=��oϘ�@�q�Y���񛛆>��m��j���Ycf��IӍ�JeCݻћ2�y�Vn�Jf�ǹ�<�yQVu�������e�z�������y[*IZ��>�AP�Ɣ76�ݻZ�Q��ݻU�T*1��J Ȉ$�"AH��+7Z�P��ϢOa��7
M��b�h*n«�#=��
zEl�s��!5X�ޤ�2�K�]8¼z3
�Ji>TIޛ��l���E}U+�͛,���!b%��α¿`�R��:e�D�����eȔ�oy�̺:��O�������ճ��*��bN0����H�!0��$TyQ	�{�.�"��ޚ��=.�VNHx��ວ���-L���t�N��.�Hf����_>��9#`��q;ԩ'+m;M�����T��	�Or��Q�<Û����#ϯl+�(b6����m��ʷ�Ɖ�nqj�D�@�5ڝ���^&-lr��^��ӑ,3Y�xZǝ�a���^� �?Kj]ڑ���O3P�ν&6��ǵ���N��@'���b���ܚVh�'��EےqAD���|���/|՟zDo�Yu�`KM&�T���{��ѥ>��dg=;�R�nE��E\L�x�>�T�{B�(h��R!a���>���2��Yc��U�f	�:��F�#�����~�_x\�_5��A����Y�!�>�})ߖ��.>�=���Y����g������J&n<D��ϧ�v;pk|yͰe��)�HY���/Ӂ��J{���b=LYu���l�S���c��5��4Ԕ��]t��E�k!\�L˔&s{���-Ջ�L����lT����)�	Q��h��{iDǗ���K�w2�움������ۭW5�ݗV�Ѷ�v�V�VJ�b�X�ѣj����(r����W~��O�=�.�B52��^��C��[_C>���>�	Z��IZ񛽩����@�J�:�G�{̐�a�)�Et�!.?���e���gT�S\5 ���ht���\��<�t�M�����0z1��4��^Z\��2(X�fv`����{��v���ȃ
�R��D	rr���-�<g�d�ԑ��=f�2o>khNfM��ޟi/=}������l;�#T��t�u�eΓ�gl ����mW�Z���GI[�2r��b���z�	�!�+���_b���BOTO�d��T@�	`=+E�3r�I�S9
�v7�?;� ��S8D�ܨ�;,�M��;/���|~~w���-��ܦ��Y�L_�KT�Z�n�]�E�]�^'\�M�A(��S�S�m
�q�!��:N�!��3Tf�Tlj�߃�b�W|��|3 �g��#�7���t�/��qF"fS#E����I�gs�1S��w�{赭�vA��9"�zQ�����)�u�n�ZF.iG���;�6�x<U/��7�w!��G�+�U�����Z��L�	1F�b& 8��|V����������7�5����:`���-�d���}hɳ�t����*�]��ݽ�u�땛�f�p�f����b"o�F�3A�;;��*p�mm0���
�c�6�k��(4]^�-�$�i�5����vu�ݴ3f�]���+j���b]Zk;�m���},N��m���q}�<k�8r��7�K�o���%�f��e�H�k���8�v�r���W��Q�olf�l���:�\ݵ�fH�m��/��K�2��5�ǐ�Q��.V@����G���9rv_Urb���w�@u��2�7�}�{l�/L�E�[}�Bw����8�N�X�j��ߘ�$��b�:�{� �o%����\&72�]������H(猔�hg[���vC���̪�ݮ���͈�O3�Vx���;��5B�Vv�Z��4e9K��Ӝ���dcO>�A7����ɓ^L����k��8Tk8��d��ד�} ���d���Q}�Y��`���1,X���kn�6v,���2�'o�.ܭڱ��̜3�+�׃^ŏ��x�5	��Q�N�`p|1	
>���F���[��s��S���E�PbbU��;F���nu��Iy¯uҫ�ң�n�,k����\�v��M��A.$f&��ì=�b��S59=�)q�0�����N*�^0�k{;7�+�����1u�:Ei��,���D!Bz�QQ��-]r�X��ﻨɼ��h�l��3��?�����(%r����ok!8�"�S�
o9tw^����y,�m?��P��x���-N�p���U���\�)�m"31p�qHc��ȫ=�y5�#k�����5�Q�s&�&�%��{sd1]����������r	�,ř�E�9���d)a�D*33R={ɞ�`VxG��L��&��V����5�x�Q�䜹l@�0��|g�!Ӧ�[Cw�)ZK�G�
S/��� ��C���Z�V@)�O��J��OK�Z,&��@��3�M�-R�fB ����שs<�����-��r��A�'��C�ik�3�g�h�oMd}�Qk�p���ӣ�����`�"77����9,p���u�̳{Xf,'��5��(�E����������&��pZ��*������o�{�[����2��n���yה;l�}X��Nᇖb��%�Ł�7B"��>rI�"qx�+��^����אT���l&	�ۛ�v��ܸ�I��"�<�&-�9;��㻾�̀gq2�L4�Tۺ�Ѩ<3�u@�;���1t��N��aу*\��,=�����,���!X�B�@�X=Z�֓��VݺyV����v �n�W���Tz;tN����,*�ejK7������B������'��h��`�I�ͻ\{�1�#�4ӧo��v�Ǐ<x�����f?]���8�D�����H�4�"I@b�H�Ri}wS��:|q�v��Ǐ<x����#"��FKE��10�$2,!���؁	5����c�8��׏<x��׽$ I(�df~�A����wBB~7h(1�S�nl�#$����37oo����;z��Ǐ=xc$$�! 0�J��aIQ�����q	#4�,��&D��4��%>w	2Y����^��Ɍ	��u���'�\ł����c`};2�_mtш�YQ�64b̑4B	����j{�/u؊�D͊D0�R|u��11!��O���!�K`d�I����LЙ�L&M�ْm|���%�6I/�p0ZC#(S*�ĂH?I�ު�R.Y͑�5A�����K�}&����p�9�Q3"ud��WZS!��P���O�I��ɥs��<'�T�*G� ���i�F� 
i�
�(H)"
�"�|���y+��yª�Vߗ>ϥ�{���x�~�R'������D�5�JNМW������Y�:N͖�޶�N�e0J�^��'�ʹ"6�З����,Cz�)��%E�Z��2Y��������t��m���O)J��<��0���2�2)S��q����T�My��[;=����y׹B/m	����:��n�<�p�"��	(�@��Ȫ�(�����C��#5�����S�hc�X���\�#L�;~R9P* lVa?�Ba6�oZȇ���G�m��\���=0ǱE"i�'=<D����ڟ�����5�-����;�.��4B��m�F��M��P�_��HϾf�!>TD�.����'⦜��[�ֆ��q��a�J�����V��C�c�b��l	�"ˉp�Խ[�P����<�Kn9.����C��Z����輻����=��}KN�-V(*������S��暨A�	�%�=��̝���hy���[�N�Գ��&:�X/=��.]5�S)���l���a��ʏ��
���I�wUig&�����\@ ��=&�ˮP7�"7Kz":wO����_3�O��{� ��3�32��İBp���u�_B���*	��{��ź6M��XQ��w���O�h�MH{��S���v�*r���n����w��6f_���E�?f�
�$#i�bi� ��)�"�(�H � �o���7�1�Q#F�3/~:�V��&Ae^�U�kOc�Y'�#�թ�!�L���eV|C55��O�3ec��"��zЂ�O�4U{g[���S��0L���@FM��S:V%RUW+k���=}U[�Kj-$rӆt9���>��)��Y�f�"�G<HSޭ�ll�X���zp��k7o�� L^gEǧo+���ǘ���"�5�<�HS�u�F�QtÔ���b�:�43���Tlg����	��003��7d�M�,τ���q���Cߨ3-S�41h�+��)��n�����7� �����������߮H����surǖ�|���st�m������V�X�C��di��߱�>Ct�0��-��'v�?���o;]�t�@5t@�� �s��PKܼu)�f���l:��7 `L���ԫ�)v�'Bzu��C�e����'e�d��<�y��g��0;*j�����E�bSXj��V ̄	���A�._H�㔧�G��j-���:���P�ݏ�5~�s	*�Ќ��Ed��1bP����8��o*�"A'J�e�H�ː��9�CҸ�����]qVm��%n�u�����#Y�9�rn�"��/�bn���iά���ݥaMwЫ�ٶӍW�`�B7ӢU�т��ꪣ��
�i�@��i���Z��m��VY�lUlU��$|>�+٧Q<�ݝn���g6���!91T�vE�"�������,���v!=ɛ>��p�٢�� ��ۻF�C�M{�s۬D��oS0,�?��ܵ�n
c���?�����1J:�˝���\���Od���pj����{:Í@#4�;���Yz�<۳e� Pz`��<ūw���n{��FuM�Oh���=R���@�!ȟ �ҝ`Z�Kh=����{gS�)�,8�1�r����%#�N.�ݺF��ɥ+���v��	Mw�Pd��Q%�ӌ(�EZ�Si�Ֆ{���Q�Ѽ��3%,H�"Xc��{�dO�G�N���\o<2�I)�Q�D�ap�=���d����7굜��+�)ZN��!>B� T!�"]ڏ���>^�P��15�S�z���F�j���oJkk����H�����Lz#�3��
zE�=K����x�v�fy��&�jl C�-�@O�g�,�<�4�scs{/���׶���1����<�{����������ݗk��P��-?,O#�V������?���}��B}��i���O��8Gߎ��i��7�+�靃.gls�v���j�����D��d�~��s�*��kj΅Ը-��\��`�;vMHP�yB��~�}�Z0�k1O�R9�/O.��u 0_17�\c�o�4\9���5�`~���p��7}IɅ�s~�}(��4��IQP�P�4�PA�4�1� d@�$P�y�y���|b�E�����t�ƨ^ǩ:�<y�yf.4��K֨�*��ح��{l�}�hB`���[{=2']P���^��-|c�zz���/-O�Dᚕ1��S�Z��di�����I,8���ු9��^�F����H��B%������z�\�]��&�1�����:r�P�����\��z200+�����x�1k��wy$�y��oW\m�EkgL��w��҇W��R9m.7�*(���a8guO�0%�3v�`=]�{�l�@�]Nٯ
&%=0��>&����b�P�>�&`BU!]�zq���TֶẰ�H�[��0�b�x�Ⱦ���ܩ^͔^���r�v���9��E;�P�����rغ2���H���Q�zl.�����\����ū�,��FCM��,Gp&��}n�(oB���x8�]*����X�w5T��H{r���{��;a�@�9U�}A����s/-:�ù�����D�xT�?W�1	�ׅ��Q�����&�u�y��뒥�y����"�6� E*�y�(��;�Q/#�5n]��a-�J���O98%�˭K�r���t}��c8c9qj;)-�VM�Ϟv���r���f��� 1]�]H�9���1�H��t�a�y{�77�w����s5{>���Ƅ^ݺ�TҬY�v�����n*��#"�:��������^�QP�ʚ���)Z�L)��Ʈ�Tܽz���B[��.Fa����8Ow*f7/���ӭ��Dkf��D�ZJ�̔AN+Dl�Ǧ����!���qq��B��淆\�����_Z�*�;�1*�tw���>��E���Z�T���@A�/]�j�&��ǭ,����@z�d�ϭ�7MoS���'��˜���{���=5��ZAw�:TV�ֵG@��p�E?�R_��ǖڦ)���"�c�F:�<��j��/��M�f��Rk��L���O�RC�1��@Hk���9���z)<P�#��x������.9a�U�E��N�V!����-r�u&/�F6���I05�Vw�|h1��Z|����X�����"�Uo?J��\\��گ��'��G�cꤶ5��Ģ69�@|O�%�f���s����F�.Si��T:��Ǿ0'(q��>; ���Wk�as��Ķt�}�zeo�y���m}�������g���$f����Z���v'���Er���#V����P��5Q�X9>jt��/�Pt�1��<�ڽ��7il;��{�K1�v�g�M���|�f�%�%Ӭ��x�wjY�Z��B/K�/^p]2R�;�F�f�D�W����Q;S������<]�H)R�Spĺ,��YH��J�Uq�4�P�KQd#M	QR4҂�$ ����|������n���惠��Q������U�!M9.\�!1=�b�)�)�MݽzG�f���Rr��B�H�|=#��B#ז�<���ɑK>�V���}�k�(�[�|E���S	��7�g��Y��p�j�5�J�楬�9.��(x/bTO *�:jE5,�ŏ]�@����qy3٨sw+������^��"��k�w�Q~B4�4(�v_����ꛗ��,b��-k��-\%5ߴ�L�`
�'�����]��H�4��ERNq�@^S~���V��j +���J2_!��xN��LR�����2m{b�����=���N�e]Z󹨫<�4�mbD����ϩ^+��'�} ��>�f̢���,Sި�4Q��\-�]7WJT1G���˄�s���1,T7�Y���lEl�Fk�^"��T��2��,ҥ�n��w����C��.8�|V��*,
5����9Z���_Rw�
�5�ksK�B��Yz��eAJOH��5�G����ad���^6@Z5�����=1��7z�;u��sb����[W�W*�㧱Q�Z�WD����k�H����O�52����8=�	��Q� ��f��
(�4l��p�-�������+~w|r�s���v-�ڻ2�Ė=�!��w<��N�jhK�j�j���C�N��Rk�n�Փ�WE�W%��SP��C@�D�Hsh�n�r�n�nU���b�P�s[�V��o?eA;����!4��yYn�Zl�"���_x�0��X���9ޖ@�^��ݐ|�hGO�	�].�=M�.�R�s�Ѱ�ߐ��[BdKk�����+^�T�/B|����tFF����0�W��^���Ւ+��^-(�`R�(:��3�tj|��}8��1��z:�4N$t�<�Ob�=���J�Ћ���Ә�B>W�&��{�G_�sJ>[xE��-,71W~=�<+P�ӡI�r>�[-$K�(X^��W�-3���������z����F)QP=Q��9端�
����f,�O��5�n
~30�d��/V�s��_�f�S9I�V9��/*�M��M�y���kܾ�(�������?q�5��˓�#�x�Ef��]���ǣi�wUC�lʂ���#��l�zǶv�t
w��9�ԥ�Z���wf�a�CY`~��FG�r-���"S^��A�E����s���1�ފ���2Y��m\Z�����{}X�)$�F�O�DM/����j5�lA�1,��IH�	�Ee�A_ƾyw�}�ܬ���>^��ke�]3W-�õ9���w7�������o;�\D!1r���^�����~"���y�{�N���*T��o��.���7�n�m9)h�oR�^�-�b�Ů�AA�p^���E���|*����W6��m�v�۷k��d�� 0�o � nԎ�n�V�o��p�Z�>�I8l���a�P�Cm��A�;�<�6\��1�^;���F�s�K��kgہ}�p����\c\+�'�΃��s�C���c�`��+�o���q^].���^�/�"�m�yk�W0�z,�>G��6�Q~`�:n$1b��N`�;�d7 *3�8�뭗i�(~/I�܊z�./>Al�	������=�����l��ɥ�맴g�;.���P�a�~��1-פyP����G1��������AxwT���vFaȻ��Uأ|�.�|�<�t��ȝ�B�L
m������'Z2S̨�R�嚘{�v7ۓ��5PɼtSIWּ3�� ��AC�Ɋ����^�0��W@��?O0�Ϭ�z�U
z��O�Õ<Gt�����2�����29�+��L�����>n똻$�m��sW��eU���/1٦�7ps����K�	
��a��(���oԷ|&s:j-�aK�MU,�&�r݈d�׉��T(f�[��gM}��&vX��[��ZX>�A��-὾��BS(FDM%�����&��<�����Y�� ��e6y."u�]Θ�u:�`\��E��"�5_̡���9��h��Be7�ƣ��W�.�੓e�]��'W��5R�G�Od*=�Ǥł��O^��;:�Rg��3{>��dB?MTH�BTIn�sY�u�r�HՊ���^��+��^&�M���p��CRkVU���u	�$�NnG�+�Ņz5�?����t���pz��M�ٍ���)����*M�"�?�%���r2ރ�|�HjH�a=46+���f�g4�>,nV��9JL
a��.�Ӓt���_�q��'��t�S۝㆙�,��۴��s���ٌ(�s��	�r~g�5�|5
�A�(+�z�{�;(�+5[�m($�L��\l�n�W�|5���N�U{(�b�J�QaMAm�5��y��xBz��j���H씱�GQ�,+�b�6/Ӭ��TD�M�[QN/&Xu[�����o8�p�)n��MR5_j|p��l�Tkhi����T��n�Y+n�<���{�U��)	]&`�q��ܥ�x��i�d�T�y���ُ+XEq�սN׳�G�[���.��5��^���$�J�xTg�EY�]7�@�e),Qbփ�S�b�l�ψ���PhOT{���=��U>�
��kzM?����ÊHO�o9	���C�5�K�uRd�\��&�<���W�}O|_2f詿m��H)S_���b^���^���ǜL�<f����K^�p-�8"<kG�v����30�[Vf]��w()\Ʌ"E�<���X@�'���ǉ4��KȽn�k�x�ϞnvI�j�c^Y��������s$�%�?f���B�aD�hJ�� I�9�y�����o>�4�}ѧ�S��#ʎ���Q�P�ꇋ����>s(�.<���a����5����+�g�K\�8��J�a>Y0~Ź�%�4 �����Tϐ^����zk7�܄Y��
^��5?%�*(�0*�A��{&�o �7�i�� ����dt�w얬���y�����n������K�'|��59��_ٮK�wn�%�`ynV�[]��YgY�(�ixX�<�~戗.���>��0��>z���P%�*�� �;f`��
����5|�1C,"-���3�X��=p	\11�\�:~�!M)3J��}����B[T��WS�O�6�R �J�ɹq3��\e�j�A�����\`��|�EL��e�-���{D�N1�X]x�P�Y�"ڷ �Te&8}�����1P�C\��1E�|j��e�Yg!�sq�e@��������{���.�&�� ��&�hz��oV��)흺-=B�}�W|�f}&� ��� SC��@)��6cZv�զ$��T�	�%U5����C�������8�m+oLʯ�.��Ǹ��`��r���}���uW9�2�"l�r�l�2�T|F�s��7�,����	�|�ك�in��z��E�f_L8ZG�I���ͻ=I����'.��<.*����cͲwWm1xΙW�a�bS#��qM�l�Z�8h��<9֙�xo�n�\:+�s�]��ŝR�Qf�䠚�s�F����g[���>��=���6�,?A4��Viap�IAw��T{����\\���g�q�;z��I�����1��)X	a��=���V������ű>	az�e���t�g jx�5������e�&L�ꖩJ���S��"��Yu3�iY]kA#s�S6Rf�Aht��"7�<H�����H�o����c4/z{E9:p�3��n'��K��?)���onE;�m�"q(7vD��)�8d�ª���sc��P������kr�Z�������Ū����Mj���;�4��г��L����w��7:g����+�c���y�q�5,6M&����E��T9Y]�u��)7������J��x+gp"˲��Lp<�E |@����+����utP!��/n��f�]u-۪e�s�.�T���c5�^#�ݎ�0@1a�CA�c�.�;z+�ǶfX�X�'��;���W(i�)(�"#clBl�ew D��0�=��x���g	0t4�u����c��3�-k�?1+� ���ň�{0r���l��'�Ȼ"�i߻,���e�}��go��q����]�ě|;�u�^i�ue�s��6����#�^g+םm�'���Z�M��]\�AJnM샸e�:jU�9��>;^��p��m����_-؏:�v�Gز�ҷ/�1�`�n�ɲ�s-�.�U�r�����#IF��Ǿ��ɘ���Kًqỡ�kU� uý�Uҹ��+d��u����!��7��i��V�5v\E\���{`v{��9t}.�.k��`<�p[)���U�� ����޷<�Uj󰮹�q�8�ED7���WntX
����n�f[�{�<x����E�ǖ��9Ey�-[pR�j�N�"ul�R����H��B�t� �్I�{�}+$j��)����	�H�vӰY�˃�D� ��!}W�g�f�Q5JS'r�΄�	 d��z�{nw��c�^�=���R{-5�&a������"��S6_b�T�%7p��j�>��z�-Wm�'7��d>���ބ��h0�
%����oq����o��R[�ı�HA��37��	�R��k�k������ �@>����&���L�DO�	&��j��y�����F]�7�S�~wݧYy	�� ��p�^\�D�J�v�1�� ��y���0�1�I��I$�i�>;|q�ǎߧ�<x��@����$$�2�@��%��F\"�6i}�4�����~����x��Ǐ<x���$�! �s�2}u̚`�#3BDl�#�n�M?���8��;v��Ǐ=s!#�� D�����,I��*Fj�i���$�#lcM��8�۷�<x��̨	!A�I$,G�pe{��(`V�<�_κ2{�0o��k���Q��[��^Hi-��O�i2A���h�X�#)

M#h�1�2Dm�H�N�c�Y$آ�X&U��F �Q�����n��#FK�%�c\�1n��D��RDYs����r���d��l@`��ssr��0�g\��L��!�m�8␘�L��\$8��0
1�%|�>��{/��Os���U9N�2/k=�i�԰����[�t�D�0=�Z�t�/.N�=�m���?���J�(Xq��6E/�M2K|�8�jL2m��7%���p,��؉1�� 	���p� ��p�R���zN,����|�hi�*1�����B��3y��Z�˝�r��$4��z�]:�#�9��q��:�H��O2�Iz�B�JĜ(���V`��=�5�>>+�讙%�3��SE0�m�o!ș��<9T�4u�	�QqA��eF��P-�mWа�lV>J�\��n�v�E�h5y4�[���v�[��cB���\��"C�Z�%E�S���ז0#��|@��"R���y�;řG^��j;�;��zv��Q��)���C�PN%�d��%��_+B�b��d�%����e-�+�J��4P��[ގj|�vtޏB�Q�cLߝ5l#���6ǌ�]�΋�{�/�2���Ķt@�W��7�,~�PKܽҁ����tޮa=�˺b��M�Ε�0e@���7_���b�N�>��1PS�מW[��Z���J�2�y��.�ȬAc�XxeC�����c��Q�Zo��>WHT&��/�0̅S<Q+i#~��1�է��Gs-%"���+�c���O�a�B����	`B�W(�`��M�7<��CѲ����;�F�ysdr1=��z��X)}����TP74e�0��C(���^��#���b�2�,���-�i3��Ĉ�m,���ϳ��m=��e=�rmoo(:�f��?+[;��C�����ɇ}lPy��[��n� �;#T.ޣ���A�n�Z��-��� �JٳzXMV����:4�)?ʪ��u͛�W2�u֚n��ɴ 7���֭T�BY����>����Љ���lp��ԄU��:��1}�K���L]��:e��7����K�+k�r��jT(vA��NK�Α�ޜO�^��N�cBAj�o�����4�8�q��{�KǦA���&�����Oo�S>A�;�����Fu��j�l�O��4�Gmn���-�ٚ��*�
a�����c��/�P�7���0�N��ژX��:s`͎�����8�G��G�� k�@Y�����Ѵ�0��!R?�����%��q��%��ōx��h�j)�=����_�͂�&���'"��\y� ��v��n��M���&�e��ͫS��z��S/ ��*�ܗq#:�$�Dxy���hp\Û�O,V�O����Φ���ތ��ν��c�o�,nS7H$O=�i��s����}9愎3�w�l�Ȓ n���{*s���RZϲmLzEAi�C^����.^�9Y��1���N���<|�������tjy~"~�k���8�/�"ΞI��P!{�|׍�ve|gSh0��8~����Ϭ���oc��V���3���yB��5=}%�<u�/�ږ�Z�4��V�9�ô��g%:�rszv��4��A��9K���^��S�ff�� �����齫�j��]:K�n�|��䊉���:ԼE9�sU�y�~s4y�\'��h*i���7���1�8T]IY��1!���R��4
�9��K���R!a&̊T�<�|��ipT��#'���:��E����C�:�֐_-�>����3����C�"�%�>?-3$Q���k���w9,�VǆƼ�1�}�$O�ō���N��x����ܬ$�oh�Y��"ض4t��s�h7V��6��k����v>��9s�bMGv�	�K�:�ֆ�+#"�2�^�ߺ����Q��:y���ۈ���OƊ��8}�@jMy�?���u�&�l��� �˥��cZ}�zؼ�nޗk�������fx��W��j�r�����1��!#m<Zɖ�A*�T?H�<�`��Û�裳�Q\�cb���G@��P�ғj�k��1?Sc��g�\�ٯxt��T9�;�:�,k	q~k�{ �bP��	�<9�����5@��+s"#F�^���f���z����R���,T)XU~�am`��৑CXWLU�ȧ�t[��ȹd�2�闼���,��*K�8�O��y�s�DJt���L�}E8̎�a#�}6Ҭͷ�hϨ��E6Y��O��إ��t��M�4��̵��h�
�y�V��i\&މ�B�0*�[E��{%QX�ӋO��Ɋܗ��&]���[(ZWY�}��HӔUiżi��]M���'�LP��.���N셻��ʥ�����߯�W���H�Y��}D��+�g�mX=}�ir�^�`dO��i1�1��쓷H��U�lX~��#����W����y��eOWa�L�O0�;0�P6�}d1D�˴���{��t]hkx�޶:���#g:����{��JK��
,r�}�D@Z�F�Ǳ	U�ڙ7�H�I��X��olgL�XݳX�B`.��<�A�5��h�V�����R ���e����ۍ=h�ͼƍ�k����F����=�gӄG�:a)ĉA.
�A�!���J�5��^���u��{unV�VS���B�`!��^��xjڝi�t��V��6�Hg�'�}U�W�V�J~��Yinh�a���Vw�m�6��͘��#Lu��8��@�%�EflO{��=�~�I1%"#�I����h��l�mΟ�;hVjs˭W�sW�������ӿ����_ �߼2��g���p��$'|�jc�;4K�'�W�4丫�{P�'#�̷R��z��3���χXt`br��@���D\������\��kz}���C:���[0�\�����R��7J��5�Y�2$]���QJ���`�O�O
:z�j�f����vvˉ8��,���ӝ[�V�کmc:N
k:NH�5˻T6"��p�"#�6��.�<�cq�3;��ɓ7���RlY�jb��:�7�� y������4U*�Y�eD=�giRL�)�:�!˵��"�޽V{~y�޸���?W*��æ���3A����{�0�'�k>��L��p�j3�ީ��v�E�㑮\�P� �v ���"n�pO�����7��i��
{+]��}����@�t_�Փ�6��	M��!2�,T)=�Wm
�����o9ק�]93�@�JXɐ�c�F���ڠψh�@�"y�z"TB*S2l�IT.��"���y5�QuM���K5wԨ��)I�%�j��M����*Ј����)8<f'����k��n�I�n{�z��Q�_ʪ��r-��e���HW�]�3PAS40&�z�5��>�d{:b�P��-u�#ܶ��i��i.�`ކ�	�fh��Ox�y�o�֍ɭC��q(Zޞw�l?q�O�eAb�O����>!��a�����g#}�W��]��;܉���;�[�ED}�|t�l�h�z�Q��L@����$QN.fei���>O��V��Q���g~d�r���|���.���/0��yÜ}�1-��D���<�yB��}�{.)?�*�������$qİ�V� e�$`�ԧ#�]oW��=w�[G�F���:^eܗ�t�,�8vV�`#Hǋk�����߷�8�t]�a��<�7�����?d�p	������f�J�ǎ���No�$�-Suň�2����~��/5�z�^�p����c1������C,a޿�C~�r�D;k~,�t�N�=/=#$��+���ž����Ƥv�CM�n�;j������n�a���������͝9�PR�p)�i�J��5m����Wv�i��;2�2�.�>��:Y���韵|����i��u�E�y�TY{���t�St�Xf.��k)��6��m[i�t�Ţ�=S.�y�h�7�DT/je_�e���V:�;yz2)u�eu�^Vd��],�����#��P8g=H`�u�K�ţ�(.�F���Յ�f�asKH�L��βa�@�)�k�C��e�N0-A#N��6q9�ï��1�]^]�6��A����Y��]�)1�
/�
�C��"e��`Mǻ<�c0��LmGz�P���ڦ����j�s_�!���:�U��h$W��P(T��T<q�?�z4�7��˓n[N��Ɍ��o�L���۳G��{ӿKiQ����*���O�צ;���\�\��)j�6O,��#V뷗��[5�%�P.�ǊT�yP#m���H��c����;vlݗӰ|�Iѻ@�A6�*���b�����4��Z��� ×c�{�� �<Q����Mk�uL�1�] �r�:�@<��^��,�A�zr�Ib�WgE��!���%׮��os��#�ȏ�7��No����M� �q�R{��V[��A��$l�sI>��_<�4Ut���/^�!�������=A���6��I���ς<ja�;JAq�5�h�c��yה�`kVj�fӱLM�L�b;��w5�w�׋��,yi��j"p}��\B���;�|7yO��&0��w;�]�A.�g#;
�u/RC��I�VQ��b�B�Hǖ�}#����'eR͏yI"�+�� (�"6'��i�����P���4���bȜ��وg]$�����5ݘ�/�_[$f��us�P�.�.�n�Qx��/1���y��S���xN���_FHh�
�!���мx���[`�TD�����Iܝ�x�"Ԍ��p;B��񁷽s���1���CJ*��칤U&�0��>��M]��Q}Q,թ�g}#���A��^���%=0�����9��g�v_G#(���tǲ��k�(ҡz�	�(S����L�&�����u�&��y%�%�]��2�h������z�c,m�Bq�U��>�� h�ǨE�aKv���"[�"\���W¢�(d=�k^c��R��Q�P�u�֮� ��	�  �g�g:{P���XlU�0a���xB�Ʀ9�9��qi�~�؆���-_c�h���o�A�c0��VCܥy��Vy#�л��}�C��!��t�`���x��gmHټ.�a8�i<����:�Zw%����1���;u��ws���љ� �.(�k
����r���暧N[����m��ĺh\�az��ڍ�dx �Z˗uc=�����q��K��^B��9V�������tͧ�\�5s76�j0},U�0X�R%r��Qۜn��yjg�g���%�eOk�i�\뻃?wkZ��Ǜ}^�bdKkH؏?�K���8�.�#A?�(�!J����74_����V���o����a���N��Ұ��j/����]!�@��Q4'�Q�T���q����j���e&Dl}q���-h���|��i���Sء��2O�#��ՕK�r��v���k^�@���y u?����_�\j�^;\�ۭ�O<�ڪ��Y՝ܘRk�xen�>�=1�����I��n��Ʋ5(6=^}�S�t��*׀����Ս�Qځ[ӥ��J����n�����֞zwx������d�[�a�R���5����0lڑS���q@q�U��<��-#����?��q�¯�jtş��+�k�e^�f\�@b�{�ʝ%�]J1=����Q䓳.��pE+��o_�Q���npH;�Xm����9beq�3;��Uz��2&���k��O�ɘ��e쮔mL��!��d����FCI&�{�b\J�����<~1�c0w|��<�2��w�k���i��f�u�鷈_�t�]f�����?�|O[��=j>h�\��W0M@e%C�1�x��8�֓�q��
�Q�SXz��g���c�Lx= _����2}�����9��3l8�@�z�LK�6��S�r��/k<=��rnu��ɥ$�1�� �~Rl��Ώ����I�Dn�F1��؅�\*Cy��;7o�1)�����g�)5�ʈZŖ��\
��lS*d������Ws�����<
�7�J��[�\����t�dl:j(*��'1���f����xv�u�¬A̱	'��k1F�Ϯ�l���)�dECs��g�6�Ca{�����4���.ȥ���j�P<����}3��D���|:o,U-I�*>=v�'���{��V�Sb�k�u#�+ד(��ǐ�P��Gپ��1Dy�_F�%�oD�VT�	��n��%����S4=�嬤��¼�*���I���Q��>C��}�����\��su1��#m�m'}���Z�C�1R�ҏL-�/}�=�����;Ek��]|n����
���#A�g@�����0��p��ј�e��Z[�۷����r�T�	�;Fg+.�#��I��!�K�z�X��@�󛿥IO︊�|�	�}O�.�7�w�a��vh�'�7Fm=��D��&��Ka�-Բ�ĳ^��ԫo9�`����u~���0��y��n�Y��¨�<���϶���]s>Ә���F;�0����� ~2�?�k�>���};�kU6�:��O@�^���.����e���T+���pN%�>��;p=�mÞխ���2��Ǿ� ��>�!�ȇ�s^�0�Y�z��*�=z�k�e#uo���t�o�V�|�%姳��SU�ݗ�]+^���?����F��=��';�بw�r�Q�D�.�9�+1����>�-���7��!�������/I�U���:`�:����.V�-Ǭ��V�n�����r��Sн��j�Q�@����
d��_5�H�|�0Mn�%'�_O��*}��^d�ftC26�e���;��^=^�� IӲ4,�ׁ�&�^�=��=�py�f�ʿn]��M��~�s�zrCG޵V½/Y����I��~�p��tFc	��pS�������\�^���t�뱩��3��1J=w)�ؙ��Ȏ5�~��{��j_��4:��L�tNK��R���Us��{`@v`��E�Bc��s��OG�r�dҒ��8/���{d$ Ô^ۙ��y�/]��4���2���n���3D�[�e�Z:Ȥ۴a)�YP�Ʊ�]��S*��2w>�p���t�ob=$ʔN��wKkEEPH�m��n-�tմlL��fծ��Μ�b���d��p�z�1��E��{qxL���)E<QL�=6�n�Ng�0a�К�XP��!�2m^�f�}G��5c���ĺxzǨ�0w{�J\�_���3�.�-����E�o{��/E�|��[�Ȟt�<��s���-��K�@p���Sj�Ζ��X7���3�^��2�Y����w�P��(=V����vY�+B���:d��W���cʃ�ㄤp�ZWI)��!r�ֱ��0�Ԕz����mިk�u�I��� �(ƫ[BM�GF�h���31��
��ou����n��8���|d:��7��e˶�*/�K���ݎ�.>w
bU[5�1VK�`�sOI���M����X�f��XY��C��(����T�j�f"E�9m��V�������#Y~�v�",Z�J���˯)�+���k*Ld����E`P�9��MX0���7�=�a��Y�= ����=��n�|��� ����z�c����價'R�2�АW�O�:��p�h't]���zA���☠O#��6��1�;|6n�o���d����Ãk��f/'�ɧ�����D[@��A�C�YW[�ΰ�H5)_�� �gN|
�zN�)F97ьٸ-��=c;4�B�.u��K9 �P�pp!���ۿAW�$M�I�����P�ғxۍV�LO3�-	s;t��W,^�c՚���.b�ٷ;&L��v�Zg{)j��K�]�4V'��
�&�e@�_R VHo:gJN���/v��XC��}�T:�^������<2 �&Q�k{vJ�傹H��&��K��$Z����5v��0�D����x�ۇ�6�)vC3��˨�=����b
�E9�.��	�'����I��VZ��ĺ�-�C7Ma2���-�\K�+C���戯�Gi�]W�s�;������A
�uF��'ϗDuj�WQnx�2�-7|{m�Vv˥�m\KB0�wl�uz���c���PI���f�"�e7/�V�N:}�W^��,��n��ݢ���CΥ�^���c�ɫ:b��)ӕ�\R�����BcP�����w�Ю���dSe�k5���~{˶��8��E�Lښ8���)�cp:7N�p^ξy��a��S� ��&�������m�	X��������9�7��S\�j$v>8Gp��'��43I�����q���`��-�z��C��'�v�WGn�^[���g��%�1����?\)�c6� 2tQ�,��ZI�;!µZ�y�{�o�-I%¤dddd$�}w�"/�����nZ6��u$�		%1��6��ׯ;z��Ǐ��8@�FFFH�D���،�S�X��i��q�<v��Ǐ=s!"�I�4Ie�!�o�����cR.�c$"HSi�>��ǎ޼x��ǯ?j#_��d����9i�����<�(�("�i�4��q�ǎݽx��Ǯ�p����JlL�ݯ޺�}�޷���NW�v�r5��j����r��Ɗ�I�5���\�\d�BQRQk��7�\��d5F�Ɖ�D���ϯ{h�ˆ��AW�(���6 )����&1�ʹh�"M>��	��T���$.\���R&Wxޏ=̳/:����T9ٓ���Z NɎ�n�z�R�5���݃����۽:���N�Z�"J�n�P����c�w+��g��w=��a���^�ֻ�c~7
0!e�_&��G�Έ�H��nX`�Zm��Pnh������gU�b�J{׾t�^E��H�w*iM'�D�>s澿N3
� D^|�ͩ�Pg
�6�U����n���E8[�-���)�W�^{�+���V�9�<��S�Y�Q&�qRۇFK��u?_n�de�9�{&�=�Ie�Zp^�'���,בy���`cm�S���(�[Y�ܮ�KZP0|<�7^qY�3{�W	��!1\�$�U�9��Yz|�:R���I���ѵ�PN$S�|�F1���.'�P�M̋���@�Y�����ls�m��J�1l$� 4p�C5y�Þk�!�}�Dk���g�Mk��<ǎ��,�S��M��e��}վ�^�j��{w
C���
�#�q1z~��>���neK��T����a��O��p��)��vz�*�Fи�q���@|!�X~�4y{���y査�M�ۏcwA~d(���MѬr}ǧ�Fg�y>Կ�m���(P@��L����Qo~����`j�7LA�`�����Yt�SgD��q�>�*�y=LK�*�5_,9��/�zq��ݬ��,V43���3X�����n=��BK^D;�̎���|x�h���چ��sn�W�1�����H)L=��c 0i��y��7����Ҍ4K��"ԴS�.}�<�+�8�A�?r��&��(u�F�W�A �2��]T�zm���s�=%鏁k�u�G���6�k��}��T�掘�d���|��4LԦ�	��j�B��"Hp��3����A��O�k�SRj�����>j�dD�قa'�
⻞[���ӻ��ۚmxj�O���>Y��A�>�Gܙ��zi镹�5��ȇ�}��%v(,�vI{����>�!�/�5�j�#��b ݪ"��;M�ލ#�m_y���v�Ωe���cvU=j˒�w^0��)�k�$���A>_zn���=��Y\�xJ��)Yo���F�_�g���
�\Α'�]�t���*߶4Ա�p'*��3�����B>��;�Pj���2!7s�']����AN)�)�٬��M�K9뺎j��W<ޑ�|k	�4�a�e5�o�@͕I�77�Ht	/�F�M�mR�<��!�r�U ���Ű�va�yl����!X��F�Bg|��*�'��U�6+W�*�={�O�whN�o���+u����2Vu�]��Q�����n�X����ь�˝J��&���zXӎ{�o/'+Wo5�Nr�� t��[s�Bz�g��=u���Yq��ƞ>�aΤ�:�n�b�&���7�nI��&Y+Z�Ԧ��1�a��^����O-?�n��=������%�{}�y|y]E����i�I�Yᩍ7�X��vDꔁ׀�M�@O��=	�Jct�I-��8�6��Vfkt*���3�;^Y�Eח�l2�_/|��A�}��HHO�����xTco��R�+u�T��^��Iq|T��L�89��*�������N�1�;��.Βڇf����0��J8q^�2�^��s`Mg�����]�	{g�ʞ`�cG�._��w��Qણ�+���ᓹ��ú'��O���-�*��1�x�{�7OlM��b-�8��SrтZCWm�k��H[[Hg+� ���0���M�}o�KF|�R&�=E��)�\�u���Aϧ=��&;1:v��c���W�#��?z�%
�?`W��D(R}��B��I�κ�3�W���1\�=�8�l�'>��3��f���D�e��W��l�y��
vF��i�Өڍg���
�������I�\5t�}DZ^3�æ�e|��5H�p���K�v1�BP���7�v�%�"�;T�j��$��9���ҝL���ӌ&��^]mb��?��u�m:�q�{����<��_D�'H|�5ל��������u�:�a)%�L���M='��䫴tIzP�=2����W��t�w��<ɚxN�3k44��]N��BԆ��6�U�l����rT���3�M�]2�=�.��xz�xxxxy��嶹Ze�����5��i��/l����֟{����!2�_�%b���ΰ��e�X�Pg�b�|������m���_tx�i!�����w��>�b4��q��f�|��Jq��Xͼ�m�W_����j���jF�+��I�Q|�|�0y��A�y�?5re�L�)�"�]�A6��<Kr{�Ž@ec��lE�+����H���. o�Y�փ�f���f���]�1gN����Ƅ�G*�Z��ܮw푷�;�|IT���b�{;ac�u�>fY�x�셍˺�4_��k|�li��v-)0����v �]&L�/�0�LH���C���Tv�$�B�����*4`>�+���>��.��1P֣X��w=,�͵m}l�ܮ�D�n&��m��ԘD��^�5Ęy��l�+���eQ�\½ڥkŕ-�c�Ǎ!<�Iew,���\�=�+3!�!Ԋxs�w������`,�$��C�1M��
��9�[h몰^Nٔ�u؎�\�ӏ^�Ij�]�$zx��`dD�BQz��3iz��'��ց^�A\�26e��N�o\Y��3G6	��~<7o�~8�-�ݵ-��n���a�Ȯ�[v vgl���CxI���5d�����n��x-I3l�����(f^F̏/;P�������6�H_b���=�������¿�;�����o�C�g�B�*��>A�3K �����Pv>��$l��4O��!���%�tM����+�R�d̾�a"��-�gv}�G-������.��.�HÑ�����)د]��̇���!,�$[�x�w�ڙ�q򚝙3x��=���F��P�o"��
B-��d�ke���z�����ك���^\��U�*K��B��t��|ź��n�q���\����z2Xp	�U��{1�]?L	J��a�yq�����)����0����N��i�hأ��52�%�z,��4���K傯��G�g������@)�vw��ٛ[�mv���C�4c��)�1,P�~6.�֭{g�ITa�>��zs6���n�����<��(Lf/C��Oȿ;�u�H�4Q��ϵ��p���)�T���vZի�.�?>{���;^���9�oI�I�����F�M���z,硦�7D$�kq��;S�sP�4!P�N'�?����^��ܶ��o�Z}�~�u����)H"�*�eɐ�Y�5�F����<jo
q��ˮ���em
��|��f3�r�w�"�ۗ�{.���C��6G��v����;�wh���YR����Ĵ�x�s*t���Z�B�*�Y��cP�fL$�K�߾�����1�>ӗ���O�O�7f�Kÿ7����z˒<<��\&�����'��z�P����kġc��Y~�x�s<~��-xn?yH�i�&��3����B�����1z~� �xsk8Э���g����Kb�S��W�7�#�}~Ϫdd)HU�
���^D;E�J�����V��S��-H��:�a{`7L����>�3:����ھ����.>�����1weMהG�����h�,��]���.X��Jq��=4�8��k�A~�-@�� ���kKD��4�܎���?�4���猵��k?�*�J��>�G��x�H៳�V��n�
�u=~ᓝj@��5J�'�m)�����{ʡ�9��;ո�b�6@%�7c�$��ε��+מ�k5�<��)��GV�' �����s����@�nN]w,�{��g6���]N����:�iT�P}#X���T��s�X^�U)5��b��3@�MFo��cw§�\Qy������g�oE���u����� 38�^��̹8�؛[6��V�n�Y���XUJ:�sF,��٬ﳾV~�t=�[Ɓr]��n�<��=�A}��Ӭ\_��&C�i�w�
:g�7q�t��G�8�G]xw���LΤ[�P=��c��w��[����+%�xԋ�oEw��R,Zb%�,�H�������~H�_�Ϸ3%o}����z�\���
�IM
�V�{�ʍ�l�I���h~|�!ҞT�J=�9Cv=�:yͭT)d�0�9Qm���,��جk"'�gD{=�x�ΞDg�<����^�l�<æ%˼'�L���)���:���M�{U�Ҷ
�[A�b����w������0+Xb�=><9�d�%�7{4" ֚|��� ���?�tWP�v�hW�9ن���!�Z��g�'6Q�����Ge���o��5y�����CLSs�B�x��{��c�X�8��I�x!����}�ĺn�}ծ��z�N���Q��A�l�	��2�r��N �+�C	O�:ڵ$3�6�C=35ۙ�κ��F�/K�~��7���߸�,-ts4�XJ~@o��]�(Pԧ ��s���mm9Y=(F<TC_vrD1�(��B�����r���"Ts	[Q:Ȳ콮x뱊��v�t0��OSO"���<1�����2}T��zq퉵[�#9��w�'�	�Onپ�N�`i���"�Q��64s�-�HS�E��6d�mٮj��"&.o�=oXnJ�k��xD�θ�i��<��M}f�3;fܹ��vE)%w���[��+�v㓥���F�(�٘X�Qs�GfhrɽG��!����Yg���I���8�ԝ^�mS�櫥]��lO6M{�Ns9���4��bG�e%��}�~*k�T��oC�ǡ���;���yw�HA�������=ӈ��F�L��P�C�O�=g��x�4���A}/��!��u:=ޙ��)���6���3���p�Q�����G��z�ޥ����oMB��=W�[q�?�B9��;��zݎ��G�T6��5��J�쑫oX<�	`k�w$Z��EMH���E�nI�Z�v�&��"���R���;��D�����������1E�Ci�a�[�'ϜD��-�	�5�B��G2�r��-��,��Sս[�S[;_�Ql}A@��~��{dG���Q�4�F���J#L�����#�֤���0G��z0��[���+��(U% ���}��cC�W\ǅ9�Rׂ�Tٽm0�7�ݽU���ķ?�^�G��#~X�P�9�I���A1�),#:�|ɦۮ�j,�36�Fԣ�Ct�&�}\�K�8�Ӧ
�E�3���Q{K��#����\ekq��T�<U�n���,���bN�հ#��|����}b��YPX��9����Z���8�H����ț��N��JH�*�T����F�Ѭ�"d�/�x�&5��	��>�h��$^���~�|�|�d�MB�Ӧڒ��-hz![��aCo8u�gK����d.g�I����e##������eR:�3{,\���޻��?����V#��F��@wt&�h���A~:i�zQV�_VԢ0�׺{�|����(��v_�Q����!�32�>��>�Ԥ��apXF���l��ضD{�M�BdK)�\���k�Q��Q��,�5O����
��tNer��_����b�~�"qx�|`��<��^:���:����I��C�c���3�+��9,f�����e�ܡ�7�&Щ''k��셛{����o�Wz�'#��)�u�4��{�>�
��-�i��-"���U�s��?`�x8��&l��V����,�,wv�<lJ�1�C���������|��僫��u�>ii&v����z���M]u	͂�Q�Q��x�J��ib%�����Wrv���e*��!��yuC��K�]�ʨWd�49v��^�	�:;�C�9�zȣᓹ!^:喨�F��KP(!m������ϛ�8����UU�rj3��Swthct�(��'X{ǱJi>S�'�O��Uȯ��!ڨX���ً�ߗY�mR��1a����)U��&���-͋��Lu�ٗ��1.�����?A �M8u���en`���kt�����ޡ�9lB�>�B.�^f���T����Ok�}�<�<2I�����n<}��in�sr���������yݼ�����.��P2�˨-��	�i�d���)�d��)X�~̌nl�<'��z�@ȕ4�:ɑ#��WV;{�(��Ű�q�][�LKߺ"K�H� eu��X���;^a�'	>��c�8F>�H�`C2�p5�A���H���ό'�Y>t�q q�����+Z�"�TF��K��1�P�UǙ�ͳWT/ ����!���Q�<r�=�M���<�V�v��\��-?%<uuc����9���pOn\��O�/���;"s�'[`�!���
<5@G؞�nm��#ݟ9��9uJݘ3'��6`k(t�Ѯ��}D�Z���(�W��_�/J���ޘ�b�M�Frp�|&!�f���0;�
b�}+�T�z*Ͳ%��i�_���y�lI��U%dm��w]����9����;�zm��]>Q��=|�^�O����������_�qF,U�)]��-��F�Ż$q� �X�3ފ���۝$n�HL3�gC��:���T0/lY�#L)�����335X��3P]WP�����=�op펃E,Bbc�ەX�a��
��f��X��p݀���p˩�eװE."[[�yǻ��욲��<������r֋�aN�M�����݋�!$�\,���[���Z�;{{'h��:ښ��W�W7ÙZ<F9}[F�}P�kF��!�>��q�����XiD!���{}�?`���f��t쇲
+���)�F���F�u�ǎ����acv������@��zn:S���
���f&��nbk#w3~��}�OdƉ�F����֕쭎L���,Q�y�ӂ�ya'���X�,jԝ�Q�M�T�Aa������9�E�w\��V��X�����9s�q��~rA�������e����m���x���P[�8t�p�ΌqgL)XV�N�L͚���}}���������Ö,��(�A	6�ƋtU�����+��Y�C��]Ǔ��:URy��ѧX�*�9hB�=��@��́�)���-�umR�A	�m¹uo+̾�����>j�č�U���jѸ��E���d�o]�YS����͏i��{&7w.��2��sfmD�;�w��V�0Eh��U^�R���vN��c3]Aox�΃Kݥ�7��7.o/�Ʒ<9r�]# B��;�1����6��~��7�s�D��9[fk�
w)X��%v��v�{�%�����0�ih`�p�V����$z b�_��4k���/yf+��Gd�2w�PA#��u�MͱupZ�uZ�o�:W�0e9,bY���8U��1@���Wx��AgX�Ӑ�KS7�Y}�i�K���[,,�ƞۋ�˷7۶�Z����BW$8��u�s���߻(��4rkg��<N�p��Nҥ���9�����'KrSV��7�ww�J���E����+�������~���p�����Gg�ǯ��,^��N�_Y;�I�5�V k���t����+K�t�Ny�N;�r�nF�_ ׷�Yx��xT����?z�9��j��C@nZ7Α�;w�m^Ca��+���Y� �Ng���}�N�Sa���3���1Wr2��B7C���!/��wo�{�<q���"������aܙYm����B�7�9�Ft�	V������87W�i̴&�����2oDwR
̮=�xy�Gt�mt~��`�7=P �7�Gx�'v�U|s-޴�R�z��	k�B���A2X�Ki��1N�])H��%���_ti�Y���*�6\YX�T�]�W�WT�bb����Wv7Q����T�@���q-r�yt��Sj�xN�*�Tu2���˨���'&u��W)�G�����v��b�]����2v)tx,>��|s�ҫ����7�w��3>b�h�%,Ga
�82A�z���\�d�Q-a�T*N��a97]���C0�0���_� cQ[�4���׏<x��x��Ǯa	$	l)1��HY��scL�"d�ʨ���I"[z���x���o^<x�뉐$I'j�1��S-'���\a(o�M>:z�<x�㷯<x����ſ^��l�F�'����>��$��cO��|q�<x��Ǐ=p�22B)�EԨ(njH��hMkp��卲F��o���A���׻���]��t��^�-�\�kDd_5ֺ`I��͍�*��&*�l�}7o�ܣ[�5���}wd�5�x�~s��DZ��}{��F��d fr;����!�6�L'D�3!��Xm8F	D��Z�;��t��0�[%ˏx�BG����;��Y��2K�Xu�u۩�,Y9���Xz�ӱ�Hk]�x,���q(-�m���Z0�&�m���!XpL0��B[x�$|�JÇeae��$`�& xI%�&�%O���.	q	�eԹ�!_�?���������^�:�X����'�촿Ak���rv�`�YKN�pw4a@�S�����g�U83��py���]�D\�����7]�.f'�o�_�(r�E��4_3�-G�/CUȆ.���eΧM��ss� ��˵[��ʀ�dJ\*�X�n������X�V��c�3Z�'��Q�p!!��u��8��p�j�'J<�s�z�\�[3�Sq;%�ݫ%��-l�(EþA��,a���]it�2hΪ����a��0���k�;X�N���(6�X��W�r��	RIVMTs���)��x�9���]ד%��H)���"G{ ��6���S�Ǩ^�`�#�<���R��6ɒx�0����Ϸ�vF�E�l�YX2H�3�bF\���Qݭ�dwI�c]Ya��+ѧ��SK�n \wu��
9���o/\�gz7���N�;�'�}F�����uƿO��e��h�ޚ��,5��F6�yMH����l�Y�Y]`p����#G|�vz΀��X0緍EpX���kMFӼ��!R��)�j�uc��u��!�%���^�,�V5&�^���d��doN�^2���>"�����zZ�E��ۊ��z������y�o7���9�V�����;��]��7ң܈��b�n���hxOl%SQ%�k&����&
�!�v��Y�/�t�{�X�͡�"[G�E�]�Yo+&'���#��,9c�Q��s�w="�����m���.�����Q��`8s>]/;�^�)�p��iԌ���ol��g?��;*AM�$��fl��q��t���U��sPn�O�̞��om���z2�%YN��i:I	d�tI�q�/�-�΁�D�G�%tf��Z�N	�5�-�N_��Mo<�����/s�G�p_o�r�Ǯ[�S�}�y�]b��緹0!�bV#g����9�$�fX���^����O��}��i̛�<,X���Y�&�l�2��)Jx�i�Eeȥ-��:`Z9s�W>��SV����l/�y��O��,��F�K9�Vz\­b0��*�]f�̡z�꫗U�t��y��<���`\����lۜ�mX/5� ��"Wɒ10k�U��u�Rs=ҳ�jP����'.���ͽ���0�Nk���t��v�`�6�&��b�r�Y��ٌj�cR|׼�>|�y���@��+���<ެ%*򒪝��O���s�8�XL:��ظ:�o�9=�7݈�=5�{pT�4�#c�
��y/>��[�\
��s�C�g�t,�\�b��ɳc��'��<���#��{����#�K�ª���� K���}}
�6W}�Z��/)M_��k��+�m�a�����Z��n��{��c1F;���>]s]�9�ks'm�Vl[�wd��JB�Q�u�.0���b#�7��ݫ�T��ONշ�?NfJ������'�*K�1y���;�����x���L���j�l�zcx+��r��7�E���d��g6��>���`��r+FK��M���bD����'�m�v�؏�J[��x��h*3R�Z���m�4%)��lЋFE�z�������u�/��/�����N��z�<bu��J�7��O7Ң�s��5b,�aUd������[/��8�����gg�	(�\�����Y�5&�-n�?6�ev�;x4I�O�8�v{%^_)e�"�Y���t�Ү���W��!1q���xxxxy��q��m��E��>��m���l)`��4.jz(^F�V3�e�e��:��Ȏ���x�2�Ȯ�{���������teM �#��1�ؾ����%�bH�婛'4%R��_�|�O���<�=~ {����C�S{*��l=벁����d�7�j��T�����fO�F��0��6�
����XzU��C�F*���*��@��v�y�M��]v�w|�^3A�S}p�,57���(Ñ���E,tz��r��(�m��a���=�����oͧ����l�ݐ�	�W��7�JOθ�Ge�^]fe^U��M�N#F���l�n�,0l��҅��+�_�ow�%���y���ec�����gG9���=���<�!��.�~�^1O��;.fVG��֞ؗ��{�^k�1IwJ�p gms+6̎�&�crbn�k*r{�*��ŽEN�t�Ր���<tr�l�WMvN�������݄U�j�f�^��V�gh���4�W�k��F :�)���5�&	-K�׶%��㩜ӵq�cIoeK�+r�ӭ	�6]����5+��D�h�i�Z80�\�.��2�+��xxU��h�*|���6����J�U�A���_ѓ�e]x?B�9&��b��JU{L�g��k�����k�Q�sZ�����c;�7�R��h7j��������N�m�ӵ|!᜶Q��vNx��H��t��-۫�Z���G~�=�|�+�Np�^Z�xʮ��ُ� D�X�$q���꺣�U�⺍z�C�{^Զ�O�\ώ�*��@R�o�4/���e�i�݊��@@D����6��&��T���v��^½~I��h;��t[�Cz��F����/*Zz����w�erg�ܝ��o�~�
PL,��\"���R:Z�ᗈ��a�����n�����m��� �����ǭ��\��s�E����;���YC����x� �?1���~���FD�@ǽ�p�Vr��\�F�sTU;��+98�=���SOj���/����`�<)y��[���	l�{��״�o�Y�۝XzK��~-�`�ۓv	���G��A��GH}0����{뽋�ߘY�h��x.J��v���6���z���<��Yt"��>�и��yAww!�t<�=��sS�=�B���\�C�xU^L߼��X�c�1�QϜ�/��:����k��>�O���dt䋠���!_��{.���a��{l���zG^��+�d�#cl5S��p��^���}>�)��<라U���}@j���ܥ|�qsn���G�ڨ�ζ{$�*/' K���w3�����${�4�q�վΕ�ǞEK�w�S��؃<Y$��E�Me��nXV�tw=���}]����7k���}�^Yљ\�e��Y�k�8�,D&��0��� r2"�M�R��i����R�9jqU�h[/�	Ǜ7��7k��{2jjp�u�'�8ǜj��6��Y�K��{��&.�:��� �&��3P�1����ZF���w�b�w'�.9��'��E��;�U���^�ndl3��tf��ꎋ�zt>��oR4qn�oG�w�����$�x8*5��o����R��=G�
��^}N��s�y��+&���d_U�n���&�ڷ��4�[�;���]6"�c��k��HE���a�K�$Ց�QKkk��qV�2��IۭKT�v�AR�߱�e�u��cq�ξ�D�%r�tj�W�
���u^P�g{,�_��X��T�W��ꋃѶWN��v���䘮��1k�|��W���uP�2F7��v��Bs��[�Z�3��5\c#\[��]��,�ܖ3YШdӞ�Z�ٞ��0Rb���l/��z�ɖ#iUk�^�����^�������m䊚sV�ujɹg`L�Y�\��0���qKc5�װ����ӣ�J��:��s��:�>ǏH��q�\��[��є M�	s�do�
��c�q�W���� \�:X��
/�.��+�}n>�C��Nż�Έ��������?2f��&���I�1}G8ՁG�C{r�VH�x.+��뎾�Z��gv�Dj�w���ȴs{�!�;��J30Kh�A�oc�^��_�sר�qU�#^+ru\L@���%��v��q���[�����y����~�x�"��ճ#�ay8dƬ�L����JA�웾�p� sm�5�M��C�������y.�#X�{"ɞ�2�PW؞J�*�{#c/���]d\��1R��!�{~��JKZ�jR�&��XW:w1�]k����F����1��y�s���Oy��{�ݼ~&�e?�b�e-��`G G1wd���c�ы7����`[��n5�	�#���Z;��	�;P8	�ͣ��wA�S�F��+*kmJ�Ъ��R�"���1�+՚��wLzw�p��$秸Y�����Mo^�6�v{%��*��<4"�+-��?SD��5���78��n����Ʊ�)�r�w+�?$�E\�������=S����EA��<od�郛�.��N�:�k��q�3��#�&=7��	��Y������%]�ۘ;����fڹe`k�� ]u��[��%��.�
�=u&Ӎ\֔���)��>�ʷ���SŬv=.��N^|'C+sK���[����O��\�� ���U���`�]� z�Z	�;�`s�z��Q�Z Y���OW��*�x���1�Mn�5��B�ʬ��m�׼��Oo�a�{
�i�N1���V��ZZ\C��xz;`r��V�Vj%���v7v�K{��S[Y;�7G`/��	_[���픺V+^QYs]g5Ah9N�N�cT�;��q�ؤ��q!��_�<<<<<<&��-O��ܲ�9�|��Xq[Y��t�c^�9���-�K����!7R�����vU-?������*B�;�E�6�$���כ�g:���o+��{w��s�uyu�lǍ��Cl����u���e���¬�ent�A��rujW�[5�Gl�'��[���F�z�&T���z�mDV��wO��Vg^k��������4��͏0]�%.��MƟsq�͑
��Vc�_�6���o%4���芒����"���0	��Bj��6M�6�J�%#=�\.�۷���OplՔ8�uA����g"�Ƀ�_��$R�C@�2��ha�F�w�H��Է|�O�����u:_n�fIѵ����0 |���X�8���;չ.��ގ��:���v���1I@����?��p�_|����u��.*9�3���Ҽ��u��$}Zy�ܻXb�fffǭ��xB��ռ3@����W�b�k���aX�D�ئi^Fv�H+�y[�3��M�x]������>[N�$��ì��I�yf�^d���N���Պ3��w����LwI��&.�knV�ou�t�2������'t�R�a˻��H��*z�c�1�������w�j�<����<�񴶷8)J��%�=ٶ�����lhE^�������6�8Ⱥ��R��ۧ\�}�^!����3��u�K9n��^�����㵑�4�g�q�/�}�)���:Q���P�����,LȈ��x��.�}x�{M�7M;��9
8	4�u�+�ʸۗpjǵF�1{J���f��[f8Ӈ�L���)Lk�Q��ء�Su�/�
E�x8�Z�sn�ֳz�6��Aȡِ�V}����KɑE8�6xL�oh�zL;�j����l����M���x��QS]�[�\o��������8c��ͼ:R��f����L�P�|��� ��>��#w���#IwH;Χ��o�\�Wr�/@QY�Q��Eq�n���HiG�L(�v��Ǖ[�j�eMŻÛ ӹ����+ުr�����W�CvԈ�R,ʗ�24�����$m�+Q�]F�v_ 6��>��mL��88������UN�����J7k;���}�k��+�F�M�~����gR�)b���Ĵp�Z�Ki�֪�V�j8s���Ƙ�}�.4�a��/��(�*-�d�dJS!R��}�2*x)ᝒ�D���*�um>\��2j�����B�b��
wxN�ީ8<W�&=��aD�ܳ{ң5w:�Q��w��]�(��mu��6�Ћ ���`yݐ�t�o*![����+�w����@��MA�U䝒������������5��$�zLZ~��\�dj���9�v�к<D^��H�4�J�77����]\��
έ��z�j�m�� #
�pI����vs����/[4�D�٥+x7I�D)�71eN�6lٽ�����f�Z>�%ƭ���w�.Is:��e�\�PU!��o�!NY�U���� ���D��J���.E����L}�P)�{oK��Ԧhu�j�HG�3�VJ����v6�%��@��=�e�oP�3@q+��+J�[�M�*����ԥ��9G��//K`��y��U{��ed|�n�Ԗ�V��ғ�e\��I�-��o��^a�A�p<��.�170���J1Z�cF���Ibn��ِ���|h����z�YFViw[%��FhZuq^2ӔA���0X��������0�y�d|g����t,,�s5�L�Z�ccG�fatLh��8�P����>�<?�-8�s"�BD��Y{S�;Ł0e�lf��1�UgbR�ݷ'^-u���32la#If0�W�΋Y�b��GU��7�Cٲc��#(Y�t�a<kgu5�5:�4��x�A3pNk0�I������b�{��Μ��|�����B����N���F����YȢ���z�P�/c	�	�v���ū/q����im�*/3f@6wn��9�
2��k�k�/�����E�;]��T�u�Fl�a���n�ּ��Gj�R�5�w��X�)cM{�vdɽz{!�6d�Ɗ� s�򓝫�N^�)eOz�����{!��e��5&;�q${xA�7V�mww���Ls-��V-�{0S��T5���;��;�����M���>��}�w<'��͘���A8}�.%Z�f��U�t�EIh���0c�2V�`���f�d�͗����ys4��> ��frL-Uk�bR�$�ۖ��a�V��ٴzBP9�E��5�>ZT�--J"�Q۷b�����9��
79}z��D��vr:&{��:~~>��7�+W`/�X����B��h2��>���tk;�1�ʘ`1���}��t��I��vDw5񮙐�����<��NsY}�^��k�yQ! wM:m��n<z���o^<x���\��*()4X�h����F��]-�ݾo���\q�Ǐ;z��Ǯ$N�j �2���������m�=m��8�Ǐ;z��Ǯw���߫�O;��cF�H� I2-1�����x���o^<x�̌���!�5���H�b��]۶����^O�Qi0%F�\�Z"�P%{�'����Y����~uՒ��QX�^p�cnk����\�-�������1N�濟:��+�k�n��Cn�\"�ni9�wv���.t�<����һ��H-@,�A0JE��ފ�莊��wW#:�:ZenՇ4�5n�QM�x�7��xF��I۝�`��fZ{`vh�(���m`=�������Vo'>�e���Q�߀�C�c]�z4s:>즐ɂ���aH*Ŵ�F.�\�&o67�ۊ���3q��t�y����iY5�х*�Q�T���������_1J6��7��>{�A.tI��ng��AY�|SL�Zc��7_`/���՞��T��=!D��F��,�iL��'0��5c�Os��`��:ы=>����ʻ�;ـ��gilJ�j��^�����O�y��2m�O_���(R�
�k�p�
EJ����U����y�,���䷽�Sv���7.�}�g���-�"��@%�e{yr4�c]��Z�F�Wg	���ʼ-#J�K��ھ���<7���޽U0�EqY�H[���;� !�1�}�V�W��0|������F�%L-�AȢ�4DWr%v����%�N�x*�#��t�Ӕv�{�t��unCC[�Z��Q#Y.ln���8�YܶLƹ���͐����S�)ߢ"�{q�s{�8k�F�\XN�G�T1ƽ���ٓh@��\Gi��	��kRc�W��{}z9�ǃ;:լ�'F�gm��B{��$�&�h���~���������}+�4q8�����uţ6y+��B�͒���/��C�γw/��h������l�A�M��_zV��f��	U��G���z�()<O��[w��3:\��`3����b���2)MQ;3�'���v�wg��I��G���0��zb16Г�%������:�l��;=�!�J���y����Jb�̽ײ����"+���VL���J�g,Uxa��ň��zͰ��>��݆��^�x����G/�0o�����%��W@c+7��_|[�n��EU#��@2���{/a5�;yn�B���᜾mur��[��5@����w����;R�54u�/��x�p�{b�H�4;�]�*���Ѭ��:9��QM2:��2wf��y⮖��d�_,t����?5�e�a�R�Sً���oq���8���w�#������ր��=�X�Nі�6Т��)J�H��S�����s�K��ۺ��[򿾝���Y�纜�l>��`�Ĩ&T�/�v]���o��N,F❻�q�G�o7{'I5RQ���-�������������6_˾�i*�8t�Fֵ��ÅQI���am��xC��3�v�:8�4GZsm_{.���ˏX[3ػ%���aǘu�z�d�)Y�#�+�������z�ni̊
\�ܭ����g�n��FD.���TU���:����N��Avʣ�]�z������t���O�W��,\y������s���x��I���
:C�\W!�]E���!�׷���ռ&`�^pQ���hޔ��6��=�q���<�U��&n��Ǟ���Y��s�1�a�][,(4Wz੺�^�Q�X�uGv��@v�ir
��1sl޼���kN�2a0#z)]��+9T�,��u]��Dt\�:�\��K�@]�<g�>|�:��Ũ�R��;��.Oy��|��·����@oK=��������m�T���eV]{{ӊ{1��T!�r�ӓq*C��<�x��xοk6�e��w�A��;�B�Ќt󃃴�fZS�ff[�CӰ {����}f�) :ު��&��;7IT�gW.�qN� �o��n��.F��qˬ���*e<��/I���:a'��f�M�w�l[:.�W�G߼<<<<<=&}:1��aC(2����
0�R� �����g������C��1�����m�����]�h����_TaJ�`��-=o�ԽS�zKOUV�"��%�G��)w�x��2�4�sX�+�uM{0��\���Y�Sݱ�m �t�FjI�ӭ�)g�-��h�^W^��Ⱥ����s�:=���2*v����+ ���_�H�����s�>XSE�~���]���;�e��&��8^j�#��'�cr�j�z4ĿwsM�8�4��`���k o�+é�}@oX�o�5ukL}?��f�FF&*+}�8'Ls=�ٌ78��g�6�m�i���ރ��k��W[����oS�5ڍmy{�N�Ksʁ�!z�F�HܷSّ���+�!1��`^��Λ����Ǿ�]��KZ9�dl��\�c�p!��k�t�#Ϻ�(���1}v&Y�QN/�i��q0����z*3�;'��0UL������f$��<v��fA��![y��-��9�Qé�F�J��P��Y�k�W�IÞSʍ���Ǘ������ e�ˑ�O~��������-�Ra�ng�C6F(��_�ok�\�� 1s/uyu�L7���G3���sz�k���B1�Z�=cdV�W����i 5w�X"�BQu��X�ۆ�[�T��`��d޾�T���MV��V��i�6�d�S>[&���鹃݆ʏ0���g�f��+�GkyM�Mܘ��s`��)�~[*�;��2I��߫f�o+g^|F(p�7�>�����=�ln�1̹f��c�u��7Cz�������TG��ٜ���Tܺ�ăt�\�Ӹ�B�<��^ޓ>��s�_݂z}��Φ���,��-Q��WO^�O����=�W��V����t���0Cx�s�fD�N�b��߮4PZ	wJE!���+�lA��'����d�н�<�>����s�!��\2r�n�d4��见톡�^!(w&���N#y�5���4(|_a�l��h܀�&�S/7��І�7���{��̼�vo�5�}#e�����g;����k�Vw3�H�R��vJ1�F�JB�=�MK@ͱ��۵FbjB�����w+�2�Ն�X��h�t��)Y΃��y���C�����9�e�$�w�R�dq8��8�i�f~��{��ǫ�--3Բd�7�V��B��b*��)GV��Tәl����W[��b@c�SY���ew�����`�߱�#:>��@%e>U�j�y�f05ʧ���4�s�����V���#��v)��/�Q�٩�y�z����]����l���Q\Zl��_#�L�G4���5�F��٬ѝK�c����ί7G��S� �ճ|�^�5qװ��x��ɮ�}�pgl�s�BC�z����f<ņ��jow�ɨ?�;�����K*��	�M(ㅉ����&�����|�9�~�_�~W�9���FY�h6`۶e����k�z_�O��9�wN_��3䒨�O옹�[#|�u���j�F�UfWY�R ���N��cn+���㙺m��v�t��|S��5[�/���vi�N~oR>�%�մt%Ιsn�ɍfQ�Dj �;p���E�aGQ���oLHi��A�;	"�"��C�l����)ku:�$�j�oc�^�ad߂�����z�a8b��(c�U��67I@�B�hgYr2�Ye��1�j��{W�ʚ�̽�R�ٖ�#+lgjv-5���~�y�uo����X�n��Ѽ�]ݮ�<��a",ύͥ���������GQ��
�E璬��������)�n���T�l�r*70�gh?H�+#!����t��$�v����*j�����ڃ��S�%�^���^Q�tS��%�py'T�衁��5j���3\X��0YK�z�X�AO��E��y�zԋ��D����цЁ�����MP+}���-Q��mF�܂�҂�q�v����������)��&+E#]u����`�7"�+�#7�>���#Ma�4
R�t<E=ۛ��Ҟw��l����r�0ƹuR!�����g��?эa���mo� ���>���zN��]9��K��;�e{͹̲9gn�>On��7�=xu��מ��WQ�vm׀��� � ^q�ѝ��2���ӓ�uA�(l�=\�.������7��O�?��n�}�1O"{��ڶ�%�γ��!2���H��F����8�q?VM��h��52���:��d�A�3L��n]s�23Ϻ�b���є���S���xxxxxxU'��A�_d���!��P2���gX�h.����k�B�.S��ڪV�y�coR1__lV��կ\Q�K�v>�<f6N���[����Oݹ+w����&g��MV��*��b-��䨩���_<Һ:�x�t��z7bA�����)�N��g�uU��e��b%R�Y]b�ז]��m�o�o����@Y�ǫRՃ�zLoT^n^N�M�u��6�] ���7���8s`�g]�6&�E*u	D���k�vKQ �2�����*�v����I=�A�@�c�^ر[�������nܧy�NK��Ԁ��1#A=��p���h���w�=	|�#166�j�SͿ��g� 8OWa�A���m{�j]�Z�V�.ys��Z1�j�\0��G�/Ӌ�QSt�����H�ñ�I�z����VCE�M�"�]���Y�&`��rQ���U��L[� ��$��;n��Y����ctۗ�ٝ;[M�V��a5���\x��6�$at7h&�i��ך��N@���t4��-�w~�@�~?���ܮ��/���I����F�e���y����ߧʒ����P$�k��b�y�I�Ys5{������#.�$U��`ǧ��% W6��^�fj�6
k���c�7,�Ϳs�E%�8�a+�:�����bK1nS��c��(ν�I��H���װ�^�)sA�S{�>Y��I<�-���~��wm�ʄ"�YmP�_y�Fi~�ByL{}Oz�Ժ}��d�W��iMA�4����^�Ck�aj�ݑ�McdV��W��<�4�y.�=S�љ��]�>ۥ�Ϻ��òV���U鞊�m'�|Q�֚���*{n�P^��ED`��a� �m�/����~�~'��U5`��.���n�Q{�A=�C�u+���WF�S�,|(9~��_�ǆ{gʩ
�wk����E����Ǧ�ס�����5 ��8�t�yN�̪�۱^�A�U9�$�ۨ�I���:8��#ۛ.eQ�=;C������ێ�ᶁsN<�#U-ub�.A]9$r��ʇ)�GǬli�ىKT��s�0��g�D�pL/KY��έi��2����IG|�����������P����(6����8���t���e�KyJ�-�$�Ta�,���t������"?�4>�qb�y�iP��Z7�������8��	SD�{�����9��2�	F�H�ϡD,��SS�..Y�v^���Z�4���'�(Y��M����~�<�觏{a�P�/$��������S�I;t���`��=8;]7��<
����sYЉd*�9�����S�e4M�hF;����8à��E�m*T��^����Gx:�PU�~�ڪ&�8s�ލ��9�վgg}L+W�\{5��}������RQ�S�^�*әLӍ1W*�����Y���;��5Ҷ:9��&�����a����Y�Z��:�.�\��"D�p�⺢B�ʸ���䯕"��|�������;��\w{�ӵ�6?���	�p["5l��t���xP#j���9�s�>�d�r���X|�Wq�ga�.e�E���}ȼ^���l��f�Mm#�,u�	R�֦��D$�6��!���}�
��#���0.��6��!wLu�^�mv��O�8�ǆL;�1�(ǲweS|�d����+pTT��iΤc��0E146q��1���l�+ݕ��H����&�ء�V`+E�=u�V��GNԩ�2��s�@��˼'�9�Ok-J�����&/w�Á��u��ո�w��`U`mK�6��ub�d�c����M[�]��(<���Q緇A�p�ˮ�s�Y5�]��-��x���a�JU��͑;�'�'�=�Q��Κ�J�>._��ｫ�q1��C����zl��%���s�b�`[&9�y���o[�=���^;�|A�K'M���*��s,e��{�]�@��{)ɑ�ð��u�-5�α����ⶾ�o)d�Y�/����m��Y��ub�V�j��TƧ�ɠR%v�����q��m�w�晞���m~�=�m�ܾ���dy',�C'Y-w9M�g��of����0ؔ#^�z%a2���A�A�+mvhXA�:�n1غ]���g�)�
�u9�&��V��ɎJy�0�=���]�%s���谨�2��Q����23y���{�����F8�r�ϩ>�9��B�LK�{05���М��un=��d �i-Ew��[M/��3�Q�����3���/���VB\���7d��$H����Eϲ�d��y�{:#�9.Es(�yw&��;���)b�6����0�'�Xթ,��5�<ї���S�Y�szy�R�w��]}��w{��&��byZPD����ZD���/�ӮQ��5`�I��-���9Cw�������F�;1Ry{��v�s/�У6wT�����tF�=}����SҰ�Ubw�r�3lrM���
�#��묆�x�/�6l�r��|�
�!0!�;T�3�9�YY�<Qw,q��M�|/�1ݸ�����[C+�Q��%���I�{A�S)STs'vm��Ūwb��X�	�;M�$R3#Pm�[�K��@:rR����U
e��,�����[�>��9���ۇDNy������̰���kc`�����RU/�Y�]�Y���\�}�&A��,�#�H��@G�ՙ�༴����bn�b�ųt��[���/����ϵ�Xz3��yl	�ޡ������do��Avwrf��#(dL�q��Vcם��.j/���m�s:��0���p�wV��v�zz���7ujavA[�nL�v��Е�o5Fp�&n4���GFnt�ve���J���3�t+$���u��n�c5����Ip̾�Y3Q�E�DJX�(�M�;���������`���b5s��� $���	,jHj!E4ӷ��=q۷n�_�nߏX�!$$��%R��]t�͸�/+����P
��P���ii�=|m��ݻv��۷����dMBA�@<�Io<�dly�^s@Zi�������v���n޽qrvT)�_�ʼ��ק���#GFFIT!�
��m���v�۷o�]�z��WjI�U�UP�Q���KF�̔nE͹^�������˜)ں�����Uȹc��rط���t+���m��t����nh�iW+��u��Q�wW4��W;�r�wA_�/*(�מ�_�r�\������9�nt���9r��ήD���u�6��t��ſn�s];6��u�}}o����=ܘ��%�c�Ye �0
0�0Q0�x�8��G���o��e�ݶ��V:���pF����XVr+8�}+Q��ol���VL"�Q&����He��3�7MVZ��ְAR�&Ri��a6�`������Nh0�l�Ȁ�xHH2�y�,���?3��P��G4� �!� >H Xx�(�H�Ur���bzl�vo�2�ڵ�e�k�e��3m��5n�=#Mc�f����.�=�3s�>\_��:�3��[F0�zz����][�y��E{{MP)��X����}��g���wk�v�G��)y�_��t
~�Y�w���TA��9o%�Q5%8����T����>��R�/`�d#M�0(Ã�}.�+�}Y!�[�r����;�Ϫŉ��_]f��K>I$B]�?�����z����zB�[/�z�S_L��m̵��Wڊ��h��<�to�p�����1z-O�[]!G\6�cJ�ף^:�"k�s?X�>�����z^w"���[���N(W��!Ҩ��훎n����}Bk�8H������r�7�a���{'��CM�S���	6P6f�(٪py�!I6�$u���*l�����ix�Ts1��aR/�(iM[.!M�()W�m���d�!�Hp�j��uX�þג��R�a��"vZ���j����
06����/"�D�p�yv��uT2�����H�s����P�o����+�_<p̼3��i����(2����1i�g�lY�{e�寪LtY�jhһ�(��`�f��4�����C���dBtߦ�������V��V� c�ꡝ'����̡W���/=ӵ�F�]܊ڬT��VΥ�3��Ѝf�r#��8𡡟|3ǷN�y㑺�=פu*U��m���B�� �$�9�.�(|���m�A��ݬw�����ֆ�g\v��v�;Q��A\!?���F��Ģz�DV\����}Ux�׮�o\�Ѷ���>na��w6�[�/�Mɞy��]yߌ��{�F��� �8U}:�\Q�K��^Q����vg=�����B�-���ww�����]�!��{���}y�L��YV�z+�S�n��m�qZ�fѓ��U�VEK~�Hއ	�m�Rt�7l�d�rvtRL�2o��ߪ-L�|�����V���WBإ}��)k�+g��AV<��N:*����;[�ݜ�猬�0'���4ڱ��&+��Ļ�ڼ�a�n��Wד�p�W�z@Kn}�{Z��ox���L�(�0���{�nv*���_2;�\�=9��9Rk;�i�eΜ$�v{9z>>��c�b��böQCT H�$<�4��qn��c;�9���o7��� ��':���`��n!�h�^t��i�H^��n����}<#z���N�����Dz�����g!"4�_,�]�"U�{uԞ�{4wT��1�q�T���M��u��|	H�HK����kM���sH���j�ɖ{	�ꧪ.�{)vyW{s��x��t���g�񦳇��y�3�k��}[��$�TK��:
=r�0��#7���Ukt�o{������:@��6�2k�<��_D��y����ВMDfS�	�y�e����=�Z��<$RE����R����������ڎ�NNf+^����t��|KІV���8��k��,y�����s�ie�D�*x�~�5n����ƅ��=#��9:���������kc��&��YVm'��eAe����"��A!^�1w"��<�F�ְw��T��)Ёq�aը�ں:���Pjyڋ֩_s;s�{�ڧ(��D�WnpZgO+����{�n0O�LC���P�ĸv|34;��Y�we]6c3c� ZR�dY͜��3kAJ��f1$�Q�n�	��e0'X���4{�p��1��<���ޚ���|���^���v��g�%�oW�
�=��\���ݍ�n�I����o$0�(����T�CO���O���Sߜ�4��s�ŻU'4b�������9���JĮ��������0�D��]4�q�+.���u������2���Nzr�s��dv��f쎺K�]���C��<g�~b��oxM��L�-�>'�G)MsZ&�{��p���Ö�/V��4��h��6/E]=�v"Hsyq�E<�Y"j�~|�f}��-���� ǣP��)�ˊܼ�:7H�녩�vg�׉4If�����HښE����v��{�5�Ed�yq���ė��B�{�k�ڍ�*���yf�\�-(4��[ې�q͂�E�u���"���mz���)U�*�׹��\���Ϩ[el�hoB��SH�We�����b��;^v����B����!"���&��Wչy[f�o��7f�J�;!�	"�{�q��$�t�:���nN˺�&�W�OC3��}����d+��2�$���O]ɍڷ��Z��	�i�? x�����T��b����{�T.H�,Q�d�s����@�ۺ���J�C�d@�x�C9#:�%*򒪼�W�|W���6���i�;nl�m58� +�KJ�e�N+8D��e�����ǯ���"1�ɍ����5tC�e�����qh͞I48��sE�i�7jk�z��wGm�ɶdd����#��:����j���]_���u�J$.�j;�ys�D����_���WD�Y!�oT���Ϲu;�V�~��u�F��]Cu\Qy��|N�] �n4��y��r5s����x㡓
%DgLB�>guⴢf!O����>��y�	�+!a��`��9�	aܞ�e�t�}Y>m�u�g(��&��5u>�_NTUu����e@1֙�,�a����,l��ϯ��dfr�݌Dʆ���{ki���ѻ��&���%���O�����ZR�z����N����w�d��t���b�Z=�Zp�d+��N��{�����C��Sۋ��i�͘Ԥ�ӮK2��[���35���#R��ϯa��oCn�>b�y�S��lb���`��L��s�^��9�g��xxxxxxW���|�߷\f9�Rc���$��?NC8A�
���K�����#]c'g�/GI9������l5�����26)�rY�twn�Ry�LИ���z8I�!���������R6�R&	�l$u�ie��p榜ზ�WstWe3��ֻ��v��\B�P�Xt�=�MT6@U�(�i�G[�"�ߤ
uN����W���7�:INp˺�bWsC�29��pwn�j�2*���u*`Vh�G��l��7�=n�vNϦ����I����=�� QUO���][ �J ~$:jV�Vh{���|�]���׮5I_��:���8���^ߛ�[����ӽ��g�yM��"ا8Zqq��ZW�lZ��R���J6(�����6�&3��O�s������=|�k�^}](�\1u'����O_��,���/vn��H;�2�ج��9i�V`�ݾ�\�.ݤ^>�npW�(���H����۟�C(r��	�`L]b���͊�ͥ��xo�+�or�&;x���G(�U�rsXt�:�˕}H	; E�]w������o7�������,��*��ʐ�2�x���c}�X`��2"1H�;>}ު�Jin�T��ߣ�v��T����]GwjC�-����{��3.4'��.a[��hu)y��������gE�3%e\�z���(>����KE�: -wm~Ʌf��4Zn��ɺ�-�*���\t��6笫P����볞�CU����c� �
�i!4���}��vz�u�ӝ��/귩ǟZ��i�g6�r��H�����F��z����}%"0��r�V���bmV�{o9���귳A�F��Q�R�*��]PS掲n���e+"z5�C�M/�j�Nn�:+k�~L�zY���=��F�.�.T�*rn%�B��sW��Ϧ��E�B�]�W���Ǧ�?�a���,�~2���V�7VoM>�1|���
��h�Ъ3���&u7������\U��`�Rh-d�8��d�����%����2I�w��ʸ/Fp��+_57\�Cu��dK��< �ꝤxUd!>[wdⷝӡ
�*lt��]�����:tNnnU�⽾���d�Y�E�2�ݦ��{"x�83������������B��q�}�\\j��5넕�;�K�K<���Q���vJW�5\;3+�f.�2t��5�׬uAL9{6%u�_|J��?�O��/�
���&$�C�<�;��넀��,����� �)��[<���u��p[��f�:npgV���n�� 5y�������� ��j5��<���Q��e�gL�ݟT���;Υ?���<6X,�>�����=qc�����v��۝9��=M{�DO*�q��fz��2�\/#��;')c��Q����2�C��"4ϴ����J�tyl߶�_Cs8e���{��{�wkS����qqtNR��m���{�g(otn��Z������m�J��8�g��6����2�T'47��hqj��9���E��U��B�ڷ�v�/��:�q��FƍqWO��o�F�f��5l/�+���N�g��5�<�v�f��yj����/V�Z�OXJ-�Ć���)�w����9�U�^�wq,提�,��9Y���7��+9磸v
m��fJ��[��cP��컃v�MBP����+]^3�{�#� n���Lg���~?��
�csZS�sr)jՈF�5D���`���bb9]t�G��=%"&��]�3�)�F�bKoM�W�0���{��y�זg�����E�`XJ�C��ɻw��+(�n��-��T��W[�7}$�5�4�a�
���ѓF�$�}ա��>��s�m�P�+�e*&�=r���\���A�꣝몐͉�w���}YOʬ��1��З�IT�+g��gw+�׭mӍ#���ߦ����+0/��'��ic�
�iغ���a�xovﻈ�6�>�K]:�k85�H��h�,���MF�Vfs�GWt����u������:c�H)�?�gV��mK��ń�Pܭx�d�y���Y�~����[��a���θ>���S�3)�x:K���v{"��;X%E�K9���k��W�Ϡ�n+��z�:�*����9��9n��1�Y��:��M�]+��x$�Gzs���3�E���D7WWa�G��f�ZUg)��KƲ�m�1l�w��D��B6v\7i�(F^�WN�%ې"�˨�s+RniRm�ء��o7���#y��ۦ���D�T�guԷ�J���v`Ţ�]��KL�zכ��*P�`�C��ƨ�p_�h�zU-��W�o�l֎@h�UqU7x:r��EGD�g�z[!�dny<{�l	S���n"����=1n�]��s{�k�A�T;f����:�z���foH��:k��Y���n�a���ѩ��ф�u�h���o�Lu��([V�'Wk���i�����OR�
2��[�S�\l�=�tdlS􌖽=�A�*�i؞���d�`Ü��U���Ug�:��p�ޣh�]�ͽk7o6�S�?��'Gm=��p�8�YA�%�طn�q
�J
U�O�tE�ԭ���C3�9k2oha߶��"��V�X,Od���J����#���Ŭ�_�W	}Y��dv�[�3㶽��u5m ר(70�
���x�?�Ú�J=��6��)Y���ݸ��k���7*�º�g�����-au��;	(t���!�R8�hڹ�N���d���b��g֬�=!e�(�r� ���ci�V�(������n���dC��n�;�^�P����G�<M�q�]�x��2��
3aE��ފ�o(m�諲�t�nʤ���ZѝݏQ5-�UN8>�����9�����kuԿ. ��Փ���'e�ڊ��]�CBm������C�k�n:�#ۇ!�4}<)���Q̽�M�MV����E����5��I�fw��T�^uN��ZV ,L��o�E�"k�!���2s�̩{pP�$,����7܄��v�t�܍x[�I�\q��X11&{Oq����Ӆ��o���en�d�0�	����1��U��z��z;kz������`;'�#:D��f�|k��e�a��y)��^�`ŉ��{M�L�.�ʋ�uu���������GiX_�_�$$D:&�b�K����0��xz��^�&��yʬ�:�~3�7qz�^�B/��,�zK,G4����"J�E�˄�p���W8���w;��cקe��ȸ·o\���=�ҍV��&"i�����w��u�C_8}��C�OFl��9�sF�=xn�T��w��Y�������E9�q���Y3r�6'����Ǜ��^�O�o皼dW�7��N�L9+�M�z��@�2�ظ3�2M�_���ݐ���i���|�k��zn@{[ץC�ol��Wh"v�ÏDbK/��dV;�׫���/<0����l��+�*7/P�f��\�d��{6��|q��ɩU�hT����#�ck[��.t���y�%�t�<wgA�Y�ͻ.���e�du�p�4V� �.s5%��,����`�R��䦦2��mi��O3�2G����b�4->���΀�v�B+�yU����aW=�w� y�'뾠yՁ�_s�+�r�Ӷ���2 V�5����ݳ��	���\v���M����)�!�5\�����Z|w�������Ͻ�[��I��Z��X8�;c{'m��ժe!�Ħ��u���m�&8t��X�=�1ϨZL�B=X�S�o{��M8��s�3(�K�ju}�����uQ�n�"/����p�:\�mB�I�v�����#x������#4��R�s�v�C^r�`��k.�R"*pɊ��5�e����x�,��7�Ϩ�N٤g'����l���
<F"�͇'��*(��9�L�Jj�t��cg%��\��{%s�AC%=%e���T��7k�7�N��$������+��Uή�lm�9�d��b���͔y���H{�B�d��)uL#��cF"��(�t��W4�����v�����׮veFB.���cb���ݍ"��n��U���Exk�.vn�z���nݻv���׮=���"@b��J7.��t���+�����E	�����Ǯ;v�۷׮�z��! �$?��)˾u��c�\�u���9���C?:������z���nݻv������Un(��\ޛ�o7 �+��j#�����]�s�Q;��")������n�N������q�Esw��grW�9y�3*
�y\����S(C7u��[ٺ]݃�|���wr'��<�
w\ �n�S2|���wu�)s�^�WR�"-��{�C�v1owsu��ǽ��׽�N\/5�mߝs|�;��פ�����Н"^�so9w]J/wJ�y��us�;��w~N�p��g~�o{i-��m�C:�.���ˉ�r��f�n^�\:�8��%�h�a>����VK�-c�]���w�ߪ�����y�8I�n���e��ܼ�g��?����齺u#K��H����V�4.2��s�`lb�}�zR\�ȥ�%���(�f<m��ڇ{[p�i�~��'��cG�9���^���*�Ǖ�[��{eI�==j��ˇzl��ō{]C!�e�><552��t\��3Z��1�I�x��i}�j2��;�*ޭY�陖Ss���mX;C��\dDbsw�޻�kή��BH�h�/G6��1-���k���a�+Ì8�f6�Q��QԞ�-po���7�~��F�}u%���}7�"��O�O�4{Z��,-f7vw��V%���z����l�-׼{}'�!�=���Ų}P_P��l�Y�(�S⦈������g�z�3IgOp<B���h��gC�����ܳz�Ҳ��u�s��D���j@����}���ף�UN�[H�y[��}��)�ŋSx�[}$��HJA��#o+7-'���Q��+E	���~J_$��u�7o�{��3T�M\m�g�܄�V�y�4�:��yϧ ��3u��L� p��%B�v�˼B-s�T��`��~�������O�o�S���޷��Z��E�=�ڊ���d�jW�}]?���w_-L���cl��Jʺ�T�=��;0J��D�s�ݺ����ؖVlv�Қ��=�����S�{|z������ ���A�q�e
��tgGvR^��s��+�g#*�I�S�}���IĔ<;��&�,ؾ�S���;R�4}ށQv�wh���W��u�N�eF��^ҍ��u�����R9����@�"(���Wx����&A\Z��Q2�b0��^fc7�֛���M�v��� �v����
��}��yi���thcX��N�я���F�/����|�"�b��ڿpZ��ULl��Dy���9m͌����c�����3�^�8oy�G��s>	��p"�
�=mg�d7�������d.��y{;ݩ]�(	[��c���d!y�{�%���dʣ4��2tiy�oE���H�*��'@�E�6^	�����!��|F�l��/a�#&���i������`�	ܒ���ZY҂޹�r��H%���K%6���8po�Jx������̇k�D� #ɱAvS�
�#�~���
���J�vj�g|$Q��'ml��[��z�ղ�78�=�� �'��2�z_���~>��RU�Ѿ[7=]���v�q-�m���{�,��l<y���yH�u1�ue��2Gn��$����%p�ʳŎnfn�#p4H`,s�� �ꀔP�ž'G��h�49��Z�!]���}���;6ok�
�{B��Τk����4]0��=.k�f\�@��(���gB�J����0k�8�<W	J�^B�Q�y~�_3�b�2�BSSσ���쌛6�?\MME�n΅�4�����w����X���և~FS�ۅ&7^��oU��&'����
M�I=�yG�4�F�$�����_v���$^@u�v�|���M%V��S�'j�7�O���VM�����\jL~ɟ{�� �ɶFՑ���u�B\JXz�b��^^�V�O\N�tv�h���g��
9"�@��(N�ҷȣu�7T��p�!{����&B^z��$ﻳ{�¨Xѐ�މ���5ǵ%�n�5J�Kc߭g�|�ś�P����'-@����v����fbKV��g>f��Gض���P��3پ���z��NG��fa�U˥%ٛ�6ԙy_��u<�5���1���s��Uy��}y���^	J4�]-t�u�dq�\��	�1��g;�����<oV�IRJ�����c�1m��'n�k
�,�Eg�d��ܨ�O�y������Z�L���B2ރ��o�
�CL�m�j�i�`��>��|���5\Qy�^Ί�=��R��v��b���=�����̘�P7M�ff�X#=*|���x�(������e�DEmܐ��N�q��y')�+�2�^���oL{.�j�����D^Q�2��'c,n�[Ds��~L���=�I��~��]�E��?LM��e����~�o�'�j����=�3��C<��½1 ��+�K�d68t��a��b~;��c�}jR8�0l�?+�MI��B�R���YI��y�Ι�e��MI�5=xzB6��y�������t����̭6��U3��ۊ�Am�]x�H+�\��r�n�<��'Z�Җ�,-��;�����`����+ ���I|�Zͽ�6ٕ����k�K/kL�V�<-�S���+j�G9�F%��;&���ܿ��/bѵ�>C�����u87b<D�	_�.~a)�B6:j�й)�i4�]��1�Xg�rܖ/�)��1s�[�g���{���K����D�[�!^��vf��^��۪��/<i�z"�qP�aٵ�n����mE�oLX�U�Ӹ�+�f[�8�u���+60�`�/�dv�}��U��.��D�b
 ��!w<���]�0]i�~=p�Ǌ��T�Q�N�lx���C֐�N�:�!�p�D�u�7��Y�s�r��oJK�q��s�Mr4�-��%���K��Y�����$�k?�u8��~��Q\h"�2���$T�+�fG�;��6���e%I�<=p�;���Dp�Z�A�\�ei�seܽO@��5Y���h<Uk`�ʻ}��`�Q��0F����ˣl>�S�ǰ�.5�st��_Wga���M�%Q��8�0#��$q����m���?Dn�傉|�o���O���!HN�2]^d6�u&��U����ʎ���nzy�̺n���s�H�=U��5ź�����TK����~vN�+���qw�/&���ʥ�2��e.T��W�H��N�N�/��^����y�o7�v���~c�?>�m�9C��vk��yY�o���p\�U+.vu᧭�'���9����ea6�n���z�Cv̴��v�Q��OM�4�4�{�X
i��M�dWs�}������lgA�m$�	��rճ����XÆ����i�ޝ�&�/��4J5�W]�L��x�֋��^e����g��i���[��`� �{��1����^�쌳��;B9�<8;n�/l�8�!z��/q"�U��u=,��z	C�OP�^G��-�Q�׹���x�k���V�	 ڞ�ǵ�Ǫ��t��\�� ��.�����Հ����u�ɷ��Ufǵ��+�'%Y�FuUx��D�	���M�n��ꌤ��z����Ɍ�s�1�Y�q%i�S��Cg]"��.Ǭ�9��kV	 ����F� V���{p�{�^�ʶ%��f�hF�-йtfYtc\8���O3����sGw�E����Զ�w@��g�7�P��w�vY����� �����$x���okl9<��p҆
�J޶fo�WH�afk�s/��3�1qŕnQK��� vs �:�t��]�����sߪ��P����}���oR��w�k��)7+��'5fG��=�����F��/�~~���{��vC��?E��6����B!�Gl#G^���Ogv���td3�ӵ��KT���-�[��d�cd�]�6����Ȟ�IR4�sqд(ݯ>�m��{Z��a�֫V�}�}u���ޣ>�p����*���؋��Wyk��Q���o�����~�_G}΁oXZ�ޑ�V��W)�dä��3���ڇWq��2:�[n9��`��,6��\zz-P�X�U�뽽��]��龜7vfE%r̃��+�"H�G�oI�'T.��]{�^p�u�=I�+æc�
����ge�:�9X��jg74�ĸ�q{*AMwƇ�U�3��{Kbp��ZW�����ax��4��!{
f�k2�c��U��a5��;�Q�'0�5s�~P�c27=���#EG�Ǭ���Y���a����S�־r�'�T�}3�L�Ʊb6v�� �no�t��V�>��k�ї�� XF�NK�G���D�f<�묝e�\:階
YB+��a�9������Rq�aY��+Xw���yH���T<<<<<*�[��A��Fv��*sۜ
7�	�Ǭ�5����Å�a�ڼ<��'�b�m�-�I=�`����)ZrVү=έ�;{;5.v�����i3�����_
��cz3��b�u�@A�Q�DeHl��x9[v��F��,Y[3���c�L��㎪w��9-1����^f��_��<z'����S�,}Շ-Ԏg
���[Afs�Γ[l�|��]���@ޛ+�3��=��7�ş�H.j�s7s�����ۈ�g���["ߠO&��/;Ե�5����kkO' 䥕�[|�֐�\�e�U �|�F��EGA;��k���j��yo'
M���l��Q<���r�[�F'u^|���JJ�1|�3a��!�����E�i��_��O�R��o2<�~wl	��=~I��s���^�s�h����or�2/�v�1��vq����rgMY�k���=��7��T�4�x�vaqP��Z� ��&�D�!�.��������u>��G0�ک�ō����%ξ<��0�-P}/���뾜����Zj����U�~ݟl�7Co��C;�!ԦJ����l��L���z�
�y�e�f��ng|�O���~�v�i�gy���`v�t���·te0\ʢV�0c*+�}�nb��;غ�V3I��u��Ў1rr�懔���Lu8�>�=a�M��O;l���17�҉{^6���Lz�G">��[��ւ't��W��:� �GP��1��+c�o3���Ѻ!�����ӨlaÛ�ٵ����zYŋqAgfT���ծJ���
M]y�^]��R��uxv��Q�d��U��r�gC ���Z��^�W��[élmw��T;�H)J��ϻj�i�1|;Ǣd)m��]��ѷ��&�d�W�	��)mx*����K}vm�W��� ��\юs�}���k1��V:q,���-�\u��q� �uyu�Cb���x�Lmr�ۉ�u~}&i��6f]��֔'�z�t�e�:Wd�vif�A��[<�q�����Q4G��qXS�}s���V\q�L�'L�����Ќ�p�����/g0f?6J۪w��b��+Q*ʉhP��P��U��U-^v�OQ�/�W�}�!��)�N&��\{Һ:;����7{�o0�~͜n>�(����B���[�6Ej�կ�)��mm
��ݻ/(��gv�V^�^:_�/�-�b#�׳a��>��{s	�Yi�������ҍ5��=�(��P��ʲ�k	�k�{�R�H*a�qMj)&y�����=C�S��(q�>�r�F�lo�|�Y���q��ũ��4���y��z�J�n�4=ǲG�H; GHb�/�=`�I�]��{q��>A�*�<��<�e���>���M�w�*���}n������P��j>�g�	4R9u�qOם�n��ZU���-��9Nws�2��,�i~��3��i��⡽^�op�<-i��Tk�:_����<k�w�/��)ﺺ�fWN�U����?�����Z�C��@Z�H����?������
����Ѣ���|=��@5�V�1�VX�V�3mf,f�1�m��5Yb��j3[MFZҬ���6e�,���jL��3j�͵,Y���-��fՙ,e���c3+Y�c-Yc��Lfՙ2c6�fjUe�f��1�-l�fL�S)��Uedɋ6�feYf՘�f[Yd�ZԳfL��L�Ͷ��Ɍ�f3,��1�k53-��X��Ld�L�f1f֕���e�5i���ʶcR�MFmi�M�+6V[R�3m�fڙf��+6�cR�����Y,�i�Mm+-Y�55id��J�m5&m���J�VV"�*@`	���>0J(�b"�`�����5��VVkef��6���VV���Y�����k+-ef�VU�el������VVV�ʲ��+41����l�@ 0t;Uue�T���+*�J�PQ �� �A� ��U ��E ��At����"��� �D)Y�����R�֪VV�JͭT��UJ�Z�YB� H4(� 2�T������R��U+5j�f֪VU���[^��ޭMF[R�ڕ�ib�jVm��e�VZ�em+6�ݭ���VmiY[Jͭ+6��f�������jU��+k����6��f֕���f��Զ�f�J�ZVVҳV�����sR֕�ZY,զ�5ib�jj3kLb�ZcR�1�kK3[_�>����������T �X� Y!��+�����p~��o����O<�����G���_V����(�ҩ�������>O�
 *��������**����_�������?�/�������?� U�����#��i �=���~o������W��?D�O����!JԳkKMZ[6��Zm6�ԫM�i�զ�jSmJʴ��5���5����ڦV�Y���ZZ�i���J��mi�6Գ[KR�-��5SV��ZZ ��$@�$D 	��iV�Ҷ�e�-MZm*ҥZmM�4�M+i�kR�kK6��5�٭IkJ�ԥm3Z�MjJ�i��5i��M�*mhզ����M�4�Q��[E��@YAT$����Ud��[QZѵ�%[X��m��jM�3V��Բ�&�2��֤��V�kK5�5i�ԥZf�3V�@� H0D��!(/����)�H����) � �ϰ�������� w���p�o��E h?:����}�kb~�K?�h� �=���?�<?B}�@_���������M�W�( ����<?�o�DQ���� U�
O��	A�V��4���a]�,������@Y�G�>�?����  �~����������/����"���A��PW������
�`/����D��$��Pm?������0�Np"o�� U�=� ���� ~��?F�h?�k��gW��"�l
��TUj��\�����
C�O�����)����C��8(���1!��G��$
�
R
��$��*���B*�QJJP(� ��B��
EBQT�JT��BUJ
�P�TQ(�U)RT*AERI*UU))IRR�P�UJ��
(��@R�IJIHD
T���QU@�*JE*=4�J���""*UD�
E"����T�)DJ$��DJ�T�F����P(�I$��
��D�����Q%DD�(Ip  d�ul�kd5�m�ΦЁ*jTյm�,�j�mn��)�MZ�kV�Kfa5]�!]���k*��*ڭ��!i��u*�)VJU�T����(�R*T �AR�  �:=C���!E������	(P���B�$H��n�C-i�l�kjU�CZVjR�m�3Z�i���:ݵ�Wv�m��ɪ�iJ�J��-��R��	@�R��T�H^   :�²��ҫ�l�e64��k2&ԭ[(4�V����Z٩�Zڭ�;�i��چ�m��MM6�͉6�Vۻ�Z�U�m��R$  �J�����   #��@�LQlX`laL+T��j�h��j֊�Y�ֵVh*�b����*+lQ�S[k[daH�T�QIT� <   �*�[V�Ejj��i�f�Pl�(�TCY��UV��kmUUj�Y�[P��UT!�(�4LCU6ĭ�EJ$IP%EN   -pj�A�DC`m4
֣�ٞ�#��@�"2�KF-�ESmem�*���A��j��6�As�	����J�#� �
V�,h�%�7*�4��R@
��JR��:P �wUn�T����wU�!��8S� H]�%ÂT�J��J����Ux � zu���R�J�"��v��gCZETgӪQ��r���C�nT�RP�����@���UΔ*��L�*]5A��$*)P��BR^  ��$ ��:7N�P���,:h�&��5"�îڀ���H":�j�4J���])GA��s�i����c�$*��DD��� �	!B  a��JWM[�p�
W:5�����+�(�h*nUΊ�)InӪ	V�ګ:U nSu�(:t���t��SqpP� D�%*( h�)�IIQF� OF��ڀ )� ��@  S�i0�U@ z�"&ʩ@ ٪4�f`1���fG���Q!r��y	�K��)ş%԰�2������}_W�|�����ֵ��֪��_�m�k[o��ֵ���*�ֶ͵UV�������-�'�
�U�t�U)X�&��Ջ�KSٲi�{����6Ηs��S�AܬƩ�9�X�{t&2���[���Ez�J���9�Fl�:MY�va�P�J�P)$�7��1K�y�J���Z.�L��f�6��\��ywCl)4)��4�;��� k�ebÊPy\eԫ�˱H�`�A��D]�7WlQY��e��ܕ�κW�	i`]5�����+8u�4�Yu7B�h֜gB�O-P�%Ӥ�R�[X�\�ŵza�{�jV��@V�7��;Z��	���w��[ՅL|�P��2�����JȊ�P��2��J�V�=�+'.� @���*O�
��v��ꨃuq�ɕ��8iՁV+5A�h���z^�f��j�e'p&Z����VQ�U��[`������ܨ�Q�lIu3�F@�^sG���jӵ���\" ֨�-b5k���ÅP���Uf�g�0,g(U(塂����Op$�����1��\�n��:[��T� ��(3��f�Ʒ(�ױ�A��i�0��sn�:��A�ETm��$(����+ݫE1��d,�r�h�t��(r�`�KYY"��@�VVK�v�������+)d��M�[A�/
M�	JP4.*f/��5�jE1�^�*���_U-2��P+����ʐn�>�UlдQ�vhm�����0��K�	�c"�����ň<W�-,5��0b9jZ�Y+i�ٮS+v���.�`�[#X4l9���&^źi��l����M���i�ɍG�Dٹ�����,5�3�+���YNQ��mX�'�P8�U�@;���5P������YÆ�J1�4��O;������y�����[�:OQz�S�ɚ���wR��]���f��9����J���&R��ˌ�ߓ��Ἠ[�Dk=n��^�2٣�}�Rv�v�4u��n�I����
q1M�m��OX���2�%�eF��k��d�D���0<�`�ud��˔r��n��TmUɎ�[�1Z��,�!�v�`tL�U�2HmYW�(G5�a!�D������S��d9�S�-��a3H�x��PR��(����bi)Y[����SP��⽫"�)�.�mC6���单�k�1�Р��"[�I�ES�4U��/!I�K��m^�'F�=�z�"�J�m,��X�Z��V�Ɍ�N@����{wf��^��*VE�(#z#2%�	Ĳ�Mt�b��az��g�p��]҂�2�eJY=��o#�w�M̕&�<Hٴt�m�$7��]�U�5#O@T)m5i)������*d����Ё�	�ŧ�oM���/�"���͵Ǘ)P��Zkj���(�ݺ�.��p���56���e�G]���E�*����]9GJ��2�
��[��pLLnԭz��6�%	2�`Ci�����EKWx�t����{aқ{HA���fP�#b�[X�{J��<�IY��M1�rX?��{+oR+�J��,�5y�e��1x5[���r��o(F�NhڻXm�����l`V���u܊�x1�a�^����J39�J�K�����f�i���J��YW�Px[�6��uZ�-�*ލ��lj��7W���u�lЂib�)\ ��+ ����h*g	��C���V��(`������(�k5���Q䱗x�ĥ��b��j��VѼ�!�*[8����Aݳ�L�s�#��P���iq��Q{N�w�4w�)렢S�I|�oe��(�j��.�8�M�S2,�mMSkT����(jI�sZz�
60��D��+6Q	]¤ߌOj�Yʱ'�l櫊Tb�6��e�5.Y�,�T�cٛ+2m�"Z5�
�n�͡X �e\�w��"f
N�VZ@��[.��F��aI ���U�׹!����PԈak���=T�dx�HO�X�,/���՜���CF������H7�Ս#��^�k6�Z[I��Ak���haݏsU+̢���J�N��T�uଶ�w�ar�[�6	����gFA��%��Q�soI;�^C�����ԫ[f�� �ڨ�p�:A�2��d�'N�t#tJ�@^��`L/TR�2���(Q�WB��JhL���&����n0���Bh;(�fع���t5 �4�*������AU���St���*���62���� �����Ȯӭ��1��B��IP�˕2[V�t�S6TC&˨��B�WZ�����N��A��Xuv�66�E-7lY���l�v�+YI��*e5�Ǌ!)%������x��n �-�.��-�R�D)S-�
tlm��.��uf�HS��Y_-��.
cZ���ˤ�⅝6�l��r^8tKGVi�΄^����j��"���ؖ���5a���n�h�n&%j )�E�k+U�U�j�7�ūX���!Ty����v�-i�eM��*VU�P D�RU�Mn�W)`��2M�ے���>f��,1��l�W�Z�6��h���/ޥ ��E�z!$9�0�v��E<�����od�4wEϞh��ә�e�ѻ	S�Zd-0
ߍ�+j����")�o �0��;M�vf)��ZGĻ���t������K��L�Z�/N�EYyKe���3@Ljܓ1���&�*
�i�t��q�������|�j*��<�	ToK�4��DB���ٲ��gXt(�=���YLH\�ghL����9��J���|�@�K�)�l�'*�wh�;����d5�twU�pb��f,Y)���owvYMb�1��+�n�+�ba�"�;f'��u�e���@;�z��X�&]����8ڣt�(X"đPʺ���֏�u6$�uk%��h�7X����u*J��z��X�ܳKH�z>i���ק�n�VReҖ��Ue�e�t�t���w롓`��
� ��HjR�.휠d�Ww��4+-S�Z�f{X�j䫌����K��&�-���zP�[�0�`�PZ:E����衹iܭ��p�l���V�̥�4�ץ���rlV�A�	<h�6n4b}2���^L�R�D������t�Ѓ��$���lFY�T��w���r��$�!+W��%Oj�yWWD�Z��4�-T�dR;A,��p�UwcCu��졒�d�ŭ ��LY���s� ����#��g�}G�>�����]���6�q9� c��˒�4��0wax��X�$710���#a,�xJ��M'j*Kh1
u���`R�;�m�"a��sr�F���ª��mm�V�ъ�B'��(��(q�eZR��d�.��\y@�b�D
�KF/�r�K�su&sC�Pn=N�����{ocפD�V�J����â������-PJ�����VKٙ�����Y"���>F�I�sfX�4�]4����];'a�Y��
��6��;nf�¿�f�I��+�`�,|���pj��e�ՍJ��L�[ kBT��.�lݸ�]1��-����o�W.fD��-T��0ec%Kx��5f�iG��J9� �j�u]i���%:Iࢦ�[e�pU�D�I��9���mB� Y���˦��d�D�x,���g~�̌
t1���*n��V:�+0�5��DV�JZ�Cr��ƫUb"�(�`饒�j�����k�Y��ö��e�Q����\4���K2���`n����9-��^ϝ	�E�	%�$ $��5�U���5ǋr@�f�1W�I�k.At�Yͪ�Ҥ��*T�X�֮�����O)�rz��MչN��F�j;I`��%<ʰ�����91��鹈J�)R���3jØv�	�f'A��4 �[(���Y����f5�X��a�ZP]���dJ��t� �)���pl�\��H!��mK���d7	�f����� qC�7Y�2�Ű͢ڼo��ck[�.�S�E�w���5v���T�k�V�xUrU�y���$L�FŃ.�%j <�Q�M0�2=�ʗ��F�f��&�֚Y�����n1�Q��5x[I��`*��0\�/15�����Sc�$�]Ff�!5���l�t#w4*�H9����+���Ǌ�����Slͱi;����oLjDF�ñ�&�a�n�^�TH�X(�[t�	J�Ay�0�J�5>�Ol��`\��2�dOjni����.0�,��ڲ^�M �Ѭ��뷭*w�J�Ж�W
v�fZ[R+%�S�2�*(VZ�x.�(�LJ��	�׳w\Y�Qe��.�3�F�ՠ:3�S�mꡗr��qt��E�֩�&�Jw5�t�jVA�'/A!Z�2��b8j�ljZ�f��A��ĂJZ�8�U�6�j;���`V�����$��rm��RBm���vQ*x�C���s0����	Ib*�0/�&36ތx荒�H�Oh�y��n�e�;z�fI.���b^Q��$V�S-�5�(!���J�:�CRS�O���n�{���ŀ�Y�n�)挀%M���а�h��Jf�E��;t�;�j��D3�r��fc�^S�b&Kn�o"�z�b�4�%�z̽�q�j�u���ՠU�����\�ӊ]�˲`YwL�+��Sr�j���=ed@���m້��P�	�2j"V�;Y�l�n̙�*j���)��͒��I��=�"�����&a�E��+&Q��S#�l���ZV����;SbDZ�Z���L[[��NC�J!��w*S)\*�[%���j�:�,b�L�.*��*�X#r��ȍ`oV(��i��,���+�<El:ìm�Fb��h��d�>U�#��k0��J��n^�C�ʏBeXL޺���Cе,cul�lf#��ڭ�m8t�R�ڤ6�֫��t���l�j���5Q�C,Fe��譨�Cx�|��B$��^��s@��6�mj�;�U�ʀ���jɤ��򻵅B�,7X�m�3I&l0��]��hm@��B�1�skhX���W2�Bܡe��V@6��"�)��1$�+@�z1��;5��g@i��m���n�ln��5
�#��Vѫ�j���b�Q���&y5(���,6f���VXWV,�G+U��l�Zk@�uR���;2Uନ�P�
8VP�$���kt�[m8m:��Y圔���+�"�n\A�$o+�t��� �TM�kY��l@�=��f&�0 �fL�R�cM���j�Z[0�7.��P�'��T�U�T����4� �e#qjͬx4�L;�m����%���-R��,3񙸘�kd�űཨ���,X�̬Vn["�cvH��+.ܧ��3t�Lc!l�y@Q47e��E]�C+D�U2�Ц���e])E[���U�v�f�+�K�\�v�d8�!��&��7]D�%����R����ӈ\�U�D@��	j]�Ջ��CqP�v>'�ۿ�+����{X���0����ZƖ`��n��n�+N�.�#S"�6��VsE�����!��m�+V��j�ܻ�y&5}�B��\)���w5ZJ�n Ƞ��P��ȣ%5K\j���Vh�b��tk�ā;4N?�mb��Ʈkz	�m�W�������e"��4@N��qq�w���0J�㗎�j�4�[�)�J?,��b�.��[f�2=aK[ba���{MQB�I �Wt��EV-�mC*�2m]�@"*�n�vNF0d�]�a�m��������֓5��̌� �J2]�\Ǆbj�)�d�̢�Tkj�� #�S�p��ތ,LSCŢ�4�@:dت�n�D��=�i����T���Y��
l���7[���ּ����s帩���i�`'E-%��E��\�2cU�mG^��1X.��V���#	�]�
I(ݐՖ��J�����A�D]aR�J��>�ԙ�SgJ
ᕕ��k�h���t-�YOrh��Ȅ'k �	*���wk܇�T���;��ٹ��]XZ���6��xn9�6��#�\e�aڲ��{Y�]L{M�OnR�����\9�,�6������+�74T֯r:s˥-��{W��"�]`@�)���\	�0��3\a��Y��S�ÄancV䥭 ��-�i�{j�J�͈��{R� U�d��śX,��B��wp�Ѵ��j���aSnL�Xӎ�6���&\���m���im����wJ,��A�1���Vn����ճ��8š�k4r�ZW!3*@b�9B�ٲ11˰�:%��a iYv�cf��m	���Xa��7)Պ�f�wP���)7tO�a.��<�F�J�Υ�m*�x"��^�j*�f+̭J�YÒM�v�!0�-Qa�mຬ6w\kaV�u�P��@KE0����)�1��]�x���h$R��ɦ��)�`�2[r��XAfH��JU�q�^ǯ������E�ŵ�aI�,�RjG[�K�9PH�
d����4�z2Z�!��Y�df��iʶ�A��W�H�����nζ�Jk�yF?�m��>��JνӶ��pG�b}V<�N����IR�4�)��yn�ס�Yje]+N�ȷk@5;j���R�o,�j��{�M���`P��J��kvؑ��0C�������¥f��g��j�,ުӑ��Z���МY�Ԑd��-H�e�էcUG#�/��en�����t�nkۭ�[���R�b2���X-;�i!g���RX(B�i6j�T�mQfG�rB�\9b�T@�Ǎ���mB��� oi��[F;v�=0��=$m^���Ѵ���U�C����P�<��v�7i�Q�!ػ..[�5�7��n�k�Qד\����R�4��e�}:C�9�H'W�<)_"�mp���8md޴�Kw���C��d|�n�\xR����5oMkh^�wi�/7y��ey�m�i�kk�X2�:XN�r���Z�׍�ռ� '�:�ZQ�k�|r������o-�nE��UI4=��<�a\��C������Nj��I�H��0�f45��C�&�h�Y�nՒ�ie^�cG��Wd��bu�(B�*��ڬ+n[K�Z)WWZ�.�z�P�+����K�忧��rd�ajQpu�+�m0������G���P: �x��Cf�D�KV�]M�����@v�4-i��ˈ�1<�r�(�#ei��׽ú����6��S*,�ysp��:X�C$��zU�7�L�T�'"�������v����Y\:�l��ғW��r�b��R��u�˛��A�u&gf6$��`r�;X�
��٤���ڑ��W8HQi���,�����Űy>��ͭ�I^9�޽}���Q��x=3|�r���ks9����w�Y��2]D(̦T�h�{S�:2�IO��Y�GX����v����ͪ�qsi�[�z,5}T�PE��(PYܮ*͊�ii�[��w]�z��j�y�b�8ٝ��q�q�2򻯒܂��N:Sd}*\N����sz���|�c�g&{�lW����x��&B��h�;OGw ���V�>۳���7G]�5�yܪ8]����ns���{h� �@D��p�{!\��76�f����*����4�.��e�v���y1C�)�w8����e�)�{yK}ˎ���k�c}̏�a�G2���o,�^��T�[��˔���u��nҐ*It��v�:�LѲ�<�ː|�rන��|}}�[�K�f��.Y�s2xgu/�ͷ��鵻�E���i�(�.8+��C��8,�ÔgL�xmFFw7�K�\�!of���nث��ޚG�\�]5�
��}YƝm���=��g7��y�ݧ��dz�;W�� �/��(8Z�G
L"���Ѵ�j�L^�}y�U�6�:H�n�+�6����N���Xr0��.�]jr�X����8�t���Ź��d�)�{zE��J�SM�+t�嬊|��UA7ӂЬagy�9Ī�f�C!���[J�-8�w���[�sf����/_m�ևY�-6�ҝ�r⦐:�Zȯ!�L�ّgT���2�c$��0�I|��"s���o�劉�6��2����U`榖�u����]hz�/L�=�xGf�X:��\ܐ�+�ǏzYt�̺t��wWĮ�dg��F���jv^b�#YM5��c��r��^&���D�ꀈ���S�u�.������3����E�[��������a2@5�\�u֨e�x#��h���WWM��r��|T�!�0��n�4���A-����3Y��Ү�\���`�Yλt�Cݥ+v�KhU���x�1��ѫ�6�A�gn�DV���a5����u�qΘ�\�bά�y�Pzj*˥n�j�
��(��kI'Q1�o�g�)��AD ��|�{ꏛ�e�Ƨ]{Y�����\:�b�؜��ǖ���,�zղ5e;�*����uh�#[B� �и����}HoIϤ�>���t���o,���;*�����:�罕t�z>��Q�J��Zs��X���PVqԨ��-��Q{�F��9W�V�8��P=�e�*�f��KB�4�M�6�w_>��[�Ȣ���s-���h����ARWP�jg{Eћ$�h��c��0R�^���u�����	݃0��tswv�R+�/�Y7O�%`x�ob�z
v��7�]h��E��rTc޼���Q���e Iʹ۾Sf9��,+��|3�m�c��u���&X���nWu�ty�*�G��YU)1�c��9��ۣC�Vq��={\ºb.�KT��[�WR��XZ��Z�LI�]%��tL����m��͗e�N
T�%��L
�<��J�/بE�n��e�[�CW��uة�$�Z��wSq������!x$Y����w�H�r�ݚ;4dJ�p.Ʋu��=Kf���q[q�(���4{�I�/��ږhopPA��ˮ;�Q|qӳd�Eh�v1H�MX�6�.n���H�f���c�����7ܜ���^mI�0�7�bhn������ʻ��]��ݱ��l�������ϐ�"@�R�*]��e���m͛Cf�rC�zgZ;/y���"{dꈕ{�P5(*Y&Uv�r	�U�_BR�y9�b�ƕX����s�Sܜ(S�n����nnq�@1x-�lIȽ�.�"p�mu]�X�yk����9���؋�IGr�
x/�٭W����lc���%j,o���O؟��%�\�lf��vecvur̩]g���m���Ѩ�El�7�p`�S�wj7[Ŗ��+3z���i�P��ͬ�[:=̀`Θ�*/��@�{`v�0Tw8�`�@)E��̾�/qLj�*9��pqZ�e����[�:��i^�֙/�{յ�e7�̝!}�0�����Ծ3!��
���n@ �ʽ��嗱�Vh�KUZ��ͺ%���'p���u�f���+�u�.K2���X�A���~���`}u�]����(bu�v28]ڼ��l�Ó��0�V����.r�J���e�X��HN}�X�DRώ8r���� �7��x1Pt�`U��#x�)�s���w-��&Ӕ=���ە�bj��&H�=W�MKT$�m�@�\�4���Y׊��Um1ؓ��|�y+.L�R��[�p|CrI�L�{soM���2D9Z�v�4�wy4m���!>�P�m��u��5�Z�첳GS]�3�K����7y���YDn�N�\ޭ�LV���0�[�՜uPDws�i��)l�g~7Kea�I>����n�w��,���<WV�A�4ou�<��f��}'+WEP6�u8��#>��;n�����]SZQoAo�u�cj03�/��GO<%�P�v�ia�r���oU^J�v�����U�)>�Fd��u�6���Hݸ�pE�v���{�����MN�*v�7o���T�����f�h�v#NK:�b+P��ﳺ�*�k�G;�['VX�#|q�Ɠ��欉3vb떵Sz+sh#xm�i�NorC�v��'7��d����A�u����[��!�ga�&X���8����柀�h�zj�m�+Ï��M��xU�K�WI�
Ow�V��2e2���4��Ǖ�۵7NMh�֍ZRа���1�ޤ�G�>9s�-���6��r�;{9J.��cL՗���f8��QH+Nn����vlŻ U�w�)�a"�"�U��늰��0p��;�Vj�%mk����C���֘T�n,W�ͪ�А����s�q�tZ'w��%�Z�`���Z�|�!#ܱ�P�l�G���)|r�E�7nGK�ui��>��.^W}j��E��#�]K�5��T�p�-�S���)�#�5v:�<��O��r����2��v�׈zl\ܿP>z��B<,�u.��^̨%�x+
�:�$�YI^�Q�¬�*��:1��z,�M��;ip��醗Fm8ii���sr�6�W	�kT,����ﱧ�}),X�зK��1D��r�*f�u�'��L��PM�v;lt*����Z*��s~Y|����V�W#�&CW�K+E<}s�e`�����Rd܉�4���opQ�=(m���)*��G�9����+����:X�j��₝��i�+�
<p�
����,��3Aט��ճ�,�)}e�aZ�$�Aį&�+<�m^�%�s�/q挠�
�N���粱��ڥ;�n�v���ZÎ��[Z��ax��.f� �ʻJer���H��j)��csf���=��{�����Z��˃�J��J9��A�p�y�[�ø���(u=u����k�В�s{0в����r9�a���v@ܻB��1md��9ChR_7���}MY 5Z��b�|��E��nX�(��Y�7�#�L��R6e��0�S�B�,��6-]�Cղ�$&i��AF��T_f�ͩ8Z]}�#��h��tffu��dCV�Ļ-�gE>�0��n�4 {-�� �K�IB����8�MΡv�t�x���&	K�Db��a��T&ƕi��\ͼ[�\���N��*�34*�X艙��C-m�ۧ��v�>�W��X��u=´�7'
J�$v	E����.�L��ҕ�l����9���7��_V���X1ʺ���9�ؾ��n�*���X������֊�6�O �c�5���x�����m�ի��4�`Z��[������ۡ,�u�x/`n�V�f�ڗ��fP���'Rm[v�Y��6��w%�'E�*�q��(�uک���YQ<����λת��C_ʴ��ֹ*��jΝ�%r�m���[R�Xyטyi�`N��2���QZMH�JwW�ku��ŷB�p��m���s�w���,-�v]"���;<��3`�8^\{�gƹ 6���w��5u�R��}ܐ�7MM[t�c��ϲ[�{������Ӥ��Ns��3��r��*)@ �T����vӵ9Eu.k(mEu�ky�`�v��6c9��vC9+W�{4��l�YKX��r���vҧɫc*�U��4b�ۇzf.��*][�%�N�ɭ����󦱫�#��&Vb���m�t�s0oo���kսc2�_va���p�`{Uyz$o����"s��=���gm=�@]]J��:Ty�hÊ��b�
�Jʫ�w���\��-�(۷�q�v��|b�5V5�=�R��fEڪ�l��V�[^m�HM��:�K��@v�{�����?k�-mv�rV�� @1�'���##[�G(��["�D�7{�R�w�S�xwOs��v�����>vyF�n
$^�&T�:ð$z8*nު�@��.��7�v$%��1L5�NNc��w�����*��n�[P�L��5��P�ҲR�AV��v��l��[���u�1�,K��]������+�S2�ʝ�{/d�}�u$�V���8p:����U|�֮'��@��ֱ�ȾW��kY���;�0SO,z�R��Tm;���<8Y�(i ���'u�k�)����'�����ut��o8S��a��&?$��[��`3�0�X���M5�����(���O_*]�Uo:�n��Kh9��F��7��B�A/��'t���H����ӽ}(qx�um<Bb��
ǒ�Yo�N���4����c�!�#u,�Ȭۤ��f�Ӻ���z>u(�[�A%�#ӥ�����ȳO.]�u:�_R�h�����v��Z��M�m!;�����m���5���4iJ���X�qE[�p��4�5�o���q9��qe�c�0�6+E�Dӹ���2�MI�X��b�ev���vA����+%q��\�����ƴ�_ǉ����+�l�YÏo;�->=�Iϯ��3��Sz���4G;c�d�Է���_����*��<��0�˶VNl4tJ�-��G��Ƿ�J:�u ��#�2�e]v%\���Jc�&I$��.[�=�fb�Dp�wx���&���G�P緖��r�v_�:[�9�s��K�E��ie*�[���Nl:3{���}�6�s��sZyԄ�C���d��-�/@(+9Y���Vc��y�C@J�w3e}���6�!����د$�5u�Qt�S�9��Y�&�}�,n�բ��ӱzz��I⧶�qZi�aqs�]	�y��իa 㥼Vd���^ww��GF��\z-�Sݴ�����KJ�_G����|�,��ܤ�t�>DS�\.]�AN��ҊJ���ۭe=Ob�K~�E;#*�٣�%%e����-���Z��G�c68�ӳy��v��:� ���(n��
��![>�ʀ�	����yO�v��9ݹ�#�C((*�-�>�<g R�Pr�s���em��6�lks��u_H9���=���XVʱ�*��,�A$JG��G�+f���s��P��{(lVT����#fe�宜ԾT`3�]��Y���m��N��;�X����-vf�8��~/6��F��vL��:�R���r�ɋ����:�u
rV��Q]fC��L��y[�����@:�h�t��wX�
��H'�3�.S��W����T��e�`���5	6��v�����]��\�:�㊷#�pT�|S´�`NW���bV`�i�tw�=���K*P��.�o�W)me:�R���_`�58��a���0:=f>Ӏcl�rk�eCHZ.gv�����t�j�T��v�+�w�:K�����\�[Y|�9QINVY/�t�wr���x���C��1����|△�󂯅Z:�tٳ���'��὘���*�F�wֵ3���Wt�י�Yqʓ�^pU|�.��zv\��:0�y�#��k����j�ݓ�4��tGWQ�3���u�����Q>6�*w+Vބ�(a����~]�͜�k�#Nu.xp;�q�,]f]vӥ�+�ƚ{Y��(Bo-Sj`�۾��;VV�}���՗�-3a�@���*�.�R��F���{�Qj�y�.��	�z;+�y[��7��k|��/��ۮ�FlVWum�
8��zMH:�s`��9+2���7rՈM�y��5Թ�]L�h���آ�S���Z�Jɨ	iu�-_Q��Ŷ�s�:�.�w̸�Rά�ͮ���L�3\Tw�D!��G܇*}���s>�W�3��ts�]�ε �}��;����֬q
+x�0%7�e_l�{4w��^b����%ʟFOLƶk��˴`�V;��ly�����iWn��u\����c*�5�ؚ�����3333{�o�3{���{ޮ����6�����6���[��#�սtʖ�����Ry�k��{D��ҕ;D�l^�H�/r�\�6'F��K�v΋}ioG�����)cE!�i.1�+�닐�*�Jf���[��q��:�԰:h����gbPם��+Ӕt��ç4Ӯ��d���Bb�N� į%��r:��v�]�8s�آH�di�}v��Z!<��yrԕ��f�-��P/�7b0J�߈J��^�V)�����d�(b��&v��;�Eb���mٳ���Om|�Պ�C����5�D��u��9��a�s�o�t�P�d�V���FNX�)�jՉz�M-O�5D��+)R�:�:�P�ͥ������Б�F��%݋��^�	�7�,w]uoq�
p�R�.��u��S�k�L�vv�@�-U�C�:�q��t��նL�u mm���sM��s�5���^M�����:�FYu��6�t
��
��h��Vţuu*5Ŵ��n��.�j(E�6F�F#@�,�K�rb�[�)o1���B��o_h��Lq�3��c��IX�Ty귚c�wD1մ��Ԏ$�����1*��ֹ����ju�6;l%���#P�\���͞昅|v�f^Q�	{�Eh�#e����ơ2V���B5�3������w[�Ӥ�3.��
�2��Ϲį%���u�JS8�&~#{B�EF���,0���
�焔�յ�|1+�W�К�tc���;�s�T77-��ոʬ`���,���~k��@�hu��C&b�p�;�z��ψ�\G��u%\�S��=&J�Ĭ��:�S���p;�i�[�4C����i�P4�5A|�r,��-����N!�Pb����S�Eg�8+:�3o�M�*!�v�f*&���h$6	|q�,	][/%�f�`P�J*+�s����AԺ$��j7ۀ�t�e�i�P���PhP���:T*h,W	i�I�g�x;�9�N$I����q�����=]����̬�Kt���윙�*�2��6��ڴ�����0��ĩ��9t�+�(�eh�r��j�@��h*�GpV�p̧u�D���]����od�R >���u\yP�qd�S�v�tr�ޮ�)y�z��9@���x��y�\.*|��ټ��Ú�۵�����G8�������Z�1$\���%��[Q^�uh].WJ��&`v�nBvJ�f���"�La�V%��l>�v�
K������@϶�[jmi+(��l;���1X�����¨��]�;"O.���0��FU��tA����p��)�y�������Ad�k����T���i�Pq�_lKE�8�#��r��yQ)FLUg8k`Owa��[(|2������To,P��2�7`�*�W#�%mY���������٣�#��i�{�P�"��{���U��2��)�DR���:ӎ7�X�wPN�0�[��,��|��j���U]aU���·�A��O6"�*���nɣ��4S���N������^c=���5�3ֈ�C����yGb�Ozj��ᬀhg-����v�w��[̰eӜ�pvM�t!A�8LT�;HЬ�^��U�f�xĊ%�j�9r��ւ^ �\F��qZ�)�����p�⹫[��"��E�����D+*���W�n�t�rHC-�I��k<5��c��r�͈<���>�8�j郁�2�����ZԦ�u��f�`��(�n*٢V�`{�j�ؒA��ܭ�_�y��Bszd�|�L����y�}��I�u�t��5���:ץ�ZŤ�E�6�킛f�fᶬrl�=i��G]����s �9�3i
5���D�r��Q��ނ����g�1�ի�4Lr���].��)��egkُ�t*DT�Y3%G�V?��Р���kE������9��>啹2�-EX�8ļ]�vk�t���j4(*�{]��m��Q����Nض�t	q�Q(��j�t��7�)��32��k�Dԫ�u5���RW/�s�I>谦X^���
,T�I��	����}�\h�ruG�gR4���I���VX���"�ئ���}����fqv��HV�"�גm�y��}3�Y��GB̮�Ǆ4�e�N�9�lEW`ܒ]��7�rwA�}/�NSuf�2C(�YC3r%�]����MD4��wp0�3�{��!Y32Ȯǥ�����VBF�D���T�S�2�r�Wc �M)�����a���k���Q|%�R���n=�e&^�*�d`,�j�B^�i�+�e��ʦSϖ�Y	�\2c��:{}�NZ=��8���h�ٚ�7�����#�W@[��w�b�B�X̲h�����7H��^�ʝ//S��޴�«T�K�,�iY��o�;j�Δ���(�Z�̽7�����..�%�Rhm۬6��T���[����F*��R7�� �٫��!YW����X��d��1�_LE��f��s��b�JMj�{��ʛ�J�[�fc�4�@59]2�v�r���nVv�d8@���>��XSuw�@hi�%e�;YXz�a��v�ms�<��'�GvJ,wt�B�Z�t��褬t���h�oq��Vt|I�HA�He��C1E�h���Z�E��,������Gͷ��<�^!�X�������BJiF�Ĥxq�γ��q=T��zF�ۭ֩��Nѽ�0V�[5�YG躄+tj+�gĪѪgQL�s,bW\π�ݽHx��م(L*�\ � ���oZe���ҴZ���;)s�ð�Uz�	\ �tl��]�e46j����w�a�K�Q9p�/�L��ܬ���KY�h�C���s�v]m̕ùq�#=[Y�n։���u�޴+wqS���de���g)d6����DvGa�k.�Ǝg"�5�&�Vú�$�8��+;/i/�T���4��ś@>�h۳��g ��ݕv���ŗp$�tыw�)�k�?� "ݫW6������y)�+1ai=�6Ї�!�j������б�S}R�'��c$�pses��ᯚ��Z��C�'��V
�[S1d���N,5�J�B�XxPYz���Ń �3qK<�x�v�\�W4�f���cqѺ79y.�@P��ɦ���,�;���2f�AB7��uh�:C;�8�Ԉ;��L�K�r�>>|���@[s)֓�:�UN�i�L�k��
N��2�F���)r�W��ګ\�:u=�8�F�Wκ��GX|G_R�]����ܗi�gy��@�]���e$�U��|�3f�YhP�i� �8�]3B�vy1Y�����W:\w]��r�4�x�@ �n���������y���ep��պCI0�Nh��N���Q�b���T�}��c��u��{��>W�1��Na��}׽G�++���{��Y���|���S7m�'�cΥ�5-�6�YWf��(vt̄3��J�!+K@e��Nc��+b�j��<�}�^������m�Lk��F�:��Z��s����Ӳ3֘ܠh\8}��D�.D))r5��	�S"��e�ݏ;1|0�W=�xhJ�n'P��$�R���A�	�n��B���ѫ����soy�la�^�5]ϸs�^�8֝�
r�;Dh�o�����z�ͭ��W��|��-��t5�z�ZbA
���KX��&�}!���! �,&C��y
���[çMqC�ʕ�k�+ʈ$����Vd0h��kS�p{�!�b��3>V^��a���;��A�3�Ӫ��b8��b�VV`�l��B�2)2u=�Mc����s+�<�W�
F[��65�`�C�-Y%�ؾ�j�#Lv$��Mqq��3��ٺoMM<;Qհ�>|��|s�v��%��Քf�E��Ķ�.��P+��&�H�nh��&�����<��1�*`�%op��(�'�MDnom��]sF�D�7��7��3�S�uN��� 	�t�e������gA4M9\I�%8k���Rr�6�Y��ArnrT�'g6ͱە�*]kT�t�m+xSL۽���Cr6irt,ie;���]����s�p�λ)��v�z��:���(r��V�Fpt"��)����᢬�b�r�eY��JV{1wB�)�Y`��]w��A�*M����ғ.��1�ՕvZ�m�*m��5,�\3y�'���sJ�0FT5��*�Y@�+�����k3��u�j��6>����sͿ�7p��V�׊�ۅqm���!�l������0��Qb�e�V�,׏Moݬ�h{�:��<+!��\i��Z� ٨d��¬	;�]$4�6]�����ma�W2��]S��f�0Z����NFH����z�u:7 ������me�*Whcx �Y4"u���R�駶������k8�b��쀃f�wV|]ۗ�z��2�;.Y;����j�S�K��Ƿq�U��N�
�qQ[���G�j�\�u��o��!W.�6�}�qzĬ�c���;��⫛�?>ǸGw֎�ٵݷ�+A�n��t� M!��B�q�]��o{wA�[�hƆi�'t�9
��P]���["��*c���SEH����f�h�;��h:�ӆ*j���=�lؕ�9�o�U��)#�w>ʆ�h�y�)�,��r�����Z�]A���k/4��Ʀ��o�R_)|�[:�B�gE4n�B��s:냣�dXr�^iB���-�EL�K�T�n�tmn����vn�B�k�}O4��q4G����[�����h�|F:]�<;WC7!f��4�q�9N]�:niy�7n]*�l`p=�j��Wnr7��.����֫�5@G�W�x��u��Hu�]�wC�v�U1�F[��퐮T��û��+�!σ\,X;3����S�ˮ�i@���h��N�)B��n��*C���QX�u�<O*��j��ܽqe�Z�r{ʕa�m�� � �u���{hT����ox]�D�ffQf�r��f�:���Z8f7Qr�r+bqܸ��K0�������і���pu��m^�}�,�=���C��ΧX��:Ii"|e� �)m7Y���Ө�W�r�T*w^�� .u���..�qE,Y���	����>�o��\�0�H��e���#Ֆ�ںZ�t��u6݊hvJ�7��otَ�.�5tn��
�� wPA$�ъ�pҳ&}t>���zr�s�e��ht����H*�����W^�%�+o��-�x\��k�J�맬�*�II˜�@v�������#�p2���B��fu��]w��J��N��Os�h�O0�x��:�z � ��r8;*<�,;k׻�S4�h�(�"([�2`�S��³Kv�+BV
��2�јB�8Wf恙h<�i��b$�tN�r�jŃe|k�p�HW1��g��:���b�I�#f��|9X���Vc
W9p���򸌎���4��+�]x�e&��p�[N��t��ZRb�X�)j�hoܰiv��Q�o�� I|q�LV@��Z�Bi�gdrt!V���eEs��.�J�Ok$inʒ��V�r��%dO.���Z	�d:��>T ��υ� ҭ[�E:u�c>�������VVV��xz��{��@Ќ<�Wx��Ӫ�7i�3�RUv+cuȰ� d���"��Q�����N�H�ӽ�C*>�M�R�8�'�ۅu�*��}��yֵ���3mK�qŗϗd��n3ms�rF'P�=�����R�vC�8JӺ㎕�p\W�s5�����G��p����̫���*S�y�ɸP��zI;�+�wK�|��B�d� �=ǩ�w�Vs����;l=N��B��4��&5ջí���Њ�u��c��kh�:�J�c$�9we�Ȅ�B���]�>��,p����A�o/���\@#Em<��$�:��ݚN%e�z��w�1S�muT�4��r&��콐&gS�o����vob�����@�u���怰�c];���%�x�Å�MeALu�R�3��jU�鯏K��G���m8��77�ε҉>� �˸�VΛe�ە!��c������t�{75��y��S��KX��ڲ#Tjm(���m���w�4���4&���s�u�؛�k�[5��.�c%�ю��� �౛q�w�7d����ʗ4���s4�F�c[n������MɈɠ�ֹdr�%�Z�FL�qe�ʁA��[��,�Z�phә�*d./+��	`I4�.�nۗHf�	ʡ�_ ���ek�YJ��<���
w�:#B��w��@�v��
�̙"�q��H���R�Ze���+��n�j�Qyd��/3S��<�3�r�����������s6ܣ�%9HZC�:�sȅ
ΧWb�w0��e�,�' [�e%�1ΰB �4�y�^:@�i�:�,�f�I�M��Dᡥ�5&����wj��i̸�n}��}��r�0�r�HWS�23�f��Q����5w�5$���~�Ҁn�_[R-��,S��S��Y�ٙ"����iY�����ʬd�-Q��p3|��e�������8����#���㹼;�Eө�#��}��5�bT]�3�6m��q�n�*���WIq�"H#��ʰ	�Q��I��Hma	�X�Q&�ft=a��I��ŕӬS��E�-��Β��Ǌ��/9"�]9d@��z��a0�8;o#�e;2�J�.����.���:崛�[6�ҩ����Ι\&_-!Y��%a���E_i���`Z�|;cW��%�q]����
��e��UR�2�U����=Y�V��#���	����@@v��{V%Ҥ�J}�|,�*$�i�c���d������t�K��:
�]8E�2�јEcsD:A���|l�7��PU����z�����.����2���4��ﾯ����������{�����ȭTPB��w����>μ��Juot���vQoz��emָ�P����3�u�4t]�/I!QI��â��j�źf�1�����ΦG$������ն���@o-iL���ȟi��]�]/ƳA<*qS���O��0�uJ�caen�,n��y�b�h�k���n1=�����m]�슭>+8V��`[3X�ݛ�jp�ф�8F���h�|�s��H]J�'��%\��]�wsz�ɩs	�m䅕�V�h[���G1��gh�}@u���e�*�&*��UJ:��b=���]��ζh�o%j�F
�Ż�y�&K��H���<�Ź%�7�Һոefm5��tF
e�5r��*��
y�Wh$qm��e@��[�e�Y�lZ�KIz(E���q�䯇���.s�
��U���hU�.:��%3%/l>Y�q�r��_gRU֫.�[-��L[[�F���qx�K�֪*���x��53���;u�����\gD,Q� +�>�O��8��]��PXE�X]�"j=����������.���F�5R:t��
�X�(w�k#�h;���.���%衴/��zp�_fvH�)ؾg:�<��v,k��'{غ'
P�w���
�����ՆPu�bowww8/a���D���q%�ۣ����qśp�wEDp�y͓;'a�g��´T/�� �T)�B�ɢ�ӝ���.Q�ws�M��	�;]��r�����sH�J.Nps�snQ˗!�s��s�����@B�]����r��.n��\:;�sQnwt'u���Qr�Q\P�gu��st���任�w���99w+�.�Iӻ�snE�\�s������NEt�ͺ���2�[�r(�˗;���r1˻��t�S�:��n�7wcs��������W(����r���wuв[�܋������s�F
71�b���w;��-�s�:���i35�71��9W\PS�s&��Lb����t��`���4Gr��#t���n�-˻�t�"wr�\��뻹K.��u�p�.�볮���Iwk���i�M3�.5҈�nh��j"4Ir썙�v�u0����۱tt,�*e1���˾�k/6^�	Λu��v��B)�z�]�V���Pl�/��q�ܧ�*�i䠲���y�|�w����7c��3@f����v̦k��Un�R�ιSwZ:���j��b�O=�GX;m>��K��窰�2rho*�=���,����3G1���yJa��Zտ@�2���.�Ol�n���e� V{�	�F�{F�+B��?vR�s�	��$K��K�Q��;UrsM���1�e��F8���:AWyT���Պ�۪�v�4�%��FQZg^%%y3o��P]�t��Z��w���<$���L1�L=^����w;;�V�ǅL<S�ٔ�x��Szh"k�z�]y��;u^�� 3�e�<��{^�-f��-��=P�ʹ���T6N�?1	�Z������xYVx �y？����!ƶRZ�]fתH~߹�9q�6�qek��5�,WPж��u֟0>�u]��9�2p�{AŹLS�yI�2�΃�5��$�K C��#E_��o��F+[���)+�Ğ�X�y/0�v_�����)d�'Z2,Ar]Ìw� lhw�$��˶���"��e-h�D^u(X�7�����n�N�7�ܛ��k����Lp����s*&6M9XE�3r��#�X�c���'0�g��nu<X�6���1�x��8h�[�H��X(Qݦ��(]S�;ymIM�9�X����k��r�J�^�s*xQ�>�o9.��Պ�|���^{����z[;������x]*GU;�eg'�zLl|@���y;��������U������&{=)a��U���0����C���ۊ�a/P@`Tw� U�pC��`�ҍn�u;Zv�n�ӓQzޅ���@�~���һ�X�U�e���0 �f`�,F��w��	���Q;k�=OW�>��>i"1�/�M��av8*�����x�ߚ���0�c�q�i�g�{�M��}��]sW`wd�P�UhL�/^)H��c����Uы*\��ؓ�Ygy�R�je���9Buͺ�n��%UK�ydyC�P�>Sj��=���5���7��i��ZY��\[�;���V�^5+����	Y��u}�` ��Z�'�kX5<��3��c�XCWDzx��X����W@�֬-[��kr���g`�;}=���n���bi��{}jrɾ+O}�^(�	?�TCG=�p�X#�'b� ���|ۯ ��M�4�q��O�����u���ﮎ�r]d��u���r�h����im0@�в��d� �7��؃��>���N4�]���#j_y���m��NcEP2��S�[���a���f��$i���orT��w3����sR��/��o�sX�8���^��	�Z]dU���xc5^����{���V�d�o�ԞH����v��l�����pڿs�t]T�tӪ'�a,)��Uޙ�ԃ���x��4���2���|�Ci�԰�ө}b�'0�����^��.�c�A��^��
��w'�q�s��2PQ:"�O�<��)B� _'�e�bp���)؇�ì��`���L��d����U��Z5Y�x$W��)�4"�^� �R������8u=�ۀ�D�]_��[\`��ʊ����0��1���X��N.�Z5�.�V�^4�-1%Թ�����eo�	��myN �|>�;����:��t�C��l��љ]&R�}5�䟖I:��,2/n�l=y%P1LHh�0��C�h��D�F���H���%Z����䥸�'mP2�Z�N�.�!yB�O]x�����+ͺCI#�>��yЃ+����8w6�w��VЭBxl{.}�uK�L��Qykb�S�z�|�s�n��_&���&��<��x�,�
iʄ6ubxeOOG���7����<�LPR�t��t�F���w��[�bı�\�]��4�S�n���᜹*_L��C	�3CCof��c�xA��þG�+����-:�:�b]Q[Ϻ��r��0(o�0z�g�����<�;q��^@�3#K�BN�X�z�ϥ���R��E�u��>��2�S5��,��+��
��V>��3|�]�c��o�����S��c�Y�r���/_&)׼-�O<�:�=��]�a�Պ������z�~
:�4�	W6�j^/G �@B���#-���R떁tc������_b�a蟀`�~�s-@O�H������]2�1:���S>ʳ8��n�'Z6n%�����.�þ����2��zd���G���;���Z>��4;���9��n�>�pQ��w�}�R`͵[q+�gzb�ך`��V	OS�y;>�c�`,��A��BO�ʧB�h�Z�~�'�w�X�drOc�GȬՐx��b<���ewZ�& c,rdo*�m��x\�?h�>�;���p�w(q5�` t�i�N/��}�cd�p�xf�
��|d�xN�W�����q<��η���xq�����5p�����Q� �[T���z<%�^5�s8�����eeh��ϻ���]��[N���������=�,Xuἅ�۞�z���q�v�mQ��y$
�*+p+�J�ՃvK��w؞�>S+�����D��WJ����sO,�wy��g�5Yܫ)�,N�����YOu嵝�3�m�絭X�t�UKJ�B
޽��lؠ�W��G8�����?���<H(w:5�@(V������h�:���^�`֞mNm	RN�N:��*J�-��Bsmq�D
���(kɅO;�9��H����$BvB�9>���>Ҩ�F];:�U�QJ�o71�^�N���ꔺ7�\�':h��Ἳ�� �[\�si�uG��S����=}���n
�Z�D�Ұa �x�L}���������;�����x��8r��/�f�^Kv�9��0���/�i�G���/+�Y��μ�P��0�ߏ�5���{B�6}vc�3�ܼm�ϋJ�z��0/�����!�wO}��Ͻ��RQ��*1p�B��ם��{�)��N���x�d~Bk�u�D@�r�Y����ٰ�]��&�N�!	Ò� ��y��?e�J�����`�G�C7��Ƀ��a��+&�U�m�������/L����Q`��w�8�>o^vv�2� ��V�B�O�vc��!��&���=���
!��jS���1Z�`�(��n
�2eon�.�Mb1�K�G"���)83d�͞Ｒ��
��9�
r�w��]{[�����śZ�.[/s���%"z�9�����S�����9��I�����<��ivp����w�!�[}�^��vDa��򦾜5�R���C�
�@s#>7�N
�G�io����A���y＜��AO�^0���&U��ڊ�T`5�2��S���^|�\� O�w>5���u�s�<�_`{��ٛ���I����3��w嫅������٤0si,k�D�n��5nE�<����&�[��h/ת�=�T����#2�zNZބk�C;�r�����*L�m�ʥZ���nd2i�mNdǠ�PM���>�޿�Y)dPʘOm�`?\~������WX~* ��<�ڝ��~x=�����Fw�`�Ʊ���;���U�����[�3�|���@��D��`?���v=�@pڝ�=j���
W�9JA�����ގ%z��)'�/^)u�ҔPC��@v�H�0w�#_#�n�����XQ�9Ƶ��'\e?j`�.�X�^��,�Z�߁�n��@Ev�����^�潧L-t!yw^�B�z�����{�׽6�{˼K=� 3�
����|���tb�C ���(��Ʒ��f�����Z�9~�$)�7[�}�mc�����YF�r7�v�T)V|�����u9��Hm㾣$��d}nt8֩��s9ގj��:�Q�,Lt��5m���X�U�Z�ҥ2����p��c	��<#n�q�7��D}���L�[v���eج�(yfJ��F2W�� =?�{�e�9`����#�tj�Q��axߍf�6�&M�T����/�W^'U��&�y�߈{oP�rKz}��8�Z�]vkѪ��C�XK:�m���j����v�{)��N��֑w��F��렇�\���vҨ���EWYc�����t� {��g*��� 7�9�`x��&!��E��w�ˣ<�Y�^Z�Q��V�ٜ����eS�xc5^�.�:�b�w"��[ǚ�jqe[ ��0�Fg�ey�v�JX����K�����Q�n���f?1���E�;��K	}.�Խx�IͿt�%r��뼸R�=D��P�n�����q��	�B�?������ڮ��u6:�=V�Jn�/���[f'�O�	�����sT��v�!��>e`�V���;��E���"��)�4"�Mk/���瓛�]����\��4��J��m��+��oYA��`:>]�����JqwJ�����V?V$�d*�%�3�v�.�N�c�a`�|�<Sn��i��n�/$�8wg]0��+�wv�i�C��\���2�޻8���ZѴΠ��p7�ʯ�lj���IoFt�U���;,#h��8Ҿ��8�Eg;� ��ǋ������ښ�u2C�����ೲf��ٜ���=�`f��TE��c�u�myN «��:���]�U�nṏj�4>d��j3���<��J/n��"���`�{����Ɖ</Z=�Q Q���t2�>��bJA�p�޸���L��x���E�Ρ�2�(��O8�;�b}�� �";N����6g^��5�=T�V���5c�;x��Z5:J�Oj!�����"���v�h4�������7�R=�}Z���!�K��ą
�i؋�n*��MT�
!' ���S�t���s��|��_�Rڽ��G`���r��y]�L�d��ê���n��w���f�Z�s�͙��}�*c�)�{Ɋ������Ø�j�0~�J�^�<'+��]E��6H��UgU��`L"c�6� 2֦P������!s��l��~Ҩڱ��xi�*�
�N������ ;����8.Є�](�^5����
�ln�� �g������ra|�U�4+;�L4܁ft{]F�a�eRNa�5�3%Y����w�E&���;���w��[F�����K��񞒰��Dhm��3HC��*$I��t��yp5��p�A|A�2
�j�<A�q�P�Y�*v����G۶��U���,ۻ�A�o#��s��ېԨK	a�*e��_un޶乃��-t���9��.�������)�6�XxG��5�q�B��lsL����5�T$�j�B֩}�&Qj���PN_��?�ѯu�E��+U�J��|%4��S�wbC�X����*��/a5�oի3Y�:�k�̾^�~�5��X7�@�Q�	8��v���S<3L"~H�VbB3⍝�����NK���8�J�0;�k�V���Q� �[H�4|ꇇq�J�'�Ǟ����O�8Ply�f��z�vW��T��t�W������X��F�t�N�/�C�Eg�
u�]�׼��
�<+»
��8�T����c�r��6�+R�jfS�����q���g��:,�xں�*y��p�!;!Y��l�`�iTA#.�]�%^c��K�,��pZ&ׇ�۝O�V4����F�N"��v��!N�ӂ�k�]щ^"0hɨɗ�����%�*����\��3J'�\ܥY�^�U��k5mu�7�z҆J�g�\��t�'tߊ^Kh���}��,�x�3�CB�|�������Y��׌ǴF
=깾�)e�>����n�r�6�w_�G�]?�Io'RA�[X؛�CMUy+M���6IC²��j6$�蔧B��x
�d�C��89e���)�&+��5��,J�|wr���Z�WK"&ynn��cd�L.�;jJ�-'���D�6+s�@����Y�j�s�;��$p��}N�T��5��`U]�`y�Ug���l\�k8���
Ќ\5��u�k	�,��Ҍ<N��BSL-wǦ�)��uu��e���FKfP��6K ����<A5=��0`�*ă�mڿk�WV�E��_��j�nZ�
�{n�[���ҧS�ؔ�ꜷ`2l%�4�Y��=����z�ې�6(	<UhT+��n'eq�#,�y�#+_��B���qڬ1�*$<�N�<J��z��9����'�Q_@��Z��K��l����[�(4�56j�ZQ�y7�.�tĪ�}u{v[�<����#�� �pw>8+�m�U�ҫ�͗�� ��[(O��"lRlu O��ATU2NԤ�u���V�m3���,k�D��b&����v��{oB���ix�}��7�u�~��,��B��Zul�"��D/je�u.����_����{k��:`�T5LCjz4g�>r]�I�:�c�3޿�R�A�����dk�J�W�wv�a�m7̭P5�8�ڝ�Vߞ%.�J���F_y�>���T~�v7�	ư*�]�vͬ
�u�G�FV��K�~�X���rMiq�ع
;�j�,��L��*��_H����e�H@A�C�R�r��Dč^r1ݒ���AÓ��&л[Pb�NM7t���JQFV���R����s�����v���{w|�K2��z
�u�E�z������`VQ��I&��^��ln}�[��c\��	s�V���v2���ԩ���Z,��ܝ��B�v����5�s�R��b��k����\�Q��S��-��6g ���_S�:��v�ы�κI+���2p 7�v�\yv���n���*�m��m> ck���)�9>���O+��.Jw�I�S�Y�`�2�ۯ�W�ƙ��#w��55]o4��.��| �C�3�/^J���c��k =Ψޅh`�[�,�Wj�H`ּN��M ����}Q�WI�B�9�b֕һֹ���$��i�8q�s�;\����s"��m�w������K��4��􊮘�`Ĺ���VZ��<�tuly�N
9��wh�'I��Gb7�:�}*��˭Z��J�r����S����6����zH}0�Q�\��rA�X6��J�v��i+m�Dm�isL���:���ZB�T��u�SΛ9��J�頛�pk{F7p�NuNʘ/�{�uVD��̧Lv_Ν��X̜q�!+�X�7���C]�R�w�)K��M��ъ�q_���Ʒytp��`J��j�+]����q»"*��b�Cm�Q�8[�;,v�뤨��8]�i��*ݐVu��w\���s\�2~����@L�c/x� �^�*�e�]�80�����4� �U3���d٬E�:��|�S�i��-���k�I��(~�N�lle�v.	q��+v^�wu�9���+U��2�)ٸj�m�NU���wnD4�r�H���kn�Ihl/����9N�35�}S//5�K�����r�u�g ����&v�;-k����S��e�!E�P�7&u�:���jl�_4;��m�b��鶯��*�C������^��F�5�Rq���:�O6�촷�+�ʶ��������fZ�(YB�ъ���[sv�.�eYo�J�Wt��6�j�.p3���_8l�rB��:c;J���R��2·�6��$d��FV+:���<�Zc�KeY&>1�īl�p;ڨ>�M����)�z��� ތ.�n��U��23����fR��]s�q�|�MP��XF�.���P�����8,Y����X�yqV���WW!;J���ww����x@�w�:&5:�1q'�s���VWwr%��K&�E��}S�����[�dPVnY�Jb��Z�h���Oz�4�p�8-u:�eh(:�3Y}2V9��Z��$�ؗv�q�:�b���j.�&��Nu�o�SD��{����;��V���"��ņw1�b�",1�i���wWK����s�cF�r� m�ڋ��wY9s\ܔ��\�n��t��L4hM�i4��((��ܠ����b.�"Ww
6,���tbC7wc�B,JP�v�)wr 9:�nj�Fdb�������vh��wc��X���2�s��HI#'w39u����0'W �H�Ē�s� �r�F'w3�wP�`�]D،Ar�FwF��r"�t�����آ��s*g.�2!9Á���#��n���.���:�&.p�%:���E'N���"H�f���3���7P�R[���63#.q1 4> ��
���c����������U�Z��RE�w����M3w��7]��T�c��,���@�m�M�-����δ��ս���ۯ�ޚ�^�{�^��zZ����zEx�+Ž���cs}|Qx��6�79|��zU˕���[w޷�^->u�m���ߞ�͹W�����ﭾ?�n3u��F�8ns�x�d�*�뙬6�6������[�\�m������v����wo������V��w�����ʿ��U�[��W�~v�;��7���/�{_�{^-�\��^/տ_��KA���y[���X9�k�!v[���Gz�|Zu~����鷍��|����n�տ~��_���n��w�*�U˛�ϾW���Z��_�=���վ��-?'op���^7/�^F�<����菍���=fy�&f���1���z֗�?�~}�o���+�^׏�;W��_���}��^փ^�?�W��+���|��η�x�{m����;�ms\��_��<��_�������?;W-����+��������!U_�V+���Z��gp��������y��{noso��/_����j~z��������o���zo��5�~z߫�h���|���k����<؊��+����|������?���W�^�7�6�(�����33�p��]Q�d�g_翞���ǯ*�w�����->u�k�w^��mʿ�ߗ_Ϳ^7�n^���/O��W��-��x��s��~����Z��ۿk�����_��h߷�ﾶ�ݷ=._�*����.��+�P]r%X'���>��?��������!|j�`���+��W����r���������ww�ֿU���^��W�o����y��^�{{U�s}m��������8k13�!��q���-�*�6��_c�����o�Xr��a�ohBC3v�4�P��������k��o������W⽭߽o������x���׋F������_Z�/kA�޺�W��U�{�uy������|\�5�����~{���{���jV\�杊���f���ʪ[�?�����^b�������z���}o�oj��K����om�ۚ�����^�ݷ��m���o-�����]��|[��r��Ѽ�x�Hn#�#����`{��ۺ���em{ݹ�@|T�AT����y��77���}[�\����������{os����������+�Z��7߽^��ۛ_�|����oo��{��/��v�-�\�Wj�?������w�?�Cʺ6�gR��.�s���5!��@T�0�軜���=�����TXx��x�v'W�\��|q	֮�eԊt�Ĳ�Ñ�;����w��`�w� �iE�$e����
��Ҕ�'�g2���Ț�7�_sj��w�2.�g���v�x��-�����v��\����6����~~��U�iݫ�������ս��>���}_Z�|_����~-�oϞ���_������W,z_[x���?����?����}����wz������߫�_�~,nU+��|���z�W����ߖ���M������o��ϝ���Ž����>�?�ʸ}��Z*��+\��Rv|�����߾��kŢ�]���W�}W+��[��x��~v�����i�}6�W����ץ�>5s^�w�zW����[~�?~z�[�ە{]���o���ۛ�������C���ߥ�a@�
-+-��������[��ſW�~����7�~�{���~7���o����W��7��ߝ�TE/���-?ݱ�z�{U˕�����>v�6��ޗ��~��w��S{�5��
v�'�$⮴�#6�뎩�>�?�??}���o�nk����{_[|x��}�Ү\�m�^|���k��+���}�潮�ֹ�7��|�~�oO�ү���wv������j�9^^u��W��u��������ޡi�-�:�h��]�㺚�#�r����c��ת[�5�� �q��{|k�m�y������>���������[w�}��[{U�s~��|׿ε�x��z^�x��Z���[��魡��q�8�{��o��06��츭�������箼k��j��/��-ߝ��W��_������\�Z7�{��?�o�����W���=-��[�~_}yW�η�x�|_��<׵_��r��������5}�T�PoP��g6�Gp�--5�}3���>��ϻ������Wۻ~�m�ە{���M��7���ݷ��ݷ�x���m���Ž�������Z����?��7������y|k��k���W��^[Ң+�p��������r2Z���nD9���������W.^�ݯ����}��}���zZ7��o?�o�x��z���6�7�no�]�������{\�W����߿|����y����Z���m��|zR� �(;u��z2EMl-hU|�Cɷwm����瞖�_�{��y��W��u{���_���׋������h��O:�-��Z/�믫z~������^|�叫�����گ����{��~��oJ��B���,T�wČ�	���ju�j����)W��)�/��j��U)�q&���|���b���^g*`��2�s��V-j���VvJ�sq����Cϛ�qq�MfE:N]��{ ߚD��6�5&��Qy[cm`��v�7~rY��T��w�܋n�����딊��n�ew�i�y���zY�3�{�S�~o����/�z����7��7ߝ]�צ�5�_��W��x�W�G~u�o��o/�~�KF���}�[�}mޑ� y�38oXfy\V����yǬ�����8��g7�ӷ�3@nc�:=�}\��޽z׋����_��>������j����ս�ھ�޻��w���~7�n[�Ͼ_����s~�����{U˼�[ûW-���+�οU���s|o_޿^?��Kgܩל�W���h����nf�����k��/����W�翾���{o�^y�7���*�ם����o���-�{Z��~v�~����_��˭�� h���36��=�=��2���u��2k8�q}�Xfl�Ǜ��H5��<~6����\����޻���^��_��wm���_˖��޾����ޯ����~m���Wּ_�{���\o0��ۺ=a�7�h�z�0������>���<����{[���W�l�����}�v�*�����y�����.~{��o^�����o����ǟ�o˿|�M�/�?o��=~-�s��m������u;zyA�3h�RaU�w�e��m{�g�'X?M�����=A�t�8f�̃x�^�Ϟ|W���_�ƽ��\�[����Z|�+�^yz6��������K����~^�|^��q������oa��2�O���pj��8��Y�@�Z�+����c̜9���y8��w��5��������5�߯=v�����s>n��~9����o���x��w��h6"/��^->v�.oA�f֩���p���w-ͻ"�^�X�o,nK�5���y����}��o%x���W�������߾^�r�����������_?�ﮯ��j-����?z^|�_����ۻ��|^���U�6���n���r�[������/Ͽ~���X�#���a�{�@o7z�g�� {ּ_�߿}[����y��5��o���x7չ���^~��ם��������ߊ�.o����y^�;|m⯟������.�&p]J+�=Z7s��U�s����.儳lN�W�x�S�\%I= �����U�ׯΕʯI<X���.4�o3�o��k:YQ5x[O���}��d�p�6�w�H�؟'AY��۔�����`Qx(ly����x�XW!%B�̣��pݬ�&�6��N�!�}+�̷ș����Üժ�ffN�:�q�k7
,�e=Adwƹ,yMd�9���>�>}����Ė�t@��0w�1*�7+V����}����u��dn�F	�Kx��k�l���N}�=fV�G�P@QӃȶ{�n[�.�Ty�E��9�J���Պ�t���6��*P���R�}�Q����x̦k�ӫu£�N;��ްW?6Q��=�E.�s��X��)��B��#�@��.�(=�Ǜ�'5PIM�g�XH�w]����/�]�+��wy�;]�`y��� V?y�r���R +B1p�S�}7�m�}�v_���2�꬚��<�`��֊?s+���h��l��͒�
v��V���)���^���� &�ƴj�dj���yY7*� �{n�]soҷ���꽩��+u���/f��Ү��7����5a¡�i�.�U�P���Ӊٔ�x�����,Y���*�bf�>ޘ��둂�L��{���@g=�_���@s#>7��g�io��C��-�d�}m��k!ɻ��Z�M� 3�D�+�iL��j���ώ��G ���υנ�Vl��}�|��7��|��ٝ��� �1g�a��w]<�9�+.��94<u�Qخ���g-���|[�Z/k|n��<��<�W�be��U���3�=3M37��9S�qϹ�L��A:��<��7��`nu-�M��ۺJr����ĉ��̊38 ����EZ@9ģq��������@��
�*�'jRe�Q�ӱh��X ��h�{����g��#{/�T�c嵦������Ax��[�p�ۦ��>H�!^1�_�E�/��2u=�Z�v���7�bm@�,j���mNdǠ�PM����e��A��X5޻�}�$Ԯ�8�*z�tk���P5��}���[Q{]���|}��q�
�?gC!��~ŏ���JX`o��]�G��=΂����{����[���plm3^�$�~����ɘ]��[�
U�J��y�z�t�p�@v�FG���L���!�)�����g��Z�{S�+�7�)���̈́W�1UH=1��0���q���0�������Û�T�/��͎��P�a;04�N��
�y�4���[���1�ܡ�3�Y��پ��x+�B��l�)w��-v[��u�wzFjW�}�_��@��F3�sc�5q���^��er�a��*�2|X�]f�|�ƥa�l�0p����W��[�[��b�L`�<�猞2�]]27@��gdB�;z�x+q��+L���[H<ק�c�[@屩%��ov�և��ҳi����;8�m�bB�u�8��XW|���;�43�JW�+`G�+�����
ܥI-�|�[ì�O%u]{R�rJ���V�!�U��xf�<�%$.t�
oX���h��*��UOe���Y"��W���`�[��֎�
��z�7�����_��ُ��U=�t+�~߻���c��!�o�qX��#8a�������]�{�k���~��|ۯ+�xgj�Z�Y�OEl׾��V�fr1�Ga��7��'�Ų�+S*��D店fX���˺p!�T�pb<E��L�S>�g%�[5\>�M�+��V��+E����k���X24���* �/p�m2�iwN���)�#>��UzCs�b���z���u\�lRg�A��W�K^�����LWL>~SZe(X@����t�n�U��D�"\��~�S�?J�㤞uE`i�>iW�KF�믯r���盺<�)��
5n�g[t�4�e�/iCh{yJzW�b\v�}[Ȫ����g˸ϩ��ލ��4j7��dp���ɣ+}�ƥ���Ngy��g�Q��c�u�myp �;�ǫ�y1_V�Լ��{շ��)�6'�9�^�r���:���:�`�{��?8(��H�Z=����P�z���P��]��λ2�c(��=�v�8b�g5��Ѡ�P�1����f�E/�H4�}��Cԩ�$���}bA�[�*n������9��PY+p���{�v�AnӺQG�m�ֶ�WmeZ]`}���U�9��C�iP����+KfV-���������{:skk`�T�}S�v�ּ�^c-�i�:�Ѕ(�.���>*m<�lAޅmJ�{�pOh�R,�!$K��yW����ikr�sa�����%S�N�Ի0S���z�I�_V&Q�m�w���r��ar�rZ�4V�L��^� N����e�&z��K��/��K�M\ �^+�ꊅ�v��PYg漮�+ןc�c��E�̻}���s��s-a˻}qM��By� �Ey(�Ҹ[B�yv�Ӈ1�J�o�imN����~���D)ٿR����y��5;�
�~o�g��ފ��[��N�����
�u�{�k���k�ݘm��+(iw�X��ꕔ��bt�!>�Jg�Vf��F,n#cEpɎU�j���(�G�	p�5}�(͉O����_==^{���SLPlȜ[��a>��+Ԙ�I���׾����e
��A�r�XxO���rvP�Ƿ:j����}�Y�/�J9���Ng�;��Y�`�{��(�?v��Z�Ji{L|���Hp�����	��JR�gk���mփ&+��|kVP��:�~Kݎg|'W�;h�x9��=@��2��0�*���Sj��ҿe�B2�V�G����!��Gv�c`!T�Q6�uv��Y����
�r�ۜk�ȷL�5JV�v��	�(��x�o"Cnx#_y���0�-Żq����E�Z�ڪ�Ǧ3S���t���'�����FwL�R)m�C�Ys�1bmШEb���@N�j 6��_�<�zP�� �#�X��G<�L�R��u����>0;�v�����ykN���]�8�ؠ�V�יT�sl��n�A���g�"�uz�ֆ_� %w&S�m`�6��W愩'kw�u�eE;�/mbҐ=o<ʞ����tלwrYc��Xf���C{T�W����<gJ�	t�Fn��Q.j���-����1�`�wL�{^i�4�a�K�Gu*}��t�a�g��say쩆H���%�rsUly{l�w6���"#�N���\�OaώR��6��^���-�w�+I�輝�{#R�ڼ��Fj^��AĲP��W��#)�@�`�|����itqA�<�IX~�����*c)w7���h�=��Q���İ�����< �~�b絜JC�h.���	!�]�)�Z�ª��\yO�ͅ��6'��Q����(��l�U��ي�\���x���g*z����H��\>�7��֥��<�w������Km�:0G� �[�㩮ワ��ruLY�[)_]J�B�L�����i�ʻ�N����3d/�h�B�3� ��ºw�[�S��&A���e�qGْ�s^�q�VK�j����{��3VE��W����Zg M[�\5P�c�ߏ���G�v����]�����~&*<��L�fot{K�$��Q�
���]�eW������O����
���Ew�Wlx�˕��ﻯ��ݑ�����Q���q��ڒ��On�)��!��_��it��2��X��	�o�K�g� 2�@l�:�J�A���у/ڲ�,��Cn-$�h�Ek�O}�P���ی�jc>���]nL�o]Ho�
���;�Tr����Ղ�sU��NA�1{��=�[��j�����cH`�����h/T�}�:Ǽ�d4�Zu�����C����qͰ���Ϫ�B�p
��hwr���o�>_,=���Պ�|�`���A���sB+L�j��"�Y��>� o?��\ G�S�xVߖv?�U=Yd���oonzmb��Ze���KE�D��PΞX�C��=�DՏu�O{E�_|s�r�O�5v���z����^�6@u�y��z�t���M�Y#
��z����k���*y�~����wI����d�f�Uw�|��5/4br�� �u�ڳX�Y���V��[�p.����w\@Ci6F�+K��t�
�R�v���κO��)��w�K��r)���Sv�\��z��t��#��eb��D���gﾯ���(}�b�[y����;o���,�嘥:Z.ǁ��߁䧚�
�4��w�}d☋��<d�nh�Î�����;��ۨO�����
w������<���ty������Iyl7y�ɑ1n�gEx`�/-��^����v\���H�,(}fd�0|�{;Թ0K�fMe2��y$�����.����s*�W�
W�^�|�Ƨ�x[�l��f�m��=�ބw2M�kg"��ifWDe%M8��ۇ7������7f�SU�,p�m���@�,~��{�8�Z�.�z�����v!��j���k'�U]H�{w�ǆ6��7��+���^�]�I^j}(���q�]�z��@�C 4�!�b���ժ�E5/-z(��0�:��k |�y�1���=��ȋu.̵�ܰ�gr�G�T�pb<E��^J��f�g%�l�0�0��WL��p�]ZCW�vh~[��>@hf�xl�΃��O���w�x��t�%b`��+�~���75���G�9`��)� �+��"�O�-z#k���0Ʊԡ�L�
L�L���[S�Ž���w�U�aV��)�ɚ^On��e�s�LY�`�/,R���ٶz.�)t����q�n�]�a�΂ݍ�#/�&��,*��� ��LG��7ħq��Bwoq�4�1�2Ս����6֡BhIu��zZ�P��)V�'[Z٥[:*s�ҡ�nm���}��79ܔ7��F��\U�=�mS/�J'+hj8!��<�����`ύs�U�Q����쩋tm������7�E��XÏ���Y�u�������J�����k	n�w���wm���<{���"/h�w���N_ϫWs�"ͫ�qEwX�,�/�K5_9���"ڨ��BJ[���T#@�v��U���sp�
ɪR[�c�V�iub���7:��[�D@���Lu���͟2�{0���c�Y��ζ`�}Ղ���7iz��{U׍gE;��x��|w�[uJ(��t�x��c�V�L�N^�=}0�׷K`l���U��� �����뭽����]2�X���e�����;�Z��2l\�T�ܸ̕�X�;F�E@� ���Q�;:��R����,�ԋ�Xj��^�#o���Hq�⚩��F�Ɂ�9ж��>/sW��/}t���M��nl�٥�Y��{*p�=��Z�݅��˽Dg_��b�NK�<��|(e-+���[}��Fⶉ�;4r6��Z�IX ��)�"l�H�N�>o�2�����,a��qr����j��7���ڣ�G���sjȘ���c����`^�`��x�X��@f���]��͎w�s*��>���o)TW�	x!�_5�w�.�i3���[X��f&�h�6�1��\J׼��Vczo(��ۺ�!�].�=�_XNv��\�S-�V��+r�}�nn� &cc\.��ϭ��T�y�oP]��4hq����%����>b���Է�Y5j]N���Ήr@
b���x7+(�7Cj�I�c� �/kv��t��F�YA�ޕ�L�Yj��=�q���{�=-҈o%�F��۷�r7����
���}�a`�k,$-v���rZx�(���0��'�*�N�Q���@��n�P�������IrPN쌥�(���C�f�wy�6^
,JI�{{�k�V�N��k����5\�,�Ý\�[);nY��7����&fVJi�\�Ú�	��(��󶀶e�Ğhf��۝(Lм�S���;X9��f�rZyP+�:G��p*Y#x��<���t����.t�;4l�+MJV����hvP�^`#V�'�gY�Ӯ�}l!L�dd�ݹ���9�_,��9�ڱ�au��VmK�Ah��0�"��ޛ��>��V�Λ���uh�w�X`���S�W�xǕ����i3:�:0���koRK{mѮ��K`eV�84���L��RzY��:�
.�#���&��.���j�iaT�I��N'[�О�����[w�lE�
��u��4 �Q�
Q�Y����I�2��L7e�ۻ�:'u����@��\L.���"��p�����u)���]wwtD.��hC9u����! ����'w܊�n��;��FNvBwt�.W)wrSH�ss�t�H"Lh�t��0#]�K��1K�8+��ܣE˚1�4n]r�B�5q9u�sAf%��%0���$��q��.�n���	۱�)���DJ��7wB	3I#"����#0ȣ��D�2A;� dܻ��(�@,#��@�ۻ��#H�H���wwu�Gv�J������bwt�Np��0��DdcLJ!�rH�Ewn�+�P�!��Q� ��C���"���v� Ļ��m�w��ԡ/:�P�9�2���ێ����s�[���K���"��G�cӭ�1ӻ�&:麑��mԦ8�����P4R̵V󥼃�O�%��w�*�,J���sx�(r[k���d��7��`q$oP��Y@���J�N��c5Æ{��W��OҮ���s˗'{{��vok�'��)ėthEڙ�@/���=��*T��6��������s�|��Z
���63۳�V�t�g�&�F�i��m�jV� ^9X���C���6��q X+}�d�
�t�c���b�ל�]���
���n�S�$�OA�rήl=2J�d(��fȌ����i/qB�&wĺP����^c-�i�:���R���P����z�9�tq���vz�"�~{�H=H��CyW�p�4����sY9hhӪ��C�'r��7v�,���{U/�e���b���~fUr_mf�b�3���4��Y�ް!:�0�m������d-t��*��~��,'ڮ�;(E]�,���n��^��ܯA����ܵ��u��8`�.��
�]�c����e{Ɋ{��)�'X0{L9��>@���X\w���vb�g��
���Ow9$o���>ҤB�jeϻ*Ʒ�[�.w��PѴ�G���=���m@Ŝd@�S�ٮ����g�F��[L�Lv��\�aʂY��:�q����rư�_6�v�(_�������>Z�́�v誽�����]��n��W3*�I�UƜ�{}�rIy^���%�ŝ]�q֋��=8��V�n�&��33{�)NJ2J��̷�{�.&���q6k�1�]F�� h�7��;���.���y����'�4�)Fo��*��=Ih�����J3bU>Cڧ�xW�/��g�xU���xw�,ٯ��B[�`}Y^��%�Z}�e�Q��;�]�4������1MrvL{oJ-����������idu�s�"���~���i�ݑi����G�Ҿ+_�����w^�,�y"X�DG%v@߃{nϣ�V13�ZԠ��W�=��l=/,D M��P���Ǻ��-~}�ȝ�������kþ�O¡�[�y�ؠ'l�Ra��|6��'ޔ1DzW ��~�u0Xy��|��r�B�]��K�-\��щ�{cg)���zm0�|N^�U�T�s�|�؅Ep��6���@e�,� ]��T�3��c�r�,��X�ي���
h�P(ӵA�M>s:���X�͵�:�� ��;�LOI�B����|8�UC�6��cTh̦�Yze˦(��2*���KM��O��H�oէ�C�Һ��Ҫ�ew ����Q���#Fe-vl����e*��V>��d�C%zto��B�:�ߝH�<��t�홥�+dk�V�;��}m��wv�C�&���I����[�|��Y�CcM��ձ<!N�z �]���/�D�]��x(�}�Oױ��,���y��{̈́����Ź�Q1�&1�����,�C�b�I�I������Hy�����d�gt��[(��b*b=����$�K�0��8�J��^$e2�n�T��4�_�U���\*e���e����2=���U�Aab��t�s��U U��î�m%�/}�� ��׉w2����
`C��-}��k�q�a8po��ۛ�ڼ�N���(N��gh�SD����u���TL�@��k������&]Z�.{ep�����D��8
�q�,��|=U����x�(�PW�@6pʡ^��B��>A��@�m[�vNYB�5d��p����������|�~X�����3C>7���=y}r��*{��r��o�ynbO~ 4�� Cf�ԢUB�#��s�������	�)��ʳ�����-���hv���BY�ԁ6� �b�{Ƽ�x^󹣸�j�#���w�@Nx����K{'I�Vj���!��#�p���0����>����l�^�����!(��r��i�=)BP��_ ���x�\�,S2�~�|p�巹^įj�I�m_1]�mk9Ë���ӛ�����:ք����Q��sk������r���o����ee�b3�w ����ʖ�=Qp82��[GO�o7���}�ݢ��S��x(�	�܈!Q8�j�_���T��o����N��t,Sj�D���r��m�L�.�K�3�����u�^�25�>� o:+@Tp[�N��o��u�>%�x�ڌ�w��w<�.��T��,TяL&y}�4|r����@`T{����n\���D�[8ʛ�j�߫��z����Ƽ*N}�y����J��M�.�'q\���k�Z����z=����g��ƴ�(yb��t�PAư"�U]�<�n���{u�p^<>��=� `����^�i�f��w��N�@�0S���V�O8��r��E6l��+WX^���=pk�f-� K�l�y�r�v�.W_w�f�W�}�]��[�� B�t��iz�u=W�����֟�ڳ]�AU����+���6�;�����..o�;��3t�yJ�WOm�^�eu�>�`�&uU�@�b����])�����`�H���wM��<���\�< ��qׄ�pS��ت{6�0iy���(�S����o��~u�&����j�eλۙ�\cR֝�2k}�-e�x+ۄ�ʇPj��=z�y�a]�S��â{3s3�Ηc��@|G��Ws,�젗a퓝�{b�i�s�س7��W�>W)�z�7�9�m𧸏Uڤ�8n>fù}}��-���	�)��U�UW�^�x��ɥ��mc��w�f�@
ղ�1�����[����tjyl�K�^�5� �� ˆZ�a4cJU�-�Wb]3�K*��Y�b7�@�'Hy�8�j_h�;ƛ5����ҧ=���J�>ŸΉ~������p%��旵R��xf���_K�u/LT���ڋ.�-���gu�/��_��R�ZH:�m�pt��gw=;,ۮw����S�v ߬���7kcm����%e��&���S�_I<��>��SJ�4����g//�z�'���'�\�oس֬�N��
4����*�l�zzW���C�����@<\;m;�sf0�y���=㦘�!-��S���h״����}�TE�����y�{�.����an�L�2��)ğ��_�ꥄ�\ju6�!�����z��I/~u�usa��*��*h3�n���՛���tnR'��x���:)�=���Z�/��Ӵ�ߙ�6�A;�w-{C]�e��?KѾ���L�acT��Ԉ���c���^1�lӫ=㹨��Z?z�c�:���U��cY���q��ݒ'.�]�+����X��F��W���k縮�$����͔����9��(�s��U�j?���Y<�6��&��W]s��%Le�WH�0�S�`5|/lƟu_Zw�Sxn�{pl�d� LF>��Qd���7��Ͱ�^����%9�?��U)��4�������huٟM����v:�/Yp�>=���;����NdkeY×W�	�T�
#Y(@D��:�U�}p���v�Yg漮˵�V������@ħR�3zCL��,O��D��pT��1��iV��u{��)畁6��np�]b���'��m�2�����K���>kt�n�(�<�R!Mje��}�xT4
a"P�}��u9�(���8'0�>����=�٫1�%�l��p,B|/L�ϱ5�A�l5Ϙ,����ɋO��vB��=��A>
<f"3bS�=�a����^{�C����Y�G��vf�&�x�W�ɼ'���g�\5�6��PV�+����Ɋt�:mfߧ�����]�f�}��R��Wh�jt�BO��t-w��m�c�v��\>�1]J���2)):tX]nc��7Ŏ�X���Q�(-�U�^3S��0x��Ni_V��r���m���\����;��<�a�}��/P��,�#mNW�0Ȩr�J�S^q5u����<GKSXT^��[Q��n����w^�S���O0v����ЫzZ�=L�aέ�O.�k���\�R����`1멽���dE}/c5��v0�I[�n�:�]��uc'X��n�F�*��o|t�|���������y㷼=i��C���C�|P:{�:�%9Ip�2��xv��<��u��B�@�;"�n���篸�/L�6�V�|��t����+���<���>�c�<��Ձ�����Kf�aW
��t�t���k����Z�;�L.5�0�V��-.�gs�����Y��7�Z4�.]��wL��4��M4Z~gI#�h (���]3�ijCt]{��N���f˒��_���W����{Ӯ�����k
�=&*T�{^ָ֨�[t�S/�i�V�v�ggk>���iܱ�7H[f��YtK%u~/d��Y���:�</�*ϭ�s0��i�N}��X�S�c>��g�j­�t����n�|��2����͋��پ�%H^,��v=xuY~P��� VW�-V~��3����'��E�9��(��ձ=����É�r��xS{�N\3��CP\s�Sxj�j�F���Y7-p=u��@�.o�U���W����s��߷S�xO�}��;V=[ŹPv#-r&�N���C�*�����I��:�tV���I󋈫�������¹�'c�V��U����o��Ǻ��hx?�Y�v�(h4{6P1=Ni�V:��O#�fl�����P��vV�GS�um%:f��ԙ܌��>��'pWc��CozҸ������O��GO����UW��f;�+-dP�J�8��E[˃��o�	��?t;���F|n��OV֤�c~��Aig����L�����z�6��3�D�+�TF���+������ @C�G�=G9M�w/Wf��3�O���c�d�K�ɔ�}o�
���vPa�7Z66��*U�;{���&�z��I�I`{]ti�/E�ŕ*�u@N��x��������i>�z�]ܨ=�^����Ȃ�V�P>�U>iV�Μ�L�
n{���P����<�^�}9�W�-�j�{μ+�dkǨ�B��qo�;�i�p��OgG�T徼�a�;��J4aQ�בּSF=	��b��<�qW�v���xߚ�}�K�d�:JM���-0��>ܦ �m(���S���K����"����u���3ۊ��Ol<���w5�!����h:;��W�!��X�P���'�8�E�*�wd8.#U�h8�Vfk��5S90��*���^�i�f��|�ک;;�h?w��s׆��g[���-�"oR-��À<�+���g��ꛘ�z*{���mq9D[ ���P�O�:jtU���S.�z�)�zXu�(�ou��~yOם9z�p#���Xm�ݷ]l(r�}o�����)U��{Nζ����}��ȏAjL���|N�3Ɽ�����7��f���4�Rhuu��z Y�z��^��~=����n��o���T��Y�}e����/4]Z�>0���H�a�����p���gƽfç��j}Xx_�/TI�~����W����R����,��g�5��L���R�gҭ!\�r�F�J�������yv����x<���V��?N�Ob��۠���o���S���m��6���ilZƪ��j.��x�(���;>U�S}����^r��]��u>����ע�{-������_{@�IC�7�ڌ�Z��F#������5F��g�ey�v�P�"2�\-@�_|�v] �ճ��R��N���,^�R� 4:6��e�A��'��A^�ēx����Y�Vp~����Q���
^3稃����
���D�m{y/�f�s��䨴ʃ�ǧHҞH쿶�ƊN�/��e��eٲ]��/��B�;pNeG78���6��wཛྷθ��q,��׵29M�Lr|�^��JT������ɥ~	g��c��^0O(��CS��YXC�-�>�x�㈁�W��w��&�絃����z1v/S��[A��^��5��֪R�����ޙ�Kۥ�
�U����{�F�*�y��+�,�;�C5ݸ1�A� ��۹}$�G˝���%���:(��S�o{��{0$m�	�Zc�w��s�TK���Vޔג��ܩ��C���*a�T�S+��@hCu����@�3m�g(�
�
�O�Og�#�&�#/[0lC���Y�k˓~�b��L߳��zB��6�F�Z����bnE����o>�w���Y�_wNN�/'�v���vy]gE����r�y�Tj/�}�kκ=H�V�f�(d�S����=��hZ�8�r�\�Y���"rV�M6�$b5��Q)&�E��5����NH�6���T�^�t��;.��̊��qf*ƛ�Y�/N&Q,�Le%�����cpz�hh�d�$���.h��
��x]�h�s��^���:紦�V�>S}�lR�г*.�����ϪҾ���Ëj�z���2��#KSXr����)�$�	f�ҳ��K�c<�-�q�NXqnuzj�3��]&�w�9xe�9��-�����J��Vs=۽�u��v�M�b�l/s�)�{�ζ�Lhn'��M�1c4��\��g*5Z���a(���c�)���x��r����ӵ\�R��gf��0��0��K�M�V����L�� �N��B�33a�=v�MEj`ܗ8eӬ���-H�J<��r��ϝe[�c"�O��Y[�����8V��N����"^��R���-*΄��د� ���3:a�Lҕ؉Noo�t�U�&|����}����� >�KOU�Ȩe@\MfaY�7�M��vE/����������C��q�Ѧ���P�Yl_^ov��]�f�+"y*t�L[ӛS�o(sœh����c��pW=�h�@a7gv�޻�T�ΗG^w��ݑ�e����0��->K�T�b�P�H��ۼB�+$|5#,V,�ٍ�xe�L����i,R���ax:��њVyi�CX!�^-�S7p���QV��)[u���X��I�y3E��w�8eM�[����>�P��'k�6>!۠m÷�N̦r�W�%u����_Wb-ZN�n�{ c@�]v�������ܹx�an�>��q�R�`-��W$ mI`�[&��(���P�\3�3���ޫw�ٽ+#��r��[�IC6����`DhVjl��H�ݬ�s���*>���`x �^q�[�A�;�-:��h�e�VR(�鲒R;��n���{{���B$%��.rZ��F��h���4
�|j��cfv��N^�}��ɮ�,�����I/z(��k�
ɡ��LǛ�++&��3��4�u�_:��tL��=�5���=�g3.3)�y�'/!�UqŰRʨ�(�x��b�����̎ZG_e�o�����(-�򻭺�V��j��ٔ8�ʮ;ڲ�p�}�PQ���F�ڻ��
S��٬,��f�$8��,�!�D�Ozo^oltv�YM�����NH��.2�\�f�p<�7�t<��]iA��l�Wv�AsҢ�����l�S���4~B�\X����c�"�[ƃ�#9vf9��u[��{(��[ ��G����<�ɍbP]�l3�4�Pl�\�8��R;�W�!�ూ�\�{V��6���Y�z�¦\�f�w�6�![��b��Vf��(�kI��w�Jl�:*�a{����8��R�*U/hp���B�bj�ɤ���.Kv)��a��;�t�f�<JB���l�a�kNc62 @I�b�h���>�q�Q�}u�ҋ��Ef�TՕ-�����w�bz]��\{�A@�fܮ����������w�J[T!��R���2�T֐J�m�Y}�"�˾�2�Os,��mvi�p��H8-�]y3/�|s�u��y:���:��>�γ����]ܫ6���d�&B���E�q`�)�^��Zc�_�v���ǝ���LM��6Q�,��&��Jssgw8�4	BHD�]9�x�3�����f�)��s�w\j% ha�+���6MΑ4D�e��"�x��4�J���r�:$H$˦3%�qf��8(����b	;�M��nwv�/�	��#����pN�u�P����0�.\�d�I,���ws$F�3����CD���(��h����u�7i��$H�%˰��##�㻤�ݻ�J�n	�����H�9����-ۘ�.қ�Y�uɦ @��!��$3"BN\�Rs�S&gu��s���9ؼ뙍y�]�&�;���H�4sr"�7)F ��b��Lwwu�P<��CJ%�����;�$�sr%)�;����&"�d��d�����W��~�y~�Mw������+��K�!h�B�| 7�j���������a�k�Kťn�z�;����fv](����������Ł�),���\"��MfRW�h�lH��5o�{&�WB2�D�߲�AYg"���d\��MZ�(�*Ki���c�$�e��*�A���>h�\;y��MKnB5��U�J��[L�����\�v�s��=���I�%m{����OmT:�Lj=[�bdn�m�ʹ��h��P=RA�"��4�����^�1�-�	2��U1�q,��״�;���ܾ:6Y�ε"�-�]3��z^���a��X�Ly��հ��Α1���He�1t��lV)�&�-��=ʙQ,b���F���W^O�H:�Ze�ה��n^,�������I脕�2�Q,bN��V�� �(x��h%�	��/7!{
��Ф�Q%-
���E5�HI�Q:�l�����*uPRqF�$�l�g�0��-��f+$��6P�I6*/,�[;�k��:���f�U��,�92d��r�䔤Є�rh�WYgW]��s�FP��V5�1ou��ϻge�\ܤ�NR��۾�W�WԷ<�o����Z����R�R[�f���L�MK���z՚Uܧ6�ܵ�NE��Cɼ��@��6�<���W��UU^ļ�� N�U����f�Ks��W(�yT��ؙA�"� 4�K��My��%]�#v���:�eY��K��_g+Jy���bQ����R2�R�{�=���g��L��Gڪ��5=��]b�_R�u�q��2�gwz�k��x���g;3�<_��'�x�G��ih�^��,�y��X��+b��)4�;o�U�v��Kl-L]Yī3����CnY�hΑ|I�gn���/FF�[,-6͹lөAeImVz6jy�� �/r^�"*�ݳ|zŦ�^|��a�Ϡ��9�c��,J��Ғ�^.�#z��`�Y���mBj9p�Ӡl>3�:g���腤˘�k)]?W�o$��s��/�}Q�����3U���2u�������H��t�[�I���e\�*�ꪫ�㖎�&�W�X�JU��O��>3�Zf��ݣ�BƋ72�)�t��6d������0m�o԰�c!�5���=]Ⱥ��e�XKϭ$�v%�-�ٜ�t|��S��.���V����4gX��]�ocN��ީO��7)�Y:���S�0�����N�r����'P�2i]�x�����G%�8{���{ޗ�h��:�j,�9��inYY�YZ{�2bJ�S��}��ёM;�֘JTY�3h�Y��ΔMX����ƗT�X�9*��WXj�(�����&n/TK4��T{o�i�RЩ��
��.�Mc���/%3�ݏU����cG���{m_M���fN���(�ϗzfV�����b�W�Y�f��d5{�OM����W(�{"��{��g�b�Ѳ!K��m2�b���+E�ba���K�>�w,�mb��1�<�3w')٥Gaa��
�1�=ꚉ>lL.-k���"чw.G֤e�N�ȺM��*=u/�fs���O~�iy���X�Ei��=鶯�u�=��8��Y<J��m/Q��uٓ�k�Ϣ�)'��x�-Wx�1�OzuG���[��n��5��d����ط-�S&��2q�׷��r
���}{�!�t��*�QevyJn������AI����nS��MΉm]1K��燚�{l\�ҩ�,Qx���A�oeuN�VHUg�c�罁c����b��TR�#��M���&@+���h[]ʇσ�%�F��X���߫ꪪ��k}K}4��'?_�������znutڵ���ukۛ�>��Z9�4��f�VS���B����M��N���D^�x�S���j�J���WMi�KVS1���.q��:ڿN|��6}���3L���e��o	����4��q`�v�dv��NZȓ����s]���z�IJ��;s쒠��������i�|�L:��!���FL�����j�=�6H)�a[�r�,��t�l+���!A��e��՞����D�²d���\gd���W��s��˭]����ﭟHs'��<�5zވ�d��U(.�/\�0�O�����J+s��'Zn���yp��^�PT�5�/mSSG�R�peC3��f<x�X�z�~�z������tM��1&bX�e�b�/8��U���[��y�J�{x���iY�u�[�1�Y][Z�#�%1�����gw�a�̊��/�t템�g���qo�s2��׾D
�v)Ok�\:�]&�4ּZ�wh#�y��"v���^�N�KC�&ؼ��
�;bP_gs��R���٣�3�!��w>;�U��}�����s�~L�X��k̾Y�Os����^���{��{�)>רo��y��p�z���oj�`�6_�y|�g��ީ��ǧ
�%�E���Km�M}4���]1L.��P�������_Q���ҵ-�Z�(i?M�'��Q~J>��6T~�^+�ih���Xqo��躣^:��[n,�;�+3VM@F�.��vMe��47e���	�_�o�ɚv(/���G�0�[Mn�=Z�(R�(�h�l�F�i�@��g��=�(�����^��c�uj8��c�U�L��ZKiIYF+M�,r.{��k��਺��&d�7v����UsTÕ0�Mx�<3V�U���LoY^�Ȗ$B��5�֓&pQ �3WI��'ڱ�=���ҩ��N�{M��.f�p�h�ڳ=d�2��}�Q�������t�4�>�ؖ,3V��kZ�͋Q4���f�6{e���xr�I�VU����ܻ-�rI��v�+�G��F�H���2�J�UJ{�>y-Y%�)�.�jQ�l��9��X�ԩ��;倒N�@jY���\��T�[(�R�.�u��(K���ؖ1ncN�������R*r��+���H啘%���S*$�9����lq�"s��A�B��,�2����/}��J$�KB�ODK2K<���}�ȭ�޺��D��b�s{#Y�{#��ݪ
Z�t֨��1T���(��y�bW(��{|��t�ѽ��z����_J��6P��I�S1x�5�f8�*����v+���2VH����Y���\Tzzj�Ӊ�b�'bKjk�Ȱg,�i7e�*�n����j�л�K�mu�^�}qъ�i	i��oE"�bh�Q���U,��U�*��z����W��R��K�_3�aU�WE*N���K&�V��B��b��/n�O8�}�.�9���B6�n���0�=ƽ��z�B�����zz�g�E�)��&m��v]:�M��\eq/=������e�����lөB�q����ь˻>�J��A&�Ĩ�[����r�������U�lΛ[��Vv�n���7V��iȫ;����~���yt���;�P��3�	h��o�2�s��oS1��v�7Vs�v�y���wF�dx��L�
�ޮ��uZÏ!����^���~����ﯔ-�z�*��_ztu�í���d�#X顨�*�Kv�Q9V���3&��guWqi�(�ۅ�l`��>��-4ƠŔ�S��i�)���̉Ug1��m�Y>H�/Ih�s>c�g�v�"g���FV�qxr�7d�4/&����Z9{�}9#��My*��(I�]�1��pKR2��fc�iquDSYG��m���k�����)�T:>GD��2�e���y�xk�0���p��}��q"�
�JJ�Y�'����Kﶊ�YDӚ��|W�X6?�[.�[x{N��)hT���^����.za���8����iz���k���t��������ݭ$�ݒ%��l^��vJ+�N���pׂ���Y���J�GUl�âC�q�T�е�t�ɦ7���-~��*>h��fz�z���z�o���[Y���1wΗ���D`�}��Έ�~g�S��_t����p��X�9�h���TQߏt�gr����
}�<�#N��!5p+7�,WԔV�k+c�q�mu)ö��.==�yV5l�\�cV��yV7�{(�Z�h�j� ���9�Z�GQ�_vb\͗���[G��y����+��J��3<خn$�l�1��'���RQ���*�jZ��X����1�b>��6z����V����R:����fw���x3��[]�G\��w����y���e���v/��5"�6Y�Z�Q����*�g2�hB��̥Y6W�U¯rΪ��(��[-�-�nZ3V��Y3I�l�L�^��9��Vb6v��ؑ��sL0�C��,v|.����!�[���Yx�sMܲ�!(�(�u���^�nh�u�K���hv�.m�l�r?^����׋�|�8ױ����%t֘���+(�i�Nd��g��W z^�t�쇋K��UxѸ�9*�26Z��z�,�JT��K�z�VK�u4��N_�/�=��u���-n}��K9;�em�k�V���Խ/ё�o9뾮�:4�z�����1-#
�c���NQ4b.�Ȼ�l�[�U���D/��?c���k��
������v+�V`��U�ә��G+*봎�e�[vMA{�nPB
�8�)��J�b2�C؅c�Y���M��^�l���mO��XN�og<�$��vw+��ua�������B2ޮC>��3L�����[��-N�x��SvpUك���鋞��������^ɝ�������l�Oɩ(νL��4��
��1
'\���KzX�=y�[y��f5�^�^�o�no��2tֈ���ڥE�]l��}5-�������LU�&�a̔ж�}{pۆ�f%��Q,�lD=[{[j��e�xT�$[���v�V��nrC�ɾY[sF�T�1��'���W�(Ǽ��y~
��i����Өj�;j�ا���w��G_��g�ީ�ͯ;ъq��a,\U�;O
kLZ�e���ǘ]ϟ��ʹT[�
����XlT�Cn�6�4���+LAd�2Q�VqZ���b�\��b��:�3y�B�8����2�a~f�r�L�L]%��k2�����r6��쳚���<=ڛ���Z�xk_%4[,�i��V�J*Ki�j�1{,��ڝe������,M�Ms���O<
к�K�-g�����HΚ��0;yGwt��]o/Ӂuj�w��E�d8Wa][���lF�ۧw��z�U�{hb!Қ��+;B�]B����~���&��^5�ZŻ�j3Y��B���9�,7aB�s�[��;�v��}��}T��l�XM�sܟC��M�NA5��SZd���[^RV�);9��;E���b���«a��K�s��M3��ԭ2��^�hX���-yj���ִ��'�2�I��|��dNzJ2j1�����/v��ɠ�1%6�D�6����Z{�2M3n����;c�ձ�媥9Qx5�g��d�tfO&���=U~/�w����^Kˉ=��j�Xho�Tۤ[�=�����[o7-����g�Q4Щ=���(��A}'ybY�׳�6�}\��ۙ���ÕQIe�;���*N���)�S��C��|���n���)/VvFL3�����&��6b�Lę�e�K��y{�Qj/;�h��d�E�r�J�zr����kn���u}kqΕ��Ak��՚�䜷(]���0��)E�-�,ؘl
;,.̴+�6*�z�z�_�L�f�E
.�=�츏^u%9���gx�ޠ7i�"�%�r^�h�C��BP�t��V���0|�K��H 7)T�g6YQU�ɀJ坝���74d�\��*�{zcsVv-х�JN\�D+U��@m^S�")�Éwc�)���y�Ӫ���5[:����O.�k�T1�/��ﰥ����s�"[�{!˙��H���@�x�Ul��chŸ��P�ܰ�f�l��P,򮶸)��)�U�o]���`��VLLr=���O��ۙXe�5	tһ����Yݥۗ�q�Vj/�� v{VܷfԀ��f��xQ���N�]Zt:�����'�x�h�JL��F��$�X�o���t���1�)=N���i9�@V��W8��3�
	u���$:�t+������.w�����`���]�t�X�X4z�!�*��i
4��4�����C>̧v�K}k��R���R8�*�]Ze�؝J���\�.c��Ӯ_[\̾�;u0	-�bT#�U��p񥒷Y��m�9�b[x��2�ɲ��[Tt�V����6��9���z֊T/��XY�ٵI�7�RE��f�H�t~tc�	(m@k���ݗL������;6�v�Ֆd�Ng &�+WX˛|K���U#BTZVs���j��ő�gg-ݑ�1[O�=��A���n�"J�j2S�9�c��9\�E,-̠����lMr�	�8%dM7�L�8R�A�����y�%��n�=*=)!C��㼆�榹C��
�b�܃F�7X��Fk�ӯy	1m'D����Tƍ�7�Lh}>�yj�p���elwM��C�fVk�aGE��(v��X�31��%�[�@�D��w5��=*�f�����Zq��{��d�L���m-����Q�����<��^.��K[�Q]�}���æ�/�v�iCK�b7�'+�ٹLY���1s?`�V��\䳪�f7c�'5*�Y���f���;��,e� ^E�ʫ[v �������C��o����0�}B����a}�M\b��}\+�K��u1{|d�
��ɍ���Z�{�.%�eQ�[����IUa�~K;���ܢt�I�˼ޡ�R�;m�뺅v_sԫo��c��-��鷫z�k����Vf�jP������\4_%�hki����v�(�tg� 98��Fl����\dڙ�	˧vu��q-���:-�;@��X7ˬ�2��;��n��:��e��W��2�s����){��_n4�v��N���SF�|�U�3e�o/�P�:R�^��\��N:�2v��}�\�r9ym��Q�r�}�KJ(��O+�qVw��dT����YlmNu�7�Zi�*yv�;��L��f���%M�v�	�����C*Uނ��I��r��n+�ʘ�,<�����Q�*+/���k2E(�<x�u�q�"��v�Ȧ91����r* �����]0�N���������J�̻�J)�f �9�H̒���CD)��I`�uܦH�Js�6)LJ8��0;��(���4�� �".눢�n먔PB33Ra2is�˩�r�Q�Y���&�7w2I�����D�J0�1wpF;��]�e$HFG��"f�II;�j34� ɱFf4�a#H���,0Б`�;!�	���Qd%$��s�Rl�YdYac0̱I%��]�I0�fPgu� H��wtːd��st�-��α�4je��hK3&u�A;�@�u�Gw)y�c���;;���C��S�)d�슒I��!�I�,d��f1��sg]$b4����ؤ�iF��h�",�%}uqwK"���^3�K�u��O&��4
��.@�')���릠��^֐cM��:����(cЍe\���(3�8I߼��{�T�Z��kU���ې��&�L�eZ�*j6&am��2�K�}��giǓ�ﻫ|ggD�����	a6���-�Y[�WLl]�/W{	)����-���͆��gz���@Η-��57�,;l��֬�kG#i�vсEwp��sF ��r*5�����b�Z얆�:�)K�nd�8NDX�dJâ�e<m�������v�C����d�#�65%!:L��c�l+Jѹ�����W<����"����Q���H�:.�>�bM͞��vwO'�rE=�a��Zc�������2t��!o,4����w�!�w�����yf�'���Z;~�ד�z�,��L2�I������ݏu�b�w?M�^�ng��������`inYY�U��S&'�C�l-�1�Cfj��B��i��x��3�x�J%��E���+a�S��K|k����m�xL�٬u
��sy���n�ѡ	�)WP�� ���z�Gg�>ol+��e�z�����hSF|��;���;;����N�{˕>̧O�������y�ڃ4��]��*�mL�2�����q.��w�䡻y��9I߾�꯲yt9{��ۇ�ZF�V!��a����,�r�x�Q�RО�Զ�h�|���޲����_�]�r���mi��8s�%�mĵ���-@W��X1[���k�7j��m�"RM���bij�J6���m��5�w����P��}�#)V+9��#h���a���+E�S�\�\����6�?o-���>\�v��qP���lW74k6SL�UɌ�%����. �B�����s�E~{��]!v�)l�6T5��؃��JՉ�R�����M����|�uC�Y��F�&}�6^^�PͲ�ޭZ��jj0���òn����x؏�՛�XO�5��c�*��C͘Qs�͖���h�*f�yIm�#ij��v�MF��Ӕ�VbVw֎-Ln���uH�Z���m�=����*���h��O�r�bhf�A(��EmBՕ����M:Ǽ�`>�{N�j��I��@Q�
�h��w���O��Z����P7�i��c���.�Wf:k.Eյj}7r�̤�e�aU��n�wcy���GK�W@��˦���|��S����6��mB�0t�7�n��̑���6�����v�Vf^�ws�7�������6�˭���Df*m�F�ҫL�Rm�:m�-��<�@2��.��['�z�#����ȼ���=<~�n%�WM��ʴ�%^��R�HA�Ȫ+\���U&3wp���P�⼉Ƈ7>���hwHo��]�O��F��2��<�cm�B�ǧ��Y��O��;c��
ؠr=��i��if��ċ3���Pf%-Q����+�.Ģ��Х9ws{ ��66���~F���f�m���i�ߪ/{��Z'�'�*T_�B�mpvFL9��P�tK�@ӫb�n3Jm�Iى�PH&��^����T�u�ӾU���l��s5-��t��F�ĵ���j��1>6�D�$ث���h��04F`:76\�E7�x�3���\�Kn�˯�+:�Zx��g�~�f���|N�;Ȏ��c��O���M����S��U��V��8�)��|fg��(�J�%����ՠq��(]t�V�� >CGl�е�x���C1�_.4
�N�E��Z!ۚ�=k��4����}y���k��s��|m�v�B%S:�W�뫲��61��gv��B�(�T�ܩ�V2[nH�.t��7��
���j����m�_7��u(���s��vg�QrѼ.l���e�q�굈��͹��d�����cg�oڼ�3�+KG���B:��Q1�U[f��n`� ����3�jѮ�6�Im�Mf%[�h�m4�ݖg5z�J��g1�R��A%s���?RXgO{-�%��^���d���#5�Qv��Yf�]iN&�K��8[p[L��&���Uz�%u�ImyIX]]�+*�ٛ�Jw+Z�'��t>{�j9Dv�G����]U��bdq'��SC-�j�nVZ�cj����)̟i�|ga�m�S1�q��}�ȣ���y�t�N$��^蟩=V��A8��1��� ��հU'Ʋ/s�]��cM��/���g�Z����w
�aWcU��S*%�C����*,�j�W3��f�^����l6�>҉d�"̞��$��̢�uލ�/ku�E��7�L�Y�� �z`�A���N��e�2�K���O`�s���T߱��~��ѥ��{��B�\i��x/v�`�%p��8-ia��1`Y�-ݮ��Β��|Njj��3z��Ķ������P��N�U|��K&p���5�]ꉃ��*74buD���S'Mj���U�m�٫�-Oxx��B�z�H�t1���w�:k7��1&`�B%�L)�
mT,�P_$+:�f�U�x�bE�Hׄ��Jcmnr�o˔y�2�۳&u����◛�>��eԋI�֋y���a��e������ͳ=ڙֳ��ء�C��WL{Qu>�;�ݚ&��Khp&m���1GL��:�"�4".m3ԬU�8+J�T���?E�/�����&�cU�淪��0�R�az{��6}i��������U]�!�Sv^^�����>�-�ܞ�7�>uP��e���Z֛q�ܴ6iԢ�/C�gk�����}��Y��6�y�^�a��|2��e���.��[�g*M���o�O7W��/w����g��p�o��O�����/oS��ٮ�^��;N����A��v<r\�:�=���C9����h������ܠ��,�ڍ��"X�0ԞV�V0�H�ݬeGgWT���������q�V��F���̎�uz�<SU���j����~e��FQyїǟ諭����PFB�9봯#E�1��Ee1�I�\�ݠr9F����#u� G�c�Y-����4>�4�%��WLڭ��{�z�)JM���O�a���J�Y��[Y�U4x^%��m��rwh[��V`V����c�6ǘ���cLI�8����q����h�m�:Q$*Ĭ+��b�������e��9��x}Z��~�+_zf�4���w�����/��9V��TF��9�F�[�A[Y�Q:���d�?b�E�K��3��g��*�����^�5]��f�P�)6*b�ؚZ���mxJ�V��$^�D�|��������]�ifMm6队L�|�a���h��L7>��W�n�'���G�����}�-�k)��ěfͅ�q2�W&2���Uq@��8��T���ޡ�����{����Ge�����p�lA��b����Ћ����;vz���w��AJwt�X�ڈ�	٪�ǫ2a�(R*�}�}9���Wcͫ��#�j� ��1h�7�:��en�|���7cgF����۫�ܣn)[J��Z���o�ή�Lf*S���2���܇�W�U[�ʧ�����/�%r�v��'��Tb�^c��"�24R�Qb7&���j�u��ފCS�^ӏ�����mgW����ͭ�Ne�Z���jNH׸����g���~������hq���NH�"Z�qS�J���3
��k�2ׅ�����V�-YF/d�p�tZ�#jrX��{jQ��V+��qx���cPM{*�L��cz���N��(�;V�ۭ�A9��k	z�� G��h}N7V1�p	T�z����s߫��fr9N ���
-�����'��Cλ��Gu!��H������{�`���'�r�x���Q�5��g*�K^�׹3*%��R}��U�|���Ϣo�N���Gf���cz�Il��5����F�؟$��Jy1w��~�c랙������$W��yAS�J����F�Щ=P��J$�y:�;X��B��f����s>�@��n��w]�On`B^<��a@,��4��f��ҜR/�{Y&�:��S��D,�2�Y%��$�ŭr��b�=:,�\o�^g�V#���ӓE����9>AQ,<���k����J]��̾��K��
�ۗhPr�pHM��ͮ�3+�t�sK3�tf\M��Ф���%I�Z�/m�54j�L鍥���F��vY�}d�?Vw�mR���x�0m2�fI6*/����oY��U7��[��y�\�u�{�A�U�Z7nm]���'٪r�q2�v��Y[��L��f�J�n��&k1�
x��5�Rֻ�X|�9Z�<�>Db����nBWNQ���U5�O�u�2�Qg�Uc���/N��f�{]"/@����-s���/̞�aa)��Z��wF����C��R�wٱZSG�{���tO�J�^��w&zz��Km��e2W��G#i���w�#0��k�9�=a�k&=��t�=!�gO(RN(Z����$�5���6׹1s��h�7W��:�u������fi��M{*���]ZKm��WmslU��U2�������M�Rt�g�-4���:�^����Yt/�[OKw��+�;}�u�*���
nKuz��7�P��`_w]u#9w�eԽ��[��F��Ri��	��+nb�30��Y�I�cȡj�.ժa=��KA����̵����P�˺z_T�m��wj;��8f�P7{:����ꪠu��1��y�����y^�OIh�s'�a�n�D�>���:��z,4�M�e�-+MeT/=%zi,ؚ�YZ{�B�i��R}���4.��묤y�oN5�O�uE���Z�UKX��&��Y~b��Or�TK1�s;�ҩ��y��JiA�ie�g^W���0;���iD��*d�D�$���'����B���z'p�R,^��/³ء�Te�����
8	����סVEfh>����k�:�?MT��k�cNr�`�����f+4I�9e\��7��U<�!r��WzDN�^$�r�[Cj���m[>܉^�K��^뜮0w8�wg]ޭ�9G(�E�K2Qs��q0֓���ϡ]�2��5��3CT�$�>MZ��ks]a��S,�i񊚃X�Zڡ����^ڱQŷs���MsapI{<�j�;�Φg;5;�Ɵ��'藴�K�㩔�3��W]/ƺ2^�9���`:��J��]�/zۮ��׮�fp�L	��K)�n����bR�yh�j���]���j��5)e�}N���旈:��r��RL<t2#<%�4ٱс�&��z�jo�9w�|:��t���g�?���=���(K�	�g�m�~�����͖�:5�&������P�뙦��zf��
�R�p�Fճ��͖�0Yl�Zm�Z�N�W�ޜ�瑮��sc��#����t�fXq����6���0�g�[L��E�o�Y�N.�r��&��W,��LR��>�NS_f��O@єǷ�#�dQ	�n:Q�������j����S�F����1�H��1iW�S�:�ƭ�HXve2�ζ]6�ҥX��pu5��z�8��U��P���u{*d�5U���}��*䬾��o�^x�����w����N���[+3�m����c�3;������'���ro�(���F:Q�(����Pb��c%�F�]���H�C�Ь����%w�oR'ٸ.)�8�*�����BPZ��C(q~WZGk��Q��/m�Wηd]x�R��VA󶯔,VQ�~�ޞ�Om0΁�PI�=��o�k/oL��A$gl����RqFYݮ�}�s������B�}ǖk��c:���O7h�э|�ʷ�V���{MTL��ػ��z�!�Z�s[�K�H�@Y»drt?K��_
���ݳ�o�ۺ��vݥnAӗh=؎,G�oQS�9Z�of�)/�х7��Q�]���l�W��\;�����Zm��;���*�]̳�VN�(>��t�iYJ�a{���N�v���u����R��]+-i�"^٦U�k�G�I���B���3w�D��%vn�.���۱�6Cϳ&�	�\�Iq�Ԍn�w�b�`J�t8��h>�����t�����
]�U.����ǳ�LKu��̗-V��E��`��3Ռ#�0W<��7��g���Vd��}$���%��u�=�bp��_b��s�^�_W�^��H��ԺC�G��G(�/�r�Fi'm'���v�uĲ��qw���njd|v��	��[9atil��W��ɉ�qhtv�}�̡R��6��)��9�tgP���98�J]�(��@X���u( �-n%d�/��"ė*um�جڽ�3�]�@���x�hA�@)����b���t�t��7�N,K�����8�+$Վ=[Kz�ѻ��B����7��S4iꮬC�	��	,��]�[L_�v)�&��eh���i["���`o8�r<�xb�^4(fU�ɇ�*�׏d����7y�D7�v)�nǙ��ߞq�<v������|񗻌�d�V��Sԍ�q�r��5��@���,�;v���EQՒu�X5+)w,(�7Ď�"��3��e��)v�����R򙠣.6�\�;����#.�j�|��`�]¬�)�T;ͫ�X�j�,��-�s]�ipVT�o��ϗa�Z�r�*J=�u[��0�Wu��ӗ�-����f�͚:� c@����PL��ƭ�n<ǚ����܅s��Fn�1�d�{&�I�}�U��8ս��zõ)���Ǯ�GV���:"M�ӳ/�֯�;XD��;<��oqXa�SxT�k�sV�
�j�\[7(�n ��4\YyO��Ɉ�*J�+mK&�;B��!��}ڍ������ĄtMýA��y�dwo�Rw8�FKղ���A��x�pT�'w8R[3��N��7Ծt�eso�Qe���n.�5#����4i��7�SΨ���e�ҳ�`���|�C̞Sj+�Cs��XLy)0��r4�J]3&^e��2��58�Nt�h[>���In=���6vb����;n��j�t.�9�Q�s%�;���x�or]s��ȤN(�����v�f;��av��Շvԧ�e�V��GC+�Ӝ���]�u���p�q]��tQ�Ub:<듺=Wϩ�*r{�c������jc����f�������_ԁB�}@P	D�iED��s'9�N�r%E$̘5j"�D���X�e�PbQ\�Ah"���r���6��L`��AELJw]w\Ƥ�p�4lfcH^uɄ�]�cHf$BNtb�Q��I��:PIH�7�F�C4�,�a(�a2�@�乹��2��	�F4L�6D5�)��
e	2\�:t��.��`2F�T��	��l[���n],�#r�x�bH@�f^vw,r�
L�s���&�`�CPa�<�г,2��Rx�"X�r�CAH&6���6B�����J4rܒ��BP�I1���3 rB�fiӃ�e�cg���Jpm���%Y},�س�w�Qݝ�2W;A6���l�C!��y[��p��Hd��Eb&^2�+ۉ �;1,�JRkDS,ɵR��+[$M��i�¨VT�s�xs\����n7&�n��6�D�I�jz�Z-�-&����h��Z����^j`ݺ�x�nn$�l,8�AfW&���r�E=�w���t�A�3/ĒsSaamGZ�<��A�s�*�p빱�a�k���I�-:��wϏB7��Թ���*����s���8���뚺��zyBt�K�n{L���~{���Y���-ʞSix�|l��Px+�z�����|YYX�j�e��,�V�.M��L�a�n51�9�9ޏ�
���C :oz��.}q�FB�e���m0��ZBQE��^��ҍB��5�վBc��lGp�U������֜f5�J��%u�L�J+)��OT��!��|��%�<U߭԰Z\p����g%]6�G-1� )������3����V�zԓn��N»+:��Y����ҍ�Z�lkn�3�q�8�H��o��ꙇ!��3�[3��[�v�S�Ҥ��r��XX����t�z~����JחL�ڰ�)��V.O �)P�y����lՖ��om
՟>[Y�n�g'�9 丛�Y�ս&ۜ�a��X�L3�8%��&}nrR�󓻷FӬS�r�^25f:l��D�ƫ4^�)/,T:�i�lZa[K�iFhi9�E�R�7�x��#^`�eT3�'��)O>1g� ��a=0sZ���t@�i���p����U91�
t�4�-		 �'��*�I�Q,�/���l,�4�ͥZ��w74z�q��\M������PH��^�
ji��=;�ūƃ�fbM��{���UM��9�a���Е����n+TI��L�|���{~��,pHVuo�j5�lJ�5���ȯ�����i��֫�S��N�X���{ K���2�{���O�sRֻ9�}�ޣT&୰c@�ķ_.�j���w6��6��	��˕Ԣ�ǘ]����2�Q}R�\���Ҥ��&BGm�ZlL��X�b4�ugJ����V��1����Mٙ�ߝ�e/?m$�Q�+/�n��8��ˍ*[OOt�r�fv���6� 7~���sl�g]L�����y�;o��2�PM=�^V�.k��Y8q� �����p��[]{���X���ۗ��0&M���DiFe��2z��Q��9���b�GK��{S=<��X|��)���G#Te=4ƫ\[�;��o{�8C�QȾ9�-k���^�d�5iԡJX���m�[��a�M]�ܙ/p�幦�a����k��NA4͏�K��$.m�h	��;g̎^��Q��C)����Zj�f�Zh�9[�uSd;��R)N��陬���LrU��e��2}���dK��Y*�V���Ŕn%���4�Zj�������]a��gl���,������`�7�0���rmb�H�
�aWcY���S�������ލ2ݍ��H��/������ab������-�A-		#�T�j��[�*�e#�����괹?���(�9qef�>'TK�%o3:��u�9&�J3��(٧6_��j[#&<�.%�
��W���ֹuZ�kJm,�!�y7_�.9���&��Y����v�٭�SiK��!�
��ݞP�ݭY;�k����M6�\}�R�󝯾������u"W^f15���ޮ��(��Z�/�.n�z�gч	�˔.���a+JK�`�u�[�4�wix��Kfm]���[e)5�b�rؚ�U(4�V��>���6��\*Z�88�{��,�9��-x�eH��d���E���5|'k�w�9<��3�/���eȨs��MLN�ͅ�q6�e��*�AZs��ZF�fv���Ȏ/l�	o��n=ȭm/P;��fs�S�<_��/���O�xp3o!���s���[r,�$�ؾL�EϠ��Z٫N��Z���,;�Nɇ��E`��'��Uח�֎F��۟99V���7:�6תjQ�<�����ɧ��z�4�vz��C���s���!�w�w&�R{N�i)�C�(��X�.�ȹM����TR[JJ�1ZsjeەAЯ�ӳHWϧnNF{�鱕����/Df*fڅ�e+����Zc���bҡ��X��=�C^I����d���r�0�᚜-Xh�Ug�U����'�P-��ޱS6�9]�)�l�oiQF��ׁ�R�\�A1�u�O*F��3՘�67]4��7�:#�غ��V�T�=���ےE�uV�g0�g>t;*��v@����.�ٹ�s�
�V�uOh��ٴ�(}� x���ّ�[��9Vi��.>�P\Vco�l܉o�h��~����{�=2_<�����4�/�f�ֈP^w%)�4��zU3q��p�`����Ѡr6�m(���d��w��N)��WTI^v'ȫi�Q,b냾�lO�����=&��X+q���[iD��*d��_w���S��i��4{<�M {Af�3gT:v,��M�f I،�P�)6*b��D�j�BV�s`����0�#�.��h��Ƶq�ɣ^�Sm2�I0�OV�E����Si9q4��k��F��4YXn&�f��8�D�����LBU�QLullJ��Tj��X\xQ�|���]b���\yҵ.����6h�(����/���T���K�ڮ�X�Ei:��|=|�V�o�����07d���b�LF��Ê ��]�};ŹS�o��c�d���+�e`Ү��l�������^l��œA�g��9n��*��Y�
���{\;"��m�,ٶ�([��
��O�<���:���)�
Z�),^Gȫ��_#|�A����T^���s�L呝}o������st�V�l�:W.��V\(N��
�F���x�$�cD�Zm�[��f�MF	�h+2��-h�m4��e<t�|j`�2sѐ��R��>�nuzR��ue�(�b��Z�X��F�cV۾E
{�SF&�wS bf|���ۈ:h�ؔ�J�2�(�ɀ� �Ut �Ne�
c*%N�t1�-3�re��U1�q.J�L��m篢;�ǻ˓��\�q�-m2��2��Fx����hss씡��y������S:�SV��G�����[Y��ò|�
B�䬷:fm5-�%$�E�Z6��L^�;�*�l+�,�{uK���G�j�aݶ�n�y{֞.�f�}�I����g�u`����u��C1T�LB��-��MܻY�ܩ�����6��g�Q>��Vnh2����IA ����;|R�Î �L��cض��a��I�l���#��K�T~^5]ݹ�r�{<+�϶��Z��l��P�M���Ypӡ�=f�H�K��6��/t�Z���Z�:�5�;:���Z�H�+nU�|���c����W	�;)\Úy+w6�aݰh��db[3+S�c�xs����d?�ɩ�zה�m�vE)��3y��c�{���T��]��V�_׼��EVr�/�j��Y�#�})uw>e����n�]����D�)/��d�o/=Cj{l]�S��]b��9�R�=���6��᥵6���)��r����J��<��Y���َ�R�q<^��¢o"�B!m/Q�?9�:�vy�����k���u��l:��u=��]ڻ�����w���M	��ZjӢ�ajj0���̯%z��X�L�eV#�	�ҋ��ؑz�T������[V�N�ʒ�5��J��w.�N��Pz���K0��x�~��!�e��9�`�e�l�m2� �	K�QF���|���m����N~�����v��9�:�3�?��>�&a֜z"�Lc[������]���Ud:j��adr��zrW�����﷑�5Ctsk���R�˖;T�1SՁ�|�~���r�D�I�+On���T�O��X��.b_a3sx�f��ޭ����qeCeJk���u�l�h5��v�g;���t�orb͒q�pL?�q=�vM�v��5qa�[{�]�x�� ٸ+�����ֺ���iV�n��f������<�b6>��,�$�V�G#Q��eN[2���=$��q��6�c?xU43ġ�g��*gH�`�v5Z{�S*$�3Sw59>e��?�p??�Ϯ����s��tD�ΔM�*d�@��eaP���M]��0�̕�2i�u^��
Y���vZt������ֹܶ}����/��_��q3[��eM~b�	1J'\-l�r� ����_��;ۅ݂�zƥ�l��oۛ˽y)&�C��kmR��	Z�)��wM�k���iaYC�	�z�ţ1�\6d��6霪���uZu�b��1S�\�=f+m%�y{�O���-�+[T��sy}Ng�c��R�Q�֢��85�#W�6��N�=�2z��V_���V��<���+[K��a͈84�G-ݚ����=	+��+��|^����b5�����qmg!�Zt�݅���jmn�(�[�V%mu���ފC���d�i�����r�pZmL�P�
V�\����۝���W��z����s�zhC	�+@:���oq�Ri�ڒ�iU�q�qu�/8f�=��r���M�Ѫ�]�ۘi�'�s!ŬK� LoR]C(v#��[y��U�XoDn�.��jOT�[��)��
��ځ��q\�R���w	��-u�x̎Xq��t�9��Ճӝ�h?`U�G<�wc�ݑ�ۜL�顨�(���+(�l�͸4Ӡly�(��D�������|�އ�w:���)]{#t֘�VQ�I�\�[��-���/wH���2f�-R�����J��V�߱5��^�����@�`�����'6xt8���9F�u*=0�<���hwHj��1�bw��o�Uf�5�9Bj�{�2�|T:�c�}�	�C��b�����݀r����N��^+��B�#lؖd�����b�l�����0r�a�Ɍy'#V�X�8�Q��1�
ZOH*بB��(�k���;Bz�����G30�Bh[q>�q�B�����b���D�j��Ř2��cyy���;0�}h��H�qf��N��%$�'T^j�����ȸ�E�I�o�"�� r�Î�Gn�YDa�.�l�[c�(f��{��N�mz���;��A��z��go�=f�5�w�١S�r�P!�7�2e$���d9Ir�:�k�v���N;�1ŵ�L��xS."WB������_]�Dy��y�ٚ&��er�����ե��Hr�\ej����5����~��Ğ��}4���b����&k1���jO��-P��.��J{].�n���<�m�ho9��16.�Ǵ�'���}���k�����Ҿ��ᠺ��E����fw&�f���ܳ�ɮU�勺���d񒗊�k����Xsdξ�N	�R'r�/�ntO����j��b�==S��씻ٓ�{9�~�Z��[�М�w��eO	��KC��Lv|��m�Ӥ#�z��=�m`<iHo��=��If��:��^��<B�b	zi��U��+�����n%�~��x���`{�N{�Z����6�f�cnc��9wu,�����*ixI�b<��e4�%]��<�b��x�z��C��_T�T_x����fWuW��p꼠 TKC��á'��c���C�F��6n�����.���/���A��;��ȳ�ڑ�MW�2%��#O�@j��}�c��FI��g��J�f7w�$���^o�l`X���)��X��`�km���r�R��)Vu��ç�Qէb�"�5�w���
�|ꠢ��ˡk�}O��Z
���\�е�'��%E��f �ɑ�ަ�M��H���#��9x�p�͍��.�i���ھ��#о�ahyxNؙ������I��p���(��
�v.�y{cr�[�'[,���]�+�A3�(�-�b� �uÞ���IG���1Y*�
1�v6��Q���'o#��ō�,�Ro4k��m{R��kgmt��G.;����Wul,�V��W���ٲS��:�*�b����q;��/��mŗA�-�Ǎ�q]��P�6"�+�G3�Ʈ��0�E�a��1�5!wne�Y��é��}��\(i2&��iq��W�� �֣�Ac&��NWk_fY�L�t{mN�\�ڝ7(���І-�y�9�բ�@o,�ڗ�5�;���)�=*�>��[M����A��ѼG���n��ݺ����Kږ�3��b�O�f�j�I��E[�N��ж�e��z�6��;:�|X6�Mg��}D��܄�֕ F�5�s8��R|�B�5JN����ݲB�����(V|r�[@2��:t���=��{�b˙ҁ����٩�x*&�F*^,���9�1�\e'�9G������aW|ܭ|��wYM�ֱ�qp�x�LcuI'P�]lU��W����,�K�e U4ŕ�-�d)Y=۷��o�S%�2o�v�|F�ЬJ&
]QAr����e�C^pw�Rf�}t�����nlN
8E+�d��-�ٕ�2�!'wj��a;�J�4<V�Y�z�;s�Y��L�la�M�c���0ʾ�Ү��������b��u{��¯�:���r��s��b��<�ne���$d�7�6F)f���]�ɬ�\�<�
���	G.`�0����D�q5ݮ��cp-`�K�����Mܸٸ����,�ó-��t���(�B lv9���o�1]WǶ�MM�]�v)�����U��.��rvq�@�h��yTU��%K�ݼJ�*q��ƥά�Z[��VLXp@K���c���VO���e.6u}k��c�D�cQ]�� �߀�Yfe^^3@f��t��~�iCf	s�6
�8��ʕ�R5�-^2xe�;
�)���ac� c��9V=�#o6]7E����wws�j���u��_ֱ�[*���:�����ǭj����\�6����R��ܩ�zSÌ�y6�'T��qd�5������[)�;z<��g�$˒+��*>�$:�vpF@���,гC{!�1��+Z�w\�m��M�u��������+1P}��L�����3��Z��L�xl�6;��s�8.��N��g����)Nt�Ԟ�Ю���2g-���U>u��1|ᭂ����\@:��N̐)yD�|V�c��yFNc���5���v�U (P*�
@P�wv��GI#QH�&d�����i4	��IJM��'��"wp�I;�2Cd��y�K�����ႉ�9v,�$�Lh�M5+�E�w-�;�MI1 y�D�ȼvP��뢅���4`�����!bsn��\�I.�a%ݷ]��x�/��$���㲉a�w<��F�4�Ć s��;r$��wp���<]M�����wH�� ��ǎFF%���☀�5ݹI�%w ��#u9ݠ&X��I;�F��;���,$����9��<��]���5�;�F��*I�P4��@ӕ���1��+�f�1���.�ې�m9ҒŮ�v��U��m�'���64']$�s��>!�x���Dܴ��q�)�_j�;}v��ѿK/��ec@����]-����1ͧ�<O�i��"Ӻ�yla+��)�� �1pTc�ֲ�V�ꚩx���"�NQ��Z7�#�r��}��G
fH�H���[s��]ҟ���Eњ�F�D:��:���i�2�^P�g1�]s��2�9�<2Jj\�5���ƫH�m��rx<�i�m��FW������3��Pn|:�5vi�����}�B�;��M��|�8r��f;�Z�z h�S�m��!���e_��J��cb�.��31�4�')2�i˽�c�y�]m2�1+]����y�<#o�q���_<㯜=��G���)�j��k��9�ӹg1��t�Kক��k��d-��V���j{e�#vٙmg;VveN��-a��-�W\�k�7B)�j��c|���6sҠ9f���8�0*g��约���-�R#)�J��2ƯH3�ӵ|�3cܤ�N�|f��8��4��ˤع���:�,�=�%���b�i(�G[e����;�bv=��n*g��P��(ҝ�3T����t�r��]c�k��g�p����}��[�	ƫ�,�c���+���c�Ƿ])���:�0��Oզ��K�-4(�^��ͮ��2ȬU���ɒ���]L�Ɣ���r��ڪ�T�,�J�5E���*������p�_��Ժ`Sז̠����0����;��w\m�lu��M�c���Q��|5Z>�^\	<�-��ѨJt��F�c�����Ӱ�s�6����i��v=�o@�Z��>�7a�[}����!>�p
�<h�f G�[j\����_�?x9݆����-Z�^���Vu"���1�����z�;+s�3ӑrj��B��5���ۀ��*��K:��&�:s�Gʐ[<0���z��h�M9��&��C���$R�iN:���i�x�~f�	�D9S��.��/�c�n��R��%ߪ�U��}��7z�&uhi.=z���rI���2Oi�$a���&�#�mTZ�eDnhQ�^�'cg]Eڟ]�]�;������S�շ<�ߠr�7T��J���ْ�h��Sج*�<ͣ�y��}Y^T��MO̙���{e�U��~���F��(�m��RY�1Ğ�*/�Q��ر�Mq-���[�W{ٝ4�:V�	�d,yc�t�~'���c�h�����OQ�4j1�'Z�׫�A�ۢLJ�s�q�睹�a�I����ArVD��_�ȳ���V���N�wF�`U���6�ި���ƍKV!�� T-2e��7�Œ�ڱV�nJ�/��ou!��Hf
��}3����pȈ��0xΘ�G�����>�45m��6�Ŧ-Xu
z͊��d�\��캫_��ke� �_lO<�t�c���fJ�B"��7�O�U�_�@w̦xn�n�:^OB�n���3���Sǡ8��1���v�݇�T�[�ͨ���]!~�:l��3�/TuB�Vj\�k�(k(ӌ1/��$4�~�ہ�q��N.![\h�W:9��칗�~�z�:�����(z��2����OF�{��b��@�����]7s��-���Ю�;E�ws>�@ȈЗ�D2қ甧2��a�+��krS=��
�/Υ�tw9��M�j&�ז�ǔ��0��хQ;`
Z�h�z���=�S:)�c��򸐦��u��m��(e�t��Mܩ�o�'9ۛ;��t�ڗnm��UZ��ī���z��>�����I�b=j���M	u`�=���6�}�F�`\c�H���{���l���׌�;�����)_`��^X�m4�BFȝ�s��+�3�Q��X�k�|[1�Z��&�L�B Q��5�Җ6�K;-rݍ-�Ӭ��b�)��F�z�X��a��h_vѬ�3;<�>Ѿ��L\���*ב����̕�ʄ�k�7�p��\�� ˧�^�+U.K�����<���5��i�=\���Zŀ\�:�_'NZ�}Q΃xS�ڴG}mZ�t���>m>�ӳwZ�k�m���������~���۫�iy�\��µI�$�ք`�.�+��Ù1\H�Z_F0)�f�g_om4k��%�M2^��`(橒+���˻�Z�c�Ste��|�[��l�
-<���y�V����S2F�]������\~���C�|@�&-<���a�s�&�;F�
���(��V%��"��;Uabz�E,�1^���Z}���0�g�,�M&�q��d�����
��g�vZ�Ә�.��oͲ�	�e]!~�3��e]�'Ǧ���f7"��o��&����G�.E߷�;䇱��ϙ,����X�o�������
�h�-�{U{�*�v��k����y�xF�eX�.��|�)������73��ҷ-�=��tZ��#�Ѯ��oZ�M֦$�jzu9�]��ߘ���Z�ɍ���^�B����G������Yv1F�'!�Ք������`�����O]6�ujv�g-�.�����!�E$i M(w�����\�qziP�ǁ� ��:�M���7=$v�q{R��F��� �5EL��Vt�i��g�➒�����g&)Kz����t�� +h�(D �m�#R�5bi�u���l�ŠtN�^h:d�|�U����QPe�2�
��ׁdkM�pp���&Ku)r�� �Vy[ٔȩ%���q��^pu)�a㕹�Ǳna��L�a��ˤϨ�'A�.��K�?�]HA_��U�f�h�|�v���9{x�V_e r�е��nHV6��r��Yᵀ��:O�A���k�7e��I�����zjk�ߖ��y�צ�3;�xq�� 
����t$�k��fn��unũ�4�u���SM4.�^�E�|e�1���:�eOM'��9��8.� {Z�r-��cJ�eWz��0a�!	`���΅p��v��e>7��5ۨ��ꙑ_rJx�R~#:�:c8�f���l�[TH�OF���Nl�[�pB���?=�DZwW�yl�m(ۊk���>���4����R��p�>˵�v�K�F�m���tӄ+��(�~���Ţ����]�U[m>q���Xz=Poz�:	/N�
'�]��s��e�'{+�g7T:U-m�w�:���Wg.9K������~��#8�����3��F�é5vk�z��9���9��w2�DLUoe��{���_�j镣�Z�����_T�~�\��"��'M�ç�X��c�1��a��VvN���s��*oz��U���j�sS������z�+�״I�>���cW��ͧr��>d�\��k�����4'�a˷����FR����4��TɧQ�o��&�J�ޢ��E]dyj��d�}|ź�"�(��)��L��͝��X���s�e��+3��lW4�{l��ﾭǦ�����#7�N�Z_D��y*i����.,*��|ӱ��^��#�u�l�������NWD�kq�fo�ɩ�4�=��?%T��&��o���O�Ӓ��YTC�c<z�[)��Ik�I[��k�	��Q��E[��*����Q�;��Q&;KMB��0ɑ��P;'A[2�sw��d���*'*[
t!��9DSw,�\��}ht^Y��*��qz�L
u%�'E��
�ـ�Æ5������~���㟭gSw�Q�
���ظu^PC��}�q�M��©Z'������Ѧ�'�q?<�bU���9�:l�	����-�tNs�kЄ����d�yB�U�u���t����OCSLG.�V�ס*#�Yԋ�8��ݝMS�I�7��/m0�X{3LѲ�uqя���p6���8��<bm���s�G�R�~����u޸L��5Wn�k��[��X��OU�T񯴈`������=�߾��9��
+� ��EkOC�8�"3Fj�mΫr�3ml��{č��EeY�c�BR�R����X��-b��<hExNS�\
�ݥ,����|�橐�WcV���+�3ٸ��㕧�V��tz�teÖ�2�w���4��B����ή�	Y�>%���Y�f
ܚ ��*	8/r��Ė�9[��Xz߹t���q�&���$���F=��#��\Z�玆A��\Z��w�W��6�1ή��\ւؖ �߇+CuL�J����/f��%�l���Et[/��vp�;6�>E���ߔu}��H�m�2Qm���B�1�d/���B,j�[h
|�Gv�\��v6z�i�O��rxN?[���F7]V�c�ѯ9�r��.��fh�߳2�hqEr�f�Yۺu�	����s�N�8�#���܎M�Ua1�LV��~y)��i⾢���mC�9r���0�ג��ސM����_/'��M�u� �~��|ߦ�~���,b���A{�i��Z?�������;����J�qzmqպ����λ�'���������z�'��;㔩<�DpŰWd�}��E��Gv���z���(ڄ��*W� lo�Z�#9�w-�E�cTF?Hz?J��sm<i�m�m�M�0�F��D L�h��GI��������l���;%3����E�����M�*n��E�>��|�wa/��*���Dl����^�ǉ���5E;���\v�qOFL�����"G�m4����j�T`+��m۷F����3�Nw"^V�s�m��{��˘�M��n�����GT*&�3f��e��d�v��Gj`G�0���:u��г3���{�m�+g�;W�JI�p��X�-h��EE�����u��{�҆_��'��Tݲ�
�:��[�p̤��3׎�îc�������1��'�� ��+W�EB]X/ǲy9�N��_�_Ym��Y\�z��z�U��l6�9�̜0(;k
�܀u�Y��*6�T*
��)�M]��ۼ����.�£;�7gL�Bn9�.k���F=��d���؇��u�'kH���\�/�Z�����{���[!�|Cn�3L�䔞��� �'ew�����,��?��ٚ�`h�=��y��eLQ���.�.������X˦��R���'E�ą3��=	[��μ����*
&�YB�������cDwv��okE�9p1�����b��(l�O����u�.Z]�����i�9X.Tv<�B'j�!lOUH�,�1|5^��\�.,��� ���q��a:��Шe����:.����?nµr�(��Ml����?S�Os�ڗ�?�ˈ�h2��j�,�̋�^�+����]�vB�zi�l���90q��0����+^�E�ǳ�Ū`Yj�J�Ӱ�ι�r��n��MTi��m;��u�Z7/��Y�#Y{{RU�k�N�·��X�S-�o��`�i�qvݩM񙄾��(��c��yP����p��#�N�}h���^+�i'0�fh77G9[���
";�����zg�m�;oyu�K�����f�V�����SMI0�>��uF�v����~��'}z�?0��ƛ�LI��ON�9��LI�����%����[�w�5t���5xA��Y���2�)��#���������������4��n�ujv��s]��V��7+g�SZ]��gO�P�8�c�`&�\%tw>�6ޮ�p����T��-L�t��؜N�+I�0�������鯡)c{�ޤ8&��fDm-�{���1���; v��C��M�
�m�'���Լ6��?e^ixI��1}g��Ro�-��V�7<�,��5�\��}]�e@�m� -z�3)���u�l\:�2�Q0�x%,6�KH3�TWdKa��$͒lm�a~ix��s]rӰ���/��qo���S4��x��"9�3��v����9f��u����aw,a��;��^|sgB�]I;[|_��.nɯ�uu	�3"���N�Qъ-b�kr�α��K�.ԑy_	$F$SJ����ͧ
�5�~�O�}i�.�˞����%��=��=��77HN!�0"��/-+m,��b��)�oi��T�u��O�p����*0#&�;@���[̕[��jr��A}�h�L�<�� U�v3r�Wr��,<���a�bV��e�.*F-c�$q�$���<��[ŗ�u�rZ������(~����4�����[j��3���d!�L�CR5R/���g۰�e�%���w=�x@a���5K�=.X�9zj �(=�~29�-�eA���ҶMd�G6U�,��#qD˛P�n��5�ی�oG�sFg6��h��u|��4��+���/�P��x��nMs��_��H���sR��UV���������uH��)|��ސ����ã�=df6fW.Yy���Z�]|��6k�-�~���j��Ǚ���m�3�6�V��}�8�|�>G������+��)�=���-��d���OBw�od "��3%[Sթ�tO92�%:�
����}�Ĭس*�{9���ʞt-��;*�]��|���6Jʒa�=lF+wb��q1�z�4������}kE}o���(��c���P�E�T �xd��s���J��rk��@1�D�����8m��"��e@>��N�{J�:��zL٨}�w���n��-�	��c}Z~6�e��GvO#g)�!_��êe;��� ��8q�k��y���N��ވ��P,�`�"���C�՛Y�p���GQ[!YbP�z�gb�ch&7�YYCC�#��V*�Dp�x�g^l��l1äk�:j�EF�V�;\s�i�ũ�u��i�ZF,�� a��j�97&wvT�����8���0�[QI��zQ��3��3Cto����|��Y��?9zά]�Y��Y|�3sx��k&;����w���8$���ˠ��t�R�E�2�.�7Pݤ�̂n+��]B���c��n��7KЗ�)ۀ�vA���e���l�Me=�ꋛ8���A������.i�:R��2�6�JBb�t�죣��~���iu�|�w`'ot�Q�����`�e�G��g8���h{��v1H�,Z��G;6���Ӆ�;����g�L-dN���4���4Z�:����c�/��=m�^�(���s��T�Q�s�;/�o�uH"i�d�s�t�&V�ͧ��#�nV��qvSv��R���ѧ�
{6%��r�Ϩq���m����-Z���^�KuJR������6��.hD��r�m	q��̹J��W�_��1Kn|��s��4�B�����w2�"���z����Sdؐ�M��qڬ�{�$Z�n�r���nd�d�Y:�v����읚�0�s�r�ztNL��MQ���QZf������Z�%�Ƀ�S:���{�VR��w��l ����M��f������1 r�h���^�n�ѹ2�֤%N����s�@٫�
�x��j�j�;�+Q�1pW��)������gt'������VQ�
Qy͐�;���L>�.�=��K��N�E�Â�1�3�^��VN�.���d%q��'@�V�F�b�p�M�Z��K �lM��n�zfD.�{�o�Ս�*&)��=u�|��RF�u�M���7��i�k���j'�t�no7n�s��7Q9X3C�ӽ34�$��e�<D]:�����|��0�u�S�$�4�����V*��;�z�BA��*j�=#��c��'ks�շ�~X��&�O�u����=�������L�}oUds[���P<s�v]�zU�s,5j��yڃ�0Z�32v/���C	 N�Fd�����NH�b9|�=/j�a�-�m[kiB�]y�����P|�G���ٹJ�����RL}E��@ɑm㣱_d�.�:%��5!�)�&�v�cw:�bĸd�m�Q]�MsZ뽓�^��Ɉ3X�-D��HD��_R{���aY�f��1��4;/e�,w;�V�ut�pL:vn��r<p���{���T�W=��\s��lwa�]���V9̝��˻�|D��#.�����U������r�c�����wa��������,����`��0t�<�;����J�[�&ڊ��7�͂�9���oGU���T[�c���8�ps�S�)o��f:��~�f�h.��{��s�t1�64>�{�����ߟ�����H��h���A��!EE2S,;��x
w^8��;]�Gu����A4$��໶�a1�F�:�!K��Ļ�4S*)�"MN\D�R��i22K��2�:��G��w#wF�b!���(�;�Q�wu��y\"̘&5�r1���%%:扐��uy湆�7#gu�9͓��ם�4�yۤ�O;��2AI�r������:�x��;�p����<�	�F�]ԕЩ�'��$�3��pֳ���1����*K�R��PԾ��v��W'��ݪ���W�˥MY����Zk>l��#6��{��X�v=�z:׶΀�k��-����b��d�]Yf��^q{�n�<������j���/����oBTF+:�}��}��ц�\��Y�b!�n���笻[�����xc��p%��n�������:�P�c�ĩa��%e���ӎ�;�5ᦌzUJ�k�ba9�:� �zv^�.��-�23�n�+��M�����ͫ��y[�s�wW�x��黚�*%��&��MMi�{MA#�{F��|�[�%��v2�1�om[�a�\�߫8Kd�t�.�!�۞x�~
p	n�Jf�a��C�}�ݚ�{�-P��g����Ks0�h����z�X󺲛��*�zY���� �B ^tq�Ǧ�J��o�����r�Q]��ނ�i���;#�˞���G^���p�5�= �7H]3|�Wl��Ѯ�7(+.b�TW=<� O?���Cѯ�pO����.��c���oH=���z���,\���*���}�t�}�wFa����s��ң�3d�z붐M0���w�4��|u�݀��G+�a�9ܙN��U
��yH�'0{X�M��ienooT��m����tW� tyd��p��
��N�5�FS����sZ�h�2�i ����1�d��-�A.��Y�GA��[��Pԯ��B�$fM8&$�˂�?6���oD�&7�|6߮��>'޸�1�+��GT/%f��w9Zua��n�ݫ�;����]���A�
#��]�A��DSg)�s~��r2�![���e�Z�%\�'�������Ѹ�r�@f��-s�Cg}	�Fm�-�)�T�9F��M�ף�2C`���(�3�%��gLGl53O@*)lO:�~�ֺ����tw9��Mڞ(��!�??aW~�sY���ʊ��H:���B�0d�f��*-\HSM���m��C-��'���F�3�\k�TD�f�y���0�o�g��\t���8��HE�q�S$�V��hK�hke�w	����:ܫ39�>w�����$F=wWSu�ۘ�N/�!Ґ��2��F��N�k�EC�UNh�:o.�OE�Yήx��N&�vԋ��UpU�)s_q >�HǇJXIj��͛x��v�p�����8��b�_m�Q�����al�j���mՁM/2�9%'�j��";��@�16�s��õ�	�䉩�σ/���m�Q�ښ;��,�����U��i�cܿ;&�Ưne���X�����OoCa)�;0����t�AU�7��/�-l�mpt��f�J;vkxt}ӭ���^�Z��YU� B��9Mͮ�c���f��^ �erk:����2�kњ]I�ʉ��kk2Pg"�����
C,�;&�Ӗ����ͻ�;���{Y���(k�����a~&�s�w��ԍT�QK���G0ޣu�۝��!u����櫚���^�5\�
��ϴ�p�V���y�B��U�	��	���h��;��[���W'����nVӏM��,'z���xT2�vc���٨�z��F.K�ɭ*ws8��ÝWw�qٞ/l��s�vM;�6�^\��oHw��{\fC-f��.�v�M3"c�e�x3�V'��;}�O`���@�B�}*x}���V뜗�0�0�fy��(����E���������f�d�=}�j#W'�o��LI��峢�cG(�=0�Vh�ћw�n��s�%���tk���O�~1M��8��=G������9=t۹ou��B:Hl���n��R�ڞ�ɧ�.Cƺ1^��Y�D�7�uL�C���4�=�#OJ.V�mwnk�Ua���n&z:U銆��Y�$�0􃲆����1��WRFC?��%�U�q�ݹ�W[�3�������R�jnHW�0���������2�xI�)�^s�HB򰽟��D�:[�!]!0֊���*�=�OY�_��G�3�y�M�,��Uز�G�EM���}�5�u(]�r�c|�%8���3��u�cp�{i(�>�um�e�F���'�N�=�m��T�%�=��ʱ��Ƭ��x�r='L>Ř9S�'��SK�����9F�t�������ͯP�8T(} �\u�;�O̯��+�ͭ��p#Yh�u�~7�M5	Q.�9�>]kݝP2����2��|�B��{I��ۄ��DP��`�.�'C�y9��:�I�3��rq�v����b�*rxEsŅB��~�T��e��Xg��҂U���~[���Nl�Z�Q�[�~s!�#e�$��c��Nh���;*.ur��e�����%��GK�K��4�t���\^�����c�7}U[�6�'r��-rzl�R����h�i�^����Ob�>G���k(RR�3��qW�J���Ѷ_�n�C|�����n�_��OE�sF ��������)O�1h�ܚ�}w.�#�^a�5j�;�uX}�c@4���(F߻�F�)|��ސ�Y�3`.���m��U�6/._)�&�Y�r�e���Ok���i<�����ո�ؐ���K���V^�9��v�_����2�20*��|&9�+���B��V������C^d	�&�fU���31����Tz=�!��G�e�
����k�s3�<C�����N��y���+���fx����^BįW]Jy��ի�qY]�[ޗ-J���ɬ{j�(Ƒ�RWn�YN}�y�|8�3�]K�$���X n�S���noI`����7��vλ��B����+��Я4�N=S��L~�ρ]t��uXo����S�r�
a͓<�7T��{��"������=���=��e�zzd�4�{5J~'+1;�sW��)��Q�k[�p��f税���YP�Awr���<d�r�Ԑi�gެ�S������F�c5�3�h��s���󩻌_����e7D+���U�;���mU5�mgwz*�P+Te)�s
Z�}ޕ�T_u;8�g�����e����i�qc�7:��Qi��/��p}�A�%����-Z��I4��E���1�8k8�ڡ���g�_�ra��mx��;̠5Pt�	��16���c�Z8\w*Cu�f�4t>�uIuH�}�1Ty�3��]�M��]M*!9��  �l�˭~���FL`�瘥&�1�^vms�s���~kI~����[s`d�?D�$���� ��{F�E-�w��)�o'�4�q�;�|t�n�$k��t��|���`� �wUpu=0��!��e#��K�9U�t�(d��)� ܷF�s����nH�I�6�h�Y�����Nԑ�P_{����)>�Z������`3�3�imlo�h�9�Ҵ�*�-��o�����a�2<�� ���r�UCQt��W�i��a�6�R�M\��	|Al̳��\vp���;���/�g�������5�����wQ�ܒ=㬔\Cm��-���Y��ic]��n����2d��~1xt�r=��?c���{k���D�V�Z�i�{�L������ם���:$���7o�Ts,���0�������ۑŲ�!zg��ZV�G	�9��r.�+xj�n؞y�fΦ�zeו>8�'��3T	�1���xit�7V� ����{�[^F�_������g�s3�؝TsoD�&3��pgŰOn�z���q��;o
c�_�<�r��	�uM���o�]뽓���4��I��xj1��$�l{(��S���Qn�ez![��s��gT]��κ7�i��fKץ�/X���6:�'J��ӌ�t��nx�n�r�B��N�����J>�swWf��8T�'�P&p:�2�b�Hޞ�,���(�:,�oˣ���*n�mɑ)�.�V]!���Ғ����<�F9���.�9�5�c��W�6.�/y�Pȹt1T5�])�[G�VY���:��-�����na=2r��Y�@�仁Γ��z�Z�1g)�����deN�yG��_�V=hv]�7�MdL�b\Pj:�*�;x��:��6��_
gk*�}8�If;�����S��)���\��van�W�Sv��n��*=T�L�J��x��n�^����Zpu�w��:S�S�د, �Y�.��ќ����s\�Z��7�$��;�ry9�oH���#�����m�s�p��fxmat�	}��g,��&W����A���&uO1���M5��G��`�i�R.��WQ�)s� �r	K��b)�d .�]e�GI�0�p�Z�7a�Q��GTo:�>���[7ڰi�VCK̪�II�{�%>�!0����OC�\ ��<&��`����H�]/K���=��/���� �y��Uf�~��4��Y!�k�Q�H���q�/����d,y��p��5R�LR�ys��f����T���;�z/���<�4�R��O���sb��ׄm�O��*;qм;Ua����m|�=ʲ򁫵��m���ʈ��Vk�qj�~�'a����Ә�.��q�
�=mU�I$ܫ���n��Z3<^�oH��
v-����~�!�c@�@�=4n�r��D��Q�kW�JM�ܻ�h�&�}g�Q~��-����{*x{ޙ�~���K�r_-�`||��w����`��8�R���縱��Y�q�����O��C�I�d
�ɧ9ݔ�ߏV���;j7[��&�,d�8V���2�p�87��Y"������SV��l7a���tP�����j��I�3E�s�*]\�*h�%v���/޸(Ү]��]5;'A����ST&�2;N�Ӹ�&\��,��������|��{Y,�4����Z�1�������dٿԗ�l%���|Ҡq��@luL%��v�������sM�".%�]��w�}���틭-;G��ў@��^�]#�řu��0�׺f�_T��m�;�K1�,��O6�sv'��e��YQ�~� f��\)L����\��b#&�F2����H�\�{���h�|����R����Xm�'�N]�K<6���,�78�0�����\�m��}�ҹi�BU��z(��c��@���\:�l\:�P *0ɍ͕km��ܧZV�� p���#y�^9ֽ�u�*�%D�����:�~�b~�-M���$	�)�����Z�L�H�|`1�4@ˡ�]I��lhFRN��׵���0oiC��\)gW��>3o�*k>h���/���w#��/��.Y�(xj��GM�m݂��\[��e�A�Ջ3O:~l��'|ʋ����B�R�52Gm	�0{%��F�K6B����w1��Cw�Ź����(�~^�:�=6>\ި
5��5��%鯎R�=��=y>��`�=�J͖����5].G�:_]�~�t�b�Z���u��]yL�I4p�S�h���4ыxg`<��Ȇ�s�u ~4Ի��2ur\���\/���N܁�u_g���X�y���vr�hv�k+�?N=�nӀ�f�7�=[��pΜ�j�h��{��m�Os�Yc�n�R	(�s� t�up�l��Fq,0���fAk�-�B������=�j�߯}e��+Yf��/�
ǟVU�-=3�YoH/W�(F�uH�P�9<�u��ٙ�O�����[���ȱ���]B�d٨����VTw��)����ݳ<'p��(�1Q�G��Km�$�?_=s�y���@|��Dp-��cL\�
f�;�d !��m�����N�&�Ď���g�9�yq�X���?{�'��fF��;2�]w�ʵ�qt+�q8�7	%�L����v���j�8���ܗwA���}�$Vrڒ�On���+yg��U=2\U�sA=X�]�j��nr���2�l��o�� O��I���z���r��W0	�.�]�/�T4TC;a���|�)�?��5�f��.�����g@��Ζ��^n�<5EI���[]R�� k�3^��%.�I�h7T:�L󘦘�)���S�bU���9�:l�	����-�x�k�[<C��N6R���c:��Ђ�ɜ��
y`��53LA]����hJ��~b������OF����6�n���u�RS�br>��Q����{����h�K|T��سޣ�]}�
U7V�ف^����-�^�WF��k�rc{���~äQ��dɪШ�N(�2뫋���]mun�����m���Λ���S��u��;w^쿡H|r����.;̶���NީϺ'\�G'�{�Y4ѕ�U\쭇\�=&p
�<�p)�������fLAt2�Me�L�?N������~�h�z��~� ?���5��*����Q�@�_	�k�u���]�b��{���ҹ�\�=Z���*B������ń�]�:�u4(�jp{|Hlҹ��*G�}�f�V;͎�~ir_'!�>��%�$k��wI��0������J����>�kT�@���*���h3ޖ}4M갩O3h����e2��T�y�B�yz��z�<��Tf���J~w��X_����z��t��c��,���X�v��Y=U���y���oDrlUӻ�0�ɸ�i7|�=�L}�ٚ5�	����Z��
]���r� ����[%��b�Lڬ��WӔm�_HΗ%2��n�a�^J��9�і�"3�4���4���F�-����d�A�X���P���\-L�h{*x�o<݌�	��*FZ�w�ʞߌ�j���`�ĥ}3u]w]R�m�v��K�w��O "�q^3�y��L��auƍ'����:�\VOuU$�ܷu��R��O��}j�-GF�|���Uc(�ì�r����������kB�!kV����[y�;{M�� %*a;��W�0'����^�S�'k��_f�}#�iX�Z]l�(���zC��A�GQ��,R4)�eh�#ꊺ��؍�ܠ�[C�1#p%x��Zɒ��7b�V�L�K�edjճ����	:u����MV�ѽ{�k�ڕͻ���P̺�u���
��ޭ�H����\�ISn�<��(���JU��O��;�5�y�>�4�ٛ$���=��e�I\\�#:gR�5;	#�z���lR�����\��k7V5>�LǍ�<�}8k�v+���[�7�:Q�+#�/F)��W֝k3�\Y8:�Pv�۫+�Vc˷17XG��Ir�[��%V�
4��R��;�E��,_��o��VD���H͎\�K�^��゗s�9t;}�ι��,���_Q�`>'W`�TS5�\���Z.����k��s:2��{�6(g>ǹc*qA�r�J��sK�F����uk��%-r�8�Q�<�K[Q��q��v�Ԇ����JW
ݾ�jW��Ӵ�]�7�����5��r/��;���4s��ۀU�v*�)�lu���f_5���"��,�����ut���W�-0�Xc�
�3��|/o�Z�^kQRq5�t]mX��&�n�X�8z�]J!*غ�ܓ�]�鋎�+�uԐ��E>�cU*�a�L^����;�E����r��RVT��yS�ʁW_�d�q�ڻi�h�Fƃ�o��	w!�X��ͼj�q��1�)<�7t��Ti��FD��M� Uǫ���:��b��f#+kp����v�����[�NK�1�57��ъ�-�}�t���u�*^K�.�Q%����ɛ͚��k�_�)>�|F�w��gV[��9���9D������i����Z�U�FwJSY����+f.F?� f�u��KD�y(�A[yD�s{�����̙[��܌�X��6�>��+��H�}����ڣW���l��Z\1ʓA�C��%j���v��9�z��\S��Nˎ���SGV����O�s$$s�j'����i��3��PӺŖ9օ;�ީ�1�Mۣ)��VLZIB{�]=֫DF�@Ø5���V��x��Yڳ��t�X���e���ac�j2^fw[!��Wauˡ��#��iA�'a��uPYȝ�t��݅�l�Tp7�vE���.��'���JY	�¥)%�x�ɪ�v���	䥘�Ǎ��kֻw��ٴ���YƜzI�"&J�\�h���*8;a���P7���ᝣ�GK����%�x��ؖ�7����vw�o=z���ܨl�w�rQ�ɦ�gB�n]�8Ks��r<�惵�w8e�W��yYy��� �W���Æ��H��wy>c����O,\4�6�Qc/�oniy�|��ޛƼ\��E�Qb�ƼY�\������5$Q�Ɉ�<�k��L�\�ݹs�6-6+��F��k����ss�n��/6CFM�u�lRE���g+x�x�K�Eq�]
H+��@(��6���+�F�ɝ���R󸍯:�#x� ���v�v^urx�CE��wm��pwX�s].��h�wv�6���&�ѻ��&CH��Llk;����yܢ�������d.I� 2һ��rᒌnp�u�yШ��
>AyZݵ��E6�ʈ(f�����ĸ�v�����4&�Ww!o`BG�ٸǛMN�X����ڗ�Jpݴ{���jNL�}\��G�{P�,2ӑ\Qg�
3yk-[�7s��-��(�ظ���yf��ƞ�1P�sQ�wR�����1a��@*)�%3����E�����vPR4��z^\�N�	�~p�������)�V�e�@a�й�$W�c��ON�_���@�?MnwfdJ�Y���q��^�Tݶ�s�����z�r��>���p9�t�A�v58��w�Yc2]i��bGz/��_����=�#i�$���ʈ�^d�A�XS� eK�\paw�s��b��uٯ��!��Nv�M4$l�gW<_q�N�w�vt��f�BWDGB 1���Y?$�"���6�7/g~g���y�tC-yc�%�3ԓ�z��q���� ��^el0��>���߇RTԜ�}� �F�酯�,:瓚%�k��?Y�s>d���Q�M�^���8z��꺀���+�nL��[bE�(�y�l�����3#��j���Fu�C�c&�KmD���<*Ij�w��^����ylif�/n���r���Y�m�O���*;����:~�ׂ�����H�#�+��K9�ٯ8�N9*̨{TvR�}g�1t;f��/� l�g;�r�P��˒T6�ٍ��V�j��H^�#*�UܭWO��3=
z.$摗[2���x�x��ԣ(�ػm[�K�i"��,���8s-��.�Ȝ�AN������Vp���G��:GLS7t�W��
�F8�c�;P*c��ݘU=9��6�%������:[J��$�]���]]!m�e�-��M�4�_~Lo~���o���>7	Lǩ�S�\�ۗ��]���p�f��-�u�������T�<���<#o;o2뜗��geb��R6��ݚ��)�=>sDysM��ׇ'r���5�T�~Sy�Qщ��vSXd,x��9�WB��[V��qn}jX�G\�7Q,z	��R��LҠq��@luL4��vymۜ0�nc�)Q��׫��O��[3�V�jl�%��ܚxB���]
��/R�'42$q����ȶ�A�8o5�w��V�S��6wК���үL7�R��$�2�^^�^��^#-��g��D�m���ݟ������}V3���׳��]Hv���s	��˻�g��4�<��\�;�**0�i�|����f�zb<��e4ס*�{=�m�t�������ͯP��B�)*(��l��n~3wíO _���L����R�]k�즚����:��:��>�t����]1q�0p��a�2ES�W]�k6��-L�����z�O�X%zl\��g_pƆn����
<��=���UM���_{��WGw���t�vk%^��"�W��Ổ����ψ�6܎�У�κ�.��q�anVS�ܷ�"7%q�пӊ�H,;@i��Uy�t����:ד�:�.������>$tZ�ff�>R��{;��%ޯ%��Ҫ��Q	��a�4� ��s�$T��|���ͧv]����.<Mg*ͩ�7��#�S��3�'����W�4t�;r�R�z^��ȓ��9�44��a'N����7�g5gS��F�E1Jy߯�8��zl|���I뮗��xw���}�m���@wxm���&��a��~f���5���ᬒ���,�������d�#)���Ǧ� �i�0��v��v�f�Fe�b+�_�7>�+�_"�>��U]z�����2ސ:^��P�����a^w�h�X�Nn^T�=D0��� i�d`�f�����1�>\�0��왊�Η��o��:��"����f������q뾋����A�{I:�zSV��	ɋ�G��m��n�k����ۻ�$�d��u��2�f���1Qn�q�n����Ц��ǯJ�8����r�����ݱ3�k:�쮬q�`�9(��T��~�rڒ�槷ri�[���'�혺����K��]D�'E�R�J��ZW�+H�>��=�� �8�!IR�:�4s��[J��M�J�kw{o=��j�a��;�k���O�E�#�K�}��V�E/ok*(�f���w�}�({�x-�؇����WT'N�Q��Y�k�.+&�����Uk˿Ќ��5��=�8��<8�OQ6��(��s �Tw.6E�몈/o�y`R��rb�2��.�����.܆{/:����)�*H[���0�zەq��~�S�O]�苆�'%�!�u�T�J�c���q)���;�9ֽ�g@O��.ǲ��E� ��ë����zU����L��*^4y�CSLA]�����%D`����h��j���W�6yc�������hʞ�Nɺ�9�3�T��'|ϰx��t6��������{R��F���:3��[<1tf;�gSF?L���x��`��@��qyf��&ѻh�LQ��}��8CgIͷWѼ��x�������͵�N�n9$�(�;���vQw麨-�87��{���if�Z���У��i�Qͭ��������`��]���$(����;¢��f���y��i�;�%��<�w��ZJ�^�B�y~�3��Ǒm`U藛����hsu�/�H�R����Kh;S�lT.�¯�z��^u���(�����G��m�x]�p
* ���U36�KulwS7����2�F=�; ��{5w(��p�e���EQ�X��gDW��{�N>��-��=�1�olu�����ؓ�FӔU`����j� mr�{w��Ŏۺ�"��/5��@�Un�����;l�$]ٹ��/�֡0}��\e��yù�p������;zTc�VAX�[ᷰE2 �82�֪��s1��� �[{�'�v���ӯL˯*m����* �=Bn�uB�xh��`X���)ºݓ����'�u�\B��T���ǲ~�������@$�ey*��Z�9��vo��%f�d�DZ`	������
#�-��7�ǲ���;.iX��5^ou��M2Ms9⾃8�g�t�"�qz��[HT~��t��nx�n�ak_	�X.7.dN��rd�ͩ�6vj0��b,�[4�q��iP
��؞ul��,&�S���Ws�Px��ڻ*.�VWB|�U��m�M���q�=чe�4���T��"��򸐤�v�[��e��l���ۭ�75�X�Z�(e�HO�ܪ{�[0�3�x��Oa�A�$"���)bSM��.��)Bʞ�9�j�H���X\r}M�#i��H�z�s�lam�v���i�6/�=��5�8g1��6�k���i�H����2�Ѯ��/Y�����я��V4ކ�o����jo�vo4�����7t��lijv)f���֑[�0t<Q���)ز�������.3J���ܺw�#S]p�D6�lLө�h�x�B�+�\�̎�9R�>��C���2�\�+���yxplpi>�oni�6l�����.- �_�)a>����1�V���q�.}��eڰi�Vp�)9�c�_5n�~:�:�N-%&�b��5���mhT��ؿ̯�sD��(�K�����Si��Iw5D�yޣ�-�&�E�`(�^�Er�h�$v�T�=8���Qs�Tf4Go!�k*��n�N�m͛���2��8��_���qO-�-�^�	�랗6*��v�G+�J�Ǟ�S��{��/q`��X��ά����]U!g@��@>j��~�l��맇5�P�i�f;#N�Y;��_��̅�\#�^{�LXQ~�WFjOO����w(r�lȾ�_��{�c@��So����Z��]�tY�P���#���<��b�fV��7�{zg�m�mຩ|b��e�2���^kmB���<�* ��:�
.#<��ykt��*n�Sy��e=;�ߝy[��I�C?0o�=I��껼x��E�ƋY��������cJ�ܥa���'�"^��L2��G�;0�=�])�vOR�9=t۷����^�[R^��ܚg�.X<k�M1^�T���H��F�.�8��u6�p�#���uº��Z�[h%����Oj�K�^���u��q�Po+f�_
ٵ!C9.s;�[J�zc:l����v����ė|,	�f�������-�)N��'P�����������ޞ+lo[��|�i��%�_j��l�փ��e`R�u�\&�t�9��#��Nn�s�˻�xn.��G2ɺ�O]�e�Ń�_�cF���ot�-����~ΐ;i�u!���7$+a�0���s�*kW�Kz�gn`�����T���Sú��Z�it���Ǡr��gH_�������B�P��.*�]^��껾�y�\ 3�}�2�aC�'��ֹ��i^���	��qo�����fzi����Y��t멬y�!:`5҈a�R�C��"X-syoB�I�5u��@k�>�f�m�gUQI8ǻw���ѕ.����5�H�{�u�K����ff�ᩌf'Z7#�V&ܼ[��7�upB��Ɵ��"Ӻ�s�c	]}M5�S	���ۂP���MG�@����[�8a�t�_i؞0�I�N��T�f)O;����G�s�T�M�$�2�VVΚ�w�ѳy������7+���&�Yc�����Y�If�_�x�FS{���r&s��jN�^�z�������[��5��~�_��YF�����c�4�����@sc��)e{釛��^��)�2�G�E����6�C���>��p�J���_u��`��x�'��66��཭6�"�����񬣹(AY+���P�I8{œ�j��p
K^զ�!��B�M��w.���Q�la��ụN��5��K�K�F��i?��������1`�v��S^�||�r�i�����n�� ����l�����9/w�zݩ�D!9�M��Es�=��Y)/���X=�pO�/�9��vi��������E����*9�q�=l-��jt̳��_�u��X}l���3�%��J�q���Z�4�Qi�v���I1���al�g���E����"������Fc�f����j&3�+}�wV]���m���� q��#���R��%{�xq�i�#���#����x������ܼ���!S�N����Ψr�D�`Sיl�
��hU�	�_����t��kE(�猽V�rb6�EpQp�^0C��}��2ʚb������ħ�Jz�8_��2P~�+n�>���+�k���?�v�m�D�?[���3�T�h�`���CT��j���y �0�Rz����ؽUU�Xܵ'_��c�{���)�z�;+���&p
�I��KĻ��t��k�0p�ܙ�<E�)#C�d��~�c.9��iۨ�4�B�3<oH�ݷ�r�UG"=C?T"�g��O�|�w���qzp*��JN���
D�Vᬮoj�b�;�F�nɵmh�&]b��a�`�tz����8���<�f�\�BЯ���ǡnFq�Y�a���P
�8�U�k7:���[R�t��M�ݼp�|�ݐ�]��b�t�on3�n��R��/sń�]�:4u��W���¦9ɂjj�Ws{Ť��{��"��oSF����v���F�^�t��m�< ο0S�]��2�9��^���4��\Z^�1_l�ݚ���Q/�P���k�=eFc����\k�y��b�L�D�����Ϸ�Mc��H]o!d(�^t�X܁���Nٱ_.�±�9����wk*�rR��vao�28���w�=�	��z�ԏw�Q�B��v0�m��c�K�b�]6M�ǀ���O�7���Ur�����-�� �_lO<��SN�.����p.��ḳ�;/cD�c�_W�U����˿��7V�붸Y�U����{�#��lR�ʑ��1�1�_:[BG���J*/�-�<k���id�Z`	�kڊ�e�d{�c�e�$�$s3A�Y��/�X�9��S�~d���%઎*�������a�6 ��%=��I�n��؞�/Z6;Vy7q�W͛��2�;E�8.e�2�#B���0�*yc�<�����, p��V8���Q�~���K����7r��:���T�r�u=�&��xh��gwVGV'r��-!����̎��*l��od�7g�Xe��=�R漯8�b3�p�z�IXO-��j�m�����ϴx{�����b�^K[�f�i쩨��1��T�]��-��6#9�J�y9u/��.ss�ݕ�z�z<��5p�^`?B�`�3T-�	ߗ �)�ʼ�ا:Fw�3�����<2�:B}��y�b:�])�Zp����u�3�ͥƺ�qk]\�	��/ޘ�[+��!�鱾c�������3vI��=-͕27�"j�1ZvT� �v;*�(绐'�|��v8�Ͷ��i�#d[3��/�˥�_��ﺪ��i�����Tux�;Ғ��%� a��E��0(\��c���Qռ�����_��X1H�樗��ţ�ﷆ��5�5���y1�x�?�)���aѢ%�?��Nh�U�p�hܽ8���6�7�i(˺�:Ջ3�w/�ȋN�۞p	��v�=/F$���b���B��^�ey�;�]f�Kds�͙�R�LR�qK��[�ɢ���Ƙz��`�Z��{�yPz8tM>9FR5fl�epٝV�UT�Y�:b����iǭ��a,z���K�ݬ�q�)Tӳ��6kz�g@�>����/=���~�TT^4����ʮɠ�bۺ$mʁ[�mq<=&c�]��k���J�I�ԃ��wn�m��J�<t�5`Qvp�f����_t���۔��� 9���Q�_�.՚Z]Ьr��cv��k�kݢ�����q�;"�<��l�l����W`�7�1L,���jTC@+����ER�([N[@ڱ�n"�֛���f:���Im�;���c�&H6�3�<2wV��(#3J�;kT+Y{f�sF�л�m�{�ǐ��lY�G۸3\�n@�&u�/�bՓ�L;�ڇ=���"e-Ypօ9%O���1-�L����V�������%ͩ��9���c��x�Iw|t��i��q�s�>�����A�o�:�h �7��+����x��~�p�1��_8�F�N�mw!(�'�gH��]n1���8��k�:�W:k��{�:]Ѷ�r��ӍF��P�0��;�Iưs
];�T�ֲ��EE��Y���=�f�T�
���XMd�8U1��t{��R7��4�Yj�\�����J�:��X*%Ι ;b�R���>0G��].SMi+'
鶛v���T���Φc�,TV�X�o;q��ͭ�I�X��4���[ytf�w!�Ծ���9�Q�\��s�l���.����_���F3����x�ױ]̥Q��d��n]!3��,��Jl�(`�Y�ȫ0rW>*�����B�u�5U�8�����FN^�W6+47�󫷁�C�?q�kp�w"�֥IW/����F�h[c���f9��w���c_.Jf�Rb��A�t��T��U��5���l�cE���qd���2A�lg�GoX�j���V;��b_245u�ep�����İ3��8m�S��al���yь�y�q���
�8���ө�2�Q��l���η��v�i͠6G�19\Z�Juν��P,�W���Ƿm�z�����t3Zκ\s+��X�̱��Q��a��k��	�r���t3%4w}6fF�(�́���	R!��U�F���ma��౬������م�cg��x��E�����Y����9פ�tmWs���N���b!�jd����V7���ˠ0������]t^9}Zj)@o�e�)�i�6�af��(oQ�b��Bҫx�JH�<z�Wr�h�%�W�t�����u���n4��>�]������6��3�3k����Z1�
8�u.�7��Y4�p���&�v�5��N�2n���3s/�v�H�V:v+/��;4jgWon�k��z�ZEC�*��*���:�8��6�pK	�{\hy�i�t���>�$�{�]G��S]�]�,ܜ�������qCM[���zr���7h���}���:ۗgf��y�c����#v��N��V}�'�gۛq�Cn���F!�)�#ȭS�E]����vß�lX��D��5+�,��$Bw7��7��������7��-��2�u���'yc�ǿo�2l��3����2�&�U*+��bJ�%1�����l���8ȫE��x����G�����?��ϟ�??�b2F(Y�3���;�K�M��#��]r���A-x��,r�r\�x��U�d��yݼr��\��u�K��.s^uэ�r�#F;�w�]7����EΛ�w\�"�Ӟ+�/;����4�䘻���s��9��<��(��x�[ɍ�-7q���"��\���wv��Kݍ�ܨ�7Q݃��9�v��
:x��Eywg���us:v���i��`��WwAwusN��s�:t��bܹ��.��\��n��ht\st��]�˦�s��l����r�Wwr�v�$�sw]����y��;���8+���]��t�wqq���^/&v�+��˚�뒎���M\��'���>�( h�@|G�M,�����g:��3tCe>۬:���@v�QWon5Ck�Ɉt�p��͗��m��E�}�P0�r��^��Hz���;���X��ù�C�����!߆�U�E���k��7�6t���
��Ռp�욹��6u�K�v��u��`U73�M.y�M�a��F
p)�,܈��_I9����x/
o���O�'�-mɳdpn)hب]!�՞�՘�r]n��=J�(m未��Q�al�z�;p��3=���%�(������u�Y���ʄ03�\�r����f����bGl~�l�W�.��7�$v����]H����1�k�3H��y>6�������<�` �wMl���Ζ[^]Hv���![���UQ|��z
7���JtIp(2a�:�B�����3œ]�y�(���׮�-����d]����-�z?h�R~�����^@��:`a��^�/���SMBTAO\�t��C���������r���O\צ�e*�g��r:��d����pMD���Ν
�w[7 ��mҫ�ȣyד�W.9��5ۨ����fErJx��@�0��@��L/�n�{�8��"�{�U�O��M޼�$X�)�������v� ez���8q���z�G��;@p��ً6f���mO�TE�E�'(��gC|Iݾǎ��Qήz��fTu�ѱ�Ŝ�W+ԭ���e�Z�'.i:�Nf
���+��.���F��NѮi�T�i�����q�羈���l1u�4�2�������kdy4rȊ�pfj�<�����7.'��GO��p�N�H�)O;��s��������K1뮗囻QDQr��݉7��
�w6��0�
hu�sW,��۽������G��_��ČҘ��T�]"�y�F��.|���^�� ��E��+�H��*�x���G{5�a�Gc@4R�[k����yZ*r�T�w�=sY�L��DV�����!���M1t���5��e_�G,�ۖ=L?<4��M$dn�Z��X���y����p�?}M�D��=���c���F	hz��W�������6g��[gEs][�M�F�Me����]��GK�]Z��tO99�5��M��R)=���<2�~�!Dm금�C����᭪���xvOg��;z�&e3�������wl�Y�jK�S�;T��r���s���w�8�Y�P�fp�8K��i�ԁ�A��|ǲ����[`svG3 ����Pz������A���L�5��[�1��q	�w�Sw�ݥϴ3�^�٨P�[W_�r���x��vu�B&q�}Y��:;܅�x�Gi�yB��|"6
b��j��d��:.�����4��y�r�WVs�z��mMgWQ!��n.}E\�	�X�ˡ�w�ˮ<�	U�c�02$8Pͬ6���k��k��6Hw5w�3���!Kb���I斀�~�^���O�=�u]i�r���*
��OE�v��ŏs�g-�q��^�i��D�?[����T�Ɓ �,����<�7׽��E���ؤ�uVWX�����Τ_7�c�vK=�wU'd�Q�ɜ������m��"[_�����;|�uٹ���9ա���4E���c.>�	�n�lӪQ+\��ZD��/u��D;2۾���/j3=ܴ��~L�Nm�B��T��?F������0����b���j��F�sjQ5���>�PH�1�Ѥ{��1̭�
:��].�������3��f؀���~E�����~�~�~���sw�T��:]L�aZ�fѫ=g1�vGv�#�;=������h��)�_�Ґ4�<�o@���N����t���f}��V/aY���ن�d��ʾ×W�x�U�Y�=/]И�n���|c���;"��b�f�.,�-v�����*�]��J�7�^m�]YUam2��ٖ�z�O9}�ӯL���&�D<�}�V������}���]7:d�@����������u
��
�i�!���W>�ɽJ��3Ju��G؍���==W���D �_����w�G�l�<�R;�q���9^`
�%���L���>�f�%c��aV1�{�-=��j]����ӗ���E�u�>:��Q�5���+�;;���Y��/�eV�*;z��Gk�{;f�2�ʑ��5B�~�޸��\��pf7���Ix�Ⱦ'+�Z ��ƚ�t�qjg���$�APlf"bM.��[�k*�Op�E����/���Bi:�q��1E�@,ֵ��ܛ���u�J��������3J�m�n[hVr��"��s>�@ȈЫ���@Nq��%}fڠ��P��ͼ-��W.V�Ǒq�[;�MC���^�Z�l�>�ȃ̪��>��|��~_��o?Dnh���Y��9�q#�W���׳���|g�7�ҝ5�	:!]vFD��W�o����]�����LB����!�鱧����:B}��#���������ϰ#�_=��BZ:��0��xja���=K�ǝ��i�4$l�us��t5�nΘĞ�YE�R�~���'�N�)�� �d�3u@�;Ŭ�o&�ԓ�z���]|�f*��ۉI�O�u�zz�y�%�*�%'�F�=�PH1�	Q
v���[xr���2\w��Z�o:���y	��
�w���J�`;7X��1`>���i����:�F���ͫ�ʶ��Xz=FWT�+WYݏ �J5��2�}���X�Τ0����&T��ΥR��;��a?i�g�l��4�.�\��CxUuFn�b���3a���}:a��'/joe�ܧr�����1�M�yE�Kшp�lHt��#Q�T�n�
�T�%S}S7����j.�#U.��.��9�u���cOt��z�鋷aNא�+�h�����a�v��3Xsb����q����bz�
���S_7,�u
�c�Pk�;�Mtd��Ka�*����2�Sv�/�^z#�
/���/�4U�P����Ce���F�ν���=5<��Z�N���F�C���'ƾ��o�����EGϲ�Y���7Z�q�N-��U��gb������0��gZ��сE�k��q6�5om27�X����8�|o����R�����]�_U�V�֧����h�����i�1��)�@��n>m����SQrnv���l����v�6v��Fg����n�(��3��<k�']̷V;ѦN��ɸál�zr>��o���+��.����RGjx�c!���P�s�Mی}x�+����5/8�Y�X*��P���Hp�F��9���{:Ym.�;^�ܐ�LTCa�,�~�F�Z�c�n���c���
ѝ7�����lz����Y�,�}6��}Ku���6�*��EC�{�@�'C��t��N�thع��p[�7	]��v�bj܉���a��؅�n�nd���ٝ�=K���w=�o�����[s��K��p<��p�d�s���m���؞��9�/?z:�<�U�[������ y�J@�%���y��SM4%DM����s`f�tJ����}�Ψ��<�ؖj:��d���9 ���zalv�x�ʎƥ�/�o4gW'aղ��9�&�m�M�uLȯ�%<kH�����$j.�T�x�׬Mn.*���n���u�.7��i�������"ӽwKc	e���Jbz^�b#ZKj�����Ԛ��$s7��֮L��oË4᥉ީR�w��:�=6,��Y�ޡ�*٬�Fj�Z/�2Oi���D�V*$�|��:�c��ܩ��M��mANE�)��e�v̈�ќ�e0�7h<��_��M]��z����Q��Gf���D�7:Ľ��^��N��{ �]��J���Ro���ڭt-X��?�'�{ a�~	zG�ݟ���cG�6T�E~�͹��esI���8[嗢�y������k{����/.��!�Zu���9��GX3/��<n���j�������L@�5)�{Q+cr��=͡w�m�e���؎im�-@��>�C��^��-犾:��;Yoy\R���a�����W�c��_C\zM/4Ӽ'd;�7)b�U�K
Ⱥ�u��`�����Ec���k�vG]��B��uj{]�O�v-��R�z�g�^���'7y��,�K��sg[*�%�6OeI1���ajg�A���K�� �-�/�m0w����B������V��x�3�6�KL��L�g�
3T���m�����z�LӅx3��k���4^]H�EN�t����qGT#<^�]0)���W�~�&���k�l�����.�VW4,�U��ڛ���t}PC��h�q�U�&�g���q)����61u��Cv���m�ylu���>�Mڞ/���ňOL�8u/00C�䡢���Eۮ kR�ꭙU*��NG6Z�Pz�`��ԋ�o@���-��U��l�nc��3�T�h۔ ���>@�b�i�[�\���X�jpH�H�����eӺ�^��h��-8�&9��-s�G�v��績�3�  ��o�2�9��
b�R��;������0ˑ��C��w�\���4\DE�w�~���bkQ���7~�1̭�
:���h���7j�����ё�:�[M[�˨�;��VM|9�d�u}�+S6!�ɼj�{w��Lg��峷��L#���Խ�>#sv��m���]
o��.�r�6��0`'�%B�6��Kl�c.�g��g�H��6�e5�hR��o>���.�KV��@��a��O��A��f�a����94ObaR��ѫ=ef0����6'&*0�lΚ�w\e��!s��.�z�� �1d>��~|��_�J���^]��]8'���J���L�-B2��_-yɩc�Ω��p�4ܸ+�t��=F����FC-�a��e�qxΪ��o6�ܫ��ҳ:m�w�A��~��V�3�mkzCSN測���,5�t�}�i�xM�չ�����6_xFc�E��Q��%s����Zʞ=�:6/;g���DK��[Z�j��)���|�xcnC,i��z���sM���g�pQy��)��E�f0p~�>?4O,��/�g������c�9�B���[���Za����8�@S�wv;����LS�V��fM��}%��6��i]M�ݔ��ЪZ<z%�n�Z=>i~�R���#Y�ce-(]�iý+lf'Μz�k�������/k���q��*'��X��mF9�x�T:xZ����q~�z-*��iyo�"!�s����\,g7G��_2�9�Necna:��>�^ہ1��Z�Τ��D�T�"�gEr̝8\��0�Y���h�I�J�g�N�y]����e���s��%v�+O����>�	� �����[= �*�e��Z���]z�r�K&^��NV��#�"NMR���p�մL2�g^+��`�_D;�|i��z�Z�*��g�9>�@O�ݒDc�7uu7  �ފ3�B��U[®�:%�0���d	�� ���5򙎳Q��B���d[��/�����e�,��\�WCg?�g�/�\����� �h�*���H�\�lC-yc�����'Y)Z�\^��b&6�Uu�I��rp=7.�M�5�5��µI�$��hU�����cO�ҪW�M
�cY�vG6�ήN9��g�����'�\s^e
�F�fH���B��s�]�4�#)�@�0�f@=�b�<�\��L�T̑��j)u??;��[Yt�pTt�1�n-�i�$�ɘ&�w	��ިv�6���c�{!��������^Y�:b���޿'��}�`C���|��33�#�F�|"�l���eB�vi��ы������j������vM;
7N�~�w�[t�lI�Z1�u��Q��:���5�GR�vi�l�Y�U���z5$��*�O�b�O+�fa������ض�.��{�1����0nluB�Xj�M�>�aՎ�&����Du�(H>U����P}ۧOS�e�G7(��αA�9�_K��V\�+�@�Z���?+�[O���k,�7T WL���fv��V�+l���9��X���{���6��`Cp=�mU�VvZp*�mX�b�;�t�n��×�v*9�a�B��S�t�n�b���z��
���B,à�S/��W%Q���⦮�V�D��Qa��<m���v�S���'��vۺ��Sg-�/mOn��<!oZ���F,�&�y�5vk:5�w�v$�J��[
X
սHOu�s��#��D�v����SUj�ݙ>��%S�N31�Q�LR�zjHS-�+����ϗ�<8�U!��*21z��/%V�n_O�StШڙ���w!�Xa�@�B�=��h�&���z(�O�} I��̾���z��l�r�u�l\:�P *&@ba��BO^���լ����0�OI�ͫ�r�sl��"�S�R.�Ү=��ĳ�u� k%(>��$��K_�;:�"�p��=��ս(+�ԓ�����_F�|��M�I��)�[�$M��y&:7h��9��"GJ�����p����?q�羈��]�M�)�o����'����<�h1K�7fv����@��{*^���M{!��˂	Q�]է����������km���ֵ���kZ���m���km�5mk[o�յ�m���kZ��[Z���궵����mk[o���ֶ���kZ�|�Zֶ�Vֵ�~Umk[o�U��m��U�j�V�m�_��Zֶ���kZ��[Z���[Z���Vֵ���b��L��9����%� � ���{ϻ ����3o ��E6�CQ4h  -��5��� ��� Ҁ�B���5
��m�j��(�s�OJ�(+lše��%V���֠f��3i��,�s�A�Mb٭2֖�f�Z�ٛ&�2�eJ��\KX(m6�m�1C-�j���j�J�Y���Kڨf��6�km�ZkU�Z�6�4���k  G�togq�E���a�tö5�Y�ʜ�v���5�R©��
:k�ժi��v��,f�  x������4��� wW( P 9΀ ��r� 
]�^=( �y�Mj�����L٭�����j�   sW�{�݄lM��낋w;�6�79à+n�Ҷ�S �XN�s�
�f���l�*"�%[x  ;�{QѦηj�UmW6���n[����u����w\ꮆN���:�V3"���i�U.��j�*鶡�fՍ�VU��� w��N����.w;UZ�;KU)u��t�X��Vڮ�wu�۰M1m�.�s��u�+vۺE�U��m���j�%��x x�v�m����n�l��iU�n��;���[T�'w�v[N�]j��ΜSfU��u�H:�f5���T���Em6��<�z����meV�u�jj���7Zr���d�5-[c���������ƻ.�+j�6�Fr:2�]�-�ز�M*�^ �o'f��[��������-�[V�;��Bӣ�T�t�+f�LjU*�m�Ά�7m�h�[�v���"���3�Wa@�MP�w:ܲ@��;����l�� �V�,�֖�cY�Mjx f�F�ێ�hs��h�w���4֝��+���f):�Zс�t]�4�
 
   �T�T��   �  E=��*I)�O� h     "�ɑ�R�4&�M4`#�CO�J�(�0�d�Fah��M&�bh�4�b=CM43D� �J!�R�`C L ��& ����1����~���Q��kk��e����^%׼o��4耄F��l"�bH"8�*KH0B$I$�"#ҟ%Z��IF2Ea�������?��~�l)"�QI#$AQeDj�D"6TE��*&%�R"2�q�e�m��0)��ۗ���@�Diғ<�-/��_�t-(�Ί�d��:�';Kwj�p�Z)*���զ��~�o��R���Q+�FP����@ܑ�O���tM8�HsFWb�����^|5��VQTu2�I�B�{�#@Y���{�B�?V�1�ݡl^�Qb�)����F�V�ε���f5�Y�tHEV̠�9O^��K]aw����{�eaE��vC���P�3Zt�52����$]�O(dL�]�x\͋r���Vp�����:渴�5[��9Ed��,Y&�ݷ0��]���	j9YQ�4ȐDr�����K�o,[����![H�n�.�
A,j���lR��j�[`�ť��V���≷ݤ\J��D�vTn�m0EG]�L����]F�{	�ed�V��*�l���%�s�.������tڵmS���Ҳ�! B�oF)٪��l�)f�ҺE�;LS@e��X#c�n:�eeZs;���H]�N�kR���,�X2��f�U���Q�Gfnh��6v&��D\Y�l��E�ٙ2�AcE����L'r�=�,1�V��.��Z�;�>i:���E�<@��o#�]�, �1(������e�q��*n��
f���I�"3-f��\�]6�h�Z1PJ���V����ŇLB�فͽ�b�n�]��ݿ���D�%�d�+*P+��6��b��,�j��D�.���;��+5s[���2e������#o��\�[,���!wq��a���Z�l�q*�V��X)Hn�׭��ƻ��5vM�V*V�O0-}n�H�ͳO�^���j�M�J� �KM��Ԧ��V^�h��H����Yx��i� P�:��C��KF�-���]��>�Ɗy�$R���JњuS����b;7FѠO�;Cs�&��U���%�Ԭ�m�L�r��ՃqX����V���^�Df��.�V����4n4�+$���l+�[Y�+��J&��r��fŲD����U��b	�C����,m֌̙K2_շimKlkt@ȅ;,�ۻ��]J�I���.�SSz�2�*��!C��-�Y�`aR�2��:�T��fiA��U�si|��emX�2����`�A���]�̜}Ie�g�jX��ad���ǘr�f�.���K�U��y�S��-�9@�u-Y�{���Jm�w��j�����㳿:R���ckZ�M'u�F�-�r\(�uҼ�P#rm�ww��p����t�e�+X�Y�T:lE��x�^�5�ݲq'/mZŪ��d��������t	̥�qX�T@���f-J�$i���6o&�ȥ�xJ���F�f��!6c5�c"Nj��b��	�nB�W�Tn� Um��x�[��8�ܧ����
m0��z�"n�ȯ�u�8L�P`�T��:F�4�N3+a�f\�U(�Y	�����Ʃر�e�"�m�j�ԹV�g72dY����:.�iv]��{�Bݓ"�u�9�>5���E6��r��L�L7X�aԨ`�%�ټ���ˇ�gQ���H�y���S�*V��<R�p���nR�� mJK;�^CSqV���sC�e���VV\Q�/��x������e-c@c�Oe0���yF�*Lm-E>t;�~2�*2���y�� .�AR��w�[�E��eb8�<�q2�f֛"�E���2�J3"сC�J��n0	Ȋ�J�[��0b���eY��R�I�� �2ۡZ�1D=�V������2یj�Wb-��n�'�Ռ�����[G-�$w2�i*ϋE`�ybOU'�n���%�M�<��ESA9/&V�P9OIW`S�`1�XP�̒��=w+ ��᱋Vƀô_ט���r����q��)[��\!D�.�r$&0U��'A�C4����7gM��8L�u��U�ٯ4A�}u0*+xP?'m���J���b7�y�Q�V[u�l�v�Б��f�`�Rfk�uh�oQTXT���Dn�i�%��h����S'�=�*7�l�4�+Ga��h ���c��G�[{J��������cXZك)b�x- ��6c ��0 ,n���\J}��d�\ї��P�)n;*��(kzm��+lL�� ֋��ww\Z BD��;�b2�nbRk�2�83(�Z��tV���m?��k˵��+d@nV(�`J;x�ɜn�襻M�`�t��NX2��76�pŷ@]�h�78̛�]�!�l ���B�XP�т�h`�"k�P�)5�VhU���	`F�*_�=�[�r�_#�9�.���DMY����]�A:(��HQ&d���8$���V���R���p�Or ݹ��� &�Tʹ	/Dt����8���$�|��oeY{x�u���a�A�E� ����� �1V\�wr�4��̵ZA횳��S���&b�/K#�*��̂`��3��X�7.�k&S:K0�3e���"ْQ�[xl�p�����#ON�6�k3#`ЩYolVРP�e���r��a�[�0+yx)jڒ�,kU s�|/���r���b�+�,��R�7kEa	b��M���f�՚S"4Dg�X1[�����.��f�f�@ZC�QT��n�_kx�Ь�T_.}V���56V]76�Z�jb��˭z����K՚�Tldk.̢,�$To/q�mVO�!�B�j\�kw�uś�k;}ׯ�u�����ĴV�<�*ΕXecxi���ڱw���i�� �� ��"v���1����w^:���*^7����J�Gv5"����h���iV1{�N[4P�6|���t�V�G@�uj��M���wQԅ�p���f������kw~�f�)�6ެݻ)�
(�@�4��))j�lu�cN����e���|2�� ���[B��'[��Ƃ"1X̟ܫ�)!7NR
P��l�2X� D�̧���t1�.d���[����4�G(�Z.���V��=M�PyW2f�9��kgV�.(�j�07�{�����7n�՜b�I�"���#�1��Հ[��뙷����S	�Ev���y�vfBy�7a/���̍�.:n�6���zlp�gtm�e�`먖*��pJw���W��,��6�٣2ZݚF9)k:	),�˩��Թ�(���Y�Y�(�I�Zɛ��4�=t�*RBa����1����Q]ut��
En��`m������iR6��	�[��QG2v�Kh��M��Ĝ{*�U�v�!��`6���P	cs^!2�[�%�r�������9�-��Y��r��7s/@�Ҋ���F+��ͳjM��%��A���~Wl�Ц;[�vNo>�)|Ջ�2c�ۋ(4�� X���F�Y.��{2�dr�J�N:���]j-��F�kG2�[u2Җ&���A�� ����R�aF���(͛ztS�{MU^q���RU�X��^2�-�$�wY���U޻8&�-f\�c�5]aϵ��.��vsA	Ía����5�)�X��Y3l�L�f����ު�c~��hm��A \�F�ܦ�Y�5Xz�B���H*��`u��������h�4Pn�°�N����+V�R���zG��=R�}k4��P�[c��r̺X�V�U�7A�m�e]=MJDM���[��ڷ.�¥��̼ͅi���g6�*�L�m,B������)C��4Xx��!n7Ko  �y�\V��#��h�CB�]����*�-;$�� �ܴ��B�P��������Q���i241�ӥ|�����ѢC�Eyj�F�-��q�ݥ��n�:��vcԝ�4�Z�Lj��e�����X��@ٮct.�ȀtV�����*�O�
�ɛt(��Ŷ�ƴ��b��$���ˣ�z�ݕ���n��v]Mz4�/o��Y�Ҡ�n�kB P;���j�ϭ�KsYܙL
xU�.j��.����4��+kS�f��ud���J�/5���fZ�ҵ(��t n��R�ط>�DS�uۉ���������6�|z/V {Eei%n�֝��+W׺�ih�ޚ�2ugl���{�n��)XY��y&����v���,B�.�Z��7)RZ�L��75
6�Ƴr7[��B�Y{�te�"�<2A���L[���vL��{��U�7Af�A�K��ap�y����GKs.�+�8r7(�v�,���Vfұv�Ь��c6�@�����;)�g1�N�Ih�/�8���idvf�uu�h�J�VԎ1��w��wr;'6���r�g����E�p���F����E�0�[	���N�J�JMW��g��%�37h��`��B%f�J�B� f�D��WΛx�:��G	�.nZ~gK��iz�aF�Z9�ޭw75�R:6�a��iO�9xq5�s�.d�.�)F�����j�����X���cU�b�8|h�/�Ҭ�{XѬ�xͮ��չo#9��'�Ʋ����)�Sӽ�n�u�J��/� �j�����w��f�4�A��fXx7m�k�Y��uf�M^U��nn�nU��9�޺@�/D��B7�st�&ջ%!���c6�n�:B��J�Ӫ�&��ڍR�������UXǱi!ޚmn����Cmd_mrL���j��q��������٥���7k	ՠ���V�wA�6�n'�h�N�]���h �i�=�N-�D�0�]�i�����u6���VZ��Zec������3*����h*hLu�t6nR/���h�c8x��dk�=y���05mR�E�3A�*n�z��N`V���aQ������m��ܔKb���llH�l��Uָ��W��G��uZ�k)���}/,�)*^u��ݺ���  tχ�����=y�ċm��mԢ��BS���(.�v�W6,t��<�%;Y�+q��B����+�4`�Ǣ;7�q�	j�s�r�D�2�t�L�A�rO����[��B�껑k���#Eۣ�[��e�Go���F��bO��津>�n��Z+:�Ґ_K u#�g:�J։gn�|y��nJ��F����'I���e��q^��ʙ:oYl�Q����o�Iw��#6l�I�c��.r�U06f�LW�(���ܱI�ի���x9$���Gw]���G�2��ڳ�����o]�6��\z��zƝM��B�qw�B���A�m�+\���%�%mkd+GJs(���_�
|sf�@��,���9��=ELpV5���3��3J;�W:/��Sܹ�ի�f��y�[ǌN���{�k�mZ�ZI�ϲ��M��#u�t`}�`)�+$�%�s���m��n�J۽���TukP����*�63L�0�n.���9R�VȬ���FF�M6GS':�CMŶ��*�k�p��%�ɮ��"s������N���U���;��W[3�W4%g�.�k�ٹ�̈́���l���j��]|���;��Mx�j������N_"�Mq��'"��:HF��M*����Xԝd��/l�fw<��!A���iN�>�U����!Gky=��+ ���Di���)���ssv8cΓ�Xl�7�!�]F�FQ�I���W77^'@�
/j^���	Թ�x+L
%�n�y��ꃃ6��:]!�s�&Lٔ[�`f��ו}wA��j���n��s]��JLj�L����pښ7㷅�n�|��F��[F�����B��1�Ac�#�T����kl���C�(���$�-�\f8A�1g8��
��!5B�߄[x;Q޻u"[7NѷJ;�S�f�ȥ�)��R��r��*v*5+�R�;C�>����5>��r'���˛w)VB�>���r���:�l��SQ!��>`�F�l�a��M��4�V%Mz���E.O%��ۣ1T� g��;�/xqmo�ۮ�ӛ�Au�{�M��Wd/���yt�	]��s�e9��r.��w��4����X*�������s�.�Bd/��	�[P��j�Zt��ǐ����*:;:�B�kUi5*�\�n�9�$|�O�q��í� T�u�B�	�U�F���T�{V�dU����eY,�\�Cܼ��\i������i��|�Ie��0Ѐ�juf^lr����6*"��q4�vȮ�c;��Ȏm]�4��6f�}�8Ç��El���ޖ�ϥ���̙�Yڼ�QLi���ɣ�q2�m���.5��u^k��(4C̪G	w6+��%�S��7K8K�͆����n�eJ�AӁ�A��hf+�H��B�_�ʽ˺�*�o*-H���<M���3n�����h]��ɺEF������y���u���nT��ܱbp�bY���>a�WD���m*[L�m�e1��:�1[Y�����j҆(󦴬wF.mY��.W*méF��j���㲲������V@<>$�A��u[m9�o���8�&�u �s��)�
ӫa^*Ѷx�j\�D�S<'r;����j�[��e\�+p -P+��ktw��
Z�bn;2���Y
�5�OUZ�l[p2H?h�$<����Nٱ�/c�Z=�_*�7�GvN�QX��G��\�"�/�[�u�֍�{��,����6�������۽���r����p>��*���!�[��6�n&���%\�2�)q u��T��)vq�U�/si�ԃ��+[��i������������D+s�[��\��cd	w�Sޭ���Zlh&]Iz���,��v'J1#�]�)�*�o��C���&z�ʭ?0��C\T���){�o7�����@��iII��Z�2^���y�o"�O�G����P}�
D�4C٫r�R�[�}���`0��]�ݘ
��ݦ�]<��̧8�,�2u�.�v=1M���ݬ()�[崇-�����JJ����tז`$5�K�F�Ճ�(H�^mZ�l�\�V7cĪ8iЛhwE�"eE��|�曌*:M-L͏n��N4�C�zY�/x�d��Ya��h��S��,q�7��(p�P�/!8���4��A֕ d{b�+:O�ra�Ѱ^r�u�JKV��֐.q0���Mؼ�/���Dˁ��mm����p���[NPyK�&��Z�A��*i���鵯hY[e�u��\U`���#EK������8+%�yx��\�%��bwr�,*�It�CEܴ����yO��3��юȢ��7�E�n�c�\��%;�Z{�-ZtB��h*��v@��EF��c�߅:;Մ�#Gu�=T��͗��3dU���ef98I����T���3y�'o`pQ��ۑ�k
�9Cj��xU	�4{-ɩKպ��2&-ڢ_v��.�R��k^Z��*�yz���;���4�1�|�� k��W�	t^�]C�ۘ*��=�&p�	��U�� ��$����ڇͻԅᨭ��4x���r��v���Fn�w:���ƞ�-�9���
�fc�إ��Z�
���v���Z�Ȼ݁/q<y
�
W����:�d��Eg]�n:�!ȷ�]5�xm�.���<�@�v�'�uԊ[�r���s`�}᫭wmо�P!k�ڹc��|�R�@El^�q�"���1y"�7��b[|@sTu�b��բ��5��p���mEԺ(I#7~\;^	+M�4p@�M�V���W|����ae=�Es-m��ĕ�u(����K�N��LV
�tm�x��O�>nٴ�n\r��-�-wٮ��z]\��*d����!���Č�ό�#;D6@�g��1ٟlH���[�����u-�*MҜ}\����2o`̕�J��+]=�3u{�$_Ɯyhjw\Đ@q����I
�j͛k���8���񎳵�w�U�&�$K݂*�|��|t̒�F<��ٺ/b:�j0���pa*(�I��ש
N��тN��d3�ᇉ���}	�&5�s��]�˭X�H��S��2��F�\��i��G��6yʮ}��迕��Z��q��<�[�p]��
)�8,װ]Z&V��!��)�A�b��[,�93*��W����R�����F���[�4�/��Vy��O#{hԐoJ��vrgy� u�8u|�3��f_U�	n*za7��ҭ�{0�:����^R��S��=g�v��w�eke�%q$���G�<��O��s��빩����[�5�Ih����)�jfa�������W�IS7�%q�	���7�s^l��k����Q桅D�X{Ce�{��ڸ0�z1����1Ne)��כ���+����_O�	�[;iz򖌸C�N���Dqʄ�<����gT����MH�l�������6*�v[���2ɌO\[{�&Sr����]C�6�B�W�Et�&H�f��d���ֱ���٥����ӽ2�K1^�z�Ac��+�<�IW�6�;����:�E�y�ق�q�Ն�˛tӽ�z�0s%k ;jK�E3�z�>ӽ��X}Snq�eS�,Ӝ�a��a��
��l�$Y��}�7:�yA�7�z�=�:��&Rݎ5gx2`���h�d��;J�1B�x��o9�H��y,8�idӜ�b�N$�g@4�޾�ݏ��]Lդ��BoR�U����Neu�ԅJ�淎�W�14���ymS�K����V�4�-6��B���Hi�SJ��2�\��t�����/�z�8�OX+�����H��J=�	����W1-_�)d9׽-��'v)5��$
z]��f�v�m�5kd�*��4�Ͳ�[�zR���M֭�.�K����Jf_]Hn�Z;wz&��7a�� +K\�V�=���|�����PQ�|;
u��|*����ێ5Kf|�.C�:hR%�!|v�0��t	X�6MT�1� ��źk�Tz�l�r_V����7��W�%�mp�O�����#���b��٦}�1'������l)3יu��۷Ɩ<	�Z���f���'���Շ.lX��w�)����x��H%[!��V����A�	�^��q����Ds��� �Yf�LZ��',NC�0��9NjeR�>ګ�����u+ih���2N���lZ�Y*QZ�y
�����1G� y�wX�$abcƑ��b3s��T��H<�<�ʻ��$q<X�I$�I$�I$�I$�I$�I$�I$�Igq�u��C�f���I�,�[SX�r��
cv�,6�����A�į;0ݴ��ӧf/����Ɵ˶»�*��ڒwiD�}n������AqS_&�'p��\�9����䦑�n��O�m˛�w�/ѕ����S�[����/_E˲T^o;����F�3N8�\�]Ǭǆ'2���{%K�l�3h��F٬���tK��T�J&������9�nPt�*B0���8�n^��r�r��ֽX��޽�U��J��]7F�9�- ��r�8��V#�,�&W5�v�N7��Čޗ�n95>l�K����]��ZT�]�'v��oe=�f����AYJɧ,�b�q���d��Io�i�f�<5�]:�I��cgv;u���4P���d@���8_Er�H�G�#�Z���h�w��$�mgF���nlvPX�t��_�?����~(?�~��-�n����D_lS,o�d"DF�k�H�h٫r����"$��������������#V@x���u���V�V\��M)[r�Y��5��f`q�0���`�E����YL�D��1B.�� )�Qͬ��R���,�S�Һ:�?ph������R�p�W��v9lgG�����vG��,��a v�W�+�B�Tk:Z�ղY}tJ3e�9��e! �q��ک((-L���R"�u�ͥ}{�cΖN����-�y�)ˮ���b���)�H����_�*��;t��;[Vu'���S[voG6���_[�nf�Fi���sc��k�t���7$J�MQ��ԗ��$�vEe��qon�1�٥�,t�?_��,Ӳ(<O�D���Ib`=GU��� <&�z'�n��!����f��v]gq�@� ��n����JgV��tQRTy*��V��;N:}��vu��Cja���<B�3/E��0(۸��/U����ۊ�9}"�1u�6u��Zy5�\�ù�`XUNtS�a�E��XY]���][H���6	t��1b���?зtj���!D���l�햹mo#.Z��''i:#ňg[S2�]C޵*�}F����[ɛ�1b͝��4���Ka.Zt���]j���N�����d�2Ȋ�T֊���nfWE�r���pZX�B�zu�E2i*[e达�kx�zl�nYΔP\�t���/��������Z���E`P�W�a�ƹjz�M�(9��7��Z��́Z{�%Xֲ*!sˌʺ-I1X
�} ��}w��(
�2��8F��a�m�M>˩�i�A{Wp[5xkb)�Jy�+��rZ|U�H�C�,�Ɛ��lWb�=r��e<��G���q��e���e�ր�Ǻ^P;����F��ա�����,}���b[�t�H��)j�.�[�&}���v�PѨ�/��]1,z��ch�#@!�W�pg�������h�69�\7R  F�l��SN}�P}B�`n�%s䫢[̽�7�����VIA�ț�"�� k�Q��TAtmR
�.���ܹ��I���k*]�2%f˲d��F>���\�N�B�`�!
��n���@a��%Ved8 
��.���&P\%까��K�6�t�Lk���˒�$V`���\N��L����M��h���'&<�m�!fș;�K_б:�ݤ�v�fӫ��|%��U1E������@<c4� ��V���uZ h��|>�I���*�X;��{9�mM�3��ӄ�6˕�_؅�������QM)B�*��
B�bL��h)��@���0L�Hҭe�=���J�z��vz0��CL��B�I(���o��sT|6�@�Eew>���LXc��u��(T�r-A�:��.�����L7�%25R�t�TU[Dܶ�1���ը�ʸ��q�m���P�a	Es��`����%[�eF�9kh��݃.�Y������N��f*� V�/�|�vQ�:��\������l�����CR�|UY���ڱ���<�K+1��\\�c��*��C5]V��&ެ׵ҞY�5`n��Y��� !C�d���h=��'�'v3TkcMB�HQ��7�/��ysqU��5Ϥ�B��R<�;�l�F#�`K���5�f�؄nG}���º�4��]�b#λU]�Mj���.��]����V�XՉ�kn�e*��uLy�\[bK12k\�2%���dǓ���^ޤt]i��r��L\�.��3�MvE�qrF��[7��j��I��W�4ik7����}l��0���KTQ�(P��l4�۳~��d�7��r�#F�CNd���g%��5̒вR�VQ��Ď	+E*t�����n�ֺ�`��ce����3�K�,�F-Ab��5���ZFud�K��$Et�\-���n����9�,(�Yj[���ش[�'���QI�[ѓڐ�D����_is07��ȧ9���/6R#76��;w-�����J�Dz�kR�oC���t:K5�+T�F�z��R�D|4٥�|��$�����ٟ��5�r�un,����+���r	�)��8��{ڈW��S���OmU��U� �E���%b�'���s�7m4�$a��Ԭ�7��Y��G��@6V��(�# ��}��j�	(s���eby�&�Nd�YM%\�`�Wn�����,ǈ����ds��c	�n��h޻Ha[0]������F$�v�\4�t�]��]tj\o�yIZx������!Ҳ�b�7m��J��3�I���b|�y���F�Nb�;��v��顆��3u�R� ���GS�dKH�}tMdj�X�r�r�m�٩6-�,�4���:r����C��ݕ��c�h�v��G`K1֗1��3m%������5�e�,̡��y��m�5�:���Qt%�g�
�lS�L:�ݍ<U@!ܙx�ei��n* �ܛ��80��d-\�d�Z�"甜�m��E_ˉf�7V0]bw6���3_�Tg���o\�TU�	8���ҔR�ʗ���	�D��o_-�ptU�@ݐ��F�JŻZWQ���F�Y�O��T���f0��v�VTw�L�+�}�Z���('S@�c-�hWp�rGAUԣ���]}�T���.�nd����2��kG^���s�Em`��%��e�V	Pc�W��������gZf�,X�C�s��� �I� 9�qm�w�g��2��6�M�V�7.Ƹu�1�	r���Sd�B����%^�Ueb�q5.�Pd�]ʆ�����p0���sڊ`��h�z�+�f���Um�r��}����ܵ��vі�K��E�5淚�ZG��ZP� �v��q��w�q�4N{�cWmb����]
K1(�j����%�v2�S�\㫶hWˎnZHSڽ�"�e��V�Cv���M�7���`�ehJ����$�,�M�Y��-�:�[A���/���Q�{�bV�U+V����Z����X���m��]vܛ�v(�5]��ƺ�o��g���km�0"T��/��T4٢1a0S��fu+�;�3P�LW1b���-��En�l�f�$�����Ŏ�G6��WSom�ՠGYfZa���ُe�\�����|�AFg1њI�O�����Ǒ�n����/e��+2�\cT�39�J����tW_%��-��B��v�O9�ӹ�ә�:_U���M�s��urI��²Ma�*[�u�����5h,���4��w��ѯ_agI6��+\o���t����.��rΖJ�˙ܩ����%��(k�0|�c-�[�2nV��ՆG�⩣f];݃�x��RI>8Xz=b�U�[��3Z�9-�L`g���g*t���N���Oܢ�ml��Ma� 9{���X��R���0s&�SN���T�#����Ut����p�`k!˸4���5
�.7C��[:��ڶ��ݡZL撘\�Zܺ���:��i84:8&4*,��"�rT�6��lxG:`��`Ҳ[��*n�A&i_�'�2����}3v��ԭ$%�4=M+�[Y�Q[��:q��
7��U��E�"#�P\n�#]�v��^cӵw�?�Ie�W��>ut� ��Bs�������y�����^:;�v�%Cn�!���;��-Xլ����ע��0�U�;
"ʩ�N�ɐ%3tb9m�T�Z7��/[�,�lةbE�d��[+�N<��gUnud]�6$w�:�r� �#�m7�^�̤�@'x��lƋ!�̺*�����]���f�Z�EoM�XT��oQU�j	ˤihVn#O�&(nf>��7�6������+ɷwyKno*�O"55�ȕ�٨�C��j]Õ����GZmm]!��b��
�Vp����0T���h+�ͫ�� �7�HWk�� d�D`]YJH,L�m^
y�7]=ƶQ+��]��s� ڍ����y�*��h6]r�ש7 �TA�ܕ�l����x*�P�k��o�2.��-+��cp��{�a�l�m9w��,YU�Pџp���X֦%�4J���I���vi,�j+̭&Uue!�Ʒm��('\HQZ�4���5�C�B��n�)�r��b���V��H,s:E
��
ϸ62�[9*�j�����^s���i�L��T+I���95u�
���*�SQ]Y��Q|�M"�P%m˷v�/Fm���:���p�r�[wS7oQ;A���+�*]
רأB�e��
m;�͠6�$��X�V���v���FZ7�|��O���n>F�	K�k�����_%���#�O
�yi���nd��>��xQ�unZ�4	(v���2�C�8#z�/(�']����H�V�4��'&���լ'�!�-�pT�V�Pe�[����g1�,��bج8U�rxr�����^4n�2�g����ȓy6됼�r�<��Mv���Vz<����հ�k���w{��/���xJ8��(��0��&�U���켧Ρ�V�J$e��۹)�z�Uyişm�@���46:xU�mMi�F���U&��0��V�9����U����~J��[gku9�u��� ��H���b|�l��K7WOj\4��`V|���Kw�Z4&�L,��M�j�S����{A+lB�[�����m���2�F���޻�� ;@v
u,�W�[j�AZfGt��W[D��:���a�o2�]�YDL\�h3V���a,v��l�w�;v�*I������.7��v~	�$��B"�+��?)<x���4`�`a-�{�7j�S7}����^~�=�� s�M9��˷I��m묑>���ZDӼ�+�WS���Ŝԑ�jQ�AD<!mk�y���A'K��R6x%� �ۢ���9���#�9�f�p����e���� �\���4�Z/Y������[���b�� y��'FPJ�<�p��+0�z����4�ݍ �ѽ��3��ˬWsk$Χ�XZ�Q��b��7%�4U�r3[�+��:v䣳y�?U�޽s�P�A�b�J"����µ�K�mY��S�u5*3DZS{F2��&�oY�]
N�ӃY��df3�+��:�q�7������;m�qe�|w9��\�Mi̭�(��o&J��L#�CC��N�ks�����;�S
M�`u��n͸B=԰��	�z��~[Y�ǯ�@����&���R�'��0rQ0����Й��MoNEIBTY�U𮃗E��P%�Ҍ�۸$��o�r0��˧Ƿ���/�ߞ�+�<�~�p���UH�EUU
�Q"	F�
���Ihږԥ����������L�b�E#mGTGm�����b�ډT�X2�J����*��ᢪ�iD�R�g�����E�Bڨ4��XҭeS��ciEK�R�%+V"�������Ƶ`���J�KHڢ,T��R����lZ �Z-AA�kj�-J��a�.+KJU[h%F�Q��Z���օj�*5R���b��[jԱh�J�j��%�F�֋[DX���cj�Z���2�4i[�(�\�ËAU���[F��M�}忦^�o���-_]q=_�'㵹��aF`���@�#�hr�k.I�5�:��4���wiN]���w��L�����ʥxU����n;�c:#�v"R�1���vK���Ps(I���
P_yB�����ۮ�teJ�h��qHOS�����5�Y{����A�S�7ێ`x�$�	]J�o5����M���*5��î���Tg�v׮� ���<+^F7=7�¶_!#A���(ń�fR�f�]-�"�i_V��i@��p��b�I*h\/(.�W���"辝�.�y܍�A�|��#�D뙣� ��	ɝ}X�>6�W��lj�wdJ8}����ðcun��c����6�zxjYo��JS#c#b���^u{W��Nt��=�g��wW׮�"�9�w5:����i�b�i>�+��ꋑ��Y�����eG�F�*j�I��}�Ҝ�f1Mp����5�iI,Ham�ic��WU���<�P���n��EI�{kKg������iM�1R�[���T�r*ţ|�޿az�|�w�ߡ��̭+�`-��U��[\\z��P�WC��)KTW��4k]^���sN���#���Ʀw����X/�z+mt<�G��N����>�U��{ ԫ�������
Jf��4�S2����E���}����~��Jr|R��\����2�r��m.��B�m{�'
c�e��&"g�p9��#FV�k�IT.�r��F���*�[�O�#��)��	W��%L]�jr/��sx\�s8Z� ��d�t�bW@	����v`e)�:��d�:.�qY��H�a"i�[f�bբ�Y6�� �@�e�]ȡ��[�a��� �+3;�5xRP;��]P�$i�v�8c�&1.Qw���v;�yqs����NrΓt�7�G�Ŗi�nf�|P$ѸM����ʯ<F��sXz/u[��������������8�޼�毧&j5E�z�#X�J�s{�O(��^
�[3Z���J[{�Z�P~=�9��δ^�z��fD.o�έ�i8�t�^roWk���&�:1�,3���[���"�lP	��&��^��������z�7�X��wTi�3P<��i��&1wrR�l����^�H��Ƽʫ�#�l?/J��7Oy�n���^u�Z4�#tVY�cji7Z���:��/�^��W!��嚵�7�n�P�O�;}u)=�	�*�+j�v�κ�ڂ������W�W$�n�p��L�}��B�I�����V�2��2�Q̤7����'�B)}됑i�$��y@�f3u���e�m(,�u��݉��*���4]�R���Ԏ�+�LVM�<T�;�O�I��=
�$��7`���`����۠-	c��٭ǚ����E/k���F,�#�5����*�����-oLC=��Ct��I&/(Bu��o1q��I������rBAe�:�7���ą��멙��k��+
j�&:�]���m6v����`܄�R�E%���g�bz�{�����o�=�!��V�d�8���Xd7������IzTr�Cc����6��ZX0���F��!��#��N�-cɾW�J�ޕe�rj�u�Nmw@�/j<�	z�b#k��OE��SPd�$ ��9��#��|�J+��r*{��j��k+�IO�x��>���Q�,'��idE[����h�Z䖉�}�����Fv�=R���f
�9��۰�{�~���|�b�5�4m��K��.���7攒I�}��ޣ��Xsc�/~��a���^�&�����^*�VŔ\�p���K-��I��]����z�F񤜅U��ў�(au�Dr��B+���75ie�q���_�f�;>�Az�1�J�����Cxy�ֱ7�ݦ���!�*��������6U��CTyE�8�F� �6�y���EPN�y��t���u�Ju�twtT77u��tM���TZ�؂�d�	+U�$���EÜ��,X:� ����.�o�%���)���8#I�s�M&���s,���6r��;�}�.��d� w��|'��2��ܯ�r�@�S���ϮF��$�=Z����qջa�c�M�]0u�V4�C:$d���<}�Mx�l^��+8z��	cΎz{�\�՝�yo�d�ܼ��
u���}��t1c5θ��O,Mk�p���I�Kȳ�ܼ�ѽ�֔�8��y��^�'��c�L���ܔM�6�#5V5��cU;ɞ��p�w=���?��WC��S{<tYhg"�Z/Ƹ��LA����n��)Mf�'lճ��p��$��C�5�׶/��9��g�9e��PŠ[t���Ix�Ŗ�ۻ��GX�2+ÍVZB ��A�k �;r�ī(�ᓷZU5��f�IG�U�u���c�g���4����:�S^�����;�8�^r%`撤��I\nW[�Cg.�מ��%�wT���=���C�pZ�.�ȼ-LվB�r�'�6O/����	Rbb�Yi�᣶����U��y�nEU=r,�Hb-!p6��K�8%4�]�^Qt���{�a?d����HtEp2	�68�ˆt�H^Ű��Gv<���=}v��8�=ίP�-���N�܅D^P�[�s�<F�sZ83"Ke"�d�r���Oooe�t�9���=z�m�i�ө;0�-�\^�	�g4!�WUK.��Y�T�i����(���/�\�t�a�t�$P!M5�ۋ�$���m_h��O:LqG*��� ��ӧGՊ$��xP�S�狡�|.254djM�D��I�9D�ɰV�;�r�ybqQ�1㊄>Ŏ��r�<c�g��t�&���b+�(�~6hF���킝�V�����jqg��o%.�h~Nʎ�}B4��C�;�s��;�����T���G>5MH������7�V��U3|�2�l�Z�-+���W�QG��zĕB�.�$M�Ά�iK��r�j�0����I�'j��;���~�7$y�Vk����6�2����?��M&B�s�-�^gT��v=~u�|7��v�9��;[N��;�Ʃp�t-	��!��B�w�coY��`��=��1a0��
���;*���j�I}����R'Y",��-m�Y,�K)��.ਜ਼�������ځ-���c"�I䮴C���	��FF}���ƺ�n��\��B�=�v=؛���	�e��4ܓ��;\#��)���O>҈{c��V�o� ���>8�C܊���gke�
�*k,�UϒP)��]�Y��M�.���J��^W���r�e�����s���Ʒ��,�"���Zjl���eF,����B��-o��+{ĒrH#[6x����V��PK��DO��~�w5cn$�Ex��J�Q�y�:�K\~Et͉dǉ?z��=>��`Sֹ��6j+�Thہ�s*�OtK�{��:�x	����z��W]�I�wԾ�DSG�z�?r�m>��v���3ܸAK�Hu2��|�����ܺwZ9����z��x��:t��i��P{�"��;}h��5����UJ�Z�go���i��[��yh��"��R�
��pII�<�gah����5��ʓdb�R#X�F�=[a����1D�q�^�[Q&�� �@��\s�X���Χjo�C��#9b��L�_���eɡ�_�uԞ�U]�v��p�,���Q<e����)�K��TY�߯�v^��1��8(>���C���+����1���l�՗��|K"u����캻J�o�M�>]��SaI�s�Ygf��F:MAV�i�p*k�vE�U*f�/)�U���N�-�l��ޘ���֛қ��X\[N�nFU͈�L�s��S�s��I�ڞ�i:�:}�~�\}f��%�M04~��"������t�꼼�'���	�������:�ukf�vFC����f�n32� 'y�����X�����٬CQ�K�)ҚΥ��:�T"��[���4��ǹG4��^Ѵ*s^s-:���� ���H��� sm�.��@���zF��J�wI�A%E�ye�4�gk����'e��:�4��5;�y6J�P��(f: ^;�2b�ܽ#I�w2]	�_>Z�h��[�6�F��d��*[b�ڰ�������_O�0�oE�(X�"�5n�@F;]5u�u���kN[+U��f��r��#5�ћ�8=��H�f��"Y��W���ŷi�/�}j�j�,2���j@1�5v+���5�AW�_j�]��<B	�Ft�]4ڡj�m�y`{�$����MԐޗ���7K��O�]ڣ*�u_pXTj��+��1�1ಳ�e^���@M�����<��~N��E��ɷ}�WԒ�=@����mJ훴V�VsBq�a���Á�j�*:����\n��ܵ�	MZV����
���"��3I��Q���#��+��ǳ6'�V_mKC��7�}uX"��j�z���N��ܙv�`v87rK��Iv��B[LΥ����4�WN��dq,=��unX�è0��vZ�W��6bѴ��bK_=;C�5�'/F�iq99��4�m.$�_�}AJ�w��{B��ʂ#Q�=�I���7�Lmn�4긑�\�	|��wQ�,әVԼ��i�<�t�B�|�	��n���#:�Wg	G���C�h�d�2C/rS�3��1R�d*�V�`��=��H��	����-XRBf���4D��2/��z"�K�H�c.����L����ѣm�]�q���b=6��l!�MB�:�6��+
��*A�� =Kr�j�8�"�(8�$���-º���[z�����JDh�ť�qG��uTE�t9Y*۠��z�(��Io��ɦ��P���a��MoN�J�M�a��ʜ��Vm�� �؈�s�n���-�)�]`p_sp��W��]� c��!l��k+KX!ZV��Z�bʕ����UE*����D��F��-���fV
-J�a�(��Z�[o�G�2#X	J��l���h�KDKmA�mQb%im�Q�ʱ*��J�JZ1�Ҡ�Q[J�ŋR�Q�*��h�kK(Ԗ��G6�IE(�Dm+��E��%J[*T��0�[B��Z���8(���`ƵV�5F�kږ�J5Q��meQ%`����*YR�X[A-�KX�m�cmF(�F�J֍�e��(�
ʅ�h��j�KmB�j7.0�hږ�����jP�JR��ED��!J�J��0�Z�VQ�mR�elKV��&)b8�֥UiZV�Ÿ�V���ưVԣC�V���j(֪+U�ұF��F���(�E�H)X#m��+�.���ߟ��KG�N�M?n���2@������o�7M�u��Z��U`�+��LX��d��H���0�	�q޼/_w$����z�wwY�W7Bm���'k�y��_*/y|~:��Z�����U���'Oʄƍp5P��_^�?k�����ڸ�s���l���5�9Fq�;]��w�sRȡj�[I�U��u2�"���+��W�Mlea{��l:ޅ���o�nq[�ؚ�%H%
�P�Ԯ��8�4Eq%��Wcʸw�,z�MW��N�(�ܠ��(���Ȇ���H�+O�eۭ�u*c� ��6�`~ց� ����G>�r�,WH�N���1#�,�[
&:��Z�i�a�Q���h8��B�Ss�"��ث!�׋>1:���mؑ�\,��Yw��^vaVH�!ǴomWH�3c�����eڒ���*+�^�m��R�U�yЋ��Ρqf��"�r�����T�t�c�@}�5��շ��l�MeS�p�wH�W=��������5�"J�N�Y�_�v�u.ޥw3�P,��3�����y<�ΡsS�E��\�F*oKP)^�o�^��&��_.y��1��
I�1ϖ�Z��{�(�p�=�97��8��>{��uu���Mv�C����F臨wd�(��H���m;���x?c�]��ᧃ��g���ק�;Vn8wu������1*�zC�3v�VΜ��xb[��v�!r~�ݮ9�S<�TP�8�_C~H���K��t-�O9�Pc됶Q،?n��4�|Y�%� �z��Fm,�1��W3+�:#\�]�_)D!!�^�d6:�|;a�/[�؃�o5/gZp�q�{����ݘ�N��88��{4YI''oi�ά#�+�1��n���"d����U��;ɔA����g����1��D-{��]���]�QoѮ�q��Ϯ���Bx�B���u����)�
y��Py^N��;7A{r��{JJ�&�s:t�1+�:WC*J�&a5�4*�Q�x)��u��]f��OH�EXXk�3{{,�iV���=�"�fF�c�������z��_������1"�}ƽu�a����9,���;����4Լ����&��(�5SSHMot_��8�;N�2M��;L��^{�w�o߷��d�	���<x�ӖM���N$=����!�m�$�O3I8͆�l�Y4��.�q��u�.~[tZA��\wd�S�FۢE�U�v,![ړ�%���4��ߋ*wd�^?�_`��'b�		�s������䳟!Zܔ	Y�8���e�!�L������� q���ІwN$��	���$�&Oi8�|̜�	�C�H�0RC��=a�}�L2M?g��g���>���Ӑ�&Y��N2|���ha<}a4��ө>z�xr�i:ɟi8�<�1!P������m$�����ޝ���^{���fvI�Y� L��&���:ɶM0�����gt����N�8�f�z̤ά��
U��`6����P�+��m�{�'}�|�L���(C���k$�x��N�Y����q`q�Ƭ��ՓI���6�^z����~��̓(w|�d�wx��LM�O�4�ɛ	��>��RP�J��{�d�a�O�*hǗɬbߵ����;���hN��L������I3��J��2�m�L�r��|��_XM0�$�Y:��,E	��nﯷu5����EG�i���4�q�� �&��l3u��Py�H�k���&�>O�P�`q3<���@�=����y�uܜ��x�wW�IYP��R�N�`d�!���
M�w����ĕ�sVE�LKa�����6{ܮ�߹�}�|�vC�C��4��&�L!<�x��ԛd�1>�XC�e'
@8ɽ�$�@֩+�$�8������~����>�:Ì��d�!�&S�a	Ğ�d0�i��$���!�x}M0&���d�Ow`zɦLoO|�����;�~[�}|´�0l"��}�}�� iܦ�}�� �W0���b//�0 ~�,����N�S�]GNrI#d�#;}�1��5)Iᚭ`&�8IXJS6N.H�x|�)��y;dRz퀤S�����6d6��OP�!�ԁ�75a�I������0=�D鋋��[��;�����z�=����>d�&y�d����`�8d�!=O�4�<eMv���d6��;Bq��'�'�6�~�c~�}��M$S�M�0�7M2u���r�����~k$�06ȡ<C�S�x���L�Rhzw�c������i�m'
t� z���ԓl>��i8��|��O2jrɶI��s0�Hyh|ʄ��a0�SL�Hq=��q��k�������$<{�`,j��4��=d6ɶ��_�:�i>t�x�:�笞��'9�Bu �,��1���Wr33KωD?����B�x��Y0�:�4��<��N�w�2d��SI'3�u'ΘO')&�����$�������2:��{���o���!߬����I���ԛL��I�C��r�(m�L�CR@��:I8ɣ6P�{�}�{�>���rt�i�M2����	�Vm
�ii4���!��,4ԓl��:��,�Re��6�\�/\s.�{�|�u��L&�;�M3(M8@+'���I�2o|�!�ӌ+d���4ɴ�'4�aְ��%}d3����xv�����0��M<aRC�6�m�d6ϙ!�N���@���
I��+'�['4�����N2i���ϟ��'��^nI��&7f0h��Wס��S�I}�ϓ5�ۺ|_�ͳ)���q�.�4�/ҁz_��0:�Og%�g%k5oD�.�.�-ܼ�2Ǩ����lǱL���H:R��uYu��a�vI^��
q���6�=�f�X(m��3����I4���=0&��t�D{� +p�a�}�9|�;'<d�w'�3>Y��I�<=�8�x�T�<�����$6��v
I1�AI��eB�/;������_}����+��n��|@��$�OSN����l2v��d<x��I�IS�qc�2�l��c8޵��H)>d��IY1���+�$�VE'���`i'�Sٛ$)�z�a6�L�d7���!�I��|�����s�9�o����w�2�l�d�v��d�u�y$�'�{�*I���OX
@�:��Hi��i�2�2v��d
{��|,�f�IH~� �9����t�'���:��ԞCv��d�yܒ|�����	'SԓL��d��OY!�w�:q��s�;�<Hql�C�N�Bi'Pɫ$C�u�OO;t���~I�� �O\���I���{�!�2���[�;�7����oG'�fP=I:f��|Ì�yB|��q�d�a���N>��N�I뤜d��=w��Hg�{��c_s<�߷�%a=ga�I�ORM��y��Ll6�XI�2i���2q���d�a���M�����O$�;�9�<�y�������2-��L�:���� q+%I>k2|���C��|C�CL�a��u$�_v?|{��e^2���;�D��?�[��.���{`O#XL��[���`��=#�>��}N�0>UF�ʞ1ˎ�����ו�����a9�3��3R%+AN����`s�\S�G�qp$��� d϶d�&{�3$3�:�Hi&K`q03l��L�ɄC��C����� 	#�ՙ�잼�^ q�{~}I4���~;a>fY2n�lk9��O��*����`#$�M�Xm�q�غ�8�r�������w��2e�ABm&_P�Ł�gW�C&,�N��p�VOP�I�37�fB�3�"�Y.�a�&���{^���w���}���%d�z��d�g|��O���x�b��ӨN02R|̰�	�6��(m�1ky����������~ϛ�5�w�+'�Y;�	�O\&L�N2|���I'ϔ8��!3=����Y'�Vɻ p<x�P�{��n����r��>�I��f�dՑd��8���6�<�q<C�&����.�Jʆ;@�$�+!��0�٧\�{�}�;���+	���Y0r�d�I���%d��X�d��I>I���!��(e�@���u	��� P��\�=��~��d�IS����Ձ���Aa�Nr�VO뙒�d�}�"ɦÌ���{�$0��P�I�;���e�����w���3�CI&P�O�6�|ΰCöe'6����N2`�1�$�&�d�'��)<}`f�r ���>0�g`���Yp>�'S):�z���{I=C�:�g��d>��8ɷ�8���w�Ƒ��C���eD��������6���i�"�bu;���H.�;aӡѝӪ�o����"+�]�f�մ�3�sAʝi�z��8b#Z툸�\�R�5�5-mZc0��^�F;��m{�?j�A�7���9���񀡄�L��R0��2d���u������fj�'�϶m�L&{M2m���8�q=�L��O
�OʑI!��=��>({���,���C6Ͱ1��&&~�u����Cl1���|�@4Á���{>md�,;%���C��ި��=4���<��d���6�	�7d=fX��8�'���I��0�|�L�J��0����_�w���;�n�&�vn�2m���Rx�]�m ��q ��*�ԇ�6�m�����f�l��y}�>�߸מc�y���&��C�������:��L'��l�����I�>�<�M�
E������>��=a�^޳�|���	�I�Xq�����&�6���Hw4����'�4�O���r�i:��N0C��2	�q
�|�^8��͙���}޻��O�6�,�@6�<��'=��6ɦy9�K���Uqȭ��ټ~$��\1��Z��޽��sk����ʼx�vޔ��R�8��铖�S��.��n��dۊ�l�R��Be����4��Ub�p��/�Wu��g!��h-�0�I3\�f�G��!�oMԗ_q�Xt����ꍱ��|��V��>�N5�t����R��eѷ�r�[N7"?�wa�]s�_�x ]6y7>?���-�������R�[mr���<ϱy&����]شl"'�jl�XA��5M�ǈ�8�b^�2E�wf`�	J7(�Y7�S毢ȭqΊ��;�i��xOQ1��,�,F�K��{*��1`Ȅ��nCZVZ���[k�7�*ϦG���l������hA�{�� ��3�iɡI���=�OQ�u³j�2c��b��tR)p6umr;�~;Gܶ0�{f�(�nU�p��o�S�����Ry�i=�;ׅ���	7���ubEױ�Tc����)�jU|�������E|����u/i�0^��z�֊ۣ\e��/`$��3�G���?�������+_�i1�z���b�sh(��C+����&���*�t�.��ާ���aw瓺�P���z�u�yߵ:;�M�j�{���b~�դ�>�/)z�_CQ[��?C���X�����g�O�U ��u2T\r�ODY[�gL���?5�B�G61�j�W�B�GT.u"W.nT����=P}��M�Lx,��麶����+��as�nyU�,{j �GH\9����è�z�W<����18�D횾��mbd?0tŲc/��=kj�7�j����V�;��~Lm�L��yup܅@�����P����a<�r3I�f�G%zi��ϕr��>����Ɠ#�裂����pQu����h&$Ktŗ�3r�+�3!������l����-0��û��o1�.#:J��x����˛F��ju���l3YN����Q��h�{wR����J�8U�.�A�l2j��Kx��ђ$�n��X�3�41�ԋ�X:��3����N�J����P�Lܲrۤ��c5N-#��е�bś�о��s�Jv2IJ��C4�&hI�wnaxy���Q@W��"냆��Cyr0��:�)z.g��x;��wƦL���PvI�}�����:n���a�`63	��������@�wHF1n�)Lyr<x�N������X�Dݲ]z�[%�r��5u�)�M��xc�9�z�:�Ժ̕;gsX�X��:}��g9��������/�+	L{6�BJ#��D�A��r����;�Z�gwZKv�e����c����hc,���D�鰽E�;n��׻��Ӷ��IVL}�J�S:Z�7�/8���a���u�[}�� �Vn�P��o�!�J���s���d��b��cfk��q�,9���X4����:�߷�㣎�$i��vF��|2a�:���h9Ro@����ù�y���D��wRu�q ��y/7B�F<g�՚j�Ãe��0����e2A�	���\�7R������)Z��V%�=�\��������j�?��e�5��q�/�*�]���d��R�FWC$�і5U*<�oն�	9Vı0�d@��@\!&��3�q>�I��Fc��.�q�d�I�^k��9����J�[�XW��w�720R�Z�d/rE�����t@�T�=+ |:�]��hi���lt�"��2�i�n�D�v,Ћ��Ga��4]]����4s$��w7.�E@�^����(����`�|�h�)U� ��'hĶv�[�;�f��㢡Kzn���3gj����N.���[P�ݥktnY��MoN�.Y�|�KL:���`�/���(v1&<¡��J�����Z���v=�������T P��m���D�F��R��F�F��j�IR��Q\�Y�d���eJ�*R��km.0`0�bZaEp��Y-�\$�E*"�LҰ\���[b�)[E��P[mdm�����J2��+j��[Tje(3R-
Q���p�F�%���TD�R�8�!EfiEKJbƶŸL �ۆᕨ�W1*�`�W
)Z`L[�6�.*���(�[R�0ˆ�ԩh\�C�1�G��Qp#l���`�iqjT��T�0���6�UfY\V�R�
ʊ-kbX�[khZ%����TJ�*֨��Zn��4*)Z�lZ���R�R�6����X#E���q��Ԣ4J#Z"�AZR�*Q-���+sj�8L.(�eh֭�U�b��B�T@YR��X�QB�.�TL�%����-E&P��PR�h���J��T.�;��c������Ǖ���V%(�Be�X�T�U�Y�kwq3�N�G(�i[�g���޵�Ȧ���yf����t������o���c(ܘ���;�=�y��,Kr+z��
��<U�k��M����I��N��W���:+�Cz��v;�U7�˚��5�3䛸�|���i��0{�����/�>���<{���\u]^�..�9^�Y^��=�B�8�!��Ƭ�.�ou@���t��d�x�.�m���l���@�d=�����xe���E@�=�[�M�]�"�0�������� 6:�b0ˣ��8���^�L��a�7;=�/��\���=�����61͘���pw��u�u�Y�/bB4�ϘoV��cJu�,��i���=z�g��b��=k	xr�?ʛ�W��{�u��5���iDC����%�/��ko�~�_vSLN¨´c��~�� =�ͧ�'�$/׸t�<4��u;yuƼ.�]�,j��j\N3A1$)J$�XGk2�ɢ�V��-H�;r��zG*F, ��&x�͛��u��"�N�SYT3�[�s�O"�,4f͑��o;zk��*�M?0�1�v�c���xy�WжF�ZC��ͭ��p�W�>�Ά�R��dy�� ��=������h�&��^���^��;�sG��7`��y.���ƭ���ud�Ň��!��y���=�+�ũQ�0v����Ors�i��c'hI��e��n��ϱY��Kf�uFf^|ծɚ�=�ͻx���^�6�=���X�ȶޢ��3����zu�,�R�z���룏(�����Q�S�f)�k�f���v!r�[y+D����֗�-�h��+J_� xx{+$��1��;ڬw+N�:u:;��mec�l��]$x�������C�po^��af����'����<+S~�"H�M;�e�z_VV����}�B���랰M���!i�g/��(��h*ht^+�_��B϶�^Vm���rhG(Wî���2��.n���Nk6h]���Y8j�(��K;�{j:��ӟc�7y��\�u�]�1�����nvW�ִ�N�E�)���cg�]�V������{�MЙ������Z��^�"�׃ƯL&`�-{�y�>Y��)/N��	�3z���1������[�Bt���}N�t�ֳ���+B� �F��YI_�Y�u䞘�T�5V�s����#v�~���Wʬ�H��qr�]�ONg�ǓYs��:�W��J��x ����?<�4�k,>.�����/]P�U�QZ�"�
W��
�ϙ�/o^u�Јؽ͊��ɬ۫�Q-�nK�\$�60�ohq����T�axU��l-��Ѻ�ݗ�^s�d���엺��#NuDa�=�1�"uyuP��x����nP�����1L��j}|���{�l/^̖�n����ԅ��t���%P*\���	R~���}�p5&�19s;��z��(A�=i��ES4��I�S��렾ڑV��k��K�yݭȆA�:�[�]�sj"H�l�e�E���V����:'�;���٬əuz�碵/;(ͽ�<= ���Y��j]
|^�����.�0��V��a���ͼ|K�L�ˑ�2h��H�e��$�W��i)������6�ZOڣ�n�H�}=ytiS���{���se�\�!��J$�|/jb�Q8�A�Cwd��u�bo$rY99�cW:�Uk���X��l��}M���fW5yJNzϧ���=����wgw���2�K��8�v.V��Qd�=sZ�"[��x�˔(�/�����|U��v���ú�;;�ūu�q��3��TE֮�M��t���KD���k���:'�T%^�����9\m����T-7��޶�=j�ơ�4�+{̺	ᱫ���@�H�w�}�CQ�#�@st�'�y5u7l���uq�h�th�B���J���vdD����ksE.�&�*U�͔��Z�@<��T�P�$A�p�J���XS�ne���B{���������A$�[�ff����{rUv��T�D���F�v��sT�9~��Y�W۩�p�nΉ�c6mT��qnj䆲ؠTt[�rkݞ���~f���5c����}jE	�!�*;J>��cو
�k�+��V����0xmFU����;=]I1S[E�*�^�·�Ph���b�GH�o?J&��j��ι�zԍ"C�bʒ�h
(�*���;�ɦ�z����d�b�봉�U��#*��|�<Z��lȇ�Xj:��C7�*�[����^s�ʁ?{���[R+Z�a���y9�Tl_M19}���{ dܗ��;�A�v_.�o����� Ϸ$�+	"��gU�Q��+/�8:WA+dYQά����5݇@��'b��vA�[���</	:������:�柎ݛ�]�O,�Q1�r��j��>�$���r
PsVsV'}�fB��65vA/U���VBQ7��p-��=�ckaʥⷜΆLf����k����OqH��(˃�kL�i����/��l[ԋ��z���ύ7dB=z�(����.߻�G�3$�k�k����`��]jy�(��iٳ�?q�D{���
���ϯ�x]AW'��m'�I�"]�*����B�:.ɫk�ˉ�2-xRR*�L'�H�#$�!*)�cxs�׆��F�)~�z����jc�U�yTT���\.��Op�m��2�Q�x%C󻥙ce�����6��g��p*�U�䰕�j4��zt|pԏ%�U�,�y+��yRAڑP��3ԍҟZ8�I�G8���xxW4�$��R�0M佦hu���3T���S$��I&5�i١�2�^T5MMb��:�]y��&��p�����
��Sѧ�H��DY��i�R^5.t���iޖ]�H�w�U����掸�vé�t�
�����^�槖��7�`��W[����\�o]5|��|��k�GzQ���]��X�JTtc�T��	��y��e�!qԱɃ�3����k���&�3����y��_*0VC�"�/�ԟ�n�3�g.��p�΢s��q��7�qX55�ld��v�x��������}��@�J5Dހ�/� ru�zi��r߾af^�r��vc|O��%�->%	������;Q��}|�P8Qh9Vt�z�vU�r>'�#X����B��{�{��l�m������;��KK	E@+O���{o9'B+v��Tn�j�W�j6���e2��b1�].��j7p<Y�3��u���;e��r�HBp�Expۡ+M�Uw��ͨ�*�Θ��n�����Ёfe�AY�Pז(�3A�U���֣��{����)���&/�f�=�rq�/�V�h�E���]L+��)��p�<��ې��^gg\�WJ��I����ݚlc�5�YRs���t�+;��[��"��9�޺ǡ��e�q��H��޶�wl1 dMM����J/���� ����Tz�b�uhW@ח��q3��ˢ�>�/61s�V�8��t,{�B�oz�{��w���wo{����Ԭ�㉉��F���\�J�.�r�)FT�b��bv���!Vj���2��l�W�|�����1>�C�]�e ��V��guv��V���y�,�;Ƽ0�T��R�¸$�c��&U�eWvf���m�*5f^:p�oO�;�q�a��a:�"���k�V����@�)]1�rv}{֣.|�P�_�*UW���";/��v�g�ݲ{��ӕA[�Z��龺"x� F�*��o쾻���פ{H �֗��Z�9SZ0W=DU�*�Z��نmi܎Ĺ6Z�����c�T%�:<�ṋÅ�_�ֽ��L���GA2�L��%8N���uA��R�6}s
���I)��V�/���/��8��@Tu�m�H�^+gD�ue�z���s���Xp��)�Z�ǔFQ
��
�&�:ǿBv��a�M������d�̉�x���1[���-�[�ͺ�*#	����wp�n�X�A��g{��_5}O�=���6�z��0�D���I{\ݶ��A���}���W�C��FeH�Z��]s���+up�Y�6S7���u/�h���o..�/i��n��i!+c9�`6/�(���\7�WQԼx��=^ D�Gt�b��בǈ��ʵ�.pډ���z�gE8�h���`Q֔�B�]@$�N#B�̃PԬ�rKB��*4���9n�Q����h�ȗ��4�!c�Sx w�c0b���V:}/�Ry���9�H�ȫ��ܷ�C̎�`� �u׭NN�.�'��v��쫫pJ*:��S*�+4s��u�P(iz���O��@yE��nn���r�I,�thr[��>KW�t�f	P�^��z��B2�Q���J�X�;
GPm�J��鋫�����W]+�ro	)1��u�`� �ı�ٺ�7�QYGsw\�~�������$�[~Uܺ��탶��bи�����`R�A�iT������>	���5��KrN�F�@����cة.�ЭUl	OR9AM(,�H�:�c��X����'=�.ՎN�K�<�Y�R��j<����֓61W2�Rb��*�%� 	\��
u�p�Ș�B����y���:,���GJ̥|�6�|'J6��X�ü�l��$w8n�x��H��9���&6�T�[�wh���.sA;܅[os��>j�Czs��r|���6��¬*Qȇko��:^�n����z��7w�R̾���M���\=���6n���VW#��rR��}5�X�ںc���0k�� �=�ps
�ΰ�1���ױP���A��8PeƂ��e>�R�gO�����tѷ�t[��|��w6rh;�QI��IM0��{����I���a͛a�n�R����8��o�h�c$&�����NnVMa�_l	2�������� ��1M*\
Z�����-`�%j��T���A�R��բ���,H�H�V��"[�
�2�e��6�)e*,�!Qa\!R\`�m�(��
�VZTPF�+i@XT����Q�clF+�*��TR�PPKn1p�m�UFVV�Q��(��F9�Ä-��eH��QYm��J�U�FҪAj�AJ�`��(UG6a��c���AkЭeH���1PY**�A)�%�J��*B�**�R1R,�(�+	R1�,�E��Zŀ�L-���b�IPCeE+)R,�l�3ha+��*��)U�B����H�ʄ�hR�%C)�YU��`�+P��*���g���}�~�W6��e����'v��P1�)��&�'A['
<nT���+�=�=��Z-��׮Ej��[r,d�
J����������e>�_�4�v�۽6NR�R�,�{�0��~U}(@.S��3�.B�%vr(d�B}B��#���V_��`�^��D�����	��f�>J	��<������ٚ��" (��j3d�e7j�s�o,�U�0�u�a9eGJ�9�	EQهF�J�>��TFX*�E�^����ι��
8��aT�\�����ڌ��Lt(0�v��WW��s�۱6�jF��"���I��ŗ\gT�بm��h�"��s}�Xz���=	��E*/kDx�m�R��>R\лB���	M�*���*g��z GC�F�8��9/�
l�x2�eG�:�F
ת�������o��<��{���G�n��Ld?��m�8�^��@'�k�c^%խ"V+R��ns���.6�
c�[WY���I���V�u��(S�Ý�`JW�S�[��Cp^.�GM�H�]�
�2�����Y�˛t+`����GÉ��*8�P��݃�c\P��+�-ؚ�����m��u�:5*��@؀�*�g�9�ON���$+=�ƫU3Î1W��F�.����^�Dy�����3g
�*P��-��˧VoƮN}PМ�b���F�jlp�x�[@�7���@�q�8��]m�,1�`2��n��ܻK���MІ碸��NHu�~��_]":�7�H����d^׭��ECܨ����S����ΛCn�~u[���,�zE,��{FT�:K
�Ѫ��rc��1Vm_Fjѕ��рu���n�)�=�^�5����!�J����7^���|>{�gK˔o��g)�퍆&z6�8�Y� �g��{�;�N14!���K1�֞rpč�6�E����C�M�^i���J��޶�f��C6o���.�E�e�s]T2I�������+x=d�ªn�wN��J�+H��)iK��x jG�c�t|&|M�
�h�j�� �5�0O{]h��B�R�ǺNrj��ͭ��S�&b6"�)�UGEҮ�����P�%x���f���v%a��!F�Ә����+�r�䴺�e��-"�AcW�������hn����"7�*�WT�^v �\��
!Vw.�����(��R&45JR
��Z��S�{��Ua���QB�g+vT>u089p�j�	�ӡ�����"S@و93=��'Ip�X&5㊞テ`J� ��vz;����Jo��7T4s��8�a��K�0���^��T���<�M@�B���a�
<�\��Rٺ0^[|)|�A�����.������¸P���G�\@T���u�E�	�����t�����q��	o�޻ђr4�T�`�sjj�@����v�nq:��nm�9u�6u!�˖�% 7�����q9[]�)��P]���c:��Iޔs`0��e2�2Oʯ����Yⓑ��|�vH�;��n�K��E����C�T�ok3*��������<n�8+�j&��	�e�j�=f�yb������L�@�V��<p�K��Z<9«<g���/f�YZn��z��� �E�pџa�I��,��k�[V�=���ܣ@ũ��L{��lz"�*�<�P*�DP�P`�koy(�Q�V��FB2:68�FY�܃	�q8t�
����2ȡy�e�'�5Am̳*;pm�Qx�ũҔ��N:�	������Q�!�zOL��}�.����<A�={��k?r�XˑR���[q��^9��ʌ#���H���ZdӲу��tD���(?+>�.v����d@ �\<�PΌ8z�Y�*���\Z���^A�����Y���2r����k3�3��5 E�p��dL��3Nݫ-q,�-��3p>Ä���z��z����ÑS+fN���$�%|
��E}�x|����}R�GH}���[��trK��ؼ8X��>�U�t�m����}�@u)б����������-��U�^��;,�Q<�L��u/���D�~�/Qഁ�::����z�Q�"����n�.��I.����t�ޗU|�9QU�~Wr7�ĺ�Y�l�"�9�)]�U�_�3Ef��6�0�ew*Y�'p���3D��=���pdÑ�:���w/�W7Ƒ�L���K�j���q{gNT���������~#��ev����=h�m{��.~bZK�z:)��`W������kGFy�ᓽ7�T"���҈ơ	!MYK�r-�c�Ƙ�j�8���������vdt�Δ���@=Ty7�!1P�������Z����^��fyS�=S 儘�j�!��p���0<�\�6-���К4'(4�1Np�&v4;�!�٩�LD8�+���uuۓ�Ns^��|��g	���}�-p)��x��3sS�('�'��}�U{Q-�}>�F;.���"�� ��}b�u�sUC����Ff�\�Z�@��	��iV���Z>����t�ЧŝL`��W\�����)�d:�	��4ts�(9���p�c���1C���}�5���V:�jt)�+h��p�S�<���Sױ?$�'�X��C��ڵyyX�%�0���h/����SH�7A^ֳ�;��D]zr>/<�XxV0��(p�;�
��AX^�������q�S5��׳<�+<�b\��5ဈ3u[�v���<��قf T81ѳ.�n�r7L�"$e�<�r�w;�Ha�z7���z4C��U�/m0���Q�n���f�I�CEz��Ϙ�5'���!O�&0C��j��0���˹�?X/6�S�:S6F{+A��v���tf.=Cnջ���;��I���뛠H����O� ��\�٦AC8a�M|��h�1`��Q��C˦mţM���{'{�M�턤\|]DR�\r�����a`U� k�P6(r�t�qwrn�R�p?S547���2�*�ܿzz������u͇�g��H��Pɔ�X�yC��Y�`��y/���=\m�ݭ��j�F����*�J,ˋ�A�qQ�A�6�za�U�s���a%��Xd�6aA|uh��jj EPX�0[���fͨ�xZ[����G�� `�!��$���hu�^u}�}��o-�܄� �O���k%Fޜ�X�tP�؁;<��D��=J���D���~�Nu8�ޥ�î��>@��C�D/�A���پ����cՐ*��L x<�p��F��'�pbq�fTD��1�\��A)�}Fň
:���c,�0v�[�<��=w�_�>�G1��h�=���}L:�9�=����l<O�c�I!�:7�*�S�u\�w�v��R�S)P��sP�KOR,�!+�hd���Jh�;�ܑ)}�xx[��ɱ�>��*fC��F�G\��B�Ϊ�<lp�	VX)\������ *�MudD��m�a��K�0���^�U)&���%�����I�<�W.C�)l���v�\
5��G[�F�l�co%�2l���1Рш�@Q�ED/��.�H�L�&yK&^����d�|�f�3�j�r�Qn�lpދB-Ɵg�<͙��:��z�����U�b�ڨ�J��I�ì��B��{�r�-mѰ̍�v2�EJ���+i�����F$f�.l�Ѭ̓���gIy�3�-ˍI^ǅ�T��ɡL`���u���<�k��#���m{���ъؿ@��#�]�f�;5��5DN]Z\�������q���[Ǽk��
���W��(7�qK���y��ζ��sw�y���B��L�U���=�������Iޔ�r�Vŋ*8�4�q۵&���q�Е{��$�B�l���f�ظ�� 2�-�Dg���ړv�(#8P7����\t5tN�Gm�"�E����dnF�m�uh8�!_�֕���} �������-�R�0ƺ��eA�$��3A\�yV��ژ0�x,T�.d�u��9���:&�9��  jr�-.$D-��ر
u`�8���l<h��b��� �fj�A�}T��M�{Nd٥J�wq���%:�9
4D�]G�:�?�@L�t���h�>v�xc��r5��jER���t���@�D��C��&�! �L�6�>r���c�����O�;��nN9���EBhk�QbpJ�&��A�I���(n��P��	x�����\X�:�b��R�"|2:��xd��'�=�>xo���S��>U�X�O�Ń�yU����$�N��1��q5�t��X�]�5pa�ڹ����&R��9"R���t�U* ;&Lb��Z�;ٵ��b���� �nQ�x�A6;H�����6�p����sp��~ܭ�q�ϧРd��1^���{.:#6J��i��bڠ�.��)m���ٚ2w���!@q1���rxa�����|�O�]~B[s%��Ng���:!4�KpI����uz�R� �p��֣T��׳�ـ�Ҍ�O����t>���@�y����7��!w�`\g5W�g1���mcy����oG�Uᡓ�?����^�=k�}m����L��U+��R�����a֟��:���yA�|)�������@��������J�#��0vt�=��UwzB!
�x	b`bŎ�)%�hD=^���+��>��#Ä)���6�9�/r�X�/OxS��ԐT�#��_*��YD�~(s�PrJ���>��NW�T�Mڢ�{(c�cXܔ\2_vؤ��(X��v	�#eA�7�D�����Ѳ�,/{�Ǖw+��1*�ɾ���0����L�����L�̠�^)����x+{u�y�c ^�k��#�bzns����)#tH?s����8W\X�蠫�(M�aa���`��LP�����_K
*��*Q�m�\�3�����a�c���n�q��@��:*�+�w��νb7Д4�˫��X���T,=!�����㮶T�������q"�`�"U�&� �ʞ���B�RV��f؎Ίf�"��Y؆b��ƶ�b�¦o4>�W)T)������5�Fǯco/vޔo]-�|kH��=-��z����V�cJf$$��%lrA5;���;�f��,�*�;�̰��9��*�[�W��@�qk�2u�1����#�p�
��<�6�]ZV$�c���!�O��.1���.2�]�������]I-�e�(e9��j��YZ��8uX�g		$)n'ܤ�Te���|�J����8H�3٨.]#��>�DLdKBZ!���kG�b7~�4�Fyӫ��]�{ X�]�!�U�J�Y�@�9�N��)�������h�0���4�v5K�����ƯEs��ln�݀�޺�5�z����z(�r.�
�¹RQvl_W*G�qMbe���{Ǎ%��|+L-^-Y�Ι��Ţޭ�"{R�HQ�b�?��C�F�}~�'�H�u\7<��9rǢPɘ9L�C1�iS���uV�)�E,���˛3�x�ǵ}���_N����K	�yj$�)Y���Gu۾��n�qФRi���ylm�6��E�W.&N�\��?<�\��i�Ѵ�G.�����z��׮;X�P]]cccw7P�k��p�騦_E��$��e�2��-��W:V��С�]���]sW�h�ڨ��UC��L�2йG+ջ�e;��ݬ@��pnL�c���:�$�v��5)+Z��T��Y+��=�:]L{�Ȑ�e�u��#$��*Nr����x<�6�Vص���/�d�t��C� qu����"ԕ�-hK-%OXV
DF3V*�	h(�EPP�0�£,X��ʐX�B�%H����m��%J2�*TL�a��EPm�Xa&)H��aZ�&���`���aZ�XAH�
(#Am*0U++��,b�E�aD�B�D͕,�`a!Y&�PP�G4�Pc0�$X
�R��m�*!X��XTXVT�QL�,�EE ��d�0�Ra������*,XVW-#�
�,(�p�X��gL�RaU�.)�k
�&	*V6�����l�����<ˎ�H������g7���@(g(v��/�%Ҡ)������O�_Va�\��N�P~xM�t���8x����Ƙ
C�B��v���\����B�F�3f"���	���.�?ˈ����{�k�u�Q��kJ���a�9�7b��J�Q���ٮH�@�m0�����̈́����/�V@��DE�*t+BW:i�7�q��x!V���\�	��ޞ4X�W+�UX�"5d�ޙ��*��
>�F�glh�d�=u�u�����X���u�P9
�僃�{��}4$j3��/D�K9f܉�8Q'�gz�j��Y�ˏ]C�����X�V=���'~\8�Y��;>���q�Ӷ%�r��*B�ݖ;�TJ�	b𠎭�j0�kD�u��Vn�maI�����^�&A�*p��H��H�Ԑ�����De�|{�AXn�)����;U�/h0��Y���][��V�6鍩������!�O�����h>t$Ln������C�#%�L�ԪrH�7�U���⛑ܠgʌ��P_9��~ә�����	3�opm�w��ocE(jD)W,I�S��Q޹p��V��SE������Q��^��V�v)Ni��𽲸R�\4j3)�AW�p��������r�-���"��Q�n,\l�nɅζ�uz8�}擡������}�2�_P��D3]uJ:�l�;CF�9���C��c�z�����  ���cc$��;dã��Q�g�ށB��I/�����I��j�H�p�ؗf!PsB�y\�	Y&��n�-;��3�Y�iȐa��͈0"|���c�I� T��� ˭�8گ������[���+9�C��_��xQ���	��+�{wJ�w���܅�tMg��
Ҭィ�P/%MуI_h��[�5|њ�Ż�gv;`TfP�u}j����vi�hC�Hx�WM�Q���V?��;����u-�8��%�b�Ml�&e�II�;�O�(�[If��J��<�JK�������LA1����7D	����+�����w�
OI�$/��V1�bp�/�zo�U�Ql����Yz�|�N�VuO�mݴӰ��X4��p��=��}j�� �U���V��6�G�׽=�LA�Q��J�
/�Q�R��rJrgB�a~�7��ӷ�Q`�L�pt,{jX�N-HޛJ�����Ya∔���O*$�����3�8�4x�Hz�����L���Տ٧��r��{͐�y���h�]v�Zd��+�I�g�
P�����X]Rb�a�@��Y� 8�Ip�@rkF
����e1��R�:JP$]���EԸM=�����uIp���Ê��t�c���@�V�X�x`"����0v�P	(��}�ٌ+��Q%zb�����OAP����j�t"�d60���rc�Q�[|e�����{k��Z�V)]I�5��o��e�3�W	�C�hvfWY�B'W#������r�\ۊ�+X?>�?ʉU�"	C�֐'�]@T�{�ۼ��wb�"��CG70��4�*+<��8Mx$7/m��70Õ!b���������Τ6�eY�^�W� k�!��o��M�w���*���$rۨ�ML7F��G�y�S�ì88KŃ��^��Ti<�ˋ^B���@�%K�R�&h^Z�| �
���	�4)v�w�t�����h�S���U{C�>�����2w��*�
��m����̸��W�E�ִs�P@�yU��\%�����	E��*^�ip�Ɉ)DO�w��=�S}j0N/]{;�WQh�͛���8��0@ϗ#S�W�A�plo�嵴���;�����TUNލ� �0hd����*�K�r/h> ��]m�T٥ہ�ku(��J~�y���#9� ���,ξ#�J����K7�#*Cd|�ѐ8�R�2"	�����zo�p ����e�[ժ�k3�A���2^�xݢ�~W�So�e?Y�����b�����U1��v8L�@����+�p2?^����1�;�eK�����W;��v]m�@;�`W�LD��Օ��zA.�{gz~y�X[�_�/�n��Z|<+AH��.<)NDd��iz��z*Yl�MS�h��8��³(%��jIV��P���ޕ�@���h�Z5k���/O8)Q�b�c�nM*����D�EN��4�Hg��(<���ٿ�I9�S�3�=�y�L1��"��J�܉g���_;5����z<��Ì�y���u�&\
�Ń.t+|��4���/�����N�xثfP#5�?*���F����ϯoK����ٝw��'�E��P(]WG���5TZ�a�(��_=�j��~�K�����v��kM\��Ь��L,Z�Hk�Wg�ͪ�9�b�;��oELze@-b�O���2i珲��#}v-�+{�k�G�C�{p��!�g�V#�wn�"�< 5��N�O���!ƀ~��b�w��.���Q[�`�<��W
������nQW���q�����,�^\8�,A���d�2qU.f���4����u�U	�,�&�#��]����%�Vk-6��W�Xp�i� ��Ë��F�L�,��C@�i'� ¯�$�:%�OA~��P_�9�d��Ә�Ѣgas�+%&[�H�{}r,I���]y��隸k>�Ї�6��2_,��X�n&��90�c�Ŏ蠯:�NL���9.�
��-kö{�
��mӂ���P1\5|�1�a����T8F5��8�^�e���R�J�4���D�
X�f�EMx��]����U��I��LEP��(1��p�D��ɇ����vxj:�u��ԩئ�0�L�H��ol�E�hD�����wz���=\þ���������:mʹ�Q��,��'Ff��"qU�A�a��>Y�Wy|��;�,0QG���J���ԗ������TmL���#%��J��+�!�C!������A�(�{�]r��1\-�C��/Ư�@!�4D��nz�0��w�ֺH(�#�=~z����p���U~5�W� ��p��)Q�pE����lq1P�ʘv�3j�F��0<J��pTv�䩈4�x�nG1l��@^!�ۖ�] '�����1N�m(9�],l�[��BmgH����*q�[��7\|1�u�V
-�b����Y륪PT��&���LK�LWJ
ec[C������y�� LL�伅�H�T	����u�sh°�l(�U�T�Ӏa9
��/�܍v���0�"fC��ٕp�P��:qaHޛJ���"1,�W���aoΦ�]+��C�`�h{�Cץd��鴧{{_�
��C�7��μ� �GǪf�ە�
��:��}{TX���d-6yԖ��f�-V�t��`]�9ɞW�=�*��H3ӴY�Bw+][���y&Δ�	��Ь7s8��A� �����̎ͬ& &0�y]۝��~�A��rc.j��w0��D�%��e]�
��Q@d��.)�F���]j�i�#n�lI���v���p1u���i(����,y^�R͋�t%��c�;�+)R�x��Ee��r�6^Y=n�lem8ѳ�R$�� R� K�B,���~Z�e4�݈���b�nmeˇy��'߱Ј�U	�N<�!�	��a�|� `�ވ�)�Ȁ��>�c4VyԆȧH+��k�©�q��~=���ZlpP�>�W�cAԈ�f��TyW�b�<L?���.3:!v�޹�I�B�q���@IˌSބ�ܭ�pc�!@��_Ϻ<$zG$�����񍹜M�)]�Ò�s���~�2��>�$��yT�&EUk91��9G� ���_�ęn�S���f��bP�2�����f���j�.��mo,Ii����!������51>�G""2GӰ{�i3us�������{��~�/u��ʵC��F�{����+Z9֨ s�X���J�þ&�¤�Ō֓ҧc��Z�O� C4�\7����r�x��� Z���N��`t��bMLWK�*�:�jP�r��&q��T��9޼�t�R�Ϧ�����ވH��C��} ����o�Ҏ��dO�ʩe?b���.�ʯ�"�O���Ѝ��U���T�%�UD)Q�iC�ޟUs��kzj\T^���B�w�wg��O�b�x_7y}{ep_i��t4 D�JP.��jY5ع�#":e;����R��9���±��~(p�;�?<s����U�w <;�hd�����b��;eK�6D9�#fT_H�W*�iƛv:	�5���ȏi��0\���w�N��� ���zU��������s�i]�o%d-v#oz̤PʵXc��k��z
�v�֝캕�Z��b�y��;P"�y��sS|	��fɉ�1)�����d�X��Р1���^ۿ\�Y�q�Sm�~C���DEx���_d'�mT@@���ٮH�Ag�)��\]
̍����:�
鈳.)'b�+��D^�)�6-:�;Y�dyL���?,���i��	� c}���<*���ﲕ�܊M��\ *_��
M.U���Z�a���r.w��b{i��,mԉ@��agM���Q�.�]~�v�ρd҂Acjro\_���R!����Ů� ^�a�Nu����d��ᬗ�i�ɧ����9��=9��a�ؕ@��գ��F .KՆ���ۼ��PP���Y}��0��YE����H�#�CN�����E@���	R��*��P_\����cM��m^��[ϓ��Hyj�t�0��C�ǎ�(�r�ۮ��>P;��X|t_�ێ���qgǨm��5Q�]������6٣4nY��o,D�	.[4�7G[����%J�XH�M۱}��X�$���^�F����T*�+)�'�W��:��6���R��9.4필V\����|�;4����.*]<s*V���IJ�ZԨ0���E����U�U�Q���-u��Y7���t]���hڣ���g$�+;rmr�!��v�9�7��G�FhXرh4pnU�m��7.6�H�5�vӕg&�	�=O��v��aչ-(W±>K4�ő�3aOV e�i>ك->�`뭕�u-�u3�y��E�O�2 ����A��lY�����y������1a�]\¶��<R4��z3�6�{!Xt]�ɘ�T����Q�k"9;U�F|�{�K&=�����F�r� #�7K\���R�+;@����ʴ��n�v���U�4�&h�����YA�KQܺ9���`Q����j�<�O�o�#x褷;
�c�!B-I���M���k\˵Gb[�]�Ғ�U�j-�v��<��ԍ�!U�v(y�*q]���$��5y�[Rkܹr*Բk�O��F2�'^io�`9�fJx3�k��1�p��G�=��8xs�A�m5�vm㼜j�9I�n,�6�;ǶXD+D�D'��>�C��/t�^o��`u���֣} u3Q&�PP��2���(��yI���-��ST�n�m�f�!Mi�[P|Y¦�����ї��Zn�����=�~�|/6��l��x�޵ R���|�m�Y�/o����@�ۀm㣵R��N�ڮQ�+bcme;�kRA�X6I��܆�$�˖��6��;'K��R�BJ�
5]�͂�J��8�<1q��+,>�+Q�+eՒ�,�]��Q�o;8��;b��9�R�[�����.�`˙�-.���uXv�E۴֙I%�m�"ouN�&��L�g]�]�c�����_,3Z�mu��jY�'0-x���|ϳ��"�g-&������VT�H�$�Jز��S�aX����QH(E�
���IY
�R(
��L2�VT�()&P�D��	��`�ȥAH����D`����0�1d�
�Z���Z�%J�(�m"�@�RV6X�dY
ʢ�Ȳ*��EZb��SJ�(�
�XE$UQFI* ��%q�1�nN`�ڶ�b�.�n͸CL����5b�N���n{]t�'m��V��`L�6[Lm���q������
��T�^ä�^�\)V��N�+^:�w�fya�ɇ	Ȣ�b+Ɣ (��X�s��{&:ڑ�X�R�J��^�0�f�٠�ː���s1Хрs�e�P�}������=�bN�!��=��5�
�`U�V���[CY0������T�rr6�n�51.D^R�D��1
���K��B�ȜMg{C%.�I!����t�mԾctT����|�W��?��H��{/�{��.o6/"�51��d��5��J	��yC��˷�[�/.���-�ī�0��B՘p!��Ds���tMg�����M��å�B�w�����d��ŴbǏ���mV�b�_ب���]yh�S��ޭʐ�f>%ؓ	D�R�����=Vh���|�XO{�o��&oo�Z~Z��y��d�V����z6���ܬ��~l�Η`Eˎ�]���{�X��֝�|���m'ۈ�$6�.!��ⰦLA΅V��r_zu��)�;�>]N"�2IyA9Zk {`��#��&"�֔.)�6D���������pvL2�l(���ꧦ��4%9)�<�	[Qr����P�����CT6z�0ʆ�mB�r㔍鰕��9O'N�D�29]ʦ#�|#����E�@�}g��P^����>)ͫ�Kb��tZ��ڹF��*�[怭v��~�L���c���	��.��qQ1���y0�"#<Q��L�b5wԩ)�D��:����c U���s�Z�4`�=��������]6���*+u#�-���6p�P`��D(;=z��(X����zi�[g����mׅ�^���W�
_ �%Et��^s����-!�
��`��E��_�6�)(�)�*��4?g��y�^�|���x:wA/����c�o��wm#�wC|�bM����<8(q����_�t�]��`Q�o�S�Z���u��IҭUi�mgYT@q��q8w�o	�&u!�9����{�� qG�j#�
c�4�c55��3�"��`&6�C��)m�h}�X\ 1P���tj��G�{
���Z1x?�:��ɽƞ�T2���E�s�uHL�˜�q��
H=b��w�TcAzbуGmD���Z*�Q[J�Z:1��E�v�I.t���ׅ�k� �J��1�=|�Cח7����xu$;��bF0m�@��
�*w�2B�mڌS��̺���y�9}���T�F	꘮�,J����Pr��f���|�f'9�'�u��Y]2����k*�;Wq�T���5�V���-�"ԍ�v��+7�t������t(b���s=3�R'�+�3[��P:�t�d\�1ٴǝ���*���gEL��)m6�!�öD�]n��Z@A�&�V�U4��i���쾬�/;j����a�	�gR�l�.��fcN�-wN������`�^lﲸ� ��Nt������� wڷ�vd���4�LgJ��_^��}��´t����'�WqG'����*�H��MF^Vo��ez�ʁ�d�9�NXw{v���k��̋���+ o4�^[˭�\|�a���M��@<�����v�b��ڿPSH�@SA�Ps���voƋ�F~�)9	L�r"v��"0t��UB�L�=q ��\/M��ng\�<i!!�ʸ���aӉ�p0;�"̸�$�RU9#H��1�g�"ȝ��J���$:���U�� �UnW��}�ݘ�{��R˧�rd�y�������W0,ڃnwt�6��I��Z>qI@Z�)�WԹ����d��,�{�� ����J�sk/UOK��p��3����� _���;ǂ���Y����]�°���Nbf��s/[��U��_l�/.�V.����&�55kj�'zE�]w��iHBoS"dw��^�<�z�Q���n�r��u��@1; ��,��K��^�^�+�z��km��z/f��>�z|2�T�U KXPTuh���q�ډ��ޅQ����0�� �P�0��[� �p�"#"!�V��f��J���
������p/�҅yJ���}]t�3����}��f�U�y�MИD�W^�ML)0�\y|��}Z=~�W�٩�l�uz9*�٘/�o"�5
5��L���6O��<+4҈���X�ec6��Ш����R(NDxTpͧ��S8q:�o�s�_A=ǋ��?E�GD��A��!'Q�c�x��h���vI};�{Ι)W��8<3(%^ TZ`^J�����[Ep+���y��+H덙��ט����D>\��T w�����x'��7\��\����{��V���l�
`#j�R��@�K️aSʓ�^���:�q��_��إ[�:¤
ᎵWW�8�Z6�V1c��v��p���WWGs`��nQt��4塻7�����qF�3���e���TQ9��G����_j-�"c��F�@�&	���Vy���߭U���[1�ɛ{=��Tu��E�d�B�&��DO/��V\K��c�߷��ܧ�6 ��q�`�>�|�V١���h�/��
4���ΐV�0��q����{8�Ɩ�c��b����]%�l��l�c��U�@2z�@���89Zk= ���y�bn��֮�o��<ySiAO��:'���br΂��a�r�<�Q
7�C����T:�"��kiB�r���9qf�/{���s�p����L��ut�.����4<A�=j�y���^�l�>�g��X��*Uz�b!V� d(!]]����T��:>��'�����yW����  g-���B�P|z�3`X ��(/��{/n]{k}��Li�v5�O!��mQLe4�n��gn��KfftHp4��\[.�z*����<�rV��Y<�^q��D��;W�Jp$Do�҇Az���]u�Y�H�H�K����[g��:��7�^̝�E^���������C����D(]&��Vži�%үWQ�Z3O;�낷����D�>�-�:�g G/!��S�~�fY�@
��m�+,�gG�]�ӳ~.��	Ƥh�
�z�W-���`@q�b��<*�B���)�+<�\X�Hsq�t�f��.�
�>Ub��yF�*�HH�T��ʼ�A|P����e��=�4��c`�=���_J���9�!3C�)��\>T]�ijA�+��6-_�ы��6����:�++����kGD݂�Z#u�sE�3A��B(HP+]+4C�� �Z����Y-�܃���{�wRѲ>��W��ʕ sHv�����'���o-v|�Aý4p�Ub3e�֬)Y��q{ڵL��A���ֽ\�&���\�%����AU�P�9cJE8LY�)�Cɯ�k�����թwf�7r+AN��/��q۱YQ��c�f�J4OT��!J��@ܡ 8�/ɥN�(�m؛R��2�a��U|k3��  ���S�Y��=ǵ�E@e��Vn�O���B���c���Dl^���+����֭y�����cǯX���|7ƣ�/�Q\tl9��&���_ �>�F���*�W����J���>_#-��^f���aK�@��6:�]��z�u;:�۲�m�Q��{M�a����\Fz�xx��gy��AX �y�f�[���R�`C�����e��Ƌ�ê0�{Ƽ(7����0�1�;���||�����B�Ùh��Y���T�Bx��@@�/��b/L�Y����{}��C���L:�c��r��
鈳.)'b�%s��F���c��U�Ih�U�Y�x��-G�pz��N�����ˆt.�J[83&�ә��ꕌA�m�v�u��B�v���4�|[���a��cvv�nOϩ�u�Ox������P�G��
�X��1�b8�b����тe:�KQmN��ץׯ�g +=��"x|�e��jA��/�u�i8���F���߮H]�X��Nxѥ��~<?d1��]��w��U�]��^�/�-v2�5a�6�QVi������Ĭ�-�jD��=P��i��p��U	� �X�@Ӄ����a/۞�>0��*�bA���z��4�рJ�/�1ז�v�f���B�˓Cn��ę�J\�0nv"���J�ݭxv����6P[�p��L�@�����t��0�u8�x�Z��ˇt�gI���Q��X�ϥ��{E���k�qX��o��=|�d����wK���3�=��T%*6
�@NDxT��!�֧�+�|�Ͳ窭 ]X���']�@�c.�[��[�z̒6'T̾px�83���=�����[����,��՚.gE6�����e�`UqsRE�v�Iy]�J�xn�䜎�ET�ߡӋ5�Nz�
I�E�S.]`U(��-�WXNe����E�ʞ�a�J� T �%Z��:�;gu���1�y�{���=�X)S.υЮ�Ȃ���f[�W-Ss�(�����IJz�ᦧ��vH�ym�Rf�_x�X�Cb��L@7��]L����XȀ�4&+�F��:c:�	�^��V�Q�j�sb�O���}۳�*���68{N&Z#�B�Y�	O�'��_���\ڑaA�"6%,��9q��6e�X6�X�+\wԽ��M��K�l�vf��.}�^JR�l��Req"�]`�狀U��\tW�WgEgEQ֩ثî(*c�~ϑXC�|�����Z/�M����^�+Ɲ��:�Zr��ie ����ty�1�1e��1ru��LWFw�'6�)o[Mޭ0A��Z^�6�^n�c^Q/�d��ۺg&Muڃ�4#Y��Sq:�%b���Ab`�F�����}\(�9-��.���/L�(I���u�i�1A�3���kn��]9
ZR����\-c��c5�dn �V��kb�h\���+*���bs#��fo9�w]��y�Qñ�˚F�W�檐U�|�RM�*��_j��j���V��ƍ<�\����yv�ڮ�&���X& ^8��N�x\�r��]ir^���_wc؅���AJ�DOC[���N^�Zgw!�����
��Jﴳ�h)���ޓS�k�t�_\e����W%Y|:��o+g"�Y���g:�R�ۡ���RR7�c|����c��Ћ�{���wm�P�|��.���2����	Ae�s�O�֖Ҷ�,���d�������+O�N��m�"�;�P���T�ct���[8��%y`t�yd-E��oSё\�c�dL��<���{k.U�9tܫ.X�G�{�
p�[P��K,���GD��N�)t�Ykd��J��/�����d�Iօ^;Jfe�E�0����N��x�x����*W4\{yZӠP���j�꼽�1U� m�Ć��͘��c)����-��
vH���:]E��M�R��c�t�h0u�]�j[i���	+���:'��F�Y�a���"2t���-��$*d�{k.�C�Պ���.�$[��� �����BZp`�4jɽ4r�Ǩ�"�Z����Y˂� �*a��q}#͸�.��粑f���o^O�n���f��O&��[���-�K�<d�Vɓ�8��[㈋�n���Ո��g�P�Wj�[�z��V�����Z��A�c�~��$�w8P�i,�Zj�<Rl���,�u��r觕���=Fr���hD�����d�����M��t�ޒ�2kL9{��31��t��-o��Ҡw6��r��n�}���4���DDAb�Q`(e�DI�P�aH�����XؤEI&(��V,QEVE˄S"�dU��Ŋ)%�k*I�RL1B�+PQE�,R(E�
�*,��+j ��0�Ha ���*,Z�a���#E$PD"2#���X)"µ�B�m,�I2�S	m�φ~5�/�o7�7O�Dlcq4����u�p�q�"�ݕ�y�<���	D����U_VOr0�0dr��?^�p**�m��p��jX��EڷwUz���A�ܐ]b�C�[��y>�Z9�"���7FOK�;wr]Ӽ�VP��l�G���<T�[!�D*��F
^��H�{C���$�|DȾ����Y���X��*��������-ջd���n����Λ<i��i��j��w�_\ZW�S5~!t�H�0 �#��@�Р����ʐ����q��]b���r�W�xf�*�T+F���*f�s���S9lX������wMׂ�����TJ��Hb���Ӳ��Ƹ�~��ȩ�~��q@��1�*ݭgD��L?��&ủM��i�bM�G�!�Q
)*�0�\# f�<%�B�g�D�S�v�u������z��J�*U�@x. X��sAȈW ^MJ����q��5���<w��&����W-�SjU�A�+r�(i׽����{��^X��r�ZԪ�̵˷V �Ь���۫�.�4��[�k2�c��f2�������,�ہ7W���n�WR(�NqΩ�!3B�+j\BW�Aܽ�-`�0�B��L��/$$9X�E/j���P���fŧ�G)'F�9����V��
4�φ���`�q�5�G�!9b��J�ʍ�*�{���%5N�����P�QQ�1�AF���N��x�0�.��Z*r��tu��< x{j��r�u�NE�(=�m"����鱋��g*�|�u�HB `���H��}��FL���+h՛��|꥿�y���u��i(J��u�P�n.�p��p����~K|뭬g`����L��"&"GJٹ9˙Q�gS��:�vM(�����EB5ʯV�yJ��p��d�4 ����炧�p�p��]<�5����)u���B^O�X{Kx��e�*����L&��+)tբ���`pV!¢4ҾY�[�jW+��*˸�eZފ��4EJЗm����*7���,̹*lv���~ =����ہ���5�8T*�v0*
��Jf�}o.��q�����y��ND2�t6e�0�ڠ�D@��2;H�4cJ��{���=Ӎ$�Ն�j�$�PڵP.0 �H��|XF����{�����nOyPϊ�p�u��vls�PZ�R�^���Ϥ��ɬ�m�Ǳ��0p�W�Z+c­aC]Z��ʬ-��@'��mҩ����oy0�9�g}����S� c�P�� c��L�F��mS��z��
�Ba�����{����.��sHlˁޮ�b�r�.d�Vz�Gp��	ǉ���}�p����~�o�3a 0.�85�Yy���l!%�G)���7��!��J%P?��l`#|6�+��YZ'�sC�TDb4X�0S� �P�/]t>T��B�{��w��n�ŪeY�핸�t1��� %��9MK����w-U���l?3O�ҳ��`j��(��%�L|wp�N�->��C�s0$㡳'�����=h���J_�	��'Cb6"L!Pn��$>�I�sۗ�w��+��9M�T�eq)$)G4�=p�tT��	9<W�t&;���+e�N1C��̶ڰfT��	�E���S �T	
(.�����q�Һ���e؍��`�w�R��(N58�.��P}�W��)��m��{�uh�����j^&��Nn�
I�E��`�90+��r0F�z���-]+~�k�1�yd� *o��cc��M�F坽8}�	��<�³�(W�|�**�p��*D'ۨ��z��,F�ҹr�O��yt�
b���Ų�p��_*��yq+ie�IX���� i�0Ɍ���h�&q_b�>�V��j�09��������Z 4`�lA�� ��Dt!���~�īC��́�͘��}|��e_H-��z��*�B�ˤY�����V_
�z�7B���0�P�͵/�U�,��[FRw��vjY�N�n! ��D�S�ӱcI�u:��-���ﾛO�4�n�?Cb�P�q�eBS��p�# d��: �ī��*��-� �V��k�ō�
���%�@�/g����x\�үC�OE��ً�
T;�0,gQ����zJ��5�=�w�ܫ����v���bĉt9g��3HK|��r���~2��l^�%��"�^����֏
�¸$�c��
�P�V�TAO�:��t�����tXk,'3�\#�D@�u�S�f��Y�	>y��4��_���W*�d5����"4A|h�Z���F���M�.-@�:WQo*aBg��.\TL`.���LZ����M�!-B��d��룬o��l�4p��kC����E�сrh2���2fZis`��݁X=�p�>)�S����@�K��$��"=�,j�б����m|��ͫ�3a��Y��h�NYV��v�|i���U�1��|�Д�-�V94���%A;+*i
J}�y�7m?�M�f19��3���t�MX����Oh�D�>v�x*����:õ��I��&��i�D�bLt����GP4�k)�/�tK~t��U�>�5}���P���QpGLA��i�u�9�ګ����^:��	&O
��U�N͊��^yR�/�W����	���.�����"xsJ/f�`(g+!ۡ�$@�U(��WPY�3�NQd��t����[�e����Ŵ����ZM�#N��L����������eo�{�X5�U�sK1PF�Q�p_�0kGl�
��q3&��&�d�.� t��+��P�q[,��^��
�G4���~s��`!Cy��\���a_@�J�GL�@ض�_��q��F8ie_����
�T��s�V٫Ru� B
���vśl�<Ux��jIb)�7��k�JsR������o�ZpkkWg�Y]���"������>w����A�c鄎T��V���b6���x؜݅�o �drIIowIm/R&����3���R��C���\�U^�������[Uȝ�`F��8�_3tb��<=����V�nE6���+1U4I(!/��
[F�a�,ѯ/��</O����0_�K��*��� �7��H�ؿ]^٨%ӀU�0mne4;�(����G�7�p7�T�>���گw���	���#k(rޔ�����i;K^�haY�J�*^#�?���lD`��=��� �ʩ�����JΨ����
T�P�L��
XF�'섉=��*�\�Ӎp ��*�i:���!���J;�"�eB3G"��Q���(�<���	Λ��drc�G`ˏ��n�]^$�['��@S�x+�ޗ��mW��Y�Z�Ҥ)��kN�5�}�Օ5�"p�ҙ�`Uٮ�h��[)��Q/�����E^iK*�ެ-n��M.a�}�;C��Փ�3��-�� ;�{(V;����"hΣ�ّęn'>�{~�qޱ�cmߧ���0,���3�El��������i��w/j�9*_J��
|�6Df�d\DV��$Uf�-�ۆ��^K�"�\��ˬ�x^�w*��2b 5�zfjha��uѵ#*z"(�����������hA�Ꮢ��*m����0��Tt�R���|)قmZ���]c��֥�m��:��b����AZ��Rܘn���!_�U\1��!-�I�5/.\`�xU^���ҵ�Ӌ]@�S�嗲ˢ����99������mR
��
�j ֨+C��ÛUw؛p&03)��:�`wC�Ƨ��Rr'" �t28���r{�X�l?���8�/~	T T�a��/>qӐ)�u��sK�����t냠�r\v�ɫ���X�3�m��3BK��D\�d����js;VA����E�^m�J%�T΀�%�RĒ޳h�@��ro�kGZ_E3�$�g�Q�7����A��׼������`Qɘ��>n
c��x�8P8�"�ϋY�����uꇀZ���D=�2��*��ZڿMk�&)�\�+W����F�b2+x���xHk��j���h�u�L����1 ���S·7GE(nE����	Imp�nHɗ~���瑢#��]�,��Z�xnY�m1B�Q���+$l��	u�:��*|S<��Y�/�<�aд�[V`	���V�K(pr���e����{���Ǿ�r�ظ�	5��³�竄�U��*��yn6j��x$�3�uֹ�rd�P����q06��1ʆ�d��X��%�܅��+)��6�ʄKV��wj�YV(� Q<�w�lWT�[nS�����vE�5P�(�����'3�þ��X�������EB��Z�R�(��/9��n0K��BSp6����yWN)��!���Q�)��$�����x2
�����b��j��<�R��9j�u>;kޛ���O�
��� ��:�g������9��j��7)�j�.�}��D ����m`�ά�H����ꑢ���B�P�uj,��N�`������]��N\�ɯY�ٮ�+��3~��tH�yxy�^u*�0����n�-b�0����S�q�{�d���=�t*���$ gP4^�dSc��KʌO|X�ٖ:N��Tv}S ��5W���� ��*��!Ё�	x��<��'p�^�Un�[4�إ�R�*^/�W�����h��ƛ�
�r�e��{W��VC��e� *4)�1�TZkO2�&��k���(|����/ؼ�R� ����m����(�����`�ڬ��E��-�i�A{�b������=C,��H���:�-�u�,}f������J��\�n�P�į�b��YH�<ɹMe �f'��ɦ���@�] ����V��4�ۼn��1:D�Cw���֓��p�47f��Ds;I:�h��PB�^��%⼢���$�g�i���Au��'4&=7����)�z�ïM�g�?qv��Բ��l�tgTʂ����a0s� ���;8�6F@Rcn���x��u3���[�n�eV��^�ڕ�ׂ�q��ڤ�"y�Vm!��Z:ԡWԐP`�R_< $K�u~Զ��z�cr��޼W����@�ʕh̘��`R"�.Y[�B�XV����ړ��q���J�臒��LL�[��2܍�N-ٗ]/�U�B��5��6u�Э]W' )���v�Ӕ�>��d)��O���.#��h�y?�Vʀ�Z\��S)3l�G�"����v�=G�!m�Kg�_��V�
AȇPL³^R�3b�j��:%rq��̬�$^7K��r��S�`cˮ�q�˘�e��<|1Ͳi�u���n�Ĕ�2mr�{ur�U��^���} ̛j"�fñ+2����㽓�ծ�`�K���$n���7V���.�ʳ��Tq]9wzq�&���%-5"T�`�8��@�:�^m����5��[pR,IpϮ8w�4������Xy>65nC�w���f�-�0��c��#�,cdI��=�}P4�ȩm�C'�����65^^=�V-�Ja&�T`W$�7c��a{|I$u�3��[�nӛ5�5F��GV�+7�#����bS�Ș��\�h��M�㹪��b��h�	�n�4�T<��FV�f�Jݛ{ew\h\�F�H�k�Zޡ��)�bʷLk�!n��	���xтM��"�u�u�(�ڷp �"
�[b3��23������M������%�r�����E|G�D}@�Œ,*	m*B����x�I�����C"a0Ԋ�`���b��a��()XJ��kLل	3l�E0��BV�+*VIF �P�����%Q���H9��(J��V,�m�7!X�U`T�+!X#"���*�`e�B�%@�>���B|�����UL^l��u��n|��[ySn#�kV�P������I&Wize�����k�FS�9���#To�U� ����Cv{�Z+��^&̡q�.���/e�̍�Lל9ʯ��J����YDz*����jr�x~y�EC�D:��Z,�}Dj��>2��`�S;��e'�Lu�Y\+���G�6P�P�#Q�ͦD�lDf����7��<dV�7���P\�k�"�/E��i-E��������(`�0m3�Ltz���A5��}u=���e�a%-Ht;��(Tǐ	|�����c�i�o>���A�_#[Ǉ��)�Ѓ�TzoP�n�f�;V����.��tzߠ��f���v0*
����j٬���|Ӝy=�6���9LU�?
_2jǲ*���E��
Cib��x��k�FcAT�ڇ���ՎJ��M���9�f�_M:�L����Ab����W���� �bw!k�@��p�+�,mr]hGu�A�<*v���F����9��۽�hpbb۷Lh�S��j�/��!�5��u�V�{.fw��	G����j�
><����2��{rU�צ������RV(PG��^�oK��}R�+
�Վu��ง�;�&�f�5tX3���;�����Y�Z�Ҥ)��4=yyX}�˚J�ª���E�p.���wѯJ�0m��^��'�&oz�]p�����ӫ��7�{Ʃo���������5���u
�5�S�՝���C�uoZ�p��!U���f���>.�q6=ZPGmQF v�����^��8�U�z��GwU
-�Z�@��1��G�>�!�I7��C���#>+4��Ly��<��3������ `�����!�
�=~�FV���Y��ۚ�_���B�<�igЎw�e�0�)@7d�_h���Q$w����Aj��m��M{F���:jwR��:�<��/6u^�"��\�;T�bӭI:�W��W�hv�دt�
Y	���T�]��~v�RmK�ˌ�p:=cgT��0Ԩ�#1=FEԨW�k,�����(30�âg,F�P��u���K�)9����M͝.{�j0�.�h�x��჆Q5 �0zw�K�=$^Y7�:�w����NQ�-r��I|QL�pM���t$d�0L�W�}�:��71O�ldW��JYh�J
C��P�@Wx�Ev�������ǁ��a�!�4F�� �(�%�_e,�ϛ���;�w��1�i�b
�y�Ὣ�h�q�xZ^�~�����l�
_%X,V��W������`�
Vj��X�z=�\��e*c�Z���F����W���4�0p�im(��l!��خ���P=�3���h��>�����<�E�U��%
��-n�ź�pq{U�.�oGZ��(�v­�$r=L_%q(� lٴ���E$�*JI�_�`g*�d�C³�0�
U�U�{�V��Z�\�攍��!a��&'#��٨��-��)����q��j�~/<^���'b�l���H��\k��6���V`��
23f�4���X�1!G`��r��ο��8@�Z��t��U��y����|n�T�[!����v��y�ӱ�ȕ��`th
Dw�׺��^X��E�gVR|t���zG�H Oī�TM`�{��|* �U� aL=�sʋ��	�������U�'M��>�в�a����ZK�����&�p�A�U:{G O�U���x~A�}XϜ��F���x�W��-5$ @T�5�F�	 V}wг���a�E���AM��sz�Q$T�[v�eٽ[]Ai��̬c���\��<xQZ�t��r��aħ-w��(hq�w�Z2�V�����e�6c�o�*rri9�7$�Ç�qP
�h����i�U
C�7A��>m�=��^��\k��i�+�����q�W�������n�m'|f�+������J/f��Prn��D*��γ��^����~�S�X�����p0F�Y�RV��˾q7�gr���.	��<��R|��z��ug4�Tj���������m�R�+����3��P���9�BFʘ���OE��ے�\�r\&�s2���(*\=�^ھ�F��gQMh���Z���:/�{�Y��������s�qH$a*�e���}.�2q�w��Cb5ĸ1s!��鑰	�����S�AAr�����,�U�ԐX�ʙ�3�BD�5&4��b��<</�P��e�4�;nkx�.ê�����Y��u���K�:�}Xn��B�\����T�T���|�; !�c1�����A_}�P�Rsz�C	5Ttn#�
r:��F_��:�Ѭ��Ѩ�/��z�i���Ţ��>���R���cC$j*����
�M��J��~]5=�I�3�+SR�5�g�P�É��Pr��;���AX �|��W=����F��m�b�C��*X�(GqW@��d�-P���ޞ`T��Z9��ӳ�J�D�j�xp���"�Ip{��Fk�� �˕�
�DzmҨ���Pb��
���كr��秒�7Bt1Ƅ�K'd�ҫ�df�(k�c�ފm�}���}h�Ѭ1��o�`��!qY�PR&�B����ֲ��6I���Eƹ1�T��1m;��!�������=���S�Jͻ���M�W�����[�N����(���֥F�*ؼn�*���<���U��}�<L5��c۷����bH�2�`�V�ii`��U�r�#͂e2�)����Ⱥ�����h��๙�N�ѱ�wYM�ڹ�"�l��o��	�ƉCl�*+Vk�>��U��;�RnE'�����c.�ùC��!J�pW=�L�m�Q���78��\�< �ag�GI!���h~>��>���<<�s�w-t�^����NJ�]m����0����k�_�Si��K��j�����ϖ�*�DFUdD*�Z4#QF�6�V�nf�I7�kN���-�F������Z��<�ꡬ�d�ZS���1~�����EVb�������r:�T��v�mcř<	�OP9�e��r��=t'�ܹ��cوg�s1<�78�^S�1å���L��>:(�C�T�e�D��!��EMPX@�S�7x�U��-�[v1����P��Y�-]b[#P�5(s� �u�]z������*mK����(��Qh�&Q*G$'�����V���!��Hn|X�Av��U��y�t9/�KS�j{»�z����
Q�Qյ�!Q�������S�F�s|5⚺����#5%k4�Y��&˞���������ik��N*��#K5���)����=Z�_	�y䄽cD����{���ڑM9�fdF����\U��
r;f�����&�v�*��4���Aq��w7DM�M�1R����u)�[�]I���4�EM����j���l��k�ӠR=�-�c#/0�2�����tbP��R&���P^�Xi�������d��K�PǴ@ꂇ&�5�A'%`=�/k0������W_k�TszҚ1�j��y�
�L�%Yw��g;�����]��O��ܗ�e녤�9��d�m�}��ޱ*��S��L{Z�\�QZ^��TǇB4Tٽt��h�^G֏��u2��9quًKЄ03Jkg���9��Fo��9�n���}診>��Hq����Ye�T��e�ue�n]"���д'�[,���yE�>sO�����T�<n���Y�588<e�C�7օ͒����|�	�S&��U�ucxUsW�&��%��;4;�^�˲E��"��<u�Rhfl�+/I����k1&ͪɫ͎�8���sHۤq2� rߴ�U�KI٭$_\،AvgI��v��/R�#P��>�u���x0z�y��7@	��+���hågۋC�T���3!���!u����sN=�[%�V����U�e;�;;�C7W<2��k�j%�.eIu��<j������;�t�F�lZ��/�5���C�ا\
��M�s�®��'{�&<�ޕ���7��w��šk�I;ά�\�������Pލ�ف�vRwpy���S:�Z:��+k���|b�om�%��z�h��X����BğuA���J�T	�ޡ'\e�f�oc3V�N �9~Ξ=�q˜����.͟f�i��y��+�u�x����'�88˞չ�X�qo���æ;��-ш��PjR�hY���E{[��p�x�:n�B�W�T� �O<(��Np�C� ��,v�]��ܙb��S4@�,՚� 1Y%KE�)Q,-����_��kt^郕]����K$�o��J���qV�h�1]r�e�������x�.V����ae\��:io+#���{L���\Qɣ��rN�IԺ���0�Gȷΰb�f��]�DğP�@���)��H���T��d��l�*d���{sv��"⍌]��Kכ�&r�o]�9%�L=��)�e])�� ��8�:��s�YA�r�.�"�%��>�>%��kh�}WC�~�'3�Z{,����"��J�������0�d���E�
�uej���X�7n��,�ז������E��ࣷxR�� 6�d�+�3�Qjb�fsW72�u�)����%��)�=�|<�*�5���k����y�tٵ�>��1t�yƉ���J�2Ե- ���R�P����lu��oNY킈�\��mQ�넰�#"��iw�s֬*V�Ⱥ�p],R�P�Pܶ����Uf�^���r��
`��WsI+v�KY�]YwNZI9�ӣ�x똂�<zA��)sL٦�t8���1�*�[���Z�=��ő(WY�:��b���}V#iV|�l���K��{cq�6��|kr8;^�?;Pԝ�\0�^�Wf�>���;L�\1�����Z�!��[CQW!���F5�G�V_��ul[ʻ�Յ�u�6h�]^`Z���uD��0���q�u:�l4W�m��%l+X�L��i$d	\�a�9�[��P�j�3���`$b��LT:[���oJ!�Ay�5H�n\�p#ld�('u�|�`�A�,mHͶuc��lnǚ\56RK��G�`e���-}:��S�=W"��oH�XMŌ@>߷5�n��l���B���I�ԕ���7�R�$�D_d�Ӛ�����\�w����G&�ʣ����bM���}�&�%i.(�Z�Y���w�vK��)¾���8��� 7ɢ���r���[���c�E�XT��
�jV�`�E�P�ڠ-�bȥk���F�QDJ�`�
���+%eJ����J³6�p�9lCR�*EKJ��0ႆ��"[
�b�e�Qd0���6��qHaZ���Kj���B�J�ѡYP���L4`��)��&SŰF�����&tw7�l@Q�1M�Bj�r�ھ����[F�C��N�Y'ܡZ0i��Ew�w�R4�	1���P �gc�weꝈ���\�I�B@4���Zv�Q�#�s=6/�9��T%�um��b���s�N���W���ɿN����bE�
��Xē�ϓ�}������R�J�-X��b�H�5{�]�7�[y�&��f�S)�vΌر��S����T�7���e�nai�}��<�CM؁ kЌF쭦��V��j�]�д����7��=�-g�G�� ��R4��⡓�~�0���$�s{E�KЧ�C7�h�]��r��d�wQ�R��V�[��G|��We!2k{A�����zD�띵���K�6ۧ>gr�����q����*�^����|�C"ǣ1��E�Ytv�.��v@giO���
	�2cSh�8x���V\�Vb�3
�� o���7]�����V��[���W��z�^(��2;�	��]ܝ�1&��/F\v�]Uf�و�Q �u5VDw2�~`:���A�=��덬����55rt�EX�����,��g������<��+��^�u��.-��R�Ѽ$:FʐumY�Qp^��Qݘ�j�X���dU�<]x��#RW出�}B�W-���k%�
�_Xotpx�	�Hc:x��NjVOcBk,A�dV�ᕄ�G76��j�:���3ό������.3ߜe�⍊G�d<�4�{fI��e���XÐ����c���K���U�5{�^z�d�/=F��Ug�! ds?X8-��+��ʝmެ�5��8kRot���_o),��)LAK�-��؞v8	5q����_h�N��q�Ř�������J�[I]�k�z[M�Ċ"�YFi��|3�߲>�����P�qRR��}���۱��]v��m������nΔ�i�q޽��YJ^�SΌ����=<�/�Y�%���q����M
;�8�"��]wE���N��
���xq�k�W;�r[yi4�US�`�R2M�=Q��g�N9�m�UҞ���{AȽ(�Ot�<����P݊Dp�u+��٦djr��v�	v���s�m��+�c��k�؅]�Ѷ�����H]{V���"k�9��}a�����p�s<� \���A�2�N����,+0)���5+��2FS�}TYG�)VnCL�ͮ�N�GG#œ�Qp0w&�S/]c��B�\(���	{�����v�m�	�����\9a^�^mG	���ઋڼ8�X;	��t7�S�K���Ʒ1������M{ҙ�rǵ��R�7���{at�Gݛ������xz��!��b���Գ�9��[�]�r�s.�mM]�^�ط���!�����O4�/�W�%bUj6]��3�{˩:�һ��ӝ��&�9��jk��yU�o�W���ߋ���ٳk�ibL�}�̠�'7��e)���̎��- �.J�u���q���o۝0��!@����f���
٩3!�C{��ԛGFfʧ%Y�Q=Ǖ{z0�0��M�E��K{�3*��9���J�)�Hjϵ�=h��Z��qQ�C��^��JA�q�j�d^0��b���Mq�neD'��HB�6��'$����i�f�Φ���w*��Oz
��U����uj���wOq$�(�y\+ē	1�8^��Ͳ|��V�Fsδ�nE��(tk�z��ݷ��o�."r�O��>)���6���5X���Y����[0�D�����[��0�sM��^�ّ�+�v��kI�N���Lwc#'�uPZ��{��V������L�\�IH���:] v2�̈�S][� U(
�=5�s_q����mwU�W�]OdQ�f;���]e����LI��٩��;�j���$(�5K�IG;�5�(,RhF6�n�S|����U��X��$Ӆ�$W��vuz���ғv F���m�[4�#�����u{d��{gG�KYd_-��y��s�w�Iu*C�JW��B9��]�wP�����k4JmX�p.x�ӁV�:�{u3斎���{�&:�{������­�t5[7S�:b���ɤ�#���1�Q�gm��9�,��{o��oŰQ8H�#FTv(G�Vo+i�E
�M2����ÞB��0o�]���t�b�a����C��R^ƫʉ1~�1��f�$���2��
�d�D�w��Rg�� ��<gt����)ǹc��?:d%�D�/&tOID�}Ywൻ^|i�8=<�`�"΂>��j��]|o	�$�f�E�+��pK�t䲏Z[|~�϶.��a��>�:4b���E�'1���u���̧���S�N��;�kr���(G>N�(L��t&�{�4_t�)����糕���:�MeA̊�B�.|e̼e%`�󨷍w^X�tLe3��l
����6�H�X�)/�x���X#cW��MQzJ*�㜢8�}���ͲV-J�R�uJ9,h���G>������:)���D]���&���j��F���G�O.;p��wn�2[��vu�cg�J�\������&�׉��.�|M�I�8)���g����N�g����؊��c��0L�Z&)�����ħ��Ǩ(�t�����^2&��\л9�Jؽ�7t����2u�U�;�*��
�7�~��_e9�Q!Ʊ)3i�Q�7�Q�mw���^�8B��Mp�}�t9���h���,+y�����N�ǂʲ�s�^��f;<�Q)G��ySή��dp�&���L�{P�s�+LQhpF�*_^�]gV�ᑶ#4��P��N2����r�B�/��S}ֽ��/�S��vV��<�ӤMt�ﳘ���V��/bo�IR3�Ή�{A�Y�&�⽛��#�tC���*�6��U���"��kTC��'��Pa�˖������ё[�����5�1�y�lK��NH�!���NN��_uy��{���+�*�El�ē�Ƥwp��[i��t�]u�9$��]|w����hgy�b��"���"�
��!h�-8F[Վ�gH7ڏ(Vb������c��vD���q���RR3b�PS�
-h��!mG8���O3O��V;�~��e���:�Y�Q�=ei���'ώKጶ�M������'ڝ����L�\���5c[n��{R=�^���J�Tɼ[���{M�ole�j+�0bo�5��SW��O��K��� ���Ρnj�GtD4���4���k�ѵ�D�B�=�Da#[;�/0��d9�g�{L$GY������t@cbT�oj4B���W�6P�h����y@G,��T7yoo�2����۪NN���ME�G�:�y��}o�ʦ��w�/�A/|�x
6��A����u��M��e��÷J�f=C��]�R�A���54��!n0���n�R�V�9j �Ȟ�`���w9�!�<��vb��f����gy��z+]B��T�95K���0�21���q��Ⱦ/]iS<�S���l�ԉCy����$U�A��Y��K&�"��>IX�-v��OQ����#�WN����\����x-5�����w�JM�tH���J��������y��N�T0V�q�[E�rN��5t��&0n��ɾm��cf`�|����t���d_Ti��L۹�i�Ba�w��	W��:���ҩLK���iŒ�2�N)�i�����Z�Q����GP�3�i�ĵ��$�!�q���SB��4�8b~��~��v_�U{�U�7ݣ��� �	��jY�0ɘ�^�-�Y7v��r|%�K�m��U�d�3$-��	���7�E�|Ү�ͣN�x��'V������R�+H]�r�)SGk��E;�Ԋȫ
��C���&ޗ�4+��۵�C�2�֋��6��יk��e�O#[E��]��b� F�$CFM���Z[���żWcA��,$�v�Cv�!f4�'ؾ��)���*��y�/8GcDٰR��21�Ь�|+i�o�Z��֚�4\R����̠&�մ���	�x��0-�ji;�d�!�s72��	gt�R�#�qQ��9"[���Zե�;��M�yM�W���Ƒ:wchY�X4��8�`15���X������lS�ySHA���Ҡ)v�3o� �%�	/v�u�3X�p�} �Be�Z�QmJ@�}ì�� �����>I�p$Ş��-���_[z�@����f��b�g"��ͽ��XHY]F�C��^�2���j�cw	gru�"[:�;���쓶^m`�vhT���	���j�Z��s��IڗW�D���:͕�E��L|������8+�*������xmZ��I��J�+Ɯ��7��@�x��]�=F�v��/�L6��&���9�����m�p'��So��݇X���P΅r;l���p8��e��jo.&5[�T#�ۏ�K��|�$��R��cI�_+G^�r��L+�s��C�����IS�R�D+��A:o��[y>�塷��%\U�����R�� ���rI��s`�wƖ�&Fa����G}�l�2�^V��M(�ۈ����u�7JJ����JvQhX[��3:��팅��qF��)� ���ӥ��Ҏ[�CqR�o�4�KQ�h��.k�1bT�"��c�������],�����h�X]y,��fVSΖ�-Q\�a6�-T���ڹI�O^	�����Ѐ�Ӈ:s��-�ٴ�֗i��|��XsZdv�n��B��d2�Eo�Մ����5����}�b�Z�"�UB[AAV�m7��DL�EUX��l
�R�TS���	X�����R*�mqj��Z �E"ȰEIU**1�b5��-F��A[���0�+V8�a�0�1UfmTUAUp�
��
��
��a-���J(�UQEQ�ȉYT`�Q\��."���#�QJ؈1TQA9������}����D�;�\��[�P�[I��ܩZ̡���&6��w6��[����}s�����F�ާH��p��v�l27��
~�ǐt0���<4���v�,kg^����-8�\���	bF5��A%�j_H6(��%��'��QU��9��*�����0V�C8M��k�@��P�1x�i���]c1:���2Ng�3�>J�^?<$��oe��.�^'�"�gs*u�����9���u�J�͝�}5y���V�]e\i���v6�.�ې�e�k��|���Y�&/Uz5f��c���eo,�
D:zc������R��è�'.a�suz���w9�%>V0�{�4�U�g����(�;6��a�#��ȩP��HF�7� �^[wX��|�#h|�l>��F۽�c��O{:���*E{c�[�&,y�1���l�Nr;fӛ"(�nt윔�|}d���c�K拼&�M�ֹNd,{y����m�f��];=��ƌ��.�4������蹞V�t/`[���-xG���Mޢ܉\����뺪J���T�2y)v�ќwJ��д�l�0ս�&Rj:�E1�Z�F&��z��������<�V�)�4BEc�WU}{m4X݂������ʻuf"xE�Ȗ�Q�+��Ķ׵�]�-q@�o%m3]uWj����X#]�\Qp9�"��I�1y���
�66zJ3Y����/YR10�y	4̓��wm��hF=6'p�P�E`����p��`M�GgH�ɽB�h+}�1J�J�0rÕ|�c^����zf���j�L��Fgi�'�.�>K�N�A���8�"�gLV�9�*Z�M���y�΋)):tl��ٯ^h��əh�풹��2-�\P�=�Z����'����d�g5@�aԕ�{�P]q�\�_V�>f����:2��zJ@�+�f;���Ep\��/=��L��)3����/�5�.����~܇�#����v���L�\����)3}]���Q�;-���*��4��m�4�Z�:;�鷳�*o�P�y �E��<�����s+���6��$��4��&�n��I��(y���1���V>��ka`�D9�I>�<PԐeGζ�Vi�q�0<Y�%�9pv(��J?<�4j�.�mMu�8�o�����lb���c.�[���v(�=��}n8�<o:��6�`�'J�h"��h��;wNVwC����7KpVI��Z�r�Wb�я�˗Q�"�ѷ�}%]b�J#Duf�7t��V֎�A��{L%���ˣ"��#j3t�è�Ky:lv	���	1Ę��z[��=+_���[{}뿫�9����yum���κ����N�Y�ۿV�VK�x{�5Xz(rYg��%[ilM����Ԅ����eX^ܯ?����į1�o��Z��u����C$U�!��u{¯NH��m<���u�p�w���OQ�1`B�t���o׻ք�K��&���
41<��n�ts세�+=���%\#���hJ�޴�xc֫��ݛ;]�w�΅VNɈ+��6j&*�8�ʅ�P#H���!˼�f�]�w��7��Ie�c��V�6���T��r�)}��N��GB=�۠0G���h=��#�R��)) g�R:`Z3m��G�8��!���y7ǽ�S�cr�+��8�*��\u��u��y��}{s���b)��IƟG�.�*�#S���Z/dYT�SO�X=T%�#��7�À�k�}i�����h����<j�/j&PK��A2�Ok��˳vdj:���UO����d�)�e�P�0n�-�t�<�O��5��8���ٲ���K<�!ZQR�[���m1y�)���g�}Y�:�ܞW��y"��)���vk\"+}�k+1wf*�#�x��v$�Jp0?��*i�{.ɚaU�_��>��K�'3�"��[�j�\���Wܗ��N~�JFMk[N�7�Ct�z�Q|o�߉������x�|T�a��^��ַ�J��iZ�$�t�qh;sH2&S��k�į���W�B�k�D���At�@첗&�-1>�u����F�y~7��h�1�4���.ޞ�������x�������॥��.n����K��Y����Գ�gM��or!�܀�*�c�=�g�WPh���k4�q�����ŷbUi/�f����l��K��{�G����i��Mv�Jnw�������py櫾u��/DK��){ؖe2����L����x�P����-9Y����T5�iʯqT'H�Q#�q{�{ưg��Ma��:�=u䠤8�T��X�x�o�q�A�rg��˚zu�&�)�F۸�+���
�\���׋�B9�#��OU���tnueG���u�1�I��x�s����J��f��q2�7sv7ǊB�clp�]�V���.�18@�z����O."������U��1aD#y���뫥67�i�׮.�M6����Z��I8��[N�z���]�	�c��L���+��ob�}AcoQ�-:D�\����av��>�ε���*���w%����ٛ��a�Y���]�'y[BE��KRy6��<$��Ļ���ث��-`�w�R���>��EX֔���W�ܮ*�޿ZSp���h�2���Oǟ�%x^�wCۄhL�J�.�1�
��1��j8��ڦ?����JZ�?r;��\�͋��zb�ٶ�[�}
�
�;[�\�r�,�Wӎ��THf�*�;C��;f�-�'�]��^v'�Zx(��WOz�)���c*U��R�{�iB��7��I�����;�[״V_([z�-f��t_�3[��LuA��Էg��ZG:�:��2�c���ϜF}|]�K���~��ăP<��&��P[�g(�����N3�<X.�`f��E�8�7=B8�h��=����g+Ol��)�Q1���B��0��z��G�gs�y�\�;S\��ԑ|	1d�����!	�˙}��DMw?TN%����]�Q�Ւf^��D�1$Q��5�G�2�G%z���5;�Gޫ��y���+*�~+x�1���9
�mNC��3ݷ]>Q���G��+��hq6V�.�'��rk���EْL�w�(��+Od������'�o0�V��8�5sW*	���K��\W$�\���Qgl!�sb��ֻ�i�5xb�VՂ�͢�XgZ/o�ۯ#^3 B�b�q0�ot��\SZ$?{xU'��5��>I�#�y�%�.��ND[���^_������ZN�=j�O=tj�NZM�BcD4g�ګk��|+8�!�(�Cڮ$y�L&�Er�{��W�.:���u���]�"˞����[��6�8/��Z�t���傋x��	�+u�8$��K�@�//Ӑ�*{py����V"'{��\R���/F]z{]�N^�.�mci@�:��fȵ!9&�S���0w���.' �K닱8)�N��TES����	���u�:���e�qmkW��r�ᵠ���=c�]����Vp��9��ڄ�tfM[}G-JV�
s��ѱ���`�7$�*�\�]�����ĩ�B��XP�����ćt#y����.���jֲ�yKJt&r��D¯x��JSq)wFwg�ŲO|=O()�0�L���vL�ȡ���X[6p)�ŗ"����M�>��bW͝�}5�ͨ"&0`��γ���3c8j��jޞA'�����8h�V\��x�r�sDMot^&�︼N���͘5�Mi���
;u�e]t��i��U�%�N&��.�ͫ7Aѝ��P�����c�&EWI��y��͒�Y��7��ΰw�YY���q���@C��@T��V������ �{Y���$A��E�T� ��ah�J�T���b`X���_Kd��++{��x&90֦�j��ր)D� �D��ZD���$�$��g�c�y�������}�`~$O�[m��̩cl��Rպ��1i-����z�D
J�՝VV�\+�|��l�IsY��}R��I��
/8��ౣf~�3���^_j�,�M[*�����
���q��9���H"?�5��[W�vI��Y%$�:��D~�I��H"?(q���Iwlq���4mX��~y�Le��ۚ��Ns��r$�;=rH�#C�#��;�Gj����3=��t���zi����,����ZLi)�嘯I�0�-n��Q�GK���3��_+���e,�W%'��H�"�7��)1�{]�/^Xd�:�D!��I�$�9U o�Y����)��.c���9�82���0mz��F�2&JUUIgL���ˋ���t<�1�^�+���jLN��Q�o����>X��61{OS�{~��>�/��ݩR��y%���xt�r72v��Go8o�ݓϲ�̸Yt�H���ս]|�uw���&$���~���_l������{��RH�#|:�%�/BQG��m�4hbh]J|���DYR֑���DQK��$A��R|���}TNUiUdt�0�=�cn	4�)��#s�FMגIFFC����(��/.��$���7J��"����3���e&#=MxS\*2��Ԗ<A��簉I=�Y��a%�7>�4�*�z`}���Dk�=.�'�bGRH�"�+�ܓ��Q�r��R}v��M�|Q�Mc�?��8"�~��M�,��z)E���OFök�Q�b%�c�F���a���I"��9��
��֋Yd�>�i�D�ى�qZK�s���p6Y�٭7�l�%ۑ�឴g��Q�/���J.K�e�M���Û�Sm��֣���Um����f���8+v�중E���������J��ݙb��N��)��n�M�Q�QeVgו�tb� ��LR;�GE��D�'���=(�D���nW����Gl�N���&�(��dc���$�T1������Ŕ��U)E�����cj&�9��ܑN$!�z�@