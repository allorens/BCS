BZh91AY&SY���t�ߔpy����߰����  `�~==�     ء{)( 4��{� �   (      @�   
 8���:i�|  <�]��x��f��hi����#�WC/��sl�M��C��\�v��'�>�*>����=��:ts�����ۼ�z<�=�Ǯ��n�ۛ��:{���d|  ��R���ܭ���{���׷���=^�����g�Ժ��n�'w��ٝ��!���Ϸ_{��[��ʻM�.�7�nu��w�u��w�޹tx   !�n�٩��(7���ݽx^�t�۠�;����w> 8#��ܷl;p���vu��-��]U��
wf��m]�\;��  c`y��w}o>۶��'���l�흶{��ݺn��Ӿ r��s���\�w{�{۹�ڻ͍N.�m��8��һ�   #د=�n�'��ե���u^�N���^J�o ��g�������p׻�i}{�ﶷ����4��]���T�J��P�P   �  �h �@     ��F��U*P=� �4@��i�5?B"IT��� ��� �0!��A)�1J��`      �L$�@%*��F�1�4ɦ��D� �@���0L�=���21��6��0UJ�F Fb` �;�Ӻw��K!k�b7�٤�&��� ��F@�>�� (�P���?�(%PQ�W A��;*���/t?���b\t��"�F(@`�@:����*I'�n ��"�1��`A,�I~��-B"�f)�C�z��!�O�׋y>�٢V�5���>��Ik��ܶ��<�
7��W���I����'pG���ݒ�7��$�lG~'>��jt��\��]����z��b��`���rZY���%5��=�ɻ5�ɤ�o$�r�:�N��s�d��ѓ�;�Np�;'vr����-�;%%�5��ǫ0m�U���C=5�u�݇65��7�M�B^�#�p�[&ҹ�h٤�	�ᾉ�E ���k�x�ɴ��=��%$���O	^d�]E}��&�Ȱ���;�D�'�A#�+�<��d����)�<> ���K4i�*��DOlD����/������(~�DNq"'^���>M���������'�x�n��?Ak�D�D�xI:H�CZH�H����D��;z""�(~����K({�:Gd�=,���"x�����
a>Bp7I9Ĉ��6k����t����3ĳEi"%q"%)8h����DMA�� ���D�����/���N?'D֒QǄ�=Y��'D�bDD�6A��&��%�'d9��'ւuN�p�&��"u<v�d#�~�z!4i{H�<$���l�n��O5%wBl�k�	�М��<���'�O�<�+��A��rY(G�v�s�8"v�t֧Nvt{�#��NT��pM�F�bwR�d=D4��D��tM�F5<^�NnN-q)�J;��}b5�"y���f�4;�#r��Y�=�~��b{ӂϺ[U6j�Q����{-8���������[��J�#ԯt~�d���R"<����{�>JI�8OYeh��F�˩ѩ��8/�"^r��f���L:�'Np��w�ԳW8s�N��;~��,jʱ&�����5r; �F�˗iw
���Н��v�#ٱ�'j"<$DX�a�6���'�#9QgK4Ϡ�Duur�	SU>GUQ��Dgj'GmO+�uQ8oq�"S��T(�D|H�)�FUDG�����Br56A��d�R���D�\j|�$�c�DG���I���Dy���ډ�kR����������˨���7��d�z����xg�"smK �|�ʩ��A�TK�'^T����"/j'��J�jY���U(F]DG^�T"kmJ ��#�TD^ԡꈜ�R�<�#�zMF��f�G�v��j'y����9֧���|���C�;��N�~�ӿD�tʁ�h:��tѪ:kz�Q�17Bj%�"76#�c���M�J���
��8#]����O�NmM��
gӉ(������y>G��&
���hң:h�����
g��$�4j�Q͏n�?pK��d��j ���5.�IIgv��Μ!|JM�)8[�/�.J����S��v|�(㢃G.����j���s�,Ʋ��;�w,�sl�0�e��]4v�g�Y���}�gV��۬�Ah}P�Q��<�G������x���H\�nG[+b7Q��{ʋʗ��ԦNz���i팋��>�����:�g5��T�j{�E�E���w�WjJ���Z_�'�o�y<���t����jY��T,>Ju}���_t�B�7�t>�_i�ߘ�w�'I��$A�>��l{6T�D��I�M}&����>�C½#:�>f3��o�X}�x:�U4C�Xϲ���O�X���;�3Y���̺=������ǡ��Q�b�܌���>�g�;>f��_��i�/:)�1z�{�.��C0+��#>��XϺ{���3�y��:s�}|�M�rMDu�(~FD�ޛ:�y�4t��pٲ%�W�#����n���K��-;������<t]�x�����Q�%|����lM��+d����;R�nxO�+�z?J�f�Q����d�G�����	�֥|��Q���!�gɿ�ƯR��ȉ����N���D�H��\4V�${)���=%j"=���OB�'���u)�J}>��JDӹH��R�X뒾Mh{6"k��bm�	���7�W��H�{)�et�����]���ʳF��%����r�hu��'�JDӹH�~���^,u�_?=�B&��[o%"me'��|�R&��D�[,ټ��h�3�w�M�Z���W'���r2[�	�eP��UK�^�$�u�5S�$�c�ʣ_#��F�T�;վ���VCԪ��U:|��G�v�Z'�H!ʉP~}U���__�j����F����H��{̮�D}�^/�e�Z'�(� �#ɾ#��:rK����By���Rh|H�US�I:q�~�l�RnYR#S�$G����U\j���A�J���U'�j"�:�?'{ �C�#��N�t�z{�5ͻ��6��a�b:a:Zt�:}��i��;Q��{��Ϋ}��y�h�f���sJ��+�V���ߦ��;����&*�Wj���v?�|����v��P���ý>����P��1��~���՝�{O�T�Myi���~��5ߣ~�������������;5�w���V�K�&2��M\�e�s��ߥ}����M�Az�n�D�p�N��ĝ��&�/�$�>'���e�_N��	�l����/DY<$�ޜ&��[
�Q�No���&vx(��#_��(��Pd��T6}m>Y�wե�Nȳ���9�j����k�\P{��6������AN��&+���w;w������Mȶۺ��y�VwY�����{�B�☳�=);���U����g݋����/�|o,h;�R)�O�]0����jl;�{~����n���{Z����w���}%������6ɜ�����W޿M���W�嘼�O������c;���l�������EWani�_X�W��+��벗�	����f�۲l;u����w�}�����޿��ߟ��ۻ��}j�]��<��nԏ����dѝ����dS�����I�Si����=��a���<;p��_:�ϭ�����~|�>��sÞ��O#}>i���s=�J9�W��������x;�5�R4�I���o@��ӻ���:u?[�́�0�����o���_��id���q���gWڤ�ˡ�{ꝩ�s��Nm�Ny�����w�9���\�ʻ�O�&=G+����񧽜��7����׻�w���Q3�y��{��~�M�]��\ɖ�f���޳Y�z�랸�	���y���})��Q����.�2wl����d<u���ƃ2魆w�L����K�{�ow�ܟv�;cc�};L�K٧�	���������3��y�g��i�����gU�K)�X.����k'�3��no�;���N��)_��w�zE����8��.N���"k�oн���޲؎��w�̿����x}�役���Ǻ���h��۷�k�z���h֎��3��E,h���Bz��'{n>���3�Z�f�v̙��ޛ�7�Q�`G�Es縲<�ʼ�eO�L�ys8��Zǽ��^��lY��N=Zw�Օ罛��S�=�$��io�:�u���vn���K���]�,�5-0p,nm��W��e�~�[�y{�q����e���w|&�i�5�K��"uڹ���;F1��^�X3�3t�m��;^ZB�d�tF��h��س��{g��A���׽b�{ �x-G���S׹�N<�����skF���@��i�-���Ǔ7�>ܛ=����;��μ����}��C;�w#��oo���K�O��3$5��w.w?��3�Z��Ħ��C;;�ݘ��fm�c�D������w�c�m���~1�=�c��k���|�t���]ڽw�M��ï�y���sp�vvif�M�M�]���
=�Y\�+��ɋ�6ۍ�w(��ᩯ�=����{��]G�;��H8ޱ�b��8Z�jb��B��Gu���ݱg�~�ӹ7�ǝ��<�ޛ�>����,կ�ۍٿ��d_��cA�9�=$z�)7����͟y熳]O��YܯV~����~ڣ�O��;"��u��o���Ξ3�X};�+�J<��b5ײ"�M�JR��i��߲���W�sx6�]�=v{��d%��R�1Ϗow�g�gv���kT��Q^��ϰX�/���M�9��}ٳ�s��]������bss�g/V�ޛه�7'��o�;߻�do��/!߮�}�Fu;:����g��uS�~�O��5mqc2/�s{��vOvh���b�����O�̞����w�.ɒ������o����K̼�}'��{Ӫ;x��v)ܿ`l75Zwt�o�z� �\�vs��~ɚ�}��
;2�����jh�/�\7f�G�vb�n|���zA���(���w���!���-���o�W�Z�����{�ݙ�T������tJ�o�`�k���;v_�^=�3�����d	؞���1�KG�v��7�9'g{ٻz��˔���}�g��y��4�2�ze��ƞ>;�N�^2\�:��>ߵ�������?{�47���쵉>Ÿ�%õC������5�����v2ٱ�DW_r�CB�����'z��\��aKm��P�k�����H���t|"�����3>��lw�_f�頻\��O��p���n�r;�������ڝvYFӴ�w��:���_HgM�ӽvu��	��g}����߇�}�g��йn����N��6Ȧ�����E�3s�q��l���:T�\���5�3;+��o�|���o�n��\?Iۛ�#��GUt�a���r��.d�9�;����f>����u�2K���;i���юhJכ#���&�L$�/m�V�f'��ty���gN羚�_/��^͙�!t�?��_��\}%O�������W�_f��`{ޗ慕��svsO�e{�o~�wN���������m����z�5�L�������+:����w�J�h�j殮�w���ʫ߷��n��'�r�N�������ͽ�����Wt�t��߾��|�տ�㰈k6��s��]������Oz�~��G�>z�?�y��^c뙛b�g�N����m��N�䍃�ߖnV�~�;ޯ��2v�g~�٫Q�=�W����z�������o��iڲ}>�3��]ۿ^ϾW�_�x�%���ӧ��z�X���V�;�=x3{��e}�������jg���+����Wb�{��.�sŴ9����j�����Mh}��{�]�ٍ~���_5����������&cgY�S�`��ӻ����=��Qا�d�n*�cK�Zy�{���3�ŝ�緞2�rǙ�̝y~�����֘=Ů}=��5�k����~��z��|��}ڱ��_ww&G�3���پ_O�} 亽,��o�z_�>������\:{{�_k��}�{�`���7w7p{��Vy�}��W�6}�wU�w�ӽϟqQ��!���۝�l��z��>kۑd�<�D^�{�t_{�y�����u0h��ە���Fx����j���H{������s�~�)�E>��ƪ�s=��:u�}o<L�~����$V�~�n���}7rAu}�~�+�|ft���w�=.wn���5��jR���lZ��������T[�ߟ�l���L�c��3�p�z!=���������HNΝ�gNpc��6O����swo�Ic�A��:��ჃE�x�%w���q�$~|��œ%mB@Q�2{,��*fخbM���mG 
֥!㯹�+9[Pb�,R�H�#bht��Q2V�j��yTE���ŐŖ�4�7)��N�B�JE`��N[�':�՗�(�ヅ�AɊ�#�d�1�w0Ơg$�WN^Y\S� ��&J�BrB��l�|(�l�+��*����Z�lG��u^G%����+�!�7k�
�DF�P�b���T�Ȭwr�1U,VGN)(�8G�8��hVq���br~j�%S��Q,L�I�$,�R���DB� �*`*;c����I6��X��N�9pm�MH��X�<�#�9	UUD�mHW�HX�NB�J���U2�!NG7j�rI"��bɕ�1�U%��K)Z�AT��s sF�[b,U����xq>Fے�(�������2q��GZ�[y��1��(F�A60#�@�TW�����r�rL�}Z�hi�쎺6(X�(�US�;���Yƨ�f\A ��ʊ&��E��C/<�bRZ�R��JJ9\v?�.86�\ ����L�PQW����5��D≍�%��d��0�We�c?L����EA��Mq�li���4x��S�#��D�NJӟ������|��� $��<Z#�R9��ݢ��3/$9:Z�a�(���5+V��3	g����V|�fd�,���E\�o�S��HmT�8ҧ$>��Ր�^<�S����Ld�IU�e��$r���Q�4>:Ӈ;���q�Q����>��q��2�r��*��&�±�h��[M��B���n��t��tQ�KJ�pM��(�۳�Zh��#��&�6�<"��5b��ղF���5��#�[�B+�cO	�axЈ��B�ԟr��;��+� ^���G�+y]��(�X"E�+��%��9ڜ+C��![u^N��G7�[�:s8̮8:��/VE&ŋ+±v���9+���1��%�z�LT�k[�}���B}h=�O;]Ŋ�W��ۜ��S��@�{�`�J!Q�ڡ����=���x^�����@*�*|~�+_������UUUU_1UW�J�j�V�UꮔU⮕W�Ҫ�UҪ�ZUW�UV*���WJ�Ŋ��Ek���U^+�UW�UUTx��TUUTUUTUU{�m �"H�% �������I*�-T��!hŋD�A���Il%�C�C�eMmU|�UW�U|������]*�UmUmWj�j�U[U��]����WJ��UU�ҫ�V�t��Ej��UUUUZUW�Ҫ�X��労��UU��>���X�@�QHAR �d�O��>	�J�U�Uګj�U^+J��b���U^�*��iUU�Uz�������]+J�WkUV*��t��U�i֩QUUU�Uz��U�Wj���Ux��U�{��{����!;T��)�d��'�BT�����fg3*��t����Wj���j�x�UWȪ����������������Ү�W�U���ZUֵ�UҪ�UmWj��]*��iUW�J��ZU]����RA�@�T���WQ��h 	QEdE	@jHD`(BZILP��)�TB@v�Td$]D��^���TU�@!>�����>���p����c���y6t�GO�lO	�<'���"'���"%��"h�H%�<'
<"q�,M	�6hCDD�"%����"%�b"xE��'�؛f�ДA8%I>A�	%�H��,K�lCf��� ����,��B"X���'��bY��AAD�&�ѡbhL�%�=���T~���Y�2�)���Ip�������I�j�"m4G���+�(�!�k	S��P ^�%�b��
�b�eS\���fr���+�I�YG,��N�*�LP|�̬pl�<T�Ȫ-�H��T�2y�9�+�N֣G���X�LAaI,T̳�4ZFIH��]���ش�'�u��T&���Pm�8���R;%Y9qe�2��I۴nX0L�¶�������5�'\�*��b�)c���, �+m���1X�Xr�;C��+S�̌��A�YT�^'fJC,m�b�IE�n�##v'[�Qa#��r�Vԩ�i��G��� ��N�AZ<���	d�N�ь���X���#�UE@Q�Q^RpQ��TE"���I(��Zm��c� VA�Sp��
�@vIcv'(��u8ו�(*�MA^ATEK�h��ՄV�U84� eI��:o((�1�q�Ń��<-7��eַ���>پ�����(��wwk�����������ݮ}�ffffb��wwv������������ݮ|}����,�çN�8a��tO���D�nɪF��,R@RL����g�ӶDN�;��S��ͱ��ŋvG�"%[qV���g 2����	9%`��X��N�K��w7\b�z`S�� �I	��l���	�q;#e�?�'����~�O�P������v�[wKeJ/C$��(�qW4\1��J�	� ����{7339�"ōU0��0T9�o1��`�(�Z����b�df���c�Q�i�ZR-����%�ʓ*9UVt/���~���:B\�w����:C����f��8`�xO	�<<C�{�������#���媬g�Tpt��������T�Z�ɹ�!�K3�$��I�N$SF�k�MZO�����M	�������x;p�����~'�H�ʤ�#9 %P�m�r�&�Q���ـ�Sw��H�Vh��\"\���j��\���������,�|�m��M��F�B���8�ċ��`��ئ��J�Wϕh����m[�3
b��㙅ʞ�,ɳA�a��J�J��c�y�T��m��z�1	%��%���M�A����W�_S(��l��t�v]���܅t�=ئ��,,ߠrv��nF۪��~Ubԃ���{ϰP	�9�ʪ��O�m��i�[h�J�珙ַ��e���U����f�|��f��/+e�������WE��ƪ�Ŭ�_-���h�Z�P���,��n,����V�rjx��LMx�����FΘ��Y)UGSN��M��f��Fʳe���e� ��}f�O#Y��Ï�͸���i��u|������E����#�c��2�j��9�ׇNK��ɝ�h-M�70����V��w-��xŃ������|z�ܪ�X*[l�����M��3LQ�J�dh��UP+����U>C��*�
W�AV��67ƪ�0Q�d�t 9jhE��T
J.�TF嘆6���6�#�rdRdU3 ���������uTpm��f)��3e>g����(�72d��¦��U�fj(�A,Ձaþ�����w�a� &�&Z�
*� đ�5jQ�r\8DNl�b1�Ǐ�i���8ۍ6�l�Ѧ���9݅S��wT�4��*���!s�0|ś,�a�eWC���{ֹX7����Erv��rtɃ>�����oP���9ŔT�󊑨D�)be��l��I`ڶJ�hܞ��6]�΋��L·'$UF ݧ����bg>6l��x���xO	�<<C�Zѩ9� �%V�7m�� �N+��6�ɦΚ�V%�q��ӻcsk�N9J5�%P�U}�D�9Pۮڠ�P�a(��)��-.�,�1�����*���H�Ro�1Ȝ//X�SUY����G�g:T���4b��F�˖ba�i���4��Zm�N6t�p��4X���W�e���&1E��ڼUV80K�	�]��oX�m�)%jD�q��J"p$��9Q�Uũw�k��|[�@yjw
�h���j�7%Æ�
�[,N̞�P�ѨQp��g=lpf�FL�Srv�Cm�k0�|C�]���}��,Ç�&�tO����E��>B4I�X:���(�x�+�Kbj(Ӣ1��˘�r�ݴ�����,rH��)2حs܎��-���V�`�X;���VV
�8�J�p� rC)���1�CQҩ_".8i1x� \�7%Ɉ'zs�n�MX�1�KV���g�1JԦ���;��T�Ƅ�0Yp�J��:Y�bj=NK٭0�\2`�b�&����V�Ĉ��
GdN������N&�Cd��)��1`��4��m��m��4Ҳ���׺`�i�DV����B�U3�&!��tܜ����o��C�=��`ܘN��{59�2g�l�a��iwe��&��{2A���x�54X��+�\�RTJV:�$CteHnA��"ژy_��v��YjL�%M����Ƽ�a�(��		FW��H�V�(�95"�~�&����}�����N8?�M�u��ë�uv�m�K�L(�&��酚�a0�h�0���x�'O>�%xG�,���>	��^���<;<T<:_�������>mk���0�F	�V*��0�aZ0�&���t|OO19�>>b&��l��ч���j��>.���l|Z���r"'�Q�M�0⸳��~Y��8�[z��Uzpz�P����x��>�g����<;�!��<X��<;<>!�̞���J<r�G��̉k����OS��g���|��bP�]u�U׬�a�z�W�Xy��O�����3�gZZplœ�cT���su��+?�����!O{ѓ�c�{����0��7�3h��h�߻�?�y{��˽�G��}�ޒ����΋c�I�G��]ܭV��=f����W㼜�9o���%�đ��[�}M�P	�o����*��������3&ff{3Ȫ�{��2}�fUffff{W{���|}�32�31�3{�����8t�ӧ0��xN������a	9�UUUUEr2���L�ڪ����I���O��.N�r	9�%ġ�h�wC�/��x���yU�5?,�%11u�K4A4Do�R�E��J���9.�%�/323����H�n�"���*�_�U�RB�%"B+d�Qx��C�⚢�i��������220d(N�f�o��\��xA�c�;Y*�z�^���N R�.�H���3B��q� 8'~�v��E��~��0b"�ц(�UX�dz�1%K��_:���e�Z|ӇmN|a�	��p&n��UU��T�~��kp���؛f�L��VlFQQ�_K'�~���Rۑn.AU�Y
r�F���>Y4���1�����$Wm�n�@��r�-�.�Uq�E9��b3������ؗ�\I�H0a/?UOV��I!��=sx�ʌEqa1)�a�p��d0B��F07g�p�0�`�!��b\�&���b&<�,L���eI�Vᨰʟ,U�Qd�V*6��6��q�<'D�`�:l���k^�ܦ�፧$�e�����LMM5B�&J�!k��~�R�1R4ܸd$�1<M��r!�tō^�z�m�@��e���zd� �Q��`ܺKD4Mav��^sʪ�!z�h�n\�ݷ"Z����TL�s̩�<F�Q!����9`�$Ct�0Y��BA��ДX��=.%hjLA�1(�J����qU��Ca��D���!��q�/���J)�!h!��)��"�(ʆR�LFO�0�0S��H�`aZ(2�6�UR]J�'c	�MA�D>�Wk��5kmc�5(�rFP�,��j����Jd�����B0CԴC�|��u��|�n��M��F�:'>0��DKn]:�����UFY"��AwsSU(�� f(XT��`�K�y'U>e���Y�}���jC0`dC<Emg�z�Q�ꙑbx��8U4�JSTa:�5���O��7�c#�dp��74a�EY�4���d���2�lB��1��H�/(��7��%g$��G	t�>+wl�����r�'Z+�"	�H��(R%#t�1H�Q,2*,2!�atY��2亁� FG=}�-�)L�.�L&��D����N:|��\i��e��8�<e���Բ�z1cM��T��Ϊ�����gc�E��R�}) �R|c�K��:!�!3��S`�|�Ҳ�,�3m�}	I쥖D`z�Y�%z�Q.թ8ñ����,C�]4�P��\HHI7��V�V7A	FD�2Q��ܳ0d��eA!�@�&"i��2fP�jP�,$]Gd��!xfSKDB!��U|l��A2}G�T�����s�>0Pr$�0��YȂ�	S.�5�̳q�
-D&Ve���?,5���S��i󎿇Ϳ�Zm��m�M:�L�~c�q�%��'�x�5d�of�~UUQD4 ~\*%��V�7=��K�*��X~��a��ƹ�js�������3Q������&q�#�Wr%��s�8�O���l���r�8n4�p!�f��\?2�9>���җ��dn��+E�ʍ*0�M+Ǵ�L�Dl�G����聢Q����� A���xHR�l��±66�#�c$7H�	Q{rV��RK$��h���c3�!ET��\���z2JB<9�	e6K�F!I-	��ފM�Yd�i�>q�:�m��mp�>0�3�_Hȹy�2f`��l��cp��R��`X�;���Ob�׋d�""uMǬ�ܖ�B�w�z�o4�I9F�P�L0���V4�ow��(��X�V�\�q��m��ջ����H��w �bǐ�i����h������6	?!ph5Tj����]��݈)y�E������h� B'	�baC4"�h��w��h��M��JJ�r+2��@�Xx�ߘ��9H$n0�sm��w�&�a��[��W	t��a������Q��Y��X�M��!��P���ɜ2ʬ%|s���$�{FM�3E�SrV7��\�di����Ăj]
��b'�@bv+��|��J~�Lϗ/&bǓJӮ���u��m��4��p���J�K�e���<UUQ���I����f�r�����.����a�^Ǐa��+ذ�#Fp�����X���3GP���Z�l���g&O=r�ta邃pTca�����g�ϐ��/����d	 rX�bE�.(��=��}��Z%I�8fh�g�PlƓ�`V2J�(�b�"�#*���~w��b��OVU,��I�fJ�loH�$Nv�����a9��i�N���i��eӁÇ����O���1UUF��JS4Y�4�R�.4�Ct�����a�*h�r��I"�8�1bɵ�G���Y;j�,0�l�������n����������h5� D?}M��M,j*�'�d^��G���i�U7Q��Q������ïc\,N�i���ī�Ж0���7�J���,��s�e��E���j�HvDG1rFR�E2���h����ɧ]u��m��4ӌ4��$��ŸnQp`���R6,5 �ǜ⪪��(�U� 9�U%���|S,]�X(
�o	
\�/	f��,G��.j����(��FX�-��-Q���C�l�Y�1�4\ͷC��y�*6�tٻ(2D�j �(�t@�b$>ab��0�%�n{z���SWT���a���g����������	ࢉ�в��D�!�p���:��Hr'�SV	0����H_IKF�Dd��?^�CD?G����с6?�~ptt?�J<`����'��������x�^:��X��p�L4a�&+a0�D�t�Ba0�Ch°�.�a0�aҰ�0����>+�8���FG���~��k����8�^.\cn0���	��h°�p�0�"C	�`�:&�4>65���x����d�t�ŕ+�+�BxU�B8g��M��'�<3á63á�͜*d�H��`h�3�pl�L+��`���	��QXHaXL4f���a0jL �	�Q�J8aZ#bxQ�'����|)�S��|(��(|3Á<`���O	��<WǬ�o��4��mՍ�?�6R��@qV�f.���}����~�ǯ:�}��ȟ��◽g�b[3^rb�f(�d��B���>8�8��4��|(�{�[L�m���U�/��9.B'�o^gM��ｫ�McI嶊��O�̰�m^�n��l���M�e`ԑEkq[8�cU?}��n`t���dvLi��g�����}㽜��#�BډE6���~�1,b�m<v��5'ү�z���~딝��E��CsgMbw>�vwݵl73�Ķ���mV>�����DA�6o��N�]��G�j@�8̞=�]��5�0%��H�q1����'�����O{q�=XL�����K�}{�vי٭��<T�s6�rd�o)~�������U�}�2��Q��#]<n��g��c8e<d˖��54��-���$㱲Ѣ�P�{�t�`��B�UXE:Ej!:KPp���.Z82b�X��ҚoX�#m��� rN�%m�����VWG�Y+r1�� �v���4誇RNZ6[D82��1��ל�*��i����G�Z�G�N��#
Հ�ڭ�h�ʳ����u��%����tCDSq�n,س=�]s �낙9!̑�J�	aI&��O����ߏF~9�32���\>�������d�̽�{��iU^�Vfg7��3�2�333�����3=��C�:t�xDN����0鳎�+Z��J�����Bu����k
67��Z*n.I�ݏ�Z�!�3�ũ���<������U@i��!H�&�dqI���8U�%+�X��θ�`�bz�m��%7�|m��rC���qEDb���d��n\�P�-&�FL��!�Q�غZ���j!�a�AA�dX�PLp٩�lO���b�\!��$,�"����	IB�C���9��S%��,�.Q�l�sX��P�*g6!��s�#�J^�@�K."C-?	C �"�=�.jP#CB ��U?���FB�"h�j���j�+j^ay��P��]W* ���RS���<!�3r���%�4̟�N�㌸�-��N6�-�i�><|a�qF3��UUIEr�Vr�/!t�g�*��X���˝ﾫn�N��	�a��C��C�آ�%æ������2)`ݺ]��9b�Dr�)�K,Y[��jP��2b��:b���G�ne��9�d�FKt�z~�|�K7�i(�d�b�7^x0��2�&�#�x�'��������2�}�,�"\ֽ���d�|uQ���#����^�:ˍ��n��m�����6xو*v�SXCWB�f��X���	R�������D��'���0lj(a��rkPf c��<��0p)�h�*�9]���SH�c�D�~/Q���xܐˍ�1LL�5Is,GKVe�r�͆!%4}(� r�����\Ht����P�¤�X�&Cp�������$��ay4�K���*`L��p8Ma����r��͜��Bũ0`��[�Kf��d�]�y�;��2Q�)t�T�Y�z�׭����8�l�Ѧ�|x���^�ZOha)����ت�UBM�K'&(��SgE�3�K?l�0>!V@��ڑ,QS���7Qa+�	@Ģ8��y�Q7ęLd�7�R�4d�D`�~N]�n��<��fO���@���&�9nR�ˍ2^#�!�3w���� s�B;�$v��I��˷M����#)����@@��*���C3��j�)`\1& ��S�Gb�z���x���e���N����0�~�rJ�w��ZX	��f,j�ׄy���V[嵴��B��׊>W��eS�j`�{���nq��1��y.��d�ݑ7J��i��D�H�-h�C���B%j/=m��m	\�tp���F
G8[wUx�c9L�]�|���[5[�A��J�.\�>��j�0d����E�ɳ�S)�i�aR�5�İ�jd�Q�e��u�ֶ�����p�%\�9L��%��9��Xǧik�©�6�!,�K.
F�md��ITT�ra��Br\���/'��]�iߒ������ M���x���7K,1+�e w�Pq.F�(�>�Xe��p�ku�j>��T�S�/!�=�0�q�]u�m��4Ҳ�/Ϸ'$�zRIc[�*��B��PJ��� �S��a��.}*3/�]7Eр<t�=�8����*\2�¡�x�����cufa��!Pٙ�LB���F�APQnCу��Ui�Ffvv.l�61��0P{�fY�h��� r/Pb��Rb!#l��p��U47�r�f�\�C�~
�İ�¢$ļ�訜2!C3f�+뺻љ�Q>'�٣!{����x�P�r\��|h��჆:&�a����:p�f�Ԅ'�˟?g{j��B�^��>��.��)�8�dh6r>���a��|�]�/1EɓRh�ٻŖ7J�%�t�X)0��gRʮlU������Oqv���a����V���=|e��0���N��u�^J�a�d��C�V��bL�=�����Sq��m���V>~�o�8�/���'�F_�u��e�t���Μf�<xފ�n���j�!�{7�%��� �~�.H�e���!�!�s��p���w�2�r�o1�KD�YlE�7Lk ۆ�����^Č(�6T���Ѭ0�����)���b�����#0�c=hj�}�p��`%�&����d:0�ܩA�ѕ�*��&C�r0k�s��ٺ�;�����I�G�S����ܙ�Ox�N��.2ۮ6�2�F�V_<q���0��jO�
�%�+Ta�J�u��!�Xō�V��8� �r�yI��qЛQ�s0cp�ÈmV���a2wb9��C5/+(�LTZ U㉸��P�����m��m	�����^u��{�wI�e�g#�n���6���,63S��Q��hѳ|��W+�vl4emV<�,��f5:�%��a�&��Y�Ѹv&!F�f��0�$�׼�TT4|��~��Y��̶04�j2�l0����r`ف�)p�fK�f��
P{�q-�n��g8s�wq�:vz��}���z�s�z�/щ�m���2ێ��2�F�V_<q����SiK�tj#�H��w��m�ڤ٭������g!��C��x�ZJ�	�`P�'O����(������C��)UEQ���h�7�!�je\�зG�l;5� ��d<w�e��e�mq�,���%|x���rd���������g����ٰ���L��f6�)��W����4�.U�er�6�JⶳN���8�]���یJ��	�a׉�l�HL&V�+��Ex|>����H�?�W�>2W���~	�xO+��u]*x���^4&��h�'�dx���a�&	�t�&U�°�MVk	�I��0��
�&c�Eb/���j��c���C��|���_��آ|(υ��W�⸹W+�\�e�'��D�<C�ч��l����jaf��VSF�a8aXL�R$�a�(�p��D�_R�x*��D�p���#�D��C�<8�
�<Q�	�!�{��쟄_���=֯�����k���qi����޾��v��P���M�w�����k��V���ݝ���.Y��LZ�3=g�}����#�w����^^Ȍo|��N�ܚ��|Vl{<���g�yi3ML���Y��&ѭvUu'}�_nkZ����᯽�r�~����_s3��9ww��335����i\�.�33J��i[�]�ffc�Uⴭ�.�36t�ÇN�t�&a��Ä>6YE�##�yUUH��h4n��?|�b�����<�-�s��]�ڤ��7%%����&BC�&�>��0�th��Y��s�n�̬�&%�L�n�k ^b[.A[��5����]�ԛ p%ey��X���s�F�4Q��_n���p,���$#  ��f��a��a�b�c�Ө�l�M{K�n<z�m�^=m�_2Ӯ6�2�C�|l��$��F-�u��UUB���u�TL��a�����:FY�4�ɓ�%>���n�Y�Ul�#����H��D�#��2�o����P��k�7[�w�b��%i�a�r��i�ٶߔ����"78j���ȹF��z���A:gŬ��(�>�@���x���|�9�����=�5TqS&��$��ק8���z㯙i�[q�q�M*����o��	�j�1�\\-�Ǘ*�q_ڿj�uD��W��$̱�J��X�pH�� �kW+�J��U4��	ښřy%jE
ݵ����W�2Q:�%emX쑊�����(Ԫ��s���m�%pƵ�����Z��@��}�1�b:��b�s�~����;.Yf��w諾���=Zs��~,���:o�Ȣhџ�a�̇�h��G�xrѱ�WUmV�2�NOA0fg&9=,�}4�[*Y�bP�e��T؂-V�]�CeZ6��p��$%ѳ�n��ӡ�>�Ba��s�����/�ϡ��q�]e�i�q�6ڲ���.q�vMk���@�'����M��n�H���Qi�n%C�32rP�b��)0r�
2ˮn�hbZ6!�夫�I��&����i��^�wv;lr)c�8�Ӫ�AX�U��Veh�y?WM�g�i:C�Q�]s�D����|`��Ѧ3���|0����mZ��9�|����i��q�0��"C��ߧڕ�ֹ�p��+�ܸc�wY/���@�I�!ܕ0d�C>j��fM�>3�)�&�����������\<ϱU��O�v����0y��^�i4Xy6}�˴��南tQp�ύ�0v�6U�G�F�W+�z�\n��v�t�c6���=;��<|��m37ɩ����|,r
غ:`�7ŷN��L��m�*ڸe�|�-8�N8�8ٶէ�b��	�.\H[�.K˱'�uUUH�r˚��\SF5��ɸ���Ѻٰ�{�6?��!.�����c�VZb]°��M���*.`�B�ʃ�pM�G{|!gƍ� m��9c3CPJo"��Q�B�����P���%͜�J�Ę�\.hNgF�d+��l� ���ԯ��kU�����,��8p�0�~0�<`�$<pѲ�NR����J���,�,r��.\��!������!�-t.8I��ME����I-u"alr�&�G�3 �g ���r:�N^[̰��
]��m���6٭HA��E�)'���
Bۢ�Ç���oG~>,�>�0>���P�X�
��2N�<��ơώp�!�t��J;�u,��E�`��N�2t�Q,O��j���d��fr+,��Qf!�
��1�FDҥs�mOv�u
	XŅ�F,���Ov��;�?Q�@�6�U�^�?V�����\u��pL0� �4[��Yu͎���4}�Y�m�>��~{�*���;*�cC'�L���Qp�pF�����	F�4i�������щ����.1��㑦���#�ns��|���,�&��K�a�(D��h��E����!�]]�HF|ڭ֌=G�4�.B�pĹ�Ô4a0X���0뱉y��W����{3�����^?��0����F������wT��LΪ���j�\�<p���[K���O�&$�
�"72k���,Ț0Q�~0��{��X��A�b�<rJ���MSeU�۶�Y�R9Wr։g�G�6C�Ȉ��:k:X�b���Dd�6�c�;���r"\�QS
�<VU����c.?�]q��ˮ���x���ْ���`�#Ƭ�]�nL�Z�h�R6�h�;<���Cc(�K�IET��6`��CN���3ا���
�ZM�PhKJ.[ee��"
�S���m�����!�p���P��j�e��!ύM������j̉p;'�85.n͉M�w���Y�Q5����Ȝ�B�Y�Q˥���tnf@�.l��%��y0d�>�#�0>��:�/U�u�m��6�d0J�$0�aBaf�J�)'���q��.8�|��1�i~W�aEa0�,�!��0�C�&$8a_a9&l!��l�l���L(�XCf��x�&��$�%Q�K�	�������k_�Ҿ����'�G�d�4xRxؘO�c�ʔ��G�ҩ�Q\Z�*���e�?+���r�Y�ix�-0�u������8�Һ'��m|_���x�\)�3S
0�����0��eI��=��K�&F����3�S�O
(��D��[(��˒�<4xL��x�_q}2׽���]�����}Bfh��;�n��(�3��[�a ���o��NOnn��T�Cw"oeǙs3dKVD�Zy�j�+o�C7�u|[s}�G�f.���{G;��^�϶{9�U�������{��4��RW�f֯SZ��������Xw�|}�e�V���yl����fu��OT���7&���E����svTz.�7���j��ܐV��Sf}�f��e �[�ٟ[��A��V�`юU�՘���c�j�ޘg�{���,��5+L��N�"�.�ͭ?u1oޑY�|���x	핸�f�L]�3�>3���mY:���,QM��N�=�WtS*��D�:�ڽ���>��+z<��v,��S&����n+��j��י��n@۟]����jMK
�>���ʂ���5�Ϧ��ɑ�7�E����5}۝;��{^��7_	4Y�4�<��,�K֧v
����3����e}�͓o{�x /O���덾�YQ�n�Ng�>�\��'y[�U%ꟾ�)�Y+�e�V9�D�"�b��,�[m4�
�r�թ�Q�J� q6ꜜlL�i�b���EYSo��q
؆헹�5S�N��vÅA��kC��DD]R�BjY)]�־x�4@�L쯹�>_��|2cK-u�(�v=g90m6"8�QL�VPR;QThjZ�m���2Q6^4X�5`��)��/�9��y�+J��.�331Ҫ�ZV�w����UmZV�.�333������]�g,�ÆΝ:t��/!ub�-7�&�oř1[&KD�x�����fUD����a�n�n�3mגbT7�TȞ���a��Im���Ss%"o(卹_.��e�#�^]�U�y�I����j��9A"�X��GZ�W�%��͝E�6b"'�����JJN�I�P�dL�|�"'/M��4uY��"�p��B��bx����~0t�à��d�,�.L!,�5B���se�E0[�i2X�"	aR�X��Ss��f-ݥcV'X�r2�	��8��X�.F*n�����I4Y����0�Ɗ��F�Z����Bp��x�㧎�<p�p��o���0��U��'H¡�*�<jbT�g���b&9{���d�nd���;��z��ܓ4C(蛯��f�{��M�� �H�/��}F��Ûh�Q��3�6t�Y�"'��˶�M+KwKb���Z�j�6YcZ:j��G�Qf�
��.փ�a�"zY�bX��C�b0��?OJ;3���ŝ0��0L0L<x<x�K5�����0Ř�˚�*������VC�m%4؉�>�11phL0�4Ud��>8"���bdM¥7��e�0ȉ߭��KJmS���0�e3�Vk%������j��3"Q�7��)Z��&��F5�L�U�Pɡ(��_���f�P��O������-��UR�n+�Zq�Zq��u�iƚ4Ҳ��|���1���b�%�n�UZH4J%�	TV'"�;��*hȜ���wj��1���6}�:&�{բ�V�,m̷�8^bbfY*�nEzQ�ǺxDK�R���J�髆 ���򺃃'q,�9�;�b(�!v�oҎH���%�L��Z��v\�z�����F��f� �'0�,O�B�M�B\�⣃M¡���}c�$¶�Ӎ8�m�ێ4���yy�U�_�gŮ�mZ�3u<k>�˕��"���#�B��ܘ�[+F)+c�*h�f;��i�cuU`GȧE+�']cQ�I��i�('P�Ӫ.��'y$��9r-�\ꪫI��l�阱3Y1�1c�Sf�(���%�2�V�D5U�.��j�!l�R����U�PįYBl1>ga�ϳ�;�ٳj�f`j�:�������76+�/%���[4Y�ǫ���r�K5TQE�:[�i.��^��1�5�m����UVj��8Y�(HCg
���L����y��5a�Ɯ|㯟:�n8ێ4�Mi�d�Iz�j^�f��*��B},��鲫|K�٨��cp�f�b&�������~��IIpɶQ�;;<Y[����`6Q�p��82̉���Q_&-���`�.T,�[���,qR?�]̩��D8vå�D�p�I-sa;7(�SУ�7��%���6�L����֤���6�n��n6�6ӁÂl�fxE�}u&XwW���ܩU��UUi!_Ha�G��}50hM��V���!�\�|t����%J�����f��[�pP����qJ��o��}]�Kd-m��V�������!�v��A�P�G�:Y�|s}�B}d>�.�fק�s'�ƚ�t���7p�bjs��!�f�SX���{�Nx��*[*5<i��S���2l�N���r�i�q�m��4Ҳ���j�;UUi!�I���5_��|˫����||vN�����7:&������\v���uû�kt��Z�tx���8;�(D�����%|*"��βP�R
�
��.|�bnk�]~.��lMK r��/3f%��=;21,M�Vl����"�p��I�`K����%�8|dӬ��n6㍴�F�V_<m����;��Z�M�j�;ϵnq�mZ�[32c�A�<�y��US�Li���调���#���W�-uYS���u,��*�NF->UUi!����%Ƥ���~���Y��%|fy\ގk�CE�U������<W�a�9+�pR�ps;**z�)L�}(�jfg������D����54oD��`L�:&Q�w��!��h�4K ���}���A4�r�:A�4W��*�+�	.vT1
2N�lF1��;�k.�����Ĵ��d���[i��q�m��iZa�����%ʓP�Uܻ�fGj��$;B�g~�(��r�j���viX-h7��[6g�8�&���ۺw�Bl�V.o�CR��K��j	�R���0��f~ڻ��thHwD���k���������s�[=|���bfi��F�s���q��.q*��h��vhN
�s�
LoFĨ�QLH#^�Ƀ��	���	�'�	�<'�O<'��<lB�DЈ�H��B�DЖ%���,�,DؚblК �D؈���H"&�D���<',M��BY��6&ġ(����	 ��6a��a�0�6&�(Cǌ0цa��� ����<x�bY��AC�	DțBlD�����}��~��J�:�^��놛g�h�=�ǏfN��������3�=}��~�h��]vN���}��_�L�ilz#q=�m�3��kj�߱f�l��{���VDL�sz~���������z�#�{�����}6,��)b�p3�����y�RWs�;����r�t�y˼���v�ڮ����3333j���n�.�333Uڮ����3.Μ8p�ӇL0��q�Zi�i�_<_�J����1�b����X���B'�!�Bo@�A97���_
�V��''j�鹳P�!�?�y����s;4'N��O�c�fE���E&<���$s�0(L�\;�"���Ǯz��/�5,��z��wĿ�`��]j�:{����4�ڽ{+
����{Gq�޶���u�m��iZa��9���2���\���I�UZHXʜ9��Q�b�Y>��W�����B���9�j�_x��M�U�i��c%.\�/�]��FU~�� ���X���]Se[C%�q�C2N�ϵ�J�9��KMkECCFOO�F��*�bg}
�fT=>��:l��>�0&��?��jZdK�����{=d�uYm�]|�N:ۏ6p���e�I�w<}1�n�TVZ��Q*E+'#|9ES%N���A��㼶Z��%��Ep�Z՘3��Yvr'%�2*@���2��pc�ІW��a`�[�,�uUU����Iq�e��.K��H�e�Q����M[;�5�6CT~=^'*��93>H���0�3e�?Jq����Zj��u�|NM~���^b�n��N�Y�3�rZԚM|"+�f`�&#;���7U�Q��2u��M|�%o"��:$+KI*��F앜 ����߹
���Z}	�Pt���'|f(�n���N8�n8��iZa���!9�iq�D�]�s�ꪫIQF���fN<>��.<��(Lұ�3�|���j_�fɸQ�7w�$��@��Ѐ��8����Ŝ{�6`MH7+�l��20���������%Y�����O�o�Ḵ�0�-��d�YW$6J?Q���W����ڱ(�36"xaRQ����k�]�]�٢c�G��:~8p��n��n8��iZa��1�����.+]��`�Ѭ+!��*��Brh�>�Mnx��ѓG�S2�,~e�(M�� ��YX�w,L�C��Ul�;�%�����]��An˫n����:}�5����مR�;�aV>����U�r2���&�Gr�t_ʩBbJ9�X|j�S�l�?QfQ��%a�::�Ϟ���q�m�M4�0����=�I3��I*��FQ�2���9�<pɌ��9b{WU欀��9�NYl9V�O�B�Y�j��/"&a����1s'���t�#��󭲮O�#���������.	˘,�6�o�ơY�F���q�x�cGM�_��U��ǩO�T�UU��hJ��_��f�yV�e�]|�N:ێ6���W�]Z�j$.��X�׷�I����L�jH��<��B�Bc�2�	�͙���ۘ����%�˙#�)��Z�u44GT�"*���d@���Y
�*������EQ&��fBVSq�jqUU���GQ���+�#i�+�M��ك��]I��/
6��YF�e�'ۆ�pɧeU*���{�/Y�ȝ��p���O�hN,���aL;r�O�\w7sSPޥ=���7�b�ᣄ�f��`��9
���y�B��_?��-t)"%�W%fLLU��Q�Y�ɳ%���LT�`�9
�C�a��X��P��,��m��6ۭ��m>i�i�_<s_N�w�G�s���$>{R�����4&��*���6?`�.}*}P�	����؈y1
�r>r|�^��ݵpﱬ3lG�S���{T��`�P��t�uF*��uH���/H�bn���W�8������&�bs�O��+�4B�$��k%A'��:<,K:�O11Bg0��6�o�q�[q��z�J���7#H�A�9�mUU��j�ل�/�����U��=���Ƴ��'~A�����O�F0��5)_5)����=4%�y�p�d�q>7�+en�Z��m�akt���77D7,����S�j���-Ι�:`Nkʨ�	�dM���ȉ=�Z���{UN���11<\��u
��6hٳ�|㭺ێ6�֚V�e�Ǚ�/<�� ��r�RV��
�Z��ڪ�BT?���t}[��B5˼^C���?|�A���,�"�����R�K˱�Kb�Yd���\%r��,N�>_P�Lό����6�ȟH�1,��Jp�ǆq�YG��k4P��Mƨ���YBfr;�3g	�J���3\�R�e��0x��i����_�~e�e֛xO	�<'����DO��"A6��:hA�6"xO"'�6&�؛4&� ����'MlD�"l��'�D��%��6&��BQ9'�!�|��BxzNN�a�Řlن�!�hD�0L<Q���b"pM	��xK� � �"%	BlM����z�7��!^��J�ΚXy�qU[M��#��w�Q���ovj=�η\&��n�"��)���9�9ᯛ��aT�If����oN��J֫_�?nX����\����:Ț��%4���^���[6�<Ƚ�c�$Fc �VA�s.�L1�e�I�p��}�[��֕$�6=�M�����b��c�I*��?��b�aݢ�rNNZ�,a~��7I�߭�c�sgۇW�w|���̎�H�b�i3��;����:4nܴ���|�}s��j%D;��-�a��w2�9LV�+��B`��c�gٚf�Z���Io'w��5�$��=�rX���*��w��J9~��s�o������._��?�� ����g=����-U~R̲t��{�n�m��qŲw-�dΞ��k��g�܈�ߞkMe����y"�NM�J䜤/)Q������4ݭRIU`Ꜯ���rXrT�r�1EA�<bt]h�ԣ�����PW�fwd����cl���|�����cC�S��K%�Z�;c�(c�V�tmֱEn6�?77�d�j�l�u��ܬG#u��,���V�dÁ��)�{����byT�q;�T��	c#��p޷N�~��v���^fffcj�Uv����fffe��U�ww��������Wm��^fnΜ8p�ӆa�a�x�Ä8'�˯v*Mݑ���d�6	���jt|v�iѶʆJ�F!;P�El�S���Uj��]EC
Z�8[D9�Ydn8!���	�[�����l�8�H�TBmF��Q4Ў m-��wͶ�o��`����v��X��`RI��3�6&�U�Xͅ\(��P��P�U4z�`��٨~XB�%:��"�Z�+����

.���E�	��RQi$><p�{z���~����YNSU���p�:YAf�/�7���S-��VV��ΰ��M8�m�6㍲���/&��E ����B
�:�mV�,�>�̢P@�s������7(��7
����j�@OMM�4�Ç!F[6M�j�Ųel��>qC��P%���-1�n��Deʈ\���"�l0�^��w�W2�W��e���ag�ᇒ"�x�V���]c�q��e�x���!⎜4{=#u�[ѭJ����UUZ�Wpk++�J��)��z�WS�^��2�)�&����"4�J�9O�̘@���T^��uw-��d-cFV�j�T���֘���Yܭ�xѷ�Ϙ~��Ѡ��s�ʱK��B��j���>z��d�Q�:�up�rϜ2�m8��'�0�:l��(��Em5$ԭ&cE�r��2e�c$ͪ����E�ڡGIUZ�=�K3�C�F�,���&K�Kqpb8ˎKV*���V��u���`p���,]��
/ĳ�\<ljxٰJ�Ql�����f%�3H�M4���,c����2]�v�E��VCd�2�?��,�4~%Ty%z�-6�,��M��l�i�i�V���y���X�e��	Yˎ�	�F&ڭ��Z�*��ǋsJ�4k��f����8���q�Rȣll��cj�l�U��0b�Gr�r�/)*��J�c�^UUhGxoyl�.
�0�s
�SE*(��sB�ý�����8Y�Ĳ����A��0d&��{�!���mѧ#����[q}��L�*�������9;kmJWA,�e��̆J�uU�-��jo{��,�̂zkb���Z��"90h��u�[m��q�^4Ҵ�/�<y��!Z�zUUhO������	Hz�5_R4Y��ь�y��Kk�4ar�M�}IE��$�MÓ��<��`����kgK�{2���X����C2�%�e2M�G�TJ,>:w�?.}e�|}^�J!>.�n\�K�_��(�L�>���P�6x��i�[i�\m��4�0���o�U#y.�}�UV�Ĝ�f�Odq��>����\�T�Ua�����d6g
�:�bQ[��}g� �d$��δr����[d��U0�q�q���Og�q�~o3@���0�)�ѣ�^C&<bbc]JLʇ����pӬ��ǯZm�e��|�L��M��l�p�	����d̵O��UV��U�]��jԫm��3s�Q�/8
={�h� �㏒�l���GF!�.�����i�n�ƞO�}��p�+`ǸW'�(�\����S'�tv�a���G������gU�ˊ��Й�/G8n����d�����y��wT���+'�rx(�;bh��̳�~u�2�m6㍲񦕦|��?>F��B>;l��}��w�J]���Z��i�:n�۷q؎fZi۳d���o!�`To�'U�V���r��윎WyD�$U��A�T��
�H��q�ş�m��T��G$�i��-n�8�%*[�1D�_,��U}�[.���0�6�7�E�̅5�U,�����E� t��3f'9���,���&��h��ll;8lѾNbt�Ygð�h靆�ì�~�@��l���ZIwr�Z�۲�hj��5+g�1%�u�Y��ҧS�lӋW,bu�.4��Ze��m�eg	�4'���(¢�]7$��ʪ�	�%H`���9G��Q�s���2oЮ}�|�8�϶�TV�+0�ɳ�pgRd2bC������g�wG*��
�]��	��n~��R�� G:�Q��u�(���������S��Up�)��f�&��H%oGM�M�Ǌ��HT�#^E�~��km>~|�:˭2�-��<'D�<l�8P��:'���Љb"tDJ�pM��6t١4A���҄ �,Љ��y��X�f�4����8l��r|�(�|��Bx؝����0��0�<a��DD�(C0�a�0��"x�e�f�AA�L�e�b#�SwT�����߼?d]��Mn<���a��{|�չu�_?�]����n�����N��0
x~~��Ok{�w9�|v�_{�Zu���&����u�s���O~�N�����:��U��S��:�����+����J��O�/vkNs�{�sJ�ۻ������x��V���333338��V���33333�*����ff�<t��ǌ:`���8C���2���Ѻ�te]OBj�e�F�|gk�0���=���O#[~Z�|�|�y7���.��O��x�ʈ�)o �9@�4�#�&��5,NR�Ӳ�W8���'Q��m
t�yL�4��l��XwJ�sWL��bo���<+%L���~�f;���q�̿8�m>:p����8pN�ѷ�UKO/׋��1�}�UV��r4e�����W�j�~�����y�*��t��T�b�2,J��Ɔg�O�=쨇����k���WA�ϖ{2C�MQ�5����37&(F7F�_Ux�j���uMx�Uo�F�vo�4�&�׶{/��o[��c�����q��m�[i�\m��4�CP���Q�	ʈ�"�"��YhD�F�'�[�ӡ3��6G-c+�׉�H�U�UVK,ܓ$ʘ���6asB����
��i�XBr@!�ՈW,�I�֪�x9T*���m���� U��J�#�j7�\�dF�����������g�΅F���0ٙ�fl*�uNJK�RU&ܥ��s��p[xb����14��14�g����$��m��g����1m�j�m�j8hA�TgI�*' fr�%�0�m���:�4ˍ�ێ6�Ǘ���CW|���~���"K"����ԸY�yUU�(�Tp� ���c����w]u���/#NM�{=3χ�3!ayʢ��>7K���/��V!(�j��"(�er�K]*�l��X���5r.�}�=��n���i����R�>��=y�պ�s��e��q֙m�N�:|x���mt6�˻wR�U�Rl���5{UUh�I	��b��(�b`���`-4��Ĳ�m���+���4�<��z��%�n�Q�Y�{��_��*��J��7:sc��V(���CD��ҎS��ʅ�v��m]p�I�l>�"z�����2_t(�J=��.x�x���kan+��ˬ�u�\mç�>,���ف�L�z�p��UZ=�]Y��s<E���ޅ�ϑN͑�+a�<*�Qj�̽��c~��~ݹ7[�f>�O���7�>���Z��1~�����c1���ڌ���F�͜�/����֦�~;[;�E���2�6~q�.�˭�ێ6�ƚV�ͿI�ޯ�׶��y��%��X�`�bۙq����7;�a�S��Y�"��V7�^�wem���,�D��nx���hu����UNH ����&E�~���m����H$��R����S.�����Ç'�!���ۆ<���$H�b��*�����h䩘d��õ�}�'F0(Ś�<��ʸ=5���1��؅�MZ�*�L�)��f[&Bڑ$ ���>�N��(Xd3<uYA�[}���ڛ���ξq�]m��?>�p~�c�;#����UZ>��T|l9}G�2"<�k�������u�٫�ޟ|{f6�m_}�Vv��vp�p�3�rkA�oڤ��X�kP�^��Iֳ��+��a�������LO^9m`oo�2�o��;��y97���j�-QG!و`Oz��]i��i��q�i�i���Ǐ�,��P�-y�F�'���ڭ9���tv��M|W���f�G��2S?*� }G�*��Pz�Gߤ�h8~���̄�F������ܖ���e��Ä�����by�HSZ��!�gi�\z����*攡���!��k��G������ԝ���S*�'��:�-��m6�N��4�1��_�	�4&=hj�%c�Q�ʤ�j���T�Z���-n6j���j�+���!���F-{������X����Yb�2a-cB���)�U,�arX�������j��=py>�Ylјr	�>�l>�j�����Ŝ0�Ի�6�O���|k�.�p������m����{<q�q��u�Zm��'���xDD��:YGDJ(D؈���(J �M�g�舉�8&��bY�f�D�"lDDO	҄ �� �<'����؛4"l�4%�4�T� ���AD�8lD�GD��0�	�0�,DD�(A��0��	�a�NY��(AADJF�M�f��M۾��nj�����ܪ��f��r'v���=�yy�LlE*���qkpvd�XDH�{�����b�]�$�Q�nE�Md2mW��1��V���潗'����we^�ov��\y[��LNrd�ztO��κ�|=s-��2��c��:��'I��ySM�:85�A��'�lb�s�䎣"w������"��dD�g��JϷ"�鲇���v��+�y�V����cR�ɕ�$[�]&��ɆcVff�9��p[��k����}�����kV���_,��L�g�U�[#+��c�qWd]왊��}�l��>s+��X��f�=�~���>����sm�1᷻o�X���ww����<�s��&���gV���hEb���Mk�����(۱�h��c�[�n�PڊB�e����iJ��INX(ԧ��qBư�1;�,�VFӭ� [L�8UR�5[D	8��mZ�أMV��Q�l�m��dQ!�7YV<`4�H�MR�,RB��(�Nƅ*"��2Bq�r�TȈ�VZD��mv�QW�㑢Vؤ�@E
~��:}�=����U[��������z���wwnfffffuiUn��������|�U���s3�:p���'�Ot���f����=�H�q���_hK��
�B�ER��c�Q�V�ǖ�l���EG5���]��VV�F�!]�B���ڥn��$*�&b+f�W�l����g�UZ5Z4>���H��hv��*rq��([L�=%N��&x?@���//��.�N��0s�C\ٰ��T�`�v{A�Y�Ύ�ߜ��+g& uダ�9�d9Cx5_"����|�ޢ	�0?k9���Fck3.�Ŋ���Yف5�M¦˜��3�u�*w��O���N,��6�m��m:ʴҴ����{�Դ�'9N~�Vl]���>gG�U��T�$pd瓗	��F��w�N2&^���e�}x��b���KR�0fjs���>�sl�h=[����ݐ-A\VJ��AțmvNB�EL�&�(g�2|_���h�#�f9Yjrl�����_�>{LF�u��m�\m��i�U���^9�4��9�U�gK7wv�M�k!���)�隙� ���)h��CKV�W�V��Ѱӱ�J6�LE��Q��#�*Ҍ4B�C���NB�>��wj�_a�Ү�e�� p2	��Q�����_�Vn�&��]�=�E�e�a�L/�������Ŏx��]i�[m��i�B���TZ�d���Q��� ��بƧa���R��d<iQ`�Wؗ����}���W�=�]i����s�!��B�*�ˋ�zw��Jv1�V�i���q��&�\G��V�8����
���C��%�d/�4`f!�
Ȋl��Ĝ���w�G�1��̴ӎ��-�xD�Hx�4pO]e*d�Ce4�
�$ʥ��MV��"ͅc�1AMl13)�d�Z�D���V�K9Zǘ����qY\i�Y\��]�fTf><E��r:�+�Ӕ3�<mX�,N���&YN[�]C�� ������)�`��&6��!�Z5s+�0�l��K�8Q��8 ��6�*�0��Պ�ѣsK���}��ɒ8M�(� ̂}5�.h1:j�ꖪ�{��GRdC���J�d�c���N118�TL��)o ��}ba��b�xq^:ˮ8�.6�m��*�J�/4͘���+J��V4`,�3A�9��&�ϙ��x��u��)^j�C���q��C@��9O�CP�ӂ������6s����n��x/G��2�Z,Y�`��r�p�a��R�F �Cu����z�1s��	������'&a���s
��"'��L̒���}!tlJ:'L�'���>,��о�=,�.de�j��Ua�����.@K�a�2>�9:C0Ƀa�c�e���3�k^=�4"�r�$p̧	3-^��d��dɃ �p�tX&����}�6L�8�|?Dɩ��䜅K�v�\y���R�Ic�]|���m6�.6�gN6'	�e�4��]���o��Q(�r�����2��%�{U�p8Q�A�ՠ�x�qb��T�{���JJ���>�ȅ����F��6vx��V��f���c]�T�!�3ʛ*��*���ļ��rL�#�>��M�k3P�(~����_z��%eٷn�_������M�a�	��'�:Cǈx飃�}a����G�0z>�Aed��#�s�D70��Ƞk��r�.�2��4�&�Ց�	*�!��eXd�<���ԧ I�Bs6o��o���V�����wsc�k���ua���/�`����0TѰ����߆�������|b���˸�z1���پ\Q���QLǨk�Q�M`˿+M82��Z��e���a���W4Dg��e̘e�]�mU�!F+���ɸt�Yl�d��)�}<|���8��\i�]i��u��m�V�V�x���Wx�Eb�Mj��K���/�UXb\�̙2Z����*���Ai���qe��|�y���"�5�e%j[ڡQ)J���&���������(&�_��uٲ�'rbYym��i��s�J��{2�Q�UW���҉$����;&�DL01AK+ꚗe�8Y�<x��:~�DO	�<'D����t��D(D؈���D�X��O��,M��͔h��DD��p�F�DnDG�X��p�blM�I(M	D�T���'�lAIcr%�h�d��a�""xN ��"%���m��q�W�=xÇ6l �M	�L��4X�=U�7|�q�rN��s	�>w���0����������z����Ft�\����J��|ߟg�|�|{���^��n�Wކ�W�w۹SS.�������Z#w�}��/#�־׽;���v�gn��ڼ��&�������.�q�{��v�wNom�]<ޞG��MVw}_��}��:�.�s.b���E�Sw�/��<�{w��\���7l�"/�;���)�il�+���:��w��o��������s3��W+�2��s�����3�U[���333331Un���33333<�U���\�����QUn���:YӇq�\m��i�V�x���m�?I��iT��驅��Ic�m�M͚���ta���*7h��s�8��S�,\;�E8&���U�BYH2;)�{B׽\���&�N�我2�E�! �;?>e�|l0H{�����M�f����7ɘj�*�rh>���~���4N�l����K��N��:t��Âp�f��y�[es���t��ep�Qvx�J����.��63��6�r�t7���V��HV[Qj�Ɗ��d��E���&���d��wcc�=�F�R�s�8Q~UD��0����K�7�׹e]��.�e�[uF�a�5G�
�N�1�]���4l6���u̴��o�:�-��m���M+L��D�W���1���S%�35�&��ch�PW��:e�]����䶒��p�n=��d��ǒ#��>�̓��d�;��mW�o��92f`�y%hv����DaX	��ڢ���[d�� qL�4JTТ�9$V�U�%�aA[�Tw�|�7ElÔA�&b��QU�0�1�+�0Y�e���LEʲ���9kbl�6K�����p�f	�b�Gg~U���jPoK�%�+!�R�J�q;�'o�q���@��j�#9Kykn@�T"��
���>��j�C3���4'L,��'DO�8`x�l�Q m��b6�����a��L��b𩸙��ѕ:`�<l1&�S�zw�MeE#0Xs�v3JN�&����9A�8YF2N�ߞ]�ڶ�t�weQp�.ʇt��Թ�nb���z�nL�����uSII\�e_M�+�-8�֜i�[i��l�p�l���u-Z���\��,�WܒI+��,h��Ռd"��B���re�(��̞>,�4=;	�5�I��e=�j0�;w���q�&]�cv�m��d�EMQ�:b��7.^�ق�6SZ�.������<�raɺQ�s#&p�9���!��1\QPQ6Y�jt�b:tɃ�L<tD������Gp�\P���M�1��b�t 9�����4j����f�8��.�X��bL�0��a"�0I_����\8�v?w����b1��y�2ڜ�m����6���
�K��}�"aþ�X�,��4�]�_����������7��El�ӭ6˭��-�i�e���7u��mǙ�ehk&�ws���+�Dh���&VJ(�0ȱ[�,m��E�Z�Yn���Z�lqVG-�h�����y5�'+S � T�jF��8%X,DE�q���E��ƶ�ؤZۊE�0����fb	���h���G+v���tx�*�tK=�1@�4��Γ�(���F�MhZ63�Cf�(ɢ�	���ɸ|fR���Tog�d�[�Υ2=.�ș�N���L��et�{K��Ջ?�^�m���m��m6�o��(]Z��sӗ�=��o�9rTX'�m��=6OqUU�CU�l*bw���|fl�<e�U�?U���'d�0e���l�'�Gܕ���FYq�l<|������co+��wUuv���B(�t�r��
��N?��!E�Ǉ�=
2���pf�LYgGA(����uewU�#ɝ�g|u㎴��e��m��4ʲ��|	]*��|���UVnsÉ��0I�E�10���x}鉰皭ç�tatB�S��z]dDn�藫��q�˕<�m��m�
�lZ���4b'L2c�&ɕ�@T��[����14���#�r0}�Ft���±��g�D�\䭔p4b��s�z㏟8ۚ�m6�niY|X#]XN��d尶�7Y(�o�$�3C��,�ڱ%W�W��� Fܒ1��a �Ȝd�F����q{��=�+ǭ;m�������������31��^��[>cߙM�F�~5��(�>��GkX}_�o��Lҩ%S�h��_v�]a���>'�<� �B$�B@��$�"�EK��g�ԛ��?�K�A��X���R�����%L�~a�{%0o�ͮ����#"��1�B���"1F �D`�*`�IeUT����TU,R�X��J���)eR����*X�����,�U�X����e,R�X����R�X��U*T��YUV,~�bR�,����ʱVUR�YIb�UU�YK�R�,����1��DF"F�YUVU*�R�*)V*��Db"F	"#Db%YUV**�U*�,U*���#� �DKB�K���Db"1$��)T�U%�UeR�UU���*�b�V*�b����T��*�b�*K)eU,R�ʊ�*�b�Rʪ��Qb�V*�b����**���������FDDdDDF�0DaHbJ���T�UUb�Qb�T���UJ�UP�F��Ȉ���ĂeR��U���UV**���"2"#D`��b �DFDD`�#""2*�J�T�J��J0D�"2#"2$"��A�YK*��U1R`UUU��D� Ȉ�A��0UV*�,U������J�T������U*�UX�1"#��A�UX��)UeEUT�H�DA�F"1#"#���$F"#��DB��(AdF��A�D`��b*��UUb���Rʃb"0DF"#D#�UYJU*�E�����DA��" ��#��Db"DF"$���YUV*�,�����Db"0DB�J��DF"#DbAb"1"#	���Db�H"1��D`��`��bA�#b1��đ�0A�0B1�b"0DF$"#""X��Ub�ʪQUTS���ȔTJ,IE!E��Ȣ�QbX%1I�E��RT�E$QdE%"QP�(�H��X��!EAE�Qd(��X����̖0��őBb�% �*
*B��,�ED������X,
((���EIE%%�!E�)�&��R(�QQ(�E
,E�*Qb(�QB�!E���E���QB��ą"�E�(�YJ0,�E���E����B�%�*T(�QRQB��F%1I�QX��P����E�
,QTYB�E�*�)�&,R��J��U,�R�%)E%��-��Ie%��K)JU,�)E)K)JU%��K)JX�R�*�JT���)T�R�e*R�*�)*�JU,��K%*�)T�RR�)JX�)e)K�,RR�)JYJR�)K)T�Ib����Y)T�J�R�%R�JR�*�JU,��U%�U,��Y)T��PȂ!wP�0 T�2 �"��X�R�K),��R�T�JR�J���),��Y)T�R�d�R�J��R�J���K%*�JU,��K�K%*�JU,���JJ�����R�)JX�)b��,��Y)T�R�d�R�Id�R�J�%*�R�e*��U,R�e*�)T�,RYJR�)K�YJ��,���E�T��e*��,�)b�K)T����JR�)E��)e
���YJ���,R�,�Qb�K)JX�Y)b�)T�JR���JR�*�R��J���,RUR��J����P�U,��T���e*�~Y�iT��K)�0yIJ,�R�X��R�)JK�,QJX�)b����K(�YJ���B�U,��eK)JK�)JYER�R��U,QJYJ�����e*�R���K)T�QT��E�K)�R� $`2�A��HHTX�X��X��E�E�,R�b��"�)T�E��B�%�K(�H�J��KX�b���U,�S�R,Qe,R�X�b��(�H���1C�`	Q�F 2���RYE(ZYE��R,��%�X��J��QE%��K),��,R�,RYEYERX��,QeK?b`��Ie)T�K�X��*�(��ꉈ�R�ZX����,�R�R,QeKT�X��U,RYE��UR�,��J�,R�X��%��Y*��,���K(�#�	 �"#F)e,UU�RrJKI�����9d���a�h�)��a�� ,�"E��DKj���ƻu���?i��x��g�o�=���������\�?����`�2t^M��7|A�rS]�R�j��x�󦎆�.����m\����E����g������J�����Qآ�����W�vߴ����Cܢ'�0vG��EP�*EI@���#��_��;O8��2�J�e�����?�@�A�F=���`)��U@v_������@0%i��4 �k�(?G�4)t�)�_$����RR}	����4-y�!�ט��D�!���K��$ ����:|%%�1^� �[� K%�)TQ*��D�@C���� +�
��
�����8�d��`Yh `:m�6�m�	WC������S��!�U$�ZUHB-$��$bĄ�
YDI1HI1La�BIiT��ZU
),w�a������l�z���U G��A����P,�Cs�?0�>_���	y��̰b��'��3b�v�">�&� v~���������9�~!�py�V��������� ����}�D? �0�{���Wb���4|��?��jx�n��:���%|�c����q�����@�=G����R���#��"�!>\��������ps����^7�b������{�:���&#]�	<�bIg����<@A����d\ zr�;�	IC�R���Qk*��5v��6��ܰ��X�,A6`I�	��U@i�׏}����v(Ѳ;eQT�-�@� =���w|T��`���������K$��yj	�>��h��N���A��$�zH?�����u@z��^�S�|_'֏�QT`|�AƏp~�~`l������A�	~�l�Uݠ$��!C�ٟ0� A�b�.3����Q ���C���=���R�r���X=fS<�q��n6ߏ0�QT#��L���TO2��A�?�C`�!���_xt���v�� Q����`w�{W"�����DO�W�l� ��tm@��dr�ɲ� �G��Z����)rY��P=�kx��$���((F���5����rE8P����