BZh91AY&SY&$��K߀pq���b� ����bF?                �^�Q��� �IT�H�P��HTU�U$$��R%6 Ԕ�B���F��R��M�ҕ&��hٽ�p���$��N��U����$TE�iMH�
I&��J���̨�!(�f��h��AR�T�U�ӝ  D
�W���pԄ C�T �:�l2uA�Z�m X*�
�Z�A�C�&���+c[0���ٳQ��U%J�R��\�I$!�
��P������*�ӥöZ;Zm�����Z����4NU(n�۬�[���Eu���i�Uٜ�v�U�S��uݼ�-��n�:�����k��JDC[j�@JQ/>����^��ɪ �n�� ��}�x�Q�7e,��^u���z4{��:m�S>��J����=Ǫ{�vP�"��s�@�F�Y�G@�ǥ �)C�i�UT#mXs�JU(y�_M��]����JP�m;��ޕ��hS���کzȕg/<��
z5���;���MJR}m�
_M����T]�UX�{�(�����S�!��E)QTTIR�J�ҔR�=ݟJQ_[a�����( t.}��W�V|{�}�ev�ށ%]�o*{�>����}�Ψzn�����D�P��}�z��P�����v�Aƞ��J���b�Rk-B�>��)@緗�(J�M��E�x��C�ƕ��>�J�{_��z�>��xOOw�i�y� PzY�/k��uٷ��eT����]ox�J�ި��b�u$�k,��JP 9}�kA������ǳ��g��zUgN��Ϯ��z �k��nz�μ 7�=�t \{��m�����B��H�N��Jk*�,7��})J �{s���W�hy�=�zP�g  m�,��-�n P7���l;��補���t\�@�(�J
�B�TAٍ��R����>�9�8P ƹ��5@�04;��a`H�M��  ��l���w. z��� �v�@�� �ڌ��F�E-4K4Sϥ
P ��_ B������^�� f�҆������
.���Р<z`ho�� 9� �0 g\*�RIF�#o>���@5� ݽ����s� m�u�oz
 w+  9�0T�G::4wn  ���@�   
    �S���D      S���(�      SɐRT�h      OM%%H`��C��b40�$�Dd��@ �  � �R��J���%6�zI��!����4z'��~�����y�'vIʗ���9R|�����>u�Ϸ���}�w;�>��-�'|}�7���� gY瞾?�"�@�'��"$�N�O�����Ղ�I Y?ǖ�m��R"$�'�(��$<�����������t��g콯�V+����1X�Y�1gb�Y�1^,�b�Y�&/��8�V,Ř�bɋ1X�.,��v�bɋ1f,��U��bɊ�b�Y1x��b�Y<Y�Ř�V/��8�V,Ř�V+b�d�bɋ1d�f,�b�ۓ�:V,Ř���8�b�f+�1X��sb�V,�f+bɋ1|\Y�b�f+Lc��bɋ1f,Ř�Y�1ۓ�'K1X��1f,œb�����f+b�gk�1gK&,Ř�LV1�Y�Ř�LY�&,Ŝ\V+b�bɋ1X�Ř��Ř�LY�1X�Y�8Ř�b�Y�1X�Y�1fE���Ř�Y1f+b���b�V+b����Y�;V+�1gk�ŝ,�b�X�b�ʬY�1f+�Ř�Y�1�qdŘ�b�V+b�^,Ř���X�b�Y1|Y�8��1X�b�j�f+b�Y��b�v�b�Y�&+�;c��ɊœdV,Ř�Y��b�Y�;Y1X�bɏ���1f+�1f+�1qX���Y�1f+Ř��1X�b�f+b�qf+�<V+�91f+��V,Ř�Y���,œb�Y�Ř�qɋ1X�Y��Y1f,Ř�,�qf+bɊŘ��1zY�;\V+ŝ�Ř�b���ұX�Y�Ř���œ�&+�Ř��1f,�b�V+bɋ1^1�8�V,��Y�Ř���b�V,��Y�&,��Y1S�'��b�b��HňŒ1b<R1H�#H�H�Hő��F,F,F(��F,�$�I%Y�$�$�������b�b�b�bĝ�1dLX���Y#H�#H�C#�#CH�##H�C#��I�$b����,�,F,�����%Q1H�#CLR1P��X�Q1d�Q1d�,F(b�b�b�$�$��&)*�����!��!�$b��'##X�##�Q1d�$�&*�I1Q1D�$�HŐŒqF)��F,��(���+C���C�Q1d�T�T�b�U1a1d��1d�Y#�X�Y#GkX�X��###LX�Y#*�b���$�#LQ1d�R1c��1b1d�Y�H�#H�Dń�#�ňŒI�!�	�&,F*F*I�	�	�&,1R��,&,F,��&,&(����&,&+ŉ1b8�F(���b�b�b�b�b��&,F,I�	�$x�b�b���*'�&,��HŒ1Q1PŐ�Hń�D�Œ1P�##H�LX�YX�bLQ1a<Y;Q1d:YX�XLY<XLRN,�b�b�b��&*�b��S#HŐ�H�d1b1b1b1I;V,��,I1H�$�������V##LX�R1I&,�1d�b�ő1P�T�R<YYRt�H�#�C1d���LY$���$b�t�F,&*I1PŒI���Ő������$ŒO$�*I1d�b�1HŃņ,$�ȓ$���Ș�I1R'J�1dŒIV$��Bb�1RI��b�qR1d1H�##�b�IVHŒI�(b�b�b��F*��RLRI�DŐ��$�T�Y,I���)��b�V,����b�ұX�LY�<\W��bɋ1d�ū&+�œLY2+�œLV,��V9&,��b�X�Y�&+��b����b�V,��V,��1�1d�b�V+����Y1]��bɊ��f,���b�X�Y��b���b�V,�S���Ɋ�b�Y1dŜc��&,b��eY��b�X�Y������b�^,�bɎ���V,��c�$�b�|W�ŝ+�Ř�W�1\V+�1X�b�V8�œ�1d�X�b�\V+NՊœ�;Y�ŝ,��Y1d�qf+ڱX�LV+dT�b�X�V,œq�1X�b�V,�����bɋ<V+�X��LWK1d�b�d��f,�TœLWK1X�Wj�b�Y1f,���Ubɋ&,�b�Y1U�1X�����&*b�z\V,���b�X�Y1d�b�X�����X�V+��N,��V,��V,œ�1d�b�^+1d��X���d�b�Y1X�,�qSbɋ&+x��+�œ��8�b�V,���ŕqX�b�X�Y�&8��œx�LV,�1�+ڱdŘ�V,��X��Ř�Y1m�b�V,�bɋ&,���Y1f+�b�X��9&,��v�Třt���;uܟ�NV}���yd����u3����В�"ͪ���ڋ4��$�zm�Ktl��2풔��z�eLO�1JB�Z��h'��ټGD8M��t2���)9��4
a]��p謓^���%^G.I��r6���*�@����4Ch�!���C������S3,���ÒLT����ݍr�<"2�:�=��m��4X�����j-h*��kf�QG/E���;{��$5/7D"7.�K�U�bW��p�op��m2N%T�dE˩#�70e���0�\yHG�Չ�XՙY��|��r)Hb'S�t�`�����n�Z~�\�`n!�j��%�Z2Ř��(��7t���]8ڕj*�d5%�Ӳc6�U,2�Gr�0`�Wl�Uk@��#%@��j�5Y7($���kܫN�Q1�Gr�nBU���`���wZ�}�,J��N���-e�h�*Ԥd�в�j��(�xo>���ϱ�2�S1�ɭ	p24��ZsrY�_]�ĒM_Φ��u�v��p�6a��b�[h褷!���5�fA��l��i����6beR��O3�M����*�\�̣Iyni0����x��|	6:��t-��@�6��sh-��<�r;�ȵ������5���PK��Zqw=LJ����$���W׳T�h��ɶ�˚��D]�5(]�ur�B��u��r�zYaD�̣{��ƶ���I�n@ۖN=35�$&7D٨썗��DZ�`3ycM�{��W�j�����[oP���tMИg2�D6n�X~�+�Ӌ]-�e5��Yl�1�wL�2�G��m�Ma���-����-Łnn,�[��F�C��K��Blו�ج��i�,�)�!�)Vd��Em�;�6#:BCK,Y8���pKY��-��l�ݷm�����d���aÍ�t͔[����Uc	�j�5�e4m���4�.�\����zi�����%����s#̕E��v��y����4�v���������-Em�f�J���D�Ș���Zm�c���-�T��м��7M�#�cI)j"J��3��(R�[b4�;.<�Ҋeni��q;�+�9{B�i� ��(��SI0ֻ��sU&��F��6�X��SIԈGr���m��ΚpP��i�2��R��V��h��-U�t�[��56ޭ��r�Z,^]ũH�5�r�D�L�|IsH����]m��e��6TTL�K��3f��Xj��
�u������OsФ��,Q�˸S���qS�2��6Tٍ�/kDY݊��3E&m�FV��0\b�_eF%^bՕr@��1���#Up���҂��ۉ*p�$���&]�rfZ�ZY��j�\�1���T��{�]E�0�<�E���qI�r�b��(=���װ��P���F�lP�B�R�j��+Q�Pll�X(d{siݚ��!I�Mj��a��<,Ff�H�3tF�d�&�Vm5W$�C��"*����O䲌�oV�lY��Sc'lm���0�}���S`�3S���QZ�b�M�i�P�Z����h#�����ڐfFi��Xx����_�t.�;�ȊB���i匊�H�wce��!%Cr�ٚ�b��xcr�����yDZ�"�̴����Y���T��T��7�:V�L�J��w�ZeX��!K<����̺��n��	�3.��۬)�@]n���b�ƈ"ܙ�-۬�F&��Mn���V�q:�TPʠ�qhu�V)�xFeC�J�{D�m�ue���0BFcz*�0o#��k*iԫ�`�/)iX!A�+��gLq��2kn����Z���uq'Ge^˄�a���1�EV�W�,Yj��6∬��۹��B�^�5]�.e�Tb�7n�h�/%�b��[�g&c��(�n�Sl*���,Ce*�r\�2�C%]Pcy<��6�``ܥ�jV�]�/~ٓd���B�q��W�-���4J�yH4�3�i���ͧ��XfÀ��h�l�:�̓c`��%�V%u��6��,e�.嵑��Z�P���e���UR��N�7�`�s
=Y�%�ǖ���*M5P��-g^cDIn��hb�ۙ:��9T	CIM��=L�`�sUسrU�DB�T�����'�`i*,�*�!�۰eF7[�[�)#�һ��\�.�\��pR���2�P(%m�*���
n��o	2ҙz��0��٭�V-���c:7q�[kTl6���/6�c��6%cE��R ��f��H�]J��p�XȽ���h�-+��Ҕ`�ֱM�t�/jU9[W���76��W��'N�i�~�^\�L�&ke�����'�"*�"�P;�2I��6�朲�A��*g�-	$�t+�'�2d�����
�t�NY�抅�niz��k.`Ko)B�?Z��m�a�fx��e@�
cͳ����UV�����\+dH�v�Ĭ���e�Gb�������5`Ȉ�Z�Aa7�6�,�ķ�:S�{Y����@�i&(�5�[A�A�2셗���)���%T��=#��&#ǂ�0T4݆�hڼ7Na�L�]�¨֜%KRX��h���U+C �I�Lf���F8kon nź�(�a���m	j��sT�W�-VfԷ����ɛm\�K��\�v�ʕ�"X�Lx�ىjN�Zs$5<��C��(Ul��JТGr��pǮv&���=��L��:RjڱX3F��Uv�Ѷ���u�a�*���e��l)Y,V,`Q�nJx�奖��kn"5����0�5�ϊ�f��Nͻ�J�7aPa�J
a�5Ol�����[YOkt�c��m�LcZ��͛n�w
-�\F����[�.�n���xF�Y+m�����W3V���^+$�sK��
��$^:�w$܄�nm���ya�� �e3��.�X��r5m=L��o&B�Y}�p�[��{YO}�η@�R�,@�	Y�����B�-0օt]ʹ�ķK�� �ĵW0��VFKu!z
�F��`�R��ݶ*�)f�2΢�Ky�.�4ZƜ��(��d�ou9I�yl1��Xn�Hi���r��]Q��Z+\*�c�j��TYf��/���emKV����b�n�:��T)	��(Jm�խ�lV��.\v�e��Cv�^�K7H)�nQ����7*:ɖ�ѻ7,�Tw�,�(LF��Wia�3b�T8�6)f�Ui�R�N�AP���'�ikcZ���6����{D鐤� qt�wm*%��0f�T�n��V�͞v �t�@��$;z�E�Φ��خ�:E��^z&���CY�ݼM��y�f�nH����ۺ���T�,�i�fm�v�ء	��
B-IG5ɢ�rk�2����+%VwpM[
�o��KIл�wG1cx¬��{0ɂ��v�ȕ��]���Ō���U�	Gp�i��pP�S(�u����XVř��V�
��o`�l�u�@��ł�dm�LxuL]��UJ[u��Ȍ'��[�Ud���	��P���0RO�(fdBԮ���]��u���:����Hե 60/&f�O\&�~ѣC�.��r7p�aT�"i:
td�A����Y���n�Zm:�l[�4C����7O04h���[W��w��͌]0�hiZ�!f���۵k �~%�)ˇN�ůoi���V�[oh��܁j��V�EԻQe�v�]Ӽe��z$��X�Wn��L�ųV��[X-p��B071��YwA^��E!)a!S�e�'�w%�M\��h[b´۰&�r�]h��h�퓬����m�G-GE�e4X�(X�ͪ����DEnQ4b{�h/f�bX�3�M�n�	�;�4eB�Z��;I᭠V�Cc0}-�y4�S��!�]L�{��$�Ux�V����r���(iA����["l��b�3ZB�+ˑ�w�$
T(hY��b7�eY���e�v@vߑ~�yLk%��թ�zY�U�ְB3^�l��:V��V�+I��2�%��$;M��B'�a�"x�ؠRh�3%3��"���cR�U���&����C�f9@'��Y�:wU-�mH/fP�d�;f<�52ʦ�&��c�̙���a�z��C210���B�(Ki��P�+�;zr7rv�(�,�KiLēw���`�8�:Yv��Q�>Sqjxd��m�£�"�	luDJz�@��Q!�w��ov��EME��ύ��z��B3Y&-�Z���܆�l�FdI+p,E��V����;ԛ����h׭�ݭ�f	J�m�wdLn[�TL�ƃ�[^��.k���W�VmY)MYaT���yb�ߘ�j�#PX�^�O놅=����f�e�a9/vm�e��&�[.�Qa��	Z�:�i[W.��E���6��c��,��UҧB���Ȣ�Yө�V���jf�2��dԃ۪�sJV�F�V9�[�释�`�F5�lf���e)^J��W0��5yE�n�mAJ��Ov��[G-��0�ʦ���sTy�)'B�F��d1U�F�T�2�����vm���UYP��f�E�p<��qL��+)^��a���9|���Mq�Ye;fE�ζ�1�ZФm����X�?V�7@˻Յ��o5�8qm*��:n	��
q�Of8&S����R��+sLe̬.�V��%�cMS�&p�%��h�%X!�j��h��p(R�hǨ��"F�s1��ݭ�@��VJL�Ԉ�k緶X2`jf�c$�bj��D̺�Ԭ�X��(��\�F�����;�u�5$zHц-k��W�ȁZ.�&JA�iД�_��Ot%2e"m.��0=H6�K4V��VVդ�I�yL�$z/KS4N�(ű�hVتt�%4�czQ����[�� �kQ���oNEY�ח{&��6H���äeDh�5�9��v����z#�G[Պ%���)zVꃻ�����ᙄ�r�!�Fm��T��HձN��+T��6�n�nzo1襔�ORD�J�%v4��Ih3�t�U��n���CI�죰"�UIyeBp�����T�J7��9�)�$�B�Rw^�V�����I��!k��v-���짜.'�Yv��[���2���6wua9I|wn�N��#"�e��n�(Z�Uw`<�З���N��ZY�9nU�N,E)b�i{.�c̎\�̖@��dnVO�ˆ���fk�ָ�(�s@��^�Pe�wc4[WokSTӸ����Q��?JͼY��P�wb��F"���IEo��`�]�i��CM�k��_9�Y�=��Y�;M�Eg���ԅ+ݻ����(5�X1��t�7���؈�E�Z��A|za���lц�w���)��MO2�2�9l���f�mK��a�xl'y�\��=��v,"���c�{RS˕��b��q��9�d������K|�ݮ���ٶ;#Ñ�T�924�
�%���M�I���V���ǅI6��^�"��iB��j}O��E�W4��B�wk�vm�:D�jl�o���[f�������]�U;��紪U�xp�~UUۼ9y{��z7f��(e�yr1��q�/�ym̿@K�Gof��-/�4 ��"_jP�m����f��#�"�>Wa���%��4�P�E	4�*�}��s{�[a����ǣ���+w���~��wx�6.w�6YC�׋`K�5��KV�{Gv�u�u���N��L��Z����E_U�;W��=��j�E�մ�̏�'6�a3�w*�}q�/���ƚ�T�|��t	G/QJɱ�G6.�����i��#�T��>���݉KnP���+u^����a؇f�x(lK3}쏷�pDnH��/-s����0W:�%`����Z�vZ�V���7�9�ke�e�y�Q�#�I�E�4a?�h��OϿ+�Ƣ�k�r�_�{p|�,�	I]x��ŗ�_C�y�Oc�Ĭ`�R}}P_KS#�N�d|��FC7yh�vW]�;�'F�9)�ϒ�ʊP=Q�1b�NS)��K.�\�m��L�^!�:�X�=��r.ĳ���SdY��L�u&ڲ��b��t�Dp�o/sRAw�s�-;�k���<Yc��.�!��7���6n�X���b�	�@��q�JL�ئ�{$�V%}{2g���ḿ�����EnԼK.�\4�+ר�F�[W�{�4�&�����z�u��8QQS�^w�Ä>��J�Y.պ_1�R#�Ǒ㹑u��P�'$�4=v���V���l��ug l�2��~W#UGi��C���H���*�~D����h��,�]Yd\�VW��v׌gB)�>K�ӕ륤Xڃ���G�K�x-���`�a=⨉�zo�!�n�!f�̻�t�Q�#N֞Q�^����e<���JT,�����v���:Ow�`O���r�iJ����q������±�{`���!�S�6f�Hr�2ߕ�|���c����5'�2�#�ex�+֠�l_���m�~��+��i�54����H���扈��y���ݤRE�h�|�$EP\6sN*T��Qq,��]v۹��j�6�a!R�ܮq��=�p�`��,)E�pb�.�m�K&kz�vZ�e��K��[��6������*� yi�tkD�޻���m�EGBr���yud����`犏>�2�eS#��Z>��Va׆3Π�]�Ό��ĹW���ۮ����Vj@�w���*�hA)��lf�u�N
"�/h�J�a���f�޻�F-��P`�,�I!��fl�.#��U�%MҶ�7�K�+7���Z�6�g��ubBl��̼?�=z���}:��3B�*�>�&1dt�Ck4�q�by�d�����zy9����u3�C�₭�2�ξ���U��Nʪ�#E�mbD�^<��ŏj���6����ԥQ�G{y �uc;�1+Hd����Mc.��,�=��q��NF�6�����7��Y��vQ徍��� of��[���ZR�Cʉ�k��֙8�/�������c�`�ؠq1�#T����J��&K���c����p��������w��F~C�ϥ��~��go2v����������v�	PD�|9��闼8�k8.(���ж��p�oz������]BFEܡ�k�4-�N�j��L<��uii�H4���X}I��^�[����r�aЃ�	�M�(�C��Y��0e�:ټ�3��n�ۨ�i��:t��cc�ɓ>�u���P�W��Rx����vé�ZN�$��c�W�(���v#��㷑s�/��3dSz�M���!؄�Fޘ�oj�@��Ww���ns�u��N�M_d�4�ooM�{ݓ&����6[�$�S5�)2��ᢤ�f`j�,�Ur��<.7��V�2�]q�ٝ:������7V*�T˩�F�&eM�+��H��8Rc���9�)�;ů7h.��n�h*���W}��|�Mnw'S��Yk.c�A� �S�x��i�:1���F/��}�R���ZrE��[y�O/�2�|:���M��M9�Y�8Xr��g��o>�qgl���@��R��N0G]N�[DEܘn<�_E��Xq���9I����;^Z�Vh]ڌޣ��Nt�ɴU1�X��w=�ԝ`s4ng&�M���y"��/�,�(�޾�ػ/DNn�z[��`�s����-���]���y���'�4�J�[� �]����@��SF�}o�7X��������S��U��c�;�����co�U0�j�Ϲ��E�X.Z�(���#���������ٶ���5�=���NҫtR5;���To�X�f�*�� Wq�@vZ���1+7�\w�uܸ[�Ð��]ۡ���3_�=�OM	��w�L�"��xJ��o�;Ξ��ݼzV���w�'���v�	7��2Ϻkͷk���.�E'W�δ껹�C�T{al#��O^�y706뜂�������y�m���4n���R��+D__4c�|�T��o1K3[<i�.�I^��V��+- �V�|�Vu���1J#)b��µVl�N�r�;��ɱw�O�T��x�f[&��y:�U������R���0^�%�qn�uь�	w��[��s����w�q+��]x�^n�p}x�uţ|��67!!����;����ܮ�v�Hlז��i��-^Zۨ*�v�5Ls��P��pv��or�ؾVƝ�Dq̓���34�5�^�UyL=�o���ϸ;a,�f���b��Wa��[G��G�y#��Uk�3���l�k�~Gv�r�"y]O�Ko#;o�9�Հ���{˨gp\�Kr�+���hZ7��<���f��x(Lٝ������*��0E7^BCC�r��n<�]�;.#�MtX�u!>U�S��	�-��6���a�p\��ˈ�B&�;XZ���Lɪ� �v,y��Hq���9wdJ!��{t\��KVF�-.T��F�����Ls{[����qz);C�����+���J�p�ٕ.�I̰Q[�U���u�>9�6u[�OWr�S��䷵5ͼ��t�z�j�t�����-�i�'kض�':QPz|٦��v�����^˺��e;H�p�����=�Qw5ٞ��O6�ɩ���c�w���cT�#�%��Ǌp�0��B)3����A&�+|*��h�fn�wɾ۾N�<'5������ nn��o�T�\t�;��^i���b6��.s�H��FuSx�2{�u��J��j��֔�.uՁ��:����Y�f��2¼�v�fQ��gb�Ⱥ���t�Q�Z�ܽ�Тb��ڍL��ZE��}�I����8���"	������k��v.�������`�~IQ���F�^j������	���rдt�`���E���]�K���s�t��8T��j��887-�
��೎��J�YcM�b�Ѩ�h���Y�Ym��̨��D�cy��>H�.���=`�'�FU�y�i�qp;�Mo'�v�Nw&�p�d�:,1�a�pڮ�:R�4���5mLW��c�hXM�̇���R�ʸ1kv� �f�s�Z�u�ǝ������,����R$&����iH��z�r��Q:W]�໻�=���q�h3���Is�s����YR��Gp۩���|��*����Vf�[��i���zh�����}��Vݵ��w�u9A�����:�&�2���$T��[F�<�No�uȅ^�.�kx��ι��+��5�Fګ�lt�1S��C姘;��u���Z[,Y;�����Q>�ȱ���n�#���u('����-��34�7M���t��t�����^;�.�$p��+
|+����Wi�rC�te�7��+$��t-�<TTc��Y/n�=֔��z��d҆�F ��,!�M�ȵĒn��>�s�I��`|�ֹ�}y6��m\9ծ
T&����,�V�k�0����e<;%����K>�s�,�C��m5&naR���$^�a�4d�--'N|B}d;/nm�R���R�����[+]CǦc��S2:zXX�^�5��m�[W�kh����8⦪Yav˶�>s,�}-�-K�R��wZe�Gn�O�U�¡�XӃ2��[e{�=޳��Bo��BU�:���+��nU嫁q��J�^�zO'���9�{�o�>!��ᚱ�>�b�;�jXد�n�/x���;`�����3���,8��}U���țz�m*�uH�ww��H��X��&M�{���wOkF���gY�6U�ѥ��;�GOq�'6{<�]wpN���W�WSzrs��V��7�Z�1�0�o������]MR�@���m�u��̉R�s��/�	[{S5�cu����dK#I]u��v�.����;S]�do��cz���6�������O��}iT��(Ool��p��4Ű�=w�(�TR��x���>[C/S�_E͎EJ�o���-ku���+�ACU�P�k��B�[�ґm��ʛv�s��(qڱ{|�3��,�9�a����=��B�2U�a�ie���G�VPsK�Co0@:�h�	���U��ھR�j���B�"��Ȧ%@kq��٫��VU�{@�7r��ѝ#���B$d+{i���'^`|��v�Uӭ+���yk��h����%�7;;*�K�n�O[�n�E%�(:�d�B0y����z�gK�ҭU�[}3,BE�]e�v�R'^��N�$�{��ګ�1wCe>݊>K���Y��.����Y��j�_��s���}�.<�-��^�/c�
ś<��d0��گi�ð�@|��:�����t�S���M}��-��=�-t3^w9R8�^�3e�%J�|�ю�t��Ґ��LAz�,�J��v)O�w�L@:˥+��'P�7ƌ��{��V�+G)Y��;l�뗒���o)4��m=]K�s��?���B92_u�7Ո��̵�:U���U�/X��S��5\q�V���7���ӯ�N;8)Gݝ�������k�U���ˊ����r��cH��//{o벸U�Y�1������Z�N�wJ��f-d��!���>�v3V��٭x8w���G�^�"԰�����n��vH;=׍1Z��m�ϵQ��M`YqJ��H>ʱ�Q�(��Gc��Z*B�z96v�J��]�Ё��r_K�t��.��Wm�(�#�xK�87	k��Q$�j�X�7ʖ�t|�:T���5�z�5�򩕍Ms�vl���;���ӌf3Y�����<�n���qX��f<�X��Asab,����Ⱦ�f��N���ϯ�X����wO9UVtq��3v�ܖ�nc�O�|���'aGj�CK�V��hwL�Û�20��\^�̧�S$x{Vk�c�=ݜu�J���S���dǴ�Y�Q�dRBM��q�-��%N݉k�Neӕ�<��-;oo�ޒ�ْ�;w��6;=���G.h�7
8p����3�'�\��wx����g���T��Za}B�ı�9Y�Jo��ښ��=`-5{iD���8�f�N�� >0Ir��8%��� �r�tdĐ}@��9-���P��*Q�CD�6�_$�1��jv��Y�L����7:���~��PR�d��(�0i�U!IɎ,�|I'��D<]�ICN�Y�5TKGa2z��v�.fm׷[�SD�wT��]�CY��]��%w
�S/OnҍVK���o��$N���sx4�n'Q��r�2r�̙bֺ蠔zh�eĦn�*��6������X�J�l+��}����.R�]X2���
\����4��2�O���
�ur`�&Ώ�K�֡�P��x�w]t�9减q(�: r�>����s����MWu;�vi��_dU@U���5�=A�e^��s���V��M�}6FZGAae^c�Xr��阢��η��d�Q�U ]���u��l��kR����(��h�ۢ�WE��it�w����=ͫ�Z��pl'ԯ/�j��\�[���m�D��֪��,d"��`=M�!��$F��䂵k�����K�-iX+Ww�Y��R���hn�}���WXXU�ҋ]*ݾ��{!��i�;�R t]Z�H�I!�,C�z�S�nus%�GAh��]��
eorN�6�9�h�Ve
#�rIdS��6`ۑ���p95HU�ݼ�J��m�l��݀`V��֋\vN����cs�_USǤ��{kD���䎸\���ϕkr��h�F�}V8�G|
ݜ#btg,���j��p����=�2l�K���9��g,�M7�I\	'�v<�\�%K�|���bHww	+:�}�3��nGϊ��;�]]{��:��E��ؼRA���,R�Ɠ��u{wTy�$���!Cw�O�tb�nmWz���f��X6�l��1�H�XAC(#\���pt*���NUso�����L5��V��|q��ǟo��D�v҇�����6��=�wv�j��cԫu��:��NlƇz��6�kԚ}�O�Q��V�.g��J��k7,�!;7�k��4K�H�(����̶0���D�{B_Un�I��4��wuwv��uU霟.�͒���n*Я#��Q����;��P�y;m�i�0�`�F9�W��aƃ��.��i|���u�N]e=����:��$��+��h������r!HU�7���S)\��к��㰍�wW�R�d�q����:�K358PwY�!�i�UM׌�en��]�w��`��X�\CO_2�e���z3����u�<�}r1͠�o^mb[�-�3�����릸J
��*��f���M�7�ֵ��ʋ�ɍe�a��8�f���^A��u��f�ǭn��m*�!��b�����z�w{��Š��[E�M�1(�W:oFVS-��]�O�Q�:Z�|�%H*m��!�Qg&ѥ`�qF��"Ib8\A^VTr��9yj�A�!H�|@��S�[Ѳ'z�W�T ����"M$�r*NU��A�c����J�I<��ؒ@���uT�9��� 10�)e񠉍�F�DF�]vInā@��\	��,vl�F��l��Hz�Ց�B�3$��)�J0���D�ϗ�xg�N��ţ6�4!I�jG"h�S�Y�"EBV���̴�K[<�H��DD�m"P&(�$��L��l�q��!�!��L���*�2uW5�`14�@�`-v��:	�˛�$�L1�6Ȍ$.>�d�DXHY��%$�������n�*�h�P	�I�N�xD"Yq��MƢ(L^��I2���7���T�h���H�hHCa�ق\Ov��7���DE\-p� R17n��a�IG������ݙWb��%� a�f�4�t��fnۗO��3�\%T�c�H��h�$������=�O�h�T�I�1;^pZtF(�!J!�Bם֚&Ui��R����@�谨k��9+3n]��Hl�qJE�%�84����q��S �R��g�}��=>�
Gm���$�"�Q66���фА��%����*�-!�L�HRP�`�C"F���*���r&�Q4Y����)�ݲ�"ș6�5i��Z!i����i4c�CDcq1��DdF
�/�N��ȫ�Q:��~x�]C���
�:d�t�����P�Y�2b��D���A�D���<G�q�$J�L���ک�1�Y���BT��H�U4�6]-��c�P�Ͻ*ޤ̒4R|1Fi�!]�[8J����%�&J�	��l�q�\~�M��0�[�]��E �41��h��	H�gf
���>"��N�"6$�6�d2�
}7f�o-����X1$I��D�M��+X��PاJN�HB������$=��P,��HD�$�
�. dI	� � �6CH��m")Z>�g��T.8�eё��a��Y&ru��s��w��O����?^������??�	��R$ ���'���7��|�s��~�➟�d�6e:՛�i
�L��Ta��v�^Y�o��Q{���fh� �rmF�fV��rJ[���}�%���h0u��Q�N�5\M���tk�o��������ԥQ�w7�Y۷۞_/5�늂��������"�"$��D�/3���������Qa�685�y|�H�vv+4*}����G��H��D��)m��V���X�院��[���˥��=���������e3+�-ܷ�n5��n��Ò�N��J��5@��N�b����'v-GC�&P�ʣh*�i-���E�����0�s!��%sohY����W�uʦ)Э�xz���=a>.�m��l8p`ݵSY������Y|�6����CoT��\B����1H�b<�t^Iw��$oU�݊ne'/UŻ0:*��D$��gک[�m�eV\2d�q�'Gs��
TK�.��:ʆSY�[��c��de�j�m9Q峥�B���_.pSC���է��7�]H;Y����LHJ��5�黾 ��V�yW�k�6�Q=N:�c}f�ft�m3���<x����c�Zֵ��k�kZ�kֺkZֻkZּkZ�MkZֱ�V��kZ��Ƶ�kZ־�Z�V��ZֻkZ�MkZֱ�k�kZֵ�k�kZֵ�kZֵ�|tֺk]��k^FƵ�kZ־�Zֵ�xֵ��ֵָ����������kZ��kZֵ�kZ�O9�}����L����=@��G�y�s%v��\�*�Kv�O�������7gi�S'�����ڣh�b�^������%�ʰ���un]�Ǌ��铣�"�AvfV_�>�}x�u{�+����W�5<�w�T�3]�5�ػ�К��S�FN���:I]xa��u�-{��mm��-H�tOnVæ��5J�F�-L�fC��j�B�[Uh!;�Xl��3I.c27�[O�>��[�����/����e�u2�!b�Lma�3�6�����,}
Ө>J0�׹vk�޾k�+:s�������j;�9��^!�'���)���V�ӨXxv�=OHr6��G�L�ɻ�L���16��%e�<xf����S�yOw'"l�Bڨw*�"�+�4���$��-�{7T���֟[�7��wOb�ֲ��Gu>$v�U�y|:t�MΏj��\�Dw!�Ϡ��g&��u��.�&�^�|��_*]otn  �C�i�;(�"劧{���� ze�V�V�EKX�B)��1��WT��K��:
��a�t񳃠����^�_���=��kZֵ��V��kZ�ƵƵ�k�kֺk�Z�mkZ׍kZ�kZ�5�ֵ�kZ��֪��cZ�MkZּkZ�mkZ�mkZ׍kZ�kZ�5�ֵ�kZ֫Zֵ�ֵ�kc\kZֵ���kZֵ�k]5�k��������돯�kZ��Ƶ�kZ�Ƶ�bI<�g&wλ�N�ן:�ΙG7V糨暧T��نV�a��
���1pԝ����;�ț��H�\�Y왣� �����u& ���R%]���#F��F��9�o9�a��c78/��y�J�f��^��']W��� ��!:�L�~�0��[��b�fc�gBE���)/�֦�u�4���K6r��i�����H�ϧ:�A�V4�OVn�W��ή3J#nP�:eG�mxu!�m��l�{V�)JWf� u�3d޻�nP$`���%r���򽴅@s��B5JeD;�tVE�M��/Y<4ODCt�j����\�&��0=����a��"^��b2�i�ش8�C��Ρ�����笞����
�����@Xn�Μ���S�!Up�U-x�> �e�)��JA�����Q���8C���	2�9өB�,X�DUA�c<���9���R�-]���I'��8�[�-����B�{[~EE�T8^k�4��]A��!.�������X�A���פ�m�a9��l�ݮ9Ąf���\��rxѸ�`�X�t�j�gj�$r����*���ך�)��vȞT��Ou1�yp�z)
#C�\hP�(�7�UI�XzKKk�{� ���*_ �i����ݚ�!F����CL�=�O��0�M�减jfC�b�rn�L6��0�꯵���F�u�����]�Wm�H���gf�!���R��t��O�.�A��%*}mR��E��E�l��fkܫ���-�&�����������[�r��Fr�r����+�AH�秷���5_ֵ�k�cZֵ�k_Z�kZֵ��k�kZֵ�kZ�Zֵ�Zֵ�ZֺkZֵ�j��kZ־�Zֵ�kֺkZֵ�ZֻkZֵ�ZֻkZ�MkZֱ��kZֱ�k�ֵ��ֵ�ccZ�Zֵ��}q�kZ����___]>��kX֫Zֵ�kZ�:�N7�ɽ���]s���$��͎X��{�v�7m�\S(��ґsi��
�j�n]�R�oU|+��ƍ�W� �D�2�����:�ʿ��6�r�5��NP��>���툮&��ɢ<���8`�Vn��h�8�
�96�ʝW��7!�\l�*r�MY��~��{�h:��Ʃ�ڭ�ɥ��3B��(��b��DQ G�����M'{/����IP��N��80�%�hB�!�uO���w��]���R�����a8���'�r����_V���=u�\�ti�%.�·���@�萧��$�P�Wn}]mN�
�W�6�uޱۢy`S����ʴ�W*����R ��F�^�׵ԉ�Rj2�`N}p����I.��5�f�,����*��3uv40A��wJ��@H�m|���3z�����M.��T���y����Yц�y6��Fǣ6,Ka���>�������]�'_�������-�c54��Z�z,�1�p�J�"�Ǔu_ț\�ڝ6IݺH�C,�Ml�����sN�H�31!��KE�b,�E��}���$P�'%��Pjd]��k�׫��1�}k���kX֫Zֵ�k�cZֵ�k_Z�kZֵ��k�kZֵ�k]5�k��kZ�<kUZֵ�kcZֵ�k_Z�kZֵ��k�kZֵ�k]5�k]��k^65�kZ־5�F��k���kƵZֵ�kZ�kZ�k^>�}}}}}kƵ�vֵƵ�kZ����������3ε�����_TwR���Y��E��~Ԃ��pq��	�f�DR�����{o��y��ӽ2k��t*=mldGL�VR�N�+k2��ST�V��W���f�C8sr�چ�j2�]4��Բ��K�"�Y>Ų�5�����v��Ϭ��t��w6HdZ���Jh;�R��Kp������%���L@{z2T���'i�v�=uzE]v�á=ݻ��t�o$��V$�sFN����T��'�)]�=�pF��u�L���N��}���r�l�6���X��K��w+��B!Х[��z[Gn�<cҟ��˛�T�O���ݮ����������m�tOq�CR��7M�WhHR��u��V��[���%L8�s{�+zM4e�qn�Cr��z�+��0F��k�t*�K�ՌZ�еW�����0N��}1�u�Y��4�]M.���z��n�ᵸs;�[���Jڹ�5�V��;eC��]g���{RlP��]�2��U��,��TJh.�Z�V�4���\�4��ʹaln��z�ž��:���#�̯{�gsL�����%�O=]�ʮ��muF�^)�^~~��?g���k���kƵ�5�kZ�ƵZֵ�k_[ֵ�kZ��kZֵ�|k\kZֵ�ZֻkUӍkZ־5�ֵ�kZ��׍kZ�k�U�kZֵ�q�kZ׍kZ�k�kZֵ�5�kZ�5�tֵƵ�kZ��ֵ�k�_\}}}}}kZ��k����{���w����~�@�,��R���u{"ڶ��:�4�ܒcR�U��a
�k�u�IOl��k�Q#]��	�{�_kt;o��(����ΧZK+��w���8lܷ��M�С-�bY��U�aO�Ț L-��A��i�T��7����x���-�$�ڬ#��R����[-+]g!���n�i����"��6EGÍ��dԖ6+��iY��7���yo-_wfu^��a�3�%��>u2�b�nR\�'|�JU��OF�t�v� �"j���`����Uhr�
�Ԧ,��vR��n�����(ө��g>$v����T��{�ә8V�N������ӭ���U9�wr%��;]Q�K�
CO�8�\�4v��:P!p�Ւee1M�������ƅ�|1�֑���Bu�4�5*��ϑѦ�n��H�J�)��M)/���\�;n�Ve�uR��sF2��H]P��[��ˮ�E݌q��FJ9����H�1p)��n�|T�$KͭR�;GA�{��;%-�\Ŭ�w~ �����M���ꁺegz���YݸEd�\�����DS\;���B3w������k�k�Zֱ�k���k���kƵ�tֵ�k�kZֵ�}lkZֵ�k�U�kZֵ�q�Utֵ�kֵָ�k_�kZֵ�}lkZֵ�5�lkZ�ֵ�k]5�k���kXԚֵ�k_�ֵ�Zֵ�kU�kZ����____Z־5�5�k]��k]���>�^g�ۙ>nߞwh�5���4��f�]�K@�.dF#��f����U�xz櫻xѮ�h0G3���\Q�݆w�,2�j��)���2�%���J[�9�&
�j��x�GD)��b킸`�,���αsP>�E���n�3I��tyP�˗ݰIx�띨�+�0tc�*=ӣj`l1�F�_q�j�M�[���hջ�==/��S�8��;l��g��h�pS.�Ub�Y��FKzo��.��yAH����ꔧQ�E�wn ^8���6�4+N&�H��+�2�{s��;N0�3{�.��Ua|a�
gH��wg+ָڗ�,v�GYaD�^F���Jg��s4�9e]aB����AUT�H����1G�r�uL��%rbL5��Di{��!E��V�ݺ���iV��v��Cm�@��4���7c���M�&�����޽��մ����)]�vP�uv�Q�6���Y��E\��T�OC�{l^��7��U��=�ڿZ坙��x|���Xe��G� ԟ4�n�����CYw��U<�X(ԪU��G�llLGV�q��'�{q ���������|�IP6���Th�2��b������^�Ls{GD�(��µve+7�V�CFk�bT_!q9w�+�.���z%�����ve΍2�"���<��mԭ�b�)t�6[�bw4�x�p�cx� ^a7�����w+[(��%K��w^�T���V$������eǻ�s�f�U���8v�qܼ:YW���mc���d���;�x�ժ�kv���N����aX��os��*"���4V�8���PH�+��9�N�(��������J�'%��؊괸AN��^��]�խ���{Eh@��2����UTʵ��P�"�םr�"�`���*h��ػ�vuW>�Ac��ڄ��������W���s%a��u�l���	!Iٗu���{�9�(�a�I˂-ͻ��S�KN���S�%��Mj�ěZ��ɝe:b��^��ɤk�&�m�곶�\�+#[�*>ε���FI8]���<���R:�WA�&��E
��N9.�py�l�����E�l��/,$wBR�@b���{�n#�a��nV���eލ����ݪB��v�7sõ[���M+1і��t!�xL̨�9W6+�E�ooP�f���s-�[9�U�U��C���
��>Z��p�t�I]Ǯ�Qzz��<㷛��3�B�{&���E]��[|r�R#Ϙl���|hY{��a�P\9K4��PN�'3�`FUev}'*�cz���V�������=��uc{��\���.T0�"�Nħ
93�����BF|l5Y���6..8���7$�F[���
����C��)��M�/}c-֫��®�nH��R6fyJ�Ví�y�+5�a����_l���|	�K�Z�;���e�w�!w])�R��5�E
���-t�լ/�m�W/���̩h�)������<�G;�W�T�V���Ure���Ԯ��/f�b(<j�a��f����G�U!�|;�vN�d�MgEk��De���3>FJ�N�4�|�>e!7%��4�*�F�m��j�wl�wq��z�\[v_bY�wi�H��F���sXt�R������͚�<|z���5C��] ��d�z���ږ4�wm��S,*��+Y'o`��]��N��������u�P�PK���2X�C5�|��p��zE	�b�vy��!�[� �990��5wmMV��澘94Y�)���%/�QY��c ������sys�Q�Z����\�X���2v��r�����Kv+�jwt6��/��n����I[Z��7�E�4�V���Ow2Ԋ�qG3F��\�5	7����Fo��Y�^y���М�(����9V�>�YR��)�V����]�uSBo���v�%.��d�̳�f8r�\j� ��\����{�X{�V�G ���mͬ��s2h.rJ�H�:ɸx�N���o]�܆�v#7/�S'Kd����f�h<�32�f�l��]N<9���}�hG(��[ʡPn��V��v��4R�m9�B��%�Bܤo�ˈG��9���e���۴�Z9VU��%����s�v�)��d����#���b�w�H��t˕g�oE��P��7}ګ�#ƚ���L�to�	�Хk��JVe.�訦��YGy��
�J��,�?���������-w_�~���ٿ�?X~��߈������Ӧ�<211�(�j�B�&Yf�E"M	�t'���)?t��m3���B���F�)#m�S�B�Ha�ꨓ*�����RN�d#���#L҂ԥDZ!�����ͻ5pb!߀eV�� �Z�K�����X�[�j�)�̔)c-�m��n�`�ME .�g]ged.)ۖK4�ok�0���z*���x7����=A��R��.Lג����>sx\�����v�����x.�3X�$��s|kW��6k�b̤��@�l�ki�x�UCD"9�ȧ$i�x#�����+X��fdã�J+�Y�jJ�l�6����Sm�݋��N)��a�O%F�nsޕ��4⦰%"2�;Y�MY�!u�\gSNV]᧮�WQrf&N	N�찾�T Zγ�,o�N�R�m�ٖ�+����c��FiZ�ha^�K:���#P�{ñv�����Ch�zxR�8V<鰰�%����+�9=�&��[���/p�y�F7�.d۰x����a�lI�xV��Z��6l��C�̛�kȴ�=����l����q��|��֍$�=]ٹ-e�fc���YY�솙�:Z� �bෛ��p�Y7-s};G��Eode�ln���d�������Mq���u9��D��e!��WF[0��J�B%�;)�X����a��b�
�[�@�O��*�]�O-^H[N(��&t!@��HT�ea��!JD$��PH�\��ʍ��6Ĉ��a�&�f�dD`�&�'#�Jl��M�k-m*e�hѤ
b��-ǻ�C\�ܻf�D�=Ƶ��}iY,#����޹��1c��ƙj�`��7WX��dU=hĶGrL@�m����QTu�b(�EA�VDf\���ɩ�ٹ�����{;;�7�"�F-�����F
��g��&1GT�,TF�-j~q}�G���)�V�q�UA{<�����nv�۶�ǯU\zI7o-NXIl��(�I�°�-B�AQT���գ
�`�{$bI�Œ q*E4�(@`B�ҪȲP���$1SP`B�
D`*�Lun!UE���&"�
�%jk,�`� Ym!�#U)l	YkV#FHWI�	�J��Ku�W����Y�\WO��۷n��ǯLe�@�K$V���mJ�U_�,$묢�"��)Ts!��H�YJ�2��1����Q��X��[
�T��r[�*�L�,��S�c����v�۷����W'ӊuK,�1�\J-k��Ҧ(�+Z�D>�)��X����f6&��P��c2x���o�<{^�Uq����O���9�VhB�*�X�H�!Y�f)�A*"�(�s,�ד�̖jxǏ�|x�^�Uq�_*}��-��V��+s&1eml�1��\b!iR�`(V%K���*0b�Z��-�EƫZ/Z:����~�f 4,UQĤZ�X�E����(�Q+m`�#:ظ�73�KH�@�2���U���3D��i��s=̙����QB�v�;ò�U���k7_e
�ڍ�(���x5���y��uwf0X�کp(�I�I���pS
��(5�D�$��O<{�;֛��������{�Ul�I�*�a�>�6W,�;�n�s��I�k�>È����r�vS�o���zRͮge��ٮ��pVfʙs�Bgc�>�ϲ�] ���-���2��ѻ�
Ҽ<7�k(d�lh��;�f���ꞗ�~S+v+f�����5Ur^Ͻ܋L; �7��� MzV���3(Шx�]�JNJO��v@J��f�ψ�����!��
'[/6���Icem-��nl�+�ښ��o{ӏ��q��+uե����ʳv�Iǒ�O��qj��^�b;�hyK�`(>+U��~�Љ/k<|�N��)h�
l�آ7��r���\y^T'��J�j�̪���#�E]���c6���P�[$%�xE)��٪{+_�����~T���V�
���=!�&<{�����y�hl��hS�#���Y�����P�1�t���\��֭ٽ+��j��e��O9�0�wA_T]J%��=)��n��"-����}%ʗwz����A���>��m^�:	įXo�ѡ%�{�W+�-_�Ow�א�kǮ�9����XS}O	�ԟ*�C���7��)�hN���ڥ����n�3<ú�~|����3{8���Ʉ��j��{�m+�Y��8T�{�������ug�z��|��vT��w|�����{�἗u��0���x˜�����ث���K�^�[����gn��/�������$2����3�`.�R{�SMx{B���t�-ێ����Y0-m�	(Ka
���J���n��lz�W$UH�Ւ����&��\�ܘ�Y2�Wmg@*���>��Z6���Ԋ��K�8^m�Y5�lE©�aȜ}Z�]-'/S{*-�br-)����h��{uVZ�wk������$5�(4Tz����U{����M��'Tݖ���S(�]�m��&a�Cevp/>�a��+��=<��}T.Y�B���ԯ��m�9[�P G���| �̥�I�B=�m��j=�fME�1P��$UN_s��Ҷ2�y��S���Ӑ��1uU��=� �4���ck��Y ��p�+<�S��^-�YW�ձ;��#ە7��5�y	����e��==u�{</��3���ߛ�;E�vg�N7x��ti���.�,$X ��/c�q�ݩ�S�.�I���i9F��v�P�PրR;0w�V,h_�j�?m��}��}��5~���
�5��rT
��"�Z��~��+h�=#���E��6����eT=���]�����j��u��J�L�i�����Ф|��w�q�ٳM��;�F#�X��G�c�~���y	����yy��My�[O�]���à�(��3fe�jZ�hh�!>�#�"�	�'a��$�Q�Pk7D���K!!��ojqI��N�>@*�}W������fz����݅n(��;�\$�d�����1ygtog��fϪ�Ƽ���)܌�I��;oC	�g:�l��ʹ�:�l�z��d��b�!�u{w�e��;��Vؽ/���UH�������?5�=��Ԫŗ!���cGJ���WX�k������'�$=�~�f��T|�ޡ�kz�P�=�x	�{��� o�D���TMN��y�8���d@iُ>CK�v�o̒W�sٞ=ݿnQT�\��i��z
���I�h�n_��V"`���{�o�z�A�i6Q	b�	�ef�Bq���q2FSfǶ�,>J]�Ӕ�M��3�1cj�Mcb�*��:y�h����� ��jV,�	�P5[�*�U<���e(/������U��d��[��l�I;�����Rs���&�k�RԲ�̰��RR#0�ny8*�04��ɩ�Yn�4\b
5@�����Xf��\\sPmW�A�,�goN�����8|�;�����{���J6]>b�Y��w����>q}�߫4�����YP�s��`sc�]�� d���־1��,�7��doԈ��*�Զ ���mE��?uq5|�d����p���k�J�'�t��5κ�u���lI3�Z��v:]����Μ� ��K=qE���Y9S>���	�3���Y�e�!%��!TA%R	+X�@/&n��S̧j����m�K����El�>2��B�-��ё�=�E�T3q�7ڽ���*�ܨ��E&�e�l(���A�H4YMQ	3�x�=�B@�iޑw^�X�IK�U$IC�6���E�Tƻ*�J�Qž��|�ӵ<��;�O �:���lH���eqt�	��_{?�h�A�_��ǻs'o�0X]������f�AN�[c��D����[�,\��T.��̢����I5HA��S�9_�h�C@�~4'�xɯbL���!��+*���2w�ץ*����_�#Xnj�M2����*������r���A�ˎ���0���|����k�Dz���������Tp�Z��~�*{;�7��/{��u�W�}��*����/u�7�|e�m�Ŀ���y{�6� &���*}�R�]v��*������ՔĐEj&����.n���U�e�\Y�Q$�ry�)s�L�}7A������nJ�҉j�������Ҽ�ʝ��
4^�z��e�>����u���K��H��q�a�sDW���C����R�GU:Y_#tZ�7��M+_���}����M�>E\��l�=���Z�iE,s�Χ}Ir��>O�X��ξ�]����ܩ�/�ӷ���Z�k�	y7����@#�c�nӠ�ůI`�Y���5c{#R�B��2,n���	�}�/������א�k7\	�ց��$�����w	VFװ4>:�c�\N�k�S1y��|�|�+F�zwӰ��|<m)���	�А�{�2�<6Kiy��-�h)���㞄٬ؙ��>z����"&�׀��	�k�Ł;X$��aG����=o Y`D�������Z�:©a`��{��}��Woհ��ٲ�>q�#"}B��v���V�R`�4�ӕ�<c���I2�H�7�Q�{F�Q�����1�z]��<0�nL���@w��ڧ��a^��ګeRG��`�ϴ�g���զ��À�[��7.����v���Tzō ���!#BahG���^&�����kiB�1E����PH򯝾O�=�9��(�S�X~�a�^����mo,�3:-��9G��ZƷ{�C����X�Wo��t���r�`����>O[�]��e*�\uɮU��eV�N�\v�<XD��J5�2�:ޜ�Y,�]��
�  ?CX�yj����H�
�k�#�,)��P2���q�z�U]hJ��-s����X�7`^�#��m逮>
��UGdk:�3�j#&Dby��jU�M>��q S����~�Z�b�5]�X�v?-�����Zk2J#�
�{�2ۡ<����J��X[:F׮�*����6�;�vG��i�p�܌��' �f�o<[02�չC%`jYV�G�|�����k5˻�N��#�RTk�ls�F�l�����M��V"�1`	&ʒBև����ʼB$<�^K.<��PJ�k�.�y�6��Q���zy�N�m��1n�Jsse��M���o��g�	��]M��i�5���\)�E�͹�[�y��l�2p��$Dc��ir���QW�ZU%�Ωe/TMϵ(��S���'6ܱb#6�)��n����o,�Z����s</#�����H�~{�sw-SQٱ��[P��ǻcĀ+WCJ*J�(������xgcΝwM��m���gq��������cXv��*U��+f����]-9��D�c��Ԁp1�������z����T�%W�/��OwJ��1�ϴrKe��{�/O��`�FI��7�B���̭�6�ly���<ꧽ�����GY#�@�8*U~����c}�.�������.k�B��������!�q�"����T���C0r�/��z+ƈ�^3�	!�TخF�O|)X�b�=�ݣ>Ɂv;_{�$Yꥑ~{kFki��O�Dl�h��O-��|�7S ���v;�n��_���j4j~��^�Mͧy�+oc���[V��@�X��:}�W
�a�N���0%�٩	{��{�h��;*�n�N��c�z��Nz�ޡ�W��X���H�	ǟK��Y���'�z-�g��dѠ�
�{����֛NUO}�5wa�W�4l�;�)z��Y "o{�\�#g ;8�T5�>���sϻ���-�㪂�b�C�V&�p�핈&�F(����YSt]��;L�"�^N"b�(��M���p�t�M{��uk ��L��v}D�EB*���;H��	�gv�9��fsu|�V�	%���T�Z�	��ـ&�*��kF=��$2Bj7��!p�'�$,��3t��f`�^j���ȤP"H{��6�ލ���:����M�����Z"c5�`@U�4��AX���6��Ƕr�H����ЊIkͥ>��1�vЎ�>S�V�>Ȗ�ߪro�����Ѵ��k�k蚁��A���wV�������6�����J�N������t�YKTN6��Í�,m6n��Kvm�n���ej���\ƕSL|}�*�er��w%W�W����S� PN�XѾ���y��?P�}�/�L�|zVA�B&Ec$��h�9Яcm�]���~kk����V1�x�V�R[���z�L���!`�i�Ih��rn9��M���^a�_�X��Ӻ�o%��:`��L1 mW��w��g��� +}�hvz9��@5��{(������I��OB+Q��lo,�"���57��5�"F����'!�ɸu�����Y��۝���e��;\�����o���j�iINU�Yn�&���U�l]wu����J� ϼ1 �6&2�v���/%|�R�;���ٖj�`��ҏf���gF�Ք�{>��t�AQ뼠�G��#����}���r�~������n�3�~+�ؐ0��iV��f�%^<��vw}�ک���"%������IY��ｂ�2Y��hFE�N�Y��*Vr!z�b�W�v�{�y��̪6T��]�U�:6�3�N��_)���w;=n���g��6���Zc��+��Y*��U� �v3��
���++Աl�ado�1��,�I��!�L�2]��l������jw�G˕_���q?y�'���ff��e'�e�Cݹ���uez�90�
������=x��r��>bյQ�o��{�x��*�$ ���h����~#,��  �&y,�,��箚�Z?E�K�̦_�jiД?�-���cG��?���oO�g�v;I�osq{;����r�@�za��:wPپ7w䫇/`�����xx�����p�ٔϗa�sM.%eVt�/���Dꎂ7�X�p�]5t�9ݵa4�H�n��n�,Wfh�r�����ݣz��w1R}4�B4{ft�7�6}t�u�r]��������a�2���w��K��3�8]�Y�d"�|T�.�
t�v�ͳ�
|j�,��g:#�.к����6>�M�l��`�}*�fe��xW��j�i��Ӭ�Zݾ�Ʀ����+�[s���>]���o�lIVw�ꆟ+3��g;���\�C��X��w"H�5���=�VunZ��]�nd)H�0NlB­�b�c������r�/o����$��Z׉V��L�Ԇ\8�$ڏ2���y��˜�����_U[�`�r��h.s��0��
r����M8A�T���+z�V*�N��VV[,�,�}��;��6���h�Y�2\��)c5���=fG����0���ng������3V�6�����QT�6��뼣�;�Aӈ�X�+q�B	Bum��]����Vх&�//��3yVˋH�MB��/��)�g
)(5z�޹gKw�9;�k�eS���P�ɶ�dD���J6�iUR����	�������v-DKV�"7�H��l����s(�Z�$���ґ�j紙�CNP�]ۏTl�l�z��^���,Ѫğ�iI$����J�k+u^����Q�؍^��`���C�Oj��F:�$x�����\�p�OT� q�#(4�]^����_.4Z)ސҝ+�]��5�9�k�ȭ�ۓ��+JE\J��w�u|�]����}ˮ��sz֙L���I{㢤|�Z.�Z0c2��xi�����7t���O�G�d
n�R޷��c��b��{���eKl.�I�6z��[Y��q���9t�î�;���o(�rIjHT���l�CZE�v+Y�l�L:E[���T����d٣���c�hƺ5�^�yt���J��Z�D��;d�^#Z���g;��!�j����qt���ۺ9/x�e�~���JI:�.��C�Q=]��^'�P���b�]�`�ΦgQ�Ne:�#U}�X6�p�ҵ2�PÍ�q7C�i:*fpǇx���]�X��]e��\�U�WC��4^.�;!v
�ΝMu�n-�hmBf�^L������nD6ޫ�f���o=��
cܧa��H���He�-w#x����	�%���E��ݻ��i�S:�SX�G�Ңr�E6P3c8��	n�y�E��ޖOR�PQE����Q�!A"����PĢ*�1�gX��]:q�ǯ;v���}k�W������P��72�5�2�t0Ö�Ό��Ur�H\J{J��t�Ǐ^<v���U��U\vވ,��
**�
���d�*�BT=��-�ѽL_�(,���b��,�f���ssSSS�����dfL�:��*�iZ�p��b�QX$D��Z[�ȩm�m�%�[+�;v�Ǐ^�x�۹�}9>�L�d����X,8�֬�a��e�En*a��<��ꭒ[=k�N�c��ǎݻlk��Y��':����A��e�+%����[eF0G�c���#"�2����572{=�����������}8vv��I�wZŋX?!Eb�4UUTX�ݮ"*#��P�� �"�,��*
��h�J��*1Y*��V�n�N�b"��`���~�|t�T�QUneE��s3%`�XUt�MeB�QEP]��<6�7����F��X�R.r,����wt���[=LZ�Op=�Q��{2�����ֵ��y�w�/~&�F$bF$bFw9��]�l� y.f{C����p凍��3�P�W�P>�`u�{�b�N3x�^k���ض�{M�Hʬ�ez�p���,}6�\�%���b�������rx"��Ad$o@	4}�6�/�w�Vs��zHO,S�Q�l��/pO��]�'��������\��S(�`i׾�=�� �׻���1>$#����K����ޒ��3V)��jx�o��wR�5�xm����E]� 
�z1��`;���3&�)�,�8�'[�L`�rx g6� ��$��ϰ�j�>�7�H���|� 7T������AWP�\�7���Y�wy������2o����xu�
l��[����ƺ�*as�3�3�4������8���ό��d06�chρ�.�̫^�`: ���x=����p/��m��<З���@�v��D߾�x�����p�� ��i��ܪXMgl{��ͧ7�C�xEA���bZ���=��o?cE�� O*�9���d9w��"13���T8��|��E-�8�S�D�xa����{��R��3;8wz��5�;'��f�s�� ާ�Y����Ml��9dPrz@���v�祼"S���0fK�FO�9��8g��cb������w|=��Ds�3cPK�s�h/V�2��2 :u�v�nZ�l����V���[ÞJ�vsy�u����Z��on\C�p>b���|S��Si����J0�q�1E�����cO�a��۽�7�%�Q��"E��:�U5e?c��qb�U��]{�w�߳}�{$x���� q��d�C�c� ���B\���C�D�=5ƀ�ynX�pKR�|w��0��R�]wp���>t#_j|��O}���̓7�5�����,		
q�(�=�҈���0�^�_g�ծ�yw�5�4Y%2�� ]!G��@'��8,7�[�c6 ö�47�Ē[Q'�׈��������m&���j t0��E��i�H�x E�O1�{��'��O��� G���$s|Yݺnf
��M��A%��1梈�����+����ʛ�
����-w��_�tc�4&w�moj���P��� ��>��Ht�]ڱ��G���d�P<���{S�h_".G�5��޿;\P<`Q��W���\O���Bza���d�X���(P�> (�����qO	��3������>�+�� ��@�]No$����=h	��爰���S	-�i��{^�!�z�l�p$��X����6�ҭ8	��(��"����bz讏
n�x�:�����a���`#�Z �z><�Q^ @��9p�g�}(�Q��`����a�/z��P���uc�*�*��WG��7����D�N�JHq�����Vf���n��*4�
��������b�KNݓ�� �b� �B���q�s-P�>9u�W ;��U�D���AG�*�gr��e��.v#����b�ɲ�(�� ��2n)��[f��HO� �M���O$<�DbF$e���[�ӫ�_��>˷��-g3���<������	�^��q�>�w}�fM�?��J�'�O���vº31��{lu�w����� �Q>A�;3���˂|��[�@,�o��y��u��Z\a�&[.�Z�7�x5��Q��S�!�j^�n�`�^�d{�>�(.p#ɜ�e]����{����-���Qܗ���C��M�+վb@T�p�U8/���5���`]�3���� �0ꁗ�z��v�*s+���|dd��>�B���ӝ@���oϤ6��L52�Č���8��Y�\�xZw�O� I��Q��p�}M�;=>8D��O~=~z|3�d����B����[��:a���3�Jv�Q���|86?i����|&FtG�?��#�:�1�*R�^\X����$�+�'����ͼ��ٯ�<�����qa\���Я=����{�#����Y����0d��	��t "��v�ƠY�5;�p�{���ɿ�!�>�q{����y��jauġ��� aH�I�-�{e/��x��Y͊7�FN{m�e�
P ����ô�����wb^�>�5V~}D��K��>�Nl�lЩO�\o��*ɕ�=���ǩ��3{�wZt��#$nuk��]���P9�%u�k'v��,�S� �F]Z����`��^�h�{IN��'���`��}9����l��o{��{�+�.f���Č�
K=��#2�w������ �����;���������d��U��C��'�E���2 �N���T�o�V�;�x���� 8�v 8���Y�5�� [�'ÇF���@�;\~�a��&�C���Hn���|mukshJ�9��Dz��������ya�y���׷�+���B{�fk`�����0
�[V{��ʜe����Qb�g^o7���a�=��~��S�lۮ�l����=��\;�"�T8S�6H�N\U�헂!��/� ڃ#f��b�A^.�+�`t��>�{���e���n2h�ء�E�ftZq[��BG�_�:p�mu>ّR�;��=V�	��
�����t���V�O���P��=n�c�Q�Y�c[809��q��o��Z�q5&�"Abx�zn,�O�����E^_�d��0���4�lq2�ӗ_;N߫y<����k$:������`0SF�>�y䦏�ӣ;]�&�CO������쀏���z DL�c��՚�Np�4���k$����À���@�l `\�@����G��uG�1n-�@��������tz{�K}2t��Ā��>�<�Eo)�y�㉤&x�:�G�SvЙӢOC�}1Bf�Uf����kSQ���OZ:��w���a�H�4��]�~��z�����ȇ2�y��|�oEnz�mv���څa�9�����)���x.i��3�Q3E>t*R'C}���ݹ����M|~HČHČ��}������5����3�<Ohn��z����=���}�4��+�x�&k�i���9�U��BV\�޹��vM�6!�s]�_� �������6y��B)� 	Y�D��p�Q��������e����w����q;����,I��&��H=��
~^o4$: >1�45�٘�6oU���GO��^%�q����:�:M�;�#��}۶MKn|�o��sjy����U�5�h/n]m`�=�C�EH[X�9�7�ʑj;�I�=� ̭ ����XD-@G�/2��ʼ��~ʼ�jY�,w�!���G&o'�`	�S�q����'�A�CCx!��a7�ou��/�2�c��0̈́���8�9�#����Ǧ�s��:�׍�ni���{9�d7X�!O7;�݌fn$#�x>x���Oͺ�Yi�����/��ȇ%Ӣ2�8�y�~����K�u;�z;٬K&D�M�;ӊY{��r����.W����y�G2��q��Y�������߀�o3H��٬m?6*R���vH���>y�oP3ߛ��*�3�n����{�������_9�"�a�V�����PLSv��x6��W��0�y��V��IL=P5{év�^���zQ�9��N�kC��}W��Kܻ;��ͮ��<ܤ�o!��0p�\騯t~'�t�$eo	�(N^o�׼}9�����LS�g�vCqjkM�̛ԠIY�m@P]\�[�2��5�^�^�u��>��̇���M��h�4�τx�c���:}�ԩ�|2��=�2�(<H�"�s����ϱ�0�	���7�R��|������,>�/"q�`i=�����W�p�1��O>M<ٙ���^=];��Z	��;�P���ᨅ"Pl9��'�����`{��D��	�yY8	a�h�uk�\�!���X��o��Cϲ��H�Yp+p��I� �oc�F��Lf�#a�
u�:�s̕�psܟkĘ���ǳ�u�(4�{f�9t B�޵�ǈ�|��q^��5Mw\'<�E�-�ߗ��}����雍RW�M��'{@%e�S6X��y�J^+�`�I��B^�ٌf���0�܁Dn5HS8O�(��c�Z�)�+>��$���_��I�ǚv���e���`?����HQ�o�k#��MޖW�5�1���������0z���x猪_>��q+;Y��>�ÆC���jT3!d�u��)��U]�7�O��y�q6n���d���S�ti��S"�[b@6�(�J�~��P�R$��t�L�nv�ו�J�y>���8��V�`W�UA9�r>·�`��I�U�7Z��;p�$u�i)A��U3��q:�]e�]'À G 4�"��m��wz�*88�q���:C�ƙ�~�='T?����>�l� #<�F�8�/�~X�$[�\�������8�1�1/������y�Tx���	J���������V�Lc�8��KG
�!����eq���K3��zG��c=<�������{u�1�5Y��;��s��^��$�R�v���I�|��pV������g�H���d���R��!�0�xge�t�;G_�Z��ݍ��6����c-�ޏ6���)�{c<$�24`[je4�B¹7Bf8�J�c���D0�]r�U�����}�1*Cֳ���ĮS�x�c7��\�oH�?[jnn-��@?^�W�ٙ��QY���/!��/�(����$i�ھfJ�71]��v��[�[�C�j����O��Ԫ��%S2�`k
�&������~�L�f#6�e���K� �H�tx4���^���5��/����ӳ���`�ͬ-��C5݁ɦrf1[\��a�Sv3�ހd��>]��c��>$If��$��lw����o ِ��1���Q�#�	u(Rt�+�nd�ҮK����M]o"c�^��e���_]�)��w]nƹWV�����ʑ�̼��,@�H�H[U�9����X�$ߤ���c�"���f���ǔ,:�Ÿw)R�!�,ܘ.�dKw�{�V�Ww�� x��<\Z}�����(�tk���0�������U��o��C�u��lƯ���1�Z��W�;&%�*{��\��8	1�����2R����%w(�?�M�����ў9I�q�yn6���S_-��f�.�dWpΝ�D	
����1�:�4~!��Ym�X�
4��z3���8�͵Bh�P��ü�ϞƬ��s\�K{�%���@���Ƽ�݁j�V��9"����>�;�s4�է��{�|N o�=:�	\Y
�
��`~�c�T��K�+a�C\;�#[�t-�P�-�Ļ^U�vNT�,&��]�\PZߛ	(ֆ:<�^K&�����̀ML^�A�6�XL\O�;���l;��D��?�xBf�����5߾a�}�gxb��J�︙���!�Nlip-x;<�rnWB����v! ��I~��G�d0�0:��*c��`�A�:q���nuT��8{��;��ͥ�޵Y�LCN����ف~K04!�?�K���My���jGek��䯫X��͛:����}����b���T���R2"� C�MQ���:�{;���r���8�W"������j�(��K,���8[�z!v罘�@�Fբ ��CVu��b�DQ�����������.��M�]�˧ؗ9\���!��3i4ȓ6ջʒ��CH�r�ַ���xz�����xBh[��LS�y�w<	����_<摖Q���GsN���v�ypX��p1tk����3��i�k r,�aT�v6��G\>�w�$�{�(�baY���Tū"��}Raا(?�Wy�q�>�T?c�}M8�������meЭ�1�T�'�g��ְpj`O{���/���W���x�������)���a21�2���[��%��yy+�.���W��d�ەP' ���ȇb�U�P=;�K���:}�U�P�9��ֿ�v�C�/��h�vG�.r"j4+�2C4b�¡f���ہ��@[�0�B`^0',cߎlp�:�r��n��Ki�3�q�f��������ù��>Ǝڏ#)>	
��AjM�3�q��
A��m�vD���ёnϕ��j�i���9�0�E��ɂPN���	�[wj�rZ"c�6��d|KL�bX[YBp�q�g�c�{ޜg#���߮Y�����*T4����W��,|d���[̳E�2�;��1U͂�-��7�a˞�7���R��Ha��;!��D����Y �|�k���gv�e�]&��6��w�8LĬ��|��q@������,���jT�F�5�H�l9�5�����[7l5yv��k���&�>{IC�I��5:}�Y��.��C?���G	������Ԟ¸~�T�����B����������75{�-�D��T���Y[�YoHm'|��JV��WV�sӚ Sgm�*��i����o7�˂��Y& ���ݢ�l�E�H�>R�x�g>�J��M|��ҦҖ!&�w����)��馞�2>@���sstk�	�3���&�B8g2�V�z��`�a�
3~J�d��`�]~b��6q��=��Q+?z�;��=��H��ocuׇ�'o�~�$S�/Upޯ7��;��c�el��n�wLM�0�w��{�:2�6߯�[K�/�~QF�?(��8�z"1���n(�h�� ��V�^V]��� �h#wT[�����j>�߈�NN?��K��L����i�v;1Y��Q�o���U7^l/U*����������8k�V���;P!�i�c�;�Ɛ������ܕ$�m��{Ջ�����볇�|��A�Fȳ�lg>�>fG5E;3�[;r�kB�{��*z���?o<��+��>^�E��>��5m3����d,��
r|{w���g~��^��Qg���I�iM4��7�K�ݬ�A�`p�X<쎆Ft�M���ܼnj�X@��˝t+v�e*�*`�N�����	�͵0�NSɍd2��z:�k8�WcE��c}��n����Z��\�b������C��oj{��G:��V���;��]�������z �҇0���;����0b֬໾��8��R>ܴ���������H�U �8)�{2nfFU*J���Q�o�^t�����s�>�HBӄ�֝��U ��S˺u�}Wn`�S�8o���
�Bղl�o�[+�j��RG����_R�nM��e����{;\&��s[Gn%NM2[CxC��f]�������jw�vfz:�pʦ.�M�'�Q���z��կ`sS����H,v5J�2��Լ�^����(R=s����R���N�A�`��)U�V_C��F/U������{3+�$������ ��SU���S��[\\�-<�F�U��X��O�n���;.��gD�B��Z�6�s�vlE�
�&P��'_>�4���uw7�R�e�[��U�J}I5�eD�<���q�*�3kdŗd�u,"U���2]')J�ò.RM����f�$�r���Q�5���'&�U���1_��Ө�*�9�"�W��i�!ա����ۺw�xq	+4:�di�a�ڇa�Z�b��A:�@��YX�7#��HV�.6�M�%����G�t�ㅲ�٣3!E:Â7��=/�pU�XjŇ��-#)x��#��~1J�kڂm3.��d�B"�� �����_�m��Tsz�ï�Wt`�G���﷚Y��-yʱOr'��g�e���0�T��v�Y�%���[�v9�ɛ+y���D��0d�,�M�^(��m�WHm�yw�ծ:��]H�9]q�u�=}N�T��Ŗ�o&�6dŦ5M�D���V֍2�EN��.���#pV�MUu�����/e�=����.�{ip`����H��~��չl�t�Q݄9(��n�WI0�,͗�&���ن�I!;u��K=Y����l���̛oyᮤr�]���<�e8��Ѯ�n��=�y��l��Y�]Wfĭ�1D0�y����ju.g[��w�`x�zye]s.�j./�eI-q�}����3�dc����(a�6�U>7��O5.�E��²��T(�B�<6Xy�y�za�BZkr��Q5���>ײX�j��S�����"��'�l�b���x��{�-䏞���Y���f�b��ey�f��n�++^���$~���������KwhU�����1���"�جB*X�P�ۮ�&u��B�d�;�;JRǕ��eLi��}������V-�=Ohup�sU��Q������p"�I	dD�m��MV`�H�Fq�d���xĨ��i�iU!AjE`�E�
���:�D�RP26��)E
QJl��>Q�`H��@@QH�#
EIEL&�9�HctQ�TI�Z�"i��D�PI�e�
QeI\���L|J�P�E2ۤ�(��
�Z&H�(����JB�jFb��HO�����*����!���Z��(,� c����O��m��ܯ�x�x��m�Z��q�}��H��!`����{e��r�Ed�Q�k-՝d�r{2d�x���;v�=k����|��%�+`v�DU��gPSHv5�D�*(�Eb�Q��ٹ������1�ocֽq\}�e���$��" ,�\�U0eN�n6#+
+
��O��s&��Lc�1���Z��q�O���ITVC���B*�X�V[��Y�9,��۷o�����1�Ǳ�����79^$TQƧ5p}g�䪅jA`�022*ϝ�t���Z��1���ׯ\q�ߖ'Ab��\��Z�`�l� �b���X���+&�W\������n�Ź@�4����c
Ȱ]��6� ��,m�b�1E5��2�Ơ(�J�eWI
0R,�\L�f%L���n��ʂ1TTa��疋��w.��q��!F�~e"�͔z�[Y˧"y��T�(�(�®�
�YZOqCu]����]�Ew���<p�j3f��i,��i��#�6L�T.3�M@äBd�m.&�#�B%2Ds.�O����� �Z���u���|������h2�j��s�G��j�Pސ k'}[ҏ�M��5n��a�`m�K{'���⧘M,�v�"O X@2�a��m��h|P+�&r�+�j6���ۅ��zoa�Z�O��":^&�5��x	��GI��:�3�f3�	ß9�m�S�_�t�8U�xε{e�����{��׋T�޳�w�>��Dm�<�.Z73��=M|�-�w� ����Nk�Nǫ���r��ؕ����
vҷ� zH���u5[���&^J2r��~n��o�tf����3��Q�`��W3������ؙU'�  p�gr��l#�\`m%�9����̻��^]a4���X��Y���빻b�����<�!f��p�Dg%b@�k���<�g�/��M?��av�x��4�S�*���?~�,�.���0���D>o�kAE��ӵO��>�"[��_�f���,�5��_�+3�{��߻���T���_�&^Z�=�.��Z��U��P�8�>~�Ai.-|�b�,�j�m'� �\���ޙ�d;�����&e�f�S	�^\��b�|]�yl����J(��~���d�u��~(e~�Fw��PRJ�$�}�5���fGo3H^�������цg-���UA����}粒���O<��B��cU@R\��9�z��\/L-��]c oY��]6j��m�J֨��	b�4I�pn)����G? �<H��MK��S]�|�i��D9�Ǭ��1�fUF�s"�X��qS��߿V�-3�k�g��ٺC|��| l���*xim�W��EmI��6P��9�C�;bjX���!H�z�O�ۆ��]�x��E���*[��	
����e�����"�G�D6��K�F=k�p���~p�0kUT>���܄=\D_������cO zM}"�<m3��фg��v6O;lai�ᩂgG4�>l^�f��	)���/�J���"�$At^s>m���(o��������X����3���(۴o��n�k��_��<[i'�l��-�n������&� �Ͻ��L��*�|O�ICh�Ⱦ�z8S1��H��G���u��0��T�~^a0���@��|ǲ��hr��u-N2�Q�����([#K�p4�,�.c�}=����'Ͱ0�8�.���&�b��I�w�<^a��u�=�q���}�P�Zm�Pm�~��Oi������mB`�
B�]��������ڞw��^��1Q���J�x�'D�;55�
����a�X�(áwӞ�tW�y�v-��xv}=U3K�/��d����ܻ+eE���Ŝ�;�J�WR��8/�Y���&�0���V����˭B��h������-������=nsm�ɬ�r���{�#%v�Z<�.�gU�&Q�DL���#*�7�;�~_��.�?��X� �rX��X��'¦�u:\x	�d�gv�M�@vY�ϼ��9� ��ds#��b5g��f{k�3�鱾b���W�64zH���Mv%/�Su��/��,Dd8o%��+O'��TCMA��1pj�q�! ��ei�Z�j���tLn7  ����6O��>�[����&ʥp-�ȳf������k��U^��� �EڞѤ���'�l��w�2Q��u��ߛ.Y�7y��Wh�E+6�}��a�hQ���t_d�
(�����-�y4��0@g�ݠ�1�~�o�g����"�;-֊=\�m��_:%�׍�3�K�X�7��<ol/{�8Ó���ցE��;�q����p�N�15,r��f�{00�)ڰ��"��z���C��shqq� %��j���L'��;�O<�k����N��x[�צj�g��g�*�q}����Ia�����
'G�@�p���r!�7��8����W�Oy�c�{�a���oCto�/;ה=��(����1��2��⛟����к�����,�����rDxC\BK��w��L�/�f�������~�zc�=w��2��a|q��|��	�k�����R�}�)D�<0�Y�?U�ʘ��L�-S�,��%�nX�����q�(���Me*�x���]O�˽+�HD�������[鐨H����d�2Iw���F��)���nD���G'�y*�s.�����{��~�s?��F$dI��0Oxx^�]��+�zJ0�b���?�|@v"ٞ��H/�Ma'�d�8�g��� \n��b��w�v�ʹ�l��aY���#}�m5���V�s�a�鋩���M�E(wf�n��t��{�ٞ�i��7>��xs&"�p�������>�.{_|jJ|���t����z�8٣������ɦU������=yyW��� %� �;��t��%�si��{�z�&�V����=��-��8P�bw��������azW��:��(ڗ���I�
��Ƨ6���ӧ��k�؍��{�ǫ+�x[k�����ρ8�9i_ց~{���Z>SΈox�5@�Wx�x��>/骹=̹������]����|���u��� c|kg���"'=�i�Ϊmߔ�!��oB�j6&*������k1��9�����sсl�� [6�(��ʣ��ȯ���g20;��S�]���7�,�fs����֖}����� ���	&qN�S��ո������W�I��r�]_W<?d�[v��,�z��v;zAqD�����΀q;:��/��;�X����5dG<�ՙR�7�L^�ppW˪�l������\�m}���
�*N
��u|��!G:�e�߸u�sY���V_(u&jȫ�e��s!��`����J��/�M�&"M1Q�""tݛ앓��]7r�ݏ��s�6_oJ�SJ�0�Q�XD�-�P:�������^B{��ۗx�R�k��a�r�$Y�G"nE"0x�nU(�T*I�V\3K���2D�"@H�0 G89�:�P���~ß�v�Se����`���Y6G������ >1  ���}9�ȅڷ����(��߲Y��m���j����]�x	#:��X�zn~��|hk0�U;���s�'��Y��&����"��-�@n/�Olgo1��f�1��{u���8\;�?ks�t`}g�Oܲ��������0�<Ls>��vj�^��p�kvZbǧ�sDQL�}�B������[����N:�h�ָ ��1�4:bm��H�Z�;�E�[/����sG6Kiz�s�O��`����m�Ʒ��'|z&����/Z{�������8@'�.m&,,[i�"�7(����ff?s�9N����Rj1`�\M]@Y�\��R�ysѳxC0!�@c����"O~}%���г��w��8�K��ܑ�է/�w���ߗ�4uܤ0ҽ{@���=r)�0s��l�o���=��v��d��>W�N���z�Y�p|8o�2L��u���k�W�~E-�ٜZ���ĳgc��^�W���D)�j��u��u���,vSA�n�ޘ�r���bM�X�w���Z�g��>'א�:a/����d�[�ߋݮ��B��u����Cc``��]/�C]G�7�$l�Z+-��ѐ��;u�u{�yh���D2�X��Aʺ�QA`�2TEX�Nf��4tw��ȯ�N���Tށ
K�+�6>�p(N�V
�ZUÖ���P�E��c�"�X�E���)B H�Mo���z;��.EFeg���+N���l��hbヒ?�����G�;�Ԕ������]��F�j�Hɧ[�{��6�q�=��\o�����菾VO r�sBg9�.6�0������㺷����?f,??}��vw"�{�\��/%�#9����,��Y�C����Dk�����N�
OR������.�����Q6«��@2.���o֞ x����*?�Bpy|K��klgt@�d��x*/3��Q��!��&�k�k���W3�z��do]@JZę��ǐO�^���uO�;�>����۲{�gĂ���t���5��#T/��T�e1Mn�5�K$��G.�����,fu۰�,q��;�����,x�G�J'��Q��g%� u�l���ӲG[O��O��K���tH��:��>����3
x`�:��K�^!��>���c�bIr{=���i,�
1���B���ϟGku}��~�L��K��A`	"U�:~l�7/s�����M�Y�	�%���s����m�ڥ���[�Įp��[H
D��_�_9�BGߕE��n��Y���fܡ�N��K�rNXپ���-��9J��ٳm3�A�����o�g�[^3r�ǼK�	<�<x���[*Rpu�Yplټ��D�:���Q�]�`�i��L�<�_+��y�\Ϲ/9�1���gw$��I��$�H�*�BwNE�9I9#  3�i&�� ��(𯻽�pަ
a)`$�a7y��AN�i+��m�"�3Yr�֑~���m���5u�+�t/e<�$o�'�Y�8�"V��̈��~�=��/��Ky��^G���Cy�'���L�^z�&M/�x^ \�L3̌�4�C|�G�����ڄ��9od�ؿK����W�߇Ï�Ϗ���A���F#���L���RA/��΁��"��ii�5/�Y�ٖl���]�@�h�_}M>�Y�q�s���~b�����*�Z����������kd���B��2�{� �?�q����{��%�����q�p�c�5�=�/ĐzA)���yy:��\us���)�B�_
���q��?���`��rE5R�<'�V�΍�!������5,�=�U��sh>���x0�D{$���Rɳ��e����gh�&��4��4��fر(��=3\j����zm�aa�M�RpA�c��)<���6E]���$��8Gy<L6C�B+�ȭS���o �^޸���1@0O~1��q�Y���z��T���y_}�f�\wߜͼΥCBȇ���7a.C4`�o��,�����%H��YRT����]�d�VÎ���6!�gU�3.��׬]j�uC�ˍ�:*�P\���Y�zK/��| ]ܨB�M�!W���䐧���j������'vI'"�KDX��I���r)9HIlow�������88&i�
0.������A����2�>��S8�'}@21ͅ>ݮzڝ���)���SQ�ј�h)pH���.�&f6e״&��1S�̼A�p�:u�ݸd������3C�M��-�ȭdl�qΆq���d�z>������g5�+��|������T_6��h���AO{Ѻ�{S�%��D�6��z����|U� %����c<>�jla��ǎ�L�����\�G�3�� <��jD����Z�����*�=Z��p���5�$L*'�|�H^���#|M�Ր��ߵ�����N 7�Y���O�u��}��tO����̣Ъ�_���c�e����Z�Dp-w�ܨ���"���|s`X�+���&7.�����g��|��s`O�2�C���zY{��4z�'3i�˾�}���{k���@Qp!nF��� D�O��{
��8g�>���Uy�_���x��|G*-z�n�g)��6~y�&%�!����������$���N����.`9��w5�����(I4�t���]�k[�0���&�/�)�yʌ��:��&�Ѹ!S��q�(0�r���Vꆵ]IZ4�[f"&k�@W��[R�N���Y�u9���_'(GF	}\�k"������X���d2Q��2�JgX�@
�(�ShE�,0A�q	B(Z����$�E>t���,�,Q%�D�He%�	74ma����s��L
|�=��KI�����rY��%���Wk��޾B�<#R���Uq�8�P�S,�n|��+aJ�����c;����0���}P�ܖ�W�il�7�ge
��d;ılk4�"���5&ގ��|�KCxd$�T���Y��:��C�����]WtQ������qkyw��v�ˮ�=y[C{=A�ɇ<���/�	�z��tޱZ¶Y#W��"�%��t��'Z���;;F!)�ȿE��Du��Fg?��g��z�q��+{(êS}���>����q�2��g�U7�kf�6y������7��:0��zs��-�-6�3�Eϛu������4�sv�c_�w>� ��uRXF������Yw��n&�����v��95��P��3�>kO�_���;���-4��5�J��Z.��]�o���Ҙ��wY�X�%�ǇQ�@@�Ĭ����Gj����,gF��w�l�f��c�g��KF���Q�&Y���o2�[�.Xsy�>�F@���hz!�f�qG:��d
6���pw��9@�q�B�q3��+�S��=�c�.����bxQ���[$���s��x�o��/*{�/٨�.3W4�]yÖIp>��+�T��_�K����J�X�<��R����o!�u��O�'9��$�E!b��$r,�Ib�,Rr��R����g-��<��T}��G5���͂�ȿ0�a,�y� �ַ-����=s���U��N�Y��o��͕O.8�^�!k��{,M��$�q4WS�<������݌V�iɉ\�M'�ނL{Y�;x��2��"k�k�u������Dai_r��H%C����0��	9�6P�/�=�w�>�v�>���݇�boa��J��[�p����to�I�齯���;-/�]�8��(i�d�j�{�;H�����(xk��(����t���_�c������̵�s�26+��gKb�fyw	��+�o����TW_1Qw�n�Y�bׁE������c�h)�؋�_n)ר_gi2Ba�@�@�˟ ��w��󽦚ǩ����w�q�Z���gϸ��Pgc5"��K��W��c:#+�!����i�h��¨\u�&Oo@�E�X�|0��F0�Yn�����ߋ�w�O���\R��9�1,��{@�P�����@���L�5�	�o�c�������6��kX�� r�9:�py�c�+������V��e���[n��uD{�3��}��r_��!;"k��˛�9s?.^���WW(����VNJƊ��s^��e�ŬtZ�CR�F�R}�Kѱ��+��Q��m��8��O��xC�oriG#D=�5���g�J���;�l�wT/����R��]�|��WSGa"�*�j�d�eІTzE^�9��S��8V�66�{Lq��|:�N9K6ض�J��e�n5���0�=�f򑇕	�^�B��3׵2VbK>|^��^pC����j	�]:/��3v�3�����+:L��xм����zs��Sg[�o���)�:omJU�N��ҕ��52��tR�TK\ڐ�+/g6A��m�|v��I3�%K���m�7�r�Z��n��Ӣ��E�N�$�تB[;���u�0T��P9-DuX-U,�L\I-u�}�:�M��SxX���3ʷ��*�1Y"N���|�iA<}�؞d�r�����������A+��X�&ڒ�R��޼b��<���寍w�5N������F���X���>�R�瓚�[f���g�Z���U��Vv���cw/������#r��/�
E�wt�P��]�T���<�1Z;�O�ӕ����1��Cs���D��o/v�"�(�R};25 ����۲s�����,��QR��,��4uW�룋P��U��I%�O�08�d+_mB�{9��0��� �||لR�װ+Yam��?,W�I�����#�֍U��{�K;���H�Kv:c���7�/�ݠ����wǋ�0�Ð3��/V�e�Δ�v�[Ϫ�T�|�˷��n����f�dcU�6k%��|uo:ˬM��J����#Cu��;YU��],���Wuw���[����������U]�֊4
v&ᢦTݡM��s�Ӭ�S��5+�u��^<q��}B�Ʒ���u��%���4�r�B�ws�X���u���*�l�h�ҧ�/�s�Im��F�Z��n�\�Jm�uo�;�:�ZQ3���7Ӯ�@1ٻ�����ni5{w�w�f�����ښ��1m<��l��skE.�/����S�+9BuA|�]M�L��/�볹*�4�������%S˛�q�CCM鲺n�N��:oz�y��zax�mܝU7�+��:��j�mn>W-/E����/V��]]r=��p
eʱ�7���4�WEe�vnY�#ǳ��т�<����{�,\�0G��]��������]UQwP��W����Gd��BU�9qt��u�RDJ�qr�0�a�Z�`���h�U̢Ƞ���O�]:v������<}�^�q�}>��
�+�Ɋ�V ������*�U�e2Âi��%�>___]<}|v��c6=z��p8�`����E��Z�<j.!�Z� �1��X�If�u{��Uy��n�1���1���'g��e�r{�e~B����AE+
���e<�b��&و�UD"�B��Ϧ榦���S���1�ǯ^�㏳���K*Kd�U���,�PQ�B*<B���b0ҰI�1�y71��|x��1�����q����V)�%>�F"�Z�������2�QPVF3��ǎ��=v���c�����q�c�;��`��e����s
����6�(�)���(e��\Z�9���&	1[B�P��V��@i��=L_T��&�n�m�*
PH�c+*cU��4aU�VR�h��F=J�5e��I
�J�Pĩ��)FEe(6�-��6�hq�Y�/���rfP�9U�FK��E
��	9�]O�Do��T�7/_30��E��m�Z4�x�������X��X�#��P��D�B�I$}��Ͽ����*}}y����9�Hn2�@w�<D�sZDTqyCM�t��a����*Z����g���?}��>$6�I�dlx��ߔU�-�5[~�M^6+�	��ݑ�s���'a����� u��E�r���O�>6�Nr�a$_o>j� ����PH3fjc0�օ�3k�궉m9�'����!Q'	9c`pXA��i���h=�R_S�ןc����}�Ap�Ce�E�}���7p�����z#@$)�/��3{�gA���(��Csj�q���w�g�.Zȓ!��0��oG��g����@i����0Np����<��yz5��G� �p�.;�1�OB6v~�$�^@M(o&"�T�Ӊ�D��،���=��PQ�C������ز��e�B�ε_W�w�� v��oPx����~��I~���^>�G�&����].Zz!��v��ki��v�%��n9�sv�=�X'���3X���2D��s�me���h�{<�&���a-吙�-�b0�ZY�g�qKW:i$��5>	��Ʊ��B����Hl���t����'Y>`�:���*������_P��Gڭ;�i��Ω�l�E+�V�x� "��A��m�UW9��8����v�yw�7Vu$n̔�k��y�������}�}�����O�(Ib���:�I��[ZIȲ!2T!�$��|�|�����Jr?���a<�0���:t�~t=T�NOx��6�ÿ�Q�s�zކ����r;�#c�D>0*ތ^�/��)Jl�/�	��5����⤕���O])�xE���]��;���,��M|��� �Zxc�f��2����n;R: ����mz	]�E��P�9�%S��6_of�~��*�$|/�/��.A���T�)	L? �1�cC�G����J$�D�Ik�gQJ.�w��g�&3��!�������=�h��]�o1�`+�^?k��l����@���ތ��f�����{BQ���5���l8�,����e�&y��Dt���N�]}u{���y���i��YF�#�� aͬ��|� �S�g�vF���Z��+�۶f���;����G�sf������-q�5�-l��X58/���Bn�����<z���0�6�4'��"8�|;��=-�� n�����:��ҭ���o+����4�fc[�{X:W6[O6O���o���5�'"��ǔ���&�X�dcYm�.�� ���U ���ָM��d��r���םVmZ����qT��w[��+��aj���k�>I�(M�U�����̃1Ҍ�2-��������]&iVVT-+A�P�p��ڧY�R�����Dnr0J�z�d[y�p�����zy�8���A�<��w��A|��0a�uE�Q8�Θ"TdelUQ��%.7%�TQE��$���Ib��$�ȲNP�$R!%@�����2L�r+Ñ�zU����fVM�x�!'?H�}��M���g⭟��̗�&����&�l��svC��H�m��z׶u��a[1��o
��o4=<���c^c�ɱ����q��\ʡ�����upݩ�2��{��*6)�ڴk���l ��8I�!�K#�7�KG��"�1+�q��~1營SgE���W�=���U����.,�|Ԥ:n���K�ٌ��Q�,�Bg�1�)h�O�[�&x7]�s[^;�R���QG|L�0�@����T�f�}H���x�i5e����ƞ�0�f�n�]#�7D���!�$���as� =t�hѱ�`H�!�v�	�����t�ˇhv��Z[6
�g��D`u�����g`��{H]�>.p�T�̷-�r�5�2���q��=Ϳ'�����@Y���/ǻ���ίw��+?P����5��l��LD��k���"�1,�|7ӌ��ٳ�3�����B����\?z=kmr`*�c7���o��')wx�7,9�c���}�m���ӄjg��Oo}�~�]�$�6�H��0Cb��dXx,~M�{�i�XI>�����X�+�H�L��Z�:D�]�R܍2����Kإ\\�.�ۯ�]�L՟�h��(�g�r���U&xG���B��5Ig-�ܴ�+���vwfM��-�s����;o���p��$��0�u�r,�X�E��'����=��{ո������sO�w�jz��փ�ZC����z���Ov�	�c3�^|#��۔�t�C��ƀ���g���$z�s����\�yǽi�~<@���w�6ǲ���M�wT(���OܮNk����1�x
w� h`�Swy=S���>�n���h���k� {�kмvW7k�s�I�[�-�i���M�2D<]/�=a����)Ó�}���'����?l_
>UywHxB>�!񅃉����6ש��úX���<N<��U���R�'�݊D�;��܁g}_W�q�z��|��xG�Us��w�d�ﶂ��u�w�ͯ�p�t��C�zP)��O�'�o_,g���N=����]t����*%�n����γ߻?4��ͪ�V��遄#Gؾ��$�8��o�/8l%���IM�t���A��v[k�wq�)�c�<n&n׃	7E�0�^�<�f�ۚf��Z���%��~��
$��ݤ_����R�|�u��n�$�\�#kcr�!��ւ��ם����(O�+)��^�<mn�)���-v�oj�F�O{N.д*5��k`�������f�����OP�N�X�*��h���ս}8u)�J��vڣ�}d����L��̓1,೎������<��? �E�$�R|�$���,X�,T�9`�["@��2yO2��*�Ö.��O�\�;@�5��7f�ߗ
A��H$7�
�߱�nѳU��q�6���沎MR����*߮\�$��.�?��=ؘ�(��/���0F�!%5=�w[�Mv�,L{z�lǌ�_]�ޗz`+��ل���Bm�}׮M�4�wG:�_�{���ݞ��>�xM��y-��5AϾ�f�\�-��v}��7��9����Gx��  a0σ^H�����^,Ci�4Q�bs 4P3x�&e�[�o�t���2�h��*�Y�י[,A�-|�c l|C���o��w�+�����!��r4���6�gh���>ς�dN���顫�6���%��|�Wߗ`�W���g�^2S��r
��g�Rè�|����އ��v���@�։�3���q�"�F�t�"9�|�0޻��M��-2����,�
�{�"�|�=�0{���+Q����)�b����ӃC5Re"�M2�����!���
���몎�ڼ����=҅��}��,��Z4Z�=�& ���XDm�N���m�98�U7hmwF��]�<@�}y�����EG�M�S��X���b����mh���ss畓��i@Ї��4N�wy�3wh��;U{'!�;�7�6�V��#;�`	 {������I$�b$�d��$-%$!XI"�����sΘs}������9:�E�ర �^��� �AlӍ��}$>�Y]*���	�X=��b���~a0�/P�U>����Z2��MG�7{7�i�w��K�V-����	�#�AGV�`��|+�������];�>�VS�3�?j����Ŵ��=@b���%��h��<fk�i,����h`��3�3�%R�@�&�$3��sϔu�0��E��B[γ�j�T�v���Rj���'Ϣ�jh���'ܮ���g G��ŋ�/%�wsG-�֪�q9���[��c���Ol��^"F���bl���۱۽P!UC;���6�u�n-�B��th����0)����<{x�����x���(��S�P�Şl����Vw�����iU��C������k�cib@��.R�_�͘�1�Y	�^�lܦJ�� ���<�o݆�)�=>J)��d(��,CO�
]1���@�8�@a���
��ַPy�9m��:Df{��b}���|�[.	qȅ��_�0�l�&G?�
���wL�����=�x�l�jl^��Nf�x���Jթ�@��>������#���ê��o��gk�U�#MZzT�NaJ��)A"����m���W&:��9v,�&��;xju�j��i�u���59~s�-�-�յ�D�ҝ�R�Se�D�	H˂Dxd&DF� �J�����^�/� ���'rK�TI�$P�eH"I�H�@H���x{�T�l�z��uH6|X�>�ul��؜
M��t�E�P	�0��&퍅Y�;�r{I]Ņ{�����m�m�1�op�Տ�7Bٺ��
:��[�O�'�P�-q���	O�y�+U���y�iN��a�O��_70���K5���]5�� Fn��P;��ވ�]<��t�y��d.�˰rH2
}����M��67��}	5����>z�ܖ���l�vכ��s��{�<(����&��y��9�7�+=��[i���["�=�Rc�Ņ�h�[i�;�wa`��n�^���4�����C99�	�ܒ��i��sH�&����}J�1�q���͝@�>(.��,0� z>(��M����z��4j�8#c�Ƕ7cu"K�c��v`R�H�� 4˱=e�ٯsX0Is�,�5��cQ5��S�>�b��J��cϪ��������n���o	�M�7K��<�ȷ2$�o���������K�R�����4/W-���d��E�7}��k�L�~
�g����p!ǖ����jw� Ƃ˓�*�!�Am����-��R�ևg�qI$�A'u��p�fJ�{G�Hb��}����c��ˡ��MA֮��m���S0r˦%��暇,��L��'����=���9���I��B$BA# ��Ȳ$�>�!ȱ�I$�,y�����}ˡ���~��kfs�k�4����/Üq�2m�	�	}9m�2����k���I�����3�/j�
���/���rq�Q����.�8Y���W�Q����qE�!��yly5����/�Y
��m$�}��j��S尅�oO�z��t`:2^�S
��:I�k�.*�aq��h�s�_��c)T�������3�^�<��[ǯx�1�~P�B���}�F�7|�)����wն+g6�!��t�>�@˾DF�{�ʎt6D�^?IW�|���%��L�fr�M����>Kq��!��>e��p���'e�<���=�]��mZ�`��,�&���<D}ƺ�C�%V��
	o;�x����*��匳�������Z1ON��m����g���B5��v�����c$���k�M0���C��um��yz���9ԡ�j��ʆ\�»��(���(J0�OEH#��wM��� 8n��6i��ڟ
�[�њk�<;�Q�3����`dN2��M��k��`>��O� �"U�!�7��ܿ)�i�'uu�0�w�>����;0�!չ�t��G8��K3"b���&�S�C{�.�=���
�f��{s�����+F���򺳦�N;�N��I^�`j!��Y4h�.�;��+���s�ƻ.w5#���_8���"� $d��H�d�T9NJ"�	�
n�-�ql�o?��1�rj٩W�6��XG����0�D|���dm�}~1�/g0x1�<���� ���9~����C���΄�aޯP�s�m��M_G��e[�n�e�m�T�S�%��#�*�Rm}�a�.y��UD;L(�r��/L���T�bw��ݭ����y�m`촅�5kh7�g�H�o����q�+0��O'��uMJ���㝸�Ń3D7�A�̍ǔ���^�\\�ۉ������x��%��CS��X�Adw1;�K9�{���$�0B8�.�Ԟ�|���s:"c��#I=z^@>q�^�q���4��>��z��!�	�>BI$��^�p�z����{zE@�eӰ/z�ᦘ��I�淞`�]j�Z7�8kӁe��w������j}��p��{Okm���y����n"p�|��oD'�s���릖k.!�9�{̄���9�tq!��l�p;���M�e��fU�3Fx.��>%�Ɲ�C�+�����>#>W�����/_&����/�Y��E;�_?S�v��Muf�	l��(E��Ѧћ\���1+T�0;I\μw��!����^Cq[��Āf�g5u���P�S�<kR}һ��so��v[�&1�]1�V'q�+��iธB�Fv��!!�D��	)@H���a1a!�!H�0@ ������$x�Uu.���&3�ߏ�1��Drz8d����-!�?�@-{�1n�e̯��F*���밶"s�����૝s#��R*Bb����0x��X$�1ۖ�sG���o�z�{;ZX�Z1�dHC-6
<_]�zpy~>���u��^i����Q��F���;5��S�1a=�l�cٺc�B��|$�䣦?����P����i)pt3�Qd�oo�+;��H��ٚ�ɷ�
�p	�3�(��4��}Myw!����}Mn�<��+�u�����5!�Yg M�����_����L��Қ'�º��o�<������u�"���~@�^zƐ9����\��.�euu����<��%��!�ؖ7=Y��	}3�$�����0-�^��=���7�Oج��b���5��Ԃݜ�dt�7�À�a�;`o�{'�lE��UwnD���;ν�� �lz�0i��0�֑q�{��5_���$I�J��а�����Y1]e\8�H�q] o���n��N}l�A*T��ݙM��{���.n�ۇ��c+�e���F�6���<T.�ք��u��C��ו�8f�C�e��}�o=}��cm�{Mӆ)r����Y�Pߟw<[������2�i���n�w��ۖ-]��fgJ�b']��j��#�9VB��m.\ne�c_u�����.����k{-�%��y�6��z��d�{�_X���d���3(@��;�R�4���7�[rNuY�6�d��Rv�P���N�����d%�k��wSV���U}vL��2B`�@�㔭ر���sj�5{�5[7Z�gz�voLV%�i-ov���^V:d���%����E1n��[6�,�1U���Zt������{M��8�]/{UL��˜(�jf��>�����G\�G���`|��LV��﷑�FD ���׈������+�Vyry��xlk�qi��#�q3�5]��𴙿P��s���A��KU�B��6�.;�m�5��q���h;��".�뫆�V��>�2����0�Bc�G�@qb9t���u���V3��ً�Ѫ�w.��ir6�oF�u�72��Y�{"��8/�;���M����-T0���Zv��۳�6f��;!��e�C�z�!Q��Hd�t؍#�,K�R��`��g���.8U �f0BA�7J`*ݢ��"�rz�l`�'\�	wB��+�7���c����b9��Kc� w�3uO�Ue��>4���j�Xۣ��ta%FB���Iv�DKww|Q�P�܌i�3c�C5	�vl����)1�ٖ��T��c�;r�4p�O�e���lH���B�7�u ��I�MXvml��Mg�>��8�DNӣ�b7�bq!��[3Hw�X���{:��hL����X��(�b�`J�7�.B�gl�m��_yy��PN�f{�"7�մw�<��R�J`���W����o&oXq��t���@�!I�`љD^�����z.�Q<��	+Ѯ�V��k�9m�At�X�x઻̔�U��ӽ:0���i��T�Kz�En@�ڞ�̛=�,�q�ɅckQ��`�����<���V�e��l�;yզ4�[��(�=��]5���F��[�1�R��3k�G#P�{7�]u^nv��Q�7N��[odRe���	��j+ͥ�+8�[є���)���s��Z��v�gE�o
IOE�Wܘr���V
XA\��[��U
�G)w�g�p�׌�C*�n&FgV_Acp}"�����V8N6���"ywG����,�c�m���d��v��yoP�0"�)o����8plUi�C��j�6�cV}�Z|j�s�2��I1��PT��xi�V�{�����)�`��["�Y�7�'�J ����t4�D6D4dvn&�D�!(���(�7/��d>7��,��%p�����3\e�F�`�!��p��d��A� ��@��$�e$X22����cE�B�n��#��M��B꛻�Dq%�dƒ1��bT�č�j���� �@�Ț@��H��i����U*�T[��Za	A�!\�Fd��q�fR�j"��u�c0��c16R�MX�"���jjv��o��<lz�^��g���;���)���5p*ԩ�*�Ɍ=s�������K�ܳ'o��^<|cǱ��z�����s�Eb�`��ܹm�BĶ�n��2�L��V
�E�Ŷ�>�K:v�^<|cǱ��z�ټ����+R�V�ZP��Ҭ��T�r�����1�+x�Ǐ���Ǐ�c�=z�\W��x�b�*�^�B`¹xL����bzٴMaW-��ҡZ�X[e��ۧo��x��1�c^�����X�B�����F1Q��f6Q��VJ$�L2�Yճ׎:v��׏>1�{�W�+Ͼ��-�\l��8!�������¢���+�U�QQ-<f�ĬR��Q����+̴qb��(ؙi��J6ڕ��sմ�[X���TІ�TR�V��t�0���Y�d�e��.7z��["�m[�WZZ�UU6��3UV��P�r��7���T(�#F��Xѣh��X���㹦ɉ��zj���b׆��]M̱��E��t�{�ּ����9)'�TT"9���,�+�Z+{7M���1<� eu�T�񴄐��*@�@�@�!t\T(H�BS%NB	��8�!,Q�D��9%�	�P�P�O���I-�g,��|��ns�4U2R���2��$u@�O�<硨|�V=x��
,��yDMZ�V�^��w��b ̥���]���;���Kz���m	��81!��9�\WϽT_� �sm͹5/R�3���4vv�ϧ�/�1*ҝ��h-7�㡅З{��X��`щ[u�NF{M�^	�4�z8�5�>���.����n�:+�|l�1%����5S�����hncYú`��vz��|�5��3wy��Y����+�C�F�*���sxB뗭��}�s5�Ȯ�H��4%�si�{Ϯ�R��c�mc��O<�����N�@K����#�I'ż0u�s��`���E@��e?b�!�6M����Ad�=�Ar��h �<w�ya��X���>z7����k�I�:V���>���1 ߽owV�l���H߇q�ϫ6Q�|Љ@u��/�zD;_0�8�j)y�s׳͎w��t��=׍������k�u�P=�@���|+�&�dW)���0����=�A�5*�蛚�UO�MF�?;����fA:u�M��|mj�R�������@>����g�����s�F��_|��ET��+�E4ϐ "�b�gsڮ��q��쵫p���2�p����Q���O	=��Á�\���.��6�-�������a
D!X
#$�D�H�*HR[	� ,!����Ͽk��/�������.�_�{��8�M!cBH5��G0����
xɥ��Y��l�7D���?R���A��n����F����nԲi�'��=E�D�h��Iۅ���M1.�D��h�?�["�$oe9'�Y�n����(�Q��{Yr��T�is�5M�v�~��\�M��p��|�o9ڮ�������������1�9�q����\Pn�T(�S�X����#��,1�l�q��|`�p�{��Y	]����h�S�P=ܺ*��M���^i���i�&\@������d�"XIQ�K�WA�D�"&H�?Q�ϳrz��g��mJ�]�}|�)�v��R���~!ؽ�T���P�v�;�b&D�ꁕ�\����e�S@֎k�ѩ�?��J�tߍm�Y3I�1���:�Ci�@���h���%o<x��~�ڷ�sg6G�;��U�����AL�x���Լ�H�>d8u��k���zr��v�|bm�Zr_��L�>s&�j�u�[��w��KQ�ښ8�G'^Z�f&�L��r��i��(��d7z#S�;�ᬚ5�M���%Wk���\���ի���&�^�پ:jA�C;g9w�%Gq^p}{�F5�;ͭ���=��v�o�����o&��3��E����P�RIb�X�9d^G�%�ZH��Ϟ�_����~Y��=�߮�	`$���o�%���t��Ybo�@P�������-��lu}����T��	��.N�Ǝ�︖���nD0�נ�C"��,Ԟ�.���!�_+��s?s�l�Fa�7�V�.�Z��'�FBba�,G�L��w�VÙ�sFPL�k��ӎ ���I�l�}jj��}΁��b�����w
`���v<O���_M͆�vCZ�a�@������,��dh�?W��&�A�S�`9ͦ@my!X�w%��%#��QaO�Oyp�f��H�;Y��A��,�I�s/��4&��l��;w�s��+�KK�����TnuPUp/��^�yN�A�p��fr$�� ȁ'<�2��T��G0��@���Ԙw���'���V�3���g[���a��Aڀ`��������v5s뭜X�`�B�+ͭmCy[�s._����W��ｩ����];1��k�Z��/��an.^��X�$��os�0�}t�N5{z>�:�u����l;�[j��뇫���X���`�5��N<����0�ӕ��}m�@�+����,�y�f���WR��U��r�Z��㷶�P�Y��2��R��Q�\�6��D��z�#)^��}��_7%�~d��������[�bD���) � fK �2HMT�:��ѽ��;-a����7V32_�	�����Y�|��$H]P����S��R�:y-����B�@�m7��_�x�'�i�C�7=�y�=̥>g]�;��7e}���,l&m�ojBo�p|�[�xƵ��|#��:19�;�7�aӺ|������ٚ�۴�u���5ޭ����`���{q�hn����lx��~W���ݿb��ٸ��~�a�=D��c7Kdd$���5u&�3���5E�X��~�f�t�&ۃn^��#���*ߓ�u��6a�!'�Bb̌b_�K��W{�(���*/7���{�[��|�a��=�>�{��S�{�D(t��1�5��c�c�4^;$3��ضD��\�؎��d?���f����9̧}-��!��}���sL��{:�C	�$�ln�Y���<6����	�;c@n�?�T@��i���	
7C������S|��!~1��fd�8\��߰;%��	���p:��αA���s�� >���yr����f�eQ�s�q��X��Sf�eU7��������O<!�x�݀Ӭ9�X��F�7R�"���ŷ����p�A�2����ѥ{�c���X�:-����f����\N��\���c� �SN�R� ����"7��0��)$�D��L�@ZwR@���c-4���a���b�$�R9d��9R��$�#!1�"����wo�On��5�,�#�j$�� Ã���v�\��(�u����������%��LM�v��z�|�s��C��X���٩��X$,�F�}���-�K�-��d����P��r�Ϟ��<*j��C:=(0i�q�a��b�5T;�if��)�����5ۆ���!����Pjx1)�&Δ��M��	u���z�P�]Ӹ.�x�4�&&	3(�F����Ƽ���^�1`V�p|���<�mϗW�9�:���Q^<5=�
H8������"[D�^��1�U����ɇ/��6��*�<��B8k���$�*�Ş�L"��"<��֫=+��>.��qD�_2���S����-թz|���ɴ&��s�є�iK�\n����?��<�vJWϰ���&�Dc��yѽmK$��� _�׺�~�^�>�R�);1zӬ��Q��6�Ts��5=�x�̆�_��9/<ӻ��[�S�_��<��8I��f�����X�i��{�A���ҥ�Y<6�F���u,"�<2�q���(��=�5��=}�.�Y�k�)c��T��57Seem��kIv���n���犒��V9��X�;���vt���综m<ߜ��7y�e��B�HH�E�,T�9�NE�n|�?/������,np�������q�`i�����@ܷ�.#�z���0����s��e���B�q�ن�����
M���Վ/ĝ掺�Zhs��8���9������m&��ٌ��b{�6�D@v�h$8�t[��d{��d�y1���tc ��}$�{��c��x����I�8�6�1wUoj�u�K<����ִk�Ø��U���[��b�l�+�Ѥ@ǘ��/I����]ܸ.�3=#�9wv��Լ�xM��y�ټ�dA��]ؼ�����$i|쀶]������΋��������!��{���{��~�nf#l�I�S	��3|�{�*}������5@��7=udk|��i�+�D�.)�NlW;��t<G1����Y�Z�:�xN�q%��&����b�"�V#_s��5|5N{��4������L���I�3���j�Y�o�@��+�>|X)�^J<�3�RYҰk�Ú��n�ўwT�zWtU5W���*ݏl�G��'SWn{����伽�e<��r���j��'ݜ:�W��>�WC?eI�޾3�-��4�w��´�n=뿌��{?#0X�7ݤ<�};!=&���Z.�z�=X�Q��b���;sd��p�r>��,���i�=j�7��q-�$���aH�`R!P)	�R2k~s�9߯?	�����{|�}��� v��c_����J�TQ����Z����XFA����\~������y9��K�.+�л�L���]׵H��ԮFPU���N�����o*�r�����D�j4p«Y�>����� �� ;zF�N6�{��'Ð&���ś�6�pv�gv�4�3�Y�Z�#��	�	���ĐA[5�%���#�҉:�x,Gu�%�لv�b��ƀv=��� D.n�c�ь���_�9Cx���dN�'�Km�b��F��Ȏ��>����+э秱&��X�H�� ��'đ�u��a�����.ӁP�˵J�Y�q�ι���	2BG֔�I��a160��3�$b�L��s8��#��7P��yE��4��)^4�{o"�9����g�ꄷ���Y����D�Z7~�¼�
���o�U	��l��So�0hֿc:��z�>\SCT� <vM�����;�����Yv�������`�D���[�%!��>�:=��br87��3��]ow��H]����yTV����Na�d���-�\*Ԙk�;�0�\}�Y�J���[��y�d4�>}��t�^������ �K�_N>Ӷ��w) oOWe��U�ۗB�S8db�+���P�W��|(0�	2��$aQd��s]y���'�P2/"��u�q���>4�l������0�����>s�S۞֞���}���<{�>�6��4x�K��ϝ�5��~b���o�~͟u�	����3��F	�����#��c`,@t��cy����ܞ>�gj�˱�-F��o=��\��[�l���� >5sp�'_Y���gS+���(g��Kݰ��.Dz�;�!!{%,�z.�H^���or�E���s�^����uD	i�xM����=$�4��r-���e��J~��,ǰ�`�s�f�����j[�5>�H�|M<�{���p@��eK�o&U��r�T�=����[��[Y�����Ā��Xj/���%/XV>vF��/j��c����gZ���Þ}��G�����i�������ǈ.�x�����,4�Wv�9y�3�>�� Y�et�/N.��[�����j9	��l��9�G��M�Ɋ��uy��� 7�Ud��Ϛ�x�m3޷Kܤ/�Ta�NN�8"+�8�r뮼���1�8��N��(-�0]�2�ƅ
��L2��͢�.��'�/���r��}{�1*���7z�Ŗ�'-z:���@T�Hܧ�bAL,�|��a:BŇ� �{�Ԋ�ww��5f�V╘��£�:f�Z��r���]��]�jWq�:�5��F��B^���L�RlV�	T�m2�"RHC�ڒ$b���g�U�O� jRPĔ��FJ�$0(�DQE��y�5�{ߌ�^�dJ��Z!6�g����#��h*�Z��]�] ��=%N-z �����3���<A��.��>��N��_����G߈��zi;߈p��)����*��=�M��c�i����"���H-���I򆱇�L����-mO��Ŝ\�N0�����Ә,�$]�(�R���ݫ��^�6�p{� &���'������<�2|��⣂e�7S4�<��AA���4y��#E[<|�kej��b���rU�
������Bg���[�+��t��ĺ�03.�y���'�3O���,Dc�������`ǡ~;��o埼�(~�nW��f5����Ԣ?'�s�ap����M���mN���[+IɈzʸ�{�fd���`5�2D~q�Ns9�N�9��\�6|��o�k%�ݞ$�2��}��+B�E��D�$Q�y�0��Ϯ�S��^�~�X����UC�?}q01������L��b���ﱗ<g"��&���4��zfE����I�R-�q��X�Y0^P���S���V@���-�7�E�����ީ]�7t�������csm��(���Z�`���|8����!'�=p�oTh ��R;�rA��vΡcq�y�c���A̦3{Y� �d��T��#:����*��{rp����D�1#&�/�|}�[Y[�Żu��̈���^Q'��M�y4�Q邼��i����[�f@����:cr��t7���.����t0���HM<�W0�1t*l4��;��1��S����ʴ/�����ȣ��㰝h��x��z14�&
�f6w=�	�������I
�ׇCA���[��l7���} � ���}L8��ֳ͞{�N�:�}�Ə{�7]�ѝ!�S��XC`,a���S/��dt�Vl�s>|n|)��Vk�Ss}��^�i�ن�F1f3fY�9�I����L�y�>�oVV�4X��PH��sKeh��ˀ�#(��|���4e���y�	<�3���m�N�x���!�9��2��y#�]�t�#\����PS��mM���d��/̀e�m��d�b�hv
�ګ�--y���Ea\�I��SǞ��0�o�;�t�κ�WKK<U�R����[��X/,����痳�y1�n���?=*u��;I���v����~X�;^��bP�)rO6��3�mX:71��,��cT�S*�����$C|�fr/T`����|�#c8�����y
�gc�)Gsڥf�C:�v���z�{�,׼��
#���R�>�qvG ��o,E�gY]�j�^��f^S/,�>(�7/���V/��':^oT���#���Z�+� $� �hїm*$<Yp��y�<�.P�K�Dvl�k.N���RR�m��ZyVY���(�Q����X��߫Ap�f35���(gu��m�I��m�v�Z�^����1&w��"Rٿ
6�����2�*�V䰋�_.�tW%TT���9j��.�p�hD"��0Iy�5݃ժ1J��9��_lgF*�4�d툀3,@�:���(�j����H�n;�I��^�))R��r�%3���Xw��r)���{kرic���gnݡ�	�nD�֚��}��]$z�R���q�W�"J-�)T��k��^�2F�N��Sz���b�ȅ�����3�׷]+^��R��C2�s�hY2��H�˫�m��)"��Z�{"0��6� �w�s�V;�}�# u(sq�ЀW�;m�eb}NP;H���,�7bOUuo��@��]�xY�Ԇ�!F�S3�h�)w%b�HQ���
�i�7v��H�������-"�2��̝"��g%���4��]D	
6�!D!��K$�E��z ,��>ЃK�й���|��~(՜}�0��H�H�Wd}$\k��>p��D��d[�X|.�QS̺f�(T߶O/����+jΑ,���`��x�^t�������b�S�-qe�3l�۱��bf����ut�o%�T4�ݠf(%�\%��N��>Gk��h`gKw[����|볓��ݰ��.�����ހѠOv�\1�]n�^`�\tYDB�7������滹�m�
��m�����"�8	2S/��`;�T�jf�m�����=�N���[ۙ�G�`��OF�N���L�����N
�m�/��V��2�$�
����YVV»�� ������.��[�Ze�c��`��Ɨb�9*`����)gQ���Y�i��M=�r�ή�D�w������]��)K{m���+3���!� �x�Շ�)\���-�W�tE.�n�lPWp��/V�Ʋ�-�9E��l�g2���R͂U� �gU�ǣq����+�2��
W���wW�%ru�īokG[����&+aV�۸l���Ţ!wf`h�����b�՗ۙ [�}s�]aͩ-��ͦwo) MЈ� UFbլn���Zֲ���N8�T[kӓSSO�x��ccת��n��圷�-hQV��ܮ
�޲t������"i*��aE�J�<���^�x��c���q[��o�H�`��Z��L�Q�j���E�;a�E"�VbTQ���N��z��Ǐ�c�U{�->k"˼���r��Y���̦+4°��݅L�(������N��z�����1���U^������b�G3"0�*Z���Tw�b��F#��ɓSs������y<�N��c>��ĩ�6��m8���0��Ec���e��(-���5�E%�E�rdɩ��������y<�'���}>�Q~~ʌb(bT� f8Uo)�鲪�7JV6���iA*�g!D񻴊����c�A���ys*�EV%�UCyY�]e*���&�E��Jͦ(����F��jcid�Ln�FzՃR���f7fb5P�ә
�0�"*c-K�y��DE���cU���&w7CX1��G�]��w��Íܾ.8m�����1���J]����8���"	-)Z��H��H1x�L>�Ks|����8�cM�k�'%S�����C�ϟ�6��Up�v����_�i�Df�3@ֆj>)����2�/P$�v�O#��qs����:�3��ev�;ݮS쨃ҕș�2q���+�YS	Q���ש
�6~ Oj��G��S���ӛ��sM[ ���uP9tݵ�=pg5l�6��x�`(�gn���-�w/s:�Ⱥ��H@��A�-z�\�o�*�υ&Wε�sY� u�
�:�ϯ��;0�n�¯����4-��]�w�\z��N~]��]��ڟ�>S��v73����3��q�u#DHœz���X:�7"C_�1}��9�Ҏg
�|X�����#����{c�̧D��k��z�l�uJ�E���l�1�44���z&�W8� gd�&���K���t)���I�v���<�����0wk٨�L&�3�ɮX3F��y�^r�g][������Y����F��������b_�'���(��+���dn��K�vD0rs��5�;	坺T��EM�}!����Z�y�<}��rwa��b
�}�/��1�#�v^�+i�"[j�wV�V���]�f�{�s��.�-�wv��܋��oG��p���#��G�H�e �o���������2 ��ѭ=��R-6����K{ha�lG)�vC#I�!���3���g(���v���k���H�r6s_���'�}ޝZ�~�b����vwX=3�9�{�z $��s����ˌ��>K7�4�U$�U]|� ����P�:NظU,Z�S���e�`x��*J����{��}0��!@�;�G0L�9�6�������/���o,l�Y�r�f��'�\3=��pY?s9�aj��i�w��4yV>�]oģ������W��{Dw���~�Ϸ��\�F��z;�r���J��}]��e�KY�i���џl^2�����b�AE�n9p����BʆvA�Hv9p�=�x���yR�o���x_n�^�St��3��f�-���`�$��G�ΦIT��Ә��]���U��:g���ׅ�Cr��}r�i��N�����Vy��^�kC�ԥ@�l��>��f7C����bԄ8��ގ̥��E�?}]�ݱ3�wkT�������^�E�K�:+d#�W��[q����SԤW�[;��UpK�cs��c�5�mn(n�f3�9]�@��D�.���=���j�]��:[�l]�\l�[�M<�D��%	���q��IԔq�L�8f�����b�%"�0[Q�
�*SRI�����(��R���F$eaH�D��^PX����ߪ�'H�e�=��f)�ۘ��]�ZL�K�<oƃ�A��5;�^/��,v�EUr��д��2;�;/Ǥ.����]l'��GHb�ӫ
M����k��Pp}�-��'��=ܠV7s�ON�$r,����_.gQ?h c��dC�obn�3?%�S��7l�����3�S
�$��ͩ�XV'��M�'	9����R��Y��0p-�0�~�wl�r��������T6a&�4|*�����5��a
�xNoI�& ��=4��haW��F�oj���vq����n0��]b`�!Oױ}�Yg#�{�Y"j�� ���:���ϤP���Oeĺ�9O�����f�w7z熕��y}�Ϻ�����B�m7�`��a�^�kBg�]3ܝ=�3C�t��}��@`Y�mn8�?�:=��<$hl�r��6�	�5��u���͌�{�wS62g�SP�&9Ohj�f�;�n�f��$7���O)w�Zj�d`S�������1k�u\E����[
G�q�ܛi�N1�Nؗc�L�o�����$��{�	�W/D�?�<a�x3��T>�ݝ�a����9�SS-�960E��s�m�[��~"�/"�/��E�g"�� `I�$U+��2�>���8[�鏡�*�V�~\���og1axC#t�G����W��x�5�D��H{��\Lns�����b�6CKTλŭP�":;�G��T77Y��)�L�`[ٳ#����ͳ	��"�������ˍ8s��xo*�u��� �j��P��{K��yMn#ӑ;�j�7�r̆ĝ��_?nZymn��[��*�r����/�W�[׼��M�f�q�cc��tz}��]�P��o@��*�r_�m�oMg|��Յ^�x�$Pᛯ�
��0vT����K��C�6�ۊ}U���֣I�Rɽ�G0��~|y��ٽ�~��f2��R����ʼ���ݦx@hD��B����hz}�w>��W�o�ˇh���g\o�2�ݍ���K�h�f$����u����,���/_,��\��ڸf���Ά�=����������֠=�v�����N�k�ڿ3���]'��{O���Ԏ� r�S����ɮ��w���*U�L��Aq{����t��5���7bOp��&�y��{�=����F�[
FQ�A%�<X��-l-�y-��5�b��n�G����L59`|��^q�
&��V������{��������@���k[8���qp��6���j���h�n��O�F[0'�������`�h'm�g-�9�:j�X����.�&�:�g��m2@a;�;C��芭�5:y����Y{�՚�)P5����»��_���y��ߺ��� �j�,"��ìl͞�v2fи����^y�0�51]����p18���[S��Y.6��j{b�"=�/�ٍ�O��t[��do����7�3nz�7���~M����K�?t�,\}U2�����5���@ۺ�J�-�/vz"{�ݓ�鼡��|�}��v{��;���w&��lFN[�=J�.����N��\{�����U-]�d��llY�g�ֶ�}�����
�m�O�y=�Kd=�T'hK��d�T������ʛV������,����c��%��TB�ͻ��wt�sՄr��a�n��_mvY5���&��:�b{�-��1���X�%wL	c�Μo�BK�g�~��p��b�ď�n�YQ�i�7�8*��E� ��qNa������o+uD�7����8��읶 ���q��3�<�M�.9��z���kyb,>���K�F6�"w����%o[��>���U��������u����3����C	t����;�wޜ	i��A/:��v����i��Ό�N�ԟ���.^v9t�)�8��Jv+|�zE�d��Wf��$4�hc�����ؗ�a�螵�t�}:gY����9K9D��q(H�v��f�˟@\�+=qU��lE�x��|L��YƼ�7���`�*\鉹-�'��Q��[�� i�v�ȝ~d����Lo>����1+���Qp�Wy�=��U���a+nW�Kz�w�E����c6��v����WO���GY�><sD�T��?T�Ф��8񙣐�y,�Jg+n�s�qȺ��ee���=�A7�3ֽ}ʿy\�Âg��w01:�$�/	HP �J��ȯ�ݐ�ǖe���*I�{a��j���]tv�ji�օe�壩�-�Ϋ��b�h ̉�Ars*R��l�I&�e
f�l��l���b07 f~q~!"E"VR%i;I�)���֌w&�}��϶(�D�EI	��ɶ��~WMp9�욟y��VnQmy�]��ɖte-Ü�<F�T�w03���y3��c�F���q��h�^f��3C����K7!���@@�M>Euz3=��f��O���ڪ�6*�d,���}P�M@k��5Py����T7[���o�*"�c����ܪ�9('�s���p:�5D�8 �!���D�	��Z��������L�Vo6�e���lvnllw.���y�ŀۍ���j0�<c���5���9�WxE���a$��kX�k��w�Y��p����k�cXv�Y��]k1�{���m�G�F�� $Ԅ[ʂ��<A�c mV���~�N����d�V�pAS�c��[����ݯ_G���>�ށ.��*(3���xY��D#�CWN7�졉��z��#���j��vy��ڵ���L(z�G�
�>ϗX땽qc��x�xeڹ��1���,�r�:��ع��G�{#� ���
֚'y�:<ŷ}o�]�����g67�������`�M�L��8�p�]���X��L��{�;��=�U�h4�$D�Xx�a�<�>'+&]̷��4��pِ23��{ [���U���ϸ����������fOf���:�0vU��_xk���Z渫���os���Gv�Rj�g����UMZ��P�޾O��;�h��Iie��hls�{�r�)����r�􅉿W��/o_�7�f�=k���ȴT_/Pg��Q4���BgiV�ڧ5��ȶ�7,�<Oud�C`��94�����D׻y�z�9�"f�j�b`��_3�5>�I.|ğ31��Wl���\�����i�d��?��tND�˰�:���gc�׵��	�Qʫ�wQ�D�$~�#z&{w���olrP�=�Ys���H�	[	�c�q���1-�;:��+]y�}^S����m��ך���`c�ygpX�����8�	<s}=��(�^��<�T"C�T]�j�t�m�Ny�՛�6P���Wf5��IR���çh�y!י�k.���_�~~�����\��.��&b�'K��5�v�Wڤ�0s��'R�u,�w*�,��_[���=�� GD!��8a��a�����X��.| ���|H3lޠ����>��a{>:D{��͹���l�������V��c���=�}n�a��9��x� �hr������[����ӕeg3��e9�1s��/l������yO�1�6-_G�ߢ6��$���=�����{�_ӄm�'߹W�I�[��;rw�s�<�{;���)�OYn$$m���@�[s�d�K�o��v6 ��S�Cv+��ݩR��9�n&Nkҷ7כ����%���w�N��q�Vf�"]d���5,57n�
���Kֲ���_	��k�^}�D�,���:��3_A�Ԩ�B(�@�>.��u~J����Ny�z!lhU�r��{��������z�v��4g��D	y�|ߨJ��&���.9[4e\6�C���X�����n�����<��`�F�q^�h��y�0?e?ک7L]�tR>�
�z_~�A|h�nKbvvIR��}����͠�]b�qg*5ھ��F���fkOQ"���o=]/_P�:}+n�L��97��΂�3K;�u�J���xY�PVFgo/3���s?�g�ZD*R $�a�`���$ H�}k+W(�o�P�h|�[��?��~���!2w���V�6GR����%�ׂ�y�'���v��SI?.�P $��{;�e��f�9�A'L�/�E�-��L�#!8���zQ�x��	��^pqG�s�=�\J���I���h<ܫox�݇�K���5~s������"�4v���d�ىvk��E`��l]X��ݽn���z�ǃ�_�pTV�l��3�ޖ��/�r6&��c�y�A��(.��>��ܪ<������p+�eD�Y���-�*"*���巼27��;CbqJn2�l|��.r��Ȏ��T0,g�5Ō��~��.qKՒ��}�O�����sy˧1���q�X���
�{�ٱ"c�8S��'-\���:S�*��;����vg�SO�O?�*ٮ���`~N-;��W���xx�Vpɡ�k���6�.�ȉ�[QF.v���������5l\�R�=��M�y,������w�r�7�blک��N
����0k��ئ�j�[ʘ����hǯR/d|3����:j�qa�a�/�'��'�v�ʺٸ7V�ɝ�HY��9�U�$V@�n��$4hL�V�*]hU�՗N�A��Ωp���V�^��WDD|�Mlɖ�4�N��*��7�	��i佷b7�W Ҙ�x(�^���
���GA��xX'e�P%�HoE]���|�X����T9��a����*�9���ئ�K�Փz�q��(,��/z饙D]�&he�]*U�V�f��L-erc:����EF���Ε��/d-���e�뷝�Drz��ǖ�r�,ob���qmZ�/��	T�ʢ�T2�5�,�m�Z�s�@���9n�In�N�k^K*��q����כ���>X���#u�E:��9�mM�\Ϻc�m��vF�E�n�0Ґ�J�-��]%�c0}��釲�N��^+�W2p��u�D�f���.D�%�{�V���W[ދls]�e2s��CL:n�O`Un�6/�n�Va�TR����Ȑ�}N��{�ve�@��#�c�ɗM,�������[j�5�k�~35�AEvMi�b] �+��m�-�d颺x�n���C"G,b�2�̱��HP�ۦ������_c��,�H�A�;hKK�-s&���wH8�)�r?+�lm)�ܸ�:�t�)n�=�Hsz�[����֋��WTP��{���kw�v�����D����n�&h+�29Z1�P�RF�ee:v//�΍��G��"m.�V���C�F�vc�2��n�1�ޕsO!y�1t�۵6���}���{OU������Q]h�,�ʄd=r���Q��[.�o��{!օ:��o>Y7b��1e�H�Wb�̬�9��[�N��g���o_�� �v&�ޥ�<y�ہ2�;���0�cΣ�C%�Q�h�55V�w	E�l�M�>"�C�,G�s��lu�D������x���=�o���f{rv�4�p�1j�V��aA¯vO	Q�鰧|�ԍjpD�k��E�|(t/�};��tK��Y��`��I�N�utm�d�*�]�`�X��K5�{d�:B�*���)�;��ۢ)�7"�^�w�tcqRM���5��W�v�=��M��v�ھ5}Fq����#9���ٯ�\c6��jO�Y��z�*���'�*g�M��O4Εg/wG+v*�(H�͛���{+pI��֠�ݯM��]6���{U�9ʓ1��b��yҠ�*�Q����6��۴z�����v�Fh"�b�4ȶ.��O;Vn�� ȔR6P&\1�DDM$[E@�N0�iAm�Ԍ[\�FX,6�-5J@�b
E�*.�!bk�$�V�?IH�&��~-R�5t9�������b�L�-���E1���L�EF�1Ѧ���̗
��lGDT��ӧM�nHiB�P',D�(��n
�Q�ێ(��j�-��&�q4.-ˆf��Ģ�E�[E�&-*����R�jba�rնԩEX �ӓS&���Ǐ>1�c^��kھ󓜜�'%�֌����4f9K�Ur���DV6�b��1��u���cǯ^<x��}�^��l�P���3(������!qb��6
)�fAƢ,�K�`�l���e��|t��ǯ^<x��lz�1�N�(��(ѵF�A�UkPcKc���TbV�nZ��v�ӷ�]�v���^��v�Եu�2���b�E�[
�][���ˈ��DP�r""(����UUN�QD�}�'��������nrp�O�Ӽh��m�kQQeIZ2�*��6�¥[b��QYl��c��2̞O'�SSSSɹ����F3�=�L�R��ūD�*��Z�6�J!Y[*i�!�#u.��#R�A6�r�W)c�mb�Kj�F#m*�e1�m��A�F�QJ��媉��LD��VV�-���X҂�b(�e��"<�kBf�1���ۍ��yu��*��eU�U-�T�b�D�cF�1d��F���$_��L�	�4�k� cm��<wN����ae��-��mom(/�2Nb��$�nN
�㮕�X�]�;�2_e�u��*�7>�u�6]:HGV�<�ES��qGF�TK�"Q�n�[�h�:��H��-
K�0� �f+H�0Qַ��wϱw���y��O�"Ei`���}����Q-.^�V��y٪O�;�C6���\�bkv� { �ƚ!4�B�GZ�aG�wd��~��ܛ�r�Nt��\���l�� ���kpg]�qY�bz��D��Zjۥg$cJ=�a��\V�/�&�<ץ��a[�7{7�;��w��c�5{����D��a����AJ}�p�Nq��&�5�PS[}�	l�{G{+�ݒ����>K����e{�r�**��)�k�f�k�7��������5>�=�HI	��t?V@�>i��ؖfO X���������2mV��57��mP�U�K��!�c���x��N7��>�c��U��7��bX0b,�,|^��^y���{Q���Sv���NԹ�Ϝ|�b��]��z2z�nrKR/{���֎�t����s��pнh�߃��c���G���fZ��ʳ��4uLƱ���w�ޥ���r�Oq��:J*R�]
��a�+y����c�v�$&������D1��2�3f�Z$7!��f�:�+l>�O�k��0H�4�FX�}�߷��߻��;�7��{�N�ά�����8�0*�onʶe��Ԙ|ת�9p=O6m�}�"�����|���ҳ*�,���z�]��μ���w�{���%��;��ޞ���b����f��E��' ���q[*�}���9���:�ʣs���[U�%fs�&9�S
F��Q{�p�n���)o>�	4/4����Lm����O'Xا�F���n���ݞ�1<t���h�&B��������LU?������E{a��M��i��,w�q�|i��=�Kֻ,�g�FtZݢ�\Ƃ��e�gCc6z�ٜ��@�Z{��yô�>�^�"L��jz�;kn�3G2.��\��\�n��p�v�i��nJ��Z��#r�;T��ܳ$�WI�ɸwk8�:X�4Gޡ�r 5
��&��P��гv+�����ys2�c+YK��q���z�};��ؽ3�N$Y�wL&Un�.ïv�����T�2X�UqԘ����Ә\V��Z	�¯j��G���#u�(Lk�==�M)<A1��V��]i*�W�=�J$D����7Vf��~������>Y{��j��ߩ�0v�3.n\&��#�Z�՗]ٜӑ~������=��G�mM/?u��u� vA�5�����V+MO'�(75��pa��	�,L��O����Ξξ�;˧�;}r�.�SMs�)Om��jr�?���{\'�I��}!�0�\�w�O-do6?��fcYV�վ]K�[	�QM�Zl�R�յWƘ?n}�y�ج�hΝ��B��6]�S�J���nb2�ު���@Y�z��d(��>�����gk�-�Q Y��H���~պSyI��81{�u�A�s{��t�\s�Ϟ�m���ۺ	]<�Z��-���f�q��ːk�彼��8k�ש�{����7�ij��x�=6<�^km�ݍ����@�]n�-���	��۹�}��D�P;�6	8��{mh$�g� nwwe��%�u���&�v��P]�]tݬ̃N�mG���y��{���՚�����O:Pen煤 ��!��%�$g��K8���3����<���[��|���Չ�����b�P�����J��l���w��'�<����@oM�-�\;�83����������>Ļlwv
s�8���=tE�x�t�po�7��I44�7��Ў�>F���
d��A�W�㹝���4��j���R���`"��	O��6Jq�Jw�2��<�<LLnG>�C�}c/��.����(g��ȨJ���ML
�2��U�����>���B�҆=��͛����w�v�h:���Vc�'��ո�Ɲ���8#P.�-�w�Yxʄ�O.�v����8�<�nvD<�*�KUFY������������T:{'c�C�^m�ԣ��q�3^D��>h����������D_���1.oea��8J2��tU�^n�;7��ϷFp?Q��(Ť1}��Y�$��@��ukRC�$���^�h�^�o:�� ��IޑC�����C�+3���{��e�ܡ!�q��ӫ`��rL��M[�M�i�F"4U��}6n�qM��um>�����aN M*ʡf��v���a>(���E<홸�zno����W��ڦmft�ڋ�]�,VYǪ;�٤�Vo��Q!!�`��K��	AT1�e�@�� �<@���-ul�O�}�t��-�����k�|�wz2;�n�F+�� �_�G�6/*'�ME�xZcU9{��F�b�La��$ZΉ���z�I#�2�n��騖���Z�Ѯ������*]���^�/_��0�X5+���R_/"g9�+��{}��NEqpg��N��
�����?h<L��Ƌ�˲ط���pAp*�l�XD�s�^Î��
 +$����St,�mVݹ��h�C�����s���ߚ�����[�u�vT,w�ܶ�4x��-�D_]��b���~�v��<&����\5M.�.k��-+n�Ƶ���O�|��A�v���V��K��as�_����%g�=�W/� E�@˼j]�����Oq�,�V۲�U�.�2;��������U����n�A���]���Yl���Ռ�$j˻�nB���U�M�t��B�Av��/���b�i;�.�O��kp:��5��Yr�p@t=;�������]�0rX��R���(�ʷ��s�ac���i�&������jn���$�k����&�)L���D�j\�<���:���r��x��q����]�yk�X[`��ﭷ�G[^��+���g�n�OW�y}4��ظ[���ϗ]��z�s�>uoz���u�X��r�ϻ���NwY�د���n��E�D��D�|#ϼ�^e��c|:_on��M���ĺ����ّ��\����F�X�x譃؝B�.��ۻ7k�$.!�z�(���7���U�K�\7U>��h������@Ε��
�Z�����s����0�r�6[�d��l�V㼗x��+�؍���n��D4-�wc�׹-LӤv�A����_����O��Ng��J��-���W0<�z�^�^}ct�][錽��.��k�i܇�����zߤY�ې�%���,Rv�٫hu����SC�T�F�Y�w'�#H�Ӄ��[�F���:��=�
��j�_�(ց��޺���.�j<��{���Ü�]���2��k��z0�i��`�"�M�����3c4A:il�{gJ�w�1N��o�ph��;L��k�e17��D ��t�97p��E�N=���)���@񙙜����ә������OT\aCCT�3��^��Aܐ��r�vi�:�9�lz��M�	��=b�cy���j5��DG],Zy�Ny�I��=祜!L*�|ﾈ��u0��8̴��nn^n�+��)������(̃�>�w��G�*��������>fk3������2 TBA㜨�����u�\�����\�'�ų�+)@m� 3��ݨ[�T����U�;
�0`i��K�=�d� �j�d�f/�����z�oL�l��W�+��R=5WQ���	�!������i琽!�g���/�h�yM����_��v0Eո���U��q�r1(��Ӑh�u`���؟�sռ\_i'���&����)�Kr�+��u)�1��`�\?48e�wk�=b���;�)���}���T�%�i;xW)x-Tv���7��eozOd�C��ѽwd�+|��w\Gn��N":�It'P��I��t��N��m`�}2h�H�/ ���?1�WJr��Ҙ������U篝W	ك���	!�&*�!n�ۜ:9���Y���Ӕ���B9boS�6]�sň�2��\5����wW��Wzox��ۯf��|nEϲ�goF�U���v܈��^;xx l�b�d�o/S��V���nG{ˮ������$������5P��������O{�C�g���b6-�^���%���~� ������o.9yg��2A��2��޿)�z��缦��^�Ҫb�r��nt|���ޫE$Y��|GC�c�guN���:�2w�d��=ˡ��VLnm@*;�V��Zyr"��7������h�c�+�n>�1�s�xY ���x�{ָ���{�g�(јI�6����V��s���<�u�I����ș;�����,�̋�a럦,�,�Ѱ�����-��n���ԣ��Lum-H��~a��z�����I�ys](��d񂮳�Gm��b�as3v�W����u��DB����![���h|}��GR�2�\_XƦC��k�r�Z�Wg�bڙ}&W��b@U����rktV�pK�-:����wax�m�"R-q��)r��W���X�N򚻻n��)����(b���Ͼׯp���!K1�%����g�^�u�B���iT��ȉwv��95�xz]TfOfA������z�u��w^cHˋ�~�Ԣ��R�T���uƬ���ͱU[�����-pGTя�����0{�m��n����&׋f&1������̎�F��Ek|��n�.��yX��j~���U�+[W��T���w�q��_����\�Od$���O�mR��H���Q��j�O�<��';f�������3nǠ[Є�7�st�?�mzP;y����g��ﻷ�n<�8�v�bK�x�|���0��@?����@��8�F,-0aӓ�z������*��u�ޓi������=��y߷<��f-l�ew�6'��+H�#u�d��6�*y�Y�f\J����9��V�0�}�� k�����c��Vכ���L��j>���ɸɑ�ۊ���SDM��5���\���,5&M�駫�"�f�x7�lǖ(����x8�ļT�,���/�*��N|�]��C9�acM�[2�����W�C�n�]�I�x�=����[	Bk-�:<��椮��hο,ݢ�l㖹�T�r���c_w�
���r_חj�������^��f��'�����y�ukq��\�O�����Or_k��}�a`kەِ��͠�3�UC:�=��C?��k�@��w>�-O8ÙÊ�N��0��皆�ޯ)ھ���rSܫgp����T�2�mʖ��ڈ;ujk���$���C6yR���gD�y*G{M�7S���ث$ڱL����DAI6!"�X�Y�vbC"�\�ȷ�	��F���l��0�]���TM'ɧJԦ��2��\���ś�K=��YyWO���x�i|�="f��.g^i�spݓا��5���lu���#͗m�U���o3L\KNI�@[����'\���@�̀+�������$��=�4��܊��`K=�����aؕ�J{�Ý��Y6���|�s��	VV��5g�X�����u[�C���v*YjU��%�H��soӧ��s*�#;�*�O��SW��L�ĵ(C+/�����vې��NJ�aM�°�Su�&����b}��n�ˮ�`סT��fڼ�:
�gk']t�x�d�G'��L��[�����a-���l}�|at���ɪo6���W��tueLa����t����g�g�Ճ�ڦ�m�ٴg�M���\�9 �K(4� �5��RqK��B���o'^oU�K}\%+��!���h*�2��d����t���F9�X�:pR���m�]985��R����κ��A$"��(Fq����I>�6�%kkF�L�����%B��{��r��/�aՠ�C�r*&�]څ�u�� q��Ɗ(��.�*���}�kHW:T���^���v���Ƕ!�}Z�{�_�+2�D3����S�l�Ҩ�e�玱k�����P��r���H�Usf��Twt,ݤ�vl�W/�/��n��p:SX���)��>��<�9GNv�BƋ����!9���$�E hBZ<���Y��w�B�).�l��{=�|��k)]�Y��י��F�wTj�L "�}�o&�(�h�J�n�^fY��_T�,*V(d��KgWY�s�{�u]mQ*�e��J��*������xZK�5��s����W�b�T(Ex-����,GVr���1O��U��b/Q(g���K�{�RQ�,�Df�Kf�d��u�e���7��R��.�Ƙ���4�J賚;��Y�}���74=p2��M��8ݯ���iҏu���J�\Q�~.���M���<�̵�H�Y%�m��_J�O��2莺m��{55�HAN�c�3`N�X�Rд��+%�R۬m\Uoה�˖�@C�'W�:��u������댭�-|@��'`�f�P�e��0�F+�
���l�f�Հޓ�:��a�wM���Y*k4�ᏸkG٘��w����ƈ����'_V�շ���7z�J�8Ti,b=]�ˢM*N�tWhmV��DW-˘��X�U,�}%R�2e�7ע:�q�/�*�ք�ɘ���r�V�e']��-4	x]��u;Zt���ts���M>����啰�7[�ev�����Y9��.���j�윛����#�Fvc�6�i��&j�9f��V��x�[��OfE��1y�z9�:E�0ZC&-H��B�j�i\��7�_r�4���"�R�(�����Tr�X�D���#n3Ϧ�2jnn}55555<����c8R0� 2��*�B���Y���鍨�YMVʶ�Ֆ��5�t��Ǯݻv�[�c8q�mR�(�P��ZV�1�׭�P�W�,�fb:�:t���v��ǯU]n��2�Z����E��X�Z�ձQQU�bQ�%PE5�q�Ǐ]�v��ǯUZڲ�Db�=KYN��f&d�i["�Tc-�QV��r���;v��nݻcױ��V�ь�kR�(���[6�=ްMZ���� ,DE�Y�T]^χ�c�nݻc��ת��,�<�&}�b�����kBȣ9J��ŋ���&�� ��J�pl�(V���E/Ԩ��J�Ѭ��}�b��
�1
�jF ��KJ�#"��EV��T�t�ٔ��SWQE=�m4�R���c�x�elb����e�y�{�o�����`�G�te�z�W��t�q8Z�I��kzN�Wձ�ܗ��.^�Vq��~s��9�),������߮�r5?��_���,w��5�q�s7S^�y�����/����ﱹ�Ӱ���ݏp���X:B���Zд�WC�#lN��;�oN;fzѰ�rf��l�%3=rj�ĩ�|̵��Jq+���W��*���R��;�߫x2�7\���ZKwdb��h@��`�JBD�I [$���+�Z��F��aH40�I�#s��Q-3�ك-<;Z]�k��@��>�ӽE[0 *�B6��� )��(�S�<�$J@�c
n�t�0���zZ�y;��1���i�m�*�測��s�d�r�Ă(O��_�T���SK膘�Ob�&���D
��Z�ԛ����IuϦ@���;\MT3�f$eg�6:a���U[�:�vu�j�[��lZ'!Gwz��~��G���-����͕.m���\4�]�a����t�a�K+J��kBP��zARJ`+z61jX��������UÇ4�����l�w[�K��W����[�p��;�E�鵢H+o�����۽ُqo1���G�#�>DԉӚ�p�{��q(\S���b�o-�	Ou_�<�E�V��]�V#��.�1�W�$���G{�q8ϻ�;��\�cY��^�Bp����r�e3��&��$�č�D"�����|e���ԭ�a��:�+{|��.h�2���t؞�;��ˤ2��'ܭՖY�9#�
���O�v�5�\i��_w�JU��m�	�7�O,u)/FY��ds=��5���M;�i��{�kWtk	ˈ�@��j�
�}��/��[�T��f�֎�4*7��IF	���7��o��z��'�z�e�C��ez����g>h<l���[��z��NO���[�nt�ykw����d�f��K����"���8�K�;�Ek�����p��3��������9��Ag]�jL21�� �7��Ƶ�>�!����7���U?�j�J�,~�cGw�f�iu�a�m�m��,��lJ��(Лݙz�U<����X��-cm���b�be�r�ȁY���pC�d��.^�4�	�7�*�P �ΤZ78R�{�e�#K���S)%e(z��6��v4G��Yڠ�tL�.l����ﵵ)�m+2�Q�k1b&�m�wN�q��2Z��#��4�28૭�U}x�]�o�P�DY�3F�@;/��Z�>$��Th���O���z;m��"w�u#���������wȎ�\�5"+U$o�*-���<=&S��י���Ս�|}P>���霗���ٍ��j�:�ٯu�&cg)^RiO\w�S��EQ[�c�p���.���]_���wU�����O.��sC˼��gG0v<[����GhC�~뗊���<Yl��F�C$T���m�X4޽�<����<��{��t�,�=V����[�_��ڹ�t���v;�Z6q�??�_Jz���z���;/���A�$�^ǭ��י��ۜ�s��u�F!T7)B�h�l��@.n,H����]��ȇO�Z���c���O��s3�� ���K*j�l����F��䊿/pϢ5�9�gr�3�/y]ŭ>�bc�^��q�&�Tb�f 3Ν~����9��/�(y씽��vt�צR/tc�쫩lW(U= rU�{"����@�j�L��v����1Au5�}�3k;m��^wv��J�3�e��N�f��P*���$x�<A.��V��� �@wn�\jRkپ����^.>���̀u�g�%�V����GZ�ٮ�ҥ�mok�^�N�gbkد�7oiK��2�f�5�[���:ґ���۰����b��/t�]�x�|��b��2V����%��r�����ǁpo�G�}4�������|�w������pm�L�J%�mk��,2�Yݰz�x�G���Yzr9E����7��w�;��S4��n<k<��^���,�����sl@9��/��Os��JrG)�B���v�ϝ�Uq���G�c��������є��K2O��}��ɵ�]%���Z����8g��S�9����F�M<@۔��+���O�+ʧVwL/E�]l����
�I̛�p��f{?R��I�SW��v���M����"P�Wz���Z����Ñ�Ƿ��iR��,������޼�3e�Ȫ�	7t��۫�Lӝ*=�Z
�<�x��t�v�\^4��g���x�S� ��q�֣��u�f� ���Ymr37t��F�ݫ���C]�uw@�*[�I�#�� H�H��7,��ȋ�|�}��PN����u���꫈�@ך��n-T&7o5���ܚ����y�#u��^��;[��|G.��j���
1O:�9�`����f�"�=)�����9FD��������Z��V���sJT�����h�1nkk��+���i��gbH�ϭeaN�����k-�,5�$L���o�C�}��!2tb�w��Cy��;���.��������r����vT�ɨn��*��"�1��/�6wY�73[7�}��7���m+�f�AF���c{���s��L����?�����{��9B��O(�K_���Ǌ��v���ă�o-K;h�^g�A�G��/a��jW�'��6Y�9�Q�y���׻���C�.���3�{�[ɉ��ޖ����\�ȇ�p�z��ʢյ��Ilq��D���`������9�<�,S��̫o�B�"��N��5yb{ڬx��J���}��YnmD�xH易1�ƪ�|� �v�/ۻ�3��=�KO�4ם�֞���W2�-P�zh�K���;-���|@�#�{�#{�5F�*�I˂�=�b[6C>;�ߺ$5w���ސ�/+^^)R��=�7�;�7�t��f�/=0�;����-��Cm���]��ˌ���歉�"��n�S��ވpY����oM��3W�v���TX�G�2`U������d}�'ar��� �� ����x�o"�]��h�w����^y_�,c�"/�櫞�qNj	G.{[�`��J��������ȴ���ݑ���N4Ĵ��c�*����JrB�/���|�B��.�/��M63u�#t�R�T3�u�hܼZ����aa9pǲ9���V�2HG�m��P��BI��iD��t�Da� �E�}sd�~P�$��d�؎�z[��iޗ ��C���3W���s�=ym�i��_���nI�(�����bm[84��ֺ�mEU�F�v�tH:ۊ�Ǥ��*��o�n�^3�ǂB�U�3�v|�
B�`"%&�������Y�|��d }�Y_���ٹ[P��7����	����ev�{��v+إfR��H�$5�����CvH��*�BB��Bm0���� j�t����
�S��s�8e\��|2�w�#��T�qO��hnd����\��^T8[�lYNP*�o��y��ўT j���8#�c�ȂA�y��ܵt�о�ŋk�ֻ�7����T��_�E`<�c��79!�tz�l����s��c�-1����k�[f׈���hcs��-��h�ӖgR߳����?���9g�E�U^�F���Mw!"�3k9����m�����S=��]lT4�����I�Y?zg�`L���h�� µ?�"�%Eƹ�G"��Y��w՛�3�:k�n������k����-����)	\�������L*؜�m#�� ��yq����2��o<�x[<nMvzF�c�[�]U��6+i�gw&?�p]�3���;��L���<hx�qI{k4W3ZY�8�e� N�����9M6�Ő)��5��`�.8K�3˧"mʗ�ڹ��2�#����*��F�{a�l��!�s�|3x�����{){��4��V�$��9ŧݙ�x�u�;��S����;��8�o_
N�$�9�	p+{ײy]���9\���>dx�wןg9��|/��k������O�z��p�b���-Vw6�7��܎���s$�A�b]�u�ڝ�>����lLo=�7ws���4cV+���ڝ��{^W_���Gty��=��{Fw�+;'�i9E�tNv�U�ǲw�\�,uv�{.�Fv�zi(n��,�2SO,��h,"}�g�vP�@���tS�\�H ��j�c��t��٭���JR�ʿE�o����j��U���A�G�� �A>�{(i�f����7��t�r�[��5�+�s;��+�Z���ځ��[a��F���s�V_~�3���9���P��bm�Щ�]�ћ[���Aqw��M�ZJ5�Y�{��"�ƥ�	Π!,#98ܒ��[/t��l�E��-��H�m�N�������ɯ�^B�V^ku얫
rn^���wrI�u���3�P���}F_��]�ߺ�}��cY���*���{u���tދ�Y�!��!�W�~�V�1�*���ߺ�g;��{���}��{lKT�m=E>�ٿZ�p�O�6ݢ
̊n�\�����^���=�x��9YP�6(x�{ڤ�9���c^u@}��L�z�3ʏ��k��Ŏ�n���7m�;O��!eׯ5�5N��<?7��8�F<P��}چ1v�l�����{�{H	�3�3�LJ���=�fnj�b���)&��8ٚ-�U_�[���@�\�%G@]UzZ��{3���{['H���O���߷�������"4�f �}���8�>�q�oo���ʮ\�2@����壐u��u���_@�^~��oX���B����3�'�7��m��t��Զ&r;��z�\x���h4s�'h�N�>���c9�ӲSIYR�Fo4
9̗F)�?�Di1d
oes1�^�rk��q�.aB2k��C=F�ԅ�ƁIl�!]�ʺA��p]����=X��X�c^�3�S]����z;c�
��u/z%ӍۮM�d��s0�$��i�?<Q�V�/Ge\
�p*��k{-��`;�Jp��.����O�K��v'x>w��fVJ�w��y�w����v5Q�f��o\�u/}`�]6;���򺶫h'�ۼ���ٛ���(Z�l���f����g�F�iK�Q�g��Z���[���2FiICR����/X-�g��]U>��F���m�V�|��z���{A,���~��}��kj2���T8�������G�cRp}��m�}��[�Ճ=:7e�9]]&�B� �p�s�Klc���`T������g�)OH���"�SF�͡cU�'2����%z�w�]I�˴C�T����o�!�������]��Q�-ncSW�1�wI�WT�ѼoR���,�L1?�P^��
B��j� �\L^��<��/L2)�[�"��?���SMc�c�ݨ�S�w`A\�:��k����Un�A�w�Z{a���L�p3ά���.Ym�в�������6�n7gs �������H3-i�]݋��g��]�����NEM�|�w'�ω׶����%k(ItnG�$+�1��e��^�'���/;��ĴE�`�f4��"��Y�����K�U�\+n�	{3��oeɱ�ٮPAf ��u�'X:ZfƸ�;�G/v2��h������N涤nDO;�����`�ky�u;o�s��h ����ά�[�FL}�}@tJ�K�w��s�Jr��}ʖ����]ź�nQ5�*��˥3�/�y�e�WQ]�.�J�6�Xs���﷫ј���1�B����M3kV6�յLi�r.�J����4�r��%J`V�������c��K�K�'%�y��+报�et��� ��v���]7�u5k�3ۍQiݫ��-Of�"*�tFܑ&ʝC3�JU�7Ϭ��U�V�GY�n���g%�{jf;��A۠�:,��ے���e]�!˳�a����U�8l(ժ�=;��z�a8�X�v�թ��B��Wb\U���RM�v`<��ǽ�anx�.�!g�}�v��D)�Y���혥n8�r>����qZ������ڪ�5�N�m��눻v�>�"`7}�V��QcZ��A�(,P���ťF��pT�D��2p��Tw+[��Rh�w�Tm��A���_�Xr!-��p۝Y)��i�"�4)*53�l���:���!;eԸl�Yv)G�T�K����-Rm;Ld�%⪼v��bP��i�n��f��J��m�{RR�U�.²QiZ����m�AMCZ7l��Fb�N��LTp��n@lcG��[.�����m�|K4%��X��Dx�<���!���Щ��'%��L���G`�P���.�|�V��h*)m��J��b�v�Q8��zeUѦ2�
ƚ�R0�>�p��#YABJ�d�`�=�w.�@��Ʃ���҉�ۘE��yLQ>\͟T�h#"���=ܿv֚�z��v����*�n�F�5��qs�-��a��}6�w���	35Z+�٨#0�J�����f%�z65�:����0d�h۵ӴL�C��ݕ�Ww�DY������ڷ��;6`�q�u�LVX�vkk�N�ع
h7Qګ:��X[�#��/V�b��1K<֎�U��N�+n�([2Ͱ��8[Y���o�e�Y6g=4fbg^'�	�qm���ķ����s�2�o��x���voڻ��`�H�}��Fg�є��Il��d��P[�i��eł�$���^\�%��h��%.���5�]*뭎rw|�kZɌ��-W*@{L��l_l)r�c�ɾ�q�gZ�p�������nc��Y+�Һ�R��n��FoV�ab�C2cvrJ��]�U���7��8��g�.�fQ;+$�����R��f���=�	�})b=-a�a�o%���u�W�Y�Á�L�`|j����m�iH���S��@U�m8��L�J��'0�f�J�l8,�.��R�"R^JEq �N"���U�R@X.T!AQ,�h��B �	H�dƂ�F���2�E���Q)�`Em��pB"D)�\
4�0�(&5H�.�	].&�eEm���A6��:P,A!M���D4��&��hL����f�QZ��-��DEEk1r�Ѿn�҈��9l?6�N�<|v�۷l~Oc�z��6�����?$ҭ|q\���Z���E"���K->aC��,ɹ��v�۷lz����>��-�N%uʈʙs1��=�������������5�y>&L���MMMMMO''��}�C�1�eJ��.[(���-�AF�mQURל�J����t��Ǯݻv�������:^��X(��"塍1�I�QV����CGV�J"#���N��۷n�ǯU[�l�,;�"�G)EU�-*���L���"�X�*�����dɩ��������{>'���w�-V,[j �C�Z���\�J�6�J��E��q�N�1E]%F��U�}$���3"bY�����c}$3TH���J�� ��aE�jTZZ�̺��ՖصLn<LD�J�Q�q*������*�l�_-`����HW�&�E�Ħ�����%D�ēh�*��u���
��`;bq���c�dW������;���3�ץ�4�����.�bZ��]l�܍�$e��F2�q6���*�	!a��������G�Tr["b������ �]������Q�Z�.�� ���Oy	��MS�s��0ԭI2�s�KOxf����oKE�y.��]�E��b����s8�?q���}��:�^����#o"ys�6�x��%�-������c���� �OQ�٪hK�Pڽ�2m���!�G\l�y�Uk��nی�#�� c'��<۬ؼ�ݐm�Q����s�5���S츊݆�!:p�#�dZ�a�Tgŀ�cw��|�a�� $��USEpgk�o;�7%c㜁�s�[>2�GՏk��r�!(���y� >|�Q'��9�e���`r��7�c���.i>{��u��}�MW��=�P9,��JmzZ��t��:��4b$�9�y�?�+�?�+��q���k�P7|q@g���]֗�6�uW�=��72Nڶ�E��0�p�o ���1���u��z�Z�;��n8��/|ۣvg�#wQOc'%�LT�d�|���Y�]��v&E4���W�:�{n�X
&�`���  P�y�A�J�ƫ%�����[\�{���V���"�Nd=��p=�;�N��y{���{a��*oy����!���7���uz(_�^��@wVQx:H�yy��F�w~�$y����îA����X����Mmj�ڂ�^7�N�������Q��M���{@#&�̓q$K��,kSRg��Q=J�#��f�z�l	��t���Q-Cn����=e������xɞc7-�	��%��m�.qZDp�+}�ԫ$-�;9޶p���pkh<�Q�Uh-�wPh7>���~V2;6usyFwn����6i��\���+�(��=Uy��mY|!6���}�c��&o:�q]�;�^��蛼㋤�mL��x�x�e�҆w����7����Fwl@>�t�شH����vf���̀��~�Yf/�]�1)|Ί~v��u�Mvj���x��I�j�6Rޭ��r��>��J��l�%SX�9�fz�(��;����ʾ��y}L�,V���I�6v��hy���~ۣ�T'���Vݫ���JGB�4(�f�/yɋ�M�kh����9�1
j�����`��f���7��%����:���qWr��6p��H��J���J{�}pV�N�Z���7ddތ ��۵�Wv��$�,�ӯ�����5H�p'z怸��p��=��[�vV�����}q���L2yއ���@ e�	��]�;<��6��jxa��-�U�yqw�q���i���b�Q�/�ݣ0OPq ��8;�L�^K��_Z����C�P�E��gS>f��q�u6[��;ͮ�݃����;rn�mf6)���8X�l�Ӑ�$޻�b*vY���O6�c���-�I4��o���wt�@R�
�fnh���~g�t���V���3��~��X�٧�WG�{E*�:Gm����x�0�K�;�4�k�����5�*�s�	�������-�?]ϡ&���؛��� �1HCd������x���eyf�w�xx7p�-���ȉ�l���8���"�r���xfӔ��E�D������t�C8���q��MD7�/�]r�.�����5��m>�:����-��Jodv�����Jby/�bn__=�e��_ <��x���ִ?���u�N���b��k�^F=��i�V�U�d�#y+�8��-͆�k��3@�n�X�.�r;j�]b�6�����dd�ʨ�aI��n� �J�;Wԕ�B.�>g�,G����\-�Em�{�jN��s�/��{���ι%$AH�wּ�ط$��Dr�_��:6��l6#U�ղ��������.'7v7�GG+��h8��������c&ffff3oXiU�R���o=�A$��e��s3Z�co��>�����av�Fn���s���eO>�	 ����7'��{}ײ�R,n_w��K�d5��_R�<R�����72�֩h:O��v7��h�i��l�ќ���a<4�6ͼ�Ǆ����ocL	R�P�|$�å=� �x�^���)d��%� �T��$g*���F���8�n�b�ᴹ�O�-��֏k�A^����Ӵ�a��u�f���#a)��6fB�m�B�2�$��4E��aĵ<t�dm�L����L��Ş�⼄%����ջ��G#r�o�'�2��76�1Zv�jd�Ɯ�"�C�a��1��2�n��[w��F����Q�
ejܦ�;������n��f�߮�)zA�j�Uݠu�TW���-dc��
l�����|�h�m9�o88_]�TV>�$��z��U��o�{|�z!^ln�%��J����|��Z��H���9S�$���&�M�㭷r�5�x��J�l�>�n)|Ϲ��ո�̟0)���u���ŧN�>U+�:7��CH�e}�]��|��K�7k`Kp�+�]�:Z����+vz�3u���p�����,;v�H^	k�Ẋf�[;���q4�W����N�=OfǄ��"u�zY*/K��cJ��a�z]�g&k�;h�u�F?�w���.ʽ|��R�)�o%O��,�D�\*��4�fh����`@uE&CA��$fD��gnx)_�}�=Q�����MS�=8��O;֍<�k"p�ֳ$��Q�y*7�)�-NFq:��M�(���'��x��vM(AKY��N_�d�k&d�꛷-�­u��c�����h��Vd���#.�*��+ĶM���k��j�S]������lc.�N����S�^7��̅�j!���.���쟔��űl[s;��|��|����v]�U��p3�XU�ag���>l\�z�-���lkP�"8%�}@�� �q�6�y@��X��l1�m݄���L�=�$͌���WO����5h��3��Z3��(�i}{+�{�j��}��*7���T��
��nVH|���ң�.��`�וQ��A��fL��F3�]M�ɗ��ˊ�N;R��ۇ�/�"s�%��<l$�#�tY֑�(�U���GAO(�D���ʺ���t�O'`���j�Sd�I�'A �hۼ�6���]W�[M��:�ȓ�8��4V�KS0a�,y�kVk��#���=�U��YT�*���Qb.�5�w��0������9Y���	�z{�{'ݱ����Ir�ٹ�ܫ+�)gg{�ݯy5qr�Z!ܱ}ܟ��u�m���׹���]�ِ�Bg#&2�9�Ul/g�+�y��B\�\�2����|��.�*����+ӎ��hodI��th�=�u"7:����L���:v ��8�k��m^r�w��5+x��:�Հ��;����5A���Ds뛻�>|�.>x��uj���g���\	�ڌ,�d�vLn��ݥ�ݦ���}��`���\���#뇦ت��Us�~X�c��\�FؒѶG܏F٫^��kx_=�⏭7��o�߄7^ܬ�6'���mim�(%���~��	c��`o������/��l��n��~gɾ����&�	����ߥҤm������>댋��/,��^<�љ�_���R=0:�P��ˉ����zv��1d��SC	K&�a���z;)��.󺘰��*d���*4^Kg��}�=΍ZK�!�MVÙ����:B�.��ڭ�=�g�!��[:5��R:�T�刕�g��`vY�ZDy���f=��Fvr5��!����ԕ���Y���KP�CK8�q�N��iT��C�۪j9qw#�Up��ŷ d�)μs%�Q�|���$��Ż��9�������w�Xw�4�HpI�'�?gt���'OeIs��Ӽ�|�rQܻ���w�#V_p[���A�ky.�Z�D����0��e�?��#����*r��U�h�vZc�Z��bx�	Z��L��35��ϲ�`������M��$a��M��{^���i�R�f�J���}F=�4��M+�z�\�P����U��3�径�A)lG�m]Ou���5�9�?y��]r�~���NN�z;2Fj�.OǙ�&��xI�:Ю�E���dc!uS>���q�	k� �F_.�k�6b��O����]��J��<�:�7nM2gjv�~�R='������f� �Y5b��;���0�nk��Sy������a��<\�d�Td����+����df�@��v�̛�����l��=��Ѽ^��to$�l�I&�;ㆽ��D�w��] /�~��j��T�GT4�_K\�.���z`އ۸DOt����YX�b��<�v��}l˴�Ո�ҷ�-��t�P�Um�����ss�a!1��{s�Q^�Z;i�{��)<Z��@ˢ&w�řV�%Z��2��W�$�F櫨l��M���4Ws����8�i�#UT�x�q�o�
�6���B�4W�@��~�����G��L�V�ۮY���e�����`�v5X���$��a��n\ۍ�pT<�u0=0�#ꨒTS��$"�%(H�B���q!��(� b��EJ0~�G9�s����L��,�~���ԃAړ
ǋ�߸j���oiV>,�[] P����h�%S�DJ����M�Cz�=�ϤdU?��h\��co�J����*�����7#t�p��H5�9�v
�3�(�����g�U����v��=����l���7�뢑o`�|�<&�V��Y��)؍i�=��0N�^7��sY�5:��ojT	�.�!��s�k�<R�����}�^�ΐܟC4������-����Ԏ|[S�n�-�5������"_әT��ܲ�ed�12��'�uT��Gci
���Ī���퐣��[��j�5 [��=��M���VW����55�Vzb��A�塣"r���%�ݍV�l��cK���4d�� �b�ٛ\���DriP�[�Iw������C�\��S���'&+=��h��+[ͩ�:]v��e���7��}�J��AW���`���Ǳ3Q��=s8UX��N��M�>t��{���jƎo�qSN;��C�!��,X��q�p�N6��{H�#�@�U�6w_a:��L�V>8�w����߻��{s�HM����U<�y�ܽ�q���f�O�-{��uʜp ��}�s�΄�si�B�_K�y�b�Ff�U���&�_l��>9���YQ�f���-�}�k�c�:��d]{vv̈�6A��K[9z�u�zn=}��p���C̽�F74�+��N;*i-����O�1ź�g��"pK��`f�[��h��Q���?�:����*����.��xFs�Xp�l���?]��ǻ�����t��V�ƑH����W��O���19�����vJ��0.^�\��e$`7�D�]���3n:0"�^��7!�Y��lЗ1���<@����u��5@�Q�ʎ2k�k�eE��z^�!t��)�P�Ωn������AOz2@ѩ�L�p�����$6�7��y��|�XVr�/����6�%tidߦӃ`����8�Y�%k&�n��n�Y7r^�Zʝ݉Lf4�ܫZwV�Igc�{���VE6�,tKɽ�X�?9���>{�Y�MiF*W=8���V�B�q�s3���� �SNHk/y����V����1aГ0_7Ү�nP�R�!�ث���oH�LmT��Ws.t��܏3���̰m� �K��}R�n�ko��}L�DM�q{7�(%�]���ۭu�%��Y�>��
�q؆�#�H��H�^y����<F�-d�Dоw�L�*��P������.�v"��L�:�\�6NԺ`ћ�]�V������+L'k5��\�&_w*�ػ!�-��YZ=m��k{�f�3���I�P��oz�)B	�me��lh3���0F��MK@Α��as�LvRa�9�-�F]ť�Sq������4LWU$"�s]4r��{��R�#e�Ps�]�e�T�'�v��U�|�=㧯OK�.��me��IW�"n���jfP��ԥs���Y�s�<���,�B)��k+�T�������ަ�r�8K �ʒn�g.X%ɛpǇ������=�<�3�̌��P�m.\V�n��Z�]����Ӈ�X �`�Y�ȐJ��`�Jծ�&
�
#T5G�#a�W��2�7r�z�vU�[��c���ޣZ5ݍ�B��ОTV7�\�|X�������	��W�^�G�!��SQ��R��Qyh|zvؗ���6��qAYA���d�ږ(Uө�V�C�ci>O� m�'��+^��vu�
���K��Z��&l;����v�n�#�U�e�ޙ��^!^�����V�o�[�k����]t���ٛ�gs�۲v��O���Hs��wД���X���{_%�aC��۪pԵp�z�,"<[��B(㵮^-ܽF]D�h��U�g8��c�)aTs��Sk4剓���1��}'n���t�;�\Z؆��)��kI�d���N��ӕe�+���C9��K1�=�4]��$T�^�@��۶|Ofrg��Y��f�l\&����Z��s{�r��[�0a�;��m��Ě�of�HhV��V�t(f�ģ�,�*\T��]>X�b�k���� چ��ف.����f�&�o*���-�w��M����z�v�l�O�E��Z,�h�ړͷ�t㆔����=5�y�F-n5��,%im��,��Kmg���J����r�Hcm�Iv�YS,�����漉 E���-�Q����A��M���(��B�R&�8MMM;;v�۶�5�lz���l�m]㓶�(��QE�,��,Tƍ�L�DKJ+��2d���jjjjj}=�K�>�辽C��mH�̿dҎ%F""����`�\f$Q`/w�4��Y��*3N&���f�����'���|O����#i�_�i�L��UWƨ���KiP�h\�gg��d���njjjj}=��3�}8O{(��u*���c>j$U��T�"������+���v�۷���+�����Y�P�(��ĬE�Q��WV�����A�v S�^�WO�v�۷�_\q��f�*�'���!X�ZZ1���KiQr� cE���*��>R�0v
�J��e�3(QO]`Q�S�V,v��KI��@X�����eh��.(U��9�K�1V"��UUU���U�u�E���EDU�"I �}
x�1��,���Cx����������{I,�R�F�����tl�f�eS��7�'�f�Ȯ) <�5�h�/��5VgP�]ѱ@.�y��y<����nx�D�m��S;��.
����_HF�}��)O@ꭏoKS�<6�`�?n�e���
�ȱ�3'Qw�����z�S��s�޼t;zk"�Æ��˻��b.�:l)��t�n�Y�]�3�7Mp�m�US����U{�	v�"I(�3_���G��,k�`}�s���1�q0b�£2�*�s������װ#+���P��8�f1���7QwL�b�)`�w���^X ��o{ow�B���Y�绡�S[W
~D�����t>�ݺ#u����Rt�(���m��eg6��+Tfr'y��=�J�����u�]�-ؓ�����[��D�n2�H@�_�o;���6�r�L*(bDW���sq�����I&ނ�}��ܓ��Y��mF9w���s9���ǋkZ���sp�rף�yU�<�uh���
}�VGc0��4��S;�8�p(�Nao�ޣ�xn�=��o�)��c���<|lW���fD(���ܞM< �$�u�z�M	`&L��r���܊Z�s�`�;oW'/ӜtUc��*������"���c���'��
n���w��m��]�'�>��qk��d��1�EX�A��<{s��Fv	FjL�,��{��=������E$�n&�
9�r��{�F��z�Zķm�]�%�^��9�.꩖WG���=��Sǝ�z�ō	G*��!�ٚ|�K�u�s�>[�/}<�2c��z1���=nq��!� �P�������	���Y>�={vG?b����۰���H2�0l>��*=��ݳ�`��ȗ�0_��������\���u[�?H�w�n����[<= �ܵs��Yj<_��}P��؎L>K�m��j��%��6���۰��2T:��C��Qo�nf���Y�V[,e����7Y�I��'A�ɭ~�8-W\gJ���m�=3��;�U��<4�WME��`otX�IR��V���L��v-����gw��V�ֹ�gesiܭ�tr�w����U�_cToi�o_v�%�"B�������hUuA�x��0��IR1!�T�a$�6��p�-T�q¨�i9!��s�G�*�|���v����h/�0�xᑮ1 ��~���/��cٴ�m��6��10"H܁��Q�F*`-�{�3�;�R�~�w��V��>މ�)���-�[�N�rg%�=�n���)n�ɟFs{+eշS�䱟���0��K��69C&�͵��_V��kM�����X�������ް/�f��q=�\�������Vkt��7������>�m�nQfU��#�%�縡�"��U�:
|�v���1T��lc�pYz�[����CY�B<�zf�u�x� ���Ws�>��~�U0��n0^ϙ�Z8Ԉ�N�]\�u��h�^���T*�,������X�"�j��T3&�ݳ�t�u{���8D�l���hΦ��Ar��Ͷt8�z��3��ތ�.Wu�>���4i�.z\�L{!��d�߻`/�/]��o�溞U���y�;Uhn�����Ԋwy�ĨL�ʧ);������U��/rY��r>�}�hӜ���K��2��]q̹�dgb=�vE�)I�ac�K�<��	n<�˪�:�T����X�G�<�� �=��6�b��b�a{9]L��Gz؋Q'z0o�I�)�Xv/�s�����$�7ĞݘS��W�����5k��"]����밺-� yy��+�����\ח�k�6#�vw(�
4�"!`^��=��������Ǡ8��#k�Wz��팝����Y�k��m]f#-W*��6u�6�v�k�jdGz6�'x����Wo�'fL��/|�
��uN�4"t3�zÙd�m���������ej�����So	��ㄊ��K6��4}O��2�T$��ٿ�����0���=}���ڟR��J4�����͕pղ��ůS�9}~om;0-��� ���|:Uщ
бN��n��5.�����Y����,U[`+�G_�2�CS�lV^�Z͍]��ۘ ��4y��G�4����I��1�7Tϱ9^��B��m+~�`�oB0������^(�+�&Ÿ5�$�{$��Q�#/��;�s$!S����tb���YXT���m�9�/7�}��)��^�5ڸ#�%�����l�����^�X���q <G����1KS���/l�I�w�����=3˅	����J%k߰a1+�~��9}w]��]�[Z|M �ng�v��!⦅M��W
'��^�;31tJ�f����Y��=;�
�N�;�zESwA��w���՛5�Qu��6;n��ʧ�!k�j��h���Q������WO�e�@��%�I���e����`$�KH��I�f�C�bS����WKT��}Ys�<Z����۪JH<������Godg�0�D^�@fι��ȗڨ���d���x�JhucF���|�!{Suխ�n����v,ҹ��w��:ۻzm0/��'���l����u�Ǭ����j�+�1wf������Y�H٘�[R��͐rr<i��|�+�>��Ł�}���ƣ\����j[:6[!��*�����Y���\E�O�fp�b8b{�f~��|s-��N��e��Sz�<q{;Ԓ��/���Z}��[��	z3�3[o�<� �	- 4��6�������4����m��Fr�^��-�:�z˚hl��tJ���{�{v�H��v�����=�xe��6�]D0��]k�z�m�ǔ��N��{Cko��ɚ��K�T�Em�{�i�p���o�ر��=>�OL�� o�\a�:�s����^fN�w[v%����X��f$�w�QJ��W[�{�j.�k����h�+r�r͵�5���+��ǜr��uez�
psl��k���1ҙf���
�\P��9��P
(Aފ�/�e�W�Ԉ��z7Q����g��l��8灰$�m]�鉨���t�E��������&�vH���ݒ���m���F�o�`]cD��gǁJ�$+yG=]h9����u��V�y���;6fz�6Gf�%S�~n�Sc�`DM.�`��T���d+��QrX#t;h������l`mF��ǨӆY�\ޘ����
�~Y]ҟ�yER�Q�`�D7�����N���4����!k�TK~Ɔ���{�Wq�$��5��-��y�瓴���̈́MO�KUxY;em(5�Ս�9t��>F�p��$�U�tQS${����E�o^2ȃ�.��Q��g���z?,��7&������ ��8M�K(4$��1���m�!A�~s�G�9,ـ����}����Sap��g���ke?ʣ��[P�\Sz��M��l[-�v$��w2��"��P���>�V��>�j���A�o�L#���}C{!,�����Z��g-�섵fr�] ?܋���jv� :�˖{\���6�>i}��{�����n+�6�l���6뜖��;����W�ʹ�Mtvh�G.Ⱦ����ɭz:*���ղ��Q s�����w燽��[ӯ^+X_E��Rf��m�b�,������~��}b+�C�#:np�_��zl͜��ʇ`��7c�:_�m�"��+���}�}����ڭ��1�����]�F�tN���i��v�B�(�JH|x7�m���w���1��f�Q�řNè��wMOngݿ5�p}pV����"�[`VAg��3��ϯim�D���=G>�|w�ws���t
�;�yۥ��$��aM﹍+{�[��Lqryx��+��]���x rk��1���r���ca[`<�/�t�х4o�Д��C�R%���&��qrs-�����_�� =�u��Շ�#�M����>h�`v ȓ�w�hĚ�m��n�����/|d|r�&
��?�䞹�_�_of�$Ǚvsk��~��Z�����-�[&��﫰�=-�M����>�ѵb�f�O���P�l"b�S�In8�A���\� �}�U-��GOK�_W�>�~k���%U�%s����dۢ�K�E��vm?n����ە+7��Y��P5W���P&.����Oi.���<௷��d�c������@��=��}@n��^��GgoG���+�ؒ�d���˗�|b�0��>�v͔+�1��f�����>����l�K����م�6���ڼd�S\�ɶ�ex�%���#Ӡwo�����]с���ǥ���T�9��LY`o�3��������bsb�R�du�33���j�o68� 9��"���] ��O'f0y��J�����I);�7�G��#�}�a��z�"�=O&��co0;05 �}>xt���&���7&0��z�3�%��6t���؝��8 �2�(:��4r�q�y���w�[����bp��L�����w��t��$��\�b�lW�7j=3����c���p�p�^�7P��}��K���ۛ��$Y`}�5H���
ʁp
N��c(����rnֿE�&�n�;��)MI�����7-���UG�4�B�>5 �i��F������d�C�y��Z�d��zGW�?�G�^�cp}}]6�nq.�P�x�g�z!�U�bn��ߕ����U��5w��vz�-��,F-*3�Y�� 4�����jUҩ奙�Gp�1��e����y]�8�l�HO�aܫ`���:H_8�����ܛۤ��"f��zګ˪�(5�=�z͔���Wˢ6כq�D� �Vr��^���9L�]V��=�ϥ�R^=G�3V������	z�4�Tԣ��l+_d���泌蠤v4��ܓ%�uq���js;�����Ќ��=y'8����ȕ���q�(qV�k��_[he�0�Wl|=� x��R��^���⚕Һ� 7�uuн���g��յӇ̻�������՞�����W�pgl��魿J���g���]e;F�,�Q*>-ٝ]���-�k�f-o-�9��^݁Z�O\�ƴ1�;�ձ���6%a�j���z=�-��A��`�Y�u� аk+��3�UV�v���]V���K=���Z��[U��f.�`ǿ0��"�j;s�M'����z�uO���ϩs�gtm���c8���Vj�oDF��s:E���t����(RI�1�-qPѺ�/��h��V��NAg�}�Xh����"7�0	4���MT�6�Y�����xȇ��ns��]�f9���I�z�
�N���_�ŗ��\�rh��Kh�Hp3S�����2<�g�*��{�����~����bDH�t$����?�ğ�P"	��N�R�D��y��L��rȓ;�&B,�,BȒ��$�,�,BȒ��$�"K",�)T�9�,Ib$�,IHX��,��YYD�D�HD�D�$���,�H�,�YX��ȒȄ�D�K"K�PI/^GrD��$%�%�Ȓ�u"�$��E�%�,�*HE�%HH�$��D�$H�$�	�$�!%�%�$�$�!%�%H�,�,IYXK"J�D�D�K"J	%�%�L�D�ITK"K�YY!$�$�	%�%�K"K�YT��Ȓ�$�D�DI,�(�%�$�$�D��$�$�BȒ�,�*"Ȓ�,�*H�$�"Ȓ��$����H��E�%DYYdIdE�%�D�%�%�D�E�%DYY�$I�dIDYX�dIDYT�dII
��%!bK$�"K뮤�:�D�$YT�dIRE�%ID�DYTE�%�D�DYQ�D�ID�dIdE�%�D�E�%DYQD��dIDYR�}�ϖNL���q ��I"-� �VO��{��;��? �����������~����~P���?����w����rH��d�����dI$?���"$,��_�?����*I������O����$��?��R~�����X�O�����R�'���?�O�'６��8��"Q!l�"KRX�[$-�!j$Kd"Ԃ����*�,��-HT��T�,�%"ʅ��,��J��T�(Yd*�[!UDUHYB�!U�*�Yb�I-�B�,�XD�,�Kd��,��Y,�I,��!R)T-,�H�P��X�!e��EH�U��YB�$�Z"���!R�e��R*�T�I,��d�T*�T�,�B�b�bYI%T,YB�)Y
�%��$�)**%"�,�J��d,Y$�I,�)%��P�d*Y
$�Y%B�Y)"T*T,�R�X�$J���B�P��R�R%
�,�J��!eB��YBʅ�H�!I%��E��Yd�Yd-H[$*�Y$�-B�E�[!j�E�d���$�K ��I,��Z��$Ie�$�� �A$�!Z"~�HI	,����y��?��'�ĈA-���$$�`�[!$_�6I��/���9-���I܍���s�"@�O��?_ۯ�O�$�"oi�q�I?�?���s��	"$��$����u�'ʈ��I"$�I�?�O�$Hs�'�d�I,����Ӓ�i<�����������4�$���?���$D��$���3���$���?���}��I��'�%O����O�ȑ~�_�I"$�I��O�w%��?T��$��|O��O쟧��Gd��߲T����DH%�U�>|��q$�Rw$��,�I�o���7��$��v�rO���H�!���7���?��I����(+$�k5z�w@!�0
 ��d��Ho�җc!�*B֨mfm�&���EJTRBB�P���SX�� ��i��	SZ�(-k5*["*%F�T�F�Di���j4�Z�ն�2�YMF�4�X�+6��̭�Z�UVe���������,�5R��֭�4��cf�2d�h͛-�2Uhʤ�R�:���ѕM-�Zղ6�a�����ն66ɵ�M��[Cd�3ḶR�*�S+4֍�V��3h�m�ZcY��Ffl����T��l�Rkl�����Z�\  ��+�m*f�ʰ�X֩���j�k6�k%����R�9�ڵ���iq����i����Y[k0tk6屚,07m.�Qhˊ;�\ʳY�����l�)�j�ld֊�l<   ��(P�B�(P^t��B�
(PnL:oV[j�2z��fEm���5+j[E�u�Y6�f[WS�J�0�wU3��ګKj��k-E�4�]YԩGKY]Z����[F-�ֳ[5��x  ׷���YJ��V�R֋V��ݴV�J�kn�V�i�����6�lN��*�fV0Q�*�5ںL���f�B��ΕUUF��VfR֭f2ֳkY��j�  ��Ol�֮]��BESv.j�̪ewt"����wf�i��5��WZ�E�i��DT�wk�6Nu3U&Z�ɖٳ
6�-�XɍR�  {�`&��tlb�UUU[m��.���aZ�ݚ�v)�[Z*Z.ڳ���[kZt��T�ε�Z"U�
u2klRʶ�A������ �t�H9m:�튈���*��8�wlp  � :t���@h�v� ��7  ���  n:e4�ڣf-i���6�63x  .� PR��u ����AE:2� t� �h �� u�5�0���� : � �;���j�,�[i��[Djjx  ��  s��@� -�� ��4  v�pA�Nr�T�'9n �Yvp���i�����M�؛)mV�$Z�o   O  Xu� h[q��:-�� 	��� �ø@P��U�  ��� 1�(
&�8  �Me�K3"�m�d��T6�U�  s� �:����  9s�N�7T2���` �� 4Pn�  �vwZPӼ�O R���S�0���  E?S�LUE�@ �JR��  c&&�M10LM�eU  zj~�O�����o���_��d_�{��|'xX��x�h���#�;:��X+�⾪�����$�HBI�!$?�HBI��	!	'��L$	 B��}_�����Ͽ����â���`�"�X�4$T�[��p��e���+����뢳.�,�ڡ�0�Y�Kbҹqt��r�����.g�ka�n�m;	^�Չr�+�X+i\ЯL�өF��f���i@R��+]��+D3���"�G5��Z+_��=�v����775�f�
�ޤ�1�En�8�b	�E>s��׺�R4v�0�;7�.���(�F���n�Ѷ��Ʃ3�MKua��xP#1��u�����8��a�F��!2��+^�f�] ��0��kt`�+f�	uS7z�:!�\u�Z��q��i'`8>�#4�3x(�pH��R��#($�L���ku�>��Sv��Y��9)7�x̽w5b��A�wYEn���B:v���S�j���z�6]����i�bK�M�S�U��*{KflR��c�+*��R�R��ݿ���.,��̚�-n�x՝&\��,X��Xщދ	fd�(�7��;Z�^$b+L�koN��ãr��JFmg*�] &�^�{���ZŻb�ġ���(�>d��S�/q}cfM<����}�/����;�5S5��,����l�t�P&i���5�%t�F�@�ˉ.d���W�h��T��-��[8b�X�Ĩ���
�GrYm��/Ȓ��2P&��f仦����YEBMKiX�!IT�ӈK�u���k�;x6�"�ѵ[V�P$����2��'OJ�z�k�(J�c�Ykr��˗��7yf��F~Gi �chPX��1�*a�!�Cp|A#&t�l��oi<jB-Ԭ׫PĲ�kdi�46��6�4�x��ԉ�TM�o
�%��^d�v-�'�PY�X�f S�`É���C�#��4vn�wf�&e�v����4��2�T� BU-�oK�tC�/dlυ�.���B6�N���m#��Ӳ�ӻ�e�����
M�=�wY�u�A�Ud�n����T�8�S����[ܕ��%h���ޛ�2ÅR�F`����S�$b��������*+�GX�u�aܧ�ʴ\�8~f֤�SDOA�>�m���r<}���9�A�ِLb���PU����	�y�<�ք���I��-� _l��em��n�[��t]uAV�
a�"�d!�1Еj�2"uK��ˡ-�[6�TSD��
�Y�"�[�ʹ2��Ã��Cy��PÆÍe�2�է����s��_�`G���ޙ��.#�^��c��[����D�46�d�t��w���ZX�M�e����@�dBM镟4�Ch-m�o.dD�X�Z9�`[�{Z5���e�o昦(�z��n�*��� 8�nBe���T'(#�Ը�^��I��U��K��P��,�M:���@#2��Di���0�x0�pf
�7��*e+�R�@���(��Y�aQ���c�v�g�<G�(��� ˝� �7p�[�.��VVVh�����8TT�"�'wq:�.�˽EIB�dc'!+������׀�)���(<j��h}�b��CR�VDr;;!�cʺ�#�M{w:��y���LI2�9�D�eE��\ՀJ�.:YJV�IH��ɯ�G`��#�o$��_��c,JG)ͻ�3d��t#a�p6�5�Ý3Ę�CD3�5�Y�{$^�FZ�cYו��q*WQnbye��VD�l�R�Ӥ��\��e%�tQh��x��*�Hv�U�[e�N�r�Xĭcd-�%��|+��|���c{X�v�0\p����1X�H�,�6�+�	�.���N�	u���R-���hb�Zw�Q*M���ZiE�Y�/n�wJ�,q�X�!T�l��hD�m5`fC���w�����rK�j�e��GH��o&��;F�V�R��3.SHV��h��#q�h<�,ԑ;6RD��n�x
Z%nT�r9 �`6%�o#wg(��z�[k脔�jY) ���f2���9t�����he�Z5nVm��Kli"N�U>��=42����M�d&�{%�A�a�k�E��^��3 C�2j
l�:X�)jf\�>��Z����%�n��W�F�H-U��`��е�Q,��s��4u�W6�4;��j��ڕ�R��%5[E�C*H��I�0��YSv�H_� Q+p��UaCmYm��P,�͠��b�j����s�SDѻ�A�
f�.̓z=F�4�e�,F@���Va�Y�)#iɥ�6RT�j��"Ю�m!��/q)�����?Rj�[�j�,�K`L�5xݼd���9H�����]o[�ie����4<���wL�*�fI��j��a5��U�G�)��n�-�ѭ9�9Y�(f�u"���X���RZ
�#2�f�M��bFi*�5z�/�9�G3q���-<O)TV���Fܩ�h�cC���(���4]�'4hiqV�x�,��/��BHhctk��A0GM��z������5��%�MMK�������oC��h�N�υ���Euw.�|k*4�J�:jX�V@���^ �q5�n�e閵�ܨ.��]JM]��u��Ұ�g�>
Fh��۰D�V�D	�[.�Evĵ�`V�ϢV��V[=�OB��ޫ�n�]�@�7�h�(a��>	N�:�R��p��ǐ@Dn��m�e�n�[eI�M��ӗA�lM�d��a1p�ܙ4�@Jʀܼ�*V\y���ʵ��v�3��T����X�kx���y�1������F��m�JE.S���+�e�R\��kM'+1j"��1r+R�y1�B� �b!�<����E]��7-z�֗)#N�Zn)���#6�E�ڭJ��u�f$%GLSwI�fM����B�oSn�_�j4����9NP,JP�6�ߍ��|-b`eJ���[)�V��ۤ�V���Â��vB��)@�Mnmj�Ҋ�d;m�W�.n
(&�YݖB@Y"��ڽџ$R���/jZV�j�\u֥���rne��<3k�CBe����6t�����cf�i �M��<�q-��F�8�mf�t��[M\R��m�oe�0h�e�[mފ&+r�j2R7iZFYL3��Ġ����KÕ2B�s�[�M�CH�+8���I��n�PYc����[z��Q����'H.#-�4:�4.�M�F����! 7uX���ja��l@�lj���r�˼���\b�q��dl��K���~��섄�r�{�X��%�zje�Ò��@Ebd`�"q�p�(��Ee����nM��+"������
a����n���M2pL��x~��5x�f�,Ī��%K�,��yi���2��B��I�T<ӳ,�ٴU���$פ[SKDZ� [5�`�'�����E,�G������_L��M�уu|�j�EL9�*N)b�(lk�Ce�֚T�.`���cx��G�Bf0�k���飔Y�C�&d��5uU�!��ݭv�&�I�Pa��.5%���b���[)m�ky���;{BͲ��f���#qf�֊%[tZ���U6�bku�x2��LF��Lӏ7jk�tbaV�A�ق�F�e2�QсRZElw���f�p�([��K��̴�u.�0��2��5�.ֱ��&���s-���F��2�Y��<@���1���2��㽟��9n�i�i5\�)���m����f��Z{B������
^e�7^�1މ�Ì ��]��icw���n�L
��Z�V�n���gVYRTO"M�qb��v4X rf<L�N��� >;���:�nAB��%��HA���aC� �O5�c��O`X%=����&�:�ٚ+ �ME��
�`���O�;�ڀ��1e���r=�v�ݺ�4�k#Rԑ��L#f5xļ�,Y�)�ƪ�J�+5=�Z��pz�Z/�T�����j�iUq�Z���'�S�-�bҶ^-ۧx
�����T��u�N�UN�)��� ;��D��p�I4^n�{u�c˱�Zr���$���1*8�5�i��3���!w������	"�D��Q��x��O dnPd!��ta�u�,��ugS�m8
������=N_����V��M��L�^�t+�ǹ�&���0��(
����<8��sk(��:nd��f��GE��hëc�.�T:۬�5�S�u���2i
�ݗMM٫�^��&�SQ��¬R%V�=v����Qˊ���-��k��E1�sᰣ5��dl��06�JC;c)D�F��Y�(���aw���K(e�y)�N���hq=�F���,�9B	��W4;0T��%���x5�1�b�B���6)EV�t�� d���I�յ�c�L��.������Z)2�˗c1XխPǑ�xR�aQ�-��[Z�yQ���J��ZvށR��"�$v6�`���ӄ-1b��"�%mŶ��:Ib�ݦiD*��<�*�1�	��[IF���M���WE���F�hNj��Yw{�ÇSi:m̸�m�㘵�X�SG%1i-C�JD�W���I�������i �^�2:Oym��h5�^;����K�v�>kI�w@���e��qn�C����'#4#�=Y�=�o	���y�Sj��E*4�Ձ�u6���	�V2�fK^Ie������e����iZ1*�!�%k6�cu��Y	Ȍ�,ͣ��N,8(�e�ܽm�Lm9J�E����B�"7R���fm�B�m�j���6��5Q�*@ɺ�8]�LE=@h*��Ô�=��F]���So590��dv�/s�������
�R=�<Ivh�E�C7Lۈ�X^��z�cW��k�E�
d�4+,�n��;��,��sS5��Ee�/E��wj������7.��'YM��1�[���L���
�z&�7V�cn�I�{[��Y�t����Sv�ؑ��b:e�y�X&d8��Y%�h��2�SjQ<x�� �W0x�$r�'���w�	f�j�3����Tpi#X�i��q�wj�ٷyh�C& ��UMw���"u.�:��̋,�he�sz�i��¼�(��m�iY2n�ak ��O, >Ig�׸��Au�4�{i�8A�6��Ś�^ztA�	�$�b\H��(\#ڀm�%�V$�c*��GB��+LLf���x1INL��� �Tx�o8���Z'�M1Zm�{��V�Co@�gA5SH���U���ڰ���{kE����*�фf�q����I
!��R=
��E�Y��\t�m;҂!Mц�!�əj�ݣ����Ѻi:�{E����i5V��SCfCRhmm
тe"��n�Sh`͔n�R��j��t.�l���w\R1�.���D9��X8� /w$Ũ�Ŭ{7 Y��V����*�;[*9�I�P٩��T�8n�aR�`nk�,C5|ʑn&���I�B}��7b�)��b�R��M�3��)��k�F�e n�Y�rh�U����*[�r�LR�'ikе��Z�!)��#ې��T;,`b�&�@*z�� )�Jۗ��jQ�$���t�� �L��F�4[�j��r �2�n�6i�<l��>Md�(���n��[N;H�7`��Sv�h�i�iNf�{t��"`�����w5@QE�`��@�br�f�W���t�z6I���i�u���C*1)��,����<��Ji��#���J�y�r���5�u��Sդ��O.|��jSZ.�	�9���%���)l[����fb�i�C-�J�������qf��GBN�l�,�,��,�͎e�wH�B`K
�W��`Ivk4[Ҷ��mώ���������
�3tb˅�o4e�I��(UՃ�R���m�k׷���B��Ɠ���k� ����kkxR1K�����Ҭ�[Rf�0c�ƹAX����)Р��.R)��׀=1P�j�̰r�U�N9k�p�t�0N��|���O�X��)6�֊r֬��-U�K�@e�V����LJbV"G��y��Ve<�&�驀pܺ��]^9.��l��Gm���b�%�� zTSv�@�{��WO�j�v� �ѡ���Y�H��x*��y6���4j���w�1���R4�wu���,�,��|~�LGB�i{�Aш��LKo6�C#e�O��7��m�dY�hYcQ�Y�̡[6e�;���6RF�]�d����@���J̶�,ʙZ,�uV���&�湒���Ob�Q&��I����u�1a��jĶoT��Z]^�s����K~8�u&7Q���[Aa���e�[B��؍,���˺c�6�޲�WzE�T��4r�]��bjǛ�9%YN��*ķ�j*0�.��s5i�4k �jśu�)oh��J�-KkE*�{Z�'�h7�&���c��B�4�kXW�3L���^��̻���,��AEi��e�[ώ�U�JG3C�˨P���*V���\Q��jĞ]j̫�%�k#2�4uEx�1h;�2�Õ�P�0�mеV��IP�M�m��V��wr�YM�)�����^7m� HQ��SL��)�hmGG"���+�n�-`�
�&d(�P��1�&���u��v��6�S�e�(��n�70�n�!6-��X�!�1�v]1GM
dۇ2��5rNO�!6������1�l?���zܫ�x�;��bՊ#��wr�s>�Y����Z���;�́���t5[�I*1�8%]�o#�cwD
Tʰ��a�}���VUn��ٻr��
A�M:f��&�o5ӨaW��OY2�']�:5������ɛw�D�LЋ�����ӷ����N3��%�8�MD-EWY�7:���Jvq3u���z�	�9>|��K�q�=�xw��]�Hs�mȻ��K�Μ:�b���"R7�rh��UCm�9�yJ��:q0�J= ljZeCq�[��r憐gs�������7�n�4� ���^�����b�X���
b��`�'�Y��;�Œ�uY�UfJwP��D��5��g�m=����7fk~|�� %�Cc�oS�؈�Zw�ek��{�����R��Žsw��z\h@����D[@�Xp5����:��$�⺮�Y׼Ng_��y�pf*��k���˼���{�ǡ^7X�U��:�\�]A�����$N��ab�V0t>����mjf/�B30�-�S���Y��R��o7u{Zw��K�jN�)4ӕc�ڷ��ne�N?px�:�D�ܗ5�-���h���S�b�v⎸f���)�C�(��G�y2
q�V���	��Woz0�3�.�ާ�첱����s��ȫ\7Ҭn]��	5���r�ԡ�;Z��t)�|�J��u4�8��4���z9/¯b�-�r�O��E<�W��g�"� {\�V�Cm�c��t�Nlٖ��>����b��v� WUਔ\�q�xԻr��wr{ѻ6���f�ױ`��a�ǆt����ew�Pxu��MI�3u�����7��Ƣ{��<Нö�Ǹ�9�c^y��м�-uk;ӳ]b��S��}�$�V�f�jouk}�bA���6!<,��a�[�s������q�]�dۗ)xo Ϡo��V#�HR�o���dk�^�pI�4��j�)�5�c�ux�;�]�Fv��ś�WSr=����Z�:;O���"�Z0��f���y��;�������8 3�m���;�G��gKMX��
�]���hV�9
L����ͲE[םo.a��Σ���\Ĳ��hx�v�T��뗩�Z2�C�
�cfE���0���:n[�N?�s�������۾C}ǇRdPV��b]s�t"x./��ײƐ0�qCj�YB:�
����8J5R8����ݤ�m����^��Y'"q3|3:�!�n����6����sdgR���Z�˵��_=�^;��E]����;J��#0�N�n��<�(�{�#)�'�����'�~=���9-�{١�"'R7�y��:B6��Y	����5[FO�$��t���7��
�d�w
7J�$���|On���T���2��֙��UN�v����Fyl� n7rn��>�{g�����g>-�߯�J^K͓7<.<�46�d�$������J���V@�O/^֭L��.��J*��j��0;���<�����<��J=[�*�-i��rT��`ݮ��Mһ'���0�V�S �׼���~km$�'u��d����&��ѡJU�kZ�P���{Q���M��p"FY�x6TU9��
�\�w5*�u		},=����(t�*A˽��0
Z,�L��|��'�f��a ��@�wk�v5#MYw6�X���a��,p@CJXᇊ
��`��� �� ��h�{�%�V<_2����@�r0窽];p�l�DA�H<y7n��F���Ty�o�y��!A�Vӗ=f�cѕ���!��﫦��娸lM�e�����{��y�����v�ce��u��V1p?,���7x\��S|��^�\�x�F�%�4�Ik���#�J�dB��=�/G�7��ݴz��2n�-��Vs�å�E.��m�$���OP5��m�T���i�K�ǋ.����Ȕi��f:�3�+b�s�Ⱦ��N�VRʣ���^û��q4��󃺻���R��:��[��E��~��t +�9�q�A&��'�#���,v�H��}}b��p\LԸ��w����a�ɒ�S�G��X�$�o��Y�9�!��,:�${�x�jB�5f�u�P�w���a�ƣ��.hO]�7Z�O���u|@s�q�i����U��Q&�އ�dڧ]1A��<�n��[�E|Q(nvebv��r�	�ůL���lu�nt�cF�|W�A�pšOW�"����+�c�6�x�$6��^���񸅻��<��^�.��r�ÿ�BY0�T���,p�z�(�&�ԛ+�ɷ2�+�N�AQߏj�n�1��u��YN�A.M҃�od�n�@�|o��kq�E�쌃Ä�ކ����٫��9
|4ǁ*l��:�E�e��5� xe��y[�_��C�{Mi�[�as2^�7$]����0�wC����q�8NSP��8C�Y�1�z�����v[r�?��[q�c��7�9&ʋ�|��2n���D�!��?lHvxI��U����d,�]������*�a4�z2S����Wa*���rQ�V�H�ӵ�r���˻��<l�<�N���R�;Ԋ�][�f{�<���l���MP�Z�e*�� ������ݵښ�ȓ�V�^��m���)�i>=�k{��Ρ��qMYmf"7�;��!M����z,^�*�G�}�B�[��:�\Į�"��/��h�}8��d�0A�dd��V�.	y�eY�u��w��<x� G~챼�ju�5h!9�'N"�kפk(aieM����]AuKzq�a-�o���m؊��ׅV�˧��)<�vG�2��叀�ⷻ%���q���Y��z�p�樂�[M�{������N�� ޺{���Eve��j����X\뷠F�̺�Tg7Yp�Q`�x���7�J�B��E61�,�8��B����N���H��e�h;[A�H���\�A��o[���a�z�}oi��X�Q�	�kF>�k	n�ہ�6'
Af��#�t��m�gh�͐<R���B���b�Wx3'�a�XӅ�F�՗��#Mj�b�ើ��<wη���^7ԙ{ܳ�C��}D���M �DwALu�_z����9���̝l6z��q���\�[G+k�1�N3���g��� Ӭ��lP�$ݶ4MȔ;�&��4���TF�Pl����&Wꕮ���vЅN1��γ"��������y�"�t/q��:>XI���]~���Cɋ��ʲ`�;��b{�hϝA�2�X�a��^Ti#ݺVM���7���8�.�;��0�V��YNښ�c���7=۬ryV�N/f�n�pｽ(�^�;6o9F���/���6(�#彁�v�^t��P�ŇZU���ꛗ
<��vV�ut__+�Ӱ�;�Vu'8Z �WH��b��y��s�ݕ��h4��\�}]�V����]f]Ș���9qo=�hF^��u�2e��٤�.��_ma�Tn@&���BxE$:�v5�eq6lk�v����8���`}���綫>�����m��k��nZa6��v]���Dy�meq�5��f��˞���F�m�ǜ�a��F�K2ڔ�c���m&HPL���e�ݚ0����C���9�k�F�v�)�[��i<��7o��`dے*�i��=Kg1v��1�Ĩ���������)�W�'Eech�w5r�$�}n��v�kX��w{�ۻ��<𽓢��}�G�ӥ��8/19�w�t�����I���)'N�t� L	��''Pm=����6nP�;�z:
�V�;��B�ٵ���7Os��N�pF����Bo<J�2�ŝ�J�(��r�M&�w.��ZU폱`ͼ�W��/�1eS��E�/���6�׽���\��L�x�Y�V��ZƮ��,M8�x3��om���a9�K�ޭ���.���A��asv��B�V��k'�4��r�[�A���Ee�/U�7��� ��D���i={���_GF��z��;�������b7�1r �QY��uӋe��o2�S��,uh�
}anj�g�� +*��M߯r���r=���U�dte����(��t�7\������z�����A�	�8V�0�|��/�J��t]��u�ĪY>�Q��!>�u^�N�v�<�+k��^u/���B�����s��;���Kj�f�9f��Ӳl�1�(���7/�z^��%���;6��������-�W��2Uf�ݶ�^վ�J�q�f�V�/S�����s"N:m*�zfYթ-D1ԧ�:Ӌ%�F4z��0���瓴�u�>�P�GN�m^�U���|�����|)�b��LtӶ���9��F��6-��+��w@���.�J1m�ct'P}h4;M�\{x����[�u�ξ�3�#4��u᝔��w���}�,�rwCw���_0����ZY2K����3�XH�s������h�\���e�Ok��E���L�ƯHk�R[ܹպ��sm&�AU���C,����OMWܨ9p�]N�;�&q4��|+�-[�3���svn��a�����H⦝�=�	R=�v��Pb��w��>\�w>�4:[�����<�/iQ�&��Ӎ.�|��{[����z�	��-�xv{9baC/2&)JVu��v�%E	�Y���;X�����E/x�׽����D��b��r �A|���^e�|n42m��,�\S6�Js.�n�֠���l���]�J|�uL�l'��g9Z���fh��b�l,�e�xB���֕u6�U�ל�v^�«(�ǣ����J��ł��eCyhM���48��7um�R7W����N�[KGJ�}���O�d����E =��R�K�z�Ų������\����t'�2���F�N���69U�&����y��%���3��5�}��G��l}�^�����&�5���Ⱡ�\r�p��-H:[�,9��;y��4+^n w�s}Mrzf�0v��^���1Ի��֢K^�p'�S�hGg�Hs}�uS�ݚ�?=�����އy��*��n��&�ID;�Ar��z2��O������S�ǴD��7���F��-Y묒E�䫲�g����+��Fx�.�y��ۿx����X9�l�gG<�\^X5w�r/\{��t�v�Oo�5$�
���H/��V�v	��r����_+�C+�wX�'n�N�
���X�9T����m����c��o��2��7�h�T�e{�E��BSL�T�C���w�n+1Q�,U�n���OC�f��͝�� .�(���E.�~�庛�8�͹�H���Y��d���h�3��f��s���H9�yl��d(�Nv���ɔN�9sY��l&^�{r��\�G��s��-���kU��K��t�]�:"6����^�r�HcQ���,��煜@�5>�uY�3�׺M�+(7:'og�N6D}�.Y�P�}�LJQ��[���{�|ͯ�f� �<���±ɫHB�o���R鑼Q���Ǳ��r:��v�y��#K��U�}��b�c�"WY�Uu�5Vh��.�MK
{-m͍@Qug��7�e�n�׾��3<ʻ�N��'
��G|�-�"$(����.�(�I�6����ƶ�K��\r��u�2��� ��+��q��V�ˤ���m��P&���wP=��f.�L�T�Z_9��b��m�%�=n���W<���貲�c2�t����i.�>�*p�d�F`���5hyw{��󣱨G3��=�K9���7���z��P�ub�Sfjz)�&zp���H���x�(cz�su���h��'�JT�6�!����hͧ��뛄��o�Nu�ە�U��泛񧪭���@R��}��`�h��Bu����5{ �_'�	�>�G�V�}�2�ҁ��`����oS�ط&�Mn]�Mk�<�2|��n�2��-^���}.-�zѨ���5�0��0z����%i��H�2�x��L�ƴ�Y�!�o9
at��kݥ��~|T5���YSv�z,����^�ȓ~_Gi�/M�S:�KӜy`�s=���t�[O��b<�˥d�)�@�3&�n�B��v�����A�����I�՟C�����1`��9�<on�_!"<X�M�D�4^�B��쵲��ͅ� ;�0�q��Wcn���j�����\&fu��6�p�{2�i��<9��D%+�e�&��/S�����[] �N�n���Y6���7�N��5����I��:��Ըܮ����J!vx��s����u���ZMl!��-�\�J$v��W���F��8��ѥE�{��VF�����>j�(+�bڽ���8��d�	ƣ�����!�C�R�͜�o-�qtg����CM�a<ťlj�2�ʞ:;Z�z^K��4���v��}��C糷<�U�h�K���e�o/RW�('��[��놔�<7�Hti�ou�`��`�Y�W)|]�>�����
<T�kk2�6��k��>�?�4��eU��O%k����JЛ��Գ����F6�S��E���v�������L^�.�ւ�ɺE��r�fr=��j[�f�I7��ѥ>Ȩ��ݛ�[���۶�d�l ��iǤ>��;��h��}���B�,�uݗ�W�;��f��&?4N�
l�wO<�7��� \�o��4���]�R��Է���i�lM�u��d<j�f-[2�\k���6x��oL�8�xq�}�p'����P�M"��giLv"��STu�Y��_S�{⨉�W}k��Qz�Z�D�6,ǯ}�f���ufK3ϻ�ȡ��M>��2;�}cs;5�����yq�Ɂ�eGq�d��H�tm�Wh<�$�]�Q�=/u����D�y$ۣ۸.ۂ1��e1-[|���[V��8���uъ�-]w����Ͽ/x���W�y�����$� �����������{[4��i��"��W0N�������*|v���"�:%kN)cz� kS�-&�L1BWr�S��x��w-��`�b���W��<�X����@��:���g)�y�]�ء��VԨ_l��N�b=���z��֭R/k2�-�9���"�ܡ���s�Ř�nM��:U*�*e�-m��X�1�.W0�ۧ(��s�5��Hn���th{�kۧ��Kh*!�)�F���}�m�#׾�v�NM�6ـ��Ad���V"�6��0a��p�W	/q��cl�� ��y%���X�V�v=ܹ�Mafp#�[QK�q+7osgF�!ք�4z��c��$^�G���Tqo��R�b�ٰz+��s#٪Pz	�[���S�L}i��<��,x2zݷ:V����R��ʺ�C�0�]b�`N�B���Lq+��Ń��Z���U1GWLL�Չ�7��Ò#�s�-�	�2�r�XW��n��]j��rR��>�ڨk�n�Gq-�ᾏ�7�ѳ�+�JHfn՚h*�$th�檅kQ��@i
�}ԻV���,�r��i�woD�`k(R4�����˲������.��P�X	ty���t��!|��ʲ)�;�)�s�|z�<#���R�to�bѶCq�=H��}�1��Ӥ��*����Ԅ}����m�������EӋ<�Y����X3e
b��s���ʁ�y�,x��M7��������A�3������']vo�4n�c��\8��l��7z�Nyx��&�O-�f�;vLW|��=��㝋�rl��3>�
�ļypR^�s	�L�ͦ�X�{�i�����^w�c쏬�cڼ�-iv�K-��F�l溴��6�g�����u�˓]^RzU����]��v|����>�#����H ݂�6������Qݝ�K�Y��/(��&��^���b�s.��ϏE�U�@*`G]'Ӻ=��9@��.Rr��ｮa�B�q��;KQ����vwh@w�c^�a��R��8
֩���f�d(>��7lq�]ut�DWq�@���K�_Gq<�x	�H1hV�.��r��]01�R����;_dY�\9��bj��z�x�H �;����"R����@�h��찞����.�cb�Y�W[v������zey�&*ss_[��Gi��lm8a�k��`y1ܣ9[��YLQ��ӳ��D�#']�S��)b/E��"f��Ƕ1�8�~m��f:}gk��v�̸
9a��+먞�,ذӨ�_n���f+�w�u����84Zs[�Z�'C6�QP��W��⦧��l��KPvk1�"�衲7tQ�� l���w-t��)���B��_%}EK����S�����sZ0/�c�
ufQ»;�tn�Ǻ�%�)p�O]w��GG�v�"睺N�Ixq>q���A%�q=�מ�3�\!�����BRp!-��Ϯ�E���m6��H���b���]@J��W+s�ї}�2����. �ZWr�8�U�������B�:To��˫d�ן4���u�yx�(q�)�4h&:L�tl�>�W���T�WP����!0����Bc��%vUg��48��wd�q�.S�J��WvZ�.}�ᗋ���G~�YuԢج�`x.�T��	!: �~'��.=�/a�K9��RZ�9�%"(��u��R����N`�����L�證��f������w���R�ND���1�N�ժ���"$�M��kmφb�2���iU�˛������SIz��]Q'f�������sx�;�]��숤\ u�-S��i����Fe��#�_?��]��eI�E��t��JB��b�e�om���Q��#������`�ڹ�O6W�+��k��\�  oht�������5���oL;��Z��́:���t��q9C�`���6oU��3��Y._V@�A�����h�!n�V.����д1J��y/V������&>�����٫]ti�*w`ΣS�����_,��w`l�k��ѳJX�F����Z�NJ<d��۵o��R�\���^I���{��r�3[o���8o����p�+�����Ј5���)Ԯ�L�(͛}txn�4~6
T�O�m��l(��}A!��]�w*Gr6����u�;��"�U� u��T�9W�K	5��5yx�����j�@���9h��u*�ky����{5Mߩ�u�Y���%<*��񦴦���fz�4��+Ǳ#�*��\� J��4jjb�e�ǻ :.Z��0�'�a.����w��6$���6�ݫfY
�}ŁY�p�Z���4��D���/�^���`�/�3����Z��U($WZ�*��\a�<ܓ9�1i�#!��@is[Ku��Gs����pz���{��!{�_���Q�HLb�ˬ¢���v�(�����*���Э�F�I�V)l��^�����`�:�>vx���"h�ZV���}�|�0��wʀ��h�ڑ�9C�Q����׃So�BLI�,���-�]�����;oOޜtT�}�GK��\轐+9�ő̝V�uH�;��2x=��c��t�Qr��*j���]�u�VvH3^r.��;���w�ޫ}���Ҷ������*���w|:`��y��V:��XV��髺��=u�/+��c�x���;�(��k3 �k�|��uܴK��dS��ni�V�X�&h��������I��3x+1�dl]+�ԑ�������	��3��r�(�9��AG��0�y��t ���b�)q���]e�ܺ��[j�a]��h5n�M�����B�{�~���<,��o���govY�jW�n��CV\�5ಋ�Gu@n��IV�i��f�-���yʰp{VI��o\ٿ)!3U)J,u��YLQ���B�m,&:��UN�_
�ə.���MVY��gZIp�E�ݞ �Ӹ(]��:<W^�H�	��j]�p�]�6��	��c�����s�<��y-Ÿ��z˖N��7�Oݞ��]BŨܤ�xˎB��V�]̼	��|il0|X8榻�-sy=�4>w ���罠��ޔ���k3�4�ew=g��M_�j�P#*$w��
80��@�kg8�Xi��F�o�jk�h��� P��I���:�'�
�5��A�.��$�QQ��*�wTe=ބB�����)��n�"�/˥��v�py��Pfs��bB��w�'SsP����ַ�����4ܫ{�:��烾6m�+g����Η˝�W�쐗D�{5z�>�cWDBG�';��
�y��gMAxC�9m��zV��cnU�f���V4���*.�A��x����h�s��ţ7�f���x�{EY�MN��s��6j+���o.��`�<�Xpf��@A���Nw��f�u�p{�(���G�C��\N�5�m�n�!UK�h@;Ғp��9��B���ΧS��5�@�Z�����n���#w��m��@��wZ��]N G���X\�qZ$�����)��E��V�Vb�ȺBw�f�G��1[Z���+�W�g�j�a��ƅ�G(��%�,4�(�qm5Zڴ��ڀ���;��+%氞��X����:-nS��v�ok C�E���FJ�4���[�����E�6}U�}����9��V�7�ދ�w�]��q�c��z;/����ǒ�����y,;��h��|�	J��]�c�oE򭨖]Z{�|9��5 ����y��!��7��Zb���>�Yմ�^G�P�]�{��]X�p�d����{Aom`g�T��|��
)�Ͱ����n0nWY]�`S+��(�X-��V�	zG��_�OT�[fy�c 
j v��m�LԘ���=�|������k�!�T�k(���R.�m�ec'���� �;��	����~t����1�pg�]ƽ���r�㇥[��X��"�2��z���k]y�h��Q���aӤ����<ڱ�7�)a�$շ�YH	�% ����=�8$�u4�`���h����,��=�_c�N��y��e]��as�}��w�{~?7|�=@��K{�<Qꦣ*o֥r��:D���m�+��V��6����Ҕ�c����G�wu��C1,���ڵo,��f,:0%Z~����4hY]��߼��mǜ�Lji�.�[� �m���
�d�|���^^�!;�}��u�����z�)3�V�r�}%1YȞ��G7��3�:h��\����%����+]�
��I�Vv�,���,P�����k\��T����j\���즓�)���x��L� ��1���׮��3kh�c^\4����^�^�����|kݏw%������7~j!�J�"�P���GGCw�=��S�W\Ԗ�u�T���n���_R��y�>xy��z����=�\�;�H~��w
~���0�����\�M�9[#`^��*�����W45�:�=�]Y�Cg/���9���J���7��kZМ^�s;;����B��Hں>��M�PY��͍oAF]�G�UۓTrrbu�����,�VŒ�bAWQ:���a��{!����on�*+:�_8:C���j۽ѝ�xC$�;(+�	�!كc��:K�Q�Mos]�5V�sb� ��3u�'�@j�x0��h^ʼ�mJ��S�֙ōr7�m}s�K�st�ά��g������b�zi��I�Ƞ��aL���9���J�e0�}�r"�BH�Ѻ4��w��z6�=��#]nS���CE;��+P\1�G���ze�@���p갠�o��9',��o��c�\��]�^�]���$Q���B�Q�y}�Վ�"��v\u܏]7uì�n��Pq�IǑ#$OZŷ�D�ǥ���of6�R
_��o�]!Т'["��knvu1־E^TѭCƺՂ@
�=j�e+w�,;z�ѫX�W��*wN�{(;c p�t�F(R���P⬙
�z[��F�n��nP'+���2�)1����G6Rz��!�J}�M�@4χP׬@(����.�W�<F�K�V��^�,�Ff�C1kt�i�����֦�NmJ�M��B\I�@Y�����sp�~@:+^C�j���va�_T���Ƅ�9w.N��T������*Ruq�a9KS�<��1i[St��l��W��n��t64�M�w�a�r<\���]qGw�6ұ��4L���a����d�;⎿
W��������ds6���=��G5���}�w:27F-]��g�v\<, �I
��9SIٍݵ�sp��]q���D܀U����{�n�پ�_y�����xk;n�oC*ܤ��o�y�� �h^������{x��px�$���tJ-��ܡ����)�ã��so(r��^�6!ݩH8�ݚ��P�����^Ҭ��XU��ʏ����#��bx ��3h��x0�zAR�����>�k{n'�����L�'��o�5��z�]����g�7�N���gq�����Eܳ�m�<�Yt������J���ԡ/|����M�mh���'�uR̴{h�%b���yY2j���ɻ�C����Ӧ^U���IqOpMvk�}�݆wc��7�p�0' *���)^�R� ���8����ef-˧9,5,LH&�OYk���������E2HFwi����W�� �'��|��/���~��g���B}��^ �(���H^��nM���$K=r�f7�Db�.c:�'e��v���� ���vL�X3�E�Fw����L�`������'z�/w�u���{�:��tf�}w��TEorΛ���g��We� vmm>	8FЕ2��+���8��"��܇)v5]�eE]H�F���ɔ������z������X�����))�1^_*l�v��&Cޛ�a:�ֳ���Þ��]����Vh�N�X���ߒwt�7�;��3A&B�e�y���Z����$W�{.^�����~�_)#i��(nF��;MU�)®�<�c7m��k�+�xi˿S'���S˼�6�-]�i^��2i���8ǵbG6yl�짲�L�=ըq�ɽf�� ,�Ri�Dp Vf���%�N��4y��syv�=]��u��|9����~7u��s��c�#�3JZ�A��
�sMo�?.�J�+93�M ]�0�P��ۍ�s�/A��5Fƞ�ա]�}5J�F��z�����^�{wt_M8s��J���\�szDC��ٳ�p�^[k�8���pݪ%�js:l%����{)½q���Hz��3�����͊9Bح�9v�d�p/L�E�N�~��M⅝kNȱ���aI=z@�w��$���}�SR�L�Ś�v�`e�¦���7�h���K�̩��]���|
 r�[�Ac�1�Ɓ�w�Vny�|�f+��{�v(4�6�nc�1�tn�j�YX�+�v���h+��i �.����ޝ\0�f�b`8�a+�p�B�tC��ާ0z+���е.��V��J�dJ�?uܼ�}s�g{M&=fL^6�_$�l/�M�c{!�r��g��n.��Q��X:t��(s�DoE���d�R�=S�����2����@���]����b�7�ݦPf���+���v������.<��6KZ��}��|4� �Tu˚�[)RٸrTY�@�4$��{n�Y)E�.��� �+p'J��ib�5�f]8Ol�?k&��v�XQc���Xc��v��9��]�z�gD&Ĳ,@ѰR{�0+ˡ�e����w; �5+i[)'!U�:�;;����W`Յ0x��v=��w��u���?��$!$�;��+���;�Ќt}S��Ņ[���Hݾژ_z���Ө$E<���.�)K�ՄL�_ʗ��۶1�&����s�4`��N7�3���͖8����}\�}z P�y�FZ�,�}�.@��l �	sM�+����(U���\7&�q��]�]-��R��`�8��/@����k+ F�ӽO�IA�^7vzUB;��@���=��#&R��M�M٤5�X�9��I����m�{&�޽�;#:>�<n�u�4Fqیr��W:�|�>���U!���]Az֌YBZ�qGˈ(I�[�Tw�w�3�xK�;��[n�i��s�}�b�=�8��9��4	E�*�`�N+�wN��"����8) 3k���	�A�^ѕ;���J�&�L�ͤ���>����cBZo�Ú*�_a�y�vB)��z�^XԇՖ)Ҥ��Nt���6�7��ud�L����wMK}�S����ſ���fb���r����F��R�Z(4���<�ـ�����w����{�7�{G��WJ
� -�8;�c@��mSZ��.�Pp����J'L[2���z,��d��=Y�]}H�01�=P����N�o�r��nF}�p �N��:V�7+;�o���ﵴ�ߜ�y�����t*����T`��V� §i���(,U�A���Q�U�+
V��ij��͙Ab��[KB�J*��Y1b���+E`�TQu+"��WYAD��!R�
1���dX[J�0X"�֩"�ʕ�ETT+><C'4Z�C�!A�T�QQ���8�X()P�r�
��5�`,
ԗ����"�k9��E��B��̪�����+��b��Ub�[[ ��H���Έ�VX-x̯�*(���[i&aU�Ȉ1�P�F,X[EEAEc�0�dedUb�ATU�*�U���s*"T�"�����u)mVT�YĢ

[l�+Q`�x��6B���rN$k�QV$�X��-��YF��U�@ �|2�����莽	���1��j��mk:�P��h��U�x�^v$+՚�Z��HU��wk��%�ߪ 'cG��&á��~c3��IhSqHRʭ1,A]i��u�u�<�l9841���[�g^�KkE'�Y�����&��p#��!p̋�Pj����mfC��u����;c[	�,�����:�tN��-2Ϫ h�{��*V�|j��2ꟲ}�V�g���t�Dw0�a{��Nt��m���?cZ���R����XX�t2ˊ��� U����Q8,2�'�S�z��xO�T��^^S�Lc���WF�����Դ�)˯Rõ����=��٠̫��0a���E��j|@x�s�_�Έ�_m�[�Ƀ�|�ܻ&��=/��x�MA����cߍ�c����a�8~x� ���_o)�w?i�+v&���=&ឥ�Y�gG�����-5��]�1W�z��h�^�Uˁ�
��M�Na�'2�_jvs$�k'����(`��8a�l`�E�;�4����k��M����I>x�9]r�e1B�f�vB=�0�O���'!����c�ȊS���kȝ'��e�h��쬨ήK�@ћ��qV�V�v���e�ռ9Ϡ�L�7��
�5�I�JN�TT��D=ɷ|x�V�3\���ԕ��n��`�gm���sB���Q�*�
:���LOc�Oq��>�䤱�;l�{���ϮhQ-C���o���d�a��cӊ�lLS�m��6) kHqL��m�&u:V혻��5�!�"�wKd�L��z=z��@
vJU2�!������p�4G�u�:�����.�ތ�`=U�l�u����f���i{.Ս����W��WyV�p�e�R�����S8ύAU�i�&6}��v-��׸�� ���m�we�e*Ԛ�k )͈��*���,�~�t�  �ӳCxk�r!������VƇ����bB�V��{N�E�:{O��g���쀣h�8���Kd���� F;�c�97ƈ�����\����W/vE��da�2���Z��Sc��i�>�a��J���ߑ�5�G[��~����y�:�㧜h��[�a���YB����Bv���KG�\y*�%�Up�W���-3�����Zy��'�ie$+&���z��/�
�
&t�,�V�1^�QS3k$��dng{=Kw��"��bc5�y�O[?-mU!�޻�Ax�:ԫ�.�*��v��Y��7ȧ�������BER�Q}�&�8�t����y�$����/r�b�i�/��.k=�3V�<SY��<J�����ET��/#ɰk׫ڻ��{�q���#C(f���Ft�mp���'��$�F�}����QN�ڽ{�-ͬ<
GZ�P������W^!����T̥����esƅ��ۯ^b׎ꏃc��kO��0��k��4���(��"u�m
��E2zb=����^aX�+�[�\���ʽ��]Ge+�R��,9d�}�%��:��'���^�g�^�D�+��~��V"�ċv��kO�X����$݊��瘘?,�Aʵ!Yx�>��'ʽ�GuU���?z�ֆR���mm�A)׷l�.�s4+{��&�g�.�Lw�Oc�4���:��������YM6��lP�kY�_/#Uןk��'�\}qo'�h�y�׵� �t.��h7J�ERA� @ڗj۔S�l��[�E�iy��~Y]݆�[��ɜ��.���C�w�kִ��q�Si��L�g��gE1U�g�h��(�%z6)��b�M�a�=vO&�z�`J׾���{��+F4>�G+f�'(���=���	1w�V`�e(n�Q��+w���A���x<N-U�^:�ƫ�z�9?"���X;�[0|΃�*_�$!Y(~�t��w���� |/l�]�Td��Y��Cb�3���\��&���5�e�EJt�гuخ�.Iȋ���_foM�qǥ+ۓ�:����j_]FJqF��:�^�Ӿ�N>�F�z���n��m���X���S�vrn��z�9f�N^��^
ӵX���+�j���\I���r�f�t�&'��}��-A�Y��~ߤV��<<\h�l��#Q`f۔iQ�֧�$�SvB�p{�����]�< ��z�Ry���1���QV��u��T뱹<�ׁG�JJ3����;��=x��!.���q�Qw-�o�1!O��-�h��:~}&1��wo����V	��z��sA����+*�P�"�~y<2���W��ڃ��Zm3]�ڽ��Xs�u�@}�f��;
l��OL��k����S�e��̊���e]����g��/xB���m���rυ�a��[7�dh�L4�;�b��ړ��t)��U�y�wp����/*�Y>�taq�Pq+��sć�Y��/�UlB����ؕ[��ٹ8���U�:���R0i�U�>�U��)�F��o��\+8����x��(���e��{����r���w��������W'�v��ŀ�~�T�{�P�;��z,�Wm��U
���5�kϻ�;�L�nz�,�u���k���a�*��(��$�;w�ŠsX>T3WR�����gx��p̗����<c��rE�_<�w��|�\Хa��y����td�u��q�	�1R�e�
@
x�V���EF���v���Qyx�z�����W���m��;��Lz�0;7��Ɨ	'�Vu{�!�Nq����z�~"�҆͜�ӛ����d�M���ca�L��
��7'��x�Ztf�������b
���ڣ���=���÷S��Wʀ�S�yx���ӂ�8/�;��E���8Ǫ����D��v8�T77S.�H�a�$��@i���1P���8�V�~����/ؕ�V�\P�^tk�_���i�@�>v�R�-�@L=t=C���o��S��+������E���Gl�iU@Q�WW�����bK��9K�^�O% �g� 40� >�����0Q�1.3���O�e�Sy�5�Yub�B�=��)�Ey3\?�0�٬N��Ȅ25��B���z
u����&�a�o�$�M�}=����A������9`)�V��r���hy�h��:yE�۪ܲ-��٢<�NOf��'u���q����,z���2�r�@vlx�Z�@n;��G���n������l�SI��j�	���s5�o��JC'd�5>�d�M��]����n��]r;hE��T�v����|<3c&>#/toT������؂��ߟ����=����j��cY��n�_m-nԻ�:���fs����k�f�
¼D�#8���:���d=�����j���x���4J.�Hz��ƣ(c� V����(���,Z>��/���<��:��ȸcQo�H���|B��	�Vb��ud�,��*vr Mx��'d+L��4{b:wٌ�L�I�;�˥*�&>�k��;R��;�ƹ�S��eu����e���f�A���A��-k�*��\_=|(ϵ���f�w��7��)�ͺ�BǤtKS�`�>�Ƹ�"$�,�N�˩����RrLBֳm;Q���%�vg�.�O�����ᅩ�KD�Nn?�^���8����S!3���{��b}���>��L)����	���Kz��h9QxvʷX8üpx&�ĽՈ�dz�_��/d��YY�X�C]�����C�N�V�/̡.�{.��3�c�����]@����܇�[F�,A� �̡�q�AB(g�6�����x�J����s�[�E�u0G�u'c`��7�U�Cv�'Q�3�� d�R@�P�lvp�h��Dg{�҈f�}��7E���fߵ0+'=X��j�1�[,
�̛�I�E�i"��?�������k�ϸ��������Ns���
��zS�@w�@���A��b�P�Vr���U:�	ƶ��s{8=�f`L_i����{Y7��0���PR�Ќ��Hۋ���y�9���u����{;*ǭ�y	��#03m�r�Z�U�y�����^y���K
��[`��"ǅ��S'��CΝw��Q�8삑�5���� ��6��w	 ���2�dU��?"���+�?�c���!M���H�k�%
�d
�Ȍ�gs�/ӫ�Y|*Ǫ����{���/VO=��7X�'Ү*����)��
����|��ڭW2ME$2ԋ}v�nF�>FE���P:�B��H��*��B��e{��?1T�=~�m�f���O=�⻨:� ;
Fp�����h�d5�[PE´�^��֞ �8�^��)�9�I�w4��I�wu��,�g�W���w���vy����]���ƭ�3�<'`�`��}�G9=B�[y~9���}թ
�X�>U����6x�X�k�����ً"
��Fg��*���|���u�6�*���p�^8;��L/�����ˇ��5y��w`S�_�#����}AV��[̾R����_JO޸��fgF@Ͽ���A��]�Fs�~�2�^/[��7�J�F�i��#�����
��촰)0�`"��^
�PU��e88M�x��Si�QKܦ.����A�X�b�]�}Vr��ˌc|�!J�N��pk'>��n����5����;8��F OI&����:�~<&;����ye^9g�<�b�n0���9�h�A{ݽr�v��1f���r�<�k�g:�_y,�]ܮk(e��N��qMN���|��}¼42�ҙ�D��LUC8֢F���i���b��v+sѕ�ߜ��7�:�p/U㝊L���?p�u,������ۺ�E2vv��g��8�묢اV��J�� ^j��H�Ik�Ю�Vm��azdY�C���rݩ�Zѷ���y�=�W���}ʗ�d�l��H:��3,.χ�����7�#^r�7\�����p��8���Uw���^�Y�n�R���R��~K�Qug�y<|,?�X\4xR�.���v�ս~��g.{�͎F {��+�>;)�{Rm���%1J�gԲ����� ��2;U\=���7�0�e0@Г�
�mD�f]F<y8⨻��Z�1!M=E�t(�U)���-y�����(Iw^��|�6YSxD�h�+�5�UD��NZE�0Ty���yj��UѺ�;���g
~�T̫�壀���O*��}�W[�u�|�Ɇ���*7ʤ/�U�53���{�
��)��3�呓�U�z�֧0��0�RjN��k)4n$��n�,}z'Ī"�7v��Ⱍ�?i�U���&Fw�&��K�/g'k�P�¾�V;�j{�w�y��Ġ2���"��s��aߐ؈�� *��~�5��q�qw<4S܉pI��Nox�}�o�c(ת��%�n��+]W7GK�=
%~2��
�X��r��[��;�6��Y�:���v_Qp��o����m,h�,D8�<��h�3L4���תfuУ=K����M�Ǚ�����Mzo�^	���+�X�\�\����l�uL-�{�mwkpZ������=W\'1�m���2�Y�>I�h��R��d@㽨�C<���u�1�$|ϝf�=���N0��CG�JG%�@J6sf�405f��2�t�C��Zi*�{(�[R���g�ǐמ��:�F�1�Q{�ϯ��{�ëo��u�U=����&�{[�z���0(��(����#"�-v���xy��<%,^ꇅ��&z�J��]yy^C�z�P���!�:�UO������7ܱѬT�r��3�U1mh&iCK�E�ݧڽ�Z�;��1O����H;*P�\7���6�~߳2�/�=��C��D7$���5,��2i�gA�b�|�|/������8t=������<$��`�q+{�q`�����7��db󴮰I���yi��t7_�gxR��1ͩ��vw��QS�E�nU�)�� VH��ɞ/��)/����y�^�5��{����+/����ȳ��]$u/�!v��mN#/� h�� ���e�#P����3��������Uzsg��6����T�Yw�(-p��,g��r�{r!L�@�X��VY�Ps�	A'����i?,W���c����5CH,յp�=2/e�n���[���|�
|��w�ܕ��}A
�n���J�����^_ظ+�=o�t��Oy�Q��:�gnN���O��tZ��6��e�,1���+�ǢU����K9 R:{�nP�y׷<y��	��#�3l��7�or��^o^d��oΡ��vz��u�Sz�hlax��p��8��R�!��]��ґ�cP������(Q�n�3�۟o.����~>���[ ��R��Å��@v³_ ׶����Z��CrZ��|g���TV	�ӻ���י�w}q������O�*�����)paS��A����޶�K��3�8K\��ζł��yk�u�0S]X#�+*�q��>�����9t| �_WƦ��4�<�cv#]M5�#h�]y�r� ŗ�X֋b�@oWqyw*���HM��k7-8f�H���wc��`!g�Pi�sa�b�ζ)�mP�â3�Kxz�uǭW-L�SQ2�t����]Tn�խWa�Q;��>2�˳
���5�U���p�ޏٮ�?|;�4:��N�m�W�E����R}K�b�jwt�<;�8��C�8D��3��B9(��F��r"��n�N����NYK+��� �����ޑ��L��[�Ap��+�
�7����읒�{�g�Lzj��`$co�ěSZ�]��3���"��i�c�ͅe�:��'�dSXh�~/����j���*l����0���@���e��-��FE�9	A���hĦ֎y@hV�a���z�쐹s6�T�mx�������a���Kl��0�00eJ�O	��a��	����J7b�y��؍f��^Jw���4� �e)��5�G��eky��wp���)'kc[�6ˋ8"j�:�csw�N����7vE���f�՚�P�-|���|�[�<U��<yώ�Df]�%�c)����<d��Vj��O��^�nȱ�h[�i�7O����o���7,��{�6� 2Lݔ�<�u*��]��Ӫ�e��;%����b��]{%y���H���4->�޴'ů<� Ըh{����1�`d���>�ͤ�E6��?"��O`^��:�I7Q��H�at3�Ee��I�^���I]|����V��9u�[�S�Վ�CUv۳��c�O"��
�[���S^6H^�4�m�96���M�V)�1��h+��^4�&�؛Dvb���4r����6 <�*h7$�B���ݝ*�gjښ$�L�Չ����f�gEum4ˀ�����	g��
6��]���>���[kg��r��̼&v�y�vQ�9�Y�B�J"�)i��*��
�\U�k��ݍ���!O\�����Fk\��ո���\�'=��b����J�氏�̹Ds����f���撨��E#Iԭ�f���{�>�t�*[ȅ;8����	
ò��;y���Vh�t\.>޷�gWxf���>�(]5��Nw5����6Ա�ŻL��H��eJ��K�Rw�xlĵ��h��%d&#ov�9�}Ԯ^��_Y�s�V�j�Oh���Q��W���Ѷ5,�I�5�֦�����)�3d˸��p�hr�U٣�=;�X��z��YG��{���L��� �L:Q�<�L�� �ע�H��{�}���h�5�a�-o���ɫ�:�be��80�D�H������GYV����s�V�E�����_vfdZpH�	ޜ��|.<��ID����O�ف��J0��i��Wh�ۆU
�to	�v8:H���
�wX~���o`Yn�mpI�m��q��zs��w����9�
��q%l�RT��m[������h8�p�sJU��݄�t�N�u]\�BPϒ6���o�q�4����lF:N������.Ls�/��Y��AE�?�TY�G�j���UX(�S�
��Y��cb)˞2Q�T�IFE@Db ��*��q�8фX��V(N2ZW�
őE��-��B6�W$�3PU[-B�r�����J�bT�^%Usvق�QEV2�""�2T�H��QD�2J'�,#���x�(���.�b(�kUPDX)N9Y���Eb�DP+�)S!�#l+�IR�V*�PXq2J��B�q�V)Z�jB�+b�b�,U��A�aS���*"��̬R�,"��I���q�#UAaĕ �m�T�efeE PF�E*TR)�Y*#"�A�2��N!DkC2V���TY*$P,EkUX*�*J���PD,S[��"�Ŋ���&��E.e����9jW�n��ͽ�����
�h[�u�y`8�U�Of=�'7Ns]�Ý'�3��l7��s�}�|�؆�6��xx�$N����O_�{�g��=O�����X���J��)�T?0�7]���|���g�ҳ�J��T��z����ɐ�������z�z��ɱ�3\O3Pl��3����R|B��%��\��8�Y��r�� ��~�d�<r�~���0�>��{�8�����w�}O����n���>���}�$I�+�;�+5ݯmYח{3ް��7�eNS�,��&d����O�T�ԝ����g��^����L�aכ��|偐���C!�g�����'P�/�;�撫g��^�P��!_��.�J-��3ͱ�+�`���������g�>9�~��T�AVNҤ��`~>�s��������'��%eg�g��	�Ĭ��y��%IY��e
��'�L���'x��E�S�U�Z�żn���.oL/5�8���`n��|J�8�`=w��>���~��d�z���?YէI�0��9퓧��A{�@D��Y����N>�-C���w���`{�{���C T��j�IE�O��Rvm��6���@jaP�]�!�=J�C�|:�N՟RTS����J�N2d�ZO��%��:�a�z�~2~M˘_��ܝ0��i��l�*O�8�������Xq��.��x��3F��o�9���g>��߹2:@�*��5��3�}Nî��v�U'���2����H/�a�Y��&C���>�S<C��(%a��׈'�T��gq�X
��?5�ί>����>���nm��(x�L���<����%ACĽ���!Ұu���2r��{�2���>'�z�ô��R}s��ZS�v�U����q'�*N���3�l�@fd�x�����l��y�8�� v�N�Ӧt�����g���OP��M�C���0��:�����Y��δ��'>�Y;=�$���g�Ϻ����~�i��/af�>���w����-�����{���}����uߵX�?Y�d�`g��|��~C�
����5�3�2z����UT���;C��^��{Ϝ�V}IY:=�|N��+�>�o���*q�/�S�z�q&B���'�H��b��k�I��ܓM;�&�e�cx�t@���Z��݀qI��oV3t��s3� Ϳt�f�!�YIB(}�Q���Ң���JSM�ˇ�v��v�un��1����K7�[�������*m�<챁jܢ�5��r��6������l��H3�s�j�����c�쟞���3̣	�fAF�� �}���J�땟Y*A}a���'i�?^>3��8��^���Ϩx�!������Ad��̆O�f��0�,��&D����_�������n��o�s~��? t����,�d���|��$�s���(N�w$<C�?!��d�9>c���~g�?$3:��!������}��7�����4sNL<�쿨�H/�l�d�!P��b/l�&g�����;@������ι<~��%N�Xq�Cĕ�Gw�q'�W�z���N��%I�x����:d��=g��x=�ѡc�p��w�2K��d�3�'�����|�v����9�:H,����S��|L��:��� �?>'ÕH/����=O�v�R���÷���̝��N$�
�����dP�32���V�9�GMf��T��m y����>��%}O�>�N�<J�ԗ{�q'�V{7�y�d<O��+ t{�q�2T�<r����8�_����v� ����=��=N#4��`��dgwt��Po0���=����8�P�=��q�����Ag��7�=�
q'�*u߽��N�<JΓ�s�� T�'E��0�+�{��&C�&~�p��'L钠��Z����X?+l�)�"��#��^��X
�a����=�@�=}a���)�?'I�!�)��'��3�ː>�I�
����Y=L��=��v���t��'L��L��_���8���=:�'e*�{X����8u�k(ʱ�P�'hW�����B�RT��^���(;d�C��8��;s>�Ȥ�
�Ç�}N��
�Rg?Y9��H/��1�'^�3�q��L���ǝ{�'a��8fhm�+��S:^ =ce�F�7ψv�C T��J�|g�3O9�%N�<J��|���*�^��XegV|���������a����i
��+����ί�}L�z��h���ש����~��xw�Agl�*O�����H)�_��?&N�Y�?h/Hx��̝�� ���>��=��&H)�4>3�2q��
� ���}��t��T��~�Md��Y��}w�ϼ��8�!��~�N��K�}WnVv���̉5�8x4b��|�ξ���]���<�O��a��_g�ݻ1>k�����T�JG� ��Lܱ�/`gTΙ2t���d�P�1Z�.Zك��������
��<���}����:��J��z��o�Y*���^RXty�33�7�[�0+>����>������x�a��OS��?l���!�᛫��hL�ED�[�1�[�y���d�=�����~J�����d��+%eVz���xN��'�W��_>rN��%gߴS��,�|�Vz�<d���]s���_���E3̃��&��Pk���2޸�+����q!�~���_ԛ���w�=�~/H�;��Y2�*���ܵ	d@�W�+�{ə�E�Os�cp��n���veU��}��\�R����B�vyO����X�WT7�p�Zw�^*�z{�zH�0&R��%y�}9�>�Z�V���*��逃Cf���׶S+����t"�oI��+E=ؚY�E�Q�w���X����uǡAį�_�Ϋ��S�W?_g���$o����y���Snǰ+��5[���$i�fQ>n����7��xo�SFູ�P���i;;4��&�+O'�Z�64!>QY6+}�����!��v-X��Y��ٻyE�:ӛ��#r�"�x�v[���;��7׼���>��,�:r}�dS���;K�.a���.Oom�bJ��`�#��#t���7�g0��nB�V}A{�u�ּ��j!"�YP�7ӱ$;�"R��]\0b\���z��PB�������·��J$��Z7� ��\�a�a�+W%�dQ<N�CʱS3!܂�8��p��'K6���t��X�Z�Μ;V�'<3�������6��������r�Iǳ��b(}�
���Ŝ]g?���iʷ��[�Â|��ǏK� �B��^L�K��[���'�/S�>�.�5t;��KGu�`�/+B�i�����9���Ǟ��A��t��L���Z9��c�7�}wD8W��GܥU��U�
��\� ��ZF����V \��"�Z����#>'�8P,%R�(p!��d2A��R�PE�k��s��4�z�����o{��oT"v��j�Q�*�2��|��K�����@^�������./M26)�ƼE���Y��#ڶc�5>�.��x(m��������6�B+`e؂0��Uw-��ƩK/lB��kԖ?�(]��
���S�|k�,���vm��=�O�����	�j޷,N]z�������Z�{^��/����xQx�������/��Mz}P���L�cq�D�Nl��͗�{�^᰼E��,A=����> �b��x��뛾)�U23M{��(.��z���j}�P[2��Ϻ�ÞJŝ[��#x�p�����{%N����М1VO{���Ә(�,9z�S�0*�J����8�P�����灵S:M�:��� �Ũ��.����V��d5��+����W�*V{����Gk��C�F���`w��F�&�w�6�q�V�gu����:�2yڎ��@�}ҝ�o/2���3BY�4N���*�a��
�,���,��ᵗhz�r�h�Ve��[��#�s�t�U���g�%�k�Yq�PqXVk���h{-;䡂9>�F���A�3���+96(��=kl�����-*��X��V>:)'�6ȫ%-�-y}ؗS�H�8�U���X��n���0;z��� ]F��O��q��7���9{Nzkw���	�w\���Z�5d�5����б]��.�췱�z02�����im;����+���O�Z��NFT�9�l�����%X��dC%�m0�:i]T��6��敯�=���7�2��Bhe��FM�PT�Cl�d����쀃C4����Eb���,[E[���5�j�c�7�{�/]�s�V�0�Q=e�{_΍���F|�����!�TC!��ÙVɎ��/+N�SWan�-Dc�E���.��z����_�U�⪖�P���0=��	z�Ӏ��oS^�����U����ά{mA�����F<�1�F��X�]Ź�({cآ@�y=��e�B�K�Be��w҃�%$;�8D���p��$����n��Å���gQ̶���>o55J�6����\}Ƿ*�kn�o]� 5���eZ4�0a���WæR���^<(�̛n�<:sA&�C�Aٛ��MYԇ|_���߻@̵�r�ܟ]���e�����U������h��0��.�Q���BS\h�!6��>��x:=��A?y��'�{+�od�U�b�x�(f�q_;�u	��fy����F�>���:�%��h	l��(���qU��-��U�I�"=��]�pI���*���*��m�1�>v!Ѫ��a�V��b�@z5P���q�.3\�[����"l�iV��C<?z�gJWo���S�{2|}�(���|3"^��5-2�㽄����W��/�#v:�Q+�*�����!X���|�pN���򭜫�o4��T����|L[����:����X��ab}iWQ.��q����'n^-/eu�w鸺�{&Y�U?->�������u�k��?z0.��3�w�������q5��Jf7��]��"aT���Hx���D�כ���XT�d��Al�X�	'�@��3�)��T[���H!�^�-I��3J��UC8��#t��4�T]���g�ߥ;�z�g�`���2�4���*fTͱ3R;P�C)'���=v�M-y�`�J��z�cQ���J���h�Ky�\w��~Wg�zB9��ː�:'p�L����:٢��%\Zԏ;���fa�h=��9qN���ǽ=��O��\���l���$�^��h�e�X1_Pw>F�B�M͟=��;��4KS����0CƩ�	�Y��ò�/�*�z5��w.���y <7-����/�٫�]⪳JK�|uo��U�)���
���5G�k��ā�q�*Z+"�E�UY�N^t�ECA��/��-7��2���)����sp\�sC@�O��E�c(�o(�[�|����(�<+�����j>�7�sVm��JYO���&ä�-��;�6 [���>h������%u�? ��*<|�Q�5�Z�JǪ�Wp����`����m��l��p�џD;!��inn��C�lW�ێqS��	ꭶ�����5�ν*�����^0b6+މ�lI�ŧ��	��+���w@;��xe�x+�Z�ٕW�g��O ����X���=�W諑�j��%H��u���z�LtI:Y+r2̳��+:��PE<���L:�@_Lh{%k���ǅ+O�^˿fS�n�ԭ�fz����'KkQ�v̨v���ƌ{N�q	�� +���*5�7��/�@#�����L �3����������婰��� t3��0&bx�]�Dg�ˀ�J&{M�N�b��7���GՀ�߭X�'�3��+Vt-%2 |:m�]�q�w��vg�>��5�e�C�vm���i*�t�s4ʛ2�ݰ�ۣ(�[i��vZ'SG����M�=�����g��>�hu���o�˂q�����u��r���}�<��Ҩ�m-ۭk��qvSc��x�ij����y����
�~d>�����1`�XM�+a~eWem�fg�c�g��'�k�m���8�Y�,������U"����v�)���a����y��]�g.պ3���F2%�`CZ<+!�;(����AJ�g�W�U�vײ��Ew���i���v��2�� 5ϝD
6�A�o�~9�����+�;�L��e[Y�ie��}i�V<Qf���[f�:��	|�̝�~�omP9�R_X���ְ8�V�d�[<¤��em�dȡ��^�z�B��:�#�S�H����VMmL�����&�w�Da����qke�3���*x�4����@��@1:��B�k��x��E�yj7�����6]�>�&`��s���]t�?A^��@j�pT�r�͓)�`��2��:W��7`Z�����CX�9�3�F��?��E�ڙ�0ۑ*F�/q�/�����B:�ی����R�|V�ʈ�N�V�Kt�*�Y�#(L����}|�Y�]][�r#^���,��׷���*/�[]o8:]ˊ�
���9����r���U���]����Y�Ͼ�.�}��O����3vh���A�/��
.:
�c޷f=�jǅ<��S�|��� �U��P��1������gh)`0�Z��4�u�����[��^�Ҽ<)�����]����sR�͸ѱ�>kZi>� ��eߤ��K��{�U�s`�{-h�?@���^�q�5�	�n��=޻�ٕ�/�ծI�K޺�ѫb���5��w��ĬY�>�Ds�����{c��v�g�E'��G!��
f�L5`F��Z��]��d+L��0K,�8e��->�z3����k��77K��bܺS�KΡѼg�P�>^����U����~z���z��l0Jy9Y��"��7(1& �S�KS�K`X�o�ظ�"I��6�XK\h���������w���Ϩ�p�{���X��`U@��-wp��3{_پ�)߮��Ϸ�7���]�хq�k�*��?����TO�z��c�`e\U���;i��n<�vқ{���&�z�r�2��!>��P��]�%�m0�:Z=E�s�h�+�~i]͉{Y�/݋1kM�ȹq�@����o~��g5�y?\�g��\�ڼ����� ثd:ݠ��:�<C�hyC��,��#�f�Nb���,7N�W�AV�g�A�ܴf�'�>�ػE�qz^�:������麋�#{�Κvo{��Gxa墛<G��Й��Lx��}�S�u�*������m��J�"J���mp��jx�u��+��<3�ީ��[<*�(��x�Ex��k�i�A:��:�ĪH��� �ʸ��nim���fE��Z��}\�������G��r������m�u��g�L��ģv͖T����:��^��zHk�2��]������1C����ަOZ��'/�hk���ЧU[�X������T�d��BZ�r�*�o�>�Uvk�Z�au��k��+y'8y�����^�FV�p���ב�����k��ah'�`��톼�z���8�ר�qr�s����iv�׭� �ǃ�ԫ�n.�~��u^���Z�R��fsƅ����+;��`��Ө���`�K��U�S�����n��X,��
]�[-�"쵆�d���NH��� ��=�Z7�ｸz���֖yT�!��W����A��$c��{����ubzl�|}�������+��kڵX��H��+o-Q�\Ԓ����!X�������g�Q}ƣ��gk�����0���Oh�Fb��!kmL�9<s6(k]7;N�."��Yn*&oM��3�Q��i����8�M�+��E��v�`	�#�Ʒ�.:�e��<4v40�c��MT���{cǴ�J��ۧ��S�n��TR�j��'��YzS��6�G.��ƃ�Q�f�]قT�o��w-@��ڠ�,�R��VX/FT\�$�jP�oI�	�}�o]�j�����We@�Ϟޙ�9� ��m)9#3�����9�]��ַ[�˽�.W�3�<�.+j�;v��ɣ�꯱*'��3ۭf��v�=����僟+�ؗ\�¸�G�R{�X�G����L{�i�Ӱ����IQ#��:K�ʂ���V�T��-��ʕ�Xz���u�"��l��y(w��b�+(�3s~H����׺ލ �L��kfp�xVI��)����b�Ȳ;ٴt�ET긾;ֻ4�$���5Yr�1v@�3	e���=t��z%��V���4��	��w̵	�z�_r�|�Zb���\���ʶ7��-i������b�/k,t�97��%-QM�x�	�
��J��(b� ��~m�*R��B�t����
�G�P��^W�}�E.�.uҲ����y�c�����/�����]:��}�z�&��W�7ԡ���}���{,�ۆ����k듯(R��߫���u\8��ubG�|��vq�Ԫ�]T�f�j�A��K�� O9w{N����C��Gf��cg�DKf*䈠�V{���� +��fkVii��(�Cp��]�9%�ի�_��uX/��:�y���{Գ/�lGj�X��jvb����^I2�ʖ�ZO,�ó�����n���|t����Ns��;nm׳�Q� " ���W�z��ܛ�
���:U�=k�ݝ�I����
&�;�����?�{NPb�p T���A'��ܻ����:ӻQ:�.:Q�XY��5S�#w[�j3�f��{�n5�G��s{�������5�}���YWR>��:Q��A�=���}ӛ�`Dw<���_��<�xW������	���[P����ة��M�d�e��{����1�q�Co���uGer�v-0�*��5�{n�|��N弢��Pͳ��*gWY�;qz�j#u��$��8{V�i�WU��gX�Ŷٻ�,>>x�h~�:7o /�osC�hʃp��R�-�+*���}J8'(�ɝ�y����Y��mI�V� ��C`����-EAK�h�7ux�r�;8�Y�n�.���b�]��8��ُ<��4�9�OcI��a]mM���@32o-Y0��JZ�B1G���6�-����;�ˆn�q�+.A�W,�����LU;��`�V�i�ϵ��:�o��ZĖ�	�A��%�	<����-�m
�5gt�`��,a�*䕋%�b��`�"E���x�B�T2"*��ɕg)�ʂ���)˴JP*[�
��J�!R��6�r�QU@U2�a�2,�aZ�VT�0.N3k*(3X����AKiPY* Ŋf�(rܕ��5
Ȫ�d��&�[F1C0**AA`�,
��#c2q��D-b�"�咃(�HadV"*U��,ڣ�IR*���`�P��(�Ub
bՃhVAAb���,P��b�dX���*J!���)�0cl��YP"E�@U֬�1R
(�R(�5��ŀ���A@X1VfDU���QR(�
*�,MlQ��V6��
d�QDR�T�s��֢M�)����WM|�#����0��3�MN6��l^we���Ϫv��M�;���DlW��	m�4���"3v�INfm���]�R�t�>�R�)����]o��-*��,�_=7�,e7W=���I�%��d�-pt(fQ3cE{���k��ƾ�f��������\[� ��T��޶r��wV���z!d:7��"��˵0w��׃�Y����-�J�k�4�רz����}���nF3�+��~G>����Tĺ����U�پ�<����#x�8O�{*��K��p����E�m�+�yyب*x�N/{T��])c��a�cN�Gf�I���8{�����#DINJީc&hP�~�YY/�}�wk*�H�E��hN�urBq��������d�:��w�b�OQ�U��tu&�����2��xVDAbu�A���9l��!�K�QG3�I�͸��Z«���=���ޟR|�e	KX��R��ϗ�*r2���#�rm��vu�e�	�@}03� b�}�	�
 1I48g���{V7�+���H�V'�5�L��p�\fە�-A��;$r!�V;�c� J!L�j$J��x�r��Yܴ P��V��!x=��o�-�~S�Cr�#<�w4�!5j&����+$�鶕>0�o�-���%�́�+2���h�`��+�M2<ۻ[�:�����3SɶW8�x���l)H+��t���>Z�+�ye�E��kX�#�Ue�+&��_}�~X��޼4E��w,z��Sx�^�X����w�
m(b��6%Q!0��hpDH��6k�2t-#Z=�@hË�ʷ��J��/��)��U��*���BV�����x�#{��I+3E�S^��`����1r�es�"��s��a���}�d�| �^�x�YLUn����'H�ɷf2��j����<i��%�7H����<9�.�W�~ W>yn���k����Z�}�!5lHK_�]Ԕ�ϰ,��/d�a{|'�~�\��:^�.՝�қ��[R�N�-lw��ׯ1>ik��Ї����,�@;����%e���3j�GJ���W���:����f�1�����Fn]�sb�d.��;
P�{���en4%N�x[ ��n�n��@�!�$���_�c"\,h�;��Ƙ�j�5s��=�1򹎙򡕔��zgS:�[�0a��O����!�C[W9�]E�;>������z]a�Μ��~�I�61�$�(ixE�tKl������U��+�X�|b�5*�/��_�ٯ��n���'�Ɨ�t�R���;��d��7��3��D�{Bp�b��v�����ɤ���״�3Vu��B��v��'�pi����sTv���ؽ9���u��L�u:�]�J�8�1M��a!w�����U���{S
sl��t�4�`��C-�[LDy��5N�����M��mQ�~�U����*����|��dS��v����p���a�t���Z=;*]�����1���Y�x�C�^�'O&}��k3Gf|��}\�}��u
���rrc=���ܽ�βʻ�g��H����J�M����S'm�KD����6C��De��L�f����̩*Fs9i�x�#篝����u�uo�K� ^�y-�}��G��}���>6���^1b�;�Oy����j�W���kC���%*3K0ҧĳkZj��o����>�l�ꏃ��_����m����ۍYoV�j֥�-�{��סY�j�׹[g�aP׶��9��mz�s���&��|�k��+���UڵO���T������HU ��{�X#(��<+�M��F��#ӍS�Kٟgf��y�yf��𱕺���oթJ������QGl��j�A�af��<&�F�z2G��Ճ<�'���u�#,����Iz��+�,���_�v����=
�]~#ݙ��`b�M��}IeKƈ5C�ht{^�q^.]��c7�#;�]r�6諭���հs55/��fO9�|����D��#����j�>��x���r�/oe5I.Ɇ�m��acj�k:�V���Zv{j�t׾�r���v�����2Vγ�fj��+�6ͪl���(n�#�[TSiQ��Nj>\/x{g�(���n����[ST{_�vX6k�kܟy�YT+"���u�Vkثz�{���=1����R���y[���mʮ9����C�����= ���-3��b��eL�E̶+jV���B�Sc��k*�|��LZ�@�o��z��iv4W��7�mA��:�u;ْ�5��<��[�� ��4�\/��:k����+je��1�Y��:���\X�hz�,���v�}M��N�-�tcq�P�,r]\��mB����}�ɓK���᳦f��x��k�i��l6`ǖ �孕	�\�=V�c��b�S�sٰ�7hI�\H��<�ܨ�fZ3��
�K���b��<X�b���QOUe����ܮ�����c�������+��dgK�;���D��}Ks�G'�������`0�N�����|�'��.�̝e���e���y��Y�w0I��˿��cYJ�m:��=�G�{]�v45�h�;+}P�S��D�qJ�+im����U/QI�C>�S�?o�jN~�ӏ�[�y��5oZ�9��m�bo��K��"���K��u��_P�޼��]��\��sFZ������~�Z��|o��_Ve��o"�7�����T�-�~�ޝi ��v��\�2Bs5��Y^u�[Yr��Vϰ��<�͊��p�}C��
[:��/d�{�\�׍ӷI�jt��֤mΠ�����鋪mq�* �Z�7dө��SB�S\-��ǭWR��	K0�;Cum��w��BF��|����j��^l�h�j�r�gtT'݀�>�;T���o��Έ���O���=�Bv�U=������<�m�h	M�{I�xo�VNѭS�V-��ɫ{PWr�|�-Y��5�	uW�ϛyg� ���l�+n[ɧ����L[W=�y{B�괥?6=�(:����3Ws�[.��AS+�@Q}n���|P=oW�,��q�T��U�.�s�GQ�_1�W.��M.�:�Z��ՇIg{(�Q���S;����kR̰�{������j�7��iž��mI�'hF���Cr<�b���|O,��H�|r�񿍩��Zgw��k�<%�㉲)gh�E��[���PX�2ѕ��Q8��W�g'�7h��^�.��v����aI�1Bs쀳@�t/��f�Y���+mD����y�7 �������m�*4�e�}U��hVs��>\�?}Y�̬KN�Iu�mҏa��E$e����Љ77	�Z�����(@��p�^.�'���J��c�;M�L���j�d��p#36��G��ٮY�Wv���s�Y��ꔽ�?#�滰�1���h�O�ʕ�6�y����m�NC��7=�gܴ<M+K{�u��L[[F�ի�В;T�^�fݕ���ǟ%y�_^�d��t&�K"߫�U�޺'Ʀmz���mؙ��^�Q̴��7'Ϻ����Y*��H?w�����g����r5�/�n����.
�@�v�w�����^2F�-�7C��ݲX�ң0Z�2L�a��iU�(�$�e��}�	G�^��Vn�û��vVELE�������ߺq�V}�u�u�S\�/.�"󐒢0a�4e..��m���k����ꦠjz��1���o��;;h���,�~Sq�����m��2�h������	����a�~�/���[6f�U��G�mQ�eS���{�w{/�$[��/jm?v�[�+}U驟���F�|%s9�Z���[�� Ke��U�^�Q�ՋVϨҏ2}.�B}��-{��:ɖ�U
�T��&L&����[���f4�x*��=*C;F�lAm��"����HŨN�J��kw�d̍����)�j�/Sn�iW��=�����.�t�G�{f�������X5}$%S�{'â�P�Y��V����<3R��f��M�m|���S68��n�fzU\®x��-C�N�y�Rv�|Րm�ƚ��b��ͯ#,�6������g���x�篝����Y=�v�q���e����ֹь�s�OP�b��W�m����>�|�Q��aY���WJ]��b��IG��(+B�g�$ƭ���?e:���*�9Np��V�6
�E|����m��,K<��y�5f������՝Sd�8�
U�ǽ� �%�������d�ܣ�3v�T���X��ld�t%��>�^R��m��y@� ]'�_dȼm/���aը��UU_|�9�~�~�s���G�AJ�5�U0�h]Kc�ܟ����_$Q\h׌],郲u���>�N�S�N����_z�^j����k�Tw��L�̜��x����!{WWe!�.����~]��)n��[S�ep�]������oW��[5ڰ�!��ߧF;){2�87�:�xU�ӛ]�݉ٝ�����Y8�S4���jM�o��{���AqT�����L�:u��{��.�s=�̂TG窳}ʎO3�6���bf�2Y���#6���i5�[:���S���,2���kMy�cY-�.h=x*�u�����o9X�ǪO{h�����6��&�hQ���Cv(�m�����^읕�fn���񑰻K��NX�|����v}�7��̡Y驰�!Z�Ɉ[��F�l��-�z�XE����I�~&�}���T���H���r�W:�D��_�c��П'Ζ���\��{9u�ޚ*8�%^6��[2�Tu�#�v���{�r _-6U������w;���|(l�sO]@�0��R��y,�&Q{l�E��*I�t�fX�^���^�-�мpR�~�磌�%��w_D}Dm�N鋏����h�9��J_��q�"�����I�:����!u=�)��b�hlp�{4ά��3��/i�	�w�&,���9����^g�^�=�Ce��&��A.�Y��Z�L�p�gE����2�w1R����i�JǤ��5��-�w�t��-,�j���@>���V�/d�EZ�Z���F֏m�������h�7y��c�{H�o�{E�@�ꥉ�G�>]R�ua~^��{{�<��\]����%��=�[��mIJ�˼�*v^���_�$�WR�<��P����)�u��^�'�-�}U��m��+�ױ+��Ur�י�Nߘ�����:��o5�J7��{⠃O��k��|��*kc�ڣP�-M����9�嵲�i���VF������W�U��ܩ���w��m����W��-�ɮ����^Ә'�I�`�C
Y���8��a���:�vv��ӗ?����կL�:���O�U�q���������/b뾉�J��P�Pn{��+� V��J:�o�����u��;n����}������f$V�)���8\t�u|���ꊙƒ�{��ݲTs�譫9��_}�}�|�D��ݚ�-�� n��q��1�Ֆ�e*�x�n�o���+�!e�}7��%*�s���*�;<6��M���6��+�N�$���ڜ������m��q�����{q[�����<���6Z�Ch�:�5��:�-+ױF7"5��-�;�V~��΄ϯ����û��צ���&b�jm��!�_KCbc�[�e�w���һ�7�;��zX]'Vf��S�j�l�d%,5'�Z���~�<5+<+�uz�����X��/2�-h;�&��0�lN��@Yh�8px����;��C˕����k�	����m)G��iҲ��6�p+��{�ќ��V%�������.�O=���xx�ơV��[�ێ8��hq�?#��@y��^��ib|i[K�����j����{	f�ϗ��	��|:���r�	b뉦V?L�~�1%�Er��''���Y�9��Z�*���	���޴�����:4�#CS�r=�^�M�.�;��]�S`�;:S�.oAO]݌�$&������V�}����ƧK�e����پ���{'��l�E�E��vS6%KW���0��G���B;9˶ݠ����'L{�wmZ�����D�s�l�}��ʂp偗{�s[��#���#/!�k�������$�e�:]��5�ϓ��*����щ��)q�ΖA�������ġ���j�i���A!�=���{n���sf�,�O��X=0c�����+�U�z��t��^��;Lq���M%MR�ze�d���3;�o.��N9�q�H�0���d��\��9�r6�X-:έ��2����15�I�F\l�$}�V#��E��+�Kgi���c�>%�X��[���/�ל����M��dk;F�s��[4�Ɯ�7J2}z^�1�Ȥ��r�F@p���n6Uaz/fu�1¡����A�.k:��K���ǫS�����|
� �ݏ{9 y�x�|z��^}��9U�"�E��'�Q}oBF�+vݕ�p�AA8XTg�������,A��4=fhk�ֳ�J|8���\@�y�X	�N�!�n��a�.$��Ŕ�g�;��1��AO'ؕc�`:bp�ղ�+	�u�TȂ��jnԇw�K sF��i�6�:�6�|���.����@R�`�TNu�]�!�v��*����k���lpf�VQ��386N!�+`�A��e rs�]�,s��m��mL���TW\}�5й���;�h`s����#�M�c��Ք�;�Ӱᚳއ�:x�ή�6��2jܮ���j�i*�j��lk����®�r�㷄�ԉ\���4Jb�svpو��춱C���g"�$���˸�)g��dH)��+:�0�m��6�K���>�Z�t�5��;�N�7� ɬ�=���l�h¨Kf� v�y�¤�Ջ��3w;	�7D5h3�׫Z�}����#~B�RR��[��������=F����=�M���\ �V���i�	�ۣz�?�����>8-��ȑ"�j�`d�HesV�,� R���k��H�����_{��,t�M�G��Ǝ�UF`��o�s�f�_����<Q��˨n��WX��ш�/��7&�[�u^�]�Փ����܌�h>�֠�Dm�N3P��qT����;�e\�qnl
�O���f�&��}{�@pF�>3�*ZV�ӥC�H�&�ٴ��#�)R�۾>=>��h�AyDXZuS�p�ݏ�&J�t�,)S�Y�~[9�o{ U����ܽU��~s�����S�T��F�2U`�*�"�a�l���U�DQA`��0E"�(*�T��X�Y
�XZQd3-�b��R
*�H�����sAE@U��Q*�Pm
**�
����1EQE�-(������AT��QE���(
���J� �+۬�JŎl(�XT��!X�rT�"ʕ3%**
eB��j,D��У ����PQԬ2m�YYDdEfa�sk��(���$*6ź̨�i++Y
)+D��DX��`�W!\�Q��lT�J����@R�P+T*
"��TRT��(*�&��k��Db�+QJ%eB�[eaP�+V�%�HT�E�R�DPY)lR*�)[�� F}�}�,~��}�%�z�=��j�%,K0����a��cc�ĒMR�O:I*ݧ*�h	����8�r�������37��'V���0�ו��H:?�;��%~�0!��_Fn�kR{�w�[��wzyO��e�)��t�2��8׸�߼ս��gؕ�e�\��}�e�9OiW�N���mH�Uw��M1��1��e*ܖYCH��תK(�(�o�u��W;���2W�k4��D�?1����=;�;ӳ_��~���ǈίsE����B8���UǼ����}�9�N����ˑ�@�cA�aUkcu��<�.�����	\�T�Y��m��nztސ��Y6�uf^�"���>�Y>�y���ca������E��Δ�������]����K�����z�{����ml��S�(����E�b�fܨz���ȵ7�ڝ�I���I�7�)����V6V�R-{t%ba��mAe�mۜg�4t��q�����'�z@��R5=��|ը4�V�:�!����%�Q��G+�����ǹ�f�W%�ֳ��|L��oh�\�]�K��_��x�뎯*9\��N5-'L����E�)�p�}�k9�Y��9a�.�>J��� ]c���ZK#���gd�M���^�d�j�Z=tU�At�=Ζ���ӵ	�k+����������$5�.�X�_�o��'�3h�͚���v��Ŭ����ח93O6���F��|����N`��%�O�/f���&_g�_�{�x3;T^�%q�;����d��Z�.Y�Q���J���_թ&��3$j�So7�8�G-{!Ͳ�R�^D� g��g��t�\j�ŝ�A�L�B��0�n�z�c��P�Nڀ�����^(o��v�܀h�T[]��k�W���W�S���sT�|�-�z���VkO�Bh݅{�(�
�I!�������^v���k���e]T[�I�Ԛ�X�ߟP��<7��.>�OJ��;������ҵ�3_���[��ɫ�5�J�����A�Έ��Ls�~ܪ�8v���n�ҪݢSk��<]%�{���_�F�k�zf���:y�vOM*�K)�*�Tf���r��
��ۯB�N)Gn[P��ήs*�yQ��^��Ϋ>����<{K�5���nI�tq�d�+{�,{=�/-�C3�ۚu�񇵜�v�n>�8{�u��X�� ��!��1��>/��h��9Q�sĎ�|e�����Ǯ��(�d�JlG�^膄�J�z�O��up�|��� ��R�A���b^}�ؿ~�Ͼ��-�/��e��7-���s!�V\�ۂ�(7q	66ͳ>>El��3lh��ی���}c���Q�M��mT��K���5;B��FQ֡�i�m��KM��05�{�����A�y�Q��}=/�>���]��Jh�;��v=�O�ê��� *y<�+=�M^�IU�����&�z�m��N1���P��Tr�վ�=Zi��E�Y�1.���w#e�B+j�����ꄈX}�1y
t�T�boe���6ϔP����m	^�>J��{~%\��n�]�^�b	bX�J�m�}��߶��T���,��퀲<K��z�U)+Pڈ�MƅΨ���qR�Ǫ�쪛��_��l�=)1$�쵖ڸ�2j]�nzG�Za��b���&z�ūް�����b�???j�!��"�ґ!5�
��I��x�� k�h�������iu/m>�S:�������W�w\�}���h*�����m��r_$�h���lmT?$|�5X+<�u�q��P�rb����v�T�v|��kE���Y��x�6�|I�2�;���o��P�b�ޅ�VWA��<����<-��S�W�UUU�_���-1[_�:��/+�����W�ݪ]K����O����9�>�������9��Y6׾�J����Ur�ן��;�yŨ�̵�$�j�=���v��a�U)�+ܖYC2Y[>Ƽ��^wJ��Я�۴��
'�
������S�ޓ~sJ�[���V#TzO\�y1A��N��}��c�3��E[����wT���^��j˔���JFQ�� �A�3��X����^}�3��o�#��j�t�;�"Mq��H��6N�*;�b�������ݔC���U��t��E��6Ϊ���u�|=������7����!���[�E�n���e�nUP�;��r��"��N�J�S�H�fGlf���F,��PY,US;XmU����M-n{�3/���>��s���)�j�16[%,��m�b���mr�^z�W�z�d,WuzT84S�h!|����1AO/N����(r9�v{w��yF6Kd�۲W|�^o_h4�@��G�hʝ]lo
�e�r����7ˉ�@?JMM�� 륈�X5��.Q���{]C��ΫG9۸VH8t�E�ct���S巫����te�3�,`.臍;�����f9�6�$�.�F��dm�ې��k�������q�����,�""-Ńo�H���󫽖���J�v�XF�a	�0[��}��E;���Y/��b�W�_�7k����~h����:]L{��/��z������z����^���H���������H�]�>�՝圼 �K�yl���J��8emy�v��C}�vy���W5|}��3x�p^�C|Q7��n���kS�clP���[4��e�{�bݺ2W��ד%\~�y*�w
QKfn�[ثMI�CYUi�74�­Jv�ȽUCu�S���ȳk"�nν>�őL겞=&�4��6wa�C�b;������4Q�h@�^���a%�3��N�=����t���q�:���s�ӊ�۫����??V���T��n?E��C~C���۵ë��J������=��?pG��	QUB�����S�����|��2q��¹����a8�F�7�,� ��k��(�.�����c%�DK�9m�-Z6j��؇���$~1I�{�y�Og�,��
Ѵ���'(ܹ�c� �_}k��<=:������猙��_1K�o+�r�KE�'^t7t;�W�W�R�o�*.�dz3���ׂ�>�p�Z�2)��ZAG��m-Ƥ�	��y$6�n����R���k�`#��<�.���Rm���Y\���k��Ka��q��bT�h��ш-�,�5�&��*�T��������)�*�`�e�/���ǹ����T�����`�<�
�I1{�ά��������`�Ru��w���/���m_�{v8���IE�#�s�+ԳiT��t�+~�}6���Vy�-bvS�q�upr!N�%�X16��I�Ǵ��V�%���Y.����f�\5�1��Ӛ���l��y��]r��Tn��	�R)#*�l�zԂV��Oj���_e0z��H�ݜ�z��y��ʃ�PTy�ǼX���v���z���N%�)Pku�Y�Z!m���q6�Z��z�ү���N�=������Vmy�|&[�mѤ�`7��'�|���A�u���V��ZEܥ]��<���V۳#Kf�A�oYcuE��:è��'+ki�7�|@���z�L���%4Gג[����8��Ed��ܡ���b��U�07�=�rͨ�_N����o<ڈ��R�ٍJ}�sY���q�!��[��,����UW�U_I�S̝�������vڋy��Z����F�vV��Z]�Ψ�y��)9R�m��fթ�P[�j�m�ݡQ��=8��=��S�n��w��ԕ�:����쌼���y�2��.�i�;��{}^��t�K�x�y��ܤԡ���n[4jxu7��FT4�#%�W-�l��yR��{�[�7���fumr�fҷ[[wX��Rۏ	K��,(n����?p���m��{�_JS�fJ983�7��l���}=��m{;��0�5���i��m��)-��֜"��Ӛz�?^��%�k�w4�{��� �}��V��h=�}�HS�~�k7�D��D����ߴ,�k{~��yv������Yi�>�M��l�Q��(����P���Pb�:�u;ْ�G��fi7���[3����^�u	�����,�h�B�J��1�Y�<u��Me{�r���d��p�܎��Ɔ�Ub��ZN����R���)[�;1eji��/���}�G�Y��ޥ\{:��
� jaa�M��s�����kgL����Q�vD[��z]����_UUW��^���ۧ�VӲp�؃��ń�l6�֩Ʋ�
�4.v�M����(�z�ъ�u�{f˵m���F�
�i1Q�+���H�I�E��^�.��gNn���^f�%��qj��e.���ܘy�PO��`;�l���A��{tU�ςwˈ��9�Ć�)K����:��^�V�|�L����5�n�>܈��Vٯe�m�,~i=�]K���ܠ_�d�ZB�Y�r�W��6�>U^����6��%s����߈^s<K���s��|aU��M�Vv�l;6,���b���Xِ��c^pd��a;��(o�wo���`����I�ٳ����r�uo��۬��z�b�<k(>w����3Q�5��n^&����7a��*Y�eB[cP�l��3hxP��*��d�&��%�߫�W3Sqh|�~;<6�t�;�6�|ǚ���8f�;[%j=�L���\�|sX��N���tl��1ĿT�����=����,�s2�s˼Geﮔ8n��~��-�Է��Ǝn��6Y6/2ӂp�2�������fk�q�V��^�M���ܐТ�2Y�� $}�3y��)c^^˔��o5�6u�XP�vv�%y���}��v���}"J����;����njo�\�6�}2�����v��̭ţ�F��.z�7�j�z��Kp9�{MZ��P�P�m��*C<n�ϧ�ݴ�?3��ٞ�S���z5�vL:�T��vkA=��έ#Sb��,��1��,j���m�Fңli�G=�|	�&Ab�m�X�]�v�أ2�-�Z6\�*_��33�yX���;Y+"Y���"�R�c)w��So�<~��6�ۮ��ňn��5F�M޾O�׿���W�S1�f�%忓~v2�P�缚�ǢOx@��9���w�����܎ס��.-�?#T�>(�]���_{�����y)X%{��.�O���P~;=�ȥW5k�]��m���L���&�7K�Q~�;|7�Ϗ���5ojr��+E�}�Fa��?S���V��z���>��{{;�RK��;BY��atd�pF�����DY����dg�i
�82���4/yL+%��T0b��N�f���(�����H d���b��WB	��l�1�]��ݦvî�Ҿ�"�$:����y���h��IƬ�{p2m��M(�cfǬ���Ų�i�T���G��Y niVT��<��(����s�es�[�7=gv�ױf��j�hW7,�Vn������M{:�_��w�s]�~��{}1�:�l�{$��H��g]�����Z���x��?[�[G�~5�����|�h����������n���v����+�S�	K0�;��7P�Uy1h|k��44�.kH���Z����
�(i��*�3mm&��a(��A�e�x-��fIȃ��b���.�s׳ո�e��O>jI��cƖ�B�Yl(���vf�TK�S�+EkF�+�Ym�=�<��BO��)��j�ɷ��}꜌��@M{�����|�Hٺ�r�>so���u�N���fA�j�<�kҢE����s90b��wR;�lf�z��]�ƞ��߀��y/J�X��ٴ����Պ�F��2k����93m.f���W��ʕW_5o�G�0k9T�+kRC�q
CX��ϵ����-Hʴr�'�e�v(wm�d�!d�B޽\{&/,���U!���\�`�|�x�){rjrm��X ��osE��N�[�٢����r�@cwPM8B���X�ޙ��E��~EX8f5����;��H�2t$�/��v�"��Qe6�
}��"Dᾨ��f&�l`���;�(ow�d��h��1)��8!ѐ<�&7����_2��~ ]&��ƞ�ȹ�ڎ�`:;Z�_pnUp������B3ܮ��4���Q��ݦ=6o���v��;>x��3u�獾G�jx�B_G��"n��nӶޓagWq-�b��&�T9��J����}�d��q���0��e�~ғ;�qgF�W�o'>�����,M�D��m�Ӽ�������Ճ0��{���4Q[^�T}%����ЧQY[��Yہ�@,���O6;��{J;�������_�KWJ�V�o����¹l<Tӕ�k{D����Lŝ�h`$K]����5n.�l�����>�G��ÕGn{Y	쁊��Ќ{+�,��(G��)����`��{�����(�#��ѳ���İ�.��u�dWX�U7Ε�ӫt!�Z�@
Yc/54gd�wb������V�F.k��45�.��uQ���� ��%�+*���nحғZV(i�W��RR���^ ��3Xw�:Ѿ��A�B,����t�����Wj��'�s�yx��ڴf��4͔������(A.&�X�X���^x�7K>
E���ѽ���7[�m�A��Z���Pa�W��-��7��p�
�����x����(��%&�;XĻ�K����@�CU�ğt)-'�{~�}F����Q��1xJ}S�©�@Bw���7���O���+��7PE}�k
���W���ְA��bi�a��;�u�p���]�$��c�={0�a� ��&U6y�"��L�8�2+����<>�"ʻ��;9΍�pH���g��<�Uu�F�-��0�o;o��"ww2�fX	[� ��y��"�������kyJ�B*���5k/��W|c U�m���y�x.���]���)�R\x�E��`ɞ�Bo��s|AuD ��kSV�'F3��� :�>�N������K�unj����W&C��� �j[H�2ܫ��yB�1�=��U�#k˶�R֏�\=�w�săX�7\�_6x��Þ{_x\0<`���ѤRi���e�bZl�P��R�mҞ�]8�@F�{��0X8�&�2\v���
�x��N���9����pW+Ni��Vrg~�JH��e�oZt%
��k����ξdnE�N2j���v3iIY+Xm���ʍM}Z� �k|X'���ռνGbT�+�1ک����V��2�n����ʝ���a>jQٗL��I�-�s��>󜷮����I�fI*�V9+* �U$Ų(ArT�l�b �A��]j�(:�3���30�X�kDR)Z!TjJ����J��
�)b�,Aj��̶�3U3��ɘ�J�օeDX�
�H�aP"������Dȳm`,�32B���X�L5\�HV(�
Q�QlZ�+�b��T�f�X�jA�W9��$�iP��ʒQ�Im�3ea5�TUP(�B��DFd��Z���VV�əu��"ԊK�P��m��XJjh�P���3C T+�(��b�ʅI��ŁR���8@�Me���	�d��R�
�e,���Y\��3#�R"As �T�ڬ�j)� ��5!���3d�
(~����$�3F0qNekϬ�,'����U��2f�;{C ��/k��3&�_Sjw�1��>�F �k����7��6�{�+gV��E�L��S&[ uz'Y��V%��|���-�^{���[KK���ST��u�F�a	��H�I�OãuY�	U�o�,���t|m�J�R��Ք�臭[Jy�}P{�ꏇ��Ox� �M�'Sr���~��{=����p�8�z���Գ�S�=����N>�cJ}L��7��gSK��Y-^��+��e�m��Z�h��Իi�-��'O S5W���W���z������f�+�\���%p�ma�#h��Dzqc�=}���q��(�m���W�N읓5C]��+�;k��U�U�yf�8�V��\F��j`��Ӛj�\,�z��ܷ�AC��	|����od�f���d� �:>~:X�o��=�<�$�s^�	�ګ�vȡ�T�m[0�a2i��J	ȳ�;=�zz	CSLj1;���ř���Y�5<'ܮ5�<�"�K$�J�U�}�a��k��a��@�/Q�a;q:t�j�@�y|1������!Ǚ��H6/*���J��B���8�T��+�{]�2��x���[�����] �5�vU�m�8'{뇡0nWq���+wv{�rUos:��v_:^��S5��ٙ�hJ���UUU�n什PL��s����}��>D��y�iW6�<����(Lݽ��d�F�C|�:Z�uL�A�W_�B���k}���J����7��+;�P�;W���Ö����6ĩ�.�����2-�垅?�v��UVm���S&�����u��3/Vv�p����)��0g�Z�m�3�*3182'M�hMDm�Q�W�)=�������6,%+L�1�=�	dϓR�P�b��K�mz���]�h�jvȍ�d9Q���5[2*�����c��f�@�oq�R/��ĸ��iw�.���ڀ�o?e�����x��Ov�c"��}������d��?#K�G�K�{i�A��e�G��>G9��s�b���c�����������ȼ=G�_�z�T���a����}B�]N��Q�3U�ثW"��T2�ݍ�ů��.�F �p���K�Uؘ-,%<k��oW�J��U�;�x9Cv�t�1�!� �υw���
��;oB��2��g�P�0f�o=���#��>���\�һ&�s�W{�(��J-�֥�����&h޼4�\�+��G{2����������������^5#��w���~�U:p������{��/������J+���n>��9'��/E^�I����n־�,ܺh�H�M��5'�^Z��nN	q�o������Y��[Ggo�wx����].�~���dI��aUR�'С��͌��u�R���Z�rߦ�߃�[Gg��{���q���VGiP���/4	��KZ��M��5��ڟ��[A�&���>�{��Ŗ�?��R;��`�j�	�גtvh��%�h���6���+/_���&����=mz�^��-�0T.u6ǚT��}-��fB��|:x��GW��~Θs��ykS66]��r�5i����}�[�%����tX������7͇i���K�e�r�)w�ء�&LL��v!������/V�5~nٷ%�~%U,����֬#gQ����s��i.�J��;�bZ�`�5w{�溾 �A(]+xf�m�3��wSM��mⒷ����E���q���cF�R���s��'��=wdh��2���-�
�����'w��,�0gc{�斦����꽘�L�f�Qk�ʺ��R�����(V��ﾯ�Ø��_�>�އu��~��=ɻn|�}sOT��z�X.��5���������S=~�e�^<��Y��G}7�qo���ib|~G������5��Ժ�{%c��l|=����ڞA�=Eo݌��{�ދ=*g�rR���3w��^��I�*[�[��
�\6m�m���$����E�N�ï_4C�7P��C~wռ�Zbٹ�=��g�V�Df u� k��>l-M�A�]��,��O�S?���$�ĕ�,�wa�C�,�w� ��B1�EM�.�$����h��<�K��>��0��~��ұ�\�
�����ɅV�M�K-����v�u�[nr)�/i���F���W�`�U��� �Ƚ�铫*%!h�{��;���]��[/�V���7o�k�#�Ϧ�������4��w�U�3f���&��a'Ge�Pݟ2�ĦӰ<��.6�ɚ�0�1\'~@�q\��*
Xp���������/#��s5��z�ˬܻɄ�ć�˥ʈ��d*7�M���n�Wo�\�̸���\i���5N�٠Y�m[x���*�z�:}[\��n4Mry����l��着���2���lN����O�2'r��d]�[U��e�
aT��r��\���}nuo}pW�V��mTd[�1��d�lU�Pi�<5ixbb�Q�4�k(+q�TK]���Z1����ؙ'ZO��̃��P��М���:�[��k-Ҙڶ>e�Ah�c,v%�n����,e.^���'v���k�9OȧQ@�q��k�XրL��s	۸��'�s�cLV���N4�e�J����+ږ�dB�l#Y��P�E�
b2�m^�}���^[r�|_�3't0��׍5K�V�1z�(l2�/J�W4�ڪvwv��
�s�O���Z>�ch��R��J���5�b�۪��B�ƣ%m�E�cQ�'J�@qnz��o���T	P׶�rךB����o�yoT��p��O��ﶵC�v��(�ճ5~YC6�n�2-8��Ϫ�P�y욯ٌ��
D<��I���u�VM\"ā���~���bg�k�1:_ Qe��B�뺗v��W�S3�ə`��|��+w~z����<���IJ̭�����:��6�_^�n-0yoU��:)4���Wv�1�ݷ�L�@6� .KKk�v�5�f���[�Z�T�w}~iP��F75���whfKz�>�%�0���q����x��4�f�/|�|���U�]4n�f*qK�������������vD�6��˻ܐ�7���T]+i;�,�a�s/VT�j�P�6�%��7��M��]��;إ����io�򭣽�{�L������G��]�͏�w޶xyߡ�GZ�h?}j��HS�}������@y�2P\�߁}���C.�4�Y?\!���n�����#���F	���>ۻ�w��Ɋ��D��-O�szu�5�n�Sl����1��"خ]Z�'�g$ �rW�5٬��O��U��P��$�؆&��,�G��,�b^��R�Ԥ���r�wR�y��%�׻T��6K�jb��R���]���"�V1Ij�����G��u�[�<M{e��Ҡ]�S�Dl{O��$el��g��Ε��W>
{�^ �+*�-[�������w��9�:�MTI���:7`f&�|V��\Q���J�֋^�Ŕi�s���X�S�W>̜�>�Fy;��Q�zG=�d
ǥ���V2���רY��Go�͵��s��$n9���]�f��Vp<��f}�х���W��w�^��g1���qG*+P5�-n�5�ְ��b����ی���\����Cd��@H�/�ױ� _�R8�u/k��:oSɁ
եɻ�媽^|���f�{��k�eN��^�=�H�����bDl�'zYwA�[Kҳ�:/��Uk��2ګ��P�(d�l
ӵ�����O�	T݃�Bj5�YڋQ��m�U)lW��F^y[>ԇ�,u�C�8�V7g^�,bl�eY/iz������ܸ��m(���)�ɇeH�Fŭ%�=m�}^)��#�i��`n�|�{��.�f���`u7�v=`���z����_�7^=]��j�Qκq�t�[(�����|�y��sVZ��d�6Q����W�,����2�E��J{��M�o��� ��جdN�B�-	!څ{����n'WBz�������aK젷H���3؟b4���	���V�:��X/R�k֣x9]iA�E%�||:��q�/]�}��%O����P�לݴ`J͇.�Q���9��N4���pw�L�����x�n7W�8/F/s/GF�Ј��_}���g�(J�+w8BڦK.�a�-��\y�u2�S1�K9�?�p�]����a>���S=�3t�ڦll����|�a�Lx�l�%,�jQuV^�a��I��Z��ɛfCi�ۧ���d�U~/�6�8��ueѣ���N��%u,�U2�{x=+�P�,�~(���X�]���_Ep]C���ڗ͹�Mw�n0ť+o�vo���ޯ����#����Ħ��xH�R����7���!ӌh�A?�}x[S$�w�c�Q�G�Y�
e\���j�8w�B�Sэ��3Ք�}[Q���5��N)77�hi�|��
_�n��Nl�f��/m?R��;<q��U�eW�NўM:^s�u���t�܆o���[>�Y�-y�B�����|�B�NЫv�څrsm�P�[^��5�'�Gq�J��ګ�D.�=8���d��؋�c��,���5m'\�a���Dsq�ދc�5��,�jo�©��K���7�o���u��m�x޺���evP����-)�VnC��6�Ź�pK��K�^څΦ{�hn��a5�^�U����}9Պ' ��	˧%/�*����­����}�W�rw?q�=K17����׳�5U��t���	����u��}tg�9�h�;bY�������i�;�t{Bl�W�{��ڮ\��5Vk�Y/$x��P8��r�!��Deњ�^�[��z��5?��� �ʵ}��������.�N����үe��1�jj��+�a�Kkɤ��i�Z�WzD�P��4�㷆?�����κi{�n-y�M��.�}���^�+{]���-.�\2\�1Y��{�.Ƿ^m
�}}�HS�k��y��]���f=�W�ƙ��V�w��r��J{�f�Ac���O��C[��F1]3ع��x�U�e4^d+�ͨ[��D,:��щ�'le��o�/�h|����#�޾{۴��4��B�.�5mRq���
+$!�nIvZ�.]�Q�1:���k����I����>j�������͑
�m"�3�����;�5��J�eK0<P�q9�bvӱy�1UY�\�df�W�*���dj�t�u:��޾�v�4�ֿ�Vʽ��n�+N���o�{��wu�fz�Ňs�lU�G99m�:��� �z�Z1*��ڷh�O���wC��ei+H��
��������o$��{�eٟ����'�8�{�=j�J=X��Z�֬�{	�T�%�N�: �<����B�z�r������}��[��^�Բu���w��2`� �yrg��o��t���>�������"�Z�H^�Ի~c�AΧ+x��׸��eJ�eu�
�K��-�5Cv��ck�V�4���)qn�J���t��&nON���3Z��uI����}��U��l_t�8��L�!�ߧJ{ݯ�٥^�ך7YCJ�R�,mG�P�ؓZvL�m�T��ܭQi񥢗�5�Е43Lb���p�/s/VV5-�b�)gdE���|����'��f�{�v�_W'7�4����{��g�zM�\���p��^<j����ݣ�V��i�n��c9�{�^�xL��_�v
��FgugtWӽ�A�)��J��/�����[6�	���e��_Uj^�Y$���,o��r��34;�i:'d$.}���u��1^�}9�{Yf;q�r���|-�7!V��F:1�SM����&�#i�3���٢\UvF�a��E��8F��/T�𧶑�C���Vo�����,U�<�֛ ��L(�����>~�ǥ���5ػ�oM�a�&X#�i�n�딟Y�j���l唐s��Ќ̽�[��_M���}�G�B��O���]���{�p�9�(;�yذ�5;!UcF�PTm]�t��9��.W�^��V��������:�ph�>%qvMS ~�t�Ϭ8(U�#�O�&L�9�X4�\崝c�M��}Z:���jdor��G��6�3a05��x���;����C�Қ�<��i�M���d��ϙ�7ܙ����;uʽN�bL�(qaɽ|�c)�	���XV[�� j�q���;U�7ܦ�R�.��Jb�B{�6�b#�=������3�:M�&V:boIf�&f���Ɨ���t��O޻�9�~���;��s��\���3��9��z�4WG�eJV��XLѧ��k�x瑺fɵAg���E�&�^��&��0]�����p�C8^�ꂱ3��m�j�/x_V"�hwK��Jv�F<�Jɘ�:�N�MRJ�;9�Z�f:��j<�aͶ��f��o��jDdY�2�,���"3�J:�I���l�

��E��|%D{Sާi5BY�SF�$[ZJ���J�kXY� L�+Y┻�zx�s[��s�j�R�Fb:c��oa��=���7ۏK�y�y�Hᘏ%�
��n�:n����������5oU��u�*���b��:�>���u;o���h�ʶ�#��kk7N�QCjK���f��4쟶@۱���7%%���:�$m�]�w����i`��w�X�ƮNݏC�����&Q��&T��$�s[�W�[��r1�l֑��J6� �ژ1�F_s�5p���AJ����}s� ��$�7/� ��أ��I��9�h)�^�z?���[�E���5b��<�Nf\S-����g��wK�����wSۀ#��ʝ�X3�y"}6F�c��o��/H�5�!�o=`���Ai%���`�س'.�DoָrˠM�7�5���RY�+q\�<�gڮ�p�i ;�#�޽i�XӖVr�=�k�}
d:��#�����EpCQcʉ���B�­��	������-}����#A�Ni4��X���I}G��x�+��X���r�MY\�H��<�Ӯ\��o� �݈�k���\��ޓd�Sz9�v�B�ty��PN�Co`�*=���N����,ڂX�I��>�U�0�z��'q�װ�����P��*�e�si��
��{̆f�³���W�;(�v�V���,�ʀ�+A��d+�Pnlխ�v�PZ���)J�dY�Ab�E�(��EUdX��*D��RkV�ITԨX�D�fKKj�.)�]IQԬm!��RV��
%E�K+QB�Z�!X����]j!p٭Rf+h-ij�m(�K���Z��J�Q\Y,H�g31��*V�ȵ!m�m�Ū"�cj�Jň�n�jk�v&-���ER��V�T�J��ѐkJ�Z�kE*��a��q�C0�6E��R�	U�T���Jȶ�хdɳ`Vm��նKFd6(�l����XT�l%J*��L����((�ڈUE�ԅ]`���˗d�A^t|���Ű�Qc�i��}7��g��#=�,���p��(T#�����X�G��-��n\����g-mFa��wu.���}�6��wu`�z��bQ�O��]��P�;{��J��J9K��x�ƴ�l��
F������|A?��!�lP�dj���Z��,�Kݧq�O/0v��74��z���,��_���Z�*��O����n5\�e�|Z��������	����#ዕ��Sw���c6�b��Nƾkۯ(x��yJSl
;4���$���{W4�[-R���k����817�s|�T~6�W��m/v�5^[� eײ���?#I?
�]Kվ�ۖ_d�ϙ��{�[�W6��x�}������Y�oW��m��YP���-~����o:�wO�n՗�S;l̉��{i���N���}���ͽ�3��+�Ѯ��Y���E���,��7=D/mS��-��pΜg����^��ͽ>�[]k�5�J��^�
���2��U�˖i��zS�Y�}������&�W6�ߞ;{�1V�@� ��vx��.�H���=�0_�����k�t���nn�
�<��`�x/T�_��x�A9_ �5t�^P���3l(s�en�|�ux�z�]?�Zp�X2�Wls�`�?['�%}��X�z�U�Ú�������=�������ם������7ܫN�7��;�}+݂�Q��}~��+4A������Q�F���C[j�!��|�~����B�����e����<�fme�c5kS�%	K��,(n��ڵP"�u��ĸ��VGyz���o�Ҭl+��d��J]M6�*$�Ȣ۶�HH�֍��ɷ�2�g�H��y*��ٙ��7�t=cwz��@���W$�����t���Rj�Ceiew,�)�U���~�)����(N�r-y���7��ƴ//'R����ʺʧ]��~�߳vĜ��T����[��)�v.w�~�c��)�k(��gf̈́�,�%�j���-a��c)w��s��ërOj���sՄZ��m������y���nM�ĽR���{�� ��p�l�X�h#P
h�>N�0�ϴ��I��mL2�&�����{K��J��}wkTG�J�w\��3�gR���S-���9�D�������Y�1���c�ރ#�V�W������>ˍ����v$����?�.�<����}Wh/㣒�T�����9��i�:*6��C���[�_w�o{�"'BU��U���1T�iݸ%���?��3[l-��T҆�����O�����ߣ���ō���{ݑ�^�kȼԋ2ܳ��0�7�k��^�~��������>5^���c��%ڷ~���-�2���o!/��6��]S��c�_�}S��`��{�噶���j�����g-%W��Cv5B��[cm�N�W����ep�I�mQ�inV��MYy�*uG��*|�PY>jA�^wL�J�ܫj��^8]���`�sޥؚl����N�Ͷ��3�؟u�(�ڶ�ʴ��Svmw3'�L1)���-�����ˤ�iBR�$��
���ܬ�r�^�o��KTX@�v׾;�4���o�y��s���[���/��[4�kޞ5Y-&qn4,�md�Z�v�����ڡD�׸��e�'2~G��86�;<e�z�$�ۉ����1�P]���m��Kj��,uȸ"�(K�2u�Tc���Û9�;N���u��a�7m��H�5��y��Ѫ4�V� i=�UK�V����åB��!Xq��J.��:Y*��c�7u�k�n��Y�iM�oWx�p�gU���%�5(���qď�1a��@�.��'�C:f��Q�]�b�o�U}Z�'9[�v�������|] *���Ƚ�!i�y�㏎E窔�ԟ��kw!Gp��7�_a��s3�J�ˎ�v�1��/��t8�Gl�2�a]�Na��ǈ׃�~s�05�5���[�jױ�9/K�����̹��ϟ^u0U,7)&Crq��j5^�j�uT.s7p�ok��er�g�/�C�6��	l؂����=-�/�Q#!�B+y����Je4;��]������ha���^a=lי�A��&NB ;6�G	���-�?��WE���d���'�
���	fJ�>N�me*Z�r����,�Y@_<�
apת@�GE�^�i~)S�Mm����fg~���n� �Y�˓�[������^׺d��2��1>jw�v�N-=��I�;�gDٻ�T�sr�{S��R�i黮岛���eod�k���ވ"��B��j�� ��9�x���gY�r�;l�c���H����"�l��d�%�2�:[)}:�Q׹�s�r���O���N�Yf�;��;��M�!#8�D5vBӐ�L��_�T9��E�_1����B�2�6}ѧ���s*���(�4.�\��4w�W���\��B#������*4V�Efb4��\���9��(�r�����ZAzL~ݝ�X�ŞZr�\�R	ۤ</-;t��ze��p�t��)7��׋�'����ox]]���J��q�����薶��r��_Q�PZw%�)l�;�����wW,О`#�SP����������"� ��fw<3s���������a>���杒ןVT2�}�|U��"�.�貳{��#s5�ui�)1�
4w�Tt�HH�c��f�qE	�Q��N��'��t�:�qmmT]�WL�sY��<y�	�H�*OT�-���<��(+���2{����
�#J�{2F�Ԥ*��:c��i��X��,��
}]T�%<s�5�Zs��G`�أ��d�u��C�0t���j��8�	�~'�6�ƙ5�7���������t5�U�T��x���.�����u�U?y�L�^c���nc�eY��B�6�t!����\�oiw�y,0��.�K)�u���'�5yGl�Ӥ
N�T2˨�1�*�x�e�=�0���/���/��Y&���"�PE,�����Hܧp���!��L��2}QsaY�����;�(y���*w1Ј��]�ej�uG9��K�'ݝ���"��w\Пv�;����Ό�f���؋/�W�
�_�?j��n��e^X+`SP$�@�ҭb�=�^��V����-��ܳQ�{���Ԯo��)�t�#����r��aHV���˿f;��-�n��O��!��E�><D�{sM*�v��t��M��J�d8h;�.�.�Ml��P�Voq��������b��4>�C@O����v6�,�چxn�������'t�2kq�L�Z�&�&�Z����ګ���m�ɖ�p/���d ���;
�QC%�*NWA�Ε�ݬ��R�s��a��jx�XJ��4y���ӽ�p5c��^tH��a�'�=,��P�w��v@��-:��뱳dv��p���b�o`;*[ME��;��4�b������-u}��{���2���(s6�lخW��_A�< >��/�����u<�Eq�6K��3�����OX+�g+]i���Ma�4�S:e?/8���Es�0;%l�\Y� �S�@��Ɖ֒����Z�5�k衳ϘZ��a����tt7Fx�s�%��H�2��~'m�Hk:Y��~��GJ�{5�pq��#�Y����u擁�=*��s�Z�e��1qz\��7w)�fm���f�����V���Cc�5��
�)��U1	�t[ys�0�q��^m������8�m�X���%T�f%q�b�M�p~���=����J_�[!�P�����&�M}�Wط,�*8�[�ޘɞw�.��/��p6�n��1ص2���b=w�۪��b7w����9�\��a��y�c�Kn��oQ�޹͇]%X�l���]�N�g�aR��#p��XR��t��U�?�UUP�k�WW��Wv���"vv\	؃�g���9q�GCMT�:����["<�sf�����r��r��5���:��wd ��.p:)�7��
�F��7��l����O�^Ry/rw���ډ~��<��s��mLO�-����T c� �"[�g�����[�Q���jc�q� ��Ulv���π�5Ɓ���3\(a����^\�1�l�n�%����6��m�~QT]v��[q��5g3'��½t�fZ��ǖl��^3�8	m�Nzo���83�n�M�w[�N����~�A��bx�_��o_����w�@�c���<�Mi-[7��_�:��	��+F?X�9�p�u��s��g_��V�r�&��k)��8���: N�g$�7hV�Vl�M'z��Zy�Z�ݷL�uÄ�z�7L�ԕ�<ӽ�j'�=�@g�����M�O9��T�W?o:�q�魦�<oY��H�4�.�}��.z���ѝE����gǜ+2��[����V	k6B)'�8��2�vYS�t[)��3�� Yd�k]:���ԍ�}ui�/��Y�i�dn���.���Bz΁3���~��������;˞ӔV⤄+�n"�Y}W�µ���oq�����wJ]~�H�j��`�_Z;O50Z���Y�Y9��Н3J�_+��)I7�e3+�O���{̚y����t'O��6�c7�VU+w�@~e�Yj_���:Ge��r2ͫcD��w9�^�t��.��SX�SF���0���?Z�����r���Ƞqd�R�K�?�Y8���2ڟ*��cs��ek�k�:*��d�����7��s���X���L�{���.19��Y�9��aK�j��b+�P��j~@��vQ0���ӑ�'��,R7>h�#'�(M�=�������q�;��^vĬ��g�9�Dq�s�9+���"%Ds�>؂�ny���dU)�0-��:ΐ�l��F�ٮ
�e��������,:`��%��{L3�F��g�=<���>�}��O?l���c�kװ�r>�J�:<���.;�*���"�2��jS=w���4�o�艖������}�o堧X�?�?�tmx�O��wD�b���⣟��(�U��Wh|�r��IG)�����C,���>����d �c����������-���欻�GX�rG���3��������2�!�WFKv�ޢ�[�S�-�0��TT=��j�v����X,:��C�`���e,�ޙ�p�y�A����vw\t+P`���X#�y�΂f�{��͹�F�ݳ��IL���1�!�uJ���$��+�o���=T�A���S��)�_��������r���K�xn���}�������n�"���p�ӽ�6[`�ȌֈPwp	囂j�p�~�
田ҷ�ų)~���w-���rtϕ���秠w��т|Z����-&��K��;��~ҩ��,���"=�a�1�Ϸf��-T^�ڴ"vP�/HͣIU핖i�7L��Q�`M;�3�wC{G[%E	n�Zn�B�,�G	�x+ו�6���[Z6%��c�9�`�~r�W��-l'��	���S�Md�>��q?Ȋ��k,�����u�OX����s�kr��(o���.Y�]0�����N�k��C&J�9�����l�<_j<S��l��4t��Lz�A�BF�F�L@�|Sb���t:�+�dĐaV\�Ǳ;g3�vG��2ԜqS]R@�P��<��[��YM$Z�ծ�P��|���Hh�3Ѷn���͙:[b2a�m?yN���b�9��R�ۯ��S�5G5kn?U�n��FI#�U�1��v�	���xF�ƙ<�y�_����:��}Je��4�>T��,*�zw��Z���J1��4�����Jt���=��Uԋ{�n�u.��>9NSy�\dEXN�� .��M��gmul'�������0OgS��^_cO��ݏ&�t�֯%+�K�����Os�d���Jb�N(�oE�jV�9W���෬8�|_i	�T$��ּ��:h�~�w�����և����|�k��ٵl�q�t�E�����Kd!b�D!>n5�@ٸzAx�]�i����Mj�8Ls��(Ӂ������r�:�(��U��0�U���\v!���k��W��<c�tN�ޣ������DX�`�$Omp��qVq�28e�E�����(qw�"�S���1�g��x�c��k�P�YsŢq�:��p?K��w+�s�m�й���t�����Y��L�SQ�7�Oٶ����I������a�\�7_>�mC\vT�-m��fn�4odo��^���p�ݬs{����7�v&�
�����jY�u�B ;^��IGa�ב}�Rp�b�v�|;no�D�l�y:t�GB�v��eZ��~jw�2���r�Ή��|Sg�u�8�iOqS�FRm̝}m{����3����=;M�-`+U-E��;��8J}�$Cޜ�����J:�%�5�?^c�4��KW^�
�r�]���
�v_@�4�a>��O@�����<��g".��^�d���5����w{��	Q��M9F�܍���� Y^٘,����f�.�ƿpܴ��߰|��Ѹ��!�UN� J�!�376v�P�s>��aj�6�p[�Su+r(-�wl�53,tQ�@ ��7Zx�A����B	p�����8�����m�3�Qlh�bMC�����99\�{GYP��1�H�B��
�f��q��*_�]���$i�dI��2����D�mQjX1mJu:`4P�v��f_W'�Nɰ	}�
直�]j��u�r�5�W�$�3��wh|gכV݇����h37(�
4�a�J�h7R���Z*u�u��ǣ$�:|7n<c|�1MR%0�{����T�C{+*�]EgsմW>T+�5k�]��RD�Z\��C%v�=��&VS�Rm��s����`�f�N>��l�"&4/���zS��78#�]���o����OR�˫1Z���Z� ֕��k*iZ!�-눂�*�|�*���h&�x��ȉ=�ޕ7����ۼ#�Ȉ~.qs����4o�"�	GW/�ǲ�\{^��]�T�h�0��D��qC�-������:�\�b�o(۬�.���T5c5r><�5�'1��HS.�w��䒳��(ɜ�d�j��a�_m�=�!rfv[eT��5ڱݛ�/��FV�D�p�qu��9�0�9���x��ۧ�]>'6��^��n��t�랻���+=n����d���+v�a=�X����<}�mDжr��Ԉ4���-�V��Ɂ�"o�k������9*̶�{�/Y�n�ď$�]>�>!�;��e��ث���Z�U�E����s��In�iɠ+SEe�1���t�Ͳ$�g(�2�}�s�RR&�?/���V�=7��]\�sc�{�f��~���H	+�2��TI�M.+&��'	��Xt��Z���c�����;UE�6�	���ޫ�@�jX�C{q,T*O�`�;�*)u���A�{Wp�9h(�}�@�oM]q�~>�ej}�3����ܱ�;9�u�����Il�;+ƒ/Sv�������pPN��a[��;o�>h�w޽Ҽ�5��-j��;4 ��]"����r�gn��S�I�0a���VL=��ȴuR2�w\�T�3���H11gqN�[kr4�u�J�sGv��q�.��CI_[7g��i���$5�D\��bT	<�)�{fفry�ZW��5��nQy�t���V�U�0jyD��\��'�'W��(�Ÿ�	ב㾓_b�k3�1v��QuS�"��.�&�}���v�ӭ�R��,���$�Vz��
�8������k۹x�(% ����/�0�կ���}�w��{o�a��r�{f°����)�2�k����	�˶i�.P`;:;VuJ�cv%��>�e�6��������|ʺe#���{v�;>�P���4��Et'd�W"�vN�;so��b܊56����s���82��A�ŀ�!W�t�y�VTj����,�՝7�9OqeȆ\��Q|���(T�F �"�k���Ny��h��\)�Y]��B�����}{ےԽ�qnl�mg�|j~���+B�5�!6�(����݊��f�k�E���m�j��*��j)iKR�(
(�۰]�AA�`b�T�MM�*��
��TdUVҲ�A������f�l���̍�D2U��*VVa
�V,�m�����*4m�u�(��-�)Ur+R*�ҵ+U����v� ��1�6�T�Z�]�ȣu����XVTXR�h�]r����Kn�DrlUh�k3��Eik
�PUX�hT���b�q����;Tu�؋�QF[E+2��F�T+0�k��B��m�B���SZQ���0f�*�����dɒ9)���k�j�[�6�U\��Ъ�m
��[����t�>�￨4u���iL��v���z����)�0��Y��*�a�39}t�0����۳KHݽP����m���6lf�܅��Ӌ=�����'B,R4y@ԫ�ͼc[{��P]��4(ʄ|��������	���ךNCOJ�q��a��v��$+�Cnfk�+��e�Y�v~*�`X�}��]i���vc�C�ߑlħ�Jz��YE^s��֗�by�,K���u��Pv�f�WOF�J�wL��x[m�i�&	�~i=�!�����8����ܪ@�iS��k�Gx��d�檩w0�U��LJ�7�#cf9�]L#s�Te��k�r盫�F����`� އ�/m���9���������(3(�~�1O�3�ŋ��N!M�,��QAG@�ZI�je��2؎L�Tߤ;���c��M��Ǫ{���5�8L��o��-vs�e���3��p�dt�	��P��?<�lHɦ���c �ܳ�.�"]�\��ϲ��W�f�4�\�Mf�j���s#�/n%'���N{������~�7��p���ôӕ���JC�X��O�(�톱�/�򦷈/�v����������x�nç�.�hjc:+�F	����.��|��M5i79�L{��KAs���1͹t�T�XIQl���4C���yf����x��v�mbΚ#2�4Qk�7:��Ж�]���)��J_�B���z��vk
U!`��8��-^��x���^�ɒ^-�py\��NJ��b�D��.�<a6@��<�͑Tw��{�̓_��E�,��`J�����<��DF{�y�������>Կ�ܮh]ل\�e�3��`\Mg�ڣQz��\e���P��:f���T�,X;M�6z��g�w����T���]q��ؾz��qqۊ [i�O�T��YD��{�G���!e�Eukcb��f�P뺛�Wv/�H�yGE�V�BS(P���l�;g_vO��:-��GI�x�5,��I��3��>`�s��6OGY}R���#���9m[1�{}�wOKpL]��<���=���%�˦�a�s^Y;��ѳľ*�%�]iy�ථ0�7�a�c�,re�p��kEF��}c�D�JnlSc�S�NV�۸	c�~9��d�ҵ@v=Ok߆ѓk�Rs�{2%�CT�5��N_1���O�Ot��MuI�ӑ{�x�,����=�m=�b���5G5�Yݟ�`�����&ZJ��l�O��z��2f��9����t�١t�Dc���y��ѐFf'�q�>S+�l=�m����1����6'�9L
����뵞q��O0�a� G�Ls�5��[�,���x�~!����F�{ɻ�kN�Kw+B��L&F�[}�9��ړ�|3�� "���[Ә��e�;$ՙH� �M�������hF,EJ�gH�\��Z�Hk�ǩVf�Y2�uln���� ���=�����$�w�e�'�%�d��#����l�ׂP����y��y��+F7�Cޝ�	��y�n�{{�esOe��u�q>��8C6��$�?9��{/�2v;K|�y��n�G��<z�l��{���	�톿0���kʩ��0���d ��:8Lyo?�_%W�3rM��i̶gD#L���kȎ×�{
��FC����n�/OA\�;]��ݤ�ʗ��3�KX?4���t�d��#M�Qb'ݖ'�#0�@z�Dڸ�1k^S�6|����-�g˶���_�<��{x�����6V�{���ە�#L�l���ON���0�zb�ŵg^f�X7��N��i�t�$+̎#V�>S��0�^�#�t|gLe�n�������S�"�D��C֞z������(onD���'���Zr�B���4��F;+����@�'�]f��~g:�xmal��r�K�3N�-9��b����O�x&�����{�T�Y����?OO
׸(��R}nw@,z�xqT������׊֭g7�z�FtCC��1�D�C��۰�M����u.�l9��؆M�/�v�󐫸��7*f�j$����z�i�mOg(�y��{@���S��Us�p%x��CVX�d:
.�mm�ÈL1z��Ń�)�வ��{�hѫ�z���v�m�jj���;����{�ҥ
�ꎂ��܄���\v��Y�'	�������-Z{�Nz�D����᥽�8���7�tϩ8⥫�H�U��#��ӕک�*�~��֬�?��>�a�#;�W6(��5��ُ����5�|S�ǔ�pMu-Q�O�
UZ��W��b��,�e�;:��rE�j�se�?��B�ձ���a�8�s���i�_t����:�#6Ꚉ�`M^`q�c�C_]��q�uKۚ
�E�6�t!�y����ηeQ{�������x��h��ڧ��)��e���:�P�=u�ʲ^.qR���Ϋ�܋�����m�j�:�(�`���#��:�*��F<r��aw��x�6zޢ�GE
{\�o
|p�Qw�{C�u� ����t�qVt?��E��9/�r�7@}=</&��o���sV�SJZ�i�2�5��(j�T�Y��y�K6�%�^�vW=�F�Kr������ɹ��4�C�Y���/Ɗ�n�"�����z��L�_8��u�6B ;j�������(���u�s�iP��{�?(6�%d?-	�_ⲝ�j�'N���9�7���)}�B�jD��?qU|��m0��9�e��p���ī�����Ū�.����.\��Csk�p^�T#�L�]���0�r�8.�b�Ϋ�ʉÊ¼G�y�ug\�"�S�{�/����M7��L	jw�3��T�8B�:$G�V�;C}~�[�����T��#��z�w�C�b�%���4��<5��]4KQ}Fi߆��t���*6$�d�̮�������8OElئθ(�_A���c�l��<��KSΧ��˙���`_h�{�gZ�Z��nٌU�h.;f{��讘����r��`�f`\ͭ$4<�H��AUV�u�Y��{^QA���f��mk܅��iŘ��ڎ��x�t��i�[m
���"�^4v�
@VvL����u��z4=Gv�0)w�8$�Fz�#����pK<M�s�":�݆��ړF�Y��[�^�,P먇-��hW�˭7lP���(<�1�s8���e�C�W]5���
�]�T�D�#,5�h�3��Xv�i�t�@\j������M��:�+�|穽���S�t�1�9���v��]B\	mp��q���w!�癹w1�Y�6�'��1�t�#1�2�4�����8�Y��e�6�s���xJI������?WX�_�q0��yk�we�`�cwZ��[H�F��<��7jUä{�P}[���{}1]��r��}��8^��R#'���N^!R���!c~���}X�4N��N��ED�us�-�s�K��`N�ʊ��Ҡ�w-�9����gsS�������?.�g�F��Q�睡s9�"8w
p�="���Ѻ����_s�ɭ吖��g���U[��3�����:[��k�!\s��w<Y��+���5���B�.e��=P{a��粽�X�i�����5J��8�'��8�Ny��������P��%�T��f��@z� ϶�
�a�*kx����r8q� ���L=�B����zɓ���%�W(�pe�,F	J����u�	j�)�Y�����a���Y̚Q�٦�!�E?!Ԡ��(��?F[�)�M�b4WS�KWD��U�E���;��E���pɞs-۶����M��)l�{S��\eD��u����D#,�����uv�9Q��g6@�
s�н���.6ȟS���4��^ǐ�:-�(�4�A�,�a�n;�לʹ#}c��Nމ{�� ,�3`N:���/�N�۷�Ȭ8+OY�kP���Z)�2�5�Z���5����k�ϡC)any<����eF�ϊ�	�K�/4��Td��H�Eʲ���s2��.я�AK
�v<�kw;����[��뫩�~&������`wb+�H����nQD�ʶ^iO�ws�r�Aǜ ۷�6���i�d�W���ơ���)���"{��P���0��i�#C,�9[@3�{��A�&#y� ���YX[$���k��j��;����P���jf�'��p5c�t��gκ�D�׸��\vƠ�'�{a�ԦD�*d�]�g�{���Λ9@5uIҢ�>m�<P��Q�h�"�(M2���]֐��8��ں)br�2Y����+�s>u��uI��ȶ؂�ny���_47l�Ea���	�|��09�_��0<*+dK!�]��?<��t��S����Ң\F�|�=��m�uQ�w�B��.��z�ѱ�o·^	B\t4.q���ׁ��Ɔ��Å�؈�oZ,O0'������[m�^���z���3|�����f8NlADz��K�Q�g��K�ζ1����ݹ������p^�k�<Kk�5�ÿZC������SO�o�R@��z&p��dptgݕu<��+0�n��m���&ںr�����2���8�E*��ec�q���k�!�!�S�q���^]��iS��g��ݖ�*����t9�Nͪ��c�����|�����lR����)~����r�M�rtʷ�W����:2^��#�ڴ���J�O42&�dUMS�jI	9����v�?}��5}��e�gP`5�����{t���F�`3ڔb�8X�O�7�{�܄�m�r%�7g)�*ĲY������9b�l�4zg
�3��7(ݫ]`�L6���x��ǿW���Ѵ\O���ϩߴ��p�[#���j�A��8�Me2{��#��췽��ɩ�x�k�n�F����3�B�V`M;�3N�oc�H�0'��ԩ_f���͕{jC��+�jth��z[)p�FT:e6ĵ�����8���M���ϭ�Ն"_����|Z�{;a��gO룄�^*]`�O�����f|[L&�W;��[y�X����z���G��1���P˹�N�Xy�43�ҥ�g��*C�~�?<��~;��Q�O�Un�6�����귓�3��t=�&�e���N���!s)Ό�����s_JA�ț��5vq�uQ����rB��)���7`�љ:Y��]�<q�'�
k�X�h��v��{�ម�t���h֠z"﵅�g�.���#��dlߏ�E	���xCm�iF󜬒ל�D(Y�x;[Zc���T�N�/Y�Lyߦ[{q�	n�ȷ0�U��l�,G�����'gv/��k�㧼���|� w��ގ�����&�.�z�9�5�d�_U��O*�'�����ڨ��]��H�}��[/�h֭�Zb.@ѻ��5��3�~u.���x��"�}���ZsX�9�0=���͕{��$Xk�#�˸��hy�wԬ)����;nv�6�}s� �X>�_L�Θ�]�5YT"�td��6i�������3.p�C������ ��]��4��2j.l$�l���w�iѺ������}aw�Y�#��[K� K2·�>�������/Ϗb��>���9���Y߉�-w2u�n��C;̢/U��-���-� �
XCc�s��ܙY�}.���yF�mC`a�3������
�sF�d��W��]�I���Z�#��! �Lpy��`��	��ݠb8n���:�[D?+O��
�_�����lU�h!���v�S���T��!s����>dj��/h	z���]����Lܦ�T�3���A�薰!Z�h�/��S��g+ct�Y��tf�8[���"-�w�tП#�v�B5Elج낎��
|��^��U,�Й�֨hȩ���e������v�-�v��\w7s�u=<+^ࣔ� �'�p��bf;�c0��&t�������Py<�/U��0�1��XmE�����Px�4-Ɩ����S�8(s�G��q\ϐ�Ц2�C�S�;>��
]�	���ז��t�v��[$?=]9t��7��[��AeJ,N�"r��ݹ+ۮY�Ⱥi�N��Xn�(qn�T��'8M��mf�;��W��5�,�e��5i��1u��`Ś�cBg��t��o�ĕڞv��Q�5����Z��	��ǃ��(���LM����{5�$�fέY|�Ù�pCl��:FZݟ�k��bY��hSu��f젶2:��[F��F!�,���e��̲�_�+���n���	΃��H���i]=%q�b�H~hT�K�j�r����/K���8���L �T����/#x��AUR�m��7c�xH�m�cy����G+7G��5����^� �e�: �P2��/����#�M�<O2ƌP��U-в�xv�vT��y�s���#�PU Cw�â��Xߨ�a��zj���k���-��c��a�qS�lr����s�/~��M�K=\���2/�c6_s�c@�����3�r�Y��;���l5���_}Mf�_��̙�٨��/�VC#Zlu]���g�����n>Nk�j��V�PJ��~qF�FK=���W/�q�8�� ]���	�S!�}v�Y��8l�������fא�Ϲn	�J���C
{�B�\�4KS��n���>X�f��E�Y��t.y@�Ϩ����y��N��v��]P�$U����`��Y[o�?�6��#���18�<=�a͕Sm�'\߷������JucH��:�zZ���P��k��^�{��HrՏ=����D�G��|
��,L�8��m��7M'2F,�â��֖�m��+Kǜ���{i�0U��T�f�dA����f�to�a�.0Ԕ8���|9�1�e����JZD w:�3K�M���NS�cKΪ��ޣ��Y��F`b;}�q��6@�.���)��&P:�q����\�皷k�q�
�Aؙ7ϹR�^#2��,�:v�mAr��5��z�\ ]tp,sh�[�۽F
3GVsB'!8,�7��H���]��`�%W
��d��좭����,�o���q�Ӫ'2��D��[�������\�$��0z�ޝ<���=�qi:�>���ؙ�e]�/�����N��)qxx%��F����']	�#F^����(�NAQ�]mq���oMo=� ���X�&��?2D�D�^������Q�ٲe�=�*}���2�Z�u�wu������N߹2xX!_8z����&E��x�}�u[!�;��T��1�=���-d��Uk�f�]Y`�<7�l�?pǆ�n���s[���J�%��u,�6	�r,;���^;�X�9%�I;����k��νgE+O�@�G���m�V�*"�^���zW��"��9���^��ED8��&1�>x�]2�'���f⮧�������U��Ţ)��E,��t��:ʿQ��ղ.Ϛ
��P��i�.�tCy�@o'"�R'G\�i[&@��\dp��,e�U�qa��;l�Y��r�n�2�{�����`ֲҏ%G>�Cͱ�g]-�q�*��9eV�'�.�t�)�,mJ��SSB�m:T�
Yf�)B�Z8h�T�<�y�Z�V2l���Ť3n@�ty8�G���k]���g�U���Y��ה�yi�dk�W�¡��mP'//f��Ut�y�I$�F���B�뷙�M��yw/1K{��+1�)�������9��Fz$lo����v {�&��\8��N����J�EZ���^
��aыsku�	�V6+�g�v�v8��{6r���I�)Co��ne�*j�Y�kaH��6�h��SF��/�� ם^���w�8=�&�u�q�^�sx\t�}��H��Y��ݷ[Es�)i��c;�k6����F�|@�(z�B�'�Ko����B�7��6o�P�Xe`�(��հ�@;������j�G��w�㭰��F(6�'bJ]���1ޮ�9@��H$B�L��1���j�ª7׻w5mf�8:�F���x͙��@��T�	�Ǌ���yJuQ���Ћ·�~u-֌��Ni`����ӕ�'֕e��w�݅o��:a��E�[1���s�=Ɗ�b�3����Ņ��fo]b��dmp���dx`������kyy�F�Κ��t:���>�H�JU�Ak�iF�V�RڬXVmbŖ��E+S6�e��]���SQ�L�n�(%ne�kdQ5DDE&J�R���4�[-Cjq�W
$�-�Bԩ72�k(�����6d�vʠ��A5�u�uɚ�\т����-�lDs���mnmjPiU,F �*U��i���C+Uu�Ṭ-�*�*.��k*V�c[\�d�mKJ,�U�TEX��*�U%J[mP��hUDT�*�T�TQkV2
�B�&�PAUQ�,"$F*�T���ư�F(��T�3��kJ���b)U�Q[J%h�Es��(�V���W4��E#R����R*��UT�h�dր��EEU�L��Q��"�[[J�@����g�;5�*��!N�a�{��~�.����AS;��3$w���B�^˦��Y��՚�Yf�a�����_X%\���K��S�!-l��ڟ`ו(g���Wl9w�Di�Zܑ���t��gX�湔OF�O:P��u��BS�����,�N����E��̓г��n��}ihj�y-���y:�lE�8�jt��S��gڶ4Kb~Ә�_:ڎ��k)�6�VfZ��3�M\T��;�x$w�!0�w"������/'��Q�P|Ʃ͝5���9"��G;Q��}�����P������nRy�������\�u� !k�u��0˿sC]ff��Mk���wc�`�R5�$iP�z0��nZ*�#7����T����ѹZ�Uz�]�R5F��0�����I\S��6{�H�Q�N���l[�-#y5i�`�y!vC�iz�h�h�#*�*�у(*=�!�}v�7�9�ݎ�CKMBT���\���u�Y�#ݳB���oC�6:-�V�^	B=�:8�q*�|Q�u=ק*�γ݀y�نl�9�q��M2�t�oe�]Ga�����#fc�t5w!�@�d-^_�PSg�WM_
r�&�[�(T�I*+2��hZ��
��;źú�v;�VJ	��ٖ������"X컙9�S�h����z�=�1�8�B`�ϥf�(��}E���4�J�I`��gV���O�~�\D�}.i��ω4�Y��	Σ����ك�~�&��������7>��n�oU���,Ϭ�8��Q֝֬�nwǁ:/lQ�5� 枞� �"���ʋ��O"�Y��t�Fٟ(�qR�Ӕݱ�w�����-�[��q�|��:��z }�"R��{���O�.N�pp�t�{9���s#f᏿^/��ۜ�;�{\��Z{�ik��}��\�)aZ�y�d���w,��nN���E^����of2�=D͔������Qq-N�����J�c�Y-��F�tC�+�U��M-���e?h��~i���s_�e�=iOL�3`C*�fӾ�-N�oVD��䨠�u�a#�ɾYq����\vY�n�Ў��d�lL�'�t���-L"{�@���e���2��s�E9��Dԅ֪{E�u��?ʾ�0K?OO
׸(��R}�;�gh�By�س�����O˝�:�ݶ�e�'�˖UϺa�:��o�=�ꞔ(�=,)�Zfݝ#��Ud����ܒ��5{����zɱT��Z���M�6�=��ð�2����$D���D�������
��FS��������K��3����s�������8��K�n�xp�4�Gۻ�d|��d<���z�4�Z���Ս�/����;� ��4.�wK�����y��-��Ի���f�(kث�mVr�*��`��g�����oE��6(W���6�q�l��ӱ0�,�xd�8܀q��9��2z��ʔ���uf�$lb��Nσ��.H�T�b���̦�i�x^�Ɨ̊Q1�&ݗkoFm�9�._�:e�U0��0���.��<�g�0W�q�W�?oM��my9����r���{�+r�kP�bs7� u>�q�g���'�:?t�s����2�.�3]G9���lI�X���]�n��_�0��B}�w<a_@�[��:���=�a��(V�Ddp�u�8�5=K$:qcY�ͧ���QfΎ.�e ���n���뎎�L�#Ͻ�!�z� �틡ѳ�\�Tj�sGnӇ��b�׮"𪷡m\�ͅ����?W;	��,�nچ�e�8	[ZC�Q2�o:�*z�(�6u�Xi�ѽ�e2Eu�a�o�fӁjru�B ;j����7i����0�����5�L��J����;D�}�uݢJej�ӽ�W8��!g������lgxё=:�wj��s��|�1�z��P�M�b4m7dN��Gq�%�V��&��4㳩�[��Z���E�j�zȈ�4��d�~�
\UuW~w Պ?+���>����]U椯N�b,`fhor)�k���5A�p#=�	�gV
�oj�\߹̾>:�b�)���2�t�]۶�9AL�i5ή�l�M��)��<j�Z�=��-�޻�H����n�~8�Do>��r��[6"����lΒ%Q}[��6�Z�Y��՜Ӌi9�9�ai��㻞�%�)lS�g�W�]��J���n�,����O92�D��ۙ&�J����Fsd�=�@[5<���N���S�Y��[37ei�l9f�����%�Klf�V�;k����ͺRk�l�	�<�Gd`R����>y9}E�[}��Q�]��1mM\�EK8�[�*����Vu�*d�?g�̫@��v=��HPU�^n+|r+�Wb<�^�]�x^������<��:�E�k��WOF����gZ˛1��&�n��K��4a����.�3������ �J� k�Go�^Fq�h�#�v�]P�W�/�TU^t=�h�<OQ��졳��� ogހ:X)�7���l����Q����/pmnU�V"�3'U�ax�VK���Cle�����:�@�t3��ӗ<��L���������3�����W6>�����s�/�@>GKp�q�A����/�=�tB�5�����ي�X"�(��~ԧ�c}G�솕%J��{�qW�����J!�*\�Î���]-��P�#�9	˭�8�Kv�#�эs�$-������Dq:����+�Y��eu����vԳâ����ws���LmL�;܅G3g]Pd���8�Λ���n�/XPۧ�2֟�<� n%5�& m�p��c7V��q��2�Nzm�m�������ag��ma�~0י������tVxl.}�Ǟz� ?zT ��:^R�¹<����#�pp�{�,Yׯt�
�)�,rx�%�����lc���J�u����q��g@ժ5���h�2�S�9��%I�Ń��R��X��)�os6���&Y����5�	Ntȍ=��
����k�<s;jP��z�\l�u��R��qG��Q����63OB�'��	f�u��BRђ�	I��,���e��<+�h�l7yt��t�y3��2g�0�`�"���V@���/4����j�ѧp�8��Ѳ.�/�^ *VY��sr���^;EK*�)<�;���ف`��R�K�?��#�����q�[:�iU��٠t�<�+�����qL�ц��k� %o-��6Y�m�wC���6b�H�ݱ]��q��mFs�3�r#���@6T����br��kv}G�t0�/�pcx���l����M�B��[de�VV+�L�+w[�����2�~=e{�_Pc
�P �N�>l�wj���
v�M���*�[#5�z���⥖��UN
��QU��P�ޚY.�`�O��p�����&޻��{}G�|'�d�UxF����vCt��i�n��5� )f�L�#�%=��)��-�56֎Q�ǉ�����c̩�0)�x
��*l~�vF��_�r� M��8a�j�?Y��i����#I=�t˼E��h��=MoCŧ��-����(Sk����Y�9��6�;�cW�)��.$%l��L8]�^�a����vYU�vG|�C��w��kփ=�Q�;{8�G�s�G��9ʞ�|i���-�F<{���a��*����ku�/�o��v�-ڞ�:r'xS�9���3tt!����?�쨸+��_wc���w��g�2SO��nw;��C�k�3��S^�4�TE�s�aL.5@�8�J8b4ݵ"}�rp�+�3ˋ�����[���:B��֞��K?*��C<��W㒷΂�柝�I�����S��*>F��gc�jǮ0z����DP�W
�	�{F��+}��f?��zu�ö�;y��t�m��Ƶv�Y���tN�_*���m�g��OM�62�V`K5;�4Jۑ�v���xf9�kf�~�;Ř�o*k�I�?�y�K�<j�����{�CA�x�����Y/b�: �x�o�X&����r+K�#���D��6�⸠`U����w.����r�P4: �l�����цSM�hãM�B#�혲��[w��}�D��"�$Y����α�周���������[_��]ϙӠVĵ0�Ou��/��}�ERM8�6pNg9[��oP�1r�g2}���ez���>~��[S�nRy�}c����U��������4��`�&3��nZ��VT2���3ea�j���OJ�(�GAT-�H�i&1O��V�>�`etw�b�?tتx�yju�=7p�-ѓ�i�v�%8��U$}�0�ҁ|P�a�Л�sc��|Fm��vW�!�~�0X��<�`>�n���c�A8�MƱd�����<�&��b�c�9>D	�/�e~T�~ۧ����2�˰�&ڶ8��v_2V�O5�V�S��*M[ۧ�� :yfҀ�]T�J�0���ܧ�7[���j5�]�E�a���U&j�+_��r��І�ss��-�;�x��{{��ϙL;,��uػ�Y	<}��9�8��(��=g�����;�Sf�3����r����bD7mp��qVz��7�D����i��9mJu�g����.lu[�[Ϭ�%�z����K� K5����E���y�vr~w�*V+{���P��)i+�o��B"6�k�Ġ�4x��پק�.���$w��KDU��t���:-�����s��:��3���߄���̬�+N���VgBĎ�S���w�T|��č�_�5ܦ�G�
����gjG[�����>�]�UzT�<8���H�>@�ߞ��o4��VY�3�p��r����a{{)s��w�{|.bk&�ɵ���4�6���Ԭ>Y�(sGv�L�]oxU�H�Id8뜄 ��0���U�W�ך��'J���n��^{���i�f7?=��a��ej�ӽ� j�����d�ٴ�:�����"��Pz��<�\��$]p#�̄vz%�j��9v�RA�ѷ��$�Զ��޷{�c�
qD��}Gr�*P�-�[6+����"�x@,}e�i�w&��o2oi� ;/n�K5<�<�tW�K�X�d�^:��k�gގ�S��s�3��IL8�7>@��*�x
1���:Ge��(͌��{��׭8�w���^������&Tfz�|;f�A�puk�mĺ��-q��,�����6������^���T��m��_+���W���)�v��LX��Z�``�?u�
2�M݇C��?n:��ȥ�/��͎gN��{'ܧ�S]T�D�FXN�O+�j��VK��0~�����3��w2��i6B
��T����i�&��ovOX=g�]_ s�{-�qdD��6��豠�z�:��{�D�o+�����l����d��.�*��o9��^��>K��������TwYO5�N�
1�})�b���Z;���Wu���F�6�4�O�<����L�C��#���D��<�c��tnjb��E�n�i��ݗs啄��-΃y��2Ͻ t�0oLt[�2��S�[�����49�������oX^�.�eq���]�;B�s�k��,;c� ����޾ͥ/M�A�"Y�&�G)�8d�D]��#�9���\ #��N�P�0��z�u<pF�C�cw���0��ON���ܩ�ܶ���-��M��׿by�����>���5J�����xզ�Ԕ�Q7eF���ny�=߻U��y��V~�A�&��~0ו5�@��=��Y�u�V����?c��`�y��v��Tn��Y+��+���<���DfC��v�%��VL~ʬ͡u���a�w�^s�z�QyS-��U��֝j�	d���xek��?R6��l��0|���j����|�,��ڞ��*o:hH�O�e�>�؝�����Ě��m�sN�֓����݂#��tT �b(�TD��u���������l��Q���m'J>)�5�[�l��T�wN�тE]����f?d4�r/��.Ҧj̟�gé�wK�kVk!x�Z�)&VX���A�7�W)kRX��V�(c7��2�I� �׃
���n�fiyY��BT�k�����D9e�ҟ*ks�Ž���yQ7�î�e2�&|�� ��f����d	�}���������5��`\���]m��/��3�
�Ѿf��t�2�(�Sr��;��0,S [T���n:�8&%	�s��vN����3;ا�	~|�>��9_@2zT����*�#�)�$�U��&3r�Vx�?����ں�գ��Oqn܌]�%팞�>l��vB�C�p��9�x�����l`wPڱ�v�N�FAi�ô̜�*�v;v=�i�W�Y�@�0Ff�+^� �?eQ�Xu�5���w� �Ҍ>�yd5R����7�
���X��c��t�-/H����շ�X�K�j ��� G�XIwЪ�0�y��c�kOc�[#�ǵ��&e,mm���r��3k����8����wS0U,7)&G�8�|����kx�,��;xK߾����G��;h��9+O>�M�S1�[z �%���O��dd�fT�rDϓ֛��n���r������Gh㍊�:��6�ӏ,� v���>�z�'r~3�Qp{��_*0�n��m���om׽����ް,�O�>��@k��p��䃟"�)��U��ok�sM��L�0{���ް3vj��zf����g��\LEb���c�dg��XN�&���η��c3����m��N�w�ս��8����=�T~�����y'�#�
Ĺuh|����	g��t2^0���n�:�>(��^4	�/�Y���,�5�:����@۝��%�{��"��ٳS��'@a	��}����hGC��lr�gv��\���ɕ�@�]���b5�{�+z�:�G��eάLVht�=�M
��0��{SbЭ����X��]Ց�����Qe��Lښ�v�Fl{qH)��D��T����VG�b1���T�����[��yz��1��и,awz(�jQ��,�����P,���&�Gܮ��]�9e��c:)0�2�Zv8^wk	�������p^����̧7VE����GE���z�=�7�ݐ�ZN��dE`|���:"#���
���
!;����U�#v�6����Wh�}�U�� s�f�9��ZMi�Σ��q��Ge�Y'wp�J�-��ݑu
��;�^� ^.��N��9f�>�����=c��L���mfZQ%aX܌�Ay�Op9��+�m��:r���'�4�aֻ�ۀ��ཹa���Q����4��}ר�/
�-]B�6�R�C\Y�_��aJ~8���v]�\=z�Õ���hk'�>^�Φ��.�nm�=�p|�L����^�����7�H�H�O�e���`+���>xs���X��	a�auA�tH�"C�էq�^ �.��AS<&S�z���%S1bgC�jʗ�O7�$���1�ضo�y��Q���#��ނn��[x���q
��C��ס@-sM��.��DEM�����g��d�S�yoQ��N��ٯ��$�aMkP3���R�`.*�;� dCg���x�q~��ЏrX@���ӷP�� geԏn�L��ª#���:"��]|OU�ֻ	Y�r�yPx����������[� �mܶwf����񪕻M�ݎK)�˘/&`�[���!�u�f6f��_ub�v^�{�v�P]2����_f����kZ�cqk�F��n�����o���j���cF!���؈�I͵1X�ל���呩�VJ�XF�6��Y# #��&�\�fE9B�Q��=3˴�u�]΂ggq�"[{��7��
�My{�N������H6U'���y��)e��&��{d�g���BR�=�p��%Aw�|٣IY�E�>�~ő��s�$|^Z���m�`��4���V�S�d�]�������;��=>o�>1���Db ~-b"݌*���D�e�mX"�QQQ���,UU�� ��b"�TX���R�#T"�+env)��*%���3
������4J�U����0b��U�R���k"�V�J���UYTU��m�ZZ�
��R� �b��T�(�*-eV)m(��U"���v�Q�
)�ŋl�T��Z�V*��V��-�#Yb �u�,Qik]ak�j0b1ZX���Z"	��reF1����[F#"��j�(�TYu�&j"[,TB�c5�+U�ʡU[#l*�-��EAQ� ��j"�UF"��X�Q`���b[Q�A��F���TTX�F������**)��Z��b*[*�ԕE"�5R�`֌bE��j�5����U)�V�u�-*���E-�dEb"(�0UEE��cR�Tj�*���/ �����&:��w">�j>��M�M3��^�����5�qК鹔�R���O�sRX Sf/�K�x�}Bt�{�7�.w��:c�[�%��� vm���)(�k%й]�GK��A�4��鈆tD�[�,���[S��)=�:��K���w�_�<��v7e��M��طzMw�F��=�q`�t�
�Q�D�8�N��a!]�Z�w���e�C<�-nδf�����V�e-���Z�	�4�e��Z�V`KS��,���c�8���7����<��"=]��r�z��8i���y��:�6ĵ0������5�lk*��9��!���6;��4�/�Kb��-��nS_J%�zxW����V���=������t����֛�n���2�M<�w�S�Z�YP�[z7L������{С���*f�Fy��#��Z�[�	ȡ�<nv}ӝ⭟ت`e4���ՙ����i�'L�'WMQ|9��91=W�@�z&�C脍8�T���$Y�f�;1�v3�ƻOw�]��錣�gM]�ڗ.y����R����O� Na{�������!߲6f��̠�Vǒϫ�4��~�5s�gJ�!�
�پk|��ݲ�{F��c6���C���#�vb����H��Vr�?Zb5�+5�.�Ϧ.���9���Цֻ�7\h�9a.d��<��n�8�osF��휸����6�YՓy���͏��B;�Er)ţg��ܞ8���Y��ݴ�CJ�3@��j_�����zM~u5�#�g�,f�EpL��o.fV��Vn9�4X���7�sL��ޝx��h��#zz`<��<vY��ηWRwmr�jf�#v��q�����VKӷq�l�!>�s�8�wd��O=ۆ<;Mp�1#�_-o^Κ��苎W6[�[�Y���&�:[���@W��q��"�>�s����R9}F�5��֪���Eb��Wxz��E�DW>a@>zy�T���9N��p�<�g����J��%eѢҕ������n�.�=0~�T�B������,e� �g�����^dJ��7j�A�?YS�-vԝ-�J�,4��d�{�Xя+U0(�����KLu���ά��n��hp}���r���T�Y�޹C`�v����dO*��熠-�E�o`T��o�����~h���FZ��Ʊ�-����9Z�Mj�,ϻ%�:ࢩ�����T�c\�܋��=�p��x���ۦ�O:�h�K� �[�v���l�w?a�S����|&���\v] ?k~\owk(�o�]�Fr���F/U��-�\%o*T��vMcv���@҂�D{A�C�m�f��_h�חo�d"��Y�:!����ٺ5���U�}a�	�	�|�yȼ}-<zxL
o��w�i��FwoWJ[��	x�v�s�m2�Y���O�`��)� ���0._��O:x=���P�(�,-\u���Vt�Oz�x�ג�_<�n[)�>�BMZe�� ���`Y�Td[1�i��|	^n=sj��nnh{͢��;��׮ tt)g�������+:�'m٬���h���?;b�ڮ�P�kpU��^�%�dt�`�3��T�2���i����H���o�ٓ�:�)�ٚ�Og�Znز�l���Cm�i�)�'�; �n�"T���j�h!$��Duv�5�:"�6Ο]�;���{��le�`�^� �e����ֶTXH�3����^�s���b��E~�Q�*�KM�B����z��P��l�P�p�]�;C.g<t�7yF��*/˿j0�C��w�gy�T�C����#����k��=V�>�-���\ 1������]�Z�Yu[�:j��9���'�灑,�d4{��hX�?����pz�Y����q䵳��jeԧ��T�ixD��?9��NyS�[4b����Q���]R�a���o�¿=uh�E�Ň>Dg�\.�D�_�@�Y�u��;����:�ǟ���o6�z �O{J<��t�Ŋm`��0o�=�C�խ�p.�6s�_C�il�4;Z��fN�Ј���*��%� �D��p��Q_�M��p/�� �l��<�t���}�%7+��J���,��;o%���fs!k��뺡��r��N��-e0�e�߅ϳ����ϙLp�i��N�nۃ����k���9��L�M��?!3�W���먠%)�}�{N���ڞ��Js�D6����S�=�x�ӱ��7�4[�sL-��9��(�3��O;3�D�+"Z�t�4��6<��!	��M�hE��kU�]FS��֣W�g���g��n���e.�e:�W�f��uDj��/4��n�mq�{q���E��J8N�Go,�t��
;EK&�R}�\Ba�q,C>-�?1�D<.{�ns-8�S���t�Fa@��9�O��z�@�ҥ�s�Z�ܤ��n�j�ڛ{u�?:�̧Qb�3 ���wT �OQ�p��=9��^㑖<�J�@p뇑~�����5�S���D]�ZѢ�頋�ޜ��N�ئ��G�F=w����L��2κ ��;�5�qFz��+Z�B u�i#]�Zm�<�q�h�#*�Tԟ��&��!�c�k�����������1f��-��YCo�{�ó˦�ˣ��D�.�����(�{����w�TS�t���%�b'=/;��$/
��&���D�l�jK���^�keTx�J�t�c�� �rg-�v��L�,i38��K�˼a@"�J]���[��/�9�?�l�︲��2�	�R�3+˵�7�r�>�a�6`�����gv�{1�����+��,���b
爣��9US}��]��Z�a������}x��6��]�����"e���첯]GaF*�� >��s_RƷ�T����B:f��s�+~s��/�x���]��7(^��-�uf�f]l�:��fw@��Zkc�{�Qg�w�<����s��ɞ"�v~7h�����F��Z_@se1��7������R<���KWNS+2��e|��S�P�o<��p�k���]4�V�eM8u�WY��(ukV��7��V3��!��ir��ʧ��3�6s�XV��w��t��4����[�T��g|[���-�͛J��H�EŃ��$\y\*0(�G)ߴ�lw;9����b^u�]�)�A�e�P�S��l�듥���B3�H��n��!�B���n�1p�{�6�2pU���ݾi����#��'�m��M��C�E�[zzYW8t��O�%[��p��+Sk�ێ3����Ŝ�9�]#,���i���>��O�r���z:8g��
*��I�M��fb� �j��o�q�z?�E�6eBE��d��s:���hd�aAs"*���� �����5��wW�[���[-�~� ��f�Q��HRJ�CkMZ�"	Jqo*Vo,��감�\˻��No"A�7U[�.�zS}$`F?d��~�O+�嚝�ךʆR�ѺE���\ƃ����2��cB��V�n�o�c�qNE���q��/�lU02�����ןVd2���:;	��$�Him�Ӯ�8��>��(�j�"v!9�^b��6X�W�$\OtءLeFٻ�|�k��iҀ�W׺no��6:�:�����R��tIr�X�c�h�ϛ��2��ܳ�GD<D�T� ��ٙ�3���J��xDqϏ��l�U0&Wa�;^Y�!�]����\�[�VG5)���[r��s�Gl�NG��ss��>�ɑ�o� e��`�Ε�V`=�㻿dT]`�ZdqZ�꡷��9�5�d�z�٘Bu��\�1�ÙK��m��Hϧ��ŹSW}L� ��q�?�o_������ol��� �t�O��"�w��Lꕺ�56�j�)��h$�"�4pV�d���^�zfm8�yfv�R�'k��>���λ��a��;g]�-����Pק�h!_��#�n/-o�֩��e�8�{�%�1��;��C�keXn7}�N��d����Z=k6����!�j���[�P���S�k-o��,EESv|��бd[��xWT���ot���X�
U����0w��z�Oc�x�5��r��) �P�\ٝ�3X�Z#8wi:�ֵ��l�];0O�=�;A���ٸ�`W;�6�6㏭~bg��:�G���+���ijVaa�3�Fa*�hǕ��ϵ/���z-�`z��&7ge��[��-�����u�{z�Fݶ#F�cD#,��#��cR�w�s�[�Ve?6��*Z;�]q�wCxױ���_��QܿJT�z��Q��6�頓ae���R�x���<h�L���O+�cS�	s�NT2T�d��0�r~ù�����ۨVE>��Y�_"���3�qc��s�`��0.Y����ϩ�;-O#�Tn��ڙ:��OVW���*o��7'a�OKu0ڎ����[� ��U��+4'��y���ݢl�]ֵ��kfs�_tGq�M��4�bT쳅��k5�~Fm��,���bY��he�%H�R5��l��a����Ȧ<�%��"<ҡa>m�������N���S��<�Ns�@�l�����N���_�,�_Lx��� �� B��jߍ�:���F��7u��t�ay�.2Λ��sU��D�1��{:m�x���ߖ���i{#�*:x���Z�%If[ͿT��v�\�k��h�+*REe���Y>�	.{wy{�zʥ�߸^��]1�p��+O�T`;s8��/�}���a���wZ�98�<����������	����� ��|����RM���l���^��xaw�z���3f�v�K�&˼�]f�u������`f_L:.'�g������*{��ʩ�����<������;��L����9̓��C�\s��/G]~�*���@l�k����~�k�O5��Ut�e�M�z�q���骾q��\N�%�S��{*WlP�+��b�1�i���Q��F:i3�In�h��{j��9��*6M��28q� vmO<^R�©�E�=�#�pp᳕�y�۹����oVk��(�$R��h�w�y��5f�~-� V��_�#-�ث��&�ܾ����M/[/Rkv��2�A���
_�@��Y���;M;�����)l�m=��U�Ql�;h��uU�i�m<���CWr�<v�}B)��O�s�&0�MN�Oa���	�s�_0q���˥;�w�m-8ܟ����t�o\�W��B�5[DX���u/�_p�lLe���J�8�h,ѧ;��Z�7؟���X�����N�E�I囝��c�8���v��D�?+0�!��6^�ga╺�4|�r(��Z�\�M#��;���I���fy�Ⱥ�l��������Y��ms���2¦3:^e^�6F�\�oR����:���Γ5�xs$Y�"E���Xѧ�۩r}���%���FRݘܫ�9�)}��x-�Tfè����0O���7?e-��~�0��SMmn*�7'Ʀ�&u���)n����/.ˎ��2�{�F|y�J ൫�H�y���μ�������Mlvo�Vw�k�l���˰v6�
��������c>a���'�ʅ3Y�f%��RDN��r4��s��3�u��*r	jO�q�{p���V�&�7����EN1�z���n6�˧�,æ ��@����|��]�t�����c֞�F��G���W5�Y��3��#��jq�����;���`Lr�B����~f�kb���>���[~�����fF�~���=�1�[]�"�9��Ƙ���]��(^�oq���Dc�ՠa2��r�WQl.6����']눖ܙB8�Kۘ�ؠ���Evs�xg>����(wԕe�,H]Ny+���(���Y�#�J���o;C���Ny�φ^���W'��u����=�~l�'Q7�Ԉ����lR�l�����?~y�Ʉ?�}t ]!��uKՈ�������vVe�+��Z�)��ȹ͹1�"�0�/��N�f�r��f1��fp��M{\Fy���{7��}Lg=гfwX?�͐���*��X�;�Ԉ����;����8r���63I4��_i}��Rgo���ޙ��~��,�씏==�Ej�T`O��њw�*]q��'��W����_�(�s�k�xe1��M�[-����f�h�eC�)�"��U
� V�X�5�T�O;�u�Ѯ�U�o=�&��6D���Ȇ��Zr�B,�S��k�R�^\"�t���]ENA�T���YT��2auu sT�q��t���GI�Lxڎ��������L��O^�c�:�2k��N�Ǯ5�%���v=t��|WL(��|jvK^�]�oF�YXyk�{�3�*zFp���5�b��s>�9�anG#-nψ�t��|Sb���t<���^}Y��[#'��蜥:*�u]��̿���x�~o���9D':(���[��YM$\4�M��Tm�������]TL򍮜��ޡ���?ynO�����Jx� N�u�y��v=�/�J����W���˻�h�1�i�z���LlOR�O	k/�1��������飰˼Cj����E�I�!���ђ�'��.�1�*ʉ��b6���.p7�����N�w��0���
�i��΅1O���Mfc�2u0���i�s8�Z���o�Bbv����v��k;�һ���z�E6���s�H�W���`Z[� a��Dz �{��{ڡ��i�jŻ�̵a�0���[��ǃ��]���[�r����ۥr�.� ��x�,)i�l�r]w@���՛/��[3Yאiw(wr�ֽ0θ;m� �+Y�/�������5ܾf�^�#>�����fś��Wnvx��W[�;'3R�qwA��%�R�ӳO*�^�ˏ7y1C����$�R�n�g�Vۗ�A�ȾP��Q�57!��ȝGg��V-z]e>4u�^߉�	���<�.�o���U�5��*�칙�#�(G>:é����&N{8g]��k.�ј�;�E��d�Π8����,�������S��*�K���Β�V�=�\f�M��_v�}�7�������v3��%���vk�s���z�}��ݧi.T�jY* ��]p��.��VɴM6��T��x �V��t��0s�u����F�O�[yOx����7%���+,�F�C���X],���FűB�꬗j�:�+�&��Y5�B��KW-w[,��+vF��9��x(��:�8�%G���đ�1�ў�gK||Q���OZ�X�ql�[.	�u֬J�tf�#���q���Γ:����G:#����x�!��&m�}%����#�_(<z�{Y�t{�x7�g�w��@�%v�=����Q��mwt�zuFѬ����׵d��O��C� �뾩��nƷ��Z���]��?��Y�[���/�{O[za�"�XJ�t�x- �s��W�˷u�6���S��W7�Smh�ۨ�˱[i�m.g��ܯqv���YؖnU�Xfq��`��j�\������>�Qہ`��W[���]��]��8j�%vA���jy��w�'5C((����[&'�n�	.ڭM⭕�f�+Iܱ���,�^*3h�X�&*�9�F=�e]GZ{�qn��&��]�S�g�����O��`9$�G�j��ՂTw`/n��Nh2@�o�$�U��V�8;h@rh�E�ׁx�����#���-�lC�R=s��wTB�z�@����u�
��r�v2X��Ԣѕ�I���f/�<�ó�wg;�>�l-�C�+ׅ���� ��l���D�֖*�m>��Ymg��q�R�t�jc�7ύO�<�sKA�J�X��n/*��N��-9Q�	Rt|�ˬf˘�Gc�dnܬU�.Ot�	�{�bv)���Ü)�8�J��i�8��Z�ps�~dW�o��L�n,'
��� ׺�V���M�W ����0w�ٽ��Eǉ	v̵���L�ˢ5^�������yx���aοvR�I{���v�>���NA!X;�vZ����&:��T$|���%��u��B�u9�����L����P��}2��+�F}T�J'�>9q�
;9&�8TN��g��i[Jq�M��1��;�;6�߷��l{��,!�n��fc��ob�
#�@������VXȭJ���EV�QeJk�*(ňơIZ����T��1-��1�QֱX�X������AEcV]h� :���2�
%���QYmDL�H(�R�EaQ�PUX.h�B�e�(-k�X�ب��u*�QJ�h��16����V#QR"�1�Z�YER�L(�V��EJ��k+�"A����Eb���h�iiXʖ���TEf*��m�d�c�֙
�"�X#fj���*���"�j�W%3(��F�XV�V"E* �u�R�����X��5�Pi���)ZVʕX�3�M��rU���1"���*T�Ab��b��J"1c$̨�"����#"��U�J���Tb.�Ԫʙ�Z�F#Z �1T+*��s�fQ�krTV���Q�(�{���|��}��;.��s2�h�u��{8��l�`�ȗ�ⵠ�>4�Y�K�{%'��� t�Fc�R� [��z䓥��?����٭��o{��t���n���x�x�v��j����b�Vl���L�<���F�h��.8my�()��Ǜ(qw�Y@c�7h2�l��Lkb���U�t�c���{�"�v�H�[P�b��>����n���ބY�Es�a@T�>���w˓����u�[�N;��?6K��n��{,���
�W���z��N�&��ݐ����!Z�V��>s\8W>���Lpy��W(�y]�GKR���?=�;M�,h�������ٛ�q@�w�3��zr!r��#V���g��u�}7�"u��G'��}�vf7G)�.������9���}E��ӿ�X�!�y��P���cg��X�D��5fs�m�����nC�/�m�A�9���	jy���\%�M��������m�{�K�TVe��gT{(������-8
uB�5_�!�ǟ��y����;>�����L<)�]=u��"�dk<=�E���c��G=�=-��j:
�a�2�� ,��c%-~�b�������wvw�������#�i�8S�lW=�R��'l�Lɫ"��0S(�Sħz9��x�_�Íeڋ�g�
���=��)#����fuǛ�{�,�0�e��\1��R�3���5(���f�j����˵Y��O�Mʝ40��g�,ו�˘�1S�IK`+�=�٠���pR����|:�I�螕L�%��C'����c�\�T�u���!BA� u�Un��i���=�#,y��d��R�]T�CJ�e���O��E:���x7L+�����tWzk.��x�F�)7��m�i��px���@�[e��i쬚�։M`�8�p�#Q�hp3��YN悳�p�F`;(l�0cy��5�	[���\S]��������`=�|ʝ��>I��̪�h�u��'�/):�����x1K�hW_��o�	��v�bp�؄xK���d:.%��g���v��?*x��?d���ݕ�m��/M��ƫ�k�S}�w�����;#�9���\Kr��ӝ@�A��s��2[���/
0�x�6[p]�q���y��F<�h���Ψ�'r���n{��r�1vu�����C'-)���ǒ[s��3��n�Kuz�6L�8ӑ��P�y����
��{,F�.�s�_9�+Ψx�h�tE�8���Z��h�5;�=��Q�w�y��}E�?
Fț�.y�������4M�ii�~�<��j�ۡ���qý�o�9ɳy�4�ݙ6��jd ��M���Ɨ<�>�������_�s=V�@6���N���rW�͍�Y�{���t�s0��w][}��0�Q�,��t[�w�۹�)
ytܥ�?�~��px�7]�	Rx�`�z:ljJ������ڟ	U�ș��`���؞�,�y�U�q�
F��݆�]rx��!��'�ٛ:�YOZP��u���	���,ꭨ�J���p9���"�zw�?a=��n�e�:J)�W���+ Y�����5�OK�,�z�6>q�k����-}mGa�e�E���2��sP+Ns�0�����:�M�1x��JY����� MK�^Z�����0���� ����.'���YDe��R�jB �[��8'�Ӣ@̷��x>��M-{��e�'2O�2z�r pV�VbL:\K��;uaVJi~ U�S���!����E�=�Bm��{�lJ�}�݌��C\����$Tl���"�t#�{Δ�ܪH�Q�N���<���h�##�Jn	j]2�)�I���I�lx�Y;�wl&�8�ۙ?@t��y�Cy�YC�#�D>f0��Ge`���rJ�6�����n�9q�)�`��B���JG;R��t���R�G�I0�98�|I��h_���~�X�rȖ���;�㣲��̜ý�+6t��(�R��R�ML���Z7�
hs�ʥ�M��k-q� �s��3]s|s�h�ىLc�"���=�6e��6t>�ofQ���郛��@�۷:����nyF�H��e#��&��7u�f��PYr��3�O��\p�3']�"fOA��.�Yk�\�Ç�N�������f�Ft�no��r�f���Y\�ѻ=�|� ���}���n:�}�Qpb�oet�Q�%eg2�͆�yf�e�9�#����Z���Պ�)��g�-�0�����x�Z*�s�v�]7x��(�B��:�/J�l���n�DX�W�OԳ�������͘��z�����3Vs�Z�k9�c�k����O]�r�]�'L�{%#�O@�DZ��Q�4�h��XI�iw:�CȈu��9Yφ�s��l�!�l ��c�=2��l��[7���(�9�)�g@j�cg��w��x�h���62ٷ���0:�֙jw�G[Ȇ��Zr�Ǧ0!���R�0�T�n�cs��ݦ�@M�tKSi�j_x�(-;���(�;��,YX�������:�Gc�lo/kL��<��s��! ���8�X]<�w�S�Z�YP�}��Z��țnÍ���U�R���5�}#�ޛ�z���anBFm���� \�)�L!���זj̆Uu�C=;��P=uc�[y~�FmKIo\b�7N��q�w)���6T�F��~$��C��s��A�FVb^XR�?K���R��S�b�n���oF�ݹ괆�6�x�v���Dc����sԱc��(�Џx^�������.h�(���������~�D閮Px�\�	N�Όc��,t{5�#'���g�a�#�R��借Ax��+�*�,��!st��z��U�(�T��H���3�ʖ��o!5܋sƜl�b$-j����z��͉�f1Bm�_��oG�����7uS*x�	}�����H���v���VY%6%ϳ�[�^�ݞ��9X�lB3z� oiwǼv�
ގ�g0�Y�=k����F|vR)��,��%~���u��Jx�q؇B����Ⲙ�9<(Dɫwq+�d���'w�_3���K�t�q�*##�W����w�~��x��ˎ�����G��~�DU�R���H˶�����{�*��[�#��Z�_����p~O�����oZ� O�������s4��Z�'�#������{.��V#0�&�D;���sdwH����ֽƵ��ަ�s�6[�}>�q�-���U<�LvL�(gf���)XO�tAi�lc��NV����1��z�`M;��k��-���x�a�1�{z�݁��_��y:��|�#��s��� �s��Ƿ�]9���!�d^w��M��n�B�����\Gd��sґ��UН�Ph�	���k+�i�;�l�޽EU�F�q�3J��d�q��Zo���Nu11opl����+/;�B��^	{݈m�;�l@��|RR`ٍ�P�~n���+�%�V��'�_Q�xolwAf(����Ԭ�8nU�:ˇ7WIۻ.r����x��{P�4��e�i�t¡�j.��vKl��Z�TH����НV�`h~��΀ttp�;p��,���P�m��rϊl	��<Z�#�*�hR�g�vx욛ݣ���l��ZX���7�"��uu2h)�hz���+��q�
22������iu{$�^�[���l|��Ց�O��	�|:���ҩ�w?eA�iMnϡd�V�w��lN���A�T�j�G7��u����n�	�����#�v��y�F61��n/0�%�n�h��S�����pŮ'�^M����eF8?m��!	�� 7�ߵ�u�Et�H�SwkEf��Y����� ��d^Fq��٢��M��7�<��Cj�o+�?h��fx��T�3��s
�>ڐ9������r�.tO���6��c������Y.c�P�Yqnd���-UYO}�p�89��]�;G��Θ���� ��a�q>��?�"݇��z˿����Q����p�ӷX;���Ϗk��wz�M�2`4�<�<ny�z{f�M���s�܎���pD��v z����n��w^-�����c����uq�r2��A��xY�� ���Q�����]-v��ɞ�M.A���Q�V�W���g�w�j������F��-�H�`����s����uA����;��ܷFKu���lh[YzX^�+q���DGm�2Kѫ([��8ׄ@��}�	�_<�s~e�%�]��;�t�B�X��ٙj�'~u=C<����W/�rӁ}-���P�m��/L����
	��U�̼̱��3��dt�fZg�c�w�\8�E�)�H�fW9M��|�沘j2͎�/9��O��5,kR�=�K��=�`�<�]}:+��鞻���(��t�ԕS<�S��i���k�\%B�|�@�ǵ��l��[���溃]J�]��+�"�(�A=6���
ȣ:P�.��gY��FP���p����s4�P[^t ;OwNa�O�e�v[���[�8��.���@I������>��L?٤m�H�����jy��}�a�k��z��x�,��I�/ P����i���0u���Ɂb_��
��_=O�l�f%�:7M#���H"T츸�����EkI�j�hM���f�S� o[�o�2K^�q�Nd2�{�FO=���'��^���-wH�:�F'_���6oQ�܀�Ѷ�f���2����$���VV�؇e�}C+U1eS��g!��.�O2b|��t}i�¥Q�4Y*�(Q�F�������z���_*Q��V�����6r��<B�D��u�	�=v'��i��0Dc�����nϨ�z.���T��ٲU������n��s�Ta��֎Vk{t�;��s:��]RDJ��"TAO}�onE�U)�0%�?a�T��iޫ�oX�s1^�k����	�X��:y�g�� ��8�5��$��U�Әz�y��0�h�M��E�����k�蜎�Ol�-5�7�|��sϷ%�u�L8�Gk�R�Ow2g�E(����`'�7���eWQ�e��/p�l�p��r��q�z[� _�U�UŴ��"7�s�H�=���ab������kv���㏎��s��"w%��rH�9l���U�q��Ý:{�\P����D�eFC������a\�
�Qw�7�{?Kn���I���2cc�v0�n��cF#�/B3ݗ'�����н��"��a��{�i����Py����U�#�_B1�JW:�w:S�ove7l�ӭ�q�����;>�6<����di7�)���vx�Mq;[-��{��6;��~5c���c�=(���ꃥ�}���(zE;fw[�D�����s.Mb��qE�Ĥt�E�ږ0n�џe_�R׋*��!�]\Q<�u�C9Ҷ�di��<vk4��&>[;�;b���8�(T�U����miQ�_wR��57*��^�,Z·�s�~�u0��V����';7[�it b��N6dk��mS�m�	'Q�t7��$u�<��]�-l!�ϱ������Z�0�9��R����;Pys��E�Xtwd�5/�Ϛ��Zr��t�b~���C�E]9�����r`nmi�b����T�s�����\Q�R�}S�ϩ�-y��e>ލҒ�EKe)��s��5�ԫL�K��W=<r�����	�w�|Sb�B:��^��j�.`9����'aي���泯�{�a:f��*Y��H����nv~F}nϡc�W��=ۇ;/,;�v�4�V{�У20q6��lS���x��Les�r������*Y)�F�d��}��q�_���7r�f���
�~'�m�iF����=�LJ�2��0�ӵ��[_���/	�����woӎ[�^��Tz7!��\�.p7��������I�2��kE��fl���mIs����oi�J��?Ⱥ��%?�׿]#����m�u��'�����/x'��#��`��+�e��߼���6޿�LP{*սR��%̈́�75r�-��S=v!��4[.�jjN��=c�ά%�<C��i�4ɽC�٫�M,�}@>D�u�Ŗ�S���h���u�y!˼+��S��X�l8�[c
�=�_k��1-@����0�C�-��oBԼ�݌�u�}����Ǥ��:�?��w�'��s���ؑ}��,�@}+���e��&�׊����>�?R���k:�_�P���4f��a�����r��~[OߣA
?~�,����U�E�WD�Q���<��E�h^#�J��,4;m�L�8��:�! �T��Q�U{�J��_
^C<ŏ����ܥ���F���d��c'����|g��d8B�:h-(>)�G�z���]���(��Mo��@��l��2��D��
��D��膔�7�6;��H�:�ح�{:�r���oF��Ւ]0��C^r(sr�<v���)� ��^��U,/��娺+�d�%��93<��j_���-Vv��q�=���Y�g�S�e;龷!A^�P�����g�6�Ξ�}dD���Ӗ���	���:4�c�J{�t����5|��tt7F�r�������mHb��=��#���n���M�i��Zs�Y�GiѼt�MN�:|�e�.~0ʃ��¸>�s�-�C��lǗ���z��%��q��
��fy���n����^u�]�������BO��	!	'��$�$��$!$�HBO� II?�$!$�HBO��$�$��@����$!$��	!	'�	!	% II;�	!	'�@��$	!	'�@��YHBI��$�$�Ё$!$�@��}���)��l��h��9,����������0r��T��QTT��
RU@�P�H$Q �l� �UJEAD�(H���
L�*�u*�QEETTRUD��	*�f�J�(>��(��skKfl4,�։U�
��![m�ئ�!V�*� [�V%� l  8� N�ؘ֘�CP�
�N c�1$m� ��l f�� ����T� �U(��
��U(� ��` n��� 1 	R!R�R����������m�CPHQ���j�1�H��Jr� �4���m���h��UR���X�Q� ��Wq�iI��Ui����SU�$�l�R�TT� �]���L�����f���"i��F�"%p��Z�BX�UZI���ڠ����1S!A�8gak�j�R���ڋLQ�*�3.�J  P ��eJ�@�C 4�b Oh�JT��bh�� 0昙2h�`��` ���T� JUD @     Ed&��2#�Sjd�D�xSmH$�(J��S M4f�`	�Ʉi�o�F�o��W]��.���	������X�(���`eF�EA@�T�?0�QEJ+��}͏��r~�&�â��Z�
*A0#�EL�Z$p±
]*�����m��j\��s�v��/��e	�fCG�{���d����H"4GM)|O[�U��M)5N��t��0ݳ��i�	&Ŷ�[y{W����^;�dCR���L&�
�[6^l���f��"��&��F�!��5L# Њ(͸�5fS�i]�w�h	����)"�ܽ���Q�p�5��%����fŅ<���4�X�GƊ��4���2�sQ�:G6�c��f�Y�sJ�7��1b�7�(�j��W�yRbٙeM��C�:�	��$��
��d�GUʺj�,�`-����5���*vU��X-%����ƦS(%�d�Uc�4P5-�H��oc��N�N���i͔�f��W�~r*U�yhVD\QX����1�h�T�bө,�$H���q��ϴ"�\{�V��˂�)��s%��ٲ+I'e-�1\*�L����ͩ�M_f���-�ἇ	����ط�
����dV5��Vŗ��v�%�.��͂�J7zu,r��[b�i�q�7���@eb
�N��5|آs&�1���u�B�]8�6(,I��5�d��T��[����P�t�!ih�9��Du��3^��z�V�8�m�T��-e��e�!&��$�܇1�3W,��(�Ui����]�$��h^����n�֬(�6&ّ�2�&SM�b�5f�k����pK�R�/j56�3�ۇf�ƾYڻ�%�.Im7IM�g�����cBIQ�yZ���Q5E-̀���䪐�4<�,�PRscBY.A�[R=w%�b*5q1�
nхY��Yz��C��]�5'�4��Z��nMMְZɖ�X��Yy�������ٓj0��L���@��5KN�y���$I�ѽw)��-ɶ��H�RR���l��;]K�ے��*b%ݔ���*^�E�bUyi��m�m���W����̆k�N#!D�T&+6
��õq�XƲ���4���D���e^���8Lڲr=uO(�ʤ�`;�ҩCA�����Mټ�gZ6�S/18��L�cwKߦ�N�#D=��(�V�#TP�8�*1����cfU���*ƌ�� H;���)�l���xd�Um_�p���,�KZ�lU���-����26�W��3E+{��Z]��78v��)=�a�Xu�f}��+n���˺;ev`���b�#wbǒ��/�̡��	�
�%㴦2��(;.àX�E݁�@�5j��#1��8[[��FrT����?e��X�[2�X��d�i��M�GJK.���pꎘ!P��e�rĬ��挗v�k+��$ǂ[��u��SV�f���:0��ܛH���:�p�^3rE��bV�׊��Ե��$�ǟ0��2U`�8�jl:�T33���u@�wUeݻ.٘Ek&��N�ii#QڭJ�=�,�!��cH��[�TPY1͂{�ƀX2L�IY��q(r�����D*z�Y�(]͆��i�G{�L�WNΗ��8g¤]�W��I�0�E�L����s&��1;�BZ��n�vN�[���f�^RBc!�����Cj�E;zuJ�3�*A�^���Dݛt͢��U"%���	b��1�.���NQŕt,6 C��ul,3+X��`m���eR��
بR�f�b5>.��ʕsN:8�S�SA~zql�5������8Fea�JIyIn�ѕN&m֬�4V�©��4FԽUxKY���Tf�'��㼛ӯ⊒�(�ݧ�Mo����i��O	��[���`T�m��Y�jRܬucQ����Ιp�n_�jֱ`ݠjGN��.=5�>��n�ڡܒè��	9#(;Kn�ޜ�(<�@�7�0��(���&�ܫ�ֈ0k��qb%b�Orc�Vɠnɺ�B���1��o
��J�^�2�H��0i������k�/U��+�5̒��u��i�9t
:-X�`�"�*�t�X�C��SM���W�0�ok�I�,��GMVM��-z�A�u�6oI�K��Td�����NK�WL
Nf��LL�.V�!�m� {�۠��߳c�1ʩR�%�M�Vjv�f�jS2�83hi��m�WR^�f޳D��&�p�`ݰ��:�b�7v�:o\&�����c
��w RՏ�(!��r�6�:��+1�S\�h��yj��D�·c�0� mڏ	���^'��ї�S�ʧ��,'w[TT�1����QK2�gH��h�L7Z��Qw��B;"�h��+����t�B�;�R#J	���¶�C�#�w/�W��n3$eX�u7r�0��-�ʹ
nb.0	�{K;Pf#K������j��J(�=9�he�A{E�,���i�##F�:�T�t�5��`<f��؍Z�)�ڑ�>�9t���[+P��;Փ�Ę�ޫ[��5��*��YR��,!f7�#dd��oXq���7 �5�VT,��o)��R�&qh2��v�ݥ׆�BIf���oUk��y7�p��iyB�׵��j��A���V2������v)�1^]3���7����%�*VV
����t��[�Zr��Z�,���z�E��1�+OՅk��E�S`�P��)S�G2: ��YX%��Qʼ����`�V�CC�Ƃ����J�&�P"�$����cSp�kcY�?k���{6P�N҂�dOB��k���C}�o'�Ib	2���.�4j(k$�N�?�s�5���w�]���r��3ƻ9B��F�(���跈K$d�|��z��䙡�;��u1��I�n�l�fS)5�h�w���xK��)�N3g��O&e�D^�M�V��MMnfM����;�a�!|-�1:)����ք::�+���aӣ^�w��i�9�7L)��NdބE=sQ���b+�V铰�s�oE�ww�F��r��}�F,�u�ȭ}�CX'UK<O<@^"��(��4�A�"��ЙK\�gvHIr��;��G���1PV"�Uыn^���k�_�J���G����t��\�ͪ��U����&���}s��e\����2�xt���56�C.��ݔ-96��)�Lp�r��٭�z�<即.:�̘I�܇D�b+gI\�r�ޓsW
��5��U��GMXޥ�E��9T#"Qh�f+�}����{�1Cf�.PW�0�G�M���T.X�w�����Mް�)�uYʎ�5�?���\
�_:}G�H��3�����uS�Hq�ژ��5@�6����.�6��07����Y��XKw�j�[Yw���#�ɽ����3!��зJ|��^�ˊG�Ȇo32S��_d�����O4�C��`ٳ�b׻�D4���Hݻ�1��<�b��Y_����x8e:�v�x��hS�sgGK�peΜ.�o�����$�h�s����n����y,���FPȽ[�@�vpe_g|t�\��H���͓*�*�����{�AFU�S �2��m����ӊ]�������Ƹ]�'0���<�lw��`xu�)�!��g3?Y94	�?�83e�Ϟ�f��#�:(�����[��=v�����Z����ۛ�\�Y�uY÷o��oZw̳�-��]�׎%��J�Psk�ʊ��q:�MC/��� ụ�Bt����n�x�M����a���V�+H4�]������f:�ma�03(YzK�R�]��W<.)8��
Q��5d	yxP��.����L�Yٌ�l�X�.i���V��p|�c
u����[�$�}�՛ٜ��]��'��(�������.����(#~U�q��x��ۖe�m�ݥ�4K��7�0-� ꓫ+����gLg�5�}:*3ô�a�x8S�,��К!M�o�僗��7��7M��6��v���K��8N���gB�X���4�ނ*�n����&�'GP��v_"K�MH&rs�κ���b��d��l��s}�tZ�+p�1��v*|c��;{C����N��dwt��/F�Uc�˱̰�fti���)T�nQ�I����Q��w<|��XkoV�'=��$W}4�3dY�p��FՔM#3��oYo�F,h5��y:�k�*�.@�7*�*חk����?M�E�\��e��:��z_3��u�;c���^�g>Jh*p�J�������w�gy�oq�}+V�+e��*$���=�BُVg�~�F��L��Q�b�V�U�P�F�NU-�͓�ݮ��H�XX�<5��q�r�c'������s
��]ӭ�#�7�N�E��ns���:��S���Y�ZIqR���ؘ+�/�Z�Gew�+�Q*�u�e��cr�n�Wr���������N^��׏�O-9~�+�|��Z��Ѽ�ckTd ͕���P�l��nw�I�y�l�ս�n��t�(�|�F���Ԫ��U`�{���5�}&ffH�X̎��4i�����U�76i�7]��cMˮ�/��:��*Z�.���}]�h偪���t��79@1���#{��)�w27��+��ز�=m��B�-nc�ه�ʼE�F���y�	\.��n:���b���`���#�P E�7�0	����ɸ�T�i��Lm���H  ߍ�-k�Kwd�T62��2�цC���	"�Dt��Nb�ھ�
��s^_"�S7+.�)7(7��ص�T9{1�)�����W���=�r��V!c$J��	J�!����]���V���=gH(���)�	��%b4�V\�m�|�_e�8��X6-+��k�� �k�:P���v��ϲ]���*A����Uw��M|Ԭ�$JE�Yb�L�����8C�]"fS��|v��	S���v��:�VYT�=o�S�b�u���#�y��볧\��\wt��Zw5��lb�#�2�5�']�\Q��՝��b,n;��=ψ�]>9�R�bv�4{�d�8�7\Dr��ܽ��]_>-՟�.�R��83����\fo��+΄��1;��b��Es��,M��.����j�������X�P�w��x��a�r�+n�BCs/IW)�EJK�2�].�t�^1��ѵ�n4o��bW:\���{�9l�Çr�{j�d��֗ujsٽ]�����L2�(M���J�ݝA0�hY��D����c���N�7�~,��"���Pou\��,�G`���~i�M&��̽�+��b��+�W�CS6vv-f��)���tc�d������Zu�6p������b�p�T�d��յ�kl���כ�A�^sf�jn�ul'/@Z���̴��ٔ���Mi�N�k���Bh>��/�Bō��_e��9ϱ��zY��J]hk0L��ڏ��MQ���{nN��S=�4a7�#鷯Y�'N8�T3�~�QSN)�j�
���@P�8��E:��M�������'�� ���>^��C$Ћ�Y�^
��3[Yw�:��A�PMr�L�
D��G=�.�������ݵ\�*B� ���e�(�����E��YV��*�P5�1;�{(��Τ�2��T�."����W��FS����_q��<�l�Mf��������_#z(bSz�Z�d���7z��V�r��ō��i[ӱ!{�v#�ґ�Ml��:I,k�!TuzW.���u��&���NHZ����C��{�F۲H*����PRվ�u$!>����Q��Qn������[8�Ɠ�ӭ3��\�`p(`Hc�����4��Nf�c3fa0���d��:4��3]��K�]`6*�f
��8�Q��g]��w�e�p��46��ݖ��U�t�$to,8����؍kǫR&�d�B�!�N�λV�ZL�M��Z���8��zvd�J���ko1�)m;�s*�Ѫ�w�t�0�$N�f]�⩚���1MͅWè;�n�-�Ҭ��j��fwQ�ۢ+\,Mӽz���b�n���� n�7Aj�/S�ݗ�*"2]�ˋ�R�R"vG�O���˯��W@P7R�8�p��=Ro	Օ�;r��_�Ԝ'inBfb����}b��[Îw[.c��!�P<�;�lJi��ʶ�����:OLM�υf	̄�|qޫ��r�R�Є���X�[WJ��+�n�t�p���e��{�w�6�[�ݱ�r!�� �k@��������"�����ZC.<��ma�T�U^uoF�u[S�7wap��f�y��X]J�W9:��j�,��J���	�!����ө7;��sc�H�8*��t�����\o��ފ���2�5W����#��dT�f�|~4m�2#Ʒ7�t�h��F��Ψ�m�6�˽���TaU����f�1pA���g���"�'����m�@4\��s�-�9Cs���l�hb�%+�O�J�7��w�ِP"�RgT8
s�i��=�[w��B�N���V�S���3/�O9gc�Z;3U���_��%��rȷ��d�u�5��aZ�xY�Oq[��P#�.�S��sz�mk#Wf�6��:���GL#rb{�b���2B�i�Q,���M�;��8:�/h�|S35/��F�`��_lp^;���r=Î��t�g�_pf����ڐ�z����m����in��13��J碌���,��m�l�os�q�]Q��4��]5�L`87*������o�򕯚{���`"lڸ�0�VN�]|�[�l�ĺ�V����� ���o8�����յ�z�Hkҝ`�~꽽e9��j�4�2b��D2�O����4�Z��	0fRצn���L m�W�d��nt�/tl"������N��р�9X�^`:L�W�E4���9�Q�:��Fok`s(]�=])�l��TW�*۩���e1�=,��	��kvYn�q�L��*>�Sl`6�Y��(m�wJv��o��v�Ci�w.���u����}m%q��t����ԣZ��A�� gT�F&�\�Oh�a�n�ː���r)e���G-�j6�t�����oop5�����4��z��wlאa�w�9�g&ذ�wKF��{��K|��[��(���J]FN��k;���[��3{��51Ƿ2������ަ�#�ec�jT����ϥ\<f�aU͵*<܆�Y�4̭.��j�{���er	�ۓ���	%`�<���*^˸�-�N�,qqdw�e	`K�;�*
�S�'�9�7��A8]��&�ҶŦ���]D�pp��vL���n�q=�}�`@�dw|�^:T�cC��T��q��	M�Җ�)��US{n
���:[·���=�C ����U��vҾn�X���1���l\��p�R�>v��(f3zZf�Nl��4�	o1���q��4��7��pn΢{�܎��r��M��dfu=���]w&�$ ���R\ �Z���fL�f��ȼ;G��Me�ׇ�1�X�`�<S�c�;�'[����rT�Bo-XV]�˪58�s*j̺�P�ړ��^��y�i�=qU��h7�0��D�j�9]:p�8:��:VJC������4b�{R�<&n5�&Q�K����Q�8!��e��bb�sPl m�.ᛤ͇���n��gl�i�L���ћ�s:0��GU%1�д���VґW$����3DL��������w�-&
��3��V9T26�´���ƚ�n�;Xr�K�_L�h�Z+Hev�^�4�F����2eJ�7��4�oEˈo�M�g7I��:D�9�ه��+��V
�M�]��.��.nsĶ���r��p����Z͚���G�,\���nvh��{��FRՎ�u��у
{���Wy]65�&��<'�@v�+��ոx�<�u���7g�s:7�7�,LHv.cLy�NU�v9��M
�2��7����e�t/v�ff�Qb;}�Z�V^)c^9q��f�;y���B�P���2+�e��;_dΒ��I�x	�u�<6�̊s�ҷZwٴ�҉o;�������VX��<�nn$�ԽOVj�/�+�EԵ_�r�yO+H7��ocE³v+"G	G�m���a�F�ѹ�8K*�bWw�LZ�NP'�`-T�(�劳����U1 �O�ճ��o�l����o�!vt�6ö�c&_�OȐ$$��_݁�0#�ۄ���E��cf`����F��~���Ǳ��a>��͝��V��kQN# |঎SJn�L7j*�!�WCe��:��N�z6��ʖ��e_wI�Nñ��o(ad�ʽ�-P�T���6��]���6�K(�#U�[ݐV�x��Lߗ4�pϡn]Z��i���K���yK!���T��0Cl�=V3ub�\��`�X��ؤu�[�8����śG�ވ<���)�� �`^em�3��(��)�2¦���+:�ew�5�E�?b�M��z����:�]�\�`��E'�LVo{V�+��f	L����:�
�@�=��[��|���TF
�,�
1`Ǆ*
�(ԬErʬ��4F((EQ��R,X���w
!��*PX"�VTD���Y1%ABڨ������QAL��e+Ec�X�b���1*[I�塉��n8�%Kl��,�jG(�S(T�eN���������y�杻�}^z�͎u�����8���ꓧM���U�VD��D<�������o��wA;� ���}9/N��7Jsf�`!]���sE��[`3f1�6��Yub���Bl��܌i��qQ },l�Sx��v*��^�>�{K�`��/b�����{2���������V�j7������8��.�����Ի��0~.�wR�gL7yڙ�+O1����v�q�i��Z��2˸��;pNӤ���!��r�V{��i�X�S�D�~�*z]�%%�u�Or�.qJf��C:�e�Ԯ�:ȗZ�<��Pg�;��.1�F��s�r�מQ��~x���k�4.�о�jѐ6ro�U���sБ0�_
*o_#9=nrk��{�fĺٞK���Ƨ�\�j��e	\�l�^*In�W�����aV��ܧ��|L�;->�,u^n�j�m��c��ֺD���Z���Ԯk�Wj]��n�H""Nf������ ��;�8|�����X��.��y��MwV��	�׈2{_��mg�]J�{ m�*,@�Z���T��7]_e�}<���J@a��^\y�����$��V���:���r�P7�#M�''ܳI2�bc*4�"���V�Pˮ�/,�����&׬e٢�`za��[H<u8��#�)��[����CR�}�,Y�*�?u�+tj���c���G#�bT`�7j� 1ZaU(Ib���V�������� ���=q�G���t%����3�=J&6<v8��v�'���LT��ˆ�g>���|���2��dc7Ո���O���������(���b�oB+����8�{�b
�������48kXnI8r����;{1��p�M��/�.NS�̤ )	Y�B5.�w�x۷,Mu��=
�`�5ԺcMC�혣e���Mވ��#����R�g�=�|�wH�W
�V��J�r' j3��9�(+����d�y���墵��h׬=RL+��њ���pOؘݤ��S�����믛W�{�h�W�@��s3��G�6�7��53qZ��o[zX�WB,yFR��]���s}�WM�fk�ή\kطs4�5�ꐄ��C���mKN)�wZ~
�9����/K��d��.��b�,v^.kk"^��O��B/��U*����[�'U��\�j;3�a��u��؇C|���z)�,y�B�q�����10�;8�_kg9ڜ�Q����P�^�ײO}�e�ȥ�{s�%�O��1��:�5�׼��A��;��ٽ�S�w�uK���c�[�uA�Y[f>��X��]:�t$�i�C�Сy��Q@p�����.:84��u�釭���3F����1���S/*ʜ`��h��Ժ�veṔn��\x���=1R�f3Ư��=���aܮ���V`�ԍ��"vc'
�kU�`��͸��G�n�dk������{[��x��%r)w��J�Ǟ<sN$�DU����yѯ`����r7��Ɵ���;]���k�<�B�(u�	��{m9���لi��q;X!�qy�fT�B�me�x��^d�w���31K���w���S�d9�K�������vj3��t#���΄zS�mm�O}K�`����
/��r�Z.�"��&*���2��{�2^jU����q�s����\������6Ll����o$��*k����Z<���N`��Ü��K����.�6y����q�y��{��+�WχuOts���k��v$k���<�3�8�Κ�ca{�������=�oe�#u������k"�C���u��:	����bqM��2�L���<����u,,��M����3Zx��ٌd�N`	+	j�޺�β���+C}�έH񄌈�w�)T���+�3�_g�KMԞ��Q��*Ћ�b�it��r��
�꽳�a�Xp�̮��Y�2��fƺ-���p��l���.Cj�7�n�y���/8yV�k1������Rm�'���>��/�/��c\~�H遵����Zc�l�d��0���vU�U�^(�3�"�ƃ��6�/{���Mt��ㅭ?���3�.�v���/��¡�ڦ%�8˦��3�O3{X����8%	�,s�#��H�S��^H����-��fK�Vvd�J�b>r)k�Bt�/$Ӝ-vؑ��j�v�>RͶ��OcO.㿷5d;�m��^�R�)�E�
C~��m��>�gsX�ҡ6�3��V<i�#`��B�hI�Ӂ_\"��9u��#��ݛ�W74�dYUS�d���j1Rl��by��8&mQ��ZN��m[����n_f����隼��
71Q��f&𕕜X��s��F��q���3�B-L�sm=#"�n+o'O��{�ML��up'0IWdR�ڴ3J.�����A+e������OZ�P�X�H��0CE*h�x0^ �Qk�H������6����^1*��7viՒe�G#g!��V~�X�#*Ȫ4i�I4~P��;�X��jۼwm���GsN��Q���	���(ur�Ăv�+$��t~��%a|���Y��׵�nk�������@r��c�a��KM�s2ȄJ̣D�Ǚl᫨ꪱ���(�X�
�޼U�oX�vpQn�$i*�a��]�{�e�#�'�*��W-�e��)B���YbQ��8�8�P[��5�G-TY���\����
�����J�&$�Tb��c��+ċ�K�%h�
� ��1���X�V��c��.�Ě���]V(kYT[`��X6��+KlXT5�-FՍ�.����O���۞v<ʜ6��q��u^��%��-������Q�>ͣ:�٭C)*1��iwS���%a`��͔/~�)k92�im��q�9�Ϫ��Ϯ>��֘�ys�����Gi
C%�ּk�t�V����Q{c�	�Q9��'H�DS��d����W:�u�h��%vо��I�{�:��vO�y�d�{2=�dPj4�7���p��|L[鏣E6��r+(�^��j����:�]�]eE�*�ږ��<��
Vl��b���6����2it�f��A*�L�C�U����^ŕ��S�6��%eP{�uz�f���G3k4�s5�nj)K�����<S)�8F����^��.�c"�ŷ��/yd`yM,*��{��Żx���WB�nƛ�'�#5#ks��J�Ss�i���������~���;�tʴ��\g5�nl�5��瓵w99�� 8��
�N~ow��������1(���wׯ|��翡�4�k�� s� ��|��	� �	�>��>��!=HgvC�'�X|�Y!�S�!۷܁�	�!�	�vI8I;�|O��㞤��'�2ä��YY�P� ��I�0��x�p�N����}��OXT��Ԑz��d9d;By� z�o�!�v�"���8���]��'lR�C��c>a�@���'I=H0��Ho�y�����^����X��ՋNC��S�,	��1!�!~��t���}�@��>��=d������	8dSC�@����w����~�8H�P���c�N>����ԁ�$>@5'&Y!FNa>Hy�s�塞�W�����s?o"���l��q��B��9hnvd�k>�]hk���ۉR/�3�������|>��胖@��� c���|{��儧�HR�C��=����z����~~�iф�'H��t�2Md<d=I� �{`ô}�~�I�I9B2p��!��Շ��,'H�VCP�{޿_7�{��'��2,��C�i$����C��,��S� $��V�׾��}��wŒ08dY>9�Md�,�Xj� ќ�01c.�N<����~:��!��C��'C��I9��p���$8�z�HN�y�}߼�d���!�0��:a� 釬�tm��I��x��&�A��2�u�~q������t�>@1$��|��	�!�@�_S�����:I1 ᓓ������y!Y�!�&&�����Z���E:�2a��x��I�=�o��=@�$���I�X)1�d��a�@�,R#gއ1菧��՟U��%�8��ҴRϨ�&fW.�
4����/sX�
����c��)B˺���^j4��y$�bC���C9� t�	HLa!�!�`�5�0� =����?y�\y쇨C��$>>�Hp�o��,'��$�r�P�2I���Om��{㎃R}Xx�3�k�'��;I^S������i$.�|�w�=>�^�y��<$�E=��	}��N�M��z�ï2N	���*���R{�\{�y�>��:a�>`j핝��Ô������v�;���Ϭ�{�����>��I��0�I]d����R'�	��r�������>�<����� c�Y3�H,��1X$��� ��;Hs��}��{	�|���$/4��g	8I7��&w�HfY!Y=a�!��̅Hr�v�y�W����>�$hz�;@��YP�$/t��9�}^h&����T����cn���1'��i�b%���u���+��6h���zF`���`��o%��hَ��ж�$����T��\�{L2�eeneꇮH�EK��4�2��1��z3�ʒ��o7��q��ص�R"�8%\��p]{�`��#�~�~��O�4�՝z\��>�b����"�������D>�R�ˑ1h�[���%���hOh��σ,������[�2�t�B���Q�w1ũ�V}64�[�I�vEΩ��d��m<Ql���;��kgW:���P،罅�jKQW�(|O-���z|ٳq0 Fn�����D(*v���^��<so�Jn�Dս�x��AP2k��3@���K��,��,��BO&��o���n�^!���I��z�,�^��Y��Ē�iao�b~ S��=yW�g�7[4}$�i�鷓���� ��<�9�/�i��_�eP�c9v���ꑗ�����,�߼Mh��(q[��;��t�KNĂ��I]'�pHe7[֏n��NcR����z��f�M�,���^=|��b��{ӏ[-�w7g��q�����W�	tϽ�Г
5�_�۠���pAS8VJ�J�����f�䞳b�p7c7)�5�T��U��ȶ�\6r1��2$�B��tm�����h땐b���*�p8�E�;9*���7�uށΤ�E�].vC�k�ҵ3���t�ux�9�&�7����L�	��ⶮ��w�-z�/����j䥾Z��b�B�};�c��Y����C�\#h�ǉ�ޢ��c,O\1�D��R(oK:��YZs��� L��7�ζ9̝�ԧǋC�Z���i��N�\�<!�COZ�X��OL�������)R�𹧼Wi�MR6��}���t�ͺ&��w������ْΨ��47�+�;Dc�R��"��׍��f���*�O�>�4���^o��4׫���I�c�3p��g~M�<U�TO��@�CF\|*gs3X��ދ����Zc~�}�V�L�+f�t `�Է"��-�)�;Q��Ѿ�1D��(��d�
ب�4j �0Eˤ��x3�V;e�\#^^�=�2]�c2��
�̢nѽrמF�����x?߫�M��l��Xq`3�ݛ6�e��賚���6wk{V;5 ��H���w�:�c�oF���Qaws)\��Z�)� 	�ٶ�4�itj��+(���HvH��I`�yl���󆪋p�����Mc���w�at��XXL�(oM�y�=BK��Ɨ�i�����,��jbW�>�vۼ"M=~�d�������F�N{��_
7�(�ÖM��%��Yy]�!��v3��օ�hQ>�E�5UyP%���eQl�.�I}b�Mo: ���_u�V)�[_�?2���6�^m�elB�7
�2a(��6�KS�D�f��HƑF`���d*��h<�DRC&r�7��ȱ&(��"M�n�Q�-B���T�����G�.}��5�j4��Ō�"����"^'F��І�*��E]��W-�wX�j���K�3UY�}Z��*�!���x�!^KÒ�")�YA�B֑�YMR�u��n%r��E�j[X�j݋�F���w#�eݔ�l���Nr
�RrӌR�&eJ%]�k�9��{����(��{l�����qEb���ei�1+��a���#h�ىH�,QAV1D�H��(�Q�Uw7+%w-��l\j\µ+a�\�e��r�;mF���a�f�&���q+�ݵ*cF�]n�CmQkP֣�k1�A6��d�[Kn�[��XcZ�e�H���&8��c33ߐT��?�u?�
i�Qr��+/$�5;���Oq��ku�
��U�jS�no�/`!k�Ľ�j��>w�Y��bQ�s�R�}S�>J[��W��.�)�9���F]vլ�[��I� �wz�lX��NZ��7�v����1��rD�g^H�Gec+ԕÂ/*��1�"$�Yx�]�;z:.����;6c���a�񼕞�SE��d�aڐS�����d�R6U����A����lHx���'Hy�k͋�uiN�ժJl�����{�8�s��_���e���pуt������]�Ũ��X�lћxa��S�w�}�~K�b�m1�ٞN>��u�p}.���<�ͭ:V��]����s}�{#Q'��x�Bp��"��f�*���GyFھ��14�U>��8�����rԓA�N4�eE*��ۿ�ʴ>�j�Y`�8i��ߒR�[w��'f��jϰnu�ɜ*ٍq�YK��\�5`<�e�}�Mrm�}��w��Ƭ��`��TÝU��kk�A�����]���y*~)r��V���FR�z���T���YdQ�����Z����>�U˞Wkp��	Ha�-#	(�;T5�yWz�M���#��D3F�#���6=�j���:ժ��D0� aX�v��eiU��a�#�x�
�=���6G�|��Q�{X;��h��!�cp��"����A�"-8zP�m����O�a~D�|�����l��Y�~��p͡G������F����h#��yRFr�Y�z�z���_nq=D�vrV�g�ְ���z=�}7��sN�6`��wc��N�C��4W��Ap��0��p(8@�VEkL�ae���~�0Α�Y�ᶅ�?jTF�b�ƅ7�Y���ׄ	�a�,�$i�f��{d<�r���uϼQ�fZ�!r|p�;zVL\��_0�n�Q��A�f�,��_v�U��}Gی/S)������ڿ���o<����>�+���ɐKCڬ���!�3�paÇZ��<j���$Yv������ޝV����^�9H�!�hQ����/�p7w~])@�83^��V3c<k/����U�%�O{/V���ƪEo���Gc.W+V���DD.i�P>����k錜�SKHC� � ���+�{=���0��K�=��<.!$VE�Y�_�W�?QhiÇ�cy�*<l�sw��ZG�6�6F�Mx���¨�~����^!��)�yi�7V��j'���U��"��hQa��qY�m�u��oz�����$_-<D8B�l���VW+� �mQ�����9"y�F���(����ݞ���S�n.0��7��2�� �{�پ�h/��҄^�-Y�ô���B�Kn�m��R���<���q�l\P��/ϑ ��8��R!�+�I%b3���E_Q��Ա }��y�o�^W���߀��:ݻv+¥˝�W�^\n��Di��%f�8���bb�Q{��]+}Z=���D�g�a?Y��aYs��l+Zp�j�{�ʎE��#Z���jvr���uP�F��z�e9�3�l4����g�_qv�Yp�lKC;0�ת�@���4x��F�\X�K���҂��f:�6��L����0�Nv�i|����o+���Q1�DY��+���Jfz������ �X�|Q�\��S�Ty���jj�:�&��������+�����*ЍWu�闳]ª�Nfn�#�����W�US��١KJ�xWTz����c��@^ ��ηQ��G��+<���J<pr뮁�/+:�/v�k�8
����u4kس�y��K�]f���F��a�B���Ưx���h���,�VQ$ia�<�Y�'T~S�׻��z�,ٿ+:��>:h�A��8y?J�_g�����b����W��Sѕ�o����gZ��,���Q�i�8s�a����HulRB��ZX6If�+�}w����i�^!�|��+:cX|��׋�~��-��sD��λ�}6������Nr�����I3�YS/ev�h䢝��[w�M�hL�Jȑ�u�Բ�%�+W����y��=�6��Y�>zu��홴�����wޮ�H�K�6x�dQ��(�6���J�������0,a긧���� ��@�}�60�h�:I�~�2��*��z��3�]����#L�0����G[�w�+���V�''%�:�a㤑G�A�P�=hl��s9�ί]`g�Y#H����l[�dJ.j�#�U3�U�z��~C�гD�x�f�ӆ��ŧ���L�+��$���s�/��o,����UyLXC?N�+SY�1��}x:��J��v0��ξ�m��}��=�F�żj~�NclF2���B��?3QY��Txf��B�CBl\TQ�jn����|�	�����d$�����A�XY]�l�잀򝾺�=H-�g( A�
bf�o��{��$̉.`��T���\aF��B%�B{�r�5o�	��$��,><BK�հmy<?5�U��nVڸ����EDձ�I�/UEǍ�"��0g���<FZ&��2��CP��j:�Ww�����i�&,�(������qy��-G;�d�du�({�hQa��m��4�럪�s76O�e��չQxv��Sg)�[�u�6��X�S��>��j��䥽�����4�%J~U�#f���J�l�"�Y$z-&μ��,��Z<��s��aHBȯ����=�f�sg����9}x�l��L#��e���=e��W�K
�z��lԧ����JAu�W���_]�:�?y3��#Sc�N���=LY{{��b�/��a���g\ayV!b�Y.��ZkH�k&�<t�j���XX!Κ�׽�DYD3g�C�X#uY���l�hG{U~�~�gCV~�Hm�`�ȻS��0��?W�Wu�����8�!��q����3��������}%[ѯ�N¹��$W���Z(-=\��W+T,����n�F����fN���ל��%1e���1�<��}A�m,y؏jx���'�˷�Pc�J7���0&S��q6뚴��3���Kk/U:i����2!��"��Nl�])��\eYt���r��U��x[ܭ�*PwT�2�,�|/F���f���Y�u8Ԭkn�d_<k�`<%]v8���,5·L1��_V%�B�6
��\ ���B{W�R�Y���[C�2����hi�1��z��I)���#=�ίu�wr����aӳ)f;�>�a�>���ʬ`�c��v�Cv�ۤ\�m4��d��\�fH�I��»E�v�he&ձ��U1]��yO2��iF���9��	�T�*��BƲ�d�ӷ)c:n�@Y��Em=W��ȩ�e��ǯqF�eY4���R���&a��˥����,������9��@��կ�0^��oR���Rv�d0���*�n���R��q�lұkFT.S0lR��[��j��1²�Qm���J��f�U1�[��\�1*KZc�Sv���Lۑ����sm����6�16�Xբ�Af\)�k2f`�bԮY�DZ���k����fR�ef51�Um��[��2�M�X�*�&���s��1�s`�K����wq�k��5�4q�ªa��<�����\*W�Z��a�19�3���<��|��O6�Oω�sC��[��ʕ����Y�4���s�<@?_��Ax���&hu�C���c����h����	T^0�6@A�MHU����B�v�p�Da�Dq��z^�vY$t�Gfb5�k���`��{MN�0Σ�ԫ7`R�V������__�.tk+E�����E]�Dh4
7���2񍥆,���,��a�}hY��ƅ7�sv�m�AWLx��J�h�x�4aгg��K�Fd��v+�dq�%*8a�CCC4@����н�+5��/ƍ|����t}�BS�L��钶$U5�5��X�ؼo��hЖk,<u��uQFq��l�QL�Ga��Q#Y��.��B�pY59��_W�}_{k�"�3p����X��D3yl?���y|i|��r!�bp� �Y�ȁ�c�\+P�ϳϼ���,��_��
����x�t�$�'���݄v���R>?*_dT_+:Q��}��B�G�����Д�DV����mp6a�6<s�xѣ�C"�K<�s2�"�!@��o��k�mx�kX��=��z�"��=��>:I��ve@�++�MF��T�],��40�u�#�/XI�C���Y[��M������Q��?��'hY�Cb���Ϧy�;}�(C����P�5eL�[=�G��{�w���>Ӆx��<4{NӦh��p���u׫z����b�����P�9 ��)��6j��<�׳>���^\p����rgM�hH� �Q�}=�h����Q���#���B��c�N��yx�K�s�-�.��a����{�>�&�o�O�Ahq��K�oG��Ç���#��D���x���,�G�HQ���"�NҌO����<%�GR�tr��
�v�������#M�7��R�XD:G4 ��y���vC$�|�p��]{�<.!$ 9X�>��V������$O[�R������:d�4&��8�O) ܭ�]0����J��8���=�����ӓ@�i|B����ǈ�m�q>��ˡw_�?k��ϩZ'�"`\sP�O�ȟyKP��|X"��s��7Qo.�����H�C�A!�½]{�ު������;�03/V���ǐ�d���]�ז�s�<x_O�-4}�
��}LQ�|w�	�0�9}x��Vj��B,��oz�ه�����]W��t�WX�ԭ����%&W�}�&p��[��2�/��u^Cqi�DW���6ha� <�6u�Ǣ8�7�IS�`��Rە�豕����v|b>���p����|�M�C�U�GQ��s��E���Dz=�'���2c��.�։���Q�g3�(q�W�[[Aj���~�Fr����В��g�Y��/�b�c��2���M�Z_Qա辆ȳ���di�m���n��ͻ�({�8~T��(���<|zv�]�Ɋ�}^`1��!t� �懍�)<#w������b��Y�ITS���Niy��؀f�q&�}ݵ��+��$ŝ��Ok#O��D{P���6 �bʹ@@㷾
�لhZG�#H��Xw˓<g �����R����d�Dr�,'�*7{���L�$�&k�ژ����4e��Q�$�<z���Ve�ڰ[[�X&�<�q;���س�U�ϫ�@���}�l���J�'�N�t󽜻�X6�}j���]Zx�)qhF��B�δi�|���w�LdǈE�CF�$��F�]Q�3�5iV��u ����Oe�@3�}���_2!yli�l�_T�T�ٗ��1�F��(��(�6l�HA�]�^�zj�UY���a��%�q�*�$]�c���/dSI7�>ld\B�D��Ε]���R�a�6A�m�(�qe���% #;ס��u�#F��yXhx�!\��!���Q`�4ZC�/syd{�Ov��]�ts���bøt�w_Dz=�}V�_9��s����P�!�{>��EXXA��}�Yv�7���'�=�ƃD)���E��<^QIZ�۩�HIDwn���F=���TAE�!�8l�;�JƲ�wo�
��2�G����x����B�㾗�8�u��<E��"�$�>:G�wV�e��l]�<~{o�kU���$���ד�k��aOX�V�r�0�4p��׫�9��z,�8ޡDY��R�0���wV�{C6l����a��%�%GM���_T��a�٫b\´����Q�Hm����i�j��Or�Y�J�T��;:V��+}�Cz�C�}X����ߒZ��UϮ����[���~��������/�?+Z��,��{��xQ�Lo-!�ŞB��:1��a���{������l��$~��o,,�ϒ�\�����qf/�C���C�--c/Ȭ���>!�E��-�����!����τ�����@���U��[�(ң�ҡݱ�^���c%ye!��� �Gh�2�@6еj��5�6�c0�\��<A�mT�nBu#�,�\a����N��V���jxqۧ��h��A�RS���9
뻲�wl����7 ����2�L���k�'t+�}_UUzo�cE�G��Aj�\ɦ�z���F�ݢM��g?0E���f/�e���#և�f=���Ȳ���&p��cc�N}r2�����s�B�#yCC[41�?y&l���}~�{������+����-C㦚��^~׽=$�9�!�(�F�c�&�,r��cw+z�Y��D!D?2"Cڅ�?"�Q��3}��1����6AQ:F8����so�-i�C��.��P���#=�R�V���~d���@!���Y��+2����!�׆=�aR�i�鹺h��FY]��q��أʝ)��bцr]�s���U�?w��,5����"0�i\_�4l��"��=ݔ.�
�� �v���;Tl���ge���y����8IV�mY�<���w)ȕ����l#L<�G��+��c�X���:���O=.���b�U{j�s�RO*�W%�Lۼ���u0P�>TB��+z���l��>����8�}�+,4H�h���s�|�����N�CX��V��$�ha8�qvNw�H�4�_x]z��������ח����<l�Fy6g�J���շ�s��ێ�7���E��2�>�ڝ���ZL��5�qխ:�S��`d��*J��y��Ze|��q��J�D�w6�]�����k��W��A7����R�yB�v�V7�%E7�;�7����u�B�A������w7ʣ�j;�iT��*��j-���w���C:Kq�Lδ��VΗE�bfY��lU��#�ڣg����:�X ��%�h�X�8�swv��'�4�>yH=��.�b��;����,QP��:���W�זހ&�We,�"X�UyO�T���5<s2����v��\��(j�Q��j�� �VP��W�s�b��,��l7�]��{��ކ�!|�Y^�S�������Qf�9����θ�����r�ʀ�v��s��ᾱft}3�K�o����v���n��u`1,_uݰ���Q+(�*r��gi��t�lV_\䨢v\K����D[�ӊ��P��"����S^�JZ�KX��K�
kw;m�2qui]K1nocՙ]:���lE���N�"�Et�]�X7fu��is�i�.�a�:"����Z��x	�]�A���ԍU��i��(^��.QAAf8T���"�k�т�!�ʁS�-�kE®��.҉��E2���კRc��c0�n�K��;�2�+m���!�2��P�[�[��2A
&�'ӆ�ehB���.8aP�W)�9�������u*��[h�[�J�\s(���LJU��n.e���\m�ƌ�-1T�b.�ev�e.a�9q�s.W̎�3-F63R��H��m4Q(\j$�Q��t*�N���'��:��Eݲ�٤�����DsI7cߖ���N]EOZd~2в	H~6��:y��<)�"z��!��B.�CD>��؛�|;rϏ�Zq!�C�8\@acW�!Dvs�e�}������O���/���. ȣ�v�^�~�!=�h?A�kXĵ��ZO2"���uԺ@T�6л+�,3�H��4`{��3�mX�V����t�$��#Zo��+Z6K�b�r�!�dP(��@v/�eR�׽���j7.`*30�ס0�'��|C�}��q��9�S�J��+c����L/��EF���Z��u�Ge\OVt��e�d�����{r��pf&��[��]�_z#�����GP���^�C����/�^�5-���$x����f��(կ#>?JTlp�[jＸ�BG�j���5�S~�(GMҦEOs*�#N�?/ i4h�k�JώJ����.��CkX~ׄ��g
?rB������l3��P����X��~������r����,�/���Dejc}��k����Ǫ��W��4b�a���XG%��cg���u����:y������ED�s�O�����x0�T|h����t��O�FT�����Ϋ��g%�Q�cbņne\�9ݹcŰAi�Jݣ;��MF\�\�� �y�}��״��S�:�/���(J5l�]yC�g��0y����CdQ`�4��oM6@֯��N����Ǝ��d�Vg������=ʉ"�B�lv.�3���g!d`�u^,B��D�,>8G�׋M�a��]X��9�wc�2���,��־���Tl���l�D㫗\�`U�|�4E���,��uN�A��ុ6l��;�4Ef:3̈́F?rN�{h�<LCHߝ1S6i6h�鶨�b���g�U�г�3Dq�R�|�8��g�LU��b�kݭ8���l���=V�MN�a6�o�k�܈��v�{*�o\��[�5���,H���G���x��U�"�DԹ�5"$SCy3�qxf���{~��8��%�"����.?a�&
�hn�<,D$C� !�����u~>$�4||M�+�������;s�ޑG�s�v��#��E<��e�i�����C�{�Yb����c�|���`p����p�F���[Vx�=�	����\[��릴�iD��\�1�]d�w���)�z��1�f��L4t��CƉr�nL�Z�Q�ψ�DsC>hY�Zi��.9BxCp�q�f��!FVُ:�����J�K&ts���9�Ӯ�}�k-'��竷�z=��k:�P�t��j�IF��M�#���c�o�k,����q�\E�#*ݙ���k����������Ӣ4קE���r&r�{�kt��*I����"���T~��a���c���!�C8��~t�"a��QW������"a�o�� �c���#+PgϦ�|D8u�>H{��(�d:~��s��acHh�!�./HN��A�Y�Ao��]�=[<(""5���;��4��6�{U����di�C�Q��|x��N�ul3�]�)����X�ִ�{�U� ����ܝ�fγX�)������,��N�ǽ���9B����MP�l��(ąr�Å�������|	|�hh#��|Y��fx�[�g�S�xK[hiw��[�0�#�Y�ō?Tl��B7|�E��̈́E�́�?e�!���͋��O�m�<��fuP�����I�ut��d���Rf6|�����.�X��;?N�ǌ�#ؙl�htB��ސ�5g�����F�Ś?j_f7gn$v{��6��8z��-$�f���!V��/:�y�M�Ha�g׬)���L{�8E�����dL�~�=U��P�E.�t�9����'ܲ�-���63���Ү�s;j�G�ٔ�8n��諭�9w�^�q�Ƣ�H����ߜt�j�x���%��=H2(�!��/V"��z���.��W������DF��6��!㱳�/�Y�.}Ix飄<@\B�D����޼��`4e���⨇�j@w��f�M�z�JlK�t��t˾�E(�2"����F4�!�fCd`��z������.�Gj>&!�Y�Bε|��j�4���`Ć�GE:p���Ŧ�z���O������[���+���j�e%C�,KN�Ҽ��8 �99�o���NH>��[R))�%>�e�_�j\T���_}��o{�i�W��!�,��4h����S����4}�4ѣ��G������O��m�KMq�5�V ��*fO�����jf���u਌?Y�d0Ѽ#�r
�uu�v;�g>X��w�}�ih2(�~dJlsc<������{�i�>#�}��d���L���I�U�a$t�3�!�`�Z�.�`��M���v�1��Gi1&vfL���J��@!�p�����Q��z��"��!淐�4��*"�ϻ����y"��y���i'3_��PB(�=�����A�H(��ۭT�AX�}]��\��ڽ-i�~5�BP�A�6&�_@���+�{���j6�����,4I��j��6M�����б��f�a�{���OS��oo]X��.W��U�@濼lƾ�E����jc�]�p��2�gya�/�d2+��^�ʭ�څ��C�6����6Q'kg|G;��i�#�՟�Ɩ��B���(N�`�E!�:���6ln'�������b���U$oLf��%9�/�	�s��2k��@nq|0w��lU��aK8��7.�r�{)��8[;���Π��^�����f�>���� w*>��lY:99(���_}��{��B������.������/��S*y��8{�C@p׹�fr�R��f��c��FU��7¡�<��c������x8(���1hE���.�[=��b}O�h�?(��p��+Is�I���b�5}{��G�!c�.���5�D���	�����X���z������Ǥ���qWX�Y���K2�S2����U�a�q�Y-�-8�'��ͼ&�mE�ܽ����t��� u.kMM�gn�fA����;=|�n���8!�9039u�t�Q�"��Wkk[*�;�g4��X��5��9n�ttD��R�ݓ{,۸v�"�MfpK�צd��P��cp.ΈNb�6�od]��	|!��v֥Y����S!�.��k{u��ꣅ�� �w��)_c�p����X�vo��vѮ���Y9t1����b�NU*D���*-�&*�pӱP6��z۟�<3+o�{Fe.�3�r�en�:���K`w�y��|L��^<��<�5֚<�a�u˳I� W7V�R���b�8�g7PA�}�(0��ρ}��r[���,���GA�d���+�p�*p=ĤcY�v᭭��0:a0���BҺg-ƙ'.�#z�z��!�]�F<0����2�3B��s[��u��r!yB���F��
.�E:�5��F�VW��c��wgz�e�F*�\��eW�%�*��wҊn�h[;ON��<��xD��wXX{��9��u��,:�X�1GA�[���_>�ti�&�6j���Պ6��jX揱׬}u�u��¯6둮b�hƳr\J4������V�˙�ۈ��D!M Hia��b�8�e�31u������2��4��
�̫ZfX�1-5��`�iB�@��#�$�|J.@�)�e��.���Z�̦Z4���\q�E�V�"�Z��n��t�i�\�5���14CZYLcJe��-�L�s6nV�ƍrU�n��L֗l�Ѫ���."i�L|�* �$3�h������O:�������^���@�LS�����W�.m�_��ځ����|立��p��l��ʪ�Ѵ:�H�s���G>��f6:��b86��[T���1<���7��e*զ,�-K��MO]E�9��x���n��F��F��@��92,&��+�B%7XV�V`q�s�~B3�h���޺#d�9K��د-���j6�LOz���,��r������pOp���W�KV�XmX*���3�ZY�����2әΛ?�;��b�������-�O�k�5Qy�풙�*SIE�ilތ�j�ĜU���_�E�8��b��TZf��'�!���s{��=M��ql�ר���>V-�{����n��^v;y�b7Eb1F;J��� ��v2��J���B�����	�R�� ��'���q��4�g/�+��閍3��
S�+��P���kGGA�kV{��)���{����骴�T�գ:�
��X�ol�#�m3��˪�6����=Tb�J�~u����	�ܠ���>�+�k�%�9�|񁏻zv�"���ڎ��܋��֙�/v�����n���G^c��ю:�B��{�9���A1e��B�P�,d�wAU���U�]
4���5Kj��U{�!�`ɴ{��N;+��N����]���AT�-�y:r�!)�>Nӽ���/1kٖ�>�O��X��+�]db9p}W�P5�}~��(+#��Qv8gc|i��y��W������!���~3w��'��a����_it�_�4}�c���~���c.@i����o~X�ܟD>.5~��o .�
gu�����Ԭ ��s�{����ա��%��B��W��&xiJ�W.۾;f�j��qT";�v�<N>GMn�������6��[��2�_WI�&?~���[]���W`�_������u&���A�ܰ�gv���WL�W����Pq?M 8��Xae�#5�B�:Z	vz���k�kO���7<���>إ΀˩�pX��;�#�<'���Z��u��H	��h������q�M�ܝr�v���ՐY����$&x��\�핃qg�.5������f����{܃àB���u�pT��=�-���K��7���ÈeeOb�[��T�Ip��IUi���7�.�PT`=@���w���V�F�#+��\9%�{�u����=Is�L�+|�'���Î|.q���f5`Y{�4�k��Cz��F��}�6"ܓ8�X�'����7=��厂��inD��n�{�TZ�'�]I3P��7R����A'W��Ķv�`����3�R�>Yg��hl&�l��D���	ϒ�J���ۑJ�Ϋ�ˏz-jQ�;��v�
t������#4�3�W�2��f�������̑xY��|��Ug���7S�x��{��b��6�4ˋ��A�����5����eHS����\"��]�3T�Q���u,�Xg�v�~�ԣ}jC�^���q�:����Io-�p�Vf�ѷ"_݃z��#������n@�h��#J�FĞ�9��0`\d��jf����1[V�|������+��h�ވ�%s1寲�w�I��{��I*��Q��c�_`��ܔ�.��f�q�W!�c�e���GV�w�՛�����Ѐ=�P�����^r=#�� �Q�����-0�&U���mNu�:n���g^����o�z�e��5�C���t|�7�}�E�|���6�җ�.U���U��U��6Y�n�N��K�f>�%λ�^aNs���9_�d�_.J�����I60��fC��O߼M�/,KΥQ=��bH��^0�;X�r�¨s�0�n��Bd��ͅ�
Zs�WN�ޔ=��n��N���9�A2m�6x���Ӷ�f{$Qb��]E�N��fׁހ���8�<��nիFbzsq�k=٠�u_+᎜�� ��35g�����O��������p��f���8�x-J:q�X����6!X��WVg6;77�.Nr׼��U_wO{����b�5F�>#`�����WU���y
�`�Kn?gl�pXn�z�5���J>4�e��˭�xi�Z~n-�&��q׍�nf�'{�-e?l���	W�WwWz�46F�Cނ���5p*8T��>g��OMd��U�
{�ۉj�:�Z�p�+t��L�Ua��������켶�מ�'q��{��@�;{�oAޗj��W=rƭQ��qfȠ���^���١�$pj�����'x���t7��"�S��	��ꐕ�w:C��#U\�{�_��WJ�g+����QN�ɗ�	���rt�%Yr����w]{�DB�Jv%���QK=v��YT��en���b������{�)%c%��/�`��ڨ�2\��-^ˤu���/�gt֬�[} 7������ݹ���'+ת 0���
"�9������I�1�|7�$�L���a�Tj��vK�E�;ſ���Q7�e�U�mht�K��`r���q�WT	������D�;�h+�4�1��'ZX �Rk��&��	XhK7%Ee�J�aT�S����,r�p9���P0�[R\�ʧQa�EUn�۸Hwj*�]Y���J�B�E|O�:��S�Y �⺆��yuXĺ6��!ȕ*�A������l���+d���ݬhkς�ta6�x�3yXh+?;�D�5W0�(�9�35)ը���A�<�m���$AVp�����1]o��6�ޓ�z<�fT�k��rU3EEJ�+k[�h*�2c1�����*�����l����̣l�kmW��f`ک��r�ۣ�X։Y��8����[s!�E֘��cG*�ə�4(��-Q����r�ͳh������s3"��X�J��(1b�.f)�Pb�*8帰EUm��Q�\�"ԬT�AUSYU�ks0R��1�Q1�dX�������]Ys�S�;:L9ہ��KVs)��؄(�:K�����.�wZ�8w���4�:�0(B2�{m���M��̹�NQ��ȱ��ŹP��q�p�+��*{��ؑ{Z�y��s���*�^Ԭ�$ߒ��ȭ����L�;@�푵�����X�Wj�K�n�<���y����]w3�S~#�&W�Dfi,ov�(�P���rRq�l�~r��G�Jo��B�e��w֮xѶj�iG���3;�pA�;�z;xxW�w~�ӏ��<wrDa����8�y5j�Ʀ��F�=�<�̠ v�V]�.I.^�1�l�ta���Z�n�pz��0*��x�����/E��Ӓc'­�i/�	��^S�~R�m��]�I�Ngf=@��X s�}�xە1j���{k:�g.Ŵe�ԕ��#WfaA�g`W�Uv��W�_w���uֳ<-uվ�wH�[���]�wtdkC�wP)�mZ���K�b߽�G�6�g�!u�M����6�����H�u�&�:��R��S�RB8n���ٔ��bR��N��+�^�d�-�l��r���c E����7����[�f�3*���B<�#����ܮ!王�^����q�VP5�]��=���
+&��z��ȧ}�Lj�pڮ�=��U�R��qp�+Y�݌���،]u�n��unXޮ��1�>�[;��s���I|���O�W��'�6~�58!�;�psL<���2O/&w�7�^�Wv����u�<�Ck�n�KdR�8\��@��dX�n�u.��^Lj��={����.� Q+��	���u���`��[i>��0���ڼ�S�������9zy��UF��:n� ���7�v�
�|�����Ku�
�9%����-�`1AC ���pT�7pbM�R��`��DDDG4�IK���9r��T�N/x�x_�F%y�4־�[�k����}ѿo�"��Rhx�6��+��ͽ���"�E2�����>J5�Ԥ��!���q�om��@&�0��<�u/^>�X~X��Ш�o��*�	��<<�0V�z����/j��q���R�k���6���ٷ����u��v�bx�uB�d��I-�1O���\,�"��U}�}<�s����
Aȅw`�N.ѣ�m}P��Xˇ���(o{�w�{�B&������L�yַ�=ST&j��������1��{��tK�hz*A�"���#$v���]Oh��y��<�'��U�6Z1{��5Yy2�6��(u��fWY�����xe*��\����d��c��s�\q�mn��7I�UAٱ���2�s���<��	�Z2���L���ԵC�S/������B7x��z��7W���[S�� #�&h���y;���������J#BN��z����[�f����+��֌5�<��$Ow*Ȭ��.�L(v��ws��dC�����������<(�8���4tدJ�
���"�m���[Z1�Oz��k}^������AK}��B��;�ޙ�fts�*q��݋�]�7t_{й���ߢ���ܵ�̻P�gw�d�s��#�ӷ���xn�}X��I<�9v��n$��4��:�r}W�V"��p�Љ�-�ͱ�ѹ����_?r�EAٳh���1�bZY��ug\�ze�=���y����L��S�0}���z�;wvzjJ��c��5N�M����$_oZ��.�1Žm�ts�.=]ݧ���'��l`����R.�u�]��s���1�~��8H�����U��sMq ����#<��Iju�0_��� ϸ�}��>�
5�ͺ�����a**н��of�����E������-?sg���7��]�(y�ؖ��{_s��obxb��L�W׻��^ڤ�ǔ.�5zMn�uv7�z�����ɘ.��Gԅg����K�ʬ D׬'��V������q�	�o@�FY]6��m ���(Rc��Mqs������g.;��n'�fTEKFν��3I�Ź�K9A�^�&�Ag`>��k��G#�u�I�#BL}-�/M��'������:ݣ.�r�����¡�_bԸvp^ۻ��u���_��v��S+�k��R���r�kr�Y���#)3OyN�5�V�o�
S���k�-��Q�Q��Z��V�z_m��p�Q�޽PW�e3}��,̏��ꤴ(�m��@o�&4��)�w�m�/	]�m!�
g#z2���J�q�]KK���7�Q��q ,��^��\^���mf�]tL�������2��>�����:���7t�t��v^B]ʻ����Jo-���Y���|2;�"=pW��_1�e����]&ձn�3�Й���R�u���x��!��3���#,*�y��':��Q�e�bW!�oN/i��Z��n��V�;��{�M&��^�)n�v�崊���F[b���㲐�����Yl�/����R�e�[��D��l�?5w�/$�J�|��&5�^4���w�e���!0fA���TnrFmӘ��&V}X�����:e����)+UN\�����a��83wwJQ�3"ˣ��
eI/
WR���r�6��t
V𪆑��$�peTX�����i<���fb44�&GF����F��+#F�V���2^-�
�ݒ
Øً!T!�����QY��U�ڛ�U]B�D�"�
�""*�EX�J��+��@b������X�*�#Z����a��*�UV;K�%m��u.fa�Q�M@����C-�\��C1�`bJ���(�j���T�*�R�+Qu̲(�
[L��PI���S�(cPX6���Z�YtW�WU��b�]ʓ�|�'6�	]�ؓGV!�7�%-�'9�<t�0�v�z}�ÉŚ�	����g^���.{aRWV�n;�_+��#�U��$Ć��ͭ�9����H�fy$Nva~O��C7����1��T��{Z�����{��r����z��Ҟ�}�W��ͨ�[q�� ��	yݴv�&31�/bhI=��~��m��G��-�֎{���^���Ω۝F*�h�Ѡ5�)�wck�\�eS�(n�Cw��:g=O���F�p+mLQ�	�X�FO&�*�û�����`���?l��|/0�:�!b��C�oݽ��6n$��v�C����F��m8\�VaB���|���}�{��L��k)!2lu�/v��iOcKws:��c0�Jf�3���"p�bh%�\m�S����ǂ�B�Z�֭��N��w�74kTl.ݬZN�����yKRU���o��2�v��y;�q2�'�mz�^V��wZ�e�Vߖ�l�oq�֘�N�\ګf	=��qVᵦ��]\��<���Z�CM�LLK�����X�|��zn����>"5<\�dS��U�W9qI� �ߦ�Ko}.z���F1�M�����g%X�ל��J�7;�}O}2����i�p��r����S���Jh�޳C�l���I�E���i��Н�W�Luv��ך�$�IC��e��
��f�w��;�Vٜ*��F[գ�9�7�3(!��½r..G���}��<8���j��*hb���/M����2h���;9�\��.����9��
�l�X�������kN��@�z4rvJ̅��+�K��e]�Y�z�n��.7�f��I�6`���:�b�����|��Z�I��I
4�_w��>oV��M���4�;���5 Ʌ��ZKN���ƃ�g^)ص��1�$>���[!@��F}�[݅v&��n�.�H��Z�r���>qt�?P���6���f9������Gi�C�R�$�^����Vpq��EV�ޭ��v��U}�+6I�e�g4���ScFM�3 ��� �ǅ���lio�[x�0V��qb�Ty?
�y����b�� �u��9�zqC7{zN���MΓ��seL���s�XOw>刽�Z#-L�Ű�on2m�(u�V��sk	�3�z�GnN�>����1�M�')��2l�腱N�7�d�y��i�j�5����q��1s�����Dxo���7,���/��'�}�$���U�V5v��3b�۾	�W��c���ݼ�/��G�6�^�e�$�]3Z�o��rxҥA�w�'@g;UC�� 0�w7�$�G7�vp�����[�N7_N�u}.ub简����f*v�p�i�}=9�0�u�2;YOvU���H��ˉ����h�WfϞ��*��U���:�u���wj��G��μܶ�Wcn,;==%aȢ���y� s�shY�0<��A�N�pc��=��9����o�$C���CJ�k�k�ձ.��uf��N��5.��Z�*�v��voj�5�`ݗ��F�V�+!�S�M�$��n��s�.� �������4���pL��G�_�u��K���˥p؏����xh�k������4�S����,ܗ�IE�b�`�(7��W�a��*{78����eAf�1x��OZ��݇~������N۔�򚽵�½r.��=��\���z���f���#q;��x*XY"��������e���zRԗ/�L���~�j
!<+֯�Y�(͇��ed�㳓���W���%a�q���ůTl�z��^*>�j��O��b8�,ه�X��8<�k
�h�e{r63|�7w��tk�fd�`zZ�5����z�w�۝̹�`%�=Hǝ�t:�T��lV��5-@dlmxRoXF���Zh����8�׷�f�����W�g�&ȸul"�àli��[�[8i��� �K�9U�R�|ni��${�H�}N&:N�Z�%�P���<��N<�a9�-�mc�o�HR�mM�U�o,fsw�uc*�b�pޛ����1�\���yٳcz�N�1t];�d�	�O͚������ώ��{����|*c�mx,�n׌�O���)��^A�o'���X=XS��4���xy�c9�e,����˽��Ԫ+6ar��}[��5f�YWL������4N���1�t4\��|'?�og�o���re�b��Nw�U��U,=��`��_ù�x��
uۣҹ�8^�x�O|�Ƶ()�����r�H�{���3�o<3#�WN��N0�R/�\�<�m\�w� �T�N]��d�G�(dW�n�%�(',�z�!hwaM�D9W�c(�A�ƴ�����=��cH��)�;dGK't�������=�:�h&��:?YuyG�u�ӽ'v�����I�U���V��&��F�MeW��O�%#t!�@F�3p�)� ��Р�ĚL'-��Pె�YR�C2�Z���8-�X;Ec&�[�����TK"��m}�)ݑA��7�:x+L7L�qY��)<�
�IJ pV,��9x(��7&<�D�w�[B����v�d�K2�.���nÐ9x�R��v)��P�xn�Xjh����5X�7���j�Y�3u7+�
��� �Q�-�lU�l�Wl��\�R(�r�@\pLb�Sib*"�*�ͺ�dUQ����Y���P��J
��`���
*��`��ҡ���,�QAL�)+���qDmJ��u�Ak+QTTE2�,Y�L�+1�����30�s)�Y��y﮽|�s���}�<��Z�]�J�s��s���r8�Gx��Vj�3Mr/�����%a�b�!,���T��i�-u�@>���ߖ�S�U兓��}�D�T��ed�T���:y�ꋐ�ix�|�{6i�YY;U\�~&1�\)�L�Ng�b�SIܭKǘ��J�v�a�ڽ���'K��N�Ͱm^\��[Po^��{
���=v�ݜ��SC��i��{­q��y���2M�w4�ef�@���{�bGؔ:5����Fӗ����T���/^��7�a�uY;��;�����E��ɔ�Ŋ�l���̠��j9ؽ=^,a�C��}���OO{��\�Zw�eff��:�>�E�FB{Q��5,)�ME!\�Ka�]Z')Ɠrz�ۻ�}-p���uB�y�k�����)d&9�ۛ�;�#w�!��I�W(�=�jK���7���U�ԕ�u�(��5�J?�d3�3^<��>�jF�|�"L��M�A����-�Y���c1-�,{�w0,�}�^����> _u���s���է�M�I�@;T�nS��glõ~ ��Ul���5V`�n��E�cg��#�s�.Q�n���}q�K��_9의L��ʳ|����r������I�s�M�
A�}�Db��+ �=��z�by%
/�l�p@���w��ˣ�����~�'�`k*���P!�: %�b�\��V�Y4ɺ���%NNz���@oq����-^�\f.V�9����K-nv�V�����7�9U~�[�	�G�M�S��e�P���%������%��]`��S��х�S�n 9sÄ�,���ܽ}�Y٘�v	oe�Q�]��V��zk��&N6\�]j�t�<N����u+Pvd�J���[j�"٘�}˻w��wV��ϭ���u1��7���Җ:മ5)�U��˛���9=q�W�T���82l��鸲�>o1ICI�K蜐��"�y�+�wk�`�5|[���uh�6o�-�l�h��v3Q�[G����,ڱ���_�vw�~��.θ��BaG����(ʾ�:y�;쥴���VS���u7�����*�i"������^W�@�����IK�����&u���ۨ�-��v v�VwC4�.��i�����qu�;wu��*�).�+���n��n�-������wZ��ՙ����eZ#3�A�[����6�n}GU��N�!��e����<�n�$7��K>#eN;YA����V{��ξ��~5�����>�w���8�p�:T����������qr��<�x����h�Ș�����c/��k�C��1�ϳ�M��rv���Sz��۔���hy�틄Ʃ���{���u^>鮻e�n�O��o���Tv�����aol�,.�1���;:[8�^���V��)��I|7���LU��V6%�c�o}��+����5at�%"�Vc�
�4{��)z�B�s�V���92�.�\�!�s����e���Y�I�J{�0��!L�C�x�u˙�wc�q!��]��ݛ�nwt�$�v; cч�5QSk�'��ܤ���kX�06�ǊcM��<�ьeF��N��$q�ƑŶR�F�j�2{�B+n
s�g3x2��-�$�m��{��izB�*hAؙ[93y�
M�g׵�v����z��\�Kܖ�.8V��%�����Z;Xb�&D�"�W�)i��\U{�$����e�cl�J嗯��}i���KzI�v���V���Z�d~V�#�oM���ߒ*v��+�cp��yDc8	�<Bʹl�/�r�<4�V�K� [���6kj="��#<y�O�=}��nz3�q�l~ݤ��ݜ\�}^�!�s|�8X�����J���N�;�=U�ut�;'�C#��V��c�_nD���Q髁�ol�o ��!���[��S�Ǚ�@�m_��!�%���ݻwG������j������m�Ŵ=�&#�	��=3�^���b��s�=�3q)^����>Z�����:�j�j�a�EY��+�����c��J5�b���N���ƣO����T��==zhc��h�M��έ�w("���s�_;���S��V2:�Lޜ��;:����HB�����Tԩ�����g¸0�[�
wi��	U&fż��TUasʥj�Fju�L	
�F��oz�0B[�[D�4/S�0��c����G�f�a��M�U���P��u�;ǛF�l:���u���*���F���Q43$��;Τ���"��i�ȋ�y���}��CǪ橅���)^k8'p�s�U������W�블]&�hh�Fq�n3�e���g��Y��b���U�idN�<��oo=��AhS�k�q����<�;]4���V&ͽ�*ɾ7�P�8v��C":�6�	� g^`=w�bp�x�M �:�ݮ\D6�m1�r�x[C1��E��=�2��fW)5W�#;��b�d���+Y�r���ˬ�WϞta��;:��!�W]vvv�׻5��0�ʝwtWHr�9g
�{��2�Ӝ-�]�"8;������3Tg�K�:���s��yf۸��H%b���p�o.	�*&�������}è���9�y�*U]%�YbW@�}�G��ɖk�ۤe�[��+p�2��N,����&�D�����X�US���"��Z���LG)��*��ed(����*T�H�cnZ��AH�+PQQ�W�*�F�e,�I�l��F0�(��E��8�b�k(�Z
b�H�H�*T�ҥ-���z���`��~6�X�)��ܰ����J-O��������2�����fߠ̍�A�U�&�b����C��P�����}���q�6���=��7�߫S�ڙ��bd���`zt�f{�mz���:/xV�՝v�)^s.���He�
������l�웳���ܧ�sp����)�yt���h_h޴;ܸn���>��׉��3@�z7c0�c��.s�q޴Iٜ��so���}�G>Q*��R�&"�l�B��4N�X�LeRk���qu�{A���p��'d��jJ���SSo���M��E�p�w����W^f�%��#� �̧�]�	���{<���x�y��Y��7Fyc�=��x�"� ��ͥ����׫���Ae���F��w���o����%,Bg�'S�s޲�s�u�%y}��v�����n���A�fK�Х,��l|{�n�R�9I	�ܢ]��r��o�c��<�VV��{���]��[N����I
���"����r�� �㈱�-Z�@�����`��t�u!�q�n�ˮ�t�Е�C·qY`���Y��^g��f#)��]p>e��r��}�.�ۮ�|�bB��!S��h�U��LAx�!��H.]��қ�R�Г����?�~{|�l��g-ͽ�f.��㧝7���o��_9H%�>c��\���0"ci�p��%��^�ifC�&��"����f���H��W<�늝[ģwawhN�wjtX��T�2�a���d�h�y�m¯��-��S��v^�!C�ezF�Ȇ%��tB����9�R�,�uZ�Of}-+}�����3�U��{��}��䅙��5+����fI�q{>�jG]9� �uf-j���qi�B�E@�u;�YӨ�w���WQbZ*$�3`���J���o.:�ba�" 8�x�AA_��qǹ��zǙ�^��ckvt]��{D��.�.�����ӏ"��y��gGm��pe��
p���|�OlA�]���bIc::%ޞ�V殞<��z��o]U�+�ϩ���u�z��9�Vw5(�oT�cFiarހ�2��!&|��1��%\��N�-�oQ��&��k�����{�e/��;$؟D���v���۪����=Yt��d�n��;��u՜�qh�@Kꅝ<#��u:��B'��k@�GG6;n����l�-^���iꕂ�f��6�0,d:�SW��wOKULP���ݔ���z�MU�ʩ��
�-���É�y��6�{�i���^z��Ad��m�w���0�y��{/��}�^7{�	r�e�^d�`��]��;v�l���n�����E�O�����}���\��������U"����h�+&���ܳ{-ܬ��hЄ��ק���t�aت<��/g.��lwC�������ע-���u����I��/�v�r�}���N@{f���7�ƮZs��5cu����cS�WL1��Ur�A.L/$;{Ǐqr������3j	A73�s�O�g.��M@4�gh������F�W�iź��e�8���ڲ9��-�S��2�-򫖣�mB�6cn����ui�]��ML��� �#.����Bh��#.��]K���9|:M�R\q��yy��0j�F[=7٨�;Œ��?v�u$َ_qQ`f�<M�h���n:R-��;�!;��G�1��^2w٩RU����';`�ĀP6v�姊�O<XZ[%m�ҹr��)����s]�s��.�S~���^���J��bܡ�A��(�v�Uv�S82��o�0]�1Ρa�Իu��}��{2O]����>o�%�Ňgkq����9��{qr�Yz����/��=�f˵��nG��كA+��a��3l��m�8��W�({C~[2��
��޹�;��M�U��<�$Y�A�SY�֧��ct��fF��w��Au3���"黠�*�{�ܛ�������YP"�__fi��^�24���!g���S��xp�]zq�Ȭ��:�{�*\�j�2�`D��sC�_\��{~�Z�sj�6o%�Z��w�^z���BUoe,��ײ@�	�n���7�B'#ѻ�c�w�/�tS��X��CH����^��~��'���XT�ԭEUW���DT�I��(���2�(��m?�����B�e��;)��������&��n�BT$��Q��$���wg�҂SS!�����?����t�P���=��)����#8K������U���I�){�!�4,��눡���:��<�P��a�>|��_����}��}on�AEO�t{Otݿ�x$��QS䐶 TT�Sp�	+C���tM���C����'�M0���>�B��0�!q�TT�����\�" �4�0Z*W�B�c%����*1��ɭ!Y��rL���@W^Ӥ'~ΉNws�vX �ә��آ���cX�	v4�w4�TPQS�C����]5(Ms��	�;|�^J�y��#�PQSKd-;�t]�v�K���ڍ�!���3��2�L� ��A��,�_��x[��O �U+�ˢX�ԙۈ�ǰ5}�X�Ol��h�@��_)�Ùn���DTvT?��Nt҇B�<��P^k9�
*jx����_MG����$�,=�<%sTT�E�PQS�������,Į�vh�y�R@r*�!c�
���ƪDD����B5�G��s��U������?1��8?�{�9Z�zb�
��Z�w4��Lo+R�(���ELZ^���]��PQR.�9	�R5=����{�ᑣa���ڟ�P� ��4�,|�@P��7����!<�C�kJ|6�/K�y"���GGeu�#`�Gx̒!���;E%|���������̏�9��C��ûѠmT���Cä�A% �q�y��^}�b�01 =�؏O��:a\��:�
*r����$�v�g<n,�w^A��b�5�d���nB�	��y&�RE?� <��X���{|�M��f
(��v�GZBX.�d߾F�Z�`���+}:Q�JT��A���J��iG-���rE8P��h�