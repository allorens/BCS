BZh91AY&SY�|�ߔpyc����߰����  aU�       J(P   �    �  ��               �    �|�ڍ	T*E% ��|	�	= �J

PEI@(^����m�����ϳ�����uz��_A���>A�{������6׬��  Aǂ�]���@Wv;a�׼������v2g�C���ݷcJ��ٞ�(�������m�@   ��   �������>�zϛv=zz�����;g�9w�{��{8�S��  8ҷ ��s��<|����b��(�����F�v��� p :� �6R��=�l(}uԃ܏��z��ѐ��9۶R�r���2z�`�� ��{�*:���pz��g�����c��ք��!��� � ���������@�-/a�c�<^<�{��F�wl�{���  �p�1�����|pm��6Hh��^��v��h=� ` t P��7�ǁ� ���a�{]�F�F���={(:�w��Ҟ�� p�g:2�z�qN��Cl�ɐ�#���`�g�|q'��<P                       (P �  �US���J�I���&�� M��!)*�ё�	�CFCFL �d�D�*�!�(�     & ���J��b10 F`�   T�$ �MO���MOj6��a�==)�x�!5)SJ��@  �  ��X�G9��V�ۘ���g������yy<o��f÷�s�G��}���&����l>L���3��8��������z��������ӏ��y�#���X֥�������'��.q�R�{7��1�a�l�Ɔy�:ʪ���?�����c��1�v�П�?���x����t��~���o���ϳ��,��i<L�c	4�&3��I��q��<�'Ro�Iǩ�ē�<I=_a�&����x�<�I/�8����$�"��I0��$�'>ē�Lx�v1�L�_bI&�ĒL.bG�/18�_�m&�I>/�I��1<I��g�%co?z�[ěx�,c)�IƷ���/�$�M��$�+8�e�ǘ�Isz��z�I��I0��I$��<I-bH�0ēԟ&�I9������'�,��m=_��)�'�Zz�~��F$�Lm&�����I�LN=L�X�-��g�XI'���|�L�<z�&���L��&�I9'��ߞ�e��qē;e�ȓo?M&RN>����"L$�/Ӎ$��q���&������6��K��稓S��|��'���$�I8ԛ|��I�Mfy'�>OS�$��	<y$�$��'�>|�Ęo��&Y_��8�ra��Od�a���_&p����q��������$�ƾ�i'��V0��D��8�I�'�'�I�L~����ēV6�'�1�I�I�I<�'|�[Ɯx�/�I&e�<a'�>�$�+��$�I��i<I��I�ɋ�y$�|��׏RO��d�0��I=�$��I獤�o䓌�ƙ�'̯�O�fI>y$�5�Og$�ͤ�$����Nm'�/�z�K�I>��/x�I���?I�i<�H��'�ROs�2�i$���=I0�y���Iq�ǘI/����Y�$�&䞤�>�$�Za$��I6���2ܞ$�؟'�$��$�a$�/�I%�~�|��$��I&�ē��i1��3$�8��1$�I�I��I8�L~���I%�I>�N~�x�O�$�N1$��bIe잤��	��bI%�p�	&��ل�14x̛�L��;�^oh���x�xPĠQ�~߰��� ���>�q�b8���cIx�I��$�q�o1�ԓ��O��RM��I�Ӊ%�I&Y_�O��[�񴗸�I�ǉ%�m8�2���I-c�>K�I�I~���{$�cI'��\��|���$�e~�O�O�I$���1<I/q���q�L��1&_%�I�Iom�ؒI�I>���8�m5�6�ė1&_$���|ǧ�ǯq��E6�F�zߎm�:Y�6{��o��1$��>x����K�bz�����Ս�_0�y��/�<N&���O���<Q�v�<��J�O1'�c}2�؟5'2�x��k�a/�$�����I-�Ot��O�q$�i��%�8��%��~���v5´���od<A�;��XÇ���x��&ZZm�m���Ox���a�z�k$�e��^4�֖q<qoN'��m3�4�Mo���6��I>Z�i��$���p�\<���x�]vYg��*�<I.bq��bI��$L���a}�%�q8�~��<I3cO^����m����<s�I4��&#I{�I&�q$��e%�I+<K�I=\ư����q�ϛ��O?I&���X�����I/�N'cX�|�s�I�K��h�sX�I��I$��Ē}�$�m��~�|�ROR��I$��4�e��I$͍�I�L}���k�$�M�=I9�&K��뮺�]u�Ϭa�Y2�{�'��V8�6����X�q<"�'#��$�K��_bI&�a$��'�/1$��$�'�I<e~�$��ƒL�q$�M���I/q$�%�m$��$�%�I$��$�ĒMX�I-�OR^bI&�1=z����RO�_����ŜI&\_c�RO�<I/q&�q�K�I=I<�ǉ'�o8��6��m$��$��/X�$�I�OO>ĒM9c<I<�2���N=I��I�I�bO�x�$�	���0�z��ox�m��%�$������_,����'��1�^/��KX�%ci�k�N$�����x������^�".ba���ĚXĜI{��z�}����z��&�\V=XǭX��IoO_/�I$��0����i5����{�I$���I�I�cԟ6�^���I�16�ek�0�>HL����>xh��9��9��/EYҬ��4�p��7g�r8�٥�Xc��^<��>|��,�14�L�2������c�ni��ceo��~�^�i<ra<m��'�������|����%�~���s��N8ǏZq2�6�����q�y&�y8�m�s���2bI���$�z�a�����'����z��p���#Kx�<O���Y|�H��"q��I=�x���$��+��/[�4�=XĒ�&ޗ�%�e$��2������\��������%�O�h��Ĝ�zKx���|�\��g���ަ^�cI8��8��ߤ�q7�L��$�bIsƜL<��LgI�a�o�/Kx�'��1����4�z�e�I�ؓi<j��x�e1$�/�Ğ��'�Ĝ|���I��z��G�1�$�i�$�s�Si/��_�[I3��I�/�a$�iX�11$�L+��Ğ�$���$��'�&�I�I6��O^$��$��x��<I2�4�OI~�I��&Kl$�a9��z�M��=I���=�I=e��$�Zğ8�O�x���I��&�y�$�$��$�Z�Rz�_��m&W�'�$��c��'d�M'�I&��?I&RjI�O�5���i�޼I6̞���4�|��m�q/L���&�ѴO1�be'�M�\�=z�O_O�$��I�}=��9D�nL���6�h�rmm�M<c�$�:z�5�a'�6��zω�?I��m<|�z��}��<�Nm*,�GW�:n�p�ߛ�ʱ�R�g������o��N6�̶��f��}���!G����]8jo���x�Cl�TD<Q<S<fx��S�|g���|���}>e���i14��&\�e�1��>_�Ĝri��ce~�$�~�i}�>K4�bO��$�S	�oX��ϗ��}����`��.cƎe<�lm�YI������I�ǩ6���=q9���߸�LI<}�ԙOU�~�_��O��&le����1�ͯ�b6��c��z��ϗ�RK��|�?�c�y�'�^2�1$�X�,�jƞ�K8�is�_~�	kO�XÉ���L��1���6�y�+�O�j��'���XKx��3�2�r������x�/�$ۛ���<}�Ikq��Iy�&1���^`���8��	�&����\�O��M>{c3�M"N-��O�ĉ&Z��	&d�}�����O���e�b}�����o̕��<�Y������;#���&��^76��a���}���; ���Uw�iW��7��w
~`{�ō�!sݸ73����;�}��M�D����(�ixy�:��H�OSdU�E�J�����7�P�D����>�:��Y.D�u���d���of5k��b��
����3���ۃ�U��;2�v��I�����u�sna�i�At���NFt����w��.��|��xw���,$=�ճ~�X���շ�H�%M�n
��tl����&��==����$:T����ei��@�`ț�?`��4��Ѻ������|fW���(��jfr[���쫗aIeA%��n�0jU���c��]Y�֓G�TV�G����<���׼������,㵓VC�fgl3��p�|����Y���O.[���\�����?!��#U~�?kӱ�̼� -+�J�a'�g�kǪ�g�ґy�~�����s��T]�߷�������o�q��)ۗ��/���۔��c�]os&�9CJ ft笣����G+e3Kŕ�4��n�<���Y�g�O��*�}�U5w߭T�/����~~u�ѢI	{��w��ʌH*?,,�W����U�)�?n���]���#~�~�o�������GJ�08d�
��b^!�����.���q��M{J��df��F~m[�,q���c�Ui'�$�m�R�JzJ���{��gJ:p�J$<�^g��W��^Z���y��
�#񧊴`��q��o�0��Y�W<<z�^'��K��y��k��oƔQ%���M�/u��j���8�:�Yj�gqOE1�\��gʻlp��f��N~{e�㹇��$'�N�?|�-��b�J<q��X�:Y'�2���7���(�uƇ䧙9����ۣ��.̙YN[ć
O:̪52{36���N��O�b7�9��nN�˻���o���>h�op�d�ׯX5x�	�\~�j��s���\T�q�{�܈ {2g6X��Sq��3/־4�#���}�ᝁ�=���z3:Vz�.�K�x��~0׃�켷���ǥ`Mn�N^��疢}C;���עv��̭��~�xV����0{<{���yz�pBN9����ב�f����ou}N���<t�'�(�4����r���qA��7
�{�Vy���'�|'�wW�NۂC��OQ^���kOΰ����	��_�x�zǂ�B��#^��x����{X� Z׏X����t��l��^~'�;�i�I�	/�N_��z�ՙ��L�n<��p+�d~;gS���y=��%ki�80�4|�z���ӍЊ��<p����\�/�Orf9�c�	d��91��_ADn3r4N�oj�s�5}*����$�W��2�?��9�?O��Yj����H�?���%�������t�z�Ņ�2ߡ��(�����f/�^8G�����߃��fճ�q���qַ�M>$�&�l�F[���V��2O\�?����s��%�7ޣ����~���e�Ϛ�vC�&i��YƶdB�D�[�)|�~�7��޵�\��V��۳s�'�����ֹc!x�D�$ӧc�~����D��t�')_>\lvQ�/`z����⛟\Q�`펨����¨8�ק��*�$=���>q�C�d2�#�Z�k��OŴPX�_9��P���GBY n�seϘZ�|q����r�Wل�;9>h������fe:�<�,��j�ë*{��v_.j\g����C�|�!�ɫӞ�y差��q�*$��_^�T�ٞƷ��}��<����e(�T��X�,��\�H"��v�א~E=4�S:W��j0��2k{Gv3�2��t��}a^C��E���H�s*`���`�>��|��\6^��(�N�[�)u�۾m�L(�:��k���#ٷ�o!K�Kuk�%ve��}�~�i`��J�"��<�<޸�#ݬ���E.u�����D�y���/�m˰L��HZJ/�f a/�M�b̥��1���#X�1D]C�RaES�<|�&���{��w��[=Q��E���eAY3-�����!9�*(�4���ه�Ǥݵ֍�h)f�)s=v��w=}��,�¶�rדD}���81x�Ru{�>G���^�rе�g�tU��L�A�agM+J�aD��!ggʥ0�L*����$4�3���l���)`x4��#քѳۭZu�whM���������G'r����Z�v�̗��(D�wL������NH���r�n6S��(�O8�<�����'X�������&�{�����w4�*�Yy��FOcWXC�^�a�-f0I����$E	Q�%�Y#-PQ�CM;|@�L��q?�WU	V6���,!��#/kxGΘ�!/�Ϸه��FI%�B�j��0���r?|�S���d��b2�)������ɡ���;�|��<�i{�V�{�}كUg��z���1�������~'V��KHao�S������&���D֯�h��܄%�YIm}���aXM���΅]q����$��[^�We>���do7�s����������n?�z�{}��W���7��ϕ~�NX�]�F:�nZ+�G��n�/9οḣz�L������!� y2W�ln��	���c3h���N�F��}�4���� l��7Y&��p��7O!�[w��É�����x��t�f~F'�i$���짳a��O�g8��S����D7���9
E��&Y��Q0�=i���j��G�LF��Y1੓p�E����&�˗s�n�<���g/^��d�g���N鹝Ib�˗%I�]�l���t���8i��a<¼���7��B�%�OԲg^h�3����nx�n�9+�\0�]�'�*�ş�=���,1�M)W�+Gc�i�Fd|Q,gO��HZY��I)Xj�c�%�c�a�+ ���x��*���+*�ܗNrsU�*���w4�Άc�O}�O�f9[;��Y�hD!�����o��x��ld���Ǐ�a��6ҎG\���ov��f'�^�<]���Og���G,�}��=W2>��p�t{��ٶd���q�D�0�p��n:�ծ�ւDnΕ�/�7�U��r	ĵ�FN_>ɼ�0�o�B�s�U��ێ[�'w[�Pw~v���������U��V�t�����x���M~��'��2a�Jy�q�����s��G�)��:v}�s�Ð#Ԉ�_�R9�n��,#]Q3=s~7w/�����c9��q
�ʊ�3�,<񁨯y��Rx��(��xi��x�R?p��Y6{_cm��>���i���N�;�CE���z��Wu�Z��振�����f5�0���,ތ��f���5�}��Ï�w��I�yYT����m����$�m<^�w[{�_�җ� NB>Y'�k������I��7��pɥF-�+7<m7c	!���`��4��Y����	͘ݔt�t��eCb%������,�k�ch(�ڴd6��"��i˘�fk�6�e�{�ZCI7{lt��N����Rj��������|��OYQX�+ ����}�4�4ޝH��K"
��r�	gRoʠ��|A.���2�cޒ7�\����=�=r���(=�L�Z{�xޣ�NG����d�jz��lf�t�F�s��EO�{�h簓4����Ĝ��Z��d���|���kי�7q�8\Aᔢ�<��Y�����<٤���r`�V�McP���,ר�t��M����L�m�G$��滌�}��{�����2nA�r�̦o�z0� �Z�q��a����E�������+M"�Bq�/�x�m�LNek$Y�f#N����N�G��J{�⦽x�y��u9�������dk�����S%����c��sՖ�w��y|�f���w���[��CG�q����G�����F�B����%�����jXۉ�4�7�b4�6�d�-�F��͵u"�|CwO���f��j�cn����=v=&븶�Av��*�i��2��6���FH�䭺\��S�R�B�nטy�~3��#�L��kE-�ݵ�[���6�x�5�ˆ�*���)%���)RsU��K���H��ΠA%�?�V���0�M���q8d��۪ѯ@��FDa�UV�4$�rb#���0 �+,h;lF}cq�p	c��
ٞ�w9��'�U�E��m��:yD�װq%�vW<��bX��rY�ќMt1�yS���N�<mk�;�TqG\'=���`1�z�5\r��=�}pe���IY��z���T�c���nu���ڕ�	2�UE�Ll����l��FB�جX�� ��$����g]��P`�+�[����T��<�R]nګ�/�2m�0s���0�#��^;�^v���u�J�Տ&�y&��Vm��Sv�g�ޫo\�ŭ�Ǖ;�}�lQ�A�d����;/>q�9y[��+���F��l��֦+6����;މ~�pjw����V/m<�����-1�;R�F�c�n��UȎ��[w����j��n�a�b8Z*�Ë��f�F�R�"�[���ѹ^W[ȝ��d�mIrZ�7-HQ�ʹ���n ���ӻ5�m ƫ�����wm�9�'�5����wO�,nx�d�,��[I
�[8ȱ0�m4]Dκ�Hֺ�^M�f�����Ǹ��]��K�Ά	R��l�>�n}�nOS11�lB'N�>	:�x�1g�cw~qqפnQ�hE��ny�6��9P�*m�wj�iu�f����)����D�J��R��m�U�ɽ�Vҗ<�Zqɭ��z!4���BI'���7cbshZ�r�;�z��P]ϲ7,�����>�x��ꗫ�8Ԏ��C�K�'��hWY%���vd�h,-5�S�Ŵ��x+�c_����r7`�k��3v��	�'h��x�l���<�ҞX���/�K!9�,:�����R�ǣ�Yl�NE�h����iy��a�|K�)�Â�&��#i\jӻX�#��ɒ�i3���$צ���Ħ���l���]��7w����|[>�;+^�SkmM&���x�Lm8�B�t�D��f���,M!���q�a�b��dy1ݽ\�aT5�d^3/��z=�f�E��U�"W8�����,�A����H�3x׺����o�����lF�%mԑL���*���Q�9R^6��r�^,bw���b��� ٯHԓ!m/#��!�z{}@�S`���o������)����]���2N����=���E
m�
�OŖ�,��0%�b�-�y��D>!�>����?Y�2KY1-"�&)b<r_��j�2�� 9G!�矯N��}yN�o����u�>�w<c�g������{���������N[���/�?���������q��[qf���nI���2Y��7-��R�mM�q1�M�c9m�k�g�?������\�UY��꼭�nUUn�����X���^UU����uyUr�꽪�U{UZ����*��^J努�וUj���՚����Ԫ��UU�����W�U�����~��?,?~?c��f��7��m�����L��ٲJ�l�չ��VlF � SJ��(�d�����{���UV�ʪ�W�yU_[���u�Uf�ꪵW�U����5_UU�����yV��U{U�Uj���U\�UU*��g9�֪��{Vj��U[�*��z��{��x�I/1l`&�1l���hI�oR���{�߽���=�UnUUn����}W�UnUU\�1UUJ���*��UUT���UUr�Uf��W�������{UZ�ʪ���sϪ��^UVj��ʪ�*��UZ�=6��&�K)�b��ՍAM&�[�9��#ԥb��u:�5e5�1��9PX������s�Q��Q����Ŝ��m��Fܚ���]Z��g8�V����ɺ���+�s�������3a��k?��?��~��=�7�����:}�+��������É$�$�M����稒M>I��O���$�&ӎ8�m��4�z�I$���ID��4�z�I>I6�q�8㍦�I$�I��z�'���I4�M��#�$�I&�	'�$�)$�$��z��I2�O�I>|�2�ēǏ�#��OSׯI�	�L'�#d���OS�N<N$�6�8�x�I����6�m��i��=I�I$i��	'�2M8�8z�a$�i�O	�L$�>L��I6��D����X��Ow��s������?;����B$v�$9�.���l��{xnUUN�����mi3�\�T��9MH����M$ZZ\G-��X�!kZ�������̒�نr�H�M��[ka������;/0�`d�X3��.���H_-tnL�����:�mtu���q%�Q��yx���}p��������f~�nwQ��&ۚ������Vdm��猬�R^�O��M�[��w�s͇�\0��A���3��,fc��b��m�_��o��ȕ��պ�<;s�"`W���{���+U�>M�������7~���� �D��^��%�%�4^b1�n�xnup�.��������e�{m�v�Mp��m��/qˡ� ݹ�"�}���/3�9�v�̼�lZ���p"����݅�ku��ŕ� �*"Y�YL]V��lYm���������u��u���m�yv��\]�[�LZ��%,��1y��w��ۈy��Z㱌�[Y�LAq���'l����.�x����P۝��g�76л�'��v�MM����E�����'tm�xz|	�$��.s����1�h�qyp�}X��v)�������q뒸�q�w���}�ls���>��N��;�a1^=���[}\�����;u��2a��J�dg[��Y9����ۤ�����9�z'�U���5uҚk�e޵ۦ�ʤ�\�Í���GGSڮpI����aݘ����ٜ�â��t%���kM���g(�á2���n�=.���<lk�P�R;L-y�t�*1�.SNQ��Ik�����G15A��t��5�\k��:�[��.�㳚x�nwf_3�f�v�0��M�,��)�^z7
��<�3Ǹ��>zm�=n�ʎ�=�HQ�^�yg�[�;�7�(�Wa��4��ٔ�k^źtwi�Ϧ��ݻ��"��,Ӈs�c�L��5�	�s�u��0R+q���b�Z��o����WB��֏o�_����X��wf^D�لL�F��qXz-�n5��7d@Nœ�НN�E֣�=.:��t\�s֪�Avr�)�����v��1�w�{��띠�l��9�f�wR�	Iz�y�;�{��������k/�w���{��\�9���9�������Y��������jkZ�!8��Q�L0���m��z�q4��$�a�蘦����r~�����$�m%f���B��;������Ϭ�Yld��g;�t�8#&m�V��޻f$]	�u���A��J��&k=\�V��u闠�p���{�ķ �Ǎ��9k���'��aj�S�v������_\t�wC���2��U^f"�k�cWӸ���z�m��]��:9C>�j�h|��]��b�p�U��!n�Ȯ˼��\���z���9�g,�>0��2L�J"�H�/�cϥE����C����V,��!X��&:6H�+"���蘿���t�����4�[���#�([��h��f�xoF�|��)X�~)�r8J�4Y�e�.��6t#4��z��4ilm���p�$~VE�$��t5�G<�ܒh�#od�W
���ü��!��G�۩&��VE[�1,Z$<�rS�禂W!�CC�Kk�Κ3eq�3�N�BS�p���x�q��u6�m���M$|>�O�����܈��7*���5x��oFΖ(��Rݺ�����R*:r�ţ�zTt�>����zʑ��?.��3��M�zo����lUf�dj(1���\`�+!��&��ڢ�.4.��ן-�ս[u"�$m&l��N}���`���fV����!��C��i�4D?F��w�6���4ql6e�E�:�Ѣͪ	!C*�Iæ��M�P�4���ӎ�m��z�q4��Ǐ8xf�3C,�ƅ^�$��)��ܰulrls��<ݭ�֎�vY��m�q%F�:�oR�nTuL�p��giw:���[i�};���4c>����-R�H8�=<��!���xngb�U���{�������a��"�
P��X5G<�Q���N8U&͝T&��VIeE�����V7�ءS��86���ڊ�i�
�c�KE_*�U��:1��E��O�Gtt�\bH���~4Q㮶�q��m'��I8�M�D�D蘦<>>K�UCrr��n|���b���n�}�Cѥ�h���xp�!Ҡ[]�uC��Y������*Ł���?ZW�t�d̰ؕ��y����hΏ7:!��0�7oy*����h�m��M��+c����A�Y�2U3D4xѢ���b�m7�rl��<tڔ��5�6�k�20�B�yC���S��Jr�l�f��P�������Z�ؙq�/2�q�_Ͷ�n���I8�M�a�X|��~|�XkzU�Em���
�K�8P���Y�B6�^���%���u�5d:ЊGa$�/�8�%/���V�j*͚�$)+t��f\K&<�USٷ�0>w<jM�m1���l��uU{��s{��Ol)�ٕZ�t�oÇ�0���-�~���E1���z���G���gv�ִ��W.Qr��]����<1R�
!�����Px�1�Y����	�I��)Ӱכ�K�!��4�e����ۄ��r�� .�ң

��aV3�ZWg	x;����Ç|&�!hi�8���m��h�e�<�>vf�K�5q����]�)9Ѣ�B������cvhvaļe��e�[M��i<N8�I������he�Y�#�~i�H�7S�Uj9ӫf�L�ɾ��	tPxgH��,���l�c�,ڱ�n�,]�`��^��l����b�2�̓��*��J�Q�+,�4�6Bը^kD�jj�.�6���/(iv��(�i����rC;p~��u��\����(�Jh2ď��Jj�X��������͔@�dK_���A���Tn��Y�+)t�^f3oD\�\r�J���<=,agK6tç�i$N8�IĒm0�2��-n�-��6�Dk{m�?N�+62��@�kϑ좊4l£h�Ь�@�1��j.P��]�m���fwE�
862�D���q�
|�
s��屿tl�Q�,c	���̺a�N�7=�ٳdy��KG�ߋ&C�8p���t�[wt=�z�A�p]A���uw���I ���M�b���9#�U!	F&h�L���hн��'9ɻ#%��8s����H�oϿ?>\c�^�뎶�m��'M$�I6�i�a���X��UC�W��-���LC������7D;Ӭr�4c�"�G[�bhbi��k��Կh��*R���w����/�� �8�����!��><���Q�dT*Ēƒ���Q��=�7�o�G�pA�
�nIa���HC�G��z-�����Sr���7�����l�6ʊ���D���lB59�PʕZ��Mt���+K�
�i�Fe77+^�Yçs��\m�\u��u"q��N#�M�����Qg��y�rGN]9(��K:z�k�؛���v��� ��9~�ϴL�0� ��)#M��-�u7g�v΢��r�i+d��y|��'��;���Nv
��%;h�����@N7=�>0�{4	�*��vu�]g����G��®� N��h��?28լ<T^1lך~$~��uRF�՚���Klc���p�l�[,�T����{2�l�#{TiM�lw�]�-�ֵ� ���<Y��H��`���{���ǎz�ƄbvZ^�T��hh�Cà���4n�������zStiN����ӨTU�<|�5�	0�o�!��R�E���t��IYCG�4�HI��O��.Eｋ���茐&$�]m����l�,�U�?'g�>:oP�<3kH`�D;����͛�������|�={��zH|6����u"q��N$�N0tD�b����t��EZ��ǔ��n��z�1>������56=�` �Ptco�貏h{X�x!O>���e�S�G� ���( �bٵc��0�t;�(�@���[�2��A@�~�w>��f����!��Ý�Y
R�#s��rz�q=���bl��A|��J-�B6Yj^n�0�g!����o�6p� sOl��K8���.�vk�����9w.�C��y�$���cI밵u/����d�?�!���a����a0�
����8p°~0�Th��a�h�a�:a0�,��<0&CFV'O+���t�+�
!�&LK0°���<0�Q�l�a���a	���	Fpx3�:a<x�o�Jل�ģǊ��0�
�	�����كф���p�,���l��F<0�8a1��ф����e<'F[xL0�a0xp°�Y��������������l�
��a��+�f����Q0�x�P�x� �$0�;YP�a�0�ڃ���0px=����lz0�8a0va0�t~:YX;o	�p�(x6<���:�α:�q�����y1'��Ҿ<QFL2<0��aXa4<0$0�<�&�o���p~ψ>(����Ώ���6�f��!��f+���#�<a82�&��0��B9�]^f��o���B�(�����P`���ɲ�DF�2#?"(����-�]4��76�F����7��T6	g�=��{����"�QTHBy"�<�nE=~�0����q���uH���J�
?-ng�����E$t#H�0�(W��yux��JI7���U:�mxut/'��ER�}��G�KM��(Ig��E$&��F����=g=_s��:y5%�������V����ֵ�?y�����U��}̛���7���33����s�������ۮ��m��H�q4��8���$:t�:���BH@@�4��lt�?PH� Q*
����%�������!pD84* ��i>&��y''�;������sS��5.u��%���c����8�ё�E�kPcH�h��*�Cc �81e�F�B�|1bF��0hxꔒ�h�ű��(.�T�^��1Z� ��?Z�����-�wm��:=��8�A��Ҫ��YD�_,�96q$`�Q@����l�c&�yB�n���tXz����nAM֙����#���ᴍj�@{m�xJ�J���(�$`�֒���7E� �N�PfclA<6_�zZ84�064(ŵ�f��Ī��i������(-��G"B���n�ڼ�F�8WAA0`��b(gI�Ӳn�v��9$;�1�%��`tb��X�x{)1
�8t���_Ͷӎm�q�m:�4�!ӥ1�~�y�bp�AD� IR!HHP��ϻ���8[��=�1:P}����Ɉ��BIl�61x�(h�4�1aGGe�8<�W��y9���@��d��qa��Pu �kf�w��4�q���˱�^�����д|Ax�"�ƀi�1�p�.6��ii��d�SG�_�
�>�mʔ�����X���Y��D��,wA܇ww1뭍l*Ke�*$)1p�Lp��<0>:�.{�J�-1hb��I+B���4������K�p+dB�M�x�Lٵ �q#u�E6�h؄�X1��黱�~ 1YiTRX����Pp�@`|4�(a���dB��wekƋ�R�{ �x����;J=�n��n��͝ ҡCCዪ�D�p8Y��u����m��D㉤�x��f!���F�,ў�]����dV��m�J/��;(���͠/	�ͷI����/Ld{��w�n�"�N�Nؓ^w���
�O.e���d��3T$��@����!�n�8W���/��c�*�j6�Eq�\mn��0��<��ֻ~Q��w��l��\G�)Q�C�D'�p�!����Q�v@F�]�ս��Q\r���e'����JfT2�1�з_�jb�b�0,� ��iZf��R�������]["c
A��lb�-��a�q���$!x�t�@<��2�:Ķ5񲕘�s��E=B���������b�Jn ��A ���0��ز���Z�J�;-BƘ4�(�]IqZ���&+��G�����60�J�`p��㎒g}�ǑM�6sF�� ���Z ��2&�ɭ��1pdCfȗ~ǒ��!VV�<1tcik��IVt�y4q���$�
�J�Ֆѡlb\`��+�p4�����}�;��Ҳqt�k�d2:ƪ������e���|;G:0��cKaeP�`���,���ٴP@>��vA1�J�t��������,["�~<x�6����m��'M$���M�0�DCE,�F�Gdz'��GoZ����������4�ų�q��ɼ'iG�f���� ��9���%��lm�UX�#M�-&^� ��ϓ
�m��L!�ғ���Г68(n�xh��a���&���p�kfObnt�q5v��Z�'�N7���j4��4�e$��ҁ�u�GF�F��L�зݹ)#L�:�� ��)S��&�"p�)�@>y��@#%)/��<�H^�0Sv�TMG3�X��q�Ռ�!�G���sTL�a�e4A�C5B�IG��D=��U�vbydވ����_q���f��i/i�@`hb!��E��Y�)���.��t �ҟP��4j�?`�AbА�J�Ʃ�Q��8�?�m��8�i'q�h�!��Y�����M���X����7���blhg���	m3Z���8@�7߁��f��h��0<��G�d0iB ̡��cI�0i-�b8RG
H��n�Cq�
�6Apm���4�b��gyqӧh`��4`�l��xf�k��oj*I]a�f���`����6�*�eQ �kb6]��M	pz'��yʉP�#0�A� ����F�D�Ӈ:�=?�/�D��"X�@�[Pb�o���C���y�\�Ɲ�����q)"��U6J�+4g�C(��A*�P����s��bmb��2�Io���Ih42�l#\)����N���C��������ym��?���u����"q��N�<t��G�h����B���c�N�R���^�S�y���R�	��sÍ�6�d�w�x��rJ�Ag�b����!^�t@�������T���7$T�0�d(cL;��^�0��G��4���a�h6�nůQR�gJ\�ޫz�f�kQ����h`x��Ih�,��2R�\����1	�x%,'<B�o��(��r|Flt�t6Z�ų���Cg+AL��)ŭ!"Ⰳ�)�:YE0m,��pة7�
Fk�9Pu2���8B4R4SOE�=:}/2tL"��Nu�q7J����BU��q�wW4o�  |���)�E
,b͎(���@Ф��,���"G�!��Gqu��13��ii�&�E"�pcd�8x����:�m��8�i'q�x�D�N��:o�H�{�T�%��RmE��k����B�A=��ך���"n�ѓ��+���W���552�?+(�!b	�XhE4�������G��_iͻ[�p{SoD��hM#�E�Ci�׍���*����Ӑ�-����l��N�"�Θ\g`Vb&I�\.��]�9/|kA%$�6�cB��Q��<�C���$=��o�t�B�z�yM�L5"�.18AX�A��pa@�=�e��F���*�0m��K�4�P�P�5�3PQ��4|s���؛�g�$D;o;8�	 ׋�H|
4�Q#�,�A�t1�&�0��m$�"��|uTX>ot�ƒ4�YP��0���9)깢�R�N$1�%F�V�(i2���xȑ��P�Z�X0:�<�G�4h��%ӻ���E��c� ��>L(l`�.���i��h[e��	Ye�2��4����/�%�X뤮������q��Hm�g�F��-���v��n\�48��,LT!0��+�a��`�i�.�X�D�X���hZ��&���J�ǼNEA��%��:C�6a��m��8�i'q�x�:t�1ӧ�x�;��(� 1��o�#�Rh=�;"������tk�A�!���f��')!�>��
���r���TU��NZ\l��Ϝ�t��ѳ`6�%�,��&/!��C��d�Q!�3�$!$�m�� ��4��q��DSe"�06!���+b�ͻ&셳5�z:sn��!����D�v�e�˥��J�-)��J�}�4W\��jA���#�#�K��ߛ��0-4u��c��!5��mI4ZTmC�dS`Т��[�t��\��KC4����l����f>h7G�4�p��B�,����6�o䓏M$�mƜ4C2Ѣ�4h���aRzTԨ�wkN�7����M���Y%Eb��ńBc8�DV������X��ze 鲂��h�����CD�dP��z:0\�T5�8��j���0�ѿ6��L_[@C������G��X0/������Ĵ�e���QE�b��(�ؚ$�����i5�S�~#�ѐ ����ll44pb(h厂����HCKL��
�|m�0��g���P�T2����(a �ƅ� F�#�cH �FlhZ���6D�Hf�*Mq�}���TB��iB��K���#%acG�H2Tr�a(`�bl�9mć�o����˯�u��uԜq�i'N4�/a��2�������JՍ����T<y�I�(�J�����(��Ť�i��Ę��S74yOD�Ge�OM�P�����Fh�eR�"L���|�i�f� 09�WJ���	YZK˵;c��|�oHh����n/!���p:4��������<�Kc���4�ǧN�7�&����A�zc��@�'��G�I�|�cT3�62�Ċ��@`p��hc�wh�qK���>�����s�4q4x��p�(0`i5{��|IU�g����:D�%���߷D�������`X���"4iߴQD!L�zII�g�D&��Q�so8d�n���-�1tiLo�7�-�Ihi`z�� �q�B?n���O��C����&�	���VL6L0�x�l�0��<V%Fp��Ѣa�0}0¸;0�C
��a�
���t}N�	��L,��|W����L'����h�
��d���a�0|0�a0����	�	!�8?��a<x�<N�c�aD�	�&&�	����oFSxp�=�����GÑ�
$0�x6a0p�h�<8LO&������a����	�%�K0�a0���L0�a!�S�aÅl{�8T0�?�C��<0�B`�t;,�a��	�������dƉ��<6|F|M����va0xt�������l�n� �&l��&!��t(��'N������p�_�a0��0�Y���	FF�C�0�:2�"��<��>�!���A�������e�ML0��	�)1ᄆs�\��tUMn�Uk�4�a��H�'gr�nӦ�t��md��W���[=>$�����X���ߴ��˫� D`o
��!,@�N	=����=��Ɖ����S������UȬ��J��+�S���J��^�x;�7g�T���+�5)KרY7g��8�ְ����B}SK9vd��Bk��Ҭ��7jۛ�a}������t�CNq���0pr�s�+Ma��j/�Ó�y�'ՍL�nV-�h{V<&g�@�H��ͳ䈶�KsD�k��W݉'��v�.�p8������hs�� ���-�����0/[qR���}Ʈ�y��[�U�!9V2\�$rآ.��<ˁ\+Nb
�XX���~!���8�\�����S�߳qɷq"�l�u�m���m��,7nV�DE���0#+|fS��Dͭץ�Kg�@iJBvX�����Vy�ey�����3\c�Bi/=Lv��SJ�c�QD�,��h���1�����ś�x�a�Φ�s�zŰY��kyhoJ��@�Ԓ����jfn��Z���&�͠ ��:E��=Sx�b#��t�Dقf8�K�[ky!�--�c9�Yq��p�I���I��ѷY@����i�i�D���\�ؤ�ݵiW�w9�q��
�8�*�pl��B*�]��:�a�½�)�cj�>�?e��r�`�4�vkt�n�]��.Uq��~S���A�����Ůcg�p;�u�!�q�\�vK�XH�ǅ����[rm����lV��tY���v���Z�%�J(���m.��J��|�9rH�= ��s��?K�Ό"�G��ủ�ө�����k9�?���{��33{���35�Ǚ����9���oKy���d������f�[��i�\u�Sm��8�i��O��H~ �:c?^�߄r^K3!v]0��c�ݳ�n���Qu'C�T��r��m�B�q�Z��7����ح�1\����-��a�Wc2:� Ӹ:�9�n���'v�k[�%��yw����f���^s�v۶�C�̻Ku�du�f��M��J|��#��'we����ѷc1i���\;]��&Ʊ�oW3�c�֞Ǝ�u0,<�v����lAs�9Ɩۚ]����'Vㅹy�ꑃ%��݈'�g�*X�D�,.�d��;s�֜�?<�/�ㄊ��&%�Ҝ?�p'�3��<����@��fcQ�[8l��$~35nJH�hg�A�:��&3��4��G7)ԕ"֒|"k�Pc0b|pG1�w�$/�H�811��|0�`��!�=�-ʢ���ļ�kvA`�cH�b� ���A�G��CK��L�P`u��cF�T�-�-��ڞ"�w��:��Ŷ�ecKh\p>��6�Wz���h��4�4�� �A>śM-��Fx`��QQ>r�d���������n��;�:���zv3�9];i]u��mI$;�4���s�q��>��Y�û��Шf�}C8\Mc4�n!q�m8؈��i�Zz���.�����uԜq4�n'�4�/a���e��Z��������
( �S�Ё�H<
|A��K�P����aLB�%�q��g�H:uB�|t��Y��h�>$0bؙ���4�Ŧs���X� ��2ZJ��@Þ�׊���]Z �3d=Q/u�p������f |4.3�*�|�Kc<\��8X�2DNt����ų�)a�Z�`ٜ�0���p��'�����h� û��4E6QfB�/m�|0�
�Z:B1��x���G�o��]���\ � ��}����g�xI���xvq-���)���|=�h�(���DF!�u�=s��ϟ=M�����uԜq4x�ç�t��D0c!�,�ETczt�8Ҧ"�&������~����'HQ�&��pzm����5ؙ5�C 0(�F�A������4�2.ta�f�F��V�=9�R��&�3c6�W��cL635;C
8��C,���Nџ�s$V�N��$�,����Cv9�����@N�`�R�o]x�ԍ���<��$6�G!��g������&1|4p���yUToDڃ ��q.�D������s��p�1BW�kz�ڕ#�o� *#�0b�(]�{!cA���!�҈>��BA�@tiX1uB�
i\n�)����[(�Řt��N�0�ǎ��I��q�^�x��_>e�����x�n%IN�( �x�,���~�)h&ph27�P�g��r�����42׿F��<��s��X21�)���[��K�.�d�H���f͝M(��!�dF]�<��_�iu�&�pވ�@,��7�!N��v`���4p�����Ǝ�\Tu�.4�*(C}��槇>:�Kơ�ϼ�P+�Ӧ��k�:�2\֜�`C�;�dql)0b��A�vWp0�Ԙ�)Y�s��+�C* 5������{�-|�i:�i��q�]u8�i&�Oi�]za�/|��8g>�R�����k#dy;$�}	�ɷe�n&�\X7�����9��e�|�����������[o��f-��i�иɫc�Z5,&���mX�f٨�cl�Ε��~"�q&���4����:�v���eaf0��ԗ����+�TO��9l�����z7v���)nk����{|��*(���B�.o�1ởO�#��j�f	)3H�f��p��Hx��<�`�����Ț�����0gq����[����_����G��΃]��L�ro�6t�s�����2�����b�tD|Ň���h�6kc(,|i�9��CM��#
3�h8�*Ň:}���g]�3f���2�ԕ�q#s�
B�LXF<?B�����A}�G6h׸����Z����/�}p���>>:||x�Ӧu�M$㉇q�^�x�/�>4�k�ҘƘ�4�2��WHoMT���͵�u۱��0`���b4Q��pz:&���ύ�,�-`�q��(�k���������*�{>a�a��G��%��C=��a�&6��o��uL�Fy��>�a�a�"��
)�
ލ��϶���v�M��h�_U��e�ʔ>��=����=/���<)���sdTY�yY�x�Ķ���}83��Y�l�}x>�h���0��Tm<:��8|�40��0����q�뮸�i'8ӌ��:c���?S��q>���тԝ�/�ðh�����;��Mv7,����A��8�E�D�6D�����tt8k����D�p������GFh0����7�TV2�A��O�O�UFit�6�Sq$\�����V���G����Y�߁�(�"�s��M�����MM,T{���Uݺ��f������D8t�t-�\���0�ݖ|�Pdp��쪪��d�8���0�6k�rh�ϼޕ�h6�3>|�N�o�|��>!�."��H8��M%�G|t�f��8a�ӧL0��u��H�N2��ǌ���,�m����G$�k{��llLW�g>�$��J�<|0�[:C~���k��u��s)�g]�rx��Нk틵�C����H�g��.��[3ó�fηZ��(w*�;��x8!˳��s�:x(|4Ϸ̒J~��za��m��hхn7�cֽ���\��0�0a�D������-��]T<�Qg�p�����Svx����φb��0x|t�Y����oE����'�㎺��Si�x:h�
CF�,ѥ�asn;n��;�y��k��ն"�i�%������5S�e���aL);��[�/<mG;fIf`8m�$�ݗU�ښ�����MS���a��b���}�hK�袜A�w~�b��}���^�����4Z����4X��CNk\q�hh��CczsM$3r�'d1vsST�*-���Kg�Jtή�5M��/�@Úc6m����2T�Z�FuECPx���\6�l�W^.��9���u!Ih��ː��A<)AcJC��C��I |C�ϕd�Gŏ��Ir��m-�xtt 3�<�1�J-����8:����ц��Rg���F��|p٤|j4�������m^ޜ�n�Uk%�[�	����4������f��eQk�cz;��?2aQ8MZ����1���q���G�0�8㎺�:�N$q�u�:t�N���I(^�T��y�����|Y��z��4w�Z9p2��pa����W�p�� 0g��L������\��@f�,��,�k`x��`��j�����R�٣���	�,IM�n�p��a>��=�O;��5���ѫ)l4�WY���tΟhΟ9��YaD�a@�3�l�}��-���J�xPÅ��4Y-Öp3�3�8k�ܨُ����f�- �͔|�pц�g����°>&L0�2<&�fV�G
�	�h�`<83
�	�F����
�d0�C	��l°�t�:>�'�	��&�+&&�&��f���_8W����'���჏aX`N�aG�e�;�0�'�Ǣa��	��+�0�a�p0�a���3��ä0x?��|#�������xl�o���&��Q�Ɇ�0��LYVY0xa0�a��	��	��fɣ��Ä���C����l�a	�F�P�7��/!�����ϏW���D!��gĳ�cvL�#��0�<�7N+f�a��e���a����|t�
:WG��}>'���3�`dxaXa0�aD���aq�LEь�/&�`�g����lxB(��J0�ݓ�̧���x=���	���������ޱ?1��P�~Z�a;�����&�ĵ��I�����ư�O��g�f���w�o�＂2��-�O���s�EFO�^3�0�(��O�i%���"ޒ8Ҥ�
�>��=�`�T��*�k䲮,KA�|~תϼ�0#���?k�}a'(<U:�Xz�>?C�bMS�G�����mߏ���o�ϧٙ���y���w�����d�z�{\��k_5����ʪ�s�w�ֳ��:�n���8㮺�N�Ӊ�:hѢ�4�;���0f.��^�(!=��Q�ѱ���@e�+P��lxp��g4�4ϸ�iCgFy�Ξ�ن�ٳa`φk��,�,���my<:s���|���'U'�U�B�mcBOD��-V��o$���p����0f�����h9�l����᱔b��!��\rJwٽm��IY��׳�Xb_�nD��k�ڃ��۳�"���@�k�)�`�>:|ksd��E�lTa��$>�K@���C~���{�g,6�iƓ�6�:뮺�u��Gq�^�<e�̲ן�g���%�^T7���PDD�<�o��ٿ�:�K4s,�c-o�I<�R�ѵ�GǗB��(�c�`��$��N[�)!U�����U.q���ӥ:-P������&B�@a�G�۬nx�8y1�ȍ7ף_6����c0�I�ҧW-��^�c�G�͔65�Vw��7L,��O��Η�JMn4�j�֩t���|<1�g|Q���S�R�>(��)��Ə���{ߖ�Z٥g>o�u�ٴh���θێ:뮺�u�H��u�B:c�K����!��^�I,/p١'qБ����/dXy�3��$���]�e�d�
xAp8kF��1�����
 �����$�eX	�"���?�!�'1���t���l�g���r���<YxQ�u�f:�o�\�@ ����?�-6���B�Q��h�?���?���L1�QS������`�S�7���D�f�������]Ͽ�x~`?����pcˇ��~9T꜇�ض4h��c+�p��,�8X�42�C#i���Ygc�����Û+�n��X���X�3��e��{c
7�C�O���x��#�j��LG��=/'����"%P^P����^xoDDO��H�?��!d��
��Ym����{��H�Zz|�/Ű��h��4/@�Y��*UXma�_�?�q�u�]N��$q��F��h��Fi���������}U.e�i��.��P����yP���@a�����7�8��(�4ٔ7FΠ��g�x�T�ȶ:LҢ!񮐣I��B>�Tb��z��^����S���7b���вW,�6��T�Z�:��,d�Jy�y��z3>n-�.�����T��e�,�GY��\8�@a��~�˩M�u����x
:p����ǌ>8�:뮺�u�H��u��:c�I�߿�J��Co��uh���f8Im� ��|���z6}�n�"<Q� ¨n\�ݛq-\���[ި�._� Ëç��	΄���Os�-�+,��Q#���g�xa턚�r1��gHWڒ���Fց����Ȯ�랧)�GN��..��壙c�<���׺6|Q��+lJN����ʦ�k��tѣˍ�"���ݮ��A��NY�HcR�P0�%�١���Qd8x��gN�0�ӎ:뮺�u�H��:���,����2p�ࢂ!xb��Sˣ(��4�R�������,�\ZJؑ�<1�a�6_���(���12ɗk�Vx{{��Yz�~cT#k�B�>K���A��,j/3�RU9A�X�d[>%�����m����)CEZ�GgO���:k좪����W��P��6Z��lvg�*Je8�0�|IcV�Y-͖x���_��7R��N�a�CVh�;��K
h�Ӎ�u�����?����u�S��>�P�:t�N���f�m�d�7,�&�Ή1g�N���s��+�G�"����B��(��%0�lku��7F6?��k��|<�]G�Nsd�s��_����%Ӎ�K�m�����&Ӓ��a�h6�I�]�
�V�p YC��=�$��QfXj
Dd`��3�R�t�%Mլ&��D�*YF\B� &�`��1�(SJ��6��"�g"�h�� ��� lnuZ ~t��c63�0�3�a�E�͞_6X�d>�ŚZ_*����(a�QR�jΑL�Ǜn8|�60��g,GY0a���IQW>n|�uRxÃ$���}�y�RV���i$��j��<w����(���*�^�6-�Z[r\2�rd�/��h�s�7LD?�W������O� �p���G�8��<]����xӬ��u�q�]u�S����t�
CF�4h�qۃ'�-�Fʚ�Yᱰc�Q��1;(پ�CiG��Y�� ໍ讐���L��>ce�a�Y�c{85�[޷M�_%���;��<=L���c(���g�oe37$�kL�
:l�\�����Lc��D�|tӛ6*IPe������~�#i���a_-aj�iψ�[�f�1�E�4�0�<Q�9U9R��U��9��Κ��|����N8���N�]u:�'�>u�B4Y�UwTڍ�ll�K���}Ը���85�W�q�������M-�4he���zIZ,�\�}�7������(�䲗�5�znX]�S>>�nCE�6v0�ܓұϮ���,���k�^�T�?�v�}�}$��h���?lI��	`���E2I%`��-Y���1�K�&a��(4U/e}��4Ȭ����*q��/�H<�Cc�z,�KC�Ϗm��kg�g0�z�������m�n��q�uԝu�]N��>q�O2��F#�<�U�@�ce5���pgt��X�}
36ߍ8mQ�7���p����,�֤�QR��l���C/3�a"��ߤ�Ա���U�|�QD ��Q�^����E�|���,(`ψ�^�<y�|t:0�`�,�g֖�C�d��4��ҋe}�̯�������0�Q��ᢈA��a���>��?c~/�N�,a�t�w��xY��4���m����O]'�&�M��i<x�I>ai���&�|�&I�i&�m��i$��M$�|�I4�z�I>I$�OS	0�Gq6㍾I$�$�(�ORe6�q8�q��0��0�L�����2��I4�I�z�箺뮺�$�$�e����O<x��	=x�I�i�	�xîu�[u�u�M��|�aL��I4�m��o�m�]u�t�I&�x�x���4�i0�8��ێ8ˍ&6��x�ԓI��8����΄lu,DKJ�!^�sJ�3V�4�����K��bxZ* i|Q_(9�`�4�����k�(��AZ�M�n�`�$3�W���2�c��5�K)��O��d�ʚ�[,v���@R��H�Ob��Z���<EX[��;�v�;ۺ,�<m1��,-]9aEO4��L�"H
qqBN1&8��4�>��ق��;�a��A����I��<�_.�ZTT�M"�BkA̴bwv��K��p!�!�U[5��~R\�A(��s�Z�aL�n�9�zZg��̅�~!Uk(3_4���]���������	��+�ǵuXԶ3�S���"XP��G��-��D";\��������*~��+2�X)��&o�C���Aǅ�]�{:�H��1�<�Tm2]�Е�Qg-$[x�E۞eBy��S:�1jY����w&��'˴N�}s�{%j�7<Qٵ��>޽�^�c]�))u$!�,����$��%ӌ�\曐�[�v5�-���˴��'<�l����%��<'���\tv4vS�����C��ڷj���c=�\��M���<vǴs�C<\B��6͸SYjV��w��m˱o�����B�5۳���n��n������Wj��g��~����k���ֵ�����ګ��{��Z��Ɲu�Zq�\q�]u']u�S��O�~(B:c���a��5�ҽ���`��7ng��=T���q�δk[g��x���1V{QU���ІP�x�գ��q�'o2*���6�X�Y%j��0ұ$Ж��Q�o6���JHK)V�X��� ��L:�J]2:Vl'f8M���}��n�����cJ�1T����k����ṕm������..x��c�s��L�k�n�m���#�U�w)RM��3&���Lȓb|��2ԏp	 �[�1w�g�Oj����{�K�R�����Bf|�J�lI""�]'zu֪�@�R}�����i?��_���^cpc|=�S�΁����]H�Hw���'�ȓ��I�����5�H�ds�t�oEP���1�m�I��h��<��BG&��8C�>(�gc+>�o�ㅌMp ����AgG�7�a���Jom�xe&�c8c�o[
/O��S�2ښ�Ɍ�ct�=>q��L6��i�P� ���w��L�����9*�H��Ѣ�<l0���n��q�]u�뮺�u�],�f��h��l;S�ѱ�c��9M�o��`�Ok��,���z ��^[�S`��l3��h�B�0ň�<hҴh���L-y3cB<��7�����Ӿ9�v88�GK7��p�J�>�Hef�dd��n�R��0�7wLr�j��V��LB�����"��p�#�#J�!c��qY���u�HMTxf�QBfd)1�!����0sE���b���G�'�8㮤뮺��]u�JA!ӥ;���8��]�EC��D)p\E��,�k���+Ll�,a�4�ç���Q��)j��H��;��5]��6���c�Cpg��vl�Pa�t��lm��P�W<͑F2�ݢ��>�����WMѵ��cח^L��*(|o;m�w��(|v�E�-iQ�ql���Vh���0�w
��k�c�4Y�H���E�,���3fϽ��3j�Uj�ʯY��j3�G�Ο���ihc#�R�f�43�<|���8㎺���]u:�,�g� �h�F�/��M�H�X�8x(���>>��[q����xVh���
���ka�}�Xp�_�>���Q����3��e�RTѭ�9�ɬ�m�tW��1p�ƈ2����4M��>�rhV0b��e6<��㥨h��!\�Б�=}a�6�k�6��᱌�))`Ŷ�:v86��I�(`�C⎽���ش0��Ѥh0��~��	��	*�"�{�����Ə4�<�����̧u�Ӯ8㮤�u�]N�믓���e�-�Q�D_��ߝ�?"���aB&�(D�B�2[X�+���$f�p�a��F�FEkQQ���
�h��~�}qnD^o[�q�X�Gqӹܛ��ՍZ1"xy��!�~�@ ����*E��Z��~�f�n�����O��Lp�8jf�`�G.�S�$(h��Q���74|BY�|�Ç#D"�ݏ���ٕ;w�3�����!Em��c8��X�d[�$�c7�\>��Y~0�-�4xχ���k=
��>4�t�ų��YG�Z6�A���|�m������4h�� �W�ݘ|l�yiqC��c�ӿR�e�%U�K�6ٍ�e��-��#����y�`��Q�(PÀy��0Z�t��5v��ՋA&ڊmM�R�{63�^=U!FF�Y�E�:I��?�q��:����u�Vx��d4h�F����mE!Q��cc`�R�l��1��}���jX d)Pt���֍#D�n�T��t�>��w"��8�΅j�a�(����l��$��60�&͝6��˟m�X��C���غXy���<�H�!�~�\��#�䓧O�<p�j��	e!�1ɳ>�G*�,����a���,��!�������Y~��^��0�-'f<0����u�uԝu:��]u�|�׌<h�F��զŦ�i����1���E"�A�Kk��o���>�/�����h�B�0����RI6ʯ�R�����h��0��d�mɸ�â�{�~y_䕮��䖸adNI!��$ae�dd���	�G}�V���K�E��q���a���?b4{��*Y����a��ٳ�(����"�p�	����<M=�R^���GY���C4YC
غ����&l��Tm������1�|��p�?�q��8㎺�����]u�|�׌<e��������RtQA��Cߩ�I���vY��|B�Q�r|�⿡�QlPP��#��ёX����c�!�v�g��:�l6�0�h���j�41��R4w���#�GC��΅�C63�tY�yn��?�C���᎟L�7s�J|����׎M�ؼ����ud����zG�X���
z�|e���!D�s�ό���Ce#c�l�æ�0Æ0�uē��묧�=x��Yz�������X�Z�6s��Ql��%���BW��i�\�@Lh��㆔@�H"Td_���qJ�F�u䋡dR��9�ʪ��$�bH�G�!1��Q����t2��71�|g'�}сꃓA�bOv��el��n-���v��:iH�O���DU���Q�aLRWM�w;C��w9~�9"8� 1��0B7o�3�=�0�=�d# +�fD?^4��,��s��h�R(����S�9���C|�͍CᔼR(���YϹ;R�Wpᵣ�>m����;��*b��-�I
0���Y�d��F�-�Ǜd|c�g�p��T0�$�f�ٛ_���{���|�ՙ�p��D�Mi]�+]�����u|���rz�/>Z:Y�>�GM�]8�cm5��)��Q�ph)�|{C���|m�۩8뎧Ru�N�뮴x�ed4h�Gi1��ĉr:|R,�&�,�@�eH�#�A�����S��Yn8g#��1�ڂm��U���b�<Y�ä(L`����ueU�g��+4Q�(a����Z(����)��|gM�e3C(�gXپU��)U)���Q�A�1�/������B�~���Z�l��3U�R6�I呾��zzzyy���k���,`�c,gŞ_r����x����0�ܝՍ{��eQ�.Qc��E�~�*�r��b�>c?��ӭ&]2���I6�M��6�z�q<x�&�N&^$��I'��|�m��I$�x�M0�q&�OSI'�$�I&S	�i�z�N>z�I2�O�$���M��N4�L"'�$�)$�I��I���D������I$�I���]i�_>t뮞<x��	=x�&O�x�O�OS�$�i>u�]u�N�]q�2�'��<I&�i��|���u�]6�$�II�z���a6m0�O����O&	�>I2���Q
<x���e�75N�M�J��ǎ�~��sd�T{&��ثaޗ\��D(J�\/���bL>�
ȡ�n,��w��A:=ޢTH����%↡�P��b"=(s�ֹx �\�[约g/�&�F;Z�!���X�Hk�r����RW{3x�x��]Y2-|:����)�<_6J�q�r8b�lV˘�V6(�:Rj��_�h���f���Л>�w�&ַq�w@�_�!g$Ҕ18�
��p��u�I5��Y�[O����Ϳ�~����R��?~����w�{���̹�w�����W9��ֵ���U���ם��z���m��u�S�:�&a�<Y��B4CG�[0WU���}܀�dͷ?8P�T2���j�3F(�4��u��~X���3��j|�4lѣ����|���%!D�U'4�|���d�u��Hqp�e�O�e�>L�k���fT���.�pc���а٣�4̱����yj�*K��h��nI� E���hag|l�����!�ȳ�^m�9�y�Y�!Ã8l��:뎧Ru�I:뮲�2�����wǗ\����m���tQA�ϴ<�x���?#��-h��x�[��i�R^�xEg��xC��2s�*�)>]Yij�������}��ϟWs��!�������F��`����C�
�������-	6Y��=Vˡ�����Kħ�A�����v���a�GIc�s�θ۪�� �A��|Z(����j����ꮍ�a��aC0��y]�w|�<t�Q��:Ӊ�ۍ��u']mԒt�4h������7Ԧ�h�����	g&e�HuD�AQ���J��R��q�Ew>^K4v:��)���`�n;8�+���M��R�g����}��o�)���qu���_{�zD���fھ��"r�`@��^��,�Fo!���=J�*sf�o�����ўs�'7�����`�<��	�/?�A8��1C$����5D�^�O*�7��0�=
;��k�M���ܕ_�/�94X���?�U*�7��H�\v��1�"[:x�K*4��x�ӉB�(��F�1��Yf��3�a�=ۗ��m�l՜d����Ϛ:l��cQ��E� �{F�!7���6�uv�۸��qf�Ԝ����m�U�7O9��Ə��`�p��0{%�EiaX@��47$ֲHl�sm��8||hه�a��I�\uԓ���e��<e���]W��#lY�o�c`�$"�6(Yc�1Qa�B�o�2�(�h��x�=�I:ǣ|ᄑ�H�(���=�V��,�D}�#:�㎺a�K�<߈x���M٢p(�f� ���s$�?:v��r��<s��A�L�]��lm	�~�?	D=F��Qs̅��eQ��e6�����飧9���;}�IZ���#�nkcŔk��͜fa���?�N��:�I�]M2���QE_��>�������"Y.g���0�ti�I��k�s���Ǆpo�>-b�٣���٭i|C;h��cz���٥����I*��������`p�.��0c.�af#FEf����%����]�հ�)c���r|'$��Є���2IUd<B�/�I:tߜ�ꪧQ3�8l�C�6}���}:��� ��.��ʔ:�:֍��h���F'C(*�>�>�=�֤�.�83C�i�ޖ����pٴ�[83�Ν0��O�]N��:�I�]M2�ǈC�N���^���N,���7~
("��&Xt��1��N|m6;�S7.��7&)ןNr_�?��
!�A������T�խ{��/e��dtpO{�7~��Ez#F����J.����}v�6�J�^!c�f�65Ѧ��oE3O����P�6��\]�F��=���sC,-�c$mk���>>�L��?�Y��	�e�#��9�RUA��i��Nc6a�������1�=?�m㬿�M���ԝu�]I:멦Yx���Ye�W8x�!���.H2ύA�c?[l|ocr��%L�^]��6Ynb1@x�nI�E"م�YM\MѴ�#��39��䑬�Y�4�5N���ۓ����i���e�+%w��߈��d�?f�G*{����c�@���t�z�Xs��0�Y]��/7(�HK��ڏ���
'ל0ҳ��(�ôQH|n�nIgǋZ����0�7f�FmY�ņ�YR�+���lt@a
1p�/���򮊫��rti�`�0M�&,q�c����0��cmSl�->6QCq��E+B3�ێ�D?E�C���[h�)[G�P�ӭ_ul.]ld0�.����F6��yi�WZ~8h�����m'S�:뎺�u�Sf��!�F�6bo�S"��b�!���z�'yr���y�1��lᡘ�rC�ą0�p����:��{[��BJ�:l:1�i�<ilgŭ�����ue��kƈt�P��u�op��'�����GJ�T���l�6��K,)���J�L���󏇧�	!
[��vxa����et�>nH:V�ha{�qm�m�4-�����ƛr~o��PQ�xӮ��i:�I�\uԓ���:B�N�(��	E��zRr�豱1��{a�tP���~���l�H�Hց����:�V�->Ұ�c6|�Bh�C4y�~Q�f����M6���q�CLYU[	�>��yῪΔ�tx�f�!�(8Q]�*�:"ъ�p\����-���Z@3F���P�-h~g�Ҋ&ى�E�7����[+a�cp�@�x�Oi��m��u:����']0�F�BѣE�<p�H��/�cbgaG�(��>,6xQ&X|�.7�Ř2֟�������C�q�+�	�r�ȴm�h�&�&y�<4�l'l;۴��)l��RS��=-�n���'��'��u|�a���fp6��񩅓���5����ۀp�w}CtW�7;$�t�+�Cۢ�F��ag��6��/c>\[ݷDhi�<B��	�	��_��S�72�}�B�5�e���N��{,���m8��SI'���$�H�I=a$�z�i=I�a&�$���x�-��ԒI4���M�����I�I$�I4�m8�$�z�I6�O�'�0�o�e&�I6�a�D�M$��ĒI6�$�<m>a=IĒI$�&Ye��I<x��Oׯa8�8��\u�z��:���$�i&I�:u�u�κ�z�e�M��oYm�]u�n��ĒII�O�	�M�$�	6��Ɇ	0�'���I��z��G�&�D��#4�D!�Y�Z���pfmC�삛
P�
�C���5s����{!8s	��L��1�X��K_᥻A\r��ۖ��(eJ4�Ɓ��
�X:�+.?�e#�ɬ���V~�r� V���qu�hWP31݊��=b0�l1�f�m,����[�����ifdT�ٯ1	����={c�X]��3��5��>��	�=�₭"�	�PGk-B�H�e>��M0D���U<X�b��lJ��	#~B(�H��n�2kYC饥�y�R�ZE�9Ό'ӫA6(�{V�A?L>��?<�BD��ւ�T��9��$�ܫ2���n��E�cY+&HL!RJ����҄��귭.j�Uܦ3 F�Jq�jՋ��6ȴ�HMĂ.�K-���ءq%h��AP����|'J�j2��B3���<w	�%JGR&U1O�GnJ�8�U,��K 0J�5$i�PA
���??C٭q���1n�U��{)u8J�z�.^z�K���TW;g=�xy\݆���T����Ɋ���DaJ�t��I�S��OEeY�b��1$�</^�Ʒ���ee�U5��-�$������2y��������]�V��b�cñy�78�l=*p�:�����@��T���i�K�ӷ��!��>�Ol�.�XY�e%i,m·��vb�klQ�l�c���_�{�_�*�W9�c��s��}�}�{��\�lw��{���W9λ��>���]m��m�]N��:�I�]M2�Ǐ2�ҏ�q�#u�T�\M�Y�������C+K���<�h�]����4g������:��F��ɵ� �s�Y�=�i���[]��vƠ�ܔ�F�<'d�sݎw� �m��T�
�/~k�=����8��;j���InҶ��'!L�n�=5雋-��0��͐t�
2Z�yk״5�Vslssیs��v�ܶ�'O��������;n$|E��`"�($���v�ǝ��q�Q� ���7�ZZc��*�*���'��Fe��]�:e/e�48�9(\A�ʊ��~�����Z�x�3�]_	����Ƌ��^<Ce�mFqpٲ��ttb���EB�J��T}�g��j�vV����5���a��"�-|>��$f�0�C��3�*:*�x٣� ��uZ���zy�����^*Ԗ[�M�HY��nYg%�/�m����?r�!�:Eӂ�6�lpc�co�>8���������q:�I�\t�Ǐa���4B��)"�C`}C�>�n�ȕ����qyל�r4���m&��1G�דchf8R,��ףvh��*i��K�͡���@�@#���g:w��E*h��_hê.�=7҆��"c��X����/l����P���%:C`�"��`�)��Z�ӢQ��~���d����irVѺ��[#S���?���a�ޞ-� B��<ܵ� V^�UZ�{2�sD&��:��1"Ւ�N�x��[ZZc\z��:�6ۮ��I�\uԓ���e��<e�^��[�Tp�gv�������8�I>O�lc��n�l"[,M� d-6A�*�i�;@�C|o��p�
��M����<�0��ߪJ�?q�<�|~�}�u4$��*�g=�d',�Ÿ���烚Z6C�;_h�3��,4u1��� R�!��cc�$�j�7�X3���Q�QΩc��B;��m�A�h���j�)ip�j�P�a�b�G���L�p��A>|���u6۩��N�㮺��x٣D!hѢ��n�;Qe\~�x�5������3ƎfT�A�h��/c�E��!f.�g���?8�E,`��Z��/���;��o7�����
Dc4{e��m�F���1xy#�-xa
kE��<���O$��E��
|���B��C�S��v::5��{G3wS���֮],6p<tL��ފ!�3��A^�sڌ$#,�Fl��3����V��]8h�~Z(�x��n���:뎺�u�]M2��!�:S�>u�0�ۙ(ۮ�Ҹ����Z�³�q����3�M��ń뱯Xu�}�}��:��1���1�N�[��vƶL��-t�{P��i.I�u�諸�N��w�v����M)h�w��0"� ~fğ5�jG���̈���d'���8ыz�w]��Y�����aۃ� 棞g�0�G!7TQm6ω|��������d67�� 5�w$��:��Ԕ����]���,�o][��Zٰg|=mY�7����@cEUh��f���<VQ�c���gŔ�X�+~v]�{���gp�p�����=Iq��L��(l��A��٬MĴP���/C �	aU%F�U1�8��<�����i6�i$��\u�S��SL���ǌ���^a�"S}6Ux�u�
9<�^1$��X2q2|��@���t�Eݜ(,�~n������^���e�ʲ���rUt� �FΈ�6T�,��q����R(�sUԻbm�l�aG���?f�p�.s��Sw��#�j]��k%�[�s���Y�w�������~!�F�)`0��pF���$�^y��0�\��Ѩ�8b�Q�al� �6�m},�x�ƛH�<c�=i��m��q8�N�㮺�Fx٣D!hѢ��=$"�����38��!��Lf׆`�Ϩ�l��s��K�X�"��n=��d�p��u}���:QJ�}c�y��'�Ϸk5��E9��油��O�D�V�?�y���?�P��:;�j�k>��V�-�L����hI�/��zL҆�g��@��=Z�d�wnߩ�g���'���T���j��!J�j�I*I��u>��<3��#�b��Tt��0�q>=u��m��N:�u�]ux�4h�!4Q(: wF���qF�֛m�g��a�gn�*���M����`�)Qy�,�^kJc�B���>5�k1�y�\؇I�j�3^ݓ~ƾ�)�Ͷ�F�x!�D`_@i 1�(�_W�|��zA%�lE�|�'y"	_~�Q�3��
 �N �fQ>�����?{�Fu�WN�E�7��<3�*�h����xZ��1��_[�Qz�����p�_~��>#/�Yz�?�m��q�]u�]u:�u4��<e�2?#���#��*n+揼�¶GR8�"�"pJ�0]��Q6�L���J��\�Cv4����������+��n0묄V{eK�������I9����;�K5�#��Ce�$��$�G쉎�өj_�X|��of-<�8Y�Rf�-&$QY����P���������+��A믎<�=5�b0���A)����/�B[u�����g� Ǉj�T�Jh����xP&(!Yꢍ"���֝x��Ph>j�GJ<XC*>�M���CGO��� ��F�F1����2FϺ���gTUT��KS!$�eIՒr������G�£
{��QQP�2"�K)lkyb�!�t�����a�B�ZKc}Z���\cz���l��(�8p��O:a��뮧]N��|��ǌ�������(�O|UA!�D�Nt�o�`l!�}�Ң�N����f�f�:l,��gCK6h��)a�m��8�`�=��z�}�1���ѱ2��B�<o��T[%\6�DQߧ������;+=Vv�t�kT���8�mV&b�>:3�!���3FFq�.�*�Β�J�k��%�dH�Rb�ŷ�U���<�h<\�J*��Hwm���ᵯ���<m�$�L&�x�I$�Ğ�I=q&�ԓ�4�M�I$�-��I�a$�M$�|�x�I&�	$�x�I&�M��8�8�a$�I��&�z�e��e6�I�Q���	$�I'�$�$�i&z��$�I��|�O&Ye�Ȓx��"I�z���'���&�|����î��[I�$�ě|�ۮ���]u�_:��_6�m��-�뮙a�]I�I�e$�>L&�8l�L8�m����L'�2�i8�<m�z�$���syÞ��~��<3�g��,G�X%�<`{k��b��}�H���|��L��9�Ė��R�'�s�3*d�PC��OQ<}AMq�!��?	�^ۿH�ީ����
�K.w�g�Y�����{��0aj��G9=�$�0��|�}�{��ww��s����{�UZ�s�wy�{���W9λ��9���]z�8�n��q�]u�0�0��E�BѢ
wM���4Axڞ��6�u�gMx�o��ǽ�M��C��:����ظv�w�$�k:a�������{;�; ���)��8�)^�R�%!���L��sA�1�hC��c����0��4���1~���;F첃A�� �Z�n���b��Fxm��϶_j��w�v�ᾄ����Qg�G+}nI����م>e��m:�q��:��\u����!Ӥ:z/��������+���jv��U��Ӟ^�:�����^^�9�1l�g��5<$W�Ͼ�+ٛ�חe�l�����q���g�,�Т5����P6W�0l8��ca����<x4hcK|pnH2�|�tR�[E<ruYK�i�=	P���Ӕ@�:mC��G��-c"��ϞI��J�A�|��,��ٳ�a��q���u��M�N��x��h��!h��o�pr���R��!��֗�n��["����{;�!z��1=�;O2.�S@����s̻^� &e����nv˷.���e�
�9�����������W6X���;�1!d�l+^��y+~|UA��<����i1�l��/�dy$c�K~b� ߵ��iMf��q$±�v�R��Z�ڷ�w4u(E�,�0`����r�L�y�cA}t�c��6?p:4|5�a��8h}�ݍCy픎p���E3E&��oA����u��D:5��̍N�}���Gh�0K�y���F�������?B:�D�K�vSi�c!�m?̚�d_8H���p?�\��`���AA͘��:��mq�GǏ|u��I��?�u�S���)���4h�R�lm6�ڌ#S~��$b���`�C����p�<qh�hSq�!��r�8*8n�$�v�����~$;��1�e���J�i�l���1֭ԶK%�����d�P�-l!b��j�A�����Ӄ�����=����If��Yj*mѧMS�){5J��W�mMQ�V�{4k>����=5�]˾�of�j
���l�f�6�6��f�O?{�cx�]q�m��u�ӎ$뎺�u��e2��Ǐe�9�~���PO�/I��zx>�73�K6��Q�����.y�����7,��&�#Ŕ��j�<���O�l�-��~�l2�&�H9��JI,��<j坲��眇㥄XȰc,!ᓧ�c�]U;!��Ђ3�m&0ʍ����!�{oR�t:��-�.8$��E���k�nÞ�GC�
����ѣ�d���6�n�ӎ$뎺�u�4x�e�4h��b�.����r�m�*Β���(�T�j6�xa�0Tp����N.��}6�@����i}�]j�f���M�TMt��Vj��6��aÏѵ�*O�f}S���_r������N��ê�N�s�?6t��X|h�8X
ȍ�.$� 5L9�R������ϛڼ�u*�}�b���\&kj�|qQzn��<ul{o�S��O�M�x��T|4�-�t�㧋<t��ζ�q&�u�S���)��H �!� �%��MARD�-��+��7۾����o���B�A_\q:K�"�ƚ��� ҁ�����/���|l�a~�ŭr�-�����&,�����6�b��/c�9Q���x�v�0E�5-.$�@"��?�����in�b����I�tٲ)��*n��
��Gr^K�N���La9�^[m��N���f��f�x�ǧ�"��x�<p�h�}Y�fm�۴Q4�gtc�?|��ts��TQ,�p���/9�iQ[X3G��Uȓ&P���>3{>
!ege��x�o�bg��)䑨��ɩ�0ic��Ψ���mi�s�߁@��a������2���Ƶ�ql颌<��[m�i�m:��Yu����!Ӥ7�~��[|ʨ$����/`�gASI��F�-uL֥[���Lyg�����h�O�=����^���nO67���#�e�Mx�2W)�c��z�=����i���3ƍ�}Ӎ�2#�p�s��k���ּݏm#��ZW����wP�GOÍ�Z�O,]]F.la���F|�t��OQ�.�ˏ㋶R�Y�l��oK�C��L�"n:e�[�����^��L��m��i8�M��04x�e�4h�xpcj�L���N���l8��C"��Tjfͮ�l�Ƒ�o����4�R���8ȡ�vh�ld�ʹ�i!ߛg��=�����$nS���Ɠms���[��S6�����h�ZO�A�w�χa��)\63��.5�(���y�8@�3�>�U��w�.�8��G�Ӫ�$8������p�.�����'q�go&S���m��4�q&�N'�:�e�׌<e�������y�?<+�ϑU���l�Idk�eA}(��C4b�H�[~�G;����-���<��F���V��8�'�t�G�����6Y���΅�Tl<s|drC<��-��C�����`�}�jQ��x�E��-�=ChA�
>�Ll)�<Y͏�GQ�M�:�Q���5��f�F��Q��BH�`���i�TB�;�2J!ղŵ�h����o��u��I$I"I$�oz�$�ĚORm4�Oz�I��4�I�I&�OQ$�a�I&S	$�z�I&�M�N8�8�$�I6�ē��M��m$�)�&Xx�M4�O�I�I$�I=z��I'�$�I$��a�Y|�	=x��I�����ĜO^'M�D��Xz��Xu׮:�.>I'������ԓI:Ӭ�z�m��L�뮺˯uԚI�|�$�>L&��l�L8�m��~�	<z�)$�F�'��"I7xX1��ME+�fW�
�CB��F���?�N!�a�jV�H0��(��vll�IOo2�Ͳ�)L9��M-([v2�Dۖz+�b�K��3���ݟ��
%z�@lP�}O�6b���߽�)e����u~B��0
������ԍ_
��+Z0DFLי�bD���V?1|���*���A!e҂���L�>Li���bZ:䀨�Ɩ�
�Tt�d�hFD���P�2��*�����$��Ө8��w����秜ul[�����f����;|�Y�I��� ����z��珞�'�E�$�K��q�,W2�[pBؙ֖�b�H�\a�r��`�YGP��Q(EAPb���7o�Rg�b+^�nM�&�i���'A4�!�A�o=�~iդ��	k�����?<cu�[B$��E��$i/�I�DFay.j�ՄE�7k~�)ӈ���h_x��t��
j�m}V1jQf&"a���J`�y���v�C5�Z�S�𢝠��nv��|u�9��J��4І.�4Ė��h�j�0�.�;�C����F&�5�3n�^A��n�2� �����n�U�g�[Zm�{I�/nu>g�Nz,bks�zv�W!�u��;0=���m��u�b����؂{s���vi�nw]�~�ȟ���L��y������)nA�]\'�����=iKq�0��v�#+�Z�U��0��k���=�{߽�[����g9�{�wU[��u�g9�{�wU[��u�g9�뮺�l��m��N8�i'���)��^0�^��?�����Tb�`IB�4�&�_̈�H��12H
`�b��J]-d5ّ[o��oKk�&:��!�˝����-���ˤ�]�õ�5Ty��/ķq�Y�X�v�j[[�$���ݑM>9����ǔ��ny�p�Җ�x���{d�p�����\ܗu��ˌp�F�=���7`�Q��g���㭭��\t�8ۮg7H[��.�<ˆWQ�_;3�?!<t[>x��B,�a�ߕPO���ѿ~����F�5�&��0w2#�)H%�մ�����h�9�>��F���Ϡ�ıtR�B��N�K��ϱ������ߖ�ف�k�3�4�C���gQ���!�`�"�EQ��Ҫ�8xӇ9�ђ�O��8L5�ځe�\6v���Q��J#�\4���(�����ib�͐�2��YTՋF���m�C(j��%<=�T 3OI+%�L����1d�ulhyßءբ���`�8}��]#f�my�<�������u�u��m��N8�i'���)��^0�^���im�u�E�z�l��L6iCz��xg4aN����q�{�6uCAa��x��t�KF��\^rIQPݭ�ik���I���+H�3Gw�"~�Y�/�*�|�7���5"r�$���,6�q��u��tB�����LӝO�gǎ����-�n�un[��������Q��9<i��:M�[o1��r��D"�Oqܫ\6P��4p�4t��u��6�q:����!e�t�m���is���3�^Y�\���ە*��uw�tn�v���6!
�$���d��Q�|�'~oP��Sm*:��|Q��+�n]�@�H.ݿn>BhB�֯?��z|.���Ç!�k*�Nԡ֌\\)5þoj�B��c1{��Y�UIG��3WS�p�2�q��9+/i�*A��n4��CԨ��ҳ��_�g���8�o��qěI8�ΰ�/|�,�t����r��6�3�����g�:|h�]4��h���~,��lzI���Kmdd�E��jV��\�|A��0PW�"���!�]�G;���D�P�S�*��&�G�6p��gM|iC�g����f�70Ö��xq�D,�ƀ�m��4�̌��((g�t�K͍C-�v�Sm��3w�����]L�����m��L�I����0f �,�~���cd�����%������N�٣C���l�$pL_W*"�kL��۫v��6k �E�l'g|�;�SM��r[�qi+���6p���f�攱fa����m�#	��,��w^�	fi.g��k��⪂z{�o��O?}|�P�ScuV��������	�=�x����ϲ$�@��)4��{e�z���J(6� |���	߇��e�4��v+�]�)�I=
<"��>-t�f�C@σ�v�qܻR�4E���.�������A�����7Q�Lo:�!�c�x(a`�k��m}�	+i<����+�Ë�D�&�c��UR����i���F�
��c3i���K�x�F_��0v������l��|��o�e�jN�%T1�e֝|�4�i��u�S�$��ǎ�0��h�,d,��r�7�ޛm�0�#ꁡ���W{��N�6Y��6��9��S���k�t��7�A7C��.<0�	���/N�>-�^��0Xh4Vݏ���xl��ȈN|~OI:k��H����Y�&,�r/��ۚ��G�GŨYP!a֛G�(��m��OC�Ѩv캮lo�c��uN�1�x��K�������e��h ��ҏ?�}t�=$�i��q�S�&�I��a�����/lcK���R�nZ�g'#�۝��UD�=���)��^:cu$gXl�(�_[��12�!�����#�aG�-iiq$�d\9C��(o~�t��x�F��I��N	?(R�Bdӫoh�m�=����n�í�n��w`i���E�F�3��.R�1��o��0��BA����ރF�i�Q����t���Ç�6����k�������e�a�m:�m��e8�i$�N�î�L$1�|x��x|E�R��w����y��k���)X޶�?�� V�ޝC��ͫ i��u
C���;�KVF�ڗ�OZL���,�M#K�yc"�d����*E*NުJ���Ã4DsE��氣��7$q��e(~(OƸߍ^�ɜ������(�k�2�O4l�Չ^Rg J��.�/�S�բl�\�_����|��QD�� T�E�e:[�֛m�]e8�i$�N�çH&�>λ�p�ֽ�o;���-�ԗ��{�m����e�d�I�ir3D8�M?��F��D����
���bBu��l�s���2AՆ[[�x�'1HJd �*��I ���q�GGR��̴����M](i�]�жV]f�F�Y4������򅍅J�0����=Y���-*�g�/v�T�u�,����.�����������>�H����!G�z�a��x����|�C�3�:t�������-�� ێr8���è!��+\��^P�˥� w��+��Tvu��-m�̔~+M�x8CF*����.}�4ߎ�|���ᝋG��,���8p���8�i$�N�ì�a�>z�fvQ>i��3~P���3�c3�w���+�e9
�U�<Ig��t�@Λ2KE�1t~7�.\�tY�à͋P՜��Q����1��i=6�:s��|t־��� ��������&��'�
H�0��)�f�t�<@R��o߇�^6i|R��_,fΪ4Q�����P�_Qg�Ӧ�eu���Gq�F�diE�ul����s�r3�e)3J�)l���7f͞�4�u��IH�I$�z��I=m&�|�M0�I>e$�8�I�^8�e$�$�$I8�x�O�I>e$�I6�	�q�N0�I'x�x��M$�oRM��a"L$�$�$�2�O�$�e$��z�$��L��|�2�/Ra6��#��OSק�$z�a6�֝a��:�����.=I'������ԒN&�:��m���뮺��^��I8�x�I�L�N0�z�d�aƓo���I�ԙI&�6�$����<�W��˫@��l.�7b�i�N��H�3҅[�%�T�ZcI�	>Q�/Tt�4��ب�m3��@�/��'ܾG�/6H9�X<���@�v����[@ s_2=�����ת� ɇu4��1���}E���8�X-�ks݂����S��o��4͸�"yu*D�b� ��*��b�Q���?
E0��"c�z��C���V����>ӞZi
���f|��^u�k�{��*���;�k9�{���UU�s��3���{�UU�s��3���_:뭶�M�믓�&�Iĝ:��0���5�m��2��HQ���8u|��E�ԟB�h�Z/m�*8p����Ϙ賝�钮˶�H���E��y�&��m��1�m�S7$%]�$�KFZ�����辯ߣ�}0�uɞ�MC�M0����gM�c��+�Ϫ�ʺ���O�o����oeXtaE{��oc������>�����4������af�W)ԕ��Q���B�z�6=��a�_Ͷ�m��'M$��:u���Qe,��[�m����Y�M8�ag��B�s��,=<�����;M��XMyC�ؖ\�b�6=#gw]���F^��,)r�P�n�6����aR
4J�4-]�sm��I��m:�L-����hts7$������F��r��fՌ[>;}M����:Xt>4r�zͣ�e��߹��ǧ�v�|4�s��I�������9�&^8�u��m��8�i<x��ǌ4A�2�,���!MR�O�ݝ�'_����zSh�!{��G����� ��p�g�H�yș2MM�Q��'g�i�6܍��켍�3�Vr!QM!18:��i��z�'c�YH��uR�w5[Bna�%�Ņ3��Xm���(���%�b�/��wi���\��hd����z;�>�!���=��B+�E/�	ѥ�	KqVv���zH�5����[�?��m��b�˘Μ6�c�y���L�fŞ:X�+9|P�[�g��3�����:�n��ml��Ps͡�Qͣ���~!�&aK��	 � �I�1��0��ZL'[�T�pxt�Ro��C^T}�m�t���
�Ԏʦgs$������fh{� �_㋇L��Y�I|�G�
8Bƶދ-��N�C��4a��Fx᳇�|�q4�I'N��X|��Ӿ\�h��EM-S�m��c�Ka���*<X��3f��a�� �}�ϢٞVik:7�� i}㉖zA��Q*��ejܖl���&���p�Y
=V�0��C�U��$�$-��SY75�i�n��@(�qxg��[-u�c��u�c�CD$6l:�E�G�n��f#�q�������`М5��1���+F���gN>8l�����8�i$�N��,0���Oxz��ǈ�������Ό�GO�tX|(�ɩ)�p��
�l9>(6��0�l��A��E�=|�B��t��]ߍu��Rf�5��Wi.���v��V�?�����)x�C���B#Ş,vvʕ���gK�~]6�Y`Φ�ͳH��ѯ2S�TC�f.й־\}���Oq�7!RA��l-q(�u�=��x�u����i���I$�u�a�X|�����Q*��"�j�$-���j��m��{gW�����43Aю͘Y�p�H~���r����N���h��6��0jFZIb]�^{&Ҍ!񣦾�3S�FŻ�$�量�U���!L{
M1=�a�o���ai}����<G�OjUV�N	�,�E�N�[M-��A������$p�b�dL�}�TJr{ގh���^�A�-��ԍ}�1�OPB�ޘF!bţ���[>!��Lm��u���I8�N��L0(" bi0�8rq�$���hy�ٻ�wQ�[I&q�E��Ze,�PJ�!�"q�h$ԔC);Q(�^�jB׮�t��It�4 �l�e��W�æ�͖;���&v�����Ys9��T?W�u�ڄ�%��F��q��!�ܭ�HG卷��X�B߹n���R)�x��o���`�L#�����j�n�Y�o��aA��3e�A���M5el���(��57f����#E�@�Y��(Dz6�y���D�p2��Q��6h���UI*���H���G�..<ya�D�ڼd��g�A���}��c~��?�-�vG���oKׁ�-.���Ҵ��|t����f����_���}��y��l��<p�m���M$�I:�0�,�(��
���*���:�ዣql�vލ�Z�����T�}gü��S��A�G"2x��˦�3t��_��'R��ꤞC9ڃr�O�:��o�n1��(�BE��Q��;�.�Vph���ɝ�m�'h+5��.֩tX��׿$+SU8�
i=�P�ߏ�p�p�ƈƮ�S����D;n�,���B�T���U$M����B1x���I�u�/��m��OS�&�q$�ΰ�2�篞����9g5%-rV��������U��%	XwV�f��%���q���G��U�J�)�#�TD���UO�y�p�zbkc�D�8c}6�|6�iRg�m���2�a�G$������aG�+(5G����r^�gN�����z2/y�Zˤ�v�v�R�/�����>J���~����l�BF���]Ŵ�`���x:p�Ϩp�E6�o���R�kDK�l���A�;���ϟ�x�,e<q�\e��m��S�&�q$�u��a�=|���S�(�<�/I�����w��1�i��(�ϠhޛT3�
5�E����XM.Ѳ�7]$lk�nY��6���3�Lh�m�i�=;��'����3��Ah�(��n4E��8�a���-���i�Ca���R[��eN��0���p���F`�g�م��|l�c䍧8lT�2Iţ��=��%Q��gN@��ųƏ�}����+�;[;��4�w�'N==����~���4���QUTkf��q��7�~��g��7l�Mm-���gN���<���ۺ�"�Bz��/��LZ�Iք(�Kd�!�8E�[D�dDDY���"h���E����m[h�h��D�dM��"Ȳ"&�"DD[ȑdM"h�,����4B&DDE�DY��Ț-�"�&�E�"-��B,��E�D[E��mdDM"h�&�h������4[DE�D[Y��DHZ$$D[[h�h�h������D�m""�$M-���DE��"�YDD�2$Mm��h�,�DE�mm�B"-�""�"&���D�dDH�-�h����E�4M�mm���h����""-`�$Z(�dH���-�"h�D[[h���4H���"��DDZ"$D[D�"kmdDD[D��""h�mb!�"""�"&��DD�dDH���d[[h��E�M�""-��B",���Ȉ�dM���<��dDYE�DD[D[h�"""�&��h��mm&DDE����4DZ"",���E����"X�"Im"��X�-�H��$Y���&��$Ki,�,�D�X�,�"�d�$KiK$HY�&�,�"Y"D���	4�[H�,�&��h�[I��$�K$�h�Ki$K$��[K,�Iĉ�$K,�H�,�"Y"D�k$I"ZD�	,�,�"Y"D�D�5��$K$�$��4�H�D�[H�Y$��I�4��;u�D�D�D�D�E�%�"�i2D�5�$Ki$��ik$H�I"D��B�d�d��I[i-$�ɤ����E����,�Ii$�Y,�-�dD�RKD��V�m"D��-�iki4�"M-�H��,ݷ��%�il�Kik5�H�,�K$$%�h��$Ki	m&�I���il�$Kiĉb�m"Y&�Ki4�m!f�M-�$��4�m&�X�"Y-��%����4�Z$�"[�KD�E�[kDKE����Y��,�-$�mf�ȴ�id�X�H���ĚIdZ�$��D�d�Ȳ�Ii$��,��֒-$�kY�ZD�d�d�,֑$��ZIm-$8�8KI"ZI%�K,�YRIXZIi$����E��ȚY"��$KI����i�JM,�D��E��KH��D��4��$K$��$Kk4�d�d�%��e�%�%�ĉd�d��ͥ�%�%�Kie����g6Y���[d�a��ƶ[�����q!ŉif�V�͜�1��2����kd٭���ckd٭�Xp5��B�ж�	�cB�B�B�!cC��C!�ͱ�l!6��[2̇��m��!f!m���d'��5��ŎCsA!BB�"�n �!���6�B�-	!,94"CY	B!�:�u�k#H�Mbk&�96�5�M5����&��4�.q�h��:��&�D֚Zi5�K�p��I��d֍&��72bɤ֚F��q��4M&��L�ɢh��i��i4&��5��hFZi4�Zi�Zi4�Zi�"k&�i5��M&���M5�D�ki�5�D�d�Md�i���&�h��2&���ɭ�����M5�)�i���֚Zh�Mm4&�k#-������ki��ɦ�h�&���i��i����k#&��ki��ɢki���Dd�m4Md�ki�k&����5�D�M[M4�2�i5��i5�Z5��2��4Mbi��������2i���i��4���5��#&�&�4Md�M4��D�[(ki��ɦ�i��i���h���M&���&��5�d�Y4M4�ɢki�4Mm4��M4�[M	��&��ё4&�����4�[M4�FD�Ml�&���i���i�&���5�К�h�i�Mb2&��i��i���h�&���DH�&�E�N�p�LY�h�[DȱD�m2�&DE�&���"-�bbh��&�D�m,LB-E�h����-�"ȑ4YB�""-��4[L։�"�"-�e���-�"h�5�KmmD�dDZ"��$-Bȑ"�m"E�в"D�Gnm���d$Y-��D���%��F�[�"E�Bhֶ�BE	D��--�"ѭm���!h�Ő�-	��d,�D�D���$YDB�"��[D���4Z&�։�E�dDY[kB"�""-E�[kh�$Z$,�-���E�DBȖŢD�DE�h�Ym�&�D"�4DZ&��։�Ț"-DD���:��d$Y&�-�DE�b$D[D�,�Ț""�4[E���"-�"Ȉ�",��E�"Ȉ����"�Ȉ��""�"-E�m"Ȉ�&�"��H�-�"�"&���,��""Ȉ�����B�DB"&DD���dDX�dDMm����h�&�h���=r�S=m�.��y5�o�n�mb�PF����4~�l6Zlm��٘�T�y��sݗ�����������~ߣ==��g��>N�[��?C�������?s�����zsvh�|�����8�������g����o����b�7_�k�|Q���wiE����u$h?��g�{��q�3a�G�3��=��o���F�M��f� ��o�!�6�mȄ�[�����}-�ݟ�y�}L1x7�e�l����3�������|^���o�֝�Y�O���<��l̈́}���<��$x�Ώ��m�}^8���6�o���Ɏ�mgZϯ<�����g3����]��7>�<�x�򏥟�|1ߞ���u�|�;�Եeo���g��{~�3��p�lͷ8�9tͷ�d�lu,f����1��gVc=Z3c���V����[l�f�\6O造A@a��!�"PM���}�ǻ��������=�ݽ�c�Z6fm䁛��P���&
�&lg&6�C�t�?y�}��}�՞y���o{�fE���������{G�7��cG8�z;�-�ao������_<�m���}M�O'C߿������y�soO�~����[w=�����޽��ַ�����>��v?����e��=���o�ߨ�����߉������&�#fl>8���5������c�����z=OF�>���g6{��ߍ�ٰ���3a��Ϳ~e������4�踺�g���W�����n�o_G��Ξe��<a����l�;����Ee�{�9�=�M�gG���m�6#GC��>M���m�pL6.���� �?̈�	~��B�H:#H9j/���S(�����zWx�g�o6�3a͏��_��|?����/�����l͇�u���~��G�-�6�=��L}'�?��=}��ރ���n�gC=O՟'\/��k}n�|����o�o�#n}y�O���]�7�������6f���=��ő6߇��~��6�w>�����Ϳ�z6ߤ���g��g�����{���f||��)��֒}�����"ݖ����f������}���?O�o�۞����v7�ӻ:}�����ӹ�7^��I��l̈́߮�������퓜ϧ>�o{���;������7��=�=���g�L}1N<�;��7MOW�Vy�{���-� �c[?-����������#��ɼ��{^�]� �����k���Kg�f��@_�?p5�;��}��fV��8pn�4m��������B�H�
c��