BZh91AY&SY0�dL��߀`qc���"� ����bB�      �*�QB��@cRh��@6�-e�mEUق�(�(
PEh���P(�m�4I�d(UV���)"�ۺ\n�_p�:UR�j֦�٦�Q�kP��[hcKSL{�樠faYe!�"H6�3amm�l�[4���֫��jV�@Km�ݦ�
R��BG�t�[L��j�7q���hm47 �s`֤VV�X%�lU5�e�E)mX�mk6���{�ml�I5f�h�J�-H�e1J��,��5C^p�(�
��   .�g��hV��4��N�� t�έ`U�� uWF��,\�GYE]�Z횪c�
�k]:m�꺭i�M�m���4-����  <��Mծ�:P�kAu;������JPu��P N��� ��� ��P]r�Ei�1�� Au��W��t j���L��f��5��[m�3"x  Ż��)��yǼ �{l��@����^� =�W��
	���yҀ �W������{�4%CF��� h�v]�  �R�b�KkfTkejV��Yo  m��e*��g��	W���)C�A�,+��L�ָ
t��mSMf5P�MҀ�)Wu��

wu@$
w:�hP����Ja�ki� ��*���7Nt �M�q�� �4 U�[p:t�
]��lh+M��V�Ѣ�]wCCJ�*��%��T�;��m��������m��5� �x =]��W 4:	˳��Zik����*w:��W:q�3u�æ� ����@;E�xP��Zj�x�@�yDm�@ЋY�F�R �� -��y� ��N*�����p�R���� *r�Ҁ�� ι��l� s[����45Ѯ���-+2K1���5�mRͳ� ��ttL0��]k��E;7  .vp uˍP�`� �\ 6�;� ��Y�C�F�I��
�K[[R�[5���� ne�Q@�w@ցuq��� ��p �F  ۣ������8n]��4�]ƁU�s��KZ6�0�ʬ�3E�ko   f�P ǧ��Ϋ �n�� Ց�(s�n  �U���˜Q�wGqT
    �   � ʔ��0i��  �LA�{A�R��0h0#	�&�
J��     ��$�RC &� L ���A����@*�2   4  %D6�2��M=F��d�i��1=OD��9�=12�5�莗�y����RFk�le�n|���םǿ�=\���航������UEAS� �
������:UE�=��������?��������-UW�ETW�T�T��
��G��/��?�)��L�fS0���&a3�&L�f2��&a3	�\���L�ds)��f29�e����S29��!���fS2��̦a3	��e�L�fS0����a3	�L0��̦`s	�L�fS2��d̦e3	��fS0���&e33�L��29��&a3)�f�fS2���&e3!�L�f���S2�̦e3)�L�f&2���&e3)�L�fS2&e3)���2��̮`��fC0��&d3)��fC2L�̆d3	�L�fS0��͘	��&a3	��fC0��c2LL�ĕa3!��fC0��a�3)�@s �dQ̠9�2�Eʉ�RaE�
��0��T�s�d̀�����s `̪��G0�Pȋ�As ��Y�G2�fE��s
�`�9�\��#�s�`̠��G0� \��D�s�eA̢9�2�Pȣ�s*�a�
.a̢�� �"e@3 .e̂��&E�#�s .e̈��2��A\Ȅ¡�Qs
.d 3 �a̨�� ̀�T	�2��\«�Us�s�3 �*.`3��Us �a 3��f 3 �� ��\��W0�s��L��09��&d3	�s�f2��&d3	��fC0�	�̆`3)��f2�̦a�	��fC0���.ds#�f`3#��fG2���&`3)�L�fS0��̦e3��L��29��ds�s�f2���&`s)�LÝu_���s�#�J���&�\?�ݢ����/v�)`�F�ͼ�-��$b˲2��ݝƪ�Mu6���1p�)�^��(3��c�ܑT�*>v�W�'E�p���Y��*ӈ�F���f��۵�RyfPu��Zԝ�J]l�.L�Z���!�$Q��"Q��x�p����Vn��URwX���[�-f9*^�HV:��*�̈́I�kb1�p�K۽��1"��gec{��5n8\Ků2�l�u��?�w�YW�i&�9$"{nÂdn�MWol�jMn�2+cF�Zl���5�P%J���m�vqYA-Ql�fZV�7�	�1Ҽ7�4�uv�:��[%��̵����FRv���5@�[�rId�$¬��������he�/r���lb&����,����[j$��{��	V����f��B�TM�m�+u4��3q���'LvZ8�5+���b��v�h:��m�3t��Źf�Q�.��YVn��Yf=��cQ,Y�6�F�v�nC�T�L�Nf ��l�e%��Ǘ�e���h4�Y�ZݡV�Y�!d��H��{�^K��a[K1;�747�	4-!�3&���b�7��qR�T�j�-<�!���L���+!Y4��JɄ��5*��Z�c�#NM�3�V�����b�M�%VR��]��7Kq����Y��Y�B\د5:��4j�uX���$!�7�ɰ�1�-j�x��(�q3�Um+&j{&�&��(��i��
&���F���{��L
w50[�Z��e�gU����`x�c��0U��uL~ڷt����Ƃ�ظB�w�+X�%�����jQ��䳙{&�c��ïU�*]V���H�B��e�;�&H�v.�5M����λ�6-�^al+�FZP�c-�2U��0�r����û�.�mD[zU�K?�i�������.��'��T�kj/kx	2�%G/V�wJ�i���;U[0`��7���%���44��l*w�۵x�]R�dҮ��5�X�Ô�`��4Q��:g�Ж�T�Ǵw�Tvr�%�ݹ�w%���{=[�M�ޢC�ހ�u��AM�x�x��gq��N�M��n8*�t�j��h*�~̼��a���`����l������z p������J�)���vj�&̅;a���Op�z��sV�ĝ��t�Y,Q�LT�OU#��4��n����mY���p�V;h����[h�����j�T���e��	��$�ו�C{��a���Ɂ�;�(<�Vh�ŷ�M�#��%�meY!�F��'-��ݕ2oj�J�3BB�CԮb��n�6&*8	w�U� ���]��Cm�74�6����	�w�r�t
�K3	70�gf5aZѶ�X.sI	��V�N\0���hJһ��1nB$Vn^��&�/�j7zn�n�i̷V�m�w�[�����u�5�=5;GYt�𵛖�[��f�X�M�S�@�7%Ӭ�JC,E5�`�Y��O)뢣�-1��^d!
RI�w B]�RLOXJ�Hۼ���D�"�a��h�*S�Wz
zI�^A��.؋M!ow2��W`�y�ҥl:l�m��2�N�*Tڴ�Ӓ��i��Qj^^�&ݭ"�"TV��a������z���T���i���$��Ѹ�v��CCjF�!�DY�)%Q*�nS��b���c���Ij��ݺ�"�R�S��[�Gv�zj��^��v�^����(T��Df�3���[�+4�q����
�i-��(5��w�*.b�ݗW{��5���#YJh�wV�U���$7P4-̱�g/0k�v�X W��	6٢�ۛy*V74�AT���5��,�K�kR6�XZ�ca(]�5u(�Gu�o��X& ���;͖�0ɸ��hy���6�z��le��$�5X���p��[&�������n��Q:^e\���h`�,��+�9�����L,5n�NnQ�ך�p���^�co��2݊�w��!H�7o)ԡK��t����l�Z��	�*��5����K�Bh2"k%�x�������n9�Rݫe,@,�e�0��TF�Yu�pɎ�m�]���@����,t��{�Z�y�cV;t�4X���Y��.�ƍ֨]�فRne]Z��P��o	����\@�@�N���X.��f��H�T�֢��\�5�8��6��[�l����,�y������^�n �u����
u�t��B�of8v�,��yIܴ����C3
���'YE�bK�����!�PT&��ʚ:��g6����!F�Յ+V2%sc�@�և�����Vᚴ�Y���C2%Y{�'�{�ۭ��n�wa2Z��$6�f��l���M�L�{��n���-4�-*�c$�m^�'���[����Th�6@b9wl�p�Lbv�a�H�Vus߲ɢ-3kmeN\�FZGT4��wAˍV��5���`Km�i�TL;`PÙ���W����i.���e�y���Q��|�Q�mk�u|��a��!�z���樉0i���TF�حX��v�����X��[D=a�	�QI�rkv��J�l��Q��;ԬSH<�ٙ��kRTFn�w/����ض�,�Ga��b�h��6\�g��O+��<���/�B?2$�v�f;�,*.fjlۄ]Z�(4�[����Af�O`m[�;[�O�Р�qFN�@�4u�5�8c0����2��9�M������(DE���Ĭ]�X0_�[̦�5��&�,��%ia(ci�[�]o���S��F��͚P��su�U�5�9Y�F��터�pX�T�Z��,yX1R�^���`��k��%EB�*�)4\U�Ϥ6wK�÷A �SE֝Ć���v�A���,j��t�D�:k2Pa��ɂm3��0���d�W7��4��-0��j'f0Y6!à�Y3i�r�%e���j"�r���3l��\�opzQ�!7(A����sjЧ���%��֢��̺ǔ0�7u �-�7e��1nc'[&i��v�@4��ow2�����)��L������ǭ�CZ:4R ��J^{����"�L�Z����8.��YEK9����"y
��sh\�{�f􅂱�K�.i4�e�y�U��lm�W�c�i������ۇ����Yq&��hPVP̤栭<7�#��r�e	�flFQ�#��
�ZYd ;�Cl��=��"�$�wj�R�Ȫ��0fM���ܘ`X��*G��r�d�1[y�j�:}��^�ٶ\��h$i���G2� 8˫��-`�ױsM��~��j�I0�k��(2q!��J�`��T��YR�+4��i��P���e���Ե��e�S)-�l��eaˠͼ1��A�bW�M�;��X�e���m
�0\C*��Y,��91����{�Q�Jj2��[�vL�a[���	�B`f-���*�
6ʹv !R(ĩwq�ղu�I�KL$�XCT�sB�,�j��i�b���u��/��B��4[V�����V+��6�ǥ��
�'X*(�l���n��H�z�Kce7k	�^R�K3dX�b:w���`ʸ�v�j*�f����U���l�DPaSf�˭x6m���+&V�(���+˰)����u0��V��n0���
L(�����^��R��V<��oeeA 9Q���ˊ�N���n���!�!V�M�(k�eQ��ł�b����5����f��%=�X�f6�S�V�.4\�%�6��%��R��u.T;jf�(ʶ�4U'�3n�"C;�h�و]��%�_���E��[��^�ܬ�k6��y�0�S* ��*7�0m�F����d�I��f	�٬r)ZU�2��D%]�F����iTm���<̐BLU��^ÏJ;��������"�x�w�k"'�Ѣ
+��R��䬷�+�0�"T,���QT�N�f�
#.�^�:���j��(���2��cc:�b���x�A`;���j����M�{����$Xs-�M\�6U�B�޲�)5�ͫ��l�l[��H:&�Z>�MY�U����Qw*�A�2`��m�gl�I�9MZU�6Y�6��`�<���ˑ����@�Z�f\�۔��ri�����2
�e�h�n�]݊��ڙo�v��)�Ԣ2k-�'%@`n�b5�nk��H1�wz�kJ՜�T�/0!���I��\�i}�RV����o�F˖�i߰����Y��b�	�H�<���(X��.�Z�". I�SKû�E�6�������|�ڽV���I@	�U3�*q�5�D�]J��<I0݋-k¢c�2��b�&�7.�嬄Bt�+aI+���E	/���ɮqnѧ��E���Η��弔�����B���s�ł�Rİ�	��5^���Č8�G��y4:��̽�qY-��pL��
&�$Y{�&Q��j	�ɖέ�D��s�,9c?���'y���+ssvv���yv��͉ǌPȓơ�7����[�/т6���9ZsaIl��Y��u�T�j1{OM�1�֪[�/w7V�u�F�����#n�n�.���)9n���L���$�goEC�V����Sg/LӬ�C�Q�Ȗ�e��M�9��n���k/f`Ӿ�n�E���QX-�G(����d����2�bP�[Y�r�\��v�mč����[�	��f@��EM��t���KFQ�OZ�\�n�r�$�M�kQ�˩5�K�����e�Iɷ6�E���V��Vi���"�:5���j�
�^�jVHRz+E,͚����B�r���l���AG���f�U1���GM��G��l����*K�P��t7|n��*��#����Z9�Y	˦�@�Q��Z�'�7���Xn��B�3E3s�c`f؈�4\�z�;�d�ۚU�C�u���&�ވ5mBt�S�(H^����"$�Z�QdÏ-m�J��s`tٸ�ҕn$�Ļ��q��7+�	�Mn�wb��h7Z�[�U���]���e�a�Třj+l	@�a�]cv��=m=�x�=T/�V���8K��2ڹ&м�	J���Ùf�|i��v���ur�g5&X�5�h�ɗj�uwj��b����ܥ���n.x�n��V�lL��*Ւ��'(��z���.�ʕ�0Okxs
7r-��![swP��-skaN�IP�����0և(f*�$)�_��Q8��b�f��嘁�2J&ȧ��5�lv�m�9��J��k�(*��)&QH[RnAe3QnC�)+	��h��a�2���7-�wQ"���6�%�MI��,�l+u�4�;�.'2�v�ǒiy3l�P�x��X]�m-�{���\�[F녎|�eQ)���m���a%,[H��N��&
W�=v*^����b���C^�W��
)�ܳcPX���pˬ���ue�f�Ŵ6�fܼtұv�-�/Tt@���Hږv�Q���Y[r�p�2�#(��SSP/kM��Wo|�[m��5��$�sW���O*�p,t^�9�6ȳ@piN
����)���;{NElǶr�T�н��MD��,̸
)�.��#�/(,�����[XY�7&�7P�Y�5n�a�֕Ȯ��	�;̗��xv	N�dw�rYd\9��3"K�|;^�Q�{&�֝�^m�ɐ����aF�����I�ȍ�B"�KxS90�v�K12]�0��B3���d5spVi`J�@��n����iZN���.A�FevdQL�E^@Bv�J���
Yn�
%��em޽ц�1V6	�$b�R5�n��L��L�ۻ�3u9�#VN�����Ѓf&��n�ָ��$��F����J�1)�x�w5�y~�("I�x�,y��#*��:ope��e�fB/&�ۿi T��95�YVc��z���Ӱ�I��%�ۭ�w/M7��(n���z�.Av-Q��J�n�kV�*�e����E[�ǭ�����[��$�y�(��'���sq��ۦ�f��]���aع�3qh��Ԝ3�xƊN�ڊ�փu�q9�Z
c~�Z�Y��u$������cg�66k�Lb;���r�rm�?�,baJ5��(0'�pmk۽Kj)z�^�I$��Ź���v,S�M��#�7�xF4�D4��Fٓ6/E�v��2�{Y�K8sw �8�[ؕiym+���p7�F��Z���*ݼ�Z������xA�3(m��lܘ-^ެ���֧6e�U����I�q���x�טZ��oc52�%r��n�rR�>�.���T6ax��G+p=�����[����e2Q��iǴe��{(�пJ:4�l��7p�Kr��A��i�՛�2�r�'Sɇ�`��݁V� ��Ul��c`r=�pp[C@y#�6�~��q�����c@�.��v
bM(��L�T�X�!�z�7�!|'Z�WNy ��,u�|�~"H�v��� �o�լ�apD�5��l�6L�".KL�0=�S�P�W�:����-���C�!�4,)��i�^U�������B��M���T6+XO4�h�.�0�-̬�L�]2����AZk�%H��9&>+$-��<J⡉�b��yb���H�}����z�X1S\qlG��
$�xle@�B�ؽ6���,c���k٥5��ȶ��嚉��:/%v�n/�;�문`Tw)��)b]�R��aKK�:��a,��2�aÊ��{0�97b9W��Al��5�7P�ﲦo������u��=��ѰDiY)5z��-ۮc�f�ʸ[�2����U��{X
�� `��}�zv�1�KΩ�$;��͚��bh���� M�q�x4��n�cD��`��n��s�?����{��?ن�������K��MC��3����_��s8ҝ�!�I�8�	���E*�\������Wfݘ�rڲ=׈N	J� �ˤ����.f���v��N���.����>N��A!�,kZ��ܠS3��5_h��ғxR��K�o5'k�*f��/�(�n	}ל�d�jl�P�*m!C)cV�7���ƴ[��C7A�]�rղ�����$�e��jVƩ)ܜf�ְ�HU�*�0v��I���h�L�1��-so,�Z��,��Wu^Uk�O���I�x0˪�YF�'d�%n�Μ��>ٖ7,g1��;@�#�lʹ��$��7ĝ��3MP���Y!���V2D�{�L��YV���8p�J��ȶ0�����
���G5��'�fr2nvu���q���'s"�K9V+лB�ީ���˩ZV�	��iv�8u�:ժ�̙d��z�4����ٸ�gk��i;�������m�����(�\�oc�Gj�`�4p٠�%�q[j�TE��:it���n`�*:k_r���.Tt2�UR��m�8�	v��e.�+��-9��e��z�N����n�>����"z���HǺ�'2�e������q�@��'ol)5����y�I=U
�ameM��Y�I.��X�D?�t�V�Ϙ���\��u7@���thD�u�������Ÿ\;�.�X'k�b� �+�m��T(G+�u�a&��%��׉U�ٮ��𳸛/%�yV�B�K�D^�����Kv���Țfλ6����=Vq���}}Cg	l�N�8��u�'�9�D�����*Xt(���F�a����򪸼��.ö��֘�;q�!�(�O�D,C�]��5���j�P����� ��O.T#<.gR65-���7�EI\4�[{je����E��m`x'C]۵b�}؇%L����	�oj�Mf�teVo��nZ��79����Ǯ����NZY¦�V�cP�}ᓗef��r��v]�Ŵ/`h㽱9J�f��a*x"ne�C��T��a����\�҇x��7a{+/-��gjv��8]�|��hR\��`ޭUB9�����:ʽ���r�[A3*�`�|;���j�k9!����x������LV!z[��(ը����Y���%���Z͑w�8+�#N���I[/�<;�N��V���|9�I�^�mk�a�F�VlN�"�;J9��۝�s�F���*���'/�/i��x�)�	Cӝ;�	�<Xr��pz�Ū��wf�*%�QZ*,�v�n��o<�B��=��2}$�l'ݶ� 1����.�Im9�P�g!u�(zǈ7�Y>T��5��$x>V��t±FA�4�2��Sm�Q�����+�α����N¢������Ҿss"����w�R���[�;���,k��l�@��;����Kn�'���H��tF���ɖ�d������.d��8g5&�'%K{.̘�Ъ�ը�nfۮ�������QA�c2�9qU��8�K�/.��Ik�XMc�k.%k��r�G��d�:)�V�Vd�x/�h�ܘ�eAl˛���R������97/��'S* ��C�T�B(,��F�O�t{0^�<������ʀ�ӛw5\n��+�����6� �L�Q�r��SU�Y�s��j�V�f	]�L�[�v��o/Fkeq
;d���w��"���7�V��C��y�W0���q��9��B��\!����n��}��f��Ya6��T�6��LQӆ7�xU�i�W �ݔOQ�!��3�Lө��cd�CY�t���=�ݹ�<b|� _�QǺ҉��R����+0�5��,�7d���h"vUjyb5J��W����YV�S˪H5J���K�+��4G�G��T�]s�[��`�e�٣!H�;�^'%�X-;��0\��zĈ�Ħd�K*w8��/+tdz8�{J�42��f�<̙��(
�y}%�=I>a��2�^���D��xc2�`%�<z�b��]��&�VV�A�#�=z1�|��m�'��ۣp��YI[�=V�Pb���q�����R���J�q��A��puB����|��,>�'So��|���c���\u�7*G����i�Q�꣹�u���רv2�/�pu֑Z��癷d�:K���dP����!}GT��u�A^�h������1sm��B�h�;�M���S��hlg�7Cf�(����s���lE���f�Zf��i]�V�'��t�e	s�	Ty%#�6j��ĳ��8�N#&���J���%臠`�	��� �����ҁ��i����+U��·s�CF]*4�s���d�ۥЇ�2����p�L5�N�P�Ut�h��q�4�A�h�-����2i&�ۺӁ7)`��:���t�+�_ofr�ˇ�Q7��8�듛��\���Y�d��F��8)� j�=�b�L�t]�U�\�м�֮��#oD$^3D�K������Z�,�:yY��I�E<�j1>��]ot$���#�8��,�Q����W�m]�\�o:��q!����:�hx_$A6�GU�&uZ}��D;\T0\�v)�T�9�w�3��r�ӽ���*b����>=)�f*�tn��åu�昒��O�X���;���o-�C0��v.s�̇&�[3a2� L���I�����9��W��n�CȉV�|Q�DŹA.D��`�å��#�]����V���i���+^4�e�UJ�W(��N�{
MU�
9M-C�s另�#'<Dq��j��ٖ�7��V&/i@�ڄ��ˎ7�ě[��w:��i[�4�X�l��a;
��	Ǡ=�Q���h��1N^��	�Ḧ�v��D��ݗzU��Sw1C����v(Ν�X6�\�n�in�`���Ƶ�d��qʆ�	Lޭd�+�<�bX�v��|�=�x9��g(�j'1�;sD�T�O!x�0v�۸�JR6;7��ă��yx���e�
�L)ki�<�l�����X�>�����Q����K���&��ma�i�!�e�m����s��zr9���(�p���(:�f�:0HJ&��j�g�oO�xy:!��҈��b��[��K�wF���`*k�L����/���0�sH��uͭh�L��K��q�0�Xk.ZJ���ᖤ��Mm̜�c�,�n����:'���`�0���dn��p�st�C:�TI4��Y(Y5��p�g7=ng\�R)��⹔��Z������enY�v��hdS����,�ur��ґbes��u�{�jX�ynƢ!�s���S�O{9g"ꆜ��U��;��N���t��ڮ[ξ��5��i(���I.'���k4��8:�r�=��{BZ�J���V��eu�8]����xY�|. ��\�vΎ�kmn�3Z"�vAS��NX-�x��/��38_7F�~�i4��M��'�oϯ'ז��C�>f�b���;����ޑ<�Vw$	�)���\�(x�9���m0�= �r�h5�[���N�V�	iG6�� ^��#�7\��.����[��匨={2�#(�������:��հ�(��	n&�����;�17(�G����yu�^^���D��v�P�#tJƫz�D��i5��v�-a˻��F!����p���g���۷J��6��y|�Z��E�k#y��mS���):PB�r�t{g	x��5)�ݝt���i�N�8D�2M�o��Y���w.�
&�Ђ����e�����5��#���*5~��u��5�ѭ���4(U��f%}B����1e����8QS:Ug�=��c� �?HO�����t���X���DR�XE8b�'���qR5Y�2L��0'xo��-hcL�����z����:27-4�_+�u��n���"�Y�|��TW<���2b}�J)Ҳ�ݚ-��6��bn(f�WY����e��㱥-i�V^1ǰ���^���F�!�;Ru��A�V�f�&l@��I��i{0󆍕k��}ւ�P֡��8�Z���w�]y�뿹��s��:���1�&��Q3�Ivt�Sf�e�&varӶ{qd�1]p���{7Y��v��wZ�s����1)�20tѩ�bm��WY�:�]����8�)�f����Oj5
p������L5���t5��vve#;T���gV�㪆��UV.+]rA�qop��r�UUu���𙼖��.���.m�A|�D	ْ���l�t�^�v����[-]�"��c�(�|��"��8G���9�x��KP�t̚0RR.���se=�YfҫB�mXƓɇ�u��'v����Ew<k�TL����a�afk�G>U���7z6��mY4UY/1���V�+���Q՞5�u=�JH�%��t!�o�i��8�in��%Un�c6�9���I�3V�3*�
D�ή��n��MK�e��1��ڳ���nWW^H�5�^[m[��D;�Z�v�Z�f�lջZl�ά�M�[p�F��&v�\j��Q�H�k�������ﲸ@��O7��z�t�0N����j�6�QLr;����a>8V�ᶇi�[�u2u�u(��j��'(4'	Ş����:4B�''V���5�N�ྣK�SA�0��X�;">���h'�oY��a��Ӿ���{]%�t�[�yU�h�U:[��9Cz�S���1\8Mk�8(L���E�1-��i�A�w�*�a�^J��E)�W�hN�1nȆ��V#;G�9��-�Z�����Y:0k��#�1�v���^QǙ,�㾙 �B����jWv�0N����Ա�y@�89wT�������顨e��*����(�
\3s�,��ΐ�+z��D���J�]�\�Ý�h#�l{������JŁw�P�Ԏ!�>5U:Y�����9�t�C��%^iJ�A˖g[]aǀ����vY��Oc��������g-��	�0=uH:��^��0�K�׍wQ�*0��Ӷ�wvS����=v9{�%�j=��S�;d�Eδ�q����q��iY�]��B�ʂl��:I^�֐+�*݋	�:v�c���*v�[Iԛ{9�N�譌(&:kҌg����=}���:V�IKъh�(��b�t�P���Yv��oc�.��E�s؍���������ՉS���й�\ԒC��l'y�Ћo#qU�SӲo�J(��"CS%֐��7��⻝���*��1I�"���/��5m-�Dzz�;o)"���s:���|�{~u�V$m�������%[�Uٛ U#Ż�nTY�j��i-q��H^a��l����N��I֎X�PZ�4z�k:�㤥`�/U0y�K��B�	}ҝ�ܻ�pw\n�J�WK�k��M���w�+��v��t�+�Z=q+#��^�hT�/8؀��4s3Z`�.�NƈZUHmW,��r��X��0���wq.p{ĕYܵU�gY�`�|I���(�2u�V%�(��t�*���k�<-p����ysS6ov�̟T��5hS=�J�'����^#��L�Y�q'_
���ó��Z�H^"�qڦ�9Gq����Dpu���(�Р��U�6�lܼ>ǎhiU�D�;	2m+-gu�^�V߼��zSu��iY��!�[�tI+r�"�#t�8��ZE�.��Z�E\u6�{{�͜VK�锶�y���J�tD�(����;�e�v�0F��Iu6i�))��KQ�ًo&��o���1C҃��-+!d�a��J=�'�Sx5\��Q�.U����&D�^�#)�CV!�+7K�����;n��T�a�Z��]�D����hFA��7��IoK4..udWґ�xrvΉ�]p)�R���\�S̮D���XvL��c���,I*j-3OWTy�֋�3�$��Z�T�+(�ܻ�b����'*�r�l(���8:��gT�;��VA�7-pv��w�:s��m���GQ�a[b�f+��+��� f�s��xi�yJQ\�����w��5@�F��z��ՙ���1�][���,�h��zg]Jtf��i�d���NY�v��S���,���ͨ�.A'Q���˕�ҕj��;N�X�g6:ď�KTļ�53��dk.\���o9��{g"� �qwC�Q�:]kI����
i���n.&Cn��Kb@�vm'�v+�8w;��*Bs5ly���˵`ĕ���c�WUqOV;�����S�p�&��,n��7G��k��u��R�e[��P��t�V*�1��\r��{�2������H=���(�0
���Ta�-�*ےn�2r(Y�{WTތ9W��p�G�kҋ��V��� �t��0��3j�D�ʒ����[cLy�`�p�y�S�[[b����w��tOr���t�!#^�[1f��8ݱ��͒�:WKڛ/+9R���0����i�ڂ�.�Ϗv�j�wM��k.ꛟd� ��{%h�'S��"�+&���|-�joh��`b�މ�w#Rg9#M��=+��N�Y�ݱ(����|_)&�C�PN��Bhm7�On��/ǐ��8��q�2p4?3��(���[�#(*a1[�4*���^곙�)�+Lz��tEFr����7��ޙ?Ma�8S�t� [R�Q��Qwo�.5�����`���H��S���%/ȵLY$��Ug�V��o���*5�^$Q�u�=B�WI�^,+$
�S�U�Λ�{˅U�fN�뮳���YmMA���~����5{ �4�h~����a����T�� '��j��7�g�:h�?rO�H�*?���Y�!��Q�C���j�����?w��S������p~���/�������~�����?����J�K_�2?�p�R�;?��$1�%"��V�unW	+�A�N��+�:B��"�k��u�T&���y2��`�#kpV"��cl⼫�#�c��}�pt��M�V��S\�ioMٜm[ɓ�r��P1	�Li�	�Q ^�j�Y����5��	�d����T�K��f ���MV�4N�o��V)�
���)���Jz�˙cYUz
��J�o7h&GW���>����mv۷x�P9����E�СuBh=��#8T�s��dn:��
�2V�Z]��h��ӡs���aGp�&7r�s�gYH|n7���Kn-�����؝uc���uu�bk/e���:�Bvtl���ѹO�-V'Su8�U�N ���j��Y]jb�S�Mُ��9.ix��6��R�pgQ���%h�1E��T+y�Xѥ55re,���$%��Ґ�������t�$�}��Q>�Pw[q:��;�����߁�5�r�TV�nQ���1KL�� �������Q�G�[�y�s�	*��ҫ+"P���|Y�M�7L�]?
=����鲐}�m��u�q�3e��]���WX�<�p�����LH��]vF̳�o���d%U*wAY�i�=�I݈��1QQ��9`�E����y��V�C,�U�ʐ�ݳ����=�K�n^����;�),�U_�������{}���<x����ǎx��Ǐ>�<x���Ǐ>�<x���Ǐ�<x����Ǐ��Ǐ<~<x�<x��Ǐ��<x�����}��o��o<zx��ǏO<x���Ǐ�<x����Ǐ�<x������Ǐ<x����<x��Ǐ��=<x��Ǐo��=��x�������}>ߧ���l�2i�J�P��*Ua�� �c
|�]L��v;�\�XV��� ԇ�����3U�\�Ľ�kh���N�lݩ\T��(���]�k��r��E���u��4n�ҳ%���آ$�P�0���B�K÷�Ժ�Rp͐�Ιg1ueD�)���]81gq���]!zQ�=��\�2|��7_wr}Ar��L�ۛ��.�/��j�Yj��v{#�+���C�f��Z;��w$���!���N]x�Wu�:�6��4���Lp׀�(iQ���2�A��UV��3n7��.c��U�IT��]�T|���`�P�R��^\ү'Ȭ�S0�� ���vi�oٜ��KcoK�]{�[Dk�'��w�]r�9�o9	j�#d��z�s]�EU�栽Vh���F
q��=��v*��P�۵�B�XoxB��gD������i��f���OZ��V�.�g�,u#5z6�����{�\����Z�%<�}y�E*�\�ir���R9�^P�U���GBkv�zp���W���K�`��rI��U*	��nfd�w�q�J��퓭�&
��vJ�O[y%���0�9r���v&/2���v�j�*�ap;˭�H�������|�
�9+20���՗״��\t$���
1��vY�o�i<u�/��f��;!�_���~y�sߧǏo����ǧ�<x���ǏO3Ǐ�9��ǃǏ<x��Ǐ�<x����ǎx��ǏO<x���Ǐ>�<x���Ǐ<x�x�~?��~>�<x����x��Ǐ<|x<x��Ǐ<|x�<x����Ǐ�<x���Ǐ<}<x�<x��Ǐ�3Ǐ<x�����Ǐ<x����<M��!aᩓ<;�,g��٩�r�l{SK.�i���c)����;Y����q�^�ﯰ��f	u�R��(cVrJ����Y��(s*j5q`��f���ǵ�����cTT�B��	�H�${t=ɹA����72���N䗭]Y6z����u��!`�-;�Ƶ���&�fn�yҕ9L�T@��c/��d�;V�X-��h���t,����ɳ�n������3JPՕ����u)�A�C�ԘS��ȱwjJ�L��pL�E;=�qo��M��tv-�)��BI5��O��h�pxԨOe(r6f.��n�}{Y�M����r0��ҵ�9yn^����}t��D̾c$��ayTl���7T�],��
�F(�htoA�@��:� "��'r����Ϊ�]Gt�c��р"�][�Ŕ�ޑ�.��$z�ǧy���5�]v�r��-��V�D�Å
$:,���ӕ��ob��5�Vڻn��]
v3$�S�{�hea$�x(�P��O�q�Uݒ����.tk.P��6w]�hӉ^ʊ��aJM�����e��;ZC㪕�F�M�n�,�Mw�=��r�#����{�Y��D�"hڱ�9[6��8�,�I�,[�i51�r�+n��u�M���*8����U,fJځ���݋�
1hx�mc��[�xT��u1/�M�'଺ŸV�ѕq�`.�;���ƒ��$�ܤ�Sz��٭��x2
'��w�
��0Z�D]���B3rve�ZN�s��{����s���� WU���ʫl[ˤ�ާ���x�voS�η�D޽���+�٠.Ȳ,.1�KEsy!��fS���[����
9j��z5BnH���8�G[]ը�XtCς�k�-�E�z�:a����-�tf�,a0tX��0��NU�U�Ùn�*ƝUwM��Ma�/c��gǮ�i�)t�|{���`�٧a��[�����e�&����$�.��oD���ڃ�VC�d�K�ou�iDY8�ՎTӵ��сu��m�|�F���V,Ha,]��#���Ƀ/��I�g!i�>GeU9w�u=eL�4��~/�Juo�Gi���~�Ũ�n#������4���sɜm��ǯ&����:K+a�gs^V^�&�o�;s6b[�˓�N=�]:ؘ$�i�g/�f�#CԶv}H]��c�	6�
ه�	қ�ڡ8�>���%�S5�gN�[��_L�M�̷�:S�� ��/��Spn�+��L
*ǩ������	݆>�,nl��MgK��7q����|�[q��v�G�P��kC�N�K�A�h�]v�8��pM-���(i)�+9�釯��M��I����9ͦjH;Z��Y��\h\nZ�WP��G�a��ȫ�����Q��}�rb�8��l��AX�&�̮X�%8u�K�F�:�}R�V��B㛓^sD;;cF����6� ���S}b�z-�J��ެ�J�JF�|�u�wi�v��cYLe/�0�u���r��g	��꺖]a��];�t�.e�(\�.����A���V�������/pތM�� �at�ҼSJ����ݒ��V��3��q�.�&s�ns���=va��m���([4�*T����^��9ڤom򷷰=2f�l�>$���
V�mޟw�nhvh9q�Z.F���YmbD�".���K�T����X���=� ԭ�U"©Up)��d��էi��x����N�^-f��]�7�l.Č�:\�/pa�;���CE�Y�\���ՏC	T�v��IL�Ό:�Y�\�r=��.vE������cp v��Ź�\�u�CB=
���P��U��C��;��3��}���A�zv�P��ŦƋ���C���D��6-�4�J����M4��ܽNS���7�}���Tm�^GG���Y����2�z�:փC���BgD�z���Z���j�܁VnAp�o+�%����b�햴X̅��c��:�cR��U�&`���ۀ�PZ�l^��;!�m��9BX�B
��X��|h�v�C4QziT�Ǟx_>���Un��j��qu:�|㎺8��HUe�z�C��Ԟ�e�ёv�
�,:T��S�}7]k[��tʢ����:��*�gJ�B�Mٷ����w+C7��Ja����lA���٪|NA���hBp�f�9��K�oV48`N��
W3o/i�{j�T����^��&�z�c-K@r�v�@��5��JC�\y*��Aة#۵��`4�n�H�Zj٭�;۬�Yy�r���o��\�b��+>�u���	UV�T���U�I��W�iޣ�F�.v�6��)X�Jc8U�%�3�fL�B��
i�.$������'*�J3 �k^)�Z֑g�wKs�U-<U�gȻۖ�:�5�U��B����CyX��3���B0u�=�36T���x�'�Jd2��b�5��Z&q,��'��ۮ�f����.��L-u�|1
�L��,�}Y��+XVS! �3�� �H���Ī��h,/tM��Nʵ.#۴
��:U��3�s����1Z��gs�#���7�Ws)���^���Ѫ�,�����*��5�	�ۮP�e���V���w�ټ%;���"��w�j�V���.���u�7�-��v���Q��]<�^�nTs[���7{��+�+G���l��S�Em8N��5��d͌Q���d�L&ƽ�:��t��@ī�L;�b��m��!odB1]�u���^fRS���owf��ȭ�tv�Wa"��aɎ�4bި���U�kv��XS4���p��SK��5�һ}��RT��Y$w
�>���t�=[۰�Pr\E�#7(m��*X7t����d+.���S���d���ޙ���Y���E��ݾܗi�v��w�1�1���a�����,Ys[t��&� �,C���Lø(�d��͊�H���A����-���G�r]�b$��
��b�.8Y�T`6U=Ǖv�u�t�����;R븆�Lhq���*�p��L�[:Z\�v'1�׼��|�8����:��{ui�ra�
�@�OB�[�3��."$j�)Q��`p_R��{�%vR;�)Z5��[���pA�#�z���!w�Y~�y�P��*\+u��U�ܽha���8"�[�N*'9n5́���h��.�Ӝlå��"�;p0XΏM����J�Y�w:nb��!��JO��`�8�Q6.v���Y�l�˽���;��=�	�X��U	1*�v����� ��D�j���oe��*!;���;
=Ӧ�4� ��q/�__Y�V��b��Y�v��%F�����ԭ���d<!���]'f��;qt�fё]ձݶ���h,�ׅa+ ���y�ȉ���*���e�����]�lW|����6^W�,c-�V�+�1"胤�W�H��Ԟ�5L�|���n�M�vK�Ȝ��D��U�'dN U��"u�C�\�m�uu�9lU�x1�����.�5�n���'-!"�ʌ�7�z ��y�����^�1��5����$|m�&���.l�v�6��%��О��}u�{��X�yi�t3E�Re5i�,�}�ܫh�東�ʷ�-����ew٥��+˦��25LyX��5)��Y=6M(+ʒ����T�-Q���m����q�;Ӷ���_B�%��M�n�^Zd2�"cD�w��+%cx�#��D���usq��KVmS�a�^9�鄆G%���uڲ#֪T��q-pۛ�ƚŎ����Xz�Vt��WN���
,l�,㠯F�}�-8@�m=�J7�ݭ���$�)e��W�0+v��pf�Z'�LQ���Ί.�t������dA\f�I���#-^��P�ʵtz���I˚w�p�}ۻ�yh����(�Q����R��fNHN���lԸ��2�]��8��2�s>M��/m�;�w@m��U\�<�JK����֐�����u%G$���	��>Ω��Kn�5��S.�,@�g1O��vU�[�C}(��J�y[��1kh�E\v�.d����ތ��J�,�u�Π�I�E��ɗ@i���N�i;Am���ںnlǖ��Z46�u
hg\�C�\��qw`"ftՒ8C7���5ޡ2W(v6g�Y�n�N��TY�mX�,@L ]D�Ab�X�FĪ�u��p%(�b�f��O"�@`���;na.i�Ԯ;����֧7����h��O�(�̷�}��~�E�d��-�v¹eT,aG��D�ჺ�>�L?:r�
zw=����ax�T�̇�K���/bEp�̤UQ.�����j2ob�Y!��u����U=c�p�y�m�����`�xdUee6������2����R[Xf73	�#9�3iB%�y�V���^�K)��.�\'�(=JK�?U��D�f�_Ǎ
��Fe$��h��aU�;�^�`h��tn������qa���Uk~"�h̨�=o�Iyr]'�oʾ͆�(_n�q��Q���ql�09��r%;�|�NN�ܻ�&8��]wJ��R)�e���*��wUE��z�vWj�oݡ�۾C��q
٫����<��t��˧�{u�duz�K7f��yw�s��U��B�$��KL�5�LU�5E�ĉm�������[�S�+�{��xT:V�9]
��d\e�b���|������<���e�[[�u
G$=}t�I�򶎍��Į��R�w]�Ejئ�_-����B��{xq�|sO�&�݄�*�燬K5D��]+d,ާ1�9&�!��nΤ��!���[&��G�s(j�?M1�����$s��}�J���ٔ����j���Iw,�r�I���^�U���v�8�˵z���������r7���pIxl��&&*Ƨ��]�1	3P����[����Õ�I����W6�����c���=�e,RB�i&tpune�e�cpcOׂ��_O#�\�B�'��:ӂ����GY���e-�����R����0�h6a0��*aSgK�(ZʣfS�Y[}\�=�$5���/�����]���cA�.eJ�ky���75���hL'Ufob�=�[��e�T�f�Ť �[|�> �^jl{�~�PY�p�ӫ���i�<
�L��5Vc��J?�0��\&S)��ӑȮ�#�dWP��u�F
07��r���� �J�o��:�*jt!V���\��rG;.q9e��8v�l���&�䢝�K�/X5� �V�^Go��f53
U�t)Y,�kt����ou^f3�u�#�(�^b35+�QÃ���B��P��yӯ���a�9=z��+��a�6tg��B1@x��֓�e���,�;[���x��|R�yhJ��� Wv[�5S�7��M�E��/nX�u!=���u�|�?>w�^����?UTW���7�{�O�������'���	/�����uDn������.�۬�VE��7T[.�AF�"�b@��~)0� ��(E�,� Lh�ԅ&tѵf욅@������D5�CQ�2	i��??�pX[�R��&������S�m;#��ۭ-���C:��V^I+s�[��6i�$K�A��U4���YYt�2�b�V�g��X�t��93F��ȥ�QܭK]B�摌[+kz�"����fR��� j`]�<�H=�%��y�dZ8�B�+P`��<	���䨲�:�����+�*&�냂._)�q�iN��s5�ຶ�����T3zT������]V�����`���=�k����n�9[W��e�2�Y�R���}O3$5�\
 U�Wj�5|M�&�S5إG�ϳ��Y��%��p�҅oU�>}�x�V��a�&��X</x�S�m�Tn�	CL���f���Teo1�s���X�J�~��U'x�C��Crnbo_B��h��n��{s:�q@ &��޷�|��ݑ��"�]m��8���B��ݫm��,@�\�)וs�܌n��	oY��M:�E�7��%�M���#�HO>Fì0��7�-�΁\%%;&�l�Վ���r\�oH���NҼ�7ja�C9�Yڎ��{�E��V̩�����}cL��a{*��)��z�4��E����nfVU'�z)�fI�U�c���b����W.�JMN�/&Z?�W�NN�W�ӹөQv���U�`�ѳW+D�
�R������X$�ЂYF �&��TI&�m�b4��Hk��Qbiˠѧ�0B�K@��&9F�U�H�?��2�f$*�(
bD1�A*T��#(DSM��-�Ca@�A��4�8���B��u�D�8�	���@��t�!9
-�[ƥP�S$%��BIQ���D�h�_�0)mF	D��]]��%Q��DEQL��Z�Z�5AE4��DAEs����o������~?<g�k��TU�T�A4UE4E�tt]F	�Ji*��Q3<x��x���~?������>p�"���K�����!� �m��RPT4R���*(-a��)��kN�b���vLW�u��URSE1D�wh��J���fb����b*)*���.�PU�ADSw�TIE�N��
*��u8�)��(���(��)�����:d��*)*!�"�
b�d(���"
* �(�JJd�ih�$�TM<a�LUQMP���T��O�;������uKEY�Oe���&��F�?.��N��E4j����U��dŭ{�u��bb֊")��Ν���)ɣb,V�c�F�kV�k@V,�j�Qb�Ul�$�b�ll8�b+:��kF���kM�cY6m�ΝK����Ha�b�#Y*"6��須����:�5�4v)v-�ǿ� �Fd(@�D�s*|73k�U���5Wy.`�q��zC\L�Q�ƾ�ޔ�[�_��Cg���`���٫��}.k88Ic��e��q2�d��)�!��"Ii��\��j���j��ѽVw��O��gc�u4�W�xf,�5PT	�ʗ�~��p���02�z�cdk�k�~�L��&����Y٧�k��$��Kzx�Y��u�y۷�H�ᢉ�μ��ƀ$�%�l�;!�����kX���}�o�b����~������x�ҩ��9T~�1�gxy�j�%w���O�ᜐX���}��b��k�tm��'Ma��kɩ��s̽�ҧ��PC7���Ǧ_�u��d7s�1�����#�ύ���G�_��8^��T��:<������I�^��{)��"�F�b-�t����7.{[�s��]C���]�^���:�a�u��P_yM�閞�L����=&\�����ظ&4^X��66.H6f���	8��!m������W�/;C����)�RS��-�_�r�'C��SUt�K7N�Q��5;�T�3��j�uuu��J�1�D�"�����d� �^�#y����ʽ�Dʨ�oe����$1��!��T��/x3l�'��U,)���ށ*�-��%��ntgvM�����W0R�(1(����/�ȫk�e��ib�v�ؾ�=���9�]�K��|*w���B��ͽ�x��=�i�]�yJI]&�x�T��!���tG����Ы�g�|T�h�$�5_Qo�7fw���G��_���Ϸ���J4UN[ι�]�X�m��=�N���w\6|�t~��7��'����Yt�U��:�Þ{�3۔��~ύ/}:σpyo�����g����̻���N��LY۹r�}V���P���p�;C\���K��}�̋���:8�c��s<
�{�٭^x`�f}3 ��+z4ޱ0�ȍ'%�h���>���-�x�i<e����������K�;�[��cS��dN�n �W;�K��� g��
y0�x$�:�V����i�E�w�h�گa��]J8f��`�>�2h��M����c!�M�T^�[HlR��b������*ٰJ�}�s���v�0 H��1%���K��w���`E�f��[Ԅ�p͏p�ӗc�Ʊ�=�a���� ͗��r�w[-ʓ�RZ�����4/�O��V��;/��_�_y�:`�$�?��ö/�C7����bO}_���=��%�Xw�>E;k���>���w�y%�\ˁkK���i�]m�-�߃�BK!9�k�;|[�П����=��cƊ��=�vF�o�s�w�-��Z��dePs^�a���ȫ.�˟c�S5�rCb��[�=�D�q��S�������u��.[��CO�:<���z��7K:O�����|$��laI��h�)f1o=t���l⇆N|���Og*V9���̙NT�\Cfzj=���m�\Ű#�����W���r{~�윀[��q������^d�G%@�{�v�_����"�����*���QMk�Jǂ������Ӑ���s�z<)��x?N�Z��_�(�
���"�Q���O��H8��f��R@~�7�K���N�r�]m9��^�m���t��f�mVymUh�|zd��G~��Nݻ�9xk��g�(��a�˷���M>�<͜I-��U>�3^�}֯��~�v��k��U�
�^�5B6�ovq�Ԟ�Z�*3��0|��A�֦8�4	���1��O� �̜�~�A�A��nX[����ߛ{�7}B3��������=^��[�NdU��.�c4�1>���΍O:�(�v���6�g�F	~x&�4hA�Tn <�.#j�Ev���3Β�w9�X�^c~�^ ��t���p�{E<�	�#�h��k��{�����ͥ��<"�x���X0y��*��w�ȡ�'�C��{+��L�w>c�1/l���鿶��*!CxyoǾ�������M=��o��΅!�lM�3c�+���z���x�m����<����2�O��W<ܬ�^�<��%�������MxY��3�3z6�8�`�� 0�Fm!�Xy�Uqޞw�����o�Ժsڏ�@��t{�hX�S������[ǅ��f���K��!}���<��'^��M��w�����2���j흖�6���NF"�vr���k��COo0�kθ����o9�r��R�S)�~�Kb}gg�<vU�1uQav��:ĪuuN��چNt� Ti���T;����n,9��nt�uj	��J�YY�'�
��;��B!/������T��K��41��:�x�a�
��?xCEk"{�r�ϢaT����y�d��i�5(��b�&׬+��.�C��o݀�M���v�W��g�Nf���,�S�t/;���$�ӆ��1�_��=����o.*�{z˲)
{��G��t{|~��o�;��yG�B�ީ���!&������*�`wn"jv��\��x�vdQ��'��6��Q��T�={�t��x�v�LY�.��w�9d�>��4�"���j{.��aF�*�dK��b�L�a�V��F�s�$@��w5�&�<^���6�{¯;�߆7����./>���)�.Dp5����z|7��2�dp��{�Eߓȷ��lJ"��z�<��
x�O�#b��3�_�S�uҵH���2ihA�9���O:��y��O�@���G����6OU�M��&��b�ER����;1����H����ćYl�I�DgtZ���=ǽ�/	��%��|��C�⡶~`���J�L�.9[��uޚ�TSU�t��+++�ǒ���uTrE�6�l^5x�m*=�eSi尰��Z��H��k�{������w��7�I�~�#p�j�[�WSe�J��xbo���'Ӆ�3���=��~Ľ������?m��y|}�I��5U`�l�b�s��^ٿ;~S�e�k�3_�Wʬ��KȳWOM
"��zH��N0Ì�#�[F�~����)�M�{�N�:>��lU=��P1�J!K6�m�+ޮ/�ī�gO{��0�$��v����l��T��'�������ǹ�
�7W�����⧟��77��t�r�m���-�! D6�w�hWG���dOt��u)�>�����O���Z��ɾ]����u[�]��_��y8lil���K�k:h��&nX�P���"3(ׄLt�ہ�H��t�Q��I=��6���Mt����r#��>��c�9PJ߈g��}��+߰7��5�/�+��ˇ��*7���Z����I�nl��mvsN����Q��Ð�BsGh�)���O|;���<���a����m�h2F�;�keS�j��Y��Z+e�X�:��0n��+�{����.g2���];:�i�6�����R��F�c�|�6�=�#z����s"��7^�����~���lng�m�m�r�z�X��� ��gh����3�cƩ�n��Lbi�@��s�$GC�E�tE�a|$���k��8�3����h��ƨ>��k�:�W>�2>DAm����;l?�u�x�qX:�x�l�69�x�oz���}��M��u$m,6<7�������qPϟ������TɠE�̠=7�ީ&��������:�b;(�:��ˡ�W��i��9�oOC��y1����viǧ��[�[��ɝ�T���u<���y���x���[}�b��uh�o5WmȂ,���h�&�������� d@��C��,.'�ܯ2�̓p�Q.(����e��zk\�A��u��0i^����M�vM��+�E*\�7Wx�}�\��=S3�)�w�3�9{�X�������VvWv����;4���;Γ�N���ȸW*f����{��i�����y5���ooE�X>�:�Zkf���]�Nܛ�����$�]X7uƺ�̅-�1t��v�G�U�j��l��v;�d�t;q(e����UA���;���,v��{����+����2Tq���f��<�*`Q���g��[^��g<6�H�}f罢��o-�y�pNh�z}\�|���R�u����^p�>y5qgز�_��Cyo{����)�ol$,L��d�3�C��@�3�wSe囖3U���W�"@��:���[u7Ubf���:I��G�^���x��l�gݚV����8\F_�K/GsT���.�z�$\v��W��4<pɯA����i����m�*�w��̌o}�(�e�X8@�;>�$�9:I�Px�m`���}�i�������2
�ۈ�j�����$��$6���!�h��`n#�����ev�\S�^
�g�������o�잲A�ꆥOI�/�W�ڵ�2��c��g�k�8�_v���c.��M�߷������mA�Ӻ�q��׺^Y��(ll�u����Y��}�>�^���	ꯄt{���v������0U߳�L���^�W�.�Fͤ��6�cbr*�}+M��+Z����Y��y%r㫪]�Z�w-Xy��M�#�K���sI{\�TOX�PE׬�����w�rj=���o2-��]�M
��z��}/g���+�<h��+9��y˝�wȶ�Tf��[�ݚ�ͦT���Ӳ��d�����گ��M�~�5ֻܡ�j{'5��$�E�����"���c�T~[=&��;�О
gm,�����]�J���>��4OPI�k=Y�"�z���4�_s��w�i��'�����Cw}�*Z�>��V���{ל�_>��Ǐ'��}(���+���À����2º#�]�������h�/��w���jC�w� ��<H��{[��{���X���V�a�Y���d�G^��쓜��7���'o���diឬ�#b�϶Y�u�U8P���߯�[��D^�[���r���$�z������Cފ������Q2ת����#w�ز����4������ο��dQ2hAۧ��5bbk6a����\�6y��g�wUR��-�ڢ����l�th�XE�s�?x�+�O�SM�l6
?Y	��"�!�f7�ƖJ�ˤ1�"s&�6�引ok�����;i�� ˷bq�����gv-
���9�Naw�"h�Ӛ��6��`�� m���	�}�x,���[o׾��z��}��My]��뗽G�@��8��� �5��[�hVnt�y5^7�yN�tS�[�OO	qV�Ip ���p?�������UAW����܁FI�2x޼��ζ���������->�mu]gd�s���=����rw������&y��k��iP�j�6�����L^��>�!��吝ɝ'n��O����~�����er�;9eI޿kk��?���.���^X(C�	�>��`�7�d��y��8�����y�������g�f|��;>7�Y�C��t�h2z*ׇv�E��9yz�R^{�׼�Z&}4T��S�������×m���Y�gy�ن�Po\��]�6c�Rú!xKak�}��<<�I�e���țy^g�a}��z,�/�
�=v�SNQ{�-̆����Q�'i�6�:1&e���o^��t�ξ�N��q(��(X�*���]n��/C�lt%"$�ރP�kp[�3�]�h������f'�\��ڴE�n@�Y9Sds��E˲��v۬Ea�unnۉ����%Ќ�ͺQԤ�{�ހ�t���w�/K��}7�+1}�Z�sK=oH�ڊ]��������F��s�o%9���Za����)J9R�̭�!�ɩO���U�/p�$�|*F�.8��ɴ�[�C�9�6���I����3*�7Z �	R-��lM]9Je]�WI�Gc �|�	\[=U��鵦s�F�O��儡U��F���szG�udm,�i���,���V��:��mn�[�����dب�Et���U��=D��X9���i>}11Y8��q��{ݶӭ�CE�q��ۜ��L�ԟQ�F�&���B��ݜ��w���D��/\�2Ǖٿn�ۃ�Q��,Tֻ��g��_@����Ɠ�v^W$Մ쉖����"�bŮ�k��_b5.��t̼�!�C*��5N�(7�6��CG*\����&]�N���3	�����&!�H,��*٩�b�4M҃{�К+t�̃P5�s2Xʆ��ӣ�3��wm�Pz��ml��1���y�P��%ˮH�=J����T�>�@��z�Ue>Z�����x+I���);�:1���8�S^-Hqwv.��ԕxz��3��.w��)�����iLns7:�ҽ=�����7s�U�ts�gH԰�x���"��U����_{�{xR��Ɣ�"�Bz�Y����v,��E-U�c�F^ʌ�[p�[z7:
��]',xV!+r���d��Őڮ9)�$w!�[�Y��e�!<��R�ݓ�V�
�5�7�S���碘�W�]���$����.�譪\���d<)���ɣg^��ݍ�Q��[)�f!���K��E7���8�Lr��+�{�����0jݥz�����tQ��'��rm��ف�Iv�4��ֹ����`Ѕ:�i��&G݂�ot3������b#
2�� 9ׁ��Q��]wa�0d����J�}���)�xje�h:�O	����%񏚺v��>Y��Km��ղ�u�:'a`�o'��,��(���C����H�3����4v����'jmQı;M�ٳƹ��ٺ4�W�Q�M���J끾k*d���C�672_Gy�ZҚZ�vs�c��O�V+qT���t���M�̾�"�z�*��n�J*�Vͭ�������X�{T-�X�n�c��i^����˯�t�y�Ml�6���N2n�+����ռ��i��\YW"����|����^e[�����ý�ǉ!*:]��N���դ���X
�(U_0iͬ�Ab��΢5$���c��w'qGDF5����Q/PDU���u���F������~�x�~?�������~�>�F��5���5�9: ���L�F�g=�QX)�&�������cE9�3f��"	ϧ�����||~?���������[b�����n�Jz�MQTy�趎��t@bQU$ơ"h+F�����M��'!;�AS�ų��� ��b&��E��X�R���;������bj����)��������"b��((����b���15E4�4��a"h(h�
���h�Ѫ����j*I�!����J��1QDAB�]���)�詊JZ+Z�

"&����b�!�!)(hpA�m�WC4D�P�PLӯWD5TD�WYEUQđUw�TI�D�u��1UUPQDEu��D�T1DSEBSETQU����^�>0N���3F܏:b5�
.�b���jQ�YE�tov��G:�ӊ��[��=yΒ��.�c:��������FѪ3��la59�m���oW����0���A!�hH�i�	���`�뤢J�*Ƨ�0�.���s��H{C�T: Ƒm�㞱�﷨sH��@3MvIa�\�7���ȼ�o&���H���;�������lKE<+B��|9��<���*~��U�w�Q m��׭NHp[VWH~��4���U�k>��`__L?�p�O��AI00!`�\zyL��j+�3��@77��^�M�5�;=:%d=��5�ν&=͍O�q�N�:� ?��YE_�/�C�G�!�\�,�d��y��{x�2���d\��Ijw�{`��hOB��HP2v$�02t��0�1	�=ou����J��1��g��%ܗM��D�K�K#U���vO0"��{��;���]�r��Z�ZM!��G)f��1�},�Od�q#z�$�b)9Y���y�7^ǳC{�2ݎv(�if���H4&f�?�hLpm��i/�:�.�������<�_���y���2��ǽ�#���
�a+�/�+#�=(�r��}��zD߰�ֻP����7'�)��]�UlK���5���3�h���*����*�9;ybK���E��=����w����p��nV��C��V7����3g�-�Z��g�I�����/@螛=w�h�q�%�$U��Y5���.1ٍ����՗ނ����91�v�G��CT:&8_��v��v�>`���'�#]t�n���vG��9���n�{�b�����_���y�n} �A��,b��/��ි'W���|����v������ɜ⇫�;����az��1�`=��V٭�� �����}X-��O[������\$$=������Qt�7>ϻ��E87��i�)��;�W��W�r1�P/a�PUQ���De�=��ʐ�lg����`�G�&��n`c%�!����k�kÌ�v����;ϒ��b��ʻ�^��7=x��${�='�/3ͼ7����!�ߚ�`�V&-���@�W]ޱV7�۵[kP�/�W�5R�ܲM�⽭�0�?�Ȍ����-�s�>�xL�� {�d_�{>�����o��?�Z�C���{��.��Id���� ��8�S/�T��c�a�0/�H�(B�����sm��dh�(x�zdATV�	�����!*�	cIuc9~o[[\�C�����o����Ts����-uDO!���-	��i�nj0y�d�ֱ�)w�`]T)\�,)�=0;���)�F=��w���[�9��`|�뾪�!�s>���]��T�$����l�j��~.X�����/u�zQ���I��R�ƒ��[�C�i^����n��r�M���D ���у��2�����	-���3L�zTC�K�SqLt����&(�ڌw�����W3W妥S�)�7�L���+�A�����%��F�H'ݒ����$�b%��ZJ���E;x��:�:�`�"�!�C��z` �[yH1�0��a�n����{�Re��& ��N�Z��>�m��ڸ_l������B�zw�xo'�l�>6��Nj`p�o�K �v�u�j8tQ�Q���P�����L��<���>����k�]�%�r���C�PC���R򟊸��Ϋ�7����x������*��W<�j�������H?ݍb������\�ؾ|���79OVm��=�)��4�'�
�~s']�U-t�����$���W+A05'yk�Ԛ�Ӿ�N�z������`1����05�}zhZ�2d?��C��eA/l�����$e�LO3U�z[����x�yU�؏38������fY ^笰v�����o��;NT��Rw�w��ۗ��U��b��=}5�Oa�u!H�x�
<�Mm11��n�fI��;gge&3{wLl*�y���=��n�����L˴�t;>��Y^Pj$�|<ĚyF����Q�����/}N�%��w�0�Q7'qa<��N �ۋ�>���m^�rZS�G���Z
���7��{����b�٥&���WV8�G�(f�ޘ�;�窢qb��9,5EC.󮺣jd=y8[��Αw_fdeF��݆a���{�2�>�o2����}@9���2�#Ļ�^J/^k��C�Q��O.�iY���ϰk��Q#�W�g��>���ٜ=���a}�1El\e<K�zd3`k��[Gd�B��X�hy��n��b��{����峗z�/B����z���S��o�����T�&��L�[��R=�ve^��(�J��z�ǹ�����y�h�y��k�S�{��i�C�[X�,�}u�v1�٘nmJ>��>�G�*��O���e	x��ͨ��#����l�T1U�h�e������J|��<c����<��Bb'���� ���5���{�콠ܥ0,�����f~u3���Z-b@8����c����G2{�����U�R��O�ۄ=������X�%�u�7E1�� �7<�
�?��9���Gܽ����2�ռ��=ۭs���n^5>f�$Á��c�L9L"�s�1�b�v������p������u�tܾ�ˋ	��7a����f����c �zl���7��������?7���A?���M���&�usx�4Gu!�w)�{!��sH����BbK��X�nEo@z��fº�wfB���{� ޻��\��ϹtQ�gH���u�n��t��5Ȳ��)m���ͧ�诒�����+�6��֠��rnH��O^�}K�����;o�A]�%�C���H�hت�gC��G5	:�<�(�c�Ӧ��5�q��0��l�Yb.)����}�����!��S�N;�8�Dk�0�����Bb[	�-l�	�aC�H^}��G��ؿT�e����A��m���Nj�[�@A_�a?��(:�1�	�P��~����������<1��趏���eH���~k���f4X(������'�������[��=�q���'��ݛ�����܀�h����Ǥ�- ����`:"صxuϚa�{�]��8��*~�t4����ie �u����{��_��@a�/�F�Š>�i�A}�oN�T?N^���$�lN�p����,&ښ���l`$C�pOB^���mi�Φi��%��r��3�S�Zy��-(�Hx��u�o-�hnhg�顳�M1���csS��~�:*��;(0l17[�7I�\S�*��lӈ{�d9��/mo>���yh0)�0>���`t�}���Q�9l��f���SΪ��'�(y�q�]�%<�F@��%t�
�ǡoV�^��7�� �d�,.@���l�ǐ�	Ū'\�<Nu�:*�=0]3�b�B	�Q,��)H��(�k�Dn>08=������	�˞-n�0��N�7 Q��w߳לh�Ea9�\@��sT�9�J��VnōO'v��Y\x��#-��u-�.cؖnֈv��r�i\ZN�r��9[�@������t���xb4��*�o�z�̣�٧ �e�7����>�����;��!�!�l�f�p��H�>����'.��H�)MM�7m�[�d:�`�Pپz�e�0P���q��-�n�1����Y��ކ7��O�"��
��kUse�fqTU
)�x���|�/X.��x/��|w@��e���TCQt�y辙v�n*�c?`�Y����u!�\F>��xj=4�OE����c!��g�9�x`<qD��3�����-lF��Dp�#��7 cd:�1���}G=7��������7s�2~<&D멩�OpC�Ww��/%�5��V�~	JO�`b2[��j��T����ٻ}�t�A�=�s���uv������g���R폲,�V�a��5�8ɺ}[`�sI~����1�`�]���71�5?�,��pbs�b�=�A�:RS��Šv��u;x��1bWVVfBye��1���!�l�K�����
#�4�&9������֟ga�5�h�Wv,�4g8�Sж�t��/zjC���G>�� w���~��D��GE�8�����g){5��y}B#~����S�hܿ5��y���8�e˱�{Re� ms��p����Y+b��s�$*���10�Ӻ[�gb���&^�Ck�*V^�W��-�<g|�> �k�	�7����y][f������fE�F@���g[�ow��͜|�y���������lh~�ɐH$��~��Z;��=���k���OٰR@<bO���g�+�p~��v��]轂*f���:��~e�cx8��Csp�#8�C6q��l��s�y�=`ǆNI�-�3�UO�9�׏&ڒ֍}`�c��;v�Ecj�!?5���p+֠K�m��cm�eE����f�D��� F���d�=�^�q��L$
�!�tS&ܘ\�=�2��_(��ek��(RXK,���f/[��Bڥ����P�k�6,�k☁��_��z�������d���t�8b%:���h_j���g�i��W����i��x�����l���-��@ׁ�V�x�����*S.	��[�X�r�*ל({K�`/����2�Ɓ�3e��-ᄍc!��r�zc��y�%���!5��z	�髜!��S��ްT["�x��ظ�������P ���|(?+k������R�����#��^z�OC��]�4ȜC&�%s�P�r���%�y�o��+ݐ�����Htks�}��=��`jnQX����ubj|XYc��/|J�aV�@�3a]k	/v���i~&���>S�rK�פ��Z;NNG�u��yԕ�h��w����%�7y���uh���݅(z��G�=���k+ʂn�����𓲹�	��&��RZۜox ���W&��N��R��Rby���m�/��׋�Zt���d���{���½����W�^[j,�!�`����X8�8��Ík�/ML`ێ�1�Z�T{Ľ��Q� ��<�;-�ʉC�,E�������4���9�0̰�T0���8!tռl��p�\�S��Y�7i1.�T�MKsQ���^�9�"]�����0<F���_�~�I�{z]��[�6i���C�z��4��C�L[��<�P����">Ш�9�+�~���|<���â�©�77���H�v��Z=N�/"��{zB!� � ܯ��ɽC�m᎟@v�F0�xX�8�nΐ���dc�2{���Q�צ�{�C���rc���
�#^k}�M�1p�z��M.u������ܠ��^�Y�YF]J��A��Nzq��j����T��~;2�r$�=�hv,���"��h7]����_{a�LT>��tW��>8p5�6�|��^���P��D&�P�(�*m(닸��U�s�{��1}�{r�ߺn�2�7J�/����?,�0/�x��ا���b��el��	DKig�}$���U�9�C_q�=o��C�d��`��w9?�'ҝ����R)�ݺ�Vk���!p0s���mm��=E��8�֥W���w�{����u�옼�wz��1_
er�țN��n���O� ��&�f�C�:۝��l�����nh���� &u�r�8���ν��>��������9���<�s��5����ˆ�����>L�u��YX�ƒcI� ���L��zh��zkD�MM?dQ�ޒƶν.�e�;)C��E��*�]`��W���e;a~�-��6�Nj����^u�	Ї�������4����Hv���X`�=*I�ͮ��Qi��(,kˤ�L���/��l����������!�x������v�bS�����,��.��vL9���s=�[�lH6/���1��5̇�qp _9�����r@p�í�G�2���Ķ*������k8��&׬K;U��AP��Nu����W���p��D.΀��s	���:�(����8�@�Δ��d�0�P�5�v����վ��S����ܳ,3�������4B/W��x����е[M��p?O�$;d��%���	CeW��D[�:�;%߷����ׁ���ֶw����A09ח�+����}��T.�>��DA�馽Li��k��Ŝӏ�++�4^[���Zƫ�q�C�CP#!4�{d����z9��5���i�hi��A,���V�Sz�M1��w��/�s����+�j�V�|�W__�	�f���d��[B1P8n=F����_��f��Z�eekK���_�ja�:a�zV��!sw��ZV��6M( R�f+��IU�i�ٜ1��sy{��ګlAT�`ֺ�Y/Q���U��\�7���<��}������wʒ�[/�)i��ò�_���R��s���bj}<�/�ӌ�)f���%�7��f�m��pDu��/!�i�a�@��k��������) ,��%o��UX�*5.ݳ��m�m|C=9/Ƽ��m��Mhħ�+�Q��z�oǩ��=���tPy�e����3�
��q���C�o�h��\��'�%�{�*�Y4i5���l���C���eGx;ٚ���q�tg�C7\�0���;`�.�F"S��[�FSSw��y��?�k��ˬ^���=���dy���=,�@Lpe7���
Gd�t�	�V_���ct�]��N�TԸ��̶nћ�^WtD��sxIGk�?��E����D&���0��:KR{o�i�n����R�+n�h�gu4_!��R�����5&�\��z�x��}��~kÐ�3��zQ�:/7h&˾ӓ���i������D�r��C��$uaDW�X�B�"~]���91M]�QQi�m�sY=CP�x�]B�*U��ޒ���6�a\�50���ю��=�~`�=�x �U�� ��b�t�mF	�r�n�d���՝{Æ�c2�Ҝ�m�;E���6ޚE!�Z�Sb�\�2v�;�u��v��Ћ�N�]ձ]̑EA��M�n�z�� =�]����
˕�[�����O���PR�N�q�ZZ���m�WA"�	��:�9��bzI�^��@�zl�9�H%�gB5��]䤠�/�/JTQS6�;�&s�/eժ�U�Nt��k�U�_-I���ow6�(��=/�	H�e�4]b#��v�F��� ̾9��*�TooI|�����ظ�H֡���-��q�ܱ7��-��TX�#}B�^1z��C�17xE �ԫ�ΝgwIɼR8��#n�K�6���杩���TU��$�������f͕+��e6��p�JND�G��}6A&n	����V@^�W<��7lp�zxe�m6�◁���ݕ�E��+I����ݬ|M�b�����(*�&e7��g���,V�~�\��΍$Ia^g�Ruw��ѥ7�yu,+�����D/VyL�K�ʓ����\Co"��,JU�����Ī�g	�<ZY���|)ne�w���,ƬTl����8e���(�}VN��.��X�̼&��ӥ�wՠ�n���.�m����
<=�lĘ��C�����I����զ��$:-���ܘF�aJ�WeS[�)5�/�թy�U��z�j��,l��ƜQ�
ӢE�iU.����Z[�E���;Y�g��b4�x}���r����X��l���jd�p��\#��p
з��3��<����[E��e��x�w����n�f����n�n�S6��1R�O>�df��ݨ�f�K�y�G	a7:��K�<�Gu���i!�\��靅��y�H�N��c:�i��u���K|w��mG��uv���4�n���Gw|y�:�+�j���.�&eh�<a�yl�2�J{z ZC�(�91ON��niu)�\�usc����^a�s����@�T��c��)�t�.�6�eAy��Ն�X��44
K"�������j��0��޾$��G�YB�Ty,$�n��p�_k����v��F�/&�YZ����2�l��2ި�m�&t���Jz�*m�o�n��\���OP�G�>�VsѮ�ە���+d�@�H�8K�kt�r�䪝X���ڥg0�6�;ܥ�K~�3��PG����W�X�n�F�'�k;/o����Ȫ�)JF0)�Ӭ�������@�m�]@�A����Χ*�	��S���5���Z(7b��b��S={T�����')��pa�,�ѠZR4Cwt?jp�Z��T:u�/̖g��y�]��H��Sv*�ر��f�q��j�+.�-_p\^�CE�@_\���r����3%��J�$���18(����I �A ��%^�TDKDMU�R����(������N|}>�o�Ǐ�������������")j��j���A�
	������h�
�;g<x�}�x�~�>>>>>>?_�אPД�4P�E|�T����I�-T�4�H�:)B"& ����(�(�"
i���)"
R��
)�����*�5SC@�AAA]"��ZR""*(Jih�jj"(��F�P�TT�UM�DDT^����T�PP��'�����%�b�������
�(��UUIHU-3{ t%LPЕQU	�@D�R1%ABDv������*ab�&��"J(�pi
JF�
�"�m+lhJ * �if����
 ���睆�%�Q$ȣ�C�8����4V���"8V�cmWM���[�/�]��!ϴX���R-���NS\��b[��5��c
����[�����r�4ʈ�x�N�,"�(�U~O���:��>��]�]_�T;L��z����۰6�p��^iC�Ռ-��Czwf���.��oMxZ�2Xu1�e�h���*qE�9���hC�nTr��bd��6h�|%���2��9d��~l�.��}�h>�JN	��
�@�LW5�M�y����N�ގ\�S�+{	(ۡ�(��<�S_b�#}�lV��4'�Iv{ť��t�l�l��ܝ���B�G�h��S�~��SS��4-��&tކ��s��⼎�Ne$fbg$\ݣv8�����Bx��vK'�a�ma���Z~��$���W�$J ��I�fDZ��� du�||�g��>4rq�?�x� ��%8��EE��l�*�%���� �+�X�<5��������U��fˠ!�^�<d[�ʚ�<�'��t�j�K����|j*. rq��*������mUd3!@����2���ٿBh�����2��QI�%"Q��,��mcf�&����7���6 �����v���z��� �A����Џ������M�C�$�����Ņ�l�g�Ɏ6��v!�p��ضvE�.�1� ���?����5�~�М��7�Gd�Y�i��cs;r�Sϝd\��]��̨&��Y��Km�yY��QՊ��>��9#���+��m�𪾥,�
�1�/�����371�qu�E|w[%}�ֶ��B���<�C/Sq�3+�k�Q�17�U�}�rЎv��Ϝ����(���P3� ���Ǟ~>��nr�[�ޗ��U����2�W9�o'r�i��`����-�;��{���mk�nCV�4�Sꤞ���.u��sb�s����zw�~yp�������+���Y�&���S�l��u/)��:��֩���yj���^l�,k��C��+�1�u��az��6��t�X0Ԙ>1ݗ�`�R}�Ϋ�U6�8��E�]<�m]k	 ���2E��50���Lʱ�FGT�ץ�{�7�71g�.����^�T//�d㎶=+^�PK��V�V��S���O�k�5K/lJd��{�0��<�����Naٖ��՜�g��:q�ʏ`Y����F.��Ӥa�r���nj��g�AW=K��U��C���^h���M��e�Uf�f�a�N�z���*$�a��Ɉvâ-�O0�m����#�g>�oڙ�#;+5��s���-�y ;�ȴ�CzA!�(4��K��g��}CX%���va�L����Č�����
Dp��)\�`f�~�ڤ��;��-C��(�+7�tg�O���|�w���������I;u�㶩��ls|r��z��TZlP�g�̗��C��\��zL�����o�E�(�UZ9���l��͸�|1W@�Prt�XkKc\u�*��v�E$�	����LӦ�UXT��v]R
�ETy��y�_=ny��Pg��A�r( ]}��-��Q�|�?\S<{�s���L]��|i�U-�Ar�������B�P�.���D�zsX��9yۚ�\:��a \�C����O����4L�C�/+c+U-�^�"Sh�tቓ�嫸��B+�~׿{�MUu۶3<�-QD"��-���|��l��(\*��9�Ѻ:�x�'��3�s��LP�"�]�٘�V�*��0 B��?|���s(����|~-��Q�~yz+�%o�_�1�eW�ze'E����Ų���a^p:+�S��'�}k���s3�mR}"Mh���#�.z���+�L=s�t�m�f�I�K�6b�v�:��w7]���.�lӹG����5:{���!���?7C����ׅ��P��Ut=��������hܻm򓷼�7n$橇-�!�%����Zc�kuzbK�����r+GF z��^Fl����wSE�p��)z�祐9��8x���k�����3�f�^�-L����	N0�٩��|vCl��/��=K�}cU؇E�]?t�����(�������>@��#�V;]����U`��_*ڛL�{�qS<��K�������9�l�k��;�c/������ݜ"-�9Nc� rI��1�����썼9�u�}d�u�}��%"���x�ͦ��m)aoqwT��^Ai�˃t~U?�	��T@����w9�ׯ:�x����m�&�e޸�����׉�i;rK�1a���g�`:F���93������af:���]��Vmm�/��=%�&iE�B�ɍvN��v�:�y����'x=X7�.��.� �p��g�̯�G��sA�����/�x�$q�vް���B�:Q�4�\�S�R�V&R��ƌ������PU����o6���S4�Aa�z��)���#Ŗ�^��7�/���rAAy/ʸ-3��V`�{����/X�?NUz���x��ɋ\����D�lؼ���Lܼ��cV����C6q>4���t�w��Ŵz}bz��OE!:�7&$-�sx�Ɗ��mg����ʊ􄐔�c��ɨZ3I�t[�1�[ռ��|({`�|a�x��u<OX8�ע���ݑ²MsP���ȹJ%�
�&��F��W=���;�.�L�N�5{ѷ83S�����¬)�D۳eLs"�H"{$��'I��Ju~]"��F���<p�htwZ��[dΎte�s \:���Ã�D,�^���o��)�a��s�6��yN�&���~�s+n���-�FW���ۭ�Mˆ���H-�
z�郁	6�Q�'u���wF��}N��}���y٣��6	C,�}�+z[�[�����T�F�I�������ҴTY�s�h�ڎ`�[��S6a�D976L��437Z˾WQ�^�5�9���ny��N�:��'���P��� <��ʤ	�ъ"u��G��?I�j=�1a�<�-�<��D|v�|��Ƽ���d�A�˟}NX�2�,�Zaւ�/���	}E�w.�a>=��l�
5����k�kD������n�n�f�tX�]խv)E�jF���y(�z�|w<f��GF����02�e�E��bs��g��3׹\�=e�詑)���'؎�ƻ���'��`��W?1�TC]�N�d��z�s?]f?8�X�z�F��wfNS�ǡ���j��K�1��=�ϫlU�"@�.k�?�p���x蚥�t�p��W�3�Öx �,Za���	vO�7�Τ���0��Š��.���=�n�����m����|�Ol�8�����b����́j��A1���|��y��醇�S:��$/������~A����~���#���������gݮR�X�r�G6�ׇ�������ǻ�X�Ԟ�y����~	A�.��֢އ���b�:��צ�}]~ͭi`���A�����pg�c�l��;��V� �x���[��ͭ�R=|pC]|��ڧԓCmG�q��$�4�3��]��E�ɧlh�^V4򉮏��8\�x(\aW���P3t��[���Ӯu��yt���\��ٻE����`3�Zxe����0���V�	����d��s����~��(�� g9U�|�����nʭ�~`��v�y`�P
ܨ�j��!?5��е��.�g���שG{�"֞���fކ�߶/}l��A����e	�'����&�2as�t�������T)Rz���g&b�0(e]Ϛ��d2�a��mu[��?�~��{��#�-�{�1k�.&�'�VfΛem�����{�����ȮBU�ߢ�u�4.8ސ_� �a�e[��:�1��oZ�:e������2��`7H��q�H�6^���O�  ��_��Oюח�0ʝ��t�R:6�O!c��-��>�0�Ry��m�u��sN.iGf��ߙ��8{`:���h�U)��R(��~$58 B�ݰ7k�G>�Oo�i0���\���j�?�IPX�Ɇ���E���m��=���X���a��9c1���F��<hY�2q�߉TXZ��2Uְ��L�U=0��g�إ�͆uU��58u�3���!��sL	�@���BՇ2q�Xcҵ���]�V�)-������n"����g��|D�ؚhV���?��5q��ϗ�'��{^#K���/}�mU����sۛ��N�b����q#�P��s`�D���X��4�W.�ڤ)���M<pe�"�f��*��#�i�{�p�R����DR�!�6�#�t�R�A��5�%{Rf��-�N������O�K�7��M�� ��r"�8A��p���<�s���O�;5�~*�+�Է5�3|b�|� �|<�о"�&��p��7œ�{�;y��Φiץ۞�m�+��0��Jz�P�q��i��ƽ�-���;א0&9*�c�����7L�4:�nXP��n7��v/"�������O.�i��ʽ�6�ƍ:�G��t]�۞���T	0?|�y�~N*�Gk����C@v29��oP�g�&�4�ݳ�T�D֩k��q�[�x�;���\�+���R���"E��b�h��>�jr�5N';�����|�:�BL�i<�U��O��9�ʆ�p�_�s��5���Rť�d��eHͨ����_��nIH�4�B�ߥvP�ј��O-L���/�&^��'��V����*��x���H�Ǚ�II`��"�]��c���	��
`8�j��Z�����g�;��z``כ� ��U��):,�ȺA�)�i8�,��˘N��n޻\�Y��z3�x#L�ys/X�f.�Ë��|$J���(�c��U�U�ǀմ���h�0c�.���>�I����Ŏ����xn:��9�%3�卼n�P�7m�eSγ��`k��`����KF:��쩪cG�A��\�cb�I�<h+W�OT����o[L=ě���ޮ�D��y�O�u�G�}WrW���&��P��=|>�A���	�� ��y�����m����3Ù8g����F>=/�
6҇VUt=Z�O�4���9�;����[�箺Kv]~�Ld�P���?�Zc�ku	�.�����9B�(���ĩ�!]��a�=��WC��di��n0��ids���\�9�u�k����r�^���wr��+��XW�eA/r��4�v�N�ezu�o��o3t*�н%90_���j21i��ktm�O���!̭�
�6��&6-����)�b�.:=�	�y�(�~�	���57�8����������S�+-��#��)����Ȁp�����1�3�y}�B߹QǛ�zn�����I�#����~XPA�O�I�/X�v���mcm�$?qù�
�M*�h.qƏVn���fu�e�}��b*c�=��&��2H��I��N�����f�x��7��/��o�]�w�z ����8�:�z#�Z@ABi����\�K�˪t#�*Ns�Or�D�S6��!�S�PH�����2��
�H�x[E�E���ힹ��廹L�.�"{�N#�œB[�C��\�5�݁�W��K�W��wWc$�����hkcD����
�6�N�HB�)����|$z���b��[����.�]�kP���T�A(R�v75�MIF��0�sX6��O��cS�D����
��> |=�����C����{�<��_����V���!<�mol%z���s�U�ow	�G)A�W���%t��v��z���o�#k]����[�+��ξ�I~f�b���7��d.��A8�Q,�ߊSL�Q�����d��ڃ�7"s7s����_ZԜ�A�9� �}����I箈��9w��l	n�l�law1��d��;ٶ���.9�ޡ�{���#�C6�������8�4���Zd��������q���z~�`�~��9���� 7��=����r!6������UT��p�v�&���b;:�Cw>6à�Z~I��Ri�%�x��Om"���
1�C���E�qDd���x�N����Z�c��BԍcI/I/`K�� Ļ�lcq>C����gNMu�y��`�:�ʡ2%:�="��;����'�>�d�ʨ�U#+�b��y��#�܊��Qf�<�:%���m����*!���ĉ��X'ߚ��AY�d��b5�{B=>��W6Ot=e$&+��J��.^yF��wn^�`�t�Bb����]������I����?+�R������������s��S5�o�D��Y��S�\��c��C�I;6����=���a�'��<�Y��a��ٕ�"���qw���RԺ�p3+U�(ԛS��U�J�r.�;5U�qNs7H|�Yo;M�3����Ӄ��"�*��\���7�����|>=�������{�Yz��5���ךx��<�$ �C���/���r9�;��t��������5�1\kwK���{@�%y�v�)�C&�����Zz�a�+�C� q.=��:��d��g5B"戝�ִ��=>�yf���+��%ޭd�J]�}kס�6�v��ym��*:%f*dx;� �Ǟ&�ҟ�3c[����AY$5$g�b�[�gO�ky�d��'o&%uZ�u�t?s���zaQ7!ʊƭPB~k;'�j����-F��cjj�`��j��Mp�x��mE��zפ;G�>��2�1<�!t�&�d�箈A���N����5,�zyYk�2�Ns�
�*��1�lQp�1�C�� ȸt��^�7	�d�����ɗ�x�5�Ô�p��Zuш�~��ʅ�a��S�]��0��ШXV��P�Ƙt���2�M���~}�L�*����7�-�v�%J�,/1C�J}�\h������@܀���Xו�;֝EOZ�/�`!�z�z]iu7�%<�)�E�x��8y^�\�.-���{~���ީQ�I��ݭ(�T�<
t�ӳ7(����g>��5��i�@�==tjB��]���L���v�	��,�13�*�IQ��3�շ/��Тow/i;ȫ�7�L�F�o�fWCs�A��%�����U
���D�{�[fhLMܡ�;	f�6���j�w���e�W��������(E!U�Q�	��BM+t�d����m���S� ��i [��$9z�f20�mYJ{i4�\Ш�9�v�!RÚ8&��\�����B ��-bS�b�3�v�Kl������;y;��U�Pq�.�%��u��F<yA��T��	2���s$��%[E�,]M9}*AMn溷�:^]v�j�Q��Ne�:HƜ� ����-�yi���:�SZmT��WR�l�A39BW���>m�KR�UV��י���U�ou︪��[� uJ�c���qDIE��_lu��z��:�
9�\pd��<�#�7�1���@�T�5��x�z�ͺ(_9�Lzi�71��p��­\qp���w|6�H5�|JAq�zXWz�AsWF�$_X|mcRY�2��κ`��P�"���mMic<V����v�iiUK �=��e��ol=4/n�M΢��Mcu3x��(R�:�t3a��fE�j��MK�W3Yfc-���s���\2�Wc��zM�h`<Q�A��.�ƬP���gi}Y7�U�v�Ҁ��uP�]�Fq�VT���Z���E�ސ���������
�ܑ�������+�=$�z���eI�3�6M���������5F��яoB���:�,�U�p8S�@�{&r)��3�ۃ(o)k�J�Z�
$��[|k���ዶ,6v툡���%��B:�	�a
�K�������rYJ�tM5��]5�Wt����ub ����K�;{���~-�!���[�ѝ�b�SF��ۢ�ohWN�B���8(�'+)�؆_:FN�r�7z�V�:ؖgN��(cB�Lt��M����*ݘ�ٻG8�!��㽋����Ӈ����U\�ݐ�P��삫�Wo>���**�л�� ��0����a�!u@���;���&�p�Y�z�,�)a7ww�^��w4��:��#���X��,��s��U\;��U���8TJp�j4�uf|�_Aj�>�ӫS��5�M�;�)�,w��w�>ḽEy@�S,o�(���Cwp��kJb�UGL�ѩeI.WZ��j"�@J��u��A�S�xM�:�;E�C 2o�����eZ�`�7oFY����J3	�u.�7N�$����eZ*�a���VCט ��Oo�1cü�ʛ�L�:IR����w�1���A�o3u�چU�X,��q}�#{����tk��b��>ڔU
T
�z���i�Y��QQ����	�����:�)��
((*�q���������������������������E�P%KM	@�U��TRS��D9�<x������������~�>��y&������()b��3USS%MU4���-QU�M	HR�v

JJJ��������J�"("b��"�������"���-SHQIC@�DD�	��UAD�4Д�1RQIE$KKICT4w�]D�%4i�KCAB�44,T�CITPRL%4%4%�D�����J�PѣCDR1�R�RRR�AM4%!�]@�DAݠ���j�� �߉�$�W�������.]*�5���Xc���G�˱����٣ V�q.��3+����NE̼�[v��z��z�=n�������U�r�'1����c~Xq���,"ZK�NP�xi0����,o\��eIb��0y��(�4��s[ʝ������)`�����y�T'�6���0��I��G1���j3ԯq����]Y�/-��+A1�P�ZWB�01����)s����y��rv�:�u�����yM:]����6��'Z�=�~�(p��h�� >�P����s���aK_�65�)�Cu^���{��&V=�P�9@�*[���^��g3�"]぀�	�� a��s=�r�^>)�e�k6]�s��
���	���3.�=���~�,�)�%��e}��J�~?���GeԜ�/�qQ�ؘy/�^���Ӱ�y^szA��8!����'[!qT��W*ڱN�1�"�S�kW�T�8�C����̟|�U���â���@_?T
��B�o�E�ثA�v�)������{Kƿz;k��0��E���#���~�>�k9�R��=t��<twt�L�׻pD,�R�Ӕ+lh뇭��.b��~�E?���0G� h>@A��?}�]ڞ>R���?Q�}��wXt��1lr�mD/Q�ljԄ�������P�dS\��f�p7F�Co:D~��\X?�<v�<,�xgL�3�6��˽��-Gjz�i�Mom���<U��o���b��9��r����,R=����,/��:�$C��8�p��޽z��������?n_���<�~*Be@ZT)=��vzw^���i흡Ʉ�w=6+iĚrwWVF�bB��Ga�j���X/�_���5B*��l�>���}��x=�� �	�h��݇�X/X2����@^���y��|k�7�Ru��d]`n�cELy�W8�E���Ǚ�ɛe��M�(�C4���b!0<�%�n��"U{��<��(�a|�Qu��Ll�FS�tOM�R���۷�>�^����`�̜28Bn�L�7ƅ;JUzʮ���R�N5n��-sU��"a1��a���]��>h�a^R�!����8&%:��,.Z^rfCe�k�I����0��C�Q���X��c�qͥ����>���o�C�Z��Wn�:�&[�骬��[yzz�����k<�8��{ �%�^�V�Ϯ�;_���@A_�s	\'�y ���.��g�����b�4yxƉ�R�����I���u>_�O���i;r1������gu�eW�y���|��O�#	�|�}:����@���{�_��c�^��{�>�?��9��U�][�y��o��wb��;�H�޻W�耪��ݭ�V�T�yq3����ɨt4�X����V[��*��]��4[4YN�U�Y������o�E�l�uS/��'�E켽H��6���q�gv�J��Y0�S�U��K"��6/�	���9�*=w�u�]������}*�t��L��t���?��?O�O:a���xQE�K�:�,ް�ޜ����H|�=�gXJ�l�<���$����%?yh��~ڑ5�1�������X��Z��[�^mmv.�֏���Ⱥ���od&iK��u��9Iwy�R����E1a�|>��/?�mZ�6&��u3���.��ƟU Ͷ�j�����3�թ�zǅ@ȧv0!g��gT�:+��u�:��y*_�-��n���C�	M����њO��{߅���L�W.��B~�p�3a���wB�O�D������Ed���'�Q,�ߊSL��Q��z�}ܞ����M��ڄ�}��/���� kENǡ������X���<�:"S��D�Y��'�6z*S��ۦ�v�m�-���}��,v�W?�1�,���;_��U�3�]@��֭&�fxu�`ᣕ�b(�!�%p�\Ú�LYz����B=D&�~���R�T�Cw��]�K?��r�o>�C�=0�-w�1�I�ߑ	����9tK�?KE�>(���E|2�_Ѵ��K�b���չ)��0�H��tⴭ�7Zk_j�T���Et	w�ۂK��;p�y����øe�L*m(�QUq�D�����mg>-��m�\�.͊a��z�0�i��(��H�:L��nf��k^�t�C���^^ �8���G��SJ�
q�<2��vi��r�k��Qx�Xä������qxwm|g`Ku�V�3��)��]d�&�ݙ>�����Su�k��I��b2m�T{<��f'�mbC��~��>GnpU��DM����`_9.���K��M�j��K�N\N��>	)�X�N9�-�����7�W���m��~�"�\g�\'���75ǲ��3d�"�/��&�4pᥩ�(zQ�㎿�h��H��`�v�
H~�P���k%���Y�B�n	�-��C�sh��.��]�O�=�ߕ
Z~�V>�e����P(�4l0ꧯً�1�*��1l�́�>��#hoI�d��3�)K���^�y��CdS����xU�*�#^X�,؎a��6ܟ ���΋cn�pB�����[8#�y���,Y����Wy�Lu��
����+�(�Թ�Ym郈���QXժO�u�N|-@�[aG\���+�vlA��Zνq���2��u[���,9�2���#�=?ܨs�����z�W��M���U1/�L9�O*�]��٘yv&��)K��8q��A�*�ˀ���/l��1��\��xa��O�١�cjUҙ��H��b�.��0W\J����l�sof<4#��I�7��ͧ�[2k�7��F�λ�����~��>��~  <�^t#M6������^6�I�5rq��\:��g�"z�"�wғ�gK1��kF���i���%��1ܝ;�u�IP�r����;"�t�PO������=�4�"�1�P�ȃڬ1Ke����%K�t�L�c���c"��Ɓ�3~T�L���"]|��O,����noq�����^�����A}�%�ꆛ꒞lr�d]`/�qsHӱ<��ة�q��9N��;<�æ��y�����^S�<hQ�a�¬���W(��*K�e����=��=��qJX!Φ I�Z�Aa�����6<{ʠ
j��z��qc�Z��%�XwS6�p�M�-T�png���Z�t�HOwމ熇c\0gAϹ�0~b�-�����д����ە���ߝ�b�]N�����=2T��>�Ow�a���(1��%~��r�S�k�ʘ2��e��1�:v��f�o.���6��ITމ����(R�sqe���d�P�yP���n,qaw��)c`,j�(��uc�Y����v�r�
�^�0����f]���8:��e��xT?�����!p`�x��S���үn�k�����<��:�-qǔ�-i]1�FK��ئ�B�Zƻ���Η�Z��E��֗����I��!��ϸɻ�*[g?�6J�94dN�/��^w�s��|�n���*��z��^�<��^���~�?��3���x{ð�+��*�n��P�8!'�y��訶F��N���szA!�%�].�Z�> k��Wql�$���/5��!q-3���%bO~B
2��d�z��΍i�	-}� ����m��g�j��Ւo���.$�psg�K)q�tv��Ίx�v�! wr��Xgo쪇����d����^�(����q~�XnB�P�`%G\=oN0�skb��t�o~(��l�*㯪�}�Jf�tz*��Rƒ��Mj��ؤ&UiP��+���y�̤��~xY�����h|�}]������X$^׸4��<���Yx�����	�T.�9�[�ǔ��ng�O/w"q�~�s;�'{���r�`pO _H�5�ޙI�x�K"�s��K�m[����{2����ss	P奈<�ļGܲ <A| �vO5��(�a|�Quv����L��{^��ތ=˛]N�AGNY�6�;�� ���Dp��^�	�o�
6҇i��ƌu=]�ln��ټf��n{�J{G鞳+~�F�~���N��Yy�]�6�@D�|�|W�0s��Cv��2�,��tI�mS;ZX�,����uW�85�������&X�#I��wZ���D��[صt�R!���⎄��b�95�k6j	�ns4�L���`��M�x�3t����NC;5�g��<�^p ?�{�w�)uY�Rq��Yy�HG��·}�t����=f'��UH�un5��Ý�!�>:=�XXb�.���z��B��sqI����K�z��5ҵ��A/r�?�qk��'�[�A�Z��EG��[���yoT�~�߅���G��v��t�+�T��(�|��}8��Lsp�Y��$?6u����W���86�xr��҅@fq`�xA.��_=.��}y!�/a����$8���F�v�����1^��&�;�dF6ϝ8wl�tK�����ϥ�\W����ma���/���afź����D�z����H؊��΃��C��]�z�oE�l��|����y�c��k͖`%�Xu%�>�O$���R�0j�1a�~�|�&+�lU��^t�O������cѯX�/hLU3m����8��y#���8�����)މ׍�q|�t�8����z�6��3��5Gl�m���}�O����M�9J���4��+�P=����Τ���x��8�}�%ש˼`f����A�Uss�	��d^�)M2<m���5���=�tz;��ۋ���3��U����b�I��c�&)w�jp��}''�K�n�ӵ$˛�R0+����nTb�l��W���tY��,���󲋡e�����[Q�'6��sj�$tj��>Y,WD�����/?�?�{�ǧ0��$����oma�_~O�mbO�H�6�sȝ�����<�DJt�f�z�k���l�4ب���F^׸��[�FSSw��q8���s���`}	��?K�H�w��s�1�:G]�:����K��5�S�DRr��E*�*��	�/O�������N�΅z��LF�4�>b'^3��ʽѷ{�l7#Қ����a�Y�|�^Ť�w_��<����H��,8}�`K2]���/��������<1/S�4�c9V���(�Z��a���z>;�t����ƚy^|�ٜ[��>E!����|G�/����7���.7�zz�l+�)Ͱ�!1t�r^�S5����B�i�d�\C�Y���<���Dud���+���������Ta+]M>;��h�W}���h�sH/��:�;t�k ��c�b>05�<��3���_~1˵�vQ܌{�}�.�����m���m�A��0����sP/��j���B�`���b���G��
�:��Y�/ڄ����C*^�4]�����|����ʇ)i�Xi|D��`������y{6���tx�?J}M7ܺ�K�fs�:�UD�J+��@��;9m�H�����W�p^��Oh��.��T!0�4�T�m��u��%�Q��m*�uk:u}is�"�\��
����Ӝq[�rk���(�3�a�ѓ}F'/v�^�������?���Uh�@�V)C}_�b�)��6}�hM�<�INW�}��0b�*򖟷�������8�le�~�&m
w�N!{sqm��j������Z�B�Ed����AZH��
�d�L�Θs5���8�|u�N����%=}צr�TV5{T����A<QvQÍ�������%�]X@U�ذ��v���O��.�9�I󵮝dՓ��S��l���Nм�����2���Kο!�P�bUԻ'�T\:��| ��A�u0��Ix7��f���c�.y��rf��D�&��'.�$�EV�ſE��ȶ�]8ށ �67;P)�W�>�*���C����c'��/L�O��Re����)�ޑ��\���oviȕ�ub�a���ACDsH�-��4�#�E�	eC��4�꒞o��(�T��9�j֑�0v���_SMH��Z�a�)ӹg�8{d-wd��<�_czD��L*�.xn�Qy�j�t�(�®�M����a�z��;;Ϛ�d<��|m���t����Լ몞4,��n+��w�e�B���/�Az��n��&��|��1pT.V齑qؒ=��5ܝ͟�p���^.4]�Ok�
���s�z��ַ��UXv���'\\�]�APTܧu���$G�j�)b�ת�4�n@�D��h�iV�ҧ3м=����k�ɾ����������y�����!
Yܥ��<d��
�XH�{�֮{p��P �=D-<`c���i���!j���5V֮���úP%�6�r�.��~)����\�7�4�ro��<5�M-e�0���M���2��3�����C2پ�a�C9*�˦��;N0��\Ys㾌�2%����Y��DSfC�r�}���>�`��bmՁ0����v���,+�Iz&���l����N�d�΢�=�Qǋ\F��c<���x��&H�O>�����푼�a��/�w�'7S�!�����:�Wי֝��m�:L��X%`����!d���Ts5��Ox*8�W�w�	�e��ӂ��k�B�wd�xך�)�t=C�����RfU��5�wuCNYQ4��U�޿d?��X�9�ז����P�~J�{`Dt[1P�)���y�PZ%��F�u��[[�;1����[�g-����D���)	�J�'�J�vMՆRf�YFo|/r�}����MϹr��,�J]"���/�_W�i�S�O�Jee�S���(9�	�	EP��t�>��I������7q�|n�<���_�VgR+��]��c���q�S�	B���d7��V(1%�Hd�b3���e"����	�e�NW�-��42��B�/�[U4��̣vx�(�ne��Rwe_e�K1�*�)̼����[���M��opY�δ�;��ǌRv
�3�W���u2uV����<�=�kFߕ��JNͬ;�F6gc�J�Zn`�����q�Xk�.�׫mA���Բ7�F�sޒ���·�HK�W���=wl��=z�KT�>˩���N���I��Y�[��b�+��ި���՘��-�B+����<A3=g#�f��lZ��sa�����U͢���6�I��8�ب�n�vWi��ݦ�K��Ξ:�%m^.���MK��;bd��y�5���jk��O7�ƞ,���i�*+�����6��8��K:�9'1����#.�m�ѵԡ
�����6V,ǡ�"�t�e�i�8�	m��)ྙD�>�N��>�o�8p#�JX��a~;\�)��MI���w}"����N���h�f��}pf�C��.��Gp8a0�R2�_uu���e�w)n�����(����1|�y7�<���
��sF;eYY���
=�kVn��5(#�opr�v�\e�,N��K����.�=�J�_aV��o\�oP��0Pxp�N��W���.�9�h���<|���[�a��M�/p������8�pN��V1�#����@T�LBB��M���Qr����B��T
��U��V9�u��q[�#��t���o�D�{'3meJ[e
�=� 3Ӫ)B��.�&s�f�sY���=�f[�Ά��JsM�*��\�T	�O*��0dQ�=)LA�wm�[�:n	Z��Sy��N�+����ʆ"]�����fp�A�b{��*�V�h�̣�dC&��d�ci_��+-�Kg׸C�����Je�S�����5���C������q�'	B���at��_Jv*>�P���>U��oc�!K�����Z�P/��m��j�{Ee�Gt�E�k�Y9����ޙ49�K[�_t�/\��ٯ�D�::���9Xc�J���L�������;Ι�r�9*����H�LA��i�k�|TZv��m��qk�ݘ�%����6���"�:5�:J<�Wb���@�e�ڼ��9i;�n�����a[�F�NY���WW �6���r�g	�L<����>{�&�ⲣ���̹YI�o�q:��`�[�!��m:�Y��c��uE!���t�ǵD7�ǜʵ�d-+��9����-��7Q�8L֠ۗ��f�o�݋����o&Jb��\��m=�	�x���j�4p�5��R6�M�6�70=�Ɋ���^��$V::;7{��5ܪM�I�A�e�T2˸YI|�^��5ҍ"RHD�J�E�+�W��OǷ�������||||||~�9)DB�QP%1M-5EP���G�zsǏ��>>?_����)=ΓX��A� N���D�w.�mEPҚMPU-�	H�CKОܝM%5T	�Iܚ�4��� �4SC����i
��B��(Bh�+T�P����!�����!�)��Z����(�J�Z ��i^���:�4'{!A��)iz�]N����;�����(�)�QABPRRą	K�C^��E5��K跬�(B�{�/]���f�;�]�X2���̼o��Ufb�t$W�f s��7kW-v�qĖwlֺ�K(�|u\�]�ղ��\���f/���K��Le!�Kq~e��@J)��%��Ox������6Yf����SS��FA�F�_��rԘ�,j�����| "�קze'Y��,��n�c(�کg�+��c���a^B2l�l��|�ե�Bu/���b�z���ey��_EL+۴?,�7�Eu��9Ҧ߹�;���R=_��R��uZT_��N�4�B`&���D���!����<��b�m��Z�q��=���O���$尅ҡq���>��-������σ�ɂ7P�F�[Qw��7��{�WRa�Z�P����~�2U��zY�KӇ�7 8��kuX\Su���Na��O����//��%��N�4z�X�kXq0���%�^��9���Y��-��W:�'�3؆����	� A�
a?��Q�������g�}�&!?K�(�[���hi�465��]짗5�)�����΂��4B/0����`�����.���<�U|��	j]��e��މ��N �P�`�����?rio�x�4,�>���y߸9�ƅAF����ļ�g��a����
hq�v-��g�C�T?W�!O��a�~0���Ruw|��6c�`��ۯ��^mNP�8�hY����R�n����u��o�;�^�L4$�Zj���u��&nV��#�&��x�k.\�i�vHm�d���ŉ�j�4Π�vi0�r�W,�p�k�s ���zZ�y��i�|/������)������~���Ζi�vJa�䲂�K�y����Zf�aqf�_��>�^}��_s�t�:"�h�̽O�&�Ҟ�c�)f�;(1�S�RG(=f�'�z�U*G"�CNd���)�]]���GK�`�y�EǥPUX�+ڊ��)��)A�Z D��J��o��*�ws�uYӰ�o`�:�o��|wC�f{D��p�{��E�\��q��K"�$u{ͥ�f��ו��Q�L�k��Xx�^YJ�~�`d�]�*a0W���'�&�2��ow�
�b���l�k�b'����#)��;'���g��>�4�R��&42+/`Ո�*N�7
��,���r%*Rr�)�⛤R�b�a�@����}��l#�&�G�+�D�gkx�����R�CZ����)�����Ry�iR:�M0<��:Х1U]w��Q/�t�<a�#_���|9	��z��	'�7o�r�k�2��Z��a�~����F4��S�|[
���#���t;�wd&>gat����@�\�����6���!���݁�)?5��o9M�fS[P�ƫ�颤w{��5u(_{
�G�����O	?�&۫�,��V&;h�CuU��#���v�F5ǬgJ�שw��L9�w���*c1,nA�{Fi��)w#�noqх����1�k�X��E��Y�W���j�v�7c{�"����?~�������n/'�Nk��\�^��wf5�����~�.��z]��}zw� Ł��{w╎ƾm�7Jk5�G=��ӮF}[��wˬ/�uq"2��
и������~[���P#�*BE����x͇>ޞ��pB1,7Ĉ�	���1�W�z0C��y��x���Bz��������^>!0q���9�hM3EڀㆽS����p������1CW=_d��>�������xc�ܶ�-���Ǐf�<a���N2�õ5�'���Lj���E�TwW��E;ƍ�2�`��ľMG��]y����4���Y$5u�f��ʓn����Sy�Yׯ��@�~r^��K��iFz�6^�TNH&򢱫T ���w��ڏdL�'.tGf�O��6/Ռ�c��eEÚ��>R2���hLIvލd�'{a�R��]�'G_Syu����X�
P���л'$=P�4L:��|�p�[7�(R4��7Afg1s�j�Y}��\3`]�[��DI��N�%B�ʿYN3t�	̋h]��K���D.�:eG_���~�R���t+�p�k�tji�d$)�W8�^0v`��I�#�U��,��u`ڝ�reӝ�٩�H����tֱ����c{�^�:c9��F�W�M��7ڌ������n��4Q��cY+���)�_>ef�|�o0W�:b{p���C�c>��d��g%�I����LU��E'�Ɓ[����&��}2m��GM�׆Z� F4��~�&�}Yv��꒞lSl��/}�ubs;��z��~Y�o^��jI�G��<�K�sˇ��,ר{����yOu<hQ�)��es�IX�*q���:�+�iM��q�Ƽچ���#��cm�t��q|�xгyW��)�)텞��|v�ۼ�\b��]�H
�X�}njp���i���3{_��	M���ۃVWtɬs�cr���2q�XzV�����*��O�؝j����8��2�2�R��+��%�Ŭd >���6���՜�l�k���(�����轆s�6�@g�׊��p�3'���|,S	��o@�����͈�nIa�q�/@����;���6Xo]V�=�uY���+�L|<���_=+cXX��do���#בe�z!����~ǻ�S��3[.3�v!�����'<"���4M�1�lg��`L���C̟|�U����C�ɷ'���i/���gPh+�q��V'7��Z�fm]I�@|�"��i�n.r���w���dp�n^�Շ>5��Q�x��9ܸ�������q�Å���5���p5T���S��wE�ӯ41����t��fl\�L�����������%��U��܍'S��zd'�/|�B	5~`�����1p��L�0Aaä���KР�<lFqQ'o�]m3��=LmU-�E����ֲ�	Q��4oF0ܘ�5�g���p�ٺ��b'���D����h��yy�\Co+�qt��:��g�&UiP��3�Z;�1��w��p��_�w2R�e�s����X@��	}^!�(�nBg����M])��Zj�3hw�w��b���zX��^b�k�;���0�D���.p�nc��_�e�:�S��%��m�卼rK�r鿖j��̜���������2D�U��0�>�lw[�-����tu����5%���v�;Nʁ��-N��ޚ
/�����	���?!ӱ���UQ̛�gY����Cyj��iOC�����+���rq.�����0t�Ǭ��n�MT�n���,j���*��QI����8Mz�лUz���s*�w?,��� �C}�Z�F��@I�?��g�{�=`�
����X�Ķ����ɜa<zV��^��\sO�ܳh���)E�k�z����9�A�o=�u�i���0F�w������o��f������:^=�X�L��u�qM��WX�t���I��v6�`u�jO���odR�lM�e��}C�.�&����`1R7ה�#�c��FЯ�����=�;I.xc���\: ��v�M0��o Vt�'�)�eO���ӎ؆P�se[[	ꩥ�u�w�����6P�L�	�ah_y_榬��`�Y�?xŽ�Jħ�ZΝW��_��E:H��@��I�Ũ�Ǟ� 円���e�Lz/#�H\
����KxNl��F��4�����- ��u#�����7Muc�?���c�څ��b�L�����ʚ�᤼��e������%��R]����~h���k�>4�;�$=s�ŷ�otGO[�2:9�FFS����O^��i<�3m����8��{����8�̢��ؙ<����b-�g���؉|�]�ܣ��uz�J��W�����b�֔�tk-B暋��ͫw�y���R?�;����/P��6�D����C��\)� tB	����zX�y�Ɛ���6�j*���O�p�5���Q�����<�ʏ��	�͉�o����c+z]F�y��b'_�炈��t	c�Mmb:皜��U����	�%,�-�*��*��ku�o5K�[��v�_�����n�[�B���~I�d������.�=�0��͌�f�����l*��!����x��kð�5}�֞���,��2��r
��n����v�������:�4�9t����؅��|~����ὖ�]v��{��=��/��&O���O��Rr���ث�sQ1e롆ϣ��wfsc��ji��7H�t�O
�>�M�1���{<�_N���Y��A������T�M0�%�*s&c<�{�Շ�O��ty��Ð�����=sM�'9^�`�(�P�kz ��{��x�7�6�q
u���&���dC���w�ܬ4~]�A5}Btz�u[]�zR~l�H^4����O��3���������&����p&t���У�e?�C��/R�/M[����h-�G\�p�ܹ���n��uy��W4����Y����c��|QӞT�30���'gn���ݐ���N���a�'1�^���o�<	�7D[(�ٷ@Ԙ�s7f�`�*Ũe蘾ub���b�m�}y�vo4��~�.�aط���A�^�9��
n�e���֥���8Sެ�bP��/�}��9Kכ??^_P����v��8�d�R홌o������K�d��)k�B�m�:�߰��D���֓^��f<�fկ>�9�!�{����/�A��ǅ��x��M��ʸ�9�S�����ɃX�9I���8��4Jړ�U^ qm��,�q���W�x��E�����V�\����t�+���Kj�)��E��^��U��0LMK$r�x�Y.tj�aݗ���v�G{G$������T��a��7�p2�g�ٳ�h�l�NT�ǘɁ���DT����X�u���6�su5�����h��IG��P%�%Ռ�c�ċ��s[��
�x..9�KP����҅W^��V���1��D �c�|�T1*��0�;qls0�LK�}~̳���_8�I��_��S�^��#�Kss�d������JP�&Jy�]�٦�[B���kS;K�^���fL��t23k����Ypqp�V�7���*�"�6��"}0ut��оsG�g�/�K֙�NH�ֲ�!�sB` ^o�K�5"�����b)�t�	�^�e<e�s �|,�;�0m���S*/��b�pe�R��ȓ�i0����ڧ�6jM�'���4�Ǫ;�#�z��	��Wd_�ӓno�5Ϩzd&��%�BN�3A��j�p��l��4vwYJK��c7�V�z������^�<{\0di����.Ӧŧ�i��g^���b��M�/�W�2q�q�Z�9/LUG0��'MV�A��_tW���xR���S�K��b�
�S��fvu��Q����{훪	cr'b���+#������z.>J�h�69�	4�t;�nU��*�&��B��݄��;:�8����@����N=��Dgn�:��Jԙ+�ڣ�^T��F���W���9�ֺފ�]R'&����/38���@u��ͷ`VW0M���Cæ��_)$�71�_d�}ݫ&�t��=��B��*�%X�	��|CM宱?|�3�em�<��bK���|�L2�t��o�3�h���AW���Ξ}�yw���l�6��A��S�dP���c6���|>���
�w\n���t��gu���41<���Gu:L�O�#c��$�<�;|�=c�l6ʵɱ�S�Mm�F�?m��̅�-B�z	\�+��4����:k1����^8����%���iJ�c%>�-�����q�e:��ޞ�ۖ�\`-~��A�Z��Rq����.a��S:hl~�5uIk���[XǦ^���lccj��Bl��BeBҡI�J�y�߲����ҿ:�W�3ݩ���(����Z������Cv(�������%:�%%�m��re�����k+"�=3�]!
2s�3����m�8f���p�範$_��BN���S"[�M��ط�i�H�7e3��:+�P{���X�a��!0X����*����*;E��E��vT���� ��i�ދ�����3;cr&Ҝ�Q�)v֨�QZ��(w�н��VLCՙ#�����K	�h7�h�糑|����l3�kj5�=�U�؄�y���iY��4�4{o3�sr�unJ�ێ���\ZӒ��0�CkWo+��j��� tѾ����&{�V�0�R���)�.��m.��4���D��".�]���C��[����u�˼�ڀ%P�����M�=\���$���}d�h�l�#ܠӦ�ZLI�ԛ'���b�2v�S:$�C�~��aͣ9e�*�=Q�b���,��%��Ʊ�A�ig�3*;3>��a�(������ϰ	�)��M0���k�*	{��+��Y�VK�t�6�Sgqf7=4���`�L��8��^aڽ��ٚ-�Vt�+9P�cS嬎��[��5��tͮ���}dv�y޼^�;���<8B/>����%�>O�d;d���N=�#v���T�q���d����^�����к' ��>;��y�f-݈Y�5R�}�u����$��Ʒ$>Y�a��|C�Z��u#㢗�J5֙Z?��v����.��3�����]Kս�mz�f��,;�YAP]Ƌȴ��4�����Y�7w��nN�Q_Xva�$s����������\T�h97QS���$v�����ƺ�}�!�«td��j��3�w=�N�/̎�༹OoC*�O��m)�1wN<���C9���ii����R�N/j)�Ѧ��#�Hb
���;��:Km�����Ú���M�T�K����fޫ}�����&W�j5�^�W[�D9���u���7
�=�Rܳ����6Z�Gi�S� ���G[���9en���GX\b��-q��hAH�����۽�:��)��*+&<sN,�&r�{�c��y�����	�oQ6p>U��j��/�{{�輽�(�I�w�P�}�Gn�d�MV��ɞ�cx������i6+�T^2mɂ��ݰ�`�f\�v"��.�͇�ҦK!���
�D��}H��W�=��7.�H�u�[��׸�B��^ڢ��[y�o�axFl-������/m�꺓�g����#���LE�)z��ڃ��JU�SlF�ӭm�}��٘�K���W����#�rL#�Z�Vq���:�uL,��j�F�������FS�ەϥھr�h޻�7T�w�E���+�/V5�3-+t��(����{��d>�:A�Qǖ6���S�l��Zg�:e1��/��g\9���xTӺ@��,௘�z�Sz�����J��W.��f9��zh��tYXJM�e	]�.�t������d9�Hѧ�q:���(���{�qҫx�w	66�U��>���K���T5�<#	㗻L�a;�[����h����5������D����o���^{1�%~�n�PO���6ܙ�f����`�UM��*ա�	1l]��ʁ%����\;��F9�@N�1��>#l^�M2��f͊g��ǽ�mJ���&����Êmax��/矪�n������>�=/x�(�"�&����W�Q̫xs��7osdg1ÊA��L�^<�-�
���c�K
y���^��׶�ں�
}�޳y��к.����\a��.�^����Ѳ�j!�/M�*��XԫIS�N�i-�(]��"�i���C��8�qht;{6�.�Z�@�)���+4D$�ѹNv2|h��s���Ɔq�w�j�������J�"��r"wr�>�;x;�5/9��Z�)Gfu�`i�*�WP�[567O���%Qm'B�v�5�wM)����T\:��y�A���p�����,��A�ӱϙs����\ͩ�'P�x:sg��r�}�m2b��h�/;��ھ`��[���q2
N�
�u1+�鏅r�J���;�0�ĦW$+x�`�Eku�wEʃ;�r�	��:U�zƼ!�(��4���)
���ˣ���e�ud#ܳ�Q��&��O��fͭ�t��ʸ)=������/�vm8��z���wM�"K�٦Ԡ���JJ��:��V�c7��T�s��a+�.ֆ���ƤÉQ����Mv习���<� |�͞�((B�H��t�RU%(�R��l�=>�O>>?>>>>>?^�"ܺ>@i*�)*�)�] R��s����x��������������<�(��)Jt:��a����--(P�A�J���)��(S�SHR)����4�SHյ��h"W�;��Z(Jz�Aݦ��*�)K�j%i�ij��;��j�{� R�THRҔ�4�4��К���tKGS�����*�-�44@P��Z����t:
M�J
_�iR���4�4� z�����w.�'�q��#[��d�!��g/;��Iū���T0NNa�ut1��y����3z.�'W�#_���~�ų��D|�����TƮT�2�K�`qw��Z���TW�q�yB���mj�hnR��oFխ��v-�=�V�ב2��vd��^�`�"���S�D�r�bz���h���#��	q����΁Ji��*4)>��g��<�ۼH0#��5æ
�^{���f���5Q���'��$�b%:�%"��F�[X���P��� ���f"c���v+'t�Z�z�L���5Ȭ�aӹ&H�I>��n�J��a�Dŗl=�d�\ӆ�fNdEf۲�Lb�
����F�W�86Ƚ�)�v)��-�$�'�h�i�,�'�W�T�E��C��+�>���� kÐ�3�����Ο�"��>��Rv��{/hΔ�\�o^e���>�F�����7H_rG��l=_=b-������/&��All���?	�$��W>���f�;�c0l �֟1���]2����vғ=�p�{�Ps:��e��=>���/����5�A�A|ǵƑK�r���BH4����M�^[N~u����y�͔,��E�uN&I��ru9��,���M��.��g˛z�n{l5ڷ�1	�����­ej����O.桰�]�ܜ�2;�!7�+e�;�����yؘ��14/��Z���]���,cL��y������m1E���lǆb��Kłk�+�uӊ�a`Ё�@�E����#���m^nU�T�;�`P��-�x�n��1W���Ю1%ڽ�]����q �/}���(t�m�pDTj����6�c<�wY�����b`��C�_9�fϯ/�N�v)HA���F���1��~�W�ԝ��־z7�xU����2�[ql��W>����iY��^������u�C��L��N��I��ꚥ�|h�
��>	_
r��� wN�nA��W���ca?��%�|��8���ߐJ+��;\<Û��P.lD��͸���˛�5�7[)b��ry���� �Z�9BeV�
W�U�Q�vL=5to���9�}�W>���!��m	��i�����M��gt�?�N�$�*�))�؍�`�5���;,�����lv�tf�kF�kzS \��T���a��e�H��*�,�O���n�I�jζ�R�$>h�ջr���Bvp���"�p���˰F<9K�!��=L��^�K,���<2'O���!m_WZ?�ץy�A��_g��K����tJ��b�����r��8yg:����N�] ep(]U���y,Ӛ_�-���fmJNO�em���ړJ�+3�PL���U��Ƌ*﫱���<TL3�?����������(dcmy�Xg�������}A;z���h��=|�����VX�!�����&|{��Q�{�yz0z����Z��|�� �/j��T5�ơ�ʉw~ȋv7|��t��__k�����vT]m�]��yP��'Y*K��c6ְ�^�ZT�x��zA�繁<���zS�����2R�e|dU��8���{�PK�)~a��r:,�[۹L&13����XJ��w�/�����|'묜���%@��6��E�j[�0t�.�eUF�YW��&�u!v�c�gR�g�<h����߬L3$�y�;���"K��nQ9���8�����L�N�zd�l�sW��~�y�4,򟚟+"�;?z��N�:��l�͎����K9��i�\�z�`�8��_����~��ϰ���hd	�B,�{t�r%�:�J�U]���&�V�ĳH����U�z	\�;�O�E�����R���ˡ���D��捷�6y?p��s��x�^izن��P� � ʆ�q��T��ь4\t�h��c3���6M�,V_U
���/�[����Ǟ�I˭o4�w��fK�S&������n>;A);	Q#��O�p  �~X)X[�6���\��;���w7jơŚf �Ю�N�n!��u�]���p��qN	���y��f3�us������y����&L�Ug� kh/�p�ώ��-����1�lq��P��R{�(U�A�,��2�W=Y���w������=d,,�Þ�%�b@����v%�,�&�Q)��5CnsrB���;��u�a��,4�k�FNc�S9|��!��'D>T�I�� ��>d{�j��l�N�ӗ�E�9֍>��-��u�m�FS�(��=��z��q �5�B`��_�)4���2�6u���f�V���NCϊ�N�X�R��g�=��ukĐuZTW��"]u�꿑��}�6D��4ܲ�&��'@;JH����Z~kJ]&���h�lݦEn]Z�M�?a~�`G�-��}#Z}思�a�Y�(_&�Q�b�K�	{���vSGLc�h(wf�~ià'`<`��x��Ý~��	�^us�X³��{A/r�_,b]C-{3}x��栎Գ}_�����q?���y"u|l4NZ�+:m��*�L�	�U�sSF�3�Q���}�>�kUϟ�L�zk�4s	���kNyW��1���U.���uq��c��'.�,�Ù�W��!��Z�kΪ���YJ��uˡ�c��o1�gM�u�Ͷ�I�|�s��&J����U�ѽ�L�A�޽�h��m�b��v2�6��P[�N��]�0�����$�y���0�w~'��~�%�	g��9�ọ��p��C�+�����7���<E`_y	2�֧�W$���ˊY��.���A�Fuciy��P�ǻ��-�A��]@p�y���r�$�>�����6-��q|�oF�k���3MoIa�䲂9Iwy�Ԅ��>�ȩ�8��,�<4�3���#Y�P��\��O��{e��297PN0,�,Gk�v��{9Κ�����:���r-�ёN�ŴzÒ�"��!L�r^|��M�����#!�+�D��R�j�ׯ#ӌ=��o�vgA@���. ^]�UDź�}v���Ge�e�9��Y�
SL�ʍ
�v��X�1>�+���_��]�S�g��^�e}�XpH�>��]Y'��N�%"��Mm`G\��p��cm�j�h�gwG<��`ք2�R�0�`c"�Y���=;�JO�!1C�J�UsG��������f-3��7�����^t)�C��/���ڏ��{���fh�OHŧ�3{Ư1�Jֆ��t3���*��'28����ή����3n�g;Z�$�lW%�%whWAT�vul��rk0���}�����ץ�|���s��]1;o�m����,k:�C�y=j��b�>�D�ڤ��3�b���&�ە��g߀����Я{Iݖ �٦4���a�Q� C��<�̵�N��u���U�\�vk�//X�ʘ��8TQ�T l�<K�0�ד��M"��D0>��?rG����A5}S�mH8-����Έ*~���f�����mKg������T{���6-ݚ1�3�C�x�}�vb�VHkw6h�;ܜ1;Z�U� {�^�s5���b�cߑ��O��֢���y�e�v�vCC��D�o������m��}��Y�Duf�n��I��]4;(��j/��P`��]1�1�4�.�g͝A��D��X0!���,z���Ft6'�^CZ�u�B�jQ� �k�>��J��ɇ7ߴx��Ǌ����� �-���*{�MQϗ�l��򥕼�p��w���E�ڦ���c[ݞ�4xٮ_@K^�l����N0���E�/U�z�6q�鼛�7I�鈭9뺷��y� �475%��W�7�l��[:y�x��,:O"�邳��Ѹ���KUtQ}�4��q��QX�䠧泰�O���'V�V��6�����?��9k+��C��*K��C����PM�;o��V��t� =h��m��;��N����"��qOS�K�����sS��g_U�x_�誫�k���Y�aU��U���>�7\V�}�WK�)�uc.F�r���:�t5hN�bz���V��4�V8�u�d㵳�Dg���?�!�Y<m����X�G�C���h��:td~�\�����(L�ҡJ�W0���8�:����>�ba�M�gB�&��NЈ}N�/dp�;%77;�I��Jua%A:��L)ҷ*��U
�S�X�Sh���`D���C�}������!�e>��n7�"}�&�"�&�&t�8�x�6+6�nq���<��N�o3 C�o��~�s�8�\;CD�EB}�i&�<,l���i�&)�u�൭h@;5�N��� E4y	�$<���˟�n�1؉3���:c2��n��Cy{Bj�BԮxj�Q{AcK�C		��@��`�i���/l�Bcl�x�o���:[j��M\�	yO�'����V�U�]<�o��=�W�2� �`bY��p��վ��m��р�W�/8Q�h	��oL�Z�N8�=+^ʂ^�K�[bu�[�ЏF����� A�?jW�0B�P���< ��a����uw��^�#�؛}/�8%~�ɑ=��kmc���Z���k�V
����
h�o-u�?|���k����:ۙ���.�X�f�&nm��5��\«�o]�>��D�5\�+0S�r�Y�$z�q�nn�xA������k/� i�A�=�r�=���'eE�a��6ZaNFGm��ι�R��̻*�����/n�.k�۪�����ǻNѦ�}��{�=h��h������a�q�2$q�8�]�Ƃ�˺	ך�}�v������]1&��v�lR���� �[D�R;��F5ǩ�����<S�mdd�o �\���p����A��_^]?����1���N����<�_A砕�B��k�o����FC�W��,�2Wl�{�š�z�"�CW��(��/sP%U�KcP�R=���A���(�p��l+`c�׹uM�{=~ð��+�lr��h>S�����T"�	���&UiP��}4��V3ݨ��ͬ"��ޚiᏕ�3�*-�k��Ny�W�l ���D��8��xMr�C3�+�DY��g�^�FS�.QV3#g1�s�:y��C�hN�|�	>_�\�D��P�fd��F���>ވ5�OȽ��c@i0ny��s	����f�	�׈���^���������X��FH9&w���9T��==kغ��r�d��<�m��L��rA{��~Dʞ�n���5��$YS��9E�气4�LdsZqL]�,�/�����%����2sA��o�<�Muwf�o[ٻp�;s#�6.�R����tׇ,���k��S��f6+�ړ�k�M=>��[ڕҏT�wz��;YңQ�m�T<Jj@Nk�($3�%R �gtt��f�R̬�����7������a����j:��>s��'��zB�u� ���
��=1���M�Ú��P��̽��K6BR;���7��";r2�71��(g�ױ���\�Dk��8u��Ķ*��L�GO����+^�1��kf_.�/v���V˽0�^3 �d���6o��#|y_����I�f�5��Ͳ�*�Su� �gf��]�a��
c9�ʟN=�j���;t����:���[�kq��uKP���CL~;�q��'��zC�M���~c��;�u������]a��4��qJ�˘�NzV��z¸p�M�'�|b�=�SU�r��w��잚k>�c��6"�����;'Uq�'0'�����Z��/���x��Uj�c6�1y}D��~.9,���]�.nu�U��XP�����k�r��~T]&~�
v�00¸��&=��m���j!�9�yO,>Y�<��t�Pu�O�Z
wдz��5��j����*�?�%�mEx��TL�U��{[�{��bt?2�K�Fq�.�ǯ[ռ�-ِo&V"X\� �\ڔTS�2s6)�5�e���� 9�b�4ꂹg[֋���f�9[3(�ܵ��'H���Ъ��	���2�^l+e�!��X%��A���Le�^�7+^J���o\����7W�,Q�h���Gsn&�#W�����q�b\��/w�s4w߯8w��ɜ&!��
(��˺�h�"�v��t���N�j��Ƚ�!;�M�fJL�У�����=�ăڙ�$�E��k�<���f�0Bq�3��$�^E�,��1��%"�ׁF�[X�9�38�;b��SZ_�i��[v*�d���L���yz���ta��9��Y����q>�I> b~n�H����9K�fe��I;˱:� @��9�a�6ད%�L4�ܲN��~Q��r��*��ە�������/�����Av���H�iG�!bkקzk|��eP����8[�*��h��L� H��z�Q������ѱl��ls�&㞙��`�B:�[���ù�ܣj��Ҕ�P����¹�������x�>H�yzKW=9�\����6-Rj{�-j�P���1���]>�gYz�������#��?r}h��v�S��8e"3<��%�rz�_;:F�BN92��u�&o���}d�)��hô�NM��R�� ���#��&K�͠��3�С�$�Wv�?� �^�����15b�i��%�VVm��t�W9��QkB�F78��m��KF�i�qp�8r�o[��;�^tf3r˩�5�q�|@*�S�,�u�o�n��o������AK3�.e�٢����9��y͋v�8�n�#�m'\�n���/�;6���N﷙�l��y$�}@��-M�\�y�����N��E�������Ԯ�TUaP���USaU�3vt7�<�<���|�LG�=�ǭ�D�ڔ���p��#fl�Q��;2�n�Ӽ����ߘr�&�=<��]���	��%=�<�g�c:1��sV�5�aI{	�Ƣ&��fHOwiGRc��	 F��5U�p�+-�t/�њ�ލ���=�fӃ�R�]��Fa+/s{΀�%٘�ٶ���Z�5�����v\�^㙎�Kr�m�`�G�7Cs��a�r�*�4��o��y�L����7BNB��w�t�wuZ�f��퍜iwiY�ڵs�'�/��gX�#��REa]�������	 i���r��8a�A��Wi�����*+�L*Ғw��*�X��Z"�W��i��6����y���2�Nd�y)�|��Z���d�o+���ڬ�y8������v{�
є�������nY���G*;}���+��m����_C���$%�^Z�7W|)0���G~�P*��)��d�øU�y&Phu���O�6���N�t��6�]<{С�+'s�]����J�f�He�t��`���7�2����Gѳ��!��AF~��P=�_H�j�W��;Ig�˙���g�鄗��.us6.�RVS��.>U�	ePc;�|'SN<d�lLX[�H��wN�`t(�Y������3XN���7�+p�������U`�:��Vf7u����{| �8P@�[��SZ2��I�	��A�%l�����3�m*�Vژ�+��	3i��$���������u�H�i�fe��s͂	��I�V�bh�Ɣ�G-�G8�s�c����,��L�y}b9X6������g��Pe�k���1.;��k�����pL�f���7܌��/I�t��b}O�l�wNP��s}���%+���d��۸��w����G��V�u����z+N�Ɔq�Ζ���Vವ@F�fE�ʎ�Øg�ڊ���a���y�1��
����{$z�ʍ��r�S}��|���B�]�U�G���Y���qi���ӛ��!��̻�6+��]�"��N7�2l_kr&
/1ͣ��љ�a�[�1]t�O8�1�����'H�Y���Y{���e7�Ġ��5B��5�t�]���`̴ڛ�-d]߁L"^�;:����X�"����6]���v�&ǒr=��&�l�ly���vs����G-�N�Y���-0h̰��\��11��n�7:�t���)���d4B5t]$F�￝���Ǡ9!O�Jh
i�
ukDK� fs����~>>>>>?�������>��ݩ)�j�(J�r�A�)F�Ol緧��<|||~?_�ߡ}�S�!�0ABk�@�M!AI�&��(A��ą	�(
6CI��5�6˥)JJhz�B�n����들��B���w=F1��#�O��	TR⤠��4�AEWX�4��B�4���ua��'rwEtZ(
�R�I!��5�4h+�:���ҍ4�U��i)Mi��uORm��r�TI&̑��J�G���Dά&��;�&.=�εZB]WO�*�$Zj�P~#��kzՓۢ�by����G�T�9ps���X���H��Ī,BB���e��W�D��twu�?��l�h�C����|�ߛָ����Ӟ OU��P%�,u���AU����U�B~������A�6��6�^��}B]*�	��*����t�;/wH���;����6�hl�g	@K�!���<�^{Z�|�
N�ů�;Z��=Ό��qG ��*�BU�A�FͲ��-�?4�а`E�I�R|r{GI*c��q]-���m����f?�SnR��~ka�j���c9~�shll|:�E�Z�ï���Y��(x�ig5�!s��2C.r��̍�B��TXSP=���#cR�8͓t�cc�)�[��3�~o'0+&v�{#���M���~�뽉E��!,��z��WDp�՚��Z���a'"�:�q�C�@.�q C��ke��O�zD�wJ��4i�R!vb]�޳k�~]?}S��OOh���@'���@���>�I���C��E�	e�ؑ�YDe��#�[�n�P����QL���<Ӌ�|6��s�K>��l��b�.u"OwPGXV���p�˭�Vٚ�2'�0���\�֪r������O�J��
�1B�������TL/c��=����4ֻ�-� h�����Z�˳�v���&�%���o)�Rf��A���ݟʰ�܏�%��l�z���r^K���ݱ�����|n�s��}�7��цB[�Q�	���
�{'�\xu���ج�ܓ���_��{��d����`�s����K�sSƁ�2q��*�
���eT�/m� sӇk^]��٦ML��y�X�����L �a��v&2�^��9��(q�Z�T��_���G�\��Ԣr���p}��R�~��@0�~&xs�-�@�=u��~d�7����\u^���hh���뉵#��	�b�����s�C0���phR�]�'��G`T{s�f_[�����%�H���l�^J�*��{C�������I��y�<�7����fJ�4�%�ak�Ǭ���^���o�">�v\̓�
��<����D�Z�����[��m�/���+�+�o��N���^lk^9!��:U]>j{�L�=3r��ڧ��m�(�����?;���YC�R�?��G�j�w����.rzm�Y@�Rq���H��p���%fӹ��~�o6��>}����;�{���d|�!�s���^�K	�"Sm�,S���wz�7�ak��w����}޿�*�V���YE�yـ|�7���{�^T�F�)�dY�zy�����+��n������}�>�H�6\��I��h�:zp�k-���G�-��Ε��gju�zq�PY����3��|�_A[,q\��{�|+�ıU�s�yJ8�^z!�^Lk�<Y.%yƺt!n�k���ݺo����D�����{��k0uc�w��p4�I��6
��5zT.�#'1�^��ϩ����tC�8I޸9"'8�&�cN�]wp5�!��Q�p/Ƚ�tS�F�
s�@�7��41�M��_E3���c�>�w��հ��B�7H8H��P�n��E�x�5�]C��r����8Dfร�-Z����ֲ6� ��%ۡ�6���J �&ʞ���-?5��4I��m��mm��"��w�m���5H,��!��-8`|���}Bl�9���(]��7��ը�0��_K���� Ou����{�E�9퐙58{���@G?��ڹ�s�B�����/��g�t;�թV�#Fwo�At�/c�a����5�f�A_��1�{�O�jM���n�א�%�Yc�,�p��ҋ�;@�(��c��q���4��f���c`3h�C���#lC8��렳$��6w'�>�#��{ˬ���ۮ�_�����JI��wʮ|IW/�[J���,$4Ӆf����Vm������$=ţ<Ƹ�v��O��;n�yo',9���`�}�NT���|�8��%�	C���ّ�GG���]u��Z7�_{���o7p:V;a2�ጉ������ɿ����5�����U@�����_%�ofH&v���:���^̄s�ѓj�.��e��ϺS4�&"��_�?���������ܖ�92�+�DB��~�3�^?|�EV�ٳ��_Q3z��pK(!<�[���S'~=����g*wձ|增�<��r��P�ӜS��{l��n��T���Q|��������T�)���P|ش��l�^��!��!�����-�;�WR\�L�un���/!��m��A�U����N0��ǯE��M��|��3�6�xapV�b9i]������Y3����'9D�/`��XThUyF��W=���{wh�������6�^���E�d��'f��gעAd�~���L�و��ґLh�J�����+�Zz�ʵ�.{hY�~���_Ǡ>^�e�����t3��a�t�I��a	����?.���zL�R�k�����d7b��X�-VEp�?�/�ڏ��/`�U��f}}�=�Qv�mV��3�Sgm4_v���恬����vi�g�v��a(�t9�i��ڨV��ս�!𯼃b�}�;�Nݹ؆ ��x�ސ����Gs�|w�D��eC�l�_r����p��*���ຟũ�6�&c)p����:�m����A��]�������q�PZ�[�u���ɇ
��	?w۞۝����e��ve�0�fs�/*�Ê��q�ۗ|ss���gX��jvГ��֎mm9�j1ɞ+:؈盥ˤ�'�2�N��G}��_P��\����,��e�td���~gA/�L�bJ��TJ`�Zخy530-l[�4v�!����C��é����`ݺ�m~/^�����j��K�1���O��k`/�3��}�a�)g�Z��c-������0d(8g�L��9���~��}	8�t�
$@�b��P���,+*f�� ��]�G�Vje1�~(�a�����0�*�^s�С�$�4�qE�bb�mm�vVQ��5�s�� �z�u�]B�te���'��*j���y����α�rF<u�n��JF{����h���[��������2�[{�e1ׯmQۭ9�SShwN���k���!d$W� ��
�!����^Ͳ�Ο9��=`�����P!�|�'.lbB_�+�v��x�(dż�%��GM&�8�I�Q.k��T�^�]�����m5�T3f��;-�e��+�H�0\�K��G]�ч����TA�؛"��i��Q�nDW����=��%��%2��& ������5o���8�4B�/.��XÎ�Ϧ�3����:��FR�c��T*�v��Ts]]W��W9�I��6v�1�V����L���ނzq+��9�*g7�(��MB �[uG��t�*�.��m�Rzr {љ/G�li�W���_�՟E�&x㝞�No���jF幟vdH�I�!@� V�X�Y��n+�d͗ǉ�ݷӚ�x��IJx�lm�����@��K�AsU\8w6<Mb�f�W���g 9s�M��R�޺3��d����Jl�5��� P��vzbz�g�HQ�]��Y*���(�]�w�J�}���d���l�ǔݱ���b}Z],U�Dq�g�w�r��`��o7��U����Nf֍:2�`D&�G�w�u�R��ڰ�m��U��Q<ݹ�g��c�Z:�*{�6*�q4�|�?�����@��U������K`m�+k�0h���ע	�KOb�@�c!�<��Fa�o(@K���|�"[���g��w6��P*K�A ̀LG�t�3�΁Ƌ9m��<��s-����~�{��>��\XjA��Gl ���7̼gi�5��njsﴢaޛ�wص��ŕ���2<��8��^���t�:��JZ��w3�y��c�[�PF�b͍���ƶ�ࡏ�N����6%�N�#���0('V|��f�{UJ����H�gm�vHl]���9�枮�|��U�v?C��y�����#�:����SNo�6����z�\vQ�7���FZE�����:
ڼ<^�4��uPϣr�{�����ص�#�l^{�d\��)�:���{j����͌b+m\K���"��0�>[�d=��!al�E
�y���=��9:&�yEO������ߪ��ȼg��r�v���eO����ZJ{��_�Qx'�H�EU>]첿M3�뀑E��n�(�dUdb�K���X"����J����-��Ǌ�?W�W��']e��;Z|o��qv�
�����X|���i����ϯ277h<)����v�Q�,�5B�P+��dƭ��Z'�QZ󦎫(�hk+���.��05MS��u^8��Tߤ2m�0��;��q��r�3��go�݁�U�F�c���yoS��
��ח��=k����7���zDF)��9֭1]�;s�DѦ���YX�J��YI��ݬ��ӯX�~շ��D&V�*t[p�/F_,���w\]x;a�)�v�����9|�o�\G^�1E%�(�2:��Ġ��z=������c��ٷ�h(�lDywgDm7U�o�y�����5�˷=�'�#��≨�T�A�"�>�����`8�Z��%:���綫`��ɳ�ݲ��{J��z<Ў���~���c16Y4~yׇ�w^s<��1��g�/~�W�H�-�ю�4P��Y�ك7�dL�_;�U��P��&��j3��c5�;=�vJ"}Ŏ�l�,�nz���4�]T��c�A���sqK�Uɾ�����Z��ۗ6Ty���ɝ�˰��j�e=�S�>���� ���H�OOP�*��`��g�x9��������48ӛjn�F�8�n,#���i^秗��e߱W\th����>3
JAm{�
iG���d��Ȭ� �r�ø�Vz:�o�D��֥`=��n�o)D����Aʹ�n�{rl��gR�bp<]�M���7�_�^�غu�5�x$�^����9�`\�KT
�R"V�hE��Vx��^t䍜gܤ��q>�>7C��V՘m�X�C�a�%#���F:Wl�L�yb����Nwt�\���P�H����ۂ�s�7������9�%�Ls��[x�P���g(zXG�����7z�範B���H��������[G���;SÅiD_E�L�R�0��E!F��:�ΐ���՞���).e�w��s�5�I������ū�xٖ�x�t�^0k������rgy�'1�k=�Ǹ���j3o_��b~�h��'�(�so�PQ�oLB��dB����*�l6owF�vf�ך)�(�u�;�k��6.�͔��7<6mL^oKmJ��p�\b&�5Vx�EN�HR��JVH�f�a^3�f޳����giy|�c��%���e��n+*�z�����Tg`�8r��1؇qw���3k�����0�07k��XM@[~�ν��y�ʢGeʅ,Т��5��g<�*��ʳ��:Ǝ^x����B�~I���w��-?�ؖ�[��(F�FH=ͪp�A�G����p����xJC�#����^/b����9���K�^���x��%��e�=9�5���!
,Gk���� ��/��q��M�\���3�]9��n!E��<�Ą8�y�L_dZf�^3�Xkd�l�Úɷ�7;�yK��f�w�O�t��Kr�9�,�����{.�.��LV���gvYdZ�H��l�;�d��뎳���m�4��t��Pt�������~��/|��!�N-]��pxwN�
�ᕔ�j�t2���!R��ʌ���纴r���<YW[�䶼;3EI��cH=a��e;.��j�q-��Nz��6�����ǅ�0��ѻ���B�H�d�b�t���I�N�?ݚ�OH$�ɃI��]�А���<�%�z�*���p{�Υ��9�T-L��<*�V@�n�0B����'�}��:�v���׻�wFi,��ߪ�2�=-T�^���x;/�ߋ�gkw,��}���\{:0�\b9��$J���=t$������ЅͰ���0C*���Y}W�3r�z���j���zDY��=W�Uz��='�����PĜ���y�U-z����[�B ��͞��ܹU���M��<�mx��z�j�:h�k��^ՙv���8�D{{�A�ޑ��@^K�jÚ�~��}\���|���g��Ή݊2��z��R�t��|�>i���H�[h����Y�:��:��"���Hm�ʠ]S0�w��;5�[2:Mp�3&!+�Q]��'y b# �V�#�NٯjjȆ539����8�(�&n�5�Y]��;��L w�oh���x�2:B��I;ڠ���(]`˫僐<Qn��;�1;J�"���,���Ϡ�me�վ[0v�&��E���wb9y��"7���޾��<����ul��z>r�*e}��f��q|��,�EV�4�R��:���8	��SE��,q���YY�O�_I8֠�)��t�Ȝ��=�Fq*�U�KM�z7#�VvY��fQ;�l����H���j'�8P��t�`94uɃe���%I�t��+��c���s��G���F]]��N1���U�`�UXK�0A>�.։%	��C�.���5�v)���g�
�b�r3��bfv"oY*8Q԰�����f�	J��n|�}\g=��&���ֱnM\r��kr��DS᠞mu��P���R=��W:�����<λ�l7� �jNw�c׫UX�e�
Amb�q\�0����:;3��f��`b��Wb��Z5�����}�A3Y��3����au�V%z���B�1gfBs(�㖃�o�PQLCzoY۩J�]%�Kʍ�
�����G5S���x�܁�7�:��<`q%�o�*lI���6����7^��
�F�˫��5�$�;%�$�.�b��3��D��}W*��zi�X
//ӯ)�b�ۏ�B)ؾ�b%3����M���}1����gS���|�YI���4��1�[Xw���ܧ�2�v>}o2�X�c���k�X\�w;�xO.8����WhL�K&ޚl7����ǘ�v�ŝ.�aꒀ�pLUl]=Åb�oZc�h�z�E㽗�_X���EJSP�c˰�b���D���p7yW����"._�J��l�V��J!ɛ&��f!��XUm��~���v��=*����O��&KY�v�qT���r�m9Δk���;ٶ$�vP�W� �(�3w�XT�XN�7�&���ٷ�&�O-Q����k��E[;v�&
�<a���\ٸ*�}{z5'�֩(�v��[ݓ��CL굝|�CY����hk@�+���u������~�U�C�w��m@p*;�LlV�q��r�C��J����;G��v�H%\�P̂��-����&�L�"�/����j��E�0<��0N҇Z;׏����cW[8*���:K�M�x4�A8F�r)L<yvvk��B���;�˹(k0e���R#w�C.Ҁ��p����=��_\{%�c_;8�M���1S�^Z�(S7�3~�i�4Iqof�$N�Msu��+;��Y���-�f�[R�\��]'}O��&�V۝��o)| �G�0W�v���p]`u��BkEUTP�����o���������x����x���@o�:�#l�f�:�WF62���������Ǐ������������J���!�Mu8�E�`�TkN�&�l����CKU�q:�A�h4�
j�JX�����s��``�Ո��۩z��;����u:(�vz�)�V����&i����&6#�1D4E�
�"$(�b�֗gD���U������Кb=cPWs���&�
(�-�D�4S$���IT�4=lTD�]{���C�
:�""���uE	�k1U#������=F(�$�	5��;��5����U�̬������c�'|wE��.�m.l6_KyU �V�:�n��ǩ�x�S��,G�e�`x
����O�{�{�1��}'~�i����G4!��8U}��zq�t�#'蠗L/I6z���=}��-���͆0C�1猾x��ɶn��Ͷ�ݺ���n5��\c��:�1�Wi�<��=Z�⯮q�0������\�6*Z�U�����m�<xr�"G�	և��M�p���;T雦f�
*�R�Dm]u�ݏ^""k��F��i�׿Q�Z���eF/s3�\S���2���P(���z&:k"�j+��	A��VfMvJ������>��"旡�k�����c���q.1��-�E�,�s�`����{i%q�ZR��%vH=w.�ul�pMϜ��e硚U��&W:*��j!go	�)�ׇ�zUO��A����c�Y��sں�s�W~8�_�~臣wB����+yHҒ��h-������7K���]�nsdJ���R�2���fD���v��1���"�3��$��S�!����ܬ�_bA���OVu�,:��L�馆�-2��A���+	G�]��$rG�3��	%�[jh�^M�'TE˙؝�C��哝�Q5Ӿ^o0���<Ĉ0qyŌ��oT�0+��/y��_�R*�<���j�C=��O/5C��x�PY6@j�G��>��v}����t�x����z���k�fbα�Qm����z]��>�0�������؂�I=�et�����ڥٯ�#�-އ#�u�� ]>4���LÏ��\���АA�^�����+u9xy��.� �Z�S�LŉD�e���2�q�U,�[��S:��Kّ6�U��?#��VW-��O/H]b��Xˬ������1g�;J�2	g�����/�g?ރ�А>���c�y��nS_�R{���6�c�v|��r��f�ZS����^�D��D�Ţb�����]�_j�fu�X��S��C?�w"��U�I������[q�-N�ݾ�p~��T�vh�Kw�����'��] ���˚���_�?�Y�Z�yR���a�;^q"D"�fGX�1n�8���ffv����J�\Q��7��ST{Cl���:���s������9
�aw;8��N��N�΃���E�����\�%&:�{Wb�m[�sxL�`H~��}uT��ӿ9>��;f���In�	6F�F�8���S�[5l���E6�t��Y�t/��9�m�c�]9�W'ӴB��$�J:I�T{2ni̊�O���G?B�������D`��#4@]�|.� {ˁUF�JU1�i9W�e��;lVvd�ʓ��(����U��b�d�Y������Ъ�#l�}V�0?iݹ��Q�O�5?��HC�Q85ns��ۨ���̊��f�(���z��9#{WQ6g��ۢ�50m�B�E�K�swO ��z~��<�2[���*�6�l�vtRpKa��ko��~#�`��V�&��������^�9d��y�F(ܻ |�����[B��P���MK�/_��<4P�$3��5�dF��~�x��z(�G�[��a2U�����7��&N��|�|��6#n����ǁ�{˺�Ύ�x���&�>N)��6'��t�!vqrQ�]��e��"�u}P�O�-}��.6M���o�ŎS�s�H*f�~���Z�[e*#��z��qi+=O��Y����U:�������ɓ}���q䓏7���(��u�iL��t�B��_߾��}'b��3=u� �����^�y�Q�@Yg&�%�LΡQ��B��M7X���o��I�nh2��ϣ�����WP��$�����V�x�x*�nc4��;�6���[T����:$��ca���;Jz�N-U�6Fm]����5ە�}گ�_7�	H�N�r�T:-Ί�a��n2ꇹ�����d`�M���5(^�{����#��<E��$D�z��6�uwZl�gi���K'z��P�va�^x�T"mu���gYh�4�cN�v�c�%�6uۦ�V���g��c_57�!C�B�F�Jt�׈W|�M]��z�r�Dn��yrw�,�8��fo��V�m@��Ps�	�#�kZ�+y���(_Oe�Sf��y��u$���T�ʏB��R.�B܅8�E�)s�����mU�C�.�q$Ŏ�V��\F��T�s FTs�GL(V�b�/���i�r�JH��^ �nÇۂ�->η�5T�{wD��ԥGZ��/��5z�"�ر���yD��V�=E������{ڃ�u��wN�޷R�e� �#\pv=�p����gkdRf:Ķgd;Ըm��y�tWqn1P{\���+���J���FF.m�vzCx���s9'e�"n#q����T�y4OW��U+�����yԊ�:D��`�d:Xŵ�a�nC���W�R�L��]P�]!5���ݷ
s<j�;�.�z�L':�0�2�9�k�+��ؤ�J��kv�pƙ����ROq�|�:�a~��vRUǤm���7ͣ��އ�
��i���դQ���+�&�4˦�j����Պ��2"A	�`GwJw-Q9�ёF�7oN���} �z��2׉z��$�LG�t�6�{�/LU�s���d��/�� ����֬��C5�=yo��0"H�<�pUW�ݙ��+���O��^Ei��D`Cz�����63�/5�Q�9����&8ɣ��b�^gBd+l�1O�g���	C��x~����V�_�v|�i�WV�����6.+m�����:���bA�^�w{�x��q�+��{q�{��v�Ś���r`F���2S�CP�x�V��]tvε1ނ:���輗�P�Y%�>F�^ɋO�(��I��Y]����q��~o��p�p���&�����#-O�i̍�|B�#n`���E�2��ɷ�w��m�m:/����Y⒴�t.��S�*���_ߖu9�ֻ�Z��鈿ɀ����s �{T. �J�M�K��f��黏z�;�"Z��Ng��?}'��[��!���JJ��#��x���{_!��-7�/3GM�=�luC��+�5p]E�6y+�"�s��,��q^�L�^�}��o���>	����H�[7�&���{�R*�w�(�2��,w���Ө �����˗�w���<ۂC��Ǟ��"�k���ߥ�i��x�'�v�s�,��y������i��5�<��0�8[�13���P��ZM�d���Ȣ��{x���-QR��	k����#��>3�5��fe�>�E�m*�˽���e��<�	�=B:Cj��e�����Cf��ڷ�ز,)�:8��"�iꥰ{�muX\��	ў�5����������S
w%r��lV�
!���w<��{��3�=��'t۝?T���x0���&8�Yy�3����j�l��G�o-)HY��n�洌�Y4M��}_P�"�ۏ�8�e�!����V�����1����f����w8m��Rì��(�V�lk�k�ڪ�st;��
�����C0��Vn1)��d��7�+�6�pD��ܣ�V�7�OkU�1���>������WC�I��ֵvfR��ǋ�z��{{";���BG"�WJF�9��X�APT�����0L5�-�r��ۓL廜W��o`��5{��H�H�Nm��e�g�v��;��7<,S�lx4��=)��>�7�܂��䂟
Q��#�u�3U&���K�w�I�&�H��@�";�H�[>�@�P�x�*����g-�3fn�i��l�V꭮��9��T�^���k�k��I�pK�<�e�z���L��#�̷���@?\uө_�ǝ!��h�������Uj���P����l� 6Ǥ�Y^&̆�x�k���.�ѧ���#>��~�m,���r�Q�Q��=+~I߮���)�է{���5�z^����A$S��Mq8*��j�䜥��"[���6JokQ��+�F��&�����p��wԘ�_`�HJ��8v��Z.㊯�r�a�����̃Y\&0��F���}@'�0r�Xq�J)J�[3�u�|�T�7@ah-`a�����39nD�"z��g���d
�E#Wt�.ǀ]�m�z�����Z���������"K�8o�f5W7uW�7��K��J�'����u�3��r����l��#���$
�
̈ۊ�J���1Օ�]�i����������כ�Y� ��7�7�.����Y���a���	��O�{�� 9�J8��O��5v3.�&v|�~I&z���@�F�u�v[;�;Ϋ^�^��eZ3�y��fz���0_/�8�D&�_��g�=��y�?�⽽�j���@~~��w�Ay�V�?[���/}yT�9����=���^���u h� �"R���O�u��a�O�pM�r�[]�l��,����\��_����_�<zq+����?�N��#��F���b���U�Zk����&ۋ	���te@�����.�iQ�r�<W5Ig4��v1oh�BI�A����z��f388e����0ۼ�.��X��;��el�]74��+�Z�UO"��e�����T������^��'�ͬ�̫n*%�X+�aߖX�9�̍�t�r��df�,:��v��4��y>�gj;UP=��j&��	) ��h@���]�l13٦�7G^�i�yZxJ�I1�8�jF废vdH�$.��,��mVGoF�	]�8�"��lq<�7�A����[ge�����f^h��ì"eSn�5N�X���.��I�v���4-�5џ\�'g���˚�g�ɵ���k:�~��]|k�f%VW<��.J���U��������Z�a��g�C0�m[�"
��f�]W��+���{��w�����wr*6yiaq�@��`�g@a�G��دL�n��}{�0ԫ���^��zi� �&���g���j^�G4;���چ�nJ�e٧��ێ�VF歡��L�oS�wl�l�s�����M/����x�o�.�_^�ק��y��F��*�VO��5|�F�5/j>�X���<�ѹW�h�`�:gw+��=μ�w
moz��8�F��9���h�:k4Y>�����n���\���P[*)*��6潜�F�Xؽ[4�m�XS��:w�}_W����'^,lYg�*myh��&I䘎�\}^��o9e=�s�=��;���E�獤�kf��[���D��<؞'��Zͩ��S�5|�O���z{�L�#�<E���ѵu��݁xH��q���Y��m1m����}ɕ���pQ~�Ï˽���wGGr	[��x~�Yc8JuO�M=��&�:��W/�Tq.���SsNge��S���t��\��qfl�]�=}Ă���"-)U�|v�ji�ճ��I2�v>�7s��w�9݄/��01������Kڡ�%'����F�&z6�4��OXcƵ�!���sa�ල>3\;�`�5>Ғ,��)��=��Rת�������k1�"�?x�>�ȱ6�[�x�
^xā�<�)E>ر�67VU�Fl����W��6E��jtq��cV��I�)�{��w<��}��Ɯ��L�L_v����	T�u�TÛg�&9Pض�frMspt�,���5]�PeF�N5z{��,>����p��m�	 aT�������Jc�,g%����48������Э��dD�zv�M��d��D���]��êI���t��h��7H�Ӆ�;T42�g̀3\PA�/g��qO�n���*�g'g"�#��{��M��fVmҢ[z��`��MP��k�x{y�X�.0Ntp���$d<�W�f��[�p���У���E�V�8�<���z��3�Z�d+$��*�K�j�v+�_S��o��cԶ;uof�29���绯���$�Y��G9�\��zf���h%��Ҳ6v�U��7���ĸL� �b���$��-CL�gl��P����Ɣ�Ui�м�.�����mР؛�)��'��9ff�ZY�1>[�!��&^z�h�t۹��)#�|��5s�R�t�on�3�� ������6�-��4��}*���T�Ô�+�,�ZHf�{�WPw��Ե�;!9f�A�w��U�;�m[�T�q�:R�[U.�IK�Q,�%��P��r��V���"��#��vNCF^'	8�[\L\�;�o�L�/�R��	}�O��f��Nfᇕ���r���ʙ��WY�����Y�4�):e��Z<�/T�#h���	�D�xj�(nA�+��GC[�U�����*f���������M����|�Y;7!��f	��޴8��]힪7�N���`�gԪ�|�|�\Uui�S�I��%��Ԥҩ�Ev��+l���[ۘ��Y1��;t d�gh�g��;�.�v���+�ƈ�]j�ۑ���2�9�!)f��l��;��C:%�=mk��sW�����w�����Ε|Vռ��Mk���o��n��8/�P�a��xB����O�(\U4(���<�iT����T��l�w���s6��Tn�>C�a��`��ж��4%RFL��{�ae,�{X�f�V/E9�cWrjm��1�Nc�VX�ˌ'����,۹���n"���xۯ�(n�=dW��^N	�����R&t�e;Ѝ�U���Żӊ��>��n/]W\v����U�*n�,���4S����G�ݮ�	ݛ�m�n�6�5�O+2hE�WH��M;�.N/����7:��=x/<r�Oj��qx	Ӵ-ԑ����CB�FL�XRT̠������\8��.��k��z÷}Թ�^1�5jț��>�QȲ���n�x�-�*5�]�)7��ӯs�ۍSU��2��Xiݍn�[�m4�52��)�w+�kz<��{ΛAfԚ2���L�E��8�Ɔ螢�RG����/uz�T�`P�h��;�)��zRw�@���e3�-����>�ӵ6�6����X�ቃH�#�nk`�N���f.ሻ����@E߉D J:�I�ph�h��"������E3�=��O�����~?���៿h��T��CMP�ADE-[j�j�F���h��z~����������~>߯Ǐ���
(>Ͱ�EUDEBRk1TM6Ɗ���F�z��1���h��=Qh����u��vY(���Uli�H����h'l��R�T��i�Q4�TEAA1TV�SQI�b ���Z�������&��qS�5z�.�E�O�j"
h(�1m���"("=m�hh4�tj�Ƴ�:���vs4TQ���h�F&�n��LU��cEE�l�Z�$*"�������f��ت��ET�՝��i$iKL�!")M�JQ̭$��q����Ase�����n��LgM�׊.��nR��Сv�w1K5���ܡ[�O��I��gs�Y���Y)�)ف�BA�1���e�b��(�������r�c=�*�6t�����֖���]]��&W�fL���WK�F�w*)���W3y�����ٽ�R�ʤ�y���;�mt�`���oC�6V�a+Z]���v���O���=�[���K8ME	Nf/%>��3��%�{\��������e���T��[�]x�z�}�}:��
����KR(��J��B�g�\+�/z/Q�zg�m�K�Uϭh=cRƾ�7�5�W��tU�A�]�wVY՛�ZR/#�;��t���8o�w;�ꔰ���#�r:�������/]��BZRX"�L���r�2�f6����ב��.�I:�[ŠUҝ�s��,tB;Z��>���!�
ʣ�oi�� l���D�n�+��=hm�qh�
�6m*�Z6YC_4m\�x��.�hWc-��6U��l!m�H)�$��uՔQ�l~�j�C�s:��u�k0N�R�5��Zk�uH��ޒxbH h3L����D�F�_RéM������0(�UV(�ufe,���)�q�a�t����Q�ʔ����Y�u��Jwd�b4x�0_t�s۠������ԇ�s�&��¾cj��o\.{wʆJ��:�B=┦���#J�����wnܙu~�Z�I��9��"�^�;k$m����#�����=��:Uu$UP~�t�K�Z�G�S���}����i��o�YgK�5�ϛ�K�#`���&̆�}��B�ܲ�[�L�捫��4�=�|��T!ʗ$ֶۢvB�>.g��v�Z��v�q�+�V����?�p���ܣk���E)S�˱�h�p�-zBnBY>����]�Ĥ%�����0F��k�($S��U*~���M"��EJD���>��������f�;5S,3<���q`���VT�Ǩ1��͗Si�"Ep�*��E긊���^2`z�N�m���C�#Bȭ9a�R�a�2�:��!����n�EW��|Lt��#�1���x��
/�}]�x�R|��a�Ȧe'k������;��r��`sfCo�p�F®X��p�b�jҳFpEa��������KE}d{U8iv�u���\&e.�T���]�6l��U��2M��-����w^;�h�X�}���{f	vq�#�h������%L��:gixv�śS�:}��g��tI�}�?b�y|nR�_q���3�p_X�!�|���-�9�����iR4�_�e����w�,�f����g�(R�ϴ���C&�^^M�b#�v�U�)w�bl����xd"瓿^zNr��z���ͅ�,�S軞�W���ً��mvDc<ܚ�Е3y�*QKP�������� S���/	�Y��Yh�J���h]�ti���y��;)�X�`�$�Q0v��ٓ�O�dPPn}	�>�*[9y��]��r���%e�$��<j��ܷR:��"�kI�3;�r�DE�=�	ȩ��
��Hޤ�nE �&@b�����N{[����W�����s��c��zb8lƩU���t�CT�65ϒ��ͫ�jo,����9h�;*������d.��=C� ���(�������{f׶�A�����k;*��:#���p�b�=��>ڇzI`u;��m��m�K�f����Śڗ*WkK��u�6�ū�u!�`f.�s��7�HV������[�j��s�����3P�u�t3x�F�p�(�=�}_{;T�����;�FxֵK�,G�V���G6z��<��
m��p�ݽ	$� �u�*�=���/� #}����1[[x�WVglM�.��/��t�{�u+U�����@�;�8S�Q�!VK�3Xܠ�u
���t�]7��;�;�6�{��2y�|x��O��p;� �P��[\{-я2săs�;�<�f|��{v�?i��xT3�`�P���F�[cז�3{��`��ц\��Y�;��j��s��gz��\�d�D��*�mD�f��sM�����wDYs�C�̛݉wri���x��=�%>���Q1�^b�GR�D�9�}w���]���fB]m6���.i��RAw����|�ͼx��b�kn��4��^Ғ��p��ޯ}ي&"rׯI��?~��a��!ȴ(<Z��3f�y�uDJ�cVW�ϳ�$R��6��
���*����K��h�F��}���B*n�>ĕ��~�+`]�I��N�ZY��7��ؖ۩VT�.�FV�n�[+�Z�LL1+�ʬ��z+.�Pr ��َ#�u����<�$��޿_�}���A��>���p�|�zS4�L+�M-�.�B{H�AN�G�I� ���w�i�}QY����L�0ǲ/Y�q��&
�]oҒ����<�:��nٺ3����9�)y�ȹ}�i��<W��/���%v@3a���,��7f����Θ�!�vE���WHd�/x���p["9tޙQukH�W��^
��m��v1ٯ<h겉����>�x�g���@~�E����֣2�㙺���x}V�%�\Qy�,�N�k������"��Eu��T_���Į�8�	?F��][�mME	O�1s��k�	��X�*��c<l��G=�,3U�.gE&��]S�	�2�S�\?Tt���=�vt�����D�e�=�b��3\z��H�G��L���"�����n�����*Ol) ��b�l3�v L`%zDLY�E�7�66�w�˼{��ŝe��)�&��<�Y��w�f�F�A#�Ϭ��o�j�Yo|/zm�팳�T��Qn��
t�����D�2ڬ�I6��:����v%��;+�dPfk��4ul����b���v�����r�qcƕ��֑Qy�ҥ�by�T��~��}_5�/GY-��i�=�JcN��(��?O�C8�	�B����j�C���m��T�Tv�l��]tO�J��X��-t������ t[({����V����C��0�WDJ�^���HH�Cx�)uל��2�L�p�n��������W�h����d�F���׹ �R��v��e&���ήn�$�)��*��>M#j���\ .�n�5�*�J"y;��2���ܣ]�8`����W�[<�NjD"�G��j-���ݍ���48�����g�$�4�UA�㮝H���A�*~fry��HN}�i٫,�*�p@6��JJ����U<uq4u�n�BҐ�WI�y�[��2��bO7���];e�V����D���{%w[�Cr�ٲ%��:~��}Cs9�#�\�9�L�:�E#wr�t�_���F�N��eA�~�7wX�H ��䭩*��"�R�wζ6c=K;$��\��;i���S9�co(���5n��_;cE��D�MO��xB�4%Isb���4��W+�Ff8�˲&F��{�/���e�JODޢ��6���p����^o7�+8~i�n��
������<dDg�k����R)n�VM��h�ͱ�8Mf�v���f��pQ}���i���~����\��-Q�ւ4gv�I=ʔnx���dh���a�#^�������R��bv�Ft��x������ ��c��Gw�B;�\b���l������A�u��B\hf�����ޖ��� �hE�7�+�����	h��n��\؇��]W/M�yחѼt�4�@��Nr3��5�^Fn�
��uo(PoN����d�M]W�1b#���*���!�u�i����o��:����
�tǞ�����"l���\�����r�	��\nH���s��=lv��ג��B� �#��W��?y4E�"�nDu�v��r�ę�&���s�W��E�8Bz}"?���ρ�ۉ#�����c��ԘKC|�y}ݴ-2���Z������w����i�<��S�.!IN9醑΍{6�s=eׂ�ɰ�������pB�3p�AjUoJ�b���i��8��o���ϫqd����z6泎ud�|^�}�ȥ�bRI&[�C��mˈNfL�-.Ųf������LJѧ�4���м"��f�F�;�P�%q-����:�8K_v1x��ݹå�[�HX	�������z���^=]%P�+��BV)M��fG_6>���j�$�)��%���at\g�v%T��J�/�lN���t�馊9�{��@hP�7!�{c��~\j#T��U	�fl����V�\�h;���_��]�(b��W�$>� f�d0�ܩ�q���j����X��u �][Aɹӫ+�{�Z�����Stzu��\A~����3�n�v�𸺁7�W���SuW���ux07:� l1ֲ{��%���u�{4�~��� iP*^2���J}x��v%t2d�p���*w�%_u�^���0D��Ti[��3��Ψ؊�k٭�#ז�3{�R��%��e�~B�T�A��SJ�R}kf?�N�/��d��3����%��Z�]b�̼��2f����F|���{�����:}%J�N�@[7%���8eЪXhU
���o3H�CT�W&#�ջ��ux��|�۶���0+2k���&�?�������}� {������<6A)�Iv��z��
��U�8 �,��R#i{,��8���v�"L��:\qX��9�x?O��C�ٲF�ЂP�rj&�أ1l*3�����wAw�.���G�z��K��)g�i�쳡Y�qV�S����]�=b�:����k& g ��F}F�h؃W+n�%�Y�����sqf3��fY	�S��=�g���{��"Gb�dP��T�y<�O�t�ݗ�#�h��14�,e�lc�u��������En=j��$�mWw����W�o���H�pj��������x���Uu�phْ;;:R�o�������	� 1`6S��,��G�:'��h�3oW�Ϣ�7��y�;ݘ�R3��_�OI�y�0{�~t�P��_گ,���/q7�j]UuȔ�jDf.�W27�t=Nĸ�Ӌ�x`㱢"	�W�ߥ&_S���oX�ᵹ'�fz-}4u�cG�*j�A�D�E��Y��{F�2�\��ΣV�,��v��OT�GS�<�w�Ό��1@�w{,�	�`���yh�6yY��b�X�'(���p_ǳ9�k�S��� �2Xy�޸6�zx��>�����m���KhMEJs1}�8*�ٓU�A��:�����,(@�ŭq�9қV݊�{��p7_:L�����_}v�j���t����v?���2 +�	�pa�Q����<��v4hӶ�x�e�1���:�?��8C�0'/
����,}���5��c�,N�l=�d���H�qk24�G�y~�l��!\�G���g^so��+�j���Y�W]��W>!r-���K��O}������5.n��δy�aU�Q*U܏.HOZƑБƜ����8���u��}�p[����1,
��15�tQ5k��B�H.�� �;�=�����;2D�.�O����;5�EH�nxX]�E��d
:��L��I�w��i���Ex�Ph.9��܍V�E]���
cU�X�^� /&��.��?=vU�E� ڥ�E�F1���"#b���;Ck��*�D`ʺJ�E�Ӈ��+8��ZG�c��J�z���8��t�,�����-r��7���q�ǱH��.�(��&ʛڮ�����3��r��%���0�%m����K�Z�HwW=���ר(��u�Agf�N��˩l͖#@�Zb�E�'Ǎޚ{�z-bV�2�L�A��ҵ�\��,X�M���k�� �ո�v��-hg%íl�w�{V�׎���Oyņ�	&M�GdE�o{���`�]�\�m`�3y+A���c�d�1��������/��Ai&�/���ľ�̨y��˅i��V��e�sH�bL�k"�V��S(��t�pF�7��洂5T���D�	i[/�V��z�k�j�P�s�d9�L7u]d��vU�jwe�x��ՎE����5�`X�ʐXy�܏Z�WPr��+]���M��*���Ќ���YĒ���H?��jn�u�|/`o���#���F��
z�æx[R����e`����&mٕ��G�q���pb'{�bk�6�:"WL����y����q|���fl�V��&�iӓ�5�9��DhKضuq��G�$�@�]E���n��9e9��r�^�)U�2gq����7/�צ|�rz�"u`��u�spֵvcf�_o[�j�Za����L7�s��yh-Ĳ�M�(����PE��m\��^p�J�	}�����r�,Ks܋ٻu�g�8X�5��X-���\WD�o��b�!�*�wFJ%�dUD���Dv���T:��vL������9��$�����2��X��2����4Vö۸��@��rX��2�O�[OUݧ�|�)��÷m_-'Q�۱;��x�7-�nl�$*i�Z�]	*�.��]΢#(v9�䙥`�lM�"��k�*�-:�veqN�G$�|���Y��i��NB;\!wabzf��%\��!���Ⱥ<��^e��(尷���:�y泑aa7��D���b<���s���wKc�ѪM�f�`9o*Tv�ÝEn�B_3����Dto��8���jCh�Ӝ�߮�9�".cǄ��6ˡJ���{;T,�1�U׉�jlvk����:�;
��0.� n��xG\����v]WWZ��2,�"�ؒ�H��( Ǹ�j��Ov���|[��֜6�3c%U[6��1�Zxt�f��\��*ˈ<�xb���^�����΀����U�Ό�h+r���Gj��.ve������ ʍKs���&ċ�)X��Wۊ��UR�����=�+`����yvs���n�eA���V�1L"�eV��Bqm����^��|U��@�0�bt76k�,[�Ֆ�ӿz���ϒ�����y�A�M��4�W�%�_9�E�5k�z8Vb�]WI�}��jn3����)K��D.�$�H$�b6qD�TTT��GV*h�MUSLUQ15ALţ����������~?�������UT�P�UUTED�E5A51Mg?_�o�������~?�������W6�)��L�EEUT�DTL���������u���UERQUT��'EIUQ5�TQEGV��B�
�&ch�"�g5l��*�*���TL�SDQ������i��(("b�A�*�"�&��CS@MD�SQ@UkIF�DLUS3C�-I4��ADQ4�DCP^�4���"������cV�
�cT4�8�Q�UEQ�*&��[UD��[U�e�!��0]�h��w��D�TETQMT�MS�%��ZJ ���d�EAE5E1B�[9�]����V�|��J��
�aoD3ک��N>9��2��(�Wp��Q���e��uZ�g�m�5�W2N=���z�O_K�o7��|�E���4*�?\�u#Lt��S;�p�މ�a�;�,]�������88���󤍺�iK�⫰O3 s����G�@چ��+`϶��i*+ܩr���-kd��Sƌ���e�u:��8N�5��%�qC��j����ޞ��)�Y\��Z�o�I��q������N�ڡTO�5�v@u�ǈΏ0�e��ƚ���ܒ����י�,��L�۹�A��L3�F?��0m��FD7[���Z�>�WO���7�=ڈ�^�WuP3��2|6�lo���C�#Uu�$��F�we�����d������Mנ��=��h5X�g9�>Q{:��Qb��ffaq��Z@�XU���=f��:E�i�y���u�l{�ބ�+�xI��ki��!F�jk��m��;=8��;Ǆ�F�h0ԙ3���h%2C�ً�ܴn���ǵ�U��^�C'�m�&Pg�S�V3��,���µ�ҭ|'m�X���lt���:�Q.�:�!GUX0bq�j�࿫������և��/���n�3*in�tބl.�؁�D�߾���O��x�g7�_>/Pk�>�Љ������GP�L�ek� �^�׾��<��[�+<:Y��\P	C�O<O���f2_�8��EKm��գ|ٷ9�l{jW���Z�4�i=p*%���sN�+�����v��Y�3*�lrJqJtW$dld�o*=u�/��[@@�ݶ���3��b�<��'����̀o����:��	$�9�}w��Q�q����������?l��qz��q�E�pQZ8G�z3a#c�"�Aҏ�Ks���ᩯ6�t΂;*u:�@��+�AZa`�- m� ����������<���9�{��\� ����d�	�����0M�;Y�ޣ���Ow�f4��g��p��;���L�gv��v��q��D�8]\�{Z��H���7�[7���˪�T-w�[��z�Y��k��*<���/�:�ʩ*���kǍ,GؑQ��z��y),��x�Q}�������,��v݌N��,��_5���X����Cy�_;fc㗊�:t�I�� �@�>��N�|s[�����8��s.f�d����\�M�V	��_��gm�sʧu�]�y-��K�U>���]�HWkBm�"�M���O9����݁���q��Q�W�7���{��X�dk�m�z��]S�23c�@q�}��9��7CTd���4t�]iRlsđճì4H��� #�� %mq�Md�lr;
�����18�NM���wU�a�諟r�]P�/��<*5h�km�ˉ;c�SU�W�l���0�]��E��X�h8* ח��g�,�%b6���2��%妧��T�{����2ï9��-D`�ɤ^Z�tS��;��������DF}u�h��5�Ws�'�
�~�Kl�E+2�[^]���3�-��ڳA�_�_���Oh��P�2|�/�l��
֢�ZR�B�v�H��#fC]̙쪶/}�B1�{a���6�Eۢ#˰��]#�>���[�sLum��6D
��I�θ�.���5l�� �ǔ�W+x�BG�Y󚗇�n�v�a[�t�.�WZ ��g]�˩0���9��j����^����2a�{�`���\�Z�̈Gx`d3up�Z&D.L�W���}��r����^��f�[faw��s9�o���r����q4���`����;��>�}_W��k�l���o�o�g�a�Ϸ��U�[~p^�Ί���k�.͋зf�>�[���Ӛ��>��t[�;��1m!�-6V����Դтɽ��6�Oo�ry_�ohW>�Z��#Qn�f��oW^?6�I�b�)�'-��i�:��:�f3as�,�8�E,�N����4��I��:�e�L#X��H��s���w�q��݊��������#�׋��Te�v���'�ֺ ]'R��9����u�+��جX;u6{;+���b��@�P����g9�`>٘
�Յ�en��̵�5h�:7�����)��wF�#�ٺz�8�g#� �|�DY�s�"&/�=�}9��Ε���o����XƝn�&��<{�ש�|���ř^�F���gV)�Wj��7�RcsI�Co"�yJF�T�_���1;T캻8	٠W�7NfȤlkE���k�A*�ty3�SԉsXj�Ds��d��ߦR}vV�j�.B�բ17u4�j�*0�ls6��n�D�YGV��EVgCE�pS�;�*�z5��b޷�����߻*���ivϾ�y�YY��7-��TX�3��z/r$'�hl�=�OA#��ӚY���W2h�>ϑ'�����~`ѯ�W}m��=���8�$h�������4{m��oF4����4�@��x<#˵M��X��z��/��g+���4-��Fw��)W�|v�}��M[8������i�C��.�9g7��
��p�}[d����I�'��UA���u�rA�q�6z/0����l
�|�T	�>][%��%��6ɞ:��6g͘��q�j�>�:�́`�9�6=[m<�*�R�icp�n<Ga���_���m
�G�S��VA��1@�ޞ��)��Х��aA�<BwW3K����y\�㝟�mp��`���<k���ۃ��w;�^�F
x�����I�`I"��5Y#i�z̀F�8(���+g�Wm�U�!ߗL'��k;J������ɩ�U��C����F6:G
3p�6�0�q��xB<HMvmΙ[|j�==���'*�7�y'�(��T����i�3[�B���{3�]���\�`�RRp*���z�m�/�5vnc�K;@k��o7�I��-u{������-Y˺x�(d�������̈�޻�^�gs�n�su��՗�p9	rn�����CQ�V��K<<��wG�w�$`cv���Tm��R@j����4��c�LۑN�SU;��u���ͷ^y5�@"�9T�D��@���Ǆ�A-g�)�l���D��to3������t0@B��D
5uW�	�븓0^����wә_��R�r���-{G,t���^��S��<�U�1;��j�9��ӽݽ{� Ȣ��]� ��D���N��8(���svD����9�z;1�����U�z�C�����Hɨ:��fH駉�ydҰ�£��[^�Z[_4N���[#\��:\J@sƫϖ�%f)z����(�ޓ</�;����1�������6^�ɂ#�}Z���r�2\F��S�|LL#l̦h=�2���`��KU��t��2D͈�ϲF�3��Y��G�"�(���orSdC��_�Za�k�Cn�:#�+�z�i����]O��`�mEuW9��	\*�>�S�M�N�u䩞�ٽϩ�B�h��;��nu���zR�Q-�)��޿_�*�~�S?6.m|7�%�+�T�x(�@�|ߠ5K�74p�){�r6t­,Et���5[���[F�dY���P�ͲvzS��5H+,?�!tz���O�"��>����ś�Щg�+	+K�C8�l��`�<���o�4�ڽ�ݼ>�96z���V��)�Э�5�������펚�91��*���Ob�y�B&E�R�&�N��8�RS��ޖ�y��Qz32�;�NA�7v��[�w����ra�^pʟ�}�9"B~��Q����d[U��kX2���<L��`�Wk,3�p`Y��x���m�2ϻ�=�*��ĳ�0�V�
�W�7����uS��g�f~�G5���3��n�ӳ{V�T6���u�tH∟q- �#�������b� =%o��e0z��Zy�������O^�4Fi�N���TZ. t3�%�-�0ƙ۝��+ؖ�x�ͽtWf�O�A�>��9���mɷV��NL�X� ���e��3z�I�-Lm=n���_f�T��e,j�'���˾��-��tB��-=%Х9��c6�ީCyL���1��'�0͔݉kru:�z�q��5�����x��n9�.t^�\b�L�޸���o�y�Ve.��yj}sNLn�'�"����]u]����� uA܀N2c}�!f��_)T.��s�;H^����s;����4�z�9�dܺ"dñt�8C�0�gtHk�%���
�7{�X�~�zg⻰=�D�<�^Dc�Z���5�lI~��1����h��}8����g��P
$�U�����	z�G*���z6�3)���!�M��m}�8ٷ�2dx��*EXn�7��t��k��5�f'ƛBA0���a�]{*bN�6`^�^�["ɓB�h���MVQ:�v�A�+�X��w��m�d޽=�s/0�t6�����W:8��K9�wd��X�ԋO\����F;��9@p_y�F)�l�ݞ���[eY�L�pq��n�b*j��r/�f��&z����q^��*D3n@�5��W�o*;v	�����&vfV��o�>�� �3��.atD������u��U��e�-���V�d�ɂ���"�~%=�����s�E�}|���rGC�0�0��A��o��S8��[�ve(Kuc���f`��f��\e�KgJ�ަ��ouOƎa��4��	q�:Cl{9�h����C�Py�U@��8{>O)6�?7.�4�~���nH��W������� L	s_Zh1�dSEKJ�2g�e�]�c�x�w��x�����h��t6+|Ƴ�O�r�����ۙz���8�>t��������t��!#�7g��*�$u>��}Ɠ����T+F�:��D�O/Q�gl�����6�.F����V��M�tc����ll�uaw2�&��b�l�|��ޡt�|�c�b�',gCޑ�}�G�X�>ϴR
��uȆ��UWk"2��DO6�ח�;O��r��Q���][.�[��p��[Π�!���*B��/��{;po�G����?���I�J���UA�����I���xfm=r��33�+O�H���8
w9�RWθ�m�<uue H��9f�:�7�ͮ�������ٍEo��0^�o��h�q�%<�ղ���W]��ִH��a�e�F�=MU�w�#+wR�Z�V�Z�4�=�ʣ[i��o�#� �6�E�\��a�ڮ�4{�O�`�&JP�0�eu��=�Ą=����A���R�.��َ�gm<V����Pɰ�\��}��}�l��;��w	y�-�{�q��|`���'~vۣZ<]>����j�p���Q�һv�k�'پ]n�Ȉ� F�dzk���B���;������?��a~�FhF�8(�Z��g1�5�6$ֿmn�M��˫�ug.��gc�(d�m��0�1eU�rau���~���v�_)��[�\��;+�wc/ ��7�A�#)���N��7��u���RY�oC��>%�X��>V�)w�[`_Y��ч����t�k�f~Nr����EM���������F�����;ǅ��u�j=S2X`�m�G���vPͶ^E��{�߼k���& !F�&��/��{ysLT[&����=��!wρ7�N�re�ۚ� H&<�S���?����~���R"�+��DA�����_���1Ѳ*�z�G��"f@&���0� C�0����C
��2�0� C*�
�(�0�0��0��C �0�2� @�0�2� C*�*�(�2���2�2�� C �2�2*� ʰ�0 C(�0� @�2�C*� 0� C ����#�222,2#�#��# �"� � � � �
� ̠����` � �� 0��ʀ� � � ʀ¦d{����   " ��]Ѐ0�2�2 2 0�� �C( C
 C* l�Ti�@!�@!� !�@&�De�Di�&������&�i�P!�&&Fb`���Q!�M�L(C 3L�C"�$2�C3*�"u�=(�7�W�C*� ʰȄ2�0��*�(ʰʰʰ�2�0�0���������~��@D�E�@)32d���������w���!|+����N�\ND��x���bu��/��n�O����TW�������(�+��QX�������@��?���'�����T?�AU�O_�����O���H�ޟ������`o�����b�P�QDXF�@� @
A�)"�e@	�  � $� $�@$$ @	  �� %a 	@D� $H@T� %@� %D��dYU�!F $!U�D% a@� ��	�i�@(��X������'��" ���P 
~��7��?��x�'���?����QQ\����=��~��z��	�=���ht =��#�w�=����*������"/���O TW�PUE�؇�0��"�����������?��������=��`������~���a��آ�+~�?���O�U���P����}�!�_����8�?��I�_����Q_�?����UEp����.̟�~��� X8��`�1�?����<�$����ETW�{������@� c�?�=�����N��/�Aa�����@W_����z���!�S���e5�b?��D�� ?�s2}p#���D���(
�$JE))T�EBU!
��R�)*OcB��" QJ�(�B���BR��Q%JJ�#l�k%l�"
�UI��	T���U(�*IQB��PPE���*��*�QR�URTT�"H@��R9���D�@$��T�ItLj���(UH(T*)TD��PR�ITJ�A
6d�CCDR�QhȢ�
B�RAWlڪJ)*�   ���[j�0k���YAT%�F���λb��J�R�wn���2�K[m(i��T����,e�IݮV��T��b�5���B�P*�J���   X�a"؉l��1���%a�z6�CC#&�7zW�H���Zm��Z6��W�|�����e5KmR����[YE�Y$��@jV�V�����SR�,,�֤�UY*��A$
��
!$�  ݬҔM���[VӭuQ��)PV�kt���*V��5%E;b�a��Z�6&���e��S*�V+kSeZ����ZZgJ� R�!	 ���� sT%Kj#�zGSFSD��df��ͰJڳ&i�H����mhѠ ��f�� )[P�P�D	$����9F�
�0�PS6قU��>��%��
F,[�i,
Ud����A��j�L ��)>�J��$R;���r��P&�P�S
P�mkF����

I��j�Pl������`�Z����V�U �QTHTQQJ� ݊UUPڵ �MY*Q��F����T^�3�
 ��+���Pm�8 Y��(�N�h �*���"��)URT�� ��} \�p�Pu+ hc����@Ε� �w� V�w%[��R� @mCu@Q�B�J�*��%I(�   ��  mCz����  �\  0�l��XҺ]�΀�	�8u@s�p(J�p� �p�P*J�U
@��I/    ��ҽ ��h5��� �8��ww
�%��픎�� (\��Ѡ9��n´��@�p |���U*��h�B)�IIJ��  �T��d��T@  �~%)P   ��*J���di�M��DLj�  �������fE�������|t]�����uCУ�jvϪ���3�=�F < ����ۗy��u�ֶ�+j�mm��Z���ժֶ��V��Vն�����?����BT0�G�� 5]4�-i��j;�Wׯ��c474��	
L%L�����QVD,�;F�7dvް�ݫ̼�t��E�mB�論�2K�J�R�%��J1Pc���v%H�ޛuhf��ٔ-*�1���bu�ֱ���t *,�t^���]�X��54���b� �P�������p�+��JMh�ȗ�����/wb���1�[�T�ٛq�R�`'OYH+���IS7���a�i-����oi˲7!M���st&),q��c@�k�n�="mV\vQ�m]Md�����s(-E�^���,�i�ӕ�Kb��uJBl��,�V$�Q�p�):ݢn-m@�%KTU��;a�It�}�2�:�mEAe!s+a�����K
vD�ۆ�m<��e�M�K	:��ǅ�"Z�!M}!u�+%^��qQv���ϯm1���-�{,loF��0Q���J�F�" éȖ��oV�W��n�˂�\�W�;��/�����!�2�#h�Ź+u�Ǆik,؊�AX��4]6�o�.��;�I"����1��Ev_��	����Mf'��V=�xe���!|�V7R���i��J��I�h����H���R��yLLӵ5��3��6�ya�݋)���UL�N �J�V�E��E\��ѫ�.D���{j���̦,0��K����hܤ��Q�L���'u�V/��V1[������f���x�Y�[�i;M�vqŗyC�V�:�K-+���1+v+��Te��� �����u�:��aU{f*vX�����(l5%&LYdnA�U��i�n�ۂ��U��2��덊b���ͫ�Mڣ��+yg �ԫJ���c*ء](C�2�H�Պ��*,��P��=�h(��ĵ�jm��J�/+0mk֠pv-��
m,Qɹl�Zw���V�-�G2��"i�eM�Xd�:F��N������;�����lه`rbW�9�t�V�.ݒ�^Ң\o�v�q��eM�9İ�[�
O*d%����FGV�8E��1�cw0͵V�2֦�HԷ�)뎈Y�#n���"�-�[.`y���EG���r*��
F$h��{�M�A%��/-n��k&味rHiE)*Z���)н�`�n�4�B�v�5�.���@mIj�(+�4ݝ������D�+m�wb(�Q2�D�^�2��nXf��!6ۛ0�6blV9����(٬W�M5���sf�5V�o@��stfPPMykv��c�	*Py���^�[��٧1bY��1Űlu��	�	K�V(�_��ݫ�I#��vu�Zs"M)p\��!9j�0���@Q;y�6�i�o�%�Uӑ%��+Y��������(�7P�2U��A�p��r5�f 4nE@���J���&���L#r�1��v#����R�]a*:V+I�=�+jRdf��feE%j9wb��7](��ٵ�̨I�Swo2C��^�b��0���D��0�٢�ЦwmX��[`3���i5�a��n��c-:��ȴKۼفӻU��[�.��c��m4I�h%9�nVeVe�D�ҩHbŎ;!ݭ�	j;pG�i���fQ6��D����<�.f�.!�H�jK
�/aC6��Ŭ!���մ�CaX��C���e=�½���r�cɻ,�a^Z�N�� ^�(,:ִ��v(�f8�^���qfo/�
�kV$l�Q�d�T�-X�k6��$p�i|�U�Y���;V��+U��5@)f)F�����I�j�4B��R��0մ�;Jl�Y�5K��\�u��&h��%p8�a#��ƥ��}�Ł�,��1م74:��xbM鍥w��m�Op|�I����M��X�0��a�wW4Z�c�u�[�q� ��l6��B��B�i�:�a�m02����{@B��!���З{b�'���+"�����X���ZY��"���� J�i��*U 4<M�.`�Jӷ-�JU�oFRJ�V�6=
C�2z�h�!^ �b�]5�Cӡa�O�ٱ�L +d�xbkf/UԳ�M�41B����i��eYZ�F�V���6�"�J̙�\˥�Ut�t�ۡ�&dp-�[��'Z�a�4m����V��[!%2�S�r�
�7YKpAc�iպT��$J�p���r���2U^X� Tm]ӫ��c�'Qy��LS��0Ҋ3^��Bh��,�Q�۷Q�],�U�M�ڟ�ͻ%�NE��͊w�=7uWN��6�Lm���QqFZ�ge !���-��*<bȃ*��kv�u6�wC��E�[	 T����������,8��|&��^ċ�d
/ �,"7HU(�����m���Rf�n!x�U�d��dPz6�hn������h�g��Am����Z:*=ѕ�m��W���jѫ6��k�3�8湶%َ��j�0�bZA��q�DT:E1�X=!h�vQ@�]bDj{d�T�A���U�]�
�X^k���SE�[t�Kq��yP/%]ҽ-���cm6@SȬJ�0*��p]Xl�^�P8�q�)�&ͺ��zjњ��6Ɨ�P��ݓ��*���ɢ3j`7�\�zشЂ��F������a���cJ�įu��-E)[�,�F�[r	w"�	IE��٨��4MfM�a�n%.���q�X�
��,j׶�C)�`��E5�A��Z��-��%�����-$�ٸj��Xе`oeD�ͫ�y��*w���m8�"]�5k�	�v;�Z\��hYuy���k�Jt��L�V���t鋹�9����$�wh5Zq����0(-L�Ƕ��ti�h5[G`�0�����]&����SJbRw��̛�Y��7Lb���B�1�mګ� 9-m��.�M��J��M��\�	��-2���6&-/�36B;&pX�!�Mg�mS
�d5c�c�V�Du$�Ph��"����YYtwi\��]Z�Q�@b+/E�L3o�Z������xh���4����d��iؠҙX�J�j*¬˲��y���3M֫�z�KB�mm��Cd�*�z �]F5�y 1۰ U�[vTI���`r�ѭw`���!��#fM���,�/&Ziթ���ēyzp�T��u��'x)�]��2ZyX��ЬU(D�^�k)��E/V��W,�� eg�4nԠ�.��k%A��C�����Mf�3�S��" �Z6LĈ̶h�EHŨf�=����
{gN*�Ǔ1)	���VT7{B����A��]n�tLjjsvd�MB*��L�RĂ1f�!�L՛��&����ǔ�I4J)�Q"Z2f֝d�a�`/�A{v@[L�bl�X���<��Y�ʎ��	Y�Z��ef�]c�q,���*��Wiʳ٫�m��T%�B���)K0ۻ܇���
���� ��֕���B��8ˠ�ixPԝe!B��-��}�"��ڒ����e�<7F��p�p��p���u&�)PQ:��ڧbf7ZZ�ڶ-o
,5�*ZoF��M&�f[;�ST�*Dv�X�E��W��f�3q�(dC����XԚ#bm#{Y��a�F<҅�u���`!v�-H�`�@��R��2V)W0�.��%�F�����AwHZud���^	E�-�H�+*R�Pa<��f���mXo$ #t��`��,�X�m<Nπ�M�ySı^%)�,�,hp�I�7Y���бG�f��Y5�� O-B��dMA6qhw�LAd�9���ЕV�Q�����eDrQ����F[��A�f<VKڌQb�YM"��E��me�Z׺V�v�����B��CJ�R�i���u(��o.�K��D��li�[6e%�i�6�.�U��e�3u�2ąv�e��[N��iY��	Z���h�F�[�6
"�	a��S~ʀS.���5�3ջ����bՍ�	l�P���SỤ̑/��R9��;����8�N˰�p��P�#`P8�7��-�ȷ�n�%Y��HQ�#�K4����+c��Z�>�  �[��bj�F ��&7K�,j�K@x�ۭ�sX؍ҨbT�@`,R�z���c ?��0�/pe�݀,�� �lJ�.��UaUĀ�Иqfj�ƣ�sktYץ�L6^5�^={,?�<7d��ʴUKx�T��V���DU�j]X�Or�;�P�H4R�u,���h$ő]����h�bԤZ�xt�so�3M4/B\D�$l�R�%��Sh�8Y�3�n�e큨=ֳV;���Kx��c'>4�&�u �%X4�۽���v+F�Ն��)ʱI�Û!���JiҶL�*ʢ�Z2֛�e�4U�qhG@̫Ĩ�5j(4i���Ԉ�(^��kS�j�M����4�ӥ���3׍�Y�E�zu��hF���S&b�!��7gh1� �:�6�Ly���C�V��Z٣-'b��4��h�M(����M�f�bM)�e+	.�#@LLK k���X�5��w��2�^m]\�Z���/uWE�'A����	+�ՙ0��`i�0�R�l%�����6�n^�x�7���J�p��m
�S��I�]6�4�驔�o&����p���� ���i��d�H(2k.-Q�&+�s5�+.�b��Yn�D���"�++js^��@����H�!p�G#(���$��Pb��ۍ�q���r��5`�`���d�X�̴��!Z��C7I�6m�V9���V��.�6�V��͎i�y/X�w�l�K1�k%�:[rє��@*s�0$VUdKP�=3(9�=,���l-ۇn���ss��n�M�Dl:Ē��g%�;�M�(V�ʢj���DHRi蛎�PY�q��DJY���	1X���3tEsh�R�;4���y�@T3�_���{a��Hw�m�(���o*V"��v�ƚ�j���F�kiBU��Қ���OP+[Y��í�_­3�� ��-��A�-Z�ݦ��[�$��0�/*��b���� %V5ͺňwH+%m`�$ǅ�v�Ӻ��f���%�l��^��1a�U�N�p�L��3��c0#�j �5����^Z���#�j�%�
V��;z�t1j�c4�.�EL��#d�� Sj;[1�!��U�*eB���v�R�;�Qn�`9x�U`:��%n�MҒ^��d�-'�2Z�յ0쥩�8�&�v�1�J�RƢ3%mᶚ�W2�eeH%-�>�fL��U�Xc�n��.)�v�;1n�B�w�Z�"��uw��D%��*b�"� �ի?Z�v�#�Y�&7*�e4`�pL����[XU�ܭR���BÅT���ٗz�T�Y&�RAJ7V��m�.��Z�f+���@�k8Yv�/`Zj�6����Cu0�C�5�Aľ�Ӏ�+HY��+FT˶�E�+
�|�kؗm9��aҮ��%�yY�j%��R�A|���ͤ�'to]*�Rڧ���0�	��b^��eu�en3����r)�+n���/�B�#3r��K�	+/j�&�� V7�*J*��"�%J�B�C-<�n�V�
��қu�3a	T5�Vlp:׃D{�
�mޑ��?c�i;�h
�m�QkM�,�53%����h����GYT��b�weݱ�r����ܻ��SN�u�Qt�4��ր�A���kE�+]������=R�!vl� Wَ�Rw�0���p^h? �6�[:UA�B��t]e�3��kMűȶV��m9�}q�X�Vh:,[o.�Z��Y*ћ+0�X�n��ѹCtV����EX�e�HTz�c��tq���WOj0k-�J2��(�6X��+j
�%�l��S��+t�kSB��
I� ����l�ųAО�$:v�{���Ղ2^�VVѥ.�yqj�Gn���aϑ4�V�.��@�-��m�@^�*|��A�V��ͽ���2��(S��`C�eG���X�k1��m$�a�3@/5��,�urȓ5$�I�j����Ǘo6`���G���D��e���\I����J�<�ico(�x,�!�b��rL��]:���X��+)����Y@7��
Ŵ�|���J��%�6���J�O0f�F�Yn)��t�l�[���嵦�1�G2��MlV��I3U�i��KMcңɐ[99�M��ϓYy��t��@n�J�ӎ�%�]]-豬C.����j�l�X\)Z�c$z�o5f;�E�4��X�M��hm�age���DI��J����&��jY���D)����]���YuL��V%k�qܒݶ�)Fj�ZsX��êRWf��5v�D�J��!@3vQy.�h���+iD�3CM�e"�7vF�ٛG(H�&�E�X�a�9��/#cbN�YmU�hx16r�#�e���/St�E�z�7xּߑ�T-�-���A��L��q+�˶r��1�D�U�𷙍�r�Dkn*�.7y��Z�u��Y;t@YhV�Y�YVQn^�(� �Z;h\�2F��2j�@SmfQ�ؕ�X/4��M�=��Rs��Wh�v-ID�sN��I{yX�cJ<P�ƒ�`-��BE�t���ۼ�n[#-m$�&FS��V�u�[�YZuP��`E`ۥG5�J�gn,�l�/$KU�Hֹee'�b�!�r��J��[�.@1�R7��]ӵiSk^]Q4#Jn�a�;��3Y ��� (��70����R"��Z&ǈe�v`f�eA��R)�8���m�̍��d�M5j�N�6�e]2ɴZ��U�Tb
5����u�Nض�$ۭ�51
ĥމ#�7�*Վ�F(��7��r8�"][��AE�V6����(�ǭt�X,�`,{;0�mk���4�F'g`�ﶖ �i�g���|�D����G��X�ۄ��dw�{�/�S���&�r�k�B�w����U]���]�S�Qm�ZB7!��לi3�#�MV���P�
n��R�b�eՕ8 ��\��`�C;��9�R�>��l��B���/\��.�3�	�bS��k郕�{��q<`�.��9T�5�o�%#�;8��Q��n��Dв��2F�K����]�e��N�h����jnG9wƱ��^�5[h��*�f�pޘ�����Wj��"�]]ʓ>[��,<��]���a�%��$���%��9��\��p4�D�{Nԛ}�X�q��B|2��m�^�FE����֟�(򈓬`�^>���]��_94��w�"�V�a�W)���,fu58:�|mے�2Ź`����i�ozk㮣�*�pa,q��f,hS��M���<����s�y6�V��ǝ�|1���Yض�u�t����U���ϣZ-�}Xx!�n����ů�R�gaosS������=^��<׋B�е�fַ�Gh�D���<�t�2*N�M幌r�w,�@6��#�8r|��^�s>��v���qQ��+���s��:��s�ř���3Ye#�z��+�����]����P���{��	5��B�����z���Jf�Y6�m�x��r:����6LӽS��權�ŝ�0����sul�;���h,�R�P��pσ�o3H����;�R�4g]jf���.�G�i�0V�`���%��hrP������k�TF���i�j�o_��lo������&Ԑ��
3ہ�s�7��v�O��� Jm��{vR�U�wG�@�o��^Z�݋���8A��պ.9V6�nv��#J�̽˥7���)���kfm�OV'w|�Ŭ��]G��-�i�K*$m<I��+~]�u�O�,M ���^�[�]�TjȽiҍ�޳�CTom��0s�-�Să��m)9���T�"6���x���a�PBZ�Q��ssn��A���Ҧtڄ���oF� ��S�0�U|~�6������/�G�M��(s�j+/�V����xBȺȘCKd�V�r��\���ڗݮT�6֐թ�m���5�]͝�a�Y|��}��e�h%��\'d��.]��W1�­�[˦V�_
|��e�Yo{��^�O]�L�jn�
�G�R=�q�+����|�Kҹ])fc�=�MqH#��%h�qH��ux�ض9�B�_o�ޗw.���rp���)2�pr����y>T&��h���ԥ��+I@^���7���x�i�p*�ʳ��.��@yj���8�C9sU'ٽ�E^�{���8�Abۛ�I�-qlu�U��1���;k!�՜�g�M_7Su�6�]I��9���S��K/�eI9-BJ��S��ސ���Wi�Nّ�Bz��1���A0Ŧ��&S�"t���u�Bk�7bp=B��(��.E4m�N.@m���n�f��rŽ[3��)�Æ�r����	���Z\����_4+s;в~&ٴʢ2٤�t���8��C��m���R�f��倀�u�ۜ�Voe�7'71���� �z)���:/V�t�af�4*����e��Ƀ&�8�	�@����$�}{�E�	X���6]�x���\�%��J�[wk3)һ���Hw��NY�����f��9��"��7��ul���v�����3�d<QT��鬮Is�Hs�+&�WhC\�J��F�$+�Z�b��j�Ŧ�r���ҡ���[��+�#����Ɨf'�W}5F���5g.D�2U�y&��a	����Ju��	ͮ�Wc[��N��s|0�������*�-;��3h%b��h��"D2ƃy��w~�jec�3��zj�T�H�h�.]3�^	��ڟ(��yʏAg5���G�.U��C,�� �>�3D�����u&b]��
��>X�Wuv��ʼ�JN�6����T��b�o���ܹ�YqI6�,��ˡB�>�X0h�j�sV�p��v���+kE�����KXU])M7e�����4���Yz�V�T�{���W���X��Jʻ�O��2�b��
���F	�f�EaՂ�L�lKw(��%�VW]�	���ƕ]¦�9��Ż]�i�3c��]e�;|��w*�k�J}(_H��t\�:^�.��д�[�Z�-N��+1��wn�r!ۧ5�8O]>4���]�zr�ǻ��PTyy�77�p�wݱ)�.u�*bI]��W&ӥzE�2`�K�X�eWb� x�C�؇V�<��^���R6���	P�:�����SUH<f)���
�z�;j�4�t��h�����iq���o ��Z��1j��I��v%S{���*�*:��oj�a�ZLX�ns�唓�}�:qqf��^��o�!�Y����m��n�n_lv�{wy�H��Κ�mi�(e��\S��"�Zkm��=�l"�،�J�eE}p�-�������oo���&\��R� K��KZ�M�n6pnv�m���ⷦ�s���>1к����ޕݥ�`<5��}V�j���~��t���O��,E��L6%�5ŀ��5:�Q����»H��%�2+gp񹥈R��a�UK��c�F�ڝ��4����r��;O17���x��t�":Q��Ycr�ҋ�+�k����t5��@�a��Mڣ�"��آ9�Y��<.��U;�6U�+���5�B���������ަa���`�w<9^=XA#��3Ui���u�h����L
�=��-�p)+;��3��	Ȫ�M�h��X_t+vk�H��Wq�ÄM���""r췗ud6y��[��&���-e�[
�p�M�ܫtV��'t"�V�q��!d̓T*7|��(H5�Kd|M��Hxh2���L��,޷��PrŢPE��2��O�����D�\K��Ag2�c�|ܻ���Ǔv�*�˨�^������ãwط��yuh�����Zs��Y��퇻�	woٸEߐ�<�}~:؎�Ɗh}~0��l��9��]ˉ�T�V�>��J�#i4{�҆К�gw$��0N��*b������C���r-�,�ш��jK5�w���E-�i��(�He��8�τQ��U��{-����糝c��W 2=ͩ���/OD`�{�%�������υ���H�+A���S��Z7����к �,��w3�vN@��K���9��V�4���i����C��ܵ���N����9��������q릵�YX��[�W�Iڴ���Z;+:�roO��}�v̄Ki�N[�2��+G�Q�;��2�0���a�w��ܵ�_��}���Z�]/q�.iB�HX�J6٤�q��P�WeN��fTu��0���ʝ��4�=����X�R���sv3��SE���=�^��|
�k:�LrH:m��w�ޛ�"S���|��������y��*����ԡ}G(/�v�y6��Eծ}�/��e��������Ҁ)ɢN��_	��f�˴�5͓qNo	c�����"��Z�+�*�U��aey��o/z��ǳ�:�h���&�ݫ�'mS�����p����q-U1����ِ!���胸��gn��	����`�kR���4Lu��)�2��&�]+��a|��/��Tу-u� 9ch5zv�<����W�U��l}hT����J#)��T�x��ੲx܆U�E�{W�[��T�,5���,����4��tӡ���w��]����ia��Ȯ��{����8Z�l�34k��%�7�*d:�z��=P�s����_��5����+4ͤWj�\�o���u� ��Dd6;����&�^�v�Mi�J]��U�K]c�قc&���¿�8�0f`e�탷�|˽d$�-[t��6M��(�x�V��w�N�Z��r5}�*��w=�����y���u{��*�m��7P�8�Y���i�jMc$��N�����V�Ak�&��j�s)�����+���b�C��Bj�_KQ���
Yk)Շ(�6��B�i}�3d=��l�	9s���%\�M�:��A&P�z,��GE�v��XVC�s�ԩ_MՋ����N�!W}���I��k�[9���i=�O;Oz�jyi��.nנ�\�<�~ɚ:"��벏Y�EW�e�/x�7��c�srs�R�6vt2���Ӗ�ԩ����s��A�I#8�b�ݱL��m�1�!&���{���^
��Z}��h�Qa���V/b��ЫM/�q��ۺK�X�;�g$E�2����y���uطE��ko{��1Z�r��ؙ��5�P�w��/�A�MP]�FlF��Y�ÝA�
v
�4�ۺ���+|�* �qTƳ������E65Va�z]ob��R�Y�1�ŧ����/�)��Ǵ-��z��U�[�,c��lD��������e�Ԏ=}�Y-�]�ΰ��<�=FP��i�a��Ia$�⵱��'t����Z��n�6d�P��7���+	���z��Ç)Q�֙����nvV�z��q!DWi���L.�t���y �:X�F�jQ�	�����n����N�)ˉ�;f���j����X:�$tE��z�|�gUe�0�!\��]���F_{Y��R��tqjk|�nK���&�cwY,E8#�[v���[�1���b�u�\]��[e͕+��Q�(�:y�s�C4���񷃡b�|1X�˥K���r6o��7��[��:�C��g;�[��s�F�)�g,���Z�:������HO.��+��U���B�g���R�J�кQ��\*J��c&t�v
׽v��_�mv��?e���q���W0��]:C����Z��:��f�:�x�s��T; 8վ�I+U�5C.���J���W�M���PN�c�4�j�(
�M�d�*r���]�͔�^�fG�.ґv�P�8aA�WK�Y��0^!K���aμ�v#���\��0�*
M��[/2���Ȥ��
Vy0��J���'�%���v���[;؝\}oY=�Cn�Z�/�|��Z��u�q�ng+xԃ���"���ȝ�zhYN �4�r�;¶���i#Y�)�@A3��lUr�x�^���ח�<�j������(tx�ei�L�TRQ�͒����;"�g�t�H��}̹4�y�����s���k���'g�p��+Qll�ۚ)�w2��w��Af���@��Vl�vX �vol�%H�1����v���:�5z��u���aY]P��v��ᕲ����c���픫��v%��|�_#�P֮K0��T��a�u��Ä���^}8�4�;x�ٱy�.YOyWu�dv��r6�3�Պ8�aA],&���Pջѫ�����[s�6v�F3���+4���'�f�p+��M)�x�!���3��[�|~�������Jz5���5e�++4*U�r��=�@v�\������3�����lG�:DB4�V�:�m�� �l�.�/.u�_u@M�t�_B���/"A��Uu��|`��Ѫ�oZF�!�eN�n"�R���QmJYSuvAZ���N|+/#cL��Pro�lJ�%������{��2��p�����
��{�C�/j�S��c/�.?��U���h��$l���.��.��55y+#�«� ;�$��Nv�T�`�V
�{V$]�:+��(���R���chu�-{h��)���9��'���B;����8ks�:�:FM��Mmk�J�6��!�\�i��|N���vW
X���2P.�V�5ql�#n�Vܪ�K�CUwB�VT�I��u�r.$W}&�v�C�T�FvZ���^��H]t�f�Jm�z�ON-�)w�X��re��lOkv>�j���5��ĭ�)������g=���XWl�o���aI�U���33��52�@�5��t׹(yS�Q�CF�asPެW�$�z��`��+4kZ"����}a;|c���.����.bۮ|��+���AoJM�lU\��ZI.���B�G8H@��AaE�~�������ѣn�X����!��W���U����݌^�z�f�9�d��Q�)�ZJ9b/0>|BqP���d� ��}�k����) n�b��=Μ���Pyw՘�$3��:�Y�S{��٣G�4zwV��j��(n�h�3x �!#:e�b��6;Jŵ[3��;ʶ�ٓ�#T�BZ�m���@Fq݁x��b�wa���*�U������;���'K��y�f�q�Jk�雖��WgM�]o�WNwvI1�V9��e�e=i�����܂�o%.ws���l��ʄU%ݎ���|�\�o+mz�H�_o-�����t<�ٕ�5rt�W�O^uٵ1�k��ۙ9i�w�]�Ym��Y�wm�2��������c�&ҕ��u@�mM�I���!��+��d���	ۜ�c�3Y�ϥU�+;BRSϸN���%,28���I]��y��i��%����>��÷Ҡ�D��->5��;�s��Ƿ�|���cT3P`�A�*���J�4���6��Y�q��곈���IW�|X��o=�A���O>�!J�;��	���_;���3�}��"#=�Q�i�89�h�w6]!�e�9��b, b ��ԫ�uu�wQl����3�;��?�̱��l�����"xt� �b��_|r��mf�2�`�A>��I	u���9[�s_-���&�����${�[#9�!��s���=�V�<7���;�-7��7���$�w[#?�+�I�,���	Z[� K<�L�Q`��g:JgI|eԼD�&=�,�R�ѳ��+7�)[�f����]ݼc]o3c��ܵ9�\���IZK�(��X�������������C�vO�@�|2&�eNA�������E*��%������6ii�	�V ���@�Kl��tI��EX��j�.�Sڜ�:���%�Cm���k&
v�j,��Q´5����&4�DUa���{Rʠ�V&�S*\��ʎ�oU�����V��z�DJ),�b�r�(F/*��m6�X��J�#�-�{��]b$�ʙ�Brer��4+���I�vX��ԫ�<'�gJ�%��:(�h0��(\ �]`Ԭ�!Vn-ʺ6^<g0�G#e�h��PL��,�Yܹ�7�uv��M��Mcq�Pۢ�6��'I��ZN�2���\K)�p�ܦՊ6z�z	[X5�������w02-}�II]�6�B�/f�9�-�}�S��Xq�M�ؗ1|��G���L
�N0����O᝝B�#*����:ڦ�M6��L��TWL:h0a�T���S��.��.-�dذ�죜�J̐J[eS��U�����:�λ,!������;ݼw}n�=���k;%�x���k��(*�A3[G#�%��7qR�C4�*]%P�x��]\a7��a�Z���2��q*�Y�
�ٗ��&1;��V��ߦ��#��v�0�T��ē��/뜱w#}\��k4�]�6�P� � �h�����ƍo�v�j!�͒��Q��������z9Qծ�]��O�e�M4��sD�V�+D��2��#XoZ��u�U��p����.��My���N��6@��m>�9[Ҙַ��Y:�X�:�*�¬C(��S�b�d�U����®��IU����;3���*?�Fa:�<�2����KmX�+)��|wX�� ����L84ڋ ��W4A�G���hTS82]hyn�4a��>��� ���T�݌Į�
G���u�5><��q����ԃ����װ6�
4ĂJ�]L���]\�BG�����4�*�ab�l=aC�7���%���]w��-t�e�i@M��5��&\��J�֚�uwi�7v���<�XHR G<]�4s����`����s0?"� ߊ,�zw�a����d<��b��$����V5G[D�����lK,`�v�_+xF=<��YG�).i��")��q��Hn�+v�<���kE;qپHt���D�uc���Qe�AdI�V�ќ� n�Я�q�W|4:u	�y�xk��R��=��칲������(���\�����n��<P�R����m�ʡ��Z/��[�Tq��Y1�y�[�9uIi�'�s��i�	 HX����K��[E�^�$CH9`K�K0!��?��_����+A��@�d�Q��î�C������#�{N���5����$Z�r�[����c���_!���߅:\�W+��+,�+-UXd�%K/�M(l=����[1d�$B�m�B���/�a��Oc�h�@�Ghu�m�|�e�W��Ԋ�]m3 �]n�Qᎏ6��:QzUګ	<��yǏS�lj��~�p��ٷ��TA�d�O*c.� ]L7Wr"�����i"�-�YͲR��F\�y�n�	�+�B�(��,��r[B�^Z,eq[���Q�w8�;�"��q>����"n���+kF��ia�	V���f��z��k/П���:J��/�����W'�J�{�����9��Pzv�����0er��M�[�}yC��!�8YƵ��ƫ�}WF�����AX�����׿lyNE��#NȳfXF�w�)����Y:�Q'����Fh��ow+9֔-���ֶ�#\�i��2�T$���B���uۍ�ҙ��j�ܫ�O36�V�6&'IKF�fL�$bْ(g(?���oS��y�;)V:���KL��B"��x�	��<�m����s���T�LEb�5����-��U��F��
��1%��]z�S'F���vA�.Q9IS�[��+�`�7M �S���e�0\k��i&�
������Ԩ������ڢ6
�(�mb����h47�Z�A�����qԝX�վ��^`�.��OF��|K���%��i����; ���᫹��$8
Œ�;8F��|���)o��X����V{��ӕuoMd���bK1��p�k\�y�M�̫`_0.�Hs����`�&�`��'1�6�ko0�1-������Y��(2��)md��<T���j����0U�gqbhn����[�Be��q���͡��=x�B]��G����dJ���ܠ;� ���,/���nW}1l�EQ0��MT�:9ۂ��,���q�R"�yVGО�3� KH�U�Y��K��mȨ]&U5Y[ ��v�t�f��s$kU����ퟄ��"[���n�v����e'��$&�۬
������Y'r��{@<y��&���k�u�����-Y1/�L��;5�6�@�s���d��S�=����诮��Z�P���Y�q�u��il��T��8Q𿹘h֜��3N>�-]���]�TDW_)!*)(����������*!�H9����+v��<�V��L;G][�[�ĝVw\eZ�u�QkeL�6�y�����U�Θ�b��MX��yS�`�k�����Ą.ɤn���n�u�lݧ��B�F�����:߁�{0K�k�*�pV!;d��D�ҁ4]7	�F�-�ܬ$�9��s�.f��+�T�ŵ�쓵���7����T�����O]�±U�=�J]����c�CG�E�`8���1.�Wu�#��t��s7���*@	A��ץ`�7Dfl}Sy��&Ue����b�x���ou��WT���Y��ܫ؄ݕb�F�+`�5���q
�u���"��(���A����;0���*�]�����s^�cڡ�wcw��8���M}`�P;4�$�w��Y���2���V�7Tȇ05��$���?��@�*�t9L˄i���$*�ܭ�9�=�ה+Gp����xnK��}�;�m���J�
aY ,�݊pά|{�F�)\˭S�Ь��� bOa�#V���3hP<tȍg<�!8���3m�A���V�*� Ft��ˊ0�!7�z+,(P2�@%]��g0��EH=�!�!�K�����YC�A��Y��B��{Y�\a*�L�WR[TNef!}KT���*I���9�d���2j�-u��m�E�u���;&>�ȵ�a�Y�MYu�+t&]6�.�w4�/J����+θs3>[N��*4�EtP6k��y��Z�M�발�>���H^�輑�+A�MX*���V:-�^�`Op\���i�i�w�JZ��NoiH�D,pi�)�Kx8[�K:@;�)p��1w�̻�صf|�D�7�:�1�)W#�
�GfT_u U�p����7��
����؎�t����ׁI,�
�`�Ca����*�p�w����M]}[HV3�B�*]���i{�,K1
ZͥYo(�]e���2\q��M�o%�$	�Vp�vZ�p�Y\�V,� �+vsU 7o�`Qe�Ԩ�B�"m�$Ő��fR�3�O���d�
��%�&F�U�kh�;b�W�����h�ãvcr�醰;L^�9
����X-1�+�9J�m�UQ%uc��e`U�R:0M.T��䥗�Z�
�Mv7��I���ޔ��Uv-��eF�.��բq�QH�N{Sm8��if�v���
� �f���!�}"�k_s"
�MO��M�|�B*�]�<%gfR:�ip3y,����`��R��2��F	l�i�	�3{V�4bAƠb���8n�EY�X���T��khՃw��ʗ]�RkyL�W�z��h�blЬ�7^XCT�V� v�,ƶ�M>Ԣ�"���]�j?N1T�V���T#�E6��
�Os^�܄��;Ppq��]��R Oiñm]���y@8,̳g6=�*�e�TB��J[ʫ���i��U_1:�7.�8���ŋ����Ȅd�g�D�7�f�麫W[I�r������$��T���f�ֆ�&V�:��$����W;�i�Q�Z.���L՞���b��I=�6�7�*���-��EhW7�۷*�%�y>���u1�Rn�9�"��b�+W-�޵�	��PΩ�@�\*h�V ���I�

��P��%hA�뛒�z�W��j�=@;z��T��i�~�$֯�b�ѱN����o�05����иr,q^�j�o����n���u�J�++�qmT�j��9�[�a�Ac�p��0(evs�N�^����[5Š�ݾ�!��f����X��u��k	�e;b#�)�klS��i��-0`��6��Y�B�Z��l��&(tXҶ��(>.ކ�e�hC��h�����%x+�њ��Ug����C���*��iF�������#5��V�BK��O���]��W�g��ȨJ9Р�n=��fʾG*�,G"�7#]�*��Ԇ���eĵ�ګiT�ς���pp�{hVv����r�kn�0ɼ�nÜ���t�Jn�y���S[�&՗	�Lm-_^PWq���B�⌴*#��[N�x:��l�j�u�-��DF�,U6���(5y�噜���]n�4�!�W�fi��&3j1B�Ҁ���8ex+e�2{������@�.������x��5n��D�x���Wc�s�^I�
�a\۹��N��@2��`%���Wf��CS����٧Lu�!�ok�NؕŌأu�P�-c�@CyP��6/pc5�����G&��$Tͤ�K����Y o-](/KY�k��n$��*�7n�	���jS97���ps�<]G��Vw:�P��,�B���Mn-��}����9��-y9�t�`�g�fh����kkE\�����V�Z�t+�[��o)5"aB/U?�<�w�����di��E[I*m��e��B�v���F ;�m�ys:3�=o���]>1�jʊ�^\�+`���*}�6�U�dۂ��02X�_;=X�������k�ۻ4��K7���q� Ӎ�#�ƶ��N�p�t�`��cp�LS�
�W��������7F��p��q�w���؂���T��pyK�m;;_�YTsv�0���,w8�w�*h�΍֮�ܫM;۹W�O�,��J���+u������ۊ�ӺV���8'�m�8U�F�(8�9H�Q�+�/	��)��t��o�@t�yc��|�7�]�p�y����i�D�6;���s�F�:.�/Xu|r�5���C3S+m}�������w]jY��/�a��ёӽ��N�&�h������QL��<.�Cz��%�J��Cg�fա���5�<��+CF<�.EVῥ��1	Ctf[Z(B�EME��ע���VWDz�л�ʆZ�Ҩ�T��-�d����
R��bu+{�7��k^J )DV���];y�#�ˁ�('F� ���̮ыNu`��,m*����	M.��qEK�,����x=gY�>"�#�����V�IV��+�ڈk�E��t�d�l�&'�^��#36�u)u�Z.ŀ�i��׽��&"�9���V��e�]�c:�5�ư�,� v�[q/MA�;T!ͫS�VWp|n���!�)cʈP�4�5ZY[��P�MI��x7	�8�F���y���!|��C��d��0N���:6��a��Q-�����c8%�s�7\��)s�h�cq��o� �O��t�ź�|�3��#�֒,&S$��[�
�
9��[���J��n��9���<)�'�Hɩn�� HԄ)n���kF�jˣ O�SB\(q��-�4��HttQA�Oݏ�Y�B�]4b��V*]H�����98�͏�FG>��j/1�;���-��]dՒ�v8j�q[eu�>����oA\��*ѥxv
�D-R�{*�B�E�x*&�����1hb��.DT���w7*0n][��݁��M`�1��v��˺]7������	��n�I��,6�ԤΛZ�O`C2�@ݴ!L
�3!H���X��;Y�Ƈ|_H���	5'�E+N�Q��;Z�73o�Μ��K��+4���um��F�����󙪊�8,>��g���% ������窉�*��6��,�2��ׄj�L0:v���P�J�7h۾DQ.)q�W^���Z�qO��u���[Y*�̜�'*kU���R���,�U�[W-:�&��Z�k:�:��9t�����b�^�x�WB�W 1WjNb�0i̝�a���hq8X@f`��v�@���2��)rAJ�-nW�ڭ�L6����z��Z��M�Ɂ��lF�*�p/70��6�O��dL�(�3�y=����=����"� g��w�_�ͽʵS�?o4Y�v@�V�}v�һ5㢊��Ʋ����5�1;ϸ��x�K����bÌ͇�1h�k`j�ڂ����N��v�TzU�+4��)��c�ڪ2ieR��I;x�����s�U��X�h�Ӷϊ$
�ȃ_�cU�Y�y��`�(J��s��ĻXH1;�|������4��h�d	!I��{���,U��k츾��#/Y\��kyp<�G) λ�+9Q��9]�P���C�m0��*���Й�o֯+�l_R.�%�
�7���wX��ƕGrѥh�j�̐#[{}W�4Ůgv�ݎ�n�h���h6h)�2�+(�9���w{g�N۫�F� }b;�7WU�&��9M�U�]H�ܛ���(�cI��V�8Ge3:���H�-еZ5�t�8���&��v���;(��t���������Xh�T5�Rv/���`��[X���%�T�&����������ޫ�J��{�=sx�/�J1h8�W5��r��<#pr���pz6rǳ�g���LT~���gY�*��|��Q�h}4<�K����0����6�hvT��o6��L�\��GwN��V����m��5cn��u��b���x+���m�I���O����*5mn<F���N�e㶛Ֆ��p���ױ%"�6����F�;:��\ʳ"��;��:�����f;j��v
۬wKW6-`*h������6*/Y���V�7['$n�7�mwdt�͈�YȆ�ut�i��"�yh�*��z��x.e�L�/h���I��ۜ�����u.�vmf�����dk�N��R��~e�VB��g>�z4���ձ��>9tmC�F>!�5b�@S��qDe��ޗ�vËi����^�v��M��g_i��mJE�a��T��M��<�@9�J�L�]k�+y�6^P�R� E#܆���
�6�;A�����tT#>���C�қ]��*p�y�����.�`�F�+&Nc:�`��_,���gfv��M�SS&�UE�8�ۖ�\N���S\r�l1��@����P]m(���ċD���iF�>=�g{��%	��:�۲Wz��G�Z;3]��3�7�63H��
ȫ:��Y9�etX��#����b�󫮲�}5p{ۘ�slδ�6�%b��n��ܱ�ﯿ�o��w��ba�e��"i���$H�Q����$�ʒ�A"q9�61��d�I�
"�4f�j+c0e&$���L�a�H"��Qb�0�"bT��Q	�%�ɒ�h؍L�Lň�$�H�IDl�H�1��6�f�*M���"#Rk���(ؓQc��bH�!d�E�[45!�!�AI���ѳ3)6E��̱�J4lF�$�ddѬX�r�
$��Q"�)�r��9��
)��b"60�ř%b��h4Y"ƃd1��ђMI�D�Td�%�d�LQS"f�-4�&�	%F1&ɤ1�H���Qh�X���4�I��L����DldЙ#H ��Ti+E��(�Aa�bf���$�#h�,�*4Th�,��e�e�ݺ=z����^����R����VjC��"�ꑞZ2�R�B��uL���I��h��>�78��ŝk��=h�@�/�S�_1ܛ'PK*��GWh�BegÞ��+�f�F�S��ݩ�8��Dڗ7�=3�ے���~^��pߴ�2|}g�q:����6�o��Y΃�:�ܪՆ�o���]�I�=`�GI�����]3���O�+�k´#�՟�~*�>�t5k�D����"z�ut/�z�2�ȧ�_6+��:�"��
�EiD��9�����_T<ï3�ڡL�R>b%�Nnˈ�}a�uJ���q�9U�EU8�Y[��Wib�-�RA�tWy�v��Y�=B���N'fQ|��V<_+�1}M<�9�Π׷M���鵷4�2+��4�MT��X�7(�<O;�_@
�G�iy9��c[�ȇ|��{|�n.�!�!i�S[ie���UiZ���&�[Ѐ?�NC;~^�1]@���+��������r���v	��=����c�-S���B���ĸC���.?:ƨ��t��c}�+�ػ��3U�<�2��{���^J�}����*��5��1�N��\G[��[��:���u�]�V�cMk;���'�7��5z���{��Łԕ����\�Bd�9�<��\�:��ٝGj�w6�ik�+{wY��n��w)cW4E�=.��h�V9v�dfv�I':����(�Ml��uI�V��^-����-v��9�i��q�.���EIF���T(o��d���Svn�u:�1���b�-9΂�r�]-������t���7�4ό%��m�՘I����q��(
x,&�Խ笡X=+Uv�:��C�V��HB\"r�cK��1�Z�t���}~���0t�Ɵ���[.�Q\v����P�	PrOu	�кu��y<.��B�ݤ���:`�@s|��}`��~�{��x-L�,�[��`8|��O2}�*�S&�nb5�j�o�#	3��*C��'���).,�[�k��뤕GbY�CӪ��ԝ�#O���(A����xf��q1rZ��O����۾�ihj,��h�Uj�$X͗6MC���J��4ת���Kk�C���O1V�c^�0�n�:��'�s�!�K����j"/\�2�A�r��CFct��{70�=iֿ=�v��A��i9�����s��V/�x��G &��3_�{��D�h2f*���N=��39�;�:����e����OF�/����0��K��ze¹D�����Qm����W�iȧU�\ 8�V�e�mu�����t�^GQY���f�Q��h֍�4��RG��Wi�/`�yo��h��$����7����z%��i�]%�YX�W�⸀��vX��N��Nq��Cn�:�<K��Es��Nz�vW����X��M�҂X:4���k�������s���6�$�5O���҃`��Vn[+ v��aH�4�@(Э�hQ�GC��kS���['Y/$�P�3���mҗ9�R*{����qq��a�)�g��
$B��/M��Jo7fb�$�g���
��!�U�:ڥ��ס��x\X��#��;e�A��j6f9莍;�:�o�m��Dp��g��WPG��1ʾ�*�Eyk�~��tC�|r���G:L3�k��pv�\"_)
K���J�b!04�`�Z]����Kz+�v��8(�������K�r��v���)y�E�$O��	����6/��=����x&��3�2��s�2��[�a9Ň3l��؄7��\r�O+��<Vr�m��F\o��*�g>*z�(�p�a7ei�ܨð碤�䝚6܁�ѡcK�$�Ou���{0��$с@�{�5g�{��6:�'+�-�*D��lMo�ш�XgdV�c�*mj���H����^��?�C1K�Mp�{Ye$�vx���|��)h�V�\7�k�(򬞢ph��@���z� (��ށ���&�g �fUL��{7��']����"�)��,�5�!F׻����N����s-�N�#��gssvU������fX�,�JB�w���;G]y�r��U��T�_݊�4��[h
���]����z��S�q�N�l;����{�����3�
f_^��h�Qk��C{~^-hz���ৎ���B�W}���
��s���7�Y(�� ���7s�lδV��-��:�L�D�#�W�u�}4FF{��8J�_k�G���@]�4c���VWk\.���q
�h	�:����� ��i�
�u�w�u׋h�B3B;�&T����<~c�_��>�Ct�&[:��C�b��G\^�\�xh��(]�5 (�q`�S��{��Qp�Wp-�ưB�X�!j�����b{w2��{�9�FyE�)���t��ρ�>!L�h�bY�"�Ϩ�O�Yz�?����G{$���.
�/mߘ������O:� �MP�_n������ȉ�-�Ǐ.�]J�������_�ݣܦv��,�t���Pu`�u�n$N�mN�ŋ�,V���C����	b�6k�m-e\9�Kݾ��[ONb��w�`��\�ӏ�w�P�S{(�m�o3�z���9��(�]qT�`[ƒ��hi� ��9>\�r_o�x)��&o�Hq�p7&�tb�S��NHKh�:� <���|=���te�7��_N��C��yoWG`��0A���x��t'%�31�d�J���h��\��_@�<�>,��e�bU)
0qp����˭-�,�$Z%Xf�$*T%�&��c2�z�C�Nl�t���[f�#��t�i��q������T���KP��ku42�Mc鈺�r�oT����T���P����k�3����s�q��WF#{h���b���y}(Wxb5��4��3Q�^D��O�Ӏ��b�n�r��u)��s�{���{W�1ԥ�L��]�Z�Fč�	eظҲg��nP�C�����7�X������>D�~�-��ε~�)�����s)��:��W��.��5n�p�C�X���ky`��r�%FI�>r\"r�iD^�k����5G��v��N/�en1R�Fk�Ds�b憹�aX2:=�X�q;2���8Szh"Uk�z����^�������o�m�42���\��S$ӛG۩puՁ�s�$��N�/���5�z�[
c�l���t�b��v�B�p�;�.�_z���Va 1�ք�m{��C��sR�[Μƫ�� ܶ����'�s���c��P��O�x��9�>�4Ws�緬]w�u��뽶!L���k3���=�⾀ҏ�������kc¥Y���o��p�@΍x1���M�N�OԵ��^y>}���谓����`>84� �^Z�YM�g�y92��+!��H[���^�8yc�ȹj�e��:�&�q�I�Ip{]t�����Ȯ�c��9��롣�LK����|ps�e����6�u��q�"��� �(��lv2�.!��y�`�����;u��E�,u�uöTzܺ
��(�OV�<s�J5(�j�8����i �S4��<�h�����W����{� ��h@���^Z�������u,���VVCu�Io=f|(�����	.�q���[�H�#L-��S9�_���=k�<��]_���qg���̦{N9�>�WoWX�.�ǂ&���Jq�rH�9{*
bx��09.uNK�@��tu|;�mw�3�I~�xo����a�,f��s�_r����	�%2h�m�G<�5Q�E�n�WO�k�1���%h!i�����Pz2X�COY���Q=%��:�TXV��s��Лû��'x����>�|�S����]0k�����Kv�p�eL��N�S�o�\%��
e�v�]K�[� K�Cw�A9�;�;5����t������1T�gM�����G��;qX6B�Z�,,	;�Fy��ɫr���l�������{;�{��+��A�PT��a���ZH�*h�8��t��1ƻ���[���XA�5����4���\<��3�ʰ��`�0��V��]ޗ�Y�
��v�{>� �O=�a�ͼ�Co3�+���U���d�hB�E���EVK�N�"8 �ol"^�u暡ٻ7.�fX�%��WM���X��uW��<N�t�Y��?7�S�U�$�]�tcyݷ/]+b��Փ".#����/�<�8�z�vg�����HUD���hf�G��MY=�|�r�Hn�D�^�uaT��Q�6ܶR����~���]����*H��g>��_����W�+K��璔��jEA��ǻXt�!�#�ڰ�<���k:�S�M��U�d�\��
��$�8��$3ʻL������^�'5�bk�h��0탻ϺRT�e���/��8a8F�6�u�5�.J4#�z@2��J��'�Y�{����W-���Q�{���Ӵ�/CJ�f�)�N=�t�J�Iꆛ���vZ5�I޽�C��>V|G��;/�G�"��`:z���Pu�����M����p5�e�9�;�RY��������wAc�Q��]���	U��=��GǎwuH�����ջ7o��|�Ǐ�K����=����&U�P<�u�OH�/�P�s�g�sK����y�E�T~�9����Ro3�����������	up
$�:����" �=&�Z^&�TJĊ�S���c�<͈ނ2�.�E2:�<��>����q!�Tp��o��2���5�X�������Z�::�=�z{��l�L��䝚6܁�D�햆\t떞_j'�S���nuNR������3G�TT��e�/7d�����8�\C��7. �4v=����t!%U9ڔ��κ�4:Y:0���n��Q^�}�<0O���'���U��o��J�/i�d�_��c�)]�L?�ƅ;<N�L�;���hđ�.3�ҙ0�� D��m%I���j�su���L���T�>>�WPr��h�s^����Y��çӌ}��q\���4�Q��8{�*��P|�i2���Zj��γ�����rPF�:՛s:��2�����u�_fs6!z�j����CR�Yǁ��x��^�̟w�q�:�g���*�*�T�����X��\�ݹ�1q�k](ssZ�v�ZǺ_m��wJj�)ԋ�lTct�)d:�S����V�q��q(��کһa��L�}Y�`Lx@�F���Y��(sP`��@]JI��U_\��)���k]ݕ/�Zyޥ��˶��������/
u�����٨k4��EAӁa9l�z�t>��|��7e��c���$;̩F�D�����4�L�������z`��bB�*'$�u^�Md´��nb?w_�M���B�GQ�J��P��0R=�v\��(>���9`��G�g�vz��s�"1㨅��ީ���ߘ�%g��F�h�r�_
�8Omg��@��פ'��9e��W2��!�a���ڿzs��8�$W[Da�T����9nL>�lo7��]�4���z�;�m���a�pr&�U#0(��/3k�]�;l¥��Q�,�1>��ME���8�]�=���(�ڲ�@�J�3^rΨw�G��S�f3����K�a^G`J�҂�4���]3�iP���Y��}S�JY/�j�W���t=y.�j�s��"�сq΀�d�z��`��BWV�.tfXP+��X�mv�eO��t<��y�4��߅�_2�0��F�/�GK'����P��k�s��."��_K^%�,PІ^�CZ1��7��c�z�:զ� i���:Ŏ��l�����Д!�t�%o�m)V�?�<���c�ܔ�9���-�:��MyVT����*KQ�N�����W���� ��&�8��8=����K��®&M!	"7w��X7b�.'��&l����ҹ�C���(~on���9d8�r�2|�]Ս��V�����������[�N����Z�_��xE��̭j�O^��<)��&��d�*:�J�k�@}B�)�g��#�����S=�^^o�T䯎]o87ozgٵ�L�C ������ǫ��O�vp��ON'f�,p
oMM~�_��߼w/nT���<�+ݟ����t�&^[�3m-;�?��}'s��-8��X���z� 7�|:t�~^_�׷�Ež�m𭔼�xe���kHf}p�G|hʯT��״� �8�n���cyMh���kU=9�>p���l�������аA�B��N�ʈ�}A6'�^DlL��k�ʞ��H,�Ң�i�o�s�84�F�ΰ���2�Tu�J�7�<�a��P�n�N��k�ϯ��3��zh�FE�r�i�1��d��!@AV�b����=L$��^���)C�b�<�s<8ʀ��F�	m_�C����q1�f���7�
�m����A�)����ΐln���o�y��v�t|[�݂�-�7���[L�G�D�����iKي��M��t��m��%euX����=�%�u> VeJ3�v�����6��j��������q�͡*R��лb��ދ�9���G����Ƞ~7Yr3�kΩ*��{r
|cn�bz� �=7IjK:fk���)a5��sK��meJZ{� S�Iˌ�=!��,��}�/���[��3����T���u˦��bȸ��vHǒ���.8k��l��4V��7���gD�K�S�ٛ�d�c�����̈��z֖�٬nP�}�Q '�H�:)��8��}�!�5Q�k�ۻ�����Vs]����%�8�q��mHl:��z-�M���m�ӟ�}�4E.W���С���%i�Z���-
�uNt:ݢ����oM,Z(^���M�/Xs8e>���ŵ_na틏 Q�E��[�!�}�Z�f�xmޠ���Q{sO��SY]��^�(;X�qn�.��N�d���t+�ʷ҅цqyٜ��I��-]��J!�N5���J��ҍ�3����11�鑈�\��%�u&�}�0v��z��5g)>z�x:�q��r�Ah��]FU�'�6��9P��JŮt���{{�;Z>���]�����G
t{r����)5Y�V�vB�t�n����a��em:.��7�fk�}R���pC7���0z������R��{\=�\�����P����L�|�du��کt#-��v,�����ڕuj��R���H����'U<aH�����N��i	{W��21�r�%|3�,2n��`_\�ŶVr�B
ƵK�3Go����9J�c����:&7O��j���{g,+Q�����Lv���3T�Ѕ�t��mhcQd�*��Y��㨃�1��Y@�gs͝���+��h�+��;����+fc#�� +;��԰QG`;�Ð�è��+UݗϪ��b)u��W9�l�m��:uF�,�}��_�Pc���e0�ES��՜ez/����&>S)q�/i��ݚh�t�np�#��mc@��+nuj���f�-v9t(�+�tl�c]�u�b57yw-a^bf:vnH]v�p�6�ַ/��m��}"�ƬfEB��y��NZ��VX/+��յ�J��s���WJZ��sܽ+�
\=�t�T��h�@�\OA��nv�M��K�x���wm����r�a|�jT{u���}2ՆD{���!���Xk�u�h�7~z���y���jGF���NM����������*�wO9�[O���|���ur��s�^I��74��V�o��u�y="��ߢW�����c��i�R����-7z3/z��X�̋I���*�໭66j�j�:�B��>�����ﾻ&6cƣ��KB+�Y�&>�4���(ь���lF�D�3`���2ѐ�F,I5�@�nr�I	���F$(LB�$B��F�أDh 6F��XC$"Li#I�a$Ԕ3F6�lmNsk�Md���+�E b	b��`���3$lEm�EIE����I%��ZA*��I��Eƹ(�L��h+R\��D�1��)!�1��S4��54Z
�J� �F�R$�E�Lj4d��5*�.L�-"�ōd)"1�1�Gb�����a,`��"�)7QXĚ)!4m"�"�E�%�*4QH6�Ԛ�EQ��s����*,m,TQ�Ih����n��w���P�Z"���WWC�8lb�o���˸�֙h�!C��w�Av�'u�:�]�0e�c�OW!V+��q��8�E�տn���+�Ѻk���z�Z��]-��5�+��[��+�scq�}W���|m��h���9�����t�w�[�|l~#��xC!Ǽ�ʈ�x�`�}�!��D5��c_�@����8���~_����K�o7?u���q��K�W�<�k�|m�sx�o��v�u�:�t�]����[��WOW\�6�Z�w����KŽ.��z�tߗֺ_���O�} ������������7Y�2_�DF��C޺��b(}􏾸nX�7���Şs��W����>ߺ�������+���Z�t�W�n׵�;vѧ���n-�x�n/�t5��?�"0G��D9T�kjv��F^E�m��SW�g��� 8�� \	���Ly@鼿~��^փ^��~�-ڸ����]��WK���<�x�k�q|x�^uս-�\W�������t�[��}�kO��=��_��{�  ��3�0���⩕�y��ǌzc�0<��gԏ���,���F@��oT��p=�1�c�{�/kF��������������>���W��t����~���t�_+�:�o�{ LxFc�q������T}�t�팬�.��܃y��F  ��2b-<��׽�]��ۊ��K�o�M����W�z|m��W��k��+�~��М#�Ǿ�x��������k�����$|}��E >�>8cfh�S#�>.��v���Tz��,�ic��T.��|�oMt�+��U��o�w�t�k�]-?r�z��ǋ�n��뮀p{c�2}�.�d8 ǌ{��w�q�#�"�D)���'}}"k���.��ʜ̭�=����`B���T��}������y޾5�j7��oK�����[����x���|W�r�hߕ�qxߕ��o�|�����ŽW]�]�#�@a@��S& ����]�X���kb�u_l{�� ᶪޏ����n�ם��O�����ߞw�6������:����[q�w�>���۶�m��.��t��s����������u˶��-�{޹x�5��]5y�����JR�r�{�[C�2� }�E�� ��"x����2�>���H�}|��s;u�-��^u�h/s�/~w�}W�9|o|꽍��z�����۷M�=�}[�tۥл�t��q�[}�|��?]_�b��~�2�/5��]�O��?�͞���� �;i,�mf=��B���i�@v���񗯱F�)%�kWQYWKnX�s`����H'&��w�*ߒ��{�;+vTz��V�r�I��w������\5�:��*t�e�{*��V'�pR�ȱɗr-����|��|����k�����������޹�v��~��ݭ����vߛs�j������]/�.���:��x�k��y��{Z+�{��X���t���:���Ș=�������'W?J���:��<c\m���]sW�ź�������\�o8����O�p=0�{�� Txx��N��ʯZ��֋��V����Z+�o�������//�c�f���Y)v�9߿=7�������W�qo�⾭Ϝ�J�t�\n�x���nu����Kt�./�����_}sһZw�}����|m�^�?_�u��7����η�zg��D}71������~�Q�.�E����������W>r����=y����/kF�W��]<WK|�9EDW���띭?scqw����>6�t�{�Ly|}�d{c|\��xDyG�l�X�0G�,ǎ�+�p�S�����w�5GX����<��ޛq�{���_�}t��y�ίK}W[t���]-�q���5���-q�o�~�w�6��v���]7s���Lws��Es�_�r�7�����WM�|xL�{b��W�N�ɑ�N�G6Μ�`x���K��w\W���o߼�ޟ����y�[��W<^6���;����͹�/w�:񷵾+���w�Z��K��]��t��-q�vۥ�ߟ]�ιtѸ؈�F}X�Xds�|���]xg��6Gw�u��˵�_��W��:[�}]+�nq�o��W�ϟ{�.����W��{�������߼뵾��x�/}y�]��WK���_��^�.5�������ۥ�� dTL{�c����>��nd˹L1����0@��7 }�}�.=���]���m��ݶ���5�\�Ϳ����t���t�ߞu]��\o����ƽ7k���}������zWJ�y�V�QF�c�g���{q�j�)���Sڐ�2>�B>�C�D�q�"$|�����?��Ѿ+��7_yoj�i�;���7�n7��5�v�m��/z���qo�1��%r.�@�sW��2��1�~��$��"�}F�;/ab�Oe����ҶkXq�G�&�t���H�}��M�nu����vߗMt�5��]���׾w��_��zv�k�]5���w��ŏ־���W���۟����>��|�A�H�˺y�a���B�"�*?J��Y:kڅd8�rCm��0W-�[Zet�ŏ�%�J��ej��h�]�Mg(��&sx.��,�yD�;:`J�oir��*������Vqw܊��̽]D+��zqۋ4'(q�=۳nY��zb�!t�u�q��	B[��_�\Lx��� T� /���_V�����Ϋ���������5�\�r�[��t��W9׾Z�~W��������~}�s7��� L{�&�� � �vM��Sy#*pF�37��m�����%����^.5�s���K��n��{��W�x�9��������^��s���濗��ۋ~^�Sn���9v���\���.g�L8�D��#���q����~����,vym�6ο�x}}�$}��]��x�k��t���}U�؊�}��꽭<����]��7�t�K��]X�|}�Dc�@p@���
 ���<�Ңw��n��m��U��t���c�܉��LD���`�o���G�"��9˵��[�z�����9�/w�m��v��_:�m�ns��|�Z #0=��1���G��	����]���-������|W�t������c�:L� �
O��[����B>g�>��x��J�.7���s|m��+��M��j7ߞ�ߕ�q��_�o�|�oM��[���^w�F�n=~�E��׍pow�:�kx�]+�{��8�:��{gɊ�n��FqU<W򾮖�־�꿛�v�+����⸷�{�b��-�ﮮ�[zU�q����]����k��]zWJ�n��e�C { ����{�@��G�c��6�p�8��AN`���?��}��>����z[���m�~󞆢�7��޺��}�7�N��.�|�st�Z�t�O��띭�]k��_U���5Pzc�L(���[�2�G���K��/h�u9Z��~�q���� 9ޯ���+�����w�^6�o�{��uzU�����O~|����ݫ����:�k��^�&.=�,�f��=�O�РTj�6�9E���Ϟy�����o?��z,ݏk(��}Zb$}��U�}}�?5����V��-��wߝ�꾫�^�����-�־+�����W>/W�<�oj�\o���Ϋ׾oͺ[��~��w�c�DR> L�D�j$���ԴK싯nwUS��|G�"1����Žns��/���5����U�����~���z��\o��ߝoJ�^.��:�+�v�7�t���Ϊ�k�\k�NX��@�`�D[���>�DDP�u����v�y��~ݏ[��L�/]_W"�bp���7w�:]�k�"U:MF�� ��r�幋W\ו�1Ȓ8]�d
R��X[mqr��ד+�/�=�4�-I��n̕i�j�q\��ut��.{��G��(M�l�4���eΝ�Д-��c��O��o7�oJ�]-����\��v�J���ל���zmǻ�6���x�m��R=P=� Y����=���n�W>��?s��^��.��9�zk��H��8�E3�{��ss����D}�<��z^+�ӾoW�+��;[����ѿ~�\���[�]-���ny�v�������n����*���m����~ۦ�[�q�}�oK����bޤ��\|���%��w�pz`Nsg�n��ns�?<�u���9˻�+Ǧ-w���o�r�o���n��7���\����kF�����ץ�_�_��5��-��]�[������+��������]9�o�P���|�D!|��������H����Q>#�$DE�sB7���o����sWM�n/��W��M7��[��鯪��:�~_`\��=XG�yWq�P���y�:M~t�Q�l����PW����:�to�jo*�G�9����g�h�8g�"���W��]tfԮ'O�l�ε~�2͉�y �؞��|��6liP�a�����Ti#�Q����vNQ�	.9�*#��k��X��N�r_�×��}��o%Mn����Kkǅ%�\P�i��N̪/���}7��'��޿�:�c;��-?{Z�ߙ)�~����9.S�r�ݥ}8���Z]VN`wX�ǅA[P���x�xΣUm�AUW�;�[�p4�h�����p�;��4k�k��{�SE���y�޽z�����=(���W�6�4Cu�Mc�{x�;@I2�&)���l}�Y�����	A�p!�y�����\|�X�W\65w3��q���G�LoeԒ�C�A�Zi�'C#�z�i��b}X;�\�(w5p��{�O'fN��6�9V�A��Yֱ�a�U ��R��]=84���t ���m�,���G`���λԬ�Z�����K-�e��W������
9�=A%o�{��/���5�PPɶP��Ƅ�ꂩ�-e7	E��� 0<-x@��}�.�����2���厗9�i�.=c��W2�:#y�f�w���EO���Q<��]��x�}9���\�lw��`:�q���zf.[w]����u\K�v�H����"�k	�K|���`�����Wl��/,�R��w*Ώ3Ը�s$H��T�.5��lAv�N�Y\p��~fS=�]�w���p�����T1��[T�����DlZ"�$&��j��ξw�����y���Krc�;�1�*z�S-��~��������b��S&���#����"�=���+�%�P��n�v�mr�¼,AͯY����qZB���ya`Iݢ1��ɡnP���Q��&�\۷ƍ&�
��2������ȑ�臇"��i#4�h�p��=���Om�0�,W�B��bxϱ64�p��,�X� oB�F��<4?i��:�#yS|�h7�Α���٬��ÜV��ni
;ƹMu��Q���q�Ey���Q�Ї7]P�u�����lr��À�����7[&�;$��Go;��j�`���ʎ�l�t;+�lW�����P�7w��{��.,m���}ʬ$+�nW���XF3����^3��m�>�=�p�����}��yU��Ln��c��n4$�W�̅��U����Q�L�6��I��Ê��y4�Ԕ���C���1aӠ�8�WM���X��~ӲE
,���&Vv�n;������l���Xg�����+%�O3̽^y~q��=v�9�Q�jNƋ�$�SUږ+t��v��75U�X2SKڪV�0�>�������Y��ec�~�Eq׶�fo]�,6�xܬBw�z�1E�S��Ί���Iut_�n���jEA��ǻXt�!�#�s��M�+�׆w�7{������{5�񯭏�$�+�T�!���+dt�Ϥ���nz��a*\Up�ň���iM~:]�.D1�c�g[�a��=��B	N���+3Ы����$��1oS'�_8�+}��z�㾁�{e�
�U��tTJ$�舄Gz �4�`�H�z!n,��ٌ�����o�"�ފ�')�rg��6����.�D��T�Ҧ�IO�sُ}Vy�o�P�}>y!>���sϞG�&𹫓�Fc�p���aP�F�o^��v��~�֋�yr�D���(nDȢ�c�ޝ�&W��Gx��βf1٥��h%�lޤ�{��e����:`�ǯ[��s>�<���rי��u�.�0���X���'�  �]�v���.�@�IH�f�lߣz��.�Fӑ��˛d���H;��@E��of?g_���貊 ����KUpA��N�v[�d;s�RG4���܁���"��
V6T9�uӧ���!���I�<OTd�hAvC���Ī\�e�c�:ݓ��m�<d�]������~�=%��l:>�*���,j� ��T�<�$T9�^�C�v`~����W���sx�3����U��.U9b�{ʘu�4)�g��w��q�[��5�e9��}�#JT�q�������f�[�2^�\�s�G=�������L���&�^���\�p��s�3ьR��~5-��[��SI�N�*5�����s��~�VF@"�]�ZGf��9��n�_y��؅��\J�j�<�G�v����~���ԞW���1Z�����
�[��8
��4�+!Ǵbc�a��}^~�k��¶/)����78��óԐ�5������(�|%4�L��𮏺A]�*R���I̺oor����ww<�0v�,�5��F��U�����垱�x%F�o���V@�zי��꤅��ۣ�s,�k�9Mu�ԣ9���;f���,�o<�̔]�|��O:k�w�2�r������V!p��Ժp*��;?}U^ː[�v�꧹Gڄ�x�!m�~xg;z:�Dx�:I�~�=���vۻSiL�}�:sS�;{�l��s�<����CƲ_��}�ֆ{����ϐ5?�뵼tv�ڃ�g������W��y���ڱW��;d��-�1���8��$����f(E�<��C��N9���]^���@���]���F9����dRn���왞4F;�'�wޥ.�=�.��+]D���}!�X��
��{9u8P�mYd��2�;4�u5�޿�d ��7�ʛ6�X��*�J���4py�i��J��G���Dq�{�.�Ý=ҷ(���nu2Xe�cT`\D�:GN����yB���ӔC��4H�O����,���7$l��hIu]D))@a^�3C,���z��i�5�N�ľ��y��۾(ٕEQ�+�	Hد^�|�ޜ\�!ѱ��@�on���9d8�1}BۓѲ�Mv�^�-;7,����c��� ���Z�XS!�9�\�����g�W��"(˻ֱ�y��o�"r{��G$s�1���{�Ի��3�]�$���6gm+4S��+�\���v��:�vb��jt5us��f�5��_7�\�6�;����΍�Υp-;?��p�7��B�%!�-MC�����]|���c]Fx�y�U��}�|Oqݗ�6���ᇉ��FNB����OC'/��E^���:�`Z��u،^��ٌ�1ΖR�z}���(�+q��
�V���{ON'f�	B�7��='�r���us:ϔ�\y"\��c�������,��P�J�8���=�}�O�;��q��VϷy���Bʊ��LV)���)��]7<m��;��� `\�C;~+��}nm�����\�j�3���b5������Ӛ|�偎�d������p�(�wM�	�K��Pǝ��:�t��������iSӬ�+K��O:��_����y���7�����A��D�Pՠ����lo�o���=�X븱�cOvޣ1��}Ρ���G�b�W��Ӵ ���H}�`<)yk�������VƊt������է.�q�W�{*��&�'`�}��;h�5���YB�z`�]ޙ����ʻvާ9�vDEC��n!�D�.5��lE�x�Ldg.5�`��G�YaY� �	��Fr�AT�d�-��H07&wn:�HEnաO:���6� �;���*a��ک�;f���r͖�ȷ�S����VЬ}:�f.�:�wja9����hm�.�����o�ξ*s�ˮ�X]���}����1��V��Nwj���xy���ùss��|���$^��94u�^C� �8���eV��U�7^����2ڻ2 �ޠ��Ӹ�=L������U0��M����f3GH�Ll�9�{�/:�1�����:+�8A�����{n+6B�Z�,,	;�F �|�з=V�juԮ3�Ѯ��~����<�1��"#�.C�#!P!�ȯW*�FiP�A�Y�{}K�2�m�x�+���"�ЯW<����Vl�
�@�ȟ!�)!��� ��ڈ��{���6{tՠ����(�����n�5���H9���>*��>���Eb����rTg�*-���Ŭ��H�bL(��_>��A�p9�����9�tXΝ�*�'�	VEL��ر<ѕ�r�9��U3b�@h���b�K,��}�y~q��=w���;��2ė�҅6=��0�^'E��������[9�i�v/u*�D"��r�X���Qv�ԍ�i7�ݜb�H���G��� �+@��(�3��~��r��G�;q�å�_�1�m)x�:K�=��A��&���5���;�vˣ�F���J��)gI�Z�)�ue��9�Jf��5�
��
q��Pf.zY�V+�X�N�nXz16��A+k��i��#s�b�p�ah5��q�;��J��5A��mѶ���2r.�F1�c{�o4r�U�:p-�I����8���r�.�ڊ�
�ܼ�&^C��{ʈ/�:�>��7]�|g;���w���R�]�h��}��k�R�r�՜�+M$�d��}����u����XS�p�q)�a��9m.��Y��P��1+Ie�ǽ;*���t��w�c�8}Q�y�ٻ��z)�lQ��ʮ�c�& �=�*���]����Cqr�N.)T�n�<��zSܬ�J�Y��#X�,�����C.*�-e8�6��u�\̔�7p�7�=����N�&���5W���/p��1�a7;M�k����o�7�@����o`�C��{��+ru����gl��z���J����+6�5�)$���o�^u@7�c#�>��Pvk�6x ���x���>9pƩ:4��f;���|
��>��b	t諰Vh�7zv��-fw\X����Y�K0*o>ũ씬Y6�O�h� v9u�PR�# �ڸ�nwJ��a<&7Zx�wt��*���34r���Ww�F�rph��#��D�*6�ﯲƵ�4�k�Y�
If�>�4�H��t�k4*-��K��U�]��T`V�v����r�h�'e
Ww�T	>n;�hm��\+2��K_e;�R���;pM�ɀGV,S(�͍+F�4�10^l�6�%���F�8��C�f�.�<�u*y+n"�ϴ�d�򓙐�IHi�+�)J�N�9z��LR-�j��x��"�n����Z� �m+��j��L�$h
��w/��D�{�V��{�W���%�DE� YmN\*���q�"�%9d�LP&��P��ř[��ѥR�3d<�E͈�Ù]���)o|'��a�%�+�R��ܝhȶ�	nf��?�k���[g)�q|����h�[؏t����g���|X��D�tۮ�W�"�)�P��-/)l߃�BheU�w"q	w��;Ur�V��\�۝�;��� ��z�-7��ir0�}�+��y�[\0���k����l)e#WMZD���(���;��/�}l;+LD�����Af�az��\�Ax�i��o�d�ɓ��`�(�sjm���N�f���meio���Xz��ɬm�S�d�صU�#���b7{$�7�L�>��
Cԡ=xF���x�z�̩�Ma.�;��SS� c�BC˴��fv�!F�E��Zq��Yj�dl�Z5�2����*!�}Ҭ�b��=	�RE�Pw@I�E�D�Ůa�%�2��Z�x���zs�]P`���;�V����WW@a#5s�����vTysaxn�AF
�-�����>�+�+	�ch�t�"-BTTcDE���h��RcU�#6
�┣Xe$l�#Xf�F��k�f(�����d�F�n5��!(�$��E0�4�qp�E��b�ې����b ��"�1�)2cE�%���[Db64#RV5.9��4X�V6qk�cF�E���"ljK2$�Q��Ƹ�Q�!h,B�J���KEأb1���pX����
���b��MHZ�B�A�����j�s�qA����c�9�h�������]��������r��T}�i��QŠ>���I[%r�[��f�jۥ�M
�]Z��@���E�[��TR�;�(��Lx  ��2����W��w����{5�|on��0tW ��C>U�u�K��`cwF��d�ӤEG���q�_�M�)?e����8k�۰��,�oa��H)V�̫�6wx:ѓ��L�6ʜ��C��b�S��G�9��Ѥϯʀ�|��<��"@�+jkL�/i��8��9�*��V�ǂފ���G�@l�ɸ;�����\�<���> .;j���^����d���z�zr3=)��^�]n��9�3L���DF��k��ѓ=5i��_.${"��[ժ^U��q�EgJ�c�чnz*H��;4C5�_�e�eO�Zͩ�@M1ƅ�/�\Y<0�pAvEzWPȰ%K�VB�u�'�-��o$S�^ɵ���0ˌ{��yx]V�U/�Ѡ]���j�e�c���P�]zf
"-,�|�;����T8��qmU8\�5&:r_��P�\hS��l;��]:�Jŕ��^���j5N�\_�Hp2,f�f���� !x��HB���u/��h�s]F����%�����n�ea�=}9�W�f�TNL�H;4pP�7��C��(�ڈi�ϵ�=�SËyn��2�1��u-����=�Kyq��pS�:��%]G��m&S�Y�yj�Ûе���3��v�ի�fu��쒫vbD��تݣ�܄~�������c���{�~�;993�MO"Q�l���5#'�꽷�{�������;���8ȃ����B��'X���O���Lؔ_1�WTqp:��j�<����íz\�Ό��S׺��o��.
,X8]
�[������^��z�&=ɏ��x�^BǦ���,Jm�|�5 <��{)�C왌�\�5 dy2���[�υq2��C�Ǣc�G��Pw�m@���c �$(��Ql7~zl*��Y%IP|7���=���	Wn��������-i3Ǜ��K7�OД�gG9�F�:�Zm�T�ߛ��$����3W-��z��s��w�i��E�=2�]\.9�mX��q�l�;Kd�ζ��]:�g<6��u�.�q�6�q��1eT�G��!3�;�\ioWG)t��^J����3IQ1����n�+�X�E�fp8�n٘��%�
����l��	<�j.��8�]�=���(w�vY֦�V1��#ݮㅂE�\�/��ʔ�J�r|��lӤpy�AYu��|��3}N}���q��*�6�U�.M+��Hf��7��b�V��NZQ$z��l:��TX�!t��ѝB��тiY3�K+Hg;V�LE�:��F����<!��V�ާR���m�5�=׉-�<]dAe��Qy�F������VA�B�S�򾯼<<7�괵:ݘٳ
?BU>��2Xe�cB����<Q;@A�Xo��
��$v
���t�;Yݏx��
.X�a@����`mUѸ�bPn\F������H�K'����AM��2Ѭ�3Sw0�/Փ"���Rmm�ۨ��}��f|�V빰�������\��V��uoJ�DxŢ���Q�]��\O�͌�W�����<����Ny���U�xM�X`�>�<M[�Z9V:U5l����nV���uׅ�ꕁi�.8������m�V��9x���w��Y-��q�$\�i��q;2����X���Z�L��Ҿ틶�^A�2��z3Ω��׷M׽oFm��j�
� 0W���lڑ�L*iָ�:�"�ª�!�c�O7<�\.vcU���3�:I�@I�t�F�7�c����g��$k5�G3Aj�=��ӃO�<�v"ĵN7=+o��FM���q-�E��]�gNZA&�����ב<~�ƨ�i���i[ボ�;0��(,���9*r{�E�=c��I�b���l����)!� κ&5«s���"yS,|
��hsN��u�kL�1)@���v�P#�
��n�g���I��>��g��,7���U.�9��H]y�Gם�O�RS;���d�!d�tq68t��� i^���P�@����%,��$}wէߠ���6t�Wt��]Rg���-����-v�m٧B�K�̌������|ۼ�:��}�HB; T�; �@[�1�H��ճ��hZ룣+6��S�%4��g-�=^q��F�u�N7@��4ϫȈFx������&�Z)ߓ��Y�tGB�����O�X��I�QO���n�"���7F��h����B�:1�.G��{,ɵFc4�?o_�W�(��T�M�AyC��)�s|��9/���q�l��C
�),�H<�"��r�iZ{�W�mP���S&���Ds��Th5s��.����~m���e"L5�׾6�S��p�T�W��ۊ͐�֫�N����m/N�s0���F�g-��� ��}��U�ZhB*�U�f�fç��T5�ny�C�u�tf��ofv�z�y�5~?���8�;U�I̟�*��#^Ä�m6��;�>>�(�t��*٘�y���fY�69S�!�1�xk��q�%V��t#ܾÝ�{yQF���+Cj;�s:nW�2�Rie4�}��Z�4�Xa�p�*�]T�����E���d����,X���Od*q�X�1�ϴ*��m���X��)�ܙ��!�fj�%��u���r��;�"J�U,ۈ�f�5k8b�x�v,}��:z<�H�����h��U	~_gj��s�S��=�b4��:.�t�fc�<4J{(�|��o�7�=U\����+�,�k��}�/�:Þ��mJờg�x�����2�3OT\���I	�@��$��íTIϺ��R�eD"��r�T��0o�<�7V��:72|�����N�>/爃���|+����#��s�0]_zx|U0w5{�ݬܥX6z1��Gkɫ�Mk>�"�(���t|�!�*�2��G�^P�ȭ�:�}'��d��C�d�B�0�\t5���x"�^��!�R�' �S;ۢ�tw'N�S��hSܭ����3�z4�~T#�_$y= B!ܰqE��M(7/1��s�۩����7�;�`>\yoEz���E�p0�n�����{M�q��=Q��ܕ:��/ѣ��4�E�`�1w���պ����r:�f�/��˰�N\�Jkl������CɶLV܃�		��T�;��+M��F�=$)���T��㸼�`W�J�+�:Y�� �Z�/jԭk�+E��KZ��у�b�k;�W��$Zo���T&�����H^�ה{b�Z�g M����{Y���ko{�/����>��M�i�e��r�+Y������o�Y7����أ��eTyW���=�
�Ⱦ��S�]��ؤv����=��>��dT���bT�5
0i�FwbsI�Qx4ϺԮ�,2��7. ��9u� ]����݁f��'�ם�)�>��t;��Z�j��`]���l\ed��2�w���j�\T)�l���U�����.*3��zA��}l'Wt�q�jF@ȿgKf�m���A���:p<�A����g��gl���\�����b���v��$Du��wYU��Kd��2�>��*�L�tEF�֚�t�uvd��1??�����T��@�#��N'�O�}2��X4�LiQ	F��:����26�E�6�s��{����{�κl�x�XV4נ8�eE�:T`���ҨE3@iO��EM9��VOAͽ���Ez���g��C�f3���R�@��ə d޳[� ���|����L�]^vwJ�lW+���dct[�Q[�<<�6_+88o �W\5=+�t�V>R8�1:��	
`�۪��[>����a���#���Lm����I(�r:[B�u�U���8J�9�T�͜�.�S}=�O��y:��ɇ+wK6�����]�U���y��.�	I��VuJ�5�A8\r����p�{����? ^ZuہoA}M����w%MbC�RFY��Jە
u�ʑ�K��巪�țݫ+UQ�<���;�v�9���R6���|+8�rc��t�Js�r��\aW��������l\��/1�=��D��Z@�_e�� 9U��L���ז�tvN�#�h�Jc�aȞ�w��;9dt7���WhȜ���"��D*G}���W���;������{"�<%kt��r:�v�i�='x/�V�X�~�	V��i�9MEqI�s���P!^�&�ѵ��va��T��%L�qУ��/�'DXs��
p�B�����{�.�7��ˢd׳,(���j���1�����3�x}Y<�R��6�(eѻ[uR�s�RYɸv)V��/�⒑�[���w|s˝D:6�g��R�!�=O'&�۾�j�]�Z+B�����Q�^��N���2�t�vey
3ޭ�ހ�7~�q�K�[)n	͑|X�.���H�(rd�+�NQ�I�d����Ez��83wBC�T�N���޴�ߗ�[���1@�{�܋���Y-�2��`�+�x(U�����Z+ƽC��|���X@q��U����\��|�_���XQ�I�2�w���(+$@T�T�!V�P�j�N^��!Q���ʻ��S��}.�-��YЂ�s-���)M�������}�/���Ҍa�Ǹ�w�}P[۶�Y�9}��x{�yգ-���b>��9iߡy�6{<׷M���c{jx�Y)Y�\O��������k�Xsi�\مe�u�uT8��b��<���<�]A��S���ne�G���0Jtn�lCp�����T��״� �KU�X8�zs�|�����j�n	[z9���",˾(���D����I��\��>iq��5GKӡ�����n���84�F��PU���7�Zo�Ա-å1TLÞ�먁��!�A`�����9��צ�[=gr7���t�V����(�����lB��s�]u���@�tP@�a!���]�\*ϣ����ۍ[�P���YRw��;�q��w��:z�3��F@�TN�&y�Qfs7u��<���^�X�
G&��FG&�B�n�"�8�D�n� �v'A���ĻۻU)��b&�(�F�v���ڱ�~qK�P�*JnzB8��}Ơ��~�|�'P�d����2��%���Y��=�Ô׼q���L��_��	��2h��u�o	�D�Nl��7qޑ����=�%�]�(�σt��Yg�ɒ��z4�Y{~�s��u.�]u�)�N�@F7! ��j�����-�0���Ք�96�]oGٝ�hg�ŉ��}ըZ�9
:��b޴-e�V;��Fo����Z�0�����HM~���xZ��v�9f�+���J�U�S�k��z��?Z�~~�]��^XXwh��50\�MdҮ��-��`�,���d<�!.����WJ����"��i"��*��A�w�6fm\�F	�:2՗���z{o�/���f�+q��C>찐�?V�y�<�
�x�6J�+�/�龣�_��N :��N,#,��*|�g������C*�b�t�wl!a�kp��=oR��)�&.sվ���Z�â�q;t�������'�j�ڮ�`s���9$7Ht؇���u���^U1�g�ѝ��R�Fx�ь,GD2��u��/�:�s�5��՞��E�2���<��`����M�҂X:SKڪ}��F�v/�՞|�u�Cj-������ެ9�����8����dW�= �U�`�xʈ�+d�Z��;�{+l_z-kڦ:^1�-1��-�JQ�ХE�\B:ڠ��@�y$�#���!q����{s|�q���Z�K���=����c�.:۰�E�f��zL�#�0s��t��f�<]�-�?L��&V%��t�f�`���]��	4�w����Ytr���o`Aд��8�93qeu�V��]�+3�.ȷ�����7n��(V�Nz��w%^�"j��W0��Ӳ��[ō�6q��JY�x =����Yi��y���C�tW���V%�]���'���g��O�<�|i���{B��LDF�kiA�/K�>\k�z+���G�@l�/k ��"+]G�"t��Z��ãq7�Pْr6I�����BJӑ�)��er�to���#DTܮ7mD�	8�r�g;"q�Ȅi�A�^3#��(�;��Zo���~P��:̐�VK�y��vt�oE�!��vh�r�F���xd��ꌟm|��K�Ճ�еﷶ����R�Y���c�8Rݻ�E�Wt8 �G�%}�j�g�@���r����~	</�K���:�V�iSg����Q�b2�\w%�[�g��p�1��yS\hS�<M�,b���Π,�NK��[�܎��5��`��s���jF@ȼ�L�;� ��kU!��]A����!8B��j���i�]�ԡ�A����p�%٠
��u�Zl��%ِ'������,���g�O���ލWIݰ���	w�׎��N���ٸ�a/���l�{P��m�T>�����Z�]�SF������U�Y�E�be&��ٮ�l]2f�K�v�㽼���PB��u�\P�X�E՗8�7��nŬϔ|��F׷�BE<t�Ŝv�W��s%�d+(��H���
^��'r�2�ݛ,k�*v��	��­���o>�t����Ol�F������!���f�P�+Cji(n�M���t�O� N���Ή�u}>V�&��v-M��aZx	�b�ڜ9��n7u;j.�]�r.�BQ� ��8���Qva2���]���b�l��P�(C��Zeʘ�E����z� ��R-��b.�/�#Ѹ�-q�H�ʽb�❯���CKB��vZ�xWJ���m�N��]�\�CyO��6��a��:u�'8�ZK�umgV����&�_H�����u˙%���-�(벀f�S��yjV�:3�j��}w�Iц��p���<[U��	�E�a :��h���;�޴�Z=1_TB�Z�*%�[��{ݩa���SRMƇZ�CGeb����Fvr�V�r�N�CEDg�������I�>�X�_�˲ܕ�7L��C5ms��.���l;�ݫ�˸%ڲ�,]I��y���6[��x�8��:��.lg���#�;A������C"��2ݲ�s��[���	B뻧o	QB �}º�����;�X�A��n��z�gk`ĂI��e���ă�M��kkB��b���e�G4
Օ;���ouM��a!�u��8:ݣ@�Sma�8,��C�*�s��i���&M���kf�.��'3vpnn�<����#�܎^	���kXg_u�B=n��_�j�ˈ@r��)W�J�V��%l��Z���������w��gS���<����:N>��:O%¶����ژDpk�t]�p�yjz0;B��uэ]4O�4��ײ�;쎍3׸;T��t8vg�!�����|p���[H�R��>�C���e���(q�� .#)���6:���
�Y����[��gp���X��s^Q�@pqU�R�F���UH#���xa1;��ve��el{�v7� ֦����0XC�Բ�)������2��n�-B�ݾ��Ħ�7j�!Iz�vjSw�Ζx��)�A~��j�z:u
d�tY�@ �G;^�%X�w�z�(ӏ�L�:��j���2!�]��R�09(�b�N\'�ҎY���+T�I�
��t^v� ��O�Ԕ�75(�'k3#�_\˓�!�Qu�s�^�!Hl���Wu=������[�j��(w��2��2ht��2k���uG��	.�^� ��:I��/�"�ظ��g8�c�zv���{w.2�9|2_S�8,��C�Avn�+ǽ�x�6&�M����E��WOt�gu� {�l�ܥ}i�nT[r�
Ժ1|2���et :ÈZ;ʗײ�^t�%e�p�u��iV�]7y%�ew�U�l���H��"��"
*1S"�g�\TY1�� ��RQ�1�F��X�E�e��eF��DV���*Ɋ6�&��������h�h�E�k�\c�\�"��Bm#Z,j6* �I��lcs��
�F�J0Q�эF����ѩ5�a	���Ci*61DE��E	�5����H�Uq����&"�Q�1�m����{���=w�������i5�ލu�96se����4�p�tND�jt��Tw����p'�*���2w���ϳ�����n�m��O1_�ۮg���n�	ޢ,i�:|�wi�PgJ�2�W��z�Y���U�S��?�l����a��"�N�9l�S�������R�� V*?w�:�=|ƃ��H�=�Iy֪vyab*���¹��Y����Qhc����=6et,.J4�J}ȳ�*�[�]g2�k��aB��^˱,�[>���c��#oD-6��c[�����L�П$h+v1�����$�Z ^'H�yU*�s<��;��)ļ7HD8�-���<{���7�O!�M�-ZxW�ԁ��î��ù����8�Ɩ�tv	N�"�K�ԫ//��u<��W;{+*F@i�7���28��>戭c
��jbS�^>�;*y���o�����L/�-쾻�Qd�D�f�'ʕ	�2��$s؞�*K�`/��p������}�
�W��v�Y�>��rT�y�r�5��$'@H�ڃ0��^�ͺM���̖�3&C���9D(ɠ3,8���cj����bPn\F����/��wd;Ȭ�燖N�]R�vҴ[{�I9��Y�E"G����5�iT�g=b���h�R�[�ӆS��U07V�ۃ2=��'0ފ�(��H��^���CV1dQ[ew)��4��-�V.9O3Ll�4�=I�6�/�����lj�����%�ڦ��J�}�{� ��A��&~�熁ɸ�S�wn_��)���
�;�+��:/B���+R	���O?-Owں���ø���F.(Z�&��_��q<{�f�����xD%��*\聣)��֩�����~�v'�^\j�V�p��Z�ҩ�g����N_m(���9Zce�+R�MZn��Z�{U��b��N�r)����`�
�̣!G�*��,�lH�os9�x�@���~�W���\��S)�W_n��y]��<n�%(>�6�lv�2���ДY��TK5��!�����Ɋ�s�S��%�C��[~��S������[�Q��,;A�j�'K��hʯT������ �]�����c����d_��N5[�,lC鈣Vs���Z��Zġ	�V�ih����.?:ƨ�=M+|ps�e�rq�Ʉ;�ki�;��c�lt2m��n
5�GD�T@��D4��:�.��D���j훷�o��������]��{-�~��@K��!$��"3��C�-&(�}9�P��C-�:�ɪ<�6�xb�43g����ږm�X$M%u��?���^~�X�u��&���Tfylx]�|DטRY��¨�pm�<�X�a�AG4ovP}�urH��Fp�.o԰���+)5:���X�����B��9u�/���3z�:��*k&�}��J:2SW�{.7��o�x�g��Dp�u}������iTP��W��9�J��в�5au���MR��[�H�C��Knr#D�x&�,��9ܷj�'jz��fus?4|b!R�z��n�����"�J��A7]�."2;ȋ���B�9�E�vM*���N�,�s>�5���dU���Ѿ�\m'��mP��,��Y�H��13s�4�������c'*�J�^:����:kl���d�y���,,j��`@[Xx�秕5xa���!��`�gU�}�ȗ�0�PP�Wl
�s�^�ao,&���`� �v�Y5[�9 ��EFI��a�}��P���֞*͚�n � ���vUXHWy�Wg����6&k��W=!i~%Ã���qz�8PY�,r��F���潯U�ГW���^E/'��
�2����%ղ'/�J*�襼N�R#�	���^U�K}���;^N�u�W��n�و��y�aJ�!��v0���v�X�T�����!_�e�^�<��y~q��B�.�^�wj��Ӫr��(�x�&zb�կ��ǭ�6k�o��������I�+�CH����pc���
�vx묰[xI���v<�	lڈ�+�Wn^5}�6[��4k/�	i�V���FV�O����WԸ��.���:��LߝB�B���p�+�<  �u��6�U������+C�V���VN��t���T��������~C��9-j8X+^����g-�x�WlF=Jd�����hu�7���A��\���-z#���D�����8����B��r���������Mk>��
i'�Q����`��l��m��﷎���){qc�s�5>�@[�<0_t�]L�_M�#�L�geU]j��~��+ĶSQ>�����-�貮��7]M��DFÒ�t±B؆Z�'mꚤ���ێh�����F" ��`؂�����wO�rt��3�8��;X{�p�z\u���T�sx�w��]bD�u�ڥ@Wx�;(b�3A�{�<�P�Q�W�C���e1j����M�Z� ��8�����E*�A�åʼc���3���vK�^{�T��ֲ�3OD�4��6܁��F���xb(q�%1�W�:%�]cKdU�y��)]�T��Y,c{�6��'SKr���Y�E�]=�?k�=��Wc^��e�:�>�ܑ�d@5|ִ�[�N�f=��V�� ��XU\�ʐKi�����3:�m�M�C5�Tk��p0�*����C�w4��}���צm<��@�1�ŇY�&��3�٧)Zu'I���� #tfbͭ����/��� ��릏 �Q]���������v9K�XsW��ϼ�j��o)�k=r:�g1���/�kf�{�VFP���s�2�/��s��]��Ke�b���K�Ӊ�՟���x]�pz�Ҋ����=Jo�ڙM¸�%s1���.�
��X��q�Siijz�߇�n{�uz]RVjf��n�R]&���Ź�)uA�jK?W�����g��~Q�o�Mj���#�q^��C�N�]��.�Uk[��x�z���
s�.��ձ%6nQ�f��M;�%�,��y��[T��R�io/k/[A����+��խ��s���뽘�����`эP�Ϭu�jV΂���[c[A����v�u�-�wؔ����EB���,HH������e��J�>�\7�!�R�~G�ec��v�:��T�#
{��a-����?AӜ�Ƽ�*���"Il&c�$�<��AA�%�u�s=�>s�m&d��7b����-������%:�2-v1��LK��)M�Ƭ�G����W��=1ۇ�p��9B~mq=O�ZH�S峚=��i��ZJ<k�^Y���#Hh{9��3�Sս�?xp�z�K�Onʯ�0�M�\hM�Ժf��)�L.�#`�}5�Z��PJ�bU0�aTfmf���5p�C��+�fĪFx���z6ÜoL���U֬�]
w%K����K�:�M{�p���ؔ�r���gh�.f�A����q�/��Y�k��]��R��<c]�9<�F�EBc9ٗ[��[�a���^��FnrK9��9�Z�w�����U��@�T�L�����o��s��5�ܫ>�iv�)��6��^�E}��B���9�:�=o�)��~�{��{]��J�.����T�_�_|���)(�t�8U�1��Xs<�6�G*ݱ�:�U��r��*�(�9d�u|&��f�X�x=��&�tP/��t�\�ݰ��u��q݁�.���ӤR�]IpuT�����k!��b�����|��S�ՠ���׭�q+M��w��y[W���R���aW�R.��8�b"j�
b��=.�'�d�ű�=A}֋�s}~��]3���m�B�}���i�B�.�>a�Ͷ++�>k� s�����HÜn��ޗ}ћ{H����5;� &��/fr�U����^u:�'Q�\B����$��@��y-���m�I�YlIW��o�˙ٹ�p�-��y�0�I=�uuM4���,�|X��K:�V�Yl>�S�y<A�,����R����wEiu��mue�Xr�`��d�t���9����?Q^>6��Baw��1ݑ�2�mཡݢ;ByΎ��`2�-}�[J�;׹��b�mƺ^~.��U�v���t�Ff�nD�btjb&�NoX�淣(ri_���`C���E�0�VE`��9f��c�=:_��TtGj�V����^\�+�s�M�;��5�"$@�����2u�vDʆ2�����rpJy5�ս��}3�y�����v�gwd�4��D����Fr��H�-nz��x2���ն;P$:�[~ck3�z�Q��g�ī���hF�yT5�ㅮk}/2&��^Lr!���[H��Y��V��������K��^J�zϮ�05����Q����/xy�6�fSYǢ�OkYp<�|w[]���&��t�!>�v�c]��`�U8[�p��^s�&p�y���fw���t�o")+��j)tTf�;4qGt����I�Z�ꭙQ_=n�{V�s��Xֱ�eX޸c��Eۣ�S��h�/��[��&!�0�`K�D����$V>h�q��汪��}�*�����f�X���t`�m0#�צ�*%���.�-7�k�k��5�|�>��,g��Ϲ���.�J;(r �P�=Bu�F���z�gNJ��VYʛV�nes����[���Vv�؍�sUI}^�@����o��$�Z���j�z�K-���y�*��aS���}�	=�yUV61�%>�KP}�����'F�/������i�6��R�t��=�e�i�5k�oT�a��뮨jV�)��=k�k��}^n���n�V�H�U}}���qA�[�B9u�Ե��}�=
�n7�-��%U�Bh@�i����X���<X����@���z���ތ�ɥa���:��r���U��:$�
oNڜ�6_��]����QF�a����ڲl$5�B�aX����NR�����,
YU�g�d���������+*�����f#���Cd	>�	V7X瘕k��TO',"�T��׽r�K����m��=��}{)���*>�x(�F��S/�۰;�6��F�{~�-,imН��f1�nN�ިLC����*:Q̓΀��+\Ծɬ�ٚ�&�Dn=��͕�O� �T�Ӊ��֢��1ܣf-mC�}/�M!�-֬�F�f�U9�^�����~IԬa�؍�s�tb���'3dU�b�k��3)<��c=��O_gs����){~ZÛr�k{[+�jq/����;h�<'����)���iN��/g����E�Pecdޮd#;����}��o�ک���5�rËG�{�����[;]b��t'���Ѿ�._�k�k���4)�&|8�XsD��(>g�&&��nq��3����ڔXT�ߥv�y�^���v�\���=B��@��/h����V�z�L>Zᅸ���M�R���Nu�dM�w���7A�x_33]��O?�U#kL*'�b�	9 �Ϸ3++NR�����O0�j�nV�j�dٯr�_����.h�>�=i�'�f�2�9Ɛf�#��m�_P
�4��Ð޹�oqޑ�/w�l[7���jhF��\,��;������l�
֞n�{Q�B?x_U��<�9�"/>����ʯbT��[�k/������]9�������u�؊wq��k�=���R+�����ؚCg�����Lj�j�_�gu�C�/oI@��cw+s�O��}�]�ٚ��3]��J���V��Q�^��(	t���w���[!�P��w�ї��q�;��^�:x黍�L3z�˄�c�L�0���6#��W����!�ZN�U��܎͋����}�چ�b�g�;Py�޻;�\ŭ9@�mb,�q���<�w[[�ݎ_�'ᱎ���UZ��ܣbR��<in	^��z��psU���_-�x�ͪ����b�MOfS�Z����1�K+އj��VR�z�o˵q��{g�̐E���=�.�|�
Z���]��q����[Ε��7S^�ݹ�c �e���X�}��UКg4+fD�9Q���2�?l�n�ϑ���]�zN˕�����.Wջ�.^gM���V^�y}H�)�#du�nJ��i$����y&�|����Ej�8$�dǕ,p�;:�Z�#ܺ�a҃5�V�:���N�]Eq�|FgǶ�z��`�Uw1S8�n�:*c}[2UB���umȎ�����wO!�n{�oM�{��h��_+�2��;wYB �v*ax�A:�.��i��w	�8��o.*�]��D%�"�ru=�Xu0��hלYͿ���R�JZ�1�Zf���
�ͬX1�\�a[IYi1(�c�;�v��HЍ�iaV8f���)V]�k�yF��sc&����t�wKw�����{�����VD��.S7�c0#�E�thnK�)l# H�[ #%X(�b_gT�ȵq���4@�ư���AȽ�܂<�ݣO`m�I�&��+n�[���.�S]��e�����x��S������02��ג���������7~����P|�1[��I��G]}X�P���H
(�X�xZv�nk;{lV4l슷���yN�j�F��pN#S@���7VW:���ɋ\w�k&^�Hl���J�͖�״&����n]o=i�Yr�Č̌���w����ڄ�^R��gNQ9w�.���ʭ��v�v�P�JӰ���3���#�G�_c<TK/��To��ggd���̫�0�M+�4\�6�wBaV"�sM�\��vE�]2m�n����af��:䀍g��O2�����ӮJ�Fe7��_eᙌ�s��%kL�ۤ<�&�SS�֞lCv2VV��F2�Pѻ؈�(rA�V:�$m�f�	;�!��p��/��B�f�pЇ6i��/{�{��dH_�϶��hrO�v$k^����xh1�p�] ����G�t�w��JoqdXRss*��P4�V*1���Vb����t�P�m��9k����G0j�d�mr�]3(S�X=���H74}�P{��.���袲�Η����w������3%�Kc�������8�3�u�.�7R�(N��@ˍV��k.�{#��#k���X�W�խ�lMt7���z���!x�؁.>j�޶�`�ʇ�YD�pm��c���kT6��<�S�=�K�u��W�@������	��-�ҍЫ�)��"u�ī�quv���Y ����z��x�s�x5�mk��5����a4w�J���N��-ڥ-v���N��(oZ��}�|����:�-��4ݺ�䝙
Nu��#��ac/f��O �lԥ���L��"���(�h&uh�u��Z(
�`��4
��`<��,�@Jn]p�[�W}�#!���X��6E��u�cܵșIK*38�zz�H����"$�����E�`x���J�[]�˻dAN����y�J�ӊ�ހn�R&��K;7�} ����TX��m&�h�E�j5h�F��h�MqqƸ7�9q����"S���s�k��Ŋ�TV5E�+qI�XōRZ�m�I�#`�-�5DZB\kq��FM���L��5��h��h,UP�T-s�܅��W���۽����8�P�t9+ �s;�W��۸��w&<r�d�L��9sSJ�s�hU���I��������G��>����Jg+1�g��mc�SF�أ2��9�fE<�36�8ħ�x�^�nz)�BEc�je��3;[/�դd�'Gx{-�5��+� �Q�:l�q�H�]����:[M��y׶sg�HU+�P����ɂ�j`�<w=����k!��˛�M����p������^�:%�{�p���
�	{^��z�k�z[�l7qZ��2_�m�9�b���Y\��F~S��v�l�W�+zrd� 6���Ra�|�d:�C��g</.�&pn�W��[`9��*�P>��.�8�b��Ԛ��֣NfVR��󕵫��m<���+P�w���7����*(򾧖��J�#R��Ե�z�
���!�q�%�H�q&�/}0�4���r��pϖz������˩oFP�ҿC�å���E2Q�뷗c�
�q�\{$z�;\�CE�F�z��;Vxpu�n=�7�eN�Tz��0(2zWy��]��6Z4��t2��`
ឬ2yV�]��u�Z��P.U��^7(��WL|P����mw;�#'z�1�2%�9�9��T����1�T�A�&�r�ѕ��/�����Ο��{FD6焭��o:[ќ�� ��z+�6fr�1[ّ�v�G6���6$utt��=�mO�c��Mյ���9%׹�Ʉ�g,y�̽ŉ>����S�����.u���{~9A��v{�MM�M��"0n=P[��T�:�N��S��U��yk�	��U�:J��	��7����k�*N���_ڷ|��aռ���U4��)iQ���my����L�K��FZ�6��{#/ݪEc�je�X���V��{{,��B�y��VFӫ�}(*%1����)����x_>�Ŧ� u��$��VYS��]��<�YQ�8�W�;�.d��1�aNP��^��Y[p�`S|���Z������yv��hPݓ�`�%�m ��>u��j��J��x.�[q���Xm��:y;��y���������υs�����hT���VFS>��/y"�"� ���x݈��I���w�/���7;'0.w(�*B����t�S0��Sз��{Cot��kU����'\8u����u����E#IP�/�a���j�����i�q-�C�ou��2���Vh]ڿ ����I˩�W�H��6��1��񅭧�⨘���m�쪨��sM%3���������ҥ�^R�_6�y��FPn�4*��]��%ຜ�Ɏ�b�[ CN*9�غ�Z�k�ސ�F�������2M��J�V�g�k�̩��W�W�W=�j�M��i
*ea������n;��X;.O!�*�_A}�C�ed^F�{w�4��-��]�ԧ6N�U��Ka]�͉T�}��0wΆE������["rR��z��Z�K;uBa���9����ؕ�B�ኇc�p�N
eO�ԭu��2X�r�VNe�+I'SAci�7���vbd�/�,Ce�U��MS� ���fº�m=}��j����{~ZÛr�i&��ooe�wk�;J�����P��SnGJ����N�k����{X�2>�ǽ~��ͫSK�-���i˵̮�/r�A���y7�57)�n �d5��R��m7ۡ��kyQ�Ռ	������;��+sh@��u	]���Ҝ7�z�;��+V��J�Z�:���>v��d@:c����C|&�g_,T��4���������Pd|}C|�<��_��'�J��F����Ѽ�N�{�ˈJ�\���ƞ�����}־�����z���>��h�8<.q���>[ۥ�>�{xb�8�p����Ԣ�%��+�l'��{g*�n��yϘ�jo��%O+�����L�{(5Ѳ�Cq�bo/ɷ���
s��y=�"��S�Y�
҈�`�L�I}^�eV%JƖ����{�k]�&��lj��o�wp�Rt���͈"8[�;�����*Erw��kY�;R����;W��y�w,vn宴���������=�w�O�/�F8����wh=��w3�����q�Bی.VP���a-�����J5�·n's��H����]�x�����m�Cl�tʈY���:YΟ*��5��o1�z�z��\�wOf��&����b��݉�T��(�z�W ��������qY��|��˱�t���,F���/�\"�-����vS�mן�B��1�/�z{)u:���V&��w�>p�P�:dփ) 9u��x�I���ɂ+�p��5ں�R�(m��<�1�f��kq�r���@��2��z���!�yɯe���˔HK\�N��;F��ӹ7�D㝭��M(�!�[��:�\���<�k��k��ک���p�e{_�/r!�Pyf��.����^Tb�*���y%���Ne��k�`���(A��X.��
k��kw85��/g�w��o+�y�ߩ�o��z�r��o���ı���!�qLb�B�5CfP<n��������N�2�k�s�k�n2�X�|�)�9Z�S����VdQv*� �L���88;�����79Q)u�ċ��C��q�Ζכ���m��u,��UR�����P�%:���uO��w��F���o.opm��X}��xI,��N+I�F��Cߵݻ�j�e�-�&�gh��С�ժ��r�fo���t��n,|�����U
V�l����$�B܍W�����c�5��u������)�0���ӪҬ8;�Hd���;�6t�9��Ef��}{+.��mz
c��:>ز"+1ḩƲzμZ�c��n�a;,���%1����������	1&��&�=����n=�\�ݚ}I�ܳ�A��s|Fs��%��)�ljP���[nq�P��B��(N�u���ڧ��Q�;�;�@t���I奍v�{��\�I\T)��1�M��8��fS�u���U0"���;��Ե�o��;oq�ؠ-���&#/�܎=��f��.�|M+��qv��Nr˩˺�ġW٥�&�h����ԣ�8�>++�|5��綬P���涓��r�\綡���Cܤ-���	c���Uφ�9`���,�]�Os�`i�0��-����z�My��i65�7#|Eζ����ugx�˧b�j����G��*�Œ���6��:���4���V�:�D��r��p�gNtʗ���N!�(�bZ���5�ɦ���Xunb��fh��`c�wRif�e0Y��ݪǭ\�.���+#/��c�aL�����SG�~G��;��;bT�]��Te�pv�þ�1q�3����N�9ו|��m�:N��.�s���/9�t2��5l�H|�pju:�����8:�VDܕ��7�,=������畁'�o4��5��c��b�8��1�_}\��C�c�֋��r3(������q�4_>�-73	%���w�Ue��;�u�{՗>��
����N �b]ƪ���=����L:��wڕ��{aV��Oga���0uP����K�3/&�Bbm
z�j�Q^�	e��_�<�z��n�[����w��=��:>T~�8�w�7^��\�;���a��am6�ڜU����Z֔��Z�U�{�.b"�6�p���T5+gT���mn0��e��V;\�����Y˩�b*7��ܢ�s�M��=���}�����h�b�3�]�ۉ۾��ĪeD.�h�}�{W=�j�M��U�}���a��p�*�|�n�[��i�=Ƞ���v�yR:auz݊`E�=���������=j��4�C^�j��Jz��y�m�ɏDn��]^'x�)��IwY �S%@�r��|��Q���>�F�Z�N2߇|�i�tu�v=��4�,�[[ڥ���
8�5$����WW�-�&�u���I��k��t���u�ox<:u7/����qZ��|��Ptơ���u}��Q�d¥(���.z��=�����8m�|��dJ�([*Q���U�n��R����e�Y5������j��0�ߩ��i�q��;9�i7i��H��d�~���m}h��R�~�Nz^���S��˕��!���)��e�a���v69��-��T���[cu:���CȎ���j'vVơ-�����C����T7�\n�z��?{�n}X�3"vs��×2騕��}��䡺�ƻ�����5i
u�}��Ӱd��u	���n������D�[q�_.�8�T�ܮݿ���;ש�t��j��F)��'52�t'�hm0���W���\������{js����(`���.�ɸ���>����HAj�cKy`c�{�Ǿ��q���R��ӹw�o0�G�+X��!lF�@�#	>�)J�ry^��w
n^Xޛ��R�k՘�/f� �쨼�;������2��Ug���un��R�R{o�=�2�@<�9��X�:+�,beko7�5kκ�8�ujщ�EgF��+��)��H�>gr�e�О�q� �����kH��x�a��p��Nq��圶��vT%�� �c�$Gv׃�Oq���zu�0���z���{�� �3h[q��[
{��fئk��9|\=�@�;�];[V��b�e��3z�}�O���]���Q2����Q������rތ�ɤи+����h�q@N�Q�����d'S�D]��{Tԭɯf��2��)���!��Ec��9�7��[����%�d?Utf�砧B6�nNzy�׳���z�6�y�=9=���~���gVo��K����H�>kj��̯e-scuk�r�� ��˷x���y�J����5m��yT5�q�"�Tf"��]ͷ
+s�7e�{eE<mн�v9K���9�s�UVn�Fe��n7/ro�N�Ng�a������2�ڄ����3��N}�5���7���ޣ�pܼ����Y���31�Jؼ�g� G*5�-��3uo��q�x�3Ru�C���9�X���¾'s.��ލ�������H ����|�A�#�^.�f��,���	"W�z�\�V%݊q��J��-w�ֳ�p�����k;f�R��:�+���!ˏۇ8�B�toK��j���|���UתEV���œtq��.Tu�.�Aޠ%�l���9-�\޾�w�.�UU��e���nun���u��[�y��a�J ��m�=�ɫ�}�F�US��Ya���-=�)ί.��V�l����'�j0�M����p~ͮ�o�c֟��{,ke�i��lL%��	���P��i�
�3���8w�}t]*[4��ֻ=�g<�z�7qP�H�Yh���z��t;�[�D-�#�]��Ե��o�:}���P��a��1��^e�������<X�>����Z�r�z2�&�u��ؔ��o�{�W��\���ݫ)�4�.+�6�}5+s/�7�Us��/`J���T�ק5�g�����v�>T�z��y�u��%���7����_,�WT���TRʻ��!W���a�osA���N5r�|.� +1�Ɖ�1�u���nu���|x��WxE��i���ǊB��G�� /Z���v��y��0Tۉ�۬G�	�C�O��w�9�������* �v;�|�.�t;o��S����=]����(^��*����;�&1O�|�q������I廣�īܮ��$*$�5o�J�r�d2v5������f�׊v(�u�77�K9y��m�#�ü�.{�Е�_hȕ�9���c��h��(��;vl�ARy8�f�H�ڹ�Uo���C����m�_0 vo-�5o_T]<JI-7�`޷��,{�[us;���fh˶]An�gj�Jm���-�a����2�'��=V�Gw�p�xp	1��g<����A_wf��uly� �pԴ�C�K��l
gFD��ej5��T�5���T �[mw΄R�b�K�T#엀=8� �N�����F���J���/;7$4�5�_V�v9��t,(	��T���M��-v\X�ҳwQ����*Tɕ��ƻ��� �#��*gV�h����@NhάW�ܨ,�t�{Y��\A ���6=��!*���C0Q��TˤZ	b/�-��D�E�Y9e^D��|�'B���:���Z�.�p�}�Oe�T�ۄu�8NF:�솤�y[����'�[S�q�i�f�U����X�%\6�F�f�wӦ�բ'�P�R�	{R��&�z��X�^��Lf��C�ơ.�x^3|����ٜ%3�Ď9r�w+K����@�a���;���xbޝ]��zJ\�g[���n���ƫ|�a+�e]'hYV!y�����3r=��6��s��i����]�]����3��BSti��3�pօ�iAwzn'����l��M�Hh�E���s��Ҩ��4�p�,gX��'VšÅG�5�ɰ�6�͚��m�U��Mѻ{y�7
������w����MdVM�RWB_.5�l��v9�e0�S������,�B�rLV�G�3��.V4���+]���R���u��$�f)��H��gf�@��8gRl��Wt���h��K}]O�{	[+^�؃M3�9��IUɄFY� ��容,Ŧz��1����LXH�H�K�qA��%T"�l0Ol8\C�g�.�7R㬺����oCug:���#���+nV�ݜ3+�ݡ���iD�&��ef_�>`�H����n�'r�lWK_n܇X]Q�j	f���N�d��\S���]3X���RT�w��R]c��鵕�1np��E����X�be;.��������Ld�C��U��W,!B�,ѳ��)�ɷ)͔ev��xn`N!'��� Pw�=ط ���|���DI�ԌH��!�ԥ��}��X�R_X[������t���Hn��(r�z�Q���5���xy�{�V=�mm*}�٥G��������x��c�71��z�he�}���]�\o���(P��>�
���q���AV6�W��F�AQkE��rQb6�V��mRX�5h�Y��E�����-�Eb��Z+M�qq�\mƣh��3�TX����DXэ��-q�_��@ �����@��.��q�J�/)�ԅ��E�Zue~�X���$�u!��xe�uǍd���+�5%tp5]iFAf�5�Gr�6���r�M�O$�x6ƻؐ5ى�xb�;H�{�A�Jp��'�q�*��ٱ�����ZN��0��lF�<�׆$k�8VH��b��bgx)�.3z{2�������/j������9�u�竳k��s�i=����qG��z���H�j�1�o�D���ڝ���^E���#�ލ��1O���e&�]�H/�Jr�˷*�RXg��8Ɏ�<I^�:A�)��$K��G��Hg�դ-������X:����[�lcޕ���Մ[��5������{˷�{[�G����ݯ�=V��u�[�6��9��jPZǣg�YJ/�W�6�9��.���#Ds9��T�z���jp˃�R^��V���������0��i�9�1Av�L�Ή�5Ρ�O�q(Gs�IK���R�E;�9��x�Q���\H&��b���]�8v�ط����]�"�'��
Uf�'r��[��2�e�%���Jĵ%�;��P.��R�N���o�'��ᐻ�����un�*o&�{n��HB��̧K'K�$
]���o�l��򾋗����7�0/z���1�U�f����T%��K�O��}�b����o;�ubu8�f�'�fд�*]#H��og�w`c����*p��v������'f���'a�ֲ�P��.���.0�lϤM#�Y��[>WK!:s+c�Ζ�er�}C�	�
��qGh<\V��1KتF�|Y�_�gMO,���n�(t�ӆ��ؔ���n-4��ЖlLB��[�b[ɡ������M�9m�sY��L^�U��̌�}=��^T����h��%�y�I�V�N��1�#��O'3s�K�Х��v�ڠ9���o�3	��Զ6�S��B]x��J��Zj�Su���+-�9��6��f�F��fC����8��_���p,t=��e�^�/ ��SМ����Sq�֮��v�םi���v9�g�Ӵz�B0Ӟ���,pծ�V����X��[��;�U��/q�3�x�����i��U���iWB�� 5-���x�E��Nn:���W���|k���~���Ͳ��3����r����}۠𒲍����>�Ʋʡӳ��4��|C}oyK��q�Vv�k��e�h-D�ԵJ���b��]ֺ�Η�u��{�΍��8������f뜅�4i�]��郬���Q��A+�Ռ-�b��<�|�ߞ�z�9��C3��s<e�YtlF�)�r_W��*��R�4���7���N�6��ˋ�:��+���##�q�}�b6A@�*�����T�T���ͭ���8_]����{~���y�m���/����Ij�G?o}2�qx^�{V
i�̻{\���x�`}��n0�K}
G{z@!�<7��7teg]Wj%�t�b5+�/��_u��V�{�o�3�%�4�*ȣ�2%���Hpk,��&g�,E�+�ץ���rT�eM+��õ��%��wNoJ�x�0��N/
;PyW�l^��Jܚ��.Q��4��v"�k�{#��f��9z&�lH]9F��Օ�4'�M�:y�{�w�δ^�뚮Õ�m|g��C����ko.i}�_�ͫV<
n�_���*$�<����#ov�@ѸEbK4��.⥚�YQ�PG�`7���q1;s7O7��jl+u�қlN*#�Q�k2C��0
&�.|T��v*�ޚ�{��h��h�W��!oT'c���"��!�9�����%,��O�՝a']akj��ʠ��ߟ�g�zm��2�\?��ޓ��R��q�7S�{X����c����q�����]չ����3��k�h\��!~��^�[Q=��;P�e�v�^ŎZ���ݰ5gDI�Q���J��w��c2�W>�ʽ79B%8�m������Z���J7�v�c$����~����M��0�
�;+�\��?�m �ư��{�(���n[�o-v�[#Z���6g�j�v�[�1�	/�m T���Q���ಸ�xS�A���떞ڜ�]eU`�Q��� s�<���/|�-99#�=2�,~��ag6�ڜlL,�؎���J���~��j����QרK
����K�Ke�CZ�g���o[���[X{�&j��f�r�*�Y�Ӡ�����yu�c(ض�B+U�>^Qʏ�s3�[˝[wID�3��{�z�֗f��T��m,�6e4Z�Ѧ;:��p:�`�5�~O��ՆD�U��Ư5�k��Ct�|�8p펀���{�wu�1�J�2��\����z�m_��nz9u-}0�wz����966���n6�Cb�"���:}�]"��z�����ɥ4%V�F���}{��7�^�w��^.�Q���lGza�iS��	=�� ��ټ_���yu{�,6���v���(�A�Q�\�9�E�rm��)�u��_�����}S\���6ƻFƺ1|�dE��c�ۈ)n��s.Y�ܚ��o7/+V�j�Vu+SͱC�V�0n�*��=�t�xz�����m�79-����ڽ�v)z��4�,tN�J��5��f�ҥ��;J��X�ߢ�Tf*o�Y��=���=��f�J�9�~8;���Y�����{�A�~�����˶���D�(M8�u7��uۦ��uY��3�F:�ͭ���h�8��U��,��Y�T�<�L��.��ۑ{$I��(=���Z9:�yHvd�K��V)���o>�5Sy�bm��]ҷ)
�a��EL��xxs�G��wC'�ɳ(��:au�{ࢩK]��R	ml�TU�Mv�sm������f��tZ���_��ܝg1��Ju������ɾW��!Z�$:����r�0��l'��v�N;��\�����G����۹cBqF��N�H5q���)E�J�ͷ���
s�ݰ�=t�|ƙ����e��{Ӱ~�� AJ���;L�
�+��X����{��Suf�6��;ag��7|c���0�v!ϊ#	v�ꆥl�����b+T��fVuSSn��;�;��2��7qP�/oH(�I�K���)}'®��f^�Y�;K%lfƱ����ꖩ��J�5���́!wl]F%�)h�ouu�kl�̪y�l&�f������o�����9j��!b�������s�*\�,��-�����C��+fąHϸ��GR�/��u����£R*����}�C9:r�M�Miølc�o�s#gv�[\�wd��"�G\��̰'�Mf-�����x,a���ݹ��{u��}6�I!�<���%�{ |�v�euة���:�q��rr�|3R�,�8fP�;��>A� �V�~u�l��ܝ��O!u�{.��%,.o^탐����خh��sN�
Ӹ�����Vh��S��lp�*vƻx�a�<Ov�v'�J~ҷ̂��Y�m��s�o�����mݱ6jG
�O�X������
h[�v�o�}f:���wΔ����0S��Ip��t����l.�,n֦K���بcw��7�]�
r=�~�M����0cj�� g�u3ҵ�%��5��ϔ�n0:����w�4o�Fcӱ�1�k�6�*�93W.-����_.���������"O�����J��uEB��k�(\��tk�U�T%�W��J�e���P���y�|H�^ǆ�^e���I>���C�v�	�V'nM��C�j�`io,GR���]��>Cg�-[���w.�%��Vr��Kb7@��a'�tu\�<�%aǾ�Ru"�ħ/S��߆0����s�ߢ�J����w@RD�G.�9�*U��,��t��S��e�ƻFm�\�B*���s����a�`�.�B��x<��`��oi5��u��s�kL��-���yY���)%^.����^�YQ][�*�q�ۑ�8�,��W�.H{{gq�vM$_)
�J]�����	����e��źw7�U��$��^:o��ʍΤ�M�nw6�x9��w��Ok��۰��a�׭�G �.��<%o38(����ɝ��^̟F��of�k� G$���ܚW�;�G�+8�6��;r�9y!��gO�-W�b��[��ς�A.s:t���J�z�'�R�];��6$*Q�7< �Q�%nI�s|�}�N]��:1ܹ����x�F`�<�*����lk�g(k�9GH�[B��̬�X����C(Ouv���PԮ\cyQ���S���5�hF�o*�����]}���'�:�K*�.�	F��KYBulm���z��߹��X�]F׆<�4k��J��tUn��So��a��ʒ�|�畣VR>�=��fs���{���/�:��wqg��h�gev�Ҋ�]��}Wˣ}���3�ֈ-u���uk��P�'�����6�A�o�-�qϬ9��:��߫������mڙ��`�z}t�_VD�G��4�F��׽�{ش������ÈeSU"���Hu�/%>�%��Q�Ĳ�ѕ:A�bu�f4��������b �ōs�T������vT�3:1�UfZ{َ���|`���Nw؜5� ����j[��|�9�!��;^��۞5a�M�E�ff0��>Y+��i�J�����a���}bZ{~
s�u�t�G��mMܠ�罼���}aq�mQu���4ooXk,ci��n�lx�&�x�F`�\�:��UCu���t-�R�5�j�3���~��z�uQ\���=n*2@�k���(��~�]K_Mx��p�����DT���\��N�N��C�q��f��#��a��;7���s��9k��a	�̐ҏ�۳��m��dSol�0��+�ѰGzf�4�l�>�B�=�;�DO}T�S\�7�סۇa(��v����E�_�k|�RA�;=����C��T�$�kͱ�ѱ#]���6r+Ru��^�읞�r��Eoy�o���$�U���b6��K�{<�٥Y��f<��n�3�u�]݋�5;j��x�b�����-S��r�5 xc�\��)��H=�h�vi˥�u\�uց�� �G��Ž�����n��9�Ǖ�8�Ρ�W�l��	\xm�L�_A�����ӸC�M�gB�[�S���Z���ک��Rw^����v趪�*��C�k��h^ջ�/o�XrFC�ǣ�׷��3���z�����Z�F�eٝ�Z]���j�{K��,����KGt�MY]P�^�mC��䱪;@c�������8ח*Ê���\�ą�FI�˶gy�C�Z�̦��}a��c��KH[=i_m[���{}��:o�<��S7+\�F1�	���ŇM��Wn���o����Zn��:�w�eL�v�����V#g�YJ/�Wͷ�/��S�E�ژ�%��Q���Q35��<�I��e*R��[����0��Ǯ�
}X�S�ݢ�E^�0��P�lGH(|�	)u����*[4Ry����ʰڪ��]sj�o'�am]M�v"�J����\%ݒ��h��w����y��B�'f僼��B�ہ1�m�|���~�ThW��]U2]��`�$���-�W�9,ݾ�Y�*E�T*qZ�Te���Xs*u�զը�Yq����rt�_5�2�)�lH����dL��ӽ�zc{��
�gM�7׭��E�N�:WL�'s|�c{�_��\��v]G����.�c��)r�V�_F�n�-\z�
���s�c���xw�[�Z�ˡˊJw>s�cݵט�TU�uN�Ț��P��=g,ȗ���ђ��7��#����pSa�N���!s�0�<i��xJٗ0P�X���ڴ����P��(vv��t*�^��]j�m��V�tȬ�޺U�2��L�J���&]5�z�v��.���P-��'Pu2V8{;����m��}���7�-ɺ�L����p�Ԥ�Z�ܢ��ԩ�]8!�(�<�I�Z��ZƗd���^���[tɰ�R�s���U��+���׶�d��'AB�a(�A]�A��i��u
-7�j���l�pn����d�[�m�kC[JS^��^&��C�1�ő�B�3F&�Mb�a��&
���Vήwe�Ę�tE̡H��<�$�!���Q��|ì#K�
�Ki��.�k[t	�m�=u��]7�;�nt��r��Ķ�j�焢P��we�`���坱9�h��t�&���W	��']P�0��Zo�������O�lr�]��8��Q�5j�(�egk�uo4"�zM�����:uw������N*g�G �|{R'1t�^cl��6o3VS}���/�WW.��/3���ؙYK�5 ��k%�Z3�C��yn�3��hEW	Gdm*ˢks!
إAn����iW�*M��2òA���;]ھ�X	F�/[��y���]Xv�[Ηc�:ܬ��7�N]J��5��_B�����s|�p��zS�EY�ʉѲ�r�:�:Wq�}�q�a�����F������
܋D�+E_�QGu`�GSHvN���Õ���]�B�aǗ�KPa�g-����ε]N���и�OST�-zƏ>�2�ҡ�h���w%�l�����lǐ0Y}Ҥ��{���<CDY�z��=K�ؕ�VDk�Bʹ�K����_U�m:��}圪�_>���s��X:�z묢�+{�\���Q7�;\]{ԍ����a"�4���a!��ݓ7z��h#G$��2����}9d�'e��J��W;����AW1�B��j��/{4gd��ͧ��l�gb�*þ�i�O�����M��e� ��,��o
������:�y)��\�I+�2�
]�u[��������\� .�6�t�k���v�E͵��Z��9=p�Zn�L:nR*�p3�f��O�+X�j�;�V����MT3�F<�o��r�-D#h@�a��2gK���3�+���������NH�w@��mfl�4��3B���k[A�H�+�K5�w�;�cIj�u��e_n'kh��c�*��u�xw�߾��Dh����F�+��[��8�ne9�G9ˋ���qp�qE	n6�)�s��X7�W8�.98�n1�0	cHF�q�C��.s���QQI0шK���j�g9���9��$qq"J1���N.s�\Ÿ�h�2h ��.+�58�6��
��k��D�qq!ɸّ�����_��bA��{hMOb�P
j�u-g3Q�()fr'�O{��Y�wk'si�aq�[���l'���e��q�ЎN9��r+�oj�i���SJٽk!�Ey�r�.���.0�i���68D��.�"�f�f����� ��9sK��C����5����%-�&J���Y�]^�2��Tm��SR�&�rt�C�����8w�lc��q*rX1��/M^�Ζ���ݺ�*���#�O,Թ�~>�nG>��`�Lս}�j�6��)�ቄfG���~��c�Fmg�ߩo?I9\�sl_\N�>յ<�d��?bU���n�f��<�ߟ�e�M������8J�]ZO33G%�2TS�����2����f����߷�ڞ��{��o�D��OQ��V6�Z��g!9o��2��u��'Zߌ9��?�̵��PJ�T����!�Gk�79Q(>���.�:�XT�߂����[�!E����kvnN^YL
Q�^.��\��Z�-�b���@�;.�ӜM䵂.,�f3�A<���6P�Y��ۘF%
k��v'�j��wI��k�[\�ܨm,�.�A���b�9��K/�}�yⴓ�6�Zw��#�%	��ev�꘴����t�1cGw� �x��WL�$�*�s�.�o��)�[�n5vg��oX���F�<�*����*��K��&oTU�����n�꧕�J���\����W
B؍���P����A�lΫ��t����֚`muM{[{z�[�<w���7b*���C��3fk:�j���ӝ�0&�l�a���e�ƻ<�3k��ar��B
���,;tG+�j*ۅ^�~"�-���寶�~f��7�3�wӶ�}�Y�p���:X�#}�1�O-����-���V!���b/v�DlF9�[����c�`��(���#`��Jۜ��E�9MZR1UX�5:��(�ܓ�����~F9F�N�n|V�ײyb���^s�%��vq����6�h,N&�m�j�׆'�p��ӛ�ܵK�8?t�w�H�eK���Y�o���XsVЍ��^�q����ng�ܺL�M�����H��y�(�6�qۈ؎B�mڨp;<�ʮ�4fԨ�Ѳ�k��eo��U�WV�x��d�тơ�	n�V�Ⱦ]�@�]�k�r��W�� �vxU���Y�b�[�cܔ7��y�$;o*-H���������}��K�Y������`s��X��k���fFs=��c�������)��̢��c��������}<~��;3�Mo�)�=ۚ�����Rx|��ZAک�KG�N߰�ڹN:�b/�F?T0z��C�tf���>I-b����9� ��}qoÎX�,���<���P�7k�J��B�դ[R�s{����ݾx���؍�����wK�T�0���SN�XS��c�=(�;]-��j�M�r�r���V��n�U��2'Vi�*� �=E��b+6���;Q�:��&��_���Ol)�{�_&r�G���{z��gكû��-J��)嵭v{X΢s#���nD�8Y�A��6�w_��J��!P��G>�s����6��%�I�l8d~ɳ����Ivd;N6��5�aO�yt�q	l_�o�N�vðzB��u��}<v5�5�$"�޷v�A��ل�_u��+�<���=1�=��Bёm�E�E=`]�(��u�R�K-cU�Mg
�
���]k����dN�Up�/Nmw	6����}�^�)<�f`:{������=O��̸�c�^�IޯV��2(�
�4�#�uF�)���0�nf���Ӱ�u�Z��Y�:[ќ��&��vᨡ��t��9�%���q�����d���:�k��w8t�T׹'@6Ƶ5щ�p�"�շ&��W�X�YB�컖�{um.�V����9�b4�q�}�k&�HWN���V��hhqd_��e�=���g�ټ��z][�^:�uMٴK��Lν�*V^�/��ڞ[�H:���;~�K�����]�o'�*-��)Jzj�su��L���i�MI�Ǜ^Uf�\fP*�*��xeW^
�Q�Ǚ��-d�	�qB{;S)�x����+{A��֖�2�Ԩ&���X��2�CqG,��<_����>~�����퍞��t)討gX��v�9���!�L_�{��j�M�;���>�s�zy��]�ļɊ�7^�	��G:����a&w�3J��gX�M���n��<�7���ֳrxG`S]p������Oa"�.�A��~�y�=�{����ihaY�]mvs�yd;���F)�'Y����\�+�4x�I{yv.�UY��ѕː��\uq�.�z�%�8����=ʁ�h�X�V�W���c��f�K���mLw$PW[c����l9�W	lGa@�|�J�a����ˏ�iŚ>�l���tgF۹�O87��-�<���P�{z@(BN*��w��,�"7k:���E̻~��4
}�![���mn2��*!eo٪�p��$��d��D��'��(q�]�>���`���z�C܊�m��oǀ�x.M߲�+��y�Pz��SB^����C�5p�C�v�X�|�݇otGDVo\�����p�?A�Q�%��&��N���}S�8e�̧y[X�j�N���哩<� �]����������A[9�y��̸Zo��Nn�X�t�}v�f�eᷔ\n�U�l-#>��ke��<;NA���Y���i|oE$2S��u��h&�n����m��zwz}] �ߝ��o}b�ɟ^��Kc'�G�N���T̊~7�������c��WS/!��0U�r�������l&����h�J�erxL�K��c�>z��7�jͬAv�S�c���c7:��`��-9��j���O_K�s��}4E��Բ�=˳	��,KyƬ�rD_>� q^����Jة�f�)K�웺��}��)�]6N�F�n=��I���7̭uPs����3�qŜ����K���4�(��dH�q�T�� �S'pj�[�ކ=
�?0s�u���N�n��w�ce_���V(���Q�����XT~�~���ِ����8tu���q�(1�W+@�]$v}��W��J����]����^��V^nSޙӶY=���Fv�]:�7���6�0���"ti��!JG����#ʗ��zw.tv��|�B����1�sĞ5�+�@ʠ���Qb%��z�tV�_�$�u|��u�q�0�x}�2�юᾟDST��V_�H�$�̠$>�NA�7��f�M[��%~��JP���]O�q���U�W�O��!���Cθ[�sX��@6
4�������h^M�3�l�>�vY�. ���3�n�Uķ|0{�;\q��;q��K�F�9��~�3�.�cM���g���<����-�>��2�Z�|8z[V�7��7:�U��Z���a6 �Xj-�R+Ո~ܷq7�J<�'I���u�n���ê��l_��ۂ �Z���9�Q}[P������p�n���s�*�S��n�Q�����=�];�XgF�KnWcr�M�r���Xyp���V�t�a����ظ|��tBw�%��Մԝ׌��Y���\�!-���ӽ�f��7[:�>9s��J&�m$;c�R�W���܅�G���\O�S���n�����)�3��26vH��m:7Eiʿ�n9��}\������۶�Va!Ƽ�F�m��� cBl�t��ёe3gg¥m`���!���7k��؏�����9Zo^T;�.��vKdѸ�������bE�N���A��oٱ)�{���s���+v�WF�-7���zw|ak�tTy�m��7���h<:�d�e�7$ۍV�p=0���e`���a�qʴ��۴�����c����Z�s����ڿG�(~��+Ʀ5�O.�{��/�8lq���Bu�������N��� ���cʩނb uo�,�C�9>���������ӹ{ ����]k�����ڇ�/���N����\f���`����"�g;��u�|�|:�l�>�X�����z����]������S1�4��W�����@�,�C�9d�r�e�?\6{���w�s�!´���$�L�uj%i�~W�]lԸ��]��qLet�Rֺ��]0n#΃/
e���j��׸�#�2�R�!S�:�K�l��-l��)�r�^k���jn]�����E@����`�^�*�g���G��;���{t��DO��/ndl=p�:��|N��y �B|�'���{QgT�}I���M�)���18�Z6��8iλ��׃�`����Y[$�����ǆD��\����'���:�u�G�WM
Ɲ���k�Hg��GnWc�oH,�x/�V�U��p.J<4���&�$Qr�O��u�!Z���*N�z�h��쁽� ��O����f�9v�ݜ⺕B��B"�� %:H�_@��k���e�����Cܲ���z�;�֍'����Л�2T��@���'�J��i~���V{�:Dc���8}�e�k���f�YyX�n��][2�%���$U�t�;�;�����s�Ч9�z�2��Ƕ9u�)�Ĳ�.|�hM��m*:�N���5���zc`�=�T\]1��:yJ{v�ÿGs��7�tb�9'f��r�k�B5���U�yO�7�T�
Ǵd�N?��7`����������C�zwt-c��}�H��I#����]��y5� i���/�yRF��
������[�9�?s�\�T�G����NgO0��7�,��/l��T����pM�й�����syZ��j�^�p�^B�~l�����"?;xd�P��YJP�o��Ӊd����}��:ɔB��Cm7Q_7��#9�; �[/`N�>�[b�j��� +Mgf���S���T� �ӓ��П+\o��)� ���.�[�@W5���;��7���#{ ���l/�u�j�����Ջ����CΪ��T�59]D��<��W>���e��.ex�s�8���Q��l���S��.Kd��\�}pԙL�]G\6�;�Y���~��̟mߘfO��)�]�r3GR�.�'��Ϫ]��9,����ι���g}
��w��#�`�^�Q6�M���V��v�����'���gK2��ڠ��١�
P#}Щn[;�ܩݫَ��N$�6i(������E��?x����A��."�{�������b������y��8/m�*3�j�x�Π�v��.rT5�%��%PC'�A�H�]TK.5חs�9���awk��N����w�a�R��c����R2ۻa��R �Ȓ������#�&`z��t�t���XL�[�-�q3�s��a�7Dz\�2�S �_t��p5���=}���.�q��`U\�,⇣��з���%;H�7��E��-����;�da]��w�^��6�n�iu=�ag���3/�A���)�r8�����˭�=��Ϡ��%}��|�\x�Y�̭O�w�A�jnk�P�U-z8��<�<F���mu�zJ��%&���TP�z�ƍ[H n��r\�}؉�GYW�)\O�]�����w\b���X�_J�X��yV�GS!#Ot���e���p1{�/{��%��5Y��y�w��2~�C�U�Γ�='�!���"������k|5S�������]��y�
��Uׇ�����w|���<�
���j#�� �ZC��K��3��v��G5��M���6�>�k�_���J���<t�遅�����~']c�Ê�G����.�-�;~���[�ub>��V�˅��a�Z�GΥ	�o}b���g����A��ޑ#;{ݗ��5���^�p���N�e��-'O�ݖ��o��/�7���V}���ךm�F|m��]�u��3~���{�Gu<38O88�S�8�d�3��}p�*����u��������`,�{��7߿<7_�H���mN��O�\X�Ma��)^�|���h�cjS<Y��u��.ޣ�n��>O+��eN����0�h��+��W�T^TK�=E�[>�5V�2��V���ԧr!��}�w��S�᰻�#n�I:j"O2L)񕈌���������t�	��R���F�O��e��7�覩�+��p>%T)�I��e��*�N���˰���n!Z�:�g+f���.}��WLA]���ְ&�b���K��}i>Bm=7
)S��X ]r#�4ӭ{�s�����2s���V]Hz9�jbfX�n>3�8��&wf�����IWn|hX�VSQΩ$��ܶ���#\ڡ�[z�s�jH�&��3�^����������Q}�2��/r�Zb@RiQ�W$;��;�9��:N��Te�7���
�r�$���涒;�|�����a�k ⁾��k�Dw�o�w>=I�^��\S��X���*����]��gM���'���*���:�W*Sx����q<��H4�6j��g:��j�#�lgvT'��z����^ҡ�S��t�)�h2�|���$�ޓ{��8,X�l(���\�s�gn-�S
񩡾kxX��ֈ�ӕ�h-ݫ���Ed'���@��r���h.�n뺟��xy�8��k�us�A����+ɹ%s��[���7jT;ʓ'r>���9���^֢��ϩZ�Ge�N�q�>��!��I��B� �l�,��}�{����`7��5���,�hwKN�;jcdjB�h��5р�9tT��yc`\�NK�t��Jj�)Qo-��έΏ-�7�`�:��¬�b��r�I�U�|�bu�Ȧ<�c;�e�{�}VyPv1P&b��O~{7[� }ꉫT%N��mA�Xs�s�.e���Uy9))i��8��S��:�����x�fsY҇��Q�v��cj�D=���L�썜�d@�z�@WT��uiWQ!5�Jг���c�[�n	�K�G,����S���@�uL畁�Vt���(����(�%�_\|���b��1)��Dj��2���q����Vw�;9���#m���7�!=��r��z.�-����ʜz����xN�a��gφ��Lަ/��3�+-��(��9�orZs�؝��#��*:$pX��x]]��Xf�E�ř��s�Q]s����*s'����.�LfA���k.R�gpVt8�r�٩��/���%�+,���e`�P�"ޤ;54�7�6�#�T��qZwd�d��M�5I��v���א�a2�u+����I�����.bWq�q�Mb��� w���h�{y�g�T��YQ+8:�i���;@|�nX�(c�/�k��A_�������h����Q��J��ے�[���C8�H�Ќ�Y�s ����#{ա�
�M�Y:�r�cf��׽K�-��:F�C�M�+ɉ]���<[�j�{��ܔ�W]��A��fVb�˫_!V&<�x1%��ʼ��+��ILX5v���ilT&�ϬW Ev��m܇T����8���W��g^Z"���Z���M	2��؛��3)5�>}��s4�W����/�9�
9�p먻����}ݛ���.+��Nr�ی��5rk�E��M��5��a��ܙ�li�\��4-)�[��9qq�1&4`&ZJ�⦅H�-DI���M\qE2��B��&$�(�a"��r��1h&i6 �@��$!�fRD�H�!$���&D1��Ȅ��)�0�C��!(�BQ24ƈ�h!&K��s��	&"F4"��HJhW_;��^�d�go�or̻�p�+���Nt�u2�E�U�������/k������oo)ۅ�P�
�+�ݓ��1I�*��=`�+��if���gޞp?r���"���>e��Q�z���U���^eL0��|��`�:΋��I�NxQn�xj�Ҵ�~n��(H���ô������<c�D��� k����%�@�oACR�|8z[V��ʇ���-
�����7tBIY��=^��w;��t�\M�%�:LO�ζ����
CM�����wQ���f�)?g^����g:�/�ς%�>a��MB�s=!#�&VӣQZr�o����_�|3�G|�l��*2��tm7\��� cBl�t���N��2����'Mx�K��n��|�J��hS�H�͕��m�mUQ�Y)�F�m���P��y2k�G�Ty@9�vN�:�ӭ
p2|�KÂ�2����ZoU���N�z!k�tn<�@:�z����b�ŝ�Vn��k�����Y��2�;�xp_�\�I�Dn���x�:{���C�g� �!𣉃uo?q	I��+���Wqvl·5Lp��W{j��Af�`9�H���Ǻ�Pl��>AÛ֣̫����;��U:�g.�Y�z��c�Gkː�iQ��������9mL��\\�4#\��]���]@&�`]8gi�BL��Q@�s u��Vv*i�uեw/x-���tS;G>�^n�B�Nْ��h��|9jR��\R����&���i���{�co*c,)d�ِ��?*�*�ė�+��X�6
�;��y-��@�[d9s��P�WO��\;���\Ft䝸�d�˙^4gj;��yn��g��W���K��;����>;.�����/��g�}j�r�-��$�X��OLk߫V����y�7�B��ѷS/f.6�	Sp�Յ����2��9l�P�M{�W{�Z��1�CעNw��3e��H(�qbOO���ʟ/*�W�������t�ޏGW>���(V���2�T�6��M�[sY�;��H�'��A�&(��8��O��訰?�c5R8��ܶ<�/]_W����C_�+��n�C�rY�D@ޣ0��I�던ZV����y��]�.4��qN'�y��|u������6]R�d��� ]4\�1)V�o��ѷPDX���k+g_�ߜP��[£.9;H�oKe�����l��f�S$�]RWNدM�N���}9[7�;[���>��R���-���*3�S�М�%�As�KBlSh�{��?oW�/�j�|�9�k��Ư*���9�K�e��<]��,Ǒm<�+W,	�@˛���hkZ:������q/3�O�MX��6��/j�o��"m=I���L��yF����븖ֻA���8��E�A�Ow<5q#�/��/���t��ٺ{��Wu�ښ�E*̔5�k������_���D6���o$��l�ߣ:~�/Ӿ�x�n&�/�I�:N���n�+��22�=5�ݤ5uW�������a��{�W{�}��
���ێ~�b�^T����=0���c��x�u���7���>Igeꦽu�}���]�}2�?�:�iz�3V�NJY4_�G��}��&Fd�دS㛼�E�5��e���[�Α6[�l߶��򪧄�5����Ǐ=�������`x��z��=�Q�*~�/�?�Ua��R�<}�*v>�~�<�'Ю[<ڨ��Y�}��3��t�	(�,R�i~�d����L�wR����>���:�`�:�X>�t��+�ѹ��T�f�H׼��%�~̩f���c� Δ.*e��RQ�C��\b�L:��?�B�ƿL�:l��ϟ�ɝ}���a��f��'��@ʧJGcn�^^^���m�Bh���Q����u:�y�-��:m�ݠ��ep^%GI=Fa@���Q��JM�<��)ΘQ�r��8ou�z�*�y`}}~Ka��ꏽ�z����>�wp���/�-��)]m�s�Z��Hb���<d�[!���U��V�ŕ�y�A���+0fei�K���s�T��d,kT��+��ݧ=}|��R]�!us��I�\�Մ~�{�5���c�N(�@-6�F[wl8Jϔ�7���23x�퉃|�������{K@�x�YV+}qE��=O��)�����:�f�S ���z��/�^���&��L0O�� z`-��-��åq���\4�IN}���ߛw��'��������e^�R��թ:��6��<�h_ԧY�|:XV�������-��Dm�U+�U��et3��-�|��h`�
�	�g�=~2���(K�tn(�ɫΤ��Yl�cd׶VQ�{��zvwz�(����D��1��n<'�k��ZC���[Y��y��ƽ2��)Y��4dz�c6U��e�ܲ��j��� :n�W#�^\�œ����=gwV�n)x]�϶���*l�E��E����yp��ޟ-t�~wHN�!�����gײ��ݝv�S��I:�
c'��Su��t�vS>�ꆤ����s+]�����/�톋��D��~�>��͞�w&Qqx��,,���\T��5���gR�����*���u8Φw�������)'Ʒ�9�;۲3]C��Z-����jnS�6�����2uE����@����>8j {���,����Egr�#�W\BޚȚ�*���J��=$μ����K{�������[h�Xo���P�:�-�0w8���]��6-gA1�@R�/O�_�=9�:���W�����Ma�J�}(�Z���j��EC���}mH��{�x�u����p�>��^vT�,��3��^�U��mP	��I��m:��c��CanȼS����0����U��u̍ߢ�I:k�<�=0��яw�ta���_�mL���ܸ�k��ѥ����!���w��R�����*�S����̳�D�T�A��g���u2����]K7�U���+z}�C+O��v��\-��^������������6_��������))���˧<+��n�`�s�k�|�N#/����:�n��{�NhF�:˽1��rx�Az���Kd��y���e�Z�KjЩ���t`�S�s��і�r�U�M�;��]:�ϡ(�qT	�bg�m����ꄔS!��:�����ns�l�K"Ƿz�e��_�9�D�Cn�n�Q.gx	;$LJ�tEmmG�Չ�|-�a۞�X�W�F��\�FZ]n�nx�� ��F�+�tڙ�fe3���UNnNI϶��l��ɇ֊����͘��>�7�KǧHj5ݨWQ0U٬�J\�f_Q{��J�v��$Rsk�Umvr�6�fZ��Q�C�sIwc�Bo��f�Na+\X�zV�+��[Ƅ8�]�z`}3+8�6�ͣ��<*�.�Ѹlr�N�F���8��&e��د�O3�u��K�~������4nt�#T2�^L�͸�ý�����59�ƙ���B6;*{���v�-7��˄�����:7�K{蠃�N`����*���C��?aZg�~%W�$|�F�ÿT��b�'\Odn��U���s���N��37��Uw��k���u�C!_�|p"}���s�9�ש���Gm������`���~9{n��8ʥx���V5V;��^W��ʘ�~'3@2��Pv+*�׶TΊ9.��r�^V�y���>u��l����E�:�亘ų�ڮ�{|/���;qr��+��k�l++'��{#P�n<�S;E@h�A�p���&��S̽wP���7y���ΟI��#76�k�C̊~�����&xd�}�L�����	Sk]X^���y�e����g��\=X�d��,_���n{�q�e�`��� �(_�=\.��ʕjhV���5Ô<�w ����V��~u��=lq��v�v��c0��Q�'�@@�$ar�O��]D�V���](�Nn��8}��u����R)��{ޗY�q��'�u�V��>��6�v_X��_k�Ǻ�S�ts��3��lZ�*ڭ�v��^nF�뎼�Vh��b�^з�'k���tTZBeѡˀ�5Et���&�r�:pj�㝏�Z�.�������M�ϣ]<�xO��7n���f�z��()�|O3�J�i����\�@�ƏO�����qW�{���>:���{��tF�;�&��S_q .����ӧӾ�xa�'V���-��+ށ����N�>.}���^Vi��.][3jd�=�ں��L\� ��tQ���I6xW�^��l�mo
���������Y�s�K�5�+! �z�U݁h�?c�>��|���$�uxTK�f�Ӟ�]����Έw���䝚)�	=�	z2������K�N[P+�8�z+��$��Y;0���]��)K�]�Hm������#ԝFT�_C�K/��q��*�NXo��X���H:Y=�L-��c�o�l9�?wz���������_�ýz���W\�U=+\�j����p޸'Kh\��q�cߌ9��~�_�_yQ;�,u��;Ӳ��j['�e3�9US�yK�SWQ;x���~�`�ˤV�0��"z�>���99u�Xl����2�Wc�A�Q*�G\Cj�}ߌ�Uk�<���߬��^��A�lj�{Oe�����Le~��mZ�u�Ns;����ƌ(ͫ�u[Qʅ܍ۜ�����ٝ���Y\X��'�#M��8�
g.8�gq��K����r������2�v�W�i��w4�؍=ͻ�Cr��s���p�K�����י���Y��;��ι���6wÑة}^�P�m�7Y�+.�o^�/V��,��ˌ� Δ.*e��TQ�C]�l;���z����-�{ы��gx�\�Mg�ީF��&|g���{���1K�ݑ\Hu���XZ��)�P[>_F:m�ݠ���Y\�\�i$�0�Y}P�fS�=99��2�\y�]ĳ}on*��R���Ny����F\7vÁD�@�\jH'ѓ���ܯN�j��`?����S.㲬.>���;�����=���o��.i��1E�0�儸� �wx� t7:�)���\moW�Jv��|��m��;;s���_U��'��s�����ﵓ�~���L}�d�	<��GY�8�T����Zuw�9�=����n{|=�w�ψ�h��f��;t%Ar{@������(J�tn(�ɬ�A�q*����.r����B#R��ҖK�PM�I��,��3�}r��+��}D#�~�������5]�[A�;��\�ǲ�{AS:m2��q+�b0�D{�4Ү��4��j��Jaq0����ӻ:fP�ށw]��o�_�T���ߗ!���=M��:��l���-̮<!t��N�$���>��}<^�"��/��gV,G�����q����j�������큥�d{>ח �t�z��Zr}���\c�ͫ�-��E�����;���wJ�q�^�N�O����Bs[�X�/&}"�����:��^)����x�҆X���^�2��i:}����T>�SOz9��ec븝�ͻ`?E�x��xʞ�B�g����>7Ŝ���a��ܟ�]_��Fu */z�*���3q�bHu���]׭�8�z�n��w�b��S��'��0�B_.�5�J�G�\�V����$��k�E��]S�C��ڼ��t��C��|�W�ʝ7Y=�axѝ�R�x��L1��xâ�n�u�3�`^8
�!ތ-�����~�K�gD*����i'KG�M����7��BW�f�~�C��q�(γq�*�p�]���O��^{�w��R�������LK��J�3�,۽�R��I��5�+��y���ԣB�V+R����B;q:�l�[>��+WkQ�ۮ>`�(��u���Jxm��g��p��n�`�G<v�ח�H+bmEF��,�@N+6���Es��"}+�zb��K�vK<�ƴ7:`�Bĥ(��i�Ǉq��A5b�3�p/)���{M����P*���
����kw�(���ޠu�Ob��.ʙ�*�Oc8y����RώS����+�%՚r�⛊��p8����|���R�fQ(���2��� s��p�Ͼ�
#�������x9b���e��`z�p��n�~n��v�%Q�`CU�$L������[�ثĲ-�%�\:Ǽ���k�-&� ��->�m�?;��S.g�	;$R�C�>-"�����B���E�Q�9W�m�3k���K��M��t���xR���6�t{��Z��{� z9(�-Qp}>�ଊ��Q��Zn#���mUQ腒�4n!�@k�#T33�|���.�ޙt��k�U2~��g��rz8#p�T�;��دDn�Ӫ�P�uZa���:7��*1����Mn�^�j��yf�K�>:=�L.��j^\�I�}�H;��v���V	�?>
y�xB�K��Yy�FgHޞq���^3�~�񿰢s�yAf�����Q~xC�_�C9���V�Ȟ�:���-�=�w���>r����}�+�Ű�t�s/�0�j�|ָ����sy�9O�`���jZ'|2��Ϭ��<ܕ�WO�Uù�p��I΋_�Ꭺ�z�~�^4w�ڿ�I���V�<J�t"h1�Sj��V�u4o���϶a*�R)V���3n�M�=�Iv,��5ӆ��c2���Ar�t�l��w�D��S�k���PAd�r�Ž�1%d�p��a,\ZKyd�H=��u��u��jF�<��Gس4m����zh�D�'��uf�R#y�tu#����f>嫂��oSv�����A]�D@�A�h���/�b	Ff��"���X�8IJ�]A��34R�K�w�JC/1
�=�y�kve`�ͬ�p=Ƅ �Y�|�+:��7�98q��l�·¦+�����+>BU��,j�#i��J���K���mɔ�o]_:�[�.&OA��)�%�U>w4h��/�� �k/��.H��4R�Gg�(5!����p�z�I(|�j�!��u�y�����_(��ww�ޠ�t���At��w��j:N;�pg([b���Eq� �nB��1��Z����"����V�aԆ�ndn����(����b6�I�)�Q����ݡK��Y��^��q8N�1��rE�G�6ҧ�+�f���&X�W�������*��S��7�] �����6��r���mMN�^�SO;7Nm�+i�������2�!c2��ҨzƱv�[�Ud�;����VZhm�]첢�M˷4��KV�7}��q����`�z��֋�s�+�멉�%!\�5-��1�H���;��v�;�*�@�c.M�>���d��I�y�0�ڸ�NQ�����qe8RҺ��a֭c[X:]ХF�����5����Gc�n+!a�Y�,3KU�ovwZ�
����`IA��{�(��j�Z��+�6V����0H�EZj�6dсƃ_�+�T��]M�.���*q3Ͳ�)<+����V��]49�y���
�	���x�:"������<@#F<AMrJ��!�ju�&���8�05}(���7-k�,6�	g�����.*yF57!�����s�S+ObO5�3)��W����T.qY��k�'0���eɦ���ʰ�o�u��-���۷�:�r�{><[�+�ތ*ŏ������ֽ����	��m-(e_b._f)Y/�ٽw�5q�2���+u_=�d�U�W��x쵊�sv_5\�3�ZG!�Ж/3n���s�hU���J"�B+�s�7oq]��B\k.���8��l����_9P�Íҵ*�������EN/>�_\���хj:TbX�Nv�e�WDz��6�����e`}��.L�DX�\E7Y�ew|�Qc��k�Θ�WH�yr��F�-��}�T��/;2��E� ���͞�t!��-��V�z���%�z�;Y�+E�w׍�t�/���$�����:_ga\�U�V2r��n`���(T���m�u�)k-H��
�!�5}�Y�>7Ws�����uo�4����$1Ns\66134�i����bBR"LHdCDd�!�H��4H�f�i	��& ��9"��#0�+�� �6$D�X4�Q��Jb$�PF3H%22l4�0Ƃ)�S�YH�4�Bc&S��\�&'I���d���+�`ѣ$�Щ�0)���$d�L�&N8&�8`�a�$ɔJ2�P$��&�8,����$aM\\�$�XLs�!B 	,�
��˗���.M��˄��73��&L��H�2�+�3��q4���a4�!CD�D�R2C���Ja��(U
 |>�P� �l��/&*w�P�`��{�S[�Ć ��e�N���ۋ������7I�v>;܃�F�"N�Ť����Ϋ��9ծ_���� ʨW�Zon\��ˀ�0�d�ܧ�{��p��;��~�3�s����ܙ�@�5���L�/$��g���·q2�b��	R���]0o�:�>N[=:�f�ao:���R�7x���S^F����q{$���'�_."����K�:���\F'lh]獰b�'�q��ҟF>�:�:��yЦ��~%�GI=FP�=Ċ��.�w��\tn�S����n�ާx���}/��W����=��a�y\'�ݻ��%�D@ޣ0�L�I�q����0��r�nF[]G��?��L�-}qW-��x�S�֍&���t�ДIS�@��Ԑ�9�_�.v�uMK �΂��+�P���q��G�ϴ�s��M�K�fm���v���{ӆ�v��$�wRs&�=$L�T�83������Fr�tz�ĳ2]�UK�r�p����G��ېͲFQ��ό�r��uxu��9�5�+�:!�7�tbk��O0jzs`U��]�ؚw}��yJ���#Q譗�$�N�����b���x-�~���S��6
W���mz�3΀Դ�Ok6��H�[ݻJ�^�Ծj�������6�j�n��^�QSދ˧��-�C�����m�و:�y�`�R�- ����K�c���͐8�Ieӱ���Ysr�up"��\��˶Mr�e����v�����u-����5�d�d�L-�9����K��g�bw��o%�U�������!�����~�=���D-t��
v}�X��T�^J'(���R|canUy��ơ��1�N�M��xNgKf��}l{�U<'��jZ���?^
��}�ؓθn�e��`Y��;��2p�����w^��d�O�ʁ^��M&Y8�u�6�;��В���pھ��8_�e��w��x��l%��5�����]Q�@u��[��2����=Rd�f*��e���O��C�R*�~/,�!��1P�|�B�e��W�l�iݳ��NM�l�*3��2�ª����T�z��z�p{�5�b�w�Q����3	��=H]L���=9m�Z��We󅿽{���������߯�Kg=��� �iCȹ,�g�*��#s�@F�èϾyx��]PVAa}Fw�ŗb~.�P���>�r��c���y�#/���~��O3�bw������
� �_�|-���=q�V+}qW�����y9v���ގ�P E���,~ɫ��ּ���\�qw} MU���p���e�4�AY�T�ї�4��{BN�����I����y������jr�f�\��v���gR���vc��u���n�s+xq�r�
��o3{�/zW/�G�l�}�}����Z��r7/w�e��3�&A�_l���	V�3��t�7�ޮ�N�1�>�h��#D��3�zwC����/��N]+�d_�d�_GT����'�M��:�{��µ�dd;�J�B���G�/\����s����/>40C�"qrx��EzVӣtWd׸��Z�K&����2��Sf���s�o��oܕ2\2��B��I���D�!i�5ߠv��vr��{��gb��SV]G*��Or�0�MQ�)RT�¸��\t�z��2�R�W��5<��TY��w՘o�z_��Zn=��ܝޕ�@tTy�!:�]
~�k�=S��Ey�L��'��<X쁓��W�����i:}�)���\?*�xc���s+*��dڐ��e^>��{O��f��lϏ}>ȉ�?P����Q�pk��9�(
�ۆ;���\]g8���F�ﶍ���u��u֣�n�n�]���T������{���Ma��Qn҇N�u2}j����X�
�V���R����}�y\3�3�~���0�Aم�TP�
4+�����E��l�{RWV�����j4ï$�w�r�<ƥ3A�eA�H{.~hk���{� .:�6����zm%�Ժ1�NI��ͫ�9��gWB�/6(�J��N��]κ��U�!��3kNe<���0������w2J�+�5�
�s��C��{}�}?���/F싈�<��?S�N�1��Y|.z�m��'L�j�����y�9�TӚ. ��m�e鿶���n��Z��1�e��7��j��}+/��/*z��t�{��&�3z1�n͂O9���rJR��z�Q��Z�z��>�!��юB;9{.����j�C�������8�nk8�
���P����<=޺L��n�Uķ|0L���%�i^��k��_��$[Rp�Ǔ�9t�х��F����F@r
[$Y<�}��(t�[�T�:������,�r_����lx�m���a=n�鿢����d��@]I��r��B���W����>�~�x�:�����|��sĵ�>���X�;��2�z�BG��j�A�`OV�4Qޞ��(�r�#6Ჹ	�j]n�nx�:`~F�B�@�7P\`Μ�Y����:ٚ ��l8����*[9F�i����?Cj���L�7۠5��r���~�]ۭ��v�S���51Ǧ���|��ᑖ�ح�X{U��I�i��6��Pqギ�~��rE�X��}�}�J�l*�����2�7�!���ef-k��(1L2p��'��`���ū8�5�I��2Ws�ou+�3�U����]��CN�B�.�z�Гn0���a"n�#{�3���x	�+5�*�W>����;qcY����5E�� �:��l�id�|=0��Vu/�U��i��VA�Z��t��t�`��e�z�s��h��x,Z�T��D��c�@��
������b�%¼��~�w���6�� U��cЪ��>�O�����q�k��s"�,��3�kF�3� �z��fz.|��Q󌝙�{���@
�r�#��nJwQ���:7���Μ��-�<u�1��^tL�q3�4g*�*�7r�4F�vL��S̽wP����v��RK6����t=���ι�.��O��q�I�XPN��S/�/mP�6�Յ�K�ǝ^���F�~k|��v?	���].�'||:�QY^�����|��NťV'��*S׫b�:<׍��|gC�3�c���6��Mc0��(�:I�W�@����&ٱ��.3�P�k�����y��Sw�����t0���\��w��H��a@�~��8�og���6�~��.	�W���j)�-��r��Cu�I�����Л�L�=,�1QQF`���
���\U�O�Y�U�|�r�s���oG�Pդ؈~	�[��4U<ü0���Nl��J�}Ӛ}�3T8�B�荖!���V ����b���g�`�5y�E;�C��ꚜz9lR��F�i���c�z;�P��`,�Y݋�Ubo���T�$8�����^��|:�q���ˎN�>�.}���^Vp�� �Z����G�p��Ze�̓��jOt�� �<+�+N��ͭ�Q�˭Ѵ��,ۅ:b����]]�h���'ύx5ď}�.vl��;^f�E9�5}7���/�S?�~Z����%���u/(��w��6ܸ��z+e��5��������koc �?i�2*�[�!|<\
�ۘ+���Uxhp���p��u7� ��?`�kʐk�OW��n�Z���^�Z���?���3��V����~�=���-t�9��%��V����s���Y"FI��GW���2��C��S�$�'�#:S7��cʪ��t�59�WQ;x���Ot��PwW��\u9��d�8r�e��8ת��̞7�������'!��=��2��je^���|�����fޣ��g2||J�::��tp\T���%ׅ[l��b��+;}�}���zx��u���X����d_�mO~%+�PgJS/����"�h��UzI�o�9�IJ���Y#KKL<|���9��+)�C���K4=&�.�:H�l��������*���Kf���̭6+:ySǋ�I{V�1�\Z�PKspN���@�-�J/d�zu�(M��"ٺ*���H��a�'LJ��S]L=�����f��fޞ��օk��.1C�3Н6{���B��1k�R���N����q����)S���[%J�g煻�B����b��x1�l�c��v���Y\�%GI<�փ��6�N�Wg)�8��*:⌦_��]ĳp�m�\JV���r��c��y�#�a�xB�6��1 ���W�#�F�M�H�5'��S�#��V+}qW��}��O��9�r0���z9��K��v9E��"�S�4����Qy�@y|=��_�Fd)h��J;=/�l�������G}���g�ϯ�8�q��N_��ّq
d�_uI�m?I��B��:�{�,,�'�nT.��i�����I�d[���A��Qd3|O!1p:�b\q�'n�s�;�+i��"��ޚ{<𩾛z�4�t.ޢm��䩒��r���F��R~���� �ZUG{U���j��ݖ�3%ßenQ�r��̸zo����]���t�00��Fhe�ːJ7Ѱ��3��u��*�����᳓Ყ<}E�z{��Zo�yp������@:7�t�x|љ
�1$#�������xU�;�7�maĭ<FQ8������th��K����4��r�ܒ�F�)����2<����=��@w���h��զ]H�Ok�W�� �v�=��J�54�.Ź�5��y�p���i��C���p�͛nlrgTc�֮,��]��pг���;�,�i��@ URg�J0ԙ~0i�ܣ:�T���s�u�k�y���w��W��H͝�|�X�C'��Q�'��>�Τ�3
G=����{0��9��*�y��ucw]{�z�gǼ�'vw�?"�pΖ�B�ZZ�3�Ϻ=����p:��|��|���wM��J���}���5mO���J�d<+y0)�錭��=��mG�*�omPxmPa`n��S�������DS�j�W�ީ�1u�9X$Y�y��N�'�ѕQ�F_��J;�]���O��!���p�O���7���F:.�9�_�<���t-��U:	;Q3�L|T+�������ER����rZ\k�'�~���:p�=lq��q������(� odA����k�ZSî�3��p�{n�猦L^�f���ߡ�^�\�Ѓ��v��'�;����v�/��t7����H�y��������v�7��{��w��n3]���)�C��7>n�I�7pt�}X��f�0!�x���˽�C+�S?��m�K�qJ�n��2��Q�(��0>���պ�n�V<v��sa��H�L��`�\�����k����6��O��������I��k��v���P�%��n�%�2{35uچ��������Q4Ww��۲�9�"�J��]:��MK�{��z��g��s��醹ox�ɫCź�_��M�� �~wQ
e̯l;1]�j*5F���C�"迏�����7E�M{.9��HTb]N�D&�~��1���-ӆ�*F�7��KxO��|iL�fgQ��O�K��WR��7�+Os�C�]Tͬ�ɢ���G(���bw��W�����$]WL3�<P�|���km���-:���W�	q�w����W_�5����ه��Tn<�@;Cw�n4�3�zY=0�>XԼ8.�V���b۱_r���oR�Uc�����]s�s@�xPϺ�S�q��`1��*����2�x�:TL��7�KZY�L�n� ^>�9U;�}��U���y\//�#��K'3�๽� ����r�c(�}ANL�����F`
�r�"��nN;����mW�s�����xF�����+�.2\�� `�L�F��J����B^�!VL�e3���:����n��y�ܽ�*��{P���N~�w/���h�Q'I��	h�i~�W��J���C�
�f�+��EQY�o:F�6U��}^�W�^8u3�#l7�J����u c�J�L�n���@�"�cVh�i3�a��J���yW�9iW���:���;�vV[����*�XYĦaUɼ�Ħ���*�T[�h�ϗo^���JV����"o�vq؝ŽFK���~}��ʿ�/����W�������ypǲ��ݴ��zK6b�NV{���)	��!�:��t�m\=�B��a�\�j�OQ���H6��إ �T�U&1O*�e��Q.�{ET����m4{\��:�p�7n��\�k�D���i5��~�����ˮ�j��\oդ�-���ǖ�������|s�n�i7�荸�v��/:���ui�ދU�5q�OK� ɨ$�h6
��0���q��|\�Kg>/+�V�5wq��P�Y�d����>�F^̒�GT��6vH�N�Uԭ824�{�*2�[���ށ*z*��p�wm�p�s����Ȇi�˞S�w�9�t���b?˰����l��,����z�%�<J�},��Ԯ���I٣mˁ���z*6_��\Q;C�n�Z�ȝ�-Ao�~��{;W�zq*��᧮�ێ�y'wB�:��`���(W��Rd�v<c�w�!����U
g|����)�1��t��ҷ����[�UOO�����V�����\u��{+����nkz��H2&_�.��S���سs��#�����e@,wE+P�@��Ch�G�(\W��v�����C��zizi��u��'%�|r!�������=˳�8����m�ve���}��Ȭw!�oe�&��Ml��Mu�vf�v6Ӡ��E1
���4/%�V%�սx��z+�-�۰�;�������d����̺δ@/��@��&�fC�}��󕝓h �صR��U�εC�eM;s�ݡ�ʔ쩕r�RU��������ð�^G�n��̭�!qu+��u�ΚP=].���1k�n@����o�0�����bH]�Â��X���w�c���v �r�:���)�v�7��]���xL�#Tʴ�sC�}O�ݭ�J��B*yo
$1�j-aE��Y0`0ǫ����D��ٙg�6�2�ɸ���@o3���F@εYM��!t��L�>X���);|o/Z4U�_	Uo�(�Sux�VY9�Io^5����{��&��d��;6��Oe��}�����j`�LZ:�Z:���e��с���y`hʅ
�{;%Wf�sI�|.���<��66���V%D�YkHHMx����wX-�ī��V@_*VƖ!Z^�����+�dh�(�z�gi��}�)�� ��>.�Dq�k4���>�w���v�eVH�T�֎7z��Wf[ğN���7:��w�-T&���������Z�����&nen�qNt%(��߅ъ���_�7�{�Î��n���ݷ��^��IvV��S�L�ݩ�����C� �]���\�F(ʵ�K;Uvͥ���fڼ�����}N�w^�y��J��K�'���m��k �H��j�~o���l�$�;+��JP�x�I{�s�|e���U�#�NJ�58�Uz�Q(U#�n����f-b�vv�t@�\e^��K�*@���g]*��*� �sq
�n�\@�n�"�9ð�5# u�=��xk��ڴv�!�_D�!�sG0��Vv�j�����]Xm���G��%��@��G�3g=�<G7�:�e�-bꝧp\����e��b���q���rc5g|�cWXZ)7�:�e�\�נE�b|��oe�=��2K̻��x��J�s�ݶ��4�;ia��s�o	��SP7�9	�v:��π�c�����C��V'{DT��)�����K��C��]��3'��b0��Z�A��Bd�2n�U��[��qf�6d5Kr�i�6]\ͤf�V*wn�]>��ә}�,#dR��:1_+��]o5�u˾gg�h����w�tzzXO�G-К���n����R����yO ��0!,g�r�ҾV��9�So�mx�GBy��|�9�u�X.��Z���fM���*�e��a�|7��v,����<�t���Z���@t�}yj��VS҈�G����o˶��ݹ����.=!�X�-�r4����Cs�qWa�>��V(�Hh�OgWbf�������dLi2��ȉ��b���ɉ�L2L�cFH�Q,@���Lѩ�Jb��`�H�# @2(ɊAA���@d�H����B�FDCL��h��F#@ �F�D�0$���&�DTH�jI�h�b-	JD��1��21"QHh�b0�&L��IIe��Q���Ȳ)�DL ��)"�!���i��*@&ѓF)ТDA6'����`F���0��DD�"	4�%�e�DheL��b��YBb$�!#Dʢ!$�F�B�cF�EY1L�FX�a��2`����%��3(��A�(P�6�$����_}|���]�{�%�[lZD�n��n�X�k`��������M��j���r���}�j�u�]+v�d;ԣ@�"Wq�`g��~`�ojտ�^0>�~��[�UO	�s�9��wPt}��v���l�q�=��y�_�q`G�a�j�!�AS�\W���Ƨ�<}�*G���Re2ɾ[,�[K��;�)fZ����G7z�w�}ߦ�Xe��w�p䤼-�KGJk�8$��`�9�+\i�xN�S���P���w��xS��|��7|��1y�S����B�.���m/�w�K�������������)���]�E��1��gX��GݞsZ�j�Y�g�=^C���9�󗏪���K�w��F̴L�7�t�?B���^�-�c�l�1�m�A�S��\�g���"a���"�4�D����	8�������Y�kn*�%+x}�5;��@-7:�g�o[o����x�O����
'�H\Ԗ��qۍuaq��r��AS�{L�=���ǤW��>ʟWO���N]���y�*i�D���w���J�	�V�����`�/�<s]�]����+,.˲՘y>v���m�N_��ّ)��uI�5���Ʌ㿍�ߦ�'6f L4��5Xv區a�����H�Kd����!�8WT���=���YM{R����D�tcU�ɩj�����g,l���qT��J}�L��U����!�=��n�Y]����;_r��H7���]IF�����ήմ����G^��Ύ��-�y�mu�����Y��ϑ+��G�T+U��;�f9؝��[;N���Nr�{��}-Qts�j�v�;\��.��2_�9`c�#q�)?\
��N�c��=@A�R�*.�QSʳ���s.���{l6����@:�큥��p�R���2�L��p�3�X�K l+��_�o��Y�@��t�7�^������|7G�ѵ�����a��j�u�П4��/�/&}{,#Ŏ�8ש��륤���}��랳����ԭ���ue���1��;ǜ>������M�hύ�rr�e��1`�������';���&5Ww���;Ȕ�� {ݗ�O�=��wܪ��ޢ,m�N���2TOȸͧ�Ү}�>�<�:t�����d�/�h!GS��;��:���N���:o�,��������qTY��W]U��� �l�atnȸ�S���� ����Y|3�����Ȯ�qqt\�qs��jO#Pg����ܨ���]�����9��;��W�p�=���|xf	���Nzc,���e>�B�F�]������j��0�B��5=�����<6��M
�kӎ퉞���F�W˸�Q�6b��/��eng,�0d"��Ֆ��]h-���\�j��g�W
�}8�n�}6�����!�|6���z	=S."@��b�[�c��Q����\4��	�I._^V\��z|}�6��i�|�G,녾��c/� �(҂�|e0:x)��R��u���Rcϕ_v�=��(��c��I÷��];�ax\�j:�d ��B�u%�v���櫃�{:����ek]���mZ�������2��NB2Q� .W�<��ޗ�=�^�}ҍ9&߫(��R+=�[�G�'��%:Jaς&�u�[���mL�3=9�M8�j�l�=���{eQ��+6����Te����n� ��ȟs���Z;�;��N>�� UN��oftS#�������*S9F�V���ͫ�+�и�k�ʇ{����v�G��'�Pˍ��&�:a�>�6����[n�L�
N7'?z�d��4wZn�~��O��z��G̨7��,ޗ�|n4�z�zau��
�^��m)��]�?=���K:re�md�����c����-t9��l3��vl�q[�8�W{��>�I��Z'�.~gK[�<�+������5u�].�͠i#���g*u��iN����r=y�A�Y�+lV��l}��<�7�jhy\��e�+�qMԵ��;�R�b �Ax�'s�y��s�X�M��w��lҎ�&��c+/oE���3�_R�~5�l���_^>�=���>��>r����}�+�������ZaM[*7���;��3��w�|{jת��ƥ�{ц��ܺȾ�I�9�5t�Uû���/*�kv�M���t^�9%��'�\L�vc�N���[*G�v\FL��s̽��ã	�Q����m�>��UC�R*����ѿMD�t�����O�_�T�g�Nl�P������n�S�F�uS��=�X[-�N���)�q�G�e�/d���,�����{Em�9Gn�<q�'���\_*�9Θ������A����)�f�\�k�t��Pa�dU�����Q�~2L|s��˨�q
״P�I�5���r<v��>+���8�YG�Xs�D��{E^�T��f=J��o�y��uB��Ew��{�w/�w�֍&�����E[P����Zډ˗�^̜�� �$�J�i~���o	�o'iAs�-�����T�H5C�f�js�)�^q*���IC#�J�;$L�\*��Zpg��f�o
�������j�X��V�E�[�� ̈́{>�]���i�y&@ݏn���^��nIZʀ+�Ǩ�w'V�f>�q�=q�{���h$�9>Xs�u*�@bh0J�t������2K-��WbM)���������q�	������W�<����%H!�2\Y��G�z�i���/h��Q(�.|�~F�|��"��T���f9�ë¥N�B��a�\�j�����{�Vo��}ΈV�]ы��vh�r�kBb�K�$�D��zam���]Z�U�������Y�7�{<Ʒ<3�����N��!ԶP��+�~�'f��2���s�[�3;�Ӫ19���u���7����c�ʩ��-t��
v|�Ս�Τ��<͞5=��G���2t����3&�^���5+	���L�G���򪧄��1�O�ægّ~7�~�2S�A~�k�k�,��a��+�3�z�U�I�Oɕ�����fn�L^�Ƕwr����o�x��:�y�q�ߝ���K��#�%%�l%��5��ʠ�s!dL���.��ҩ^���k�@��F;C�\˃��3���׬�խi��'��n����^���xVRo3HV�R��k�÷A���z0�`��P����g���B��1p��(��t��� t��͹A�ܯԙ�Ec����n�
^���b��x=�%�����v���U��C�'Y�.��}7ד�^����s�p̴�Y��]l�C�����u����FҾpnX嫸�Dv�V�y��er��vᖯ�7�,�d�e���n�a�KhK`��Y���q�1%-Ib��:�
����p�X+z�ɶ�N����+�8�md�$ZN�!������d �T��2��;��\��eRڊؔ���CS�raռe�p�:��g�6��"�˾�l�P��5���J�W���4Oj)�-�q�@iM��zfw��gT��%ޔ�jN��vF]:�f�L��@{&@s*�nL��q\Q�� ֱ6���r�:p�8��L�7��E��6۸���ݳ"��G��� m2y��;>m��⏮<ҹ���8�9��!oY˩�o����Ȕ����j�j#��;�?TΓ�NLm��=��Q�2a�e*7G�M\v�r��o��rR�j�?B7;�m�d	�љr�n=R\oy�2��d/�1蕵�}[9W�e��q���mMQ厀um�K���Ѩת�����|+��_�,��|���ȧY�(�/O}�*Jkʻ߉�;6r����نyu�x�T_в�	�}�}b�����x�Kp)�c��KI��ݔ�v� �F�U�[Xj�:n�ƿ�*ia�CN+�Y��'o�߯4�H͜��N�쁓�\T����cb���"�G��G�	J�9��4)!]/���(^۟ـ��cr�9������\�S�<��j���v�����=�uI`p��s|��Z7Q�Y��S)ݛᲚ}K����G|]���L];'k�q�w��NH�q��;������n_o] /\1Ω���3��\ws�D-���h�wl�^��U��LC<���Eײ�	�>"v@��}�W���|���t��|�n�7����ʝ5Жv��!���==�=���fc�h�T;�U�iH	t@ڠ����G��P�H>�;�Ƨd���8[�|�gK��=���t�����3�
��/��P%����K��юC/3��:��w91������_Oޤ�Gz%��^Ĥtt��T+��Jb�66�Μ�tn�5��3���ڙ�_\G܋ΐ����!y��2���(҂�@G�iO ��ϣ�a^{)�n�>���r�P�)���;\u�����v~�d>.K5�G*3�B�o�!��!�S��[%O�Ғ ��e����p����7��o��7N���2Q>oT�]蚭�5�̱)�	�12�������:�+[�#�&�An���|7۬�ms��Lu�5$'8�2�k�29��D�K�tn�ӕy�ͮB�-.�F�M��r/��	�o)��������7Q�פX�e�G綢�Ț<x��N�}=�si�.�O;����3
���p�lFS:z�|�
篯�C����Jm��c{1�ɘh��t�$k1��˱\�x��R��B���L;�>�%��2pK.�xu��� �B�kZ䀹���R��(�׵�q�~8̮��2;�\>��R��*�;)������&�Q�:���7@k�B5C/헓&����Ca�>��8/쵶�%�j}5�g��q���Z��j�μ��$��ǡk�to�T��w�oK�>7������X��C��sS�����1�m�4W:d�6�wۿ=Ξ���Dc�/�+vl����8دp�g�8�F1	���1���wv+)�J��[�����cЪ��>�T��Ϛ���k��o�o:z���.�W7ʖʎ��'���_�ax��
ng�IL���H^��GK�ܗS�;�#7��S�Z���=�&.��P�fS�ڧd�Ĩ�/�
��R3ň��e�W��%8g�t��/��{q��e��%������=�i��w�o��.|ft��&t+��}1{j��޲9��)^uX�y�.V�5�T�������ވv��M{���2���k�(	�B�3�m{�~�{�.t��t��άN'L`�xy�:���SX�?D��B:I�\L��Z�� �����ܓ5D0%w:P��]�Μ?��e p�� �=��:�Bƅ}���eo�|��
�f�Q��v�!��Z�J�)R�A��7��6bjƃbY�;�z���6_'�%�j���竣���ˢF+<��v�s���rva�@�~$<����KT�ET���[Mߦ0��=ΝM�+{�\n誜���Q�a��!���Wd�������*�[�p�����n�i8�qu](%^�S;�h�%~dy�V]�$���@�� ��A����������D�P��1���z{��lg��ߴ�,��㛼�]y����(WT��4���\T�824�{ԑ�N�R���oۜ�2FHq~ݮ��|K>.|�~F�4ɌW.zl���U�Y�B�{�+��\�{��7=�W��5�M�-7��p�]ы䝚7�r�k���z4�2ONh���ӕQ��ߙ����J>z��Ra��6�N��[�e!��w��U�!T�P?Ew2Iۜ�y�;#��bf�5��2Ǧ\	�1ҧ<s�^�ٽlhܫ�7�S�它5q�V캪3 �9�~y��75��z7A�_�G��NT����2�]z�5+	���L�{o��|���=6m�T�]�y�>ν�O-h��p�����ߕϤ���`��+�3�z+�Zl��'���|��t��׃퓃D����,�Y2������}v���X̋qݫ�s]>��g]���'���R��	<���]�0A�h��.LP�Xd{�M]�՘�es񭛏�]�u���>W���֖l�ދ�V�6�ö���Ɍ����������O��6_3��ec��Kר��y3�a}'Nؙb�KGO���s�{G���s��ͫ�<���*P�j�E�W\���̈́���ʝ4=��t¼Wc�l���7��|-͞�u��!��6h5���.1C�3�	�g�N�=��0��Q'���=;w�}w9��j$�fc���EL�7�t�/Z^��in�{KG=��Z� ���zC=��`���1u��\Q<_�t���0�L�
ACv�D���QJR����5;�h�nD�����Oa��;�L�8���~�%R���I@L���ҡ[��s9.�%������%���V��'��n�ˊuhͩ�Q��#OW� 8Jt��쪕@l���~�t;��>�.3]!�:H�s�g<N�n�r��2%�Bށ�A��8x�D����#>]Jh:��såkz�ˎ]l!��Yd3h���z+U\e���/����d��3��*\M�9����j�Pt�Y��T�{��K��R(��ֶ���V���ŵZ����UZ�o�֫Z�uZ�km���ֶ��V����j����֫Z��j�km���k[o��U�m�ҵZ���j���+U�m�����֫Z��j����֫Z���Z���kU�m��Z�km�Z�km���e5���0$��!�?���}������(��P ��EPU �P �BJ�(�T��@x 9ȪUUJ(�
JI(��TJ�))T��*%UH@)
���y�D�D��UTT�QP�@����)*T�R�HJP��T���Ғ�V�s��M�H���(صPj��@��6ڲ�-��*Fcd[F��m�tHJ�,�T���q��tU�Sl�Y� �   �   -`   � qںwfv�K��Mj�R���2�*�U2��1�ժ�Lm�be���Vkl�,j�dkEE	�*��n̻V���f�+1f�ݝl���@$46��b������ܮ�(ѤD���jQ�k�mV�&��4�ڒհSZd2 U6�@�օ[iV���3,���l�I24�P��pQ��ѣU��E[P([(m�l��h���jiT4��M���4e*��(��4�([P�%ST� @�*�܁�l�CB���F�U�eR�EV`h(� 0:)]aSM� �4h��P���k"�V��e���+(Q�����B��R�-6� l�mU�Sl��FXҚ�Ԉ�h�"RkV�mii��͘T���E�0�����0��@�&��AU� -��le�Vͪf�Ƶ�Bw�% �R  E<&m*���?T 1  h ���)*���&���44��1 T�bL�yF!�h�Dz���O$"��&�RSQ b 2 4@�12dф�14�&�) h�&��=�4z�(a  44M���?ng��s�?N�����ysǙ�F���κ�H�f'��Y�@�q~T�A�I"u�!�|��U�y$�)Ǽ����CA�?��m���*($SnRI$�-P�F�@�CeD^*���
��!�#��.َ#��+s���� D4qI�K����/����A}���9��
ݏ��9�`a�w���������99�ş��6gg�g:�����XcN�sTڹj�@w�(��0e�U�n�B�4��h8F[ŶMh�J	��Q�!�n�\�Sa�%f��s2�s%���R۫;N���!��d�@��V57t��jbɹ2�T�ͬ7�mGCșq�3�@���i����Z�]�V���VB�	� �଻�5�%(�i�� � ��.�Х�@�"t$�HոS�{vI�$� �ƣ��aT�HV����f��0V�,Gnٙ��]2V�L�KFYtt�iU�1�'Ɉ�4�ݑ�6��0��Z��nػ[&��7�c	˥V��E�Ce̽Hk��,�qj��a�M���m�f�]��{)C�YV��ِ����E�����c�Yz�d��kl�/@�T�Y%�E�+��`�n�Q��c����c�[8V��u³P��0��[,���N��{l�M
�*�YP45؄��E��z�暈�wnG�eˁ�ߖġ��� Nf���� �B�f}�C�&�9FZg��v�5|e�`��naY�����Y��u�B���1�ˆ�Z��4޼�R�,3IZ�V�ĈosL,aSW�	���Ēhk��E�='uf<'wt��7whL���VYߎݽZ��ܫ:E^a�a%轣��:tJ
L�^�	�*U+6+{-<bZѬ�W��b��pF@��݌ٔlZ[�C�Fb�0^ܳM��0�ݭ,*�8u�$�����,R�g�EѼz4��ka&�`8�#(�E�׸E�b���Fyj��U�5K[1b_ڷ8;�`6z�T�M�{�\��E[��7P�sV��՛4/qa��0J�p<����Rʀ%[Z+-L��#u鹢�4{�;H�J��ӝA0x��٤�-��צ��D�HR;�k�S�Fw��kV��q �@�K���Fa�
�n�zr��0�3Z���4NeԺr�[qM��h�hV*z�=�H�aҸv�i+z�������5�طÖ�)�Wb����lm����љw1X�M�[j$j%��,��۵��ޥs�O�CU���!&[f��;`��ۢluW����R9i�d����[�y�R<��.8�����4��}V�aۺT:�lѾoQu¦��$^F]��p� �mD虖S��P62��tN��!�0����;�
�&\lme�C�:-V-�ofk�cFfI���e\��<KfՀvL2�V�aWj�5�2��[���[V�-�H�fl�32��6f�4/kp�w�qfF���\[��q-Nb��s�r�E��-kub�i�I��TOf3�n]�1k��&e��-^�#6ŕ[��ͦ�#�t�NMU ��lvܲ�a���x]����	IE�n�[�N��1r��v��k9L�	�VrnS�u�t�.������+T�h$�;:l��E_�4Ҽ��e�Ҳ�Y/���b2�\�x����O8��4ޛ�ia�B�I�)xDGr$�T�ԫh����nΛͦ�jV�vws�v`K(Y��.]	u����L�����ʁmL8�
$��w7,WB�,�Wg+pd�f��]a�Yt1ӷ��P�Ɍ\���wi2.�������C۷!���g$U1njk.���\����������{�[��j����gRN��`��Ӆ[C�b�NbE��6��C7��Y-�A�ݗj�x��u[p�ò��b������6U���4X�'or쥅C�E�YYV�Fj��0֖@LV��y���}�����ϕW�c�,XwAù�2n��5na�:ɤ�����u���w�Y�����a����P��XSZ�+��?+����:wF�Sj�����tQ��V���Ցe�ĝ�2fZ���	>���Qx��������T�]B�ڼ�%�gIm���Eb3[�fR��F�����&#���a*V;sE᷷�2s(S��M#��͛��U��SNE��[�Ig�goEb&��b����D��{YwdL���iӳGk`���	e���Af�7$��v�V�H���j0$��W*ֻ�	�Ӿ�q(���f��Į��3(��������FF�kK�G �P'" �F��TV�lݒ]w3W�M��h���xx����٩zr�v򘬺l#��m&͜�ٸ.�ݙ���8�0YAT�ڗ�ds3�9{9A��[�:+wCY5oeL/Q1�Pۻ؍e7Y%���̖p����e7�����#���Q�V~��+T�I�]��϶�i��wg��4��e*�N����t���wZ��D����`H {>ŰC��[��`��B�7��P6��@Zʎ�	�8�S6���V�8��F(fkfVZb����`�HǸ��!�o�?n�Y ��՜�.��E��|~\
�Ֆun�x��adU�=������j�J�8��qh��J@,��2�JF�Ӵ���L�jc�`�8ln֢�V7�&�BȽi�m�U,e+ݜ+1�ipH������v�JBjGn�5G���	E�`	�--������Xh���dgҥ�J!V:��؍�g~[��c���&�L�Q�()W2$K�+:����q]�(	�q���_�v�>5���g�i�������M�#j�H��ZNv�$śf�"C,!h�y�Ս.��]\�P�lL�M�Z�eǚ&�5�!Th
@>��v��hЮ�%�x��&��-JڻM'���-P/&�]+��.�!�n�1 �@�m�O$u(]����!F��e�^�g�5�n����ԩ$n�Inj�̨�c�Y�}qk͘���Pí��M�^��TV.�Y��bys*à�YTl��Й��e4m����ʰ�/$�*L#FH�C��� HQ2M�,#+&���eʫ�O[���e�F-x/Nd�f��ǻl�}��a��b���6E�)\/`�oj�d���S.��7f�%,I�5A�̰��7n䬎������N�o����;����5ŝ��4De:tZ���L��B�[�-�f��=��_
��o�i�(����R�)n-�5�bѢ��[oYb���f�<1�	j�OVPǜz�VS��`���ҁ�)����;%4F���,�9�܇!9��큱�Db��Э�X�b��#j�&������;:Ǌ�|ڳ5�n����5O
���8V& �)[6����1ժ�{kr%g�b;���^�pTk$���)*�%���aК��i��І����:Yi�T������a��k[y.M��"�H���2�I��f�6��@��Ye����`SV�������z��#x̎��2�v��\���&�[5�8!�CZ�q$ƺ�F�7릒��D[�{K�N�%(�3
��9U�̔�Jb��v+a4,�˒ķ`���(P�c��i��bC�D��22�n�q����4��m��e�Ò7/*��X�^fu�o4�Of�e��O
�F�� .���َ��6�P�7Rw����%�G6�J'Z�Yu��-S���D���KWaky�Vrxr�2�PaQR-��eM|���ҵW3$���ƞ�;$Y�	*�0�Hn��Z�2
zt�K�o�F�a��&�[ff�1�%X��%\F�Z1q6�汵o��K ��ݤ0�Љm��1"(hz³�x�J��Zݧ#�ETpm��x�}��8��#E�62��ܸp��(���$f�j�w	�7�V�kDˬ�:�����4�%�R(�̻����"X��'	�t㛹F�dI��;�Cfb��]�D�mCϗ)�^U�T-�:�:Cm�<M�����Π[���iCJ� ��V4	xqZ�k�2�����D��8�Du�K�������YvIto/oI���`��\ƅ�X��a�Vm���/,;U5����KB��k�£.��:�u�'GI�
��'��1���0��N<Ӈi�� �g��z��� #����a����=��Uw.@                                                                                                                 �                                     &@����*�u$�!KeCƔO@�Qr��	{Y���A��!OvnզX�Z���*���B��l�
�VV�2�����Uj<�v^5�90o�l�I[$�N��};%�\��X�W��*�\�h{��4E��3�[yX3�p<*sA�ܬd)�v��b�p����5����F�N���`��9R�Jl�7�����o.�8��w{�Q:�JI�/p��×_5F��|�<��Y��r�;��ѲpVh�J�.��𫎆̚��w�lkbA�����oTZ씆d��}�f^�SN��i6��
2�<�k�4�X��o�j�1�C�{�����l�&R�ҙ$>�	�5k�ҳ\����':f��<ټ�@�u���5�'_T��3j,��*QB���kj� ��QX)f��	�+9QՎ����ބ�.�=�����&ӹ�\\(��sEG^f�Q���.� _��`�P�v@�a=RMk/2�5H��Q�T�%�U������vߖ�-ö�����vq�(�k�Xڇ;U��E�#���SM��*p��ꩻG��O*
�XY�ɚ��&����SP�����5�Y{��]�TiQ�2)����y�m]ℑR�h;;:b�eT����ǭ����(Z�9ʋ�.E�ЕnڎV�ip�C0��|�:�:�;b�o:0ҴFYɊ��%f�#�i��n��gW r����*�g�sn�mJ �3g+�۱nE�Z+0J,Nw���"��S������`�[2�f@
Π��ӣ%G�맹��=�Qer�e��:4��ף�xc0j��ۢv���w�i�f�Z��������jj\�)D�M�Sv�'ecj��m���J����6kP����#b�r�JQD<^�Ք%iۘk2���B�Ŝ2m�<g1q���V�5n<�J�
�G�`%:WZ,@+��Pj�Wxѫ��֌�v]�kd�1�ůIhA�z�@���f���Vr�d����0�!��C-��T���%Pl���b�c­ҽ1��]%u��0�<�E�;z�,M�Ir��`�9�W"�q]����F���c�+��'bR�Py䖵��]Ayb�u�io"�@qa���Aua�{��:՗���-����9�K������ʼ	���Y/ɣ��ր�6LWݷ���GN3�����':^�2�$����yt]�Z�nB�>���U�2���\0.�@:���\ӽR��.`4>[o���ǸV�4�K'G	t2&V��ꀪL)���Nc�.t��Ǎ]���=�@�T]n���b'.����òF';�����OE�Mp�$��,���iV��㤝Vxj�|�	��V�n������l)�)a��ttO	�Ff�/7��f1�[�p�U8�:u�����\��[4���h�y��I��X��-]}�t�Ԣ�i����5�S�:���֝vq��s+���E�n-�H�մD�l$��Rs���pd��l�iO�� $ɩ��4r�l�y��>�-;�m=u/��i7�5�·s"����4��w�n.�U/a]����GdV�ӜiQ�,[���՟<��y`̖�)�ُ�3J!g(���p�����9`��������,֐��	t�}�;_�����\+���j:��潷*YOm`Ȇr���*"`�+�o:�����#9r�K͌q42�@j��:W�
'�t��xyD0ˏC�\ G�ɸ�oUf�Z�42#`m[��t:B�������%�k5k:���7�!ҟ�/e`i0�:Ē�bV�A���P�E�X��P|��T�<x8q�Z�D�$b��T�"N�H��37e�V#-���N�ڑxƁ2.M������i���$�I��p�M��-s�=�b�_Z';�r��8� GSW��5ZoW#U�qTY���L�	��|�f���ڙ�bct��D��,t�N7��6G�N��m��,Ǭg2�vV��n'�Ad{�^C/T�2�����̗��i���nc�{���}3-:Y�D�mge��[:F�<r���B�?#���֏:S���e�AZ���X���=zq���X�B���Y�Vd=z�an������z4�n�h|d��Y��k�Hf�ovл]
��JF�sLP��$��]Av�R��:ú/PtQ��M�]�굟,d��]���"�j���<V+�xNݮ�OE�^�Dـ��ɕ6��kM�h8%���N�Ϡ�֋�b����'J�9{R�0�:oh�6�h��;����Q��R�R=w��n	��X��;(�6IDiŚIMڴ���?L�@�RYZ�y}ȼ=+���,����4�TZ��m�}�����ub.��;�_�Mf���ɹ\�
x�̼ޔ�v�7ca�L�|A{�U"y���mnlL�\�����8����2+
��h����j�wbcK㧞�u�6B������e����b��Q�#��ǋ(��u�����%{[��zJ�{a���1򣳉�KfVL��'U�ݴ��̋�;�l$���+��+�%��>�}�rC���.yp�o�S:�+cd�#����2�SPj���>�1v@�Wۚ�iզU�����嵼2Ow�2�նi�� ���Z5b�7W[��y[�K1��'wP�a��:w-�G@˓��/6��`عƹ��p��Mkpai̛u`l6��Z�����O(V��b&K�;;���$4�q�+Z�^���eakf�va�k�w�h�ť�Y��\�p��s��}�i�Q.L��
��gV@�}�Twus\Z锷a���;�Zz�P8U�I��f�Xi`/N��E��j��u!x�}���oo�Y�j��/x4op\���3u�Bj�����Ì57�W?�q�E}a\�Z
���z��g�lڮ���w�qe1���na���y��;�'t�,��dWd0�F��n�Gb�u��&��I�iz\RR�`ŲB�eX�8͢�u����]�`�]���e��G�ݴWae�2��vރg��h���o�����&��=�&��(t�ӄ|浜.��9
8�R�X��:�c�V-���u�-цX�{Ϲ�=�.����g-s7�k4as9	���]f(���H�B��Rd�4��DС��6�r�-�p7�U�8D����)���9Z��9�x��z�I�s��c�״u�8du	�s�)��l_;��{��RCq<j�=��M2뺈縹C��l;��e�a�K^bn���79���悈a�h���Fm^�'���έ����똂ر �3mZݙl�U�(�R����Y��f\ⱍ����wL��h�|@U��9�NDZ��9Y���پ�^���N�~l{vr'^c׃�x6Ukb�v8V�B�L�kZ����*�-�wt�׎�u�(r�k����0��?��z#�����Y�P�
��L�b�f�
Ի�J�2������Gf!�۫�9��n61����ؙ�iS�+9�Ȭ��}�;mt=��#���N�����T5��{q�\X��/�y��d�Ds݋ҹ�lVԱ��hB|fWJ/)q�hF6�ZX��o=��F1f���Q��]=[փwR;���p�/�h�p�r5�8�:�@���6�\#79�[V�0�ٻ�pGs97�W*Wr)���Ka���iKV���oJ�ĥ���PnF->�E�3P7ٙ�����Wk�IiԂB��(M�/� �\���7��0�x�r,��v].[7/GmkPXP�Ԭ���&��6ou'N�#�*�z�UǺ7���-f\V�/�C�fԨ��s��[��N)�4l՜V�zw1                   �     ;��M�:��:8�nyP �H@                 ?�����>?����G�����7v{jW�
����H�ܴܨ��{�����p( �~������;�π_�x�g��z�i*M
��]�����k����f��wv�fɾ������b$ݒ��	�B7SrΫ���֞��t����cؔ�J�f��\���ǧi+�)h��#K��|M�A��S�s׼M(���ӥ!궳P�X�
���$*��Zg+��F���dR�e��AV�F���Y�D̵mXd��J���u��.�O�T���N^]�n��2��]6�-�Ph!*�չ��N2=q�9��:]�*v��Y`�}�8L�4�Y�1��]iv�m؊�%���j�a3NV{�+�ݻ�usY�t����r���͕�+��t���'�ެ�q.$i�0�6Z�W�V�;wx���r��=		��[t��fԏ�e�3j3���S��5lZ��{Р��v�wP]�V0v�P"���[kP�|U�5Ҥe΃�����#M@/��1"UbVg�P�k�V>���� �7j���T��&л"��%]e�'��T��r�Tʔ��C���q+9B��潧A�A|���
+I�����\��ߝf���Rr�[������eH�]&)|s:J�EK�E�8�?�{�qf�{r���<��/K����%��N��� �k��0P=B#N��mojVsL��t�C�N�
8TJ��ō�˛tɳ��=��G(r3+A���L�^�2��v#�q�WB���3c�rO���4����1���*�ѓE�7��}���O6bt��TA�X�y�*�d�'ON��3z�gJw��(�#�YVN#u�㼔��m��U��\�=���ܔY�f>�r�4�{fVA�f١��ܤ�5{��y�fg1�xv�T�6���܀aj�?�y�m�;X�nU�ݶ�`�pfܙ@�g{��Z��Y�GWq}�U��a����]�w.�"
]��3���.*�㕊澺\b=0Á|oz���م�[Ϧ�����ԙ�l�)k��r��1��9�_��.�"�ꖛzh���[�P��w��E��Zni#>�D��#ʋ�ծ�ͼ�a�reoʟ#2R�.��]M����K�&��9�.���ڼ1Q�I#�g#�S�:V��Ɏ빞=���l���{��T�Ǵ����Y,�AY�,['"MC|� �-el�h�ˣv+gRː��<�Ur���nk�qY������灂CMm:@en��n�֬�ن���ݕ�*7hen�X�4��[֚5/mi�Q�X8�Mtr��'�#oF�;y��X�n�J���RǶ�Ҥ;t�'o�k*�D�j���6���
���6N��)����E7�]�f�խ���n��%&)-�=�v�v���4o��h>}N-��ԡ�f�<ͺF�J�7g��fV���8�u��|C��2�i���yrS�J��;sMX�b�.B�tM�Ò��R�q=��y^�?����.�*��q�ss���.=;ux�:�W);I��,\��O�fI�W�Ҍ7���.����G7G[�Мn���O2'0^�ܧ�r.����8��[WX�n�V��,,.�MJ��n��4�`��\�|$�X�:_S�%�E�I3�MϹe���jd"�+�%��$.b�d��;%��Uu3�#�4
b��\��@�T���]a��X�/Kʶ���ُ���(�v��/�4��2�GZ6
M1��m�9Cc��]��T�G7�Fp�N���Y�90��J�ʼ����h��:[�|z�ҷ���1:�^ӊ ��,s�=��3r��m!F��7�s1#�2����6��1cj�A�@�fm�f�)	��|�6��X��K�&�Z�]�ΑY�Fp9���]K�r��̻�
4��O�,�˘櫽/��X�J���P+7���,��CJHf�e�%0���ٍfȣ.��)p���4v�iYX	��4�	���K�e�Hn� I��W�:�q�k��4��k4�d#��廎�2�*���Ve`�h	#,�;�ɋ��):L�ib��,T
Y��k+�GA�d�UVC]�A�K}�B��[v�5�����ŶH i��&�f���6s��h3�fJ՘��S뒱N�9-�'���t��!��M�g���ZN֛��$�&O��Е���N.��hU�r�&ʽ\Hl=|p�m��.bv�.7��tvV�+ˢ֕9�G����IP��Q�b��p�#7+����{��WS��\AWQ�H�k6�<:>��e�6�.�+eK��8B�㦖�۽�ǔս� �etw�4l�8�[��R��h���X[���U{�/#��7�r'�
p�=؈�f͈أ��E:�%f�z��2���H�R��`�P�$��ˇ%Bx����7nM�f��o�wd��d�b�&cj��{5SR��1*��\�yF۬ܤx�i�B��˃Xv��R5��N�de���n��pgiu�`�w
��j��)p�0җV�c�'��1������?��ڮe�3n8�)�y(��R��WW*v�)V�8e�m������PK��4-P��m��)R�2M������qr�ɶC�
���wF��j����A��Y��㕷"�&�]���BnS���]�R:e�x��$ؼ���7����ӧ1ȶv����2YÈ9g*X#���,]j��i�=@"�@HK���C�t�惴�p���!)�X�h�RS/x��G�8n�p*yN[��U�_Fa��ʐ�q�ˬ6�2���w�a�k�`>�s\�Yw�^w5ӯ{D9��#����e�kE֭�p0T{t��/.t��h֋�׻����ᑆ���t�3&㇥ദ;�pKV�;���ؑoQ��[{��zڻ��+�ˬ��S��a�xh(m�A�ټ��U`\Me+���)*m��r�7�j�GD��,p��˖�P(.��O,�O$Z�����?5���C��^<˷d,�
1w�18��(�Ka]��.XԮ��nX�w�I͝��L�uuJseG;��M%]�v�y��s0�U��ަ�m�:No�FϚf^^Q"�Z%'�;��;��w]�ѷ�Sl��F��l�v�\��j�v�V����O���"*�+��K�gt�7��zI�#цM�+@��ך�,�R��7�J�d���d�*ٲ��3vB�=�H��g���7�M�E�׽��F��[Yu��آ���nM���0�t���xO�]-����,�3�K�K�>��\��*e���2n���L�na��/
3��R9�ϳ�8R寶�/6����Bnl�GD��j��5}؜&f0�8���|� �!������[ݸ�0�YՁs")�����ү{i�.��Z4�,�f���7��U%�$s08�h��hy�e��c�(idv�]�{s�`�d�B�WN��l){)::�tGJ�lPy��z�;۸S��Ɍj۸��)k7l�G�u'w�2Ig{��Y�{�Ht�H�z�ٕ����/o-%O^���zE8�=l̲ �-�0V.<:N?nf���Wr:bo�3Y=h�W��Q�\d�O"�D���*ZX�9C��C]���:;�������;Z�@�a�b�^a����t�����)���5r��tWmaݓ1YS.�Vm4��nVT��R��0[ �ǹV����OO7h�}"���=t)�3N��J�qP��R�&�u��<곻�GDu���m�U�IFm�����y^���H[�@�h��s^>Auv��3p��;[���>�L'����FeO�toT��؋m;�
���f�;ܟVî�u�ō��q�L�MsUayK�yXj��9��\�T�����2��M��on����,5wՀ�2��Q֥B���R�{hEy[�[6q��Y�9M�1U�YiUoC��!¯J���u:]U�4{e�\�^KY/�f:����l%���*;��k�绪v�Xn
f�s�ͦ��!���J�f_�7���������UA"���ښ�-�:C��f�	�k�Ǿ}���            	ɱtV8Z��@�̎�C�B�6���� �8�c��u��6��c-�6�M��+l�%�hoan�:��d�V���E�V��F�kHB�Y&R�gŀ��Ɵxoس*�FbApV��z.V*Q�F>��{;|�r��"_(�"ȬbR�';�t<����(�ݳ�0M���כN�{�`+A-���{ԣ}Kc���	�3��Lq��oM��R�_=�,Zi�)<������|8�K�]��jWW*-�3�5�E-��(�K���)u��T����ܮ|��ȲT��_l��_R�ͦ�X�����Q���~�wSU���yBt�������n�w]��v��q�>���:ug-G�}H.����	����p-��.��k+pL��N�45w^)�*نQ�o��  � ��g빏��?4�@'���H��@Ҕ	� �D<{�����u(^`� PHP4��KEj YD�QBU!ATyM	B4ҝ��=�>�H��a	�94�!��� d��@��P4�H4�!Z��u*R�=A��H��4!Œ4��@ʁ�y��
Z�=�3���<����H~���R,-���)�Vv++���]I�*���P��ot�����c������W0�:��C>��B���x�K��6q��w�^������/8N�+ټ'���\y\e3CbXr첢M�zrdt%뼹��7 f���&���.�o7we�W#W���'O/[R��7C{�m�+z�*�����	��\nZO~ˆF���gccA�����q���=Y	��Y3����`���:�d��+T5���"OBm����Sj|���յw���
���q�W�by.pGN��nxz�����J����sf!�/������4��4���!%���;Cr_j+� �r�aϛ_2Z�3�[�..�E�p��Ngj�5yj�.���h��F���6�zVW׽y���m3u���[W�^r�=>Qڕ��dde9-G�g Ün�{ؽպy��viV�e.��Rqo5W�l����u\��=ҹ\�}�a�yA����}B�^��k��|�޾�;�NO��f�VOw���t��ʗ^X��=��|��m㚸���?TH�	�}�77}�M��5��1=��{������%ܴa/*�8��w��y�WYwыЦ���? ���8;eJ�
�+�,��:�z���c^Lt��vy.�{�=��<�26l
��,p�_��Z^�f+0ܥ�wگQ5QW_l����N�Y��\ʽ�O��o���	row/-f���?z��M� 9������~υ��
^�/c���5�7۞���r��c�ޯ��G��xU�M�&$�{�5����r\�����e�hQ�4{f{�y*��󼻞�]Qz�*��֖���Pת5q��ya�Zq�r�I�6K�������s���u����\L_y��+���Z�$۪wͳX�^�Eb��J��괚��T���Rْ���{��ة�������7~�+��7��r���-����^�}��Z;H!��4O��E����\�;5��b�<$�C�g�I��1�7���Zs.r}]�s| �݉+fo��[��#��^>B�_)ԗ�@-ҥ�q��x�R/������=�H3<v��	��W:?r���֪���� �<��K7骎����F���[[�k�S���r ���%�(y96O��^���)��k5�[)�a���Q;�оK��4�6Tscމ,~�>��L���{}صsb����M�"��u��~9�R��RY�͇�^�dso#.�y�{�~�c׊���ߏos>���`_>��'7�٬�gظ�F�b97���~�/����p��װ�J�g����>�T6��A#G4��݊�{R���{��&l��q�o�3S/)k*a'XV�3sխ�{�^n�\i��lP<�<A��̹Z���Q��R�ݸ t�ꥻ��V����ɞ3G��,�N#_��|8GV�C��1�C���e�I��VO^����[I��5zrM���9�5㓴8��:����櫈�5}�ܒ�^xכ�"���v�OG�]SU�w�jw6c���F�Y���p�+�ELy�{w\�OڙFҘ���֞L==T���ʾl��i���}{�!�p��+U�\�f�� g�j٨!a��x��(�#yK��.+}u��۳�9��^������N3�v�ߥ^�=��Vg�1V���ܬk�N�$�k[@v�,u	���ɐa�����WS�������D��x�ۥzUv��q�N`XK�L|�d��0��m�y^j�t5.R$����<�e8������u��\f~�rTٺ����?,Vp����ei�������ůC��,^sW�߹��o=xB��|F�}Y׺�z���{`�˹�Tm�Eᒽ3���Fɭ�;��}cA�t�<U�����|���9'��M�ϓMk�w�]����t�Fy+�����Z��u\��Ufsh�
]lQ^���o�^u�Ӣ3�jb�ڞ��{q0�*�]��{>�O��w�������r,yO�М���p��5l�	�Sy��_En�����ǚ��Sl�+2�v� ��WSF�܏WŇd0�Xxd�{^̬'�.h��#r;T"mg�	8f�&4}+m�����Ӟ�sV���$����s�C�9g_٪경� qo���g���O��:�Kje��*�&׹���~UjeE���Tt*�Εލ�6O����;��.�l��qj��r�.r���;X�|�w<�V��e���E[H�:d�@�y�W?{���^!�o˵O�	A�/7�ݾ�ث�/3&��������L�����x{w�t�.6��TQ"l�b��Nl��r�{�W�G��ya�co����b��łl�Ub�.��ؔ]�"6�.����<ڱ��)j3���nrsG/f�XHyc)̸CZ�oc��ko�Y�r�@����w[]$X�V�O��'�Rj�I�J0��R�7}�y�FtϤhg���/n��q���}uN�ȟq9#2%s���Wk~-筞̞m�z���
�@kyX�����ߡ�oy��=v�t*p㾽���^p8n��%�OW�v4#���z�xs��f؛��>NA=��V��{o�U6�F�oFK���]��5�n<NuS}��ǂ�B�o���G)#\�����W��)�����~;��5͵1Po=���N���~�2w�y�͜w�q�4z�1ï�l9*WR������3��vC�q�n��d
�R�2|�˹%��\��	���G�=i7ʹ�f�Ӓ{��+W��m��v��j5yz1�'sނ�x�µ���� ŰL5���?9��ʖ�M�����5�<���sz�����GX�V�zw�x:�^K�i�pc5&�|߷jޞ�	�9���֢�K¡��=��M��6��$:=9�!?}[Q}�y#ܺ�m�j�Γ���wx��5�Sp9».y*PZ6H�_.^�K�����Ƒ�Ղ���y=�kCg��do�x��qZ,�k5�'7m�{�ǫ'�[/|v?q�;V.�Xb�wp��r}k�\�=���L����{��n43)������=��}��mr�BV5�����ؓG/s��OrR�
�r�-􌱲��� q�SҮ-o��2���m�0�k�{7��+ӵQӤTllv�뛬���};σ��z���>����q�A_Sˊ�\WU۸1�Ll{���m�G��Kn�j��Y]t4�\Yp��d���0߳;���d_�Қ���&��kH�k�E����qU���+_p�Sv�ɝ���[�ڍ�t�]j�q��L���M9	�Y5n:5W�_�tt����xc?}2yw#O*F�]v�룒�5������{w݈���e�ܺ�1t���G2���H}����5����8�~��?�:9��8��E���|ȡ���#n�}�a�,�|��]w_7�t�u��	I��^�b��4T�ݚ��nE����-�о
����(�"��PJ�f;�.4�c������z���6�P�����/���"mIB=�pPbZ�L����|��;�,�3�Z��83�<���\2����9�蜮�˟YYܚĪ�B�,=PhPU�c�/O)��S~�W�v)SӬ�{'$�]�bX3(3��g����ڮ(����J�Q*��[]��w���,l!V�Y���nY��䬥��s��+K��0��3��aӲ�YQϝ�1A	�E38�Y���D��kp��/��EUG�5�ti�~�r%W۴��۽�;A�[W�9�ܔ$�)����C�{���<e"]���3y�c�m�8C�n�i�ǽ�;+�b
������RF�zbo����e�>^�re��?�?}����            �J�q���#ӷ��B����\�L��&��lR�����☒�krpͮ�R��2C��KR���5p��ú��5hV(�)�������X�]�]W2N�g.��M�a�r�@�1P܌���IQ��XW5�v+���C:"���Z���4`�u�*��z����TO,ΌP�v�������c-ISv�XB�b��H�;�J��8�"B؁<������b⊥���]��iy�Pp����5���=4v.  ~���)2�R�������u�V�@W>�M��5�GU���6��SZ��i�#��\�Pbd��uWJճ5]vӴ�P���̋@�msUn�	DsWm�*�F�Sv�����ջӯ�\������Yǲ��    o{���;�A�� @�JC�ԃAM ��

~��CSHU �-"��MF@��� �d!T�G'̯-Q̩�*s!�Ps9-̉�̙SCHR�#@U(�5!�S!�r���p:�8$
�zκﯺ���.0Nζ���ꏦ_;mb�L�����7�PY���S���ʹ�����ek�K���ַ��;����M��?8������<�߽��Wx�_�y)�N�M�\��ЅO�^_�W�z�����o���ÌG��{_�B%\f�������}�r����K���!]^����:�b���{�|�
����8�����^織�	��}�@�ei^�P�/};���.�\sg��i>�׽?{m��7 U��~��f �]���~Z�q5v���wY�T׊v��8�;R�{�����e�Ͱ��9��]�?g*"�Z�|�V�ǹB�#��^����9�Xj�%�5�SXCBV�t�o
�X�w_�������V��l�bF�J֔����-�$�8��)���m�%��v�����u�<�/S�IF��T/��&����M�I��Wv��kM⮆�����^�}�g��qV�H���l�Or~���[�<�<%|����h�{BBN{�h��~��/��*���-_��rk��S;w=y�{��
��%��}�f%m�������|�'�7WW�S�${���J�ϹC����p~��W7�?s��T)�;�ٳ׵�?V��fw)?}�_���g~dg��
�}� ���ևߤQ���Uy���]o�t����N�:�B�����o$��oƷ+>/�G�12���ZA������'_��TB���ou�3��k���6���u�)QyБ�� 9��VZ��i�Ky��>��磌O4���/������ �OB[�}㜨/�Ø�]=s�U|�e�`�@�m:-=CB�s:��A�Y�Z)�a�o]��[��#�*.������A\��)���U���;�z��S�a�%����O�W���m�������a�UN�e+����y���5�=4���>�7^���ƌ�IrsޯUM��\�N�W�㻃5��ͧ{��{�dn�u�/�'KQZn�Y��\w����恴�����(�Fj����Tk��oo�G��I�A������~f�ny��rF^%΁*��.���������~͓ꖼw;�#Ÿ7eЋ7eC��|�����2� �������+��N�m��Z�]l�{�N��s������w{�g��w�j�ek�Q�V��M��[8�9�G�\c^����t[t�j�^{�s̅��P��!{e8�w�l�O���.�>Pn����<��9�����Cr����O�Ò���>��R;��::��P�����+�@{�F@�g�{�����g=�����2S����>�w'>{�(]=���!���^���ԩ�2�G�=��S�p�d��O��^{����>��w�+��Nd;���^�e�2W�4�� 8�KK�8����8�䦞08��.>㾹�M}���=}���G����(;�(�7)��`�����r�
G>irܯ����!I�]\N{�;�;����oϷ��bn�w!�j���>�p�@�>�>�C��`��y�/��@9��w���<���oߑ��C���W����Gu<Bu�{)��/}_`'3��<��t��n]ù%�_����Z�<��y<�rߚ��}h���K���PVA,D�<�>������bY��ҘKջ��y�f3]rl�5e�(��4�r��'������y��S�z�Gq���CY�ǳ��	��15)�{�����yrd����7/p��z�#�/���{瞝K�w��`����C�y�WP<G��Q�ة��7)�z=�w!F��{��;��s�c�:�}���u��w#���_%�_e���S�h �S�ԅ u�g��x��C��#���~{��ߣ�u!G��C�;�/�w'~c�~�����]�ܯY�#�'`u9 u#�s%|�q��ߜy����|�{�_�}!Hk��}���S�|��p��P�C��<�˾���x���f-)ԜeǞ>��>��>��~Cpw!�b'Q�+�ΰ<���7/���]����;�ܾ@s{#�^��y��C��z�Ϻ����|��u��c�)��/r�;��qS5���^�rf��_���y�]ș!��|�tk[������]F��P���d�b�'Xp�!'�˼Ol���'p��� qu�<����;��י��{���߻�܏0��x��� })����x)�xy&HR��GZ�w/q��'�H��e>7�G�o�~ߟ{���8��S�Xw#��)��)�=�z��vu�I��!�b�.���98¾�>����_����-�B�D��tQ��Z��p$���~��p�=��^26G}�x��k�3�wD�f3��y}dh\&nf��h*[yP�`�ރr���������w����~�!u�R���� Qܚ�r��@�|Ġܦ��r/p���5�/�0��ν�x�>㞻��W�{���e5:��>�ܧ�r2N|�JÜw	�'b��	C�
ߟ}���޷מ����s����?Hk0W�������G�8>�9�%9�=��w+��X{}�܅&s�]��=���s��������_~�ˉ^�x���� �>�6kc��ܦJy�΅�d�T�;���[߽w���
S�5'r�.�9��~}�B���.B�8���B�:���O$|�P���y��M�|�3�o�����C�>�P�A�yt��}/���C�w/g�/0�� `�Hk1�W���T׺�W=�����~����'0w�n\�=ø;�!z��~����p�/���Np^$5�#��S��C^��u�6qs���~��}�~� �\g�}q�r{!O0��u�>J�'���H�+��;���ޕ>��}�}ϼu�={���<������
:����0S5��!���'��'=b�K�O��'��{�����7���]w��5�q����'1�h%8�ZW�O`�B�e�K���'��Ҟ���9��_$���}�z���x�g��֯�.>�5��o�rW̷��p�㨤�T�_w�9|�c�OxR�l����E��T�HT^����0(eb�S����rF��)�k���� P�k}��~o�? yj�� ?�'r�G]�M�2�x3܅+�>G>�� ��_�a:3pC���fg]o>�~���S�_!���G��=��
w�S {{�pd����C�1q��<����=o[���ߺߛ�R�n��.���!�.�����/q��x�K����⧇���.w�y'��w�����������������o0C�=��N���^m�αS�X}�>�5#��nSr�}�HR>��7�}����w����>;�}��Q���::��pps�WP<�A����qa��(7	�� ܾs�'�ߛ�z��>����t��K��C������`j��9���p�9ҧ\���=�ϾמkϺ�޾�ϒ�$}���]FH�Ϛ\���Z_n 2��u�S�Mb}h��>���=�(8י�;����}����}����9�4o�B��JO��� ܽ�8�N�iz�ј�J�{������>���=�=�׿w�ߠ�S�x/s'�� �x�!J{:��_%}�w�����r��x7Rf"}e�����ﯹ������G�>�!<�:��O.N�C�4}�OS�
S��e��}�:��<{��CŐ��o�;�M{΢���c�t	�ф��V�M���^��=�b.�wO�{f���W����?������g���N�o��RId�r�lZx���r�"v^b��L�C�ޙ�������S�������B�P�����T�`w)�}���;��O$��:��䏇�w/��u�N.��}��q�7�{�Ϻ�$>�- f�N#�Nǩ�{�n\w��P�S�
5�#ԛ���<�<���=�ޱw��}��κߟy�.����^n5ޅ4���d�q��f w���!�.��܅!�1;��Nad��w�wy���~���wnW�<���G��^.��T�xp�f'Q�P�A�Y��=��;�'��?y���ל��瞻�Ϸ�/�3�O`;��p܉�7R>^J�]�`���X�Ϙ4�Rk0O ܅+ԞO�U��[���x������:�)=��O �^�����MG7R>K���|��}}�<˽����u��u�_���.�mc�u׬������w�A�y���b��oay�W�k��pI����y����1�n��ߝ�e�l�DЍ�Zk �^��r����/�7Y���=�!����d�4ӳXD�3ǥ�Q��eoS��\ر�����O�s󟄢���_�S��Q�uu-��wKѧr�2��q2㙽�}�U�@iQq�=�����9盿ǧ�28��X�˲rav��.�E�k��u�����:���Wm5�_7M����i���^�5�{�6K��g����w�Jʛ�(h�.g�Y��X�41�ڲ�έG���2,w���=���Ҿ���z������G���*ܚ��R��d{c�r�'P��3{gmw��O�&,�N�~��+cӞX�}�}mrM��q{d`vw۞���v��3���M��u�J���{p���Uz�ƾ��e����vjsHG��DǄﳯ�Q=Z�k�p5�Y�Z�B�l��
���j��������gi���0�Nl�@�8��&cP^��\M䨞��� �¢P��(�
ҩH%�J�J!BR��EQE�DS�~���ڭ��˯�<\�ȉ\��мZ�
&g9�%�ː���L�潯(�؜=���߷K����t�3���~�$��}k<4� 3�"$�-Q���w(����`�0Y삠~����n�+�Mh�q�8yҺ�~6�Ux�סT�����$�ɏw�X�&�ڷ�yw���͉����G5u��$2�i?�|V\�.�4����&��fR���k����0���=�
�k��δ�yY��Oӹ=�/u{���EPs�Z�F�}/9��F�ʂ�$8�f��*Tл���M32m�ZN��upX���k�
�������k�*]����q=�/��;��m�}�R��C.m��αټH<J�J�+��)��+��J52fc˸v���q��[B���ͽ;���[��B^�"���|w,V��b��w�9񽵈�5��+5`\�Z��P^*9\��X_�jc�U���ܮ��n�E}��'�ڜ�yݷu"�e���z�<S�h]Ϩ�\�WV��+���z4Ӧ��A�O��Y1)L�jS�r��;l�#����Y}�T��_2B�=u�X�^��9B�S��]�C6��i��&���eЭp����'�[��u�f��Mv8-c���t9��-#.��]�\�Pa�T��:Z�r��R���z�`��P��ک�y�7W�������߀           Nt�"��y�.�j���Ka��J;�4�p©��淜�L�-�O���X�G��R�KL�&4�ô7k�>�UVAnѕ��*�ES5s�;���2��t�n�!�m��[�p���\�Aem�S�n����۫���\��ו�VsɆ���Ww��]��L��7t&�Ɵm����V�/����`ȝƮ3p�5i��~�:fJ�v�Se��6��4\=R^ڥ9�����vC͓���m��[$�-���q��s��B��4�>�>Ӥ��/BF����,���\�^L����(Ɓ�vs��5�,^�x��c&)+Pq�֠�c��k�k�<&�s�O�'7Wb�Sr�+� ��:}���lq�%��9��]p��í,�JNw�9�B��=���    ����}��LD~� /�� \���#* �)���MBj2���(�@)��J�?jVS��� ~ 2JB�R�9
�Q�-B�/.@�(q�%�F�\����(NdrR.A�NAY�-U"d��R��"ҥB��c!�i���*�u�������ė�ff�u%Ht���N8�Nn�Dn\Hs��ݏ�j�W�U}_UU/y���O���q�����B?:�߶9�??0���3���&R�K��d��'��e��Izq��9V}]N�qm��.��Na5�i���O"Eu[&C��_T�GA���Zhl�w���1�����Z�T'��6�{[~�R�R�y~v��s�;���v�R�K��zM��^�����>��a|wʲ�d���h⻱O�����^�9���-�E��^�����j�=X3�=	v�wv���SH���y�NEU���S/�o�{?���2�P��sU�:�ۙ���84ݎ�GGK�F`�2�.�&"o�gZ����9Re��ǽe�5z��]�렎�uI���ͬ��DG��M������P�!״�h�g��o���!��׵��йdj���W��Ɲ��L��b�}Uv�:��(ϸ���O7���ʹ��)&�l�k���F��b�t\[f�O�O�Ԟ�e/��k}�j����ӗ�!�r�4u�Q~^}�����$��F,���g��5`U���l]{+�7���1�ď� �t��[����q���gw�מ�OuM�Y���ܬ���[�.�3�\�p�~�O7�ӗ�=>ۖ#}��z�
rt�s�$\�sPGx��G�=�a�̦�m�w6��c<�Z9�~��b��OS�U��Ϛ�e�QoA��:��+�N�
���*�O����W�UUU-�^����#�;�����~[�բ˫��絇>��v����r��k��k�/�S��Cvx��z2}E��;HK�u���X���l�q5�z�F����w�7Y��O:�/�VƟ��z�OJ�:���W�v�U�G+�f�ǖ\vm����WB��\`{_�N=
�Ø�{u��^��w��������</�O��i�G�\����tͬ���Oz��;=�N9vS���=f���>J{���0�B����['n�/`ṓM=Nō)ם�쾹�M�Vl;�EE��l�7��cG�]���=W���6{�"�;�٣����kՎG,o��/Ҿe�ha۵�y>�">��ִ6L7}o�y�x~��R]�W���y���
�{�g'���/FN߭yZ��c������Щ{�~��l���V�<�l�-��y�R��5��{�x���[�>ECt/��zS^١eޑ�S��A�aK���o+߃���;����/��=3���W>B�E�1�]����䤈{)���Gp�N]W::�a�<*{�o7���~��ٵ�2�HkIT��f'w%�j��Cl}$�/��Z�������}����Ss����퇏��ܾ7Ѳo�7�\m�ӽ���ʐ�YM�xa$R��><ԭ6*5DԚ�M�p�AE�̮�Q��1���qH�'L��}��}���rmB��g�DյG;���t�3��׽��[�$/o8)0�Y�ӑ�^�Eɫ����*}��V��=Y+}���ó(��rg����Y��gVdۜE�wC|7�-�S}��^گ�>O���y>'�grd&��UoT^������Ǳ������,7�i���=�P�U�{:*s����h��>����S�C�K�FH�*�Lc.y)�w:c�$. ]��ہ���ozv����0���-�a��^�n{�Ҹ[fF��CyG�]����f�v2��A(6����b���.�q%�o�k	=D��9��og^1�Vk��mM'�Ѽ�3hAr�j.v����<w��<q��Z����>����CM��<����Ϧ�=�th�Xi�����7��M�)��+}^��[��[�-[��S�ܚ>�jj4*�:~�M���΃"�d[�Ϥݠ�{3���uEw��md�����Ӊ�Bw��JgN���km�>��{���/EoN��Si�c.���~c��o<�Nn{���IcUt�އG.�O����ڑ��{����f����t�&�X2�6��-u<'*�7�Z�"�yl�}�j�n�aW�<�WDsM)E������M/z����o+>h�<��.X�TC�ޭ�g%���\�.8��^Pȯk_j�͌hD�w�2Y6T�5����.V��sz��U_}_Qֹ�=5��onF�<�.
u(��{��f�h5��9;��LG�����q��Za�TB�5���ԟV�G)V���i,^���npBgl��YǾ�Ĩ���ݻ�/������w�<�Ǣ�L�|B�d�6���}��'��t��;bn,5~[ϟ��S���zc�r*��<�.1���Y����fP>��`������W�3�,���"��j5���.�B�^��k�"���bo���m�Q�ؕ��V٬u���T.��h/!���-w����r�y{�c#M���HBr�K=�6�D��8��6Z]C�<k֯v`�9Z�q�#75""�[c��ǖ�])���>���ƛd���V/E{������H�3p�չ��n���sՙˆ��w�����~;��Z�P����pz�2{\[��\�z��wbW9$�i��S^�ɥR�o=c�͕�ӕ~�o�{i��<��1Y펽�ao�׸��ͷ�5ŗ�{
Y��z�p��m��V�u7c9�.n��9�ʯ{#̥5U�ޡ-�F��o�Ի=�{"S�¶MhxF��U���u5�f�Hk\�V��zS^��׼�>��ݷG����f�0iV���?����q2�z`�O:H�!vlwat���y^��#%���Tuc34Ֆ���
��nc�u(������/k/�3�s��{û+���t����������M����٭ߕ��s<����6Q�d�2G��ff���պ/��/ݭV{�������a�>¨��pүZ�{��[�i5�p���?�o�������\�T>ƣ7�F{�wO1��:u:}��;�*M�_��}�LR�7+�}ιtbf��ۥVfsI]�����p��u]C�G��ڃME�����qŉ�o��<�QW��b/�&ՙN��ٱJG^Ճ�^�����ʷu8���I7�FҲ���Q�oH�sV�=�n�xZ�]/'e�d����@�D��߷��-Ww#y�P-�(�}y��x���%]5J�h��N��;!F�\|l��,�+ 4D��G舏��~��g~�hw\i)�X*�Eڡ���%�'������[�k�sFH�vD�����ֻ�@���y�Z�;�`dj�/�x�jL����Oߨ~�>N�ĭ�}w���v��?b~��߱w^��5����MzM��^�Z�i�7����EＭ�lH�ֳ�}��<�^M�'>���<��G�2�5����� wWE���]?u���� \uަi�Jv�3�}��}^�����둲��&97����5xr�K����tU2�1yվ���l	�����
��Ц�cv�ްk��2͗	������n��(l0_f�q��8��Ѿ�kp�վW������bP��TxՌ Ɛ��1]1e��	&���=Αa5F�I7���w��-��8o�����ɑ0|+����=��.nag��v=��;R��#Fp��̣�&m��g��œ�X��U
��hv��Ǡ��[f�XHCdokm6T7k�@2.��"�Wc@&�ly����f�3W]h/�W.K��F����6��i��mK�x7��M1��ծnvs�+�V�ؚr�Fe���ݗ������\�Z�f5�(n�W�dq�$>n����l��eZD�d�Z^)��92�jk��)�֡�%�X�
<x:s�g�{gWaV���ZLm[�(��L��J�,0���t#[�66��O*舍𛺠�"��Ȥ�l_tt�����Z�s`            �A~Eƒ�.��L�Y�ê�̽�o3#!�ז�BT,��@�{��#ٙw;/�0rjTˠrmkW�V�@ǂd�'6'#B��<��
$�����w���+`���̄U�6h3�����Z�vCm�&=F�[��#�v�"V	���տF��OJe_jUn�@��8=�M����5�$4m��j+�H.xZ�BK��J;�pM�J�nY%�z���<��ȇ�y���KD����S�a���5%��s;���j�m�X	KNiw�IU�0����M�0Wә���r�
o��e�{A��[�Q���2Qu��ϡ��]�ݩra���N�|�s],�T{�x�u�+���*��ɮ�*�x�������IWǨ̅��{+=� � ���%N$�B��(��Ƈ�rJ��y�P�4	HP�d?J��e(�bLP�KOrd(u�%�(�{�2S��) x���
�Zj�3XcB��-U!�KT4�E D<��%4W2�KKIUA2��W�|��ӛ�Na�喯�5	��)��t��}Ʈ��7�o+1MyV\�f��5_G��v�k���	��}>��=���� �Gu���5�rl�V9u����g��U��� ��̞��{�D|�`�Օ6]o+�j��Yl�yI����ô(�G.��Vw�X��0�%Ɍ9���O�αd��=q�S��e�D����P�y��~/t�:=9�*�.}��[m&��^�L��ڳR}��EQ��[��*��NK�s΍��vZ�����j=︃����'u��K�_l��GkF�L�n.�#{zw��ҩ�^雰-[�g���J:��Q�f+�Fv��lU��G�cd�L��R}���4��^�����\�^A���wBU��3�c87�ʸ7b�F�2�Wj��:�UW��Ss����!���!E8n�_�[�bwY��y�g�6�j��E�Lr��ڞ�{j�]�Y��Ę;����hn�L�:��%n�����x�l�Wj����$�{�!>�GX��k��6����v^[�U�m��2䢉7f�|	OG^\J-�����:�0�UkɃSO�M���_y�`[Ќ���)�id���v8ڼ{��_m�N^;��V�a��qy�t_�l����e�v:^�"kR��]�ɇl{͖�z7Cmg'q�n\���i�Ev}p����xSY�,NT�Y��
~Z�q�/���ݻ�KAׇV5N]N4�2�C�]��_@�~�I�$.5W�����D{<6�k�	��=_��X�������/�??O8�߅i��/�;�{04�����[�?E���w���2��N=2ׇn��9?zq\�������FS
�����E�f�ꕣ�a�6�&xVu�*KV���٪��[�5:��7l�=Q"rreb뛽��M�?�˹|�/j3ݐ{삙��I�۝��� %�=.+���y<X�����"^rC���Q�"϶
��{�|�W�6�+�y03�9�u6j�?V'Sϲ�>��7��<�&��Y}�T�2�����ݧ��m𭚗m�u��Oj������ܷ�|�b�p�j���}Lܬ⌶��%N�kN��UU_9����~G�1��Ҷ���v��Qy_�S{����������Wq�@X��P��Z3%����ȿ%^_'�	ϕ��b�Bw�s����F�B�$���~X��O4o�=u�v�u��I傫_��)9zH׻Sk�L��Gt(Uk�ڲ�Z^q���٭����Ǽy���¯S�~��gt��3�5ޗ��c������<+�y��@�=�ξY����lxVfnֺ}Y�G� .i��D��h01L_��5�B]=����H�3������V��(��4�2м������v=^	nzdd��gi�=h��;�9�5!����R�j��k\�lQ��10��U�{�{�~��G�g��py�:�Ó������{i�=ꝯL5�&�5���6��W�P��)���{	��cƖٻ����}�e�=uPxz� L�WN��,�3b�����.zc��v1��tţ�����]S�X]"ņ+�r���I��fu���:��솪�7�hWuӬ��O�\>,G��w7��꿓���qfI�8`��Ƒ��0C�>ˁ�|)����ҘeeS��k��7�G�������{|�{�h򺂎ᝇ6隬4��utmu������_<�z����/z2��Ȱ���e��6���4�8�����؛���f�:~�sp	�-�k��y���v�Y�Y"��	z��#~�I%Gs��h!:��A�eֶ�����u��Ř��s�r.ǳZ�;���>�\�>�*��
X�]��f?�U}�{ɦ�������˸yJ'�0��J����٪�kp���Y�J���PC>'���+�uy��_�m�ܶ)F ���d>��ݑ"ɫ�����b=�
ф��X��}ή�%="��[Y^�C���� h�t�l��;U�kڞy{�[�֣�^�mf��⇅p#l����D��X���G��<ow���ދ+�B9����]�.� �#�H���[S�8���]�[<��b�.
�ߪ%��w�d�.�TqU��_��鸔�HDd
���&�t�C^�`]3@��1u����;�s~x�Y>3�j��7�i��lL�{es��W�-�b	�^nȤ/g��Ŋ�5zxM��]�ж�����=�,Dg�eu;��n�[��HEktMue�nr%hܳ�l_^4Vbu��璐��N�ń����s�N��ߪ����#nzH�֋R����b�{fIR�,�׶�2����j=��`U����`]��7�q�-Q�H?]���n��f[��w8����Jٌ�aO���^�R�?�����@o�� <;4�C���Q9�0�B�X�f/kv�����!��@��N���j+�
���b��;՞7��NQ�S%�g�(!�:M/ۖ�����ہ���{�OacB���^;�j�)�Wp
���<�����L�:��O>�1k{#"τ�����Hh�hW����9o�OҕA��eo���k;�\)��)�i��e��_���=鐀��<+î�NE�T��=].\��D��m\�띷4���BnԂ�Wg=Tfs�Z0��@Í��X:!�r�|,U�W0�� x�Y�7y�7�Z�JtG$z*Y���uq��%�O���>�z1��џ�f�8epU�\+��Z;�N�U޿>����M>MwK��L*��4N�g�2a�Z���ͣMZ�:%��xeS,]2�?k�=U~ Q��AX)�&1��qw��:�����F�R���#LZCr��;�	Cԕ�������L�g�V���a#��4V"C<�X�3�ܽ����sŌ&�0S�Hx��&�B�����[�=�g��WU^Th7��_x՜>��U,��z��8�����r:�X�W�*���@��-�S�3��y�i7=�46{a5{�i��@�OƱ�b��O��a�#�ow�{�.F[�Tl��*¸4����4h��)�г׻3���"��|��lL��k(Q�V:]'���t�(q\X2E�A���
�L:��앮�7���طs��l���X���!݃������4���e��a��o��!�r��^�����iu����w�aa"��8Wf�͚�:�7�����r�z�\:r�"���}t��{o	�ӖP�wW����W���/j��2��� &`d��[t�49�Yu�q���%���&iک�R��h�;��B��b^f@��@�H��ܝ�^�|��6�V��b�C�#M�A:�YW�ѽ��O�n��8�s����tX��y�3O�9n��rw��G5sίyѦ��W�;�X��T����Z�u�Q3����]S�X Ū�M�{��ނ�s J^+�}2���5�z\���fB��^�'z��R�ԙ�}��u��c8����L��[��%�u����Fk_��``܇�6/!��r���Zˮ�N=��nK�2���ڰ�'$/�("���4;���1`�Њ� ���HXu���}A�!��c�u���>F���0b?�i��.��C'\�1��~��Fy�AW�u�5��X���t,�s{=6����y�7�p`{m	��c��y,a��RB��tq>>������<�Ez��� l�����x�,���7�נ��m�9�� ���];˔,W��+Kg7�)�G�7
����uo�bH~��]��\H�D�}�}�(|-5S"�h�Cٻ$m٩ZW�3L�>'�
O$��F[
��N�����97n�}쩹}�
l�� ��E
m۪%�Nf�#���փ|K�w���K�X�,As&��`W�#[�ovG���0����#M꿯�|+�]���ba� � o�K�}�t3�8>z�����J0�5��J'[r��亍?h���M��Q�Mh���)EV�u._"jvm�mǜg�q�����N�֎�����MG��^�֯Nl����sYvz|�x��"w�����K��̎p�p�%"�9�wNmc�X�kxq�^-��k<k�=v]��,syo��8�f�t.�7�$��e��;5���ʵ��C����"�5�#2��x�}k��u*�2�S�#^��k�s3���v^4�'Bk諞(_��J=�[���i��˺�T�6�q��Q���tG��*CW�%1���6�zC��;�׭�d�|Y�Ӭ�$�K��R��]�l���@��d��a�u`�r�\�YY���J"d[�k�e�iep�w��k,���2%���"g0�R|&�"��tBy�.��B49QGwG�ʭ�$6            �Vpe�v�ݪz�K��w���䶥��\�IJ���9[V��7K4��qWl5����q��ؕwl=CiZ��q�G3GC����D,�}�u�f`WA۷E�}l��+&�i}��7���)"�.�]���_�ȼ��	w�eJ,�goBM�̶{��Y��%�o��C�o:a٩;TG`��ޑ�["-Z�=W3%9L٠\���/kmA�n'���oBh[��Dڤ؇W7D�C:�B�Q�����*VeK�hH�il�чǓG��g�i�ۙ��oTT�#�PJ�����^m�
��C��w9#�W�K񻵠����sʹy�!�)̡��Z��1�3"��`���N(�S�GY�Ru�YH^�5��t^[�$��T�98��p���n�x   �c������Ǩ23��&
G�2[xd'���sEP�-d�Z���ƒ���8�`5;�0���j��r))���3QN��Uܧz�;���b�"���"�i�;��"�8����b`�j+�*�����*h�rh"?�q�~g�q�us��fw�~���"��#ZiڅD[˹EQ�p��P�Li��_�A���of=?�UzV����].V<oMx��x�����麢�0u?��
B�A�z"MR��߮�7d�f��ۦ,.y����d`x��/��P���N��Ъ2�v�:�N�����Ni�1���_�.Z��NS5�c8���B�����u����{���X�P���օU��ܿ����@��]yu3�k��OK�XJ's�k�_g���xSu�H]
�F���s��\}D��Z5�~�w��[�c��v3mO�p豤�/-�JO���O�"2���H���5���X��@�b5�� ��Щލ6y���.�'袯
�k!~*�� ` 0�#Ɯ����C>����{YO�S�=���+�lwxt�/�+�;�i���Bl[��˖��7ϥZ@h.GX�e��ն[���\���޴�P�e'���F{���X=C�s��Y��%o]V����K3��p�X�4kS�.�����s��z)Z��nb���-���
�B��/zI��Hߥ�
���V���W�m���L]B��˫L�7���ɾۯv �^:+��&/E\��=Jy׮�nK%�K�a�Q�Na��R�c�
�`B�;#-";E�`�S"mn��#��*<4��VeW(郟��4�;���Y%�����g}J�qB�d	B�]�i�>�E^/d����ޮ��k���HPG���k��� U˭i�[˯iQ��=��s���~�_��Ͳ<���T<*�i�Y)W������{������eM�/|p�� ��ʃ�5[tǉ��	ziF���"�6��v�_G�s���j�o��D��V.���MoW��*�������p���[;�K�ԊwLՕ!���47�G�N0��?}�?I�S�<��n�U3^��˦p����vT������W{�l[{_{h�7Q덼*�6s��h�J�[�5������\'�9��c��3�٥;4A���72
�������^���-����.0G�8X�s���әPj�a-uW�����ɂ\]�{>�&o��I^v�
ެ��y��!e�W��{��{�$����H>$P��t����5{��V�Ӻ�=�[�]B�Y�/TU����⇆,U�u3�K�`U��,_9��.�5�bsϮχ��~��Na �|5�<<��p1(pYt�ϖ�h��H�%_�]<�ke�*ٮd
�
T�f�nI�jԵ��>%6\l��lT�E�)NUҠ�햏�%,�����0
��EGl���(���%+�o�wG����������T��0;k�R��ު���<���]���nvB�enhQS�{ӋI��9�S��~����Ʋ]s<>�t`@��.��K����&�S9���5�r�X�w[�9���G{���i��!��\��ٖ8xR���v��G<kv�4��C[�;��׫��� A^z�l��G��!�qb��UǄ��Mc�������͙�~���u���J����0!T�a��/��鶧�=�$��i!��PQ���ßu�ˢN�����6��;�^izJ�^�՞\PP�R���F/��H];3O<3�z��e{i�F�2�S3�[�>�s���|�s��;�)��8���r�qEԹ%��];˔/�^
�[��":�������Uz����  � ��HnB�����/��{j�[��+�l�N���W1J�]hiε��%�1atX��(.�i�&���ӊ���T�{�ENT�ݬ�a9�$�WQ�ͨ�����-9���+<�1��5����'��Ѣ��[>��ϯ�N�=��oH���ݺ0~��������f��@���N~�����M�Ɠᐡ�^�զ�-
@��,L0Ab
)��_[f眞�������4����
�%��ba� �/E�����*��H��̮ް�֚�5��3�I��R��Ӽ����i�*��X,0�e]���[P�k$�(o�˞��?{Z~����2!�&��0�V�ں��Y�aa�a%���^��v��D�#��[s/��~��I��c;�(����Vٸ���>(x�Xl����և��[���5���N�}��q���°�4V�8��v0gKc)���*E���-{�c9�N��^�E�)�g�\�>��r�ޱM��A:a�NڹM�sw��)&�˾�zL��&4��bA�@;˞es��6S�6�����*�=�{���m1ЀƓ��6�����u{w()���{ݗ�nh8��ߦ��Wpyx�4��1��!�z�zvT�##M���>F��#��a:J�ŕh=˥��#4��n󰽽���a�ğ���VW�o�V�B�00 0�t�!��t#��ܽ%�9+4���nEJ�gYw�D�44V 4C���\��fOu}ꈊ5~3��~:<�
�� ����?@�#J�&�ސ����H]L՞Gh�����L]W���캱\}oխ���\7ƣ$X�>c��W�i���"�P��ׁ���F��6�x��ѧ,R�`C�W�]���pwYcMh��{�2%�nzqWu�`W��fB:W�<�`�.׻���nnʲ8�E��A`�f���Pu>�YW��tT��1Q���}��XhN�u��YѥN����[)!���lB��u�X��|�t��?�To����%��W@����0tk&[�ok.�<ٕ���l��Ld�9��(o[o�o���HS�.�d�|�3����~����|sO�������I�2�\]��ޙ벆a��^{��/Y��<Mw�^��)�<M\,�:>������zgu�c:4i3xt4�⇃��E��uxm[�$���ٛlT���L�@Ъ�ͥj��ۃq[�@�1��?Iv��V��E�5=n_�v_��B����'O2wg��irfd��s7��M�-C��'�3��;'.���`#s�3˓��xp���^F <<=�	��/��_C^_u�!��Q�����,�Pa�P4��$P��@h�O
u{��������{�����:"����{�04��}qrZ9��Y�y<?z��m��%z\z��V��B�I�o*[]�>�\��r-w�zk%hQ9��P���f4���g�wWT��L��Pc(�b����F��&�N}e�2��ؓkފ*��φ�s�^��"� L�2`�L�8K�����;��@3����ӵ��b��d
U�X��́YY�9��&ߣBǴ�wƟ���Ab
BS�t�,-�z&2�?Y�z�3v�.�y~�>U�atM��*�:j ;�B�v�����?;��5�xx]��C�;�@8h��x`����+en����<�*��:��4��e=w�k4�C]nK�\����h��P��l�ׅQ�^ζ.�o'6�I]5:������̈́�֮=q֨U�����s���Ӥ��S���@��b������ǆ:i!�5�w��0���V�s/��x����#x�*�f]�g0�q�\�Y��	�{���T0���(p 	sn���e���y�if<��/# ��^���7(&4T��U�M�M�-���W�>{ؚm������f!� �И��1˭F*�*�v�=���G�iz�� T��ub �Dz��m�(�+]ǻr��'��rq�)�
��9|<���iG�^�;ݴ�7�Q���d�o��S�?8k!0 �(1��~$2i
U�o�x�Ǭ�E�|�r}�w]ꬷ�X����ut�ȴa<0�&�ؐuy`�nw���E %��VA��yƷ�k�ZkMR���=5u�/|����=��C+}lb�Z����������APW��v�=��Ɉ�A����u^�#N��׌��c<lL4�bXFy^��&�p�@�+G��˱[��Iや/޺�`��+]���֤z	�^J
=���C�킓T����S�wu{=QV[�Ez�l3�%w˪�(Z�Ȇ�U�7{8�����:po�W4�x�mp���[3n����PDA�'dT{Eʾ�|�s�֧��1����(6녲�+,� xC.�M@G�	�[[�D�OT��0����
�e��ƽ$�Ƴ�w����5�'���C�½gB~Ã��Z ;4�9���t�kW��ɱ�n�����QD�B���V�	,�v�R��GU����<�]`� 1��G� ���&�e�I���f�?=�'��O- �E� �޾KO�:�S��~z���i��bE
�TwVMp�t�2����.��>~���V���A��Uf��+p�#J�Y h�!���t@�>��.�����\�`�f��>� xMT�Z㬮�ON�-����u0뭺�����Z��n\�\-����YW4�=��g��Y���`uD �c�֞�cLu����2�E����q�1(w
@5����w̥�2�]gT�����v��j���3�/�-���&("��f���A̛�t��Z�e��l�ГBIk��M̙y���s/��J����g��q��E��7������gr�ZR�a$�y��e<笲�Τ����qB��ە��Mq�w%7kb���ь�i��_}{����"|�<Ͷc��)Т7�++o�T�@�3soty�fq�e-�p��1݁2�g�a�p�ɘ>a�"yf�v13�YңfL�Âޒ�9VzR�TnZ�Kn��V�ގ�jŢ��9�7�hYu�8�w�Ze4�@&m>�[{���E�mb1�q:���Wxl�wk%͡�c��*H�u�+N(�SG�V���;&s:��R�
�x+ْ(_NV#{���4�             �
+�!y�}��֚��<��K��^�y��sՀf���»�lve-t��eFL*�jz�U�՛�(q6�UӃ]K��\���7�Vk:�L�#��CR�9��;\��K���2�<���A8V[�-,t���
=O�h� �)�.��D���N�Qy�j�*�X8=��Z�!�'L(S�v����,+���L.�����P�u��2��0����5��[��V�{�-��ugE�k����^VnKm7�h9ɳz���%Sb��ЕvW3��90n�]h�����J�M�n��̨�*y�[��݈J�r��KX������jG��>�šN�JQ��s�M�����9��S��{@����b��A��U�'�^r��Fe_q��ݿ��]� H ����QD��fMSEQIUL�9�{&T-sIMUU'��P�ˑO3�AE.s���C:��z���9!�E�泉'��`r!�.`˘q�ŐQKLT�M�6u��
����5'<`��0�*(��^�9�_�뿾��-n�~��<gg\��y���Ê�{�T\k/.�98��R5	Tx��� ��m�Sʪ��=��9Z�^���*���]h����,�s�k!I�7�.9�L�;&�L׎r��u���k�Bg>[֗����64�|)���)d1�e�U��W�VX�I�><}�!�ͥ$cO�E�� �7�X����`WP�U�C���gw�=�y:I
Ã�-����	�%�F�ن���q>5�V٘�?y�n�W��]��,��W���
(��{�W%�d�aN�O�lE��TԙQ��K��W3k,��>��sb>V�29�
�}�,g]׆�kn��]�W��A���$`|��:� ��t��;J�k"6���N�\�3bg�n���C�g�\5�l}Hm��8��v���������B��1
t�*���:��}F���Y�>���wJ��U��#�3\T�F�Y��+gFu[ba�u�4y��ol��MVp���S�;O�UP��0�L~�ng=}0*�ԟ��Ә�����*x��V���8�t�B�/�J޺�9lgK�v��neA"ʈ�g��R1+�,} ۻ�*�ڦ`�I8�ʟm%PB��s܋Ag��N��^R�Y�0z�!:�O����/�ue��֐����x�3~�h�	�:�>(0(1[�ύ/m�5�nψVc��M�]��W�����?a |��2`�`7bԍ�zIS��f����-a��f��+�  Ǭ{�/�$��&��z�Eu:0L��&T)�E�o�g�V�8�)�k�˿�/q���'�J1n� ��s������z���,�*��B��A�9 ����x!�}�^��h^+&6O=�@��\�sI</-���l����}�T}�)�3w�i&>}�����M�aI򜲕im��Q�M��S�|o5��: ~��A�B�> m/):��p��Tzra�/�+./ǚI��ݰ-D�ၲD^e׸��ׂ��5iF`�s̽��q�N�Ll>�X0�8}��d�����{��H<�
a�V\۰���z�<)3V:Q�q��{�4F���lh�y�<�ѡoaz��a����o����z_a�k¯޿�*�"2�����E�͍�e��5�Tp��b�#���p{r��4W��Cfz����K���tޯW\�T�j��X�P ?���U]��čD��q���˽=�s���>sr��aC�ӧvE�	ᄱf��)�/;}�'p�W_�h��������}Y}�<i���
*��׉;D�X������4P�vۮyڲ�s*���L7��&�2����&g^۽J��@v�D��ǌ��w1��R��+�#�OW�V��]Ǩ=����=��ڴ��w�%��pb�֭��xxpB��)2�&<�ݴ�?�Ɇm�M��/3)���=������axؓL�fwH���Z�=���)%�2�U��\�xޚ�Ư,q+9��K��il�%�RȈ�V)�5U�{u�����@�;�����q�z� �YĲ�� f�%���]3E�%l�-y��сj�5}nb�[��Nn�au�U�˸�+�����3������ӂuK�I��1�΅����bv�[��uh�|Mw��U���'];�v0et�3��
�e��K��ܗ�hb�Ռ�ġ��3F��NL�ګj��y��s�i��-��S�A�J, ��������ގ�c��lw}}Ջ��Ohܡ�3�VA�I,���{�w��e[q�N����Mx���|ȭ�Y'�8t�ك�EܠY`g4�۷Ӛ�1f��3�5'���O�y�kQϛ���������,��Wq���� {�u�C{�ko��n�i�$i+؝��g:��ĥ���El��v曬<93�j
γN�b����\.��������權���Ƕ��<=+�i>�
���ڱ�uQ�G��,R�T�z��UY�m���S�EM�h��D��7�6蛎.�`��Z
�
�T�v������MQzL���ᔍ��O
?X
�/¬�Q��$V[���"�a�1h�Z �fd@Q���j��=u��5�������r7�Hd$�����:0]2�hֻ0������YO��J;��Y��Zb��5	�����XH~��V����9}�m+7'Y�.[YӨ�(9��έ_;���n�re	D��:��]�^X{,�%kb�KzyL�^�S8+�Y}V��.͐B���� ����9�߲*w��FC�mdUt�z}W� �m���𢝀[(���ԙ��doa��p4������������O��oW�[~s�n�`̡<^�:/N�4ׇ|uѾ���SMb{��'Ac̰�5�/�
L���5�]x>���^d����v�n����E'-��
�;���u�X�%�K�p,/��V{�9���+D.�Ib����#���}*okUF���}w>5��Q���>�\!&�1���>�Â~>�%��.���O1�A��K2��u=K���@�㬀��O
�H>���rJ>�������a��$�I��0�b�5/e��(*#q���Z�y9��Y^0n�?Y N�0z�J�^�P���~��f��k6{EP��ܔ��ܝ�wC�m糙�غ��xz���N����9�;v%�N��* �"'u�+szPs{��W��y��N�3~Ċ��¬�U�)��@�@�W�}�ϻӧx`��A�z8@��?��dR�$�R
yYYOf���l���OՑg��73�;lA�c�&��U�b�8�츕���ۀ@ ��a�7I�˓��=y�y�L�"���o����m��xW �d0X��<VPb��CF��B���*6�r���0`��LnT{j�d��.��^�{k�þ��Q��EB��85�U
�C��5�	c�QX@e�{};�����YáV]iWc4�
�N��h�y"<�,��?`5�{�*��j��f1V�)[:��:=e��6}[{�ޥ�:�~��^Gl�HU�u(��Fm����
��Ǯ�b�؉�	������V��i
��yS��,6��ǫ��50��/{J'rp�ƹwKk����+IO{�Iwx��+*�I\us��?}EĤ�k�~�k?KB���7�At]�7.�R���=0���؅Mi�N�w��^���e_����!v�0��ͿCPW"�n�a�ҙ�9�t���wV�'�U)��Jp;Zk��܏mM�9���}&�+4�a���a���
U�_�����:5�VɃ5_�#Y���B�٧ח�#���%
�&�%Wt�����#N�����%���{�f�6H�F���}�@�+ w�ߕ��f��z˺g�Zn�'�Udב̩u�d��#x�V/����]
r�����:
��$�CMxxA\/�h֫,�V��W�y�ڗ@wp�#%�)�����}Jk����(13Q�8k���R�Zn���W���@��.�� �6�%;�S���z�vP���R<��#��w�i3"��[K��宂hEy��J�p�e���l^����8��ƫ��?_�����Hb:�R�����o�Ժ��p��+b�����ۥu뱃:[X�`�旣l��8 �:7A����Uy�U��NLF��"��R��Hq����<=���!�$E��i㠨x{��:�jn'��1�{�1�K��?:J���V��I�Y왗���(� �i�V�=�,�+��n)#H+�bU�����I�|C5đ�����fm���@���
�l
�������xA^O&��"���f[�-�c��G���7�8������H�\�WZt5�;��gES���q=�zO��G�h�9�h�!b�����+M�p��T�q
�^V�āw`��Ϲ�]d���3+>�e7*�<�*�ᷘy�=� ��	9k9C]�+*�V���q�ӫfemsUmn;�����Gٝ�s��H��0~����ꆔ e'd1��D�;�y���`�,q�Ӏ�шZ �^�+2)e_����������z�՛*�
��Z�L@ƺ00��W�{�5�5)=4�^�~�E^����>5�`���׆�׹��S0�A7�dl��Q8;���xk!�OV�^{{��;ۖ���0x6H��+��b�s+Å.����$�\<�e� C��=:؂��8Lκ��<i���������ʦn��������6+����J;�L:�\;ټv�3�L�^�\q��p��E��p�O@}!.b�f㢎��<5�5�Lh�~��埫�9{��2������"�ƌ <�����XU��c�/	m�y�����8[�[&�kl`5h��˶ggs<��9Y�ev/(Ì��j�F�Vp��B�>��N�e�䧟
��Y] ���_!�E{w��D�[�����Zy�Z�k���Vl�[��iJ��	�11S����Cy�v�ۻC��-��!;>��A�\��"���u  X)�Հ�6z�k��V曬;kSTA�o�����`�k��W��^�W$�+1�Z��ކR�㸥2�]�+٧r��� 6f����ACZ����K�B1���6�,N�9��ʵ�Ʌ9�gb���`UѬ)��BZF�L�1Y|(T)aXfP�s�-3�!͏x�
�nt��>�B�
����<d�%X��ƾ����"e�v����m_tƪ���+�g�C���!����             R��z�#��^f%XLMC��3�W���[�c�f�{"����hc��),SUr58�ΚM�ᖛ;{���l��NC+Z�u5�.�"�<�O3u�H��=z�[�'���]�o2������;�$�n�g���yݯ�-i��j表��*=;�=k�s@U���^oR�Fl�ɴn��	��wW(o���A�{����v,��wE�ܟ̈��
�-t���ص�x {ۢSmKΚc]!�xP|^�/�ʧ�=��[�׸ e	�mˣ-�CΙ�0vTh�R�Zu�2��J+ɋ�K��z��0�z���I5����ɗ�s[�0���1���OiVT�@ta5�:׹����۝Z��1|�ԩ|�����ܐ���\Y;{��{�y�   ��c~����+�2H����)�\�\�r�(�c�k�u�������d�n�8�!�*f���g��V�5�Ye�ŉ��ee�q9.���̌2��,8ǝaF����X9���ʩ*����iL9�F�2�<���j#	ɉ��i���G9�pd�q4k�r2��� U�Bo6���
���\���ݪnӘ�R�� R��\��y��O9tx�G�y�cp��߮:gf�e��`���X��Ӯ3ƟQ5�r��V}���XA٦�`�(W �2�g�G�C�⟑ݍ�%oe��?![�wWJ�NȺ�LY��]y]<���{���������Mh���e���
�jZ�E� ���W�>�ow���=�@,0!���Eo�5�Xh�+Y��������p����lV�q�xT@���qR����}>qP�V���f�}���?`�3�]CNA��盱F�9W^�؀��a�F郗�Kʸ/��@dOq�H�NECݘ�
@VL������ӵ_�5hc�`��6���ٯ3���ޗP\ }��}xl��9��pc��k�5uhyӾ�y&Pv
fQ�l����̢�]��)aI�=�L��3$�yv�7_K�]���|s.EQi�Cw�Ⱥ�y�u�O�}���������� ���z�n��n\c3M-:K��������ӫ�>��U�e�1[�		3X(ס�Ý7;-�GΘ|X�>����-�xN(T�.�h�}��q��ް����F�t�p�4�FkDc��Pl�u��}�{�N[↊�w<<zȾ5�lK4���};�k��� �>⚺cx�wUu���� ���Q4��hG_yuF��f��0�]�0�_O�^�\\4�C��&�0� uy�ۏ���PC�c�`�]�6����6v�x�ۂ���oT]�\Q3=����n��t�U�/� #�ƉA�,�ߙ��>X��ʇ�M���,;{?_�z�q�Ή��=��|Ep&��[�yw�sAI_E6��qG�&bܻ,RՐ,�v��fV��ts�����,��{؋f���x��$�?�_|bS���+������«��HW%2����\�^w�&;+p�2br���Ѭ��� A'd_�@���a��ۺ���/I"�^�0VBI��}�H\0R�&�j���`xR�R�]��.����ܹr��r`�5q�L\<�'!Q7�)�.vw�I�յ�:�W���VB���<~��f�lx�f�b�:�yg�B�ҿx�]�lS˺�����rj�&�&�\�Jc0�K�+�u�.�xm���� �&�b�Ͻ�l��{w	P��VK��y;3=茿N&��c�����.S�fJ �)r�i�⩻��~ᤡ�����d����#Dpt5w*�GU��v����Q�<Ş��Jߚ�<q'�Gy�C��/ln�������1x5%�����v�k3����R��;̙B�A�VN�P�&ry�k���=��:�_�#9�m��1ӥO�UN��}$�����~5���8�l+;�6��~�b��Mjʩ�(C�x�c��Է���y�����z���U�����G��4�F�+��MgVx�t)9�RI���t2���I�Z X�>b,��W#�v���ȑ]�\�a
p�4�2C
����+t��{���H��VF�i����ut��}�� ��7Hvg����U��"kl�>��vA�0�A$�k�|��W��Yޢ��W��)���
���H���'�����!�Y\xY(c�g�����i].�)�{�=��v��D���C�'|�x��ׅ�b�s+b&����b���+ޒ�f#enh�t��ʈQ��T\R��J�t��	��#�-���6Gl���v�Q¦�dL�b����\�:��t脖��#y���{��ߝ�*��0Hvu���Ä�5���Q7c#s��zm{
�C8��oz����X�}x,}M�]�����#M`�V+b�0;�~WI6�Ã���~��h��I=��:<(�+��
��`]b��5���?7��p{�6܏ء�5!�4����W��[y�2�z�&m��胪:s����\e<��@�X�pyD�&_�!���I=$�/���޸;�?kY��$�d�Ƙ��t�Mw�-����?M����ω��r���0� �����Ǟ�[��&��:G�<V]G��뮢�Lt��$��4�z�=��@���w��K�x��U���c��,m[��}�j��W��#��n�Q�N��1��On���3/9e������`�Q��z��ޑD�B��s"��7�#R�t�搜M�s��+��5*�7{/ȟ�-@�Z�~�+
�;Y"m?H�<�K�B�
�cQf郗>4�߮�޼��M��7��6W��]�ۘ����xn�˾��^E\�����ic��su����NأSƮ��WP� }�p6H�^�L���z7j<�7�y9��VK�q��Q^U��oG�y�1=���\�Q���>0.4�"�n�W��oeD�����*�
#�����f���P�/m��5�Nm�?y�X;Oz\��B��p��eY�Go�n�lS�R�l6`�W���_�ZG���lK4��} Gi��$�e�`��H���E��!I��.��.���IG��)�*�:_���������E�p���e��ndg�/TT����[Z5�:��Q���5n�ÿ	�i�[q��׉�o0�jțĴ�[��>��6���v�6c�>�X�Y޺U/z�q�ZM?���=����%Q0
Fk��T�<��
�?i�}�j�����T���F���:h�fj�F��c�YX33ק�z6A�5���b���x.��h��]]au���4�O��y��(e��l{A��2�+����]��4�ч`a����=%��������(�pM�Tn�DTz}S�q��k�nב�Ju��7𡆸@�p�kQ!Y5>�d?-]�� (߮�X����5�X;�z̠���{�5Nm{n�K8k�;�
��*�Ŏ�ai�<~I�� G��Ѽ4�ӣ�O���R�V�p��+b�����4��[�~:<��n.4��-VD�̕�C���9����p�n��_&w�W�;*��ā����lځH�qp��
��޾M�3�?����'=7M~�
�8�t^��ᤡ��5|i:�R�u���UnW]���\����q�e�
, ��v���r��RE�4��>��
B�r��kƵ�q?��(<���{��!�-�tl��t�UiC��ʭ�[�
^������j�1�āG�q�.��݄2�]z\���+#�䕽pdd�}`�9�M�B#��,Ϭ!\,�.��Y2�}��q���n`�ɨ��X�=�CW2Gs�.�pWB�1q]=W�2�W>����k{��G��x�4F�ŧuh��)��Rl�Ϟv]=��x����M��emU���<�i�j�d�G��T*��I}v�a�%�5z`��wV�Ţ�ЮO��z���%��"�0e��[Uiu��x6�6�n�!���\�na3{�f�!eF�nA�s	��]ݘ��s���f�����bC"�%�<Z��מ��ٓ1�&U�UG躼�>��d���ۛ���Qrq���*oU�$U�)V��ߎ| �z�#�x^����>��״�!��5��\x �ͩ��c͍�~in>�=}��N���E�X��1����DG4�kÃ��ߛ�mw���H1]��b��X �$;:�ʆ�a3�x������}^�6`L��qA�7]B��i�ۮ����u��社����@�xS#��CR_s5��`}����z}Ì���_�
 �]2�AW���Wi�z������˧��esޏ+��'�ݷXu����>��vs׾����9z�]1�[5�,pVi 6|*��\([^��زk٫7]��3ڸ%�`�]>b�-�NYY�xc�6�-�Zѳ�fb� V[�v�ɫK���F�����H�����y���Q;O��Q����L�8&V�����!X�F��!2F� &��ITK=�=S{����֍s�ӫ*7�
���n�X�s�O'�@i��MK�]0��/J�Ge��Vh�)������^��^�_��,I��.>�F�f�*�Ee�zuo+�6���n�tkҮ����i|����(ug��ך)N�rBG�`򢅣^��_)q�"�`�%�O�w�o���z��h(>>R��S�D�ڙq*o)�1���S`W�%����f����	B�.\��q�<��99�q�W[�Vu��5Ӄ�^��]
p���v=���X�;���5)&>�d��B��Bq�E7J�%L�
���)׿/���y�����w�X{��:ھ�z��I�8��㵋m��{�BU3�O�7�p8�<o�+#$�f����7�ڹ�Y#�Jf�7C����l�j��|��ѷpc �t����`�{�m�[�4�v�6m2�_8��o3r&�X�q ��n�9��=�W�o`�0eԦ���{���@�`����v�ay�D-��%N�_3�8�b��=�����A>�GV��;.8x���F��|�$���u�{�晽���)�.o�I��ݶs:���Yu5�.=�;2�����/N�!`��gM.Nl��eMɺ�>�4��4i#�SZ�W|�qܠ�	�����>}W���R��tѨRnJ�:�5\w���z������Pu�wt¡˥j7����\Y� 6!�u�/N�*�s:��w�%�\�=C+��h<5r[D|C�m4�j���em-�cu"7ب�Gd�GG B@        I$� Jk�|A3���췑l9٭^э�Lgp*WR���$���i�z�t"��r]A3�[���PG�VZQvP�]��<�Tr-��S�1F�mgDm��*Bi���r�ЁWt�=Ժ��v�B�2+vS��bQ��X�亹�s�αe�c�e3ݹ�����b*��JC�{%7���{��J�+)�i��{[�!=	;�������ް.�4܂�Μ�}]����LZ�⡂;�0V��.�G��v%�-��*X�S�ڼ�x\�2�I�2�Q w�Z�Vh0%WGWذ�2L"]�e���Fq���s�<���u<�B޳���3E�{�-����V��̎������I�i10���y#���-�])E��i5~���	��a��  ���{�����Ң���"h+1Ȫf��^���SVe9RQT�f���UDk0���Yag���q�U�� ��td�TN2Q��<ÑA�QTZ&*��Pd�TUd�W9�ADjƢ&���\((��ȉ)���1�����H��Ȧ9�-`e1EMSMTCUM��bDEfM�T��0g9�w́Q$�]u�^�Y�Y�p��V�٫g�i�]��A�5f�	{��ل:�nGh9����I�iZ���V2�tP�lt,(G��3ǽ�/x���!�ۗ\2�Zj\��Ti��@�*3LA^�}�}�r��95�֏'�����vLB���0�� ���ۯ��}&N�U<ϨX8rZ�GY��Y��$��=�Gy��@ƀ+"Z*#&߇���η0��ifGv�����]pd��%�����υpW�e�_Ə���c�Qg�5<�وԷtF��G��`�W��_q�;f�=��/7'!���W��0F����p�2�������l��Y{���G�ZX���LK?v!\4�˹��x�����46Y�r���CK��f�d�'u�
��ufX��4#�<
�V��ҽΫ���ZD��� �S&�ѱW��%��f5�[G������m�h�;��ҽDfXﻰ��ܢf��f�}A��{�+�`�l˯�X��d�f��C+�
�C Wo�]`����}�n�����_�~/3�EN�l�낽fP�٭XK&űy�bW�K�æ��"��Y��W���'՛&�~�m�lˍˇ8W��dM4���]�X�a5W�����弤�t�"�#^�|+��c��{���a0TQ^$ߣ;;}�w:C�|�6�a4i��MQ-�וr��z��9;�{ů[�K���y���҄��
B�z��Z�f�~��yk���;��1��I��Q#ˊ��C�J�YU���p��^��o'�յ��!h�:e�$�5��S
��7}��qF��჆�f}a��d�tMj�E}���9��؛�ħ��.vƁC����#�p��]��O3&�׏yau-=��vY�v�`�:©�pphʛS����L���M8�_�'�9'��{-Fx_�5]�`�`�Uփ�kFԵ<|Kk�wsQ�Y��V��:՗V-�5��<X�.��Җx�II��@w�F��]���]^0x������U�|gzG4�^�0Q����0�i�`�w�f���CZ��6}Zǭli�f÷-	�wF��cExc$�]01M���/:DX�����$U����`���B
�������8�4�դ
�u�4#O/ |�9�o�!;�V-��iɖ<�f�WBT˃�*$DsH�vvE9K���}�̬�<)f�x]W�e� ���u���&]�������u��.�[e����B�ڌ�٭�V!�׮��uD7cκ\�����욘>[�>Aj~��;�;�E�j����U�376�=�fK|aΖ`������D�\q�,�?D-��ow�>����^��-F
�,<+b�X�N��
�*�!���=B�m��}}���A&�eL�����զ�7��]~���ӭ��Uxӆ�w>b�ڳ]x������;���C�p!�����N0 �][ u�,L�k�{7�~s}?�?
�\Df��^��c�F����$���1B0�_���ցC�$k�iͼ�kE������ˮ(���0q����x�תYS35� T����"�e����5�;|1��ۻ�W�zx�s���E�¯�c�������������GC\xyU֋ޣFU����K�l���#��yzCC=��� ʯQ�F� R�&Z�5����B�)��k9x��e�	Y�ww��[��5l{J� If׻���u_u3���m��:�/�� xt��R�@.V�j�f�����?��Ή�z-�����t6\S ���B����k�> ��7��v+��^P�t��M�G�Z�P�[Ǉ�ӵrո�I�Ȫ0��ױ\Y׃�@�=~�ǯ�D�(�&¡�~mG�SڏS�w�
��5VD��Yu��!\��y$����z���Q[Qs|���+β(��tj��b#دn�����P4~h���ǡ�4��)�W�p�B�;����2�e2���Z��f/w�8Q����cp}ynvN���7ԍC�(}XR3�����V��w�f&��ݛ��/H�(xa5.��YWu¯��{{?Mz�m
x�ݺ}�l�p(�5����
=�DxT�C�U�o����h�|�`�wM]�F�;*�Ǹ��j�q����Ɏ| �\Wf;�w̭��% f��Z���S�b�vvM�Y�O9���Fz~���'<�׿m�9HӷtTh��E
{�L��AG'b���v���ɏ;cBM�߃yY���9�Wؼ�;�˵y�g�>�eCbebY�}����p�d�{�^�o����!!�5��dC1�@	�~Ç��<�y���c����*��QZn��жj^0R��{wA9�m�R����@aW�Z��y��ʇE�<)�ψ��%�yt%i�F��xt�Ǩ�����`d�o�j�P����^�Y��=�)���^��s�[�o}�$Ǯ��&�m�mMW�Fr~�s]�W������n�}-��B������5<��'5�����.�N���3p�.per�����훤�R7��8⻵"W�f!�z��JD��Y}�U��$y��f����ʽ���o��ǝ���kpqw^oy5�8L-�u�ON���7�ۚ�F�O=��BнN�EqU�C�J��4�}��`淬x���BS�&w��.���mv��Q�m�?n���<�n��X;�ڞ��o�����x�E�uIj϶!��΢���6�G]׊j���9�佐�'t�F繶"W�t%�y��9=7A4��|�(W�q���5��.���Y=�^%0i:��`VG����ۏBɬ]L��Ƕ�(�y'm����/�T����uI3͊����;�����t���DY\���u^1�uC���4��t��s�7wxAn�z��*��|�eΙ���ߺ7�u����dt,�U�r�����7��=�&�-��t�:ނ�5R+ȵ��U�cCs�Q1�'�f���wr��
�$����=���{��/����2��9�x�
�ƚ���P7�T�_<U���t���\��S��7�PL���χ;�պ5}÷�ql}���z�M͗ӧ1��枺=x(f���.T�4��f�׹/)Vl��j����O�<�{����xQ�E�-~h�k�Z|�E�Bk�R����}����W�t=�d�CN�ptݼ���c6֕�r�g�ХtjaA��m>pE�T0��h �׃Ϛ��^�;V�R���gn�^,�fF�>�%�O��v�ۋ���}q� �J��w�nW���?{zh��Ѳ}�^�9������S*�=�LM�q/���B���wU7��s]J�3�X���2
���;�#�ݛw���yg^���i��K:W>���p�r^9�뫶q�;"㎊��!9�N]��O��9I���ob���k�2���ZKy�Fc^���,�_]q�:�&vw'.���M����G'��դո��k�]�z���U��l�{���6?&�MeK�O�7���V+��m��ep�c�گ+�Y�T~�.n�x�e�:c{�q�hu�{ےn�G1�i�J�2lY��(𽴩�Q_\*É{�.��N�ܿVfy	��aocю��N�{o�բ�4������w]"Ľ�nz��{Εz�g�Mk�q��ԫn(�j{{��s�I��3o�r��H��m/��?P̉\�G�=���h8u�߮��n�7��;ǾC��ٚ�Βzf��pu�R��՛�t����W\]���}��y_���bs]*�8�V�����l��Ӌà�4+�QЕ�r��gڌxw06qF��uw�:�3]������o8�(Ngķ�����9�f����Ϋ���{Cux��f�W��z���;w/�
�:�^U����Z�9ռ��-9ɽ7
�b�H�F�_mJc;޳Ai���Ò^�Q�X��ee��]�S�e^oH�C�%���譲Zp��+���^�mu�����|:��4���3��w�D���������N1�"P�;\z"v�P���9��M�u��W\��X;��gK��}�]�#�d��5��Z������l$ Â�J���#X���R8��5�8>}��__L=�k��	YDu�B��*�yj�8�4��*{C ���͆�,up���	q�b|��{Y5��GOZ�:��J��B@�;!ޤS9ͨ"v�|m���Q(�Ģ	gq�tٽ֖��2_^P�l����:�e�̫/�wIc�Mʛ�R��a�,� U��vN��>���	��v�h�f���}̝�            &A*P�NX�k��qu��R���m��D�<&�,��1�^ˮ ÿ��Ņ��ñ�!칐�Ք0�N;�qq�Qo9���gR�{2�qS�*�����Kv�P%�E�<+V�����͍�����|�L��%���������,R�dݾ	��ޠA�cEIz��Q��q��d�E��L�z��j�.��Z'l5���Y��ΖD���ɇ�g]�-�R������}v��,���u�rJ��M��3����N�"���Y��K����<�uc�QK�8�a�U�E�aI��r�w.�����uo�͌6��uj1�GnO�1��4�Hc���xH�ٝN�0�V4'\qs,�P�w���d";.��	�E���I1۪R�2P�km`{.��   ���QS����T�TU@DQW��QWfcT�G1�U��T�UTPT�QD��XQTD�ETĕTQ4�AĜ�� άI�	���"*��*�(�!2j��q�j���)*����Ne�Vc-M%,AE5�a@[�0��.p�lJi�b�d�'�2"��*��" ���B��� �2ʘ�f(��j���ʚ��ri��j��a�IJD��@TTP����\kX�ӯz=��.r�Q�v�ŊN�u��V���ڔA[����G�7���?�������<\X�F�\Z��G��÷������n�noR�d#Nڳ�}�Oc�ݚ��Q�b�.�i����=����rHk�Tf���S��������߳����<���Y(�-���9�,iǛ����w���mq4g(��j��{�b�e�_%�I��W1�@��dcN/��(�T�F���T�=��<�_����Eɏ6�/����m�?j��7�Jp)������T�c��-�{tQ�_*�a|x������y"���-Ƌ�d�ڮ3�@��p�*�E�Y���B�k�����<����SI�ҵձ��ڶ�qSYe̮��1��QJ�ͮ���h�y���m�������/3��߉����R�B���/?o��:�[�3p����iLa�]�ZN��t�As�����b�xf�6&ev���6�ҽWJ.���������ȣ��z���6dtiSO9���}���4�
K:\]����G���+�U�Z36-������tyF����Tv0>����=��:���M�[�k_.�1)#�R÷���b�{��^���l�<�=���9y���~��ۨ�?۾ �`�r�Y�7s̺�F�r��U��زG1V�-d��q�88�rD^
��E�t9���&
'+��]Y����_�*��9���\�ތ�zR�����*Q]T��Y�ՠ�����\c��r�����EA�p��kb�+I��i��{�k��sP������C�ޓ�&5Y���n�:����i�\�%�y�r�0k��y"W�5ޙ��׆���lgg��s�z�zb�K}w��կ�	���Ķo"�~������p^��Ҧo+{�ò�j9L�kK�Q<��PW���m����$�Vڵ]^�n�O+EY����<ߠ��^?y���n�y��2��� �ZO�w����啳3��q��Zt�7U'�Q[A�&r����d��+�]����s\�6�9݊���ArHA�kh��{+j�B�J��ۄ�"v�����î��f\t(�'�orb��X��O\k�~��Ğ���m�4���Ri��>�w�^#+��ù5<}��=�P�4���c��g���ܾ�n��	�r�U����N�~���Q+��ا{���ᔷ�R{#�So.϶(�'Vy��F��ۣZtl׹�5�7��U���WV��DO}�H�+�i^��������f�V���?q[�����^x�Fc��G�}^��F���geY�D��/ԥ�B�&-rr@�+"�@됊��Q{��� Y��}9�E��.(Wu=ťb��(����7��Z4��B�wp�V��{�I�=���z	�0������KW󣑺���u�\���|5��iW�ex�ҩ�O����Y��7%j�Uw��3���wg���xR�Vzw��v*�}o/
�Vy�S�d~��}�]��^O}�aK�<��B�b�^�$�U�
�H����Ӕ���X�s��g�JIެ'��쭔U�y�����SR��Yo+x�ߜ�.}��Y����O�w^Ǫ�s{�ˏoK�ދ�woY��O5�)�Av��HJe��tX�,ʛy���a�e2]�Tk�����
���c	ת|#M�*�OՐ�m�:`����b�ug��G�o��	4�s���XW6����ԓ��Qw�/N��O���'�*�����sl������{ǹ���Vxנ�>��N�NCQ/Pi��٨���W0y��E�۽�?�5��wJ:�G�Y�	�����d`Ӄ�i(،sQ���W�Y�q��rkɾqzMsuv���G�ߙꃝ�g�F�շ=ܫj^��ek*y�rF��S�4A�/}�8}':w�\���4K�������Ύs�t(�\����qپ�,��2ֲb��O��
ފv_�{j5�O^��1��U�y�ʬ7u��k9�j��MښZ���V�N�d�Lɲ�޽��i��i�qߗG�p'1#���:A��QBg����l��c��^*"��x�����+@;$�2����9�����R�<]o+�K�8�<y�?Hϖ��_V��70l.�WёU�{�ӹ�v�\a渺7g��S�ý�U�Dy�T<e�[�u�; �Et4R@@ر?z%�d]6�%���I�|�\E����Sޥ���wH׻#^�꣚��׏|��ƽ%{դC}�N���On?c�+_�;s}�6i������߽�/"U��63�{��	�.�.<���V'	}��r%�*��ѯ'G��[�K��Y'wf�xI�4�豙��ܻeY�=Z�f�lzUa��X{K_m��sPw�O*��Ѓ5v�K�/\z#�#]#x�2n����ۧ6&��oO(����v�c��|�в?eC=��S����s��k�ի�p���dCǊ=�1�[Qзʢ�o���R~��ؽYRׇ�7)-���Ǟ�5*��w5uc��S]yk��x��0�n:����~J�9��BgQ�9f瞃�W�y��@0��٫�zpg�&���Tf��.| w��*3]�����g�;.0�ߞ�v��u��{�m��'���o��.z�{�m5�T��9e�_E3���.�ϼ.�����U��냱D�E�i�k��Fv�届p��;�vbɀm�,e�e)9ˮ,gkp�ت�ͭ��b9U99ڡ�1�cL��5b��R�x��������m�y�MԿzE��+���Q�7~�sh�J� ��ӗ���Og��_z��=�����p�z6��{�~~Ӆ��}�����}��/�ާ�q�n3#g�Y�F��w����l��|�ў��*2
eG��/z��g��j<���]&異��wNl)�iAS1�'lV*|����rI�<��(��:��L�@������=�F�$6}���H����v�s=��ٽu�ٛ\�<z��M8�u[ �=s�m+�D�x1��&kd�՚���x���p�*������s"B�ؔ�Ty�ue�1���5��QI��zѾꂮ�h��\��5��<�82sf+�b3V�ǀ���r��{3zf�?x��u�濖J?-��dS��?km�}s��-�h$�U���ɯ.Oѯv��c�;�v(k�B;�x��*}�u����^y�6��X�{u�;r���O��l�zd�27s�It-��:���J��.9�S���;�בY=�T�YIK��nϟ{�!c�oy%g�����ƽ@>�G����?j���\Z�5��>������Wߏ%E1R�*�����ݮwP�r�n]��K�<yQrM%z9ot[�<+�Aah&wM^�XްhmtU�6Q}���N.�_YܣX�"0�2����&��-��4��1T�_p9 �.��<��&�3��%`�!� ��j��A�L)�
=�����gA�#u�j�s��Ý��S'�*Ht*�EӒX�(�*���u����5�>í�}�:��C��d�[Ŝ��t'/QE}���e��ko)�}La�J�ܘ�����M;{ͥ;'�)����}�>y�(�k{�7��Ӧ2�[�����n���+�%���e�A��z�*�h���4:�8OA	�Z��Y�j�V��>=��y/zI[�1Ǳ�y�f\��zsK&'���Sr�fS.��T��=t�EB����S$|�6�7�4�B��o(��[>�ݼ��ë:��
��2���$�I$          䋚�U9-Nli�15B�XknT��(�+��fy	�I햩�ڵ�쫎�XC	�:�*���S"�ۭZӄ�q.�V���U��#�yQ�cS��z���ά?��"7V�ޤ(�Q��jֹ\jL�`.a�T0��B粜���PQ;� 3��Az�-a�u��^�eIm��wC�*��CY�8�P��Q���C+OtS��B��.@We��!sn#��3WT9L�]̜��e-���[7i�`��Ҷ��ݖ�U5�L�)��ջ����/lbu�we��z�����#S���t=1��;��5}�aI�����(ȳ�epđv�j=��� I��8�"*$�v`�i\��t�.�� �.\�}�[:�s�kɯC�����(-y&�߸    �B���D}333�aMD�x唍#IJ�\��\���)j���"��r�L��j�"bC�^gQHHdS@�%!ę dd)y���Y�f"�5TKՄ�-	͐u&A̙RSC@R�SJ��a�Z�B��%#@I�Ă�5�΃!"A�h*�9@Y�7�.�-B��/aR� P�U_|}B�8�@cg޵�Y�/�#+��8~��@���ӭYG��c�_����=�@��-���Q��]�*j��{uqMo{vbm�`�L���6�Pa�ב�(�b��В]����[/.�П���m��+5�;F9���t����{7~�ܨ��V��.Ɉ�7[��?y2:�*�t]�紐vW��f�F��x���Y{9�s�����חa�����,�lM���/WN�u|��o��hdÈ����_3��e�[��9:�F.t�2�aoq����x�ώ:=3Y�]����.q&�ϯ��lS�^q97>{��G[w��s�ߖa>�חm*�ǅ�{�gد���A�/�x29�/i�9Ĝ(�q,����*��ͩ=�;)X��ͮ�yH�Z�~��2R5��a��Hq��'v�ܦ�5��x��<���^��eĊ ��Tƫ��͞��ٷ;8�c8u��.��9�O�\���\Fk����Ɛ��;���e;�9��(��v��O��(���}3nj��E��ɝG�6�z��z��1u�#���IA�Q�ME�_�%?�<��]:�vc�QQ�8�Q��=��P��Z͇R^g�i��df&���gj O-E�6��_Jw_��]�Y��� ů圣>M\,��̙����&yT�T{{|4��ߊ��|@�]�J�/���С��>�L�{ٮ.�椺Il���e>�|��#:ofe�{�9[ �����_V�	�*��S56'i�'mFܙz׵��wY:�vN6�^{�|o����[��8�n"3Ol����R�^��=��?��ć/E�ޏ`�[���EP~~Ü�,���B~BM��Y�1.���=ە�i��׺y+��}[qF�<q~�U����gz��/3^�WV���{�'s�+�xa�9Gf��ȖS��#���q��Jh���6�)���~�ϼ���E$�i��^[�O�gs@�cV:{y�_\eg;��99����k�����}H[y��P�O@:��З��_�-�N�2��[���K�֊�]wO��2[˕�	Q�݊��;�V��z�	���",�3iXq�z��f��E�d�a�M^��;B�����x�w��]�*X[�E�̞� A{F��M��nTt8Ε۰�&��o�\a;��{8�zOHR�sd.��4�He�f���eꕈ����?��rk��*�ʭ[X����`���5�gxM�#��3�W��뤘��f���Kܣ�j��
;Hs���d��[�+��|^�������f�Z��|�ƿ�$�q��a�pu>дu�©W-����Sј�z��]q�6��q1�g�$�:h,z��'�)���Oz�8��W!�,���D�(a$�w��<"�fo\��q8��e.J��R4�7�=ɬ�#1���>��ռ�4@�����>�9;��+�ؠ�o�M�x�Ƥ�]�d��S��r[oE�.ry�kH�z������_��=�yS��;���&	c:﷎��I�c������'��^���N6�7���zk�T�����Mtg�Clǻ�4��[���ˮו���-���e�_L���t*�Ν�C¨-a�m��ת��0�F���SQ]�[{�����'��N׎�L[���x�ҷ��j�rj�\I��˸~;<S���c�mw$���k��]�����Ժ��Y8��	{0T\n_��p�WK��DF�D�ãzn��8�Tu�t/C��)�ww$�hi͙,��2��M��1u	li��*�뾇sONoś���M���6�/k��5�(߫����^T��� �E�����a�+��=q՗}�z&}O�Ķ�8�.0\���Ӎ�.ZX����1�V�zkk<VjMabV{+�mǩʛ�ʴ��V�D�5��TsRBq�q��l{��[H��Dƣ����=�������2��qZ�гT���W)9^ܞ�>�]�h�7*k[�Bm��+)?���!��H����z\'�4Ð������Pny%�N2/����n"�3Ҕ��us=�O�^�p�J�{Z�\�*�沝����Y5%��;�s�B��\|T�t�[�:i�]����V�Ay�6��j�bi������zz�߇z����r���EP���q=�{}�I��K��N�F©W��m�ڻv���M�6��U��j��M��,?_�黯k�m��:o�?D�W�u\����yԽ��2����J�w�͹�g���^=|���d���M9���s�Nkڅ���?sJ��$P歍��Pe��2���G�m�^���]��M��g���h:�Je���$�홳��OS�ٚ�P���"Vɫ�w=q��V��z��������342%Ч���(|��	(�Z�#������P֝�yz��0'���$�t����x�άjd���t�n^� �(bmQ �m�X���Pn���0N.�$�������io��ߞ�`���Kp��{��� ���Ҏ�u�m�skڍ�ѩ�?N}������=��=�m�y��դW�����g�!�s�tg$�8�}�c2'\���ۢQ�|ߊ<cY�;}�g�����B�Ε��X�8���fo�&������Msn@���������9��*̗9R-u-wO{�`Bǧv mM3y�R��=�����=jN�P�ɼ�ɨ�;'!LW����i$�N���������a훜�h]a��3dٹն�F���s2����D�W��}C�!�ru��ҝ1��|�T1�F�]���8�;p�rov�ǝ�7H۬��b9��J`�=Je������c2f�rò���t$�RJ֬f�7�2���ݎ]x�7xW1�Fuw�՞U>c�<Uz��y,g=�p�ۮ�["���4��?P�h�����_`�����Y�op�d�r��邎Y�6o�]�ꊴ�kIU7t����{<[��gYǤ�g����6S��O����U/c�w�{3$8yQ��@�m=ޥ�2��k��υ��W��7�Ʋ.���B���z�5o1_�����&c�k��R͆�R+q�eꃛ�2������ƝX��^{~������9����\��Q�T���z�d��O�J2��HG�4�2��h�#��*����5^�d���;�T�9f�I���=<�:˞�'}�%73�^ś��N�����]׶,����Y��aӧ3^dR���*�c��M��^�:��>P��jOH|�]"k|�r��m��7읊�*ir�豐��<�k�د�Ѭ�3�Y&F��vYO�s��{�7���*�*����\��7��g��o��r����D_E1����}��ޝ�>q8�=I6Ue(���?	�k٧��\u��}Nf&ߟ$z���+8��o���-��������e�%�3  "�9� ">�i �k0���H���SA��h5�~���?�?Q���=zG�o�4���*�V�"Aj$�T>W�D�9�.X��Ĺ��?Bg����<t��b�)�b�����:��HC�IU���i��KpӖ쵞�k��f�I�YJ^e&,N8(��J/�ƃ�;�<�0;�4��G��N���{�j®��Tbg�s=DC�#W��b�n�4��II3؀�|��0�!�C�ETZK�G�XtFŎ'�'�=(�����v?i�bvNd�go�CA�����Y�IJP׌����H�H����#9rY��]F�1EiG�f+�E�0�[�|��c��Ҏ�s��g�;�|�e-zW5'��
hn�i����3����;"8  D8O�ht������F!�0�C4q�~f��Cn���6= �e#%J��,����ǃs���{��-zT����Jbn=�&��N���?s[�����g��g�e����*X��c�-%MKÁ�#k'$~�����d����-�]5B�,fG��ގΌ����U�o�~#v��6��$�2�9z��7S��I!ñRQZ8���E'����bh.�>�a��vhE�-im���� �~�>�)��^�':���8.0��%��$��SC�#k�FM��A���
H!�:/���'��UfBEI��b��H��e@��v{��u���؏�	�z���ЇP�	��9����W�|�|@R����kH�#�I$��`W��'�RIF��py�'���O���{b>)�p��nM�#���&�J��Ԣ���'�Y�j�Q�Z%�#�F#Da��֒I$!��7���[�Ux��Y>��"� I��˸���}a�M��:z�&�l�Ļj==��Fy
3��➮�/��v��ڡ���t���FFn�5(�~u[<=���KQ���;��I$��gb8�(ÔgǌUͶ��F�=9�Sq�ۼ���G]E�lY�fVᡊ0�ǭ1H��TJ���J�yK�!q��h��^S�ɾi�9o��):�ɾ)2L�Q��d��YI�T1�����{��Fت��������[b&��9��ܑN$%�ހ