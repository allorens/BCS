BZh91AY&SYA�e���_�`q���#� ����b+_            �                                  zР P(�� t���   �TC � h`,P h �@P 
      (�      y�R��HB�*�����T�U(����UR�����(URR��QA")�EID�(U�����@�����J*�*^�����Q;���;���M��
NuJR�*�;u@�l�@��DG3Iw%aЮvr.f�   �(� &�l�5%
^Z��qѭPU���]�)R(�n� �w���P	�<��;ЕS���;� o0�@;�\��  ���JH���U)(
T���S�J�W���y�i�`�x�� r�r ��@� ����Ӟ���h�g@O�` g9ꨥ����0�u   }URL�����׼�J+�C�0����@q�{ -ԑ��9�ް����@ T  w� ��*A
�A@ D��D�| H|��`=z C� eܒJ� m�^�<��@� ;��`��$���y n΂  P �Yw�� �� ���_9J`l9 d�݀:��{ V�	 	{ ��<�� ��� ���Q�})J ��%(*�E*�ER���%� �>�h����g�Of�T��
��aǰ{נ{�����:���Cu��   7�%P ��XT� �$�`�1 rJ�݀=��xz����䡻 :�@ ϒ�( �ԒD�@�) !(*UUO���{ l ���� ZRUV c�
n��<�9t�� y�x��x ͏=�q�B�
>=%% `���� :�UJ� { y����{= FEN 6� v@w`�6 x          �� �J@     )�&�������� ��T���5 �    �%D���@     ��JH�U2`      �4ID��MM�4�b6��M4�>�������¤�k���7a�v��A�_�A�b�*+�Ȧ��QQ^PAT�UQ_��;?��f�Q_���#��������>�����>��z_��S��QX?�*�����<	�!>�������<�� �`@��d@� � 4¡���M0�j� 4ʉ�PM2�i�]0 i�L��i�L
`P� ��P5D�ax�t�!�J��@2�i�L�错 4�.��]0 i�SLeWTJ/�eW(�]Qc"�a �'a �i�8`TB�2�L��t�i�t�a�!�]0`4�i�L!�]0�a�	�f0�d4˦]2�8�`8a4�i�L:a�L�a�.�t˦]2釆�)���0e�&�t��8`�0�La��4ɦM0i�L�`�:d��t��0�Li��L�`�&��4��4ɦ3�i�L0�L:`��4��0i�0i�L�`�&�4ɦ0�L�Θ1�L�d��4æM2i�M2i�La�.�t˦0i��L�e��tæ2i�D�&�tɦ]0i�L�d�&�t�0i�L�0�Ld��4�1�M0���2i�L�a4ç�L�˦2�L�a���L�3��e�.�42�L�a��L:a�Ì:a��tɦ0铆�&2�L:`4˦]2i��4Ɍ:`��4˦M0�L:4æ2i�L�a��4æ�0铆2i�L�a�!�`�.�8e��t˦LL:a��t˦]2铆tˌ��8��L��t�i�L��t�i�a�.�0a4�p�a�M0�L:d��4æt�.�4æ2i�L�d�&�d��4æM2i�L�d�&�ptɦNtæM0�L�d�<3�d�&�4ɦ]2i�L�a�Q�tɦ2i�La�&��4˦2i�L�a�8�a�&�q�ɦtɦ2i�L�e�<3�\a��0�L�e�'�Ld�.�4æM2�L�1�\a��tæL�a�&�L�&�tɦM0�L�e�&���&�tæ2i�L�e�&��2i��M2�L:a�$�e�&�tɦ]2i�L:a�c�t���t˦M0�L:ntÌ:a��4æftɌi�L�0�L�t�i�gL:gL�d��4��tæ0�Ӂ2i�L�a��4��M0i�L�d�i�`��4��M0i�L:`��4�2i�t��M2i�L:`�&�t0i�La�&�4��2i�L��2i�L`�&�4��M3�M0i�N�	�L�`��4��M0i�L�gL6�1�L�`�&�4˦@�aS��t���A��dGTJdBdGT@.�Q�
:dL a��0i�\`GL��]0+�$GL��TH���]3Q:�tʁ�$WL��]2��Et��I�CL �At�.�A�(�eGL��QL"i�0�Dt��0�%WL�feL��Q ��t����2�Tt� �e ��i�2��uD aTBi�J����uD��]0��tʎ��Ȏ�Q� �eGL��]Q�`GL ��*�˦tȏ�0#�%L�0��%L�i�&t�.���Ttʎ��
:aGL(��4�.��]0��AtȎ��
�a���'�����ۺ'X�����{0!�V��*ar-�ޭ�&��<Nv�# 8�����4=S��gfp�����R{7OP5�%�K�4c|yty\ˉpNv��u���۶	�ܖ^�oe�N�Ն�]�[8&�9�c�踲ҕgo<qv^��>-G���w���B��u�c�l添�+j'�\�r><�����{�As�g$�:𤌢da�UIGm�;�gZ�!�A{�0��׵vs;�f����;�ŀ���V�e��C	��u��๸��_ �L��f&8I������i7�	Z��o�ظ�wH3[W��b8\��u�8�^ӓKf
����ķ�f��3I"#>5�'�2 ��0@L�8�[9��gdD�u�3��\ha�=�#�i�F�b���X�h�g;C�k��nn�T}��LS����+�b��!~�{`ĵD�3t���>ٚ�ٺ$�5d��[y�n+��|q��8kx��VN8��霧]壁�d�n�<=Ǉ9=�xS�*�՚�p���<�:h�<�{h� ˸�+c�Ѱ���n�1��td�lȮ���>6 ��b��5b�MqEq����xf�2��ӻݕ��R�Rrd�km�~��h�2���hmn}���L$�[y�8�˂(�3���9^x���[`��[�f���묜w;���kɈ\kZ��4�Lص��Xxs#{{���v��rò�Y����m��7����1�ͧ@MO���9��<
�,^�w^22(:.�$�N��*t'�f���@vt=�l��j�an�!|V��,ގ	Ǡ	��;�F���=ܹ��cgf�E�T0���]f��IMŗy)�e�dT���ŠV��j�K�#��.	R��������ۂ3���bk�d���N��*]�c�\S�A��n��&��ui�8+�*h�7��^u�qb͂`#�4P�웏��m���Yd5�r���L���S�ne���xQ,ڹF��3^l=��*/�^���<�,�z�;	�q�0YGE1n+��ʳ����u���2c�b�>--;�c�c3#Z'��W��e��.����:�GA�.�bs���L� ��E1���w��J��"/{����g,%�[�Q�/�qa���ݯ&��n�4j�r.U�n���βn#�]e�'x��=������!��幽��Ef�\���b���f�i����������欓z��D7^�م����W��N�q�pȶ��+�i����N[��pb���ۧ/G�I�<�`���ѱ�y�1�m�Z��&��A�h�f=z��{��Cy�� ߒ݁�p��ڗ��q�~�����L�\�]sC�FH�	d���Ҋ���3;U<���d`K�sz<cosx\ш�¦�ۮ��TZ0%�`BY�gǜ-QE��� Q�Tb�5e81pwzd �-䲭��׸7I�b�� fm������2b�N�x>YިnS�7�*��+�$�����wU|s��게t�-WDd��œ8S��{�9)i=z�I���ol�t��)�E�(���b��bMnM�R����Z,`��-��1]�N@��٬���M�|�e�ozn�rM˂�{cߤ�봇�w�c�l�7��z5[Ƿ�#�Q"�U*�8�����"��^��c7rL���u�|�in�&3{����7GI�:�'����T����Jkͧx�k���ݓ�+w{�7nt�,���.��e,^��v]Z�����F�0�9p�F�Vm*ëv��e{ܡ��Ku��z�\8p��ܦ��Ep����+�D�..5�K贼������b�{f��R���٭�Nʪ��Q�:��F�sXJ�˲����	�-��y��\{��ۘ�H9�g��F�Y�]�Woڥ��I�>��;�7��U�A���Y
]w4)��ZO�bm�x]P�*Г
w#���Wwq�:�G��y�v֕÷}�^0E.p`�9+�C�z�ˠ%�+��@r5toC���]��e�Sq��d��Z����b�Ӡ3)��N���!V�=�r��~K�׍�؛���<�[��˖�s��R�hyݫ�-�u1Z���w8�g��tb�0Zm�oX��f|�.%��c���]΄=}�v���m�.(��N��8�\(9�^k��f��C��v�^��Тǚ8_K��s�9A�c���}�îr�ѽ�Z@\�pr��6�����*�,Rns�7�l	p��´k،#���X������PW1{�ӄ25d�:�]/A���ٵʋ��{(cR��6�(͖�IV%��s�ji{\:�y+ٽVvj�4wP�}!�
�F9�U�5LB�����x��a�7m��Bq��\��g-����z^�Rl���8��)n�� lB��ͩf舝�37y��X ���)c���6��X��^Jo%��d��9$W�.]��`��Aہ3���4|�dhRf�1`b\���s�{�8�˴p���s�٪�u�҆kp�eܜ�	�F.��aA�f�Ȱ����o!��owm��8��b�%���d>]���庱k]ˤ�e��۹��(�/}5���(@	���Qg2�iv˝�^�|N�U��lR�3�[� f�@�F�:��/5ߕ�2yp\<Uxy��7F��oh��'��;�N���-�z�<��f�'Q�����օuu;���U6�oa��$��ʨ@I)Ol�}iڬ�W4���.&ɭ �0k@�xE���dZ�1~]�ɗ�95̚�=����8�)°�»J���#��Xi�׃�	�j��=�Fj˧XT�&t;�=�t����Q��N���_�7 <�d��������ǎ���i��1��(6-[��ӓ�/�&̑��n�ِNջ!��iBL5�F������{�8��j�6)3�t��z�ه��po[`5�a�u�OP�<8l�FbÜhc�����j_ZF���0��v���iâ^\^,����ǥ=ɇWi�8��o
ii�X\��	��8]7
�[�7���<�N��2�|�s�U�;%��kʊ�Q�H��v��pѩP�K��]�L��(��'@�W�n�qO�|� 6h(��,��z��e�H������g"�=sc�ja᫻FK�&�n-��v�v�֞Y1�uo>��7_	��3[��L��BoGp�'C���"����H�_vV����Òղ��T]pr�0-+���O����A�<�a�W�����f]�M=���M�c��ʣ�G7&�hulV�����M�{7;Ao����|�0�g\��>�)�_�}�lꭇ� �9�$�[���"�3;��X�b�[�h������l�n��ersz�\�tɚS�8a�&�@[�f��7K �ۯG�.�˫:n��n��^/!ut��=�&/ehs�k��{9�^��i˯nڴof�=�;4w��ZH���}6��#�d�������zq�ms����Å�]�^B��m�Æ �fw96�!�S�F��֋T���<���Ĳ<�B�M��sB��Pзa�n��������г`'����,k��9ѵ�x����հws|��f��?��{��8�i+Ź^ەל7������v�����]����U�Z�,�$����5Ƙn�
ixb���$�j��&�W 1{�o���g��I�"q��D�٢M��].-kvZ�V�"�����;�Bu%e��
��\#L*���JsMᶼ3�1MuѮF�#a�^DT�M:�e���v�M3SwP�򺱅�s��S��ԓWcj��x��:�+Zk�����6^ d�v���٩h�f�-q���PM41���[��E��6	װ�Sڄ[�ޘ!�u|�{�~�"����#[n���Թ�ɺ�t��BEt�={�>���;�kdq�ŷ�N{��fwrz���tk�+N��U�ͅ�3yH��_n�E��H���9�<�dS.�k��;*C]���;rW�v�5<t�`�����j�8s��.�O*%�z���qDD����&��1�%tZ�s{��2椢�F�ڻ$��}[��	�W �D� �����k��}��s���O�q���v�i���*G���;q=Xm���:�gQ	%fwu6�@��q��B�99�Ѫ��"���Vb�i�Ʒ�У�F	;�ce���ެ�8�ٮ˓$6�ZC�sgc3�����:1�,��[��̋v�� XQ̜�ӧ�w@�**i���*����J�i\���,nHb�}2��\�$|xmO���7��G���Q%��ӳ��5ӝ����t�FX_<Z,L֞\�G�q�{�9H�&��&���gf�R�;����&�z�j�ΔGZG)������x�i`��88��Ö��3m��t�Z�e�8���dy��N�i�k��L� �ڱ���*��ӷ��4�y�s��lwR�X�k��#&�"�Μ��DZ���e.׷J�MZ�h,���QiA�Z�*����v�����ޯ�݅`�;&`���7~'qr�A4z,�p�zݦ���f�����Z4�(+���X���C����r=u޺.��6\;җk�8��~u�H��r;�'ge�?�_�wXc��+p9�On�:�a�;\�2\��A�7k�w^ݏ���� �����]�7s�t[���3�$��܎ޛ�>���FT�7��8[/״�:�G@;���}�"��2t�@V�-Ӧ�&�̖����V�vIҹ`ǋ���c���*vH
�R�;��0�y�{.�n�0i�+�
��O.�$h:�ۑQ_v%��۫{�"lV�].�v�s��n�0n*���61�ǐ�ߞkiU>��uX��q�#��ȵ+~\��l�i�x.�"��������m�0^B�6���������G9���Xз�+!��
Z�9nWj����P��3{e���F�/L|�+V�����z�|��(�]���q��J!��i������:Jޡ�a�U�؊��z:��hcA|�=�㔓�i���K�i��^��K�Lm&7N[h�m��[���Zww��qW{d;�1L��r�"Zco�{�F��w9�R�Հ�Y:M�9��j�daS�rH�<�l�M}8�K;����GIR��wr>H�rU��wx��ez{@7a`Ӄ�P>>%z�	���;��N��/�Xr^�N���F,}0�O8���/�n�[X�>O�Kg2v����x���G7��;���7��]�g>N����\�鴱�Yr6r��,�3n��<os���@�����8��l[-k;�$ V"x��&�:��p�I9�C�،%ZZ ѳ��ʘ�ͮ'�+���'t�Ť؈Z�W���A0��拴<�>6�#r��� #�Б�G!��Iy;�8 ]����۝�S�{޾���s�4��Ꮘ÷��,�عr��}���QK^d�vK��]���qE7�ɝ�+�ww��s�NɏV��fQ���.>��P>����O���氿��}^sE�8���CY	"`���7o`dŦ���#�xa�"˩ хԛ��,�b��u�gH3�:wl<��{N�,h;��5I��R��8�B�s�*5�"��\��W2���]���\��v��Yw�����VU��74Boe�ď
��6hX�moBgvwb���K�eO��!�7o����=�a&����EK��(�|U�Z$�I��a���Գ����I-��0!�O�}ߓH��i\Y+�|�����p���{NLx�K�oD�j�Id�i��{ՙu����IG�o�O�	��_t�u7��4�N��$%����RA�ID�OS�t`d�8)�G�L����$~<�ڶ���	������=��$S�[0�ID��� �ID�Q$�oJ�B������B>��.+ j\��q��0����pH7��N��C�A� �����=< ���>Ԍ���-��xx��#+�����l�����X�:��v�Ѥ�(&�	d�i:L&�鬿e��Y#�n��g9/Ӻy�z��i���������1��(�M'I�a�)	�t�Me��O�D�|L$�I�f{�̟݉;F�%���t�IL	d�)D���J%ID�[��2a!��t�/Y�w�l�'��|J>M�H�(��M$�0�J'����6�S&I��Q0�N���t�\�=��C�2�/���x��}ϡ&s������'��`���b���Z!�L:��pY6��i����>�p�z`D��}�'G�=�t�6mD�x�����]�2�N��g�CO3��C*����n��y�Ƴt�;��Ȓx�J1��{��;�&�i$�L:�I�o���̤m���$�t�K$���.>�w �	d��L=.>9�!O���������c��=�x���:M&��0�I�I%r��jj��Sp�l��;8\����0�� ��I(�Q(`�	8�0q0�%	$�Y:i+ ��r(J' ����I$����/��Zz=ؙ,�I$��ct���O	D���S�"	>>�����2i�a�����t�����vq���k��N	
!-'I(�\��'I%�&�<��N	�i6�d�����i$��O��|hUnx!�x�Ǳ|e.e�q��ZF��k���ԖN�����jީx�{��Y��0�R�&ĕ�ɑ�邱��)A$�I$���:J$��i(�]7{���� �Y3)��,8����{��W���������4o����W�)>�Qr�@���Q(A
(B��G%)U(T�iA
@�DL��hEZDL��UrA2C%��D� �� ��R�hPh )J�Z�C T�A�ir ��J()ih�P(i)iT)*�\�L�R�)h�
T2�B��V�
PJT�D� �ZE�@
P!2)E
 W$\�h@B�L�C!P�\��rQ�R�JP�R�@�P�
@D}��'�q��@����<�O��oXp���3��;����rɺ��S�{ծl�9��8vO�Xsq֮̗>� ��&nĤ<�%�6�38�6�^o�;@��r\G�d{��^���=$���4�����N����}\B�#�ǯq:�8^I�H<����S�x��:������p�EG1Ԟ��.xˇ�u#fwܧ�:�au��S�2�9�#r��Ό<�}��Y. �Oe2y/:������;Ǩ���;8μ�N<����BR�d�V+��N�1�m�_A�=�:H����ww��ױ:y�U�����O1l��%��7
�b �Ci �^��g<!��<�R;��~bMww!�x.��8=f!�ڪ �?�w�ADP���_g���'�������q��/���>�,/�5���{��{��6`xqzW#��Kww�Ў�}׳Ft���f���ｫR)۫�B��Ԇ<A&2/����nV��A�P�V��~�a�.�����
YX��e��|&q��������{�{�/"��7l�yf��}�@�#}K������������EC�/x�ba�D�ڎn�,��˺9��7�a8j�.3��������aB�P;�|�d䒫�Ŕ�{�7׈�/[����Rg�T��{Ӈ�=��
*ol��ht*'kM�ۤ�O/����>
�Ђ�n?o��x���Ѡ���^��]/���Kc�}�r];�@'|-��wfy��n{]�Yҡ�Zާ��#�sz���|���(q�z>b�1�K:�z��Ǭ�zywx�i޶���k3���Cب~{�i�<=�O5��#W���/|>9���w��vxB{ˆF�nǋ}1ޛJ�~>D��B!�xg�d���bg�{�{'��d��+�vz�xqR���{�����]�̦�����F� ��b�$}�o�=�n��X�߻��o�����w'��8�5�t	�^n�.�1�*x�����Ne��ǷMN�owa^�\g���m�����3�o��>��۷oNݳ��nݻv��ێݻv�۷n���nݻv��۷oݻv��˷nݺv�ێݻv�۷�n�۷nݻ{v��÷nݻv��۷n��zv��˧nݻyv�۷�nݻv��۶v�۷nݻ|v;v�۷nݻv��;v�۷����^]�v��۱۷nݻv�۷c�nݻv���Ƶ�&��G}gm�nitN((��{[�>�����ׇI�#�-�}}�:o�S�K��ƛ�q�ćA�o��4���gs��y�����ʚ�ѡO�x���4!D����SO��d��>���	sJ��g���wu�.@�pv���ۦ�9a���}:���{�Zْ�4m�6�w� TU���e��^�]�����n��sr$��۳��=��N(���ǲo��7G���	�W����:���?wN�=��۱s�x��b�l��Âo'1�"�ffy�\T���$`�}z�U������%<�}����8��9$�o*�̕i���x/L�Ox�3ǫ�ӵ+�'n�d�{G��aJ�0sSئ����5No�<�sg�bw��9�F��W7H���v������ ��cN=����_-��k���>��-�s{"�����6��A�������dI�v�E%뗷L�{&��Kz9�����3O���Z�f���f��9�u�c7H �h�,�,f#:����5��n���R��̒��l6�}:9�{�N�3��oa��51�J�=����B����to5����x���.�t~���Y�T���P�����ϻ����v��۷�nݸ�۷nݻ{v;v�ێݻv�۱�۷nݻv�۱۷nݻv��۷�nݻv��۷n�;v��nݻv�۷�v�۷nݻv�흻v�۷oNݻxv�۷n�]�v�ӷnݏݻv��ӷnݼ;v�۷oNݻv�ӷoOOOO/.��v��˷nݼ;v�۷oNݳ�nݻz�}�OV����wם�.���C�g��
���*;dnx��^F{Kl��k�9ӧ����.#�2nx��?w��f�������9ff �ٚ�VU�0�<�W��ɹ���Ȫ��MT�/�%��(p�L��q��wV��X@���2�ۇ�읆z�C��"d�һ�My�u��Y��A[��j�gy�u�N�Ưnzy?s�\��e�v��{�����i~�]�Ϲ{���ӎ(���p�p�y�8fԽ���3j6Dn�<:�C.DK���k9��w8�O=������qg��q�&���g�~0�y�����H/%��[����f�ch_"����+ч��f�XF���!�y�Y����^!Ð��YW�&1�������>0^��$1�8X���C`��C���wo�eF׾~��b�\����:�g��:AK��ˮ��0�����s� �����;�}��{��t�S�� ����u�M�����b��2��ro�^�=.��ս���������oM8�C�;�??<���|Lo��3��p	許��Z�o33�`�.zr���f����N���BL�vaM���;�վ�g�vP}�ٍ��8���VQOK= Xї�d���3H����u�����^>��۷nݻv흻v��۷nݻzv�ێݻv�۷�nݻxv�۷nޝ�gnݻv��۷n�۷nݻv��۷�v��۷nݻzv흻v�۷n��ݻv�۷n���nݻv��۷n;v�۷o.ݻv�۷nݻv��۷�nݻv�����������ӷn��v�ۧ=��g����{=��?��FK(�[\�H����_�]�\�_y���N�����]Ӂ��$/sZSz�=�j��O-���\������|��3uKs�l��ˁuV�F^R�H%�\�r�d�
§#'��G�L�@sC��V"=��ǽ���	�߈k��	1�4"�),[=1���V���S�_I�k�z���D��w'����nyUq�ϰ{�DK���+�=������0��;�Y+{����/��t[Q�r!�X�^�A�=�q�07=��h-�o����;�/�׷Z�b9�{)��{ÛZ���ϧw���{�o���ݝt�;c���ѐt�N��٢����_d�	�=Vw_k� �|:�3����O�5�^aj��w9�,lj�ǆx��}H�٫Ӳ���"�'@<�ý<{�|M/�?mAw{�v���2�f���8�՞׾�N}�وbWa��O�{op�s�)�T�n�{o�>G(����N�n�ZAt�3��5��7����_�O��4L�vaab�G
|#u��%�4U�N�/�v?I��=ٻ3�Ji�?���Y5q�D���5.,�ɞqo����6�٣P���Ϸ�ٽAF�8�B_ヶ�\��xR���Lﻤ-����C�/��[��=7�l������~��||v�۷on�nݻv��۷n�;v�۷o.ݻv�۷nݺv�۷o.ݻv��۷nݽ;�v�۷nݻv;v��۷oN�]�t�۷oݻv��ӷn�v�۷nݽ��v�۷nݻv;v�۷nݽ�v�nݻv�۷�l�۷nݻzz������v�۱۷nݻv��۷�v�۷au��ᓛ�G��>�z�f���Ū������X�b�~�� ܠ�d\�MB4N+��ħ��s��n��V����]� j��������/W�4,Ufa�[�z�)��^��J�=�۸u@-{&��E�q��E�?.�9�7��>��F!��~���3����~ޛ�������6�\}����V�/��b{�k'� ��������۝o9U�7����Ŕ&^1f��غ��e�{�u��o��>���l^2&u�s��x�>O��3V��x�^���'N����?m�S8{���r(Eoo�i.�O3�+3w����t��9��"�J�j:~�=�f����c�����]���������{O���x}w�z�U�'�F���H��x���'�{�g�<1�3R񛵲��[�MW#��.8���nx�՛���a�{�D ��Ƭc誂*H�0�"���d&1�<�<�=��?p�d���Ip��b�rRLϰu�`�e�s�t�����u��.޻���='P3W�^%Np����dh�v��0�l#o̬x��J���$|~�]7�p���/{{��q����^�=�e�_l�Y������vo�ކg{s���= k�S�<Tz��M�w�����Sb��±�w�:�'O�n�yNx�����Hi׀�<}����k���4xor�ڽTpܘ;ǜ�_�%	:&<��>�O��T�}�a��Ww��3���(Ʊ��e�ɥY�N�sڛz�6������%�P�x��y��g��ޛ��y�0��rZ&��c�ɼT"r[��R++�Ioy^*m��y����4?^eɥkY���{}��>�>{b��J{�'��&o����2m*��{g�`�(���JCV�)��ix�x��i[��}�{�\�碿��K���7��ۉ+��!s�'k���+��{(�痙C|�dEA���ކyd5�r�S*]ꪜTJ&}(5���p�Ά�m낁	�>}��c�08E�	�.�X�����K6��ðj�����z83zm~|��P��٫_9$�_'�$0t��a��佼��{�D�>|�;�t}�9�z�s<��<ф���{=0��]rn�Fg�X�g���p��z�žNH(·W�U�ɰ�<S����޳J�ЮY���L���e��G��[�&�|���ɫ�oE���ˆovD���&��X��v����gy*/�äv�= {+����}2M��獰��_�����N�^)P�q-OG�x�r;h�qS������}�I%�'���rb����u^���C}���_1��� 7&?<�N��|(��t^�n�i�ļ���Y�k�̇�WS",&į(�flyY�ڵ|;3P]��B�Db��Ɨ�%�a��� ���=�yE��ٕ���7Qk>�i�����HQc���<82���ٻ#7N�-���3k�q�ao�z�^
h���5��+�_v�e]�7���f%��Sn?k�q�b��2�x���8��GiA$f{V�pѯr�,t[�t��/����׺a�ݫ�s��I�eÝ��3��b�^���gowmS=x�LeYg!�j�_,�伳`��\y��Qf����\�M/�)[3tiBb���ryH6�R+�w������S�O�D��kl��E\Z�Ӳ�:�Q����(׭(�SPa�|G����O���Y����.ưf}�
���H��*���<���5�7�3����]�r� �djpÿzwkے�o�6^�+�H�B�2Ɠ�����A�{�T(�9P۾�7H�ņθݬF���6ǈQ�Hsf�Q�u9����kۃ.f�}ގ�xXX��� 9\�:`���PI���r���~��O�w��J��'������}s}�­]���qb�}q�&0�Vfpo�n,	��
��f-y�������q��٘�O>c����ۜN��wc�<�|�%��J���&c�q{&�y%���N�O7��Wb�hr��|Gy�6�����>��а��v��Ae��ޏ&�5O}4=�c�'���G�x�^�?[����l�ɍf��i�_j��1�� ����zT���(Ӟ)Խۛއ.�N�\�C����On��-f��/*A����M1`Y��|�#��m��������xI�#�to�1�����s�ٴ�a�j�z��{��r׾ˉ۫t�t@�.���jZ�5v�H�iڗx���?P�R�y��C�l�����9L�}<U(	�\R6�k��/�$�����DCax��:OmᏮ���W�]��������]������z�M۽���ufa��ͼo����&��zo�ͤ��<��5�����p ����[�7�ι�5��8x��pM+��PB�x�ww7&�Qf�O���}���ɜ|8"�� ����}`Qv^�}�e\*!^��{-˔��u`�:��,�d10�m���{�����jd���T��8�>a�qA	�ռ	���3���_���:m�� �ޡ��x����\��{c\�๻τ�HJʻ��mv���.J����.��Yx�2%'|e9'$]�b�x&����8�k� ����O���{�rc��E	��_ {I޷{6;;����Z�lY�y��|B���{4�=q�����pcJ��o�[rł�2��p8�D}N�dȽ9�3���`���'>���݋�z]�f� i�Y�$�PT\�am�w�m����_��=�N7=pWEm��w���(5͍{ײ�/�n�)y�۫bY<���K���a�tϣ)P��2m[�]��W*���B�ԅ�}���۹��j??I��y���@|珨��<��o)�2z�� ��{V���6��6��K~�8'�f罚d�s�����c~���Q�������7��!�q��Ք���}�s@Ї������]�4u#�M�v�ӊ�C�|o��!<���U�w������E�L�����iaP�_���ٴAa9LB�PGݟf���܌g�q��o�V�m:�]k�s���������}��݈ކk}�G�ល�1��L��kGY�E�{
睇۾c=�Þ[�h�^K����ǚJ�{��#B�罬��?u<���{a�=�������˷;a�ϑ�o��עy�O������{�Qz���	������:����<=U�W=og�^�C~�<w�Ѹ���̊L��>Y�VC�>{��nR�����)&���p��V�Oxn�=d������)6�:�o���ݽ�^�s��rf��>s��;4#���b�n��.`b����W�)B��E�snq�a^s;'����c�9�e�����=z
�v�B߽YG�<���������'���0�VaB�p\�R^-�mݐ�0K�͸���-p�5asׅ��_o�3J�a<<縝�
Ǎ�����^��N�}��Ƀ���#L�����B �౾�������{h�'^vb���l0�}^.
��}�Y��W�6�=>�e�Z�n*��K�{-�^�ǧya~_N	��N$F4�os3X�9�*�I	vg�\��A�&��x����[�`�ww�y�C�r˓��z.!�Й6�w���)Ǡw�<�5�4=��K��ٵ��{h��e�ؙ �ܛ�_
_�e`�751���Եvǵx�Pz��y�nVGOU�KZzI��t?s�'n����L*IϪ�s��l:=t5���	fF3�%Nvpf�p{�{�Nw��2"ԋS���V��y��w�����z�3ێh�w�}���7�=�z�M�/'�^Ny�Ҳ������+%�"�ٟcV}J�|����7����1D|09;�_��xm��q��������������'r�ƀ:Ӿ�Me�H3�<8���O��V�vlRo����r�5��>o��g��� �����������?����U{��?�������H��I��e%�]��zY��	���)X��m옗s-���NSKp&��&�.�aۨ�T�u�ifs��u���E4jݯ�y�|9_�]�E�Fh$�ު\2mu���n�3��pƚ���yr�&3��ɖ .nd�-�)0�x����:�ȣV.�9�j1Xƛ*˵+1t.�^0�70l�'j��a�mk�Y���W�<ܮ��i6��@���t�|��9��<ܗD�i2��`�cse��¼�5V:a����A�M�.�mL�X4A�1�.\����1x�\��3)+�4��i�0l�Y@.Ж��IT�ZU�%kS��4Yr��+k.)f���f��k�i-c`\1�-v� m�8X\�e�A�T!@q�XQ���WQ-WL��Z\�� -���hB3�ZF�6�/�b�.	���j԰���2�� �E����,IV]��M��C]�u���up�V�^�A�q�l�қb���1J1nvn�!!K����#i6I�m�G2�14l`F�s�cmj�i\kbJq�Z�Gv��	H0���5B��Pe֯�J�1� Zf�	��0��;���2ј��䉲 �'M�wE���m0� �[��[�a�`���B���v�)@Ma\Z��ֻ�,�+K�ڑZQԬ;�%v��Bk�m�����-ڲ�K-�c��Cnte4�h©5s*U�M�J�ݪ�7�0�ZK޸fc�b��&�0�l^���$ˀ��l�KX�)1[͋��0��h!��u&-�Y�7�Q�1��v�6�x1�q)�24�ɒe&�:h:�B���Bf9�tMV���Q�#+S�͊6B$�k�F��lm����؛��k-6 eM.͖n�y`b�(JKq��Y��ȍ&3����-���
؛g9�6�[�Z*�.l*�V��l�;!֚��Cmp�"�LY�Ke �)�j mxaQ��]v�6�YaĥS��P�$��\f�0�K6�s�k3���Զ�h�JG\�nKXm, �4��q5L	.��g�E-�c2�j��XA�9$m
杞�B�XV���m�ivV�	�+�8\�ńeЫ�L�0�,��V�u�Z����(u:�v�Tz�HB��ut3F9��mi��4�U��0ڕ�%��	Jl��Ò�������]�p@�Z/P�t���H�*Tf��Kh�LZZ�]���(����pBm��0��v�V��J�4�e�0�n�uV.وC�	�%X�K�*�WUn@0i��5hq6�JC�.��ٳ6Z������)n��X($W�C�Q��1�4n!)
WKB)�2B�@6����i�19#���P��b9�8yԖ��m	����Y�ll�:��	�PcZD�&�k\�)��!M���]�vЕ.���9�;9jFz�5ݪ;4��p�5K�f��f\4��.��8���v�W/n[-�%.�)ɣ����P-� �8�b��M&m�Ym����j]#�mB��;J)6c��2��)p��{g�@ڵ氚mp�9��m�f�V,�n�r:\�)F!KpZ��VQ�v˭F�Z&��k���[Ի)b�n��TڻWf5P.MQ��)`�h�`�ڦ��[k���Jcٴ�,Ѭˁ#^�:��N�2� d��崌pkb�L�8�u�)*k4�(M@�3δX��qt�m����&�j�%��%j�FmeCm@5�q,czlۄ�ݪZF3\U�5jM����S1WQ��%ٴ�.2l;j��:��&�"f<�%o,.�2Ūg0�:�1AZ�1���-f�jڮêJV��M.�֗BUm�V�m��ͳm�X��v���ڬ2]It���[,֙,q��fr�L�XX�+�vJ7%�j���sn���aE�r�	�k��M.֙��Z�4е�C1�lL�F��&t�bd�{ka1��	]-rE���v�XK4���+��6�"��ي���,�I�i�Q u�W�&.uQ�4/:hgb2�ImFYKVe{[&4˦��&�˖[��b��
`�[5T�����.�4��8K�u�+2��Mm�,�Hk%͔*ם("�e��`��8U�,F�x��bh�щ��3��J�kqj��{�8b�;�b�	^6&V��ɭ�Q1�Ŷ��+�Z��2�Ќ(�\,�Z�R�T%�My���IV�YI�1F1�h`�u�v����V�M�4��.@6�2�Ypuΰ�ζ�Цi�l�QH�:\�t�t��[�L`��S`��qJ�P-��&6�\$�h��\�̷�p
����Z�n%�pa-���S�UcR lF�%G�ݻCV��T���\�˖lB�@�F]�@��JVd�"���2�l���3��� �2˩�-�Z6��<�Ι����*E�-�b��av�W���ld)���ar���K�7�����Wf�ALI�u��ֺ4��"e.5WTvt���MEk�H���Ib��.�R�l��MoeK``�,�d��+`ػ��D�\�(j�)E�� K*�m@��փ�l��6�-lr�w0#�M	���r�b�Զa%��Fd:����#Ub��]��:R��8%�79#�K��"k��+QnVŷk�q���$��j�.�h�B�`Y��J�[ζm)mM-�����W=L���Gce1��lK�]�2�ѱ�evk4`�/a�a�fW=���l��!m#�]�s(�Srh���)������6�9���5�)Cq�v��L,ۊc4��u���b-H�5v��dt�������:�ɪ]�7��+��,m�Fb�e���[�W5G�@FD�u��M&�xm5e(^�&�%q2�sZ��Ч�2e��[1�QJT���(�: nHr9P:�p&�k�+�%54o&]G�ePcl��cl�a�`r�P�I��6�+o:�l���ƪk�����1�ʰ�����(��b��3h���VL���Q�4kk,BnXS36��.���Va��Л0���WvTtٚM�[\�{#[qn��1:^�Z�X�j]Am�&B̖���݃h��*
-�@v[��Zf3b��CC%3.��yKA�T÷Y�m��� 5ZbY]biT���n��ڵʔɡ�/c�+\5��tQ���A��W�F�xt��kl��d]t�{m�#v���f�NY�F\lMkPHJ�\ح���W8q��b�؁�34�M�k,#]����f�lˎ(h�]VZ�L�f��u��0��L���s�mf.`�G-r��������]��	�����M�&-4{BS6�ZKtY�[�Be֔�6�SK�����
jJ4��[�H�<KS:ڊ�ݝ���&uF��T�uάLɵ�qΖ�b�ڰ�i5�r+���M�.D� ��:m�-�m��3�����eKq�	��Xͦ�@��+��1.�e�H�fvl Z`F�ӳm��&�P��cq��5��a�Ҁ<d�YQ�HS]J��sSJ2��[(��	v`�ۆ������V�1��\������t5b�f�5mZڦ�6:�"ՠ�V
v�+t�JV����p�*)��[KiF��)��k��l�RГnl-�f�=�Qqa��,3�e�fv�G[3h]5]2�b�c��:^j3M�5�5�)]&�����-�dmS�\4�R��3ɵ�DH-*@��vh�y&�,�cKP�Kq]�bb��J
қY�1���ݞ\a��j��P�0�r��q`��Ƅ	����ļ\�Y�0�n�5�U�̷�R͝K�)�S[��#�EyŬc\�q�h��[,�Ð��憱��u�A�Q�`�C36F0-�d1t���]Z��X�c��t�c]�����DM��t+[L�خf1��\��0c6�UuXא�ԇYo\�-��)���BS���� mH����;Q�bf�X���]kcλR& �1:f��BX4�-��Z�U�iK�1&lX��C6ma1���J�&�	F�밶��G�R7�@�k-�F�t�)����a.�����	�ФsKr���t��8\�h�H"64���g9ن0TI�m(b�7Vk3�{H�l֢�eA�k����q4N�=bZ����h;h8"U)�nб�PT�M*26v��F⃵�X�X�6��1�0p��Fc�#���\�l-e[�`�Fѳ)��`�^6f�&��gV�t����Qe���<�e{ZŹ�K���aepqf��v��Q-�ccV:`[l�jF����1�P���*�:��h���+]GcZ���(�thƙ&�UM������t�]�vL���f��nfu�����c���sb�V**���!P!��ԩ���{PX�E��F�.��t�vh�۪إ����.�V9�Yt��3�������6�5�ܦ�X5A4�J�tA!�sm�rKJ���U*E��k�R�Z�[���B4��|7��T���W@�KtZ �[1q3�u�4�X�m�Jb6�#���]��^O<��. -��A�����R`�ɦi]�01���-eW���+�YVlkv��p$`�j6]�!5�6�v��4z��K34��Rˇu�Yq�`
��u�[�6(�D-K1�3H�Ōn�[s`Fհ��]e	�k6��e�6�/Q��3hmԶ�)N%�U�iek.��i�r ��͸58n]���n��a�� �meFnє�S������V�z�k���\L�JL��Kt�q�>J�Rc`�.ى�����uɃY�@8� �!�3m�0�H�0	���eƢ �·:a�M�r�\r@-�^����"����"���8I!Aܧ�g�xt��8B�A,�-�_����}���ǧ��nݻzv����x������28:t������v�t'��嶠2�Q˧�Ƿl����۷oN����T$N
I�rBG(�8��;��9�,�������,�2#��O�N����۷nޝ����*���
��Y�m����%��w�n�^��ȲV�v�.��,�������o�����nޝ�����뎷S����j�m�l�,�b��6�l֓�(�m��ۋ�����K-t#�t	<�u��|��gE��wZ[��+��]ݞ�{fei�]���(��U��N�e�V�t���N:褩,�f[�\���{�<�:���vv�T̲�Lͷ~������i}2���mu�:�6���V�%�罨+��٤��Ee��K!z/H(�!:�4��đ�;Nݭ�9�Qm�-���ާ*Х��ڦ���^�^���o<�%�oo�8
ܳ����������|y��vg%m�K�;׶����Z\t��Zے���|v��u������;�I������.L�̾{�q[j#��;){YpD{c������o������Π�s�������N��iG>j�""��{YQ�U<�窫��]�fqpZ��M�;�1�ˮ1
�X9Q�1�b@8��Q8&���PDM��/�\���a0s��R��X�Bh�������ݬ�H������Y��(����l��K6�J$@]Em�JT5���rަ�&��KSm��hZmXb6�0֨b]5Ʃ���y,C�3�A;[�ґ�o!��ceP��䑸�)��BP�X�7 &�a�3Z]��f�m�,���i����Me�A0�;�b"�aZF�����mh�C,8;4��,-�nG@��--�a��J]cl�m^�@���k.Y��˒696z�k�P������,�U��`aoZڌ�1�6ڸv����R:Xc^Yn�Yr
.�`k��Ɗ�M[j�з�Ye��$��ѕW3WA���L%ѷ�_��R��t�3f͖���s���4Ae��e�JA�me
�K�%�kJ��d%�CYf� ���	a.�.��K�U	Y�5��	��Լ�CK	��@�Z2�.��p��ulq���7��\')��||�5�:anr��Uj�	[�I�:]^t��:1-�:,�2Ь�F-�]�\���6ѭe�YVj9�Ɯ#m[t�ʚbY��@34e@;La�]\��X�⊘�k&�N���J�LR�a�:�l��&��ih̒��N!)��Z�ݣ.�2��df��W�H��K����JbM�lkMh�
�(�T�ۮ���f�ד3L�m+�5�qX��6�eÑ� 2��f�jԆF���ri����SVQR�:��[XQl��K��kc4Йylu͵0���a�,	�����q,m鍳�c�¥Lh�֋�N�D��Y�bg�p��V�R�$`و�b�#�]c�a�t5K�)���u��U3�Aچ&�,pALQ�&4&LJh�˨��Ӯ1��+���4ٍ$Jj�aIQI�F��!e�٥`&���D��,��m�.��[�Jz��wwr��5<\��<E���s!/^��޲�+,"֭���Kh-6ƭڷ�Nb[(�b�B��)Z�HJT�F���Q�����*��%Z�ӗ��`C�Ұ�Rȕ�ԣU������Ջ+Z�ӠJ�H�$j����KH��JJ�rͩ:��J�A����\�?�,�p�z��B�
�D�eEdR£��6��m<�����u��s.�����򫷈$�������Z%M�pH'�錄o����Kd'�����VA�j̝L�T��@$�EU�zx[PN	(��1�ݯ8��zQ跜9*\TG�ָ^�Ҝ���*�Up6Q$m����1r}>}��.��@����#yy�Q~����@��I��apI;��v�eQA{����C6�r�	w��qO���i���_�[óz���l�ȟ$	�m!�5Qp\�5�C茋. �Z-� �8�m��&�%�]��52��W:�@�:7]�'�Vt3�g,���5W. Տ�H�T\��J]�>V�<��@�[�^"�pdId4����_� n夾3<Lg�@�S<3u��}�J��^ cg]�L�y���j�노6f&m�i��"�g>Q���q��c˶���YZ#�_�M����-�r�{z��־��Nݪ��;:,��Lj��Ej����F���f���_�������pxX}�+���^�%݂̈����+U��|@�T\O����d�e��[Z���%Ӡ��gY˂'�v6}�Ϊ�Lo�1p u�9FԨc�$��L�]���������~JAKL#�H��i���J��9�\�Ki��J]6M-÷�֚��߾��Q`,�
�GIkX8�%�|q�^�@�϶�C���<`>z;E0	l=�'}�� ��Z$cO��{^-�ہ��+W�z����DΓ�?�����"�E��½?!S�n" u��V�l̗���-9hT�5�G��׾���C�U%�۷r�=�.���w��<�s����2�={����!�v��>X�}����A;���tŝ;gE�<&5PY+���'ʞ�@�	���7�x���2w*���u�����rCM��8�0O�Z�	6j�iϭ;�O�� �X�'5��%�abuP�؍�������n��1Gm46�`��c5��m�9a�6�θ�	e��:Nĺ,3ޭ�ƸpI
r2@J?��j�,���Y� h�L4O�zt��\-��o&i�2����XZ�H�6�0�>ʋ��^���FO�K��P+��#e��vL��_�"�/��@ǎ:��!1�s��n�<�|��&��~��k�Ė$e<J~�b`�x�������=FSarͷ�4q����tI5)������q8�YfZ�uj�o�)��7���s�����Ժ���Frr&�L��"~��́�>��o�Me��<X6�S����`� ���*��"|��f��F�?�>�Xx�9��
i2*e��f,��P���Лf�gs����2E�4�Cl>K�}_և�L��o�=L ����l�"O��0p[ج������8�Sn�]��ܨ�i$%����ǘ >a����Ŀ�&�+`��N��
"�c�������{�{�^}%���{V4�xx��K-������a��%�{�R�M��#v�8���;V賲gr�.����Z�(C!��)�.l�H�}8�|\V����K��3���$L����H4�aM����������=�&��0zq�� �����̍��эH\�n�nf/[���H��Ɠ4ڞ2�d��沖lK�{�>�tX��C�����]�����ujY�B=s��o�����OF�R�hN���|:�Lk�.�g0,��
љM�@��v1�vE�Zn�S.���E��V�.�f4JfJ6����cc#6���2��D��(�MV��im�B�7�֭ΰD����5�a�-�릫��㵀��qmT
#���l�Q����rY����u#1�.� k�UΏ49�,��uСT4s��KL]B�a��-�%��- ݫ��ġ-�|��}�־a��&n��Sl0�f[��c�f]�j:�������W��QU��oe�gM����xߐ�3�`��@������M�R&Z�H����S�e��rB|S�8̢�{zȍ�U����"H��G�����ڬ�h��0�<���z�e%?iB��'��H0p:��R��UfA&��� ߟ�3��P�i��-����~�����
��vH$�ׂ��^�4����=>DDӇ ��}��Yٙ�EܽW���A$��dW�(���v�E��ۇ7䉪�� �}��cP���)�_��ٿ����j&�3m��/U�� ������e.��%ƪm�s��<=H�|��}�\l�[9p I�{y�/Mx�����Ƀ�du�`�?O��}�JMe�=��E�;���Pem�hoD3�NAsU+����k��W:����Q����g	��q�0׎��&����f:Ǜ����`�\��D�L��r���o
Ƨ���@�f���MF��1���C�rC�����5_�9m�}!��RZ�`im؍��|�5o /[K�s(ĺI����4�.�{2��'�0� ������T5f�?W��#���eL��'�#ԧV�v�9y��iH�C�̒w�^[N��YUc�#joHkYz�P����\3��2�բ�ch��Jԁ]����/
(��e Kk6������^��gfg	r�¼�Z��eo�x�N�pd��;'f+ϑ F�apI/�8�e��O��\��?=�������n۸0Dlٺ{����vH'���-4p�
x�G��~��c� ?�^�SG����e��Gv�o�㣦hQ��ٳNe�j��{�r����/��.�j����{_p���͝��3��h'�zݩ�g˂A#6�9-�!���9!^ja��Y��4|I|Z��Fr�9$���k*��\�z�o`b��a 汛t�EÆi�f�A ƾ@�t"���%:����}��Ēc`C���2u�4�xjfHȶ�v����Xr�\ ���)��#m����&Q���Yv��mɰ���(�o/y��t�1��̓��$g�a�L�)��j��Zm��'�����,�Bi&A-�3w�H3,LB&2�VW�<nI�8��J�f�0�M�6�'�?x�a%4�;��;���J�:6�g8x�u%��4Ә�$��C���m�y6��vvA;�dƪ�g�F>��Ppb���y#�';'�0�/�w���P3BL�Of��?�d���*�u����ڰ�O©�~��xy+o�]��-�5l�G��%&\ҰI� �Ec���c������oU'�帙¯��&�qXN�N8rA&��= ����^A��d�7@��}��I��[3�֚]l�V8v��&��m�m��nX�W��Y&i	~�i~ ��x�)u,��#�� ��������C�j����wc"2������3� T����,jh�V�cFS��1�I$*���	����׳"���V��H��d��Iܼ@"AW:��Vl��Wq�%P��kӈ��m�=>��L�̝��{����X�rَr���s�T	��A;m���Dl&05��ܴfs����?I��[��̴�)�h�����]0�F�4
�մ�@����|gU�n�
57U���ؔn����(����x~�w=��^I�v���C��o���qj%xg��8'�w��z�-ar�P��ɼ<Kb��CX�݆��WF�!�$�.�*Ț.�N,#.ʕ�RkI���`�e�l݀r-�{�C��,Eo+�qp�:j.vY�Q��-��`1�45��]C:�9��t�����H�T6%�jF��hVZ���,ņZ�;$�(ۙF-3e��[)�z����e8�X���T���dc������Ռa%%ײ�۶9�H�������y��_vFf�۴1�ucXe�^ra���SU�sr\��7)T_�(1e�6C��w��z��	7kK�Kyf�x�����zj3dZ/y���,���H�Ѵ�r�p�����ϡ��>|T�� �H�X��
y(�9����ހn#2�������q�2��DSl�7��Hi����-m� Aܷ���n���6ᓲwI'r�@�m���"1�a�5T�!�q�����66�k*�4��]�嬹$4�I$7��>R~����?k�'�I��yTC\9�>V7��A>'w\9 ��x'�Ͻ��?���q��,�}L���eE���q��I�.��v�]�\��I���:-���qYr"郒	2ē{�J�f��4��۸�ɘ��1%��%5Kf��	�߰H/�=�S��o��T��x�9��9�Q�=}L��.6�����h�%�wr��r}�>��[/{Jf����#}���"7a���X-�	���Av�.O���jˢ��4�Ӹs�(m�I�^wwUQ%�����`�� ���Ap���L^&�`��vE��کe�F<�c�� ��'r�E�"����:w�[�XdŨ.Hh��,�;���s�g'"yy^�u�7%�H|Ĳ�O�jm.�^�@$�wu����\:�Ǝ�߻�pab ^&�T,�f��a��j�21�ε�`�_'�|��[m���u#Z�q>H7��\$���{n�8�l�Ï@^�� �D[�z�NN��wf)��Z%5�3X��ݝ����`X��j�I������9���&:Hvy�T1%��%�^�L\@�w�$O�������h,�����C�
+$c<����tz�{��ަ/���z��	ӹ�VC鷸onw���v���&�V�����y�+�K����۝3Tbs�rS���7j�~�z��䱻�:,1����;��o��/sz�xw%������
LI�F�a��n7^�~�w�ދ~��ѭ���_�ᢐ�d��pR~�h��Ưyt�95^���]A�q�޵�AT��.�ܾ�$�C�:���/{<Wg{��{�V� �g{;ǽ7xf�������>�'?���|7S�{��Ű��٧V��w?U�,���52O�1���=�=x.�'����bӻ|��= Y�rg������ /ۨ��,"&���*���Il��=��;���xIQ|�,s3\�vg����z�}��G�y�����-��߯_n`e���o��KL'�@t��Qo�w�^z��;�n�g� 6����?	�;���a.Lm�Ϯ�Vڼ��k����«F+�v{ۨ5�w�ޞV��炳m-*��
]����Jy��|y����P����s�k��{6�Cپ�q��A>����a�nr�~������e��/i�Ǟ���|�8�rX�[����r{ݙ��_��
d͵l�U�o�`_h�L�~1�p��z���5����ڮ�u��q?�g��g����W����"���ǹÑ��V�A��E3�3Nt��w�H>��?x�g���7�*j��u0�hS�������1qs�:㎻뛽�إ�7d%%1�:�i�j��"k 0���2R���۷�l�����۷ooooo	�����QG8�|ݔS���BQC0L�*"ف�ES��v���۶{|v����������"x�-�⣍�eY�d\�Sfa.�"�v��Ԕ�wd�)͕Dx������=�;}}}}}{{{{x*(*�3)J���ZQ}���lI�� ST>>>>��_������=����{u�Dr E�G'QwfVl��q�Tw'=���*�̯2 ��N䎈�2rN)�s��ė��8w��rNw�gd�]�E����w�@Q'GNFV%ם�~�O���8�������k�:S�����Ey�Ǟ��ݞ~.�8:8H�){XRBN|Vq	Cn�S��@uft���ߺr��L)��]A�(O����u�s�!��)Y	�o�>hr�~zo��V���G��<�ކ>�k��w�����)JQ�3}a�	�K�c��'�3z��2�%�~|ך�wι�wָ�y͊d-!�:����Bg�y��d�ڻ�ww�S��{����ޢ^�$xu�:1�<��*�O�`"�25�w��:d2r'��hrYr� ��淬���\��y�>��5��p�$���:3����=�ăC\�,�4R��mQ6�Me`������M�����Z�VkVz>A�>q�9��:�2\ �7�[���!�dFBa�ލ�G��b<`+��PD�K��aFa��|w�C����!2O~q�C�����n�H��3�! g�@�:�@yx׊>�$C	���*�6˨���7/P���=����2R���[�JP��:�_1�fg�Dr~^��$x4E.����0l�G�w	��<�ǺN�%(��O~q�.�2��<JQ������Q��ǜ��d�NJd��3���s.A������I�@k~]�]�P��#����~Uhk����k��~A��'^q�g�>ać��x|�_.iJ�%3\p{�|��{�o8��8i���iڍ�K���%����=�H�QP��qI@�7h����w\�=�Jͻg��G�����c;	$Y>	@��xL�-|!郋�����'Ԁ�[�$5���p�G������a��/NFw󎣩z�����ﾁ�w�z��;�� �@�}��h>�x���t'��E�\��������C�Q&2�{[n�!4J 궦�We`GiKh�RZ�����~���%�pIx��=��z��f)�`�;��ԥr�dd�F����:��2z����}z������y��J��:!޽�9�$���峧%��ʑ�#�@���}�/yמ����7�Crq��rC�2C�<��s.�y����t��oߝh��R�.�Ǟ��n�/O�y�;�B~}}��.�w�&'O����Ē�Pd�'7֞�^��\�:n��t����R����<���G��R������Jd�>|�A��dx)�]�ݙ�`ɜ4�
>�o�[��Xs�_w�S!iL3���5rBe�&FHdb|��\�ԥ)OQ����>{׆s���5�-�\�$<���1�����ގ*ֵE��c�{$���:�tI�-	�d�7Ǻy'��F�S�b�xx#��#��z{�H�=\H�d���Z��R�����|׀G���;��"Z&qպ,�^/�+���3�y�����w�J��|V�7��s��0�B��j��5���ק1��`�*�o2"��g�(!ZZ�\�j�g�z���3?�-�]d�*ikKKF�tz c5��(��eaٌ:�4e9s�3����qce�\��UЬŎ*����Zh�`�^�`]w=��U�e��-��[]�1��Xf��ƫ��l[�;S��l����a�e�6�F�
iL�Mm0�Z�����u��f��̐��CBQ3���B!�2�`S1i3��WU��v����ձ5!��0h��_]$��B��T%6�*Xav�v�����R=C�Ю,,c��.wO�U�� �p�8M����+��08�d�I�G���藨2\���w�>r9A�5��E�5��_��'λ�T����FE�#��m)3�K1u$�	 �>w��'7��u�����{��!����T�{	��9|�9���H�~q�@��#�/:���Ϧ6yd(��U.�֩;!�9��{�Z�h�Z������Ϝy�'D.A�o���y��	��>�[�َe�N�9� 7��z��Bud&Ja�w�s�!�X� ���<��|!2/AdQLŝg��oH��wr}�1�ˑ�rl>�g����@dˑ�y׸u/Pa.I�����?:��L�������/����吏�mP�p�Ha���o����K�f,��8Q$xe�u�i9.%31L3���s#�g�����׮���C#��>p�R��@d��׺C �\�r�ߞC��#��g��n��x$��xp�Ԃ>�HQ�����3�2�ģ��պ,�n�C�Lڃ�k�@��Wh`���D<�{�|n���N��r\ �7�=���!����{�����c�>>�<-���x �y)k�i�R.��D���w���$�;���o���xl�-\�ח�4M��!���Qx�A��k�:�����kro�:�>v4�P��#��z^��d�S�]"��B>^K���$P���j��~�@"��j�� �	��G�w�-���ԫ�{�{Q�zIcR��ΐ,�А$,���4�óq�	 	6gc0!H q���	O���.��(���!�����~�-��McX��B��Z���mh�	� ���d�<��$��	=�>mg�`o��4%�	!���IƸPHJ��2(�bΠSR��"@d/�̖,ې�ͺ�Ӽ��~�z�%��
	&�3]\�PI��->�S�ZZ�=�l��I� a{���zͤ��b݄X�0�u�m�-c�2��ŕԢ��!8t�@��O�ӳ`Y�,��W�I�q�D�
�ޖ��38�����E�{ճMP���H�[p"�ub�t��ZBN��^R\��pǌ������2 �IG�fD��qwKH�)*���%R�� �=6����.��� ���G���e������ܧ�ܜq�Q�+g�RY�2!�+S��b�m>���P�S;�t�c�@v`ɞd��h2ޖ5�]d�J1bEZ֝4��'��1��r �� z=\�B$�Iu}=�����h�SY)Y�� �O��+���d8c�ޯY`�	=C��J@%m]-&����n��D�Tl��ls��89�$'�i��;%;�T@:�k<�|�'9cǙW1�M;�s�z s�Hxv�`&;�^Vْ��(���С*'��^�.�Չ'߇���-N��Z8�un��W kl�R�\�:lmm2����Owfs��p�)���Br�p�!�H��ה�I'�0�},��ZP�����;���2}�"0$��=��'�~+�e����r�?�h�E�=襐ꦻf�� Dc��$%
j�i�K�Į��P�y_�)�us��({��C�}uF�B�tIa*A�.���h$�Y�� J	p�с�'���]X�	/$�7t��%���n	�����k�m�01���ʠ�=�$�y_k����2^�m�	$�@Od��m4(����&���Ҫ��z����Ie�����׃of�H�m�X��wY�N�ٽF���6��|�M���ɖ?[�'ノ8���@44 H�	�љ�|u�u-�aE�q:��@W�R��I$֯�«ͷ���޼�/O��骒@$�`	"�[�;��O؅�SF���P$���\��Lv,��p��g��J�ܶ�:i�����յ-�%�ʕ������3��W�8%����k�o-x�$�9��}�$

����'-#�iCD�L�J����8n�'D$ɓ�R��U�Ŋ� WEXy�f'�;�	$Kz�G�Zw2��_���<4�m��vL���U@W�글Ȕ�e��! ����p��Ng������VT��J��ݭЈ�
AWZ�@NQ���@���.��y�ӻr���'I$Ա�̈�·%7����z(����Y5��%s ��!BJlF��\�v.V�ٝ��% �yS/1̺"�%��v,X������T��@ �6�3ɋ$YwKA�w��Pۆ<6��؆�	���=��K�ʿ{�7���e��Ay��7m!�{�
^��$�>��O�����Y�}]y��1��S�})�?N
㍈�,�@$�� 4�B4"4"q�=���sn%��ؙ)xmmՊ�5��թHJ�#�j˶�E�Ć�d�Wffi4t.�[Hde�cB��.�]5p�E�8�`ҙ���#@���S@�m؍јѻ��6��Aq+��l��kZb[��j�����Y�� �؂�h Y��c�IJҙ帹��lU�3k�ͱR��Mu�5-)�ɒ�];_��ꏝ��f:6�ij�Ģ������X%��(�v�T4�{�|��߽���F��$�;�I{e��y~Y�" �����[����� {|h�����Iې��e�;�.��N�UQ\��C�@!-�G�;˝I����I$���D��K.��{��ՠ5����
b�̩�;��@4�"���`�%����{�%�D�H.��$��)T�7;�d�;��P��ͧ�����zI)(}w�&A$-�e��s�o'uU^�k̘zqY�� ��	{���A�wvA�G���u���<�Y˞�y��uq��jw�gy���b|��e�˃2��%m�-2�I/f�:��5���w��;���a�d"�mv�%�Lijmv5I��^�r�����Z�W6`��>�7�#2����g %̖�ꗔ�S�W:'=[��6��x�Y��!��[���`$JOo��Y'g	'����WDJ���/Ҷ̤���y�<���Dn4>g�Whz=��5]��*Z����B�qx�W�0�����|�<���;��w�wY:�����B��"% �Ă� ҡJ�"�N>�̒���*d$���7s} (H��R4�{�l`�|�nV[:����Wa �ۭD�|�*�c�$�	[^I,����z �ZTG���@)��S�@�\�|����C9���H�[�E�lļE�xz`$�]5L����	���D���z�{_%�f����r�$K���<�k:b�N���t�!�	 �e���YU�719|�xo��E��-�T$�9�Q2�IO\�	�}����oo��N[����G(���ᙙYb$�؂.�p��m.F͑r���},`]ݐA��[�
5�TJD�.xd�D޸H�I��i��޸�#G�ĩn�R��K�׏��|���p��ñp��Ʃ]��	(�k׶���s�_sJ	7�&W͐�hd��/1���E%�y��k;�m�:��X��c`�8I8w ��U.��A%䧵�I"ȺU�ڥ����k}��7R�V�+�ަ���^������M�E�譶�܇�L�)$���L��ܛg"g	w�,J	}��D�	�p�P�qT1�q�P�D�P�P�P	�@z�w]�W� ��l���̗}��b�w0t�@�K���5�X�BK����$���T����W��^î�I)��@\��a����My`�n>�@1㔮�g!�0w�Nl1��1 �k�)v��ջZ}���>8H6�:�̐-؁)#�� R�]:j{w��n#�`�]y��Eӧ!Ӈ~pz�j �-i�u�]5լE'���}{�K��q����-���-�Oj�7�.��;���+Љ@$�� ��Y������#��<��-���@-�y2�n)�t�A�#� ��{ D�t$!C9"�<��<2A 	C}��d2^	/)� O�R\'��;���sj-�Z�r�ظMB�e��%~f �z�  �K�g�:W����S��B�E����f`=ę>f��MD��Jt]�z�̽�����;�-���P	$�!�z �o2A%]�Fd��U˝Eo>���*��"�0w���MΦ��p|��F�Y��w�{J<D%5�o�!'2&c)<�Vޚ��c�E��}�]��P'��2hA�q1�p�@��D�K��xyW� mS� ��߮�ӗw �P.���z���'~Z�;��X!�"]����pP
|�!�G�y�2.{�3(���n�>hK0�&jZ��N�/���K�?4i��1���ZV��.�F)��Ə6ݕE�{��K���ɉ�Y���~��BA$��ǘ�
I�kt(	^��
�^�]S�&K˳"c�}�f`���A´�*��4��_�3��@��%$�g��I47�0nl�ٙ �_ً��`z|R{f���NK�r�:���;U�/J�����Iw��d{�����`�6ֈ&BG1�Tʿ&	g.u	,U��ñp���qw�� ��n�+�/$|��_aBI$��l��Ӏ1�|��n�2���5S�)�w(���I=�!ṢoK`#���{��4����������I��!0M�{�x�/�����(Pn��bId�}%��=��W�F�����TN#J��w����6���d�b���>�ܬgz�������ڣ�W<uD��3�o�Kz�dŜ�9L���Q��؝-�3y��/��{{�q��V9j	(� ^���0�^�y��=w�%�۪p}�{��Bj��sd"�乌�;��#�{Z5�3�Ig鿯LX���6:y%sԍ��F�C�"�����:�۸�1�N����~������m�N�8y�o�K����5��{n6l�ӷ�L��d�(h����Ց��t]�n�yK��q��A��d�W�M1�߳�[�`ｾ���?OzK8��K~�c;��kR�Om�j�>|c/�9ޝ��i�����unt��Ip�Y<��{�}p3�P����J�&G���qa۟������ �?O�˽�{{�zx���~������ ������`#�l�f�G���t���F���Qs�V.\�/��;����{�=��_/%H�CT����>>ᬝ7��1�j�j\�i뉗��gQ�;%Ӿ|�{�^rמ����J���ɣ=Ζ�{��D���w�ށp��~~�*��+z��]��5Vy?eA�=��lE�V����e2P*qM�0�y��{��d��G��������Ǿqzѫم���ӑ�"���\@����
�H �H��i�A��b�\�)�+���D!�а� `'%?qZ7��bx8Y޹hUL�yben�4�3DW�O�ݍ���i�sp+}3�<Y |AOm�lrH)NwҴ��UMD��������������������UQD�Ms��Q�[9EA��v�EUT8������=�;v���������`H貳���6�p�&YU9�c���������۷nݾ�>>8E@Uy1'gbw's�sk��#�W���O����nݻv�����KJ^`�)YALTu9/�s�R�򳢼�J�:)�����.uiQ�k��IA������)Z8�ʄ�e���)(j���x�Ȥ��JC�Ȩ��e��ޖ�V�tQ��飒:�+:���e�r�we�g\D�y�u�y�<��0�KsWJ�q��w�<�bR�-�Z/����̤&Е�V�bh(K�i��E��m�Ma�AZ��l�"96�m�����%��Ki�\bS�a�l.�Ն)�ڔ�l�#D������m�S��[f�4r�.����L՗2�0����!a-����6�7�Hh�v��ƌ��fV9��ԩA-�V���+2M��U-b-�n�t�����@6�0��Lp��"�t5�h�/l� G1B�q]�I��s�h�%����,fe�0+�7 fYxHGq��i%�H�E�[����uֳ1@"��nq��Ρ�L�lj[�S	[��/3k�5���1����%�l�[H�++�VX](.�4)�؄�YJhL�E%��"��E���٣u�kC��4����+#���i������p�v��ce�j��&u��f��F�Ҧu�aڏB����:.[��q��t��r���-�#44Zb,H@�����Skpf�!�CMln���;<Ff�U�miLѤf)lT�ISa&Fk-��8ΖS7UJ6jjݝkY���]�	`G���	ie\5��cl�\�0�\�-G�����w\�͒�詶�фXZL[V�!e�ԥpB�v��е����]b�-t6�Vl�trV��� �����v�Զ.t���7��u����;04�db�,7�ZK�e���p� k-˱��XݦkKXKiPa`
��.ڙy��j\]f���CVaUiaW3���E�P�ZаR�����K�&��@��;q�K�Ɏ{*�XgFh.����TIx�,ƍM�aj]���ʚ���;Ld&&�m�U�FP�[�mJ����6��!Z�͒�)�n�rU�,f�%��p��J��К݀�+�-Vl���ST��ٵ�P-ʄ��䵩u��A�ηc��|<f�)a(XK��u.�&���B��q|�<"�ԉ�EJi��İ�"E�����"[�B�5dq���D�q q� �Q'TL��qEL�)O<�OW��n#�ڶ�@ab�B&#�&jbܵ�%�67^# +��8"A���p�BQ���۪U��^�Lg0,�(��Ymv�"����k�ш#�!�x��r�"40;i�E�ؔ��\�F$��UƋ�����%]��tI�V��X�`����!H����6����k��C1Wb�:ع��"c8òK�K�f�U3����>��ߦ���}6s��BZL�itԈDʆ�#�ւ�J%��Ĭk%�*��B�K�L]ܒ�|�6�?��I9�c��^v/=|�1)�U
�$â�O�P�߱A2W�С��|ʭl��X�g%Ģ��/З�cw;�Wf���-$���n�} ����gh��6{������(:M^��,�2d�[�Gg���	 �帀!Kl���}X�:��;���
C �kd(��[�$D�iNK�r� S1]S�̂Ų`��j�K� J���2A$sܠ:n�>#]�|����RJEŕ`�p�8MK�
��0#��f�D�7J.�Gm�-��Ip�
<��(�k��"��x�g7B�(�Җ�ivj8���x�۝�e�7&�-V�B�C"[W\ib��Bl�B-�dͤ�wE8N�஖�0��wC�R^��+=4����7{#�5U���'�i���߳e��� �+=l���!���OK'j�pXs���b�R�{LKbj!�]" �6�;W1����,��`^M��DvS���Z�-�gg
�Ӌ�H$�` "�8
��(�<>�$ҹ�dI$���=�T HR���Rz����4�
�mD�n{�mդ�˒�,]1�K��7�8��K��TH	��.�����f��0 '�Nڠ$�5v�!�Ao?J�,';�fp̙;��U)�q���D��	$�}ۇ})�&��@I�.�:k{���Jq	$F�y.�Y5g���,�,�e� ��`�}Az���p���Gl]o�gtvf�m�L$��}��"��r�R:��cj^�6J��E�����y���je��$���+���Z�J,7����2QV�0:p]�N&������D�7R�#���˝JM��;�Hhq� v��_��K����C1�ӄ]��;׍P�6�!��sn��m^y�w\9Ĕ30�9�Ԑ�%��>@��K�nR��'��ϲ�q� ,3�I�n��9A#�V�c$R�6��ˎ�d�0���p��w��Â���i?1^Oz�����������=\�wy��%�J����T�PY�r@hI�S$�T�i(������30�'�[K��U��� ���,]���K�i���m��<UX	 
·i"ZP	$�{[zZBD��:�'��.^}n�)	�zb�1f��j����D��u�p!���fM$��^�I ��햏$�Kk�D#�x�U�n�6	 �y?S�ɨ��q��ˡX[�%��sٺ.��	�Q�tû��{a��t��E�bj��PH�;��ř/$��G����=�u��]g��b�PL���[v�HIՂ�p�
>�y��U�{Nc�?l���|�������hIy$��E$����d�k_++k��Sy�Y嚋wI8.�d,���I _�s�L$�J{pl.Ϊ����?�}��Q䗔��������`���;��	R���&6�t���1I+�o��Q�a>��!"L��k���ߦSrݻ��,�H��U��w��v���IٰOxm�{Ø4y�"��)�ٓ�o�be�ʭ��3<�Ț ��� E%i�� �pW$Bq���)) ��-��?�H;7�ܗ�z�O��!�f'�mc1�3�^�roG����&����M���Ml���h0'�={�磭����b�h"�[t^4�f1�G,���3�p��$����N��ݔ�8G2 :%���I �I{9���[V�C;��Ɛ7[ֶ!��L�퀼�q)�g)ˇE�%��h��oTV��i9�f�|���(P܆�fo$��~�2�=Ύ����=�1;���<�dS�E�A�� @��Hz�RҒ^Ik��;Z�4u�jG�� ��ES3.��Pk!٤�wt���"��*�9�ܵ�y�	$�%�H$�y�f�t�@J����s��|� N{�%�0ǽQ�):�A��P@*�ږ�^Kcǝ�G���� $� �6J��+�-]�Ѐ@W��C[R��%J̚jUt݁rC��o��ܨ��޾,���f@�X�H�ܴ�>9<s�ۑ��d�yd(^����f^��i>�`/���{^w�Qk2+3����J,〆J$㊡�8B+@P���O��=jϋ�i,R[3�Qml�0�+���ՙ��Kc0���6n�5�m�j��Wv�%�t΃1��q�W�.����XU�a��D�b�m6�k�Zi��`����qx���K�!lu0�K\#�X�4\#��k��w792RU�m`��/+�j(�ݔh���ꝡ�iY���
f]"�2��s�k�xte�>��� yc_L �F��Q�P�an�FQ+�bg\Z��l��V9���=z�S�̲:˹�vo3�.��k�����g�)$��swK�{L�7Tb��H���W�M=��wS�vR�M'� b%ɶ^���b;l��FÈ�!���T?R�]�fI{Y��$f5h4<f*��|xe2�vr����a(�J�j�&<����$�։ٷ��H1��UH���o;@I�xڰ]�N�P���5cַ�r�q�PGs Jm����f>e�;��y	5�:ޘ[�b�}h��^@7� ;��ʥ!�f��L�܃2�*׃�)%�9�G�"�lȈg.�$��-L��>���	���o.��c����p �&����K&"�$�ѵ�f��r�љ7
�h�
?Ǒ�y��CJm>��׺DC��N�;��w7�$�6O��$@8w�0�I�� 	td�DCFy�V��y?� �.�h�f��c ��gr\@��"���kl��"w��`ׁznk��s���}�=���}��g��:]zKN��"�j�N51{�_����PӍz�o$N��rn�����i��e�G#�
̊ػ���KZb�2�������5��j�Cn+�eJ�bE�M��>N�t)���Q�$�8&BR�S�*� N8��% U�
d
����{�u6b�~In2� y�$�5} �I>9�k�.��Jy�o�����r�ʪ����I.�q���@)ykKy@~J�8��Y�/$�v�@@"N�8�	z��jwI�9(����Փ�5�y�q�/嬜ռ �|�f�x	,�3yo<Rݼ0]��CP�0ދ �I3����8qˍ"�h+�}p>�>����n���v�ղ��n.���U��t4��K�`@�RH-��@H��$�
������3���t�J�n�0eKc "ij�ً]k|���n�%�?�_��y"@�����Iv�Z��k���G�[�pV�!�$A]�0O`��3�A'r���e��F��f�*cU�u���$���L$�s�  �	q���۷�n�H7���ZAټ�一�oa=0�\�y�y.ƺ��䗐c�ԍB�۳[��>�u���]٢8���@9�X$G���ln�3�d���V3q���	����^Ό�sq�Z������>���"c��
N8d4"�8""�JR�0$��y�<}bI%��;� K��H/���i�� ��r���^����ĩ%�]�ª��ی�O���$�Ki���!.;�ӽܡKC��3�	�ӦO����d�Y��;��;�6R($M�[V#u�(s���%rI'*Dϒ+�%�t�QM�`#��zIۥ�;�"�	�h�A����L��iD%�5Ż1%xkX���&[V��]h�3�$��E�'��e]�|�.BB|�Mcu�I( ��}~���פn�q-����	#����D�˿�����o&���H�&E���L�ދ�� $�Iu�ҙI,f����!�%��__Dlq�-��+7�S�.�N���%8�r�|�) �Ǐ:^H���6��[�J|���ԤJ(��;@�f6_� ����q 4���u���_ �	���攀I(�n�b}^2,n����ID�f���쇼��Q.�;7J�ҍ� /r��L�P����,��E�}s����8m�s�>��Ӈ]uk����da} 9+HOӊ!�8��%
�8���8�� (4 A% ��ј
���@4��;�r���T`�O~�HS068�.�ucj�<��&hu�o ��I$�v	*�0���SB�������i����@)cE'e�3��&+
4K�b��h\�͓9s�|���j3h�T��12�;�i>E �׀�$��]!-�<6�&�&���  �Ir톄��F�BæEó*y�ňI{ɷV�[�C)�G�v4��� �����lh���ؔ��B("�\l���T�����������&p\0w+�C��5�̫9�Hy �J:�������y��`��9$�̺��@
���rΝ0)���Q����3�~P- �@.5/�I��Dx���3E���;,���j�^�{�˻@�30,n1����q 1�\X��Iv6T��1駥���\�d�v�t4$�I[��0L��Z�ԦU]�[���L^��>T5ං�M.g�;lu��߱�ᘉ�����{Ь��~��w�i=�&�|��޳}hAe9m����	���!8�c�*�N8)��E(�DD�'��ϔvb�h��(˴�q����M�����m&�mM�ZR;1+k0��Ŗ+��l� Vb8��i�뫄�,s���!E�L�X�6"��к��M�n�Rѥ�k,ku�V���DRQsl5���U�̬YX������%,��R�uՒ�V�ڋ[Z�ĺV���a`/:��b����k@S]��J�S4��K�R
Y~y��C֛�فU-Qjj���V�a�e5	���]����s�}�?���9A�ҁ���~`���`b($���ր�y�9X౧2���-wC@J|�L�@�	y�X�;���)�*�]Y!��Tr�#�3ǡ�H-� ��FH�	 �[�Ԁ��0��7�F~�˱�	?���;	��6�0�1p�*��@D��Q�ƐS���%�^`X�Ç�$L���@O�\jr�:g%�a臧��AF�
	$�)Ø30�05���������q
n��k�� 4o0f@-ڀ���40t��D��8ӌ̒��؟2���;��q:+*@[�G�o !�1��Q�$��n�@5deN�]�LR��0p�μș���,E#�M�E�c,5in�i��O [}����*�d����p�@$��6T��W�[����V5c[��ma/���Oku)����۞p����z�O[@�K6AMK���nG���v#�ȷ8vm�E����G�W������_����v���g�+}�mDٗ��$ٗ�y���<��ם�*v
3��`c�8�#�8�%ЉxG� *�}�	o�����Gj��>�y��I�$4յT�<1U];�LY��	.J�<ĉ>��q �q�)���7.,��67��I�t�#�����G�-�а�Y8we#�I=]i���7Y$���r�3�o�	��'R=�爮�C-���tv�B��s�;3������	s�"7u�4�3S���$�؂!�K��5M��g{E��E���vP8�H`$�gᛦ)���f�� �R�h�V7[凿�>��EY����������]v��WD����S0{s��]�wz*7�N��p�f|g:���u�}N�B�X@$����ω�}� �D��ڋ�kl!I:�p������ߟ8痧1�<�<���PB�涋䙛�����ȶz/����Oa��)k���OLG���?@Ø����V-Ěs-��ur303��=�8���x��z�Ip�G#}��~^%����`�=��/�c��wȌ�z�V���.Z{Lߌ�l�ݣ���W����WU ����w�\G�{o���9��>�	����:������}�t���\�/��v����<��d$����=F�?R�%�=2�7��,>��y�g�����p�z�y�z���w��{�?$R[�.�r���ؘ8+�o�A�.���̱r�_�\����S��4��d�������-�o'?m�u�W����+͙�t�3�x_�n���5���n�{ykUg���B��������$8���;{.�/�ds���g>��P�Ohr9������{s��f�gz��o��}����qoP�������h��G3�`w��u8�����M���c�������g}��V��>����r�5����]�K��G��W��&w{�n�����}U޳d��ovm`v!2����������Oa�
�K�Oz�w�D�`��'�6�Z�]��S�$��.��MG~�Ov-y�"�3w���3̈z5捴x��J]a�.�1}|/��G}PήM�i��&}���{�����~oP Ql���Nv�G�Z(���Ǔyc���zu�pa �,�<�FM�x�
l�9!�ق�����εɝw����`�aE�C��GG_ó�������������v�۷oo���zx�k6�<��ʣ�듣����ݻv��=�;v�۷oo����_�;�8�J����Y�+ �1��O���nǷ�nݻv������ePt������=�tT��KEo2��2�۷�o�Ƿ�nݻv������|`SUIAF칵�]�y�;E�t�5�y��PQ%��tw}3�:Dꊾ}{�we[��8����.���J(��)����u�q�_��tI�뭮+�ͭ���D�ʦS�2k%���q�RwQ��i�� :�{q\�	�p�2hT(R	8����aIw�x$���G�+�X�bgffrRNĊ��N�}w�/[��9�O ��Ȁ �3�R�/!	ͱ;���mE	�@v�;��@�97�@�ԔK��J�3I�q����q 7WR�Sz�{�})��t&f(�.����7&���6�$txXغ�16J�<_���O�.+;7�%���H��1�� �?B�ր�}���yY�� ��k�
SL6w��át#�UpJ�D��E�E�W<�$+nb> ��H@%^`m���Pv��k��=��'�	]6 ��<�J�i�v����@$�ޛ�>�]h�$�׾p���.�Ȋۈ�0W[73r� �t�A$�t�H'��_E��v�+��e�!b�L�~�N��P��T�l&ځ!���tڴ#������R��/�[L1��]^)����~��3��+	HN8*c�"��y�}�xă7��Wܠ������I;�e�J~S���A��3�o���
������1 �<��	$g_D)���cc�h����T��2E;аNc5זX�,/kF�X�kX۶8��ݚ�vg�>8]w��>�Ig.��w�x�V���X�U��oHξ��8ǩ�{�c;V�	�Ԡ�|ӅbvgE�h붸��	v�.����ua �I��m  �2�f�@�SU��{ۧ�}Q�z��[$�'{��Ҽ#��q���W5 ��Z���z��{����}!�f+(��0,�;� Ftמx�zH�t��	#�2 g� ��L�g�^�%^�~�$��\;�t�� Gm=���ژ��FZm�]�A�s�!���	��p/�[��*�;�Ir�]S��8�W3KM@�W9��6&�厫1o�i��IyO����-poe
VE�y	��a���>I��d�.>��?Nd	8�d�8�.7��<~�D��	H�{�c]ڌ��Uj�M.��F�i�.���Ƒ��KIZR�lŦe�ڰ�ڰ��0D?Ğ�M�t)�6�V%��+���0�F�f6�4me�9m���fg(�f�<4t:���3�/;�͈j�R�֝��vۓ(L��Q��:[V����&4fи"���m�)�ш�MS 8݅���R�U�M^2e��&`��h��v��JѕdʙJ쀁�5k����˨�ϻ���t��IIс�{�D1�$	�׀|ck��zd�ܩ�-��R�ܬ�1$��^{}�r_a,�ݓ�+�%^�u�L;L�L:'YL�A���?���do��	�y���6*����u�/k�ZvgL�i����]�Z��@!V<��gGv%�yW��ΈB �	WSי���IwI��N��χW5�ٽ��Z�]��k��G� ����D�sِݝ8ë5�
�؀[Ȏ���'�@��T>'|�;^� �ɺ5�(����h_�ot8���nL�g�-���^2�{��]�−�W���H��������gK���8t��U���w$:wd�2m��{/" wy� ��j&�sy ձ/g�%��Fr�O�l]��NLI����$ǀڃ��hn�-N�"���+"Cȥj%��|s�HaN�s�ӷuy���{�꼽��n�yo.7N���s ��O���#��2rr�y�`y(O� 1��'L �q@2�`�&��� Gٳ���Jw���_�'��"$u���ӻ'vS �@��D A��@>����mM�Nȶ�FX>���	��^ H��2]��:tX;!3��&b{h~w/�����0��oSz(�T�C��݇i�ϒ׹� j�v�vI��N�:y�<�� 	[���ǆ�ި%��\�H�ֺ�4�·����ϓu^f�:�i�U�+�c7Z�YCj�
�^)X�����.�M������'�v�_^Ϡ�f� 	u��v���XP�6�]쿰��z0	��w.�d��%z���q���|z�U�a� ��K��}�>�:�����Y����[^�M�b�22t`U����z��"7t�ws��������q2!ĸ��ax/mLVbk����Ѫ���=4���>GCx���l���ɭ��1,xlr�5J�x>��y
c�"c�@�(����Սd��}��@��m�� �e�n2��ӻ'vU �@��U��"�M�"�5�$	�$���> �<�4�շ��[3��I˗��Fͳ�ggE���{�H���|�\Z�;�Ī�ϋ\�| |:�b ��<��pDm"����8������7%�][���X��p�MQ�n*����<��B��w3^%}��r]�ft��$��7X�`�B��y�$������m��$b������ ����$�+D���d��Ȍ�.��v:]���v'#Y��w��'ٛ1>>�~��q��\��w��x�+��3ɜ���]�<F���@#�E��<�ٵ5:4	��tG�'n9�_�[��\&v!��R�n��\�e�Aj�x�$�������mޜ��B쐝♖;OX�$�v����,�����x�l}�M�d2���99�x�o��NZ5�,?w/�Ӄ]wގ<�~�o	�G��7؉?N(c�&T���	8�&HC@!B��箹� ��;<�sL���P�@�e�����Uڶ����#Ḃ"l^/j�¹� �oO8���i��,�<��N[$���Xӽ\�5�f�npR��ÔF4������;Q��k��aD2wr�����d�Kn��q4����I �=���G;c�Qݑx�r���	�Gh�b��$�2z�^	 6��n�6Z�i�>���	�P �1~��s
���/5�1�3�,�;����~�3��@k�̫m�,[	U�}��������	я65w)�d�YD���k�ע��BE�D���� �F��.����F������f�� �u3q!q�<q��Έ,���^���H$�����w��<)$u�G����������`�/7��Y�ɝUb1�8n��uf�����1��.�"�ݾ�
g�sR:�ZB��2f�{ģ���bZ(`���d]��/�����$-��q�t8�N���$�$��߭�$�ؕJDFb]�\�L��\��8�TS3�Ii��u3T� h�3pʪ��$aY�n�M�v,$�,�VRX:kT�+c)Ⱥܹ1�I����0lQoU��Z���[N�i�Ĺ�ٱ&�7: �ux1��g�J�]xP�lŋ]k���M40j�[r9Xٍ�.��Q,6���SG\�"T	N���B���͏&�򴠹,���KK�˪.�v206�jZ�ҋc���D�Ch�j<�;�gv]"|���tD��įwk� E�����^�& 3u@>*�jp�;���X>��q Ե$.��aM��3�+�g�Ws�N�tG���]r2qVK6<sf��]1fgd��H��@�|3��9�'w#I�����0ϠA$���  ]�MNCS1�3�,�;��U+/�Ntm\�Gh���� ��8	�$�}��-��z����ף�y��0� ��D�w(8,�R��ul��@��� ދ$��''���^�ȓ�}]�!�=S����a��#�F�81v��ٍ��V�b��vDm
77f�G������g��3Hd>���^��<$�n�� H����Q�L�3MUV����=�����|$��r"|�|��E��3�)�_���!�9��}nv0ͯ��t+=�G�ƣ�ط�yO�O*��}��I��}��y
���[��[9E�������vaY�}!����&S�&8�d�%4�BI���Z� �$Xϵ�AGȐ~��z @l�k5B�{[{jp�;���Ӯ���|Ӌ��9�a15LD��Ӄ��Gv�@� #�: �*�n��,�ٓ��y��`umAw�17���P�I�}x�'��B�ӷ6/!Gf�g�z`@O�Ǽ����v2�*vz#� �{&��{Ta����=�G��Ny"|O3��@��<���z�?g����>��A�f�4Ȧ���TH8!��5[.y�U��h���-ߵ���,����g� Aݝ�E��x ���cc
�ъ`7��<@ �U�]�1.��92���
�Jͽ�
���	��qpOw[�A�Ю�۪�T�6�;:gfR �_���I��c�$*f�1�j�)	�qt����=�`��Kd��^YۊQ"b�:��#j#(!0W�h[�=Z�>x����^c�~��oӂ�����\T��e�7�7��x����mg,S�(;!���m���[�@��I$nƚ j�!���dw��h�^��E�	��.�2v.�*��[�����v^���5�^�ܩs ��{�$���N?l��sv�O�NQ��򇢱ڎ���+1F\M�L�L2l<����C%.�e����v�5�?8�˦�y?t�?�kм@'wZ�"@$���"�f�ϣ�k���_żM�= x�YE&�H8,�R��ulA�x�*�dmF������{2k���^�v:����+�o!YV�܄�N��:��<�'�@����D/+�8;�r&����/�K0���ă��@#_A�''gN�ʤE�ۅz�6� 醘�@9w�|�g����.}�6�}����P����k7�3O���t�j�a׫�{�*TB�s���[��(�XXC�����>y�g%�}���8.8�S��89x�!�>�|�*,]��B���A �8�@�j��u��Lk�@��$�}���S�z5�EO���t�;��8N�V�@tn�F�h�,������K	�܎�"�>x���s��f�'�;�_59W��'���: LGq�l�����f=�;5�����;�gfN�d�9=2�'� lkA�W�{�� �}���q���Y�g#P�+�)�&A�Lckb $O��|��Q�[|lc]�9�Q�c 7����}�	=O�r�qTK�܄�L	ʬXxc".�^���Gt���$?��f}�H�����bΥ�M��"p�8��-�w4f~������j��~�ےc�"���o ����1ˋ{�� ��Sqoq��15�U!���o�@u���,}�t�k��ӽ��up%�_.>H�ȸ��QgF�}�;=x�Z�����e\sn�|4����d�"6�{��у���}�M�y?,I��|Z���$�0e,���g�=�j�s���H�����W�2�9���5dηr{�����|�yM����|����)����̈�܀��3O������<��W���۪vw��a�pgDm1���{(KN����w>h�g�E����{B6-�����q>�,o���~+]hSG��ERS�}�zg	�97��M=L������8$��s��M�Q�,�'�S�h�1��T'/�H�C"�q�#uV�u"Cf��4zK�k��=�	�A�.>�ge��L��`0?z��f��h,ܾQ{��ӗ_c�+��;�zh����]��ɸ�#H�:��{�bQ�E�D	~�}�����Ȯ��sr_,�N�)�qq&�|�k���N+�� �-^]�O������|rl��x�1��w�M��G)���/���۳�AU��u�-�!�L(s7�t���^$r:��U�f��޺�T���vzw>�~�鏜�����X�
={�,�|�rSpc��ެ������­�ǭY=�J�Gu��cd��x_8DWv�]�MX�,�(,ҷ��:�_Q���,�n{|��s[s�� ;�x�:DNmI8]߶�{NxQw�D5��gr��+
�C���3���"����>�Ft9l��!�9�~g�5�����cX�m��_�=���Ӡq^�))waD���NF�yg�`A������ݾ>3�nݻv���|x!"�;�+�Q���I�����O��l��۷nݾ=��9��]0�5�ʚ���T%4dRd��K�����}v��ݻv�۷Ƿ�ǁ�xURAUD�Hd9KUNK�nݻ}{{g�nݻv������⢷BwDPAY������N��N��'qȝ�2�%6�]�'��m�{gI�l��*+���F�y�u��(���Ͷp�pyQo>�U�V�"(�㬬'��-]�h��-��9�Im�C;I�u�9_�_7V�t�'s[ŠB�	@���T�{^ntz�����V� L�K�h��FV��l��Fia�-(��c1mp�G3
j�Q�ћ��v#Z���GF�4f��)�a��5�ƕt֘���	H�okZ�+&�[��mXVQ��<j­n݅�j�j٠MuX�V,G"���S[K2�b�h��-ʍ錃R��b;J�ch&��k8!r��R�Ii��!e�+`B��FӁأ�ٰ#c-���e�a2]*��$���M]��Z˘��v��QlV'm�ѩ���Q��6�Zؐc���gʖ��liIf�3&L�X++6\�]M.��SK(���.�J��6�b��65M�ip��6VY�),͖�p��59�4^��:�Q]i��H:Д�&L���<qYoj8�t���^qKV0��bk-��u�tA���q�b)6cYH�\1a��Q.A쬰����P�f�R͜Im;!l���lvfD��\�J��1�SY�&�cT��Zk-֏i���a� ��^���1�̭�څ�yɈ�n+3��Y�B�`XU��ѹ hm0eښ�MF$i4H�b��Yq%���X2���X�+e�m��5��eƎ��*�&�M5�SX���ZqarJ(��U�Qa�T�˺���ښ��A���^z �Y]t�(1!�my�X��a�ch�x�J���cX� Y��r݋��p�e%DtMA����sfSKtt-�h�m�h�C\�e�
^��+��	b�x�1�4��ņ����������� &�*rS��6�2e
ڛa�m$�V��؉4efmQ �.��o\Rѹ�Pl�C!HGJ�;Z�PH�{F:i�d�r��vјI��y���l]H��X��+.i�a[���|Ec��ȩF�%���+(�ub�[ڍi6
�Fj�\�Vmb��g��G�-T��seVԗQ��J��sÜ[.2l4qc���C��`U�*ٮM \�jD0�օ5K]���� s1Y[��q׳ac�c?̝����;q��&q�rB�������q��jk��]���hA
�6	�-�4�sv+���ݜ2��Ml�&؄n*)�5m"M�Fi0�%+�
7FY��e�av 9�Q��h�J�SU\�fnmD2�3flNvD���@` Ą���N�-�T�h`wl���i�M�ImSL�֑1��W�h���L�W.�fvոfI����3babEmib��]�o�Ʋ���`��=P��JK6�R��Ko:���	�h8��R�O��\�,���}o�[h�: ���Ԡ������	$���/i,����$���6WE�������>�ӯo��vz ���J	$h'm/ 7�a��-��k��ٙ�� @������)���Kǐ]��y�Eo>+�zI10�����@�n�!e,y.
`�ğGmƨ���?��Q$���A�)ucO�vs������羢F��� `�\m�;���q"96*�l�_�r�t�|A��xd�y!x�j>꾌�Ԛ2��*)����ljŤ�M5����r��	��A+��dk�3v�s��|�E�]��/D�t��ݙp��Ȁ3�J��e��I�� �x�g^y��o���$��zPHk�L��]��F��@$��A�샅��>�r�.�uԝ�vɻ{���F=��Tk�m螕�cm������%��Eb��y��껾W����U���~�Lq��q�r#� �	�u( �_���Jq�q�k��s��\��N���p�2v��y��7ۏ�k���Kω�X'���}�N��g��\#�wg.ɝ��Α���ȋ�p'�ő��<���$���Í:36�	�j�t�JT9�0tb��
ީ�I5��2k����I��}Io%����+B|0��wN�ָ�e�*B��]��\9]�X�M�.��{��XR7f&0���rt=����	����*�fWJ(��PO�+� �w�Zɴ]ػ:eR��TB�@��wS�ɀ�l�װA� ���B"�@@��ODevrJi��z� �z��.ΊӒ����D��1]

��2pl<<��6LJ��R�uԟb��flkKHM��௰1Wẑ�(�:UK���jHE�X�-A���������]�E�re�y����#[��񙙙�ۿ���ڈ&�ٛ>�k��Мۥ�S�fN�M���.�awa�S>��A���" ��-��IuKonS�*��OTH%�5]��&v36���|I�[p��1�w�(%���2I ��@�w.� ��}��B!�5?%�
]�tj�	!;�r�]�9��箱�c��A�͹ �1E��co}�ϩe�o��%0t\wy^�@$o# o�Gku�<ͣkn*�$"�����1 �	��x/�hu�tCyӹ0*�Z{Pc5�����V�L��{��Iq����֞B
��{O���"��{<l6��M�����)�=Ӂ~�"�O($�	5U�@9پ#|{'�@+����$�]�f���:(3@�뎋�5�&��$���I&��|��=��P/k�_4ۻ^�RHX��,ƜH�=9�֓o�ao�}��
��ࣽ���k��9r{Y5��n~��5�8�ɨ�h�j��C�W���� ��";#H��˚�vb��ü�il�bI7ې)���z�ĉ��tߎ�!.֋P[�w��eQ����A:�Jvb������m�L0��Y�,��j�q�0R��-P�.�O�ϟ)�"��gr���p
y�I1]@bW���N�=�-��F Zr��B���������K&!�`�Uzz� ����k�J�q5���A{1I �w< H,A:�7u��NH����_�<EۇD7�;�Tr�^���{_\�� ��ܭs�<Bd��v��	�k�-���1�'p�E݋�v2��*�wot��s�>.��I3]��O�#��2�Hq�B�B<�������i��{�5�񬎈�ڼ���Y��k[��z �v��,Ws�.��o�0�
!45�=$41��1��u۹=$�xb�} �<�3Ք��K8�I�c���v����co�6��3"Y�3���+=�>> ��ס�҆�cSg�F]�R�B��3K0�$���Y��`�m�a,%+l�Vhl��|�Ķ�Fj���7��P�$KpjSPXcgX��W2��0��u�)f,��-1��ц���Ye8�%e��M�2�)�Y����j�*ԫ��2e#�ڨ\�0���0��nxv4��n�f4�aG�a�"ŕn�ݖgmo&�،��Z�lQ��?^y�n�E���1�0��3kjK��V��7��a_-��e�*Ou�:��_�~�t�E�m��%��l�7�gd<q"G\t@�%T{��#0!��@'����;U��˻�Y��Ɍ��ޅ�[`Tq�16��F|�g|�H�;�� $���H^5}Yi��>Td�>0�J��!�`���z� A�|~���IΗ�fX��yD���(�,�ي���0m�	;OG�]�����N��d�Y��_����S�<s��ȂA#�����]���͆�A>�Ύ�Q��6Rwr�;�|2-�!yO�r�����Ǽ�Ct���}I9˩@�-�]�ۆ�ۉ�Z�C�9�L;;�v����4j��Va�@�����X\�P���a#��鯞����P�L���7�꟠���&v6@%�_�H�FQ�9���f����D��3]-jIيf.�U�� O�|���m��B8*oipP�?)�Э�n�(Z�׹3�o����7�"�	�.!sizp��L��`��L�pUյ��S��p�89��r&ff�~�]�A��؂|wWR�	��|���LED���]���s�FZ{���eCjk��j{gr�J�Y��]aa��AX��	�ԁ�)uLC��ѹ"z�:�F��P��	 �M?���-��a ����4�
;+�� �� F�q����ܘG����gkߎ\2��"�� �Ϡ�W*��H'-���~`���3����oa)�1I�t�$�Fݛ(\���Z]�-V����T�.��o��Sm��X��wr�;�V�n^Ibڀ���olA/1C�dj���Q�x��4��3�p�'�"<	�=����%�v �5����0H7p)��c	Q�q�b\�椙��b�݄I�]J'������헯��7q��0���]��y��8������
 *�k�`%�2��q��p�%��͉z�N.�Zl�:���b��'�Ԛ<�E��`���-�h��6�(>�3�?����]�"��`1�Puֳ!թ�'�Է]���C���d�@+Θ�],K�q��ΈpB�K�`��`����� �fD7I,��[ԉ���x������b
���m�"���*��v~�5aL1-F]Ķ�(�nnф{j�R�L�g�k�yӹ0;�5Y�v��N�C�i�mv�w����X��!{��!3�0h�	3�L�Ƞ�M���f�wv}�γ�ܙ��x$��3WL�$�nb�=���ƀKMpcN�2w.�']���D�yy���w�Y����n<x�o˯�Ϯ�
�tY�&Eüv��Z�z�FgF�[�$��x$�W���	�.����|�Ҙ�*�[�7�x��Mp1��*�Bk����h՗�wK���u�kR�&�M�r�{
�ވ�o���_~��g���~3335���<��s�秦�5�gsh;�
��SS�X3���� fߞ  W�wT|��b�ʙo?���}C�P�~ѳurB�m�lD�klY���F�-�4�5�{;U3��Z}}L}qc�3��=��x$�GfD{�Q�A����l*��]��I'��=�}L`w$7�3����c�N�M;>DuL˽�I�=�$�[��
�b����{�54��{���d�4v��:,��d�VǠ�^Tw��׉wtK�&�KE��Dr�\@8{�����Ɲ�b�\3L�tD�v�n{U�Mtc� ᫩�ψ���`c�o]KC��f}�!ߍ�2`����D�2{�����ۂ9 )����G[٤�����|N�ڇ$�FwdO�䇍g˞i鷵i��c՞|���tѳOCN�t�?����Y95�݅�*�\��_���M�z�$2EY�}O��,=���r\\'9�q�E���~0d��'�����@�m�%a���6�7R��]���Eŵ�]��\�j�c��k�
W(9\]�c@��M\	6ֈ��)
µm�[2��]eiM"�u��+c�P����T�����M�����N�kL�M�,mœ��-[�����es�����6��8��Th�iYx���6�%
�����t3vЖ6�|_/Q�mK(˚��(Z�����|<`yOP���d��#�s�yNէ,f�,��T���שv��?z��F"�,�����q̛r	��{&N<{"Yݯ�RoT@½�v���1r���L�^]]�z��ђ��u�f�V��[�wvDG�ǽƔ�?q�n5S��J:n�8!�]���R��Đw;^ c�)�յ�����k�&�gݼ� _��7L�����ʕ�k��%�k��|��������s�m��)c���Hng� w�����wE�85^׹��%�Hz�O.����� O�_�O�${��"��'ǯ�#�A�����?1W�i��eb���Kۨ�ר�h��m	��+������;�L2p�Ӄ�[��1 ǒ{q�A-�hoBYx�����Ct�_��3DP������,��'��uG�m���r-5mu���F��IR�e�0��ΫC���չ�SY���/"�Z��������������ۻv�ޒb�D{��������3�9|O�?}D H9��/��q��͡1U�˽PG-X�:)���=2��	� �d�G��iV��p����k �EotW����� �ࣸ�bAvpXVz��w�@AW��%�: �A>�+� �x�CDI��9��N�߭�&Io0�',$�8`�hP��=���ި�wƇF�s�1K�� I�ɏG��T9/��7d̫u��������5�nt\�etQF��)�YY�^!�˒Z�U'E ��W
�!�h.]���w�ix�7���ػ����⮊h?^���L������(<-����h�v�.��}e� �D{�f@�K�n�a��5�3����;|�(@�p:<H�y=�C�w$3;��n����J�I�$=��O��l�f�(�Cs��%��A�2�!�ƈ��Q.^[�0��/C��D?)�Y�(�0�#ϳ�\�渴��-����B�Y��������ޖ��^���ʳ����j���ɴ�_k����&/F/??m�c��䘎=�ڶb�����0�:1��nh��}Pպ4m����w���e�*IƿX��O�~�1�L��z%3rS����Ru{�v����1|���9�t5V��{Q�g+�4�x��>�^��bM���jX�K�W�L����y� ^��]|�3�:�n{y��>�Q=8/�����Ӆ���^�'a�V��㈜.?K�;�b�{	�~����;�y�i=�'�Δd�7d�󰘾��Y:g	�p�Nŵٽ����=����"&4��qR�fw��$v3é��7����&�ǟ3�x)���3��Jf���b.༛�7;��\;X���·���{|�W���瀍E���ߞ�%n{����<b��+�\�F�l|�>z/��S����{����7�+ֽ��{(S��׻�rUOh�������R��._1��}j[�<��}�4�b݁jP�`ǜ��0��þ)��1�=�u��ݼ����@�����%M��OW�6��6;�!�r��R׮��W����|�.��<=w��J�S��`�7p`f��f7HEx�q�/gOi��h౓���q@f�B 	Z#��y0%�\�y�&H��� �����C��={Ғ���N��� ��N�%�yM��9r5D����f�ό��Xv��%�9��+`��$���P"|��M��:�t�����bXn���>"�@�?�'Ŏ]�鯴�����LNH�{���{������;� ��X�[�O�Nd�9O��߿>\�N��%�) $!!	-�b�Y9Y�ӷn�^��۷nݻ|{}|s��X�ẒY�AZ���8�0�̜�
 �۷oN�_��۷nݻ|{{}x�i������m'���o=,��:(�����������nݻv�������_���[ki�B�ݡ_���`�,j����2l�"[�����nݻv��nݻ||{|8ujx�b������;��N�H���j_6�B��9	Y�QΝ�6� $��+e��ٍ$ߏ{�8�H�͚kYpۖnL��~���9�L�Y�m�cTGqYkk
�ս�����/-^ۣ+�6bÈ��8���*-(�2+㳶��2&��6�,���,���b�ͣ��������fg������w���y"�����I`���0gE0."D��(�����I퉏z	 ���F�w:L��7��|� s7a��gg� ���H=��,Q�ƫ`[.I�� O�[�@i$���4wC뮈=.�E�X n|��H��[$y�D�W0�Y�xt�SvWn�MU��A��=�5�Y�p����'��˟6�z�༵,����[�(YW��*�%�Kdz$	��Q�(��4bI�.�h]s ��ժ�~e�+kk$A���J$���q"Igص����:�� _��	��;g�x���Y��7�|s2���f�2�f���^�g���;���� ����s�	g;���w$&w1!�j��A��}W۠�m�D Đo{\A>=]5�7M5.�w^)GQt��,�Tb�)d�'<6uԧ�
�{9�%U<�o�ۺ�����:y���Yb��q>{���ϳ|��k�p2������c�T&��k� ���Ř3��'UHH'���A�z#j�'Ca'���̽(��ܞ��G]��Üw���e&|(�S��_}z�>g	]cWBl!e���fx�	2�fݛIr�Sf�4W+�߿�d*�mw����?~�ʝ�ĝ�9|�I%�v��y8���[�5b�^�	��x�;E���̉=p ��3�e��B���Đ�ܘ�A�� �H3�V!ݷ*��*�NL�"�覚7Qq�s�H8�/SuGF8'�r F�HSщEEئv,��0{�05�t��\6�rg�	�>��#3f �q��[��B!+�}��,�1������6&�}�>���z��Y���h̶Mל?�4�q�P'�o�<#<Q!����O�G�ky?8\n��.gi0ԙ�*�����1R=��r������jY��`��I�_)���t�3�n�~����ݷߟaO2f�1��#+Η�u�}�＼|�t8�8��!�C���6�^U6�����[k���4ʱ+0&ٷP��%���v��m��Q�����I�L���(���J��1L���@�b�Ȣv�@�GL\��X�S�u�乧b�5�b��5�6���:P&��Zc�9o��/]��D�J/�[-�6i��1��Ͳ�X�A�;�5ҫ�z䲦�.���U�V�K��&��������`�̚����y,sD���Y�"��2�!�sq�T�����R�G8�f�f��&K�	Ê�߀7 G���ڈč]��	�&���7
:�	$��@ZIZ��@��7~<fv�SOkkR!��%)��q�I��x>$�������=/�uN�(WVNw3�4
���{��k��=�5���_�+s���ͨ��D�u�B�B����gtSD�������	���i@|	$x�4����u&V�4�tFl�^��.��xWnǧ҃�e�v.�3�fy�'na�/!{��v�	M�E�=Y����J	'��#ś{Wj<�5���h~-��ut4�.�ʩ sl*�-���(�Wh���+��I�1c�\�.������n��^�A��x&�:���C��eY��ܪ�ǋ}V�
#�erf,���q}�J�:�w}舳�����m�����g�cȷD:Ժ�@~������^�l5�ŗo�V�F��=�p���*�E������yy// ���x;q��!}�=C	���LU��ƴ���ޅ��l0v%N�̃���1���A �Y�yri^!��ޏO6R��D{č��BtcX,8A�˃>=5�$8TIj�Q�� -�؂H��*�l;ɚ�c��TF=a�ˢ��&���*�A5�O��$u�l��W�}x� �H꼈=�=oQ����a�!^oׇӘ���&�4*��5bѶT�:m�$���������v���ϋ�K��vw�*��y��#⳱��WS<x��uO��΢֐}ٙ]��n]���'�� uwZ�W���٥ϬA������������hr�}Փ(u`uGX�f%�pD��\ze�A=��gn����NS��������A��忟��E�?zZ���3�;.*�9o�m\{=���Z�6�m�cԦ�H���C42�̐>�F{��^^K���觙B�ɽ�gB��
K��^j�B]��pPt�L@5G�^���3:yP�Q%d��'��h ��'<�ku��֍��ټ:�(�:.#��\an-�����QI���]�o���M�z ��ǄNOt=���7L�~>{�*���7[g��J�N���@�p�lڤ]���PY�e��phwI3:I�w{.z �@�){�~$��~�%z2���_scǵ IYr���Ֆ�rY݋��Rf�T$�����}9p���Aoz"	���B�~�b�9��	P��Hg7��9g�;��O~��ŕ��(�8�[��!b�� �^��#˩@$hk�331p���vӘ��Hm#�AK���FS]C |{����:'��S�p�516������O�e:�>�.N�?#7��_n6ċFiS<��7+
�[h2��u5�ᶙ۽������Ogs$Hϰ�\�Gc�srf|q��&t��s�x����L�ua��G��{}vxK�u�a[���<R�P$�_D�����T����y�(����g����PWF4̺���F!3-���k���y�>�/�pE���J�p� �S�y g����O5�G�sv�6Ĺ��v�F�͇�g9��$G�9l�3'd��OG@�8c$el\S?]z0|m7dY�HW��;�;�!j�����n�a���vK;�vx�|j�"	�u�Ayn(��>E�sFh���X�I<�� �ݖ��&,�DA�f�dM<�-�6�$�k�dI9�$��zb���fM�o�׬�A"�:q�$��9tD�Q�B ����p���/%���b �7sрK�2�b	�%���/����4�)�*A���� ��& :9�<+��8�.̱E�MM����l��I�q���M�O�lN�X;G�����o����g��~v�ׯ^�d�窄�k5am�l콱ty�D���j)�֫tјk
�b�8�f+KW��0l�ͭ6$qfö��`új���5�Vˡ�ٺ��%�Yr�Ά���Ị,�!-��0�(��1�)(��8L@�1F��)�PU4m�эsp�U�X�m�)�t�ԃ��cf�b9��g\8շsN���KB�YM�w������یh�F4ԕ�\��C9��arZ0�r.,��*�ڍj��׻�����eIA�ܝ�-�0�����H��d�fqaQ@�\��[�_nDZA�u�a(;8A�ȓ�Y�� �2��c�o��K�Q�6,x��$��S�	�7u�_�u����&��8��fN�7��E��Z�����~������7�͜d�k{"<	$����� �.K��wy�g��=�y���(���9� �������Ďm��	��c�Q!���"���7� �E�m��b��ć�{/ǖ5B���q�Q���ETG��@D�d���7������<��,��]�l::n��K�Ta����It#A�(nՁ^�n��J@����L1d��g.��5� �e@�A-��3�F�9�wL�c����;"u�')grfAȖ���nR��m��9N��g#�=�Ɨ����P��s�(=��qK
�ˌS�h��Bey�gDr{؍X&�j|�pt�Nh!�ľ=3336��{󞂀%�U����`�Dyuvj��l���v�Fu�8(;8A����D�=�P�n��sW(���D�ͨ��F�=q��gg)�;$�L�WD+��t�Q���&|���|I�$��D�:���㓥Я|H4�� �v�,��vvN�#'Z3�� �m�����%����"��y<H'�^��H���aچ	�f�D�\��;S��L�GA����j2���3k�nՁ��/,��B\�:L�;�>0�ל�3G���g�������X"�-��#�{^� 3�~�dPb᜺�]q ���w2�D՞�z�&�����H�ށ՚o�P�]nRt�vw&d�l�c��R��z��H<���*tJtCb�qtU��pz��ƣr��b���S���䤰<�ddᱮr��!f�����<EM\Is��&�G�������y�<H$f[�����m�ڙ�A��H2Edo3)�ڋ[/�53�\� @$���ҳ���G3ur�lʎ��g�y����ٓ�Mު��5�O]�Bɟ��`�Gݝ� ���s�1�|�h��=�=�X>�]w6�.6!�+���z���c6,ȖXh��K�$�v!��(��|��,`��m�l{�͗�r�'3���uuL�������9��$��d: �`��;`��ؙ�Jl� �^yoGjmh�A$�N�<ψ�y.��q�#�l^=ydw�z9�A�r�z�=]� ����⎩����[��7�Hٯ0��s��S���grb�_��͹b��%��.����V�$�ꪏ),o>q��S��gq�w����U[��u%�R���8��g`������3'ƻ��eOx��r�ʌ��|+U�ؑb��8�B�m��翿�f�̱��NEdAusT+���/!��-N�DT���O��TG�{w�̃x�5�W�s�J�e�f�`6�n�ͲEmJ��X)z[F��MD�B���窀��1��L坊t[��sy/����s��
�Y�����<yy^��oB~�
C,���{��m�|ru=�����O�%9�	'���`$�;�v�>˃=�9 �.,t��;��Ou��z����╡w���]�|I���G����8��Ġ�9u1�Nn+�S��<A���$�b F��Dmo8��<0t˦-{,�������Lf:)��vg�l6߂>$���۬s]�l�$#{� �c�|�`	�� �"��A!�H�4u<b5U+&Z�2�����{p�`�q\�r��#}wV{���>�l�e��9�ӷ��$���������R���O"V�g#~x�%�����6v�n����ױyP�f�/g3��c�sKg�&�e�`�x(�!�k�ݻ�]IfW�)s��}�)�wE8�s���7�C��g�_��)�H^���o���L�yQa�xb͵�d|�xכ|�E2��׆^�b]�i����)�mMiuy���S�d���_�dʆ7�`Y'w����o�����8����iG.����$<9�z�8�{��nf$o)hۡxN���������hvk��>ر�#�l�sS�������N|c���ܐ]��C�k�����rYا�yZ�h<�lN�Sw� ��WWW�qg�l�;��}}�|�>8��h�|�eX#	C&�^d˙��n�!*�2�^t���L��Otv���n�M����u�|����ӯ��#�2�w�^,5=���1O#�&\�Z���´&���я�F��3ާ����x����&�3_�p����s�_U�{��0Z��"Y�kYN�{1��d�Z�̀ڨA���~�~�=���@'��3_n�����b�s��Ӗt`���o��f�}�ۃ}Ό��K=���|���L.YQ�E��?�Of����
�!�:|����=�}�^*�a��]�^3�D�q�%&I^_a��^L���~Eb�6wv�j6^+&�gg��MaT�kN~Po�|�,���{�+���A&�������n20��{ئ+�`�$���~/5S�X��JAp�@�������aj�ߑ��-��U:�e3vۣ��m�ٔvVp�a���������]�v����۞O��m�X�+k�::[-����=n㐓:~���؞�v������]�v����ہ�L�I���m�kI`v�l6��q�mB@t&��nݾ��;}x}v�۷���>�s�khEDln9��	֖'D��v��`fg��ݻ|}{|v����۷o�������H�V�a9��6��:�+#��+�0��v$!�!6Ħ֝m�)#�[m�܈;�������疅m���Z�i��n3qȓlB-���� ��������'m��M��Rkem�9��_7om>4�Ũ�����5�M� �{x��q�ծt��Ӕ�9�.G:C5��
HD�O�lK�7FdN��mk�sbm�蜊}��s���vΏ�w��^�{v3�$+����}�}~������|i��q�J+��WX��%��,����k2�J���JjL١vLc.��q��6��%�\[RkZ�F1��:���T�8�%*��ca�RT�Z:h�jKn�b�aa���І�1�+Īmk ���B7XG9��3�_'��3mWYxΙGms�z�e�1�(��1l�=i�J2��sf���FK �^5��6��� ��#Z�J8��Hѷ��ܻ�����b���K�])�uo!�x��nDX����-�핊�Y�Xk2챸�\[���LU8Qri�:%vz��88Ҹb��n,�I[�a^��7Kp��n�ZC8E3��ֈM���:'9�hu�l�
��ئ����+z�m���PҸ�Ar�xR�X�#�V�K+��if��hZ�R�:[]h��s�2�C`!ՕJ�M$m�%у����-p���']0�KY��v�٘P�Ȋ6��ta��!�"� [Zȱn��#`�\�,��B)<|M
�MkmgM[1���Tn�Y���b�ަ��eed��^��j�a��T�����\�q���b6����,\��6]��HL��:˥b�*�#��ֆ��hi,T�h���ɳ�jPI�����e��*:
�&5�dÌ�*k���#�� ��Km�13 ��#]/�0���X91��i���b�0� ��Q�7�tWM�C:�1HWѥv�[Q�-�yn�16�!
��;�΂��f�16X�1{q5��[�)5�)����o,i��*�]T�˴��!�B�iGGRVkbթi5���p),.K6�+F]e�����hQ�F��i`KM�qLY�qG!+rb�JLh�Uq2���W3x�lOR٢
�6�#����\\�@a�k0�m�������L6d4eQ�(�X+xf����`�wXµ�mg�x�㛍�)v �З6$�CB��4�y���^�R�kȘ�]454R�h��ćqĚ%B y�aR��S%+���ڻ�����qN�����r�R�V��pk�kn�6U�,��Di�C�]��f�lsKy#[�@]Yz����aHn#�J�F�Ydȵ�X�U�ih��s
��Dۗ&�a�0r1�2ݦ抻R@�Xb���0�+��v�VU�3\�sE��[æ���CgF9�+�VXMve\�����αu���A�߾�=���کM�5���3KbmF�E+���sJl;3o�>0����#y�� ���@��=Y�� �7mP� ��胞[��y[�|��;}0 �mF�+��-�9gd���UQ�$�j�3⦎��IG��)��k��%E`����]�-�xP`�ٝ����֋DEy�˷�hO��'��B��d�\��ɹ8��`�*�z q:Kc��f�bA|��ۺ·|=���G���>�6� H=}46��f���$zpN�tȰwI���P�ˈ���œ2������D<?BG���B �WTC���@�:�I�ӂ.*���dhn�ֽn�%�nKw!rX�V�4W+<���>��tY���3�bB]��[A�	;�� �LyG���s�yj�͘����~"yG�N��o�&k�gtX�8NK��z*��M�
�ϯ�`'��z˹e^u3v-��K(��m��3x��J �ɀ�f$�6h�1:�U9�C�����w���y����333�i�랷�ϣ�dq��>� �F���5O�Z��C^��;��c��E0�-`[��� ��������jY$-��״d��؀L+����;��쓧vB�ԕsUTT�C��$�u�g�xg��~��I��T,���g�j��$;
�˝;1`�ƽTc� (DgkUzZ��zQ�vo��y��O�&�& };�Dwj�j����������ؠ���h�64�x��.���.l�p�Rm�\S�N�,f��0wIù�ٷ���Iv�ٯJ;#��3zkS���m��A&�"o���2fL]���[���%��]�8K��O�&=W��O�y��m��f��y/��gtX��NKȓ�WIv��$�J��&Y]T��~���~^{����E��w�ڊѮ�e�T*?���u��[�O�.x~�ݮx��~�8�=dE�홙�<w�V��I$�lǣ�����GyL`����g@��k |�������M�A��1�^s��>�܊QJ�:�q�e��쓧v��+�O��$��x�ϝ����fA>�����j0Gu���&��d��J_~�ǟ�_�}�������Q�d��t��\�r�Sn��BgEo�~���߾���(3��A�� o1��y/�ݾ�ª"i�I
%�H�� ��j0�:V%���'��� V��ק??t?������ ��ݗ8�^pt�u��z@K�^Q��Y�b��	>�[ O���u�!��~��[�dF�����j/���D7ͫ);�Ν�9/A�ڶ�i׸M=��w]� D}[yy"
����f��ɯ;��d�N�n�F�[[�<��m��w����D���2(�r:��ܾW���+7�:��x埶y�\�<�O�|��33��|�w7v#�r���JЦ��$�g:c�;5m�������[��`���B�j�h����~��dc�c1$[x�(�H Pu��u�
Tq��,���ἵ�5k`�ϮZ������퐻c��b!ǘ^��8�G�WK�z��ĸzB��S�F˺~��Z-R���\ ��d��ۆ���Z�m˽��D	ă��d�v�b�q��?n<<Vq�}A�V�E��N���;b�A�ۈ�oҶѱmϔa���t� �	����o�^�
A �x'�ڀ��'9V g��` �)�%�s�Go=؞�3�b�g�y��p_���?�,6��II�i��x�sQ���k.;�d���A&n� {���|���0^�1�H3Q�>�7�������2n��8>��b��J�n]6�Cr�o�4Y���{3$DM�#%��݊d}>>>>>>,���q.Dr���.Z�*�7�r�(m*b\�"6��r���U�k��шё�k-*�1���.�Ye�-�v4��f`��6�9h�ن,d��������Bk
!Iv�ar�&���ql�ZDP��wl�[l��´�b��FkbTήt�FR��2�v�2g#��cj�&�u���k�*����22�x�!��Z���<��x�pJ֌F�VQL[�JF	MѸ�\݈���� �>�/�SFw!-�����%��f��$��j0w���w�3Tm�� ��r��F9���"��Do4�n��k����{$�|	9�Q$���oF�ܫ�*9��W�qZ���\ �ʪ���A ��Tx;	�G+U9K5�C��l�$��^K��� N��Z̓'r�;��ӷqʸX�z�� n��'�M�Y�$�d=����Jق0�踌�l["�Y��8'� �Kd"H7����h-^�΀ �b�<ϱ �:�= �N��AT����YAL9��]-p�f:ƤZ�l��F7f�Mɚ�MY�<��!�0r�՜��'.圗���� ���k�|�̈$?ls��PF;V�1Jq��/�EFDx�Ucـl?JV��G���	���A�c��-\*��Bq嘻�~s���}��o7�z�5���/F$��w>���ob�;!�����_}�w��@��O[�g���!~������(����
�u^�3335wך��>'՜�`H��x�z�<��UϺ��^wd�����i����q�|H9��_y�wmf '��H2�؈�yKB�N�.쐙寯~S{�p�ŝ��Jn�Iv��@���{��ȟ]֬�Dvҁq�c�|z}��1	��1ْgb�����M�H|qd�k���ͽ�Թ�`�t�q��+���Ot���<6�[�TS���K�hwr�^E2�R���W �y!�`4ee،eX�QuW���.s��`��fp��Ȗ��$��׏A�V�D��Qنq�86?�С��$�wD����d�ó���軟J9ҞV`��`�Ыgq��� |;��b	"�� �nWm�\��oƬE�\�΁P&���A]/ yăՎ:%��m	1�Q*���e���?L�݊���!�/G�V��-�М$���1�� cf;R�*0K��u96��|yfff}~|��( U�@$���q>_���W��"�鄃��y]4�g4��L�#���㼐�$O��Dx�6��������o ��<O�ͱ<�,.�K���d/{�{u�ۙ��͊Y��{!��]2I'��x��{#��z��k�L8N����~%sDe��@��ښ�����ݫ��n���^����j��p�Ǻ�� M�L9�[�f<���v�h��=�m� o �� O�{=�t32`���=�}�Oε�:����A$�dߦI5w�d�)3]#,r�z��4D\��6�U�Ӧ.�9/�@�V< 	5\� �>��GE��&Fz]U�����Dz�$;��ǵ 0GR�%˸g`T��t �F5l���0�Ј'�]�&��э� �E��N&�S�y��l藙�d*�S�+F͕2�Q�@�WĄwcO��]Y����|�W���g�u�����g6i'�{�tRy<q�DQ��B�s�h�8�������G��{"b%�e�N��"��$�i0	���q�2Z���=�����ĂFֽ�<�����e2j�~�Y�#`������0�ҍ�92��[4e&f���w�un�..�K�Γ̔��U�$�ǸA�goL�|кf��\�c��b/�'3S$��;�v5��ۈ�1��%�K��l<A;���A>�� �bA�'�#x?�������L��`�ݜ"&ND�@{�� �L����dGVlA>�ײ�{o�	Y�i�:b�Ӓ��趢Բ�cu�0{�C�6B%��^f̒I��ꮑA�X�����v��2��.]8v�D�tNt�i�p�
އw�w������'��� �A�舻�ŉ|�!'���HN)��Ibς:�;�;�B�?f��ڎO1ڙS?��C�&�.��cVF�uoNW�v3-�^ym?w�8�8�/��|�+�mC0�h+�u��+Q��j\e����:cv��`�L�0��!�q���,-�ii����8��c��e��t���4҆r7���10�nY�I`��0�v��L�d����Kns��h[�:[��"!!C��mB�(�J�n6 cK*���&��.�����&�6��٫4����qX6R6ų.,�}?}yOSpڕ�.����V#a)ÐY�����f�jl˚z�����̝fE���k��<�"n��g��b}>Q����\�"��\���5��*�"<w���wpY2r�H�i��AC.i�؄Z;3z�`"=y���>�$7D@ ��ގ�"��ζf)�Ӹwc�4�F�$ە�q�&��78���#A>�܈$6�b3ӱ��wg
$�l�����;O�̽~$J �F�T�.��q|�)h^�=0$w�-�<[�w8�Pe�߿�������3���r"�h~�]<H;�1�����G�"������g����h��5�06�h�#V����4�f3%�M
������=��G~��#X�n�Tc�|d�m��@�H�wDY�b޵kp�6,g���%J�-�/N�3S2t�wHUx�kT!�P���g^5T<��y3��,�o{k��ڤ���s)M)"��?`�O��̕1q+Z"%�DE��=�z�||||@>;����et���梼`��HL���%;'��Ol�"G4�	
@n�g��>����Q	8�����d��r	$��ǠH�� �ػ��i��h_����`c:g��R�?DQ>$O�z0ψ�)��q&�v�l��H7]p �r8���မ7�w"��x勊�~�%;�L��3E�<��z W���hWv����*s�����=4l�ms��(�Z�ٮ�h�+�V�l�\Ы�w�� R|>m~5���?��>y��ףǵ�����v���LS�q��o�;`7����g1�|�!r�K�N��d&FWW8�$u���Z�s���r阞�	��z0	'v� tL'���4l>�w����2t�wN*A]�0�dO�˖����f�v�W3��z��1�ʋ�hk����g;^�
>�:���Vl~�����*��������q��W��>wȰ���7���fS����S�`�����!�o8a�=}3��T�����9�=�#"���G�T�+������Se�y��G,N?! ��h���G��/��-��`�E��6���]�u>˝��l��O��3[:��㫽��-�4}=�Lo��n=��f��-�� S��?�Y�^y��ї��yt�a���q^�)�z���<�0A�)�'���я�{�����;�{r�yg��A�r7�{��^q��p��)���&�����w���U��_/�����kq��`꽯�!�]+]yӏ������eA$��9�W�<DAyW��p�۳����4���x�����^;徚߻�4/v�_�Z�)��Q�H�#��e��t۱�|���y��}R����pj�w�=�qy���W���wz�i��M!O3c��<G�}�@=�}���"9c~/eo��{��y���Z=WE�wIG�MW���'sAyfw$7��ɂ��})����]U�ro����]Nn�{���'N���8�p�٨�ݣ}3�ɏcx�;(W?y��*�~�.˗_�~X���ﳆ��R�!��_���C��� �/����=���Z >��x����/����Y���h����P���v����|"6��=ݟI7��|}�{-8$��o�@,�șۥ-�Ba�3&AN-4�V�=�;|v������۷n�|"�i�����kfP����)�#8�ӈ�o]�v��������nݾ>w�}�ǵ���~�dBs���$��k�݃���-kD�"rص�TUDm��������ׇ�nݻ||~������6�(�$&Z.��gh��Iq�Ŷ��~w���z��������nݻ|||s���2�%�|^_IH��ۂ�jʹ�ӠI�iIÓ19"�&ڔ;l�${iޫg�D�#���;�e�I.9.H��},U�IB:r�$��[��8����ܖiC�Q�[l�A�m�[��l٬�^���w	�k~��QG:�նqgm1����~m����q%u!I���$��vJǶ	k��N$����H�)[h�ehY/�0L��c�矍]��ߍ�����%���Z��,ҙ/�m��z��6�h�'��ZH�D*�bقk�|�_�\�1�Q����h@�;I�H�7�L�ݝ��;����`�eG���b/Ugs���p�'ϯ|�g��S���|��OY�￶4�gͺ�H�.�]�.�d1`���M)�J�Z�lʪ��z'�~� �&s5��A\�B$���A �F�L@,�Gyi���|)����Hՙ�&-󭖺t�Ӡ��:kv�'�(�;��UO(u +��u��GW<�*;"�����X�'%ܸM3=ޯ3+:b�&����f&���G�#o2 �v�^<7�*�i�V6����q��������x ����p+Ɓ"���6Iɼ%4���;��+*�R{���ő����ľP�5��lfbݛ��v#!�m��
t�`E�M]2.%J��n�A�������|||Gx����:X�9t�7u_�/�Tn�\f��t��I=�. ���RY�iv��L:r�	w#���L[!Hi�ZLZ��ۨ�jX�,i�m|����� õ��wgd�]w�n���9YPO��n�݆��B!�����^��������
}i��!��4�/�qw��Cc��].ۘ��@�n�|�QT�{.�#Gm~�5�2�N��t<�d���>K�u�W��$�;����`��2������H��O��`�J�lX9)Ä�OLs�c�g�G6n+���[ϟ��U�A'���K�U�:UU�
~ȯJ�kvN�Y0wu2h��yω�*�w��{V?��5�Q �a��K6�#�Fl]DAp�2KI�S-h]p�6Z�$EYO�;A������8$���D��"�	�2IA��FJeM6I`��v�F��մ�q�f)p���������a�vw��.�pmL���v|�m)M����kVZ��:��@Õ�s��4f]��V�h�1��l�ٮ��aoG��M@04Z\,���ih���Ā:�՘u�,�u--n/9�V�	ԕ��:U���54.U@�fh�ca�1Y�l閑�Kheٌ�F-cY��]�Ll��	Yhkr˳kT6�,��2Q�\��������������#�z�!6)�]I�(��Jh�\��L�X�ci~�����q�0�C���+>/�o�l�S$n�D��U�ҏX�� M�f��Hn�m��9fr�ʭ��N���}����0۰	2�頂7��}(�u��c"Ǯf�2�f2'2\�NĄ��L����rEngD��~�n�y���w�	�+6�$�_@��܂���t�Ӡ��(t>w��ɉ\,��Ѿ�(��9���I;]9Q�-��p x�[A6ysJp�4��tA$��t�O�c�D�H�s�@t�8����:�:?!��w������e�H4�xVRE%l�n�q�W53,�]
�����uRL�7���Y3�0wu�5��!|�� �t�x��̹��<�O�A�� �1�J8�C�E�;����z��Ǧ����|��'Gno�ZNzj7rD.�M��>�]��B{�R��]N���9�C��n��a�bF�Mdz�||||||h�v9-�]�A�o�� ���/�/]��U��4�ݜ�9tbdv�A�6Lz����ouKF+�㗺�o/)����{%˲t	I�4�9�]�����l��y|B�ʁ���;�躳�˄�{1HUT�:r��y0�����4��WfT��Ξ�-.8�HG��@�Gm�����ś]W ��� �IѸb ]�J�:��\�dгMA��l�]���4��������L�89�``�0O4�En�^#yO) ��|�%��\�ی���_}���읜�`��g��~� �؁�o��'WD9�A#�j����e�9���+�pv&���9`��<ޡ+� ��Mr��A�v�;V��u$d2K�Jv���<zF����i���O��<=7;���ԁ�E})�{/��j�S+���gw��";(��/m�"x�������_�ڶ��G�� 	�C`��!ȶ�$�%f�m��%9��;���X��D^\A$z9�ǉ�"�t����n�3$Gn��U��&���'@������j�ā��p���VQ�ņ����@8zu��7��j��O?NN3�=���|��\�b�ڱ�p!�+��փ��k41*��k�4��34`�ȶCd6?��f���G�7���Ͱ/����AIC��<�O� ��~1�l4�V9)���N���$
���j�2;q�{|�W/�y#�����l���$E�>����~�d��wQ'��"	 �v8�]�S��S��fׁ$��~0A���D rxBV��v��H1��f�}3���F?��O]C� �y��A'o�W��X̵�$]�m��]͚�y���|X���[9��y�8L�� ���gk��s��t���������i���0��
��ᒣ��d#7�� ����?BVE�����%L+ݝ���ǓH.A�0�SI�QDd�#~��w���������SI�u�[1�L��ܲB�C5��n\F�F�d����@-��{+�L�� !��"hP���w���d1WWI��@u��ky�E2�I����@f��ٜQ֊eeT;SIi�N�61��.���~\�����8�A;TB�|�#�?=��_L|/�bW��.���D�#���In+aVd\&���O����N�\L�Q3��~ݓF����0rS��z�:=2��H|@%C����/\D��Y}I"|�:�@_S$��vS ��j��غ���@���<I ]�DG7��tp���/!��"*,RZ�r��vS%�j=�q͑f�<kH�Քw�3�ޕ�ْ�<OG=�=��r#8i"j���d]婆LZ�����ǣխ�vTO:���S��U.��~÷U��V�*��:�0����AZιї<�q�u�%Y��$�q��<�[7��-[��[*7a
U�ki�B��r ��ΰV�Q6�g;h�8YIa�2��$�� ͌�Fau���
�GV8��f+(A��Ƃ��b��32�*A��e�e����VhRl�v�*t�r$qHKe9�h7i01�d�5�J�cn-��,��E�ɳ��NTr�8�[KF����\묙ۈ�Enu��E��������p2�+r�tMe�37X-�n���>���Y��;:d`�wO��,���	�n7�
��^>���G�]C{P'�"p��r��AA;���*�k!6�jG=;��"|�5�9O���[_��o���b���^���2rrA3�wd�A(���@����z�Ēz��<@���&��9X^p�;Ba��"�+���&纉�E�l  ��!����@'�]�n(�="l[:�
��v�[kvrY�;4
����O���m�v�ə�|!ir睽��D���"-��� ������G�`ڠ`cs�E1)��Dȳ��m�a1���]�w\��묨��|����K�^���>}������D�����k78�,l�^+`@&c���;�d��3:e9��wI����>�.]'��}�4�ӷ8�nṱ=��_$vj�Np�GQ�����>���޹�7t�{W�ݹ��Iݳ}���3W��N���u&��
��*��$>>> ��GO���X�`�B�z �n����n��6	��.���x@��Y�I��An� �sg����q�f�� �o��[��r��<��V��s����-T�`�����H���p�/[=�ǀ=��`"�"&̢9ՄI
ި�K�E鍛�3$G7lW��Dǯ64�$�^�|F�LB��J����@�訂ny���ċ8�M�ŷ"�愖:1q��ʰ\8|x����5ε�e�~~�����^<u�+��O�:�<l{�9�կ]��[�!V;�^I&�2q2]�`A;Y����4F�{9�<� ���^�H�x��r��}�������V�d�33�S Ou�=y=�;��1[o��9�縛�N�U	?L)u7�/{N��.�Y���fe-d˾���mG|.�Wˤ�.�ĥW(eF9є�5�"
f�o�������綒�-㕗��OWJ���;���� �o���zz쫋���u�``��瀼�}/ ��-����N��L�̵ۃ�,���g��HA�����⇪n����T����D��q�ͧ��=�9�ר]�ȸno �ݐ�GhfƯ<ln�V���ŲZ�K����c���_P�YVrC$&̺���o�䀤E����=/���-S2���d�|z�b�ɴ�Æw�->[R���Cs�."�d���@$̗�䗒�gTq�&�c�����6	�{�����3U���l�#�|WP��<��n ����	t��4�9��L�ft�	�Ӭ�j����_ɥ���}��d�g{ 0�M�ԋr��Qum�ꓰ�"��>]������qW�ݲ��A�d�u�2j(�2�K8pW�ح17V��٠�<|||���IǨ� ��=�Ν�%�W����^2�ポS5ɢ�tKN(" s�����z"Q��^�*�r���e.�LS2,���6h]Ƈ)�ڵM).X�[���	�$��oTх%��y0?	.���YKy ��=�>o [{b<g���޺[�x�^.����lUA���ش�u�A0�����Crࠌ}�n˺�]Ti�,B�؏o����t�q��k��3�3�p��٥z|���$Ю�dμ����)I^���$5/f>$n�C�X���gL��g:��L�^{�׆���O�WdA=�W�����=m���|5!o�<[�sPH��ɜ�����$z��B��o���*����q e�@A����/�������c	9�����P�1l[^%g{��U�D��S�h^�˜7ޡb~A�i�f���^u���ҹW���F��D��٬���si�Ƹ�L��:�v[}u��אA(�7���6�;Ưm��Ѐ*3���Ｗ��:u&��}ͬ�.x�ML�"��^�}��)��̤��ӦqFh�m�~�X�W������q��-�hP��&���휗�{L��C���Y}�ym^ђ�ObJ4���h��8^9�]Ra�{�3oo�䏾K���n5�uY=l����ܺ���^;���:�zΜރ{����B�_&��n��>���{Q��OA�䑜��~�^��2��߅��[締^ ��|�_{czM�;9	��t�dupe�v�f�
�)N���J��c��.�R/f�4���7u��k/&/z�ب`��;�H�y�}���۹�H���jDo� �D`7C�b��"�I�wQ�0�}���FzuD`ǩ"��0�곮�*!�z�y���zgfN�T�(���,
����e]��w��#b��x^+������q�7��Z���v7��:��"��(���*_T�J���{�;̚�n���3_�^[�r���/Z����i��Ւ�`O߽�q�N��(>���b�=��׋��8a3�|3��e[�9�@��`��s;HUfA�4��d��<3�Y�za���ݣuRoZ��d��0�o[��|�s/p#eٳz'WhS���U��>� %y�knĶ���!mb�+Zfl�6���&�+*�+=z~��_�Ƿ�o��O�ݽ���{�D�Lr��1ʊKܗ�r�\��[��lݹ�9)pG$"�EPA��Wv��������������߾���^��}��fƶ�H��J/bÑ�r!̈�,�m�Y�s��YI@�0��2s���n�__���}v����뇉ʋ,�s���& ��v�jf�JFg�E�H�m:(�ٵ�˟}�޻v��������n���ޜ�(��6D�D��s�v~<��P�k&Չf�@��u��Ŷ��2�"�۶��K-�qM�e���	'9�ɵ�6�N��x��I���Z/��ڲ�����2�S���ma�$pr�$�m��s�(	��p[v�����m��nHe�#��$q{���GH��&�Z3C��k	Kβ�����D�j�m��p�m�6�r~��ysv����
mZ#nΑ8Dr�$�k���±%��9��y��h��������&�`]��0135�Ԗ��ǞOC{,AC�ɵefvC`+�%\�L$"���
hG)�FdD6�fR� Qb�!s)y�Z�d
�`mt.�-�� n�ͣ��8+�A�D�ܓ	�:�iH��������efJbX�;%��pBn����2�uee�!���j2��i5�A
�����0�f�:�ЖZc�"�K�\�.t�\�2��GP�W��R݃8�ڴ�0UY�&l�]
���E"�bZ!�K�3t��P��vq!6Q�0+)��嘍��ZV��6�b�3���� �3L��rvK,.�I�n�s5R���a1���a5������hF�5	�KṾ���$Q���K��Q������"��ы��j��sz�e"3eZ�m%
�GXԸĸ.��ԡ��55�\$Mc5�R)YY��X"M�B�����
�� ��ui������`6q*Lՙ��ZG�aY��s)*�ml�r�Q#�nL����t�-���[��PITau��Cl��u�Ќ��D�iV3.h�����K�élI���Km����(��0�5(�uC�]��Tܚ��4e������F�*b��؅42:\��F��mqH��B0T�]�h� ��5�p�X@�l�t 	c4�85����t�#D�,�ݡ��M��(l�h&5m�+��]33���֚�h���rט�����Z�Y�R��]�:�\Re����P�ԭ����@ơq��;5iW\� �0a��Z���F)q�Ō�&E1�t�Ib[qsv	�H���V�6$�&$MH�݋v˦�`�s	f0�V)2�!�º�dde���1U���5!tfk��d�; �&�԰�+	� �t��+�m�r�u]�&�5�Mh�X⼦�ʌ���KBu�b�h���	x�d=y�u<����+b�l7�!Rr$�8m6�Cq��/�,��k���e�T
�z�|qćqϑ������JK������ґ������3qc���J���̄��+w�0V�gJ�e7ѦR��fT��M�l�D��Z�e0C��e��ƣ��t)c�z�.0@hm���m�G%�l��8�C���`������k���X:�2k�AɢM`j[0F�mr"���Q��jя1���͗ �֋�%ԅ2Kr]�,���>0-�<d�b�-�Xd�0���f����%�j]��U-�g/������acX��������D1$�v8�C�<��nuDx�����h��md�Jo���a况��	�qy�"	���=Q��C|c�ݱ>>�� �
w�gdK,�XH�u�,\3b�=[��������8�.vW�u��
�3�A ��@�m�{N���fr�Љ�+������jp��2j�A$�H��ͼ&�1�o:5sQ �t%����vt�2zuQ g� ;qp���]6���e�D��H����F��ٞ�?%>?-%��8v@&,t�lv��,��6%�FaH�lY���q)�f�BE��L�w��"�_�D@>'��m�a���Trז�l�'<��xG��u�wfr�A���2k-��y�-��笖I��V�s|g)���܎]��� �����\���i�!�f@�8�v��W��x�ѝ�]������o8�r}2��=w��	��}��N�������Z�T����]��F��h'�t��%�r}ȩ��@�=]㳚B�G�Ezȅ��h$ϝuqʸq�L(�;⁭�q �]6��Ho]�%.��j�W_L�����_�ިI^Hc�N��3��$-��y�E�O>�c������}�S��gN��4ϊ�Q�*+����q�=��L\9Yx�y��$�W:�'���y� �3���������9��L�*!�sr)�k��ra��e����:u��
CYs��wL�O�* �ؔ�w8L�b1�ԛ]��|���䇮8n��,��(B�� �y>�n�<d���S��Cx�F���v�R'/�t	����9�l�1 t��wfr�A���2w.��>=��$�V�TӜC��+����3!���'�g�
i�^�I�i�39�������q&n�:��Ul����.ӯaޏ�����[��8�imC@��@n�D7m�̠��� sM�\n��MF9� �g�s�I3y�$��e�X71� ����ޛ�X9p�]�U��]3 �eVGLUT�cߦ���� �}]�Iy�����1�n+i�1��G�Y�ٜ&34,NѮU��lW\�Z���(���O8���W{�Ko���67+39vo}�Q�����y$��\�D-�8�u�?/��&�h �}y��L������ ��q"Ny=�#�$D�S�	&�F-� �����@�B�5�q�	��z�,�gd�U
ۈ�M��|�>o$c���jP/��^`�����I�~�G�ٜ�S�ၑ��dȭჼP��b�}�;A�i�^5�64�f��f+������b��.r�R��:��^�R�f)�6�f����M| ��H `ޫ;�@!m�/����7��uι�8߾\y���2�8�#����z<�.���8䓽O�G"�dǛ�M<�w�q8፜����%�]����5�%q���Z���7$طD�˂�b�ٝ�a,�0[���\3b���qf-q<�D��]�\���]ߞ�\��M��ݬ���] �dsǣ+t����4
z
�W@bOn�L푛=Q��y$�/�ѓ!��'ӭ<������⩽�	Wf[Y܆�ؼ�1ӱr�O�2���B� ݺ�Ì�}�`�r�"�uO)�$CPA0r�;%-�ճ�6�7s�|{_�$�i
ƬQ�A=]���*�$j�'�G�ٜ�S��
1�n|�=����k�P���,�5�d�y��{��8Dk���;w�X�[�j�<��$q��A��rF��Gr��q��d�!�2�и�X�L\`l�9��4u���0�
Ɲp���Iio�8��w�'��H9nÜ�k�9���m�,�vV=���a��
���k���'et�����Xu��®j�ءI��a�Ƒ��z�]	t��3X����nf���F��RK�ƉX@5��g���Rjl� ���ِ�qk-�G�����ƆM��Rl��`,0S����v�nmNc,���%���3x��[�b�·hMa�$��I��e��m�h��2�\*�m�eXZ���1t�a�M�h�6�(�R�5�n�ŝ�����A�S��O����&^mJ�	� 
���zB�+��]�i\3bЉ�}U�{���~�����ٛ��Z�Mm�Dx�@#m�G��'[Z��s��tg[������7���Q��H5�� �
��bdG3X��HV3��W�F��B �����3���ܼ
�Z�7@�\��� Ӭ��(�&���H=�y�����L�G+�i�)����& e>���'��"vkn�$�
'��8��H'+� I��=0�C7l,�K�G&,�B�;R���Wk��S�f��e��Gel4���$%���3�Rd�?����$�ǂ�P�%�+eC�4uN�˅R���5�K^����� ���c;�[0~�ȟ���_h<�^K*��{^]����e�N$���D������[J���d3ۈ�w$��0=���>>>>>=kz�x�s� A �w�	�
x���*_�1Tc	yhmɀ�>Oq��&\3b�"@�ف���A�����g4=P(�{fR�7�܈��vߢ���fgv	�ٚW��#��^}�q`��[	�����dkJ�,@��'ջ�W�e����Ý�p{��N����9 �Q�I�`	�� ���y��Y��A��M��<�y����fp�ɨxL-:�FhJ�f���ŷnV���YM/ωK����Hp���ʜ� ��5W+�*�=<C�"'�l\ۉ�Aϱ�;'g];;"�$��O�a��/:��}�$ �S���KĤ��Gt0W���&#h��)�K0#�"Aǻx$����H,�/X'�nF�����wR5ȟ!��Z�oe[��>x|��<$z��}�v�g�����N�w�y��gXn���w=k�k|Έ2�{��3331ǳ*#�'��2�|\�Z��[�ӴRo;�Eش�������{6Ȳ	//W����h�'k��U�WW-��DЪ#4����$��A�;�N��� �������x8�ܿv�z��}=��Ii4�y�\Fx�Z�x�m[%z	lp�&E2Yy.1+����Q��43��&�WT�`5������`���wwL\2w/�<gg��!�k!ϭ"F�DAwn��뉩M`��^��E{�a���ï��9)�%�Ul@$�1�Yޭ��m��q��Vx�	�h�i�&D3m�B�T�1F��OQ/='��;'H�)����r�A'/��$Q9V��2m^8ӓ��Iݑ�FhQn򘱁q"h�fJ�;�+Fo�(�k��w�"�!����S��])�r�*n���������4���9M�ݫ�I�Ou�}�vx��6���h�ߖՁ��]��D�l����9d5-�oL�������x䧯z������.:�sb �nsoR��,�ɲ�A3ב �:ۢ'f3ob�������KQ��ħ� �pG9n5R�[j�2ݬ�.�T�&kU�s���w.`�gv	�ٚ	)���ns��O�!o� ��ۑ��M��i��=M��W{� ��fk��f;��Vv��d��IannvD�y�+In�A��c���"�S�zz�cNa��>�!Vcq`ߛ��r7�&tRD���I븈 �����$�t@�y��Z�I#kz���J�/�:vE2Nd��������v�	 ���� �{�W3k�[*5� �[#��-�zf`G�H�Zn��ObS�Cy������@**�(�H;� O.�l�闹�L�O�7OtX[*}�Y��5���%!���x�e�l9��=u����צ��>��f��M��m�'�����7q���陙��s�U�8��B�iQڒ�s��b��.�F%���#/f��[�W%���=������R7ba���E��8Wckm�A^\[@�;�<����U�jK,s4�����s2D�]��!�aG��(R9�2�����2B4�G�6m*ZJ���Lmc�J� ���5.�tH�����6���A�LV�ŕc�&{��5�'��)�rRy����y��.L�U-E;HH:Й��f=��nq�����-���)^l4fow�Y�o!9�8Hdy5s7�_��P\tnsۛ'��@�a�-ׇ��vl�gv��� �����n�ҽ9�锅gOzg���i�SR��U�}/�=䙷m�س��̃9��J�$�Z��amʌn�^H�o2c�~Q����`�6��rK7�;:*duV�S<7T��a�� � ��Aw�%9E��>�� ��].S�dS$��A�q�>$�v8h�S��V7)v[��R��䁌Ƭ���	$v��x������6h���Q�ɛZ���\h��9t�ׇ:P2�-t�g+�a��\�����U�O��o1�>ɺ�_�{��P�>J�b#�=ݲO6�/�BĻ@�0�ƛPHn9H���V�w�KEl�@a��4����c+.Ȝl�r�ȍ�>o��Ր�����d�h����r�R�O{v����ِf��\��ٙ��qξsU�E_7�>gu�/W>�x���d���u4,����ӥ�;�N���&(*�Mt��#�|��vk�7�9g�b�Q�J�� ���	��D�um�v)��N��
s��%	�4��x��=G�����Y�H�t�3�]HGI�IMР}�O9)7�;�)���؏	=�s�O���:j�|������L�lG�$�����ۧ��e�g�h�^^'���S�O/%�b�;�Tř�.��5���.��Jjm��U�a!��|��+]K�c�ڻ�$��ǂI��D���2���G�|���D�lA<����]��&(��<zzr'gz�ӻ��C	�� �� �b�'l�S���Csbq']��4
�g{$�9��>�39�����'�_;X&�Dd�B@{e��fn��_��F�D곎˝��䝤؃%B��M�L���&��8�X'���/���w^�wN�r��Ycx�w�w�<��('��L��w=���S��aM&"��x�`z��6p0����*	��ϸ�����ۺ�������:u{;e��Ű)�՞_y��`L"����^�}|��+��q��{���}�>�}�Q����	�o����jv�!�l-�=�M8s�[����"
��������=7'����gaE`�<��s�tb=�����	��>�e�A�[�c8׆�(}��������{r����8����8'r�ʗY��-�{^ͣ|�˽�������j��ba���7w5 /��{!O�;:o{}�>ξ�ϗ�מ�޴O{�=հj������}�������4P3�tL�y9��*ۛ�Q
-WƱ�˕�橉q��W�S��{���rv����~� �zh�v�{�ܙ��^���%d�,�$c �$�b�dи��/��Zs�ׅW��Ǥ�Ӗ��L���o��e��S������{N{ƙ�9�x�	�՝�]��ik�^Yؽ�-���.
��4��/�꽲���酑7fV5�V�s*�_1�`U�E��ܜ*���0߶I,��g�����2 J�%�{��m�/Q��K2g%U�idj��)W�2���̲p06�2�d�ܒ\�ZΝf�<�Ok9�ANJ�l�[�;�ߏOo�������v����͆XeY���嶑�rtENL��@���y�[g|V�DWQ�^>>>�}}||v���������熧��0�j��h����(��@�m�bӄ�$�Qv�����������������ۜ�fQ��bd��TDV4����Nq�|ݩ� �y�,;mM�?}��]�w���o��__^_]�����`�5Hq�Ӈ��JAC�nD�BqHW�Iy���Ȅ'9	Ey�:�@�Y!�'��h������R\�	N��������q[l��t��Q�rI8P{b"E#4
+�Ry������8��#��E_�� >���pGB�_���hT�!GN6�#��Ò~�c�9$'D��'"|W߱)$S��P��զ6��LԄ�D�1^����������|�zB�1�!�,�d���ٚGJ~2��[�뉖Fܐzz\A]lG��v��@��7���-� ����ӄ��'r�.�6� ����͇`۩�)�Z��Ot�$���DO�$o7Z��'��hT���R�]3���1f�ZE�,���q�Fd�3��
TD�����s��r�o8g.�Vf@�I��|�^�/��pי����R��G��n��+�)Ӳ)�p�w��2��pMg84�Dd��߉��on[_�I>�
�n-��y��R���6�`$+��N�	d��W;��"k�u�Ng͹�d�dd@ �;[���g]N�ዠX8f�T�]
��s�V��nn`$������Om�]���(�m78)G�}�b�C��^�ޛz!��R	鈊"f�`���ݳnu�t�۝x�F��j���/����C�;�������=ĚǷy=ͬ,�݃;�3\�Z�C�fm�x9����+1shH�n���;�����x��$fyk��r��m��ER̩��M�]��Kbg�U�ík�Ίu��,˶�\�p�8d�\��3s� ��YX��l�Z�'˩YZm����Ɓ ��d8oD��P��v!�9p�Mu==�=s�B�;g+)�k��� ����p������9a1�c�N����}5t�:vE2N�W�)��F���Đ�˲ն�$�c��'�YpI#��'�4A�5��%��Ll�*u�5�?�r��L][�$�鵁����#o�� ��r��n�sԤዄ�M1-�`�K˫�"\�I�_:����!��8 �nD//gtȅ;l�*{�6C6��!q�i9V�ަй|v/��$�Ӧ���qU�u�c��ђ�*��.Y�L�e�6f�fS@�_�������\�����T˓P�ԋ���#�:�15fK+J=n ���43�q�jaH�ݢ+,��;K�L\��X�7^AB&Ѫ�#V�bXJ�a,�خZkU��+*A��m�-!Z�KvZ���6āVɢ�K�@n�Z-�K�;�2�b�˵��l��
P	��9+m�H��uԭ�X.%��b��-fg-��\�ѥb	Z��e�J�`M������'�t���άe��e�͎AD�ڳ;3�R��5�b�X���}���b��;�3p�������	���wJ����Fl8pNy!U�H׶]8L2g2r��	;��\��H/�f� @'�;� ��#Fd�^��a���v!�9p��W\@ߒ+2n�h��
Q���j��9 �ܸ�=�0!��k�N�&I���sL�y[|��drou[3#��	潹��3���7�U�q'U7�7s�䛴�K�BY8������H�\]ɽJ'qŎ}��O�z���A/��-|�2���:p
�����i5�&��K3�2������&ź$1±�F�eH��Ĝ1p�9)�g���"z= �d�x�LQ$��53�.��'n�/�� �u�A�W���wt��X[���|���j���9�lL�'�
��OQt�rz��%dG�XO�E�&�M
s�;ۃ���\��kD�}��(�qǻ�x�Z5��y74�������|z�I$�@��� �n����I[=��q��Clu�9g�K'r��Օ�5A�XC�|�*Ť�vWT���;䏎n�\��k[��웝Eb0w#��'*�	�'8�Q�A�^Jݵ���ݻ
Kvlu���Z��
i��Ѱ�g`��'�I�c�,�dtH5�U�L5�ю#�y���	$]���sk�[ǥ��N�0�od�M��Qb����X�2��l��݉���Y��)u
�a&�/���~��1?�%���� �;��!�$����*��ڙm�����g�Y�<��LZO�pC9)����#yf��T cC�/^a��� �ݗ�^H�+��(�{m�v��fq�\�K�yb�x�dr/v��k�%���%�u;�j�2+�}�b�d\!A�f~�۽O�F=��~;N��~Y?������M��߹�����	�����wy�4|������\DA>Yn]�3�Iܴ�yuu����tޕ�O���D��ǀI>;�(4c��`�:Y�����JA�;�3=�	7�1��8Qjۺc�H�-� q�����yY�]�����"����*v����7AT�p|�;�Eӧr�k\5�шsj�[H]r"�co#��1����34�;<a�$˷�D�oT@5c��s�UI���Dv�A�(�랷t\�N A1@�VFJ�LUE)�N���У�N�<I��G�3ݥ0�;����Qi?���Bd]GDH|��{\����D{cx������=t���V��k�Z����'w)�P�M��2��|F�c�oQ>$���qH'ݭƱ�_��k���]\����yB1��mV)�Lb�qf�Pj�5f������C!{;B�=1.u���p+z���,���Nc��3�17����Hg��,��$�X�F�M��,4��s]<=A�4c>�B ����=�ܣ��Fvij&[Xt]P4X�Y�3��"�m@̮b���b��K�!iu+l4˕���P�?PF��;�^嵊���1�	5��� �FG4d�C�8�>@���� �Ol��3��r��%"^;p:hx���6~����O<[�B[� @�F���-uG��Ρ?����M7�v	�4�!�(�#Ns���yC�t��J�e������m�z�^�ܠ*f�3��M��~{c8�ZH#�.=ў� ��������9�޹�9� ��w�3�ֳ.�.�S@�����c��pl���cU咽ۓ3~D�j�=~q'69�g�Z��6�\\�*�v�����v9��W�aK���E�M �iF���k��r����+{N�_�}毶KY�d �ʪ3�r�~�>s��<����٢S��X����q�t�޾�=߉yձ����3b�t^&�a.3f���	U��6;ζL%�sq.2C9c\&�cÝ�-��f�nФ0��I�[���YvM�����Mj���6��J��EGPH���` �cveWjD6���� �[)��٫�-�T���3j	�uvl��:��5����i2�.�R�kSM��q3��^���翬���~YtQ{B4��`�r�������5�ej��6g��)�nx;��ˤ�Y�zx%���y�c�$���[� �p���b�xާ&pl�Y�K�33�q �M���#=��*`w�˓�A-��&{v��[�����)�:L�8x �o�9<��ǀA.��
4t���pO��R�NA�qd��������N A2Iu�O���V'�}�B��$��ݼI=�=�_wyh���\��E��g%4O��"����Mq��j�ǥa	���ywuW�[�ʵ���EI�,|k�n����b�YF��KL͋i�����M6^$;{2��;���M����%���A�^��61��0*#����y� w�X;3�Iܴ����{۱c�}��$�������b�D�ޛpS�_��m���m㝺S���ط��=�R�B�ȘyS{6bПcU3B'��>> �4��#�G��m�Ezǭ�o[�+%�--~���WoF�L3����Ӆ39��I7�0 I��^�&r/u�TH'�7q�{z^=�ܮ�'f�p�*���ca�>1l��z��I7B�ə$<�Q�T0	n��
�N;.L���]b#�s��ޮ�S�s���]#�	���$���Hs�'Wr�j�nWs/5Z�q.i$J�a�R��d���Ѱ��ll9#���9-�b%���c߇��3�lt_��rSoM��] ��H�ܜ��gZ��ӠU���&�� ���vt�]æx&�+��'��5(#���f<z$=����8 �Nݤ�:���<m�\�0vg.��h�gA�눏$|pտ������['�G�/���ac�<מ�8���ǜ����J����	��#9�b�lܨ>�	�j�&�����z||<���w�I���R�N���Aغp�z��'Z��6Z���&|����!9�?�msߢ5�0��c��f���ك�E�<Ƀ��6x�{|��+5��H-/�0nW�9;�p�Պ����> :�8�63E�q�be�4њ�(�Wkja�T�u3��֚��}(�L�k����� �
��:�<B�5tG�O^cfS^�ތ�JU��麒�tK9)�g��	*E�c���B���_.	$��O��yf�<�X"T��}[R�s�7 �y�vt�]�v�s��m�xω7q|�zmT��>� H�W�9;��'��Kfr�;����ݴ���쿒7���{K�$��ӝ��Y��ݗ�-��{�(����ت�������/o�G.yv���wLѨ+� ��,���!�\�I�D��f���.�Ӹ ;$����(�>�Yn0������Y�';^�x�k�pI1Դ��N��МL�C+��~��<na�'P[<�:�8�J��q.�sR81�� �x�R��k���(ɫ^�-�m;�Ic,���/��b��E�8�N�/o���[*���hgp�{o"	�gp��ӈL��_� �$�oY����� ��FI&xr��A��K���å��ְ[טx��.��@���1��`�	�ymuO�/[=�»c}��Ǡ�F���N�LA�<ֻ:�.�Oz����RڦL������@�	�y��d�s[��OK�m�1}Q�WZ\0vg.���������`;��3�+�9�$�nL@$�?����]f#�(���� A�����p�#~���D09�N��Y���X hd e�Ri�Vi�`I��f�����Y�`U�� ���Ua�!� ��e!��Y�i�DBi	�Ai�Vbdd�	���ha &�T	�i�dU���Abi�Vhi��BE����& ��&�a&E��@�&�ViBT���!&D����f�i����BT�h`HR`&�V��dHR��`e	
dRV�� f�� ebD�� `�� D�� `H�� na�� D�� a�� a@�dH�� aXaC�� �HHAHHHHHHEHN1T������������������@�A5� ���09P(�0��ȫ�"�0���+�"����+(�"�0*��+
,"�0��ȫ �p����+"���0���+���0��S�`HJ�*�0
��!�"842��ʫ1!(�40��ȫLL"�� �CC "����L�+��Ą*�2��@�+ �� CC*��2�0���J+�0��C2��C("
������ë���QA
QPdfO��g��������yd�?���?��p�A����xp����������N�οQ�~� TW�?p~�����Q�E�����F tJ~����_�� 
��~_�=�b�oOg����a���������?E�}̂���$��(��+H+B+#�$"�
,��B+!(��
,2
ʐ���
�ʋ ��H��+$"����2
Ȱ�� �� ���,(�*��� A+(H�B���,H�J��,$!,�$��"HJ���
��!HJ+P�B�"�H��4
+H+J
Т�"�"�@�"�H+B����B+��ȫ��"� ��+*̂��Ă��+2*��H�$"�B+
��)�+�B+ ��+��"��������D APJ �
���G�8����hP|��x�����ϯ���*+�~�������o�<85����������c�z�>��O�@���??��k�M��ހ
����P�}?�w��*��������BTEv?��L���Q��?���A���oI����G��a�h@�@����������w����>'�fߟ�|7��~ϼ�C^l? � }��������*+�����W�E~�9�?#��B��_N4�� X'�������A׀|O<	0���@�:��;{?�������__��~�Q�X0>��(����΅_�~A�~���
�2��8a���� ���9�>��. �     (      � P                   � wT�����S�B����I@@D�@(R� ����(�@�  
 �

$'�                                    �          ��� d��94����iJ2�2��� �� ��gY@���<   <� ��` @4�ӖQ!K��0j�����\�h���p 8:QE`ܲ�J���*�h�������*��p�AB�JX  8         � �LF�����җf�\�(U'YN&�U%�  5E�u�T(�4S�$�iT/^��Ф ���*�f��H�P�  �g��W-m˨J�� 5�[k�n�*W7C�+9��)7�޲)z� \�JMvb�s4]{�^a�<���@�T��  �        ��4\�uZ��`�j.[���ӡm�� �Tl��P�hq�9�R��{�{k[O �ڔ9���ir��
("�x  ��yj�[m9��H�� v�Rں�)Na�&�91]��s:Ut�p 6��ˬ��shN�i��:LӖ��U��Kl�V�  x        ;��quA��N��m�C38��Q�� �,ں�b\l���\�\ۈ n\ 5$�;����au42��A�  rxڅ^�\�H�� u(���)�e�5��v��5�U)u �v�9�viCstUѣ���@(���    p        ���M Q�ݜ ��:AX�u]r ` m��� d  P   � �� � 0 ���W qF�1�:
� �t�ˡNv�9t 2G�@jy4%*�4 �~#�%�Rh�Ј �'�U JR   j��&T��hL�i@�ʕD  ����ӎ8�W�p7J_���3	x�`3KA���$ I:�?���$��HH�B���IO���$HAE7�5<��T���;�qzZ�Ŋb�����V��:���m
`�JjQ�7��.v̐���6���}�a�w.YQ3[#��o��bG�wΏ���)�7�n��������]U{ÔX�7%�S�5�Ŝ�\�ܬ��"/4О8��D�b�$�ݗZݏ�n����d��H��;凔-߯@��k�h��;jٯ6ex֮\��Pz뛧�9�Ѐ�OS8����3s`4k*�MĖ�I�_njO>D��I󽮷�V�fܯ�L9j�v�L:{�ZR��5]���k)�Z� :s�m��&�]�)�ĺQe`�X���g�"���Z9$l�W�:]e�x�5Z�d��L�Ɯ�T�%G4R[¤[��v)�(ùs,E�]�DͰXYD�iԲ��	�\�Bn%��CV9�r#!fr0�}�轑�-��
�8��e9/���oXqAi�i���u����,�� s�٥��j
�[.�j�C9�b��B+�|�u�j��כ���}pЂ��D4��W�,���d;�=��Sq\�6ønFUc�� 5�uヰ�7P��Gs��w@����'d^G.��KZ;LV9Wv8�������gq붂ս8.��v�_�^�����\�Q�:hSI��ޒ�oLۛ�R�k1` ,���b���zTdǈ�CV�;*��3%o���h�Y�Sˈ��0��v,�v��4I�{O��vp������+��"�r� �b�Sy-zǌ�*@�!�\�nY�M�ou�V�7Cǐ�j�ڈ9ۺ���PR�{�����sS�����q×6�Sɥ׋�Q8��w:����S^�j�v 'i=�o�>��\�d#�Ը�k��r��Ϲ��M�5��F���KA��������>{P�RkӂS�Q�Vd�g =OS�2ۼ�8���sL�-���)���!�x��B��;�5�������ú�S�\:����v��!�and�L��y8P��l��WoC����= +f��&�;��k(��t;!#��A��w�+�}�����v����o�D�S��']�����}���m+9!�w��7	���{���u�n�b�L������U�dY�k}q�o���u�E*I�VJ�vM�t=�p��s�����}\+� �{Wv�䅮�-��g$v��M<;��v<�Oچ��v����}Uz�Yw�J>�^��wR]�m+Q�@��e�n���c�.�sps��p`la{��|M�2v7y�J�5hW�����\��8:ɽ��
L��o^��6-u,qLyy|�㐨����}h=��ԡ��v ��:� 6U�ݼN��٣6>ȟw0�l��ކ �չ3sB��M={���a����6�כtf� gm\�7=�i���Y��JE$6d\H�	���UAĻ��oby���Yog^�����|ʘ�n���,�{��t�Vtxm��\��SwT��/r����7�1 ޣ�4�1p,v��u=��.��]-vh��U�p5��/g��A>�'��k�c,h���3v�Y9t���Q.Y�7�[�)��m��ܦ�բ@�M�����#B��́�ڞO�pJ0��
��4@�:�{�I'�^K�/n�W`�۲B�ltEm-��޲M�x휴>�Ю)��5�f [2�Q�*Q7�DQ���3���g�7��l$���O�"������p�|�b=�Y����qs��/RTl���'Jz7�i�ǥ�esgi/w>|k�%�6��������Vs|B�0LEwk���һ���\��=,�4hǄ>K5T��d�KŦ
���^SX�&M�.��.�+�`�oQ���H�딪�O��g`�5���ǔ��=5��ΰ��-!v18�C�w��3vd����۷4"��d�{�V���޸�M�lX��pJ��`�U�t,+�`��ux�n�5B�w��Ζ���qm��"ѢJ����3�������x�ϮwL�2�ծ��U��o��%�����!z��܂�+���{����<���r����X�b����{ü5���~��t�M���I�z�d.d˛d�Z�0&�[�x�'�@U�i�ʌ�wN�Zxg;{�\y5�[sl����X͇C�r�����B�1W�F�I�F2HĨ�H�n}!C�O�)�rϴ��-�S\<	⫕��#6�;��&먑��KZS�oa��V�.x�\�=㥚qvת���=�<���>�_��(��Ѭ1M���3n;�������i&u!@#��/>�_v��.#�MԮ���:�j�o�ꎄ7�Eئ��x'��d�Vt|QO7�+����1�e'FK�v]�#�ุ���M%�i����.���ޓw�f��h8�v�;p�;%ѻmق��'sD���YǬd��dD��2�-�Ő�硤�v��u���)���sPR�K���%�Du�):gF)��w��#��J��\��;��q8{�8��F�W���lt[���'����}8��f�.̛��vߍ�fqҔH>`|+͘{븦wm��c&5����&��l�H:+�;qv���\�h�3kD^�D�Fk�{m�]z�-(v�'�Y�o����]������P���
M8S�p[K�+�<�y��R�h��ɢ%,�����f����4U�"�@�-�
�vv�����X����,i婡�5�g49����\�c
���xH���6Ι,���yO,�;
�Ӕ�JZ>�U���5ώI�ոf��f	�٥���.��2�tlGv	bB���ѻx���٘4
SC�;�,��׌�&w���
fDq�T;{{�v�6��j��,	� _5] �'�q��n��uR0�6d��B�h����&v Vr�ou�t.vS6��W̗�q����&rS�B躃@p
��\BA$[׵Gӫ4vw��)y��y�#h�=k���I� �{~A>�T���Wۃk|i�ܡ�Zm�hb���z�����4;xН!1-�r���/��j`$���޻��M���6d�Ӽ�N�J=��e�������j߸����Ԗ�ћ�M�>",}L4�{�bٔ;��ș�lZ~�e�4������C���#�'rP�{We�I �1����kM�WI�k�����8�5��l���d�d�4�{�Mʮ��շ@���CZF'��Al�q&Q�*�&�JX�w���ݜJ��uhmqC���/;�SMoc����g,}�I�j�����kL4`�lR��^NRFy��bv�:�a�f�Ȣ�Oj���՚��(�F��Q�۫�-���z�u������A3�^-����FW�穼:{���͚��%�;��Y��٥.����z�W3rW�:��1�ԥ/�8��gf��%�&A����YpV`x"�x"�pr�֜0�z����xy[^�.�z���k}�]s��ݯ_��]T��ݜ����c�2��I����Κf������:.ة�ٜ�xwK5�A��n��
7]�}�DM"a��v�M"��w�u��ʈ'f���α{�ӓ:7�i����ߗ��������''�q4B6H��Zr�t��ʛ�r��x���P.� �u�"o���qZ���.
����i[���d���3�q�e�����>�]cZ''�͖*�\=�iM�=7Gp���k'�c��i�VNK��-[��'GP��H�؎%}�X� � �&��l�_QS7웉�.l{� Ц�gwu-���+Z�9e���m��z�����jX��{��gt�i�t�6�ie�/P�X����/\khG.MM%��V�.��Ie�eˀ5��O5�q�]O�`2;u9;؋�)�X���l���@�~+�f�q�'I���z-�t|_�v���B�.
��c�x������GM2mK�{ٻ��{�ׄ�x^��AΖ���nc��毟J\��&ѹ�Gb�����{���z����Aª��rD��p��[�0!��,iWk˒��n�1�Ni���6�S��
j�+I��i�"����Q�q/�g��xos���%��q�;�X���e;��(k5śub�,}�h����C��Z}�	�p�#��G�'����Z&��TF��*��E]�/f�E^L)�1ݿȧ
�U��lZ^�s�jYӓ*��<Ө\���ZR��@�3f�r.x_1��Et,�
:˅	�'�u�ZX{�pnO�ty��N�l�:.E���o�%Ⳗ�t���GL�T��&��I��ȳl�oN>��>��
�(�鹶�˹{��}�b{��3�imI�^�`j� �MNݳ��p�^��J�Ȝ&J�ν"���.��>�How�A��8�#�{�bᚶލ�`��	�Z]�Ḉ��=�o-&��
A>݋��7�:�{�E�K�U� ��I3u=��s�'D:o,� T60:~�����n�#0��~��=��9�;}]Rn����{dS�i]��B�	sM(�-� M�h��j�1*ڈ�A�я������S�b�̱;�k�������ڲȴ�k�^kl�&�NapiE�VÇ�To5�4(�l( �dٍ�C_աQ0�7R����쫱��4<��c�_ҳ܆�;�����>Q^�=���7�9E{��f�Y\��2��:dٯ^^#�B%GvqC)<p��8���'Sj����f���ώX�t��PY�V�C���Yr���e �݃�L���B��S�8뽃pj��a+A�"T�=D�/�����r�aK��R�=��r�2r@k��͛f݂��nmC���U/%1U�/X�۽��ذ��;�dT,�Д�:����)���R I�x/n��\9��r��ˊW��Lhe>������-��ѐa�o9�A:ɮ�0(���`�;�sYO�5�@wvwb|�pe�5|����"�.�KV�=�7r��<}Ծ���mІ�l��n���O�f��v��Q�`e,���vq�X(�����Cq�AA�[����=�����#z����њc��8oM"]� �8�F��]�V�:��z�-��~�+�����u��/ψ�wL�����X7�:�a�Đ�.떬w�9���&�x#˷ü&���fAbũ���y����8�r��ܒ��f��s�p��79\$�帑��l����[^�d��8*ѥ�`N+�a޳�!��6=���i�Q����9�s`���!�;d�3^B)NŇ����n@{B$&o$	K'��	�YP
-�z����-cx����w�Wd:7��ӎـL��̏qU��k�:��t�y[�޼
0��;5R�;uV��q�R�)��ס;Uђ����U��a�u��b�WL��2R�i�:<Xy��K��L�9�zu}r����<f� �s�ӏfܗ�fi��p�V��_1����ˋ�F�Kժ.,PC�h��)R��L�E�/���|
W��s�w�~S�o�Rjz��8��=t��n��^�F��kNJ�6�Ѻ�"�ݸy}R3�{Q�T��2<j�wP�Ю��\��!�\_n:5��^ը;�2��ۊ��I@e�a��o,�u�ϊ����7����N�"��cw�R;Unt�,(�-��ޗ䷧u��a֦q�
c%tn�!{�^b^��Ǳ�ӄW��r������Ex�'�x;{wN�3���$o=�v�V�=.�Jk�VE��A�W�,bu��0o&m҅R��:¼�b���G4wM���(2oF[aga�,S!]y�ǤnT�gO���A�A�;]�y�D�Ǹ5�,�y��K�{_d���^W*�h�[�8�5p�Ҕ��@�%��oq�q,֣�(|4=�{5�����=ݶ��D!�KG�P�M
��l� wj p.�إm6>�7�2E��WY��)ϒ��tc;N5�\q�iS0\�&ފ({eך��j3l�.)�K�V�κ!G`Ñ�;wIs� ���9�
:ģ:�:���TK���q�\���󚆍�D��zc��gQ�:@7X��:���@э�����qĎ=��@�6̫[���Brlb9�zI'�k�)�`�`;"˳0epAN�[Hd�8�Ű�U���d
ұ*Hu��%zog&qK��CY���d8Lw�ƭ�tA�i*�����"x ME��(Qh�,xXph�l�
&��ld\��}{�Y�9�)�.��b�{G&*0�p�xJ^P�4Q�͋41s���cS�|J}���8q�c��:�����viMnoNr�m�Y����hp��q��Q��N]�8wW�Avr�v]"��B ��uW�w�@f�D	�>3���jf�Ȁ�Y�r����Xj�f�h��"5E��ȩy �Q�);�f���۴��Ή=��Q��w.#�N\*�3�o�Ȱ�yn�Y�c]��m�@�����L���E��q{qHݝ;�;y��N�s�eE��܄�D�2n�ۛ�-r���G�JN�z��K��ۯ�����Q�ػ/ "�*���qLo���en�e��sIw�����]X_ܞUwM�G5ٵ���B�oLO�M
�&�Ь�,�M��u�8i�1F'j}�8��K�Fg,޻�c�S�M�yh�qV���
DѼP���%U���@�����	 ��,"�E( ��@�,�T*@ )!��"��YB���I+ IYI,$�@����IRBB����I	"�B,	(@%@	%H
E$��$��@X"�H0R(I� �E  � �a! 
 E�� 
��XB�DI
�B�� �$�XE�@ +$� 
H
HB$+	$�
 @RH�,P� ��XI��$+ a!$ �ABI!$��P�E��	R@+ �*B���"����`
��I+ X@ T� ��H�$I,$d �� B �� ����g��Sm�5��i�8�o�sL��=BF"��倕���.d�~�򀉛���DC�e"C8.'qfd-�ڇ�Wj�����n��=w����o�e8Ȕ*��%����B3��;i��K*�R����I��O�giŚ��4��uٖ�.lH��Fx>�w(^t-�pH~"�0��M΀�fSwuNu���ƞkx��T2�~8r���ڧSӳP�K�[�n��<��|�rJ�8!��c|Ռ��x�;!J!U�cgcv�6%Ӊ���-e�^�Y�A˰o�^���u��~���ZwV����T�ό�:*݄��^n�,�/�}��}�]z�͓Y���᱀cFB<=]�)�O+���[ј���\�<}Dc����v3��ry��8
��9op;�^��t�������	[�4�x��&=Ѻǀ��cu�3w-Ԛ��� ��Е�tNn7���^z�1�{��ҭaygz	�H�?s���{כ+u!"	���F�,8׸<�L������)�q��O`�-F�ׁ[��ǧ�ó�ч6�O���b�­�N�rb;0�rs�U <ܛ��.�O׋��ý��\B��޷����-��m`N�҅��ܢK=��|�4ll�v��@y������W��9�= }7Ch�xn��] #�kx��ʘ&.���}곱��p��$��X�Ou,*�!~,Rݸ�Lwr3g,\ed��l�G �Ly\�ș�c�.�7=�)��#�@|qb�*˾؀�^��7jc���E�u�	R7޻~����B����suN�o{�)ݹ�C������&�F&��$���o�f���� �
�5'��
��S��͜����Mܙ�b�a똼0�{�i��V��:ж���]k�Q8;
f��1!Ψld�mG�a�Z�m�����;1�-b�P�yr��RW!w\��+�ϩ7Uy:v,}�<{\k�'(zsʔ^�=�k�N�w�_��R�01����.�slY����W��v�h�=�ۊ0�ϴ>�y7h�Vlؽ�V$�<pٓ~*u�s�n�[�`�,۞�
�w%������D���V�lrl��x��n��A��o"I�t8]qq�<B��8oț��__�9���F����Ht�o_ Xx{�Zz� ����;s�� m����){�V�	�cؗxR�e�m(�mf���<�vx����S?w���e���X�;�{;��K�b�Y9sj@Ft��1�T�gjK}�Dh��q�^s�4��Y��=�e�B�e�e���P�/&w/4뷆S;������3���:;�ަn�&�<�34�*�7��,/"���r��ߊi��چ��Y�O$Vd�۾rxøM��A��������k���u�Y炿V�T��jm��������K�%_ps��L접�kQ�hyYT�xG=M���z'�w�B9^ռ_�)�n��l���u�gnq�Ђ�$ߣ���oq�:ǽ���^��&�[���wa9�{�����P~G���;���զ���j���^���y�N���E��`���Uh��w¸�t�F<���[�`l}O��[��5Vֽ��{�h�ݖ�ɑ�'U#f	�U1���szS�R���E���}௄�����z1Z�ٓw�z���⃚�{U��y�N��^Ax��=�l�&r c��t�N�w/z�Zx�U��'t����V���Xˊ�d8:V"jm��鍗T5�v 䓞t;�����Gҥ
�w���VޗG�oqy�0U!'�J�(�{�f�n�s���w2��;�$pD��l�$��;��(,�f3Xb�bg͜�l9�ց/��!
��L?S�n�)][�����!y{A��]�Bw�A��7�7:
>kT�Nr�gj���[Y�/6z R��oi��B�P=�iߣ՜w�M��{̋�:��Bs{�M1�m���R�K�YFL̨����,�*�j4cu�W��ccu����y���qa�����z��ܝR�_zz{ݍn�>�v��/,��{^i��<F����7V�j�o�]�Ք��Â��'�NxbԱ�՞ݾ�l�]|��uO7��a���M,oOy��Cs�s[��զ���1b�����1�6D��g4T�s�K�Br��l(��P�g��s�g��{[9ꓽ����qt�;�;ѹ���0��t���ͮy��(�.7^K{��a��(��^X߽�ZLK�O��[;^�"���:A�Ֆ?iW���w����3F�
�:Ы�xa�A�/$�#1��[|�Jǻ�V�wb�vE�}�d�:n���z���6uo'}F�싗*��|r=��<�0��9�H_z-*�JdM�*�uθoHȩ��mߜ�͙�ĉ;aVD6Xfq�0fSJ`d9ka[zN��V;��
/sQ���9�o�n�ڨrv���M)�r�z�o��Ȭ27,J�1���L������ؖ�ƛ�`3ȿ�yU��N�b��h侖L�.�|!�]
�F����N���/���E���5��Ɲ���=���{<���>�����sh��Oy$����g��ٲ�q4�2�z)�=��;7�$��:�<�V��+�����u�w���{�g5=�Pf����R��k�hg%������S��=�=[�P���sϑ����7� FA'��o�tU_#Y�p�F�~�PZ��@^��V3����]��"���ya[e��3d�i3���c>۹1o���t��=Ae�y۔��x�v���QY�5��b6jܻ�Uě�3-4mD����&���z�^�ۺ�v��8���������������ށW�O��wӦxw��f�A(����9qQ�f���r�L��&�&�CѮ�����w���Ƴr�LgIk-�{�у��luI��u����S3�������\[���ܴ�����9<6q`�l�]X%^���_M�x������/�{<B�, ������Y���w�)���;���u��d������n�X��o^�\yNnzyb�����Xe�~�Á�Dm�>ӸR��r�_vۉ���g���O�xEl����=���ĩ�Y5v�~6��D+��{5]���f�79^ÂM;�W����`r�]��<@��3��=2Ĺ+�����T�ɜ��=
�T�="����|�ӻ]͜b3A��"�*��+�)�s1��kn�t�n�Lj��݁W-,��W{y�j>g��p���u���j^�Ax2#ok^�)��d���TM�/��g��۫���{y�վ4��9	5�XB{a�_��*a���w�{]@&Po.1�ν�
��n�CR"�cD��c<�vF�x�ٍ�	�Zc���������u��<�쀂ڶ,���e���Z�.c��f�r�O��Q���B����6O7�z�.m�uN����k ����wrVc�{N=s�j]�g����嵎�{A��z߶�+P�do�<�����5n�R������f��K����;��j��{UA�� �)��ף��sfd�o������ԛ���'��Π�<Z�����[�O�xE�O���v��{O�d\����䷽�s�_wN�R��J�v��E�����b�[8h]�i)��$`��g��l+�����Ov8��l�}�_3�8�n칻��3�Q����כj���#����'F�Mr�e�D���o\��IC��=���s]�=���\�f�X �z\*gW�
���r@6��δ<�ľ�@���G{�ź�[8�3So�j2�,�㾞܅������"H���^���[n�u���w*p�������F�׾�xK=�����ð���K�F��v��=���k��4[�6�Ic)���/3�{��s�+�X#���{�+��J^��ћ����w��׋5���%�ysѼ��rՁ�޳D�j|�o�>�ˈ)�Ԯݞ��� аX�M`+~�2���z;&!��������4_;�9�[�љ8 ���֎���XS77OW�ּL�pї;�j����71�W�4���e����k����<�tK��n[��2�������᳏qP���㰧gF�J�4�S
��WX�8�]�xxrV<t����$dݯ{}��o�<h���x��Yyg��^�_�Ǉ���y}��@��k�י�ǔeit���E�C��R�+��d�W�������S�/���7���)d���1ԃ�y��G�m�W=;�n.�ν���w��|��I�ٽ��eDHy� �֞�1獪���
���Hi��a�����s�J>1���1�z����r��D����c�'<�̞��'���/)�NN��l˹�d@ga�L;h�2Q%)�9}�sؚ�^{�<!��b���?N;Ȝ�=�����b�ˮ}k���O�z�^&{���Gb�y�|_�y����[�����^�^M¼#���w��5	֭E�x�����W{[�����uU�^��nra����߷��p"��tw7ޮ�X�Q�y�ї�>��Ul㬦j��'�u?���7ƭ����o���r�E		z��E�!9^r�����?s��Ξ7=�(S>y�3sm�����I)A�����n�k�����z���UY^^0Q���\=��)���D!ּ��j
4���{��?W<�wbG�X�#_�u�󻫔�L�d��%�.��ze�����/4�`�܅xw��~�Zt`�)��;��s����s�X���o��Ѣ��α��޵R���y�޺����TٕX���n[<�9V��u���{�)�r5���5�m���D3f�{m���ݭ�4�4���u�ﱻ�������4j�D%�["}LHn�:療	��h��==b�1�����Ӟ�"t�n$L�曳$<���Ƽm��b��秽���60xaY��E\��J5�^�>�-LO'w�ؚ��L�~����#�7�������Ѭ��X=�[�O��)�*��8"��*�f���o;���ġ�z���R�d�~��[$�Ͱ�y��k�'�!�6���u�\�o���vZU+{^i�����%D�Z��Nlu۹a;� g�P�:�m��huz��j���S_��;��wҰ۹���iS�ἩC6t�8��y#�g
�P,�Ӫ�m�n�����;Օ�E�o5�5���;������#+���-�#=_��B�4Y[��o��݉:�/�6q/�< ��ͮ�3���5c�0:1Jz�ʝ9��.FQzܱ����Z_h#��mL��1�m;�/D�Ә�gr(�����<��ڋ���?�N糕�s�u�Ϯ��5x��t�6�՝�޳�܅�{���V�73�g����{5?x
"�6cʛ*?d#v�g}{�n��ው����7=�G��7�!Snn,/l��e��0�xdA�u�"ߜ�'>�<��������ݬ��HGw�������N��fS���(��{L�O��K�%�/"{�w�p�A��w�+=����^�h���=>��r�/�Q����븵�߷#1n�>T�Y�)�z����F�s���uN�Ó��)�.�Uz�*zS����ιE����Zx�������&z�l�q]�N���|����h�[�mx՛�LM�ޜG�ɪV���.��[J
n�zrw/Ng��ǧ�znK��ׇ��Fr/�W�Y�;�<��S=���}�&*˾=�
w	z���� J�tL>�{�x�6���>���^��;�Y�xw��:�;�Gd����I;�դ�Ӄ���R���"r���3��{O�bO���Y�ݻk�.���1͑n4�W��ތ�v�[2jۜ�Pogg��3|���7�!�쫴7�P?�H����7|�G�:{ ��=]�=�<�p�q���G�GK���t ʹ3_wn�=dn�g�,�8�t�&{��^��^6pa������n3^:������������{D����"��'=��n5�,F��j�
/"Y�gn�q���xϴ�xq�I;HwXV���p�a�MZ�*���Am&$��o�v��v<}�G�x�8��Yۜ�1����'��I٫9F�6��Aݒ1�|�����T�yG�i�O�}��c;��C���)^��Nn�d�)�����?i�3R�8��+g]��Yb>�r)Ö(�y���\q���9Z}^��7��]��R6�e�vE�;�`8�j�E�T���xх���-Dֺz�f���Tm52X0��ua}P�p�u�͍y��{zu���B��崎�����B"��1� �F�n.^�$k�!�=[&=��[�K���lS������,��{��9�퓷oR��#\\:����.k/R�����x�)^o����6>�#}+wM�+���b��z�f��HY�yw���/�K�̒�~�����)�=ؤ�o�:�����>D�{��t�::�X�c=ق���y||�+59[1!3m�G���p�Bس,N�6z\*�wi��Nu|:����O+�<[�o�8���O�y��{�}�\G�}�C�_w0�����Se���Ƚt#����^z;n�שs�9��ȷ��8|����w��<o�g�}TZ%�l^� ���	���n�SiZ��<��h� �c��9M��NŞ��L��/vY�ܼK+�R}���{�p�
-������E�ݾ�!�b�w60T���gV�Θn��ǹ�t�3f�s5�K�bt��j��N�m���HU��Ġ�; �|�+E.nWۗ�m^�v�nx�<���}9�����׺�O�1F�@N�DW��哋Ż�bܞ�p6aݹyDWh;n_�~�Ok�QE�E��7S��OAC9�h��mXs��ֈ�6����{���{���{����~�-���j�m�6j��l�W[�n]v���������8�"�1��Ҕ�5�\7�Z�huxݹ�p��m�1Η��۬ۓ/<m0�䛏C�6ތ�$�Q����qK�ֶ�\X�y. �\$`���5���G�g��aM�]��5��y@�
DL��nܤ{q�qs����d���7;�Hmm���7u�>n�l1�y2ܙ�������7[�vU���vxm���֍�%����k���0O�0t����;x�k�ˀ9�cMm̓wA�������"�8�ydj&�Nq��Ӷ��'s�tvńkur��W��X�q�=�h���^y�ͼm�����z��/n�\	���`���_n�wQ�{NOX7nx.S�Vs��\5����r��ɷ���I�e�h%���_f�ݝ[`�Y:���Ď�\����;����t�l�e�Gcs����ۥJ�ڊ��p��Pq�멛qV��S[��h-�'�\��k���-q����Q�`�v�\qֶ@cv��Pb����y�7�*�;R:�{qλ4r	�8�rِ���f�K�[�S�n�#��٨�:��@�v����rv�G�u/jp��� 5�t�[�U�B�X��Ҽ4���f�m��=:5�·���1���v��18�n�7n˳�h��<����v�ۺ�ݶ����G�ϳ����r�����څ;6溞�S)Im�<n�qP��'s<	=E�����[X���;Mv�wZ��=�x^�� w�vgvzC�Y��kr���n6�]�A�M\z�X9{)�g��������u��my�X5�+�"t\��v�K�;	����8��O��]�l��v��2O�=v�`��n3Ԥ��y�	n;eݝǆ�q�c��<.�m�s��L�<a��<��۞�+m�rn}-ąv�g`��r=��;C�}Hu�\�v�1�t��jN��[��g'q�M5ס#n��$������k,�ϷS�n�5��w��iLl۠(V��xm�;v�b�wa�M���7T���=��-��Y��g���ڳ�w�=[���7`��a�<��d�3�{�-n��!��F�g��N��!�OB�6�
���Q��:�����'6���=5��r\w�˷\l6�<�Y�:ݹ�ۋl���܂J\r;Ƹ3i<W:T���Y֔ͷ�gx9�	���u���F���V׉��x�ݻu����M1=�Ԝ��u�4�n۱�<0>�#V爹�nvݞ
r�$W��s��d;.��l�8�O��[t�6��q��/Cu�V]���!�:�܍y�[���E����C���.���.�L1Ѻ�"�n�a������C�ҩ�л���Қ�n�x��t�ո����B������)ۮp�����-�=�݋�㵳��&N�q��mb�cv������!��;\��%��r]>9:����uѮ.��<��Ln5�77kb����gx�nܚ�n�L���q���ܶ���ښs�2C'>�Cr�akn������GGi��G5�`^��wN��������!�
"��h��y8��n!�b�n3�.�݌e]�E��#�}��u�c��qs�˷Il����y�zŭ�m3m��=�w<���us��s�6�sD�4�G=�n�e1��c/[���Ӟ)z�@r��j��d�n�W�l9qս;m�8�FN���ac��x��y yC�0�/�b7���y3ӫa�����&��v�[���1�]<^=�:u\�.��I=��Nޒ�<v�vzU�8�#�36�V��]p�tg���u��n��=�vj��k��F�Nm��=�;'`�4��c\�s����ǔ&�� ����.�(3�	�4�<n_ �睍���vx�܉s�y���d����n��㍦܎:�։_m�u����Gj��.ǳ�/s��κ4�$�!���rk3�c��d�X�U�ۓ��4�����Gk�j6#����ɮs�0ـ�:̉ �u�M��F-&y���1I�8�τJ��1��`�B��EB�7[c��t=e�1��v.���3ظ�V����u���x<E�&�g��۝��NwD����Q�ѹ�6��[����JB̯Z�={q�����LO=�y������xN�0=����ۇ���\jx�D�q�E������Ga��$n'��j������`�=�s�r��m]ZؤuMvۜ�=�9��'i���;��\{j���q&v�\u�����]v����[�1���s糮X9.���l�Ƚ����;k>�k\���8�:�	N�ny19�>z�(;uG;��s�]l!���6�8���<ݺm���;N��c=e�_Fܚ��/!��:zd�73��2�뇕�ls�!��nج�1=:�x�.m[ی��#l�������N�F:5�nܽ�D�ڔ����h�k�ǻuب��!����;;���+Hx���[[m�������OH͝^Yn�JnW�<p�;���;v�MJ��)�d�� �ά��4���i;&��[rr+�g>���Иח�Ny�`h�y8�'F��_l�=�z���늸γ���m���G%nj���`�8]��m�V���,��9�=\88/<�۱��H;==����pǰ��k��=z �ïl��GL�̆wr�U���s��c�n-���[��f�%Þ}[��S�7d��ɜ��.�c:�5�ێ8��ϋ�ֱ�[�Z�Zu��<��g�����s܇`HƸ�vX��rl���]�x�[5��k�]sьv;Nu+L�u�{yw/�tnq;jδ%E� F���G�����<s�Z���tC��A혫e�Kkn���v�Ci�;,�Br/"�m�y�<Q�[l$���<�Ϧ0��6a�憏m�<)���c�����z�t6��bQ�p6.�dxD�dnc@v�a��s���^.�a��;��m�<q��v�M�n1`͕��-��e��n�:w��N�z��7��q�E��C�[[�7���81���6�X��QO;v��/=�@�ψ��.s����m9t�;Q����N�&�F��p�=Uf���-�&ۡk�]���En{Y�ۚ�8�ɌA���;i���ٸM'�ۘ_(�[�u�Gu��\���Fv�6�s�ۛ��wUW>ܚd��'+:�C�8棷/6���<����!�n�xql�#��]p�������4�ŷ<m���g^ɼݽ�NH��îq`��LwnN�5���3l�R��o:��
��=�{G/v�ny�"�a�p��ս����!ͦ�8r��Ͱ����u!��`��:έf�z�cq��ɞ�s�p���zN������Սbn�&G��cs�F5�6l�)xq=��<a�6�/m��M#3΀�ȼru"���;i2s �<l.oN�m]�m{s�\\vN��6�t!�FC����q��D�cr�A�eGu��V9��]��N��`��Ř�ɞ�y���Z�ʝ��Lms�2��u87`�l�O�\�4sѷ�v7evoH�#�HoZ�tZ.|��;��7hKqih�su�㎍ڃ���FWt���e�;��k���wpu�|�aFk�׷fϳ��s���VC��ۓZ�N�-��u�k�X�YN��;a�I��Ϩ1�<�r;��I�]��b�ݜc���m�;y���u��9�xy�� -�]�.��g�;[��ٓ��i&�Ŷ46}�i��N�.�6� b��cl��:6�Ccw���:�Gg���&�V��ղ[�+hC
�Z�Y��v:��c��@¶ì�l�hb�n�է��\s�)���\:w;n�˯s87������0^���:�9�˜X.,��;����w+�� �mͩ�u[l�@^h��垓��3���B���Y�W���n�A�	�+�5�)����l�t��i���Wt�:���;;[bv܅��ѻ'��:ݹz��]��K�u�:�7l�E�k�i��v�=:�{Y,�,n%�x�S�m���q�A�t��˪�v�B^�i�s<�vx6!I1���!�rX�z��m[bk���z�����{��K5�y��@�=�ׅc�֚ܪ�����֎M�n�.ݸ&;`��N�ۭ �L$m8t�qě�{��[�6��]���T��Y����k{\6����<Z�=��x8�ɫ�󋞋�����}<U�	���\ey�= {��\Vޒ����v&x�v�ݝ�6�;l���������h�2秴��;;n��ۋ��wt�����l�v�=Rv�͊������۷OH���Y�-k�n{ݳ�Ui�ݚ�%�ű!���ޛ]s�Xъ�c�p[p��ˍ�:q͝vݖ��ŋ�:��>]��\�u����1i^-G#عxW[���b�@8$J��gn�GP[A���{x,�c*[xN|q�cv�Nj���]�!�1ع�x�g�rg[K>ɷn�v\�,�͎�n�<��R�G�q�`�px=�x*�퍹�2�E��/9�٭"]���{pp�'v#7��S�np��av�[�����6N��SDX�Gs�fܝn.�g�=u�]H�k��:dz�[��(�Z�on+6�n��e���챬�kn�1�cnC��sۢ�W!��Ѯ�:.�vY�mf�{k�ֳ��6㴣�۶�#��!�:8�c�p��'��ݢ2u��5�C�q��OWgt��At�Кw8�9�wk�����N�@%��(�÷cF:5]3��s�n�QކY��Ɖ�6�^s¶w	��.,[Q�r���9�Z^:��$wD8��C�����o�f��L��mƅݛ����F��z����u���=m{r�����D�j��U���v��̨��zKvkf5�:5&�n�9ƸW����g>.�N8���'���<�\k3ڻ�.�ݱN�)"-=OK۷n{cn.����0��Ԡ�[AZ�Z(�EV%h�m��T�22ڲ�[PF0X� ��b��e���m���Pm��1�b��Z�Z�Z6" �Ȃ���*�J����Q���(*��DA�cZ�ZKb[P����J-+PmiTTV"���%�,R�("�b�,E��**"*,U-�b֊De�B��UT"1TY�4J�DUA#m�E,V(���*
(����K*���A�ȥd�Ա�U�h���l,QH�
�
",UEcDcm�(�
�mE����*��DTm��DETEDEA�P[eb�Fڂ��b��UE-��DDm����Z�-h,��TAZ�*PQ�X ��-�Rae��6�F[e�5�"�kU�R�@���QV�"��TAX���R*�0R*"%�DU��m+kb�cZ��Ȩ�"�Ŋ�b�E��Dc ����$�:�s�g[�{hu��[�Ý���51��V۵�0vz]I������9`�vkr�m��n2W8�j��ގ�<�q�3�[mř��Ż�u<^�u˶���Xr:�u�ug�3�^��=s���T��&���/y�sgV�Aݞ����d����인��1����o�e=����ɸh�ӻr��N�v�����6�g����qK���'<���E��ۋ��;����r��L�{v��+��terv�=ӱts�����]Gf��n���7&�����t�v^�K�b�hD����`u��ǣ�h��\R�cU�uwu�u������q�n�M��P����i�&����i�xU�]��x���vn�r�����̼��E��c�g֛gm���l�󮂃�dvWq�7m�����''=):<��q��^���,�q��^�o;�O������N훈��g�������nڡ��ڒ�ti��;�FToQ�6�^���щ;	Ή�v[���x��nt�,=�$;l�v�'q�.v���V�6��[�s��e2��=ny糨��\9�nG��(�c��|�^��[,��|�������ֶz���ݭ��P�e���Ѹ��n-q�ē�b�xGz�6t�`��h1�y���g�G<�nsĹ�3͞;�u�D%=5��z��^�Y�Ӻ8@�#�����>�˟��a6�[�wa���;�95,j���Ç���b8:n��p���c���h����2�z���^�v�S9t� ����q��3�gQF;��Sgol�3�+�8�C�vՓO�o�s�s �v8�㳙�!\m��k#zs�pqnčո8S�����vm�[��]xs�+�q����`��[2�K3��,�g\ݹA�g]r�{E��r.���u�g�y�V�� u�J볺"]��r�j���nۦ�d�]��պn�����{��X�7�v������L�0��n��;lQ�v��pm�ݰ�M��s݇;�S�����g��q������Ôݹ]����#�v6��2����g+�� 	����l�7n1���܂���<=�0��v�6�9�le�nO\q�U��^�]��nۑE�&�9���e�����ێ0��r��yp��9�n}�HK��x�[���������$P ��􈉬2>�}\Y��o.����9�6N@6��AnG�wFJ*�ӈ-�É����9�	wGH^2b�����;1�{V��Wjl
T�
!U�˪��#� A��ȝ��B �ts�$�=4H$���n8�D$�B)�ГS[w|�jQy~$��4H$����y;B7*n���|دL��
Z� ZpY0�5F�c�b;6�^�C[�f�Dv`53w4	!fGH@�b:�h�:�&L����Dv0P��A�	�sa�:N}�N�v����=���x�Ӈc�ۿ~����t@(��ۗW<	 ����A>���я6�����ĀH+66|L��mx��f��^רL`Rݒ&�s{`����x`���TF;��c?�wM�R�ތn��8;���B���f;�%�,��p%��S�d�v�p���U���7>��Vs�$�וD�W��D:������ �VH�&ـ�P�-ɮ��H1Ovhf�՛�%u��A�Y�ҁ�>�w�D�h@�BI����.����Rb�h�:b�I�k��$���ryTcB�!*���3��@JF!4$�V�Q��zk�{�{1M��㍓�O��W�y�M��ӛ��Y�c�p�FB����6�.��-��������)�xۇkZm�=v���ڛ,�m���2	1�H�{��P9�2X78�S<�l��−D[�� �""8@(����}8%t�?^DWGb$�cޡ@��=TH2��[���S(��^!���g����Gs��� �Ga{��ce{�S���C`���|�bд�"iN(n�	��!��
�2a���
�kV��n�CL`���Ŷ7dʺ{wG�$ƽʠI#��Ux�K��[,&T2b�����N�A�}�D|{fzhI]Ѷ7\��`U:H����y��A1���뼪IY�����`*b�����Pϧ��%wF���`��<�!$S��zfMt�x�m;��Gmv���g�/d�=X�m�>�?w��2bp�C����� ���$��ɹ���8o=}9t(�{=TO��DYp��e�Tj'\�|��vz���s�H'zgj�$����,�"�0��f��5:2T)F"0@(��nD���	�]���*�>�0�.��7��Q �
�� ��!-�0[*h�e�9�a�{B3}4A�����>��_%�?��U�]؏�ʫ������Ś�����n�:���;�B�*����H�:F���r.*<����'�4�*|삼����[�n!Y܀�m��P-ɮ�bI*��Q}��.�$��˩�H]���s��V+��&UWd�@4� C�C��P�Gc6�v����&u�Q���+C�w�����������%�\&�*��AY�ĀH�!s���yy��&�Ze��� �Vw9 ��er���$*b���Ɯ%)�㎅�ݘs7���$�ΟH%s��*����=ڨ���$-y�����8,�j�j:��J�"�ӽFjg_6��f��
��>>+��Rh�F�(��C-؞��Vuk9�t��|or\��A>T���'��U��ίZ�r	��D%`�d�0���^��s�@펪�����}R$�U<���>��"����L�O������N�D൜Sg���K�k�#�VHu	�Z�6lZ
၂Ƚ�p�xy��s�F��XR���㵌p답�i��]��у)���h&�M��t=v���;q��9�խj.m����]�k��l;����ju�vq��ʼ��{x㜵�=z/]�R{�͸�d�iӴ���4��8�m���QWrK�;v4��۸2��z,5ƹ��y]F+d8�v�8����O^&5��{�i=�v��bM����zv7l'Y�@sA�^Q�11]�3����1���Ė��,��nvw;�y��!��s	F4�2�2[�so�B���$�w�uPz��]{x�i���i��oy���W�<
 @���o(�뵳uY�t�cO�!oOUx��몁&HT��g;&�C\(d�I�l��j��I7κh��̅�|���^�H��림HZ롖�AP�j���c^v��73��0E��W��;�l׉!wF�휊�Ǡ(ٺ��P���C��s9W�+�����$DLt�m�묭�#��H�|Wtl�y7*�A2P�d@*�q1[U�u�eQ�qch���v�k>��;������B�$�$0[+x���
$tul׉$����=���D_:��;�r��z6�����0��C���nA���Da��͝��u�LfUBܛ����cY�	1K+k�RN%��剬�_7���{��%�\�}����{vo1�MrNMl�H"�j�#��es��4�h�Fa�4���9�1 �$	x��+o� U��0}��5g��(�zG�M�VЯz:4��1�!C%2��0�m�\^-ڽarWZaY�	񘙩�I# �/��� �N������rK����Ζ�Q0�&�SgĘ읡]��N�5W]4&㣧�	�9Bi>ȥi���lD������N  �3��D�̾9�u�`Kn�,�!i����r<}����H�	�u9sđ���H'���@�S��龪����}U(� �$0�eU=��D��g&&��c*k�z5�I�w�^$�qBb�쌛$]Ɠ�8b DKr�F�>)�Т	1�$��4^�"�!P瓓-ۙ��K��d��s���]{��
�vE�/q�Z���p&���ڮ��:w�QI�v:����QW;P��tt��*���3ڀ)s��kyM�	;�>�deD� �#�r��{�m<��.���M�o\t���|(d�\Bp}S�V(�M���%�gm��DI�f��I$�ʪ�F�V� k�Vv�sq&�+,��۾� O%t��Jwl��E��Q]����|r.��򥢈-$v}�s��D@L2ɐe��7��Q�$�꭪1Wlq�'�t�3��H>1W�4	�8��\$C��	����|K�[�t���s�I ��T)Do7�8�:���9VE��{vh��"�Cq}�Zj���ڏ�Z_�{o964��ڪ�wUuQ7Q��0[b @��b��Ӯ��k����nW���w��ExWf�ʍ<0�"U���i{�����pr_{�'���(bm���7�`b����N�ѲioZ��U��/��K��^�D��s<��,P��
��$kAc�TB�b�OnUQ>${�Ni�����$��B��[B�vk���!q�N1I(��R	����O]��� t�9�wN탈k{2py�����qP���q��7wUD��[4���p�y5&��|;����	'�q���(s��D@pYd�x�m9� ˇv�mK����γ�� �:ٯ�OFk�>;��goػf�4�8��[H�	�}7�0�Ѽ�|\�=y���r�$o:�I=�H�ɂ�@�d�a �P�sk��aS�15f�	7��4���GE����와\[��5s@��m���nA�r�F������d���P�O=�> �}�s�@*wBB:�P|�k���a�4��\�1T�Z�I�rtYܙN�E���['�ڣ�b1Z/���rvS�3ԃ��g�M�J'� ��Ef�=rv,m̗E�7��۲�Ӆ!�2mn��H�<�r�ś5��;Z�u6���n�|��.��w+k���xxŷ.���)�ʴ��w6q�3F��rżT�<�U�� �a���}U��]�ܻl'[xǎ�㰼�xչ��M`y�Ʃ��ݮ=�B��
p��61�>��L�K�q�xnxLټd�9���s�hN.�m�u���3t��ltA�n:\K@��ݭ����ޠG���n�:Qŋ�md�P$�o9�$���(d(ܨ��͚�B����$N�� ��O�%���>����c.6<��D��ʺ��I$�}�$�H�s�@��9��Gt��r����#\�"��&���~�y����3���!�9�y�	"��I�r��P�����C��	��nWM�n�6U�|cz���|O���P$���u��	[��k���O���! Y0Y)TVOW����S@���Ќ��`���	��U�F�mP�1�}��.[��Y��WH���6�D&�m8��u�ۻsG���M�T;;�54�<vݶۏ�����7l0!��x��9� ���Т	�v�QL�]�g�� �H|�*�"���A����*���Ux�"(!Zr�
��w�rhs�r�5!�Fw?ç��Q���A51���xoe+�m?���Pfjz ��1Q}3щ��6j.�I>x�(W�]�SDGh:����+�$�K�H�d�0S-�pD�n����H*�jh�|^L˓�н�[4	v�H%omUD=�9�J" 8,�j�S�x��y|	r��Ě���$��,ު�Ot��g\p�����$�P\4Hp�a8y�8�O9�V:�l_>}�h H�꺢I;j��{�X6�9د�������~���Aw#r�C�dPɏ������5`�=��8;����N{�g[{��t�Q�����$;�gǥ��!VН{�@����U�1��a�`��s�{�\�r���6r�TtdLG.�w6	�+w��@� ��S�1x�DV�$n<"4�1��P�9B�_=� �F?������~���|(�t<�=2�Hn���}�w��}�/'9>2��ϵS��܆k�cy�TFo�7Q��4Gz�l�����3��&]c�[����I��c�x�)���}�n7QvBQ���^��O.Ey�u2����,7ݭ(�Z��g1�G��wv�0�w��z]޹���D;�{c!yم��|��wWf\������a �x�m77��I>kaI�����l��)6~�,��EIY�<]��=��Eت�!ݫ.�dΆ����ރ(���P���<"����O]�]��lB�A�tJ�$U���{�w�����;[�vn����v�����R��:��M<a�ڤ񄈗�U�l�GQ�pL	7�Cn=�&�q�׆N����������r��y%����t��RO3no���)���\!L�2����{*�#6*���{FM��4����4�۫��A�nd�4!���0�H�wM�S��
�ry��:z��̽m�Ʒ֪��Uo�[��d�y�z�!���d2]LcUIf�o$'.�!��K�]�hK���^{'�$��%�^�����=�[F�@�X�RӘ%��]˻%���	ѝz���Ü�z��oi�b�G��N�9�V���5�v����BA���݃&�#ۯ��
94����[
Rrw���s�������ykܺt�V/E;��������<��g�=��Z����ݼV��qp����va�#.vs*nh�iԙ��vSf�q�KV�3��-͖u	j�a�'����IX)DA#F(�1������kTb"�UDUb��((
��("�DT1A��6�EUQUQ��((�F*�DV0ekm�*Ȣ�*+cR�"�iB��Tb�T�VDF1ATV"���U-�X����PDUFZTAATUEk%X�mTUX��X**��6�m��Uj�،+%`��"AAF�*�PUR+mb�eZڅE��U"�EX(�(�%j��"("������,R
����X*�(�`��X�m�F�("EX�Z�AX��J�"�V҈5�#$U�1QDdkTA@b*1
VE��"�bł�UH"(�1Db�*�b���"
#"��1b�"*�*�`��Ab�V,PEb�F,��#b�"�UU�#��*�`���Q�H�F**�EE",UQE"�"�E������X��{��,X��o3�N�A)%��n�$�V���nc��WT�>9�R'Ē�w*�xa�UT֒*�n�C�'\�D�h�S�b|C�ݪ��p����x+ �ǕU�I����;���2�S�Ȧ@)	-��j(�u���϶�( �y�݈p躧\�{��߽�@��,�6��fUI��rI'�k&�WgS��!�Р��rf�R"�D�d�����P�-������eyr���H$�$�H絔+�z_r,l��N�u߉��1��6��nA��s�H�u�� �N�29�3�cWP�s�	$ާ$}�k(U�AFP�<Ѫ�����iF�l	�^'���A �O���==�0�	��r��:2��ҋ.��P��^�D�P~����s�j�+vumVn
�L�aFm5�r�$����:�;��M�Ё�!�'�RKAlC�$�;^�	��[��,u���gP���	����'�����R���jS9up,�c[p�EA���(2�Nzы��c�m�q�N�u�_/ns�:�XVt>���~�0,�k����A>8��E��U^0��v&��/w*��Ld�|O;����JGay�L��3ەC�Z������O�	>&��U�GOmU�QٺC��X�b���@�`�J�O=�D�z{�h��y��e�}���Fu���۪ ���P���&��X-ϏR�wCmA�\ݰ_a��323ǧ�ꏉ'�9�TH$ŵkc��ӣ`��Z��W���
�5@v��W�$�z��/��ȣ��]\�$��H$�ͩ�y�K��j/ w`���_Q�A�|/U�Ȕ��ٷE��BK�W��Kt]��7�ױG��x\��nk4gCS��yP,�Oyդf��i�A8���o����Ѷ�v���,�&�Ou��4:,������|�n���{pd���m�o��8ؽ�Gg�V�E��v�����$��׍����n���;\�n����у5����8��lfmSѦ֓�{^;qGu�\4��[�͇issrm�;v�2&d헜���m��W[5��9�#��ɵdծ۳���tݎq����uZ�jcO�=���՛����w��=s��1%�ݻ��~��} �T�p��f�j��M��$�G,ځJ�gVH.κ��H'�z��I� �1��&�:��B��a���3D���s^$�x�԰A;=�0�vE�6��D�@5����Q>���O��>7��`5�X4������͘��gЄI!"������n��W_MA><s�$�G=ˮG0��4s�~o��ǩ�U��t����{1���׫3,q��0OMuM'Ol���n]P'���r2��e�V,�5��u�:d�g����g���:n��F���5��XӁ lB	�Uי�T$�g�e�H$�˪��ıM�s���g\��I�!Y+*A}~��(�u��U�T�p� �B>s�>|�G�U�?q�y�A���b��	\M��7�}����
<�9L�v`a�o�=�;ǖ�W/(|�枎g����3�rnQv�A��c�_��;�y��h��!iHT�߱�����n T�������P�8�YY*��ˆ��:��p�3���D#��(�~L� ;�dw0�
���i%�T�B�ϻ��8�2Q� �{�y��Q�������X5�{���H6�$�ݹ>G�6:
�">p�*� 	���Q	�\*�Z�V $�}��G�ﻣq�HX��`���{�~�8Ã
*J�߹�I�+����W��L2�VWW��ؚ@����b��8r������}��8<`Q�
Z ����U�!�G_͇�n���"���Ӧoq�����
��{���6�Y�J�C��;��pIX~��l��n�%���
_��j���<Y,��<M����f�ٓn��s�;<X+g����'�f�.�}��½���@�M�T�!Xg���P�'P(��߹ݜ@�J������_�p~�T���\��H[a����C��Z|w��0t�.1�b���q'��ߴq8 VX�Y�^��{Uα��^I������&��%H,)��߷0�°�
��{�Ѵ��VJ�����n���F~����ԜHݲy*��*2�*�+��|2��@�x��HP���;�|
B�B�_�ۻ��A��O�����,��Ϊ���j�nX8{��H�����&�Ts��޷GNC|eq���87��`I��;�?���I�}�{���O�
�@����~�8�2VX�P�o����9����o��ssL���a\����7�}s����+k���%���P,�s�8�XjA}}��5����7��z!��^3�>l�P
��8w-��k_~�e���d����}� d˥[���^<H�'�}w{p�
�RT�����NVJ��FW��oRm4��a��ow�}�~2���&�a��5��me�[;J���6���0cR\�ѩ�}_�c�r孹��	Xk���h�9��)i
���=�w{���@������~���w_oP�Ag�J�;�s�8��G�64��J��s�υ~\���4��'�{<���^�F>5�Z�x:Ý����q���T�����%`Q������H4)�~�}�K�A]�xl?�|>;��_h�I��g�1�p8�{�~�G�����%~���m�I
$�)�j�?c9����C�0�+
�����ĜB�Q�����{z�������[[�s�R	 h#��rGۘ�uU�|5!m�u�h�)i
�Zw��)��R��3��~�8��>��~�l���u�u��i�+R$�>7**U�5挅�<�8o��Th���A��&b�o+X�)�����f�O}�����7�vm�4�u�	'��g�%B����{G�$�)���*`��74��a����jRn!RT+�}��8�2}�Bh�+g�� �@��Ȣ ��	�
���w�R
A��}��ڇC�6�kzdtL|�/+��&��7s[�l2fy�tM�;�x���s�&�=�=*|�~�������7-��s{�����*Aed�o}���B��PIXg߾��m�V�߿w����������8�d���2����(����ů3���;8��+{]�AH{ݻ�>��'�?o�Ѿ�B�B�0+O��op2�*P@���~���Ă�2T+-|�Цmun���r0�dy;����i�ar8�2�_]��@�O�*J�a�w��8�2XʁR�k���s�������Ϗ |%H,����z� ��>�ܟ
6|;��I��m#>��=vl�#�5_/\�|Tw����Vhd��{��6ɤ,IR��~�6Ì*AIA=��8���N�~�����8�(��|����?)� ��l�k�e��˜b�R��0(�<@���U�<w�b�c��g���5�p
Ә�~���*T
�?���C��*�����O��"��'ǳ�"�}�]��:�\�'3yz��*/�!9��Ce�ɘ�{�3�w��+��v72w��b��\_�ٙ��zC
󮵴n�:�{]n��n�;Fa�:+������4�y�sӵ7�>|��~k��7�5��;\�1�IZ���Oj��ϔ6ɳ�K��cb+[�ۏN����SD�����-��*�e5���ۗ�$V��B��Ы��˕W�����.��0�w��q�Ѷ�p���=������\c�}�+���m:�gn���ї�Fq�Վ���8�N0p�x�Ӌ�J�4�X�_�[�[�x��ֶ9���=���Ÿs\��m ��k��a��
��Xg�{���%e@�P,����A`k~�}[~��>5���85�����R������ǐ`V˼�=�\d�8��w)�'���E�>^>�>}o>�����+�{����q�HX��RVϻ��Ì80�,aRT�����Ad����k�;����;/<�]�O��I !�~!#oņ�nvq�Xk��tx�R��~��򐶐�`W�m�����k�c���� T��L��ߵ3�%e*�}�,�`�#�J��m��b|_]��3��c��*JT�
ßs��6��ʁR�Y�����%`V�(���oP.�������{H[a�e��Y� ��~8R�I����@5���F��
�2VVJ�{���ɤ=x�֟~'�pIX]����8Ñ�aF%O�����8VJ2�VW�~���>��b���(Ą�[<��RU�^�ʓ���t��׮�W�s��Aϳg�9��~oӿ�rb����ǅ�X~���P��R
���Ѿ�H-�
����S`�SW��=�\ۭ���2͂w��ڇ�2VQ��P����H,7��Ÿ��ksr:����sA�Ib'���`��NƨA��>�ٗw����ƈ�sx`�L<'�=a�|�k��<O����=����Y���YԦ.e֗�E��)�7:��߀��Y_�h�g+*�S����8�Ĭ������H)��kk���{��]φ�>�NB���1p�^���������@��%ed��}�4@^#Ȁ�G�����K��No��aR
J	���q'
�FT�����P7�?1k��&lnvq�O��=�ӓ}�p5O�3�>G� 	�;���R��_��ޠe6�R�
�>��ڇ�{�~��o�|�FJ� E��"��'���=%��Q�b�2�c
���h64��*K�3��H��>�\	�{�|�Y�G� w�H�%H,
׷�ޠe 3��~�
7��teWQ��`���m,��o\�n�4�͹6�m�Ν���r�D��Q���Hu����N���0�n0{�Q mmd�#�g�+(�_�����B��T��>����g�q_i����G���̓�9��Y(����u&�i��g�F0�.!�Q@����U�l����k2�\b�@��Eo���^B��[�{]��؁YDǿw���pd�����t�}�����h�<���	D(h��3�G�ς-}�!��I%B�Ǿ���JʁQ��d8�S���1PT���������������;�*�����}�� �}���	���<��Z���:;ss^;��o}�w�~0�x�$�H�����X�~���It���?�w��ǌ
M9
>-D1m�>�@꯳�Yk߱����=��q�d�g��!��
$�,����Ì9��*��wF�9L��>��}��&�+%U���Rm6�}���Z�1ɛ��@�����t0(ԅ�k����.�{���d6�W^��I�*T
���چ����,C��;��r$�-��9��ӯ2��y1�ԡ��a&�	�GO��vqݸ�!	\v���]���QW\{v�_���q�ږ�-�=��¯�}��l6��T��V�~����H(J�{�s�8��+|g��u��A]}�jwH4�-��=��jx0+~����q�[�8�Gp8�I����8�R3���ͷ�s�H�}�h�ɴ*J��+
c����q ��
���{��Ĝ�T���}�~��w��ֻ<��w�>���Y�P-�&�CP�� 
��]�W X6��R�?k���)
�[�1O(a.���$� �>���m��%H(X���wG�������b!�%��>�%�\�z\�׾�u{�ɋ�e'�*��o���q��P;�s�6�Ĭ
5�Z��~�:��(�y�L�w��W%o��_)�6\P"c#�<F\��ǽ�V� �hC����M�\��F�뿳2����?�	k���R����|,߁��NB�ĸ��n ׀dQ���{G82T��_��4���}ǧ�ֱ��y�8��V���Ci�#
��}���N!Y++%�������I !|R�ؖhP�@�H�`��1�8�=]Ɏغ!ɹ��+�g���>�(����}�i����7>:��+{_{A�x���-��=�|�!iHV�+�~�Q "�G�M�}�>�F�gL8�Y�J���tq ���~G?8��-q�e�хw�~��l2��Q�g�n0���k�߀�ષ���y*A@����� q+��F���{P6f�R�����<�>�׿wP��o���	0�0R�DX#�v^Ȳ,�VVJ��^��a�J�IX}�Ȟ�yA��+����>� | f��m �N2���{Rm2�g{�W؂�2�qB��(���U�/���{�p��a��
Zw�{F�R��
����nq�Tǿw�C��s;ǻ��o��dY�J��~���O|.^6"�
Q��~>��sA�ID*J!Xc�w�g9������{c_J�Ĩ�u�l�A`q�
���׵d� Ґ���ߵ$@jF���m6�3?hB2*��"�`��N�n��V�͆�\�2�����	���Wbpzq^�no�ࡏ�����	��O�]_Agp^8�:�*N71�2.���[~�G]���jq�S��mf�A���?��KlZ��N�J��,�@�&�%ZuSP'Hx�t�p:�Zg�{EȂxN�8b��,�����F!x��~���Ӆ�z�n��=�W�Ǌ�ؑ�tw�y�����sF!n�ߕ�t�W��?:n�]�r�%?^5#n��9m���{���̺�����s՛A��~���cu|���(o�x�������m t�øm���skܖt��G�ݬ�x��|p����ru�x���}�]����z�ц��[��6Q3uk�ŏ�&yaĤ@��B����pZ�Z'ʽ7,�A{H��vGi�k�f���\ٝ��s��O��3��)��M����}x��96�@�_y���!���]�u��w�ڙ�z�v�t�����vN�P�7o�gV����m�fAA��>��2�U�j{���ױ�j�"�ˀ�N�f����4P���l��5��F��'�^�ڪK�}�A:W���<�k�������I����Q�w"\n���F�:�ش��fl�����05�����U�7�;핵�w_G��J��C+&,��{}�ścdJ�q�)H-�J���أ3&�[c99r��>&͘�~�/y�n�j��,�ږv�|�3�9ZDEH;�kI�{Bl)ww1^�J�"�A ���cTb
���PF,U1EAQ�� �"��"��(�EVE��V0U�"�"""(�"��
1H,PX�""�UEEEAb�
���ETQd`����,�UEF`,H�TDEX*"�* ��
,Q(�E�TU�������+E"�*�*�����X����Q��b���"�E��E*�E��EU�EUb�ETE��X�"�1��1cX-jADE�2�

EQ���dDYb�1V��
�`���X�����V"
(�(��M�oϯ���5���n;i.n�46۬<�����7��|�F���(�9M.v�KO���\�a�ۋ�^v��۱��ٸy���Ύ�����ܸ;]ڛv��f\��ǯ)u���{]�0�j-�%�7�E�����ǌkv8�:�������	Ϸ���p/�p�5��\�s��s��[���vz�=�v��ƺ�ڈ9�x�u	����>WQ��`�y�+�k��[�cn'd��f�{N�m��ΞK���y��Stv�ъ2t���a�q��$�n�k��x��]X�z��A���غla��i=��ݳq�S�8��6��L�{7����'7qBP=�9�Xc{�nh��x��<Jo[a�Q���7'[^͗��x�`��W[=��'���f�G<���g���<�^wg�9zRvOc�8.��{�6o;bqpm���ٌ]3;�nձcs�\�K�Tx��U݀�ǵټ�MvLu������['	;
p�ks�>t��]ݜFz� �5cw���!�v��$�'<HGcɧ{&ȯ5��� �<%g%Ǳ����9���Փ�ە���h�q�b۞Ncp��m[���Ê�uq��`�r����ˮ��<+X�s���Qu�Su�wRv'8s��C���=z��������]�W�IH�I��ˀ��a:�6�^�k���³A��x3��qɜQ���yX���uw2�Rc����cu�T����ɓ�E��;����ă=<��]�
P�� uO"�b�����m��qs��G0Lc����l��q�Y����3'<�t�������%8M��x�Ϟ^��9w�oY����sSP�g1Ƃ�v� -4n�ʜ��8�����Gf��r㋳۞���cOP��f��2����쵍n���
��e5i�/��u�W;����]�Rۮ\�ۮ��.�:�u��-MO*n�GMF��g��[�c9u��A��Q��ZW,��8˻pqv7F�K�<#s�u�]ׇ�C[�z����w���f��|����t˸��:��H�R��N&5mɞ�=���c���F�����	�v�8�;Zۧ4���Nx:,\7�N6�7snՈyuN���k��f#zx���4������^p�ղ(p�V���u�/X�ۃ�p���C�^@]콨��8�:�]G'��.�����n�}�f��@�#*�<���s�:ɵ���8��y2ӗ�f��v�)�Z�K�V^�rOF2��u�;v%��n�.^�۾��ܾ`���n �<#����E� D��2W�q�j�$��=��ja�°ﱣ��>�Ӑ�LD��}�H,����2��ƽ�6�@���6a�33W(���Aa�g��tx�R������������=�i��h������
n VQ1���P�8�YA����x?xӎ׽���ԕ���~LS8��-q�e��
����e ���9߾���H(*�sg���9���9����5���<%`V�,k��^�$�B����jx0+~����a�L'��Y�ݕ�,�_:�u����J�2W����l�B�*Aaf>��nH,8¤�����Ĝ�߫8\�\�y���L��X��x׵&�e��u�n&qqs����Ұ�5�jH)� ���E�f�~�'c�jE�"�xY\k�w���m�@��1�{�C��%eJ��߻�G�o��?g����|�V� ڊ��,��G[ص�lu��] ��.έ�c,��������g+Ձn��w�+�X���e%*J!Xc���g
J�Oo����J��o�߳�:��65��oz��4��l�ǽ�>l �
����6���5�w�O���Vb~7���ƽ�q�~}�yX���3�7�W�:+��=w��{�)���7��܍�3���<��z�ɜe e�8ED�0�"&k�=�<$I��ߵ	*Aa�������Ì*J���h�Ad�+#��./inzM����C :����H�J{8�ȕ����A���HR�=�{$U�!��C���q�����7/|�@�P+(����P�Ag*!���"�G��[�H�#L$
�(�a�»�>��ߞ��]��N�T�!Xg�o���A@�P/�}��8�ħ� Q���+��o�w�}Uװ6��N����a���5<�������3���j]��pI���4q8�R����}�@ͫ���4b�Z<��+��p�AH)8�߽�Gq
�FVJ2����P0��|<�>���5�����Y��qu�$�X$:G�0��OR��)9��x�&�F��c������fI�Q�v��9�}�0(5 �~�}�F�H[HT���7�@�n T�r�����gɜ���8�2T��C����qJ��|r�q��[���8Ñ�{�eπ�=@���T��_ O�K��tg(2�Q*�}��@�VjA{��o4�i���fk���ϡ�뿧�N�|)S��`�����A׀dP$����8�@�������7���B�J�V�z���x�>����gT	.X��t���V}�D��6VV�FR���e�4�X�v��*2-6=s��vޟ��͝��?�B^{�?��aR
��h�ND+%Y++����6�@,�U�-��^a:@B>�WH�gY1���X�H(��{F�)
с_}���h( VTǾ���� �k�s߽����,���M��O�~�x�Ѹ�t�s�� ��>��v��	e����� Y��͡Ă�����^�$��c�nO��>����u5	p0\$�m�,��8��"61d�;<��5܊�24�1��>�?�o���qL�s���8��������e+(�_�����J�Xc�}�P���G�S����d|���G��}�"�9��eH/{�fM��/���f�g�s�\lP7�9�w�<`Q��3�ώ�":vEo��IQ��oWui����jg++%C>�}��y���}��y%aNwo�Wq��ͷ91�q��s!���T*K�1��G#8�FT
%@����4�w&A�#Gp� �B>x��G{�f���-�����8�Wy�z�p�7πdW���}�,����gGn�Ϻ��d����>��c&Щ*V�߷0�0�%��{��p�/��Џ�xl(�q#.M��\�ݷ�*��km'w��2x�e���#��u8�/?��������k� o���6���ܕB����9L%�� {߀�O�VJ����ԛL�Y�?r���d���%a��wAǌ
H(��d��!����]��.�>�:��M�*e��wߵ3���2T*׻�G�JÛǱ�c�����������昺l�k&c�/6����=��z��v�:�0\E��;θzx+g���~���!�K��C)�x���a ���a�{��8�2Q��P({^��H,�:�t�e�5x|�ϧ�SC����>��L6��}�q�S8�	w��={�܋"� #�}�}y���MK�x�����2e
$�Q%a�w����°��IS��h�NVJ2�z���gt;7�;��7_O���@lh�0�8.3���b�Xs}���0(ԅ* d��"��x"<	�ެk�/�Ug���@��L}߿jgJ��P� }?vH���#��U/��Na�I��g���E�e��}p�A�G���(�a�{�jd�e@�P,�_w�� r%`V��c~�?߸g< ��V�υ�>L��%�lbop2����h�Ag̕ ��7�L��~�_��|8���a%a�{��6Ã
��%����I�+%ed�+ﱿjM��p�x}���o8w�L~��8v�a�<ך�G�4w���x��ቨdG���V�q����2"�T��j��_�D����ɥ�,�Bl��~k��[���]��t�xѫp��Jyܷ��[�l�`��k�ۍ{\�J���eP�ap��IؒyrN�k��ٵn{!h'F{q�n];N�4[�m������*v-N�=n^:��n+q�z�$����=s�z��*�v��(��=qۍՅ��JP�n�l�س�����7K7]mԜSv��+>8�Q����n�������v#��P�mfN{X�I-�������B��0<�}~o�Jc�����:�����k��8�Z���{^���!m!Z����߷	���|~�����'9�wP�Ag*���h�Aa��|�a��1Q��-���+�c�h6�)(�I�߻���Q1����o��h�g+*A@�k����D�
5�A������ Ґ���1}�o�|=�1��P����ޣ����78�����Ѵ�����d�����Ci*D����>�\�*�s.��υ����>�>��dRN!Y++%_}��Rm2�N��`�6�Q@��ʹ����#Ou�cR�9�o�7�HZR�
����a ��
ʘ��P�9�����}�v���2̲T(�?~��8�Xp>�\-7\	(f+�υ��"�2�
>I`�IP�1������'߸?�����O�8����Ѵ��Rﱮ�L�)Kg���q����|S�1����_vٹ���qӓ��և#�vv��4��$�sn��9�G��O����?m��iܕ���<�Y���8�Y�J��^���a�*$�/3���8�X}�w{ƾ׵������ID���I�B�Q�������Rn&P?q�]�c���Ɍ������6|�}��n���_l\-{���w܋��u��.h雝�D��s���R��g�lί}��u���b�ڷ�D'+Q�3�,ʉ��!%�ֿsF��JB����ہ��@��3��چ��J�J�Ϸ�胑� g��@�<��F�����27�R���h>a����Xw?��"���y�G� ��9��Wσ���>@��(���o�����^�ܟ7��Cw����j
j�'��߹����νﶛǻ���%e+���ld��*IX{=��Cl8°�*J'���Gc��?}��ϻw�Y4��FW{���6&P/cE���.��N� 
#��e\�f�!K@����7�������w��!\�
��sϷ	�
�YS��jg#%e*�}�!�%a�ݣ�����g~*x�x��N-� mE�i�/\�[�<�r�C�z��[�����w�KF7>��z0�{���l�2��RQ
��{�چ�9R
���ݜ@�����Ƹ���g�R�c{��H)��ם��fπEyL�_2Y�e� �u�T�$�����r VVJ�_|{}��{q�������6ɔ*J����?��p�0�%O{}�$��������.r&T��혧��7g���Vr�8em2c;8��+k��Aǌ
5!K@����%!RX����}�c���?�g��Ά/B��*�:��I��Ӓ�ҏ+��DT�����h���D�:����ڹѹ69�N-4]�O���ζr�D��I��s_�0�� ��g���q�++%B�����8�X/�B�"$8h�W�>�|��~�>�����|��yDD�۾�Dz��|=���3��eH(�~�F��X��������q�q�
Aܰ׿~�ǃ����o[sG8�7�'"O~�����@���YY+�q���&P���������C	+
w�;�Ì8¤�߾Ѵ��Y9_}��RlL�/>�?�GzE`���Cl�D?D&A;�]%]�qѭ[���"ճ����W8=\��������3�۟
��?~��h8
A@������-)
�l��߷	��Q�㌷[g1Ͼ��pd�������6������\��0�TCN�,�X>����G�#۷��O�����y�G�q���X����l�A`q�
��c~���)�g��h]�&���H�&�9+!��ac8�
�I�k�h�r������b��
yGð�̩��Q���~�
°�{]��i8!R%e}���I�0�f�?�S�\���$�~���u�������R�~��ѾR ��Z~�z��T��@#�e��Q�i�?�_��*��M
��&���E<q���f��&/�S��m�jסzO��Xe��y��T�b��BM���W�,�j�{�0<�����g�����?�J�C�����q%ag��_�?��L��cp����>���l0��RT+s��G�G�s��<��<:^ΠpJ�C�?~�g8��F����u�����wP�A}���??h��w��c�~:��{7o=�4�����	�쑳m=&n}FQ��~��ߧ�$1:?����>�����x@��d���{�c&
V���a�aX~�;=w�7�{���?}������Ѵ�!R%_wy���L ^��L��s�s�@ؕ�9�sAǌ
ԇCY�5���������F�)JB��_{y�T؁R��L{�=�q�+(�P�M�|��g@{U2,��y����hC%g��6Ì+�~�4a%�*�=�=��8�FT
���~����}ׯ?c>�����F����P6b�m!m�����8�0+o3�}�sq�aF8� ���vȲ8l�iw`g̕������J��*%ay���Ì8°�¤��{��q&>����G�c�����ȏ[ڙ �X�B
,2J,C��=�O���捝7q�i���w�>�B���� ���ꊤh�ͮ�ۀ�΃4P�)�FtL�qu��%�t:��G7]l�*�Ҍ�y�닞��[J�u�f�[�m��1�:��u�;��  ��'81�e���H�&$��H�t�f�Ji��M3�\����]s�qs�"K+ru�g�����ë<�9�ݛ>S�,�uL����؍���������
�g�7*�뵣�n�/'1��:���r-��ι�sUƄc����t6Y�nݧW�Z����3\�cn�3�'���98�.܇&8�6���!X<��h@'�v�L�6v�:�V��ۈk^��=cfl�n�ܸ�C���"'��C��S/l���n>�?������Ã�n��|IU��(��B�۪������z�ܧ$J쭪�ʹ`� ��)���6�G�T�Of(k+1L�;r�u��A]��D�|���P7��'Of��g1���r�AhD0ˆ�LH5[U"�U��� e�Χ=S�v'� �H������ٞ�I���p�9�v҆���w��bv�h����P$�W=]va�8�){�L��ARʍ$�	�
;rsĀH=��|oc{j"X��WvM	��۪'���� �`�c"k���X-��� �o���]�uu���kj��=X��ulgS��9^��ߝ��B�A)�z##s��V�\׈'��������C��ٿVn�Q8��%אfB��z����s�%�n#P�
���D��5%�J����ir�s�z�2���E���E--c�-�F�.�Ȍ�of��mŇ�V%��m\�������#���@%g�eW�/$~��5�;Uޑ�N{��>�6
� �����H��l���ۛM0��G���Y��m�A�>�!���u65b\��e�m&&�W�ww��k��XN�[��!��>�ͷ�';;1��կ_vԄ�S�U�Kb�'�	��I�m7Y��A9����#�������G{�Xƀ �gS	��fb��뺶�F��`(AH�����Dx�
����y��^�|�u����n����������*f*�'�|�`�:�`�O{ݙ��y���vgb�R�Ss��RDA�z�FM�P�A�K��=9�v�<��wWӪ��vzڐH �η��>���3	�0T�5~�	��)��`�EBD�1.�����Nw�� 	$խ��3WqW�x�$�a��EMo�=�}�������~Ń�N�եӣQD��v�wS�<�_s9��T���iɁ供ޓ�o��Z-�$橵Lƹ��r3iǡ����m�(D^��O�fO�:՜H����m�{�� � N�\P5y��nM���xfK����=�gU]:���������F��Ѻ��9���3ҦYR�����,o��O��t��9��\�v�5Ԥ�����{���W���q�tnws&�b�foq�Y�'NT���x.+�ַި�`ާ�|��'G�4����1v.��b���lձ�;�� ��'��ր6%��0Uĩ;��s�єys�TtL�d^R���������$oQ��NSd�t^�9nEe��F�O�d�����I���#��,{�Q�����|��7�ϡ෨�ʫ@�r��/;�l��������.<'oN���� �'��{̷V,�@tr��R̝�8����}0V;*�.9I�徑矺�︄��t�4���rh�#viz7�<��;��oU@�]�9����(fp�{�)7�V{�'�����t/c	�<h�^����#�]o��ichf�tJoXx��j+�'K��|G���#�Ƒ~�ج󆱝��<M��1�8eۋ:�^8�9w��;�ǧ���;Z������������}��_��Hꪏh�:����9˨�T��Oz�xK�fB�r�g?&�s;۔�y|nҧ���Qw�x���vw������α���*��H��Z*�(��"�QQ�"���,DD�Jʈ�EUb�*(��A*�PF[E�Ub�EF1VR��"�QQb"�V�
��RV��,XE��F��2(�EUUc�Dc��"ł��UU��"* �Q*J���H����e���(�UX��,U�"�"�FEX,D"�ر`�����V(�* ��EX�1��ZUUb�U�A�UEQQ���-�)TE��F0TDX���U������*(�QATbcb���"�T`��U�("�*"�"�E�Q��l��b(�F#�V*�,Q���UX�A<BC\��n�����s�q�S����n�6
Q**bjB�.�*�Ed�õ��#����Wy��$0������B@%_�=���[L~;e�a����k��H\h�0W�e�p�b�]�ff 'vr�����+��OOm��>���H	���0���6�Λ��_�����;�=�ˢ�ɵ���'���olq�r�v]����Q�6>��?]�[�j�*��/2�d@�}�k� �XȂ�g1�yN�ϒ1�Sa��n#����)0�(�Oc'!p�ۈ����V� �S���b Ol�hB)#X��9L�[�I�b
$2T��֗����  ��h w��Zs����� �o�3>�۔��}喡(�B')�=��WDNu�d^� W��ŀ ݖ�� ϩ��R,`&w����س�خ�z|�E�c���<�o��������|I��7A���ޯ���Uwqnj�4M�n��gR�uh�BFep  <
?%}��q~LIH�LT�W���_ �y�@p���XzM����I!_�y��J�_T��df╶1y膢��o\DV�F�yaÆ�!ٝ���\<�t���3�}n�y��0�eUu�PJ;m�5� %�9�Z��o����fbQ�n��mGA��!A.lM%�n��zW��g�f;�����'�-�CHgg6�
˨�[��p{�z���v�S%(B)S�O?S` �{��l��EEdU�a�a���|�1�ni"JB����M���A�K��|�:�D�������K�Vf��� #����
{���Z軸��'j�W�B�(�P#0D')�'��w���sŅ�뮴y��S�=ݷ��kl�	�{�0�ѫĊ��U_v��:o#(:��K��ܯoh��X�y���y�eL�����,r��V�;�9��(���譋�0:�����������88��vzi�%����S�\����jrrbӶ��{r�׮�lLA��,R&��2�۳tQ���S[�q�q������طM��8;�ƠMn��X.�+d��og��4&�S��h�9�=b������\�����e�why�y'�l8�ג�,pkr�N
�JLrg����C�������^6ǫBۛ�=#կ]W]�G]��7]E펧,[\�O��rN�P�cY1�g���A;+ڗM�ݑ�>�����{�L��]_���v��D@������ޟs�n���鰁 ,�k�~3�$Cd1,Uw�wv�	(��.�F=ux��7�����fD`D�,Q��w����x���A�V�ĄT�T�B�oq O{��` �7��[��7�Lmޒh$�ܮ�$�ٝw~I�J8���@���Q;���sȸ�p�7�R�Zn ������۔�)ƦV��FY�6������p�ؒ0(2	paӯ)�ͺ7�J;��#v�vP�1� J2��o��}����uA'm�W�a�76�(oC�b!ܙ��^��^���k�P"9֭t��;�ў���7=�!*tQ0���u��kM��Vw��� '�*�긋�����d
�{s1 6uFN�2�
TIM�;ΛH����_�'��//�R��h\�KP��mȔ"�֭�<��1�uE�	���;Ae��%v�bR�u�P���7�%J"���MҌ��� T�~M� �߽�3"'��[D�w��P�N��Q}'z4gH��bQ�y�mǐ�r��@����g}��'������fb ���l(l�K��H�4@u��wz�b$$�_z�dA�z��p�DY�����o�.�޻�$�Q3p��@���R�RD��w]U����[XJ�1���fg� ��M��.�cl�̎�E�3J���O�mр�-0�ϣ�_GgKm���kw)pv�6.���>��s�{���T������"1We[��w�����2�����I0�	���&۹!*|(�RTĺhgs��-���/G����n]�԰� ][�� B�v6���m���]]Q'���b��A;$ʂ�S��]_���6��݊�4tG=J�X3�/��NL=b(JF��z��[O�B������O^͘}+6V͗+]�]̻�²��Į�y�Ը������ r.��	 As��RD����U�Hn�\�"!�M����wә����Lƚ�A+��$�Kޏ�d��g��?6�נx��V�`�yґ�[,���RA�\�y$���n:8Q��+�/~@%��[�� ]��q]���@)��Go�L]L�"c�m�wo'^\ro/n����
\'n�<h���[�1���
p��@������TA"F�\�4O����PY���,0�V�#� d��};���` qc�������ng�{���Lul�Z���V�AG����*�f�b@|=����-�z��$�1�p��&�S����i6|
��n1 ���W8�G�y�� !n�6��_{73 ��0N�8�L4Ӫ]�N�ڝ�V�/+v�zL�0�	��v��s�0 ��dDN��ƽ�Ku9��X�uL={���wfv�Ѐo!��N2v���\NK\��F.oD�:z��,��*f�u[�����\�o4�j�ǳ=�w&..�ǈI v�Z�߾���{���qi��d*�%6�g��� z�*���dT���˷� _�;3 ���m����s�"6\^�,Kh���k�Ne�i��2t��h��v�� �!R	7 ��0A���l�$��*�����m�"/}�� ��ܷ��Q9md`��[L����V��<��N!��/q����'���p砜��TI(V����$�^\��I܋M�aA���$��D��P��AONmشJK�[�h���~N�]�o�S��  O=����m�$��1�%�����5U��j���&S�]�oy�ŀ��:�*��on<��96{4[�`}��n��$68��a��L8i��rN�{q�tgk�6��� �����A{�m !on;��V��&Zµ�ؤћ���*i�x1/�&9v�a' [�ܸ���ɩ��[����,�1!c5z�V;[h�c�"Vd@ql��r�R�]�M�ڶ��;u��:Cn�YC�冸z�q�3��n{O&l�v[��۷g��;;����x�[�$1��%{lN�[��-�8������>.3Ξ�e��	�qm�u���ַ+��.��rb������`8��t����3t�ݏn����P��/U�.[<l��%���k�ޖ�{v���.�+ s�m���i���d�h"�1u�W��)-��k���HL�J�tL�ɰ�rIi�J!�/;�����a&Ɂ����q� ��U���(��v��>�S��~�� G�r�V�X2)U$��ҷ';�6�����h�<:O+��a �ܷ ���C���a�WY��q�|�*a����&���7�"�cI��'o:��s����m�p���D@���w*3&��|�t��J�%X���pI%V����D>��ae8�.o�վ���D���eE"��	�sl�������ӿe�x�]�p�Y���������EI��t�nv������s V�!�޶��cGA� s���F�]=&-۳!�N��������S中|��:q{q� ���s01�������{�]�7�@���m3�>\Da�I�`M-�������*e2K�DvNL5��NN�긙�O�w7e�����V7ϖ�ݦ�/���R𩰱;����C���"��K�y��x{�����y"F}�3A$S�n�X@���Dǽ|�3}Z���TTʚ�&�`�^]���y��8�tқ�u�\V��U�  B��m� �vnݓe�%Zj�Xtk�^��Y������I�"����{�봒�c���$�׵T�,��@�`��"�2�{�� ������uü%��� >���m ��w[��ïr��ؽh�[hFP��1s��Cm�1��A�C;=�m�[=�Lq���n���%�x�m������bC�$QH����m���x�^�\4��	؉��|']ͤ�I![ݷw�i*�F��К-�4m�l�坯<�Q��� �۹�׹M�ў�+�d�:��I����*ff�Q�k�o��ܫ`| �:��}�Aʥ���c��ܹb�.�ß2{�[=��Z��F?�7=���%�n�^;2`gF�P1�h7'�P����:}!$1���5�m-߽ﷵ�m/�ܦ�U��T*j��M�Z�#cc	6�< Wvsϰ> ��-�@ ���wٹ. @�{��S�eԧߌã^R�A$�uU�|NU�(ŕ��7�m�U���7��P޻��z/Y�S�Ԋa�
�AAC>e�qv疍*펻j�Cq=Ļ�nt��<�/*w�����hR���������ً�>�ʶ ��v���;�u|]{'���π�׹M���|���DS�	�u�C��zze\V7׏0 u�[�
���R+�)r �ȧ���%�JV#a����sAv�:&�I����Cz�����Z��D�ܦ�@oc0���EL�T���F�<Ʃ��.�ef�q댺�")���4����&�B{7n��j}1^��v���K�^ƐlL{P�d�ݭ�3�'s8�K��y���J������;�����>4z�;Ք��ޢT�����s{ߤ����罝�[s��Wbp�m�b�3S$�S�n����S���1^���A|,����+�n�b$�0�'�E�#� �q�R�h@g�.�����޺s�>y�.{^�c�~�~����J�Uq9�|��"�����n����fM�vuΎ͢�]"�2�A [ۍ�����DT�S��}{������]�B�����A��mE��[�zv��g{�'z�#��PB<�DS��'���πAyݯ0>	�'����c�<�Zn��%  2���߀���f �΁�ڪ���J�)�ݎ�\Dz�Y�j��V^��DOv�� ���SWY�Y��߀B̿6�=�EL�T���H�癟, W�հ��M}�/6���` /{�3��6���}�w>�q��z]�C�E{6�ı('�*���t��Y�h��~@w�������oiAN~4o�uu��2�UD<��*�oӆե�ܫ�$~]���J���q�/�˽w����os���U�z���,�k�aE�<!?g"�s˼-�ZS;��,�2q��T��F�i�EL�`�Ҍ�ТfAro��ޗӎ�Y/b��yn�qμ*Vh�b4e�\�{w��=r;L���`Y�{��<X~�:tV_8���Fr��W��G�|�G��$��v̡rK�9YI޷Ǩ��<
���n%��z��{1��%o��>�<ϱ�w��6��.s��4z�)�2�m4浳x���ۜa�7�t]�;�jWSs�r"��zo���(���bp8�|�.�.��zV���g{�G�2�i��|��'�ǧ�l˳b����}��KO1��O��@�==w�+��e�H��w�����%�{���y?��8�lh^��9\��z���`�ߡ�pyb~��,�"[�=�� t��n�2�[R=���^�
��-VދVsbFPN�h��|�9ph�ϲ�T���]�_��X� �����,�Ư�u�h�:�Q�w0��K��Y¯}��]�ܮ��x`.	���Kz�.��<8FX�q��R�l��s9',���5`����/��<n��r=D���_�C��@1��g��C�85�����`z����F���W�s�0{G��I�~η�VO{=�}�����PؖT�U�VD��Kİ˚iY���|LTTPE""��(�"��(��*�#AU�*�
"�b*<����EV��1V(*$

"EU��b��PTcR�H�#`���X*��F$U(�(�E�*��,dU"�b
(
,�T��Y�Ȫ�F) ��QdEUUb*+Q@b�U��1cER*�`�##DUU���E" �`��X�`!iX�
EU"ȱъ�*�,b��1b�`��*�EV("��(,F"
,��b���"�ATPU"�����EUb�U0EE(�Pb
�`,U���QQ��Ŋ"�H�F0Eb*����o��������_�F���V�u�t[�\���7�J��������@��0�u��B�i���ny��9݉:���>��\�v�Gg]���z�������L������[�����ݓ��|�ܮ$睵jݸy.��Ww�ntb:�ݻy��W/mקDv���n�掵r����6��ǣ���vg�ƴI�zɺػ��ݻ|�>��և����h3��W�5�ru;:ܜᠻj�x�<ƞÆ�<g�s���n��i|�\�t9�3���d�&��<wYz:�\�l�՜݅ۥ�aFܼX��[z��IKWL�wk���<n|�L��S�x׬Gl��}���뀶��p����8:�����N㢱ZBܸ��^�v�:��%6Nz��8��g�����㡸�5�u� �Őˍ��&u�+�BD����r�9�V9�Hiy�ͻAc�I��+�C��&v.ˀ�hy����C'��ٮW�Ք�z6�vW8�]��p���MyݺM7\�v�x��n�p���83<=s�fW��"�Η�.n�^�.�v��V��ݻS�����]�+5e�X�7)v�v�\��=��h�l�w�m�]�<c�l�]�mr��N��u�*��;�e�+�\7��8ݷ\�=��\���hQӧ����iwd�Hx��v�N
x6��9ܜ^}��xm���g�is�%���Zf5��z���Q��K�\m�a�5�T�vW�U�1ŝ���콈{j|���'�q�֗��շ�ս��m5㕱N�m^�*�`t6��شV�˻7nĽ���w��&ղ[�����=�4���0e�XG�YZ�nnڙ�pd8u�իw'����k���N�v����<x�=;��K�2;�lq֜R��u���vuݱ�5��F���Vauַcm�&�y��Ȩ���{{,�<fq�r�9�g{V�
���v]v��I7�ۊ���!d)f���ne�؋E����[Ƣ������\�p��ܷFD���8%�sZ�w�ޞ�|�һ�����;mfzlZWU;=�GU��q�
@�v��'f�F�$�wo<�WO1�r9��qv���`�W;�����E;u��N����|Z�������<9k�2��7sO+����G#Y۞{pN�X�Z��q�x�o���Ö3��8m�:���+��"�{oI��[vu0��3Ü���� m�m�KuF��Z�bt��eȱ�t�sh��-�h��h��,ݹxp�q
�1<��97���Ƚn[���"m�b�$.��U/$�W�n�� �W=���/r��]e$)�m�"�v�`E>UU3P��)�+������u�8��5r/ޭ�$�}y۹���i��4��BY�}��v�U��, �B(�)�/ow1` Ϫ�DD=�w���ׯ��Wokq\��C�����yH"��M}��r�vvl�K^^U�i�^}[5�������U��30�h��UU�Қ�%�{�)��ݽi�U��D���0��ت��}�� V�tI&�����)N��u[ټ0Y�)T;��r^��㧷GM�A�f�ͩ.��q��b���ضa��7�ÑLC,�(`���w�w` ��>�h���m�뽁\�0M^e�$�yZ�J7�3A��Q4�B�o>l@���ON��a��\$jh@��tW�;����yYvkuܽl���TV�ov�]��~��5V���W�ם-��v����ϱ[���,�V����Y���L���z}�p�2滫�H5Y�)���&`��Mf�h���_4؀)�d��Gz\<����	^W9$�H���0Qu�$�*$�N�/�����b��DK̫ Q�|�@��ۙåk�r#Q~������$#�AE:`���n""s�^}��P�Itd�p�9�\0Y[����}=���B<�Ebq{R�Br���8�i�Cn�Gc<�n9����չ���1�ڧ��=����ٿ���b��N�yfM��$�K�{�*�	��[ς����Pdx�ͦ� B���L>��P�R�����fg<������ǟ:� ��ݴ���v�b �E����{k��E�H���5TM&�.Ǎ��{ݯ0%��μ�a[�Q']C�a��2eWB}�7��`�2K����˯�r�}`&�9뛚��ۓ;C��	��c�p�ˌS��D�x!s�T)�vn��*)t���E))�L���ϝ�0{�3U�H����^I�ݻ&�Iu�S�f��3���� �����&�BX���R��V��q�}�m��Oֽ鯽y��|�!���۹�� |t����nl��+��"i�M��
���]v��۬=�����R�ZQj�^��ZBw8��L Z.�"o3��I �_v�X �_e�����ɂ���M��kx�?q_{�Bo��Z����7t�3ێ�{�`��x�<�i���v��G���&�k"���fM�u��W���;ݪ*��U)��<��H���V�  �S;�a�������	����b����
�ТڤI5H��i6q�����z��Cv ?_����6�-�� ��ʋ=D7�{�S1uz�o�3ۜ�.wF	����Uwb��qxV
.(�̳��ޭRzZǴ5��j�m{�G���� ��	 �L5��pB�F�}���|����t��N�/�ّ�}��!�,���&��k�o����7q��[]f�ln�y��KG�<�O)�9�TD�"��!:()T�J�[\^^�f :�*� F_s��կmz$�w�}$$�/~�̓L��ʀEEN��z��{!euNfc�n"8׹n���!����e}q�v��R��'=��2P�8!0�N�.ۧT �z�g����#�w�s[��"u�Sh @|.���oyC�����SS$���y�~��#��_�հ Hy��@ ����mg��csFz���R��rLv\��e��lN����+��s!ԦUw;���Y��h+�;p� ����d	 �������G����&�f ���e��wj�Ƭu�1�z�{���Q�)�@d����j��v&����p����C�|qo���7v��s��������e������tsӊ���.��[��,�,J��݈�Fyۃ�������n�#�6����.�)���Z�j���N���8ظ�j瞍�<��=�Z��l�i{eS�Ɖ5��6����]"���[�����pv�����6풞Ŗ�[g�sݶ���u��N&x�\�r$\�$�<��.U����hV�;��q���Gg�Oo ���� �ŋ�v�u�C���AOϿ��?rPK׊��_�� � 65�N�>O{}��>��U�r��{M�� ��z��f:(&�ӥ/�n�=zvr`UJy��� 9���;}��%ƭܬ�]�q%���!�L Z.�%���������W�>�t�����q�ͥd';.�z}>�D���Jj���]��}\��J�-C�n��'����{��'�S|�V��NQSELJ�
�ٝ癟` ׾�a~Oo����s��tWe�@|��n#> �ͦ�F�o�v'�E �B���a�ѳ�5�"�u��:?�;䝻=��MvMnwa[��X���M��$�]Ц�A(��<�@�^m�h�[��<���(�9��h	��f`
��!�UL���q@&�]W�A,��c���鼅Z�ޙ��F��ٹܽ�7]Ԕ�	l��5/!���vf��mM���}Ef!d=�SB�J�
���.�h^��u�-���>Z���8W�: �����`	 �כM���\�T-�Q�N{�k�u�U_LĪt�.��3 ":�� s�q0�9��I[ەZ%�z�^�xJ0��&-N�U�8ˇq[m��� ����F ^m�h�;����5p�v�;*���v���Í8���&!��B�u^I$��j���l�L;��Ɋ%z���ɰ�٭rI���S�M75M��8��BLÄ[��aAnA�6��`������ax�Pݽp�x�W=��s������x��*��fVr=�y����[@ �]�s�\�yWW���:��$�o*�b2�m6(��U1a)LDZ�{^vj���|�	 ��ۆ Gx����Ŏ�:�/%K���lGP��Ijb�%W�S�Ufӈh���n�Y�3��d����+�ʟ�2�M'����]��ݭɃ1v�s>���=�zz������=�N;��s��̭�>}5�zO3�)��'c�� 6k�I=����We*e��~�0�:�{���ܛ�z�'���l�lN�PH���ܻ����;W��6�I)��U�ޒ�"`���^KmgP���1}�Tbp�1|��`��T�ѠI/,�=T�%�ܻ�%:�]ԝ��,�@?'0b�+˘�mnn��ۭ.vGcѧf՗�G��V7N�$P�����BJDR������o��/_΀��f`6(�u3��ǆiӒN��j��k:���M�hw՗v�H�9ں#�S�  g���C{ٹ���\�c�UCv�u��s���Q�d���&�T�H+L��@|��y��޺���sTW��r�;�������n]��WAQA���a�tk�&��G+C���z��֙���m�Qӝ���yֹaN�]r-��ۜHc�X��O����c9F��	"D^<�����Ѧ$Gv���%�*���3����y�����,�}9�G[uI�,0�o�"��=Y�v�H�u�k�FA��{�Q���������#���y*��A5��8p�ZN.>�=���/<]�B����dT�+�#���(�T����W�E[\�ݺ�a9��� �ֲ�U�bN�f�nNzQ&/�j��ק8IBaˈt{T��%u�vY�;r�Y�ݩI ��o^��D�w5���T&�����Kz���M7	
�g�d�	�Nv/sD ��˙K����v�D
}���H:�u�!��IPa���6*�H=��=sy-t�_<�@�^W1���]���?_���o8�����I��9߂I����J��"�'�R"m�M��t���Y1�w�v^I,���M$Gd����#v����t�:b�DC���,<��S���V���2�v|r��vi�N�ƚ�3��<��0�U�E^�B��G(u�&x�6��|�qXqvU�^[]���Ӈp�Λ�v�t�&v.�;1����D���S=��m�Pٹ��:����*�{'7tp��-Y:�������v�{['�ˍ�����Ņ_g���m�n��v�:�X:��e�z�kJh�^p
�]���<ul�eݸ��n;s�lR�����ũ[6�BpmÑ�.���:\=���svvZ�U���/J],���{U���"!��
80�o�"��)����Aד��� ;���{ٓ�ً�W˔�=$����?�/̇�-���/�"�T�$:�
�wf��iǙӺ�  ^W1����qDd�~�ܲ'����7T8IBh�ˈu@.ً����[�����{��d?8oN� ��M�𳯝����d�*����HQ�����l�����9�n�����l"9۹��M�ǚ�#Q�k��z,�TUA5���� ';u��j27N�!��5{n"�|�!����E{lQ�fo2�>�R.Ӽ>*fַ&���vzX:,�ttk�On��zB�a(�`�X8j�Ȓ��Ä��NoW� F�7b �;w3���Nq����̧e��o��du�XD㈙i��@P�EyOV�Ѵ���ș9KM�3v�G�ҵx>Dv�y����f�%��Zb�x-Ӓߴ`�X�&�I���4���,��6��3�lYORB��Ní�{]�5}V��G=�`��[� \jRr�d���e���s�%{��0�8���t�8�擰"=]���yn6�:G,�����$J
�V�zQA.y�Ua$3X�M�JD6\C�]�[;��)p��Tk:Y$з��v$��\�tWgOFżGBIA}�^���q��&ɪQU0Ci9�3 �9nF�~��}3s�Zpd=ۨ����� #��[J�sw;��f��p�p���M2������ȍģ���x�8�Ƚn,~o�9UB%EUT>��n���׋ �]����F�����.�������U��B��4�E�0]�{Q�Ԁ];l�;��=�H��N�Wn�D`k�nH>���?@WE^�8c(��(�&�P[5�wix$OsS�'	8Of\=���:y^���_L�Ӗ���o8ߥm�`�[�Jd�֍*6�慌i�˽�i���Șn�����xoz����A���(�o=���"��ʴ5T��Y3��"Ӛ*w,/�*�<��޲��gSF��i��ä��]1jḝ��Z�֤���l�msB������ҽ��� G}��ۑ[��������R��%A�[
�uh��f�f'"�B�M�U����\X�~tl��s��n���Uץ����N�n���&u��{7������!�X'z*iO��LB���?h�/�t��ZD]w�v���;L��{��Wb�j��pBz��U%W�c7V��t>���[*��~0���<�W̀�;�����)��9z��V�ɼ)��r~����5��s�{/<&i]X��S���Ǿ����r�s�t�X7��i{ӄ}�^3=��7� %�aB̙���ӿH��Ц�Ľ�{q��V��;�h�}��^��^du~۹��^	�.<�U��|�)�&�2�"7���w�k�[����5�����f�V/���Dk��zPn��5� ����9I���z�2�o�q���znm��s�H�.V�UHܶn#M��6"�����r['bl8B;�F��^���ۮQ��󅋉FU��^ �����~���N4W��7@1-
�g��]y�D��ٞ���/Lg@ˆ���2O<u�����՝�[%��u��g��ǋNI�!0w�f��ܔ�[�:�ۭ���3�^�@ٰ`Z�ml�]��p�L�+/$�X�{ �e�gxk����ݿh��J0UPU�T�#��� ����X0F+1(1X�b���(�*��TQ`�Tb#+AUTF"��`�,`�,��EPR,UQ�A���P��UR*���+"��F(���*�`�QV(� ���R�J�EDTTQUdX�֬T0�����F
(��DD�AD�YZ2*�-��UV
[�D���������(�kF��m���
�Ҋ�Q�QF��@e���("+)�� �cU" �*ZTQ����TPDQe�J��jZPPPDEAD�*2ڪ���TQE���jJ�(�V�+bŊ1D`�QkUQQ��A���kH�U��(�-V0�X�J�QEDDm%T��ETkjX�j�F��YY+"�$#^�'��g{n�$J]�U�W�#�(-'�%G��^N�����Է[x�b� =α� �����ʄ�{�q�{�n�>��N���U5l��m� �cw�SJ%d{�'����� ���H>����g���O�P}0;�_Bp�~a�0!�g���֞���ۗ��N�a��	�۳q�������z3X���5�u։':��"RJ�nS�U����{��Wg�0�F�d5y�QT!��-��4N�U~�Ifr���6swv��XD7�� �>FGo�D4K�*5�r��G�����ь
�8Nh*�&*ᢷ'ͩ�H=޺h"&olT�{rvkr#~�q�""2;�n�*<	<X���j:Yg?zc"m^1w�]n� vt���w�4�۹h�Ɋ��t���&M���%7�.Y�z;ڷ����WM�Ƿ��=�F�i��`�k��uoN�Tϛ�=�"�fƓ�-�����q�"6
�'�7��q W���ܸ���ʸ/~v{���"#��� �����&<tǶ���/�Տ%�A�Yz�
c6��v� �]�/����8�j"!z	 �x;Sb�Xe��ם8���]4�@*�n�b��Jsi��-[��~ 6=�mX��$MhҳQ�A�6~vL��5C(����}�{���Ow�0>�۹�z���{��{I!9�QT!��-��5H��˧�+��� ���}'}�q8I���ۦI4�7n�$רtH��C��1;�b�OHW\eٹ)�ךw)���� ^�=�~U}V�]��ThD�ͷ���Ƥ��3_QJ�2����` ]�l��C�t>��N�K��	!��dߒ<�ܓ��z�b+�R�m����Ҭ�3��n���7���To�>�� ��������?5�ީ�\���7�VW�I˜�/�{�<�T��7[��j�u�i#l����Q�sq��CK�-����v��qڇ��v�ɖ^�[��닥1;�=�3�;2&۳�s�z�&�b�u�8�W���l��
w�9�����x��WR���]�<`����)n�c
�]M���؂��L�ׂ�8�gp8d�'���ݧi޶���{u�2s��a�)�ֳv�#ՉuT�:;=�p�3uȕ�Zk��J[��q�v3[��.�匉�\�jn��<%�j�Ͽ͹w~��Oբ�=����>�H :�-�A�'�����]4G[� +���&|I��qC�"�,��T�&�PI%�%�>������F�>��3> u>��� U�x�ە�ˇ��K�78��n��3��� ��l	Ƀ3�nwk$�ݝvM�$���&��U~pK`��RZf�$.�l��s�J�w�`$ ��n�������{9 c�������C��f�IW���� A����0��Y"�� >����A��o��d_s�~w�5^�At;���v�Ý+�tp]3='S��rԽ�C\��nì�TX�`�	GwxB�D�[5rv�����V�DD_s��aN��x�9͝�ۻ	$�Ǹ꼒��	�# ��EL�h{��9L���}K}U;��ys-ڞ7>���U� ί���"a7�hY�2���.�En��@hNb�p��}�t��~�����L�5�4��<���[uu��`|@.��q�2+�Y4�O,�u�^���c�����́4LE*�����w�� ����� �_ �g���|� �H�ͦ����UJK�8��[n[j��˻��۲��}��� ��` �K
�u�	����f�O)�� ��i���8+��f?8%�[fs�q���^	o�^,$������<m�q����@�]����߭C�K#�ﲼ�OU�,v�i͎�iގNw3�/E�����q��Z��q��Q{ֹ���N���s�$�I���Q$�-�m��!\�w�P֞���$PH�}�^��aو�@��)���6���^�S���sS�����IGV부+����du���(wi��]&�@	�PK7u.�N9��)ϳ������ ���`�1b�JjhC��؝@�j��S�wv���n=�\�t[ ��lS��� *M��_Ayz=�2���ZsJ!Ti��$���2o���@!uw6����bӻ�!��,��FK��ɵY�؛�� ,筸����7���n� �XP�*�������{��A)���3h.̻��I,��$�9��P`���h$��u��"R�u^HFnRx�t�͒�R��a���-'����5��n7ch��=�|y-�۬����~��.���6������$M�Ϊ$�H��I[s�nd�#����` 箤�%�{�w� �Y�'*>�iPS�W����Hϭ�ڍʤ,|�� �����_SaAt<[�G�Mz��ؘDעb(�[�[���h��d�I ���=O�
�^�u������ w���I��h��bH,�I=y�㟿D���̃��,�	<��M��d�Ѡ�����嵥�������#�ݷ��۩�HU	���ͦ�Y�������[����bC�I���J֙��۬���LC5=�" ��o����R� ��)ãђ�I���9���b캬�V����z��A�|z+�=}��w�q5:�������wQ�·�n����m����z.�qø�۳�	����N�����ų*%Q@T����g��3� {���  >�}Κ���չ��ݿ��ݙi$�Y�N��x�l�&-�T�Ӹ�O��2���Voy�����n zs���ZP'�t�gs�м�"*��$��yq2A"l��Ѐ�m����~���N"a��B^(��Da��r�L�m�1��ﯽqk$��\C�x��M �&���'=vn^�nɼ���Okd���3)�%J����;��`^w<X�4��D�vf[�� �6���^��$'�q��r����p�
����kq�#0�Ԇ�b/Ն+j���Y�nr܁�Z[^͚+�%��~��I�n}`Giu��+����jf�d�Z:�ͱ�b9㷴�l2;
�{�.v��ll�<g�S�۴�n�6]�����az.0]\e[��B��oV��z3�<���Qr\�[���u�[e��-�qgz��c�j�c�f�Elrv��؍Z�1�v��V��z}��#�����|����f�3��s퉃�׷���#;��ض2��V��ʜQ�$���Ԗ��f�:ۤ�H۷�;gg1��cj�n�c!m�A゠���������)Ó�㟀Iy"x��
�|�;s0>��
���l �n��{�e@��
L�h�~�ϰ`��{[RL�ި��ޫ��i��� ^v�`']����;����dF��3p��ӂa��5A.7wU$����� u�~�q���[���7d睹�Q�'*TW��z:D�\��*�&��ԗ���ڢI=�ɋ��s]s��	;U5(9�
�UB��Ƌ����@|׵l+19���{@\^7L"���f Gm�]$���ҭP�1�9i��D(N!�7��9c���t�՜������ݻ�#���v�~}�������T�*gg��i�@��� �{n",�US.����d1�sx�V�l���e�漺r�PIy'٫ץ�T�щw2�^\m��W1z6��y��ۚ'��w�m���u+���e��f�1g�D�''OW2�nt(vʛ����bc]p���������Zm:�3�Q��1 ��I"ڈ3Aw]e߭Nmk�I$Ky��vJ���|�@s�����{M��E�&�QPL0[f���۸��3���I'3yY��	�ͷz7�s.�}K���2-֐���]Q,�"&	$�b�8w���xH{�x��gGx2O����|�wf�a�|z7�ڳ:��z��Q�k�h�M5@�ZRa=�j˸u�;^�Q���ݮs�s�ܡ��W��U{uյ�ӑw�ٟ` �6�� ��{͒�Uy��f-^���ͻ��Ao^�`}�<y�(TT˖�8�杈'�zHq9ѕ���}��@}��n� >G�{�� (�����]>�0u�p��ؚ�$��%A3N;���� :7n�I&EP���8�kq�r����T����Y2��f�'"�n\f�;u��V=����5��ø侀i�{����Y�j1�]��s�����@ ~�T)$��h��T���)�����y웓���g��QWrA~}V���΢c��2�oח]������;5�J���� -������� �����7�h!z}��ݷ�ѷͫ ���ݙ�.fۉ;������B�Ԣ&�m��.uc����`���n�62�I^J0H���DlIM��x'w��G�����>�?{�0+ޙޥ�#wM��8�^I-==LщȈ�6K�7J��g]�$I���OQ����$�@{t�y�ݙ�	����]�[�#� �@JUD�i��]D0��sϰ> �Z�V��f��]]�'ĒI��y� 
����m^��AA3Vήt��+=�}=^��g�Go]4 ���0;����j�ߊ
�����YU'�2N��>-�W}��{7���@rkK*菇<��ݻ
v�y����W��n��3�B��ˁ�r%�f$��:kzhJAm��
�� ���l���b�H ���m+v�Ε�]N��e��a$�םwi�fs�#�D�T��K%�T8e\�P���b"v��Z�r�n\�c���Jr�[���=�a�i�a�������I{y�0 @w���!��E�fe�z�"c���I!�y�d���IM��q<���gh.FO�.]� �����$I��rI��m�[{��m��=5,�ODDP!�Xa��yWVmݤ��]��@y�� �r���\�.{s	�_7a$Hٚ��"sV�J��������=Q[�n��"9������ ��ݢ���v.�'˂L��yvO\m �1�FQt.}N� cu�q�p��y��o7����H�$���g�!�͂��ίx�	�{��<�<_L�؆�.�"}��vO}/sb����f����Rʄn�TY�Y��Y��'rs#4�I=��g���ŏ�a^��t�<���F&<�١���^wv�Nu�)��+�QW@�V��G��1�0��5�����"��=�X}ܷZ���@�x�{Wf�~�\����{K�ǣ��n>��Z/�B����Ty�;��9K��	��9ڑ�t��
�6hnƳ�]j�2�kl���?v��d��p�t�`��}�W�S��9�G���ڒ�=<�2mD9�	����9�Df=H�������6I���7��T޲�������֏���O.���y��ի��7��d�i��zi������/7ˡ#jkJyD��2nM�%�$͚��ِ�{�����C욲K�.OIX燧YT�[�X��ٴ,��Tc��!=�Mm����v΢�tMw����6K�#��'z6�BQ����ʟ����������o+G���u�Bc�g�k�I�}a�{b�Q�\��Y��$+(��ݺ�j_h������p���t���G_ωzW5���ѩ`����J���={�W�u}ޫؖ�{M��ϵ/j�g����Iޢo��ɉ:��}AYυR4����ޭޜ�K|$g=z���T�M#���mCrD�����Tl�"��b����/o����P�)d�����S�s�z�ʪ˩�G�������DG���ѧ|L��E��+��ߝ}6%E"�B�6��Ѷ"(��(��,V-����Dee���,�VU��lR����J��*���KYm*�QD��EiT*j��d�V�TQJ��Eb5�V�KeAQ�P��ET+UDDj[E*DAjE"��)�VQ*,�(��iiam������l�Zѕ��ImP���,���R֑U�B�%�j���K5�d�U�m�Y"Z�m������XV
��Ķ�V���(���iB�d�ҕ�m%�F�XVQmUjV*ʒ�TVJ�ZT�1�Y*Q"Ŷ�
�+�-�,[J-h#(�-�)FőAe�(�%V�#�R(+m��V*�-ʬ�lE�Y����Qh�����RZU�(�J@�
@^7��i�q8	x��z��&���Gu��g�:�����$��v�m���\cNE�����:wN�]�oE�6;\t]E�}�/!����uĎz��ۃx�=�����#�=��n��Z�vy.q�1Wn:Hi:r�,�0�������vw�g[Ep�ΰ`���8pZ�p-:+�U��략rs�n����np;b�96��m�uF}���3�Ʊ�q�h2�ɸ:���R���x;]�l�񹣱���<dvyw�2s�k�d�E���aى��m,gf����.�ω�cg�n��v��8:�d:�s�g��m���rl����S���r��ڹ�;��Tuf�#�"��㱨}v�.����s���]v���^\��`0k�Nֹ퓍�<�7"�+�ⶶ��]�2� ��cu�:��;.����WA��L���;n��u�]���5n^7�]��=ˍ�<c����v�`��������zg�Q^:w@��ܼ�,b7<p���"���u�s����u��܍���fn:3�t�n(�ɧ�4�3�Sm���D6ù�Ӻ��^;u���:
�5�y6�nͷm���F���z�{�����*���ݲt���E��z�x�;ed���,��������Mv�J�N3��ܛ<�ݩ���>����=��;m��r�,���7@�^�o>�q�������Ǫ��mn��k���q����<S��)�ۃ��Ά�Hsnt��msn�ѻZ�w='�u�ӓ�+��j�!��cf��q�ix�egl��-5]\��uӋf�Xꝺl���|+��@m���ټ����w8Z����T��m�Z9Wp@D[��Į{<�Y���g=$=��<���N��^'�sc%��a��&ƒ�&tN��Y�<s���Z�,�p� ��t��ylGL�>a׾\�h��z��v�E��vݑ{n6���ۤ��0.���h{��ݢ83�xúi����:_`���K��l�s��E6�0�l<��`ŗyxY�ݎ�8�n�g�����:Y��;��2�ޭ��	���F�-]����v��V9�v�w�����Z�j�;ۮ��p�q��n駄���m�\�[)#���/97L&l�{9���n��n{8��q.�5���»{����9�6��۳װ���#n�����-�]s�vI��ѥm/���<���o��V2۵o4��Gл��7��v��.��E ��a�&����%�Sj!_�9�b�	�|�$���IM�#�j]��]�BNO�?k⿄h-ŧH��T�lfe�E��Y._?n�XD .�����m�dDs�z绮�[2��k<�GѾ��1
�	����o��F�i��fY�XUe�g�����G�����Vzdj&(�T�	�3��绔�Dg�r�@���� DOku��7sn(������V�Z-<��@J"*�r�8���7�u�������ܫ��	z;]� ��ݪ���հ��L�Y����/2�:�9��b]2wU�9��Ň����sb��eG��۳������SSB&����ey� �� ����[����az�l�Sh @#cy�`��tD�
�)*�%�����0J�ˮ��6��w{�~�TDt����2��7V�1;N`��E�I�|��b	>\���֍ؘ�O	��c��N�F��T'��x����� v��f ��{3޺k�s������v�-�i�[��uIq��u䗒�f�ϰ��K�l���VƠ E�ڪ�	/�ݻ&�^<0�B^�`�~�~Ź��=U�D{c����@$���� �6�g�%C�^U�s�����Qva#Q4*U��c���G^u[�5��F����S��y �x�!�nn�� �כM��q���>�Q���Z����C�3d2�j����9+�7mQpM��+�m�.^g]�����_�@D�UA2k3�RJKz�jť��+���0���S�W^�:;�ݐ �����*ק�a8h(p��.q$��>{
�`�I�yy�d�k��	���s�D�I���(�g�ᢊ����� H=Y�l���q��u��9
�wv���TV�Є���98PRٗ��hYp���{m�d�im:v��_l3�g�d�������̚c��R,r�;�c.�+-��D��mU��<�\�J3�L&�-0�s^KM]���r�b�t�[�"7u�Ł� ufۆ ��7�饝E�ِ��ew�����<��B��$�h�������SW��$��6�$��9�d�I ���� �_7c���/�{�&����v�4:S<v�Y-:�s���B�A�i܃��n�3�$�`���ݭP�i&e7��Nc�"��:��@E{�����*�m\E���I>$�'�����NO*S�@W¥C8�杁ї�t:�<lKݼ��%t��i#e��J($36�I�7�3o��B��n*(�o��7�DDlW��f����{��	󩰃��]���N�����*�%�����{/)v=�먴 o{�q"�t����j�Ҏw'�F?e�cڽ֮{���){��{8A��n{��@���1��9����#e'TuN��r�ʼ��v	��'����6��I�5PXf$�6ꃡ�4�@ �o����S}���<�����sn�����1ޭr��������(���0x̯&{^�v��;I�����Ƌ��GB�OϽ�f���7Z3���O}N!��N��@.��s"&��z7q� ����l""7Nv���	rL4�2��z���֐K$�=�&��~�~��> 3ƻ�� ]���π�0s2���6h�ky�6v1�$�Q�c�k�Ѐ�7��y� ��G��}��` q�� � �wۙ�S�H�P�fP�D:��4�y�r"�˿pT^��" ^���b vfӉ��.Ģ�,�w���.��i��5Q-�>��b�@�m[Q�ܫ�����6���@)��9h������O7'EV.S�w��ɸ����˹�S�wr~y�H���\蔊Tr�G�'g�˫���q^���[���'�����ꡦV�q�XL���i0���l��۹7W�v:��V�v���s��ƍ��ԑ��lV9�x��������qX���{[�v��YWgY}��w\���\a��H�ۇQ��d#��R��㭵���hx; �\V��C�=���0��.S@��9M�8ɞ/nr
��V۱�/k+�d;X���l�W%�8���M���=�t�����vyݙ���:6�	�G*��f}���僌�>|�X�ʝf�[[������_�l����-�WB�I%�ٵv |���a�{5z^[��^���b(�\F&I*$N��?O4h$�p�9�mdd'�{�$J��ۻIy$VGR$�_;t�LF�8���E0�	�4f��	Ց�P �������c�Y�}��ndF �~�����ژ$� )P9h�{"VN��25vt�C�v<�@ 5����z�_U�P������p=���{=$�T�jfj&f��v����۝'!��{|��7}�� �y:�Љ&�c��v�]��ꞁ�
!6IO�I�%����r\�F�%�M�A�Km�6%7Aq�-h �wO"T� ҩȷy��U�I$�K��y-a�zܮ�8_�{�3 y��Ojnh�MP��U�;3N�H�������%��/Qb��%,�E���_}�<���^�ݻH���l�;a��J�E�αFFˊ���=sEվ��v�ף�	$�<�p�e{������y	�	3j���߉#�x��Hh:�q�î���"#սM�1U�뗇;��ھu^H��������\"�-����ۺ�L�����;a"gs��D��=�A"W�6��^�{:bf�K���.�N!�OHI>���"�-�u6 ��n<����w����E���p����]RE��6�왰ɺ�����v��Եa�Rj���U�ڹ4�����u뢼��.cѝ��@_���,�W�/��VU� �{O�"�׹���l�9�J
s�h$PI�:�[q��l��'B��ˢL��Cud��w� �3o��@ >�k��@��-0��=Y\��J;E*d��H�sT���l ��y��DOޏD���*ԗ�t5�˫�ww��O�������a�mO�,+ͤo�nx�w\�Q��&�,��|�$~y;����Z꼑%vmm݄�2x�0*,����L��$9�@��Q�!%亲�z��ݚ�F��}M[��{g}o'�|���^��r�"��`(a���K��nł�}���Ԧ�S1�dC��v���^H�n9��.9�u37�&a98�t�JB&����I�]J���o�wX^:ܼ�)J;���&	j���6�	A���0 .{�p§�+j�`m\�Ԑ ���� {I�52R���U2S�ܺ�|�7�]����&n�G�籸���M���An��ؙ��v��1ɧzx�T�U��U6���� y�մ� A>=�g�'��nm�>�wf�bA�j�{T7Q
fhA7T[u{t��30��#�sw�c�>�6�43�[�u��'8�MnJ�G!<Ed�fZ!��)q�6���5��,��PMm�����;��f��
�4ؘ'׮����-7\[��0?a.��p��I<.jp�B�I�s�i"s�*�y"�e��|���M� |��ܕuT_������Ϳ�G.ދ����.oe�C�μs�v"�n;^A1q�&�+ߟ_����Y�8�c��gc��y�o�����ߝ�=S�����_{3 @y��@<�A0z��X>�֜�B���\��7��~K �Z�����ے -�{�o��{�ڐ^Ӎ����QS*�Jl�S�a��v4�<���;�=��[3������ڶgl�r	zsdJ��&�Kc��dl	ά���h��V�"���D����,�3��E�NgSh9��B�jD���̜nD�۹�0�To��G9 .���a�Ȇ�������	����<�BYsy'�ܭ�ۻ�{��r]{u�x�L��o���k`?}-����ߌθu�9b�����/��h�E�K-@�[.	�.�7�w�\���d�۬;{.��Gt�]벼J�#ə��k��lwd�v��TB�fr��1A	����]!����mp�v�	�6�.�]�6j�V�����^m/];���؞{ ���1�y��X��ϯ0��Dc!۫\�ƶ���=dm�g9��|c��A��m�6�wA7�ֹn�n��u�\��ͯ6�N�/'v,��[Wn$\���cP��l�X#� ����m{qv���:�J��2]~�����@����v���AEK��nz�'v&�vh~�M�{�i�8�2e�ED�iP���ۗ�~��J1ޜ�-D�%����Hz��"v����C�y0�����3��PU��0�4�	����B�H%�յ~�J	s�1��	��L+�< �띲!����+�q�53SAR������7/!\��B�� 76rƒK�.ͭ���)u�:�5�Y�ӸXIױ�B+����$��AT�e߰�{3��72p�3=jL� ���0 ��^�b��Ϋ��b�us�	��O����@��.�秘� L�N3^ͅb.���!12�4"�{�N��P�H*��e����n�y����3��x�eEV���� ~���|I�g�$�UPK�"3��	nwN��}#�%nWj�w"���f@����m6b��u����s�9T�JQ�3*\�rD�\=�	�uk��r���E'%�wʩ�e�2�!����s��[ς �쟵�@���?VZ����*��t�q��.b*%J�U8h��nb�@gy��'���d8��F`�q2�$�B�kn�$I��sI/U�* !��L8iT���l^��Yt�#޼����`$f��?� Fs�{nkˢ�}� ��y�H�k�h���
�UE6v��a�s�������ϱ�f|�He�:��(+ꍤm�׮jQ�$��vN���݂JP��$I�����랧!]r�݂�a�&op� �a&IP�S��~�|�fu[ ��ZƁ�n�l��{�7[��כM�Sژ�!� �
�m�nD���a�<�m�{�� �כnA#+�[� {%��/0��s�%'�JT, �D)t�f�$�t����I&}��!5�G��jP�)�ZB��f�VH�zΗ�V�A�D�x���\
T��ǝ��E�Y`��͋�c��4U�Bh����8���!AsE=�XT֫���v�-�Q�鲢��d�g{�N<���ND����s�'�W �����.�����P��Kݨ�0�s�Ux�^���`�<��U�kf���Nȝu���v%'�w5��u!4�L-��bv]�#.�24)�@�b�p9P%�y���+�w=H\o��Bu��9��Q7qX�OǄ{������t�2�k����7q���MW#'+��3�w�;��.��w�磥�Lx`��Hn�zc���+���k�tNzp�Sbd7�;��}����gPRz����	�{�絹@�w{d�]˭Ou@ҩ��vS��hA�eť��4��Ηǵ�M+��wR����[,������!}��[�}�e��Y!�9��f�F�+%9��E�:����T�ۢ��V^җ�e�n��t3�x�.��2�n��t|΂@�� ��nf���sB���0{�׾�^z5|;|z�T4���;ө������]88p��Z�?7�Z�����q�}�4�|�7�����K�Y�.��ƭZ��;��B��m호�3��z�nг�t^�Y��%y�mک�뫄^��q��,� sM�.k���;��8���r5�o"5>��Y�V�8����}ѻ�D^>�ͣ�:��*�֧�Yh��x�R��s�A~:��o?X����	9�VQ�V
V,�щmE���l�lP��V�JȢ�X[j[J[U���Dm�
���k(�b6�0��m�ikVT�
Q���h��������6����eeF�Ab�iZ�i[V��l���J��F5����ib��DDAJ"�Q,TFEF��"���BڡZ�A���UVJ���"#��kh�T�m�R��Bҕ�aE�������J�-eb5
�V"ZQJ�%�U����e-�-(�)�Ҕ�B�ZQmTA�6��jV�����[mJ�m�Z+QE��kb���j ,E`����Pm��-������j��R�cd�U�Z#Z*6���J�[A�� [b)l�F������D�QQebK-+-��%-�H�UB��DJ6�+[hX�%�k+h�T�J�j�ʬ��A۟7�"#�:��D	Gkj�&�%�B�JU(�p������N��$�T�ג$��q�QA"P��۾����7J���uA*�$�M��y����z�a�[���up�@|e�bw��f �A�2d�������n�պ���\�n�ܫmcu���
R:SS�LRۃ����}۳��������H7D�W���$�<�mS$�ͭ�������u��{���:q�Gkt��0��%C
*���ˣ`%}P7'|y��1��W��@}�=�XDw��x e<��98��~@)�Lu����
�l:�Ɲ �k׋�������yj�t��b@u�舃��s1 ���F2�BT�:�t󱺎��@��{�:� �׹� <�yn�1ł�y��
�����d�l���U�y�#=��o6{?H�
�ǻ:�o86��.N�C�3��]�R���R����]G \n��"h6Z*̔���ym��شJ�]W�I�
�
7G�x�o]4 ��3	 ���l��U@��k��(a�e�/�	4�G%v8�v�B��F�C�rug���n$Fٻ����+۸��&�H���ݭ؂#{^�X"��A.������6� ��ʯJ$�;g���@V\��&%&ᨪ\�P@|f�WTe�(��릀�m��`I$��uC�S�y;���Nf�ٳұ_���*14v^]�I,��m �A^�F8��^�g�;o��� �}M��Յ�B
��f
��i����{����� 3_y��%���1l��z���f��{#�\�{Uݓ`<���(�a���J�'����$�����)�{Ya���{/.�%��ˮsH" B��m&x�)N�Т+�h�w�]�
�Fc2��q^~>��/c��ˏ~V�#�4Ե�;��w]���#��n��W�s����a�|B^(�5�;B��_\���μ7���b.�{*A�m��8kq��]��vLO3�:.�]��l��ك��3�qx�v�9�m�\�ɍv9�h��;nk�ۖ�헵XW2W;�:���; [`���u�|��Ap��g�-in����x��^a�D�AnŲe���;=������ox.ۆ�5�mW3ۖy/kF�[����Ύ��rݷlm�Ӈ��:�Z9��[�:�c�.��{u�p�t˜q�U�Y	�Ç�j�2�Z% �]s�  FWk���^vϓQ���3_f~I�z�܅
	����HM�]��WJ�I���{��|�{3m�@,�۸��i��3髚���y��|�4!0�)4ي���:&�D�y�$��ϔ������� �ٴ� Wki�̯�LUHE(&�Kh|��cw>�s�&����F����ٟO�kwo���4HsёL��p�eT�S�Z�ϛ{^���A�ք��~� ���!����a!nT���QB'[��	��%����u�
7��j+٧0�n;��x�]�Y�)�������QH&�\���7�  ^��؂ ]׻���ˬ�pm�䷈ܲ�:mD��o�5�D��)UK�v^�0����.u�� ��V�W��黽/:w�[�ܱ^{���ȳb���/�{}gY����"d��F���� b���%k��S�WW� �@(��v� ;�u�@ �{p��΋�ۭ��H�SE}U$9h��lA�{��פ)��^�� [[�B�^	/�ݻ&g�Є�$�f'~'������Q�v�'��l@|���b�ϩ��F�'��N]D���*�-�{|�l�L���˱h �U�ޓ�*x���2y�D/U�߾ ���3��:�A�M{����wٝ��C���X�����u��<2��x�@_�w��E:�qmnwn��������+���/6�&ς#}�^a }�W/r#������<�����3
�Qs$ǕU*��A����S�`c�9f��Y�0\̒N��n�&����i#j�w2�PQ�}���e$2�(("!�sJ�\�ns�q�ٝV������woZ��ػ����_^9x8��c�0F{;��_�o�
S(;�zx���CW�=c�����~�������	򰅻�_D�^Au�dF�=�>۶ o��x�@���}JfT�?D�IX+���n�:��D׀�n7 vgU�CY]���*��Ѻ�db�s٘N��M�M6b�.{�����Z^mz�P��˵G��DK���� �:�A �y�1aYe�n���)�ḁX��䈆�L<y�5m�'`��=��._M̻�leY�{�bd�0�����<�	e�90�
�t®i{��q>��	~�� �ˮu^Is�t�!6Ȉ���KM���C��\�G��Q)o���I?���?� Ȯ��4å��IB���<��81!��P��X�RI$���t|Uܪ���������|���D4 ��[L$���L)����U.Z;/v���=��&�YݎI��I�z��������u�Ν�XC����5�=N/�I���9<�m���9��C50�l{TSq�~n�
n���}�ƮΝ�s��˞s�p���Y��9�%[�" A6#��f	��U/$�[ӻWiϷf=���6"�Wm�h�Ws2 ;gv��W���9����0�$ᨈm��Ӓ�,��gnɎ�Y�Su�W;�F6w1�q��_��ߜ�"`��&˞Z�RH�C�l�  ]����^Ժ�;�~��e6-��I�w��l�L���=�u����=��M��uux�A[��H���ݻ�$�z;T����.��$�>M�W�UB��S5M���i6 �{�0)�k�ˌ�8��[[ͦA���wi'����*m���A:�uP㩸�k��$�s�� �^�f :��:�fo�N��C�7m�J�Z���mÆ[��e�mݢR]7�kȯu��|���Ǵ��u��I���&$J���x$/��f�Ö:�Y����k���Buw��d�)w����a�z���"�^W�|ƽ9#��|n�L­�~s�9ipLY<,CdDi��{��2T�VA�DS9yUb88�ݳ<굖�e����^���I��O-�E%p[`�\f#�N���t�db��I�Ûu�=aM��v^<��Hv�D�a��%�g��Ɖ�4Ll���Z�/v�v��ӕ�q��K��v�vz�;aօLB��� [ny]���j��Ը���ۧ[�I��ю�4�cn���p*GT2����7����sc�:������H��i9�<y�<��\�ƞ���wY�r���pn��?�Dj�5TF�����z�[�@c�h!�Y�{���{^���m��`�YB���H�)U7�׾���Ȏ\/Iܪ��S{��> >��� ��?�̐I\��~j��y�+<͈����0�*Q4����NT�Iy!��}�g=];WN�7�[����	.��TC���_�l��!�$mU^��uj���]��� �{l�I%�-����vI~���cq	[1�2�c��T��I�>��o��v`����y�� ��8�`+��F;�
�.T�u6F"�QQ-�uɳv�][�\�"��;\G0����8�7�-
�M��c�\�]�I/�U�]��N��Wޑz��s=�nf ���}M��3fIDA�"%��E$&��U �{�	M�q;��c� Sw�n�=bE!�
ù��*�u	9T�.噹�.�^�K��vykg��u�}�"�fԼ�w%���T[X�:1�c� ��=�� Y]���0s��Vd�� �v�=]0B%��NJUW�{�q �m{[b���6w){}�*�u�[�� �c�o��,�٪H]��CL80�
QTv^[�sеnW��� N�U� ���v��n�̏-Sn!�q2o����^���W��B��S5M�[���؀��n*N�����r�z�0k�� �'���$���{EP*�Ǯ#���x���NA@9�L�y1j7c�aֆ�ݷ\���Gn:�+�[2t�3R�T����o�!�z�RI$�۵�dϼ��\7��%�݄!ew���j%�fdS2\�޿6�|��{|/}o/��i ���ku���]��2""={9Y���'��ݓF�DJ���)!7�UB���� ��dЮ��o��"��f�,#5y�t��޻�Ykv�p�����,�9����O�-}���w�9��aǮ�U:�[�T��mnF/ՓvM�Q$�cΩ&�Kݛ[wi)��m&L'	��N�Pq�6A-�6��4I*�sM���ۯs""1�y���̙��$ߐ��42��h&0�
QU�Sٗb�#*�;�W�s�ꋌ��=S�T	�휪���l�׶�����Ͽ�����Bgɹ�㥮0`n�ȤOjP\ݻ�^ˣ��c�c1ŏ�����׆������꽙��D���Q�L;�Ҏu@ks���/:�{��@���,��L��9�$B�ڊ����ۻǯ__(��=���@���Q�&���7��棲��2�m��iH��ʢA#Ǫ�dA&�TvLD��%B���ʢAU(���(��B�a�w�o�u���w��}D��O��I����FFs�pv7��R�5�*&�y�����1�!�S@�w|�+5h�3tyS�{��Y�i8x�QLH��W�I����jGxM�Kh@0���u�\�OkͯTVĐm�q/�X�>�گFUFH@���1S���l���pp0r"DA	!��{\E���:��i������Y..�Q�w]��_���a��h�|+g.��A���D�}��j��b���謺E�F�;����a� 7ϏV��*���nw�㽑^��O�IؾگNt������2��V3(-2�����Dn3��3��F")���~$�z�6B�t_m
Pab�P��hCm)�������q�� �����v;��۳rk�熹9�^$�lt�՜TD"P�m�U�P;�74n��&�+�@$D��> ��ݪ�$�����x���s���3ZQ'i��TXf"��'yh�@�+ސM�;P�?nE��-�{K���kh�.�3=dB���9:��L:��f^�����`��k#r���V숽ג6r���3�(褧��B̾&�`���ļX�Ӽ�z,�:x\�{�:{���N�q�c�m.-+�+����x�=�S���I����T�-�~ܝ̚d-�
�lm��U���V�@��C(n�bdE���r�>�\{<fU�~��R<&���� ��a��@�hOq���;�;qZÙ�)�%Iݗ�G���"�a5^;���0�����n��	�c~sPw�(<�Vlm����t\n�V�ѷ��V���q[=�p���НS��%
�\naݯiV6�M��m�#�b`ƪ]9��^[饷/N~�ܺ��x�D��͈��hҭ�Ud��:��wtV�w�X�ۇ�t��ȇ6"c^�r�ɵ�}s�5�q�N\:��LMx}|���ˁ�����F���]1�jt�k�$��L��j����͚���������B8�|���>��nʘs�vTДX���<=���]���jzR��4?\~�8�F�O��u���t��n�֩t�r�z0<�6��ŋ{^��~���0�X't�;���ݭ�Dt�[���L�;�K�!}��yc`e|�5��=��8�}���{���.�=ƨIC}�sHݟb]v�/b$MY�����ƶM/K�⼵;�%��C���f�����༸�	�G}�~��U���-PF�Q��T(�Q�!QemlRQ
"�DQKYh�R��E�����D�jE--�֊������TVҫR�ie����,�em)V��*�V�[E��cm*���#�m�Fմ����(2�Q��Dm�J�ie`ڪԢ��R�Kh��EF5m��-�*QJՕ�T�b%KlZ��+l�*R�h�X��+Z"*��X�+m�YiAbŨQ+V�iZ��V�D[j��+UDcR���)KE��*�����kR��[V��mUJ�6TE�%J�V�`�+*��#Z�XTE�#*4Z5�E`�Q�b����(ĢVҊ�UD��ֱ�ֈ��ږ�X�T��R�U(�ZiH���QEkUV"��J6�b�2�T��4E,J�F��6��|�ں�Gu�C��v˂#���'����.�7뮡u��t/v�����!k�f���퍳b�q�yT�x#�9.+v�拞�XX�S��c��'X]���7��;zϖ�J���m�ͷ	�5n�;�˸�/�;N�����n^ֱ�ђ#Fn1��/'�f@&j^�s�y�$/�����갇�x�'�� [dob�lt��x��е���6r�Ք���v��s�CQ���v�q�{�	��6񫵭ً��	�3Я�`p�6���κ��j�S�<u��soO]K�@B�Ǉ���hs���j�;vv�ϥ�:':���=7]���,�v�������v��r�X�j��\c�zM�v�Ma]���Z�^�v�vڡ��M�/m̛\V�c�Z­�-�7d;ne:e.^6�\஬T9��[����n�ݴg����v������*�5��Eی�\�5�êDK��[5L�dqW�[nO	4���6�'�7 ���+�Y�m"�#<���x���v�iC9�rF5��I�<��<h9��`�b6�N�q��ӻt>u��\��=\��>�rN�Ȕ�)�	��[=�ݎ�k�Z�R�m�[#��96�A&�m=����7&�z��nΠ�}s��^M��v㍎�)ټ�����m�x3���u�s��&��t��<�Ƿ<�nn �y�v��������`�8r����W��h.x�� xώL��ݻ6���l��x[g&&�c��.�m���܃K��Ph,1�\�&�m��\=�ym��g����]�MԻu���Q��j9N�P�(Yz\�Շ�r�Gq�[N��y�\v��
�ńA�A��s�f��1���jx:�n��D丳�c��q�u�:�i9��Y-������
�۶483���=q��h���n�r��ܬ=tD�qv��Sgn]�q<��L99:��n�j�øg�y��g��#Ŵr�t�G2�[gg�t�O^�B����t����y�n��5:�۸�Ŵ�=Wc��5y�v)�dl��ִ�Kb6g<��`yZƷW]m�gTu��v�n������曷m���Wv��MY���5ܜ�1��YtD�'`8����X9c�q�lv|���c��5�Rf˷�w-�Cȏ�5�t��]��4��K���n�=�29��;�l��qN7�ś6wS�����{^�m9��g-�A�1�rS���7:��̽�C{�.wn۶~�??ma�]PXo����|I����H�ٺ�ⶊS�eoV+�鉐��#cwj�O�E�r�m4ч����s$��ވ���gL3@�Qٴ(n�РtgÝ��;�w�w�T�0ك���UX�	�f�>+1�Cxwm�@��ު�ݛ�A����`�U^1Y,u�f�S�8fo� ���
 �}��u@�UF���N�&�T�\���HPab�Pm7Ce�g�*�� �Tl��8�H5�L[�� �۳u^$:�4���۷���A+{A(]��X��[b��sunL�hԜ�뮝��!&�b��QJ������D��sD��}�OL���/6��"�Ź۪'��t�Q>���YPa�PXn@<�.|W�t&�nk���s��OK��Vb���ۘ̾cD��lƓ�;��y&�4[�aVK�Qn*u��6Ä���W;+ɐ~��1C�veOO�:n�|z�6@@�M��ؗ[�|H���!8hÃT:�]Q>$���A
�ti�l��s7�Ff�Т@=7grL�+��bp܃շxעq��Q\��%��Mx�H���$��yұ����w��sD�z"-�q�
��+#�A�&{V̜�e�k�E�mP$M��:/:��,'ڷ`u��wP�`�a���gW7A�2�u����9��Џ=�Gl��Ų�x�?7��h(6��!��M��H;7d��y�@ץ��FI�g:n�� ��t��]�),8r���o���x��b[1�{��_c��@ɷ�A��B����xt&E.�	�fT��a!�r{&*Q�ѻ��$�;gz�����@�S�f�;@Ig=+x��V�����+wc5��W��뿄ճ�x>���-�S�q<+�j�C�Y�����m.�Y{�	'�&�x�l^uP'$wF�0T0�1����넵�v����:��'3��ȂI��ڠI7ӷC���vN��D3WqS�o�̲�l��C�����>$�N��,�Wq�0g�"s��lgu
�v��=�7I�����/�����3��K�F�;Mֳrj����63�<W:�2��(D*��Q���W���\guQ$/�n��D��Z�ڬ��Ù1ҁ'c�j����(M��j9�NI��ն#����q����'��T>&�v�I�\$4�D��=�_"�3�aUx���H=��>�d�Rs�Μ�6	��&�'�v�5yr�)��pP�!�=�����rH@�YyU� �Gl��x�9���Y�Rbdwf���y:��	]�FN�w�,K�Z:�Dɩ�M��*w.�,g�LC�V�#�<�}�%���?AAe;�g��_������0���l�{�f�$��\H���U	��TI#:{*� ��k�$<���Zei�JM�j�Dm����6�<T�n��'�9��(,��L����|�	����kj�h�og�h��B���c��l��E�v�Q$�N�Q1�1l76�1K� �t�ɩ���S�A>'�w*�H� �Z���P�7�9ـ��+"ABn��\�d�$�k�$��4�g�vv6��� �fM�P$���uV��/�aM7��g*�	�x�'{�$
�ư�I�wӧ�c�:��:%d�U Hyr�I��pP�!�ۨ�70RZ��<��f$���$n6 �9��q�b�&}keD���K���[��w����w�E��r@���O{���e�}��l�)b�T�����1D�&Y3�Q��ٵ|��k��t�R*�ٻ�����q��'X�AAֹx���n���r��r].��IE�N'#�����6ܵ��圈ݜ�65�c��D����`��g�eV�{>v�oQ���M�\����|v!9�յ�=�i�N��n��Y�e�E)��=j�4�q��-�wV��i1��-��ӵ���x�ɝ��s7=�y�<�:n���2OJ���y���8�p��Ek�ѳ�t��4pF�Ɏv�n9�v��ڍs>n��s�������Wn�h����� ���0HW=T=�xEn��	2��{�T	�����̴D6`������nK����  ��U�Ux�k��љ�w.�⯔�dp�pZh����	"�'�� iJx�aL�ʺ$Ѱ� �\��%��AB�Ce�}7����o&9m����>;S�	���H�{Q#��`�܀I�p��ED _�8eU \�m
�U�׎hT)��wF��,2@$v��Q'��f�9�s�) p�H���J����ّ�t=�J]�S[��	�n�y� qsv���Yi0�N
�1y08�v�P�	 �꾪�V�N��Pw�������;�Ql�&�um��[}��S�u�4���]�� �v���<��*�sڹ�w�WI'=E��y����p[۪�.5��H�l¶�Z�Qkkc��sܪ$�龯UhYW����d��!��n�5b���o���y�=5	��w�;Ě�}5�Ot�M��rf*hD�(����OMӝ"�2sT3g.����ڠH$�`BW*�!�v�^'�g.�"�!#C�!�ԇ�}U�I+��k9=�e�Y�$��gj�H9}4I�g�w6�D�������j�E�t��{!��qZ�r=��v9C* �	RZt(�L��������(�B�a�tMY���k �e��'�/�W��%��$�!7 �T0I2p�#��u��DE�_U	�a�|����Sz���+�Ơ��"!���feU	7I���ٮ=:a��n�V���nO"Ko�����zA�b��ڨ;T�$P�ة�m�T��L�"��5v1�$`�Y"�p>y�o���62�� I��d�i�)�"��qCC��!"!Y[5�O�$tkGEv�Q�ɬ��yQ�k���޻�^Y�LT@p�%Q@76*"�kz纮vbjq�Q�9���|n�	>خڠoi�%�|�������p�3A�Du�sur6:QŹ��y����q��tϓ9�=��������guD�/.x�v�|I=O����j�tV���UD�v�GU	@&�ÆUP�f���w;�7��G\^N|Aő�ӳ^'���B�F67���"{���0�LB���h�A���A�7��go-��teh$�����s�^78v�Pl55ٙU�,�|�ogXM*,O�zr�A#c�k�T����N��r��(�=��$�L��ܑ97,ڝ��jq�C����1�"6�NM���i���'�v��o���\C��ěj_��fJq�0\CPԃ�s��d��j/`���U�k��F?"obK �kg*�$tumP%�@ڷ��cw��K�x���0y����d�Ll���U��� X'�4 �{�a��ф�8i)�U-h�EnOP�H=[>��=#v.'�MA�R��og&�첑����Ԇ�����]���TK\g������ �������P-��F�i��B"0+�2�K�͚$�ut�"�b��T��O$�͞�D����5����I��-�=j�sH��h�2�����P&�+f� z2�t�p�H Tv�Ux�ӥp:��"!�U]��T$���!�s���g��ok*�"㫨Q �,i��4�`���U�g�ۚ'	ۇ��kw��;	�o����6{�ν���W���-Y�Gr@T�M��!C������U�%���\)�
�u�o��\��N�Kcf�y̛<�6S�mϛv�gN@xW�i�Fہ����Rci��۫\nz��uT���3v1�;�����9���p յAu�U�S�{.z�,�����Ѹ����{T��^�g
�Ŏs����V}x�2q�Uc�k�� �Hx��]ʕ���ܔ������\�ۋ�M�<=u���9�r�m�T�{q���{i�n�V��D�)�7n�犞����L��5�SZn<����M�~���Dٻ���V/ލ� >|�7�[�T��5H5n��
��7[�6�eH'��j� z0�7��総F��P"`����P��Ԇ���OB։ ���,�#{�z7+^��#c'�Q �,h�
��-�b�vV��Sَ�A����I$�G	��{D��%�`H�uT	��5���6[�v�4I��С�4��m,�zn��$B��	#y����Y����f�@��l����P��Yd]��.؋��3��.��ǅ��*>8���_]���ݹ���6��G�/���~E�v��gGM�x�H9_���"Q�)1�pY���Nx�lo�y��~��n�D�/q�hI��ە{���\���B����L=��s���{{B!��ν�C-��UF�ld<���FbW�u(�M�y��s��A#b0�A;���r���J˷�y�|����	Ux�\�>5�;TI5�tS�t�UZ�g�7Z7�v��f\�"چ�m�����x�"P�kD�z�v�	���"o����MUR�1L��)����$��� ˝贪있��Nu�$E�,�O��z�@o:ڣ.�H1�=�z�9IX�B�CF��"��lx�),(v��q�̻$5�{9��&�nݱ������$�-�7�����v�(�@;ζh1ݓSm��/�ƻg�W�� ��Hp��UיUD��:��)�{�1H��F�V�1�]���n��5l���A����P�2v�E�qճ@�A�m�	�wI����wS�S�Nl��ؾ��h�B�ܸ���1=�x�A�Cƞ���<y|[���ǻiy�q�]�/v�S���{�^����P7�d�*^\��c�&t�Lo��b�{=;T�6��ä�㺠����v���I��JA��oJ�	  �}�}ƦIa7��/J���s\��ͭ�<�뷳��"�</ڒ^TY1�l�h�2)웗Z��h\h����ʪ�g�5i�5���L��4��}����'y� w�{ܷ�<:�R+a-�Е�E=��7�N����z�S�	S�9�rX|}��lǔ՚�O�T�]&�{W&O}�%��}F��n�	�����[�0Ό�w�:��b���^@޻���-�x,���>�ܯ�8���|~ko���}� �|�;�O"́�.�B��x�'��=�ZL	'�1�w�v�~����v]�tLk$�ծ�i��Ј��oz�������H�v�#��u�	�k�}�yK��w"�8�����s��u�eܙW���kӲ�.��^s{cbD�tYf7e��n=��0%ù���<|�TK��&�^䋃K\�ȫ��y�/�p�z;/V^a�OԴ�
!eqY1vot޵�ֶna�5<o�t�=��-"��+h����^Ē�x\��6���_xX�.���(۞p����s��q�~����^&�$L鯜��Ѵ)2eB�Ϻ���e͠7��9n��s��g���7[��v��X=�.�^O�%|:�^�C��a�.�{��Ķ��0  ���Dm("Ԣ��j"*�F"�(5-�JŨ��*�ЩQkDjmj�K,cYEb�F�B����"2ص�T�D�k�+X��,V,m�����R�EUT�5(�T��[-��%�X�
�[eQQX�m
���hV(�QB�h��aR��-`Vѫb	*-E�F�5�*�Q��R��ѭ-���U-*��eF�J"��*�֥�����Z���Qm�J�J�#
�V��("�iPUZ�5)m�l�1
�B�TDPDX�ik#X�6
-UDe��QUjQ��Q����"�"[DX�(�֊��j5*�F([Em�UU��D���	m����*,j4��b��F�ʕE*626�[kKTATD�#��b�����b�֤�Qd���бjT�*�V(�h�"�j��� �����ɯOG^�|�Ti�A�i8J�KVq��lNu�>$���׉'ã/��$z^�WH"}ۛU^$�-s0�j,�O��ڢI��Z֙ˊ���򼫪���OBƫ a����WTE SpN��+�vMv�m�x�r�^L�M�S��[F��݌Asb��rA+�%��gx��گtu�׈$�FL�5�:���]B���ڠO�0��!�(��M�=}d�	6"�����]��$�����ѤH#��(��L�Of�[�$!1�T;/.�I����@������#K���|H����@=>GۼdJ1	8(�2kn����x!�D>˚�$�z9��b�v������W����
�r�N10�9�Q��搃U���d�<�ǓQ5Lhܗ�:zzN�"�	�":.�N�m�+�+�u��7i���5�uN�$v�]W�]�R��p�CI�T���L_N׫wS�{
�H'ݙ�^���ҁ�>��ڢ���|�:����!�<L:}'���G�7ur+�k˗�9�nސs<C��L ����˜'	��e�k��ʯ�|�G$�\���=�2�*�W3��U{���@�"��Ԟ/�}��bP��L�-9U[�3�;d�H��ڠ��E[�=�;0r꤅�PI0����r&+gj��3�q]��/L�ggA>7+�G^�
�'6�Q0H�pUv�Ԧ����wvI�.�:|�&2�����rJ��_d9싘�A���G՚dJ�1	d���Q�m��׋>��o�F��NŹ"I�WeUA;ӷT`ج���O^��d����^C�Gs�(R��a�J%�$�a&m[;��W�3V���u3#hV�{����o^�s`�X���N��"),X��x2��{C&\�7;ctS*�t�'WX�n)�gg����=�m�L[Z78�-�i�!�@�m�tr��yӓs�ڸ��z]��J�]�c;ՠN�t	{oHm���m����\l�T��gۍ�n������){i�x�/<�w47W+����'i�� Jݻ'&�0փ��^�\�Z��IɹI
�ok�y�t�ˮs٦v���=�8�V�5&C��sN.����rl�����C!���·���!��*�S>DA�Ω�A��r`�٫�{T@���x�/z�� e�p�&T6D8q/�r�\��M���qH�ު�O�ӷU�L$�e��k��z8��T�Д#p.!ª3��B��IDU�ޖ���E��P$umU�������BnA��[=;���ȳ �[��(�N��UH�F�1��r�Ăꯦ�< �A


�YYTO�8�6B�k	ۭ�wθ}�u�D�Hޞ��A�F�S�s�n+�wP��Lh&�X��M� �m�� ����؏�_>|݅���\�҃�/��O�B,BE6K?��� �og�kĀO��>zGrcOm�݊�;�<	'�v��7��pAq�UET��/�T���/�ww���ݜg.����j��E�^�y̾�ˣk9��+\=��w�r6�:pZȊn�i�P�����|H'vv��$�}!r�LuU�S�O71�g�z�t�̬m�Sl�p�1�N�����zh�����A#�z�� �}(�H+%j
�8UFo�2�ع����O���H��zD���̥�lHM�rm�<�{3�h*�86�6��!���x�/��o�hL�R�!��5ճ���veQޥ5���WC�� ���6�1����^�gt���sm;�ګ�ڤ"�7�;�T�o
	�]M���AǑ�>�ٕ@ˌK8EY�K멛��Ѳ�:Qh�E�H��dS�ٲ�_hH����<|}>�GfW�=���v��WUэ�B؀�(@M��c����۵D��B���o�p|��;ڋ	��8��f�x�%gf�rsI�
�O�
;f�ڠ�i��2�z���
��bm*&�z�$}����݇ ��[� -�\ہ&���sܞ;%��d�[S ��d�LE^Ux{����p5�a���s>��b��A@��
����D�����wy�)R�a�d��xd�H#�����j������8��|Z�3�f�ѝ'NI9�d�ф��E����;c%����{�2��1
q�����]�D�7��{2�^vae���r>'��B�~yȍ0�'WM�����NyյŌ�_� �[��]խ�N���~w
ɞfo��	"��&�fMUmТ	��M�	��"goYq�G� ��� ��4	�(E��Ѡe�=W�7{6�H=��T|H�>��A����쵃^b�9c��^�R��Ƣ)ֽ���㝺��v�b?ww8���XF�ʥ(�V���5�w�e�@sһr��� ���)��kkG�}TbƸBI�6�K�ܪ�A����EX�j���7�^'ā����� ���WH�8�\+�%Y{vZ@k��bA]��Bs�5㌮���Q����`�!^�I����yE�Zq�����tqZ�u9�k� �������A>�}T(V�\6b�'o�2Q;mFn�5g��V(�I�{SG��(3ف��f&���=�:	�<Ў�� w	o������p`��~3��d
�@�׵TH$�tl��ҥ$�!$�-z��[�3���y4	�>&; �Ds��� �����<ô���;� Z��L�"3^5>Gă�kՑ�rB��{�mP$|cr:P �y4=���V�����s��W�>�������
(����Ҟ%[�nCk/��k�o���,����y�ޕ��q�{�^J�B6ʡ��n�mYq������w<p��w���pMګ�ҩ�ܜ�s�k��rS�A�0����|;��ώe����^ڎ-���F�Bvͤ۝чq=6;+�<4c���b:�Y5�xD:�J�����ۺ��a^�ܧ��T�`�v�\\G��Ӑѝχv�v���vw=pW�ѳ�=\�GDg	ں��cOo;I ��Y��^��F���E�^�ܨg]s�◢!qFqD�u��:�*Zw.��܍U��F�6��4�/9�=��߽��I�F�U?�{TH'�7����(V\Z��,Ӟ�I�w6�BQ9��E;@�0`�	�8S^3�{#yϹ+�ܢ�^nT���Fs�>$��yTI�7�����C����j@M���Ȓ<b��z�'�ٳs�l=��������"9�P���a$�@��ߝ������sdox�UD�GĂ}�hW��s�zr�)quϫf4���2+�LAQ	1	١Z��cp�B�꾷R� sW�&�.�$�#�mz��s�^.���F!���ϧ������	"0b������!]�%�:�s���#�.Eu�6�v￯�����g�uD��D�c^uQ���P��Y���b,�����x�;�d@��@aC!�q�aoHޛk{�F�^���)�U�q��O�K��;�'�}3KH"}����Â0n�2,>XO��j�L������!Z�� ���T��|A�~����W��#��k�ΐ��/>"��#B�!�h�9��D�{���$������SN#NLs�G��MGȃm��ߋ����r5.gJ�|q�uQ��n9ڠH'�wF֧�eP�E~%�6�9T{TƄ(���~��P��!T؞��f����G9��O�aQ툔/lL�~ȸP�@>���Y{n݋��8D�L%@v��;�-�ݸ���7��H$��D��4��nF��{�D�J�zdJq�S�٪�
co*�$�q����@�� 8!�hJq��5]2쇉f��{u��$v�ڢA�6P ʣ*�w%�U� ȁ1��Y�ܼ��O��]���Xr,���}�u��k.��խ5�Q헃�ո�hn��kCTv�F��-�8.l��E^�;���Pd�*����]wK�2E��bH�Ah���<H$f9�@!wF��
+��h͙콺9�:v8���ݚ$!n>2	�>�w�0kD̊y��S%��Ux�XO�!�0�.$]ђ$�=��c9�)�����:ʠ	+��^1������t@/UǺ���4�2|�E�B8I����NV�{Fx��p(O����9���ß��ߟ����=��+�̪��#�Ȓc��׌Q]%�A��Eo9'������ԂH�M���j�n�D��B��˜$��L�H&9�UNۻ��Y2b2��Gd���{-1�m�����9�РA��s�8�5u\[�'ĕy(Ds��$�f!pm��a�>}7ն�$��y'�:B$��E����=Y�'b���[@�L�D+F��D6���u��%��	��&�t����k����;J'1�Vz����嘝��f8�U�vݵ��t�%�
K��$��j��^У�;��׎�t�����A� �qfI�$E=�H$w9��;)v�������:/KƮf;Z�m����p�|����5�g0L@�|I��'�k�C���[�̌2	1O�h�O���W�df3G!��N�5�:B婢'9�҄�EWN]N
b��#d/�*�I=�z���j�3
����`,� �BLD"�-	5U�B���=4	�'�nމ�}�Dp�
��2x	�S��$���P�-|�C�f��C7Ho>r���s׻���������U|I]Ѫ��6-h�;�����x��*s,[jngf��]����U�^�y�S3�k���Q�}��$ I?�H@��H@��	!I`IO���$�Q}�TA_�W�HO�@�$��H@��B��$�	%�$ I6$ I?�B���$ I?�B����$��	!I��IN$ I?�b��L���͖Eտ � ���{ϻ ����о �z��UV�J$���+`��B*H���JT�J��U@�J��HIJ�$�h�J�)H(�  �J���I�)AH@I �*U*T$QP�R���%*�T"BUE`(�����U$]��@      (                        � q@     m�D|���>���j9+W-R�o����������账sjQ��D:n���n R�Z˙�1�7��UE
	K  9��ī�}z���n� ��0�7��ڮ���/'�������^�;����ޯ�:�}n�۹�׽{ww7W���v��"���� �        �����{�u[n��U흯7���u���u^ö<{U]�u^�ٽ�y���b���π�)MU�w}�Ί(���^�%R�� ��]�:%T�ԤR�������4�zΞ�U=�����G�[�>#]�uI���� �}-�J�1�}�9D����7(��t)�ty��@�U$@� ��     ��>�h�ۭ����W���%��i���7l-��`�N��Ѷ�Γ{�y���ꗪw��{�Kz�yfv�y�"
���P��}��]��������:T�s��U�������GN��y��OF� ����ͽ�q�[��
Ww99z�*�UP������ �     ������{r^^�V��g���z�� :�nN�mw��E�^{Cƶ���v� ��9�^��m����L"�5%B�� } ���ϯ;�7{,��ޔo=�\ky�p�:�3޷zv��{�זn���{6.�6��mu��[U�*�   =      �*�oq.�Nm�oU��7FZ���We�k��Uۖ��SNv�1�Nf��d�M�iF� .���l�ٝ��{��E �[�����R�嫑�>ǻ���6U�WK3[�R:iu��M��R�� 4�v�]3��Nv�cY�FN�k���j�      T�2JT�  � & ���~F"R�@ `0���O�*��*� a@ j��H�MD� 0���b 4�!�*� 4     �PA�HИL���G���=OSC�6R}?�����f7~�8�[�~�$>��k�͇��ˀ|rf��I$ ���b��s
~P� ��Y�d�@3a	 ����S9��BjH9�l���O���O��@��8 ���CA !Q���		��H�e��
�$ ��H}?�v��~ ���c���_�� _Q'�
8��c���,C'䇶������~�!�,/�������T�(�nˤ�ѻի#v�$��������M�2v��6Ej6�<7�̓]�.�d���fX�q��+v��N�Z"&˺�X!�E����(����^�J�{,�a��!��,�T�[��	_1���Mm��,�|ky�9%k+.��B�w�O����M}��z$��~M2#CP컗�D�
�@�RM���yA���҂�P�=��6��^f��32eͰaW�+v��yN#�c�V�n�)��V7ZhŠ����ׁ���{$h-�h�b���ش�vQ�Z�r���,�bK�����n�ֶa�L����;؅�[�޸��P�$��ʼ�5*0����>,آK���I�Lb��ԧ�'��Xi돨���u0�{��9ZkI�(�T]f��Ԇ��p�F������� �bsi�/cV_�V!"���GI���eɶc�9����#�VV�9�M�d쑳P�mHބM�.U��5��ⷈb���m�>m�������CT�v0Kk��Ų^&�cs��̬T�����I��2Z;�T�x�L;�F�إ�ڡW����S{t0Чj����KP��ɽ�֋����-51���V��|��˹vhDv�����)��k2�'R��)�[b�����SGU�Mh0��L�J��B��3h�oV�@ia��hm��c��R�"�F��2Ve3-��$��f�s�A�)��U�g۲�ͅ��{!�#Yf���K���U�Ϝ�:��L�}���A��ɛv��v�c��0�`I��y�
��^r���r���]��1?��U�$���S7hA�u��ˤ���Vb�P�)]U�*�̓*�x��L�UE�2���aP<z�@2�K*��Uk��ӹ�d�cIWR!�dr�T��x�궠�
�W���$��%4���[X��rkR��b�֫mf[,ѻw��Sw�F+��Ie�������ҙr�s�x �j��X�����'��ݔ�
Ӷ�S@�E�EJ5�$�R��6}�8�E�ONRۢ�ku�w�Q�E-Ġ��$��i��l,�@�1�H; �����3h�ǋvVA�m�V$XA�RiE�l:/	�e�ơ;{�[���:�n��kM�ʸ�1��ܬ��#�`А�W�`���X��+�у+%dIٹ&�b���H�����6��4�xdqb�����LW̦֠.�Y��յV�q��3Rƾ�ؾ�,�S�]\0f�-#�bspL��j�X�7f�����܂�w���'�\(�F�PJ��3u֣�ݪK"8��W�"	D�����:��ҭ�"��r\E�uB	�$�+�S.�hbgu�����k%��)�f�>�P�r8"�&�y��c;�D��0@E�W*��a�1�i��wI�X�����5���z��ɇ��!�I�6�P98��e�	�w{B�O/n�Q��5��);Q�Ѓuݥ��ӛ�	��J�lU�cgv���n��sk�OdF��m��\�V(Y.� n�5���K�_�Zn&�C,��������tqbԣCh�����֝��4�`���Z�1����c���+2d�Z8�YJZp#FFSo:�����b��pjq�J��4sc�+rH��0Mg��4A�E��J� ���Z�kkr]��̀ñ-��D�0��6kpj�Q�&��ӑ�����,V��:)���G�f
m)b���5&���6��h�!�Ù�A�Q��cNT��V[���d9*�պPȅ��ؕ�4;�1�ߜ��fPD!���F䖴��߬@�d�;Iݲrg�o0A0]j�	Wf���4��Ꭸ��a��'�w�
T�U�-aA%hRV��U�`��[1X�3A˼�G]T���D��0s�����pS4kU-+*��{njۻ,(�L2�f�	i���=&��kn��A�ot��e��B�57��,dj7������zmM�6�%Ͱ�m�j3Q֬J=�R�Wz�ið�v[�E7��P�V�:����Ɔ���ԓ�+B�+�-��7��DN����ͪj���
��l�+d-Ժ�l�hf<�ӄCO�5wpBHʍi�6ĪW�Ŷi��#�Y%���Y��%�7X��&�kYw��4�a�3��n]bZ�=�
=q�:�A�lөN]�����&81�ԕ�ĸu��X~P�:��������^�%Ha�V��{���f�2D��st�N�������֎E����Y��:s6�[�L*WJ�V�3BӦ�JQm�h�x"�/r�SThB��t��)7��*x7q���KwU�sW7P��\Y2�S�.��Ҩ��p��M:h3%�xl��X�]`��Ra�`����Q�h�˺2cGaY�j@5K��e�5]�{A�i�X&��:ӛ�GY6������bn��Q����c Ƣ�%Jk�E�e|VM����zVt*g-�Ҹ*:��h���C!j=�������Ӹ�w�A�9��J�5����ն�;�jdW@ǻ���C!Q�9X�5n�S^�)��+cwIBY4he��V�ز^I1ǐK����U��"�`��co^V�T`��E�]����+)=0\�Yo-�d���d=R]�]�6e[�N��״V��^D�i�
�fYt���2`f��`c�Ej��غ��r��n�\�h��Z�A(YP2�H13F&�(���ta3j�6��p��ŧ(*�'�@%3J�xhۂ��m&�н���U*����Ǆu�+�j��:��K�]�qƃow]�o-�a��[T��7�&kn�2<4�恦�<w�Y5	�-�26��/Qس�8m�P�o�u�I�M�oH�u���L�٬\�B j�JZ���-,73Znh�����'6��0��,�������i3;q�ef+�X�Bg�֡,��zkqV7ui�S�Ш� ~jPځ��*�N;�Ғ6_K;I�q*�g�q�
�(�,�eb١ԩ��L͆���K�e�Vl�Ɏ[��,�3f���&�V+tcq�Z�����:��[V�A��5ݴ�ۇqQ�wTƚ��� r��ZPǴ�����Q�e�oB�L�Br�l$�Om�fe�:{
qV��H�&TX̂^�.��7{��X�R2����J���\�e�2���H�*�++4�*+�J�h�7��2�}"G5U&\9UMj�:�OnS;�U�O��%쩍b1��r��ld�%۹�X#0f�t̆�4f*�ݠ���
�Y���K�-8N�eմr�Ӵ�YK&�r�H�BSt)֑���37*���jb���2ܫ�t�J�,�j���e���N�4V%YN��̉����*`3F����ڬ��ڲm�F��_i0Hʁ�rR6VP�L崰͕�'�2�2��c�Q��sm�ףH�]=���(�.A����v�əF�9��e���͢��+U����ܓ"�E�mJT���w�,�
�B�̽{���wL�U�؉`��i&)d82�m�\����	��U��YHc�ȭ�BJ�&���M���\����1d$q�K./�����.(�V��(��͠R�)�3��Wm�0��.��{cJJ�k/l�,of<WLi�n�F���nY�i3*��V:�	U0�,�b8�4�Qw��<rƧwrm�#�h%+VTֱZ�YoN-�������[-��R�)V74�Tsj�D��'u#�o�*���H��a5-Mh�K3'�7FK�� �"��#k�xN�!�r�'kn99GN-�-���!!Ssk7�Z70Sl#��!��S�q�x�e
HF՛�m��"f�P��a�׆K�Mab�G����I���VeR�5�/�]Ÿ�0lJ�a���x^�d��m�
�D�j��	��ƅQ=��L�F��-�u��4���7o(R���HJx�x�Rfΰ�V�Z3]h��mɑ���u-\!h8�Zt &�2�p��$:�-���DV�l���&Lx��#J�������V�Dh5����׻{��UHШ�8��V��Ѷs1�W�L�L[�c8Uq|��������L�����P+7wv-ǲ�8@:3%I6k�r�JDZ{GH�%f]�L�)�"�6���!���ga��>��9>p�+>��2b�2S{��E����Mdc��J��e�x^�h)ZPcd릵cq	��L���H�BJb!��^(0�ɐ(,*�,[_`//6Ӻ�^nS����Vr毳-���ַd9A̺!�q$m^�U��:+ԫ.f6a�Nf��uYb�nƕؽ�-V ������d1�N�w�bq����#kE�� �x�fk��R:m����ͳ�
X��AIZ�d���&�n�#�W�r,�p�8�O��#Ӻp�ɥ��$�s^*OM	�"pD�LYj���e�N`kH��9�q(�s0��
8� މ�P��n���A7PxX���L�T�T�XF�ƍ�����-%Tt��V\��?�����/-�s4��W�����ӵa��t���a�6�f
�G[fSwdX?As&nMͽJ^ᡌ��D�ڐ�N��K5m��B�:�K��3f:R��Q
��ĆV��^����bV��UBl���$�t���](�͡Q�@M=E,��̊���uPAY���$�ʖ*;A좖k��$�M�uU��q�4���b����4�љEޣ #]`����	EQ��a��g5+
���Zt�Jɇ*�k3<Z��fS*���@�j�G��XBS�,�[W����U�͕1�;zތ��ݵw
�"��G�)ܺ�ZƆ-홌���e�XU�Yq12��,�%��-Ua��-�.����i����k,];9�Q0Td��F�au�t�(h�傆�5��
̛3pA��U��M3SX?vh�*$��Y��ke{�UVj8�a Q��t��t�4�㛍��0[t�t ���˭�>ȡZooJ�=oKѲ�*Ԫ��(�Uʍ�%M�$��Kd.��(�ܐ�On�%�B�{��p�V�J�plS�Nޙw*�cҚ�����%�,^�{1������{���q;��g*��l�e�YI��q��jӔ��6�inm����a����h���}���FoB25��̍^��z�!�?�⦆ޫX�M.�$r�oG�7Z��q9Rf�ť���q8��A�4H�բr�6�ց�)�e]4�㍀��p�pm�X���h�V��P�X����$�4M�.c�omW� [Q�o��{��G^:kq�V�d�Ӫ6n����ƨG�ђ��5J�v��N�E���$��g2��+nƠ����9i�'3��2�*$����%M���Q+!#Uh�� ��ǌ�/�B��+m�-�7�҆3n�6�.��f��T����T��f	UMe�d,<����(0`���ה��4`�,+cn�"�Dn��=��c&�F���b��q4�f �0SxP"�Q�z5��@���/oQ�H*�vr�JZ���]���/��B�f��"�6�$cSd�&ᤝi���%ґf��2f]C I���ɷ`����Q Ȍ��Ϩ0�U��.*e+�++�;7�(�, ^:
��I��4V����5Wv��[�1B��
�N�.����1�i�K h\S��h��)�Y������1e-ʊ���S;z��kn���**гt�
*b�W�&�~�u�����a[�.��SP�J�.GI���]`���t+r�8�9�m�d�"�m���VkX̂�N-�Ĳ�������H=��&+�����A�M.��,m�.$r�D���aHfұ@�KT1��F���IEIL�����bsz����2��I��#���;�US!�Sͽ$�ؼ�U� jC��1���qJU��ߛ���c�G1ު�-M4!.j�܏��hzkV�5��mލ9�JwZ�k�we+un�j8
���hX����\��q�nT�4���.��������
��q'��R�U/�5��J�az%�.��\��S,!фIcudGl�2���zR�0ὖ¬8.尩)�t�o)Qn�*�GRv��+@��i���M�lh��V��K�Y)vu��f:�z�Y���k>�?#?'��x��	������q��T@N���uѽ?���vxt'R��Aa$��,"��!P � ,��$�E���X@���d� 
H)!E T�$+B ����HH,�R*��@�(E,���d�$�+ R ���Ia$��� ��Ad�$�d�X��"�+ RI��A@R$XYJ�* Ad(XI$�	P
BI����
 (`V (H(@+��
�TE�$Y	$P�� ���$�$ Y $
�*B�$$Y$� , � Ad��Y�}_��~O}>��/�����'��� �� ��=΀$!!>W�B}�=�V���d� $'�?1�w�}����L��O��S�<�����d�:��;[�詸DU;����/K�C2�y,eh���U�<�k:�"���C1R��v�7�_@K��;}2�e+�j�-��N��1dU3�]@�恰mi�rv�"�}�_.Ŏ�K��[��M��y��r�i���m��G�ƫ���(��U2��ƻ��T���B��
k�C�V�[Ϡ�LVɕ5��A��v�+1�):�P�����8�B $�<�Ϝ/R�$�Fp�`*�n�F2�I
��S� /G�Ȼ�9����K��]��AY�z��ל4�k��g\���:%48Gma!(��3 �u5/�y+vZuvQ�Y7#=�l�mem��7-�ae������˻i��s���i��ǯ�吮XUÈ;c�i�ѳv9R�b�P�(���(�з2�Ca
�`��{I��{�I{�9Lhۖ��E��[�Ǖr��ɸ��6�7�EY;���������%�s���6mG{�j�w�1�'Y�րK� ��䖲�۳0IGVm�����׽�2�2�'7�������j�܌t簭��y���ƉF������R���N�N�.��z.9k��s�djr�ur�u�����M�1AN�N	N��ϲc����c�B�7w`�9J]�tr$��PT�[��Tߺ��P��Z�Eۭ�������܇��Z؍P���ѫA��up�+�kȆf
��#s��r
]���p��@��%� E&PW�kmRH��o7
�!�^�nO���!n�R`�z�%�Bu��x�D	ikԔ�-˕�qψ�΍9>��bW����V5��J��[�;"u6�s�N�%/�^P�,�W"{��F�b�/_-���%'[u�S'��:��)Sa�����󾹜r�m�c��-i����]��lXJ��Kԣ���S�+:�pG5kMg-9�93����7Z�E�KSl���C��g�������Q�uڜ�1a��%�7WV��l�*BU����sI���P5.�׸r("�g ���#��"ݕ���y9�AWv��͙O��6M���$*�SJlYK����(�z=�S#mC7.�]����9j�D�ϺAg�����'r](�}�y��O,�9��ud,��f��7�M"�ڔ�+Y�lc���];��qa;uV{uj��KE�Aj�+��Dp�u\�J��b�ܮ����=�}L�{D��p�Cгna7D�їD+=��4d�ڨ��Tie��ep�]�ǅb�j��A�����oF/���c"�b��L@�+����^}pR�h��v�M���=l��a�hZ�M�����م��͙Aب�E��/,�˱mpjܵl�ɹ����$
����`����]8D�D��.���x/fǤU��F��U}jp���.��d��������7l
��\3�/*d�����ƕ���J�ܴ��tp�ĺ+6�vFp�N4���/��0*쫐�Ex����ī��̧�D�z魻x��Ɛ��]W	��w�����c�o>��7�9��{�q�xh����'Pz�V� �++K�����;���	�Ѝ5*�x;�{��
/	n-x�6�J�o���ޞ��K��0eu�ҥ��^�6T�Ý�Dea��*��[�!5˅=�0٬����u�H�ٓ��h����,CR�udhk��f\�0���ì��'	�]�WId�hSw 5c-�SyFk���mM�}L�2��]����`�����,{p5z�QŅ�s�ʤm��V;��P9� �+0Ӱ4Z�!�ݸ�a��p4_V���̺�9�2�oz;�Kh����L2�Q<��4;)nl���I��C9�Ϡ�UD���5�<�"9����|� pKe_*���%hC;s��&;��L�$���������9�W�����CoR�6��n�ɯ�m�+�u�ؖm=�YAM�����T3�6J� n��4��{�H�G��g������O�K�b��!�Y�f�]���U�n����ϗi�!¬��]��c��ˇ镙e�U]t�H)z+�r�W�C���n�M..Qq���t�Ww��l�Q٥ܣ(8����2h��m϶�	۽�N�:���j]�;EYC-���#%fN�����+&k\5�Ԏ���u#yggء	a�:q��I,�= �F�i�5_	���NA��7�+]H�X�̦��+[WQsO�a:,���!�v6ҍe��\2���4q^�J�H��Y�e�d��7����M�nl�P�b&:�S�;�ڣqgBr�	п�;: ����n+�}y��Ge���P�x͂�✑�J�0�r�3�V�&s}i�3p�����)�2�f���5�i�(�2�Ӈ��躬wG%�j�T�n�;���Z]��7V�:K���.#�G�)��k��)f
b`%��05k��F��QzQ�E��Lju���`���x�ur�<���Z�[鶊*�v�7zD++)�])���pV!:�#������a�j�'�C$�{�!e�(yMmn�FY9�pn�k��Û.�����n�i��j�� �}�§qTك4��OlSx��ÿp���H��+Z4�myF�+u�aO�x�'#'*Y6�N7`���]g5�bn2#f� �ګѺ˲ W|���4�^���]O^s&�Ϸt�nc��*�|�.�w�W��1��=v�@���0T���k,�yMn�i�=08�΃��ed��
��Y�E��l>�S�â}+78�}!�\�fI��7m�"���򚌖4}�KH'-t;����2-�qAH��W,L-��������L�5�]�XqU�֛w0R��w[Ѕ�H;���XB�`m抺y�����}*�uG��L�n����mep���"�Mm�ɺ�UV�[��{�ghOT4����㜒���p���ޛ�|ᆹ�˾K��j��qǻ��6���-"�v���Զ�NA���SK�,n'���T�uld�%�L�)ZGlZ�1/�6�Ҟ�
�F<��t*�8�;�I\�;:�m�mZ�4Rz����6�(���UY�7_b�fM��y�^U|�}P��� �zC|&q]�K���٘���rw�����a�n�F͟�7Ip���M�J�5���X���n�&5G�w%�`�������ƥgaTS��Ia��v�s4z�Z:�N�<J�K\�6,7`�:�^D�c��r�2���ZU��d�7mm��JXb�wo�&Vi��v��s�����
܌I�>�[�6��gn����ťb��&K��&��Բ��F�.N�͙O)ҽ �/��p;�����15m����`��)Oq>�YF���*Tw�h�iΉ�����Y�n�&��wt�(��8%�^k:���'6ZDet̔����H����x{�_.݄PGoy۱z)�q��:��Mb�Rw-�L�������ɷn����m�����ntU�0~�b�c�c:���������1�&�V���D������S��3`꜑����T��RK��̮�pєփJ�C�[6;|���b{�Uͷf�3@}�����w*�Wiwً��y��%�K�l,�)�]knb�n2��y3�-;V��\�r��Lv
��Tr*��wz��={k���Z�Jی��>.g3]�Xc��uaձƈ��Wg_Ԫf�u���3����:��X���Wh<sY��BŸ�����Q)I�n�w�����j�9���rI�]-�P�fE� ��t4iљ��lñ�4^)q�l
򳨼[�N��d��H���^�P�˼n�\�wj*��)N
]�k��9_g������ӑ�F�/�'$�&nS���I���+��3O eoa�lQt6�n'��x~zIz�|;%'&��(�Ϲ��ќ��7mY6_Y��n+b'1�EUgܧ��{�w\FĊ�r�	cE�� �ř��V�fEaa�rok�Qi��3��,���A���r���om!��e��eĕc��b�Q5�:fo&G9V.�pJ��n��[[��|��=��,�*�٩t�E6�\�M�M�	��~t&.����:��וT�ݦ��d�\��L�Vuts딓��D��k�7����sq��B;�E=<�m}M�Op�7�\#i
���ȭl7�(X�\[.��S��s޸k�Ԅ�J֛�y\����Fv�@w�]�sq˪L8�w�i`2��"�Y�7�m����)fK\0��뵜�-
��W=)>�-&6��u3*�Z�p��p�w1"�2�M5���1�\�u���}Qfay�f��&���.��'z\-;��,â�j--[�l��L��ƘżG�]���]ہn
�jKn�ꙮN�܈�@�GOXtj�7���Ffݺ��.�+�u��9/
�Mٗ��0F�/�����Ϊ���]�2��Nf%�ah��Gs1c��q.��՝ϋ2E\fɸ��x����t
v�땅v��]N���m��EGA�zh�U�7p�2��hu��.ϭ
�bρ����e�Q��ա�v�.�T�G��`맊��f-Ϙp*�s��i�:۵/i�J��z�1�W]�υ>M�JU�ι��m�g&,a]�抷wy�'�L:�7�a��Vnr��@��ή��5�
�g�ia��#:U��^˔��ck�QfJ}aU�Z�F���є\��#�����,]l�*,�΢�1Q�;�:,]��[W>ǫjY�Z�W�mV��5�c�x]��mq�-uj��&�G����2�����g0w���m�xa��I&n]R�&�Dj�.>�C[���23	jG�3�y7P�2V�oQ���]���T�
�/�RF��=.XB��ޗ�3~}I�A�&�G���������wh��}�;I
,F��o��FLho���H�e�1P�d0N�j����z�����՛ٰWG��0�����9M2�˻� �|i�VU�椣 �c���
r��.s�m�츱�3���f�����ũ��ך�8V0��K��L�L��[@�&�9q	�m�o�,(���9+p���mJ�8��I8�}���#�N�U �,^�D3�ۺ����^�]��wln����VU\Ca���8�G�����މV���5�@��������_ 28Y���3���gy}t�M׉f�T9��E�P�p�B��7�~`�Q�%�E;q(�0�)�wq=KDu�R�t�&�6�(Z�}]����u��vv-ӸѳR�u���N�Y=ntӹ��!�q�5�Q�#��i�]w����p����f��Olf�l�vK�9z4�R�����%X˳[L��Ya�L_k��̦�Ka��-͎Uͽg��[�+&�̽=���esU���Tƃ����,c�`��.u2���(��T�[�|H9���ԍh�a��u�
��` �Q_*�Y��_f�ܮ����d����{�r�"z-!R�ve���5��Z�JG��� @�̨[R�3�������\ܼ���E,7k�F�0�V�Y��.k�/���0��	�{)�k��r��|ֱgP��f	�X6�����ٹ,��L��,ns����-گ�cwwO�,1�f�x��'�*���W3:�`�	\4��lM�g�m����ik]���ѳ�"��wo�"�	գ����4i_N��D͜A��M�$"9u�$�Vf�R�'��k�R��7W��q\;f7׉�z�$����k�{�X{�(u���̊��7n�����*PN�B��3z:w�
��h/�6�WV�2���k����#y��L�X���B$�q]���G�a��<�������YK�R�
\v2,L:ڏ��S�hA']��X��ݝ��7�.�æ��1c���,i�}��ֲ�����˖���'=�K�kZw�lWu�q�$z��<�F������K.ʜ��}voI�((��N�:�f,��s@̠��%bJ��˙ה�Vs��l4���w�iFbw[a\�-t�7m�x�^m'�*�S��q���V�wX� r�ob0�)b��ͽ}�G�xr�b��V��ManCX��)x��Y[C8Δ����k�$�+�YPVf�h��|]���� $"���l�$��4°00v/�B�/�(�D"�8��i�*���gR7Z��5�tg=�����V��{=��ݣ�rm�7d�o;d���ss��z�a�[�{l�����v�x���:\z��mȫui�bz�w[��k�5�çF�нG�\/F6��v�����磱w4��	�q�����Vy;m����zUA
��|����
�!e��8��p�Y�n�ֱ�w��F�4��i��q�,]x�3���� ��i�C����Q]����k9�F�7n�����-㮭Û�#�������n7>v��k[Ɗ��H-x'/.tf�zxݶ�q�;[�ܯ;���;w\�6�E�獰=�lu����Kz�;�SnՊㅻ�l�9��#�}�2����==n��و<�e)m�S���b�؝�٫t.z��F��c�9f^��8y�/�Y������/=��m��vƦ�n�7���r�qgrz���v�9ʊ�A+7.����Zڡ��<��W�g� �>5�+�%�����g���:�'�c[$/���q��=���ܻ�c�G<z�R؍[mr*�ܼ ��`]����� ��n8����7l�y�+��i+=�m�[��s���@�"�,rp�.t0�Un{`��nݬ�7F�v���u�fS��oε�ju�ct�۬���E����{*�gg�Z��6����G8�o:ョ=�;����+�b,�˷l����k\�� Ӻ�g�mݯLv�����v��=�y��]�3:��qj粳�|Dv�Α���:��W���Ӷ��p`0�a��̧;Re^qq���̻V��v�qƋ��]<���yy�	��ɞ���Kn�.��5�ܺ�5�4zA�N�u��16��Xힹ4v��v�1�;#�
s$vj�r�q1���\�%����j���޷j��Vq�m�2n���;]b=��Ȝ�'	�bܼOl�1J4��og[��Nݱ�S۪����c�½qټKksu�c�����[�\�l,q����!��y��Żq퓒����L�]7�"�0�3�V��b#C�v�;�C�;[K�Q�`��{g��
��y��ܱ�u�ݨ�t�I�ݍ�kO5u�W�v�:7F�
6�u#פD���m뎡�0����_��M
' 
�+�룃>�J�������9M�݌뛮��î���!��^�r����K�gm�dy�۲8"]���"X��&��C����v�#�r���wn����8�ڮ�1<\�%�	���/�띩��1ulFu�(�˒��d��9g�.��3�![vV�x�X��]��X�<ۍ�͸ ��P�����k�h���6yנ�c�������V=,c[�݂�ml�u=�0�H^c�`ݱs�kv^�yͼr9�<�[���7���v�ul��l���ώ������շ8�s������
σ�p���G:ٷ�N����n����8G�*[W3����'�4��э�v^�'��������f����-�m�c��ƞz']����'^9��e!K]tn����z8�^y���v,Z�%M�+���z�v�����qv٠+ԉy���<n�8V{v�ݥ]:{:[�Yj�u�F�n6<���chm��9���(^�M>ݭ]F-���7]h��n���F�����88$� M�u��t7q����G��v������@����W`|x�O'8yBݞ5x���;p`��\2tM���Gt�����V��;p��k���<8���3�S0&���OQ��ǳ�mU]�fk�2fږ��py�*��7z�\X+\z����]�v��^-����Ufk<֬���n�q�<ӌ㶮q4�H����e�vD�D�Gv(L;"�����5� nG.����]���ѵ�*w��\���%�$Uwn���'b0x�5n͇�uu�㌰[�:����պ�t��C6��ގT^nSu{t>�1�3�^�	�v�ӧ��s@�����M��\<=��������r>���������V+�U�Kg�D��;uu�GvÍ���%���9OT�tq��M��6�EuO��ݟ#=��ݶ|�Dp�����XN��ñ���6k�g�8�� ��	��͎+�F9m��3q�8�v�X�sSS��B���x�#;S�Yȗf{]ٸ,x�y��wg�P2���=�ëeWi��������5�ON��n�n
7�{qӶwomp8�\<k�8���7m�nݞ#d<���ݒ�rd�CXȾ��]�F�5�J�\��q���]�h�������m�ʼ+�q�m:;Lut�q�Nw'�G{m۞7�kc�g.ہM����lǗ��]�����9F�q�u�7a�i��[.�;@=��s۲�i�ubÅ3�G0s��N�h�"y���vk�=��l�n:��<u���m�����՚ �S;a�����yG���W�	ň����h�����g�*� ,\����7S6nK��T�ϴk!	�v=�˶q�=ۋ3��u����[�����ɸ=�Q�lc�mn�P8:�hy�u�BT�f�+t�b�ځ���n��cn�볱^�<�[n^���.un	�z�b�ݮ��Z�s��	��WLl�07A�9����Yڰ�Û��qk0��^͊��wOX�v�s��Ok��XR�2rۊ�R��0�/���7=W�+�� p�]<]���X$�=g�nMn�l$����/nyN�]�::-hˈ�6����[�A���&-�)عf^�:�� 4]Y�۱�m��ٖs��=dK�ۜ��d����p��n�WXi���Gu��	�*m�¶t�����g��a����Ϸ&��˵���8�윗d�ϷN��ܨA��[v�֒ݍɣ6�x�n('�e�<Wlnڍ]�`��4��ѹ�,����MVt���1��o;^v�g�/5��j8˱���Y�mь-\{sN��NkQ�����t�݅a��gF�v��.����!�v��{�<QX����xb�ln����q��m	�v�4bc+��DEz��Nw��O�7L#g7[�W�ur��E����6<�ty�wpUku�F������V��t6�9ۋs�[.�(��/�m.�\u�	���k�n�ݺΔ�uk8�l�q\���|�s�^\r��k��8�=�����|[�U��F�n�]���`�i5[=��v�1��;�%<�q��
��ƷtC�ċ��tL�S����B����8ݵ&페4pt��.��m���M���Y�7Wv�Ռ�;����X�v��J�Y[/x7t��Ԅ��\�p�Gg�Wsn4�m�c���ݽ.ζ,��v���n"뼵us:�8�������y�*�m�c���Ǘ��+8s��X�Rnˮ-jy��W��ClۇT�m�ϩ�[�Iэ��m�=q�#v�k��K�휃��-��aPU�g��v:�i�N�r/Gc��x���6E�b^�v:�;K�p�Nu�{��8��t<;Q��Q{f�Dܚ'��16]'H��(�G��5pc`�(�n�:J����;�SF����qq���A� �i�"�=C��@�n�$��T�Me���;�ż��1�#����+c�2��R����;]�6��66n�F�^��ȝ�x=�g���M��8:U�λ)v�պ�q�wm:�ܨs���iݡY9{&�t���Ӷ#k`�<�{;C���z�L�s�m��G�n:U�+�7<v�`yxݣ1�������H..%`;ps�:������ �rv�t�6�P�����R��گOn��øv��[�N�ޘuO9�܊����&�7jiI4�׶+d��������X�Ʈ�[8��.Q��v|���A\F7E�{�@d�ޜ���\%V^y�l�N��N��"�s�F��i�>R�U��$�i�zz{W�������+Z�n�H3O\��fຎ�P4���K�[�+�����e��8�� -�UUUUUVt�1�3�5T͌�;���G�p�y�n��g�Qv�c���]f��u�+��ӷ�4+�խ��Y�������㛟l�pX����a��\N��=�,kh�D��ū�k��+�gFM���ڕ+�lo�v^�����;���5�=b�݌�ֺX;>�g��dF�=kS����.tǓkD^m���Ў��b3u�ǫ������k����5ɴ0���������Sדh�=�quؼ]�����7��Ĝ�9${v�����.�lՃ;Q�.���zN�\]�n��N��l]ev��G�<*ՁΎ�R33��]���®�y���sg�e�t�/]5ss�c+ϑu��c��ݻ�[v	�8���i�۠ؓ;<ќ�X�Äz����֝��N�S���Yk$���$ ��vU&�R,ÌR�+"�F1BT����,H�`���C���np�`J��T�R
T���Za��)*
C$��a�T��ӖT����Xa�e�8,V""DI�E*RVa"�jg8��Y&1fd�+"�0�dˌe�d
)X%E� ��$��T��
E�-+ �E&Ra�bE�$�Tf�(��"�-���J����Ȁ�0�����J�J�a*T�-�U@�	B"(T��E�bHe�B((G�a`��HT �,Z�"� �

H(H�dU�a*B�*�� ��2��H�VAa �T2V,�H(*).�����dwkS�8J�dbJRVM.ӷV�ޣ9Jgr+Ikg��]���Y;�ݰ�O=)�gZ��r7�N~r��K#�QF�#X (�D�
75�v�nu���X�=rm<c=�S�n�q@cg�+Xw��7�]v���n���r�]ۑ.�%1�k��9�<\���!�uu�cWJm���r�*��nɮ��G7k�]ql�H��Inɩݺ$�^��g N�p�ŀ�ook�{[v�;��.C�aؖ��ln{b9�j6�uv��N����.�k�U]��89���wQv����W��۱�cC��;!qs8-��1
��N���o�k��؉s��p���hc�7 	��N,{A��v�w���-���T�WF�;�����r:��ڛ��'X���]7;�����¦nw��:�g����ٶ���p��ʻ���̧k���k����ݷV睸�FP���V���j���Onn1��^�X���da��8n�Ů�;`a�9�0q�^/)�v����q\q��]� j�q��o�^���w>uى��u���ʇ1����-�]���z1��/��]��5���(�=�4<:Gf�\ջm��n|Jݎ��E�>�rv۷ώ-s�x��m�m�Z;T��x7�mz�ۭ��s���Q�q��c��M�c���ی�ܴS�z�Q�u�ٶ>N� 2Y㢷U��&5v�v6�.ӌݺ�g��^w��GX�]r�9U�\dl`7�;��jq��]c@�6�Ƽi^_l՞�ۮ�������k#&8��v�k���Z�J檸�]&��ݗ.qc"[�������><\n�K�Ϩ74[;����p;ŕ�N8�N�Kմ)U�zӤ��y���N%l4�W�����{ќX��ni���."�ԭl��	�F����6�"F�A�����;���{re��"���{e8�;�3��g<��o' �GA'���"����n�cl�������rl(��O�"g�cd��0�ݹq��{��ȣ�7�����7g�����{�^��;�ay}��a�۲�b�"���Z/����))S$V�/�}��[�t��7OTQ �L���֟��w�o[緦����1`+qA�ҫdz���x>l�l�o=+u�m� ߕ��D���,d�'L�oV^�oz�۾����RI`Z=6�x�����A��w�R�{���� �zf@-��tQ�"�����/}���{OY��8���Ո�h�&Ō�D�>�5�h�{�7��6��=�J�]���AA�M]<��I$�=�s�Lc�0#8n|I8�Q&���&����#�&Wt�����n˨��݇V�[qu\��䵹ږ<G0�b2%^�y=K[�h��x5�p@����&�$�]�~���3�fkω��!���ޮ��G;�rʙ"�����{P�'�{�
}��I��[J�fr�b�m˝:dH�� Ō���gT���ݪ4~���ϱA留z��jTue�J����Y��~$�d���tI�<��$wF���i\�zW����I��Y���I?���*D��R�����I�O����$�h���WY����z���}�E,7�� �=��c;�́	4U��v�ѤA�N��;tB�;�e�R
[ut�{�o{ ot�TjG�^�����I'=��!��<bXU������Mg�U�Q+%��!ŭ�����9c5�؃ YCWC�k:��~�]���W���i�j6۞�y��6d��D�F�g��N�ַ5�TI$���t�Bx�$�kv��]L̘߽W��DO+ۣ�;�I&�?gw�ITH���� @���:��ǉF��}b�򁻬�N���HI&��{� ��Y��ܭ��������Z�h���7ا���7-y��جwf�T�SK}3$�%��=C2��K'U�VNGGs�cWm�~���&�N�IU$���z���&X�J�Ʉ�9�=S3E�M�<n�5y��	 ����I������/k�o��ֹ�1�}	$��y���� ��V;��z�����n~�|f�k��������^�]/~�`�cv�p�1K��a�փ/D݃:�t��LP����>�[d��������� Ü����+o2�</�4�Q�󑁰��^o^u���89i��=����'�g9�_��*�4I$���D� ����h^d��u��i�7h
�ˤ32`x��=  ~��|�b���7� ���h�O����(ө��`�A�y�On��zw�m��}�*�6��e�>�gw�ހE�}���9:���
R�m"]X�7$=<�R����;�ui!^�)$t��ٝ���9��)�M-]Ϊ�U�_j�ϝ6r? �w�>��h��c�:���G|L�s�\�vhچ��Oe�`���Q���Q'�m�v�5D���9�:��g�%�eP�z��)�S)��&T6�gF��:����G�%b
䃱Ki��?y�B+!h��ߥ��;��H /���{�#��~��/�f\�ަ�T�}��J�Kn������ծ_c�\��ܗ` >��Gn� ��{��%�������m]zߧ��[���l#�Zj����֨| g��ʄM�R���^���M�z)��﻽�����vG`
�������)f� =����@_{���oh3��TN���D�π]��jh0Z�6���wYx��}$�	�����=���;�Dqԯ~$���UB	$��Z�\���{n�K�hJ�cS:7���kR7\�d�Ή�i��,̸݊��Y�$��G�B�0�K���s��UCd��ݬl�w�O�i�3�T8�j��D���<�ٟd1Ϲ�{�'+mu�u�����k���k�5�Rg=�2vˮ���tpN�;s]���C㴽q�㭦��o^k����w�@P�`��͓d*�xqm�6ܜ[��j��O6:�f+��v��Nۧ�\��NA����T���R��q6��6�b����^�W�nۮ�=���jW!�)n�\1oN��Z�smZ���\<��a6�~�uL�I�T��ĢI#7׈�U߃`�#pɮ�v����i�c���)h�w�J���Ω�I��, q&���|I$���T�>qk�6N���f^/�T�ݮЕ8Kn��{�oil�y�pa#C��z^]�����}������(�)��)�ɥ>��F��N��o�%?Mr�4I�p�� �4Ͻ[/�����4_��$<+H��X&�	I�N����$�؝#wEW�n� _������3 ����_}�sӾ���|�o�=ȫ���A���e����eC��a���n�\l�����\i���7g��g��QyU�Ė{��&X��ީ-͵�o{�:s�x�*1uʢR�����85����2�����n�֓������4m���NݨU��]��0�v�؆�7�r^�G��:����j^~4�;xՋ�֮{�����9�1�G���&Y��;�V;�vv�6�-��	GKeoZA���o���W��������l�s{Hgzf@-��[�i^4�*�n�߽��[,��.�� )��f�{z�@ {�wz�}ћ�xw�1�3�`-wY��Wu����7T�$�w9
]��׆���D����D�MW��x�I��{�$*��W�����߬�S�H�3���zn�b� q��w;��נ�[�9p��ulO�U�����Z_ }�Ӥ@$����@m��p�/��UHb��{z������$E�ώ{7��@>f�xT���~�%#��6��I��9P��h
>FR'&QU�_Ʃdz|��P@ ����6����'�w�.}����5��E����*�<���j�/I���3�㉿�OYggx�hb��1sm��_����v�������-����6�%moZA�x�˯3�� �{5A ����Z��<��E��I�������}��7��R�%�WD����� )Η���警@?rỳ�b�t��D���z��bޗa1���HWȔIe��'��h���K�țx.�:h�D�QK�m�OXG ����_7dO�w6 ����H�Gv��kb�z��b�t��J}�p� ��Z�%��M��3�ַ��'d�&�5^]�$$�|R �#�q����po�ǯ>�Ӳ��-��n��-�N�&�y������|�� s�����|Y���j3��6����G=��n�C�q�[�$�Ot���OĒMV^��D��4���9����ۃ K}�N���D�:�uW\5�|(�X�M��8\څ�<G�Xv"�j=Û����>�ɚ6���X
L��d���>�D�N�\N��A�'�Z�e��J$�0��?i��2�%uov+{��q^5'T��Q�lr�@�,RB�����#��;�h��:_�pr�d����a-���w�oO �qL kݻѤ�_o���=��cl�s�}���5yl�IWuY���쁒?�E�6B�E�4I���_�� 2D��{]�����=��EJ��a��32`{�y�� $�5�46w������1`��۽�֎uJ'c��-֑����p�ϕ�0�,�Uh����e�@�{�����v8�G'�bX�����/.�g�m�V@W��UC��-+O����%ߴ�D��5Ӳ2�O_�3~�OWO=��yR�
՞��������y�jӳ�f�2��'-A�е�\�_���������5�Z6�������t��a�8�Q��,j�Mq��G�R����|W��ƥ�f�&�.�='�h-��<�]�N��b��l��ј�a�6����v�imW:�2��p��]��V�aN.tq<,��%5�k���2x'B�r�㛫�)�uƜg�i:N���܏-�����;��������v`L�Y�/�Y���[��ܼ��'h��4���p�X��)�n��:�Yd*Ž��������!�d� �7�'d�I5��l���N�-P��6j�vo�`π�}w�@|��++&�1�7��Bm�j�]�k;��uhI��nF@d�]�l	D��N=����2�G#	\��Ľ������{� !>�=;��ֽ�sh�D����9�>��P�-2x�=�Gv=��H�X��W'X@ ���! �|s*˗�������~n�h�{�(����O��k\�|�0�Lԁt��F�`�N�q[$�N{��*H���uz�o�ń��dn�����v6Y���밶���,!U�Pn���h��(ڱ� ~��:����{��IW�)}�G>mp�%�v�$�9=��:t�څ��moZ�!�g� Skrmr\��Ne��M�7��6�����9{�cy��fy���^ͭ�7h�-˂�I����[�J��-����K�MI?d�t��4HG|R �92i�8�\��"�Xx��%�+�����  Ý�0����V{|�@ �����f�z���6�)�ʷ"��6����=��۲�6{�� 
�� 1ދ8f?yH���2�$��s������F&�h���[���|~��X.ڱ�Ȑ]ｽ��2w�,�O��]ݨ�f�l^7��3���F��m�<o8j���&���V�6��M������~}�����=��!$�%yU�ı�E�yGƇI�QQ��BĄ}�:�������ޙ�kn�4N�b�L4��GК$�IW�)|H��G�:'�V�Fx��%{����S#-QKkx�w��|~��ۃp�`t��l��ߍf|za:�]]罉�/Y�O/H�d�5tVk��i�Ƣ�$���T��35Q�ˡ�tj�h���o���;�oNؤE�M.�-j=��sD�W���f ���Ƹ�߈:��w�N�%f.�u�i%���\��Lwy�uS]���a�'A�/)��p��ϵ^�N��hgW=��$E�V�T�#���z�����;�o���C�����=��G1��O^�,��7ӊv�*�Qj�lS=�Ugp���P�/��ZC����u�� /Su������PRAR�1��^ڲؾ�>����ҭy];77��s��V��nv�o:�
X�} yʇ>�L����ܹ�N��=m��kf3�R�H��R9��E�;fZ����:%e�_)���dW wMVF�i:z+H5v�ˮy�������(�ᨪ'�l(�)�A�OR�]�v�ͻ�)�O�b�Ǉ�G���vˈ'%)��X'���f^* X�z\˲���n�0��>U�F��]$�r��r�X�j3��@i�Jܭ���trG+�^$����u���=ҵ�Kq��{�|�NK0�MYǗM������/GhW*�6t�#��J��9�siuW&�RI�Z��J�2���Ɯ�5�	z����dnDre����Yge�n�I�ڸfǗ�j�g+)�ÎU��Wmq���n�(�w÷�G>��N��d���&�qX
���U	b� :�TY
,X���U� �`&V-� ���"�����`��$"��B,"��AdX�"�+	P
���PPDXT�AAaY	X�*�H�@X,"�U�*$XE����B��R����sa+"�d(�

��X#H�
EXE��� �B��"DA,X
)�P�`��R
AVDH �
F ����$AbȱAA�#�,�,
ʄ��E �H�@X��@X�`"

��
)"��H

�Rp�9�s�����V���ޮ�zo<�
T�m��E���y�s�ߦ�N�C� �5hI�3����I~��N̤V
G%���L�f���Ɲ��89\��#��֒ %~��!ճ���2лe��Ā|}��� ]��!�j��9
�h9w����������-Kl˶˭nuk���s�#.�~}}{�Su7%����|��߷�X k�{���~Xmq��p�&�� p�����Z}�쐀��~�eUܳ<^TH���~$�}�I�-f����s/'0b�׊6���֑׾�Z� �}�ml A���V��z�?{���h�GϽ�CΝe^�-R;ky�s��}l�vi�3M�Eju���{��$����}՗�	'|�ɦY��kU�n#�b�w��L���noBw�.�(},��i�N��-Gs�r�g�k�W��?~�����hy�[+��۫�_ߵ�@$��¥��u�6�]�9��+6�koo;���IB���Z����Ӗ���U�Gn펀:P^+��Z�]){��OX89\�=����#s��� �Kng��p�qs���gu��n���]Rt�7�%n��b�i�{=@}� ����������E��~�����Yf��QE��wb�B��LA8�������5n�w����Y%g�$t�h�N�*j���v�_�{d���r�	+"�o��v���vu��U6-�l��l��ݷ���txg��4'��� ���O�&��cœW��޹i��8���+�,�P0������֣8��B���R�a,JѭƔ�]rݳE.��um�m��?��N��D�{(&v�n;
��<p�V�Ol�a�<[��aШSf�i筻]v��9�1��9wW<�Q]C����l�1�]��wb�.�WlМp���۶�G]���4ln�]��\�oDc��Pq�ƲZv�\�9�;<��A׋��ڻX���%�#���[&n.;\�z��F.�qs���-�n���9:�h1��g&���&lq��*'\,����G�:݊�Ko2{m+  U�n�{y����b�������� ��a缺eQNJ
eU�v��)�y����|�]eO{W���Eە�m�Λ���s&�2]t���� d��A}ϗt����~�}���� �o{���~�Ks$���F��Z��R�߹>����` �sy�	��O<��:�Uͦ��Ѥ�����۾�@�m����'x���8�繙 ��yw}���gn���ɧ�}��D�V�:��\��ֻv�u�f��ha^1L�_���}�;W(�B�kh�=�r����o|y�+����CϺ&L�]�ew��������^�H�j��X_jβ��qb��;��r�Y����+���jr-S%N�������˃�S���5�}b��������¥@#�o��!��{�׬����Z�
I�]}�	{g]�I�|�Kv���s���6 �yRy�f��hU�o���F�
��H9{�`=����U���#َ���́�1��A����m�暺LJO�]g�H�xO��v��+6��w|���s��̈)�!������]\��awJR�U��s:v��*����˨SD��5]�s� I�ް,y0MQ�5J������X�5�QA�Zd�<�rܚoz<�v�y�p������+6����������79�79%�ct�j�x���Z U�i���Z��v^c��uט�SԘ�� �����!B
�u�yz¢>˞6���9������ɾr���=3����!F�o7� �o߳M���+̝ݥk�)&w�;�)�>Z��y����d/�L\��_j
��C����X�#�UƚuB�N�a7��{l/��{6FM4�y�� ��{��f]O��G]9�-�eI�r�E��v�\�A˴�h#p���F������ߍ���7�o��_��{���]s�Z�O,��iZ+�rZ��}5P��n��y�t���.z|�d��P�H��� [�o3Y�UQ�w������*��N��0�$���� ��㧴O>�u0���
���n����i?�M<���<��� �2�I��n}��������k0l�q�`���=�p�_�OĹ¢��+#�F[�u7@���S8�WGzh�YPmb��K/)l�<�5�v��ן#�$�8�ήE��><�.P�2�ߟ�t_�9ܹ� FO2p
��F���y"G��+�,����7��1���#	Uq�ZP��"rdݸ;b8���k��-֑ Xo&�W���
:W�x��@���x�]�m���N�X�5�Є���3	U�j�*h�A�S�E��h�-ze��t>�n��
���@y85��RaT;3��*�˳�S�^mР9��P*:�V|] lݍ�B����KR�R-'I�	���W�I��|w�0> }ʐA�����a��9Z�e;W}�N��p��6�x<���l�k%tn6�<��m�� �_��g=O㼝�F��Qп��I4��q3`�G�4��Ԩ.܅�q��7QٕJ��@)��G�i�0�ʈH:~�>�流ؿm?3r�Gs#2@�b�N&#aN�̯�[�Ƕ1�=���֘Ҭ����s�=�m�l�;;a�X��u۳��!��X�H������>^ۏ/m7��zw�#�=���ps�t��s&����1��Y;VێI��v�ݞ϶�58�.����NzKx�ml;k�����g:���z!|��`���c����;O\�5gO(�LTQ� �;]��E
�������(���s�5��si�ׅ���-�^�t7=�0���X��z�SM�e�Z���������o*�*/v ��W����{3��T�*)SN��*u�$ٞaH��u�z.�A;~۴@+��`�[9�MR�tS�̍��a�d�U� ��뿬�A7]��#����ܹxc�7\����q��y�I����B��蘘{������ެH .we���y��ius{�B��W⦬�v9*+
�_������;�R�A�7�q6�}}}c�GNi�t���[�s��7wy�9�y~F��梥�Fx��V��#0�w�]�J���D�#U3�!�٘f�V<=[��]�
�&2��:_��4�]B���7���S�6ڙ�� '.��p�����Is]o߃LM=yfyϏz��z䦽����9k�T���"iӚ���`��x�5f���b/92~3��$���J�tlV�ܧbd���� 
�tl
�޳�"�w��tj�6{�)|�M,�{w����]�<��S2��x^��}��u��9i�^קV�)$��Ս�],���e��B6s�aJڎ�*t5h�����;p�%�G�kA�}��.��pi3�v���77ۘHwW^4٧�i���󀢆��r�ā^﹘��m�AǛ5'�3ء/mRtRO�M%a)��$���vA$sr�{����a\�OVW1��v<y�s�7\��f'�m�\��΢��N^2����^����t�#cM���[�9�u��%�"��/���y� _{���h���`���>������f^ϻ�=�=x �=���Y꤆���j��k礅�}��{E4M*i�e����H(o�"�]mPI��N����5����z�X��M��S-����ۣ�JTB�%m�f�$�tD�*�GA�Q�u��*��UNk6;��� +��b ���hݸ�]�u�M{���A^��,���WԉlӒ�$���|�\N��������@e��A�{|�޾^�.��R7C�uK��OW���A�gr^v���7�b��s^�7{4�J;-h�H�_�L�o�{��E��qpV��w}��}�V�RJ��z��yۯR��m/zػ��q�-uꏂŽN��Jzg���{�1��O��nu�N��uf����G��2���_�С%������?f����X*��־h啯�����s:��+���A��`���ù�s�׵�<�����),�Il"���t]B�$8�|�[.55-��HUw����2QWj�����x~j��n�#�x���NL���9/����f%A�0���z�f|G��L�}���HP q�8 ���:L�W��mo���WfbX6S�Ε�����o>$ۜ�JTh��H�'�e?W�w�3;wj��uK��O0��P9�@��n�H��s+}��5h�S�s"��Ӝ���J���Y w�η�ezu�ke,�A�V?a���L�	�&@W����_/�v��1m��`-2��I�:vgq���7)�P�ܲ	Y0<7�9��/�^^U|Z<��ۮ���LM�����&�iqr%ޕ����AV���cAqub��W|�+�F?��*�ڶ�\K���g�j��K\�or���w�*ǐ�;�c�ZE�gMa��z�v�1[�w�,��T�����V���/8e�d:sB�.��e*g�!YOt�]x��M^�*6��r���uԕa��������%�o���nL_��X�ã9g{1�@v�b_��N��Et5��k�h��4W|��˯M���C�[��G�\o/b��ۋ"	�C/��ej�r�`��#��K���GeS��:�b�U�&���Pn�����o	GUh�0-$��g=��8�vY9t9�0%*C�3�ht.0���lF�	ďE�r5�v)��.�i�jt��+Tù�!2q�6S�l�K��!��ǚ�2��ܮ/�����I��޽�5ڡb�I�#�Ų�t�ڌR�לu��֥�w Cq��r腇��Ie�diԦ$7>�{ik�`ݺC�u3A�e����p�h����XE^n��/��ϒ�����ɠwqti��ޮ[+��k��a�e�-�VM#;�;���-��ۮws�$�/�/��࿡a�'+�y
�ԡuB�Y{+U��_K06,�F�;�������fv�E���
@YaEX��H)��YdU��,X�R,���(("��H��H��������@Y`,��$XE����BT
�Y)R�+Q�
��10���X�@X�l�*��l+k��V�T��Adjʂ #+"�TRE*+	*IY�(�`���
L$*A�#i
�T������d���(�[b��k%E���,��+�Z�V�TR���<��۞y���c:����^���h#c�&�5/���n�՜s3�{v�1�]n1�\v8��vo6!З==���[=q��:#�7*���mp��j�{m���8槜�0�D
�m�2����{]�q����ṁWm���:��#l���5���kp]C���8-FdvU3��[��\r�X����3�%�\�\ s�7+���g����Vzت�t��X�hv܆�6��]��v�t����f����$���W���Sj�/;�yi���p��S�͇;�H��NG$☮�Ƭ��q�۝7G���gq!mI�.E4m����yx���n����m�G�l��.��6+=y�-��uۭ�fw�q�L����vr�X��NE����Z���N��n��۴py�:u����ƺ��ۊ��<I�2m�)�Z�ۗ2�烐�ɰ�.���)}�,N�\��oQm'l�v`4i���e� ����X�����u�{��'��ٰ�m�;q�W�:tpx��ܵ�X��ɞ�ܧ.��7v�fM�u��m�V���x-ۋ�q��0[p��ٶ'�f�9NJ�V���^w\���F:f�	w:�F�j�$��u�Yɑư������X�.{p�J/7>slƈ�a����I�1�`����=G�-�o]�;[�RZ��{nq�q�q�N����p񀱲�^=��alWh��h��mr'j��L;�r�7<�y��*��+��k��	�6�����{u&�w��u��r�<Y��n�� ���)�-�ս�<�&<�k�9vۮ��h�q�k�yMv:έN`��v��3Pj�]uX=c6����n����.��:�s�3lp��pG(Źy�
X�N]���k�u���g[og\�+�=�t�Hs�G����{������n����鍎���9<��˹��5� Mw���x�>q�37N�:�mW����Ӷ��jػ��|�`2�3�4�]�鱞,��o%N�=�cGi���]��.Jmգ�F1׃cI�Ʀn]�dzeSd�7�Ƥ��c�1���8������S=�հY��\�)��8��g�����qq�9�S�����[�l�T��wk���)(.S�e�u�T�x�a2�X{]�~�����*����L�h�Ͼ�9���@����W[���h��_�`�?wL2.��*�i�e�;뻲�َZ����wޭ��� ]����}ݞG{�/��眽Ն:ϫ>a������\��$���C��n�hk�����=����{.:�l�1)��rZ'���VTeP"����
���YZQ]�Wc�u ���� ��]Mu���ۧ��5��
����}����^ ���Ⲵh�m]�7Q�ew�R�u@�t��A�H0���nqBU�レr�;�=]���������ǖ뒥��� ��\Y"��f���/syk��^z��ȥRɜ|��z�1�,�����O���d��˞�y��x��{�uJ�ix��a|5����-d�"�Ny�*���o��?����
���o���ZY_����e̠f�s�����HI�A��F��`B+���r���k'y<���}b�%b�	,�D0��Ref?LοS��o����_�F w����˓����ɧG	�M6S��r$/}��R�%ҹ���݋���A�==���=���ms�� ��+���j5a<5�&��� l�ņ1A:�ZR�+z�!;k��e��d�v�FvZ ����F�W�����I�~�b�
�������b�m%^��{3���;=���X��9)�w{��:���~��I�y7%�E(���if!v�4-�7�� <�b=��N���J��;4;��ɺ�Ą�+�3T�X�8��B��rOk����^$�fO�y��1��~�Q�'����~�`�?���NE�@��Tnϥ��v�l��3��`�2N��A>����,o���+}�`��DFg�s3`�u9;���k��������d7;��y��^���e��+�"�#RR;m$;j_]b�z�t&5��΢�x����������P؃=Z��ܼ@�6��`.��e�V��۽���X��^�H��X0��b�����[O�A���~>}���*��f���[�CC�ɯl�E�����0���	�R���L�'ݽ����<��g�Yڂ�t�a6���r�f�Hv|I�_z�	��w�*���-
�=�M���{��6}a��%�>7�K5�н�����K�s�ey�&��y�~��w>l��Wì]r�u���?�����ӳ7���B�&�[��]زB?�5�;�3�GzVQ*�w0	���qbi��;�7百f�s�yl��k]�ݞFK����6ܔ�J�V'R�vK�
꒣�~�}*�M:�n��3 B:��d
��s��N�嗸3�F��G9� �6S�`�|��T���o�� ��a�T���i2���Φ���I'a\�֊�۲w�����u�V�9�A��]��y,�a:KcR6ꨝ�oϽ2;v����R g���{��U~�E���&f��~ê
i�T�mfS�Oý�����7N�� �v�7���
��7/�s��k�N'�:Ֆʚd7�;#k-����x�l�hp�޺�5�H�)ۼ��7N<�4d���Q��w6��*U��e����s��Q
�H_��qg&5�۰;϶ys��5Ƚw=����>Q]����I�;�*\kv�c�n���n��w���۳�c�q��9Ļm�D�F�΢td�-�b1(���v��3�ׯ;A�۶�{\i�y;e`^�Gkj����<x���p�B�<M�TӴ���˞��!��e6�sk[j���m=�7N�]g2;��;u�h�F�8�<�-h�K�������sgtR��ZG��;��3qOr�᷽�,	dL��u�2�k�E:��-���)��ɋ���ā+ܦ۾�b[�´>����~ڽ�`kj��e9 ���3}��,�/�Y�^�$u�ki�;�Si7���־oy�	!�+T�f����b�f�r����{�6�A�����C
]���2C�:56X��IX�~��I>s���w�f�	/�23;�x	$�����{9�dm�RA��A�ۖ����v	1.�7��*�)EQR�U[���-�M��M�'�M�$�ϽaR�������yy�#�&�����RA�n����R������ hIn��Z����
W��!"� �j����ѫ�œ*+}HE��*,өEV�B����B$Bo&lHj�]�������調g/� G~�ܼ@|��V���d�u�^&	5�;H5�V`��3$�����,��2�遹��� <�����h��a��T�-��L�`��3���zՄ�U�[Ÿ��.w��'�n���b�%R��.�Y���v,�<Ü�2���|�Xk�j��M��^滬�k�_ώ4"F;Z�9 ��>V۲W����9��{���TV�FU/5��Z��I�ۘ���Z�
�i�7<�N�o�}������.��]��MU6��K@g����ܳ���אsv��i���_$6}/_�[��ZТ��O�[��XEw\1!o/ܰ�`��z[b]Zv�܆��KꚊ�՝DI�%rKݖhs�Gq���`9 ���;�7��&{�:���J!D|��]߭+D����)�,'U���S}�]V��J�+��B����{ޏ���s�u�#7������67'!o�{����o�.�w����e�$�{�����n[��1�B*�h�i���y�W;�_�|�>��I`[A~��Z�n���	��E4��:�v �j��}��d����K|y�o14ڧ6)��x-�l�j�oو�E�9~�W��:���m�3�k(�z?������)����ˑ=[�)���iV�OM��~���u���fq����<��D�{sw,o�DS���w]�u�YH7�1 fsy� ���\ڂ��h��xo�X[���,XwoX�p����o�1꫕٭��/�9�fN7M�5�WO;�W=�v�ߡB�QQ����$h_�����V~���BAS�_�L4{u���$�& ��&}�{��=�����:���!�ZW����yT�7]�lH,Ӻ4kc�R�Ud*��<߾�uZ��]�L�o}��I%{�v��N�~��S�I9Ӧa;v*�^h�E�K0]�=��ײ�خ׼ �wI�	{��g��3^����#Y NqV�H��J��	��R3W��;f�$�.oL� ��;�eDct��t[Y�1�מ��jfcd�e����Rz�H�{#gk;{���y���B��u�y�.e�Ý�L6§|��6��R.��C2Ƀ8�����{� x%@���Θ5�Z�S=��@���B��_�갨}TEw����9�W!-1%�+v��#��_?�e�l��#ty��ղ�l�WV�O����L�@��n�X��r�
ڿ�������������ۧ&ۗs��̛U<�_]�vq.S�9�GZ�vݷ5�c#p'k��F�仅�ͱUz�5�=,vP��I�c�-]����v;u���Ӽ��Tm���!m=�67lH[�<���=�k{p����s�T���=t�q��G�h��*��W�����F[v礡s�>��Z�ۏ[zq�V4�q����s��Ϟ���c��IZ�w*#lms)l�w�~}}��8�tc6���O9����u+(�YY*g�s&ȓi�V�k��R
O:˓�aRy����'L�����'���b	.��FE*lnmI	a$#�敢�
fT/Wݚ���O�]�=��H) �Z��M�T��'��Ȳ"D�!D�K��o�x����Z(A��x��k�*hj��\D)=� i&����zי4�2Q��T���8�����|��Z����
ԅ�ל�@ٺA�!Z��\�2�S�`C�X�l���%�����O����yw����ν�C�+
0�)z׺�Xi�IA
��9�<��&7�5{��J߽ ��s�j:,R��Oʧ[����6t��5��5��t���Q.�~���Rqw�?Q�������J!)��YI6 VT�k��)	(��-��ָ(A$�~��ך��\~
�����C�x[�:��q���Ou'Y�٢�ښ�6��_����{��Թ�s�i�#
��{�lCi �}׹43L���@���gL���=�1��3�]�7i�]��7�AH,M#����!����샣j�CX$���-`�yG{�����1T�\�~#g�.�?s^�徵��wLy]}�X��ݺ�ۖKm�o*�:�]Yk�P�����u1���>���2�w�>�B�*Aaoz�P�0�*%N|{�掙:eH,��o���[�;s�j8,R������i���X��>�4:H[HR�9�=�F��+X�
�߇~cι�Z��m6�R��K�y�e�*IP�{�y�\ ����&��R�����\ S[�C�u�9���}'hT���zɡ�d��	P,��|�gL����-5�y�1�{�}����!X;�3�+��E���2�[uX�bK�w��^@�����T�<� i��x�z㾉��V_u�C,40�*�s�4m �N�T�=�I��@αӿ�:�����Ş�S�X���VYsvm�<�7:{O],�g�Qk|?'	��v�.�����s�R��!m �w�9捤���`T�����X$�Y/���['L��wz�6i��RTs�y�i�Z�>����Ý�L6§|��Ci��p^yz{_r�{��{ָ�dD�$IH�I{���6��jAHP��=�@ٺAH/:��}���p������(��3M~0f���`t�$����'H�2VQ�����6$�IXQ�`�[�����Y����ݣ���M�7�K��}ǐ1bٝ��1.b����<G+��ʙ3������l���-�:��_�i�����]ÍI��	jf�%ϯ4�7��yu��nZXJ���ǁ�v�v2�K���ds�=>�p�@�j�w^bH�A���"����*����`�[����&Q�Qq��cr-y�j������uѮ��Nq�C��;dB��Û����C���Vn�ʓ2%���+K� �&4��Э��u�{�.�nT{(���D��yyܯ��{ ��0:{֌�w{"Mq]�6ờw$X��ޑ�f+�7>�{X;����r ������1�s���޹ںjM���a�뒦ɣm �P�ݓhv��$¦�fV�t'X.�����;��r����CG#9��涞-[rQP����՗o9��{A)oʣ�0+�%;��j�k����%�:�՘u6�M\���Y�k6�Xyr:��lw}�[{�t�b��w���JȻ�r�tޣ�"X��r�h���]�U�Is��o��c&ݣV5�g~ӻ1�Gu���׎L寔��v�]�B_�Ot?z˻9bF(SY��}���6vEìH+tf��tT�iN]��u�&#{�ˀ�\��iud��A�g���Ѯ��Wβt�r쇓^:ۧ[�̽vy��x����XU�;a�����-j(
�h��*
�JȌ"��--�kTI+,XQ�E%J�F��Ҥ��`*1eV�+
�
�*�UJ�.)b
�B��m�)jJ�P(�X��IPiE
�l��lXT+R�j�P-�,"�j�dR
�*ZU�����X� �ʪ��+
�RT
���b�X,DX
���d�	R���J�[eE!X����@+*���J"�����R�6��L�a�hV�Z��Iu�̆|� �������GI�����"Ϸ�Q��%�/��j���RBX�!z_�!����ܿO=�BؙP�%__�Ѵ��0+X7��&����N��ff7˻�c]sÍ��4�#旳=�[-��˜����B�cP��¦3�d6��T+%ea�ך��dE�z��߯��%��)���b���,jB�o�s i �u����?DI��T������%�N�A�봋"��Qd��#oO&竢�u�Z���8���$���8� �pu��:H,钤�<�&�m
����azƹ�a��T���{����U�R$��}����"H�H�$���{̓bm|��K�T�09�4m ����H)��g��G@sy�7�!RX7�=�H)�
�'X�3dD�H�D��g�=�{����%[�;k�/��$+�z����qC�V(@���K�6��+%��<��M�A@�(���9����9[�%� P�g��@�AH.���a�Q�R�d�-�Rr
�9�Ip\B�Ͼ�	�߶|����f�*AMy���$�IXV�:Ƽ�0�R
M'�s�h钛���6W��V�_�),��?.��	~'o���ہ_���x$s���2s��?a�;�D�˲�Fǔ�0<�����5�X�w����|���$���v��T�����I�6�����q0���s�HK	!}/敡�(S2���wֳ��H���Õ��-�~�m�`T�k�t�h( VQ:ƻ�0�� �y�9捰�a�k<��3������&(j:�	j��`m�m̡\=�-��R�+���� ��O|��_��j_߲Ci(�d��:��&�2�R
%1�}��pP�y���޾-瘡r&W��d$��s�0à`T��3[�eL��$ňQ�^m��JH�DI��8�|��v}��}k�Q�S�!L�:��0�AI�*J	�9�4t���"%$G�;ߥ�y�^��+��Q�`���'�'X*�Cu��%�HU>���P�����y�}�i�
�����5�o�;O
�@���5���%Bĕ�}�6á�aOu�oY��1C�L��)��i^�>����԰Q�B�VV��0�AH(9����M`V���y�3�K�x޶kò
��-��
���N���>�0*v��5�{�O++%e*u�ɂ��������7��!4B��\0�C
�P9߾��l�2�X��F$\�~j2�J��u>�~�_4�2}<�Ý����+:ݚʟt���ؓ��3����f�sm�� �l��N�8,�t�9�G��$ �*�盛26���ڥpgmrc�ulZx��S�8�5۰�s�xV$�k@���iy5��&���"�W$�sI����� �V1X�陟�ʬnQ9�r"��7=��<�y��m��9�<�nnM�ۨ�O	�0��§m��b\ZP)M��A�s%���y��p�ն�Yx�n����lnn�Z�q��p5��F*���rs6���!.��>��v"
��sVr�uP����o���@c9sq��V�5�w<�hr���,�{߾h�E!Z0+X,:��M���[�w�5��3��A���
��%H(T7�~y��0�(w�f���q�rb�p�PaS��I6!Y;�N�<Ώw�N�{q�O�JʁD����l�R�-:��d��
A>��|i���oz?�:~���F�)�[���@Ǟ��O++%ed��y�M��IXV��1�z9��oϷ-�C=aRT*}��4m��VJʐS|��H��W�o�K���6t��5�/��\t�9�Z��o���ݤ-�y����HV�
�Jo���lRR(A�ʿ�*"��w�g���>V�p �臝y�4tá�aC����T��s0�p�AO=ֲ�����2��o�ȍ�>}e��#�JP�IN^}�\`t��H)�ý��)
ë���?��V��d���	&`~t���lu�^}��8�[�}n2���G[
�q�U!(WHT~]]���L;��r$�{֎��
�R
o�y�i6�IXV�:ƹ�a �}�\��w)c��+~���%���k�$E����7�9�4�����xr�1�7�+cXys̆��-�&}��-� H�ߔ��Tz�gwg�m�
����xp͖�
gI�@y����yQ�v����vcˋoY��|�	/�מ{��k���ߍ�؁R�VQ:��!���P�ιz-�߾�|�����<a$)�q�Ԏ�e���\!q�T����m �k��JʁD���>ˬ~���/�$P�B}�Id� Ґ�C�sӦJg~��.Z��۬I1`���m���?}:�mԮ��`y��ɨ0��w�d�FD�{ޠg�kX뾧02��7̓pM�k{�m�U�Y1i����S�������9�6�W:�x����@��`T��w�4�S`�YA9�bf�*IP�y�9掘t°�1����Zg�V�L���Tb��X�$��$�n ���ͷ����US�����8�r8��	�/m�K�IP��eaL�%��$�)����.�	!!�_����_k�(]-1�~d���؇��ӦKٓ~��&&f݁�t���}h�:@�����w����;����ߞ��4�Xx°�k���haR
J	�s�4t����YY��^u�q�{4��䝉�
_YՔ8&���8���B״��(@�K@�<���+c�`T׽>���I�X�>�����_�n-�Ĳj�s^��/��7z>��2]�Q�\�+�}19����4e��}U��N�*�E| T����<�+4�P�J�Ϗ�|Ѵ�ý�y�Թŷ&.5��aS/~i5{�ϭ�������R(A]|ճ	 �_:��l��jAHRӚ���k�g������h�^��¤Wv��&��7V�b�
����$T���S��ܛmq��y=�����M���+9��P�40�%�����$N�Y(ʞ��d�M�c���|�Y�iw���ak�u�����C�Ds��2r$��%,qEU�����uTB)d���ɿ�q��8� �-�y�w�}�h�����o~i+!%"|���RC[�³C%B�J��<�z:a�°�x�eSs.(w	�/�v��!,H���>��.��K�XS�E���$F�)�����MH)i��@�� ���v��z�3
�0*_�}<\d��ͻ��s>�֎��
��Yc%O5�2lI��+{��Y���Q�IA
��\�h铦VJ2E׿5��JT��YC��h��U ���C��X�c7}���ֺ�Z7��
�k��$�aֱ��(�s���56`,c>��.�{gv��v�\��9%,�{{�=�8��������*lrSe��gʏW6�'Sj�oJ���ߚn��>I�:C�T(��;�:a�aX_:��u��8m�n7�t¦sό��6��Y(�ë�2hfX�g��>�mzB���b�%�T���^� i �R�u�s0æh�l����X(�#m�\�u�� �뗤]��;qZ��;�=H+���N��y�A$���%ZJs>y�i�#%e*s^{�4��T�!Lr��D+D)M���{�>�R�S)�}�Z:d�eH,�eOu�d�h+����K�T�a	p�O��iPP��t��X8z�뻮����4o�B�0*AO<�2�h,@���7��D�<��Y��on����������
B��;eQ�7.�C�L��)5���m
�YXyw̚fY(2�X�=��'}�y�ׇLZ��R
y�y�7�A���C�k��0*Y�Wo����\9n����[Ѵ�똼�6Y�J�S�﬛�6�XV�;��¢��P�%��o�a\�.�:m�0��$P�}��V$�'�j����[vT�×�v�!ai���6�]gg��[�N����Js�w�6�R7�י����*{�|����z�M X=��{��wpŖo7$�SY><uq#��>ѓ�S�>jx�>�=���]7����poxN�O)�vf��en�l�5���1�J����qEcS�p�j��{u���v�W8�1�l��;<���t�w6x�]؅�GZ6u�LWO;�[]sA������X���ܭ��yុ8����ی��X&�y�YX8kU�H���aҷ-�N*�c��ᡶ'<g�蝸����9b�XE������j�:�u��W��3l[��;�ޓ��L�Wsm�)�;�X̊���'��[Щ�t�vס���[��>��2������j��2�J�d�+��ɦe����s�4m��5���=����C�i���@�n�iHV�{�{�a�`T��E���˦�LX��ݵ�B�%g^�����9�L���yHv$�+
k>j���Ib%�s�4t��$D�$���keMf�]���豤���㉞A~��im��#�Ը�d-�-�s����HT�����cZ���^Q�o��y
�YS�g�³L�
$��=�F�t°���t�ۜ�t*s������^��;���C��=�+&�T��N��l� �"�3+o�4�V�z���-���B1	y�p���Jz�;�SSCn��:{�w֎��
�2T��k�e`��O��̾w�R}�=�0P�c��¤�B��{�9排'L�������%�$�~���qN@�qO6wG6�'e�q��Y�rF��X��t��?_�㞡nL\���5��cY8H[HR�;���i�Z
���i7Ǿt^w�y���,N�ϙ�H(i%B�g����B\Kو��I.�tL�B��){�IX�����9��3�e�f��o/�iμ��tY���3Y�5����n��ዲ>[��ji����C�5�9�T�����h���,jB�Nkό����HW%�γs;�`�G��
"���������k �m&3���:@������&ěB��,aX;���q�/��f��
���Ib�y�4m �t2�VT����IL_��K�RK��pP��y��sԪ����E/�R^��ְP�����
��{��l@�P+*s�#��k>�7�� ��$J`I���
B��굷5B�7	���R/�x��, P����Ew�y�{�+��h�^�ם���R
B�Ou�f���u��0]0*y�w[����\��e��JUH',�	ES���\��:�7r�*x�摓Cu7�p�&�O�,�(��ygI ��<�ObM��a�6� �d)}u��sz�
(]����DqY(��YS��܁��u��pd�-ɉl�$%�������(R�T/4���Ɏ���ѿi
�[=׾�&�*T
ʝsz���������4t9��x�Xzs���[�9�-��:a�
��9��!���Xu��L���4���]S�˸O�]nC߭3b��pX%���j=��*�I���;G+u��B֋Y}S���C�ְ�o��M�������o\���>��_g�9 �>�->5�d����a��� P�]g�jkQ2�\�X�bJ~{��Y��T��[�䖑���%'�|�D�B��,V���0�(��/o��XD_�I=�O~�c�E�(@�7� X$��t�}D��D��X(A
kͥ�$P�eB���z�
vvS7����AN��I�H,���`�Q��RT=�h��
þzu�1�u��I���b�һHۊ!���Kh�GF�Ѳ���������5�e�U=���	�l�J~�V�M���D6��T�Þ�94��FT��O��}��%�HKܵ㸟��ء���7H4�+y���Jg����LJc6���&9����t�R=5��
sѷW���O��܁�7VaXS�oZ��L*K�,Ns����N�Y(���bs�g8����u�y�x	����"����C�-1��{-K���P9���}JB� ���=��y����o�4�D
�@�;�y�h*IP�{�=�GL:V�ͣ��; _-���!�}��{��Ͻo�]x�OFVs�ɦVJʁR�]�ߞl��X�i��@�y�_���5�}�^��silUE7����נ�{j׷,�Y2ᑡ�+�4�0���я%ҧ�E��Z�u��u��Ē���C��5�)W_�+S^S2���X�b�(���k���J��S�^{�i6����c��)��+�V�Y�T��߽�捲tʐY(ʜל�6�@����Y�u��;~�vݫL���6MsF�i�^��WA��nWO5�攏�u5Je�|�B_B����e�,���h�E!Z0+FK=�~���(�K�Q]T� ��/�[�,��P���y�{捰�aX{�u.q��q��n��aS�ky�m%)����4��=���V�DJ"D��@��|�͝0:k�!m=׼�� �B��w�y�y��
���8�1�1�]��t���}h�:++%e��<׼�CbJ+7����1���[�y�C
��RT�}�掙:ed�+%S���&�h��7��ŭT�b��H^6����/�6{�-b��iho���}�h0+X)޽��X,R(A����A_7��PВ�P�\�0�V��|N���1mơ�0���́��B��WIs�W{T��yw��bĔ�H��=�l��X�
Zw�=�H;	P��|�� ��j����;�2~�/(u�,���,ާ��y����N.���l��
ٷ+]M2G�Dv�ʘ�
��2�7�[E��\Kq.�-.�7�n�8-���L;de6{�?��ԅ�pŝʳ(S�s:��=���g!����Z!�Ut�U���˒9˻{2m�a�{��M_U�Nl�<]A+�������Ud�b� =�iorhA�DT��lD,�ga�pE����-�/P����E#�߃nG�[ɣ	����\-��K�{aP�9��{y���]
���J�$pV�^dt]l�t9k���\t����ݶ���������h���vJ�����}Ϊ�4������9r�f=�� �֭�	46�w4кi���曗�i���e��s}�Ѳb~ԕ��j�u�Rl�5��v��έ��P���T�mV���ݲ�5���|jG��p8�;�o���k�f�۱8���Ǘ7&Mi�u���r>�`��9x,-�6�Yx
ݥ{Պen�c�u3� �a8�Ӹh*,��+/�ɦ7�ks!|L8�{|D8����8��X�.�.��vJ��D�0.�+7���i4EaF����^�"a��_U�s��D.=x�g����]:�]�w|��j�fM�n�*(�M�֩����ے��˷�+	8�����&Z]�����U��yyF�Jλ��.Ǎ�g���r���!yǉ�ׯ��r͌���)P���(�8��L*ᠱ�
[�0���\R�,DR
T
��`��Fc��d�
�X���%�YP�V�R�±`�����Z��,�K�9�b�fqJŋ�U��8AB��ʊ
T��
Ũ(a0���G+X*�d�֌"ɖX�QT,DC.R�ED0����ܸ`�nL`a$�\%G.\,�ec["����J (�����0͞y��|<jL��	�eݞ��F=�<���t�j6�Z��t�F�'[��>��W��"`ɝ#�'=�{vN�i���_pmM���&����6��ښ��/�~�m˶��h�L1�[۴b��t7>6�7G�&�[����Հk6W/���bѻq�wv��g���äA�.6N:zX���x{4��n��3tM���U����5 ��HA��cs��m�/���;�������A�v�+ny�::tͼ��F/㎨��aks�$k���:�fi��m�������]�OB�u�a�W��*%�j�A� S���˹.:`���c�D(���VU" ��:b��f�q맞k�7D�Ylx�ܝ�V}����Pq�ݹ�q��3��r�����n�2c�u͜�;�3��Yw(϶^���i��3��Y�s�F#��=����8���<�vڵ�����%�W�0�t�iۇ�ۘ�۬\� �f�;(a�ZL���WnL���[�ex8�Ξ���psx�W
��;���s�g8�[�%1�|S�_3+�H��
q\�����]�#q �q�gv7]@���D]5Wc�m��⍽;���q��˚��]�F��<Vx3��ZW^�î�n=>=�����}��6c�T�\�!n�����7S�nSuǒ�N�.1k���j�8x�s�� �</Y^�γ��6����4��q��$żj���~$��X����kE<h�n׶�O/5�m���17���,G�k�]$©������c:N�us����F�[��9���ى��"�H�Ŵe�WUbw=�C�Ld�ͥ�g�{k\�λ{ ;n�r��JJ^�]�^�<5I�!�;#X��ڸ�M�u�"&M�d����i����w�b�?+�v�k�5	��z.�<�[<h
�����׍Ƹ{���^_qjz8�`|������q�#�u�筬����N�9�$l�=Aǎ��J-���#��NM[2r'a���M�bS��<"��(���+�.6!��	�s�:�;����^�I�x�	ۭC�L��mA���ࣵk7�]b��]�M����7oC�����q�s��\����C���?�{?�m�1O����c=s�:N�
�2VQ��5�6$�IR
g�kPXi�Iw������a�g{�F�;eH,��9�s$�Zi#?w�o��Ȃɥ��[L.ܷ�H�]P�$D�����ƾ���-��g��H-`T�́���+*g�k0Y�J�T7�=����3�|����}�eu�i��	���,60��5����K*Aa�9��Y(ʂ�)[y��n���z�ڸ(@���i�� l7H)���L
��fp*��MV 4�#�~��4�ۧ�^3������:ed�:���m&б%H,)�w�Aa��ID*=�h�'Z^����6�;d�2�VTƽ�I����`K�\�T�b��HZ�m+D�����|���R��M�f�� z�R�םh��*T
��{��f�J��*C���4tá�a��������|�g2���;�����{N�5�.��]���R�kz������,�O�/?���j���m�J2��^g&�+%��B�%��o�a	r	!'�/�g۸�Ƃ����yf���h!����H/��j�~P+�bJ�����Zkɤ�DI�T��"k�R�#�s|���ݖU͊�(j�F���~u=S- n��2��ػJ�W-��]��p�z9�F�v�d�s���Wo��Bo���(�)I
XVϟ�aR
J����N�$D�"H�ήW����X���#p���d�4�B����-��H?�t��I;b���d���wݎu��
�֚;��^{��.A��N��Gh����ٷ6�^jA|��� ���{Wݷ�mz�֍��W
MP�m^	�s0&>���er��}�ww����msNQ���5��xvڥ��AX�PMF�tQl3�9���yܧU)$N�k�\��FQ�[�6z�6�g��A>}�+yUc"��ͱ���>������穭r���5ъ�:7@P���
���L�5Zl�9}AQ^P)�Ҫ�넒|�;��\8�&#�ʡ�}X��+���u�9G��K:*��"*�P�K�����"���2���e����(�?{s�?�~�e��4bi�SK0�L�O��4�������B�۰
�p��|�cا*u�@NP�]�X��X=���T�`�qf�le��^�و��y�@�5�����]ϳ�ܔ���Z99��a�����:ю�YR���HJ
�(�q>��eT&�ܞ�ބ��` �֚2���e|�k� ���$��yٮ�M:4�j���Ov�	�zz����zo7�{_u�AY�4}yy�Fn����r��2�֜��,m��J�ͦ�e��g%�����q��pVkMv���S3Ln�v����v�1]��͵` V��${���]¼/o�0&'�e��d�!�{R�����=ܪ:���w\�̼I˳��A$�Z�z�64_�3�ם
v:#���A��߾_� �=v?��_UJ��\�d�I�A����%I�Y���κ��m݈U�4�>��3�Ce��<�m��¦�U���4�qL
Q�(�B�7<\�Wv�a�ZҴ����6����7B�5���ŀ��� K��fbW���d�ϟ"Ѓ_Zp�����#I���=��H1�Z����_X ;&}�;���<���#q�>�'H�RK���T��V�HD��Z���*W��	~a�A��ݘ2�${Q��RY��x��w�!''&	�sӳ �=�+7���n����a�5�]�*�L�����g��	>s�]�w���s��wns{�� ���.���Wb\���xy��qv�=3���"���{�1N�:ǋق�ŏ)����vo\M��w�˛s��"�F%-G�$P�O:�=�����Ж}�C]e��콶���7.��nsph���6�i$�n�/=���']��Q.sn8�]q�V]O��4�ɍ�w@��M����.M�=��ٽ%Y��Wj�m.x��W%�bݻ��X�I��a��a圜��\�g��lV�j{B�kh�Ć�D�u���ڕH{n�����2\�#
r&؛d	��X�9x����)5�s�T�m�t��Oē�z�c��VgF#�0	${zfa#�r��cI�E:V����V!�{��=� ��30�9�1`�ޗ�=�����eR����.��$}��ìt^�р�D�e� 9��FhTp��2�/��3е�>�b���<���@y��B�[W�6.T�S�>�����PZ�&�0o�K��y��y�=�F@)䍰*�7�mOn��;�����	�%��m��N7V�õn�0.��==>H���ZEJ+��*��^�s�@����}���A?,��+k�zc��s@1���ĄUB��X�J3E�X/fc�zu���ab�,b��b�J^��]�Ⳅn哭S�]3����o>/���W�b���5�Ea�=�|���~�`�>p��W6�@������	�T�1��"�!��]�`��'� �Ur�<��� F��բVkN'�&�%RuU5�6on�*�t���*�^�`	Wx�@
�o��v7q䲛�����!@��C�	�F��\X$�v��K����w���]�wp��� ���0���^�w�.?f)y�w�ѩ�i37�󓈾q鷫>�]]/Xt��C��'�m�MW>D׺�+'�J =������x��\RzϦ�� �ˈ~q��A��|��~�9�K�~G�u!@ư�tn�y��c]'�E�_!�ڭC���B�,�aM�G���	.j�X�Ox:�ۏL盼�J�qj��=;<��{<�^B�t��<9_
F�}��	&��C"�A�b[uk�Ӓ���_�9}�����Z _o��`ys��d�����\�㯞���5��6��aI�{o	���ީ+n,��A:;�j�PcT��UH�H��Y�]��H'�m�k9��F�q�{,h+��3 ?{3Ϟy��ŏ�~qP�!��Q�M�nӲGk�a͛sl�X�͊������0�\Վ4�Q���`| ��$l��U�`��y�|�fg���MV"}��،���`�(}�gy*��َ�S�c�tYP¯�E����ـ��}��S�W��U�.$��f@>��!��A�h�)��*����,��'ʾ [��@P=�؀τ�U�y�H��Ң��9y�:�[:��:3���M]\.ݵ+��N�f��*LM*n�s���<�?}�>���	������~����˘�7�~j��N��`K�����h�Z2�r��}�S�)m���Ej>�؉Tg��:���w/iz.P.j:�Gg5�瀎�S�&���w�k��k�vՐ!,u��Vn��1^����33#}��̥]l�M��mѳx�wSF�W{��yt����  ��v1֎	��nw��N����.�T}�m$�a�޸��z�D���{˜�YW����ݸ�#h��s�f�T7Cn�&���en$}w�A�&{]�Oѭ,H���)�B����bB�J~A�pۡ���H��K�N$w��y���!��� �6�N|(ow����g�%�nq�D���؍_M	T&�8�J��l�!���ҕYi�G�믏;�-�����1���{�;��Op��X	Е�Ͷ�v�N3���lΎ,I���i�@b.csmpr�����ݶ����ch^�صF���_h'�xGxܜt׍2]�.�ۮfy���N��k|/�ε��n���s�c�����R�r�-�"1�Y�:7����F�� �f��7j"m�5�GS�n�&�[���\:^9���僝��h{<�2��s�Ӭ��L�K�Y��R[(�R��u���-��)?��w1bh������
s6��^�+D콗W	�M�7G�N��6��0�'�>�b���$�P�A"wz`��_R��v�Տ��V�h����;P�o{��x�E��:���&�3�G]pho�{��!�5a*��T��)w�wg>�^�� ʟ5 ��{������vg�j��b^.�*�n��\��b+�����{�{wh�C�g�&ɘH"?y���7�N���R"ZJ�U#D�&4��f$ l�D��^81(Gju�[���ώ�j��~L�Z�A��{y���w�J}��f���`�Nl�0��N5U�M��N��^�b���[Ŧ�zeC�W}Lj�x�F7gf�<˅�Qv���:���Q^�ĊlD�h�J�mn���U}&�����H3����V����G.��ST�4�Vl�.�!��  ��S�:,F����B;��|*}�&ۢU6�V����/�.9Z��|���� w��>�ПV��)-^o�(�PuwБZMi?K덽h���\�S�\�( 9��h�Z-]�����)��Ƀkc���h��v�t�N󳝗��s%�kN[�������M&::�ͽŀss��eh��S�'	����,�����j��I�.Q.j�M�_m��&�w�c~�D��`�Hkł1˭o����H�M�U*�I��Z�K�>���*�?���2W�,9�)��J�Q�t���S-r\Z�����q�u0vS��-�*����[��+N�I������r�G#;�i�yX�֣��ַ�����V�-�φRUzb�a��ɜGyR�R�ub���ż\������eT�Ȯ�}{��!�
)2�s�P���A�ǗaȤu��}���n�KK˺�0�%�ʽ�������:s�'38
֍4��Lv[WHf�Oo'.��!�Q���:y,���ΏN��g�E���(.קkx5K뗕7u��L��ϫ�u�MށB�q�n�v���jgv:���bI�N��)�GϚ<��C:ڰ*fK}3��MBb� e�˷��0���[yD ����FؾQ����_.8���raɕ2.��vnѫHjؐ6���M$��ڇ2����.�Yy�՜��wYQ��Q[�1
`R�:��t�V��.Ei[CZ�7i���A劙`��/�LW]�@�k�W��2b.��M�c��7�6�vs�X�=5n-'�G�M��)rS�-�Igue#�R��X�):k�ɮo�{��y�*F%��Ie#���yWm�5��}� gn���c��Y�
b�r����T�-��w�R�.�J�`�`ѩ������sm��R��Yʕl-��î�A���������>�OAm&�[J�~Z�U��ggv�k�RݼB���,�b��[b�q��t>$�U���TP-�kH�sJ�ڥ�,+-�.��Щs�%��jJ�Q�
�����\Z����e��g�����[l�1��- ���0���q�A�Qچq�p�X�.
�B�p�J���eq����m��v8<y�=������n(�L51K%�-*e� �%AG4P+&+F����KJE08C�V���(�V6Z�ql+
2�\)R�U�r���cp�c��� y�U[�"�����Q�*.6ڭq�B�U��Q�	�`�aX�¦qE���1�U��Y��"��R�
���QG�/�� �9׸�!by�f&����Bn��t~�m��~m����M��2�.��\������R�|oY�:�M��{1�ޫ���;h�>��TP~���m�T�I�o�y=�1�OZ��~${��g�`�q�Empj�ѱ4��(}#���X�2�t3;aup�����-o��gT�$V����w���� ��v�B�l��|'�T���*Q8�4�e&�����!-U=���Y���m�C${��I�^��A������ykq�uL�֙���׽�s=|�>~Y�~ �jH&{�3	0�G��'Jϔ���y��~Ș��V�G�=����}�\�P[���ڌ��N��Ӛy0+��;V�t`�{XVf�t�9��:�9X�[`�,Y9�@�ؾ(�p�]%�u�W���~��3�dЛ�B�i^y�g����/�
X��Ebe�zzL�A ���r^�5s�F�S?T~��2�Lv�6��vE�.cvc��r�T�P��y�w2�6�A�G��$��z'@@o��6(�M��{+(
�'���ƯA��$�4Ҽ��}e�������Ѐ[�os�z�.ͷ����fX����L� �M5^]�!��I�g�k�{��ĂFI&`$����C��U}T*�,�Q����氱d�y�xh|yr�A�]_�Ə�;�*�k��S�j��yQm'�t��=����Ʒ����{��71 #���B2�����ܫ/�jΝ�����X͔���GO���yu�2��+\iQ����Z�!qZ�R�y������}�]�)�EQ������Y�4�k��#���s�GVT�v�];��uXlg��ln���
<���㭸��Z�{[�|�e���9~l�c����{vS�נ8��n-p<uA��7[�T/U�%�2ue�^�Ŧq.��Kb���<b^g ������L�pmɪuy�uڽ6��x��T�z���;�gu��a1g\v6�F�Q��U�<�wuϛ�Wg���A�*!hժ����7\G�N�'���	�^�5�_�>�=��-	�v����� n�ݑ�*�.�ӗ)����ӀD����oo��ٷݽ��y�$�'��[IM��A"���
�%9�]V#k{dv�x��Y�[��i����h�9���C�i�3JMJ�i�	{�%fc��l?z��� !<֚��s1�g��ܚܼ�~�4</ʨq-P�t�LI�t���A^V����.� ���~�����=�S��^l��%UE_�Ҥ(Q�m�����q�8.�1�خ����iI,�{�����_�'���f6�ݤ�{��f��o|��/g�۶�!��0���5U#)L:�����,D���qԳ�wFWi��-��-�;j�o�wx��ӷ�>�{.�)yJL�+S7\�X��}���鍊x����<������|ߢ�!�Z`	n��f�9O��;W{~�9%`u����Ԉ�-w{�c>$��{Z�C�l�}�0@�﷘�&����e�.�27������Qv�0A'�o�s	 �{�{�&��f�j붘%�^O(�q4�F���$��b���)����
�{�� nw�%��uy�m�s�/f5��۴u���\��!ٜ/rKѓO
��0�O��׈-P�t��ɧ���0�_��9��'7�8 �sy��=G��Rc7�ϱ�pP�r�fw��]�7#�X>��u���Y�_��U(��n�G�N��7���==E���nk�שaD%�g���|��敝]�\��t�5|��{�ȹw%K��/[S<} 7�/=�õ;�|�T�E}
!B'��	o{�3 ���du0!)4K-�6O(;�n.S�!��^@ @���`^m,/�]�lC9�ԛ^�;�i6g�1Ö�)5^����=�	{_nBn���h�%���ݸ���fn�2�7��Fl��y�B�@�n8uJLk�΂��֮��VcOOTe�~���>RԶ)�N���^�8��
���g���3����d�wوD�n��죵hS.j��:`*�9<���-����qc�z*�w�m��k���4�\��jF�Ni���i�/����~}��N���@��Z /5Ü�:͛'��.���R.��s� >^T��i0��3ћ|s��wx��Y����:5����䠣jAo*]m��]���jl�"9�h�iZ5Pfi4�k�)��Vu�n��ήq4�?� }��t�v.�Jq4��-���B>�7���jN\�ƺvt���޾݄^��	n��1�m�����<��Y��6�^ޏB�W�ݣ������oYN�\�X��*�__�o;��D����rŒA���A �{�x\&�5��=�{3��U6�a�q�Z+�[U���^S�.��_��� E�p�{ۙ����VV{ڗ,iֶ���ѵcjЦ\�.MW G7���t���'��ͿX�|֘#�����F/T��CM+5������NA���&��I�痢�$��ݶ�Y1���A�c���G��]�����m��F�B�;��jR�����.�?_�N��?Gޱk;����-{6RjӆPx�27�<N�z��`��^�~ݥ��<���Rۓ''���G��_Ea�廐��""!�����q!�ώ�m�utͽkiD�x`}� nv�_�炍u��\�H�;�ܽ�:D�=G�e�5��8�����^�ָ�LӇ˞���9��l���ݗmT�+ۤ5T-h)�f����7����x8�=�8�On'5,k;Z�Z��ί��!���7�]��'p���Í�Cs�����ػ;��OnK��HVQJ�������/y>��rn��^� ��ݵ�#�v�s{�5���M�3"�A�K�i�̃���/n��#H��b!oy�̄P;�P�zq�٫U\]Ԩ�v}}W�6�Si���fA[��.u������L	o����X��A�J�ƔP��|�fc��ݞ�=�%�$��޻$ Y�������bűtb�IM�6�_�W]�,g�2��	�a�:��=���	+Ӯ�$g��n,���eVT؈@m�b�,���ٷOl�b�΢k����u���i!`�j�א�R�u\�=�fd+}��n0φsPj�_���$�Ry�h	�V�v���=eM���&������3����.h��y:X�j�dy�m�Z�Xg9듺�u��{j�b_n�Է���ު�}�S�7��$O���U|1������}�+o�.Urw;���S|E�W�D���|���w)�@K��i�'.Un�x�]�ݠ3q��S��ݶȋe�=}�*���lm��,hB]�i�ۻ��^�8�����۲�]�|�}T�fJ �$���Q�떶V�.�0����{�����A��s�^���#
��Kk���qvc�6�ۇ[�bvZ��Gde^\}8�-�[d]5o���Ӄ�G�w��^��b�'�ww���HX7���L�_4�=繘O���Wdﵾ����Y͜{w{y ^�����w�Vj�E�>`P�Jѻ,i�n��H�^���N�ųc$Y�/J�;��M������n��ުSXT��S���Ƶ����fz�l�*�7��v�ݿ(������:�E'�| �����wՃ~�{��_B�UMl���@�?���:�`�}�&����W�S��O|�\_ď%^K�U6R-��%��Y �����>������4}��,'ⷽYt�f���������d�	1��CC�਎^�V��6TH�\(�y{Ӫߋ�W6	���n���\������\�gVv�1����s/+
Β�n����,��1��|4q�.��?g�L�I+{�,m�u#�vW��F.���S�1)��f �m�`!�����W�9b�9��dEs�qb�J���$l���z��z﫞�7m� ��$��>�����g���;���-P��b�v=҄�,o�M���zϷ�n��d����B©s6���2�
�Tf��}߾���ߦz�X%�BK���Y���?�U��y���ޚ�Kݓ>�T���������E�Rg.���F�&�;�<���Tq�,��%�Nn��+�rI�e�����%zu�d ����}�U���KJst(U����_��L��iTtL���v���ޟn^�E{�w �6�b�J�]z���Z�'إ�	�uԎz��;�mH�v�.��!L�չ?W��/�3��k��[m*+�e{ۙB27H�M��� v�h���uso��2ie�U�M��X��T��	)Y���o{����wu>��� O����OEe�}��xg˧�n�gOh�!�]���dL��
�K�x�w5��7�oM�ܴK@�msmV�Yb�FR���S�9X�:/��q�����9)��5�+�1�^�W)��b�y���*����ِ����b7��d�!*����:��:]�����5������`�nv@J�����r5������}nN}��t^͙Xgm7M�!'�}��ыHl�i���WB�,���]َ�ĭ,|�'�T�|6n�w��n�.�٩u:�x��O��蒋�w�=O�f�;��݈��s�;3��n�U������V-+D3`�ӹf�i}�F�Y��i���k�S{�Vb�8&�+�V)S��$,��8"C˹�Uf� �J���ɴ/����T@��rpsn���������rݔf�B�O��{,Suۂ�V�Uϳ�䚋8)���Dt�#R]�gN`@�+��k-u��BԮa�O��ľᥲ�(�Y����w�o^��֯�m��w(�"��Վr���1��B��̚E�������~��`	�sE-�E���e������f*��s=ܶ��E���*T�om<�3�k��k���D�9+��Dw#�|W^QOd�KYh��ӝ�c*	\[�����ޅ1�L��$�����Mǎ�*C�a4�uU��Q�T30V7y���׵�Y׳> ��|&�JA��"`V��iR����K`��qj��-c�bEE�`Z�Sڥ�ҵ�����[[jQ-�`�,��j�h��1K"Ņ�0b���-�E�ը�Em�����,����U<q��yOc�F<�<�.	YlV�KS��8eDh�����l�8���81F�ѥ�kB�R�U�.�UEVb���TR��Z��LR��a���ZQLb�b"�����ҋT�[b[U���+L\3�ڭ�Z"-m�"Q��F�F�J�qb֫mTKX����E+hҰ�0am��,RҶ�b5�Zm���7Z�4��JQqp���ҭLYQŬ(��X��j�jPVb�cT(�����n�����4�[q3p!v�P�뭬s���m<(e��Q/3��.�7	c�+�K?��k?�GOzҷB�����w��Dݫq���]g<n./���N5�f��yf5��b��w7gr�^���&S������=7Pm�m�{;�����D�����"�]aU�Dt,9�g��t����wP#������,+s��qF���>9�֭��Ot��D\�ݲ��v�u�G>r73� �[�Tv\v�;=N�s�"ES4�n��:���$��أtr�keym��-��x7cs�[r��m��'yøN�xQz_Z0m���������؞��p
i�uۥn���
�{p��۴t�M�ۧz,Y筲Y�k�:ݫ<󰣞�;��tm�=�TL��o�"����m�V�?v��v�����;9\Eڠ�ճ��ǭ��s3�8.Ϭ��keݻ7a�h�W7ORX0x`�]�m����xx�¹ĬNst��-��n��=r����m�M�:��b�0�90����pF��ᛰs��vvx�k�/���/�Gn3<���e��<�,��G]���Ak,�{9�69[�n'8��C"뫲�n�h��)������^,8���X�#ԯ����۞���|��s��mP��?�8G�0��rO��i��m���l巀���s�,n6r�l��5��;i1�a��Hn����	r�/c;�0mu4��ˎ�÷���x�-�Oga�1��͌�Q�v���f�h�;R����c����vl�w3�ك�������������}��ұUS��_]��f	�Wъ ۵g��%��\8q�K�]lr]P�7[=�o>�6���q�w��瓚��oOc����<8�H/Z�7d��g���$���}��>\.;\r:�'lp��s6�y�%lQ�x-���6P�v���M���`cqŨޝֶmyL�
F���\9^-���m���mf�PF���H_�<KX�%���z��lŢ$���>`�ݖ�7p�|O9�պ���N��p�؛��Y���5TW��uU��� �G\<��`�79	��Ut6�m�d�m���\�n7-��v��Շ�P���M~dR����"�u�ٶ� �ﻙ��^	��ߎ����VX$rU�KRli�ӫ����ݕ�f��;�w�c$���c�r�١�k�Y�Yc�z2�&
i��Mv� 9���G�̲v��}��=6�=փ���#��J�%�c��{w����aWt��e4 9��s  ��^̗�7ӑ��9nO�p([E�K���|c�]���D���E,����u@Cܼ�i塟q�Ep�Z��`���*���&�c��r�L���54�{��N�-���L#����@Aݽw_M2�<쾒R��37ۘO؋��B	%�y�;;dT+�{�0<Ux *���{j�"������U�ލC�-g�Z����I�
���٪��m �9�����>�;/�>��z'A��|���~O���n��Sp'�*��S^O�0� ﯮ� ����ׂIu!	g;�fݽ�R�[�QLB�ef#��_��;X�/��Z�H�ߝ�A��^wo����S��a#��A6�[�
�v,ny3��u���Ő#�f!�ߚ��֜˕��h�ө��u��у���%#�	oW(t���TCI�Ro��{jv[T誇U�w��!��� ��_��+R{PL罾\ y{����
M�,�L�{���{7K�w��	��݂y�
���>�^����15UU��on�^v� G�9����	���wC\�z\�����]��u:㡴$����c�p�O��衭앜�+�b�W�\����Z�3��(䒸L��<	�}w��d��}J�Ӧ��שw_Uʿ%;�@9��I�'ee���F�xRoǮD)�����"�+���~#}鷟��@y�ڸY�7wܼG�Q]�ξg�/�/�k��r�:q�A�׺cf������cۂ�kY������-�2���ݥbV�4�#}��^��N��O{�}��j9n�.�F$R��P�S���<�]���A�u~�U�˰��V@�kM �n�5����g-�\�"芯2Se5�A��y���@�^���ro/��Vm&����(sͩL�ƝUf^�s"��du�@_}M+��3"��^O����ݤ�&-��{�u�(f�R�-����7Y[(]5����j���<������I}�wy��HW��nVP�e%�&�����0����ه���0I=�ۃ ����57%O���/7P�-L%���iϨ9V:�Ħ�v^ǃN�'[�=Qh�I�=�Po�)2�u%�~$�{��	��v�+px�7�4#���1����%�*)�ۻ���5�S�Z���t��s�S��ύ��$�<�X�K�R�E��)�S��	gz��H&�wޮ��0�vOf` ��ޱf�M��@Z��x�f�w׾��Oyw�I">��J����JVg~ݓ3	K(}��1�4�0���XWg��_0�@�o{��n��s�X%yi+��d�����_>���F������%��c���oP���½�{�7�l	,~��׃�w�*�]�^��8���A��
���bwe�Zޤ�Deœy�*%e8m�n܀6x���m�r�ayɻp�N��h���b���X5�۝gɻb����^s�kqx�tGnc���0���í� 7�v7sԛ�Z�!bמ͹��}r�60��u<uM���y�˺�ܻ�B�zl�
L�k�nk���&]kf#q�l���a�B�s�vl�q���M�@��Xd����a�Cza�Yw������re?�M{�� �9���J�����v�e-(=ٙ��=Yc<7� �$�e`�����86?_��	#�s���M��֫s�����θ�6E1ѽ�R��Om���n�$���Ղ��S\�k�b��S)�N�f5M%'��:�����X��$�W �����:���Vw���`Y �&��N`���� n�L6dն�����	U���w}���\�67���s��� �>c�K��su�?�׏�_��$����c�Xt�uw}>U�8���qL��+B1�Z�ww��=M����sn|���+�y֍�-kD�M�Zj��}�0�~Ş=�)W�{u=������?��(�Ȇ�7à�
;):���҉l�_83FMw'n��8��KӁE�������!T '���3���V�K�y�ϭ��c��L�R�$������A�F-�C���h��������)�i�X�Cړ����������(}�{[>�ԟzx-�[A'yq`�{�V��lԦS̉��dd~۱n�S<������d�ޘ0�ް.[����Ψ���A
�jv���ױ>=v۞�z툝���bp�����%\\[���(�Se*�Q��I����y�*mA��9��%���L�N/U�>N�L:�l]�� �X��_�׍]p��N�@~۴��{:�t'�q�	R��\k{��k��60��V<�����zK�"�=jV�c٢��݇��5��C�Yέk�1_M��r��v��5*��>ʺ�g��������&NJ��f�����jƳxk��J&�x*��vr�\�Oǽ��`$>�E^�+���*)�kG�|�S��;.Q�")q>�2�k�ȃ���kj���<�vo��W���DD�?V�̋�X;ߧL,��s���\=��N��7W���׮�!���놪�Кt&S��30 �ݻ����H��v�/6�>���r�:��>ӎ����V����w��#o����r��  ���pK(;铏���^W�tO�5%4�ϵ�;n(c���{���� F���Ёd��:o&���	�[j���{��g��$7���I�L������$��,�[R��GJ��3v>C3��T�]����fG�݊�m!�����Q:i��܁�VE�bFY��Ù4s�33�}��]�Xs�Qi�(�c��*���ӻ�i"��o��\|�`�v���9~�{-�T
�@��my�tT��z�č�n�k�z�I�6%3Z�w�ɂiK�%��=�^=�P�#�+�[[xϻ-�<}��O��?�uc�~�6دJ1eV.�>�(
��2A#��3>$�\�:��d�
���tU4�>>mwӥ�$W��}u;}}�� G/����x����S�����s�ˎ>��wG�V����3!���3�g���|o����e�9{�a��kNq�T_��({�d���t���u��^��L�R�7���h��]�D��Յ'��\eQ�֟v�ׇ�8�%��Z���_x��3�������:�=}FH��P���ൊݻ;y�^(ۭps�Ͳj����1m��y��.&�^۲�X�m��]�;v�z�Ϡ�B���.c�,cb����C�ul���a2#:���ܛn@�=�9.�S��Y�U���
�I���F���ޮ�]�݆ە#c��jn�6r�LaF{)���m3��/�I-�@�f���3͞` y���n��yzl+��Yt��{��i��Re��W�#��[ P�^H]9��w�9N��	�v���;y�DR2�~�˟&{�?U������7��@���G{]�]�+�JԾ\j\4��������^�VA ��'�}�62�a$�L�I=�����!qZ�4���?X��)u6�j>N� ��
/ru�g<w۷��@�}{�[tk(qN�R� ן�Y$7Y*�P��z�׷o��J7��hH2of)g�7��"��J��<h�����z��s֎�O)��U@rYeU�R��_w|�� Cb:Ս����Z� 2oe���Ž�7ݘI'e��Ki�F�2��&��n�+
��^"t��Y���uWKս@��p�h�S5u�ȕm�3�ɔ
����^�xc\4�{=l�aЕN�h�#�p(n�HPex�^�#�C=z�{+T�˸xw֦�D�A:F����ߚ$�$��c�j�wă=~�h�7��^�]j\4���������T�~}�h)���B �ݮ�����H7��������_$��4�>+�D���//3k���B�뿉�}L��)�*ח	��D0N ��&�F��R)��Z��Z&�c�P#\��YC�t:��'^ڰ����w�[����_���%B����@q��M@�Ai�ϻ>~[���-����z�P�5�W{ݭ�7��̔Ӥ-�tɒ�� ��Z�{���%�?k+�|n_��ܼ��w5�AE���u ͞��op���E���85��LM<̽���5b<�u�z<6����*s�囸������v=�����/R�6�1L|���Ѹ�a[anp��6ᬵ��.���UՋ�����u?݋v��S�<䲉6k�������+" gĥ'���B�r�t����Wn��
���A�m7�(�"�[H���� �u��7]�F��+�5�����h<���,��	�W��1���q]�h��U3ϺY����yw���v엎���Lr���ᮈ�n��@�e�$g<7o��n��6X�����ص�ӎ�겲]���8�X�O]d��r^Wt�y��/��WJ�c:*�]�'t}�^ȹ2wu�(m�ܳ��{����ҙs���MTe�|�M3���n��P"��EX����X$���*Ex�v�n�̼l�p�`���ce��z=��ٚ���fr�t4+
ƂtEo:]]b�j�w���%��W7r_q��tjZ�x��|�7�;Yk��)gG���
�#x�:�Pt��*��ũ�=�Z��次�y�	\�k*�eNЏd�q��^�;�f���he�H�s�����7w�2�lr�gz�|�[=Vs��B���\�+sE�;����q��G[��v�Cڥ��mJU[0�0�UF2������J�n���.1�V"%��
�0#�Q1-qq���LL	YL�.a���-
�KF�H��
*TT0�p�Z,�,��F�
�(����EiB�X�ҪR�V5mm�A��1��[m�mib�D�����
V��F��0mZ��Bڸ�QUڴh��Q���4�%h����-�)[c���g�B��Ŷ��&mAV8R�+����ʰ�\Z�lj�Z"��kF�j6�kmkj��" �.-��0�8/.���\888�Qd�-D�m�1-��ŉVʕ���U���J�1E�jJ�&��ek�cJ�2���@�ʠ�k"0pY�T��Qp�(�S1J��P1�.1�2��j
�X�iY(�Ä&*ґeQEBڥH����)�׷"ŝ��;������J@�����&wH�j�����0 ����o���Nܸ����2�gkٙ������Ƹ��,�,�\��h!��s  �^ڼ��-���U�U�2'e�>n�\!��:]����\i�jt�VJIo�w��V����=�⦷'��$H�_��6�����t��d�=��0^����j��������g'M&qQ�Ϻ'�����B��:����ڛ�[���@��y{�O���_�X��j����.�=�����mX���e�%�%Sd�yՎ�iVV	�}����߮�$�墓C�z������ҡ$�ju����Rd�:��xd�n�\��W�G��d��s�K]覫%��І6��Xp?�wY��\X��X6E)��ә�i�ι�u���2�Bsw׈A�^ڴ yZ�P�����M�Ӳ�G��Q-�l�z�P�-�����F��96�"�����~}�>�����=��;��V�V�w�9}3�6��#_>���`�L����LJ�����4�Q��z�~�?94�@|ö�������gf������T߮N��9)��D��Š|�����-�ۺ|����@�V���$�3Cu*]:�Z��v�e���%Y�˵b@�2�v�{8_����$r�ckj[rJ�<�;R�I ow��8n.�|䷛Ʃm��hW%��s2	Շ�L�܎j~�0�5�JT����?�2��ܺ]��k�����YwZ��}�ʖ��Ƴ��'����&ͮ�uf�U��h]��-�')�%����1\yt�f�.��䣴e]�bS#���Y�kۅέ����S����nn;���N��_��J|�Uɖ�nvT�����v۶RKq�0m�Z5�͘�4�1^��a�,՗�3��u�;^��S�ً/n�m��<i��v�-�ٺZy�uX�g�c##�l�y[I���tv�5n`�ĺ�.z���Y�[�tN*��;%�[}����RM�~�(����C��G�z��#�OpX&�x�HH#	�*�n�{י�D\ޜ���^Mn��@
��4 �����٠�&x�O[�dx.Ԩ]٧N��Wh�A��m�$����.��>$�+F����	{ru:rP�/0�=��R��3FM�9�'��읷��A�~�9^냇S��`���)5H��SM_�N�ρ���g��hԭ�?ll���>�}�:��������4�d[j����ݨC���8�w�h���q��gWR��vuWeJ��Bxm����y����*�.Q�s���A����j�wЬDR�.&oً��έ{Ϲ~�Cx�y�d6�j2��co\Z�]��.����g�����m�������������9P4���� M��H1��,U�ϥwaSK �Hv��TEK̍��b�<����X��N���ww��:�_��*�)�r�A=��s�o��� Ewy��o�� n�2��	oǮ�J,�d��s4����L)˼+^ڋ O��5]Sf���g����H+g��!��`��{R�e�)��� �1���g�6븮X�����.�Ηz�&�SFzw
mSDSMys�~[� �C�����7r��>}�3 �V���i8���PL��6(�q��f<g��� s�v���A��{�~�X��+�Rǹ�ş^�m'�~~/;xeૄ��u�ׂ������8�n�|ݙ�z937I}�6zM>c=(/N�Nـ�ڞz�V[�h���%k�ҫ]�x�z�C���!�cD��*�n�y�3=®u��L�۲C��?O{ۜn)ݝ�,���?z�����:C�T\"}:89���_3����7�܀�n-��h{ۼ�b��{iI�����f�n�g[GT��7��n>M�;=!�^�aҭ{����8��Ǌ{\��'�$ ��{s],-B�;�˿�奒e�j�E��U^�\!뼴���u�Hqid{���CW�t�s�]Se���l�@P��buB��8�mΐ,
�MK��K�������o*f�QNje�������̙�[�mH
��^���[�FTV�r�w���Y��P��t�r��V����W�\�=��-���H�O,���+�l��}��B���ƴv�MMx3�B�aR��:�3!W���q�h�X#��7����=�X����'��q��]��� \Bn6GF.݋���sREc)d�IV-{�A�5S����� ��ܼ@���v�s�mw�F�NƬ�A#{�s	�R�ꁆ�A������=xe�v隙]D {��� ;�`�qr��w+T�x��W:�S�������� �I[�do����K>�x�:{o	$��]��Fy�T�T/0�M�(b��}Rȃ(���&����@c�FK���PIP��j�CgEb���q�{3�^��[�'�c���y�fnd ��\\<�Ӳ}~�g��:t�w5��6g:;J�}+���Y�M=��{+׊�:��	��r�R�Z�ٷI�ŸҺ��K �]��%ϷV�@�.�|\�5�۷NЧ7m���ӄ���:2s�ڮ���۷]u�{%��v��;n۳�^|���q�k=�dJk���;fG�v���=���� sn�=���l������u ��m����7QP��eӆj
ù6�v���oi��8�K�
��
�"�{e�=�Mn�W[>Uݧ�ƹ,h�]n.��H �U6��s���]REX���돿��+��7�\w���mŢ�h��>��w�pI}޻#���h�K��W�Q ���G;x:��^A}޻����8'y������y�y�^����M�y��{p��r�@���-_w��3��M���V=a�_)���(��V����hm��EҠ���X�A�\X$���^p���{v��$���3��M�H�w�Ԧ���/�]-M'�.�H�����������d�Gl�]��űv�s��&&H�e����H��
B�&�U����X�-���yq���h���xj�&��׷��P�9v,	�	�k��K)�K����*Psy�(�-?xU�5�H�u<��j��o#����):ׁQH�{O�-;֫bԃ���l0��+�W�+q�ֆ�,b� �$��w�g�N+}ؽ��o>ཁ).������O��swݸ�Yu��L�۷��h���{��]���n)60c���[��d��V"����ژ	�����N���M�=98�+r���6���_)���tV��$�'L�~s޿�k��C.��x���/pٳv�u��۱+*�q6���Y�[i�+](�����MT����� �oo '�m�+�h���V,��P���4
gM5vh�qu�:�YC{ue��OOt� ���B$Z�����졧��:T¥�ޯm�b�E{�iZ���l[�$�d^\���% ����aӰ�d��x�X����Ì-�*��-^�(��jՎ� ��3 �T���#�����,�D5�]=�{�Nǭ: 
��|�ex�{M�$��Y�EP�3�e�Ek��Nz�6�6�=�5pׯ3'�(��(����%��x�fis���d�z��%���t�Wl����<y1��xS��������Z�������f���o��2{�BI$��TH/e�%ǝ��s�:k�����/��`oKj�:���3cRXI>�#ʹl�M�~���g$���}D�z����i�}	�qN�(�d��_,�F6|��x��e]��b�Ow��{z�ص��b,�s��+p�ۚG���q�s^����{�� ��p�������ݾp�S=Wb!F�b@�(/7���+���Uk�\s�g�]���Rn;}s"���x�S��c_>�:I�N~7g��&ST�<��{��؃�ﻭ�9�D���p�p 4d�߉$��w��������s�^N0����!4�y�e�I[���cZ+�V�K%N�P*�7�]��+]us��qI�n/�����t��y��I5=�;e��V�L�L_N�_��ŗU�_{Z}@��}��a��cg����Q&�'}�t��=锖]^��{��'pp|�0�O
F]�uU�WOwf���Z�����{9ρ��{& �G���>���߯�h�̻��'N!�ԗ�gSYP7�r����w����z�pž�Cb���Dؠ���Z	�����yzI! �8{��2^Vx�H6�?a�+N��IP�I9��EWޝޯ.K:��lĪr'6�WT��fݖ	��^Z�2�P��)�iG<gb�i{��^w h\h'�=ZM�B�hI
U��L��K���yG�d��X�%�󴙦ퟁ������wr	���|7�Z6u��!�Z�\�4!!�|m����_/���s:^wry�Dܓ^��"���zĉV��ao����h��oS+�<����N0�庻&�Y��ڠy�$aJ�T�n�:��sJ�5�S~�)�8�]4����AQ_R����4B^Y�s6�M�o_�Ԑ�Y�3�w���H4,y�0�۪hX�8t3ϛ��tٻ�3wV�r�0>�Ґ���5��3��:�������[��A�s�5��5�A�;��6�9�[��e����ғ�d\Ĝ���6E�[�iP�k��&�gNfZ���y�u)bt'*w7�}x��	4�Ԩ�	������m���	��ا��;M�v`���QT�ުk�Ü���{�_Ha���&�\����z��)�d�Q��t_w6HvZwٍ�h�g��T�ѕ��{8ΕZ3
A�Gi��2��!9V�'���x����J�u�����W�ut��bB[��׽�kv�;ēJ���}I�ws\ur_#�]ǰ�36�5e�@��&t|�0G���V�E�5�u���]�������S�1���'Uf̾l2�B��(�p� �,Qp�.0\Y���2�,�,EF��+��iR�p��+*a&-�,Y��J�d��Q���T�qT�ZQJ�\%`(�C
2����Z�ŀ���
��D[r�U�P��V%�*�`��U�#-������2\P��X��QX�*2�E"���X��-P�����Ŋa!Ra��1i"��(%���Ab�\5�[j)��*��Qb���n�H��*���p"
�mEL�j
EX�X�L8K�	h6���j�,�Ķ���"01j� 4��P�K\Y��*�j���1IRE�)dQL6
J�EPŰ������
Db�h�Y.E0�*�aR���ZE���ߞ�xpb�5f�&��z8�>���'���z4�lƇv����Vy�n�Y�<MR����x��vt;	��J��nA^������q�YCQ�����������:)j<���N���s�jU6��mۣ�=e����[e��v�.�m����̓���2E��6u�n�Wv�m=[�<�#��Ogk�x��j�@6��5q�"��� ��u����B@�a�n���lh���9��k�4�X&�v���ޜ�Nb��:�i�;&���I�qں�M]���hԏ2�G5-q�ܞ] lc�<��2��q����:����f�#�1��>�m�M���[�#���u�zܧ��/7n,v�E���.f7P����N0�6çi�Y��n<%���=!�x'��ۛ �4�G�m ++h� ���!�n��㴼7�5m�#��Y��WHm��m��;�m<�( ���ڗ�{O�#q��4��y�nx���t�����i�[t!�z���/ou��j���s��Y8���^���=�.�	�u&�N.#ͬ=��:������o�V�S�2��SO'n ��N����^���p3���]��7����9��v��nvq�<s`���v���|v��[�uӹ�u�2���� ��.oF1���V�\�;Z�%�n�]�l�0�שx�2�e�<�z�x��ue�sm����0��u�b��ڢ����pkPZ��^�2�;���5[�S(h��X�=�+ͣ������c!5�]H�]:�N�Z۵q�nb��6��}��%ׁ��v�%\��j�}q�n	�u;nz��*��U3Nn�y0p�۲Çr�좴zۗu�&��v��Ԝ���v�ǆ�����*�����sr�NM��\�),�=#�s<���lu�q�Dv��n��y8���}���X�c:��/^N<sͮ�7tۭT���8�����kn�r����NM�%�nN�J��y�/*��p�f��a�8�Rln���F�x��OIl]f�n�UݹGG��z�نx}�qx�puͦf5���Avm�ۍ�W7RS��;c�?Cu�*�A1V�]F��k�P���.�cfG�N�ã�m+mVU����߽�<2�R�����f* �}�o� }y|��7ubs�[ҧ�� �����
\�E>��]Z�N�g� �+_��=�2����O��wH�Fm�`
�n�mE]>t�w�_|I��\�_�ߋ.��������� ;T2k�>$�#���!��Gr��X]��yT�P��WH��=����N�u���@�RO� BO�x$I$�>�˯?Wn�=:Hk�V�}��s.ᙤ�� q�v>w�Y';�󘀚��J$�H�|0TK�h���4������݈nH�'S��\q�T�`�'Mv�qn��gq!v��N��Ym���Mx�[|r^f{�M�~_�X~�TJp �����{�`J$y_�:|�	9WXr�6tg��I�x�5:�L�|�N9\)Ma�t�R��9j���恺����~�$�,���4fE��c6���&d1��n��B�G/^ ��X��U��[Յ�����ޟ��Z�W
�n�޼THkń�H�E������LX1 ���o'}g��w�ˬg3��j�br��'��$�7���@4�j�_h���<#X6GQ&����[�O*������dm�{��[�<�q�>�m���zO�?Qk� �?w[E|I$�G���*k��+�\;U�z\�n�":A�k\ڳa���y�vJ�n �8���j?7ƺ�� �esX�ݲ� ��Q��Ow{���s�9rJ��6�iI;��IĻ�D��CC��w33���ol��*������Ma�|�=�������9���s7w=;����o��8�˱!�+H�H��͉�&��"�׵��q��f"WCCq��0�4����}�`�wPY�m���4�l����+ۖ��͉�S�����3�j��N��Z�A��O�?f�AQ$���s�	��u��+G���hͦ����A[�D�I~�s`BI+}h�nX��tI��3/b�쒡����=�kO����O��h:$�1�D�=�{��A@ ��bXk����s}�|\���IYs��tt:�yY��z��I���+,���ͯ>�uT�PR���?fe�A�s�����a]�J�����<�X �v����ڿSE
m2��<�z*���f��Xf�th�������4J�Z�A's�6,��~�9}TH��D��C(X����zI%Bh�D��X� .�v/m��'�IS��l`7���8�t��R+,�0�g{7�����8�A�{\�� ،��`%��;���G� +!6�ǬAd�J:�p���Q�!��;�]yھ�u�]�N��I�舅��٘)�ow�r��������;	��i���
�MI}���~$�J���_v�n"y�}�<�gI)]R�i�8v��6���Tc6̧Es��Zީ6��s���~���/ŗ�ȗ������<�r�Ğ����O,�ݙr�a��zF ��L�ٵ�T"�J�]#���J��k��n�7|��&�4I+���$�y�Y�m߼a�K�.�{���{�ݴ=�sJ�-���|�����O`� ��y��{������Ń]��� �;�R�@�Ye��{33����WO�yBI>���~$�}�$�E{��,��G��8��ԯ>�֛�J��=?e��|	+{��Be9�{����WzI�<�*$�g=L2OĒ���>��̩Ǩ5sb�W�۳|��*��=�v�8���Z���p\��m��U��2]�(í��j�V |�U��^��G:�kݭ��E���-	�wn��`W����[�$�zE]�\njn�v�=�Cu�{'��d,nm�	��
;�q����gm�b�����ә}�ü�[lf�9�#��2�a�=��U�f�2FZ�y"!�4*\Ӝ��!v;+��:��F�؈
آ1�竚5����_��U�㫈���A\ևx�����"8�(!�*�A�bN���=!�#gie���_|~�S-�?|w�����sH g��>%��o��|q��x*&zZ���3�٧�>�]���6_��WD�����}�o���b4I�OӞ�I��r|rp��߼^�,�ش�x�RDG(ǎ���6H���r� ���[�'�H{�$�q���3��w��{��S�B+,��4��g����w��p��ۚ@  ����� :sǳ=����%�oo���5[Hhcvwי��H=�V�����67@ϗ�&j���ű�s�a����5w��Ob��'}����s�n���2s�ӱ����l�ۛMg7~�Ͽ�Θ�Z�>��  3��u��Nx�������Htsݏ�ɀJ��a*y�B>��[���y�gnyy_�յ���"V��KC��t����m[�f����I�$��-�����~t�}��h������B���� ����[@�g<f	6kK�c�5��;�,���Z���������$�8w� �yP�9�_��D�#�﻽������X��x:���`ǌ�+�����ӱt�M��� Me�Q'���/��s�o/�%�o�F����J�m�]�2�Ь���눌��(�w�=�	?NS�BI&�^��A$������3O3��s˱F]U�S�rvm�bj�:�����n�[1݃�t$U�~���qn�]r�x߳{ޞ�7O{>� �2%���+	X��{� 9}�s7��e0�i�s>��Y�P���W�נ��]��	�I&���/�4I{쌰>��|�^����y�Ɋ���ڂ��H!� �7������Os%�l3�<�l�E�ț6=�.�o:�&\ں#ė��u�O�5{)��A�v,����v�/�a��GP�Ϯ�䏻b�� *��D ^�#,���FX���������F�y�l ��@{�#,�I<��+�����{�e9���|B)�����i(  ��s��V'�@��d�����=�d�M}۞�Oӯ�mD߻�tO��%�tv��h��+��a�˭�)iM�����w�����+��@��. ���i( ��}��|^�id� v�f@*�nFY&�g��W�g(`�y���rHCZ7�C<��u�pH5�]�����n��UI�X7<���=�����MUV�,�<�k�ZzA�ﻭ������4wdKȒ�<c��Q ۑ�I�J3��w��
b�t��[P[�wݴ���nk��7� >	�N�|����Ί�����7i���c/���:�;�*ruqw���g��T7���_^hx�NZ:w)�W!)���+�:�c�]�&�F��m�|*��s(�o�ZM?�oS}�n�UF�^ �Ѣ�w,��n6]Q$�����X��,;��qv|�Sp�!�6��kc\�҉&�,���>��J�N;S��z�^�I )#+��%��H=��u��9�M���w�{�����?.�F%x�Qu4i�e��=wn�U1�Ok�s��/� :$ž� �I�V��"m�h����\*��tP�i0Ye7y��r1>$�z�h��
璾q鄀Q��{����s�0>�Y�vYj��d���n���c�j���l'���I%wZ���NZ��H�G�}鿶]���ڂ������ o��N���u7V�zID�M}�"	%�2���S�}���cbn�gE 2N����d�P�X�y�b��|��!r���&�oޒ�f�/�|m�Қk��N�ꖡ�!����6�MKw?��qS���Q8�Wm�5�����'[��8�p�G/�={szz-\sOmn80q��$XƋ�^x��ϱ���vY�w�-�5ۃp<v�:���5���4�Y��<�Ad�ҸN�����ʗ3���`��l���z�ĺ�N825��].ug�>��y�34%�UYŵ���֞��D6灲)�R8�T�K��Um������<k�\��-�=���H�w� ������mm�~i�`BIW���D�ſ^HH)#+��'rwZ��~~�ֳzg=�zy� �~�S�de�h��aR��=k��mWj�kɣH6�/,���H=q�D�[=��F�s�Qo;ً���F��״.�%N��btw�ɰ�-B�!ٸ��^U��I=�dd ]��ȼ�2=�`�I$�KH'q��ܢ��dz}�����9�w[U�aǟ�q'�jZD�'��" ���I
���pO?M�ﰑDX`��{�
�n����񤄻-k2��N�*�h�����1ϤNE��;���Ē^���I]ړ�j��<���D��H�N���{Q��C,���iw����(�^�\:����*Yt�Y�K���Ҷ�����[}�x�M��t���h9P_gYG�x�aj~�:��oN�g��b��w�� y��O��~0�y�p�m�W�a�mI]�g��r��w���� �ͽ�����{��&��눿� s�s��T<���m&]�'�1t�^��Լ��g���`|�A��yw+׹_,|H�v�F� ����ieN���=ݹ$&� .����V 6��5�I$����0 7���=��-X�A-}�3�m���ª�cGK�a.�~	���c�J�a����QJ�={��ֵ� >g��ml ���=������єI�M^�+{��v(Z=i|wؕ��h�9c=��5���z�Y$��yo�� ���Ńo��K�}�r�f��J��X��Ǒ-��0L��\;����.Ӝ����������Iͺ�\�u��]�H�) �)�B���5ZJtٮ[0�����8���wV̚]��hf��%Е{�Bf@�S���{��em�vK��;nT���Q�X�u���Z�"nr��/����(�n�]Wv�6�����&�-�w���a#r��WD�����d7��\�!v��dn|۽�}�]�G= 0�X\EQݻ�<VV`�,�K�p���jPoe,��ƶњb�3��%�J];7�{{~��pQ��(\5+GJ��XCs��+X��B��d�mm��{O���g��f1�:���{��7�
��HW`��mv*ŁE���*E���1����8�S�3\9u���=Ƶ���2X'�\5,�-&j�������t��b"�Ӗ%����%��Y]�%o���7�����!2�1��}�#��o`��-�o�k�f�I���U����x�b�tjuwMQ.���3h��ES��v
cx��j��G:L�`V�Z9Θ�u+2��p�NU�v�ʋ�5��XV$�18�b��V��\��f|K0�5m��	e�"�=���_�&�]ǲ���[���L��k�x�U�d��}�<+zf�t���<چئ�}T�l��'D�hw��G�+�1d��ups-i�َ�9��%;�Qz�f�Lib�V5z���V���3�ު��79�u�|v���y'-��W � ��X�"*��L&$�8B�6ũFa�Z�b�����őL$*��ecU�Y�T��Ab��DB��E@Um�"J��
�d�E�d�
HV#\8�-j�iJԮ�m%l`(
a*�R�n)UIm��
�Щ�E"��\S�Qegt��q
�U`�ͦS��F),X�B(,�Z�Er���0��m��Dv�)�����-dAE"��fPB*1j�b�TYX)�ŕ0$��R(�P1j�TFa�J̵FA,
���RE�S6��D���V�Rp�)mF+%b�AJ�h,
�Qcl��.⊲��+P�qB�I�j)m%T�E�`��d,J�*3,$��fɔ%E$�z�~�ym�޵�|뮫h�s�>�Ϸ�rAFH�VN��s����� ��׷�� H9阀@k���&/7����E���O���Wc2�4 �Ɉ 7�q;'��}$�c���$�D��H�S�de��!���koi�dO� �+h�l��J���Ͳ$j�.z��-,T��V�]o�~m����7��{��%yZ Oݑ�zMެ�K/E������0'�f��g]T��,�ZG=�m���~�xߔ��MQ$��|R$���tH̔��Cnv�BiVb�`���M�}Ħ6�ټ���V��/#�BB;��M=�F@t���"��������71�4gs�D�I쌺$W��;�'��W���b��t��T��G�q]�YD��˩�W�3���n�{���*��qMwB9����^R�}솥AB���YCG��f�fϹ�zB4H�Vz����%{{��ԓ	H�%d��攉 �{#:H�3��w��5��G�����jE�����#���7g��4�Сy����v��9�sY�߿ϭ�ꎢ+d���i[�{~��@@w�b9�eng������F�?o�Զ� ��~�Z�� ���ge\���V���"�$�<��$ �+�-\��IZ��t�EQe�i�=imY4I��}�s�@ ��un�Þ=s� ��]�� ��w����Vg\dQ�h�﻾�>͹w�׶��� o^�w��ٓ�9�K�׽|�f�����>����.�T۔6�䷻�!$���8r;�)`Y��2�$�{�$ U���'#�~�~��Y�3�d*�P�5�"|�O����W_.�z߳������r��1gr��ܷV���u\���4&�d24}L{�q�7�;�Ts�n��1��un�7/=V�A��i�bm�f{y�xC��{6�6�|x�v�b�����Źvu�p��=u/Y|+��ӻ[�z9KRs��s�� �ê����X�:�']SNK�&k9٤�{[�0����W=sz%82����Ֆ��.�����gPBrݘZu�LAv�А��%"%,I�u��(5Q��B��-��N�4H�_�=�Y �>{��T&�$�{�CS-M1}o�e����;�~^��4C�i2�4Ɏ�i������r{�٥�{�$$Enx*Dz[��9���"`��U�`�A7�Sۛ��MU_/b��Qۈ���IǸ�'�U���ilb��y�«�WH�U����|۔u[!h�Ko��*D�M/g� ��Guپ��u�`^�{	���dQ���h'g�����4����<�i&�G�%j�o�D�}���1z��Ϟ�|���c�f�j���7Q^��s�R܊ƟN-i�������e�3�_s'{�{`��� k��Ѥ
M�Ɂ�s{��h�WgH�P_�r�
HZj��;��=���������GG����w���nE���gA-'|�{:�R���;GJ�`�����	��E`�M�N�ؤ��Ytd��1Nb�К$��	Q }쌲I;y������oL�ڒr�0�L����Wu���M��_qU=�����ߒ��x�����]��>�Բ�$S1���J����_��h�9쌺$�J�{���h��1d�����Ú,*A������3�I����}esgG�^a3/F"I'���$�w��<��t癇��=j!y15l��h>���t�,^'�>x=���wf%�+Ge=����E"����銉$��ê$������|�s{�7�g0Ń ߧ���2���YlS3:7�ޓ�M�`���V�d�]�Ā]���4�9�wzo`���ޮI��P�9��-��� ����zgu���h�=��$�TNgqg�)}�^���~�m�7X��
Or�.��w>ζd�[�yW�:�o�{o;[�כ�1��^��7��'�]���Ϫ�!o{����t�`*����▿L���Vz���E�I��� �V�t�7�js��\�9g!�t�rk�
����ˡvj�:��>��'�Y�+Qu�t���۰���nZ���;�$ �K���'�>w:�����4_�:N��@�r�i6���:
K`�([d%Y��OB*�few�=7`D��s` %S��J������%i�}� =�s�����u`e��l���=�fc��􇎥�H�=��`|59�0`=vd�p��؉�oު�j�m��x�R���a$����I&���C�rgm���I��S�3�g%�$-5\�{��� A�{���  �;�3� �]����~�02WKX3ź��h�eߒ�dl�(�<sx���i�]tA����1�F�>�b녃�}���OOv��K��b��eE���o���|o�i�VWfC*�8V1k	?N~�O� �w�8 	��tNŇ$i��+n���"�Ðmh�u�q=��^1���[W�:��"n5���������R�x����l �5��0 {�2��c���x�R�h������T �~5�׋+Ǚ:E�	mZ|��`����k�l5�[����k�&�4N���H��٬�$�5�㽪zo1�1Wa6�v*V����w��=9�P6���+s�T���ޢI#�~
��K��t7"��-��-�xv罹�yo~6��|I'}|0D�N�dI:����a�y+�=��q׊�z�K`
HZk�0���	�M�����/9W���E~���D�{�j�H���I���+z+��iwFSs�w����e]�.�L[Ztzh&!W}gdK�)Z6�'�p&�f��3Y�����m�8��~�ӏn��m)p�u���	��#������a�����v��CM�Ov'�jqP��t/W!ykrЏi8�=�Yr��ζ�5k&MD�c�츫�D��@�x����b����(����sֽ����[��@�1�Ō=������Tק[[�l�)���p��9CB�ŝϮ�4^p����JT�*��3	Hҙ4>�Փ��i�OS̜pݠ�tQ�(ZӇ��~}~=��@Z������o�9̏@ �w�ֶҋ(�j�$z\~$�m�������-��R�i�k{���9�=CE�v�mI;��v�4H���!���{��Yf}z]�h���M�0��n��7�ﻭ� A7�5痯8�� f�� Q��tbT�Q�&��ˡ�Cd���O,6���-X d���Q >�=+��7���x�7���{�+m�Kn��'��ޞ� 8o�3��>�u��$�/|� ��l�F�����qna���9�ݣPR������ne��<Z�pGm�kU��El���(KM���Z�@ ��{��� 8k�ςË�G��[>�<�Nw��۽t���$��hb'B���7~�x_�PH��q��J��e<md��V���b?O���:&�/5*���^���`G��Y�Հ�y�wZ�� |��İ`/om_y{x�77��E�~IJ�-֎wnIP��5D�TI�hz�A�^��H w��u���9|��/!�J��:������'lP�{{�{�rI�ݎll@,���@ �{z��d�����=��ˈ��H'bv�==�a�$��^?]�5��w�sޒ|I�M����K>�x�2�`=���x��;�SLn{N��]/M�Wl\<ۛD�oP���N����m��m�R�3�h�����@c�2Nm_�.�h�OZ���z��齃�O<�6�Ka�-2���uH�[�����7Vbo� �inpJ� �Ͻ2M}�#*X:��N�wz�r�T2�e��ܘ�x~��_`|�g���r��[��Fn"��c���4�e�Oos�Q�c����w��_�B'676���ԍvNuj�F>�fHE����Du��`�<Ȁ3�G��J��t���o�^bv�s�ꩼڪ��sEo ���W_ E�}��;��r�w�k�Hz@�ҼW��z�O��"���  ������^+q�ʒ\��;�f` -���t�@��w�E��y��oar�c���b���]��0+e�D�gn��B�oc�$�(�<{�p;��� ����z��d�e�A��b��-��t�V��b�������^��B~$�}�w��I$��:$�3��r� X�yu^A������D�Y��v[$���]�u^�/���il s[�,�o��݀�wz� 
}��ݯI͒�)�4ګyTz�d�N�A �\�����ֶ 7��>}�^�,��;{rɬ�����h/1
��6�k�v(ec9��lu��4�<ɑ%�6ə,ξ�u8����5�`����{����wY�ǹ��߉m�}�8��3��+�t��WI ��*~$�J�^��Qה��!�,�Լ2�uض�Pq�ⲝqj�E��m�YzY%m��]��.tR�0�G=P�f3���T�{�v y�K�.U�\���'���߳���I",G������,�k�K��"I4I���'Ē@[��&Do���:了���T����Kn��%����0�r`�9弧2�ww�R��I��t`>*�����Q6�����S/�:��n1k�����Ѐh���)h��>��gK�?	+8�UB�����^;<�l��l�JÓ�M���\���=ˈ���w���j�s�ܙ��_;�5o�?3�?`�~�S�j(,_�a !Z~_� �~�����f��F͇?H`�d(cX�������>�'�kf}��,�C��41���5$! b�$ tX@�:���D�!~)��	C�3;��YP�,���>�0�����E�=!<��?�����i@���p=�Qrh�}y���!��;2C��������ჰ�&��/Ru�р��u��C�@ ��؇��������"I�� ������ HO�@��������?������]���?��?����C�O���h>���4��xH HN���U�x�>�""5!��?��`�>���"C�����?Hzԃ��SFB��s�!���?$>��:~?��{ܸG��� ;>�{k�\L?�;0���4� }̄$$(I�$��R�%�(h>
t���#�w����.��O�����I��U��T�~0>a>��g�k��?q��B��g��h>��L>��Hk����������x?���燯�7���}�e �_�,����?I���!��>�����l�S�����{�P�!����Ϸ�7�~�E�>rh'���G` �>$�����?�t}'� ����=���?x�D��4�O������e��BB!L�	 		�!�d���x��B~-�H}F ϓ��C�$������	���&ϖH!6�� �A'�b`~�H������	 ���,�'@$��}a�4Or��a�V�� ~`�B{�D�$�ܳ��I����t�d�`����d� ����>��?q�C��@B9�?O�I����~�����'�����!�D�����O��������#�G�D0?3�	��|��a�a�HL~p�d3�_W�;����	 		�����>o�/�!iH�����p`H HK'��o����C�@��x0�`~_��}>'�	��C���!���!�����Ɉ�`&���|�~��?w����C����~??�;�:'��������a !1���>���5��_�G�v�0�O��Q>��>_0�AŇ�|�����4C0
Ě$?C�B0!?��~�� ~Q���~����?Q���B}�}��O�l���>ﺓa�GaI;�u�ۈ�ѹ�"C��Iˇ�	Ϝ��.�p�!�d�