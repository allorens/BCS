BZh91AY&SYw	���y߀`q���&� ����bD^�   �}��*٢��`ֶ�m�B��Z�AJ���ƳY���ĭ5FkJ�*�B�����P#l�Ҷ�V�*�U�*���}�pe�Ke�қ*M6�Cf)�֍�m���[[R���&kem�,F����m,m�JT�B�ե�f��[VX5��F[k�I��z^�Z�Zƪ}���Ij��Ryu\�j�U���,#f��V�U��ahVF�ml��l3amUf�ZլM%mkP�X�$+f֦�m�m��՚����ZV�eBV�    ���w5vk�k�öt ��IWU76�r��N�].�%���iYۣv2��hs�F] ݗmڜ٥��!l�֥VM��-�HŶ�5��x   9�}�ۧIJ��e޹z�*�,q�E)'���J���{����(wx^�UTU\����R����<��k^��}��))}e�ݽ�JT�{�*�M�
f�L��Z%J��   ��|�F��g����R��_=�ޯ7f�UQ]�W�����9���v޲�9��G�=!*��﮾g^)y��N��駹{yꉬ�R��*;o{�N�kf�mR�Z������   ��ҥRJ�m���Um���;f&�����lP-x��R�[j�;ٽחV�2�7z��Tۮ�ҕ�.�)�{���=�{A{�۔5��{2^;ՖٙF�l��ѭVTڭV�  �����!#����Y+٥"�z��J�s���+x���E��ڮ<]6��9���ow��T�n�%9�Ǥ(
Wn�
I��O{��R�%*W�֊[,���[Y4��   6{꾎�dJ��.t�Mv�;޵{ԩR��ޗ��L�*^ǚ8\etԻm�YޡR�v�ox<z��R���w�� ���{Ǫ�Uٺ�u��*Uwn]�l�Y��J*�Vfm�d��  �������=*T%#����*R�{�w^=묥$��緼�KMM3z{^�J�!S�����mR�W����ίv:���C���޼�z� ��J��f�5�i��-[
1�  ��}4)En�sZ�������+���[���8z�Uzpz��3���z�F�޼q�]���w�R�gE�t��=�հe�5�e�mcP�Sf��   >�>�_^���]�u Vs��=
�]���E6�X�t	S�Ws�]4q�xQ�A<�w@��ܣ]��ю�h��OQ��mVm6��U��Z��   =�} �z�ր��s�UU���m�{�N�J��ǏZ�Awzz��������u����Z�=j���=t>     ��2�)D��F	�0&&&M4�S�R��FM4`� �i��14"����( 4  @ E?	�)UO� �    �@�����!&  ��i�`�)*jI��!��C���4�#��|����w�i�I�KS���9���;o��~�N#��_��Ǿߏ��6��]����� �|6�����m���ᱶ���m8�����/���<�cl��!U?���������?��}w�O�}?l�?l�,��Ck85���m��!�ɃY�� �Y@Ŝ`�,�ŝ�Y�&� �,�8ŝ� �mg,�k!���Y�;d�Y�8�q�&��d�Y� ����L�`���M���vس�k!�ɀ�m��k85���lp�,���,�ŜcYk b�6�q��`�,�g&�gv�� cY6��861d��,��&66������g�,�� b����lv��l��b�lY,�l91����8��d�m�8���,�1�8��0`����!�bɍ����Y� 96���mdƳ�YYY��Lk;�6����k;mgl��`�`,��1gm��q���md6���M���u�5�b�?Qf��3�]��~E����GNam!��[��T�B�H��J��/r����K!��SMCu�i�
���Q�0�~�B�;�5f&n12=��� �D����r�*ׂ���%m��c��S���vGCjK%�:�n�Ǫ&kd�ۙ�X�QD�7��u�$mi�Wb��ϴ�U������u� ��:��s0G[Z՚����	e+�B��j�[��ݔ���M��z�dW*�4s.��0�{a��QH(zL?2���(Q��d��:�;6]޻�Bg�سa}	W����4�t�ڴ.η{�\C��{*I�*�S���
�j�m`ԂK��������ph6/�M-j��[۰:���N�Xk{+��R�Xh=;�M<�$��Dy����Pڛ�J�1��Puae�a��Q�2X��Y�ժY�����otR̚##v8��|,�?��U�gM�q�����н�*��i�e��]dz���Ǌ<����H�]f�·*�����s�m����m�u�%c���n<�[��id{�19b��,�[�ZU�T���O~I�sjC�sq]��}Û���p�K�tF:5|~Yɐ����(R��V+�{�h�&f3/[�.�"�Ӎij�Z� ��&]�%�3�0�uV��}k�٧V4��qh���ihl�XzŒ�(5�Cv�k�ct�9��}e#�ԭ��ded�Y�y��\v)٢٣�ËQc�N����'sw>�{j	��W5�-����
7!N ڟ`N�G�RrR��*��eXЦ���Z*Ɠ7��V�ɂ��XZ��e�Z1�D�%��h#Yk3�)[O[	�}M��C;i�����ކ��1�a+
2���"�׏B�\�%9o[��[)e��kA��1m�kedyJp�U:T����k+]�h�?��ּycNkj�ER�ˋc
�i�S��(tcW2����6��������5.�H��H�⺰U���E��:�VK�z팉ڥ���Z��9�(I��H�=�?Kv顴����Ó~�Z��L��I�Y�5�5�aץ[�:>h��h�	6
�Z�{V��k(;��0��m�(��+N��0�<qY�<�B��;�@�4��^��ܧ�ʗ{L-sc-�F��Z7r�MF�(R0
EJ�v�<�/Y��*��Sv�^V1��yA�Zu����i��(Z�/�o��k^�I6�q�c�L��[����P�@ʕ� ͓M�˭Zp�M�0�aT��.��˷�a5���/E��	�*5�f��BU�G2)���j� 5���'�Q�x\ P��� ��0�l�[�a�[��WiZ[J�͘�ZWd��cJ6U�"n�1SY�Q���z-�����GfS����k]���F�J
�{���[6�-V^U��%�(���c�VH;���YL�̩Bڊ�Q�*I����vZ��=l�][�f5IѺЍ�[�G$t1Iu���LRi!)�*ݔKt�'D�4�X.��I��ݪ��T�Ym��h�K��R��g�l��#(+�U�����r^�a15�H��ӧ+�����[�[��3��yVݥ��Z����IC^�*!��7�\$�4�����i��oK��͢�E��둨�.V�[	EB̧�6SfDe���H�Z�����vS�#�*3��Q�ˢkH�%�D\V^ˤ��ۨq��u�SQ���2�[�v6m�/b���5��ߛNC��x�y*�p�|4��{Oh�����"��9�ɻR�����B�vc�!�4���e��6cSb�C,8iλ�t�Ha��ؠWY��+%Y����	��e�O&XQD�Y{i0um^�E�YN���o/Mm�Ua����7sU`x�f�YU�,^����2�#�r��X�^-J3���Vϒ� ��F�4�b�n6��B���WP2m=�$+3"�9�[�^\�1�oX�-B+���GYU��!��r-�TA���H�����z��<���	�� ���F�8�Ěo�K0�1�D���mV���3�J�e=BS���4�͛�Ū�un@bm�kX�b��Q͸e�V�f��w�Fj)�X�%e�kI���������:tN#y�&�㚩���eJ�X��Z��$��`U	.�&��݂�\kokZ�&K4�nʇq��&`	�B�JX��DC4	1��{a˲um�VQ�O�,�n��w�7d��$*V�[{Z�iz�����
�5�n��Q�bZܻ�+oXx>��Qz���3q�i��N��&]��e�z5�@�(��;��u�1�z^��4�M����`7W���m-K
ebV��j��f������5f�53w1=e�R��b4�5��s+A����+ǭ�Ӱ���ra#fY�[����H��4�m��3�z�kE�r����z^������i@*�$nm`B&	8r�p�����Vӕ��/��6�r�m�ř�Se���Y%f���e������n�������ǡ�Q�Ǚz�A�"�A�}˩֠��r��M�c�Hj���fX8n��sp�EJgMa�7tT�5?�6�2�P8m\KZIn�;%�ɔf}�(�{,�� Ûk$u�I�H�%�4p��Z��r�7o�f�Qm��Ү�ϑλ�K�PiwoU#W��/ Q{L�ە�����iX��ʍ��1�UwN�l�E-1�-��8�jݙ˱Gu1"�@h��n�ƒ���x&+�y����ϴ�J-��.Z:+ձ,���^�sE��M9�v_
*R��x��3/`L��3�Ah�Q�F�fܣ��/P-�%#�P�軲U�w���VޅZ�
�̉ٓu!i`����d���f1D�e]�C�EKtͫXf���k���Ʊ��l����Ӕ/(j�Be=��6ZR�̪�6:ڑA�$�e��B5��J�,8�!�E@��uL3��t�*4�9����V�b:��v��g��Q�a�S�@�0Se���o@*�:�n;R��<�ֱL�{����W�<���.��bnS��ق�0|,�wL"R	�t�ܖX��n��/ٔ�rjZ���Z�%fZNK7kS!��.���ƺ�J�,˹��8�6!�q"���b�Q����R�+I�QSib�;�+ë^i˺D�N����vB�"7��6��-�y��X�ecx�����x�;�
�c"�Q��B��������je���D��{�]K(Bwh�[���[�r���{Y�H����<� qmAy��R�#hk˫2T �N'yz���6,�Rw��%<I�"�E`�;�5��g7i]E�/�#����O�#�dsF�{Z�b�]iT0�Qā�ݬ$��;m>��M�����޴n�rmX e�(^�N$���Ex��ڼx���J�i�V �e�iښd�I�1Sxi�j�fQF�'7/Or��Bh���F^7�Rt�n�i��}��4��9�b�xZ�zڢ[L]
������{�5��������x���d�MQ7�(�.�I��@���v�@|��w�X�޶��	�+�y(�X���m��`���T]��ݰh�~dh�k���V��yX�ڣ���&�s�q<�h���)b1ޤmfK2V�́�V��V�Xެ���z�٣��E�ӊ��s226���J<�ɹX6�1��bp��b�t���V�+�ʝ�u3i�k�Pꕳ��X�h�i<�.kU���;E� �����U�b���.UXR�͇dА�uU�r��B��PbF�{6գ�Äe*Xܨ�wQ�ua�^����s�ߒreL�c�u��-ջ�"����ۋ�f6��\��(�6�n�� ��h:A1VF��I-%N��Q01�(1�%7WC~q��Ѣ�)[n�Ҩ\h �hY�Ea���D�m�lhP6U�5�6G��	��z5�YwM����N����hC*mmk� wkK^PjR9U���PƉ�s�S�#S+������T-�9�T�m��R�(`t�)%+G1����(�?jG��7]]�R��5��i�Ȯ�����¶��o�ں��Z[��$�%��V�r���#�6�=t���H�-�t헿lJ^
L*p椖�$J��z���VnRx�")l
O�q堖`�f��[�M�̩���-���yS6
�L8JvVU�8Ѹr�)�*�wj�1R��]�M���t�Ҫ:��A���Y�5��p-���IG$��1���[�=J�p�[��'����ɽ�i��;Q�si���(؋Dh+K\1��.R��V�Tg*͇��Q��6ۂ��[sUCM楋.���um�Yfn�N�`�wvMf:u��t�\%��K
�L�(����GּZV���\Z08�n57sp�kè�lh6�)�j�Z-CV��N��)33.՚�%dq��o ���1'{��լFKx�f�+`3ۼ��
�IS�
t4�i�JW�u&M��C/wU�R�!$�B��̣��S/q,��T/����$�[Ya)ۺ:rٶ��ۥO6�k×x�!���4U��Uxi��{yM�4m���@��tsessi�KTh�mu�,��5�i���5�!��#5o+6�<�F5k6�S3S�ul�[M2�m�/qMƮ�Ɔꖰ;�2]�xM:{�-��0$韮𽳭�l��R�����Q6�L��fVV��]:�������ͥ�DӸ�!��#do̭�A%��e��{x�ģ�3L����;D�W>�ɔ�.�U��e1a�����z�N<�Z�M슘����v�)Ol�y�h�و����,Y�Oh,Sn���';aںժ�3J�Bѥ�Nq�)L�(�˙�c�� 
���4�-���6	kF^�Ě�a��ȁ�اcKD䊃��	km��FZ�)�1P݊�IWS�i�v6�G1n��;��ر�����mT�֛I��E�~������ƕb�(���D�@u+p�0�x�V5q�7y�^�d�,R*�
�d�vR�ƣq8��-�9�X��Hh��[D����M��壴�9��5�b9r�b+�1e�4�I".�6�ZU��d7@3R��1XU�"�S�T�NKU�g6�T�����9���VE,;J��F쭨�֣�f�Z�W�q���������ֶ�(Ή����~�/��)��t�^ݑ��Z^� �
�R�7j�T�wh��Jol�Զ"�Ǣ� �]��e:{񕱘[W�|]-	n����]��tW".�f_�p�쭶.�R�JCA�|�	���9��.3��a96C���K�X���.��k��j5�R�7H���H��UJ�N���@�Zǅm̐�[�I�~M���5��)�-�۬��	�l���ʵ�!�nk�Em�]n�a=�K�P
�v3[i�c.Z�ї{wY����3
��H����m��<{c8��[{�#NN cN:F�]nj�j/�N�0D��w6nb��C�-^aWM��(]n3v5�9��F/��ڷ���Zm�&��[Y��;����K��4�A�r�e"��ًHk���j�2mn��#��@��e�$�"�t.�9��՜ń!����6�K�z��&�HOܭ�k��|��k&�v.*]��YRk�r���4�-�3u2�nI+ !i��c��n��&��H���3NS+3A?\����!���`ԝ#b���*�#�d��,d*��e�8���L.�Ƕ^��f��\ԣ�ۏB�i��YlbXz^LE�y[��7Z��4("���QzR�5,��8Dա��Q˭��tA��\ *r6���,](܌����+c'm�31��0����^�[Q��A�Dw�t�áި[����]nf�����Dg�d�i�{�юo��^�Qꥹ�����i2-o)+�1�-�0�b�(�z�0�.��U��4=qj7����ſ�F+9r�Ƃ��-�T���Lz�n���eh�R�q�7/1��Z��M���-m^��^�Q����t�`�oF�[Kn�����2`�si)pYp|)�d��8�,��昩��gW��r<2�I�ܬ`Q��`�V�y���$kdܵz�4,�,�����4y�l�$c@�<v7f�ާ�	 J�41�-�ѻ��ل�i{�*��Ct*ǹ�����GL	Ƶ�ً2-ƶ�ĳL�yj�[/�jơQ��V��5�J	cxHBF^sa6�B�iXROo���ȅ3��:�-,_*�����@���ݡRZZ.�5�����um�ϲ�̔��1�dSEXM��2����f=�R+1�DYj�1<G0�i�3tX�$��ҕz� ^�W�[A����UM*U)���k̉<���ZH�kC1\�Tǆ�V�[JS�%�rk�h�x�@r�M$ʗy�J�Osf�j��#(��)l�EA���꧛i,ٻ�+��	!���\P�m`Vmn^Edѹ��W�{E,��O�^��HaKqpP����Q%5��Ӂ�I��a��raH�XZ�T4�(���,;�M�u�E��j�T�M�"�uniz]���*y���4,�ٖ���M�#�i����J�O+~�u����[��M5r�e�)2i�<�t�˔I+����wf� Q*T�²����T������e�iAi�d�pA�Z�j���4��n4�կ̥u���
kπF�4�&�Jk�@�Vt�ϲ^��߄y`*�w��mB��j^�X�e�j!d%������t�3Vq����4��k�z�u�˾�P����2F���Fܭ��ϛR$uYk{@�_aʸ/�\�Y�Թ�A'M�,����,���g,mjι {�&�ea����,2٨Y<�,�#ʔ�����7��R�P�S��4���������镚:f:�\�7FC��j�'3�n�ݼtt^[e�3s �o������<"n�ye��r������#y�@?���0}���\:m
�O������V�WHEnjR�����en#k2ܘkB"�̻����p��wU�g��(KQm�H��ڎ�(�t�� �SS���������ڰ{�d�s�;��2ټ�#m�%[w�}C��yS��m��u��wRPۗ�>ޙ�[b�G����:��A�e�,������s"�C6Z
ݺ����@c�PT�N��J���շ͓/�ʐL}36�jo���*\�خ�l��*j�9X�Q=�1�J+w[�@Y!����h]c@9��ʹ��
�[���[�r�	�]�<���;�Je��d�!��`H�EQd`0�g�o溒��>r�{�ރ��1���}��H����Ã�ynS��\��.,��K]0��{��$7���C�[�ʧj�|@��k�-�S����3:�Չc��X�K�1wh5��^V,1�,u��3���ӹ�8V5�Vtk�;8���L��U����Em�[�>���,v�]�=W���MJN���K�v����]�K�9K>q�eC���a�Ez++	�16i�ף�ާ�������e:��>�]��]fZu�@�Z;Tqb�Y�&�ER�N6�Z�,5�n�r�S`�n/Vn�S��]ӧ��ʙ%�M�X]]Nř;ktD�:�#KPq�+���VL�gG��n�H�ҫӊ����@�sV/$��l�P�z�6a�J��D�MWcm�q�B�o�*-p��Y'��N�G��T�B�#dL��	�efmp��x���1/��d[���[�4d�:���N`�qK@���F=T��}Q2.�4�
%GK4�m���u5.�v��:�]���ɻ��^wT[ͱ�)Ʋ�K�wZ����j���5�)�9s}�Nױ���=�)Q&go�L� ��Tf�Ɵqՠ�k��E(��G$���bF��t4�U7C�(��6j�L�-%8��)s7|���/�B��9�YȀ�ɻ6�\9��ZM������hkھ��d���,0;t�d���j������b贵���$�Qt�)�R���V�|��'�����'t��}B�]�����{,���':x�*�YSqVUX��[յ��pR��Ļ�K��{I��R�ekUj��\,�pL��d��b� �S/����ۧz�Jޮ�1l3��K�ݦ��9e���:�ջ
<NQ{$���7Hu4m-%}��ZH�[����na�����I��y1��uT��U��d�}/z"V�n�ׁ�^�2{��t�J�J]�5M�R�H1�y��*xZ�t��֍qk�
� �Y�r��n)�g��[��ک����6��;�H+ϕ��H����.ug�j��#̝�.hŤ0kYN�K��5�VF����k2��K�嶯����6���\�l���W�qo&�,X`�w�	oi�ޔ����)6/k��w)�T�x�Sot�=�����8�j-j�����uע8��z�a��[b��{w������w1��j;�j��ȍ���&ݑ[�pA)"ꥍ�k �[h���y�cY]P�j�.f!O��-��̠P�H�)��ݴ�S#��GX�F�Dtn�{�d�W��e�wX�7J��	�1TksLU2�j�&Hm�eY���_s��]>-ץmm�'�	��f��q��\;����P���#��B��2 Z�C�Ös��Ii���طA�>�Bz2ً3aGJ��v�\ݑ�:O�]���XP��e��g4�dr
w�y��{M�U
ׂ�;��,���J.g����z�Z����vj@�'z�{ܲ]�Gi�ҭ�Uǭ�=���Cg��5��;q~s�e9�8�R՗���["���ݑ1�<1K�Hrl�DNE�fX����'u��m�ʶw$H��zo9��WH���]f�C,��2�����P�jZ��n��	!
ئ��p��c�d�1h0�YzJQr��bܬ�Sc��;��S�=��%"�}�N����Nr}׎:��Ŏ�!��Gi��m�z�ڋ���t�h��2^�$b��
o����s�B�-����ƺ�/�*8��F�&�1��^Q�Є���O)d�=�Q$4��7Yyն���&�7\\W�[���u�
��/wWm-��mҧy�8]��#��w��`n�sx�og?�����!7�MU�������(��u�WK���q2���}��I�q���`։��)�c��^Ṳ����Ű�� �ed)��c5a���,޲H�:�sI�2��X�\�8�ʛ�Z�kGj���`|�#�Aq� iN��ő�-S<�ڸ���f���q�Z�+`bܔ��/rɀevD�T޳A�nht2��j�\��k����.Zuf�R�Z�S��U�t�1��{#�]*������t�<�[\�UdF2��	�ޅ��=��w%�kU-r��In0m+}�����mS^� ޟ�p��#���I`�(���ח�M2��m�nK{�Sv�'Z���ҳSh�^��v��2��$wG(f�ݓx�;���K��z���V�η�S��^s�����Z�h�v�ʛc5f�_%��dV��DsR��եӗ9&.-�!�j����RU*渍v�0�s�h꺵%���D���T��BZ6o�����Y�lg ��%r��w4���0K���8��{(f�ba�U�e�Զ��V�k�]��0&��z�ɸ��8���P5M�u�f�-<.����]��O����MS��ON�('�76eY��6��/b�3�ȴ�v;��m�rh���������2`v�v�r*�R�ep9,�C�m����T�:g���o�ߪh
��V5i+
�,�'����h�6@�x�M�Vb����]`ɱuT!tN�d&�[3L\�uБ'��J̼SHZ;1��b�V��{�HUI}���Ѧ�DMK�85���^={y�Ƴ�.-�x)u��U� V�i8��F�&H��7���y�jڽg^l�3]&���{7j���+,�WR�y����o*�p��nek�R3k�,��yv� }s�'hAe�ܽ��Q�ͼ��*�$�e�ǎ��-�J@Ė��J���[]8��S�SGa�.����sGL���R�B$1k8'�Ci�����.aw�iؖ�c%�k.N0_U��2�*�S��a�7����.L�3&���o���MP��m��,tT�#�e�!*Yq���n\�^�����A�.����W��v0�{1z����<������d�n�`l�o1%%zS��>Új��p��'eE�����	Y	�[�Ĕ�n�v�*ݴĵ�&��Ѧ%����n^��u.�����W]]�n�����#3��nF�`�0��*J~� �ߪ�������S����Oy�Y�i��M�)�:N��\`�/�[e��F<�Q)�
�i�'8i�gD�]؝	ۥm�n�*]3RE��[Zy	/��}u�YY�=Ύ]Lnfm�T���!ˌT�[�B�9��ז�ɹ���X�Q�n;�x�ypg҄B�	�.�Bs�oK�����k�v]vK�a1]Kmu-;����%m.��u}һeKJ���󠤣m�ۉ5���DI�κ�WE"2��GWnb�;���m�����@���F�����˾��q}��\��1-�݋>`�޾:ѳm����I��T���G�e��áR�1q<kCh��4̵�(��d$��t��s�j�f��'�7��shY��U鴲^3���ݫQ
�쥤$�ۃ�o<޶���{ee(͝fjGp�K�5u�ֱ��v_'YIA�r�cm��^;h�J��?�K�k���dzp:��@]�yJ�'�p��=�c0��U��jՕW]2����Ȗ{ggK�H�J��ս5���ղ�w�;ov��;��Uv*&��S�����j]�3rC�X$�h$&�;�:e`P����N��Zp���y�U�M��uH�¶�)͍V ^�Y�Vt]���̗b�F?�Yx�S/J���I3���We�Y��I+���D�`�OL�K�)U�i.��]y��Sz�,mR{`�粝��tGss0�s�Q^҃]A]�fV�1pAL|�8�u+sԃRt����tRc]]ur�b��,S�J�鷹�q�����t���p6�dY��1<��dy\*}���5��nV�!s�l�+�$F@,m?������Xi��+sZ����]i�;&Q`d�>���j�JGy۶7��w9�ͺ������f�V���t1�kx�GE���1��ĆXA%]�=�����X-�Ƅ�:ogl�B��-�و�̮��6-ۥ���T�P�bZ�{j��	��v�\�4NX�;:oX��V)]�*sn�rQ�N�S���^}y�#�
q��,�)<�l��u�g��"TAEI����!�ً:��Mt�(�t���]n����oX����([n�E�� ]�[c���fQ<d��w13�mv�k{�J9m�I
XqU�k�e��s3Yb�:��]�����n�X�V�F5����i�\��p�0�D�}��]������톛{��%3#���YH.¦�]ct�WFZ��2n��N�t��E!*o�m�b�eK��W:�7{0�o��Z����re��z�I�u�lW��"�R��&��h^`���E�^Ř��/-���s1U�DH9�"��Ʋ�v��J���[�e%z"��s�
����*�׬+a�T�FY�ކ�p��/�W�Ž:�lZ��Y�[t��ٔ�_e��Z�#x�nr���.�5��kt�0z<�.�9q[�u.���eq�{�A�r��nd#-vm�DkI����{�Ku�	�����*��U��a:�Խ�tXV���gV���N��ѹ�����r��M��"Cg�M��R�j]�:��lW"�e��:z���Ÿ�nk�\Mt�l�^r�GS���b�mdʼ��x���k�*K(�C\3��r�̺1<�]w���gה�k����Il�@��e�u�إ�O�巩A�%�j�gawW�(b�Xn%�����d���nĔ-Χ��z�Rۮmn��������{r�o�
%#�z��(��wyDd�k:V6�j�|��X�4��X�#x�	�6�}V*��3ٰ3�m�ʋe�l�W/��������$;^.[�u�W)���1�w$�I��WU���m�@񬅝�(��1�o�N
�G!�\��oW#ݼ-vt���;su��Ϋ�IY[V�l�DոX8���n�oW�٢�w"�1�����������i*aU4�����IoW&Vs&F ���up��ז^��Kn�U�o�����.��rĆ�5MeDԥF��έj�]Yq<Ht6��睴S.�t�R����u֤��<��5�5ĩ��m�ieh�t��7�F�QH�����y"�]��kBwR(�n����f�:�n�N5h3���7� ,!����d�)G�fA��L��P�Qg�6f�QO��}��'�v�亵b�3ӡ|2f���u`�~�}���
�	Q墶��9�5b魰�n�I�^�lg:��-1����)\]�;r���`у\��j�W۪��4�[ZY�MB�-�r�s7�t���T_.�*���@����o3d&�vR����)��!.�W-�3Z�*�<tB��N��)CX	�:�.���T�vF�Q�B��={��tU�{�L�y:�n��9� T6#Ƈn�Pǟm�i���i\�,�W9Fu�*�;ԛt+p���2���S6���Y���|��ֶQ%4j�ܦ
z9v��Su�'*-Cе��eq��{34[�:�[��V�@��c���ybCR����}�i�-�fg>M�AH�P����Q�w�C"��+Ntፅۋ��E��)�/m����Jˬ=e��2C�i׳sr�=�8/!"z�eNogW�f-*n�f�f�x�7$��r�a�T��ws�Eٚ4��ٮm��;B`��LU:�,k�$�^��6#��fV+�Y���2�q�8�ޫ�g@��O3�5���D����N�,��0���N����g���h`����o�2��(�=Z����4�2�����ZYƣ���:2�rj�^f�>3!Qn���9���\��h-��_j�#�\���5u�՛:nNgZ�5��Uԯ4C�us��VBR-�IV8�����
B�oeظ'y�1]Ǖ%>2bJ�z@���^tR�`#6�������'��40:��J��6h���Ws��k��ql4���Kɍ�;t��p����ۥk$�e�h�n���toZ]��S�e�naB�Wd�p㭭�Ռrhj��͘ʱ.��*���N����pVU�8�����P��v����9�h�����N;}���ϝ^N	��n��a֭-�K��pw#�xsGwr)P����:�:5��,��{ͬ�{h%}�Wp�)�ųR��`��/:>F�F��%�}|�E��cE��g=��B�έ18�Sb �/��s)m+�}XOd�L�]m���2�Ӧ�Oڏp��:��{'7N����'i���:{�;fhx�Zyx��(��
�뭓rw9��e�0N�he�⹭�^]kǑ�r�Ώ��ٽ8�j�n25.��?!�����R�vt٥��'9�z䰳b��kU:�S6�w{!�v(g1�H��ٜy-�"�C�mtg�ѝ���g;%�c���}I�t�T�u�f6�˸�|���1�2��n���@Qd��`Gsky�	6��V�9[Dk�wK��W
��ԼM�[7:����^u)��V��Q�m�7���󾚬�bM�]q�{m�%+x�9|���=���DнT>)P! ��F�e�6�,���l=Łʋ�@5�(�@�t�H���V����#�Si�v��ر
#X�ʻ�wzζ�ݫ���=֩��ƃ�l0U��D��q�EEDY�KB�6�w�1���?q����� ���G��>�����y������?����Y�W��_s����i��=.�Qf�'MpcbF�t��ikղ�}����uB�$��;Axo+�I1֙[����r�dTܷ�.���k�I�\�^ޜИ=G�g�r�]���r࣢�V�,�E�W���Rܹ��5��'Ùc [n��V,�)ˏj�j5P��\�έ�����A+U�O"���眫���l�W�=��i�-��f�(�Y]:�Jp2k���A��"qX̝+�w��G�%L�Ockg+�I���uGf�h޻�v��.�5k�s�u�� �n�詫P�_��+s����d�9�h����X�K?�Uh�������K��c����uXAI��2qu���]���wEN��u|�B� �::���yj�&�6�h��-v���9�e�A����{X��e�w�Tz[�ics�߲�TGL�FJ���l��83
�1�a)c0���J�Ȭ�]ʮ�f��ZKsm�Զ�]e)E6��Ϲ��x��Mԅ<;��y+c�Q��������'Zˣ2U������ڎ��V�;�. ������˩���9�,�����u��WTKMA��:gS��
U�G���jV&�,�tP�}��6��b؂X�����R�b�����(�l_j�l�[r�UØlR�0��A�2�
���\��#6��[�n��_f�QP�:4����;X̊�^�>�O������}>�O���=��w����{���p�{���w�����}��o�����}��o�����}��o������}�O�����G�ā� *���Ē��z"�:����F�x���������|��6j����ˊ��l�肕��o;Mip|.�I0:4z��Ĝ�s:�.�]AY�������r��`ܭ��E�&�cI�]PD{�!� i�2���mΊ��{�E�O��]�T�3j���5��B�	5Ǣj�L9�M�`i3UK�\��EU��ޱ��ol�sS:�r"���ǝ0.6��}�wH����t޽��G�;OA��@��{bԧ���mvZx�=Q��s���ȗB�m8F܎��|��`T�,67p������u��]�˷v��@�*=�A"e����eCG#ǳ9���;�4�-Y�c�T��m�����kܪk�-v榋�b���u!R�l�f���Az�r�,��.	ֺ�����ٝ��D�r�����e�S�P�S�������Vk�b�)���Aи���5�!v��5�M}R��%QT��c��o��h=�	���W";��wV��;ep�cHv��/�c�n�Eh����p�Q�n�g�֮�[��M�}F�Fnh�B;��f��K��qa��.M�-�f����U�%�l�V��-ݧ��}�:�l^Jaf۵�g[�E�s�Km��?��%vmˮs�TNo*�
D�L��j;;X�1���V�d.W�����o�5�,�N������~����/��������w����{���w����{�>�w�����}>�O�{���w����{�����{���w�����}>�O���oM�!��[�;�A��yز�µȖn�67��qЄ�VV֝k#ϕ#`u��cm4�}��&r����K!s]�ADm���`U3h1�Amun��4З�wX���
���p�A�y	&��ʛ!݁���S�;9� ܑB��C�-Qh�_G���r��ob��l$���m����\�}�+�ק�Ҕ��>��jc�ݠT2;ݼa�.]V�Gf*�n���F��qE��g@Nb�����ՓGRq	];�o3U���mICk�p�CW���|A�+@ҫ��>J�D�*7FB�����������E,��|n�f.��j��y��כ��ѳ������؁�\#t����� �᳍�1޵����>�M��%I+:0Y��_�>76�*,j�=�o6�جp`�4�6�U�PT�%��Y�+{fe'�f����L�}jE:6��\�J��&Kyܰzr˨�&�;�
����E��*6$&��5X1��dк)�g'x�/F��ަ��l��_J�~Uq(z4�W\f,|42��KX|���LA�۫&$B^��3�;�|�W;]�Ʀ����n�)�p�dv���^��G�yh�n��y��W5eoEV]7�-���Iy��F� ���[���{�t��{,T�<k�:�L��s����=w��f�G;�����ޮs}iWv+��"(١��tP̫qR�g����]�Z_R.��C�U�Q����`�)"����E��#(]3��[���xpά��.����io);�hP�"�Ṯ��yˤ��Ҡɗq�kZ�h���{T��7('���isGv
�R���{i��{.��+��WY����ĕָ�y�a���Bq+�����zJ�$�r��;���g�/�{*B¤+:��f%�G�Ss$�IVպh-�7n�qС�@�@e9�=�̢Z5�#˖^�v�����ӨvmXX���1t���ìvb����w���NF�cw�ΫY�ڮ��&w=�ɥ#��b��I"LG��+�_;��Z )�S�|�Lu�u8D�aC��r�`R�d.5�Mꜷ�K�]�����^�Z�D�Kv*TЊ���T�
0�5UqUn��U�Xo��Csc��K�	�@��_����Q8��Ꭶ�!j�i�w�fZ@c7��wp���	`��]C�����_V��*ّ��1���eiU�C\����T���)u-�XuS9h
|��7V���w�uX�:��s}���Nv�לJ�P�>����$6i��s�y� :hݵ��'yұ|�`�o/r:Fˊ��[�yfE�U�S%��%�]��I��:�����w}}X�@5���SV��ՐX"��d�ԫ+o
0��y�����ջ\��N�K��NN&+��M,�X��	�x抏f⼷x7�\� _be��;&b��se�xP2�q�1}|��o#n�@J4�T�vo���i���k�-�q������4�uf�E�z��֚��r��%Wduz�w\W]�L�*ml&��G�X9�z)���{���cnX�#��Ejb�f��XP���;\�4ر1������7U�8�5�iv�&C�u�z$HZԽ;w��UBi������T�]�9u����Hl�iC��Z�#���t�P��c��\�X9���f���&���(g�*$���WpPd�����Y��ҴZu)�X��'��ɶr��fݭp�|zΧf��μW�f�rj���������,�=��Nr!��9�d��Fޢ.��ioo��/*'y��B��7(\�+�c�w�1�JN:����Iջ��8쓊���G8�+w)w"�Hx1q�4�4�2
�-b��[H��5`r�z$��Y��L��w?����H�EU�F���]ec71,m6sw�>R�'��;��ŗbH�c�b��4�o@�A} �l�L�t�9��feY���\|�OWi;A�m�K���.=�Ԓ����"�tP�ڭ�����JG���O�	h�wٲ�dyv������d�v��|ݿ�h�s��>�(wA8{��-Vw:͵�X�C�k	t�Ǆ��Ef� ���hΎ>�o��*�rbӛLm���hu�̀D-QV/���Kh�Y�Y�c�s�j���ڈ��Р3^�ڰ���\�D:�
#�sv�h�K-��:-:j���e��kfY�){�[0���J9�3kt��t\�����,�֮
�:O���I{@m�R�k78N�;�ҩ���h��>��J��Z�,�"�k6u�Qh`h{���9v��Ky�I�kL��H���,�4� s�j-G>�`R�%��w�U���@�-Ҿ.ٚ�C�KOi�%b����9|��z�8�Ф!���Q��;B�kqޫ��S�P���i�����HɎ��\Ƭ�j��Bhwp��r��7M�o�qTR���^��f�P+E�r��&LŪ�鮟4�v%���ӎ����f���	�ֹܺTc��ׄN"��i-�=�&*a����%�6�D�5�
Q�,�:�)�YR������]Z�44�ҝ\����!tӺY]Rt2��4��kj�ˣ�m�'���H���ѷ��+R�y]A��6�ѠB�s�-f��:�j������=�:Mw���<WMƙ��x.���`�X	U͓en�qt��c:�IgEJ���>�mt�D] �F�����zc�;:���!Y���[�Gnq�1Zc��V�Yu"�f�`�U����h���9K{�Z���͉����+^�ٛ|H�^:jڛZ@��F5��.��	}l��N���7��<�A�m��a�����(���a�x��%Ky��+NM�2�j�i괲��d�*�hd啭K\$��<��#�}tzӽ@gB'���*�5� ���4��� 5����]��@Μ�Tj��R�%p�k�$U��M�Z�k5�F7�M�l^%gV��Z��Ɔ���6�����b�'�	{Hq��S����!��&c��Z��I���C�[s;��KWݯ�yIo"�nWU���s�,饂���m�A`n�������LG7w9�'Z:�aO�Me��L��������cܥ0��\�㊦X��r�sٙ+k�\�,��9;��&�f/U֨�U�t�ݫ���M��v� -�u����]S���NCR:ec�}�1L�5oM��4r4�̈�G$�5X�j�yċۥ%�E�9-�'1�֊{��`�)����h��ڞ=�[z ��d���7ip��yl��;ֆ1�qR��b�}'�Iْ�]vg�]�-��[DP�V��phc�\[�e���G�*��j*
��+�z�y�#���;ąpq(�X�Аu#Z`��|kB�ÝμIt��o7ǈKf�d0�9���T�x����}9Z�ݒ����xf>f�cX6�~�G-
ڏ�J�|N������"��c3���Y��:�$��e��ܻRǩ>�.�n5R���@ka�_ugX{W`5�}v�*yi:j��]u
ie���n� ��j�E�G�H��ǻ E�Ƿfޠ:Nްo/������vy����H�����B�x�+�N���#�U�e��mÜЮN�Vs۵���G]'Xk�Jms�).�^[<�-Q���.���n�YM�l�����ST�ڒrJ��ç}�����j����c*�֭��@:0�07�<�O3�fїZWZ�������Skz�uu�5�W7Q�k�g�(�d�w��l�����+l֕���|bqs�N��x��o����:wd%����8z�����}���T�f��� ��N.�ŋ��o�+,�bG�{i��u������X� ����U⥙X��5�C��|�Ka�ID+�.��e�+�Z�q�L����N��.,�`f����i�ۧse���#�阆����ٰM��
������cn�~� Tl�6�6�j���U,�mvrc��x����4*�S9��v&i'GC�\E�u����d<8�#K�6�X�r`��W��Xu�<�#�w�a�]v�Б��U|�������\u�ͅ_;97cgnm�+Bȥf^2�ꏍv;{z&lK��7B(�����D�d��3Z�\��7�.$�;��$��$܎K�4��4��pYII����t�x����P��8j�/��"�p2�ӊ�*�N�T�AKkhqͰyȻ���p|oft2:��>��ˎ�&w&�TF@X����az.�/���ƀ����tVrvgA���������WV�9Pv�C��kt���o3%��,����f8�t�G{z���i1�%1���T˂L@a�lM<�K�L���Z4��ͪ���������1Y���yY\2�v�JT�K�l���ϗD��!l���nūI\<���r����c����;S�v�/k
6 CH��z� tc:s#�H����R�G���B�4�Ħ�u�6�y����B}h��s�g���B�3X+d�T�;z�n�pj������4J���E�oY�)]u���6�/�];L��=�V��r@#0��a��Y�j��B�F4�i�*�*�	<�Զ��0��&a��s�V��Lu�i<�k�f^�|Q��*cjQ��7�	�ʋ*'3����G ��R�R��W�,�����pnq峂��q�r��.������p�9\G�pS�f�����$�/t�7��,^�D�飚��	5wx�������i�.��ɴ���)����'�2%��������G�M�R�;b��<ox�f�v#���`�څ̠�n�eo�v�\���T�9]I�:�WQNE�}�lM�wT�6�u�Tc�Q�4�����O��u:��"��;#o��[���vE�+`qũ�;͠{�5J+Tc�V�|�$�f�ok�"F�ȃ�T@��b������0ޙ�Y��:��1�]B)F8&j��7��T�n����z�X��:���䛡
�Y]�n�R�n0�����<��Y��=�ql<�w�����ӦMsܮ4��1�����Ce��E_�j]Nj��Y\h�:��J:�2�U�;��ݜTs+�īo���&�2��+�7)���⤖���&�KX�q��j&���p��R�4W4�e�[��[Ar���� �u�I���8�Ǜ��l�]}q%]�VƲ^������Gk��s�İ3�J����#1�c�O,�d����VYw]��"C���X{sn�^�ЏF�x:,5�XR5�7sjM%�Q�	�Q��.^Wp�jD�s�z�������3����BU��N���B�nL����Fm�T���5�|���ζ��;R���Iw�Qu��Y���[���ݱ��:�%�
�]�T�Y�NѮ,��ό�ܒ�GN�d�|B趑u�\JDT��%�ܒ�B�橊i��e���ur�l����Vd
A��Wk#�K�Ą�;�e�k,bIaf���b�5�
	���˘�tO,�C/z@P16[��"�,�����˳r�.�Т[��uλ7��t4=e�W���!.1ɝ(�Nl}%� �>�c+X�f�ė۴�\����E.�3xkZ�������&�&`�OM�������u�������������������{����{�� }_(wx�%�|�������Wצp}���s��;Y���tN�N�Bbe'�_��6'tZ��d��ڶ&VlS�v�6�g���|y���D;n^B���\IF��
�Z���$k\G.D�d'�^��#%l�>�E��ք���fE��O�u�.tW�S)�D77FG�'L���%�.�%�ܸ�Tˣ������\�©���˙�`��9M����k1�U��4u`7�.�[}� m����w�;�=b���6��v�,�yA��Щ�|�\v`ah(��C3����T��Ϥ���m���-){!�2�!��Y��(�����]�5�v�B��d�tA-fv:�l�E}0��5���h
�S��\bN�X%����î:���ײ���4��yw ׉��Ue�K�{����ô��so���9��Y���
�v�Ȇ�Z�J'��e�Oq�[�(��*���^��M�xAVoV�c�4�i]���s���0>�=���sSZ7l:|���ĺ�i�27�Q�����)�=Yku.�x��[W��w-�+rSE�
�i9FQs'�L������sDx���P�;���z۫����%�N�.▜oo"l#ۮ���[�G`囉A��7�T��m�����d�̭�)*ەe�}R�k6"��.��Ah�3��dJ��5��n���n�����d����U�B]p��VT�{�����S��̢��I��r)A��Ǌ�7���m��7��}_��Z)�/R��nhd|�G�Tz�G=�Y�$�(��Ŗw<L�
�[�oo����o��r�AQ8g4Gw��+�E��J��r�#���/
ᴗ��'�{p�U�+i2슼�qCA*(�
�b�ww(�(�G�%����(Q/�\򈪋�iDD_Y�]T�uݳ�As��qɔ���h������S��T�**���M�W�]�b��M�_�:��\����S���^_G���ϕ���\H�s^�y)��Օ=���������F㈒���a&p��I �P'^�:�^�'xb}"�c���Eyϻ��b�
�EE�<���{��W�dE̤���OQ:\�"�T\��ؑ��֜����=�PU	˔QE��s#(��Yϯ!ϙ�9��Q�l�:{���EC�v��r�=G��9Urap�e�^g�J���8��9�vE��_w_l~;�?���g�����Nõ\�&5s�w�J�l=;v��FR�+��;ف�S-��O���ȋ�E�uO:Y��w����;����У�: ��	��**�oR2��	�:oo����G��??�;�M�x�O{mx|��Y����b<ʴ��0sܩ\�$>����=�썟k�>��r�T��Ĳ�v����������1�|ؓ>Տ����t�,�S>fH}9W���û}ȧ�z]�,m�wgym��~��6�pr_�<�W�j���|j0�.g���_J��Op�Nr�����W��vW��zvi��}\Ղ���1��a�^��m�����4g	׶�����<KA�;�I�� ������>�N��y����s�����QU3ؽ��>��I�������k}���\��h�|�m�jy���;���z��{U��a��a; Q�3�;�,���SoT^��AR^1�8�T��J�2�<�U]�>���of�n��xy�Ej��V]���<#)V��^�e�WTʀ�3_�>�R�IрV_�&p��z��ItZ�Zh,�v�O0UՍ�RJ�m�̤M�/�m�F;,�\��m�T�q
v��hL�/^�]����渺7���X��Y|�<�F�Y%�����L�+wI�2Es04�U/K�[g��yd��������qQF����ʺ�Ds��Z�g���n�x���et��(�<�c�Fs�K4������W^�uY8�>�������x�G\���_>sH'�I�3���{ 8��c�o�X۳Yx8�Dݐn8s���0;wy�q��.L�y�@&�O����6@g�3���bks�<���g`��}�9�u�H�f����{Sz״�MQ�]�a��9(͆�j�4l5� mNY��/�s�/C�+���=�oe�h�=�a0�zh7� �I�ыѮ�ґ�}���������=�<)z�nJgE���Z�cg=��c���{%Z�����g|g7����7o�Z�ꋾ�A���Ȭ&������=��
`ܹ���s�n��.�I���Dwp�܀9��8밙�<�?KǛ�e��(�ҳAx.M�ǻ�8_3X��V?k.�D�[���A�t�4�T��ul��Uҧ+,�q�+���}b��Z^w��.����9���Yq�:�+��Ǆ�g�`�;���#�����n�M4����4����Y<�+'�on�;�#:�����ի�w&k��<}��o]�I��q�Z�Uw{��`4=�-�>k<*���+���w�wO�����G��ޟ_Ե�t��˞��/�e�������n5�c�;���:}[�V����l�ӹ:��>�T�.��N��e��J���Kg�ֺ���eQ�/��3�繎��nkW�5�	��B]�M�9]�݇���n}&<�!������?L\�G�X6|�� ��m\�����#ߪy�zc���{-�{�C�����
��9GؠN���:��x�)=]�j5P�^�����^���T���7��ݛ=�~ً�.K*�Á���}u�{>���s�p�v��xO�[z����J5筷�-��,r�x��T��^�ꜭR"�3x:�z����n��jR^����_M�x�{����������*�g_Oe^v�j�M��ŷft�^zo]�زf�ƣ����㵢 �MsҎ����1����(���6��ѭSˎ�	4�^��6�qm,Z���Y,
9WX�h��{��wRޯ&d^��u�^N)�a��u}�����yw1�3h���w�)+Z��*δ)]G�V]1�0Y���t�OC��L�eO���y�o�7Z��E����1���<5����:�xD�����ח��}��o�U=	�C�RA�w�*f��pl]���hɨi7�n3sϰo���Y���ܛ*z���7�%�X��ݕ�A�z��#�Epʲݞ�����=�TO�eD�޼?kpQ�~]�v���/`cAw>}��p;>�|(n�����/'t���j�"��n��j�	��'{6�y����3�*�Si_�t�Ҟ6�+�}M�)�K�s>Xw{���V���zic�b>����[��W�^Iu�*Y�h�z>�_�$
4w�q���;աd@Dy2�qY��O�%�fr͊9�ư'��g[�Qݺ�7ӄ[l��EV]��Vi�s��m�ߐ��e\b�oOwa�by�������M���9��;WdR���S��k�e�]��`�V�ٺ��ѱGt Cv�-e��%��b�Yr���WF�:H}W�W�9a��3�+�ٚٺ�}iƁ�ӓ��]���އwq��@��n�|��׹'9��*��#s�E[c7e���C.AJӼ���^�=P��sB�0:��� !������.[��Ʋ�C�R��nzc�<��}QX��9lgB:��L�Ԫ�խx�=�.z��h����Ѥj����L��T<��j�x[����}I.o(�ďzW���ǜ���}6���1!���f}W�=��l��v�D;9���z�����#��ώ��&�*��>{c|:l��BBj�ᚴ�泥>�����<|ޞ��=�^���/p^�/b'�T@f1�_��?+=~y��3�/�\WZ��Y�X�z�S��}��y6F��@s��x��a�*?W��/w��9�M��TXq����7^<A���;B��o>��+ڻ���$o;�z u#-o�:��u��|����R_�� �uõ���i&��}���4@&�k��7-S�y��>�mN����j�S�&����}mO�S�X��d�߉���mz:�'�C
�K6G�������'��n�;]�^~x����e}��y�ߥZ�w�� ԝ��?lH]tC,f,+Z�Z��{�}�k�ؗ>��,�u4y���U�n@�g^��L!k���n�I0���ڶ��0�G��N�hÕf�l��تVqܷQM��6G06�u����U{Zs�@-?IR�=���w	7��G�gd3��Q=��&M�CukJh��^�U���}���I��=;��R�������s��L&rѹ�x�ݛ���j얆1�ݛ"c#�g��^�&'�u���9`�Q�Y�(3����w�x�
�_�WK*�1Qλ~ʾĨ����+=�[C|�7�'F�o����_�{cG���(��^�WO�_�} ��uX�;�9ݍɩ��ק+����C���>��K��6���i�WL��@�l���Gˢ���H(�>�h{W����=�LI!��eŻx�6ߍ�5�3����"J��^��"Ř�ƍ҃چ,�A���F`�!\o�G�ss��{W{F���q�������(�}Ɯޮ��"��VD@��`��xm���W17H��e�3����y&�����W��g��7��vDU�S��b����*����{7�vdݥ	��ỉ"{"�f��՘-�r$ZB��r.��%����.��N���{d�)��Oeo@�}�a'5�h��;��c�I2*�]K:P���W�yp���ri��6��cVj�fZ����
��+�b�ꌊ�z��)w��'�uzY}B%�<�[E�<�����LY��s��2�;�������j�k���څ{��x�o���{��>�ڽ���4¯y�뽙g�0z*�>�A�v��n����s�V�Vv��}K�Nze	~�立�y�?�ڜ�=w����A�5Fe�v��^��������e̋oǨ74�̱Ƿ����y1���7��̮w�y�=��V���Tr�;	c�� ���uh>���5���,�X������u�+B�9e�ϳ��9�����Π�g����܄��A<wHv�t3d{; 9�w���y�q�׈5��OW�ٲI���g|��[�z�I�G��pW�կ�k����GL�rq�K�ÒO^P�ͯ�7�ޔ7�]j��3ʑ#ӥ�K��<��W(�¢����[��y�w�y���JU�m�w�����#��-F]b�yOz�D��~�~�0dB�5����wLѴs�-�{���\%Khh.��8��3Rx4�D��{/ q>�;��@�Z�6�̹�k�h�-hԛ�86Υ�h-��i'aJ�W�ﮟ<�w_5�����q���>hM��H�xj�^����_�{�mk{Ə�� =�5'���ݧҞ�C�e8;�J�c;�̊��k�8�O���nz���Y>T���~�;����������J�~�~oޫ�M*�kP#6��z�Ό0�G�WS�9s5���]){�:3����Ԏ}$����Y���P���>�WO�y����)۱n�����y;��|�y�_���]ѿ��:��P�k�_c{���_��^�)/\U��i��`�����.��'���2t�M�o(�=���˻���=�Y�רUi�����io���J����ߪ����9�-��<0���'k�[�u�����C.�u�pvU��JR��~o�u���m9���e�L����s�Ww�9�]��0{�)un����^����X�z.�'�6;n��2�}9�*l����{/�ۆ����y�[�a6�Z�6����|s$Y`U��;�ʙ{�z�����,㽥9� rt�����"T�v/co:5���Xz�k������$�A��W8&���wt��E�2��ت囫7t~9ԝ�"�y>���w���h����p�#��*Ϟ_� �6����V�%%��%/w�Y[7�jzG�z�.����C��V��Z׽���k$��~l��үw�������9�۠M���ޟw����kth��
.lp�jp��z���{�ߤջ���'����o��-Lw�p���d��r�c�h��0�[5'�l���כ�!�S\l7$��iLsw�9�]���eʧJ
X=��k˶��$���R����a��um�5̈́8�;�@d�=Q�C'
"�◧;۽^Wj���]@����.�7�I���^�j{)y�a�Eb�Ǳ���
����3k��P��^.�Iy�Vk��J�̥���E��Ƚ@�>��9�|b^J��v�g���;���ػ�L���b���Le0�|:�(�V�9��){A*��Z�Ɛ��w��cn	R��߽q���3nv�!.������hV0��;��xѓy���hN��2(�p;�%[5�c��kn$N��Q+y��lI:��ۛ/t�pO��X�U���\崩�f�4��]��uA���7S����>�-}�dݎ#��q��р��U�u-����.�����whH���w�rQ��(�k��=O�߱��m8��ų���N�z���9UvjZ�:�ܝ��'ET�����=L�y�|��y���~m�{ڳ�tL�ۙj�����y7���B�Ԧly���u�^^:����п?mC�o�meOy7~$$Ɠ�\�쵄��㛝ӐF��ޮD�"�v��Wt�/�^-����h}� �����T����[1�}�n�vm�c2�Ns�2q���ƪA8��grpWf�r�c f3��L9,�ĭ�������%+�Z{p+���2��Zҭ;���O�U80/L�����)��,�N����~���~�E����lc����љ��K�t���|�xx{���YR�*�����O��J��Y���;eZ�/�yˊ<V�nx��vWm�Ј���j��8$�L2��!Y(�u��pn�7�b|��ZNBsh�X<���v���`:f;Q��ͺn:��Yg{k�R���_E�B���Ves�ŵc&�鍞�]Ž[(RP*C��Dy��m�B��쌢y]v�Ubv��V]ܧvV�w8��x)K�*�Z�L��@��YR�YRI�3��r̀�嗤�M�vQ���;�v.������xXh-��R�sJ�:�$��F�1��.A��ʖn���&reN�Gn}ss�iͼ��;v7��޼r�ݨb6��j�]&�9���[+�%p;��&��dI����a}@�`e0�r�}J]f�Z�Fmc�8T�j`���κ[V�e�86={k�d4݆���a�ݙ*�n�� �"��*u��x��m �Ki�Y���2�͸���&��E�6�8��䏓\V<k��-� ,�ϣ�E��a�ܾ,>I��5VwZڱt���f3a7��]�̧�l�&��Ѱ.��V�0Wv���g^��jM"��7#T��K!qX��g:'|�"E���s6�d�Է���ܚ3�}���.5Ǹ<2�%Q���dv�����C/�n�S{Ikuơ�a�}6�&me�ܩYP�p
k�f<�`rTb[{х=z1�f�0-��c�o(��Ot�h�1�Vo���.�hW;`
˳n�-�Rh�Nt��M��gl�:��ڛd�ݹ�w˕E6ӡ:S;g��	⫂]�oj��j�X�tuӳ^?}^6�C�]��M�s�щ�K�P�@D����C�
X wb� ������l|�����ʘ�
|��cd�U��f�:��t���M��qI%��C0A��O��/�&C��F׬��.�P�:3��љ���d�'nf�\��Z�D���OP����U��{%��֭D�k�1]I_S�˚K�ܤ����C���gS�FL�:��-�yx��5�	�ﱻ�pbYy��d�4ȸ���N��;�i���qT��1k<+j_���;��Q�)�D�O�el!��,�(؀�:V�����j������/F��'�1-vMSS�_KZ鷕���S5rme��ZU��p�/��IS�/�r�y�u�X��W���j��t7!����h�R2��ѹ�T�e�v�F����B��r�b�Z
)Ck(85ջ�E�H:uF�:ye��Lj���������	�EmuM�m��Og\���	
��=tN� ��c 5����"��Y>�Bm��s�GW�Z�8F�w��A��4a���ܔ���ڎ5'�f\�Um�/v���D؍X�@��{��;��8���vj���i�����+�cy�n	���v�-�[ ��9�W��s8�o���Rݬ+v�؆�����я�'�/Xy�N���v�8fo�A���h\z8۶x�7(Z]-��-˸T[�y��|�JR�͐J��B�*�߸������Y��dz���$�z9Q_0�G}S�<��s��-���rB��{v��o����
�}�~�rL�e�B&�럮%��!�wdz�J�����;م�<��/Dt]Bn}���������������=['��QL�OR꺅n'�QG$�'�v�J'+�:y=�EyШ��s�A"�T�FENw�o4�r�D:�-�L�����%wϞ�yxm\�^��z9G�Ĺ�{�է�UT�L�s�+�8��*�q�^vW�;�2(wJ�UX�������73ʖDr:��s̠��vBd^y���Ӽ�9W�N\�Ke���ȧ:q�Pr�T�H\
� 룅(�Ʌ��W)
�D��@G�t*���ۻ�V`D�w�V���t(��.�9�>���E���'ӹGaDE���Ĝ*�t�)gseE�r�C��P�;�ЍTU9�Эi*1��wP(�1e��C�""�^�U�I�2<��\��>>���{��u�R�θ�Й�z�meń�gC�6�7�)Q�1�5y��i��NKT��H������{~�ԍ�����\�i���Ⱦ�ށF��ST�x�>�wd)��S|�T.w�����͉���g�-WE�i= +��X�m��۬��^%�`��Ӈ�5N��}�+��V�4>"M ��\�p�qf���9~��4feT5n�h�T��A�C�6�!W��5unE�vxـ���%0���s⮩|8n+������W�PĦ�|����z�LCMgrf}����޴�ވ���(�~6MT�G0��+͗;6���H)�VU�<����?\�]���h���m��G1k]ɷU��nW<+�[�E�ׂhTxuC\�u;���he&,j�zﷱ�H-�V�
���l��s�;����%�}	U��P͎pM㐦Y��߲B|��fKȓ[�q*`'&�Y�ϭ������T.p��~E�%t��YV�Z��=m���K�mY!���Vc ً�h��ΐ�C�rn�@�ؠDm�U�.Oڠ�R;��A�8)�oV<u]�����u�grj�R�:|�k=a�����$�ּ;!�ʥ��E��{�)+�B��u�'W��K�)�����c�R6�%{ci��X87��I�s��[�a��X�`\6���R�gw�plC�X�չc;-f����>r�f�n=�xH���bR��ܗ}s��+�rZ�[��Z�H�2Q���k5��L�ه�{�u:sx��>��^�R[lr���]��� �����3�ޯL4i�m�l|�o��&�&a���aw9�e��׽25F�5���{i����أ��U����Ͽ]��ǿ00ڝ�>�auҮ�߉T�n(�t�Z���{�W5g�@k��F�' �<7�s
�����J�TS�C&�bӿ���N97�Ke�J��3�ؔ'�C� >c<�f��4��kb�VH�6�i�*�W�=��͠����x�w�L�1\-��ˢv�lI�M��d��dh�rj�1vG"���r>����oCg=������/���1sF�iv��7M��'��F|��У45�"�o۱:�E;slt
���nl����Y�������VI�RA���i����c1�����F`͖�����1,�b���5�AA)�z�J��Ȧ8��
j�Q&TS�= ����"�*���<!v.�iY��3��G[ժ�a��+���e�B�Q}����{T�iي	1x��T�����I��~�����(p����^�yy����Z!u��}ur�<;����lPܶ���)���ޡ�����or(H��ғEN�le01�"�V�m�W9Y��j��
1����;+i���n�
��.珚[�2E��ԣW�.��g׀^�2�D>�W5�6�� �h�ioG��6s�ύWQ�i�"x`���,֢����P���5Źw�Yz�����Km��ZcJ!�	�=>m�>��"m�2�b�2z����{������{I���]׷}��/�6�yA\q�}{�q�4��T><ː˫�$�p�f�w(\v���5�KŐoV���C�����y'�c���W����4�}1^��-�<F3�eς\��zǔ�Kx���Jc{��Tc��j4�RU)�t�	���<�A(VZ|��98p���\F�b��u�_�_��E�.���l�A<�����U�p�Aij�S���G�z44zӊ �-`J��WJr`��{ɚΑ���qH	��-Bfs~��@��b�ĪR�qG�<ԟt��Q|o�[�+i��^<'�!���Zk�᳈W��'v�qN �n��}.hTS)��-�$����^�<�dP66b�]
ɜMч"�4�/!�!��,0ώ�1��4y��
��D�:[eN�n~���zd��g0�:�swߘ���ρ��^��PC��ʀ�H�.�t3�d_h!Lh.v��f���D%I~����9�=�,����j���kh|`h�H��i�7gfk?W�#�ei\&������'Yx��dkh�dWJޏ_oiYd!�u7����rG��zڊM�;Y�θ�ؓOL��(�i��u|4����e����;Q���L5uI�@�L���ag�����eÔ��g�����<�����#�i����Zb��ɮ�\�n�"t�s�a��C[Cr�!�EG\�(���A�>	(�u&U��zV�"v����nݍe��-��z�P�m"�'+ئ�c]RCdIa��=�Ih��O&/a��4$�£W.���.��v3�*����Bh� ��UЬs�9F_J�qpj�q���q�I�\�0�e��?�4h���:�T�M��U�b	T�����z�fB��y�ߧWk��F���e
WP\Ȣqg7f	�����v�4�x+��6�Z.���L���q�'�v�aFX!}2[���2.p�m��WX{�v�U�T���|�.a���aݝ�&Ƽ��뼳ÝXmÒz9Q/~s�0*a6��m��N�X�7�XSE������n�w,����ۓ5������7d&�a�>��j\X4���(�O�`.�9��R���T�ݎ(���'Y�Ǵ�颓��gwG�k�;C"Yv)������YU��(�]
$v2ʠ�e0iU��s"����y��0Ƨ�{���j;�\ǻ���ϙ�\�̙�e�ڇ(��%��9ۙp_�
<iEse�k/�VЩ���d�{:�»1��p�Us���)�Vm[R&�t����,nU��8��.�/��{���ꪺw�IY+ݙ=���L�a%U���k�T��M%�oJ�ƺ��\,[bQ�i;aO3�))]�����:9i��?9Я�`���`3`�c����0�	����(KA��3f�;�ZɃQH=�i�ʞ��%�i��iO��	�������s�:�zzX�uf`��ǺʹN��&�Kv߈m���LeѪ����P=T���ߝ��z!g���F�/���e����0Y�a��g/����5��(I�r]��ω�����aw(ȶ�S5}Ƙ��Ȃcd�y�hy|��z�v���N�	��!0Z�{ \v���O09N�u��-��摂|��p��q��`��h�k��)��8W&���E�G:Fb^�]\{E�\��r/��Ba�����	����=-��Ge�Q!3r�b��n=9u-������z~OBj=�^��~�z���Wc�Bf!ee�4ki��]r��y�=i���A5��ݘc�<�m��i��S��peTE���w{��L�����ӦO�?zJr�de7,�M�1ˋ�,���m�_T��.W��gfx����S&�$�m͡A<e��o6�͝�0>(� �pe�ڬ�7�¤��!h�v�!�d�X�+�RG����L��5�3l-���fY���%J#ZN�8y8���.÷7�s���U�J=��;��q7���+Zf�,��꯿�+&��m��T;�����Gh�L����+J��,��r�U���2�9��ٲ�T
T$h�#y�����ͷ�y��hO��x��o���ha���cХa�e�[-Y*������N����%U蝌��)�3k����_�M@���v�䨳�!DR}ݝ�)�CM�k��@~�.�{nG!&������;�n�.�Ϡ�E��Zb|�/T@f|��h��nD��|]�^�v�A�ݹ��D��lLwu�Ú^�A��L�:;�醍4���%����b�M=3�[/"�K�V�SBr�Y�B�<s�d����}��O�a��3�T�|�Gx_	5O��eŧ�H�%R�}
2�ke�n�W�,K6��1̬�P1T�Zv���5On^���Z�r��8Z���9�2;|\Χ���#A����zJ03�k��J/�Sf��,���A����P����Є��ӑ�3��7�K�dq�ӽ{��j�6�{��]���
8��T�tΘ'��`;>��bC�+��ͬx�W�g	�2 F�cnv�����Χ�/�sn�v�j�����^�֎&5S�� �XԻt@�]z�T���F��n��0�1�U��wY�J8fkNn��Y�8���0Yv�
�¹�IO�־�X�`�ecWf�;ݽ���GQ�s�5S�2���ki���3y��o�r6�4��5tl�e���6oL�%�0��C�i~Z(ك�(��O�+�V:��&��;����.���[B�.�G*�3j�r�C?�'!���j�E�"��d�6	�{�J� ��1N)�{N���3�� �t9N�b0!��Sn��*���]�y7����]�WXwaﮜ�B#:�e�F���S¥c���2��QEՂ��r��l4�kW��K�D5bq�$?�CNf�6J#)���v����2�#�s�b:%65�	�=�QI�mȬ�rj�b�c�={�$l����pC*�#�C���P��-C��ʵDq�w�z���O�3zSJ�9��m/l��n����v��>��	|� �|xbv��C@�2�7�<�*ڂU�24�7(�̮s�<S.~�Ҡ_�֬�l	Sy1^/�!�����}����A��ST��	B�T֪��U]��<��L,�&(�y���/�uE�ӝ 1�cf�qB2�;�����#���C�ǝc�p'��P�dÉ�p�aԌ�D�sD@6+��H9��k�4E�w�]�i�,�K��-[��/����l,�q�|��V����/p:�k�@J�kB��b$x�k�LTZd~���{��r�V�n(W���7�w�H�Z��,�;>U�X��R�3C4qK�̤�dfn�X�bЛ{����o�2蕚b��nv������f����z����a�_LB~h�%֊�t_g�H
d��<e�>�k����,�\�A�p@��vٺ����86
�����9��2�1���S)9�[�L{S�*9�:Q|5�(s�K�B���F�p2�:dh�6��tg9�ѐ�N�b�Pkv8+e�l�8A�T��Y�=Y"T�	�����(?eR��z!{ρ����u딬y��@o�K���g�Ⱦ3!��ۜ́�^J�y�E�'�kL�U�C�1��ag��3��=@r��$=-��Zۡ��F���WM!T�;����k�̃��~D��d��ܞC
mQAі�s�V`�cl]�z�[:P͎f������Q�^Qj��cZ���R��}	�0�
~a���.qM��� �QA_DNv��s=C&�r+'��A�OF�b;�按pZ�@�c�L���#��O�m�s��C]8��M��Ds0�ەm~�nS٪_qd�_���s:�^�O\��wJ�m"��Z4��g7R����רq��F��P��+�j��%�%i�o@��e�^`
gɸ7,�"���*Q�rP��%��r/�n��z�;Y�ޚ"N���.W��&U���x����KӼ֚* ��Y�`[�+S���sku����,��(�Ԉ�E�F^��M��٭�υ�Jv������z&,��8��>��ggS��_���9EA�. �Ϸ����?���_�ۢ:c9��Ħ��e�US"��X�c.q����y�+�#t�h�"���*�.�G��=�,q�� Ӈ�;�ϡ�%8	���LN�M6O�����m��KE�==�fa&A˦s�6�^�� #r]��U�	M��6���7�C��.(���N�"��h�h��Q��Z�7FN���s�3vy��LS����w~8&:_�dK.�U-�NЊ%W'�(�_�����l% �|,6o�wF�:���O@�>n#Hq���i�t��bJ��2�#qQkc�L�gyB�p���r����^�	��b�-�L;n��灬�wa�����B�r�0[���|ΚVwKOF��K�RNw���j��R5Z�Z���71�Dh��ym�F2�=o��@��k��xW��Jl3�rW�)㓼���yQ�^i�����꺈����b�H:m;=D�Ǫ��E������ ��ls���05�{
 ��20h�N*�؈3���⫽ Һ�V�o5�"�1p1�c�q�p���O6@^��Q"��;������F�t���V�wf�Kة���F���.G2��7�n��]:����}��$�P-��l�Y����=%$M��{Ҡ�p�5�뀬i�sLw��,���e��/��ȴ��V���w����e��V����#f4�.fuZ�DN�Y�+����C�v]�L�G
l�7�??>ߟ���~���F����ϳ&·#�..<qq���m��>��Y�1��/t(���X��m^��`hCz]�i��A7N�D�{8m�A���4K�g-�wB�E�g��B���5q:�0�t�c�&82�D��W$43Z�E�<�L���\�;j�V#$S,Ñ����*�3]���Z��{�CK:�BrbM���1i�ŕy+�^�E��]���."�׏Ti�',�Gk�f:�s��)�3�I"��W�ad<p(���>.3i��-�䢴�y�N�R�mk]���|��v赣q0O$Ж��#%����ڝ^)�c
Q~*-98��엇7
�����XI����6��zs�}R��hg���#�.9�73�Yڀ�J�X�r��<7!�Isvg:�v6��c��^�#As�W#u�U�8�͆6E��h.��a�=E��Z`���W�UȢ��c7���Uj�����={onhV�mM�Ia��K��0_t�Gys��mt�ma�좰>J�����&�=�jBr�:��@��ܶ�H�����f�x�Z�}���w���(eo��J[ø�T�m��7���� �<���Y�)���z�D��̥l̓&�r��vv4������S2R1�H뺹�ڮ�jv<��+�N����vi���4�ݭt�$y��Qp�������krt�H]���f80;q5��&颫f��L�ԛ	ך�$R�SZI�m�{H�}!ş2��Q��E�]q�T�G��X��A�7M,�����!�
���\�ۼL���!�ѐ��N�vݜa��e)��]�=�*�r�Ma@�
�9�)� /;(C��mn�Mr�*�!�I�mO��l���#w-Y�;���%����X�T��V��0�ub	�s�gI��4�Z��hѮ�y;ɫV��)+Q��Y��F}��]Ѿ���P�i��x�з��c�o3{����+��H�T�Bư�N���F�]���!W2�mƈ�i-�$��r7hU��m���8��ͫJ����֬� �X+�������6���.�j��Z�9������󚛭b���v�<�3#W�'z\Ry�ሪ�o�n(O	�u)����n��2�C}z���2�gy5��ׇ��0�+�t-?_f.T*)iV��v:�id,<�:]��N�_�ncy�F���+��u &�(�חٴ����������uo%k�ݭokV�3�� �ҲAJ06S�NX�>�n�4����w=u2#�I$��R���x=���7�[Y�5[�uZ��\�S+�E��X��Ѡ��$�&�����2���u;�wޠ.,RK�gɗ1BcȚ3�K����S@^��4�&͑n�
Ҍ��Mb��c���u���D�v[TAYȺW�8��.�5f!��7u�iѣ��3�[�kD�`e�-��Y��ܞ驎ڰ4���N�M��O�*�n��jn�J
!0��V�ֺr�ʓ�޲89��V���2�X�V�V��k�"-<,�˒�)�K&��QLnl���+i��:S��q���lʖ8b����&��:�n�gFfN��]ڶ�,]Բk�)zP���Tӵ�P ��9PU����뾶�SΤ�e����%�`�.'�2�:���ʁ�Ә�]t���v^��N��&���/p�uM$F�jY�S�υ�@m��X.bU)@�P�6�Sj��Fc��u��t�W	r*t��c�م�D>ƹ�H��c4d�f�.��J����c-Bu�S�
Jts����O������,�'h>\3���缕d�M�zu�
���-^�v����Y]��q��3;��md�SgُXx���	/eGz��6Gm>ue$쬋�ei���2���n-��i�͆�X��Q�Q^��]��<��
��镻��K�QH��R�upT���!�9���g�ԫX��G\ѧ�����SR��:ȖC�9�=͓�ۆ��E��1�ĵ��F�0J�F�{G+ �B �-�`�l[�_z�����	�v7�j�4��{�2#��y�_oV[�1"�e4��"��z�$k�Ѿ;�~+8�M:q�̒�Kg(�.Qe�ȴwlB0�*���
v�o���o���/���e�Q�YI˕s�>76K&W����G��]�I_��Qݾ���|�㲯�ڴ��8T�'�Q<ȋqn2+����[�>���\#�:GVһ֜�&�Z�Hwq����i���NTT�Z�q�)�C�D��w{�
vEB�N����(�"���o
�]�>��ۄ�����=Ԩ�������B\����^���^p�n}��ϒWt�>`T�G֞*���^�I8}�r��UA����Ra=~�<�S.�q��'� �d�"��HN�$D_��l�p��龻��.>�q�,*�\�x��G.z�yDQ�NU�9s��氾_@s�<;��ٞ�QϏ�>����Pŗ������>�q�ʵS\�g�
�-�O��f�Sׯ{��S���gϝʊ+�Q)�\$�t&��t����TJ��?���}}�}��H����3��W �u$@��r�W-��!�+�/VK�F�}\��.,�nM�+&i�Ņ[R	�s&���EU_�~����Ɍ�9\� .aw����~?/OIᑩ�Kν���z/ �B�U �V�AF}K#ƥ��tK5�˃4�?-01D�ח�u�gXS�0��Z\1X������3���H��61Цx�|%ز�T�C��x�!��6���۸���m��
��o���#�|`����x�w'!�MZ."˺9cS�^.�Y1�h(�rs��.�;�ϏZ_��N˸�^��FcB�m
�r�۹4��L����S�P���(�|Y;���z^!�I�~Z)U(����z��q�F����H�n�&�\O�u������0���r� ƨ�*u�1<9�0ƺ�竑;Q/���-��Fq�ӡ9�ca��L�5_B��R���	g�I�b�r�:\ǭ�r�4�n*�h���N�h���m^��2��8�u/�f��5ZP��_:`��'�sUCFj�=��)]�����g,�C�[.G\�{��C�LϹٹy n�����c�h�ս�#KvP�Nno)<�WO��y����"��G����"Ĵ@�Q�)N_�����û�������iE����!��`�4�y.g��0i�,ZX=�
��G[�e�=��f�U:�MV]9>��z`3N#|�λ��`x����yE=��s0yef-�|�tvi"�9C��p��Hu�7n�� ێFF���{��o3Ɨ]�t��^�l-�������T�r쉑�A2�����~����c�2�/��ȕ�*�m^P�rr�Ķ�d�* �!?P�b�{�����EԴj&��1d.Ti�����)��r�b��lƎ��y��Db�����-sU'�)j��Ӱ��Hl�@k�y��?a�Ì�n.�T�]�Fh�_�+q0�YɆ6�˕�(�����t���pi��u�<���Eh�'�P�j���Q���F��N(�]kzL���&�/��dK@�Brx�h��:�/��B�ĪR�7`ߍ:{��}�:���c��5��Z�sn�*`��ָ(ΐ�T���4:��&cS�ۛeB:L���U��;`f�e�7����a����#�S�~3�0ނ�0��c�43��[-Q!"���$�0�sn�hO���*ؾ��	�kz�3㙘,^�C���^EOz_���D����5��4v�e��0w����`~cۦ����k�.��Ϸ��Qq�V�k�8x�eӾ�d��A���繰���n��I��}q���;��r�9L��`�T��r��7�Wt�kj�Y����c�N#�R4)Ջ���Q9�׺�-Oa�I�����Oo,!5���쮠4�ڮ̬w��<n$��g��T�ֵ�F%˺�k����Ml>�{.Pf�WSY���l����b�iM���wZo��Q�YI	���ve�J�*��y��7�f�f o3x��YV���ߎ�a(;b�_�uxw�m��'T����t�0����%���;$;�B8{�tS�I�X��$46C�y,^�+�	{~��E6R��\5L�i���"�����H��U���~�3�v֢�Qԣ�N|���a�ꑧ�e�W����ګa8���d$�r�`��`y5u���*�i�e�%�Q�V�&�!Y��țl�<�M��r-�[�5���*�R�2��I���S-���m��j�1Qqp1�1Lkk$E)6
6���&Gn^��^�: ��B9R/nbS������Ԫ�տYَ���?T��U�8/)�xԎ��;�9�v�BH��@d2��n��-G�O#l���O�2��O����n6t�D��~d%@�g����*#�4�;E�m(q��_s�<�?�rsYvD�Fn�僜j��d���zL���[cH+Kt��ghwPs]��,&FSM��4�V�<(j�y5�Ԭk����N��ϒ}��C��M0Fрͽ>x��!��9�m����MN��'fFN���̜�u2�-�P�=(f^tR�2rF�.�$��4]�����#s��`f�W���䴺�R6����JQHm��)���Y"�j�P��[��
��\R�n��h[���I��E/��1aW��Y�V�І�R
����������~�L�6D������A�1o�#��k%*���%��֫��$��W�v4a�s�@ր��4!\�e�PP����3p������]�U���`�/���y���G�(�b0�S�K��N˵�1�n���`�Y�S�.aсR��;c�G�t��F��Dj&�t5�(�D���n�H:RJ�qK�v6D� Rf�8����ᯔn�3i��A�q�v��h�Ұ���f=miM�qʙ}	��QVX����:`� !P�l,�~�w��C˩g�]$�ll�bwD[n�ڪ���Z�ޢ2P}�rF�hp�%�����W&Έ',�p۴�GQ���m�W^$�鰟�n���
Crg[�^�!ԣ�G��
�W$5�.�^�$�.͞P�,� n�9te_��R�mF&楶�]N
�t�	���IeP��e��f�[�E����Yq��Ʈ.hA�H�]��à�]bj�<z�1I�:��B�ؔU�9a1������"�L�����#?��ui�;?<�BZ�2m���}5:��ǡOa�$�u-"�ܡh��P���.(=̥��Gŏ�����*�^4�O�Qp��:mG����N=�z�͚���h�Vz;�I2i�U�:���m�`��֧57��,=����§T2���8h�\w;�,L�O�b���wPe���J���3U(����&�L�&80M�6�Ͽ���ߗ��J�#� �[�8ܾ9���g���z�}�̎�(שL"9:�W	3D���;�9�(�.�������^�Hw�*�a,5������>���A�h�VQvH;>�4�C�?@���J��rK�	�ܺ,tƶPH�bb�&�)�?�W��[�+��߱v\����j��
�)�ۚh[X`�׬ܦtys�W����<s�{$��w��j�^V��u�v��y����4�g^c�л �I�߱O3����1:��a�^���I�#�ջw�*q�Yt� 8��y��h`Kh�c�y<hu��i�ƅ��ciN��]ֻ��>�m:o'_4>���ܞ�2�Cān�@�yݩ��c����V����7�{{����2^�ֽ���eߺ5�"n�5u�H���h�]*ZQ�ߝ �r�C�Dg���{���=����t�ؠ*s������I��-�)t-�=���N��*��sΓ��裶���P˴<����Y��k����p��ܝg���ITS�;��S�'ŗ��~ۮ����4���$�mk���߭�gw������
|�!��ٻȳ��u��ިwQ���r������ے�7lN�y-�u����$��nG��N)A��*�"���񇾿w����w~?L�dCa`�����uqz��"����K�8����X�UP�,�a�%6�FD�V��w�r�r��q�ۛGu��93u��J2yD{�v�UDZ�b���U��xV%+^�A�=Z�O�%e�Ԫ.�q�;rِ�H����ܑ��5�ڮ�{r��D�X.���h��&���171�h>�B;�	�����)��pd]L�s���e2W-Y^m�'���#��;gP��qlY�mV�jF��\y@���H��̃��ϥG�q[b��XL/(m�r����ZD1��hd��1���qݗm�A����-�s���r��#yI.�!'E�����{!�uSe4tS���Pl�؅�o�� ـ�cxMf��XZ��t%�e�CS�ay#��aC�Jb���˳��%(VZY��rM�;+'v���h�3qG�r3�F��Sn���,m��1�	�y��؞�2⅛U�,d�8�0x�q��D�xgn�O���tbAE�3��`LF�5	�I��{�gJ�.׭}�QuQ��D�W:���|���w��ZW(�->�k��}�0ނ���`�>i�D>#�/!G�6xx���PIz�"�/ߟ��?M�׾���%��d��+!)��=�	ڴ�sa�l�vޝʎ���R����.9`s��,����⮘N^�pO���������qXe�ٶ3�9��CVZN�e��b��< �vi�ڔ�l����nf���Jf=j�N��+tDB�~�?W�C�_UP�{��� x0` �{�c+RI;vN�!���>E��z�5M�@q�h/@`�d�4�=�E�5~�TtN�Xe/�4oT����⻴t��E���k1Ȧq����t[���<���]��1�#�����hF5�����Pzp�x2�1�ї��uݻ���|�oC`�S6'��ʝ�g�:��J{�Ķ�F��i}�l^��a�.-17	��4,"ow#�<l�C�	��Z=�(0��0���Ix%
��e�d�h�@��ꈖ�9	�z�S��V�;bd�tX�|=gߏ�*;ޫ�]��]^���ܷ�t�q4S��V}2ȵ%�[FED��2�.�*}Q4�S"��=��K�1�걍�:�C���
��=3���n3eWN  p�ߔV�3^Nܞi8J��!1/i�i��"���Sb�����x)E_r�����3Q�V�.͓!Y�K�'�O1ώ�F�Ok���L��2`�W�[k�]�wD ��@\��)�Z��
�Ʌ汚�t}�ڋ��
g�FW��Z+�.Y���l���co�W<��^�0��Q"�>������x3���0���H��{/V�1��~��m���W\Sn�'��%��\M+W��x�~���H�=�{|���6��S��O��m��Aܗ��	�JSw(��)q���u�o�ӛ/`.�8���tum��57 �dj FR
��O��o��7���}�  �o{�{��R��l��{j�e�\[T�E�ƙv֡Ä��4_��;8ڗT�(�O͘��Ɂσ�b��;��f�Qн�y�v����J8+�z_��c#���z��#�(f��˔���%M�����R脊X]�ͣ`���$�Z�iP?�׭�K��i֖�Lg<J�a�����R,f�^��e<��ѫ�C����d���0�c�Y�36�yT�K��Z_$&8ׯ����C;m�y��'�j���L3-���)��l���; T��
3�M���|�c�!�K���Ƴ:Z�u��s�9���`7U=Ύy���F�r�	��=�����w�2my�Yt4�V����{�dY��R�<z02/�#S�x�CE]�E8f����]�=*8����[C��@/��@Vx8i��������<�l��;���2}�En_<��+m6�]��u�f~�(Θ' [
���(Bb^�U5ǣL�et5'Uv�Cf�r�ݵ�����v�J�L�kڬK�t�F=�I�>;�Nf��j:��C�����;*�.���(��mI����I��t�IX1�S��?Z�L�s&������Zꛦ��nj��F�
���t#2�pyڱ[J�C
��%t&��kk�k-��J����(%5W.$ؘ�K��=
��:�𽨭t����:�/�r����ğ���7������=Y%Q3���%�/v7�ְ�TרYR��T�mr�%�1\��֞��L�\e�����}ms/I�N=��'h��BЌ�Lr`iy��	�����R.��W22��N
�b�r�g�z�:�N���WcPi�^w������y�߭ݲ}p@�]@؎�:�	�N��tRsh�m����1�T�gn����r��7���>��y&��9A-��->�������a;Unm�a�̇yxY;�-�^�(yK�_�����g~�mhV_!<B9mv4{�pC����	f����̃��_��OݡH:�e�&�C*�/��5��xE�b�&:�����۰.��\��#]@����]�c6]q\��q=k�YK����i�;u�w�؝L������3��^���H����"����곔���1�b|�����{$�4�Г�s}�nE�mkNV��cƞ�C=��0a�I�w�I:�0���6'�Z���q��F�2�ح����V�7������E�M�4T e�����|��2���6��b-�41�����B��oZ�"�΢;���f:J<u�դ+Rx/���S�J냴2�jJ�vr���e���y�\�c��(v�ח_���w�M���,�j�X���*�ɨc�B9r;�`)'������^[�c��gP�5S��m��3�o�������y��/nq��3���s^�g�a� .<i�9�6����ɷ��{7U�4�Ǧ�#��
A��^�+��2����D��,�<mDZ,�4:(98���! �m.�OH��y�#6��0&:�	�t�=�} nz۞3���-�)t,��(Θ':K3�a�7��o��.we��b�������`�a5��X"��K=�8������@a\��_�\�a�Mê�6�B!��0��'������]"�T�z��qM^�[A,Ի͘A�=���`C^Sn�2�6ģ���C���~H���֌;i}󫴧���V�4���*ͷÜǥ<�S��Dm�
�m�6շ}�0�:H�C�c
j���vUs�=΅��@��ǭ�߯ߊy��?� �O~�}�v�9�+v�2/xyˢ��S�_(�-%e�BGbCϝB1��g���.ʌh"j�ks���ؾb���5S)9§ț���V�(m��sc	hnᡟ�.���L?\�4bߤ�l�:B�h3W����$���1�9��>
���F�f���}��v��r����u0v7�o	�WHR84/5�{�����T�tS�\S@�4^�է)\֎�렵N�X��p�ዉ���KՐ�窮����T2��5�;}�h��ȑ�e��f,N�_�g\X�[6N�2)1']�q�W�p2�b��е��ގˬ�X�v.�%%�q,����ڼ��q����[�؆j�[V�e������.�J'a3I�����vg�si���Ox�ո7a�7���O�*�w@��-����L���n�be	tZ�؉��������X�dU�w�9nb V8��:&��Xo�������P'�-�WK-��4	)ӣK�N�T��w��Vgmo"�o�k�*�{�:724��`RR���\�.t�WZ�2��].;D��Z�l'��.�w�ϫ�IfE�3��s�!��s78�S��cz�]�àF(�;�w�A�,h�
��f�#��p�\��-ڣ	n��庲��-�h�A_T6��g,«o$�l�ź��B7�1�.mje�ɜu5tފ-���r���kg�EH�_.�b�b�%�n���'MTyBu���1�j�R�is��fb���V8j�y�]Gy�R՛R܏�o|��z�<�Ɇ�r��׏EB���A`T
j�O�j,����Ms[M��{�ms_�K��l�w�,�V��h���5chV���~�|�5a��x8jӳ�
���\He�f5N�$ӫ0�e�p��L+��c}��ie5R!�r�-��\;�c����t�fg��Ad��P	�K��B��|�5qN�v�ꊎ�d�����7T�e':���7D����nq�}t�
lJs�Y���o��:7{Φ�.�	�qCǦ�"�9z�S��H�F%�UnPy�ʈ���r��0��,�w#3��r����V�P�Uz;h�\䧼{�Ԏ�٣�%jF%�(u�y�x�mꏖ��g6�v�E͈ů�T�Nu}�+h�oڄ�d�����&i2K�0��h!ڒ�Cz��Wk���{SnWssY�{������;NI��.!�z1]u{�2:�0�ٗ*��;d(-��4��Ȑz�9^�Ӥ�{�WSJ�����r��PϺ���q�l��J6JH!�ǻ��gN�{Ӎ�Bv��rY����2�R�1�&d/SWK�ۻM���Ц�Jr;��k�_.M�J�S����ĭ��[
�cQ#��S��7[�Z&I�����/6C�r��]��ܕG �2��iJt*��w�ҿ�hxE<�ǡI�.��7H����$��L}&Ψ��p�N�I��Ѣä���+Z�ҽ��Rc�j�
��u@�������fm;�:��6ST��di�u>��?2\�rtw�y�똄î�%���t��l�Sm_By���.�T�9��}��S*�z�xA����Q��\�U_�,�I]��q���(�ȯ��u^I��㷷��}o��I�\(9��G�9�X���9AUrη
�=}�}V'�q�!�N����7���g�~*����Q��#��h�q/�<\���ʲO>�U���	4����w!�珞�RM��Q3��qv䐫p��W>~�8�I�9�w=ݗ(�__^��Iz�N��E_�a�?V���ӛݸ�/w�U��Q¹�S�v��DEy�3�
���3�S΄�^�rB��M�ò3QGד��
�c��E��<�: B.��y��E]W'u�J�OS�9EW�V��I�乷�p�C�&�9)�s�w�ʣ��U99�⢮��7�ǅ�N�NWR����w�!"�d$'B#�E��!��(.����� ��#��I�� �@��Y�Eӹ;�ϊS�F��L��K��*��d���}�h����(om�)��+t��%
Y2]��U���"������ x��K#s�Zw�帊������߃��u��C�d�8�7�)Sړ�]�qH�L7�Ŭ�;|]�{Z�&��=�)�`�m�T�p�LnC��M�֮���V��<��N
��7�ٍ;h�E�OI�
n����f�<�y{f�2�&�����2hN,'9�b�e��σ��N�������b�J\l��ў�y�z֜F��k�??:��*p��j��L�C��v�vC �)�L�>#����m�md�L.[-$>���h�R�^���/�t�3I���%�����oap����x�	����ٌ�Db���~��{&���<k��`������5��g�38�;���_��X�s�t�+�";E&u�Vfち����8'������,�8��b�S`.Zgg0�&��
�viv������v�*18{��sώ0�z�9��H�5��d��ݼQ��so��V���FzU0e�m��GO?�����¥#���3އ*����T��/`��T��w�*wC�����I#�-hjF��ӕ�V�A7N�GK�|��y繎�-�2�$w<�,�`+��oo�;Op5MbT=�V�y��f�iחU����MV�CEL��	CL�V�ԩi�	wz�^Lպֆdʓ�ګ�:,VgֹMy�&�����y�-����������=F�D�?Oq�w�{`��|l���1]��������o7���3x  ��Ȅ;���<��uj�)��2جCL�˒���b	� ��Ĥk��Π��'�MYS߇N��C���{�m�P����i�^*���WtԲ��j6J�,�ݜjAI�踪{��U���C(�h+I�v�;p�_�Kg��&�2���8M������2`lJDN�h�T7dgO!۩��y߅�r.�ۂ�-���/��F�RkͦL(R�����X2�w.i�з�A�yՒuB�x�	��!�z����vM|Z��4���TS��`�x�Tʙ��.�sn�t��=Xd/b�Ci���>���U�<�%�+�:I~;d>CO^&<�U�{Va4H1/X�]�d�2#�{P����L����d�ۆ}��<4�0��x�3��D&�k��7iFn�u��1����T�^�Z��S,m@�PS�u�* ��B��h�fސ�43w@s��N�
w�6C�A�|����G	|ؑ;���::nZ�3I38�Z�ۈ0��������V��_5�j�N�Ϫ\q~2޳(�l6�ؔr���`ϫ��Cǒ��^�?Dߏ����c9��:��$;��3;���ct;tδ�^�Y�O;�kD���\��mn�4OP�b�QX��v�t4�*��F��vZ�>��I���Ԯ��Q��&��9�o`m4�'-a��,՛K�)}ΑSn�R��S�D�A���HTJ��T��������m��٫�<��~x >�{�����<0���ܜ�K��a4=��l}wf�\�v�0:B�/X�d�V�28(4��&i>�ș�Yb\]�m�񛪝~���]Q�(OR#:���� ��-^�TW���v�ưT�6�I�!���v���!�$su���(���A�tgL�<K��kK�h������^~Iɬ~�{{���9q��	�DH����Tד��n�;�M�.ц�@���Z�,%�O�x!\�8�j<n�;^�Y�f�B�2|�#%�\�����%�Mo�Ā4�vW�j�o;�`�&�K^�r\�Q�L]HI沮��蕮F��iD�l�8�Sm�����2\�kҙ����!6{�`���$P���Ɋ�4�r2�;��e9{@�tI�����آ�8�)Ol_XZ�1Q���6��sW�X�W���J;x<���x�`Kߑ�/��v)����]�B��wbU`��SV�������%���ӓL5��ɇ:��@�X��?�|���Qp��Oe�b����~���x��N�"����H:����%]cC_�d�ヌs߽��?:�h�������C��i���[�>�͙��<�$.M��RY{�_�7����[yn�m;�ʆװ�+=&yh�=�V��ЗM� g�-뷜qP7F�{Q�Y�u���8`��ѕ���o"2�⎿�UU}��W�C���{����{���iQg���c�]�7p`�m��;���_ڵ�a�Z]R�尒��X$K՝[��)h�hM�4''}R'�{�j�a�/f�4'�Q�-��Ԙ�6�@쉃�w�9B��Oq��J�";�c����J�2gLy�:Z��J��A�*��}�̷ppz-�2�F<(�P>�c�Q0C���
�N+�|ۼ�xr���"5&�9"�0�UW�oZF��h�2���-Hy���H�Β!�Y�kZP/	�md#�fn�ڎj	?R�������<ZN�A���á�6�y�h6/��Ǽ\��d�
�[K*Yy 8ՙn��sMq9��"�C7*�'Ǟ�GC��=���zG���%<d���5�13������0�˷�!�-�ڏgp{=ʤ��)���í|ʚΪ�����1�<s!����z��*�Cq�S.sJ`�ǒ~`�#"[4˞'���m���V{��:T���8���ö��P����%=d�]���a^��{aP��bj�����ju�a��,���� �:���k}����Y
P��c��S�_�m� ��B�u�T.Ѭ��օ�����(,��L�R[��Ź�:��۰ٗ	�&� ��+�k�}2�J,v�q�p�;r�� W$w#R����wt(.v�e���x >�0oxx7�x�M��J%pg��y��$v��a���C���T"1��>�/�ς���L�r��W�G�SP���E��_�mׯ/a�Ow�B�ʬ�~�m�
���C�z��N5'�-��-�''{bUem�:���˧Y5A�E���/��N/�,������%�p�5�%�A���g�9��0�RO*
`�s%�mΆ��\�m�H�Ys���>�v6�����[U1jX@zx�6�:��c�D�L]�C9��A��CS���<��i0�0��#�*S.�tO6���8z����E*��1�q��A�b�&����6a��6cLnby���Y�\���������3r�kq��V6�4z���x��#�>�ii�t�������vw�E��K�O�u��xh���pv�q�L�:��8��Q|Z[\��q��mi� �4�\��:�~S��6B�ۅ%��H��j~�~���7虁�w����oav[�ؘ�J����Ϡ5E��d���L���J}Q#��F�Q��p��'��F�{r��׮R��ڨ��5�ˇ�Si�fD�_䐶���8s�h��<jخԔ���)�!j�:Sꓬ�{oX��I���P������?P�=�$�_���C��1C=O�v��)�5S' ��c�,X7pκ�'�f�;I���&�gkq��M��Ke�"c#� <>� <�`=���6]^���#z����?C�G��G����2�� e�/��� T�	���
��0+���˖�(9�� ��w�;Q^�Ů&㑯aY��ur�֞D�'t��Gsd�m=�H��o1�a��@���[6�������>��I�ʭڞ�>Ã�u�C5��|���(#Ss�"��Q����M��4{���N��3�S�~0Z��g�[D�T�xfYʐڟN���.�U1AT�׉	M�&��WB��T{�-����"������ͷ���g���H׾jpeS������QC�@Gk֢Q�OC׌ܮ骼�$��6N"z,ʂ"y�]E�p<�;�,z�%�+� �����D�	�L�
�d\�E�cu�]Xc*�\wU����B�����Jy�e�n_[�l���nC@8M��+�����a֔�^ .p2�e�n���=ϴy4tS�ŨDz��`�OM�2hŤ<�E�CX��O�Q�2��v��c��);�:+9�d�%
γ
���v�`}��84;��:�uF�~�^���X��ک�ʚ�䃩�:y�e]�d�AI[̀�"#$!e�ሡ6v�7���ȳDK���Ѝ�x�
4)�_B��8u,���s(rQ u���3�M�t���_M6����}��hq��<�
��H�b�o����Џ:��tB]ɬ�pe�vk�|�;����y�=�����w��K�:[��-���QB(k��r]q��aBӜp��[ZX��Z�jd�HX3��D>�X�M�yT۫.��a����\�?#�U�(~����^���.��猛���/p��@5F'�/)�P��֑�V�;��~��ȵ^f� ��6x,#��#�d��[�Ξlq±�0��ݤ?��f�	狁���F�e�C��2W�����:��Jy'��߻p��/oK�8�Ty�0����r���_q��G��Qs#Y4��_�<;�ܕ*�s�O���ƟlD�e�X�E�p-�~"�|�3����z�M�����mË����o'B7(��!���E"�|�2Q���\X�\��%AO�&�!��1��F{�=�]/NO�D]̸���C�(L2Yt�!�P�+�
7�I�>jy��6�h�Il�d)����s��ța�U]�S�^��Q"�خHh���w$M���v�.�=���Y�Z�gJ��T5W�$S�R
zɩ��c�0�&�-D�3�DW-���E!4�x�U����Qӄ_�u����"����Fdn�r1�C7x�j�Y����tn�p7�Lfա��Gt}�}���dv�1�զkȸY����(���{XZ�;j৯S��m��]�'Po�͏bz�^�E�{� /0���� ������5�=�1ˈj,;^<�Ш
��|�H�d�M��Y��V��*��n�]���;���3����U��F9��s%��ȶhJ ɷ�����CTƧ�[\��ےO8n�;���NN.�{ji���� �{,3�SO��a������Ě�.��s�N��V�W)pD6^�T
�*���*Gk��e�S�@����ި\R��ݩ�W7��Ts�hd�Yp�uN���ڝ�oT�+:�=�^��pT2]t���I'6o���/.s쉦��E�Z���iއ�ӛ���Wc󘞨Aѯj��۞=\��l4���`��K��b�90��d��� �����3<����߳��]Ja��g;�>)�n�ŹR�33�~��Tm���?5�@g8�}z�	�kpH�Al�{�O7ף��ZF��ޮ�~ڥ%�%�Z�U��:�#M����-�0�  �#��p�b����)Mb�X��v򹎺�B�lj{3�C��e=C{��Ff���H��:�f��R'�
"um'����mh�����$�g�Tdy�T#�b��.Jv(�]�0N6 ��J���vq^S��Y����;������wTb/n��Yk�c�xfI�X�Cƺ�Z�Nm乻:u!!bC׹x�i��띉��[�Z0it��2��%��  >�x��oxxx�w�����c)��Ԩ蟞 0y}^�*���z^x�]�Daʡ	<�
2�`����'��焕l���7�wE&2Q��x�1sC��[F��������.`F�WD]��ȩ-N��e��3�Ow���rW5h�N*��)<6�e�7h�UC՘A��
�E��d��Z�O����BĦ�(�L7lS���ʖ؏\0�3�{W.��ȫ��r���i�B��5I]�Y��^t'Z��/;��zϼq��eb}�p�a�\����\3I~s�LJ~EcY��y30�����5����wL����I�ZmG˖�J+L�,-t�	�=gP{"��=e	L���,��6�Un����%�aN�c���*�KЫzU�7B;[C]郇ڽb�N�F�W�1��nAFd� �%�e�p���� ��q��	k^(.=��n�z����r��E��a�n�jYJb{
F|]�C�;L�a�f�#y�,f�m�t5ny��k�N�Oh6�W^�+�7U
�|��	�c�8e����At6@�	��c�<���+�ɗvwY���k6���B왺N�:�q�i�>V�v�:�:8i������+5�6o� 9�� 0�m�dQ���dM<J�����~[�r��Y=��=�q{t�ft�[,��V�]�T�8-�t[�����BQ�w:u���n峹�J�-�z�s-ۏ�2�={��}� �xx ..�t��LV�"�┦G<�y�↶}j�} ����Zx]6���lv�+��:T{���\�^]��8����֣�=,�����`�d<�~`� :��F,Z3;Ԟ&��)���8s�X��QL�:S{'U�¤�E��z32���6���
��G�z�NF��M����t�0�Z�\�s��e��V���9�����8|���)MQ��?uô��J�V"���)Ȳ�V�8�z�.83[v�bb�e�ag��3*��b
��uW�C�l������S�G�[�DL����IOu���}�
{�Jw/������L�O��ã����&�ؠ�y�::��Z��2<-�439����y��� �t����ev��Ҕ��m"�˺l=0CmE�FW���p�Ի�v���[��# ۭ"ؼ���`9�/=6vJd,��rϻ�B��g��ҡ�)f�R�f�X�����lA4)�-AT�UY�ΊO�g!�H��X�C�L�[L�̫�k��S�^%K'V1�]y=�ʺ���e+޹ӵʍ�Z�?R��h�('p�t�ocwy(F��w^�,��}5^m�i3���{����^�F,�
�وfM�v7�<�R�o��iT�*����oM��0���:;׎^����zz��T�+u�Ȯ�s����K`tE˯�k��54,S���+7�'�����xg;��ڹ�Bʛ����]D������y�'���G�uggE�����u���;��d��8��C
�r�E`9e��cnҚ�s���J�������"�Y��)'���pR[ �qB�r7Ζ��f������J o]�F� WJ�æ�Vи���Qi�5y�Y��������S�s�Iw���׈m�c���=���t�Q�4�s�&TW�r9gy;�7��ΝC��y
!���>�ػ�B"������DL���쬊f���ϵbw� C�wR}��P�;�������ýQU�U^kw����4Y���\��ז�n�C[O�z�T�W���� +j�8�N�C4+��!4wbw��n����)S��=ը��i��uh|��.�d"Z[W(l��.�<���k�L�Y���ħz�١l��'\�Ճ�V��f�Z�4��Z��=٭�ݛ�璕V��ͺ2> эN����\��7w�:��W5Z�Ar�]�Lp�V�V�ZY�Sӫ�����	K�R4P� .?SĖ<�*�)�b�]ʋv�x�6˷��R�x��5���O�b�(fZ�^��֒��-�
|;��$�]R��:��`� 'ZŘ����wA2�����n,Y|;Z��Zf|���y�;��e����ʵG �[[{8���/�24���m�i:��i���M�{��Tٛ��闤���h�ДA`�R�$����J�*g%��Q���>j�v-:����
7gv<}�\0�Y��9yx����5!����w8'�J�Xo������uM)wa���nV�9*)r�=�ﭩ1ZC��%Ʈ���W�{�;�qts E�t�����]Q{�HwA»�q[昇��A�&���f���N��t��R�nr�����-�;�]W,+�*׵�$fP5-e��4��]�ku#�Nu9���KIj�{��54��1]J�����h�U�y����S6�õ�qD�r�i������{F0N��Q[�%��'����/�lL��Vͷ�vX�M���Vc��\���Ğ�br�KXG+�1P����Sd�jt��e=�Y��j�;.ʹMi�%Nǥ'��g\��˙WhI�Fv�v��}J�{p՞NN�c+�����\�*˓��55Ղ����V�^�����
 �7�
.���ԄC0�t�k:���e���t�Ⱥ�t�����/:ҽ�6��rR.�L�ͦ4�7�4m�+snRM�g��!_p��˳��3!�����ӳ:�[���*���t�%����qN�u��(���9[|�:�}x��{��z�ٹ�Ow>�Q¢sN��M&w�tIE�H�z�Q�
.���ߦ���7�������q�zR�vQ��D�R,+Ne'L=c�]���7��|7�P�ҋH�jH�e��Fna�v>t��<�塟w<̡3�V���G�G-M".��y�B)����q�Jڪ�ja$��E�'OWDA>�����'-W�:��:.�M9T�BZe��r�I+^+r���4
24ʄ(9qP3m.�Th��t��q֕AVFi:.�䝗s�;�9�t/8��Lʺ�$O78�H�����U���V��]stZE��ʜ����q�.(���E����w[�70�"Ϋiȿ�w����S��̽���h-o���+4�Sk/J'.��N�]�o�M�F1�X��豽�o���][�t�m���f|��������m������~�~����'�x����^]�=z_�>P�4�����fS"T�.~+��^&*#X��z>qw
����Ю��r�فC6n(6�j�,��C�n���jf%�A�L���;2���V�ra`�K��C����*�@a}~�����uZn��G��iHBsJ2j7s#�#��MR�,�4��*_��2yB���n@�4��}��t[�4�.�U�lF�1]j����i�oO�0��G'*#��q��3��2��	אŝ8�݀v�λo=���W�A祌�B"1�X2�|p�kk �U-V�k��Tsr�P�؅K����g4u���E���]�y놡L[�A:�,��"��!�3f��{G->�J��	��
��`�ˑ&{sq�-�DRlv`��l�b2v8�qg�\ṛg݆�:���t{l�e	�X�0r~��n��n�qA�5�!���9�,����\�C6�e���`P��	�5�g�qKnl��_�2v����3Jd�L�����"Q�z`CG�܋�b�[��+<.W'Y$˫d��3U<����v��Ts4����E���]ݹ��㫥��`���3��E�H�bѿr�����\5��
���<۾n�(��]�m�d�ԣ����6�梆�� �AT�ܥ�.�R}�״�_@�m�wEL\��zQl��\Au�j��h�v������� y�� Y]��A��%3\���v'�w�mZZ�<�R,ODm��8 �iq��l=]��4�;�y���ކ��#�
5>�p���.+7���v�L6���X�T!���(��n��u�֩Bٮ.���:�ï��^��CQ�ɬ`O'�u�ԡ�YK��lW$5&ܸ�B��kF�leŦ�N��L�Xe����B��)�L�����Y����Q,�7l�q����u����Պ^�s�o,E=��&B=f}Iu�%��W�-l���q�.���D���G7X�ˢ��;?v+.u�*(��X[Bڨ$�5��c\Ւ�o<�Bc��ّ�7��K@f��R�iw�q�2'j����TZrquڵV�[������]3�0���{�&X�4�U��U�Nt0��@8�U� wE��`"�;�|�U�f�jW"؍pn�ޒ'-wt�;����Ў��]i�AL����]����oK�=��;l>�%�MӍ��r���
Y��<�j$�x4�b�<�}֙h1�L��|�R)�v2�jBr�:���Dm�Z�\>�m(��V��sJ��]�:t[I��_:�Aj��/k6t>ʑ��%@��8��1u,�G�8/z�,:�ޮN��K��8K�ǚ�/-�7�������{��靚�q�LD�ukȠ�.͉9.�쾭����^��ź�e�A��s-���ְ>�y��<�`<=�
���E}U���~���O|[YC�0v:�>�W�zסdU��#��Z5���age��zc��V�ҹ(�O+��}���w�ds8b��.;PǤ棛�Li����*��Ζ��І/s���J2-��H}^�3�Rz`Q��hv$psI���zl[�&��f�]Ñ�^<�KO+��k���~����Z��?gґ��dﶊ��k�!���j���g���u�V��($� X�܏n��9�v1�I�sئʡ	<�
2Ӝ�i�t��$����3�[ʟf�
6P�+���������Z�v\#@�v@ۦ@XJv�wD��߈9�h��r�o&��'�Z��ǩ���/im�ܢq���7c�V��̪�t%�8�^n�6��=�!��wyf��.Ȯχ�}T=�Twq��#�e8��s��@M����݆�4w]Z:�A���yG+ܮZr�T�i֮�{e�[,Ű�>�:�L��P�L��m��Ú�l��{<���-��\�:籗�l���M�j+nHk�AF�X�vYj��a��X^c=���)�K�W�I?z
�S������P�k��֢�^Jn��,ɓ�~Ǿ�s@ܢ����ŀ�f/oD��aS�(�z�Nn(7+\;y����5[v�X�̀�|���Vk�T(&Kt3��,3�����|>���������sζ)HfX����[�c}:ɶ:M��e'�O�)u�͈Y#k��yU���V�z�F��pY�� BR���'��@!���f�ܥ�3):��2��سV�L��V$(�v�-�]^�?l1�ܔܽV�Ά�,,S"�n��[�y�y��I�q�LS��9B#�C�5�MMe��Tu��Q)��V�������7I,��;*��üo�ٶц��܉OK��QGN���n�s+��f�Jt2\��|�8�pO ����t[?;�=���k�Hf̵(���ܽ�U��J�.7K�6����↡r���n2������a�r0]U@Z�S�=T�Qh�iy
66xz{�6X�m�c�^M��a��q7���Y١5hΡ���j�[�&!�_P��IՊ3�>�8�o��<�_�߄k�9[fW����Xk���"{��e��͚���� N���?+�Bm/��K���k��[�h�vucn�>jhz"�Ǩzu�sQ��DL��⦲J{�mq�����݀�{&a��#�*�Ὗ�/ϫkw��:��C�8q��t������R�]��j�5�,��S�Mߟ|��'-������X���Pn/�����y˝F��̘��uF��wC\�62A(S�$S3����]+��F���Uۭn1`�DH�ߑ�wYԂ)���#�}��y� 7�������ܸ���W��ߟ������0��r�hO�﮷��1�� T�Y�������0�vlf��؜l��#7�rP��8ѡ9�7'L��rئ�c�HmrGSc����j3}��Ba��'f�>��B�.D���[+��T��P��E�	��Yb���V�~kM�����.lƿV��y���>s��"�@����m_�X�S�@�,���.�6��fX��^���$���R�g�l�����'DT@l�C����^*���3pT�~?{tA.z����~�"Xe;�����=9|��y+�a]�on�V���M�PE����>�~^[C��$^�d=4�v#D%T��ז�Zt2�[�"��h�h�pe��	��B��cY�ٷdwpn-�|����f2Ef�׭	��R��*y�w�tV'ђ�B����80u�v|�����2;��͇y<�s��H�E�䘘t�v�oP�v�P���ܗ\B��CTl��_���C���,w��2e�.�޸�귳�◥�H��Ǯ�[dn*-m`�SYX ���v=�?��dc_2J��O|�u['gf!�\T�-�pW��9oF���T_��A\������$Q��f�-�7�)w�%g�u�ha�[`�y�T���jߴ|�ݦ��hHE�&m�ZfI���H�,s�Ml�[k2���s�Y[[7�b�7����N�Vbw,rZ�Уa��}_>_|�o�eKfN&���?y�Ph�Hy�~�0cJg�١[��p��ᔽb=�x<��4�p�4*��
�.��4t3�`s�[
�pF��>�(���"��􍘤�b�y���*����ciy���r[f'���O�A=��8O��r�dX��Kֻc���سJ:e��]��h�H�M���aw���i=1a�0hlw"�K�l��WrGB�ێK���Ýˆ�;6�spCP�]�����^�v��J)'�
;f��0LQ��걖c���L=jh&�~�1/a]���feT5�ʝ��R�7���a�'�50�l��@D��ãV�wK9��bqa7���^8� �\m�_�R�q6k�h�W(��Q�a�/�̣��f�9��HI�{�\ek��6���DV�0�~�"YY�a@�������a�4޻�1�C11�Է��v�-�I,�mF��S�PCC&��GYi> Oƿ���l�h=�:5��7f��[-ö�t	�Ny�.�Nml�l�%7�w�[a�6U##���NF2m`��΀�;�����5��fze��,0Oݝ�϶����)Z��A�ҿS:���K'�%��g��her�=&�%��>�؟k>�dc��>����9�\�r��B�r��	���j^�l�GZ��� �P�p(%�E�z��p�@n����xx�������wq�K�V��0��$�c
N?������/k֪�kP���ǲ�3�0J2�렌�g�mM�׏q3�H^L���t�^˂'�*,��*Q�t�\��(u��lU����\u��f�?4R�[Y�Zq�nh ��M�^���c���Y���]��^�okc5�S��1�HJ�k$�:D��0_t�Gz��-:g֝�F�GA�ڄ�ɽ���(��+]C�!�u!�����o��=��Cʻa��s	��З�t^��c�д&���N���z]��ɬ��}ɕ��j����/�z焭�0�u�qK _\qC��m�r��u����Y׬u����9P��%�)��htT��z	E�Q�h�@�`sI{��V�hF+����c71+Y	��{#ا���6�`/n��y��34\1�_<���z;�~ˬ�uѽ�nu�aE1�b
+��A-�d��z�Ŷ����`o���#�IW)�t\l�l%����;6��v�c�q�o%��a����63���i�����Vc��ܝ��fZT,�l�ڪ��-j]�L9u�ܦgjsz�)�_]��u�	��:����{���qS�BEN����Ѡ}��e��*�O_�E�[z�m+{Ռq,�r�.�*����;/�R���Z��ܨ����ؽޝ���A�;2���
�-ə�8��m��u��￟���¾��="�wwrOU̥��Uӳ�ݛ���G�TH��v��NIOS�z��ŲF껇��z�J�\�Kr�nyD6âcC)��/ɷrڢ����6z]�N9CL�E���Q��U��'��������ݵj�f�{.C7�B��l��[c�c
jj����{ �=t�/:�v���}�����$�E4�T�եб-��-5i��YrՕ�oU2ܒ*܌K)`)ޅ򃺅X;y��s��G�݈�-n��W��4�\����4k�bJO�G�w5,�/��mׅ-��g�8����&�\x��.ݩ�A�0y�[p������*M7C�U"��ʪ��bU�z�vf�N����/t^]�9�O�FA�{�x-.9�������ބ&��g+�z˵����h�)TT���ԡ�Yi��l3����r�o�i��<=!Wp<2�+6Z:��Ĕ�q"�)�ի��������N(�8ArZ�p��8tJU��I�c���J��5�d־K���(�F��:�.2��]<�Q���=qkM.pސ��]�lL0|i��-W	�%t� ��D��;i���_�.��l�̛귩�<惍4-�@q���+�2�6(o٩fW�Efś$
c��W.Ρp�����7Z��z�F,�w�g�:�E�����8�s��m��s&>� )p�ŝ�Ѳ2�u�M��{���oxy�� 
ݨ�����7��-=	�IԼ�����$ڡ�T�ȯZ}��d`��{�]�r#%�C��T7w;M��1v_�l1���G��
�f���MΪ�-��6���$���=�d8ŵ� A]�n�Ѱ�gq�n�+�`�nnv�Ǿ0�B6=Lhl{mN
�D,��H���L�ٝ{��H��#�斠6��	nz��ipp�;���,D'�-���װ�2rX@/}-�!t����]ЕӉܾz����H� �X��E����|u@t�4H��6�X��wJc�B����7Ob���@p��y:a�˄4\��,c˪Hhol9���3�ݾ)��<!y^�m#?g�	����l�3Ck9L�|�y�R�C'�KM�T�e�sMNCM�uR���1A2��D6>��>�C'n�+ٯ�L�ƴT�~��i�X�X��UQv��έ�6n{H�xM}�ʣd��3�X��N�M�i��4#�K
�t��l�Œ�a.�W���N��p�7� �s
�Qy0(^4Rz�Əi�v��	�=�CG�Py�����/O64�w?b¤�d�{n3r�eV]NK5)�L�^�,�NP��q�O8�����Ĉn�9ն姣+q�r��|R���+Y��|�V�m�3�sgTLz_���i��g�w����N�Ԏ��^Qb��}����x{�e�J!Sv\���s����qT�ܟdڧ�8��*�L�~PF�麬�>F�12�S���7�Ϝ9жY�����ť�J�G��pZ8/�(VtT'c�F��`}�q�W��t�^R{��])����a��ȖS�j�;	�B�Uד�q]i�# ��㤓jk��L]�۬��!a3������b �vT�n��KSԪ���
�`9l`S&'��:{ТS�y̼�^�X
�]�����s��0c�lЭ��߱G}9�䡋�n�郙�7�0/n���G���u�Z�|e�='�FwP櫴(Æ"��\Mbogf5����YA{G������XW���O	���ƞ�gq��S���r����)7dm�Szzq�z�OY���I��	����`��Q����'�0\M��i�;�;,\p������uTf9�6U-i��������V�3j�n�v�vr�v�g�;�74|R,ODoL�9'X#u*� u�#8\DZ�>�f��UCP�N�EI����i��;�)����G2.H#�g �mlb��X�+��7�W�R\�b�ͩ���P,y5��`�q�N��
$��b�Sx��y��cz%��Da�,���t��N��P6]4.N}j,|�+´��.��)��̓VtA�r�T�h�";��[y��0�O.�ZY׼�R`�ћ��]����}��b=�(
�,L]p���]{��uf_G̘�-�o��5V��#Y}�H`%�B����У75�X��&fs1�OCw�rTYӲ]�_fe�j�\�S( ���M	������i�ӥ%�k�fS�{]if|k������:j��s�$��7W{�VL��������\�0�x�N,7�7��3�°��M��.��{�����
U�q�u�a���U�������r�N��O[��F#w�ޭ��J���|84�D3�f�1��S��'s��.W��=�T�=L/�n�$	'>٥:ܭ�P�:C��[�����k�x���Xd֠�c���'Wu�,r7���_ �c����o�͡5�zWVl}]�kt��&���}-����ɑ���mt|^!0n�MN?��!K�:7��ݭl���.��]ZѼx���-�R�:�S&.��u��/�=�!c�]75@�{�l��]�ا	}G)]�t�&K��d�*��ǜ�Ȭ��v��S� ��u\+����Lu�LJ�)tO��=w7yc�O��W"�doH��� i�+t0.��]M�{Q��ɡp-8�#�+n�G.�K�ĩ`
��\��>�"�{+[����.lR���y�]��0��iڻXT
���%��Я���gZ�.���F����6�l�^8y�����k3*e��T+�dr����^Lt�R��F��\g���{��+�dDe�u31��b�6��R�Ww���v=��o(l�6�ؗ��[I�Y+(�Pܛ:��E��g�f!���b�U��շ�ʲ��3tխk��%ZvU;91�F��޾�/8�Y��RĂ���V/UaR���թ�'L�2$A��F����Y��@K��z�Zs"Ɲʚ��홆KԮ��x��K����n3��B��ש����W�=���]edұ�`�r��^���K�+3y�o3w��GS��>Ԝ��5�{!.
�kw)�|��2C��E��D�ʱG+�>bu<%��#Zʝ�^Y9Z����j�U�R����WD4va_1:�Yر�*dٰI"�k�1\�b��[�n���%��M�[z&!�OkhI&ئ��Ӏ�l�w���f��e[l��r+��eqwE��vROJ�֞C��Mz�fO�/i��]�o�5.���q���hB�'.���M�Y��0�B0��ie[�)mҔ�+��ݤm�����Px��7�FI�|����n��Y�`��)	#:&�Q~P�/��L��L��MM�v�7��|�2��Vh�Uq�Nt�L�HФ�Ь�"N�f�\)�H]r����#8U������o��*�����9�e�;�t����XXf*�;4(��宅r��3΄�DW*�W�I�h���^w<T�Ny�"������U�eHJ���wW�{��^�I(�U����/<;.E�Y(-tiPS��wt�f#SHBLOq�Ô��9���D�̂�r�N�B#<�:�Ȏբ���vܨ(�6��x�b7;�N�=���)�b�K+�*�����r]5���{��:�zG���1��3�,�=͑ꈢy��VB���nGv�:�r��rHI����KG:���=�uJ��*IG9q�w(�̲e'((�W�W ̕z9ϋ{�n������He��.�XT$�$�V���Y��ۜ��-���9غ7{�rI��L9cq�IV�*��C)��-��A�����
�����5D�Y0q�N(A�8Ϗ��a�6�"=�5�mɶ��U��b��IfO2���4��.:.��=���ި!��ӼO=;�z��yr�]"�eԂ�k2���iu��-{1��y�)|���.a�ybLp��Ho�E��~Yf�
��C�VK;�*|���=f's�����.�G>_q'n&�6�r���FH�הz��E�y%7�ѱnr��U!��d���K?vm>�����"�z(`��|�����a`>EŇ�(������˨^ښa����U�����k޾7����o�ne���'N٧�/e��J�Y�@EE����#@���e~���ҫn��	Y���(Cb���Dc��%�E��1�0D6Vj��늤_ٜ�}F�c�j븺rDR�Q��H�B��m�*m�`H����lv���#�φ���Sv2�-��'G;\Ig���:t�](�C���p�@�K�P��wm��:��r�3Ε�q ��" Xu�j���Y�M���U&c�9z�Ϸ�]^��6�� ~�1,����Wv��|�#��niǥ4-���\E��h�pR�R���ȡM�fc�+L5,' �/)
���b�2��k���]E�&�uK6�<���7mE���1Fb[����;g[����+V+�z�h�]����|p.��=R�e+���sk�������������|��=�Y�����+">Ǥ�2yP���q�41��F��zT�5 �XgOE�6�$��!�Δ9�b8H�l�9�5��=��6�9�8��;��<�h��q^sb\�M`VW���;{|�Y�2��<�.�NX���F��n�s'�;��m��1�.�ڃ_4naR��FT^%�^�e��A��ɽ�Ȯvw�B�}0V���*?KIf�ߛ��i]�+5��1��X�[��n-NѠ/&+z)ʟk�bxfs`�CT��F`͖�-X��Vi��ё���[���K�]6�I:a�X��QD�lQN\n�6zٝ���ʙ3֗�y8ye�/�YMn͏�/����ެa^��ˠ����l�Ӕڦ�H�W�e�Z�ź���	uAje
�y#eK�&<�Lϩ��>��X��Ai�a�,�j��7��[rlU/5���Q�S��h�����Vx�
��Ce�J0p�������Q�ܲZh�����%Y�j�Ӽ3��<���q̵�%�A���ރ&`����-������BEN��¬ݼ��p:B�_��G��]����vV�-Z:Lt��t�I����P�Ӆh�oegb�n�
�[{���(h��n#�)��w��Gc�*����ۅ�y���Dvo"t�L1/.�E����6f8��m�lN�;&kaw]�C�����w0$ΗY�QdI5���}�>��� es��E3�Vۅ������_��g]��2��`����7M�Gj��3F�T�m����dn��h�X!�r���o�a�_E�P��GC�0ŐM�At5�!�eX��l�8�s�NP���aF���Wa�.:ͪ�
2[� �y�"$�����7RZ���d�r3�)W����	����6��Fq�TN�T��ө��w8�*p��)��Av�f���1K`^�Z�z֛[��ӭ53��QL�;���$ڡ�t������@��Z�����OT)�Owp��t���i3a����<���#Pb�h_K\K&Q��nb��xq�ksBG��`k&�5�4A�\��b�gp����F+��2/������(�e��FX��Wr���Jk�u.xl�k�X
�M�Q�u�D�뚈��0"�*p��3qȊ��p�z1G]ڞ#_۞Oe�OS�lqv.�Cb��
�`�9M�'��
�w���߃F�w�2���˭�������4K�����S��"�z��Ȧ>�Ō��zT�,WLշ0�����S^�]�q��vR��M�/��au9�'(� �	�Ɣ���J?��eOw��վ�lh�k9�3O���EP6ڞ;�m'̠�:�*R�K4��p.u}�9�S�	�]\�6{[����K�U�j��z�̭۸���j���<>� �o ='v9���3��=�l��D6T���U#F&(f҆�L4Q�A�77��h]�&��ˤ��E*��`D��9��_�1��~
�?��ʫ��r�IY���D���Kh��o��j#]@i�U�5˒�0坃C�|L��K���CB�mb:$�i`�pꄮ�8�}�%��c���cuz�(7#;��nU<�a��hvAi�r}�mis�����9�:��'d]yL!��$^������z�:�Ƅ�A��t�i��?sA֨:�w��Vێ/^�猢ጩ��(�O�cTsh�c�Bpa����M��ι����*�FUh}l��$Ѱ�8���:6Ը�{l�����D��H�zT[?<��#wWYX��6���d�;O��,�1A����.����ؔ@�N�S�'Ѷ�foX�:�KC��W]��� xT�*����
�s���ޟ)���� �n�Ц�Q��2J+��#�j�3�N������6'�#g�0����l�;��@*��F��-fQ���������7~/�z 7Z���ug��(�PY��e�N�ݚz���]�]���
���	�'D�;g\;,lںub-=1��]ȅ�v�q0��=�����@*c\Rhf:kiν�{�zy�tGk��E���f���_>�����=�Df��ܔ4tb�(3E�*}��~=�A��H=r���v�3Ͱ��%�C����S��f��v��φ���r�z�z\��R��F1���޼Q��D������!EF�_�[������6�ӽt��ν]ά�}���n�A��.�2[�C[$�~�(�qY@!nш�w�جAD��Yp����c���h�ݻ��a�8$2F���m�����ʾ�������z��Au�����'6K�aZ�����ˉ��^Ģ�eCba7$�Q��������{V�Z��c�2���O<�J��g��9��"X+ڐSϫv���1�!�.��������&�tt�����ɶ�ʦ6VV�Sb�r�(�Z��Ш�ꆹw�$V�lNK�y�֪k7��ط67�b�}�@���]�(��e�(��h�EY�J0�x�)��:��I�!̧�及�j`-&�	].ݻ6�1�-�J�ҥk�����6��~���,Vq.i��~M>��˵������~p�O����gk��J�Xs	�>aR;����F��V{�:|9���iCT�ymQ0�|ZC�,RA��`�a�eY�ø�4#|Z�������S�/z�utS"�["����;7J�\J��l�Ŗ���{�S#+W��چ�x�z�WPox:��.�e�2�;�	x�SnX���-7�.1 �W����C��}��Wˊ�16���nD7��4F8U/����4!L�w�$M���*�`S=�r����Y�������P��l�r��������!��n����ã���:gqCH������{h�ڝ9{��ret�U>���+��T����ײH�q������pcO���Yw[=���f��]V���R.�<�0���6�[>��LW6kg�k;�w��>�ܞDstlð�B"r%)Ɠ2���{��R���zs���L�q�41��#A��>y(��0pܧ])O��,�<�]#7����D1���|�ڥ/do�����}���c��ص�#Rb�ot�,��`��*���H*Z�t~�``󝺧�[��s,�]�'0�>������Q��n��*�q�3����[!���v�O�,�������Șk��K�n0Q�-9k����Y��q�,��`r� �6�����S�Ƙc[R�qȸ�-"��y�Gcw2E�bv[T�A%UZ����0\[�_�Eu<�q^ۨw=4�	Qͩ_�X=R�~�.?�T���53Rw=R���L�?ʞ�~˲;��i	Zj�+(�9��W)�]:֮�[���Φ������C�ǍN�oz�
w���0����͗��6��������N8�c�����+x杽��s�&LZ��e��V�T���T>]����7�xz�WԔE�Tj��P���u6¸�:�]P�M��[�+oܫSV,���:�����*/�jvU������0=g��?@������K�C;�2����Q�.��5���$㩱� Rj$�T��B4�n�͏c�:؆�I�E9fRr��P��E��fQ}��"C��-x��*�kSۼ�6Q^J�YW��NK8��c�͗�f�70v��`7S�5AN�]�r��T6��5�*��Oǟ��b��|$���������cJ�!ina�r�"�]
:C�b������R�aLR�(4�0�#i�[lˢxm2uE����w0m�H&��Cb@'O�+t�/\�M��3
jǔo��6�:>�j���H�du��$Z��zj˳�-`?Ef�;m2lYj���O��Bq(	��-^����@^c �V-.�.2�˗B�w8�*p���\�?VKAS���kA�3��t̝a(5�N�l���`�>陘���)����-����G=GY�k�4LeꦄZ��V&��9�D�A�i7�����w��y�:v8+f�B1�t_�^sMz�T���>���.�+��@�cpZ����AJ�T�驓P�1�@�f��R�G�e<zk�"�	�lj��9n<Jb�S��0�W7�C�����my�+�C�:�q��q��u�w���#FM��aGhk��h��AP�����M�MS*ޙ������̥y�]A�bq{���y�D-������q��{�s>?L�l1ba��ͥ�vׇFDL��xfO�0�ȑHi��n�@�7Rv��L���i�s��ag�`i��T�ƔD6=>� ��w�;0��wO|k������7]����^�X��%�����A�Q5בi'�M�i�)����
%�H��΂��d��M庈���/9���=�ͅ�A�69�7'L�p���b�%�.�!���hhSh�*���R#x��B|�ꌴ�1�3Cq(�cY��B4����R�dF�����|�*�f����\�: ��СR��A�d��s"}�]E����Qp���>�\Z���Z��[��iz�X�N��5W�fIs�d�2�n�12=K��2AmmF�QjLi�6
��],�m�,3)�p��E��m�2�;rz�v��r������\�; �������wӒWQ��Ь1AvЪ��f��yN�P*�7vV�Ad�~�3p��\[L�;І��L"!��sv��'a�#�gC�d�/���2���*��nf��`GE�%
�
R���v�$5��g-��1+��<�a�����T�E�����;X�b�z;�h�T�ա��^��]J�P\����0���C�+��2,4�;��}�2f'iR4�f-ގ�αЦ],�,qͰy�V5MK�Yb^�b�b+a�kǮ˖���?{�0o7�<�o�J�AЊ��=�"!>5N�k��e=��[�ļ��J�O~1�)�v?n5�@����t��R�������.�]��:���O�D&ޘ���ܥe��>�R��fN�S��d��ᅰ]A�\o�K҆θ^S��v�;!��F�`�t������(L!�6h=t1&Ig�K�3����S���jҧ�L7l�	�t���;�c�a�:�0F��f"A�Q��a�u�A���!������"ڀ�Rq�<	�u�׬�5�jܶ��	�.�3�kZ�|1��8j��n�Q;5�u���i���Ⱦ(�Ngܺ[;�6Ǟ��I�2�aQ��iF�A�1��5����N)M[L jQa���>�.O-"w��}ᔪ~�����P���9U��`G
�Џc����������^�����q��?{�&�5���޼�B�1q/U��S U�����\Y;����Q˦�/��w�M�Q�bQ>��/��ߡH�[4�}�-�&Q�a�ި�x�jF]�t�5�\ݘd��T��HW3����a��`��X�W�>ѹ��k��>�-CyJp�Dݸ�J��:��т
�:��o���v���'=E�ĄJߦ�n�h�}S���/@hS[�k�vA��vf�B�
!��C�_��ѹ�k��opSޝ���W$��޸$�J�4�t�h>�3�����Xޜ������ G�j�S��MR�F%k߱B����M�
[v݌�0L���.#�X.p(U�k�/
'
��][���A"P�d"�!�_^�mהV��ފE_����7�=��F9����]\���̞8�LZsM�yz���D�Q� d����Ψ\Z��)Xo�E���Ek4���6�.�1I`�����N�)r�_�R�h}��~p�M>�����\����S��?F�N���h�����܅ۮ=�ɺ��t��C�npV���4CQp�6V��/T���J�E�=	m���K���2�+�<x���5�����;�ma�^u��cb� �2�a�l�iҦ8h�x
�3����2]��=�AlO`�%���h�"]�1�����(��ΟxɁC/���M���_�v��-%ЎF��%Ra�1O3��O��
Q{��^y��F�%�Wh��۾?���)vC{w����X��F��I�gW�'~K�c+�h?P�t�e�G���P�wTNn���[��0��H��!��Ba�Y�k_Cn+�fwhu���z�,7}�(�5�o��z
��5z�]�;��v&yV��Em)�.���2uK)i���c9��.�����*e�p�{w��z��]�{�q�`�2q���!�k�z^*p%��#��]mk
�X֙����<��X4�3V1�ה�u��e4(ЛN��f H�HsԊY��G�+��^Tb�$�mEe����e��,��V�v.����}R��.>�N��s�v�lƍw�u���c���vqa�he#J�a9rhnef<{�̍�n�aU4��0`Ȫą�;e�ݓ޺Ӱ�-��uچ.�T3^-�n:�/	A��C��-ڎ-xOE]���������Sۦ8r��v�h�Y�僓oy�������rLn]�n-�o:�s�������i�%h�v�Õu�¸��H�]�)ިQ�]
|�=T��i��e^޳��o��)�Ǚ&�X��o�q,N�w7+v����<59Z��qL��pɗtW�ַm�h�%o<��Ň��d9(�\L�O�씚Cg��e��ދ8(��ī��-�s�Ӯ��W��-����_>�ԅ�Y���\�.�A��oJ�̺HH�Q��'D�	Y��"�b���(�j�6�[7���&ܲʡr�&O1m{{�G�)����+u�d��/{&�S<���(+7I�[Ⱥ����\�2�&���]��hX}J��{P��Hk�l�9���%k"�=s�!�p@��ǈ����ZW�³$N�%wp��Z��u�w&u':i�
�{*eG��T_4���w��KD��r��7����x*�;�:9�e���wvW0�ݮ���ɧ����+۲o��f�x�{.���THg��z�VY�9Ay��QrB��Ur��I�tܬ�/7;���n�u�٧��%;��X�(�咇d4XA��`�ܮ}Acf��{,=U��fN����h��Ԧ6~IR�ߞa[�U�93]�#�Ҍ:��[��G"/���gk��ri�b�7��V����ۇ59g���X��Y2���}r����utF�*(N�P�V+��.4٦��Fp�zd�e���EK���Cz_wHPܭ
Ξ���e.�&���	��):������ݩ���U�Yi�qr:]��ԪwM�*�ʺ�5�5�ղ�d�v�=P�빤�d*�qm�;񽱅��9�OEZR��\�Q���4�3� �Fb��^7�Y������j3��C��e�դ��	�p4ܷK�N���D�<B�ǉ�I4]��co9k-�+0�ɽ�kˀvf�[/Z�)KYؑ(�a�ዩ�(��0��9�M)he��ՙ���Ύi��/\uС����f�w�~$�):�E�f!�wl�q]�z�Dx�,4�g l!:�u��jľ�4����Vl�,�we�W��黗.������r�|vS	�Y�{�t�������b�gX��Ux��,;vzK�RU��޶��!�\Sh���;����6��N��~��=k�<y_�:�"?$v���J�%*������A��;��F��*���ȻH6�*��dWv���|�7����s�	�P�RȑfKB) �Q)
�g�%��JH��|�7��/ĕ4�*Ϊ���qVRJ�?+�����3� �t�Y
��N�FbVuZAg���I��b���4�C[N��"�������<���7�7*��V�PU縡Ȩ()""��9P���t��ᥧ�L�#���X��\݋���QғYn��zK]��C�S��癒N��r��_{�㛥ܫͅ^m�L��!f�x:��/G>w���D�Uz���QH���B�P֔tZ�T�����fP\H��73�E�y��y���]�!V�b���OVG.�)Լ�	�$�� � #[��D�>Xs���U��}�op�5q׋���;zȉj�v�(f�{�"���anc�/���ֵV�s���<�a�=R9��7[T�3
�.?����8��.�;�����!�2@�ӛ>��5�#�6@�Y��u ������s�p�ٰBa���':|]��gt����M~c��4/9H���<�٣�5�rw�M�h���0����RA�j�r���1<9�"��i��#��x���F��x�)�6�;C�;��=�A�APC*Ȗ����yM��Ȝ>ʫ��4N��t�]�zo�g���5�%5/;��� ��[Ř���X�c՘A�=n���W"r�V0��umD=�#���3���)�7���`�A�l7��Y���fS�1黩��(gs���O(�2˖�3��-�BY���qE��$���#�C���&Î@�59f��W�[̚-o
SU|��!�c�bWVq�K�4�6/�������;�o32K�Թ���h�2�K�^��9݊/79��M�Ҙ��=H���_(�C*��皇�:.��w�PZe��ӱW�\F	xԏ]�M|�TQ���W��W�(r<���t^򅆯_�Q�f���Gg���܇��q~�}�U�}Y8���Y����f�5�itP�f�iӥ�XV�Rb�1��!� ei �oV��dKn�	h2B��ޫ���p[j"�N��]c�3ֻ~�p@d���*��g�{��l�H��Y���.h��|����G�*B�P�_��+�)��{����<�a����$�4����&�/X�|������їf�hn\��~���p_���,O����2ϦgWt͑�c2j��Bb��t��G�;8ػ%R�x��=z�w8¢ˈҮ�U��7s5��-�+a}bX�3C��m��\�'��E2��[ěT0��X7o�j����u1ɺ���s)L��;�aіn!��a���1�0�A��஡sL��)��]�\E�+r(������T��oW��A�=3'��t����:DN���ҟ1�OO66�һ�h��
��֮�C��^~.-�
�M@��C��Y���l68&4�nzn��h��7J�p��N��v�ۻS^�~D�j�L7�ښ�E�AF��V�/��Qq���tC����蘳qc���R��/`���T��~��ئ�c��E�Ͳ���ݩdm��lrD�b�.<q�,��F`��9W47�ljP��BԄ�(ե)�ϗ���/�L�g�� �ƑU�O�.����S;�z���Փ^-�
m�*WP���}�9?v�{}�'{W}8����k�u�ԜnvK��J�4�e]L*��K.�� ��r~<׺��=�u�qP���R�Wbꊅd����|��JwkԖ���Qt��[��2c�ד�cfzv`��gW�#���R��$AݭC�����C׍�f[]�2��d�3�)�4~Ea��V�u���pB:�A%dn.w~z�9l��a`��,T�9��C%]M��rz�v��r����/�K�Ǜ��KDѓkOd�d�M���2��;��E��Jt���ۼ8���Γ�m��s��ч-�'�9{h�MNѧ[��so��K��J��d�/���2��0�Q�a�ĝQ�m��y5L�����ٹxD��\��4�7 ��;�>�I���ȖS��Pޞ�b����K�zy� &��x	�j����n#Hvƀ{Ks������ͦ��>kQ�jWM�De�����<"i&8�m�t��E��#'��͆.�����1��x��\�`��j�]�*?�����uA.Q��'�jTx^��-�.��(p�B=�E�_�_�/ܣoϔ�vlYͻ���9j|�@�Zz��@�ȋOt	�vG�,��MzA�w-\�˻6�a(f��Zf13�UK����2s[n ����hr�ŎzC2��g���#����A��k@ĵf��g�,1[�\�h��ޥ$\��P	W�2a�u�f���nܝ�]�rw��CFX�%�PWH�7m�~&��N��ެ��緹�Ě��] ���	��;��w]nڸxWS!�P+P���k�<�D�u�R��>�22z>ۡ�_����\������p1�>
�	�¢�ʇl5��ݽ����8-�	i]��v�#��BV���}�<X�ٓft�:62��)z�����ɍ��d�����F=M[�݇�PT��t�ͬv����a�:N5�l	t���xUy�>@�{t_=5꡹5�	��Uŧ�j_jv'W���K�82�TH�U5#.�.�\��<��H��)�C;ӍZr�R쾾z�#q��������1i�ɲ�z�F%QbsϊqˌiN�&���֒C���\�v�u���N��2i��}q��s�yO�#�-�����Qc\�r��ހIR�2_of��D�`��d��ނ2ΰ�m�N�\Z�B���Qi����껛|~~iO2�ɍ��RØ���@�ϲ+�#A,�Cy�d�"��=dh"7R��.O3É��ܝ[KAv�x�h#As�W#�UІ4����t�Zf0�E����ힹ���"�D@���;4�<vUr��Pu�'�r�m��r�]�v�K���G�lxn,�`��s	���Lޛ�)��􋇇}S@3j쬘>޲�4)m-�N�f���ë�:{H3�B0�p�Ďc!�%x�J����v=B������W(X��^���/.��2�r��֨��7d"!�%�]%(�˵V��Mw��Q��o潷�`��9Z�P�q��7�����0v�y��rI�6CǠ���f����d��WT ����)7�&.M�@��;�)�4ځ7��Y���f�i�?t2T�\�OE�;��J��lb�g/kc�D���_8�}�#�n��B��	nf�Z1���)�k.Q�,��(�:��ۜz58Б�m��%Uk��213�Tc�*��g}�v��!�� [�=Ĉ�h���6}�������m���ms.���Z�ףX����E�/)��� �z`���v]�v!����a��p4�Ƕ��߯��1<�����!'My(Ǽ��L��-�[�P���Q�0Nt�h���F�xz�n��!>LG�]N���T]�5��C 9�9fO���ʤ�ڢ��mOsa��CTuT��E
YX��yzٹ�.k.I�B^�ŵ�����5fcA(A���-��I*���63�Q�7�������D^� ����,�EP���u
��++�ř�Kߋ�}��(߹V0�7�v�K[(��k�)��w+��V���9G�S�3Ǒ8�76|���
�t;Mz��:�UG��Ƶg~�e�~��H̒b�X���[�$]ˆ�������Ǔ��z��aw�m�23�rl}4��&�ɕ��v�up]z)�Y��,��U��' ʺ��0�����}7n����^�M4�m4�k=Qŗ]�]K�r�/nu���P�/�����~�����3��k'���qv;�����v=A���4�N41��[5��ԣ	f���kp��n\���.�$��&|Q��/�\��v�����C�H� �|xb��!��;�sD5em�Q�z���fA(�(���!i�d�����)���[N����^r�Ҫ.��?i���h�zY��!�0�+^S�映��S	jSr|1R�v����P���}HÒgwg3ka�q
�*k�8ʚW��j`&%�c�<�'�U�hˊmW0�d�8�0�1C[>�(!l����ĕ]�v��+Ĵ �1�)hw.Z��2�����b���j�uoL'>����Յ�����陻4"a_L�3*���j����V3lg`t �|ש����E2���-�⡙��v�6��	��m����t��@C��5T��9F4<�Έ�8�q��g�=���d�SQ���vɰ��t]&dE�+��YWn���M;K�Hqё'g��A��ܣgz�8s���eltte��,:�pe����Z���2�p�_��$=8��e�\,5\'�O���B�̽L���n�G�Z�r�ܜ�h�ri_u��t$cJ���ƞ�XT/D7L*t-��W��P���G�6չ7�P��t���Sz\�6i�4^ZG�T��0e���p.;�'6_$r�!�5f�+�J��ʸ�<�5y���Go��(�[+_Y���:s��~D��d����QA��Q�s�UɁ�ٚ��G���|f��
��9��ۻ2�ծXÒ���4[\0uGΣ9kpN�I�X�[RCF[V/r�3��8VCb�'[��w�͍k���$��p�=���Y�qhݩ�6x�T�������Ш� T}�f��E�cM�����WfYk�A��Bi�׳��ۮXȕ,_�b�e�1V7���ld�1F�Ze���0�@Va�"m-�O�ޣ��(s����wD�^Jd.<��^�!�<��ݦ�ʗ�l{4KM?p�"�^-�8IDOC��>����ٲ$�'���]��]��9MՏ#3^Ek�/O;̕�������L�G��0k%�֭�cݽ+�Q�S��2w�tV'Ѿ��z/ɇn��s�_d�Н��3�i��/�gwGƸòٳLk�zGa1B(�\�\�6e��2���I�^�)ö��42È�:q�D��D��82%�H����*e�qIje�w�a�x������+2*�w{n_lc��l-;�T��ZH��h{o�l�"�k�%��Ey֕��:�]X��]����	&A����Ҵv��z9R��NrM�/�X��PnV\C�s^#���0"��5�X��j���{&e.��C"�����{�z{��ǻ=,�(	�(,V-�*]��b3�a'v<�<��|�����K�&U]�Bb�j#דʬ_%2�j4�������w�D{|�t�hT{Ύn���h��M8�e'���|ٰ4�����#[���ޓ>�g��4�ק�ܳ�n��/\i�]ҍ�A�4L�)��]����q�*��k��!۩�(8N"c�u()�O��TE�׫/W�3^^gvl$��b�[�N���~�Z�<��/���Q'��;���ibuӕ]�5ꖶv��*�~SW��.��t"le
��9��{uq���T�iĸ̴-7Q��k#���]�l�D���#c�J3�I�%�0�-Y��Q��ȥ�X��V!���]�&��)r���%���Y�TH��rCCZzI>6L�G0��Φ��ߗF<���n��"Z�R9<�ͼ��ΧZ����x�Bg�̎�Qbsأ��,19h�'@�(�3�ֲ�F�˚\B"K�_8-�mmq�'ɊN�}5E�+�Kf�f�﷭��j���C�s+Z�FⱰ q��}�JZ�*�&ٻ�܌�J�r޽yƮ �U�I����P�M5d[p^�[\Q͗yX��h%�C���	��o�xʅ�l�ڲi4��lU��V^^)��Z*.Rsyַ�mk�wsKI��-��ʈ85ǋ�CsA @������/���e�D������&��Gf�~JK���ݯ2�'�\`�j�7�Ց�4�k9�:όS[��o��Uw4�\Ki�xw�oSl+�*�i�x�Y�q���F�<dډ�u� υ�a�Β�TT�ΛN�gU�^�}��q�$�2w�s�]Ϸ�#}B;G�ge���?+=YQ��r��G7�c��%�����UZ{�t"�ڳ�k�L���~̨٘l7}w����d��>�G�:�}�]Ί¹�zVc���"�*�q����U�̋]o���p٭ 1��ײT�;@�-��c�/3���b�vɫͽ���h6�o�c�������f��]>'ܚZ���4�o�l���,y���L�,h1�l,,%�����"�)��\I�1��_���^��\��KP�U����� 5e���uE�Z��������f�C��k$�v��\��pߜ�~ ��6j�xR��Ԥ�i� b�cP��p�e���]fP��G�S;&�ལ�[Q�rX���Q�[���7�s �v{���=����:�v�#���a�&ۮ�ƗZ���m$�cDS�ݡ�lfd��M�
Cd"�
�jU:�M��yO
0��]���݋��E�H6���i��/"�y��yNV*�I<�1�`|�M��N� �#x�q�^��\t����R[^y�'+������g���=�p�~��SI�T�E��)���r�Sތ*s9,�T��1+/�w���wmuE�'��U�){��m�	�!���	�	d�4��#z��G˝��r��RK ٸ�[�ݾz��r�'�BѲ��`y�����oxFC7ɗ�!�$o�V풶B��Pi�}�r�1�]�Ղv�Ӽ{#*��(�������䉔Q��qIE�nO�6�;nl<\�������2#Hg�C��G�n�H�s#�M������aݧ����	���!�gE4!���C-�������ƉJ/�kX����ݺNI�3��/
���:�ʎ;(�dPm<�q�(�4*s��g�;��o+2����pV��]&��U��ը;|j[i��b���� �{��.[fk���\7�Y�kW���ގA����)c�-J��j�+y�t����Ǉ�0�nK��6�r��=Υ�8�[��Rw:�<�i��@�e��j��A��5�͢I�(�U֞�ޝ4M�w���K�:���چ��r�]Yȵ v�7���X���,�A�)"��_��s�C���}!��j'�[�=7��=��y�8�Ō�NT�V7��|�+�ݱee�b�t���b/�A]^�Ο��[���ZX���`�`����k9݌?<�*y�LP/�+sU���R�$ܽZ��U�-p�X	e���4)LK�Xj�qZ��Au)J͕t�D��N�]/����\B�����k9l�z5����G�pp�.��B�����"���N��p�6�omjԋ�߳S�5�_�Wa=�R��3u2tV��d*[y�g谗�ܦ����F�Yxܒ��4�eV�HdT���u/�S�0a�h���W��^F�맍�ɻ�Eˆ�wgj�n4�i����90��FP�>�@txM�㇭�����Q��R�f^�¹S�L���ԫ��)₷&�߃����^������/jS��V��]|�����4��F@p۔�N�pS7�+lh��u:���FN���B����o�'��:�ʃs':Ů�X�"��%«OF��tx*F����%�MGv��y�;53y�k����i[��2ₗ�Яknm��r���5�Ḁֱ!���#^�C���\�´����B:��:�Y��  _\����,���uw�ؠCX�Ҳ�Ctt��Cvti�(�ini9��W[��Mj��ۡov�A�t+
5�]�n�u��Hr]�y8���C�d�g�#no��m��{�K��p��/i7DM��m�n�/����X�R���d9�	��;a)3����V�uڔ�A�($6���5L8������z�[�������b�#���y�W޷W[�
=�#�kV���[-3����[(/+Ñ��#����]�K�xF�Fь:��Bl���;�`�>8�3C�&��@��1>$
T�L��;�3f����a�l7ܚ6U���J� �}L�E��0ntQs�ϲ����_RhS�p�kz-ZnDn�86�q��4t��Ak��.�=\e��T�2Ծ�ȧ2G��ĩ]��v嬸�gj�ck�J�97-9��z��Md�W}�Y4�+���(��D���W(��,��n;�)/r��ۦ��ܮ�W2�krk�h�Y�>���*�`�+��ݥ�v�Υ�!so���p�A��m����6&;��6 �I��W6�|[��
�ͣt���+�-cpr���^wґ�Y�J����6�U�R�b�}�bxݭS����:Aʑ��ins�K9
�]:���7�ض��=@�uL1DAЪ#� �EYR����i�Mb�C��!o��M��o��㻁ew��)[Ԏȇ	<���2�s�V���n�7��}o�|At�J8�%�YDVa��J��M9���o:E:�$kN���I�^�iOqe���*$2*P�Q�4�t�s��ZS��b*Gw��*F���d�=^�ϟ'+솝:�y�Ui���2�]LP��Ӕ�n��D��*]y{�(���N�Iwp��QJ$����d_\r��2I�z8@�Z�t�(�����TE�)E�R�.*�r"HT���x��������{y�k\��\��H�99.��'�E��u"�<#Ѥ]�<����*����(+̲̉JSms�CIy�J�h�U��$��#u��/		�����$hRM�T���@�ll�;�:M��3s
��d����(�p��WBp��F����t봘�a��%��&4n
��`��7��y�:\���2W��[��z�v���z}��+�t��~��b�mjT�ZO��|��7C�ϵ�zg'�� ��aƻqhlJ`m���CC�Ƿ۽SY��C�w?��N�s����"=��y�V�c��3����!�zI�v������18}J���s����p���t�R��H�l4���`��۫8�÷\l��}<�5blO7��KG]���SO�$.kƓy���w���f�[����d^���iC�uл��̧��LIG�3e��e&P�%�I/U�tGf��L���إ� 1T�f�va���j4&*��@�"U�s�c��=��D�r(��`����g��;ś�ݎ]�FM5�EUk�R�"���,���7kKA$�jN׬���Y�����l�]��j��xٜؗ>�Vn�zyq��r��� $h�:�-�74�ʼ�|��C�8���ٕ�#FP�<�M�¹H\y���Z6�VN�}Շ��U��wN�{�<=�V��-��-���.��+��j�����3[�շ��ؓ��w1��*e6v�Vƈ���J$�igw�3u�9�Z�Z�f�V�o���3}�\?@^�8N�S�5H�J�0���5�����*��S����p�x�6���v��	:�^���>���=|��4{����m9��՝�~9��ųs�;.������~7N�����[8oO���Ga0�JS �$V#�ߜ��G �������f_�3��*���އ�[L/KV3L�`��gG3zZ;'b�<LM��ܲ�tZ��M�#a����7�w�Cf)S�E�1X����L�@L���U@�շ����*��Wx1����Gܓ�M���HI#f.���Z�ŧz���FM����k,ݍg������c�5 �)�4�v�2!�۵/�,b"�l͋0;���؛�G<�2�;�iKtP�-%�U������:X(ǿ�Ŭ�E�����`�ٍ}�S6Yi�۹�a',�8=N��밆�c,�l6)��=	)&�UO>���������/���u���[I��+{LEWj�X) �
�^
�}3䳅�O=�|76Aw�҇R��|d��ޙ*��AT��oL핺��� l���&�XIFqda+�B���ȣ_J�b���;:�J���Xi��i�3WTWx�es��n�NO��I�Ƚ�;��nt���;*�Pڤ�m��!�!����|�*S0i�)w^l�p�u���x���(��#� ���V�}�ܻl
�5M��R|<:��U����f���U�&�v����X+u+h��)^V��.Y�����p�_�&R�:xk��6s̸ȵ�~�x6ʳ<N)����(+Y�H�ڊ��9�7�� 2}4� AM�/����
�c	d�'�i�ػ��&F�=�zk�/ھ���^�x@�5Ȃ��q���3n*aU��ٓ�-����ږ���o�v�Voj(4�|í�AOEѮ��U[����"",�h��tO����_>䀑�� ����L�A!�Y����d��L���$Da�Rl��u�3p�h+���(�%�Gc6�#h;������פ�d�CO)�e�	]L�n��w"��s[�Dƪ`G[�꓊w��U�\��&o$Vi�F&��fT*�"�҈�W�ѭ�����uI���V��g;b�V���L,��q�$�^<�.���^'�
�xP�X�{��֬^�C6�E&���l�}�����}&��4��'���|-8e]��
w�<���,.U{�u�($��[�1���d�"��J�����j�X�0'�x���A�����k��1�>�5�n-�ϲX2Çs{WsU�:�������cwM}(ǻqz�����,�ѐ�A�L6�8d����+�H��U�{X�.NJ2���S���/T�As�Y�OCiT�u�p9>Ş�䨙�[F1������SŠ-8�lS������%!�5�E[9���cש�
�X��VC6LΞ�!�Gtŝx�5� 閛C�I���r�[4`���y٤
��6������	>�A�?���1<��T��s[cP;>�����7���3{�L�gE��)��w@lщ�g���J*&�:�a]l�;�']�e���x��Z'J{��/mVL�r�O��#>k��m�#��泉b�{�G:�I;�{��j��'/�D�[YJk3�Ǘ�c��&l��$6X,ޅb)��v`�{z/�^Z�I���{/^�9�6zQ�z���9q�U���O9=�w��{��^��;Y����\��o���z>�zt����S g��9"�)Q��N�M���R�E<��8=�;�oXn�Ny�xU�����]U3Y��_d�������_4���0�-3A+d+9����ӓ|�+;L��9��̧ �!�p�u�h|�H�O)u����U	۞���<�ӣ�ɐL��B2�4G����7b�5~����"��Mu-E�`(Oe���{>DVY��F�%�B�O�h6`���m�t�I��h���:S�ꗸ{��7d�DO{���:����.5
n����33gdFh���7������V�nugKOFl$�b�d�Y���PfsN�v�,qa�a�4ivO��T�Y:�ts�Q5;����:;U�m>�Z��<��im2�,⁋�	�ª�m�7܈��;���[ s���/���`*U�b� ��Y�㷢�2�D���e[�^,&'!g�gFn�z䁔����r�d`����f_�4����~����eb��{�Rs���Y����}�^'Inx�.�	z���)�Sᐻ����u�Ơ{ɑ��֫tH������_K�yf�e#I�����4藯[T�����l�(���㝃�7��8!Y�o���.�V��{����w{ww7N��.c�zc{Ո �Q����7/�{��f�u�Ϙ�:+P��f??�s{2𝸹�m5z�U�H�ӳ��.1���U�m2����e��ݎSA﩮���؈zu�I^�tk�[FA0n�@�jN՛[^+2�;ղ�k���.{l_BG���ӛO��b�N٧���&�*J�Y7SK�Pk�j�WNFdȞzݝ����O�0�d�E�C��i}K���J*f�&��g��Zp��M�q��y�u!��?��p["�giv�(�L����b��q7����*���ޞ��x$��i����;٘u�7��ǆ�~2�$�/���(Vj�wۙ�=�ٲ_������V�G���D2�0�dD-��q��c.V�o�|"�vi3K,�ݢ�~�B[$rm�}��4��3E�v�zl��/2b,�&6/z��RSI����G��c�J�ށ�x9��U4*rYX됔R�6=���� ���l٘�Sƾ���e��"ֈ�f�	�^Q�n�ۦҸ���9{.���{5��|����܇^l�*��t��d"�۴ގ�����eA���T`�&99Kk�+*���8�(_>���<��:�%}x�B�_N����k�x�ضD��rscwR�On50<�c��W��x*`���屹0�t5z���ܦ7��=`3Y�nbi�:����^`��˔���^/u۽�傊�g��C��0;1�0��9]Ul,V��@ܚѝ�fKognR��
�!�K��EH6o���X6v==#�ę��|�b6@�/=܃��s+��٣�:�_S:��q`�F�®o��&��fp3O�@�F�rqP�d�A?$�HLT�����˺or� C�N�j�e�wAn�l�o(�"Ok���
�jV�\�Ur������ۙ�Eӻ�n�Oo�kP�@�SY^�O�n�L��1I���Uw�"�u��.ng]��:{{�ɪ�DΑG���l��lu.���r^ӈy�����]]�|M�z(����㻗L�	�䅵� =�3U���a�ە�-��n��i_�x ߺ�,�1��U������9A7:�fg[��#�$Ѣ�[�R�F���M�92��Q�n�ʬ������!���뛛n�O�H��[z�[�h^���;r6])�:���v�C�13�o���o[?\�<OPb�W��lr�]Y>��
��fC>�X�@���i�*7;�a�DJ�T��4�¢}ƻ���.\�Y亲_x���}�;�/.�F5���"�bu	��*s���4�P4������V� ����M!�IK�q���f����F����7ȫ"ַM�{��o�R~��9[�}����_}�xc)����m���Ð��t�Z��5�;sz�������mPg�*dw�@q�y�͈Ϡ+7�R����w	�t)]��͙�|�,w�f��4��C�p�<z6� )ځ2��g�V7XkrWRv�����A�����>����קA��
�T��z�ms�RM�����z��M�
AHE�,��T�{z��@׵�[�vM�f�Ԟ�<l�;��-6���i�Ô�r�	#%���<�� ʕ7\�V6�~$�f1x��edo	��D�c�M���`���AoB���O�򟅚��g�0�����ʜ�v���ϡV7q��Bҕ|]����t�a�yY<v�L�pcm1���ѝb׉�e�W/�x&�dY�p!yr���{]��-y.�#R�j�OTM�^�K&� �9�p��z����-�v��ٴ��{1�������E�L@��n���-�Y��ö묎�X�+�e�W���g���22�z��=�tf�XD55ԫ���5x�����{	H�����*��q�o���.n�Ӵ�륫el�w��3sReݬ�F�,�۾M^��0��0=���:����y+�	+���ح�;�y��{e�_�o\�0׼��K���WX}�Ss8����g<�L�R^u�?�F@6��C�ޖ����'���'åby���Wj8e]V-�lۋ�A�R0�m���/-��>􈂍'�ݜi�� `�ít��U�]pw=5[�����Y|���)��{�6���zb5n��cO�c�[��ݞ�Z׼S�����>����;� ��1��KǸZ�f��nǽ~��PU��g@+k�Z�o9�q�_�/RV��+tD�.�̒�!��m��p���m!VM����(�ȷpa�oi��V�fG!�/j_(�[2ژe�e^��t@�f�cPg���u�־*@l�b�ڛ"�6�R�E�\�ʋ#��&_1ƞ���O�R�KdGC�l68��ǚ�̓�,9�u����|�w2��Mj0�/{�,����>�="�"ť=���7Y|�{�W�u���PӸª���z�f���%��|��0(�p�]�^3�3��)�b,��à6��bN��{��h4�@Ͷ��Cj���5�1�LKٸ��F�s"+3Ud�usݍ�{��>�=	.=��=j�~�
6��|bF&�_ϻ*���Ug����ѷٮݙ5]��j��QKJW9�u��-�6Ż��7*�=n`>E�謬�
�l��i�vG��wJ��AmZ�=����Q�1��l�ʨ��������	�;F��*�Pxe�򬁡�8׉���F�9휏��íW+צ��4�]�=�0fw��f{"��r�A�s��Ժ[��|�wT1"�6�mR�؊ˢ�]4� r�t�6ϣ���P;�wg��ۢw8Z�iٍ�,2I[�e�f��R�õT��:��w^һKu�p>��7( �Ƈhy����!ۖ�vfDSn�O���V(�35��p8e͑bTU��#���]u�F�6��m�,f�gX�p�Wm!.�rba�w�W�H+�����7k��[{֨�t~�y��JڟZXn���VJK�s�;���q�k�i�&j�����J���n��Y�Hl�O9J4,�1[�n�����f�U�C�i��<UGt�]��%% :ƌ��%�d��q-,%֮�SK{����8�\�}X7pi�]��Z�f\���c/���KA[��j�y�|9D��Q�ZQ+-�G*�:��O#����h�oA��V�evǰUbZ�:�Ï�������c�b��;��\��m���{�Z�fd̺� ����(o:=�Jw����7l���奣w:��3����WW@@�R���*e:k��Ν�R� iX,%/ݲ9�UK��QT�[- 1��aІM�V���ިF]��]���G��9r�j�RKK���w.��[]���$��*s���n���*��ɓ8��zxF1�Y�x�ov͜��R�)a��fgJb�Fv$��Xy�Z��'.��;*kn
K�|Qb*���	���S�zw1an>Tp�z�=�{l���u,�,'�.�w�tun�`�x��t�U��Y���+͵-?�t���cXӛ�e�
�B�e>�d�f`�^&��eH��s&b��1@0�g&�i
�7�Q���/�VH�]�|�H1�ځ�]��l +p�H�7�U�*w�<J'G��Ver�[�yh��������*�U:�s���h�1���kU�ìm�����3+�+�!儈K>�Ҏ�y&�
���P�Ӝ�NPPt�vqug6V^B��gP���G���X�u�b价�c{b��J7��m'�y
����K�����Kn�u��HY�1�'3���*�'�Gg|k+�F(�r�Y����=�^���e-"�2�#��xc[x��a�ҭ�-)[Z��:�\��T��8�jlɺE��֚W��Z�5�r���]v<��-���.��4W��]	�7���*�ĥӁP&E'�gl�m�1�I��������-R����kZ�]d�if2E��Z��Q�"B�3��[[��i�S�����Yv�/�_����rM)3E$2��M�@�SO�pu�Ӻܟnn�:��a,��n-'����O�>m)�_fZȠޮ�x���CM(h5}�Ҹ^�>��9�.�N�oHV�(3RE�x��cӶQ� r;
ZТ�C�LT�uu�ԣ��.pw�R���G�tJ�ck.AՒgtˡԀZ��oS*� �-
w����d:���WT�Wc$e�|F���e���7kz*�^,�;{�j�]��+6��-�=ڷun��7�9�(���Ï6�lX\�H�L���C�C$�Q&�(��]X�b������&���\��C#T���p�J�Eu��M-+��*�w/�q*�����|�7�]�	�Va+4K_!�Dt�K�K�y����X��@�Z��CWws�U���|�7���)WM�*�+7��I+�!���iQ{���OoZy�y�Qݻ9Gև�S�w��2�HW�#�NQ�KSD�
>n���I
��C�(�0�i��\�u�0��ǣ���(���n�ET�w7�x�����=��z�E�fh�鋢Qz�*]�ݜ�$Lx��hs��'*�\�a��$��(�ݹ�<��������ӟ\�s����^HOz�ٻ���r#�x�"����y�n:�p���r�=���.�E��.�乑AqrC�*��'��U��;(+�p+֜�	E˪*EuNNVANHG�w����IЌʤ�B��'pJz���U��}{�tnDOݕ�z<���O!$�'$��רR��{����hp�DZ�ww����ZP}UudW��iO)K:TUD\"��\1f�`�   @;�a!��qwO^���ˢ���1�вA�1cC+��pZu�/��u� ogtk�Z�2�,�M��`u�uXi3�1$
�xf�q�P�B�#����Og$��aЛ0��\�2��~�L�k�pyQql���L4tn$��/A.R�w����Q��-�c8Y��:V�W.S����ck�]23�D���ƫ���QZ��d(���Lc��xmI^N)�)��+�;�ݦv2�(�S��; ^��ؾK+�u�ӝ�KOx0��1�ᓪ�V�t�nv�8Ӿ�>upy��/�s��k��nYd���Wn;fŞ#geZ����t�S��z�7wH�F`,230���#��oT����@��Q�G`C�I�c��Bm̅�pɜ:���U$DHFେ~���0�Ƕߟ��N\�a���K`*U��2��8�^ݘV�gJ)�Z�E��3f.V9��"'0�WF��=o&�W><�$lڤ�mkN^����`M��;W��q���ى�*}�{M�4PO b$ji�R)%�-��4��)[���/�l�5x8��'��|N�!�t"��N���F$3,H�i�Ҙ�����9�(jfn���n՗X ��n9lj�u;q��¼ƱǶ��U�Ħ-ɋ��X)��)�M��|�9c^Y��)���[t9���v���t0<}�1H�x2~,����I���]]]j[4��E���i�~nub�Z �K�u�e������ze�����B�7ky���/(&k4]ǲ�NO]q��ӻ�IU���(XәN�ņ�k�BBp|��2�5�X�*�7��ӷ]�3��{Iɬ�Kk��<�ږ̇)�D>[����%�bd��3�9��2��O�"PO+6�VB������w��8�Ǫ���<zv�����ۻoT�8}
��7�����>�(�N��F{k��9�n있x����6�ZLgl+Mdȇ]0x���1��ċ4�=�H�L���j.������t�܈����@�fqn��F(��2&��/����r+/ع�GMZn{me����զ��>��?}#8[l���c��ǟqt�\(���^^D�=�7{w�۳j:���-��Sҕ1���0�ch�S�rk�VhvH�x�-P�4��mc�פ��΅�Kl��N�u��#~����4i��l,��wy&�ٹlpvj^ԥ��J���+¹�׽	6�9�8g7M��3J���(��ڰ�w���Ni�i��vb�i��u8_�����yy]-��Ӥ34���)�Dt�)Χ7V�S�T?���~�ʇ�[�%�oi�h�/A����?�'��teӼR��g�W�r�tK�!
�2�Oq��c�Rdk�����0�zi���3�5�웚�ӶZ���e<Y9�o�jFah�[��C���#D8��/ZNsdG�~#�gH-S�S]j����N����Fmiw�,��I0��[b����Q�q������Iv������T�E0�GFTOXĖ���A��"X,�����}�#z��ҝ��=��j��n] ?KPEB���u���ͨ�F�gs��U�Y�9|����/����S��[N͒���wb�Z�!��3rb̲����~�=Ў_�������5�-4#�ƎJ�jn�r�^ٺՃx�
#�ٗ��s�P䌆0�2�lI./�l��[�ࢥ���໶~�
Sb����F��Wlz��]#�h�*�4�M�<E���l�ȅ���g,3;�~Gk>���A�ﵾ϶�N�C,�E2lK���\s�:�3ζ���Qi�}�g�W^)��z�"��T������U��5I&��ww_%��n�ա�����sp���V��@͡�0v��k/9G�	3=�~0O���'���n���]N^�o��](��� �����n��c��ܙwv+m�u��l�e�>s���ٍ�p	bw5�q�2�=AV�C���#����3�ue��P�������ofI��UJ�m�f՝�n#�gA��ү�me�����t���@��mM��bø��*�q����H����f8�iǱ�j�f`a��K"*���L���ǳw:�6b0o2���+4P������(/���O�3sE�U�}�@|���g;/��e���U�Վ�:�Ϙ�\�����☳M�[�fΜ���ٰ{��oRl�G�%�EwT$�D٪�ڛ775�M���M�a�3��,�m�l\*�Z�ݲ8��1{d�gR��P�R{��fU�����7J�nڵ��5B���/]����^S4�ਃ��s�6��:wtg��v��=۹עjʲ���� �@MZ�7Ftր��;n��y���Xe�b�j 3w��zg�����}C��O���LFcLuM���M�2��P�8h�lX7���I���i!R�ى7g�Y��oj1��w^
��gd��	����<���P��F���;��R�ܣ�s���	Aw�A�$���̛T�*�o:��4�S{�k�e���2����l�b)am~:	�����+�H�g��'�i����}��Y��) 9^D���F4s5G%���֌�ԶF�r-a���n6eݛU�s�3q;�d����/dW���w�S@~$V���f��6 ��D��c��n��:�{O�qޢ�qY]���xB.GOXg|���4aʋ8�=l�U��p�x��ΤvJ���|�U?h#��݀�L]6T��x��<p�L9���1t:���۔æY�y-�u]'>��*���K9̓="��r��L��z1z�vǏr�Dc���w%�α�SLq��EetZ�:�uk���kq#w�NU��A�%��]W(gf~ՖO_w3�ۧ�ky6�G{��GL�����[��|G����ծ���x�f^���5�},��+CS��w����7j�m0k59��8�W2]`+�f�N���ZΣ�'�v���Ï���~^�2��W���m�u4Z��R`��2G����-�̀���97%�q
Nb�C>�g7F���'�e�Lʾ��sD%��:��g�p8К uF@�}̵�t<)�VTK�^b͢�K�e���_�F�ql�HcL�l�ں
�yp��5Ѧyj��{ox�4-(�/�ŴFH<�
�k�:�p�:dlC;]�:�"�N��4��"�ȉ���8N'0+
衐�t�RNԙ4�
x��:����pe�^�W�}uQḖ_!ȋR�%�l���AS�d���/d~��K鰛���RO����	y�)��#�ay����\�<6)�[r�4�����ӧ�NW%,hl�X��MP�����Ʋ{y�s!���=�GRA:W���@��4���w@��a�ky� ���F����r�x�xp���x��$���l���(GR���Ȭ�wh$ߝbi�<�N6����T�(��h��)ޕ�ˤ��F䄍�P�jr^�VrJ�k��n�T�A�'$�x��b�=0���(hW��_
�J�S
cy}5���K�R�=�@s�Ѻ'[Vd�!�9>�w��9;�wVL�� r�:�n괶Y�Cz�N��Lu��h�F�Dt�1W��+���)���F^f^��VB`�a��g+a��˕h����T;4��H�����LK�5sQ=P�:�sj�mv?|
�t`p���6}zDBF��Un��Ȭ��;а�̺��<�sjJ�_O�m�3����i��.ܔŁ�0�)F�v�^+��h�W��}G����[��1���7��]��I�hti�(��_�p�W$bJA�M ���t���8bN��{������	Q�ۼ{�/��|���@��]h�q����yTO�X�!�7m�9��;Z�pnW���.��T��|pfz���8�1Z����F��'lk;FVn�5��HΗ�7�N�=�EP
n�n�w�/>�E�'�0�L���mU��#��A�r�ަli��͹�b�Cܙ����"������k:A�}g�����oLU�J��d댑ˆ����Z=)3U4[ ��6�x�q27}��7g�Q�׉�=���7JEj��4�����΋N�J7d^z9ر����/J.�^V6rU��+2��1K�65ʖ��bnE�r�Em��r����Rj�K]�x#f�����U���l|w��/�vrH߆t����ASS=vU��¨�2�m�9����]?v��w���C�����Ў|�����J�@F�ݱ�lue`�&�'��b�;�Yb�WA��
�"��<��@r��zJ�|�'1���幩}�ރ]:�=C�v��'���,�F�J��S"ZZakT���}���<n	6���dI:�K2�gś"ߣ�H�N�S7.�������|�����J8��j�	f~Y���Wi�RgGz�έ�����j�Ҭ��)c�j��#P��#L�ilS~�4�˚<���K1�y�fb: |�T;�-��]!���� ������.љu�0v�����4W(�Vǳ)*��{�����foM��sB�:.;���/��z�v\=M�.4/�g����Ų9����%�F��ʺ��k�����,d�
t�2���/"�
#�nKv� ��㏜}tm��8��{R�^�����e���S��$0Lô�0����X���v���05�l���_�Nlu,]��ZX�r=�fL��fi�[j�Kn�V�1�d�ɦSX��{R�Q �`X��N�̻��C���u�.��Nt$��DYSb�<�������.��:? ���{3E3�J���q��i�N�\�⺊���oG^�SD��ݍ͖���z^F��!�k�,�S)�l2�AZ���sy׼K�L�B5;yX�b� ^�%�����qH��\�[h�x����>덩.��rP&�s��PSJQ6��̦F뵮�{Z1sl�{n2��ϝse��xg#g��a����/:�kr�XS���f��{��3��ϴf�M�2Ց�u!�]�	s=����Qvs67�{{�D�w$�$��U{�V�jc��r��Y"�g��i]=7"ʚ|���}aSy����wgPכT8�O�7��=l�d|�(R�yώ��9�TC��-���[���,1�{*�[�s�*ߴ�6�g�~_���^̫��L�g&�u��Ҕc�It��K(�SuQy��0s�\�3���MW|������^����ƅ<�W��&q�p�B�Z�]i�C5�5j��B^G�*����-�}�*�I���4y�Z�4.»�6z�'Z߄A����Llm��sӣ�u>+ue�������O���uX�oj�i���(=�ޟ:%ߒ�3����]vx�&w����j*�4��םZI�~���/<�i�h�(�m�* �ӵ�س����E<�kM�&���sk�q���&��{\0�e�"1R\�fwe�/'*!�M��F�Q����[�9<��GPd����S�jNfU�`�y�k-����Z8�9�;V6��Z�)(1�S�ؤ<-����mu���wػ��.�d�{���3%�w�E�<�$�f�T�N�U�X��86�˱�'8�<dvUh�T��v����RC$��u{/nt\���|r���ɀ�J�]�#�od��Jd�[��H��T�Զ��G/�Y���5U��~���CF���&�'��*�[T�T���G�?	����>��֫�,����]��q��8Z�KN
��	DE�M�����6y"i���K�X�]cW\a:��fҴ�s���}�<.�+u��l�K
Y��/4�-�mbIgL�s&�>Ѹ�Ҹ!�n������]99E�V��/6��#/y!Z�t__#���J��'��/�,ٳF5R��5�ޛ�ؖ�S4�=h�^е�S��yTU�nTV�wFi5\)�ӻ�L�֗����j�I��\��dX:��E�#M���әB�L�h;��������p���KJL��A��m�]��r�x��٫�*�J��J���{�2��-_$M.���������u��z�fzwp���suQ��sVl4����mu��\ܶ5oW>M!S�2����V�9��[1;t]�!B���;Q\�.�"*;�*�o��C��D�en�[��ꬰr�];X�>MańGG8�$�� ��Yz�Ҕ=P�[�u�0�hWV&Ne<	��ԫ��X��&I�����M�](im��*)��wv����J��I3k"��MPr�M�|�J��X��%�3_m�봈n�b�tU�iq�����6y��ҢYbYݬ>�9U�+��]��~�G�����A�����f�U��/4�ǀf��t��-F�Qՙ'O5:��� ���bvY���hRG��k�B��B��w\X/�`��g��M�Sj�1�J(Gx��6˺V��ɶ�SJ
űC`��\�φ��V����L��Б8�1�L�T��VWh������a���i�!+k'�g�Ӂ��H��7��Vk<��Wd�v�ֺ�S��,r��s{nb.��9K�Z>�l�ƵCw���n���N�rݩ�q�2)Y�t�v���#�l�3��E�2��`T��eS}����2��%�}�7R��������rV�J�5ʃm�צ�䮁��E�L�F\���}AWfS�J�7AsLQ��N�9�ԋv)���Y���#v��q�ܹ�gS��4�T�V��O��J��Ӧfl��R���'
H�Š՗����7��X���Z��K����S7ej�rg&U흹�hm�巛����菥�T�\�X�f�^v�6�y�dVc�ôNE�)������|;B�H��F�I�$��匔fn�ݶ.��ȫm�(���%��Hk�2�ZMd�KJ�<����A�MW&�b�lO��h
���`��{w�w�aQ�l�O+�F��N�wy@9�VTN��kzv��&֚�"PR5ۛ�ϲQ�1�U�����]v�}͘���+S5�Ǭ��gdu� Y�/[�2�������vT\Z<�:��d��S�Դ�tƺC�k�\�mh
`���Wt������k���4ήP K�<�}B�'VШ�EFmlN�������V쨹�6��	�H^���1,ѷ:�r�T���t��B+��A��gq��en)l�W^���:�Pڸ���M�g9�4;�D\9/�
9v��PNi������G���9�Y�sD�;�t[��~����!����(�Ȩ�\�Eȸ�Gp��Gh�_wp�f	(�G)P�	�v�n�7��|�h�O���Ep�b�I����+����A;�ȹ�Ioj�EU_SD�׺D}s'f��*rNABe�ǘ�&�J"����./���w8��3�Q�����z������Ҝ.�Гz<�<�#�k���!OP�\z�i<'qruy���Ԫ �P�y����͔|ʢ�oqq��.p�B1����s�
�\���Az!D_QE�*��%zI�w(�|Ȃ�r�*4""ג��!�P�"������h\�GG�:��;����M�=y�صc�� ��*�����YE��bDV�ya��q��(ԺX�H��z!�z�P�����Ⱦ��;9�z:�(����gE�IDIE�!	�<�0�9Y��rB��GL-�� �u绮A���ve�n;v/3u�:݃�c&[�Ҿ��^��Z�K�f}�%����h9ջ�^�j��&���PQag]�lf�f�!Wn�w��G�駬gӲU�W�X�[-���ܦnLE�U��e��4�ei����CH;�O�,aIn��>�J=���;�>l�ٝvO7����gnM
�wd�`[6��o�՞]^�U�afW�[�N��>�}qmB��a�M�rs�"�_կ�VVe*�u���C�q�]"�tn'�aڠT4��ʃF3E��d��d�Ð�}�JxvF�p�]OCn�ٌ��*����l��*Ȗ���X�1�g`����{��|ݗ��E�_�s�i0���״���ۢo������ >m�\���)�k6��ט��S3ڻ~�7��g���������w��r��]���ro�ݸ�=���$�L������v�%�{	�4e(��P�6�Ou�@��ʣ|cg�!�<z-��
G=�{�7��JUߟ�3<�q�����SI6Y4-D�d:m^�%��tv%<Y®:4]c���)Rk��qJ꬇R��0�G��������2G��]�,d�[�^v��43w�����YgaŔ��T��ȣ���ɱ��v��/)u��N��VBkhZ�$������z�r�����.G�o���0�o� �J�9��p��BJ`'rw~;#\z�� fS�ա�E���K�5g+v�z�E�e^�L�hL���;-t�B��Q߀8po'���lѪ�5�rR٧�C!�g>�m25"���;fMݤJٵ(��dr��mU{���A��7.�B�䈚�TV��:2j�8�n�h	�g�H�R��^���1��t�V�R�ƶ�V�d9m8��˘�"�>��^&��~(򵵒)U�[�&�]�u6�f���v��s��v%�H�OŲ`��Y|Z�_$l3�>�'����ϖ��ټkx�@��K�᭞��ig%���u-K�{u����P�KD�����v#_3y���{��6�a���=,��d���d�N��OG��x�~��s���Fî���|u��׌ !�7Ea6��hS�ܺ�X�w�K��y���~�z��1��u­wV�M�lk�ALj�^ҹi郺� 0�=�z:l�ƶ�s�X���Ħ�]͎|EEw�a�Q�Q�(�Jޑ�o���L�W�]\����ﱘ%��3�7��b�����Z��u�P� �{����|�9p��*�ĥ�K��W��2��57Q��h`ֶ#�_'v���0��w�!��(w�f7{���k+܋\�ӛ���^!��ŉhٗB�q�{\���`�9>�X�PVkj����XPsݐcA�v�ôݶ�<���M�|h&_lϠ+6/�ų�~�=b�������W��=����AoQ����V�q:���QMQ�8�NЕ��w�Sl�z���k��q���m�����	݆u������F�#!�!9��x�$s��Nd�x�-�����W����1�u�a�޻#ww!�ii�>��>s}@iS>�@��RҪ.���9o �~3�=z�[ ���y��^箙7f��m�
 �h�[�9��,t"���jz�h8��f���
ιM|,�R�~�<h䥳��MQ����C�1��:��!Q���=��YN���5'���7��u˗�����Z�ɛ��?��<vk���>t.ϲ��nD�n+..yRun�q[��EIw7o�!]�vs�7��Y�Ӹ�V���K��>=|wrf#�X�@L�u7(�+�h9�e�YT��z��OL��{�k�U�Q���K3�z��X��wW͸�O�P՝�H������.-����6g��s��Ǚ_ 1���#[#v��6�I�1����V�-l[��+5�����{��[&oc����G�Zh���{|.��m���.V���^�;��v��/6h�y�漡�n���>K�ץ�;��c`m����+�tV�����ͽG���Z����c�4Zk�C�]�}K�����䫫|�5x�.�o�͖��;�5n���c4H}���v�4O�\v���	�N�oB}�~|�6+6�f�v읎�ګW�6A��#�7H>�-�wO��	��әYq7/ګ{l��>��'�u7��؃�$���@�`�^�1k,8#��5UB��{�|'�����س�^G�[d���� q��|i��wMxǈ�O-X��4��&�5~�u=]ʮ�ui'҅kJ�Y������b�|����������Ί�i��t�in5o����j�(WnbƖ���}{�6���Ӎl}����s��&���'�$��zU�c��Su2ƾ���Ê��c��:ι����"u��0+v��=9�/>�-p�:��*�\gb�$<<K�̓��6�c��J��^.Mm��%F��v�Hg��Ձ���Λ݇��=��
v�ڂUK U5t���s^�S�c)tM�3�M�vsu�����%=��ej��.��FC]��q�"�Y���C$]R�8�����7^$��2v�qV�*�J���N��`(���̕�}�M���6C���S�#Lc<������/(Z���Ǔ�XklJ�䪛�|l��܃岑-�Y|(n���䒿'��`��]Y�y��s��pe^1:��{r�+��!��
 ��n�Y��\l�Z���ρ>ò*�x���:ݙQ�3������s�>��n66Ү�c�US=��i{��#r"owe��\�I'��E�M����a�e��R7����m�dktŹV$E�yٔ�
��h[3�w�������7i��)�M*�Y�֬�a���|z21a���B��'Ƿ��v������|�b�J��>Ѱ.�y��v���3&�ݩ�)k��D��aEӟ�f���*��Ls�����={׿����\�}Kv�i.0�"�dw��͂�m�X-Zn�!�7���F�uY5rS���,��E��u�*c�՞q��Щ�$� l�V�3OS��E�=M��q�q�[��"�Oh��i�i�pĜ/Aͨ��W�T]��>�3'~�F:��?��^b�pU�љ��@��NSH*��쎜�/v�����l��R���3�����Yx�Y��]�}�-���S��t�g6'D��;dW����mL�Mfґ]U��Z��#�g���fm�"*�t�m��{fs�ߵGb�@�'�{m��k�����^eOsWN[vҞ�k�~§�b�)d�UMױZ�V���&i��E��4Lemw6讹r���P�4�s!_)mZ��,��U]P9��.)����|�൞�cQ{��F�F	K)d��C�3�ۥuf�]��g��M���JF�cBzu� ����W�%[9gO�v�0X�kz�W����+4�N4�x��f�32���*q.�4�شt;V���ޔ�d���Q�ᷕ����{�����:�>R�q�Ys��1��*�gt�o ���H�:O����u��1^5�[0E�ث�|�8ES&�&��U�� 6d��>��ȿng��](�r��r�6�e-�Y4t�����駆ח&F��Yd���.1�!����ý���y������w$"q:�,dd�J�|Y���x��ӹ��{��8C�=�/9�^8�w�:��(��d�ٞ[�_u��]Uyxi�^O���%��M�I�J�2�՗�ΡM�Cs3Uj��=�s�.z����z�#������Fl��|���Q\�4���v&�˚i�ͪz���eS��bs�$�)6�nSm�ݔw��L9�lt�0n`,�7#{CI���Uw��=���d@Vg�/�n-�������M�:���j�x�|�ǰH*��4=����a�x��b�;a�C\{I`�c��/��wy([!�J��#L�a��p�;�4�ж]�'w:+F\k�A�^�؛�,��:t����nv���q���؈�K3� ��c��hWyLܳ]�-��c�\x��OӞE	H�l����l8�K1��𼈣pWi,��9�\���[|��B�i�n>\�j�+��<%����¯8��t��K��B^c�R�Y�;yi����$uS����f"b�CQj����ǩ����)�|�6� \m�X�cC�s[q�]�Q]��Q�@���v���j���: jwv������G=�9-J^���Tz�\�SD�=
�@��Aʫxg�t�g)�nr���#nb��n;���U 7RʎM�-<R�iw=|a�S�6Z���jj~3�@�܂j��٬�Y�S�HV�â�m�T���P��w��C�q�%YT���U��+d	��8�K=Ô��t�?sa%N��.���Z�������X]�ˍ�GV�	+�yԆ�.ê�2�r��2q�/C��9����nr��J�Adi�|��}�}���1�w��3X��*��=�r�~͘}�m⪵�>�:�Wu�I�n�S��f��2�M�M� q�"x!_��p��?��:y+< ����٨g%��C��o��m���5nX\�tm�j�t� 
ܨ����$����;����v����T��W�V��X�њY�HLU�Q��Yw�<�� [܍s�Tnf`C��۪��R`81�`su҃��)rq�8>�̹���qS�����g
&�tP��1f��R>��~޽������×C�tUʆ!��0����\���8H~�V��H����:� ����O��5�d��MjN��-U9�׽Y�\��MB����n�-P�P�qW�^T9����r5���t��J����b���)V1ݻ#N6Ϲ�<Z�P�t�Y|�jDm����g�s4�%'��6c��<�\l��̗��H�Qy�lqd!fjڢ�c�x���=07�����-J�/����Xs�(3ZP.vZ��c�qX�WN�h���9��=����n��:6��O��'�ֿ�jP߭^h��W�}�F�����W8UFzջƠ�S��v�-C��T�A��]�u��z
����2n�.ɣ<h�*�p�<�X�lVn����U�ʱ�A�~��>Un+��:ur'�Y@j;���Ud�E�\e�4pg�}\�/*�s(�W�-[X+�=[CX����Yf�^^jb
�:Q*�"܎���A���&*�S;���+�O�B��}}OB1��2�vŐ�̝�:lN}�WZ��D@-P�C'_\��Ly�:���d�C5w�ú�?O�m���۞�6+���%e��ߊ�l��^8����İ��b{'_�G&W���~��`�ٸQ�}>��η���n�.�=��t�k97ef�B� �x�ݮ�gX��oE>e%�e� �/7.�0ۼU�ѵ]'�N��w���	l����a�fȅ�" �]_.�)�,'^Y�6x�q��J�\��ˠz�p�m��7@�7�Q�j�Ø}�'��ͭ��е*;ԧ�#��{�e�ya�E��u������dRj2a&R�r�d���ԅHj��n��I%^=Ō��NSn�u�5p���\@>,������oZ�W�]KhW@h�q^�6�4�;�}�5n�	���&a�`w����:�����Y}��p���.�:�������r�3�����ͻZ���c��,ca���?7|�~\wϟ> �������7��q�c�cm݀��w�q�;m�چ_���};��&�ɱ�L�0	��2l`�`�@�.q�3�0&q���1�g��}�Ý��;l ��� L�o;`�˝�3� �ۜ� +k ���m��� w��ڭ�&�p�m�d�m�;m�L�m�����l�� &v�l�  L�m�gm�ɓ&v�l��m�gm�&�l�� !��3� L�m�d6�&L 	�4  �6�d�m�L�m�d 3������l��m�gm�ɝ��!�m�L�m�gm�ɓm�L��3� &Cm�d�m�!�2!��ɍ�L�g`?����C��B>?��� lLm� �� 8���_��/���������g����������������a����ӊ���|�������lm��?�����ױ��m����cl����o��C8���;���6���6���A����{݄����}��o��������83~�m��m�c ��0CM�`�&� ��c&0`M�0	��!��3��g	�� �m��m�q�����cm�ˍ��m�ˍ�˃m�& 8�bpc��p�7������ ���P�v��������w�
�����o��}�����n���=���;���?�����̟���x�m�`��o�~������~��8��cm����o����o��6��6�����lm�����b�{Ѹ��/�}c�7N��������6����w�6m���������~����~���}������������1��6�?`������6ߨ��~�0x��o���`�c�`�����o}�������������6�X��s��c�b� ���C���m�-����m����6߱�����^���6����;��}o��p��b��L���M���-� � ���fO� Ēw|�U)AT
%
T�D�)�T�QU*Q
%F!I$�Q�Qk!T���)$*)%*�J��@"T$��ʙ
�I2�Vzn�VY%[jE*F�h֨Z�[0U,�i�l�ɖ�j�Aj�V��Va�1��a*��l��ME��f�j\�m����o\�f�mZV�X�E�L�cSE��Z���(V�e6Y�mh�
�j��eh��2ml�%L�,�Cf�QM4)R"�J��,�m�յ��Ѳ��-m��  ݷ���[
����Ze�&AZ��q֕�gN�l�Y��n�A@��շ[e��#q��VL��S�p�: m!�6�J�[Ut�m��j(�Kh�j��QW�  �ox����B�
��)BD�
=�C�;�}�С�=�"D�
��B�����b�[ͮ� 5[wi֕�Û���[mP`��b�-]nm�m���I�m�in�*�mh�K%��E���  ���(U���(��]�l֛`mu˱M[��6j�lm�����U�kQ�� :�U���P#w7f�AT��e�F�>�����ʲm�l�fQc+o�  �zPP�:��8�Z�ڔ��sF��Ҧ����24�(U�Z
���[
 �]�N�6�⨩ጠ
��0U�MM�kL��%%2I�͛W�  nǢRCw(N����t�]S" :�\��.�Z)��#Wq�(WV���P��gN%U@�)�M57;�6�fd٭�]�  ����]��B�*�a�P#-�TB&�PM�0h]`-+���HU�5�+k]ܡ@���U@�pd+ Z-wk�����-h�  �z�(�k U]:�*3�QE�U-���(\���QU�v�EUD��]B���s|I)V���UJ�)�H��m��M�ڬU�l�M��   �>�|T�/�N�)J��s�u �S���מ�P���b�*������wc�+{��*J�V��&�8	猡ґQyq�t��A����l���ض����   ;�}JR�T>�x{j\�{�B��t^+����T⺠�F��UURUOz��J��ԕ�W:))T*��w�%W�w5W8��B]ש��ք4il�l3aZ��   g^�DR�כ�*�Ku.�*����(^�� ���Qםꠗ`kW��Z*���y��օ�T���DGlPμ���*�� "y�%Q� hb)�IITi A�~�����)����~%*��  )�̪�i�42I��&*�  3S�~߷����-����r9�����`��g��K(����j�K, ���__�������j�}����cm��cm����6��66m����1�p6�����?���|����5iF���ʋ ͉*��� e���:׉�@���2��Զ�#N�ÈBZŀ9�Z��p��7�n��WM4��͠���Dȭb�C-ԁ��J��J�p�� b��5hf(i�oB7i�m��̬6������[G)�zj'�FK��l�&�G~f��
8�њX�7Saݖ�'Gjt���4v�єM<[B�:^"�h$�����������5������S�TEn��#���J�J,%�Ӳ�b�2f'R�ݦ(�;w�fa���Ha��4�t��b]4�dw/Y,��Z�^h�pIi�#4ˇL��cs]n(� O�J3��K$qa3A�,�Rj',�������� ZM�9�S���P_Pj���(�i��v��:�Y��.H(Mbe��]�!b�eER,8,�t�,uຼ"��Z��,[��hF�:��9;̌�g4��<����up�2]]�Y{cv�"�7,�ʍ�y��M�Ѝ��mɏt�@k�Y$VQ,�0cW>Vi����t�e�;�҉=!�s;��˦�v�fޤ����9u����ٶ&�v���qZ2޽-�b�jS�p�NCT�+�KC4VQw��ʦK6e��ܛ)7ӗi#�*�y��{6ͬ���cq֝&h(���]&�Eҗ�Ei��5)YN�/N���I�'�,]�F9V!���8��3�R�"�k�[�7sS,�)�A�u���+^V4f1kIE8��b��5��8Ӡ���x���rf�UЅe��m"^42��P�T��[�����)kk)m���r��^A���ȳz]5���,Q[�Z�Yb�,7-��#E���x�/(Bn�ĭZz�f�A���0�0	��or��Xb���m,Y����(!0lPcA����D	/@���%B�f�ٕ}���@0	$���I�nT���+͊@���bbk/d��Y�
�y�z�%2�L�d@b	G��6��RU�W���EGe��A��Zljn�x/+"[o��K	Jh�hn��l�Y�'�!��oRRjF�6�u��������V�f�"��^-ִ��b�9�,�n7+Sv�.Q�w�wބ��41!	P��d"f�ߙ���C9eMG�:��8U<�,��DI�U�u�60e��m<u�N����(lK�bv�òk�I�ú��D��f�=��b=��sAgVmiR��pU��bU�Y��R-�Gn�O^2w#q�c�P�Iy��[�m⬻;��ONTrT�4�v�f��9P�2X{N^A���,%� �n��	<��;I�Z��	=Lh(T9��VZ�U��d�e/�����Y��P�[��)�n�`�ܘ�CU����MF�$:b�r�M��:�j��+�fV�U�0�r5R:0�1�&
��3Q��e]�v�gǖ��P"�T)���;�0�J�X�:z������6�	y vM]e�v)�{�KK{B��%��Ɨ\�H��k����IW��<�^�LhSʙA��!�S{�Ӭ�ǥ�{�*��;�!U��O5Y��	���mǶ$m�&�]���Z�D�3U�2��k����c.D�x�0��˦��Z4�'W�X%e��ΐ�D�2^`�s8N�������J���z7�1�ILR�P��]��Y��S��B��	�$�-���A9��t&%ˎ���v�M�yF9��mn	i=��X�TP
hRGm��˟aں���f�¶�H�1ٺ��Ñ�i�Uf/����b��أ6Q�^�l��e,�0�x)	R�-�(�R(B��cNk�wQn;�Fem+O3�iǔ(L�02�+e�;�5"�#�..˩D�Ձx����B���gۺD�۬7D�H��)[�`jh(��R��[����0S
/�c&��X�ˎ千>qV��޽U4�HR����J�KJ�U�[�u���iӳ5ۼ����-'whM��`���C���jUbE,�zd�W{���I4�SaG��V��v�O���DՏDw��&��R�[���4V��{Ad����i�0!�b-���T3hL%��VЋpl��!h��f[��,�e��q��F��`l!7M���+�i7{	Z��؞��U�����6�8�'Aȝ�չb���+2u��l�軨T�0�ݹ
i~�
�R_ 7P��6�%�ő��D�`��)T�=G2}3M�J!e�RRYsi�� 0�G �VZ�ܬ�Ri����dx�ц3 ���v�w`З��a�jLУ�)*��â�^13sD�VMH�nT����(���:��&�5.e������dhi�(M�F�%�1[K�KFV^e�n!�c����1�S.����&3��;��1�@e�(��y-��Wu	h�F�^CL-O3楋)h[d�W����Wۇ��ǟ]�޽T��ɸQ�7U:	]C1%��r��Cu(�������p�T.�=Gn�͸�M7���֛V��9Xɶ�.�\Y�[���F�S�n2�P!ӨB�V�fm눝 ^�?���t��Z�qP�Ï�$��C�B����^=w�OV!�;F�P�i� ���r�2Ux&�Z�]�щLD���P[�%�[�{�� YT(MqI�u�T�u{���"�!;w-9�Z�������	��h�!YCVnG.���u��Uh=A�Z�;��/!�i�ow-�4%�*�%�Jʫ�$
p&�����[��:hwNBEnP$��oD�����
��Mf�(�vز�[2�L�ֳ��ֶ?�E7\�VK	�ed��y�n�{c7�嚷4n�����h[����eĞr��跪� )ǛdPw�YFX{P\�;�i��酠�0j�D�7k
��5ǐ*�{�� n�v���rb`#�ۧ_bKSfj��J���s^�� -��R/���s��Ms�i>�� �B�S�/.Br
�S���6�n*`VB�Zvʤm�n�8P�c,d��T�쳻��[���n�#[�+i^%����Ne�Ob��c�����®��F��� ���F�!2��X�Ȓq����b�ˤ�ɄAy��ˍcX]&�YZqLl�i��	M�Q�&��21��Ѻ��q��fk��1�	eV��`��{-]�fbm�;�˥�A#F�n���e�Ge������:�~�=̼�X�k(^	�H�B��|䥣Y{�v�:n�[���hܒI�3�6�ۘ���aL�6��M�V��3D
y��V�`��-��ʎcVjk��֭ʱ�H��e�J0��e0�b�4Z��h���������tq#X�p�Xv$
����e��PX�è�)�KcyVj�兒�q�;s��hl�yyf�"���l�ٮ��*��oql��cd9i˧P��sY(Cul%H3@ĭ=Ȭ��A �V��	��lXe&U��F�f�-��:m�Q�+��f�P���RT��pJ&���iC&S�&Z�m��F+oX��u#yW��V�6W;����ӿ�5�32�+� �n��2�t��wM،�߷r|Զp���`Y�W�IZ��6�J�zp%���S�d@��|d�2�f�Z�I�*ɣo D��J��!�#Wu�j�E�,Y6"��P�e�C`gn�.�7�5�VK�
�Ƶl�t�6�+�ي�EMbZ���`t�l?@4�1���

�X���V����&O��ur�����jὮH����Ռ�q�N�5��J�O,�,X��-�5,��
�ITwwLk,j��8�o�pYRu���@٫׹a`��*Q}����Jzm"^�򴏖����#�1%n�[�*0T��5����z]
H�F�{W������#�E
��]��&�V'1��-�W�شsF�]�6(�
�S�0ާ�-Xܫ4�D�Ȳ2����vҽߵȍ �D��f�b�R�sU��-'oP�l�Sw�6��aU���u�����$�
ʸ��]&na�W�zB�1�ߎ jM�d���"ƍ��h;Z�Ec]6@��S1�7!jT6sCI��r�dҁZ��Q�֝bM����s	Y�֚vDJDPʂ�&���B�y���g"Wq�ܴ��y�6&i�x��5�9*�6���d�+&��#�����@5!L�p���,V戩�z�*�����=��ҡ��I������:0g��ެh٧���̡�U�]3X�"D�;yy�ڭQX.`ƨi- �ܢf���#�I�N�1i�y�5�٩��P,�fnR�oh��%��G�d8���t-�x��D�*�LF�P	��IN�e��ua.�����$�n�q�B=��f�U�פ��
��;,,n9��*�*�FGr�rn�t�+*HT����Hn]=�EA��$�,n��M�*�xul�r���/#����0�)�/)��eۼ_em�������C�p�h%p�Џ�5΁{%�n��`��N�)��1�V�t7[Y�W�<z�fk�E3��b�^��v�5&
/`+.���h,ӏu�h�ѧ�7V��08��fJu#���Vd�WsiիLd�"E5P��j�VRm8.KiT��v��5�v�+tn}v)���v�J�n�:���Fݤ�s75j��l����`�e�$�K0�4�c4*�����YX\Š�_F�h_k�|Q�B,Ix�t���<QҎ�B�D諱u�M��|�Q;,{u3)�F��
u�2���3X��X�H,M���3sc8�{��x��,�M]L�-_�����c74B,ޭmel�D�������d����i2bf8n)SbYtq�t$�^�ֳYV2��ѥ�!rí�0�Kw���To*bgMiU�ܵ���:ԬD&i�,�7w�അ+[E�q�MJU�WgP�w��iV�}�~�[�g��XS+ÃI�Pm:W�����)�A�eS{Z�Ro6�I|-a��t*�ZrĎ�`�S@�ކYC[$V���(��[������WQ�;B�ZU�v6+�uS�� a%�W�1n���;1�C/+TZ�iH����U���	u�ї���Z�	������#E֣�U��s����#mY���Ci��ьLpԢ+m)y�^Ȯɚj�#�f�H^-�)ꪟL�W�ʅ�Z�"+oD'�(E�7�U�cI-������w��[����a4�fhݺ�3�Ag�bP{����g]�
��t!�ŧ�Me(<"����,�؉��l��ޭ�H�zŉ
��n�e�j�V�N��j�	�F����X�h1���^!��*򌂎�T�;v�Q�w�QL��i�ˇhfKAn[SYV��R�����9Q��4X�f��SQ*�Ct�T�ASج���f�6��aV:�m,={�p��Z¬HGr�Q�B��1�؇"vh��|� �
�&O�a����[2�^H��f�Zr��!W4�V��gͬ���Ӻ.�d�H�7*�EP9��v]i��c����S�3*�6ZԎ,.��*Q�n7�y�a_^-j�G^�	o�j7���3^n��V' $i!X���eLR]57$�*,�up9�9{A��������#1��u��R�[@�72�:�xՁF��7W�G��Ke�mKB���743z�����P�ʭ�XXց�XD�]j+w(�
�Ä�t�)�Һm}9QC,W��`4չY�
�AQ*�4�%�ܬ��u���;��u76�GOn��{B��h��F�ތ8��g�w�6B��q:�i���{�>����9Q�Af���{%���]_�k�N��B��V���\[���c�)�ۘ%��Xt6��du���(�U#��b)6���6
�P��8��v���6��V�:&��������I�&�6;�աH1NV��E�	{
×�d�ֆ0�wMgv��v�V��� ��3^F� ���&�GZ.����5Z��ը,\�
���*�-VW�j&@V��L�,[���+rɋ"�ŕ��b��r�k��8�Qk�6�&3�J��7l�M�A��՘�6�Ds9��	�H�IfR�K�ѽP�F�V�+��u���na��!�EBj�J�'\��#�Z�F
"R԰9Pdc��tc0��n���1��)��qS�)�m�rR��iݱOs&^���r U���)�@F��{���-�����R��`�@o%��^��C���鎈Z!u)α�Vлn'�[�+Z�1ls%[���3ƒ�&i2QDD��J�@3h�k,fl�ye�PU�f��[�		�Hyu$��v�= �7"��)�7I9MY$�#-��Sl�[(R�kc��$���\@�����!&��iF�VKݛZ�%6GMdXg�@+R�'��$�9t��7�	2N�@�d��O�a�׍�;��������m���%�ǈ	V������G� ��Wj�QN���x�ī*��ɋ	�S��v�W�y���PE�m��[.7z��[����&�b��X͊#�?GG��r�4�1��s��t6�J=n���cx�Vj����z%d�j�T�Z��Wd
e@gdW`_�1вYi4�s����3;KQ��.����LR�z�K�B�%L�&��2��@��3�3$
��M��y�V���n�Y���N�W"�t���b�M���&��\��l��p+e�pTd�ʋ��c��z�vq��%#F�Z���ڼT��aR���*Ω�IzK:ۿ���k3n��E�Y�E�K�)2�qH�-�M��a�48����f��q���ż9��% s�O�!�b��ѥnO�����4,l�m��R�5#O(�C��@F9x݇�zm��d��A���G�3�����C���c�c����}����o�9봹١L^^V�Ԏ��Im�ٙ[dخ�Ywz/�dR���:o�U,��=%����;x�*�%��0�W��a�T&l�g��PVt�}ckm�j��uq��է�o)�t�dǆo9�\���LO����YC�^vKE;����"뭈yuu���U�����x���j2�mX��`�� ��`y.��#Z8t�}�3wp/H����mNo��I�{��{Q�y�l�]%�@��o��Cf�[���n�K��!��yy9���|����=���A�ft^g7�q�}�|�W7Z�s������qէ�p*�u7�Q���5����Ù�1>��)��<�Ev7H���S�y�6��yKr�R�l��r�'W��%����SzVy,�FuÆ��(�|7�pƇOL�/0\Jk{1޷�pR�,7������EI�
K��*V�M��� ���<�ɲ�Fj��t�"M��D.S������q�=�ίDN��:�d!���e�}Pg9N_��?���'����ﰿU���n"���n�ꨯ4�G�"=;2�3d�6��;`鴷��e�%�{�yj��>� I��p?�#���[W����J`=\���(�[۶�[VV�Ĉ�9�m^�n2�Ga�Ʈ�ڻ�����`���@���C)�]��7��=���Wղ��|:$�˱�:�co������{oMmHo����-yGa���2����佌T�^=�p_M^��;D=�٢��9����Z�%���s;�ωL�U�`���)�m�
��d��$�>VF4�k�$�Ic�Wb&���t7��j�� ��t�Z��-Wrw�Ģg�\"�5�3�U��NZ��j�^�����R{R�s2�j�NU����vp~� o����`�&�{�`К=��VD�:\	-6����3r,���w���g�wU_a}h/uU�n��wC*3���"^��ZSO�9��U�f�:�>}}	�)�䒲:�!�*Ų�)�طP#E�P�κ��y�Am�����xD¸���pǨ.�H���dde%>9Y
�̪�=qM�C����_�A��,�p��+�sv]A0g���ga�>��w
l�9�l����z���v�_����О��!���72�&���1��9���MQ����Z�>��;���nJh����h	����W� �Z�v�֊�Վ���J�̗;6�ަeq�[K6��	�aT���_����L�4h4�@��Z�7��k5�;�*ĥ�(�6.�����2`l}2�vr�����h���ܻB�0�m�����<���xշːy�s�/�ά<wOM��$�n��i��P�_;5���ЎP4�{n@���. U���s��T����2��[S��aK33u��Ԉ�n���L�<�a��p,�b>��ُ�5�V����N���� b�np��n�V2y��:�D��	y��[{�tu�w02��Q+9�'R[b����8���|c�BHG�7ܱ�Ljt��yW�U<�:C�4��5��}��I�a�<wD	��h���h�c��L�ʳn�!�6w��9}�W��+��pc��u�q�䭶̊\ Yt�#&��6�f\�ėc��&멽�p֤��$��8��g	��0��Ŗ%��S�  7Ɍ�Ӝ:���=SM�|5&E��Mp5��f��;����]�ͻ�Z%c���f�y���u-aӳ/4�ť���՞\yn��`��D;@9r�80<ַ5��9��ʝ��ݧx�=�GM�5��o��*%`� �n\��Aay^ �Y�d��Xo�{��ހՁ��9or�˩���b���iw��f`�;!�NҊ�Vs���Pv#��ItD��Z�����G
���v:V�cv:ܗH9�*ӻgH`��O� ��t���v���q8�s3J�͚�mC���\[�۶J�p�#�������D��VQJ".��hFu��s\�d���܂n�H�V);k�h�c-�6�b�ۙ��p~h�Fn��28����Y��+d4�h�w
��h(�ձ2���q�!E�%����V�u*v��M�ȶQj�ۈWs�!�����'���ּF��]�21�[4(��י�̲##VӷsYL.쳵�{p�ػqn�,����;���ޠG�����k�D��K��ֳ� O��ɋ��j^��ކ�}Ʋ�?*�ݝ�\����}9:���!A��c��j�r5|P)�_�'LҬ�u� ��v��#mb�8�!�(�]�:\���D�ŵl3�[{i5�tn�E�f%
B���s��s2[�88�n�Ѭ6�m�hE���3n���)
�1�|���L�4Y�/�-sI>����_XA<�ˆ���f�x�z;��p�Z�&�D)����H�Jo�u��������Y�:�zȨ37�^�V׽Yr��g�P������U:��3o{7W6���.�D�Ǹ][�*CA�g]+/"jd�KT������B�f�n��B�Tb_C��"v�BQ�}f�q�T;��c�욉�2{/	/Cܖ+6�)��o�%�f�8�Ԣ�1���i��TIq��I�}�,��@l�4�;��o���c�r�V�ƛ��z�9��c|�=N���P����� $��h+�#3G���d��x۹��f���Ғ�K����&fjoF�\�G�{ D�aK�j�V��y�@������L�b7���T�S�8� �9K47&�U�Af��� '6�AN�]F��6ݎ�ɝ���GaR�i����S0 ��0R1�Yʐ�VqA=�O/�+�.=ZQ���`4t$�ܻ;��t�r�,]/���'o��T`��zTƕ��B=���qo�/��j��%"8Ǧ����E�	m�O���Vf+7h}�:C>un尕
�0_�r�=�:� t�^��-Kl�+[���������&����f]�`����T�{C��C�]���7޹���z���^�ނ����u����1E5��F��]��2�tNgj;���c,ʹqd�#��7z#�qV�&].���]H�����m'lrx�Z��y�-ܹ�G� �齜���M����ͳ�ZKO�R�]] ��⾇7��Z��
��ۘ��IY�]�3�*q�/<a�P��H�݃��X�.J�83-*�뷪$�zk��ő���*���]DŋWups2���=��u�|Y�5<�@�ʡ�S��hU�C�����%�72����]�����h��x�9&
+��ANx&f��0ެ��urmt%H��{@2b���/+Q⯧��8��FT�t��'G����L���������&A<-���v��4������1U�S�}13�Ru�s6�t�����c���8�܆�Y�Մ%e�*Y��Sq�'�-���2;u}�vH���v�K-m�T�7V�6��z�u��Z�r��`N{#O!��n�˦����k���鳽��)��ͼ2�<�'�R#�1�{�^��M}7��X�����O7�����xP3�@��Z@�y�K��ܡ���S\	�������ݕ�:�9�+>�����tT�讍�W^f:NȦ�I�E[M�-�����4�&��}1{צl쩗�}HG���i,����R­����l��#H֍�c$Ӽ�D�wm�keBC^bO��=�X�G,c{�df�Ծ �H�oba����
d6ou�:�au�mo7�2^W94"C
�U���*�7.��Y�W(�ŕu
��`���hc�"�q�8^�H���t�
�>��͚%k=gQ�k�'�M|���BU�v�L�	��M^rW���ڻ�D^ن�@�rY�g�}�|a���j��	��'-�t$<{iޅ�s��Ă�N%�Uڳx3�T�ro��]Һ(ϋ�"v���Fu���-����r�/w.e�*�����\2�0Ώ��{PG_�b$n��T�<_uh�7�x+"��c�A��������ģinAÉ����c:S�I%u�-����F�oy8���nϧJ׫��L��=25�l�������U���n�+	�ҝ8~Y��A�ggQ�*r��&���6a�)�� ��2��}�ԏݒ���8��9�"i�3`�y*���lj��	�`�Y��~��Q�����s*LV�n� w۝��ˊ�aB�P*�Y����x(V/�R���,y�)��.�8�"v�b�%��«z�c.��V#��b�Gf��v��DQ<�.�N(���l��p;�Lܹ���gu������,��V�T:����⎜:ϑ��]� ��Ar�Ij!X�;\6E<���ڙM��aM�H�'�Lʌ�}R�-�ڶ��N�^9Mu/�V�^�o��K���3���:&�pc�b��:�[��z�/�vI��o��]a��b�75&$�V[���i�ti�M��Y\�B̧HG�jtn��'Q�7��Wrc��l�b��K����ø��e���.�K�e��4����O�9q�އiFzg�(N�s��p�R����4�R�z���`"4\�qոU�ݷ�bj�q(�]�E��!�]��S�ݴJ(�(�9�\�+]wP�5;^�c�c�q���J�xu$(�m�,k2�W���b^���s�yu8�����3mXͦv����N%�����;x&�>-�y�8��o�NYTɗ��u%LQr�a��$�}V����m�%�]��:�l��:�A$��u8�	:2!2�T82*Q����:	1g-N>&G�(�"�c�w�Z�]f���9qtH���;2 ��^}W�[��A��r���0j���}W�c�ձ��%��Ux�<Wm!)�v�(j��p؋����Fe�r�Fb|�eD��QL=�Y�V�{}��n��h�]�Q�5���b@&b��ʲ�ƙt��0���n�itb�bu�nz���o��1N�3��Ϸ,�N��	��d��⨓fqj�� :�w5���|��,&�l����\'�3;�����;,>�Y2uS�x�B��Ҩ
���7�)�|w�,����r�ۤ\�q���E>��vVrj�t���B��y����^.�c�pmT`�ͽv��x��81*e��<���e��Ф;��8�my�Ƕ�}�Trz �kޛ}�ʍ�1�r�sq�u�z�>�s�1�9����5_['�vvt�*ۖ�72L�n�9R�0H'���&@��K����n��ptdm>Sh�-�V�������(���U8d]��d�L���ڳK����ȝX��|�t�hK���{DgoL4)��t�VoD9V�2j�>�0u]{�H�W�oӦ�D9���5.f�����N����-= ���.�=-�O7B������V]l9jt�e�0�%&�m�9��bm�4�h�5)�^�â{a�0����ހ_Qu�Y���w �'���t��u|����*Ch�����o���Oi�|�!�qy`��7�j��Y�Ӵ����g��o��r�Q=1���sw�X��H�[qgTo��6�P������ng{���W��z�E����;|7��&[��h�s���[2;�1uor�(�y��%��H)Lp���;��KH��d��k
\`ue*ۭ���-%��h4�Ho��Ψ�8��%%��p�W�cn��`!N$cI*�6VL��Q�]�}�K�s,}������W��)eB~w��ͭ<��P;���Bk7y���e��V{z� ����I[w�I�+���C��뿇�hѮ泩S]h��^�"q�Q���c��K����՗����R.,;"��=0Dd���O���F��f�L�6J��[)�d��f�2Tؒ�|1��ڗd��67�g��\�g\����n�*��^���sr�(��{�`�pǐ�-��_u��CSJsc�>�w+���ʐHB ܒ=�N�S�m����t�ƿ{�fd}���Ю�`�0�����GJ��d���F�j6�x��{c�e�(��ns���Ë�h���������x=;�&�m�)Ul3F�8��i���v�$���x2r��S�eK�}����t���n���K�Խ�>>��t���m�ѽ��E朗�_o	NKx�4���v�ή]��Y�iS;�������t��-�7���}�j�vǛZ�ģӴ.�>�%̄�Q1�ѠQ���b�|�t�8�����S��i�9}�k���2o�^M����]g�I^y�����
3ك���6 �'qcFs
8����T+�e<ܘ�n�=Yņ�m�N
��ι����B��,�8���a����(7�W��!񢍷}��#˺�fc��Lᛴz��xT��rrm�&>H�66�>��l��y�g3m7R7���/�6��b��i�2wV�&ͽ�y,��9�n��4��e����>�0��lFh4�Zď[�v�,Rώ�2��,�]]�>s]��`�o���69wJ��Qe.��dE���{p�A=��3wI�ٽ2Q
��i�v����|u[��-�^h,�
w)ʗ�{��X�k^��T\E�]�����r��>��6���rF1�V3�u�պ�N�X�x��wLCh�RE���B�Z��܄s�a�D%��M�P[����uj��պN������T��:�_6],�&��X�0!|������$R�m�ڮ����+�����-vf�!Z��	����P��2�.�Ӌ�q9��m��8[y��"�}8˴�|vfV�I��qb#�w&;�Q���X;���L-�!��7m,엹���4m�kUv����^��`w�,���8��A6F�y��pE��D\.�/�W����������*'�����ll�c`������Ǐ�>>��>|��}�Ѿ'�t�3"���o�6e3Ì�l$:�]I)���.K1�i����D��g�4��m]($�E��@��JP �hSxS�m��ˮ+�G�ü�6eH�����؊�A�ç���n��N�Iz^U�iW��1`�u\��@�
�c~B���Y��y.f"`�ȉă�'����a�&Šօ�kT[��S�M�؞�q��]�2RAQ��.�v-9���R���|�w�
n�ul�մ���<�7qNE�s��Y]��f+0>I�WÌ�Qv�]սlNj�Dj�zǘ�����Ç)ga�6�&C�ъ���xqQ��Դ��9�V�t���#gj`$�x�F���-u�����^�+d$h�.�O��á��վI#(��L�j�p3�s-�`�0$RU�;)i��0�	�p��}/�;f�T�IN�p[.��
91��ik��h�SJ������,�;������|i�q�H}�-u$f��5�Hز1���!'�|+��x*&�}���׹��3������^���}劅��f��w���]h|�f@E�Mc�����r��s-m��h��=z)�+M�����_�
zwuӨO
��#<�\1Y(aB�_"r
�\'\�5���2'=�V���M��;j 2����)��R��|w]�I��M���o�<�����_=��Hg���,�ycģ[|��r�I�5v�������Q{�)V�g{F�e�.�X34g�n&5��X[Yk�/�z��m�oJ��p�e3u���|.:nx�ܡݟ8~�+F�R�[]uқ�Ct����p�IP���W0�t:�� \�����Si�}5=��9�!4�s��r�7�cle���-e�s�	+�\jW�y�k-�=����lw:�f�A��I͒�5���M�ܼ�dbG�V!�*�b.5^�F���f���,Ws]�3|j�J�{���^;�����|�v��5��<厂��W�`+4BS���ܼ���U���;��b̹eo%�ٚ��iz���@��A�Y�.���M��y��5����.�xX�`��}c]�ba��)�.�.l�
���q�sCu�(�Z��7�;��"��- ^��R2u<��!�ow9��ģ���k֠{tu-!�Lv=aXwj|72�bY0t��c��M�������ϱM�Lc\�v���e��B��۔�z̂<��͗,��O��3�!^��xGx���.vQv���-�ks��tbQ�^�� �ts�d7���Y�M9M��7�\e�C��>J�>��{bv}����}�8��^�s��;oi�5�	��0�gv�&:�e��4�=��2B<)�m�y�eU����Ϻ�4в֦_#{}�לZp����U��N�\ިA�6(��C��Xq��jJ�����١fb
d}]�O[=�_gs�yr2�"�thg;|ԲU�ڴ9�WYSw&t�\T��|�^��⿠�v��󅋊�+���b�h,�Iώ�r@�����KR��5#�E��[��f�'@����B�xg7��C3j]���bt�4�1�{�&�I�����,1'۶t;UH�e�vT�g��F���.�wͺ'�(��r
�=�+�3�]�J��l�Z;(-!���W��̏:�S�xz�(�	s��x;cK��%̆k�|�2/H߅:њ~뾹��z��6,���	��r{�X�e�������7x!��:2�ʲ�-�
��	���f��ChG����j�6WK��eu�1���z�;w|���+���	)u�;
�o�W3OI+��
�O�urm��`-���������x�$pm޻�h�L!ut�HOxAn���Ӫk���j�� ���5�vҳ3�q�#�J��gBx����n÷Av菂�ǅN��������[�G�PY������L۾o��vM�{��r���urWmX�l��J
��9j;KF����l6̬�1Th(� ��}G���̠����ۏ�������tT;������hQ��t�� ����c7�ԼYGk�3)'1]v��>ݲg��u�]$��B�WI���V��A#vs]��9����v+P磷A\$Jq-<�}ɼ��k ��۠8���<8�zE)�N��*ޟ����o��E�Ӕ�X#J�ѹ���V��^K9���
���r�:&��vPWKxgI�$V_*��[ƴ�\�]�dd��gL�cj2�V�H���/{�˥P0����ӛ�d�����3�v�@�c�/E��� Ak/
��+݅X��4;��Zm�{SC�u����A8�����$ ��fb��L,7��&���O�ݍ��|G]�g���}w\]P.e�²���ߝ]�e�6�̍dJ� ��rҔ�KRT�s4�jv��:��ʨ&w8,Ȅ��lzg�uN�ߎ�!p�Wf�d��_G�2B)�[�:�Pqk$���dK���1�Ú+9֭˚c�^9ʎ<�4����E{Νvق���]t��'d=c�,��(ZN<@)Y��!��`�_u�"^��H��
ǎ�'���^�� ��J�=��Z�Q�œ��X�t_f�I�bn�BY�M$=��q�df�j[�1���e7\�擗��-�h[����>W o5������:�ɉ�˹����NKp�gZ���}��g�y����q�D�Z7;bz��wW��;�Q��VóSC�Fp�̲sU@�[�dն��+�|�j���%��M�!��Tɏ�&���gBVAVOs������O_Vp�d�Nkӯd��G��:ݠ�;ad���W.��;Ly�^cyr�%|(������d+�MǛ.5w�C���NE_Tp�U��{�n�m�	�b��ѽ�:���T�JVнQ�ݙx-#\�;C�:I*Dm���S�j�=��u�����g��Ƙ���������}�y�U�#vE֨�����iǿl�܃�h�[��A>��z[��;J�hd���^1�����X���f����Ip�%^�֛��-�=�é�6&��V�z�z�<�p[��
���`��x5Ra��-hͺ��,�8v:Z�@�����hU�$Vgۭ�go:�{�ػ��[T"Xz�ڷ�m��cyBc�.۲�)kݏK�֖��؞!��
�з�(�������oIO�������t[yqL,@�h��S����TY�/`��%�ׇ3��ħ'֘�~�r��(u��>��q���G't��k�G�Yp�n[\�T.�9Q��_J[����VS�͊��[��<�f�pPS��U:	y\0��u�:#�h�MƑ4�*�K6��ƹ�{z����M��K���KGNP	�}���:�X����!w�;Z9�a�������!N�Λ���w�{�����{Ub>*���=ܹ��4\��0�sK��*-�n�+�}I�W�Xw��b����D;���v�s����0y��燵8b�K$�q���3��|�f�,VU���8���k��ZA��ց�S��@�1V�%%@�*[f�޹�3�r@II���l:�������Ǭ�{�M��]̴��ۂ��q`�VE�����-����X��[ţ��K9��.�V"�e��L�j���=-M+�0�c\3��vZTq(�_��cn	��KW��줖�kⷓ��N�v��T�u'����/(Gf�O�cz�r��}�V��i��ѻ��J�]���n�oA��#%�d���[;K�׆�5�ܚJ��.�{�1���o���%S�J{�)���WG�3b�����DB�0�0+0�P�;�3n�n���ݷY�&��dYXS$��܌Wi�'���+�pق$������R��H=�gS�l�&V�f�7-�҅�e�����c�f�52y�+N�fop���S͆�:܌G�Pf3i��V�"_;�����W.�s���7>,�^����8XU �(�z!����9gk���Z@�l\щ��0�B�����s6��β[[�5&Rۜ��Nv�۰���/�ܾ��t{��zí�~�\��!�7;y�Wtj�PT��V"�Mm����ɂ���ǧ��u�H��I��\�ꐺ���1"
�]�4>�ȋ���H��Mun��XWq��&��)�j�-,_G{����X��+E�ƼZz=�PK�1'&t��+r����o�З-��7��s�F�0��J��X�I�ҹ�vڋC�N����wÃ���c&\y?�q�;c؋���[��ޞ9�o�C��nn�PV�"��W�d�ˬ�xM䲋jM��ֳ7�ӛ#w��1徖1�ə�=K�"����<��'�	,����SR����G'5�q����5}�na�g�]�m^���ѕ�����u�u�����ᴞf�\�n@XO[R�䢢�����31(qgJ?]��V����wZ�.Ëb�اi˫AX�����=��L���{a7o��פZ3���1Q�	��Nܻ�H��Ҧ�ÕT�j�w�Z����bH�h]�Ħ"�_.��w��$݅�c�f���s:ݱ��0]��:(�$T��c3 um�4�p=���r�a|�_��&���5UOOB.��VI�l�A^�PZ�x�����Ή儡��Sՠ�[I-�yn���3��a��{�g{��т����\��.u�!�\Ȩ]K�ί�nb��j[�M��G��J�Ra4�1It�k�ݲ0WW``�k5�����u;-D�8lг�!���rWat��tz�'��@㕅����B&׻w.>��G��%��iޯE{׈�s5��_I����X��v��^쾹p�zE�x�j��e�X��N]:	7J�u�D�j,R�̶:ٽ�W[��e���N<{����U�9O���Y�V&{�e�%Ӳ�ܪ�bn+èo��3�����ڹCm8�N��K[�}���A��YTV]X�4�|0��GkL�W�&�9nb}�H)Kf�D�Z�L�"bn�R���'{'A1jHa:T��>|�s���c��(�+��s[4����A��r.3�N��W�{"�t�Ǩqf��d���A���y����y�PW9U̟!�8��bԜ�9E�R�Vq���.�-u����ŏ�Y�U�5�N�'�Z='0=s���c@V*��Mw��:��*eW8�c��K��Mt';)��5�r�l��&V�� IsS!m�X]�gus��WO�2ʾ3+Q�% Z�6[�M�.��&�+&��Ԫt��{����uf�ܮ�����{��k ������s�|(��*��8Yry���Ǖ��������,ev���;ݱ��"��r�Ģ��BY����۩��M�e��V(�v�8�+�3kY�֓��������M�@�=�b��{ҏ����Q��΄�	5���x��Wڗf��4ծiRc���xN�k]���a{nCN�eg �E;��y�;M�v���;4�s.��.�S'}k�����k�j�Ct	�y�:诒j�vِ���Ǎ�첞�zk����+z�엯VpkrdMf�����U!D�˾W�9N�6��ޛq4lճ�V�YW��tؤ7K5sg�J2�&4�|��s۲T��ϖ�4��W;�6�6#��k�ܥp�p�Yo��8�N����l�TEs9h�`����Բ���Nփ�3��kj r�<%*e�������L
���[J�*־c쮮y���l$�{�[{�{���B�E�mv��������
�q�]E]��}��3m�k|��$��!�Z.Vn�p�u�Y�6��Rs��r��an6��}�7�,�s6��LqP�,}�n�Ɔ���:�&Sյ�l8��ܚJOdW:gG�z�dV�*�um��Hi̫u�B�0�ID��t&Zq�:{�r�ʶ5w[��&D�81�d;��Ѻ������,U�;�l]��[�su1��Cx���k�MQ��9�Cj��T7�y�P����2�zN_r���.�vi�a�s{�eL������C���XǻD�Fp���E@�.�F^�h�6���@b�(�n.��w��7-^���1�'��rD��ˤ�t��C;��{~��.�e����'4��n��mr�~=�m��h���0�A�GT�Ώt�އ����-�v5��U+δ�b'&�����r����[@e�CV��7���0�4Y��j8Rʖ���F]�ǜ�M�Zɽn���Fv���s]ก�Vε���Zƒ�-L�wI�q����i��p綛�R��@�-�:�܎�4YлS�����u�BȰ-�G���*v����t��
g8�H})��+8u�+p����,v�wA�Vb���m���̜�ɵ#�m�*�4�o1\������U|���ʻ(�<��V�ݬj^�Ƭ�)�Z�jm�T�r���ˎ�A.��r�3�:�^��/.Yv�+-����{K�!��󳁏pw�.ݦ���e}�L��K<�c�*\�ƣW�й7)��d�/U�q�[Fc�*��vv���p����v��b.�|������}E$�sl+�\1u�n��>[ږ�(�dZ�d��3p��u��]�d�RM�=u�]�������梵�z�8C�w:v��D������nf�~tZ�rS�M�8k�q.ʊ����|�����ٻ��'gE�it�{BΣSA�nxj���z��0�$�b+�O��<��)��C	;X��V�ku��R[�2�Ħ%g<�Jl�eɐ�Y;V}-+�Ï}��:]��e�5/��ҭ1�e��g��/�b	i�[8������S��[)��7���؈�n#�Y�S�u�4�lM�ȑزvu�Y�����n����Xy��R3��e����H
@K � ���@ɜ>�Ljɺw)n��W�W�U}_}�}���&%쀥k�.��p;���5eGs���G�Kޤn�4kz8>���i`�[�!�-��R��ǝ�Y٢��P�9{��t�.��Z�y���W�0`�f�_JǱ�Y��*�le��S�bl7Y�R��A�&q&Z��C����B�����JZ5�*9OՇ�G�Þ���[��Nqj����p����Qod��og�� �T�ؔ��Q襜E(��E\��Ƭ�e�����'Y�b4�xH�;�qPK �NV/9W�����`�LPf��/Vu�5�r���-f��9���ٳw�iq^��Y���0S}:�5P�m�'R�s�%�㼺�S\�����P�sz��������� Uѫ�� �.�W]:^^.��9��WE�̹�p7x��K��Ca�<�0z�;�/�M~+A�Kُ<nͫ	*]��VcZ`�|�շ�=��b����8B����2�6˫KLqL��ۘhm=�*���O�^C�'P�`�;6�h�M77����h�hc��ۤsA�m仂�����(؍���o�M ��l��MdQs)�3g�b*�g\#^ɯ�9O��:�&Gݣc��f����	3����;i��ʮ{ۖþw���0<
^+�n�v�h��q�A8N���૵L����4f�㵄��ep�����éq ������L�tNw�M�>v����T��V�ݕ�7�˸�_d �[K�Ps�櫘DUQEW�y*��wIEF��na�������.�e�lC:�"��йN`B�EWs�9���^��xG���\s�ps�N���-%Owt�L�Ўx�ʫ*4��\
#B)0�te�{����8�f��9
a�M
�\���9y!���8��:�f˜��1i����sģTL@�U�'"�J�wUQ�G#4�Y�3/D��9,��iRU)�*�	E^Ip�/�rԂ���t��5U"��U%FU��KҒ��FV���q/K$�0�E�w""<��"M��e��xFdU^{�"��l�JLw;��^eeEW���4*�J�+	6��LM�&��4H��,Ң�!��HQ��=ȴ=7<T.k�{"���+4I<�8������!V�m��������χetm�b݂�yˏF��R�,�7(m��B�'^�w*W9��oM��X[H��n.��6���9w�Zy{g�9�d'���Oo�x+�s��S�~Cj]j�{[U�:��컥1�+�&��=�Q�"���yd6H�!������ܩ���>gk�V�
�m.7K���o6r��aZP���uP��z��P�I:8���\+��c��o�q_�8aK]�\hIo����]�nZ��S��g���{3��[בx�аthu�Ф�V^tU풠�D���^;�!��Rnt0�p��[Q�9�C�ZoM{�Q�z�0kK]�+�'�c�k_X]ًd�ǙB�tV�� C��`WLSrE�{h@��߷��*�5�c"�]Lw`��T�����<�}C"�V�h�I@K���B�L�f1���wV��^I'�z;u+ku������Uv�FN�ip��S:<����_���{v(G#��Ӱ<�;W�+���v� ĎO���7���x�;���P@��R��-��!�[0�s�����3����|������XS)��Lh|^����q�V�Z],@W�%�3��Vr����м�\�#/�R�P�ɑ�����d��p�Q������Q�J�#x�\-Yz�w�'�l�l�;��GM�e���$����R�������zZ|��Ƃb�dտm���s��R�ھ�7�9t�: ���>���x(5�Z��Z�V��j�Z�b+&dc����~�h�8��n_�jy}6*�Y:�2��4�鳃bx
i^�TZMt�pL`�j�Nw<����Z(_6�׮'�� ��7o!�6�z��<A��W��,��yq�27n*���Y8:Kn,��#es��
܀��nzo6M5���v��d��v�����Em< $s�0�J�K�L�<�b{lodI����m��u�+�?FEq<��K��th��4},�wT
gt�
�&*�c�ފJ�Ղ�yƭ���"� jmY&��8�Og���rB�1�|��{LN�g%][o4m+ï���扅�\������r��v�j ~�N�3+���Qu�$u$��Kva�ä�Ln	�%��fO*~�4)�;'޺��:��[e�y����,n�,J�t�^U9�:�&��<�u� W�K_��%'" l�uyh���+��[Nzwr*��>�s����:q�rzo�
6��;�bp����k�M��C�B��b�ʍ#�Έ�$�1��xsgfSB{�!��3���=|�w�ـE�u�J�3����$�G{}��`j��*����t�8N ��˟V�s�OWۯf����z�%��(o�7.v2Z���������hAԢ%����I�YC��;3��u]ʱ��mn3ґ�#��!-_=���C�^&�<�wl糈4t���x��a�'�x�V�]�u�k�X���v���jT��Ú��k�jk,��wC�!0�����P�H�%�ћ)dι�ɧ�w.�n�f�$�d�q���ݰn�g�����W�}�x��ģ@�U %b:��j��յ�k��fg�^��g�$-�l�=�KҼ+���m#]�G�ƕ
��uץMۗv�4��%�ZC�V���p�+��UȘO<U4X��0c���y�zT��C5R{V�ث�[�M��˶����:��b5`�J��������1¢�E1�&�G8�y�6k0��٪aƫ�b�d�W]5��}a#��PyN��
2g�A�!C��C�Z�ҝk�Y��Rr8��طj�\7U+�v(����T����j�l/ ��_Q���M���;�bn!�[�~f4G
-�g��)��t�H�j�o���#˺�+�yr3�ȉ�Y{~��𮵱;C�R�0�s%��Qݐ)K'�#��p�.V�JZ�/�Ey���݈6\��-�.�H���9�
�ܺ*�L|#�mQQ����\a�c�|*�%�1�6)Sˮ��!b���S�c��R�P������{�����˫D�y��J,˺�{����q��9��=]�
Ou��xf^��'*b�=������-PV����>�<LP��V�٠�{�y���N�nʷ�~s�"��'�<4ZVi��Ra
�j�|Vl�l�b�)"e�M�U�v,8&�>]'� ��A�s��ok�{�-̩t%<����ޱ}�%��t��9��w���c����Z͗_�*�q/�������x�|�s����t��P"��b�Jq 6!�ee�1:�Q9��Cog��Q�~�ɌƉt��i�ޕms�:�v;ezW_�^
�{�7��*`vC�b�E��q�Ir�{e�u�Ck]zTB�ȶ��Q̺�!>[ɦP�ɘ�P1�1��;Sy⧦2΍n놾�<b�K����&Y��^i�n��etW4xT\�"���j2"�]�71�.��v�nsz�����\wD����Q%Sq5�r��1Ȫ[w	��������^�^�7�;��K�7U��Y�}o�O_�VȬ�\�Z�Y�<|�;Ǹ�JWH6=�8~�+e��òJlg�ort���q��Pr]DC�T�G���m��H4"��a�f�x�ᜌ����FBVV]wH�f'����g9��7v��8Sg��V9�wjgl7��l��7]+<V2u�R��7"�י�-��C���2�Z��<�3��1�=M��,C�#J-o���x��pG��ǅ�#]4�/P�]	�Ͳy�r���@�m{%�5���dG8T��>�4�W�9(e
��ϻ �d�/�3�]����h��{A�-l�����,j<-�zy_�| �K��S����؈�a�grI�ޅ{�K�YRo�`��� :
G��H<�j�!p�hEx+,n���*��:fȚ��-in���D!����\�T��k�pW��iu���"�{V���s�1|�N����z�!�yA|k�4�e�dk��t-.��&��bi�vo�]�g��y�UȄ�u�6Ԁٸ��~��I,"z�B���^W��fRa1}2�0�@�l��M�{��ٽ�/=p���K�U<�q�>������{hzٳ4�G��+:���1o�+(�<z(x�n��%�Ìr���޷�ĩʌ���9�E�'�t��1=�4�Jф� ;z����[�uV�C�| ����<��K��r�nH����p�hۇ�~�!l�5��p�:��ӫ�G�=��"����mBf�Xˬr�R�sK}Pfv���K:���2G��gG_`o�w�vc����c�ffYܱ
�2"�{ ^\���we�Y�@�I��Env�w��(c�MD\:��9'��tY��IY<�^UI��f�����~x%�#���^��Χ�C>X��u������ʾU��3/M:ԩ5&��]ie�	q�o���OB�r��g��u}'��]�eP�HRbɒ���#tH=�� ������
�.L1ې�ۧ�C�c:v� ��xh9)�L���V���Qƹ�]֝���Ģ�)u�R���ei{�3HƎ�茐'�N��e�P���Xü璝���K�ΎO*�;�n��#��pdwM�/�«w���mTGf���%�2�u�	������7��k�����EoO<\w6��pv��9]�w�3�W��gsE�o�5���1�gk�2��1��,8LpwknW�e�	)�q��� K�Eօ��h�e墱3���fG)f�t������V�Û2����%>뉴xnU� ]�K�N�y��zE�|��y����r<�Ip�N�1*wd@)��;�wqiiT@�F:��݋���p�Mz��.�E��Y@u���b �ai뛤"��
�(��7�2��\���䢫ҩ�z{�K��g��]�����aWc����It���M��)R��T�{�#�B�*���t�D�h`q;�5lO&3�ݚ�d�޵Х�7���y�JӾƦ��Sz/`�:��A������vM�s -Y��8�;���`Շ_)LW۝��ڱ�ȶp���f���{2�ٮ�����{��i�����%����$F��!Z��ȭ��8�Jb���0:��6M@c�(;�*�X`�0�H��ey© ��`�{��q��@v��v�;^���a�q�Mf��g&U�a�I['� -�`_C ȣjo��z�O+�C�R�?�v��D��*�g�|�7ݲ����`
��r�j�����N�w��O�.��(>��[�N��>u���jY�8kU/
D�����+V�*s��&���p;N�۟y�������V7b"��\��uQ;=���1�by�7��۔&��z�1G]{.5;`�=��q�7M7��p�4@n�ԃs��b�C�仵��;��^h��U��%{�o#�ֵ�>����^��v;nq����1����_0�w��/{�J��
�q%�Jk4��fT��D���e��^��nXݖ1��X��ۛ��?C��]��Z(T��
����f�%*�ps+hJ��<�"�uي�1sC7�X�ө!�0L�{��Y�$I3�u��%!�|� �<wz([�O�����@�7&�(of�W���6�X��Cl�V�R��=?o��KB\(�^Sa�o������7�$nw����"0�^�Y�y� �lu<z��ӻ��W��?ŘO�5�X�e��HJj	���s�	���\D*B���W���@��X��_g1&/���|�24j�N
���p�T�ٹ���P���+�˸��蓉�W*����H�cn�IЙ�As#��#
��ydU��%�&8mLLs/e� �H��k�y�:K�S0\��8C����§1nr�L�3�����Q;�i'��[�:a���~���8'��Ј-Q�X�Ȏ4��B��\�[9����@=�=��Ck��5%�n��e�>�A�^�裮�o0��"�1p�)[L`����0��V�al>�<�-����۱"�h�9� Co`͎`�ok�{��R�m����;=���8��]?o�9Z�Us�9��ڧy�wp�{(`��t��*{ �SX�ʱ���qm�Ywc�*N/e�����j����s��nD�}�~�s�o�&0Pc��e�Þ�a����m���PwG�L�Xn��#T�:�\1�q��<�q�?�b����.Voz��ҭ��C��Z��w������W�8�^���GA�J��]%x �P�W-.�c9�o��u��q��.�-t��vb���גV�C6�̺�nzu�7ۦ�RztG.��y)1Em^Ny�;3�q@�r�v�n<�V�@�Q;:%ZT�b ZZ��L@窟ȣ���=����.q����1|��]�ҴɆ�K�DP�ɘL���������:ˈ��q|�4`�w0h�Lu���[����'�%V��ѷYIih�w)I�F��@\d�"�f=�O�����sW]6
ø�#��1��=ԅ�NQȀw>+ �(� �|�C�{*;���X��l�&����滅����i����̺b�d#���I�z]H� �Dp�{���LwW�9/��^�R�6����s�<�#�-��l�(Y��R�{f�c�<�٨��=��;��职�������¸ƯƠ���7��NDk���}��ls컉�o�s,��9���.�14t<6J�|ep���*hEx><1�0�õo{y�j��	��dQ �"�Zz�@Zjؘ�][F���&��LV����9��rWK�|���.*41@�7��L� C��QyDu[��Q�i�!w�'i��mJ[8�}�A��E �(�+�)8�9|�t�����C2�z�4�i�՛a$�TЃ����º�n�*�}a1Lm�+��U����g+e�r�unX�(p&��I�|%�oK�2���;����ȝ��m%z��/�ݙ�wz�)M�y݅��W@%���_m�ޏ�
�-�畇�7-��°H�qD�\B���忻B��>�����Oׇ�& �fui�gɗ����>��<���9����S��۸xQ�~� u���ř��D��[}a��{[b�A���pH��Τ�T�mW\p��tt�<�����*¬���3Gzwly
�:aC�k��n�?��< ���Y�
����1M����~j�m*��r�x<y;Io���=���	�$;-uW�O��U�lܔ �~]nϖ�d�PՆ	R���}.JW˫�R�w�C��Bp@�fu��._�.'�)xx�ݹ�!ˆ^�݊OcUX���awu-/L0��y�s�4[�ód	����(��v�w��mo���˕ܠƅ;�)0ѹ�V�=�e#��cE#\c.7�;- �� W��A#@.[��t�=D�k��KE,���"���Ȁ���Ξ��ޅV�צ�p�0��%��KD��Kݵ;��v]�5�4h�TY�V�.�"U��C�U��{N�A`}_1��]u���5r���Ç���:o�#�m�эTN�Ba��Li���!����1^a��6b����-SF.���Š����gX�('��{&��ر;Uٓ��vh�	�z� u�eE�N�u; �x0:W�2����`fn�g���>�����<qwRW��-є��iP�e����.\�+c����{}���bxV�9�Y'��i��۠�5���wZ�`:W`ZVJԩE-��u�m�}�WY��Î�����3q��䅂�hA��Nh������<�nC�U��9V��<��Zt�T yØ}�o-��O��dў���$xp��5ذV7ے���3ً�)�iGp�� ��U)&��ab&�ݮf��q���P���nu/R�鑶Q.dH�ב�G���-�1�Ӄ��"*///���>�`eZ�a����xt���
2��k��lҁڵ��i���ho[]Z7���ιG��I=�JF�f-`(J��Zk3ty��jQ�1��m��	�]�:�w�c�*ZI��p��$�tl ���*a:1ef�:���oB�}"ˑ�v^,��N�Í�����kV��/���k�`]Ձ�K�*�-wc��zv�|b�',�i���f�Hn�{�g��!�9��n�{Zj�b|'eQ��j<�и��jo�<�)I�^���yԈO��"%��,��i�E��8��j��-���n�c��`�i�2�ȅ�w늡lf����+7-��&c�WׅD�L��F���g=�?_,˷���`O��D����"B4�t�rUK�N�۶�r�1>�8�p���m� ��Ⳝ����3��.���t5����쎸u;1�+�`TWF1k��{�u���hвxu��4���9����F�!�h�[�=y�&��/b�+Y��}��q;�w5�S�θ ���1�W^��s]�%_V!:>�`���6�բ����EU�O]2�>D�̥AD��j�B,�pM��ul��Y*�ȼ�J�QƊ�h�t���Q�C{j�WU�官/�����u�l�nu�Rm�&��"tR�C) r�k�}���p�k�z��y9��,���3�{ohp�&�F�>5��u�;A�M>Nu��"إ��v��h��W���f_p�{#�ԥMchAx��t!��v*-m�m�pJm�giB���&��A$��[��oL�Wg�,��Щk��s8=�@>?s�G����z')*įz�����j��T# �|,k��(mP֭C��)�Ԩ�3(%��{�����{��gam�jsw0���݊W���oFe��냞�U6����h�/m�W);+��á�9A9�󧖝���L2t�����t�-��к��}�D�5 N3��Ly�m�\�Z�f���q�1�g��o^�jgoW�-t�<2�yr��N��qå�j<"nmm�0��aCI�E.�өM�I;�����t�k{UM*�.MS���
��8UfsT�n�̄ԜJs]�|w�&%ҍa����Qs�_/��y;ßr"���,�����F*���\�K$UCZN��ieK���bQ��9��4�4���D��
UW*U7'vt9�W6��{tKʤ�\�RЫ�#��YR�D�X�F�Q]Й�0�)29y��`UU��"�C*��:�9N��0DBT"*�-κE��G���Z$z��"dH^*�桢�kCJ��="�:"�4Trp�Idr�g"s!�2�M2�4(L�(�4�tG4I�J�\R���:%Z�wq��MQ��)����t���=iݖ��)��S����������%Fl�r��/K�#�r2�%hU���y���aDI�ӪP���^����dN`�B&"�s�"�e\�tr��@�u��S�K=�L�
r4�L�l���gH#uqw<\P��5�WC,�
h[��^����#�]ұ.rNZ��z+�3g��N"�
�}�+*�c�Cyr�]39 �Ԝ�^�	��m�����:�⇹�q-����v��Z{��9��I���H�؄V�ڷ.�nH'D+�,F�q-�K�����@C�b'�|��� Y["o��s�����ÂC�}OG���<�&�G�~C�}C�����¡�ğ�������|C���+�'���D's��!�zDB�=��}D(������ЄE��"@�
�oHN��y�|�����Ӽ����?<�L.�����ʛ�<�*�S}O�όy����;��'���94��}w!�=�����aTߝ?~�|w��߀���vv�K�f�oOޑ",G���< ���7;~���<��BN~&���zM����Wϯ޼�7!8~�c��-�'�9��-��O�i'v]�7�/֓�\�G��?����n�ƚ��X0)�2ܟ��.�o��˯��ӟ��0s���yރ��ߺ)�\~O��ߐ����>�?'!���������tﯣ��7�ێC����+�����xL/��v������ԑr��4�.�Z��ͷ�f��(zG�D{���W������ۏ�s�����!�4�!��㣓�8���F��w�����ǌ���������	������㓜�;�O�{C�򑽍�m^����ō+�"$����#�S�����U��H��׎���<;ry������R?�ro�O�o���>��C�k������>��}����T���߿���p)�'�����}u�N�ݬ�9�0��H�x��������'!��nw�>;��OG��)�S~OO!�=!Ʌ��opxAw��nCϿ���7�$����=��P�N/��Ǉ���z߾�����y�#����(�ɿ�못��$	'���|����˴���޼m;¸{?���n}8�9�><��?��]�7��G��A�0���=�'���I��s���9���ӂ">G�G��v3&K�B0��Nfg�<����>�x|��9��������g�ݽ&On�����M��O?~�����8����oo+���M�	���9�x��<!�4�On<G�����?�=C�������|�qj��mW5�>���zG��z"��"#���=;�Nv��}�{w�9?��w�߻�aT>8���<�_(~���%w�i���9M>�ӷ{<q���i���x�����,m�Ͽ��������ϑ~��U�h���ȻD���g��e��f�)v.���C�7����lͻ����q���J���)ug�6�o�R�Od�n� ���{y�([7lN{�����a����g9� }��e�2tU�<ss��&sv ���}�Zpz"DB#F">
�׏�<��$��r�����<&���>�?'��O z���P�������s�^�������r�߿����]�|��O�s��K��Aw��nGc}��W��+o� �غ��P���(C�>��� �͏���\I�}����Ǿ�;����<8������6���c�]����Ͻz4{�Lh��b=Y#�.]�}��/�|���������!Ʌ�~�S�!!⌿�';�xO'�y@����|v�~&��C�������c��}�I����{�|�A�7 xK��v�����ߧ�DP�=�$G�����許�U���vj��F����0{�?�n7��",G�����<&>��)�7�˹7����&�'��.��3�N�S�]��'!����ߐﱿ�~?�I����4���#z �k���K��8�RY>��~��F =�<G��BS�"�CM?�����yM!!�5���^LyM�	޾x��o=��rS�AΜ}~�$���I��y��90�����S�z��1<ǡ���{�+Hecq���~y�U��k~��="#��G˦! �P����!�>�������q ���7z� ���Г��=���oN���@�|O��q?~�{O���n@���<��xE��ϗ����s��j�ל�����X�D}��Y����^���0yC��!������=&xC�?�7��s��~��&����~�<3���>��z�y@䝿�}��yw�Ï+�*�5_R\+�읹�Ӎ��l�h��_������>��"=""+��<"�����}n��	������e7�'ۏ;��?'��w�߼^��G�������vﱿ>�{�n@QM�W��W�zG�A������Br��}�����?��_�P�;ێNN@�������/HyL.?����>��90�<��>8��w�׾������>'�X����}���1&��������}N~�3��*c럄�zjc�_��\�2�-��Ͽ�~�����]��I.}x�4��_����'��'��x���'8�����yL.���z=���O�90��V?;���q���q ����8��$��_~���o	�!;��w�/�o�����r�6��5K�%�L�Q�FѠ����L���1sx�M�\�6kG>�������7O&Ta���Uᨋ~����L���2��.E�\��q�,��[�*���s���^-k8"�T����V�=������؟���z�i?��9_�	7�8<8�O��k�^	)��7�nEӴ���m�ܮ<�&���m�=u���������������{|&��;}���»t����G��&(2"����<��t�_�/������o��>���s���ɹ����<)�]������&���Oe�ߌI�i��"��������|v����݁M�	��;�����&!LU�?��܊Y��)� �����������;��7�ü'���p"����w�~v�7�����}C���'}?~�cù��ry/�^�	�P��}�ǔ�=������9T=�7�b#�D!#Dp��/vs����֬wvg�?{�G�Db>�b*��<ǯ1�:=#!t��޲b!���97�~v�C���q�S~BT��M�>�8�q<�?@xC�S�y��ߍ�=&�>�����
�+ER�	����;
����M,_d�$~B<G���"${�Q��x�����x��}I7��G���v�ߐ�X����;�{��q8�lz�~~����@���ߝ���"��o�l������� ���������ݪv}���Ϻ�b@o�Ї��CЖ̓r|NL)�{���	����z<X�v��o�������s�ˎ@�����Ǘ]�����>�U�P��������w�G��Ϗ���z{{�G-Vs�vp���DH�=x�1��B=�	?��>w�p)��>w���m'���!����;x��Ӿ�_c}|'���aW'x����.��2���"$y�E��T`�@c��4��Z<�~Q�z)�0Dh��� ���c��>��M�{������������P?$��i�}������o�H{�|{�yW������ӵ����&�8�>טw�i$��>�ʦ����q�@#k6���ٟ/��X�!"G�G����ǧ��>''���ߝ�=&~Oe����@�w�S~t��!����c�8�]���_����I������&���9Ӵ��	��>����#�����}g��ݶ�R����8G�<��~����iI���	���X����	��C��?�	�|����o��90���M��������U��N<y��P�_�ރ�z�y
���������(�[Pjѽ�L�Z��	� ��b��t�Q�&]Ѐ�㝵�Z��]��qml�+��ݵy�T�kS�`���m������|^֨�rZ]ԛWĸ�3��Ybugcy9���\��rk��7 �����,܈�ᗑ��ȗv���w�}~&��9��U�������P�=�O���i��u������w������7�$�����߼�j�Ss�~�����s��'�������<8������=��<�J�+쫙��E,��|w;�u�?i0��������0��v����{O�Ŕ�]�ߓ��S��&��?�I�hs�u�?P������< }I�>��?S�&�����G���#��]��0�ik� �zv������oH&�8��=����aw;I����w�iP��&����>'��o�����w��'&{?x>;���q���*oΐ�O��LP�@z�_��9��_���֌9|�=�+��D{DD!{�'�y�����H3~���_�o�o	�!$�?<�����zC�Hy>��<<�"�e7�/�o��
�S}B��I�7��LB">#�"�H���h��i��B��6�e����{{��و��Tz(�p�=~�HxL/�wߜ~ON�r��x��:w��n~����=!�0��_}x7tnC�|B~�;w�=8�ׄ�"����D���W�DW
� /��7�!�?����@������� G�~�a��^#O�π�	��x�	�|���k�X�}���n��U���p�;�����?\���{���zOI��]���� 
G� x�<D 29����o͆��i|��DPb!�D�=��ǨDB@|OA�/���ɿ;�����ךp)��P����x�����!�5[x�����}�~v������zT�����ᯈ���+������QA�k�������.�����J�,D������C�p�4��f��Cg�,_�	�]����2x0�䍄������G�Z����s���u�������݉�a#����o�KT�-�ٿI@V�ݟc�V�o Zz����]��b����]o��k����N8Jvv�����1����F�;�Xu��s����r�9�1t	���R�yem];ę��D*�Dk��Vu0K9����4W�g����T�
��ͣ+�k��{j��t�yzцi�Z)��N\Ώ{�򬬚��w�7t*"[ʈ\��4����6wҸCkv�}���k�x�tl��X'��m+KFe
��Nь��R���f���/���W��ӷX�@_��tTԧ<�2��v�N5v�dc�1���&n"yՆ*�7)���ɍ�q��0��x�(�!��3�r���e%��k@�s6�J�&�2x1��C�n����=�zkʓ�*��=�K�*��9v1���l#��K�QdW�wB�L!��enΈP�֊ͫ��������g-��1��tO�����j�2�7�HωЕ�u�Ζ�c��[pz�\p�o�"	��K�x�[��Rro��`�nH����嚅 3";���V��G2��~�v�:����[+�.5~s	��wXcw��R@#�zeF
���{�":L3�ﳲ�{5�,�l�����z��b�\�.IW swD��&fai�':a۝wNfp������ӵ��Q�ˤ�^1�}1�)��2�ڕs1�ʙ���|٨�6��L�Ĵ��Ac����urN"Eh�&�}���΢��k��/qp��p�%L7�$Ċ�ʝ�y�Ss3��b����w���yߧ'n�s��� �;+��Y�7��t��Je�꺜��u��i�0r�QP��	z1��Nꋬ��p��o��=�d��l؉��rb�Վ��(��9��ߖ�/mg��A��*���3'�Ҁ�����7����Q���lʤ{NE��?��5ҕ�zo\�3Qu1�����teu=��_v���4�Fw�����([X+���t<�!��7�+�G��0�YM��bu¾}�Q��2�Q7���+�(�u�0��a��l�'��6x]�Tp�Q���EeKX�ݹ�q=��x!}Z�h��{���EBy�4F��كW+Hj6y�C�;n�����\dΩ��B01ϭ{�����q�cX��o��h�>�v1s���4�bs�*
�&{��_E\<D���5���r��7������c��(��s�DO�Z9j�{�K�c�J�S�U�}�8dzzk�H	�N�d�a�,���
���,`��p_2F�md��Mt]#˗�������d�C�tMVy���Ws�!<9��KT�Љ*��2J��̎ծ�F�=P���S���\1�jO .��% �T���$x�Q�/�[i7,���nݭĨ�Ψ<b�g���9���c��n�H�ꠅ~�o�z�����?�#<&���6�:� ���ܝ@`n5F^=}ׂs���}���̗۸��g̃�5˫|F�]
3�p%�|�I/�{��Qg�f��B���8ͳ��^�T�t%ϻ3����/Y��WY�)Y�e/�.�Qv����!�4�'ns`���Xb��4-9��٨����DΆ�jc�
 ��)ԑ��T��:���e����@�B�]�>yQ�ߦ&7.Y9]0� �Y�����U��yU�67�E�U���mN�M��}� @@=�	;�Ӟ��zm!||.���S��Ɛ�{�x�%%��@��T�]�$b��,qb��9��jei�Q�l�y��<�Ug�yv���U/����
󀳴�0�sTந;� n��A[�mnx&��U'��j.���qv��fǏق�0]��>���c\�e��6��ye7�c��fu�V
�7�1Lɕ��5y�{���5�*�7��S9�S�]C�N�N7!��e���Z?A�)]��k�ԘOZ��rꡣ\J��D=��+k��V�`s�#��֣���O��������M���_k���0�
˓�\�1sXP��Tb�1.wCzS<T��L8�e�[˜�v%��o������xԫ����ZU�5��d��ב����j���Qu,.��W�mR���F8��q��>q�<��}z���7:,[�R�@/�m:����\�-]��e�'��;�[l�e�=)�=^�ep^9l��^^Zem�e �f]W��c��ܰ&Hz�@��:v��J�q*C;��ލ�x�r�s����.u5Ӡ3�װ7�xol�騒�Sq5�s �"�-��T�����{M��6�'�\��Xxo�1���͜�`Vq ��Vy!�*�W_aWgZK_��QR�����=���#��3�9B*�yC#�i�B�^�z��&�N�	�z�����މ�@��F7�xh��N�1�:[7}�iuC]kk��.f�����b*����z�b|�"��W��g��SZ�a(���φq�=�zyC�8>w�!q��x���$�^���zn�7��*U�	�VW:�D����ߠ��2����ڢ�dJ������׊t�Nk�����Hn��Y�"�J�� -6���)�A���[|�f69�	���Ʉ*�q�����Cro,��*+����xf����ҥg���Qݳ{��jvd�%)�G�		�Q�<�8�P�>�$�پ�B19����y@S�8�S
�Z�(K���Qs��I�]҃�'���`#UN����@v͚��ܦ��u(*��4��j�-r���P��0{3Ԝu�̠Ͼ$�.,�+��5.G�b��9���0S�A4[)ǖWG3Bo`S^;�{\��9w}r'�t(�]��-|4�}{ -�Wc�=��Wek'�CM�܌d|5u���]]��;BxE���/����%%ޢ�����yX탃���B*�Sn"{��#U��1NT!���eV��
��M���wnA}O�o�kb�{�n�h�����B²�s���`T)�nH�w��3%���.E-Z({q�ɻs�vXv&�Y�#�}���/^L*�[d� �Ք\���ӷ�U&�%v?.���9�{�ֈ�&��1�a|�����\,����/�����̛���B{�����Œ�X=��N�����u��Q�P�~��G�fȓJ����>>���c��ɴy��~ݪF��	���V��~|貑�jc�w��U�uձ�����Y��M��R�Y>5��eZ�º�A�7~w�Z8!���n_<���D�]��F���Y��1�6��U��th�C���<�ԕȅnth�����iu�N�o�kg]c�V��삮q���~췐�f�P<��zLlt�牎���԰�ۍ�U_�1ꋨ�!�e.9�R^9x:S"��3p���cjBF�ȿA[OZ�}�!�]�R�3:�C� <o���1�1.���nI�����lf�wX�V!^�6�/8�n:���8�Q�6?e�\Q��OA���#3 ��oYn�|�r�l\\T��[j�+�h��Jʫ���YZ��|x�V��  ����]��5g�?������4�ooWI����¼�o"I��{8�n��H�%OI��8EA����l�w)w��ۿ�[ؘUs�BUYDrf��K\�.IW w7�Ib ���^�8�&�JϷ�6���r��a޺�3��x/��3�5\4
[5[���3禢T��庄jqtl��a.K�`$I~g�xn$ƆfavFT`U�18X!n.���<Q�FN��YG����#�j���&�2����"�^DՃ�g��8��4������X�Ka ��Tb�f]n�sy�;�����F�*@������%%�rR�\��^���X�竳mNS�Ó��z�����r��a�=�+L�J@��+@�>u�g�u�q�e��溞m}&��X�x�g���> ڵ���O�:�骜����".�M��9a������Ǝ=�0d*�奞Usho:�v�l�O2��MD7��� 櫌�
(	���Wޛ��`w>{Z�9)�E^�+�%�h���~��>:�!	�ʫ쮼b��H��k|r�k�����1s������G�b��ۃ}�l>�nU�xJ3o'��7W��O�hϧq�c�7�W������K�0+��m@X�f��|'G� k��1�7��V�V��>V�hSL�P��9,x�*t�5��%\{s�������*u������j(�m:���K�c�L'��1c�j®��t.�]tg�3�sb��
��k�:�[�S`r��X�x�\��S熄�V';밠ޚ[����T�x�7�4G���ȯ���a֘5q\�7N���!��O��f2�]�]�c�r�`�O�K�ӷ�[��6꺳r�:�m�!�u����-D=�)%�y֛w��t�ʥw�&T�4�m�\pQ�Mr�"P��)*�b
��ޚ!�뺲��߫;�6C�� (�x�W�-�+�n^�)��݉����z��v�
�z�Wb6\r��_9��{�t�.R���[N�/le<�(P	>-@]��*ۻ�{�z��K
e��4.������J�F R��]&�����L]�Y�z1n�>ӂ���c�'�Ja>R�m-w{����dGq������%��e;�m�,�|�Y��NNɺ:���:κKu��7L�9�ȝb+�M�x��o?��W2�p����5y��{-�.��]b�t�+룗ы�Qc7R��=X�V�)�8��!;�4V��1��x�%�Z�z
���������w=�|s��sm��\��,^���T��@�3(���u�|�N�A�`���;�"���*�b�Ju~Uhŵ���2%P��0�Y����d�"lݺ���e���n�G��Q�cR�7j>u��.i`��?��9��b��KfZ\���*���8V��Șsn��J�#	�H3:e=��"�2.ã ��wVw�w{X�����	� xe�Υ)�j�:�MڡZ�O��_?�؄���)��V��́�����;�J���u��[)�b4��l���we<O4�A�a�Ĩ۔u#R�m�����`��_neئ(�/{�{�}�]c������ap�xy!��M9Wql���H�w�NnES���fĕ�*mt��S5�o2�z�YN[��Jm4��#�LM+]I����m���~�q.K�.v�4�J{X�u�,��W�!W)S�6�GF��J�U�����Q�`�����RB�55�r.�%��t�B�����.�Y$�2�8��|ӐWQ�"70��c�w˝ɔ6�늢<5���ú��+�� �<�p9* :���vp�#ڷ���F��Omwg�Ʈ��Ek�(8��(u��E�)R�m�(�%��㗎��a.�F�Q��7���M&_?z͐`y�$�
鉺}[u���1��#j��=�OD��/����V���Ck��دa��;_qˡ�y���'Ь�^X�ݭ뵼�0<G3�Q�Y�U�U׀&J��X[t~�� E��
��R1
,�%$�Mܽé���f��L���]1	Z��Wv�=��
�<wRO\���w<��bd%���.�ۨU�k��n�x,D�u�W��P�wq��/+2���E��c��;�Gunn�^�N��ڮ�mK
%%vg����wvE�^Q쳑�d�\�]�ʹ.��3n�]w�G�
�9�.E�=ĽH�$Ѝ�P�㺉Y�JE]��1Nu���"2�TSKU5K4L,��,����f�YJ��2�wrΐ�F�U*''t��T�Hu%�wqr�]�u!"��<S�Xj�R�T$P�[*K-iJft�n��ȭ�0*��\�2��u
�E�E	J
fQ"l�RD�!(�C�s��T))�&a���Pi��p-�������asN�TZIb(�Y�S�����9j�T.jI�Gue��A���<ܤ�,����v�N'2ͪn����-�@	?@j�)i���6n�˾��82������,�gKq3�ـ�$����XN�fD��wZ�g�+_V;����"l���u\���������,�k9H����iLe�s�(��p��MU &�x�n0�F�e�&�X쬛��1�	�Qv�.�ٶ�F+����K���`�Y>�9�D�g������������6`��ܔu�I)��:=��f�,E�!x�X��v���ꠊ��' �My|��:����%�������2�z����}���N�;��ߠ�V���y�#e�*
n����{jkqU�Fʶ�
��&
�F!��[�I�����L�Lߋ��/��¯��ȣm���,������[%�L1�鉄���W�����5*�Up���F�-~U9NS81fI�!�����"�N���j���%�C��u�d�.�����܎2��"ĪO��H�Ӳ1�Y��)$�K��A�䘰P�9	�k�+K�Q�l�y��S�vxW��f��1Z�e�[�r45�&�`�c���-�`�b
 ���8d���W����Y�+�%5ׯ+%�� ��&y��c��QɈ�[wp�\�?�1���1��s����2��v�:Ւ܎P-����a��'�cۜ`T8GƷ5KW��UŮ�;��@��R���|�"��{;�}ź�~7��}i4G�����
ݾ��N�K97[�\*L
9�Na3S�[��F�觷��t��%�]��,����9)�>��������9m߸������f���Z��LN�3�"c����V�D�ݟcYG��������TI���Q9Z2�*��6r;Us���Ϫ�����-����C�(y�qs�l����{|!%�9,C뉄.��C2f���\�Fr�b ����{,S�w�c����a����{'����Nh]�U#PV:J�ōe'}[w�F:&��=I>�u� 2�'����ъ!�1�j�a��{Z�<;�_T��u�
ܬ-�w�;��rǖ��P�q�����S�^�<�vC�cE�W�(+2#7�@��:��u9��YW���q��
���Yh��H<w�놃����7M���sN�Μ��br.�d��]�� #�����[t(�bE��B�#�!O\���o�*�tz��ljxѓ�ם	j���~�KG6b|�"���<�a�*a��[L+�5~5�G�N2�l黗D�-:ogk7##j{�귇QՎӑR�󏉤�Y���ҸyUVz`��Q�� kGd��지�~�~���b)���tm�7���\��7+λ�oU����SR�����pZ�S6�c�Q6�>��@[��Kj��(=��^N�,��ý�`���6��Jl^�]�3�e��wn�	ݣf�ε�[�%�9��A�5[���ﾪ���$�7��F^�D�U��d�V:�[Y@�d������T�kCn�g���7w][ӵ/��͚bᾫg �@G\,��"�� I�7���TNNֶ�򍝾�[�.�!Ch���u���U����H_����6���.�1 w��n48��/w�J����c��f�4��gRg!�����b���6���X��b�d�3����d�e�q�:��ӣk��Q��Ϊ+E^*`�΄T��j��]���o6�nQ.{;�P�'6��̆*z���/*r�
�����8{T�����L�r�%�ۙ��FbB������~鰩�ϐu]���������Cb�ycЦT=�6�4��ﻕ���^�K,zֺd�3��{����j놌}��^���	B���JXу#�Iwj{u~k�5xs7I��N���ܸ�p��(`��GOf�"�
ݮ��ݒ�-�c���m�ü�F�[0�<��YX[)�
�`�q�1���7Gp��Oְ{ K�����ⳗ��"��ɡ]�R�{����yL�I1�Wi��}��������D�g2�r9y1k�)IGt7�O/ ��c��ap��4B��T���v=Y�������q�!�\���o`<�I�6�t��{ޏ{��n6ҭ`a���	��b��\k7��Z8Wv6ǵ��ޡ�6�u{�#��H�����{ї�b\'��4G�IEH�T�q9g��]$Gy[�:$%j�o(��f��5˴�<�%i���;�4�5���p��٢�����*_�]� �N��G>�x�b�ڃ�,�$\B�I��"��*�*!6.��W�BFk�
���'��x_�<�m�+�s����{��C5�*!4�&��&n��y��o�ѐ��-F|�iOG{�̡�7������,���A������_!�5�m\1�\�3&Ґ:��t�XqLp4��k 
.��t�Z$!g֍���e�4Ler�71~n|��~a{Z�^絷!�;2s�>�=j������k�n�e���/G&�Qʬ�'r�(�3qZ�eCHva�u������뵐B��e#�r}Kކ�f�:���l<��}��b@G E��A9�['� l���*!����,Y�5�k�^���Ek�����V�����U$W~~�<�c5�k0�wX�Y�\v�a�Dn����Sc�ţ㱷��pl����3�l΅�!��v\�LY�tdO6��l���u�s��)����c�6�p�⤲�G6��(������t���0�]�_q�Q�V���{��m%B��3&8~��G�OS (�&�9��j��>��B�+�r��:τܫͯw9�ٸ�c8�ȗ<�)§p�2Z�:b-���K��l`�wUW�~���o��wF�`�F���gNX�q�"��b�CG����KK<�|���R �e���`眦{NxX�0M:�/#`��L-y����M��W{���p"�wŃ��xp����ƴwR�Lt����r�"[&���O���QA'+�cw�}��߄�Le��Y���"��R}S�Y7�0���p�4BYt�8�K)�gw�q ٰ�e�|)q���O^�@�ʳ�䲨����}������_-љ"o�iw�����򕶴'���]��y�]Bౙ�����tQY�BSPO �d�rcuq��j�}�7�z� �i�>�C�Y�>����rr7���h��X���.�~w�(՗s'z��﹀;q{�G8�GWi�!�w�֙�.f�n��1�86E�c��]��ɨ�}ݠ* ?j�K&�kE��*�:����W��|��O��{ވv:�n`C����:ph��@�Z���,���Arډz�E�ZO%���<�PG�r%A�8̈̓�hUQd�Sq�8��Y��
Y��*�q��ùhZy����3���L��
��&,��_5YSE�tGmnF���:�x�ơZ:I9�1O*��������ۘ�[��u�͙�'&#���R��Z=��_e��i>�H_��/�A�j�[�f�R⊘����mHnn$Ł�T<����m.���e���X���],� ������o��|��������ڠg�˰�A6 	�rx�x�7/�ls8�fG\�7V�o�+��D�Z�� ϫ*7��1��u�9b4L7U�,������U��W�Uj��g%o�<��wM���^��|Bş{6Pjg=�bK�z�r(�nN������_\�0?n���)窯���@)4h���\�LV���w:�ϫ��ʇ�EG-�g��D�Et>�ٯ�^jl\�*��6���19�t��"a�(C�B�氡y3T@�@�p����-�P��_S�P��OLd+�p�_�5�Q����1b4�L�IC�s8�X��hX���>�|��Y��P�n������������&���덑=5P�E}[|�X���^���/l��]���o�y��&r%5~����x瑎�tƉ�l�u���� ��[x=��u.�z_x�u!�݈Q[>+��YŃNv�.�6�q-[!���,TL�~�u����)�i�iع.�M�v�ɽ�O�yΤ��v����]��X.Ru���A|���:��7��������5bW:�K*��X:t�J�Fz#�����j�_]+�� v��~x�E8wǧ*`�O�B�e��;0���P��:��^	=�#�	v�u��q �O���)�
���0����S�D�t���s/�P)Ev�[�u���<�C�2�N�rP:`�*��3�w�*����a[��B%(�|栃7��y�u��H�8G%�˝��ѯ=4"�J&:G7���H��Q�����*�u玣Yw��Khkw��Ü.�A��V"�;<[w�+�y�@G������1�ו)��Yͽ�c�x(�������{7E�'C{4���<� ü�*!9" �7�s�9����T�xu.���%��E��5^�FҘ�II����mH��yw�
�$��]�������l����
uz�.q���35҃O�3��`#�T�g@���o٬��^��kU[Z5�Wp�k�g�J��aVpH���L�Ѐ�J�C#��엷�Aw�� �B1��ܫm�1���&8eD�Be��>�aY{���X�w�n�̲vЇ�'9g��(�S�"9�n��g��:7��`�g�f��Ҳ���g~��5�J���&���y*Gv�ﻨW���A��%z����VgAX\mEy�2��6�au��,��D����|b�'(�#t�jqQY��M����� k�����W��Eio=$E�G���E��N���{�+���!k���l�]����Y�R=g�7����W\��5��w�7���΂9��x��ݟ\v�dߙ�gw9��j�گG{����3���e��ȟ�`~���ѓ��J G�p�;E)��1�}0�nC�#���{�x��;�]���z&wS���a�a��Zޫ�~ɔa������ea��2�ד��J�)�r��J�r#w!��KX��:K�_5��e�)�[��~|F�S Ȃ�c�1����
g��۫��O��ث�d��̺8��w}�@���<9��]@�0��ܼrjj���j����W�pu��,3Z�c:q����FIД�I�<�a��yݙ��md=�89��H!�P�=J\��$R�]�!���r
��L��雅�f4D$n����<�{3�B�]��U��/��;�ט�MM��������� ��tE'�I�X�60�*��7Ӝ��h�4z�*wd��9 ���3^�o��.OD��:V̤'�6`��3y������[Wu%���)�ٹ�9rN���V�VU��uއn�۞���T9yQWzG�ց����E�¢%�}v�+=��9Y���}٘#"�7��9XŞf�U�V�/t�����������G��3�\M�^�$*1�}x�YހP�\�5Ϋ7���ξJ��+$�o5nJ�_<2���pX���}��D}��33�*0*��&�!����R�dc��j�)��a.��h?q��+��i׺�ރ� ��;R=�%,y�Wf�
��xS��(9Þ��'7���lg���F�a��S8��R�Z�(`�w���#�O��9)c���uku�k�+���͜�ޘ�P�[=9��`�r��'0��j��oL�J@�]rp��i��*P�t2�<o4ء�\J�y[p�%���و�mt���]�s�Ƴې��&��)��J}�^9�p�vsUHG�HXO�Z>q;=-,�K9�5y�s{у~{I�㕋�i�zn�n��;NI��v�:`�+t�����|�*�B��R����G�$.g-j�u�p׮�P�}�D�8��>5�Q���g�8e
��N��5�|L��p��¼��؜-Zz�饺v�W�������%i��r�ߕ]�TpL#�S9�k�O����5�:�.���OQ�U���Y͘U{�(�/�V���+>��W���%��:ӴT釤��l��#��$$� �U�.Bo�.emDG��D1G�=;w���R=�3tㆵQKoz�G�,^�r���R[;9�6�j�og	[���VH�L����ꯨ����O��Y<9�Ҹ�
���Q��KӹՑ�L00�y@!t�fӑ4��<��ni�ɻ�^şe�%�=����ŉ��u\��M׼���/Ԭ9����,��V����5؀˂�@�sf�����;�v�f��$�oӼ;(���o��s�	��b���D;uNJ'"Lp�9��H�0��1q���'ht
��GwsӨuek;{0�����\�suPqK'�!q[1���M*}���>c}]W@=��bڴ�f��4=���;�v
��n$��<����`-.�裮�o0���us���[�/fK�(B���CE�f��&mHx��db ��'� ��-:�v+s���[��S�zP�/�v�߳i�oLp�^��L�y��7U,�P��a���2�ȑ�"wko]|���L�����sv���W���WK�}"�w#�s(���鮙���v��V�&���绔p�B(��P�%�dЭE�����7���^�^>����<�Ct�:�mo ���8λ�`�C���"�B��Lt�֍���j�\���:k8��إ�i�C:��@���9�3�p�_z��F`Q�m���BDr%f�[/3z@�/�A�<s�''��|lo��!9�;m�7KJ����ݠF�9�qU�у��=���k98L��|����T�!>�m�{Y��ޭ\�Lf����o;K��X$��x�57[�Qr̖ѧ�:�ZG��4����`t0m�:�K��2�}m��5�� S�8�@C�#qb"����r��>��ҭ��i�V �˭YH��;����K�dD�5�n�S�=g�ϽVXr��%��ҥG�k�#)^}�mC͐1����JD��ŋ��-�����ݱ)Է�a�oq6�:m��b3�r����b�D� r�Dfm~N�(�KÚ��p\ˉ���s���wa�r�1Y�/c�ɌI蜌:-yې��)���_p5�b�����J�Qב]&Z�K�d�r}{�WG�k�>��h�S��h&,n"v�q2���&��W��t���*f�d��[┆�\w��tV+=�>6e��@b�T��3�~{���P���VА��n:��_bz� ���zG٧!}��-��֞ʘ��}5ޝJ}�0���	�]�chxA�~R��3$�S���(�o�R��I��d����E��OP���+[���qnص�֬��oV)�:a��j9b�\e�[����{>�+���Ԓ��m�_v�杁�ᱢq�q��IJ��M#N�O��Ul���Lyk��˅:�b
v�VV&4.x�'�����t||��z_��pf�R�鶫q��ӄ#Sr�IHLӇ�u�h�,صu�}(�'��&�|���;�"E"�i�Ӳ�͏V�Y9�#I��̕��
N\�����yKU����>x񹨻�p,��b�H�����.�7O`�[l����,F �_��f���C��>��Uf��|^ĔN{��ػ�D�.K6)�ɡW2����#6�G!���*3&ۖ�I�&�E�<P�b��}i�"��:r�x\j��@���~�q��Ѯp=��-j��;�Yh���u����ˡ�X�|�e�b}�'r�]�9$+P.���XPָ�iJ�u	�X�;�OAA�׶�����
{�Uo^���|�La��m���P���L����"�@�Xa·�pq�;�	�t;tt�I8s�V���z�q:�v�ǭn>�%?��N�u��>� ЅA3w�oD���������G���hc�r�<�E3�3���u�*�En-Q�ݣ��*�Ag��-�Olh���
����x�Go�޿_
`e�t�wV����#�xȣR�C�	��Ny8첷;���z瓑X*U���IJEY�!��������YR�B��꣓�FUi+��	 ��f�[����bit+���=	���D�X%ewwu!t�K*"P/q��v�fa�1:j{�p��9���ba!���%���s�7U���s�Lr����5	1jbbI.��R͚Y�#r]��TTV��snNY��'���32���iF���R�-9r9t�U���Ъ/%ښ�f;�Ȫ9҃�*f�[YR��D�41K�UF̍�Y��J�"��U�҉�q�+�2��.��K9�!�s�9f�eG"�D�UBwp�<�xz��U)�Ss�#)3eU�Xr�K���W7%0�N��*�S �T�(�NJ�`�j��r<L�5d���)NyPs��sS���P��,\ \����z
Q�M���r�/@v(�:y]��O�f�b���Y]R^��7���4�7����{�����-��f�@����)t�SL��i�G�{eR�}���&a�����������ʹe�v���J$�`IJ���aQC6���eb�;��F��t�w�����<ն9n.4n�J�BļV5M�q]wь��iP��p�wLj��Xn��܂t��J	M˔��1r�s-�YP����m�&rSW���¢5�f;*Xb�U�ӔDoe(T�1��3���KZ=ۉV���V���:|����\����{ez�M�C0�9B)]�}[
B�k&��n� ��Sڡ�\@ B�N�W�� Ve ьӣ�OQ<�$bj!\��l;<r�lH���1��������Gx��R���k o�Ç�xIi�J�Vj�鉭iŚ8�9k�w��4�޵�U�{�j
��q5�ӑR�ut���:Ы��k�m�,��h��='���B*,�
��@w��0\@,�������=����j��\�V��y��i��l����������-��
 v�x,��s��]��<K������xl����h7F�s�K����fu=��FcMjkׇ�,�j�2(�ݪA!�ޓ�]���"Y�b�c�ޛh����k�IVN�C��z�._t&���zODm�h���Ѓ��/�Jq��n^f��I�(mlo�u�x.u�g��g����}U�UT���n.Vˋ�3>3�6�H��Z��Z^�F�)��Ԉ�N���͉yu���{m�o7E9Q���p$=8N����Hc�ו��g���WJ�]����*k.�,�����[��W��wh��tmp�5vy���K��S����W�!7_�P8}:i�*��7��4���)������Oi��2�*�YluҰG��.���QGѽ����]�?b�)�nH�'����F���[���a����{�n�n���t���$�yygFH�q��(���T,tɸ�cƧ��G���[�>�0@� I�X������w�%���S62����㔢��6����ҡ����ۦ����0�Ɏ���Sͻ����v�}^@ �Ѡ�H�w
�&Q�/�f7);�A�g���F�BZaL	z��N�����8�suʯ��@--b�����9V�p��,���~znK���u�9�vq���l#�n���[�p�Fj�TF�3q�2�᤿���)T��Y�b!�[>��6n���Z�I�G�ӖV����r-�sdp�2g�lʸ��um�J����5��`�T�t��%ɤ咚��W{q���îej[4\G,�y�;�m��c]�j�u�o�Yf���	s�b��t�V�9�L���DDu�k]�>{��D}��;�w���ӹ��>n�C��LW�y"��z�R���[�<������m,�:�\p�J�w���1q�@�^�Ȧ雅��cL��j@����īKb��4(��ÐKGw�1I�q7���c����o��
;�����9#����Xb+�
�S�p ��<J�^��y��`3|\�^]F��Η�6>/�m�q]�S��7�
��W1Ց���#��?*�W�ZW��5w�\lɔ�ê��'���i�=0�|�Şv=uA�K�����5����vڨ��&�&i�N��5RąA.�����ND��k+���V�=���:ǿ{h�B��	�Mo������[ڷF�nAE�j�n2��&�jfV���>n����O����W��O+�O��j=Ӡ��o���VR��x<�S��+�:�2S0���3zdRRє"��{t�=<����1^ �@��%��jJY�8~ǕK���[?t���Z��?�?��=�=��6��'��\];c:v��;�L�Ŵ�f��&u润�C���.�}�N��K��6TCz�g�Q�%�� �I�w%)�&�W8F�-P1��	�l U5ݠ�N��\��/�"k{h��Vz=}���I(+��G���4��w�q_{gh�舻3���q;=3^U>�C�3�����0sj��q7췩E�6P��=H=ݟyJ�7R��a�pׇ�_y_�#��6��jhS��rr:ޥ-�i�G�	�|wa�>7k�2���g�8L|zfP����<���q�{��q`��ٻA<�Kꙝj��g1F���r�oi��T���8�o�7������� �h
�/�y:=�[ڇЋ�B�1ı���`hn��RQ彁�Xs��J�g��J�HY,�T��`6x�\^�u�F�ħɕ��
�>3��7v�7��7��2K��Z��U *�@K&�`��.b@E�v��L�cn�ngBeT
��9Mu��$��}�7_X��7��>�"�ʕ"�
��
�� ���j��D(�u���EAf�C�]�-7��.	��֦�U3��t�w��@�EqW7^�,��]Q#N'�FaR��u�ov��k��Hm������gTNI��u zc���2���M�.��Y2���7����hn����G&q1[��vgJ
h�AΩE��{,]֫:�.�%��7����9��sʙ������@���j�KzM�K���c�)y.u�]�0�?��+�].�4��YK�����P]�K+:f�=�G앨��� ��X�Q:|kGٹ�1u��UW��V�yȻ��6���*MF�o�L`���������H� �O6�M�vC�5���+ڻϸ�Z^���I��~O}s*\ل�7�hbUR�9��[��c�����:f�f��Sم.k/`!��0�²D1]�`w읭�͔>S9��!0�:�Q0���U����]n��xz��ߍT8�0p�~�\�u��n�M��T9΢��x۩r�gs���*2���.����� �K�D*�+�k���vxY5��-Aʾڙr����Z2H�bYc�M1 [R�ū�~o/�c[e�f	Hߤň�a3N��Ĩ�n��]�?)W�߾���}���C�F2���:��鍵W~�p�
��A��=��\�Z��Nz�__�k��ޕ�
�s*�m�&Jj��Xxn1�c��)Wu�[��*xOC��jiu����@8�.�b�CQ�Ȭ�Ǔꆑt���3	8"z^�]3�#�g9.�R*�q��)�(�@i5y���
���5+���h��ϓ�8�$�{DFFmv����u�ߗ�ᆳ�oɫ�W1�f%V�J��-�7ґ�.
�1��7��;J�? ���Z��w�9����-o�9fCp�Ф�$T�!�Xm��Q�V��+t��L=���u��j]W�}�kS�9-�0�<d��;��U��}�V���\�����1�%��g�;�P��˒�D+��T���Z�'|v���^VP�[��l���n��μ[Cm~)mC�G��7�O+��=i��wY�����V��F�o��b�dx<�7��į4{�#���������GA�ހ�d`�#I\t���Jye���
��pLMk��q�ݾ5EF���Ȅ�]j@�PP�TD7�Ȩ�\b�$f���'B��T)�Z3�l�ǵ�w�{D��4T%$F.u4u�@4eӸ�O���7��w�F�5��I3�{,��HC�ו�W���CL��J����T9�50��u�M���#
�ԢD��ʎ�����yG�Q�+�T����.pP���ť�6��ʭ.}� ���B��n8F{��5r�U�{gLs��,���^�'w.z�MW���JoL���qX��,b[�3�˭�
f��g��m�w��U���9&���+�q���s�ǹ�!Z���X�.�g�\�T3��G;����E{����M�Wgv��r;��t$��A�V����$����G�hL�ܸv"��I^�\�!��R�(�=�<7�E�*��b���KWb������wQ�ݑ��6�؋��'T�\�Nl��v�-x�4r�ǮJr:a�Θ�LͷoL�I���{��DU^s��2�=<���<0���,,U^ȳ�DܱȞ*�gF�o��aڌw�ǜ\���[3�;�2�����\�ȍ�$L��H�P��2�0��eD�U����=�ն�:y��<�&{N�V4,5=Y·��ZZ�y�� ���6tp����<MY��Gе��p���M�޹�gF�z��/MZ�y�#�c���@��wB��C���o��1�OyB���]g���ٞ���dgs�X�p��t�7H��%�1�d���}���A-h/�eK�ӛ��	
�wm�`��BƺU"��n����=Ĉ�f�f��d5ٍV�1��n����]��R;��y��i\M˨L�S��u�̸u�Y�c���x��]��(2���"��Aנ��S�sL�%iLk{P��ȗ83%iVf�N�-=%ľ���'Y��Ϧai��O;m�����xYrj����bɄ�V��\s�>7�Sa߂�$�D��#30�eFe��������j�o���3�.{�9oY�7Wf�I���oM���u$;��Ww�m�3pp���^�~�N<�e*�w��z79��lJ�L;ʳ՛��]���>�a��)q4s+u�n`UvP��`]���}G�G����;�iK����(�^�m�Y,2ƶ�I��Y^v�k���NϞ�,�mo�
���g�|�l�F��꩕�m'�0�S��Tݵ%p�k�n�o�`����=T�T��rl��7R��F?m�j>�9�;�)�p�����I<��Vp5գ��Ր��a`�샎�.s�q����=��lT<źGp��˭U;�w2\���s�Ս^��߇{Y=�i�qG+�:�7.�KqFMUt�9k��r�T׼ڮ=!�Ǟ�ˇnGC���Ρ��v�B�>� ��ng9���6- �uF���;{^S]�p�>�������݀!d�i��%����7���S�N�|�4���fsoj�Sq�+mB��+xf^ɒy?4�S>�>�%��F���V��)�p��W��5)�9�w�[z�US�������*�3�	p�[��5t�O��}���(x@�u�ǃ�pN��4���!��sh�^��h�ʼ��,e�m̠qV�h^����Z�]���YV���`�C�u���<�ske��658�8Wu:���fi�]�v�d�h�z�)>�J�l�Px��a|��E���K����KI����JP�舏����w��G}����U�Kj%\a>���.�;S�n5%A��Z�e<;9ѕ�l�~K�U���	M;�����חf7;�j�p�����m���j�s���3�]�7C!1�J��=�nc���g�M9է�5��ˇ��g���AV�wW�>�spf!���0V�R�/���'3^�_E���l���֜x�W=����RU6���t������&o������YF����W�k5p5ܞ���q�k�s��3r�4D���}�j;���v������|�ťw��uLB�n'!%w�C{�078?b���������z-�����US�U��'�dJ��Js�	��a<z:�������;&>�8���ܶk��[���5�8e�Ό��s�kb�'���v���}bJ&���ۖ׷3����A�1�y�3�`vi	���%ײD<��u�!��n_^�t��R��%{}bu�'Vo�F��9*���b�����)��js�P�$�ݥ��f'կ�/`�_1s�vm<f���TX�b3���ɋ�B�)B������p�������2O<<��ˌM��\n>}G�*�� u%�Ԑz�r-�7;�ы�[��8��u�T-���Cw��wg����k{\"��jVsP	\������u��Rb��*X�U�|�4��F�j�}d�=C��Z�ތv����F�g`%¢�YkGD걛�v�GZ�(�Z��e�Ե�bQ�2i�VͲ�w;�삧����pՏ I����l���9�%Kdj�m�W�q��-ؚR�]�z*y)��pޞ����M;�o(�����Biu����n㟭ؤY� ��k�oR�2s)��^�b����$��3�_SaC��J;늸���I���n�O�W�h@=y�Kk׃��Ŏj;��Tr�3W�\��l�_N�W�213�[~���:�u�^Z��U�����/��{[��+��-�hpL�h��ʅtm
iJP�.d�,f�,�@{+�eǔ�,���>1����wO����m	��1��TlHu�G�I���B��y�����r�aR�2�M�ō��i�F��w��N�V=ۃ�̍z�q_gu~/�R��z����_���:���tu�ܻ��ꁸ1� �ɂl��`~[׎�X�~�IǮ%|"9�9FV|��Oc��J1K���ڕ��;B�d�kb�t��Yh�@F��p�塉�w�Rm�H�#�`����]մ����Ey99��":���Z�.Ք6�Z�4���d�����C�L����=��&��ގ�.����A*����� �F`B�X�5��ݫ�����Q�i$B7���+��[[>]zv��B��kh^��Vf\;�!��#l�a{w4M-�"J��t{#�Π��-)��FI)�5�`��*�M]8�J�x�:w���N�n�ԐK�֍E���{c�k��,g��G����<�[�.��H��Tw�0<��}�nN�h��x��dNL{�����eei׭^>�;"���n�n������>�����Cv����z����Wn�v���[�eM��|�",�7��ޔ��������KW�W�S-�je�©ڹH`Gy�˟aF�uP;�Uo��}�H�r��=ɔ��i][��w}�0�[PgR5p#���;���Uۘ������Ww��-�9���Y�7H4ˉ`[��M;�sSr�KQ,a�E����#4	Ũ��l�����m-�8a��صQ�� Ȗ�1��������I^Ç�-�ޮOj}�&���E��V�x�]%T�Q����]���s�+*��w�`0Ɨm]6����E��⹜'�4(�v(�!X�u����!�-�7�z%�W,.o0L����Ę���u�Zؕt�6+&��+^�L��5��Y���˱w��EU��"\���R⯽>88�Jc��I���+�,��uy�rD쵡 /.�[�L_ϓ���2n�9��2]�8��I��+@�2���[���0GT�@u��E��k/;!���Z�Ty'Jȹ�@��bִ�S7r���vb|��t�2���s�x+0�|��]�\7�hC��n2h�٭4�$�k�w"Y�-S�K*A���$�T�]�%Xi3۰t��:�ۊ_$7v�<����{Bһy�7��s#:SN�]vE+�L��sV*�(8j�2�� ��JN�;����/X�&�B�A��>K���x�uő�Hv>x��wrHB�[��*����:g�{�$�U�x���w����i<݅��
��^��sۤԱ`be�;F�<yf�iT���d�ثjZ;8>ͺO����f�
6����y��������܉u�r�e���5�Vw�J���)a��� �JȲ��a%��VB.f�ic�s���.v��!�����N�{��u6�;o��]}�(�C��+O �뎞I���)�e#|�<=���]@�Y�,��V˞����	������y�nn�;�2�D��J6����+�i��^d�Z��diEn���C�<��fJ���ZG�+�9�A��zU�����9ȫ4U�<I�'H������U(���N��9u	(*���]ЏM	���$�UrO)e������鸮Q^�Tz㋊jH��!8d�^��e	Ԍ-Ve�]B��ӭP�\�e:����燢RFV�B�CJ�==\�R]�,SN�&�Kf�wg���]ҫ�꒒�HE����V�U�
�h;��&�����J���p/2��h{����Ďm:䜽B1Z"@��!�"J�(���儺8:&�t��H$ʰ�.���w��fb�P����I]#�<Rs����4+�](��V�*�*J
�"��n㜏*sćB<��I	L��"CZrL�$詹}�"�� �lM\�J]\�y�Ď;:x�eJ=���|C�糗��3I� �x;jԘ��b��'��
�n�D�_�����U����T���v_�����,��K:�p�B��y���d�ܰ�O���{�����:ݾ�]1{�s���SM���7+�vQ�b��a�0�|������u��)�kϩ�������>�~�7�{!��J��=�x�՚������w���i�mz�p~ԣA��y�oCW�=Vw��۾���k�a�cj[��Ug�ˢ��M���^�9~J�}��OG�ܧe��ў}��d�/�Ԩ1Z�E�Ml�5ʌ���2s��o�A���;�L�>��K}]���|�ʄσ����=j��>I°y����c�~�܍/W6}�4e��酪�ŗ��lcv��u��nHp�ksw�[٨<�M����Ҕ덳�#��/Ex{'pPȩ�Q�aK���?D��޻�ߖ��W�(���{å}~�Oψ��BV;˜��j�B˥(��R�3�K|��ZW�g$ʱ�L�8}�q��x*ޠ+u����LdZ�Yv_��sL#�ŵxwy�>�h�M̝��>C|���J2�'%�vq0`���^�Puib2�wv�Oc
gj�y�Bl�1�[�3{K����z#�BIv�o	�;�Y�nb�ak�]w�Sq��z�'z��ao���A�Qr�p���Ӽ<=w�:��p��x̾++ܙ�w�p�7Vvν�:��qq�e�uCv�8L�F�ע�S�gر� Q��xru���?-w;ɉ��P�.�:�hm\AZĮ��Sdؘ�4�.�*�VY.���{Σ�Pԕ^mA�k)�`LF����uR��O,T����{�}�S�n:7�n5p5�2;��~�����Z5p�SD7u���N��/��Q�x1�<Uf�ݩ�g8�YM���p��3~j�)�'=�:��M�{3ͫ]�/<]�����:������cc�v��9�1��x{zoR
\.i&�;��]^_n���e��(��C~to�y�x��[��J��m>�b��{��v��;'�ƺ�n�=:]E�*׈I;a01��7N�JJ�iN_P�N�ڃkܩQ��ʮ�{��\E��{h#�w�:��ě�Q�đ�Iw(�֮�7�����6���)L��Y}���#��a�ԏc�<+b��!���ŗƁ��'�D���y*!%�C&jk+��Y�ɻ:�L������f�I��^=-�c%o�{���5��kq��J�nC�}y��0`OKc�H�)U�Wb��O���;��N�e&�[��v�{^�;8��ެ�]KC��(���ms���N�|3��e�4���R�ȍŻx�%"4=&�{��8K���8cy�J2�s>	p���-h�]���`����}��gi��8YMV؋x��1������xZ�D��F�6ks��ۗV�u� ��{��gTbբ��;�CW�(w��zO��n:5�_S�~]��W�m(u}J�]�{7W��M�e?s|��;�9��wMؘLp���-�+��E�����pa��n�Ȏ{�9�-����9:v��yd;�4&93�⭽��)v��˭�켷��Zg����{ܨ:�6�p��U�"��蚮��t4m��˚������'yko�������=��ө�jŏ��c��庍\"���V�J0��T�ψ��ͭt�츮��vK���*��?s����F���G���72�nb��(Gi���N��i��&���XD�k͏(��'#ɍ��&��b�YF�MऒYYx��fj�~�����Ҥ7]9j�۪��;_�Y~?,�8����ߘ�)�=g�K�����;m,f�f�9=�j�2�~�+S�ˡ�.;G�>��s�u`��UͶ�[�;+�ģV��`k1��饸6�:�ex�}q*�T�0�&yn�(��ԕQ�1�s��͋Ze�7��mD=��v;��۝�t\!so!���g��։s�6�X��r�S{�������;{Jk��� 3S�4vt���GIBS�8:;��D�Y���.��Z[��uZ������
r�ۉ~���h�p7 �k*
Lu�T��W'�S��vgo"�ݴk����=�w�e�l%�loT��x%¢�Y%m:���IeI�z��[ݭ=ٴ�i[�i�Bz���'�����/�]���ɚ���^̻\������V�!���y�g�v��	���o��k+��KΚ�{J��X���*ZʝE؛�	��.�=�_�z;L�W[�h�~���.'Ƶ��2b�=���;#��Q��/YJ��;[�+2���2�"e�R+v	�Gf^����[�Ȏ�V�Szv����u��(�H��ĸ���^��A}4����z%~���D��<y5���X����.8��[�-+p���S�sf�UG\�<��r�m&��C(�	`��A�ܚ���n8��$��7��{{j��u�!z��I��ʞ�3w�\��y�j��A��g,��G}�߼����4�ӯu�k�M- �!���Jm�~+�+���u�&�߷��i�R���&w|�]�9�6_\��`]�f�P�?�~s��޸�pOQs�lE�8�R�F��q��e�üʍcr��-�U�|�*N�=��&���rս����Ka<��n���[� �gb�A��]܋���W�+�j������]K�t���=�?yy�<�M�s3\�2/wϦu).Ԟ�\;p�m�Oa��Btm�:�-5��GMO(�ǟ(jт�w{�[����+���L�����C_�j�J�}�Zn>���aZ�v�ri�z�<"eޅ7jݎɹ"���9^آg�z�mb�;�;�p3 �c4�il�8���+�T��ꃴ��NĦ�p�7Mwn�ܻxQ眒ӹ�xp�q�,�5e"�Y�z�����5[����2ϲ��!�#�����ꍪ{�|- *��qՖ��ݞoQX^A�;�Ҡ��� ��EYw��v[�9X�g6�|�Yx�n�6�ox��z�2�ӝ��c^Ғ�YZny8�离ɩ�/����`ԭ��ic��~Ɔל��Y@\Wt��I��cTD���\.u�qU�v�>��B�� �x@.�%����}ݠ+0�0� CYF���Z� .���&��/S���U�+r_��wն;8�����b}JQ�ev׌/�"��[�a<������V��^��9�=$�߽��56�ހ.�Џf���Ó�.�n]�"V��^2��\n��=�0��j�rf[�zʷP<��x�tit��b� �M*KvW=H�<}ڝ{���T�&�m%.��&1�r�[��䛓g:鼤�u����^gU���|^��%M�CRWq�ѣ�}�x���>��N���C`�7��=�9��z���`�)X� r>���H�%K�"b�R�c]��mb�ܳ��kz�1��jY�pK���Tk�����Vvw�E>���U�R�'�>|@��_
i�홝�ɷB]q��Ո�����A�VO;���� ����
���P����]�e�W��v��9��tн��
��m�U��ڵ5��mӝk)c�͗»�t�A�{G�>��u/�w��ڕ��O:���7��8�Ż�Ϻ�_M=��C/
6�'��.��z|��'Dmx�Mw��ihɉ�ZW���|��'���[~w�t;����Pj�$�b�y��U��5�8��9\��U+����C���S]��pҡ0�V�K�L[ѮF%����½|��O������ȍz�����W���8mM9����]�s�265T��
�����OZ+qٖ���pm�kL�Zs���"-���p���BR6��f}W�/~��y����� ~4Nm�%�軗}:�;UՊN^>�x72���g~޾�]��_��T;n/j�]�8��m��ŵ����Y�`��b��b&�(�ح���b��@S���}򺝷��D�	�Ɋ�����k�Su�P[���Z�Τ�=�:#�<�a�Іܱ�k6��`Ѱ�X�xQY�]��OmJl8�h�ϊ�R3���]YϜ�+/�%^�;BL�K��ޓ�i��X�rv�C��.�;h��z=�ӼԲ���7s_�/ϥm����Ӱ��py�+us�� ������Ӎ�<ٳ�L��Y"��I��v����\���W��-�dU�۹��݁�<s�7}!��j�AŴ62�g���پ\��-�v�Rچ��7wM�k���כ�
5PSNX�]x���w��׏k5p5z�7vԩ���Q�6):�]�9�)@Cx8͍�wN����W�-ex㽣�{Jťw�%b�zuH�Ӭ�$�_9Ā�q�X��Z;�,���j��s��h\v�⛟�O�]�Om�|�l��(�Qz�k��بy�E�{���V�ޡv=�bx�����<�-�輅{��*_X�-ť��ߡkb�'���u��my��.)'�]�o�vw5�S7cjyϯ������e_�NTbkn�ې��h�&�5��+�z��j7��_�����z|V�P}:�E�T����;���2k�ժ%�A<6l�ת�M?l3�:y��	ܮ�ՁQ-4��Yj�D�u� �0S���y�Ww���=��h��w��6��{�,x��P�)�Q�k�q�#�R1Z��:�M������Ǉ(<!B�o�=��u�H��-|�5:�|*G�%�������p�^���K>���	U��u��Pxlk�Pe&/��,��F�9�p�S�=Y4��q2uX�[.�N_E��e=�a+����8<+�^���ْnjV��s�K�ˇK�٨�ҽqگdӤ��e\Kh�v-���|�k��7��jUnq<ڨ�jMy�%~4+p�:��	��G��!P�i9��mU�ݚ�g���]�q�4���[��[y
sr�D-��yM�@z��!G�* ��b�V���}��L��m]�9�#�ӪУ���/��r6��-���Kj/O��e.^͓�Zx���-jr\>����}e]8T{��+]]W����֖Tް�-�[Own�����]��6�9�=~ה� U�c
��vW�'u��9Y}B�̀y����vV�S�x�7�5*nڜ\29��C۩n�汹z��HP�Ou��Z_q��+z�������b�s��.|�!��g2�����AJu�Z�yvr��1�L�\o8�ݼ'�l�:�d���b�+��v���<3}eO��=ko����nx͆<<GC���'	;Y�J=��Y�xg����������u��;����b��O�s��M��|��[vuz�b�L\f�f��}Z��a���w78�������[-�x_&M�Я*�z���ԎN�-�����~m��=�ojX=�GӴ>��WG
sV�+��a/�t8��u���>܈��P��{�z� ��\4��V��DN�I����vn4Kk�|�{;�΍�煬�m>��
k�n5B������u-]���]wI�d�}(~�o���ܻO�z4���({�ۍ��m���z�9*n���:�!!>oi�b�nZ��k��of��W�;w^�7M���SCW�$օ��j�YO�9��Q=3�]�\��h�X������'C/_]NB��]��3V���9eX���%5�0���8&�q�{n��Q�R޲�P;{Hk��E��R���j&�z
컃�w�)���N�I�ݱ���/_En����{r�g���)&�b&%�s�C�빼�s���%��K��=�a;�_��Y+�mc3��]�Cct��]ŉ
�޴An�&��mB�Xw��Ǟ�Y�>�=����r[o�Q70�F��\uC��4g9�]�Q���K|�@9V����</nF�'+�^�����Ym�d�����
TU�۬�t�ӕ5�ư�N+����{4��wr���*:�f�,HLu�^���܁�|���R�*1I5�^su�
�F�2�kh��&�f���ʻ��̇Gӆb��	�Rδ���0�q�ha����՝�'��.�tK~�b醥�}'.oFZ�b�T�<���eQ��ڄ�D�I�}W��%q ��_.���q'��^��j��L���<w��>6�h��G,\Lf�w�^̗U�h0��a������)��I�[�xy���2�h���Dm�}��3!�2�~񃣥�uH�{��'�w�'c)�Xy]�U!�:��s�f�������3"�:�솕�L,P���^g��*ZT�|1�'^8);��w��*xz��<56򑖋Z-a��_rۼ��Is�dPAVm<��n�_f�ӂWh_9W21�M4�%m�0��}(�5�C���jXp(N�eo8�O���0���4�'e�Nj�ž���-a��<�Y��{�Es=�����ӌ�ѝ�m�[�㐺��x����U����윴űܭ�er��q疩 p�,a��ר:x�E������J���Vi%������)%t��&ݹ[�^�g�n��b�˾f�����8e�����z��x{���<oN�wL��t5Vu͉�X9�
�[����0qs���]s̼�/Lu�Ak����L�;�L-@r���;�*U��{��u^�[b�k�΅�=���x-bJݸMb/�4���U�ڧ^�^Σ�Y�	g������_�9�2�˱﷙��R@pqb<�l�w(�}d�8`nX���S����|^D����K{�|�˧�5��+U��%xz�O�.8s�7���z��+/&��tw�٭�ϒl.��F�:����k�5+ΩN����ʰ�t-���5����o����+�YՑ�3�V��In���c�}���I���}�&M�<�p�KY�3>4umuj���uҚ��n��^%Z7U`t�M�_]ҬN�l�mh��3��${�r��2p�ib%'8��j� s�����Ndta^M	m=���`��t#[�46���C�&���
�R6ͮ�mv��ݱ&��Ԥ �fn��jb�.�X�Sݖ�Er���3<��h�hٱb�1l-��*c"����:9��k���Y�a�I�MCis��%�{�v �w�v�٦9,C-��E�t�M�
5�ck��n�gJ�����ZJє.ތ��s���J
 �9LX�L!�Q(�;��d�������PA���#&�[��^����GtB��Y�Q����EI�H[K2����Y%E	�2GP�Uw\���p��RÉek�^`�j)e�S�����D*Q���W,"��z�*������P�$
�%�p痩��*�6iZa�TFEbrNFee�3P�R*�J!�e��I�����,��sM)
�Ȋ,Ȉ��WԈ�֜��J�f��VK)�Ҽed���ꙩ"m;H�ER�*��KR,Ô*!Yf��,�|q��>zy�\�,�HTχ��V��*��Qd^�ڨ�E�\��i�QYQs<��;�!*p4���Qe\��f׈8ꪖi��\�Q�Z$ѢE	&����t��[)�sj����lagF�=�7�uմ��,��1��ju�G�g���6���p��Z] �Ty��}UK<Tپ�x����b]K��J;a�S'�oQ�����.�tn����{�����g�������jOB�&9�+^ͱ����lR`mۺ����{�;�X��:��A�5%T7�'���p.����A�Q(�.���g�j��E.�^=�����	KX�K�z�fd�1�y�}{���\�]�Z2�}�ս[�X��>���r�z�����(�R܏$���z�i=���I6c�w#;�����=�qF:�:s(T9wQ��%TgBm4���K[�_M=��c2���'����q�S���xs+�M��N����6*'��3[���u]���V4=���Q:	��t=��FV㳜�r�R����[�ܩ��o�ؕQ�+�sUU(iOn4b����;;�W���YI�O��o/-ۆޏ���c+
�;{j��J�+b��yf��^s�^��@6i[=ö�4�^���D��şw�Y82ȸ��*���,6�˫��x�C��V{�Sq3+�r�>�A�!B���Z�EG���dF��G\��뿻�>}��!d!@���	�4�A_������l[����S��L��e\J\39����q]�z��Z,$��[�(��K(WS�ݨ�N����U��u�<��/OO#�;�m��Ǭ���	k�\^�w_���~�4��rʸ��K=]3��R_��NK�����n]��9�3�w��=Mz'�,��q��#��
,n��(�El�t�o�6d�ӿo&�_rG��g{��d�ps!�v�bS,p��K]gl>ޖ����ޚe�΋����Ԝm��d��^t��Owo ���[h>��@?-L�J���uzޙŎW<Ԩ��5%��ѳ �|)ձ�%�|FF&r�o���C�����u��To��z"�7njF�]�۳�f�4�Z7����P|1��j]_;��r#ܴ/��H1K1�ܚ�f!��uJ��tm��%e7p���&��q�=h��~�xv��D�:�����#�_��Z/Q�0�I�Gw���x�\�:��6o9}�rk�;�P�b���ޙO�75/N0h���O���83_��<�S;X���aW��u�@�Gg#�����|楹C�����t%�cK֗|���}*ӻ��#Rt+z_��֠lmr|{.�g��U}VK��k�7�t�D�5�8ɈX�Yo��ݸk�Fh��I�I�*�׆�si͞���k}���4���\~��g�b��{�
�j!��Λ�r+�����\2�9�d7�,e�ږ��Ԫ�'q�q�'�Ǽ���R�BkU�}��$���R&޺���W�אz`��^�ӭU�Ke>��8�s�Q�b򲹅��b+k}Ξt)�W���Pz|v5Ԩ>�����PI����W%�v����~�{K2�bsM��L%��#z�%̝����Bζ��V�F\�ڻ-��}��ɥq�;U㌚t���ey,�{�.��[��_(�֏\�e\|MU�x������MAz�᧨<��^�c6��q�9@웭�y��:��f���J�y�v�@N|�s�/��@wÊ�=�Bf�U�f7�KM�s޷Z�ts���WmA����k6�y��A�{������kiPe�^�ןx���B=����ЧI2��i�}j���1�:�/*r��w[�P���Z�g�
*6��
/��l���������z�# �,��1C7�^�)���e��W�T���;���N����;~�琭ՉLp{ ������<*��ɧN[а��8��T[��Vݎܩ�����yU�>�*� 3��X��y��A#3��Rw��9r�JI{���9]������u���X��:�
� ���­�5����q��w/�b�*u��	e����Zڞ���x3�@��@C��5F+��L����ϡX�Q����ae6ţ���=w��1�?���I��N8���7peB��>�Wg�3j-(\�o{�Ws��G�eY�%e���=RzmN�|ս�n+�{(��k΁��U��\�y8��=v�z�O3�ޏړ�����EW/��Y�5��j��U�.ƥ���}^�E����3��C�-�M-�1J��p[^�;'�_:�"���#�U}kWǢ�h�I����>|��p�m�����6�J��1� D���Y�.�Ñ���f�{2�b�o2Rk�Q5����v7ufR�Û��t^�ڎ�o�yfg$�k�:�{y�g��M�c�>٧58�N���1LC~F
��PF�	��D�9��Nq��W��S��ɼ47�៽�DA�כһ1����ډ٘��
�k.��KU����8וi���K�Gv��A-��Y��X~K bU�#�]�.wp�r���/���qD߭ѷiGm%[c�c�팟R�j�U�C[F�6���/�}ZZ�CR������zYǭ��
څ4]�G�WuA����V���]w�
�����sç�n�ߪ{�k��;�!Tv�`&8d�%l�Fh��5�n�����[�peQQ�W�'m�&gb�c�+@�Co��5�;89�8�X��g����y�V��b�f;S�r��%o�Pv��bq�y�W�.��Ko` ஠�ʃ���*�ǵ���Q�R�5% ^��HY�Kn6�)��A�q�/M2���w��v���m�j>���i��yy)��Ty�a)wߣ~�{�ey�N��[�`��to����k?WY^B���W������o<=%��!�P3���-�4-_���튐��[��������et�q�H�0�6_���an�9�N1EN!q��,=.�n�������)����wa�w����q��{�W;�1T�31��KW\l����x�=|�j�Z6aw�KV��y��oy��=���3* �y�I5Y��"�qc��gEN8�-Q���ˎM���w��K�ڡ���@P���iS���k8�(��b��;H^�Y:|5R�-e��ny���=�-d[8l�n��$����vJ�5��w���JtSա;�p�cgR<�m��z��٪D�SI�Ab�P��Q(ĥ¯�˅��=c�ݶ<�<p��7}+�nEVt�u+���]�20D�#T���9.����	2��⣍�gv�Bf[������u^8ɧH�y�K+��WM�{jr��L���3Oe
V�j�y�]�oS�[H��í��q��؟R�xY]�Sڈ�ا��ќ̶V��Ŭ'�e�ٗVWrmc�SP���.㩻i��J�������2���a�k*v���8�f���e{��a�{�z�i�Q�>bkn�⁭��yrt�ݳ�|�*V�c�˸�BB��prD?eٱM��!������k
����;o`d\�_RŽ�E�u����p�ҁҷ���R=�zt��0�2�F\�n>��%srrХv\�P�+�ՙ�)u=Yb*��w������T�8������2�]��N\��"<V��1�*�E�����v��Ko/�ޜX�W=�H�,s��{tnR�����g���Ru	�K�@_���os��U�j3W6[�Ǵf�����u�M��v�ن���u��5zq�z�Ǜ�MM��V��5;�Bs^)��Y��󂮚�����޽=��o�����!�O�K����Wv@�f=����E����3�j��C�Z/��{U�fo5o2l==3�>;'E�w���"�.q�ǧbG�gF���w�	�A�ˠ�	������{=K�-��T�&��m�w��D.�ų�P}���sx��*z�D�Zq�,= �O��)��ou� ���kҢu����i>���xĩ�9�.��u�ݿq|�#��]-��U��C�@܈=�TJL\�޸�8+��O�y�5j���{=����/Bݸƶ��7]���o����U�'Y�o�����[�P��o|���j��P�z�Z��գUb,��w�b��{}onnpڔ�Yp��T)�3�w�����b�C:��y���b�|0��͢%��IV��YVr1NX��*�y��K�g��LhWY�ȏ9�B��S����s�{��Ƴ���{�Ns�ޟ+��&��as��P�&)��4c������˟WH�v�G�7�Z�/ބ�.wp��x��z���
��*�k��BÝs�V�c��~�ï�Pc��+^_�����ZKX4XG,\e�X�u:�����k�::↞�	n�t�\�o�9�K�ك��� 8������*������~�[]a�|Gl7`&8d�Pk��W7�.ʛ�G��4�=��ɽӎ3V�'�;~LL�6������`O���+]]��bc��G<����J�/�/s���`3�߾�r�w椪z��r��u�u�:(!��lQ��iE�����D^NW��F�%M��֎q��M앩��DT�=�M*��.9��=�GսUٵ��E뉎�l_��ò�b{ܢ�N�?JL~���ꨋ͍ZچҨ.�Ys���Qk|���	"��}��Gx�,OO(E%�	��۫��n.�3�X;n�&�,�nn�9Iu�	�wdi�S[̹�0�[<yC�W��l�"o�z5^(�CfB\t����t��kb醭,�9nn�c0�@�,rU�w� u�p\�*��c��{z�ܿSK��-����D�[C��<��곍��:����kQ���Rj0��;�+�z�=��y�͇�;� ���jTu��fz��|�v�-�C��9y�c����[i�c��
U����אyܖ�ɮs|��[Q��7W!W�W�e�h��e���mf��j�46�h
����w���.]�0o8�ccVK�K�sV��ϸ���{��Tm��a�ʷP�#��l�*�%#R<n>�����h�ŝ2��U�[���0i-���^C[�}.���~�נ�S]0��ُ#���٫�����ƻ�ݭ\�j5�v���z݈��Hp�+��'\_*ڊ��G�淲��k����{��y2�WOq2��B���&4�Ԉ���l���y��U�V�\vǏo���r������>�n�P�]���G��.��9֣r,�f��AU���v�.��svΩ� �yJՙ�f����:��!��:��swQ�̘+��[3�Y��oқ:�����SݘGS�����l̨��p�;����	}�n�3n.�x�]��:������� N�np�������V�{�t��KJ\p�ܵ��N{Czm����=z�����֜�f�"�4�_\Q�]+��gn�����eU=�R⼊�(����{.�˭����0M���,�;��F�G;��kV��EvQ�u�z�ד��駵�vî�h̽���ra��ޱ���ֵ�ΥB��fO+�������G{}��=�5��3�#6�s�Zبy�w<�sUӱpmDu��m�vf���Ȏ��Ǿ��`U�9sy�h{��uy���7v��	V-i��\�	ex#p:5���$�'+���J��}��oK����DjZ��q��K���VA��{ƢT�b��*Kl���io+I�1�b�]�ڬ.���r��W�ƅ��P�B�u�Gҗ
��h�uk�*��e����39;o��x�n�����������ݣ�Vb�.M���ڛBV�#|P]�V�p+�r�]4��C�Ts.�{41��ղ�|��˃zyM�sr���nE����\׭dk)�6�$�,	��"A�8��ׄh"E�S����|#���wu��*M��P���+���y��$�����K/���krD��wX�n͈��LT(� ���z�*���vkG���:/65Pj����j�ni]�{0�g)$�L�ɻ��wJ�)�2e�	����L��k%Z՚c�:5�=̻{�x��o)���ڜ�j���D���m�pD�����jy�݆��j�i�5�e�4 �DtiP���ɹe���hE6�<�
���c�B�b�ox��є��)}��w3��C��ϔ�Ƅܥy���#��J�a�y��\N��h�(1J]�a��\��{}6�N�+ܨԃ�P�a�׫b)&gVq e=>읏o#�Z'O�68(��R�L�0�Ffά����	���M�|�X}wkN}}�Q˚���o��C^��gI��£\�v�n���hr3��tI[�l��y�O>ϬQ�yv�i5�"J�>��B�z��*�`#;m(8[�\^�	|�l��^����
=�Ht�V�>}�$�=cs�{���n�Ɉ�{Ι�8�6I7t��Fi��5��|{�5h��q[����)U��'q(&���f�K3+b��,Ì�즩o�T`U��'���ocE�ȸUR���ʔ��3�<�g4��-�����V�N}ؙꀹ�Ѡ$0+�n�,��<(�u�z�_ׄm�,�oe��ܷ�rg&h���־ha�.�;Kt��K�j�M�;�8c���7`F�L6��/��Y��kl�{(9��)9��f���R�`Ws�n�f`.�hOt�a�ۆ5�w����$����`h<�мD^>U��	���fQ�0+�̰=K�-_y�^��{��ωd2�"\�̨�h�q��S�hɽ]����
A�}�������X1K�q�;�hl�'d�$%�C��{�I����b�W�h c��iO�v>�m�{���)�/(y�d<��ϓ�iIM�Z��v�Ι�,�g^3 �+^�x�k;�hؔ@�ͩ���Һ���1���B�[��]y	5������C!C�f��d�K���;��^>,���^�*����]m�Q�g0sR+��mm'�u��o~�>Aڧ;1��b����!�K���a�k6:8���9��g9Q�`R:�+
��P1�r
n���|��Ϗ]3SV���j��d��e���}�\7�;	`Qo5L�����%i]ow�����e�ǅ�޶����B�?mf�:����#�K��^p։���4z�v4S��k��7��iF)7*�a��FP�7�Ѽ8�A���f�jb\�Ow���-+���o�]��޼�(.W�� le�pAv�q8�@�ˮ�}��i6��8G
2F��@��k�)U��k4��b*+�_*���²E{Nw+�PV�s�EUl�T��DqSS�<��e�M�Þ���a��*Z!�BH�j�ef���xE9QVI&E�R��"TV���H���*h��n���,�B5hd�B�J�4V�X�$�Q1Y�zR���`mYZ�j�R�ҬI2�BfRTy�x���烔b��.���u�I�U9f�Va"�*>:�Pym
"�9�|ws6E>:��,NE�ŎN	�XjH�Tmg8���Zr�t�J$8E9��Ȩ]r��]�N����u�yN�^��YE\�F�i�����/�/C$���8�*��ӄ�H�$��ʓ���E��b��A�I�Ŝ��R��XV)*).�)S9�(T�ru���ݼ;�qY:�?  � �G� 1�x�vj�m�)�1��k��M��F����/)7���:a�,�4C|�%�f�(�_�{�}t�g���!;)���N��`�����<��?�R�T���=%7�8�r��nY^K4�Lt}j]�MoF�mN-���ω�q�������w����+t2���I�	w]�l[�R���]�/�57�E�Y��D��uQ5��SP/���s��VE���Y�������Zĭ�[�&���++����vu����x7V*��dbg.6�qƉ+][Qy�V��b�4��_�b�N�v^a��82�d���r�ڪ��o�T6{h��TW�f��6�{���4�/p=�T-mݭD=�6[�w�]}�Ye��8��c��]�������k7z2��-�o�x���)��h��vu:���777+\Hz$Z�Un�����ط9Q��^t��\ث������uP��T3�94�3�ޮ����;*Z�w1s����֮u�[��o�)��}UG zff��\��oON���ˡ)��7�T;�36R�c��+dR�Dr&��r��ojƛ��D�l�1w(��[�2zr!K4��v�ѧ8��q�e���*Ŏͺ�Ǎ�S�gJ{,hJ�;o�����`TmYt�����z+�nF<m��7���8�qV��7��V"2&���8���K�RjkU�����x.㒠�'Z��2'�11��D���Էgnu��W�-�>[��>{ٳ�����&|?o��N.�A������}�4�������-%l6��=�;���WS��R':��'r�q<��^ř_[r��{��w2��y�9�z�\c��t�h�2���N�G�O�.�Y^Վ%\c�W���s}��D=]P�
��N*��f��i��y��Gs��V�.�j���.���Biu_j�1c�,8���M�=U������\'��݉�,��L-�`�V���6 v��5$�K}�s��E�"�ч˦\>��y
� a1�K]^4��x:`�C�Y+���~�I3�zs߻�-\�6��t��9��Z��v�<՚��ͱYY�t[�úg8bF�n��/j*�%��R�c�J��(�N��P��I���L�[��-��ҕ�@D=71����O,�跡�N��զZr�Y>�/~s76��J�u��;)j��$��,J��<�s�ێ����r;S�Wn�-QW	���]���}����NG��xN[AzlE�:��������Q0�7mN.�nޟ�\�E����.q��I��֏E��[�xo8�y��c��PHඅS�젳a��@n�q�{��M{4\�;m-}j����0��p���<u{��;�{�I={�ڞ�ݱy�r�����؞Fo(SM��+��,��A��le��ڽ�����U������HU	���dZy����Y\K���#��H[I�t�5|�}�ޣ=y���j��WZ�vyM#�as�e��߱��<*�%�^�O��)osۋv᷽BDԝ���z�6�;��z����R�B\*����>y=�3l奦��Hmv�\ᕶ"�?v�r��S=�����09���&����\����v��7�:?���it¶V��^�tcQ�Ap�:+37��������|7��[*�4I8�.���9�:��8ώ���s�n�����e�Y�X��g�1b�3Ħ���Y����yJ�4q������qS�e��c���>��=OroPoo'�N���~��J�߂�gk2��q=s/�ɢ�Žjc~�3��q�����G[y
��(��FW��G<��ev\�U�*q$�<�섮������}N�<L�W	�	���D��/zu,�c����.elC>^^f����my<���>
��x�u\^TZT�F�$�` -
���K�-l[�1��OyPtԕy�2�6v�͇!ԫQ�v��5���i����hS�TR⼊�*gVS�q��l�u��z_v��=Y��[��kk[vUOY�����V8�%��ѹ\^.����OW�ֳ�2�{���Ҿ� ���ta�a�.$�6���Q�k�ˌQ��=������o��q��V��m.*�y�>W&��K��.ڭ��ns�cӊ9\u���%�-�W�y����O_Rʚ�%JTP0M�Hxo��}ײ���ؕn��@2�C�� C���H�^р26z͏V�  ����fv�������|���"�.Y�K�s+vv�4k5x�:��k�y�q�}��[�d�p!��4۾����63��V_;�/z�z1�.���Ac��6�\֬b}�e\j�Q���=i��)����������jK9A�~ε��|��و-q�Pbw��K�RvS�w��j��Qq��1[�uJ�]8��[�	��S\�8�[~P�`lk�����*^Ѕ=�Ne��;��6�G,�!4���Qi��Ct�j:R��02��3���ŭ�5�s�\���v_���W�4��\7�^��#M�*�BZ3j�Wο-{��a�[[
�nL�Z����jum"ri���SE�����;7qX1�`}����<�[ڈ0��W��ٗVW�5�_S��[uҽ��BmYA`�K��㏕ʞL�}^��0V�[^��ɯ^'ݐ�*
)G8�%^`OVN�r 7q��c��/@>�4IZ�-���zv#9�N�����L����j�y��*�9)�x��c���;E��ڢ�V�3ϙ���������������Q��_A0�ʋ>xM�wn	뙢+b�ͳ{@�3e�0�ݍ��7Z�t��7Iʇ��m��0�c�0��
��Ϗ't�9�f�����������Cww�����B�P�t�X�c���k�;677J�ՖS��_rw��9	����=w_|�Yk���jr�GJ̰��ǵR�Sj�ťN���Vr�x��K3Բ��͆�d��4wV��Wb�:������mex�]z.s��Q�g8ե��/Ck����o�f�^]�6��O{6������ī�\ⱌZ�J!s��-lTO��yzi�. �N:�j#�����v;��]�����B�[:�n��2�6�d�]V$b}���q�p��.�ݐ;OH6��V?v�>9xw�<}���s�y.������)�>[���g�
:����O�r����;��ٯԹ!E��[_tye����qi^8[��FӦ�8;�MT�5A��e��ٓ�]=W*=͙�Me��W�;���U�q�׊0E޹�ߤ�T��Е�a�W_9$���q�è�TJk�`s��ִ���ϳ�}X�р�Rj=��n�EZ;��ů09{���<��R����N�R�XﲯՅb�md�Oݻ���]6���5�+,�y7��{��	�.�N���^��&s�ڠ��V���.�c�J�V�	���G���F�ZuB�6d�>�O*
�ծ�\�Pi��юF+t2"��л7�9�l�������H�{D+��oo�y=­O.����M>���B�C)K<.
�0�i��%ԭ��zԸnq9��Sx�N�sgil�]	�AWP݁0���z����P�I陸yo���.͓�R���i&��y)u�
���:���y>�����!����"�kI^��1r���Q���RUy�;M�>4���rGe4��܋���t�7�U��)v�V-�)0n5AJ��G%ZпD�f�_Ko��lY�9�ʰ��[��K:~�:y���~�����(r�I���{3�9�O;K���is�����W5kj����q�9�(�*��w	��E�
�y��M�0��{�����&����y�v;+�ƙ�䣲hF�����U����<C���޽Oqy��G;[o�wd�K5�lS�Z"Q�K��+bC�9���c8�Q�����kZٝX���jH�}�)�F��,�%�{��V��XqP[���ma8�Vn���|�����)]�����v�f��5�噎qt�>����vʻb�<�V��n�~�����\λ�Vo>�"{ƫ�'g�<�(|��nb�^��@I����U�{��T�=^����ͬ��=j/��YEך|�Yx�n�n�l9��W[z�&�5H�p���#am3��.d%½��n�r�����m�v�]9�J:�[/s�!��y�u�6�X�Yo�@~����{MOo���>,*8)�wSwU�֍q]�5
_u��㌚t�TCl*�`����3V��<ms��W*󐻚p5f1ɾ�e�p�GsOa�a��"� ��4�Y�:���v�5��0��}ۙ��+^�η��<Lߊ���jkE�)��8:k��ѡ��kjn�}]�qc��yP��be���jX��y�ү��o���`/�FG�z�ƗT^b��}��j|�9X���<����.@#�7TN��`kX9����җ�W��d���ѯY+nM`QX�U����/y�{���`馲�m���7-l��ld5�����)Q�Ҡ�pn\��&��8�zz	 ����k尋{AV7z�6��_�Y��n�a��l7y۵�XB�R�
x��S.+����.+X��4yv]BT��1��&�Z�ҕb@t;��q���}�����V���7ޙai���0��פ�%߻��%L25��jM\3�x�
{I�gc�o��8���sn*����#��e���K��t���)	�K���8¸\��Χ����o�܋�����;��uA~�"�%w��z9���l��g�$"T��x9�<�������P�N������N���&�����J�y�R��@j��m�b��nK�z⩀&��b�&u������e�����V��_wf�}�}t5�	�����m+�S��w�2x��9�7�L��0=9/]�`��q���FT��X�_�'�����߾�4t*��)�,�y�f�����'�� S��Q��Sٵ�t�;��Y��c���\�[{p�t��3(n��8>��nݹ�9A� l���S�����녳�K���:��ó�yiسM�%����ޡ�v���uH�6��쩸4ןF�f%P�=�LLwU�Q�,,!���;iKƩI���V|4��3>U[��*3�le�}��}նa��VT��e"��0�@=6���:�N�=�ڵ�ޗ)����������z��f�Ɇ�4U���E��G{:�<�4�ʺ|�=$��j��n�g#���]>f���ݱ�|M��85y�
���k�ژ�M.�U���������¾$��Ύ����Dx����IS���s����y��-ݭ�9��b�W�y�q��5pC�"e��L>;�	���hߴ��vycB�������w�B�
�A��p�j�`j�^�U�,\@w4&��Q*{�6�ݸW�WI�iR�M�50����u���;��yu>���'֝L֔����ᓄ�/���e��h����o�V�ݍ]-��S����\�&�4�v�fC�HG@��gCwU�+(`����ȳO��4~���]߱*��iR���	�Mxg�ziS+����s��ڑ���-Yp��3q6�j^�ս���AX~�)����^MiC>3�k�7�������"�ݧ���W"��?�_r�ԭ�����r�P�]��/�?a�dUB�Y^�7�U<��-���Fѩ���yo]s�K�j��}¾����ΐ�~��W�R������>�Wp�2g\��}	7~�r=�y~��]��qZ�Tf'KO�t����/���*�[}A�����԰�Ξ�u�k7/*�]�k7�$�4�s�̚0�|��:�/�������s/h!|W�ej�s�wXQM�¸�W�e����U��.��<�kM�����V�.9jtD0n>'��J�oWu�� r�,�*s 5թ�iru,�%��>5�'R�s�i�{�n��!S�4�ŉCx"�혎,�)��V�k8uf%D:��6�Zv���SZ�|�b����c�of��}o��`��D霉r4�wPĞU��;�(������`��a��{����K�d�v�f�����o*�à��I�``!�I*�L��Z�6�Jށ� 9T��.�M"�3���G�_�E�O��bv)w�3�n�mN��7�k�O�,H��3��t���'������N�j.BӚ�<�e���:���[��E��i�83WK�9�l�]F�h�g����&fY*��ü6D�5������8��e.o���L�x#}-ŏ�Щ�h��WW��>��N����X�:F��(fE�Cv�k5ݸ�ͧ)���Kg{`c%+2����ޣ�@�y�t'i۷�醅𛕏��]܅��&ڥ�,���XXMH��a���N���Mr8�v��P�7Szpn��|�E[����%}�)t��ï�w�M�_��2�f�@;J1�z��1�{j����8�ѽk�=]y���YV�����D��{M��{κjb�= 6Y�)[d¡�Va��ı��=�YLzg�Uc��hU��/�{'���ú��r7]ܘ�{۠�l}�� ��Ȏ�c_A�"�d���rɎ>�gz�|
\Ll��L��]�FnSE�yKD�Y�oi�I�l׫F�p��K�E!�EnS��h��;���:�8�׼67+EÆ�xBÅ�ڴcc`&�n.p��w3%R�ڻ�7�ۇiթz�Z�Z�J���!�fA�h���Ô[��8��:�t�������|�+�䈽�u�A�}��Q�o�ݕ͍e��QcD�7��.���Y��e)x�=����K�|�HQ; �dw�4h�W8�����n����es3��!�Lk��q�V���\~�T�Q�Vm���vv'�
��yKkR�gn3�����U�n*m��l�L�On�LZ6$H*=Kt��*|o�� �^k�؝��ٛ�r��s|��QDB+�'Q��Lw�np����S5t����^�}פ5Ձy�n�&"�D��r��Pý��T�/�'{C�����곷�Sʁ���D#��>�OVZI����"���/�h*����Ԩ��
�x�n���0OV�����=���u��#V�h���a;$6Wd��LK1´��t��y�1\���(���{3ؒu�cd��"@�f��c9+�R�}G��� ��h��i|	������FW�s3
=�����}����s	/ה��9-%��9�~���D��ϊ�4<�<�WP�u�$K��C� �&�F�QZ�TH*�$�Q�T�Iiu2���.V��&QFGP��!dE��Vu�%�G9s%���eJ"VH��eK�ψ��4$��UfE�fjZ�)W.s�[�k!��9�jʙDT��ť��I��Q*F����v�vyA(���^!	��A�E&"JkC �X�UQe�*���
�����U��Ԣ�\R�U�DG �3x�U^aV��jK^싕DD(��*��Q��E+KkM�(�Q�&"Ht9"Qud�	ɞ�kXU*G-Z`��B�Qvi�Υq
��&&���歕r8QE�D3����&Xe"ԸTf+JL*���
���ڬ��.�l�L���,�=K���Q�EJ��̒ĵ
�i�Eu+T�ST(�$�K��$�ZH�E�.PD�����""��$�*�ʪ���TUW)�+�$a���Əe#�*I�6\�c��X�t�"�<l

��ny
�W��d���ڱ;�.!�Ӷ�Ny{���VH�L�֛X���7���T�ì��#��'��C��g��ٟ�u��� �}��*-���q5�$�=���rd׫x���^�g�:�O�i�8U�3̭Өw��I�H�Y�!�=�j�w�gj��:\@��(i��]��"�{!m��K�:nr!5J|�kEFC� ���Y��j���ݯ\t�q���0p`�U]B(s�����!m�W��$(��D�?C���n}�p�[z��٧�%��/#~�5�ϲ��,�.�-��|jИ�S��NG�h�����_Ѵ$��:��W����n���Ҽc�0�� �}�@��Oze���`���qW����3��t���:7��V�����n�d��I�����T��eL����C?&�3��EPM��3W&�'�i'���[D:��L�׵�JX��vn6ڦl�z�_*��Ҷ���8�U;^Ε�橐<�#��7N{<rV�a��+uV�7J]G,��8���z���M���A��o��qV1ؿ��1~�	Xo�%��;P�����i�;��_7�lQ	[�:�e�#�B����z������%�O�`�;�R�W}�L��[���ǎ�<��s�3qك`4
�W)���a��{�z���~s���<�󕷋��3�H�f�����f��;[�q��'Y�:'N)V�*���7ɱ�*�ه��4`\�������-��l����F�Ԡ��O9~�mn`���=w?L��c�����T���:��\�·��*Ѣ����{� �+�d�G�Yf�V���+�o�V���tz��8��PS�}P�oH3�C�q���_��ڮ��E�����s���Z�q���{�}p���+���(ݓ�f����w�<�����3��N�>�/L88�xdUs��]�z�}c�*θO��:z>��q���欶��ڛ_';�����!]V̛:����S޺�Y��w+>����ͪ|1�~Q�y��d�yy٪�g p��J�����5'G}qT��;��G�y��uSЧ �'���wA�������c����kbC�s���0���¸�B��x��1�"n0���|��p�=�{r��;��xl<�t�%���ߢ~��������B�� ���#q_M
�+�Ah��{�8��n�����s��Y�ߓ��p˭�C�ܟM[�~�!�H��`t�`f��&3-m���r����GQ����ZW�)�������/@������ybm��%:h.���;î��APr�2�j��b�����b&sIEF������r�Mg�g�9���DU&<۠�]&:"�:�m1|_{Z���wP���פ�p�S�tǜ�,No�o�A���]}��[��q\痀EX�S�sow<����mW%Vy�y4�nLS��~���4|p�>����G�.;���ʪ0�R��s��m}m!�?^-n���[��K�4A�Y���X����%�iՓ����c���oB
>�z�OW�;6�v�k��ӳ����EB�O
%�w��W�#��#&���Թ�D�ZB���'>w*�fl:��j��3��L��U.nɡ:�B���\�^eB����(��]Q�B���k����� �ۍ��ӝ���3]�訆��.�/Y2�e���vX������}ػq����M����}�L�Yo�c@��.�q-I����w!Eq��?���8���{�om���Ul���ɟw�O�����-v�?Cӿ6wE��6�i�r����ӿ*��un/����+�F>�����Ir�
lc��L��]�2w��-�5:��^�# �ؽ��^��ֺ�#���MJ�t��N�u�)����K=�[��<������@���ݲ���]Π/���Eh���9��]��q�MF�F:D��9I� ����X�*�l_��(
۪F]
���[�+�t�y}8�"V�T}C$s��L�b&}��.HL�r��4u��J�������O�����Rdiz[.\o�]�h�l
��fT2�{�Wkѷ�˜l���^]�u��9��K��s{��v6��P��X@��x,�R��!G�a�q-���>���Vt�^�?o�7n>��ujج�T�r�8�7E1�g[�����ض�;��V��h���8èu�T����A�C>�2���ߧE}��nK-Dgn��@ڬ+d1p�f�r�s6(�=�\aR��|���,�I;�ە\���
�j�o2��Q�2q< 3���
���]
%�ؼ=ZǽT�}]$#�!�>O{Һ�K͊�S;}f�Z�S�Vj��K:��"�1}9 .fs��� ��~��/A�|�Cg�P~��.@�����ܾ ����9��ec���NOHh�A0�T[��[^��L{��O�����5W�w9%)�s�\>��Ǽ_���a�b����5,w��6�ل��*KG"���x:�<�Hqa �[�ZV**!s���ک��+��
��N��������{W](��Ǩ��-��;��������Z�T�o}�CL��J���]��YG�����ػx�i��~�8{��O�*r�y��~�d�7��_���`'_\|9���+�nn��D����;(ދ��U|��s6m<k�mAЊ�ɂ����i��dJ(��;�`��ќ�fB��K�����M�1���+'�]��j5+Q:	����ur4��	�4�%6�8B}j%�m��_7g�� �gXoN�O�@�����wڐ3S��*:q+Z�(�"���w,�hOi�?#�;Qus��;~�Ӭ��<���_|Hx�������g�����A"7�d�ʐ���h������+�*����m�Yuo?���/��S>]�h�)X��}y�#��/pC�W�7l�7q}|:�>�-��H\fIF�b���QC�λ��#Y�������KsB���6t�������h��0��E�q��د��%Q��Da�A_K��Q������__O�q�[��6�E˅�I�)�;�������;����_\_<��:��Hb���o{Ov�ʾl� n�U�MJ�������R>I�lS�=M�w��p���̷�(���_��Z��~����C�٣�)���-�K���X���w�S|��7I�-��U�����R��<g��Bw�CN|n@!�눙��.���,9�~̏>�[>�f�J-�X\�c�-ފ��׶���i�����Y�0��$�b^��s������ޚ�z�oo>ϔ���$J���Lg��t��n�3*�X��UG�%ó���J����>hu���O'L����y3w+�%WX��ʜǍ<K���up5�\���ڈ�t���ʳZ� �p.y�6Vgõ�"��|^G�zȨЙ�R,.U;I?=�"���#�xp��M�fk��xg�5rs&�GL�=Z6����:�+x`��혺��^�6�����/�c���y��
���C���%�R�"�S)� z`pƨm� eΧwr7}��u�o�T�_�������oӿ���ݚ�\G*f�_�ک|B��7wL����пv�ό�`4��!�w񺍫9��)do��]��^D#R�j����o���.���T��|��-8"�9�VeR>Ӓ�c��-�u-~�>���
�~ M�=�v��0O��F�bw��|�3�����~���F��e�r�`���k�'�­�9���j�dO�Z���v�g[�O�e�\1�WU��V���tz�S�	SQ�>�3n���� W�ڿ\��tx���S�p|Tϙ�Σn�`\?!���;���p�������|}+����Ms�r�|�����1զ6��q����:����'nZ��CtW��W�[����������湞CCbg�5��,
=�aF�S�綥q��-��u�:�c"�~4��|����2~Mg)U��[��_m�adlL�G�b�L��`����;j�#��ͳq��ʷ"�$�5�8�{L�7���za˂�6���ٜgQ;��ŏb�Ul�o��!n�֞��VK��R�BG����iG�B��&��l=ܠ�b�)�A�e־C�7x�ᯝ>;�.�n�YH;�9V�����s��mg���ܯw�\��%wb1\�%@ڛ`e�c�]����S��*:t+��RM@3��Ә?RU�\Fa{8c�oj�e�>�dS�^�pt{}�=��As���`h�?���R�t�'F�顿b}�+>ה5m��+������m}C�S���p�Y�qV��p�l����V�Y��d.�3�WQ ��ؘ液����58��S_uȉ{�㴦/�y>u��\1��J�t&J�we�z��׶�<�}�'������[BLW1�����}���'Q����f2�s%��O�*}���]�X�R�����{0��D�u�n�m�0 �i�+����FX���	�4.������fh����N�ùH���(}C��LJK���B��+��Α�r�˭jV��uvwL�=/�)M�TP�mT���eܹ�rH���p�;4�/���;�E��3o�隯{�»��A�ͮ@ڇ&�jr#��,!�\w��]ŭ"�F�8`
V�^�"�YB����)ngx��q�Q�g+�o�!�d{�����㜈L�G��_TV��l�^���[׵�t���pwA
Ȳ|:f�d�N^��C=�K왧��{���t�����Fh�Eݑ��/k)���`Z(��jb�OrI	��4���Eqg�6sC��4�3�eJ���:ԇ��۴�C�T=�;ҭ�;�Ѹ9$��yɢ�)���L9��y�!�&rs�z�p�7,m�N�q�ZU�K���_ϗ;r0Z
v9�|6����}^ڼߋ��}�_����(>ڤ>�dօ7�a>`y���r���.<�z�Z2�����<A��}s�~��\m�ݖx�X=Ą��������γ�Em�''RL\PZ�o���x!��kT��_Cw����$ǬH�����Q�&+]����7�|g�U�7������ԡ4�d���F�O�#̩�n��yU����l��� �8~R�|�<��n�����Ë�M^�H�=�`���ۇ�'I���k>�̹�9A=����灢2�g×f%_ ���j'j���'
���!⸚o�H�}�*L���E�b1�*��Y�����tm��K�T�b�`��%�]F�b�x��7�H<�(mK�F.~�~3�u�7����7����@Ղ�,~r� Et���^�D��>����3����aѺ���ڱ�-�Z>�(}=�l�y]"�ɞ�o2�rzEA+GY0�T[�)mz�ꄎ@�n�y��gnm��'hܵ�<c�ځё:��:���2�up�����C�����	��>�m��7HrLԻ�po?�q�)�,���Ý0���eu�9�J�6�Xw>�o
�K�;���_{��g�h���NkҘ,8�e�
�fi��\��+�T��N�(9�\[O����>��v��1������TR�E��L��Yw>�� �;n1Ϥ�D�[��N����J����^z�*����<T�&��)���.W;��O���mUC�OЯ�q��mN�z�D�~��?i�(eNS\d�����h�9�s�
�R��޷��?*��/�G�C�ݳx}ku�<=v`�]�I��!���ڋ���J�֕�@ߗ�_�]�/�ܾ�rpnuB�z�L`W2�>�=�<��vzL�/l�Tu��B������E��55Q���k�UwX�ी��n�F�߯�m��7r�î>�--��d�@b��z�:��� ���CB��%�M8���;"�Q�UQ~�����Lo�<�З��GG�:���P��1u���3'���������v@2��+�:Û��I���Z��c�я
�}W���雬���P��.�ᙓ����%���_Q<7n�|�ԇ��Ÿ��"9^$�,"�O5�髿4u�R�b�g��j��(yy���P����Z�6U*�H�蜘<����l�3��n5گ	�9o�f���Q��qh��5�r]j޳:����4�Tm'թQI�Wb8+@�wE�ÕU�2Mw�n��wIZۖ�e�����^�<�2�q򀐨fw�dd �D�a�[$wF����>��W«>����=�GW��~��Դg�L�t���B��H���0�]u�g�{���e�s��y��o]N�[[�wֺСq/�h�}����`h�����
�h� &=|`rAi]L�8������]���d��!1��\_�W[��שHP�L�z��������y`�q�=��h��C�/��	1Zw��9xg�/�LTm��]���/�|VT�[y`^�&}��0٧�����tN���^���HT=G�_{�N�j���Q�i�֜�u�)LyZ뺽�{aǴ�8�F���������6���;�F�H5�j]�ʮ\�e8����}�;uN���g��8�*:-?U�ȕ�&+\���z�������iY��I�X� u����w�)���}3/�盎S%�
4�y��ss�U�}?`b��V-� ~_��)�l�4e1�v��Φ�� Y�x:}�#�nfj!zݰ2:��2_��R�$�큃*q����{E�
�6�6�e�>�=

�X��)�b�$�A0��5�wf�)�;�ϭtT�y- ��A�cλ�0hy��>6�0/-�$�wt����ٰG�QܶO'�m��	���Q���~=a�s�����9{H��
�>�?!���`4�<�GT��[Ξ�)àL�U��t���_�{U�O;=�S<8u�bwA��0͙8��xw���L�	:^,�W�`ny��1����<�vDS�8��C���F�ݱ����;��v�a�9��e��~��-ȏ
ӝXKG�]�Mk�B$�c+6��r^G���*�	m�+�t�QT>T���?4�����C@��t�T����z�zq`��诎^da�"�7��-W[��&lP,���,+��Wi��߁���)Mv���ֳ��
��O{8��⇋�sGa�Xc]s�F�b�v�m�/}�#�p<+�b���%��@5WL�aK�m◕sv	k��-S�>�PXVm��[,4��<)�d��y�^N�O���7��3��u��_�m�}X�i��\"�ä9�m�V�Dڛo|�Yi�>�gK��s�s��`Ր��ovI+���;݃�Z����S���ZƩ��>��Ű�ܽ�)<Y$�����$���8���C��.��P�*��X��LʃO�Q��BԐf�Gu{G/��1v�Y�Mi>{W)s��D:u>��쾹u���u�ۘc�RufN���L�%\�e��Kv��$=��ۇ�>�$���:8�;�љ*�TB���ϧa�	�(��rg�o�v�s�ɚ3܃ǣ6�م��x냫��)j��4Қ�k��ml�NW�*eih*��F�-�Z����o��'ۖnEU:X~�Kn`�!�N�]dŧqb;r��Am��a��3,��*1i�(����\X�u��̻�N�h�Ē�`r��x`�
������V5Q�uw��,-1�g���5�5�����ͩێ��B{AB̫{�u��;� 9�^��mO*��c��c�덞�����s(����ĬRk�c��lU�l��I�޼t.�W�c;�2�	r�6�d�8m>���ff̝��;�	N�oVnv���bV
�'n�b�z¥��1/7�2�ᱜ��FCb�1������������|��v����xl�A�[�����R��#4�ͷ/�]����:��]��] ���0�DY��\�����ռ&'�>)b+�v-�+rwtΘx�T�;t�sV�!���Ǹu�W@�o"ػ�J5uv�e�����間z�I� �xCZx�	���El��׏M�`�������bM� �r�\��ԗ#�v�F�C��1s5`������N����{���v���Շ�Üd����)iDQG2�EEf��L�\�:I�Ꜻ���HNH�TW���4OZNM(�邬��5�D�Q28G���bslC�*��Ej��9�q*V�^�8�2*"9r"��%�wZ�*�9ʮUYs�".S"��ʬ�L���.Ȫ/Z�DqZȧ6�DHT����G�s�(�Y䲨�T�]�DDJAB�J�!\�]2�DQ�z�IG�u��\���w1/"�t�:Ȫ����]Փ�r�%*5*��A�r��9�E8s��β��T뺖)�V�UT)B��s*�XZE�B"̊8{��	�t�N�S�)"��*����c�D�ȸ�T���T�W3��rwqtHۻYʢ��y���K3:F녦,�X�^Zp�����#�R�s*T��Uȋ��T�5��"�.ZG��tB"+�!B�E����,s9U�ig+���Qa%Đ�J�	�J���Qܥxx�J�� �e�*�7��}�Dy�rz.wlֶkM��넷I�7�/�:)��}S��VFe��qG�[�x	W��T���S��J��9ݘ������q�R6n<O��\�6�]�-�֡ݭ�.6���nN���t�}>�̪�ד��=��.F�Ӷ�d�1go���}�ӗ���轜�P�%]��':��k>��� r����,߰������T���)�ۖef��W��:���4&g9��Wht�V�|x�7Pb6�	�G̩ت`LT�?xS.�����9q}�=�tZ�)Ff�ˬ.4�N}��nCt�#G�O�Q��#*�D�:� �7H��>�=���ksig[�;�{U��PןdV'I8{�w3�nݹ��Yy ����} ��-����Y;�v��5[�H������^��(��\Uï��6'���K�ݫ2�,�W|z��y-�������P�wW��{��
}l�χ�3萧�3>��L\cJ��A}ؘ��f����2�U�)uIܺ6r3�|d�5S�d.#���H���3��2Ƨ�1��Lf4������}��k�n���ӳ�+O0�N~%C�&�\e|LM5[GY�n�#LmI���t��
���*��kt�XIð�����!�}jf����#��g�艽X���A��e��p���w��v3|�.J%�da�o�K�S�ڥ��D���vﻋ���e���.^]���*з���])�0�c*�e���gm��z���Z��\r��(�d��B�Ԅ]b�����ѫ���?s�||FK��H�����D���uo�xG_ю���{�/p��ywE����6��j9ا7��ک��eܹ��hM}̎��s�Q���#uy�H�Z���=�=�@/6�1p�e�ƪ��25�N�z��(]�}��r�zw�f�gӝ��\�u}ct�P��h�����y���9��������8���P�6��Q��1�)�vZ�9�d��<K�>\�d���V����Wo������-v�_���6@�{�}���t�g��p�l�`�������������>b��L�d.ys�#z�"v�^	��ݔ�ޠ%ݒ>���{b�B���#�Q��R=^�0�;�����~IN`>�ύ7֖ۛ��q]�]v#s_���}ξG���j�6�{�PZARC�|j��07M b��F��}�}�)dˇ��,ڨL\��g�J���|ei܈�(���S�Yy@����5Ċ�or���[���?z�
ޔ�J��{V%�U.��eўehf�9�un�YU������8�]��^�#Fd|)8���D&!�[v;j��l*[;l	�+6;�ބ&:�{)����WV�����ͱQ��H����h��u��tn�9�\�{��,�Xuw�duk��yc���H�{�0�]˖ 3����G�w�Т�o%����Hoݪ�Y�lƟ��Q��˺��.xإ��۽�����{p����sbA�#@�;y�ϖӕq��[� �{���[�M�-�n�~�:>Kk��=�H�3��"ܳH��1�;�LLS��H�2Ƃ"���^W��PԳkZ��Y�c}�:�7�
���d;�����A)eh�"9��u!Ĺg9nq��Ux��[=��zn!?�t�}V�|������ky6&�28 �C��־�j������Zߘ�K���[��Q���;��q	X�����V��L�6�T}~(���wnQY��H��姻�2��h���=�9*�0z3ԧA=�K��2s���Ϫ���!��^��}+����@Q�v���vQ��?��Q'�v�k�����tV���w���`Kw�Cݸ����uU���iv�ѯ,�O\{Y�O�e#��Kz�[���^*�p���vT�;sb���f��s�pBڽrF?��'#�\:�YhP��+B�w�x~YP����[F� �.�H���S)��h^�Y��$����x/�(��d8�C���5�:���v��u0i�h���j�J����{r��ŒA�+�/y{����k��J�{�pPw��@����##�!���.]��ْ��2�o77�k��h���v�g�V��|��}吝�����C�WM��'��)���y]Fe��F���`��ۜ�~{4�n�o	��^��C���G'oF|��;}.7E��{/���A�V%^�!{r�"Fߖ�~s4�T�uNdޫ�xy+h�f�8�v�zLv�x[2��հ�h��3�_C��+~�P�>3:�L�;̋�=)��.�9����p[���vD}�\� +ӣf)}똦�?���p����A��L��,���a{؞+�����D+_M[yo����Z���ј6�p�8�"$JGl�)]WP��z�ry�"�3�7��{Ն��9t�����ToS��7�N��xzBQ�s>��v�ͷL\,�~g�dɾg�{��ջ���f�A^������8T6.!4�{I��<���<ٙ~�s�UH����*ƣwtު~���>���'�w���Ǽ3��h��Tu��b�#�2Y����Ŋ���}��4� C�>�x�j���"n����vV��~=��~���js���{��Lq�@���,Ҫ�Ök���dᇲ���S� 9q� �����&wٿ�g����Xlk���ݠ��FP�b�'Ρw�%;�`�G>{��Z�V$�dY�y :a�v��Dz�-+,u$4"�̓V+8)W-��Ơ����S��y�]�Z�����sЗ<��u&�cZ5�\�w�[�r��U�4 ����B���.�����.t��>�{iK��Y$g��{<^���B�bK�._���_�!mz�^DJ�'\����k�~?-lW�'��'���k�����'�{������.#:�fk�ۖ�+H�3;�C�����9~�h���C¯t �R��j����{����W���ӛNdt.��>'k���r�N�N��EhVN�T�V&U+��]�n�t8���\ez��}G~>.g��˝L�v��~>Cw�7q�.θ���k::G�'/<,絑=/e��%�\rF�S�Xk�\a>f,�(f�S�N����i���v\%1#1Z�߱����脵�<�E�<JD�lت`M�|X�����Ԡק��}݀�eg�F�#%��ϘKU֠>�:>]�|�}e�r��7���@��I=2���`^˱V����r���>Wt��;EwХ�bFO}���G������*�*u
��Tj �λ�4�g7<�dmcr���V����v���on
X�������33��ݻs��At�H�O�yy���h�����U�2��7韕(z��Kk��^��k�s�ۭu��e�MW��-�����A�Z�}{�lW�.U̥�����������S1���m˓]/	��ղ���gM�|S�e];ꭊ��$�[VL�z$�K~����١P{�y?#���(�x��.�i��C�M'n̘�MuB|]�t^�7ܗZ��$��,:�T+�����v�i\/m1�s@D�7{�c��}�U������+��Ȩ��W�a�ك�.�H���]Ƕc*���/E�:{V��_v����p5m�O�L����� ��
0��|LLSU�u���-c>Ϙϧ��^����g������2U/HB�컡$Rbx_�&�^V����~F����u�m{;-�����}�zqT�5U7��� ����s(����r�e��oX?o�s�$N�]�����4�|2��L}�6�����ڄ�7�nr�(pϵ�N�����J�7 ��W�ee`��{�=��ŖJ	ڜ�d�l�l���,	Y�����C�������zr���|ȭq_wm�6�'�ߧ�CoӴ�^MiW��ׅ���g"=�έt����s~R�[h�B�>�,�Wq�K�\>�<b�`��r^��fp��3��t���ZT����?4��iuΉa��u7���4��ȝ���fM�:�h�hpp�l�f˩�M�G,%�&e��nYt��Y�V�䗁��#{�u�m�1��|V�����j�X�-]`�c��Y�K�e>�v�������f����wlQ�2��2mw�D��N;��5�OF���m_N��m�b�0JF�K�zf�}���	5�з �N{<�6ѱ�6�_�iX�g���>�_#�ﲾ~uv�����H,ؙF�%���!�Ǫ�y�Y���-_����p��)�����y�C��L��������ۭY���������j�lv~���i*r.0�	yU�!ԟ\8c�v3,��?q�=�7����~�8gsRp�v�>�_uPE�f�����\�M��;�}D'��SRF78�s~̃��{ԕz�-��i�
�n�cL�����uJ�A+��r�9�}_��d��S�F�cLo�]��s�`��_Uj
r<�'n,�Qn����\7�&�(�����v>����2W�j)g%�u�X��k�𭞴�!Ӆ�[�p+� k>̂��v"e�W2�O:ў��[X�Y�w,���}����Jg�	��99��ҫcU2v����O&��d ���1U-�L>�vuX�����8�y�G[��������%/��f�Z�����e�²��^B�g��y��7]1Y�����ܬw{��n�u����V#�F��"�!�����V��5��u��XC�2˘���8s�Ǟ��')F���@�M��I�rz'|T��Y2���|riы�A~���m���X��Ko` �CIV��7?y��߲w�5���39�X�������;�ʙ����;d/e�?Pk��q֌�UE}�5���Ӟ��;s����p����Zn3]~s���]�؇�N#��b��Բo:[�.߭���_vU����1~��Oh��\=g�.2��7�5�jw��;�kݪ�l��][���IaH����J�C�y�օ`��/�f�꾜�=����y�Tc��v/��S>x�݈܅���|���O_�e���C��Y(����U��7��R�^���q�⇧Պ��>e�W���ê�=�Ȼz=���[��*9?,r {s�yA΀T^I��v�7�Y}�}H��( z�L��]¼<����I���}��xg͕�H�I�|]Q�~ُ�/��ֻۡsTPw���\{#��!�3'�A�3��L�;̋�ޮ����{��Kә��j���J��;�*�C��z,�w2��#`i�޸�t* Hp�a{cY����[�]V��Z����
���;�u3���y�u9�W%#���)]WP��B�d�����[u�����|; �;�1���$�MD6�BP66
($씕s�hӻ��B�:V�7��c���]�<� ��C[��g��couwq\]��z^t˗޾�u5,�ai��wۏ{M�I)8)��i�1�۳i�2�."��eY��̷���Z�Y�W�RG�Ŀ�#���H������v�ӌ�P�$4�\$�gFr�϶�HX�~���
���>{j��;�p^�b]���ߦe_����ǳ\�jvD��=�&�pߜ+��$��Aq0>o��1N{N��;�"��~�O�p�>U_�g�;�z����[;��V��_{{,����t�>*�n����u땤�y1����T*1<d���%�{ �zA���;0�ܨ|�'�>��H�{�Caw����.t��>�R�9��m[�w=�s,�8�M�;##uc�(�;�U��,ev�/�+t�8�nMY�Q�6B���.��<�{lI[�9�5TW�k�����jn�צ���.e���R���X�9_,�G侨w��)�9�s2�N�	�pТ̃��鑭�Zz:5�$�Q��]n����7�~J����V�a���c�<n�} br��,�gs��w��[�y_@���rgR��OV��1���[`�X�w���X���>U�f�9:R;=�Я�s�UNS�sf�c�'������<�l��v���Q���t.^��y�>�1c�{���[���fZ���)�-��T�h��6�7�m>��v�O��鏽��������/1r�4�JJ<{>�E\[&��׽�%w����Ю�������xA٣����j�G�Z���R7�s���"�,\dο�v��d}?qS������h����&�N����-d<�����<�Pb7 >IS9Gx05��'j:�]������<�6�b4�9ȍ-ߧ<���l��5\p���q.�x��zE�㓃��>Wڻiv� �:����?nC낍k���A�c<}Jw}
�rS�N}�����?TP��b>홼�vgʾO�J��hT���d�~�}pQ�x��_�}i���G�K��;U�(�ǲ��݊�oab��_���_� �0j�P�_���{BaE��}K���zA����ۿߣ���[��o��艧T礂;�10�U�&b���@��9����=�.�jM���}�}�6�y�V���̜�,�O\7�&j`p�G\�[q����.�PN[8L溮}{^��z��y�6�u�ө�c�u5�K���Ț�BP5/��7P� �[�O�����.��]t��a}Μ��/O�m_Å��5𸆪�ک��]˜��hMs#�z>�kΘ�J���h��V�`���fc ���m
��#]�N�D�� �R��!�v�o2��tl��
�u��
]!s7O���*Gm7)�������j{��	�Q��{%"����oQ��}||K�TC»8mv���{v�7~���<�Н��
3e W�{�c/���*ie��ƍaQ�7��C�Ԭ����+�*BjU%Y�!2������ZŃ�.�.q��ǔ�onZLO��7�YڸN��=�.�ù,�Jg5��s���hG�m
�n�X:��J�׌����g�wl��m�����{��/;g�V�e�����C'kx����0д��
��g�ܮ\��G�,�V�T7|b���r��K{F��}+R�m�˔f-3���|F�2�0>���B�N�^WS"��{���o3^����P�]�W�O���;�ѭf_"\�K�Py�K�hr����h�Z���0t�O��x�vIn_Gl��I��;0�r�7ġ��ĳ9*=��H],�:�g}v�f��hV涄|���ѓ��iX��jg!����W�k�:/	1�u�nd�o�{���4�^�?����7_[ǯ�\�0Q�B�n�j'9����;h6�q�qOg�rc9W��
$Qv.yy}�M
�oD��k�7rl�a�K�6v��n�b4@
�|�S�����/0g"՘���\�Е���'(n;��v�5
�U�Z�� &�l�!�{n��E"뷼9ۜ�(,\��ܴژ-�P�u)�|��@R�Y��G�c:pfW.u�e�u&nz�rΪ�����V0L��R�޻W1������T���r�B���a�PhCRm�䢒����O]�[���z宰�{"����O�wJˬ�	]�X����	�-<�i�U,{S��7M
��K�^iJ�+�.�)���@�5ٛ#��nqo30Z��[��iLbj��M�]n(�+�ښ9P�8n>�a�a���;�l���=��}�w���1�9(3]v��u(��=y�v���}����p��S9lw6�����v�q7'1e:�(|���]9�E��Me�:��B�WY �����ӂ����+S5Wte�ᡦ#�����.w�_Y��2���[�2�&	wf=KK��i��]��د��eo�|&�]o^�6)i��mv]�l0�˃����#�k��3�T4�Q��e��v�;l`\:�k�mG��U0���:ú����F¶��'�1�;2XP"��DB�C�)M��K8�u}Gh�����#q����RNZ���}Z�u�T�qݤ{`�pӃ��!!�Y�:ݚ�]l˘^nmǶa;OA}��mo�G�{��y�wm�vg	��V�1ou�_�inwvkQ�D$�.�1��h�w�D���1AO7{Ըܚ�U{A�r�G(������K�`��}�nk�{�9(2��ʹ�LDh�}T�ُ�{fxh�Y��s���@I�����yܜ�\s����(���P���.�+��櫩z��������B˔z'���B�@�"����D��E��"<�=q/�9NV	�&]V�.����W����[�#�j҈�8V��I�e蔒䃺8^G���T�Z$r��'Z:��M��Hc��E(�:�twwnx��N�z[/18���Dq�=�r��N��n�"9Qx)�Ay��)�QW��Y�e����W�R��I���rwm�9�k<騄�Zja'��ԫ3�R�6�����J&T:�����+�QvW�G��8�Z��YS:�:u�\��W<�]̉��ّ���9�ˑ��r��	����]EBr-ԋTM(sG9��J�(�Qk���g�&�uj%��F���IU]

���"/Y��]�ec��U����'��	�:E9�9)��u���I�J���9������
ֹ4�:S��/P%ef�VM����Cɾ��7�F�jy��K�{5rγ3��:�.-�|�����m���\�	������r�?����a�p4�ڇ�ע��p�n�2��uA�4�!���dT���5Ԯ�-����ބ>�����Y*{�ϊ��rUE��7�*_��iz�9���P����x=~�v+ه��h��G��늸_m�6�ǧE�O҆��1�gJ����F}7��m�!��
�������S��x��q�J��m�0�`��S���F�7׹B�^��׽��k�8\����r�`K�/����u���=�"�F��!`L&=��m�C��d��vi�������hvWnd�m*��v�dC�O��;�ۆ����>�ӷ�N�ؖ��K���lO��^�?O��Q�������-���O����g��;�ӟOB��RK~W�f3�f�eA��'1�>��D)x��E'��|�Je�=����y�_Sg~!��Z�-8��]j����.�4�;*rAd�#��+�P\�M�%��܇�B����Q���r���~\ g�ՎN}�a����3�V�\,c)�� @Hm���EҢ��;��|s�c�"�1Z���h^�U���+�]��Y�s��V�f-���"pX���fq�����/
��D��x���񌵁������q]32�ƃ�����>�}�E5�G�#0_&�#���1:������s�O!i=�}���^���#�s��\m�(S&�ߘ��&��i�6>�E��g�y��m�@\�ۏL�Q\h�}&�ER4�w�U;���N�L���'�?�:Ht��lK��;��L��y�&���*	Z:��5�ۂ)^�;ܷ�:O`1;��~���vB5M���U�>j�^������hL�
U�+������̳��3�h4�͢z�l����Ezzi�5ᯮl߾��"(!����}����46��ǽ
7�)�/�D���Ĭ�3��،���6�Q�Lp&���i�d8}��j�ȥ�tr�薏JB��o����|.s����D�����|?_�wO����]~s������e��G;���/��܅.�R;]O�=ʹ��m�1}��q%��f���������Z��1֭5�#��]�5_�T=���#�M�ޏ�Z-���k���ƹ8�@��>���;���4�N�_ثl\A�,���F�-.�c�o����Y|�`�2)v�Ɍ�7'��}�=�L�¦谫�}����	�Ϊ3�v�d=)��D<��K����%O���S֢���`��el5x��Z~�{��]{v)st���x*>;�F[n�SB��\����A���e��	l]f����N���Ho%�O�*2R����u�@�D�Wn��ޫ��td��W��Mf�B&���i�R�b��,�APyVn%j7�	4>�[E����m�R�7��_�\����)��)���ү�7J�&�'t��y��x����z~]-�J�o��e���OH��0(���a�H_��F^�n,,fG���k*37�K��{�K���~�������P��gx�3�$8���z-�\n�l��繴�o��o�$;���C=�T����l7S>�yo!�}P�w0
�d7���!/�h�}Չ�������wk��ȼ�>�*�ZF����9����w3�v�ͷL\ ��=Z}^2mн�Ƿ�j�ƫ��ā�~��⺾Ñ�ws�Ba&��N���dt7Y3=��{�/_mD����.�_>�u��M��M�����	�7�=�Ǽ28��Ƀ�����ɋ37�^�^�Jr��ׇ��L�O,_ �Q����c�.��i�Q���c'���ȩ;{j��{�;�BBj���6�N��#2�"U��d�7_�n��ͽ�~&r��!�"�+�z������\^۞�n�6�qm�:/�W/"VP�5�O`�g��9���\�f�b���;�D^���f�1���9��}�z��غ���2�/-WS��M������Z��1�����uްk+�%�n��]���C�<�0N���ض�y���`���C��h5w�w�y������"Qh�U�m�oA�P��k~���K���ȓOaY��3�s����}hΦ �7[檋�25���T���ɯ����<�5��Z}~V�F������̪���ŵ<N�li^�s3P�n���8cW¡�m���Դ$�̑��/s�=.������|T��z�0��<�3�����Bt��xq�l�Y`�cr����܏�3��ȼ���md�:.%��]/�^�'�ş*�0뫟u�T�@q~�s�]���4�C�}M���XwE���>[eÄ�n\�=qT�����~����^׫����m5/NO���=�r�:Z����c��W��n��@=C���L�x��"�H�\�>Z�����p�w	�_+Kw����7!�s���2�w��:��H�?eA8���ٛv��`v�Z �Wu"o
��}PQv�P� �!�ji�w�k��n�9}̺T��u.A��s�p�.z��/�C�j	������x�H��h��QȼJ���֑Ͼ��g[�p��^�-	ϻ����5X���7o�E����/���,:�T+ŗ�2B��̎�L\cJ����l:9c�����^��qlQjT�<d���<��e��9��5���<���?��Y��p.۹>��4�m4%��ZҤf:�֍�n���jg�N9�:	�-L�ݳ���h7�������uQ��Ğ;���9�ia�|�R]k�a�)u��;��Y�f�$-Un�s����N|GI��y묛D�8��9�]p�����xzֳ=obg�yaQ�w�>v���piu	�4���HB�u��`��E��T�u�n�m�0 
�+{ ��{�7���T"�w�>�h�ruld@j��\�tD���'dWĭo�qq�ٝ������׹���	�"���]nvR�4�2B��weܹ��Bo�� Z�>^���V�Wv�����A�r�^{�
��S�q�+�7�	�o2ܷ3,�ߪ�l26�옛�V�{��P�qq�E��h��9p�J�7�zr4��L߳��Q����W60���r��ƞa">�(����5��m�6������;,^�&�����i�\�wӊeϛ蘪������3��/e?�����#﫸߾X�*��l�X't����*��}���ޖ� ,/`p�~u�iv��h����}t5���!>�"�-�}��ܤ�
/��n"K�{{$N�F���5�Y�+�/��L���ef>������S�����=�:���+���Whh_�;޾��zb_�%Q*,'�o�G���ed���U�P���urc���uK�M��S�|LɁ�^�C�ʤ�f��1w������C��L���
���qms�ی���QD�\�d�(�9�Ox�U���KG�3�&����<5m�vP�������{$��E���$�]&c��U�%2���?����(:��g�� �<��zs3�.Ԭu[��j�u+9�B_P��i���	U �gY�
M%NE���<69>�y>����"D���̍��Ƭ�Q�ہ�/�"�[�v煐��)
fw�)�MWaR��B���l�^v�wv��z�cb=}��z��ǐ�e������멙�:íV
dĬʒG��y�]��góOO?��Rl��:r�ps�1�gِE[�m��/��b�
��A��m�Y���{�3˧���N���/���zԅ�u���Jr=!��;��S��,����R��C�Q���������>��q~��b5M���U���ps`���t�??���T�n%�Ep���d�52�0h1���!T_ղkK����M�1���6d���7}�h��䕩��~�׹��d�5�T�̱�E�����N�f�6�&�)c��h:��]'��B�bw[��T�ϒ��7��wd�pߣ���ӑ'�v�k��+�*�;� �z<���Ru�Mk�_�>JR�]��ꕳJr���'��2WL(݋/Ȭ�3�Ǘ��kv-���y1%þo=Q�4��f��j������ʝ�G����]�.Q�%X�-:��Y�q�ܮ�=d��χd��\򂾔4m�\�܁jZ(�����������] n;��}�V*�{gL\G|'�ܖ���+��j�ݣW���ϝ���i�{�3�=��j��"r�\5[;p�/���ގ����J=��{	�#ߧM������`���C��[`y�Z�݈܈Z��o����!�'Hh8֝�,~]�=O;��'��XC��\��t�λ�q�U^Dx��,껏f�oF|��;j;E2B,}�R�Ÿ�7��ZGn;�]�#�6D�Q3�@��S�ꇹ)�����\���J�ʵ��7����:g�>��)��]t�j�(�%��}T���;̋�JBs�24i*�Ef;~��}�	�:�Wm����d�b�[�/E��p�8ԡp���gx�A=s�t�$�jvr���~�@>�{!���c���mR�����:��7o!�q�.H����x��f�m�go��%y�z�Pݮ�� >�՗�*T*t���HW�g�V�\���6��`���\�Z,�g~��h��/��8KGw!��7pn�L`y[#��-�3���@�qA��T��T�˘�x�}zw'&�P(Ѡ��W	�tM��OC|��x9�Z=Z�@���kW�&3ۆ�>�#�MK\�km֫����(G)�8�^��vo���H^U��e��c)��P�k��Ѫ[�::����3ٷB\[�g��T���K���Ho�D�3��.\��8z.�@%O@4_������q�?x?�q�	��3ԞX�G�Y�0����1���27��~=r���.}����,V�E�(���F�/��1pک|r
ʙw*�\�J���õ�+[��V����q�yӿHX�v<�C~�R����9U���+#"�H��uX�j�"{�+�K�;mZ��8�fXj�;����V�B���] �ٶ�f�+v��+��f}�����^����D��ohcFrR�-ж���	�N1�ꇂ��B��W�hLi���s3km�'#㬳q�x��7��s�c�K�Ԝ�3���g���������=h�f:��X��|�B�S;-v��|���:+�^��߉�2jp#���uGq�⸫�ݶx�$n�s���nMixN�1�:�0h�y$�;����N;�[���7�X���q�YE�<JF���T��\�Ņq�GR���>k��}��oK��s���w+�=ڧ�}��z._\{>��c�6&Q���*P��ٯ}T]m}���[Rf 2��WKm�4YDv�
�Uցr�#{:��.p�Ż����Z�uZ�Շ;�7��k��R��Wg]��q��h���=�uuz��kx�Z��g��[�\�4b�����*�E�ҷ���dy��_g��N:L��)3��	�T�)Нd��M.�}Nt)A�l:�}�~��{氪��^�>�8�4��ԉ��+��\i�ۆ�����wΦrv��b�}w#ԛ���y4�T��$JF���.)��	WH�+��%��1�N���&�a}|�:V>V��'G�����?Ihr`0��P���s �]/�*��+�oo�x�R�ª1j�Z�N�$~��s�ፙ�X��%�	Z<�0c�_X����]��R1��)���S�F������/��f,>�d�g&z�o0L���`�7+�u��!���*���%.p�I/���Vң��:�cud�O�: 5R����q.�H��RvG��u�Ek��;�^��xy����^����U�z_��]nvn�Nn!���/zWc���7	��/�bv_0����2>�R���;�nS�0���ϴ. ���1%�nr�(p�Wƨ֚a_�E��̲������e�{"^P�q�G�\���8����r��g�c���2~��8�9���j�v�4L�;SOf����·u��%�N�(�rok��I�B��f4 �ݲ`6�m�8^d+�+سyM�V;�by����Dt�욌�Qo�CsS���8*����q�D�2�<ð��LY8�H�F��o���kcT�J� �:��̞Zs8�`|��u������0}�X����,��l�w3�Y�Nb�>����~�v���4�\\B
}K�܅�zF�7[���ElC��-`��q%��L�mt���{9���Gvvf���Ĵ.�L��˞\�B�l	��OF�>�oΞgN��{�^d������7��w�W��������Q�1QS�	���9t�X#W:~�qln}��Z��4/�[�Ǭn�{9.��|��D���Rf]��0���]������YXG��;�9 j�I�S���R}��}B��Un��9E�d���M�Ri*r.# ��I�y=�^���C��}��kh�٧�'�9�Z\ӯ���~�@l׏H���\�M�%���I��r٭���ۋ��']���_�;HF��/3>n�¬f�
f%!�%GHa���5 ������+lU�8�1�ir��_I⫘S�_�'���Wp&�F���#,�
���9;��s�?*�bb�ii�%����:��#�%�3~������~������>I���������o������M��h��1��&������6��66m�ɱ�cm��c`���������͍�o�66m��6ѱ�cm�66m����1��&�����6��ll��c`���������c��v� ?�b��L������XN� � ���{ϻ ����7���(J �Q@P��R@�*�H����D�P�U*�@��*T*ED�H�P�D�	UPD�{q"�	D�B��*�$�"��@�I
�T��IH�[4�5�A
��B�$� J���ld٠��w*���*+�T�%H�*���
�@��H�"�V�l��T�%D!$TB�D$�H
��%shT$���  .ꁠ-U��0�E30�QF���5c ��TX���3 ١)R�Y�EeJU
�fMiH�P8  ��T��6��3M�53�Q�V:QE c��
(us��E(�QGgm�
(\��
(�q�E �gi**IQSC*�R��  dP9�����J� Y2��� d&� (m� �@(k@6Khl�@Qa��!C�  'AUu�b�6 Sb�*�H44��
���ƪT����F�ԕX)j��T)$�I�J U�  Y�[ji�m�h*��f�R�0ؚ6U6�HX�hh3e�[ֶ�3UR���Y���J�ږ*[[T�VYZ��D�UUR $�*�A�  'v���j��kfօU�mSE��V�4��ɳm���6�R�Ī��`T�cj�kT�X�̓j����T�SVD�%R�U@$*.  �"!R��j�E�SE���l�Ԡ$���U�j�Z�TUQ-ZҤE����ڲ V����M��Ui��PUB	JD���p  Z�@�k�J-�ZSjj���5YU��+U5���Q3Y��k��m� 6V�mVUKMA��*k*�RP
ْ����  Fi��MkŶ�H�4�CUZ��QSmj�ښ�kRh�6�)��VV�H��E�����2imX��"HJ%EJ��8  �d�R�+�ԫl�0j-�ZXRR��E�m#m��i�j&U�lUi�,R�T��2`     ��eJI(�� �44����a%EI @     �~�bP�d�P�F���  "��	R�1��FC LF�!�A��ڞ��C@� M2 �I*�2Lhѩ������6���E�Dn���K!��[dJY��# a)f����{ֿ@I!	��0�2HI!	���$�RBI ?PH HL	�8�!$�&I���������?��z�f�F2�@�B*�ʐ�IN$��Y I$�'h~����y�F��O�~_����$���O?n-��A���m�]��ƍ
��`^�_��W>�E�Շ� ��u���BXM��owY�L�H�.TW��,3�y�d��4;n�:�M�r����TC(]+"T܈�-�#IgqX��
a�9��ݠ���лjۓ6��P1Pݖ ȩX���y����5kbҙ�Bʼ�j�"��-ױ�r��3"�kqjV[Ѻc[@8�m`��n-�zL��"*��"�.�v(��R�Z���UkNLyuy��1{L}wzl�N;�c35�E$����t��a���;Y�z�[�.Q���4ӫ%	��q�s)�wc�Ջ2f�P��re��n���|lf�E�-�Vn�(���)d��.��Y�hmn���ٛYJ��%;�mdU�ݚ �of���a7�XEd�֘���Ȧ�E���A�͙����)����
�+�{���6<q�Kr��5P0�Z[�f�m��0�F% ��\0Tp�}3tn�YI�d؄n"�M|f(2έ���Som<`[�A��k�Yb4&��pR��f*�����R@&6���0 �A�����d�ɸ�ܤP{�-�H�!���`j��[��^ژ�eEX[����w"�8��0�٫�Q;�Y�-�u.[R�}�Ӑ$w��̖�ɉVں��S饖+� �k���M`b74�uٺa�ň BF�K�orZ���	D�K[�������]��2#�L�"T�KNY�!;yL\�)���^���g�q;N�{Iv��YY�fL����b�*�� т�L��U�3u��r����c;Z�"sa�wilp���y��,!�ӈ�3jݭ��0q�u�Oe�R�kbN��{�Lܤ�ދ��6��I˺'2 � ͢j]ހ��q�s���d.�koc��'�#z��e-�Pa�F5�P�?#bQ@�@�����1fَ��nΐ���6��"���3�#�/��J�����S`�b�n}�~E,Bن1����u�ŏ�:P��C
�!�_Z��Z�b��S���V IZ���6���6&��S��,aK;�,lfl��2�b`)��דe���[��6����S]*�z���vP��i�<Y�%�/7[�p;ݥu 4��l%��2Q�[�:�ud��yei��SY��ݳK2�^�7H��Z`'�-,RL���y��Z�c[�U�!�N8�+�-�ׇ�`���ACn͈ڵ�se� V�*�R*�ÙN��IP1�QK�H��N��������5�a,b��U=.�t.�7M��� mi;��<��w�U�7K��3Xm�5�%�)Y�������t/6ݑ����.���05�%!չ��[��+ @5����Of'��ݫ-O�fB��a^���(#J�
�J4hh4h3z��R�5R+�0��&j �������%rUf�^�jGEm��;,ޙ��Y (k���I^:�]hI'��M`��3��Z��̠ɲP�ޑҴD�;�����XR���r��[��d{i7`���o��d�ʻ��[a�E�I���ifb(��+�&k��s��'W�I{-��\;���J��C{E{�l�9{��י ��j���/!�ig\0�� ,��m-�UnS����SZ9{o���h���)��`7gs/���ޅi<��M�Z�l�[9��R4)���M�yZ,hWY�à���8
��,�҃�r�#Jj1���w"�;n��q�ܠ���)K-ʎ���X��V�%i	ٔ�;8
���taP�O�(K"��f�u5+��E���:�0v��ZA&ڡ�����#�]�\��O[����ZD�$)����F��ے�{���/]�2�%���GD��ݍ�V)�{�׍G��n-���X�3j��V�bowooHY|!NqTu�si�7�(	��t�W{daɁk��d٭'3bq��b�m�A"���*�Ce�b��U�
����m*�vJKe�wDٔe���mڱ�s�J��֌��8a�+6%�p�J��]��y3tw�9�rY�Ɓu��T�Q�&*f��I�V�Db9Xn)��v�"y��Z8U��p�v�=�Y4f�L��&
mۧi��#tm[XjM���l�&`�Yb��nSƶ�eHJ@iq}�����y�����=
�Q��˚6���B,���R�W���[����Y;�h �\*+ĳj�&s`,A�=j���P�*L;��L;�u�T�O�j�!�Ŧ�8.����)�!��:, ��7J;R^ŭ
�Y[H�
Tcʹ�F줬�	�o3㸦�ˏc�j��G����K2�wUcZq;��YDM�9�Ln��A.!2kݡ%(C(Y��Ъ͍h9�ީg䧵�B�v�fкM$]
YsGʖ�N̚A�uY��c�8�m S1�	V��VE�6�ٲdr�����T�v��%�]毠+C��K4H�9��`�7on0�� �P��q��&ks�nbU���Gp��кdP�)*�5�pi%'��Uw!�P�%J���c)Ռ�xPBQ�ǻ�.Y��	 6��劙�%T�I,ո�pjo�(�.KA{x��w%�M�35��Q��Qn�<;k*��)�����Z1 �OlBql��n�.Pk_�0o+Rbą sF��YYV�qai�O)Aw(`�lШ�pe%`Ō�B��6�
��8��CX���aa.��V֛a��SHh��@4����`�*[�(:v�L�LI��lV�l�-@��j���Ȕy��m�u���Z�{�ae^qB�ݹ�⶞X��Qͼ
&��sic�y�9j��d�A.�ǚN=5�Bl2���8�v ��U�v�
�
�m97mXV�U���!������pA� �{�y3'��e::6��`	ov�]j�����K�	���4Ƕ��Q���Dn�����R��;�H.�2r��z�B ��gX]j�I,x��9,�NU�q��X�[,m�EZ���T[3,Gt��Ib����2�o>���80t2�m:��)��
Q�\O/l�*�O4%��p[�2�mܒl֭7c�l2���l-���	��-XUU�/0���֛y,̴�8���v�1�"�Dn���n�=�t��R���b���G�]��7&}d�����eH!��*����U�
;XH�������U�k�Żq���ji���')��Lk�+�L�^ӇTl�sw�e�jhX�d	%7��o1%DPi��A���+��ڬ?�w �T�x��(�S�SSƚ��{[0��7,�g>��osj�����F�-�XĽ ���������,��V��2Iݷ���x�+�!�˖蓮��!���+l� m��l
R��ve)�BNڬ�ҭ �n��(3��u�*�]Z.aUd�v�QFVP�%2����Z˥9e�����w���%�16¬L�p!�L��KU��\�tw]��{��)�hɽu�O�2A%�e������[��X��W����cI��P��F�a�Bm�q�i��T(�#7�͋�i9M֓�/wf5l�n�|��hZK-ڽ�t�
(�0�KwhH��&8,��oJSԮ��K϶�mȡA�4�����I�n�����Y�͗�$v~9T�dy�YQˢvj#���ĂYz�z�$21����[�%��GD�kE�jOwA�V݊����e�)���&ڸnJ��]�0')��=Slз͢�*J��LI���U���X�b�YPL���W�r�i���"���ɵ���{���(֔�nZy5Ҧ*-�Ki !F����d+��$�8iLI�/^f�YEe�f�Y,T�[��N:u�P9fS7v�J��,-��76�1��ֶ��qf��Z� �ڼ�+j�e�6�b��,�GL�N�H�,��+w"�yX"�V�´�9�ƳC���39���*E�9��6�a`P�9e� ���ۼ��&Vl��U���̦H���;����dp�P^�-#R�`�ӻΩ�U��ȝ���4��	J͢]$�ԕn����*��Q�B&��c�f|��[��e��6�f^
̼�v������(-���x$P�6f�;ݼ��H����Th[5R�Gg"��&
6���l��$�8j�u��賂S�g7ՈI�SY��*ڽ��n*=�ئi�.�����^� a����z�l�m9����Cܖ.��,�%��W)@���� �[��3*]�3rE��b�6�K��j�n��0���\�`[+eց�:�͍f)�L�"�0^��7F��;�qJ�C�BPS~���h�C+c�����LS��Pa�; Y[K*�j<ߜ���n�P�I�-��kr�{��V᭤��j�J��l��B/��^PYK�^8��E@��Y���/t,��JOM�w@��. e��w������2ɻa#n�]�M3v��U]R��B�L:(��ojV���;{/p�Y8��n�H:�V�ͻ�z�����Z(���`�o-�E��bBQ���h�?fЍ�j�$�u��C^�f�h���̼��K;R
pc���SÛ�Veǘh/��u1-T�ز���.��Қn�G-��[SM^�a!fe^Z�Ȃ��	�][�m4+o6��Fe��m�V�Хa8���r��0�����:�VR��`��Lf�շ�(�ڷ�<ܼw{H)���H@v^�YY��mV�4�f9�+�CK��6�撵fS�`4ИsVm��M�Q3ƐNj-�A�∭�&mn�!c�;[J�d�a<YI}"H��� î�^m( ��$L�Q�iaXv-`��ł��\�u4���m���v�e�{'�'ה�:a��n�3rA���U��N�KgƘ�fڤL�p喲���S+� ����2��҄�^�������& T2��کB�!�eF村J. �X^K��\�R"CP��L����0�k�kB�OB���঒�e=p�
�ր�n���m�$N�To�����������ޓ6�k�@.IVHt[�fc׺�W��vlm��b^J.�;�(��]f��.3X�!�����א��4�����b����.ȉ
9e*(��y��@�+/P���øe-���̶Ўk�Tn���g �N��0�"�D��-X���b6L3F�j��R�B�4ڇ`^�-�r��bL�{�	32n��]��Y�����GQ��Z�Qb��D��ۖ�{u��@�ْ���ڬo�Z(�Z�v�����e�cn�Q�U1+b�r��k �ڊጁ>yj;7�o!-y4��	F���׸�cA$�o�AdNL����������Y�vZ��boe��:�n��Na���+F�v��s��]��S�u*��[O+7%F3],
�^��k2L�3X�:#�"��5xsVV�U���1�+x��n 1�q^��*kz5�!! l��G�]���M*[�OX�/h�H�$�A��ܛfMy5��t)��i�·6�BG$��T�l�PҺ@��ɂ$��E5Gw�P8ja�fh��ڲ�*t2���Ƶ�A�(��)赌��%��F��Qvp�Cp�;nm�]�:1K��Z��%[l�Bq$�'�:j�=tq�ص}�Ke	Rȇ�H>�6����[��9�Q����9��.u˫�����Y�b��4��5��(�Ѹւ�c�kTZ;�X�]4�y��V	�ԏ��2PRR,d[���3"�5hґ���P��ʝ��� �f���%��d�c��Ɲ1+l��ffn@ܔ�P�P��j�ږ��*�ҥ+��#S&�9�E��J-�B��ge���Wn�M�vS�B`N�	Z�״p+:vKd�2seƜ`�n9��4M2���e�s�F���,m�����؛��w���R���Ѯ�kܚʇQہ ����^7GF%.n��nذ۷���I��f5�m�I�@V]є.�TD�{�)�w��CUiZKNx�Ub�-�/mVe֊Sx�ހ1�iT�5�XMd��Eb���o.���2L7��L�-J�G)��<���C��O۷�5�Gc"S����զ�B���D~߯��wuDJ��%ڎj�*koz�p��ݨ4���c<����d��{�R�Χ7���91�*r��ލ� ���%��YwS�����T�q �a7�4Y�*�)ِ%��w�.N���#��4��9I˸97�{��tv����;�u��R7�ۺ��!��\_g��Kdۚ�;.u��ԟV歝Cn�gea�X���H�<Z�V��eݵ���34J�ivӣ��_qY�%m�̢��=�^Y����J)m��=�Y{j���rIi��*����szbV��v�a+�v�dʲ�i`�K2��1}L��*`&���ŕ���u#T����ty_^���2��T[����gV����LLQl�� �2˔X�5���
�\-;�e1�{m2�uC�^����TGo
e����ݮwQ�N���*o%�u�)v��-\�lR�@�D��c���R�*#:9[�!�X�Hܺ�x�P�;�uc"�f�X�h�x���&�'A�i�}�G�k��]��8��`�oF��:t�����x#�����f<o4J��r�c��@���Q�f�us�c)u�6�2�_"�;��,��۩�8�A��i@��N���Vǖ%)�N墸�ߤcg ����v~��P�)~'��L��e9�'�wvnV�ߏ�8�!ڳ�_!1�x/�.���M���r嗶�� t�<��Ǎ[�8������ѧ�NN�/Qm�mX�G5ZY�䧩�02cz���iܧ��͐-�9�u��>��,)���;��N;u�wB����z��#fN�e��� �ڹ{�J�[C���>�˘�u8����y�M�`V�#��`[
�@�!);���qd�SF�zh�\6X�|bQuƭ�*;\�3+i�]\)2𡅬K����k��/.��6��L&�o+#͙��]��_V쌹s�_d�"S����vU^$J��Sk-�Z�B���wbÏ�zK�tue=��B,�k��>��sZ��R������f4�s4��7����_"
(�d(�`WJ�����uR��='v+�/�ٴz��N��4rQ�_om��TW�Jq�k�3>X��阒jv��3X���|;
��v�me*��\��(ܖs��[�Ku��ȝ���L��M�m�V�U;�O��*G���ڳp���+���b�	��SV���ZN*wb�DMlWC�pݽ��ƅ	�^;�&�o�䀗�G�ua/I�^s7n��T��n��=зc�D���oQ殃�c�D��3v;ɋ����6Q�����S�;t�0�������'#g�t��vj���]�tk4��*W�y�jJU.}�k�Zƒ�Y:X%.߷�"�?!u����G(3(؏p���$���V����'fD�M(�c$u/3���iD����{�O]+.7y�%��sF[�x��f%cvoL%b)oS��q8"��lw��1�
��I�&s� Z��3[nK��+��;�c�-gM.�Nڵ�BAu���3��zF���1J[̞�%{x�jՆ�]Z�L�R5��PX����fc�ۜ�}�&5ul#{���yέ���Y��xp[�WeҧV���^p�n*�hc��Ӌe�17ڳ�ٖ�����®��w�hm���Ί�|���v��m'��L�|�(]^KDR���{LB�4�v��l�J��/�;e�*0��^�8jZ�o�����u�\9�k�Ν�r�*�x�̬����P��Q�7����&T.-Mk椛�;��Xi�(Xɂ�u�s�ʙ��;���;�`�l�9�|\3�-��YҊVmK�S�-��{���I}D�����r�{;]�z�b�Y\cg����7D��ვ�k{Kl$���|�U�S��f�XVݵpo�<�R����^�����u^]��pA:�m��JYe��w#���H�Պ��Nt��3Bz%C�Y�vM��/i����Z���Ԫؙ֛�v�i��5�Y���O��Da�2B:낛��]�z����敧��̦�yF�ѣ�OS���y�,T��z�[�Ǯܜo45}ݢS�v�X�6�Ui�B��Kt����kf�FC�Y�`7�@���6�EZ�Hw
��]�c��֡��o+�_._(�F8�oN�y��j�P�QU���e�^�H���B>�$�xɬ�F��+�+�+�زhgN�;�ʶVG�� �Vt�1N���{���v>N�h���eZ#��$��T�h�Z�\F�:��fO>v�О��SU���c��R��oc��7�b��Nq�Vp�t#�W�ĪS�i�y�e[�(���le
�X����>��j*�Zp's$��N*u�Au\�B�<YB���hR������]�DԺ͵;Pq{2ٖ�Z9�ir�Cl�^� �61�\w���1̡WS1g����ǒ�k��,;)����`W��衏�r=ԕ�����J��f�rg:Sl,P�ε}y���u�·�:���`<�w�����9Qܫ�F�y�!���6gT+B��<<��ڗp�GN�d�9�,���hˤ*���ͽ�����+]�N�[�}�����8-��^���]�!W�qXfcO&f�RMO�V;n��2�xr�=��IP�{�t��Y�+9:�2W]��j
���w����95���&�wP���ݝ��`�;�̷8'�fr;c��W6��MAx��ZUlU�o�WX;�i�h\�־�G��V�'|o1U֣��!:P<�g���[!Z�W��`�"��ݩ500�p��S�l[ȹdɎhϥ$bCiDէS_J��=�`5)�X���Q�͞�23}���4���H���7�Ā=�7��,��dY3rnĸ�U�[�9�jgW�7k�96�0��$C����[�e"��ܫ���(�0W��nt��5i���Rr�����J�fv�ښn�l��[шS�#6����\*J�7��`����Mߜ���pe
H�ZfGJ�������79g1�o�������-�����������.^=�����d��c�=�)�7o%(�uaDN��~�R�Ѵ�w��NO�]��s���Fr܋;J��DyBiY�8�w!0ӕ-mf���e�u=��#�)�V�y�mՐ�\x�4'b��ͼ��3���}�F�� z1��hÎ�:��p�p��7�٥���$��ϸ��΢�]"�NyH�Z^����";xMW<�Z̫�
Ô@<f����@e�ߍ-��+*nq�G ��F�5ݑi�&��.іoxL�������т�:�'7Yr�$s���W0������A�$�ս�6&&N{h�KC��P�^�7�H��j%�%ު&���{��̼���]�Әu������	T)���%�v��me�W�n���EK��M�m��nLz���<����6|P�ǋ���2�T��I6�;Y�q��sT;q��P�2��D�J��u�%q���H�hĒޝ0�b54�u��+�re�]З���)�F2�,�(7p�.:aݍ�p1u��l��8����Y�����}Z�#HZ�H��m���N�����S�_>w+e�T�u�Ԯ��3K}k�ыEt�Jf�`��ꉟ>��n�k7�+C�̋�n�5�B�Qh����u�.�`�dy}��#EX<]��@(�N�g9�E��t�u�Ъ΢d$p<���dL���Z�� ,g�)>l�)ޜ��|�gw0&��u��dm��h4��y�!��5kY��5����F�Sgv����%�B��n�s�ߺ��q.�
H 
�Ю�`6~�\GoPt�m�D�0CJ�e��샦������ήm��,Vӧ���k�d��ՑV�;�Kr/�h6�-�K���v�$pΜ�"�,�#�h�uT�$�cJ��y7���&��Ҟ!�J�D ][��U�ݱ9����7+a�g��t�8�p�9����Z!�&��� [����܅U��: s�Ա�^:o����0
{C�nSy��̙���jf�*sڌ5z��!��P�</��{5���"_#��n6����mm���\[4�6u4��8h���*u�R�N���.MxNL=]YN���c�9��q<<:�u��pj�\J�J�� ����+@���T>��[��X:����¯�.�C΁uq��.,[�YZJw|��ռg�v��%���Xh,�\`[ԙ"���)��CQG�5��*�6Hy��CULZ��K%J琏��vr�����T�_�c�Ǫ8)ǙЭt��3�'1R��������!��̔�f��^���#o�7]B}�@�3>�ɮ�jZ�Xj*H�nYk��\-R`l�1u����;ULi{mh��i]q1��e�쵠 *�4��ٍݨ��xN%*�jy uǘF')1�r��b�dRΏ�s�heڠ��t&mbc�]r����*ϱ��b��=u���<cRM�+5il�\��&Zްo��<�s��Xp-��o�Yݟ^tH��'�I�߻�@f���U�k�Ƅ^����e,QR�Cs�2 �]M��+�&NPYy�c��誴���DT����������\����T�0��Y���t�!����Y\��ُz�u�c^�C:��fʢ����CD�i�]}�IW��s(`�F�TW�8�J����;5�/N�R��i+eY���Huq��,�=��9��
T�������GJ�^8��_���ݕpƛ9�X��*.V$�ȍ#�UÔ�R�ϒ�����m]�%U����&h�ޛ�Y�"�u5��cUJY���d-���έ�;���̜X)�hlK�TX��D,�����������謲ͧ����#?n��K�1SW�#�V�y���3zg3��~�zCC�-:	�V����j�p[�y�L�ɖ)�ʝJV-ɫ2jy)�'bO[B�u̒�S�����<���|[o���ըUs�4�����/�mD�n�u7i�O\�8�E�.��=�I۰e"�
�o9��.ՋG'>��z�����M�S-�����/�ѯ7�r���-�ԛAb�^L)��ʀ���l�F�t%+"�<є���O�m���t��R���Zgm<Z���t�%Z7�h֧�Iy.]Z��WiulzWj�W�Kfmm�x�5Ls&�fF���_U�	��u�M�8�S�����'c�uq�� �/o^��9.�C`�چ=����C�tXX]KY��Oz�m���l�|�I�Xi�Il��4�^[�J�Ql�(<��e�3��z2�GՁn8]e\E�/3��ᮌyo��vɏ.TZ����p�%� }H�}k��b��ѧ�;*+đ{�p�Ԟb�"Ժq���;�	3�2V�M������;�ugc4m��-�#�ZHe�ͮ�ʆTR�j���Q�׍��|���z��bjVA<�N�9�t�,�ܭ=SM����&,�-�XJ���&�ʹ×��]|+a�[�`bv�W8�$U����oz���*H�o
��I~n��)_�����s�G�&�=k*\N��] ۣ++�"K�������v�V�E�9�`�W҆I�G�F��I9�Ce �yV_ RK�.�6��L�Ź{��d]S{�_jFo[��.qF�q}r�k6l/�������bP62�3;6���ԟ'�R���K���A�/��5�ݭ�Ч0(���D�>̾�]y1�{x���4��m7,TZ��� ��Rᴩ��53��Ip�ǚLޭ&�}y��@k�H�\�2�ٶ�J������ջ�7�[�����X���nFWb{��,ǔ�6�nn��dd��W��q
[[���zo��s���I��kV��d�,����u|;�����]��o;�Z�벻zb��v-I.ܤ�R�)�X�bS+'z���vZ����(�:����n���v�a1�z�=����P����
ݤ��Y�^��Օ�J�,��p�Ml]�d1WT�k�WKPΐ3ǞL�f�i*8�Z�]�j���Lt�+�k#aַټK�;�G!o��!��̺g���p'��z��g�޲��.Gȹ��k��0_R�.$�C/�v���GLAT瘧.�	�5i�%3zmZ�Wm�7�j�xU�x���GP�zr5F5��&�}�c!����� - ���&�,��N�"���=J�E�VIDHI!	������P @���e�������BHBa��<?�����������ν3�־�_+���v�Kv�o�]�Q�����hf�ˇ��#��,�f��n\4�]�2�����X�%P�c��v���=6�KĘu�R�������UcC;'ٰ��w2�|�i����.�m�:\�*)Ư���{����r��б�N�홠�u�b�t�wsa��8��Y���g�ø���f+�n���)��Gj��v����3�x����^Pj�E2��c�V(�b��\�d�i�ۓN���ۊ��yo+�W�6)�-J��� ��&�d��ZNV��\���E����+�~��J꽢$�ܔm�4$h�	����V}nQ��e�xm��>���lj�<]btӝ�f9i�Bt-��طR���%iR������J�a	�8�7{P�T��Z���ڇ��d�;ѷ7B(*S����a��ܳ]waɝ:�y!�/�5}��U�Mꃹ%��'�[8a�{��9����S� �*c�Λ�e��VaۈGu�Š��K����qn�9/.�f��Ef��V��m��U�:�9�^ol���a��yxl9X@��o1��dXxb��^�
 	v~�y-�,��8j�+��Sԥ�IUΝ�/e���c(��;A��Yì�bi��e4A����b,�Sq����SwZ ��MΥ��ɹϊk�O�}�#U/N!5R�zVbH�*f��_�cFj�V��'�;�{Ǔ���k�f$̾實��������;�@NWv�kf���ˡE�-[� �����,R�u`�s��0M�]/$F���=ǳ�Ta���ܡt1:��࡜؝{�GKK/�玮���v�QV����e$�+%���f�,;H�8�j�/a�6\0W�r�[huLU�z�LY��%u�K)�0�l��lbI�F�v�oîp��/�I�8]_u��&�\v![m�X��H���L�۔X��4�MV-Y��EV�!�э6*vsF	(�2zk��&�e�j@-������Z̾t�]��$l3���.\��x,L��!��R�on�P����M�����PAB*p8]�Z�7�����U�HM͂�W�i��κ���Fl�u��˅it#gu|X���-�{t��K]YNn�SIYJ�m�D�`�/P�0E0��;�j�1r뭧z�L�h����i
�I+	"�`��h��{e��̋�gu�Z�YZ�<]�����9���˖��{:^^��tcI-/L�:E�jʡ.�Q���V�y�XlF�`��[A}�Y*�w^`�Qj����A ��萞y5Y�JP�R����Z�Z�rL�"������$@���U���	��1�邴$��իB�n�52e6�һ���]-��XK���s�Эs8�\�2邔��e^J�Vեz�"g�tNT_�6��
ez�p��wEk�	�][��D(u
;l=��h�t�}5��;���g��E�5�7@�\)l��Zp�`8�ݫz�O��dUc�yZ��|��.��q���-���y�塃5mr�O��
ߓ�㕈]&+�b�܂��	z��޼���P�3�y;a�[�&M̤�lu�����}*뺲0;M�o"�LC�9v�ˠ>h}��#MӖ�S���Mk���%`P%^Vb��*<�f��jް�y$�4�_S���Zyg:сu3Kv�����BibU�t��u2�T�vΠ�tu����h*�� ��+�q���/�|p�4c�k.t�Gn�'Z�̠���H_'6��v��T6��c�)���N���h�`��[N(Fg1�e�kn��Qum�u!�yo@x�RY,��n#V��̴@�=���]�֤�5N��X.�5lʙ�s`�����b�����'�9�J+�:B@r^�vC��V=�]N����&T��[u�g {t�U:�Yf�S�F���Pe�щ�ˢi���s��*��n�a}��wGD�}ܩ��gN�Z!�+4�j.��`U^(qԄ��H单6C�v8=/��F���]6�T�Z��=�͗қYz�Ⴋ/��sG0abʮA�/9��R}y���1O��&�(�VC���7��S����(�����5ز�mr9lAq�;<��xwmC\���7\�c�VB�(��0�Gx�g�R7�3�}��w�սV�)� >�ʚ�9� �/�4��w�Ks�Q�ҷ���5�[n����;曠�K��DB�Lf��sV�R��CL깦�Η0��l
"��	�G�*ͮ�N��w׵�[����L����,"!�D���ŭ:ѭu�){VڹIțg��W�^G�m"),���s&��R|�t��T�΋�8��+�^�N�R>V�C\���y�-�[L�|��*�맩�9��{����QSzf��7d4�`�j��6R��ũ�HH�AZ;r��̨O!j����'y,*uբ��Uo;��e���&��V)Ǌ��Ƴ-�@tnbi}�av���6-�9�G#�\�7_l3���Cv��ɫ)j,x37]�%_3R��8�rŝ]2��q�ZT ��ֵ�f� ��,oOGu��o>�=�Ե��N��U��¦S�)�/0�m`���:�ALw�W8��{��@U���Zˋ�.��|;yl4y )m�9Yfg^wo���F�1m��f���MgE����x3�20N�/Zf<�愦��(]��z"��x�6��+Fp���V(�,豙�s\<-N0�Ӂ��	���$��p-�Q[4[�h��e�} �]6���^]��rs��X�ŋ�����Yt�3�w�y3E	���fu�²�,��&�Z��ܳr�55;�8��D1	�̡�=N�Vٮ=�L��(�06j��ĺ^�~]d�գ:��v���@Kvs@���
�̽+Q:��uh5u�B;f�jy7K�A��E�3����ÒU���z�%�{1�\�d����ZOq�Tλw ��uU��'o�,Ϛ� ʐ���wB���MN��%V���p�%��4�C5w@���t
|NQ-b�7&���t�W.GBݼ���Ma̾��vNE>�:�D���I`�����ݩ]��]bb-���9o�)�(O������y&ɦ�_m�c��m���Y3C��v�����N7OxNn�mmS�r�㝥����VQ1v���	Vh����β����ۃ����{���6��i�*�-��{>��R�!��;R
���	�n.)��-�+ZLruuHv]]J��P�t�	�vh��˖v��H���<�M4�N�����9;��Hb!��hXQ�K�l���xqi����Q�)V�.���b���H	��j�%�A�h�����=����R�]�S91VD���Ī='/9�*"B�t���x&rԄ�ґ�Fp�ulz�8�qk;v|���>|^ҽ�ɴwt��������O�����G���B�Z�x�EC/r��k���V��Nŕ�ed�_�n�k@r3y�1���*�Q[v��G���ląmȬ��Gm�3hj�5EL�`(Z0y���[g��5�J��V#V��9B=�9b쩼�����¼i�1"�.��"�P+E]��h�3r+<���hXYsĕ�Pu���Pf⨭[��K�u[�S��Z�
M	��<����V�
Qv�zٷ'gVes�.
��Q�D�Bf5�(9�H�r�R����`�	5'na�t�]��Yczm�����i� ��=R�%�oZ�bi�u�jE"ډ�-w��l�8=��p��i�#��U�������{�ݍtp̪5ɕ��V�>D�n�;(�X��gf�"mq֨�be�[q�Z��gm��B"�p�ӣ���M�&�I6�e!�6��sw�%ڢ/���Kd���JGe� �Uk+`8�)�d倍"TD�t�77Xz���7��V.]k����=�B���I�2ZܣO_ss5ȁ�1(�Ύ�0e7ن�mJ��m�6���m�'���ȪR	�.y�!@Э�^�Hq�X^d�孢�ʌΈ5�3��9h=9%jt<N&�+�-�ϸl³WTF�v}��Yy�����t�dC��Y˗__�ISl�؞�u��q���/��t�N����S���O�=r�	Q��S�W�*�F�}����[�V�H���׊�ok�����CkX��b�Z��,m=[�Z��829��
��
v�dwV���d�e��r�d�d|�9�GX�t��.�kf�ܶW[3�,ݬ"��Юx�s�MW
˛L��g��6��0���+���/��u]f�t��m�=��I�ȍ&���)��[�O�f�YV�7�VVj���t#
P)�F5D�Fu��49�Vj�ĳ%��93bP�%I��"=�Qk���ZW6\�TScѱ�7�	��ù)5P7G���J��K]��'tu$����0��KYL1G(�++�
[��9��:.�n����)Q����D��猺!�;�	���g�;��sF]�A��6�hqڮy��lὊ�Bݝ������Y ]G��5Mbh�9[m#��� KV�u�v�]�;F�����R�ҳ�],#���ee�r<)�rж��f��j�.l����H��$Ӵ+je�e�w����t�|U��=�t�{qk���hX��q*�|k�'R�t%8�I��I�F�b��1��N��f�@��t6+�:L��A���*��g�C���N3�<攋9�ۛ���Z��n�GPU}tE"oCv+�#����۲��U}�I�0�
�yikz[�B�H�_Nv�7�ѶȒʶ��Ş+yv�ZN#QN*g��;�X�=��K��s=Rm�P��#��L;�Uk��H5.���m'�U�zI�F�bUɤ]���cZ&���etF��h�m�h��:��CF�+�N��ʺ�I�栍̶�x*i�s*rʬ�]�]6�TŹ#�t�d�2� k�WFk�v�ܨ���R]�
�����\I#��N�2Jغl�]���5�28N��N�D����v��+Z�Pnh���.v]�ٰ厴k�].�� lW6�R;���Qv	[���y �`���%�P���$*�s"=�i�ֺf��kq"7�覐�L�mV����v_JM�6�-���f�]�x�rж[�S�ݙܪ�����4���ݝ��;0���b1a\�[��.���>v9��̖(�ôWQ��1BZJ�t����aŢov��|��vҠ�1�lgGSz�We,���:�U���]͋ޤ;�H� .�D�+��<F��v5L��o#tࣔ:M��0WIWI0��Ի X��u��[/l��E��ct�uB��A��ݘ9���q�b��=[�v�=����5+&����s��J���)�`/e���$G%�tLNPei)�%]2��Ͱ��9��ub��ڢ4��Pu̔@�ntM֕��9�!me�5SV]l�jB����n��(I}�8_)�,=�:QL@lX�ٷo�L3h��j�F2��n��T ��9���cP���:s�
̜z�V�gS��WXw&���9=\&_d��݃S��Ϻ���
؄�0��3G�ǮˬW�pd���'!}m�u+�y�m�n\�"��b�V�S$�6���%���#�{�˔o�5}d���|�����<���}���u� �d�؝��<^��ON���.�Zf4V'm U��Zq�*���z��9�luݎ;���,SX4�COʏ�qG�@�t|u�&k;φ�t&��f6�4��u�˜/�)��p�eX�8XѪ*�	Rk����3{)/��7����4��f��K3�J�`%bi}��P</�tpw�ŏ�,b�jܷԸR�Ł��U��*8B&��B���]{�f��P���@��)��V�,��%��=N}x��;�P�NZwZ�Y��b�CH��)խK9˙/���>��n����`��s��2��k�
�-
A
$��\�+%�۔bA�XjĽ�e4��`K)�V9e�75+vy��|{a��Gնz)l��&;]9���dwҮ�����#E��Mх�Dt��G�� lУ�LÒR��}j:��l�/�{ϔ�940L��B,|*���r���.�ѳ�S�r?~{����߿�z�Ο����$��A��P2L��Iw�\��Q��y�9�}���z4s�<�����SP�al�I���L�Ǎ�Lj���I���O7	�8���B���Cw��́2:�m:=q�0ED�q]S:�����iy��#"�o^�E�&d,� ��c�Ά�*�(�v�WB��Ut����.b	K�'�]c%�(�z�p��u�ّ�FQ糛It���7���ޛ7�Aܴ��G1�4+��q�l�;�L�{�-^J3-�@�z'(2��k��;�|��i.tYA�� uxʘ:$x:�6�X��ˋ�fϯo/a=&R)c�|MNuvre6S͊�gB[�7���PX�{8b��|�nV�U�"�<j���w_M:fVop��v��]$�0�;j�{w��Y�|�Ppva@oNb=L��r�ޢ���Q+t�48Co!X�s�jU�εQ%׈�{x��
ιZ+�bZ&R�����)�i�zW}8e`���=��Y�`X+�4�*앏C�Y ��l+Yb��S��ϲ�k�V���r��v���#�JK������Y��C7�\�0���ء�1EO;�1��]a�����c��*^i�ιLu�*1Jۇ�_r�YGZ˙�m0Õ5-��nR�\%Mx{��J��:�O$��i�rk������ˎ���:8����x�>���)��S�x��\�_7ݕ�^�]�=����}���P��QU�h��Lf(�ц�]dƍTU�������pW�c�UVe�f\3-M%qU5j��,��Z�SN$�e
�\��UPz��Q3V�J�ڸ�B�ke�*�ҵQ5d�m�*���-�����j#�11#R�����U�UUq�"���q��iu��r�.h�Dcb�aj��[u�4�b�Q�,b�3
[�1�����mr�k+��R�QTE5l�+TYDY����9���.��&�-�(,+b�-]&"���c�Աm�Zъ+Z,D�5e�b̵4R��#�c��(�-lAQs2��iJ�bj�U�U���W)Ub�h����Q�QP�PAn%�W�8ؠ���&�b��Q��5J%qʕQZ��!@r�������=^k?��'���R����v
+r��s'��s�s��1v���9���JBJ%���z-�%!�?����'���je-���R�q|�ӓ�Y!�
�wJ/��fuTv�F��}�*��ۊ�#�Du�k�[t�ú�L�<��{'��7�o+�؏�� 4�]7 ��P������ay�&:nV�F�p�����&u�p��M��O�;6��-mC
�T6%P�qN�W�I����6'y��;Z���7ڭt�m{tB��J�W̸�f�j]��B$���4yu(|�u�p��օ�c|��w�ѓ���U��%���=G/]���V��^�G=��	=���ѕʇf"%�Q�ұ��F���zJ��B��g��r'F;���4w��+�=*#�S�R|j��޺ʢ���@�@�7�*/9�{��n��N�/E`���V�;�'1q��~�� Ѻ�W	���V8.���Aom�5���+�Ԝ`	��s�U�N>�{j�hOm�lGA=[��bw^a��Zw����=�;n�]a�P���i4t �fR;ҳ�/��+B9D�p!�^U���CX��X�-�� ��\u�mk��"�j:�e9=��J��JÔ{C�V�<)�J*�X#�+�������9��1�:�_��_
G(L��>�Y���E�[l��g)�Ҝ�u���{�ܷ�����@�n����t�0闘�zsno���db�9�O-��J��X��!�ph�rw��Ś�i�w���F�E��N�܍R���7��^��
.�{Q�Ly1��;X���oP4�����⏚G*����VvF�����+9Hu�(r�HlO�d���DP<G*�J���"���5K���2�5��89��!�yY;TU�p�ːrp�V�3vg5b����;b5���|��P8B
�w���.�3��f�秮��ӡ�Z\�22���Y,�j��ɭ��L-��Ah}Eq-�H����w[.����3��ͦȴ������Ԕ:�*d2�jP��*��
{�����n�0��m�%�wS���({�fPG�㣽;!V�[����d�99�4cK���9��P�}�}��\��ل,q�Y[��U9B2�/w����'q�onP���'q�j2����7�ܜ��ݰ�꽘������dd�t�����uec�ڜ�ng����-�wS=������|&�Ao.P�m���R���]�e\��<5���o˞m��ݬ�V+*���W���S��=�a�KK[6�d1����:���m�&��G����f	}#��{���N�kȹߊ��k�{g�!���u�3�5�9\�3T�Zk.��&�,�;�Qj;)Si�S��ԩ��ؖ�n�l9����K0O���u��s�����s�[Js�Ð�Ɉ�Rnk��I�a0�h�x��*��w�^�KNpŹ�z�Bٓz#FNI/%ot4D�Y<���~���a'%X��٣^�z3q�}�W�2�O�=��9U��UNR�y�uL�$���7�z��uqCC;����k�:Y�G7���h�z����`]�`D���8���`��r(�]�;�U�����8���G*ʨQI�t؅�~���E&bUc�?fi5j�R>m�)<�@�'Ä�{E�Uz���X�v�^1�z���6��]-�h��'�;y0i8�&n*�-0jSG���o�g}B�r���vѡ�	�H�a�50r�"���yWS"�?oGP�[B(�E�G�f�yH��ޡǳ7���|_{��/�C$�o���"Mӻ�[xe-�T3ֻ3Ӑ��OZq�]���%���4`S�DN:k�y��C9���i�uj�ٹ=y�Qv���;Џ5�8Ƙ*�}a���7Gl��6���5�!g�>��^�1��	<J����n���E�X�q��ƻd�@toU���1�FiX�C�Fa�@�d���8U�3�9;�)��z�Yl�;����ݜG>�NK5b�R����`0��r1��9�p9���:`����ZRju�,Dg� ��-��fz��v�3��y{�:���O ��d��p�ʉ��N�&��>��|�߂j���F����W]�&�Al
�^�T]q�Η�ɕ[3�>qt{ܮ��T�ޖ�m�.�A��.n)��D���*=\e�Sr9���mK}ϻ1U���z,�p�v�?A@��R�[���h��Ԍ�}�4Y	<�gӖ|��,?o��(��=o�::�$�������x��q۫���P6�� ��KG/ԞH��R���;�R/6�-�A⽷��\t��_;�n"��}��0��L������)u��]p8�a��zx*����9z{7/�rp��1�1M8A߸U�.f������k��2�J�F��,Yʝ�c�b�9��C7�W*�H'�6�}���m[������xy���fY��@.�.�ѿ.u�L�L�϶�U�&urM��}`�w:�M ��Ng%!�%2g��*q2�s� ��7p�V��#s���Pj.b���¡��&�y��I�otڳ���pݜN�j������Oa�e�p���"��Ј��C+�V��j���/����6�#-�/;Q�Z�U�R�W�*���6�c�u�y�(���o8�#��z����w�v�Zr˔��R�v=2������ZqB�tus�\��^>e��r-h�E8R����O7�siwX�<M�N�����9g''�A���&���n@�bz�:�݊\��Ņ��mu�OF�y̻�9����䭍��z�t�l�Ms�M
$݌���{I���(rҒ�]��C�\�b�"��y����ѯ|&�xz�?tHWǹk�*�N8w����s-'����Q�P+����MD�;�f��dh�[��Z�"�e:^Z��<=�v���ʽ�,+����p<�.\C�\�t��4�Q��gL'z��u&�� z�HQ�$sL��#2�V���T�7�}V�s��ذ�}2�o�!�N�]�V�^[hj�w#�AB�����RC��+;z�C41�[j��_;�<㒼ޥ����S�"yE�8LlX�x���=G����׆�ei�ͻL^ه8��'�'��lxu�j��Ÿ�D���]����;*w�25��"y�c��yS�B]{��jf�LH��I4�V�(��ǋ�Bu0�3E�>u���lo4e�6�W����Ѫ���-�� {a�7����ѯO#�9���N���]`	c�dI��t��B����U��T�v���i���ͦf]_���`s��&m�o.�ЫN3��[ӛ����s����s4��Ί�>���u�^/KB�b̶�u�DO%;�N����ާ�����s�E������1@��9R���e��>=�geՇ��]D, )[�t�U�
D�<~�y,D�!�I���b�]����;<�����]�|m�Wm�Ts	�;"z2�+����)9I�a���	��Ң8�������GV2����!Z��vc��+im�[����Ջ�����v�j�"�\�yXR�N-��Yj�#죏��2�\n!~�Zg�8�FR�8@�;���o����.%f]6ʧ��0Lw8"��_��<�G"}�b�ٕݨ��z���;���8~��A�B΃���lq�b�4�m�E������i)5J`p}�A8�؅�jI�&�T0`#���ȓ��Yn��y�Ԉm��O$R�{E�4�a(�]�����b��������zª�y'Z>�O�sIî�m�8j,:�V��0Qp��U��l�8��a	�#x]�÷u�;wO�#��v�5m,UA<�)s�^��w�+��Á;�&Sܛ Gug�mq�-��*�r�/�#��W��� ,��"؝ck(.aC�q��voo�+���ަ���D���/y!��"N^��l6�6�7��$��*������ҵ˵�j���鷝�c}g�89�h;��lM�eGCMwE�r�S��'�V��X�^�C+:�����m|�7��eX}0.�Y8�O$n��V��l��'����}�ڇ�SQ>X�--2Cx�� �#�VVk��Uώ.�54�b{`Oi�rPB��o�75:�7��8�3����,���w�c`�s�P�h�˧k}��%��5ŢX���_�3W��S�m	F�����[?Ic�>��" �A��7������Zdl���\D���m�W���{��R��t�9��k�;~�\^��fNS�רn��Ê�Y.��$蓍]X<���
�P��Dv8�IƳ��X[w�x�Q�/yQe+r��B��U��dی~�y�����lz+�)�fn�f��}F����j�����omS�������<��;sY��j
���$�f��h���JGޒ�0Y�o@�����-�5�Po��^���B{���6����"�k:#;
���h;��!������f�}�Q�w���/�\�6Ѿ�GM#�)<��M�[\N��w|��U�����M:��j������b�klQ�&щ�j�$^�!�:���J���VS�3�_[4���<�g!�a�w�N��1�i����&���Xv����6h��rn1�Q��,Ws�K{�:�!{�;*��S��,E�֭���w#Xs��G'�,-�m�n�}
�_Gi��j��6��D�M��SǬ�t����-��C�!c�k0�N�m@��!�ٺ��X�����xl���=Iƅ��Eׇ6�f񻘩�3�7J�}KJ�7���%���
�E�s����B��‼]�fv���S��G$��oR��ʣ�8UМ��
q��4~��}�W��1r��굨��с�2֬u+���7�W�c�&�w.+�p:�er(����E���1�3��y�u��_f��
�t;%iһ���!�j��h^��,%G3'-��*t�X}�=md/���,�r�Q�.ͫ3���(�2���ry1B�qT
��� `]jv��]Wy̝}Wu{��)�Y�tö�����Z[����9Ykp8:�����Nq��y�JFe�[�*˝T�(�v��]�Pyώ!ԕ�;2�3ۙ/��X�4�+׸W��u'�QF��j*Ž\w.�ኻ�,�J�_[ˢ���L���r���'AwefsBK�w]8� .��Wm��ݱ]�"�� �-��pws�gD4��+�_!Y�i��U�������>аX��6���+F��h���ٝ|�u2�d�2���~4�!��:-Wx��IckU�W���#����� 4��'�^��v����B�j�:��Gy ���r�tO�:�.۳�f�Hk��{c��fެ��hΥ9��ޜ��FQ��ǫ!v�Xx�ˬn��z��V����B�
'��&Ƙ�f:ʕ��2�bSy&�p�=R�ޕ�s��%g{UM2-=m�8�q٣�d��!���r]�pJ0�NQ�+(kN�x�e\nn���]`An�X�B�N�\�����$8
��u��Bg4�)2m�J��qv���V ��P�����$�o�Ub�#���oF�+]eZ�k��f.����T�rg"�C��M�
�	���hm����Ź���3$�g'H-�&���pe
�+�������m�W��p�r�lM�;��q5� GyՑuw�1S�d���J�
�m㴌�0���2�˛a�T4`�`��4�9��F��۱v�����3�@�Q�
�t�Q�;L#� b����r�R��֖B�\l�5�b�����-�G>��ISb�ͫ�ff���W1�v�whk�����{`�w�U, ���S����v�V޷/�{_��6لD��;Q=�*;E�N���t��n�.��ȩ6Hֆ��uZmڂ�L�q�V_�\�xh��Rk��]����4�ɚ�j��:Qxb_%f�OpC%'o768T�s�D�Z�<�n���F�2ƌ���̻���˰�uo�'�F�%,&:ܬT��Z�1��׬��ur�����v�7]LT0���Tj�'y�\z���'@Wvw7����8l�)�W*��n,���>
�%����|/�H�i��4��FG-Q�X��{i��w�)wy�$7��3�[�$�v9�9����)q��a�d�f\��5��������J�VY�(��Z�E���*���-���� ��Ut��b�i��NLj+j��ֈ�t�bʕEF�"*�#��Ɋ�(�Ɖb�ƭ-J*�*��V(*�5B��ȩmq*�,1���������E��i��TA�Q�
[b1b��L�(����UQT �"�" ���!X �eu��0+D�j��,*Q%B��-1*��"�ڀ��d��4�UAuiV
���ˊ��Պ,�.R�$�Qm,Uf%b�0SICIb �֡���b���R[E+S)X��86�ITM[��*���"&��a�"
�W-`�*c\�+1&%Er�����,Seut�"5��D1��ab,m�e(��*1Ĥպ��3Y]"&�Ɍ��UekQ_�����W����?'���ud��x�eGՓs���4'O��r� ��о�1��
�H�稜�'��c�X�;9�ћE�얰���s��>����x�]�	kӦi������"�1��qJ��2�z�'U���n��RM�;��1�6����/,�J^J���H�������7k�.s���GS�K��t9�^.���F|����$m�ـ%������
s���.&-EC�b*��${���N9�/:Ĳ�p���7��aj�����Vtu^���p�	���q'�'��=OR~�j�֤�!(�ᠢĬ� R��鎑��k.���Ck�����;b}:�Ղ���}W�R��;����w�}��z��6�{U�y���aBvj�(4␗\)r6���=�e�ǩs�<i�d>��~�.�C� ��ѓ1���A��NI������4��p��FP\�9�O"|5ݼ�Q
_.�����Q u�Im7޽��3x�Yʪ�87�����}��bU����ȭ��|h{����B�F��N���f>�ށ��.ӗccjn�cRg8�*K��T޹��.v�Eq{�a�̫5M�Zm��/#Z��7}[e3�l��*C��쪛���܈���y��Sdn�K̬����YK��r�z�l-�l�A�*�eQ{���*��b��Yx��4rtF����]{��N���漊�$��Wָ���D"�sn+	�cP��j3YZ��V3�p����snkj���j.sdݬΠ`�͔�}�P�J�\��}/'\����{M�:��NƋ�#��>�Nv���c>k�Q��љ�W���zs�r9���v����t./]NU{{����LK/s3l���/���K����b��G2c��)�W����>�3���e	ֈ޴F$r��T
iEy8�W�a,]�5�&]/#J�1<�j��^o���gJ���a�iU����#3�Oa3�S��Ҩ��q��}�CW�k������1�K4�)%�<Gp�VS�f�}���.u�E�22��S;C+1s���Nӗݼ�*�
J\��r��#�3ַR��f��("�T�bq.nj�w"x!�v}g3��<]��2cX�W�<��zêo"��A204�c2uX�3F�a�{�­��L�b��#w���r��Sf/y�{]&w�,֦���α��o�sM��/���Z��y�R箽��e	��Hش6���R����f!,gvA�Q�O�'�*��>�t���1�
�3�v�������HY����	=��ʷ�8��Fq�sq�#{�RuXN^�%H7�2ۃ֨v�V;Ĳ�[�t:�Ȉ7���\��r��=�/�]Q}����g5((�=�5���"�3�Y�$Ҽ�a���"7�L�x��N<W��t9'k��*�ٞMn�T3q���]$
N4�tU�/�X�l�1$��`�́R��w���2"$�q�Lɯ8ӑ^�SI7��n�)\����>Uw�<YDc��ñŋ���:��bO�k�����nU�,���S$t5ټ����[}W�k9���t��������>�k�ީČWbWH=���um���&��x�,��1ݲ_�=��x����⯍������NB��D�����.x�Q딱�]R�oq��,H��5��Ut���p�9A>�Y�*�o/Y�n��ĤZ�
�Պ9�w�Or��W�`�9"�ܮ/-*�\ǘ�bD�����)���3��{����
�[��xʅK^��h�]{[��J�[ʬ�n�i���������&Z0槷�����i8B���ga�	<G]����Ъ��yiE���w燢�!�d�N����X�
��&Zsy!�J�F谜d��OM���=������Ǖ��$}�W�>Ĕ͞��� ��XtÌ���<���E���)8���V����'v��;@�-�o VJɟ^ڒm�G������z~��}��5g�L�l�k	��I�>By�;CL�`tyd퓉8���$Rm0�̇:�M3���8�ֲsy!����`V��z���^����E���e�J�����+rKk8��v��`�Tl��vf�2���J�/c�'
{�;��2{�xT��';�Ɂ���@�Z��7�+L�]|�E�O{yW�ʲ�J��(!���fun��\n�t[�;	'���v�ըN�)6���@8ɞu�l��哌��/�i��,�~`$�N3�	��,7�$�7݇v�����"WՅ�Z﫥]m0c�(�0$��tP�02}I�>d�gz�<CL�r�γ$ڲN���&�d��t(�L�g������p�xK���3�;溼�M0�d>a�x�v}���3t�I�$�^�Ri$�C�2q�C�O��$�'\�m�:��{�L���i_`N±�^oS[6�0l�Zp���!�����I��	�!���RN3u��N�O��Hv��<C8�X�q'�o�z��yխf��v�y�o0�O�������8���N0�8�o$>`m��O!8�����<d:�3l��Qg�����O�CS,�&�>E��bh�[�߹��������Z�����$� hι�7l��0Ӵ����i:x����>���!6��hgl�ͽy�I����6�7�]=���fs�9���Z�b�9l�O>E�A�8ɮ�֤�2tf�O�M����:N0<Cl'L�=<�,&��o�Л�&�xɌۮ���>η�y���s���k��	<B��`��6�����,����d��=@��]{�B|����ēi�RN���&��hT<"<<���}��R�y���Z�v�hi�w����bBq
���0Qd�C�Y7l'yM�x����4���'�u���M�ެ�L�<�-B�b�����%1}��x�﷨��I����:d�@��y$�fn�m�����d�I����f]�x��1�lRiyd��<�����z�?��^mq�3��)���`|�0hM��@\̡t�C��&=����!g&�!���-���n�[c�Sɳ`��9n�j�`Lԟ"�vGiݒ1�r���?���b���B�-9�z'lgZ���j]���5q�o�=�{��Y�'IѮ�l��Y�����I��2d�R�C�<d�Y�5�!�
����m���,�0�k��6��J�p�Y��v�߼c���)������]X6��jr�z�f����6���'H�<��Hv�m�7Hq��6�q�G�޻ֵ��z��������I^�N�3 >I��2J�5�����tÉ:Cl;<�1����H�q=�xE�bxn�`wl���
��Lj	��<湗��=���ýҰ�2p�M>!8�e�靲k�`k�jN����2q�I����M2m��H��}�2LCTn3�+��ql�y����	��;tï����gצ����v��+	���w�l��;�'��Jɵ@�I8��}}u���G>z�{����=���r�x�ya�RM!�{�A�O��I�i4��� V�^QBm�<g�:d��l8ɮY�I�e�h�����]ՠ�o���Я�� ����|��L݄�����7Մ�{��<}Bw�p� �k��;d�|E	��T=a�N��1	���A��MY�R>7����q�}�P�=㓩>d�:��`m��o�q5�2z�a=a�9�����;����$�Ęɤh�Vv�s�u�|���c~γ���=}ח��;g��C�d�Y'�<�xN2O�6ɻ`zy��0��<:�06���o��z�О���$�1��W�by�t������[�E��NҌ��!X��a̤<I�&��	���$ݲO��q�lN�m!�'|�B}��Y�i0�\�\ޞ���fu�TW�c����Yr*�+gz7��v�ul��ӸUdK@�N��K���JZ��B�}�a"7b�e��i,�HŖe0`X�j�@�L��{H��N雈2K�ǣi��`���}��7�7�*�Gԧ�c�������޳��U;�Ԙ���	����m�|�E��P�l�'��T�e���.I=@����3G��I��G�@=N����<���u�s�w� )'��q	�N�̓�<I�m���OP�<�hm�OB{l�'���E������H<�
����י��>q�;�]kmc��@v���ͲN���ϰ��u�8��1���O�tɌ�8����0Qd�f�b�ԓv��'�Ƞ|���1v;7#�_M���s�{�nX��<�a+��3�e��O������I����L�!��d1��0��&Ь�7�*,&�k�Y=��_���}��{w�Գ��=�{#���y@�q�i��Bm���,�	�4wd>g�:gZ�N�m5��6ͲNs�d����C�=��T�e��m���j���|�Z����;I����O���%v��Y6�f����^�O��aĚg��$�
���8�m:�d8��R�܏1U[,/�oC�)T�}�0<�ީ�>vC�
���z�OXO��$��55a�$��]�O�d�&3i<��
bC���0�%O�8�㭝}׽��8{����H�O_r$�	��T�2�xsxC��5$�&�����I�КgL�/��%f�d�>a5�y ���>���T�h���)�S�G���t�������a;f��d��d:9�
��&0��
��v}zJ�m�ԝ��'�P�C��� v�}:��޺y�����o*�9_{�q���{�Dzty@�&�8�_`C�ϼ��VI�u��8���;`v��L<�����!��;ghM�gƺߗ��:�V��ﯜ��T�|�c�NFU�뻽���~�������%��;��_Z��]�%*9�#v:7{[xaX4h�����.K�x�RG�6]�X4#�t㙑s�w�r�Gǁ2_jGrt��۸Ko��F�~{ ���� �k�� ͙6���jw@�&�9i���&�����~Xq�I�!����Rv�9>�ǽ��U3������W�LD����M3�c!�d��ܟ0���d�E$�~`m�ć^Xz��M�oV�'ܳ׉'�7ϰ6���C<�<�]��}�O���e�l�9��N�'�h�i��4e��i��8��Pdɭ��<I�,�E����2r�zÌ����@�p��;]���w��]��0�0��p��C�]�O�,����;��m��5�!�O�aє��8ɮ���5�'-�z�wd���`y�7ߒ"['��s4�1����(P�=�!�y����'S��8��n��|���`��I�u���I���<I�Xte!�M�u��'������Z��u�9�����߷�����M��x��w���;v�&���o��[!�%f��~�P���u��>a6���'��+�>P<�{����r�Q9���͡$���<`s��'��v�m<5d�'O03�y;� ,&{���'l�{�I�:d�6�>� (w�d�!�'�9�ٖ|�X��*�ܫ?�z�Dp���=���d��iya��	�n�3��ͲM����~�v�:�}�l٤��I�:d�Y��~����}������M$�s�(��'��f_P;d��:��`q'OW9�M�:;d6����FY�	��X��{�vI�T��ߤf�m���Wu�w��l�{���Ę�:��q
ɭ��$�O�Rx��8§������N��'̆�Y�!�N�#�x��o��U��fD����1S��%��Z3���|E(�l�N���;�M��E:�HO̳��UzZ�h]�D�e4����ʙ3�1��y�v��}Q�����(&:wc��g%)��3M�Nl`�!*���ි���_���s6���MjJw-�3W&�=ԗ꿾���.�j��8Ͱ�'sy�L�"���'v�f� V#l���t��o��ԕ�&�V@YL�|�y�߯6��VB\>幖l��Q�{c�����z�d<��j�>N]�q��X�
��&Zݐ�%a��a8��"<*Ǉ�Uxz���q������o>��z�+8{�'H��L=d�8��퀦08��H��v{���h�xd�Нs���Y2��݁�����8��~�}�o3o�h�{_x�x8L��f�5��N�h�xN���t�2q��vN�8���I�M�y��VI�u7�8����7d:a�bg��sY��׿sܹ��@�
Ó��P�`h�x���e ��ά�$�}�$�8���&2|�'h$�N3�'HN}�x;�{�<��c��WWbЬ�X?k��ڼ������	��X����$:}�QBq��Rv�:f�ިOL^��� u-�j�0�XN2mN������d3����n�ϫ��YO��=�!���>�!���C�{��'���I�$�S܊M$�0��j�x��4u�I�MN��m�]��y�����=�]k���7l���NZt}�H|��:>�O^$���9�<d9��$�1���$��:�X���5�!�N2u���}�U*>P�e�Bh���Y�e��zt��<�Rr�'�l�$ݰ3���&ө��!��ѿz����<����9�d��_k�d�'S,Y<gi�ޮ�ϵw�y�o���Ov��,*CĞ����u���d�=yd�ݤ:�P�i:x��̒}���!6ɻ@�;d��:�{� LxCΙ���~ɂ~3[;���K�Ď��b�̺"!OiC͆�%��6n�(�_�ϲ��[�~wS�*���L=λ�*��.'�����k[��"����v��=���e��qzn���Ѵn�a��gX4�w!�~�������n�C��R��P�=I�&�a���>d��5�'̗�O�M��:�>a�q��a:g������Z� td��:��Wz�|z_Q�W�|�{���;���1�<���Vw�
,�hh��&�dl��N�ԟ04u�	��9���I��T������l
�y�f�_ʗ-c����a9�j$� w:�$�2bNoq����`��6��E��a0�mğ5'R� q�OXO��y���� e��Z'u��ϗq�O�q�s�d� �=C�$��������}}��N�1u��Rd�u�,��0�Om$�.�>a�̘ɶ�4�9Ҿ��6v>W��R2v��{�#�p�������'F�'�Vh�p6��N�s!�N�!���I�&"΍oq%I�v9d�a��,�0�|�s{��W�uoz����}��ι�:Iɫ'�%f�	�C���M05Հ��&ӏ'�Vy����,��a�N�`k���-��7�8�P���=ל������^k_��l�>(=���0��}a�IY��O��S���6ð�P�N&�E��߻��,�i�o08�ݲW��nq�(/����J���� 8���RÇ��XM�h��M>!8�e�靲m��s\�4Ͱ�}��铌�	���~�E{�㷜���uz��}��̂4�����K������ox�Tq�2P9yy��7K���6�`c-��4��Wf���ϳ	�t[Ͼ��_�(~�=u��)�%~WR��vu�[�
��+.��ujǓ�=7��7���v���ut&��s�<�F9��Vg:&V���+�a
��R�q���=ur�'tl�Ʀ}�x{z5�>e������W-�l�ru^��ߞ0�ζp72Ù:	���M��WTͧ���\-�3�ZT1h��kf$����tf�as��u
���f�X�3��)��*�;����JK�/��{Ív�����a�]_�K���	9�0��]ۮ��'�|����N�
�!e^n�:�:�r�ٔ�v�.	������u�S�飝�Ôo����)�&��w\6��MZ���s�b��3�z��w7�J2�9��/��qǷܹ��:�hmѽ���r�@�+�m�-ehp�c�9
c>FE���p�My]Ǯ�.r1��0��.�豖�v���{�ue���L�C�:5T��{F��o2��:��Z<ǒ I ��eqB������we��;ӇP��� �u;���[�$���m܃9W��'k�7;�Es�E�1�;pV�����ut?odzh��պG%�b{��=���Ô���s�j�n�n�%<+�NB�E����m`�4���h�\w�T֩g�Q������?oP���tnloR]�1R�g.�+A]Br8���͑�X���v��*4�=ɨ;�K�}�46of
(n�g*�C��c�e<���g��l��wii5��	6�$����d�p�;���k��XNvA �EJH�\h���;��	E�
��bh��
��Q?i�)���5I	*)�W�:B�v�ΫbT͋��D1���	&ssZ�3���w�M�cfD%�8VU+#2�2�t��Eh5�����cX�fYH���d�aޕ�m�	��%F�9x��\pa�v�f�F�S]����TX�.QAe�.�H�зb(Ѭtk��ۢ�P7|�F�5�yts*D`*
��ؔhif�tlNU-֔j�^�w�t�N�J�Bъ�&�7c��" P���v���ޛ��`�׭���:�b_e8*�m���i4q��]�)ujJ��,� Yt�sט��������ԓ�Ct���S�
���d��bb}���P:q��ZԻ�c�;X��CD�g	��[z��o�������Q�v�[� �k����=MS��V����w�*����'un-�ŕ�ӷՒn�uF���h��໤5G�+��نB�"sg�};Q�������
����tv�F<���A �Q�U��Q�PhUE��QcQ��.�
�K�ĭQR)�*,PR*�J�TQb[[J�b�3�Tm1�aX���j�*iUDĒ�֫�t�%��J�֩�q��R��6�L�QEET��[Z[e�Z�#"�Vb9�1q��+lh�VJ�-2�2�����YQ�˘Wk.6
��B�
�KAul�W5U��j�)]2��֖�1H��-J��QF�:���	D�m��j�1`��TY����殁DQ���UQr�X��	�b��"�5���YZ�
15h�[1TX�R�iT�����(,b �K�DZ���YmXbV�f`�Q�,ť��cQ"�J�����JU�UE"�A�b�TTF�%aU�b��b�H�%B"c]9�A@Pm�l�%�b���--.�r�%
�X(���r��?ٕڈ��f"�y�{�tՙ�/�eŷ�[�k}ir�/#}Ρ�ŕ$����5���I��Y��� z������������S�jG�k��c����c�9Ō�g{2�������&j�ߋ�W���J
/^��ڽz�x#s6b`��=����z����$ֻ�Txm��QY��+����S�\�*�/N�)=���]�۷S�ս[�s���j���	�������]�	]ѻn^I�ئ��#D�bT��lv�n;y9uކ�bv�u]�1n<��ϗW+~AZu˩Ы�׷;6dc9�2ȵ�J;�&�̞��n��^�*���xyˊ��Hl�΃3�:h�'[I�p�t�j��܎��J��ų �(��=ꛊTb§ͺ-�	�'3L�L&E����jgR!�pX�H���f�g�j$�^�֓��!�	�q�N:�Ϫ�����M�`�k4%�$�������L'Y��*�]��)�>��l��ّ�ˡ6`�Jݗ��A[/��oH�fr��ڇ����_�7e�Ҥ���-DvZ[h�s��bܰ��S3�[Y֮}��H��:��i������}_i=�F[��7����0k�!h����spo����4<B�={=:5��"̥�rϟE�W�q@,��v�oD�G�\Ճ}��.-�	m�wF<*9c(W�9�Ī�����Y^���,��D;]�C�f����/^�kc+���x� r�ݮ̈́�)��V�'�d�;�e�-bt��U�&�_^]*�FZp}���˟wfD��[r��yڸ�`2V���WT[��u���R<Ϲ����s�)zU��jhĄ�!&�)�3�Hahn�����vT�	48���I����q���dblNW']&���Y�Ȝ��7����<Z�ٝ���)հ�M)�jFH���޾�ynf9�A��=fg�Q�|��';��� �)p�}#B�z�GM�*�p6f
3x�������y+U��8�5*]vq�T�VhC2��Z�Ԙ"nk74d��Z��*�ZV�ѫ�r��r4�2	�_F��˟L�����O�66�s.��u�����r��z��Q��M��U}��;u7��s3�Z�b<���8r��]�'};��'�.>�@uwL���R�Ln8a�GKSY	^�����H�.�_���aQ�x�a�+��Q
tn�Vm��&�fzz��ue7������i�ם�s���
J(!<�Eˍ�]���"�]Ԍ�
��|�1����v�kOaՂ��"��J�X�Nê
jfR�wB����ҩ���
x�JC5~�vI�L'r4W*¦�oyq�1O2&���nƉB�9S���&)����^NE�V�����-�M��'��4u�,�2��m��[��������j�vz�6!1�:�%Ȍ*������e��uA��d7w���e�Wsj�jʹ�n���09�¯Օ@�@�m�����g��S��M���z:ڰନu��o�.zq�7���vE޷����8��U����g>�}A&U�ʮ|�O!�n`�}#OW-o�woZ��`YKTxv�jdwp�Z���n!8���HH;�Z�kgg\��_{�{�o�;�{6�de�����d,ܒ�F��Fcw�ʯM� ��f�jP��Ѣ�̕��޽�<��׶�;�*��Ӕ��Wg!Lm�o�׵������Q�.EV7n_m��`J�Ҟ��|�/IOҫ�'�����XJ��>ռ�;��6�w�&�76�������0H�|�P.����3ǵJR�����s��r��to��ʳ��|���w��W�����F<�V���ݮ8ƈ�j���-����!+:����%��j�8�:k��;��sH�YL�>����:CA=gF,�Vy�,�~���-2��Ԟ/�d�ȡ/���ӹ�pbQ\5�Ȝ�fK��"˸`ƺQ"�h1�CX��	������� h��7joN�6�x0sB�+�[G�KN��f�#��\��=�}���Sg�i��+����J�gn�����aH�o��~��W�s�"���Ժ;���v�kH�v	��[���NPŔ�e���,� ��N)�D�n,���{��9�[*?	�2܍�W�k.]y:�[�k�tK��J������fLW����D�EM:\e��ܤ.æ%+Α��*�h=#���삔e�}<b}��)[���M͘�ůˇk���K�5����.{���I��ge�#�	nk
ۥ2���̜6v���/5�n+�]jG-k�[���G���E1���z����+*����N0g%�=oޚ����p�/d�����^s��ylDΥ﷽5w^'�ǌ���~���pL�}.�ٜL=�%��F�Gǅ�'�u�����x3;
�z�^�g�+���\�=
�dSAt�Z%M:�==���T�i�)᧖��ӵ�1��_ �8k�!ŇjWu/���\轙�S7
=0��fl|˗�v�C}im_[n����Bt��<q{��O�=}��I��HĪ=\I�I,Q�۹�6�M>�V���wPI��mK�����֐�m�B�ל�ұ(R�����9*Y1|�ԅ�6��8jY�ܳ�_�� T��I=9�7����	�V��
�R��<������G�]v��[|�~��fG�&>Tt�f�;�oZ8�ʰU@�҄P��q�af�+V����g��CT�B�	ajX�8r�[.o7��r�0J�*��B�G��q�AhKp@��{���u����RqHL�E_9z_Pn�w��X&��\��/��6��D�W1%;���(4��t:���㖶�s<���G��a�gz�Y�K�φ�&�'�|�d��$q���*빩����u�=��w@�de�-��;�5'�j���k*+��׻���1f��[kN�u��os�;Q+��zG1�
QG�9F�z���4t��"=WTz@��W��������̳x����
��e����S��f1�#b0LgW�dY���dn��;Q�5M��U�\��#7tgI��&��oo[��V�%l�^i@ĩr�\�$����	nf�|3��+����Rk�!����ܭ߿@{�7�9s�韌X�W=���j�]���
ڜ��QU��jzϥ�w�|��%=֥b�L=��/�C1���`N��A����3n��Y�^��[_;vT�#���]��-�#g�!�ܻHT�Q�tf��I�x��<|�H�z�i��B���*M�A_uNz.k�	{�N����O��-�q���U�Eqda��A�WVFS�.zhjtDe]m�h�����	�΃�Ǖ[Yɔ�8ʸ{wnWLfSM��{�Sj��T��f?K={G2�T/����^��V�}���/����]ʮS�RP�+2&\mWa"UX�ZW��g1cFѾ�^iY:��Ua':�HBUp<��;����Ȅ&n��N���m#bU67�A2851M8� Ӻ�fb��1mlt�;��1l�M.0��x�<5�jl��Z��w"	 ���!m�}�e#"��6S�3	<-X��9�����t��9w7z� Lr�t�|�;F��S������О��R/��7uuǕRt��	Q�2�s9��W�{�=`�U���\<�l�5�,���<'/9.r]䈳��z/�R��B/��&'��}1ʬ@�1]�-�[щ���b�dD?f��c�M]Q�]3���=��=t�Ҧ��9[N�چ;��#8á׈ˑ�Y�n�xP�l�i��[ ݤR]n3//�׉,5�j��ׅNN�^���i��Sݷ;��R6m�9¢�����{�k�i{Ʊe�(���O�� �pbo�}�Y��׼�r���&���[��6q�:�l��g0X� ��F��Dr�Ucwp����ԳSO��q�;(+�w&dX�����]qڌH��o��:/4�ijm�t�����"7�9���Df�q^���jޮ����g�-�}MN'�<�%����#z��e�Ĭ�їj&+8E+�cy���]Ϭ��il&i����5�('��'b��m�^���M�&��+�b�����å*��[�����TU�g}�<< s���}%#�~Op���
�%�~X؟J΀��V�1�7���]wJN���⏚G*�fD��:C`iV����v�v�\ܵO����2�0N�y����ȪN��n�&�����^�|-P��R����e*�{<�	�Xon�t8ط7�v�����:]���,a��g*T �nS���K��lw]��&�?F��%71�q�}�������#�oD)d�s��9�jw����4�#��$i�"J�;X�Z:���f�-�j�V'Ӣ�1�n�Y���k2���.���2��E<��ҧx�F�M0#��A��������w��b��i�}�ۼ�vм�JnX;�!^�N3R��.��z�8mW��Bi=�{ԤK�[+�%��D��=�~ܻ[W/�|�wl��
VF��Q;��[�α&��+�-b\����OH�Ӄ��f��r�h�\g�
�eұ�W-V�c���9�v�#��7en.z��Ǚm��s�W[
_xx{� �_Mê�S�7C���j�گBJ}a(�^;\R��ehƮݷ/��v��=���I���H۠&xW��P��;q���+.��0�K���m�X��.�)�V��[�\dh��B�o�5K*�l�o���Z#��1��Q�*琍��
����c������!�/��}�N^������k��{�0FJ\g�9q^��X��_.#�﷝u��.2�~;����TE���ϧs�!Y%ϗ�+���f�ѱ>��2���H�Q�c9"�僂�&�:��u����ײT����οfv5�k��g�i	���׏;-1�f ڜ�I���'��W�Ӑ�WD�U���<.V�K_Zk�;=�0Bc�D�0�g<�\�N3�!��Z$�?@�[�'��>� �u�۽[;�J�a�e�2��y��a.�8j��9)hw���j9�QȖ�ޜO�Wk�-U��:�,�Â��+����7���2&%t8�:��<��`�&�=D>��^az\�et��e����[�:�{���p�j��+�x���ךݪ�7�RT�������k����J�{�^/�+��'���1�7]�r�̗��X�<4��u�*���Λ�iJ�wu��,���T�Ű;�vġ�$��Z.����.|]ˡW��ݱ�d3��MM$V�gr�������?A9C�m�e3�5+��IL�%`2��
��,����r�ltoE�s���j��B�5���BҺjQ��uj��}�Kp�κδ�c7���]�@,��<��Ig��3��)�4/,*�q�r�쎘�u3*L��ε�@	�D��n�P��n�G-S�Þ%D�.�#.���}+S*�^M�[R��q�YV��\C4�Z݁e������'nҭ5ɴv�\U�m��e*�:7���\�ݾ�	q��żj$�gJ-P��}c��;nu�k	Dq�θC�<D�:F���DT�"�wJ���f���҆�l��9�
�8u깓�-�kD�}(Âq}�j�K��1Mxk�$9b�>�ڌ.qtF��)���{�x��=��?�8��Ǟ��s�y�v�<��D��1�.B��~-V4��wr/���>-�HV�cC�wp��x�;�K_5Ƌ�;��P� �� lȵ<�M6�h��K �˗n�̩�7y���s�ߨo}�	rV��a��Aza�7h�nP(] =�엯���Q�����T�`�h%��C��#��I���Tt� n��w��Tj�.��#�BTӺ��+��D�c&O�T�:v��;Z.���V�ˊjʘʲR�i8PU�C�$\(0]6�;������N�c
CN�jqK��:1�fo%��mŇKY�fdI�w
2���㗨@	�2���*w�f-�seZ�5�z��^n��`�.��{�<퇵���#QvdX(�q�s�h�yY���`�)�R�l�"uz���y��|6VU깏1��z��ɳ)�ubc��D��׫��u'f�+�n�J��O�q���j�9���bܬS��"�:�u�I�4,gt^#�J�}�G�����Jn�L}G�����=o�ռ�{w�C%0��+��x���]��0�ųr�u���J��l���k�ٛ�v�]QN� �j��98EV�����.�-X�{J##"�h(�q�[J�E�"�X-KTKljGUb�"����TS�ɉfKEUX�F�+ް�"ʍ,5lG)U�I��Q%DYmV,�a���VR�J4AEU�bb�c�%X�!Pr֡\d�V�9[h�W)���U�X�����9�S2�X��1
�%f��J陃d.�cA��9J,]Y(�ЖB*j���@M�h���LPR�V�5��R��V�����4�ʪ,1�h�RUV��4�!�5�mr�D�8�VTm��f�M1�e�J�q��F[����)�P�

$��+++�lq����6���*0Y����aCdU*(PYY�麥�U�]f.+i�q�fY,EbȈ)i`�R���
5FU�`QX�akS̥H��C�4�Xi��eJł�J5��S*�^\<�b�y�fcYS�!SO=Bv��Ƃƚ��sn�1����Twώ����T���Q��]��V��x�h����k+~��p鲞z��&&��=�w8DO�Uq*�iGj�?	*����ˤ[`��uV{�̭�&�D���K4�2!�wv�Nm���P�hy�ŗ=����O �UA�u��k˗vRþ���E]���l殺��E }�n��ۇ�=������������i-�Y�.Ў��OJ\��6�CW���v�{��r�btNW�ѭn�)"�q�k�:��q����eq|��&�)�z]��<�Z@��q�1X,�qi%��] Uq��B���ɾ5K�C�r���A��@��So��tʸ��bc��U��T��:n��8�]�W*Z"��$���Q'xp�����b�Ώ*KW�9R�,����W��v���t�� 9����(G��[f�w�.�O�Ư���G*�oS�k��U���G�2���b���I"�w��q�ѵ#N��&�����������'t&����[�5���!�o�5���e]�W 9��]�v��:��/N:;yz�>��vVo��%�KR��o��^w��YT�29���8tH����Ѵv&D�6�)XJ���b�N�k��;�����q^�v����iX��K�~��h�sr~�T�E	��rF4�e8�%p�XWf�M�B����[�;wH~}>a�6%S�(AP����(6�U�����2����Q/����EeSz!��S����v����}/�R50��De¿n8�|��8�X�ux�<Ttp������Ց�o+8��"�WrC؉��Ų�aVn�>ͮ��l)�8�k�^��,���<w��������u�WYU��+�������77׻��;8խ��y�y:�����=���K����r{���]f��Q|-8�x����k��}^3�k���%�~�.��H�'�� �M�n���}���R�$�n&1 �B��%��pT�-_ �9D�$�i�F�_�ɔ����֜���Q�ʂ5:���ν��R�����������v��	�N~Ju��h��F��irR_8�Ň���~z��U�I�v�{���U���_R��g�ċ�iB4N�[����O�<�,;�uv}t�U��n+.x�T3�!��z�7�BV���C�\�z���ʾ���!��7��w8�-�.NNn>(�Y���'��Ⱦx@���Wiſ%�6&VtP���@]�,��ڈ�j�r�.yY��@�(�rr���J�P(�1V1nw;:m+�0��N�L�
h�2idP�I�#O$ku��� �3�Uݠ��*2Em(lK��N�U8���pʯ���)���j�.��zx�G��X�����)ˑW��+1φd;[��L������4o�%0б�D�EM:W����WXJo��+�3>��j�����p�cw�Q�@������gU��NY�;���5y�7�O���=q�Ѝ��W\&厇r��ƺ����0'�T$;c�k��y��N�ޝؓ�x�VDn�޴(��T�V��<�7/�Z�kz�$D���k�o��h��]ͷ��@�r�Rhʝݺ�ͺ*Q���/���[{j4����˫}XV��gV�E�r�5Wpy���.��Ɔ'��sF�³��1�)97P�өŝNk�&���3������2Z{ع�M���Y�݊Uk�7��쒍�D�5u�xn��J+5�V�d���:΅;�hQ�(�a��a�.�fHWS<#!�y�U(b{��ى�Y���iv��yZ��F'yB�
�����,6��;�ZU���P�+dbھ���+���l�
�U�3�%{���{�w�7�+�\����[���ϲ���)i�n\F���+�.{y�uR��c��v8>��倽��9BNsy��Օ�rb5��Exg��Ζݗ��[4�/f]�&�J��no<ԧ���Ԕ���w9�ʬ.�1�m�XC++��f��[]-Ov�i��v�B�{�r�*�Iz�#ʴ�I�S4[�S�p�)E3Z���;�6��ڸ�	j᝷����MӴ�d�8�~�)w�6&Vq��2���Vz�;ʈG����^[\�٬wU�\�A�!>Bz�\uS�B�_X�|И����k�>�Ģ��c;b�[0���ɉN0!3�Mfǎ���]���׹��eĄ徇ɸ��.��V\�4�C�;�z[���ۓԖ6�Θ��뙖�@pr515�O ��ɠ� a|:�P�::��پƥ���Y׮M��)��Hy��
:٣]<���]���O���X�#�M?T%�8��kӯ^40�:�FF������t���m>�y~Kv��{�C��j��2%���[W/��M�0{9_��wܸ���{q��*�Ӕ�ġf��\�������+6x[�3[Џ.�y��׉�22�u���p�\�:�/.��̌�W%���e�ُ݊Wme3�Bq|",�[�9O���f��':o�ټ3tq��eI�T�s�:�6	u{ҕ��ϥ_A�ݺg0&A������K�K�T8�*�����;vڇ�������W2�L��IḴr�]�x{�{�j���&���E>��� �|���:��l�q�YRk�C�t��5�D�b�"S�\D���x��/�[���p��Y���ǚ��#�q����B���G�C�;2o�u���	R]���iw���#��W��u{G	���΀<�-Xp�9��SF��y�W���*����1�xdH���s&%�q���_f�ř��fmM�.�ҫ�w!�[�ĵJ�v�Eg��<.p��~z.�DZ*q���mߡՆ���p�-Ʀ��o8;�9
EI�AWbU��18��j.cbN�0N>Y}����P�l���M�ފzl���(P��SG�|}Y(���m�I�պ,���<��QM{�����x2��](舃:�Իogn3m
����p��T�e�y��c�%i	l�կ��"�Y5�8;K����%�3-�����Cq+jSz�8'����n��ee�V+3���В�=�xx'Z\��C���F}�ƈR�F���
��D	s�YM��ok�g�g�pcǚ烵X�5�ۦ����*rS�{x�)$��Ԩ鳬l�F���*/��簮�hq���R�}�/9��)-y���6��*ӊ7���N5���|��̊3�8�S��i�M�����N�6�S�#��Q�X���3F����k�o��'{�^��0؞�N���ˣ�ݢ3��A��Ҟ9�6ۅw�ҲU��Pl*���B7�\e�7|"�G�w��8���x��)[9�	-�`t�V/*o���#b�\�)BZ}��2
�里���r���=޼^�g��sM�w�żO��z�u���x�J�G#��.i�)�RQ#.���ґ����,ɓ�EG�{�
>�$S3�]�/Jы{*.�A�m�2��$&���jo���[7�m�G��H�Yk��1b��l��<X~��_p�[�>�iG��)��J"�ؚ�ې��-J�}� �&m4�X�?;�����=]p���:�n�,�kn�)�%^�w�&�z�V�ƽ��G�[�2���h�o��0��K�e���;�B�2�v���̒#�u!t&����/�]WQU�!�Ĭ*;Ή�R�Oh:X�L�cmƕ���V�4�Z�5b�G����+���H�>�j�Ġ���Ѫ]���v�n%|kn�({8e���k5
\���0��A
���6�3�՞ս��ռ�D�ኜl^]��Ȗ&��@cd]�͋Z��Jn	���YyY��q��kw��P��T+���o<��x�=Xk��,y�f�u�|�)���E"
�늞Nlp��X�g��0R��&ߖS˪*��K��1�yg��E]�����%oeF��eI�pX������N�1�׊.:5J�<��Kw2��=��v�{6�w?,���=���X��9O�gʖ���_����`��/dm�	�Ӯ�3��h2����Y���-�5�X��.�����Mv���K]�Vs��r��`�m!j�
n�/k�ƲMC��vx��]�X�FX�^�U�S���9T�����.1��1�R��3�v��x{޲S䓼���g���q�}A@�Y��U=��;@�!��ң�����/-p	p���{�>|�5��7��-��ت}u�v����iR�=�D�Q�����ͽ,�*,L���y��T:�,g�`�9*�P����¸1��`�#uƵ��+��F/mV!���޶
�=�{�(@8��w���O���4�@�ӣ���=gf��Q�#z>�?z�ќxxo���$t��~��U*����]b871��䭛ˍ���|���<YwV��B�W��q�X���*o�h�Ŵ�5�ӗDʊ)@iއcei#`[K�S���g:�1p���wBP�������)5�VO���ގ\'�N��;VTL?j�%E���HND���+��C�3qS�����N9�דw��q�t�zj^��ZT�>֟��5�� �50E��̵3�P#�ʄeLF��}���"�%��%R�@�~^��P�ɸp�Pkj�Wt�	�)[���W�����2�h��a>���ĚXo�ǔ���gN牜v���`Yn�&kSjv��.�c����k!�d��icw X��7������:\iܚ=�'�S_غ����,o�[\��l������Yϓ/iٜ�>KN��J�4C��!�5��e[=�������e�����`\G�=��?K�Ne�S�hز��5\��I�6z6��W�h���.\ Y< ,�]�-rFͣң�v�+��~T9�E���{WG#��b�� �����be���f7�q�y�ؙݥF��m!nyD��4�B��(��i�!��n��D:���0wi>g3��_W&w,]�G�z�'�c��AugG��Ǉ_	�j�g��˩u�r�Wqn�4C��u��W�T�8:��ps���ˉuV�1�Ui�}*���v	�$������o�m����|J�X+�*]@��-\}9�yN>G��X��k������itq5��Ed��R4"��u��t(��~QK|f��x�] 	�I����"Tcm"�L�n(O���/�P�[D
#F` h���o��:�;��Iے6�pr^��*	�*E���):ȡ���O��pP���z�z�M]��C�#W)}.렧`��0UdWo�z�j�j=H�������S�=��.�6Vr��o)�JF�j����.j��:=x��e��\�Y�PqR�l��r.�a�f�u�0L(�飜��{�x��dg�n���C7/�� %=��a��-��{�\�2��P�����Q�}�]%�x�+��.��'[�U`� 1�<L�DS��i��8��"e��ԍ5���(WK���`�$�k�RJ|H�T���3�Q�ep��*�p��6�Ź@����X6�f�j���KC���E�����܀�g:WU�'#+�b
P}ctsWn+Z�6�nGKX�M4!Kᴱ\�o3w���p�V���-�Gq������u,���x��V�-��ܣ�Ue���d�w�ʽ&ӹC�9�qc�-��ekys(���}���!0�N.S�#��5^����&g>�3+>u�c���]�岱*��9|� �7�,o{��5�'_JY[˧v��OE��N��H��;۔�8n�rU֒�n�.=��*����9���t�c���@� ^;����Z͹ճ�LGq���݊���ǀ$�v�����v̰3��u0s�v+�h��.�˧>f��>l�j#x�Īv@�&�s�4ֺ�7+n3�
�=]K��M��H�N����1�L�QoN���@_X���t�1��7��d��pM�鱺ة�8���G��s�'S�y�}D��u���]�+ɷ�;Y�0��V��Z�9��Ǚ�#I��'��%�dڠ2���p�N�혦f�0Y��(}\H�)�XGb�+�ӳPGq��v��k�+.��r��S��gfA�l�ȼ}�8�oN�iWѣ4v��8:��K�0����+�錵��˔���4�,�C3gj��k��>q���J$�ZL�f6ۭ����y]�j��:˸���M��^Lz�V�2�*ة�H�77
�hV�o�f1!G*Ŗ&u�{j��hS�>�����܍���]�WM��K�^���&	7� ./�%r�:�o�
m�Pf�sx>]݈X���g]>c7��D��I��n.[y��eEg[�S�9�);��wt�}4��1d���$�Y$�]L�X�*��,U����f�0��.nHG�ueC1�+"#ԹWt��R�4���;Fh�"˭޵ׯ���͖f���4lYM K���4�;�q%K��cjjT���<�x����L�{ǧ0��ջk��)V֥j���	br�KN�]��hó�s!�}V¨�n�����{گ�P�� (
�"�j[�+��6�VV����b��kU�%�,�U�j�VQb�ks(.5GV�VТ�hҢ:kcp"�ڬP�`("%J0Em�R+h[h"2��̃��$�Z��n\H�
c(�B�*T
ʬV3-ƬUcX�e�mգ�TYYPR�Ak(�R(TP��Qm%)IR
6Ɣˌӧ31�V���*�h�����n(4̮%��5�q0��lD�-���)J2��h�Z�[**��*-�X�i3#m[)Am�-����U�ee�j���R���j6�-(TV��j#��X5-�(U�i0Lek%�DB�[H4j�r�f6��F��V���Ej"��@P���eb����chQ�)F�eGZ�����BĴ��hŭeDLB�
V�ij$�	�[��Ck�n�%'h�-�'�dX��[|/���<�{�Z��Uܭ��'X�x�+�@�	��ŭ�xx{���}���;v".�T��S.dv���3����V6 �Of�\LyS�u�R]FWv�.��d>y.��H�Cmrcgր\_��/��R�>U(M��r~�wK��w���5�ve��T!��A��T&���"��nr���ٗ~� 8���$�͊ڿ|S�X6ՠ_��A[a�i��*�p�yU��$tٗ�!'m��AZ�Qa�D-��X��'�i�~�AU���l��2:yQԺ+\v�e�
�聑j_M��d��Y���GFF ňqc����}=Y�/t���v�[3Dc�1t�^Pb269�$[���{�6qw�a���������X�������o���<}C*π
���z=k}+e�u������x���G���l?(U#l蔱ptgS�����k��NH1��X=ë�)|g�Z���W�ZxX��$.u��R�P!Z��#8��N\O	�W�(u� �����%��A�{�7Q�빆�^pb�˷��Qִ(�C�,�\nw�Vg�qo�f[��������Z����O!�[y�N�om� ���xN��u;/��T���<\�RE�ds1�!��r�]O�xz^u�E����GGܨPV�h�<b>�+g�pF�ХGuB�qsC���e����R��l ��>�C6��q��q��z)�RTN��5���{ ��+2� ��y�LA'3$l��x�`��T�1m".�öVMb��.�wax���T���ޢ�5ȟ,V4��@i���͢,hᵥ�5�b���4��ú{T��|�!m�d���GIK��S��%�TX�#� �ș�T^���L�*�ox�۲-	}��$D���&B�p����.H��/�À���Q��S�<������{�.���BA��P�1p���@���u�P|$셢�#����@���eR�im��z6�f�'���GP�7�'��
�/Ψ�DpyMXؔ�ڊ��?����䲳1܍�ʠ���/�C�:�9����=�l ��ؾ��|�ܽ���y(9�%�~��+���Pv瓧���P�6#&�#��71c�AZ���ez�f� v)Jq�~^�����z|�֔��nZ�C���z��(X����r(_BC!=}|������ڐ�ҭH��7�8yF ��x�-"lKs��ַDdܰ��W�.�_xx{�'�fi�D���J+�3$����m��!�K� 8�����*#0!=�U�������}1�y��p��"0S���Jp@ʚ.�-��ͥf��N�j�ŧ۩b+�������O����X]^���J����X����8��q��vmiS/�OF�Jd�x�ӑ��⟈�3=�Bf6*hs�NzNz��5.�X�^u�vu��d(
w���{5z�D��9Qb����r�%�Zs�g5
�k;c�
����=�C�2�J��3P �[=U(�(l�L�F<I%�Ӽ�AO��h�GVAxx?�7L�0j8ϲ�p��z�Sy�x!��H�Η~�GGk�0����o~5�Դ/�������W����JS%����}X5f�eYlf��S+XP-�PE�lH�R��t���871��
�wU!���uj�����:���}\[���X��u�@�D@��$vN]=o,{�N�8����ɗ-���N�ٺ'fN�un>�9�,�L/j$�����BZ�
��״�Gxm��IM��Y�e��:�.ua޹*C��QU��wRD��YTWa�m���:Y�u퉽�2�ҨojJ��	99��}���Y����9u��C��`S�s��Ä��wB�6u���AB���-��7v*�@\�w;�2;�ɞ�k��!�.r"d`N��׷�!X��E��XE�{�o}���q�ս�tX`�:蘯g�����ĕ�0(&G���X��^
�s����:P�v�B� \�o��fɂ��x��f+���eymO&�d��K	���2��Ҷ$XKN�j�+D��)̗6ѫ�����e
鴷�����+j���*2Xrռ��PcR�%����sQu,\�7�����w�iU(@wհsiÛ
�!ߕs�o����V�B0],O��WW/B�_^��rIF�(d\p��)�����|u�F�.��A�wq��94�cY�7�m�H|�cj}Ip�N�I�X�٤�=<�Æj��Uj^�����
��k;�J�X�k�u����T�-����ˉvi�N������i�M^�����ة�̢1�A�,�Yr�NZu�P���J��#lf46���U^J�-ž���[��K�³:A�O_:v��p���2���.�k�D���[GP�������܍��F'�M�]�)��[7�������綗=���'犰p�ʕ+�����U(�%K�t\ש��t�����m��{���!�3����/$�zI�W�B(b�D�	9�I��7Ң�����q�iy�:zz��4�=�n-*q�]�i��=~���WF����)2���	�K׽ݠ5��=Ak�41�v�*�Ϲ�#'"�gb��ʉ!Њ��Ǚ��+'�`�����M���h��N�g��Ud���1���=
��󆨊��L���ѵ�p#ޤ�e��-R�@!�
���;tl./�T�ީ^;E�� s{�Y�*�~�Y����mWQ�]E��4�����������Ró\
�����?{�$�X����>���q �
�~Ճ�E���V����s��=�3�3��<=BCG�q�'üp�]�:�t�o팎��%�TK�<Env��osZ5��/�6�ѓ�]�EîҮL-u�<�cb��T���{wL]纅_
XZu"�b�ѩB3�W\a�Xﷄ�����J:������O=92>u�^�s�ת����$�{�z�Vs���7��wZ�^S���e�ot!�cB��&%��8%�3�I���v�u@�9E�}�eo燽��z��N�vd�NE|[*1#�B�N�8�J�c���x�t�O�N<QB{ӹd��;�tM:�v�xsԴ9���� ������v�<dA����g� F�����K�۷Z��n�Q�BE��p�eN��}V��P�����0�[��#�D�o��}�����P:,1�$-uή*U�Z�����Kg���ӏ�[r5�]�}ޞ�v��K��Qqx�W�i�Q��ڗ���$���3$P����͍By3��5�6��s�"�F�V看��O�#M�E1*'���b+�!�jB2���}l�{���%�<Lϑ�t����*��]��
ϧs��|�=���\9���ԡE�}�~�A  w�U��k�EZ<9&R����/wIH.b���w
U�W��r�r���[�t�K��Q�O���=��ƿ���a��v�r'���1C=:��.�a��g���J�J!g
�P@��r|]	�!lm��w>�X�rɢ�R���p�#�.`�ق�aw��fRgΥ'�/٣��=�7uJV
��j�L�yW����y�N0}������P�ON��H�x��RdS���W��夗Mq�7}׹gbP�T���I-�k�J�劤:�|V�����/���^*��ptWE��D�҄W�S�\�����琚�E�b�"�*7>)S�}�;޿cŐRt�!��*�	L�͆��*Hd	멅h5��uRǯ#�ڥ�����v3lX\WHo	/g��!���PyS�����0�l �C��n[��g��d$}�PdJC=�F�S��X����m�{Y�mo���S�{;:�h�D�ϻB�yKG�eO����{��k�:�^��*�ip�l4g�T�u'���e�f����W^:4��U����O�h�~X�B3eC��*�W�^v�SٺG�l�y�aP���z1�;n�C&E�X��6�U����O�ҫ�2S�%��,ߩ�铽N1�yj����zr/͢��,l�!����\�~�Y��s����k���F�葯�ʃ��[�B���
e����-�r�Y�Tc���רڲ
�����5�i
��`u��.���K�%�t&y�J����]�
����E@��%�]Md<�~q�˭��[�0��$�Z��͊ށ�XOV�F���l����%π�+{׼f�D��e-h��u ���\�W`�}��d�#��Dsz�kU5f1���w�+:�}� ���\�L��3�OG�'�G����x9��I�a�|+�uz���ZZ�h~� O7��gܚ�{����@UNg�v�+����S0��
\+�2P�gA2�^�]�ֻ�{������F�Nh�"Hr
��!
ّB���S�C�5�������i�Y|�J���4�ly|��ƽ�	C;�`UƄ���1�#�r�j.���sn'(�C�J�t6FIt�Q	Ո�	�EM"��A�VU��Ͻn��_AV ~J���*2:3��.o&*E�EL�9
'V/��@��=J�B��Nw��+�=Y�h�T�H5�-'���+��Z�z�S51B��DHN�9Ȗ�'r��� M����A�B���xx�vn�(�[�ɨ@���c�N���-��a���n��lS�wk{��.|�z��	Y��6�sP��Y[��(�An���bz�]r�cr��9����{B�!,W�y�� xeLO�S6��]쿧D�;ˉa�;3,�[��m�q4ͥ�։���0;}k_n=<�^�fdn�v]:���l�Ap��vr��W��|�hO4i+���Jk��֏��d��/*kOu;����|�p�	ӜO��DJ�V^w,_�����������ݝ��IB�Vu(��
HWj���N�l��T��ʠ�C\�������~�9�i+�Q���Xc�U���+<y�=
/�u�F �v���C��fC۾���x�{�BC�Ɏ�tpʩ�T������h�����c��#�c�}f��k���X�9��5Я�u����j���4x��<N���:wW\v���&�`阖�kEs�R� m����u/)�ʁ^~��.�o�˾�a�yL�W��Ǣ�o&�ґ���]�TUC�WW���0���=��v����r���*ls���g=m��.M{���bN���Y�M�)��c� �{+���{��\� Ҹ��Ƀ�l*ڧ��`���T��9��P�7���
��GF:��G�*���/
����馒T`c�۵�y���4�ED�*�!e�Z� �4J�<�ʫA��~�NZ��%7i%�|G`y��īks���i�e!��af�R�״�vqO�6)�E��Q�)�]6�_����ё���[D�_�v����&�������C�@k�.<�;�oh]|Ε5±�RU+������������Ƙ[��� ����FTM�.eq~�%K�T/$�4t�79�7m���x֚����a�!;��h1�t�?pV����sՃ�
^��4�z"�7��N��_M��1�QV��,Jㄺ�*�����+c#��Y
�JPx(x�U/ʓ���N��d�p	����/�_1��~��v���eB��Ȗ҂C;�cʽ����ްn�"�B�����nw�����l��?T�&n��Wh�\�Tެ��6�o��?�u-�S��+��g&d[��Y��g_��E���]|B��v�!�BE��/U:��9x����ēC��+��mOd����I��~�g��~Z0A�$.u��|�Ti;@���pcX���޸�|�2L�e@`��ڸ.�yR�ǣ��~�����Q�:�*���.c Eb�g;7��H���H�ʅ5U����u긁B�����=��_��1C�쯠��ڌC��6�h����"2�@xuݍ�]��2�n��4�{���Qm[�yד���TJ��]����[P�U�Ƽ��ҍ���u+�S��x3i�f�峍�=,����/����YU%F�K�t1�/����E��Nʐg^��CƩ9{��@�=� }}S��fVG:�Tq^v�OB���5;�̔��If�eA���¸:�6	��!ek�$�0��WdW�͡Н)���5���B�F�X�����o	�`WpE=�Y��,^"�u�R�n��S��l�ߘ7K�N�؄ȧG|^�]�����w�Ё"jcgk�����L���@��W�_1xo4
�%B�Ael��y��c��lG״�C|�`���䅎�
�ڙyx���ٜ>��U�eʃ�oe`�ݑ7����䮃Gm���t�x�����7ٕ����^��an��fʏ��d���UI�R�'�{�U���8�S�[�cm՚#�&5�5�\����s��/m�:��xV��!���u�Ƥ�A�ȶ�'�6��m˩�zfj�)�fu�dݵ�yA�����;r����c��7v�C��V��]�E�=f�J)a�K����z/��N��x{)��Z@�!�*ǲ�\����у/��ȱ��\u(�2qK6a�̠��A-gsVlokX�U|��s�J��oOV��*�K�ݰV�),qM�� ��}���N�g�9��~�3��v�7o0�mj�rBU�\��P����n��֘<jHCGr����V<��w���%�ˮD���ɧ��
�L.ZRn�<� �u��Ya��
�XBXb��6Ml��IVH�r��d�V-dw6����>�kGl��-�p0���9�u($j�"��e�9�F��P�*�;�N�]��P�� 6=&��s�rK�ۡYק���8[�8��$A��`rV`�z���c��(-����b��u:H�XE����4�
U�Y�s^4��v��hL;�E�#�m�v
�T�X�E��	Zr$4�դ�4Ky���}��q��e6�s�v����]9v*i�W�:Z��aN��CR+X��b4U��g�h�W��:˚���Sk���&\��p'��H���wJ��t�fᮂa�Wg@�F`Ρ-���r������� 7��#�Sn+� ŚÕ� ���@.�6�{K��@�r���n�TU^�5%���;�,t�~�:�;�N--�X�e���M�G��WR�p��pR��)'ˋ��%[�ݽ�k-��B��7gS��5��tb���C��7.��S��ʉ�{n�x=O�@��)ȝ[�:�WMN���y9��29M��gWR	h�gN�6�ZyJ���\����=-Sqs��6��F���@j�-��J\��ǭ	��]V�\�n6��������֍�F��kO��%k%eh���ԕ+Zж�����T�%2%
Ȍ�W,�l*+�uB�����iq��*��-(�\ʕ�kU��ZҦ��2ږ�-�c*�"˙S&VىSMf*[J�
��Z�LDֱ˦�[�0CiQ
�U*4e�Z��\�.e�PL�
[bԨ*�l������"Ԏ�cq��i�R�����ZV���Mj�	jҖ6��D�m+��[mF)m*
[b2���J#r�m��s+ڵQKW2b�qj6�LV���QG30C+eB�K��F����0����*c��µ�2�-�[R�emm���Ķ�m
V�m
*Q�e1b\ɂF�Bڵ�c�(ְF2�VV��F#*X��m�J�,EZfX��X6�DLK��3**�(�߹�w��iϻ���K8�b���B�;�+�Q	���ǽʰ��Go�%�rD��6q�W��#κFP�:�a�{�s7�r�vFP���8 D�u�W�zW[X�:�`S�U�3�тI�5͒�ө��l_��*�2�.h�D��CχJj'G�/�B����[�����X.��T0ql*���9]���+��q��D���ȱ�֎g8��lz��1���X>�R�tz(N5N�>�N$����N�.H.��8Tt8����kRO�+���Qb2�UňW
�`�r."+�S�B$z��&*蕂��:�B���~�x,W�K�T8��"�Y
�(bgRw�9�b���?V�G3J�SѾ��vq���B�
^ȉ�S&9�(�U"�X]xJ�l�i�㛞hp�����[�� �VI>��!W�5�Pk�[�ؼ,��6i������0�݌�1�D����W;����:��+:=R�X�ٓWUp��gc*P�ͧXA�C�`�0�A/�y&zT䠷����L���0G���wK��ثE|��9��( 9������h�u<�Q��*����RS*�6Y���{�� rh�ML�ņ+3$�^��c^�yyE�n�%]*�l��Sg@��ת����%�����X֬�;Bb=!-[�[Z�W;n��\/��)Ͽ+���J]���l�ھ�3��P���x��m������S5q�M\�a!E��L��m�j+cV�eX�nv2��N�q��P�VG���ȶ���K�g�61;X��TO�y]��d�3��C`�(��eA�*Qo
r�[�b�v3ge�w�%�=���ހ��6<��u`�O��d��(-��G��,m�*Z{��`���`�z����̺Wm�Id�
PB�(	U��J�{ٕ �w�#�WY��E�=0�������C��u6���
3�.f����*!N�yxIT9x?��(e,��e����iA�S
R�=r��tZ ȗ@�ߨ2�6$J���U�q/�9��o	ۚ�cf�9/f�r
��؆����ء`�"�����\H�C΅���|�U�>�w�^C^-h~<)W�.��;v&HҡA���	�EI �q84��d���� �^�H1�,'ͯ���ӝ�LT��t&f��+��1QJWC�2J�[�ͥ�ۗ�2��^��'ݔ}�^LQVp
���Q����T��8��J�x>Zr���<Q�����3O>̝�H�J�P�+�+�0��i�۫��meV�)���^�9����8�`�9�c�����)�1�O�ҮX���E�uٗA��J�P�kg^/��$�b9�.�cTT��Q�1Cr���AH5�A	��8_�W��ؐ�=�h�5E���t�̫�YBU6Pu��@|4K=�IT�P1��r��=�m��qk&h~��i0(��{2-�;������\R��q1�3mm z8���hz�q??{j�f�V�J�*�=���ls�260,��6�Q�16���3j�Z��Ǟn�Z�$�Q�6\��21K��Jߕ�C��s��ʮ�W�S�\�u�H�s�,�#oԢx}t�$��`uP�
���r����vov����4���E��]�u�I��k����9���1�)-�j��X�����1{��4���5�o�J��ц��M���:���+b�y`�h���|'�b��e��);-g�\ Uشwӕ�a/�h�4tE���q=*
�Q��UNVF��{�3��/��oNz�����X�1��y��	I�W���;���C�-�F2����Q �uӺY��i�:B�����K�{z���{�e��܅�Dr��r�r���3���R���+"��)�U}v5�>Nw9�򪪪�}͈$�\��G��2�����A�꼎�4��5�&����鮪iA/u��a0��LG�D�2��Tm�(9+dҡ�g��"r;�3�C0qIm�%��>�<����<���@c�ׅ�z0X��!�qv���pm;�^f��8��ZB�gf�S��&\!K�Z� A�
��3�����u��TS}��rw�/#X��b
U1uCT�H�>Aa��U,��E�b�z��F70;Y�,=в^��@���3!��ʜ@�h1�@����Ben��K���9ir=��Y5�2����1 �.��'=ʠ>�A���SiK��K=[ef4Q;S�	��E+DfU@�'�Z��Q�eT��߁BW�[�g�w�)��ԧd�j���~kn;ݣ��ѲX�y!���qċr��X�޺Wm�qwSu�Z\Fҡp�9Y�8u:��<�BǀP���} 8���i�q �6g��x߅6�L�6�ַ}Ga޹����3��.��a"e��J����l	��#L�T:����v�x��nn��oV���:�r3�\&w��&��!@�+���p��LՔ����=��v���x;=��}�ы�J��:q�o�:�z�Ǥ���+i��tj�ʩ�hw���y:�mQ�S,�q�w�m���6S0�e� ���U�ü���7�b�I筜�~s<F��8���R-=
�ʖ��zd�%E	��"
�g(X�M�<��N`�&#�4:Ut(ѽV�ƖFv#
zn3ͣ�O�a���{��k��c�B�WQ�
���|5�q�ꗧ�u��_*��`V};�D{� $z�K�vl��s	��4���`�^����aH�L\N���K-=#y�����w����i7�!���P@=J慔GL��|��*�y`\c��%��Qc}���ch�{׉E�P�X=[:��j,CR�����]{KKQ�oʍ����'	!����{�w��!��gѱ4+��t��Dg����̟p�����]*�b�/���<t���	�ʀC����KS�J�!A��L�EdT�@��4�z޸��Gl0GL�xRT��;am�-f�\���M}��j0*����^4�e���\�1zk��/@��m���ٹ�p��+^	0�=��R7�A������d#��{e�V7���'xF�CiNNJ�O/��;)',��م*n6d���๧!]Pq�ͭ�B���j���_z{tꃪҧg%����E�k�@1㦮�\2�ر��F�l�C��i�ȗX���}ʪ��\��X[�Df�g�L�)pT*�IA�����T�yN��.�ݏ�X؈˓	�TF��{Ӂ�tLd,)�\���3����]�1I������5�p_�w~��K������3�V��@bj�֕p��|rJ���ao��Ai�>��(��㤫������U:��î�|t�f]*x��e���"��=m�e�T��2�P��!8��PF*Qo<�P�S٧c3Y�O'���į����*;AQ���W�HV����_�F��A`s�ǥn��Ytnn+��G<a*m.C�]X<e���lL�lu��ܺ��I&���lbx��L��Z�h�%�o����hG�&^��M��ZN�w���RY�uf�<��(}�긏��a�z��]�9۱�"�`<:3΅�{-���^�y�A�*�Hr����Z8Zq50���ź.\/���C�'��tT̥j^�Q�xl��b��j�m���u�m*�te�W���/���6�O;�rW���4���ȳe�t�1q�NÅc��8�����A�-�p�5U�`4�v��&�8{k-�r�.�{˄���2:��c�X��Ve>tƈ�>Y�e�C��s�AaS�Yԇ�h����d
K�ue������w��I��޶ޤ���h���>� �Qz|�����c�+�x�B4�ʌ�{S#1QR��s���tS�XU�����V-U]ax:�,R�� �-W���~yE���)�!���x��ެ��h-��u�(���D�٨!���W���6U��y$E��鹙UA���y��U�SjsqЂ���`Q��^ċ�ZwM`Tƈq~S�..�`e/0�Ng���s5��11��y[E�S�6�gˋ��=�q�a7��%���ڈq�*��qnx�<����ۺn��U����ҡNpʡ�T[�r��q6�LNOz����"��LXkS���$�#b��es�"�EY�Qc���$U��:w�WEb�+x�U��nﯲҘ��Ze���E��Zu�Hݛ|��]���d���2��{�[B�P���}Q2Ч�� N�m�L����ۻ'��ݞ�м�/1��ֻ29O�1�)] Q�-bc�|��}J��
���r:��8+��%ԃ��2�+̠Ǩ��<8V
߼�dT�*<�uE]
�T]:S/o�`��K��3��h0��V���u���3�]q���X��z�}I�>�-Ż�Ϲ�p�Ж�ǽG������3WYc��)�����8ϰ@�����s���^<�����ꚧ��	�_V����ִC�i��=~��wS�d���\�y�P�VQ��tN����pu-u���W>7��B]�~qž��{|��[��*�j�Wڨ#���)��>Z�c]��ΰ��K������E�@�ըE��6��}Զj�?�/�Q�|N�*� t-���Z[׊�Wk��̔7QG CA�����̟!.(!'e�P���ʄ�p}\19ގ�v�s��syA���MCu�Z��V������Ȓ�®Ӄ����<���i��R��7�e2���pUh��������k2�]V��X�k�lr��rP	��˲0�h\��t�&Ԅ��>�hVj!�y�jt[�|kN������$���_^��ӎd7�WL̚��o������6=�Z�3���6ȵ ̸�FC�TB�wu�����d��0g��@3�U�8A���s���]��A��e%�ʥ�V�xU�[BY��
7��m�~���5-I�}z��'��쭹u;�ˀE�Y����rB��0�k)v���X�nnj�޽���D"tQ���� N��hWA�LA.";
dT�7W���ͭ0�%���U����ȧ|C�F�f|~P�h�>:����!�{
�{��1�h�#�(:�������s������>�CU��ѫV��&Xǩs��"������ּ��=pO�ʖ�=8�Z>�Ҵ�8!]�3��꺲ִmQBDt����#�WB����7��u�i\@)��=�ӗ���*ޕ3}�ݦ��(h�C�`靎�#�A db������{��j6�bqme��U/�i\դ\L~�=CI�働����|;)�/��ؔ;�
�0��;b��Í-���wd:m�޾Dj��x�?{�dh��s��͑]���j�ЋOuk;fs$�벃��v_p�=7��цTo/P�H��H��ɑ�㭫y4OD�������{��}�Kc8�d}�T����C��U��q/��:I������'����0�qm�~��9ô4h���>V��Xr*Ė���ԩğ!4+a��fs��^���8��>��|��1b=��ؚ�qb�B�!�������?U�
߳�K���ک�K��Bk�
�]�*lڃ.��8P�(�)�'���CR�����%�^�����V:%���'��k�U�a�z�D9�v�P�Q�{��Z��m+��S/�+�n�T��Pl�)�ϭ��||;&���p���d�]�le�e3η���Tk�Db�v8B�ȳ/�E��J(@̒j�[u�u(@�T�N�ٻ�լڽP��PQAI�}���ެ}]���;�྇>0U��!�J&t��IQ�&L?VqB6:�fӇ(�w=.5�ҹ�z�*x+����Ȼ�S����!k��"5,[���t��O������ ��������h�"�h���{4]?����r�ӓWF��[
n�Mwr��e��@V�Sdu�[zV蝹��܃[�S�v��T>&��P�i`dzzf�����V�wk�廮�$�v�_e벷͌��f8��R*]���gN�n��6)5��fi�H���[_^��-ِq̈́x���wZI��1YP\Y)�훴�}��P{|s���P8������<ڏl�#�άl���xC8t�h�]<��oD�n�hh<NT�Ĕ�t:��S ۃ���G~YG>�F�M����à���i��p���k{t�9�5u��Y�Ux,.j:|�e�U��pM�����w�W5��	�o�\�aW�i2/FRc�����6�Z�u.r.wM�,�y<����U;h�+��\Kq^�_d<��s��y�8�S�Lc�>'��Gv�G'y)c\�7��V^��u�Y�N�A��uv�N1�
�o�K��<��+(���m� �ͽ�:΁�Q�ԆvŠs���l�O9��#���5�|�*۷��^�1a��De��X��҂�@_ù1�gP�L�,���ʂ00���^H�����<+���˟t�`,N��ء�d���4s�R��l<:����Wε�[���N�� )2����NtZ��t�z��̂�-��U�9�{���jy���^�	�M�+�Op寈�yl����U��oIaJ@d�iJ:�/J�Vr�[H71���
1��Ö2,j�9�mb�Z�y�0)=�ɭ�*,�M�����b��`hYwB\\�� �v)RYsr���J9r���`�b�۟ʸ���R*�-�)IB:��h�Ģ;\�.�;��6���ՠn�U�Z�W��WR� 4�ј� CJ�Y�J*l�bs1捈	ur@\T�C)5i`��-�%]k��P0%ٗVKOP�U���.��!}�m�W��i�WI�Ę�KY+�R����[y.�D.Po �o0 ��*� �y,�`�2���,2肌u�R��Lr7�*�шSG��#C��*2������t^<�XjNCzkqJYc�Y�ƺ�=��;��򓣣�l+˽%��$l�s��k ��8�`!;��6m�+A���hٜ����7���o��*�rFW*ᥪ]��T���T.�_5��:]�zt��:aV��~�G�l�6n,��e��O��T����k��_W2�:��g��S{]�Dg�'�a�@i':�i3��qQ�8��q��;
	����ˍ�Y���+^š�l9y�:0�=,�fsT�1U����*V�q�2iݬy|�(�EQյlbFжږ��P��\�q�h�F�T����mj��U�R�5�YZ��nV��Q���DV��ь��ڔJ���3(8X�PUq���Bڵ�Z�������)Z��V�9��UL�3"��j���RYp�"�3�.%�UX6�)����Ԩ�EQE1�9�0B�a��!J)Kl���cK���-qŅ�����T��S2�Q�*-�T�J�([KlPLs
V�5UeJ%j*Ȱ���-�6Z2��h�KlR�KZ�#)kiJ�
0�҂�k���⡍��e�J�ʈ֥Dhŕ�[F���T�+Z�e��J�amZֹh���Tj�������LI�Z���u׹��ν�_;�����N*.�FH5�M9��t��8�q�,7f�]�
���][���Z��^���2��&��m詶`�Gmn2f�� ���\�jwU�,[� 	��-�'�)A?B�+=F#��?R�oZ��~�'�δR�Vl�/x�A��nm�/��橦:�M م=(K^�[X��T�]�G@e�� # �/3T��{��ӱc��	W�����]Gh/�,0��W%@�M�Nd���޼���QC�����#8�3\��9�r�XM�^�:�r�Z���m��[�\隋����Q�Tn$od�dIB�ߤ<
�b}��18q�$���8���D���e�r\��n�d3ꮆ�����ء`�V��O:�޵��}OUm(Mq�D*J�����U���3�Ä=�t$�ڸ%�h��v:羫Ц��!HX�l�GANֆ��<l]H��L�K�39
�=T[x��4]��c݊�.�:���,R�H5�WD�x�=򋗹6��=n�����n"��Q��fm��������7��%R��A ct�i]K ;Ƭ�U,J 9$�Bz�n���˖����f.�V.F�6�d)�>�KQ�U�YY�R��"�H8��.�ug8��/6B��I�'8���U�i�X%��{2�jyO\�`�f��@{�����$hI���;�\P
s%��������u�G�^�+��ά��Zp�^�(sh�5�̼�b�Zw$�[/mMu�/y���7��q�3l�tV1d� �)q�*��͇�G9�!��ë��8��s����}[�Ǧ�͇��*]H�X#b�W\�H9�F�D��u<�Ύ9��g��]�e�}��X���ސ���kD��ʞ�K��c�]�7e����lh��mS�-��C�a�,=j"�s�6��nЭ�S��
���**Bůp�P���'�=)L�?/C�Y�
�:;8�L�K	|kEs��uxC�NG�@J��?9�+������x��k�����@]L��X���7R��^#����Q'(k����r��9��4+���a7��j�>��<C�9^A���9m��V!�\F^�C�;W�_��Չ���P�WD
#�@��t<넳�,��Vu>5��4��'8���Q@�Ok��5��;�k�n�b�f:7�W"�c�y�E��(��$)<wd5�U�:sk}.ұN�$�f1�A��Yu����a!7mE�v@D�y��j�w:���>Ux��/j�����%[�ML����Q��v(E)pr��>��)(V�FW��B��U�{�>;2^'��m}��kܡ+�{
�����K���Ғ�E$@�1�N�9����åF1�NO�Њ�ņ�!��5�\�B\PBN˱T/&�h-�b�O-j+k�T�;	͍P��}��R� 5j&�U14�:�,q<U�1���}0�8z�|^�u?�3�(A��u�[�б(w��ʠ>�hs�؁Ow�Q]a�e�6ܭ�uJ+�l��$8����\�/��#o��]�;r����{��%�j�4ġ���Y#����Qz��A����njR�t�XJ��=j{�sS�i��Һ�C,���'`��+��t�OA�"uk��uDA������]���"�<�����O�fc*\]m8jq"�&Suw�͹��!\=�s=ciC�9 �#��V;nC�����aP������`��M-7#s���=N�J��,S{WD�D/�����Evcz�H���\v�X�r�o�8��;��_]v��<&��Oij�u����[���)�[ǖp�kA:���*ɓ����c�y�v_b�z��N�:68�zy�W�}��#}^�O)(~#�]�W'�����}��A>��b__b��a��lR�}�1��qVv%�}B�Q��R:�������g�E�Uno]�U�
���5��2���-����B�}���;A`gzLmH�"��a`���,˾�\u;���R��X�v >͂.��6Y�-{����:J^X8ς��Dχ3�}jͶm�TL&*�(;'�һU;�<Q
d��'�hS��S`��Trr){�����-�L�'�|�	q�DC���"gQQ�EX�f`H����Ap���Unr)��f$@��W;��eК(� 9��!��.6&���B�"܋��S��<�L�هgJHq+�A{�,עVo�����Y���>��o�'YN��Ч�r����j*X�>˩�A��2c2(!�9i!���,us9p��Ǯ�,��z^C-}�E��B�n}^�A
�Ơؔ�o�^^�z�i�bc�}}���ɢ�p�QA
���U�˽��7s��*���㱂1��DF�f��lt��9M�C��F�cI�ʓM�v����o����vN�,\�9X��4�x�9�MҢA�n�l��TJ��˟ �E38.Yg��xC���+\�S�0�j7R�X��g��[�\>�*RPx9�<D"�x�������KD\(�򃈊&��ln./z�ϫ�`ù�1�)I�=}a0�J}��$К��U�m�9����K�,�b�Q�����y�Ee���on�`[�+S��t2�C�Y!�Գ'���N:4�*f�\[�y��;D�x�ӑoj;O�d�R<��M)|�S�č0X��$���E
�H��TT��2W��<ұ�k.w����c��{
��ډsTw�N��*��� dmv�hW���yP]����L�C��~�B�Y�9-{�&mC(q�����n��U���^��^�4g��C��1�P94{�k5�W��7�wQ��y`�go���΍������|'�:Z�tK��;����L�x��o��3��t�Y�Ǳq<�"&$:�x"��8�0!�ڳ�d��x���x�b):Ƞ�w3
؉ij�)'	6���ߔ��J��g�F�j�ڐ�k�{�WJj�qʺ���;��z���"����|��w4��ۥ�@T�ź��cU�_hvN*,�@CB����t�!vj`u�٪Ⱦ*]��Y1�'�{�قR9h���_{ކow�sg�~"�D 5��M�N�
t����B�D�p����$]�joV�9N�խ���Vog�F��4�'��!\�w����b�><dq�E����c�p��&e��u�3�m�dT�JLRȯ�X�B�k�>�E��ux� ��%4�-�׼Abo�p$j`�#�{~��҇BE���i�=�e^��h�R�3֓F�ቋ����0�����!���#CZwMcU1Z%�,z�7��	�-�-eQ�Ӓ���
���q.
Z���=5y�^�PX���$�v�f!:پC{M�4���U�2�x/�'�3l��±���1~>�(����9�jbP*�Ī�}6�w(�v6}�3`�^>ƐT�J�?�\ ls�� c�U���t�}��"�ɓٶ�(��k���H�����$Vф,Ut8"ؠ\��Qgb��mU�;��F�8�a=�tV�u�\������p�Ui8�Sp�X7�]=2Z�RF�Խ���o���M���yћ��N�e8�	�����9�k�s����V
�T&��52_.��m�/;�-�{m����o��Q�yܢ�Kz���A#x_7;8�H�ùg��^B��ミ#�r��\n���t��v<�x���LxM:ϥ_0�5�Jq;8&T�)P� %
15�]��ɱ˗��o��|}�5�
ue�q`S5�Ɍ���c��4 ����F�G�'������n����_h,mb�עF�"�L�8���d�[+���w���^k��(Q���0E-�Sʸ/�P}��H�C`r�=3M�d���]�g�!�V􆒻ؤ�"�ˉr"e���#@`��>ZT�Z/ݔ%{���Q���ĭj�cQ2i��U�M� 5^§�����%����薂)R o�X^f$a����{<��14+�ᰀx�*����`�M��2p����~��X��<xI��BK�77�j>�t:�[ȸ�VTI�����<���3F�`�[�	B�ʭ�T����g�C���^��,A�8N�e+�gu��>�>��X>�dYm��N6����6��\[��\6.@����F����Vk�Y�����z뽆xCF٣��խ��ҵ>��p��)8�g�Vq��oA����-C�vg�,��� �=&�[6bf���g�UD�̮=�sqM7�w)����;
M#
�S��[���P�w&qc�ns�7�Z4X�Hgҏ�����8+m� �����Y�f(ղ#�S]�-�F�,��j\r�=�8qV#s�L#jǽt��Z;x�|�Ι��-;+({�> (lw��[�N{�ezk�#:[���
�m��Q��ao��z�n�7jV+�O,���+n햐�ÿC�����j#Hʤ�A)nmkJ����@U< �����o�ҙQ�m�k���Zzg�3�.y��gG�!�R�nMWdK�#"�c��� ��QtGY.�(�=��m�\@t��:�zW�@l�9߹5�w\�;�l���P��Gh"l ��pk��փ��]�Ӱ�:-r�~ɚ�cG��I�[=�8lR�΢1��W�x��Q�O�4~"����I:����Ҏ��8^����T[�j悐�S�pؗ3T�b���Xx+�W�]=v�C�^�𬡶���UdL�*5ȫCT�H��T�HBj�wc�;մ�\m1��*��V�0v����� u���vv�B-H;��k�D�^h'Gu1-�Ǥ�V��!\�칌@��_k��f���w�θ*|/�^C�P�p	ٔ��^gE�+�gB���ْ���%����������I�мE�ҏ���
��9�9x]	^5 ��v@������<�EV?�	����������'����н�Hp��=�/�V�Vu���DpyMXؔ��x'�sƮү�T�x�pv^�u3٭�W3�h+Pe��1�׊֟��h1�3�%z�yxs�o�_t���坪5����.�f�������B�u��}vTJ/�ͣ|��;WKs�]̙�������^ :<@ԍ��J�*�Ș�jB8)�Ԭmt�#>�e]��`���fU�����Y>��K��6VOF>gb�^t($O[R�QKc�,D�R$l_�tɆ iT�}������Y��\ym���4����Ό�����x+t�4��A��b�P�r�T^γï}�lXڱ�NީāP�+�Ϊ[5`j=�C�	����&�uM!X�U�m�Y�mq�ml�g/z�9�Pf�Keͺ�M��uP�U�:�����0����K@�x+���t�Mf͝>�O/8���w�xN�e��4"�e;���|��ˡM���;&cNJ�@�;���r��y9�<�xz�w���mo��KS*��#jO�
P�p��[D�p nD���|���{��x!᭭���:�`)��3�k5�������u-6g�*�S�������ٟ��qwS��b��B�գ��x=�.a|h�9U�]ul�~G��y��o����b�k���O/�|+������0{�����`k'j��9��me�u(��q�F��,BZ�>HpVxVuZ�`
��2M�A���z�s}F2#:�@]}���ӡH`֕��Mh!;Zy�s����AgM��A\#!��b��;�Ǽ�ˇ�`�^�b��ޗǷJ�4� ��z�Qf��2��_(�w��u����r8P~��]�uZo�~V�{*��7�ϒ�Qg�����'6�1{Y��=��V/bE��t�S1�6�C�sI%n�B�{/g�c``�DdL8�/)�{���������PXUTv�R�.�����Px]ޙ�r��K�oP`�1#[]�;�o�j�n��蓛�eu�U�m����O�v	R��q�y Z^�{����a���s���^̃�������9wv�G��*4+u!p��&�g9�I��m�bnrY,^MK�v`a�8�4e���a3�#�9l�+#�Ilbb(u�q9��:��c��4��l�6b���#D�/G"���gi�EI��MF�:I
[���n� H/I� �u��y� 6��4�Pɐ�4y�qf[�۵!� �m���g���!!��YN��+)��452���)1V43P�n���<MnF��矲�ɕ:AW��&>�8w.�՗J({S�+\�����x���+T s})cʵ,�sw1��R�79�.��7L�@,���EG܌�w��iIw]��Yѝ��X���#�Of�4�R���U�hY�&�5����n�������˓yl3k6�?1�JAܙ諧E5�v[�e�I�>����eX�[<��z���%s�Tko���2���w��z�x2`���93�<��^�i��;k��Z�o"�[�m]
�UL��
\c*u �q�C��.�-���-[@�/>3Op�Vp�,T�=w{�yN��������Yr�w F��9�@�]�}e��؍ m�K�[	fW	hR3��U��@����J%�ӹyV�`�y���	9T�������c�>��Y�J���2���)L�>�5%����tev_k"D��ka�u%Z&ڻ��8m 4*���u��ۦD��.���u��p܋61k�}8V��qIss,�judV��WA.�(�7�&/���V����xD���T6( ֛�>ܫ�vH1��cVʱW�q��Q8"Yr���F�e�V��P.�h[��F�iƬ�`�Ŋ�"6L��Р�<V��!:ZU`��xjp�E2!���5�(;UW� p�A�U��fX|e�#�,��h�����Y+hxc�L.�;b�t����v�í*$�(&T���ʹi�>1�@�qk�1�^�Zn��E���x�vhq��J��*�E�;n�7�Eȳ�ܫ�K�Y!V>p��(.��겄��˰O6_gm5k��U�E0�|�(���1��E���j����RwC��&�T�3�;�Y:.�����z��p��!�#�Y��v��{�zEv�@ÙB+B�)mGj�`Ci�#� ^�"��S�Ĝ(fd�d0<4!/��mR2P�,�(�+�跋�ƤZ;u �La㥽���cUJꗅGn5ˉ�\=�+6\u;n�\c���u4�ysL܃�p�2�@`�H�D}D���
����U�F1DT�hVTE-��,�m�[�PFb��iJ��cjR�E	P���4�D��Z�Q�T����(ƶت�EP�ڰX��V�aEJ[Z�R�Q-�-�T�ڵm��T-�ms0\IYX��kHն�.Bր֕��ѹf+��Ŋ�.XUq���-��Kj��l���Ki#Qm��j(4��e�aSԭ��
UcF��+[J���\LQ�ִm�Q�6Ъ2(�*�W2���QVF��b��E+�,�KT�U�\̘�jc�ic�(����2fb������",eJ�E��j����
R��2�T���s�����Ԩ�
*T����2�ZQ�~�4E�s1��p��G�����X���|pR���}��9�ʔ���T;�ٍՙ*̚����W6_.J�g.==�_��ɨ
�B#p�V3�����.et�<�j�Tm2]����p�zX�u���cgT�>�\�4*�lr� es���eg���grD��2Vp^�u_��~�/Ʒ��ymz@0:�;d�C�����
��̸Ɓoo:\@���Q���p�z��R������)��e���V��,�uzv��_����n�A���E��]Y�4:��g +��ޮ*��>İ���-��7����t�b��{	�X�8�K�q���
�P�������;KG���G�<U{�l��ű��|�G҅9���z���x�[3��3���]>�?;�%}��g��Q;n�H��J���W�z�����7�kW�����9�:�����zxR���G�xG�����#���)�kE�KxIG���}�s��L��z�K�9�$WR��6"ڧ�VQq0�˄��KAe	�p�%J=���ܘ6�G��j��w�M��z�wT�`���U������K���|xի��b{>}i�<D��{��漺;ׂR��D�K��a:�+�z�v!ǩIv&XĖ�{$���[���|%ݸ����!d\�h�6v�N�Ⓨ�����j�p��
B��d�K���LXj�q�.��ľ���@�6��3
�w���fO�o����x{�e:�����\D�n�fn&^何�.\�/X��C�Ã�>E���Vꢧ���J�6<=R���`%˂�-�-�i�.�����P0ldx:�X:RS�wxHp3j����,7��j����6}ڧ���]���m����U�۳~�t|73�M`s���^�[���u���7}G1sg���r9ģ"��d�=�͞]�m:n�.gg`�������1�K��׻٬�i+w*�Vu��À�+�W;�\�q�����\���+�[���:���4��a�R��/V6�9��B�#]	i�p�l\0!�u1|�jY�Pr)\���BءB�mJ��g���9�<<���bi��0����l�j�u�f*�niđ(B�>��+������$u�=2�T۞�C'������xh�d��U ̍ds��"59�Nr�yt�z��-��	��k-=���uwFdG��>���RG����ؒ+�����p�SX�7E���]p�\^���u�|;3lAK��#nK���ܽ[|�2��7R��*�ئ�7�(x_Q�G� :9�F�:^�+�dڮok�=�M�Z�&U�,t���q}7]De>[
ۯ�F{���I񱧅(7f��{�n���#��v\a��NmM��U;��݇2�5�����qUjgE�E�o8��Ȭ�i������e���9�~>��j�	iӉ͡����a�0�� ]?n|+&T�.O��')B�ɥ<	pL�ؙ�bB�"�;;݃����+��N� z�,�QU�C�]�$,�3�-��"��.b���Ļю6����֖��s*H���Y2}��RC!���0��5����R��Y�"�&��!�L�!���h�Nc�8�N=�!Mv�j%���o��#(1\6�Ao��l5/5T�4�wRJW��H�h���`ܭu�6��0͇�C�QP3$�����4�{3<���z���kh;ġ����p�U����WE�ߡ䅚�2�42�E%u�4/��\(6re�@j�.�Ӕ-w��k;S���X�	R3B�3�qǺ��4� �uҎ�S�#vc��:�A�lQ%]jҮ�o�	417����{�ʈ�BX7Sn��ʸ����x�œ�ܰ��Nε�N�׸��a�\~�������>�7�ᙷI�ﯗ���<n��?GEY�n��Փ��V9��zi����W��&����ѪT��q�Z���%ԩId��9έ�0�ڎŭE��v)�4�t�>�F����5��n_>%pZf�k{��C��t;�E�T�j��ৣ<�g�T��y�HV������"�2I��׽=1���=�(S��u��κj����)Sz��BTB��8�mT��J&%�?�ӗ֢�cQ��WG�&�+�\33�E{s��3�"���g�]�P5롨B�}ʎU�i>����>5A])&,?�.���_t����*;řs�12�˿G��<0�P���#+���ˮ��t���K���݅[�F��)��5i��J�f�P������DW/��WL�lZ�N��pY��77�(a�o��wm��r�:Z�(�p��T��Ě���1c�XO��B�É�ŽT��i�Ϸ��/}��P�m���Ŏ�
��ՌmƠ��r�+0cj�+Gm��ue]��39B��j,�D�\.A�ِ�Q�6��ǲ�a�Ed'q6�G:c������t'3�n���x�=��+�t|{no.sW�'1�/E�sN�F5�RiÉ��ȧ��
AU}�;�-=�ʓ�jb�ۊ��� ��> Vw�R��������Ͻ����V���3כ��b*&��P�l?�U���F����򨆗 �L��>}�1�x�*B�$�fj+����:Û.,T�
l��&[�5Fl�r�᰸��sQ��'�EiVf�B����8=��E�s�t�Á��%�3�W����%s Oy��_�y�HOVPNz/ͧ{�\Q�T+�T�5�\��	�#�ܡ�1s�k\gƝٻ[*e����zowюGl���L���B*�rjU]75UC,.���6�f吮�� i\�r�s��E*��j��0i�:뮅AM�V&2(h�~/2��~�K3lJ�"�h�K���=�������>ϼ�#����W�֥����xO1�f�{��b�ԩJ���ǆT��E�8���:�Pd�`M尰jU���_�,��%�ja�7��[z����+܈�Z�Y>��wd�.��ofsF���g%�\r����D����{M�In����49hۺ�����i�n�P��ӳ���(��5?�_Y��Î���t�U��ӻx�wG`>ឰ��\�:��z�pڠ`޳PY�fYt��؜/�֛q�g�ձ��}��FeN�T���W��(p� T/Ad�w`G�� �f�B��r�\8e�}��ҡ�gh�i]钝�ŗ¬Z���(\"�ތ�����m��b��u��:�9$�2fv\��b��R��E�R\=A��ؾ�D5�`�'����yQ�G�xp�G�� ������1a� �ƪb�$��9��s�u�ef-sĿm�|&�]��^Jr'�Sb.9�j�&��!b�q0���u�w�m���V�5�p*�V���R2���\4��i���ń=OPh�;����aS7�	��W^�A[���0�hkƚ̯]��f,��Z�^��7���J�r2H�E�gzp9�ظ���>
�C��Y<�01`~�g�����988m��'a8�v1͏Cf�,=�+��W22 h���ض�"/�M�Yt5�#Q`xP7�Ɔ�{��a��ܒ�8d�s���'cA�+%���p���z2����K·���\Xpu�u���nA�����Q�\J�}�_h��UN���ݛ��IV��+��V��� F9�#\{���xv������4�V�,yu�> (lw+��;
�:�u��m^�U�k)��x��:I3�8
��WA�NeX�p�O��\+Y�V�ۇ�C���gjtl��N��j�VJ�j��$�ԡT�lWA�JeE��qˇ-�G@s���z7�Mol%wGr2�.��lOL�CF4�Q�uWPt+G*~N�.zO	�U�OCե�O��Hb�^��
ϯ�u�M�*$�0!�O�*�"̾�u�7׻�����ԍ��2�ٵ���Z�ۿs�Ϲ�F>Y
�S����>�p�Kˇ��=V$Q$���o���Er:9���3��V�ب���в�S'�������E��u�y?t�&����^	у�
0��U�$S�2M��.�D��Yy�yZi�U��[Ah��POT�'ʊ��8@�2��7G�:�C���ѥ�6{=�V�B��Ӣ���%�RU�Z��])!e}���v�S�EO���&�ֵ�U���£;9O�X�(�U/�J��A�k0����Y;�+��VW��̨`v�}�mo:~�,�٣��O<��R�0s�J���U�+���d�Ww[1����֭�����x%�P��`q`Uy�&Ӌ�7�8�k�]�;#�l�u�#�VS}�m;ys\�KW��"��5���eh�f��\m��ج"��Z#���X:%�\
�͹���,����g�w�B�,�����SC��{��nW�B��pC�������p�J�Qkf��]z6昜����0�k6
�vg��lc;f���_�N���^=����R�rPh�]��h���xz�� 41�[i��������SY�T_�=Obd,R���p@ʚ��xi#6�9��p�rk��\����
�r�nV�f{6T0�;n�B�(�ڠ� ��1@�t�tb�3�\[,f�0���y���#y]��*��Zv�qI�.:꣧ ���u=�B�@N$t�2�s
������ܔViB �^�TڗY1�R��;�Ŏ:%*;AQ6:�����I~�5����X�]F���+��T�j�<,�z�R��:��k(J��Q�}�?r��e�>Ä�\2�cGF�J5�:����㐌��Nff�NR]���
7�7YƣPq�r��w���$���#�fB��WT�1��L�����x���wR\�pao�'s���+�m$$����Q%���Q�+8<M�/	/	���eq�Y�w�K�¥��d�W܏Η���{����p���������G��(yx8E�^��;����im�G#i.���1t�XU���4Er�P�k�5㩖�VJ��C)A��F�1x.�<Ƣ�Dc3�L�-K���pE�s�RAv�J��B���,'��#�Ƿ�y���&]�cC���b�7"foy��L���p�"�p�!WX^h�]f���{i��`�3�9��,D��1@����\�h�/H~��T�>����F�%״"*�ٞ�;���#0X�9�T���a��[�ܣ_��0�!�ZL
J�D�U�<H��9w!�X�s�݂ٱָ6=wS�+�h��5�zn��P�R��i{�.Pq�>�w�Ows���J��F,����>+P
^9�l�/�|+\o�Q�X�
�9
���zZm�[6�Td��ǥj����
��c����Ҷ�,O���Y=N�hγ��Z�4(���[�w��q+��V����eCT��� 8��63.��b�%>�z�����<�)a ��`!�ܠ0wL�"��u�v��)���V��a
�쳎��o��.��jt�NY���)�x�OSޥ')8�̋��8X�tP�c֣T��OB�8���:�Xu����]8+h���w�|��˄j�4+	: �u,yZ�{�����~r�:#������7%s|j�jq�H/����H��t���P��%D�S+$P����ͧz��4�iLOC�ѹ!�n�]��1.�}�V+�*YAQ>��"��ќ_	�8�T���_0(�n�n���k��i��K.��I��ԫ5�9��?e
4y_���f��>Z����3gCb.�(M��|i���:��&O��.0���%É�ft��	��1
����s�S���fs�ڼ����3�.�"�j�L�����|.���*#{/u��	>!L�gp���ZT�c]�x�Oΰ��½��b-�gf��S��&\d�L����ogg����,ߩ,Q�C���6��#�t9�L�ШX����1YY��c����A���v��t��%V򢝹�P����{H�^��_G�@�f�]@[	Z��� �.��j��3�o}S������"�osm�H;���n�r��*Ç�hiP�qBj�k+)��vs��e ��]:�ffGC��y�uӲ�Ȳ��w�:"��������5�$*�]e�K�|C㣪r��h��M8��jhИ�zE��|����gOz���sU0�x��0J]s�qN�.˦��0�yZ�x���(��+۠Uzo�1,�o$��l���Xym+���'���OH���2m�v�n���W 6x׼0%J�eN��׋/
eiL�
҇a�R9�w�ޥ�pd��q��5+Z�J�3��qw�ܬ��aڷ�֍9j:��wI��/Bk�N��*f^�v9��-HS�0�nc쨀� .Ɗ��u�O�z��;r3�:՛y#���;V�wuw0ɕ`�V��w&hު��<��[o���*�R5n�ʸ����/���X��+��Ҡ�Ǵ�4�)};hꏅSq!���7k���؇dV*�s[Ɉ���)�G]������������.ނ���n�;7�&n�6�YVE��' ��n�9�@�r`ə5K�"��9�������o�h�V,�'�N.xR[m�hK\����#%���d�{�.�0���m�"��V�u�^.���v��5buf^�.�}E}Rj��g��*[�*�;SvD�b9�wʻs�KI��h�]��_\�gJ����Z�mT���Ȃ�d�����\�엸#������K`GR�t�{���A�$&P��o3�\b�rm=��v4U���x��Usk�A�)�ӒԺd$E���6����@��vȎ�e�k���{x�\�*v�a��Md"���Dn/��J�/\�ckNH �����ۨ�ӷF�Y�N0�9)G�鍖���-֢df��*L�(��"'�l .���u�|����^wW%�B�b�P��)��n�X�t�pU���@y�
:�U���(�ZJ�hЕ��vڬ���ͼ�]�(�p٥-[���X�ұغ��Z��P2yV�z�U��v��6���l#�6�/2����oK�u:ʻ{%v��wP�\�v�仦;M��<Qz>K��/6c����*躕�۰��l�S�o%o�z���ï�X�ιҠ�r
��{bJ�Y��Cw�rTnKӜ����Gy��']����1Z����Ȗ��h�i��w1�ʜ�V����~�����2�Z�UcmTb���*miDKJR�)i���6�Z�E1�F8Z(ULn6�m����U�6�m�d�*ԭmm�ڥ1�̵�YD̢�-J���l���1�KiT�P�`Ҙ�1�R*�����e�&6�Q����,E�Q�EYKQ�ʠ�e10Qj�eˌ�8�PX�Ԯ�-�ET���-rࢢ&YA��2����""���Apm���Dk�����[�����\�V%�B��(���8��-��m���*6��ʣ[�1�" ֕-J5��\˂+���3&TTm0��,�Q���Y�EE�*(嬮8��W32ZQQ��3�*」J-���R�eQQ�E�J�E
-̘����EKj&2U�	*9EA[k��ªQEn�ׅ���}��{:�宻�U�M�X����㹀��7#ǥ��/�g�i}q5a� =���*�|��h���wb��1]�~Ix�Ă�Ey^����!ٳ�:t(��h�Ơ#��TAI���Y����E��\,V��L-�k ���UY��N.�~u����Ej���c��Ws�No�uY�z��<��bWg�����J�� �.�qe��Crw��-�){Ɯcn�X�Fܸr}��9�;�y=娉>t.�5�5�
�uK��%z>�-y
�=��l�H�j���N"��J&��g�<*�C�!�Ȝ#��z]�6��=�>R�OZm�a�R�8�v�G��f�c�tz:V�>�1�Cxk�q�i~�o:%��6�Uҹ�J�R�
#h*F�\�X��T_�Ӄ��\J��3*q�W�3;m*�0�p�������Y�5�C(Ҫ:���
��Eqٞ���M\�6x�k_<�v�mKx�aT@�Oo�U�M�Uh^@x*��������6�8ߏ?K���9�7>bx��4T���ڮ U�d�]s\�Lw���'��gJud�K���:��%s��-�{FJ��^�9r��5��哱in@�mv�v���.W��yS�e(��w�����5y�]��ZZs�im�r&��v1d
���gJ��٬5�]�M)��f
�V�`<�w��k���}�ۦ�
�֍��85(�Lo\�1c&��8,ّ�?��a�><1w�Z7��Z�k�*C&{�i'��5b��&�W�ﶍ����
�8V�G��}Z�E����5!��Qw�J�t��&��"��E{�dh���2�t(�(�1�T�\%��ѕ����1גG��Y��,~ <�ER��ؐ�U;(ej޺���O��:0K���������Q�o��bca�q�S9�ȩ>dxWY#��i��%��A�R����=y�wr�&�H}����0���AS�d�{��Z`"�����ܯe���|�D�4����e��3�6+��Wܫq�&vg�d�a�}%iW^���o+y�.���;`����4a�����C�����w�TA)�Խɥ��@���{4m��e��YKB���Ш������
Z�������G���i�6��F�Ű����֏�ٗ��=
9 ֒>�����~(F��S��/�g���v���U}b��m����r�X��H�Qls/�Z��b�.����`'f�=7e���#:ִ��07|�&2����qG�x�����+I��C1�U���-�U�5���`'w�:1�d�~V��tdN�!3|P�I��]+��F����w�:뢆7]3^����)�Q���M4��@;0�E���T��bL�GO�W{^;��=�Ǜy�a"��@*�w=́�(t.���u�(d��J�f��Z3�Ma����B�V�ZX<'%��4w6CL\����ٺ
B2)�"u9�K�Wr��N�o"9x��)ey`�e^��T�t�I�;:������7=�薤���!�ᾋ��1�
~��� 4�n<$^<�6<,vRz����}�y���5k"��qt7�#�<
������6MJ�|q6t:��@>���z��3���{3�_C�Ϫ��IK���pE�s�D��_ �)�N��;�`�z�錸�}ENDL�Ј��b�'V#|�VB-p�!u.��u�$]k/;���P�X�c��]wM�鈖%D@Z�!�����&�$
��y���NjT�����h)�ʇ�c�_v��?c2����fŶ��|�)�[��p�WЉ�|���»��v:��p�M�ɢ��2G�(�\�[u�C7���]#����6>U�p*w��K(㙷9���茻�t^�j���8&�u%���д`��J�,N6'��-������|���T
�:WMN��U�gW;ֶU��Ź�׫��>�B����0�D~�ʜPܟfю{���%��i"'�Lڙ�9l�b�ܞ�֝�8#��_u�(b,xR'�}v���pC�{�9�f�R�1�OC��U
{� XOv`W\�v�J6���M`hF�c�0� �[���27WPX��h>�W��<5o���]ysb��vf�%n*�+�k1�x;��܌u]
�`�Xd
�{���צ�Vxhˆ^�>����:;$Bh��-T+2H��]WB�n�n�ʱ�.b�r��Y���HN3Q��2eƻ����\0�{3�u�
�����z�á�.M����R�u\b���o��Z�k�	����H�9֣��+Au�����g�d�U1����]�rC��.g�u��|&��p���F}���
��P�꺈p�Q5�4������ͯ^�u�ia�um�[�N�D^�k~v����:��Z�<��̦�sT30uk��$፻�R�ӝ�Y��aJ8�Fծi
Ss^��y:�Jٛ\�gnRT��RqBNRq�T���#i_��}e�N�
}�4�[]w�rۃqB�8�t"R�a_M��Ƞ��<mg��1lH�FO�Т&��)� �6d��Pl�Լ�Qq1��5<��3���T��!��ly���<H4/��0���g�1A�B��FN��O�"V���\��夽��>�0�%V�t]U���,8*tD�ި���inI׽�9nH���
� o�r��l:���)e��P�"���f[�<#��v/�z��%z 9}����x2}��k��+�q\?f��w9.K0����݁��@s:"��R�;K�1kY�9
͟�0Y�T:�<d{�S���yw�Y�YFs�FCf�b2q�E�0�����)��B\�H��_.I�e�>QX����14�|}C������j僰K������j4��syMU]G�-ӡ�d��q��&M��q��^%����tz;�Z����jL�9�A9�@�@n<[NږV"�V,r/{P=@G#�}�t;�k3���^ֱ[9�G2�H���ŝ�q��}�����pPa^+}�E��Tú��;T��$����謾(f�K�Z���y��Hw��7��9���.�U����sc����Η2C�[��Z���'!W��^%a�>EW�T�F�"�d�X/�̨ᮜM���[̄�gm�q1��hуLV4a�h���Atz�*YB��A�Nho��9�[��\퓅ft�L�=u�lj��b1�'׊u�=<������<���c]yKݛg��?yj��i���]��@+�g���xo�^�}���}KDaB5ƞx��r�hؤ=GWC�h�Z7��L�N���#��������u�$훹��������V��R僄^Z$��N�gE�ك�Μ4_ez�;�H?z������w���:(�T� ��J��+'C|���g�
��t|���;��]+�,�=�V�ea�(xx@R��_�ER�.�l�����E;|+�v�m5n��\��;=�d�f�vdLt1
#���{��FR�
=H�X��e�&WUWOo4��Vb�~�od_a!ō��N�P�Yަ���d�pV�E�+�̓8��+=|���ڀ֌�e���[J��r��Ѵ�Z(�����ļ�1�@��<9;Y+����k�����z��]�wQt��+�=s]�X�^E�%��0��c�8�طB��U\2#���N��E����#���������kA�h��y���+n��*B�+2����mpux�=S�DA�M�>�F��GOy.��8ʺ��T�U�u!\��E8�\���@���li�<"�\8#6�9�Y����|��M����}���=���(;>�'f����B2�(F�FU޽���U��J��ҦZ��v��v����z�����na���K��Q'n���&����V�п?F����ڙ���ݲ
�W%����f�OF���g���!��f��y�����t+��є�"=G�%)��u���桴�j�ab�q�G���=T��u`�K�����DX�ѭ�Ҋ��f�㵷{�������\��͂�\?LA�H�+(#�G/�>Kġ�Z3�k�[�W5�-�]]�X�9!��=�p]8(L��W�hE��GW��/P���`+�?:�yײ�d�b5��Tk�	J�M�o�DG�f'��5��ࠋi�C�t ��$�Yyݞ^�V��Wx̺W��y��r���w����墑�ATྥ$Y+��d�If���V��[�vF9q\z��[��Z�S�z��E����E'Y4T�+��`�G��t>��Pn�&�y�ԝ6v�?t�#�a�2ci�q����x�N���/�G��X�O�?n{�A	~j�^:'ޯ'�U��/��@*�`�c�;���*eC��
-�g)�}|���%z1�L@�b�iD��Bѵn�9ğ)���c�<���Sz�N�9���x�}�참?���4��'��ʬ�ǰ����@{T��\9�X$���{s}�+�$?&��V9
�\!v|�.T���w���4�~��{�v�OOk�U%F9�}�����26�˓��Ei�9�:dܸ	��0gVQ�|����'
˳Ӽ#�Nc6�9�+��aPq�^��r�+CGa_T��^��j�"����ؿG��xA�%/ֲ{e��y��a����Y�z<�����$mܱWF:�T���tu8�EL����B��V�F	�{$z����-R�Bλ�3p�	b��i�}�=nv�s;$�nEY̾��b���pPVfZ�^1�]��v��k�2-�����yƳ��}��^�6�3�t(좍s��=;[��-$�l8�f9��k6}ڻ+/��;]�ZV*��U~T��\�ڔ����VʙX$QjQ����鑹_8P������C��h�d`�s[/�U�*��A� d=B�-�p�^\=����n�N>��ߩͻʝ��7�<��ƾ��g�F����f%��G=��b�,Bt�5rP=�_�'%�
�ک����Z3�m��9q:1���1}
3�U�
����g����x�Bxj�bь�	���!��U�n(S���C���E�O޻��삚'�����_.�s�N�V&d���&�[T�hZ�@u�ʑOw���i/�pq:�KȅB��	�$\�%-�D�d;j���fv
8/�8�س��[b�Xl@%��X��};(^����]�:��~����cͫl	�n��u����@���k�S�N����J������)z�o�jªzVK�dT }��v�9��p4��"ldR����JqWs���w���r'�9��\��_<�t�D�sj��p���L��'�(��l����3ޡ�U�	����b�E!����y�9���k����/���x�͔�݅��f�.w_mvm��}��B����-Q����i+:w;��8w�|H�	*����+]V��,M���b{Q]�}@Z�5^�o/<��Knϑ���Q����G{$'@�	U\pZ���M�^}�X揖Iy��]*��80�>o�FO/P�> g���P�eo�ʽ�|�Fu��.�c��>��`�qR��DG�n�&�Z'���}�B�QT�/4�B7;q�qv��uѱb�R]�FءB�	�U8��Э�/�̨t��ꃆ)���l�+[��HA/��tp߹y�2���=C����U=A"<�X�5v(w����7SC�T�C�X�ƺ��O��z)���Y�p�p����2#+՛i,�ӗ��˄e���(��h��!w{U�
�d�:����}}�m�j��ݫ�r.�6X<g�xSO�"KF����U�IH]�[�WO_�yܬ*$0��O(��s���:�!E&�	�`�7����������e��m��۹nrG��Q��8�fpk�����Y�U7��Ȧf�$NNV����	��2�͊�˄Fx�&;MuJ�)꽬���妸�.�Щ�"�{�#6���?�rf�Wso8��=�]�aTyҮrj,�.V�95 r��[#�*N�s����ٵ7Dwgg͝�k3�����V��*�u���{|&��L�[gf�9�'�w�k튺��Ձ��3���U�GP��XI�N]R�ԕ��ڣ���WRu�5hm���6�;��/D�q�}�̰��M��T�p7�uφE+�{��rPV�T����Nl"<u�w<��zv�!���3���Z�2�*ȫ�QQ
��t"���W��1)��n�ǵ�Wp)�J_c+t��v�\������v2uA�)�s�J�[/��7���h��;S9Qr�XݗHVI([:�U�{A �v�-��oi[�d	�e=zU���ͭ��;�}6��T���ΐ��f�nX�d����?Tx@��� KRjR)B��x��Y��&��i$�+8̖�#�z(ޅ�0�U���J�^`�}y��X��� 5Y��ѻ���q�w�K�o������C:��t��!����,���\���wY�;�]b����.��YV�%أ�as�J�ru!�vE,��\+^��n靌R������Q�K<ޝ]-+f�uE��ǵqdi-��oi�Z�K��b>�jR� ����-���-��/���[�-S�h���&���-.��U�|�^�{)��IlN� ����z��:>7��'�j=���1]��W����p	)ӻ�'Dq'�O��gR��Έ�fZQq�x�fu,��wQ��m��ݸ��R�Z�p.(�[uk&�t�:����YC��AV�1fއtr��o����Y
�e	kg`��X�+�&��9��T��(.�ywj�Mv���:�����W�y��}��u�����\Del�vVhx�'yxE	���L�F�Y�Rs�f�@���V�Aɓ+1>�{K�X�9�w%8r��-�n��KL�j�s��i�e��uփ�y�U������R�֋���l�E��t�륓��ڙ19z\ܻ�`�޸ٛ���xV�.��la�M�?K��������؛�B�΀5u�,��҈�8�v�qR�
K��g��[���!� x�k806�%(ց�5�{�|�e,��rcˮ�=��Q�pli��N-,���ۯ�z^�d,uu^7k���n���$�IN���I����f���L.�������$��^H��u�ռ%�Q+E̸���9�������&"��B��KTr�V�"�kn\�S.8"�im�Qq�r�I�a��R�4F��Z+Kh1"(�mE��DJ��R��3-pZ�q�5�mS2Q�FTjT�5q���\�1�[3�PQH�ъ�[K-�P��`4���j8�̥��0֪9�ƈ��.X��֚e�#���˫�T�Ժ����-˃�0��-Lj�DiVQ�Dճ-Dk1�����*���Yf:�e�rPFT�کZ1�+mպlA�DX�����E�-�*�0�ur`�n�1b�CN�q�3�!�c�5qQ��)WC��(���5h�X���e�V�e�UM �Q��(c���]f�T���f�k�QJةiR�iƸ�sWL�X1���M%�5�KKk��`QE]aQM[Lr匶�3*�ڵ�c�f4���.��eȰ�B�b����h(��,��Ι/����P�T��+I�[n�lەg����kN/��ٝ9h2�e����ـ���tX�=I��u-�]�T�	�ј!@�&�h����R�B����_uj���if�e�p���=Z�������(xx@.^�QT����Uhr�=ܘ��s4�`4��ګ���fo)�S�s(�6f&���Q	��4�_�xR�Dx=��p���wd�ۻ�&W�kbOQR��^�B�%Φ�\|,�^�'^�Ag?ML��g�vBEp�r��(-��w��D�C0د:���������u	�-f�>��<}h����ݡR��:¤/�X�˾{�eō�d�8�ޛ�ꡃ��yv�R�tr�U^�$�w�mҋ��$#YK�T?.?Bg��x%[[B��xn���?nt��%��J�ڒo\^��K^��w��krD�Pq�5�{�0�T�c{��sfxE�:�L߇K�C����`do�5}��2(_L)�b���_V�[W��o,i�Y5��
�}4�g�HΧ�2
U�E��y5a�j*ݘr�S��o�tSݹ#�N�w��K�^̵�����\�Z274�l[��*a�z�B�)YK�'8�kx�+9<��y��^��l|a�E����go�gu��4��tQ�ȅu8����h�e�>��(^�:f}�V��L��&��s�$y��0��eΎ�<�mJEp�$V�K�1��t?���=�D�K��kW��tOk���W��������p�<<2s|",h�u�e��S�ˎ��䧇6�cw-eѻ�,)�Qc�T�k����V8�e��}��G�F.:U�UI���[���k���c�ې@ޥ�lEEЛB�@c�
%B,`\�����κJ�e;<��j�(Q��%��ñHۛܘȲ�ءe>Ѣ+�j�w�M�63��o1G�1¥xe(���\��n\dO����&�� �����(��r� b����U�'��u�@��|o�1R)��PA:�D�Tㅡ�D^�q=��%�=YG�B�>4�_b�b�Y�r�o���\	���;%�W��9�ž6Z�=];r���^z���T�8]	�ÞS��Lzb���W��a�`ʮ�wY��Ң5��`Q�=�"��fU53ĸAN츘��D]��nA���o��)�Q�ݢ�n#6�3����il�Dꭖ�²֎h
J�����7y����]qaGm��5�Ϯ�M�J��;MuH!]W�wXo]�����C])�uoa黈��z"wF��(��R�Z�0�b�D��Cܮ���{���zFFŵ�rN4F��i�8�2/nCr��I��%Gl��2�
�siÛ��jC��x���9a������N����yU�9ŧ�Uþku=N�8}B�=�_¯��[w��Ҵ�F���3�:��#7F�ƽJs��vغ
-Lq:8?Q��y�Z;�ϡ�NPh��=8�˖祕&\�~]��|}ォj�uqR�'JV��n�n�ʿm��z��ұu�<�3���Y����f����ut:��P�X�O%����(<�b�u����۾S�h��!�7��q�t�D�^!G�@��q'�;�3��K�W��y�7�~��;���|=yn�짷��d�E��[f�K�]@����X����M�$JU��օQ�����b�>�!�N<��Yq(�Q\�`������,H�0Ɖ�����5���qo:�N�u�7(^�{Y����^��&
�:�9-,�w�VgX����{bLY�`n�2W�j���g��]�]fw��/�^��n�l�������S]kF:U�o��ө�v�"�,Li���R�s�9
��,��c)�ȕ}ϝ%
��ӷw��{�Rՠ��xm��E/�r!a��FUB8�~��|�Q6�^ص��fx�ַ�N]��[ �`wP�� %Nd�Tî�0�%V򢝹Ƙ�\^q�cO,LFE��oh!�4� �VTIj�vE��쨘9-Ț�gEi�ŧ�֧E����MFs���� {mx!�{�	�j�O�k ����U�X��d��M��w�'�8����}�_"�ܱbE¯v?B�g�� ��D@B����"�h:���l�A��3�FǝM|0K~�N��Fe�As����Z���\f3B�r�%tE1[ғ�լ�M�a�-y16�D�R�o��5S��6h��h��ŷ�=G����\�����"�ϸ���<+c��De8s5��P�e�{]%�j���7��
��9���Br�Hvt(\W�Lp���$Z��d�}��ܪi$��Μ靇Δb��ʴ�(G�ѿ�Pᤌ�CMuߥ�*KhsU���Xjj�G.�F�Ya�� d 7��=�R��i���7���xp\\<2�Ս˽�w�*o�E�["5˧RX�6�oQo�ɈX�}5�醞�i�D:�ɓGw����%r��=���ٽڷA+��y� ��H�%�L�`SnH�CNq����s������s�]zCʋ.��N���Z��� �ly��~Ty䭺i���]�:J�*d��尭!��fgz	��;�>Cd鉆�t�R�aM�(	�t�z� ��s�@xV���bI�]�[hT?�q"���'�%���aD��:HQ@��DH��3-O��UD>ū9�_EE���~�PpM�N�>�B(p�@�Y3�|]K������ϼCDjK����&��z�	{��O�X��t'��������V�V�U��E��3j;7���m��]�)�*QJ�M/>�� �C���;��XGʼ*��tlz�]�h~�h=�,nOD��jE�$8��P�����bj���>j+"��C�L���m��k�
��s6�\�=�U�����-یɦ$�׫j�}�Q{Ml��T���r������38�|6͋f}�,���H_Ud8�U���N����q&Zwbf����R��\r�FiBd�g��}��;�W!4��a��ì����CȬ�B���ta��om�}��@7.pA�S��8F�ah�(�Cf:o����\��B�ŵqZ�of��Y-�r���"����h�K䠶�f׫ޅ�V�;��R�q��Ԥ�S@�v/p���p:�3�fI֛fͬ��P�T9>wj���Ԯv�Ȓ9
أ����"�7GaΠ2�;�;V�����]؀^�b6/z��ާݕ�'`l_��~���N#hQ��y]uË�ǉ.J��u��T��� ��k���\u��sZV����=�(�(�P�B�����pz��s����*�^z�C��߳�
�]*&r9;w�B��+6Kۺ^��p�Qޡ<"�*����RT\�D�\����s�9L�8�c^��7Zr.�JM:%װW[�{�MкGV/	���b�
���/����a��p�	�W��`墢�M��8��ʕV�`�[o	�uxOlpf3k��k��v�m8p�o�9z��R�Ld'94��L���FD���-�ںK{׷77L�A0�@,e(���dd���>n�J�a7��� �W@3�]�t�����w��9�gF�c�i�A���e����3S]ǯ���[��gJ�t1Ms�r/B+��Z�����]s��(F����ESp(�+.9Yu�:uuvm1�V�7k��7�	;�)f�wp�;!�ś�LA�,'����EM�2����`�q����j+�Q�'}.g���^Q�_m>�b�mtL4/��x:���>S+9��q{��hmJ�9���`��}��89�T�d�6'����1�ky��%���I�޴q�k&hy�al�m;ّa�̪jf7��(ݗS��E���m�O�e��/��h��P�ʲ\]�{B�#CZw$�B�b%�m�MX9��b��7���F���(O�16��nTl=�f��j��̲5ݢDmf�Ige��j�^�'����r�
��s'ށ�zO]�8��v2���U �n�=Y�ZSk���<6���X��txd�-y[iw���$�s=eU�>�:�%���n����
gܪ�H�m���tpߧ�<����B����'y�'׍�[K���B�B��{
�z���\*������O�-y�XͯT��I��OTt^��F�[�b�<�2:LK v������+{�(0Q�i��f��$�w��2����(��\����s���R��9=�UQ����k�ф�M�gJ�u[1�i�J�B�bp,SiT�"7���\�R�3�����߾y�7HL�ne���h}�,�fl�{��*� ?X3�ܢ�]e[\ЂM��ٞ�N�ˌ3�C��'*�������r4`}���OWB2_L����xX������{	��{��ԣ/|�U�JhWzlC�9��"G�W��VQ�N�#e��Z^tكa�/:�N��{��&�y����!�R١`��a�����h"��
������w����y��hm��K�k:Ԣ0E�bk�S��2�9/��Er�4R��fy��Ds��z�g=S=&�a1��1�� )�����*
�îҰ�ϑ�ce����h.۫��˃�Y$)�-N|,!�z���~Wx�o��������CE����%K����� �]A� �>�`�[�б>����3����E��m�fk+�,�=YG��1d2�#���b�>͠���u��8�H��8l�n^zS9��+�a�o��fʻ
���r�7�	�/�Ӵ/PL��W7�`.������]�S�fG�M<T��8q�F�,h]�n����ے�W�rv���7�=�%��V ������^��X1��m��M�r�jU����]�+X%��.��^�hH6�䣩V*� l�ᮤ��#�X�ִ�q�s��$��XmI�q#d��=寡���~��Uc>�Ci�{\�S8�^�+�<�zx������s��ls)S�ɬ����hZ�h.���]��'����oR5�����^>��(�S��_чs��AvCX����5�.La�c��$zlC���Gs�+_`t����j.��'�bP.��7�u�c|��x�eE���Sds5Ժ�|����9Vz�PIE'�CbD�腲��e+	E�yr's�AZ��v��m�)<�,X'�h��U�|�\�*�Q�o��9uL{v�o"�Z	��<�������c�q{t�UvGeg��	
�&Q6�L�<�8�Pl���ˉ���U�ZIԴ�E̼�ͼ���*� �/���w��dq 1�z:��k.��� ��Ϙ�J���wS���\�����X�e`*�^��m�t�et���RV+���xD��/u1%;��\��v:����w��sı0�I~�41D�G�WM�!��LMryq}���֕=*�����#-6��n��٬��Kc}���DỺ��\5�6�7{c�4��`J�d㡶��:��B����I��+څ��[��Hx�,%�H�#C9*��-�]դ�$_dƕ��GgCkM�Ozo8Y����ǁg��xy��9��t]I(�ep���Z(�=X���i�C3ip�OC�T͵���j*p9L�N4�tP�v�F9WK���pmK^l�Î�)5Y����"F�,B5g�����6��fС�Փ4�]�L���sI�jպR�ԫ|�x��k��o������O���OΕ����|-�������HHBO�%�IINMS�����-��,�_�Қ����G���f���	 O���!uMxkP�aAB�>ua���C��g��u��'p�Y/�?̟�) I!	��E�<���?����������?9�N}?��a�_�Q��H�՞�׾�,<��هq}?(P�l�yד^}$	$!?�M�����~�����$$����$�I!	��?Q"�ɇ�9��������̟��'�'�tS�_�{����S�O����@i���$�����[�l�����9�3�Od�C��0C��%;����Y��O�/X�/���[�����s�!�?�����M�ø���"O�?�;2HHB?t�C_e�:?�;�$������h!�zU	�d�����s?���<����tr9 I!	�NöB�����u�����y��&�C�����A��܇k�������k���?�%?�������;�ޟ��Y I!	��n� �����{����~�����vj��'���6�!?��_��?���~�������~��=��s�������C������HHB~�������"������:���P��'��,��	$���9?��$���)��"z��!��l��^��?�������?�v��BI!	�v~�U���Ƀ�h?�=��|�I$�#:):<'�~��:&�����,��$�ɐ;���-��tk�
	$!>�O����?���?Q I!������A��~�?S�?���>����6~p���	�	���0�5c���D0#����������!�������C_�����$�'��~]~��"�-(����`�i I!	d�n���f��h�������?�~�~�	�����NΡ���
_��X`�C$����������>|w�@�g���_����=�����~?�?�IO��'�ߺ~��#����;��?��>���s���)����~�����N�����)$$����$�ԉ�BO����O�~������HI!	�	����v�;���;�u�сי��Ύ������	���~��������)��x