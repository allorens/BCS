BZh91AY&SY\�S�:�ߔpyc����߰����  `����T(
   =>� �  uO�렊@R��D��Q-�TIPVتF
�qި=v��1���` �      ����}u�w����[�;Mz9vt�� g��ϣ|ե�;��w}�/l�5{t]��]۶5�!\� �@ {�m۹wcJ��sL�;����ܶ�j� 8>�����û����<��d�X�9ݺ�� s��� ��s�t�1�������Ϲ��w�y^��  ��Zw�=ǫ.���wap�{=;l�R �${� ���ݻ�k�g��ͽ�t�rn˻wax��۳�9�׺�}�s7|:;5�ۯ����P@ �o5�u�{×g�����/om��7�<޽o^��˾�����vŞ��m�  �       Q *� O 4�R��``L  FFC&�i�H��R#	�4�dр& 4�JcU44 �      ��*T&& ��` �4�$�BC!4��h�T�6��i��oS�jx�*(��������#L!��0 &i�~�$D�Id@dU$�I�$$�}c���B�~�x@ S@Z,�"����w0���E � )��������sqB�����Z��*� ��U-� ��䒂T����UQ0@NQ��$�@O�TQTQG�~a���0��	s$ْ�6~Bl��+|���U��o"�����5ө�	�Z�tG�=:n�:�Μ6u�8�0o�?`b`N�tc���,&�
"؋����jL&P~e����*����%��.��xSR��)����ŽJ�e�@X�41઒ŝ��t������nj�FuS@b\%P�B�&���XQ�r�vU6���C�^0.ÝI�+��2g�0�;0�%��c:0c8-�Q9$��b�0�`�4H��,B
0$�>��Ia���H�e,�h����֬l�Kz:!ՇF\W��]riɾ�g^/�[�ƺ��ưtN2kX,k$�{(��	�0�k�S�����G�2����:�5�$�!������`�H0��6&:�tS��eze,9�;�l��%V�a�cC1�Љ"Ĉ����v�cFh��0�hoـ��p��p0��Y,c1@�h=�B���1W@�@g��D���&H9��[�t��Mü�r���pN�'ER5ь3��m��4\2�K%: �MI�2!�����>�5��XҶtf2�
���Q�&��׺��i3�R3�%��)�L�q��'=��!�f@"�fC&�*�9�\��3DSCr$�{�~�$*&|`R �,cm��%�I!��FҚ9�gIΉӧW�z:��WW�;��A��(k�X��]Z{,�v���1�5d��&L�n��E[���K�C���.C�H4,�&�$��ɸ�&�?i�4��Ұ��3T�ӂ��.˓��A~�$�/B��S:RӚ[46�V�Չ]2NݤjI3fhՋ��1RgIt�s'pҴ����j.RU�p�����L3���ZR�+
Ri�L��6ay��:L�E�FIbQXX�;�g(�����Ta�N�N��ɆZe+,(%�Gl�(R�қ0)�|Y2:L�*Ѭ�S�����4ʦfR�)TUX���d�A2t�ԡY9D�/IzV�-���0M��D�Ix^��[*��ef�sd�^�[�Ŕ4�K)2��XR��4��فL�p�&�"����қ27��gq��w0��o
xu�Z�&	d�8Mf�Ē�BxSd�kȴ�RN(��(�үiu%
,2:IĒ����h��`����ef��Va�/1&K�+l��D:8&����O�!��2b!�u��F-�-��-��I<Ej-��:�L�;RK���di-�V"�$�IXnJ�^^�X�i�L��S��7EY/J�+[/5�Y8ZԷM�ҳA���z^���n�v�{G�a�����N"�%��.;'JZsK�I���6wN��%#�I�3�7f؋,[�*q�`gS50��:o����n�(>x�{�8N���,4rS'%�Ce���t�IE�����KdS*��eM�������l�XRuAK5$�xE�A�M�l���U��1�F�)�p[$S4�&i%*��E
,Q���	����ZmbYd��l��e��.$�$Y"�/	Kgt[9'F3vn�Q{em�p���4K)2��XR���f�ٚe4l�&�M�K�{�S��Mg�e]��+0�xV�&	�Y:N��a�YJl�mjY��I8��zUiɌX�cXݸ�� Xͻ���ec/4�g�,e��-zV�c$�Z$�Q$i �$�.�x�z�m �KJd�D�*���x^��I���i��I6��[EXL���'!�����I�+Q�Ej,7i)��d�d�*hԴn�K&p��ke�9����-�Ҳ�#�804i'Cf���
�t�
�T ���Q�v2-1ŕo�֞%��իnFr�rP�I�m-�R8�X�f�,݆r2�\��`��)�CC���6d҈Ґvh86p�06X�Xb�bِ�R�ԩ�LE4���EjHK2QRh����>l�FIB��(Hv\j8,4Xh�Ɇ2����� �I1�^s@Ι"�!�vU١�I�E��d�$�L��%�m*�R�^,cIPh������b(�E!>a�B�!���2���D ���v�N����f^��-��ʡ�A(c$����'F��&�f�	aA��i���_��2J"��!р��ؐ��IQ��~�pX�,k��]@-�p: �hS���!���e�_�ђb �`Ptd@tX�ie=)��J���a�bޥOJ�Ŵ��@��h;���R5RMQ^~��~d$�	�S$�Ҩe!q����V�Ɗc]�ݕ^bl�����|��N�:���	}�����gv��$c80c#�# ��LD��m0_�+���p��K�u7�^v׹��lkcxE� 1g	������aICA�>�!��y���Ӟ�X	���B��eC�����O�K�v=��~,$��I �8�nfٷ�!���n]��L�A��.
�W�F,^$t�y6����:��zZ����q9�p_����8}{���$�K�fe<kI�$Q��∧�� ��!���&A='�1�/��fC�JC{������5\=�o��]1�%��9�OI/7od��� >�@�d< ���;�e:wd��KL�8B�/d�Ov��w��HS��8h��ݐ邍pT�4��q��>�$q�/�?�(ٳ�4I�jn�%l��"��G�"v �I�E�t�B��ǇېN�ۊ_Oo��`3}�hy'
Q�g��tu�aǣ%��܋7i3��(yP]�ؽ����0��/�,���T�I�J<3�4��o�ON�\>U�)��$f���{���%o'�=���9)Iy�t߬� ,�=��5�Ν7��.��n��H��?YϤ=9� �`~ߥΚ���O���i��N�gǄFI��_ӿ����4��&����e���_�Ӧ.��צ�uϲ��q'���~����_RW��fl�x?7|�|��� �f. ��~�����e����.�z2��2Cӄ0���:t�H�<3��ڼ��ȓ����͓� �?~���p� ~�0�ొ���� =4fN�aE��Vn&���Z��~:hZG�1ªR���_���L��c��ŝ�b�EfN%y�9Q]��6.I6}�i��B:f�"~1eIrQw,�y���xBA���R��*��œ�}��w����4��� p�,��b�?�fI(��I�jMtU#�G���o�����;���w�(s�$�'���:z:?
MM���ޏ�10�!��~��4�����~����z� ��&.�9��IȈ�g�G���~;��8�'wa*f���U�t��bqf��r���7l�xwhh�\�5���XxBJ~�?I�Ӈ�O:�!�:|t������[)D�.��/7��(�&	��>S�Ҧ�ڗ��ڍ(���eK!�CF~�i:,�|�t�ݞ��FI'I��"zm���l�8��t�e�1'A�e�&��g--DudQ��D�e<4e:B�_Jzp�<=!�B��)��ӧN�NJx�����'�݌�y�w�wgM8B�G{��\`3�n�|��J|b��<ߦ��g��#�>���}N=��{df�G�'���6\�9ѽ�7J3��q���S��/�)Ã��~]���0?T��}�o ���{�D��W&��9��ӡ��<<��.���gw�h�ؘ҉���wNMŜ�����q��`Pp��[���b�"�*&� ٓG��ׇ��CO_ t}]��NàW{T,g���0�����{9�i`�e�we�$�Q�0Y���;�ie��K$|��8}GN�$ы��B�⦩L�I�*�1N�I�zi�Ej}=�!����k<��� ��J�� )D��qGk#o6n�\l�>��0~�i{�hi��� �i���6���^��q�����dd���F�#[��ia�מ9��4 t�v�?�*��w����K�(t�qYG�$ ��\RS�������zA�Ń�{`�=YË �FtƑabyL�c �J:t��3'L���wT��Ȁ�9{潷|8����4ջ�=�g�L�{o�9����p�:HxxR�M<�<yŒI��fH�,s6bc-ʘ���=윜�+�1g�<<^+4����Ɯ,�f�FK�rt���f�'���ӕT�0tȳ�g�f�t�!�'�$�TJ,�wv'$Ś���:IdU/"!U�RK������US݃Ʒ6��e���'Ja��:g���d�8w"�#b�͓�pX��;OM<ݐ� �WpQx���U�9vQ�Z1��w��|�λ��u^���ڷ��Y����<�wF|p��/��=�~:e���
2jpY�R7m�QW$�M0u�1��p�15um����D��O0��g~�̫�h�%L�$�7f!���!O�JhO=T<Z�V|�U�f���R>���"�"j����!ӂP��M'$�H�`w���_�g���rU�l��Q<|6������������ޕCOl�F�i�"���ӛ�d1i϶D�=?Y��e?����t��I��L���O�<1w��|�~��t�}�AJ�\K|�@�_s��X��(�5#�h����s:gɮ�7�]���hZ�������2����|��+�b��v���>Ay��!�����~N8j��*�A/7�M��q�b]3JiD����z|~1e�m�W�_&���0��	cZT���o�/��V'�	E�O{����tؐ�˦)���]�7�mO&�5�t��B�.���wc;W1�Q&��E�;.O��$k�:\ֿ�*SL��j095���t�Z��5�j܁�͉ջ�9�L�Ƌ����O����R���XI�����ɥ  ϶[�)@��h43o[tb�E
6�h�)�+RUr�k}#Hs�@��`��a��$�+��X���x|�hl���G^�o!EA�^Y[7g�Nb��Z�w ��gЏ.�ֻ[�\:C{�Y3(��`F�n@ܺ�!��q�4Q�Lgv�>nw9�HJ���U���Q���"����/��! �4C�w*�s̩Y1���޼�/N�#�v<u4��P�5��a7j�W7a��CPm�JVj�aT^��iN6d�<R���ږkSk��X�TU*���)ƍc%�"����}�IZLh�����j�
MB�7e��IR�eN��1A��!w��&R921(!!Y�Q-1��*!εED�US5%���[�--	.��Չ�/�YRVt�bc1Z2�p� y(�A���Z�	�C����A��*�����0v!��.J-��mQ��N����lJu���[�=a���o�(^5u:���G��0!�ÙwzL�d�Q�!YJZ���Y�e��E[��W54�N5ט���$����ڶ�_?��Y������PG���'��_ ��A����@�|�~��A�����J|H?g����+_���cf��.��0�M�wUT���m�m�M��m�l��m���oYm�e����m����Ս��6[m����m�m6�t�r�m�M�,��r�z�6�6��g��"^Q� �PE$I  @m����Ѻ�t�L7���ꪛoYm���ܶۦ�m��0�m����m��m�wv�w\�ۦ�m��0�m���۶�0�m�m�a�ܶ�v[m�m�� {� ���<TBE*
�E$BD�+�YY��[m�nm��uuUM��6�m�i�ۦۖۆ�n�-��z�m����m����[���m�m�m�m��m�a��oM��opm������{��}�{�戒�C4�����wr��x�usm�{6�6ꮪ�m�e��m��m�m�m�M�-��ݶ�6�v�M���^�m�m�m�M�-��ݶ[m��-��m��m�ݶ��m�n2@���O��$�  �<r�����p�o^&�n[���m�m��m�a����m�ݶ�ܶۦ�r�n�m�m������oYm�ݶ�ܶۦ�m��0�p�m�!��m�{4�m��< ��ʃ�'{�g���w��}�{������tꪥ�m�m�m�m��m�a��oP�mݶ��vۆ�n�{���1���m�޲�m�m�m�m�L6ۖ�t��p�o^&�m����R���䨩h|O�����B$�?���?���� >ϐP|C�+�_��o�O�x�'m��2�
�N�:��2��^��6����FOJ�ӧN��]u�]q�]x�]z��UӧN�u[6mU�M�î��:u㮲�׎:ʺt���Ya֝u�[u�x�׬:��m����]z��u�]z��^+n�ˬ�ºy�1��O��{2>�Y�N���)\�]T�7�X�C��Q�XF!	�GfQ�$uH9��D6&�6�rX��L*A!��"�C� t�^�WW�b�֚��؜�^�-[v ���ZR6����+,@���c*�w
�@#��j��§AQ@Q�^֪�-�t\��2�떩[�ku��3rd�Dj:�.B�JWGcx݊'aUV4�q�H�l�󵍊�9D�ڒ��6m׶�@��G�Z���FJ���&ES�i�n!+��@	�q�� �,l������N2���̃����5	l��e�eR�M9,2F�Ӣ��E2����aE(���,$btbpBt�c�%DrT갣U�m�n(Eq�Ъ��R"�9���"�U,VF���\����le���9��57בN���ޕ����(�p�c�J��M�C��vV�ɯZ
7	OZ{�8�ح�Ue�M��d�厺8:Z��F�'X+()k���ʙPF�j�-DfH"�6�N�퓛)�dkT�<m�D�T�����4�H�@"��1\*E	cp�*iS˻��ص��芚hN��qZR(�e�	�˻mRH�D���CFX�b��)P�R��V��RJ�ʜ��
�ʛ��V(V��x;B`ױ�[�i�����$�aq�uH܅p�����d�"�A�Hڤ��}�X�幪����E2���D䪻[rA5�RV�TЫq7F�8��Q�k��k����]��DЁz�f�[�V:�J('$2�Z�eUV������r3m�G�'+d�(�aq�)$�d%+�RZ�&�Eq�W[��p��f�#v��.I0�R6�HH��j�kv�7I���2Iu�R'�2�m�f�RG��

� �i�J���N�dNES�2�ڨ�	ǅ$h�fj�JE���htx�B�h��T4�c�N&dmT��nٍ
����!d���lq:�i�nd'��b6UYem�G1�DJ�������ZV��T�"�j�dl�(�����G���U\R"V¨X�v"8�D�MZ�U���l�(+�i����&�]
�]��e��&*��c��NZ�E��%��6J�	0m��$����lqM�jm80���C-��6&�l�j`4��]�A�5
E��Oc�nF�WDݍIb�C�$+c#V)�Pdb�c��qƓ��7jr��D`��Al!J��HEm�&�m)5	 a���l
��DUمN
��X�mMʐF캚SZ�QܭZ(�B�
&�:�w���MŢ��UUuT�4Ц1&Q5e+��1�m��juEQ��WK�;�7dIYT��!�]��Ƥ�TZ�nBiBܪPBFH4ЛVRH�����6��II�"��Q	8�U�����;ƪ��ȡI�1����[#j�<d��` QQ0��0���33=������%<OwwL��ao����S��wt�����xx䣉��陙����	Dr=��33<3�{�	Dr=��33<3�������p���UV�����AP�畢�۪'�nl��~�H:�d�)[�)���ۈU�t����h���6�j�FABrKN]ӖTB�L�(]�UUq����T�&⒄�U���ؚт+r�u
[P����VQ��"��chL��jF�"X��e�(Epجn�![[���$E�R
���n0e�2V�6<���-��9 �f�c��CcM�`��*
B�� ��<)S*��tV*�B�+�EI��d�bmP�,_%� 2Y�թrFK�K�b-�H#r�pR%�j)U"����!M(��"]#g&-�P�4�S�������-�f��T���WpQ�\ދ���f]��5F��ĝ�$���d�+F���ӎ��i�6!$f��;����ܐX5��l`�8 @���miVY����X�n15V�7F�O<IG(�9����}�$��,�H*ă0��Ơ�`�ʚ�Dd�!�Q��Ѣ�⧪8B�H!b"f�Ym��I���I ���7��w$�q�bI�]jR�]���Q)w-�j�!�c�R��T��v��g~��W>��\>�9�A
��;�ƑecC����a�f�0a�Unyj��Ղ�q<ߵ|�}�䴒����8��3�"H���`~�|�4����#�7M]]BU�+]�5j4�K:]є�n��4�"Y5i	q6����Q�$�2h�y;x�y����P(KH��+̨���7uNc$���<O�o�.�p5,��+����G%p-h��P��VDƈ�¨�aLu�8��1Z5S$ˊ�D4B
�,�TҪ)*Z�Li������$ad���$�!bm�9�Վs��6H^3-���a��!BnŚl�4bV�T�*��gQ�`3�ae�I�i6B5
���pW���0Ÿ���ȱt��U�Y��l8@�4���.�l+T�kb���y-ӗ�!��+\��Q�5jɪ0w��ܻlam��_LQ����Sq��V�2v�}����`�B�2[d�e��)��gOA��}2*����1���E�w[��ݯ�D���=D����LS9Y���G�о�� �-*��U9�f�_|�7���^�����+w��+Bj�j��En���,�e��Qe�����,�4��/��%6<�lBbk�!,�`Yh�|Wqn|��eŸ�F���>��9�Ͻހx�w�mW���6�,�<mX+D��=_zE�o�h�خ�J]�oFN���9�����'�NvZ>G�R�-��ǰ�Qؤ�
ƥU�U��a(�Pڨ���K��!Z��AZ�t��d�Le�H�*vU*�+��"�R�J�N�@8��l�!��t�b��_�1��4���ukZn��kt�F�=�ɴT(4��i�R@Iѹețm1
��d$P�,AēU�1D�r��泜FBl��,�!�"@H%�2g#$�`p�jU;)0p�pܱZ�D�'�lMѿb�yƅze�� �(��zūmK�ъF�1I3���F^ uLnRn�ٺl��Q��rf<;	`�	q!�xph�7������>�$����� ��<0��|�>7D��#^��QȈآx�����x���x�	��h�����>�ǈ|'G��x#��+�G��t(�Dt"h�Z�dО0C��2>���	�:C�t|<���"xQ�+�G�<8Õ����'����d<<<O'��Hx�2r.̓c���'�N����t|t�v�<��h�>�|Y �(������}�X�>��^�������vg�g?O/�����_7��wv�8�wLյ�vp�%Q��]лJ�7�-/�����7w9L�h},� �0�~� r����33���IA�{��ffxgw{�DG���fg�wp	Dû��fg�ww�Q���陙�����꩙���Ɔ�-8�0ʴaƕ��իV��*��e���[mVC�E$F,��@ܥ���ljHIFX�h l����R�)IN-m�{'7.�8�ꬑRL-��LI�l؅r�$�-��Tތ&ƍ��N�h$�" :4C���E���]3I�'e'b����e���8HA,����]��!x���EQ@<4Jh�Te�Zn��#��!H��	��-;�ԑ��UDuaE��݉�5�C�SD՚L�n��̡�{n.���򺱷B^+�.��5|g)�#�.�V�s0������BX�|(S�LG���δ�-qX2�MT�⯡ǟ��[��%tZ�۬Оpnr$o.�ZX�f�,� X��`�FT��(W!#R��i�r�r(�dq��,M�De�Ж�3-VR�N�%M��dMd#j�iF�~����0YR��!G��	���[=�_ׂ^0K�M�sxI%&Se.�>�s��x����H'% �"<"���czŹ�r�L�x�8E�<A2�}����˔�+t�b�"��JV��J�|���2�Zw���`��.(kر�c~oY'�mQ����>efa�B@�	d0Л�.�y�*ba1{�������(�V@A�d�)�#r�6l��Q�+ġ,,A�ى�ˍm����!������/t,N�]Ď�v�YV**-ة�T�&Z�V�U����c &J7G�I9)�y�`&�6aF�b�4|5mؙ&۱�ac����$�	#ӃE�]IFj�JI�9d��b��2�OD\��g�/#S��n)֞<e���8�A,�1>r�ֱJ(��Q�i�n���(0bF��y�W]�a40w}�n:�Mș`�bƨ�x������c�^.�Ep@�W�fT��f�-����J1��z����ݚ��̥/	�Z4\�zD�Np�C�7��� �&�U�U��tA	s�h�,\8�K!����w%�x�]DQFD��v�oRI�����ԑا��������˹��Ęe�IeB�
�P�!h8
8�U����E�{���n�|D�*)�	�c45�bi�UwŌ�vQu���c�0P&�m�.�lF��%*݂��w-&F>b;cxcX)2�i2U1�*�&�i-�6*m�C��Ŝx��Yhh<hHA,���ϤΌ^�4wu���~.3y���$.�H�q,]�i�a�6%	X�)��`�LLT����Q#-�溔1��We	�m
m+�5A
�J\�Jn��Dd.�|�I��a�[G�ib�׮7i�M^D�a:�}�X	��G��!.�ǵ��~�EO0�nfc�����LG�#@]#�섄(p[�3�QZ�>��j�EWVg�7��=���]���,k�QX���g#l$��"���z�l���l���L��#���m�[8~qX2�$!��GLc��H���f$̋V�KضK]WtS����țH�2Z��/*���|�Q0DJ#�ɫ#b)Q8���wU7]�x��G~[k�䣖6��_�14ǰk%��7K$M0W��}Yb�1�F�"���~ά��{�A,�6Dl}�4 ^�`�2#҇�|^Q$��٨�MY�c��a�G8��Xa�.<���I�3f~\���I�31�a��Q�F"i���I15ܕUP�93I⒃1��o4z��	Th�f��b]܊Yr]����s��r�B�l��2��0D���zFC����FA)":��7�_����g}�\lh�Y3
`�&���p�0oU���=�ѡ-ٺ�|�]�)�<d��M	,��Y���[�Ri��%�P�H�#�	�ˆ*b����$��B>CR�(K"
1�J�t�,S�\�#|��7$,��r���8M%Sn5�R"i�d�h>�!JZM�,�6�CQ�F�gYHI�����bLr��I�:��쐖'�i/�:M&���Hd����d884O������$����YB�<(��y<H'�G�c��D�T|"n-#���<(�|0r"6(�k�K'�G�'�!<'����	���<'���[:OD���Q�z���Wįh~!6";6B��d؟��r?x�zC��Iᮏ��dl�<(�Q=J�U��Á���|O.��d���<'��I�����������<r;!����l�<x�G�I��M�&��`SŖx�A�d�Nő�BI����d>{z�A�Yv�"'Rz6��8`�,U�E�ub��T`ʨ�Q�$�B�q�o]�+�.k��/��QC0�(�W8s*|��;kګ�s��m�ȉ�1�UE��IQR�ṼRz'�m�=�xH��������mב����d��Ua�$(
��S�K��������	��+լDQ�Y2&\ɜ(�x�P�l�`�d'J�'����}O�:3}�U3������ʪ������ʪ���(�û�����s�S<;��*���>p����϶�b@�8X! DQ4�J./����@ �Q�k��\Lm�	"�DNB�-2�f8�["j (�j�Ge��\����A\RG$��&��#����@�tƪ�i���T�[$m8�E��VD�j�T�Ƅ·[��\���A�
�(�V�ʝ�V H��15$v�I�'\
�2A�X��У��.���vCGG�K�;�+h������U�#Tl�W�R;y*`ԮEͫwa��&�p�I%(��BEL����t��G\r�&
�0O+w�L�5G\�'R[+D&�h��ѕ<�#
�+�'j.<�Kr�U�A9=)G�-r�aY��i��uݖ��kE�6����lx��	�:�f��;eU�k�Y�$B~+uFh���:�"nS����9^��& �Q�[�$$�Og��w#G�os3n�5;c�)�ś��1P���{v������("&,4��\?O4��V*���]-��b���ͤ���0��X�&��rљ��8���6q�`���q߱�l��]�
4�T��,]���G���2	2��O{у!߄�b���2q����o^�8��=�H��l�v�oz�\�*��a.�hM%�n���Y�B���8K�����rx �>�ǘ��̠^�#���S	r�J�I��4�)�`���K �c�M��6í��qX+,��F\{瘆�,��jג_�1j�%�&$|bB�&�J�񤧏���3�y� ݄ɑ��������3�����{�D�u&n�Q���k��5��0��cL�)�oʙ�Is�S�iL�w��w۞���
lh�M	,��Y�_5�}C�/0L`�b���ۊ��q0�L?B�#���Zb�^��� ���$��+�f��@9X2Mت|�|��Cj����a�e���HȘ)�(�K!���%��C=l/���GCk4#᷵U%�i�4k�Ը-$�&2�&��g^nX仆���na�辿<a�������4e���s��ڨb�ܡ[l�5��i��Ɔ�@�btэh7	�	Uc�� ƫ�`�1�,�IF�B�"�Ģ�X�	%�U���S���}��/sUU�u[Jn]��^3��m��@��.z�����ŀ�b]=��'�Y�@.�X�(�D�`'�������%̥���Ĭ���Y%��)�azi�4��C[qE�`n�S�SO(���#J.v`�����B@K,�0��\��k�m��ԫ_��e�Z�QMM�L^LL��Q�M�Q�XwV�>"�0��ub�@#E�:v�Vm�CIs���îf@�`����d:�d�r�i�.+�÷�(=�IT�V�L��-���;��)[�t��M��J����-�Y*�_9v~a��y6�.�t��XVMq�_2���%Nժ�̑�`Yt3�ᆋ��@t�MP��1EF����a��U*�j'pYc�i�5F����'I����� y�����_ŌF�b�r�A]��%� X�>������-=ʛ�4x8���]�-�.�ǇF۸�m���͞8��dї>��P��i�q&��e��-��j�R�K�v�X�p�Zތ�1�� v1�C�E���U)Z\��[Ob (�̒S�pq�p'��Ԓ{O2P��2j�k��O����e���̼fb\�J�61<jr9��4�Î�B�T����ڕճ_��l�7�"n��Q4H���X�9ɩ�C�"�"`�Z���"����R���eQ�r�qث��mDHu9$r
�Q�T���+JBK,��.���b�p� ��ђC�
�m�����R�vI#j]3�2���~��R�Dl�_J}ZᣔY�~��ZO��� �&G�b�)��;�I'�ƫ��h�@��Mꀆ�r�6�����28��dїM߭�X��z��'k$��jb���5�^]�n�{Bu��n�Q uY���q�	�S\�*�T�g6N+>�cn}�c�հj$ic�)�U���8�=�+��2:^'�����ݜ�N8̂�Z���z�CC�DѸ�ݿg���	����A�Q��|'��Ðk��<Y�}��D���|(�>0Q<(�¯�&	���Á��L�%xvx�������p|l�|��Q<(�U�+�hEt|Yb&�[;2C���?	��Wó�<'�������á��N��I�F�O_<&�xtl��'��	���:O	��K��t�&��	����G��G�:>:N���hpx��e��Y��q���8ϧ0�&.d�A:Ҡ�+M0,���^�G��-��׍첓�:T�gI��#I26�9��!�߮�"KE�R���Woni�gx�pLZ+ƧeW\�L� bK�|��Y�.�.�3�xR�"	ي���DV��(����vD�4��/j��:��,f|�����s�V���9UUß"�����ʪ����wwNUUp�ȭ<;��r���>Ei���������w�]z�֎8��e�R��~�ܶ�.�d�Q���V��죛�̍?oS����N=��6=���WK_gB�\�ܑ��K�:uﲖ"@&^&-x͡8�x���*n��x;�Mw��Uf�L\��r�Wۢ��M�8z�}��]t���XVZUe�:���4x��I.�-�v�X�n`�a���Xٞl9�������$\)!q�m�3�;՟�g���m�^q毿m�5E��?6\�e�Q)��6t��j��1�]�B�D�]ٓH��q���$���l��Ϫ�{n.1w��d{��g8�GV
²Ҫ����R�&%ج+�tQ��ı�OJ8�Z�tǎJ�N:JWKdj���5#ly"�E,0r8V��F��+Z����c���յ[�6�eփ�&>�g�S�&���
��d�h����&��,k���j�-�frssr�<܄��L��徨8�clR��r�kWmmƚ�&Z8��,����?|!9����r@-�Ӧ�&\��<Y��ѡ $��h���
R��j�V"�F���Tj�[�ʅ�"5ah͐e�:G��DvPu,�19^ܖ�I��̦O���5��x��וujA����S�1H5jv¹F�m�c��#Q��X3��4'��rG�o[���P�_��,Q�^.5wBX�[�':ܠ�1���6�[�3ܝ�MQ�|�޲����d����f�t���lOyɻy�W����9;�H�b7o���Ԑ�S���$fT驚��wXk�V�����	�Wf�dFdؚ���E��X��0;��~Ef
�n�� ����u[�d�9��aÀ\�N�P�2�c�$!��1ɔ�?q��׆��Zo�ڑ�9n�ki����k����6ٳ�Ղ���Ue�49��eS��̾^�@��M��@z�n�d儦h�&�̣�@�z�j��I{�@'��:�rP�V�Q�b> j�byWLr���$$�L6�4�ƥ�����-����i�O&=ۛ`;��� ��f(O��A,��f�\��d^V��6;�Vȭ��b��`<������ܿ-ԗ�\_��26x�e�R�2(��0b��zl���r��Cc���)�-����c�pq/�� K�,��`��۾֌&8�i��.S�&�n���:��i���l��LϞG�����u�����j
x3}�Nn�?��S��^r��� �%%Ou�6�	T���R;U�nIe$�X�Jdm�Z���U�QQ��Zʑ+.6���V9m�0�؞D�(81��l��4Y�<P�,�zNt�����0����N��$�)���m:n\�d��F4X�VBq��F[�psCr�TPK�W%I{T��']��N��"��J���<���Hݖ_�EU+Yuz���(�B�}d��.�����&Ͷ��u�V\z�w^�#��1qSCάK�g�Z�T�Y��.˲Y��� ��� �m�od0���K�}4�4��{;�_m�{Vw4v���jj0�le1$W�ˊ>���Ե����$p�)@a(���r�2ԕ=}����>z٣�Ղ��,Ѽg�v6�̙"B�(��o����EDf(�}B�bX��6p��2],�Q������we��.�r(K�l�a� õʅר�F��G�דBf9����M�JG|m���Og&�8��"��8��6�	��1�-��c�1&N��g��uEi���`�+��m��X�ՏH@��9p�^S���w}��i:�tX8�%�w�ѝ��ޮ`�Zƨ�e<P�2����m.�&[�8ll��x�`&�����v;=G����&��Œ���O���Y�>���|8'E^G�H�E��JG��|(�������C�xp>	��<&���'�pO���
>|(�D|(�káUҿ�7�lO���|&��|<��<=<C�l�����ТX��+�W��6x�<M�d��x�:=2OG�t�6b.W������v6O!��|N�'G�Ӥ���9&���<66|��#�����+L�j��>-����~��9����U�Sw�m����̫�ԧ�J8Jvr�.܁�����n�kL��� �C��sPW���|*�i}Q˨�zsf��ěєT����2*j�$2#+�B�V�T�K�\��ۘ�;|"x�z�+1	�R1;

�s7,%l+��@���O�*��
53!1\��n)U��W�\9@
V��;n����*��>%���wT�Up�����S�Uû�X{�wuNUW�Ia�=��9U\;�%���wT�Up�(Yӭ�a]iU�Iٷ�][X-��ds=�թ�U+�\U��[AV�;�j��B�&�#-p�m�v�DW"���+)*�� -��A�j#cTV��8�"$W�yY"cn6ے�I`�962k�k�&뱺�[������B��mcPmR�K)Sc"j���٭[e��ȥ�ǃDu��1T�ۮ�R��d�*�U�̪�W\�8��[%��BR
Q�JJ��\qYSMѦ�C(�h�ݴԪ�ۤ+
R�;jȅw%��\h�!J�B�6d2��%T�	�L�ET��,Wct֣�t���$v�M5lT�-Pm���K������A�(B�0j���Ռ�.(Y��_h����x��H��|lU���H3b������ቇ�T�͙2����k�p*�hъ���g[�.]�������-s)��b1n&���Q��=>mX+
�.7�~o�*�r�|Q�y}d�],�R4\��M�2Y+G6m6��Of�pr�M'e]X����_P�f��L��I+�ȓ���<&$�d�u9G�Z�/�����wF7B�+��ʘ=��jB˻���R�~>6x0 B	��f�`�<}Zn]�a7���{��3n��(g�J�Ѭ{�L���8S��<���dmMC�%Z��y��\���2�࿉ Q+m�W�Z��kP�d�|�L��L�N�X�i5C�^!������S<�5F#���8���V�p��l �h��fn�-cf(ٟª��ɒ�W��V���Z�DH�dg��K%�,����j�G i)Js��J�7��
���i�G�!�0]9t:��=������Gv�(�����C�s^�x�'�ǺB��t�,������:�W2�	�� ����+qt�"�E�!ˈ�I�iDEz�URٿ�զ�{�Z�s�,{6�4!ͨ�h�؜ye݄b�*4Imk�-�.(!��H�Uq�-4@�CVI���t�}�ɶ��RO����̽���'2�1���8-�7�O)G�8Quu��g ��l��K�X�-#�H_-��6ဳT�.7�\"jN���j{�i��h��9�P��"��2zm�0��Ze�}Y}�;�c��yE꯰0����b�#%9=��
a��}�T�'��,�7�۝\����Ïc:֛���VL	���_�ƫM�Y�ZM��!��ށd�d��+���Wr٠�;�W��ڷ<��IOWo\�zUZ�Z�l�[4X`6d�&�H`ѽ�i㫫E��C��՚֠��Vq$���^ �0�.a���|�0�.ƞYh__�@g˥R1�e�n�i�㉙%ٝQ�1F���oa��Ͼc$�k!f��n�jU����[.�ܩĊ�	5If��Ø0�
jG�Wm}�q��Ʀ����)�Lpc�L���\7y$�oN�&���G,(!��R@:}E���f1r^1<4l5CVr���x���,gF1�4U��:���X���;��C,��r�*��2p&��#�>	���`&�ə�o-LqV�ٽ�<1�7c��ٛ��I	'��b7[�|yѻ�;���7i���j�^=d���0�HX����	�ˉ�pTk8D堯)g�o�ݫ��kj�����I[��� �TuZ�Ce�G)-�J�[����n7 ����*ܴ�����0Uԅ`�����vX�ɉ�)��I�ѳ�Lt�dp��Y*I	�t�e;:��)f�z]��>27�S)AQ�Y�g�m��cJ/d��k4�g�c��d�V�HJ#(�i�牽y8�H^�d�����/βl�la]Ua�g�o+�,��V.�%��)>���Wo'22���{I�õ�ˣ���s�m�SD)8�����l��{ٷj��cuH2U\r����^fLP��c�-fG)���令�A�ٜz��N|�Ɓ��ȣ��d���GD騸<L��D|Y!�"x
>�	c���|'�!���ti8A�F	�:(���:(���ª|(�">â�^��Bd�	�<'��tM'�"A�Q��G�����DG�DК|J�p?�h�����	���C�2<,�|��|BA��+�^<OM�,��8M'HO!�:`�{3��6O;l'���u|N�'G��6z>6\5���>���0}^u܍)���8��}A����>?.y�NR��	"
�<�@Ⱥ�Ca�x�	���FE���ׯg�ZFT
|d��^Bq��D.��ɋ�5AD]�E��`W�[R*�#I|w��NUWû�X{�wuT�W�IY����S�\;�%g��wUNUp��;�wuT�W�J㻗wUNUp���A:"CG�������NQ�?���	��)xm.�u��u%w�I;��.��3��떙䵚����LF��9q���mz�����g.*���М����s�:��켜���Jk-����4a/}\��_.2��Qㅁ@1A �` �,<���)��2�b�+&��4���d�7������c��0�1HȀ�&(�l����w�Z�ä��,M%�xB\�i�L�!�&zMg6î�zH�o��l��)���SZ�=t]}�,�*�=m�+�VW�hQ�_|�8��.��M����mq�k}I+x�h��ɮW���Um���I\�C�9��0�	]J:J�@Z����$ݮ���7��DQJ��Eu4A6��6��K|3�h��;s�-����1�}d��]���2V����\���sAtoy���!&k(_����j�͢���d;f��ZI�T	����b�UT#(���j���l�4��	��CFH�pD��ϙ	6���\/��@�f�p�0�K&Z�aD�@pФO�B��b�H�����U�ޙ䧔��@G�B�<��kJ�'����̒e�d:�9��GqT���?�?�%�����j2��q��׆�!I�:��'��m�1��M���>���G��`����|"CU����MfŌj���cw8��i��S��76n8���ϳ�kF�j
2A'�b��w=��w<�}�����N�[l��{�	O<d�~�7l[�5��f�m�Y��'�nh�2�0zHB�S`{ƴff<�MI�c�l�������$4&�֦��ŗ��vl��W�_���a.��{P�,X�(i��鹘���ܶoy�2�>)�S=��Ii��I�r�͈I	���V��l;��ɇ)s$]bO<�ͥwG	��"tD����^.�֊�G���ۥ`�6>�@\+mċ�Ir���d8����I��m��#�J֝j�Z#�D�)S�$N�!k��
R�ٌb�B��56��SHt�ס�HK�H�-õM�'�ŗ��[�v�v����l�Y!$d���(���!����ip��ْ&�oO-M��7Ԡ�T�"��P~¤����T`��Iv<�To5a�d�US��8�xA2&�Hh<b�8�.2�y��ɣ����f5�цJ�y�����]{�+���}X�����R}���!1[��+��t}��FH)�7��g�ÄL.�n�BUU�Zpt�K*f7��m~��q���M)�)�4"CD9أ�e��.q��|ѽg��@>{����$�A��ۿYJ,�;K��&X�o�!�õ{h��S˳%�oͲ��p�th�5�>�S���]zJ2@�ܕ(�Cx\�DGs�;B�J F��p�I��q�. `6 �B$4O�S`�(:#��	ƍ����~2���馤UY"�����6Q�i�$����;��X)���K��h�Q���<�ӏ�%��B���ZҤ�d2�#��^�J�P��A�Q��A��Y6>8N��騸>&�b��,�<D|	�G��xa�x|0|>��Q���Tz"'E�'D$z"5�'�d���|'�&��d|'�Hh����ا�|?E�	�Q�
�%'�\�&DG'�46|C�0?�����"�5���C���|(�i�(�U�įxl�<9<p���x�2<<D���5fɣ�<z/�c��>:O	��:x�&�E���a0x�>�1<I�4iL��M8�����$%!wr$��/ [�T8�޾�n�������\UsūY���r����E'�wY�F���H�k0��`��"�X�b�$����­.� ��t!�>*�A/�Kn�Y3Y��R�H�[�.�J^m�W�I�PĤ��zs���x6�;"���=�"NEJ��ۛ��W��꼯�E��@��0�
*jCB����S�\;�+]���UYUø����U9\;�*]���3�9r�K��:fb��ʗwtv����x�g��+j�4��������%��.LV)*�E��kؘ�ERb��r�D�"��V;u��*m�UZq[QG�E�E FGS�ɌhO(㭖�([��إ�UV����v�:[�Z �F�iʭNalr��E%MЎ:W!�D�@�FT<��eC,�v�탊��m�N��Lr���LR�k�!�v���,���N5B4��)��JӢ"�T���ɗwv�hv4�!�9���Bc N���v�r��DA$q�T��v�U�7Q�T�ZeoĒ�Б�94��UEcv����dRJ�U�,2ESd��YdN(V&宖K���-Q1�,�j�i��/&��2P��{-�'�X8a�c[2��UW��m�S��n�x�yj��C��D����d|ĳ9���w�c%�Uˢ�zx�N��?=�0uM�R������j9co��nm��pb�����t��;�����5���!��4�\�w<]˚����dQ��q=��UN2��^�"y.�N@��4�՛�i�c���>�[i�ߣn6��6hA2&�Hh��s�9��sm��.M�=o$�E�#��`u�c,M�r;%�	u�x�Y3����Mm�u��m���`�Z7��U�)�I�J,�s$�1w�n�3�%͸:���9�W>SG����8��Ӈ�y�V�F$�,�ؗ���V��2j��z�����Ey�E$!"�i5X�V�G%|v�n���>C)W�N��t�b�P����V,�+�~�o&������ڎq��U$�/&��R��h铂V�B	�K��/;P�8Q�N���rr��!\����h�z�&:�ڒG��ITm��H�0e��p��H�m2W"�8ڒ�14�ZYЅZb�H�������գ���oi��d��!&�q�6r&�'/t��6z��A�k-%�%K0�Tp��oՕ�T����"8H�Wy�x%����c�����ww�p�8/VO5���lꉪ3���T�ꕵ8Ï�N$�~�e���si-�A	P�;1��l��0��9��v�C�w��L��mN]���9����Q�儱�T[N�B\�{v��L��e�h��ܐ�Gt�j����)�v�d��ːt &D4CE�x�r*�����U`_H6j����`U;���|B�$�	�<�x�!Z��7�z2ȪŴ\�K$���Q!�(4�i���h��YH��A��W<"�P����V]��^Z'�����8��K�w�e�o$��d��yhժ0d�$(W�U��n�F�-����d�#E����܊�2�,MUa9U���Dm\�����"��m^{mh�I�JV�Xf�ɣj�9E�����x����xf�]���b�%���in��eե��(�,��$��c���`b��C(��4��b��%F43!�tI�=	Ȃ6-����6�@�bu0BLNYDr�����%��m�Զ j������X�QON�i�6������$\D#¯$�Ŭ�8.�4�u��+�<T�╵8Î]� 2Hx��5=�$W0J �#ȀTP����DMD]EKż1-�V�@/*�֞�Y����#�3����	�����K!m�B\n�q�|W+���\�)8M�wI���6��#�ǌHC�o[��v��L�lZA��>�UT�fܚ�i��M2��8|�mN0��q��qL��%�Z�['�3UT+{
�T�+�T�e�A�J�S$��KB�5q���[k"�(T5q�l�6�N
Z�l#x7^�4w�_h�ıHj�d3�k��ŭn�.�9$��si�VXy0�,{���/��ܶi����^�<.��hֻ��e4�2֗�S�h�圛f<�c�l?8ڦΩ[S���=?vJIv�x�7&&�_� �,��5edSㄑ����L�ģ풽F(��bv��$E"�:�.�k��5ܩzdY�J�����X�:�O��6�:�.?<q�o[e�.�WN���:u�Xu���U�����������*��U�\u���׎��׍�����
��lі������5�����]x۬��N�N��:�.�ӯu׍<u׮�ˍ�ۮ��u��u�]z���m�Y:º'�!�7��aā�J�֪$T+��!mm�YLb�m���N�k	KJCj���)�(ir��Q���D�1	(��h���Tb�\��3�s��}�S)Zq�[�/�iS��hF������Pu���+M�5��q �Zh��R�GϹ(�.ؔ|�Z�f��	E��B����E���i>�kML��_~�,�K��1xaS�����*�Z�H>�ċ5�t����9��|;�*]���3�;�*]��337�;�*]��337�;�*]��337�:9r����33}í�ǏN�[S�9>�3�6i>6K��`���'���D��E�)s@Jȭj�"D��iT�I�]u$VJ�(�.�&�ɒ���J�(��Qs	�����㔒��i��S~��3/�m���+j��1��V�ˋ�I�z����1Fh�]Q!��+��OAm.��vˢ��{$�<�x��lnX�>O8+;�@�(�:�Jr](<G>��R���l\�C0���d2���޴c4�*������2����R���0�0�*���iz32'�HB��"����Y�=�#V[l�*�u �R���R:�p"�EF�M�L��(�U��0�J�*�ݰX�4�֜'Se�:�2ݽR](�D��.��\뇎�$�S	�<ʏ��ݛ�������mK����@2�Y�~����ZkwK�p�m\q���V�U�g^o;�'�D�L[ia�.jm�R]݌4kp�ܞ^��ǈ�(v���51H,)Z���������5T<}Ϙ�	g��o�?g��c�>��B�P3�LJ%�m�c�Ƴ]����F#%:�T�e�G���-;��-:7�zӍ��)[UWq�ͳ�sXkǄ�v�ǖ;d�W��l�ƉZ,5Fhh�,�JR��\�-A
�,���$l���d!�bI�)��ۼ4g��h��O�I!{�Jh��4�.Bb;:ˍ�R���0���a�a����U�L�����@.�.�<�Lc(�Պ�)�Ѭ�a��cH�]��%٦<}�L����CVr�,�Ƥ�/
r`0���o�)�������lƣQ���llꕵSZB�X���2�8+�L	J4����*�T��'�Ng����
-{���hR�)l���#�Eeh����ܛ���`IG�+��$jD�ǜF��^�;��)d�ߋ�#&�mU4P[ˋr��S��g�=~ܣo�+�~������.��h<>m��)mQ[#)�qL_l�W���xY�=|�oT����8��.w2�l|�|�MW�ҽ�t�6�6�M�ŭ�:I�����K$N��Ѧ�y�lc��l�<������R'�ɇI0���;ts�2I4�\S�夺�4h""h��8�z��M����w�U*�ܳb�2G�ܷ�K7\7Gh�i���>ݪ4�,����ǟ/1u~ũ�乽��rYm���ΙN��B��u��4V�M���;��^:����+j��0}"�V*���_֭�%�8仯&�8w����E�w�s�(��P���L�N堈S�l`��nL�ۑL���گ8�������5��T4}J#P�5�^�G���$�l�}9O����x|��ج�|i�:ӎ�q�޶��]a]a]:eӧ]u��:��/Nzzzp�z||t�]W]u����u㮽u�n���:u�W]W�8i�|����>q�篘|�׎:ʺt�:0C0���2t1�d���,m��u�x�]e�]z��6� 0�0ܱaH
�Ȉ�^�qV�FU�^Tjr�ڡB�(�X�-���.�4���^�.�K���/��n.E¸�V�P��R�ē�l!\^A���M��+Ө�oƻ���s��X�{�F�7 MMM�f�;��&��?��Ϡm"���&���N��WVL�B�@5VLZ�6cj�*j�U�f`�`G�|�7������WwwL��g�zOwwL��g�zOwwL��g�zOwwL��g�zOwwL��g�� 0 @�����uz��v2���J11��m�-v��Z�U<��J��A���AE�t������8�-q�ڭ!&+*���`9!lc�d��rc���nX�d�_	�n�cs�UZ4D ��`�)$�\h�:ӐQ�8R�D�R�S+���6��du��kʝ�a\���m;G$j2�� ��Aѧ�r�A�Zio--Dv6Z�N�&���u;���F�*g.�Iqn�\���E`�`���%���7H�&J�u�v��m&0S2�*�+h��uR+b	�[��mN&!���ڊ&G��ϒɏF����N��ȫ�����V�*Ƣn q�H��5#Q�"�����xd��CC$rH�`�V0mg3;���%�90�BIw�n���%Id�t�#�ζS�1�66G��>	�����j6Bh�$��Qr���1dvϷ5=���V��a�n�R���J2zx�8=oq4��Y�/��:��$��W�Z�F���n4f�D8bU�,����EXo�n�Y�L���g��,�4]58�}cQ�^:�d4 �D4b�bmX&B���p�]�	Äb^�wv�$�`zEي�����mG�����T�%jش�$���v��a�hÃ�n���b���䐅���\t�o2ӯme��8��╵Uq���
��RB��gzM%�q�e�N�ɮG�K��K�ѭ�����fy���ר�s ���Bf_�4b�E���0]l彸�L�4�� m:RWݮ<4�vNG��Z��U��8�mTE�#o����y�гN+�3:'$<|>K9w/@po����6 �X��)\��UU���#�2�KS�l�������*�H���,n8�Q�6�c.�<��W¢.��)f��wi�h����ܒ��M3��c	��n��r�)Ӛ���V���_���%�4�p����)�i�W�/�UU����:�mP�J7�dď�eT*��iIsN��SM�h�����Ry*wf�i�n���,k�u��Yuӵ���%]�[M���"#v@��:h�p�t��)���f�����j�X�b��,�d,���+j��r��e�Y��3s)�;����,�r�4��_	۱5��i�i���v�KH;1�P�W��L!a�s���T��I���O8~R�췷8����㻤޵d�A��-��#�ںg�S[�GjƋ;�o����2��46z�mU\a���0�CPNm*���l�p�vR�,�R�W(�	�Qq�RY%�/p���s\��m���0�c�����}����8���	�	�)Ӊ���kZ�iib��Kb�VM>�a���Ep�F́��A2"&�Y�v���u>�y�M�9=?q'̓8g;��Ⱥ/i$z�J�@Ƅ�U�D�	Yc��A��	Z��
��q�;`�����:5T�'"1Ǌ� �RD�	q���j3򸻑s���I&���I����\�LrI2a2�,����SGK�`�/g)N��#��KjIH��DM�9�u�3G�ut{���j�h��L0���ꕵUd��i�d�]$e1��84�}tݜQtd��/}f���vd�G.�Gr�~�c�u�SS5w5}�\W����s���F��*�n��������I�-k��w����*Q*s'�wGgq���Z��b=a]?Wzӎ�x������XWXWN�:۬:�-:u�ǭ+����2��:u�����:㮼u׮�m�UӧN�h��Wm_>|��Ϝ|���:�㏙W�ON����uzӭ�z��㮽u�e���u�Zu�]z�׮�x�n�����z�c4�M��&p7K^��j;v/Nf�ʛ��s�T���T��R�2�\Z}��ϻ�"㼒��J�/���w7jP�L��mh@d�DlL�C.�Km���y������33�������33�������33�������33�������33���0 �	`� L���wY
����'�G\���;Y4ztt��5��K����k"h&�*-e����7qy��7;��L��$J��ԝz��g����I�AŸ�?.��k�Vj�Jڪ�yj�LL'�Og����d�k��<�
����y���K�,�ՒQRz'L�!c8�s `h��~��B�!����e�ü�6��g�rR���K���S)�吆D�	�4K��}r�"� 35:���1@�Z�gR�cWl�܂!dUZ+���ʙ`����m���J�i��v����dcDI�l��-UTx�ED��'+M���HQ�*��l���!U�k��(��1����d�%����a<�����q�ޓ�zX��gǚ.��:/�w1�?/:w"#Ȁm��$r$ؗ(�<�t`�|��H�|Y����+j��D�,�o���;ZXW(�?wfI[.�F)����*iU_#P>���CR�V���3w9٪D<L5X=~Ff�Q��|ڂ��g�\d����Į��4r���z�����	�&o�P;���l�d4 �L����^2��Z��+��C`�l��@�f��ç$�`Kn��*7r�#��EМ���{��>�lr�>���tŒ�7�*��đ��txޫd2B��.B��ӐnD�`Y�ƞ������YJhLq�$�)��ն�[S����>оl�K,�w�O9��m8�7,�)��%��7�ˣls&Ι!L������/�,��~���P�{�3��wSkĳxU�*r�Km���)+��(��YZ++���'db+q�Z���ƋT�r��.AW�n���m@��?b��R7��bBq�Q�S&
�!�B=�y�a�&ݑ:��*�{$��Uc|��ş]�z��}�D��"��A��Z���W�%�!C����/&�Q(P�hѓ�N%ӌJܰBI4�&0S���)5Eq��%�&ss�>�6�VzJ�e6��RC[�4W&8襑8�μ��G�1|,>1}��7��=&d�ɕQ�a�0`�J��?�����鷞����wTt�j�4�x�q��UJ��	��G4s�0���/�������be�y�vq�d��QO��dx��2l�UV�v��W3w-A ��RkK��a�0b�vD����+��B�#�qS�]]�G��Э��<�x�u�f	SWuv咸N��c.S������ؒ$"I�I$�HQUD���~����q���@���~�bB"��"�DX08�Ƿ�S�k��J�U*�R�Q���4�R,&�0E�R()JE
EH�Y$�PT���ARPT��RX�IPRXE$��E�(��i�QPQPQAE�QHQHQbJ,IE�Xb�bI(�QD��E���Qa(�E����f��E�����������
,�QfU�5#%J,�QRX��E�J,
*IF�I%�,IE�(�
,IE�(�(�Y$�
FXX�EAEEE�J*B����TEI(�%AEHQIT�$Qd����
?�H��Q`��VU�
�`b�%��A��#Ă��M YE�YE�Z,P�$�E�,��,Qe(����Z,QeP��)%�X��,Qh�B�b���)E��T�E�,Qh�I-
(�E�,��Qb�)%�(ZQeRK(�E�Z,Qe(YE�Ie(��(�E�,Qe(��X��,Qe
�YE�YE�9��RK(X��,QeKQEQe$��(�E�,��(��)%�,�b�(��(�E�QHX��Qb�(�E�,��K(�E�X��(��%Qb�T�eQb�*X�eK)Q,T���K*T�b��*��,��,Qe(��(��)%�,QeQb�(��QI,Qe(��YE�,��Xb�0�,��,�eQe)
�Z,P�X�ʖPX�b�J�*YR�K*X���X�eJ*X��X��,��%��K)E,���K�K(�(��R�,R�,���I,R�(��X���K)b�YJ)eR�,R�ȥ��J��YK)b�K)e�K��)e*��3��R�,R�R�$���J(��R�Ib��QJX����Ib�EE�AT�R�R�(�K)h��R�K(�Qb��ie�*�(�1�K��*�)b�K�K�I,���K)T�X�ņjCR�,R�b�)T�EK%)T�E�U,R��)QE�Y)b���R,UUJ��U*�X�JTUU�X�%,T��J�X���YUR,�U�QVJX��*�EU�Ub�KQ,R��,R�KKK%Tb�X��HR*IH�B�AH�Đ�RT%�R,B��1!H���JE"�d�"�H�
E�R+4"�(ʓ��R,�R,��T��d���H�%"�
EI)G��;�f���+���Ƅ�2R����>lTI	E�D@a	�#�W�'��5����7��g�����#������c�>������������?�=��p2�֐�>[��(d�/����~2��O�ڽ���X�Ͻ?����t>?/�.����UD�A��������`?�A�(~�A@?�@��UD�(S,���'��_���}�h��Hd�1(R��A?��� �>����!�>�� ����Ϙ���h�O�	 a++C��>�?ո�R�f'�L��������5��i�k��u�&�|����T��+�K.�ı2��m�~��,J"��bDd�ՂH��IB��E���'�m I /�~�
hi��V��jm��{
�{��?I����*-@!�
�KERD���&		$�UB-D �����?��L����������'�?A��8 �0�����8:�?�}�_��HU��hT��_�_ϟ�?�8��������:��t;�������߸��>����`(�?�|BK��>��?����'�4~��������g���o��_a��p���a�����  
\�a����|��+�����Vr?�&����q����)n�O�Q@0�k�#�6$�~��z%��$`))��<��#i60�d7q��J!�	M� �c�Y��ch��'���-�M��!ت�%)�y�H�?���}K��
�'���!�DR~d�_�_��C�?����·�8|���>��'9�ڧ�?�>Ф�G��~N��`~Ԉ�����w����N��UQ>E!�G����b�PTM�`?�h�������	�?�>��� ۑ�e\��
BᏰn\�˖,-��V��`~�/��}���ۺ`K~S?�lq�;� ��e?��H����Q�'�>���)C`�~V�v��������/�@��d�`R�����4�����T@���S� C���������A@>A�K�C�~��K���f�O���rO���~"�*�,��߂k����w$S�	�;�